* SPICE3 file created from singleRail.ext - technology: scmos
*
* drain/source ordering enforced by hand
*

.subckt NAND2X1_LOC a_36_24# Y VSS VDD A B
X0 a_36_24# A VSS VSS NMOS_MAGIC ad=0.6p pd=4.6u as=1p ps=5u w=2u l=0.2u
X1 Y B a_36_24# VSS NMOS_MAGIC ad=1p pd=5u as=0p ps=0u w=2u l=0.2u
X2 Y B VDD VDD PMOS_MAGIC ad=2p pd=10u as=1.2p ps=5.2u w=2u l=0.2u
X3 Y A VDD VDD PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=2u l=0.2u
C0 B Y 0.10fF
C1 Y a_36_24# 0.01fF
C2 VDD A 0.20fF
C3 VDD B 0.27fF
C4 A B 0.22fF
C5 VDD Y 0.57fF
C6 A Y 0.08fF
C7 Y VSS 0.20fF
C8 B VSS 0.19fF
C9 A VSS 0.30fF
C10 VDD VSS 1.73fF
.ends

.subckt INVX1_LOC Y VSS VDD A
X0 Y A VSS VSS NMOS_MAGIC ad=0.5p pd=3u as=0.5p ps=3u w=1u l=0.2u
X1 Y A VDD VDD PMOS_MAGIC ad=1p pd=5u as=1p ps=5u w=2u l=0.2u
C0 VDD A 0.20fF
C1 VDD Y 0.39fF
C2 A Y 0.08fF
C3 Y VSS 0.07fF
C4 A VSS 0.37fF
C5 VDD VSS 1.52fF
.ends 

.subckt AES_SBOX INPUT_0 INPUT_1 INPUT_2 INPUT_3 INPUT_4 INPUT_5 INPUT_6 INPUT_7
+ GATE_222 GATE_366 GATE_479 GATE_579 GATE_662 GATE_741 GATE_811 GATE_865 VDD VSS

XNAND2X1_LOC_580 NAND2X1_LOC_580/a_36_24# GATE_579 VSS VDD INVX1_LOC_452/Y INVX1_LOC_453/Y
+ NAND2X1_LOC
XNAND2X1_LOC_591 NAND2X1_LOC_591/a_36_24# NAND2X1_LOC_591/Y VSS VDD INVX1_LOC_69/Y
+ NAND2X1_LOC_591/B NAND2X1_LOC
XINVX1_LOC_402 INVX1_LOC_402/Y VSS VDD INVX1_LOC_402/A INVX1_LOC
XINVX1_LOC_413 INVX1_LOC_413/Y VSS VDD INVX1_LOC_413/A INVX1_LOC
XINVX1_LOC_468 INVX1_LOC_468/Y VSS VDD INVX1_LOC_468/A INVX1_LOC
XINVX1_LOC_446 INVX1_LOC_446/Y VSS VDD INVX1_LOC_446/A INVX1_LOC
XINVX1_LOC_424 INVX1_LOC_424/Y VSS VDD INVX1_LOC_424/A INVX1_LOC
XINVX1_LOC_457 INVX1_LOC_457/Y VSS VDD INVX1_LOC_47/Y INVX1_LOC
XINVX1_LOC_435 INVX1_LOC_435/Y VSS VDD INVX1_LOC_435/A INVX1_LOC
XINVX1_LOC_479 INVX1_LOC_479/Y VSS VDD INVX1_LOC_479/A INVX1_LOC
XINVX1_LOC_221 INVX1_LOC_221/Y VSS VDD INVX1_LOC_20/Y INVX1_LOC
XINVX1_LOC_232 INVX1_LOC_232/Y VSS VDD INVX1_LOC_26/Y INVX1_LOC
XINVX1_LOC_243 INVX1_LOC_245/A VSS VDD INVX1_LOC_243/A INVX1_LOC
XINVX1_LOC_210 INVX1_LOC_210/Y VSS VDD INVX1_LOC_210/A INVX1_LOC
XNAND2X1_LOC_10 NAND2X1_LOC_10/a_36_24# INVX1_LOC_17/A VSS VDD INVX1_LOC_12/Y INVX1_LOC_66/A
+ NAND2X1_LOC
XNAND2X1_LOC_43 NAND2X1_LOC_43/a_36_24# NAND2X1_LOC_43/Y VSS VDD INVX1_LOC_31/Y INVX1_LOC_49/Y
+ NAND2X1_LOC
XNAND2X1_LOC_21 NAND2X1_LOC_21/a_36_24# INVX1_LOC_29/A VSS VDD INPUT_4 INVX1_LOC_30/Y
+ NAND2X1_LOC
XNAND2X1_LOC_32 NAND2X1_LOC_32/a_36_24# NAND2X1_LOC_32/Y VSS VDD INVX1_LOC_87/A INVX1_LOC_41/Y
+ NAND2X1_LOC
XINVX1_LOC_276 INVX1_LOC_276/Y VSS VDD INVX1_LOC_276/A INVX1_LOC
XINVX1_LOC_265 INVX1_LOC_265/Y VSS VDD INVX1_LOC_74/Y INVX1_LOC
XINVX1_LOC_287 INVX1_LOC_287/Y VSS VDD INVX1_LOC_287/A INVX1_LOC
XINVX1_LOC_298 INVX1_LOC_298/Y VSS VDD INVX1_LOC_298/A INVX1_LOC
XINVX1_LOC_254 INVX1_LOC_254/Y VSS VDD INVX1_LOC_254/A INVX1_LOC
XNAND2X1_LOC_54 NAND2X1_LOC_54/a_36_24# INVX1_LOC_61/A VSS VDD INPUT_0 INPUT_1
+ NAND2X1_LOC
XNAND2X1_LOC_98 NAND2X1_LOC_98/a_36_24# INVX1_LOC_95/A VSS VDD NAND2X1_LOC_93/Y NAND2X1_LOC_98/B
+ NAND2X1_LOC
XNAND2X1_LOC_76 NAND2X1_LOC_76/a_36_24# INVX1_LOC_77/A VSS VDD NAND2X1_LOC_76/A NAND2X1_LOC_76/B
+ NAND2X1_LOC
XNAND2X1_LOC_65 NAND2X1_LOC_65/a_36_24# NAND2X1_LOC_65/Y VSS VDD INVX1_LOC_68/Y INVX1_LOC_69/Y
+ NAND2X1_LOC
XNAND2X1_LOC_87 NAND2X1_LOC_87/a_36_24# NAND2X1_LOC_88/B VSS VDD INVX1_LOC_87/Y INVX1_LOC_88/Y
+ NAND2X1_LOC
XNAND2X1_LOC_409 NAND2X1_LOC_409/a_36_24# NAND2X1_LOC_409/Y VSS VDD INVX1_LOC_335/Y
+ INVX1_LOC_333/Y NAND2X1_LOC
XNAND2X1_LOC_217 NAND2X1_LOC_217/a_36_24# INVX1_LOC_193/A VSS VDD INVX1_LOC_116/Y
+ INVX1_LOC_128/Y NAND2X1_LOC
XNAND2X1_LOC_228 NAND2X1_LOC_228/a_36_24# INVX1_LOC_202/A VSS VDD NAND2X1_LOC_7/Y
+ NAND2X1_LOC_52/Y NAND2X1_LOC
XNAND2X1_LOC_239 NAND2X1_LOC_239/a_36_24# NAND2X1_LOC_242/A VSS VDD INVX1_LOC_58/Y
+ INVX1_LOC_99/Y NAND2X1_LOC
XNAND2X1_LOC_206 NAND2X1_LOC_206/a_36_24# INVX1_LOC_182/A VSS VDD INVX1_LOC_177/Y
+ INVX1_LOC_178/Y NAND2X1_LOC
XNAND2X1_LOC_740 NAND2X1_LOC_740/a_36_24# INVX1_LOC_583/A VSS VDD INVX1_LOC_581/Y
+ INVX1_LOC_582/Y NAND2X1_LOC
XNAND2X1_LOC_784 NAND2X1_LOC_784/a_36_24# INVX1_LOC_614/A VSS VDD INVX1_LOC_605/Y
+ INVX1_LOC_607/Y NAND2X1_LOC
XNAND2X1_LOC_795 NAND2X1_LOC_795/a_36_24# INVX1_LOC_625/A VSS VDD INVX1_LOC_615/Y
+ INVX1_LOC_616/Y NAND2X1_LOC
XNAND2X1_LOC_762 NAND2X1_LOC_762/a_36_24# INVX1_LOC_595/A VSS VDD INPUT_6 INVX1_LOC_18/Y
+ NAND2X1_LOC
XNAND2X1_LOC_773 NAND2X1_LOC_773/a_36_24# INVX1_LOC_601/A VSS VDD NAND2X1_LOC_773/A
+ INVX1_LOC_600/Y NAND2X1_LOC
XNAND2X1_LOC_751 NAND2X1_LOC_751/a_36_24# NAND2X1_LOC_789/B VSS VDD INVX1_LOC_6/Y
+ NAND2X1_LOC_750/Y NAND2X1_LOC
XINVX1_LOC_6 INVX1_LOC_6/Y VSS VDD INVX1_LOC_6/A INVX1_LOC
XINVX1_LOC_606 INVX1_LOC_606/Y VSS VDD INVX1_LOC_212/Y INVX1_LOC
XINVX1_LOC_617 INVX1_LOC_617/Y VSS VDD INVX1_LOC_617/A INVX1_LOC
XINVX1_LOC_639 INVX1_LOC_639/Y VSS VDD INVX1_LOC_639/A INVX1_LOC
XINVX1_LOC_628 INVX1_LOC_628/Y VSS VDD INVX1_LOC_628/A INVX1_LOC
XNAND2X1_LOC_570 NAND2X1_LOC_570/a_36_24# INVX1_LOC_444/A VSS VDD INVX1_LOC_436/Y
+ INVX1_LOC_437/Y NAND2X1_LOC
XNAND2X1_LOC_592 NAND2X1_LOC_592/a_36_24# INVX1_LOC_459/A VSS VDD NAND2X1_LOC_832/A
+ NAND2X1_LOC_592/B NAND2X1_LOC
XNAND2X1_LOC_581 NAND2X1_LOC_581/a_36_24# INVX1_LOC_454/A VSS VDD INPUT_6 INVX1_LOC_3/Y
+ NAND2X1_LOC
XINVX1_LOC_403 INVX1_LOC_403/Y VSS VDD INPUT_0 INVX1_LOC
XINVX1_LOC_414 INVX1_LOC_414/Y VSS VDD INVX1_LOC_414/A INVX1_LOC
XINVX1_LOC_425 INVX1_LOC_425/Y VSS VDD INVX1_LOC_425/A INVX1_LOC
XINVX1_LOC_436 INVX1_LOC_436/Y VSS VDD INVX1_LOC_436/A INVX1_LOC
XINVX1_LOC_469 INVX1_LOC_469/Y VSS VDD INVX1_LOC_469/A INVX1_LOC
XINVX1_LOC_447 INVX1_LOC_447/Y VSS VDD INVX1_LOC_447/A INVX1_LOC
XINVX1_LOC_458 INVX1_LOC_458/Y VSS VDD INVX1_LOC_99/Y INVX1_LOC
XINVX1_LOC_277 INVX1_LOC_277/Y VSS VDD INVX1_LOC_277/A INVX1_LOC
XINVX1_LOC_222 INVX1_LOC_222/Y VSS VDD INVX1_LOC_145/Y INVX1_LOC
XINVX1_LOC_244 INVX1_LOC_244/Y VSS VDD INVX1_LOC_17/Y INVX1_LOC
XINVX1_LOC_200 INVX1_LOC_200/Y VSS VDD INPUT_1 INVX1_LOC
XINVX1_LOC_255 INVX1_LOC_255/Y VSS VDD INVX1_LOC_255/A INVX1_LOC
XINVX1_LOC_233 INVX1_LOC_233/Y VSS VDD INVX1_LOC_45/Y INVX1_LOC
XINVX1_LOC_266 INVX1_LOC_266/Y VSS VDD INVX1_LOC_266/A INVX1_LOC
XINVX1_LOC_211 INVX1_LOC_211/Y VSS VDD INVX1_LOC_211/A INVX1_LOC
XNAND2X1_LOC_77 NAND2X1_LOC_77/a_36_24# INVX1_LOC_78/A VSS VDD INVX1_LOC_21/Y INVX1_LOC_92/A
+ NAND2X1_LOC
XNAND2X1_LOC_55 NAND2X1_LOC_55/a_36_24# INVX1_LOC_62/A VSS VDD INVX1_LOC_9/Y INVX1_LOC_92/A
+ NAND2X1_LOC
XNAND2X1_LOC_66 NAND2X1_LOC_66/a_36_24# NAND2X1_LOC_66/Y VSS VDD INVX1_LOC_70/Y INVX1_LOC_71/Y
+ NAND2X1_LOC
XNAND2X1_LOC_11 NAND2X1_LOC_11/a_36_24# INVX1_LOC_18/A VSS VDD INVX1_LOC_19/Y INPUT_5
+ NAND2X1_LOC
XNAND2X1_LOC_44 NAND2X1_LOC_44/a_36_24# INVX1_LOC_50/A VSS VDD INVX1_LOC_25/Y INVX1_LOC_40/Y
+ NAND2X1_LOC
XNAND2X1_LOC_22 NAND2X1_LOC_22/a_36_24# INVX1_LOC_31/A VSS VDD INVX1_LOC_1/Y INVX1_LOC_29/Y
+ NAND2X1_LOC
XNAND2X1_LOC_33 NAND2X1_LOC_33/a_36_24# INVX1_LOC_42/A VSS VDD NAND2X1_LOC_20/Y NAND2X1_LOC_24/Y
+ NAND2X1_LOC
XINVX1_LOC_288 INVX1_LOC_288/Y VSS VDD INVX1_LOC_288/A INVX1_LOC
XINVX1_LOC_299 INVX1_LOC_299/Y VSS VDD INVX1_LOC_299/A INVX1_LOC
XNAND2X1_LOC_99 NAND2X1_LOC_99/a_36_24# INVX1_LOC_96/A VSS VDD INVX1_LOC_94/Y INVX1_LOC_95/Y
+ NAND2X1_LOC
XNAND2X1_LOC_88 NAND2X1_LOC_88/a_36_24# NAND2X1_LOC_88/Y VSS VDD INVX1_LOC_6/Y NAND2X1_LOC_88/B
+ NAND2X1_LOC
XNAND2X1_LOC_218 NAND2X1_LOC_218/a_36_24# INVX1_LOC_194/A VSS VDD INVX1_LOC_192/Y
+ INVX1_LOC_193/Y NAND2X1_LOC
XNAND2X1_LOC_229 NAND2X1_LOC_229/a_36_24# NAND2X1_LOC_231/A VSS VDD INVX1_LOC_20/Y
+ INVX1_LOC_32/Y NAND2X1_LOC
XNAND2X1_LOC_207 NAND2X1_LOC_207/a_36_24# INVX1_LOC_183/A VSS VDD INVX1_LOC_175/Y
+ INVX1_LOC_176/Y NAND2X1_LOC
XNAND2X1_LOC_796 NAND2X1_LOC_796/a_36_24# INVX1_LOC_626/A VSS VDD INVX1_LOC_613/Y
+ INVX1_LOC_614/Y NAND2X1_LOC
XNAND2X1_LOC_730 NAND2X1_LOC_730/a_36_24# INVX1_LOC_573/A VSS VDD INVX1_LOC_571/Y
+ INVX1_LOC_572/Y NAND2X1_LOC
XNAND2X1_LOC_741 NAND2X1_LOC_741/a_36_24# INVX1_LOC_584/A VSS VDD INVX1_LOC_579/Y
+ INVX1_LOC_580/Y NAND2X1_LOC
XNAND2X1_LOC_752 NAND2X1_LOC_752/a_36_24# INVX1_LOC_587/A VSS VDD INPUT_5 INVX1_LOC_55/Y
+ NAND2X1_LOC
XNAND2X1_LOC_774 NAND2X1_LOC_774/a_36_24# INVX1_LOC_602/A VSS VDD INVX1_LOC_599/Y
+ INVX1_LOC_601/Y NAND2X1_LOC
XNAND2X1_LOC_785 NAND2X1_LOC_785/a_36_24# INVX1_LOC_615/A VSS VDD INVX1_LOC_603/Y
+ INVX1_LOC_604/Y NAND2X1_LOC
XNAND2X1_LOC_763 NAND2X1_LOC_763/a_36_24# NAND2X1_LOC_763/Y VSS VDD INVX1_LOC_51/Y
+ INVX1_LOC_595/Y NAND2X1_LOC
XINVX1_LOC_607 INVX1_LOC_607/Y VSS VDD INVX1_LOC_607/A INVX1_LOC
XINVX1_LOC_618 INVX1_LOC_618/Y VSS VDD INVX1_LOC_618/A INVX1_LOC
XINVX1_LOC_7 INVX1_LOC_7/Y VSS VDD INVX1_LOC_7/A INVX1_LOC
XINVX1_LOC_629 INVX1_LOC_629/Y VSS VDD INVX1_LOC_629/A INVX1_LOC
XNAND2X1_LOC_593 NAND2X1_LOC_593/a_36_24# INVX1_LOC_460/A VSS VDD NAND2X1_LOC_591/Y
+ INVX1_LOC_459/Y NAND2X1_LOC
XNAND2X1_LOC_571 NAND2X1_LOC_571/a_36_24# INVX1_LOC_445/A VSS VDD INVX1_LOC_434/Y
+ INVX1_LOC_435/Y NAND2X1_LOC
XNAND2X1_LOC_582 NAND2X1_LOC_582/a_36_24# NAND2X1_LOC_635/B VSS VDD INVX1_LOC_479/A
+ INVX1_LOC_454/Y NAND2X1_LOC
XNAND2X1_LOC_560 NAND2X1_LOC_560/a_36_24# INVX1_LOC_434/A VSS VDD INVX1_LOC_406/Y
+ INVX1_LOC_433/Y NAND2X1_LOC
XINVX1_LOC_437 INVX1_LOC_437/Y VSS VDD INVX1_LOC_437/A INVX1_LOC
XINVX1_LOC_459 INVX1_LOC_459/Y VSS VDD INVX1_LOC_459/A INVX1_LOC
XINVX1_LOC_448 INVX1_LOC_448/Y VSS VDD INVX1_LOC_448/A INVX1_LOC
XINVX1_LOC_415 INVX1_LOC_415/Y VSS VDD INVX1_LOC_218/Y INVX1_LOC
XINVX1_LOC_426 INVX1_LOC_426/Y VSS VDD INVX1_LOC_426/A INVX1_LOC
XINVX1_LOC_404 INVX1_LOC_404/Y VSS VDD INVX1_LOC_224/Y INVX1_LOC
XNAND2X1_LOC_390 NAND2X1_LOC_390/a_36_24# INVX1_LOC_319/A VSS VDD INVX1_LOC_317/Y
+ INVX1_LOC_318/Y NAND2X1_LOC
XINVX1_LOC_245 INVX1_LOC_245/Y VSS VDD INVX1_LOC_245/A INVX1_LOC
XINVX1_LOC_212 INVX1_LOC_212/Y VSS VDD INVX1_LOC_212/A INVX1_LOC
XINVX1_LOC_278 INVX1_LOC_278/Y VSS VDD INVX1_LOC_278/A INVX1_LOC
XINVX1_LOC_256 INVX1_LOC_256/Y VSS VDD INVX1_LOC_256/A INVX1_LOC
XINVX1_LOC_289 INVX1_LOC_289/Y VSS VDD INVX1_LOC_289/A INVX1_LOC
XINVX1_LOC_234 INVX1_LOC_234/Y VSS VDD INPUT_0 INVX1_LOC
XINVX1_LOC_267 INVX1_LOC_267/Y VSS VDD INVX1_LOC_267/A INVX1_LOC
XINVX1_LOC_201 INVX1_LOC_201/Y VSS VDD INVX1_LOC_201/A INVX1_LOC
XINVX1_LOC_223 INVX1_LOC_223/Y VSS VDD INVX1_LOC_223/A INVX1_LOC
XNAND2X1_LOC_45 NAND2X1_LOC_45/a_36_24# NAND2X1_LOC_45/Y VSS VDD INVX1_LOC_32/Y INVX1_LOC_50/Y
+ NAND2X1_LOC
XNAND2X1_LOC_89 NAND2X1_LOC_89/a_36_24# NAND2X1_LOC_97/A VSS VDD INVX1_LOC_63/Y INVX1_LOC_80/A
+ NAND2X1_LOC
XNAND2X1_LOC_56 NAND2X1_LOC_56/a_36_24# NAND2X1_LOC_56/Y VSS VDD INVX1_LOC_59/Y INVX1_LOC_62/Y
+ NAND2X1_LOC
XNAND2X1_LOC_67 NAND2X1_LOC_67/a_36_24# NAND2X1_LOC_67/Y VSS VDD INVX1_LOC_62/Y NAND2X1_LOC_66/Y
+ NAND2X1_LOC
XNAND2X1_LOC_23 NAND2X1_LOC_23/a_36_24# INVX1_LOC_32/A VSS VDD INVX1_LOC_7/Y INVX1_LOC_21/Y
+ NAND2X1_LOC
XNAND2X1_LOC_12 NAND2X1_LOC_12/a_36_24# INVX1_LOC_20/A VSS VDD INVX1_LOC_1/Y INVX1_LOC_18/Y
+ NAND2X1_LOC
XNAND2X1_LOC_78 NAND2X1_LOC_78/a_36_24# NAND2X1_LOC_79/B VSS VDD INVX1_LOC_79/Y INVX1_LOC_80/Y
+ NAND2X1_LOC
XNAND2X1_LOC_34 NAND2X1_LOC_34/a_36_24# INVX1_LOC_43/A VSS VDD NAND2X1_LOC_27/Y NAND2X1_LOC_32/Y
+ NAND2X1_LOC
XNAND2X1_LOC_219 NAND2X1_LOC_219/a_36_24# INVX1_LOC_195/A VSS VDD INVX1_LOC_190/Y
+ INVX1_LOC_191/Y NAND2X1_LOC
XNAND2X1_LOC_208 NAND2X1_LOC_208/a_36_24# INVX1_LOC_184/A VSS VDD INVX1_LOC_44/Y INVX1_LOC_174/Y
+ NAND2X1_LOC
XNAND2X1_LOC_720 NAND2X1_LOC_720/a_36_24# INVX1_LOC_563/A VSS VDD NAND2X1_LOC_720/A
+ NAND2X1_LOC_669/Y NAND2X1_LOC
XNAND2X1_LOC_797 NAND2X1_LOC_797/a_36_24# INVX1_LOC_627/A VSS VDD INVX1_LOC_133/Y
+ INVX1_LOC_612/Y NAND2X1_LOC
XNAND2X1_LOC_731 NAND2X1_LOC_731/a_36_24# INVX1_LOC_574/A VSS VDD INVX1_LOC_569/Y
+ INVX1_LOC_570/Y NAND2X1_LOC
XNAND2X1_LOC_742 NAND2X1_LOC_742/a_36_24# GATE_741 VSS VDD INVX1_LOC_583/Y INVX1_LOC_584/Y
+ NAND2X1_LOC
XNAND2X1_LOC_775 NAND2X1_LOC_775/a_36_24# INVX1_LOC_603/A VSS VDD NAND2X1_LOC_97/B
+ NAND2X1_LOC_775/B NAND2X1_LOC
XNAND2X1_LOC_753 NAND2X1_LOC_753/a_36_24# NAND2X1_LOC_753/Y VSS VDD INVX1_LOC_588/Y
+ INVX1_LOC_587/Y NAND2X1_LOC
XNAND2X1_LOC_764 NAND2X1_LOC_764/a_36_24# NAND2X1_LOC_764/Y VSS VDD INVX1_LOC_48/Y
+ INVX1_LOC_117/Y NAND2X1_LOC
XNAND2X1_LOC_786 NAND2X1_LOC_786/a_36_24# INVX1_LOC_616/A VSS VDD INVX1_LOC_85/Y NAND2X1_LOC_786/B
+ NAND2X1_LOC
XINVX1_LOC_608 INVX1_LOC_608/Y VSS VDD INVX1_LOC_608/A INVX1_LOC
XINVX1_LOC_8 INVX1_LOC_8/Y VSS VDD INPUT_1 INVX1_LOC
XINVX1_LOC_619 INVX1_LOC_619/Y VSS VDD INVX1_LOC_619/A INVX1_LOC
XNAND2X1_LOC_550 NAND2X1_LOC_550/a_36_24# INVX1_LOC_424/A VSS VDD INVX1_LOC_420/Y
+ INVX1_LOC_421/Y NAND2X1_LOC
XNAND2X1_LOC_572 NAND2X1_LOC_572/a_36_24# INVX1_LOC_446/A VSS VDD INVX1_LOC_116/Y
+ INVX1_LOC_230/Y NAND2X1_LOC
XNAND2X1_LOC_561 NAND2X1_LOC_561/a_36_24# INVX1_LOC_435/A VSS VDD INVX1_LOC_431/Y
+ INVX1_LOC_432/Y NAND2X1_LOC
XNAND2X1_LOC_583 NAND2X1_LOC_583/a_36_24# NAND2X1_LOC_636/A VSS VDD INVX1_LOC_41/Y
+ INVX1_LOC_54/Y NAND2X1_LOC
XNAND2X1_LOC_594 NAND2X1_LOC_594/a_36_24# NAND2X1_LOC_594/Y VSS VDD INVX1_LOC_93/Y
+ NAND2X1_LOC_331/A NAND2X1_LOC
XINVX1_LOC_427 INVX1_LOC_427/Y VSS VDD INVX1_LOC_427/A INVX1_LOC
XINVX1_LOC_449 INVX1_LOC_449/Y VSS VDD INVX1_LOC_449/A INVX1_LOC
XINVX1_LOC_416 INVX1_LOC_416/Y VSS VDD INVX1_LOC_416/A INVX1_LOC
XINVX1_LOC_405 INVX1_LOC_405/Y VSS VDD INVX1_LOC_405/A INVX1_LOC
XINVX1_LOC_438 INVX1_LOC_438/Y VSS VDD INVX1_LOC_438/A INVX1_LOC
XNAND2X1_LOC_391 NAND2X1_LOC_391/a_36_24# INVX1_LOC_320/A VSS VDD NAND2X1_LOC_391/A
+ NAND2X1_LOC_391/B NAND2X1_LOC
XNAND2X1_LOC_380 NAND2X1_LOC_380/a_36_24# NAND2X1_LOC_460/A VSS VDD INVX1_LOC_117/Y
+ NAND2X1_LOC_379/Y NAND2X1_LOC
XINVX1_LOC_213 INVX1_LOC_213/Y VSS VDD INVX1_LOC_11/Y INVX1_LOC
XINVX1_LOC_279 INVX1_LOC_279/Y VSS VDD INVX1_LOC_279/A INVX1_LOC
XINVX1_LOC_257 INVX1_LOC_257/Y VSS VDD INVX1_LOC_257/A INVX1_LOC
XINVX1_LOC_235 INVX1_LOC_235/Y VSS VDD INVX1_LOC_235/A INVX1_LOC
XINVX1_LOC_246 INVX1_LOC_246/Y VSS VDD INVX1_LOC_49/Y INVX1_LOC
XINVX1_LOC_268 INVX1_LOC_268/Y VSS VDD INVX1_LOC_268/A INVX1_LOC
XINVX1_LOC_224 INVX1_LOC_224/Y VSS VDD INVX1_LOC_224/A INVX1_LOC
XINVX1_LOC_202 INVX1_LOC_202/Y VSS VDD INVX1_LOC_202/A INVX1_LOC
XNAND2X1_LOC_46 NAND2X1_LOC_46/a_36_24# INVX1_LOC_51/A VSS VDD INVX1_LOC_52/Y INVX1_LOC_21/Y
+ NAND2X1_LOC
XNAND2X1_LOC_13 NAND2X1_LOC_13/a_36_24# NAND2X1_LOC_13/Y VSS VDD INVX1_LOC_17/Y INVX1_LOC_20/Y
+ NAND2X1_LOC
XNAND2X1_LOC_57 NAND2X1_LOC_57/a_36_24# NAND2X1_LOC_57/Y VSS VDD INVX1_LOC_9/Y INVX1_LOC_50/Y
+ NAND2X1_LOC
XNAND2X1_LOC_68 NAND2X1_LOC_68/a_36_24# NAND2X1_LOC_69/B VSS VDD INVX1_LOC_72/Y INVX1_LOC_73/Y
+ NAND2X1_LOC
XNAND2X1_LOC_24 NAND2X1_LOC_24/a_36_24# NAND2X1_LOC_24/Y VSS VDD INVX1_LOC_31/Y INVX1_LOC_32/Y
+ NAND2X1_LOC
XNAND2X1_LOC_79 NAND2X1_LOC_79/a_36_24# NAND2X1_LOC_79/Y VSS VDD INVX1_LOC_26/Y NAND2X1_LOC_79/B
+ NAND2X1_LOC
XNAND2X1_LOC_35 NAND2X1_LOC_35/a_36_24# INVX1_LOC_44/A VSS VDD INVX1_LOC_42/Y INVX1_LOC_43/Y
+ NAND2X1_LOC
XNAND2X1_LOC_209 NAND2X1_LOC_209/a_36_24# INVX1_LOC_185/A VSS VDD INVX1_LOC_133/Y
+ NAND2X1_LOC_152/Y NAND2X1_LOC
XNAND2X1_LOC_710 NAND2X1_LOC_710/a_36_24# INVX1_LOC_553/A VSS VDD NAND2X1_LOC_710/A
+ NAND2X1_LOC_710/B NAND2X1_LOC
XNAND2X1_LOC_743 NAND2X1_LOC_743/a_36_24# NAND2X1_LOC_780/A VSS VDD INVX1_LOC_6/Y
+ INVX1_LOC_137/Y NAND2X1_LOC
XNAND2X1_LOC_732 NAND2X1_LOC_732/a_36_24# INVX1_LOC_575/A VSS VDD INVX1_LOC_567/Y
+ INVX1_LOC_568/Y NAND2X1_LOC
XNAND2X1_LOC_754 NAND2X1_LOC_754/a_36_24# NAND2X1_LOC_790/B VSS VDD INVX1_LOC_45/Y
+ NAND2X1_LOC_615/B NAND2X1_LOC
XNAND2X1_LOC_721 NAND2X1_LOC_721/a_36_24# INVX1_LOC_564/A VSS VDD INVX1_LOC_531/Y
+ INVX1_LOC_563/Y NAND2X1_LOC
XNAND2X1_LOC_798 NAND2X1_LOC_798/a_36_24# INVX1_LOC_628/A VSS VDD INVX1_LOC_255/Y
+ INVX1_LOC_346/Y NAND2X1_LOC
XNAND2X1_LOC_787 NAND2X1_LOC_787/a_36_24# INVX1_LOC_617/A VSS VDD INVX1_LOC_301/Y
+ INVX1_LOC_387/Y NAND2X1_LOC
XNAND2X1_LOC_765 NAND2X1_LOC_765/a_36_24# NAND2X1_LOC_770/A VSS VDD INVX1_LOC_20/Y
+ INVX1_LOC_79/A NAND2X1_LOC
XNAND2X1_LOC_776 NAND2X1_LOC_776/a_36_24# INVX1_LOC_604/A VSS VDD NAND2X1_LOC_164/Y
+ NAND2X1_LOC_241/B NAND2X1_LOC
XINVX1_LOC_9 INVX1_LOC_9/Y VSS VDD INVX1_LOC_9/A INVX1_LOC
XINVX1_LOC_609 INVX1_LOC_609/Y VSS VDD INVX1_LOC_609/A INVX1_LOC
XNAND2X1_LOC_540 NAND2X1_LOC_540/a_36_24# INVX1_LOC_413/A VSS VDD NAND2X1_LOC_181/A
+ NAND2X1_LOC_190/A NAND2X1_LOC
XNAND2X1_LOC_595 NAND2X1_LOC_595/a_36_24# NAND2X1_LOC_595/Y VSS VDD INVX1_LOC_35/Y
+ NAND2X1_LOC_249/Y NAND2X1_LOC
XNAND2X1_LOC_562 NAND2X1_LOC_562/a_36_24# INVX1_LOC_436/A VSS VDD INVX1_LOC_429/Y
+ INVX1_LOC_430/Y NAND2X1_LOC
XNAND2X1_LOC_584 NAND2X1_LOC_584/a_36_24# NAND2X1_LOC_636/B VSS VDD INVX1_LOC_11/Y
+ INVX1_LOC_58/Y NAND2X1_LOC
XNAND2X1_LOC_551 NAND2X1_LOC_551/a_36_24# INVX1_LOC_425/A VSS VDD INVX1_LOC_418/Y
+ INVX1_LOC_419/Y NAND2X1_LOC
XNAND2X1_LOC_573 NAND2X1_LOC_573/a_36_24# INVX1_LOC_447/A VSS VDD INVX1_LOC_328/Y
+ INVX1_LOC_393/Y NAND2X1_LOC
XINVX1_LOC_428 INVX1_LOC_428/Y VSS VDD INVX1_LOC_428/A INVX1_LOC
XINVX1_LOC_406 INVX1_LOC_406/Y VSS VDD INVX1_LOC_406/A INVX1_LOC
XINVX1_LOC_417 INVX1_LOC_417/Y VSS VDD INVX1_LOC_417/A INVX1_LOC
XINVX1_LOC_439 INVX1_LOC_439/Y VSS VDD INVX1_LOC_439/A INVX1_LOC
XNAND2X1_LOC_370 NAND2X1_LOC_370/a_36_24# INVX1_LOC_301/A VSS VDD NAND2X1_LOC_370/A
+ NAND2X1_LOC_543/B NAND2X1_LOC
XNAND2X1_LOC_392 NAND2X1_LOC_392/a_36_24# INVX1_LOC_321/A VSS VDD INVX1_LOC_319/Y
+ INVX1_LOC_320/Y NAND2X1_LOC
XNAND2X1_LOC_381 NAND2X1_LOC_381/a_36_24# INVX1_LOC_312/A VSS VDD INPUT_3 INVX1_LOC_20/Y
+ NAND2X1_LOC
XINVX1_LOC_214 INVX1_LOC_214/Y VSS VDD INVX1_LOC_17/Y INVX1_LOC
XINVX1_LOC_225 INVX1_LOC_225/Y VSS VDD INVX1_LOC_17/Y INVX1_LOC
XINVX1_LOC_203 INVX1_LOC_203/Y VSS VDD INVX1_LOC_203/A INVX1_LOC
XNAND2X1_LOC_25 NAND2X1_LOC_25/a_36_24# INVX1_LOC_33/A VSS VDD INPUT_6 INVX1_LOC_34/Y
+ NAND2X1_LOC
XNAND2X1_LOC_14 NAND2X1_LOC_14/a_36_24# INVX1_LOC_21/A VSS VDD INVX1_LOC_22/Y INVX1_LOC_23/Y
+ NAND2X1_LOC
XINVX1_LOC_236 INVX1_LOC_492/A VSS VDD INVX1_LOC_236/A INVX1_LOC
XINVX1_LOC_258 INVX1_LOC_258/Y VSS VDD INVX1_LOC_258/A INVX1_LOC
XINVX1_LOC_247 INVX1_LOC_247/Y VSS VDD INVX1_LOC_62/Y INVX1_LOC
XINVX1_LOC_269 INVX1_LOC_269/Y VSS VDD INVX1_LOC_269/A INVX1_LOC
XNAND2X1_LOC_36 NAND2X1_LOC_36/a_36_24# INVX1_LOC_45/A VSS VDD INVX1_LOC_25/Y INVX1_LOC_29/Y
+ NAND2X1_LOC
XNAND2X1_LOC_47 NAND2X1_LOC_47/a_36_24# INVX1_LOC_53/A VSS VDD INVX1_LOC_33/Y INVX1_LOC_40/Y
+ NAND2X1_LOC
XNAND2X1_LOC_58 NAND2X1_LOC_58/a_36_24# NAND2X1_LOC_61/A VSS VDD INVX1_LOC_31/Y INVX1_LOC_54/Y
+ NAND2X1_LOC
XNAND2X1_LOC_69 NAND2X1_LOC_69/a_36_24# NAND2X1_LOC_69/Y VSS VDD INVX1_LOC_45/Y NAND2X1_LOC_69/B
+ NAND2X1_LOC
XNAND2X1_LOC_700 NAND2X1_LOC_700/a_36_24# NAND2X1_LOC_710/A VSS VDD INVX1_LOC_63/Y
+ INVX1_LOC_89/Y NAND2X1_LOC
XNAND2X1_LOC_788 NAND2X1_LOC_788/a_36_24# INVX1_LOC_618/A VSS VDD NAND2X1_LOC_788/A
+ INVX1_LOC_468/Y NAND2X1_LOC
XNAND2X1_LOC_711 NAND2X1_LOC_711/a_36_24# INVX1_LOC_554/A VSS VDD INVX1_LOC_551/Y
+ INVX1_LOC_553/Y NAND2X1_LOC
XNAND2X1_LOC_744 NAND2X1_LOC_744/a_36_24# NAND2X1_LOC_780/B VSS VDD INVX1_LOC_50/Y
+ INVX1_LOC_117/Y NAND2X1_LOC
XNAND2X1_LOC_777 NAND2X1_LOC_777/a_36_24# INVX1_LOC_605/A VSS VDD INVX1_LOC_606/Y
+ NAND2X1_LOC_307/B NAND2X1_LOC
XNAND2X1_LOC_722 NAND2X1_LOC_722/a_36_24# INVX1_LOC_565/A VSS VDD INVX1_LOC_561/Y
+ INVX1_LOC_562/Y NAND2X1_LOC
XNAND2X1_LOC_733 NAND2X1_LOC_733/a_36_24# INVX1_LOC_576/A VSS VDD INVX1_LOC_565/Y
+ INVX1_LOC_566/Y NAND2X1_LOC
XNAND2X1_LOC_755 NAND2X1_LOC_755/a_36_24# NAND2X1_LOC_791/A VSS VDD INVX1_LOC_63/Y
+ NAND2X1_LOC_755/B NAND2X1_LOC
XNAND2X1_LOC_766 NAND2X1_LOC_766/a_36_24# NAND2X1_LOC_770/B VSS VDD INVX1_LOC_69/Y
+ INVX1_LOC_89/Y NAND2X1_LOC
XNAND2X1_LOC_799 NAND2X1_LOC_799/a_36_24# INVX1_LOC_629/A VSS VDD INVX1_LOC_412/Y
+ INVX1_LOC_460/Y NAND2X1_LOC
XNAND2X1_LOC_541 NAND2X1_LOC_541/a_36_24# INVX1_LOC_414/A VSS VDD INVX1_LOC_415/Y
+ NAND2X1_LOC_541/B NAND2X1_LOC
XNAND2X1_LOC_574 NAND2X1_LOC_574/a_36_24# INVX1_LOC_448/A VSS VDD INVX1_LOC_400/Y
+ NAND2X1_LOC_516/Y NAND2X1_LOC
XNAND2X1_LOC_596 NAND2X1_LOC_596/a_36_24# NAND2X1_LOC_596/Y VSS VDD INVX1_LOC_461/Y
+ INVX1_LOC_462/Y NAND2X1_LOC
XNAND2X1_LOC_563 NAND2X1_LOC_563/a_36_24# INVX1_LOC_437/A VSS VDD INVX1_LOC_427/Y
+ INVX1_LOC_428/Y NAND2X1_LOC
XNAND2X1_LOC_585 NAND2X1_LOC_585/a_36_24# NAND2X1_LOC_637/A VSS VDD INVX1_LOC_31/Y
+ INVX1_LOC_245/A NAND2X1_LOC
XNAND2X1_LOC_552 NAND2X1_LOC_552/a_36_24# INVX1_LOC_426/A VSS VDD INVX1_LOC_416/Y
+ INVX1_LOC_417/Y NAND2X1_LOC
XNAND2X1_LOC_530 NAND2X1_LOC_530/a_36_24# NAND2X1_LOC_548/B VSS VDD INVX1_LOC_45/Y
+ INVX1_LOC_99/Y NAND2X1_LOC
XINVX1_LOC_407 INVX1_LOC_407/Y VSS VDD INVX1_LOC_99/Y INVX1_LOC
XINVX1_LOC_429 INVX1_LOC_429/Y VSS VDD INVX1_LOC_429/A INVX1_LOC
XINVX1_LOC_418 INVX1_LOC_418/Y VSS VDD INVX1_LOC_418/A INVX1_LOC
XNAND2X1_LOC_371 NAND2X1_LOC_371/a_36_24# INVX1_LOC_302/A VSS VDD INVX1_LOC_9/Y INVX1_LOC_41/Y
+ NAND2X1_LOC
XNAND2X1_LOC_382 NAND2X1_LOC_382/a_36_24# NAND2X1_LOC_391/A VSS VDD INVX1_LOC_84/A
+ INVX1_LOC_312/Y NAND2X1_LOC
XNAND2X1_LOC_360 NAND2X1_LOC_360/a_36_24# INVX1_LOC_294/A VSS VDD INVX1_LOC_211/Y
+ INVX1_LOC_281/Y NAND2X1_LOC
XNAND2X1_LOC_393 NAND2X1_LOC_393/a_36_24# NAND2X1_LOC_393/Y VSS VDD INVX1_LOC_47/Y
+ INVX1_LOC_48/Y NAND2X1_LOC
XINVX1_LOC_237 INVX1_LOC_237/Y VSS VDD INVX1_LOC_66/A INVX1_LOC
XINVX1_LOC_215 INVX1_LOC_215/Y VSS VDD INVX1_LOC_32/Y INVX1_LOC
XINVX1_LOC_259 INVX1_LOC_259/Y VSS VDD INVX1_LOC_259/A INVX1_LOC
XINVX1_LOC_248 INVX1_LOC_248/Y VSS VDD INVX1_LOC_248/A INVX1_LOC
XINVX1_LOC_226 INVX1_LOC_226/Y VSS VDD INVX1_LOC_80/A INVX1_LOC
XINVX1_LOC_204 INVX1_LOC_204/Y VSS VDD INVX1_LOC_204/A INVX1_LOC
XNAND2X1_LOC_15 NAND2X1_LOC_15/a_36_24# INVX1_LOC_24/A VSS VDD INVX1_LOC_66/A INVX1_LOC_21/Y
+ NAND2X1_LOC
XNAND2X1_LOC_26 NAND2X1_LOC_26/a_36_24# INVX1_LOC_35/A VSS VDD INVX1_LOC_29/Y INVX1_LOC_33/Y
+ NAND2X1_LOC
XNAND2X1_LOC_59 NAND2X1_LOC_59/a_36_24# INVX1_LOC_63/A VSS VDD INVX1_LOC_18/Y INVX1_LOC_33/Y
+ NAND2X1_LOC
XNAND2X1_LOC_48 NAND2X1_LOC_48/a_36_24# NAND2X1_LOC_48/Y VSS VDD INVX1_LOC_51/Y INVX1_LOC_53/Y
+ NAND2X1_LOC
XNAND2X1_LOC_37 NAND2X1_LOC_37/a_36_24# INVX1_LOC_46/A VSS VDD INPUT_2 INPUT_3
+ NAND2X1_LOC
XNAND2X1_LOC_190 NAND2X1_LOC_190/a_36_24# INVX1_LOC_166/A VSS VDD NAND2X1_LOC_190/A
+ NAND2X1_LOC_184/Y NAND2X1_LOC
XINVX1_LOC_590 INVX1_LOC_590/Y VSS VDD INVX1_LOC_586/A INVX1_LOC
XNAND2X1_LOC_701 NAND2X1_LOC_701/a_36_24# NAND2X1_LOC_710/B VSS VDD INVX1_LOC_50/Y
+ INVX1_LOC_206/Y NAND2X1_LOC
XNAND2X1_LOC_778 NAND2X1_LOC_778/a_36_24# INVX1_LOC_607/A VSS VDD INVX1_LOC_608/Y
+ NAND2X1_LOC_496/Y NAND2X1_LOC
XNAND2X1_LOC_745 NAND2X1_LOC_745/a_36_24# NAND2X1_LOC_781/A VSS VDD INVX1_LOC_48/Y
+ INVX1_LOC_586/A NAND2X1_LOC
XNAND2X1_LOC_712 NAND2X1_LOC_712/a_36_24# INVX1_LOC_555/A VSS VDD INVX1_LOC_549/Y
+ INVX1_LOC_550/Y NAND2X1_LOC
XNAND2X1_LOC_723 NAND2X1_LOC_723/a_36_24# INVX1_LOC_566/A VSS VDD INVX1_LOC_559/Y
+ INVX1_LOC_560/Y NAND2X1_LOC
XNAND2X1_LOC_734 NAND2X1_LOC_734/a_36_24# INVX1_LOC_577/A VSS VDD NAND2X1_LOC_475/A
+ INVX1_LOC_564/Y NAND2X1_LOC
XNAND2X1_LOC_756 NAND2X1_LOC_756/a_36_24# NAND2X1_LOC_756/Y VSS VDD INVX1_LOC_589/Y
+ INVX1_LOC_590/Y NAND2X1_LOC
XNAND2X1_LOC_767 NAND2X1_LOC_767/a_36_24# NAND2X1_LOC_773/A VSS VDD INVX1_LOC_6/Y
+ NAND2X1_LOC_79/B NAND2X1_LOC
XNAND2X1_LOC_789 NAND2X1_LOC_789/a_36_24# INVX1_LOC_619/A VSS VDD NAND2X1_LOC_789/A
+ NAND2X1_LOC_789/B NAND2X1_LOC
XNAND2X1_LOC_520 NAND2X1_LOC_520/a_36_24# INVX1_LOC_405/A VSS VDD NAND2X1_LOC_520/A
+ NAND2X1_LOC_520/B NAND2X1_LOC
XNAND2X1_LOC_586 NAND2X1_LOC_586/a_36_24# NAND2X1_LOC_586/Y VSS VDD INVX1_LOC_74/Y
+ INVX1_LOC_119/Y NAND2X1_LOC
XNAND2X1_LOC_575 NAND2X1_LOC_575/a_36_24# INVX1_LOC_449/A VSS VDD INVX1_LOC_447/Y
+ INVX1_LOC_448/Y NAND2X1_LOC
XNAND2X1_LOC_597 NAND2X1_LOC_597/a_36_24# NAND2X1_LOC_597/Y VSS VDD INVX1_LOC_17/Y
+ NAND2X1_LOC_596/Y NAND2X1_LOC
XNAND2X1_LOC_553 NAND2X1_LOC_553/a_36_24# INVX1_LOC_427/A VSS VDD INVX1_LOC_413/Y
+ INVX1_LOC_414/Y NAND2X1_LOC
XNAND2X1_LOC_542 NAND2X1_LOC_542/a_36_24# INVX1_LOC_416/A VSS VDD NAND2X1_LOC_542/A
+ NAND2X1_LOC_336/B NAND2X1_LOC
XNAND2X1_LOC_564 NAND2X1_LOC_564/a_36_24# INVX1_LOC_438/A VSS VDD INVX1_LOC_425/Y
+ INVX1_LOC_426/Y NAND2X1_LOC
XNAND2X1_LOC_531 NAND2X1_LOC_531/a_36_24# NAND2X1_LOC_531/Y VSS VDD INVX1_LOC_48/Y
+ INVX1_LOC_76/Y NAND2X1_LOC
XINVX1_LOC_408 INVX1_LOC_408/Y VSS VDD INVX1_LOC_117/Y INVX1_LOC
XINVX1_LOC_419 INVX1_LOC_419/Y VSS VDD INVX1_LOC_419/A INVX1_LOC
XNAND2X1_LOC_372 NAND2X1_LOC_372/a_36_24# NAND2X1_LOC_372/Y VSS VDD INVX1_LOC_303/Y
+ INVX1_LOC_608/A NAND2X1_LOC
XNAND2X1_LOC_361 NAND2X1_LOC_361/a_36_24# INVX1_LOC_295/A VSS VDD INVX1_LOC_230/Y
+ INVX1_LOC_235/Y NAND2X1_LOC
XNAND2X1_LOC_350 NAND2X1_LOC_350/a_36_24# INVX1_LOC_284/A VSS VDD INVX1_LOC_274/Y
+ INVX1_LOC_275/Y NAND2X1_LOC
XNAND2X1_LOC_383 NAND2X1_LOC_383/a_36_24# NAND2X1_LOC_383/Y VSS VDD INVX1_LOC_313/Y
+ INVX1_LOC_314/Y NAND2X1_LOC
XNAND2X1_LOC_394 NAND2X1_LOC_394/a_36_24# NAND2X1_LOC_400/B VSS VDD INVX1_LOC_53/Y
+ INVX1_LOC_117/Y NAND2X1_LOC
XINVX1_LOC_238 INVX1_LOC_238/Y VSS VDD INVX1_LOC_238/A INVX1_LOC
XINVX1_LOC_216 INVX1_LOC_216/Y VSS VDD INVX1_LOC_47/Y INVX1_LOC
XINVX1_LOC_249 INVX1_LOC_249/Y VSS VDD INVX1_LOC_249/A INVX1_LOC
XINVX1_LOC_227 INVX1_LOC_227/Y VSS VDD INVX1_LOC_224/Y INVX1_LOC
XINVX1_LOC_205 INVX1_LOC_205/Y VSS VDD INVX1_LOC_65/Y INVX1_LOC
XNAND2X1_LOC_191 NAND2X1_LOC_191/a_36_24# INVX1_LOC_167/A VSS VDD NAND2X1_LOC_187/Y
+ INVX1_LOC_166/Y NAND2X1_LOC
XNAND2X1_LOC_180 NAND2X1_LOC_180/a_36_24# INVX1_LOC_158/A VSS VDD NAND2X1_LOC_176/Y
+ NAND2X1_LOC_180/B NAND2X1_LOC
XNAND2X1_LOC_16 NAND2X1_LOC_16/a_36_24# NAND2X1_LOC_16/Y VSS VDD INVX1_LOC_6/Y INVX1_LOC_79/A
+ NAND2X1_LOC
XNAND2X1_LOC_38 NAND2X1_LOC_38/a_36_24# INVX1_LOC_47/A VSS VDD INVX1_LOC_84/A INVX1_LOC_46/Y
+ NAND2X1_LOC
XNAND2X1_LOC_27 NAND2X1_LOC_27/a_36_24# NAND2X1_LOC_27/Y VSS VDD INVX1_LOC_11/Y INVX1_LOC_35/Y
+ NAND2X1_LOC
XNAND2X1_LOC_49 NAND2X1_LOC_49/a_36_24# INVX1_LOC_54/A VSS VDD INVX1_LOC_21/Y INVX1_LOC_84/A
+ NAND2X1_LOC
XINVX1_LOC_580 INVX1_LOC_580/Y VSS VDD INVX1_LOC_580/A INVX1_LOC
XINVX1_LOC_591 INVX1_LOC_591/Y VSS VDD INVX1_LOC_48/Y INVX1_LOC
XNAND2X1_LOC_702 NAND2X1_LOC_702/a_36_24# INVX1_LOC_544/A VSS VDD NAND2X1_LOC_45/Y
+ NAND2X1_LOC_332/B NAND2X1_LOC
XNAND2X1_LOC_724 NAND2X1_LOC_724/a_36_24# INVX1_LOC_567/A VSS VDD INVX1_LOC_557/Y
+ INVX1_LOC_558/Y NAND2X1_LOC
XNAND2X1_LOC_713 NAND2X1_LOC_713/a_36_24# INVX1_LOC_556/A VSS VDD INVX1_LOC_547/Y
+ INVX1_LOC_548/Y NAND2X1_LOC
XNAND2X1_LOC_768 NAND2X1_LOC_768/a_36_24# INVX1_LOC_596/A VSS VDD NAND2X1_LOC_768/A
+ NAND2X1_LOC_768/B NAND2X1_LOC
XNAND2X1_LOC_779 NAND2X1_LOC_779/a_36_24# INVX1_LOC_609/A VSS VDD NAND2X1_LOC_513/A
+ NAND2X1_LOC_697/Y NAND2X1_LOC
XNAND2X1_LOC_746 NAND2X1_LOC_746/a_36_24# NAND2X1_LOC_781/B VSS VDD INVX1_LOC_76/Y
+ INVX1_LOC_145/Y NAND2X1_LOC
XNAND2X1_LOC_735 NAND2X1_LOC_735/a_36_24# INVX1_LOC_578/A VSS VDD INVX1_LOC_393/Y
+ INVX1_LOC_490/Y NAND2X1_LOC
XNAND2X1_LOC_757 NAND2X1_LOC_757/a_36_24# NAND2X1_LOC_791/B VSS VDD INVX1_LOC_50/Y
+ NAND2X1_LOC_756/Y NAND2X1_LOC
XNAND2X1_LOC_521 NAND2X1_LOC_521/a_36_24# NAND2X1_LOC_521/Y VSS VDD INVX1_LOC_26/Y
+ INVX1_LOC_54/Y NAND2X1_LOC
XNAND2X1_LOC_554 NAND2X1_LOC_554/a_36_24# INVX1_LOC_428/A VSS VDD NAND2X1_LOC_106/Y
+ INVX1_LOC_118/Y NAND2X1_LOC
XNAND2X1_LOC_532 NAND2X1_LOC_532/a_36_24# NAND2X1_LOC_532/Y VSS VDD INVX1_LOC_407/Y
+ INVX1_LOC_408/Y NAND2X1_LOC
XNAND2X1_LOC_543 NAND2X1_LOC_543/a_36_24# INVX1_LOC_417/A VSS VDD NAND2X1_LOC_318/A
+ NAND2X1_LOC_543/B NAND2X1_LOC
XNAND2X1_LOC_510 NAND2X1_LOC_510/a_36_24# INVX1_LOC_400/A VSS VDD INVX1_LOC_398/Y
+ INVX1_LOC_399/Y NAND2X1_LOC
XNAND2X1_LOC_598 NAND2X1_LOC_598/a_36_24# INVX1_LOC_463/A VSS VDD INVX1_LOC_464/Y
+ INVX1_LOC_465/Y NAND2X1_LOC
XNAND2X1_LOC_576 NAND2X1_LOC_576/a_36_24# INVX1_LOC_450/A VSS VDD INVX1_LOC_445/Y
+ INVX1_LOC_446/Y NAND2X1_LOC
XNAND2X1_LOC_565 NAND2X1_LOC_565/a_36_24# INVX1_LOC_439/A VSS VDD INVX1_LOC_423/Y
+ INVX1_LOC_424/Y NAND2X1_LOC
XNAND2X1_LOC_587 NAND2X1_LOC_587/a_36_24# INVX1_LOC_455/A VSS VDD INVX1_LOC_456/Y
+ INVX1_LOC_40/Y NAND2X1_LOC
XINVX1_LOC_409 INVX1_LOC_409/Y VSS VDD INVX1_LOC_409/A INVX1_LOC
XNAND2X1_LOC_373 NAND2X1_LOC_373/a_36_24# NAND2X1_LOC_373/Y VSS VDD INVX1_LOC_35/Y
+ INVX1_LOC_80/A NAND2X1_LOC
XNAND2X1_LOC_362 NAND2X1_LOC_362/a_36_24# INVX1_LOC_296/A VSS VDD INVX1_LOC_242/Y
+ INVX1_LOC_295/Y NAND2X1_LOC
XNAND2X1_LOC_384 NAND2X1_LOC_384/a_36_24# NAND2X1_LOC_391/B VSS VDD INVX1_LOC_48/Y
+ NAND2X1_LOC_383/Y NAND2X1_LOC
XNAND2X1_LOC_351 NAND2X1_LOC_351/a_36_24# INVX1_LOC_285/A VSS VDD INVX1_LOC_272/Y
+ INVX1_LOC_273/Y NAND2X1_LOC
XNAND2X1_LOC_340 NAND2X1_LOC_340/a_36_24# INVX1_LOC_274/A VSS VDD NAND2X1_LOC_88/Y
+ INVX1_LOC_201/Y NAND2X1_LOC
XNAND2X1_LOC_395 NAND2X1_LOC_395/a_36_24# NAND2X1_LOC_395/Y VSS VDD INVX1_LOC_63/Y
+ INVX1_LOC_100/Y NAND2X1_LOC
XINVX1_LOC_239 INVX1_LOC_239/Y VSS VDD INVX1_LOC_239/A INVX1_LOC
XINVX1_LOC_217 INVX1_LOC_217/Y VSS VDD INVX1_LOC_217/A INVX1_LOC
XINVX1_LOC_228 INVX1_LOC_228/Y VSS VDD INVX1_LOC_228/A INVX1_LOC
XINVX1_LOC_206 INVX1_LOC_206/Y VSS VDD INVX1_LOC_206/A INVX1_LOC
XNAND2X1_LOC_192 NAND2X1_LOC_192/a_36_24# INVX1_LOC_168/A VSS VDD NAND2X1_LOC_192/A
+ INVX1_LOC_167/Y NAND2X1_LOC
XNAND2X1_LOC_181 NAND2X1_LOC_181/a_36_24# INVX1_LOC_159/A VSS VDD NAND2X1_LOC_181/A
+ NAND2X1_LOC_179/Y NAND2X1_LOC
XNAND2X1_LOC_170 NAND2X1_LOC_170/a_36_24# INVX1_LOC_155/A VSS VDD INVX1_LOC_153/Y
+ INVX1_LOC_154/Y NAND2X1_LOC
XNAND2X1_LOC_28 NAND2X1_LOC_28/a_36_24# INVX1_LOC_36/A VSS VDD INVX1_LOC_37/Y INPUT_1
+ NAND2X1_LOC
XNAND2X1_LOC_39 NAND2X1_LOC_39/a_36_24# NAND2X1_LOC_39/Y VSS VDD INVX1_LOC_45/Y INVX1_LOC_47/Y
+ NAND2X1_LOC
XNAND2X1_LOC_17 NAND2X1_LOC_17/a_36_24# INVX1_LOC_25/A VSS VDD INPUT_6 INPUT_7
+ NAND2X1_LOC
XINVX1_LOC_581 INVX1_LOC_581/Y VSS VDD INVX1_LOC_581/A INVX1_LOC
XINVX1_LOC_570 INVX1_LOC_570/Y VSS VDD INVX1_LOC_570/A INVX1_LOC
XINVX1_LOC_592 INVX1_LOC_592/Y VSS VDD INVX1_LOC_93/Y INVX1_LOC
XNAND2X1_LOC_714 NAND2X1_LOC_714/a_36_24# INVX1_LOC_557/A VSS VDD INVX1_LOC_545/Y
+ INVX1_LOC_546/Y NAND2X1_LOC
XNAND2X1_LOC_725 NAND2X1_LOC_725/a_36_24# INVX1_LOC_568/A VSS VDD INVX1_LOC_555/Y
+ INVX1_LOC_556/Y NAND2X1_LOC
XNAND2X1_LOC_736 NAND2X1_LOC_736/a_36_24# INVX1_LOC_579/A VSS VDD INVX1_LOC_533/Y
+ INVX1_LOC_578/Y NAND2X1_LOC
XNAND2X1_LOC_703 NAND2X1_LOC_703/a_36_24# INVX1_LOC_545/A VSS VDD NAND2X1_LOC_388/A
+ NAND2X1_LOC_336/B NAND2X1_LOC
XNAND2X1_LOC_747 NAND2X1_LOC_747/a_36_24# NAND2X1_LOC_782/A VSS VDD INVX1_LOC_53/Y
+ INVX1_LOC_54/Y NAND2X1_LOC
XNAND2X1_LOC_758 NAND2X1_LOC_758/a_36_24# NAND2X1_LOC_759/B VSS VDD INVX1_LOC_591/Y
+ INVX1_LOC_592/Y NAND2X1_LOC
XNAND2X1_LOC_769 NAND2X1_LOC_769/a_36_24# INVX1_LOC_597/A VSS VDD NAND2X1_LOC_763/Y
+ NAND2X1_LOC_764/Y NAND2X1_LOC
XNAND2X1_LOC_544 NAND2X1_LOC_544/a_36_24# INVX1_LOC_418/A VSS VDD NAND2X1_LOC_373/Y
+ NAND2X1_LOC_544/B NAND2X1_LOC
XNAND2X1_LOC_522 NAND2X1_LOC_522/a_36_24# NAND2X1_LOC_523/B VSS VDD INVX1_LOC_31/Y
+ INVX1_LOC_99/Y NAND2X1_LOC
XNAND2X1_LOC_500 NAND2X1_LOC_500/a_36_24# INVX1_LOC_392/A VSS VDD NAND2X1_LOC_844/A
+ INVX1_LOC_391/Y NAND2X1_LOC
XNAND2X1_LOC_533 NAND2X1_LOC_533/a_36_24# NAND2X1_LOC_788/A VSS VDD INVX1_LOC_93/Y
+ NAND2X1_LOC_532/Y NAND2X1_LOC
XNAND2X1_LOC_555 NAND2X1_LOC_555/a_36_24# INVX1_LOC_429/A VSS VDD INVX1_LOC_220/Y
+ NAND2X1_LOC_555/B NAND2X1_LOC
XNAND2X1_LOC_511 NAND2X1_LOC_511/a_36_24# NAND2X1_LOC_513/A VSS VDD INVX1_LOC_41/Y
+ INVX1_LOC_51/Y NAND2X1_LOC
XNAND2X1_LOC_566 NAND2X1_LOC_566/a_36_24# INVX1_LOC_440/A VSS VDD INVX1_LOC_155/Y
+ INVX1_LOC_250/Y NAND2X1_LOC
XNAND2X1_LOC_588 NAND2X1_LOC_588/a_36_24# NAND2X1_LOC_638/A VSS VDD INVX1_LOC_395/A
+ INVX1_LOC_455/Y NAND2X1_LOC
XNAND2X1_LOC_577 NAND2X1_LOC_577/a_36_24# INVX1_LOC_451/A VSS VDD INVX1_LOC_443/Y
+ INVX1_LOC_444/Y NAND2X1_LOC
XNAND2X1_LOC_599 NAND2X1_LOC_599/a_36_24# INVX1_LOC_466/A VSS VDD INVX1_LOC_45/Y INVX1_LOC_467/Y
+ NAND2X1_LOC
XNAND2X1_LOC_374 NAND2X1_LOC_374/a_36_24# INVX1_LOC_304/A VSS VDD NAND2X1_LOC_322/Y
+ NAND2X1_LOC_373/Y NAND2X1_LOC
XNAND2X1_LOC_330 NAND2X1_LOC_330/a_36_24# NAND2X1_LOC_331/B VSS VDD INVX1_LOC_264/Y
+ INVX1_LOC_265/Y NAND2X1_LOC
XNAND2X1_LOC_352 NAND2X1_LOC_352/a_36_24# INVX1_LOC_286/A VSS VDD INVX1_LOC_160/Y
+ INVX1_LOC_271/Y NAND2X1_LOC
XNAND2X1_LOC_363 NAND2X1_LOC_363/a_36_24# INVX1_LOC_297/A VSS VDD INVX1_LOC_293/Y
+ INVX1_LOC_294/Y NAND2X1_LOC
XNAND2X1_LOC_341 NAND2X1_LOC_341/a_36_24# INVX1_LOC_275/A VSS VDD INVX1_LOC_202/Y
+ INVX1_LOC_203/Y NAND2X1_LOC
XNAND2X1_LOC_385 NAND2X1_LOC_385/a_36_24# NAND2X1_LOC_537/A VSS VDD INVX1_LOC_35/Y
+ INVX1_LOC_100/Y NAND2X1_LOC
XNAND2X1_LOC_396 NAND2X1_LOC_396/a_36_24# NAND2X1_LOC_396/Y VSS VDD INVX1_LOC_32/Y
+ INVX1_LOC_45/Y NAND2X1_LOC
XINVX1_LOC_207 INVX1_LOC_207/Y VSS VDD INVX1_LOC_207/A INVX1_LOC
XINVX1_LOC_218 INVX1_LOC_218/Y VSS VDD INVX1_LOC_218/A INVX1_LOC
XINVX1_LOC_229 INVX1_LOC_229/Y VSS VDD INVX1_LOC_223/Y INVX1_LOC
XNAND2X1_LOC_160 NAND2X1_LOC_160/a_36_24# INVX1_LOC_147/A VSS VDD INVX1_LOC_148/Y
+ INVX1_LOC_149/Y NAND2X1_LOC
XNAND2X1_LOC_182 NAND2X1_LOC_182/a_36_24# INVX1_LOC_160/A VSS VDD INVX1_LOC_158/Y
+ INVX1_LOC_159/Y NAND2X1_LOC
XNAND2X1_LOC_171 NAND2X1_LOC_171/a_36_24# NAND2X1_LOC_333/A VSS VDD INVX1_LOC_32/Y
+ INVX1_LOC_48/Y NAND2X1_LOC
XNAND2X1_LOC_193 NAND2X1_LOC_193/a_36_24# INVX1_LOC_169/A VSS VDD NAND2X1_LOC_7/Y
+ NAND2X1_LOC_13/Y NAND2X1_LOC
XNAND2X1_LOC_18 NAND2X1_LOC_18/a_36_24# INVX1_LOC_26/A VSS VDD INVX1_LOC_18/Y INVX1_LOC_25/Y
+ NAND2X1_LOC
XNAND2X1_LOC_29 NAND2X1_LOC_29/a_36_24# INVX1_LOC_38/A VSS VDD INVX1_LOC_12/Y INVX1_LOC_39/Y
+ NAND2X1_LOC
XINVX1_LOC_571 INVX1_LOC_571/Y VSS VDD INVX1_LOC_571/A INVX1_LOC
XINVX1_LOC_582 INVX1_LOC_582/Y VSS VDD INVX1_LOC_582/A INVX1_LOC
XINVX1_LOC_593 INVX1_LOC_593/Y VSS VDD INVX1_LOC_259/Y INVX1_LOC
XINVX1_LOC_560 INVX1_LOC_560/Y VSS VDD INVX1_LOC_560/A INVX1_LOC
XNAND2X1_LOC_704 NAND2X1_LOC_704/a_36_24# INVX1_LOC_546/A VSS VDD NAND2X1_LOC_317/A
+ NAND2X1_LOC_704/B NAND2X1_LOC
XNAND2X1_LOC_715 NAND2X1_LOC_715/a_36_24# INVX1_LOC_558/A VSS VDD INVX1_LOC_105/Y
+ INVX1_LOC_544/Y NAND2X1_LOC
XNAND2X1_LOC_726 NAND2X1_LOC_726/a_36_24# INVX1_LOC_569/A VSS VDD NAND2X1_LOC_152/Y
+ INVX1_LOC_554/Y NAND2X1_LOC
XNAND2X1_LOC_737 NAND2X1_LOC_737/a_36_24# INVX1_LOC_580/A VSS VDD INVX1_LOC_576/Y
+ INVX1_LOC_577/Y NAND2X1_LOC
XNAND2X1_LOC_759 NAND2X1_LOC_759/a_36_24# NAND2X1_LOC_759/Y VSS VDD INVX1_LOC_206/Y
+ NAND2X1_LOC_759/B NAND2X1_LOC
XNAND2X1_LOC_748 NAND2X1_LOC_748/a_36_24# NAND2X1_LOC_789/A VSS VDD INVX1_LOC_7/Y
+ INVX1_LOC_543/Y NAND2X1_LOC
XINVX1_LOC_390 INVX1_LOC_390/Y VSS VDD INVX1_LOC_390/A INVX1_LOC
XNAND2X1_LOC_567 NAND2X1_LOC_567/a_36_24# INVX1_LOC_441/A VSS VDD INVX1_LOC_409/Y
+ INVX1_LOC_412/Y NAND2X1_LOC
XNAND2X1_LOC_501 NAND2X1_LOC_501/a_36_24# INVX1_LOC_393/A VSS VDD NAND2X1_LOC_498/Y
+ INVX1_LOC_392/Y NAND2X1_LOC
XNAND2X1_LOC_534 NAND2X1_LOC_534/a_36_24# NAND2X1_LOC_534/Y VSS VDD INVX1_LOC_49/Y
+ INVX1_LOC_63/Y NAND2X1_LOC
XNAND2X1_LOC_556 NAND2X1_LOC_556/a_36_24# INVX1_LOC_430/A VSS VDD INVX1_LOC_386/Y
+ INVX1_LOC_387/Y NAND2X1_LOC
XNAND2X1_LOC_523 NAND2X1_LOC_523/a_36_24# INVX1_LOC_406/A VSS VDD NAND2X1_LOC_521/Y
+ NAND2X1_LOC_523/B NAND2X1_LOC
XNAND2X1_LOC_589 NAND2X1_LOC_589/a_36_24# NAND2X1_LOC_592/B VSS VDD INVX1_LOC_31/Y
+ INVX1_LOC_119/Y NAND2X1_LOC
XNAND2X1_LOC_512 NAND2X1_LOC_512/a_36_24# INVX1_LOC_401/A VSS VDD INPUT_0 NAND2X1_LOC_308/A
+ NAND2X1_LOC
XNAND2X1_LOC_578 NAND2X1_LOC_578/a_36_24# INVX1_LOC_452/A VSS VDD INVX1_LOC_442/Y
+ INVX1_LOC_451/Y NAND2X1_LOC
XNAND2X1_LOC_545 NAND2X1_LOC_545/a_36_24# INVX1_LOC_419/A VSS VDD NAND2X1_LOC_545/A
+ NAND2X1_LOC_545/B NAND2X1_LOC
XNAND2X1_LOC_320 NAND2X1_LOC_320/a_36_24# NAND2X1_LOC_320/Y VSS VDD INVX1_LOC_45/Y
+ INVX1_LOC_89/Y NAND2X1_LOC
XNAND2X1_LOC_331 NAND2X1_LOC_331/a_36_24# NAND2X1_LOC_331/Y VSS VDD NAND2X1_LOC_331/A
+ NAND2X1_LOC_331/B NAND2X1_LOC
XNAND2X1_LOC_342 NAND2X1_LOC_342/a_36_24# INVX1_LOC_276/A VSS VDD NAND2X1_LOC_342/A
+ NAND2X1_LOC_342/B NAND2X1_LOC
XNAND2X1_LOC_353 NAND2X1_LOC_353/a_36_24# INVX1_LOC_287/A VSS VDD INVX1_LOC_250/Y
+ INVX1_LOC_252/Y NAND2X1_LOC
XNAND2X1_LOC_386 NAND2X1_LOC_386/a_36_24# INVX1_LOC_315/A VSS VDD INVX1_LOC_316/Y
+ INVX1_LOC_25/Y NAND2X1_LOC
XNAND2X1_LOC_364 NAND2X1_LOC_364/a_36_24# INVX1_LOC_298/A VSS VDD INVX1_LOC_291/Y
+ INVX1_LOC_292/Y NAND2X1_LOC
XNAND2X1_LOC_375 NAND2X1_LOC_375/a_36_24# NAND2X1_LOC_376/B VSS VDD INVX1_LOC_305/Y
+ INVX1_LOC_306/Y NAND2X1_LOC
XNAND2X1_LOC_397 NAND2X1_LOC_397/a_36_24# NAND2X1_LOC_397/Y VSS VDD INVX1_LOC_6/Y
+ INVX1_LOC_83/Y NAND2X1_LOC
XINVX1_LOC_219 INVX1_LOC_219/Y VSS VDD INVX1_LOC_7/Y INVX1_LOC
XINVX1_LOC_208 INVX1_LOC_208/Y VSS VDD INVX1_LOC_208/A INVX1_LOC
XNAND2X1_LOC_161 NAND2X1_LOC_161/a_36_24# INVX1_LOC_150/A VSS VDD INVX1_LOC_151/Y
+ INVX1_LOC_152/Y NAND2X1_LOC
XNAND2X1_LOC_150 NAND2X1_LOC_150/a_36_24# INVX1_LOC_134/A VSS VDD INVX1_LOC_46/Y INVX1_LOC_65/Y
+ NAND2X1_LOC
XNAND2X1_LOC_19 NAND2X1_LOC_19/a_36_24# INVX1_LOC_27/A VSS VDD INVX1_LOC_28/Y INVX1_LOC_9/Y
+ NAND2X1_LOC
XNAND2X1_LOC_172 NAND2X1_LOC_172/a_36_24# NAND2X1_LOC_174/B VSS VDD INVX1_LOC_74/Y
+ INVX1_LOC_99/Y NAND2X1_LOC
XNAND2X1_LOC_183 NAND2X1_LOC_183/a_36_24# NAND2X1_LOC_190/A VSS VDD INVX1_LOC_11/Y
+ INVX1_LOC_48/Y NAND2X1_LOC
XNAND2X1_LOC_194 NAND2X1_LOC_194/a_36_24# INVX1_LOC_170/A VSS VDD NAND2X1_LOC_16/Y
+ NAND2X1_LOC_39/Y NAND2X1_LOC
XINVX1_LOC_583 INVX1_LOC_583/Y VSS VDD INVX1_LOC_583/A INVX1_LOC
XINVX1_LOC_550 INVX1_LOC_550/Y VSS VDD INVX1_LOC_550/A INVX1_LOC
XINVX1_LOC_572 INVX1_LOC_572/Y VSS VDD INVX1_LOC_572/A INVX1_LOC
XINVX1_LOC_594 INVX1_LOC_594/Y VSS VDD INPUT_0 INVX1_LOC
XINVX1_LOC_561 INVX1_LOC_561/Y VSS VDD INVX1_LOC_561/A INVX1_LOC
XNAND2X1_LOC_727 NAND2X1_LOC_727/a_36_24# INVX1_LOC_570/A VSS VDD INVX1_LOC_252/Y
+ INVX1_LOC_350/Y NAND2X1_LOC
XNAND2X1_LOC_705 NAND2X1_LOC_705/a_36_24# INVX1_LOC_547/A VSS VDD NAND2X1_LOC_486/B
+ NAND2X1_LOC_526/Y NAND2X1_LOC
XNAND2X1_LOC_738 NAND2X1_LOC_738/a_36_24# INVX1_LOC_581/A VSS VDD INVX1_LOC_574/Y
+ INVX1_LOC_575/Y NAND2X1_LOC
XNAND2X1_LOC_716 NAND2X1_LOC_716/a_36_24# INVX1_LOC_559/A VSS VDD INVX1_LOC_202/Y
+ INVX1_LOC_248/Y NAND2X1_LOC
XNAND2X1_LOC_749 NAND2X1_LOC_749/a_36_24# NAND2X1_LOC_749/Y VSS VDD INVX1_LOC_585/Y
+ INVX1_LOC_12/Y NAND2X1_LOC
XINVX1_LOC_391 INVX1_LOC_391/Y VSS VDD INVX1_LOC_391/A INVX1_LOC
XINVX1_LOC_380 INVX1_LOC_380/Y VSS VDD INVX1_LOC_380/A INVX1_LOC
XNAND2X1_LOC_502 NAND2X1_LOC_502/a_36_24# NAND2X1_LOC_503/B VSS VDD INVX1_LOC_394/Y
+ INVX1_LOC_395/Y NAND2X1_LOC
XNAND2X1_LOC_535 NAND2X1_LOC_535/a_36_24# INVX1_LOC_409/A VSS VDD NAND2X1_LOC_788/A
+ NAND2X1_LOC_534/Y NAND2X1_LOC
XNAND2X1_LOC_546 NAND2X1_LOC_546/a_36_24# INVX1_LOC_420/A VSS VDD NAND2X1_LOC_525/Y
+ NAND2X1_LOC_526/Y NAND2X1_LOC
XNAND2X1_LOC_513 NAND2X1_LOC_513/a_36_24# NAND2X1_LOC_513/Y VSS VDD NAND2X1_LOC_513/A
+ INVX1_LOC_401/Y NAND2X1_LOC
XNAND2X1_LOC_579 NAND2X1_LOC_579/a_36_24# INVX1_LOC_453/A VSS VDD INVX1_LOC_449/Y
+ INVX1_LOC_450/Y NAND2X1_LOC
XNAND2X1_LOC_568 NAND2X1_LOC_568/a_36_24# INVX1_LOC_442/A VSS VDD INVX1_LOC_440/Y
+ INVX1_LOC_441/Y NAND2X1_LOC
XNAND2X1_LOC_524 NAND2X1_LOC_524/a_36_24# NAND2X1_LOC_545/B VSS VDD INVX1_LOC_53/Y
+ INVX1_LOC_479/A NAND2X1_LOC
XNAND2X1_LOC_557 NAND2X1_LOC_557/a_36_24# INVX1_LOC_431/A VSS VDD INVX1_LOC_388/Y
+ NAND2X1_LOC_557/B NAND2X1_LOC
XNAND2X1_LOC_332 NAND2X1_LOC_332/a_36_24# INVX1_LOC_266/A VSS VDD NAND2X1_LOC_111/Y
+ NAND2X1_LOC_332/B NAND2X1_LOC
XNAND2X1_LOC_354 NAND2X1_LOC_354/a_36_24# INVX1_LOC_288/A VSS VDD INVX1_LOC_255/Y
+ INVX1_LOC_258/Y NAND2X1_LOC
XNAND2X1_LOC_321 NAND2X1_LOC_321/a_36_24# NAND2X1_LOC_324/B VSS VDD INVX1_LOC_17/Y
+ INVX1_LOC_69/Y NAND2X1_LOC
XNAND2X1_LOC_343 NAND2X1_LOC_343/a_36_24# INVX1_LOC_277/A VSS VDD NAND2X1_LOC_250/Y
+ NAND2X1_LOC_843/A NAND2X1_LOC
XNAND2X1_LOC_310 NAND2X1_LOC_310/a_36_24# NAND2X1_LOC_335/B VSS VDD INVX1_LOC_9/Y
+ INVX1_LOC_48/Y NAND2X1_LOC
XNAND2X1_LOC_365 NAND2X1_LOC_365/a_36_24# INVX1_LOC_299/A VSS VDD INVX1_LOC_290/Y
+ INVX1_LOC_298/Y NAND2X1_LOC
XNAND2X1_LOC_387 NAND2X1_LOC_387/a_36_24# NAND2X1_LOC_387/Y VSS VDD INVX1_LOC_90/Y
+ INVX1_LOC_315/Y NAND2X1_LOC
XNAND2X1_LOC_376 NAND2X1_LOC_376/a_36_24# NAND2X1_LOC_376/Y VSS VDD INVX1_LOC_395/A
+ NAND2X1_LOC_376/B NAND2X1_LOC
XNAND2X1_LOC_398 NAND2X1_LOC_398/a_36_24# NAND2X1_LOC_399/B VSS VDD INVX1_LOC_322/Y
+ INVX1_LOC_323/Y NAND2X1_LOC
XINVX1_LOC_209 INVX1_LOC_209/Y VSS VDD INVX1_LOC_209/A INVX1_LOC
XNAND2X1_LOC_173 NAND2X1_LOC_173/a_36_24# NAND2X1_LOC_173/Y VSS VDD INVX1_LOC_74/Y
+ INVX1_LOC_134/Y NAND2X1_LOC
XNAND2X1_LOC_184 NAND2X1_LOC_184/a_36_24# NAND2X1_LOC_184/Y VSS VDD INVX1_LOC_75/Y
+ INVX1_LOC_93/Y NAND2X1_LOC
XNAND2X1_LOC_140 NAND2X1_LOC_140/a_36_24# INVX1_LOC_127/A VSS VDD INVX1_LOC_118/Y
+ NAND2X1_LOC_140/B NAND2X1_LOC
XNAND2X1_LOC_162 NAND2X1_LOC_162/a_36_24# NAND2X1_LOC_163/B VSS VDD INVX1_LOC_147/Y
+ INVX1_LOC_150/Y NAND2X1_LOC
XNAND2X1_LOC_151 NAND2X1_LOC_151/a_36_24# NAND2X1_LOC_152/B VSS VDD INVX1_LOC_135/Y
+ INVX1_LOC_136/Y NAND2X1_LOC
XNAND2X1_LOC_195 NAND2X1_LOC_195/a_36_24# INVX1_LOC_171/A VSS VDD NAND2X1_LOC_41/Y
+ NAND2X1_LOC_43/Y NAND2X1_LOC
XINVX1_LOC_573 INVX1_LOC_573/Y VSS VDD INVX1_LOC_573/A INVX1_LOC
XINVX1_LOC_540 INVX1_LOC_540/Y VSS VDD INVX1_LOC_245/A INVX1_LOC
XINVX1_LOC_584 INVX1_LOC_584/Y VSS VDD INVX1_LOC_584/A INVX1_LOC
XINVX1_LOC_562 INVX1_LOC_562/Y VSS VDD INVX1_LOC_562/A INVX1_LOC
XINVX1_LOC_551 INVX1_LOC_551/Y VSS VDD INVX1_LOC_551/A INVX1_LOC
XINVX1_LOC_595 INVX1_LOC_595/Y VSS VDD INVX1_LOC_595/A INVX1_LOC
XINVX1_LOC_370 INVX1_LOC_370/Y VSS VDD INVX1_LOC_370/A INVX1_LOC
XNAND2X1_LOC_706 NAND2X1_LOC_706/a_36_24# INVX1_LOC_548/A VSS VDD NAND2X1_LOC_692/Y
+ NAND2X1_LOC_706/B NAND2X1_LOC
XNAND2X1_LOC_728 NAND2X1_LOC_728/a_36_24# INVX1_LOC_571/A VSS VDD NAND2X1_LOC_728/A
+ NAND2X1_LOC_728/B NAND2X1_LOC
XNAND2X1_LOC_739 NAND2X1_LOC_739/a_36_24# INVX1_LOC_582/A VSS VDD INVX1_LOC_168/Y
+ INVX1_LOC_573/Y NAND2X1_LOC
XNAND2X1_LOC_717 NAND2X1_LOC_717/a_36_24# INVX1_LOC_560/A VSS VDD INVX1_LOC_304/Y
+ INVX1_LOC_390/Y NAND2X1_LOC
XINVX1_LOC_392 INVX1_LOC_392/Y VSS VDD INVX1_LOC_392/A INVX1_LOC
XINVX1_LOC_381 INVX1_LOC_381/Y VSS VDD INVX1_LOC_381/A INVX1_LOC
XNAND2X1_LOC_525 NAND2X1_LOC_525/a_36_24# NAND2X1_LOC_525/Y VSS VDD INVX1_LOC_17/Y
+ INVX1_LOC_58/Y NAND2X1_LOC
XNAND2X1_LOC_514 NAND2X1_LOC_514/a_36_24# INVX1_LOC_402/A VSS VDD INVX1_LOC_403/Y
+ NAND2X1_LOC_136/Y NAND2X1_LOC
XNAND2X1_LOC_536 NAND2X1_LOC_536/a_36_24# NAND2X1_LOC_537/B VSS VDD INVX1_LOC_20/Y
+ INVX1_LOC_99/Y NAND2X1_LOC
XNAND2X1_LOC_503 NAND2X1_LOC_503/a_36_24# NAND2X1_LOC_503/Y VSS VDD INVX1_LOC_69/Y
+ NAND2X1_LOC_503/B NAND2X1_LOC
XNAND2X1_LOC_569 NAND2X1_LOC_569/a_36_24# INVX1_LOC_443/A VSS VDD INVX1_LOC_438/Y
+ INVX1_LOC_439/Y NAND2X1_LOC
XNAND2X1_LOC_547 NAND2X1_LOC_547/a_36_24# INVX1_LOC_421/A VSS VDD NAND2X1_LOC_527/Y
+ NAND2X1_LOC_528/Y NAND2X1_LOC
XNAND2X1_LOC_558 NAND2X1_LOC_558/a_36_24# INVX1_LOC_432/A VSS VDD INVX1_LOC_390/Y
+ NAND2X1_LOC_558/B NAND2X1_LOC
XNAND2X1_LOC_322 NAND2X1_LOC_322/a_36_24# NAND2X1_LOC_322/Y VSS VDD INVX1_LOC_50/Y
+ INVX1_LOC_395/A NAND2X1_LOC
XNAND2X1_LOC_355 NAND2X1_LOC_355/a_36_24# INVX1_LOC_289/A VSS VDD NAND2X1_LOC_355/A
+ NAND2X1_LOC_331/Y NAND2X1_LOC
XNAND2X1_LOC_300 NAND2X1_LOC_300/a_36_24# NAND2X1_LOC_301/B VSS VDD INVX1_LOC_63/Y
+ INVX1_LOC_114/A NAND2X1_LOC
XNAND2X1_LOC_344 NAND2X1_LOC_344/a_36_24# INVX1_LOC_278/A VSS VDD INVX1_LOC_217/Y
+ NAND2X1_LOC_344/B NAND2X1_LOC
XNAND2X1_LOC_311 NAND2X1_LOC_311/a_36_24# NAND2X1_LOC_538/B VSS VDD INVX1_LOC_35/Y
+ INVX1_LOC_99/Y NAND2X1_LOC
XNAND2X1_LOC_366 NAND2X1_LOC_366/a_36_24# INVX1_LOC_300/A VSS VDD INVX1_LOC_296/Y
+ INVX1_LOC_297/Y NAND2X1_LOC
XNAND2X1_LOC_333 NAND2X1_LOC_333/a_36_24# INVX1_LOC_267/A VSS VDD NAND2X1_LOC_333/A
+ NAND2X1_LOC_333/B NAND2X1_LOC
XNAND2X1_LOC_377 NAND2X1_LOC_377/a_36_24# INVX1_LOC_307/A VSS VDD INVX1_LOC_6/Y INVX1_LOC_308/Y
+ NAND2X1_LOC
XNAND2X1_LOC_388 NAND2X1_LOC_388/a_36_24# INVX1_LOC_317/A VSS VDD NAND2X1_LOC_388/A
+ NAND2X1_LOC_176/Y NAND2X1_LOC
XNAND2X1_LOC_399 NAND2X1_LOC_399/a_36_24# NAND2X1_LOC_403/A VSS VDD INVX1_LOC_50/Y
+ NAND2X1_LOC_399/B NAND2X1_LOC
XNAND2X1_LOC_141 NAND2X1_LOC_141/a_36_24# INVX1_LOC_128/A VSS VDD INVX1_LOC_126/Y
+ INVX1_LOC_127/Y NAND2X1_LOC
XNAND2X1_LOC_130 NAND2X1_LOC_130/a_36_24# NAND2X1_LOC_130/Y VSS VDD INVX1_LOC_121/Y
+ INVX1_LOC_122/Y NAND2X1_LOC
XNAND2X1_LOC_185 NAND2X1_LOC_185/a_36_24# INVX1_LOC_161/A VSS VDD INVX1_LOC_162/Y
+ INVX1_LOC_163/Y NAND2X1_LOC
XNAND2X1_LOC_163 NAND2X1_LOC_163/a_36_24# NAND2X1_LOC_467/A VSS VDD INVX1_LOC_58/Y
+ NAND2X1_LOC_163/B NAND2X1_LOC
XNAND2X1_LOC_152 NAND2X1_LOC_152/a_36_24# NAND2X1_LOC_152/Y VSS VDD INVX1_LOC_53/Y
+ NAND2X1_LOC_152/B NAND2X1_LOC
XNAND2X1_LOC_174 NAND2X1_LOC_174/a_36_24# INVX1_LOC_156/A VSS VDD NAND2X1_LOC_333/A
+ NAND2X1_LOC_174/B NAND2X1_LOC
XNAND2X1_LOC_196 NAND2X1_LOC_196/a_36_24# INVX1_LOC_172/A VSS VDD NAND2X1_LOC_45/Y
+ NAND2X1_LOC_48/Y NAND2X1_LOC
XINVX1_LOC_541 INVX1_LOC_541/Y VSS VDD INPUT_0 INVX1_LOC
XINVX1_LOC_563 INVX1_LOC_563/Y VSS VDD INVX1_LOC_563/A INVX1_LOC
XINVX1_LOC_552 INVX1_LOC_552/Y VSS VDD INVX1_LOC_543/Y INVX1_LOC
XINVX1_LOC_530 INVX1_LOC_530/Y VSS VDD INVX1_LOC_530/A INVX1_LOC
XINVX1_LOC_574 INVX1_LOC_574/Y VSS VDD INVX1_LOC_574/A INVX1_LOC
XINVX1_LOC_596 INVX1_LOC_596/Y VSS VDD INVX1_LOC_596/A INVX1_LOC
XINVX1_LOC_585 INVX1_LOC_585/Y VSS VDD INPUT_0 INVX1_LOC
XNAND2X1_LOC_718 NAND2X1_LOC_718/a_36_24# INVX1_LOC_561/A VSS VDD NAND2X1_LOC_591/Y
+ INVX1_LOC_469/Y NAND2X1_LOC
XNAND2X1_LOC_707 NAND2X1_LOC_707/a_36_24# INVX1_LOC_549/A VSS VDD NAND2X1_LOC_707/A
+ NAND2X1_LOC_707/B NAND2X1_LOC
XINVX1_LOC_371 INVX1_LOC_371/Y VSS VDD INVX1_LOC_371/A INVX1_LOC
XINVX1_LOC_393 INVX1_LOC_393/Y VSS VDD INVX1_LOC_393/A INVX1_LOC
XINVX1_LOC_360 INVX1_LOC_360/Y VSS VDD INVX1_LOC_360/A INVX1_LOC
XINVX1_LOC_382 INVX1_LOC_382/Y VSS VDD INVX1_LOC_382/A INVX1_LOC
XNAND2X1_LOC_729 NAND2X1_LOC_729/a_36_24# INVX1_LOC_572/A VSS VDD INVX1_LOC_538/Y
+ INVX1_LOC_542/Y NAND2X1_LOC
XNAND2X1_LOC_526 NAND2X1_LOC_526/a_36_24# NAND2X1_LOC_526/Y VSS VDD INVX1_LOC_41/Y
+ INVX1_LOC_586/A NAND2X1_LOC
XNAND2X1_LOC_515 NAND2X1_LOC_515/a_36_24# NAND2X1_LOC_516/B VSS VDD NAND2X1_LOC_704/B
+ INVX1_LOC_402/Y NAND2X1_LOC
XNAND2X1_LOC_559 NAND2X1_LOC_559/a_36_24# INVX1_LOC_433/A VSS VDD NAND2X1_LOC_517/Y
+ INVX1_LOC_405/Y NAND2X1_LOC
XNAND2X1_LOC_548 NAND2X1_LOC_548/a_36_24# INVX1_LOC_422/A VSS VDD NAND2X1_LOC_529/Y
+ NAND2X1_LOC_548/B NAND2X1_LOC
XNAND2X1_LOC_504 NAND2X1_LOC_504/a_36_24# NAND2X1_LOC_507/A VSS VDD INVX1_LOC_17/Y
+ INVX1_LOC_145/Y NAND2X1_LOC
XNAND2X1_LOC_537 NAND2X1_LOC_537/a_36_24# INVX1_LOC_410/A VSS VDD NAND2X1_LOC_537/A
+ NAND2X1_LOC_537/B NAND2X1_LOC
XINVX1_LOC_190 INVX1_LOC_190/Y VSS VDD INVX1_LOC_190/A INVX1_LOC
XNAND2X1_LOC_356 NAND2X1_LOC_356/a_36_24# INVX1_LOC_290/A VSS VDD INVX1_LOC_288/Y
+ INVX1_LOC_289/Y NAND2X1_LOC
XNAND2X1_LOC_345 NAND2X1_LOC_345/a_36_24# INVX1_LOC_279/A VSS VDD INVX1_LOC_220/Y
+ NAND2X1_LOC_261/Y NAND2X1_LOC
XNAND2X1_LOC_323 NAND2X1_LOC_323/a_36_24# NAND2X1_LOC_325/B VSS VDD INVX1_LOC_93/Y
+ INVX1_LOC_103/Y NAND2X1_LOC
XNAND2X1_LOC_301 NAND2X1_LOC_301/a_36_24# INVX1_LOC_248/A VSS VDD NAND2X1_LOC_76/B
+ NAND2X1_LOC_301/B NAND2X1_LOC
XNAND2X1_LOC_312 NAND2X1_LOC_312/a_36_24# NAND2X1_LOC_336/B VSS VDD INVX1_LOC_62/Y
+ INVX1_LOC_69/Y NAND2X1_LOC
XNAND2X1_LOC_367 NAND2X1_LOC_367/a_36_24# GATE_366 VSS VDD INVX1_LOC_299/Y INVX1_LOC_300/Y
+ NAND2X1_LOC
XNAND2X1_LOC_334 NAND2X1_LOC_334/a_36_24# INVX1_LOC_268/A VSS VDD NAND2X1_LOC_334/A
+ NAND2X1_LOC_334/B NAND2X1_LOC
XNAND2X1_LOC_389 NAND2X1_LOC_389/a_36_24# INVX1_LOC_318/A VSS VDD NAND2X1_LOC_537/A
+ NAND2X1_LOC_387/Y NAND2X1_LOC
XNAND2X1_LOC_378 NAND2X1_LOC_378/a_36_24# NAND2X1_LOC_378/Y VSS VDD INVX1_LOC_309/Y
+ INVX1_LOC_307/Y NAND2X1_LOC
XNAND2X1_LOC_120 NAND2X1_LOC_120/a_36_24# INVX1_LOC_111/A VSS VDD INVX1_LOC_112/Y
+ INVX1_LOC_113/Y NAND2X1_LOC
XNAND2X1_LOC_131 NAND2X1_LOC_131/a_36_24# NAND2X1_LOC_140/B VSS VDD INVX1_LOC_20/Y
+ NAND2X1_LOC_130/Y NAND2X1_LOC
XNAND2X1_LOC_186 NAND2X1_LOC_186/a_36_24# NAND2X1_LOC_331/A VSS VDD INVX1_LOC_164/Y
+ INVX1_LOC_588/A NAND2X1_LOC
XNAND2X1_LOC_142 NAND2X1_LOC_142/a_36_24# NAND2X1_LOC_142/Y VSS VDD INVX1_LOC_54/Y
+ INVX1_LOC_69/Y NAND2X1_LOC
XNAND2X1_LOC_153 NAND2X1_LOC_153/a_36_24# INVX1_LOC_137/A VSS VDD INVX1_LOC_138/Y
+ INVX1_LOC_46/Y NAND2X1_LOC
XNAND2X1_LOC_175 NAND2X1_LOC_175/a_36_24# INVX1_LOC_157/A VSS VDD NAND2X1_LOC_173/Y
+ INVX1_LOC_156/Y NAND2X1_LOC
XNAND2X1_LOC_197 NAND2X1_LOC_197/a_36_24# INVX1_LOC_173/A VSS VDD NAND2X1_LOC_52/Y
+ NAND2X1_LOC_56/Y NAND2X1_LOC
XNAND2X1_LOC_164 NAND2X1_LOC_164/a_36_24# NAND2X1_LOC_164/Y VSS VDD INVX1_LOC_26/Y
+ INVX1_LOC_395/A NAND2X1_LOC
XINVX1_LOC_575 INVX1_LOC_575/Y VSS VDD INVX1_LOC_575/A INVX1_LOC
XINVX1_LOC_542 INVX1_LOC_542/Y VSS VDD INVX1_LOC_542/A INVX1_LOC
XINVX1_LOC_520 INVX1_LOC_520/Y VSS VDD INVX1_LOC_520/A INVX1_LOC
XINVX1_LOC_553 INVX1_LOC_553/Y VSS VDD INVX1_LOC_553/A INVX1_LOC
XINVX1_LOC_564 INVX1_LOC_564/Y VSS VDD INVX1_LOC_564/A INVX1_LOC
XINVX1_LOC_531 INVX1_LOC_531/Y VSS VDD INVX1_LOC_531/A INVX1_LOC
XINVX1_LOC_586 INVX1_LOC_586/Y VSS VDD INVX1_LOC_586/A INVX1_LOC
XINVX1_LOC_597 INVX1_LOC_597/Y VSS VDD INVX1_LOC_597/A INVX1_LOC
XNAND2X1_LOC_708 NAND2X1_LOC_708/a_36_24# INVX1_LOC_550/A VSS VDD NAND2X1_LOC_708/A
+ NAND2X1_LOC_697/Y NAND2X1_LOC
XNAND2X1_LOC_719 NAND2X1_LOC_719/a_36_24# INVX1_LOC_562/A VSS VDD NAND2X1_LOC_719/A
+ NAND2X1_LOC_666/Y NAND2X1_LOC
XINVX1_LOC_383 INVX1_LOC_383/Y VSS VDD INVX1_LOC_383/A INVX1_LOC
XINVX1_LOC_372 INVX1_LOC_372/Y VSS VDD INVX1_LOC_372/A INVX1_LOC
XINVX1_LOC_350 INVX1_LOC_350/Y VSS VDD INVX1_LOC_350/A INVX1_LOC
XINVX1_LOC_361 INVX1_LOC_361/Y VSS VDD INVX1_LOC_361/A INVX1_LOC
XINVX1_LOC_394 INVX1_LOC_394/Y VSS VDD INVX1_LOC_80/A INVX1_LOC
XNAND2X1_LOC_516 NAND2X1_LOC_516/a_36_24# NAND2X1_LOC_516/Y VSS VDD NAND2X1_LOC_513/Y
+ NAND2X1_LOC_516/B NAND2X1_LOC
XNAND2X1_LOC_527 NAND2X1_LOC_527/a_36_24# NAND2X1_LOC_527/Y VSS VDD INVX1_LOC_69/Y
+ INVX1_LOC_103/Y NAND2X1_LOC
XNAND2X1_LOC_538 NAND2X1_LOC_538/a_36_24# INVX1_LOC_411/A VSS VDD NAND2X1_LOC_13/Y
+ NAND2X1_LOC_538/B NAND2X1_LOC
XNAND2X1_LOC_549 NAND2X1_LOC_549/a_36_24# INVX1_LOC_423/A VSS VDD NAND2X1_LOC_531/Y
+ INVX1_LOC_422/Y NAND2X1_LOC
XNAND2X1_LOC_505 NAND2X1_LOC_505/a_36_24# NAND2X1_LOC_505/Y VSS VDD INVX1_LOC_26/Y
+ INVX1_LOC_32/Y NAND2X1_LOC
XINVX1_LOC_180 INVX1_LOC_180/Y VSS VDD INVX1_LOC_180/A INVX1_LOC
XINVX1_LOC_191 INVX1_LOC_191/Y VSS VDD INVX1_LOC_191/A INVX1_LOC
XNAND2X1_LOC_302 NAND2X1_LOC_302/a_36_24# INVX1_LOC_249/A VSS VDD NAND2X1_LOC_302/A
+ NAND2X1_LOC_299/Y NAND2X1_LOC
XNAND2X1_LOC_324 NAND2X1_LOC_324/a_36_24# INVX1_LOC_256/A VSS VDD NAND2X1_LOC_320/Y
+ NAND2X1_LOC_324/B NAND2X1_LOC
XNAND2X1_LOC_313 NAND2X1_LOC_313/a_36_24# NAND2X1_LOC_317/A VSS VDD INVX1_LOC_74/Y
+ INVX1_LOC_89/Y NAND2X1_LOC
XNAND2X1_LOC_346 NAND2X1_LOC_346/a_36_24# INVX1_LOC_280/A VSS VDD NAND2X1_LOC_292/Y
+ NAND2X1_LOC_346/B NAND2X1_LOC
XNAND2X1_LOC_368 NAND2X1_LOC_368/a_36_24# NAND2X1_LOC_457/A VSS VDD INVX1_LOC_11/Y
+ NAND2X1_LOC_271/B NAND2X1_LOC
XNAND2X1_LOC_335 NAND2X1_LOC_335/a_36_24# INVX1_LOC_269/A VSS VDD NAND2X1_LOC_370/A
+ NAND2X1_LOC_335/B NAND2X1_LOC
XNAND2X1_LOC_357 NAND2X1_LOC_357/a_36_24# INVX1_LOC_291/A VSS VDD INVX1_LOC_286/Y
+ INVX1_LOC_287/Y NAND2X1_LOC
XNAND2X1_LOC_379 NAND2X1_LOC_379/a_36_24# NAND2X1_LOC_379/Y VSS VDD INVX1_LOC_310/Y
+ INVX1_LOC_311/Y NAND2X1_LOC
XNAND2X1_LOC_132 NAND2X1_LOC_132/a_36_24# NAND2X1_LOC_137/A VSS VDD INVX1_LOC_89/Y
+ INVX1_LOC_93/Y NAND2X1_LOC
XNAND2X1_LOC_110 NAND2X1_LOC_110/a_36_24# INVX1_LOC_103/A VSS VDD INVX1_LOC_104/Y
+ INVX1_LOC_21/Y NAND2X1_LOC
XNAND2X1_LOC_121 NAND2X1_LOC_121/a_36_24# NAND2X1_LOC_121/Y VSS VDD INVX1_LOC_114/Y
+ INVX1_LOC_526/A NAND2X1_LOC
XNAND2X1_LOC_143 NAND2X1_LOC_143/a_36_24# INVX1_LOC_129/A VSS VDD INVX1_LOC_130/Y
+ INVX1_LOC_12/Y NAND2X1_LOC
XNAND2X1_LOC_187 NAND2X1_LOC_187/a_36_24# NAND2X1_LOC_187/Y VSS VDD INVX1_LOC_48/Y
+ NAND2X1_LOC_331/A NAND2X1_LOC
XNAND2X1_LOC_154 NAND2X1_LOC_154/a_36_24# INVX1_LOC_139/A VSS VDD INVX1_LOC_140/Y
+ INVX1_LOC_141/Y NAND2X1_LOC
XNAND2X1_LOC_176 NAND2X1_LOC_176/a_36_24# NAND2X1_LOC_176/Y VSS VDD INVX1_LOC_35/Y
+ INVX1_LOC_89/Y NAND2X1_LOC
XNAND2X1_LOC_165 NAND2X1_LOC_165/a_36_24# NAND2X1_LOC_165/Y VSS VDD INVX1_LOC_58/Y
+ INVX1_LOC_76/Y NAND2X1_LOC
XNAND2X1_LOC_198 NAND2X1_LOC_198/a_36_24# INVX1_LOC_174/A VSS VDD NAND2X1_LOC_57/Y
+ INVX1_LOC_173/Y NAND2X1_LOC
XINVX1_LOC_554 INVX1_LOC_554/Y VSS VDD INVX1_LOC_554/A INVX1_LOC
XINVX1_LOC_521 INVX1_LOC_521/Y VSS VDD INVX1_LOC_521/A INVX1_LOC
XINVX1_LOC_510 INVX1_LOC_510/Y VSS VDD INVX1_LOC_510/A INVX1_LOC
XINVX1_LOC_532 INVX1_LOC_532/Y VSS VDD INVX1_LOC_259/Y INVX1_LOC
XINVX1_LOC_576 INVX1_LOC_576/Y VSS VDD INVX1_LOC_576/A INVX1_LOC
XINVX1_LOC_565 INVX1_LOC_565/Y VSS VDD INVX1_LOC_565/A INVX1_LOC
XINVX1_LOC_587 INVX1_LOC_587/Y VSS VDD INVX1_LOC_587/A INVX1_LOC
XINVX1_LOC_598 INVX1_LOC_598/Y VSS VDD INVX1_LOC_598/A INVX1_LOC
XINVX1_LOC_543 INVX1_LOC_543/Y VSS VDD INVX1_LOC_543/A INVX1_LOC
XNAND2X1_LOC_709 NAND2X1_LOC_709/a_36_24# INVX1_LOC_551/A VSS VDD NAND2X1_LOC_698/Y
+ INVX1_LOC_552/Y NAND2X1_LOC
XINVX1_LOC_373 INVX1_LOC_373/Y VSS VDD INVX1_LOC_373/A INVX1_LOC
XINVX1_LOC_362 INVX1_LOC_362/Y VSS VDD INVX1_LOC_362/A INVX1_LOC
XINVX1_LOC_384 INVX1_LOC_384/Y VSS VDD INVX1_LOC_384/A INVX1_LOC
XINVX1_LOC_340 INVX1_LOC_340/Y VSS VDD INVX1_LOC_340/A INVX1_LOC
XINVX1_LOC_351 INVX1_LOC_351/Y VSS VDD INVX1_LOC_351/A INVX1_LOC
XINVX1_LOC_395 INVX1_LOC_395/Y VSS VDD INVX1_LOC_395/A INVX1_LOC
XINVX1_LOC_170 INVX1_LOC_170/Y VSS VDD INVX1_LOC_170/A INVX1_LOC
XNAND2X1_LOC_539 NAND2X1_LOC_539/a_36_24# INVX1_LOC_412/A VSS VDD INVX1_LOC_410/Y
+ INVX1_LOC_411/Y NAND2X1_LOC
XNAND2X1_LOC_517 NAND2X1_LOC_517/a_36_24# NAND2X1_LOC_517/Y VSS VDD INVX1_LOC_41/Y
+ INVX1_LOC_404/Y NAND2X1_LOC
XNAND2X1_LOC_528 NAND2X1_LOC_528/a_36_24# NAND2X1_LOC_528/Y VSS VDD INVX1_LOC_11/Y
+ INVX1_LOC_50/Y NAND2X1_LOC
XNAND2X1_LOC_506 NAND2X1_LOC_506/a_36_24# INVX1_LOC_396/A VSS VDD NAND2X1_LOC_242/A
+ NAND2X1_LOC_506/B NAND2X1_LOC
XINVX1_LOC_192 INVX1_LOC_192/Y VSS VDD INVX1_LOC_192/A INVX1_LOC
XINVX1_LOC_181 INVX1_LOC_181/Y VSS VDD INVX1_LOC_181/A INVX1_LOC
XNAND2X1_LOC_325 NAND2X1_LOC_325/a_36_24# INVX1_LOC_257/A VSS VDD NAND2X1_LOC_322/Y
+ NAND2X1_LOC_325/B NAND2X1_LOC
XNAND2X1_LOC_314 NAND2X1_LOC_314/a_36_24# NAND2X1_LOC_317/B VSS VDD INVX1_LOC_79/A
+ INVX1_LOC_69/Y NAND2X1_LOC
XNAND2X1_LOC_303 NAND2X1_LOC_303/a_36_24# INVX1_LOC_250/A VSS VDD INVX1_LOC_248/Y
+ INVX1_LOC_249/Y NAND2X1_LOC
XNAND2X1_LOC_336 NAND2X1_LOC_336/a_36_24# INVX1_LOC_270/A VSS VDD NAND2X1_LOC_538/B
+ NAND2X1_LOC_336/B NAND2X1_LOC
XNAND2X1_LOC_369 NAND2X1_LOC_369/a_36_24# NAND2X1_LOC_543/B VSS VDD INVX1_LOC_31/Y
+ INVX1_LOC_114/A NAND2X1_LOC
XNAND2X1_LOC_347 NAND2X1_LOC_347/a_36_24# INVX1_LOC_281/A VSS VDD NAND2X1_LOC_297/Y
+ INVX1_LOC_280/Y NAND2X1_LOC
XNAND2X1_LOC_358 NAND2X1_LOC_358/a_36_24# INVX1_LOC_292/A VSS VDD INVX1_LOC_284/Y
+ INVX1_LOC_285/Y NAND2X1_LOC
XNAND2X1_LOC_155 NAND2X1_LOC_155/a_36_24# INVX1_LOC_142/A VSS VDD INVX1_LOC_143/Y
+ INVX1_LOC_144/Y NAND2X1_LOC
XNAND2X1_LOC_144 NAND2X1_LOC_144/a_36_24# NAND2X1_LOC_147/B VSS VDD INVX1_LOC_63/Y
+ INVX1_LOC_395/A NAND2X1_LOC
XNAND2X1_LOC_111 NAND2X1_LOC_111/a_36_24# NAND2X1_LOC_111/Y VSS VDD INVX1_LOC_41/Y
+ INVX1_LOC_103/Y NAND2X1_LOC
XNAND2X1_LOC_122 NAND2X1_LOC_122/a_36_24# NAND2X1_LOC_122/Y VSS VDD INVX1_LOC_50/Y
+ NAND2X1_LOC_121/Y NAND2X1_LOC
XNAND2X1_LOC_177 NAND2X1_LOC_177/a_36_24# NAND2X1_LOC_180/B VSS VDD INVX1_LOC_54/Y
+ INVX1_LOC_74/Y NAND2X1_LOC
XNAND2X1_LOC_166 NAND2X1_LOC_166/a_36_24# NAND2X1_LOC_169/A VSS VDD INVX1_LOC_79/A
+ INVX1_LOC_48/Y NAND2X1_LOC
XNAND2X1_LOC_133 NAND2X1_LOC_133/a_36_24# INVX1_LOC_123/A VSS VDD INVX1_LOC_12/Y INVX1_LOC_84/A
+ NAND2X1_LOC
XNAND2X1_LOC_100 NAND2X1_LOC_100/a_36_24# INVX1_LOC_97/A VSS VDD NAND2X1_LOC_86/Y
+ NAND2X1_LOC_88/Y NAND2X1_LOC
XNAND2X1_LOC_188 NAND2X1_LOC_188/a_36_24# NAND2X1_LOC_498/B VSS VDD INVX1_LOC_165/Y
+ INVX1_LOC_588/A NAND2X1_LOC
XNAND2X1_LOC_199 NAND2X1_LOC_199/a_36_24# INVX1_LOC_175/A VSS VDD INVX1_LOC_171/Y
+ INVX1_LOC_172/Y NAND2X1_LOC
XINVX1_LOC_90 INVX1_LOC_90/Y VSS VDD INVX1_LOC_90/A INVX1_LOC
XINVX1_LOC_511 INVX1_LOC_511/Y VSS VDD INVX1_LOC_511/A INVX1_LOC
XINVX1_LOC_500 INVX1_LOC_500/Y VSS VDD INVX1_LOC_500/A INVX1_LOC
XINVX1_LOC_522 INVX1_LOC_522/Y VSS VDD INVX1_LOC_522/A INVX1_LOC
XINVX1_LOC_555 INVX1_LOC_555/Y VSS VDD INVX1_LOC_555/A INVX1_LOC
XINVX1_LOC_544 INVX1_LOC_544/Y VSS VDD INVX1_LOC_544/A INVX1_LOC
XINVX1_LOC_588 INVX1_LOC_588/Y VSS VDD INVX1_LOC_588/A INVX1_LOC
XINVX1_LOC_533 INVX1_LOC_533/Y VSS VDD INVX1_LOC_533/A INVX1_LOC
XINVX1_LOC_577 INVX1_LOC_577/Y VSS VDD INVX1_LOC_577/A INVX1_LOC
XINVX1_LOC_566 INVX1_LOC_566/Y VSS VDD INVX1_LOC_566/A INVX1_LOC
XINVX1_LOC_599 INVX1_LOC_599/Y VSS VDD INVX1_LOC_599/A INVX1_LOC
XINVX1_LOC_330 INVX1_LOC_335/A VSS VDD INVX1_LOC_330/A INVX1_LOC
XINVX1_LOC_352 INVX1_LOC_352/Y VSS VDD INVX1_LOC_352/A INVX1_LOC
XINVX1_LOC_341 INVX1_LOC_341/Y VSS VDD INPUT_5 INVX1_LOC
XINVX1_LOC_374 INVX1_LOC_374/Y VSS VDD INVX1_LOC_374/A INVX1_LOC
XINVX1_LOC_363 INVX1_LOC_363/Y VSS VDD INVX1_LOC_363/A INVX1_LOC
XINVX1_LOC_385 INVX1_LOC_385/Y VSS VDD INVX1_LOC_385/A INVX1_LOC
XINVX1_LOC_396 INVX1_LOC_396/Y VSS VDD INVX1_LOC_396/A INVX1_LOC
XNAND2X1_LOC_518 NAND2X1_LOC_518/a_36_24# NAND2X1_LOC_520/A VSS VDD INVX1_LOC_69/Y
+ INVX1_LOC_76/Y NAND2X1_LOC
XNAND2X1_LOC_507 NAND2X1_LOC_507/a_36_24# INVX1_LOC_397/A VSS VDD NAND2X1_LOC_507/A
+ NAND2X1_LOC_505/Y NAND2X1_LOC
XINVX1_LOC_193 INVX1_LOC_193/Y VSS VDD INVX1_LOC_193/A INVX1_LOC
XINVX1_LOC_160 INVX1_LOC_160/Y VSS VDD INVX1_LOC_160/A INVX1_LOC
XINVX1_LOC_171 INVX1_LOC_171/Y VSS VDD INVX1_LOC_171/A INVX1_LOC
XINVX1_LOC_182 INVX1_LOC_182/Y VSS VDD INVX1_LOC_182/A INVX1_LOC
XNAND2X1_LOC_529 NAND2X1_LOC_529/a_36_24# NAND2X1_LOC_529/Y VSS VDD INPUT_3 INVX1_LOC_35/Y
+ NAND2X1_LOC
XNAND2X1_LOC_326 NAND2X1_LOC_326/a_36_24# INVX1_LOC_258/A VSS VDD INVX1_LOC_256/Y
+ INVX1_LOC_257/Y NAND2X1_LOC
XNAND2X1_LOC_348 NAND2X1_LOC_348/a_36_24# INVX1_LOC_282/A VSS VDD INVX1_LOC_278/Y
+ INVX1_LOC_279/Y NAND2X1_LOC
XNAND2X1_LOC_359 NAND2X1_LOC_359/a_36_24# INVX1_LOC_293/A VSS VDD INVX1_LOC_282/Y
+ INVX1_LOC_283/Y NAND2X1_LOC
XNAND2X1_LOC_337 NAND2X1_LOC_337/a_36_24# INVX1_LOC_271/A VSS VDD INVX1_LOC_269/Y
+ INVX1_LOC_270/Y NAND2X1_LOC
XNAND2X1_LOC_315 NAND2X1_LOC_315/a_36_24# NAND2X1_LOC_318/A VSS VDD INVX1_LOC_41/Y
+ INVX1_LOC_479/A NAND2X1_LOC
XNAND2X1_LOC_304 NAND2X1_LOC_304/a_36_24# NAND2X1_LOC_307/A VSS VDD INVX1_LOC_59/Y
+ INVX1_LOC_206/Y NAND2X1_LOC
XNAND2X1_LOC_860 NAND2X1_LOC_860/a_36_24# INVX1_LOC_681/A VSS VDD INVX1_LOC_211/Y
+ INVX1_LOC_321/Y NAND2X1_LOC
XNAND2X1_LOC_123 NAND2X1_LOC_123/a_36_24# INVX1_LOC_115/A VSS VDD NAND2X1_LOC_123/A
+ NAND2X1_LOC_123/B NAND2X1_LOC
XNAND2X1_LOC_178 NAND2X1_LOC_178/a_36_24# NAND2X1_LOC_181/A VSS VDD INVX1_LOC_62/Y
+ INVX1_LOC_145/Y NAND2X1_LOC
XNAND2X1_LOC_189 NAND2X1_LOC_189/a_36_24# NAND2X1_LOC_192/A VSS VDD INVX1_LOC_93/Y
+ NAND2X1_LOC_498/B NAND2X1_LOC
XNAND2X1_LOC_134 NAND2X1_LOC_134/a_36_24# NAND2X1_LOC_768/B VSS VDD INVX1_LOC_93/Y
+ INVX1_LOC_479/A NAND2X1_LOC
XNAND2X1_LOC_156 NAND2X1_LOC_156/a_36_24# NAND2X1_LOC_156/Y VSS VDD INVX1_LOC_139/Y
+ INVX1_LOC_142/Y NAND2X1_LOC
XNAND2X1_LOC_145 NAND2X1_LOC_145/a_36_24# NAND2X1_LOC_148/A VSS VDD INVX1_LOC_58/Y
+ INVX1_LOC_80/A NAND2X1_LOC
XNAND2X1_LOC_112 NAND2X1_LOC_112/a_36_24# INVX1_LOC_105/A VSS VDD NAND2X1_LOC_775/B
+ NAND2X1_LOC_111/Y NAND2X1_LOC
XNAND2X1_LOC_167 NAND2X1_LOC_167/a_36_24# NAND2X1_LOC_388/A VSS VDD INVX1_LOC_69/Y
+ INVX1_LOC_586/A NAND2X1_LOC
XNAND2X1_LOC_101 NAND2X1_LOC_101/a_36_24# INVX1_LOC_98/A VSS VDD INVX1_LOC_96/Y INVX1_LOC_97/Y
+ NAND2X1_LOC
XNAND2X1_LOC_690 NAND2X1_LOC_690/a_36_24# NAND2X1_LOC_690/Y VSS VDD INVX1_LOC_541/Y
+ INVX1_LOC_338/Y NAND2X1_LOC
XINVX1_LOC_91 INVX1_LOC_91/Y VSS VDD INVX1_LOC_91/A INVX1_LOC
XINVX1_LOC_80 INVX1_LOC_80/Y VSS VDD INVX1_LOC_80/A INVX1_LOC
XINVX1_LOC_534 INVX1_LOC_534/Y VSS VDD INVX1_LOC_479/A INVX1_LOC
XINVX1_LOC_523 INVX1_LOC_523/Y VSS VDD INVX1_LOC_523/A INVX1_LOC
XINVX1_LOC_512 INVX1_LOC_512/Y VSS VDD INVX1_LOC_512/A INVX1_LOC
XINVX1_LOC_501 INVX1_LOC_501/Y VSS VDD INVX1_LOC_501/A INVX1_LOC
XINVX1_LOC_545 INVX1_LOC_545/Y VSS VDD INVX1_LOC_545/A INVX1_LOC
XINVX1_LOC_567 INVX1_LOC_567/Y VSS VDD INVX1_LOC_567/A INVX1_LOC
XINVX1_LOC_556 INVX1_LOC_556/Y VSS VDD INVX1_LOC_556/A INVX1_LOC
XINVX1_LOC_578 INVX1_LOC_578/Y VSS VDD INVX1_LOC_578/A INVX1_LOC
XINVX1_LOC_589 INVX1_LOC_589/Y VSS VDD INVX1_LOC_100/Y INVX1_LOC
XINVX1_LOC_331 INVX1_LOC_331/Y VSS VDD INVX1_LOC_62/Y INVX1_LOC
XINVX1_LOC_386 INVX1_LOC_386/Y VSS VDD INVX1_LOC_386/A INVX1_LOC
XINVX1_LOC_375 INVX1_LOC_375/Y VSS VDD INVX1_LOC_375/A INVX1_LOC
XINVX1_LOC_364 INVX1_LOC_364/Y VSS VDD INVX1_LOC_364/A INVX1_LOC
XINVX1_LOC_353 INVX1_LOC_353/Y VSS VDD INVX1_LOC_353/A INVX1_LOC
XINVX1_LOC_320 INVX1_LOC_320/Y VSS VDD INVX1_LOC_320/A INVX1_LOC
XINVX1_LOC_342 INVX1_LOC_342/Y VSS VDD INVX1_LOC_342/A INVX1_LOC
XINVX1_LOC_397 INVX1_LOC_397/Y VSS VDD INVX1_LOC_397/A INVX1_LOC
XINVX1_LOC_183 INVX1_LOC_183/Y VSS VDD INVX1_LOC_183/A INVX1_LOC
XNAND2X1_LOC_519 NAND2X1_LOC_519/a_36_24# NAND2X1_LOC_520/B VSS VDD INVX1_LOC_51/Y
+ INVX1_LOC_145/Y NAND2X1_LOC
XNAND2X1_LOC_508 NAND2X1_LOC_508/a_36_24# INVX1_LOC_398/A VSS VDD INVX1_LOC_396/Y
+ INVX1_LOC_397/Y NAND2X1_LOC
XINVX1_LOC_150 INVX1_LOC_150/Y VSS VDD INVX1_LOC_150/A INVX1_LOC
XINVX1_LOC_161 INVX1_LOC_588/A VSS VDD INVX1_LOC_161/A INVX1_LOC
XINVX1_LOC_194 INVX1_LOC_194/Y VSS VDD INVX1_LOC_194/A INVX1_LOC
XINVX1_LOC_172 INVX1_LOC_172/Y VSS VDD INVX1_LOC_172/A INVX1_LOC
XNAND2X1_LOC_305 NAND2X1_LOC_305/a_36_24# NAND2X1_LOC_307/B VSS VDD INVX1_LOC_6/Y
+ INVX1_LOC_89/Y NAND2X1_LOC
XNAND2X1_LOC_349 NAND2X1_LOC_349/a_36_24# INVX1_LOC_283/A VSS VDD INVX1_LOC_276/Y
+ INVX1_LOC_277/Y NAND2X1_LOC
XNAND2X1_LOC_327 NAND2X1_LOC_327/a_36_24# INVX1_LOC_259/A VSS VDD INVX1_LOC_260/Y
+ INVX1_LOC_224/Y NAND2X1_LOC
XNAND2X1_LOC_338 NAND2X1_LOC_338/a_36_24# INVX1_LOC_272/A VSS VDD INVX1_LOC_267/Y
+ INVX1_LOC_268/Y NAND2X1_LOC
XNAND2X1_LOC_316 NAND2X1_LOC_316/a_36_24# NAND2X1_LOC_318/B VSS VDD INVX1_LOC_20/Y
+ INVX1_LOC_81/Y NAND2X1_LOC
XNAND2X1_LOC_850 NAND2X1_LOC_850/a_36_24# INVX1_LOC_671/A VSS VDD INVX1_LOC_663/Y
+ INVX1_LOC_664/Y NAND2X1_LOC
XNAND2X1_LOC_861 NAND2X1_LOC_861/a_36_24# INVX1_LOC_682/A VSS VDD INVX1_LOC_486/Y
+ INVX1_LOC_681/Y NAND2X1_LOC
XNAND2X1_LOC_135 NAND2X1_LOC_135/a_36_24# NAND2X1_LOC_332/B VSS VDD INVX1_LOC_63/Y
+ INVX1_LOC_479/A NAND2X1_LOC
XNAND2X1_LOC_113 NAND2X1_LOC_113/a_36_24# INVX1_LOC_106/A VSS VDD NAND2X1_LOC_768/A
+ NAND2X1_LOC_107/Y NAND2X1_LOC
XNAND2X1_LOC_146 NAND2X1_LOC_146/a_36_24# NAND2X1_LOC_148/B VSS VDD INVX1_LOC_45/Y
+ INVX1_LOC_117/Y NAND2X1_LOC
XNAND2X1_LOC_179 NAND2X1_LOC_179/a_36_24# NAND2X1_LOC_179/Y VSS VDD INVX1_LOC_45/Y
+ INVX1_LOC_100/Y NAND2X1_LOC
XNAND2X1_LOC_124 NAND2X1_LOC_124/a_36_24# INVX1_LOC_116/A VSS VDD NAND2X1_LOC_122/Y
+ INVX1_LOC_115/Y NAND2X1_LOC
XNAND2X1_LOC_102 NAND2X1_LOC_102/a_36_24# INVX1_LOC_99/A VSS VDD INVX1_LOC_12/Y INVX1_LOC_92/A
+ NAND2X1_LOC
XNAND2X1_LOC_168 NAND2X1_LOC_168/a_36_24# INVX1_LOC_153/A VSS VDD NAND2X1_LOC_164/Y
+ NAND2X1_LOC_165/Y NAND2X1_LOC
XNAND2X1_LOC_157 NAND2X1_LOC_157/a_36_24# INVX1_LOC_145/A VSS VDD INVX1_LOC_3/Y INVX1_LOC_25/Y
+ NAND2X1_LOC
XNAND2X1_LOC_691 NAND2X1_LOC_691/a_36_24# INVX1_LOC_542/A VSS VDD NAND2X1_LOC_691/A
+ NAND2X1_LOC_690/Y NAND2X1_LOC
XNAND2X1_LOC_680 NAND2X1_LOC_680/a_36_24# NAND2X1_LOC_728/B VSS VDD INVX1_LOC_58/Y
+ NAND2X1_LOC_331/A NAND2X1_LOC
XINVX1_LOC_92 INVX1_LOC_92/Y VSS VDD INVX1_LOC_92/A INVX1_LOC
XINVX1_LOC_70 INVX1_LOC_70/Y VSS VDD INVX1_LOC_6/Y INVX1_LOC
XINVX1_LOC_81 INVX1_LOC_81/Y VSS VDD INVX1_LOC_81/A INVX1_LOC
XINVX1_LOC_535 INVX1_LOC_535/Y VSS VDD INVX1_LOC_20/Y INVX1_LOC
XINVX1_LOC_568 INVX1_LOC_568/Y VSS VDD INVX1_LOC_568/A INVX1_LOC
XINVX1_LOC_513 INVX1_LOC_513/Y VSS VDD INVX1_LOC_513/A INVX1_LOC
XINVX1_LOC_557 INVX1_LOC_557/Y VSS VDD INVX1_LOC_557/A INVX1_LOC
XINVX1_LOC_546 INVX1_LOC_546/Y VSS VDD INVX1_LOC_546/A INVX1_LOC
XINVX1_LOC_502 INVX1_LOC_502/Y VSS VDD INVX1_LOC_502/A INVX1_LOC
XINVX1_LOC_524 INVX1_LOC_524/Y VSS VDD INVX1_LOC_76/Y INVX1_LOC
XINVX1_LOC_579 INVX1_LOC_579/Y VSS VDD INVX1_LOC_579/A INVX1_LOC
XINVX1_LOC_332 INVX1_LOC_332/Y VSS VDD INVX1_LOC_137/Y INVX1_LOC
XINVX1_LOC_387 INVX1_LOC_387/Y VSS VDD INVX1_LOC_387/A INVX1_LOC
XINVX1_LOC_376 INVX1_LOC_376/Y VSS VDD INVX1_LOC_376/A INVX1_LOC
XINVX1_LOC_354 INVX1_LOC_354/Y VSS VDD INVX1_LOC_354/A INVX1_LOC
XINVX1_LOC_321 INVX1_LOC_321/Y VSS VDD INVX1_LOC_321/A INVX1_LOC
XINVX1_LOC_398 INVX1_LOC_398/Y VSS VDD INVX1_LOC_398/A INVX1_LOC
XINVX1_LOC_343 INVX1_LOC_343/Y VSS VDD INPUT_7 INVX1_LOC
XINVX1_LOC_310 INVX1_LOC_310/Y VSS VDD INVX1_LOC_20/Y INVX1_LOC
XINVX1_LOC_365 INVX1_LOC_365/Y VSS VDD INVX1_LOC_365/A INVX1_LOC
XNAND2X1_LOC_509 NAND2X1_LOC_509/a_36_24# INVX1_LOC_399/A VSS VDD INVX1_LOC_201/Y
+ NAND2X1_LOC_503/Y NAND2X1_LOC
XINVX1_LOC_162 INVX1_LOC_162/Y VSS VDD INVX1_LOC_62/Y INVX1_LOC
XINVX1_LOC_151 INVX1_LOC_151/Y VSS VDD INVX1_LOC_479/A INVX1_LOC
XINVX1_LOC_140 INVX1_LOC_140/Y VSS VDD INVX1_LOC_11/Y INVX1_LOC
XINVX1_LOC_173 INVX1_LOC_173/Y VSS VDD INVX1_LOC_173/A INVX1_LOC
XINVX1_LOC_195 INVX1_LOC_195/Y VSS VDD INVX1_LOC_195/A INVX1_LOC
XINVX1_LOC_184 INVX1_LOC_184/Y VSS VDD INVX1_LOC_184/A INVX1_LOC
XNAND2X1_LOC_317 NAND2X1_LOC_317/a_36_24# INVX1_LOC_253/A VSS VDD NAND2X1_LOC_317/A
+ NAND2X1_LOC_317/B NAND2X1_LOC
XNAND2X1_LOC_306 NAND2X1_LOC_306/a_36_24# NAND2X1_LOC_308/A VSS VDD INVX1_LOC_31/Y
+ INVX1_LOC_395/A NAND2X1_LOC
XNAND2X1_LOC_328 NAND2X1_LOC_328/a_36_24# INVX1_LOC_261/A VSS VDD INVX1_LOC_262/Y
+ INVX1_LOC_55/Y NAND2X1_LOC
XNAND2X1_LOC_339 NAND2X1_LOC_339/a_36_24# INVX1_LOC_273/A VSS VDD INVX1_LOC_64/Y INVX1_LOC_266/Y
+ NAND2X1_LOC
XNAND2X1_LOC_840 NAND2X1_LOC_840/a_36_24# INVX1_LOC_661/A VSS VDD INVX1_LOC_654/Y
+ INVX1_LOC_655/Y NAND2X1_LOC
XNAND2X1_LOC_862 NAND2X1_LOC_862/a_36_24# INVX1_LOC_683/A VSS VDD INVX1_LOC_679/Y
+ INVX1_LOC_680/Y NAND2X1_LOC
XNAND2X1_LOC_851 NAND2X1_LOC_851/a_36_24# INVX1_LOC_672/A VSS VDD INVX1_LOC_661/Y
+ INVX1_LOC_662/Y NAND2X1_LOC
XNAND2X1_LOC_125 NAND2X1_LOC_125/a_36_24# NAND2X1_LOC_128/A VSS VDD INVX1_LOC_93/Y
+ INVX1_LOC_100/Y NAND2X1_LOC
XNAND2X1_LOC_103 NAND2X1_LOC_103/a_36_24# NAND2X1_LOC_768/A VSS VDD INVX1_LOC_53/Y
+ INVX1_LOC_99/Y NAND2X1_LOC
XNAND2X1_LOC_114 NAND2X1_LOC_114/a_36_24# INVX1_LOC_107/A VSS VDD NAND2X1_LOC_108/Y
+ INVX1_LOC_106/Y NAND2X1_LOC
XNAND2X1_LOC_136 NAND2X1_LOC_136/a_36_24# NAND2X1_LOC_136/Y VSS VDD INVX1_LOC_6/Y
+ INVX1_LOC_49/Y NAND2X1_LOC
XNAND2X1_LOC_147 NAND2X1_LOC_147/a_36_24# INVX1_LOC_131/A VSS VDD NAND2X1_LOC_142/Y
+ NAND2X1_LOC_147/B NAND2X1_LOC
XNAND2X1_LOC_158 NAND2X1_LOC_158/a_36_24# NAND2X1_LOC_210/A VSS VDD NAND2X1_LOC_156/Y
+ INVX1_LOC_145/Y NAND2X1_LOC
XNAND2X1_LOC_169 NAND2X1_LOC_169/a_36_24# INVX1_LOC_154/A VSS VDD NAND2X1_LOC_169/A
+ NAND2X1_LOC_388/A NAND2X1_LOC
XNAND2X1_LOC_1 NAND2X1_LOC_1/a_36_24# INVX1_LOC_1/A VSS VDD INVX1_LOC_2/Y INPUT_7
+ NAND2X1_LOC
XNAND2X1_LOC_681 NAND2X1_LOC_681/a_36_24# NAND2X1_LOC_685/A VSS VDD INVX1_LOC_41/Y
+ INVX1_LOC_137/Y NAND2X1_LOC
XNAND2X1_LOC_670 NAND2X1_LOC_670/a_36_24# NAND2X1_LOC_673/A VSS VDD INVX1_LOC_48/Y
+ INVX1_LOC_99/Y NAND2X1_LOC
XINVX1_LOC_60 INVX1_LOC_60/Y VSS VDD INPUT_5 INVX1_LOC
XINVX1_LOC_82 INVX1_LOC_82/Y VSS VDD INVX1_LOC_84/A INVX1_LOC
XNAND2X1_LOC_692 NAND2X1_LOC_692/a_36_24# NAND2X1_LOC_692/Y VSS VDD INVX1_LOC_26/Y
+ INVX1_LOC_51/Y NAND2X1_LOC
XINVX1_LOC_71 INVX1_LOC_71/Y VSS VDD INVX1_LOC_35/Y INVX1_LOC
XINVX1_LOC_93 INVX1_LOC_93/Y VSS VDD INVX1_LOC_93/A INVX1_LOC
XINVX1_LOC_514 INVX1_LOC_514/Y VSS VDD INVX1_LOC_514/A INVX1_LOC
XINVX1_LOC_569 INVX1_LOC_569/Y VSS VDD INVX1_LOC_569/A INVX1_LOC
XINVX1_LOC_547 INVX1_LOC_547/Y VSS VDD INVX1_LOC_547/A INVX1_LOC
XINVX1_LOC_536 INVX1_LOC_536/Y VSS VDD INVX1_LOC_536/A INVX1_LOC
XINVX1_LOC_558 INVX1_LOC_558/Y VSS VDD INVX1_LOC_558/A INVX1_LOC
XINVX1_LOC_503 INVX1_LOC_503/Y VSS VDD INVX1_LOC_503/A INVX1_LOC
XINVX1_LOC_525 INVX1_LOC_525/Y VSS VDD INVX1_LOC_80/A INVX1_LOC
XINVX1_LOC_300 INVX1_LOC_300/Y VSS VDD INVX1_LOC_300/A INVX1_LOC
XINVX1_LOC_355 INVX1_LOC_355/Y VSS VDD INVX1_LOC_355/A INVX1_LOC
XINVX1_LOC_377 INVX1_LOC_377/Y VSS VDD INVX1_LOC_377/A INVX1_LOC
XINVX1_LOC_344 INVX1_LOC_344/Y VSS VDD INVX1_LOC_344/A INVX1_LOC
XINVX1_LOC_388 INVX1_LOC_388/Y VSS VDD INVX1_LOC_388/A INVX1_LOC
XINVX1_LOC_333 INVX1_LOC_333/Y VSS VDD INVX1_LOC_333/A INVX1_LOC
XINVX1_LOC_399 INVX1_LOC_399/Y VSS VDD INVX1_LOC_399/A INVX1_LOC
XINVX1_LOC_322 INVX1_LOC_322/Y VSS VDD INVX1_LOC_79/A INVX1_LOC
XINVX1_LOC_311 INVX1_LOC_311/Y VSS VDD INVX1_LOC_35/Y INVX1_LOC
XINVX1_LOC_366 INVX1_LOC_366/Y VSS VDD INVX1_LOC_366/A INVX1_LOC
XINVX1_LOC_152 INVX1_LOC_152/Y VSS VDD INVX1_LOC_586/A INVX1_LOC
XINVX1_LOC_141 INVX1_LOC_141/Y VSS VDD INVX1_LOC_47/Y INVX1_LOC
XINVX1_LOC_130 INVX1_LOC_130/Y VSS VDD INPUT_1 INVX1_LOC
XINVX1_LOC_185 INVX1_LOC_185/Y VSS VDD INVX1_LOC_185/A INVX1_LOC
XINVX1_LOC_163 INVX1_LOC_163/Y VSS VDD INVX1_LOC_76/Y INVX1_LOC
XINVX1_LOC_196 INVX1_LOC_196/Y VSS VDD INVX1_LOC_196/A INVX1_LOC
XINVX1_LOC_174 INVX1_LOC_174/Y VSS VDD INVX1_LOC_174/A INVX1_LOC
XNAND2X1_LOC_307 NAND2X1_LOC_307/a_36_24# INVX1_LOC_251/A VSS VDD NAND2X1_LOC_307/A
+ NAND2X1_LOC_307/B NAND2X1_LOC
XNAND2X1_LOC_318 NAND2X1_LOC_318/a_36_24# INVX1_LOC_254/A VSS VDD NAND2X1_LOC_318/A
+ NAND2X1_LOC_318/B NAND2X1_LOC
XNAND2X1_LOC_329 NAND2X1_LOC_329/a_36_24# NAND2X1_LOC_355/A VSS VDD INVX1_LOC_263/Y
+ INVX1_LOC_261/Y NAND2X1_LOC
XNAND2X1_LOC_841 NAND2X1_LOC_841/a_36_24# INVX1_LOC_662/A VSS VDD INVX1_LOC_652/Y
+ INVX1_LOC_653/Y NAND2X1_LOC
XNAND2X1_LOC_830 NAND2X1_LOC_830/a_36_24# INVX1_LOC_651/A VSS VDD NAND2X1_LOC_108/Y
+ NAND2X1_LOC_142/Y NAND2X1_LOC
XNAND2X1_LOC_863 NAND2X1_LOC_863/a_36_24# INVX1_LOC_684/A VSS VDD INVX1_LOC_677/Y
+ INVX1_LOC_678/Y NAND2X1_LOC
XNAND2X1_LOC_852 NAND2X1_LOC_852/a_36_24# INVX1_LOC_673/A VSS VDD INVX1_LOC_659/Y
+ INVX1_LOC_660/Y NAND2X1_LOC
XNAND2X1_LOC_115 NAND2X1_LOC_115/a_36_24# INVX1_LOC_108/A VSS VDD NAND2X1_LOC_106/Y
+ INVX1_LOC_105/Y NAND2X1_LOC
XNAND2X1_LOC_137 NAND2X1_LOC_137/a_36_24# INVX1_LOC_124/A VSS VDD NAND2X1_LOC_137/A
+ NAND2X1_LOC_768/B NAND2X1_LOC
XNAND2X1_LOC_159 NAND2X1_LOC_159/a_36_24# INVX1_LOC_146/A VSS VDD INVX1_LOC_9/Y INVX1_LOC_66/A
+ NAND2X1_LOC
XNAND2X1_LOC_148 NAND2X1_LOC_148/a_36_24# INVX1_LOC_132/A VSS VDD NAND2X1_LOC_148/A
+ NAND2X1_LOC_148/B NAND2X1_LOC
XNAND2X1_LOC_104 NAND2X1_LOC_104/a_36_24# INVX1_LOC_100/A VSS VDD INVX1_LOC_7/Y INVX1_LOC_12/Y
+ NAND2X1_LOC
XNAND2X1_LOC_126 NAND2X1_LOC_126/a_36_24# INVX1_LOC_117/A VSS VDD INVX1_LOC_7/Y INVX1_LOC_46/Y
+ NAND2X1_LOC
XNAND2X1_LOC_2 NAND2X1_LOC_2/a_36_24# INVX1_LOC_3/A VSS VDD INVX1_LOC_4/Y INVX1_LOC_5/Y
+ NAND2X1_LOC
XINVX1_LOC_83 INVX1_LOC_83/Y VSS VDD INVX1_LOC_83/A INVX1_LOC
XNAND2X1_LOC_693 NAND2X1_LOC_693/a_36_24# NAND2X1_LOC_706/B VSS VDD INVX1_LOC_21/Y
+ INVX1_LOC_45/Y NAND2X1_LOC
XNAND2X1_LOC_660 NAND2X1_LOC_660/a_36_24# INVX1_LOC_521/A VSS VDD INVX1_LOC_516/Y
+ INVX1_LOC_517/Y NAND2X1_LOC
XNAND2X1_LOC_682 NAND2X1_LOC_682/a_36_24# NAND2X1_LOC_685/B VSS VDD INVX1_LOC_45/Y
+ INVX1_LOC_586/A NAND2X1_LOC
XNAND2X1_LOC_671 NAND2X1_LOC_671/a_36_24# INVX1_LOC_530/A VSS VDD INPUT_2 INVX1_LOC_7/Y
+ NAND2X1_LOC
XINVX1_LOC_61 INVX1_LOC_92/A VSS VDD INVX1_LOC_61/A INVX1_LOC
XINVX1_LOC_94 INVX1_LOC_94/Y VSS VDD INVX1_LOC_94/A INVX1_LOC
XINVX1_LOC_50 INVX1_LOC_50/Y VSS VDD INVX1_LOC_50/A INVX1_LOC
XINVX1_LOC_72 INVX1_LOC_72/Y VSS VDD INVX1_LOC_9/Y INVX1_LOC
XINVX1_LOC_515 INVX1_LOC_515/Y VSS VDD INVX1_LOC_515/A INVX1_LOC
XINVX1_LOC_548 INVX1_LOC_548/Y VSS VDD INVX1_LOC_548/A INVX1_LOC
XINVX1_LOC_537 INVX1_LOC_537/Y VSS VDD INVX1_LOC_537/A INVX1_LOC
XINVX1_LOC_504 INVX1_LOC_504/Y VSS VDD INVX1_LOC_504/A INVX1_LOC
XINVX1_LOC_526 INVX1_LOC_526/Y VSS VDD INVX1_LOC_526/A INVX1_LOC
XINVX1_LOC_559 INVX1_LOC_559/Y VSS VDD INVX1_LOC_559/A INVX1_LOC
XNAND2X1_LOC_490 NAND2X1_LOC_490/a_36_24# NAND2X1_LOC_557/B VSS VDD INVX1_LOC_389/Y
+ INVX1_LOC_86/Y NAND2X1_LOC
XINVX1_LOC_301 INVX1_LOC_301/Y VSS VDD INVX1_LOC_301/A INVX1_LOC
XINVX1_LOC_312 INVX1_LOC_312/Y VSS VDD INVX1_LOC_312/A INVX1_LOC
XINVX1_LOC_323 INVX1_LOC_323/Y VSS VDD INVX1_LOC_245/A INVX1_LOC
XINVX1_LOC_334 INVX1_LOC_334/Y VSS VDD INPUT_6 INVX1_LOC
XINVX1_LOC_367 INVX1_LOC_367/Y VSS VDD INVX1_LOC_367/A INVX1_LOC
XINVX1_LOC_356 INVX1_LOC_356/Y VSS VDD INVX1_LOC_356/A INVX1_LOC
XINVX1_LOC_345 INVX1_LOC_345/Y VSS VDD INVX1_LOC_345/A INVX1_LOC
XINVX1_LOC_378 INVX1_LOC_378/Y VSS VDD INVX1_LOC_378/A INVX1_LOC
XINVX1_LOC_389 INVX1_LOC_389/Y VSS VDD INVX1_LOC_7/Y INVX1_LOC
XINVX1_LOC_131 INVX1_LOC_131/Y VSS VDD INVX1_LOC_131/A INVX1_LOC
XINVX1_LOC_142 INVX1_LOC_142/Y VSS VDD INVX1_LOC_142/A INVX1_LOC
XINVX1_LOC_186 INVX1_LOC_186/Y VSS VDD INVX1_LOC_186/A INVX1_LOC
XINVX1_LOC_164 INVX1_LOC_164/Y VSS VDD INVX1_LOC_134/Y INVX1_LOC
XINVX1_LOC_120 INVX1_LOC_120/Y VSS VDD INVX1_LOC_84/A INVX1_LOC
XINVX1_LOC_153 INVX1_LOC_153/Y VSS VDD INVX1_LOC_153/A INVX1_LOC
XINVX1_LOC_175 INVX1_LOC_175/Y VSS VDD INVX1_LOC_175/A INVX1_LOC
XINVX1_LOC_197 INVX1_LOC_197/Y VSS VDD INVX1_LOC_197/A INVX1_LOC
XNAND2X1_LOC_308 NAND2X1_LOC_308/a_36_24# INVX1_LOC_252/A VSS VDD NAND2X1_LOC_308/A
+ INVX1_LOC_251/Y NAND2X1_LOC
XNAND2X1_LOC_319 NAND2X1_LOC_319/a_36_24# INVX1_LOC_255/A VSS VDD INVX1_LOC_253/Y
+ INVX1_LOC_254/Y NAND2X1_LOC
XNAND2X1_LOC_831 NAND2X1_LOC_831/a_36_24# INVX1_LOC_652/A VSS VDD NAND2X1_LOC_274/B
+ NAND2X1_LOC_301/B NAND2X1_LOC
XNAND2X1_LOC_842 NAND2X1_LOC_842/a_36_24# INVX1_LOC_663/A VSS VDD NAND2X1_LOC_184/Y
+ INVX1_LOC_651/Y NAND2X1_LOC
XNAND2X1_LOC_820 NAND2X1_LOC_820/a_36_24# NAND2X1_LOC_820/Y VSS VDD NAND2X1_LOC_820/A
+ INVX1_LOC_649/Y NAND2X1_LOC
XNAND2X1_LOC_864 NAND2X1_LOC_864/a_36_24# INVX1_LOC_685/A VSS VDD INVX1_LOC_602/Y
+ INVX1_LOC_684/Y NAND2X1_LOC
XNAND2X1_LOC_853 NAND2X1_LOC_853/a_36_24# INVX1_LOC_674/A VSS VDD INVX1_LOC_44/Y INVX1_LOC_157/Y
+ NAND2X1_LOC
XNAND2X1_LOC_127 NAND2X1_LOC_127/a_36_24# NAND2X1_LOC_128/B VSS VDD INVX1_LOC_6/Y
+ INVX1_LOC_117/Y NAND2X1_LOC
XNAND2X1_LOC_116 NAND2X1_LOC_116/a_36_24# INVX1_LOC_109/A VSS VDD INVX1_LOC_107/Y
+ INVX1_LOC_108/Y NAND2X1_LOC
XNAND2X1_LOC_138 NAND2X1_LOC_138/a_36_24# INVX1_LOC_125/A VSS VDD NAND2X1_LOC_332/B
+ NAND2X1_LOC_136/Y NAND2X1_LOC
XNAND2X1_LOC_149 NAND2X1_LOC_149/a_36_24# INVX1_LOC_133/A VSS VDD INVX1_LOC_131/Y
+ INVX1_LOC_132/Y NAND2X1_LOC
XNAND2X1_LOC_105 NAND2X1_LOC_105/a_36_24# NAND2X1_LOC_106/B VSS VDD INVX1_LOC_101/Y
+ INVX1_LOC_102/Y NAND2X1_LOC
XNAND2X1_LOC_3 NAND2X1_LOC_3/a_36_24# INVX1_LOC_6/A VSS VDD INVX1_LOC_1/Y INVX1_LOC_3/Y
+ NAND2X1_LOC
XINVX1_LOC_84 INVX1_LOC_84/Y VSS VDD INVX1_LOC_84/A INVX1_LOC
XNAND2X1_LOC_683 NAND2X1_LOC_683/a_36_24# NAND2X1_LOC_686/A VSS VDD INVX1_LOC_79/A
+ INVX1_LOC_31/Y NAND2X1_LOC
XNAND2X1_LOC_694 NAND2X1_LOC_694/a_36_24# NAND2X1_LOC_707/A VSS VDD INVX1_LOC_479/A
+ INVX1_LOC_340/Y NAND2X1_LOC
XNAND2X1_LOC_650 NAND2X1_LOC_650/a_36_24# INVX1_LOC_511/A VSS VDD INVX1_LOC_500/Y
+ INVX1_LOC_501/Y NAND2X1_LOC
XNAND2X1_LOC_661 NAND2X1_LOC_661/a_36_24# INVX1_LOC_522/A VSS VDD INVX1_LOC_514/Y
+ INVX1_LOC_515/Y NAND2X1_LOC
XNAND2X1_LOC_672 NAND2X1_LOC_672/a_36_24# NAND2X1_LOC_673/B VSS VDD INVX1_LOC_145/Y
+ INVX1_LOC_530/Y NAND2X1_LOC
XINVX1_LOC_62 INVX1_LOC_62/Y VSS VDD INVX1_LOC_62/A INVX1_LOC
XINVX1_LOC_51 INVX1_LOC_51/Y VSS VDD INVX1_LOC_51/A INVX1_LOC
XINVX1_LOC_95 INVX1_LOC_95/Y VSS VDD INVX1_LOC_95/A INVX1_LOC
XINVX1_LOC_40 INVX1_LOC_40/Y VSS VDD INVX1_LOC_40/A INVX1_LOC
XINVX1_LOC_73 INVX1_LOC_73/Y VSS VDD INVX1_LOC_54/Y INVX1_LOC
XINVX1_LOC_516 INVX1_LOC_516/Y VSS VDD INVX1_LOC_516/A INVX1_LOC
XINVX1_LOC_505 INVX1_LOC_505/Y VSS VDD INVX1_LOC_505/A INVX1_LOC
XINVX1_LOC_527 INVX1_LOC_527/Y VSS VDD INVX1_LOC_224/Y INVX1_LOC
XINVX1_LOC_549 INVX1_LOC_549/Y VSS VDD INVX1_LOC_549/A INVX1_LOC
XINVX1_LOC_538 INVX1_LOC_538/Y VSS VDD INVX1_LOC_538/A INVX1_LOC
XNAND2X1_LOC_480 NAND2X1_LOC_480/a_36_24# GATE_479 VSS VDD INVX1_LOC_384/Y INVX1_LOC_385/Y
+ NAND2X1_LOC
XNAND2X1_LOC_491 NAND2X1_LOC_491/a_36_24# NAND2X1_LOC_491/Y VSS VDD INVX1_LOC_41/Y
+ INVX1_LOC_99/Y NAND2X1_LOC
XINVX1_LOC_335 INVX1_LOC_335/Y VSS VDD INVX1_LOC_335/A INVX1_LOC
XINVX1_LOC_357 INVX1_LOC_357/Y VSS VDD INVX1_LOC_357/A INVX1_LOC
XINVX1_LOC_302 INVX1_LOC_608/A VSS VDD INVX1_LOC_302/A INVX1_LOC
XINVX1_LOC_346 INVX1_LOC_346/Y VSS VDD INVX1_LOC_346/A INVX1_LOC
XINVX1_LOC_368 INVX1_LOC_368/Y VSS VDD INVX1_LOC_368/A INVX1_LOC
XINVX1_LOC_313 INVX1_LOC_313/Y VSS VDD INVX1_LOC_89/Y INVX1_LOC
XINVX1_LOC_324 INVX1_LOC_324/Y VSS VDD INVX1_LOC_324/A INVX1_LOC
XINVX1_LOC_379 INVX1_LOC_379/Y VSS VDD INVX1_LOC_379/A INVX1_LOC
XINVX1_LOC_143 INVX1_LOC_143/Y VSS VDD INVX1_LOC_54/Y INVX1_LOC
XINVX1_LOC_132 INVX1_LOC_132/Y VSS VDD INVX1_LOC_132/A INVX1_LOC
XINVX1_LOC_165 INVX1_LOC_165/Y VSS VDD INVX1_LOC_47/Y INVX1_LOC
XINVX1_LOC_110 INVX1_LOC_114/A VSS VDD INVX1_LOC_110/A INVX1_LOC
XINVX1_LOC_121 INVX1_LOC_121/Y VSS VDD INVX1_LOC_11/Y INVX1_LOC
XINVX1_LOC_187 INVX1_LOC_187/Y VSS VDD INVX1_LOC_187/A INVX1_LOC
XINVX1_LOC_154 INVX1_LOC_154/Y VSS VDD INVX1_LOC_154/A INVX1_LOC
XINVX1_LOC_176 INVX1_LOC_176/Y VSS VDD INVX1_LOC_176/A INVX1_LOC
XINVX1_LOC_198 INVX1_LOC_198/Y VSS VDD INVX1_LOC_198/A INVX1_LOC
XNAND2X1_LOC_309 NAND2X1_LOC_309/a_36_24# NAND2X1_LOC_370/A VSS VDD INVX1_LOC_31/Y
+ INVX1_LOC_199/Y NAND2X1_LOC
XNAND2X1_LOC_854 NAND2X1_LOC_854/a_36_24# INVX1_LOC_675/A VSS VDD INVX1_LOC_258/Y
+ INVX1_LOC_409/Y NAND2X1_LOC
XNAND2X1_LOC_832 NAND2X1_LOC_832/a_36_24# INVX1_LOC_653/A VSS VDD NAND2X1_LOC_832/A
+ NAND2X1_LOC_433/Y NAND2X1_LOC
XNAND2X1_LOC_843 NAND2X1_LOC_843/a_36_24# INVX1_LOC_664/A VSS VDD NAND2X1_LOC_843/A
+ NAND2X1_LOC_843/B NAND2X1_LOC
XNAND2X1_LOC_865 NAND2X1_LOC_865/a_36_24# INVX1_LOC_686/A VSS VDD INVX1_LOC_682/Y
+ INVX1_LOC_683/Y NAND2X1_LOC
XNAND2X1_LOC_810 NAND2X1_LOC_810/a_36_24# INVX1_LOC_640/A VSS VDD INVX1_LOC_602/Y
+ INVX1_LOC_639/Y NAND2X1_LOC
XNAND2X1_LOC_821 NAND2X1_LOC_821/a_36_24# NAND2X1_LOC_835/A VSS VDD INVX1_LOC_17/Y
+ INVX1_LOC_74/Y NAND2X1_LOC
XNAND2X1_LOC_106 NAND2X1_LOC_106/a_36_24# NAND2X1_LOC_106/Y VSS VDD INVX1_LOC_53/Y
+ NAND2X1_LOC_106/B NAND2X1_LOC
XNAND2X1_LOC_128 NAND2X1_LOC_128/a_36_24# INVX1_LOC_118/A VSS VDD NAND2X1_LOC_128/A
+ NAND2X1_LOC_128/B NAND2X1_LOC
XNAND2X1_LOC_139 NAND2X1_LOC_139/a_36_24# INVX1_LOC_126/A VSS VDD INVX1_LOC_124/Y
+ INVX1_LOC_125/Y NAND2X1_LOC
XNAND2X1_LOC_117 NAND2X1_LOC_117/a_36_24# NAND2X1_LOC_123/A VSS VDD INVX1_LOC_68/Y
+ INVX1_LOC_74/Y NAND2X1_LOC
XNAND2X1_LOC_4 NAND2X1_LOC_4/a_36_24# INVX1_LOC_7/A VSS VDD INPUT_0 INVX1_LOC_8/Y
+ NAND2X1_LOC
XNAND2X1_LOC_695 NAND2X1_LOC_695/a_36_24# NAND2X1_LOC_707/B VSS VDD INVX1_LOC_32/Y
+ INVX1_LOC_53/Y NAND2X1_LOC
XNAND2X1_LOC_684 NAND2X1_LOC_684/a_36_24# NAND2X1_LOC_686/B VSS VDD INVX1_LOC_20/Y
+ INVX1_LOC_49/Y NAND2X1_LOC
XNAND2X1_LOC_640 NAND2X1_LOC_640/a_36_24# INVX1_LOC_500/A VSS VDD INVX1_LOC_491/Y
+ INVX1_LOC_493/Y NAND2X1_LOC
XNAND2X1_LOC_651 NAND2X1_LOC_651/a_36_24# INVX1_LOC_512/A VSS VDD INVX1_LOC_498/Y
+ INVX1_LOC_499/Y NAND2X1_LOC
XNAND2X1_LOC_662 NAND2X1_LOC_662/a_36_24# INVX1_LOC_523/A VSS VDD INVX1_LOC_521/Y
+ INVX1_LOC_522/Y NAND2X1_LOC
XNAND2X1_LOC_673 NAND2X1_LOC_673/a_36_24# INVX1_LOC_531/A VSS VDD NAND2X1_LOC_673/A
+ NAND2X1_LOC_673/B NAND2X1_LOC
XINVX1_LOC_52 INVX1_LOC_52/Y VSS VDD INPUT_1 INVX1_LOC
XINVX1_LOC_96 INVX1_LOC_96/Y VSS VDD INVX1_LOC_96/A INVX1_LOC
XINVX1_LOC_30 INVX1_LOC_30/Y VSS VDD INPUT_5 INVX1_LOC
XINVX1_LOC_74 INVX1_LOC_74/Y VSS VDD INVX1_LOC_74/A INVX1_LOC
XINVX1_LOC_41 INVX1_LOC_41/Y VSS VDD INVX1_LOC_41/A INVX1_LOC
XINVX1_LOC_63 INVX1_LOC_63/Y VSS VDD INVX1_LOC_63/A INVX1_LOC
XINVX1_LOC_85 INVX1_LOC_85/Y VSS VDD INVX1_LOC_85/A INVX1_LOC
XINVX1_LOC_517 INVX1_LOC_517/Y VSS VDD INVX1_LOC_517/A INVX1_LOC
XINVX1_LOC_539 INVX1_LOC_539/Y VSS VDD INVX1_LOC_47/Y INVX1_LOC
XINVX1_LOC_506 INVX1_LOC_506/Y VSS VDD INVX1_LOC_506/A INVX1_LOC
XINVX1_LOC_528 INVX1_LOC_528/Y VSS VDD INVX1_LOC_35/Y INVX1_LOC
XNAND2X1_LOC_481 NAND2X1_LOC_481/a_36_24# NAND2X1_LOC_555/B VSS VDD INVX1_LOC_6/Y
+ NAND2X1_LOC_294/Y NAND2X1_LOC
XNAND2X1_LOC_470 NAND2X1_LOC_470/a_36_24# INVX1_LOC_376/A VSS VDD INVX1_LOC_372/Y
+ INVX1_LOC_373/Y NAND2X1_LOC
XNAND2X1_LOC_492 NAND2X1_LOC_492/a_36_24# NAND2X1_LOC_493/B VSS VDD INVX1_LOC_63/Y
+ INVX1_LOC_117/Y NAND2X1_LOC
XINVX1_LOC_336 INVX1_LOC_336/Y VSS VDD INVX1_LOC_20/Y INVX1_LOC
XINVX1_LOC_358 INVX1_LOC_358/Y VSS VDD INVX1_LOC_358/A INVX1_LOC
XINVX1_LOC_303 INVX1_LOC_303/Y VSS VDD INPUT_1 INVX1_LOC
XINVX1_LOC_347 INVX1_LOC_347/Y VSS VDD INVX1_LOC_347/A INVX1_LOC
XINVX1_LOC_314 INVX1_LOC_314/Y VSS VDD INVX1_LOC_206/Y INVX1_LOC
XINVX1_LOC_369 INVX1_LOC_369/Y VSS VDD INVX1_LOC_369/A INVX1_LOC
XINVX1_LOC_325 INVX1_LOC_325/Y VSS VDD INVX1_LOC_325/A INVX1_LOC
XINVX1_LOC_100 INVX1_LOC_100/Y VSS VDD INVX1_LOC_100/A INVX1_LOC
XINVX1_LOC_144 INVX1_LOC_144/Y VSS VDD INVX1_LOC_137/Y INVX1_LOC
XINVX1_LOC_133 INVX1_LOC_133/Y VSS VDD INVX1_LOC_133/A INVX1_LOC
XINVX1_LOC_199 INVX1_LOC_199/Y VSS VDD INVX1_LOC_199/A INVX1_LOC
XINVX1_LOC_166 INVX1_LOC_166/Y VSS VDD INVX1_LOC_166/A INVX1_LOC
XINVX1_LOC_122 INVX1_LOC_122/Y VSS VDD INVX1_LOC_119/Y INVX1_LOC
XINVX1_LOC_111 INVX1_LOC_526/A VSS VDD INVX1_LOC_111/A INVX1_LOC
XINVX1_LOC_188 INVX1_LOC_188/Y VSS VDD INVX1_LOC_188/A INVX1_LOC
XINVX1_LOC_155 INVX1_LOC_155/Y VSS VDD INVX1_LOC_155/A INVX1_LOC
XINVX1_LOC_177 INVX1_LOC_177/Y VSS VDD INVX1_LOC_177/A INVX1_LOC
XNAND2X1_LOC_800 NAND2X1_LOC_800/a_36_24# INVX1_LOC_630/A VSS VDD INVX1_LOC_538/Y
+ NAND2X1_LOC_800/B NAND2X1_LOC
XNAND2X1_LOC_811 NAND2X1_LOC_811/a_36_24# INVX1_LOC_641/A VSS VDD INVX1_LOC_637/Y
+ INVX1_LOC_638/Y NAND2X1_LOC
XNAND2X1_LOC_822 NAND2X1_LOC_822/a_36_24# NAND2X1_LOC_822/Y VSS VDD INVX1_LOC_69/Y
+ INVX1_LOC_99/Y NAND2X1_LOC
XNAND2X1_LOC_844 NAND2X1_LOC_844/a_36_24# INVX1_LOC_665/A VSS VDD NAND2X1_LOC_844/A
+ INVX1_LOC_406/Y NAND2X1_LOC
XNAND2X1_LOC_833 NAND2X1_LOC_833/a_36_24# INVX1_LOC_654/A VSS VDD NAND2X1_LOC_482/Y
+ NAND2X1_LOC_833/B NAND2X1_LOC
XNAND2X1_LOC_855 NAND2X1_LOC_855/a_36_24# INVX1_LOC_676/A VSS VDD INVX1_LOC_542/Y
+ NAND2X1_LOC_829/Y NAND2X1_LOC
XNAND2X1_LOC_866 NAND2X1_LOC_866/a_36_24# GATE_865 VSS VDD INVX1_LOC_685/Y INVX1_LOC_686/Y
+ NAND2X1_LOC
XNAND2X1_LOC_107 NAND2X1_LOC_107/a_36_24# NAND2X1_LOC_107/Y VSS VDD INVX1_LOC_69/Y
+ INVX1_LOC_80/A NAND2X1_LOC
XNAND2X1_LOC_118 NAND2X1_LOC_118/a_36_24# NAND2X1_LOC_123/B VSS VDD INVX1_LOC_74/Y
+ INVX1_LOC_80/A NAND2X1_LOC
XNAND2X1_LOC_129 NAND2X1_LOC_129/a_36_24# INVX1_LOC_119/A VSS VDD INVX1_LOC_120/Y
+ INVX1_LOC_46/Y NAND2X1_LOC
XNAND2X1_LOC_5 NAND2X1_LOC_5/a_36_24# INVX1_LOC_9/A VSS VDD INVX1_LOC_10/Y INPUT_3
+ NAND2X1_LOC
XINVX1_LOC_42 INVX1_LOC_42/Y VSS VDD INVX1_LOC_42/A INVX1_LOC
XNAND2X1_LOC_652 NAND2X1_LOC_652/a_36_24# INVX1_LOC_513/A VSS VDD INVX1_LOC_348/Y
+ INVX1_LOC_460/Y NAND2X1_LOC
XNAND2X1_LOC_663 NAND2X1_LOC_663/a_36_24# GATE_662 VSS VDD INVX1_LOC_520/Y INVX1_LOC_523/Y
+ NAND2X1_LOC
XNAND2X1_LOC_641 NAND2X1_LOC_641/a_36_24# INVX1_LOC_501/A VSS VDD INVX1_LOC_203/Y
+ NAND2X1_LOC_267/A NAND2X1_LOC
XNAND2X1_LOC_630 NAND2X1_LOC_630/a_36_24# INVX1_LOC_488/A VSS VDD NAND2X1_LOC_628/Y
+ INVX1_LOC_487/Y NAND2X1_LOC
XINVX1_LOC_31 INVX1_LOC_31/Y VSS VDD INVX1_LOC_31/A INVX1_LOC
XINVX1_LOC_20 INVX1_LOC_20/Y VSS VDD INVX1_LOC_20/A INVX1_LOC
XNAND2X1_LOC_685 NAND2X1_LOC_685/a_36_24# INVX1_LOC_536/A VSS VDD NAND2X1_LOC_685/A
+ NAND2X1_LOC_685/B NAND2X1_LOC
XNAND2X1_LOC_696 NAND2X1_LOC_696/a_36_24# NAND2X1_LOC_708/A VSS VDD INVX1_LOC_35/Y
+ INVX1_LOC_395/A NAND2X1_LOC
XNAND2X1_LOC_674 NAND2X1_LOC_674/a_36_24# NAND2X1_LOC_675/B VSS VDD INVX1_LOC_74/Y
+ INVX1_LOC_532/Y NAND2X1_LOC
XINVX1_LOC_75 INVX1_LOC_75/Y VSS VDD INVX1_LOC_75/A INVX1_LOC
XINVX1_LOC_53 INVX1_LOC_53/Y VSS VDD INVX1_LOC_53/A INVX1_LOC
XINVX1_LOC_97 INVX1_LOC_97/Y VSS VDD INVX1_LOC_97/A INVX1_LOC
XINVX1_LOC_64 INVX1_LOC_64/Y VSS VDD INVX1_LOC_64/A INVX1_LOC
XINVX1_LOC_86 INVX1_LOC_86/Y VSS VDD INVX1_LOC_86/A INVX1_LOC
XINVX1_LOC_507 INVX1_LOC_507/Y VSS VDD INVX1_LOC_507/A INVX1_LOC
XINVX1_LOC_518 INVX1_LOC_518/Y VSS VDD INVX1_LOC_518/A INVX1_LOC
XINVX1_LOC_529 INVX1_LOC_529/Y VSS VDD INVX1_LOC_145/Y INVX1_LOC
XNAND2X1_LOC_471 NAND2X1_LOC_471/a_36_24# INVX1_LOC_377/A VSS VDD INVX1_LOC_370/Y
+ INVX1_LOC_371/Y NAND2X1_LOC
XNAND2X1_LOC_482 NAND2X1_LOC_482/a_36_24# NAND2X1_LOC_482/Y VSS VDD INVX1_LOC_11/Y
+ INVX1_LOC_63/Y NAND2X1_LOC
XNAND2X1_LOC_493 NAND2X1_LOC_493/a_36_24# INVX1_LOC_390/A VSS VDD NAND2X1_LOC_491/Y
+ NAND2X1_LOC_493/B NAND2X1_LOC
XNAND2X1_LOC_460 NAND2X1_LOC_460/a_36_24# INVX1_LOC_366/A VSS VDD NAND2X1_LOC_460/A
+ NAND2X1_LOC_409/Y NAND2X1_LOC
XINVX1_LOC_337 INVX1_LOC_337/Y VSS VDD INVX1_LOC_58/Y INVX1_LOC
XINVX1_LOC_348 INVX1_LOC_348/Y VSS VDD INVX1_LOC_348/A INVX1_LOC
XINVX1_LOC_359 INVX1_LOC_359/Y VSS VDD INVX1_LOC_359/A INVX1_LOC
XINVX1_LOC_304 INVX1_LOC_304/Y VSS VDD INVX1_LOC_304/A INVX1_LOC
XINVX1_LOC_315 INVX1_LOC_315/Y VSS VDD INVX1_LOC_315/A INVX1_LOC
XINVX1_LOC_326 INVX1_LOC_326/Y VSS VDD INVX1_LOC_326/A INVX1_LOC
XNAND2X1_LOC_290 NAND2X1_LOC_290/a_36_24# NAND2X1_LOC_334/A VSS VDD INVX1_LOC_79/A
+ INVX1_LOC_35/Y NAND2X1_LOC
XINVX1_LOC_101 INVX1_LOC_101/Y VSS VDD INVX1_LOC_80/A INVX1_LOC
XINVX1_LOC_112 INVX1_LOC_112/Y VSS VDD INVX1_LOC_17/Y INVX1_LOC
XINVX1_LOC_134 INVX1_LOC_134/Y VSS VDD INVX1_LOC_134/A INVX1_LOC
XINVX1_LOC_123 INVX1_LOC_479/A VSS VDD INVX1_LOC_123/A INVX1_LOC
XINVX1_LOC_189 INVX1_LOC_189/Y VSS VDD INVX1_LOC_189/A INVX1_LOC
XINVX1_LOC_167 INVX1_LOC_167/Y VSS VDD INVX1_LOC_167/A INVX1_LOC
XINVX1_LOC_156 INVX1_LOC_156/Y VSS VDD INVX1_LOC_156/A INVX1_LOC
XINVX1_LOC_145 INVX1_LOC_145/Y VSS VDD INVX1_LOC_145/A INVX1_LOC
XINVX1_LOC_178 INVX1_LOC_178/Y VSS VDD INVX1_LOC_178/A INVX1_LOC
XNAND2X1_LOC_801 NAND2X1_LOC_801/a_36_24# INVX1_LOC_631/A VSS VDD NAND2X1_LOC_801/A
+ INVX1_LOC_630/Y NAND2X1_LOC
XNAND2X1_LOC_834 NAND2X1_LOC_834/a_36_24# INVX1_LOC_655/A VSS VDD NAND2X1_LOC_513/A
+ NAND2X1_LOC_677/Y NAND2X1_LOC
XNAND2X1_LOC_812 NAND2X1_LOC_812/a_36_24# GATE_811 VSS VDD INVX1_LOC_640/Y INVX1_LOC_641/Y
+ NAND2X1_LOC
XNAND2X1_LOC_823 NAND2X1_LOC_823/a_36_24# NAND2X1_LOC_823/Y VSS VDD INVX1_LOC_58/Y
+ INVX1_LOC_206/Y NAND2X1_LOC
XNAND2X1_LOC_845 NAND2X1_LOC_845/a_36_24# INVX1_LOC_666/A VSS VDD INVX1_LOC_531/Y
+ NAND2X1_LOC_845/B NAND2X1_LOC
XNAND2X1_LOC_856 NAND2X1_LOC_856/a_36_24# INVX1_LOC_677/A VSS VDD INVX1_LOC_675/Y
+ INVX1_LOC_676/Y NAND2X1_LOC
XNAND2X1_LOC_119 NAND2X1_LOC_119/a_36_24# INVX1_LOC_110/A VSS VDD INPUT_1 INVX1_LOC_21/Y
+ NAND2X1_LOC
XNAND2X1_LOC_108 NAND2X1_LOC_108/a_36_24# NAND2X1_LOC_108/Y VSS VDD INVX1_LOC_63/Y
+ INVX1_LOC_99/Y NAND2X1_LOC
XNAND2X1_LOC_6 NAND2X1_LOC_6/a_36_24# INVX1_LOC_11/A VSS VDD INVX1_LOC_7/Y INVX1_LOC_9/Y
+ NAND2X1_LOC
XINVX1_LOC_10 INVX1_LOC_10/Y VSS VDD INPUT_2 INVX1_LOC
XINVX1_LOC_21 INVX1_LOC_21/Y VSS VDD INVX1_LOC_21/A INVX1_LOC
XNAND2X1_LOC_686 NAND2X1_LOC_686/a_36_24# INVX1_LOC_537/A VSS VDD NAND2X1_LOC_686/A
+ NAND2X1_LOC_686/B NAND2X1_LOC
XNAND2X1_LOC_653 NAND2X1_LOC_653/a_36_24# INVX1_LOC_514/A VSS VDD NAND2X1_LOC_594/Y
+ INVX1_LOC_513/Y NAND2X1_LOC
XNAND2X1_LOC_697 NAND2X1_LOC_697/a_36_24# NAND2X1_LOC_697/Y VSS VDD INVX1_LOC_145/Y
+ INVX1_LOC_206/Y NAND2X1_LOC
XNAND2X1_LOC_675 NAND2X1_LOC_675/a_36_24# INVX1_LOC_533/A VSS VDD INVX1_LOC_347/Y
+ NAND2X1_LOC_675/B NAND2X1_LOC
XNAND2X1_LOC_642 NAND2X1_LOC_642/a_36_24# INVX1_LOC_502/A VSS VDD NAND2X1_LOC_416/Y
+ INVX1_LOC_405/Y NAND2X1_LOC
XNAND2X1_LOC_620 NAND2X1_LOC_620/a_36_24# INVX1_LOC_482/A VSS VDD NAND2X1_LOC_528/Y
+ NAND2X1_LOC_613/Y NAND2X1_LOC
XNAND2X1_LOC_631 NAND2X1_LOC_631/a_36_24# INVX1_LOC_489/A VSS VDD INVX1_LOC_386/Y
+ NAND2X1_LOC_631/B NAND2X1_LOC
XNAND2X1_LOC_664 NAND2X1_LOC_664/a_36_24# NAND2X1_LOC_755/B VSS VDD INVX1_LOC_524/Y
+ INVX1_LOC_525/Y NAND2X1_LOC
XINVX1_LOC_76 INVX1_LOC_76/Y VSS VDD INVX1_LOC_76/A INVX1_LOC
XINVX1_LOC_65 INVX1_LOC_65/Y VSS VDD INVX1_LOC_65/A INVX1_LOC
XINVX1_LOC_32 INVX1_LOC_32/Y VSS VDD INVX1_LOC_32/A INVX1_LOC
XINVX1_LOC_43 INVX1_LOC_43/Y VSS VDD INVX1_LOC_43/A INVX1_LOC
XINVX1_LOC_54 INVX1_LOC_54/Y VSS VDD INVX1_LOC_54/A INVX1_LOC
XINVX1_LOC_98 INVX1_LOC_98/Y VSS VDD INVX1_LOC_98/A INVX1_LOC
XINVX1_LOC_87 INVX1_LOC_87/Y VSS VDD INVX1_LOC_87/A INVX1_LOC
XINVX1_LOC_508 INVX1_LOC_508/Y VSS VDD INVX1_LOC_508/A INVX1_LOC
XINVX1_LOC_519 INVX1_LOC_519/Y VSS VDD INVX1_LOC_519/A INVX1_LOC
XNAND2X1_LOC_450 NAND2X1_LOC_450/a_36_24# INVX1_LOC_356/A VSS VDD NAND2X1_LOC_426/Y
+ NAND2X1_LOC_427/Y NAND2X1_LOC
XNAND2X1_LOC_461 NAND2X1_LOC_461/a_36_24# INVX1_LOC_367/A VSS VDD NAND2X1_LOC_411/Y
+ NAND2X1_LOC_413/Y NAND2X1_LOC
XNAND2X1_LOC_483 NAND2X1_LOC_483/a_36_24# INVX1_LOC_386/A VSS VDD NAND2X1_LOC_252/Y
+ NAND2X1_LOC_482/Y NAND2X1_LOC
XNAND2X1_LOC_494 NAND2X1_LOC_494/a_36_24# NAND2X1_LOC_558/B VSS VDD INVX1_LOC_20/Y
+ NAND2X1_LOC_383/Y NAND2X1_LOC
XNAND2X1_LOC_472 NAND2X1_LOC_472/a_36_24# INVX1_LOC_378/A VSS VDD INVX1_LOC_368/Y
+ INVX1_LOC_369/Y NAND2X1_LOC
XINVX1_LOC_316 INVX1_LOC_316/Y VSS VDD INPUT_4 INVX1_LOC
XINVX1_LOC_305 INVX1_LOC_305/Y VSS VDD INVX1_LOC_41/Y INVX1_LOC
XINVX1_LOC_338 INVX1_LOC_338/Y VSS VDD INVX1_LOC_338/A INVX1_LOC
XINVX1_LOC_349 INVX1_LOC_349/Y VSS VDD INVX1_LOC_349/A INVX1_LOC
XINVX1_LOC_327 INVX1_LOC_327/Y VSS VDD INVX1_LOC_327/A INVX1_LOC
XNAND2X1_LOC_280 NAND2X1_LOC_280/a_36_24# NAND2X1_LOC_542/A VSS VDD INVX1_LOC_53/Y
+ INVX1_LOC_206/Y NAND2X1_LOC
XNAND2X1_LOC_291 NAND2X1_LOC_291/a_36_24# NAND2X1_LOC_334/B VSS VDD INVX1_LOC_45/Y
+ INVX1_LOC_204/Y NAND2X1_LOC
XINVX1_LOC_102 INVX1_LOC_102/Y VSS VDD INVX1_LOC_100/Y INVX1_LOC
XINVX1_LOC_135 INVX1_LOC_135/Y VSS VDD INVX1_LOC_62/Y INVX1_LOC
XINVX1_LOC_168 INVX1_LOC_168/Y VSS VDD INVX1_LOC_168/A INVX1_LOC
XINVX1_LOC_146 INVX1_LOC_586/A VSS VDD INVX1_LOC_146/A INVX1_LOC
XINVX1_LOC_124 INVX1_LOC_124/Y VSS VDD INVX1_LOC_124/A INVX1_LOC
XINVX1_LOC_113 INVX1_LOC_113/Y VSS VDD INVX1_LOC_47/Y INVX1_LOC
XINVX1_LOC_157 INVX1_LOC_157/Y VSS VDD INVX1_LOC_157/A INVX1_LOC
XINVX1_LOC_179 INVX1_LOC_179/Y VSS VDD INVX1_LOC_179/A INVX1_LOC
XINVX1_LOC_680 INVX1_LOC_680/Y VSS VDD INVX1_LOC_680/A INVX1_LOC
XNAND2X1_LOC_846 NAND2X1_LOC_846/a_36_24# INVX1_LOC_667/A VSS VDD NAND2X1_LOC_846/A
+ NAND2X1_LOC_846/B NAND2X1_LOC
XNAND2X1_LOC_802 NAND2X1_LOC_802/a_36_24# INVX1_LOC_632/A VSS VDD INVX1_LOC_628/Y
+ INVX1_LOC_629/Y NAND2X1_LOC
XNAND2X1_LOC_857 NAND2X1_LOC_857/a_36_24# INVX1_LOC_678/A VSS VDD INVX1_LOC_673/Y
+ INVX1_LOC_674/Y NAND2X1_LOC
XNAND2X1_LOC_835 NAND2X1_LOC_835/a_36_24# INVX1_LOC_656/A VSS VDD NAND2X1_LOC_835/A
+ NAND2X1_LOC_822/Y NAND2X1_LOC
XNAND2X1_LOC_824 NAND2X1_LOC_824/a_36_24# NAND2X1_LOC_836/B VSS VDD INVX1_LOC_35/Y
+ INVX1_LOC_204/Y NAND2X1_LOC
XNAND2X1_LOC_813 NAND2X1_LOC_813/a_36_24# NAND2X1_LOC_845/B VSS VDD INVX1_LOC_642/Y
+ INVX1_LOC_223/Y NAND2X1_LOC
XNAND2X1_LOC_109 NAND2X1_LOC_109/a_36_24# NAND2X1_LOC_775/B VSS VDD INVX1_LOC_41/Y
+ INVX1_LOC_80/A NAND2X1_LOC
XNAND2X1_LOC_7 NAND2X1_LOC_7/a_36_24# NAND2X1_LOC_7/Y VSS VDD INVX1_LOC_6/Y INVX1_LOC_11/Y
+ NAND2X1_LOC
XINVX1_LOC_22 INVX1_LOC_22/Y VSS VDD INPUT_2 INVX1_LOC
XNAND2X1_LOC_643 NAND2X1_LOC_643/a_36_24# INVX1_LOC_503/A VSS VDD INVX1_LOC_410/Y
+ NAND2X1_LOC_595/Y NAND2X1_LOC
XNAND2X1_LOC_687 NAND2X1_LOC_687/a_36_24# INVX1_LOC_538/A VSS VDD INVX1_LOC_536/Y
+ INVX1_LOC_537/Y NAND2X1_LOC
XNAND2X1_LOC_676 NAND2X1_LOC_676/a_36_24# NAND2X1_LOC_679/A VSS VDD INVX1_LOC_534/Y
+ INVX1_LOC_463/Y NAND2X1_LOC
XNAND2X1_LOC_654 NAND2X1_LOC_654/a_36_24# INVX1_LOC_515/A VSS VDD INVX1_LOC_511/Y
+ INVX1_LOC_512/Y NAND2X1_LOC
XNAND2X1_LOC_610 NAND2X1_LOC_610/a_36_24# NAND2X1_LOC_612/A VSS VDD INVX1_LOC_474/Y
+ INVX1_LOC_475/Y NAND2X1_LOC
XNAND2X1_LOC_632 NAND2X1_LOC_632/a_36_24# INVX1_LOC_490/A VSS VDD INVX1_LOC_488/Y
+ INVX1_LOC_489/Y NAND2X1_LOC
XNAND2X1_LOC_665 NAND2X1_LOC_665/a_36_24# NAND2X1_LOC_719/A VSS VDD INVX1_LOC_6/Y
+ NAND2X1_LOC_755/B NAND2X1_LOC
XNAND2X1_LOC_698 NAND2X1_LOC_698/a_36_24# NAND2X1_LOC_698/Y VSS VDD INVX1_LOC_69/Y
+ INVX1_LOC_117/Y NAND2X1_LOC
XNAND2X1_LOC_621 NAND2X1_LOC_621/a_36_24# INVX1_LOC_483/A VSS VDD NAND2X1_LOC_616/Y
+ NAND2X1_LOC_621/B NAND2X1_LOC
XINVX1_LOC_66 INVX1_LOC_66/Y VSS VDD INVX1_LOC_66/A INVX1_LOC
XINVX1_LOC_99 INVX1_LOC_99/Y VSS VDD INVX1_LOC_99/A INVX1_LOC
XINVX1_LOC_77 INVX1_LOC_77/Y VSS VDD INVX1_LOC_77/A INVX1_LOC
XINVX1_LOC_88 INVX1_LOC_88/Y VSS VDD INVX1_LOC_54/Y INVX1_LOC
XINVX1_LOC_11 INVX1_LOC_11/Y VSS VDD INVX1_LOC_11/A INVX1_LOC
XINVX1_LOC_55 INVX1_LOC_55/Y VSS VDD INVX1_LOC_55/A INVX1_LOC
XINVX1_LOC_33 INVX1_LOC_33/Y VSS VDD INVX1_LOC_33/A INVX1_LOC
XINVX1_LOC_44 INVX1_LOC_44/Y VSS VDD INVX1_LOC_44/A INVX1_LOC
XINVX1_LOC_509 INVX1_LOC_509/Y VSS VDD INVX1_LOC_509/A INVX1_LOC
XNAND2X1_LOC_440 NAND2X1_LOC_440/a_36_24# INVX1_LOC_348/A VSS VDD NAND2X1_LOC_440/A
+ INVX1_LOC_347/Y NAND2X1_LOC
XNAND2X1_LOC_451 NAND2X1_LOC_451/a_36_24# INVX1_LOC_357/A VSS VDD NAND2X1_LOC_428/Y
+ NAND2X1_LOC_451/B NAND2X1_LOC
XNAND2X1_LOC_484 NAND2X1_LOC_484/a_36_24# NAND2X1_LOC_486/A VSS VDD INVX1_LOC_17/Y
+ INVX1_LOC_45/Y NAND2X1_LOC
XNAND2X1_LOC_495 NAND2X1_LOC_495/a_36_24# NAND2X1_LOC_833/B VSS VDD INVX1_LOC_45/Y
+ INVX1_LOC_62/Y NAND2X1_LOC
XNAND2X1_LOC_473 NAND2X1_LOC_473/a_36_24# INVX1_LOC_379/A VSS VDD INVX1_LOC_109/Y
+ INVX1_LOC_235/Y NAND2X1_LOC
XNAND2X1_LOC_462 NAND2X1_LOC_462/a_36_24# INVX1_LOC_368/A VSS VDD NAND2X1_LOC_416/Y
+ INVX1_LOC_367/Y NAND2X1_LOC
XINVX1_LOC_317 INVX1_LOC_317/Y VSS VDD INVX1_LOC_317/A INVX1_LOC
XINVX1_LOC_339 INVX1_LOC_339/Y VSS VDD INVX1_LOC_245/A INVX1_LOC
XINVX1_LOC_306 INVX1_LOC_306/Y VSS VDD INVX1_LOC_145/Y INVX1_LOC
XINVX1_LOC_328 INVX1_LOC_328/Y VSS VDD INVX1_LOC_328/A INVX1_LOC
XNAND2X1_LOC_270 NAND2X1_LOC_270/a_36_24# NAND2X1_LOC_271/B VSS VDD INVX1_LOC_232/Y
+ INVX1_LOC_233/Y NAND2X1_LOC
XNAND2X1_LOC_281 NAND2X1_LOC_281/a_36_24# NAND2X1_LOC_285/A VSS VDD INVX1_LOC_6/Y
+ INVX1_LOC_206/Y NAND2X1_LOC
XNAND2X1_LOC_292 NAND2X1_LOC_292/a_36_24# NAND2X1_LOC_292/Y VSS VDD INVX1_LOC_48/Y
+ INVX1_LOC_134/Y NAND2X1_LOC
XINVX1_LOC_147 INVX1_LOC_147/Y VSS VDD INVX1_LOC_147/A INVX1_LOC
XINVX1_LOC_136 INVX1_LOC_136/Y VSS VDD INVX1_LOC_134/Y INVX1_LOC
XINVX1_LOC_125 INVX1_LOC_125/Y VSS VDD INVX1_LOC_125/A INVX1_LOC
XINVX1_LOC_114 INVX1_LOC_114/Y VSS VDD INVX1_LOC_114/A INVX1_LOC
XINVX1_LOC_103 INVX1_LOC_103/Y VSS VDD INVX1_LOC_103/A INVX1_LOC
XINVX1_LOC_158 INVX1_LOC_158/Y VSS VDD INVX1_LOC_158/A INVX1_LOC
XINVX1_LOC_169 INVX1_LOC_169/Y VSS VDD INVX1_LOC_169/A INVX1_LOC
XINVX1_LOC_670 INVX1_LOC_670/Y VSS VDD INVX1_LOC_670/A INVX1_LOC
XINVX1_LOC_681 INVX1_LOC_681/Y VSS VDD INVX1_LOC_681/A INVX1_LOC
XNAND2X1_LOC_803 NAND2X1_LOC_803/a_36_24# INVX1_LOC_633/A VSS VDD INVX1_LOC_626/Y
+ INVX1_LOC_627/Y NAND2X1_LOC
XNAND2X1_LOC_814 NAND2X1_LOC_814/a_36_24# NAND2X1_LOC_814/Y VSS VDD INVX1_LOC_643/Y
+ INVX1_LOC_644/Y NAND2X1_LOC
XNAND2X1_LOC_847 NAND2X1_LOC_847/a_36_24# INVX1_LOC_668/A VSS VDD NAND2X1_LOC_847/A
+ NAND2X1_LOC_820/Y NAND2X1_LOC
XNAND2X1_LOC_858 NAND2X1_LOC_858/a_36_24# INVX1_LOC_679/A VSS VDD INVX1_LOC_671/Y
+ INVX1_LOC_672/Y NAND2X1_LOC
XNAND2X1_LOC_825 NAND2X1_LOC_825/a_36_24# NAND2X1_LOC_837/A VSS VDD INVX1_LOC_50/Y
+ INVX1_LOC_91/Y NAND2X1_LOC
XNAND2X1_LOC_836 NAND2X1_LOC_836/a_36_24# INVX1_LOC_657/A VSS VDD NAND2X1_LOC_823/Y
+ NAND2X1_LOC_836/B NAND2X1_LOC
XNAND2X1_LOC_8 NAND2X1_LOC_8/a_36_24# INVX1_LOC_12/A VSS VDD INPUT_2 INVX1_LOC_13/Y
+ NAND2X1_LOC
XNAND2X1_LOC_600 NAND2X1_LOC_600/a_36_24# NAND2X1_LOC_602/A VSS VDD INVX1_LOC_41/Y
+ INVX1_LOC_100/Y NAND2X1_LOC
XNAND2X1_LOC_611 NAND2X1_LOC_611/a_36_24# INVX1_LOC_476/A VSS VDD INVX1_LOC_9/Y INVX1_LOC_477/Y
+ NAND2X1_LOC
XINVX1_LOC_23 INVX1_LOC_23/Y VSS VDD INPUT_3 INVX1_LOC
XNAND2X1_LOC_644 NAND2X1_LOC_644/a_36_24# INVX1_LOC_504/A VSS VDD NAND2X1_LOC_597/Y
+ INVX1_LOC_505/Y NAND2X1_LOC
XNAND2X1_LOC_655 NAND2X1_LOC_655/a_36_24# INVX1_LOC_516/A VSS VDD INVX1_LOC_509/Y
+ INVX1_LOC_510/Y NAND2X1_LOC
XNAND2X1_LOC_688 NAND2X1_LOC_688/a_36_24# NAND2X1_LOC_689/B VSS VDD INVX1_LOC_539/Y
+ INVX1_LOC_540/Y NAND2X1_LOC
XNAND2X1_LOC_633 NAND2X1_LOC_633/a_36_24# INVX1_LOC_491/A VSS VDD NAND2X1_LOC_123/B
+ INVX1_LOC_492/Y NAND2X1_LOC
XNAND2X1_LOC_677 NAND2X1_LOC_677/a_36_24# NAND2X1_LOC_677/Y VSS VDD INVX1_LOC_35/Y
+ INVX1_LOC_479/A NAND2X1_LOC
XNAND2X1_LOC_666 NAND2X1_LOC_666/a_36_24# NAND2X1_LOC_666/Y VSS VDD INVX1_LOC_26/Y
+ INVX1_LOC_526/Y NAND2X1_LOC
XNAND2X1_LOC_622 NAND2X1_LOC_622/a_36_24# INVX1_LOC_484/A VSS VDD NAND2X1_LOC_619/Y
+ INVX1_LOC_483/Y NAND2X1_LOC
XNAND2X1_LOC_699 NAND2X1_LOC_699/a_36_24# INVX1_LOC_543/A VSS VDD INVX1_LOC_21/Y INVX1_LOC_145/Y
+ NAND2X1_LOC
XINVX1_LOC_89 INVX1_LOC_89/Y VSS VDD INVX1_LOC_89/A INVX1_LOC
XINVX1_LOC_78 INVX1_LOC_80/A VSS VDD INVX1_LOC_78/A INVX1_LOC
XINVX1_LOC_67 INVX1_LOC_67/Y VSS VDD INVX1_LOC_92/A INVX1_LOC
XINVX1_LOC_45 INVX1_LOC_45/Y VSS VDD INVX1_LOC_45/A INVX1_LOC
XINVX1_LOC_12 INVX1_LOC_12/Y VSS VDD INVX1_LOC_12/A INVX1_LOC
XINVX1_LOC_56 INVX1_LOC_56/Y VSS VDD INPUT_6 INVX1_LOC
XINVX1_LOC_34 INVX1_LOC_34/Y VSS VDD INPUT_7 INVX1_LOC
XNAND2X1_LOC_452 NAND2X1_LOC_452/a_36_24# INVX1_LOC_358/A VSS VDD INVX1_LOC_356/Y
+ INVX1_LOC_357/Y NAND2X1_LOC
XNAND2X1_LOC_441 NAND2X1_LOC_441/a_36_24# NAND2X1_LOC_545/A VSS VDD INVX1_LOC_48/Y
+ INVX1_LOC_54/Y NAND2X1_LOC
XNAND2X1_LOC_430 NAND2X1_LOC_430/a_36_24# NAND2X1_LOC_451/B VSS VDD INVX1_LOC_586/A
+ INVX1_LOC_342/Y NAND2X1_LOC
XNAND2X1_LOC_463 NAND2X1_LOC_463/a_36_24# INVX1_LOC_369/A VSS VDD INVX1_LOC_365/Y
+ INVX1_LOC_366/Y NAND2X1_LOC
XNAND2X1_LOC_485 NAND2X1_LOC_485/a_36_24# NAND2X1_LOC_486/B VSS VDD INVX1_LOC_50/Y
+ INVX1_LOC_99/Y NAND2X1_LOC
XNAND2X1_LOC_496 NAND2X1_LOC_496/a_36_24# NAND2X1_LOC_496/Y VSS VDD INVX1_LOC_26/Y
+ INVX1_LOC_62/Y NAND2X1_LOC
XNAND2X1_LOC_474 NAND2X1_LOC_474/a_36_24# INVX1_LOC_380/A VSS VDD INVX1_LOC_321/Y
+ INVX1_LOC_328/Y NAND2X1_LOC
XINVX1_LOC_329 INVX1_LOC_329/Y VSS VDD INVX1_LOC_51/Y INVX1_LOC
XINVX1_LOC_318 INVX1_LOC_318/Y VSS VDD INVX1_LOC_318/A INVX1_LOC
XINVX1_LOC_307 INVX1_LOC_307/Y VSS VDD INVX1_LOC_307/A INVX1_LOC
XNAND2X1_LOC_282 NAND2X1_LOC_282/a_36_24# NAND2X1_LOC_285/B VSS VDD INVX1_LOC_99/Y
+ INVX1_LOC_145/Y NAND2X1_LOC
XNAND2X1_LOC_260 NAND2X1_LOC_260/a_36_24# NAND2X1_LOC_260/Y VSS VDD INVX1_LOC_221/Y
+ INVX1_LOC_222/Y NAND2X1_LOC
XNAND2X1_LOC_271 NAND2X1_LOC_271/a_36_24# NAND2X1_LOC_276/A VSS VDD NAND2X1_LOC_271/A
+ NAND2X1_LOC_271/B NAND2X1_LOC
XNAND2X1_LOC_293 NAND2X1_LOC_293/a_36_24# INVX1_LOC_243/A VSS VDD INPUT_1 INVX1_LOC_9/Y
+ NAND2X1_LOC
XINVX1_LOC_137 INVX1_LOC_137/Y VSS VDD INVX1_LOC_137/A INVX1_LOC
XINVX1_LOC_148 INVX1_LOC_148/Y VSS VDD INVX1_LOC_32/Y INVX1_LOC
XINVX1_LOC_126 INVX1_LOC_126/Y VSS VDD INVX1_LOC_126/A INVX1_LOC
XINVX1_LOC_104 INVX1_LOC_104/Y VSS VDD INPUT_0 INVX1_LOC
XINVX1_LOC_115 INVX1_LOC_115/Y VSS VDD INVX1_LOC_115/A INVX1_LOC
XINVX1_LOC_159 INVX1_LOC_159/Y VSS VDD INVX1_LOC_159/A INVX1_LOC
XINVX1_LOC_671 INVX1_LOC_671/Y VSS VDD INVX1_LOC_671/A INVX1_LOC
XINVX1_LOC_682 INVX1_LOC_682/Y VSS VDD INVX1_LOC_682/A INVX1_LOC
XINVX1_LOC_660 INVX1_LOC_660/Y VSS VDD INVX1_LOC_660/A INVX1_LOC
XNAND2X1_LOC_804 NAND2X1_LOC_804/a_36_24# INVX1_LOC_634/A VSS VDD INVX1_LOC_624/Y
+ INVX1_LOC_625/Y NAND2X1_LOC
XNAND2X1_LOC_859 NAND2X1_LOC_859/a_36_24# INVX1_LOC_680/A VSS VDD INVX1_LOC_669/Y
+ INVX1_LOC_670/Y NAND2X1_LOC
XNAND2X1_LOC_815 NAND2X1_LOC_815/a_36_24# NAND2X1_LOC_846/A VSS VDD INVX1_LOC_6/Y
+ NAND2X1_LOC_814/Y NAND2X1_LOC
XNAND2X1_LOC_848 NAND2X1_LOC_848/a_36_24# INVX1_LOC_669/A VSS VDD INVX1_LOC_667/Y
+ INVX1_LOC_668/Y NAND2X1_LOC
XNAND2X1_LOC_837 NAND2X1_LOC_837/a_36_24# INVX1_LOC_658/A VSS VDD NAND2X1_LOC_837/A
+ NAND2X1_LOC_837/B NAND2X1_LOC
XNAND2X1_LOC_826 NAND2X1_LOC_826/a_36_24# NAND2X1_LOC_837/B VSS VDD INVX1_LOC_62/Y
+ INVX1_LOC_93/Y NAND2X1_LOC
XINVX1_LOC_490 INVX1_LOC_490/Y VSS VDD INVX1_LOC_490/A INVX1_LOC
XNAND2X1_LOC_9 NAND2X1_LOC_9/a_36_24# INVX1_LOC_14/A VSS VDD INVX1_LOC_15/Y INVX1_LOC_16/Y
+ NAND2X1_LOC
XINVX1_LOC_13 INVX1_LOC_13/Y VSS VDD INPUT_3 INVX1_LOC
XNAND2X1_LOC_601 NAND2X1_LOC_601/a_36_24# NAND2X1_LOC_601/Y VSS VDD INVX1_LOC_79/A
+ INVX1_LOC_53/Y NAND2X1_LOC
XNAND2X1_LOC_645 NAND2X1_LOC_645/a_36_24# INVX1_LOC_506/A VSS VDD INVX1_LOC_468/Y
+ INVX1_LOC_469/Y NAND2X1_LOC
XNAND2X1_LOC_634 NAND2X1_LOC_634/a_36_24# INVX1_LOC_493/A VSS VDD NAND2X1_LOC_334/A
+ INVX1_LOC_494/Y NAND2X1_LOC
XNAND2X1_LOC_612 NAND2X1_LOC_612/a_36_24# NAND2X1_LOC_647/A VSS VDD NAND2X1_LOC_612/A
+ INVX1_LOC_476/Y NAND2X1_LOC
XNAND2X1_LOC_623 NAND2X1_LOC_623/a_36_24# INVX1_LOC_485/A VSS VDD NAND2X1_LOC_615/Y
+ INVX1_LOC_482/Y NAND2X1_LOC
XINVX1_LOC_24 INVX1_LOC_79/A VSS VDD INVX1_LOC_24/A INVX1_LOC
XNAND2X1_LOC_689 NAND2X1_LOC_689/a_36_24# NAND2X1_LOC_691/A VSS VDD INVX1_LOC_41/Y
+ NAND2X1_LOC_689/B NAND2X1_LOC
XNAND2X1_LOC_656 NAND2X1_LOC_656/a_36_24# INVX1_LOC_517/A VSS VDD INVX1_LOC_98/Y INVX1_LOC_508/Y
+ NAND2X1_LOC
XNAND2X1_LOC_678 NAND2X1_LOC_678/a_36_24# NAND2X1_LOC_679/B VSS VDD INVX1_LOC_535/Y
+ NAND2X1_LOC_677/Y NAND2X1_LOC
XNAND2X1_LOC_667 NAND2X1_LOC_667/a_36_24# NAND2X1_LOC_720/A VSS VDD INVX1_LOC_69/Y
+ INVX1_LOC_527/Y NAND2X1_LOC
XINVX1_LOC_68 INVX1_LOC_68/Y VSS VDD INVX1_LOC_68/A INVX1_LOC
XINVX1_LOC_35 INVX1_LOC_35/Y VSS VDD INVX1_LOC_35/A INVX1_LOC
XINVX1_LOC_79 INVX1_LOC_79/Y VSS VDD INVX1_LOC_79/A INVX1_LOC
XINVX1_LOC_46 INVX1_LOC_46/Y VSS VDD INVX1_LOC_46/A INVX1_LOC
XINVX1_LOC_57 INVX1_LOC_57/Y VSS VDD INPUT_7 INVX1_LOC
XNAND2X1_LOC_453 NAND2X1_LOC_453/a_36_24# INVX1_LOC_359/A VSS VDD INVX1_LOC_354/Y
+ INVX1_LOC_355/Y NAND2X1_LOC
XNAND2X1_LOC_431 NAND2X1_LOC_431/a_36_24# NAND2X1_LOC_434/B VSS VDD INVX1_LOC_74/Y
+ INVX1_LOC_206/Y NAND2X1_LOC
XNAND2X1_LOC_497 NAND2X1_LOC_497/a_36_24# NAND2X1_LOC_844/A VSS VDD INVX1_LOC_31/Y
+ INVX1_LOC_75/Y NAND2X1_LOC
XNAND2X1_LOC_486 NAND2X1_LOC_486/a_36_24# INVX1_LOC_387/A VSS VDD NAND2X1_LOC_486/A
+ NAND2X1_LOC_486/B NAND2X1_LOC
XNAND2X1_LOC_464 NAND2X1_LOC_464/a_36_24# INVX1_LOC_370/A VSS VDD INVX1_LOC_363/Y
+ INVX1_LOC_364/Y NAND2X1_LOC
XNAND2X1_LOC_442 NAND2X1_LOC_442/a_36_24# NAND2X1_LOC_444/A VSS VDD INVX1_LOC_48/Y
+ INVX1_LOC_100/Y NAND2X1_LOC
XNAND2X1_LOC_475 NAND2X1_LOC_475/a_36_24# INVX1_LOC_381/A VSS VDD NAND2X1_LOC_475/A
+ INVX1_LOC_380/Y NAND2X1_LOC
XNAND2X1_LOC_420 NAND2X1_LOC_420/a_36_24# NAND2X1_LOC_420/Y VSS VDD INVX1_LOC_93/Y
+ INVX1_LOC_99/Y NAND2X1_LOC
XINVX1_LOC_319 INVX1_LOC_319/Y VSS VDD INVX1_LOC_319/A INVX1_LOC
XINVX1_LOC_308 INVX1_LOC_308/Y VSS VDD INVX1_LOC_21/Y INVX1_LOC
XNAND2X1_LOC_272 NAND2X1_LOC_272/a_36_24# NAND2X1_LOC_541/B VSS VDD INVX1_LOC_41/Y
+ INVX1_LOC_49/Y NAND2X1_LOC
XNAND2X1_LOC_261 NAND2X1_LOC_261/a_36_24# NAND2X1_LOC_261/Y VSS VDD INVX1_LOC_100/Y
+ NAND2X1_LOC_260/Y NAND2X1_LOC
XNAND2X1_LOC_250 NAND2X1_LOC_250/a_36_24# NAND2X1_LOC_250/Y VSS VDD INVX1_LOC_69/Y
+ NAND2X1_LOC_249/Y NAND2X1_LOC
XNAND2X1_LOC_283 NAND2X1_LOC_283/a_36_24# NAND2X1_LOC_286/A VSS VDD INVX1_LOC_35/Y
+ INVX1_LOC_199/Y NAND2X1_LOC
XNAND2X1_LOC_294 NAND2X1_LOC_294/a_36_24# NAND2X1_LOC_294/Y VSS VDD INVX1_LOC_244/Y
+ INVX1_LOC_245/Y NAND2X1_LOC
XINVX1_LOC_105 INVX1_LOC_105/Y VSS VDD INVX1_LOC_105/A INVX1_LOC
XINVX1_LOC_116 INVX1_LOC_116/Y VSS VDD INVX1_LOC_116/A INVX1_LOC
XINVX1_LOC_138 INVX1_LOC_138/Y VSS VDD INPUT_1 INVX1_LOC
XINVX1_LOC_149 INVX1_LOC_149/Y VSS VDD INVX1_LOC_117/Y INVX1_LOC
XINVX1_LOC_127 INVX1_LOC_127/Y VSS VDD INVX1_LOC_127/A INVX1_LOC
XINVX1_LOC_650 INVX1_LOC_650/Y VSS VDD INVX1_LOC_92/A INVX1_LOC
XINVX1_LOC_672 INVX1_LOC_672/Y VSS VDD INVX1_LOC_672/A INVX1_LOC
XINVX1_LOC_661 INVX1_LOC_661/Y VSS VDD INVX1_LOC_661/A INVX1_LOC
XINVX1_LOC_683 INVX1_LOC_683/Y VSS VDD INVX1_LOC_683/A INVX1_LOC
XNAND2X1_LOC_816 NAND2X1_LOC_816/a_36_24# NAND2X1_LOC_846/B VSS VDD INVX1_LOC_58/Y
+ INVX1_LOC_645/Y NAND2X1_LOC
XNAND2X1_LOC_827 NAND2X1_LOC_827/a_36_24# NAND2X1_LOC_827/Y VSS VDD INVX1_LOC_49/Y
+ INVX1_LOC_145/Y NAND2X1_LOC
XNAND2X1_LOC_805 NAND2X1_LOC_805/a_36_24# INVX1_LOC_635/A VSS VDD INVX1_LOC_622/Y
+ INVX1_LOC_623/Y NAND2X1_LOC
XINVX1_LOC_491 INVX1_LOC_491/Y VSS VDD INVX1_LOC_491/A INVX1_LOC
XINVX1_LOC_480 INVX1_LOC_480/Y VSS VDD INVX1_LOC_480/A INVX1_LOC
XNAND2X1_LOC_849 NAND2X1_LOC_849/a_36_24# INVX1_LOC_670/A VSS VDD INVX1_LOC_665/Y
+ INVX1_LOC_666/Y NAND2X1_LOC
XNAND2X1_LOC_838 NAND2X1_LOC_838/a_36_24# INVX1_LOC_659/A VSS VDD NAND2X1_LOC_827/Y
+ INVX1_LOC_658/Y NAND2X1_LOC
XNAND2X1_LOC_657 NAND2X1_LOC_657/a_36_24# INVX1_LOC_518/A VSS VDD INVX1_LOC_128/Y
+ INVX1_LOC_400/Y NAND2X1_LOC
XNAND2X1_LOC_602 NAND2X1_LOC_602/a_36_24# INVX1_LOC_468/A VSS VDD NAND2X1_LOC_602/A
+ NAND2X1_LOC_601/Y NAND2X1_LOC
XNAND2X1_LOC_635 NAND2X1_LOC_635/a_36_24# INVX1_LOC_495/A VSS VDD NAND2X1_LOC_428/Y
+ NAND2X1_LOC_635/B NAND2X1_LOC
XNAND2X1_LOC_646 NAND2X1_LOC_646/a_36_24# INVX1_LOC_507/A VSS VDD NAND2X1_LOC_646/A
+ NAND2X1_LOC_646/B NAND2X1_LOC
XNAND2X1_LOC_679 NAND2X1_LOC_679/a_36_24# NAND2X1_LOC_728/A VSS VDD NAND2X1_LOC_679/A
+ NAND2X1_LOC_679/B NAND2X1_LOC
XNAND2X1_LOC_613 NAND2X1_LOC_613/a_36_24# NAND2X1_LOC_613/Y VSS VDD INVX1_LOC_48/Y
+ INVX1_LOC_62/Y NAND2X1_LOC
XNAND2X1_LOC_624 NAND2X1_LOC_624/a_36_24# INVX1_LOC_486/A VSS VDD INVX1_LOC_484/Y
+ INVX1_LOC_485/Y NAND2X1_LOC
XNAND2X1_LOC_668 NAND2X1_LOC_668/a_36_24# NAND2X1_LOC_668/Y VSS VDD INVX1_LOC_528/Y
+ INVX1_LOC_529/Y NAND2X1_LOC
XINVX1_LOC_14 INVX1_LOC_66/A VSS VDD INVX1_LOC_14/A INVX1_LOC
XINVX1_LOC_36 INVX1_LOC_84/A VSS VDD INVX1_LOC_36/A INVX1_LOC
XINVX1_LOC_47 INVX1_LOC_47/Y VSS VDD INVX1_LOC_47/A INVX1_LOC
XINVX1_LOC_58 INVX1_LOC_58/Y VSS VDD INVX1_LOC_58/A INVX1_LOC
XINVX1_LOC_25 INVX1_LOC_25/Y VSS VDD INVX1_LOC_25/A INVX1_LOC
XINVX1_LOC_69 INVX1_LOC_69/Y VSS VDD INVX1_LOC_69/A INVX1_LOC
XNAND2X1_LOC_465 NAND2X1_LOC_465/a_36_24# INVX1_LOC_371/A VSS VDD INVX1_LOC_361/Y
+ INVX1_LOC_362/Y NAND2X1_LOC
XNAND2X1_LOC_498 NAND2X1_LOC_498/a_36_24# NAND2X1_LOC_498/Y VSS VDD INVX1_LOC_74/Y
+ NAND2X1_LOC_498/B NAND2X1_LOC
XNAND2X1_LOC_432 NAND2X1_LOC_432/a_36_24# NAND2X1_LOC_432/Y VSS VDD INVX1_LOC_26/Y
+ INVX1_LOC_119/Y NAND2X1_LOC
XNAND2X1_LOC_410 NAND2X1_LOC_410/a_36_24# NAND2X1_LOC_410/Y VSS VDD INVX1_LOC_336/Y
+ INVX1_LOC_337/Y NAND2X1_LOC
XNAND2X1_LOC_421 NAND2X1_LOC_421/a_36_24# NAND2X1_LOC_448/A VSS VDD INVX1_LOC_89/Y
+ INVX1_LOC_261/Y NAND2X1_LOC
XNAND2X1_LOC_454 NAND2X1_LOC_454/a_36_24# INVX1_LOC_360/A VSS VDD INVX1_LOC_352/Y
+ INVX1_LOC_353/Y NAND2X1_LOC
XNAND2X1_LOC_443 NAND2X1_LOC_443/a_36_24# INVX1_LOC_349/A VSS VDD NAND2X1_LOC_97/B
+ NAND2X1_LOC_545/A NAND2X1_LOC
XNAND2X1_LOC_476 NAND2X1_LOC_476/a_36_24# INVX1_LOC_382/A VSS VDD INVX1_LOC_378/Y
+ INVX1_LOC_379/Y NAND2X1_LOC
XNAND2X1_LOC_487 NAND2X1_LOC_487/a_36_24# NAND2X1_LOC_489/A VSS VDD INVX1_LOC_32/Y
+ INVX1_LOC_93/Y NAND2X1_LOC
XINVX1_LOC_309 INVX1_LOC_309/Y VSS VDD INVX1_LOC_49/Y INVX1_LOC
XNAND2X1_LOC_273 NAND2X1_LOC_273/a_36_24# NAND2X1_LOC_274/B VSS VDD INVX1_LOC_45/Y
+ INVX1_LOC_137/Y NAND2X1_LOC
XNAND2X1_LOC_284 NAND2X1_LOC_284/a_36_24# INVX1_LOC_238/A VSS VDD NAND2X1_LOC_284/A
+ NAND2X1_LOC_542/A NAND2X1_LOC
XNAND2X1_LOC_251 NAND2X1_LOC_251/a_36_24# NAND2X1_LOC_843/A VSS VDD INVX1_LOC_58/Y
+ NAND2X1_LOC_106/B NAND2X1_LOC
XNAND2X1_LOC_295 NAND2X1_LOC_295/a_36_24# NAND2X1_LOC_346/B VSS VDD INVX1_LOC_63/Y
+ NAND2X1_LOC_294/Y NAND2X1_LOC
XNAND2X1_LOC_262 NAND2X1_LOC_262/a_36_24# NAND2X1_LOC_786/B VSS VDD INVX1_LOC_48/Y
+ INVX1_LOC_68/Y NAND2X1_LOC
XNAND2X1_LOC_240 NAND2X1_LOC_240/a_36_24# INVX1_LOC_207/A VSS VDD NAND2X1_LOC_240/A
+ NAND2X1_LOC_234/Y NAND2X1_LOC
XINVX1_LOC_117 INVX1_LOC_117/Y VSS VDD INVX1_LOC_117/A INVX1_LOC
XINVX1_LOC_106 INVX1_LOC_106/Y VSS VDD INVX1_LOC_106/A INVX1_LOC
XINVX1_LOC_139 INVX1_LOC_139/Y VSS VDD INVX1_LOC_139/A INVX1_LOC
XINVX1_LOC_128 INVX1_LOC_128/Y VSS VDD INVX1_LOC_128/A INVX1_LOC
XINVX1_LOC_662 INVX1_LOC_662/Y VSS VDD INVX1_LOC_662/A INVX1_LOC
XINVX1_LOC_651 INVX1_LOC_651/Y VSS VDD INVX1_LOC_651/A INVX1_LOC
XINVX1_LOC_640 INVX1_LOC_640/Y VSS VDD INVX1_LOC_640/A INVX1_LOC
XINVX1_LOC_684 INVX1_LOC_684/Y VSS VDD INVX1_LOC_684/A INVX1_LOC
XINVX1_LOC_673 INVX1_LOC_673/Y VSS VDD INVX1_LOC_673/A INVX1_LOC
XNAND2X1_LOC_828 NAND2X1_LOC_828/a_36_24# NAND2X1_LOC_829/B VSS VDD INVX1_LOC_335/A
+ INVX1_LOC_463/Y NAND2X1_LOC
XNAND2X1_LOC_817 NAND2X1_LOC_817/a_36_24# NAND2X1_LOC_847/A VSS VDD INVX1_LOC_646/Y
+ INVX1_LOC_312/Y NAND2X1_LOC
XNAND2X1_LOC_806 NAND2X1_LOC_806/a_36_24# INVX1_LOC_636/A VSS VDD INVX1_LOC_242/Y
+ INVX1_LOC_533/Y NAND2X1_LOC
XNAND2X1_LOC_839 NAND2X1_LOC_839/a_36_24# INVX1_LOC_660/A VSS VDD INVX1_LOC_656/Y
+ INVX1_LOC_657/Y NAND2X1_LOC
XINVX1_LOC_492 INVX1_LOC_492/Y VSS VDD INVX1_LOC_492/A INVX1_LOC
XINVX1_LOC_470 INVX1_LOC_470/Y VSS VDD INVX1_LOC_99/Y INVX1_LOC
XINVX1_LOC_481 INVX1_LOC_481/Y VSS VDD INPUT_3 INVX1_LOC
XNAND2X1_LOC_603 NAND2X1_LOC_603/a_36_24# NAND2X1_LOC_603/Y VSS VDD INVX1_LOC_20/Y
+ INVX1_LOC_54/Y NAND2X1_LOC
XNAND2X1_LOC_636 NAND2X1_LOC_636/a_36_24# INVX1_LOC_496/A VSS VDD NAND2X1_LOC_636/A
+ NAND2X1_LOC_636/B NAND2X1_LOC
XNAND2X1_LOC_647 NAND2X1_LOC_647/a_36_24# INVX1_LOC_508/A VSS VDD NAND2X1_LOC_647/A
+ INVX1_LOC_507/Y NAND2X1_LOC
XNAND2X1_LOC_658 NAND2X1_LOC_658/a_36_24# INVX1_LOC_519/A VSS VDD INVX1_LOC_486/Y
+ INVX1_LOC_490/Y NAND2X1_LOC
XNAND2X1_LOC_614 NAND2X1_LOC_614/a_36_24# NAND2X1_LOC_615/B VSS VDD INVX1_LOC_478/Y
+ INVX1_LOC_479/Y NAND2X1_LOC
XNAND2X1_LOC_669 NAND2X1_LOC_669/a_36_24# NAND2X1_LOC_669/Y VSS VDD INVX1_LOC_586/A
+ NAND2X1_LOC_668/Y NAND2X1_LOC
XNAND2X1_LOC_625 NAND2X1_LOC_625/a_36_24# NAND2X1_LOC_631/B VSS VDD NAND2X1_LOC_66/Y
+ INVX1_LOC_245/A NAND2X1_LOC
XINVX1_LOC_15 INVX1_LOC_15/Y VSS VDD INPUT_0 INVX1_LOC
XINVX1_LOC_59 INVX1_LOC_59/Y VSS VDD INVX1_LOC_59/A INVX1_LOC
XINVX1_LOC_37 INVX1_LOC_37/Y VSS VDD INPUT_0 INVX1_LOC
XINVX1_LOC_26 INVX1_LOC_26/Y VSS VDD INVX1_LOC_26/A INVX1_LOC
XINVX1_LOC_48 INVX1_LOC_48/Y VSS VDD INVX1_LOC_48/A INVX1_LOC
XNAND2X1_LOC_411 NAND2X1_LOC_411/a_36_24# NAND2X1_LOC_411/Y VSS VDD INVX1_LOC_100/Y
+ NAND2X1_LOC_410/Y NAND2X1_LOC
XNAND2X1_LOC_400 NAND2X1_LOC_400/a_36_24# INVX1_LOC_324/A VSS VDD NAND2X1_LOC_393/Y
+ NAND2X1_LOC_400/B NAND2X1_LOC
XNAND2X1_LOC_466 NAND2X1_LOC_466/a_36_24# INVX1_LOC_372/A VSS VDD INVX1_LOC_359/Y
+ INVX1_LOC_360/Y NAND2X1_LOC
XNAND2X1_LOC_477 NAND2X1_LOC_477/a_36_24# INVX1_LOC_383/A VSS VDD INVX1_LOC_376/Y
+ INVX1_LOC_377/Y NAND2X1_LOC
XNAND2X1_LOC_433 NAND2X1_LOC_433/a_36_24# NAND2X1_LOC_433/Y VSS VDD INVX1_LOC_74/Y
+ INVX1_LOC_137/Y NAND2X1_LOC
XNAND2X1_LOC_499 NAND2X1_LOC_499/a_36_24# INVX1_LOC_391/A VSS VDD NAND2X1_LOC_833/B
+ NAND2X1_LOC_496/Y NAND2X1_LOC
XNAND2X1_LOC_444 NAND2X1_LOC_444/a_36_24# INVX1_LOC_350/A VSS VDD NAND2X1_LOC_444/A
+ INVX1_LOC_349/Y NAND2X1_LOC
XNAND2X1_LOC_422 NAND2X1_LOC_422/a_36_24# NAND2X1_LOC_448/B VSS VDD INVX1_LOC_20/Y
+ INVX1_LOC_90/Y NAND2X1_LOC
XNAND2X1_LOC_455 NAND2X1_LOC_455/a_36_24# INVX1_LOC_361/A VSS VDD INVX1_LOC_77/Y INVX1_LOC_351/Y
+ NAND2X1_LOC
XNAND2X1_LOC_488 NAND2X1_LOC_488/a_36_24# NAND2X1_LOC_488/Y VSS VDD INVX1_LOC_145/Y
+ INVX1_LOC_199/Y NAND2X1_LOC
XNAND2X1_LOC_252 NAND2X1_LOC_252/a_36_24# NAND2X1_LOC_252/Y VSS VDD INVX1_LOC_62/Y
+ INVX1_LOC_63/Y NAND2X1_LOC
XNAND2X1_LOC_230 NAND2X1_LOC_230/a_36_24# NAND2X1_LOC_231/B VSS VDD INVX1_LOC_11/Y
+ INVX1_LOC_41/Y NAND2X1_LOC
XNAND2X1_LOC_241 NAND2X1_LOC_241/a_36_24# INVX1_LOC_208/A VSS VDD NAND2X1_LOC_237/Y
+ NAND2X1_LOC_241/B NAND2X1_LOC
XNAND2X1_LOC_274 NAND2X1_LOC_274/a_36_24# NAND2X1_LOC_274/Y VSS VDD NAND2X1_LOC_541/B
+ NAND2X1_LOC_274/B NAND2X1_LOC
XNAND2X1_LOC_285 NAND2X1_LOC_285/a_36_24# INVX1_LOC_239/A VSS VDD NAND2X1_LOC_285/A
+ NAND2X1_LOC_285/B NAND2X1_LOC
XNAND2X1_LOC_296 NAND2X1_LOC_296/a_36_24# NAND2X1_LOC_296/Y VSS VDD INVX1_LOC_246/Y
+ INVX1_LOC_247/Y NAND2X1_LOC
XNAND2X1_LOC_263 NAND2X1_LOC_263/a_36_24# INVX1_LOC_223/A VSS VDD INVX1_LOC_31/Y INVX1_LOC_46/Y
+ NAND2X1_LOC
XINVX1_LOC_107 INVX1_LOC_107/Y VSS VDD INVX1_LOC_107/A INVX1_LOC
XINVX1_LOC_118 INVX1_LOC_118/Y VSS VDD INVX1_LOC_118/A INVX1_LOC
XINVX1_LOC_129 INVX1_LOC_395/A VSS VDD INVX1_LOC_129/A INVX1_LOC
XINVX1_LOC_663 INVX1_LOC_663/Y VSS VDD INVX1_LOC_663/A INVX1_LOC
XINVX1_LOC_652 INVX1_LOC_652/Y VSS VDD INVX1_LOC_652/A INVX1_LOC
XINVX1_LOC_630 INVX1_LOC_630/Y VSS VDD INVX1_LOC_630/A INVX1_LOC
XINVX1_LOC_685 INVX1_LOC_685/Y VSS VDD INVX1_LOC_685/A INVX1_LOC
XINVX1_LOC_641 INVX1_LOC_641/Y VSS VDD INVX1_LOC_641/A INVX1_LOC
XINVX1_LOC_674 INVX1_LOC_674/Y VSS VDD INVX1_LOC_674/A INVX1_LOC
XNAND2X1_LOC_829 NAND2X1_LOC_829/a_36_24# NAND2X1_LOC_829/Y VSS VDD INVX1_LOC_69/Y
+ NAND2X1_LOC_829/B NAND2X1_LOC
XNAND2X1_LOC_818 NAND2X1_LOC_818/a_36_24# NAND2X1_LOC_820/A VSS VDD INVX1_LOC_647/Y
+ INVX1_LOC_648/Y NAND2X1_LOC
XNAND2X1_LOC_807 NAND2X1_LOC_807/a_36_24# INVX1_LOC_637/A VSS VDD INVX1_LOC_635/Y
+ INVX1_LOC_636/Y NAND2X1_LOC
XINVX1_LOC_493 INVX1_LOC_493/Y VSS VDD INVX1_LOC_493/A INVX1_LOC
XINVX1_LOC_471 INVX1_LOC_471/Y VSS VDD INVX1_LOC_114/A INVX1_LOC
XINVX1_LOC_460 INVX1_LOC_460/Y VSS VDD INVX1_LOC_460/A INVX1_LOC
XINVX1_LOC_482 INVX1_LOC_482/Y VSS VDD INVX1_LOC_482/A INVX1_LOC
XINVX1_LOC_27 INVX1_LOC_27/Y VSS VDD INVX1_LOC_27/A INVX1_LOC
XNAND2X1_LOC_648 NAND2X1_LOC_648/a_36_24# INVX1_LOC_509/A VSS VDD INVX1_LOC_504/Y
+ INVX1_LOC_506/Y NAND2X1_LOC
XNAND2X1_LOC_659 NAND2X1_LOC_659/a_36_24# INVX1_LOC_520/A VSS VDD INVX1_LOC_518/Y
+ INVX1_LOC_519/Y NAND2X1_LOC
XNAND2X1_LOC_637 NAND2X1_LOC_637/a_36_24# INVX1_LOC_497/A VSS VDD NAND2X1_LOC_637/A
+ NAND2X1_LOC_586/Y NAND2X1_LOC
XNAND2X1_LOC_604 NAND2X1_LOC_604/a_36_24# NAND2X1_LOC_605/B VSS VDD INVX1_LOC_74/Y
+ INVX1_LOC_586/A NAND2X1_LOC
XNAND2X1_LOC_615 NAND2X1_LOC_615/a_36_24# NAND2X1_LOC_615/Y VSS VDD INVX1_LOC_31/Y
+ NAND2X1_LOC_615/B NAND2X1_LOC
XNAND2X1_LOC_626 NAND2X1_LOC_626/a_36_24# NAND2X1_LOC_626/Y VSS VDD INVX1_LOC_93/Y
+ INVX1_LOC_586/A NAND2X1_LOC
XINVX1_LOC_16 INVX1_LOC_16/Y VSS VDD INPUT_1 INVX1_LOC
XINVX1_LOC_290 INVX1_LOC_290/Y VSS VDD INVX1_LOC_290/A INVX1_LOC
XINVX1_LOC_49 INVX1_LOC_49/Y VSS VDD INVX1_LOC_49/A INVX1_LOC
XINVX1_LOC_38 INVX1_LOC_87/A VSS VDD INVX1_LOC_38/A INVX1_LOC
XNAND2X1_LOC_90 NAND2X1_LOC_90/a_36_24# INVX1_LOC_89/A VSS VDD INVX1_LOC_46/Y INVX1_LOC_92/A
+ NAND2X1_LOC
XNAND2X1_LOC_434 NAND2X1_LOC_434/a_36_24# INVX1_LOC_344/A VSS VDD NAND2X1_LOC_174/B
+ NAND2X1_LOC_434/B NAND2X1_LOC
XNAND2X1_LOC_423 NAND2X1_LOC_423/a_36_24# NAND2X1_LOC_832/A VSS VDD INVX1_LOC_11/Y
+ INVX1_LOC_69/Y NAND2X1_LOC
XNAND2X1_LOC_412 NAND2X1_LOC_412/a_36_24# INVX1_LOC_338/A VSS VDD INVX1_LOC_46/Y INVX1_LOC_50/Y
+ NAND2X1_LOC
XNAND2X1_LOC_445 NAND2X1_LOC_445/a_36_24# INVX1_LOC_351/A VSS VDD NAND2X1_LOC_237/Y
+ NAND2X1_LOC_318/A NAND2X1_LOC
XNAND2X1_LOC_401 NAND2X1_LOC_401/a_36_24# INVX1_LOC_325/A VSS VDD NAND2X1_LOC_395/Y
+ NAND2X1_LOC_396/Y NAND2X1_LOC
XNAND2X1_LOC_478 NAND2X1_LOC_478/a_36_24# INVX1_LOC_384/A VSS VDD INVX1_LOC_375/Y
+ INVX1_LOC_383/Y NAND2X1_LOC
XNAND2X1_LOC_456 NAND2X1_LOC_456/a_36_24# INVX1_LOC_362/A VSS VDD NAND2X1_LOC_184/Y
+ INVX1_LOC_217/Y NAND2X1_LOC
XNAND2X1_LOC_467 NAND2X1_LOC_467/a_36_24# INVX1_LOC_373/A VSS VDD NAND2X1_LOC_467/A
+ INVX1_LOC_358/Y NAND2X1_LOC
XNAND2X1_LOC_489 NAND2X1_LOC_489/a_36_24# INVX1_LOC_388/A VSS VDD NAND2X1_LOC_489/A
+ NAND2X1_LOC_488/Y NAND2X1_LOC
XNAND2X1_LOC_253 NAND2X1_LOC_253/a_36_24# NAND2X1_LOC_253/Y VSS VDD INVX1_LOC_69/Y
+ INVX1_LOC_479/A NAND2X1_LOC
XNAND2X1_LOC_220 NAND2X1_LOC_220/a_36_24# INVX1_LOC_196/A VSS VDD INVX1_LOC_188/Y
+ INVX1_LOC_189/Y NAND2X1_LOC
XNAND2X1_LOC_286 NAND2X1_LOC_286/a_36_24# INVX1_LOC_240/A VSS VDD NAND2X1_LOC_286/A
+ INVX1_LOC_239/Y NAND2X1_LOC
XNAND2X1_LOC_275 NAND2X1_LOC_275/a_36_24# NAND2X1_LOC_275/Y VSS VDD INVX1_LOC_234/Y
+ NAND2X1_LOC_274/Y NAND2X1_LOC
XNAND2X1_LOC_264 NAND2X1_LOC_264/a_36_24# INVX1_LOC_224/A VSS VDD INVX1_LOC_225/Y
+ INVX1_LOC_226/Y NAND2X1_LOC
XNAND2X1_LOC_231 NAND2X1_LOC_231/a_36_24# INVX1_LOC_203/A VSS VDD NAND2X1_LOC_231/A
+ NAND2X1_LOC_231/B NAND2X1_LOC
XNAND2X1_LOC_242 NAND2X1_LOC_242/a_36_24# INVX1_LOC_209/A VSS VDD NAND2X1_LOC_242/A
+ INVX1_LOC_208/Y NAND2X1_LOC
XNAND2X1_LOC_297 NAND2X1_LOC_297/a_36_24# NAND2X1_LOC_297/Y VSS VDD INVX1_LOC_50/Y
+ NAND2X1_LOC_296/Y NAND2X1_LOC
XINVX1_LOC_108 INVX1_LOC_108/Y VSS VDD INVX1_LOC_108/A INVX1_LOC
XINVX1_LOC_119 INVX1_LOC_119/Y VSS VDD INVX1_LOC_119/A INVX1_LOC
XINVX1_LOC_620 INVX1_LOC_620/Y VSS VDD INVX1_LOC_620/A INVX1_LOC
XINVX1_LOC_664 INVX1_LOC_664/Y VSS VDD INVX1_LOC_664/A INVX1_LOC
XINVX1_LOC_653 INVX1_LOC_653/Y VSS VDD INVX1_LOC_653/A INVX1_LOC
XINVX1_LOC_675 INVX1_LOC_675/Y VSS VDD INVX1_LOC_675/A INVX1_LOC
XINVX1_LOC_631 INVX1_LOC_631/Y VSS VDD INVX1_LOC_631/A INVX1_LOC
XINVX1_LOC_686 INVX1_LOC_686/Y VSS VDD INVX1_LOC_686/A INVX1_LOC
XINVX1_LOC_642 INVX1_LOC_642/Y VSS VDD INVX1_LOC_65/Y INVX1_LOC
XINVX1_LOC_461 INVX1_LOC_461/Y VSS VDD INVX1_LOC_50/Y INVX1_LOC
XINVX1_LOC_450 INVX1_LOC_450/Y VSS VDD INVX1_LOC_450/A INVX1_LOC
XNAND2X1_LOC_808 NAND2X1_LOC_808/a_36_24# INVX1_LOC_638/A VSS VDD INVX1_LOC_633/Y
+ INVX1_LOC_634/Y NAND2X1_LOC
XNAND2X1_LOC_819 NAND2X1_LOC_819/a_36_24# INVX1_LOC_649/A VSS VDD INVX1_LOC_53/Y INVX1_LOC_650/Y
+ NAND2X1_LOC
XINVX1_LOC_494 INVX1_LOC_494/Y VSS VDD INVX1_LOC_338/Y INVX1_LOC
XINVX1_LOC_472 INVX1_LOC_472/Y VSS VDD INVX1_LOC_79/A INVX1_LOC
XINVX1_LOC_483 INVX1_LOC_483/Y VSS VDD INVX1_LOC_483/A INVX1_LOC
XNAND2X1_LOC_605 NAND2X1_LOC_605/a_36_24# INVX1_LOC_469/A VSS VDD NAND2X1_LOC_603/Y
+ NAND2X1_LOC_605/B NAND2X1_LOC
XNAND2X1_LOC_627 NAND2X1_LOC_627/a_36_24# NAND2X1_LOC_627/Y VSS VDD INVX1_LOC_11/Y
+ INVX1_LOC_45/Y NAND2X1_LOC
XNAND2X1_LOC_616 NAND2X1_LOC_616/a_36_24# NAND2X1_LOC_616/Y VSS VDD INVX1_LOC_26/Y
+ INVX1_LOC_100/Y NAND2X1_LOC
XINVX1_LOC_280 INVX1_LOC_280/Y VSS VDD INVX1_LOC_280/A INVX1_LOC
XINVX1_LOC_291 INVX1_LOC_291/Y VSS VDD INVX1_LOC_291/A INVX1_LOC
XINVX1_LOC_28 INVX1_LOC_28/Y VSS VDD INVX1_LOC_7/Y INVX1_LOC
XNAND2X1_LOC_649 NAND2X1_LOC_649/a_36_24# INVX1_LOC_510/A VSS VDD INVX1_LOC_502/Y
+ INVX1_LOC_503/Y NAND2X1_LOC
XNAND2X1_LOC_638 NAND2X1_LOC_638/a_36_24# INVX1_LOC_498/A VSS VDD NAND2X1_LOC_638/A
+ INVX1_LOC_497/Y NAND2X1_LOC
XNAND2X1_LOC_91 NAND2X1_LOC_91/a_36_24# NAND2X1_LOC_97/B VSS VDD INVX1_LOC_58/Y INVX1_LOC_89/Y
+ NAND2X1_LOC
XNAND2X1_LOC_80 NAND2X1_LOC_80/a_36_24# INVX1_LOC_81/A VSS VDD INVX1_LOC_9/Y INVX1_LOC_82/Y
+ NAND2X1_LOC
XINVX1_LOC_17 INVX1_LOC_17/Y VSS VDD INVX1_LOC_17/A INVX1_LOC
XINVX1_LOC_39 INVX1_LOC_39/Y VSS VDD INVX1_LOC_84/A INVX1_LOC
XNAND2X1_LOC_468 NAND2X1_LOC_468/a_36_24# INVX1_LOC_374/A VSS VDD INVX1_LOC_346/Y
+ INVX1_LOC_348/Y NAND2X1_LOC
XNAND2X1_LOC_446 NAND2X1_LOC_446/a_36_24# INVX1_LOC_352/A VSS VDD NAND2X1_LOC_704/B
+ NAND2X1_LOC_418/Y NAND2X1_LOC
XNAND2X1_LOC_435 NAND2X1_LOC_435/a_36_24# INVX1_LOC_345/A VSS VDD NAND2X1_LOC_432/Y
+ NAND2X1_LOC_433/Y NAND2X1_LOC
XNAND2X1_LOC_424 NAND2X1_LOC_424/a_36_24# NAND2X1_LOC_449/B VSS VDD INVX1_LOC_50/Y
+ INVX1_LOC_80/A NAND2X1_LOC
XNAND2X1_LOC_413 NAND2X1_LOC_413/a_36_24# NAND2X1_LOC_413/Y VSS VDD INPUT_0 INVX1_LOC_338/Y
+ NAND2X1_LOC
XNAND2X1_LOC_457 NAND2X1_LOC_457/a_36_24# INVX1_LOC_363/A VSS VDD NAND2X1_LOC_457/A
+ INVX1_LOC_301/Y NAND2X1_LOC
XNAND2X1_LOC_402 NAND2X1_LOC_402/a_36_24# INVX1_LOC_326/A VSS VDD NAND2X1_LOC_397/Y
+ INVX1_LOC_325/Y NAND2X1_LOC
XNAND2X1_LOC_479 NAND2X1_LOC_479/a_36_24# INVX1_LOC_385/A VSS VDD INVX1_LOC_381/Y
+ INVX1_LOC_382/Y NAND2X1_LOC
XNAND2X1_LOC_254 NAND2X1_LOC_254/a_36_24# INVX1_LOC_217/A VSS VDD NAND2X1_LOC_252/Y
+ NAND2X1_LOC_253/Y NAND2X1_LOC
XNAND2X1_LOC_221 NAND2X1_LOC_221/a_36_24# INVX1_LOC_197/A VSS VDD INVX1_LOC_168/Y
+ INVX1_LOC_196/Y NAND2X1_LOC
XNAND2X1_LOC_210 NAND2X1_LOC_210/a_36_24# INVX1_LOC_186/A VSS VDD NAND2X1_LOC_210/A
+ NAND2X1_LOC_467/A NAND2X1_LOC
XNAND2X1_LOC_287 NAND2X1_LOC_287/a_36_24# INVX1_LOC_241/A VSS VDD NAND2X1_LOC_843/B
+ INVX1_LOC_238/Y NAND2X1_LOC
XNAND2X1_LOC_298 NAND2X1_LOC_298/a_36_24# NAND2X1_LOC_302/A VSS VDD INVX1_LOC_41/Y
+ INVX1_LOC_62/Y NAND2X1_LOC
XNAND2X1_LOC_276 NAND2X1_LOC_276/a_36_24# INVX1_LOC_235/A VSS VDD NAND2X1_LOC_276/A
+ NAND2X1_LOC_275/Y NAND2X1_LOC
XNAND2X1_LOC_265 NAND2X1_LOC_265/a_36_24# NAND2X1_LOC_267/A VSS VDD INVX1_LOC_48/Y
+ INVX1_LOC_227/Y NAND2X1_LOC
XNAND2X1_LOC_232 NAND2X1_LOC_232/a_36_24# NAND2X1_LOC_240/A VSS VDD INVX1_LOC_79/A
+ INVX1_LOC_145/Y NAND2X1_LOC
XNAND2X1_LOC_243 NAND2X1_LOC_243/a_36_24# INVX1_LOC_210/A VSS VDD NAND2X1_LOC_243/A
+ INVX1_LOC_207/Y NAND2X1_LOC
XINVX1_LOC_109 INVX1_LOC_109/Y VSS VDD INVX1_LOC_109/A INVX1_LOC
XINVX1_LOC_610 INVX1_LOC_610/Y VSS VDD INVX1_LOC_610/A INVX1_LOC
XINVX1_LOC_643 INVX1_LOC_643/Y VSS VDD INVX1_LOC_100/Y INVX1_LOC
XINVX1_LOC_654 INVX1_LOC_654/Y VSS VDD INVX1_LOC_654/A INVX1_LOC
XINVX1_LOC_632 INVX1_LOC_632/Y VSS VDD INVX1_LOC_632/A INVX1_LOC
XINVX1_LOC_621 INVX1_LOC_621/Y VSS VDD INVX1_LOC_621/A INVX1_LOC
XINVX1_LOC_676 INVX1_LOC_676/Y VSS VDD INVX1_LOC_676/A INVX1_LOC
XINVX1_LOC_665 INVX1_LOC_665/Y VSS VDD INVX1_LOC_665/A INVX1_LOC
XNAND2X1_LOC_809 NAND2X1_LOC_809/a_36_24# INVX1_LOC_639/A VSS VDD INVX1_LOC_631/Y
+ INVX1_LOC_632/Y NAND2X1_LOC
XINVX1_LOC_473 INVX1_LOC_473/Y VSS VDD INVX1_LOC_76/Y INVX1_LOC
XINVX1_LOC_495 INVX1_LOC_495/Y VSS VDD INVX1_LOC_495/A INVX1_LOC
XINVX1_LOC_462 INVX1_LOC_462/Y VSS VDD INVX1_LOC_261/Y INVX1_LOC
XINVX1_LOC_451 INVX1_LOC_451/Y VSS VDD INVX1_LOC_451/A INVX1_LOC
XINVX1_LOC_440 INVX1_LOC_440/Y VSS VDD INVX1_LOC_440/A INVX1_LOC
XINVX1_LOC_484 INVX1_LOC_484/Y VSS VDD INVX1_LOC_484/A INVX1_LOC
XNAND2X1_LOC_606 NAND2X1_LOC_606/a_36_24# NAND2X1_LOC_606/Y VSS VDD INVX1_LOC_470/Y
+ INVX1_LOC_471/Y NAND2X1_LOC
XNAND2X1_LOC_639 NAND2X1_LOC_639/a_36_24# INVX1_LOC_499/A VSS VDD INVX1_LOC_495/Y
+ INVX1_LOC_496/Y NAND2X1_LOC
XNAND2X1_LOC_628 NAND2X1_LOC_628/a_36_24# NAND2X1_LOC_628/Y VSS VDD INVX1_LOC_53/Y
+ INVX1_LOC_90/Y NAND2X1_LOC
XNAND2X1_LOC_617 NAND2X1_LOC_617/a_36_24# NAND2X1_LOC_621/B VSS VDD INVX1_LOC_47/Y
+ INVX1_LOC_58/Y NAND2X1_LOC
XINVX1_LOC_270 INVX1_LOC_270/Y VSS VDD INVX1_LOC_270/A INVX1_LOC
XINVX1_LOC_281 INVX1_LOC_281/Y VSS VDD INVX1_LOC_281/A INVX1_LOC
XINVX1_LOC_29 INVX1_LOC_29/Y VSS VDD INVX1_LOC_29/A INVX1_LOC
XINVX1_LOC_18 INVX1_LOC_18/Y VSS VDD INVX1_LOC_18/A INVX1_LOC
XINVX1_LOC_292 INVX1_LOC_292/Y VSS VDD INVX1_LOC_292/A INVX1_LOC
XNAND2X1_LOC_92 NAND2X1_LOC_92/a_36_24# INVX1_LOC_90/A VSS VDD INPUT_1 INVX1_LOC_12/Y
+ NAND2X1_LOC
XNAND2X1_LOC_70 NAND2X1_LOC_70/a_36_24# INVX1_LOC_74/A VSS VDD INVX1_LOC_3/Y INVX1_LOC_55/Y
+ NAND2X1_LOC
XNAND2X1_LOC_81 NAND2X1_LOC_81/a_36_24# NAND2X1_LOC_81/Y VSS VDD INVX1_LOC_63/Y INVX1_LOC_81/Y
+ NAND2X1_LOC
XNAND2X1_LOC_469 NAND2X1_LOC_469/a_36_24# INVX1_LOC_375/A VSS VDD INVX1_LOC_350/Y
+ INVX1_LOC_374/Y NAND2X1_LOC
XNAND2X1_LOC_436 NAND2X1_LOC_436/a_36_24# INVX1_LOC_346/A VSS VDD INVX1_LOC_344/Y
+ INVX1_LOC_345/Y NAND2X1_LOC
XNAND2X1_LOC_458 NAND2X1_LOC_458/a_36_24# INVX1_LOC_364/A VSS VDD NAND2X1_LOC_372/Y
+ INVX1_LOC_304/Y NAND2X1_LOC
XNAND2X1_LOC_414 NAND2X1_LOC_414/a_36_24# NAND2X1_LOC_415/B VSS VDD INPUT_3 INVX1_LOC_7/Y
+ NAND2X1_LOC
XNAND2X1_LOC_425 NAND2X1_LOC_425/a_36_24# INVX1_LOC_340/A VSS VDD INVX1_LOC_341/Y
+ INVX1_LOC_25/Y NAND2X1_LOC
XNAND2X1_LOC_447 NAND2X1_LOC_447/a_36_24# INVX1_LOC_353/A VSS VDD NAND2X1_LOC_506/B
+ NAND2X1_LOC_420/Y NAND2X1_LOC
XNAND2X1_LOC_403 NAND2X1_LOC_403/a_36_24# INVX1_LOC_327/A VSS VDD NAND2X1_LOC_403/A
+ INVX1_LOC_324/Y NAND2X1_LOC
XNAND2X1_LOC_211 NAND2X1_LOC_211/a_36_24# INVX1_LOC_187/A VSS VDD INVX1_LOC_155/Y
+ INVX1_LOC_157/Y NAND2X1_LOC
XNAND2X1_LOC_200 NAND2X1_LOC_200/a_36_24# INVX1_LOC_176/A VSS VDD INVX1_LOC_169/Y
+ INVX1_LOC_170/Y NAND2X1_LOC
XNAND2X1_LOC_299 NAND2X1_LOC_299/a_36_24# NAND2X1_LOC_299/Y VSS VDD INVX1_LOC_20/Y
+ INVX1_LOC_114/A NAND2X1_LOC
XNAND2X1_LOC_255 NAND2X1_LOC_255/a_36_24# INVX1_LOC_218/A VSS VDD INVX1_LOC_46/Y INVX1_LOC_145/Y
+ NAND2X1_LOC
XNAND2X1_LOC_288 NAND2X1_LOC_288/a_36_24# INVX1_LOC_242/A VSS VDD INVX1_LOC_240/Y
+ INVX1_LOC_241/Y NAND2X1_LOC
XNAND2X1_LOC_277 NAND2X1_LOC_277/a_36_24# INVX1_LOC_236/A VSS VDD INVX1_LOC_46/Y INVX1_LOC_53/Y
+ NAND2X1_LOC
XNAND2X1_LOC_233 NAND2X1_LOC_233/a_36_24# INVX1_LOC_204/A VSS VDD INPUT_0 INVX1_LOC_21/Y
+ NAND2X1_LOC
XNAND2X1_LOC_244 NAND2X1_LOC_244/a_36_24# INVX1_LOC_211/A VSS VDD INVX1_LOC_209/Y
+ INVX1_LOC_210/Y NAND2X1_LOC
XNAND2X1_LOC_266 NAND2X1_LOC_266/a_36_24# INVX1_LOC_228/A VSS VDD NAND2X1_LOC_786/B
+ INVX1_LOC_229/Y NAND2X1_LOC
XNAND2X1_LOC_222 NAND2X1_LOC_222/a_36_24# INVX1_LOC_198/A VSS VDD INVX1_LOC_194/Y
+ INVX1_LOC_195/Y NAND2X1_LOC
XINVX1_LOC_611 INVX1_LOC_611/Y VSS VDD INVX1_LOC_611/A INVX1_LOC
XINVX1_LOC_644 INVX1_LOC_644/Y VSS VDD INVX1_LOC_199/Y INVX1_LOC
XINVX1_LOC_633 INVX1_LOC_633/Y VSS VDD INVX1_LOC_633/A INVX1_LOC
XINVX1_LOC_655 INVX1_LOC_655/Y VSS VDD INVX1_LOC_655/A INVX1_LOC
XINVX1_LOC_677 INVX1_LOC_677/Y VSS VDD INVX1_LOC_677/A INVX1_LOC
XINVX1_LOC_666 INVX1_LOC_666/Y VSS VDD INVX1_LOC_666/A INVX1_LOC
XINVX1_LOC_622 INVX1_LOC_622/Y VSS VDD INVX1_LOC_622/A INVX1_LOC
XINVX1_LOC_600 INVX1_LOC_600/Y VSS VDD INVX1_LOC_600/A INVX1_LOC
XINVX1_LOC_452 INVX1_LOC_452/Y VSS VDD INVX1_LOC_452/A INVX1_LOC
XINVX1_LOC_474 INVX1_LOC_474/Y VSS VDD INVX1_LOC_48/Y INVX1_LOC
XINVX1_LOC_496 INVX1_LOC_496/Y VSS VDD INVX1_LOC_496/A INVX1_LOC
XINVX1_LOC_463 INVX1_LOC_463/Y VSS VDD INVX1_LOC_463/A INVX1_LOC
XINVX1_LOC_430 INVX1_LOC_430/Y VSS VDD INVX1_LOC_430/A INVX1_LOC
XINVX1_LOC_441 INVX1_LOC_441/Y VSS VDD INVX1_LOC_441/A INVX1_LOC
XINVX1_LOC_485 INVX1_LOC_485/Y VSS VDD INVX1_LOC_485/A INVX1_LOC
XNAND2X1_LOC_607 NAND2X1_LOC_607/a_36_24# NAND2X1_LOC_646/A VSS VDD INVX1_LOC_26/Y
+ NAND2X1_LOC_606/Y NAND2X1_LOC
XNAND2X1_LOC_618 NAND2X1_LOC_618/a_36_24# INVX1_LOC_480/A VSS VDD INVX1_LOC_481/Y
+ INVX1_LOC_84/A NAND2X1_LOC
XNAND2X1_LOC_629 NAND2X1_LOC_629/a_36_24# INVX1_LOC_487/A VSS VDD NAND2X1_LOC_626/Y
+ NAND2X1_LOC_627/Y NAND2X1_LOC
XINVX1_LOC_282 INVX1_LOC_282/Y VSS VDD INVX1_LOC_282/A INVX1_LOC
XINVX1_LOC_293 INVX1_LOC_293/Y VSS VDD INVX1_LOC_293/A INVX1_LOC
XINVX1_LOC_260 INVX1_LOC_260/Y VSS VDD INVX1_LOC_68/Y INVX1_LOC
XINVX1_LOC_271 INVX1_LOC_271/Y VSS VDD INVX1_LOC_271/A INVX1_LOC
XINVX1_LOC_19 INVX1_LOC_19/Y VSS VDD INPUT_4 INVX1_LOC
XNAND2X1_LOC_71 NAND2X1_LOC_71/a_36_24# INVX1_LOC_75/A VSS VDD INVX1_LOC_9/Y INVX1_LOC_65/Y
+ NAND2X1_LOC
XNAND2X1_LOC_93 NAND2X1_LOC_93/a_36_24# NAND2X1_LOC_93/Y VSS VDD INVX1_LOC_35/Y INVX1_LOC_90/Y
+ NAND2X1_LOC
XNAND2X1_LOC_60 NAND2X1_LOC_60/a_36_24# NAND2X1_LOC_60/Y VSS VDD INVX1_LOC_47/Y INVX1_LOC_63/Y
+ NAND2X1_LOC
XNAND2X1_LOC_82 NAND2X1_LOC_82/a_36_24# INVX1_LOC_83/A VSS VDD INVX1_LOC_21/Y INVX1_LOC_84/Y
+ NAND2X1_LOC
XNAND2X1_LOC_437 NAND2X1_LOC_437/a_36_24# NAND2X1_LOC_440/A VSS VDD INVX1_LOC_63/Y
+ INVX1_LOC_134/Y NAND2X1_LOC
XNAND2X1_LOC_426 NAND2X1_LOC_426/a_36_24# NAND2X1_LOC_426/Y VSS VDD INVX1_LOC_114/A
+ INVX1_LOC_340/Y NAND2X1_LOC
XNAND2X1_LOC_448 NAND2X1_LOC_448/a_36_24# INVX1_LOC_354/A VSS VDD NAND2X1_LOC_448/A
+ NAND2X1_LOC_448/B NAND2X1_LOC
XNAND2X1_LOC_415 NAND2X1_LOC_415/a_36_24# NAND2X1_LOC_416/B VSS VDD INVX1_LOC_339/Y
+ NAND2X1_LOC_415/B NAND2X1_LOC
XNAND2X1_LOC_459 NAND2X1_LOC_459/a_36_24# INVX1_LOC_365/A VSS VDD NAND2X1_LOC_376/Y
+ NAND2X1_LOC_378/Y NAND2X1_LOC
XNAND2X1_LOC_404 NAND2X1_LOC_404/a_36_24# INVX1_LOC_328/A VSS VDD INVX1_LOC_326/Y
+ INVX1_LOC_327/Y NAND2X1_LOC
XNAND2X1_LOC_212 NAND2X1_LOC_212/a_36_24# INVX1_LOC_188/A VSS VDD INVX1_LOC_160/Y
+ INVX1_LOC_187/Y NAND2X1_LOC
XNAND2X1_LOC_234 NAND2X1_LOC_234/a_36_24# NAND2X1_LOC_234/Y VSS VDD INVX1_LOC_53/Y
+ INVX1_LOC_204/Y NAND2X1_LOC
XNAND2X1_LOC_201 NAND2X1_LOC_201/a_36_24# INVX1_LOC_177/A VSS VDD INVX1_LOC_64/Y NAND2X1_LOC_65/Y
+ NAND2X1_LOC
XNAND2X1_LOC_223 NAND2X1_LOC_223/a_36_24# GATE_222 VSS VDD INVX1_LOC_197/Y INVX1_LOC_198/Y
+ NAND2X1_LOC
XNAND2X1_LOC_256 NAND2X1_LOC_256/a_36_24# NAND2X1_LOC_344/B VSS VDD INVX1_LOC_219/Y
+ INVX1_LOC_218/Y NAND2X1_LOC
XNAND2X1_LOC_278 NAND2X1_LOC_278/a_36_24# NAND2X1_LOC_843/B VSS VDD INVX1_LOC_237/Y
+ INVX1_LOC_492/A NAND2X1_LOC
XNAND2X1_LOC_245 NAND2X1_LOC_245/a_36_24# INVX1_LOC_212/A VSS VDD INVX1_LOC_35/Y INVX1_LOC_46/Y
+ NAND2X1_LOC
XNAND2X1_LOC_267 NAND2X1_LOC_267/a_36_24# INVX1_LOC_230/A VSS VDD NAND2X1_LOC_267/A
+ INVX1_LOC_228/Y NAND2X1_LOC
XNAND2X1_LOC_289 NAND2X1_LOC_289/a_36_24# NAND2X1_LOC_333/B VSS VDD INVX1_LOC_58/Y
+ INVX1_LOC_199/Y NAND2X1_LOC
XNAND2X1_LOC_790 NAND2X1_LOC_790/a_36_24# INVX1_LOC_620/A VSS VDD NAND2X1_LOC_753/Y
+ NAND2X1_LOC_790/B NAND2X1_LOC
XINVX1_LOC_1 INVX1_LOC_1/Y VSS VDD INVX1_LOC_1/A INVX1_LOC
XINVX1_LOC_612 INVX1_LOC_612/Y VSS VDD INVX1_LOC_612/A INVX1_LOC
XINVX1_LOC_667 INVX1_LOC_667/Y VSS VDD INVX1_LOC_667/A INVX1_LOC
XINVX1_LOC_645 INVX1_LOC_645/Y VSS VDD INVX1_LOC_588/A INVX1_LOC
XINVX1_LOC_634 INVX1_LOC_634/Y VSS VDD INVX1_LOC_634/A INVX1_LOC
XINVX1_LOC_678 INVX1_LOC_678/Y VSS VDD INVX1_LOC_678/A INVX1_LOC
XINVX1_LOC_656 INVX1_LOC_656/Y VSS VDD INVX1_LOC_656/A INVX1_LOC
XINVX1_LOC_623 INVX1_LOC_623/Y VSS VDD INVX1_LOC_623/A INVX1_LOC
XINVX1_LOC_601 INVX1_LOC_601/Y VSS VDD INVX1_LOC_601/A INVX1_LOC
XINVX1_LOC_420 INVX1_LOC_420/Y VSS VDD INVX1_LOC_420/A INVX1_LOC
XINVX1_LOC_475 INVX1_LOC_475/Y VSS VDD INVX1_LOC_53/Y INVX1_LOC
XINVX1_LOC_464 INVX1_LOC_464/Y VSS VDD INVX1_LOC_51/Y INVX1_LOC
XINVX1_LOC_442 INVX1_LOC_442/Y VSS VDD INVX1_LOC_442/A INVX1_LOC
XINVX1_LOC_453 INVX1_LOC_453/Y VSS VDD INVX1_LOC_453/A INVX1_LOC
XINVX1_LOC_497 INVX1_LOC_497/Y VSS VDD INVX1_LOC_497/A INVX1_LOC
XINVX1_LOC_431 INVX1_LOC_431/Y VSS VDD INVX1_LOC_431/A INVX1_LOC
XINVX1_LOC_486 INVX1_LOC_486/Y VSS VDD INVX1_LOC_486/A INVX1_LOC
XINVX1_LOC_250 INVX1_LOC_250/Y VSS VDD INVX1_LOC_250/A INVX1_LOC
XINVX1_LOC_261 INVX1_LOC_261/Y VSS VDD INVX1_LOC_261/A INVX1_LOC
XNAND2X1_LOC_608 NAND2X1_LOC_608/a_36_24# NAND2X1_LOC_609/B VSS VDD INVX1_LOC_472/Y
+ INVX1_LOC_473/Y NAND2X1_LOC
XNAND2X1_LOC_619 NAND2X1_LOC_619/a_36_24# NAND2X1_LOC_619/Y VSS VDD INVX1_LOC_45/Y
+ INVX1_LOC_480/Y NAND2X1_LOC
XNAND2X1_LOC_61 NAND2X1_LOC_61/a_36_24# INVX1_LOC_64/A VSS VDD NAND2X1_LOC_61/A NAND2X1_LOC_60/Y
+ NAND2X1_LOC
XNAND2X1_LOC_50 NAND2X1_LOC_50/a_36_24# INVX1_LOC_55/A VSS VDD INVX1_LOC_56/Y INVX1_LOC_57/Y
+ NAND2X1_LOC
XINVX1_LOC_283 INVX1_LOC_283/Y VSS VDD INVX1_LOC_283/A INVX1_LOC
XINVX1_LOC_294 INVX1_LOC_294/Y VSS VDD INVX1_LOC_294/A INVX1_LOC
XINVX1_LOC_272 INVX1_LOC_272/Y VSS VDD INVX1_LOC_272/A INVX1_LOC
XNAND2X1_LOC_94 NAND2X1_LOC_94/a_36_24# INVX1_LOC_91/A VSS VDD INVX1_LOC_21/Y INVX1_LOC_92/Y
+ NAND2X1_LOC
XNAND2X1_LOC_72 NAND2X1_LOC_72/a_36_24# NAND2X1_LOC_72/Y VSS VDD INVX1_LOC_74/Y INVX1_LOC_75/Y
+ NAND2X1_LOC
XNAND2X1_LOC_83 NAND2X1_LOC_83/a_36_24# NAND2X1_LOC_84/B VSS VDD INVX1_LOC_35/Y INVX1_LOC_83/Y
+ NAND2X1_LOC
XNAND2X1_LOC_427 NAND2X1_LOC_427/a_36_24# NAND2X1_LOC_427/Y VSS VDD INVX1_LOC_74/Y
+ INVX1_LOC_479/A NAND2X1_LOC
XNAND2X1_LOC_405 NAND2X1_LOC_405/a_36_24# NAND2X1_LOC_406/B VSS VDD INVX1_LOC_329/Y
+ INVX1_LOC_259/Y NAND2X1_LOC
XNAND2X1_LOC_416 NAND2X1_LOC_416/a_36_24# NAND2X1_LOC_416/Y VSS VDD INVX1_LOC_145/Y
+ NAND2X1_LOC_416/B NAND2X1_LOC
XNAND2X1_LOC_438 NAND2X1_LOC_438/a_36_24# NAND2X1_LOC_544/B VSS VDD INVX1_LOC_32/Y
+ INVX1_LOC_74/Y NAND2X1_LOC
XNAND2X1_LOC_449 NAND2X1_LOC_449/a_36_24# INVX1_LOC_355/A VSS VDD NAND2X1_LOC_832/A
+ NAND2X1_LOC_449/B NAND2X1_LOC
XNAND2X1_LOC_257 NAND2X1_LOC_257/a_36_24# NAND2X1_LOC_259/A VSS VDD INVX1_LOC_26/Y
+ INVX1_LOC_479/A NAND2X1_LOC
XNAND2X1_LOC_213 NAND2X1_LOC_213/a_36_24# INVX1_LOC_189/A VSS VDD INVX1_LOC_185/Y
+ INVX1_LOC_186/Y NAND2X1_LOC
XNAND2X1_LOC_246 NAND2X1_LOC_246/a_36_24# NAND2X1_LOC_342/A VSS VDD INVX1_LOC_66/A
+ INVX1_LOC_212/Y NAND2X1_LOC
XNAND2X1_LOC_268 NAND2X1_LOC_268/a_36_24# NAND2X1_LOC_269/B VSS VDD INVX1_LOC_45/Y
+ INVX1_LOC_90/Y NAND2X1_LOC
XNAND2X1_LOC_224 NAND2X1_LOC_224/a_36_24# NAND2X1_LOC_227/A VSS VDD INVX1_LOC_41/Y
+ INVX1_LOC_117/Y NAND2X1_LOC
XNAND2X1_LOC_202 NAND2X1_LOC_202/a_36_24# INVX1_LOC_178/A VSS VDD NAND2X1_LOC_67/Y
+ NAND2X1_LOC_69/Y NAND2X1_LOC
XNAND2X1_LOC_235 NAND2X1_LOC_235/a_36_24# NAND2X1_LOC_243/A VSS VDD INVX1_LOC_205/Y
+ INVX1_LOC_86/Y NAND2X1_LOC
XNAND2X1_LOC_279 NAND2X1_LOC_279/a_36_24# NAND2X1_LOC_284/A VSS VDD INVX1_LOC_50/Y
+ INVX1_LOC_479/A NAND2X1_LOC
XNAND2X1_LOC_780 NAND2X1_LOC_780/a_36_24# INVX1_LOC_610/A VSS VDD NAND2X1_LOC_780/A
+ NAND2X1_LOC_780/B NAND2X1_LOC
XNAND2X1_LOC_791 NAND2X1_LOC_791/a_36_24# INVX1_LOC_621/A VSS VDD NAND2X1_LOC_791/A
+ NAND2X1_LOC_791/B NAND2X1_LOC
XINVX1_LOC_602 INVX1_LOC_602/Y VSS VDD INVX1_LOC_602/A INVX1_LOC
XINVX1_LOC_2 INVX1_LOC_2/Y VSS VDD INPUT_6 INVX1_LOC
XINVX1_LOC_613 INVX1_LOC_613/Y VSS VDD INVX1_LOC_613/A INVX1_LOC
XINVX1_LOC_668 INVX1_LOC_668/Y VSS VDD INVX1_LOC_668/A INVX1_LOC
XINVX1_LOC_646 INVX1_LOC_646/Y VSS VDD INPUT_1 INVX1_LOC
XINVX1_LOC_679 INVX1_LOC_679/Y VSS VDD INVX1_LOC_679/A INVX1_LOC
XINVX1_LOC_624 INVX1_LOC_624/Y VSS VDD INVX1_LOC_624/A INVX1_LOC
XINVX1_LOC_657 INVX1_LOC_657/Y VSS VDD INVX1_LOC_657/A INVX1_LOC
XINVX1_LOC_635 INVX1_LOC_635/Y VSS VDD INVX1_LOC_635/A INVX1_LOC
XINVX1_LOC_443 INVX1_LOC_443/Y VSS VDD INVX1_LOC_443/A INVX1_LOC
XINVX1_LOC_421 INVX1_LOC_421/Y VSS VDD INVX1_LOC_421/A INVX1_LOC
XINVX1_LOC_432 INVX1_LOC_432/Y VSS VDD INVX1_LOC_432/A INVX1_LOC
XINVX1_LOC_410 INVX1_LOC_410/Y VSS VDD INVX1_LOC_410/A INVX1_LOC
XINVX1_LOC_476 INVX1_LOC_476/Y VSS VDD INVX1_LOC_476/A INVX1_LOC
XINVX1_LOC_498 INVX1_LOC_498/Y VSS VDD INVX1_LOC_498/A INVX1_LOC
XINVX1_LOC_465 INVX1_LOC_465/Y VSS VDD INVX1_LOC_245/A INVX1_LOC
XINVX1_LOC_454 INVX1_LOC_454/Y VSS VDD INVX1_LOC_454/A INVX1_LOC
XINVX1_LOC_487 INVX1_LOC_487/Y VSS VDD INVX1_LOC_487/A INVX1_LOC
XNAND2X1_LOC_609 NAND2X1_LOC_609/a_36_24# NAND2X1_LOC_646/B VSS VDD INVX1_LOC_63/Y
+ NAND2X1_LOC_609/B NAND2X1_LOC
XINVX1_LOC_240 INVX1_LOC_240/Y VSS VDD INVX1_LOC_240/A INVX1_LOC
XINVX1_LOC_251 INVX1_LOC_251/Y VSS VDD INVX1_LOC_251/A INVX1_LOC
XINVX1_LOC_295 INVX1_LOC_295/Y VSS VDD INVX1_LOC_295/A INVX1_LOC
XINVX1_LOC_262 INVX1_LOC_262/Y VSS VDD INPUT_4 INVX1_LOC
XINVX1_LOC_284 INVX1_LOC_284/Y VSS VDD INVX1_LOC_284/A INVX1_LOC
XINVX1_LOC_273 INVX1_LOC_273/Y VSS VDD INVX1_LOC_273/A INVX1_LOC
XNAND2X1_LOC_62 NAND2X1_LOC_62/a_36_24# INVX1_LOC_65/A VSS VDD INVX1_LOC_66/Y INVX1_LOC_67/Y
+ NAND2X1_LOC
XNAND2X1_LOC_73 NAND2X1_LOC_73/a_36_24# INVX1_LOC_76/A VSS VDD INVX1_LOC_66/A INVX1_LOC_46/Y
+ NAND2X1_LOC
XNAND2X1_LOC_51 NAND2X1_LOC_51/a_36_24# INVX1_LOC_58/A VSS VDD INVX1_LOC_40/Y INVX1_LOC_55/Y
+ NAND2X1_LOC
XNAND2X1_LOC_95 NAND2X1_LOC_95/a_36_24# INVX1_LOC_93/A VSS VDD INVX1_LOC_18/Y INVX1_LOC_55/Y
+ NAND2X1_LOC
XNAND2X1_LOC_40 NAND2X1_LOC_40/a_36_24# INVX1_LOC_48/A VSS VDD INVX1_LOC_3/Y INVX1_LOC_33/Y
+ NAND2X1_LOC
XNAND2X1_LOC_84 NAND2X1_LOC_84/a_36_24# INVX1_LOC_85/A VSS VDD NAND2X1_LOC_81/Y NAND2X1_LOC_84/B
+ NAND2X1_LOC
XNAND2X1_LOC_439 NAND2X1_LOC_439/a_36_24# INVX1_LOC_347/A VSS VDD NAND2X1_LOC_180/B
+ NAND2X1_LOC_544/B NAND2X1_LOC
XNAND2X1_LOC_428 NAND2X1_LOC_428/a_36_24# NAND2X1_LOC_428/Y VSS VDD INVX1_LOC_41/Y
+ INVX1_LOC_206/Y NAND2X1_LOC
XNAND2X1_LOC_417 NAND2X1_LOC_417/a_36_24# NAND2X1_LOC_704/B VSS VDD INVX1_LOC_53/Y
+ INVX1_LOC_199/Y NAND2X1_LOC
XNAND2X1_LOC_406 NAND2X1_LOC_406/a_36_24# NAND2X1_LOC_475/A VSS VDD INVX1_LOC_93/Y
+ NAND2X1_LOC_406/B NAND2X1_LOC
XNAND2X1_LOC_225 NAND2X1_LOC_225/a_36_24# INVX1_LOC_199/A VSS VDD INVX1_LOC_200/Y
+ INVX1_LOC_9/Y NAND2X1_LOC
XNAND2X1_LOC_258 NAND2X1_LOC_258/a_36_24# NAND2X1_LOC_258/Y VSS VDD INVX1_LOC_80/A
+ INVX1_LOC_145/Y NAND2X1_LOC
XNAND2X1_LOC_247 NAND2X1_LOC_247/a_36_24# NAND2X1_LOC_248/B VSS VDD INVX1_LOC_213/Y
+ INVX1_LOC_214/Y NAND2X1_LOC
XNAND2X1_LOC_269 NAND2X1_LOC_269/a_36_24# NAND2X1_LOC_271/A VSS VDD INVX1_LOC_231/Y
+ NAND2X1_LOC_269/B NAND2X1_LOC
XNAND2X1_LOC_203 NAND2X1_LOC_203/a_36_24# INVX1_LOC_179/A VSS VDD NAND2X1_LOC_72/Y
+ INVX1_LOC_77/Y NAND2X1_LOC
XNAND2X1_LOC_236 NAND2X1_LOC_236/a_36_24# INVX1_LOC_206/A VSS VDD INVX1_LOC_9/Y INVX1_LOC_84/A
+ NAND2X1_LOC
XNAND2X1_LOC_214 NAND2X1_LOC_214/a_36_24# INVX1_LOC_190/A VSS VDD INVX1_LOC_183/Y
+ INVX1_LOC_184/Y NAND2X1_LOC
XNAND2X1_LOC_781 NAND2X1_LOC_781/a_36_24# INVX1_LOC_611/A VSS VDD NAND2X1_LOC_781/A
+ NAND2X1_LOC_781/B NAND2X1_LOC
XNAND2X1_LOC_770 NAND2X1_LOC_770/a_36_24# INVX1_LOC_598/A VSS VDD NAND2X1_LOC_770/A
+ NAND2X1_LOC_770/B NAND2X1_LOC
XNAND2X1_LOC_792 NAND2X1_LOC_792/a_36_24# INVX1_LOC_622/A VSS VDD NAND2X1_LOC_759/Y
+ INVX1_LOC_621/Y NAND2X1_LOC
XINVX1_LOC_614 INVX1_LOC_614/Y VSS VDD INVX1_LOC_614/A INVX1_LOC
XINVX1_LOC_625 INVX1_LOC_625/Y VSS VDD INVX1_LOC_625/A INVX1_LOC
XINVX1_LOC_636 INVX1_LOC_636/Y VSS VDD INVX1_LOC_636/A INVX1_LOC
XINVX1_LOC_603 INVX1_LOC_603/Y VSS VDD INVX1_LOC_603/A INVX1_LOC
XINVX1_LOC_3 INVX1_LOC_3/Y VSS VDD INVX1_LOC_3/A INVX1_LOC
XINVX1_LOC_647 INVX1_LOC_647/Y VSS VDD INVX1_LOC_9/Y INVX1_LOC
XINVX1_LOC_669 INVX1_LOC_669/Y VSS VDD INVX1_LOC_669/A INVX1_LOC
XINVX1_LOC_658 INVX1_LOC_658/Y VSS VDD INVX1_LOC_658/A INVX1_LOC
XINVX1_LOC_477 INVX1_LOC_477/Y VSS VDD INVX1_LOC_92/A INVX1_LOC
XINVX1_LOC_466 INVX1_LOC_505/A VSS VDD INVX1_LOC_466/A INVX1_LOC
XINVX1_LOC_444 INVX1_LOC_444/Y VSS VDD INVX1_LOC_444/A INVX1_LOC
XINVX1_LOC_433 INVX1_LOC_433/Y VSS VDD INVX1_LOC_433/A INVX1_LOC
XINVX1_LOC_411 INVX1_LOC_411/Y VSS VDD INVX1_LOC_411/A INVX1_LOC
XINVX1_LOC_400 INVX1_LOC_400/Y VSS VDD INVX1_LOC_400/A INVX1_LOC
XINVX1_LOC_422 INVX1_LOC_422/Y VSS VDD INVX1_LOC_422/A INVX1_LOC
XINVX1_LOC_455 INVX1_LOC_455/Y VSS VDD INVX1_LOC_455/A INVX1_LOC
XINVX1_LOC_499 INVX1_LOC_499/Y VSS VDD INVX1_LOC_499/A INVX1_LOC
XINVX1_LOC_488 INVX1_LOC_488/Y VSS VDD INVX1_LOC_488/A INVX1_LOC
XINVX1_LOC_241 INVX1_LOC_241/Y VSS VDD INVX1_LOC_241/A INVX1_LOC
XINVX1_LOC_252 INVX1_LOC_252/Y VSS VDD INVX1_LOC_252/A INVX1_LOC
XINVX1_LOC_263 INVX1_LOC_263/Y VSS VDD INVX1_LOC_259/Y INVX1_LOC
XINVX1_LOC_230 INVX1_LOC_230/Y VSS VDD INVX1_LOC_230/A INVX1_LOC
XINVX1_LOC_296 INVX1_LOC_296/Y VSS VDD INVX1_LOC_296/A INVX1_LOC
XINVX1_LOC_285 INVX1_LOC_285/Y VSS VDD INVX1_LOC_285/A INVX1_LOC
XINVX1_LOC_274 INVX1_LOC_274/Y VSS VDD INVX1_LOC_274/A INVX1_LOC
XNAND2X1_LOC_96 NAND2X1_LOC_96/a_36_24# NAND2X1_LOC_98/B VSS VDD INVX1_LOC_91/Y INVX1_LOC_93/Y
+ NAND2X1_LOC
XNAND2X1_LOC_74 NAND2X1_LOC_74/a_36_24# NAND2X1_LOC_76/A VSS VDD INVX1_LOC_41/Y INVX1_LOC_76/Y
+ NAND2X1_LOC
XNAND2X1_LOC_63 NAND2X1_LOC_63/a_36_24# INVX1_LOC_68/A VSS VDD INVX1_LOC_12/Y INVX1_LOC_65/Y
+ NAND2X1_LOC
XNAND2X1_LOC_52 NAND2X1_LOC_52/a_36_24# NAND2X1_LOC_52/Y VSS VDD INVX1_LOC_54/Y INVX1_LOC_58/Y
+ NAND2X1_LOC
XNAND2X1_LOC_41 NAND2X1_LOC_41/a_36_24# NAND2X1_LOC_41/Y VSS VDD INVX1_LOC_17/Y INVX1_LOC_48/Y
+ NAND2X1_LOC
XNAND2X1_LOC_30 NAND2X1_LOC_30/a_36_24# INVX1_LOC_40/A VSS VDD INPUT_4 INPUT_5
+ NAND2X1_LOC
XNAND2X1_LOC_85 NAND2X1_LOC_85/a_36_24# INVX1_LOC_86/A VSS VDD INVX1_LOC_26/Y INVX1_LOC_46/Y
+ NAND2X1_LOC
XNAND2X1_LOC_418 NAND2X1_LOC_418/a_36_24# NAND2X1_LOC_418/Y VSS VDD INVX1_LOC_79/A
+ INVX1_LOC_58/Y NAND2X1_LOC
XNAND2X1_LOC_407 NAND2X1_LOC_407/a_36_24# INVX1_LOC_330/A VSS VDD INVX1_LOC_331/Y
+ INVX1_LOC_332/Y NAND2X1_LOC
XNAND2X1_LOC_429 NAND2X1_LOC_429/a_36_24# INVX1_LOC_342/A VSS VDD INVX1_LOC_343/Y
+ INVX1_LOC_18/Y NAND2X1_LOC
XNAND2X1_LOC_259 NAND2X1_LOC_259/a_36_24# INVX1_LOC_220/A VSS VDD NAND2X1_LOC_259/A
+ NAND2X1_LOC_258/Y NAND2X1_LOC
XNAND2X1_LOC_248 NAND2X1_LOC_248/a_36_24# NAND2X1_LOC_342/B VSS VDD INVX1_LOC_53/Y
+ NAND2X1_LOC_248/B NAND2X1_LOC
XNAND2X1_LOC_237 NAND2X1_LOC_237/a_36_24# NAND2X1_LOC_237/Y VSS VDD INVX1_LOC_35/Y
+ INVX1_LOC_206/Y NAND2X1_LOC
XNAND2X1_LOC_226 NAND2X1_LOC_226/a_36_24# NAND2X1_LOC_226/Y VSS VDD INVX1_LOC_26/Y
+ INVX1_LOC_199/Y NAND2X1_LOC
XNAND2X1_LOC_204 NAND2X1_LOC_204/a_36_24# INVX1_LOC_180/A VSS VDD NAND2X1_LOC_79/Y
+ INVX1_LOC_85/Y NAND2X1_LOC
XNAND2X1_LOC_215 NAND2X1_LOC_215/a_36_24# INVX1_LOC_191/A VSS VDD INVX1_LOC_181/Y
+ INVX1_LOC_182/Y NAND2X1_LOC
XNAND2X1_LOC_760 NAND2X1_LOC_760/a_36_24# NAND2X1_LOC_800/B VSS VDD INVX1_LOC_69/Y
+ INVX1_LOC_593/Y NAND2X1_LOC
XNAND2X1_LOC_782 NAND2X1_LOC_782/a_36_24# INVX1_LOC_612/A VSS VDD NAND2X1_LOC_782/A
+ INVX1_LOC_611/Y NAND2X1_LOC
XNAND2X1_LOC_771 NAND2X1_LOC_771/a_36_24# INVX1_LOC_599/A VSS VDD INVX1_LOC_597/Y
+ INVX1_LOC_598/Y NAND2X1_LOC
XNAND2X1_LOC_793 NAND2X1_LOC_793/a_36_24# INVX1_LOC_623/A VSS VDD INVX1_LOC_619/Y
+ INVX1_LOC_620/Y NAND2X1_LOC
XINVX1_LOC_4 INVX1_LOC_4/Y VSS VDD INPUT_4 INVX1_LOC
XINVX1_LOC_626 INVX1_LOC_626/Y VSS VDD INVX1_LOC_626/A INVX1_LOC
XINVX1_LOC_648 INVX1_LOC_648/Y VSS VDD INVX1_LOC_395/A INVX1_LOC
XINVX1_LOC_637 INVX1_LOC_637/Y VSS VDD INVX1_LOC_637/A INVX1_LOC
XINVX1_LOC_659 INVX1_LOC_659/Y VSS VDD INVX1_LOC_659/A INVX1_LOC
XINVX1_LOC_604 INVX1_LOC_604/Y VSS VDD INVX1_LOC_604/A INVX1_LOC
XINVX1_LOC_615 INVX1_LOC_615/Y VSS VDD INVX1_LOC_615/A INVX1_LOC
XNAND2X1_LOC_590 NAND2X1_LOC_590/a_36_24# NAND2X1_LOC_591/B VSS VDD INVX1_LOC_457/Y
+ INVX1_LOC_458/Y NAND2X1_LOC
XINVX1_LOC_434 INVX1_LOC_434/Y VSS VDD INVX1_LOC_434/A INVX1_LOC
XINVX1_LOC_445 INVX1_LOC_445/Y VSS VDD INVX1_LOC_445/A INVX1_LOC
XINVX1_LOC_401 INVX1_LOC_401/Y VSS VDD INVX1_LOC_401/A INVX1_LOC
XINVX1_LOC_467 INVX1_LOC_467/Y VSS VDD INVX1_LOC_463/Y INVX1_LOC
XINVX1_LOC_412 INVX1_LOC_412/Y VSS VDD INVX1_LOC_412/A INVX1_LOC
XINVX1_LOC_489 INVX1_LOC_489/Y VSS VDD INVX1_LOC_489/A INVX1_LOC
XINVX1_LOC_478 INVX1_LOC_478/Y VSS VDD INVX1_LOC_80/A INVX1_LOC
XINVX1_LOC_423 INVX1_LOC_423/Y VSS VDD INVX1_LOC_423/A INVX1_LOC
XINVX1_LOC_456 INVX1_LOC_456/Y VSS VDD INPUT_7 INVX1_LOC
XINVX1_LOC_220 INVX1_LOC_220/Y VSS VDD INVX1_LOC_220/A INVX1_LOC
XINVX1_LOC_264 INVX1_LOC_264/Y VSS VDD INVX1_LOC_58/Y INVX1_LOC
XINVX1_LOC_253 INVX1_LOC_253/Y VSS VDD INVX1_LOC_253/A INVX1_LOC
XINVX1_LOC_242 INVX1_LOC_242/Y VSS VDD INVX1_LOC_242/A INVX1_LOC
XINVX1_LOC_231 INVX1_LOC_231/Y VSS VDD INVX1_LOC_206/Y INVX1_LOC
XINVX1_LOC_286 INVX1_LOC_286/Y VSS VDD INVX1_LOC_286/A INVX1_LOC
XINVX1_LOC_297 INVX1_LOC_297/Y VSS VDD INVX1_LOC_297/A INVX1_LOC
XINVX1_LOC_275 INVX1_LOC_275/Y VSS VDD INVX1_LOC_275/A INVX1_LOC
XNAND2X1_LOC_75 NAND2X1_LOC_75/a_36_24# NAND2X1_LOC_76/B VSS VDD INVX1_LOC_32/Y INVX1_LOC_63/Y
+ NAND2X1_LOC
XNAND2X1_LOC_42 NAND2X1_LOC_42/a_36_24# INVX1_LOC_49/A VSS VDD INPUT_1 INVX1_LOC_46/Y
+ NAND2X1_LOC
XNAND2X1_LOC_97 NAND2X1_LOC_97/a_36_24# INVX1_LOC_94/A VSS VDD NAND2X1_LOC_97/A NAND2X1_LOC_97/B
+ NAND2X1_LOC
XNAND2X1_LOC_53 NAND2X1_LOC_53/a_36_24# INVX1_LOC_59/A VSS VDD INVX1_LOC_60/Y INVX1_LOC_55/Y
+ NAND2X1_LOC
XNAND2X1_LOC_64 NAND2X1_LOC_64/a_36_24# INVX1_LOC_69/A VSS VDD INVX1_LOC_29/Y INVX1_LOC_55/Y
+ NAND2X1_LOC
XNAND2X1_LOC_31 NAND2X1_LOC_31/a_36_24# INVX1_LOC_41/A VSS VDD INVX1_LOC_1/Y INVX1_LOC_40/Y
+ NAND2X1_LOC
XNAND2X1_LOC_86 NAND2X1_LOC_86/a_36_24# NAND2X1_LOC_86/Y VSS VDD INPUT_0 INVX1_LOC_86/Y
+ NAND2X1_LOC
XNAND2X1_LOC_20 NAND2X1_LOC_20/a_36_24# NAND2X1_LOC_20/Y VSS VDD INVX1_LOC_26/Y INVX1_LOC_27/Y
+ NAND2X1_LOC
XNAND2X1_LOC_419 NAND2X1_LOC_419/a_36_24# NAND2X1_LOC_506/B VSS VDD INVX1_LOC_45/Y
+ INVX1_LOC_49/Y NAND2X1_LOC
XNAND2X1_LOC_408 NAND2X1_LOC_408/a_36_24# INVX1_LOC_333/A VSS VDD INVX1_LOC_334/Y
+ INVX1_LOC_29/Y NAND2X1_LOC
XNAND2X1_LOC_216 NAND2X1_LOC_216/a_36_24# INVX1_LOC_192/A VSS VDD INVX1_LOC_98/Y INVX1_LOC_109/Y
+ NAND2X1_LOC
XNAND2X1_LOC_205 NAND2X1_LOC_205/a_36_24# INVX1_LOC_181/A VSS VDD INVX1_LOC_179/Y
+ INVX1_LOC_180/Y NAND2X1_LOC
XNAND2X1_LOC_249 NAND2X1_LOC_249/a_36_24# NAND2X1_LOC_249/Y VSS VDD INVX1_LOC_215/Y
+ INVX1_LOC_216/Y NAND2X1_LOC
XNAND2X1_LOC_238 NAND2X1_LOC_238/a_36_24# NAND2X1_LOC_241/B VSS VDD INVX1_LOC_32/Y
+ INVX1_LOC_58/Y NAND2X1_LOC
XNAND2X1_LOC_227 NAND2X1_LOC_227/a_36_24# INVX1_LOC_201/A VSS VDD NAND2X1_LOC_227/A
+ NAND2X1_LOC_226/Y NAND2X1_LOC
XNAND2X1_LOC_761 NAND2X1_LOC_761/a_36_24# NAND2X1_LOC_801/A VSS VDD INVX1_LOC_594/Y
+ INVX1_LOC_505/A NAND2X1_LOC
XNAND2X1_LOC_772 NAND2X1_LOC_772/a_36_24# INVX1_LOC_600/A VSS VDD INVX1_LOC_388/Y
+ INVX1_LOC_596/Y NAND2X1_LOC
XNAND2X1_LOC_750 NAND2X1_LOC_750/a_36_24# NAND2X1_LOC_750/Y VSS VDD INVX1_LOC_586/Y
+ NAND2X1_LOC_749/Y NAND2X1_LOC
XNAND2X1_LOC_794 NAND2X1_LOC_794/a_36_24# INVX1_LOC_624/A VSS VDD INVX1_LOC_617/Y
+ INVX1_LOC_618/Y NAND2X1_LOC
XNAND2X1_LOC_783 NAND2X1_LOC_783/a_36_24# INVX1_LOC_613/A VSS VDD INVX1_LOC_609/Y
+ INVX1_LOC_610/Y NAND2X1_LOC
XINVX1_LOC_5 INVX1_LOC_5/Y VSS VDD INPUT_5 INVX1_LOC
XINVX1_LOC_627 INVX1_LOC_627/Y VSS VDD INVX1_LOC_627/A INVX1_LOC
XINVX1_LOC_649 INVX1_LOC_649/Y VSS VDD INVX1_LOC_649/A INVX1_LOC
XINVX1_LOC_605 INVX1_LOC_605/Y VSS VDD INVX1_LOC_605/A INVX1_LOC
XINVX1_LOC_638 INVX1_LOC_638/Y VSS VDD INVX1_LOC_638/A INVX1_LOC
XINVX1_LOC_616 INVX1_LOC_616/Y VSS VDD INVX1_LOC_616/A INVX1_LOC
C0 INVX1_LOC_103/Y INVX1_LOC_109/Y 0.03fF
C1 INVX1_LOC_41/Y INVX1_LOC_462/Y 0.31fF
C2 INVX1_LOC_523/A NAND2X1_LOC_662/a_36_24# 0.02fF
C3 INPUT_0 NAND2X1_LOC_690/a_36_24# 0.00fF
C4 NAND2X1_LOC_108/Y INVX1_LOC_101/Y 0.01fF
C5 VDD INVX1_LOC_342/Y 0.28fF
C6 INVX1_LOC_417/Y INVX1_LOC_410/Y 0.08fF
C7 NAND2X1_LOC_475/A INVX1_LOC_230/A 0.03fF
C8 INVX1_LOC_255/Y NAND2X1_LOC_603/Y 0.13fF
C9 INVX1_LOC_400/Y INVX1_LOC_99/A 0.03fF
C10 INVX1_LOC_206/Y INVX1_LOC_556/Y 0.03fF
C11 NAND2X1_LOC_669/Y INVX1_LOC_45/Y 0.01fF
C12 INVX1_LOC_449/A INVX1_LOC_45/Y 0.07fF
C13 INVX1_LOC_51/Y INVX1_LOC_134/Y 0.21fF
C14 INVX1_LOC_107/A INVX1_LOC_99/Y 0.02fF
C15 INVX1_LOC_119/A NAND2X1_LOC_129/a_36_24# 0.02fF
C16 NAND2X1_LOC_48/Y INVX1_LOC_51/Y 0.06fF
C17 INVX1_LOC_465/Y INVX1_LOC_47/Y 0.03fF
C18 NAND2X1_LOC_17/a_36_24# INVX1_LOC_1/A 0.00fF
C19 INVX1_LOC_603/Y NAND2X1_LOC_89/a_36_24# 0.01fF
C20 INVX1_LOC_560/A INVX1_LOC_432/A 0.06fF
C21 INVX1_LOC_435/Y INVX1_LOC_435/A 0.00fF
C22 INVX1_LOC_293/Y INVX1_LOC_661/A 0.01fF
C23 INVX1_LOC_553/A INVX1_LOC_361/Y 0.02fF
C24 INVX1_LOC_410/Y INVX1_LOC_48/Y 0.03fF
C25 INVX1_LOC_266/A INVX1_LOC_134/Y 0.04fF
C26 INVX1_LOC_190/Y INVX1_LOC_86/Y 0.01fF
C27 INVX1_LOC_118/Y INVX1_LOC_117/Y 0.03fF
C28 INVX1_LOC_85/Y NAND2X1_LOC_35/a_36_24# 0.00fF
C29 INVX1_LOC_666/A INVX1_LOC_99/Y 0.01fF
C30 INVX1_LOC_384/Y INVX1_LOC_385/Y 11.46fF
C31 VDD INVX1_LOC_199/Y 2.74fF
C32 INVX1_LOC_438/Y INVX1_LOC_6/Y 0.03fF
C33 INVX1_LOC_574/A INVX1_LOC_6/Y 0.28fF
C34 GATE_579 INVX1_LOC_452/A 0.02fF
C35 NAND2X1_LOC_636/A INVX1_LOC_15/Y 0.07fF
C36 INVX1_LOC_133/Y INVX1_LOC_667/Y 0.01fF
C37 INVX1_LOC_238/A NAND2X1_LOC_542/A 0.07fF
C38 INPUT_0 INVX1_LOC_463/Y 0.15fF
C39 INVX1_LOC_533/Y INVX1_LOC_578/Y 0.09fF
C40 INVX1_LOC_20/Y INVX1_LOC_442/Y 0.91fF
C41 INVX1_LOC_370/Y INVX1_LOC_683/Y 0.70fF
C42 INVX1_LOC_420/Y NAND2X1_LOC_346/B 0.01fF
C43 INVX1_LOC_556/Y INVX1_LOC_242/A 0.03fF
C44 INVX1_LOC_80/A INVX1_LOC_679/Y 0.07fF
C45 NAND2X1_LOC_184/Y INVX1_LOC_413/Y 0.20fF
C46 INVX1_LOC_1/A INPUT_4 0.00fF
C47 NAND2X1_LOC_768/A INVX1_LOC_679/Y 0.03fF
C48 INVX1_LOC_217/Y INVX1_LOC_63/Y 0.25fF
C49 INVX1_LOC_420/Y NAND2X1_LOC_274/Y 0.12fF
C50 NAND2X1_LOC_24/Y INVX1_LOC_7/Y 0.07fF
C51 INVX1_LOC_228/Y INVX1_LOC_199/Y 0.03fF
C52 INVX1_LOC_395/A INVX1_LOC_476/A 0.03fF
C53 INVX1_LOC_53/Y NAND2X1_LOC_413/Y 0.11fF
C54 NAND2X1_LOC_173/Y INVX1_LOC_460/Y 0.01fF
C55 INVX1_LOC_97/Y INVX1_LOC_600/A 0.31fF
C56 INVX1_LOC_575/A NAND2X1_LOC_152/B 0.00fF
C57 NAND2X1_LOC_532/a_36_24# NAND2X1_LOC_532/Y 0.02fF
C58 INVX1_LOC_116/Y INVX1_LOC_486/Y 0.17fF
C59 INVX1_LOC_373/A NAND2X1_LOC_334/A 0.00fF
C60 NAND2X1_LOC_101/a_36_24# INVX1_LOC_32/Y 0.01fF
C61 INVX1_LOC_406/Y INVX1_LOC_48/Y 0.00fF
C62 INVX1_LOC_30/Y INPUT_5 0.04fF
C63 NAND2X1_LOC_616/Y NAND2X1_LOC_67/Y 0.01fF
C64 NAND2X1_LOC_79/Y NAND2X1_LOC_243/A 0.01fF
C65 INVX1_LOC_206/Y NAND2X1_LOC_420/Y 0.01fF
C66 INVX1_LOC_21/A INVX1_LOC_83/Y 0.00fF
C67 NAND2X1_LOC_356/a_36_24# INVX1_LOC_58/Y 0.01fF
C68 INVX1_LOC_510/Y INVX1_LOC_199/Y 0.07fF
C69 INVX1_LOC_383/Y INVX1_LOC_510/A 0.02fF
C70 INVX1_LOC_47/Y INVX1_LOC_666/A 0.01fF
C71 INVX1_LOC_586/A INVX1_LOC_69/Y 10.05fF
C72 INPUT_0 NAND2X1_LOC_274/B 0.03fF
C73 INVX1_LOC_321/Y INVX1_LOC_145/Y 0.03fF
C74 INVX1_LOC_312/A INVX1_LOC_117/Y 0.14fF
C75 NAND2X1_LOC_528/a_36_24# INPUT_1 0.01fF
C76 INVX1_LOC_45/Y INVX1_LOC_347/Y 0.03fF
C77 INVX1_LOC_312/Y NAND2X1_LOC_148/B 0.03fF
C78 INVX1_LOC_516/A INVX1_LOC_98/Y 0.01fF
C79 INVX1_LOC_37/Y INVX1_LOC_90/Y 0.01fF
C80 NAND2X1_LOC_391/A INVX1_LOC_117/Y 0.06fF
C81 INVX1_LOC_290/Y INVX1_LOC_632/Y 0.21fF
C82 INVX1_LOC_412/A INVX1_LOC_242/Y 0.46fF
C83 INVX1_LOC_80/A INPUT_1 13.25fF
C84 INVX1_LOC_512/Y INVX1_LOC_58/Y 0.01fF
C85 INVX1_LOC_256/A INVX1_LOC_504/Y 0.01fF
C86 INVX1_LOC_361/Y INVX1_LOC_375/Y 0.00fF
C87 INVX1_LOC_386/Y INVX1_LOC_453/Y 0.04fF
C88 INVX1_LOC_431/A INVX1_LOC_600/A 0.41fF
C89 NAND2X1_LOC_24/Y INVX1_LOC_32/Y 0.04fF
C90 NAND2X1_LOC_673/A INVX1_LOC_99/Y 0.02fF
C91 INVX1_LOC_45/Y INVX1_LOC_328/Y 0.03fF
C92 INVX1_LOC_395/A INVX1_LOC_90/Y 0.05fF
C93 INVX1_LOC_49/Y INVX1_LOC_378/A 0.63fF
C94 NAND2X1_LOC_545/B INVX1_LOC_93/Y 0.03fF
C95 INVX1_LOC_400/A INVX1_LOC_98/Y 0.33fF
C96 INVX1_LOC_558/A INVX1_LOC_9/Y 0.08fF
C97 NAND2X1_LOC_516/Y NAND2X1_LOC_274/B 0.03fF
C98 NAND2X1_LOC_140/B INVX1_LOC_361/Y 0.16fF
C99 INVX1_LOC_266/A INVX1_LOC_65/A 0.03fF
C100 INVX1_LOC_142/A INVX1_LOC_168/Y 0.02fF
C101 INVX1_LOC_47/Y NAND2X1_LOC_273/a_36_24# 0.00fF
C102 INVX1_LOC_194/Y INVX1_LOC_178/A 0.10fF
C103 INVX1_LOC_347/Y INVX1_LOC_348/A 0.00fF
C104 INVX1_LOC_587/Y NAND2X1_LOC_755/B 0.01fF
C105 INVX1_LOC_312/Y INVX1_LOC_69/Y 0.03fF
C106 INPUT_0 INVX1_LOC_148/Y 0.03fF
C107 NAND2X1_LOC_498/B INVX1_LOC_114/A 0.08fF
C108 INVX1_LOC_20/Y INVX1_LOC_482/Y 0.01fF
C109 INVX1_LOC_171/Y INVX1_LOC_245/A 0.01fF
C110 INVX1_LOC_11/Y INVX1_LOC_681/Y 0.01fF
C111 INVX1_LOC_40/Y NAND2X1_LOC_51/a_36_24# 0.00fF
C112 INVX1_LOC_270/A INVX1_LOC_9/Y 0.03fF
C113 INVX1_LOC_268/A INVX1_LOC_6/Y 0.01fF
C114 INVX1_LOC_93/Y INVX1_LOC_98/Y 0.10fF
C115 NAND2X1_LOC_285/A INVX1_LOC_99/Y 0.03fF
C116 INVX1_LOC_282/A NAND2X1_LOC_348/a_36_24# 0.02fF
C117 NAND2X1_LOC_289/a_36_24# INVX1_LOC_98/Y 0.00fF
C118 INPUT_3 INVX1_LOC_328/Y 1.46fF
C119 INVX1_LOC_76/Y INVX1_LOC_114/A 0.03fF
C120 INVX1_LOC_11/Y INPUT_1 2.73fF
C121 INVX1_LOC_145/Y INVX1_LOC_671/Y 0.15fF
C122 NAND2X1_LOC_106/Y INVX1_LOC_367/Y 0.00fF
C123 INVX1_LOC_69/Y NAND2X1_LOC_808/a_36_24# 0.01fF
C124 NAND2X1_LOC_27/Y INVX1_LOC_54/Y 0.02fF
C125 INVX1_LOC_507/Y INVX1_LOC_633/Y 0.02fF
C126 INVX1_LOC_671/Y INVX1_LOC_661/Y 0.03fF
C127 INVX1_LOC_663/Y INVX1_LOC_671/A 0.02fF
C128 INVX1_LOC_160/A NAND2X1_LOC_169/a_36_24# 0.00fF
C129 INVX1_LOC_544/A INVX1_LOC_6/Y 0.74fF
C130 INVX1_LOC_323/Y INVX1_LOC_63/Y 0.03fF
C131 NAND2X1_LOC_388/A INVX1_LOC_252/Y 0.05fF
C132 INVX1_LOC_137/Y INVX1_LOC_496/Y 0.00fF
C133 INVX1_LOC_105/A INVX1_LOC_105/Y 0.01fF
C134 NAND2X1_LOC_76/a_36_24# INVX1_LOC_211/A 0.00fF
C135 NAND2X1_LOC_336/B INVX1_LOC_242/Y 0.12fF
C136 INVX1_LOC_516/A INVX1_LOC_338/Y 0.02fF
C137 INVX1_LOC_119/Y NAND2X1_LOC_273/a_36_24# 0.00fF
C138 INVX1_LOC_219/Y INVX1_LOC_6/Y 0.00fF
C139 NAND2X1_LOC_750/Y NAND2X1_LOC_60/Y 0.00fF
C140 NAND2X1_LOC_333/A NAND2X1_LOC_720/A 0.00fF
C141 INVX1_LOC_385/Y NAND2X1_LOC_555/B 0.03fF
C142 INVX1_LOC_291/A INVX1_LOC_531/Y 0.01fF
C143 NAND2X1_LOC_673/A NAND2X1_LOC_557/B 0.03fF
C144 INVX1_LOC_370/Y INVX1_LOC_682/Y 0.12fF
C145 INVX1_LOC_300/Y INVX1_LOC_684/Y 0.01fF
C146 INVX1_LOC_270/A INVX1_LOC_62/Y 0.01fF
C147 INVX1_LOC_44/Y INVX1_LOC_178/A 0.07fF
C148 INVX1_LOC_304/A INVX1_LOC_411/Y 0.00fF
C149 INVX1_LOC_58/Y INVX1_LOC_194/Y 1.20fF
C150 INVX1_LOC_463/Y INVX1_LOC_498/A 0.03fF
C151 INVX1_LOC_390/A INVX1_LOC_98/Y 0.07fF
C152 INVX1_LOC_12/Y INVX1_LOC_100/Y 0.19fF
C153 INVX1_LOC_21/Y INVX1_LOC_652/A 0.00fF
C154 INVX1_LOC_301/Y INVX1_LOC_35/Y 0.02fF
C155 INVX1_LOC_201/Y INVX1_LOC_399/Y 0.00fF
C156 INVX1_LOC_211/Y INVX1_LOC_9/Y 0.13fF
C157 INVX1_LOC_372/Y INVX1_LOC_74/Y 1.02fF
C158 INVX1_LOC_306/Y INVX1_LOC_46/Y 0.02fF
C159 NAND2X1_LOC_835/A INVX1_LOC_69/Y 0.02fF
C160 INVX1_LOC_682/A INVX1_LOC_159/Y 0.00fF
C161 INVX1_LOC_93/Y INVX1_LOC_338/Y 0.11fF
C162 INVX1_LOC_213/Y NAND2X1_LOC_106/a_36_24# 0.00fF
C163 NAND2X1_LOC_788/a_36_24# NAND2X1_LOC_274/B 0.00fF
C164 INVX1_LOC_169/Y INVX1_LOC_480/A 0.04fF
C165 INVX1_LOC_49/Y NAND2X1_LOC_632/a_36_24# 0.00fF
C166 INVX1_LOC_69/Y INVX1_LOC_157/Y 0.03fF
C167 INVX1_LOC_53/Y INVX1_LOC_645/Y 0.09fF
C168 INVX1_LOC_12/Y INVX1_LOC_74/Y 0.03fF
C169 NAND2X1_LOC_755/B INVX1_LOC_62/Y 0.03fF
C170 NAND2X1_LOC_542/A NAND2X1_LOC_280/a_36_24# 0.01fF
C171 INVX1_LOC_501/A NAND2X1_LOC_689/B 0.03fF
C172 INVX1_LOC_12/Y INVX1_LOC_483/Y 0.02fF
C173 INVX1_LOC_7/Y INVX1_LOC_190/A 0.16fF
C174 NAND2X1_LOC_704/B INVX1_LOC_92/A 0.07fF
C175 INVX1_LOC_46/Y INVX1_LOC_9/Y 0.62fF
C176 INVX1_LOC_254/Y INVX1_LOC_79/A 0.03fF
C177 INVX1_LOC_304/A INVX1_LOC_41/Y 0.01fF
C178 INVX1_LOC_35/Y INVX1_LOC_41/Y 1.40fF
C179 INVX1_LOC_211/Y INVX1_LOC_62/Y 0.03fF
C180 INVX1_LOC_179/A INVX1_LOC_6/Y 0.00fF
C181 NAND2X1_LOC_719/A INVX1_LOC_6/Y 0.15fF
C182 INVX1_LOC_507/A INVX1_LOC_496/A 0.04fF
C183 INVX1_LOC_557/Y INVX1_LOC_66/A 0.02fF
C184 INVX1_LOC_519/Y INVX1_LOC_670/A 0.01fF
C185 INVX1_LOC_89/Y INVX1_LOC_245/A 0.07fF
C186 INVX1_LOC_665/A INVX1_LOC_50/Y 0.03fF
C187 INVX1_LOC_44/Y INVX1_LOC_58/Y 0.18fF
C188 INVX1_LOC_31/Y INVX1_LOC_90/Y 0.11fF
C189 NAND2X1_LOC_305/a_36_24# INVX1_LOC_9/Y 0.00fF
C190 NAND2X1_LOC_62/a_36_24# INVX1_LOC_98/Y 0.07fF
C191 INVX1_LOC_154/A INVX1_LOC_245/A 0.00fF
C192 INVX1_LOC_335/Y INVX1_LOC_462/Y 0.01fF
C193 INVX1_LOC_505/Y INVX1_LOC_50/Y 0.09fF
C194 INVX1_LOC_592/Y INVX1_LOC_79/A 0.03fF
C195 INVX1_LOC_513/A INVX1_LOC_588/A 0.06fF
C196 INVX1_LOC_62/Y INVX1_LOC_46/Y 0.58fF
C197 INVX1_LOC_501/A INVX1_LOC_245/A 0.02fF
C198 NAND2X1_LOC_663/a_36_24# INVX1_LOC_669/A 0.00fF
C199 NAND2X1_LOC_341/a_36_24# NAND2X1_LOC_231/B 0.00fF
C200 INVX1_LOC_376/A INVX1_LOC_373/Y 0.03fF
C201 INVX1_LOC_13/Y INVX1_LOC_46/Y 0.02fF
C202 INVX1_LOC_439/Y INVX1_LOC_443/A 0.23fF
C203 NAND2X1_LOC_475/A NAND2X1_LOC_170/a_36_24# 0.00fF
C204 INVX1_LOC_58/Y INVX1_LOC_347/A 0.07fF
C205 INVX1_LOC_301/A INVX1_LOC_412/A 0.46fF
C206 INVX1_LOC_482/A INVX1_LOC_297/Y 0.00fF
C207 NAND2X1_LOC_790/B INVX1_LOC_94/A 0.04fF
C208 NAND2X1_LOC_118/a_36_24# INVX1_LOC_79/A 0.01fF
C209 NAND2X1_LOC_249/Y NAND2X1_LOC_142/Y 0.02fF
C210 INVX1_LOC_75/A INVX1_LOC_9/Y 0.01fF
C211 NAND2X1_LOC_528/Y INVX1_LOC_79/A 0.42fF
C212 INVX1_LOC_560/Y INVX1_LOC_249/Y 0.02fF
C213 VDD INVX1_LOC_459/Y 0.35fF
C214 INVX1_LOC_479/A INVX1_LOC_79/A 0.20fF
C215 NAND2X1_LOC_161/a_36_24# INVX1_LOC_542/A 0.00fF
C216 INVX1_LOC_653/A NAND2X1_LOC_832/A 0.09fF
C217 INVX1_LOC_600/A INVX1_LOC_615/A 0.16fF
C218 INVX1_LOC_446/A INVX1_LOC_519/A 0.04fF
C219 INVX1_LOC_62/Y INVX1_LOC_75/A 0.01fF
C220 INVX1_LOC_301/A NAND2X1_LOC_336/B 0.00fF
C221 INVX1_LOC_521/Y INVX1_LOC_185/Y 0.02fF
C222 INVX1_LOC_165/Y INVX1_LOC_45/Y 0.04fF
C223 VDD INVX1_LOC_53/Y 1.34fF
C224 INVX1_LOC_412/Y INVX1_LOC_634/A 0.01fF
C225 INVX1_LOC_586/A NAND2X1_LOC_419/a_36_24# 0.00fF
C226 INVX1_LOC_266/Y INVX1_LOC_45/Y 0.03fF
C227 INVX1_LOC_317/Y NAND2X1_LOC_315/a_36_24# 0.01fF
C228 INVX1_LOC_560/Y INVX1_LOC_248/Y 0.28fF
C229 INVX1_LOC_576/Y INVX1_LOC_561/Y 0.04fF
C230 INVX1_LOC_625/A INVX1_LOC_616/Y 0.03fF
C231 NAND2X1_LOC_58/a_36_24# INVX1_LOC_178/A 0.01fF
C232 INVX1_LOC_20/Y NAND2X1_LOC_707/A 0.07fF
C233 INVX1_LOC_76/Y INVX1_LOC_482/A 0.00fF
C234 NAND2X1_LOC_523/B INVX1_LOC_362/Y 0.09fF
C235 NAND2X1_LOC_475/A INVX1_LOC_681/A 0.02fF
C236 INVX1_LOC_355/A INVX1_LOC_134/Y 0.01fF
C237 INVX1_LOC_20/Y NAND2X1_LOC_493/B 0.01fF
C238 INVX1_LOC_312/Y INVX1_LOC_586/A 0.03fF
C239 VDD INVX1_LOC_460/Y 0.56fF
C240 INVX1_LOC_359/A INVX1_LOC_638/A 0.05fF
C241 NAND2X1_LOC_781/A INVX1_LOC_586/A 0.01fF
C242 INVX1_LOC_53/Y INVX1_LOC_510/Y 0.07fF
C243 INVX1_LOC_134/A INVX1_LOC_80/A 0.00fF
C244 VDD INVX1_LOC_43/A -0.00fF
C245 INVX1_LOC_224/Y INVX1_LOC_304/Y 0.02fF
C246 NAND2X1_LOC_466/a_36_24# INVX1_LOC_638/A 0.01fF
C247 NAND2X1_LOC_525/Y INVX1_LOC_99/Y 0.07fF
C248 INVX1_LOC_395/A INVX1_LOC_98/Y 0.01fF
C249 INVX1_LOC_617/Y NAND2X1_LOC_710/A 0.00fF
C250 INPUT_0 INVX1_LOC_159/Y 0.03fF
C251 INVX1_LOC_607/Y INVX1_LOC_237/Y 0.06fF
C252 VDD NAND2X1_LOC_400/B 0.02fF
C253 INVX1_LOC_435/Y INVX1_LOC_392/A 0.03fF
C254 NAND2X1_LOC_331/A INVX1_LOC_493/A 0.00fF
C255 VDD NAND2X1_LOC_346/B 0.01fF
C256 INVX1_LOC_578/A INVX1_LOC_304/Y 0.01fF
C257 INVX1_LOC_419/Y INVX1_LOC_400/Y 0.16fF
C258 NAND2X1_LOC_79/Y INVX1_LOC_619/A 0.06fF
C259 INVX1_LOC_596/A INVX1_LOC_367/A 0.07fF
C260 INVX1_LOC_522/Y INVX1_LOC_633/Y 0.03fF
C261 INVX1_LOC_118/Y INVX1_LOC_608/A 0.23fF
C262 INVX1_LOC_438/Y NAND2X1_LOC_294/Y 0.03fF
C263 NAND2X1_LOC_513/Y INVX1_LOC_61/A 0.10fF
C264 INVX1_LOC_617/Y INVX1_LOC_383/Y 0.03fF
C265 VDD NAND2X1_LOC_274/Y 0.21fF
C266 NAND2X1_LOC_551/a_36_24# INVX1_LOC_578/A 0.01fF
C267 INVX1_LOC_449/A INVX1_LOC_293/Y 0.07fF
C268 INVX1_LOC_315/Y INVX1_LOC_35/Y 0.04fF
C269 INVX1_LOC_300/A NAND2X1_LOC_493/B 0.01fF
C270 INVX1_LOC_614/A INVX1_LOC_53/Y 0.12fF
C271 INVX1_LOC_139/A NAND2X1_LOC_707/B 0.00fF
C272 INVX1_LOC_578/A NAND2X1_LOC_444/A 0.04fF
C273 INVX1_LOC_194/A INVX1_LOC_76/Y 0.02fF
C274 INVX1_LOC_435/Y INVX1_LOC_93/Y 1.16fF
C275 INVX1_LOC_435/Y INVX1_LOC_283/A 0.07fF
C276 INVX1_LOC_142/A INVX1_LOC_137/Y 0.01fF
C277 INVX1_LOC_122/Y NAND2X1_LOC_542/A 0.01fF
C278 VDD NAND2X1_LOC_406/B 0.01fF
C279 INVX1_LOC_439/Y NAND2X1_LOC_261/Y 0.33fF
C280 INVX1_LOC_105/Y INVX1_LOC_45/Y 0.03fF
C281 INVX1_LOC_19/Y INPUT_5 0.01fF
C282 INVX1_LOC_85/Y NAND2X1_LOC_235/a_36_24# 0.00fF
C283 NAND2X1_LOC_79/B INVX1_LOC_198/A 0.00fF
C284 INVX1_LOC_414/Y INVX1_LOC_387/Y 0.01fF
C285 INVX1_LOC_288/A INVX1_LOC_372/A 0.03fF
C286 NAND2X1_LOC_324/B INVX1_LOC_504/Y 0.01fF
C287 INVX1_LOC_203/Y INVX1_LOC_245/A 1.16fF
C288 INVX1_LOC_587/Y INVX1_LOC_268/Y 0.15fF
C289 NAND2X1_LOC_57/Y INVX1_LOC_12/Y 0.05fF
C290 INVX1_LOC_105/A INVX1_LOC_126/Y 0.00fF
C291 INVX1_LOC_117/Y INPUT_2 0.02fF
C292 NAND2X1_LOC_399/B NAND2X1_LOC_398/a_36_24# 0.04fF
C293 INVX1_LOC_117/Y INVX1_LOC_126/A 0.02fF
C294 INVX1_LOC_586/A INVX1_LOC_157/Y 0.03fF
C295 INVX1_LOC_21/Y INVX1_LOC_379/A 0.07fF
C296 NAND2X1_LOC_45/a_36_24# NAND2X1_LOC_274/B 0.00fF
C297 INVX1_LOC_17/Y INVX1_LOC_344/Y -0.00fF
C298 INVX1_LOC_578/A NAND2X1_LOC_167/a_36_24# 0.01fF
C299 NAND2X1_LOC_399/B NAND2X1_LOC_403/A 0.05fF
C300 INVX1_LOC_96/Y INVX1_LOC_58/Y 0.03fF
C301 NAND2X1_LOC_403/A INVX1_LOC_7/Y 0.07fF
C302 NAND2X1_LOC_229/a_36_24# INVX1_LOC_96/A 0.00fF
C303 NAND2X1_LOC_333/A INVX1_LOC_566/A 0.01fF
C304 INVX1_LOC_21/Y INVX1_LOC_35/Y 5.69fF
C305 INVX1_LOC_254/A INVX1_LOC_318/Y 0.08fF
C306 NAND2X1_LOC_341/a_36_24# INVX1_LOC_80/A 0.01fF
C307 INVX1_LOC_587/A INVX1_LOC_69/Y 0.81fF
C308 NAND2X1_LOC_331/A INVX1_LOC_500/A 0.01fF
C309 INVX1_LOC_469/Y INVX1_LOC_372/Y 0.02fF
C310 NAND2X1_LOC_505/Y INVX1_LOC_351/A 0.05fF
C311 NAND2X1_LOC_733/a_36_24# INVX1_LOC_674/A 0.00fF
C312 INVX1_LOC_549/Y INVX1_LOC_145/Y 0.09fF
C313 NAND2X1_LOC_685/B INVX1_LOC_58/Y 0.01fF
C314 INVX1_LOC_596/A INVX1_LOC_93/Y 0.01fF
C315 INVX1_LOC_80/A INVX1_LOC_50/Y 5.32fF
C316 NAND2X1_LOC_231/B INVX1_LOC_275/A 0.04fF
C317 VDD INVX1_LOC_368/Y 0.21fF
C318 INVX1_LOC_7/Y INVX1_LOC_453/Y 0.09fF
C319 INVX1_LOC_254/Y INVX1_LOC_417/Y 0.36fF
C320 INVX1_LOC_53/Y INVX1_LOC_103/Y 0.01fF
C321 INVX1_LOC_137/Y INVX1_LOC_99/Y 0.06fF
C322 INVX1_LOC_566/A INVX1_LOC_188/A 0.18fF
C323 VDD NAND2X1_LOC_451/B 0.12fF
C324 INVX1_LOC_609/A INVX1_LOC_137/Y 0.01fF
C325 NAND2X1_LOC_526/Y INVX1_LOC_26/Y 0.02fF
C326 NAND2X1_LOC_727/a_36_24# NAND2X1_LOC_274/B 0.00fF
C327 NAND2X1_LOC_791/B INVX1_LOC_69/Y 0.20fF
C328 INVX1_LOC_20/Y NAND2X1_LOC_847/A 0.12fF
C329 INVX1_LOC_11/Y INVX1_LOC_428/Y 0.08fF
C330 INVX1_LOC_413/A INVX1_LOC_17/Y 0.08fF
C331 INVX1_LOC_686/A NAND2X1_LOC_586/Y 0.00fF
C332 INVX1_LOC_435/A INVX1_LOC_294/A 0.01fF
C333 INVX1_LOC_254/Y INVX1_LOC_59/Y 0.01fF
C334 NAND2X1_LOC_318/A INVX1_LOC_9/Y 0.47fF
C335 INVX1_LOC_53/Y INVX1_LOC_346/A 0.03fF
C336 INVX1_LOC_51/Y INVX1_LOC_90/Y 0.09fF
C337 INVX1_LOC_671/Y NAND2X1_LOC_260/Y 0.03fF
C338 NAND2X1_LOC_516/Y INVX1_LOC_468/A 0.07fF
C339 NAND2X1_LOC_403/A INVX1_LOC_32/Y 0.00fF
C340 INVX1_LOC_384/A NAND2X1_LOC_274/B 0.00fF
C341 INVX1_LOC_11/Y INVX1_LOC_50/Y 0.33fF
C342 INVX1_LOC_254/Y INVX1_LOC_48/Y 0.06fF
C343 INVX1_LOC_31/Y INVX1_LOC_98/Y 0.12fF
C344 INVX1_LOC_42/Y INVX1_LOC_46/Y 0.01fF
C345 INVX1_LOC_293/Y INVX1_LOC_328/Y 2.00fF
C346 INVX1_LOC_406/A INVX1_LOC_99/Y 0.00fF
C347 INPUT_3 INVX1_LOC_224/A 0.00fF
C348 INVX1_LOC_147/A INVX1_LOC_58/Y 0.01fF
C349 VDD NAND2X1_LOC_60/Y 0.05fF
C350 INVX1_LOC_32/Y INVX1_LOC_259/Y 0.03fF
C351 NAND2X1_LOC_667/a_36_24# INVX1_LOC_50/Y 0.00fF
C352 INVX1_LOC_555/A INVX1_LOC_35/Y 0.01fF
C353 INVX1_LOC_607/Y INVX1_LOC_212/Y 0.08fF
C354 INVX1_LOC_54/Y INVX1_LOC_543/Y 0.39fF
C355 INVX1_LOC_58/Y NAND2X1_LOC_418/Y 0.14fF
C356 INVX1_LOC_387/Y INVX1_LOC_303/Y 0.00fF
C357 INVX1_LOC_219/Y NAND2X1_LOC_294/Y 0.01fF
C358 NAND2X1_LOC_773/A INVX1_LOC_207/Y 0.03fF
C359 VDD INVX1_LOC_636/Y 0.21fF
C360 INPUT_1 INVX1_LOC_374/Y 0.01fF
C361 INVX1_LOC_372/Y INVX1_LOC_79/A 0.06fF
C362 INVX1_LOC_556/Y NAND2X1_LOC_542/A 0.00fF
C363 INVX1_LOC_47/Y INVX1_LOC_137/Y 0.02fF
C364 INVX1_LOC_166/A NAND2X1_LOC_313/a_36_24# 0.00fF
C365 INVX1_LOC_32/Y NAND2X1_LOC_707/B 0.23fF
C366 INVX1_LOC_298/A INVX1_LOC_340/A 0.03fF
C367 INVX1_LOC_120/Y INVX1_LOC_304/Y 0.11fF
C368 INVX1_LOC_492/Y INVX1_LOC_475/Y 0.01fF
C369 INVX1_LOC_346/A INVX1_LOC_460/Y 0.01fF
C370 INVX1_LOC_49/Y INVX1_LOC_303/Y 0.01fF
C371 INVX1_LOC_448/A NAND2X1_LOC_274/B 0.46fF
C372 INVX1_LOC_12/Y INVX1_LOC_79/A 0.03fF
C373 INVX1_LOC_65/Y NAND2X1_LOC_201/a_36_24# 0.01fF
C374 NAND2X1_LOC_169/A INVX1_LOC_242/Y 0.04fF
C375 NAND2X1_LOC_787/a_36_24# INVX1_LOC_301/Y 0.00fF
C376 INVX1_LOC_587/Y INVX1_LOC_49/Y 0.24fF
C377 NAND2X1_LOC_274/B INVX1_LOC_145/Y 0.03fF
C378 NAND2X1_LOC_616/a_36_24# INVX1_LOC_178/A 0.01fF
C379 INPUT_7 INVX1_LOC_25/A 0.27fF
C380 INVX1_LOC_53/Y INVX1_LOC_635/Y 0.03fF
C381 INVX1_LOC_256/A INVX1_LOC_114/A 0.00fF
C382 NAND2X1_LOC_387/Y INVX1_LOC_551/A 0.04fF
C383 INVX1_LOC_194/Y INVX1_LOC_245/A 0.45fF
C384 INVX1_LOC_69/Y INVX1_LOC_6/Y 0.06fF
C385 INVX1_LOC_679/Y NAND2X1_LOC_843/B 0.02fF
C386 INVX1_LOC_21/Y INVX1_LOC_79/Y 0.01fF
C387 INVX1_LOC_523/Y INVX1_LOC_58/Y 0.19fF
C388 INVX1_LOC_520/Y INVX1_LOC_89/Y 0.01fF
C389 INVX1_LOC_137/Y INVX1_LOC_119/Y 0.01fF
C390 INVX1_LOC_632/A INVX1_LOC_479/A 0.08fF
C391 INVX1_LOC_62/Y INVX1_LOC_115/A 0.07fF
C392 NAND2X1_LOC_851/a_36_24# INVX1_LOC_655/A -0.01fF
C393 INVX1_LOC_338/A INVX1_LOC_41/Y 0.00fF
C394 INVX1_LOC_509/Y INVX1_LOC_479/A 0.03fF
C395 INVX1_LOC_506/A INVX1_LOC_376/Y 0.02fF
C396 INVX1_LOC_417/Y INVX1_LOC_479/A 0.49fF
C397 INVX1_LOC_100/Y NAND2X1_LOC_615/B 0.22fF
C398 INVX1_LOC_479/A INVX1_LOC_491/Y 0.03fF
C399 INVX1_LOC_387/Y INVX1_LOC_9/Y 0.00fF
C400 INVX1_LOC_345/Y INVX1_LOC_114/A 1.23fF
C401 INVX1_LOC_62/Y INVX1_LOC_349/Y 0.01fF
C402 INVX1_LOC_202/Y INVX1_LOC_62/Y 0.03fF
C403 INVX1_LOC_254/A INVX1_LOC_90/Y 0.01fF
C404 INVX1_LOC_32/Y INVX1_LOC_114/A 0.03fF
C405 INVX1_LOC_479/A INVX1_LOC_59/Y 0.28fF
C406 INVX1_LOC_41/Y INVX1_LOC_360/A 0.01fF
C407 INVX1_LOC_421/A INVX1_LOC_502/A 0.04fF
C408 NAND2X1_LOC_333/A INVX1_LOC_79/A 0.05fF
C409 INVX1_LOC_49/Y INVX1_LOC_9/Y 0.10fF
C410 NAND2X1_LOC_615/B INVX1_LOC_74/Y 0.09fF
C411 INPUT_1 NAND2X1_LOC_843/B 0.03fF
C412 INVX1_LOC_100/Y INVX1_LOC_66/A 0.21fF
C413 INVX1_LOC_479/A INVX1_LOC_48/Y 1.29fF
C414 INVX1_LOC_44/Y INVX1_LOC_245/A 0.03fF
C415 INVX1_LOC_387/Y INVX1_LOC_62/Y 0.03fF
C416 NAND2X1_LOC_847/A INVX1_LOC_655/A 0.73fF
C417 INVX1_LOC_170/A INVX1_LOC_79/A 0.01fF
C418 INVX1_LOC_526/Y INVX1_LOC_636/A 0.05fF
C419 INVX1_LOC_45/Y INVX1_LOC_109/Y 0.01fF
C420 INVX1_LOC_49/Y INVX1_LOC_166/Y 0.01fF
C421 INVX1_LOC_258/Y NAND2X1_LOC_123/B 0.10fF
C422 INPUT_1 INVX1_LOC_625/Y 0.13fF
C423 INVX1_LOC_74/Y INVX1_LOC_66/A 0.09fF
C424 INVX1_LOC_387/Y NAND2X1_LOC_844/A 0.00fF
C425 INVX1_LOC_338/Y INVX1_LOC_473/Y 0.37fF
C426 INVX1_LOC_49/Y INVX1_LOC_62/Y 0.12fF
C427 INVX1_LOC_95/Y NAND2X1_LOC_506/B 0.33fF
C428 INVX1_LOC_531/Y INVX1_LOC_223/Y 0.00fF
C429 INVX1_LOC_49/Y NAND2X1_LOC_844/A 0.03fF
C430 INVX1_LOC_95/Y INVX1_LOC_45/Y 0.05fF
C431 INVX1_LOC_361/Y INVX1_LOC_92/A 0.07fF
C432 NAND2X1_LOC_409/Y INVX1_LOC_35/A 0.00fF
C433 INVX1_LOC_100/Y NAND2X1_LOC_601/Y 0.11fF
C434 INVX1_LOC_662/A INVX1_LOC_645/Y 0.06fF
C435 INVX1_LOC_675/A INVX1_LOC_346/Y 0.03fF
C436 NAND2X1_LOC_242/A INVX1_LOC_604/A 0.03fF
C437 INVX1_LOC_100/Y NAND2X1_LOC_621/B 0.04fF
C438 VDD NAND2X1_LOC_383/Y 0.47fF
C439 VDD INVX1_LOC_555/Y 0.21fF
C440 INVX1_LOC_414/A NAND2X1_LOC_553/a_36_24# 0.00fF
C441 INVX1_LOC_80/A INVX1_LOC_275/A 0.33fF
C442 INVX1_LOC_629/Y NAND2X1_LOC_173/Y 0.05fF
C443 INVX1_LOC_435/Y INVX1_LOC_362/Y 0.03fF
C444 NAND2X1_LOC_786/B NAND2X1_LOC_60/Y 0.03fF
C445 INVX1_LOC_483/Y NAND2X1_LOC_621/B 0.15fF
C446 VDD NAND2X1_LOC_107/Y 0.03fF
C447 INVX1_LOC_438/A INVX1_LOC_80/A 0.01fF
C448 NAND2X1_LOC_372/a_36_24# INVX1_LOC_362/Y 0.00fF
C449 INVX1_LOC_395/A INVX1_LOC_596/A 0.02fF
C450 NAND2X1_LOC_710/A INVX1_LOC_375/A 0.03fF
C451 INVX1_LOC_45/Y NAND2X1_LOC_427/Y 0.01fF
C452 NAND2X1_LOC_43/a_36_24# INVX1_LOC_176/A 0.01fF
C453 INVX1_LOC_410/Y INVX1_LOC_383/Y 0.03fF
C454 INVX1_LOC_20/Y NAND2X1_LOC_231/A 0.01fF
C455 INVX1_LOC_400/A NAND2X1_LOC_76/B 0.01fF
C456 NAND2X1_LOC_498/Y NAND2X1_LOC_307/A 0.07fF
C457 NAND2X1_LOC_498/Y INVX1_LOC_545/Y 0.03fF
C458 NAND2X1_LOC_524/a_36_24# INVX1_LOC_412/A 0.01fF
C459 INVX1_LOC_596/A INVX1_LOC_362/Y 0.07fF
C460 INVX1_LOC_395/A NAND2X1_LOC_318/B 0.06fF
C461 VDD INVX1_LOC_213/Y 0.44fF
C462 NAND2X1_LOC_345/a_36_24# INVX1_LOC_384/Y 0.01fF
C463 INVX1_LOC_272/Y INVX1_LOC_586/A 0.01fF
C464 VDD INVX1_LOC_439/Y 2.89fF
C465 INVX1_LOC_586/A INVX1_LOC_486/Y 0.33fF
C466 INVX1_LOC_584/A INVX1_LOC_17/Y 0.91fF
C467 INVX1_LOC_438/A INVX1_LOC_11/Y 0.08fF
C468 INVX1_LOC_293/Y INVX1_LOC_651/Y 0.13fF
C469 INVX1_LOC_614/A INVX1_LOC_555/Y 0.03fF
C470 INVX1_LOC_276/A INVX1_LOC_651/A 0.05fF
C471 INVX1_LOC_85/Y NAND2X1_LOC_789/a_36_24# 0.00fF
C472 NAND2X1_LOC_13/Y INVX1_LOC_318/Y 0.00fF
C473 NAND2X1_LOC_209/a_36_24# INVX1_LOC_6/Y 0.00fF
C474 INVX1_LOC_406/Y NAND2X1_LOC_541/B 0.01fF
C475 INVX1_LOC_395/A INVX1_LOC_177/A 0.03fF
C476 INVX1_LOC_295/A INVX1_LOC_235/Y 0.02fF
C477 NAND2X1_LOC_320/Y INVX1_LOC_45/Y 0.02fF
C478 INVX1_LOC_428/A INVX1_LOC_391/Y 0.01fF
C479 INVX1_LOC_295/A NAND2X1_LOC_361/a_36_24# 0.02fF
C480 NAND2X1_LOC_457/A INVX1_LOC_32/Y 0.03fF
C481 INVX1_LOC_335/Y NAND2X1_LOC_120/a_36_24# 0.01fF
C482 INVX1_LOC_11/Y INVX1_LOC_441/Y 0.01fF
C483 INVX1_LOC_564/A INVX1_LOC_50/Y 0.03fF
C484 INVX1_LOC_312/Y INVX1_LOC_486/Y 0.20fF
C485 INVX1_LOC_404/Y INVX1_LOC_46/Y 0.03fF
C486 INVX1_LOC_51/Y INVX1_LOC_98/Y 0.10fF
C487 INVX1_LOC_554/A INVX1_LOC_89/A 0.01fF
C488 INVX1_LOC_578/A NAND2X1_LOC_454/a_36_24# 0.01fF
C489 INVX1_LOC_166/A NAND2X1_LOC_704/a_36_24# 0.00fF
C490 INVX1_LOC_425/A NAND2X1_LOC_143/a_36_24# 0.00fF
C491 VDD NAND2X1_LOC_698/Y 0.00fF
C492 VDD INVX1_LOC_544/Y 0.22fF
C493 INVX1_LOC_315/Y NAND2X1_LOC_837/B 0.05fF
C494 INVX1_LOC_20/Y INVX1_LOC_321/Y 0.05fF
C495 INVX1_LOC_266/A INVX1_LOC_98/Y 0.10fF
C496 INVX1_LOC_297/A INVX1_LOC_281/Y 0.01fF
C497 INVX1_LOC_62/Y INVX1_LOC_297/Y 0.03fF
C498 VDD INVX1_LOC_662/A 0.05fF
C499 INVX1_LOC_166/A NAND2X1_LOC_188/a_36_24# 0.00fF
C500 INVX1_LOC_33/Y INVX1_LOC_18/Y 0.00fF
C501 NAND2X1_LOC_237/Y INVX1_LOC_600/A 0.06fF
C502 INVX1_LOC_417/Y INVX1_LOC_12/Y 0.02fF
C503 INVX1_LOC_206/Y INVX1_LOC_183/A 0.13fF
C504 NAND2X1_LOC_715/a_36_24# NAND2X1_LOC_137/A 0.00fF
C505 NAND2X1_LOC_49/a_36_24# INVX1_LOC_183/A 0.00fF
C506 INVX1_LOC_587/A NAND2X1_LOC_835/A 0.02fF
C507 NAND2X1_LOC_324/a_36_24# INVX1_LOC_633/Y 0.01fF
C508 NAND2X1_LOC_551/a_36_24# INVX1_LOC_686/A 0.01fF
C509 INVX1_LOC_586/A INVX1_LOC_6/Y 1.15fF
C510 INVX1_LOC_12/Y INVX1_LOC_59/Y 1.05fF
C511 INVX1_LOC_566/Y INVX1_LOC_50/Y 0.01fF
C512 INVX1_LOC_35/Y INVX1_LOC_474/Y 0.23fF
C513 INVX1_LOC_45/Y INVX1_LOC_199/Y 0.14fF
C514 NAND2X1_LOC_45/Y INVX1_LOC_502/A 0.10fF
C515 NAND2X1_LOC_187/Y INVX1_LOC_197/A 0.00fF
C516 INVX1_LOC_155/A INVX1_LOC_76/Y 0.07fF
C517 INVX1_LOC_438/Y INVX1_LOC_100/Y 0.05fF
C518 INVX1_LOC_51/Y INVX1_LOC_338/Y 0.97fF
C519 INVX1_LOC_580/Y INVX1_LOC_49/Y 0.02fF
C520 INVX1_LOC_367/A INVX1_LOC_520/A 0.03fF
C521 INVX1_LOC_18/A INVX1_LOC_29/Y 0.01fF
C522 INVX1_LOC_192/Y INVX1_LOC_79/A 0.01fF
C523 INVX1_LOC_625/A INVX1_LOC_400/A 0.33fF
C524 INVX1_LOC_210/Y INVX1_LOC_274/A 0.02fF
C525 INVX1_LOC_12/Y INVX1_LOC_48/Y 0.15fF
C526 NAND2X1_LOC_707/A INVX1_LOC_494/Y 0.03fF
C527 NAND2X1_LOC_788/A INVX1_LOC_74/Y 0.01fF
C528 INVX1_LOC_35/Y INVX1_LOC_481/Y 0.02fF
C529 INVX1_LOC_444/Y INVX1_LOC_35/Y 0.03fF
C530 INVX1_LOC_634/Y INVX1_LOC_638/A 0.00fF
C531 INVX1_LOC_52/Y INVX1_LOC_41/Y 0.01fF
C532 INVX1_LOC_419/Y INVX1_LOC_99/Y 0.02fF
C533 INVX1_LOC_604/A INVX1_LOC_79/A 0.01fF
C534 INVX1_LOC_446/Y INVX1_LOC_405/Y 0.06fF
C535 INVX1_LOC_145/Y INVX1_LOC_159/Y 0.04fF
C536 INVX1_LOC_312/Y INVX1_LOC_6/Y 0.03fF
C537 INPUT_4 INVX1_LOC_29/Y 0.03fF
C538 INVX1_LOC_45/Y INVX1_LOC_272/A 0.00fF
C539 INVX1_LOC_80/A NAND2X1_LOC_388/A 0.03fF
C540 INVX1_LOC_283/Y INVX1_LOC_661/A 0.09fF
C541 NAND2X1_LOC_318/B INVX1_LOC_31/Y 0.21fF
C542 NAND2X1_LOC_307/A INVX1_LOC_47/Y 0.08fF
C543 INVX1_LOC_76/Y INVX1_LOC_9/Y 0.29fF
C544 INVX1_LOC_367/Y INVX1_LOC_50/Y 0.11fF
C545 INVX1_LOC_442/A INVX1_LOC_100/Y 0.16fF
C546 INVX1_LOC_662/Y INVX1_LOC_672/A 0.02fF
C547 NAND2X1_LOC_332/B NAND2X1_LOC_137/a_36_24# 0.00fF
C548 INVX1_LOC_625/A NAND2X1_LOC_289/a_36_24# 0.01fF
C549 NAND2X1_LOC_332/B NAND2X1_LOC_274/B 0.03fF
C550 NAND2X1_LOC_779/a_36_24# INVX1_LOC_54/Y 0.00fF
C551 INVX1_LOC_134/Y NAND2X1_LOC_449/B 0.02fF
C552 INVX1_LOC_54/Y NAND2X1_LOC_106/B 0.04fF
C553 INVX1_LOC_31/Y INVX1_LOC_504/A 0.07fF
C554 INVX1_LOC_206/Y INVX1_LOC_109/A 0.02fF
C555 INVX1_LOC_455/A INVX1_LOC_298/A 0.14fF
C556 NAND2X1_LOC_333/A INVX1_LOC_59/Y 0.02fF
C557 INVX1_LOC_261/Y INVX1_LOC_602/Y 0.03fF
C558 INVX1_LOC_596/A INVX1_LOC_682/Y 0.07fF
C559 INVX1_LOC_407/Y INVX1_LOC_46/Y 0.01fF
C560 NAND2X1_LOC_498/B INVX1_LOC_62/Y 0.01fF
C561 NAND2X1_LOC_106/Y NAND2X1_LOC_692/Y 0.01fF
C562 NAND2X1_LOC_13/Y INVX1_LOC_90/Y 0.02fF
C563 INVX1_LOC_442/A INVX1_LOC_74/Y 0.08fF
C564 INVX1_LOC_6/Y NAND2X1_LOC_378/Y 0.01fF
C565 INVX1_LOC_312/A INVX1_LOC_245/A 0.01fF
C566 INVX1_LOC_674/A NAND2X1_LOC_853/a_36_24# 0.01fF
C567 INVX1_LOC_438/A INVX1_LOC_231/Y 0.02fF
C568 INVX1_LOC_614/A INVX1_LOC_662/A 0.07fF
C569 INVX1_LOC_361/Y INPUT_1 0.06fF
C570 INVX1_LOC_84/A NAND2X1_LOC_84/a_36_24# 0.00fF
C571 NAND2X1_LOC_190/A INVX1_LOC_387/Y 0.02fF
C572 NAND2X1_LOC_333/A INVX1_LOC_48/Y 0.13fF
C573 INVX1_LOC_11/Y NAND2X1_LOC_388/A 0.07fF
C574 INVX1_LOC_76/Y INVX1_LOC_62/Y 0.24fF
C575 INVX1_LOC_58/Y INVX1_LOC_252/Y 0.03fF
C576 INVX1_LOC_376/A INVX1_LOC_99/Y 0.46fF
C577 NAND2X1_LOC_307/A INVX1_LOC_119/Y 0.62fF
C578 NAND2X1_LOC_324/B INVX1_LOC_114/A 0.01fF
C579 INVX1_LOC_25/Y INPUT_5 0.00fF
C580 INVX1_LOC_48/Y INVX1_LOC_188/A 0.01fF
C581 INVX1_LOC_170/A INVX1_LOC_48/Y 0.00fF
C582 INVX1_LOC_379/A INVX1_LOC_26/Y 0.07fF
C583 INVX1_LOC_7/Y INVX1_LOC_422/A 0.12fF
C584 INVX1_LOC_502/A INVX1_LOC_99/Y 0.07fF
C585 NAND2X1_LOC_513/Y NAND2X1_LOC_417/a_36_24# 0.00fF
C586 INVX1_LOC_405/Y INVX1_LOC_145/Y 0.01fF
C587 INVX1_LOC_89/Y NAND2X1_LOC_753/Y 0.07fF
C588 INVX1_LOC_74/A INVX1_LOC_333/A 0.07fF
C589 INVX1_LOC_35/Y INVX1_LOC_26/Y 0.19fF
C590 NAND2X1_LOC_274/B INVX1_LOC_503/Y 0.01fF
C591 NAND2X1_LOC_27/a_36_24# INVX1_LOC_63/Y 0.00fF
C592 INVX1_LOC_183/Y NAND2X1_LOC_84/B 0.38fF
C593 INVX1_LOC_100/Y INVX1_LOC_116/Y 0.08fF
C594 INVX1_LOC_115/Y INVX1_LOC_41/Y 0.02fF
C595 INVX1_LOC_324/A NAND2X1_LOC_403/a_36_24# 0.00fF
C596 INVX1_LOC_77/A NAND2X1_LOC_615/B 0.04fF
C597 INVX1_LOC_627/A INVX1_LOC_133/Y 0.04fF
C598 INVX1_LOC_526/Y INVX1_LOC_74/Y 0.01fF
C599 INVX1_LOC_298/A NAND2X1_LOC_823/Y 0.01fF
C600 INVX1_LOC_488/A INVX1_LOC_48/Y 0.00fF
C601 INVX1_LOC_376/A INVX1_LOC_47/Y 0.08fF
C602 INVX1_LOC_49/Y INVX1_LOC_624/Y 0.01fF
C603 INVX1_LOC_41/Y INVX1_LOC_350/A 0.01fF
C604 INVX1_LOC_116/Y INVX1_LOC_74/Y 0.07fF
C605 INVX1_LOC_199/Y INVX1_LOC_89/A 0.03fF
C606 INVX1_LOC_93/Y INVX1_LOC_519/Y 0.03fF
C607 INVX1_LOC_26/Y NAND2X1_LOC_448/B 0.02fF
C608 INVX1_LOC_100/Y INVX1_LOC_328/A 0.02fF
C609 INVX1_LOC_26/Y INVX1_LOC_620/A 0.07fF
C610 INVX1_LOC_671/Y INVX1_LOC_655/A 0.00fF
C611 INVX1_LOC_405/Y INVX1_LOC_433/A 0.06fF
C612 NAND2X1_LOC_587/a_36_24# INVX1_LOC_74/A 0.00fF
C613 INVX1_LOC_371/A INVX1_LOC_666/Y 0.04fF
C614 INVX1_LOC_79/A INVX1_LOC_66/A 1.13fF
C615 INVX1_LOC_145/Y INVX1_LOC_620/Y 0.03fF
C616 INVX1_LOC_79/A INVX1_LOC_296/A 0.01fF
C617 INVX1_LOC_255/A INVX1_LOC_100/Y 0.02fF
C618 INVX1_LOC_361/A INVX1_LOC_90/Y 0.03fF
C619 INVX1_LOC_555/A NAND2X1_LOC_647/a_36_24# 0.01fF
C620 NAND2X1_LOC_267/A NAND2X1_LOC_71/a_36_24# 0.01fF
C621 INVX1_LOC_376/A INVX1_LOC_119/Y 0.07fF
C622 NAND2X1_LOC_239/a_36_24# INVX1_LOC_275/A 0.01fF
C623 INVX1_LOC_89/Y INVX1_LOC_652/Y 0.02fF
C624 INVX1_LOC_50/Y INVX1_LOC_91/Y 0.00fF
C625 INVX1_LOC_100/Y INVX1_LOC_179/A 0.03fF
C626 INVX1_LOC_31/Y INVX1_LOC_346/Y 0.01fF
C627 NAND2X1_LOC_274/B INVX1_LOC_242/Y 0.00fF
C628 INVX1_LOC_255/A INVX1_LOC_74/Y 0.07fF
C629 INVX1_LOC_100/A INVX1_LOC_223/A 0.18fF
C630 INVX1_LOC_223/Y INVX1_LOC_41/Y 0.32fF
C631 INVX1_LOC_424/A INVX1_LOC_404/Y 0.00fF
C632 INVX1_LOC_184/Y INVX1_LOC_9/Y 0.02fF
C633 VDD INVX1_LOC_629/Y 0.26fF
C634 INVX1_LOC_179/A INVX1_LOC_74/Y 0.01fF
C635 VDD INVX1_LOC_320/Y 0.21fF
C636 INVX1_LOC_200/Y INVX1_LOC_206/Y 0.01fF
C637 INVX1_LOC_63/Y NAND2X1_LOC_201/a_36_24# 0.00fF
C638 INVX1_LOC_69/Y INVX1_LOC_636/A 0.07fF
C639 INVX1_LOC_438/Y INVX1_LOC_450/A 0.03fF
C640 NAND2X1_LOC_69/a_36_24# INVX1_LOC_206/Y 0.00fF
C641 INPUT_0 INVX1_LOC_584/Y 0.02fF
C642 INVX1_LOC_482/Y INVX1_LOC_485/A -0.00fF
C643 INVX1_LOC_627/A INVX1_LOC_581/A 0.06fF
C644 INVX1_LOC_133/Y INVX1_LOC_581/A 0.02fF
C645 INVX1_LOC_426/A INVX1_LOC_596/A 0.17fF
C646 INVX1_LOC_174/Y INVX1_LOC_190/Y 0.09fF
C647 INVX1_LOC_224/Y NAND2X1_LOC_180/B 0.03fF
C648 NAND2X1_LOC_795/a_36_24# INVX1_LOC_615/A 0.00fF
C649 INVX1_LOC_202/A INVX1_LOC_12/Y 0.01fF
C650 INVX1_LOC_435/Y INVX1_LOC_51/Y 0.05fF
C651 VDD INPUT_7 0.08fF
C652 INVX1_LOC_618/A INVX1_LOC_98/Y 0.05fF
C653 VDD INVX1_LOC_659/Y -0.00fF
C654 NAND2X1_LOC_322/Y NAND2X1_LOC_325/B 0.10fF
C655 INVX1_LOC_578/A NAND2X1_LOC_180/B 0.05fF
C656 NAND2X1_LOC_475/A NAND2X1_LOC_307/A 0.04fF
C657 INVX1_LOC_99/Y INVX1_LOC_388/Y 0.00fF
C658 INVX1_LOC_224/Y INVX1_LOC_188/Y 0.08fF
C659 NAND2X1_LOC_208/a_36_24# INVX1_LOC_366/A 0.01fF
C660 NAND2X1_LOC_249/Y INVX1_LOC_35/Y 0.47fF
C661 VDD INVX1_LOC_679/A 0.00fF
C662 NAND2X1_LOC_45/Y INVX1_LOC_17/Y 0.27fF
C663 NAND2X1_LOC_767/a_36_24# INVX1_LOC_366/A 0.00fF
C664 INVX1_LOC_438/A INVX1_LOC_367/Y 0.01fF
C665 INVX1_LOC_596/A INVX1_LOC_51/Y 0.07fF
C666 INVX1_LOC_53/Y INVX1_LOC_185/Y 0.02fF
C667 INPUT_0 INVX1_LOC_274/A 0.01fF
C668 INVX1_LOC_366/A NAND2X1_LOC_240/a_36_24# 0.00fF
C669 INVX1_LOC_53/Y INVX1_LOC_45/Y 0.44fF
C670 INVX1_LOC_20/Y NAND2X1_LOC_342/a_36_24# 0.00fF
C671 INVX1_LOC_625/A INVX1_LOC_395/A 0.09fF
C672 INVX1_LOC_257/Y INVX1_LOC_352/Y 0.07fF
C673 INVX1_LOC_298/Y INVX1_LOC_299/A 0.01fF
C674 NAND2X1_LOC_467/A INVX1_LOC_522/Y 0.01fF
C675 NAND2X1_LOC_788/A INVX1_LOC_350/Y 0.01fF
C676 NAND2X1_LOC_498/Y INVX1_LOC_503/A 0.03fF
C677 INPUT_0 INVX1_LOC_209/A 0.00fF
C678 INVX1_LOC_560/A INVX1_LOC_35/Y 0.33fF
C679 VDD INVX1_LOC_571/A -0.00fF
C680 INVX1_LOC_31/Y NAND2X1_LOC_76/B 0.14fF
C681 NAND2X1_LOC_791/B INVX1_LOC_272/Y 0.07fF
C682 VDD INVX1_LOC_542/Y 0.22fF
C683 INVX1_LOC_597/A INVX1_LOC_366/A 0.27fF
C684 INVX1_LOC_666/A INVX1_LOC_600/A 0.04fF
C685 INVX1_LOC_424/Y INVX1_LOC_439/A 0.00fF
C686 INVX1_LOC_551/Y INVX1_LOC_134/Y 0.10fF
C687 INVX1_LOC_412/Y INVX1_LOC_354/Y 0.01fF
C688 INVX1_LOC_51/Y INVX1_LOC_504/A 0.07fF
C689 INVX1_LOC_384/A INVX1_LOC_377/A 0.03fF
C690 INVX1_LOC_578/A NAND2X1_LOC_444/a_36_24# 0.01fF
C691 INPUT_3 INVX1_LOC_53/Y 0.03fF
C692 INVX1_LOC_400/A INVX1_LOC_65/Y 0.07fF
C693 INVX1_LOC_393/Y INVX1_LOC_50/Y 0.01fF
C694 INVX1_LOC_218/A INVX1_LOC_386/Y 0.03fF
C695 INVX1_LOC_384/A NAND2X1_LOC_595/Y 0.02fF
C696 NAND2X1_LOC_781/B INVX1_LOC_168/Y 0.04fF
C697 VDD NAND2X1_LOC_258/Y 0.05fF
C698 INVX1_LOC_17/Y INVX1_LOC_114/Y 0.01fF
C699 INVX1_LOC_255/Y INVX1_LOC_360/A 0.00fF
C700 INVX1_LOC_395/A INVX1_LOC_208/Y 0.02fF
C701 INVX1_LOC_268/A INVX1_LOC_566/A 0.27fF
C702 INVX1_LOC_406/Y INVX1_LOC_385/Y 0.03fF
C703 INVX1_LOC_62/Y INVX1_LOC_192/A 0.04fF
C704 NAND2X1_LOC_324/B NAND2X1_LOC_321/a_36_24# 0.00fF
C705 NAND2X1_LOC_13/Y INVX1_LOC_98/Y 0.01fF
C706 INVX1_LOC_442/A INVX1_LOC_350/Y -0.05fF
C707 INVX1_LOC_21/Y INVX1_LOC_324/A 0.01fF
C708 INVX1_LOC_288/Y INVX1_LOC_686/A 0.04fF
C709 INVX1_LOC_404/Y INVX1_LOC_49/Y 0.03fF
C710 INVX1_LOC_65/Y INVX1_LOC_93/Y 0.03fF
C711 INVX1_LOC_626/A NAND2X1_LOC_513/A 0.01fF
C712 INVX1_LOC_448/A INVX1_LOC_377/A 0.11fF
C713 INVX1_LOC_402/Y INVX1_LOC_670/Y 0.18fF
C714 INVX1_LOC_448/A NAND2X1_LOC_595/Y 0.03fF
C715 NAND2X1_LOC_315/a_36_24# NAND2X1_LOC_267/A 0.01fF
C716 INVX1_LOC_35/Y INVX1_LOC_369/A 0.06fF
C717 INVX1_LOC_605/Y INVX1_LOC_492/A 0.01fF
C718 INPUT_0 INVX1_LOC_328/Y 8.73fF
C719 NAND2X1_LOC_788/A INVX1_LOC_79/A 0.37fF
C720 VDD NAND2X1_LOC_545/A 0.01fF
C721 INVX1_LOC_366/A INVX1_LOC_6/Y 0.02fF
C722 INVX1_LOC_341/Y INVX1_LOC_55/Y 0.09fF
C723 INVX1_LOC_45/Y NAND2X1_LOC_274/Y 0.00fF
C724 INPUT_0 INVX1_LOC_518/A 0.03fF
C725 INVX1_LOC_608/Y INVX1_LOC_99/Y 0.01fF
C726 INVX1_LOC_447/Y NAND2X1_LOC_179/Y 0.06fF
C727 INVX1_LOC_201/Y INVX1_LOC_205/Y 0.00fF
C728 NAND2X1_LOC_673/A INVX1_LOC_600/A 0.01fF
C729 INVX1_LOC_201/A INVX1_LOC_274/A 0.02fF
C730 INVX1_LOC_17/Y INVX1_LOC_99/Y 1.60fF
C731 INVX1_LOC_80/A INVX1_LOC_117/Y 0.25fF
C732 VDD INVX1_LOC_653/Y 0.76fF
C733 INVX1_LOC_438/Y NAND2X1_LOC_631/B 0.05fF
C734 NAND2X1_LOC_768/A INVX1_LOC_117/Y 0.02fF
C735 INVX1_LOC_459/A INVX1_LOC_348/Y 0.09fF
C736 NAND2X1_LOC_516/Y INVX1_LOC_518/A 0.00fF
C737 INVX1_LOC_8/Y INVX1_LOC_7/Y 0.02fF
C738 NAND2X1_LOC_669/Y INVX1_LOC_298/A 0.01fF
C739 INVX1_LOC_91/Y INVX1_LOC_275/A 0.05fF
C740 INVX1_LOC_20/Y NAND2X1_LOC_537/a_36_24# 0.00fF
C741 VDD INVX1_LOC_327/A 0.00fF
C742 INVX1_LOC_6/Y INVX1_LOC_486/Y 0.01fF
C743 NAND2X1_LOC_318/B INVX1_LOC_254/A 0.09fF
C744 VDD INVX1_LOC_666/Y 0.54fF
C745 INVX1_LOC_271/A INVX1_LOC_153/Y 0.54fF
C746 INVX1_LOC_89/Y INVX1_LOC_197/A 0.01fF
C747 INVX1_LOC_400/A INVX1_LOC_479/Y 0.01fF
C748 INVX1_LOC_421/A INVX1_LOC_232/Y 0.03fF
C749 INVX1_LOC_442/Y INPUT_1 0.07fF
C750 INVX1_LOC_442/A INVX1_LOC_79/A 0.07fF
C751 INVX1_LOC_524/Y INVX1_LOC_95/A 0.02fF
C752 INVX1_LOC_53/Y NAND2X1_LOC_837/A 0.02fF
C753 INVX1_LOC_139/A INVX1_LOC_62/Y 0.02fF
C754 NAND2X1_LOC_615/B INVX1_LOC_59/Y 1.14fF
C755 INVX1_LOC_446/Y INVX1_LOC_280/A 0.07fF
C756 NAND2X1_LOC_93/Y INVX1_LOC_91/Y 0.01fF
C757 INVX1_LOC_277/A NAND2X1_LOC_106/B 0.00fF
C758 INVX1_LOC_116/Y INVX1_LOC_350/Y -0.00fF
C759 INVX1_LOC_597/A INVX1_LOC_6/Y 0.01fF
C760 INVX1_LOC_523/A INVX1_LOC_135/Y 0.05fF
C761 INVX1_LOC_400/A INVX1_LOC_318/A 0.02fF
C762 NAND2X1_LOC_538/B INVX1_LOC_242/Y 0.08fF
C763 INVX1_LOC_502/Y INVX1_LOC_502/A 0.08fF
C764 INVX1_LOC_451/A INVX1_LOC_46/Y 0.46fF
C765 INVX1_LOC_20/Y NAND2X1_LOC_274/B 0.03fF
C766 NAND2X1_LOC_615/B INVX1_LOC_48/Y 0.15fF
C767 INVX1_LOC_11/Y INVX1_LOC_117/Y 0.26fF
C768 INVX1_LOC_306/Y INVX1_LOC_7/Y 0.03fF
C769 INVX1_LOC_602/A INVX1_LOC_50/A 0.03fF
C770 NAND2X1_LOC_342/a_36_24# INVX1_LOC_655/A 0.01fF
C771 INVX1_LOC_164/Y INVX1_LOC_50/Y 0.03fF
C772 INVX1_LOC_32/Y INVX1_LOC_303/Y 0.00fF
C773 INVX1_LOC_206/Y NAND2X1_LOC_237/a_36_24# 0.01fF
C774 INVX1_LOC_50/Y NAND2X1_LOC_333/B 0.11fF
C775 INVX1_LOC_361/Y INVX1_LOC_50/Y 0.08fF
C776 INVX1_LOC_17/Y INVX1_LOC_47/Y 0.17fF
C777 INVX1_LOC_12/Y NAND2X1_LOC_615/Y 0.39fF
C778 NAND2X1_LOC_123/A INVX1_LOC_347/Y 0.03fF
C779 INVX1_LOC_585/Y INVX1_LOC_173/Y 0.04fF
C780 INVX1_LOC_17/Y NAND2X1_LOC_557/B 0.00fF
C781 INVX1_LOC_297/A INVX1_LOC_245/A 0.01fF
C782 INVX1_LOC_281/A INVX1_LOC_50/Y 0.24fF
C783 INVX1_LOC_300/A NAND2X1_LOC_212/a_36_24# 0.00fF
C784 INVX1_LOC_340/Y INVX1_LOC_479/A 0.02fF
C785 NAND2X1_LOC_649/a_36_24# INVX1_LOC_66/A 0.01fF
C786 INVX1_LOC_384/A NAND2X1_LOC_372/Y 0.07fF
C787 INVX1_LOC_54/Y NAND2X1_LOC_128/A 0.37fF
C788 INVX1_LOC_383/A INVX1_LOC_666/Y 0.04fF
C789 INVX1_LOC_361/A INVX1_LOC_98/Y 0.15fF
C790 NAND2X1_LOC_111/Y NAND2X1_LOC_775/B 0.33fF
C791 NAND2X1_LOC_299/Y INVX1_LOC_114/A 0.00fF
C792 NAND2X1_LOC_399/B INVX1_LOC_9/Y 0.11fF
C793 NAND2X1_LOC_673/B INVX1_LOC_199/Y 0.21fF
C794 INVX1_LOC_7/Y INVX1_LOC_9/Y 4.04fF
C795 INVX1_LOC_201/Y INVX1_LOC_44/Y 0.02fF
C796 INVX1_LOC_261/Y INVX1_LOC_50/Y 0.03fF
C797 INVX1_LOC_49/Y INVX1_LOC_480/Y 0.06fF
C798 INVX1_LOC_69/Y NAND2X1_LOC_720/A 0.03fF
C799 INPUT_3 INVX1_LOC_368/Y 0.01fF
C800 INVX1_LOC_48/Y INVX1_LOC_296/A 0.01fF
C801 INVX1_LOC_47/Y NAND2X1_LOC_435/a_36_24# 0.00fF
C802 INVX1_LOC_155/A INVX1_LOC_32/Y 0.01fF
C803 INVX1_LOC_411/A INVX1_LOC_411/Y 0.01fF
C804 INVX1_LOC_412/A INVX1_LOC_92/A 0.01fF
C805 NAND2X1_LOC_710/A INVX1_LOC_479/A 0.00fF
C806 INVX1_LOC_12/A INVX1_LOC_13/Y 0.01fF
C807 NAND2X1_LOC_822/Y INVX1_LOC_659/A 0.03fF
C808 INVX1_LOC_268/A INVX1_LOC_79/A 0.30fF
C809 INVX1_LOC_79/A INVX1_LOC_116/Y 0.03fF
C810 INVX1_LOC_17/Y INVX1_LOC_119/Y 0.28fF
C811 INVX1_LOC_184/A INVX1_LOC_86/A 0.08fF
C812 INVX1_LOC_49/Y INVX1_LOC_169/Y 0.03fF
C813 INVX1_LOC_31/Y NAND2X1_LOC_52/Y 0.11fF
C814 NAND2X1_LOC_837/B INVX1_LOC_26/Y 0.01fF
C815 INVX1_LOC_543/Y INVX1_LOC_44/Y 0.02fF
C816 INVX1_LOC_17/Y NAND2X1_LOC_66/Y 0.01fF
C817 INVX1_LOC_93/Y INVX1_LOC_95/A 0.00fF
C818 NAND2X1_LOC_307/B INVX1_LOC_47/Y 0.01fF
C819 INVX1_LOC_35/Y NAND2X1_LOC_626/Y 0.03fF
C820 INVX1_LOC_586/A INVX1_LOC_636/A 0.00fF
C821 INVX1_LOC_159/Y INVX1_LOC_242/Y 0.16fF
C822 INVX1_LOC_502/A NAND2X1_LOC_276/a_36_24# 0.01fF
C823 INVX1_LOC_448/A NAND2X1_LOC_372/Y 0.12fF
C824 INVX1_LOC_145/Y INVX1_LOC_280/A 0.03fF
C825 INVX1_LOC_32/Y INVX1_LOC_9/Y 0.21fF
C826 INVX1_LOC_555/A INVX1_LOC_507/Y 0.00fF
C827 INVX1_LOC_439/Y INVX1_LOC_430/Y 0.14fF
C828 INVX1_LOC_79/A NAND2X1_LOC_432/Y 0.01fF
C829 INVX1_LOC_256/A INVX1_LOC_62/Y 0.06fF
C830 INVX1_LOC_208/A INVX1_LOC_26/Y 0.15fF
C831 INVX1_LOC_42/Y INVX1_LOC_184/Y 0.01fF
C832 INVX1_LOC_44/Y NAND2X1_LOC_753/Y 0.05fF
C833 INVX1_LOC_62/Y NAND2X1_LOC_259/A 0.00fF
C834 INVX1_LOC_13/Y INVX1_LOC_7/Y 0.02fF
C835 INVX1_LOC_145/Y NAND2X1_LOC_372/Y 0.00fF
C836 INVX1_LOC_41/Y NAND2X1_LOC_606/Y 0.01fF
C837 INVX1_LOC_300/Y INVX1_LOC_69/Y 0.03fF
C838 INVX1_LOC_274/A INVX1_LOC_211/A 0.23fF
C839 INVX1_LOC_431/A NAND2X1_LOC_488/Y 0.11fF
C840 NAND2X1_LOC_336/B INVX1_LOC_92/A 0.30fF
C841 INVX1_LOC_54/Y INVX1_LOC_66/Y 0.09fF
C842 INVX1_LOC_54/Y NAND2X1_LOC_248/B 0.00fF
C843 NAND2X1_LOC_307/B INVX1_LOC_119/Y 0.00fF
C844 INVX1_LOC_32/Y INVX1_LOC_62/Y 0.29fF
C845 INVX1_LOC_69/Y INVX1_LOC_100/Y 2.25fF
C846 INVX1_LOC_255/A INVX1_LOC_79/A 0.07fF
C847 INVX1_LOC_93/Y INVX1_LOC_588/A 0.06fF
C848 NAND2X1_LOC_486/A INVX1_LOC_479/A 0.00fF
C849 INVX1_LOC_69/Y INVX1_LOC_74/Y 1.08fF
C850 INVX1_LOC_69/Y INVX1_LOC_660/A 0.13fF
C851 INVX1_LOC_519/Y INVX1_LOC_128/A 0.01fF
C852 NAND2X1_LOC_388/A INVX1_LOC_625/Y 0.02fF
C853 VDD INVX1_LOC_490/Y 0.28fF
C854 INVX1_LOC_58/Y NAND2X1_LOC_231/B 0.33fF
C855 INVX1_LOC_100/Y INVX1_LOC_667/A 0.01fF
C856 INVX1_LOC_63/Y NAND2X1_LOC_227/A 0.02fF
C857 VDD NAND2X1_LOC_16/Y -0.00fF
C858 NAND2X1_LOC_164/Y INVX1_LOC_395/A 0.12fF
C859 VDD INVX1_LOC_299/Y 0.21fF
C860 VDD INVX1_LOC_353/Y 0.05fF
C861 INVX1_LOC_291/Y INVX1_LOC_90/Y 0.03fF
C862 INVX1_LOC_584/A NAND2X1_LOC_122/Y 0.01fF
C863 INPUT_6 INVX1_LOC_334/Y 0.01fF
C864 INVX1_LOC_395/A INVX1_LOC_65/Y 0.01fF
C865 INPUT_0 INVX1_LOC_266/Y 0.00fF
C866 VDD INVX1_LOC_55/Y 0.76fF
C867 NAND2X1_LOC_475/A INVX1_LOC_286/Y 0.00fF
C868 INVX1_LOC_206/Y NAND2X1_LOC_180/B 0.00fF
C869 INVX1_LOC_404/Y INVX1_LOC_76/Y 0.02fF
C870 NAND2X1_LOC_331/A INVX1_LOC_76/Y 0.75fF
C871 INVX1_LOC_269/Y INVX1_LOC_586/A 0.03fF
C872 VDD NAND2X1_LOC_829/Y 0.19fF
C873 INVX1_LOC_115/A INVX1_LOC_638/A 0.12fF
C874 VDD INVX1_LOC_97/Y 0.46fF
C875 NAND2X1_LOC_45/a_36_24# INVX1_LOC_449/A 0.00fF
C876 INVX1_LOC_21/Y INVX1_LOC_447/A 0.06fF
C877 INVX1_LOC_603/Y INVX1_LOC_206/Y 0.07fF
C878 NAND2X1_LOC_249/Y INVX1_LOC_214/Y 0.01fF
C879 NAND2X1_LOC_787/a_36_24# NAND2X1_LOC_249/Y 0.00fF
C880 INVX1_LOC_257/Y INVX1_LOC_67/Y 0.02fF
C881 INVX1_LOC_418/Y INVX1_LOC_301/A 0.03fF
C882 INVX1_LOC_424/A INVX1_LOC_451/A 0.03fF
C883 INVX1_LOC_381/A INVX1_LOC_586/A 0.10fF
C884 INVX1_LOC_202/A NAND2X1_LOC_615/B 0.01fF
C885 NAND2X1_LOC_333/B INVX1_LOC_275/A 0.02fF
C886 INVX1_LOC_20/Y INVX1_LOC_38/A 0.05fF
C887 VDD INVX1_LOC_391/Y 0.14fF
C888 INVX1_LOC_434/A INVX1_LOC_444/Y 0.03fF
C889 INVX1_LOC_449/Y INVX1_LOC_453/A 0.01fF
C890 NAND2X1_LOC_164/Y INVX1_LOC_284/A 0.14fF
C891 INVX1_LOC_17/Y NAND2X1_LOC_475/A 0.11fF
C892 INVX1_LOC_604/Y INVX1_LOC_395/A 0.54fF
C893 INVX1_LOC_418/A INVX1_LOC_134/Y 0.01fF
C894 VDD INVX1_LOC_431/A -0.00fF
C895 NAND2X1_LOC_249/Y INVX1_LOC_118/A 0.07fF
C896 INVX1_LOC_84/A NAND2X1_LOC_391/B 0.19fF
C897 INVX1_LOC_206/Y INVX1_LOC_478/Y 0.00fF
C898 NAND2X1_LOC_790/B INVX1_LOC_620/A 0.03fF
C899 NAND2X1_LOC_180/B INVX1_LOC_686/A 0.01fF
C900 NAND2X1_LOC_93/Y NAND2X1_LOC_333/B -0.03fF
C901 NAND2X1_LOC_56/Y INVX1_LOC_666/A 0.30fF
C902 INVX1_LOC_239/Y INVX1_LOC_239/A 0.10fF
C903 INVX1_LOC_551/Y INVX1_LOC_318/Y 0.15fF
C904 INVX1_LOC_137/A NAND2X1_LOC_610/a_36_24# 0.00fF
C905 INVX1_LOC_584/Y INVX1_LOC_145/Y 0.31fF
C906 INVX1_LOC_355/A INVX1_LOC_504/A 0.01fF
C907 INVX1_LOC_54/Y INVX1_LOC_412/Y 0.11fF
C908 VDD INVX1_LOC_18/Y 0.37fF
C909 INVX1_LOC_49/Y INVX1_LOC_638/A 0.07fF
C910 INVX1_LOC_449/A INVX1_LOC_384/A 1.56fF
C911 NAND2X1_LOC_332/B INVX1_LOC_377/A 0.01fF
C912 INVX1_LOC_238/Y INVX1_LOC_46/Y 0.03fF
C913 INVX1_LOC_206/Y NAND2X1_LOC_387/Y 0.11fF
C914 NAND2X1_LOC_768/a_36_24# INVX1_LOC_596/A 0.02fF
C915 INVX1_LOC_373/A NAND2X1_LOC_634/a_36_24# 0.00fF
C916 INVX1_LOC_412/Y NAND2X1_LOC_173/a_36_24# 0.00fF
C917 INVX1_LOC_293/Y INVX1_LOC_53/Y 0.03fF
C918 INVX1_LOC_166/A NAND2X1_LOC_317/B 0.01fF
C919 INVX1_LOC_412/A INPUT_1 0.08fF
C920 VDD INVX1_LOC_94/Y 0.30fF
C921 INVX1_LOC_17/Y INVX1_LOC_502/Y 0.01fF
C922 INVX1_LOC_686/A INVX1_LOC_188/Y 0.07fF
C923 INVX1_LOC_213/Y INVX1_LOC_45/Y 0.03fF
C924 NAND2X1_LOC_184/Y INVX1_LOC_547/Y 0.07fF
C925 INVX1_LOC_407/Y INVX1_LOC_76/Y 0.01fF
C926 INVX1_LOC_412/Y INVX1_LOC_257/A 0.24fF
C927 NAND2X1_LOC_242/A INVX1_LOC_69/Y 0.26fF
C928 INVX1_LOC_547/A NAND2X1_LOC_259/A 0.15fF
C929 INVX1_LOC_661/A NAND2X1_LOC_260/Y 0.03fF
C930 INVX1_LOC_456/Y INVX1_LOC_55/Y 0.01fF
C931 INVX1_LOC_379/A INVX1_LOC_235/Y 0.14fF
C932 NAND2X1_LOC_32/a_36_24# INVX1_LOC_43/A 0.00fF
C933 INVX1_LOC_586/A NAND2X1_LOC_720/A 1.27fF
C934 INVX1_LOC_210/Y NAND2X1_LOC_79/Y 0.12fF
C935 INVX1_LOC_448/A INVX1_LOC_449/A 0.05fF
C936 INVX1_LOC_35/Y INVX1_LOC_235/Y 0.03fF
C937 INVX1_LOC_63/A INVX1_LOC_145/Y 0.01fF
C938 INVX1_LOC_20/Y INVX1_LOC_159/Y 0.03fF
C939 INVX1_LOC_51/Y INVX1_LOC_520/A 0.01fF
C940 NAND2X1_LOC_513/Y INVX1_LOC_66/A 0.08fF
C941 NAND2X1_LOC_592/B INVX1_LOC_47/Y 0.04fF
C942 INVX1_LOC_617/Y NAND2X1_LOC_602/A 0.03fF
C943 INVX1_LOC_257/Y INVX1_LOC_347/Y 0.02fF
C944 INVX1_LOC_65/Y INVX1_LOC_31/Y 0.20fF
C945 INVX1_LOC_317/Y INVX1_LOC_317/A 0.03fF
C946 NAND2X1_LOC_387/Y INVX1_LOC_396/Y 0.71fF
C947 INVX1_LOC_449/A INVX1_LOC_145/Y 0.04fF
C948 INVX1_LOC_395/A INVX1_LOC_95/A 0.01fF
C949 INVX1_LOC_295/A INVX1_LOC_304/Y 0.01fF
C950 NAND2X1_LOC_186/a_36_24# INVX1_LOC_76/Y 0.01fF
C951 INVX1_LOC_196/A INVX1_LOC_48/Y 0.01fF
C952 INVX1_LOC_670/Y INVX1_LOC_669/Y 0.00fF
C953 INVX1_LOC_546/Y INVX1_LOC_63/Y 0.02fF
C954 INVX1_LOC_206/Y INVX1_LOC_491/A 0.07fF
C955 INVX1_LOC_80/A NAND2X1_LOC_76/A 0.01fF
C956 INVX1_LOC_17/Y NAND2X1_LOC_38/a_36_24# 0.00fF
C957 INVX1_LOC_371/Y INVX1_LOC_510/A 0.01fF
C958 NAND2X1_LOC_698/Y INVX1_LOC_45/Y 0.01fF
C959 INVX1_LOC_542/A INVX1_LOC_513/Y 0.03fF
C960 INVX1_LOC_131/Y NAND2X1_LOC_342/A 0.02fF
C961 INVX1_LOC_288/A INVX1_LOC_347/Y 0.35fF
C962 NAND2X1_LOC_336/B INPUT_1 0.00fF
C963 INVX1_LOC_42/Y INVX1_LOC_7/Y 0.10fF
C964 NAND2X1_LOC_595/Y INVX1_LOC_503/Y 0.18fF
C965 INVX1_LOC_468/Y INVX1_LOC_504/Y 0.03fF
C966 INVX1_LOC_307/A INVX1_LOC_50/Y 0.01fF
C967 NAND2X1_LOC_537/B INVX1_LOC_100/Y 0.04fF
C968 INVX1_LOC_555/A INVX1_LOC_522/Y 0.04fF
C969 INVX1_LOC_511/Y INVX1_LOC_137/Y 0.14fF
C970 INVX1_LOC_17/Y NAND2X1_LOC_43/Y 0.04fF
C971 INVX1_LOC_566/A INVX1_LOC_69/Y 0.07fF
C972 INVX1_LOC_166/A INVX1_LOC_633/Y 0.34fF
C973 INVX1_LOC_134/Y INVX1_LOC_46/Y 6.08fF
C974 INVX1_LOC_300/Y INVX1_LOC_586/A 0.09fF
C975 INVX1_LOC_89/Y INVX1_LOC_336/Y 0.01fF
C976 NAND2X1_LOC_592/B INVX1_LOC_119/Y 0.23fF
C977 INVX1_LOC_93/Y INVX1_LOC_670/Y 0.07fF
C978 INVX1_LOC_556/Y INVX1_LOC_35/Y 0.03fF
C979 INVX1_LOC_406/Y INVX1_LOC_420/A 0.08fF
C980 INVX1_LOC_11/Y INVX1_LOC_178/A 0.00fF
C981 INVX1_LOC_11/Y INVX1_LOC_251/Y 0.50fF
C982 NAND2X1_LOC_548/B NAND2X1_LOC_531/Y 0.02fF
C983 INVX1_LOC_442/Y INVX1_LOC_50/Y 0.07fF
C984 INVX1_LOC_45/Y INVX1_LOC_653/A 0.01fF
C985 INVX1_LOC_47/A INVX1_LOC_46/Y 0.02fF
C986 NAND2X1_LOC_520/B INVX1_LOC_502/A 0.03fF
C987 NAND2X1_LOC_697/Y INVX1_LOC_550/A 0.05fF
C988 INVX1_LOC_145/Y INVX1_LOC_186/Y 0.26fF
C989 NAND2X1_LOC_97/B INVX1_LOC_89/Y 0.09fF
C990 NAND2X1_LOC_457/A INVX1_LOC_75/Y 0.10fF
C991 INVX1_LOC_51/Y INVX1_LOC_519/Y 0.05fF
C992 NAND2X1_LOC_781/B NAND2X1_LOC_781/a_36_24# 0.00fF
C993 INVX1_LOC_47/Y NAND2X1_LOC_616/Y 0.07fF
C994 INVX1_LOC_456/Y INVX1_LOC_18/Y 0.02fF
C995 INVX1_LOC_80/A INVX1_LOC_58/Y 8.16fF
C996 INVX1_LOC_586/A INVX1_LOC_100/Y 0.25fF
C997 INVX1_LOC_511/Y NAND2X1_LOC_829/B 0.08fF
C998 NAND2X1_LOC_690/Y INVX1_LOC_41/Y 0.01fF
C999 NAND2X1_LOC_768/A INVX1_LOC_58/Y 0.01fF
C1000 INVX1_LOC_607/Y GATE_662 0.04fF
C1001 INVX1_LOC_11/Y INVX1_LOC_608/A 0.06fF
C1002 INVX1_LOC_417/Y INVX1_LOC_255/A 0.10fF
C1003 INVX1_LOC_166/A NAND2X1_LOC_308/a_36_24# 0.00fF
C1004 INVX1_LOC_551/Y INVX1_LOC_90/Y 0.03fF
C1005 INVX1_LOC_155/Y INVX1_LOC_188/A 0.01fF
C1006 INVX1_LOC_507/Y INVX1_LOC_474/Y 0.03fF
C1007 INVX1_LOC_335/A INVX1_LOC_498/A 0.05fF
C1008 INVX1_LOC_531/Y INVX1_LOC_169/A 0.00fF
C1009 INVX1_LOC_586/A INVX1_LOC_74/Y 0.14fF
C1010 INVX1_LOC_89/Y INVX1_LOC_440/Y 0.28fF
C1011 INVX1_LOC_166/A NAND2X1_LOC_119/a_36_24# 0.00fF
C1012 INVX1_LOC_415/Y INVX1_LOC_6/Y 0.01fF
C1013 NAND2X1_LOC_457/A NAND2X1_LOC_271/A 0.02fF
C1014 INVX1_LOC_312/Y INVX1_LOC_100/Y 0.03fF
C1015 INVX1_LOC_266/Y INVX1_LOC_211/A 0.07fF
C1016 NAND2X1_LOC_274/B INVX1_LOC_375/Y 0.01fF
C1017 NAND2X1_LOC_32/Y INVX1_LOC_6/Y 0.01fF
C1018 INVX1_LOC_318/A INVX1_LOC_31/Y 0.09fF
C1019 INVX1_LOC_361/Y NAND2X1_LOC_388/A 1.49fF
C1020 INVX1_LOC_11/Y INVX1_LOC_58/Y 0.29fF
C1021 INVX1_LOC_80/A NAND2X1_LOC_342/B 0.01fF
C1022 INVX1_LOC_255/A INVX1_LOC_48/Y 0.03fF
C1023 INVX1_LOC_397/A NAND2X1_LOC_237/a_36_24# 0.00fF
C1024 NAND2X1_LOC_825/a_36_24# NAND2X1_LOC_720/A 0.00fF
C1025 INVX1_LOC_47/Y INVX1_LOC_497/Y 0.14fF
C1026 INVX1_LOC_328/Y INVX1_LOC_145/Y 0.03fF
C1027 NAND2X1_LOC_140/B NAND2X1_LOC_274/B 0.03fF
C1028 INVX1_LOC_49/Y INVX1_LOC_665/Y 0.10fF
C1029 INVX1_LOC_179/A INVX1_LOC_59/Y 0.01fF
C1030 INVX1_LOC_682/Y INVX1_LOC_370/A 0.17fF
C1031 NAND2X1_LOC_708/A INVX1_LOC_168/Y 0.01fF
C1032 INVX1_LOC_93/Y INVX1_LOC_253/Y 0.01fF
C1033 INVX1_LOC_469/Y INVX1_LOC_69/Y 0.05fF
C1034 INVX1_LOC_277/Y INVX1_LOC_662/Y 0.07fF
C1035 INVX1_LOC_6/Y NAND2X1_LOC_294/Y 14.21fF
C1036 INVX1_LOC_35/Y NAND2X1_LOC_420/Y 0.06fF
C1037 INVX1_LOC_47/Y INVX1_LOC_230/Y 0.03fF
C1038 NAND2X1_LOC_324/B INVX1_LOC_62/Y 0.04fF
C1039 INPUT_1 NAND2X1_LOC_847/A 0.09fF
C1040 INVX1_LOC_137/Y NAND2X1_LOC_780/a_36_24# 0.00fF
C1041 INVX1_LOC_93/Y INVX1_LOC_63/Y 1.49fF
C1042 INVX1_LOC_145/Y INVX1_LOC_207/Y 0.31fF
C1043 NAND2X1_LOC_181/A INVX1_LOC_69/Y 0.02fF
C1044 INVX1_LOC_360/A NAND2X1_LOC_605/B 0.35fF
C1045 INVX1_LOC_17/Y NAND2X1_LOC_627/Y 0.02fF
C1046 INVX1_LOC_555/A INVX1_LOC_508/A 0.02fF
C1047 INVX1_LOC_31/Y INVX1_LOC_314/Y 0.01fF
C1048 INVX1_LOC_471/Y INVX1_LOC_50/Y 0.01fF
C1049 INVX1_LOC_543/A INVX1_LOC_86/Y 0.01fF
C1050 NAND2X1_LOC_775/B INVX1_LOC_41/Y 2.23fF
C1051 INVX1_LOC_657/Y INVX1_LOC_656/Y 0.20fF
C1052 INVX1_LOC_117/Y INVX1_LOC_319/A 0.03fF
C1053 NAND2X1_LOC_121/Y INVX1_LOC_497/A 0.05fF
C1054 INVX1_LOC_581/A INVX1_LOC_613/A 0.06fF
C1055 INPUT_0 INVX1_LOC_109/Y 0.03fF
C1056 INVX1_LOC_390/A INVX1_LOC_63/Y 0.04fF
C1057 INVX1_LOC_277/A NAND2X1_LOC_248/B 0.18fF
C1058 INVX1_LOC_117/Y NAND2X1_LOC_843/B 0.01fF
C1059 INVX1_LOC_105/A INVX1_LOC_666/Y 0.02fF
C1060 INVX1_LOC_69/Y INVX1_LOC_79/A 0.23fF
C1061 INVX1_LOC_486/A INVX1_LOC_90/Y 0.01fF
C1062 NAND2X1_LOC_637/A NAND2X1_LOC_591/B 0.20fF
C1063 NAND2X1_LOC_835/A INVX1_LOC_74/Y 0.02fF
C1064 INVX1_LOC_31/Y INVX1_LOC_588/A -0.03fF
C1065 INVX1_LOC_117/Y INVX1_LOC_91/Y 0.03fF
C1066 INPUT_0 INVX1_LOC_554/A 0.00fF
C1067 VDD INVX1_LOC_54/A 0.00fF
C1068 NAND2X1_LOC_108/a_36_24# NAND2X1_LOC_248/B 0.00fF
C1069 INVX1_LOC_491/A NAND2X1_LOC_609/B 0.07fF
C1070 INVX1_LOC_206/Y NAND2X1_LOC_180/a_36_24# 0.00fF
C1071 INVX1_LOC_193/Y INVX1_LOC_410/Y 0.17fF
C1072 NAND2X1_LOC_331/A INVX1_LOC_139/A 0.00fF
C1073 NAND2X1_LOC_799/a_36_24# NAND2X1_LOC_173/Y 0.00fF
C1074 NAND2X1_LOC_790/B INVX1_LOC_291/A 0.01fF
C1075 INVX1_LOC_241/A INVX1_LOC_669/A 0.04fF
C1076 NAND2X1_LOC_242/A INVX1_LOC_586/A 0.02fF
C1077 VDD INVX1_LOC_677/Y 0.36fF
C1078 INVX1_LOC_588/A INVX1_LOC_473/Y 0.10fF
C1079 NAND2X1_LOC_544/B INVX1_LOC_66/Y 0.01fF
C1080 INVX1_LOC_607/A INVX1_LOC_547/Y 0.04fF
C1081 INVX1_LOC_160/Y INVX1_LOC_271/A 0.01fF
C1082 INVX1_LOC_454/A INVX1_LOC_602/A 0.07fF
C1083 INVX1_LOC_182/A INVX1_LOC_85/Y 0.00fF
C1084 INVX1_LOC_190/A NAND2X1_LOC_85/a_36_24# 0.00fF
C1085 NAND2X1_LOC_54/a_36_24# INVX1_LOC_99/Y 0.00fF
C1086 INPUT_0 INVX1_LOC_126/Y 0.03fF
C1087 NAND2X1_LOC_24/Y INVX1_LOC_206/Y 0.39fF
C1088 VDD INVX1_LOC_275/Y 0.23fF
C1089 NAND2X1_LOC_543/B INVX1_LOC_17/Y 0.47fF
C1090 INVX1_LOC_288/Y INVX1_LOC_594/Y 0.00fF
C1091 INVX1_LOC_418/Y NAND2X1_LOC_373/Y 0.01fF
C1092 INVX1_LOC_566/A INVX1_LOC_586/A 0.00fF
C1093 INVX1_LOC_607/A INVX1_LOC_651/A 0.27fF
C1094 INVX1_LOC_395/A INVX1_LOC_670/Y 0.63fF
C1095 INVX1_LOC_446/A INVX1_LOC_93/Y 0.19fF
C1096 VDD NAND2X1_LOC_84/B 0.01fF
C1097 NAND2X1_LOC_10/a_36_24# INVX1_LOC_66/A 0.01fF
C1098 NAND2X1_LOC_690/Y INVX1_LOC_358/Y 0.01fF
C1099 VDD INVX1_LOC_444/A 0.00fF
C1100 VDD INVX1_LOC_343/Y 0.21fF
C1101 VDD INVX1_LOC_535/Y 0.21fF
C1102 INVX1_LOC_335/Y NAND2X1_LOC_690/Y 0.01fF
C1103 INVX1_LOC_405/A NAND2X1_LOC_520/A 0.09fF
C1104 INVX1_LOC_603/Y INVX1_LOC_94/A 0.03fF
C1105 INVX1_LOC_381/A INVX1_LOC_486/Y 0.07fF
C1106 INVX1_LOC_294/Y INVX1_LOC_381/A 0.00fF
C1107 INVX1_LOC_287/A INVX1_LOC_51/Y 0.01fF
C1108 NAND2X1_LOC_732/a_36_24# INVX1_LOC_523/A 0.00fF
C1109 INVX1_LOC_270/A INVX1_LOC_318/Y 0.00fF
C1110 INVX1_LOC_375/A NAND2X1_LOC_602/A 0.01fF
C1111 NAND2X1_LOC_545/B INVX1_LOC_551/Y 0.03fF
C1112 NAND2X1_LOC_122/Y INVX1_LOC_99/Y 0.03fF
C1113 INVX1_LOC_150/A INVX1_LOC_496/Y 0.01fF
C1114 INVX1_LOC_364/Y INVX1_LOC_363/Y 0.24fF
C1115 NAND2X1_LOC_322/Y NAND2X1_LOC_325/a_36_24# 0.00fF
C1116 INVX1_LOC_20/Y INVX1_LOC_377/A 0.01fF
C1117 VDD INVX1_LOC_638/Y 0.39fF
C1118 INVX1_LOC_522/Y INVX1_LOC_474/Y 0.05fF
C1119 INVX1_LOC_617/Y INVX1_LOC_371/Y 0.01fF
C1120 NAND2X1_LOC_786/B INVX1_LOC_615/A 0.00fF
C1121 NAND2X1_LOC_537/A NAND2X1_LOC_52/Y 0.10fF
C1122 INVX1_LOC_412/Y INVX1_LOC_89/Y 0.03fF
C1123 INVX1_LOC_651/Y INVX1_LOC_145/Y 0.20fF
C1124 INVX1_LOC_537/A INVX1_LOC_356/A 0.01fF
C1125 NAND2X1_LOC_704/B INVX1_LOC_251/Y 0.05fF
C1126 INVX1_LOC_435/A NAND2X1_LOC_620/a_36_24# 0.00fF
C1127 INVX1_LOC_271/A NAND2X1_LOC_267/A 0.63fF
C1128 VDD INVX1_LOC_357/Y 0.21fF
C1129 INVX1_LOC_463/A NAND2X1_LOC_686/A 0.09fF
C1130 NAND2X1_LOC_320/a_36_24# INVX1_LOC_47/Y 0.00fF
C1131 NAND2X1_LOC_387/Y INVX1_LOC_397/A 0.23fF
C1132 INVX1_LOC_551/Y INVX1_LOC_98/Y 0.10fF
C1133 INVX1_LOC_93/Y INVX1_LOC_374/A 0.03fF
C1134 INVX1_LOC_140/Y INVX1_LOC_470/Y 0.01fF
C1135 INPUT_0 INVX1_LOC_199/Y 0.76fF
C1136 INVX1_LOC_127/A INVX1_LOC_47/Y 0.03fF
C1137 NAND2X1_LOC_387/Y INVX1_LOC_94/A 0.01fF
C1138 INVX1_LOC_435/A INVX1_LOC_84/A 0.00fF
C1139 INVX1_LOC_271/Y INVX1_LOC_32/Y 0.01fF
C1140 INVX1_LOC_412/Y INVX1_LOC_501/A 0.03fF
C1141 INVX1_LOC_500/Y INVX1_LOC_501/Y 0.14fF
C1142 NAND2X1_LOC_637/A INVX1_LOC_79/A 0.03fF
C1143 INVX1_LOC_134/Y INVX1_LOC_363/Y 0.03fF
C1144 NAND2X1_LOC_789/A INVX1_LOC_366/A 0.03fF
C1145 INVX1_LOC_90/Y INVX1_LOC_596/Y 0.02fF
C1146 INVX1_LOC_444/Y INVX1_LOC_489/A 0.02fF
C1147 INVX1_LOC_447/A INVX1_LOC_26/Y 0.03fF
C1148 NAND2X1_LOC_780/A INVX1_LOC_54/Y 0.01fF
C1149 INVX1_LOC_213/Y INVX1_LOC_293/Y 0.02fF
C1150 INVX1_LOC_395/A INVX1_LOC_63/Y 0.35fF
C1151 INVX1_LOC_89/Y INVX1_LOC_321/A 0.03fF
C1152 NAND2X1_LOC_427/Y INVX1_LOC_498/A 0.13fF
C1153 INVX1_LOC_17/Y INVX1_LOC_469/A 0.01fF
C1154 INVX1_LOC_310/Y INVX1_LOC_35/Y 0.01fF
C1155 INVX1_LOC_517/A INVX1_LOC_50/Y 0.01fF
C1156 INVX1_LOC_466/A INVX1_LOC_495/A 0.02fF
C1157 INVX1_LOC_42/A NAND2X1_LOC_84/B 0.03fF
C1158 NAND2X1_LOC_766/a_36_24# INVX1_LOC_53/Y 0.00fF
C1159 INVX1_LOC_617/Y INVX1_LOC_89/Y 0.10fF
C1160 INVX1_LOC_89/Y INVX1_LOC_119/A 0.01fF
C1161 INVX1_LOC_406/Y NAND2X1_LOC_292/Y 0.01fF
C1162 VDD INVX1_LOC_274/Y 0.07fF
C1163 NAND2X1_LOC_57/a_36_24# INVX1_LOC_178/A 0.01fF
C1164 INVX1_LOC_307/Y INVX1_LOC_41/Y 0.01fF
C1165 INVX1_LOC_344/Y INVX1_LOC_513/A 0.00fF
C1166 INVX1_LOC_261/Y INVX1_LOC_111/A 0.00fF
C1167 NAND2X1_LOC_271/B INVX1_LOC_41/Y 0.00fF
C1168 INVX1_LOC_21/Y NAND2X1_LOC_706/B 0.15fF
C1169 INVX1_LOC_99/Y NAND2X1_LOC_406/a_36_24# 0.00fF
C1170 INVX1_LOC_137/Y NAND2X1_LOC_708/A 0.12fF
C1171 INVX1_LOC_412/Y NAND2X1_LOC_544/B 0.01fF
C1172 INVX1_LOC_6/Y INVX1_LOC_29/Y 0.04fF
C1173 NAND2X1_LOC_384/a_36_24# INVX1_LOC_9/Y 0.00fF
C1174 INVX1_LOC_49/Y INVX1_LOC_134/Y 0.10fF
C1175 INVX1_LOC_69/Y INVX1_LOC_632/A 0.51fF
C1176 INVX1_LOC_586/A INVX1_LOC_79/A 0.17fF
C1177 INVX1_LOC_202/Y NAND2X1_LOC_165/Y 0.02fF
C1178 INVX1_LOC_417/Y INVX1_LOC_69/Y 0.18fF
C1179 INVX1_LOC_655/Y INVX1_LOC_664/A 0.05fF
C1180 INVX1_LOC_287/Y INVX1_LOC_90/Y 0.02fF
C1181 INVX1_LOC_32/Y INVX1_LOC_480/Y 0.06fF
C1182 INVX1_LOC_164/Y INVX1_LOC_117/Y 0.15fF
C1183 INVX1_LOC_45/Y INVX1_LOC_653/Y 0.09fF
C1184 INVX1_LOC_117/Y NAND2X1_LOC_333/B 1.16fF
C1185 INVX1_LOC_607/Y INVX1_LOC_199/Y 0.21fF
C1186 INVX1_LOC_284/A INVX1_LOC_63/Y 0.00fF
C1187 INVX1_LOC_80/A INVX1_LOC_245/A 0.03fF
C1188 NAND2X1_LOC_20/Y INVX1_LOC_26/Y 0.15fF
C1189 INVX1_LOC_69/Y INVX1_LOC_59/Y 0.07fF
C1190 INVX1_LOC_51/Y INVX1_LOC_588/A 0.06fF
C1191 INVX1_LOC_318/A INVX1_LOC_254/A 0.02fF
C1192 INVX1_LOC_91/A INVX1_LOC_94/A 0.22fF
C1193 INVX1_LOC_587/A INVX1_LOC_74/Y 0.03fF
C1194 NAND2X1_LOC_48/a_36_24# INVX1_LOC_328/Y 0.00fF
C1195 INVX1_LOC_49/Y INVX1_LOC_235/A 0.08fF
C1196 INVX1_LOC_579/Y INVX1_LOC_245/A 0.08fF
C1197 NAND2X1_LOC_710/A NAND2X1_LOC_601/Y 0.01fF
C1198 INVX1_LOC_312/Y INVX1_LOC_79/A 0.04fF
C1199 INVX1_LOC_32/Y INVX1_LOC_169/Y 0.46fF
C1200 INVX1_LOC_300/A NAND2X1_LOC_641/a_36_24# 0.00fF
C1201 INVX1_LOC_548/A INVX1_LOC_63/Y 0.00fF
C1202 INVX1_LOC_69/Y INVX1_LOC_48/Y 1.31fF
C1203 INVX1_LOC_117/Y INVX1_LOC_261/Y 0.06fF
C1204 INVX1_LOC_326/A INVX1_LOC_46/Y 0.01fF
C1205 NAND2X1_LOC_645/a_36_24# INVX1_LOC_376/Y 0.00fF
C1206 INVX1_LOC_300/A NAND2X1_LOC_665/a_36_24# 0.00fF
C1207 NAND2X1_LOC_299/Y INVX1_LOC_62/Y 0.07fF
C1208 INVX1_LOC_493/A INVX1_LOC_338/Y 0.01fF
C1209 INVX1_LOC_41/Y INVX1_LOC_633/Y 0.08fF
C1210 INVX1_LOC_476/A INVX1_LOC_46/Y 0.00fF
C1211 INVX1_LOC_167/A INVX1_LOC_338/Y 0.02fF
C1212 NAND2X1_LOC_755/B INVX1_LOC_90/Y 0.04fF
C1213 NAND2X1_LOC_569/a_36_24# INVX1_LOC_244/Y 0.00fF
C1214 NAND2X1_LOC_833/B NAND2X1_LOC_259/A 0.02fF
C1215 INVX1_LOC_468/Y INVX1_LOC_114/A 1.20fF
C1216 INVX1_LOC_58/Y INVX1_LOC_374/Y 0.03fF
C1217 INVX1_LOC_11/Y INVX1_LOC_245/A 0.10fF
C1218 INVX1_LOC_31/Y INVX1_LOC_63/Y 0.31fF
C1219 INVX1_LOC_211/Y INVX1_LOC_90/Y 0.25fF
C1220 NAND2X1_LOC_104/a_36_24# INVX1_LOC_63/Y 0.00fF
C1221 NAND2X1_LOC_529/Y NAND2X1_LOC_631/B 0.04fF
C1222 INVX1_LOC_203/A INVX1_LOC_197/Y 0.01fF
C1223 INVX1_LOC_298/A INVX1_LOC_272/A 0.02fF
C1224 INVX1_LOC_74/Y INVX1_LOC_252/A 0.01fF
C1225 INVX1_LOC_46/Y INVX1_LOC_90/Y 0.07fF
C1226 NAND2X1_LOC_646/A INVX1_LOC_473/Y 0.02fF
C1227 NAND2X1_LOC_184/Y INVX1_LOC_62/Y 0.45fF
C1228 INVX1_LOC_100/Y INVX1_LOC_6/Y 0.92fF
C1229 INVX1_LOC_459/A VDD 0.00fF
C1230 INVX1_LOC_157/Y INVX1_LOC_79/A 0.01fF
C1231 INVX1_LOC_317/A INVX1_LOC_41/Y 0.00fF
C1232 NAND2X1_LOC_184/Y NAND2X1_LOC_844/A 0.05fF
C1233 INVX1_LOC_166/A NAND2X1_LOC_433/a_36_24# 0.00fF
C1234 INVX1_LOC_204/Y INVX1_LOC_621/A 0.04fF
C1235 INVX1_LOC_63/Y INVX1_LOC_473/Y 0.07fF
C1236 INVX1_LOC_384/A INVX1_LOC_109/Y 0.07fF
C1237 INVX1_LOC_79/A INVX1_LOC_225/Y 0.01fF
C1238 INVX1_LOC_58/Y NAND2X1_LOC_843/B 0.36fF
C1239 INVX1_LOC_183/A INVX1_LOC_11/A 0.11fF
C1240 INVX1_LOC_199/Y INVX1_LOC_211/A 0.17fF
C1241 VDD INVX1_LOC_308/Y 0.26fF
C1242 INVX1_LOC_75/Y INVX1_LOC_9/Y 0.22fF
C1243 INVX1_LOC_58/Y INVX1_LOC_625/Y 0.03fF
C1244 INVX1_LOC_58/Y INVX1_LOC_91/Y 0.01fF
C1245 INVX1_LOC_124/A INVX1_LOC_479/A 0.01fF
C1246 NAND2X1_LOC_374/a_36_24# INVX1_LOC_442/A 0.00fF
C1247 NAND2X1_LOC_475/A NAND2X1_LOC_370/A 0.07fF
C1248 INVX1_LOC_448/A INVX1_LOC_109/Y 0.07fF
C1249 INVX1_LOC_578/A NAND2X1_LOC_457/A 0.01fF
C1250 NAND2X1_LOC_573/a_36_24# INVX1_LOC_51/Y 0.00fF
C1251 INVX1_LOC_145/Y INVX1_LOC_109/Y 0.07fF
C1252 GATE_579 INVX1_LOC_434/A 0.33fF
C1253 NAND2X1_LOC_597/Y INVX1_LOC_505/Y 0.04fF
C1254 INVX1_LOC_62/Y INVX1_LOC_75/Y 0.11fF
C1255 INVX1_LOC_570/A INVX1_LOC_523/A 0.39fF
C1256 NAND2X1_LOC_764/a_36_24# INVX1_LOC_366/A 0.00fF
C1257 INVX1_LOC_224/Y INVX1_LOC_482/A 0.02fF
C1258 INVX1_LOC_75/Y NAND2X1_LOC_844/A 0.09fF
C1259 NAND2X1_LOC_526/Y INVX1_LOC_413/Y 0.06fF
C1260 VDD NAND2X1_LOC_548/B 0.03fF
C1261 NAND2X1_LOC_274/B INVX1_LOC_92/A 0.03fF
C1262 INVX1_LOC_600/A INVX1_LOC_388/Y 0.33fF
C1263 NAND2X1_LOC_637/A INVX1_LOC_632/A 0.06fF
C1264 VDD INVX1_LOC_635/A 0.21fF
C1265 INVX1_LOC_301/A INVX1_LOC_67/Y 0.09fF
C1266 INVX1_LOC_207/A INVX1_LOC_366/A 0.32fF
C1267 VDD NAND2X1_LOC_237/Y 0.30fF
C1268 NAND2X1_LOC_45/Y INVX1_LOC_519/A 0.03fF
C1269 INVX1_LOC_20/Y INVX1_LOC_584/Y 0.04fF
C1270 INVX1_LOC_17/Y INVX1_LOC_409/Y 0.02fF
C1271 INVX1_LOC_62/Y NAND2X1_LOC_271/A 0.00fF
C1272 VDD INVX1_LOC_451/Y 0.03fF
C1273 INPUT_0 INVX1_LOC_53/Y 2.50fF
C1274 INVX1_LOC_21/Y INVX1_LOC_307/Y 0.01fF
C1275 INVX1_LOC_335/Y INVX1_LOC_562/A 0.05fF
C1276 NAND2X1_LOC_374/a_36_24# INVX1_LOC_116/Y 0.00fF
C1277 INVX1_LOC_68/Y INVX1_LOC_286/Y 0.09fF
C1278 INVX1_LOC_410/Y INVX1_LOC_371/Y 0.01fF
C1279 INVX1_LOC_442/A INVX1_LOC_634/A 0.03fF
C1280 INVX1_LOC_21/Y INVX1_LOC_97/A 0.10fF
C1281 NAND2X1_LOC_764/a_36_24# INVX1_LOC_597/A 0.00fF
C1282 INVX1_LOC_207/A NAND2X1_LOC_240/a_36_24# 0.00fF
C1283 NAND2X1_LOC_498/Y INVX1_LOC_519/A 0.03fF
C1284 NAND2X1_LOC_516/Y INVX1_LOC_53/Y 1.69fF
C1285 INVX1_LOC_32/Y INVX1_LOC_638/A 0.07fF
C1286 INVX1_LOC_586/A INVX1_LOC_511/A 0.00fF
C1287 INVX1_LOC_418/A NAND2X1_LOC_545/B 0.01fF
C1288 INVX1_LOC_224/Y INVX1_LOC_194/A 0.02fF
C1289 NAND2X1_LOC_498/B INVX1_LOC_134/Y 0.10fF
C1290 INVX1_LOC_276/A INVX1_LOC_101/Y 0.01fF
C1291 NAND2X1_LOC_537/A INVX1_LOC_318/A 0.09fF
C1292 INVX1_LOC_45/Y INVX1_LOC_97/Y 0.00fF
C1293 INVX1_LOC_228/Y INVX1_LOC_230/A 0.03fF
C1294 INVX1_LOC_206/Y INVX1_LOC_259/Y 0.03fF
C1295 INVX1_LOC_289/Y INVX1_LOC_290/A 0.15fF
C1296 INVX1_LOC_586/A INVX1_LOC_632/A 0.07fF
C1297 INVX1_LOC_51/Y INVX1_LOC_670/Y 0.86fF
C1298 INVX1_LOC_20/Y INVX1_LOC_63/A 0.03fF
C1299 INVX1_LOC_76/Y INVX1_LOC_134/Y 0.23fF
C1300 INVX1_LOC_417/Y INVX1_LOC_586/A 0.05fF
C1301 INVX1_LOC_584/A INVX1_LOC_513/A 0.10fF
C1302 INVX1_LOC_560/A INVX1_LOC_411/A 0.04fF
C1303 NAND2X1_LOC_527/Y NAND2X1_LOC_457/A 0.03fF
C1304 INVX1_LOC_340/Y INVX1_LOC_526/Y 0.03fF
C1305 INVX1_LOC_377/Y INVX1_LOC_519/A 0.04fF
C1306 INVX1_LOC_651/Y NAND2X1_LOC_260/Y 0.00fF
C1307 INVX1_LOC_586/A INVX1_LOC_491/Y 0.01fF
C1308 NAND2X1_LOC_780/A NAND2X1_LOC_677/Y 0.02fF
C1309 INVX1_LOC_391/Y INVX1_LOC_45/Y 0.01fF
C1310 INVX1_LOC_68/Y INVX1_LOC_17/Y 0.04fF
C1311 NAND2X1_LOC_181/a_36_24# INVX1_LOC_45/Y 0.00fF
C1312 INVX1_LOC_51/Y INVX1_LOC_506/Y 0.03fF
C1313 INVX1_LOC_586/A INVX1_LOC_59/Y 0.06fF
C1314 INVX1_LOC_278/A NAND2X1_LOC_850/a_36_24# 0.00fF
C1315 INVX1_LOC_431/A INVX1_LOC_45/Y 0.00fF
C1316 INVX1_LOC_46/Y NAND2X1_LOC_42/a_36_24# 0.01fF
C1317 INVX1_LOC_124/Y INVX1_LOC_126/A 0.00fF
C1318 INVX1_LOC_410/Y INVX1_LOC_89/Y 0.07fF
C1319 NAND2X1_LOC_79/Y INVX1_LOC_145/Y 0.01fF
C1320 INVX1_LOC_206/Y INVX1_LOC_204/Y 0.02fF
C1321 INVX1_LOC_51/Y INVX1_LOC_623/Y 0.38fF
C1322 INVX1_LOC_586/A INVX1_LOC_48/Y 0.22fF
C1323 INVX1_LOC_90/A INVX1_LOC_12/Y 0.03fF
C1324 INVX1_LOC_245/A NAND2X1_LOC_590/a_36_24# 0.01fF
C1325 INVX1_LOC_302/A INVX1_LOC_166/A 0.01fF
C1326 INVX1_LOC_412/A NAND2X1_LOC_388/A 0.01fF
C1327 INVX1_LOC_270/A INVX1_LOC_98/Y 0.30fF
C1328 INVX1_LOC_438/A INVX1_LOC_379/Y 0.01fF
C1329 INVX1_LOC_375/A INVX1_LOC_89/Y 0.12fF
C1330 INVX1_LOC_523/A INVX1_LOC_568/A -0.02fF
C1331 INVX1_LOC_374/A INVX1_LOC_31/Y 0.04fF
C1332 INVX1_LOC_293/Y INVX1_LOC_679/A 0.00fF
C1333 INVX1_LOC_89/Y INVX1_LOC_546/A 0.01fF
C1334 INVX1_LOC_634/A INVX1_LOC_116/Y 0.01fF
C1335 INVX1_LOC_285/A INVX1_LOC_145/Y 0.01fF
C1336 INVX1_LOC_85/Y INVX1_LOC_543/Y 0.01fF
C1337 INVX1_LOC_45/Y INVX1_LOC_18/Y 0.01fF
C1338 INVX1_LOC_607/Y INVX1_LOC_53/Y 0.15fF
C1339 NAND2X1_LOC_332/B INVX1_LOC_105/Y 0.03fF
C1340 INVX1_LOC_207/A INVX1_LOC_6/Y 0.01fF
C1341 NAND2X1_LOC_165/Y INVX1_LOC_76/Y 0.04fF
C1342 INVX1_LOC_202/Y INVX1_LOC_318/Y 0.11fF
C1343 INVX1_LOC_442/Y INVX1_LOC_104/Y 0.01fF
C1344 NAND2X1_LOC_168/a_36_24# INVX1_LOC_586/A 0.00fF
C1345 NAND2X1_LOC_148/B NAND2X1_LOC_149/a_36_24# 0.01fF
C1346 INVX1_LOC_94/Y NAND2X1_LOC_506/B 0.19fF
C1347 INVX1_LOC_686/A INVX1_LOC_259/Y 0.00fF
C1348 INVX1_LOC_323/Y INVX1_LOC_99/Y 0.01fF
C1349 INVX1_LOC_31/A INVX1_LOC_18/Y 0.03fF
C1350 INVX1_LOC_17/Y INVX1_LOC_600/A 1.23fF
C1351 INVX1_LOC_45/Y INVX1_LOC_94/Y 0.07fF
C1352 INVX1_LOC_398/A INVX1_LOC_32/Y 0.01fF
C1353 INVX1_LOC_312/Y INVX1_LOC_48/Y 0.04fF
C1354 INVX1_LOC_206/Y INVX1_LOC_114/A 0.12fF
C1355 INVX1_LOC_684/Y INVX1_LOC_685/A 0.15fF
C1356 INVX1_LOC_602/Y NAND2X1_LOC_864/a_36_24# 0.00fF
C1357 INVX1_LOC_619/A GATE_222 0.03fF
C1358 INVX1_LOC_84/A INVX1_LOC_93/Y 0.17fF
C1359 INVX1_LOC_319/Y INVX1_LOC_245/A 0.01fF
C1360 INVX1_LOC_444/Y NAND2X1_LOC_415/B 0.03fF
C1361 INVX1_LOC_437/A INVX1_LOC_385/Y 0.06fF
C1362 NAND2X1_LOC_523/B INVX1_LOC_46/Y 0.06fF
C1363 INVX1_LOC_51/Y INVX1_LOC_63/Y 0.10fF
C1364 INVX1_LOC_451/A INVX1_LOC_7/Y 2.43fF
C1365 INVX1_LOC_330/A NAND2X1_LOC_679/B 0.04fF
C1366 INVX1_LOC_463/A INVX1_LOC_588/A 0.08fF
C1367 INVX1_LOC_266/A INVX1_LOC_253/Y 0.01fF
C1368 INVX1_LOC_298/A INVX1_LOC_53/Y 0.03fF
C1369 NAND2X1_LOC_591/a_36_24# INVX1_LOC_32/Y 0.01fF
C1370 INVX1_LOC_639/Y GATE_865 0.01fF
C1371 NAND2X1_LOC_638/A INVX1_LOC_497/Y 0.03fF
C1372 NAND2X1_LOC_48/a_36_24# INVX1_LOC_172/A 0.00fF
C1373 NAND2X1_LOC_545/B INVX1_LOC_46/Y 0.01fF
C1374 INVX1_LOC_452/A INVX1_LOC_453/Y 0.11fF
C1375 INVX1_LOC_140/Y INVX1_LOC_79/A 0.28fF
C1376 NAND2X1_LOC_336/B NAND2X1_LOC_388/A 0.00fF
C1377 INVX1_LOC_259/A INVX1_LOC_26/Y 0.00fF
C1378 INVX1_LOC_35/Y INVX1_LOC_304/Y 0.03fF
C1379 INVX1_LOC_513/A INVX1_LOC_537/A 0.01fF
C1380 INVX1_LOC_20/Y INVX1_LOC_347/Y 0.13fF
C1381 INVX1_LOC_412/Y INVX1_LOC_347/A 0.20fF
C1382 INVX1_LOC_595/Y INVX1_LOC_35/Y 0.02fF
C1383 INVX1_LOC_288/Y NAND2X1_LOC_635/B 0.02fF
C1384 INVX1_LOC_555/A INVX1_LOC_633/Y 0.02fF
C1385 INVX1_LOC_395/A INVX1_LOC_669/A 0.03fF
C1386 NAND2X1_LOC_318/A INVX1_LOC_351/A 0.03fF
C1387 INVX1_LOC_266/A INVX1_LOC_63/Y 0.00fF
C1388 INVX1_LOC_442/Y INVX1_LOC_117/Y 0.07fF
C1389 INVX1_LOC_47/Y INVX1_LOC_519/A 0.05fF
C1390 INVX1_LOC_45/Y NAND2X1_LOC_489/A 0.01fF
C1391 NAND2X1_LOC_692/Y INVX1_LOC_117/Y 0.01fF
C1392 NAND2X1_LOC_27/Y INVX1_LOC_11/Y 0.03fF
C1393 INVX1_LOC_93/Y NAND2X1_LOC_67/Y 0.01fF
C1394 INVX1_LOC_20/Y INVX1_LOC_328/Y 0.35fF
C1395 INVX1_LOC_93/Y INVX1_LOC_129/A 0.02fF
C1396 INVX1_LOC_277/A INVX1_LOC_662/Y 0.02fF
C1397 INVX1_LOC_84/A INVX1_LOC_390/A 0.00fF
C1398 INVX1_LOC_20/Y INVX1_LOC_518/A 0.03fF
C1399 INVX1_LOC_366/A INVX1_LOC_79/A 0.00fF
C1400 INVX1_LOC_321/Y INVX1_LOC_431/Y 0.12fF
C1401 INVX1_LOC_410/A INVX1_LOC_12/Y 0.00fF
C1402 INVX1_LOC_566/Y INVX1_LOC_245/A 0.05fF
C1403 NAND2X1_LOC_318/A INVX1_LOC_90/Y 0.07fF
C1404 INVX1_LOC_451/A INVX1_LOC_32/Y 0.10fF
C1405 INVX1_LOC_522/A INVX1_LOC_335/A 0.27fF
C1406 INVX1_LOC_46/Y INVX1_LOC_98/Y 0.00fF
C1407 INVX1_LOC_607/A INVX1_LOC_62/Y 0.04fF
C1408 INVX1_LOC_317/Y INVX1_LOC_41/Y 0.05fF
C1409 INVX1_LOC_17/Y INVX1_LOC_484/A -0.07fF
C1410 NAND2X1_LOC_190/A NAND2X1_LOC_184/Y 0.23fF
C1411 INVX1_LOC_370/Y INVX1_LOC_49/Y 0.04fF
C1412 INVX1_LOC_68/Y NAND2X1_LOC_231/a_36_24# 0.00fF
C1413 INVX1_LOC_32/Y INVX1_LOC_665/Y 0.33fF
C1414 INVX1_LOC_145/Y INVX1_LOC_199/Y 1.03fF
C1415 INVX1_LOC_488/Y INVX1_LOC_49/A 0.04fF
C1416 INVX1_LOC_686/A INVX1_LOC_114/A 0.04fF
C1417 INVX1_LOC_99/Y INVX1_LOC_659/A 0.13fF
C1418 INVX1_LOC_272/Y INVX1_LOC_79/A 0.06fF
C1419 NAND2X1_LOC_791/B INVX1_LOC_79/A 0.02fF
C1420 INVX1_LOC_79/A INVX1_LOC_486/Y 0.02fF
C1421 INVX1_LOC_170/A INVX1_LOC_176/A 0.01fF
C1422 INVX1_LOC_317/A NAND2X1_LOC_267/A 0.01fF
C1423 INVX1_LOC_119/Y INVX1_LOC_519/A 0.27fF
C1424 INPUT_0 NAND2X1_LOC_60/Y 0.01fF
C1425 INVX1_LOC_157/Y INVX1_LOC_48/Y 0.16fF
C1426 NAND2X1_LOC_448/B NAND2X1_LOC_422/a_36_24# 0.02fF
C1427 NAND2X1_LOC_333/A NAND2X1_LOC_171/a_36_24# 0.02fF
C1428 INVX1_LOC_183/A INVX1_LOC_35/Y 0.03fF
C1429 NAND2X1_LOC_334/A INVX1_LOC_259/Y 0.03fF
C1430 INVX1_LOC_376/Y INVX1_LOC_504/Y 0.04fF
C1431 INVX1_LOC_432/Y INVX1_LOC_245/A 0.01fF
C1432 INVX1_LOC_202/Y INVX1_LOC_351/A 0.00fF
C1433 INVX1_LOC_513/Y INVX1_LOC_514/A 0.01fF
C1434 INVX1_LOC_164/Y INVX1_LOC_58/Y 0.01fF
C1435 INVX1_LOC_323/Y NAND2X1_LOC_66/Y 0.02fF
C1436 NAND2X1_LOC_561/a_36_24# INVX1_LOC_9/Y 0.01fF
C1437 INVX1_LOC_492/A INVX1_LOC_9/Y 0.02fF
C1438 INVX1_LOC_58/Y NAND2X1_LOC_333/B 0.17fF
C1439 INVX1_LOC_54/Y INVX1_LOC_309/Y 0.01fF
C1440 INVX1_LOC_93/Y INVX1_LOC_496/A 0.19fF
C1441 INVX1_LOC_79/A INVX1_LOC_252/A 0.03fF
C1442 NAND2X1_LOC_181/A INVX1_LOC_6/Y 0.01fF
C1443 NAND2X1_LOC_521/Y INVX1_LOC_420/A 0.03fF
C1444 INVX1_LOC_202/Y INVX1_LOC_90/Y 1.42fF
C1445 INVX1_LOC_207/Y INVX1_LOC_197/Y 0.69fF
C1446 INVX1_LOC_261/Y INVX1_LOC_58/Y 0.03fF
C1447 INVX1_LOC_166/A INVX1_LOC_301/Y 0.00fF
C1448 INVX1_LOC_53/Y INVX1_LOC_464/Y 0.12fF
C1449 NAND2X1_LOC_706/B INVX1_LOC_26/Y 0.06fF
C1450 NAND2X1_LOC_274/B INPUT_1 0.07fF
C1451 INVX1_LOC_492/A INVX1_LOC_62/Y 0.12fF
C1452 INVX1_LOC_75/A INVX1_LOC_98/Y 0.01fF
C1453 INVX1_LOC_100/Y NAND2X1_LOC_294/Y 0.05fF
C1454 INVX1_LOC_166/A INVX1_LOC_41/Y 1.37fF
C1455 INVX1_LOC_6/Y INVX1_LOC_79/A 0.55fF
C1456 INVX1_LOC_54/Y INVX1_LOC_479/A 4.48fF
C1457 INVX1_LOC_288/Y INVX1_LOC_462/Y 0.05fF
C1458 INVX1_LOC_6/Y NAND2X1_LOC_631/B 0.03fF
C1459 INVX1_LOC_49/Y INVX1_LOC_90/Y 0.09fF
C1460 NAND2X1_LOC_334/A INVX1_LOC_114/A 0.03fF
C1461 VDD INVX1_LOC_465/Y 0.27fF
C1462 INVX1_LOC_641/A INVX1_LOC_454/Y 0.09fF
C1463 NAND2X1_LOC_111/Y INVX1_LOC_41/Y 0.14fF
C1464 INVX1_LOC_100/Y INVX1_LOC_206/A 0.05fF
C1465 INVX1_LOC_257/A INVX1_LOC_479/A 0.07fF
C1466 NAND2X1_LOC_332/B INVX1_LOC_109/Y 0.00fF
C1467 INVX1_LOC_328/Y NAND2X1_LOC_269/B 0.02fF
C1468 VDD INVX1_LOC_572/A -0.00fF
C1469 INVX1_LOC_418/Y INVX1_LOC_92/A 0.02fF
C1470 INVX1_LOC_319/A INVX1_LOC_245/A 0.01fF
C1471 INVX1_LOC_159/Y INVX1_LOC_92/A 0.07fF
C1472 NAND2X1_LOC_637/A INVX1_LOC_561/Y 0.00fF
C1473 VDD INVX1_LOC_292/A -0.00fF
C1474 INVX1_LOC_446/A INVX1_LOC_51/Y 0.05fF
C1475 VDD INVX1_LOC_107/A 0.00fF
C1476 NAND2X1_LOC_750/Y NAND2X1_LOC_749/Y 0.04fF
C1477 INVX1_LOC_3/Y INVX1_LOC_1/A 0.01fF
C1478 INVX1_LOC_202/A INVX1_LOC_586/A 0.08fF
C1479 INVX1_LOC_376/A INVX1_LOC_348/Y 0.03fF
C1480 INVX1_LOC_92/Y INVX1_LOC_90/Y 0.02fF
C1481 INVX1_LOC_531/Y INVX1_LOC_41/Y 0.07fF
C1482 NAND2X1_LOC_342/A INVX1_LOC_240/Y 0.06fF
C1483 INVX1_LOC_445/Y INVX1_LOC_445/A 0.00fF
C1484 INVX1_LOC_301/Y INVX1_LOC_363/A 0.01fF
C1485 VDD INVX1_LOC_515/A -0.00fF
C1486 INVX1_LOC_191/Y INVX1_LOC_366/A -0.05fF
C1487 NAND2X1_LOC_582/a_36_24# INVX1_LOC_632/A 0.01fF
C1488 INPUT_0 NAND2X1_LOC_383/Y 0.11fF
C1489 VDD INVX1_LOC_492/Y 0.49fF
C1490 INVX1_LOC_374/A INVX1_LOC_51/Y 0.03fF
C1491 INVX1_LOC_20/Y NAND2X1_LOC_536/a_36_24# 0.00fF
C1492 VDD NAND2X1_LOC_325/B 0.03fF
C1493 INVX1_LOC_84/A INVX1_LOC_395/A 0.19fF
C1494 INVX1_LOC_180/A INVX1_LOC_366/A 0.06fF
C1495 INVX1_LOC_490/Y INVX1_LOC_293/Y 0.02fF
C1496 INVX1_LOC_1/A NAND2X1_LOC_2/a_36_24# 0.00fF
C1497 INVX1_LOC_74/Y INVX1_LOC_636/A 0.07fF
C1498 INVX1_LOC_444/Y INVX1_LOC_453/A 0.03fF
C1499 INVX1_LOC_438/Y INVX1_LOC_385/Y 1.24fF
C1500 INVX1_LOC_20/Y INVX1_LOC_266/Y 0.00fF
C1501 INVX1_LOC_193/Y INVX1_LOC_12/Y 0.01fF
C1502 VDD NAND2X1_LOC_673/A -0.00fF
C1503 INVX1_LOC_446/Y INVX1_LOC_53/Y 0.13fF
C1504 INVX1_LOC_523/A INVX1_LOC_136/Y 0.00fF
C1505 NAND2X1_LOC_486/B INVX1_LOC_547/A 0.01fF
C1506 INVX1_LOC_578/A NAND2X1_LOC_302/a_36_24# 0.00fF
C1507 INVX1_LOC_255/Y INVX1_LOC_633/Y 0.02fF
C1508 INVX1_LOC_64/Y NAND2X1_LOC_60/Y 0.20fF
C1509 INVX1_LOC_228/Y NAND2X1_LOC_72/Y 0.07fF
C1510 INVX1_LOC_288/A INVX1_LOC_53/Y 0.07fF
C1511 INVX1_LOC_395/A INVX1_LOC_129/A 0.01fF
C1512 INVX1_LOC_395/A NAND2X1_LOC_67/Y 0.02fF
C1513 INVX1_LOC_76/Y INVX1_LOC_318/Y 0.14fF
C1514 VDD NAND2X1_LOC_482/Y 0.07fF
C1515 INVX1_LOC_618/A INVX1_LOC_63/Y 0.01fF
C1516 INVX1_LOC_502/Y INVX1_LOC_519/A 0.02fF
C1517 INVX1_LOC_242/Y INVX1_LOC_109/Y 0.99fF
C1518 INVX1_LOC_53/Y INVX1_LOC_384/A 0.07fF
C1519 NAND2X1_LOC_380/a_36_24# INVX1_LOC_366/A 0.00fF
C1520 NAND2X1_LOC_331/A NAND2X1_LOC_594/Y 0.02fF
C1521 VDD NAND2X1_LOC_285/A -0.00fF
C1522 INVX1_LOC_278/A INVX1_LOC_282/A 0.00fF
C1523 INVX1_LOC_560/A NAND2X1_LOC_775/B 0.02fF
C1524 INVX1_LOC_76/Y INVX1_LOC_16/Y 0.09fF
C1525 INVX1_LOC_3/Y INVX1_LOC_6/Y 0.30fF
C1526 INVX1_LOC_300/A INVX1_LOC_266/Y 0.13fF
C1527 INVX1_LOC_140/Y INVX1_LOC_48/Y 0.18fF
C1528 NAND2X1_LOC_756/Y INVX1_LOC_97/Y 0.01fF
C1529 INVX1_LOC_416/A NAND2X1_LOC_552/a_36_24# 0.00fF
C1530 INVX1_LOC_552/Y INVX1_LOC_254/A 0.04fF
C1531 VDD INVX1_LOC_351/Y 0.21fF
C1532 INVX1_LOC_414/A INVX1_LOC_6/Y 0.01fF
C1533 INVX1_LOC_400/Y INVX1_LOC_670/A 0.03fF
C1534 INVX1_LOC_288/A INVX1_LOC_460/Y 0.01fF
C1535 NAND2X1_LOC_318/A INVX1_LOC_98/Y 0.17fF
C1536 VDD INVX1_LOC_168/Y 1.75fF
C1537 INVX1_LOC_396/A INVX1_LOC_586/A 0.04fF
C1538 INVX1_LOC_317/Y NAND2X1_LOC_267/A 0.04fF
C1539 INVX1_LOC_474/Y INVX1_LOC_633/Y 0.09fF
C1540 INVX1_LOC_45/A INVX1_LOC_25/Y 0.01fF
C1541 INVX1_LOC_366/A INVX1_LOC_48/Y 0.18fF
C1542 INVX1_LOC_450/A NAND2X1_LOC_294/Y 0.00fF
C1543 INVX1_LOC_53/Y NAND2X1_LOC_612/A 0.03fF
C1544 INVX1_LOC_596/A NAND2X1_LOC_643/a_36_24# 0.01fF
C1545 NAND2X1_LOC_759/B INVX1_LOC_26/Y -0.04fF
C1546 NAND2X1_LOC_273/a_36_24# INVX1_LOC_509/A 0.00fF
C1547 NAND2X1_LOC_791/A INVX1_LOC_53/Y 0.01fF
C1548 INVX1_LOC_53/Y INVX1_LOC_145/Y 0.14fF
C1549 INVX1_LOC_211/Y INVX1_LOC_596/A 0.00fF
C1550 INVX1_LOC_117/Y NAND2X1_LOC_493/B 0.17fF
C1551 INVX1_LOC_224/Y INVX1_LOC_9/Y 0.07fF
C1552 INVX1_LOC_607/Y NAND2X1_LOC_148/A 0.04fF
C1553 INVX1_LOC_607/Y NAND2X1_LOC_107/Y 0.06fF
C1554 INVX1_LOC_175/Y INVX1_LOC_172/A 0.07fF
C1555 INPUT_3 NAND2X1_LOC_84/B 0.39fF
C1556 INVX1_LOC_20/Y INVX1_LOC_105/Y 0.04fF
C1557 INVX1_LOC_307/A INVX1_LOC_178/A 0.47fF
C1558 INVX1_LOC_180/A INVX1_LOC_6/Y 0.01fF
C1559 INVX1_LOC_84/A NAND2X1_LOC_83/a_36_24# 0.00fF
C1560 NAND2X1_LOC_791/B INVX1_LOC_48/Y 0.78fF
C1561 NAND2X1_LOC_97/B INVX1_LOC_252/Y 0.05fF
C1562 INVX1_LOC_162/Y INVX1_LOC_496/A 0.04fF
C1563 INPUT_0 INVX1_LOC_662/A 0.01fF
C1564 INVX1_LOC_355/A INVX1_LOC_63/Y 0.00fF
C1565 INVX1_LOC_272/Y INVX1_LOC_48/Y 0.05fF
C1566 INVX1_LOC_274/A INVX1_LOC_600/Y 0.01fF
C1567 INVX1_LOC_562/A INVX1_LOC_26/Y 0.09fF
C1568 NAND2X1_LOC_822/Y INVX1_LOC_59/A 0.01fF
C1569 INVX1_LOC_323/Y NAND2X1_LOC_43/Y 0.00fF
C1570 INVX1_LOC_578/A INVX1_LOC_9/Y 0.07fF
C1571 INVX1_LOC_117/Y INVX1_LOC_517/A 0.03fF
C1572 INVX1_LOC_97/A INVX1_LOC_26/Y 0.05fF
C1573 INVX1_LOC_6/Y INVX1_LOC_610/Y 0.01fF
C1574 INVX1_LOC_209/A INVX1_LOC_600/Y 0.00fF
C1575 INVX1_LOC_84/A INVX1_LOC_31/Y 0.33fF
C1576 INVX1_LOC_45/Y INVX1_LOC_357/Y 0.01fF
C1577 INVX1_LOC_384/A NAND2X1_LOC_274/Y 0.02fF
C1578 INVX1_LOC_345/Y INVX1_LOC_134/Y 0.03fF
C1579 INVX1_LOC_325/Y INVX1_LOC_326/Y 0.14fF
C1580 INVX1_LOC_54/Y INVX1_LOC_12/Y 0.09fF
C1581 INVX1_LOC_32/Y INVX1_LOC_134/Y 0.07fF
C1582 NAND2X1_LOC_523/B INVX1_LOC_387/Y 0.00fF
C1583 INVX1_LOC_597/A INVX1_LOC_48/Y 0.27fF
C1584 INVX1_LOC_521/Y INVX1_LOC_655/A 0.01fF
C1585 NAND2X1_LOC_65/Y INVX1_LOC_44/Y 0.06fF
C1586 NAND2X1_LOC_39/Y INVX1_LOC_47/Y 0.12fF
C1587 NAND2X1_LOC_756/Y INVX1_LOC_94/Y 0.04fF
C1588 INVX1_LOC_202/Y INVX1_LOC_98/Y 0.11fF
C1589 INVX1_LOC_249/Y INVX1_LOC_353/A 0.01fF
C1590 NAND2X1_LOC_710/A INVX1_LOC_69/Y 0.02fF
C1591 NAND2X1_LOC_13/Y INVX1_LOC_63/Y 0.04fF
C1592 INVX1_LOC_224/Y INVX1_LOC_62/Y 1.71fF
C1593 NAND2X1_LOC_325/B INVX1_LOC_103/Y 0.02fF
C1594 INVX1_LOC_140/Y INVX1_LOC_472/Y 0.01fF
C1595 INVX1_LOC_47/A INVX1_LOC_32/Y 0.01fF
C1596 INVX1_LOC_160/Y INVX1_LOC_153/Y 0.06fF
C1597 INVX1_LOC_69/Y NAND2X1_LOC_541/B 0.19fF
C1598 INVX1_LOC_21/Y INVX1_LOC_166/A 0.03fF
C1599 INVX1_LOC_282/A INVX1_LOC_453/Y 0.03fF
C1600 INVX1_LOC_549/Y INVX1_LOC_50/Y 0.19fF
C1601 INVX1_LOC_98/A INVX1_LOC_90/Y 0.01fF
C1602 INVX1_LOC_366/Y INVX1_LOC_46/Y 0.05fF
C1603 INVX1_LOC_681/Y INVX1_LOC_159/Y 0.02fF
C1604 INVX1_LOC_166/A NAND2X1_LOC_655/a_36_24# 0.00fF
C1605 INVX1_LOC_578/A INVX1_LOC_62/Y 0.15fF
C1606 NAND2X1_LOC_775/B INVX1_LOC_603/A 0.02fF
C1607 INVX1_LOC_651/Y INVX1_LOC_655/A 0.01fF
C1608 INVX1_LOC_680/Y INVX1_LOC_66/A 0.01fF
C1609 INVX1_LOC_258/A INVX1_LOC_376/A 0.04fF
C1610 INVX1_LOC_302/A INVX1_LOC_41/Y 0.01fF
C1611 INVX1_LOC_31/Y NAND2X1_LOC_67/Y 0.03fF
C1612 INVX1_LOC_636/A NAND2X1_LOC_591/B 0.02fF
C1613 INVX1_LOC_602/Y INVX1_LOC_340/A 0.11fF
C1614 NAND2X1_LOC_169/A NAND2X1_LOC_388/A 0.01fF
C1615 INVX1_LOC_307/A INVX1_LOC_58/Y 0.01fF
C1616 INVX1_LOC_76/Y INVX1_LOC_90/Y 1.60fF
C1617 INVX1_LOC_159/Y INPUT_1 0.10fF
C1618 NAND2X1_LOC_532/Y INVX1_LOC_516/A 0.14fF
C1619 INVX1_LOC_315/Y INVX1_LOC_531/Y 0.07fF
C1620 NAND2X1_LOC_601/a_36_24# INVX1_LOC_376/Y 0.00fF
C1621 INVX1_LOC_384/A NAND2X1_LOC_844/a_36_24# 0.01fF
C1622 INVX1_LOC_193/A INVX1_LOC_93/Y 0.09fF
C1623 INVX1_LOC_150/Y INVX1_LOC_479/A 0.01fF
C1624 INVX1_LOC_145/Y NAND2X1_LOC_274/Y 0.01fF
C1625 INVX1_LOC_58/Y INVX1_LOC_290/A 0.13fF
C1626 NAND2X1_LOC_195/a_36_24# INVX1_LOC_6/Y 0.00fF
C1627 INVX1_LOC_558/A NAND2X1_LOC_411/a_36_24# 0.01fF
C1628 INVX1_LOC_54/Y NAND2X1_LOC_521/Y 0.03fF
C1629 NAND2X1_LOC_165/Y INVX1_LOC_32/Y 0.02fF
C1630 NAND2X1_LOC_166/a_36_24# INVX1_LOC_63/Y 0.01fF
C1631 INVX1_LOC_49/Y INVX1_LOC_98/Y 0.10fF
C1632 NAND2X1_LOC_467/A INVX1_LOC_41/Y 0.18fF
C1633 INVX1_LOC_496/A INVX1_LOC_189/Y 0.01fF
C1634 INVX1_LOC_6/Y INVX1_LOC_48/Y 1.59fF
C1635 INVX1_LOC_315/Y INVX1_LOC_528/Y 0.01fF
C1636 INVX1_LOC_404/Y NAND2X1_LOC_271/A 0.00fF
C1637 NAND2X1_LOC_836/B INVX1_LOC_40/Y 0.12fF
C1638 INVX1_LOC_568/Y INVX1_LOC_9/Y 0.01fF
C1639 INVX1_LOC_47/Y INVX1_LOC_513/A 0.28fF
C1640 NAND2X1_LOC_329/a_36_24# GATE_865 0.00fF
C1641 NAND2X1_LOC_383/Y INVX1_LOC_211/A 0.01fF
C1642 INVX1_LOC_410/A NAND2X1_LOC_615/B 0.00fF
C1643 INVX1_LOC_248/Y INVX1_LOC_353/A 0.02fF
C1644 INVX1_LOC_207/Y INVX1_LOC_600/Y 0.16fF
C1645 INVX1_LOC_32/Y INVX1_LOC_65/A 0.03fF
C1646 INVX1_LOC_21/Y INVX1_LOC_531/Y 0.07fF
C1647 INVX1_LOC_12/Y INVX1_LOC_388/A 0.00fF
C1648 INPUT_5 INVX1_LOC_341/Y 0.05fF
C1649 NAND2X1_LOC_677/Y INVX1_LOC_479/A 0.03fF
C1650 INVX1_LOC_213/Y NAND2X1_LOC_495/a_36_24# 0.00fF
C1651 INVX1_LOC_677/A NAND2X1_LOC_451/B 0.01fF
C1652 NAND2X1_LOC_274/B INVX1_LOC_50/Y 0.07fF
C1653 INVX1_LOC_281/A INVX1_LOC_245/A 0.01fF
C1654 INVX1_LOC_513/A INVX1_LOC_119/Y 0.01fF
C1655 NAND2X1_LOC_184/Y NAND2X1_LOC_833/B 0.03fF
C1656 INVX1_LOC_293/A NAND2X1_LOC_359/a_36_24# 0.02fF
C1657 INVX1_LOC_153/Y NAND2X1_LOC_267/A 0.17fF
C1658 INVX1_LOC_566/A INVX1_LOC_636/A 0.75fF
C1659 INVX1_LOC_63/Y INVX1_LOC_361/A 0.12fF
C1660 INVX1_LOC_476/A NAND2X1_LOC_816/a_36_24# 0.00fF
C1661 INVX1_LOC_261/Y INVX1_LOC_245/A 0.12fF
C1662 INVX1_LOC_425/Y INVX1_LOC_75/Y 0.04fF
C1663 GATE_662 INVX1_LOC_655/A 0.03fF
C1664 INVX1_LOC_304/Y INVX1_LOC_364/A 0.03fF
C1665 INVX1_LOC_137/Y INVX1_LOC_645/Y 0.02fF
C1666 INVX1_LOC_199/Y INVX1_LOC_242/Y 0.07fF
C1667 NAND2X1_LOC_294/Y NAND2X1_LOC_396/Y 0.02fF
C1668 NAND2X1_LOC_493/a_36_24# INVX1_LOC_9/Y 0.00fF
C1669 INVX1_LOC_6/Y NAND2X1_LOC_629/a_36_24# 0.00fF
C1670 NAND2X1_LOC_846/B INVX1_LOC_655/A 0.08fF
C1671 INVX1_LOC_89/Y INVX1_LOC_479/A 1.28fF
C1672 NAND2X1_LOC_192/A INVX1_LOC_79/A 0.01fF
C1673 INVX1_LOC_376/Y INVX1_LOC_114/A 0.14fF
C1674 INVX1_LOC_120/Y INVX1_LOC_62/Y 0.01fF
C1675 INVX1_LOC_520/Y NAND2X1_LOC_843/B 0.17fF
C1676 INVX1_LOC_20/Y INVX1_LOC_109/Y 0.03fF
C1677 NAND2X1_LOC_319/a_36_24# INVX1_LOC_479/A 0.01fF
C1678 INVX1_LOC_301/Y INVX1_LOC_41/Y 0.03fF
C1679 VDD NAND2X1_LOC_749/Y 0.15fF
C1680 INVX1_LOC_46/Y NAND2X1_LOC_416/B 0.01fF
C1681 INVX1_LOC_567/A NAND2X1_LOC_513/Y 0.04fF
C1682 INVX1_LOC_459/A INVX1_LOC_45/Y 0.01fF
C1683 INVX1_LOC_501/A INVX1_LOC_479/A 0.10fF
C1684 NAND2X1_LOC_525/Y VDD 0.04fF
C1685 INVX1_LOC_20/Y INVX1_LOC_95/Y 0.01fF
C1686 VDD INVX1_LOC_583/Y 0.21fF
C1687 INVX1_LOC_100/Y INVX1_LOC_74/Y 7.94fF
C1688 INVX1_LOC_20/Y INVX1_LOC_554/A 0.00fF
C1689 INVX1_LOC_560/Y INVX1_LOC_51/Y 0.00fF
C1690 INVX1_LOC_100/Y INVX1_LOC_483/Y 0.01fF
C1691 VDD INVX1_LOC_167/Y 0.06fF
C1692 NAND2X1_LOC_299/Y INVX1_LOC_638/A 0.10fF
C1693 INVX1_LOC_270/A NAND2X1_LOC_76/B 0.02fF
C1694 NAND2X1_LOC_368/a_36_24# INVX1_LOC_51/Y 0.00fF
C1695 INVX1_LOC_574/A NAND2X1_LOC_152/Y 0.01fF
C1696 INVX1_LOC_374/A INVX1_LOC_355/A 0.02fF
C1697 INVX1_LOC_479/A NAND2X1_LOC_544/B 0.03fF
C1698 INVX1_LOC_174/Y INVX1_LOC_395/A 0.03fF
C1699 NAND2X1_LOC_503/B INVX1_LOC_600/A 0.17fF
C1700 INVX1_LOC_79/A INVX1_LOC_636/A 0.07fF
C1701 NAND2X1_LOC_69/B NAND2X1_LOC_378/Y 0.01fF
C1702 INVX1_LOC_68/Y INVX1_LOC_273/A 0.00fF
C1703 INPUT_6 INVX1_LOC_6/A 0.32fF
C1704 INVX1_LOC_402/A INPUT_0 0.00fF
C1705 INVX1_LOC_84/A INVX1_LOC_51/Y 1.72fF
C1706 VDD INVX1_LOC_137/Y 1.14fF
C1707 INVX1_LOC_127/A NAND2X1_LOC_130/Y 0.01fF
C1708 GATE_741 INVX1_LOC_522/Y 0.03fF
C1709 NAND2X1_LOC_710/A INVX1_LOC_586/A 0.03fF
C1710 NAND2X1_LOC_438/a_36_24# INVX1_LOC_92/A 0.00fF
C1711 NAND2X1_LOC_548/B INVX1_LOC_45/Y 0.01fF
C1712 INVX1_LOC_250/Y INVX1_LOC_249/Y 0.09fF
C1713 INVX1_LOC_425/A INVX1_LOC_119/A 0.06fF
C1714 INVX1_LOC_412/Y INVX1_LOC_252/Y 0.03fF
C1715 NAND2X1_LOC_271/B NAND2X1_LOC_275/Y 0.03fF
C1716 INVX1_LOC_586/A NAND2X1_LOC_541/B 0.07fF
C1717 INVX1_LOC_45/Y INVX1_LOC_635/A 0.02fF
C1718 INVX1_LOC_516/Y INVX1_LOC_508/Y 0.00fF
C1719 INVX1_LOC_291/A NAND2X1_LOC_357/a_36_24# 0.02fF
C1720 INVX1_LOC_20/Y INVX1_LOC_126/Y 0.02fF
C1721 NAND2X1_LOC_122/Y NAND2X1_LOC_302/A 0.02fF
C1722 INVX1_LOC_45/Y NAND2X1_LOC_237/Y 0.24fF
C1723 NAND2X1_LOC_143/a_36_24# INVX1_LOC_412/A 0.00fF
C1724 INVX1_LOC_608/Y INVX1_LOC_428/A 0.03fF
C1725 VDD INVX1_LOC_355/Y 0.16fF
C1726 INVX1_LOC_587/Y INVX1_LOC_206/Y 0.03fF
C1727 INVX1_LOC_428/A INVX1_LOC_17/Y 0.07fF
C1728 INPUT_3 NAND2X1_LOC_548/B 0.43fF
C1729 INVX1_LOC_169/A INVX1_LOC_369/A 0.03fF
C1730 VDD NAND2X1_LOC_829/B 0.01fF
C1731 INVX1_LOC_301/A INVX1_LOC_199/Y 0.07fF
C1732 INVX1_LOC_166/A NAND2X1_LOC_710/B 0.02fF
C1733 INVX1_LOC_98/A INVX1_LOC_98/Y 0.08fF
C1734 INVX1_LOC_243/A INVX1_LOC_381/A 0.07fF
C1735 NAND2X1_LOC_467/A INVX1_LOC_358/Y 0.00fF
C1736 INVX1_LOC_80/A INVX1_LOC_197/A 0.03fF
C1737 NAND2X1_LOC_780/A INVX1_LOC_610/A 0.09fF
C1738 INVX1_LOC_76/Y INVX1_LOC_98/Y 0.12fF
C1739 INVX1_LOC_134/A INVX1_LOC_159/Y 0.03fF
C1740 INVX1_LOC_560/A INVX1_LOC_317/A 0.03fF
C1741 NAND2X1_LOC_498/Y INVX1_LOC_670/A 0.12fF
C1742 VDD INPUT_5 0.57fF
C1743 INVX1_LOC_554/A INVX1_LOC_655/A 0.05fF
C1744 INVX1_LOC_564/A NAND2X1_LOC_753/Y 0.01fF
C1745 INVX1_LOC_435/Y INVX1_LOC_387/Y 0.05fF
C1746 INVX1_LOC_596/A INVX1_LOC_363/Y 0.03fF
C1747 INVX1_LOC_588/Y INVX1_LOC_577/Y 0.05fF
C1748 INVX1_LOC_558/A INVX1_LOC_520/A 0.04fF
C1749 NAND2X1_LOC_513/Y INVX1_LOC_6/Y 0.10fF
C1750 INVX1_LOC_356/A INVX1_LOC_505/A 0.15fF
C1751 VDD INVX1_LOC_2/Y 0.21fF
C1752 INVX1_LOC_250/Y INVX1_LOC_248/Y 0.03fF
C1753 NAND2X1_LOC_331/A INVX1_LOC_513/Y 0.26fF
C1754 INVX1_LOC_523/A NAND2X1_LOC_611/a_36_24# 0.00fF
C1755 INVX1_LOC_80/A NAND2X1_LOC_285/B 0.02fF
C1756 NAND2X1_LOC_107/Y INVX1_LOC_145/Y 0.10fF
C1757 NAND2X1_LOC_768/A NAND2X1_LOC_285/B 0.05fF
C1758 INVX1_LOC_206/Y INVX1_LOC_9/Y 1.33fF
C1759 INVX1_LOC_435/Y INVX1_LOC_49/Y 0.10fF
C1760 INVX1_LOC_11/Y INVX1_LOC_197/A 0.07fF
C1761 INVX1_LOC_80/A NAND2X1_LOC_106/B 0.10fF
C1762 NAND2X1_LOC_768/A NAND2X1_LOC_106/B 0.14fF
C1763 INVX1_LOC_603/Y INVX1_LOC_35/Y 0.03fF
C1764 INVX1_LOC_544/A INVX1_LOC_680/Y 0.01fF
C1765 INVX1_LOC_648/Y INVX1_LOC_9/Y 0.02fF
C1766 INVX1_LOC_586/A INVX1_LOC_149/Y 0.04fF
C1767 NAND2X1_LOC_498/B INVX1_LOC_338/Y 0.07fF
C1768 INVX1_LOC_377/Y INVX1_LOC_670/A 0.03fF
C1769 INVX1_LOC_53/Y INVX1_LOC_598/A 0.02fF
C1770 NAND2X1_LOC_122/Y NAND2X1_LOC_637/a_36_24# 0.00fF
C1771 NAND2X1_LOC_174/B INVX1_LOC_579/Y 0.03fF
C1772 INVX1_LOC_572/Y NAND2X1_LOC_728/B 0.12fF
C1773 INVX1_LOC_585/Y INVX1_LOC_12/Y 0.05fF
C1774 INVX1_LOC_110/A INVX1_LOC_134/Y 0.05fF
C1775 INVX1_LOC_76/Y INVX1_LOC_338/Y 1.24fF
C1776 INVX1_LOC_20/Y INVX1_LOC_199/Y 0.12fF
C1777 NAND2X1_LOC_325/B INVX1_LOC_105/A 0.03fF
C1778 INVX1_LOC_377/A INPUT_1 0.02fF
C1779 NAND2X1_LOC_591/Y INVX1_LOC_579/Y 0.02fF
C1780 INVX1_LOC_575/A INVX1_LOC_492/A 0.00fF
C1781 INVX1_LOC_213/Y INVX1_LOC_145/Y 0.06fF
C1782 INVX1_LOC_206/Y INVX1_LOC_62/Y 0.18fF
C1783 INVX1_LOC_137/Y INVX1_LOC_509/A 0.00fF
C1784 NAND2X1_LOC_595/Y INPUT_1 0.00fF
C1785 VDD NAND2X1_LOC_234/Y 0.20fF
C1786 INVX1_LOC_530/A INVX1_LOC_46/Y 0.00fF
C1787 VDD INVX1_LOC_647/Y 0.21fF
C1788 INVX1_LOC_53/Y NAND2X1_LOC_128/B 0.01fF
C1789 NAND2X1_LOC_140/B INVX1_LOC_105/Y 0.13fF
C1790 INVX1_LOC_629/A INVX1_LOC_74/Y 0.01fF
C1791 NAND2X1_LOC_837/B NAND2X1_LOC_826/a_36_24# 0.02fF
C1792 INVX1_LOC_9/Y INVX1_LOC_242/A 0.03fF
C1793 INVX1_LOC_596/A INVX1_LOC_49/Y 0.07fF
C1794 INPUT_0 INVX1_LOC_653/Y 0.00fF
C1795 INVX1_LOC_558/A INVX1_LOC_519/Y 0.01fF
C1796 NAND2X1_LOC_501/a_36_24# INVX1_LOC_100/Y 0.01fF
C1797 INVX1_LOC_89/Y INVX1_LOC_12/Y 0.10fF
C1798 INVX1_LOC_395/A INVX1_LOC_135/Y 0.05fF
C1799 INVX1_LOC_517/A INVX1_LOC_58/Y 0.01fF
C1800 INVX1_LOC_413/A INVX1_LOC_392/A 0.08fF
C1801 INVX1_LOC_17/Y INVX1_LOC_359/Y 0.01fF
C1802 INVX1_LOC_206/Y INVX1_LOC_529/Y 0.03fF
C1803 INPUT_0 INVX1_LOC_666/Y 0.07fF
C1804 INVX1_LOC_372/Y INVX1_LOC_501/A 0.03fF
C1805 INVX1_LOC_418/Y INVX1_LOC_50/Y 0.04fF
C1806 NAND2X1_LOC_387/Y INVX1_LOC_35/Y 0.10fF
C1807 NAND2X1_LOC_638/A INVX1_LOC_659/A 0.07fF
C1808 INVX1_LOC_686/A INVX1_LOC_9/Y 0.07fF
C1809 NAND2X1_LOC_708/A INVX1_LOC_189/A 0.04fF
C1810 INVX1_LOC_183/A INVX1_LOC_324/A 0.01fF
C1811 INVX1_LOC_54/Y NAND2X1_LOC_615/B 0.03fF
C1812 INVX1_LOC_381/A INVX1_LOC_79/A 0.07fF
C1813 INVX1_LOC_99/Y NAND2X1_LOC_606/a_36_24# 0.00fF
C1814 NAND2X1_LOC_516/Y INVX1_LOC_666/Y 0.10fF
C1815 INVX1_LOC_344/Y INVX1_LOC_675/A -0.00fF
C1816 INVX1_LOC_100/A NAND2X1_LOC_673/B 0.04fF
C1817 INVX1_LOC_300/A INVX1_LOC_199/Y 0.73fF
C1818 INVX1_LOC_320/A NAND2X1_LOC_558/B 0.17fF
C1819 INVX1_LOC_381/A NAND2X1_LOC_631/B 0.12fF
C1820 INVX1_LOC_197/A NAND2X1_LOC_433/Y 0.07fF
C1821 INVX1_LOC_221/Y INVX1_LOC_283/A 0.65fF
C1822 INVX1_LOC_504/A INVX1_LOC_49/Y 0.08fF
C1823 INVX1_LOC_468/Y INVX1_LOC_624/Y 0.73fF
C1824 NAND2X1_LOC_698/Y INVX1_LOC_145/Y 0.01fF
C1825 INVX1_LOC_649/A NAND2X1_LOC_819/a_36_24# 0.02fF
C1826 INVX1_LOC_439/Y INVX1_LOC_433/A 0.09fF
C1827 INVX1_LOC_17/Y NAND2X1_LOC_52/a_36_24# 0.00fF
C1828 INVX1_LOC_577/A INVX1_LOC_636/A 0.02fF
C1829 NAND2X1_LOC_387/Y INVX1_LOC_620/A 0.07fF
C1830 INVX1_LOC_54/Y INVX1_LOC_66/A 0.06fF
C1831 INVX1_LOC_255/A INVX1_LOC_349/A 0.05fF
C1832 INVX1_LOC_320/A INVX1_LOC_79/A 0.01fF
C1833 INVX1_LOC_566/A INVX1_LOC_74/Y 0.08fF
C1834 INVX1_LOC_686/A INVX1_LOC_62/Y 0.14fF
C1835 NAND2X1_LOC_841/a_36_24# INVX1_LOC_99/Y 0.00fF
C1836 INVX1_LOC_47/Y INVX1_LOC_670/A 0.24fF
C1837 INVX1_LOC_35/Y NAND2X1_LOC_845/B 0.00fF
C1838 INVX1_LOC_117/Y INVX1_LOC_77/Y 0.13fF
C1839 NAND2X1_LOC_27/a_36_24# NAND2X1_LOC_557/B 0.01fF
C1840 INVX1_LOC_7/Y INVX1_LOC_90/Y 0.00fF
C1841 INVX1_LOC_358/Y INVX1_LOC_41/Y 0.04fF
C1842 INVX1_LOC_335/Y INVX1_LOC_41/Y 0.04fF
C1843 INVX1_LOC_21/Y INVX1_LOC_41/Y 0.25fF
C1844 NAND2X1_LOC_301/B INVX1_LOC_506/Y 0.59fF
C1845 NAND2X1_LOC_520/a_36_24# INVX1_LOC_502/A 0.01fF
C1846 INVX1_LOC_628/A INVX1_LOC_74/Y 0.01fF
C1847 INVX1_LOC_54/Y INVX1_LOC_178/Y 0.09fF
C1848 INVX1_LOC_32/Y INVX1_LOC_351/A 0.00fF
C1849 INVX1_LOC_588/Y INVX1_LOC_26/Y 0.02fF
C1850 INVX1_LOC_102/Y NAND2X1_LOC_106/B 0.20fF
C1851 INVX1_LOC_167/A NAND2X1_LOC_633/a_36_24# 0.01fF
C1852 INVX1_LOC_6/Y NAND2X1_LOC_615/Y 0.02fF
C1853 INVX1_LOC_79/A NAND2X1_LOC_720/A 0.07fF
C1854 INVX1_LOC_592/Y INVX1_LOC_44/Y 0.05fF
C1855 INVX1_LOC_63/Y NAND2X1_LOC_449/B 0.04fF
C1856 INVX1_LOC_501/A INVX1_LOC_188/A 0.03fF
C1857 INVX1_LOC_670/A INVX1_LOC_119/Y 0.09fF
C1858 INVX1_LOC_32/Y INVX1_LOC_90/Y 0.21fF
C1859 INVX1_LOC_58/Y NAND2X1_LOC_847/A 0.01fF
C1860 INVX1_LOC_681/Y NAND2X1_LOC_372/Y 0.07fF
C1861 INVX1_LOC_42/Y NAND2X1_LOC_85/a_36_24# 0.00fF
C1862 INVX1_LOC_41/Y NAND2X1_LOC_267/A 0.13fF
C1863 INVX1_LOC_47/Y NAND2X1_LOC_832/a_36_24# 0.01fF
C1864 NAND2X1_LOC_111/Y INVX1_LOC_128/Y 0.00fF
C1865 INPUT_1 NAND2X1_LOC_372/Y 0.03fF
C1866 INVX1_LOC_199/Y INVX1_LOC_655/A 0.16fF
C1867 NAND2X1_LOC_833/B NAND2X1_LOC_259/a_36_24# 0.00fF
C1868 INVX1_LOC_167/A INVX1_LOC_588/A 0.01fF
C1869 INVX1_LOC_469/Y INVX1_LOC_74/Y 0.10fF
C1870 INVX1_LOC_6/Y INVX1_LOC_614/Y 0.01fF
C1871 INVX1_LOC_67/Y INVX1_LOC_92/A 0.31fF
C1872 INVX1_LOC_482/Y INVX1_LOC_245/A 0.03fF
C1873 NAND2X1_LOC_301/B INVX1_LOC_63/Y 0.25fF
C1874 NAND2X1_LOC_435/a_36_24# NAND2X1_LOC_832/A 0.00fF
C1875 NAND2X1_LOC_123/B INVX1_LOC_347/Y 0.00fF
C1876 INVX1_LOC_169/Y NAND2X1_LOC_619/a_36_24# 0.01fF
C1877 INVX1_LOC_279/Y INVX1_LOC_445/A 0.03fF
C1878 NAND2X1_LOC_753/Y INVX1_LOC_91/Y 0.18fF
C1879 INVX1_LOC_100/Y INVX1_LOC_79/A 0.22fF
C1880 INVX1_LOC_531/Y INVX1_LOC_26/Y 0.04fF
C1881 INVX1_LOC_465/Y INVX1_LOC_45/Y 0.01fF
C1882 INVX1_LOC_77/A INVX1_LOC_74/Y 0.02fF
C1883 INVX1_LOC_100/Y NAND2X1_LOC_396/Y 0.01fF
C1884 INVX1_LOC_47/Y NAND2X1_LOC_418/a_36_24# 0.01fF
C1885 INPUT_0 INVX1_LOC_490/Y 0.03fF
C1886 INVX1_LOC_133/Y NAND2X1_LOC_820/Y 0.01fF
C1887 INVX1_LOC_79/A INVX1_LOC_74/Y 0.68fF
C1888 INVX1_LOC_596/A INVX1_LOC_297/Y 0.00fF
C1889 INVX1_LOC_479/A INVX1_LOC_461/Y 0.16fF
C1890 INVX1_LOC_62/Y NAND2X1_LOC_609/B 0.03fF
C1891 INVX1_LOC_177/Y INVX1_LOC_395/A 0.03fF
C1892 INVX1_LOC_566/A NAND2X1_LOC_591/B 0.03fF
C1893 INVX1_LOC_682/Y NAND2X1_LOC_457/a_36_24# -0.01fF
C1894 INPUT_0 NAND2X1_LOC_16/Y 0.19fF
C1895 INVX1_LOC_74/Y INVX1_LOC_460/A 0.01fF
C1896 NAND2X1_LOC_318/A NAND2X1_LOC_76/B 0.03fF
C1897 NAND2X1_LOC_475/A NAND2X1_LOC_391/B 0.02fF
C1898 INVX1_LOC_84/A NAND2X1_LOC_537/A 0.00fF
C1899 INVX1_LOC_425/A INVX1_LOC_410/Y 0.37fF
C1900 INVX1_LOC_301/A INVX1_LOC_53/Y 0.03fF
C1901 INVX1_LOC_119/Y NAND2X1_LOC_418/a_36_24# 0.00fF
C1902 VDD NAND2X1_LOC_307/A 0.19fF
C1903 NAND2X1_LOC_271/B INVX1_LOC_235/Y 0.01fF
C1904 VDD INVX1_LOC_545/Y 0.43fF
C1905 INVX1_LOC_3/Y INVX1_LOC_29/Y 0.06fF
C1906 INVX1_LOC_211/A INVX1_LOC_666/Y 0.02fF
C1907 INVX1_LOC_45/Y INVX1_LOC_666/A 0.00fF
C1908 INVX1_LOC_580/A INVX1_LOC_577/Y 0.01fF
C1909 INVX1_LOC_340/Y NAND2X1_LOC_426/Y 0.02fF
C1910 INVX1_LOC_65/Y INVX1_LOC_270/A 0.07fF
C1911 INVX1_LOC_628/A INVX1_LOC_629/A -0.00fF
C1912 NAND2X1_LOC_43/a_36_24# INVX1_LOC_11/Y 0.00fF
C1913 INVX1_LOC_202/Y NAND2X1_LOC_76/B 0.17fF
C1914 NAND2X1_LOC_142/Y INVX1_LOC_651/A 0.14fF
C1915 INVX1_LOC_185/Y INVX1_LOC_492/Y 0.28fF
C1916 NAND2X1_LOC_45/Y INVX1_LOC_435/A 0.10fF
C1917 VDD INVX1_LOC_419/Y 0.26fF
C1918 NAND2X1_LOC_613/Y INVX1_LOC_235/Y 0.02fF
C1919 INVX1_LOC_590/Y INVX1_LOC_97/Y 0.05fF
C1920 INVX1_LOC_510/Y NAND2X1_LOC_307/A 0.07fF
C1921 INVX1_LOC_51/A INVX1_LOC_17/Y 0.00fF
C1922 INVX1_LOC_295/A INVX1_LOC_482/A 0.13fF
C1923 NAND2X1_LOC_13/Y INVX1_LOC_84/A 0.07fF
C1924 INVX1_LOC_438/A INVX1_LOC_159/Y 0.04fF
C1925 INVX1_LOC_530/Y INVX1_LOC_530/A 0.14fF
C1926 NAND2X1_LOC_249/Y INVX1_LOC_166/A 0.06fF
C1927 NAND2X1_LOC_69/B INVX1_LOC_6/Y 0.43fF
C1928 INVX1_LOC_596/A INVX1_LOC_76/Y 0.00fF
C1929 INVX1_LOC_308/Y NAND2X1_LOC_673/B 0.03fF
C1930 NAND2X1_LOC_98/a_36_24# INVX1_LOC_50/Y 0.00fF
C1931 INVX1_LOC_375/A INVX1_LOC_252/Y 0.05fF
C1932 INVX1_LOC_191/Y NAND2X1_LOC_789/A 0.31fF
C1933 INVX1_LOC_400/Y INVX1_LOC_400/A 0.05fF
C1934 INPUT_0 INVX1_LOC_431/A 0.00fF
C1935 INVX1_LOC_20/Y INVX1_LOC_53/Y 0.19fF
C1936 INVX1_LOC_224/Y NAND2X1_LOC_265/a_36_24# 0.00fF
C1937 INVX1_LOC_425/Y INVX1_LOC_578/A 0.04fF
C1938 INVX1_LOC_629/A INVX1_LOC_469/Y 0.00fF
C1939 NAND2X1_LOC_379/a_36_24# INVX1_LOC_366/A 0.00fF
C1940 INVX1_LOC_84/A INVX1_LOC_27/A 0.31fF
C1941 VDD NAND2X1_LOC_342/A 0.00fF
C1942 INVX1_LOC_556/A INVX1_LOC_118/A 0.09fF
C1943 NAND2X1_LOC_756/Y NAND2X1_LOC_237/Y 0.01fF
C1944 NAND2X1_LOC_673/A INVX1_LOC_45/Y 0.01fF
C1945 INVX1_LOC_17/Y NAND2X1_LOC_173/Y 0.01fF
C1946 INVX1_LOC_269/Y INVX1_LOC_48/Y 0.03fF
C1947 INVX1_LOC_54/Y INVX1_LOC_442/A 0.07fF
C1948 INVX1_LOC_413/A INVX1_LOC_362/Y 0.02fF
C1949 INVX1_LOC_344/A INVX1_LOC_686/A 0.03fF
C1950 INVX1_LOC_400/Y INVX1_LOC_93/Y 0.07fF
C1951 NAND2X1_LOC_97/B INVX1_LOC_80/A 0.28fF
C1952 INVX1_LOC_160/Y NAND2X1_LOC_267/A 0.32fF
C1953 NAND2X1_LOC_130/Y INVX1_LOC_519/A 0.00fF
C1954 INVX1_LOC_65/Y INVX1_LOC_46/Y 0.01fF
C1955 INVX1_LOC_584/A INVX1_LOC_675/A 0.02fF
C1956 INVX1_LOC_335/Y INVX1_LOC_358/Y 0.01fF
C1957 INVX1_LOC_288/A INVX1_LOC_561/A 0.04fF
C1958 INVX1_LOC_381/A INVX1_LOC_48/Y 0.07fF
C1959 INVX1_LOC_300/A INVX1_LOC_53/Y 0.07fF
C1960 INVX1_LOC_556/Y INVX1_LOC_337/Y 0.26fF
C1961 NAND2X1_LOC_179/Y INVX1_LOC_80/A 0.11fF
C1962 INVX1_LOC_605/Y INVX1_LOC_35/Y 0.02fF
C1963 INVX1_LOC_139/A INVX1_LOC_338/Y 0.01fF
C1964 INVX1_LOC_185/Y NAND2X1_LOC_647/A 0.00fF
C1965 INVX1_LOC_442/A INVX1_LOC_257/A 0.86fF
C1966 NAND2X1_LOC_532/Y INVX1_LOC_51/Y 0.07fF
C1967 INVX1_LOC_80/A INVX1_LOC_510/A 0.07fF
C1968 NAND2X1_LOC_661/a_36_24# NAND2X1_LOC_679/B 0.00fF
C1969 INVX1_LOC_238/A NAND2X1_LOC_136/Y 0.02fF
C1970 NAND2X1_LOC_387/Y INVX1_LOC_291/A 0.01fF
C1971 INVX1_LOC_21/Y NAND2X1_LOC_655/a_36_24# 0.01fF
C1972 NAND2X1_LOC_488/Y INVX1_LOC_388/Y 0.03fF
C1973 INVX1_LOC_298/A INVX1_LOC_55/Y 0.00fF
C1974 INVX1_LOC_400/Y INVX1_LOC_390/A 0.03fF
C1975 INVX1_LOC_586/A INVX1_LOC_493/Y 0.18fF
C1976 NAND2X1_LOC_242/A INVX1_LOC_79/A 0.03fF
C1977 INVX1_LOC_320/A INVX1_LOC_48/Y 0.00fF
C1978 INVX1_LOC_490/A INVX1_LOC_235/Y 0.02fF
C1979 INVX1_LOC_568/Y INVX1_LOC_575/A 0.15fF
C1980 INVX1_LOC_185/Y INVX1_LOC_168/Y 0.02fF
C1981 INVX1_LOC_12/Y INVX1_LOC_194/Y 0.77fF
C1982 INVX1_LOC_184/A INVX1_LOC_46/Y 0.02fF
C1983 NAND2X1_LOC_513/Y INVX1_LOC_557/Y 0.02fF
C1984 INVX1_LOC_384/A NAND2X1_LOC_178/a_36_24# 0.01fF
C1985 INVX1_LOC_580/Y NAND2X1_LOC_334/A 0.13fF
C1986 INVX1_LOC_625/A INVX1_LOC_202/Y 0.02fF
C1987 INVX1_LOC_551/Y INVX1_LOC_253/Y 0.17fF
C1988 INVX1_LOC_679/A INVX1_LOC_145/Y 0.00fF
C1989 INVX1_LOC_449/A INPUT_1 0.04fF
C1990 INVX1_LOC_92/Y NAND2X1_LOC_76/B 0.01fF
C1991 NAND2X1_LOC_285/B NAND2X1_LOC_282/a_36_24# 0.02fF
C1992 INVX1_LOC_679/A INVX1_LOC_661/Y 0.02fF
C1993 NAND2X1_LOC_513/A NAND2X1_LOC_412/a_36_24# 0.01fF
C1994 INVX1_LOC_377/A INVX1_LOC_50/Y 0.01fF
C1995 INVX1_LOC_54/Y INVX1_LOC_305/Y 0.02fF
C1996 INVX1_LOC_80/A NAND2X1_LOC_128/A 0.03fF
C1997 INVX1_LOC_6/Y NAND2X1_LOC_541/B 0.43fF
C1998 INVX1_LOC_33/Y INVX1_LOC_35/A 0.00fF
C1999 INVX1_LOC_21/Y NAND2X1_LOC_267/A 0.07fF
C2000 NAND2X1_LOC_595/Y INVX1_LOC_50/Y 0.00fF
C2001 INVX1_LOC_551/Y INVX1_LOC_63/Y 0.04fF
C2002 NAND2X1_LOC_707/A INVX1_LOC_245/A 0.12fF
C2003 INVX1_LOC_374/A NAND2X1_LOC_301/B 0.01fF
C2004 INVX1_LOC_628/A INVX1_LOC_469/Y -0.00fF
C2005 INVX1_LOC_632/A NAND2X1_LOC_638/a_36_24# 0.00fF
C2006 INVX1_LOC_11/Y INVX1_LOC_510/A 0.01fF
C2007 INVX1_LOC_31/Y INVX1_LOC_344/Y 0.02fF
C2008 INVX1_LOC_686/A INVX1_LOC_624/Y 0.01fF
C2009 INVX1_LOC_54/Y INVX1_LOC_116/Y 0.12fF
C2010 INVX1_LOC_207/A INVX1_LOC_79/A 0.12fF
C2011 NAND2X1_LOC_720/A INVX1_LOC_59/Y 0.01fF
C2012 INVX1_LOC_580/A INVX1_LOC_26/Y 0.02fF
C2013 INVX1_LOC_390/Y INVX1_LOC_62/Y 0.23fF
C2014 NAND2X1_LOC_493/B INVX1_LOC_245/A 0.01fF
C2015 INVX1_LOC_117/Y INVX1_LOC_549/Y 0.01fF
C2016 INVX1_LOC_255/Y INVX1_LOC_41/Y 0.03fF
C2017 INVX1_LOC_333/Y INVX1_LOC_93/A 0.01fF
C2018 INVX1_LOC_304/Y INVX1_LOC_295/Y 0.01fF
C2019 INVX1_LOC_32/Y INVX1_LOC_98/Y 0.35fF
C2020 INVX1_LOC_93/Y INVX1_LOC_125/A 0.01fF
C2021 VDD INVX1_LOC_623/A -0.00fF
C2022 NAND2X1_LOC_635/B INVX1_LOC_259/Y 0.01fF
C2023 NAND2X1_LOC_307/B NAND2X1_LOC_413/Y 0.07fF
C2024 INVX1_LOC_301/Y NAND2X1_LOC_865/a_36_24# 0.00fF
C2025 NAND2X1_LOC_174/B NAND2X1_LOC_172/a_36_24# 0.01fF
C2026 INVX1_LOC_12/Y INVX1_LOC_44/Y 0.03fF
C2027 INVX1_LOC_566/A INVX1_LOC_79/A 0.03fF
C2028 INVX1_LOC_257/A INVX1_LOC_116/Y 0.51fF
C2029 INVX1_LOC_145/Y NAND2X1_LOC_258/Y 1.19fF
C2030 INVX1_LOC_174/A INVX1_LOC_223/Y 0.11fF
C2031 INVX1_LOC_435/A INVX1_LOC_47/Y 0.03fF
C2032 INVX1_LOC_261/Y INVX1_LOC_678/A 0.02fF
C2033 INVX1_LOC_65/Y INVX1_LOC_75/A 0.06fF
C2034 NAND2X1_LOC_388/A INVX1_LOC_159/Y 0.11fF
C2035 INVX1_LOC_53/Y INVX1_LOC_655/A 0.17fF
C2036 INVX1_LOC_421/A INVX1_LOC_93/Y 0.07fF
C2037 INVX1_LOC_654/A INVX1_LOC_62/Y 0.03fF
C2038 NAND2X1_LOC_317/A INVX1_LOC_92/A 0.05fF
C2039 INVX1_LOC_69/Y INVX1_LOC_349/A 0.01fF
C2040 NAND2X1_LOC_106/Y INVX1_LOC_105/Y 0.01fF
C2041 INVX1_LOC_561/Y INVX1_LOC_636/A 0.02fF
C2042 INVX1_LOC_384/A INVX1_LOC_666/Y 0.01fF
C2043 NAND2X1_LOC_333/B NAND2X1_LOC_753/Y 0.09fF
C2044 INVX1_LOC_54/Y INVX1_LOC_255/A 0.03fF
C2045 INVX1_LOC_312/A NAND2X1_LOC_528/Y 0.00fF
C2046 INVX1_LOC_417/Y INVX1_LOC_100/Y 0.03fF
C2047 INVX1_LOC_261/Y INVX1_LOC_686/Y 0.01fF
C2048 INVX1_LOC_66/A INVX1_LOC_199/A 0.01fF
C2049 INVX1_LOC_432/A INVX1_LOC_9/Y 0.03fF
C2050 INVX1_LOC_633/A INVX1_LOC_6/Y 0.01fF
C2051 INVX1_LOC_80/A NAND2X1_LOC_248/B 0.07fF
C2052 INVX1_LOC_89/Y INVX1_LOC_66/A 0.20fF
C2053 INVX1_LOC_80/A INVX1_LOC_66/Y 0.01fF
C2054 INVX1_LOC_134/Y INVX1_LOC_75/Y 0.07fF
C2055 NAND2X1_LOC_768/A NAND2X1_LOC_248/B 0.00fF
C2056 INVX1_LOC_32/Y INVX1_LOC_338/Y 0.02fF
C2057 INVX1_LOC_398/Y INVX1_LOC_100/Y 0.01fF
C2058 INVX1_LOC_100/Y INVX1_LOC_59/Y 0.06fF
C2059 INVX1_LOC_89/Y INVX1_LOC_296/A 0.09fF
C2060 INVX1_LOC_328/Y INPUT_1 0.06fF
C2061 INVX1_LOC_632/A INVX1_LOC_74/Y 0.07fF
C2062 INVX1_LOC_117/A NAND2X1_LOC_84/B 0.05fF
C2063 INVX1_LOC_63/Y NAND2X1_LOC_252/Y 0.02fF
C2064 INVX1_LOC_509/Y INVX1_LOC_74/Y 0.01fF
C2065 NAND2X1_LOC_398/a_36_24# INVX1_LOC_11/A 0.00fF
C2066 INPUT_1 INVX1_LOC_518/A 0.01fF
C2067 INVX1_LOC_21/Y INVX1_LOC_209/Y 0.01fF
C2068 INVX1_LOC_97/Y INVX1_LOC_211/A 0.13fF
C2069 INVX1_LOC_619/A NAND2X1_LOC_234/Y 0.02fF
C2070 INVX1_LOC_69/Y INVX1_LOC_420/A 0.07fF
C2071 INVX1_LOC_17/Y NAND2X1_LOC_488/Y 0.06fF
C2072 INVX1_LOC_117/Y NAND2X1_LOC_274/B 0.03fF
C2073 INVX1_LOC_448/A INVX1_LOC_666/Y 0.02fF
C2074 INVX1_LOC_479/A NAND2X1_LOC_418/Y 0.03fF
C2075 INVX1_LOC_100/Y INVX1_LOC_48/Y 0.26fF
C2076 INVX1_LOC_58/Y INVX1_LOC_77/Y 0.27fF
C2077 NAND2X1_LOC_285/B NAND2X1_LOC_843/B 0.02fF
C2078 NAND2X1_LOC_409/Y INVX1_LOC_40/Y 0.01fF
C2079 INVX1_LOC_59/Y INVX1_LOC_74/Y 0.03fF
C2080 INVX1_LOC_17/Y INVX1_LOC_354/A 0.00fF
C2081 INVX1_LOC_17/Y INVX1_LOC_441/A 0.00fF
C2082 INVX1_LOC_103/Y INVX1_LOC_502/A 0.03fF
C2083 INVX1_LOC_79/A INVX1_LOC_350/Y 0.00fF
C2084 INVX1_LOC_63/Y NAND2X1_LOC_759/Y 0.01fF
C2085 NAND2X1_LOC_386/a_36_24# INVX1_LOC_74/Y 0.01fF
C2086 INVX1_LOC_62/Y INVX1_LOC_432/A 0.01fF
C2087 NAND2X1_LOC_106/B NAND2X1_LOC_843/B 0.02fF
C2088 INVX1_LOC_496/A INVX1_LOC_196/Y 0.03fF
C2089 NAND2X1_LOC_542/A INVX1_LOC_9/Y 0.04fF
C2090 INVX1_LOC_399/Y INVX1_LOC_69/Y 0.00fF
C2091 NAND2X1_LOC_686/A INVX1_LOC_49/Y 0.00fF
C2092 INVX1_LOC_50/Y INVX1_LOC_280/A 0.03fF
C2093 INVX1_LOC_50/Y NAND2X1_LOC_372/Y 0.03fF
C2094 INVX1_LOC_469/Y INVX1_LOC_460/A 0.01fF
C2095 INVX1_LOC_74/Y INVX1_LOC_48/Y 0.12fF
C2096 INVX1_LOC_386/Y NAND2X1_LOC_416/B 0.73fF
C2097 INVX1_LOC_483/Y INVX1_LOC_48/Y 0.05fF
C2098 NAND2X1_LOC_424/a_36_24# INVX1_LOC_114/A 0.01fF
C2099 INVX1_LOC_89/Y NAND2X1_LOC_601/Y 0.04fF
C2100 INPUT_0 INVX1_LOC_615/A 0.26fF
C2101 INVX1_LOC_46/Y INVX1_LOC_588/A 0.00fF
C2102 VDD INVX1_LOC_388/Y 0.21fF
C2103 NAND2X1_LOC_491/Y INVX1_LOC_100/Y 0.01fF
C2104 INVX1_LOC_235/A NAND2X1_LOC_271/A 0.04fF
C2105 INVX1_LOC_74/A INVX1_LOC_93/A 0.20fF
C2106 INVX1_LOC_300/A INVX1_LOC_636/Y 0.03fF
C2107 NAND2X1_LOC_544/B INVX1_LOC_66/A 0.01fF
C2108 NAND2X1_LOC_558/B INVX1_LOC_79/A 0.00fF
C2109 INVX1_LOC_434/A NAND2X1_LOC_560/a_36_24# 0.02fF
C2110 INVX1_LOC_652/A INVX1_LOC_114/A 0.00fF
C2111 NAND2X1_LOC_528/Y INVX1_LOC_226/Y 0.05fF
C2112 INVX1_LOC_41/Y INVX1_LOC_26/Y 1.64fF
C2113 INVX1_LOC_41/Y INVX1_LOC_128/Y 0.00fF
C2114 NAND2X1_LOC_331/A INVX1_LOC_206/Y 0.03fF
C2115 NAND2X1_LOC_434/B INVX1_LOC_74/Y 0.02fF
C2116 INVX1_LOC_63/Y INVX1_LOC_634/Y 0.07fF
C2117 NAND2X1_LOC_249/Y INVX1_LOC_302/A 0.02fF
C2118 NAND2X1_LOC_88/a_36_24# INVX1_LOC_65/Y 0.00fF
C2119 NAND2X1_LOC_45/Y INVX1_LOC_392/Y 0.04fF
C2120 INVX1_LOC_76/Y NAND2X1_LOC_76/B 0.07fF
C2121 INVX1_LOC_400/Y INVX1_LOC_395/A 0.03fF
C2122 VDD INVX1_LOC_286/Y 0.41fF
C2123 NAND2X1_LOC_626/a_36_24# NAND2X1_LOC_626/Y 0.02fF
C2124 NAND2X1_LOC_846/B INVX1_LOC_92/A 0.02fF
C2125 INVX1_LOC_546/Y NAND2X1_LOC_498/Y 0.01fF
C2126 INVX1_LOC_462/Y INVX1_LOC_114/A 0.16fF
C2127 INVX1_LOC_201/A INVX1_LOC_615/A 0.34fF
C2128 NAND2X1_LOC_373/Y INVX1_LOC_53/Y 0.12fF
C2129 INVX1_LOC_554/A INVX1_LOC_567/Y 0.03fF
C2130 INVX1_LOC_577/A INVX1_LOC_566/A 0.07fF
C2131 NAND2X1_LOC_45/Y INVX1_LOC_367/A 0.01fF
C2132 INVX1_LOC_412/Y INVX1_LOC_80/A 0.12fF
C2133 INVX1_LOC_65/Y NAND2X1_LOC_318/A 0.08fF
C2134 INVX1_LOC_68/Y NAND2X1_LOC_97/A 0.01fF
C2135 VDD INVX1_LOC_608/Y 0.21fF
C2136 VDD INVX1_LOC_503/A 0.00fF
C2137 VDD INVX1_LOC_17/Y 2.53fF
C2138 INVX1_LOC_267/Y INVX1_LOC_564/A 0.16fF
C2139 INPUT_0 INVX1_LOC_275/Y 0.01fF
C2140 INVX1_LOC_198/A INVX1_LOC_180/Y 0.02fF
C2141 INVX1_LOC_20/Y NAND2X1_LOC_383/Y 0.24fF
C2142 INVX1_LOC_435/A NAND2X1_LOC_475/A 0.04fF
C2143 NAND2X1_LOC_391/a_36_24# INVX1_LOC_84/A 0.00fF
C2144 NAND2X1_LOC_45/Y INVX1_LOC_392/A 0.10fF
C2145 VDD INVX1_LOC_650/Y 0.26fF
C2146 NAND2X1_LOC_317/B NAND2X1_LOC_307/a_36_24# 0.00fF
C2147 INVX1_LOC_490/Y INVX1_LOC_145/Y 0.24fF
C2148 GATE_741 INVX1_LOC_581/A 0.03fF
C2149 INVX1_LOC_11/Y INVX1_LOC_412/Y 0.03fF
C2150 INVX1_LOC_558/A INVX1_LOC_670/Y 0.00fF
C2151 INVX1_LOC_53/A INVX1_LOC_26/A 0.01fF
C2152 VDD INVX1_LOC_601/Y 0.46fF
C2153 INVX1_LOC_679/Y INVX1_LOC_651/Y 0.22fF
C2154 NAND2X1_LOC_45/Y INVX1_LOC_93/Y 5.12fF
C2155 INVX1_LOC_80/A INVX1_LOC_119/A 0.00fF
C2156 INVX1_LOC_617/Y INVX1_LOC_80/A 0.07fF
C2157 NAND2X1_LOC_788/A INVX1_LOC_89/Y 0.02fF
C2158 INVX1_LOC_166/A INVX1_LOC_122/Y 0.03fF
C2159 NAND2X1_LOC_854/a_36_24# INVX1_LOC_638/A 0.00fF
C2160 INVX1_LOC_202/Y INVX1_LOC_65/Y 0.03fF
C2161 INVX1_LOC_206/Y INVX1_LOC_169/Y 0.07fF
C2162 VDD NAND2X1_LOC_307/B 0.41fF
C2163 INVX1_LOC_185/Y INVX1_LOC_137/Y 0.03fF
C2164 INVX1_LOC_586/A INVX1_LOC_176/A 0.01fF
C2165 NAND2X1_LOC_383/Y INVX1_LOC_300/A 0.01fF
C2166 INVX1_LOC_290/Y INVX1_LOC_641/Y 0.03fF
C2167 INVX1_LOC_625/A INVX1_LOC_76/Y 0.02fF
C2168 INVX1_LOC_45/Y INVX1_LOC_137/Y 0.00fF
C2169 INVX1_LOC_324/A INVX1_LOC_324/Y 0.00fF
C2170 INVX1_LOC_11/Y INVX1_LOC_321/A 0.03fF
C2171 INVX1_LOC_586/A INVX1_LOC_349/A 0.01fF
C2172 INVX1_LOC_524/Y INVX1_LOC_99/Y 0.03fF
C2173 NAND2X1_LOC_498/Y INVX1_LOC_93/Y 0.08fF
C2174 INVX1_LOC_99/Y INVX1_LOC_59/A 0.00fF
C2175 INVX1_LOC_400/Y INVX1_LOC_31/Y 0.04fF
C2176 INVX1_LOC_312/Y INVX1_LOC_680/Y 0.01fF
C2177 NAND2X1_LOC_249/Y INVX1_LOC_301/Y 0.11fF
C2178 NAND2X1_LOC_180/B INVX1_LOC_350/A 0.04fF
C2179 NAND2X1_LOC_537/B INVX1_LOC_410/A 0.00fF
C2180 NAND2X1_LOC_790/B INVX1_LOC_153/Y 0.02fF
C2181 INVX1_LOC_536/A NAND2X1_LOC_685/a_36_24# 0.00fF
C2182 NAND2X1_LOC_318/A INVX1_LOC_479/Y 0.01fF
C2183 INVX1_LOC_367/A INVX1_LOC_99/Y 0.07fF
C2184 INVX1_LOC_256/Y INVX1_LOC_504/Y 0.03fF
C2185 INVX1_LOC_442/A NAND2X1_LOC_111/a_36_24# 0.00fF
C2186 INVX1_LOC_448/Y NAND2X1_LOC_274/B 0.01fF
C2187 NAND2X1_LOC_184/Y NAND2X1_LOC_843/a_36_24# -0.00fF
C2188 INVX1_LOC_442/A INVX1_LOC_89/Y 0.27fF
C2189 INVX1_LOC_566/A INVX1_LOC_48/Y 0.03fF
C2190 NAND2X1_LOC_513/a_36_24# INVX1_LOC_99/Y 0.00fF
C2191 INVX1_LOC_560/A INVX1_LOC_411/Y 0.01fF
C2192 INVX1_LOC_93/Y INVX1_LOC_142/A 0.00fF
C2193 INVX1_LOC_211/A INVX1_LOC_615/A 0.11fF
C2194 INVX1_LOC_604/A INVX1_LOC_44/Y 0.03fF
C2195 INVX1_LOC_560/Y NAND2X1_LOC_301/B 0.00fF
C2196 INVX1_LOC_510/Y NAND2X1_LOC_307/B 0.00fF
C2197 INVX1_LOC_442/A NAND2X1_LOC_319/a_36_24# 0.01fF
C2198 INVX1_LOC_366/Y INVX1_LOC_7/Y 0.01fF
C2199 INVX1_LOC_516/A INVX1_LOC_99/Y 0.02fF
C2200 INVX1_LOC_287/A INVX1_LOC_202/Y 1.54fF
C2201 INVX1_LOC_93/Y INVX1_LOC_377/Y 0.01fF
C2202 NAND2X1_LOC_249/Y INVX1_LOC_41/Y 0.06fF
C2203 INVX1_LOC_586/A INVX1_LOC_420/A 0.03fF
C2204 INVX1_LOC_526/A INVX1_LOC_261/Y 0.17fF
C2205 INVX1_LOC_547/Y NAND2X1_LOC_258/a_36_24# 0.00fF
C2206 INVX1_LOC_170/Y INVX1_LOC_586/A 0.09fF
C2207 INVX1_LOC_577/A INVX1_LOC_79/A 0.08fF
C2208 INVX1_LOC_449/A INVX1_LOC_50/Y 0.08fF
C2209 INVX1_LOC_400/A INVX1_LOC_99/Y 0.01fF
C2210 INVX1_LOC_363/Y INVX1_LOC_370/A 0.27fF
C2211 INVX1_LOC_392/A INVX1_LOC_99/Y 0.03fF
C2212 INVX1_LOC_438/A INVX1_LOC_280/A 0.07fF
C2213 INVX1_LOC_114/Y INVX1_LOC_675/A 0.03fF
C2214 INVX1_LOC_602/A INVX1_LOC_340/A 0.05fF
C2215 INVX1_LOC_183/Y INVX1_LOC_72/Y 0.02fF
C2216 INVX1_LOC_106/Y NAND2X1_LOC_108/Y 0.01fF
C2217 INVX1_LOC_679/Y INVX1_LOC_105/Y 0.00fF
C2218 INVX1_LOC_206/Y NAND2X1_LOC_615/a_36_24# 0.00fF
C2219 INVX1_LOC_431/A INVX1_LOC_145/Y 0.03fF
C2220 NAND2X1_LOC_184/Y NAND2X1_LOC_253/a_36_24# 0.01fF
C2221 NAND2X1_LOC_318/B INVX1_LOC_32/Y 0.02fF
C2222 INVX1_LOC_202/Y INVX1_LOC_479/Y 0.00fF
C2223 INVX1_LOC_270/A INVX1_LOC_63/Y 0.00fF
C2224 INPUT_1 INVX1_LOC_352/A 0.01fF
C2225 INVX1_LOC_662/A INVX1_LOC_132/Y 0.04fF
C2226 NAND2X1_LOC_331/A NAND2X1_LOC_609/B 0.45fF
C2227 INVX1_LOC_504/A INVX1_LOC_345/Y -0.05fF
C2228 INPUT_0 INVX1_LOC_274/Y 0.03fF
C2229 INVX1_LOC_315/Y INVX1_LOC_26/Y 0.03fF
C2230 INVX1_LOC_555/A INVX1_LOC_474/Y 0.04fF
C2231 INVX1_LOC_51/Y INVX1_LOC_373/Y 0.00fF
C2232 INVX1_LOC_84/A INVX1_LOC_480/A 0.07fF
C2233 INVX1_LOC_514/A INVX1_LOC_332/Y 0.08fF
C2234 INVX1_LOC_17/Y INVX1_LOC_103/Y 0.18fF
C2235 INVX1_LOC_93/Y INVX1_LOC_99/Y 3.16fF
C2236 INVX1_LOC_504/A INVX1_LOC_32/Y 0.07fF
C2237 INVX1_LOC_20/Y INVX1_LOC_662/A 0.10fF
C2238 INVX1_LOC_385/Y INVX1_LOC_6/Y 5.87fF
C2239 NAND2X1_LOC_615/B INVX1_LOC_194/Y 0.03fF
C2240 INVX1_LOC_554/A INVX1_LOC_92/A 0.75fF
C2241 INVX1_LOC_145/Y INVX1_LOC_18/Y 0.97fF
C2242 INVX1_LOC_17/Y INVX1_LOC_68/A 0.04fF
C2243 INVX1_LOC_202/Y INVX1_LOC_318/A 0.00fF
C2244 NAND2X1_LOC_111/a_36_24# INVX1_LOC_116/Y 0.00fF
C2245 INVX1_LOC_117/Y INVX1_LOC_159/Y 0.05fF
C2246 NAND2X1_LOC_775/B NAND2X1_LOC_444/A 0.05fF
C2247 INVX1_LOC_381/Y INVX1_LOC_385/A 0.01fF
C2248 INVX1_LOC_662/A NAND2X1_LOC_847/a_36_24# 0.01fF
C2249 NAND2X1_LOC_724/a_36_24# INVX1_LOC_92/A 0.01fF
C2250 INVX1_LOC_427/Y INVX1_LOC_387/Y 0.01fF
C2251 INVX1_LOC_47/Y INVX1_LOC_516/A 0.02fF
C2252 INVX1_LOC_89/Y INVX1_LOC_116/Y 0.13fF
C2253 INVX1_LOC_50/Y INVX1_LOC_186/Y 0.02fF
C2254 INVX1_LOC_188/Y INVX1_LOC_507/Y 0.13fF
C2255 INVX1_LOC_447/Y INVX1_LOC_69/Y 0.01fF
C2256 INVX1_LOC_469/Y INVX1_LOC_48/Y 0.03fF
C2257 INVX1_LOC_442/A NAND2X1_LOC_544/B 0.03fF
C2258 NAND2X1_LOC_448/B INVX1_LOC_259/Y 0.02fF
C2259 INVX1_LOC_105/Y INPUT_1 0.12fF
C2260 INVX1_LOC_328/A NAND2X1_LOC_404/a_36_24# 0.02fF
C2261 INVX1_LOC_35/Y INVX1_LOC_204/Y 0.05fF
C2262 NAND2X1_LOC_548/a_36_24# NAND2X1_LOC_531/Y 0.00fF
C2263 INVX1_LOC_406/Y INVX1_LOC_665/A 0.00fF
C2264 INVX1_LOC_675/A INVX1_LOC_99/Y 0.15fF
C2265 INVX1_LOC_549/Y INVX1_LOC_58/Y 0.01fF
C2266 INVX1_LOC_208/Y NAND2X1_LOC_503/Y 0.12fF
C2267 INVX1_LOC_183/A NAND2X1_LOC_397/Y 0.00fF
C2268 NAND2X1_LOC_174/B INVX1_LOC_261/Y 0.03fF
C2269 NAND2X1_LOC_148/A INVX1_LOC_655/A 0.05fF
C2270 NAND2X1_LOC_181/A INVX1_LOC_48/Y 0.07fF
C2271 INVX1_LOC_390/A INVX1_LOC_99/Y 0.01fF
C2272 INVX1_LOC_421/A INVX1_LOC_31/Y 0.07fF
C2273 NAND2X1_LOC_332/B INVX1_LOC_666/Y 0.51fF
C2274 INVX1_LOC_335/Y INVX1_LOC_26/Y 0.03fF
C2275 INVX1_LOC_632/A INVX1_LOC_79/A 0.07fF
C2276 INVX1_LOC_54/Y INVX1_LOC_69/Y 0.11fF
C2277 INVX1_LOC_21/Y INVX1_LOC_26/Y 8.10fF
C2278 INVX1_LOC_321/Y INVX1_LOC_245/A 0.01fF
C2279 INVX1_LOC_479/A INVX1_LOC_126/A 0.01fF
C2280 NAND2X1_LOC_591/Y INVX1_LOC_261/Y 0.01fF
C2281 INVX1_LOC_295/A INVX1_LOC_62/Y 0.01fF
C2282 INVX1_LOC_293/A INVX1_LOC_671/A 0.11fF
C2283 INVX1_LOC_509/Y INVX1_LOC_79/A 0.02fF
C2284 INVX1_LOC_93/Y INVX1_LOC_47/Y 0.15fF
C2285 INVX1_LOC_369/Y NAND2X1_LOC_296/Y 0.02fF
C2286 INVX1_LOC_253/Y INVX1_LOC_46/Y 0.00fF
C2287 INVX1_LOC_417/Y INVX1_LOC_79/A 0.13fF
C2288 INVX1_LOC_99/Y NAND2X1_LOC_9/a_36_24# 0.00fF
C2289 INVX1_LOC_369/A INVX1_LOC_41/Y 0.01fF
C2290 INVX1_LOC_516/A INVX1_LOC_119/Y 0.01fF
C2291 NAND2X1_LOC_749/a_36_24# INVX1_LOC_63/Y 0.00fF
C2292 INVX1_LOC_77/A INVX1_LOC_59/Y 0.01fF
C2293 INVX1_LOC_586/A INVX1_LOC_611/A 0.04fF
C2294 INVX1_LOC_204/Y INVX1_LOC_620/A 0.00fF
C2295 INVX1_LOC_79/A INVX1_LOC_59/Y 0.03fF
C2296 INVX1_LOC_58/Y INVX1_LOC_463/Y 0.23fF
C2297 INVX1_LOC_63/Y INVX1_LOC_46/Y 0.25fF
C2298 NAND2X1_LOC_196/a_36_24# INVX1_LOC_63/Y 0.00fF
C2299 INVX1_LOC_328/Y INVX1_LOC_50/Y 0.07fF
C2300 INVX1_LOC_89/Y INVX1_LOC_255/A 0.07fF
C2301 INVX1_LOC_556/Y NAND2X1_LOC_136/Y 0.01fF
C2302 INVX1_LOC_257/A INVX1_LOC_69/Y 0.08fF
C2303 INVX1_LOC_325/Y INVX1_LOC_443/A 0.50fF
C2304 NAND2X1_LOC_558/B INVX1_LOC_48/Y 0.00fF
C2305 INVX1_LOC_77/A INVX1_LOC_48/Y 0.02fF
C2306 INVX1_LOC_518/A INVX1_LOC_50/Y 0.04fF
C2307 INVX1_LOC_47/Y INVX1_LOC_675/A 0.09fF
C2308 INVX1_LOC_79/A INVX1_LOC_48/Y 0.20fF
C2309 NAND2X1_LOC_775/B NAND2X1_LOC_109/a_36_24# 0.00fF
C2310 INVX1_LOC_204/Y INVX1_LOC_621/Y 0.35fF
C2311 INVX1_LOC_267/Y INVX1_LOC_91/Y 0.01fF
C2312 INVX1_LOC_17/Y INVX1_LOC_635/Y 0.03fF
C2313 INVX1_LOC_116/Y NAND2X1_LOC_544/B 0.02fF
C2314 INVX1_LOC_95/A INVX1_LOC_49/Y 0.02fF
C2315 INVX1_LOC_93/Y INVX1_LOC_119/Y 3.47fF
C2316 INVX1_LOC_93/Y NAND2X1_LOC_66/Y 0.00fF
C2317 INVX1_LOC_376/Y INVX1_LOC_624/Y 0.02fF
C2318 INVX1_LOC_26/Y INVX1_LOC_181/Y 0.02fF
C2319 INVX1_LOC_7/Y NAND2X1_LOC_416/B 0.02fF
C2320 NAND2X1_LOC_274/B INVX1_LOC_58/Y 0.03fF
C2321 INVX1_LOC_507/Y INVX1_LOC_491/A 0.02fF
C2322 INVX1_LOC_559/Y INVX1_LOC_74/Y 0.91fF
C2323 INVX1_LOC_675/A INVX1_LOC_119/Y 0.06fF
C2324 INVX1_LOC_223/Y NAND2X1_LOC_845/B 0.03fF
C2325 INVX1_LOC_551/A INVX1_LOC_90/Y 0.01fF
C2326 INVX1_LOC_65/A NAND2X1_LOC_441/a_36_24# 0.00fF
C2327 NAND2X1_LOC_246/a_36_24# INVX1_LOC_669/A 0.01fF
C2328 INVX1_LOC_206/Y INVX1_LOC_638/A 0.08fF
C2329 INVX1_LOC_345/Y INVX1_LOC_346/Y 0.03fF
C2330 INPUT_6 INVX1_LOC_454/A 0.09fF
C2331 VDD NAND2X1_LOC_88/Y 0.01fF
C2332 INVX1_LOC_662/A INVX1_LOC_655/A 2.26fF
C2333 VDD INVX1_LOC_433/Y 0.26fF
C2334 INVX1_LOC_62/Y INVX1_LOC_139/Y 0.00fF
C2335 INPUT_0 NAND2X1_LOC_636/A 0.00fF
C2336 INVX1_LOC_183/Y NAND2X1_LOC_84/a_36_24# 0.01fF
C2337 INVX1_LOC_148/Y INVX1_LOC_58/Y 0.00fF
C2338 INVX1_LOC_79/A NAND2X1_LOC_434/B 0.01fF
C2339 INVX1_LOC_561/Y NAND2X1_LOC_591/B 0.02fF
C2340 INVX1_LOC_525/Y INVX1_LOC_91/Y 0.12fF
C2341 INVX1_LOC_49/Y INVX1_LOC_588/A 0.05fF
C2342 INVX1_LOC_531/Y NAND2X1_LOC_420/Y -0.02fF
C2343 INVX1_LOC_41/Y NAND2X1_LOC_605/B 0.01fF
C2344 INVX1_LOC_63/Y INVX1_LOC_75/A 0.01fF
C2345 VDD NAND2X1_LOC_592/B 0.01fF
C2346 INVX1_LOC_438/Y NAND2X1_LOC_555/a_36_24# 0.01fF
C2347 INVX1_LOC_206/Y NAND2X1_LOC_701/a_36_24# 0.01fF
C2348 INVX1_LOC_199/Y INVX1_LOC_270/Y 0.05fF
C2349 INPUT_0 INVX1_LOC_549/A 0.04fF
C2350 INVX1_LOC_679/Y INVX1_LOC_109/Y 0.00fF
C2351 INVX1_LOC_242/Y INVX1_LOC_666/Y 0.03fF
C2352 INVX1_LOC_75/Y INVX1_LOC_90/Y 0.02fF
C2353 INVX1_LOC_37/Y INVX1_LOC_36/A 0.00fF
C2354 INVX1_LOC_199/Y INVX1_LOC_92/A 0.10fF
C2355 NAND2X1_LOC_45/Y INVX1_LOC_362/Y 0.07fF
C2356 INVX1_LOC_686/A INVX1_LOC_638/A 1.25fF
C2357 NAND2X1_LOC_498/Y INVX1_LOC_395/A 0.10fF
C2358 INVX1_LOC_395/A INVX1_LOC_570/A 0.07fF
C2359 NAND2X1_LOC_299/a_36_24# INVX1_LOC_634/Y 0.01fF
C2360 NAND2X1_LOC_843/B NAND2X1_LOC_248/B 0.00fF
C2361 INVX1_LOC_193/Y INVX1_LOC_586/A 0.04fF
C2362 NAND2X1_LOC_241/B INVX1_LOC_273/A 0.03fF
C2363 INVX1_LOC_681/Y INVX1_LOC_109/Y 0.02fF
C2364 INVX1_LOC_206/Y INVX1_LOC_398/A 0.01fF
C2365 INPUT_1 INVX1_LOC_109/Y 0.03fF
C2366 VDD INVX1_LOC_232/Y 0.21fF
C2367 VDD NAND2X1_LOC_616/Y 0.03fF
C2368 INVX1_LOC_20/Y INVX1_LOC_320/Y 0.01fF
C2369 INVX1_LOC_266/A INVX1_LOC_400/Y 0.03fF
C2370 INVX1_LOC_392/Y INVX1_LOC_502/Y 0.00fF
C2371 INVX1_LOC_65/Y INVX1_LOC_76/Y 0.09fF
C2372 NAND2X1_LOC_173/Y NAND2X1_LOC_122/Y 0.03fF
C2373 INVX1_LOC_410/Y INVX1_LOC_80/A 0.06fF
C2374 NAND2X1_LOC_525/Y INVX1_LOC_293/Y 0.16fF
C2375 INVX1_LOC_80/A INVX1_LOC_375/A 0.24fF
C2376 VDD INVX1_LOC_108/Y 0.21fF
C2377 INVX1_LOC_206/Y NAND2X1_LOC_697/Y 0.07fF
C2378 NAND2X1_LOC_45/Y INVX1_LOC_548/A 0.02fF
C2379 INVX1_LOC_393/Y NAND2X1_LOC_179/Y 0.00fF
C2380 INPUT_0 INVX1_LOC_230/A 0.07fF
C2381 NAND2X1_LOC_457/A INVX1_LOC_35/Y 0.07fF
C2382 INVX1_LOC_590/Y NAND2X1_LOC_237/Y 0.01fF
C2383 INVX1_LOC_395/A INVX1_LOC_99/Y 0.15fF
C2384 INVX1_LOC_271/A INVX1_LOC_154/Y -0.00fF
C2385 VDD INVX1_LOC_497/Y 0.27fF
C2386 INVX1_LOC_320/Y INVX1_LOC_300/A 0.01fF
C2387 INVX1_LOC_11/Y INVX1_LOC_553/Y 0.01fF
C2388 NAND2X1_LOC_242/A INVX1_LOC_396/A 0.01fF
C2389 INVX1_LOC_32/Y NAND2X1_LOC_76/B 0.07fF
C2390 VDD INVX1_LOC_230/Y 0.34fF
C2391 INVX1_LOC_577/A INVX1_LOC_48/Y 0.01fF
C2392 INVX1_LOC_425/A INVX1_LOC_12/Y 0.49fF
C2393 INVX1_LOC_20/Y NAND2X1_LOC_147/a_36_24# 0.01fF
C2394 INVX1_LOC_362/Y INVX1_LOC_99/Y 0.03fF
C2395 INVX1_LOC_287/A INVX1_LOC_76/Y 0.03fF
C2396 NAND2X1_LOC_334/A INVX1_LOC_638/A 0.07fF
C2397 INVX1_LOC_78/A INVX1_LOC_51/Y 0.05fF
C2398 INVX1_LOC_11/Y INVX1_LOC_546/A 0.00fF
C2399 INVX1_LOC_677/Y INVX1_LOC_677/A 0.19fF
C2400 NAND2X1_LOC_45/Y INVX1_LOC_31/Y 0.36fF
C2401 INVX1_LOC_432/Y INVX1_LOC_321/A 0.01fF
C2402 INVX1_LOC_206/Y NAND2X1_LOC_203/a_36_24# 0.00fF
C2403 INVX1_LOC_586/A NAND2X1_LOC_461/a_36_24# 0.00fF
C2404 INVX1_LOC_521/Y INVX1_LOC_50/Y 0.01fF
C2405 INVX1_LOC_379/A INVX1_LOC_378/A 0.09fF
C2406 INVX1_LOC_424/A INVX1_LOC_63/Y 0.03fF
C2407 INVX1_LOC_35/Y INVX1_LOC_482/A 0.04fF
C2408 INVX1_LOC_118/Y INVX1_LOC_66/A 0.03fF
C2409 INVX1_LOC_304/Y NAND2X1_LOC_613/Y -0.00fF
C2410 INVX1_LOC_395/A INVX1_LOC_568/A 0.01fF
C2411 NAND2X1_LOC_498/Y INVX1_LOC_31/Y 0.10fF
C2412 INVX1_LOC_570/A INVX1_LOC_31/Y 0.44fF
C2413 INVX1_LOC_54/Y INVX1_LOC_586/A 1.63fF
C2414 INVX1_LOC_405/A NAND2X1_LOC_642/a_36_24# 0.00fF
C2415 INVX1_LOC_53/Y INVX1_LOC_567/Y 0.03fF
C2416 INVX1_LOC_395/A INVX1_LOC_47/Y 0.21fF
C2417 INVX1_LOC_21/Y INVX1_LOC_369/A 0.25fF
C2418 NAND2X1_LOC_69/B INVX1_LOC_100/Y 0.37fF
C2419 INVX1_LOC_547/Y NAND2X1_LOC_253/Y 0.12fF
C2420 VDD INVX1_LOC_35/A 0.00fF
C2421 INVX1_LOC_395/A NAND2X1_LOC_557/B 0.03fF
C2422 NAND2X1_LOC_475/A INVX1_LOC_390/A 0.02fF
C2423 INVX1_LOC_438/A INVX1_LOC_328/Y 0.07fF
C2424 INVX1_LOC_421/A INVX1_LOC_51/Y 0.01fF
C2425 INVX1_LOC_301/A NAND2X1_LOC_545/A 0.02fF
C2426 INVX1_LOC_468/Y INVX1_LOC_134/Y 0.05fF
C2427 INVX1_LOC_548/Y INVX1_LOC_63/Y 0.02fF
C2428 INVX1_LOC_578/A INVX1_LOC_65/A 0.03fF
C2429 NAND2X1_LOC_88/Y NAND2X1_LOC_786/B 0.03fF
C2430 INVX1_LOC_602/A INVX1_LOC_455/A 0.03fF
C2431 INVX1_LOC_530/A INVX1_LOC_7/Y 0.00fF
C2432 NAND2X1_LOC_790/B INVX1_LOC_41/Y 0.15fF
C2433 INVX1_LOC_362/Y INVX1_LOC_47/Y 0.39fF
C2434 INVX1_LOC_257/A INVX1_LOC_586/A 0.10fF
C2435 INVX1_LOC_237/Y INVX1_LOC_58/Y 0.01fF
C2436 INVX1_LOC_80/A INVX1_LOC_662/Y 0.03fF
C2437 INVX1_LOC_335/A NAND2X1_LOC_681/a_36_24# -0.00fF
C2438 INVX1_LOC_126/Y INPUT_1 0.09fF
C2439 INVX1_LOC_53/Y NAND2X1_LOC_696/a_36_24# 0.00fF
C2440 INVX1_LOC_80/A INVX1_LOC_61/A 0.01fF
C2441 NAND2X1_LOC_184/Y NAND2X1_LOC_523/B 0.00fF
C2442 INVX1_LOC_4/Y INVX1_LOC_3/A 0.00fF
C2443 NAND2X1_LOC_152/Y INVX1_LOC_6/Y 0.14fF
C2444 INVX1_LOC_89/Y INVX1_LOC_146/A 0.01fF
C2445 INVX1_LOC_427/Y INVX1_LOC_386/Y 0.16fF
C2446 INVX1_LOC_530/Y INVX1_LOC_63/Y 0.04fF
C2447 INVX1_LOC_376/A INVX1_LOC_45/Y 0.08fF
C2448 NAND2X1_LOC_527/Y INVX1_LOC_134/Y 0.02fF
C2449 INVX1_LOC_342/Y INVX1_LOC_602/Y 0.44fF
C2450 INVX1_LOC_561/Y INVX1_LOC_79/A 0.03fF
C2451 INVX1_LOC_298/A INVX1_LOC_635/A 0.33fF
C2452 INVX1_LOC_301/A INVX1_LOC_666/Y 0.07fF
C2453 INVX1_LOC_548/A INVX1_LOC_99/Y 0.07fF
C2454 INVX1_LOC_395/A INVX1_LOC_119/Y 0.01fF
C2455 NAND2X1_LOC_714/a_36_24# INVX1_LOC_376/Y 0.00fF
C2456 NAND2X1_LOC_498/Y INVX1_LOC_128/A 0.01fF
C2457 INVX1_LOC_17/Y INVX1_LOC_360/Y 0.12fF
C2458 INVX1_LOC_578/A NAND2X1_LOC_604/a_36_24# 0.00fF
C2459 NAND2X1_LOC_97/B NAND2X1_LOC_333/B 0.01fF
C2460 INVX1_LOC_255/Y INVX1_LOC_26/Y 0.03fF
C2461 INVX1_LOC_395/A NAND2X1_LOC_66/Y 0.06fF
C2462 INVX1_LOC_21/Y INVX1_LOC_603/A 0.03fF
C2463 NAND2X1_LOC_318/A INVX1_LOC_63/Y 0.04fF
C2464 INVX1_LOC_451/A INVX1_LOC_452/A 0.04fF
C2465 INVX1_LOC_47/Y INVX1_LOC_683/Y 0.15fF
C2466 VDD INVX1_LOC_598/Y 0.40fF
C2467 INVX1_LOC_145/Y GATE_222 0.01fF
C2468 NAND2X1_LOC_106/Y INVX1_LOC_53/Y 0.08fF
C2469 INVX1_LOC_285/A INVX1_LOC_292/Y 0.23fF
C2470 INVX1_LOC_373/A INVX1_LOC_41/Y 0.76fF
C2471 INVX1_LOC_619/A INVX1_LOC_601/Y 0.15fF
C2472 INVX1_LOC_604/Y NAND2X1_LOC_503/Y 0.11fF
C2473 INVX1_LOC_321/A NAND2X1_LOC_494/a_36_24# 0.00fF
C2474 INVX1_LOC_504/A NAND2X1_LOC_652/a_36_24# 0.01fF
C2475 NAND2X1_LOC_836/B INVX1_LOC_333/A 0.02fF
C2476 INVX1_LOC_90/A INVX1_LOC_6/Y 0.01fF
C2477 INVX1_LOC_59/Y INVX1_LOC_48/Y 0.09fF
C2478 INVX1_LOC_376/A INVX1_LOC_348/A 0.04fF
C2479 INVX1_LOC_54/Y NAND2X1_LOC_378/Y 0.01fF
C2480 INVX1_LOC_45/Y INVX1_LOC_502/A 0.19fF
C2481 INVX1_LOC_577/Y INVX1_LOC_26/Y 0.04fF
C2482 INVX1_LOC_625/A INVX1_LOC_32/Y 0.02fF
C2483 INVX1_LOC_385/Y NAND2X1_LOC_294/Y 0.03fF
C2484 INVX1_LOC_25/Y INVX1_LOC_93/Y 0.01fF
C2485 INVX1_LOC_31/Y INVX1_LOC_99/Y 2.54fF
C2486 INVX1_LOC_163/Y INVX1_LOC_491/A 0.02fF
C2487 INVX1_LOC_680/Y INVX1_LOC_6/Y 0.01fF
C2488 INVX1_LOC_361/Y INVX1_LOC_510/A 0.15fF
C2489 INVX1_LOC_100/A INVX1_LOC_145/Y 0.18fF
C2490 INVX1_LOC_166/A NAND2X1_LOC_307/a_36_24# 0.00fF
C2491 INVX1_LOC_412/Y INVX1_LOC_625/Y 0.03fF
C2492 INVX1_LOC_379/A NAND2X1_LOC_632/a_36_24# 0.00fF
C2493 INVX1_LOC_353/Y INVX1_LOC_242/Y 0.02fF
C2494 NAND2X1_LOC_418/Y INVX1_LOC_66/A 0.13fF
C2495 INVX1_LOC_654/A NAND2X1_LOC_833/B 0.08fF
C2496 INVX1_LOC_377/Y INVX1_LOC_128/A 0.01fF
C2497 INVX1_LOC_442/A INVX1_LOC_347/A 0.58fF
C2498 INVX1_LOC_172/A INVX1_LOC_50/Y 0.34fF
C2499 INVX1_LOC_198/A NAND2X1_LOC_243/A 0.17fF
C2500 INVX1_LOC_176/A INVX1_LOC_6/Y 0.29fF
C2501 NAND2X1_LOC_267/A INVX1_LOC_603/A 0.02fF
C2502 INVX1_LOC_542/A INVX1_LOC_495/Y 0.00fF
C2503 NAND2X1_LOC_498/B INVX1_LOC_588/A 0.18fF
C2504 INVX1_LOC_256/Y INVX1_LOC_114/A 0.01fF
C2505 INVX1_LOC_340/Y INVX1_LOC_74/Y 5.87fF
C2506 INVX1_LOC_280/Y INVX1_LOC_281/A 0.09fF
C2507 NAND2X1_LOC_122/Y INVX1_LOC_354/A 0.01fF
C2508 INVX1_LOC_98/A NAND2X1_LOC_94/a_36_24# 0.00fF
C2509 NAND2X1_LOC_147/a_36_24# INVX1_LOC_655/A 0.00fF
C2510 INVX1_LOC_492/A INVX1_LOC_476/A 0.01fF
C2511 INVX1_LOC_298/Y INVX1_LOC_674/Y 0.27fF
C2512 INVX1_LOC_235/Y INVX1_LOC_41/Y 0.01fF
C2513 INVX1_LOC_168/A INVX1_LOC_62/Y 0.01fF
C2514 INVX1_LOC_76/Y INVX1_LOC_588/A 0.27fF
C2515 INVX1_LOC_202/Y INVX1_LOC_63/Y 0.07fF
C2516 INVX1_LOC_525/Y NAND2X1_LOC_333/B 0.09fF
C2517 INVX1_LOC_123/A INVX1_LOC_31/Y 0.01fF
C2518 NAND2X1_LOC_309/a_36_24# NAND2X1_LOC_267/A 0.00fF
C2519 INVX1_LOC_277/A INVX1_LOC_69/Y 0.00fF
C2520 INVX1_LOC_491/A NAND2X1_LOC_646/a_36_24# 0.00fF
C2521 INVX1_LOC_649/Y INVX1_LOC_667/A 0.01fF
C2522 INVX1_LOC_199/Y INPUT_1 0.03fF
C2523 INVX1_LOC_493/A INVX1_LOC_496/A 0.02fF
C2524 INVX1_LOC_20/Y INVX1_LOC_666/Y 0.42fF
C2525 NAND2X1_LOC_491/Y INVX1_LOC_48/Y 0.01fF
C2526 INVX1_LOC_167/A INVX1_LOC_496/A 0.02fF
C2527 INVX1_LOC_31/Y INVX1_LOC_47/Y 3.66fF
C2528 INVX1_LOC_21/Y NAND2X1_LOC_626/Y 0.03fF
C2529 INVX1_LOC_523/Y INVX1_LOC_66/A 0.02fF
C2530 INVX1_LOC_26/Y INVX1_LOC_481/Y 0.01fF
C2531 INVX1_LOC_31/Y NAND2X1_LOC_557/B 0.04fF
C2532 NAND2X1_LOC_410/a_36_24# NAND2X1_LOC_410/Y 0.02fF
C2533 INVX1_LOC_32/Y NAND2X1_LOC_52/Y 0.01fF
C2534 INVX1_LOC_679/A INVX1_LOC_655/A 0.03fF
C2535 INVX1_LOC_89/Y INVX1_LOC_69/Y 5.59fF
C2536 INVX1_LOC_35/Y INVX1_LOC_422/A 0.06fF
C2537 INVX1_LOC_387/Y INVX1_LOC_63/Y 0.03fF
C2538 INVX1_LOC_99/Y INVX1_LOC_473/Y 0.01fF
C2539 INVX1_LOC_93/Y INVX1_LOC_15/Y 0.22fF
C2540 INVX1_LOC_6/Y INVX1_LOC_420/A 0.23fF
C2541 INVX1_LOC_58/Y INVX1_LOC_340/A 0.01fF
C2542 INVX1_LOC_253/Y INVX1_LOC_49/Y 0.00fF
C2543 INVX1_LOC_170/Y INVX1_LOC_6/Y 0.05fF
C2544 INVX1_LOC_50/Y INVX1_LOC_224/A 0.04fF
C2545 INVX1_LOC_662/Y INVX1_LOC_102/Y 0.08fF
C2546 INVX1_LOC_74/Y INVX1_LOC_155/Y 0.00fF
C2547 NAND2X1_LOC_722/a_36_24# INVX1_LOC_636/A 0.00fF
C2548 NAND2X1_LOC_237/Y INVX1_LOC_211/A 0.03fF
C2549 INVX1_LOC_58/Y INVX1_LOC_212/Y 0.03fF
C2550 INVX1_LOC_116/Y INVX1_LOC_347/A 0.01fF
C2551 INVX1_LOC_300/A INVX1_LOC_666/Y 0.03fF
C2552 INVX1_LOC_49/Y INVX1_LOC_63/Y 0.11fF
C2553 INVX1_LOC_47/Y INVX1_LOC_682/Y 0.17fF
C2554 INVX1_LOC_75/Y INVX1_LOC_98/Y 0.09fF
C2555 INVX1_LOC_31/Y INVX1_LOC_119/Y 0.24fF
C2556 INVX1_LOC_399/A INVX1_LOC_199/Y 0.01fF
C2557 INVX1_LOC_31/Y NAND2X1_LOC_66/Y 0.04fF
C2558 INVX1_LOC_47/Y INVX1_LOC_128/A 0.04fF
C2559 INVX1_LOC_63/Y INVX1_LOC_642/Y 0.01fF
C2560 INVX1_LOC_53/Y INVX1_LOC_92/A 5.93fF
C2561 INVX1_LOC_179/A INVX1_LOC_44/Y 0.07fF
C2562 INVX1_LOC_46/Y INVX1_LOC_669/A 0.01fF
C2563 INVX1_LOC_117/Y NAND2X1_LOC_372/Y 0.18fF
C2564 INVX1_LOC_502/A NAND2X1_LOC_276/A 0.03fF
C2565 NAND2X1_LOC_503/B VDD 0.02fF
C2566 INVX1_LOC_222/Y VDD 0.26fF
C2567 NAND2X1_LOC_290/a_36_24# INVX1_LOC_26/Y 0.01fF
C2568 INVX1_LOC_278/A INVX1_LOC_220/A 0.07fF
C2569 INVX1_LOC_255/A INVX1_LOC_347/A 0.03fF
C2570 INVX1_LOC_584/A INVX1_LOC_463/A 0.02fF
C2571 INVX1_LOC_69/Y NAND2X1_LOC_544/B 0.03fF
C2572 INVX1_LOC_119/Y INVX1_LOC_128/A 0.00fF
C2573 INVX1_LOC_63/Y INVX1_LOC_92/Y 0.01fF
C2574 VDD INVX1_LOC_127/A -0.00fF
C2575 INVX1_LOC_329/Y NAND2X1_LOC_406/B 0.00fF
C2576 INVX1_LOC_434/A INVX1_LOC_278/A 0.03fF
C2577 INVX1_LOC_664/A NAND2X1_LOC_843/B 0.03fF
C2578 NAND2X1_LOC_799/a_36_24# INVX1_LOC_288/A 0.00fF
C2579 INVX1_LOC_45/Y INVX1_LOC_388/Y 0.00fF
C2580 NAND2X1_LOC_475/A INVX1_LOC_395/A 0.07fF
C2581 VDD INVX1_LOC_249/Y 0.21fF
C2582 INVX1_LOC_366/A NAND2X1_LOC_205/a_36_24# 0.01fF
C2583 NAND2X1_LOC_45/Y INVX1_LOC_51/Y 0.04fF
C2584 VDD INVX1_LOC_325/Y 0.33fF
C2585 INVX1_LOC_505/Y INVX1_LOC_479/A 0.01fF
C2586 INVX1_LOC_90/Y NAND2X1_LOC_98/B 0.01fF
C2587 INVX1_LOC_21/Y NAND2X1_LOC_790/B 0.05fF
C2588 NAND2X1_LOC_498/Y INVX1_LOC_51/Y 1.05fF
C2589 INVX1_LOC_50/Y INVX1_LOC_109/Y 0.03fF
C2590 NAND2X1_LOC_451/B NAND2X1_LOC_428/Y 0.00fF
C2591 INVX1_LOC_552/Y NAND2X1_LOC_318/A 0.00fF
C2592 INVX1_LOC_570/A INVX1_LOC_51/Y 0.07fF
C2593 INVX1_LOC_150/Y INVX1_LOC_586/A 0.52fF
C2594 NAND2X1_LOC_704/B INVX1_LOC_546/A 0.03fF
C2595 NAND2X1_LOC_13/Y INVX1_LOC_400/Y 0.03fF
C2596 INVX1_LOC_453/Y INVX1_LOC_220/A 0.03fF
C2597 INVX1_LOC_463/A INVX1_LOC_537/A 0.53fF
C2598 INVX1_LOC_206/Y INVX1_LOC_134/Y 0.23fF
C2599 VDD NAND2X1_LOC_393/Y 0.00fF
C2600 INVX1_LOC_602/A INVX1_LOC_26/A 0.04fF
C2601 NAND2X1_LOC_48/Y INVX1_LOC_206/Y 0.01fF
C2602 INVX1_LOC_397/A INVX1_LOC_398/A 0.31fF
C2603 INVX1_LOC_95/Y INVX1_LOC_50/Y 0.01fF
C2604 VDD INVX1_LOC_248/Y 0.01fF
C2605 INVX1_LOC_561/Y INVX1_LOC_632/A -0.05fF
C2606 INPUT_0 NAND2X1_LOC_325/B 0.46fF
C2607 INVX1_LOC_395/A INVX1_LOC_136/Y 0.15fF
C2608 INVX1_LOC_554/A INVX1_LOC_50/Y 0.02fF
C2609 GATE_741 NAND2X1_LOC_467/A 0.02fF
C2610 INVX1_LOC_373/A INVX1_LOC_358/Y 0.01fF
C2611 INVX1_LOC_405/A INVX1_LOC_46/Y 0.03fF
C2612 INVX1_LOC_206/Y INVX1_LOC_316/Y 0.01fF
C2613 INVX1_LOC_21/Y INVX1_LOC_103/A 0.07fF
C2614 INVX1_LOC_434/A INVX1_LOC_453/Y 4.65fF
C2615 INVX1_LOC_44/A INVX1_LOC_190/Y 0.01fF
C2616 INVX1_LOC_308/Y INVX1_LOC_145/Y 0.01fF
C2617 INVX1_LOC_259/A INVX1_LOC_188/Y 0.16fF
C2618 NAND2X1_LOC_543/B INVX1_LOC_93/Y 0.37fF
C2619 INVX1_LOC_542/A INVX1_LOC_536/A 0.00fF
C2620 INPUT_3 INVX1_LOC_175/A 0.06fF
C2621 INVX1_LOC_607/Y INVX1_LOC_107/A 0.02fF
C2622 NAND2X1_LOC_592/a_36_24# INVX1_LOC_47/Y 0.01fF
C2623 INVX1_LOC_426/A INVX1_LOC_47/Y 0.07fF
C2624 INVX1_LOC_579/A NAND2X1_LOC_173/Y 0.03fF
C2625 NAND2X1_LOC_505/Y INVX1_LOC_99/Y 0.23fF
C2626 NAND2X1_LOC_764/Y INVX1_LOC_623/Y 0.01fF
C2627 INVX1_LOC_608/Y INVX1_LOC_45/Y 0.01fF
C2628 INVX1_LOC_34/Y INVX1_LOC_1/Y 0.28fF
C2629 INVX1_LOC_65/Y INVX1_LOC_228/A 0.01fF
C2630 INVX1_LOC_214/Y INVX1_LOC_547/Y 0.02fF
C2631 INVX1_LOC_206/Y NAND2X1_LOC_165/Y 0.01fF
C2632 INVX1_LOC_244/Y INVX1_LOC_423/Y 1.46fF
C2633 INVX1_LOC_515/Y INVX1_LOC_515/A 0.01fF
C2634 INVX1_LOC_17/Y INVX1_LOC_45/Y 0.27fF
C2635 NAND2X1_LOC_475/A INVX1_LOC_31/Y 0.22fF
C2636 INVX1_LOC_51/Y INVX1_LOC_99/Y 0.10fF
C2637 NAND2X1_LOC_187/Y INVX1_LOC_140/Y 0.02fF
C2638 NAND2X1_LOC_183/a_36_24# NAND2X1_LOC_181/A 0.00fF
C2639 INVX1_LOC_686/A INVX1_LOC_134/Y 0.02fF
C2640 NAND2X1_LOC_164/Y INVX1_LOC_32/Y 0.07fF
C2641 NAND2X1_LOC_638/A INVX1_LOC_59/A 0.12fF
C2642 NAND2X1_LOC_673/a_36_24# INVX1_LOC_169/A 0.00fF
C2643 INVX1_LOC_489/A NAND2X1_LOC_631/a_36_24# 0.00fF
C2644 INVX1_LOC_21/Y INVX1_LOC_235/Y 0.07fF
C2645 INVX1_LOC_435/Y NAND2X1_LOC_184/Y 0.11fF
C2646 INVX1_LOC_375/A INVX1_LOC_374/Y 0.00fF
C2647 INVX1_LOC_409/A INVX1_LOC_58/Y 0.03fF
C2648 INVX1_LOC_384/Y INVX1_LOC_278/Y 0.01fF
C2649 INVX1_LOC_53/Y INVX1_LOC_679/Y 0.09fF
C2650 INVX1_LOC_406/Y INVX1_LOC_367/Y 0.01fF
C2651 INVX1_LOC_412/Y INVX1_LOC_258/Y 0.00fF
C2652 INVX1_LOC_184/A INVX1_LOC_7/Y 0.22fF
C2653 NAND2X1_LOC_180/B NAND2X1_LOC_775/B 0.02fF
C2654 INPUT_3 INVX1_LOC_17/Y 0.01fF
C2655 INVX1_LOC_76/Y NAND2X1_LOC_646/A 0.00fF
C2656 INVX1_LOC_65/Y INVX1_LOC_32/Y 0.08fF
C2657 INVX1_LOC_395/A INVX1_LOC_96/A 0.00fF
C2658 NAND2X1_LOC_331/A INVX1_LOC_139/Y 0.01fF
C2659 NAND2X1_LOC_393/a_36_24# INVX1_LOC_328/Y 0.00fF
C2660 NAND2X1_LOC_403/A INVX1_LOC_324/A 0.09fF
C2661 INVX1_LOC_145/Y INVX1_LOC_635/A 0.01fF
C2662 INVX1_LOC_601/A INVX1_LOC_207/Y 0.16fF
C2663 INVX1_LOC_396/Y NAND2X1_LOC_165/Y 0.04fF
C2664 INVX1_LOC_566/Y INVX1_LOC_674/A 0.02fF
C2665 INVX1_LOC_438/A INVX1_LOC_224/A 0.02fF
C2666 INVX1_LOC_617/Y INVX1_LOC_361/Y 0.07fF
C2667 INVX1_LOC_89/Y INVX1_LOC_586/A 0.31fF
C2668 NAND2X1_LOC_13/a_36_24# NAND2X1_LOC_267/A 0.03fF
C2669 NAND2X1_LOC_737/a_36_24# INVX1_LOC_145/Y 0.01fF
C2670 INVX1_LOC_51/Y INVX1_LOC_47/Y 0.95fF
C2671 INVX1_LOC_154/A INVX1_LOC_586/A 0.03fF
C2672 NAND2X1_LOC_179/Y INVX1_LOC_442/Y 0.03fF
C2673 NAND2X1_LOC_163/B INVX1_LOC_58/Y 0.01fF
C2674 INVX1_LOC_84/A INVX1_LOC_46/Y 7.85fF
C2675 INVX1_LOC_448/Y NAND2X1_LOC_372/Y 0.01fF
C2676 INVX1_LOC_21/Y INVX1_LOC_81/Y 0.02fF
C2677 INVX1_LOC_619/A INVX1_LOC_198/A 1.23fF
C2678 INVX1_LOC_98/A INVX1_LOC_63/Y 0.14fF
C2679 INVX1_LOC_53/Y INPUT_1 0.80fF
C2680 INVX1_LOC_625/A NAND2X1_LOC_226/Y 0.32fF
C2681 INVX1_LOC_449/A INVX1_LOC_117/Y 0.07fF
C2682 INVX1_LOC_126/A INVX1_LOC_66/A 0.00fF
C2683 INVX1_LOC_255/Y NAND2X1_LOC_605/B 0.00fF
C2684 NAND2X1_LOC_339/a_36_24# INVX1_LOC_63/Y 0.00fF
C2685 INVX1_LOC_20/Y INVX1_LOC_94/Y 0.16fF
C2686 GATE_579 NAND2X1_LOC_480/a_36_24# 0.00fF
C2687 INVX1_LOC_586/A INVX1_LOC_501/A 0.00fF
C2688 INVX1_LOC_173/A NAND2X1_LOC_845/B 0.04fF
C2689 INVX1_LOC_76/Y INVX1_LOC_63/Y 0.07fF
C2690 INVX1_LOC_490/Y NAND2X1_LOC_269/B 0.02fF
C2691 INVX1_LOC_287/A INVX1_LOC_32/Y 0.00fF
C2692 INVX1_LOC_395/A INVX1_LOC_475/Y 0.06fF
C2693 INVX1_LOC_686/A INVX1_LOC_65/A 0.02fF
C2694 INVX1_LOC_53/Y INVX1_LOC_292/Y 0.58fF
C2695 INVX1_LOC_254/A INVX1_LOC_99/Y 0.01fF
C2696 NAND2X1_LOC_775/B NAND2X1_LOC_444/a_36_24# 0.00fF
C2697 INVX1_LOC_51/Y INVX1_LOC_119/Y 1.01fF
C2698 INVX1_LOC_547/A NAND2X1_LOC_258/a_36_24# 0.00fF
C2699 INVX1_LOC_273/A NAND2X1_LOC_786/B 0.19fF
C2700 NAND2X1_LOC_457/A INVX1_LOC_364/A 0.03fF
C2701 INVX1_LOC_587/Y INVX1_LOC_35/Y 0.03fF
C2702 INVX1_LOC_51/Y NAND2X1_LOC_66/Y 0.42fF
C2703 INVX1_LOC_316/Y INVX1_LOC_342/A 0.22fF
C2704 INVX1_LOC_129/A INVX1_LOC_46/Y 0.01fF
C2705 INVX1_LOC_607/Y NAND2X1_LOC_285/A 0.04fF
C2706 INVX1_LOC_139/A INVX1_LOC_588/A 0.01fF
C2707 INVX1_LOC_435/Y INVX1_LOC_75/Y 0.43fF
C2708 NAND2X1_LOC_43/Y INVX1_LOC_31/Y 0.07fF
C2709 INVX1_LOC_524/Y INVX1_LOC_353/A 0.05fF
C2710 INVX1_LOC_575/A INVX1_LOC_477/Y 0.01fF
C2711 NAND2X1_LOC_137/A INVX1_LOC_556/Y 0.01fF
C2712 NAND2X1_LOC_461/a_36_24# INVX1_LOC_6/Y 0.00fF
C2713 INVX1_LOC_66/A INVX1_LOC_252/Y 0.03fF
C2714 INVX1_LOC_443/A INVX1_LOC_445/A 0.03fF
C2715 INVX1_LOC_117/Y INVX1_LOC_186/Y 0.03fF
C2716 INVX1_LOC_435/A NAND2X1_LOC_613/a_36_24# 0.01fF
C2717 INVX1_LOC_293/Y INVX1_LOC_502/A 0.07fF
C2718 INVX1_LOC_213/Y NAND2X1_LOC_106/Y 0.11fF
C2719 INVX1_LOC_640/Y INVX1_LOC_641/Y 0.02fF
C2720 NAND2X1_LOC_416/Y INVX1_LOC_379/Y 0.01fF
C2721 INVX1_LOC_586/A NAND2X1_LOC_544/B 0.03fF
C2722 INVX1_LOC_369/A INVX1_LOC_26/Y 0.58fF
C2723 INVX1_LOC_318/A INVX1_LOC_32/Y 0.00fF
C2724 INVX1_LOC_54/Y INVX1_LOC_6/Y 1.99fF
C2725 NAND2X1_LOC_530/a_36_24# NAND2X1_LOC_66/Y 0.00fF
C2726 INVX1_LOC_455/A INVX1_LOC_58/Y 0.00fF
C2727 INVX1_LOC_58/Y INVX1_LOC_352/Y 0.03fF
C2728 INVX1_LOC_666/A INVX1_LOC_211/A 0.05fF
C2729 INVX1_LOC_556/Y INVX1_LOC_107/Y 0.02fF
C2730 INVX1_LOC_435/Y NAND2X1_LOC_271/A 0.10fF
C2731 INVX1_LOC_199/Y INVX1_LOC_50/Y 0.03fF
C2732 NAND2X1_LOC_545/a_36_24# INPUT_1 0.00fF
C2733 INVX1_LOC_47/Y INVX1_LOC_254/A 0.01fF
C2734 INVX1_LOC_397/Y INVX1_LOC_32/Y 0.23fF
C2735 INVX1_LOC_35/Y INVX1_LOC_9/Y 1.36fF
C2736 INVX1_LOC_79/A INVX1_LOC_155/Y 0.03fF
C2737 NAND2X1_LOC_615/Y INVX1_LOC_48/Y 0.05fF
C2738 INVX1_LOC_596/A INVX1_LOC_75/Y 0.02fF
C2739 INVX1_LOC_366/A INVX1_LOC_619/Y 0.01fF
C2740 INVX1_LOC_80/A NAND2X1_LOC_528/Y 0.09fF
C2741 INVX1_LOC_26/Y NAND2X1_LOC_275/Y 0.12fF
C2742 INVX1_LOC_378/A INVX1_LOC_488/Y 0.02fF
C2743 NAND2X1_LOC_503/Y INVX1_LOC_63/Y 0.05fF
C2744 INVX1_LOC_565/A INVX1_LOC_41/Y 0.13fF
C2745 NAND2X1_LOC_647/A INVX1_LOC_476/Y 0.12fF
C2746 INVX1_LOC_108/A INVX1_LOC_63/Y 0.00fF
C2747 INVX1_LOC_579/A INVX1_LOC_354/A 0.03fF
C2748 INVX1_LOC_80/A INVX1_LOC_479/A 0.28fF
C2749 NAND2X1_LOC_768/A INVX1_LOC_479/A 0.16fF
C2750 INVX1_LOC_117/Y INVX1_LOC_328/Y 0.03fF
C2751 INVX1_LOC_375/Y INVX1_LOC_666/Y 0.06fF
C2752 INVX1_LOC_555/Y INVX1_LOC_92/A 0.01fF
C2753 INVX1_LOC_50/Y INVX1_LOC_272/A 0.01fF
C2754 INVX1_LOC_379/A INVX1_LOC_62/Y 0.14fF
C2755 VDD INVX1_LOC_423/A -0.00fF
C2756 INVX1_LOC_35/Y INVX1_LOC_62/Y 0.74fF
C2757 INVX1_LOC_93/Y INVX1_LOC_353/A 0.01fF
C2758 NAND2X1_LOC_307/B INVX1_LOC_89/A 0.00fF
C2759 INVX1_LOC_69/Y INVX1_LOC_44/Y 3.28fF
C2760 INVX1_LOC_211/A NAND2X1_LOC_72/Y 0.03fF
C2761 NAND2X1_LOC_853/a_36_24# INVX1_LOC_79/A 0.00fF
C2762 INVX1_LOC_438/A INVX1_LOC_109/Y 0.34fF
C2763 INVX1_LOC_11/Y NAND2X1_LOC_528/Y 0.24fF
C2764 INVX1_LOC_11/Y INVX1_LOC_479/A 0.20fF
C2765 INVX1_LOC_31/Y NAND2X1_LOC_627/Y 0.01fF
C2766 INVX1_LOC_315/A INVX1_LOC_74/Y 0.05fF
C2767 INVX1_LOC_424/A INVX1_LOC_405/A 0.31fF
C2768 INVX1_LOC_608/A NAND2X1_LOC_372/Y 0.16fF
C2769 INVX1_LOC_32/Y INVX1_LOC_588/A 0.21fF
C2770 INVX1_LOC_62/Y NAND2X1_LOC_253/Y 0.14fF
C2771 INVX1_LOC_379/A NAND2X1_LOC_269/a_36_24# 0.00fF
C2772 NAND2X1_LOC_788/A NAND2X1_LOC_533/a_36_24# 0.02fF
C2773 INVX1_LOC_6/Y INVX1_LOC_388/A 0.03fF
C2774 INVX1_LOC_518/Y INVX1_LOC_9/Y 0.01fF
C2775 INVX1_LOC_618/A NAND2X1_LOC_498/Y 0.01fF
C2776 INVX1_LOC_646/Y NAND2X1_LOC_843/B 0.06fF
C2777 VDD INVX1_LOC_217/Y 0.42fF
C2778 NAND2X1_LOC_632/a_36_24# INVX1_LOC_488/Y 0.01fF
C2779 VDD INVX1_LOC_190/Y 0.21fF
C2780 INVX1_LOC_351/Y INVX1_LOC_211/A 0.04fF
C2781 INVX1_LOC_653/A NAND2X1_LOC_123/B 0.08fF
C2782 INVX1_LOC_6/Y INVX1_LOC_619/Y 0.01fF
C2783 NAND2X1_LOC_701/a_36_24# INVX1_LOC_121/Y 0.00fF
C2784 INVX1_LOC_368/A INVX1_LOC_368/Y 0.04fF
C2785 NAND2X1_LOC_640/a_36_24# INVX1_LOC_62/Y 0.00fF
C2786 INVX1_LOC_412/Y NAND2X1_LOC_567/a_36_24# 0.00fF
C2787 INPUT_0 NAND2X1_LOC_749/Y 0.04fF
C2788 NAND2X1_LOC_433/Y INVX1_LOC_479/A 0.65fF
C2789 VDD INVX1_LOC_72/Y 0.30fF
C2790 NAND2X1_LOC_475/A INVX1_LOC_51/Y 0.04fF
C2791 VDD INVX1_LOC_356/A -0.00fF
C2792 NAND2X1_LOC_751/a_36_24# INVX1_LOC_85/Y 0.00fF
C2793 INVX1_LOC_662/A INVX1_LOC_92/A 0.14fF
C2794 NAND2X1_LOC_592/B INVX1_LOC_45/Y 0.01fF
C2795 NAND2X1_LOC_261/Y INVX1_LOC_445/A 0.01fF
C2796 INVX1_LOC_266/A NAND2X1_LOC_475/A 0.11fF
C2797 INVX1_LOC_32/A INVX1_LOC_84/A 0.01fF
C2798 INVX1_LOC_449/A INVX1_LOC_448/Y 0.13fF
C2799 VDD INVX1_LOC_519/A 0.43fF
C2800 INVX1_LOC_435/Y NAND2X1_LOC_486/B 0.09fF
C2801 INVX1_LOC_206/Y INVX1_LOC_318/Y 0.01fF
C2802 VDD NAND2X1_LOC_296/Y 0.01fF
C2803 NAND2X1_LOC_528/Y INVX1_LOC_231/Y 0.02fF
C2804 INVX1_LOC_374/A INVX1_LOC_76/Y 0.03fF
C2805 VDD INVX1_LOC_323/Y 0.20fF
C2806 INVX1_LOC_279/A INVX1_LOC_452/A 0.01fF
C2807 INVX1_LOC_502/Y INVX1_LOC_51/Y 0.03fF
C2808 NAND2X1_LOC_537/A INVX1_LOC_99/Y 0.01fF
C2809 INVX1_LOC_206/Y INVX1_LOC_455/Y 0.04fF
C2810 INVX1_LOC_617/A INVX1_LOC_362/Y 0.05fF
C2811 NAND2X1_LOC_788/A INVX1_LOC_252/Y 0.16fF
C2812 INVX1_LOC_4/Y INVX1_LOC_5/Y 0.01fF
C2813 NAND2X1_LOC_142/Y INVX1_LOC_101/Y 0.01fF
C2814 INVX1_LOC_614/A INVX1_LOC_523/A 0.03fF
C2815 INVX1_LOC_578/A NAND2X1_LOC_545/B 0.04fF
C2816 NAND2X1_LOC_638/A INVX1_LOC_395/A 0.01fF
C2817 INVX1_LOC_202/Y INVX1_LOC_560/Y 0.15fF
C2818 INPUT_0 INVX1_LOC_99/A 0.03fF
C2819 INVX1_LOC_229/Y INVX1_LOC_65/Y 0.03fF
C2820 INVX1_LOC_68/Y INVX1_LOC_524/Y 0.08fF
C2821 INVX1_LOC_577/A INVX1_LOC_155/Y 0.01fF
C2822 NAND2X1_LOC_746/a_36_24# INVX1_LOC_48/Y 0.00fF
C2823 NAND2X1_LOC_475/A NAND2X1_LOC_267/a_36_24# 0.00fF
C2824 INVX1_LOC_224/Y INVX1_LOC_98/Y 0.12fF
C2825 NAND2X1_LOC_781/B INVX1_LOC_93/Y 0.03fF
C2826 INVX1_LOC_409/Y INVX1_LOC_93/Y 0.05fF
C2827 INVX1_LOC_454/A INVX1_LOC_674/A 0.18fF
C2828 NAND2X1_LOC_183/a_36_24# INVX1_LOC_48/Y 0.01fF
C2829 NAND2X1_LOC_393/a_36_24# INVX1_LOC_172/A 0.00fF
C2830 INVX1_LOC_450/A INVX1_LOC_385/Y 0.03fF
C2831 NAND2X1_LOC_543/B INVX1_LOC_31/Y 0.45fF
C2832 INVX1_LOC_107/A INVX1_LOC_145/Y 0.00fF
C2833 INVX1_LOC_45/Y NAND2X1_LOC_616/Y 0.05fF
C2834 INVX1_LOC_45/Y INVX1_LOC_232/Y 0.01fF
C2835 INPUT_0 INVX1_LOC_137/Y 0.06fF
C2836 INVX1_LOC_340/Y INVX1_LOC_632/A 0.07fF
C2837 NAND2X1_LOC_108/Y INVX1_LOC_99/Y 0.05fF
C2838 INVX1_LOC_578/A INVX1_LOC_98/Y 0.10fF
C2839 INVX1_LOC_405/A INVX1_LOC_49/Y 0.03fF
C2840 NAND2X1_LOC_763/Y INVX1_LOC_117/Y 0.01fF
C2841 INVX1_LOC_442/A INVX1_LOC_252/Y 0.07fF
C2842 INVX1_LOC_463/A INVX1_LOC_47/Y 0.98fF
C2843 INVX1_LOC_553/Y INVX1_LOC_361/Y 0.00fF
C2844 NAND2X1_LOC_573/a_36_24# INVX1_LOC_32/Y 0.01fF
C2845 INVX1_LOC_127/A INVX1_LOC_105/A 0.01fF
C2846 NAND2X1_LOC_537/A INVX1_LOC_47/Y 0.02fF
C2847 INVX1_LOC_560/A INVX1_LOC_603/A 0.03fF
C2848 NAND2X1_LOC_770/A INVX1_LOC_63/Y 0.12fF
C2849 VDD NAND2X1_LOC_846/A -0.00fF
C2850 INVX1_LOC_409/Y INVX1_LOC_675/A 0.08fF
C2851 INVX1_LOC_666/A INVX1_LOC_145/Y 0.02fF
C2852 INVX1_LOC_361/Y INVX1_LOC_375/A 0.03fF
C2853 INVX1_LOC_372/Y INVX1_LOC_80/A 0.21fF
C2854 INVX1_LOC_68/Y INVX1_LOC_400/A 0.05fF
C2855 VDD INVX1_LOC_659/A 0.04fF
C2856 NAND2X1_LOC_580/a_36_24# INVX1_LOC_452/A 0.01fF
C2857 INVX1_LOC_521/Y INVX1_LOC_117/Y 0.03fF
C2858 NAND2X1_LOC_13/Y INVX1_LOC_99/Y 0.10fF
C2859 NAND2X1_LOC_710/a_36_24# INVX1_LOC_166/A 0.00fF
C2860 INVX1_LOC_370/Y INVX1_LOC_686/A 0.04fF
C2861 NAND2X1_LOC_612/A INVX1_LOC_492/Y 0.02fF
C2862 INVX1_LOC_459/Y INVX1_LOC_50/Y 0.01fF
C2863 INVX1_LOC_117/Y INVX1_LOC_266/Y 0.07fF
C2864 NAND2X1_LOC_107/Y INVX1_LOC_679/Y 0.03fF
C2865 INVX1_LOC_17/Y INVX1_LOC_293/Y 0.17fF
C2866 NAND2X1_LOC_165/Y INVX1_LOC_94/A 0.04fF
C2867 NAND2X1_LOC_732/a_36_24# NAND2X1_LOC_152/B 0.01fF
C2868 INVX1_LOC_68/Y NAND2X1_LOC_289/a_36_24# 0.00fF
C2869 INVX1_LOC_355/A INVX1_LOC_47/Y 0.05fF
C2870 INVX1_LOC_206/Y INVX1_LOC_351/A 0.12fF
C2871 INVX1_LOC_14/A INVX1_LOC_16/Y 0.20fF
C2872 INVX1_LOC_53/A INVX1_LOC_53/Y 0.05fF
C2873 INVX1_LOC_584/Y INVX1_LOC_58/Y 0.02fF
C2874 NAND2X1_LOC_616/Y NAND2X1_LOC_69/Y 0.03fF
C2875 NAND2X1_LOC_13/Y INVX1_LOC_123/A 0.00fF
C2876 INVX1_LOC_275/Y INVX1_LOC_197/Y 0.03fF
C2877 INVX1_LOC_11/Y INVX1_LOC_12/Y 0.07fF
C2878 INVX1_LOC_400/A INVX1_LOC_600/A 0.04fF
C2879 INVX1_LOC_206/Y INVX1_LOC_90/Y 0.15fF
C2880 INVX1_LOC_547/A NAND2X1_LOC_253/Y 0.11fF
C2881 INVX1_LOC_171/Y INVX1_LOC_6/Y 0.01fF
C2882 INVX1_LOC_103/A INVX1_LOC_26/Y 0.02fF
C2883 INVX1_LOC_213/Y INVX1_LOC_679/Y 0.02fF
C2884 INVX1_LOC_53/Y INVX1_LOC_50/Y 6.38fF
C2885 INVX1_LOC_395/A INVX1_LOC_353/A 0.02fF
C2886 NAND2X1_LOC_381/a_36_24# INVX1_LOC_117/Y 0.01fF
C2887 INVX1_LOC_468/Y INVX1_LOC_98/Y 0.05fF
C2888 NAND2X1_LOC_148/A INPUT_1 0.11fF
C2889 INVX1_LOC_378/Y INVX1_LOC_378/A 0.01fF
C2890 INVX1_LOC_116/Y INVX1_LOC_252/Y 0.03fF
C2891 INVX1_LOC_586/A INVX1_LOC_44/Y 3.25fF
C2892 INVX1_LOC_581/A NAND2X1_LOC_708/a_36_24# 0.00fF
C2893 INVX1_LOC_103/Y INVX1_LOC_519/A 0.02fF
C2894 NAND2X1_LOC_673/A INVX1_LOC_145/Y 0.01fF
C2895 NAND2X1_LOC_557/a_36_24# INVX1_LOC_600/A 0.01fF
C2896 NAND2X1_LOC_791/B INVX1_LOC_89/Y 0.01fF
C2897 NAND2X1_LOC_448/A INVX1_LOC_259/Y 0.06fF
C2898 INVX1_LOC_25/Y INVX1_LOC_40/Y 0.06fF
C2899 INVX1_LOC_155/Y INVX1_LOC_48/Y 1.93fF
C2900 INVX1_LOC_93/Y NAND2X1_LOC_302/A 0.04fF
C2901 INVX1_LOC_649/Y INVX1_LOC_6/Y 0.01fF
C2902 INVX1_LOC_355/A INVX1_LOC_119/Y 0.02fF
C2903 NAND2X1_LOC_130/Y INVX1_LOC_93/Y 0.03fF
C2904 INVX1_LOC_391/A INVX1_LOC_80/A 0.03fF
C2905 INVX1_LOC_7/Y INVX1_LOC_86/Y 0.01fF
C2906 INVX1_LOC_366/A INVX1_LOC_179/Y 0.01fF
C2907 INVX1_LOC_84/A INVX1_LOC_49/Y 0.06fF
C2908 NAND2X1_LOC_542/A INVX1_LOC_134/Y 0.02fF
C2909 NAND2X1_LOC_677/Y INVX1_LOC_6/Y 0.00fF
C2910 INVX1_LOC_587/Y NAND2X1_LOC_837/B 0.27fF
C2911 NAND2X1_LOC_612/A NAND2X1_LOC_647/A 0.00fF
C2912 NAND2X1_LOC_285/A INVX1_LOC_145/Y 0.01fF
C2913 INVX1_LOC_460/Y INVX1_LOC_50/Y 0.00fF
C2914 NAND2X1_LOC_32/Y INVX1_LOC_54/Y 0.00fF
C2915 INVX1_LOC_235/Y INVX1_LOC_26/Y 0.07fF
C2916 INVX1_LOC_137/Y INVX1_LOC_498/A 0.05fF
C2917 INVX1_LOC_89/Y INVX1_LOC_252/A 0.03fF
C2918 NAND2X1_LOC_619/Y INVX1_LOC_480/Y 0.02fF
C2919 INVX1_LOC_134/Y INVX1_LOC_376/Y 0.07fF
C2920 NAND2X1_LOC_399/B INVX1_LOC_63/Y 0.05fF
C2921 INVX1_LOC_193/A INVX1_LOC_46/Y 0.00fF
C2922 INVX1_LOC_62/A INVX1_LOC_46/Y 0.01fF
C2923 INVX1_LOC_149/Y INVX1_LOC_491/Y 0.01fF
C2924 INVX1_LOC_11/Y INVX1_LOC_391/A 0.03fF
C2925 INVX1_LOC_63/Y INVX1_LOC_7/Y 5.21fF
C2926 INVX1_LOC_255/A INVX1_LOC_252/Y 0.07fF
C2927 INVX1_LOC_491/A INVX1_LOC_633/Y 0.02fF
C2928 INVX1_LOC_63/Y INVX1_LOC_228/A 0.07fF
C2929 INVX1_LOC_49/Y NAND2X1_LOC_67/Y 0.02fF
C2930 INVX1_LOC_69/Y INVX1_LOC_656/Y 0.18fF
C2931 INVX1_LOC_256/A INVX1_LOC_63/Y 0.01fF
C2932 INVX1_LOC_145/Y INVX1_LOC_168/Y 0.13fF
C2933 INVX1_LOC_63/Y NAND2X1_LOC_259/A 0.00fF
C2934 INVX1_LOC_531/A INVX1_LOC_9/Y 0.01fF
C2935 NAND2X1_LOC_704/B INVX1_LOC_479/A 0.03fF
C2936 NAND2X1_LOC_619/Y INVX1_LOC_169/Y 0.06fF
C2937 INVX1_LOC_300/Y INVX1_LOC_685/A 0.01fF
C2938 INVX1_LOC_328/Y INVX1_LOC_281/Y 0.31fF
C2939 INVX1_LOC_457/Y INVX1_LOC_636/A -0.06fF
C2940 INVX1_LOC_11/Y INVX1_LOC_170/A 0.03fF
C2941 INVX1_LOC_93/Y INVX1_LOC_484/A -0.00fF
C2942 INVX1_LOC_153/Y INVX1_LOC_154/Y 0.09fF
C2943 NAND2X1_LOC_532/Y INVX1_LOC_46/Y 0.01fF
C2944 NAND2X1_LOC_787/a_36_24# INVX1_LOC_9/Y 0.00fF
C2945 INVX1_LOC_6/Y INVX1_LOC_199/A 0.02fF
C2946 INVX1_LOC_174/A INVX1_LOC_531/Y 0.00fF
C2947 INVX1_LOC_544/Y INPUT_1 0.18fF
C2948 INVX1_LOC_386/Y INVX1_LOC_430/A 0.22fF
C2949 INVX1_LOC_345/Y INVX1_LOC_63/Y 0.01fF
C2950 NAND2X1_LOC_376/B INVX1_LOC_46/Y 0.01fF
C2951 INVX1_LOC_242/Y INVX1_LOC_230/A 0.01fF
C2952 INVX1_LOC_89/Y INVX1_LOC_6/Y 0.06fF
C2953 INVX1_LOC_54/Y NAND2X1_LOC_192/A 0.03fF
C2954 INVX1_LOC_32/Y INVX1_LOC_63/Y 0.34fF
C2955 NAND2X1_LOC_388/A INVX1_LOC_199/Y 1.46fF
C2956 INVX1_LOC_81/Y INVX1_LOC_26/Y 0.04fF
C2957 INVX1_LOC_169/Y NAND2X1_LOC_618/a_36_24# 0.01fF
C2958 INVX1_LOC_298/A INPUT_5 0.25fF
C2959 NAND2X1_LOC_606/Y INVX1_LOC_114/A 0.19fF
C2960 INVX1_LOC_662/A INPUT_1 0.08fF
C2961 INVX1_LOC_671/A INVX1_LOC_664/A 0.02fF
C2962 INVX1_LOC_520/Y INVX1_LOC_212/Y 0.02fF
C2963 INVX1_LOC_338/A INVX1_LOC_62/Y 0.03fF
C2964 NAND2X1_LOC_175/a_36_24# INVX1_LOC_636/A 0.01fF
C2965 INVX1_LOC_157/Y INVX1_LOC_44/Y 0.06fF
C2966 INVX1_LOC_254/Y INVX1_LOC_319/A 0.01fF
C2967 INVX1_LOC_214/Y INVX1_LOC_62/Y 0.01fF
C2968 INVX1_LOC_197/Y INVX1_LOC_274/Y 0.06fF
C2969 INVX1_LOC_44/Y NAND2X1_LOC_825/a_36_24# 0.01fF
C2970 INVX1_LOC_179/Y INVX1_LOC_6/Y 0.11fF
C2971 INVX1_LOC_62/Y NAND2X1_LOC_837/B 0.76fF
C2972 INVX1_LOC_607/Y INVX1_LOC_647/Y 0.06fF
C2973 INVX1_LOC_62/Y INVX1_LOC_360/A 0.01fF
C2974 INVX1_LOC_41/Y NAND2X1_LOC_444/A 0.01fF
C2975 INVX1_LOC_368/Y INVX1_LOC_50/Y 0.09fF
C2976 INVX1_LOC_354/Y INVX1_LOC_74/Y 0.01fF
C2977 INVX1_LOC_410/A INVX1_LOC_100/Y 0.02fF
C2978 NAND2X1_LOC_34/a_36_24# INVX1_LOC_395/A 0.00fF
C2979 NAND2X1_LOC_833/B NAND2X1_LOC_258/a_36_24# 0.00fF
C2980 INVX1_LOC_664/A INVX1_LOC_664/Y 0.03fF
C2981 INVX1_LOC_273/A NAND2X1_LOC_227/a_36_24# 0.00fF
C2982 INVX1_LOC_659/A INVX1_LOC_635/Y 0.09fF
C2983 INVX1_LOC_183/A INVX1_LOC_41/Y 0.03fF
C2984 NAND2X1_LOC_322/Y INVX1_LOC_395/A 0.15fF
C2985 INVX1_LOC_447/A NAND2X1_LOC_457/A 0.03fF
C2986 VDD INVX1_LOC_445/A 0.00fF
C2987 INVX1_LOC_389/Y INVX1_LOC_41/Y 0.01fF
C2988 INVX1_LOC_280/A INVX1_LOC_245/A 0.00fF
C2989 INVX1_LOC_46/Y INVX1_LOC_76/A 0.01fF
C2990 INVX1_LOC_183/A NAND2X1_LOC_403/a_36_24# 0.00fF
C2991 NAND2X1_LOC_71/a_36_24# INVX1_LOC_9/Y 0.00fF
C2992 INVX1_LOC_405/A INVX1_LOC_76/Y 0.00fF
C2993 INVX1_LOC_412/Y INVX1_LOC_412/A 0.05fF
C2994 INVX1_LOC_560/Y INVX1_LOC_250/A 0.12fF
C2995 INVX1_LOC_20/Y INVX1_LOC_459/A 0.02fF
C2996 NAND2X1_LOC_773/a_36_24# INVX1_LOC_366/A 0.00fF
C2997 INVX1_LOC_435/Y INVX1_LOC_224/Y 0.01fF
C2998 INVX1_LOC_9/Y INVX1_LOC_488/Y 0.10fF
C2999 VDD NAND2X1_LOC_97/A -0.00fF
C3000 INVX1_LOC_479/A INVX1_LOC_319/A 0.04fF
C3001 INVX1_LOC_560/Y INVX1_LOC_76/Y 0.07fF
C3002 INVX1_LOC_266/A NAND2X1_LOC_543/B 0.66fF
C3003 VDD NAND2X1_LOC_39/Y 0.01fF
C3004 NAND2X1_LOC_13/Y NAND2X1_LOC_475/A 0.39fF
C3005 INVX1_LOC_271/A NAND2X1_LOC_337/a_36_24# 0.01fF
C3006 VDD INVX1_LOC_574/Y 0.21fF
C3007 NAND2X1_LOC_690/Y INVX1_LOC_542/A 0.12fF
C3008 INVX1_LOC_395/A INVX1_LOC_88/Y 0.01fF
C3009 INVX1_LOC_117/Y INVX1_LOC_109/Y 0.10fF
C3010 INVX1_LOC_96/Y INVX1_LOC_586/A 0.58fF
C3011 NAND2X1_LOC_122/Y INVX1_LOC_45/Y 0.03fF
C3012 NAND2X1_LOC_546/a_36_24# INVX1_LOC_362/Y 0.00fF
C3013 NAND2X1_LOC_545/A INVX1_LOC_92/A 0.04fF
C3014 INVX1_LOC_438/A INVX1_LOC_53/Y 0.07fF
C3015 INVX1_LOC_312/Y INVX1_LOC_118/Y 0.03fF
C3016 VDD NAND2X1_LOC_147/B 0.03fF
C3017 INVX1_LOC_206/Y NAND2X1_LOC_545/B 0.01fF
C3018 INVX1_LOC_586/A NAND2X1_LOC_685/B 0.05fF
C3019 INVX1_LOC_578/A INVX1_LOC_596/A 0.02fF
C3020 NAND2X1_LOC_46/a_36_24# INVX1_LOC_80/A 0.01fF
C3021 INVX1_LOC_560/Y INVX1_LOC_559/A 0.05fF
C3022 INVX1_LOC_604/A INVX1_LOC_80/A 0.07fF
C3023 NAND2X1_LOC_516/Y NAND2X1_LOC_307/A 0.00fF
C3024 INVX1_LOC_554/A INVX1_LOC_117/Y 0.03fF
C3025 NAND2X1_LOC_475/A NAND2X1_LOC_860/a_36_24# 0.00fF
C3026 INVX1_LOC_666/Y INVX1_LOC_92/A 0.03fF
C3027 INVX1_LOC_446/A INVX1_LOC_32/Y 0.07fF
C3028 INVX1_LOC_238/A INVX1_LOC_556/Y 0.01fF
C3029 INVX1_LOC_20/Y NAND2X1_LOC_492/a_36_24# 0.00fF
C3030 INVX1_LOC_206/Y INVX1_LOC_98/Y 0.39fF
C3031 INVX1_LOC_404/Y INVX1_LOC_379/A 0.03fF
C3032 NAND2X1_LOC_317/A INVX1_LOC_251/Y 0.27fF
C3033 INVX1_LOC_84/A INVX1_LOC_76/Y 0.09fF
C3034 NAND2X1_LOC_391/A INVX1_LOC_586/A 0.35fF
C3035 INPUT_3 INVX1_LOC_325/Y 0.28fF
C3036 INVX1_LOC_147/A INVX1_LOC_586/A 0.01fF
C3037 NAND2X1_LOC_596/Y INVX1_LOC_513/A 0.10fF
C3038 INVX1_LOC_256/A INVX1_LOC_374/A 0.01fF
C3039 INVX1_LOC_51/Y INVX1_LOC_469/A 0.09fF
C3040 INVX1_LOC_248/Y INVX1_LOC_45/Y 0.03fF
C3041 NAND2X1_LOC_325/B NAND2X1_LOC_332/B 0.06fF
C3042 INVX1_LOC_20/Y INVX1_LOC_635/A 0.06fF
C3043 NAND2X1_LOC_403/A INVX1_LOC_322/Y 0.23fF
C3044 INVX1_LOC_205/Y INVX1_LOC_366/A 0.01fF
C3045 INVX1_LOC_312/A INVX1_LOC_312/Y 0.14fF
C3046 NAND2X1_LOC_165/a_36_24# INVX1_LOC_94/A 0.00fF
C3047 NAND2X1_LOC_780/B INVX1_LOC_6/Y 0.03fF
C3048 INVX1_LOC_552/Y INVX1_LOC_32/Y 0.02fF
C3049 INVX1_LOC_259/A INVX1_LOC_259/Y 0.01fF
C3050 INVX1_LOC_564/A NAND2X1_LOC_333/A 0.00fF
C3051 NAND2X1_LOC_475/A INVX1_LOC_380/Y 0.15fF
C3052 NAND2X1_LOC_331/A INVX1_LOC_572/Y 0.27fF
C3053 INVX1_LOC_374/A INVX1_LOC_345/Y 0.01fF
C3054 INVX1_LOC_578/A NAND2X1_LOC_442/a_36_24# 0.01fF
C3055 INVX1_LOC_53/Y NAND2X1_LOC_513/A 0.03fF
C3056 INVX1_LOC_406/Y INVX1_LOC_442/Y 0.00fF
C3057 INVX1_LOC_366/A INVX1_LOC_194/Y 0.01fF
C3058 INVX1_LOC_20/Y INVX1_LOC_230/A 0.06fF
C3059 NAND2X1_LOC_475/A INVX1_LOC_361/A 0.07fF
C3060 INVX1_LOC_235/Y NAND2X1_LOC_275/Y 0.01fF
C3061 INVX1_LOC_206/Y INVX1_LOC_338/Y 0.07fF
C3062 INVX1_LOC_288/A INVX1_LOC_355/Y 0.00fF
C3063 INVX1_LOC_686/A INVX1_LOC_98/Y 0.10fF
C3064 INVX1_LOC_522/A INVX1_LOC_515/A 0.39fF
C3065 INVX1_LOC_137/A INVX1_LOC_6/Y 0.03fF
C3066 INVX1_LOC_602/A INVX1_LOC_342/Y 0.08fF
C3067 INVX1_LOC_54/Y INVX1_LOC_381/A 0.10fF
C3068 INVX1_LOC_419/A INVX1_LOC_442/A 0.01fF
C3069 INVX1_LOC_62/Y INVX1_LOC_220/A 0.32fF
C3070 INVX1_LOC_521/Y INVX1_LOC_58/Y 0.01fF
C3071 INVX1_LOC_80/A INVX1_LOC_159/A 0.04fF
C3072 NAND2X1_LOC_399/B NAND2X1_LOC_399/a_36_24# 0.02fF
C3073 INVX1_LOC_406/A INVX1_LOC_384/A 0.05fF
C3074 INVX1_LOC_289/A NAND2X1_LOC_355/a_36_24# 0.00fF
C3075 INVX1_LOC_313/Y INVX1_LOC_12/Y 0.01fF
C3076 INVX1_LOC_613/Y INVX1_LOC_137/Y 0.03fF
C3077 INVX1_LOC_105/A INVX1_LOC_519/A 0.03fF
C3078 NAND2X1_LOC_673/B NAND2X1_LOC_616/Y 0.07fF
C3079 INVX1_LOC_80/A NAND2X1_LOC_615/B 0.60fF
C3080 INVX1_LOC_7/Y NAND2X1_LOC_414/a_36_24# 0.01fF
C3081 INVX1_LOC_266/Y INVX1_LOC_58/Y 0.03fF
C3082 INVX1_LOC_397/A INVX1_LOC_351/A 0.06fF
C3083 INVX1_LOC_300/A INVX1_LOC_230/A -0.00fF
C3084 INPUT_0 INVX1_LOC_502/A 0.07fF
C3085 INVX1_LOC_584/Y INVX1_LOC_245/A 0.09fF
C3086 INVX1_LOC_323/Y INVX1_LOC_171/A 0.06fF
C3087 NAND2X1_LOC_378/Y INVX1_LOC_365/A 0.00fF
C3088 INVX1_LOC_595/A INVX1_LOC_18/Y 0.00fF
C3089 INVX1_LOC_434/A INVX1_LOC_62/Y 0.03fF
C3090 INVX1_LOC_575/A INVX1_LOC_35/Y 0.26fF
C3091 INVX1_LOC_651/Y INVX1_LOC_58/Y 0.09fF
C3092 INVX1_LOC_76/Y INVX1_LOC_496/A 0.04fF
C3093 INVX1_LOC_366/A INVX1_LOC_44/Y 0.03fF
C3094 INVX1_LOC_52/Y INVX1_LOC_62/Y 0.01fF
C3095 INVX1_LOC_133/A NAND2X1_LOC_847/A 0.12fF
C3096 INVX1_LOC_114/Y NAND2X1_LOC_121/Y 0.01fF
C3097 NAND2X1_LOC_498/Y NAND2X1_LOC_301/B 0.02fF
C3098 INVX1_LOC_393/A NAND2X1_LOC_274/B 0.01fF
C3099 INVX1_LOC_462/Y INVX1_LOC_638/A 0.01fF
C3100 INVX1_LOC_35/Y INVX1_LOC_480/Y 0.01fF
C3101 INVX1_LOC_31/Y INVX1_LOC_600/A 0.10fF
C3102 INVX1_LOC_80/A INVX1_LOC_66/A 0.11fF
C3103 INVX1_LOC_11/Y INVX1_LOC_159/A 0.00fF
C3104 INVX1_LOC_51/Y INVX1_LOC_353/A 0.00fF
C3105 INVX1_LOC_501/Y INVX1_LOC_498/Y 0.08fF
C3106 INVX1_LOC_90/Y INVX1_LOC_94/A 0.03fF
C3107 NAND2X1_LOC_315/a_36_24# INVX1_LOC_9/Y 0.00fF
C3108 INVX1_LOC_272/Y INVX1_LOC_44/Y 0.07fF
C3109 NAND2X1_LOC_635/B INVX1_LOC_685/Y 0.02fF
C3110 INVX1_LOC_229/Y INVX1_LOC_63/Y 0.01fF
C3111 NAND2X1_LOC_791/B INVX1_LOC_44/Y 0.04fF
C3112 INVX1_LOC_541/Y INVX1_LOC_513/Y 0.04fF
C3113 INVX1_LOC_11/Y NAND2X1_LOC_615/B 0.28fF
C3114 INVX1_LOC_413/Y INVX1_LOC_41/Y 0.02fF
C3115 NAND2X1_LOC_324/B INVX1_LOC_63/Y 0.28fF
C3116 INVX1_LOC_205/Y INVX1_LOC_6/Y 0.02fF
C3117 NAND2X1_LOC_521/Y INVX1_LOC_367/Y 0.19fF
C3118 INVX1_LOC_35/Y INVX1_LOC_169/Y 0.04fF
C3119 INVX1_LOC_670/A INVX1_LOC_371/A 0.16fF
C3120 INVX1_LOC_93/Y NAND2X1_LOC_708/A 0.01fF
C3121 INVX1_LOC_406/A INVX1_LOC_145/Y 0.00fF
C3122 NAND2X1_LOC_846/a_36_24# INVX1_LOC_655/A 0.01fF
C3123 INVX1_LOC_11/Y INVX1_LOC_127/Y 0.05fF
C3124 INVX1_LOC_607/Y NAND2X1_LOC_342/A 0.04fF
C3125 INVX1_LOC_491/Y INVX1_LOC_493/Y 0.09fF
C3126 INVX1_LOC_69/Y INVX1_LOC_252/Y 0.03fF
C3127 NAND2X1_LOC_706/B NAND2X1_LOC_693/a_36_24# 0.02fF
C3128 NAND2X1_LOC_79/B INVX1_LOC_210/A 0.01fF
C3129 INVX1_LOC_6/Y INVX1_LOC_194/Y 0.05fF
C3130 INVX1_LOC_11/Y INVX1_LOC_66/A 0.14fF
C3131 INVX1_LOC_14/A INVX1_LOC_338/Y 0.02fF
C3132 INVX1_LOC_58/Y INVX1_LOC_352/A 0.01fF
C3133 INVX1_LOC_21/Y INVX1_LOC_183/A 0.07fF
C3134 INVX1_LOC_99/Y INVX1_LOC_480/A 0.01fF
C3135 INVX1_LOC_469/Y INVX1_LOC_354/Y 0.01fF
C3136 NAND2X1_LOC_400/B INVX1_LOC_327/Y 0.08fF
C3137 INVX1_LOC_11/Y INVX1_LOC_296/A 0.01fF
C3138 INVX1_LOC_63/Y NAND2X1_LOC_226/Y 0.01fF
C3139 NAND2X1_LOC_130/Y INVX1_LOC_128/A 0.01fF
C3140 INVX1_LOC_17/Y INVX1_LOC_682/A 0.00fF
C3141 INVX1_LOC_21/Y INVX1_LOC_389/Y 0.01fF
C3142 NAND2X1_LOC_488/a_36_24# INVX1_LOC_600/A 0.00fF
C3143 NAND2X1_LOC_325/B INVX1_LOC_242/Y 1.24fF
C3144 INVX1_LOC_335/A INVX1_LOC_58/Y 0.03fF
C3145 INVX1_LOC_346/A INVX1_LOC_513/A 0.21fF
C3146 INVX1_LOC_298/A NAND2X1_LOC_425/a_36_24# 0.00fF
C3147 INVX1_LOC_565/A INVX1_LOC_26/Y 0.01fF
C3148 INVX1_LOC_117/Y INVX1_LOC_199/Y 0.27fF
C3149 INVX1_LOC_50/Y NAND2X1_LOC_790/a_36_24# 0.00fF
C3150 INVX1_LOC_12/Y INVX1_LOC_319/A 0.01fF
C3151 INVX1_LOC_174/A INVX1_LOC_41/Y 1.41fF
C3152 INVX1_LOC_421/A NAND2X1_LOC_346/a_36_24# 0.00fF
C3153 INVX1_LOC_603/Y INVX1_LOC_531/Y 0.07fF
C3154 INVX1_LOC_447/Y INVX1_LOC_100/Y 0.01fF
C3155 INVX1_LOC_176/A INVX1_LOC_79/A 0.07fF
C3156 INVX1_LOC_17/Y INVX1_LOC_112/Y 0.10fF
C3157 INVX1_LOC_662/A INVX1_LOC_50/Y 0.03fF
C3158 INVX1_LOC_100/Y NAND2X1_LOC_602/A 0.01fF
C3159 INVX1_LOC_600/Y INVX1_LOC_274/Y 0.00fF
C3160 GATE_662 INVX1_LOC_58/Y 0.01fF
C3161 INVX1_LOC_47/Y NAND2X1_LOC_449/B 0.03fF
C3162 INVX1_LOC_419/A INVX1_LOC_255/A 0.01fF
C3163 INVX1_LOC_69/Y NAND2X1_LOC_827/Y 0.02fF
C3164 INVX1_LOC_62/Y INVX1_LOC_115/Y 0.01fF
C3165 INVX1_LOC_349/A INVX1_LOC_79/A 0.01fF
C3166 INVX1_LOC_291/A NAND2X1_LOC_96/a_36_24# 0.01fF
C3167 INVX1_LOC_44/Y INVX1_LOC_6/Y 0.03fF
C3168 INVX1_LOC_403/Y NAND2X1_LOC_136/Y 0.01fF
C3169 INVX1_LOC_54/Y INVX1_LOC_100/Y 1.26fF
C3170 INVX1_LOC_62/Y INVX1_LOC_350/A 0.01fF
C3171 NAND2X1_LOC_545/A INPUT_1 0.99fF
C3172 NAND2X1_LOC_334/A INVX1_LOC_338/Y 0.12fF
C3173 INVX1_LOC_89/Y INVX1_LOC_557/Y 0.01fF
C3174 INVX1_LOC_145/Y NAND2X1_LOC_234/Y 0.03fF
C3175 INVX1_LOC_93/Y INVX1_LOC_369/Y 0.07fF
C3176 INVX1_LOC_6/Y INVX1_LOC_48/A 0.05fF
C3177 NAND2X1_LOC_833/B NAND2X1_LOC_253/Y 0.07fF
C3178 NAND2X1_LOC_387/Y INVX1_LOC_531/Y 0.06fF
C3179 NAND2X1_LOC_171/a_36_24# INVX1_LOC_79/A 0.00fF
C3180 INVX1_LOC_54/Y INVX1_LOC_74/Y 1.61fF
C3181 INPUT_1 INVX1_LOC_653/Y 0.14fF
C3182 NAND2X1_LOC_614/a_36_24# INVX1_LOC_74/Y 0.00fF
C3183 INVX1_LOC_361/Y INVX1_LOC_479/A 0.07fF
C3184 INVX1_LOC_119/Y NAND2X1_LOC_449/B 0.21fF
C3185 INVX1_LOC_257/A INVX1_LOC_100/Y 0.08fF
C3186 INPUT_1 INVX1_LOC_666/Y 0.11fF
C3187 INVX1_LOC_223/Y INVX1_LOC_9/Y 0.15fF
C3188 INVX1_LOC_180/Y INVX1_LOC_616/Y 0.99fF
C3189 INVX1_LOC_328/Y INVX1_LOC_245/A 0.03fF
C3190 NAND2X1_LOC_66/Y INVX1_LOC_480/A 0.01fF
C3191 NAND2X1_LOC_286/A INVX1_LOC_669/A 0.04fF
C3192 INVX1_LOC_261/Y INVX1_LOC_479/A 0.15fF
C3193 INVX1_LOC_338/Y NAND2X1_LOC_609/B -0.01fF
C3194 INVX1_LOC_457/Y NAND2X1_LOC_591/B 0.00fF
C3195 NAND2X1_LOC_333/A INVX1_LOC_91/Y 0.55fF
C3196 INVX1_LOC_507/Y INVX1_LOC_62/Y 0.01fF
C3197 INPUT_0 INVX1_LOC_388/Y 0.04fF
C3198 INVX1_LOC_224/Y NAND2X1_LOC_76/B 0.00fF
C3199 INVX1_LOC_531/Y NAND2X1_LOC_845/B 0.02fF
C3200 INVX1_LOC_107/Y INVX1_LOC_109/A 0.01fF
C3201 INVX1_LOC_409/Y INVX1_LOC_51/Y 0.32fF
C3202 INVX1_LOC_89/Y INVX1_LOC_636/A 0.42fF
C3203 INVX1_LOC_153/Y INVX1_LOC_91/A 0.09fF
C3204 INVX1_LOC_150/A INVX1_LOC_45/Y 0.11fF
C3205 INVX1_LOC_152/Y INVX1_LOC_586/A 0.03fF
C3206 INVX1_LOC_20/Y INVX1_LOC_465/Y 0.09fF
C3207 VDD NAND2X1_LOC_391/B 0.01fF
C3208 INVX1_LOC_20/Y NAND2X1_LOC_170/a_36_24# 0.00fF
C3209 INVX1_LOC_266/A NAND2X1_LOC_322/Y 0.43fF
C3210 INVX1_LOC_375/A INVX1_LOC_618/Y 0.01fF
C3211 INVX1_LOC_523/A INVX1_LOC_185/Y 0.03fF
C3212 NAND2X1_LOC_788/A INVX1_LOC_80/A 0.03fF
C3213 INVX1_LOC_68/Y NAND2X1_LOC_505/Y 0.00fF
C3214 INVX1_LOC_457/Y INVX1_LOC_566/A 0.04fF
C3215 INVX1_LOC_206/Y INVX1_LOC_596/A 0.03fF
C3216 NAND2X1_LOC_843/B INVX1_LOC_212/A 0.00fF
C3217 INVX1_LOC_74/Y NAND2X1_LOC_428/a_36_24# 0.00fF
C3218 INVX1_LOC_20/Y INVX1_LOC_107/A 0.01fF
C3219 INVX1_LOC_257/Y NAND2X1_LOC_307/A 0.46fF
C3220 INVX1_LOC_68/Y INVX1_LOC_51/Y 0.00fF
C3221 NAND2X1_LOC_498/Y INVX1_LOC_551/Y 0.10fF
C3222 NAND2X1_LOC_336/B INVX1_LOC_410/Y 0.03fF
C3223 NAND2X1_LOC_700/a_36_24# INVX1_LOC_375/A 0.00fF
C3224 INVX1_LOC_425/A INVX1_LOC_586/A 0.01fF
C3225 INVX1_LOC_45/Y INVX1_LOC_356/A 0.00fF
C3226 NAND2X1_LOC_457/A NAND2X1_LOC_658/a_36_24# 0.00fF
C3227 INVX1_LOC_428/A INVX1_LOC_367/A 0.10fF
C3228 INVX1_LOC_20/Y INVX1_LOC_666/A 0.01fF
C3229 INVX1_LOC_20/Y NAND2X1_LOC_229/a_36_24# 0.01fF
C3230 INVX1_LOC_625/A INVX1_LOC_224/Y 0.01fF
C3231 NAND2X1_LOC_788/A INVX1_LOC_11/Y 0.02fF
C3232 INVX1_LOC_206/Y INVX1_LOC_504/A 0.09fF
C3233 NAND2X1_LOC_324/B INVX1_LOC_374/A 0.26fF
C3234 INVX1_LOC_442/A INVX1_LOC_80/A 0.09fF
C3235 INVX1_LOC_395/A NAND2X1_LOC_316/a_36_24# 0.00fF
C3236 INPUT_0 INVX1_LOC_17/Y 0.10fF
C3237 INVX1_LOC_547/Y NAND2X1_LOC_496/Y 0.17fF
C3238 INVX1_LOC_45/Y INVX1_LOC_519/A 0.02fF
C3239 NAND2X1_LOC_505/Y INVX1_LOC_600/A 0.03fF
C3240 NAND2X1_LOC_175/a_36_24# INVX1_LOC_566/A 0.00fF
C3241 INVX1_LOC_250/Y INVX1_LOC_51/Y 0.01fF
C3242 INVX1_LOC_45/Y NAND2X1_LOC_296/Y 0.09fF
C3243 INVX1_LOC_160/Y INVX1_LOC_154/Y 0.01fF
C3244 VDD INVX1_LOC_670/A -0.00fF
C3245 INVX1_LOC_323/Y INVX1_LOC_45/Y 0.01fF
C3246 INVX1_LOC_395/A NAND2X1_LOC_708/A 0.03fF
C3247 INVX1_LOC_554/A INVX1_LOC_58/Y 0.02fF
C3248 NAND2X1_LOC_506/a_36_24# INVX1_LOC_586/A 0.00fF
C3249 INVX1_LOC_312/A INVX1_LOC_486/Y 0.00fF
C3250 INVX1_LOC_29/Y INVX1_LOC_334/Y 0.01fF
C3251 INVX1_LOC_586/A INVX1_LOC_252/Y 0.06fF
C3252 INVX1_LOC_11/Y INVX1_LOC_442/A 0.74fF
C3253 INVX1_LOC_602/A INVX1_LOC_53/Y 0.13fF
C3254 NAND2X1_LOC_152/B INVX1_LOC_136/Y 0.06fF
C3255 NAND2X1_LOC_516/B NAND2X1_LOC_413/Y 0.09fF
C3256 INPUT_3 NAND2X1_LOC_296/Y 0.02fF
C3257 INVX1_LOC_587/A INVX1_LOC_656/Y 0.04fF
C3258 INVX1_LOC_118/Y INVX1_LOC_6/Y 0.06fF
C3259 NAND2X1_LOC_16/Y INPUT_1 0.01fF
C3260 INVX1_LOC_20/Y INVX1_LOC_681/A 0.01fF
C3261 INVX1_LOC_400/Y INVX1_LOC_46/Y 0.03fF
C3262 INVX1_LOC_84/A INVX1_LOC_7/Y 0.18fF
C3263 INPUT_0 NAND2X1_LOC_307/B 0.03fF
C3264 INVX1_LOC_428/A INVX1_LOC_93/Y 0.06fF
C3265 INVX1_LOC_459/Y INVX1_LOC_117/Y 0.39fF
C3266 INVX1_LOC_398/A INVX1_LOC_35/Y 0.20fF
C3267 INVX1_LOC_62/A INVX1_LOC_76/Y 0.01fF
C3268 INVX1_LOC_383/A INVX1_LOC_670/A 0.10fF
C3269 INVX1_LOC_21/Y INVX1_LOC_174/A 0.00fF
C3270 INVX1_LOC_510/Y INVX1_LOC_670/A 0.09fF
C3271 INVX1_LOC_139/A INVX1_LOC_496/A 0.02fF
C3272 NAND2X1_LOC_516/Y NAND2X1_LOC_307/B 0.12fF
C3273 INVX1_LOC_80/A INVX1_LOC_116/Y 0.04fF
C3274 INVX1_LOC_251/A INVX1_LOC_134/Y 0.03fF
C3275 INVX1_LOC_522/Y INVX1_LOC_514/A 0.16fF
C3276 INVX1_LOC_402/Y NAND2X1_LOC_413/Y 0.03fF
C3277 INVX1_LOC_17/Y NAND2X1_LOC_123/A 0.00fF
C3278 INVX1_LOC_20/Y NAND2X1_LOC_285/A 0.02fF
C3279 NAND2X1_LOC_704/B INVX1_LOC_66/A 0.05fF
C3280 NAND2X1_LOC_532/Y INVX1_LOC_76/Y 0.01fF
C3281 INVX1_LOC_84/A INVX1_LOC_32/Y 3.75fF
C3282 INVX1_LOC_447/A INVX1_LOC_62/Y 0.03fF
C3283 INVX1_LOC_367/A NAND2X1_LOC_659/a_36_24# 0.00fF
C3284 INVX1_LOC_53/Y INVX1_LOC_117/Y 0.34fF
C3285 INVX1_LOC_551/Y INVX1_LOC_47/Y 0.10fF
C3286 NAND2X1_LOC_697/Y INVX1_LOC_35/Y 0.01fF
C3287 INVX1_LOC_193/Y INVX1_LOC_79/A 0.02fF
C3288 INVX1_LOC_107/A INVX1_LOC_655/A 0.03fF
C3289 INVX1_LOC_451/A INVX1_LOC_35/Y 0.03fF
C3290 INVX1_LOC_254/A INVX1_LOC_600/A 0.04fF
C3291 NAND2X1_LOC_56/Y INVX1_LOC_31/Y 0.01fF
C3292 INVX1_LOC_446/Y INVX1_LOC_502/A 0.04fF
C3293 INVX1_LOC_11/Y INVX1_LOC_116/Y 0.03fF
C3294 INVX1_LOC_523/Y NAND2X1_LOC_820/A 0.02fF
C3295 NAND2X1_LOC_195/a_36_24# INVX1_LOC_176/A 0.02fF
C3296 INVX1_LOC_266/Y INVX1_LOC_245/A 0.13fF
C3297 INVX1_LOC_154/Y NAND2X1_LOC_267/A -0.05fF
C3298 INVX1_LOC_20/Y INVX1_LOC_168/Y 0.07fF
C3299 INVX1_LOC_167/A INVX1_LOC_99/Y 0.01fF
C3300 INVX1_LOC_176/A INVX1_LOC_48/Y 0.08fF
C3301 INVX1_LOC_35/Y INVX1_LOC_665/Y 0.03fF
C3302 INVX1_LOC_210/Y INVX1_LOC_198/A 0.03fF
C3303 INVX1_LOC_80/A INVX1_LOC_255/A 0.07fF
C3304 VDD INVX1_LOC_282/Y 0.21fF
C3305 NAND2X1_LOC_174/a_36_24# INVX1_LOC_156/A 0.00fF
C3306 INVX1_LOC_134/A NAND2X1_LOC_545/A 0.01fF
C3307 INVX1_LOC_32/Y NAND2X1_LOC_67/Y 0.22fF
C3308 INVX1_LOC_522/A INVX1_LOC_137/Y 0.03fF
C3309 NAND2X1_LOC_184/Y NAND2X1_LOC_250/Y 0.05fF
C3310 INVX1_LOC_206/Y INVX1_LOC_346/Y 0.04fF
C3311 INVX1_LOC_6/Y INVX1_LOC_610/A 0.01fF
C3312 INVX1_LOC_277/A NAND2X1_LOC_250/a_36_24# 0.00fF
C3313 NAND2X1_LOC_20/Y INVX1_LOC_9/Y 0.01fF
C3314 INVX1_LOC_117/Y INVX1_LOC_460/Y 0.05fF
C3315 INVX1_LOC_171/Y INVX1_LOC_100/Y 0.05fF
C3316 INVX1_LOC_551/Y INVX1_LOC_119/Y 0.01fF
C3317 INVX1_LOC_607/Y NAND2X1_LOC_307/B 0.05fF
C3318 INVX1_LOC_80/A INVX1_LOC_179/A 0.01fF
C3319 INVX1_LOC_578/A NAND2X1_LOC_458/a_36_24# 0.00fF
C3320 INVX1_LOC_54/Y INVX1_LOC_350/Y 0.00fF
C3321 INVX1_LOC_655/Y INVX1_LOC_100/Y 0.01fF
C3322 INVX1_LOC_662/A NAND2X1_LOC_513/A 0.01fF
C3323 INVX1_LOC_113/Y INVX1_LOC_74/Y 0.01fF
C3324 NAND2X1_LOC_180/B INVX1_LOC_41/Y 0.03fF
C3325 INVX1_LOC_163/Y INVX1_LOC_62/Y 0.01fF
C3326 INVX1_LOC_413/A INVX1_LOC_387/Y 0.01fF
C3327 INVX1_LOC_89/Y NAND2X1_LOC_720/A 0.12fF
C3328 NAND2X1_LOC_333/A NAND2X1_LOC_333/B 0.04fF
C3329 INVX1_LOC_11/Y INVX1_LOC_255/A 0.39fF
C3330 INVX1_LOC_633/Y INVX1_LOC_114/A 0.02fF
C3331 INVX1_LOC_522/A NAND2X1_LOC_829/B 0.18fF
C3332 INVX1_LOC_649/Y INVX1_LOC_100/Y 0.09fF
C3333 NAND2X1_LOC_400/B INVX1_LOC_117/Y 0.17fF
C3334 INVX1_LOC_421/A INVX1_LOC_46/Y 0.05fF
C3335 INVX1_LOC_652/A INVX1_LOC_134/Y 0.02fF
C3336 INVX1_LOC_54/Y NAND2X1_LOC_181/A 0.01fF
C3337 INVX1_LOC_522/Y INVX1_LOC_62/Y 0.07fF
C3338 INVX1_LOC_99/A INVX1_LOC_242/Y 0.03fF
C3339 INVX1_LOC_376/Y INVX1_LOC_98/Y 0.10fF
C3340 INVX1_LOC_384/A NAND2X1_LOC_255/a_36_24# 0.01fF
C3341 INVX1_LOC_581/A NAND2X1_LOC_782/a_36_24# 0.00fF
C3342 INVX1_LOC_170/Y INVX1_LOC_48/Y 0.04fF
C3343 INVX1_LOC_523/Y INVX1_LOC_6/Y 0.07fF
C3344 INVX1_LOC_188/Y INVX1_LOC_41/Y 0.03fF
C3345 NAND2X1_LOC_20/Y INVX1_LOC_13/Y 0.12fF
C3346 INVX1_LOC_603/Y INVX1_LOC_41/Y 0.03fF
C3347 NAND2X1_LOC_184/Y INVX1_LOC_63/Y 0.03fF
C3348 INVX1_LOC_675/A INVX1_LOC_359/Y 0.05fF
C3349 INVX1_LOC_502/A INVX1_LOC_145/Y 0.08fF
C3350 INVX1_LOC_477/Y INVX1_LOC_476/A 0.20fF
C3351 INVX1_LOC_510/Y NAND2X1_LOC_418/a_36_24# 0.00fF
C3352 NAND2X1_LOC_141/a_36_24# INVX1_LOC_47/Y 0.01fF
C3353 NAND2X1_LOC_274/B INVX1_LOC_510/A 0.76fF
C3354 INVX1_LOC_117/Y NAND2X1_LOC_406/B 0.02fF
C3355 INVX1_LOC_62/Y NAND2X1_LOC_646/a_36_24# 0.00fF
C3356 INVX1_LOC_686/A INVX1_LOC_346/Y 0.01fF
C3357 INVX1_LOC_419/A INVX1_LOC_69/Y 0.01fF
C3358 INVX1_LOC_599/A INVX1_LOC_597/Y 0.00fF
C3359 INVX1_LOC_93/Y NAND2X1_LOC_768/B 0.23fF
C3360 INVX1_LOC_69/Y INVX1_LOC_234/Y 0.20fF
C3361 INVX1_LOC_627/A NAND2X1_LOC_797/a_36_24# 0.00fF
C3362 NAND2X1_LOC_187/Y INVX1_LOC_79/A 0.05fF
C3363 INVX1_LOC_176/A NAND2X1_LOC_629/a_36_24# 0.01fF
C3364 INVX1_LOC_277/A INVX1_LOC_100/Y 0.01fF
C3365 INVX1_LOC_199/Y INVX1_LOC_58/Y 0.58fF
C3366 INVX1_LOC_376/A INVX1_LOC_141/Y 0.12fF
C3367 INVX1_LOC_54/Y INVX1_LOC_79/A 4.99fF
C3368 NAND2X1_LOC_507/A INVX1_LOC_100/Y 0.01fF
C3369 INVX1_LOC_17/Y INVX1_LOC_211/A 0.07fF
C3370 INVX1_LOC_646/Y NAND2X1_LOC_847/A 0.21fF
C3371 NAND2X1_LOC_285/A INVX1_LOC_655/A 0.13fF
C3372 INVX1_LOC_411/A INVX1_LOC_62/Y 0.01fF
C3373 INVX1_LOC_31/Y INVX1_LOC_369/Y 0.07fF
C3374 INVX1_LOC_62/Y INVX1_LOC_295/Y 0.03fF
C3375 NAND2X1_LOC_387/Y INVX1_LOC_41/Y 0.07fF
C3376 INVX1_LOC_58/Y INVX1_LOC_499/A 0.02fF
C3377 INVX1_LOC_89/Y INVX1_LOC_100/Y 1.10fF
C3378 INVX1_LOC_49/Y INVX1_LOC_373/Y 0.02fF
C3379 INVX1_LOC_50/Y INVX1_LOC_666/Y 0.03fF
C3380 INVX1_LOC_133/Y INVX1_LOC_554/Y 0.01fF
C3381 INVX1_LOC_183/A INVX1_LOC_26/Y 0.11fF
C3382 INVX1_LOC_89/Y INVX1_LOC_74/Y 3.30fF
C3383 INVX1_LOC_224/A INVX1_LOC_245/A 0.00fF
C3384 NAND2X1_LOC_843/B INVX1_LOC_66/A 0.59fF
C3385 VDD INVX1_LOC_616/Y 0.14fF
C3386 INVX1_LOC_31/Y INVX1_LOC_223/A 0.20fF
C3387 INVX1_LOC_100/A NAND2X1_LOC_263/a_36_24# 0.00fF
C3388 INVX1_LOC_31/Y INVX1_LOC_348/Y 0.42fF
C3389 NAND2X1_LOC_274/B NAND2X1_LOC_477/a_36_24# 0.00fF
C3390 INVX1_LOC_63/Y INVX1_LOC_75/Y 0.13fF
C3391 INVX1_LOC_206/Y NAND2X1_LOC_76/B 0.07fF
C3392 INVX1_LOC_501/A INVX1_LOC_74/Y 0.03fF
C3393 INVX1_LOC_479/A INVX1_LOC_356/Y 0.06fF
C3394 INPUT_0 NAND2X1_LOC_88/Y 0.10fF
C3395 NAND2X1_LOC_845/B INVX1_LOC_41/Y 0.01fF
C3396 INVX1_LOC_562/A NAND2X1_LOC_719/a_36_24# 0.02fF
C3397 INPUT_6 INVX1_LOC_34/Y 0.01fF
C3398 NAND2X1_LOC_271/B NAND2X1_LOC_457/A 0.02fF
C3399 NAND2X1_LOC_317/B NAND2X1_LOC_314/a_36_24# 0.00fF
C3400 NAND2X1_LOC_120/a_36_24# INVX1_LOC_638/A 0.01fF
C3401 INVX1_LOC_95/A NAND2X1_LOC_98/B 0.14fF
C3402 INVX1_LOC_100/Y NAND2X1_LOC_544/B 0.06fF
C3403 INVX1_LOC_224/Y INVX1_LOC_65/Y 0.07fF
C3404 NAND2X1_LOC_797/a_36_24# INVX1_LOC_581/A 0.00fF
C3405 VDD NAND2X1_LOC_516/B 0.03fF
C3406 INVX1_LOC_41/Y INVX1_LOC_91/A 0.01fF
C3407 NAND2X1_LOC_786/B NAND2X1_LOC_201/a_36_24# 0.00fF
C3408 INVX1_LOC_185/A INVX1_LOC_53/Y 0.03fF
C3409 INVX1_LOC_74/Y NAND2X1_LOC_544/B 0.33fF
C3410 INVX1_LOC_578/A INVX1_LOC_65/Y 0.02fF
C3411 NAND2X1_LOC_475/A INVX1_LOC_551/Y 0.10fF
C3412 NAND2X1_LOC_537/A INVX1_LOC_600/A 0.03fF
C3413 INVX1_LOC_301/A INVX1_LOC_99/A 0.02fF
C3414 NAND2X1_LOC_373/Y NAND2X1_LOC_325/B 0.01fF
C3415 NAND2X1_LOC_475/A NAND2X1_LOC_304/a_36_24# -0.02fF
C3416 VDD INVX1_LOC_639/Y 0.35fF
C3417 INVX1_LOC_402/Y VDD 0.35fF
C3418 INVX1_LOC_206/Y INVX1_LOC_530/A 0.02fF
C3419 INVX1_LOC_366/A NAND2X1_LOC_460/a_36_24# 0.02fF
C3420 INVX1_LOC_287/A INVX1_LOC_224/Y 0.01fF
C3421 NAND2X1_LOC_613/Y INVX1_LOC_482/A 0.13fF
C3422 NAND2X1_LOC_39/Y INVX1_LOC_45/Y 0.10fF
C3423 INVX1_LOC_193/Y INVX1_LOC_417/Y 0.00fF
C3424 INVX1_LOC_625/A INVX1_LOC_206/Y 0.02fF
C3425 NAND2X1_LOC_45/Y INVX1_LOC_211/Y 0.05fF
C3426 INVX1_LOC_257/Y INVX1_LOC_17/Y 0.10fF
C3427 INVX1_LOC_238/Y INVX1_LOC_35/Y 0.00fF
C3428 INVX1_LOC_626/Y INVX1_LOC_137/Y 0.15fF
C3429 NAND2X1_LOC_795/a_36_24# INVX1_LOC_395/A 0.00fF
C3430 NAND2X1_LOC_243/A INVX1_LOC_616/Y 0.01fF
C3431 NAND2X1_LOC_788/A INVX1_LOC_374/Y 0.01fF
C3432 INVX1_LOC_393/Y INVX1_LOC_159/A 0.01fF
C3433 INVX1_LOC_418/A INVX1_LOC_99/Y 0.00fF
C3434 INVX1_LOC_400/Y INVX1_LOC_202/Y 0.04fF
C3435 VDD INVX1_LOC_267/A -0.00fF
C3436 NAND2X1_LOC_791/B NAND2X1_LOC_757/a_36_24# 0.02fF
C3437 INVX1_LOC_33/A INVX1_LOC_25/Y 0.12fF
C3438 INPUT_0 INVX1_LOC_198/A 0.05fF
C3439 INVX1_LOC_17/Y INVX1_LOC_288/A 0.14fF
C3440 INVX1_LOC_174/Y INVX1_LOC_7/Y 0.00fF
C3441 INVX1_LOC_254/Y INVX1_LOC_412/A 0.01fF
C3442 INVX1_LOC_435/Y INVX1_LOC_282/A 0.02fF
C3443 NAND2X1_LOC_507/a_36_24# INVX1_LOC_35/Y 0.00fF
C3444 INVX1_LOC_364/Y INVX1_LOC_35/Y 0.03fF
C3445 INVX1_LOC_384/A INVX1_LOC_503/A 0.03fF
C3446 INVX1_LOC_412/Y INVX1_LOC_372/A 0.02fF
C3447 INVX1_LOC_293/Y NAND2X1_LOC_363/a_36_24# 0.00fF
C3448 INVX1_LOC_294/Y INVX1_LOC_297/A 0.07fF
C3449 INVX1_LOC_677/Y INVX1_LOC_602/Y 0.00fF
C3450 INVX1_LOC_51/A INVX1_LOC_93/Y 0.02fF
C3451 VDD NAND2X1_LOC_520/A 0.00fF
C3452 VDD INVX1_LOC_331/Y 0.21fF
C3453 INVX1_LOC_17/Y INVX1_LOC_384/A 0.07fF
C3454 NAND2X1_LOC_685/A INVX1_LOC_358/Y 0.01fF
C3455 INVX1_LOC_268/A INVX1_LOC_566/Y 0.15fF
C3456 INVX1_LOC_581/A NAND2X1_LOC_738/a_36_24# 0.02fF
C3457 INVX1_LOC_45/Y INVX1_LOC_513/A 0.00fF
C3458 INVX1_LOC_62/Y NAND2X1_LOC_216/a_36_24# 0.01fF
C3459 NAND2X1_LOC_498/Y INVX1_LOC_46/Y 0.07fF
C3460 NAND2X1_LOC_833/B INVX1_LOC_220/A 0.27fF
C3461 NAND2X1_LOC_321/a_36_24# INVX1_LOC_633/Y 0.00fF
C3462 INVX1_LOC_570/A INVX1_LOC_46/Y 0.03fF
C3463 INVX1_LOC_20/Y INVX1_LOC_137/Y 0.23fF
C3464 INVX1_LOC_367/A NAND2X1_LOC_413/Y 0.01fF
C3465 INVX1_LOC_21/Y INVX1_LOC_324/Y 0.06fF
C3466 INVX1_LOC_206/Y NAND2X1_LOC_52/Y 0.03fF
C3467 INVX1_LOC_315/Y NAND2X1_LOC_387/Y 0.10fF
C3468 INVX1_LOC_53/Y INVX1_LOC_281/Y 0.14fF
C3469 INVX1_LOC_155/A INVX1_LOC_271/A 0.03fF
C3470 INVX1_LOC_584/A INVX1_LOC_49/Y 0.08fF
C3471 INVX1_LOC_395/A NAND2X1_LOC_284/A 0.05fF
C3472 INVX1_LOC_21/Y INVX1_LOC_603/Y 0.53fF
C3473 INVX1_LOC_54/Y INVX1_LOC_610/Y 0.01fF
C3474 NAND2X1_LOC_331/A INVX1_LOC_507/Y 0.01fF
C3475 INVX1_LOC_206/Y NAND2X1_LOC_686/A 0.02fF
C3476 INVX1_LOC_400/Y INVX1_LOC_49/Y 0.07fF
C3477 NAND2X1_LOC_379/Y INVX1_LOC_35/Y 0.06fF
C3478 INVX1_LOC_552/Y INVX1_LOC_551/A 0.06fF
C3479 INVX1_LOC_53/Y INVX1_LOC_251/Y 0.07fF
C3480 INVX1_LOC_448/A INVX1_LOC_503/A 0.13fF
C3481 INVX1_LOC_35/Y INVX1_LOC_134/Y 0.08fF
C3482 INVX1_LOC_304/A INVX1_LOC_134/Y 0.00fF
C3483 INVX1_LOC_21/Y INVX1_LOC_43/Y 0.01fF
C3484 INVX1_LOC_378/A INVX1_LOC_490/A 0.01fF
C3485 INVX1_LOC_254/Y NAND2X1_LOC_336/B 0.21fF
C3486 INVX1_LOC_419/A INVX1_LOC_586/A 0.01fF
C3487 INVX1_LOC_446/A INVX1_LOC_75/Y 0.04fF
C3488 NAND2X1_LOC_755/B INVX1_LOC_99/Y 0.03fF
C3489 INVX1_LOC_607/A INVX1_LOC_63/Y 0.01fF
C3490 INVX1_LOC_47/A INVX1_LOC_35/Y 0.01fF
C3491 INVX1_LOC_341/Y INVX1_LOC_59/A 0.12fF
C3492 INVX1_LOC_206/Y INVX1_LOC_519/Y 0.11fF
C3493 NAND2X1_LOC_670/a_36_24# INVX1_LOC_600/A 0.00fF
C3494 NAND2X1_LOC_390/a_36_24# INVX1_LOC_199/Y 0.01fF
C3495 INVX1_LOC_17/Y INVX1_LOC_145/Y 0.35fF
C3496 INVX1_LOC_566/A INVX1_LOC_89/Y 0.07fF
C3497 INVX1_LOC_201/Y INVX1_LOC_274/A 0.35fF
C3498 INVX1_LOC_80/A NAND2X1_LOC_148/B 0.56fF
C3499 INVX1_LOC_126/A INVX1_LOC_6/Y 0.03fF
C3500 NAND2X1_LOC_184/Y INVX1_LOC_387/A 0.03fF
C3501 NAND2X1_LOC_41/Y INVX1_LOC_35/Y 0.02fF
C3502 INVX1_LOC_417/Y INVX1_LOC_54/Y 0.03fF
C3503 NAND2X1_LOC_173/Y INVX1_LOC_675/A 0.01fF
C3504 INVX1_LOC_322/Y INVX1_LOC_9/Y 0.08fF
C3505 INVX1_LOC_413/Y INVX1_LOC_26/Y 0.21fF
C3506 INVX1_LOC_203/Y INVX1_LOC_74/Y 0.00fF
C3507 INVX1_LOC_603/Y NAND2X1_LOC_267/A 0.01fF
C3508 INVX1_LOC_21/Y NAND2X1_LOC_387/Y 0.07fF
C3509 INVX1_LOC_540/Y INVX1_LOC_62/Y 0.11fF
C3510 NAND2X1_LOC_521/a_36_24# INVX1_LOC_392/A 0.00fF
C3511 INVX1_LOC_24/A INVX1_LOC_653/Y 0.04fF
C3512 VDD NAND2X1_LOC_227/A -0.00fF
C3513 INVX1_LOC_566/A INVX1_LOC_501/A 0.07fF
C3514 INVX1_LOC_54/Y INVX1_LOC_59/Y 0.03fF
C3515 INVX1_LOC_80/A INVX1_LOC_69/Y 0.56fF
C3516 INVX1_LOC_446/A NAND2X1_LOC_271/A 0.02fF
C3517 INVX1_LOC_99/Y INVX1_LOC_46/Y 10.41fF
C3518 NAND2X1_LOC_165/Y INVX1_LOC_35/Y 0.02fF
C3519 INVX1_LOC_579/Y INVX1_LOC_69/Y 0.12fF
C3520 INVX1_LOC_51/Y INVX1_LOC_369/Y 0.07fF
C3521 INVX1_LOC_588/Y INVX1_LOC_259/Y 0.03fF
C3522 INVX1_LOC_276/A INVX1_LOC_106/Y 0.01fF
C3523 INVX1_LOC_53/Y INVX1_LOC_58/Y 0.17fF
C3524 NAND2X1_LOC_187/a_36_24# INVX1_LOC_99/Y 0.00fF
C3525 NAND2X1_LOC_187/Y INVX1_LOC_48/Y 0.18fF
C3526 INVX1_LOC_412/A INVX1_LOC_479/A 0.08fF
C3527 INVX1_LOC_145/Y INVX1_LOC_601/Y 0.02fF
C3528 INVX1_LOC_53/A INVX1_LOC_18/Y 0.03fF
C3529 INVX1_LOC_54/Y INVX1_LOC_48/Y 0.21fF
C3530 INVX1_LOC_617/Y NAND2X1_LOC_274/B -0.00fF
C3531 INVX1_LOC_569/A INVX1_LOC_655/A 0.02fF
C3532 NAND2X1_LOC_376/B INVX1_LOC_7/Y 0.03fF
C3533 INVX1_LOC_105/A INVX1_LOC_670/A 0.32fF
C3534 INVX1_LOC_12/Y INVX1_LOC_482/Y 0.03fF
C3535 INVX1_LOC_32/Y INVX1_LOC_156/A 0.13fF
C3536 INVX1_LOC_211/Y INVX1_LOC_47/Y 0.31fF
C3537 NAND2X1_LOC_307/A INVX1_LOC_242/Y 0.02fF
C3538 INVX1_LOC_49/Y INVX1_LOC_537/A 0.09fF
C3539 INVX1_LOC_498/A INVX1_LOC_497/Y 0.03fF
C3540 INVX1_LOC_431/A INVX1_LOC_431/Y 0.02fF
C3541 NAND2X1_LOC_347/a_36_24# INVX1_LOC_50/Y 0.00fF
C3542 NAND2X1_LOC_707/A INVX1_LOC_479/A 1.83fF
C3543 INVX1_LOC_127/Y INVX1_LOC_361/Y 0.03fF
C3544 INVX1_LOC_50/Y INVX1_LOC_18/Y 0.01fF
C3545 INVX1_LOC_11/Y INVX1_LOC_69/Y 0.52fF
C3546 NAND2X1_LOC_299/Y NAND2X1_LOC_299/a_36_24# 0.00fF
C3547 INVX1_LOC_573/Y INVX1_LOC_330/A 0.01fF
C3548 NAND2X1_LOC_292/Y INVX1_LOC_48/Y 0.17fF
C3549 INVX1_LOC_442/A INVX1_LOC_625/Y 0.07fF
C3550 INVX1_LOC_586/A NAND2X1_LOC_231/B 0.07fF
C3551 INVX1_LOC_51/Y INVX1_LOC_348/Y 0.03fF
C3552 INVX1_LOC_53/Y NAND2X1_LOC_342/B 0.08fF
C3553 INVX1_LOC_198/A NAND2X1_LOC_215/a_36_24# 0.00fF
C3554 NAND2X1_LOC_301/a_36_24# INVX1_LOC_154/A 0.00fF
C3555 INVX1_LOC_47/Y INVX1_LOC_46/Y 0.18fF
C3556 NAND2X1_LOC_698/Y INVX1_LOC_117/Y 0.08fF
C3557 INVX1_LOC_44/Y NAND2X1_LOC_720/A 1.10fF
C3558 NAND2X1_LOC_557/B INVX1_LOC_46/Y 0.03fF
C3559 INVX1_LOC_656/A INVX1_LOC_659/A 0.03fF
C3560 INVX1_LOC_421/A INVX1_LOC_49/Y 0.03fF
C3561 NAND2X1_LOC_336/B INVX1_LOC_479/A 0.03fF
C3562 INVX1_LOC_6/Y NAND2X1_LOC_814/Y 0.01fF
C3563 INVX1_LOC_62/Y NAND2X1_LOC_658/a_36_24# 0.01fF
C3564 INVX1_LOC_62/Y NAND2X1_LOC_496/Y 0.10fF
C3565 NAND2X1_LOC_513/A INVX1_LOC_653/Y 0.01fF
C3566 INVX1_LOC_92/A INVX1_LOC_624/A 0.02fF
C3567 INVX1_LOC_419/Y INVX1_LOC_242/Y 0.20fF
C3568 INVX1_LOC_469/Y INVX1_LOC_501/A 0.03fF
C3569 INVX1_LOC_117/Y INVX1_LOC_662/A 0.14fF
C3570 INVX1_LOC_520/Y GATE_662 0.09fF
C3571 INVX1_LOC_41/Y INVX1_LOC_504/Y 0.07fF
C3572 INVX1_LOC_100/Y INVX1_LOC_194/Y 3.13fF
C3573 INVX1_LOC_588/Y INVX1_LOC_114/A 0.12fF
C3574 NAND2X1_LOC_324/a_36_24# INVX1_LOC_62/Y 0.01fF
C3575 NAND2X1_LOC_775/B INVX1_LOC_62/Y 0.03fF
C3576 INVX1_LOC_166/A INVX1_LOC_114/A 0.02fF
C3577 INVX1_LOC_119/Y INVX1_LOC_46/Y 0.03fF
C3578 NAND2X1_LOC_66/Y INVX1_LOC_46/Y 0.03fF
C3579 INVX1_LOC_199/Y INVX1_LOC_245/A 0.08fF
C3580 NAND2X1_LOC_433/Y INVX1_LOC_69/Y 0.46fF
C3581 INVX1_LOC_116/Y INVX1_LOC_625/Y 0.03fF
C3582 NAND2X1_LOC_325/a_36_24# INVX1_LOC_242/Y 0.01fF
C3583 INVX1_LOC_89/Y INVX1_LOC_79/A 0.46fF
C3584 INVX1_LOC_388/A INVX1_LOC_48/Y 0.01fF
C3585 INVX1_LOC_327/A INVX1_LOC_327/Y 0.02fF
C3586 INVX1_LOC_93/Y INVX1_LOC_441/A 0.02fF
C3587 INVX1_LOC_93/Y INVX1_LOC_354/A 0.00fF
C3588 GATE_479 INVX1_LOC_244/Y 0.00fF
C3589 INVX1_LOC_501/A INVX1_LOC_79/A 0.07fF
C3590 NAND2X1_LOC_349/a_36_24# INVX1_LOC_655/A 0.01fF
C3591 NAND2X1_LOC_503/B INPUT_0 0.01fF
C3592 NAND2X1_LOC_475/A INVX1_LOC_596/Y 0.00fF
C3593 INVX1_LOC_31/Y NAND2X1_LOC_832/A 0.23fF
C3594 INVX1_LOC_65/Y NAND2X1_LOC_86/Y 0.01fF
C3595 INVX1_LOC_675/A INVX1_LOC_354/A 0.02fF
C3596 INVX1_LOC_255/A INVX1_LOC_625/Y 0.07fF
C3597 NAND2X1_LOC_292/a_36_24# INVX1_LOC_280/A 0.00fF
C3598 VDD INVX1_LOC_546/Y 0.21fF
C3599 NAND2X1_LOC_164/Y INVX1_LOC_206/Y 0.08fF
C3600 INVX1_LOC_438/A INVX1_LOC_490/Y 0.00fF
C3601 NAND2X1_LOC_750/Y INVX1_LOC_395/A 0.10fF
C3602 VDD INVX1_LOC_392/Y 0.32fF
C3603 NAND2X1_LOC_241/B INVX1_LOC_395/A 0.15fF
C3604 INVX1_LOC_606/Y INVX1_LOC_395/A 0.05fF
C3605 NAND2X1_LOC_45/Y INVX1_LOC_530/Y 0.00fF
C3606 INVX1_LOC_206/Y INVX1_LOC_65/Y 1.75fF
C3607 INVX1_LOC_74/Y INVX1_LOC_347/A 0.17fF
C3608 NAND2X1_LOC_741/a_36_24# NAND2X1_LOC_122/Y 0.00fF
C3609 INVX1_LOC_3/Y INVX1_LOC_334/Y 0.01fF
C3610 VDD INVX1_LOC_524/Y 0.21fF
C3611 INPUT_0 INVX1_LOC_273/A 0.40fF
C3612 NAND2X1_LOC_475/A INVX1_LOC_287/Y 0.00fF
C3613 INVX1_LOC_301/A NAND2X1_LOC_307/A 0.07fF
C3614 INVX1_LOC_301/A INVX1_LOC_545/Y 0.04fF
C3615 NAND2X1_LOC_164/Y INVX1_LOC_396/Y 0.10fF
C3616 NAND2X1_LOC_475/A INVX1_LOC_270/A 0.16fF
C3617 NAND2X1_LOC_331/A INVX1_LOC_163/Y 0.01fF
C3618 NAND2X1_LOC_537/A NAND2X1_LOC_56/Y 0.18fF
C3619 NAND2X1_LOC_637/A INVX1_LOC_579/Y 0.08fF
C3620 INVX1_LOC_400/Y INVX1_LOC_76/Y 0.07fF
C3621 INVX1_LOC_619/A INVX1_LOC_616/Y 0.02fF
C3622 NAND2X1_LOC_331/A INVX1_LOC_522/Y 0.05fF
C3623 INVX1_LOC_85/Y INVX1_LOC_366/A 0.41fF
C3624 VDD INVX1_LOC_516/A 0.04fF
C3625 NAND2X1_LOC_208/a_36_24# INVX1_LOC_85/Y 0.00fF
C3626 VDD INVX1_LOC_669/Y 0.32fF
C3627 INPUT_6 INVX1_LOC_57/Y 0.01fF
C3628 INVX1_LOC_32/A INVX1_LOC_99/Y 0.01fF
C3629 INVX1_LOC_416/A INVX1_LOC_301/A 0.21fF
C3630 INVX1_LOC_419/Y INVX1_LOC_301/A 0.01fF
C3631 INVX1_LOC_150/Y INVX1_LOC_511/A 0.01fF
C3632 VDD INVX1_LOC_392/A 0.00fF
C3633 INVX1_LOC_412/A INVX1_LOC_12/Y 0.01fF
C3634 INVX1_LOC_434/A INVX1_LOC_451/A 0.20fF
C3635 INVX1_LOC_255/Y INVX1_LOC_188/Y 0.03fF
C3636 INVX1_LOC_11/Y INVX1_LOC_217/A 0.09fF
C3637 INVX1_LOC_211/Y NAND2X1_LOC_475/A 0.01fF
C3638 INVX1_LOC_449/A INVX1_LOC_393/A 0.03fF
C3639 INVX1_LOC_421/Y INVX1_LOC_442/Y 0.04fF
C3640 INVX1_LOC_30/Y INVX1_LOC_29/A 0.20fF
C3641 INVX1_LOC_84/A NAND2X1_LOC_384/a_36_24# 0.01fF
C3642 INVX1_LOC_80/A INVX1_LOC_586/A 0.18fF
C3643 INVX1_LOC_249/Y NAND2X1_LOC_123/A 0.03fF
C3644 INVX1_LOC_206/Y INVX1_LOC_479/Y 0.00fF
C3645 INVX1_LOC_21/Y INVX1_LOC_269/A 0.07fF
C3646 INVX1_LOC_400/A INVX1_LOC_228/Y 1.08fF
C3647 INVX1_LOC_51/Y INVX1_LOC_558/Y 0.09fF
C3648 VDD INVX1_LOC_93/Y 3.35fF
C3649 INVX1_LOC_312/A INVX1_LOC_381/A 0.06fF
C3650 INVX1_LOC_625/A INVX1_LOC_397/A 0.02fF
C3651 NAND2X1_LOC_122/Y NAND2X1_LOC_123/A 0.03fF
C3652 NAND2X1_LOC_486/B INVX1_LOC_387/A 0.36fF
C3653 INVX1_LOC_599/Y INVX1_LOC_366/A 0.01fF
C3654 INVX1_LOC_20/Y NAND2X1_LOC_307/A 0.01fF
C3655 NAND2X1_LOC_475/A INVX1_LOC_46/Y 0.03fF
C3656 INVX1_LOC_295/A INVX1_LOC_596/A 0.20fF
C3657 INVX1_LOC_35/Y NAND2X1_LOC_249/a_36_24# 0.00fF
C3658 NAND2X1_LOC_750/Y INVX1_LOC_31/Y 0.00fF
C3659 INVX1_LOC_206/Y INVX1_LOC_318/A 0.02fF
C3660 INVX1_LOC_299/A INVX1_LOC_673/Y 0.05fF
C3661 NAND2X1_LOC_45/Y INVX1_LOC_387/Y 0.03fF
C3662 NAND2X1_LOC_677/Y INVX1_LOC_610/Y 0.01fF
C3663 INVX1_LOC_602/A INPUT_7 0.02fF
C3664 INVX1_LOC_166/A NAND2X1_LOC_314/a_36_24# 0.00fF
C3665 INVX1_LOC_201/A INVX1_LOC_273/A 0.02fF
C3666 INVX1_LOC_312/Y INVX1_LOC_80/A 0.03fF
C3667 INVX1_LOC_362/Y INVX1_LOC_371/A 0.03fF
C3668 INVX1_LOC_420/Y INVX1_LOC_31/Y 0.01fF
C3669 NAND2X1_LOC_521/a_36_24# INVX1_LOC_362/Y 0.00fF
C3670 INVX1_LOC_32/A INVX1_LOC_47/Y 0.07fF
C3671 NAND2X1_LOC_318/A INVX1_LOC_99/Y 0.03fF
C3672 INVX1_LOC_206/Y INVX1_LOC_397/Y 0.04fF
C3673 VDD INVX1_LOC_675/A 1.02fF
C3674 INVX1_LOC_272/Y INVX1_LOC_599/Y 0.27fF
C3675 INVX1_LOC_11/Y INVX1_LOC_586/A 10.28fF
C3676 INVX1_LOC_442/A INVX1_LOC_361/Y 0.03fF
C3677 NAND2X1_LOC_336/B INVX1_LOC_12/Y 0.00fF
C3678 NAND2X1_LOC_840/a_36_24# NAND2X1_LOC_260/Y 0.00fF
C3679 NAND2X1_LOC_45/Y INVX1_LOC_49/Y 0.17fF
C3680 INVX1_LOC_21/Y NAND2X1_LOC_24/Y 0.03fF
C3681 INVX1_LOC_380/A INVX1_LOC_62/Y 0.01fF
C3682 INVX1_LOC_269/A NAND2X1_LOC_267/A 0.44fF
C3683 INVX1_LOC_20/Y INVX1_LOC_416/A 0.03fF
C3684 INVX1_LOC_224/Y INVX1_LOC_63/Y 0.07fF
C3685 VDD NAND2X1_LOC_334/B 0.27fF
C3686 INVX1_LOC_383/A INVX1_LOC_93/Y 0.08fF
C3687 INVX1_LOC_578/A INVX1_LOC_253/Y 0.01fF
C3688 NAND2X1_LOC_242/A INVX1_LOC_44/Y 0.09fF
C3689 INVX1_LOC_206/Y INVX1_LOC_95/A 0.01fF
C3690 INVX1_LOC_564/A INVX1_LOC_69/Y 0.00fF
C3691 INVX1_LOC_409/Y NAND2X1_LOC_301/B 0.03fF
C3692 VDD INVX1_LOC_643/Y 0.21fF
C3693 INVX1_LOC_25/Y INVX1_LOC_333/A 0.01fF
C3694 INVX1_LOC_300/A NAND2X1_LOC_307/A 0.00fF
C3695 INVX1_LOC_304/Y INVX1_LOC_235/Y 0.00fF
C3696 INVX1_LOC_93/Y INVX1_LOC_510/Y 0.06fF
C3697 VDD INVX1_LOC_543/A -0.00fF
C3698 INVX1_LOC_206/Y INVX1_LOC_314/Y 0.03fF
C3699 INVX1_LOC_119/A INVX1_LOC_159/Y 0.00fF
C3700 INVX1_LOC_683/Y INVX1_LOC_371/A 0.41fF
C3701 NAND2X1_LOC_677/Y NAND2X1_LOC_679/B 0.17fF
C3702 INVX1_LOC_53/Y INVX1_LOC_1/Y 0.27fF
C3703 INVX1_LOC_578/A INVX1_LOC_63/Y 0.07fF
C3704 NAND2X1_LOC_498/Y INVX1_LOC_49/Y 3.08fF
C3705 NAND2X1_LOC_616/Y INVX1_LOC_145/Y 0.06fF
C3706 INVX1_LOC_530/Y INVX1_LOC_47/Y 0.10fF
C3707 INVX1_LOC_85/Y INVX1_LOC_6/Y 0.03fF
C3708 INVX1_LOC_11/Y INVX1_LOC_312/Y 0.11fF
C3709 NAND2X1_LOC_176/Y INVX1_LOC_100/Y 0.03fF
C3710 INVX1_LOC_51/Y INVX1_LOC_187/Y 0.14fF
C3711 INVX1_LOC_570/A INVX1_LOC_49/Y 0.08fF
C3712 INVX1_LOC_557/A INVX1_LOC_63/Y 0.14fF
C3713 INVX1_LOC_17/Y NAND2X1_LOC_260/Y 0.03fF
C3714 INVX1_LOC_32/A NAND2X1_LOC_66/Y 0.01fF
C3715 INPUT_4 INVX1_LOC_60/Y 0.01fF
C3716 INVX1_LOC_377/A INVX1_LOC_510/A 0.02fF
C3717 NAND2X1_LOC_804/a_36_24# INPUT_1 0.01fF
C3718 NAND2X1_LOC_503/B INVX1_LOC_211/A 0.17fF
C3719 INVX1_LOC_132/Y NAND2X1_LOC_342/A 0.01fF
C3720 INVX1_LOC_410/Y NAND2X1_LOC_274/B 0.00fF
C3721 NAND2X1_LOC_318/A INVX1_LOC_47/Y 0.00fF
C3722 INVX1_LOC_118/Y INVX1_LOC_100/Y 0.03fF
C3723 NAND2X1_LOC_148/B INVX1_LOC_131/A 0.01fF
C3724 INVX1_LOC_293/A INVX1_LOC_651/Y 0.02fF
C3725 INVX1_LOC_139/A INVX1_LOC_373/Y 0.00fF
C3726 INVX1_LOC_503/A INVX1_LOC_503/Y 0.06fF
C3727 NAND2X1_LOC_595/Y INVX1_LOC_510/A 0.02fF
C3728 INVX1_LOC_468/Y INVX1_LOC_506/Y 0.38fF
C3729 INVX1_LOC_20/Y NAND2X1_LOC_342/A 0.26fF
C3730 INVX1_LOC_375/A NAND2X1_LOC_274/B 1.70fF
C3731 INVX1_LOC_442/Y INVX1_LOC_159/A 0.00fF
C3732 NAND2X1_LOC_176/Y INVX1_LOC_74/Y 0.06fF
C3733 INVX1_LOC_546/A NAND2X1_LOC_274/B 0.02fF
C3734 INVX1_LOC_136/Y INVX1_LOC_46/Y 0.01fF
C3735 INVX1_LOC_402/A INVX1_LOC_117/Y 0.03fF
C3736 INVX1_LOC_20/Y INVX1_LOC_376/A 0.08fF
C3737 INVX1_LOC_377/Y INVX1_LOC_49/Y 0.04fF
C3738 NAND2X1_LOC_543/B INVX1_LOC_634/Y 0.01fF
C3739 INVX1_LOC_208/A NAND2X1_LOC_241/a_36_24# 0.00fF
C3740 INVX1_LOC_145/Y INVX1_LOC_198/A 0.00fF
C3741 INVX1_LOC_352/Y INVX1_LOC_440/Y 0.31fF
C3742 NAND2X1_LOC_475/A INVX1_LOC_75/A 0.04fF
C3743 INVX1_LOC_405/A NAND2X1_LOC_271/A 0.01fF
C3744 NAND2X1_LOC_519/a_36_24# INVX1_LOC_502/A 0.01fF
C3745 INVX1_LOC_361/Y INVX1_LOC_116/Y 0.07fF
C3746 INVX1_LOC_206/Y INVX1_LOC_588/A 0.05fF
C3747 NAND2X1_LOC_368/a_36_24# INVX1_LOC_75/Y 0.01fF
C3748 INVX1_LOC_169/A INVX1_LOC_9/Y 0.03fF
C3749 INVX1_LOC_609/A INVX1_LOC_550/A 0.08fF
C3750 NAND2X1_LOC_541/B INVX1_LOC_420/A 0.02fF
C3751 INVX1_LOC_599/Y INVX1_LOC_6/Y 0.01fF
C3752 INVX1_LOC_93/Y INVX1_LOC_116/A 0.06fF
C3753 INVX1_LOC_89/Y INVX1_LOC_509/Y 0.01fF
C3754 INVX1_LOC_145/Y INVX1_LOC_230/Y 0.12fF
C3755 INVX1_LOC_417/Y INVX1_LOC_89/Y 0.05fF
C3756 INVX1_LOC_197/A INVX1_LOC_347/Y 0.03fF
C3757 INVX1_LOC_387/Y INVX1_LOC_99/Y 0.02fF
C3758 INVX1_LOC_395/A INVX1_LOC_645/Y 0.17fF
C3759 NAND2X1_LOC_148/A INVX1_LOC_58/Y 0.01fF
C3760 INVX1_LOC_542/A INVX1_LOC_41/Y 0.01fF
C3761 INVX1_LOC_93/Y INVX1_LOC_509/A 0.20fF
C3762 INVX1_LOC_442/Y INVX1_LOC_66/A 0.07fF
C3763 NAND2X1_LOC_107/Y INVX1_LOC_58/Y 0.13fF
C3764 INVX1_LOC_337/Y INVX1_LOC_9/Y 0.02fF
C3765 INVX1_LOC_406/Y NAND2X1_LOC_274/B 0.00fF
C3766 INVX1_LOC_58/Y INVX1_LOC_69/A 0.12fF
C3767 INVX1_LOC_89/Y INVX1_LOC_59/Y 0.03fF
C3768 INVX1_LOC_682/A INVX1_LOC_519/A 0.00fF
C3769 INVX1_LOC_6/A INVX1_LOC_6/Y 0.00fF
C3770 INVX1_LOC_69/Y INVX1_LOC_367/Y 0.03fF
C3771 INVX1_LOC_53/Y INVX1_LOC_245/A 0.06fF
C3772 INVX1_LOC_137/Y INVX1_LOC_627/Y 0.01fF
C3773 INVX1_LOC_49/Y INVX1_LOC_99/Y 4.49fF
C3774 NAND2X1_LOC_613/Y INVX1_LOC_62/Y 0.19fF
C3775 INVX1_LOC_35/Y INVX1_LOC_476/A 0.01fF
C3776 INVX1_LOC_93/Y INVX1_LOC_103/Y 0.03fF
C3777 INVX1_LOC_364/Y INVX1_LOC_364/A 0.04fF
C3778 INVX1_LOC_468/Y INVX1_LOC_63/Y 0.10fF
C3779 NAND2X1_LOC_426/Y INVX1_LOC_505/Y 0.04fF
C3780 INVX1_LOC_100/A INVX1_LOC_50/Y 0.04fF
C3781 INVX1_LOC_62/Y INVX1_LOC_169/A 0.06fF
C3782 INVX1_LOC_89/Y INVX1_LOC_48/Y 0.38fF
C3783 INVX1_LOC_617/Y INVX1_LOC_468/A 0.05fF
C3784 INVX1_LOC_188/Y INVX1_LOC_26/Y 12.11fF
C3785 INVX1_LOC_273/A INVX1_LOC_211/A 0.07fF
C3786 INVX1_LOC_154/A INVX1_LOC_48/Y 0.00fF
C3787 INVX1_LOC_603/Y INVX1_LOC_26/Y 0.00fF
C3788 INVX1_LOC_213/Y INVX1_LOC_58/Y 0.05fF
C3789 INVX1_LOC_635/Y INVX1_LOC_59/A 0.00fF
C3790 INVX1_LOC_80/A NAND2X1_LOC_248/a_36_24# 0.00fF
C3791 INVX1_LOC_145/Y INVX1_LOC_35/A 0.01fF
C3792 INVX1_LOC_43/Y INVX1_LOC_26/Y 0.00fF
C3793 INVX1_LOC_35/Y INVX1_LOC_351/A 0.01fF
C3794 INVX1_LOC_361/Y INVX1_LOC_255/A 0.03fF
C3795 INVX1_LOC_84/A INVX1_LOC_75/Y 0.10fF
C3796 NAND2X1_LOC_542/A INVX1_LOC_520/A 0.03fF
C3797 INVX1_LOC_682/Y NAND2X1_LOC_464/a_36_24# 0.00fF
C3798 INVX1_LOC_17/Y INVX1_LOC_242/Y 0.07fF
C3799 INVX1_LOC_581/A INVX1_LOC_62/Y 0.08fF
C3800 INVX1_LOC_367/Y INVX1_LOC_247/Y 0.15fF
C3801 INVX1_LOC_62/Y INVX1_LOC_633/Y 0.14fF
C3802 INVX1_LOC_501/A INVX1_LOC_48/Y 0.01fF
C3803 INVX1_LOC_491/A NAND2X1_LOC_220/a_36_24# 0.00fF
C3804 INVX1_LOC_316/Y INVX1_LOC_657/A 0.01fF
C3805 INVX1_LOC_452/A INVX1_LOC_244/Y 0.12fF
C3806 INVX1_LOC_134/Y INVX1_LOC_364/A 0.01fF
C3807 INVX1_LOC_35/Y INVX1_LOC_90/Y 0.13fF
C3808 INVX1_LOC_360/A NAND2X1_LOC_604/a_36_24# 0.00fF
C3809 INVX1_LOC_17/Y INVX1_LOC_487/A 0.03fF
C3810 INVX1_LOC_47/Y INVX1_LOC_49/Y 0.39fF
C3811 INVX1_LOC_520/Y INVX1_LOC_199/Y 0.02fF
C3812 INVX1_LOC_74/Y NAND2X1_LOC_418/Y 0.01fF
C3813 INVX1_LOC_129/A INVX1_LOC_75/Y 0.01fF
C3814 NAND2X1_LOC_557/B INVX1_LOC_49/Y 0.05fF
C3815 NAND2X1_LOC_387/Y INVX1_LOC_26/Y 0.02fF
C3816 INVX1_LOC_317/A INVX1_LOC_9/Y 0.01fF
C3817 INVX1_LOC_14/A INVX1_LOC_588/A 0.04fF
C3818 INVX1_LOC_41/Y INVX1_LOC_259/Y 0.03fF
C3819 INVX1_LOC_145/Y INVX1_LOC_598/Y 0.22fF
C3820 NAND2X1_LOC_448/B INVX1_LOC_90/Y 0.03fF
C3821 INVX1_LOC_54/Y INVX1_LOC_614/Y 0.00fF
C3822 INVX1_LOC_469/A INVX1_LOC_634/Y 0.03fF
C3823 INVX1_LOC_620/A INVX1_LOC_90/Y 0.01fF
C3824 VDD INVX1_LOC_615/Y 0.21fF
C3825 INVX1_LOC_280/Y INVX1_LOC_280/A 0.01fF
C3826 INVX1_LOC_523/Y INVX1_LOC_100/Y 0.07fF
C3827 INVX1_LOC_662/A INVX1_LOC_58/Y 0.12fF
C3828 NAND2X1_LOC_569/a_36_24# INVX1_LOC_443/A 0.02fF
C3829 INVX1_LOC_655/A NAND2X1_LOC_342/A 0.14fF
C3830 INVX1_LOC_556/Y INVX1_LOC_109/A -0.00fF
C3831 NAND2X1_LOC_707/B INVX1_LOC_41/Y 0.00fF
C3832 INVX1_LOC_519/Y NAND2X1_LOC_542/A 1.72fF
C3833 INVX1_LOC_469/Y INVX1_LOC_347/A 0.02fF
C3834 INVX1_LOC_350/Y INVX1_LOC_347/A -0.00fF
C3835 NAND2X1_LOC_148/B NAND2X1_LOC_843/B 0.02fF
C3836 INVX1_LOC_665/A INVX1_LOC_6/Y 0.52fF
C3837 INVX1_LOC_62/Y INVX1_LOC_490/A 0.27fF
C3838 INVX1_LOC_49/Y INVX1_LOC_119/Y 0.20fF
C3839 INVX1_LOC_400/Y INVX1_LOC_192/A 0.02fF
C3840 INVX1_LOC_117/Y INVX1_LOC_666/Y 0.07fF
C3841 INVX1_LOC_49/Y NAND2X1_LOC_66/Y 0.37fF
C3842 INVX1_LOC_44/Y INVX1_LOC_79/A 0.09fF
C3843 INVX1_LOC_69/Y NAND2X1_LOC_843/B 0.04fF
C3844 NAND2X1_LOC_123/B INVX1_LOC_168/Y 0.18fF
C3845 INVX1_LOC_63/Y INVX1_LOC_621/A 0.24fF
C3846 INVX1_LOC_479/A INVX1_LOC_77/Y 0.17fF
C3847 INVX1_LOC_446/A INVX1_LOC_578/A 0.02fF
C3848 VDD INVX1_LOC_37/Y 0.21fF
C3849 NAND2X1_LOC_615/Y INVX1_LOC_388/A 0.00fF
C3850 INVX1_LOC_69/Y INVX1_LOC_625/Y 0.11fF
C3851 NAND2X1_LOC_334/B INVX1_LOC_635/Y 0.02fF
C3852 NAND2X1_LOC_249/Y INVX1_LOC_556/A 0.07fF
C3853 VDD INVX1_LOC_395/A 5.74fF
C3854 INVX1_LOC_368/Y INVX1_LOC_245/A 0.01fF
C3855 INVX1_LOC_69/Y INVX1_LOC_91/Y 0.01fF
C3856 INVX1_LOC_41/Y INVX1_LOC_114/A 0.17fF
C3857 VDD INVX1_LOC_162/Y 0.21fF
C3858 INVX1_LOC_79/A INVX1_LOC_347/A 0.07fF
C3859 NAND2X1_LOC_847/A INVX1_LOC_212/A -0.02fF
C3860 VDD INVX1_LOC_362/Y 0.22fF
C3861 NAND2X1_LOC_242/A INVX1_LOC_96/Y 0.02fF
C3862 NAND2X1_LOC_543/B INVX1_LOC_270/A 0.01fF
C3863 NAND2X1_LOC_567/a_36_24# INVX1_LOC_442/A 0.00fF
C3864 NAND2X1_LOC_287/a_36_24# INVX1_LOC_669/A 0.00fF
C3865 NAND2X1_LOC_239/a_36_24# INVX1_LOC_586/A 0.00fF
C3866 VDD INVX1_LOC_678/Y 0.21fF
C3867 NAND2X1_LOC_45/Y INVX1_LOC_76/Y 0.05fF
C3868 INVX1_LOC_588/A NAND2X1_LOC_609/B 0.00fF
C3869 INVX1_LOC_51/A INVX1_LOC_51/Y 0.05fF
C3870 NAND2X1_LOC_475/A NAND2X1_LOC_318/A 0.08fF
C3871 NAND2X1_LOC_780/B INVX1_LOC_610/Y 0.07fF
C3872 VDD INVX1_LOC_683/Y 0.30fF
C3873 INVX1_LOC_84/A NAND2X1_LOC_20/a_36_24# 0.00fF
C3874 INVX1_LOC_395/A INVX1_LOC_510/Y 0.57fF
C3875 INVX1_LOC_275/Y INVX1_LOC_275/A 0.03fF
C3876 INVX1_LOC_564/A INVX1_LOC_586/A 0.01fF
C3877 INVX1_LOC_319/Y INVX1_LOC_586/A 0.01fF
C3878 NAND2X1_LOC_778/a_36_24# INVX1_LOC_547/Y 0.01fF
C3879 NAND2X1_LOC_498/Y NAND2X1_LOC_498/B 0.01fF
C3880 NAND2X1_LOC_373/Y INVX1_LOC_545/Y 0.12fF
C3881 NAND2X1_LOC_88/B NAND2X1_LOC_88/Y 0.33fF
C3882 INVX1_LOC_560/A NAND2X1_LOC_180/B 0.02fF
C3883 INVX1_LOC_36/A INVX1_LOC_76/Y 0.01fF
C3884 INVX1_LOC_570/A INVX1_LOC_76/Y 0.03fF
C3885 INVX1_LOC_222/Y INVX1_LOC_661/Y 0.01fF
C3886 INVX1_LOC_192/Y NAND2X1_LOC_336/B 0.01fF
C3887 INVX1_LOC_301/A INVX1_LOC_17/Y 0.07fF
C3888 INVX1_LOC_206/Y INVX1_LOC_670/Y 0.19fF
C3889 NAND2X1_LOC_173/Y INVX1_LOC_51/Y 3.79fF
C3890 INVX1_LOC_614/A INVX1_LOC_395/A 0.08fF
C3891 INVX1_LOC_86/Y NAND2X1_LOC_86/Y 0.01fF
C3892 VDD INVX1_LOC_189/Y 0.35fF
C3893 INVX1_LOC_459/A INVX1_LOC_50/Y 0.09fF
C3894 NAND2X1_LOC_69/B INVX1_LOC_54/Y 0.03fF
C3895 INVX1_LOC_446/A NAND2X1_LOC_527/Y 0.26fF
C3896 INVX1_LOC_438/Y INVX1_LOC_442/Y 0.19fF
C3897 NAND2X1_LOC_636/A INVX1_LOC_50/Y 0.00fF
C3898 INVX1_LOC_203/Y INVX1_LOC_59/Y 0.01fF
C3899 INVX1_LOC_566/Y INVX1_LOC_586/A 0.01fF
C3900 INVX1_LOC_20/Y INVX1_LOC_286/Y 0.03fF
C3901 NAND2X1_LOC_475/A INVX1_LOC_202/Y 0.03fF
C3902 INVX1_LOC_679/Y INVX1_LOC_107/A 0.02fF
C3903 INVX1_LOC_191/Y INVX1_LOC_194/Y 0.02fF
C3904 NAND2X1_LOC_567/a_36_24# INVX1_LOC_116/Y 0.00fF
C3905 INVX1_LOC_412/Y INVX1_LOC_352/Y 0.03fF
C3906 NAND2X1_LOC_780/B INVX1_LOC_48/Y 0.01fF
C3907 INVX1_LOC_542/A INVX1_LOC_358/Y 0.01fF
C3908 INVX1_LOC_203/Y INVX1_LOC_48/Y 0.21fF
C3909 INVX1_LOC_335/Y INVX1_LOC_542/A 0.00fF
C3910 VDD INVX1_LOC_31/Y 1.62fF
C3911 INVX1_LOC_602/A INVX1_LOC_55/Y 0.08fF
C3912 INVX1_LOC_297/A INVX1_LOC_381/A 0.05fF
C3913 INVX1_LOC_410/Y INVX1_LOC_159/Y 0.03fF
C3914 INVX1_LOC_51/Y NAND2X1_LOC_413/Y 0.58fF
C3915 INVX1_LOC_468/Y INVX1_LOC_374/A 0.01fF
C3916 INVX1_LOC_11/Y INVX1_LOC_140/Y 0.04fF
C3917 INVX1_LOC_670/Y INVX1_LOC_242/A 0.46fF
C3918 NAND2X1_LOC_45/Y INVX1_LOC_108/A 0.03fF
C3919 INVX1_LOC_308/Y INVX1_LOC_50/Y 0.01fF
C3920 INVX1_LOC_98/A INVX1_LOC_99/Y 0.01fF
C3921 NAND2X1_LOC_122/Y INVX1_LOC_145/Y 0.03fF
C3922 INVX1_LOC_586/A INVX1_LOC_367/Y 0.03fF
C3923 INVX1_LOC_273/A INVX1_LOC_145/Y 0.00fF
C3924 INVX1_LOC_435/A INVX1_LOC_45/Y 0.00fF
C3925 INVX1_LOC_454/A INVX1_LOC_69/Y 0.03fF
C3926 VDD INVX1_LOC_641/A -0.00fF
C3927 INVX1_LOC_617/Y INVX1_LOC_377/A 0.01fF
C3928 VDD NAND2X1_LOC_675/B 0.01fF
C3929 INVX1_LOC_76/Y INVX1_LOC_99/Y 0.20fF
C3930 INVX1_LOC_80/A INVX1_LOC_486/Y 0.07fF
C3931 NAND2X1_LOC_786/B INVX1_LOC_615/Y 0.01fF
C3932 INVX1_LOC_228/Y INVX1_LOC_31/Y 3.63fF
C3933 INVX1_LOC_300/A INVX1_LOC_286/Y 0.02fF
C3934 INVX1_LOC_617/Y NAND2X1_LOC_595/Y 0.01fF
C3935 INVX1_LOC_206/Y INVX1_LOC_253/Y 0.02fF
C3936 INVX1_LOC_20/Y INVX1_LOC_17/Y 0.36fF
C3937 NAND2X1_LOC_337/a_36_24# NAND2X1_LOC_267/A 0.00fF
C3938 INVX1_LOC_678/Y INVX1_LOC_684/A 0.15fF
C3939 NAND2X1_LOC_697/Y INVX1_LOC_522/Y 0.01fF
C3940 INVX1_LOC_651/Y NAND2X1_LOC_106/B 0.02fF
C3941 INVX1_LOC_335/Y NAND2X1_LOC_596/a_36_24# 0.01fF
C3942 VDD INVX1_LOC_682/Y 0.21fF
C3943 INVX1_LOC_246/Y INVX1_LOC_367/Y 0.01fF
C3944 NAND2X1_LOC_513/Y INVX1_LOC_89/Y 0.07fF
C3945 INVX1_LOC_393/Y INVX1_LOC_69/Y 0.02fF
C3946 NAND2X1_LOC_140/a_36_24# INVX1_LOC_47/Y 0.01fF
C3947 INVX1_LOC_206/Y INVX1_LOC_63/Y 2.76fF
C3948 INVX1_LOC_17/Y NAND2X1_LOC_473/a_36_24# 0.00fF
C3949 NAND2X1_LOC_638/A NAND2X1_LOC_755/B 0.05fF
C3950 INVX1_LOC_510/Y INVX1_LOC_31/Y 0.72fF
C3951 NAND2X1_LOC_396/a_36_24# INVX1_LOC_63/Y 0.00fF
C3952 NAND2X1_LOC_748/a_36_24# INVX1_LOC_366/A 0.01fF
C3953 INVX1_LOC_321/Y INVX1_LOC_12/Y 0.03fF
C3954 NAND2X1_LOC_545/B INVX1_LOC_35/Y 0.03fF
C3955 INVX1_LOC_106/A NAND2X1_LOC_113/a_36_24# 0.02fF
C3956 NAND2X1_LOC_498/B INVX1_LOC_47/Y 0.06fF
C3957 INVX1_LOC_274/Y INVX1_LOC_275/A 0.00fF
C3958 INVX1_LOC_123/A INVX1_LOC_76/Y 0.02fF
C3959 INVX1_LOC_11/Y INVX1_LOC_486/Y 0.08fF
C3960 NAND2X1_LOC_176/Y INVX1_LOC_79/A 0.01fF
C3961 NAND2X1_LOC_520/A INVX1_LOC_45/Y 0.00fF
C3962 INVX1_LOC_356/A INVX1_LOC_498/A 0.04fF
C3963 INVX1_LOC_54/Y INVX1_LOC_634/A 0.01fF
C3964 INVX1_LOC_21/Y NAND2X1_LOC_403/A 0.00fF
C3965 INVX1_LOC_103/Y INVX1_LOC_683/Y 0.00fF
C3966 INVX1_LOC_315/Y INVX1_LOC_204/Y 0.03fF
C3967 VDD INVX1_LOC_473/Y 0.14fF
C3968 NAND2X1_LOC_23/a_36_24# NAND2X1_LOC_626/Y 0.00fF
C3969 INVX1_LOC_595/Y INVX1_LOC_310/Y 0.02fF
C3970 INVX1_LOC_47/Y INVX1_LOC_76/Y 0.17fF
C3971 INVX1_LOC_17/Y INVX1_LOC_300/A 0.17fF
C3972 INVX1_LOC_442/Y INVX1_LOC_116/Y 0.00fF
C3973 NAND2X1_LOC_533/a_36_24# INVX1_LOC_74/Y 0.00fF
C3974 INVX1_LOC_635/A INVX1_LOC_50/Y 0.03fF
C3975 INVX1_LOC_335/Y INVX1_LOC_259/Y 0.03fF
C3976 INVX1_LOC_395/A NAND2X1_LOC_786/B 0.07fF
C3977 INVX1_LOC_502/Y INVX1_LOC_49/Y 0.04fF
C3978 INVX1_LOC_602/A INVX1_LOC_18/Y 0.09fF
C3979 NAND2X1_LOC_174/a_36_24# INVX1_LOC_99/Y 0.00fF
C3980 NAND2X1_LOC_845/a_36_24# NAND2X1_LOC_52/Y 0.00fF
C3981 INVX1_LOC_317/Y INVX1_LOC_9/Y 0.04fF
C3982 INVX1_LOC_442/Y INVX1_LOC_219/Y 0.10fF
C3983 INVX1_LOC_396/Y INVX1_LOC_63/Y 0.05fF
C3984 INVX1_LOC_35/Y INVX1_LOC_98/Y 0.16fF
C3985 INVX1_LOC_253/Y INVX1_LOC_686/A 0.02fF
C3986 INVX1_LOC_11/Y INVX1_LOC_252/A 0.03fF
C3987 INVX1_LOC_681/A INVX1_LOC_681/Y 0.01fF
C3988 NAND2X1_LOC_475/A INVX1_LOC_92/Y 0.02fF
C3989 INVX1_LOC_59/Y INVX1_LOC_194/Y 0.03fF
C3990 INVX1_LOC_80/A INVX1_LOC_6/Y 0.06fF
C3991 INVX1_LOC_409/Y INVX1_LOC_634/Y 0.21fF
C3992 NAND2X1_LOC_768/A INVX1_LOC_6/Y 0.09fF
C3993 INVX1_LOC_679/Y NAND2X1_LOC_285/A 0.02fF
C3994 NAND2X1_LOC_498/B INVX1_LOC_119/Y -0.01fF
C3995 NAND2X1_LOC_383/Y INVX1_LOC_245/A 0.03fF
C3996 INVX1_LOC_686/A INVX1_LOC_63/Y 0.07fF
C3997 INVX1_LOC_375/A INVX1_LOC_468/A 0.32fF
C3998 INVX1_LOC_412/Y NAND2X1_LOC_438/a_36_24# 0.00fF
C3999 INPUT_7 INVX1_LOC_58/Y 0.08fF
C4000 INVX1_LOC_612/Y INVX1_LOC_137/Y 0.29fF
C4001 INVX1_LOC_202/Y INVX1_LOC_153/A 0.02fF
C4002 INVX1_LOC_194/Y INVX1_LOC_48/Y 0.01fF
C4003 INVX1_LOC_76/Y INVX1_LOC_119/Y 0.07fF
C4004 INVX1_LOC_360/Y INVX1_LOC_93/Y 0.07fF
C4005 INVX1_LOC_500/A INVX1_LOC_147/Y 0.24fF
C4006 INVX1_LOC_12/Y INVX1_LOC_77/Y 0.19fF
C4007 INVX1_LOC_158/Y INVX1_LOC_31/Y 0.11fF
C4008 INVX1_LOC_166/A INVX1_LOC_303/Y 0.06fF
C4009 INVX1_LOC_31/Y INVX1_LOC_509/A 0.04fF
C4010 INVX1_LOC_588/Y INVX1_LOC_587/Y 0.06fF
C4011 INVX1_LOC_661/A INVX1_LOC_664/A 0.20fF
C4012 NAND2X1_LOC_198/a_36_24# INVX1_LOC_178/A 0.01fF
C4013 INVX1_LOC_291/A INVX1_LOC_90/Y 0.07fF
C4014 INVX1_LOC_93/Y INVX1_LOC_105/A 0.05fF
C4015 INVX1_LOC_47/Y NAND2X1_LOC_446/a_36_24# 0.01fF
C4016 NAND2X1_LOC_24/Y INVX1_LOC_26/Y 0.07fF
C4017 INVX1_LOC_51/Y INVX1_LOC_441/A -0.00fF
C4018 INVX1_LOC_201/Y INVX1_LOC_199/Y 0.00fF
C4019 INVX1_LOC_11/Y INVX1_LOC_6/Y 1.39fF
C4020 NAND2X1_LOC_94/a_36_24# INVX1_LOC_94/A 0.02fF
C4021 NAND2X1_LOC_43/Y INVX1_LOC_49/Y 0.06fF
C4022 INVX1_LOC_312/A INVX1_LOC_79/A 0.00fF
C4023 NAND2X1_LOC_820/a_36_24# INVX1_LOC_655/A 0.01fF
C4024 INVX1_LOC_679/A INVX1_LOC_58/Y 0.00fF
C4025 INVX1_LOC_355/A NAND2X1_LOC_832/A 0.01fF
C4026 NAND2X1_LOC_391/A INVX1_LOC_79/A 0.05fF
C4027 INVX1_LOC_49/Y NAND2X1_LOC_276/a_36_24# 0.01fF
C4028 INVX1_LOC_44/Y INVX1_LOC_59/Y 0.03fF
C4029 INVX1_LOC_54/Y INVX1_LOC_633/A 0.03fF
C4030 INVX1_LOC_360/Y INVX1_LOC_675/A 0.17fF
C4031 INVX1_LOC_586/A INVX1_LOC_625/Y 0.02fF
C4032 INVX1_LOC_326/Y INVX1_LOC_46/Y 0.65fF
C4033 INVX1_LOC_335/Y INVX1_LOC_114/A 0.03fF
C4034 INVX1_LOC_361/Y INVX1_LOC_69/Y 0.10fF
C4035 INVX1_LOC_406/Y INVX1_LOC_450/Y 0.01fF
C4036 INVX1_LOC_21/Y INVX1_LOC_114/A 0.01fF
C4037 INVX1_LOC_69/Y NAND2X1_LOC_333/B 0.11fF
C4038 INVX1_LOC_44/Y INVX1_LOC_48/Y 0.18fF
C4039 INVX1_LOC_312/Y NAND2X1_LOC_843/B 0.01fF
C4040 INVX1_LOC_31/Y INVX1_LOC_346/A 0.01fF
C4041 INVX1_LOC_79/A NAND2X1_LOC_418/Y 0.13fF
C4042 INVX1_LOC_298/A INVX1_LOC_659/A 0.02fF
C4043 NAND2X1_LOC_677/Y INVX1_LOC_614/Y 0.29fF
C4044 INVX1_LOC_555/A NAND2X1_LOC_697/a_36_24# 0.00fF
C4045 INVX1_LOC_518/A INVX1_LOC_510/A 0.72fF
C4046 INVX1_LOC_119/Y NAND2X1_LOC_446/a_36_24# 0.00fF
C4047 NAND2X1_LOC_836/B INVX1_LOC_93/A 0.03fF
C4048 INVX1_LOC_484/A INVX1_LOC_486/A 0.17fF
C4049 INVX1_LOC_542/Y INVX1_LOC_58/Y 0.19fF
C4050 INVX1_LOC_261/Y INVX1_LOC_69/Y 0.07fF
C4051 INVX1_LOC_382/A NAND2X1_LOC_476/a_36_24# 0.02fF
C4052 INVX1_LOC_103/Y INVX1_LOC_682/Y 0.04fF
C4053 INVX1_LOC_166/A INVX1_LOC_9/Y 0.07fF
C4054 INVX1_LOC_282/A INVX1_LOC_244/Y 0.31fF
C4055 NAND2X1_LOC_847/A INVX1_LOC_66/A 0.02fF
C4056 INVX1_LOC_650/Y INVX1_LOC_655/A 0.03fF
C4057 INVX1_LOC_89/Y NAND2X1_LOC_615/Y 0.02fF
C4058 NAND2X1_LOC_509/a_36_24# INVX1_LOC_26/Y 0.00fF
C4059 INVX1_LOC_31/Y NAND2X1_LOC_786/B 0.01fF
C4060 NAND2X1_LOC_646/A NAND2X1_LOC_609/B 0.06fF
C4061 NAND2X1_LOC_111/Y INVX1_LOC_9/Y 0.45fF
C4062 NAND2X1_LOC_753/Y INVX1_LOC_272/A 0.02fF
C4063 NAND2X1_LOC_369/a_36_24# INVX1_LOC_634/Y 0.00fF
C4064 INVX1_LOC_193/A INVX1_LOC_75/Y 0.01fF
C4065 INVX1_LOC_100/Y NAND2X1_LOC_814/Y 0.01fF
C4066 NAND2X1_LOC_475/A INVX1_LOC_297/Y 0.01fF
C4067 INVX1_LOC_166/A INVX1_LOC_62/Y 0.03fF
C4068 NAND2X1_LOC_192/A NAND2X1_LOC_189/a_36_24# 0.02fF
C4069 VDD INVX1_LOC_426/A 0.01fF
C4070 INVX1_LOC_31/Y INVX1_LOC_635/Y 0.03fF
C4071 INVX1_LOC_99/A INVX1_LOC_92/A 0.04fF
C4072 NAND2X1_LOC_184/Y NAND2X1_LOC_497/a_36_24# 0.00fF
C4073 INVX1_LOC_479/A INVX1_LOC_463/Y 0.04fF
C4074 INVX1_LOC_49/Y NAND2X1_LOC_627/Y 0.03fF
C4075 NAND2X1_LOC_136/Y INVX1_LOC_9/Y 0.10fF
C4076 NAND2X1_LOC_836/B INVX1_LOC_621/A 0.09fF
C4077 INVX1_LOC_63/Y NAND2X1_LOC_609/B 1.17fF
C4078 INVX1_LOC_79/A INVX1_LOC_226/Y 0.01fF
C4079 INVX1_LOC_574/A INVX1_LOC_570/Y 0.05fF
C4080 INVX1_LOC_531/Y INVX1_LOC_9/Y 0.00fF
C4081 INVX1_LOC_224/Y INVX1_LOC_560/Y 0.62fF
C4082 INVX1_LOC_404/Y NAND2X1_LOC_271/B 0.00fF
C4083 INVX1_LOC_418/A NAND2X1_LOC_322/Y 0.02fF
C4084 INVX1_LOC_26/Y INVX1_LOC_190/A 0.37fF
C4085 VDD NAND2X1_LOC_505/Y 0.13fF
C4086 NAND2X1_LOC_274/B INVX1_LOC_479/A 0.05fF
C4087 INVX1_LOC_567/A NAND2X1_LOC_704/B 0.00fF
C4088 VDD INVX1_LOC_51/Y 3.44fF
C4089 NAND2X1_LOC_543/B NAND2X1_LOC_318/A 0.00fF
C4090 INVX1_LOC_454/A INVX1_LOC_586/A 0.08fF
C4091 NAND2X1_LOC_735/a_36_24# NAND2X1_LOC_457/A 0.00fF
C4092 INVX1_LOC_206/Y INVX1_LOC_374/A 0.06fF
C4093 NAND2X1_LOC_580/a_36_24# INVX1_LOC_434/A 0.00fF
C4094 VDD INVX1_LOC_266/A 0.54fF
C4095 INVX1_LOC_442/A INVX1_LOC_412/A 0.16fF
C4096 NAND2X1_LOC_475/A INVX1_LOC_76/Y 0.04fF
C4097 INVX1_LOC_273/Y INVX1_LOC_620/Y 0.05fF
C4098 INVX1_LOC_393/Y INVX1_LOC_586/A 0.01fF
C4099 NAND2X1_LOC_554/a_36_24# INVX1_LOC_367/A -0.02fF
C4100 INVX1_LOC_603/Y NAND2X1_LOC_790/B 0.02fF
C4101 VDD INVX1_LOC_365/Y 0.21fF
C4102 INVX1_LOC_133/Y INVX1_LOC_575/A 0.00fF
C4103 INVX1_LOC_224/Y INVX1_LOC_84/A 0.02fF
C4104 INVX1_LOC_222/Y NAND2X1_LOC_260/Y 0.19fF
C4105 INVX1_LOC_447/A INVX1_LOC_134/Y 0.01fF
C4106 INVX1_LOC_392/Y INVX1_LOC_45/Y 0.12fF
C4107 INVX1_LOC_600/A INVX1_LOC_596/Y 0.03fF
C4108 INPUT_0 NAND2X1_LOC_39/Y 0.04fF
C4109 INVX1_LOC_20/Y NAND2X1_LOC_592/B 0.03fF
C4110 INVX1_LOC_564/A INVX1_LOC_272/Y 0.14fF
C4111 INVX1_LOC_301/A INVX1_LOC_545/A 0.01fF
C4112 NAND2X1_LOC_543/B INVX1_LOC_349/Y 0.00fF
C4113 INVX1_LOC_524/Y NAND2X1_LOC_506/B 0.14fF
C4114 INVX1_LOC_412/Y INVX1_LOC_67/Y 0.01fF
C4115 INVX1_LOC_601/A GATE_222 0.06fF
C4116 INVX1_LOC_68/Y INVX1_LOC_287/Y 0.00fF
C4117 INVX1_LOC_21/Y NAND2X1_LOC_457/A 0.03fF
C4118 INVX1_LOC_410/Y INVX1_LOC_377/A 0.09fF
C4119 VDD INVX1_LOC_500/Y 0.21fF
C4120 NAND2X1_LOC_336/B INVX1_LOC_442/A 0.00fF
C4121 VDD INVX1_LOC_40/Y 0.36fF
C4122 INVX1_LOC_45/Y INVX1_LOC_367/A 0.07fF
C4123 INVX1_LOC_445/Y INVX1_LOC_7/Y 0.07fF
C4124 NAND2X1_LOC_176/Y INVX1_LOC_48/Y 0.38fF
C4125 INVX1_LOC_578/A INVX1_LOC_129/A 0.08fF
C4126 INVX1_LOC_412/A INVX1_LOC_116/Y 0.09fF
C4127 INVX1_LOC_384/A INVX1_LOC_519/A 0.04fF
C4128 INVX1_LOC_435/Y INVX1_LOC_379/A 0.02fF
C4129 INVX1_LOC_76/Y INVX1_LOC_136/Y 0.01fF
C4130 INVX1_LOC_54/A INVX1_LOC_117/Y 0.01fF
C4131 NAND2X1_LOC_45/Y INVX1_LOC_32/Y 0.07fF
C4132 NAND2X1_LOC_637/A INVX1_LOC_261/Y 0.01fF
C4133 INVX1_LOC_400/A INVX1_LOC_45/Y 0.40fF
C4134 INVX1_LOC_392/A INVX1_LOC_45/Y 0.05fF
C4135 INVX1_LOC_404/Y INVX1_LOC_490/A 0.01fF
C4136 NAND2X1_LOC_704/B INVX1_LOC_252/A 0.01fF
C4137 INVX1_LOC_36/A INVX1_LOC_32/Y 0.02fF
C4138 INVX1_LOC_269/A INVX1_LOC_603/A 0.03fF
C4139 NAND2X1_LOC_498/Y INVX1_LOC_32/Y 0.24fF
C4140 INVX1_LOC_449/Y INVX1_LOC_218/A 0.01fF
C4141 INVX1_LOC_206/Y NAND2X1_LOC_836/B 0.18fF
C4142 INVX1_LOC_93/Y NAND2X1_LOC_506/B 0.15fF
C4143 INVX1_LOC_417/Y NAND2X1_LOC_391/A 0.00fF
C4144 INVX1_LOC_448/A INVX1_LOC_519/A 0.03fF
C4145 INVX1_LOC_361/Y INVX1_LOC_586/A 0.13fF
C4146 INVX1_LOC_93/Y INVX1_LOC_185/Y 0.05fF
C4147 INVX1_LOC_436/A INVX1_LOC_452/A 0.01fF
C4148 NAND2X1_LOC_336/a_36_24# INVX1_LOC_98/Y 0.00fF
C4149 INVX1_LOC_103/Y INVX1_LOC_51/Y 0.03fF
C4150 INVX1_LOC_586/A NAND2X1_LOC_333/B 0.07fF
C4151 INVX1_LOC_412/Y INVX1_LOC_347/Y 0.36fF
C4152 NAND2X1_LOC_765/a_36_24# INVX1_LOC_26/Y 0.00fF
C4153 INVX1_LOC_93/Y INVX1_LOC_45/Y 1.63fF
C4154 INVX1_LOC_435/A INVX1_LOC_293/Y 0.03fF
C4155 INVX1_LOC_85/Y NAND2X1_LOC_789/A 0.01fF
C4156 INVX1_LOC_281/A INVX1_LOC_586/A 0.12fF
C4157 INVX1_LOC_254/Y NAND2X1_LOC_538/B 0.03fF
C4158 INVX1_LOC_412/A INVX1_LOC_255/A 0.13fF
C4159 INVX1_LOC_596/A INVX1_LOC_35/Y 0.03fF
C4160 VDD INVX1_LOC_204/A 0.00fF
C4161 INPUT_7 INVX1_LOC_1/Y 0.15fF
C4162 INVX1_LOC_145/Y INVX1_LOC_519/A 0.02fF
C4163 INVX1_LOC_153/A INVX1_LOC_76/Y 0.00fF
C4164 INVX1_LOC_169/A INVX1_LOC_169/Y 0.04fF
C4165 INVX1_LOC_147/A INVX1_LOC_491/Y 0.03fF
C4166 INVX1_LOC_261/Y INVX1_LOC_586/A 0.03fF
C4167 INVX1_LOC_607/Y NAND2X1_LOC_147/B 0.04fF
C4168 INVX1_LOC_134/Y NAND2X1_LOC_606/Y 0.08fF
C4169 INVX1_LOC_492/Y INVX1_LOC_50/Y 0.01fF
C4170 INVX1_LOC_51/Y INVX1_LOC_346/A 0.05fF
C4171 INVX1_LOC_99/Y INVX1_LOC_7/Y 0.07fF
C4172 INPUT_3 INVX1_LOC_93/Y 0.06fF
C4173 NAND2X1_LOC_318/B INVX1_LOC_35/Y 0.00fF
C4174 INVX1_LOC_563/Y INVX1_LOC_272/A 0.09fF
C4175 NAND2X1_LOC_790/B INVX1_LOC_91/A 0.04fF
C4176 NAND2X1_LOC_391/A INVX1_LOC_48/Y 0.04fF
C4177 INVX1_LOC_320/Y INVX1_LOC_245/A 0.01fF
C4178 INVX1_LOC_63/Y INVX1_LOC_94/A 0.06fF
C4179 NAND2X1_LOC_498/B INVX1_LOC_15/Y 0.03fF
C4180 INVX1_LOC_451/A NAND2X1_LOC_415/B 0.47fF
C4181 INVX1_LOC_566/Y INVX1_LOC_6/Y 0.12fF
C4182 INVX1_LOC_372/Y INVX1_LOC_372/A 0.10fF
C4183 NAND2X1_LOC_710/A INVX1_LOC_89/Y 0.09fF
C4184 INVX1_LOC_43/Y INVX1_LOC_81/Y 0.02fF
C4185 NAND2X1_LOC_370/A INVX1_LOC_242/Y 0.02fF
C4186 INVX1_LOC_248/Y INVX1_LOC_440/A 0.01fF
C4187 INVX1_LOC_444/Y INVX1_LOC_453/Y 0.02fF
C4188 NAND2X1_LOC_837/A INVX1_LOC_59/A 0.03fF
C4189 INVX1_LOC_45/Y NAND2X1_LOC_334/B 0.00fF
C4190 INVX1_LOC_617/A INVX1_LOC_49/Y 0.02fF
C4191 INVX1_LOC_456/Y INVX1_LOC_40/Y 0.01fF
C4192 INVX1_LOC_249/Y INVX1_LOC_242/Y 0.02fF
C4193 INVX1_LOC_255/Y INVX1_LOC_114/A 0.02fF
C4194 INVX1_LOC_654/A INVX1_LOC_63/Y 0.03fF
C4195 INVX1_LOC_412/Y NAND2X1_LOC_439/a_36_24# 0.00fF
C4196 INVX1_LOC_58/Y INVX1_LOC_55/Y 0.04fF
C4197 INVX1_LOC_46/Y INVX1_LOC_600/A 0.03fF
C4198 INVX1_LOC_53/Y NAND2X1_LOC_753/Y 0.15fF
C4199 INVX1_LOC_345/Y INVX1_LOC_99/Y 0.03fF
C4200 INVX1_LOC_648/Y INVX1_LOC_669/A 0.03fF
C4201 INVX1_LOC_84/A INVX1_LOC_120/Y 0.01fF
C4202 INVX1_LOC_21/Y INVX1_LOC_87/Y 0.03fF
C4203 INVX1_LOC_32/Y INVX1_LOC_99/Y 2.54fF
C4204 NAND2X1_LOC_677/Y INVX1_LOC_633/A 0.01fF
C4205 INVX1_LOC_403/Y INVX1_LOC_556/Y 0.01fF
C4206 NAND2X1_LOC_353/a_36_24# INVX1_LOC_154/A 0.01fF
C4207 INVX1_LOC_277/A INVX1_LOC_672/A 0.04fF
C4208 INVX1_LOC_350/Y INVX1_LOC_252/Y 0.02fF
C4209 INVX1_LOC_254/Y INVX1_LOC_159/Y 0.01fF
C4210 INVX1_LOC_89/Y INVX1_LOC_155/Y 0.03fF
C4211 INVX1_LOC_137/Y INPUT_1 0.10fF
C4212 INVX1_LOC_626/A INVX1_LOC_6/Y 0.07fF
C4213 NAND2X1_LOC_829/Y INVX1_LOC_58/Y 0.00fF
C4214 NAND2X1_LOC_542/A INVX1_LOC_670/Y 0.08fF
C4215 INVX1_LOC_617/Y INVX1_LOC_518/A 0.00fF
C4216 INVX1_LOC_47/Y INVX1_LOC_7/Y 0.01fF
C4217 INVX1_LOC_17/Y NAND2X1_LOC_622/a_36_24# 0.00fF
C4218 INVX1_LOC_367/Y INVX1_LOC_6/Y 0.03fF
C4219 NAND2X1_LOC_190/A INVX1_LOC_166/A 0.00fF
C4220 INVX1_LOC_413/A NAND2X1_LOC_184/Y 0.03fF
C4221 INVX1_LOC_442/Y INVX1_LOC_69/Y 0.29fF
C4222 INVX1_LOC_117/Y NAND2X1_LOC_84/B 0.03fF
C4223 INVX1_LOC_669/A INVX1_LOC_242/A 0.07fF
C4224 INVX1_LOC_145/Y INVX1_LOC_659/A 0.04fF
C4225 INVX1_LOC_313/Y INVX1_LOC_6/Y 0.01fF
C4226 INVX1_LOC_338/A INVX1_LOC_338/Y 0.01fF
C4227 INVX1_LOC_501/A INVX1_LOC_155/Y 0.01fF
C4228 INVX1_LOC_170/Y INVX1_LOC_176/A 0.01fF
C4229 INVX1_LOC_651/Y NAND2X1_LOC_248/B 0.01fF
C4230 NAND2X1_LOC_467/A INVX1_LOC_62/Y 0.10fF
C4231 INVX1_LOC_406/Y INVX1_LOC_280/A 0.01fF
C4232 NAND2X1_LOC_97/A INVX1_LOC_211/A 0.00fF
C4233 INVX1_LOC_589/Y INVX1_LOC_32/Y 0.01fF
C4234 NAND2X1_LOC_538/B INVX1_LOC_479/A 0.05fF
C4235 NAND2X1_LOC_376/a_36_24# INVX1_LOC_41/Y 0.00fF
C4236 NAND2X1_LOC_615/B INVX1_LOC_77/Y 0.02fF
C4237 INVX1_LOC_376/Y INVX1_LOC_506/Y 0.04fF
C4238 INVX1_LOC_47/Y INVX1_LOC_32/Y 0.56fF
C4239 INVX1_LOC_248/Y INVX1_LOC_242/Y 0.03fF
C4240 NAND2X1_LOC_820/A NAND2X1_LOC_843/B 0.03fF
C4241 NAND2X1_LOC_557/B INVX1_LOC_32/Y 0.03fF
C4242 NAND2X1_LOC_66/Y INVX1_LOC_7/Y 0.08fF
C4243 INVX1_LOC_50/Y INVX1_LOC_168/Y 0.13fF
C4244 INVX1_LOC_11/Y INVX1_LOC_557/Y 0.00fF
C4245 INVX1_LOC_173/Y INVX1_LOC_199/Y 0.02fF
C4246 INVX1_LOC_202/Y INVX1_LOC_353/A 0.08fF
C4247 INVX1_LOC_421/A NAND2X1_LOC_275/a_36_24# 0.00fF
C4248 INVX1_LOC_79/A INVX1_LOC_252/Y 0.10fF
C4249 INVX1_LOC_105/A INVX1_LOC_128/A 0.23fF
C4250 INVX1_LOC_674/A NAND2X1_LOC_665/a_36_24# 0.01fF
C4251 INVX1_LOC_26/Y INVX1_LOC_259/Y 0.01fF
C4252 NAND2X1_LOC_387/Y NAND2X1_LOC_420/Y 0.02fF
C4253 NAND2X1_LOC_822/a_36_24# INVX1_LOC_656/A 0.00fF
C4254 INVX1_LOC_188/A NAND2X1_LOC_212/a_36_24# 0.02fF
C4255 INVX1_LOC_345/Y INVX1_LOC_119/Y 0.66fF
C4256 INVX1_LOC_303/Y INVX1_LOC_41/Y 0.23fF
C4257 INVX1_LOC_253/Y INVX1_LOC_376/Y 0.00fF
C4258 INVX1_LOC_32/Y INVX1_LOC_119/Y 0.03fF
C4259 INVX1_LOC_492/A INVX1_LOC_135/Y 0.01fF
C4260 INVX1_LOC_32/Y NAND2X1_LOC_66/Y 0.07fF
C4261 INVX1_LOC_587/Y INVX1_LOC_41/Y 0.14fF
C4262 VDD INVX1_LOC_618/A 0.00fF
C4263 NAND2X1_LOC_307/A INVX1_LOC_92/A 1.62fF
C4264 INVX1_LOC_621/Y INVX1_LOC_622/A 0.00fF
C4265 INVX1_LOC_479/A INVX1_LOC_159/Y 0.08fF
C4266 INVX1_LOC_204/Y INVX1_LOC_26/Y 0.02fF
C4267 INVX1_LOC_63/Y INVX1_LOC_376/Y 0.33fF
C4268 INVX1_LOC_49/Y INVX1_LOC_353/A 0.07fF
C4269 INVX1_LOC_301/Y INVX1_LOC_9/Y 0.01fF
C4270 INVX1_LOC_513/A INVX1_LOC_464/Y 0.20fF
C4271 INVX1_LOC_306/Y INVX1_LOC_41/Y 0.01fF
C4272 VDD NAND2X1_LOC_537/A 0.00fF
C4273 INVX1_LOC_6/Y NAND2X1_LOC_843/B 0.08fF
C4274 INVX1_LOC_376/A NAND2X1_LOC_123/B 0.19fF
C4275 INVX1_LOC_26/Y INVX1_LOC_82/Y 0.01fF
C4276 INVX1_LOC_62/Y INVX1_LOC_411/Y 0.01fF
C4277 INVX1_LOC_419/Y INVX1_LOC_92/A 0.01fF
C4278 INVX1_LOC_26/Y INVX1_LOC_114/A 0.03fF
C4279 INVX1_LOC_228/Y NAND2X1_LOC_537/A 0.06fF
C4280 INVX1_LOC_41/Y INVX1_LOC_9/Y 0.22fF
C4281 VDD INVX1_LOC_216/Y 0.26fF
C4282 NAND2X1_LOC_449/B NAND2X1_LOC_832/A 0.02fF
C4283 INPUT_6 NAND2X1_LOC_1/a_36_24# 0.00fF
C4284 NAND2X1_LOC_593/a_36_24# INVX1_LOC_638/A 0.01fF
C4285 NAND2X1_LOC_228/a_36_24# INVX1_LOC_586/A 0.01fF
C4286 INVX1_LOC_666/Y INVX1_LOC_245/A 0.02fF
C4287 INVX1_LOC_166/Y INVX1_LOC_41/Y 0.00fF
C4288 INVX1_LOC_395/A NAND2X1_LOC_378/a_36_24# 0.00fF
C4289 INVX1_LOC_452/Y VDD 0.21fF
C4290 INVX1_LOC_454/A INVX1_LOC_587/A 0.03fF
C4291 INVX1_LOC_62/Y INVX1_LOC_41/Y 3.01fF
C4292 INVX1_LOC_479/A INVX1_LOC_468/A 0.03fF
C4293 INVX1_LOC_554/A INVX1_LOC_336/Y 0.01fF
C4294 INVX1_LOC_395/A NAND2X1_LOC_506/B 0.03fF
C4295 VDD NAND2X1_LOC_13/Y 0.35fF
C4296 INVX1_LOC_41/Y NAND2X1_LOC_844/A 0.03fF
C4297 INVX1_LOC_510/A INVX1_LOC_109/Y 0.42fF
C4298 INVX1_LOC_395/A INVX1_LOC_185/Y 0.07fF
C4299 INVX1_LOC_505/Y INVX1_LOC_74/Y 0.09fF
C4300 INVX1_LOC_633/Y INVX1_LOC_638/A 0.08fF
C4301 NAND2X1_LOC_636/A NAND2X1_LOC_636/B 0.17fF
C4302 INVX1_LOC_395/A INVX1_LOC_45/Y 0.73fF
C4303 INVX1_LOC_533/Y NAND2X1_LOC_122/Y 0.15fF
C4304 INVX1_LOC_33/A INVX1_LOC_33/Y 0.01fF
C4305 INVX1_LOC_20/Y INVX1_LOC_127/A 0.15fF
C4306 INVX1_LOC_84/A INVX1_LOC_206/Y 0.17fF
C4307 NAND2X1_LOC_13/Y INVX1_LOC_228/Y -0.00fF
C4308 INVX1_LOC_362/Y INVX1_LOC_45/Y 0.07fF
C4309 INVX1_LOC_84/A NAND2X1_LOC_49/a_36_24# 0.01fF
C4310 INVX1_LOC_409/Y INVX1_LOC_115/A 0.00fF
C4311 INVX1_LOC_20/Y NAND2X1_LOC_370/A 0.00fF
C4312 INVX1_LOC_445/Y INVX1_LOC_424/Y 0.09fF
C4313 INVX1_LOC_121/Y INVX1_LOC_670/Y 0.01fF
C4314 INVX1_LOC_133/Y INVX1_LOC_575/Y 0.03fF
C4315 INVX1_LOC_68/Y NAND2X1_LOC_318/A 0.07fF
C4316 INVX1_LOC_203/Y INVX1_LOC_155/Y 0.03fF
C4317 INVX1_LOC_20/Y NAND2X1_LOC_122/Y 0.06fF
C4318 INVX1_LOC_459/A INVX1_LOC_117/Y 0.06fF
C4319 NAND2X1_LOC_122/a_36_24# INVX1_LOC_632/A 0.01fF
C4320 INVX1_LOC_451/A INVX1_LOC_453/A 0.16fF
C4321 INVX1_LOC_438/A INVX1_LOC_681/A 0.01fF
C4322 NAND2X1_LOC_636/A INVX1_LOC_117/Y 0.10fF
C4323 INVX1_LOC_95/Y INVX1_LOC_525/Y 0.01fF
C4324 INVX1_LOC_206/Y INVX1_LOC_129/A 0.03fF
C4325 INVX1_LOC_212/A NAND2X1_LOC_245/a_36_24# 0.01fF
C4326 INVX1_LOC_206/Y NAND2X1_LOC_67/Y 0.00fF
C4327 NAND2X1_LOC_61/A INVX1_LOC_31/Y 0.05fF
C4328 INVX1_LOC_395/A NAND2X1_LOC_376/Y 0.15fF
C4329 NAND2X1_LOC_467/A NAND2X1_LOC_163/a_36_24# 0.02fF
C4330 INVX1_LOC_395/A NAND2X1_LOC_69/Y 0.01fF
C4331 INVX1_LOC_581/A INVX1_LOC_144/Y 0.02fF
C4332 NAND2X1_LOC_332/B INVX1_LOC_519/A 0.03fF
C4333 INVX1_LOC_300/A NAND2X1_LOC_370/A 0.09fF
C4334 INVX1_LOC_38/A INVX1_LOC_12/Y 0.11fF
C4335 INVX1_LOC_290/Y INVX1_LOC_263/Y 0.13fF
C4336 NAND2X1_LOC_475/A INVX1_LOC_32/Y 0.09fF
C4337 INVX1_LOC_425/A INVX1_LOC_417/Y 0.01fF
C4338 INVX1_LOC_442/Y INVX1_LOC_586/A 0.07fF
C4339 INVX1_LOC_293/Y INVX1_LOC_367/A 0.07fF
C4340 INVX1_LOC_239/Y INVX1_LOC_132/A 0.01fF
C4341 NAND2X1_LOC_318/A INVX1_LOC_600/A 0.15fF
C4342 INVX1_LOC_549/A INVX1_LOC_117/Y 0.15fF
C4343 INVX1_LOC_449/A INVX1_LOC_406/Y 0.00fF
C4344 VDD INVX1_LOC_380/Y 0.22fF
C4345 INPUT_0 INVX1_LOC_670/A 0.07fF
C4346 INVX1_LOC_11/Y INVX1_LOC_269/Y 0.13fF
C4347 NAND2X1_LOC_122/Y INVX1_LOC_197/Y 0.09fF
C4348 INVX1_LOC_193/A INVX1_LOC_578/A 0.02fF
C4349 INVX1_LOC_548/A INVX1_LOC_45/Y 0.01fF
C4350 INVX1_LOC_602/A INVX1_LOC_635/A 0.03fF
C4351 NAND2X1_LOC_525/Y INVX1_LOC_50/Y 0.07fF
C4352 INVX1_LOC_273/A INVX1_LOC_197/Y 0.07fF
C4353 INVX1_LOC_396/A INVX1_LOC_96/Y 0.23fF
C4354 INVX1_LOC_68/Y INVX1_LOC_202/Y 0.00fF
C4355 VDD NAND2X1_LOC_668/Y 0.04fF
C4356 VDD INVX1_LOC_361/A 0.17fF
C4357 INVX1_LOC_17/Y INVX1_LOC_562/Y 0.01fF
C4358 NAND2X1_LOC_541/a_36_24# INVX1_LOC_6/Y 0.00fF
C4359 INVX1_LOC_20/Y INVX1_LOC_248/Y 0.07fF
C4360 INVX1_LOC_449/A NAND2X1_LOC_522/a_36_24# 0.00fF
C4361 INVX1_LOC_575/A NAND2X1_LOC_725/a_36_24# 0.02fF
C4362 VDD INVX1_LOC_196/Y 0.21fF
C4363 NAND2X1_LOC_516/Y INVX1_LOC_670/A 0.01fF
C4364 INVX1_LOC_393/Y INVX1_LOC_6/Y 0.01fF
C4365 INPUT_0 NAND2X1_LOC_606/a_36_24# 0.00fF
C4366 INVX1_LOC_206/Y INVX1_LOC_496/A 0.07fF
C4367 INVX1_LOC_222/Y INVX1_LOC_655/A 0.02fF
C4368 INVX1_LOC_129/A INVX1_LOC_686/A 0.06fF
C4369 INVX1_LOC_11/Y INVX1_LOC_381/A 0.07fF
C4370 INVX1_LOC_312/Y INVX1_LOC_442/Y 0.07fF
C4371 INVX1_LOC_412/A INVX1_LOC_69/Y 0.07fF
C4372 INVX1_LOC_53/Y NAND2X1_LOC_610/a_36_24# 0.00fF
C4373 NAND2X1_LOC_758/a_36_24# INVX1_LOC_26/Y 0.00fF
C4374 INVX1_LOC_31/Y INVX1_LOC_45/Y 0.67fF
C4375 INVX1_LOC_155/A INVX1_LOC_160/Y 0.01fF
C4376 NAND2X1_LOC_697/Y INVX1_LOC_581/A 0.02fF
C4377 INVX1_LOC_392/A INVX1_LOC_293/Y 0.03fF
C4378 INVX1_LOC_115/A NAND2X1_LOC_302/A 0.00fF
C4379 NAND2X1_LOC_755/a_36_24# INVX1_LOC_53/Y 0.00fF
C4380 INVX1_LOC_53/Y NAND2X1_LOC_285/B 0.01fF
C4381 INVX1_LOC_167/Y INVX1_LOC_50/Y 0.19fF
C4382 INVX1_LOC_502/Y INVX1_LOC_32/Y 0.03fF
C4383 INVX1_LOC_202/Y INVX1_LOC_250/Y 0.10fF
C4384 INVX1_LOC_176/Y INVX1_LOC_172/A 0.02fF
C4385 INVX1_LOC_307/A NAND2X1_LOC_378/Y 0.00fF
C4386 INPUT_3 NAND2X1_LOC_83/a_36_24# 0.00fF
C4387 NAND2X1_LOC_775/a_36_24# INVX1_LOC_160/A 0.00fF
C4388 INVX1_LOC_63/Y INVX1_LOC_253/A 0.00fF
C4389 INVX1_LOC_130/Y INVX1_LOC_99/Y 0.92fF
C4390 INVX1_LOC_53/Y NAND2X1_LOC_106/B 0.01fF
C4391 NAND2X1_LOC_775/B INVX1_LOC_134/Y 0.03fF
C4392 INVX1_LOC_11/Y INVX1_LOC_320/A 0.02fF
C4393 NAND2X1_LOC_457/A INVX1_LOC_26/Y 0.03fF
C4394 INVX1_LOC_656/A INVX1_LOC_59/A 0.01fF
C4395 INVX1_LOC_133/A GATE_662 0.04fF
C4396 INVX1_LOC_293/Y INVX1_LOC_93/Y 0.03fF
C4397 NAND2X1_LOC_307/A INPUT_1 0.03fF
C4398 INPUT_3 INVX1_LOC_31/Y 0.76fF
C4399 INVX1_LOC_12/Y INVX1_LOC_159/Y 0.05fF
C4400 INVX1_LOC_248/Y INVX1_LOC_197/Y 0.03fF
C4401 INVX1_LOC_581/A INVX1_LOC_575/Y 0.23fF
C4402 INVX1_LOC_375/A INVX1_LOC_518/A 0.08fF
C4403 NAND2X1_LOC_43/Y INVX1_LOC_7/Y 0.05fF
C4404 INVX1_LOC_117/Y INVX1_LOC_635/A 0.03fF
C4405 INVX1_LOC_53/Y NAND2X1_LOC_591/Y 0.03fF
C4406 INVX1_LOC_625/A INVX1_LOC_35/Y 0.02fF
C4407 INVX1_LOC_374/A INVX1_LOC_376/Y 0.35fF
C4408 NAND2X1_LOC_297/Y NAND2X1_LOC_296/Y 0.09fF
C4409 INVX1_LOC_117/Y NAND2X1_LOC_237/Y 0.01fF
C4410 INVX1_LOC_522/Y INVX1_LOC_476/A 0.00fF
C4411 INVX1_LOC_250/A INVX1_LOC_353/A 0.02fF
C4412 INVX1_LOC_513/A INVX1_LOC_145/Y 0.03fF
C4413 INVX1_LOC_335/Y INVX1_LOC_539/Y 0.11fF
C4414 NAND2X1_LOC_336/B INVX1_LOC_69/Y 0.00fF
C4415 INVX1_LOC_48/Y INVX1_LOC_252/Y 0.48fF
C4416 INVX1_LOC_54/Y INVX1_LOC_176/A 0.19fF
C4417 NAND2X1_LOC_513/A NAND2X1_LOC_647/A 0.01fF
C4418 NAND2X1_LOC_704/B INVX1_LOC_557/Y 0.05fF
C4419 INVX1_LOC_76/Y INVX1_LOC_353/A 0.07fF
C4420 INVX1_LOC_651/Y INVX1_LOC_664/A 0.04fF
C4421 INVX1_LOC_340/Y INVX1_LOC_461/Y 0.09fF
C4422 INVX1_LOC_117/Y INVX1_LOC_230/A 0.08fF
C4423 INVX1_LOC_640/A INVX1_LOC_641/Y 0.01fF
C4424 INVX1_LOC_137/Y INVX1_LOC_50/Y 0.07fF
C4425 INVX1_LOC_608/Y NAND2X1_LOC_106/Y 0.02fF
C4426 INVX1_LOC_506/A INVX1_LOC_504/Y 0.01fF
C4427 INVX1_LOC_683/A INVX1_LOC_66/A 0.01fF
C4428 INVX1_LOC_419/Y INPUT_1 0.03fF
C4429 INVX1_LOC_31/Y NAND2X1_LOC_69/Y 0.03fF
C4430 INVX1_LOC_400/Y INVX1_LOC_75/Y 0.07fF
C4431 INVX1_LOC_17/Y NAND2X1_LOC_106/Y 0.03fF
C4432 INVX1_LOC_21/Y INVX1_LOC_306/Y 0.01fF
C4433 INVX1_LOC_18/Y INVX1_LOC_1/Y 0.06fF
C4434 INVX1_LOC_636/A NAND2X1_LOC_590/a_36_24# 0.01fF
C4435 INVX1_LOC_100/A INVX1_LOC_178/A 0.13fF
C4436 NAND2X1_LOC_720/A NAND2X1_LOC_667/a_36_24# 0.02fF
C4437 INVX1_LOC_402/A INVX1_LOC_520/Y 0.05fF
C4438 INVX1_LOC_315/Y INVX1_LOC_62/Y 0.09fF
C4439 INPUT_0 NAND2X1_LOC_201/a_36_24# 0.00fF
C4440 INVX1_LOC_68/Y INVX1_LOC_92/Y 0.00fF
C4441 INVX1_LOC_267/Y INVX1_LOC_272/A 0.05fF
C4442 INVX1_LOC_145/A INVX1_LOC_40/Y 0.03fF
C4443 INVX1_LOC_153/A INVX1_LOC_32/Y 0.01fF
C4444 INVX1_LOC_21/Y INVX1_LOC_9/Y 0.08fF
C4445 INVX1_LOC_35/Y NAND2X1_LOC_52/Y 0.04fF
C4446 INVX1_LOC_315/Y INVX1_LOC_529/Y 0.02fF
C4447 NAND2X1_LOC_775/B INVX1_LOC_65/A 0.01fF
C4448 INVX1_LOC_80/A INVX1_LOC_100/Y 2.28fF
C4449 INVX1_LOC_155/A NAND2X1_LOC_267/A 0.06fF
C4450 INVX1_LOC_99/Y NAND2X1_LOC_405/a_36_24# 0.00fF
C4451 INVX1_LOC_517/Y INVX1_LOC_137/Y 0.08fF
C4452 INPUT_1 NAND2X1_LOC_342/A 0.03fF
C4453 INVX1_LOC_47/Y INVX1_LOC_110/A 0.04fF
C4454 INVX1_LOC_634/A INVX1_LOC_347/A 0.03fF
C4455 INVX1_LOC_32/Y INVX1_LOC_96/A 0.01fF
C4456 INVX1_LOC_54/Y INVX1_LOC_170/Y 0.01fF
C4457 INVX1_LOC_31/Y NAND2X1_LOC_837/A 0.72fF
C4458 INVX1_LOC_559/A INVX1_LOC_353/A 0.03fF
C4459 INVX1_LOC_358/Y INVX1_LOC_62/Y 0.03fF
C4460 NAND2X1_LOC_148/B NAND2X1_LOC_847/A 0.09fF
C4461 NAND2X1_LOC_288/a_36_24# INVX1_LOC_655/A 0.01fF
C4462 INVX1_LOC_444/Y INVX1_LOC_422/A 0.13fF
C4463 INVX1_LOC_80/A INVX1_LOC_74/Y 0.49fF
C4464 INVX1_LOC_35/Y INVX1_LOC_519/Y 0.05fF
C4465 INVX1_LOC_21/Y INVX1_LOC_62/Y 0.18fF
C4466 INVX1_LOC_100/A INVX1_LOC_58/Y 0.01fF
C4467 INVX1_LOC_49/Y INVX1_LOC_484/A 0.02fF
C4468 INVX1_LOC_17/Y NAND2X1_LOC_123/B 0.40fF
C4469 NAND2X1_LOC_267/A INVX1_LOC_9/Y 0.88fF
C4470 INVX1_LOC_11/Y INVX1_LOC_100/Y 0.23fF
C4471 INVX1_LOC_632/Y INVX1_LOC_259/Y 0.24fF
C4472 INVX1_LOC_508/A INVX1_LOC_476/A 0.36fF
C4473 INVX1_LOC_21/Y INVX1_LOC_13/Y 0.20fF
C4474 INVX1_LOC_502/A INPUT_1 0.53fF
C4475 INVX1_LOC_555/A INVX1_LOC_9/Y 0.02fF
C4476 INVX1_LOC_110/A INVX1_LOC_119/Y 0.03fF
C4477 NAND2X1_LOC_190/A INVX1_LOC_41/Y 0.02fF
C4478 INVX1_LOC_518/Y INVX1_LOC_520/A 0.20fF
C4479 INVX1_LOC_81/Y INVX1_LOC_190/A 0.01fF
C4480 INVX1_LOC_179/A INVX1_LOC_77/Y 0.04fF
C4481 INVX1_LOC_11/Y INVX1_LOC_74/Y 0.15fF
C4482 NAND2X1_LOC_274/B INVX1_LOC_66/A 0.06fF
C4483 NAND2X1_LOC_500/a_36_24# NAND2X1_LOC_844/A 0.00fF
C4484 INVX1_LOC_479/A INVX1_LOC_345/A 0.02fF
C4485 INVX1_LOC_41/Y INVX1_LOC_87/A 0.13fF
C4486 NAND2X1_LOC_409/Y INVX1_LOC_93/A 0.03fF
C4487 INVX1_LOC_17/Y INVX1_LOC_485/A 0.01fF
C4488 INVX1_LOC_421/A INVX1_LOC_75/Y 0.09fF
C4489 INVX1_LOC_17/Y INVX1_LOC_92/A 0.10fF
C4490 INVX1_LOC_223/A INVX1_LOC_46/Y 0.03fF
C4491 INVX1_LOC_496/A NAND2X1_LOC_609/B 0.09fF
C4492 INVX1_LOC_54/Y INVX1_LOC_611/A 0.02fF
C4493 INVX1_LOC_617/Y INVX1_LOC_109/Y 0.07fF
C4494 INVX1_LOC_518/Y INVX1_LOC_519/Y 0.09fF
C4495 INPUT_0 INVX1_LOC_616/Y 0.00fF
C4496 NAND2X1_LOC_274/B NAND2X1_LOC_601/Y 0.01fF
C4497 INVX1_LOC_100/Y INVX1_LOC_102/Y 0.02fF
C4498 NAND2X1_LOC_433/Y INVX1_LOC_74/Y 0.01fF
C4499 INVX1_LOC_435/Y INVX1_LOC_434/A 0.02fF
C4500 INVX1_LOC_409/Y INVX1_LOC_76/Y 0.03fF
C4501 INVX1_LOC_505/Y INVX1_LOC_79/A 0.06fF
C4502 NAND2X1_LOC_317/A INVX1_LOC_546/A 0.06fF
C4503 INVX1_LOC_191/Y INVX1_LOC_85/Y 0.00fF
C4504 NAND2X1_LOC_32/a_36_24# INVX1_LOC_395/A 0.00fF
C4505 VDD NAND2X1_LOC_152/B 0.03fF
C4506 NAND2X1_LOC_249/Y INVX1_LOC_651/A 0.01fF
C4507 INVX1_LOC_301/A INVX1_LOC_519/A 0.00fF
C4508 INVX1_LOC_412/A INVX1_LOC_586/A 0.12fF
C4509 NAND2X1_LOC_505/Y INVX1_LOC_45/Y 0.01fF
C4510 INVX1_LOC_579/Y NAND2X1_LOC_591/B 0.02fF
C4511 INPUT_0 NAND2X1_LOC_516/B 0.01fF
C4512 INVX1_LOC_68/Y INVX1_LOC_250/A 0.03fF
C4513 NAND2X1_LOC_331/A NAND2X1_LOC_467/A 0.01fF
C4514 INVX1_LOC_264/Y INVX1_LOC_495/A 0.01fF
C4515 INVX1_LOC_51/Y INVX1_LOC_45/Y 0.28fF
C4516 NAND2X1_LOC_756/Y INVX1_LOC_395/A 0.12fF
C4517 INVX1_LOC_85/Y INVX1_LOC_180/A 0.00fF
C4518 NAND2X1_LOC_242/A INVX1_LOC_80/A 2.05fF
C4519 INVX1_LOC_68/Y INVX1_LOC_98/A 0.09fF
C4520 NAND2X1_LOC_516/Y NAND2X1_LOC_516/B 0.01fF
C4521 NAND2X1_LOC_271/B INVX1_LOC_134/Y 0.02fF
C4522 INVX1_LOC_68/Y INVX1_LOC_76/Y 0.01fF
C4523 INVX1_LOC_588/Y INVX1_LOC_638/A 0.07fF
C4524 INVX1_LOC_3/Y INVX1_LOC_6/A 0.00fF
C4525 INPUT_6 NAND2X1_LOC_3/a_36_24# 0.00fF
C4526 INPUT_3 INVX1_LOC_51/Y 0.03fF
C4527 INVX1_LOC_293/Y INVX1_LOC_362/Y 0.19fF
C4528 INVX1_LOC_402/Y INPUT_0 0.01fF
C4529 INVX1_LOC_579/A INVX1_LOC_533/Y 0.18fF
C4530 NAND2X1_LOC_260/Y INVX1_LOC_445/A 0.05fF
C4531 INVX1_LOC_127/A NAND2X1_LOC_140/B 0.17fF
C4532 INVX1_LOC_250/Y INVX1_LOC_250/A 0.16fF
C4533 INVX1_LOC_425/A NAND2X1_LOC_129/a_36_24# 0.00fF
C4534 NAND2X1_LOC_271/B INVX1_LOC_235/A 0.01fF
C4535 NAND2X1_LOC_336/B INVX1_LOC_586/A 0.08fF
C4536 INPUT_0 INVX1_LOC_435/A 0.03fF
C4537 NAND2X1_LOC_543/B INVX1_LOC_32/Y 0.07fF
C4538 INVX1_LOC_308/Y INVX1_LOC_178/A 0.03fF
C4539 INVX1_LOC_516/Y INVX1_LOC_517/A 0.01fF
C4540 INVX1_LOC_402/Y NAND2X1_LOC_516/Y 0.01fF
C4541 INVX1_LOC_375/A INVX1_LOC_352/A 0.04fF
C4542 NAND2X1_LOC_164/Y INVX1_LOC_35/Y 0.37fF
C4543 NAND2X1_LOC_122/Y NAND2X1_LOC_298/a_36_24# 0.00fF
C4544 INVX1_LOC_560/A INVX1_LOC_194/A 0.03fF
C4545 INVX1_LOC_250/Y INVX1_LOC_76/Y 0.03fF
C4546 NAND2X1_LOC_66/a_36_24# INVX1_LOC_6/Y 0.00fF
C4547 INVX1_LOC_20/Y INVX1_LOC_579/A 0.03fF
C4548 INVX1_LOC_395/A NAND2X1_LOC_673/B 0.07fF
C4549 NAND2X1_LOC_45/Y NAND2X1_LOC_184/Y 0.05fF
C4550 INVX1_LOC_80/Y NAND2X1_LOC_79/B 0.17fF
C4551 VDD INVX1_LOC_581/Y 0.21fF
C4552 INVX1_LOC_20/Y INVX1_LOC_519/A 0.03fF
C4553 NAND2X1_LOC_14/a_36_24# INPUT_2 0.00fF
C4554 NAND2X1_LOC_636/A INVX1_LOC_58/Y 0.26fF
C4555 INVX1_LOC_564/A NAND2X1_LOC_720/A 0.02fF
C4556 INVX1_LOC_65/Y INVX1_LOC_35/Y 0.06fF
C4557 INVX1_LOC_47/A INVX1_LOC_169/A 0.01fF
C4558 INVX1_LOC_614/A NAND2X1_LOC_152/B 0.00fF
C4559 VDD NAND2X1_LOC_449/B 0.04fF
C4560 INVX1_LOC_45/Y INVX1_LOC_40/Y 0.01fF
C4561 GATE_579 INVX1_LOC_453/Y 0.23fF
C4562 INVX1_LOC_373/A NAND2X1_LOC_707/B 0.00fF
C4563 INVX1_LOC_551/Y NAND2X1_LOC_413/Y 0.23fF
C4564 NAND2X1_LOC_721/a_36_24# INVX1_LOC_298/A 0.00fF
C4565 INVX1_LOC_134/Y INVX1_LOC_633/Y 0.07fF
C4566 INVX1_LOC_106/A INVX1_LOC_101/Y 0.13fF
C4567 INVX1_LOC_412/Y INVX1_LOC_199/Y 0.15fF
C4568 VDD NAND2X1_LOC_121/Y 0.07fF
C4569 INVX1_LOC_254/A INVX1_LOC_45/Y 0.01fF
C4570 INVX1_LOC_558/A NAND2X1_LOC_659/a_36_24# 0.01fF
C4571 INVX1_LOC_308/Y INVX1_LOC_58/Y 0.02fF
C4572 INVX1_LOC_549/A INVX1_LOC_58/Y 0.09fF
C4573 INVX1_LOC_250/Y INVX1_LOC_559/A 0.01fF
C4574 INVX1_LOC_237/Y INVX1_LOC_66/A 0.01fF
C4575 INVX1_LOC_84/A INVX1_LOC_432/A 0.02fF
C4576 NAND2X1_LOC_788/A NAND2X1_LOC_274/B 0.57fF
C4577 INVX1_LOC_595/Y INVX1_LOC_311/Y 0.02fF
C4578 INVX1_LOC_384/A INVX1_LOC_670/A 0.04fF
C4579 NAND2X1_LOC_180/B NAND2X1_LOC_444/A 0.14fF
C4580 INVX1_LOC_202/Y NAND2X1_LOC_56/Y 0.00fF
C4581 VDD NAND2X1_LOC_301/B 0.47fF
C4582 INVX1_LOC_193/A INVX1_LOC_686/A 0.02fF
C4583 INVX1_LOC_617/A INVX1_LOC_32/Y 0.00fF
C4584 INVX1_LOC_137/Y NAND2X1_LOC_513/A 0.11fF
C4585 INVX1_LOC_372/Y INVX1_LOC_345/A 0.02fF
C4586 INVX1_LOC_300/A NAND2X1_LOC_334/a_36_24# 0.00fF
C4587 INVX1_LOC_117/Y INVX1_LOC_492/Y 0.01fF
C4588 NAND2X1_LOC_107/Y NAND2X1_LOC_106/B 0.12fF
C4589 INVX1_LOC_544/A INVX1_LOC_683/A 0.01fF
C4590 INVX1_LOC_140/Y INVX1_LOC_471/Y 0.01fF
C4591 INVX1_LOC_21/Y NAND2X1_LOC_190/A 0.16fF
C4592 INVX1_LOC_599/Y INVX1_LOC_48/Y 0.03fF
C4593 INVX1_LOC_469/Y INVX1_LOC_80/A 0.00fF
C4594 INVX1_LOC_80/A INVX1_LOC_350/Y 0.04fF
C4595 INVX1_LOC_523/A INVX1_LOC_655/A 0.61fF
C4596 NAND2X1_LOC_325/B NAND2X1_LOC_112/a_36_24# 0.00fF
C4597 INVX1_LOC_46/Y INVX1_LOC_489/Y 0.03fF
C4598 INVX1_LOC_617/Y INVX1_LOC_199/Y 0.07fF
C4599 INVX1_LOC_357/A NAND2X1_LOC_451/a_36_24# 0.02fF
C4600 NAND2X1_LOC_45/Y INVX1_LOC_75/Y 0.10fF
C4601 INVX1_LOC_53/Y NAND2X1_LOC_128/A 0.04fF
C4602 NAND2X1_LOC_503/Y INVX1_LOC_600/A 0.25fF
C4603 NAND2X1_LOC_506/a_36_24# INVX1_LOC_396/A 0.02fF
C4604 INVX1_LOC_404/Y INVX1_LOC_41/Y 0.00fF
C4605 INVX1_LOC_17/Y INVX1_LOC_681/Y 0.04fF
C4606 INVX1_LOC_558/Y INVX1_LOC_46/Y 0.05fF
C4607 NAND2X1_LOC_331/A INVX1_LOC_41/Y 0.12fF
C4608 INVX1_LOC_448/A INVX1_LOC_670/A 0.06fF
C4609 INVX1_LOC_411/A INVX1_LOC_98/Y 0.13fF
C4610 INVX1_LOC_503/A INPUT_1 0.01fF
C4611 NAND2X1_LOC_184/Y INVX1_LOC_99/Y 0.15fF
C4612 INVX1_LOC_17/Y INPUT_1 0.13fF
C4613 INVX1_LOC_213/Y NAND2X1_LOC_106/B 0.28fF
C4614 INVX1_LOC_467/Y INVX1_LOC_537/A 0.15fF
C4615 INVX1_LOC_437/A NAND2X1_LOC_563/a_36_24# 0.02fF
C4616 INVX1_LOC_21/Y INVX1_LOC_87/A 0.47fF
C4617 INVX1_LOC_307/A INVX1_LOC_6/Y 1.32fF
C4618 INVX1_LOC_681/A INVX1_LOC_117/Y 0.02fF
C4619 VDD INVX1_LOC_291/Y 0.21fF
C4620 INVX1_LOC_255/Y INVX1_LOC_62/Y 0.03fF
C4621 INVX1_LOC_312/Y NAND2X1_LOC_847/A 0.04fF
C4622 INVX1_LOC_326/A NAND2X1_LOC_397/Y 0.09fF
C4623 NAND2X1_LOC_600/a_36_24# INVX1_LOC_50/Y 0.01fF
C4624 INVX1_LOC_417/Y INVX1_LOC_419/A 0.01fF
C4625 INVX1_LOC_326/Y INVX1_LOC_7/Y 0.08fF
C4626 INVX1_LOC_318/A INVX1_LOC_35/Y 0.01fF
C4627 INVX1_LOC_147/A INVX1_LOC_149/Y 0.08fF
C4628 INVX1_LOC_584/Y INVX1_LOC_479/A 0.02fF
C4629 INPUT_0 NAND2X1_LOC_227/A 0.00fF
C4630 INVX1_LOC_183/A INVX1_LOC_324/Y 0.01fF
C4631 INVX1_LOC_573/Y NAND2X1_LOC_679/B 0.28fF
C4632 INVX1_LOC_51/A INVX1_LOC_634/Y 0.00fF
C4633 INVX1_LOC_31/Y NAND2X1_LOC_673/B 0.11fF
C4634 INVX1_LOC_397/Y INVX1_LOC_35/Y 0.01fF
C4635 INVX1_LOC_513/Y INVX1_LOC_537/A 0.02fF
C4636 INVX1_LOC_197/A INVX1_LOC_653/A 0.06fF
C4637 INVX1_LOC_11/Y NAND2X1_LOC_181/A 0.34fF
C4638 INVX1_LOC_208/A INVX1_LOC_208/Y 0.01fF
C4639 INVX1_LOC_398/A INVX1_LOC_531/Y 0.04fF
C4640 INVX1_LOC_551/A INVX1_LOC_99/Y 0.00fF
C4641 INVX1_LOC_80/A INVX1_LOC_77/A 0.01fF
C4642 NAND2X1_LOC_847/A INVX1_LOC_241/Y 0.04fF
C4643 INVX1_LOC_159/Y INVX1_LOC_66/A 0.00fF
C4644 INVX1_LOC_54/Y INVX1_LOC_611/Y 0.01fF
C4645 NAND2X1_LOC_704/B INVX1_LOC_74/Y 0.01fF
C4646 INVX1_LOC_80/A INVX1_LOC_79/A 0.36fF
C4647 INVX1_LOC_95/A INVX1_LOC_35/Y 0.00fF
C4648 INVX1_LOC_234/Y INVX1_LOC_48/Y 0.06fF
C4649 INVX1_LOC_338/Y NAND2X1_LOC_606/Y 0.18fF
C4650 INVX1_LOC_166/A NAND2X1_LOC_308/A 0.01fF
C4651 INVX1_LOC_579/Y INVX1_LOC_79/A 0.07fF
C4652 NAND2X1_LOC_531/Y INVX1_LOC_46/Y 0.03fF
C4653 INVX1_LOC_292/Y INVX1_LOC_601/Y 0.00fF
C4654 INVX1_LOC_439/Y NAND2X1_LOC_555/B 1.06fF
C4655 INVX1_LOC_376/A INVX1_LOC_50/Y 0.21fF
C4656 INVX1_LOC_117/Y INVX1_LOC_168/Y 0.30fF
C4657 INVX1_LOC_81/Y INVX1_LOC_82/Y 0.97fF
C4658 INVX1_LOC_66/A INVX1_LOC_212/Y 0.02fF
C4659 NAND2X1_LOC_301/B INVX1_LOC_509/A 0.05fF
C4660 INVX1_LOC_513/Y INVX1_LOC_496/Y 0.02fF
C4661 NAND2X1_LOC_355/A INVX1_LOC_639/A 0.04fF
C4662 INVX1_LOC_69/Y INVX1_LOC_77/Y 0.07fF
C4663 INVX1_LOC_95/A INVX1_LOC_620/A 0.03fF
C4664 INVX1_LOC_11/Y INVX1_LOC_79/A 0.67fF
C4665 INVX1_LOC_587/Y INVX1_LOC_26/Y 0.03fF
C4666 NAND2X1_LOC_413/Y NAND2X1_LOC_410/Y 0.07fF
C4667 INVX1_LOC_551/A INVX1_LOC_47/Y -0.00fF
C4668 INVX1_LOC_6/Y INVX1_LOC_482/Y -0.00fF
C4669 INVX1_LOC_99/Y INVX1_LOC_75/Y 4.00fF
C4670 INVX1_LOC_32/Y INVX1_LOC_353/A 0.03fF
C4671 INVX1_LOC_502/A INVX1_LOC_50/Y 0.12fF
C4672 INVX1_LOC_607/Y INVX1_LOC_241/A 0.03fF
C4673 INVX1_LOC_62/Y NAND2X1_LOC_220/a_36_24# 0.00fF
C4674 INVX1_LOC_506/A INVX1_LOC_114/A 0.01fF
C4675 INVX1_LOC_410/Y INVX1_LOC_109/Y 0.06fF
C4676 INVX1_LOC_201/A NAND2X1_LOC_227/A 0.00fF
C4677 INVX1_LOC_59/Y NAND2X1_LOC_231/B 0.01fF
C4678 NAND2X1_LOC_677/Y INVX1_LOC_611/A 0.00fF
C4679 NAND2X1_LOC_846/A INVX1_LOC_655/A 0.04fF
C4680 INVX1_LOC_479/A INVX1_LOC_186/Y 0.34fF
C4681 INVX1_LOC_99/Y NAND2X1_LOC_271/A 0.19fF
C4682 NAND2X1_LOC_697/Y INVX1_LOC_613/A 0.20fF
C4683 INVX1_LOC_652/A INVX1_LOC_63/Y 0.01fF
C4684 INVX1_LOC_285/Y INVX1_LOC_26/Y 0.02fF
C4685 NAND2X1_LOC_720/A INVX1_LOC_91/Y 0.01fF
C4686 INVX1_LOC_49/Y INVX1_LOC_369/Y 0.08fF
C4687 INVX1_LOC_675/A INVX1_LOC_112/Y 0.05fF
C4688 INVX1_LOC_26/Y INVX1_LOC_9/Y 0.08fF
C4689 INVX1_LOC_554/A INVX1_LOC_553/Y 0.04fF
C4690 INVX1_LOC_545/A INVX1_LOC_92/A 0.02fF
C4691 INVX1_LOC_47/Y INVX1_LOC_75/Y 0.07fF
C4692 INVX1_LOC_63/Y INVX1_LOC_11/A 0.29fF
C4693 NAND2X1_LOC_433/Y INVX1_LOC_79/A 0.12fF
C4694 NAND2X1_LOC_528/Y INVX1_LOC_328/Y 0.47fF
C4695 INVX1_LOC_49/Y INVX1_LOC_223/A 0.05fF
C4696 INVX1_LOC_100/Y INVX1_LOC_319/A 0.01fF
C4697 INVX1_LOC_62/Y INVX1_LOC_26/Y 0.10fF
C4698 INVX1_LOC_463/A INVX1_LOC_45/Y 0.15fF
C4699 NAND2X1_LOC_537/A INVX1_LOC_45/Y 0.14fF
C4700 INVX1_LOC_13/Y INVX1_LOC_26/Y 0.05fF
C4701 INVX1_LOC_224/Y INVX1_LOC_400/Y 0.07fF
C4702 INVX1_LOC_100/Y NAND2X1_LOC_843/B 0.14fF
C4703 NAND2X1_LOC_601/Y INVX1_LOC_468/A 0.10fF
C4704 NAND2X1_LOC_844/A INVX1_LOC_26/Y 0.02fF
C4705 INVX1_LOC_133/Y INVX1_LOC_668/A 0.05fF
C4706 INVX1_LOC_529/Y INVX1_LOC_26/Y 0.09fF
C4707 INVX1_LOC_566/A NAND2X1_LOC_590/a_36_24# 0.01fF
C4708 INVX1_LOC_400/Y INVX1_LOC_578/A 0.17fF
C4709 VDD INVX1_LOC_551/Y 2.12fF
C4710 NAND2X1_LOC_475/A NAND2X1_LOC_384/a_36_24# 0.00fF
C4711 INVX1_LOC_450/A NAND2X1_LOC_576/a_36_24# 0.02fF
C4712 INVX1_LOC_79/A INVX1_LOC_231/Y 0.01fF
C4713 INVX1_LOC_355/A INVX1_LOC_45/Y 0.01fF
C4714 INVX1_LOC_160/Y INVX1_LOC_271/Y 0.01fF
C4715 INVX1_LOC_364/A NAND2X1_LOC_458/a_36_24# 0.02fF
C4716 INVX1_LOC_133/Y INVX1_LOC_668/Y 0.01fF
C4717 INVX1_LOC_454/A INVX1_LOC_29/Y 0.01fF
C4718 INVX1_LOC_228/Y INVX1_LOC_551/Y 0.13fF
C4719 INVX1_LOC_441/A INVX1_LOC_634/Y 0.01fF
C4720 INPUT_0 INVX1_LOC_367/A 0.07fF
C4721 NAND2X1_LOC_231/A INVX1_LOC_586/A 0.02fF
C4722 INVX1_LOC_580/Y INVX1_LOC_577/Y 0.17fF
C4723 INVX1_LOC_145/Y INVX1_LOC_616/Y 0.01fF
C4724 INVX1_LOC_206/Y INVX1_LOC_344/Y 0.05fF
C4725 INVX1_LOC_298/Y VDD 0.38fF
C4726 INVX1_LOC_628/Y INVX1_LOC_629/A 0.14fF
C4727 INVX1_LOC_551/Y INVX1_LOC_510/Y 0.10fF
C4728 GATE_366 NAND2X1_LOC_367/a_36_24# 0.00fF
C4729 INVX1_LOC_293/Y INVX1_LOC_51/Y 0.03fF
C4730 INPUT_0 INVX1_LOC_516/A 0.02fF
C4731 INVX1_LOC_482/A INVX1_LOC_235/Y 0.01fF
C4732 NAND2X1_LOC_526/Y INVX1_LOC_387/A 0.00fF
C4733 NAND2X1_LOC_753/a_36_24# NAND2X1_LOC_837/A 0.01fF
C4734 INVX1_LOC_133/Y INVX1_LOC_476/A 0.00fF
C4735 NAND2X1_LOC_66/a_36_24# NAND2X1_LOC_294/Y 0.01fF
C4736 INVX1_LOC_558/A NAND2X1_LOC_413/Y 0.02fF
C4737 INVX1_LOC_290/Y GATE_865 0.01fF
C4738 INVX1_LOC_663/Y INVX1_LOC_445/A 0.01fF
C4739 VDD NAND2X1_LOC_252/Y -0.00fF
C4740 INVX1_LOC_570/Y INVX1_LOC_6/Y 0.01fF
C4741 INVX1_LOC_617/Y INVX1_LOC_53/Y 0.11fF
C4742 INPUT_3 INVX1_LOC_27/A 0.23fF
C4743 INVX1_LOC_492/A INVX1_LOC_570/A 0.03fF
C4744 INVX1_LOC_418/Y INVX1_LOC_442/A 0.03fF
C4745 INVX1_LOC_420/Y INVX1_LOC_46/Y 0.03fF
C4746 INVX1_LOC_20/Y NAND2X1_LOC_147/B 0.03fF
C4747 NAND2X1_LOC_486/B INVX1_LOC_99/Y 0.09fF
C4748 INPUT_0 INVX1_LOC_93/Y 23.24fF
C4749 VDD INVX1_LOC_486/A -0.00fF
C4750 INVX1_LOC_606/Y INVX1_LOC_46/Y 0.01fF
C4751 INVX1_LOC_444/Y INVX1_LOC_218/A 0.00fF
C4752 INVX1_LOC_519/A INVX1_LOC_375/Y 0.08fF
C4753 INVX1_LOC_344/Y INVX1_LOC_686/A -0.01fF
C4754 INVX1_LOC_271/Y NAND2X1_LOC_267/A 0.02fF
C4755 NAND2X1_LOC_249/Y INVX1_LOC_9/Y 0.28fF
C4756 INVX1_LOC_579/Y INVX1_LOC_632/A 0.03fF
C4757 INVX1_LOC_428/A INVX1_LOC_387/Y 0.01fF
C4758 INVX1_LOC_634/A INVX1_LOC_252/Y 0.01fF
C4759 INPUT_0 INVX1_LOC_675/A 0.09fF
C4760 INVX1_LOC_288/A NAND2X1_LOC_718/a_36_24# 0.00fF
C4761 INVX1_LOC_43/Y INVX1_LOC_174/A 0.11fF
C4762 INVX1_LOC_68/Y INVX1_LOC_32/Y 0.13fF
C4763 INVX1_LOC_446/Y NAND2X1_LOC_520/A 0.03fF
C4764 INVX1_LOC_375/A INVX1_LOC_199/Y 0.03fF
C4765 INVX1_LOC_41/Y INVX1_LOC_638/A 0.10fF
C4766 NAND2X1_LOC_332/B INVX1_LOC_670/A 0.05fF
C4767 INVX1_LOC_358/A INVX1_LOC_537/A 0.01fF
C4768 INVX1_LOC_335/Y INVX1_LOC_333/Y 0.12fF
C4769 INVX1_LOC_80/A INVX1_LOC_59/Y 0.04fF
C4770 INVX1_LOC_107/A INVX1_LOC_58/Y 0.00fF
C4771 INVX1_LOC_167/Y INVX1_LOC_117/Y 0.04fF
C4772 INVX1_LOC_367/A NAND2X1_LOC_859/a_36_24# 0.00fF
C4773 INVX1_LOC_381/A INVX1_LOC_281/A 0.04fF
C4774 NAND2X1_LOC_636/B INVX1_LOC_137/Y 0.08fF
C4775 NAND2X1_LOC_545/B NAND2X1_LOC_775/B 0.01fF
C4776 INVX1_LOC_35/Y INVX1_LOC_670/Y 0.07fF
C4777 INVX1_LOC_238/Y NAND2X1_LOC_136/Y 0.00fF
C4778 NAND2X1_LOC_128/a_36_24# INVX1_LOC_6/Y 0.00fF
C4779 INVX1_LOC_298/A INVX1_LOC_59/A 0.02fF
C4780 NAND2X1_LOC_690/Y INVX1_LOC_338/Y 0.16fF
C4781 INVX1_LOC_45/Y NAND2X1_LOC_668/Y 0.15fF
C4782 INVX1_LOC_80/A INVX1_LOC_48/Y 0.13fF
C4783 INVX1_LOC_607/Y INVX1_LOC_669/Y 0.06fF
C4784 INVX1_LOC_11/Y INVX1_LOC_509/Y 0.02fF
C4785 INVX1_LOC_435/A INVX1_LOC_145/Y 0.07fF
C4786 INVX1_LOC_191/A INVX1_LOC_181/Y 0.00fF
C4787 INVX1_LOC_601/A NAND2X1_LOC_234/Y 0.00fF
C4788 INVX1_LOC_54/Y NAND2X1_LOC_677/Y 0.04fF
C4789 VDD NAND2X1_LOC_410/Y 0.01fF
C4790 INVX1_LOC_467/Y INVX1_LOC_676/Y 0.01fF
C4791 INVX1_LOC_166/A INVX1_LOC_134/Y 0.05fF
C4792 INVX1_LOC_437/Y INVX1_LOC_452/A 0.01fF
C4793 INVX1_LOC_418/Y INVX1_LOC_116/Y 0.00fF
C4794 NAND2X1_LOC_775/B INVX1_LOC_98/Y 0.10fF
C4795 INVX1_LOC_679/A NAND2X1_LOC_106/B 0.00fF
C4796 INVX1_LOC_6/Y NAND2X1_LOC_272/a_36_24# 0.00fF
C4797 INVX1_LOC_604/Y INVX1_LOC_208/A 0.05fF
C4798 INVX1_LOC_11/Y INVX1_LOC_59/Y 0.03fF
C4799 INVX1_LOC_159/Y INVX1_LOC_116/Y 0.00fF
C4800 NAND2X1_LOC_307/A NAND2X1_LOC_388/A 0.02fF
C4801 NAND2X1_LOC_475/A INVX1_LOC_75/Y 0.23fF
C4802 INVX1_LOC_32/Y INVX1_LOC_600/A 0.11fF
C4803 INVX1_LOC_291/A INVX1_LOC_95/A 0.04fF
C4804 INVX1_LOC_503/A INVX1_LOC_50/Y 0.01fF
C4805 INVX1_LOC_93/Y NAND2X1_LOC_123/A 0.06fF
C4806 NAND2X1_LOC_317/A INVX1_LOC_479/A 0.05fF
C4807 INVX1_LOC_374/A INVX1_LOC_652/A 0.22fF
C4808 INVX1_LOC_17/Y INVX1_LOC_50/Y 4.15fF
C4809 INVX1_LOC_560/A INVX1_LOC_62/Y 0.11fF
C4810 INVX1_LOC_580/Y INVX1_LOC_26/Y 0.00fF
C4811 NAND2X1_LOC_413/Y INVX1_LOC_46/Y 0.07fF
C4812 NAND2X1_LOC_677/Y INVX1_LOC_611/Y 0.01fF
C4813 INVX1_LOC_581/A INVX1_LOC_476/A 0.08fF
C4814 INVX1_LOC_58/Y INVX1_LOC_492/Y 0.00fF
C4815 VDD INVX1_LOC_634/Y 0.24fF
C4816 NAND2X1_LOC_111/Y INVX1_LOC_134/Y 0.03fF
C4817 INVX1_LOC_545/A INPUT_1 0.01fF
C4818 INVX1_LOC_11/Y NAND2X1_LOC_195/a_36_24# 0.00fF
C4819 INVX1_LOC_372/Y INVX1_LOC_347/Y 0.03fF
C4820 NAND2X1_LOC_391/B INVX1_LOC_242/Y 0.00fF
C4821 INVX1_LOC_11/Y INVX1_LOC_48/Y 7.91fF
C4822 INVX1_LOC_117/Y INVX1_LOC_137/Y 0.14fF
C4823 INVX1_LOC_442/Y NAND2X1_LOC_294/Y 0.11fF
C4824 INVX1_LOC_310/Y INVX1_LOC_204/Y 0.01fF
C4825 INVX1_LOC_17/Y NAND2X1_LOC_389/a_36_24# 0.00fF
C4826 INVX1_LOC_602/A INPUT_5 0.05fF
C4827 INVX1_LOC_49/Y INVX1_LOC_489/Y 0.00fF
C4828 NAND2X1_LOC_595/Y INVX1_LOC_66/A 0.03fF
C4829 NAND2X1_LOC_24/Y INVX1_LOC_183/A 0.19fF
C4830 INVX1_LOC_147/A INVX1_LOC_493/Y 0.01fF
C4831 INVX1_LOC_169/A INVX1_LOC_90/Y 0.03fF
C4832 INVX1_LOC_575/A INVX1_LOC_555/A 0.29fF
C4833 NAND2X1_LOC_720/A NAND2X1_LOC_333/B 0.12fF
C4834 INVX1_LOC_76/Y INVX1_LOC_369/Y 0.05fF
C4835 INVX1_LOC_165/Y INVX1_LOC_479/A 0.01fF
C4836 NAND2X1_LOC_548/B INVX1_LOC_245/A 0.01fF
C4837 INVX1_LOC_681/Y INVX1_LOC_230/Y 0.02fF
C4838 INVX1_LOC_253/Y INVX1_LOC_35/Y 0.13fF
C4839 INVX1_LOC_675/A NAND2X1_LOC_123/A 0.04fF
C4840 INVX1_LOC_58/Y NAND2X1_LOC_72/Y 0.18fF
C4841 INVX1_LOC_566/Y INVX1_LOC_79/A 0.01fF
C4842 NAND2X1_LOC_520/A INVX1_LOC_145/Y 0.01fF
C4843 INVX1_LOC_492/A INVX1_LOC_568/A 0.00fF
C4844 NAND2X1_LOC_174/B INVX1_LOC_561/A 0.10fF
C4845 INPUT_1 INVX1_LOC_230/Y 1.94fF
C4846 INVX1_LOC_419/Y NAND2X1_LOC_388/A 0.21fF
C4847 INVX1_LOC_285/A INVX1_LOC_273/Y 0.00fF
C4848 INVX1_LOC_266/Y INVX1_LOC_479/A 0.08fF
C4849 INVX1_LOC_65/Y NAND2X1_LOC_71/a_36_24# 0.01fF
C4850 NAND2X1_LOC_267/A NAND2X1_LOC_265/a_36_24# 0.02fF
C4851 NAND2X1_LOC_527/Y INVX1_LOC_421/A -0.08fF
C4852 INVX1_LOC_298/A INVX1_LOC_93/Y 0.04fF
C4853 NAND2X1_LOC_591/Y INVX1_LOC_561/A 0.04fF
C4854 INVX1_LOC_54/Y INVX1_LOC_89/Y 0.12fF
C4855 INVX1_LOC_35/Y INVX1_LOC_63/Y 1.03fF
C4856 INVX1_LOC_193/A NAND2X1_LOC_542/A 0.04fF
C4857 NAND2X1_LOC_370/A INVX1_LOC_270/Y 0.05fF
C4858 INVX1_LOC_255/A INVX1_LOC_159/Y 0.01fF
C4859 NAND2X1_LOC_586/Y INVX1_LOC_259/Y 0.00fF
C4860 NAND2X1_LOC_307/B INVX1_LOC_50/Y 0.04fF
C4861 INVX1_LOC_32/Y INVX1_LOC_484/A 0.00fF
C4862 NAND2X1_LOC_147/B INVX1_LOC_655/A 0.02fF
C4863 INVX1_LOC_518/Y INVX1_LOC_670/Y 0.03fF
C4864 INVX1_LOC_364/Y INVX1_LOC_363/A 0.01fF
C4865 INVX1_LOC_432/Y NAND2X1_LOC_558/B 0.06fF
C4866 INVX1_LOC_230/A INVX1_LOC_245/A 0.00fF
C4867 INVX1_LOC_62/Y INVX1_LOC_369/A 0.03fF
C4868 INVX1_LOC_623/Y INVX1_LOC_621/Y 0.15fF
C4869 NAND2X1_LOC_370/A INVX1_LOC_92/A 0.58fF
C4870 INVX1_LOC_69/Y INVX1_LOC_463/Y 0.05fF
C4871 INVX1_LOC_42/Y INVX1_LOC_26/Y 0.04fF
C4872 INVX1_LOC_301/Y INVX1_LOC_665/Y 0.03fF
C4873 INVX1_LOC_257/A INVX1_LOC_89/Y 0.01fF
C4874 INVX1_LOC_675/A INVX1_LOC_498/A 0.07fF
C4875 NAND2X1_LOC_803/a_36_24# INVX1_LOC_6/Y 0.00fF
C4876 NAND2X1_LOC_107/Y NAND2X1_LOC_248/B 0.26fF
C4877 NAND2X1_LOC_285/A INVX1_LOC_58/Y 0.01fF
C4878 NAND2X1_LOC_190/A INVX1_LOC_26/Y 0.06fF
C4879 INVX1_LOC_63/Y INVX1_LOC_620/A 0.03fF
C4880 NAND2X1_LOC_433/Y INVX1_LOC_48/Y 0.24fF
C4881 INVX1_LOC_298/A NAND2X1_LOC_334/B 0.02fF
C4882 INVX1_LOC_63/Y NAND2X1_LOC_253/Y 0.62fF
C4883 INVX1_LOC_670/A INVX1_LOC_242/Y 0.10fF
C4884 INVX1_LOC_134/Y INVX1_LOC_363/A 0.01fF
C4885 INVX1_LOC_300/Y INVX1_LOC_261/Y 0.02fF
C4886 INVX1_LOC_479/A INVX1_LOC_352/A 0.00fF
C4887 INVX1_LOC_58/Y INVX1_LOC_351/Y 0.01fF
C4888 NAND2X1_LOC_309/a_36_24# INVX1_LOC_9/Y 0.00fF
C4889 INVX1_LOC_489/A NAND2X1_LOC_416/B 0.16fF
C4890 INVX1_LOC_361/Y INVX1_LOC_100/Y 0.43fF
C4891 INVX1_LOC_139/Y INVX1_LOC_496/A 0.01fF
C4892 INVX1_LOC_338/A INVX1_LOC_588/A 0.00fF
C4893 INVX1_LOC_11/Y NAND2X1_LOC_629/a_36_24# 0.00fF
C4894 INVX1_LOC_58/Y INVX1_LOC_168/Y 0.46fF
C4895 INVX1_LOC_79/A INVX1_LOC_374/Y 0.01fF
C4896 INVX1_LOC_213/Y NAND2X1_LOC_248/B 0.00fF
C4897 NAND2X1_LOC_165/Y INVX1_LOC_531/Y 0.02fF
C4898 INVX1_LOC_400/A INVX1_LOC_211/A 0.17fF
C4899 INVX1_LOC_335/A INVX1_LOC_479/A 2.08fF
C4900 NAND2X1_LOC_285/A NAND2X1_LOC_342/B 0.03fF
C4901 NAND2X1_LOC_274/B INVX1_LOC_69/Y 0.07fF
C4902 INVX1_LOC_682/A INVX1_LOC_682/Y 0.04fF
C4903 INVX1_LOC_54/Y NAND2X1_LOC_544/B 0.16fF
C4904 INVX1_LOC_399/Y INVX1_LOC_44/Y 0.02fF
C4905 INPUT_0 INVX1_LOC_615/Y 0.01fF
C4906 INVX1_LOC_381/Y INVX1_LOC_443/A 0.11fF
C4907 INVX1_LOC_46/Y INVX1_LOC_645/Y 0.06fF
C4908 INVX1_LOC_211/A NAND2X1_LOC_289/a_36_24# 0.00fF
C4909 VDD INVX1_LOC_596/Y 0.05fF
C4910 INVX1_LOC_261/Y INVX1_LOC_74/Y 0.03fF
C4911 INVX1_LOC_74/A NAND2X1_LOC_95/a_36_24# 0.00fF
C4912 NAND2X1_LOC_558/B NAND2X1_LOC_494/a_36_24# 0.02fF
C4913 INVX1_LOC_257/A NAND2X1_LOC_544/B 0.00fF
C4914 INVX1_LOC_292/Y INVX1_LOC_598/Y -0.00fF
C4915 INVX1_LOC_224/Y NAND2X1_LOC_45/Y 0.96fF
C4916 INVX1_LOC_62/Y NAND2X1_LOC_605/B 0.01fF
C4917 NAND2X1_LOC_528/Y INVX1_LOC_224/A 0.03fF
C4918 VDD INVX1_LOC_416/Y 0.21fF
C4919 INVX1_LOC_49/Y NAND2X1_LOC_832/A 0.02fF
C4920 INVX1_LOC_584/A INVX1_LOC_206/Y 0.08fF
C4921 NAND2X1_LOC_45/Y INVX1_LOC_578/A 0.10fF
C4922 NAND2X1_LOC_249/Y NAND2X1_LOC_371/a_36_24# 0.00fF
C4923 INPUT_0 INVX1_LOC_37/Y 0.09fF
C4924 INPUT_0 INVX1_LOC_395/A 0.25fF
C4925 INVX1_LOC_400/Y INVX1_LOC_206/Y 6.74fF
C4926 NAND2X1_LOC_516/Y INVX1_LOC_395/A 0.10fF
C4927 VDD INVX1_LOC_287/Y 0.39fF
C4928 INVX1_LOC_79/A INVX1_LOC_625/Y 0.16fF
C4929 INVX1_LOC_79/A INVX1_LOC_91/Y 0.03fF
C4930 INVX1_LOC_557/A NAND2X1_LOC_498/Y 0.08fF
C4931 INPUT_6 INPUT_7 1.39fF
C4932 INVX1_LOC_335/Y INVX1_LOC_638/A 0.07fF
C4933 INVX1_LOC_201/Y INVX1_LOC_615/A 0.08fF
C4934 INVX1_LOC_288/Y NAND2X1_LOC_801/A 0.18fF
C4935 INVX1_LOC_442/A NAND2X1_LOC_568/a_36_24# 0.02fF
C4936 INVX1_LOC_395/A INVX1_LOC_586/Y 0.03fF
C4937 INVX1_LOC_228/Y INVX1_LOC_270/A -0.00fF
C4938 INVX1_LOC_53/Y INVX1_LOC_553/Y 0.00fF
C4939 INVX1_LOC_392/Y INVX1_LOC_384/A 0.01fF
C4940 VDD NAND2X1_LOC_755/B 0.25fF
C4941 INVX1_LOC_68/Y NAND2X1_LOC_89/a_36_24# 0.00fF
C4942 INVX1_LOC_400/Y INVX1_LOC_686/A 0.17fF
C4943 INVX1_LOC_561/Y INVX1_LOC_579/Y 0.00fF
C4944 INVX1_LOC_53/Y INVX1_LOC_375/A 0.03fF
C4945 VDD INVX1_LOC_211/Y 0.77fF
C4946 NAND2X1_LOC_513/Y INVX1_LOC_80/A 0.02fF
C4947 INVX1_LOC_53/Y INVX1_LOC_546/A 0.10fF
C4948 NAND2X1_LOC_788/A INVX1_LOC_352/Y 0.10fF
C4949 INPUT_0 INVX1_LOC_284/A 0.09fF
C4950 INVX1_LOC_438/A INVX1_LOC_17/Y 0.08fF
C4951 INVX1_LOC_224/Y INVX1_LOC_99/Y 0.17fF
C4952 VDD NAND2X1_LOC_728/A -0.00fF
C4953 INVX1_LOC_198/A INVX1_LOC_181/A 0.16fF
C4954 INVX1_LOC_20/Y NAND2X1_LOC_391/B 0.01fF
C4955 INVX1_LOC_435/Y NAND2X1_LOC_496/Y 0.23fF
C4956 NAND2X1_LOC_561/a_36_24# NAND2X1_LOC_475/A 0.00fF
C4957 INVX1_LOC_523/A INVX1_LOC_567/Y 0.02fF
C4958 INVX1_LOC_178/A NAND2X1_LOC_749/Y 0.09fF
C4959 INVX1_LOC_607/Y INVX1_LOC_395/A 0.27fF
C4960 INVX1_LOC_201/A INVX1_LOC_395/A 0.07fF
C4961 INVX1_LOC_578/A INVX1_LOC_99/Y 0.03fF
C4962 INVX1_LOC_564/A INVX1_LOC_59/Y 0.00fF
C4963 NAND2X1_LOC_780/B INVX1_LOC_54/Y 0.03fF
C4964 NAND2X1_LOC_331/A NAND2X1_LOC_220/a_36_24# 0.01fF
C4965 INVX1_LOC_552/Y INVX1_LOC_35/Y -0.00fF
C4966 INVX1_LOC_468/Y NAND2X1_LOC_498/Y 0.01fF
C4967 INVX1_LOC_261/Y NAND2X1_LOC_591/B 0.02fF
C4968 INVX1_LOC_28/Y INPUT_2 0.01fF
C4969 VDD INVX1_LOC_46/Y 3.25fF
C4970 NAND2X1_LOC_789/B INVX1_LOC_198/A 0.03fF
C4971 NAND2X1_LOC_148/A INVX1_LOC_133/A 0.02fF
C4972 INVX1_LOC_468/Y INVX1_LOC_570/A 0.01fF
C4973 INVX1_LOC_530/Y NAND2X1_LOC_621/a_36_24# 0.01fF
C4974 INVX1_LOC_392/Y INVX1_LOC_145/Y 0.13fF
C4975 INVX1_LOC_257/Y INVX1_LOC_93/Y 2.27fF
C4976 INVX1_LOC_319/Y INVX1_LOC_48/Y 0.01fF
C4977 INVX1_LOC_442/A INVX1_LOC_352/Y 0.65fF
C4978 NAND2X1_LOC_592/B INVX1_LOC_50/Y 0.02fF
C4979 INPUT_0 INVX1_LOC_31/Y 0.97fF
C4980 INVX1_LOC_298/A INVX1_LOC_395/A 0.01fF
C4981 NAND2X1_LOC_391/B INVX1_LOC_300/A 0.01fF
C4982 NAND2X1_LOC_528/Y INVX1_LOC_109/Y 0.32fF
C4983 INVX1_LOC_224/Y INVX1_LOC_47/Y 0.10fF
C4984 INVX1_LOC_54/Y INVX1_LOC_137/A 0.05fF
C4985 INVX1_LOC_629/A INVX1_LOC_261/Y 0.00fF
C4986 INVX1_LOC_465/Y INVX1_LOC_245/A 0.01fF
C4987 INVX1_LOC_392/A INVX1_LOC_384/A 0.01fF
C4988 INVX1_LOC_393/Y NAND2X1_LOC_181/A 0.54fF
C4989 INVX1_LOC_145/Y INVX1_LOC_59/A 0.02fF
C4990 INVX1_LOC_312/Y INVX1_LOC_683/A 0.07fF
C4991 INVX1_LOC_358/A INVX1_LOC_676/Y 0.11fF
C4992 INVX1_LOC_20/A INVX1_LOC_35/Y 0.09fF
C4993 INVX1_LOC_420/Y INVX1_LOC_49/Y 0.04fF
C4994 INVX1_LOC_257/Y INVX1_LOC_675/A 0.14fF
C4995 INVX1_LOC_584/A NAND2X1_LOC_334/A 0.15fF
C4996 INVX1_LOC_58/Y NAND2X1_LOC_749/Y 0.12fF
C4997 INVX1_LOC_578/A INVX1_LOC_47/Y 0.07fF
C4998 INVX1_LOC_510/Y INVX1_LOC_46/Y 0.07fF
C4999 INVX1_LOC_557/A INVX1_LOC_47/Y 0.08fF
C5000 NAND2X1_LOC_750/Y INVX1_LOC_642/Y 0.01fF
C5001 INVX1_LOC_586/A INVX1_LOC_463/Y 0.10fF
C5002 INVX1_LOC_93/Y INVX1_LOC_384/A 0.07fF
C5003 NAND2X1_LOC_525/Y INVX1_LOC_58/Y 0.44fF
C5004 INVX1_LOC_20/Y INVX1_LOC_670/A 0.07fF
C5005 INVX1_LOC_53/Y INVX1_LOC_662/Y 0.02fF
C5006 INVX1_LOC_492/A INVX1_LOC_136/Y 0.02fF
C5007 INVX1_LOC_45/Y NAND2X1_LOC_449/B 0.01fF
C5008 NAND2X1_LOC_166/a_36_24# INVX1_LOC_160/A 0.00fF
C5009 INVX1_LOC_396/A INVX1_LOC_80/A 0.03fF
C5010 INPUT_0 INVX1_LOC_128/A 0.08fF
C5011 NAND2X1_LOC_143/a_36_24# INVX1_LOC_99/A 0.00fF
C5012 INVX1_LOC_288/A INVX1_LOC_675/A 0.04fF
C5013 INVX1_LOC_84/A NAND2X1_LOC_619/Y 0.01fF
C5014 INVX1_LOC_45/Y INVX1_LOC_480/A 0.01fF
C5015 NAND2X1_LOC_331/A INVX1_LOC_26/Y 0.18fF
C5016 NAND2X1_LOC_531/Y INVX1_LOC_76/Y 0.01fF
C5017 INVX1_LOC_150/Y INVX1_LOC_501/A 0.00fF
C5018 INVX1_LOC_406/Y NAND2X1_LOC_346/B 0.01fF
C5019 NAND2X1_LOC_734/a_36_24# INVX1_LOC_79/A 0.00fF
C5020 INVX1_LOC_363/Y NAND2X1_LOC_464/a_36_24# 0.00fF
C5021 INVX1_LOC_21/Y INVX1_LOC_665/Y 0.03fF
C5022 INVX1_LOC_614/A INVX1_LOC_46/Y 0.23fF
C5023 INVX1_LOC_392/A INVX1_LOC_145/Y 0.00fF
C5024 INVX1_LOC_65/Y INVX1_LOC_223/Y 0.76fF
C5025 NAND2X1_LOC_616/Y INVX1_LOC_50/Y 0.13fF
C5026 NAND2X1_LOC_56/Y INVX1_LOC_32/Y 0.00fF
C5027 INVX1_LOC_682/A INVX1_LOC_51/Y 0.01fF
C5028 INVX1_LOC_193/A NAND2X1_LOC_323/a_36_24# 0.00fF
C5029 INVX1_LOC_116/Y INVX1_LOC_352/Y 0.03fF
C5030 INVX1_LOC_167/Y INVX1_LOC_58/Y 0.01fF
C5031 INVX1_LOC_406/Y NAND2X1_LOC_274/Y 0.10fF
C5032 INVX1_LOC_364/Y INVX1_LOC_301/Y 0.03fF
C5033 INVX1_LOC_603/Y NAND2X1_LOC_387/Y 0.07fF
C5034 INVX1_LOC_273/A INVX1_LOC_399/A 0.02fF
C5035 NAND2X1_LOC_491/a_36_24# INVX1_LOC_9/Y 0.00fF
C5036 INVX1_LOC_106/Y NAND2X1_LOC_142/Y 0.01fF
C5037 INPUT_0 INVX1_LOC_473/Y 0.01fF
C5038 INVX1_LOC_168/A INVX1_LOC_496/A 0.01fF
C5039 INVX1_LOC_557/A INVX1_LOC_119/Y 0.03fF
C5040 INVX1_LOC_432/Y INVX1_LOC_48/Y 0.12fF
C5041 INVX1_LOC_448/A INVX1_LOC_93/Y 0.03fF
C5042 INVX1_LOC_367/Y INVX1_LOC_48/Y 0.03fF
C5043 NAND2X1_LOC_308/a_36_24# INVX1_LOC_98/Y 0.06fF
C5044 INVX1_LOC_93/Y NAND2X1_LOC_612/A 0.07fF
C5045 NAND2X1_LOC_199/a_36_24# INVX1_LOC_63/Y 0.00fF
C5046 INVX1_LOC_662/A INVX1_LOC_133/A 0.06fF
C5047 INVX1_LOC_256/Y INVX1_LOC_63/Y 0.02fF
C5048 INVX1_LOC_586/A NAND2X1_LOC_274/B 0.10fF
C5049 INVX1_LOC_84/A NAND2X1_LOC_618/a_36_24# 0.00fF
C5050 INVX1_LOC_93/Y INVX1_LOC_145/Y 3.06fF
C5051 INVX1_LOC_145/Y INVX1_LOC_283/A 0.07fF
C5052 INVX1_LOC_21/Y NAND2X1_LOC_308/A 0.04fF
C5053 NAND2X1_LOC_13/a_36_24# INVX1_LOC_9/Y 0.00fF
C5054 INVX1_LOC_53/Y INVX1_LOC_646/Y 0.15fF
C5055 INVX1_LOC_628/A INVX1_LOC_261/Y 0.00fF
C5056 INVX1_LOC_481/Y INVX1_LOC_169/Y 0.03fF
C5057 INVX1_LOC_54/Y INVX1_LOC_194/Y 0.55fF
C5058 INVX1_LOC_76/Y NAND2X1_LOC_628/Y 0.01fF
C5059 INVX1_LOC_633/Y INVX1_LOC_338/Y 0.07fF
C5060 INVX1_LOC_661/Y INVX1_LOC_283/A 0.03fF
C5061 INVX1_LOC_183/A NAND2X1_LOC_8/a_36_24# 0.00fF
C5062 INVX1_LOC_191/A INVX1_LOC_26/Y 0.54fF
C5063 INVX1_LOC_17/Y NAND2X1_LOC_63/a_36_24# 0.00fF
C5064 INVX1_LOC_395/A INVX1_LOC_211/A 0.07fF
C5065 NAND2X1_LOC_697/Y INVX1_LOC_555/A 0.06fF
C5066 NAND2X1_LOC_432/Y INVX1_LOC_345/A 0.09fF
C5067 INVX1_LOC_317/A INVX1_LOC_98/Y 0.22fF
C5068 INVX1_LOC_17/Y NAND2X1_LOC_388/A 0.03fF
C5069 NAND2X1_LOC_775/B NAND2X1_LOC_442/a_36_24# 0.00fF
C5070 INVX1_LOC_382/A INVX1_LOC_381/Y 0.15fF
C5071 INVX1_LOC_301/Y INVX1_LOC_134/Y 0.29fF
C5072 INVX1_LOC_586/A INVX1_LOC_148/Y 0.00fF
C5073 INVX1_LOC_340/Y INVX1_LOC_505/Y 0.19fF
C5074 INVX1_LOC_442/A NAND2X1_LOC_438/a_36_24# 0.01fF
C5075 INVX1_LOC_312/Y NAND2X1_LOC_274/B 0.03fF
C5076 NAND2X1_LOC_334/A INVX1_LOC_537/A 0.07fF
C5077 INVX1_LOC_675/A INVX1_LOC_145/Y 0.07fF
C5078 INVX1_LOC_418/Y INVX1_LOC_69/Y 0.01fF
C5079 INVX1_LOC_35/Y NAND2X1_LOC_836/B 0.09fF
C5080 INVX1_LOC_298/A INVX1_LOC_31/Y 0.03fF
C5081 INVX1_LOC_188/Y INVX1_LOC_491/A 0.09fF
C5082 INVX1_LOC_53/Y INVX1_LOC_273/Y 0.00fF
C5083 INVX1_LOC_69/Y INVX1_LOC_159/Y 0.07fF
C5084 INVX1_LOC_214/Y INVX1_LOC_63/Y 0.01fF
C5085 NAND2X1_LOC_141/a_36_24# INVX1_LOC_105/A 0.00fF
C5086 NAND2X1_LOC_403/A INVX1_LOC_183/A 0.02fF
C5087 INVX1_LOC_665/A NAND2X1_LOC_541/B 0.10fF
C5088 INVX1_LOC_137/Y INVX1_LOC_58/Y 0.10fF
C5089 NAND2X1_LOC_427/Y INVX1_LOC_479/A 0.04fF
C5090 INVX1_LOC_49/Y INVX1_LOC_371/A 0.02fF
C5091 INVX1_LOC_62/Y INVX1_LOC_235/Y 0.43fF
C5092 INVX1_LOC_100/Y INVX1_LOC_307/A 0.12fF
C5093 INVX1_LOC_45/Y INVX1_LOC_291/Y 0.01fF
C5094 INVX1_LOC_137/Y NAND2X1_LOC_636/a_36_24# 0.01fF
C5095 INVX1_LOC_356/A NAND2X1_LOC_428/Y 0.00fF
C5096 INVX1_LOC_681/A INVX1_LOC_245/A 0.01fF
C5097 INVX1_LOC_11/Y NAND2X1_LOC_615/Y 0.06fF
C5098 INVX1_LOC_523/A INVX1_LOC_92/A 0.10fF
C5099 INVX1_LOC_556/Y INVX1_LOC_9/Y 0.23fF
C5100 INVX1_LOC_134/Y INVX1_LOC_41/Y 0.43fF
C5101 INVX1_LOC_543/A INVX1_LOC_145/Y 0.00fF
C5102 NAND2X1_LOC_520/B NAND2X1_LOC_271/A 0.04fF
C5103 INVX1_LOC_507/A INVX1_LOC_50/Y 0.01fF
C5104 INVX1_LOC_63/Y INVX1_LOC_118/A 0.01fF
C5105 NAND2X1_LOC_463/a_36_24# INVX1_LOC_41/Y 0.00fF
C5106 INVX1_LOC_638/Y INVX1_LOC_686/Y 0.00fF
C5107 INVX1_LOC_469/Y INVX1_LOC_258/Y 0.02fF
C5108 INVX1_LOC_81/Y INVX1_LOC_9/Y 0.27fF
C5109 INVX1_LOC_54/Y INVX1_LOC_44/Y 0.07fF
C5110 INVX1_LOC_208/A INVX1_LOC_63/Y 0.01fF
C5111 INVX1_LOC_117/Y INVX1_LOC_376/A 0.07fF
C5112 INVX1_LOC_442/Y INVX1_LOC_100/Y 0.05fF
C5113 INVX1_LOC_69/Y INVX1_LOC_340/A 5.89fF
C5114 INVX1_LOC_339/Y INVX1_LOC_46/Y 0.01fF
C5115 INVX1_LOC_35/Y INVX1_LOC_669/A 0.01fF
C5116 NAND2X1_LOC_755/B INVX1_LOC_635/Y 0.04fF
C5117 INVX1_LOC_41/Y INVX1_LOC_235/A 0.02fF
C5118 INVX1_LOC_89/Y INVX1_LOC_501/A 0.03fF
C5119 NAND2X1_LOC_320/Y INVX1_LOC_479/A 0.00fF
C5120 INVX1_LOC_116/Y NAND2X1_LOC_372/Y 0.03fF
C5121 INVX1_LOC_319/A INVX1_LOC_48/Y 0.01fF
C5122 INVX1_LOC_26/Y INVX1_LOC_169/Y 0.07fF
C5123 INVX1_LOC_556/Y INVX1_LOC_62/Y 0.07fF
C5124 INVX1_LOC_117/Y INVX1_LOC_502/A 0.12fF
C5125 INVX1_LOC_671/A INVX1_LOC_100/Y 0.00fF
C5126 INVX1_LOC_361/Y INVX1_LOC_79/A 0.11fF
C5127 INVX1_LOC_518/A INVX1_LOC_66/A 0.03fF
C5128 INVX1_LOC_116/Y NAND2X1_LOC_438/a_36_24# 0.00fF
C5129 INVX1_LOC_223/A INVX1_LOC_7/Y 0.31fF
C5130 INVX1_LOC_32/Y INVX1_LOC_369/Y 0.07fF
C5131 INVX1_LOC_105/Y INVX1_LOC_680/A 0.01fF
C5132 INPUT_5 INVX1_LOC_58/Y 0.45fF
C5133 INVX1_LOC_510/A INVX1_LOC_666/Y 0.00fF
C5134 INVX1_LOC_54/Y INVX1_LOC_347/A 0.01fF
C5135 INVX1_LOC_26/Y INVX1_LOC_182/Y 0.01fF
C5136 INVX1_LOC_261/Y INVX1_LOC_79/A 0.03fF
C5137 INVX1_LOC_59/Y INVX1_LOC_91/Y 0.01fF
C5138 NAND2X1_LOC_415/B NAND2X1_LOC_416/B 0.04fF
C5139 INVX1_LOC_578/Y INVX1_LOC_74/Y 0.04fF
C5140 INVX1_LOC_360/Y INVX1_LOC_634/Y 0.08fF
C5141 INVX1_LOC_48/Y INVX1_LOC_625/Y 0.01fF
C5142 INVX1_LOC_48/Y INVX1_LOC_91/Y 0.03fF
C5143 INVX1_LOC_69/Y INVX1_LOC_468/A 0.03fF
C5144 NAND2X1_LOC_491/Y INVX1_LOC_319/A 0.05fF
C5145 INVX1_LOC_345/Y INVX1_LOC_348/Y 0.01fF
C5146 INVX1_LOC_65/A INVX1_LOC_41/Y 0.00fF
C5147 INVX1_LOC_3/Y INVX1_LOC_454/A 0.08fF
C5148 INVX1_LOC_31/Y INVX1_LOC_211/A 0.08fF
C5149 INVX1_LOC_424/A VDD 0.00fF
C5150 INVX1_LOC_89/Y NAND2X1_LOC_544/B 0.64fF
C5151 INVX1_LOC_49/Y NAND2X1_LOC_488/Y 0.06fF
C5152 INVX1_LOC_479/A INVX1_LOC_199/Y 0.16fF
C5153 INVX1_LOC_531/Y INVX1_LOC_351/A 0.02fF
C5154 INVX1_LOC_153/Y INVX1_LOC_90/Y 0.16fF
C5155 INVX1_LOC_100/Y INVX1_LOC_664/Y 0.00fF
C5156 INVX1_LOC_255/Y INVX1_LOC_638/A 0.02fF
C5157 INVX1_LOC_674/A INVX1_LOC_636/Y 0.05fF
C5158 VDD INVX1_LOC_548/Y 0.21fF
C5159 NAND2X1_LOC_45/Y INVX1_LOC_206/Y 0.15fF
C5160 INVX1_LOC_224/Y NAND2X1_LOC_475/A 0.07fF
C5161 INVX1_LOC_58/Y INVX1_LOC_647/Y 0.01fF
C5162 INVX1_LOC_531/Y INVX1_LOC_90/Y 0.02fF
C5163 INVX1_LOC_12/Y INVX1_LOC_109/Y 0.10fF
C5164 INPUT_0 NAND2X1_LOC_707/a_36_24# 0.00fF
C5165 VDD INVX1_LOC_530/Y 0.29fF
C5166 INVX1_LOC_206/Y INVX1_LOC_36/A 0.01fF
C5167 INVX1_LOC_206/Y NAND2X1_LOC_498/Y 0.07fF
C5168 VDD NAND2X1_LOC_318/A 0.23fF
C5169 INVX1_LOC_427/A INVX1_LOC_217/Y 0.05fF
C5170 VDD INVX1_LOC_268/Y 0.39fF
C5171 INPUT_6 INVX1_LOC_55/Y 0.01fF
C5172 INPUT_0 INVX1_LOC_51/Y 0.24fF
C5173 INVX1_LOC_409/Y NAND2X1_LOC_299/Y 0.02fF
C5174 INVX1_LOC_320/Y INVX1_LOC_321/A 0.14fF
C5175 NAND2X1_LOC_516/Y INVX1_LOC_51/Y 0.00fF
C5176 NAND2X1_LOC_503/B NAND2X1_LOC_785/a_36_24# 0.01fF
C5177 INVX1_LOC_434/Y INVX1_LOC_434/A 0.01fF
C5178 NAND2X1_LOC_704/B NAND2X1_LOC_513/Y 0.19fF
C5179 VDD INVX1_LOC_563/A 0.00fF
C5180 NAND2X1_LOC_498/Y INVX1_LOC_242/A 0.02fF
C5181 NAND2X1_LOC_780/B NAND2X1_LOC_677/Y 0.12fF
C5182 VDD INVX1_LOC_115/A 0.00fF
C5183 INVX1_LOC_143/Y INVX1_LOC_142/A 0.00fF
C5184 VDD INVX1_LOC_363/Y 0.21fF
C5185 INVX1_LOC_422/Y INVX1_LOC_423/A 0.05fF
C5186 INVX1_LOC_374/A INVX1_LOC_256/Y 0.01fF
C5187 INVX1_LOC_307/Y INVX1_LOC_366/Y 0.01fF
C5188 VDD INVX1_LOC_202/Y 1.30fF
C5189 VDD INVX1_LOC_349/Y 0.20fF
C5190 VDD INVX1_LOC_550/Y 0.21fF
C5191 INVX1_LOC_206/Y INVX1_LOC_99/Y 4.84fF
C5192 VDD INVX1_LOC_381/Y 0.21fF
C5193 INVX1_LOC_395/A NAND2X1_LOC_612/A 0.02fF
C5194 INVX1_LOC_114/Y INVX1_LOC_686/A 0.02fF
C5195 INVX1_LOC_404/Y NAND2X1_LOC_275/Y 0.45fF
C5196 NAND2X1_LOC_332/B INVX1_LOC_367/A 0.09fF
C5197 INVX1_LOC_137/A NAND2X1_LOC_677/Y 0.00fF
C5198 VDD INVX1_LOC_550/A 0.00fF
C5199 INVX1_LOC_395/A INVX1_LOC_145/Y 0.19fF
C5200 INVX1_LOC_228/Y INVX1_LOC_202/Y 0.03fF
C5201 INVX1_LOC_442/A INVX1_LOC_67/Y 0.04fF
C5202 INVX1_LOC_603/Y INVX1_LOC_269/A 0.00fF
C5203 INVX1_LOC_445/Y INVX1_LOC_452/A 0.03fF
C5204 INVX1_LOC_450/A INVX1_LOC_442/Y 0.02fF
C5205 NAND2X1_LOC_239/a_36_24# INVX1_LOC_396/A 0.00fF
C5206 NAND2X1_LOC_475/A INVX1_LOC_227/Y 0.01fF
C5207 INVX1_LOC_51/Y NAND2X1_LOC_123/A 0.03fF
C5208 INVX1_LOC_54/Y INVX1_LOC_118/Y 0.05fF
C5209 INVX1_LOC_428/A NAND2X1_LOC_259/A 0.03fF
C5210 VDD INVX1_LOC_387/Y 0.49fF
C5211 INVX1_LOC_438/A INVX1_LOC_230/Y 0.72fF
C5212 INVX1_LOC_393/Y INVX1_LOC_48/Y 0.08fF
C5213 INVX1_LOC_362/Y INVX1_LOC_145/Y 0.03fF
C5214 INVX1_LOC_63/Y INVX1_LOC_220/A 0.08fF
C5215 NAND2X1_LOC_785/a_36_24# INVX1_LOC_273/A 0.01fF
C5216 INVX1_LOC_317/Y INVX1_LOC_98/Y 0.04fF
C5217 INVX1_LOC_80/A INVX1_LOC_634/A 0.01fF
C5218 INVX1_LOC_257/Y INVX1_LOC_31/Y 0.08fF
C5219 INVX1_LOC_396/Y INVX1_LOC_99/Y 0.09fF
C5220 INVX1_LOC_206/Y INVX1_LOC_589/Y 0.01fF
C5221 INVX1_LOC_402/Y INVX1_LOC_20/Y 0.03fF
C5222 NAND2X1_LOC_332/B INVX1_LOC_669/Y 0.05fF
C5223 INVX1_LOC_523/A INPUT_1 0.04fF
C5224 NAND2X1_LOC_124/a_36_24# INVX1_LOC_115/A 0.00fF
C5225 INVX1_LOC_448/A INVX1_LOC_683/Y 0.02fF
C5226 VDD INVX1_LOC_49/Y 1.95fF
C5227 INVX1_LOC_418/Y INVX1_LOC_586/A 0.00fF
C5228 INVX1_LOC_206/Y INVX1_LOC_47/Y 0.38fF
C5229 INVX1_LOC_446/Y INVX1_LOC_31/Y 0.19fF
C5230 INVX1_LOC_586/A INVX1_LOC_159/Y 2.97fF
C5231 INVX1_LOC_26/Y INVX1_LOC_638/A 0.07fF
C5232 INVX1_LOC_206/Y NAND2X1_LOC_557/B 0.04fF
C5233 INVX1_LOC_434/A INVX1_LOC_63/Y 0.02fF
C5234 VDD INVX1_LOC_533/A 0.00fF
C5235 INVX1_LOC_20/Y INVX1_LOC_435/A 0.98fF
C5236 INVX1_LOC_266/Y NAND2X1_LOC_615/B 0.03fF
C5237 NAND2X1_LOC_122/Y INVX1_LOC_50/Y 0.10fF
C5238 INVX1_LOC_686/A INVX1_LOC_99/Y 0.09fF
C5239 VDD INVX1_LOC_642/Y 0.21fF
C5240 INVX1_LOC_21/Y INVX1_LOC_134/Y 0.37fF
C5241 INVX1_LOC_52/Y INVX1_LOC_63/Y 0.10fF
C5242 INVX1_LOC_298/A INVX1_LOC_51/Y 0.03fF
C5243 INVX1_LOC_288/A INVX1_LOC_31/Y 0.07fF
C5244 INVX1_LOC_605/A INVX1_LOC_523/Y 0.04fF
C5245 NAND2X1_LOC_546/a_36_24# NAND2X1_LOC_184/Y 0.00fF
C5246 INVX1_LOC_353/Y INVX1_LOC_440/Y 0.02fF
C5247 INVX1_LOC_84/A INVX1_LOC_35/Y 0.27fF
C5248 INVX1_LOC_523/A NAND2X1_LOC_277/a_36_24# 0.00fF
C5249 INVX1_LOC_395/A NAND2X1_LOC_490/a_36_24# 0.00fF
C5250 INVX1_LOC_435/A NAND2X1_LOC_473/a_36_24# 0.01fF
C5251 NAND2X1_LOC_475/A NAND2X1_LOC_493/a_36_24# 0.00fF
C5252 INVX1_LOC_568/Y INVX1_LOC_136/Y 0.01fF
C5253 INVX1_LOC_11/Y NAND2X1_LOC_710/A 0.11fF
C5254 INVX1_LOC_406/Y INVX1_LOC_439/Y 0.03fF
C5255 INVX1_LOC_93/Y NAND2X1_LOC_332/B 0.42fF
C5256 INVX1_LOC_586/A INVX1_LOC_340/A 0.03fF
C5257 NAND2X1_LOC_307/A INVX1_LOC_251/Y 0.16fF
C5258 INVX1_LOC_384/A INVX1_LOC_31/Y 0.03fF
C5259 NAND2X1_LOC_318/A INVX1_LOC_68/A 0.03fF
C5260 INVX1_LOC_312/Y INVX1_LOC_159/Y 0.03fF
C5261 INVX1_LOC_589/Y INVX1_LOC_396/Y 0.50fF
C5262 INVX1_LOC_115/A INVX1_LOC_116/A 0.14fF
C5263 INVX1_LOC_67/Y INVX1_LOC_116/Y 0.01fF
C5264 INVX1_LOC_9/Y INVX1_LOC_49/A 0.01fF
C5265 INVX1_LOC_99/Y INVX1_LOC_14/A 0.52fF
C5266 VDD INVX1_LOC_210/A -0.00fF
C5267 NAND2X1_LOC_16/a_36_24# INVX1_LOC_6/Y 0.00fF
C5268 INVX1_LOC_173/A NAND2X1_LOC_52/Y 0.05fF
C5269 VDD INVX1_LOC_17/A 0.00fF
C5270 INVX1_LOC_93/Y INVX1_LOC_125/Y 0.51fF
C5271 INVX1_LOC_400/Y INVX1_LOC_376/Y 0.00fF
C5272 INVX1_LOC_206/Y INVX1_LOC_119/Y 0.21fF
C5273 INVX1_LOC_383/A INVX1_LOC_49/Y 0.04fF
C5274 INVX1_LOC_206/Y NAND2X1_LOC_66/Y 0.03fF
C5275 INVX1_LOC_510/Y INVX1_LOC_49/Y 0.07fF
C5276 INVX1_LOC_47/Y INVX1_LOC_242/A 0.07fF
C5277 INPUT_1 INVX1_LOC_519/A 0.05fF
C5278 INVX1_LOC_435/A INVX1_LOC_300/A 0.15fF
C5279 NAND2X1_LOC_723/a_36_24# INVX1_LOC_74/Y 0.01fF
C5280 INVX1_LOC_35/Y NAND2X1_LOC_67/Y 0.01fF
C5281 VDD INVX1_LOC_92/Y 0.44fF
C5282 INVX1_LOC_129/A INVX1_LOC_304/A 0.04fF
C5283 INVX1_LOC_444/Y INVX1_LOC_451/A 0.39fF
C5284 INVX1_LOC_670/A INVX1_LOC_375/Y 0.02fF
C5285 INVX1_LOC_412/A INVX1_LOC_100/Y 0.07fF
C5286 INVX1_LOC_417/Y INVX1_LOC_361/Y 0.07fF
C5287 INVX1_LOC_47/Y INVX1_LOC_686/A 0.08fF
C5288 INVX1_LOC_288/Y INVX1_LOC_259/Y 0.27fF
C5289 NAND2X1_LOC_393/Y INVX1_LOC_50/Y 0.01fF
C5290 INVX1_LOC_55/A INVX1_LOC_56/Y 0.00fF
C5291 INVX1_LOC_81/Y INVX1_LOC_42/Y 0.01fF
C5292 INVX1_LOC_451/A NAND2X1_LOC_578/a_36_24# 0.00fF
C5293 INVX1_LOC_54/Y INVX1_LOC_610/A 0.00fF
C5294 NAND2X1_LOC_140/B INVX1_LOC_670/A 0.20fF
C5295 NAND2X1_LOC_351/a_36_24# INVX1_LOC_292/Y 0.00fF
C5296 NAND2X1_LOC_260/Y INVX1_LOC_283/A 0.01fF
C5297 INVX1_LOC_592/Y INVX1_LOC_53/Y 0.00fF
C5298 INVX1_LOC_635/A NAND2X1_LOC_753/Y 0.02fF
C5299 INVX1_LOC_103/Y INVX1_LOC_363/Y 0.23fF
C5300 INVX1_LOC_54/Y INVX1_LOC_365/A 0.01fF
C5301 INVX1_LOC_17/Y INVX1_LOC_117/Y 0.37fF
C5302 INVX1_LOC_261/Y INVX1_LOC_632/A 0.08fF
C5303 INVX1_LOC_59/Y NAND2X1_LOC_333/B 0.04fF
C5304 INVX1_LOC_31/Y INVX1_LOC_145/Y 4.25fF
C5305 INVX1_LOC_12/Y INVX1_LOC_199/Y 0.04fF
C5306 INVX1_LOC_166/A INVX1_LOC_98/Y 0.03fF
C5307 INVX1_LOC_683/A INVX1_LOC_6/Y 0.02fF
C5308 INVX1_LOC_119/Y INVX1_LOC_242/A 0.03fF
C5309 INVX1_LOC_352/A INVX1_LOC_66/A 0.08fF
C5310 INVX1_LOC_442/Y NAND2X1_LOC_181/A 0.01fF
C5311 NAND2X1_LOC_635/B GATE_865 0.03fF
C5312 INVX1_LOC_25/Y INVX1_LOC_93/A 0.02fF
C5313 INVX1_LOC_48/Y NAND2X1_LOC_333/B 0.07fF
C5314 INVX1_LOC_442/A NAND2X1_LOC_439/a_36_24# 0.01fF
C5315 NAND2X1_LOC_531/Y INVX1_LOC_7/Y 0.44fF
C5316 INVX1_LOC_586/A INVX1_LOC_468/A 0.01fF
C5317 INVX1_LOC_74/Y INVX1_LOC_618/Y 0.14fF
C5318 INVX1_LOC_81/Y INVX1_LOC_87/A 0.08fF
C5319 INVX1_LOC_551/A INVX1_LOC_600/A 0.02fF
C5320 GATE_741 INVX1_LOC_62/Y 0.02fF
C5321 INVX1_LOC_198/A NAND2X1_LOC_235/a_36_24# 0.00fF
C5322 INVX1_LOC_602/Y INVX1_LOC_659/A 0.01fF
C5323 INVX1_LOC_676/Y NAND2X1_LOC_452/a_36_24# 0.00fF
C5324 INVX1_LOC_686/A INVX1_LOC_119/Y 0.01fF
C5325 NAND2X1_LOC_334/A INVX1_LOC_99/Y 0.13fF
C5326 NAND2X1_LOC_336/B INVX1_LOC_100/Y 0.03fF
C5327 NAND2X1_LOC_122/Y NAND2X1_LOC_448/a_36_24# 0.00fF
C5328 INVX1_LOC_69/Y INVX1_LOC_352/Y 0.09fF
C5329 INVX1_LOC_370/Y INVX1_LOC_301/Y 0.01fF
C5330 INVX1_LOC_49/Y INVX1_LOC_509/A 0.00fF
C5331 INVX1_LOC_268/Y INVX1_LOC_635/Y 0.03fF
C5332 INVX1_LOC_51/Y INVX1_LOC_464/Y 0.19fF
C5333 INVX1_LOC_448/A INVX1_LOC_128/A 0.05fF
C5334 NAND2X1_LOC_260/a_36_24# INVX1_LOC_671/Y 0.00fF
C5335 INVX1_LOC_76/Y INVX1_LOC_645/Y 0.01fF
C5336 INVX1_LOC_318/Y INVX1_LOC_41/Y 0.00fF
C5337 NAND2X1_LOC_307/B INVX1_LOC_117/Y 0.09fF
C5338 INVX1_LOC_105/Y INVX1_LOC_66/A 0.88fF
C5339 INVX1_LOC_93/Y NAND2X1_LOC_128/B 0.04fF
C5340 INVX1_LOC_313/Y NAND2X1_LOC_615/Y 0.04fF
C5341 NAND2X1_LOC_628/Y INVX1_LOC_7/Y 0.01fF
C5342 INVX1_LOC_32/Y INVX1_LOC_187/Y 0.39fF
C5343 NAND2X1_LOC_274/B INVX1_LOC_252/A 0.02fF
C5344 INVX1_LOC_617/Y INVX1_LOC_666/Y 0.63fF
C5345 GATE_662 INVX1_LOC_66/A 0.01fF
C5346 INVX1_LOC_41/Y INVX1_LOC_16/Y 0.01fF
C5347 NAND2X1_LOC_555/B INVX1_LOC_444/A 0.13fF
C5348 INVX1_LOC_53/Y INVX1_LOC_479/A 0.31fF
C5349 INVX1_LOC_626/A INVX1_LOC_614/Y 0.00fF
C5350 INVX1_LOC_435/A NAND2X1_LOC_269/B 0.02fF
C5351 INVX1_LOC_328/Y INVX1_LOC_328/A 0.16fF
C5352 INVX1_LOC_386/A NAND2X1_LOC_482/Y 0.03fF
C5353 INVX1_LOC_99/Y NAND2X1_LOC_609/B 0.00fF
C5354 INVX1_LOC_43/Y INVX1_LOC_190/A 0.01fF
C5355 INVX1_LOC_47/Y NAND2X1_LOC_334/A 0.10fF
C5356 INVX1_LOC_89/Y INVX1_LOC_44/Y 0.05fF
C5357 INVX1_LOC_58/Y NAND2X1_LOC_342/A 0.01fF
C5358 INVX1_LOC_93/Y INVX1_LOC_242/Y 0.07fF
C5359 INVX1_LOC_116/Y NAND2X1_LOC_439/a_36_24# 0.01fF
C5360 INVX1_LOC_378/Y INVX1_LOC_63/Y 0.11fF
C5361 NAND2X1_LOC_333/A INVX1_LOC_272/A 0.01fF
C5362 VDD INVX1_LOC_297/Y 0.49fF
C5363 NAND2X1_LOC_274/B INVX1_LOC_6/Y 0.05fF
C5364 INVX1_LOC_210/A NAND2X1_LOC_243/A 0.20fF
C5365 INVX1_LOC_192/Y INVX1_LOC_109/Y 0.01fF
C5366 NAND2X1_LOC_606/Y INVX1_LOC_588/A 0.02fF
C5367 INVX1_LOC_63/Y INVX1_LOC_223/Y 0.07fF
C5368 NAND2X1_LOC_836/B INVX1_LOC_657/A 0.01fF
C5369 INVX1_LOC_502/A NAND2X1_LOC_271/a_36_24# 0.01fF
C5370 NAND2X1_LOC_334/A INVX1_LOC_119/Y 0.03fF
C5371 INVX1_LOC_254/A INVX1_LOC_211/A 0.02fF
C5372 INVX1_LOC_390/A INVX1_LOC_242/Y 0.00fF
C5373 INVX1_LOC_69/Y INVX1_LOC_280/A 0.03fF
C5374 INVX1_LOC_69/Y NAND2X1_LOC_372/Y 0.03fF
C5375 INVX1_LOC_224/Y NAND2X1_LOC_543/B 0.31fF
C5376 VDD INVX1_LOC_158/A -0.00fF
C5377 INVX1_LOC_32/Y INVX1_LOC_443/A 0.10fF
C5378 INVX1_LOC_49/Y INVX1_LOC_635/Y 0.05fF
C5379 VDD NAND2X1_LOC_764/Y 0.01fF
C5380 NAND2X1_LOC_543/B INVX1_LOC_578/A 0.02fF
C5381 INVX1_LOC_206/Y NAND2X1_LOC_475/A 0.09fF
C5382 INVX1_LOC_273/A INVX1_LOC_275/A 0.07fF
C5383 INVX1_LOC_199/Y INVX1_LOC_212/A 0.01fF
C5384 INVX1_LOC_247/Y INVX1_LOC_280/A 0.10fF
C5385 INVX1_LOC_41/Y INVX1_LOC_90/Y 0.10fF
C5386 VDD INVX1_LOC_250/A -0.00fF
C5387 VDD NAND2X1_LOC_498/B 0.31fF
C5388 INVX1_LOC_241/A INVX1_LOC_655/A 0.05fF
C5389 NAND2X1_LOC_595/a_36_24# INVX1_LOC_362/Y 0.01fF
C5390 INVX1_LOC_320/Y INVX1_LOC_410/Y 0.02fF
C5391 VDD INVX1_LOC_76/Y 4.25fF
C5392 INVX1_LOC_257/Y INVX1_LOC_51/Y 0.09fF
C5393 NAND2X1_LOC_544/B INVX1_LOC_347/A 0.05fF
C5394 INVX1_LOC_425/A INVX1_LOC_193/Y 0.02fF
C5395 INVX1_LOC_446/Y INVX1_LOC_51/Y 0.04fF
C5396 INVX1_LOC_266/A INVX1_LOC_257/Y 0.03fF
C5397 INPUT_0 NAND2X1_LOC_13/Y 0.03fF
C5398 INVX1_LOC_228/Y INVX1_LOC_76/Y 0.09fF
C5399 INVX1_LOC_404/Y INVX1_LOC_235/Y 0.20fF
C5400 INVX1_LOC_288/A INVX1_LOC_51/Y 0.07fF
C5401 INVX1_LOC_426/A INVX1_LOC_145/Y 0.00fF
C5402 NAND2X1_LOC_163/B INVX1_LOC_586/A 0.02fF
C5403 NAND2X1_LOC_583/a_36_24# INVX1_LOC_99/Y 0.00fF
C5404 INVX1_LOC_463/A NAND2X1_LOC_686/a_36_24# 0.00fF
C5405 INVX1_LOC_66/A INVX1_LOC_109/Y 0.51fF
C5406 NAND2X1_LOC_88/B INVX1_LOC_395/A 0.16fF
C5407 VDD INVX1_LOC_386/Y 0.43fF
C5408 INVX1_LOC_384/A INVX1_LOC_51/Y 0.07fF
C5409 NAND2X1_LOC_788/A INVX1_LOC_352/A 0.05fF
C5410 INVX1_LOC_287/Y INVX1_LOC_45/Y 0.01fF
C5411 INVX1_LOC_563/Y INVX1_LOC_635/A 0.06fF
C5412 VDD INVX1_LOC_559/A -0.00fF
C5413 INVX1_LOC_296/A INVX1_LOC_109/Y 0.01fF
C5414 INVX1_LOC_542/A NAND2X1_LOC_685/A 0.01fF
C5415 VDD INVX1_LOC_29/A 0.00fF
C5416 NAND2X1_LOC_750/Y INVX1_LOC_228/A 0.01fF
C5417 INVX1_LOC_459/Y INVX1_LOC_372/Y 0.00fF
C5418 INVX1_LOC_255/Y INVX1_LOC_134/Y 0.00fF
C5419 INVX1_LOC_206/Y INVX1_LOC_25/Y 0.37fF
C5420 INVX1_LOC_21/Y NAND2X1_LOC_110/a_36_24# 0.01fF
C5421 INVX1_LOC_428/Y INVX1_LOC_217/Y 0.49fF
C5422 INVX1_LOC_625/A INVX1_LOC_97/A 0.02fF
C5423 INVX1_LOC_287/A INVX1_LOC_271/A 0.01fF
C5424 INVX1_LOC_301/A INVX1_LOC_93/Y 0.10fF
C5425 INVX1_LOC_542/A NAND2X1_LOC_685/a_36_24# 0.00fF
C5426 VDD NAND2X1_LOC_503/Y 0.16fF
C5427 INVX1_LOC_554/A INVX1_LOC_66/A 0.10fF
C5428 INVX1_LOC_20/Y INVX1_LOC_367/A 0.14fF
C5429 INVX1_LOC_397/A INVX1_LOC_99/Y 0.01fF
C5430 INVX1_LOC_607/Y NAND2X1_LOC_108/Y 0.04fF
C5431 INVX1_LOC_45/Y NAND2X1_LOC_755/B 0.03fF
C5432 INVX1_LOC_445/Y INVX1_LOC_282/A 0.00fF
C5433 INVX1_LOC_206/Y INVX1_LOC_153/A 0.02fF
C5434 INVX1_LOC_99/Y INVX1_LOC_94/A 0.00fF
C5435 NAND2X1_LOC_176/Y INVX1_LOC_89/Y 0.18fF
C5436 INVX1_LOC_51/Y INVX1_LOC_145/Y 0.17fF
C5437 INVX1_LOC_76/Y INVX1_LOC_116/A 0.03fF
C5438 INVX1_LOC_510/Y NAND2X1_LOC_446/a_36_24# 0.00fF
C5439 NAND2X1_LOC_241/B INVX1_LOC_32/Y 0.04fF
C5440 NAND2X1_LOC_592/B INVX1_LOC_117/Y 0.08fF
C5441 INVX1_LOC_65/Y NAND2X1_LOC_775/B 0.00fF
C5442 INVX1_LOC_586/A INVX1_LOC_352/Y 0.00fF
C5443 INVX1_LOC_84/A INVX1_LOC_531/A 0.01fF
C5444 INVX1_LOC_206/Y INVX1_LOC_96/A 0.01fF
C5445 INVX1_LOC_561/Y INVX1_LOC_261/Y 0.00fF
C5446 INVX1_LOC_93/Y INVX1_LOC_533/Y 0.03fF
C5447 INVX1_LOC_185/Y INVX1_LOC_46/Y 0.02fF
C5448 INVX1_LOC_45/Y INVX1_LOC_46/Y 0.07fF
C5449 INVX1_LOC_335/Y INVX1_LOC_455/Y 0.02fF
C5450 INPUT_3 INVX1_LOC_211/Y 0.02fF
C5451 INVX1_LOC_367/Y NAND2X1_LOC_541/B 0.12fF
C5452 NAND2X1_LOC_370/A NAND2X1_LOC_388/A 0.00fF
C5453 NAND2X1_LOC_451/a_36_24# INVX1_LOC_495/A 0.00fF
C5454 NAND2X1_LOC_403/A INVX1_LOC_324/Y 0.00fF
C5455 NAND2X1_LOC_498/Y NAND2X1_LOC_542/A 0.07fF
C5456 INVX1_LOC_396/Y INVX1_LOC_153/A 0.02fF
C5457 INVX1_LOC_54/Y INPUT_2 0.04fF
C5458 NAND2X1_LOC_677/Y INVX1_LOC_610/A 0.01fF
C5459 INVX1_LOC_159/Y INVX1_LOC_486/Y 0.16fF
C5460 INVX1_LOC_38/A INVX1_LOC_6/Y 0.15fF
C5461 INVX1_LOC_20/Y INVX1_LOC_93/Y 0.35fF
C5462 NAND2X1_LOC_39/Y INPUT_1 0.04fF
C5463 INVX1_LOC_224/Y INVX1_LOC_353/A 0.13fF
C5464 INVX1_LOC_111/A INVX1_LOC_497/Y 0.10fF
C5465 INVX1_LOC_434/A INVX1_LOC_430/A 0.13fF
C5466 INVX1_LOC_44/A INVX1_LOC_7/Y 0.01fF
C5467 NAND2X1_LOC_156/Y INVX1_LOC_186/A 0.18fF
C5468 INPUT_3 INVX1_LOC_46/Y 8.55fF
C5469 INVX1_LOC_298/A NAND2X1_LOC_668/a_36_24# 0.00fF
C5470 INVX1_LOC_318/Y NAND2X1_LOC_267/A 0.05fF
C5471 NAND2X1_LOC_498/Y INVX1_LOC_376/Y 2.05fF
C5472 INVX1_LOC_360/Y INVX1_LOC_115/A 0.01fF
C5473 VDD INVX1_LOC_184/Y 0.21fF
C5474 INVX1_LOC_395/A INVX1_LOC_242/Y 0.99fF
C5475 INVX1_LOC_166/A INVX1_LOC_596/A 0.03fF
C5476 INVX1_LOC_519/A INVX1_LOC_50/Y 0.05fF
C5477 NAND2X1_LOC_363/a_36_24# INVX1_LOC_50/Y 0.00fF
C5478 INVX1_LOC_53/Y INVX1_LOC_138/Y 0.01fF
C5479 INVX1_LOC_570/A INVX1_LOC_376/Y 0.09fF
C5480 NAND2X1_LOC_789/a_36_24# INVX1_LOC_198/A 0.00fF
C5481 INVX1_LOC_126/Y INVX1_LOC_66/A 0.39fF
C5482 INVX1_LOC_50/Y NAND2X1_LOC_296/Y 0.02fF
C5483 INVX1_LOC_117/Y NAND2X1_LOC_616/Y 0.46fF
C5484 INVX1_LOC_575/A INVX1_LOC_556/Y 0.01fF
C5485 INVX1_LOC_145/Y INVX1_LOC_40/Y 0.09fF
C5486 NAND2X1_LOC_333/A INVX1_LOC_53/Y 0.11fF
C5487 NAND2X1_LOC_521/Y INVX1_LOC_53/Y 0.02fF
C5488 NAND2X1_LOC_391/A INVX1_LOC_89/Y 0.03fF
C5489 INVX1_LOC_20/Y INVX1_LOC_675/A 0.07fF
C5490 NAND2X1_LOC_467/A INVX1_LOC_338/Y 0.00fF
C5491 INVX1_LOC_442/Y INVX1_LOC_48/Y 0.08fF
C5492 INVX1_LOC_588/Y INVX1_LOC_504/A 0.04fF
C5493 NAND2X1_LOC_818/a_36_24# INVX1_LOC_66/A 0.00fF
C5494 NAND2X1_LOC_820/A INVX1_LOC_212/Y 0.01fF
C5495 INVX1_LOC_54/Y INVX1_LOC_252/Y 0.03fF
C5496 NAND2X1_LOC_662/a_36_24# INVX1_LOC_508/A 0.00fF
C5497 NAND2X1_LOC_513/Y NAND2X1_LOC_413/a_36_24# 0.00fF
C5498 INVX1_LOC_79/A INVX1_LOC_618/Y 0.01fF
C5499 INVX1_LOC_193/A INVX1_LOC_304/A 0.00fF
C5500 INVX1_LOC_254/A INVX1_LOC_145/Y 0.01fF
C5501 INVX1_LOC_382/A INVX1_LOC_7/Y 0.03fF
C5502 INVX1_LOC_20/Y INVX1_LOC_390/A 0.03fF
C5503 INVX1_LOC_300/A INVX1_LOC_93/Y 0.07fF
C5504 NAND2X1_LOC_606/Y NAND2X1_LOC_646/A 0.03fF
C5505 INVX1_LOC_46/Y NAND2X1_LOC_376/Y 0.01fF
C5506 INVX1_LOC_449/A INVX1_LOC_69/Y 0.07fF
C5507 INVX1_LOC_544/A INVX1_LOC_105/Y 0.01fF
C5508 NAND2X1_LOC_339/a_36_24# NAND2X1_LOC_786/B 0.00fF
C5509 INVX1_LOC_53/Y INVX1_LOC_170/A 0.01fF
C5510 INVX1_LOC_411/A NAND2X1_LOC_538/a_36_24# 0.00fF
C5511 INVX1_LOC_117/Y INVX1_LOC_108/Y 0.03fF
C5512 INVX1_LOC_89/Y NAND2X1_LOC_418/Y 0.21fF
C5513 INVX1_LOC_410/Y INVX1_LOC_666/Y 0.10fF
C5514 NAND2X1_LOC_376/a_36_24# INVX1_LOC_183/A 0.01fF
C5515 INVX1_LOC_93/Y INVX1_LOC_197/Y 0.02fF
C5516 NAND2X1_LOC_755/B NAND2X1_LOC_837/A 0.21fF
C5517 INVX1_LOC_578/Y INVX1_LOC_48/Y 0.03fF
C5518 INVX1_LOC_586/A INVX1_LOC_280/A 0.06fF
C5519 INVX1_LOC_172/A INVX1_LOC_328/A 0.02fF
C5520 NAND2X1_LOC_307/A INVX1_LOC_245/A 0.01fF
C5521 NAND2X1_LOC_336/B NAND2X1_LOC_558/B 0.00fF
C5522 INVX1_LOC_548/A NAND2X1_LOC_128/B 0.01fF
C5523 INVX1_LOC_586/A NAND2X1_LOC_372/Y 0.00fF
C5524 INVX1_LOC_17/Y INVX1_LOC_58/Y 4.99fF
C5525 INVX1_LOC_134/Y INVX1_LOC_26/Y 0.18fF
C5526 INVX1_LOC_117/Y INVX1_LOC_230/Y 2.57fF
C5527 INVX1_LOC_134/Y INVX1_LOC_128/Y 0.02fF
C5528 NAND2X1_LOC_79/B INVX1_LOC_79/Y 0.06fF
C5529 INVX1_LOC_209/A INVX1_LOC_69/Y 0.03fF
C5530 INVX1_LOC_411/Y INVX1_LOC_98/Y 0.14fF
C5531 NAND2X1_LOC_336/B INVX1_LOC_79/A 1.56fF
C5532 NAND2X1_LOC_463/a_36_24# INVX1_LOC_26/Y 0.01fF
C5533 INVX1_LOC_188/Y INVX1_LOC_114/A 0.03fF
C5534 INVX1_LOC_532/Y INVX1_LOC_48/Y 0.01fF
C5535 INVX1_LOC_300/A INVX1_LOC_390/A 0.01fF
C5536 INVX1_LOC_199/Y NAND2X1_LOC_615/B 0.05fF
C5537 INVX1_LOC_63/Y NAND2X1_LOC_606/Y 0.05fF
C5538 INVX1_LOC_44/Y INVX1_LOC_194/Y 0.10fF
C5539 INVX1_LOC_105/A INVX1_LOC_49/Y 0.12fF
C5540 INVX1_LOC_26/Y NAND2X1_LOC_241/a_36_24# 0.00fF
C5541 NAND2X1_LOC_13/Y INVX1_LOC_211/A 0.02fF
C5542 INVX1_LOC_21/Y INVX1_LOC_90/Y 0.10fF
C5543 INVX1_LOC_145/Y INVX1_LOC_204/A 0.01fF
C5544 INVX1_LOC_619/A INVX1_LOC_210/A 0.05fF
C5545 INVX1_LOC_304/Y INVX1_LOC_9/Y 0.14fF
C5546 NAND2X1_LOC_276/A INVX1_LOC_46/Y 0.02fF
C5547 INVX1_LOC_117/Y INVX1_LOC_507/A 0.04fF
C5548 INVX1_LOC_366/A INVX1_LOC_620/Y 0.00fF
C5549 INVX1_LOC_298/A NAND2X1_LOC_668/Y 0.01fF
C5550 INVX1_LOC_602/A INVX1_LOC_598/Y 0.14fF
C5551 NAND2X1_LOC_318/B INVX1_LOC_531/Y 0.01fF
C5552 INVX1_LOC_555/A INVX1_LOC_476/A 0.17fF
C5553 INVX1_LOC_685/Y INVX1_LOC_632/Y 0.12fF
C5554 INVX1_LOC_47/Y NAND2X1_LOC_542/A 0.07fF
C5555 INVX1_LOC_199/Y INVX1_LOC_66/A 0.16fF
C5556 NAND2X1_LOC_683/a_36_24# INVX1_LOC_513/A 0.00fF
C5557 INVX1_LOC_579/A NAND2X1_LOC_448/a_36_24# 0.00fF
C5558 INVX1_LOC_634/A INVX1_LOC_625/Y 0.00fF
C5559 INVX1_LOC_424/Y INVX1_LOC_443/A 0.05fF
C5560 INVX1_LOC_89/A INVX1_LOC_46/Y 0.07fF
C5561 INVX1_LOC_569/Y INVX1_LOC_6/Y 0.15fF
C5562 NAND2X1_LOC_307/B INVX1_LOC_58/Y 0.52fF
C5563 INVX1_LOC_41/Y INVX1_LOC_98/Y 0.17fF
C5564 INVX1_LOC_35/Y NAND2X1_LOC_409/Y 0.01fF
C5565 INVX1_LOC_69/Y INVX1_LOC_347/Y 0.03fF
C5566 INVX1_LOC_53/Y INVX1_LOC_212/A 0.08fF
C5567 VDD INVX1_LOC_423/Y 0.14fF
C5568 VDD INVX1_LOC_192/A -0.00fF
C5569 INVX1_LOC_31/Y INVX1_LOC_242/Y 0.07fF
C5570 INVX1_LOC_35/Y INVX1_LOC_135/Y 0.02fF
C5571 INVX1_LOC_655/A INVX1_LOC_283/A 0.02fF
C5572 INVX1_LOC_211/A NAND2X1_LOC_72/a_36_24# 0.01fF
C5573 INVX1_LOC_304/Y INVX1_LOC_62/Y 0.02fF
C5574 INVX1_LOC_93/Y NAND2X1_LOC_269/B 0.08fF
C5575 INVX1_LOC_213/Y INVX1_LOC_479/A 0.11fF
C5576 INVX1_LOC_376/A NAND2X1_LOC_440/A 0.04fF
C5577 INVX1_LOC_31/Y INVX1_LOC_487/A 0.02fF
C5578 INVX1_LOC_62/Y NAND2X1_LOC_444/A 0.01fF
C5579 INVX1_LOC_32/Y NAND2X1_LOC_488/Y 0.01fF
C5580 NAND2X1_LOC_542/A INVX1_LOC_119/Y 0.03fF
C5581 INVX1_LOC_183/A INVX1_LOC_9/Y 0.07fF
C5582 INVX1_LOC_446/A INVX1_LOC_447/A 0.23fF
C5583 VDD NAND2X1_LOC_770/A -0.00fF
C5584 INVX1_LOC_389/Y INVX1_LOC_9/Y 0.10fF
C5585 INVX1_LOC_41/Y INVX1_LOC_497/A 0.03fF
C5586 INVX1_LOC_119/Y INVX1_LOC_376/Y 0.06fF
C5587 NAND2X1_LOC_754/a_36_24# INVX1_LOC_206/Y 0.01fF
C5588 INVX1_LOC_643/Y INVX1_LOC_655/A 0.04fF
C5589 INVX1_LOC_41/Y INVX1_LOC_338/Y 0.13fF
C5590 INVX1_LOC_6/Y INVX1_LOC_39/Y 0.01fF
C5591 NAND2X1_LOC_543/B INVX1_LOC_206/Y 0.42fF
C5592 INVX1_LOC_74/Y INVX1_LOC_77/Y 0.01fF
C5593 INVX1_LOC_484/A NAND2X1_LOC_619/a_36_24# 0.00fF
C5594 INVX1_LOC_301/A INVX1_LOC_395/A 0.08fF
C5595 INVX1_LOC_667/Y INVX1_LOC_669/A 0.00fF
C5596 INVX1_LOC_361/A INVX1_LOC_211/A 0.02fF
C5597 NAND2X1_LOC_832/a_36_24# NAND2X1_LOC_123/B 0.01fF
C5598 INVX1_LOC_26/Y NAND2X1_LOC_791/a_36_24# 0.00fF
C5599 INVX1_LOC_183/A INVX1_LOC_13/Y 0.00fF
C5600 INVX1_LOC_6/Y INVX1_LOC_620/Y 0.00fF
C5601 INVX1_LOC_659/A INVX1_LOC_658/Y 0.09fF
C5602 INVX1_LOC_317/Y NAND2X1_LOC_76/B 0.03fF
C5603 INVX1_LOC_653/A INVX1_LOC_479/A 0.01fF
C5604 INVX1_LOC_616/A INVX1_LOC_180/Y -0.02fF
C5605 INVX1_LOC_85/Y NAND2X1_LOC_205/a_36_24# 0.00fF
C5606 INVX1_LOC_32/A INVX1_LOC_45/Y 0.01fF
C5607 INVX1_LOC_454/A INVX1_LOC_340/Y 0.15fF
C5608 NAND2X1_LOC_249/Y NAND2X1_LOC_692/a_36_24# 0.01fF
C5609 INVX1_LOC_116/Y INVX1_LOC_109/Y 0.03fF
C5610 INVX1_LOC_276/A VDD 0.20fF
C5611 INVX1_LOC_544/A INVX1_LOC_109/Y 0.00fF
C5612 INVX1_LOC_65/Y INVX1_LOC_97/A 0.11fF
C5613 INVX1_LOC_68/Y INVX1_LOC_224/Y 0.03fF
C5614 NAND2X1_LOC_543/B INVX1_LOC_686/A 0.00fF
C5615 NAND2X1_LOC_498/Y INVX1_LOC_253/A 0.01fF
C5616 INVX1_LOC_584/Y INVX1_LOC_586/A 0.02fF
C5617 NAND2X1_LOC_750/Y INVX1_LOC_229/Y 0.01fF
C5618 INVX1_LOC_20/Y INVX1_LOC_395/A 0.51fF
C5619 INVX1_LOC_468/Y INVX1_LOC_409/Y 0.03fF
C5620 VDD NAND2X1_LOC_399/B 0.01fF
C5621 INVX1_LOC_224/Y INVX1_LOC_250/Y 0.04fF
C5622 INVX1_LOC_463/A INVX1_LOC_145/Y 0.07fF
C5623 INVX1_LOC_279/Y INVX1_LOC_452/A 0.01fF
C5624 INVX1_LOC_259/Y NAND2X1_LOC_801/A 0.07fF
C5625 NAND2X1_LOC_332/B INVX1_LOC_51/Y 0.08fF
C5626 VDD INVX1_LOC_7/Y 0.84fF
C5627 NAND2X1_LOC_318/A INVX1_LOC_45/Y 0.43fF
C5628 INVX1_LOC_438/A NAND2X1_LOC_296/Y 0.02fF
C5629 INVX1_LOC_512/Y NAND2X1_LOC_685/B 0.05fF
C5630 VDD INVX1_LOC_228/A -0.00fF
C5631 NAND2X1_LOC_537/A INVX1_LOC_145/Y 0.05fF
C5632 INVX1_LOC_206/Y NAND2X1_LOC_638/A 0.03fF
C5633 VDD INVX1_LOC_256/A -0.00fF
C5634 NAND2X1_LOC_780/B INVX1_LOC_610/A 0.02fF
C5635 INPUT_3 INVX1_LOC_530/Y 0.22fF
C5636 INVX1_LOC_523/A NAND2X1_LOC_513/A 0.06fF
C5637 INVX1_LOC_266/A NAND2X1_LOC_332/B 0.01fF
C5638 INVX1_LOC_578/A NAND2X1_LOC_302/A 0.04fF
C5639 NAND2X1_LOC_7/Y INVX1_LOC_31/Y 0.06fF
C5640 INVX1_LOC_417/Y INVX1_LOC_412/A 0.02fF
C5641 VDD INVX1_LOC_345/Y 0.21fF
C5642 NAND2X1_LOC_475/A INVX1_LOC_432/A 0.02fF
C5643 INVX1_LOC_206/Y INVX1_LOC_505/A 0.00fF
C5644 INVX1_LOC_563/A INVX1_LOC_45/Y 0.01fF
C5645 NAND2X1_LOC_669/Y INVX1_LOC_586/A 0.03fF
C5646 INVX1_LOC_301/A INVX1_LOC_31/Y 0.01fF
C5647 INVX1_LOC_449/A INVX1_LOC_586/A 0.07fF
C5648 INVX1_LOC_395/A INVX1_LOC_197/Y 0.07fF
C5649 VDD INVX1_LOC_32/Y 3.21fF
C5650 NAND2X1_LOC_108/Y INVX1_LOC_145/Y 0.01fF
C5651 INVX1_LOC_45/Y INVX1_LOC_115/A 0.07fF
C5652 NAND2X1_LOC_383/Y INVX1_LOC_12/Y 0.03fF
C5653 INVX1_LOC_412/Y NAND2X1_LOC_123/a_36_24# 0.00fF
C5654 NAND2X1_LOC_140/a_36_24# INVX1_LOC_105/A 0.00fF
C5655 INVX1_LOC_202/Y INVX1_LOC_45/Y 0.00fF
C5656 INVX1_LOC_228/Y INVX1_LOC_32/Y 0.02fF
C5657 NAND2X1_LOC_731/a_36_24# INVX1_LOC_6/Y 0.00fF
C5658 VDD NAND2X1_LOC_286/A -0.00fF
C5659 INVX1_LOC_51/Y INVX1_LOC_440/A 0.01fF
C5660 INVX1_LOC_121/Y INVX1_LOC_47/Y 0.02fF
C5661 INVX1_LOC_360/Y INVX1_LOC_76/Y 0.07fF
C5662 INVX1_LOC_428/A NAND2X1_LOC_184/Y 0.03fF
C5663 INVX1_LOC_686/A INVX1_LOC_469/A 0.04fF
C5664 INVX1_LOC_369/A NAND2X1_LOC_463/a_36_24# 0.02fF
C5665 INVX1_LOC_417/Y NAND2X1_LOC_336/B 0.29fF
C5666 INVX1_LOC_421/Y NAND2X1_LOC_346/B 0.01fF
C5667 INVX1_LOC_117/Y NAND2X1_LOC_122/Y 0.03fF
C5668 INVX1_LOC_586/A INVX1_LOC_186/Y 0.05fF
C5669 INVX1_LOC_117/Y INVX1_LOC_273/A 0.00fF
C5670 INVX1_LOC_153/A INVX1_LOC_94/A 0.02fF
C5671 NAND2X1_LOC_493/B INVX1_LOC_48/Y 0.02fF
C5672 INVX1_LOC_42/A INVX1_LOC_7/Y 0.01fF
C5673 INVX1_LOC_570/A INVX1_LOC_477/Y 0.03fF
C5674 INVX1_LOC_47/Y INVX1_LOC_253/A 0.02fF
C5675 VDD INVX1_LOC_612/A 0.01fF
C5676 INVX1_LOC_387/Y INVX1_LOC_45/Y 0.04fF
C5677 INVX1_LOC_134/Y NAND2X1_LOC_275/Y 0.02fF
C5678 INVX1_LOC_442/A INVX1_LOC_199/Y 0.03fF
C5679 INVX1_LOC_200/Y INVX1_LOC_9/Y 0.01fF
C5680 INVX1_LOC_96/A INVX1_LOC_94/A 0.31fF
C5681 INVX1_LOC_49/Y NAND2X1_LOC_506/B 0.22fF
C5682 INVX1_LOC_261/Y INVX1_LOC_340/Y 0.03fF
C5683 INVX1_LOC_425/A INVX1_LOC_89/Y 0.03fF
C5684 NAND2X1_LOC_710/A INVX1_LOC_361/Y 0.02fF
C5685 NAND2X1_LOC_616/Y INVX1_LOC_178/A 0.03fF
C5686 NAND2X1_LOC_79/a_36_24# NAND2X1_LOC_243/A 0.00fF
C5687 INVX1_LOC_206/Y INVX1_LOC_353/A 0.02fF
C5688 NAND2X1_LOC_13/Y NAND2X1_LOC_133/a_36_24# 0.00fF
C5689 INVX1_LOC_20/Y INVX1_LOC_31/Y 0.39fF
C5690 INVX1_LOC_121/Y INVX1_LOC_119/Y 0.59fF
C5691 INVX1_LOC_266/Y INVX1_LOC_69/Y 0.12fF
C5692 INVX1_LOC_45/Y INVX1_LOC_49/Y 0.49fF
C5693 NAND2X1_LOC_781/A INVX1_LOC_186/Y 0.03fF
C5694 INVX1_LOC_322/Y INVX1_LOC_63/Y 0.30fF
C5695 INVX1_LOC_651/Y INVX1_LOC_69/Y 0.13fF
C5696 INVX1_LOC_268/Y NAND2X1_LOC_837/A 0.01fF
C5697 NAND2X1_LOC_110/a_36_24# INVX1_LOC_26/Y 0.00fF
C5698 NAND2X1_LOC_275/Y INVX1_LOC_235/A 0.00fF
C5699 NAND2X1_LOC_145/a_36_24# INPUT_1 0.01fF
C5700 INVX1_LOC_361/Y INVX1_LOC_383/Y 0.00fF
C5701 INVX1_LOC_93/Y INVX1_LOC_375/Y 0.03fF
C5702 INVX1_LOC_119/Y INVX1_LOC_253/A 0.03fF
C5703 INVX1_LOC_11/Y INVX1_LOC_176/A 0.17fF
C5704 INVX1_LOC_586/A INVX1_LOC_328/Y 0.03fF
C5705 NAND2X1_LOC_574/a_36_24# NAND2X1_LOC_274/B 0.00fF
C5706 INVX1_LOC_649/Y NAND2X1_LOC_814/Y 0.21fF
C5707 INVX1_LOC_53/Y INVX1_LOC_66/A 0.07fF
C5708 INPUT_3 INVX1_LOC_49/Y 0.02fF
C5709 INVX1_LOC_51/Y INVX1_LOC_242/Y 1.01fF
C5710 NAND2X1_LOC_93/a_36_24# NAND2X1_LOC_333/B -0.02fF
C5711 INVX1_LOC_435/Y INVX1_LOC_41/Y 0.01fF
C5712 NAND2X1_LOC_267/A INVX1_LOC_98/Y 0.10fF
C5713 INVX1_LOC_286/Y INVX1_LOC_245/A 0.03fF
C5714 INVX1_LOC_300/A INVX1_LOC_31/Y 0.35fF
C5715 INVX1_LOC_155/A INVX1_LOC_154/Y 0.05fF
C5716 INVX1_LOC_84/A INVX1_LOC_223/Y 0.07fF
C5717 INVX1_LOC_20/Y INVX1_LOC_128/A 0.01fF
C5718 INVX1_LOC_596/A INVX1_LOC_301/Y 0.07fF
C5719 INVX1_LOC_266/A INVX1_LOC_242/Y 0.13fF
C5720 NAND2X1_LOC_285/A NAND2X1_LOC_285/B 0.04fF
C5721 INVX1_LOC_197/A INVX1_LOC_168/Y 0.07fF
C5722 NAND2X1_LOC_76/a_36_24# INVX1_LOC_74/Y 0.00fF
C5723 INVX1_LOC_63/Y NAND2X1_LOC_496/Y 0.20fF
C5724 INVX1_LOC_358/Y INVX1_LOC_338/Y 0.56fF
C5725 INVX1_LOC_513/A INVX1_LOC_50/Y 0.21fF
C5726 INVX1_LOC_335/Y INVX1_LOC_497/A 0.06fF
C5727 NAND2X1_LOC_616/Y INVX1_LOC_58/Y 0.04fF
C5728 INVX1_LOC_89/Y INVX1_LOC_252/Y 0.03fF
C5729 INVX1_LOC_335/Y INVX1_LOC_338/Y 0.00fF
C5730 NAND2X1_LOC_673/B INVX1_LOC_46/Y 0.02fF
C5731 INVX1_LOC_21/Y INVX1_LOC_338/Y 0.22fF
C5732 NAND2X1_LOC_702/a_36_24# INVX1_LOC_6/Y 0.00fF
C5733 INVX1_LOC_413/Y NAND2X1_LOC_844/A 0.01fF
C5734 INVX1_LOC_199/Y INVX1_LOC_116/Y 0.07fF
C5735 INVX1_LOC_347/Y NAND2X1_LOC_808/a_36_24# 0.00fF
C5736 INVX1_LOC_154/A INVX1_LOC_252/Y 0.02fF
C5737 INVX1_LOC_213/Y INVX1_LOC_391/A 0.02fF
C5738 INPUT_1 INVX1_LOC_670/A 0.04fF
C5739 NAND2X1_LOC_775/B INVX1_LOC_253/Y 0.03fF
C5740 INVX1_LOC_63/Y NAND2X1_LOC_266/a_36_24# 0.00fF
C5741 INVX1_LOC_103/Y INVX1_LOC_32/Y 0.03fF
C5742 NAND2X1_LOC_395/a_36_24# NAND2X1_LOC_294/Y 0.01fF
C5743 NAND2X1_LOC_517/Y INVX1_LOC_405/Y 0.09fF
C5744 INVX1_LOC_339/Y INVX1_LOC_7/Y 0.09fF
C5745 INVX1_LOC_32/Y INVX1_LOC_68/A 0.03fF
C5746 INVX1_LOC_183/A INVX1_LOC_42/Y 0.00fF
C5747 INVX1_LOC_11/Y INVX1_LOC_170/Y 0.02fF
C5748 INVX1_LOC_54/Y INVX1_LOC_419/A 0.01fF
C5749 INVX1_LOC_596/A INVX1_LOC_41/Y 0.03fF
C5750 INVX1_LOC_54/Y INVX1_LOC_234/Y 0.07fF
C5751 INVX1_LOC_93/Y NAND2X1_LOC_622/a_36_24# 0.00fF
C5752 INVX1_LOC_53/Y NAND2X1_LOC_601/Y 0.04fF
C5753 INVX1_LOC_345/Y INVX1_LOC_346/A 0.00fF
C5754 NAND2X1_LOC_786/B INVX1_LOC_228/A 0.05fF
C5755 INVX1_LOC_17/Y INVX1_LOC_245/A 0.12fF
C5756 INVX1_LOC_346/A INVX1_LOC_32/Y 0.08fF
C5757 INVX1_LOC_6/Y NAND2X1_LOC_225/a_36_24# -0.00fF
C5758 NAND2X1_LOC_318/B INVX1_LOC_41/Y 0.02fF
C5759 INVX1_LOC_504/Y INVX1_LOC_114/A 0.10fF
C5760 INVX1_LOC_633/Y INVX1_LOC_588/A 0.03fF
C5761 INVX1_LOC_588/Y NAND2X1_LOC_686/A 0.14fF
C5762 INVX1_LOC_282/A INVX1_LOC_663/A 0.01fF
C5763 INVX1_LOC_366/Y INVX1_LOC_41/Y 0.00fF
C5764 INVX1_LOC_625/A INVX1_LOC_531/Y 0.03fF
C5765 INVX1_LOC_402/A INVX1_LOC_479/A 0.01fF
C5766 INVX1_LOC_47/Y NAND2X1_LOC_498/a_36_24# 0.01fF
C5767 INVX1_LOC_49/Y NAND2X1_LOC_837/A 0.19fF
C5768 INVX1_LOC_255/A INVX1_LOC_199/Y 0.03fF
C5769 INVX1_LOC_177/A INVX1_LOC_41/Y 0.01fF
C5770 NAND2X1_LOC_148/A INVX1_LOC_212/A 0.00fF
C5771 INVX1_LOC_507/A INVX1_LOC_58/Y 0.01fF
C5772 NAND2X1_LOC_136/Y INVX1_LOC_520/A 0.10fF
C5773 INVX1_LOC_166/A INVX1_LOC_519/Y 0.02fF
C5774 INVX1_LOC_54/Y INVX1_LOC_665/A 0.03fF
C5775 INVX1_LOC_62/Y NAND2X1_LOC_826/a_36_24# 0.01fF
C5776 INVX1_LOC_507/Y INVX1_LOC_496/A 0.01fF
C5777 INVX1_LOC_179/A INVX1_LOC_199/Y 0.71fF
C5778 NAND2X1_LOC_615/Y INVX1_LOC_482/Y 0.00fF
C5779 INVX1_LOC_77/A INVX1_LOC_77/Y 0.01fF
C5780 INVX1_LOC_426/A INVX1_LOC_301/A 0.01fF
C5781 INVX1_LOC_463/Y INVX1_LOC_74/Y 0.15fF
C5782 INVX1_LOC_372/A INVX1_LOC_74/Y 0.11fF
C5783 INVX1_LOC_376/A NAND2X1_LOC_470/a_36_24# 0.02fF
C5784 NAND2X1_LOC_294/Y INVX1_LOC_450/Y 0.02fF
C5785 INVX1_LOC_531/Y NAND2X1_LOC_52/Y 0.01fF
C5786 INVX1_LOC_73/Y INVX1_LOC_395/A 0.02fF
C5787 NAND2X1_LOC_846/B INVX1_LOC_667/A 0.02fF
C5788 INVX1_LOC_26/Y INVX1_LOC_90/Y 0.06fF
C5789 NAND2X1_LOC_274/B INVX1_LOC_100/Y 0.07fF
C5790 NAND2X1_LOC_373/Y INVX1_LOC_395/A 0.62fF
C5791 INVX1_LOC_301/A NAND2X1_LOC_539/a_36_24# 0.01fF
C5792 NAND2X1_LOC_274/B INVX1_LOC_74/Y 0.04fF
C5793 NAND2X1_LOC_249/Y NAND2X1_LOC_249/a_36_24# 0.02fF
C5794 INPUT_3 INVX1_LOC_297/Y 0.09fF
C5795 INVX1_LOC_395/A INVX1_LOC_553/A 0.03fF
C5796 NAND2X1_LOC_537/B NAND2X1_LOC_536/a_36_24# 0.01fF
C5797 INVX1_LOC_20/Y NAND2X1_LOC_592/a_36_24# 0.01fF
C5798 INVX1_LOC_20/Y INVX1_LOC_426/A 0.46fF
C5799 INVX1_LOC_554/A INVX1_LOC_146/A 0.26fF
C5800 VDD INVX1_LOC_616/A -0.00fF
C5801 INVX1_LOC_266/A INVX1_LOC_301/A 1.56fF
C5802 INVX1_LOC_68/Y INVX1_LOC_206/Y 0.91fF
C5803 INVX1_LOC_409/Y INVX1_LOC_686/A 0.07fF
C5804 NAND2X1_LOC_322/Y INVX1_LOC_686/A 0.03fF
C5805 INVX1_LOC_479/A INVX1_LOC_653/Y 0.00fF
C5806 NAND2X1_LOC_69/B INVX1_LOC_307/A 0.36fF
C5807 VDD INVX1_LOC_424/Y 0.43fF
C5808 INVX1_LOC_446/A NAND2X1_LOC_658/a_36_24# 0.00fF
C5809 VDD INVX1_LOC_229/Y 0.24fF
C5810 INVX1_LOC_317/Y INVX1_LOC_65/Y 0.03fF
C5811 VDD NAND2X1_LOC_324/B 0.01fF
C5812 INVX1_LOC_533/Y INVX1_LOC_51/Y 0.26fF
C5813 INPUT_0 INVX1_LOC_551/Y 0.08fF
C5814 NAND2X1_LOC_498/B INVX1_LOC_45/Y 0.01fF
C5815 INVX1_LOC_98/A INVX1_LOC_45/Y 0.01fF
C5816 INVX1_LOC_428/A NAND2X1_LOC_486/B 0.01fF
C5817 INVX1_LOC_412/Y NAND2X1_LOC_804/a_36_24# 0.00fF
C5818 VDD INVX1_LOC_130/Y 0.00fF
C5819 NAND2X1_LOC_516/Y INVX1_LOC_551/Y 0.03fF
C5820 INVX1_LOC_76/Y INVX1_LOC_45/Y 0.10fF
C5821 NAND2X1_LOC_475/A INVX1_LOC_296/Y 0.01fF
C5822 INVX1_LOC_69/Y INVX1_LOC_109/Y 0.03fF
C5823 INVX1_LOC_206/Y NAND2X1_LOC_130/Y 0.04fF
C5824 INVX1_LOC_103/A INVX1_LOC_134/Y 0.01fF
C5825 INVX1_LOC_206/Y INVX1_LOC_600/A 0.19fF
C5826 INVX1_LOC_279/Y INVX1_LOC_282/A 0.03fF
C5827 INVX1_LOC_20/Y INVX1_LOC_51/Y 7.76fF
C5828 VDD NAND2X1_LOC_226/Y 0.04fF
C5829 NAND2X1_LOC_776/a_36_24# INVX1_LOC_80/A 0.01fF
C5830 NAND2X1_LOC_790/B NAND2X1_LOC_165/Y 0.02fF
C5831 INVX1_LOC_442/A INVX1_LOC_53/Y 0.02fF
C5832 INVX1_LOC_238/Y INVX1_LOC_556/Y 0.01fF
C5833 NAND2X1_LOC_768/a_36_24# NAND2X1_LOC_332/B 0.00fF
C5834 INPUT_3 INVX1_LOC_76/Y 0.04fF
C5835 INVX1_LOC_20/Y INVX1_LOC_266/A 0.06fF
C5836 NAND2X1_LOC_453/a_36_24# INVX1_LOC_638/A 0.01fF
C5837 INVX1_LOC_278/A INVX1_LOC_453/Y 0.03fF
C5838 VDD INVX1_LOC_110/A -0.00fF
C5839 NAND2X1_LOC_558/a_36_24# INVX1_LOC_230/A 0.00fF
C5840 NAND2X1_LOC_586/Y INVX1_LOC_638/A 0.05fF
C5841 INVX1_LOC_51/Y NAND2X1_LOC_605/a_36_24# 0.01fF
C5842 INVX1_LOC_325/Y INVX1_LOC_46/A 0.09fF
C5843 NAND2X1_LOC_20/Y INVX1_LOC_84/A 0.01fF
C5844 INVX1_LOC_602/A INVX1_LOC_45/A 0.02fF
C5845 INPUT_0 INVX1_LOC_493/A 0.03fF
C5846 NAND2X1_LOC_324/a_36_24# INVX1_LOC_374/A 0.00fF
C5847 INVX1_LOC_559/A INVX1_LOC_45/Y 0.01fF
C5848 INVX1_LOC_300/A INVX1_LOC_51/Y 0.07fF
C5849 INPUT_0 INVX1_LOC_167/A 0.12fF
C5850 NAND2X1_LOC_399/a_36_24# INVX1_LOC_322/Y 0.00fF
C5851 INVX1_LOC_51/Y INVX1_LOC_197/Y 0.03fF
C5852 NAND2X1_LOC_513/a_36_24# INVX1_LOC_401/A 0.00fF
C5853 NAND2X1_LOC_759/B INVX1_LOC_63/Y 0.02fF
C5854 NAND2X1_LOC_231/A INVX1_LOC_59/Y 0.00fF
C5855 INVX1_LOC_530/Y NAND2X1_LOC_673/B 0.10fF
C5856 INVX1_LOC_335/A INVX1_LOC_586/A 0.03fF
C5857 INPUT_0 NAND2X1_LOC_141/a_36_24# 0.01fF
C5858 INVX1_LOC_266/A INVX1_LOC_300/A 0.36fF
C5859 INVX1_LOC_401/A INVX1_LOC_516/A 0.02fF
C5860 INVX1_LOC_366/A INVX1_LOC_195/Y 0.03fF
C5861 INVX1_LOC_20/Y NAND2X1_LOC_267/a_36_24# 0.00fF
C5862 NAND2X1_LOC_155/a_36_24# INVX1_LOC_137/Y 0.00fF
C5863 INPUT_0 INVX1_LOC_486/A 0.08fF
C5864 INVX1_LOC_108/A INVX1_LOC_45/Y 0.01fF
C5865 INVX1_LOC_288/A INVX1_LOC_359/A 0.07fF
C5866 INVX1_LOC_447/Y INVX1_LOC_80/A 0.00fF
C5867 INVX1_LOC_97/A INVX1_LOC_63/Y 0.03fF
C5868 INVX1_LOC_616/A NAND2X1_LOC_243/A 0.02fF
C5869 INVX1_LOC_53/Y INVX1_LOC_116/Y 0.12fF
C5870 INVX1_LOC_21/Y NAND2X1_LOC_318/B 0.01fF
C5871 INVX1_LOC_288/A NAND2X1_LOC_466/a_36_24# 0.00fF
C5872 INVX1_LOC_21/Y INVX1_LOC_366/Y 0.00fF
C5873 INVX1_LOC_84/A INVX1_LOC_295/Y 0.34fF
C5874 NAND2X1_LOC_370/A INVX1_LOC_58/Y 0.00fF
C5875 INVX1_LOC_340/Y INVX1_LOC_637/Y 0.01fF
C5876 INVX1_LOC_257/Y NAND2X1_LOC_301/B 0.07fF
C5877 INVX1_LOC_54/Y INVX1_LOC_80/A 0.19fF
C5878 INVX1_LOC_21/Y INVX1_LOC_177/A 0.00fF
C5879 INVX1_LOC_41/Y NAND2X1_LOC_76/B 0.21fF
C5880 INVX1_LOC_312/Y INVX1_LOC_105/Y 0.03fF
C5881 INVX1_LOC_273/A INVX1_LOC_58/Y 0.00fF
C5882 NAND2X1_LOC_672/a_36_24# NAND2X1_LOC_616/Y 0.00fF
C5883 INVX1_LOC_117/Y INVX1_LOC_519/A 0.03fF
C5884 INVX1_LOC_579/A INVX1_LOC_117/Y 0.03fF
C5885 INVX1_LOC_397/A NAND2X1_LOC_445/a_36_24# 0.00fF
C5886 INVX1_LOC_293/Y INVX1_LOC_387/Y 0.03fF
C5887 NAND2X1_LOC_635/B INVX1_LOC_676/Y 0.91fF
C5888 INVX1_LOC_163/Y INVX1_LOC_496/A 0.03fF
C5889 NAND2X1_LOC_106/Y INVX1_LOC_367/A 0.02fF
C5890 INVX1_LOC_85/Y INVX1_LOC_179/Y 0.00fF
C5891 NAND2X1_LOC_164/Y INVX1_LOC_531/Y 0.09fF
C5892 INVX1_LOC_171/A INVX1_LOC_7/Y 0.06fF
C5893 NAND2X1_LOC_169/A INVX1_LOC_48/Y 0.04fF
C5894 INVX1_LOC_174/A INVX1_LOC_87/A 0.00fF
C5895 NAND2X1_LOC_779/a_36_24# INVX1_LOC_137/Y -0.00fF
C5896 NAND2X1_LOC_498/Y INVX1_LOC_652/A 0.02fF
C5897 NAND2X1_LOC_501/a_36_24# NAND2X1_LOC_274/B 0.00fF
C5898 INVX1_LOC_599/A INVX1_LOC_601/Y 0.01fF
C5899 INVX1_LOC_435/A INVX1_LOC_681/Y 0.01fF
C5900 INVX1_LOC_293/Y INVX1_LOC_49/Y 0.07fF
C5901 INVX1_LOC_237/Y INVX1_LOC_100/Y 0.01fF
C5902 INVX1_LOC_285/A INVX1_LOC_69/Y 0.00fF
C5903 INVX1_LOC_490/Y NAND2X1_LOC_528/Y 0.02fF
C5904 INVX1_LOC_330/A INVX1_LOC_335/A 0.07fF
C5905 NAND2X1_LOC_540/a_36_24# INVX1_LOC_17/Y 0.01fF
C5906 INVX1_LOC_449/A INVX1_LOC_6/Y 0.32fF
C5907 INVX1_LOC_257/A INVX1_LOC_80/A 0.01fF
C5908 INVX1_LOC_602/A INVX1_LOC_659/A 0.02fF
C5909 INVX1_LOC_435/A INPUT_1 0.07fF
C5910 INVX1_LOC_11/Y NAND2X1_LOC_187/Y 0.16fF
C5911 INPUT_0 NAND2X1_LOC_410/Y 0.02fF
C5912 NAND2X1_LOC_619/Y INVX1_LOC_99/Y 0.01fF
C5913 INVX1_LOC_616/A NAND2X1_LOC_786/B 0.00fF
C5914 INVX1_LOC_11/Y INVX1_LOC_54/Y 4.95fF
C5915 INVX1_LOC_110/A INVX1_LOC_509/A 0.17fF
C5916 INVX1_LOC_65/Y INVX1_LOC_531/Y 0.14fF
C5917 NAND2X1_LOC_13/Y INVX1_LOC_242/Y 0.02fF
C5918 INVX1_LOC_63/Y INVX1_LOC_633/Y 0.02fF
C5919 INVX1_LOC_107/A NAND2X1_LOC_248/B 0.02fF
C5920 INVX1_LOC_366/A INVX1_LOC_207/Y 0.03fF
C5921 INVX1_LOC_328/Y INVX1_LOC_486/Y 0.05fF
C5922 INVX1_LOC_294/Y INVX1_LOC_328/Y 0.03fF
C5923 NAND2X1_LOC_320/Y INVX1_LOC_69/Y 0.03fF
C5924 NAND2X1_LOC_646/a_36_24# INVX1_LOC_496/A 0.00fF
C5925 INVX1_LOC_47/Y INVX1_LOC_251/A 0.04fF
C5926 INVX1_LOC_670/A INVX1_LOC_50/Y 0.01fF
C5927 INVX1_LOC_59/Y INVX1_LOC_77/Y 0.01fF
C5928 INVX1_LOC_128/A INVX1_LOC_375/Y 0.06fF
C5929 NAND2X1_LOC_180/B INVX1_LOC_62/Y 0.03fF
C5930 INVX1_LOC_342/Y INVX1_LOC_69/Y 0.06fF
C5931 INVX1_LOC_366/A INVX1_LOC_597/Y 0.00fF
C5932 INVX1_LOC_369/A INVX1_LOC_90/Y 0.09fF
C5933 NAND2X1_LOC_673/B INVX1_LOC_49/Y 0.07fF
C5934 NAND2X1_LOC_106/Y INVX1_LOC_93/Y 0.03fF
C5935 INVX1_LOC_469/Y INVX1_LOC_372/A 0.01fF
C5936 INVX1_LOC_541/Y INVX1_LOC_41/Y 0.01fF
C5937 INVX1_LOC_346/A NAND2X1_LOC_652/a_36_24# 0.00fF
C5938 INVX1_LOC_35/A INVX1_LOC_1/Y 0.02fF
C5939 INVX1_LOC_551/Y INVX1_LOC_211/A 0.02fF
C5940 INVX1_LOC_188/Y INVX1_LOC_62/Y 0.03fF
C5941 INVX1_LOC_251/A INVX1_LOC_119/Y 0.06fF
C5942 INVX1_LOC_63/Y INVX1_LOC_317/A 0.00fF
C5943 INVX1_LOC_344/A NAND2X1_LOC_434/a_36_24# 0.00fF
C5944 INVX1_LOC_625/A INVX1_LOC_41/Y 0.02fF
C5945 INVX1_LOC_544/Y INVX1_LOC_66/A 0.01fF
C5946 INVX1_LOC_47/Y NAND2X1_LOC_424/a_36_24# 0.01fF
C5947 INVX1_LOC_418/Y INVX1_LOC_100/Y 0.00fF
C5948 NAND2X1_LOC_545/a_36_24# INVX1_LOC_255/A 0.00fF
C5949 INVX1_LOC_69/Y INVX1_LOC_199/Y 0.13fF
C5950 INVX1_LOC_12/Y INVX1_LOC_666/Y 0.06fF
C5951 INVX1_LOC_100/Y INVX1_LOC_159/Y 0.15fF
C5952 INVX1_LOC_300/Y INVX1_LOC_340/A 0.03fF
C5953 INVX1_LOC_17/Y NAND2X1_LOC_597/Y 0.16fF
C5954 INVX1_LOC_347/A INVX1_LOC_252/Y 0.07fF
C5955 INVX1_LOC_117/A INVX1_LOC_46/Y 0.00fF
C5956 INVX1_LOC_328/Y INVX1_LOC_6/Y 0.03fF
C5957 NAND2X1_LOC_274/B INVX1_LOC_350/Y 0.01fF
C5958 INVX1_LOC_248/A NAND2X1_LOC_301/B 0.00fF
C5959 INVX1_LOC_662/A INVX1_LOC_66/A 0.01fF
C5960 INVX1_LOC_261/A INPUT_4 0.03fF
C5961 INVX1_LOC_6/Y INVX1_LOC_518/A 0.03fF
C5962 NAND2X1_LOC_619/Y NAND2X1_LOC_66/Y 0.01fF
C5963 INVX1_LOC_159/Y INVX1_LOC_74/Y 0.09fF
C5964 NAND2X1_LOC_547/a_36_24# INVX1_LOC_502/A 0.01fF
C5965 INVX1_LOC_93/Y NAND2X1_LOC_123/B 0.03fF
C5966 NAND2X1_LOC_181/A NAND2X1_LOC_274/B 0.17fF
C5967 INVX1_LOC_318/A INVX1_LOC_531/Y 0.01fF
C5968 INVX1_LOC_69/Y INVX1_LOC_272/A 0.01fF
C5969 INVX1_LOC_47/Y INVX1_LOC_652/A 0.02fF
C5970 INVX1_LOC_6/Y INVX1_LOC_207/Y 0.09fF
C5971 INVX1_LOC_242/Y INVX1_LOC_361/A 0.02fF
C5972 INVX1_LOC_100/Y INVX1_LOC_212/Y 0.03fF
C5973 INVX1_LOC_26/Y INVX1_LOC_338/Y 0.09fF
C5974 INVX1_LOC_397/Y INVX1_LOC_531/Y 0.13fF
C5975 INVX1_LOC_166/A INVX1_LOC_588/A -0.00fF
C5976 INVX1_LOC_660/A INVX1_LOC_340/A 0.03fF
C5977 NAND2X1_LOC_285/A NAND2X1_LOC_248/B 0.20fF
C5978 INVX1_LOC_225/Y INVX1_LOC_224/A 0.00fF
C5979 INVX1_LOC_586/A INVX1_LOC_109/Y 0.06fF
C5980 NAND2X1_LOC_283/a_36_24# INVX1_LOC_669/A 0.01fF
C5981 INVX1_LOC_675/A NAND2X1_LOC_123/B 0.03fF
C5982 INVX1_LOC_6/Y INVX1_LOC_597/Y 0.01fF
C5983 INVX1_LOC_95/A INVX1_LOC_531/Y 0.02fF
C5984 INVX1_LOC_662/A NAND2X1_LOC_848/a_36_24# 0.01fF
C5985 INPUT_0 INVX1_LOC_596/Y 0.00fF
C5986 INVX1_LOC_185/A INVX1_LOC_523/A 0.03fF
C5987 NAND2X1_LOC_274/B INVX1_LOC_79/A 0.07fF
C5988 INVX1_LOC_95/Y INVX1_LOC_586/A 0.00fF
C5989 INVX1_LOC_652/A INVX1_LOC_119/Y 0.02fF
C5990 INVX1_LOC_62/Y INVX1_LOC_491/A 0.32fF
C5991 INVX1_LOC_312/Y INVX1_LOC_109/Y 0.25fF
C5992 INVX1_LOC_93/Y INVX1_LOC_92/A 0.96fF
C5993 INVX1_LOC_47/Y INVX1_LOC_462/Y 0.06fF
C5994 INVX1_LOC_554/A INVX1_LOC_586/A 0.01fF
C5995 INVX1_LOC_100/Y INVX1_LOC_468/A 0.05fF
C5996 INVX1_LOC_20/Y INVX1_LOC_463/A 0.27fF
C5997 INVX1_LOC_20/Y NAND2X1_LOC_537/A 0.08fF
C5998 NAND2X1_LOC_763/Y INVX1_LOC_366/A 0.01fF
C5999 INVX1_LOC_266/A NAND2X1_LOC_373/Y 0.18fF
C6000 INPUT_0 INVX1_LOC_558/A 0.03fF
C6001 NAND2X1_LOC_552/a_36_24# INVX1_LOC_578/A 0.00fF
C6002 INVX1_LOC_375/A INVX1_LOC_624/A 0.02fF
C6003 INVX1_LOC_374/A NAND2X1_LOC_831/a_36_24# 0.00fF
C6004 NAND2X1_LOC_516/Y INVX1_LOC_558/A 0.04fF
C6005 VDD NAND2X1_LOC_299/Y 0.03fF
C6006 NAND2X1_LOC_534/Y INVX1_LOC_80/A 0.01fF
C6007 INVX1_LOC_68/Y INVX1_LOC_397/A 0.00fF
C6008 INVX1_LOC_68/Y INVX1_LOC_94/A 0.34fF
C6009 INVX1_LOC_21/Y NAND2X1_LOC_76/B 0.07fF
C6010 INVX1_LOC_20/Y NAND2X1_LOC_114/a_36_24# 0.00fF
C6011 INVX1_LOC_206/Y NAND2X1_LOC_56/Y 0.03fF
C6012 NAND2X1_LOC_336/B NAND2X1_LOC_312/a_36_24# 0.00fF
C6013 INVX1_LOC_20/Y NAND2X1_LOC_108/Y 0.72fF
C6014 INVX1_LOC_340/Y NAND2X1_LOC_707/A 0.01fF
C6015 GATE_579 NAND2X1_LOC_580/a_36_24# 0.01fF
C6016 NAND2X1_LOC_763/Y INVX1_LOC_597/A 0.00fF
C6017 INVX1_LOC_84/A INVX1_LOC_173/A 0.01fF
C6018 NAND2X1_LOC_756/Y INVX1_LOC_98/A 0.07fF
C6019 NAND2X1_LOC_45/Y INVX1_LOC_379/A 0.10fF
C6020 NAND2X1_LOC_45/Y INVX1_LOC_35/Y 0.03fF
C6021 INVX1_LOC_374/A INVX1_LOC_633/Y 0.33fF
C6022 INVX1_LOC_395/A INVX1_LOC_567/Y 0.04fF
C6023 NAND2X1_LOC_505/a_36_24# INVX1_LOC_600/A 0.01fF
C6024 INVX1_LOC_20/Y NAND2X1_LOC_13/Y 1.04fF
C6025 INVX1_LOC_410/Y INVX1_LOC_230/A 0.07fF
C6026 INVX1_LOC_397/A INVX1_LOC_600/A 0.34fF
C6027 INPUT_0 INVX1_LOC_211/Y 0.01fF
C6028 NAND2X1_LOC_267/A NAND2X1_LOC_76/B 0.05fF
C6029 INVX1_LOC_438/Y INVX1_LOC_439/Y 0.39fF
C6030 VDD NAND2X1_LOC_184/Y 0.39fF
C6031 INVX1_LOC_560/A INVX1_LOC_98/Y 1.13fF
C6032 NAND2X1_LOC_820/Y INVX1_LOC_668/A 0.06fF
C6033 INVX1_LOC_616/A INVX1_LOC_619/A 0.01fF
C6034 NAND2X1_LOC_506/a_36_24# INVX1_LOC_96/Y 0.00fF
C6035 INVX1_LOC_492/A INVX1_LOC_606/Y 0.01fF
C6036 NAND2X1_LOC_710/A NAND2X1_LOC_700/a_36_24# 0.02fF
C6037 INVX1_LOC_85/Y INVX1_LOC_205/Y 0.00fF
C6038 INVX1_LOC_45/Y INVX1_LOC_7/Y 0.17fF
C6039 NAND2X1_LOC_498/Y INVX1_LOC_35/Y 0.07fF
C6040 INVX1_LOC_570/A INVX1_LOC_35/Y 0.13fF
C6041 NAND2X1_LOC_740/a_36_24# INVX1_LOC_583/A 0.02fF
C6042 INPUT_0 NAND2X1_LOC_749/a_36_24# 0.00fF
C6043 INVX1_LOC_508/Y INVX1_LOC_517/A 0.00fF
C6044 INVX1_LOC_45/Y NAND2X1_LOC_259/A 0.01fF
C6045 INPUT_0 INVX1_LOC_46/Y 0.10fF
C6046 INVX1_LOC_142/Y INVX1_LOC_186/A 0.01fF
C6047 NAND2X1_LOC_763/Y INVX1_LOC_6/Y 0.01fF
C6048 INPUT_2 INVX1_LOC_27/Y 0.01fF
C6049 INVX1_LOC_182/A INVX1_LOC_198/A 0.04fF
C6050 INPUT_0 NAND2X1_LOC_187/a_36_24# 0.00fF
C6051 INVX1_LOC_85/Y INVX1_LOC_194/Y 0.00fF
C6052 NAND2X1_LOC_13/Y INVX1_LOC_300/A 0.08fF
C6053 INVX1_LOC_224/Y INVX1_LOC_187/Y 0.09fF
C6054 INVX1_LOC_150/A INVX1_LOC_58/Y 0.00fF
C6055 VDD INVX1_LOC_498/Y 0.21fF
C6056 INVX1_LOC_541/Y INVX1_LOC_358/Y 0.01fF
C6057 INVX1_LOC_679/Y INVX1_LOC_367/A 0.01fF
C6058 INVX1_LOC_409/Y INVX1_LOC_376/Y 0.01fF
C6059 INPUT_3 INVX1_LOC_7/Y 0.91fF
C6060 INVX1_LOC_602/Y INVX1_LOC_59/A 0.01fF
C6061 INVX1_LOC_406/Y INVX1_LOC_451/Y 0.11fF
C6062 NAND2X1_LOC_379/Y INVX1_LOC_310/Y 0.04fF
C6063 INVX1_LOC_335/Y INVX1_LOC_541/Y 0.01fF
C6064 INPUT_6 INPUT_5 0.03fF
C6065 INVX1_LOC_392/Y INPUT_1 0.05fF
C6066 NAND2X1_LOC_537/B INVX1_LOC_199/Y 0.11fF
C6067 INVX1_LOC_32/Y NAND2X1_LOC_506/B 0.23fF
C6068 NAND2X1_LOC_790/B INVX1_LOC_90/Y 1.00fF
C6069 INVX1_LOC_45/Y INVX1_LOC_32/Y 0.85fF
C6070 INPUT_6 INVX1_LOC_2/Y 0.01fF
C6071 INVX1_LOC_133/Y INVX1_LOC_669/A 0.01fF
C6072 NAND2X1_LOC_585/a_36_24# INVX1_LOC_245/A 0.01fF
C6073 NAND2X1_LOC_603/Y INVX1_LOC_469/A 0.09fF
C6074 INVX1_LOC_21/Y INVX1_LOC_530/A 0.01fF
C6075 INVX1_LOC_523/A INVX1_LOC_58/Y 0.01fF
C6076 INVX1_LOC_587/A NAND2X1_LOC_821/a_36_24# 0.00fF
C6077 INVX1_LOC_345/Y INVX1_LOC_348/A 0.01fF
C6078 NAND2X1_LOC_16/Y INVX1_LOC_170/A 0.01fF
C6079 INVX1_LOC_442/Y INVX1_LOC_385/Y 0.12fF
C6080 INVX1_LOC_625/A INVX1_LOC_21/Y 0.04fF
C6081 INVX1_LOC_7/Y NAND2X1_LOC_376/Y 0.03fF
C6082 INVX1_LOC_586/A INVX1_LOC_199/Y 0.10fF
C6083 INVX1_LOC_367/A INPUT_1 0.08fF
C6084 INPUT_3 INVX1_LOC_32/Y 0.15fF
C6085 INVX1_LOC_317/Y INVX1_LOC_63/Y 0.23fF
C6086 INVX1_LOC_415/Y INVX1_LOC_449/A 0.01fF
C6087 INVX1_LOC_206/Y INVX1_LOC_369/Y 0.07fF
C6088 INVX1_LOC_537/A INVX1_LOC_357/A 0.01fF
C6089 INVX1_LOC_431/A INVX1_LOC_12/Y 0.00fF
C6090 INVX1_LOC_85/Y INVX1_LOC_44/Y 0.01fF
C6091 INVX1_LOC_35/Y INVX1_LOC_99/Y 0.20fF
C6092 NAND2X1_LOC_370/A INVX1_LOC_245/A 0.01fF
C6093 INVX1_LOC_53/Y NAND2X1_LOC_148/B 0.01fF
C6094 VDD INVX1_LOC_75/Y 1.96fF
C6095 INVX1_LOC_20/Y INVX1_LOC_380/Y 0.33fF
C6096 INVX1_LOC_269/A INVX1_LOC_9/Y 0.68fF
C6097 INVX1_LOC_435/Y INVX1_LOC_26/Y 1.78fF
C6098 NAND2X1_LOC_755/B INVX1_LOC_527/Y 0.00fF
C6099 NAND2X1_LOC_114/a_36_24# INVX1_LOC_655/A 0.00fF
C6100 NAND2X1_LOC_122/Y INVX1_LOC_245/A 0.03fF
C6101 INVX1_LOC_402/Y INVX1_LOC_50/Y 0.03fF
C6102 INVX1_LOC_93/Y INVX1_LOC_679/Y 0.03fF
C6103 INVX1_LOC_626/A INVX1_LOC_54/Y 0.02fF
C6104 NAND2X1_LOC_108/Y INVX1_LOC_655/A 0.06fF
C6105 INVX1_LOC_166/A INVX1_LOC_670/Y 0.00fF
C6106 NAND2X1_LOC_318/a_36_24# INVX1_LOC_600/A 0.01fF
C6107 INVX1_LOC_20/Y INVX1_LOC_361/A 0.06fF
C6108 INVX1_LOC_450/A INVX1_LOC_405/Y 0.02fF
C6109 INVX1_LOC_80/A INVX1_LOC_89/Y 0.15fF
C6110 INPUT_4 INVX1_LOC_69/A 0.06fF
C6111 INVX1_LOC_516/A INPUT_1 0.02fF
C6112 INVX1_LOC_549/Y INVX1_LOC_48/Y 0.08fF
C6113 INVX1_LOC_586/A INVX1_LOC_272/A 0.03fF
C6114 INVX1_LOC_298/A NAND2X1_LOC_755/B 1.89fF
C6115 INVX1_LOC_625/A NAND2X1_LOC_267/A 0.02fF
C6116 INVX1_LOC_669/Y INPUT_1 0.03fF
C6117 INVX1_LOC_54/Y INVX1_LOC_367/Y 0.00fF
C6118 INVX1_LOC_53/Y INVX1_LOC_69/Y 8.97fF
C6119 INVX1_LOC_43/Y INVX1_LOC_87/A 0.01fF
C6120 INVX1_LOC_203/Y NAND2X1_LOC_231/B 0.03fF
C6121 INVX1_LOC_435/A INVX1_LOC_50/Y 0.08fF
C6122 INVX1_LOC_99/Y NAND2X1_LOC_448/B 0.02fF
C6123 INVX1_LOC_672/A NAND2X1_LOC_851/a_36_24# 0.02fF
C6124 INVX1_LOC_607/Y INVX1_LOC_46/Y 0.05fF
C6125 INVX1_LOC_402/A INVX1_LOC_66/A 0.00fF
C6126 INVX1_LOC_206/Y INVX1_LOC_223/A 0.09fF
C6127 INVX1_LOC_192/Y INVX1_LOC_666/Y 0.01fF
C6128 INVX1_LOC_99/Y INVX1_LOC_620/A 0.03fF
C6129 INVX1_LOC_376/A INVX1_LOC_197/A 0.07fF
C6130 NAND2X1_LOC_130/Y NAND2X1_LOC_542/A 0.05fF
C6131 INVX1_LOC_325/Y INVX1_LOC_245/A 0.15fF
C6132 INVX1_LOC_65/Y INVX1_LOC_41/Y 0.33fF
C6133 NAND2X1_LOC_184/Y NAND2X1_LOC_843/A 0.05fF
C6134 NAND2X1_LOC_834/a_36_24# INVX1_LOC_476/Y -0.00fF
C6135 INVX1_LOC_80/A INVX1_LOC_501/A 0.03fF
C6136 INVX1_LOC_206/Y INVX1_LOC_348/Y 0.06fF
C6137 INVX1_LOC_257/Y INVX1_LOC_634/Y 0.19fF
C6138 INVX1_LOC_435/A INVX1_LOC_431/Y 0.00fF
C6139 VDD NAND2X1_LOC_271/A 0.30fF
C6140 INVX1_LOC_391/Y NAND2X1_LOC_521/Y 0.06fF
C6141 NAND2X1_LOC_24/Y INVX1_LOC_9/Y 0.03fF
C6142 INVX1_LOC_589/Y INVX1_LOC_35/Y 0.07fF
C6143 NAND2X1_LOC_538/B INVX1_LOC_79/A 0.02fF
C6144 INVX1_LOC_568/A INVX1_LOC_35/Y 0.01fF
C6145 NAND2X1_LOC_106/Y INVX1_LOC_548/A 0.22fF
C6146 INVX1_LOC_172/Y INVX1_LOC_100/Y 0.06fF
C6147 INVX1_LOC_17/Y INVX1_LOC_293/A 0.03fF
C6148 INVX1_LOC_11/Y INVX1_LOC_89/Y 0.22fF
C6149 INVX1_LOC_47/Y INVX1_LOC_35/Y 0.35fF
C6150 INVX1_LOC_372/A INVX1_LOC_48/Y 0.01fF
C6151 INVX1_LOC_300/A INVX1_LOC_361/A 0.07fF
C6152 NAND2X1_LOC_712/a_36_24# INVX1_LOC_555/A 0.00fF
C6153 INVX1_LOC_661/A INVX1_LOC_100/Y 0.01fF
C6154 NAND2X1_LOC_557/B INVX1_LOC_35/Y 0.02fF
C6155 INVX1_LOC_145/Y NAND2X1_LOC_759/Y 0.00fF
C6156 INVX1_LOC_93/Y INPUT_1 0.15fF
C6157 INVX1_LOC_267/A INVX1_LOC_50/Y 0.02fF
C6158 INVX1_LOC_381/A INVX1_LOC_280/A 0.01fF
C6159 INVX1_LOC_11/Y INVX1_LOC_154/A 0.06fF
C6160 INVX1_LOC_172/A INVX1_LOC_6/Y 0.07fF
C6161 INVX1_LOC_522/A NAND2X1_LOC_828/a_36_24# 0.00fF
C6162 INVX1_LOC_89/Y NAND2X1_LOC_667/a_36_24# 0.01fF
C6163 INVX1_LOC_677/Y INVX1_LOC_479/A 0.00fF
C6164 INVX1_LOC_105/Y INVX1_LOC_6/Y 0.00fF
C6165 NAND2X1_LOC_827/a_36_24# INVX1_LOC_59/A 0.00fF
C6166 INVX1_LOC_395/A INVX1_LOC_92/A 0.31fF
C6167 INVX1_LOC_93/Y INVX1_LOC_292/Y 0.28fF
C6168 INVX1_LOC_366/Y INVX1_LOC_26/Y 0.01fF
C6169 INVX1_LOC_301/Y INVX1_LOC_370/A 0.06fF
C6170 INVX1_LOC_504/A INVX1_LOC_26/Y 0.07fF
C6171 INVX1_LOC_500/A INVX1_LOC_145/Y 0.06fF
C6172 INVX1_LOC_502/A NAND2X1_LOC_416/Y 0.08fF
C6173 NAND2X1_LOC_486/A NAND2X1_LOC_484/a_36_24# 0.00fF
C6174 INVX1_LOC_633/A NAND2X1_LOC_803/a_36_24# 0.02fF
C6175 INVX1_LOC_80/A NAND2X1_LOC_544/B 0.61fF
C6176 NAND2X1_LOC_274/B NAND2X1_LOC_649/a_36_24# 0.00fF
C6177 INVX1_LOC_35/Y NAND2X1_LOC_66/Y 1.04fF
C6178 NAND2X1_LOC_274/B INVX1_LOC_48/Y 0.03fF
C6179 INVX1_LOC_240/Y INVX1_LOC_242/A 0.00fF
C6180 INVX1_LOC_69/Y NAND2X1_LOC_274/Y 0.12fF
C6181 INVX1_LOC_599/A INVX1_LOC_598/Y 0.00fF
C6182 INVX1_LOC_159/Y INVX1_LOC_79/A 0.75fF
C6183 INVX1_LOC_62/Y INVX1_LOC_504/Y 0.07fF
C6184 INVX1_LOC_6/Y NAND2X1_LOC_846/B 0.08fF
C6185 INVX1_LOC_148/Y INVX1_LOC_491/Y 0.02fF
C6186 INVX1_LOC_210/Y INVX1_LOC_210/A 0.01fF
C6187 INVX1_LOC_58/Y INVX1_LOC_659/A 0.07fF
C6188 INVX1_LOC_54/Y INVX1_LOC_319/A 0.01fF
C6189 NAND2X1_LOC_504/a_36_24# INVX1_LOC_100/Y 0.00fF
C6190 INVX1_LOC_89/Y NAND2X1_LOC_433/Y 0.12fF
C6191 INVX1_LOC_554/A INVX1_LOC_567/A 0.00fF
C6192 INVX1_LOC_211/Y INVX1_LOC_211/A 0.01fF
C6193 INVX1_LOC_31/Y NAND2X1_LOC_123/B 0.07fF
C6194 INVX1_LOC_492/A INVX1_LOC_645/Y 0.24fF
C6195 INVX1_LOC_54/Y NAND2X1_LOC_843/B 0.02fF
C6196 INVX1_LOC_328/Y INVX1_LOC_206/A 0.01fF
C6197 NAND2X1_LOC_615/B INVX1_LOC_666/Y 0.03fF
C6198 INVX1_LOC_444/Y NAND2X1_LOC_416/B 0.03fF
C6199 INVX1_LOC_405/A NAND2X1_LOC_271/B 0.16fF
C6200 INVX1_LOC_54/Y INVX1_LOC_625/Y 0.42fF
C6201 INVX1_LOC_46/Y INVX1_LOC_211/A 0.15fF
C6202 INVX1_LOC_653/Y INVX1_LOC_66/A 0.20fF
C6203 INVX1_LOC_531/Y INVX1_LOC_63/Y 0.07fF
C6204 INVX1_LOC_69/Y NAND2X1_LOC_451/B 9.00fF
C6205 NAND2X1_LOC_301/B INVX1_LOC_242/Y 0.05fF
C6206 INVX1_LOC_31/Y INVX1_LOC_270/Y 0.09fF
C6207 INVX1_LOC_190/A INVX1_LOC_9/Y 0.01fF
C6208 INVX1_LOC_3/Y INVX1_LOC_34/Y 0.03fF
C6209 INVX1_LOC_31/Y INVX1_LOC_92/A 0.07fF
C6210 INVX1_LOC_79/A INVX1_LOC_468/A 0.28fF
C6211 GATE_479 INVX1_LOC_443/A 0.11fF
C6212 VDD INVX1_LOC_607/A 0.18fF
C6213 INVX1_LOC_505/Y INVX1_LOC_461/Y 0.03fF
C6214 INVX1_LOC_100/Y NAND2X1_LOC_372/Y 0.11fF
C6215 INVX1_LOC_51/A INVX1_LOC_578/A 0.04fF
C6216 VDD NAND2X1_LOC_486/B 0.01fF
C6217 INVX1_LOC_41/Y INVX1_LOC_588/A 0.08fF
C6218 INVX1_LOC_591/Y NAND2X1_LOC_759/B 0.00fF
C6219 INVX1_LOC_426/Y INVX1_LOC_596/A 0.04fF
C6220 NAND2X1_LOC_249/Y INVX1_LOC_596/A 0.03fF
C6221 NAND2X1_LOC_24/a_36_24# INVX1_LOC_530/Y 0.00fF
C6222 INVX1_LOC_409/Y NAND2X1_LOC_603/Y 0.01fF
C6223 INVX1_LOC_594/Y INVX1_LOC_675/Y 0.01fF
C6224 INVX1_LOC_288/Y INVX1_LOC_638/A 0.09fF
C6225 NAND2X1_LOC_331/A NAND2X1_LOC_728/B 0.04fF
C6226 INVX1_LOC_203/Y INVX1_LOC_80/A 0.02fF
C6227 VDD INVX1_LOC_673/A -0.00fF
C6228 INVX1_LOC_578/A NAND2X1_LOC_177/a_36_24# 0.00fF
C6229 INVX1_LOC_301/A NAND2X1_LOC_102/a_36_24# 0.01fF
C6230 NAND2X1_LOC_790/B INVX1_LOC_98/Y 0.05fF
C6231 INVX1_LOC_6/Y INVX1_LOC_109/Y 0.01fF
C6232 INVX1_LOC_145/Y INVX1_LOC_596/Y 0.13fF
C6233 NAND2X1_LOC_331/A INVX1_LOC_188/Y 0.00fF
C6234 INVX1_LOC_593/Y NAND2X1_LOC_801/A 0.09fF
C6235 NAND2X1_LOC_79/Y INVX1_LOC_366/A 0.04fF
C6236 VDD INVX1_LOC_492/A 0.58fF
C6237 INVX1_LOC_401/A INVX1_LOC_51/Y 0.03fF
C6238 INVX1_LOC_435/A INVX1_LOC_438/A 0.01fF
C6239 NAND2X1_LOC_475/A INVX1_LOC_35/Y 0.06fF
C6240 NAND2X1_LOC_324/B INVX1_LOC_45/Y 0.03fF
C6241 INVX1_LOC_287/A INVX1_LOC_160/Y 0.00fF
C6242 VDD INVX1_LOC_467/Y 0.29fF
C6243 INVX1_LOC_84/A INVX1_LOC_169/A 0.03fF
C6244 INVX1_LOC_53/Y INVX1_LOC_586/A 0.48fF
C6245 INVX1_LOC_554/A INVX1_LOC_6/Y 0.08fF
C6246 NAND2X1_LOC_45/Y INVX1_LOC_118/A 0.02fF
C6247 INVX1_LOC_21/Y INVX1_LOC_65/Y 0.00fF
C6248 NAND2X1_LOC_534/Y INVX1_LOC_374/Y 0.13fF
C6249 INVX1_LOC_567/A INVX1_LOC_199/Y 0.01fF
C6250 INVX1_LOC_395/A INVX1_LOC_681/Y 0.01fF
C6251 INVX1_LOC_662/Y INVX1_LOC_107/A 0.03fF
C6252 NAND2X1_LOC_791/B INVX1_LOC_285/A 0.03fF
C6253 NAND2X1_LOC_845/a_36_24# INVX1_LOC_600/A 0.00fF
C6254 INVX1_LOC_37/Y INPUT_1 0.01fF
C6255 NAND2X1_LOC_475/A NAND2X1_LOC_448/B 0.02fF
C6256 INVX1_LOC_257/Y INVX1_LOC_46/Y 0.42fF
C6257 INVX1_LOC_384/A NAND2X1_LOC_471/a_36_24# 0.01fF
C6258 INVX1_LOC_412/Y INVX1_LOC_355/Y 0.00fF
C6259 INVX1_LOC_395/A INPUT_1 0.36fF
C6260 NAND2X1_LOC_781/A INVX1_LOC_53/Y 0.01fF
C6261 INVX1_LOC_312/Y INVX1_LOC_53/Y 0.00fF
C6262 INVX1_LOC_384/A NAND2X1_LOC_643/a_36_24# 0.01fF
C6263 INVX1_LOC_678/Y INVX1_LOC_602/Y 0.01fF
C6264 INVX1_LOC_502/Y INVX1_LOC_35/Y 0.03fF
C6265 VDD INVX1_LOC_513/Y 0.46fF
C6266 INVX1_LOC_17/Y INVX1_LOC_526/A 0.01fF
C6267 INVX1_LOC_169/A NAND2X1_LOC_67/Y 0.05fF
C6268 INVX1_LOC_446/Y INVX1_LOC_46/Y 0.07fF
C6269 INVX1_LOC_291/A INVX1_LOC_99/Y 0.07fF
C6270 INVX1_LOC_392/Y INVX1_LOC_50/Y 0.39fF
C6271 INVX1_LOC_65/Y NAND2X1_LOC_267/A 0.08fF
C6272 INVX1_LOC_45/Y INVX1_LOC_110/A 0.01fF
C6273 INVX1_LOC_395/A INVX1_LOC_292/Y 0.01fF
C6274 INPUT_0 INVX1_LOC_49/Y 0.14fF
C6275 NAND2X1_LOC_741/a_36_24# INVX1_LOC_49/Y 0.01fF
C6276 INVX1_LOC_134/A INVX1_LOC_93/Y 0.01fF
C6277 INVX1_LOC_366/Y INVX1_LOC_369/A 0.03fF
C6278 INVX1_LOC_17/Y INVX1_LOC_197/A 0.03fF
C6279 INVX1_LOC_373/A INVX1_LOC_338/Y 0.04fF
C6280 NAND2X1_LOC_391/B INVX1_LOC_117/Y 0.01fF
C6281 INVX1_LOC_21/Y INVX1_LOC_604/Y 0.07fF
C6282 INVX1_LOC_626/A NAND2X1_LOC_677/Y 0.01fF
C6283 NAND2X1_LOC_106/Y INVX1_LOC_51/Y 0.02fF
C6284 INVX1_LOC_448/A NAND2X1_LOC_471/a_36_24# 0.00fF
C6285 INVX1_LOC_360/Y NAND2X1_LOC_299/Y 0.00fF
C6286 NAND2X1_LOC_317/A INVX1_LOC_557/Y 0.01fF
C6287 INVX1_LOC_384/A INVX1_LOC_46/Y 0.02fF
C6288 INPUT_0 INVX1_LOC_642/Y 0.01fF
C6289 INVX1_LOC_35/Y INVX1_LOC_136/Y 0.00fF
C6290 NAND2X1_LOC_516/Y INVX1_LOC_49/Y 0.09fF
C6291 INVX1_LOC_448/A NAND2X1_LOC_643/a_36_24# 0.00fF
C6292 INVX1_LOC_595/Y NAND2X1_LOC_379/Y 0.26fF
C6293 INVX1_LOC_531/A INVX1_LOC_99/Y 0.01fF
C6294 INVX1_LOC_524/Y INVX1_LOC_50/Y 0.18fF
C6295 INVX1_LOC_50/Y INVX1_LOC_59/A 0.53fF
C6296 INVX1_LOC_683/Y INPUT_1 0.02fF
C6297 INVX1_LOC_614/A INVX1_LOC_492/A 0.04fF
C6298 INVX1_LOC_676/Y INVX1_LOC_357/A 0.00fF
C6299 INVX1_LOC_459/A INVX1_LOC_479/A 0.02fF
C6300 NAND2X1_LOC_434/a_36_24# INVX1_LOC_638/A 0.01fF
C6301 INVX1_LOC_378/A NAND2X1_LOC_632/a_36_24# 0.00fF
C6302 INVX1_LOC_395/A INVX1_LOC_399/A 0.47fF
C6303 NAND2X1_LOC_756/Y INVX1_LOC_32/Y 0.13fF
C6304 VDD INVX1_LOC_660/Y 0.01fF
C6305 INVX1_LOC_367/A INVX1_LOC_50/Y 0.03fF
C6306 NAND2X1_LOC_331/A INVX1_LOC_491/A 0.09fF
C6307 NAND2X1_LOC_704/B INVX1_LOC_89/Y 0.34fF
C6308 INVX1_LOC_586/A NAND2X1_LOC_274/Y 0.01fF
C6309 NAND2X1_LOC_791/A NAND2X1_LOC_755/B 0.02fF
C6310 NAND2X1_LOC_755/B INVX1_LOC_145/Y 0.03fF
C6311 INVX1_LOC_45/Y NAND2X1_LOC_275/a_36_24# 0.00fF
C6312 INVX1_LOC_338/A INVX1_LOC_99/Y 0.03fF
C6313 INVX1_LOC_686/A INVX1_LOC_359/Y 0.03fF
C6314 INVX1_LOC_418/Y INVX1_LOC_417/Y 0.00fF
C6315 INVX1_LOC_293/Y INVX1_LOC_32/Y 5.45fF
C6316 INVX1_LOC_385/Y INVX1_LOC_278/Y 0.11fF
C6317 NAND2X1_LOC_79/Y INVX1_LOC_6/Y 0.02fF
C6318 NAND2X1_LOC_669/Y NAND2X1_LOC_720/A 0.01fF
C6319 NAND2X1_LOC_97/A INVX1_LOC_58/Y 0.23fF
C6320 INVX1_LOC_417/Y INVX1_LOC_159/Y 0.07fF
C6321 INVX1_LOC_211/Y INVX1_LOC_145/Y 0.03fF
C6322 INVX1_LOC_126/Y INVX1_LOC_6/Y 0.01fF
C6323 INPUT_7 INPUT_4 0.02fF
C6324 NAND2X1_LOC_673/B INVX1_LOC_7/Y 0.02fF
C6325 NAND2X1_LOC_148/A NAND2X1_LOC_148/B 0.09fF
C6326 NAND2X1_LOC_4/a_36_24# INVX1_LOC_7/Y 0.00fF
C6327 INVX1_LOC_556/Y INVX1_LOC_98/Y 0.17fF
C6328 NAND2X1_LOC_43/Y INVX1_LOC_35/Y 0.01fF
C6329 INVX1_LOC_563/A INVX1_LOC_298/A 0.01fF
C6330 INVX1_LOC_287/A NAND2X1_LOC_267/A 0.14fF
C6331 INVX1_LOC_536/A INVX1_LOC_496/Y 0.01fF
C6332 INVX1_LOC_552/Y INVX1_LOC_531/Y 0.02fF
C6333 INVX1_LOC_254/Y INVX1_LOC_230/A 0.07fF
C6334 INVX1_LOC_278/A INVX1_LOC_62/Y 0.03fF
C6335 INVX1_LOC_53/Y INVX1_LOC_157/Y 0.03fF
C6336 INVX1_LOC_516/A INVX1_LOC_50/Y 0.00fF
C6337 INVX1_LOC_17/Y NAND2X1_LOC_174/B 0.01fF
C6338 INVX1_LOC_12/Y INVX1_LOC_100/A 0.01fF
C6339 INVX1_LOC_199/Y NAND2X1_LOC_820/A 0.02fF
C6340 INVX1_LOC_160/A INVX1_LOC_32/Y 0.00fF
C6341 INVX1_LOC_381/A INVX1_LOC_328/Y 0.08fF
C6342 INVX1_LOC_193/A NAND2X1_LOC_775/B 0.10fF
C6343 INVX1_LOC_549/A INVX1_LOC_479/A 2.20fF
C6344 INVX1_LOC_17/Y NAND2X1_LOC_591/Y 0.01fF
C6345 INVX1_LOC_366/A INVX1_LOC_85/A 0.18fF
C6346 INVX1_LOC_392/A INVX1_LOC_50/Y 0.03fF
C6347 INVX1_LOC_145/Y INVX1_LOC_46/Y 0.46fF
C6348 VDD NAND2X1_LOC_98/B 0.01fF
C6349 INVX1_LOC_159/Y INVX1_LOC_48/Y 0.07fF
C6350 INVX1_LOC_496/A INVX1_LOC_633/Y 0.06fF
C6351 NAND2X1_LOC_635/B INVX1_LOC_505/A 0.00fF
C6352 NAND2X1_LOC_503/a_36_24# INVX1_LOC_26/Y 0.00fF
C6353 INVX1_LOC_17/Y INVX1_LOC_173/Y 0.00fF
C6354 INVX1_LOC_153/A INVX1_LOC_35/Y 0.01fF
C6355 INVX1_LOC_551/Y INVX1_LOC_242/Y 0.10fF
C6356 INVX1_LOC_206/Y NAND2X1_LOC_832/A 0.03fF
C6357 INVX1_LOC_80/A INVX1_LOC_44/Y 0.07fF
C6358 INVX1_LOC_578/A INVX1_LOC_441/A 0.05fF
C6359 NAND2X1_LOC_557/B INVX1_LOC_531/A 0.03fF
C6360 INVX1_LOC_20/Y NAND2X1_LOC_301/B 0.05fF
C6361 NAND2X1_LOC_673/B INVX1_LOC_32/Y 0.03fF
C6362 INVX1_LOC_54/Y INVX1_LOC_361/Y 0.06fF
C6363 NAND2X1_LOC_726/a_36_24# INVX1_LOC_655/A 0.01fF
C6364 NAND2X1_LOC_147/B INVX1_LOC_58/Y 0.01fF
C6365 INVX1_LOC_284/A INVX1_LOC_284/Y 0.05fF
C6366 INVX1_LOC_543/Y INVX1_LOC_198/A 0.03fF
C6367 INVX1_LOC_662/Y NAND2X1_LOC_285/A 0.02fF
C6368 INVX1_LOC_386/Y NAND2X1_LOC_344/B 0.11fF
C6369 INVX1_LOC_442/A INVX1_LOC_666/Y 0.72fF
C6370 NAND2X1_LOC_152/B INVX1_LOC_655/A 0.06fF
C6371 NAND2X1_LOC_396/a_36_24# INVX1_LOC_443/A 0.07fF
C6372 INVX1_LOC_96/A INVX1_LOC_35/Y 0.01fF
C6373 INVX1_LOC_93/Y INVX1_LOC_50/Y 1.38fF
C6374 INVX1_LOC_51/Y INVX1_LOC_329/Y 0.01fF
C6375 NAND2X1_LOC_686/B INVX1_LOC_537/A 0.10fF
C6376 INVX1_LOC_31/Y INPUT_1 0.17fF
C6377 NAND2X1_LOC_296/Y INVX1_LOC_245/A 0.00fF
C6378 INVX1_LOC_586/A NAND2X1_LOC_451/B 8.95fF
C6379 NAND2X1_LOC_482/a_36_24# NAND2X1_LOC_482/Y 0.02fF
C6380 NAND2X1_LOC_694/a_36_24# INVX1_LOC_479/A 0.01fF
C6381 INVX1_LOC_54/Y NAND2X1_LOC_125/a_36_24# 0.06fF
C6382 INVX1_LOC_213/Y INVX1_LOC_69/Y 0.18fF
C6383 INVX1_LOC_387/Y INVX1_LOC_362/A 0.01fF
C6384 INVX1_LOC_361/Y INVX1_LOC_257/A 0.07fF
C6385 INVX1_LOC_449/A INVX1_LOC_100/Y 0.07fF
C6386 NAND2X1_LOC_318/A INVX1_LOC_211/A 0.14fF
C6387 NAND2X1_LOC_403/A INVX1_LOC_9/Y 0.01fF
C6388 INVX1_LOC_586/A NAND2X1_LOC_230/a_36_24# 0.01fF
C6389 INVX1_LOC_49/Y INVX1_LOC_527/Y 0.02fF
C6390 INVX1_LOC_655/Y NAND2X1_LOC_843/B 0.20fF
C6391 INVX1_LOC_625/A INVX1_LOC_26/Y 0.25fF
C6392 INVX1_LOC_598/A NAND2X1_LOC_759/Y 0.06fF
C6393 INVX1_LOC_675/A INVX1_LOC_50/Y 0.07fF
C6394 INVX1_LOC_80/A INVX1_LOC_347/A 0.08fF
C6395 NAND2X1_LOC_179/Y INVX1_LOC_502/A 0.01fF
C6396 INVX1_LOC_172/A INVX1_LOC_206/A 0.04fF
C6397 INVX1_LOC_20/Y INVX1_LOC_291/Y 0.01fF
C6398 INVX1_LOC_658/Y INVX1_LOC_59/A 0.05fF
C6399 NAND2X1_LOC_334/B INVX1_LOC_50/Y 0.02fF
C6400 INVX1_LOC_51/Y INVX1_LOC_92/A 0.12fF
C6401 INVX1_LOC_6/Y INVX1_LOC_199/Y 0.11fF
C6402 INVX1_LOC_294/A INVX1_LOC_26/Y 0.01fF
C6403 NAND2X1_LOC_148/B INVX1_LOC_662/A 0.16fF
C6404 INVX1_LOC_676/Y INVX1_LOC_495/Y 0.09fF
C6405 INVX1_LOC_67/Y INVX1_LOC_74/Y 0.18fF
C6406 NAND2X1_LOC_616/Y INVX1_LOC_483/A 0.00fF
C6407 INVX1_LOC_35/Y NAND2X1_LOC_627/Y 0.01fF
C6408 INVX1_LOC_586/A INVX1_LOC_636/Y 0.01fF
C6409 INVX1_LOC_35/Y INVX1_LOC_475/Y 0.01fF
C6410 INPUT_1 INVX1_LOC_128/A 0.00fF
C6411 INVX1_LOC_62/Y INVX1_LOC_453/Y 0.03fF
C6412 INVX1_LOC_79/A INVX1_LOC_345/A 0.04fF
C6413 INVX1_LOC_208/Y INVX1_LOC_26/Y 0.36fF
C6414 INVX1_LOC_42/Y INVX1_LOC_190/A 0.18fF
C6415 INVX1_LOC_328/Y NAND2X1_LOC_200/a_36_24# 0.01fF
C6416 NAND2X1_LOC_186/a_36_24# INVX1_LOC_491/A 0.00fF
C6417 INVX1_LOC_266/A INVX1_LOC_92/A 0.89fF
C6418 INVX1_LOC_11/Y INVX1_LOC_347/A 0.07fF
C6419 INVX1_LOC_41/Y NAND2X1_LOC_646/A 0.01fF
C6420 INVX1_LOC_479/A INVX1_LOC_230/A 0.19fF
C6421 INVX1_LOC_116/Y INVX1_LOC_666/Y 0.07fF
C6422 INVX1_LOC_62/Y INVX1_LOC_259/Y 0.03fF
C6423 NAND2X1_LOC_86/Y INVX1_LOC_180/Y 0.01fF
C6424 INVX1_LOC_41/Y INVX1_LOC_86/Y 0.00fF
C6425 INVX1_LOC_202/Y INVX1_LOC_211/A 0.02fF
C6426 INVX1_LOC_484/Y INVX1_LOC_486/A 0.09fF
C6427 INVX1_LOC_277/A NAND2X1_LOC_843/B 0.02fF
C6428 INVX1_LOC_653/A INVX1_LOC_69/Y 0.01fF
C6429 INVX1_LOC_452/A INVX1_LOC_443/A 0.18fF
C6430 INVX1_LOC_255/A NAND2X1_LOC_545/A 0.04fF
C6431 INVX1_LOC_326/Y INVX1_LOC_11/A 0.01fF
C6432 INVX1_LOC_253/Y INVX1_LOC_41/Y 0.02fF
C6433 INVX1_LOC_82/Y INVX1_LOC_9/Y 0.19fF
C6434 NAND2X1_LOC_480/a_36_24# INVX1_LOC_244/Y 0.00fF
C6435 INVX1_LOC_100/Y INVX1_LOC_328/Y 0.10fF
C6436 INVX1_LOC_63/Y INVX1_LOC_41/Y 2.67fF
C6437 NAND2X1_LOC_81/Y INVX1_LOC_85/A 0.15fF
C6438 VDD INVX1_LOC_224/Y 1.83fF
C6439 INVX1_LOC_662/A INVX1_LOC_667/A 0.03fF
C6440 INVX1_LOC_347/Y INVX1_LOC_74/Y 0.07fF
C6441 INVX1_LOC_89/Y INVX1_LOC_91/Y 0.03fF
C6442 INVX1_LOC_49/Y INVX1_LOC_464/Y 0.01fF
C6443 INVX1_LOC_424/A INVX1_LOC_446/Y 0.02fF
C6444 VDD INVX1_LOC_578/A -0.00fF
C6445 INVX1_LOC_434/A INVX1_LOC_445/Y 0.03fF
C6446 VDD INVX1_LOC_557/A 0.06fF
C6447 INVX1_LOC_62/Y INVX1_LOC_114/A 0.06fF
C6448 INVX1_LOC_459/A INVX1_LOC_372/Y 0.16fF
C6449 INVX1_LOC_301/A INVX1_LOC_551/Y 0.10fF
C6450 INPUT_0 NAND2X1_LOC_498/B 0.00fF
C6451 INVX1_LOC_570/Y NAND2X1_LOC_152/Y 0.33fF
C6452 INVX1_LOC_188/Y INVX1_LOC_638/A 0.07fF
C6453 INVX1_LOC_567/A INVX1_LOC_53/Y 0.01fF
C6454 NAND2X1_LOC_93/Y INVX1_LOC_524/Y 0.16fF
C6455 INPUT_0 NAND2X1_LOC_339/a_36_24# 0.00fF
C6456 INPUT_0 INVX1_LOC_76/Y 0.18fF
C6457 NAND2X1_LOC_762/a_36_24# INVX1_LOC_6/A 0.00fF
C6458 INVX1_LOC_557/A INVX1_LOC_510/Y 0.07fF
C6459 VDD INVX1_LOC_358/A -0.00fF
C6460 INVX1_LOC_578/A NAND2X1_LOC_124/a_36_24# 0.01fF
C6461 INVX1_LOC_412/Y NAND2X1_LOC_307/A 0.03fF
C6462 INVX1_LOC_51/A INVX1_LOC_686/A 0.02fF
C6463 INVX1_LOC_435/Y INVX1_LOC_235/Y 0.04fF
C6464 VDD INVX1_LOC_568/Y 0.21fF
C6465 INVX1_LOC_118/Y INVX1_LOC_80/A 0.07fF
C6466 NAND2X1_LOC_43/a_36_24# INVX1_LOC_17/Y 0.00fF
C6467 NAND2X1_LOC_543/B INVX1_LOC_35/Y 0.01fF
C6468 NAND2X1_LOC_746/a_36_24# INVX1_LOC_549/Y 0.00fF
C6469 VDD INVX1_LOC_468/Y 0.65fF
C6470 INVX1_LOC_257/Y INVX1_LOC_115/A 0.00fF
C6471 INVX1_LOC_206/Y NAND2X1_LOC_621/a_36_24# 0.00fF
C6472 INVX1_LOC_80/A INVX1_LOC_96/Y 0.07fF
C6473 INVX1_LOC_410/Y INVX1_LOC_99/A -0.05fF
C6474 INVX1_LOC_224/Y INVX1_LOC_158/Y 0.01fF
C6475 INVX1_LOC_20/Y INVX1_LOC_551/Y 0.02fF
C6476 NAND2X1_LOC_299/Y INVX1_LOC_45/Y 0.07fF
C6477 INVX1_LOC_603/A NAND2X1_LOC_76/B 0.00fF
C6478 INVX1_LOC_449/A NAND2X1_LOC_501/a_36_24# 0.00fF
C6479 NAND2X1_LOC_173/Y INVX1_LOC_686/A 0.02fF
C6480 VDD INVX1_LOC_227/Y 0.26fF
C6481 INVX1_LOC_578/A INVX1_LOC_116/A 0.02fF
C6482 INVX1_LOC_679/Y INVX1_LOC_51/Y 0.01fF
C6483 INVX1_LOC_11/Y INVX1_LOC_118/Y 0.01fF
C6484 NAND2X1_LOC_56/Y NAND2X1_LOC_845/a_36_24# 0.00fF
C6485 INVX1_LOC_250/A NAND2X1_LOC_123/A 0.14fF
C6486 NAND2X1_LOC_381/a_36_24# INVX1_LOC_381/A 0.00fF
C6487 INVX1_LOC_438/A INVX1_LOC_93/Y 0.07fF
C6488 INVX1_LOC_319/Y INVX1_LOC_194/Y 0.98fF
C6489 INVX1_LOC_20/Y NAND2X1_LOC_304/a_36_24# -0.00fF
C6490 INVX1_LOC_424/A INVX1_LOC_433/A 0.14fF
C6491 INVX1_LOC_617/Y INVX1_LOC_545/Y 0.05fF
C6492 INVX1_LOC_395/A INVX1_LOC_50/Y 0.27fF
C6493 INVX1_LOC_272/Y INVX1_LOC_53/Y 0.03fF
C6494 NAND2X1_LOC_791/B INVX1_LOC_53/Y 0.26fF
C6495 INVX1_LOC_603/Y INVX1_LOC_398/A 0.07fF
C6496 INVX1_LOC_201/Y INVX1_LOC_273/A 0.18fF
C6497 NAND2X1_LOC_318/A INVX1_LOC_145/Y 0.02fF
C6498 VDD INVX1_LOC_120/Y 0.51fF
C6499 INVX1_LOC_551/Y INVX1_LOC_300/A 0.10fF
C6500 INVX1_LOC_51/Y INVX1_LOC_681/Y 0.01fF
C6501 INVX1_LOC_353/Y INVX1_LOC_116/Y 0.25fF
C6502 INVX1_LOC_580/Y INVX1_LOC_259/Y 0.02fF
C6503 INVX1_LOC_362/Y INVX1_LOC_50/Y 0.03fF
C6504 INVX1_LOC_617/A INVX1_LOC_35/Y 0.04fF
C6505 INVX1_LOC_441/Y INVX1_LOC_93/Y 0.05fF
C6506 NAND2X1_LOC_184/Y INVX1_LOC_45/Y 0.08fF
C6507 INVX1_LOC_536/A INVX1_LOC_676/Y 0.01fF
C6508 INVX1_LOC_51/Y INPUT_1 0.41fF
C6509 NAND2X1_LOC_335/a_36_24# NAND2X1_LOC_267/A 0.01fF
C6510 NAND2X1_LOC_780/A INVX1_LOC_137/Y 0.04fF
C6511 INVX1_LOC_416/A INVX1_LOC_119/A 0.03fF
C6512 INVX1_LOC_80/A NAND2X1_LOC_418/Y 0.27fF
C6513 VDD INVX1_LOC_644/Y 0.26fF
C6514 INVX1_LOC_614/A INVX1_LOC_568/Y 0.01fF
C6515 INVX1_LOC_409/Y INVX1_LOC_652/A 0.06fF
C6516 NAND2X1_LOC_136/a_36_24# INVX1_LOC_50/Y 0.01fF
C6517 NAND2X1_LOC_589/a_36_24# INVX1_LOC_47/Y 0.01fF
C6518 INVX1_LOC_526/A INVX1_LOC_497/Y 0.24fF
C6519 INVX1_LOC_446/Y INVX1_LOC_49/Y 0.07fF
C6520 INVX1_LOC_596/A INVX1_LOC_556/Y 0.01fF
C6521 NAND2X1_LOC_582/a_36_24# NAND2X1_LOC_451/B 0.01fF
C6522 INVX1_LOC_18/A INVX1_LOC_55/Y 0.01fF
C6523 INVX1_LOC_11/Y INVX1_LOC_312/A 0.08fF
C6524 INVX1_LOC_266/A INPUT_1 0.06fF
C6525 NAND2X1_LOC_387/Y INVX1_LOC_398/A 0.01fF
C6526 INVX1_LOC_11/Y NAND2X1_LOC_391/A 0.02fF
C6527 INVX1_LOC_683/Y INVX1_LOC_50/Y 0.02fF
C6528 INVX1_LOC_288/A INVX1_LOC_49/Y 0.07fF
C6529 INVX1_LOC_447/Y INVX1_LOC_442/Y 0.00fF
C6530 INPUT_4 INVX1_LOC_55/Y 0.06fF
C6531 INVX1_LOC_286/Y INVX1_LOC_525/Y 0.01fF
C6532 INVX1_LOC_465/Y INVX1_LOC_479/A 0.04fF
C6533 NAND2X1_LOC_164/Y INVX1_LOC_26/Y 0.41fF
C6534 INVX1_LOC_551/A INVX1_LOC_45/Y 0.00fF
C6535 INVX1_LOC_45/Y INVX1_LOC_498/Y 0.14fF
C6536 INVX1_LOC_17/Y NAND2X1_LOC_179/Y 0.01fF
C6537 INVX1_LOC_93/Y INVX1_LOC_187/A 0.03fF
C6538 INVX1_LOC_133/A NAND2X1_LOC_342/A 0.63fF
C6539 NAND2X1_LOC_148/B NAND2X1_LOC_147/a_36_24# 0.00fF
C6540 NAND2X1_LOC_354/a_36_24# INVX1_LOC_347/Y 0.00fF
C6541 INVX1_LOC_54/Y INVX1_LOC_307/A 0.05fF
C6542 INVX1_LOC_11/Y NAND2X1_LOC_418/Y 0.18fF
C6543 INVX1_LOC_503/A INVX1_LOC_510/A 0.15fF
C6544 INVX1_LOC_384/A INVX1_LOC_49/Y 0.04fF
C6545 INVX1_LOC_468/Y INVX1_LOC_509/A 0.01fF
C6546 INVX1_LOC_81/Y INVX1_LOC_366/Y 0.03fF
C6547 INVX1_LOC_361/Y INVX1_LOC_371/Y 0.01fF
C6548 INVX1_LOC_550/Y INVX1_LOC_145/Y 0.02fF
C6549 INVX1_LOC_555/A NAND2X1_LOC_662/a_36_24# 0.00fF
C6550 INVX1_LOC_413/A NAND2X1_LOC_525/a_36_24# 0.00fF
C6551 INVX1_LOC_254/Y NAND2X1_LOC_72/Y 0.02fF
C6552 NAND2X1_LOC_457/A INVX1_LOC_62/Y 0.03fF
C6553 NAND2X1_LOC_185/a_36_24# INVX1_LOC_491/A 0.00fF
C6554 INVX1_LOC_21/Y INVX1_LOC_86/Y 0.28fF
C6555 INVX1_LOC_54/Y INVX1_LOC_442/Y 0.10fF
C6556 INVX1_LOC_625/A INVX1_LOC_603/A 0.02fF
C6557 INVX1_LOC_662/A INVX1_LOC_516/Y 0.02fF
C6558 NAND2X1_LOC_137/A INVX1_LOC_670/Y 0.00fF
C6559 INVX1_LOC_552/Y INVX1_LOC_41/Y 0.00fF
C6560 INVX1_LOC_53/Y INVX1_LOC_6/Y 2.56fF
C6561 INVX1_LOC_550/A INVX1_LOC_145/Y 0.00fF
C6562 INPUT_7 INVX1_LOC_69/Y 0.09fF
C6563 NAND2X1_LOC_475/A NAND2X1_LOC_71/a_36_24# 0.00fF
C6564 INVX1_LOC_50/Y INVX1_LOC_189/Y 0.03fF
C6565 INVX1_LOC_449/A NAND2X1_LOC_181/A 0.03fF
C6566 INVX1_LOC_435/A INVX1_LOC_117/Y 0.07fF
C6567 INVX1_LOC_374/A INVX1_LOC_41/Y 0.03fF
C6568 INVX1_LOC_266/Y INVX1_LOC_100/Y 0.03fF
C6569 INVX1_LOC_547/Y INVX1_LOC_62/Y 0.27fF
C6570 NAND2X1_LOC_27/a_36_24# INVX1_LOC_178/A 0.00fF
C6571 INVX1_LOC_203/Y INVX1_LOC_91/Y 0.01fF
C6572 INVX1_LOC_381/A INVX1_LOC_224/A 0.04fF
C6573 INVX1_LOC_387/Y INVX1_LOC_145/Y 0.03fF
C6574 INVX1_LOC_20/Y INVX1_LOC_500/A 0.03fF
C6575 INVX1_LOC_53/A INVX1_LOC_31/Y 0.09fF
C6576 INVX1_LOC_270/A INVX1_LOC_242/Y 0.02fF
C6577 INVX1_LOC_651/Y INVX1_LOC_100/Y 0.01fF
C6578 INVX1_LOC_345/A INVX1_LOC_48/Y 0.02fF
C6579 INVX1_LOC_442/Y NAND2X1_LOC_292/Y 0.06fF
C6580 INVX1_LOC_165/Y INVX1_LOC_74/Y 0.19fF
C6581 INVX1_LOC_448/A INVX1_LOC_49/Y 0.04fF
C6582 NAND2X1_LOC_710/A NAND2X1_LOC_274/B 0.02fF
C6583 INVX1_LOC_184/A INVX1_LOC_26/Y 0.28fF
C6584 INVX1_LOC_45/Y INVX1_LOC_75/Y 0.03fF
C6585 INVX1_LOC_21/Y INVX1_LOC_63/Y 6.18fF
C6586 INVX1_LOC_640/Y GATE_811 0.00fF
C6587 INVX1_LOC_266/Y INVX1_LOC_74/Y 0.03fF
C6588 NAND2X1_LOC_274/B NAND2X1_LOC_541/B 0.04fF
C6589 INVX1_LOC_31/Y INVX1_LOC_50/Y 1.64fF
C6590 INVX1_LOC_49/Y INVX1_LOC_145/Y 0.45fF
C6591 INVX1_LOC_482/A INVX1_LOC_62/Y 0.02fF
C6592 INVX1_LOC_341/Y INVX1_LOC_342/A 0.01fF
C6593 INVX1_LOC_98/A INVX1_LOC_211/A 0.00fF
C6594 INVX1_LOC_267/A INVX1_LOC_117/Y 0.01fF
C6595 NAND2X1_LOC_274/B INVX1_LOC_383/Y 0.01fF
C6596 INVX1_LOC_84/A INVX1_LOC_531/Y 0.11fF
C6597 INVX1_LOC_361/Y INVX1_LOC_89/Y 0.03fF
C6598 INVX1_LOC_89/Y NAND2X1_LOC_333/B 0.07fF
C6599 INVX1_LOC_43/A INVX1_LOC_6/Y 0.01fF
C6600 INPUT_4 INVX1_LOC_18/Y 0.01fF
C6601 NAND2X1_LOC_389/a_36_24# INVX1_LOC_31/Y 0.01fF
C6602 INVX1_LOC_662/A INVX1_LOC_241/Y 0.03fF
C6603 INVX1_LOC_604/Y INVX1_LOC_26/Y 0.01fF
C6604 NAND2X1_LOC_619/Y INVX1_LOC_484/A 0.01fF
C6605 INVX1_LOC_76/Y INVX1_LOC_211/A 0.00fF
C6606 INVX1_LOC_86/Y INVX1_LOC_181/Y 0.01fF
C6607 INVX1_LOC_93/Y NAND2X1_LOC_388/A 0.09fF
C6608 NAND2X1_LOC_313/a_36_24# INVX1_LOC_47/Y 0.01fF
C6609 INVX1_LOC_35/Y NAND2X1_LOC_445/a_36_24# 0.00fF
C6610 INVX1_LOC_194/A INVX1_LOC_9/Y 0.03fF
C6611 INVX1_LOC_42/Y INVX1_LOC_82/Y 0.01fF
C6612 NAND2X1_LOC_542/A NAND2X1_LOC_659/a_36_24# 0.00fF
C6613 INVX1_LOC_686/A INVX1_LOC_354/A 0.01fF
C6614 INVX1_LOC_686/A INVX1_LOC_441/A 0.03fF
C6615 INVX1_LOC_45/Y NAND2X1_LOC_271/A 0.07fF
C6616 INVX1_LOC_35/Y INVX1_LOC_353/A 0.34fF
C6617 INVX1_LOC_63/Y NAND2X1_LOC_267/A 0.12fF
C6618 INVX1_LOC_25/Y INVX1_LOC_657/A 0.01fF
C6619 INVX1_LOC_444/Y INVX1_LOC_244/Y 0.14fF
C6620 INVX1_LOC_469/Y INVX1_LOC_347/Y 0.02fF
C6621 INVX1_LOC_20/Y INVX1_LOC_634/Y 0.04fF
C6622 NAND2X1_LOC_137/A INVX1_LOC_63/Y 0.00fF
C6623 INVX1_LOC_6/Y NAND2X1_LOC_274/Y 0.01fF
C6624 INVX1_LOC_513/A INVX1_LOC_245/A 0.03fF
C6625 INVX1_LOC_145/Y INVX1_LOC_210/A 0.01fF
C6626 INVX1_LOC_145/Y INVX1_LOC_17/A 0.01fF
C6627 INVX1_LOC_209/A INVX1_LOC_79/A 0.27fF
C6628 INVX1_LOC_128/A INVX1_LOC_50/Y 0.00fF
C6629 INVX1_LOC_141/Y INVX1_LOC_49/Y 0.01fF
C6630 INVX1_LOC_47/Y NAND2X1_LOC_686/B 0.02fF
C6631 NAND2X1_LOC_586/Y INVX1_LOC_497/A 0.13fF
C6632 INVX1_LOC_319/A INVX1_LOC_194/Y 0.00fF
C6633 INVX1_LOC_59/Y INVX1_LOC_203/A 0.01fF
C6634 INVX1_LOC_74/Y INVX1_LOC_352/A 0.01fF
C6635 INVX1_LOC_17/Y INVX1_LOC_66/Y 0.01fF
C6636 INVX1_LOC_172/A INVX1_LOC_100/Y 0.02fF
C6637 INVX1_LOC_194/A INVX1_LOC_62/Y 0.01fF
C6638 INVX1_LOC_242/Y INVX1_LOC_46/Y 0.06fF
C6639 NAND2X1_LOC_300/a_36_24# INVX1_LOC_376/Y 0.00fF
C6640 NAND2X1_LOC_313/a_36_24# INVX1_LOC_119/Y 0.00fF
C6641 INVX1_LOC_47/Y INVX1_LOC_223/Y 0.00fF
C6642 INVX1_LOC_620/A INVX1_LOC_353/A 0.23fF
C6643 INVX1_LOC_107/Y INVX1_LOC_63/Y 0.37fF
C6644 NAND2X1_LOC_557/B INVX1_LOC_223/Y 0.11fF
C6645 INVX1_LOC_280/A INVX1_LOC_48/Y 0.03fF
C6646 INVX1_LOC_557/Y INVX1_LOC_199/Y 0.04fF
C6647 NAND2X1_LOC_605/a_36_24# INVX1_LOC_634/Y 0.00fF
C6648 VDD NAND2X1_LOC_86/Y 0.25fF
C6649 INVX1_LOC_361/Y NAND2X1_LOC_544/B 0.03fF
C6650 NAND2X1_LOC_844/a_36_24# INVX1_LOC_6/Y 0.00fF
C6651 INVX1_LOC_69/Y NAND2X1_LOC_545/A 0.99fF
C6652 INVX1_LOC_282/A INVX1_LOC_443/A 0.03fF
C6653 NAND2X1_LOC_503/Y INVX1_LOC_211/A 0.03fF
C6654 INVX1_LOC_347/Y INVX1_LOC_79/A 0.02fF
C6655 INVX1_LOC_100/Y NAND2X1_LOC_846/B 0.02fF
C6656 NAND2X1_LOC_836/B INVX1_LOC_41/Y 0.05fF
C6657 INVX1_LOC_117/Y NAND2X1_LOC_227/A 0.06fF
C6658 INVX1_LOC_69/Y INVX1_LOC_653/Y 0.01fF
C6659 INVX1_LOC_328/Y INVX1_LOC_79/A 0.03fF
C6660 INVX1_LOC_395/A INVX1_LOC_275/A 0.07fF
C6661 INVX1_LOC_148/Y INVX1_LOC_149/Y 0.03fF
C6662 NAND2X1_LOC_45/Y INVX1_LOC_447/A 0.03fF
C6663 INVX1_LOC_69/Y INVX1_LOC_666/Y 0.03fF
C6664 VDD INVX1_LOC_206/Y 4.10fF
C6665 INVX1_LOC_446/A NAND2X1_LOC_735/a_36_24# 0.01fF
C6666 INVX1_LOC_479/A INVX1_LOC_168/Y 0.09fF
C6667 INVX1_LOC_482/Y INVX1_LOC_388/A 0.00fF
C6668 VDD INVX1_LOC_648/Y 0.26fF
C6669 INVX1_LOC_206/Y NAND2X1_LOC_596/Y 0.28fF
C6670 INVX1_LOC_301/A INVX1_LOC_418/A 0.08fF
C6671 INVX1_LOC_320/A INVX1_LOC_109/Y 0.01fF
C6672 INVX1_LOC_438/A INVX1_LOC_395/A 0.10fF
C6673 INVX1_LOC_206/Y INVX1_LOC_228/Y 0.03fF
C6674 INVX1_LOC_584/A INVX1_LOC_540/Y 0.08fF
C6675 INVX1_LOC_44/Y INVX1_LOC_91/Y 0.01fF
C6676 INVX1_LOC_26/Y INVX1_LOC_588/A 0.03fF
C6677 INVX1_LOC_242/Y INVX1_LOC_75/A 0.02fF
C6678 NAND2X1_LOC_276/A NAND2X1_LOC_271/A 0.06fF
C6679 INPUT_0 INVX1_LOC_139/A 0.56fF
C6680 VDD INVX1_LOC_143/Y 0.21fF
C6681 NAND2X1_LOC_234/Y INVX1_LOC_273/Y 0.01fF
C6682 VDD INVX1_LOC_396/Y 0.34fF
C6683 VDD INVX1_LOC_242/A 0.12fF
C6684 INVX1_LOC_20/Y INVX1_LOC_596/Y 0.01fF
C6685 NAND2X1_LOC_373/Y INVX1_LOC_551/Y 0.03fF
C6686 INVX1_LOC_301/A INVX1_LOC_270/A 0.03fF
C6687 INVX1_LOC_65/Y INVX1_LOC_560/A 0.07fF
C6688 NAND2X1_LOC_475/A NAND2X1_LOC_315/a_36_24# 0.00fF
C6689 INVX1_LOC_257/Y INVX1_LOC_76/Y 0.07fF
C6690 INVX1_LOC_145/Y INVX1_LOC_297/Y 0.03fF
C6691 VDD INVX1_LOC_686/A 0.00fF
C6692 INVX1_LOC_446/A INVX1_LOC_21/Y 0.07fF
C6693 INVX1_LOC_347/A INVX1_LOC_625/Y 0.07fF
C6694 NAND2X1_LOC_88/B NAND2X1_LOC_88/a_36_24# 0.00fF
C6695 VDD INVX1_LOC_80/Y 0.24fF
C6696 INVX1_LOC_446/Y INVX1_LOC_76/Y 0.02fF
C6697 INVX1_LOC_625/A NAND2X1_LOC_790/B 0.02fF
C6698 VDD INVX1_LOC_609/Y 0.21fF
C6699 INVX1_LOC_20/Y INVX1_LOC_416/Y 0.01fF
C6700 INVX1_LOC_547/A INVX1_LOC_547/Y 0.07fF
C6701 NAND2X1_LOC_781/B INVX1_LOC_35/Y 0.32fF
C6702 NAND2X1_LOC_486/B INVX1_LOC_45/Y 0.04fF
C6703 NAND2X1_LOC_394/a_36_24# INVX1_LOC_35/Y 0.01fF
C6704 INVX1_LOC_193/Y NAND2X1_LOC_336/B 0.02fF
C6705 VDD INVX1_LOC_14/A 0.00fF
C6706 INVX1_LOC_449/A INVX1_LOC_414/A 0.03fF
C6707 INVX1_LOC_20/Y INVX1_LOC_558/A 0.07fF
C6708 NAND2X1_LOC_710/B INVX1_LOC_670/Y 0.02fF
C6709 INVX1_LOC_510/Y INVX1_LOC_242/A 0.10fF
C6710 NAND2X1_LOC_307/A INVX1_LOC_375/A 0.68fF
C6711 INVX1_LOC_545/Y INVX1_LOC_375/A 0.00fF
C6712 VDD INVX1_LOC_452/A 0.22fF
C6713 INVX1_LOC_266/A INVX1_LOC_134/A 0.07fF
C6714 INVX1_LOC_395/A NAND2X1_LOC_513/A 0.07fF
C6715 NAND2X1_LOC_307/A INVX1_LOC_546/A 0.03fF
C6716 NAND2X1_LOC_68/a_36_24# INVX1_LOC_54/Y 0.00fF
C6717 INVX1_LOC_540/Y INVX1_LOC_537/A 0.01fF
C6718 INVX1_LOC_17/Y INVX1_LOC_412/Y 0.04fF
C6719 INPUT_0 INVX1_LOC_7/Y 0.00fF
C6720 INPUT_0 INVX1_LOC_228/A 0.01fF
C6721 INVX1_LOC_142/A INVX1_LOC_522/Y 0.02fF
C6722 INVX1_LOC_20/Y INVX1_LOC_287/Y 0.01fF
C6723 INVX1_LOC_679/Y NAND2X1_LOC_108/Y 0.01fF
C6724 NAND2X1_LOC_122/Y INVX1_LOC_197/A 0.28fF
C6725 INVX1_LOC_191/Y INVX1_LOC_195/Y 0.05fF
C6726 INVX1_LOC_192/Y INVX1_LOC_230/A 0.05fF
C6727 INVX1_LOC_20/Y INVX1_LOC_270/A 0.03fF
C6728 INVX1_LOC_446/Y INVX1_LOC_386/Y 0.07fF
C6729 INVX1_LOC_301/A INVX1_LOC_46/Y 0.08fF
C6730 INVX1_LOC_584/Y INVX1_LOC_491/Y 0.23fF
C6731 NAND2X1_LOC_744/a_36_24# INVX1_LOC_48/Y 0.00fF
C6732 VDD INVX1_LOC_342/A 0.05fF
C6733 INVX1_LOC_203/Y NAND2X1_LOC_333/B 0.05fF
C6734 INVX1_LOC_416/A INVX1_LOC_410/Y 0.06fF
C6735 INVX1_LOC_12/Y INVX1_LOC_666/A 0.00fF
C6736 INVX1_LOC_405/A NAND2X1_LOC_518/a_36_24# 0.00fF
C6737 INVX1_LOC_602/A INVX1_LOC_59/A 0.18fF
C6738 INVX1_LOC_100/Y INVX1_LOC_109/Y 0.03fF
C6739 INVX1_LOC_438/A INVX1_LOC_31/Y 0.07fF
C6740 INVX1_LOC_400/Y NAND2X1_LOC_775/B 0.07fF
C6741 INVX1_LOC_80/A INVX1_LOC_126/A 0.07fF
C6742 INVX1_LOC_375/A NAND2X1_LOC_600/a_36_24# 0.00fF
C6743 NAND2X1_LOC_379/Y INVX1_LOC_311/Y 0.19fF
C6744 INVX1_LOC_386/Y INVX1_LOC_384/A 0.07fF
C6745 INVX1_LOC_492/A INVX1_LOC_185/Y 1.99fF
C6746 INPUT_0 INVX1_LOC_32/Y 0.07fF
C6747 INVX1_LOC_68/Y INVX1_LOC_35/Y 0.01fF
C6748 INVX1_LOC_76/Y INVX1_LOC_145/Y 0.11fF
C6749 INVX1_LOC_20/Y NAND2X1_LOC_755/B 0.03fF
C6750 VDD NAND2X1_LOC_334/A 0.20fF
C6751 NAND2X1_LOC_786/B NAND2X1_LOC_86/Y 0.36fF
C6752 INVX1_LOC_300/A INVX1_LOC_287/Y 0.02fF
C6753 NAND2X1_LOC_174/B NAND2X1_LOC_122/Y 0.03fF
C6754 INVX1_LOC_188/Y INVX1_LOC_134/Y 0.07fF
C6755 INVX1_LOC_206/Y INVX1_LOC_346/A 0.03fF
C6756 INVX1_LOC_617/Y INVX1_LOC_503/A 0.01fF
C6757 INVX1_LOC_300/A INVX1_LOC_270/A 0.00fF
C6758 NAND2X1_LOC_152/B INVX1_LOC_567/Y 0.06fF
C6759 NAND2X1_LOC_261/Y INVX1_LOC_282/A 0.00fF
C6760 NAND2X1_LOC_704/a_36_24# INVX1_LOC_47/Y 0.00fF
C6761 INVX1_LOC_51/Y INVX1_LOC_50/Y 0.34fF
C6762 INVX1_LOC_590/Y INVX1_LOC_32/Y 0.02fF
C6763 INVX1_LOC_20/Y INVX1_LOC_211/Y 0.02fF
C6764 NAND2X1_LOC_591/Y NAND2X1_LOC_122/Y 0.21fF
C6765 INVX1_LOC_412/A INVX1_LOC_257/A 0.14fF
C6766 INVX1_LOC_554/A INVX1_LOC_100/Y 0.03fF
C6767 NAND2X1_LOC_690/Y INVX1_LOC_496/Y 0.01fF
C6768 INVX1_LOC_286/A INVX1_LOC_32/Y 0.01fF
C6769 INVX1_LOC_12/Y NAND2X1_LOC_72/Y 0.01fF
C6770 INVX1_LOC_405/A INVX1_LOC_41/Y 0.56fF
C6771 INVX1_LOC_80/A INVX1_LOC_252/Y 0.10fF
C6772 INVX1_LOC_266/A INVX1_LOC_50/Y 0.00fF
C6773 NAND2X1_LOC_475/A NAND2X1_LOC_474/a_36_24# 0.00fF
C6774 INVX1_LOC_681/A INVX1_LOC_12/Y 0.02fF
C6775 INVX1_LOC_340/Y INVX1_LOC_340/A 0.10fF
C6776 NAND2X1_LOC_743/a_36_24# INVX1_LOC_54/Y 0.00fF
C6777 NAND2X1_LOC_188/a_36_24# INVX1_LOC_47/Y 0.01fF
C6778 INVX1_LOC_20/Y INVX1_LOC_46/Y 0.03fF
C6779 INVX1_LOC_12/Y NAND2X1_LOC_673/A 0.07fF
C6780 NAND2X1_LOC_383/Y INVX1_LOC_6/Y 0.01fF
C6781 NAND2X1_LOC_184/Y INVX1_LOC_293/Y 0.07fF
C6782 NAND2X1_LOC_130/Y INVX1_LOC_35/Y 0.03fF
C6783 INVX1_LOC_35/Y INVX1_LOC_600/A 0.12fF
C6784 NAND2X1_LOC_336/B INVX1_LOC_54/Y 0.15fF
C6785 INVX1_LOC_300/A NAND2X1_LOC_755/B 0.00fF
C6786 INVX1_LOC_117/Y INVX1_LOC_367/A 0.07fF
C6787 INVX1_LOC_560/Y INVX1_LOC_41/Y 0.03fF
C6788 INVX1_LOC_386/Y INVX1_LOC_145/Y 0.03fF
C6789 INVX1_LOC_513/Y INVX1_LOC_45/Y 0.01fF
C6790 INVX1_LOC_122/Y INVX1_LOC_519/Y 0.02fF
C6791 INVX1_LOC_103/Y INVX1_LOC_686/A 0.01fF
C6792 INVX1_LOC_449/A INVX1_LOC_48/Y 0.07fF
C6793 VDD NAND2X1_LOC_609/B 0.09fF
C6794 INVX1_LOC_602/A INVX1_LOC_93/Y 0.00fF
C6795 NAND2X1_LOC_704/a_36_24# INVX1_LOC_119/Y 0.00fF
C6796 NAND2X1_LOC_332/B INVX1_LOC_49/Y 0.07fF
C6797 INVX1_LOC_353/Y INVX1_LOC_69/Y 0.00fF
C6798 INVX1_LOC_211/Y INVX1_LOC_300/A 0.01fF
C6799 INVX1_LOC_99/Y NAND2X1_LOC_606/Y 0.01fF
C6800 INVX1_LOC_69/Y INVX1_LOC_55/Y 0.04fF
C6801 INVX1_LOC_411/A INVX1_LOC_99/Y 0.12fF
C6802 INVX1_LOC_11/Y INVX1_LOC_252/Y 0.03fF
C6803 INVX1_LOC_206/Y INVX1_LOC_635/Y 0.03fF
C6804 INVX1_LOC_357/A INVX1_LOC_505/A 0.19fF
C6805 INVX1_LOC_53/A INVX1_LOC_40/Y 0.03fF
C6806 NAND2X1_LOC_193/a_36_24# INVX1_LOC_211/A 0.01fF
C6807 INVX1_LOC_117/Y INVX1_LOC_516/A 0.02fF
C6808 INVX1_LOC_675/A INVX1_LOC_111/A 0.02fF
C6809 NAND2X1_LOC_123/A INVX1_LOC_32/Y 0.01fF
C6810 INVX1_LOC_117/Y INVX1_LOC_669/Y 0.03fF
C6811 NAND2X1_LOC_107/Y INVX1_LOC_6/Y 0.73fF
C6812 NAND2X1_LOC_391/B INVX1_LOC_245/A 0.01fF
C6813 NAND2X1_LOC_829/Y INVX1_LOC_69/Y 0.03fF
C6814 INVX1_LOC_375/A NAND2X1_LOC_602/a_36_24# 0.00fF
C6815 NAND2X1_LOC_527/a_36_24# INVX1_LOC_234/Y 0.00fF
C6816 INVX1_LOC_400/A INVX1_LOC_117/Y 0.07fF
C6817 INVX1_LOC_300/A INVX1_LOC_46/Y 0.03fF
C6818 INVX1_LOC_69/Y INVX1_LOC_97/Y 0.00fF
C6819 INVX1_LOC_586/A NAND2X1_LOC_545/A 0.02fF
C6820 NAND2X1_LOC_318/A INVX1_LOC_242/Y 0.01fF
C6821 NAND2X1_LOC_444/A INVX1_LOC_98/Y 0.39fF
C6822 INVX1_LOC_291/A INVX1_LOC_353/A 0.12fF
C6823 INVX1_LOC_556/Y INVX1_LOC_520/A 0.00fF
C6824 INVX1_LOC_12/Y INVX1_LOC_351/Y 0.02fF
C6825 INVX1_LOC_48/Y INVX1_LOC_186/Y 0.18fF
C6826 NAND2X1_LOC_32/Y INVX1_LOC_43/A 0.08fF
C6827 INVX1_LOC_662/A NAND2X1_LOC_820/A 0.05fF
C6828 NAND2X1_LOC_840/a_36_24# INVX1_LOC_664/A 0.00fF
C6829 INVX1_LOC_35/Y INVX1_LOC_484/A 0.01fF
C6830 INVX1_LOC_100/Y NAND2X1_LOC_698/a_36_24# 0.00fF
C6831 INVX1_LOC_32/Y INVX1_LOC_527/Y 0.01fF
C6832 INVX1_LOC_53/Y INVX1_LOC_557/Y 0.05fF
C6833 INVX1_LOC_198/A NAND2X1_LOC_204/a_36_24# 0.00fF
C6834 NAND2X1_LOC_387/Y NAND2X1_LOC_165/Y 0.02fF
C6835 INVX1_LOC_230/A INVX1_LOC_296/A 0.03fF
C6836 INVX1_LOC_607/Y NAND2X1_LOC_286/A 0.04fF
C6837 INVX1_LOC_93/Y INVX1_LOC_117/Y 0.42fF
C6838 INVX1_LOC_134/Y INVX1_LOC_491/A 0.04fF
C6839 INVX1_LOC_129/A INVX1_LOC_411/Y 0.01fF
C6840 INVX1_LOC_444/Y INVX1_LOC_63/Y 0.03fF
C6841 INVX1_LOC_586/A INVX1_LOC_666/Y 0.03fF
C6842 INVX1_LOC_439/Y INVX1_LOC_6/Y 2.52fF
C6843 INVX1_LOC_662/Y NAND2X1_LOC_342/A 0.09fF
C6844 NAND2X1_LOC_427/Y INVX1_LOC_74/Y 0.03fF
C6845 INVX1_LOC_49/Y INVX1_LOC_503/Y 0.05fF
C6846 NAND2X1_LOC_710/A INVX1_LOC_468/A 0.01fF
C6847 INVX1_LOC_578/Y INVX1_LOC_89/Y 0.01fF
C6848 INVX1_LOC_84/A INVX1_LOC_41/Y 0.06fF
C6849 INVX1_LOC_47/Y INVX1_LOC_295/Y 0.01fF
C6850 INVX1_LOC_193/A NAND2X1_LOC_111/Y 0.06fF
C6851 INVX1_LOC_54/Y NAND2X1_LOC_803/a_36_24# 0.00fF
C6852 INVX1_LOC_342/Y INVX1_LOC_300/Y 0.18fF
C6853 NAND2X1_LOC_834/a_36_24# INVX1_LOC_655/A 0.02fF
C6854 INVX1_LOC_166/A NAND2X1_LOC_532/Y 0.00fF
C6855 INVX1_LOC_20/Y INVX1_LOC_75/A 0.01fF
C6856 INVX1_LOC_31/Y NAND2X1_LOC_388/A 0.05fF
C6857 INVX1_LOC_347/Y INVX1_LOC_48/Y 0.03fF
C6858 INVX1_LOC_17/Y INVX1_LOC_664/A 0.07fF
C6859 INVX1_LOC_293/Y INVX1_LOC_75/Y 0.07fF
C6860 NAND2X1_LOC_294/Y NAND2X1_LOC_346/B 0.02fF
C6861 INVX1_LOC_117/Y INVX1_LOC_675/A 0.07fF
C6862 INVX1_LOC_493/A INVX1_LOC_494/Y 0.20fF
C6863 INVX1_LOC_69/Y INVX1_LOC_18/Y 0.24fF
C6864 INVX1_LOC_202/Y INVX1_LOC_242/Y 0.01fF
C6865 INVX1_LOC_578/Y INVX1_LOC_501/A 0.03fF
C6866 INVX1_LOC_79/A INVX1_LOC_352/A 0.01fF
C6867 NAND2X1_LOC_657/a_36_24# INVX1_LOC_510/A 0.01fF
C6868 INVX1_LOC_89/Y INVX1_LOC_532/Y 0.21fF
C6869 INVX1_LOC_328/Y INVX1_LOC_48/Y 0.03fF
C6870 INVX1_LOC_534/Y INVX1_LOC_514/A 0.00fF
C6871 INVX1_LOC_117/Y INVX1_LOC_390/A 0.09fF
C6872 NAND2X1_LOC_720/A INVX1_LOC_272/A 0.08fF
C6873 INVX1_LOC_544/Y INVX1_LOC_6/Y 0.01fF
C6874 INVX1_LOC_26/Y INVX1_LOC_86/Y 0.01fF
C6875 INVX1_LOC_172/A INVX1_LOC_79/A 0.02fF
C6876 INVX1_LOC_46/Y INVX1_LOC_655/A 0.02fF
C6877 INVX1_LOC_662/A INVX1_LOC_6/Y 0.08fF
C6878 INVX1_LOC_342/Y INVX1_LOC_660/A 0.01fF
C6879 INVX1_LOC_300/A INVX1_LOC_75/A 0.00fF
C6880 NAND2X1_LOC_607/a_36_24# NAND2X1_LOC_609/B 0.00fF
C6881 INVX1_LOC_587/Y INVX1_LOC_62/Y 0.03fF
C6882 NAND2X1_LOC_152/B INVX1_LOC_92/A 0.97fF
C6883 INVX1_LOC_137/Y INVX1_LOC_479/A 0.19fF
C6884 INVX1_LOC_513/A NAND2X1_LOC_597/Y 0.01fF
C6885 INVX1_LOC_53/Y INVX1_LOC_636/A 0.07fF
C6886 INVX1_LOC_49/Y INVX1_LOC_242/Y 0.03fF
C6887 INVX1_LOC_48/Y INVX1_LOC_597/Y 0.02fF
C6888 INVX1_LOC_63/Y INVX1_LOC_26/Y 1.16fF
C6889 INVX1_LOC_100/Y INVX1_LOC_199/Y 1.42fF
C6890 NAND2X1_LOC_165/Y INVX1_LOC_91/A 0.03fF
C6891 INVX1_LOC_426/A INVX1_LOC_438/A 0.06fF
C6892 INVX1_LOC_32/Y INVX1_LOC_211/A 0.10fF
C6893 INVX1_LOC_523/Y NAND2X1_LOC_843/B -0.00fF
C6894 INVX1_LOC_49/Y INVX1_LOC_487/A 0.02fF
C6895 INVX1_LOC_32/Y INVX1_LOC_464/Y 0.41fF
C6896 INVX1_LOC_41/Y INVX1_LOC_496/A 0.00fF
C6897 INVX1_LOC_199/Y INVX1_LOC_74/Y 0.12fF
C6898 INVX1_LOC_507/Y INVX1_LOC_475/Y 0.05fF
C6899 NAND2X1_LOC_824/a_36_24# INVX1_LOC_621/A 0.00fF
C6900 INVX1_LOC_659/A INVX1_LOC_657/Y 0.03fF
C6901 INVX1_LOC_79/A INVX1_LOC_224/A 0.01fF
C6902 INVX1_LOC_58/Y INVX1_LOC_241/A 0.00fF
C6903 INVX1_LOC_62/Y INVX1_LOC_9/Y 0.26fF
C6904 VDD INVX1_LOC_390/Y 0.22fF
C6905 VDD INVX1_LOC_290/Y 0.30fF
C6906 INVX1_LOC_13/Y INVX1_LOC_9/Y 0.01fF
C6907 INVX1_LOC_418/A NAND2X1_LOC_373/Y 0.08fF
C6908 INVX1_LOC_26/Y NAND2X1_LOC_214/a_36_24# 0.00fF
C6909 VDD INVX1_LOC_94/A 0.00fF
C6910 VDD INVX1_LOC_4/Y 0.21fF
C6911 INVX1_LOC_438/A INVX1_LOC_51/Y 0.07fF
C6912 INVX1_LOC_224/Y INVX1_LOC_45/Y 0.03fF
C6913 INVX1_LOC_447/A INVX1_LOC_502/Y 0.09fF
C6914 INVX1_LOC_619/A NAND2X1_LOC_86/Y 0.02fF
C6915 VDD INVX1_LOC_654/A 0.26fF
C6916 INVX1_LOC_24/A INVX1_LOC_51/Y 0.04fF
C6917 NAND2X1_LOC_406/B INVX1_LOC_636/A 0.03fF
C6918 INVX1_LOC_578/A INVX1_LOC_45/Y 0.07fF
C6919 NAND2X1_LOC_526/Y INVX1_LOC_428/A 0.00fF
C6920 INVX1_LOC_490/Y INVX1_LOC_586/A 0.53fF
C6921 NAND2X1_LOC_16/Y INVX1_LOC_586/A 0.10fF
C6922 INVX1_LOC_224/Y INPUT_3 0.01fF
C6923 INPUT_0 INVX1_LOC_229/Y 0.01fF
C6924 INVX1_LOC_21/Y INVX1_LOC_560/Y 0.09fF
C6925 NAND2X1_LOC_531/a_36_24# INVX1_LOC_99/Y 0.01fF
C6926 NAND2X1_LOC_753/a_36_24# INVX1_LOC_50/Y 0.00fF
C6927 INVX1_LOC_84/A NAND2X1_LOC_362/a_36_24# 0.00fF
C6928 INVX1_LOC_259/Y INVX1_LOC_638/A 0.00fF
C6929 INVX1_LOC_12/Y NAND2X1_LOC_749/Y 0.34fF
C6930 NAND2X1_LOC_543/B INVX1_LOC_350/A 0.01fF
C6931 INVX1_LOC_607/A INVX1_LOC_293/Y 0.02fF
C6932 INVX1_LOC_413/Y NAND2X1_LOC_523/B 0.27fF
C6933 INPUT_7 INVX1_LOC_1/A 0.01fF
C6934 INVX1_LOC_353/Y INVX1_LOC_586/A 0.02fF
C6935 NAND2X1_LOC_249/Y NAND2X1_LOC_250/Y 0.03fF
C6936 INVX1_LOC_409/Y INVX1_LOC_360/A 0.00fF
C6937 INVX1_LOC_601/A NAND2X1_LOC_223/a_36_24# 0.00fF
C6938 INVX1_LOC_68/Y INVX1_LOC_291/A 0.52fF
C6939 INVX1_LOC_454/A INVX1_LOC_656/Y 0.10fF
C6940 INVX1_LOC_442/A NAND2X1_LOC_804/a_36_24# 0.01fF
C6941 VDD INVX1_LOC_56/Y 0.21fF
C6942 INVX1_LOC_73/Y INVX1_LOC_46/Y 0.01fF
C6943 INVX1_LOC_33/A INVX1_LOC_595/A 0.02fF
C6944 INVX1_LOC_20/Y NAND2X1_LOC_318/A 0.04fF
C6945 INVX1_LOC_410/Y INVX1_LOC_503/A 0.09fF
C6946 INVX1_LOC_69/Y INVX1_LOC_615/A 0.00fF
C6947 INVX1_LOC_418/A NAND2X1_LOC_524/a_36_24# 0.00fF
C6948 INVX1_LOC_446/Y INVX1_LOC_7/Y 0.07fF
C6949 INVX1_LOC_45/Y INVX1_LOC_358/A 0.27fF
C6950 INVX1_LOC_51/Y NAND2X1_LOC_513/A 0.02fF
C6951 NAND2X1_LOC_763/Y INVX1_LOC_48/Y 0.02fF
C6952 INVX1_LOC_586/A INVX1_LOC_97/Y 0.00fF
C6953 NAND2X1_LOC_558/B INVX1_LOC_109/Y 0.05fF
C6954 NAND2X1_LOC_475/A INVX1_LOC_295/Y 0.36fF
C6955 NAND2X1_LOC_45/Y NAND2X1_LOC_706/B 0.04fF
C6956 NAND2X1_LOC_356/a_36_24# INVX1_LOC_290/A 0.02fF
C6957 INVX1_LOC_259/A INVX1_LOC_99/Y 0.04fF
C6958 INVX1_LOC_173/A INVX1_LOC_99/Y 0.01fF
C6959 INVX1_LOC_381/A INVX1_LOC_53/Y 0.07fF
C6960 INVX1_LOC_658/A INVX1_LOC_59/A 0.01fF
C6961 INVX1_LOC_79/A INVX1_LOC_109/Y 0.04fF
C6962 INVX1_LOC_118/Y INVX1_LOC_361/Y 0.00fF
C6963 INVX1_LOC_257/Y INVX1_LOC_32/Y 0.02fF
C6964 NAND2X1_LOC_790/B INVX1_LOC_95/A 0.02fF
C6965 INVX1_LOC_421/A NAND2X1_LOC_271/B 0.01fF
C6966 VDD NAND2X1_LOC_542/A 0.19fF
C6967 INVX1_LOC_395/A INVX1_LOC_117/Y 0.24fF
C6968 NAND2X1_LOC_842/a_36_24# NAND2X1_LOC_260/Y 0.00fF
C6969 INVX1_LOC_266/Y INVX1_LOC_59/Y 0.16fF
C6970 INVX1_LOC_300/A NAND2X1_LOC_318/A 0.07fF
C6971 INVX1_LOC_20/Y INVX1_LOC_115/A 0.03fF
C6972 NAND2X1_LOC_249/Y INVX1_LOC_63/Y 0.06fF
C6973 INVX1_LOC_300/A INVX1_LOC_268/Y -0.01fF
C6974 INVX1_LOC_162/Y INVX1_LOC_117/Y 0.01fF
C6975 INVX1_LOC_21/Y INVX1_LOC_84/A 0.19fF
C6976 INVX1_LOC_446/A INVX1_LOC_26/Y 0.07fF
C6977 INVX1_LOC_540/Y INVX1_LOC_47/Y 0.03fF
C6978 INVX1_LOC_266/Y INVX1_LOC_48/Y 0.01fF
C6979 INVX1_LOC_76/Y INVX1_LOC_440/A 0.01fF
C6980 NAND2X1_LOC_527/Y INVX1_LOC_45/Y -0.01fF
C6981 INVX1_LOC_537/A INVX1_LOC_495/A 0.05fF
C6982 INVX1_LOC_362/Y INVX1_LOC_117/Y 0.07fF
C6983 NAND2X1_LOC_525/Y NAND2X1_LOC_521/Y 0.13fF
C6984 INVX1_LOC_114/A INVX1_LOC_638/A 0.02fF
C6985 INVX1_LOC_20/Y INVX1_LOC_202/Y 0.03fF
C6986 INVX1_LOC_288/A INVX1_LOC_32/Y 0.07fF
C6987 VDD INVX1_LOC_376/Y 0.21fF
C6988 INVX1_LOC_666/A NAND2X1_LOC_615/B 0.02fF
C6989 INVX1_LOC_139/A INVX1_LOC_141/Y 0.06fF
C6990 INVX1_LOC_360/Y INVX1_LOC_686/A 0.71fF
C6991 NAND2X1_LOC_804/a_36_24# INVX1_LOC_116/Y 0.00fF
C6992 INVX1_LOC_85/Y NAND2X1_LOC_748/a_36_24# 0.00fF
C6993 INVX1_LOC_412/A NAND2X1_LOC_319/a_36_24# 0.00fF
C6994 INVX1_LOC_531/A INVX1_LOC_600/A 0.01fF
C6995 INVX1_LOC_12/Y INVX1_LOC_99/A 0.01fF
C6996 INVX1_LOC_89/Y INVX1_LOC_618/Y 0.03fF
C6997 INVX1_LOC_45/Y INVX1_LOC_93/A 0.01fF
C6998 INVX1_LOC_81/Y INVX1_LOC_184/A 0.01fF
C6999 INVX1_LOC_596/A INVX1_LOC_304/Y 0.02fF
C7000 INVX1_LOC_680/Y INVX1_LOC_683/A 0.00fF
C7001 INVX1_LOC_99/Y NAND2X1_LOC_496/Y 0.01fF
C7002 INVX1_LOC_384/A INVX1_LOC_32/Y 0.04fF
C7003 NAND2X1_LOC_377/a_36_24# INVX1_LOC_63/Y 0.00fF
C7004 NAND2X1_LOC_56/Y INVX1_LOC_35/Y 0.02fF
C7005 INVX1_LOC_173/A INVX1_LOC_47/Y 0.01fF
C7006 INVX1_LOC_158/A INVX1_LOC_242/Y 0.06fF
C7007 NAND2X1_LOC_160/a_36_24# INVX1_LOC_491/Y 0.00fF
C7008 INVX1_LOC_145/Y INVX1_LOC_7/Y 0.25fF
C7009 INVX1_LOC_586/A INVX1_LOC_94/Y 0.03fF
C7010 INVX1_LOC_490/Y INVX1_LOC_225/Y 0.13fF
C7011 INVX1_LOC_53/Y NAND2X1_LOC_720/A 0.07fF
C7012 VDD INVX1_LOC_40/A -0.00fF
C7013 INVX1_LOC_367/A INVX1_LOC_608/A 0.24fF
C7014 INVX1_LOC_115/A INVX1_LOC_197/Y 0.00fF
C7015 INVX1_LOC_685/A NAND2X1_LOC_864/a_36_24# 0.02fF
C7016 INVX1_LOC_266/A NAND2X1_LOC_388/A 0.03fF
C7017 INVX1_LOC_372/Y INVX1_LOC_355/Y 0.09fF
C7018 INVX1_LOC_677/Y INVX1_LOC_69/Y 0.14fF
C7019 INVX1_LOC_602/A INVX1_LOC_31/Y 0.02fF
C7020 INVX1_LOC_202/Y INVX1_LOC_300/A 0.07fF
C7021 INVX1_LOC_579/A NAND2X1_LOC_591/Y 0.08fF
C7022 NAND2X1_LOC_392/a_36_24# INVX1_LOC_9/Y 0.00fF
C7023 INVX1_LOC_202/Y INVX1_LOC_197/Y 0.07fF
C7024 NAND2X1_LOC_707/A INVX1_LOC_501/A 0.03fF
C7025 INVX1_LOC_547/Y NAND2X1_LOC_833/B 0.15fF
C7026 INVX1_LOC_588/Y INVX1_LOC_344/Y 0.23fF
C7027 INVX1_LOC_248/Y INVX1_LOC_440/Y 0.01fF
C7028 INVX1_LOC_451/A INVX1_LOC_453/Y 0.02fF
C7029 INVX1_LOC_374/A INVX1_LOC_26/Y 0.08fF
C7030 INVX1_LOC_20/Y INVX1_LOC_49/Y 0.25fF
C7031 NAND2X1_LOC_615/B NAND2X1_LOC_72/Y 0.01fF
C7032 INVX1_LOC_250/A INVX1_LOC_242/Y -0.01fF
C7033 INVX1_LOC_400/A NAND2X1_LOC_76/A 0.02fF
C7034 INVX1_LOC_58/Y INVX1_LOC_59/A 0.03fF
C7035 INVX1_LOC_35/Y NAND2X1_LOC_708/A 0.01fF
C7036 NAND2X1_LOC_706/B INVX1_LOC_99/Y 0.11fF
C7037 INVX1_LOC_448/A INVX1_LOC_32/Y 0.12fF
C7038 NAND2X1_LOC_567/a_36_24# INVX1_LOC_347/A 0.00fF
C7039 INVX1_LOC_17/Y INVX1_LOC_674/A 0.07fF
C7040 INVX1_LOC_685/Y INVX1_LOC_259/Y 0.16fF
C7041 INVX1_LOC_93/Y INVX1_LOC_281/Y 0.03fF
C7042 INVX1_LOC_367/A INVX1_LOC_58/Y 0.17fF
C7043 INVX1_LOC_76/Y INVX1_LOC_242/Y 0.07fF
C7044 INVX1_LOC_117/Y INVX1_LOC_189/Y 0.02fF
C7045 INVX1_LOC_402/A INVX1_LOC_6/Y 0.03fF
C7046 INVX1_LOC_254/Y INVX1_LOC_419/Y 0.01fF
C7047 INVX1_LOC_32/Y INVX1_LOC_145/Y 0.26fF
C7048 GATE_579 INVX1_LOC_244/Y 0.35fF
C7049 INVX1_LOC_548/A INVX1_LOC_117/Y 0.12fF
C7050 INVX1_LOC_373/A INVX1_LOC_588/A 0.00fF
C7051 INVX1_LOC_374/Y INVX1_LOC_252/Y 0.09fF
C7052 INVX1_LOC_7/Y INVX1_LOC_433/A 0.06fF
C7053 INVX1_LOC_63/Y INVX1_LOC_369/A 0.03fF
C7054 NAND2X1_LOC_796/a_36_24# INVX1_LOC_6/Y 0.00fF
C7055 INVX1_LOC_412/A NAND2X1_LOC_544/B 0.00fF
C7056 INVX1_LOC_53/Y NAND2X1_LOC_103/a_36_24# 0.00fF
C7057 INVX1_LOC_172/A INVX1_LOC_48/Y 0.00fF
C7058 INVX1_LOC_289/A NAND2X1_LOC_355/A 0.11fF
C7059 INVX1_LOC_20/A INVX1_LOC_26/Y 0.05fF
C7060 NAND2X1_LOC_697/Y NAND2X1_LOC_697/a_36_24# 0.02fF
C7061 INVX1_LOC_459/Y INVX1_LOC_74/Y 0.09fF
C7062 INVX1_LOC_76/Y INVX1_LOC_487/A 0.00fF
C7063 INVX1_LOC_516/A INVX1_LOC_58/Y 0.06fF
C7064 INVX1_LOC_439/Y NAND2X1_LOC_294/Y 0.03fF
C7065 INVX1_LOC_300/A INVX1_LOC_49/Y 0.07fF
C7066 INVX1_LOC_669/Y INVX1_LOC_58/Y 0.09fF
C7067 INVX1_LOC_117/Y INVX1_LOC_31/Y 2.43fF
C7068 INVX1_LOC_93/Y INVX1_LOC_608/A 0.03fF
C7069 INVX1_LOC_522/Y INVX1_LOC_475/Y 0.08fF
C7070 INVX1_LOC_547/A INVX1_LOC_62/Y 0.00fF
C7071 INVX1_LOC_285/A INVX1_LOC_79/A 0.00fF
C7072 INVX1_LOC_400/A INVX1_LOC_58/Y 0.20fF
C7073 INVX1_LOC_381/A INVX1_LOC_368/Y 0.03fF
C7074 INVX1_LOC_392/A INVX1_LOC_58/Y 0.00fF
C7075 INVX1_LOC_53/Y INVX1_LOC_100/Y 0.32fF
C7076 INVX1_LOC_20/Y INVX1_LOC_92/Y 0.01fF
C7077 INVX1_LOC_42/Y INVX1_LOC_9/Y 0.01fF
C7078 NAND2X1_LOC_615/B INVX1_LOC_351/Y 0.01fF
C7079 INVX1_LOC_376/Y INVX1_LOC_509/A 0.06fF
C7080 NAND2X1_LOC_521/Y INVX1_LOC_406/A 0.05fF
C7081 INVX1_LOC_478/Y INVX1_LOC_351/A 0.11fF
C7082 INVX1_LOC_435/A INVX1_LOC_245/A 0.01fF
C7083 INVX1_LOC_63/Y INVX1_LOC_603/A 0.00fF
C7084 INVX1_LOC_559/A INVX1_LOC_242/Y 0.03fF
C7085 INVX1_LOC_53/Y INVX1_LOC_74/Y 0.03fF
C7086 INVX1_LOC_93/Y INVX1_LOC_58/Y 0.34fF
C7087 NAND2X1_LOC_307/A INVX1_LOC_479/A 0.03fF
C7088 INVX1_LOC_50/Y INVX1_LOC_196/Y 0.02fF
C7089 NAND2X1_LOC_178/a_36_24# INVX1_LOC_6/Y 0.00fF
C7090 NAND2X1_LOC_387/Y INVX1_LOC_351/A 0.05fF
C7091 INVX1_LOC_478/Y INVX1_LOC_90/Y 0.02fF
C7092 INVX1_LOC_80/A NAND2X1_LOC_231/B 0.11fF
C7093 INVX1_LOC_593/Y NAND2X1_LOC_800/B 0.06fF
C7094 INVX1_LOC_300/A INVX1_LOC_92/Y 0.03fF
C7095 INVX1_LOC_551/Y INVX1_LOC_92/A 0.10fF
C7096 NAND2X1_LOC_387/Y INVX1_LOC_90/Y 0.01fF
C7097 NAND2X1_LOC_165/a_36_24# INVX1_LOC_91/A 0.00fF
C7098 INVX1_LOC_167/A NAND2X1_LOC_123/B 0.31fF
C7099 NAND2X1_LOC_190/A INVX1_LOC_62/Y 0.05fF
C7100 INVX1_LOC_193/A INVX1_LOC_41/Y 0.01fF
C7101 INVX1_LOC_419/Y INVX1_LOC_479/A 0.09fF
C7102 INVX1_LOC_460/Y INVX1_LOC_74/Y 0.21fF
C7103 INVX1_LOC_625/Y INVX1_LOC_252/Y 0.04fF
C7104 NAND2X1_LOC_274/B INVX1_LOC_420/A 0.28fF
C7105 INVX1_LOC_79/A INVX1_LOC_199/Y 0.06fF
C7106 INVX1_LOC_6/Y NAND2X1_LOC_625/a_36_24# 0.00fF
C7107 INVX1_LOC_491/A NAND2X1_LOC_221/a_36_24# 0.00fF
C7108 NAND2X1_LOC_376/B INVX1_LOC_41/Y 0.04fF
C7109 INVX1_LOC_124/A NAND2X1_LOC_137/a_36_24# 0.02fF
C7110 INVX1_LOC_376/A NAND2X1_LOC_118/a_36_24# 0.00fF
C7111 VDD INVX1_LOC_594/Y 0.21fF
C7112 INVX1_LOC_26/Y INVX1_LOC_81/A 0.02fF
C7113 NAND2X1_LOC_217/a_36_24# INVX1_LOC_442/A 0.01fF
C7114 INVX1_LOC_185/A INVX1_LOC_395/A 0.01fF
C7115 VDD INVX1_LOC_121/Y 0.21fF
C7116 INVX1_LOC_133/Y INVX1_LOC_570/A 0.00fF
C7117 INVX1_LOC_376/A INVX1_LOC_479/A 0.02fF
C7118 INVX1_LOC_291/Y INVX1_LOC_292/Y 0.01fF
C7119 INVX1_LOC_682/A INVX1_LOC_75/Y 0.03fF
C7120 INVX1_LOC_300/Y NAND2X1_LOC_451/B 0.01fF
C7121 NAND2X1_LOC_668/Y INVX1_LOC_658/Y 0.04fF
C7122 INVX1_LOC_20/Y INVX1_LOC_297/Y 0.03fF
C7123 NAND2X1_LOC_424/a_36_24# NAND2X1_LOC_832/A 0.00fF
C7124 VDD NAND2X1_LOC_142/Y 0.01fF
C7125 INVX1_LOC_502/A NAND2X1_LOC_528/Y 0.00fF
C7126 INVX1_LOC_376/A NAND2X1_LOC_468/a_36_24# 0.02fF
C7127 INVX1_LOC_91/A INVX1_LOC_90/Y 0.03fF
C7128 NAND2X1_LOC_475/A INVX1_LOC_271/A 0.12fF
C7129 NAND2X1_LOC_409/Y INVX1_LOC_41/Y 0.01fF
C7130 INVX1_LOC_206/Y NAND2X1_LOC_506/B 0.13fF
C7131 INVX1_LOC_206/Y INVX1_LOC_45/Y 1.39fF
C7132 INVX1_LOC_121/Y INVX1_LOC_510/Y 0.05fF
C7133 INVX1_LOC_195/A INVX1_LOC_366/A 0.03fF
C7134 INPUT_6 INVX1_LOC_45/A 0.05fF
C7135 INVX1_LOC_433/Y INVX1_LOC_406/Y 0.09fF
C7136 INVX1_LOC_435/Y INVX1_LOC_413/Y 0.00fF
C7137 NAND2X1_LOC_451/B INVX1_LOC_74/Y 0.00fF
C7138 NAND2X1_LOC_217/a_36_24# INVX1_LOC_116/Y 0.00fF
C7139 INVX1_LOC_48/Y INVX1_LOC_109/Y 0.01fF
C7140 INVX1_LOC_384/Y INVX1_LOC_445/A 0.03fF
C7141 INVX1_LOC_206/Y INVX1_LOC_348/A 0.05fF
C7142 INVX1_LOC_510/Y INVX1_LOC_253/A 0.01fF
C7143 INPUT_3 INVX1_LOC_206/Y 0.06fF
C7144 INVX1_LOC_224/Y INVX1_LOC_293/Y 0.02fF
C7145 VDD NAND2X1_LOC_603/Y -0.00fF
C7146 VDD INVX1_LOC_296/Y 0.21fF
C7147 INVX1_LOC_396/Y INVX1_LOC_45/Y 0.20fF
C7148 INVX1_LOC_446/Y INVX1_LOC_424/Y 0.04fF
C7149 INVX1_LOC_677/Y INVX1_LOC_586/A 0.07fF
C7150 NAND2X1_LOC_79/Y INVX1_LOC_180/A 0.09fF
C7151 VDD INVX1_LOC_332/Y 0.30fF
C7152 NAND2X1_LOC_770/A INVX1_LOC_598/A 0.09fF
C7153 INVX1_LOC_224/Y INVX1_LOC_160/A 0.02fF
C7154 INVX1_LOC_45/Y INVX1_LOC_686/A 0.07fF
C7155 NAND2X1_LOC_271/B INVX1_LOC_99/Y 0.01fF
C7156 INVX1_LOC_20/Y INVX1_LOC_76/Y 0.25fF
C7157 INVX1_LOC_587/A INVX1_LOC_55/Y 0.01fF
C7158 INVX1_LOC_602/A INVX1_LOC_51/Y 0.03fF
C7159 INVX1_LOC_206/Y NAND2X1_LOC_69/Y 0.01fF
C7160 INVX1_LOC_118/Y NAND2X1_LOC_692/Y 0.01fF
C7161 INVX1_LOC_442/A NAND2X1_LOC_325/B 0.33fF
C7162 NAND2X1_LOC_99/a_36_24# INVX1_LOC_96/A 0.02fF
C7163 INVX1_LOC_395/A INVX1_LOC_251/Y 0.12fF
C7164 INVX1_LOC_395/A INVX1_LOC_178/A 0.22fF
C7165 INVX1_LOC_581/A INVX1_LOC_142/A 0.03fF
C7166 INVX1_LOC_628/A INVX1_LOC_459/Y 0.07fF
C7167 INVX1_LOC_629/A INVX1_LOC_460/Y 0.10fF
C7168 INVX1_LOC_21/Y INVX1_LOC_174/Y 0.01fF
C7169 INVX1_LOC_242/Y INVX1_LOC_192/A 0.01fF
C7170 INVX1_LOC_53/Y INVX1_LOC_566/A 0.07fF
C7171 NAND2X1_LOC_331/A INVX1_LOC_514/A 0.05fF
C7172 VDD INVX1_LOC_477/Y 0.26fF
C7173 NAND2X1_LOC_790/B INVX1_LOC_63/Y 0.09fF
C7174 INVX1_LOC_33/Y INVX1_LOC_35/Y 0.21fF
C7175 INVX1_LOC_406/Y INVX1_LOC_232/Y 0.00fF
C7176 INVX1_LOC_21/Y NAND2X1_LOC_79/B 0.01fF
C7177 INVX1_LOC_616/A INVX1_LOC_145/Y 0.01fF
C7178 INVX1_LOC_676/Y INVX1_LOC_495/A 0.44fF
C7179 INVX1_LOC_602/A NAND2X1_LOC_805/a_36_24# 0.00fF
C7180 INVX1_LOC_300/A INVX1_LOC_76/Y 0.10fF
C7181 VDD INVX1_LOC_139/Y 0.36fF
C7182 INVX1_LOC_449/A NAND2X1_LOC_541/B 0.32fF
C7183 NAND2X1_LOC_164/a_36_24# INVX1_LOC_273/A 0.02fF
C7184 INVX1_LOC_169/A INVX1_LOC_99/Y 0.01fF
C7185 INVX1_LOC_76/Y INVX1_LOC_197/Y 0.03fF
C7186 NAND2X1_LOC_505/Y INVX1_LOC_117/Y 0.03fF
C7187 INVX1_LOC_562/A INVX1_LOC_47/Y 0.00fF
C7188 INVX1_LOC_133/A NAND2X1_LOC_288/a_36_24# 0.00fF
C7189 INVX1_LOC_80/A NAND2X1_LOC_768/A 0.03fF
C7190 INVX1_LOC_20/Y INVX1_LOC_559/A 0.01fF
C7191 NAND2X1_LOC_317/B INVX1_LOC_47/Y 0.02fF
C7192 INVX1_LOC_553/A INVX1_LOC_49/Y 0.01fF
C7193 NAND2X1_LOC_493/B INVX1_LOC_194/Y 0.01fF
C7194 INVX1_LOC_362/Y INVX1_LOC_608/A 0.02fF
C7195 NAND2X1_LOC_299/Y NAND2X1_LOC_123/A 0.01fF
C7196 INVX1_LOC_29/Y INVX1_LOC_69/A 0.05fF
C7197 INVX1_LOC_117/Y INVX1_LOC_51/Y 0.90fF
C7198 INVX1_LOC_84/A INVX1_LOC_481/Y 0.01fF
C7199 INVX1_LOC_459/Y INVX1_LOC_469/Y 0.11fF
C7200 INVX1_LOC_99/Y INVX1_LOC_633/Y 0.03fF
C7201 INVX1_LOC_583/A NAND2X1_LOC_679/B 0.01fF
C7202 NAND2X1_LOC_16/Y INVX1_LOC_6/Y 0.16fF
C7203 NAND2X1_LOC_179/Y INVX1_LOC_519/A 0.16fF
C7204 INVX1_LOC_115/A NAND2X1_LOC_298/a_36_24# 0.00fF
C7205 INVX1_LOC_395/A INVX1_LOC_58/Y 0.36fF
C7206 INVX1_LOC_379/A INVX1_LOC_489/Y 0.09fF
C7207 INVX1_LOC_609/A INVX1_LOC_581/A 0.09fF
C7208 INVX1_LOC_602/A INVX1_LOC_40/Y 0.12fF
C7209 INVX1_LOC_551/Y INPUT_1 0.03fF
C7210 INVX1_LOC_162/Y INVX1_LOC_58/Y 0.01fF
C7211 NAND2X1_LOC_325/B INVX1_LOC_116/Y 0.36fF
C7212 NAND2X1_LOC_331/A INVX1_LOC_534/Y 0.03fF
C7213 INVX1_LOC_11/Y INVX1_LOC_80/A 0.26fF
C7214 NAND2X1_LOC_331/A NAND2X1_LOC_800/B 0.14fF
C7215 NAND2X1_LOC_835/a_36_24# INVX1_LOC_59/A 0.00fF
C7216 INVX1_LOC_416/A INVX1_LOC_12/Y 0.01fF
C7217 INVX1_LOC_45/Y NAND2X1_LOC_334/A 0.03fF
C7218 INVX1_LOC_362/Y INVX1_LOC_58/Y 0.01fF
C7219 NAND2X1_LOC_317/B INVX1_LOC_119/Y 0.21fF
C7220 INVX1_LOC_47/Y INVX1_LOC_169/A 0.03fF
C7221 NAND2X1_LOC_210/A INVX1_LOC_145/Y 0.02fF
C7222 INVX1_LOC_6/Y NAND2X1_LOC_783/a_36_24# 0.00fF
C7223 NAND2X1_LOC_738/a_36_24# INVX1_LOC_575/Y 0.00fF
C7224 INVX1_LOC_375/A NAND2X1_LOC_657/a_36_24# 0.00fF
C7225 NAND2X1_LOC_557/B INVX1_LOC_169/A 0.00fF
C7226 INVX1_LOC_424/Y INVX1_LOC_433/A 0.01fF
C7227 INVX1_LOC_586/A INVX1_LOC_357/Y 0.01fF
C7228 INVX1_LOC_53/Y INVX1_LOC_469/Y 0.05fF
C7229 INVX1_LOC_628/A INVX1_LOC_460/Y 0.17fF
C7230 INVX1_LOC_367/A NAND2X1_LOC_496/a_36_24# 0.00fF
C7231 INVX1_LOC_678/Y INVX1_LOC_58/Y 0.01fF
C7232 NAND2X1_LOC_303/a_36_24# INVX1_LOC_353/A 0.01fF
C7233 NAND2X1_LOC_152/Y INVX1_LOC_569/Y 0.01fF
C7234 INVX1_LOC_614/A INVX1_LOC_477/Y 0.05fF
C7235 NAND2X1_LOC_331/A INVX1_LOC_62/Y 0.08fF
C7236 INPUT_0 INVX1_LOC_75/Y 0.14fF
C7237 INVX1_LOC_47/Y INVX1_LOC_633/Y 0.46fF
C7238 NAND2X1_LOC_142/a_36_24# NAND2X1_LOC_248/B 0.00fF
C7239 INVX1_LOC_567/Y INVX1_LOC_46/Y 0.01fF
C7240 INVX1_LOC_459/Y INVX1_LOC_79/A 0.02fF
C7241 INVX1_LOC_69/Y INVX1_LOC_635/A 0.00fF
C7242 INVX1_LOC_566/A NAND2X1_LOC_406/B 0.04fF
C7243 INVX1_LOC_349/A INVX1_LOC_159/Y 0.02fF
C7244 INVX1_LOC_372/Y INVX1_LOC_376/A 0.25fF
C7245 INVX1_LOC_21/Y NAND2X1_LOC_532/Y 0.02fF
C7246 NAND2X1_LOC_707/A INVX1_LOC_461/Y 0.14fF
C7247 INVX1_LOC_49/Y INVX1_LOC_375/Y 0.05fF
C7248 INVX1_LOC_69/Y NAND2X1_LOC_237/Y 0.03fF
C7249 INVX1_LOC_548/A INVX1_LOC_608/A 0.00fF
C7250 INVX1_LOC_32/Y INVX1_LOC_503/Y 0.00fF
C7251 INVX1_LOC_31/Y INVX1_LOC_178/A 0.04fF
C7252 INVX1_LOC_81/Y INVX1_LOC_86/Y 0.03fF
C7253 INVX1_LOC_417/Y INVX1_LOC_199/Y 0.07fF
C7254 INVX1_LOC_188/Y INVX1_LOC_338/Y 0.07fF
C7255 NAND2X1_LOC_326/a_36_24# INVX1_LOC_376/A 0.00fF
C7256 INVX1_LOC_639/Y INVX1_LOC_639/A 0.15fF
C7257 INVX1_LOC_459/Y INVX1_LOC_460/A 0.01fF
C7258 INVX1_LOC_21/Y NAND2X1_LOC_376/B 0.03fF
C7259 NAND2X1_LOC_169/A INVX1_LOC_154/A 0.00fF
C7260 NAND2X1_LOC_104/a_36_24# INVX1_LOC_178/A 0.00fF
C7261 INVX1_LOC_84/A INVX1_LOC_26/Y 1.31fF
C7262 INVX1_LOC_169/A NAND2X1_LOC_66/Y 0.01fF
C7263 INVX1_LOC_469/Y INVX1_LOC_460/Y 0.03fF
C7264 INVX1_LOC_591/Y INVX1_LOC_26/Y 0.05fF
C7265 INVX1_LOC_183/A INVX1_LOC_530/A 0.02fF
C7266 INVX1_LOC_137/Y INVX1_LOC_66/A 0.07fF
C7267 NAND2X1_LOC_531/Y INVX1_LOC_35/Y 0.03fF
C7268 INVX1_LOC_199/Y INVX1_LOC_59/Y 0.29fF
C7269 NAND2X1_LOC_184/Y INVX1_LOC_362/A 0.34fF
C7270 INVX1_LOC_431/A INVX1_LOC_6/Y 0.24fF
C7271 INVX1_LOC_58/Y INVX1_LOC_189/Y 0.00fF
C7272 INVX1_LOC_119/Y INVX1_LOC_633/Y 0.07fF
C7273 INVX1_LOC_47/Y NAND2X1_LOC_308/a_36_24# 0.00fF
C7274 INVX1_LOC_134/Y INVX1_LOC_114/A 4.99fF
C7275 INPUT_0 NAND2X1_LOC_271/A 0.07fF
C7276 INVX1_LOC_556/Y INVX1_LOC_63/Y 0.03fF
C7277 NAND2X1_LOC_467/A NAND2X1_LOC_691/A 0.01fF
C7278 INVX1_LOC_496/A NAND2X1_LOC_220/a_36_24# 0.00fF
C7279 INVX1_LOC_53/Y INVX1_LOC_79/A 6.43fF
C7280 INVX1_LOC_105/A NAND2X1_LOC_542/A 1.53fF
C7281 INVX1_LOC_199/Y INVX1_LOC_48/Y 0.44fF
C7282 INVX1_LOC_575/A INVX1_LOC_9/Y 0.02fF
C7283 INVX1_LOC_47/Y NAND2X1_LOC_119/a_36_24# 0.01fF
C7284 INVX1_LOC_447/Y NAND2X1_LOC_274/B 0.00fF
C7285 INVX1_LOC_6/Y INVX1_LOC_18/Y 0.05fF
C7286 NAND2X1_LOC_716/a_36_24# INVX1_LOC_353/A 0.01fF
C7287 NAND2X1_LOC_448/B INVX1_LOC_187/Y 0.01fF
C7288 INVX1_LOC_59/Y INVX1_LOC_272/A 0.01fF
C7289 INVX1_LOC_105/A INVX1_LOC_376/Y 0.06fF
C7290 INVX1_LOC_451/A INVX1_LOC_422/A 0.05fF
C7291 INVX1_LOC_506/A INVX1_LOC_63/Y 0.01fF
C7292 NAND2X1_LOC_274/B NAND2X1_LOC_602/A 0.01fF
C7293 NAND2X1_LOC_121/Y INVX1_LOC_50/Y 0.06fF
C7294 INVX1_LOC_31/Y INVX1_LOC_58/Y 0.51fF
C7295 INVX1_LOC_11/Y NAND2X1_LOC_433/Y 0.48fF
C7296 INVX1_LOC_7/Y INVX1_LOC_487/A 0.03fF
C7297 INVX1_LOC_498/A INVX1_LOC_498/Y 0.19fF
C7298 INVX1_LOC_665/A INVX1_LOC_367/Y 0.11fF
C7299 NAND2X1_LOC_308/a_36_24# INVX1_LOC_119/Y 0.00fF
C7300 INVX1_LOC_292/Y NAND2X1_LOC_759/Y 0.02fF
C7301 INVX1_LOC_632/Y INVX1_LOC_263/Y 0.01fF
C7302 INVX1_LOC_54/Y NAND2X1_LOC_274/B 0.03fF
C7303 INVX1_LOC_213/Y INVX1_LOC_100/Y 0.03fF
C7304 INVX1_LOC_80/A NAND2X1_LOC_244/a_36_24# 0.00fF
C7305 INVX1_LOC_17/Y NAND2X1_LOC_528/Y 0.03fF
C7306 INVX1_LOC_93/Y INVX1_LOC_245/A 0.06fF
C7307 INVX1_LOC_460/Y INVX1_LOC_79/A 0.02fF
C7308 INVX1_LOC_32/Y INVX1_LOC_242/Y 0.07fF
C7309 INVX1_LOC_608/Y INVX1_LOC_479/A 0.01fF
C7310 INVX1_LOC_407/Y INVX1_LOC_62/Y 1.09fF
C7311 INVX1_LOC_17/Y INVX1_LOC_479/A 0.22fF
C7312 INVX1_LOC_270/A INVX1_LOC_92/A 0.05fF
C7313 NAND2X1_LOC_119/a_36_24# INVX1_LOC_119/Y 0.00fF
C7314 INVX1_LOC_413/A INVX1_LOC_41/Y 0.01fF
C7315 INVX1_LOC_460/Y INVX1_LOC_460/A 0.01fF
C7316 INVX1_LOC_518/Y NAND2X1_LOC_659/a_36_24# 0.00fF
C7317 INVX1_LOC_179/A INVX1_LOC_351/Y 0.03fF
C7318 INVX1_LOC_380/A NAND2X1_LOC_475/A 0.01fF
C7319 INVX1_LOC_675/A INVX1_LOC_245/A 0.07fF
C7320 NAND2X1_LOC_186/a_36_24# INVX1_LOC_62/Y 0.00fF
C7321 INVX1_LOC_35/Y INVX1_LOC_443/A 0.17fF
C7322 INVX1_LOC_390/A INVX1_LOC_245/A 0.01fF
C7323 NAND2X1_LOC_294/Y INVX1_LOC_325/A 0.11fF
C7324 NAND2X1_LOC_698/Y INVX1_LOC_100/Y 0.01fF
C7325 NAND2X1_LOC_334/B INVX1_LOC_245/A 0.08fF
C7326 NAND2X1_LOC_816/a_36_24# INVX1_LOC_655/A 0.00fF
C7327 NAND2X1_LOC_307/B INVX1_LOC_479/A 0.05fF
C7328 INVX1_LOC_662/A INVX1_LOC_100/Y 0.20fF
C7329 INVX1_LOC_647/Y INVX1_LOC_66/A 0.03fF
C7330 INVX1_LOC_520/Y INVX1_LOC_241/A 0.25fF
C7331 NAND2X1_LOC_192/A INVX1_LOC_653/Y 0.02fF
C7332 NAND2X1_LOC_724/a_36_24# NAND2X1_LOC_513/Y 0.00fF
C7333 INVX1_LOC_551/A INVX1_LOC_211/A 0.03fF
C7334 NAND2X1_LOC_582/a_36_24# INVX1_LOC_677/Y 0.00fF
C7335 INVX1_LOC_293/A INVX1_LOC_282/Y 0.00fF
C7336 INVX1_LOC_373/Y INVX1_LOC_41/Y 0.01fF
C7337 INVX1_LOC_62/Y NAND2X1_LOC_833/B 0.02fF
C7338 INVX1_LOC_46/Y INVX1_LOC_92/A 8.32fF
C7339 NAND2X1_LOC_526/Y VDD 0.30fF
C7340 INVX1_LOC_20/Y NAND2X1_LOC_770/A 0.16fF
C7341 INVX1_LOC_41/Y NAND2X1_LOC_691/A 0.02fF
C7342 NAND2X1_LOC_781/B INVX1_LOC_522/Y 0.04fF
C7343 NAND2X1_LOC_457/A INVX1_LOC_364/Y 0.15fF
C7344 VDD INVX1_LOC_168/A -0.00fF
C7345 INVX1_LOC_75/Y INVX1_LOC_211/A 0.00fF
C7346 INVX1_LOC_397/A INVX1_LOC_45/Y 0.06fF
C7347 INVX1_LOC_206/Y NAND2X1_LOC_756/Y 0.09fF
C7348 INVX1_LOC_94/A NAND2X1_LOC_506/B 0.01fF
C7349 INVX1_LOC_12/Y INVX1_LOC_388/Y 0.07fF
C7350 INVX1_LOC_206/Y INVX1_LOC_293/Y 0.09fF
C7351 INVX1_LOC_405/A NAND2X1_LOC_275/Y 0.01fF
C7352 INVX1_LOC_265/Y INVX1_LOC_495/A 0.00fF
C7353 INVX1_LOC_45/Y INVX1_LOC_94/A 0.00fF
C7354 INVX1_LOC_257/Y NAND2X1_LOC_299/Y 0.01fF
C7355 NAND2X1_LOC_239/a_36_24# INVX1_LOC_80/A 0.01fF
C7356 NAND2X1_LOC_457/A INVX1_LOC_134/Y 0.01fF
C7357 NAND2X1_LOC_231/B INVX1_LOC_91/Y 0.07fF
C7358 NAND2X1_LOC_543/B NAND2X1_LOC_775/B 0.03fF
C7359 NAND2X1_LOC_836/B INVX1_LOC_41/A 0.05fF
C7360 INVX1_LOC_20/Y INVX1_LOC_276/A 0.04fF
C7361 NAND2X1_LOC_140/a_36_24# NAND2X1_LOC_140/B 0.00fF
C7362 NAND2X1_LOC_756/Y INVX1_LOC_396/Y 0.07fF
C7363 INVX1_LOC_177/Y INVX1_LOC_21/Y 0.01fF
C7364 INVX1_LOC_250/Y NAND2X1_LOC_303/a_36_24# 0.00fF
C7365 VDD NAND2X1_LOC_635/B 0.26fF
C7366 INVX1_LOC_560/Y INVX1_LOC_603/A 0.01fF
C7367 VDD INVX1_LOC_640/Y 0.21fF
C7368 INVX1_LOC_586/A INVX1_LOC_635/A 0.33fF
C7369 INVX1_LOC_301/A INVX1_LOC_32/Y 0.03fF
C7370 INVX1_LOC_516/Y NAND2X1_LOC_656/a_36_24# 0.00fF
C7371 VDD INVX1_LOC_536/Y 0.21fF
C7372 INVX1_LOC_206/Y NAND2X1_LOC_673/B 0.08fF
C7373 NAND2X1_LOC_97/A NAND2X1_LOC_97/B 0.00fF
C7374 INVX1_LOC_606/Y INVX1_LOC_35/Y 0.02fF
C7375 INVX1_LOC_586/A NAND2X1_LOC_237/Y 0.00fF
C7376 VDD NAND2X1_LOC_619/Y 0.00fF
C7377 INVX1_LOC_193/Y INVX1_LOC_159/Y 0.03fF
C7378 NAND2X1_LOC_45/Y INVX1_LOC_166/A 0.08fF
C7379 INVX1_LOC_617/Y INVX1_LOC_519/A 0.02fF
C7380 INVX1_LOC_119/A INVX1_LOC_519/A 0.00fF
C7381 NAND2X1_LOC_475/A INVX1_LOC_317/A 0.00fF
C7382 INVX1_LOC_84/A INVX1_LOC_369/A 0.03fF
C7383 INVX1_LOC_586/A INVX1_LOC_230/A 0.07fF
C7384 INVX1_LOC_510/Y INVX1_LOC_251/A 0.01fF
C7385 NAND2X1_LOC_38/a_36_24# INVX1_LOC_169/A 0.00fF
C7386 INVX1_LOC_142/Y NAND2X1_LOC_156/Y 0.20fF
C7387 INVX1_LOC_80/A INVX1_LOC_131/A 0.21fF
C7388 VDD INVX1_LOC_654/Y 0.21fF
C7389 INVX1_LOC_176/Y INVX1_LOC_323/Y 0.98fF
C7390 INPUT_7 INVX1_LOC_29/Y 0.03fF
C7391 INVX1_LOC_20/Y INVX1_LOC_228/A 0.02fF
C7392 INVX1_LOC_418/A INPUT_1 0.03fF
C7393 INVX1_LOC_53/Y INVX1_LOC_632/A 0.07fF
C7394 INVX1_LOC_166/A NAND2X1_LOC_498/Y 0.05fF
C7395 INVX1_LOC_366/A GATE_222 0.03fF
C7396 INVX1_LOC_166/A INVX1_LOC_570/A 0.03fF
C7397 INVX1_LOC_558/A INPUT_1 0.01fF
C7398 INVX1_LOC_11/Y NAND2X1_LOC_704/B 0.04fF
C7399 INVX1_LOC_374/A INVX1_LOC_506/A 0.01fF
C7400 INVX1_LOC_292/A INVX1_LOC_69/Y 0.21fF
C7401 INVX1_LOC_417/Y INVX1_LOC_53/Y 0.03fF
C7402 INVX1_LOC_54/Y INVX1_LOC_38/A 0.15fF
C7403 INVX1_LOC_17/Y INVX1_LOC_372/Y 0.03fF
C7404 NAND2X1_LOC_548/B NAND2X1_LOC_529/Y 0.06fF
C7405 INVX1_LOC_577/Y INVX1_LOC_156/A 0.01fF
C7406 INPUT_0 INVX1_LOC_513/Y 0.94fF
C7407 INPUT_2 INVX1_LOC_83/Y 0.03fF
C7408 INVX1_LOC_312/Y INVX1_LOC_230/A 0.02fF
C7409 NAND2X1_LOC_513/Y INVX1_LOC_199/Y 0.07fF
C7410 NAND2X1_LOC_184/Y INVX1_LOC_384/A 0.17fF
C7411 INVX1_LOC_250/Y NAND2X1_LOC_716/a_36_24# 0.00fF
C7412 INVX1_LOC_504/A INVX1_LOC_188/Y 0.07fF
C7413 INVX1_LOC_53/Y INVX1_LOC_59/Y 0.03fF
C7414 INVX1_LOC_20/Y INVX1_LOC_345/Y 0.03fF
C7415 INVX1_LOC_584/Y INVX1_LOC_493/Y 0.21fF
C7416 NAND2X1_LOC_534/Y NAND2X1_LOC_274/B 0.01fF
C7417 NAND2X1_LOC_13/Y INVX1_LOC_117/Y 0.10fF
C7418 INVX1_LOC_62/Y INVX1_LOC_638/A 0.12fF
C7419 INVX1_LOC_400/Y INVX1_LOC_411/Y 0.03fF
C7420 INVX1_LOC_17/Y INVX1_LOC_12/Y 0.20fF
C7421 INVX1_LOC_51/Y INVX1_LOC_157/A 0.04fF
C7422 INVX1_LOC_106/A INVX1_LOC_99/Y 0.01fF
C7423 INVX1_LOC_20/Y INVX1_LOC_32/Y 0.19fF
C7424 INVX1_LOC_175/Y INVX1_LOC_32/Y 0.05fF
C7425 INVX1_LOC_578/A INVX1_LOC_682/A 0.03fF
C7426 INVX1_LOC_395/A INVX1_LOC_245/A 0.03fF
C7427 NAND2X1_LOC_467/A INVX1_LOC_496/Y 0.00fF
C7428 INVX1_LOC_53/Y INVX1_LOC_48/Y 1.45fF
C7429 INVX1_LOC_51/Y INVX1_LOC_58/Y 0.07fF
C7430 VDD INVX1_LOC_11/A -0.00fF
C7431 INVX1_LOC_80/A INVX1_LOC_374/Y 0.01fF
C7432 INVX1_LOC_432/Y INVX1_LOC_11/Y 0.03fF
C7433 INVX1_LOC_607/Y INVX1_LOC_492/A 0.06fF
C7434 INVX1_LOC_259/A INVX1_LOC_353/A 0.07fF
C7435 INVX1_LOC_588/Y INVX1_LOC_99/Y 4.30fF
C7436 NAND2X1_LOC_387/Y NAND2X1_LOC_318/B 0.30fF
C7437 INVX1_LOC_35/Y INVX1_LOC_371/A 0.01fF
C7438 INVX1_LOC_466/A INVX1_LOC_537/A 0.03fF
C7439 INVX1_LOC_174/Y INVX1_LOC_26/Y 0.00fF
C7440 NAND2X1_LOC_383/Y NAND2X1_LOC_558/B 0.04fF
C7441 INVX1_LOC_400/Y INVX1_LOC_41/Y 0.03fF
C7442 NAND2X1_LOC_184/Y INVX1_LOC_145/Y 0.10fF
C7443 INVX1_LOC_300/A INVX1_LOC_32/Y 0.99fF
C7444 INVX1_LOC_211/Y INPUT_1 0.03fF
C7445 NAND2X1_LOC_540/a_36_24# INVX1_LOC_392/A 0.00fF
C7446 INVX1_LOC_303/Y INVX1_LOC_665/Y 0.00fF
C7447 INVX1_LOC_508/Y NAND2X1_LOC_846/B 0.12fF
C7448 VDD INVX1_LOC_462/Y 0.40fF
C7449 INVX1_LOC_326/Y NAND2X1_LOC_397/Y 0.01fF
C7450 INVX1_LOC_32/Y INVX1_LOC_197/Y 0.06fF
C7451 INVX1_LOC_276/A INVX1_LOC_655/A 0.04fF
C7452 INVX1_LOC_547/A NAND2X1_LOC_833/B 0.20fF
C7453 NAND2X1_LOC_592/B INVX1_LOC_479/A 0.01fF
C7454 NAND2X1_LOC_325/B INVX1_LOC_69/Y 0.12fF
C7455 INVX1_LOC_54/Y INVX1_LOC_159/Y 0.08fF
C7456 INVX1_LOC_446/Y INVX1_LOC_75/Y 0.02fF
C7457 INVX1_LOC_17/Y INVX1_LOC_391/A 0.01fF
C7458 NAND2X1_LOC_185/a_36_24# INVX1_LOC_62/Y 0.00fF
C7459 INVX1_LOC_612/Y INVX1_LOC_550/A 0.01fF
C7460 INVX1_LOC_54/Y NAND2X1_LOC_782/A 0.05fF
C7461 INVX1_LOC_15/Y INVX1_LOC_633/Y 0.01fF
C7462 INVX1_LOC_167/A INVX1_LOC_50/Y 0.00fF
C7463 INVX1_LOC_582/A NAND2X1_LOC_679/B 0.01fF
C7464 NAND2X1_LOC_596/Y INVX1_LOC_462/Y 0.00fF
C7465 INVX1_LOC_84/A NAND2X1_LOC_626/Y 0.00fF
C7466 INVX1_LOC_418/Y INVX1_LOC_257/A 0.01fF
C7467 INVX1_LOC_6/Y GATE_222 0.01fF
C7468 INVX1_LOC_17/Y INVX1_LOC_170/A 0.01fF
C7469 INPUT_1 INVX1_LOC_46/Y 0.13fF
C7470 INVX1_LOC_551/A INVX1_LOC_145/Y 0.00fF
C7471 INVX1_LOC_384/A INVX1_LOC_75/Y 0.01fF
C7472 INVX1_LOC_588/Y INVX1_LOC_47/Y 0.66fF
C7473 NAND2X1_LOC_274/B INVX1_LOC_371/Y 0.00fF
C7474 INVX1_LOC_130/Y INVX1_LOC_242/Y 0.05fF
C7475 INVX1_LOC_500/Y INVX1_LOC_58/Y 0.15fF
C7476 INVX1_LOC_58/Y INVX1_LOC_40/Y 0.00fF
C7477 NAND2X1_LOC_274/Y INVX1_LOC_48/Y 0.00fF
C7478 INVX1_LOC_446/Y NAND2X1_LOC_271/A 0.04fF
C7479 INVX1_LOC_166/A NAND2X1_LOC_306/a_36_24# 0.00fF
C7480 NAND2X1_LOC_708/A INVX1_LOC_507/Y 0.02fF
C7481 INVX1_LOC_166/A INVX1_LOC_47/Y 0.11fF
C7482 INVX1_LOC_498/A NAND2X1_LOC_427/a_36_24# 0.01fF
C7483 INVX1_LOC_267/A NAND2X1_LOC_753/Y 0.01fF
C7484 INVX1_LOC_254/A INVX1_LOC_58/Y 0.00fF
C7485 INVX1_LOC_80/A NAND2X1_LOC_843/B 0.11fF
C7486 INPUT_5 INVX1_LOC_18/A 0.01fF
C7487 NAND2X1_LOC_768/A NAND2X1_LOC_843/B 0.01fF
C7488 INVX1_LOC_117/Y INVX1_LOC_196/Y 0.05fF
C7489 INVX1_LOC_358/Y NAND2X1_LOC_691/A 0.01fF
C7490 NAND2X1_LOC_123/B INVX1_LOC_115/A 0.00fF
C7491 INVX1_LOC_81/Y INVX1_LOC_81/A 0.01fF
C7492 INVX1_LOC_100/Y INVX1_LOC_679/A 0.00fF
C7493 INVX1_LOC_652/A INVX1_LOC_509/A 0.05fF
C7494 INVX1_LOC_531/Y INVX1_LOC_99/Y 0.06fF
C7495 INVX1_LOC_502/A INVX1_LOC_159/A 0.10fF
C7496 INVX1_LOC_537/A INVX1_LOC_41/Y 0.07fF
C7497 INVX1_LOC_632/A NAND2X1_LOC_451/B 0.07fF
C7498 INPUT_5 INPUT_4 1.66fF
C7499 NAND2X1_LOC_755/B NAND2X1_LOC_827/a_36_24# 0.00fF
C7500 INVX1_LOC_156/A INVX1_LOC_26/Y 0.15fF
C7501 INVX1_LOC_588/Y INVX1_LOC_119/Y 0.09fF
C7502 INVX1_LOC_80/A INVX1_LOC_91/Y 0.82fF
C7503 NAND2X1_LOC_318/A INVX1_LOC_92/A 0.01fF
C7504 INVX1_LOC_80/A INVX1_LOC_625/Y 2.73fF
C7505 INVX1_LOC_145/Y INVX1_LOC_75/Y 0.10fF
C7506 INVX1_LOC_35/Y NAND2X1_LOC_488/Y 0.01fF
C7507 INVX1_LOC_31/Y INVX1_LOC_245/A 11.41fF
C7508 INVX1_LOC_488/Y INVX1_LOC_489/Y 0.06fF
C7509 INVX1_LOC_166/A INVX1_LOC_119/Y 3.19fF
C7510 INVX1_LOC_62/Y INVX1_LOC_665/Y 0.03fF
C7511 INVX1_LOC_35/Y INVX1_LOC_645/Y 0.00fF
C7512 INVX1_LOC_479/A INVX1_LOC_108/Y 0.01fF
C7513 INVX1_LOC_89/Y NAND2X1_LOC_274/B 0.05fF
C7514 INVX1_LOC_421/A INVX1_LOC_41/Y 0.15fF
C7515 NAND2X1_LOC_815/a_36_24# INVX1_LOC_655/A 0.01fF
C7516 NAND2X1_LOC_410/Y INVX1_LOC_50/Y 0.00fF
C7517 INVX1_LOC_41/Y INVX1_LOC_496/Y 0.05fF
C7518 INVX1_LOC_589/Y INVX1_LOC_531/Y 0.03fF
C7519 NAND2X1_LOC_528/Y INVX1_LOC_230/Y 0.19fF
C7520 NAND2X1_LOC_111/Y INVX1_LOC_119/Y 0.02fF
C7521 NAND2X1_LOC_286/A INVX1_LOC_655/A 0.05fF
C7522 INVX1_LOC_54/Y INVX1_LOC_39/Y 0.01fF
C7523 INVX1_LOC_561/A INVX1_LOC_74/Y 0.01fF
C7524 INVX1_LOC_47/Y INVX1_LOC_531/Y 1.70fF
C7525 INVX1_LOC_145/Y NAND2X1_LOC_271/A 0.04fF
C7526 INVX1_LOC_609/A INVX1_LOC_613/A 0.33fF
C7527 NAND2X1_LOC_557/B INVX1_LOC_531/Y 0.28fF
C7528 NAND2X1_LOC_231/B NAND2X1_LOC_333/B 0.49fF
C7529 NAND2X1_LOC_448/B INVX1_LOC_354/A 0.01fF
C7530 INVX1_LOC_49/Y NAND2X1_LOC_123/B 0.03fF
C7531 INVX1_LOC_47/Y NAND2X1_LOC_433/a_36_24# 0.01fF
C7532 INVX1_LOC_100/Y NAND2X1_LOC_545/A 0.00fF
C7533 INPUT_0 INVX1_LOC_224/Y 0.10fF
C7534 INVX1_LOC_239/Y INVX1_LOC_131/Y 0.07fF
C7535 INVX1_LOC_118/Y INVX1_LOC_215/Y 0.01fF
C7536 NAND2X1_LOC_545/A INVX1_LOC_74/Y 0.33fF
C7537 INVX1_LOC_405/A INVX1_LOC_235/Y 0.01fF
C7538 INPUT_0 INVX1_LOC_578/A 0.07fF
C7539 INVX1_LOC_317/Y NAND2X1_LOC_475/A 0.02fF
C7540 INVX1_LOC_100/Y INVX1_LOC_666/Y 0.07fF
C7541 NAND2X1_LOC_271/B NAND2X1_LOC_520/B 0.04fF
C7542 INVX1_LOC_49/Y INVX1_LOC_92/A 0.07fF
C7543 INVX1_LOC_182/A INVX1_LOC_395/A 0.03fF
C7544 INVX1_LOC_388/A NAND2X1_LOC_489/a_36_24# 0.02fF
C7545 INVX1_LOC_344/A INVX1_LOC_638/A 0.05fF
C7546 INVX1_LOC_73/Y INVX1_LOC_7/Y 0.05fF
C7547 INVX1_LOC_425/A INVX1_LOC_412/A 0.35fF
C7548 INVX1_LOC_301/A INVX1_LOC_130/Y 0.02fF
C7549 INVX1_LOC_270/Y INVX1_LOC_92/Y 0.02fF
C7550 INVX1_LOC_603/Y NAND2X1_LOC_76/B 0.01fF
C7551 NAND2X1_LOC_638/A INVX1_LOC_562/A 0.03fF
C7552 NAND2X1_LOC_229/a_36_24# INVX1_LOC_586/A 0.00fF
C7553 INVX1_LOC_410/Y INVX1_LOC_519/A 0.03fF
C7554 INVX1_LOC_224/Y NAND2X1_LOC_123/A 0.07fF
C7555 NAND2X1_LOC_322/Y NAND2X1_LOC_775/B 0.05fF
C7556 VDD INVX1_LOC_35/Y 1.58fF
C7557 NAND2X1_LOC_756/Y INVX1_LOC_94/A 0.08fF
C7558 INVX1_LOC_53/Y NAND2X1_LOC_513/Y 0.21fF
C7559 VDD INVX1_LOC_304/A 0.00fF
C7560 INVX1_LOC_442/A NAND2X1_LOC_307/A 0.07fF
C7561 NAND2X1_LOC_780/B INVX1_LOC_549/Y 0.07fF
C7562 NAND2X1_LOC_830/a_36_24# INVX1_LOC_651/A 0.02fF
C7563 INVX1_LOC_442/A INVX1_LOC_545/Y 0.00fF
C7564 INVX1_LOC_578/A NAND2X1_LOC_123/A 0.12fF
C7565 INVX1_LOC_547/Y NAND2X1_LOC_253/a_36_24# 0.00fF
C7566 INVX1_LOC_561/A NAND2X1_LOC_591/B 0.00fF
C7567 INVX1_LOC_173/A INVX1_LOC_600/A 0.15fF
C7568 INVX1_LOC_228/Y INVX1_LOC_35/Y 0.21fF
C7569 INVX1_LOC_584/Y INVX1_LOC_186/A 0.01fF
C7570 INVX1_LOC_217/A NAND2X1_LOC_482/Y 0.05fF
C7571 INVX1_LOC_431/Y INVX1_LOC_596/Y 0.76fF
C7572 INVX1_LOC_11/Y INVX1_LOC_393/Y 0.07fF
C7573 VDD NAND2X1_LOC_448/B 0.16fF
C7574 INVX1_LOC_607/A INVX1_LOC_145/Y 0.02fF
C7575 VDD INVX1_LOC_572/Y 0.28fF
C7576 VDD INVX1_LOC_620/A 0.07fF
C7577 NAND2X1_LOC_27/Y INVX1_LOC_395/A 0.02fF
C7578 VDD NAND2X1_LOC_253/Y 0.12fF
C7579 INVX1_LOC_55/Y INVX1_LOC_29/Y 0.72fF
C7580 NAND2X1_LOC_241/B INVX1_LOC_208/A 0.00fF
C7581 INVX1_LOC_419/Y INVX1_LOC_442/A 0.00fF
C7582 INVX1_LOC_272/Y INVX1_LOC_635/A 0.26fF
C7583 NAND2X1_LOC_486/B INVX1_LOC_145/Y 0.01fF
C7584 INVX1_LOC_84/A NAND2X1_LOC_19/a_36_24# 0.00fF
C7585 NAND2X1_LOC_537/A INVX1_LOC_58/Y 0.04fF
C7586 INVX1_LOC_418/A INVX1_LOC_50/Y 0.06fF
C7587 VDD INVX1_LOC_621/Y 0.28fF
C7588 NAND2X1_LOC_540/a_36_24# INVX1_LOC_362/Y 0.00fF
C7589 INVX1_LOC_558/A INVX1_LOC_50/Y 0.07fF
C7590 NAND2X1_LOC_383/Y INVX1_LOC_48/Y 0.07fF
C7591 INVX1_LOC_312/Y INVX1_LOC_681/A 0.03fF
C7592 NAND2X1_LOC_307/A INVX1_LOC_116/Y 0.07fF
C7593 INVX1_LOC_373/A INVX1_LOC_496/A 0.03fF
C7594 INVX1_LOC_134/A INVX1_LOC_46/Y 0.06fF
C7595 INVX1_LOC_522/Y NAND2X1_LOC_708/A 0.03fF
C7596 INVX1_LOC_395/A INVX1_LOC_520/Y 0.05fF
C7597 INVX1_LOC_495/A INVX1_LOC_505/A 0.01fF
C7598 INVX1_LOC_545/Y INVX1_LOC_116/Y -0.03fF
C7599 INVX1_LOC_84/A INVX1_LOC_81/Y 0.01fF
C7600 INVX1_LOC_614/A INVX1_LOC_35/Y 0.04fF
C7601 INVX1_LOC_427/A INVX1_LOC_387/Y 0.01fF
C7602 INVX1_LOC_512/Y INVX1_LOC_463/Y 0.02fF
C7603 INVX1_LOC_358/Y INVX1_LOC_537/A -0.00fF
C7604 VDD INVX1_LOC_518/Y 0.21fF
C7605 INVX1_LOC_335/Y INVX1_LOC_537/A 0.07fF
C7606 INVX1_LOC_580/A INVX1_LOC_47/Y 0.01fF
C7607 INVX1_LOC_442/A NAND2X1_LOC_325/a_36_24# -0.00fF
C7608 NAND2X1_LOC_108/Y INVX1_LOC_58/Y 0.01fF
C7609 INVX1_LOC_381/A NAND2X1_LOC_347/a_36_24# 0.00fF
C7610 NAND2X1_LOC_475/A INVX1_LOC_153/Y 0.15fF
C7611 INVX1_LOC_664/A INVX1_LOC_445/A 0.05fF
C7612 INVX1_LOC_542/A INVX1_LOC_338/Y 0.01fF
C7613 INVX1_LOC_361/Y INVX1_LOC_80/A 0.06fF
C7614 NAND2X1_LOC_498/Y INVX1_LOC_301/Y 0.07fF
C7615 VDD INVX1_LOC_79/Y 0.21fF
C7616 INVX1_LOC_80/A NAND2X1_LOC_333/B 0.11fF
C7617 NAND2X1_LOC_45/Y INVX1_LOC_41/Y 0.03fF
C7618 INVX1_LOC_586/A INVX1_LOC_168/Y 0.05fF
C7619 INVX1_LOC_191/A INVX1_LOC_182/Y 0.16fF
C7620 INVX1_LOC_524/Y NAND2X1_LOC_753/Y 0.02fF
C7621 NAND2X1_LOC_782/A NAND2X1_LOC_677/Y 0.02fF
C7622 INVX1_LOC_17/Y INVX1_LOC_159/A 0.01fF
C7623 INVX1_LOC_299/Y INVX1_LOC_300/Y 0.09fF
C7624 INVX1_LOC_466/A INVX1_LOC_676/Y 0.00fF
C7625 NAND2X1_LOC_548/B INVX1_LOC_6/Y 0.03fF
C7626 INVX1_LOC_51/Y INVX1_LOC_245/A 0.06fF
C7627 INVX1_LOC_12/Y INVX1_LOC_230/Y 0.07fF
C7628 NAND2X1_LOC_858/a_36_24# INVX1_LOC_661/Y 0.00fF
C7629 INVX1_LOC_18/Y INVX1_LOC_29/Y 0.04fF
C7630 INVX1_LOC_40/Y INVX1_LOC_1/Y 0.03fF
C7631 NAND2X1_LOC_334/a_36_24# INVX1_LOC_674/A 0.01fF
C7632 NAND2X1_LOC_184/Y NAND2X1_LOC_260/Y 0.75fF
C7633 NAND2X1_LOC_755/B INVX1_LOC_50/Y 0.05fF
C7634 INVX1_LOC_358/Y INVX1_LOC_496/Y 1.13fF
C7635 INVX1_LOC_17/Y NAND2X1_LOC_615/B 0.07fF
C7636 INVX1_LOC_625/A NAND2X1_LOC_387/Y 0.02fF
C7637 INVX1_LOC_335/Y INVX1_LOC_496/Y 0.37fF
C7638 NAND2X1_LOC_307/A INVX1_LOC_255/A 0.19fF
C7639 INVX1_LOC_579/Y INVX1_LOC_261/Y 0.56fF
C7640 NAND2X1_LOC_703/a_36_24# INPUT_1 0.00fF
C7641 INVX1_LOC_80/A INVX1_LOC_258/Y 0.01fF
C7642 NAND2X1_LOC_498/Y INVX1_LOC_41/Y 0.22fF
C7643 INVX1_LOC_54/Y INVX1_LOC_352/Y 1.73fF
C7644 INPUT_1 INVX1_LOC_349/Y 0.00fF
C7645 INVX1_LOC_595/Y INVX1_LOC_623/Y 0.09fF
C7646 INVX1_LOC_211/Y INVX1_LOC_50/Y 0.00fF
C7647 INVX1_LOC_378/Y INVX1_LOC_489/Y 0.06fF
C7648 INVX1_LOC_103/Y INVX1_LOC_35/Y 0.03fF
C7649 INVX1_LOC_434/A INVX1_LOC_443/A 0.05fF
C7650 NAND2X1_LOC_781/A INVX1_LOC_168/Y 0.04fF
C7651 INVX1_LOC_11/Y INVX1_LOC_361/Y 1.08fF
C7652 INVX1_LOC_449/A INVX1_LOC_420/A 0.03fF
C7653 INVX1_LOC_310/Y NAND2X1_LOC_836/B 0.02fF
C7654 INVX1_LOC_266/A INVX1_LOC_245/A 0.00fF
C7655 INVX1_LOC_11/Y NAND2X1_LOC_333/B 0.03fF
C7656 INVX1_LOC_670/A INVX1_LOC_510/A 0.39fF
C7657 NAND2X1_LOC_570/a_36_24# INVX1_LOC_444/A 0.02fF
C7658 INVX1_LOC_6/Y INVX1_LOC_451/Y 0.01fF
C7659 INVX1_LOC_35/Y INVX1_LOC_68/A 0.02fF
C7660 INVX1_LOC_11/Y INVX1_LOC_281/A 0.05fF
C7661 NAND2X1_LOC_370/A INVX1_LOC_479/A 0.00fF
C7662 INVX1_LOC_685/Y INVX1_LOC_641/Y 0.05fF
C7663 INVX1_LOC_17/Y INVX1_LOC_66/A 0.05fF
C7664 INVX1_LOC_442/Y INVX1_LOC_234/Y 0.01fF
C7665 INVX1_LOC_480/Y INVX1_LOC_169/Y 0.04fF
C7666 INVX1_LOC_211/Y INVX1_LOC_431/Y 0.44fF
C7667 INVX1_LOC_134/Y INVX1_LOC_9/Y 0.07fF
C7668 INVX1_LOC_76/Y NAND2X1_LOC_123/B 0.00fF
C7669 NAND2X1_LOC_667/a_36_24# NAND2X1_LOC_333/B 0.00fF
C7670 INVX1_LOC_418/Y INVX1_LOC_89/Y 0.02fF
C7671 INVX1_LOC_564/A INVX1_LOC_91/Y 0.00fF
C7672 NAND2X1_LOC_325/a_36_24# INVX1_LOC_116/Y -0.02fF
C7673 INVX1_LOC_50/Y INVX1_LOC_46/Y 2.80fF
C7674 INVX1_LOC_89/Y INVX1_LOC_159/Y 0.13fF
C7675 INVX1_LOC_686/A INVX1_LOC_112/Y 0.03fF
C7676 INVX1_LOC_377/Y INVX1_LOC_41/Y 0.03fF
C7677 INVX1_LOC_469/Y INVX1_LOC_561/A 0.00fF
C7678 INVX1_LOC_419/Y INVX1_LOC_255/A 0.01fF
C7679 INVX1_LOC_183/A NAND2X1_LOC_400/a_36_24# 0.00fF
C7680 NAND2X1_LOC_106/Y INVX1_LOC_108/A 0.02fF
C7681 INVX1_LOC_166/Y INVX1_LOC_134/Y 0.06fF
C7682 INVX1_LOC_176/A INVX1_LOC_328/Y 0.16fF
C7683 INVX1_LOC_657/Y INVX1_LOC_59/A 0.01fF
C7684 INVX1_LOC_497/A INVX1_LOC_259/Y 0.01fF
C7685 NAND2X1_LOC_41/Y INVX1_LOC_9/Y 0.02fF
C7686 INVX1_LOC_93/Y NAND2X1_LOC_753/Y 0.07fF
C7687 INVX1_LOC_62/Y INVX1_LOC_134/Y 0.37fF
C7688 NAND2X1_LOC_514/a_36_24# INVX1_LOC_89/Y 0.00fF
C7689 INVX1_LOC_49/Y INPUT_1 0.28fF
C7690 INVX1_LOC_347/Y INVX1_LOC_354/Y 0.01fF
C7691 NAND2X1_LOC_307/B INVX1_LOC_66/A 0.21fF
C7692 INVX1_LOC_76/Y INVX1_LOC_270/Y 1.04fF
C7693 INVX1_LOC_517/Y INVX1_LOC_46/Y 0.01fF
C7694 NAND2X1_LOC_707/B INVX1_LOC_338/Y 0.03fF
C7695 INVX1_LOC_413/A INVX1_LOC_26/Y 0.01fF
C7696 INVX1_LOC_99/Y INVX1_LOC_41/Y 2.44fF
C7697 INVX1_LOC_298/A NAND2X1_LOC_823/a_36_24# 0.00fF
C7698 GATE_865 INVX1_LOC_632/Y 0.01fF
C7699 NAND2X1_LOC_770/B INVX1_LOC_26/Y 0.06fF
C7700 INVX1_LOC_298/A NAND2X1_LOC_291/a_36_24# 0.00fF
C7701 INVX1_LOC_76/Y INVX1_LOC_92/A 0.07fF
C7702 INVX1_LOC_670/A NAND2X1_LOC_477/a_36_24# 0.07fF
C7703 INVX1_LOC_58/Y INVX1_LOC_361/A 0.01fF
C7704 INVX1_LOC_681/Y INVX1_LOC_17/A 0.20fF
C7705 INVX1_LOC_35/Y INVX1_LOC_635/Y 0.03fF
C7706 INPUT_5 INVX1_LOC_69/Y 0.03fF
C7707 INVX1_LOC_47/Y INVX1_LOC_301/Y 0.03fF
C7708 INVX1_LOC_58/Y INVX1_LOC_196/Y 0.01fF
C7709 INVX1_LOC_6/Y NAND2X1_LOC_92/a_36_24# 0.00fF
C7710 INVX1_LOC_183/A INVX1_LOC_63/Y 0.21fF
C7711 NAND2X1_LOC_755/B INVX1_LOC_658/Y 0.05fF
C7712 INVX1_LOC_153/A INVX1_LOC_531/Y 0.04fF
C7713 INVX1_LOC_170/Y INVX1_LOC_328/Y 0.02fF
C7714 NAND2X1_LOC_285/A NAND2X1_LOC_248/a_36_24# 0.00fF
C7715 INVX1_LOC_368/A INVX1_LOC_49/Y 0.06fF
C7716 INVX1_LOC_123/A INVX1_LOC_41/Y 0.01fF
C7717 INVX1_LOC_93/Y INVX1_LOC_652/Y 0.01fF
C7718 INVX1_LOC_49/Y INVX1_LOC_487/Y 0.05fF
C7719 INVX1_LOC_338/Y INVX1_LOC_114/A 0.02fF
C7720 INVX1_LOC_89/Y INVX1_LOC_468/A 0.04fF
C7721 INVX1_LOC_96/A INVX1_LOC_531/Y 0.04fF
C7722 INVX1_LOC_74/Y INVX1_LOC_18/Y 0.01fF
C7723 INVX1_LOC_47/Y INVX1_LOC_41/Y 0.24fF
C7724 NAND2X1_LOC_292/Y INVX1_LOC_280/A 0.10fF
C7725 NAND2X1_LOC_557/B INVX1_LOC_41/Y 0.01fF
C7726 INPUT_0 NAND2X1_LOC_86/Y 0.49fF
C7727 INVX1_LOC_65/A INVX1_LOC_62/Y 0.00fF
C7728 NAND2X1_LOC_534/Y INVX1_LOC_409/A 0.02fF
C7729 INVX1_LOC_186/Y INVX1_LOC_611/A 0.02fF
C7730 NAND2X1_LOC_545/A INVX1_LOC_79/A 0.03fF
C7731 INVX1_LOC_317/Y NAND2X1_LOC_543/B 0.01fF
C7732 INVX1_LOC_63/Y INVX1_LOC_109/A 0.00fF
C7733 INVX1_LOC_41/Y INVX1_LOC_119/Y 0.12fF
C7734 INPUT_0 INVX1_LOC_206/Y 0.17fF
C7735 NAND2X1_LOC_261/Y INVX1_LOC_220/A 0.00fF
C7736 INVX1_LOC_75/Y INVX1_LOC_242/Y 0.16fF
C7737 INVX1_LOC_79/A INVX1_LOC_653/Y 0.20fF
C7738 NAND2X1_LOC_24/a_36_24# INVX1_LOC_206/Y 0.00fF
C7739 INVX1_LOC_269/A NAND2X1_LOC_76/B 0.30fF
C7740 NAND2X1_LOC_516/Y INVX1_LOC_206/Y 0.03fF
C7741 NAND2X1_LOC_631/B NAND2X1_LOC_625/a_36_24# 0.02fF
C7742 INVX1_LOC_79/A INVX1_LOC_666/Y 0.03fF
C7743 INVX1_LOC_206/Y INVX1_LOC_590/Y 0.03fF
C7744 NAND2X1_LOC_396/Y INVX1_LOC_325/A 0.07fF
C7745 INVX1_LOC_434/A NAND2X1_LOC_261/Y 0.01fF
C7746 INVX1_LOC_233/Y NAND2X1_LOC_271/B 0.08fF
C7747 INVX1_LOC_586/A NAND2X1_LOC_749/Y 0.47fF
C7748 VDD INVX1_LOC_256/Y 0.21fF
C7749 INVX1_LOC_409/Y INVX1_LOC_633/Y 0.02fF
C7750 INPUT_0 INVX1_LOC_242/A 0.03fF
C7751 NAND2X1_LOC_746/a_36_24# INVX1_LOC_53/Y 0.00fF
C7752 INVX1_LOC_3/Y INPUT_7 0.01fF
C7753 NAND2X1_LOC_526/Y INVX1_LOC_45/Y 0.03fF
C7754 INVX1_LOC_288/Y NAND2X1_LOC_761/a_36_24# 0.00fF
C7755 INVX1_LOC_393/A INVX1_LOC_392/Y 0.00fF
C7756 NAND2X1_LOC_791/B INVX1_LOC_292/A 0.21fF
C7757 NAND2X1_LOC_516/Y INVX1_LOC_242/A 0.00fF
C7758 INPUT_0 INVX1_LOC_686/A 0.12fF
C7759 INVX1_LOC_590/Y INVX1_LOC_396/Y 0.03fF
C7760 INPUT_1 INVX1_LOC_297/Y 0.14fF
C7761 NAND2X1_LOC_391/B INVX1_LOC_321/A 0.03fF
C7762 INVX1_LOC_21/Y NAND2X1_LOC_45/Y 0.03fF
C7763 INPUT_0 INVX1_LOC_80/Y 0.01fF
C7764 VDD INVX1_LOC_357/A -0.00fF
C7765 INVX1_LOC_629/Y INVX1_LOC_632/A 0.05fF
C7766 VDD INVX1_LOC_214/Y 0.39fF
C7767 INVX1_LOC_200/Y INVX1_LOC_670/Y 0.03fF
C7768 INVX1_LOC_97/A INVX1_LOC_600/A 0.29fF
C7769 NAND2X1_LOC_390/a_36_24# NAND2X1_LOC_13/Y 0.00fF
C7770 INVX1_LOC_224/Y INVX1_LOC_145/Y 0.07fF
C7771 INVX1_LOC_438/Y INVX1_LOC_17/Y 0.06fF
C7772 INVX1_LOC_607/Y INVX1_LOC_206/Y 0.09fF
C7773 INVX1_LOC_549/A INVX1_LOC_161/A 0.07fF
C7774 VDD NAND2X1_LOC_837/B 0.05fF
C7775 INPUT_0 INVX1_LOC_14/A 0.01fF
C7776 NAND2X1_LOC_534/Y INVX1_LOC_352/Y 0.01fF
C7777 INVX1_LOC_171/Y INVX1_LOC_172/Y 0.01fF
C7778 NAND2X1_LOC_56/Y INVX1_LOC_173/A 0.15fF
C7779 VDD INVX1_LOC_673/Y 0.16fF
C7780 INVX1_LOC_21/Y NAND2X1_LOC_498/Y 0.07fF
C7781 VDD INVX1_LOC_118/A 0.00fF
C7782 INVX1_LOC_21/Y INVX1_LOC_570/A 0.03fF
C7783 INVX1_LOC_607/Y INVX1_LOC_648/Y 0.06fF
C7784 VDD INVX1_LOC_208/A -0.00fF
C7785 INVX1_LOC_463/A NAND2X1_LOC_689/B 0.05fF
C7786 INVX1_LOC_201/Y INVX1_LOC_395/A 0.09fF
C7787 INVX1_LOC_578/A INVX1_LOC_145/Y 0.08fF
C7788 NAND2X1_LOC_728/B NAND2X1_LOC_680/a_36_24# 0.02fF
C7789 INVX1_LOC_160/Y INVX1_LOC_99/Y 0.16fF
C7790 INVX1_LOC_53/A NAND2X1_LOC_18/a_36_24# 0.00fF
C7791 NAND2X1_LOC_751/a_36_24# INVX1_LOC_198/A 0.00fF
C7792 INVX1_LOC_20/Y NAND2X1_LOC_299/Y 0.56fF
C7793 INVX1_LOC_99/A INVX1_LOC_586/A 0.01fF
C7794 INVX1_LOC_17/Y INVX1_LOC_442/A 0.07fF
C7795 INVX1_LOC_438/A INVX1_LOC_46/Y 0.07fF
C7796 INVX1_LOC_206/Y INVX1_LOC_298/A 0.04fF
C7797 INVX1_LOC_625/A INVX1_LOC_269/A 0.33fF
C7798 INVX1_LOC_224/Y INVX1_LOC_248/A 0.01fF
C7799 INVX1_LOC_169/A INVX1_LOC_600/A 0.94fF
C7800 INVX1_LOC_206/Y INVX1_LOC_498/A 0.03fF
C7801 NAND2X1_LOC_710/A INVX1_LOC_53/Y 0.01fF
C7802 NAND2X1_LOC_164/Y NAND2X1_LOC_387/Y 0.08fF
C7803 INVX1_LOC_320/Y INVX1_LOC_48/Y 0.01fF
C7804 INVX1_LOC_53/Y INVX1_LOC_508/Y 0.01fF
C7805 INVX1_LOC_563/Y INVX1_LOC_93/Y 0.02fF
C7806 INVX1_LOC_543/Y INVX1_LOC_395/A 0.07fF
C7807 INVX1_LOC_607/Y INVX1_LOC_242/A 0.07fF
C7808 NAND2X1_LOC_636/A NAND2X1_LOC_192/A 0.28fF
C7809 NAND2X1_LOC_409/Y INVX1_LOC_41/A 0.01fF
C7810 INVX1_LOC_586/A INVX1_LOC_137/Y 0.03fF
C7811 INVX1_LOC_174/Y INVX1_LOC_81/Y 0.02fF
C7812 INVX1_LOC_38/A INVX1_LOC_194/Y 0.03fF
C7813 INVX1_LOC_516/Y INVX1_LOC_137/Y 0.04fF
C7814 INVX1_LOC_686/A NAND2X1_LOC_123/A 0.02fF
C7815 INVX1_LOC_43/Y INVX1_LOC_184/A 0.01fF
C7816 INVX1_LOC_530/Y INVX1_LOC_50/Y 0.04fF
C7817 INVX1_LOC_463/A INVX1_LOC_245/A 0.26fF
C7818 INVX1_LOC_65/Y NAND2X1_LOC_387/Y 0.08fF
C7819 INVX1_LOC_678/Y INVX1_LOC_678/A 0.01fF
C7820 INVX1_LOC_312/Y NAND2X1_LOC_862/a_36_24# 0.01fF
C7821 INVX1_LOC_45/Y NAND2X1_LOC_619/Y 0.01fF
C7822 INPUT_0 NAND2X1_LOC_334/A 0.00fF
C7823 INVX1_LOC_371/Y INVX1_LOC_377/A 0.07fF
C7824 INVX1_LOC_570/A INVX1_LOC_555/A 0.08fF
C7825 INVX1_LOC_442/Y INVX1_LOC_80/A 0.14fF
C7826 INVX1_LOC_603/Y INVX1_LOC_604/Y 0.06fF
C7827 INVX1_LOC_76/Y INPUT_1 0.94fF
C7828 INVX1_LOC_447/Y INVX1_LOC_449/A 0.18fF
C7829 NAND2X1_LOC_575/a_36_24# NAND2X1_LOC_274/B 0.00fF
C7830 NAND2X1_LOC_750/Y INVX1_LOC_223/Y 0.00fF
C7831 INVX1_LOC_268/Y INVX1_LOC_50/Y 0.00fF
C7832 NAND2X1_LOC_685/B INVX1_LOC_463/Y 0.03fF
C7833 INVX1_LOC_513/A NAND2X1_LOC_644/a_36_24# 0.00fF
C7834 INVX1_LOC_551/Y INVX1_LOC_117/Y 0.10fF
C7835 INVX1_LOC_335/Y INVX1_LOC_99/Y 0.03fF
C7836 INVX1_LOC_617/A INVX1_LOC_166/A 0.01fF
C7837 NAND2X1_LOC_69/a_36_24# INVX1_LOC_63/Y 0.00fF
C7838 INVX1_LOC_21/Y INVX1_LOC_99/Y 0.14fF
C7839 INVX1_LOC_124/Y INVX1_LOC_669/Y 0.34fF
C7840 INVX1_LOC_617/Y INVX1_LOC_670/A 0.00fF
C7841 NAND2X1_LOC_169/A INVX1_LOC_252/Y 0.01fF
C7842 INVX1_LOC_686/A INVX1_LOC_498/A 0.07fF
C7843 INVX1_LOC_449/A INVX1_LOC_54/Y 0.10fF
C7844 INVX1_LOC_17/Y INVX1_LOC_116/Y 0.10fF
C7845 INVX1_LOC_270/A NAND2X1_LOC_388/A 0.00fF
C7846 INVX1_LOC_9/Y NAND2X1_LOC_249/a_36_24# 0.00fF
C7847 NAND2X1_LOC_475/A INVX1_LOC_41/Y 0.19fF
C7848 INVX1_LOC_93/Y INVX1_LOC_197/A 10.96fF
C7849 INVX1_LOC_490/Y INVX1_LOC_79/A 0.05fF
C7850 INVX1_LOC_11/Y INVX1_LOC_442/Y 0.07fF
C7851 VDD INVX1_LOC_495/Y 0.36fF
C7852 INVX1_LOC_400/Y INVX1_LOC_128/Y 0.04fF
C7853 NAND2X1_LOC_383/Y NAND2X1_LOC_615/Y 0.69fF
C7854 VDD INVX1_LOC_364/A -0.00fF
C7855 INVX1_LOC_150/A INVX1_LOC_479/A 0.09fF
C7856 NAND2X1_LOC_513/A INVX1_LOC_46/Y 0.07fF
C7857 INVX1_LOC_116/A INVX1_LOC_360/A 0.00fF
C7858 INPUT_0 NAND2X1_LOC_609/B 0.17fF
C7859 INVX1_LOC_680/Y INVX1_LOC_105/Y 0.01fF
C7860 INVX1_LOC_502/Y INVX1_LOC_301/Y 0.07fF
C7861 INVX1_LOC_561/A INVX1_LOC_632/A 0.04fF
C7862 NAND2X1_LOC_152/Y NAND2X1_LOC_846/B 0.15fF
C7863 INVX1_LOC_330/A INVX1_LOC_137/Y 0.05fF
C7864 INVX1_LOC_53/Y INVX1_LOC_633/A 0.02fF
C7865 NAND2X1_LOC_16/Y INVX1_LOC_79/A 0.01fF
C7866 NAND2X1_LOC_307/A INVX1_LOC_69/Y 0.03fF
C7867 INVX1_LOC_575/A INVX1_LOC_575/Y 0.19fF
C7868 INVX1_LOC_93/Y INVX1_LOC_124/Y 0.01fF
C7869 INVX1_LOC_105/A INVX1_LOC_35/Y 0.34fF
C7870 NAND2X1_LOC_541/B NAND2X1_LOC_274/Y 0.02fF
C7871 INVX1_LOC_171/A INVX1_LOC_35/Y 0.32fF
C7872 INVX1_LOC_99/Y NAND2X1_LOC_267/A 0.47fF
C7873 NAND2X1_LOC_527/Y INVX1_LOC_145/Y 0.00fF
C7874 INVX1_LOC_662/A NAND2X1_LOC_149/a_36_24# 0.01fF
C7875 INVX1_LOC_62/A INVX1_LOC_556/Y 0.03fF
C7876 INVX1_LOC_602/A NAND2X1_LOC_759/Y 0.02fF
C7877 INVX1_LOC_21/Y INVX1_LOC_589/Y 0.06fF
C7878 VDD INVX1_LOC_488/Y 0.51fF
C7879 INVX1_LOC_206/Y INVX1_LOC_211/A 0.43fF
C7880 INVX1_LOC_603/Y INVX1_LOC_397/Y 0.01fF
C7881 NAND2X1_LOC_13/Y INVX1_LOC_245/A 1.06fF
C7882 INVX1_LOC_76/Y INVX1_LOC_368/A 0.04fF
C7883 INVX1_LOC_593/Y INVX1_LOC_631/A 0.04fF
C7884 NAND2X1_LOC_294/Y INVX1_LOC_451/Y 0.02fF
C7885 INVX1_LOC_335/Y INVX1_LOC_47/Y 9.14fF
C7886 INVX1_LOC_628/Y INVX1_LOC_261/Y 0.01fF
C7887 INVX1_LOC_21/Y INVX1_LOC_47/Y 0.37fF
C7888 INVX1_LOC_76/Y INVX1_LOC_487/Y 0.01fF
C7889 INVX1_LOC_174/A INVX1_LOC_63/Y 0.08fF
C7890 INVX1_LOC_145/Y INVX1_LOC_93/A 0.00fF
C7891 INVX1_LOC_21/Y NAND2X1_LOC_557/B 0.01fF
C7892 INVX1_LOC_428/Y INVX1_LOC_387/Y 0.02fF
C7893 INVX1_LOC_382/Y INVX1_LOC_385/A 0.15fF
C7894 INVX1_LOC_47/Y NAND2X1_LOC_655/a_36_24# 0.01fF
C7895 INVX1_LOC_566/A NAND2X1_LOC_806/a_36_24# 0.00fF
C7896 INVX1_LOC_167/A INVX1_LOC_117/Y 0.01fF
C7897 INVX1_LOC_581/A NAND2X1_LOC_780/a_36_24# 0.00fF
C7898 INVX1_LOC_17/Y INVX1_LOC_255/A 0.07fF
C7899 INVX1_LOC_89/Y INVX1_LOC_352/Y 0.01fF
C7900 INVX1_LOC_107/Y INVX1_LOC_99/Y 0.12fF
C7901 NAND2X1_LOC_707/A INVX1_LOC_505/Y 0.02fF
C7902 INVX1_LOC_46/Y INVX1_LOC_327/Y 0.01fF
C7903 NAND2X1_LOC_387/Y INVX1_LOC_318/A 0.03fF
C7904 INVX1_LOC_298/A INVX1_LOC_342/A 0.20fF
C7905 INVX1_LOC_387/Y INVX1_LOC_50/Y 0.03fF
C7906 INVX1_LOC_419/Y INVX1_LOC_69/Y 0.20fF
C7907 INVX1_LOC_20/Y INVX1_LOC_75/Y 0.08fF
C7908 INVX1_LOC_17/Y INVX1_LOC_179/A 0.07fF
C7909 INVX1_LOC_356/A INVX1_LOC_479/A 0.00fF
C7910 NAND2X1_LOC_387/Y INVX1_LOC_397/Y 0.03fF
C7911 INVX1_LOC_17/Y NAND2X1_LOC_719/A 0.02fF
C7912 NAND2X1_LOC_388/A INVX1_LOC_46/Y 0.03fF
C7913 INVX1_LOC_21/Y INVX1_LOC_119/Y 0.03fF
C7914 NAND2X1_LOC_174/B INVX1_LOC_675/A 0.05fF
C7915 INVX1_LOC_117/Y INVX1_LOC_486/A 0.01fF
C7916 NAND2X1_LOC_148/B NAND2X1_LOC_342/A 0.03fF
C7917 INVX1_LOC_21/Y NAND2X1_LOC_66/Y 0.08fF
C7918 INVX1_LOC_49/Y INVX1_LOC_50/Y 4.09fF
C7919 INVX1_LOC_504/A INVX1_LOC_114/A 0.08fF
C7920 INVX1_LOC_382/A INVX1_LOC_378/Y 0.00fF
C7921 INVX1_LOC_6/Y NAND2X1_LOC_647/A 0.01fF
C7922 NAND2X1_LOC_591/Y INVX1_LOC_675/A 0.04fF
C7923 NAND2X1_LOC_387/Y INVX1_LOC_95/A 0.01fF
C7924 NAND2X1_LOC_655/a_36_24# INVX1_LOC_119/Y 0.00fF
C7925 INVX1_LOC_54/Y INVX1_LOC_328/Y 0.03fF
C7926 INVX1_LOC_188/Y INVX1_LOC_588/A 0.03fF
C7927 INVX1_LOC_25/Y INVX1_LOC_41/Y 0.55fF
C7928 INVX1_LOC_612/Y INVX1_LOC_612/A 0.01fF
C7929 NAND2X1_LOC_791/A INVX1_LOC_621/A 0.20fF
C7930 INVX1_LOC_417/Y INVX1_LOC_666/Y 0.07fF
C7931 INVX1_LOC_145/Y INVX1_LOC_621/A 0.00fF
C7932 INVX1_LOC_41/Y NAND2X1_LOC_276/a_36_24# 0.00fF
C7933 INVX1_LOC_300/A INVX1_LOC_75/Y 0.10fF
C7934 NAND2X1_LOC_545/A INVX1_LOC_48/Y 0.03fF
C7935 INVX1_LOC_376/A INVX1_LOC_69/Y 0.19fF
C7936 NAND2X1_LOC_184/Y INVX1_LOC_655/A 0.03fF
C7937 INVX1_LOC_421/A INVX1_LOC_26/Y 0.15fF
C7938 INVX1_LOC_204/Y INVX1_LOC_622/A 0.01fF
C7939 NAND2X1_LOC_837/B INVX1_LOC_635/Y 0.00fF
C7940 INVX1_LOC_380/Y INVX1_LOC_245/A 0.01fF
C7941 INVX1_LOC_100/A INVX1_LOC_100/Y 0.00fF
C7942 INVX1_LOC_361/A INVX1_LOC_245/A 0.11fF
C7943 NAND2X1_LOC_737/a_36_24# INVX1_LOC_636/A 0.01fF
C7944 INVX1_LOC_69/Y INVX1_LOC_502/A 0.08fF
C7945 INVX1_LOC_666/Y INVX1_LOC_48/Y 0.03fF
C7946 INVX1_LOC_117/Y NAND2X1_LOC_410/Y -0.00fF
C7947 INVX1_LOC_31/Y INVX1_LOC_652/Y 0.02fF
C7948 INVX1_LOC_103/Y INVX1_LOC_364/A 0.00fF
C7949 INVX1_LOC_31/Y INVX1_LOC_483/A 0.04fF
C7950 INVX1_LOC_90/Y INVX1_LOC_9/Y 0.07fF
C7951 NAND2X1_LOC_333/B INVX1_LOC_91/Y 0.11fF
C7952 INVX1_LOC_491/A NAND2X1_LOC_633/a_36_24# 0.01fF
C7953 INVX1_LOC_89/Y NAND2X1_LOC_438/a_36_24# 0.01fF
C7954 INVX1_LOC_556/Y INVX1_LOC_76/A 0.02fF
C7955 VDD INVX1_LOC_434/A 0.14fF
C7956 INVX1_LOC_15/Y INVX1_LOC_41/Y 0.14fF
C7957 INVX1_LOC_191/Y INVX1_LOC_195/A 0.00fF
C7958 INVX1_LOC_32/Y INVX1_LOC_270/Y 0.05fF
C7959 VDD INVX1_LOC_52/Y 0.21fF
C7960 INVX1_LOC_62/Y NAND2X1_LOC_221/a_36_24# 0.00fF
C7961 INVX1_LOC_531/Y INVX1_LOC_353/A 0.04fF
C7962 INVX1_LOC_507/A NAND2X1_LOC_646/B 0.06fF
C7963 INVX1_LOC_32/Y INVX1_LOC_92/A 0.12fF
C7964 INVX1_LOC_49/Y INVX1_LOC_658/Y 0.09fF
C7965 INVX1_LOC_62/Y INVX1_LOC_90/Y 0.11fF
C7966 INPUT_0 INVX1_LOC_390/Y 0.03fF
C7967 INVX1_LOC_491/A INVX1_LOC_588/A 0.07fF
C7968 INVX1_LOC_680/Y INVX1_LOC_109/Y 0.01fF
C7969 INVX1_LOC_563/Y INVX1_LOC_395/A 0.03fF
C7970 INVX1_LOC_435/Y NAND2X1_LOC_457/A 0.03fF
C7971 NAND2X1_LOC_475/A INVX1_LOC_160/Y 0.01fF
C7972 INVX1_LOC_400/Y INVX1_LOC_560/A 0.07fF
C7973 INVX1_LOC_206/Y INVX1_LOC_288/A 0.07fF
C7974 INVX1_LOC_346/Y INVX1_LOC_114/A 0.02fF
C7975 INVX1_LOC_435/Y INVX1_LOC_547/Y 0.10fF
C7976 INVX1_LOC_604/A INVX1_LOC_273/A 0.03fF
C7977 INVX1_LOC_145/Y NAND2X1_LOC_86/Y 0.01fF
C7978 NAND2X1_LOC_269/B NAND2X1_LOC_271/A 0.10fF
C7979 INVX1_LOC_257/Y INVX1_LOC_686/A 0.02fF
C7980 INVX1_LOC_202/Y INVX1_LOC_275/A 0.02fF
C7981 VDD INVX1_LOC_115/Y 0.23fF
C7982 INVX1_LOC_21/Y NAND2X1_LOC_475/A 0.07fF
C7983 NAND2X1_LOC_331/A INVX1_LOC_134/Y 0.00fF
C7984 INVX1_LOC_412/A INVX1_LOC_80/A 0.00fF
C7985 INVX1_LOC_288/A INVX1_LOC_686/A 0.04fF
C7986 VDD INVX1_LOC_350/A -0.00fF
C7987 INVX1_LOC_431/Y INVX1_LOC_297/Y 0.04fF
C7988 INVX1_LOC_541/Y INVX1_LOC_542/A 0.00fF
C7989 INVX1_LOC_434/A NAND2X1_LOC_556/a_36_24# 0.01fF
C7990 INVX1_LOC_206/Y INVX1_LOC_145/Y 0.37fF
C7991 INVX1_LOC_428/A NAND2X1_LOC_496/Y 0.03fF
C7992 NAND2X1_LOC_307/A INVX1_LOC_586/A 0.11fF
C7993 INVX1_LOC_224/Y INVX1_LOC_440/A 0.01fF
C7994 INVX1_LOC_404/Y INVX1_LOC_235/A 0.01fF
C7995 INVX1_LOC_445/Y INVX1_LOC_444/Y 0.02fF
C7996 INPUT_0 INVX1_LOC_432/A 0.07fF
C7997 INVX1_LOC_412/Y NAND2X1_LOC_603/a_36_24# 0.00fF
C7998 INVX1_LOC_3/Y INVX1_LOC_18/Y 0.00fF
C7999 NAND2X1_LOC_475/A NAND2X1_LOC_267/A 1.22fF
C8000 INVX1_LOC_45/Y INVX1_LOC_379/A 0.07fF
C8001 INVX1_LOC_428/A NAND2X1_LOC_257/a_36_24# 0.00fF
C8002 INVX1_LOC_545/A INVX1_LOC_442/A 0.02fF
C8003 INVX1_LOC_602/A INVX1_LOC_333/A 0.02fF
C8004 INVX1_LOC_35/Y NAND2X1_LOC_506/B 0.04fF
C8005 INVX1_LOC_185/Y INVX1_LOC_35/Y 0.04fF
C8006 INVX1_LOC_45/Y INVX1_LOC_35/Y 10.57fF
C8007 INVX1_LOC_435/A INVX1_LOC_321/A 0.18fF
C8008 INVX1_LOC_577/Y INVX1_LOC_99/Y 1.16fF
C8009 INVX1_LOC_410/Y INVX1_LOC_670/A 0.00fF
C8010 VDD INVX1_LOC_378/Y 0.21fF
C8011 NAND2X1_LOC_93/Y INVX1_LOC_49/Y 0.10fF
C8012 INVX1_LOC_416/A INVX1_LOC_586/A 0.01fF
C8013 VDD NAND2X1_LOC_686/B 0.01fF
C8014 INVX1_LOC_375/A INVX1_LOC_670/A 0.19fF
C8015 INVX1_LOC_428/A NAND2X1_LOC_706/B 0.11fF
C8016 INVX1_LOC_6/Y NAND2X1_LOC_749/Y 0.03fF
C8017 INVX1_LOC_419/Y INVX1_LOC_586/A 0.11fF
C8018 VDD INVX1_LOC_507/Y 0.32fF
C8019 NAND2X1_LOC_710/B INVX1_LOC_47/Y 0.03fF
C8020 INVX1_LOC_438/A INVX1_LOC_49/Y 0.08fF
C8021 INPUT_0 NAND2X1_LOC_542/A 0.07fF
C8022 VDD INVX1_LOC_223/Y 0.22fF
C8023 INVX1_LOC_602/A NAND2X1_LOC_755/B 0.02fF
C8024 INVX1_LOC_686/A INVX1_LOC_145/Y 0.07fF
C8025 INVX1_LOC_401/Y INVX1_LOC_516/A 0.22fF
C8026 INPUT_3 INVX1_LOC_35/Y 0.06fF
C8027 INVX1_LOC_620/A NAND2X1_LOC_506/B 0.05fF
C8028 NAND2X1_LOC_313/a_36_24# INVX1_LOC_510/Y 0.01fF
C8029 VDD INVX1_LOC_667/Y 0.21fF
C8030 INVX1_LOC_237/Y INVX1_LOC_523/Y 0.03fF
C8031 INVX1_LOC_76/Y INVX1_LOC_50/Y 0.16fF
C8032 INVX1_LOC_84/A INVX1_LOC_304/Y 0.01fF
C8033 INVX1_LOC_45/Y INVX1_LOC_620/A 0.03fF
C8034 INVX1_LOC_45/Y NAND2X1_LOC_253/Y 0.01fF
C8035 NAND2X1_LOC_516/Y NAND2X1_LOC_542/A 0.04fF
C8036 INVX1_LOC_320/A INVX1_LOC_230/A 0.11fF
C8037 NAND2X1_LOC_547/a_36_24# INVX1_LOC_51/Y 0.00fF
C8038 INVX1_LOC_556/A INVX1_LOC_63/Y 0.21fF
C8039 INVX1_LOC_407/Y INVX1_LOC_134/Y 0.03fF
C8040 INVX1_LOC_51/Y NAND2X1_LOC_753/Y 0.07fF
C8041 NAND2X1_LOC_45/Y INVX1_LOC_26/Y 0.08fF
C8042 NAND2X1_LOC_543/B INVX1_LOC_41/Y 0.02fF
C8043 NAND2X1_LOC_391/A INVX1_LOC_159/Y 0.04fF
C8044 INVX1_LOC_335/Y INVX1_LOC_25/Y 0.11fF
C8045 INVX1_LOC_76/Y INVX1_LOC_431/Y 0.03fF
C8046 INVX1_LOC_224/Y INVX1_LOC_242/Y 0.54fF
C8047 INVX1_LOC_581/A NAND2X1_LOC_708/A 0.08fF
C8048 INPUT_5 INVX1_LOC_1/A 0.04fF
C8049 INVX1_LOC_288/A NAND2X1_LOC_334/A 0.07fF
C8050 INVX1_LOC_584/Y INVX1_LOC_501/A 0.03fF
C8051 INVX1_LOC_115/Y INVX1_LOC_116/A 0.02fF
C8052 INVX1_LOC_577/Y INVX1_LOC_47/Y 0.01fF
C8053 NAND2X1_LOC_318/A NAND2X1_LOC_388/A 0.00fF
C8054 INVX1_LOC_442/Y INVX1_LOC_367/Y 0.07fF
C8055 NAND2X1_LOC_710/B INVX1_LOC_119/Y 0.01fF
C8056 INVX1_LOC_5/Y INVX1_LOC_3/A 0.01fF
C8057 INVX1_LOC_99/Y INVX1_LOC_481/Y 0.01fF
C8058 NAND2X1_LOC_720/A INVX1_LOC_635/A 0.05fF
C8059 INVX1_LOC_89/Y NAND2X1_LOC_159/a_36_24# 0.00fF
C8060 NAND2X1_LOC_516/Y INVX1_LOC_376/Y 0.07fF
C8061 INVX1_LOC_444/Y INVX1_LOC_99/Y 0.05fF
C8062 INVX1_LOC_524/Y INVX1_LOC_525/Y 0.08fF
C8063 INVX1_LOC_569/A INVX1_LOC_6/Y 0.30fF
C8064 INVX1_LOC_428/Y INVX1_LOC_386/Y 0.01fF
C8065 INVX1_LOC_545/A INVX1_LOC_116/Y 0.03fF
C8066 INVX1_LOC_2/Y INVX1_LOC_1/A 0.00fF
C8067 INVX1_LOC_308/Y INVX1_LOC_100/Y 0.02fF
C8068 INVX1_LOC_578/A INVX1_LOC_242/Y 0.04fF
C8069 INVX1_LOC_342/Y INVX1_LOC_685/A 0.05fF
C8070 INVX1_LOC_31/Y INVX1_LOC_197/A 0.07fF
C8071 INVX1_LOC_267/Y INVX1_LOC_93/Y 0.03fF
C8072 NAND2X1_LOC_677/Y INVX1_LOC_186/Y 0.14fF
C8073 NAND2X1_LOC_636/B INVX1_LOC_46/Y 0.01fF
C8074 INVX1_LOC_76/Y INVX1_LOC_517/Y 0.01fF
C8075 NAND2X1_LOC_498/Y INVX1_LOC_128/Y 0.04fF
C8076 NAND2X1_LOC_97/B INVX1_LOC_93/Y 0.02fF
C8077 INVX1_LOC_551/Y INVX1_LOC_58/Y 0.01fF
C8078 INVX1_LOC_166/A NAND2X1_LOC_130/Y 0.03fF
C8079 INVX1_LOC_43/Y INVX1_LOC_86/Y 0.02fF
C8080 INPUT_1 INVX1_LOC_7/Y 0.00fF
C8081 INVX1_LOC_117/Y NAND2X1_LOC_755/B 0.03fF
C8082 INVX1_LOC_293/Y INVX1_LOC_654/Y 0.09fF
C8083 INVX1_LOC_360/Y INVX1_LOC_360/A 0.01fF
C8084 INVX1_LOC_376/A NAND2X1_LOC_440/a_36_24# 0.00fF
C8085 INVX1_LOC_617/A INVX1_LOC_301/Y 0.00fF
C8086 INVX1_LOC_68/Y INVX1_LOC_153/Y 0.00fF
C8087 INVX1_LOC_586/A INVX1_LOC_502/A 0.07fF
C8088 INVX1_LOC_89/Y INVX1_LOC_67/Y 0.03fF
C8089 INVX1_LOC_274/A INVX1_LOC_395/Y 0.02fF
C8090 INVX1_LOC_84/A INVX1_LOC_183/A 0.04fF
C8091 INVX1_LOC_211/Y INVX1_LOC_117/Y 0.03fF
C8092 INVX1_LOC_421/A NAND2X1_LOC_275/Y 0.02fF
C8093 INVX1_LOC_431/A INVX1_LOC_48/Y 0.01fF
C8094 INVX1_LOC_80/A NAND2X1_LOC_847/A 0.08fF
C8095 NAND2X1_LOC_862/a_36_24# INVX1_LOC_6/Y 0.00fF
C8096 INVX1_LOC_188/Y INVX1_LOC_63/Y 0.03fF
C8097 INVX1_LOC_93/Y INVX1_LOC_510/A 0.07fF
C8098 INVX1_LOC_662/A INVX1_LOC_508/Y 0.00fF
C8099 INVX1_LOC_54/Y INVX1_LOC_172/A 0.09fF
C8100 INVX1_LOC_68/Y INVX1_LOC_531/Y 0.02fF
C8101 INVX1_LOC_603/Y INVX1_LOC_63/Y 5.28fF
C8102 INVX1_LOC_93/Y INVX1_LOC_440/Y 0.16fF
C8103 INVX1_LOC_377/Y INVX1_LOC_128/Y 0.02fF
C8104 INVX1_LOC_51/Y INVX1_LOC_652/Y 0.05fF
C8105 NAND2X1_LOC_709/a_36_24# INVX1_LOC_600/A 0.01fF
C8106 INVX1_LOC_17/Y INVX1_LOC_69/Y 0.50fF
C8107 NAND2X1_LOC_174/B INVX1_LOC_31/Y 0.03fF
C8108 INVX1_LOC_137/Y INVX1_LOC_6/Y 0.04fF
C8109 INVX1_LOC_100/Y NAND2X1_LOC_846/a_36_24# 0.00fF
C8110 INVX1_LOC_545/A INVX1_LOC_255/A 0.06fF
C8111 INVX1_LOC_617/A INVX1_LOC_41/Y 0.01fF
C8112 INVX1_LOC_32/Y INPUT_1 0.11fF
C8113 INVX1_LOC_117/Y INVX1_LOC_46/Y 0.71fF
C8114 INVX1_LOC_298/Y INVX1_LOC_58/Y 0.17fF
C8115 INVX1_LOC_211/A INVX1_LOC_94/A 0.01fF
C8116 INVX1_LOC_366/A NAND2X1_LOC_234/Y 0.00fF
C8117 INVX1_LOC_133/A INVX1_LOC_241/A 0.03fF
C8118 INVX1_LOC_93/Y NAND2X1_LOC_128/A 0.01fF
C8119 NAND2X1_LOC_192/a_36_24# INVX1_LOC_62/Y 0.00fF
C8120 INVX1_LOC_93/Y INVX1_LOC_525/Y 0.09fF
C8121 INVX1_LOC_184/A INVX1_LOC_190/A 0.48fF
C8122 INVX1_LOC_100/Y NAND2X1_LOC_237/Y 0.01fF
C8123 INVX1_LOC_99/Y NAND2X1_LOC_420/a_36_24# 0.01fF
C8124 INVX1_LOC_493/A INVX1_LOC_58/Y 0.00fF
C8125 INVX1_LOC_9/Y INVX1_LOC_98/Y 0.21fF
C8126 INVX1_LOC_275/Y INVX1_LOC_79/A 0.05fF
C8127 INVX1_LOC_99/Y INVX1_LOC_26/Y 3.56fF
C8128 INVX1_LOC_167/A INVX1_LOC_58/Y 0.00fF
C8129 NAND2X1_LOC_788/a_36_24# INVX1_LOC_376/Y 0.00fF
C8130 NAND2X1_LOC_545/B INVX1_LOC_62/Y 0.00fF
C8131 INVX1_LOC_487/Y INVX1_LOC_7/Y 0.01fF
C8132 NAND2X1_LOC_387/Y INVX1_LOC_63/Y 0.07fF
C8133 NAND2X1_LOC_274/B INVX1_LOC_252/Y 0.01fF
C8134 INVX1_LOC_406/A INVX1_LOC_6/Y 0.03fF
C8135 INVX1_LOC_531/Y INVX1_LOC_600/A 0.09fF
C8136 NAND2X1_LOC_663/a_36_24# INVX1_LOC_66/A 0.00fF
C8137 INVX1_LOC_523/Y INVX1_LOC_212/Y 0.06fF
C8138 INVX1_LOC_100/Y INVX1_LOC_230/A 0.07fF
C8139 INVX1_LOC_481/Y NAND2X1_LOC_66/Y 0.01fF
C8140 INVX1_LOC_444/Y NAND2X1_LOC_66/Y 1.24fF
C8141 INVX1_LOC_492/A INVX1_LOC_655/A 0.02fF
C8142 NAND2X1_LOC_858/a_36_24# INVX1_LOC_655/A 0.01fF
C8143 INVX1_LOC_491/A NAND2X1_LOC_646/A 0.04fF
C8144 INVX1_LOC_435/A NAND2X1_LOC_268/a_36_24# 0.00fF
C8145 INVX1_LOC_99/Y NAND2X1_LOC_608/a_36_24# -0.00fF
C8146 INVX1_LOC_67/Y NAND2X1_LOC_544/B 0.09fF
C8147 INVX1_LOC_89/Y INVX1_LOC_347/Y 0.00fF
C8148 NAND2X1_LOC_549/a_36_24# INVX1_LOC_6/Y 0.01fF
C8149 INVX1_LOC_410/A INVX1_LOC_199/Y 0.03fF
C8150 NAND2X1_LOC_489/A INVX1_LOC_48/Y 0.01fF
C8151 NAND2X1_LOC_448/A INVX1_LOC_354/A 0.09fF
C8152 INVX1_LOC_62/Y INVX1_LOC_98/Y 0.22fF
C8153 INVX1_LOC_240/A INVX1_LOC_655/A 0.04fF
C8154 INVX1_LOC_41/Y INVX1_LOC_505/A 0.09fF
C8155 INVX1_LOC_93/Y NAND2X1_LOC_477/a_36_24# 0.01fF
C8156 INVX1_LOC_352/Y INVX1_LOC_347/A 0.07fF
C8157 INVX1_LOC_501/A INVX1_LOC_347/Y 0.03fF
C8158 INVX1_LOC_399/Y INVX1_LOC_199/Y 0.15fF
C8159 INVX1_LOC_193/Y INVX1_LOC_109/Y 0.04fF
C8160 INVX1_LOC_47/Y INVX1_LOC_26/Y 0.62fF
C8161 NAND2X1_LOC_192/A INVX1_LOC_168/Y 0.16fF
C8162 INVX1_LOC_63/Y NAND2X1_LOC_845/B 0.01fF
C8163 INVX1_LOC_513/A INVX1_LOC_479/A 0.13fF
C8164 INVX1_LOC_120/Y INVX1_LOC_242/Y 0.03fF
C8165 INVX1_LOC_555/A INVX1_LOC_475/Y 0.01fF
C8166 INVX1_LOC_500/A INVX1_LOC_58/Y 0.57fF
C8167 INVX1_LOC_63/Y INVX1_LOC_491/A 0.14fF
C8168 INVX1_LOC_130/Y INVX1_LOC_92/A 0.02fF
C8169 INVX1_LOC_166/Y INVX1_LOC_338/Y 0.09fF
C8170 NAND2X1_LOC_686/A INVX1_LOC_114/A 0.00fF
C8171 INVX1_LOC_62/Y INVX1_LOC_497/A 0.03fF
C8172 VDD INVX1_LOC_447/A -0.00fF
C8173 INVX1_LOC_62/Y INVX1_LOC_338/Y 0.10fF
C8174 NAND2X1_LOC_45/Y NAND2X1_LOC_249/Y 0.07fF
C8175 INVX1_LOC_6/Y NAND2X1_LOC_234/Y 0.00fF
C8176 INVX1_LOC_224/Y INVX1_LOC_301/A 0.03fF
C8177 INVX1_LOC_26/Y INVX1_LOC_119/Y 0.11fF
C8178 INVX1_LOC_26/Y NAND2X1_LOC_66/Y 0.03fF
C8179 INVX1_LOC_119/Y INVX1_LOC_128/Y 0.36fF
C8180 INVX1_LOC_508/A INVX1_LOC_645/Y 0.00fF
C8181 INVX1_LOC_301/A INVX1_LOC_578/A 0.03fF
C8182 INPUT_0 INVX1_LOC_594/Y 0.10fF
C8183 INVX1_LOC_58/Y INVX1_LOC_634/Y 0.07fF
C8184 INVX1_LOC_76/Y INVX1_LOC_275/A 0.01fF
C8185 INVX1_LOC_79/A INVX1_LOC_274/Y 0.00fF
C8186 NAND2X1_LOC_516/Y INVX1_LOC_121/Y 0.04fF
C8187 NAND2X1_LOC_88/B NAND2X1_LOC_86/Y 0.05fF
C8188 VDD INVX1_LOC_163/Y 0.05fF
C8189 NAND2X1_LOC_322/Y NAND2X1_LOC_322/a_36_24# 0.02fF
C8190 INVX1_LOC_438/A INVX1_LOC_76/Y 0.07fF
C8191 INVX1_LOC_206/Y NAND2X1_LOC_332/B 0.03fF
C8192 INVX1_LOC_134/Y INVX1_LOC_638/A 0.01fF
C8193 VDD INVX1_LOC_522/Y 1.81fF
C8194 NAND2X1_LOC_704/a_36_24# INVX1_LOC_510/Y 0.00fF
C8195 INVX1_LOC_20/Y INVX1_LOC_224/Y 0.41fF
C8196 VDD NAND2X1_LOC_20/Y -0.00fF
C8197 VDD INVX1_LOC_489/A -0.00fF
C8198 INVX1_LOC_21/Y NAND2X1_LOC_543/B 0.11fF
C8199 INVX1_LOC_20/Y INVX1_LOC_578/A 0.14fF
C8200 NAND2X1_LOC_45/Y INVX1_LOC_369/A 0.03fF
C8201 NAND2X1_LOC_249/Y INVX1_LOC_99/Y 0.28fF
C8202 INVX1_LOC_617/Y INVX1_LOC_546/Y 0.03fF
C8203 NAND2X1_LOC_87/a_36_24# INVX1_LOC_395/A 0.00fF
C8204 NAND2X1_LOC_48/a_36_24# INVX1_LOC_206/Y 0.00fF
C8205 INVX1_LOC_291/A INVX1_LOC_45/Y 0.12fF
C8206 INVX1_LOC_438/A INVX1_LOC_386/Y 0.14fF
C8207 INVX1_LOC_402/Y INVX1_LOC_553/Y 0.28fF
C8208 VDD NAND2X1_LOC_606/Y 0.05fF
C8209 INVX1_LOC_118/Y NAND2X1_LOC_595/Y 0.01fF
C8210 NAND2X1_LOC_750/Y NAND2X1_LOC_266/a_36_24# 0.00fF
C8211 INVX1_LOC_224/Y INVX1_LOC_300/A 0.16fF
C8212 VDD INVX1_LOC_411/A -0.00fF
C8213 INVX1_LOC_224/Y INVX1_LOC_197/Y 0.03fF
C8214 INVX1_LOC_17/Y NAND2X1_LOC_537/B -0.02fF
C8215 INVX1_LOC_374/A INVX1_LOC_188/Y 0.03fF
C8216 INVX1_LOC_655/Y INVX1_LOC_651/Y 0.08fF
C8217 NAND2X1_LOC_467/A INVX1_LOC_147/Y 0.07fF
C8218 VDD INVX1_LOC_295/Y 0.01fF
C8219 INVX1_LOC_560/A INVX1_LOC_99/Y 0.08fF
C8220 NAND2X1_LOC_231/A INVX1_LOC_80/A 0.00fF
C8221 NAND2X1_LOC_43/a_36_24# INVX1_LOC_31/Y 0.01fF
C8222 NAND2X1_LOC_780/B INVX1_LOC_186/Y 0.02fF
C8223 INVX1_LOC_447/A INVX1_LOC_103/Y 0.00fF
C8224 INVX1_LOC_45/Y INVX1_LOC_531/A 0.01fF
C8225 INVX1_LOC_578/A INVX1_LOC_197/Y 0.00fF
C8226 INVX1_LOC_76/Y NAND2X1_LOC_513/A 0.03fF
C8227 NAND2X1_LOC_152/Y INVX1_LOC_53/Y 0.14fF
C8228 INVX1_LOC_607/Y NAND2X1_LOC_142/Y 0.17fF
C8229 INVX1_LOC_11/Y INVX1_LOC_215/Y 0.02fF
C8230 INVX1_LOC_374/A NAND2X1_LOC_645/a_36_24# 0.00fF
C8231 INVX1_LOC_677/Y INVX1_LOC_632/A 0.00fF
C8232 INVX1_LOC_412/Y INVX1_LOC_93/Y 0.03fF
C8233 INVX1_LOC_614/A INVX1_LOC_522/Y 0.30fF
C8234 INVX1_LOC_45/Y INVX1_LOC_357/A 0.00fF
C8235 INVX1_LOC_384/A NAND2X1_LOC_478/a_36_24# 0.02fF
C8236 INVX1_LOC_17/Y INVX1_LOC_586/A 0.18fF
C8237 INVX1_LOC_301/A INVX1_LOC_120/Y 0.00fF
C8238 NAND2X1_LOC_20/Y INVX1_LOC_42/A 0.09fF
C8239 INVX1_LOC_552/Y NAND2X1_LOC_387/Y 0.01fF
C8240 INVX1_LOC_45/Y NAND2X1_LOC_837/B 0.01fF
C8241 INVX1_LOC_158/A NAND2X1_LOC_388/A 0.01fF
C8242 VDD INVX1_LOC_508/A -0.00fF
C8243 NAND2X1_LOC_317/A INVX1_LOC_89/Y 0.06fF
C8244 INVX1_LOC_150/Y INVX1_LOC_335/A 0.11fF
C8245 INVX1_LOC_373/A INVX1_LOC_496/Y 0.15fF
C8246 INVX1_LOC_425/A INVX1_LOC_418/Y 0.14fF
C8247 NAND2X1_LOC_529/a_36_24# INVX1_LOC_46/Y 0.01fF
C8248 INVX1_LOC_45/Y INVX1_LOC_118/A 0.00fF
C8249 INVX1_LOC_459/A INVX1_LOC_79/A 0.02fF
C8250 NAND2X1_LOC_372/a_36_24# INVX1_LOC_303/Y 0.00fF
C8251 INVX1_LOC_530/Y INVX1_LOC_117/Y 0.01fF
C8252 INVX1_LOC_425/A INVX1_LOC_159/Y 0.03fF
C8253 NAND2X1_LOC_755/B INVX1_LOC_658/A 0.01fF
C8254 INVX1_LOC_312/Y INVX1_LOC_503/A 0.03fF
C8255 INVX1_LOC_412/Y INVX1_LOC_675/A 0.02fF
C8256 NAND2X1_LOC_34/a_36_24# INVX1_LOC_41/Y 0.00fF
C8257 NAND2X1_LOC_507/A INVX1_LOC_266/Y 0.02fF
C8258 NAND2X1_LOC_756/Y INVX1_LOC_35/Y 0.04fF
C8259 INVX1_LOC_277/A INVX1_LOC_651/Y 0.02fF
C8260 NAND2X1_LOC_636/A INVX1_LOC_79/A 0.01fF
C8261 NAND2X1_LOC_177/a_36_24# NAND2X1_LOC_775/B 0.00fF
C8262 INVX1_LOC_335/Y NAND2X1_LOC_638/A 7.18fF
C8263 INVX1_LOC_51/Y INVX1_LOC_260/Y 0.01fF
C8264 INVX1_LOC_683/Y INVX1_LOC_510/A 0.02fF
C8265 INVX1_LOC_369/A INVX1_LOC_99/Y 0.03fF
C8266 INVX1_LOC_165/Y INVX1_LOC_89/Y 0.05fF
C8267 INVX1_LOC_171/Y INVX1_LOC_172/A 0.00fF
C8268 INVX1_LOC_17/Y INVX1_LOC_312/Y 0.42fF
C8269 NAND2X1_LOC_318/A INVX1_LOC_117/Y 0.99fF
C8270 INVX1_LOC_53/Y INVX1_LOC_176/A 0.07fF
C8271 INVX1_LOC_605/A INVX1_LOC_199/Y 0.03fF
C8272 INVX1_LOC_448/A NAND2X1_LOC_478/a_36_24# 0.00fF
C8273 INVX1_LOC_409/Y INVX1_LOC_41/Y 0.03fF
C8274 NAND2X1_LOC_475/A INVX1_LOC_26/Y 0.01fF
C8275 INVX1_LOC_206/Y INVX1_LOC_242/Y 0.14fF
C8276 INVX1_LOC_205/Y INVX1_LOC_274/A 0.01fF
C8277 INVX1_LOC_159/A INVX1_LOC_519/A 0.61fF
C8278 INVX1_LOC_617/Y INVX1_LOC_93/Y 0.07fF
C8279 NAND2X1_LOC_322/Y INVX1_LOC_41/Y 0.06fF
C8280 INVX1_LOC_269/A INVX1_LOC_63/Y 0.08fF
C8281 INVX1_LOC_395/A INVX1_LOC_485/Y 0.01fF
C8282 INVX1_LOC_224/Y NAND2X1_LOC_269/B 0.03fF
C8283 NAND2X1_LOC_727/a_36_24# INVX1_LOC_376/Y 0.00fF
C8284 INVX1_LOC_504/Y INVX1_LOC_506/Y 0.02fF
C8285 INVX1_LOC_46/A INVX1_LOC_46/Y 0.22fF
C8286 INVX1_LOC_160/Y INVX1_LOC_353/A 0.19fF
C8287 INVX1_LOC_439/Y INVX1_LOC_385/Y 0.12fF
C8288 INVX1_LOC_556/Y INVX1_LOC_125/A 0.00fF
C8289 INVX1_LOC_130/Y INPUT_1 0.06fF
C8290 NAND2X1_LOC_399/B INVX1_LOC_50/Y 0.14fF
C8291 NAND2X1_LOC_171/a_36_24# INVX1_LOC_53/Y 0.01fF
C8292 INVX1_LOC_490/A INVX1_LOC_489/Y 0.08fF
C8293 NAND2X1_LOC_308/A INVX1_LOC_134/Y 0.20fF
C8294 INVX1_LOC_50/Y INVX1_LOC_7/Y 0.03fF
C8295 NAND2X1_LOC_673/B INVX1_LOC_35/Y 0.00fF
C8296 INVX1_LOC_519/A INVX1_LOC_66/A 0.03fF
C8297 NAND2X1_LOC_39/Y INVX1_LOC_170/A 0.05fF
C8298 INVX1_LOC_300/A INVX1_LOC_227/Y 0.04fF
C8299 INVX1_LOC_417/A INVX1_LOC_31/Y 0.01fF
C8300 NAND2X1_LOC_850/a_36_24# NAND2X1_LOC_260/Y 0.00fF
C8301 INVX1_LOC_47/Y INVX1_LOC_369/A 0.07fF
C8302 INVX1_LOC_79/A INVX1_LOC_624/A 0.02fF
C8303 INVX1_LOC_412/Y NAND2X1_LOC_62/a_36_24# 0.00fF
C8304 INVX1_LOC_382/A NAND2X1_LOC_415/B 0.01fF
C8305 INVX1_LOC_20/Y NAND2X1_LOC_493/a_36_24# 0.00fF
C8306 NAND2X1_LOC_749/a_36_24# INVX1_LOC_178/A 0.00fF
C8307 INVX1_LOC_194/Y INVX1_LOC_195/Y 0.10fF
C8308 INVX1_LOC_80/A INVX1_LOC_77/Y 0.17fF
C8309 INVX1_LOC_202/Y INVX1_LOC_117/Y 0.03fF
C8310 INVX1_LOC_614/A INVX1_LOC_508/A 0.05fF
C8311 INVX1_LOC_638/Y INVX1_LOC_632/A 0.02fF
C8312 INVX1_LOC_273/A NAND2X1_LOC_262/a_36_24# 0.00fF
C8313 NAND2X1_LOC_24/Y INVX1_LOC_63/Y 0.01fF
C8314 INVX1_LOC_435/Y INVX1_LOC_62/Y 0.04fF
C8315 NAND2X1_LOC_457/A NAND2X1_LOC_458/a_36_24# 0.00fF
C8316 INVX1_LOC_53/Y INVX1_LOC_170/Y 0.01fF
C8317 INVX1_LOC_551/Y INVX1_LOC_245/A 0.11fF
C8318 INVX1_LOC_69/Y INVX1_LOC_232/Y 0.01fF
C8319 INVX1_LOC_666/A INVX1_LOC_100/Y 0.02fF
C8320 INVX1_LOC_649/Y NAND2X1_LOC_846/B 0.18fF
C8321 INVX1_LOC_46/Y INVX1_LOC_251/Y 0.17fF
C8322 INVX1_LOC_448/A NAND2X1_LOC_542/A 0.07fF
C8323 INVX1_LOC_46/Y INVX1_LOC_178/A 0.09fF
C8324 NAND2X1_LOC_669/Y INVX1_LOC_44/Y 0.01fF
C8325 INVX1_LOC_596/A INVX1_LOC_9/Y 0.07fF
C8326 INVX1_LOC_89/Y INVX1_LOC_352/A 0.00fF
C8327 INVX1_LOC_435/Y NAND2X1_LOC_844/A 0.03fF
C8328 INVX1_LOC_261/Y INVX1_LOC_290/A 0.00fF
C8329 INVX1_LOC_68/Y INVX1_LOC_41/Y 0.07fF
C8330 NAND2X1_LOC_493/B INVX1_LOC_319/A 0.02fF
C8331 INVX1_LOC_686/A INVX1_LOC_242/Y 0.04fF
C8332 INVX1_LOC_548/A NAND2X1_LOC_128/A 0.33fF
C8333 INVX1_LOC_345/Y INVX1_LOC_50/Y 0.00fF
C8334 INVX1_LOC_575/A INVX1_LOC_476/A 0.00fF
C8335 INVX1_LOC_110/A INPUT_1 0.03fF
C8336 INVX1_LOC_545/A INVX1_LOC_69/Y 0.01fF
C8337 INVX1_LOC_32/Y INVX1_LOC_50/Y 0.24fF
C8338 INVX1_LOC_548/A NAND2X1_LOC_127/a_36_24# 0.00fF
C8339 INVX1_LOC_624/Y INVX1_LOC_98/Y 0.05fF
C8340 INVX1_LOC_280/Y INVX1_LOC_31/Y 0.01fF
C8341 INVX1_LOC_448/A INVX1_LOC_376/Y 0.10fF
C8342 INVX1_LOC_502/A INVX1_LOC_486/Y 0.01fF
C8343 INVX1_LOC_63/Y INVX1_LOC_504/Y 0.24fF
C8344 INVX1_LOC_117/Y INVX1_LOC_387/Y 0.03fF
C8345 INVX1_LOC_20/Y INVX1_LOC_621/A 0.21fF
C8346 INVX1_LOC_366/Y INVX1_LOC_9/Y 0.01fF
C8347 INVX1_LOC_79/A INVX1_LOC_635/A 0.05fF
C8348 NAND2X1_LOC_833/B NAND2X1_LOC_253/a_36_24# 0.00fF
C8349 INVX1_LOC_596/A INVX1_LOC_62/Y 0.02fF
C8350 NAND2X1_LOC_299/Y NAND2X1_LOC_123/B 0.01fF
C8351 INVX1_LOC_399/A NAND2X1_LOC_226/Y 0.01fF
C8352 INVX1_LOC_209/A INVX1_LOC_44/Y 0.04fF
C8353 NAND2X1_LOC_56/Y INVX1_LOC_531/Y 0.00fF
C8354 INVX1_LOC_54/Y INVX1_LOC_199/Y 0.12fF
C8355 INVX1_LOC_17/Y INVX1_LOC_225/Y 0.01fF
C8356 NAND2X1_LOC_325/B INVX1_LOC_100/Y 0.07fF
C8357 NAND2X1_LOC_558/B INVX1_LOC_230/A 0.02fF
C8358 NAND2X1_LOC_192/A INVX1_LOC_137/Y 0.02fF
C8359 NAND2X1_LOC_273/a_36_24# INVX1_LOC_74/Y 0.00fF
C8360 INVX1_LOC_431/A NAND2X1_LOC_615/Y 0.02fF
C8361 INVX1_LOC_100/Y NAND2X1_LOC_72/Y 0.12fF
C8362 INVX1_LOC_117/Y INVX1_LOC_49/Y 0.24fF
C8363 INVX1_LOC_25/Y INVX1_LOC_26/Y 0.01fF
C8364 INVX1_LOC_99/Y NAND2X1_LOC_626/Y 0.01fF
C8365 INVX1_LOC_41/Y INVX1_LOC_600/A 0.07fF
C8366 NAND2X1_LOC_130/Y INVX1_LOC_41/Y 0.00fF
C8367 INVX1_LOC_128/A INVX1_LOC_510/A 0.02fF
C8368 INVX1_LOC_366/A INVX1_LOC_623/A 0.01fF
C8369 INVX1_LOC_555/A NAND2X1_LOC_611/a_36_24# 0.00fF
C8370 NAND2X1_LOC_509/a_36_24# INVX1_LOC_63/Y 0.00fF
C8371 INVX1_LOC_58/Y INVX1_LOC_46/Y 2.51fF
C8372 INVX1_LOC_79/A INVX1_LOC_230/A 0.00fF
C8373 INVX1_LOC_244/Y INVX1_LOC_453/Y 0.08fF
C8374 INVX1_LOC_41/Y INVX1_LOC_64/A 0.01fF
C8375 INPUT_3 INVX1_LOC_488/Y 0.02fF
C8376 INVX1_LOC_257/A INVX1_LOC_199/Y 0.19fF
C8377 NAND2X1_LOC_673/A INVX1_LOC_100/Y 0.01fF
C8378 INVX1_LOC_383/Y INVX1_LOC_666/Y 0.11fF
C8379 INVX1_LOC_74/Y NAND2X1_LOC_72/Y 0.20fF
C8380 NAND2X1_LOC_267/A INVX1_LOC_353/A 0.98fF
C8381 NAND2X1_LOC_331/Y INVX1_LOC_495/Y 0.14fF
C8382 NAND2X1_LOC_274/Y INVX1_LOC_420/A 0.01fF
C8383 INVX1_LOC_595/Y NAND2X1_LOC_409/Y 0.02fF
C8384 NAND2X1_LOC_376/B INVX1_LOC_183/A 0.02fF
C8385 INVX1_LOC_53/Y INVX1_LOC_611/A 0.06fF
C8386 INVX1_LOC_93/Y NAND2X1_LOC_268/a_36_24# 0.01fF
C8387 INVX1_LOC_376/A NAND2X1_LOC_437/a_36_24# 0.00fF
C8388 INVX1_LOC_86/Y INVX1_LOC_190/A 0.03fF
C8389 INVX1_LOC_47/Y NAND2X1_LOC_626/Y 0.02fF
C8390 NAND2X1_LOC_707/B INVX1_LOC_588/A 0.02fF
C8391 NAND2X1_LOC_7/Y INVX1_LOC_206/Y 0.01fF
C8392 NAND2X1_LOC_708/A INVX1_LOC_613/A 0.01fF
C8393 INVX1_LOC_301/A INVX1_LOC_206/Y 0.08fF
C8394 INVX1_LOC_644/Y INVX1_LOC_655/A 0.04fF
C8395 INVX1_LOC_74/Y INVX1_LOC_351/Y 0.01fF
C8396 INVX1_LOC_6/Y NAND2X1_LOC_255/a_36_24# 0.00fF
C8397 VDD INVX1_LOC_540/Y 0.29fF
C8398 NAND2X1_LOC_847/A NAND2X1_LOC_843/B 0.19fF
C8399 INVX1_LOC_45/Y INVX1_LOC_220/A 0.33fF
C8400 NAND2X1_LOC_274/B INVX1_LOC_665/A 0.01fF
C8401 NAND2X1_LOC_66/Y NAND2X1_LOC_626/Y 0.01fF
C8402 NAND2X1_LOC_455/a_36_24# INVX1_LOC_211/A 0.01fF
C8403 INVX1_LOC_6/Y INVX1_LOC_623/A 0.01fF
C8404 NAND2X1_LOC_838/a_36_24# INVX1_LOC_658/Y -0.00fF
C8405 VDD INVX1_LOC_271/A 0.00fF
C8406 VDD NAND2X1_LOC_690/Y 0.01fF
C8407 INVX1_LOC_371/Y INVX1_LOC_109/Y 0.00fF
C8408 VDD INVX1_LOC_173/A 0.00fF
C8409 INVX1_LOC_114/A INVX1_LOC_588/A 0.02fF
C8410 VDD INVX1_LOC_322/Y 0.21fF
C8411 INVX1_LOC_546/Y INVX1_LOC_375/A 0.01fF
C8412 INVX1_LOC_347/A NAND2X1_LOC_439/a_36_24# 0.01fF
C8413 INVX1_LOC_65/Y NAND2X1_LOC_100/a_36_24# 0.00fF
C8414 INVX1_LOC_301/A INVX1_LOC_686/A 1.89fF
C8415 NAND2X1_LOC_45/Y INVX1_LOC_235/Y 0.10fF
C8416 NAND2X1_LOC_67/a_36_24# INVX1_LOC_17/Y 0.00fF
C8417 INVX1_LOC_20/Y INVX1_LOC_206/Y 0.39fF
C8418 INVX1_LOC_394/Y INVX1_LOC_274/A 0.03fF
C8419 INVX1_LOC_449/A NAND2X1_LOC_575/a_36_24# 0.02fF
C8420 INVX1_LOC_68/Y INVX1_LOC_160/Y 0.33fF
C8421 VDD NAND2X1_LOC_496/Y 0.02fF
C8422 INVX1_LOC_617/Y INVX1_LOC_395/A 0.10fF
C8423 NAND2X1_LOC_134/a_36_24# NAND2X1_LOC_332/B -0.00fF
C8424 INVX1_LOC_89/Y INVX1_LOC_109/Y 0.03fF
C8425 INVX1_LOC_117/Y INVX1_LOC_297/Y 0.03fF
C8426 INVX1_LOC_594/Y INVX1_LOC_677/A 0.02fF
C8427 VDD NAND2X1_LOC_415/B 0.01fF
C8428 INVX1_LOC_257/Y NAND2X1_LOC_603/Y 0.04fF
C8429 INVX1_LOC_438/A INVX1_LOC_7/Y 0.07fF
C8430 INVX1_LOC_75/Y INVX1_LOC_92/A 0.28fF
C8431 INVX1_LOC_32/Y INVX1_LOC_275/A 0.16fF
C8432 INVX1_LOC_578/A NAND2X1_LOC_524/a_36_24# 0.00fF
C8433 NAND2X1_LOC_390/a_36_24# INVX1_LOC_270/A 0.00fF
C8434 INVX1_LOC_206/Y INVX1_LOC_300/A 0.11fF
C8435 VDD NAND2X1_LOC_775/B 0.07fF
C8436 INVX1_LOC_20/Y INVX1_LOC_242/A 0.03fF
C8437 INVX1_LOC_578/A NAND2X1_LOC_298/a_36_24# 0.00fF
C8438 NAND2X1_LOC_271/B NAND2X1_LOC_270/a_36_24# 0.02fF
C8439 INVX1_LOC_401/Y INVX1_LOC_51/Y 0.12fF
C8440 INVX1_LOC_442/A INVX1_LOC_519/A 0.00fF
C8441 INVX1_LOC_206/Y INVX1_LOC_197/Y 0.07fF
C8442 INVX1_LOC_549/A INVX1_LOC_491/Y 0.09fF
C8443 INVX1_LOC_147/A INVX1_LOC_584/Y 0.02fF
C8444 INVX1_LOC_364/Y INVX1_LOC_134/Y 0.01fF
C8445 NAND2X1_LOC_520/a_36_24# NAND2X1_LOC_271/B 0.01fF
C8446 VDD NAND2X1_LOC_706/B 0.02fF
C8447 INVX1_LOC_255/Y INVX1_LOC_469/A 0.01fF
C8448 INVX1_LOC_554/A INVX1_LOC_89/Y 0.03fF
C8449 NAND2X1_LOC_335/B NAND2X1_LOC_267/A 0.02fF
C8450 NAND2X1_LOC_475/A INVX1_LOC_603/A 0.05fF
C8451 INVX1_LOC_20/Y INVX1_LOC_686/A 0.56fF
C8452 NAND2X1_LOC_636/B INVX1_LOC_76/Y 0.07fF
C8453 NAND2X1_LOC_503/B INVX1_LOC_69/Y 0.01fF
C8454 INVX1_LOC_6/Y INVX1_LOC_388/Y 0.03fF
C8455 NAND2X1_LOC_142/Y INVX1_LOC_145/Y 0.01fF
C8456 NAND2X1_LOC_516/Y INVX1_LOC_251/A 0.01fF
C8457 INVX1_LOC_68/Y INVX1_LOC_21/Y 0.03fF
C8458 INVX1_LOC_438/A INVX1_LOC_32/Y 0.07fF
C8459 INVX1_LOC_374/A INVX1_LOC_504/Y 0.01fF
C8460 INVX1_LOC_34/Y INVX1_LOC_6/A 0.01fF
C8461 NAND2X1_LOC_764/Y INVX1_LOC_117/Y 0.16fF
C8462 NAND2X1_LOC_342/a_36_24# INVX1_LOC_80/A 0.00fF
C8463 NAND2X1_LOC_179/Y INVX1_LOC_51/Y 0.02fF
C8464 INVX1_LOC_570/A INVX1_LOC_556/Y 0.06fF
C8465 NAND2X1_LOC_108/Y NAND2X1_LOC_106/B 0.01fF
C8466 INVX1_LOC_412/Y INVX1_LOC_31/Y 0.45fF
C8467 INVX1_LOC_21/Y INVX1_LOC_88/Y 0.01fF
C8468 NAND2X1_LOC_475/A NAND2X1_LOC_309/a_36_24# 0.00fF
C8469 INVX1_LOC_545/A INVX1_LOC_586/A 0.01fF
C8470 INVX1_LOC_361/Y INVX1_LOC_412/A 0.98fF
C8471 INVX1_LOC_448/Y INVX1_LOC_49/Y 0.05fF
C8472 INVX1_LOC_587/A INVX1_LOC_17/Y 0.00fF
C8473 INVX1_LOC_93/Y INVX1_LOC_410/Y 1.59fF
C8474 INVX1_LOC_654/A NAND2X1_LOC_260/Y 0.00fF
C8475 INVX1_LOC_122/Y INVX1_LOC_47/Y 0.03fF
C8476 INVX1_LOC_51/Y INVX1_LOC_440/Y 0.47fF
C8477 INVX1_LOC_280/Y INVX1_LOC_51/Y 0.10fF
C8478 INVX1_LOC_245/A INVX1_LOC_596/Y 0.03fF
C8479 NAND2X1_LOC_318/A NAND2X1_LOC_76/A 0.00fF
C8480 INVX1_LOC_295/A INVX1_LOC_145/Y 0.05fF
C8481 INVX1_LOC_9/Y NAND2X1_LOC_76/B 0.53fF
C8482 INVX1_LOC_17/Y INVX1_LOC_486/Y 0.03fF
C8483 INVX1_LOC_68/Y NAND2X1_LOC_267/A 0.05fF
C8484 INVX1_LOC_214/Y INVX1_LOC_293/Y 0.02fF
C8485 INVX1_LOC_278/A INVX1_LOC_63/Y 0.03fF
C8486 NAND2X1_LOC_331/A INVX1_LOC_338/Y 0.07fF
C8487 INVX1_LOC_21/Y INVX1_LOC_600/A 0.00fF
C8488 INVX1_LOC_117/Y INVX1_LOC_76/Y 0.84fF
C8489 INVX1_LOC_586/A INVX1_LOC_230/Y 0.03fF
C8490 INVX1_LOC_366/A INVX1_LOC_601/Y 0.01fF
C8491 INVX1_LOC_635/A INVX1_LOC_59/Y 0.00fF
C8492 INVX1_LOC_21/Y NAND2X1_LOC_369/a_36_24# 0.01fF
C8493 INVX1_LOC_398/Y NAND2X1_LOC_237/Y 0.01fF
C8494 NAND2X1_LOC_106/Y NAND2X1_LOC_486/B 0.00fF
C8495 NAND2X1_LOC_122/Y INVX1_LOC_69/Y 0.07fF
C8496 NAND2X1_LOC_616/Y NAND2X1_LOC_202/a_36_24# 0.00fF
C8497 INVX1_LOC_273/A INVX1_LOC_69/Y 0.02fF
C8498 INVX1_LOC_530/Y INVX1_LOC_58/Y 0.16fF
C8499 INVX1_LOC_439/A INVX1_LOC_385/A 0.00fF
C8500 NAND2X1_LOC_332/B NAND2X1_LOC_542/A 0.02fF
C8501 INVX1_LOC_45/Y NAND2X1_LOC_686/B 0.01fF
C8502 INVX1_LOC_122/Y INVX1_LOC_119/Y 0.01fF
C8503 INVX1_LOC_366/Y INVX1_LOC_42/Y 0.00fF
C8504 NAND2X1_LOC_510/a_36_24# INVX1_LOC_600/A 0.00fF
C8505 NAND2X1_LOC_336/B INVX1_LOC_361/Y 0.29fF
C8506 INVX1_LOC_390/Y INVX1_LOC_242/Y 0.01fF
C8507 INVX1_LOC_185/Y INVX1_LOC_507/Y 0.03fF
C8508 INVX1_LOC_54/Y INVX1_LOC_53/Y 7.26fF
C8509 INVX1_LOC_492/A INVX1_LOC_567/Y 0.02fF
C8510 INVX1_LOC_126/Y INVX1_LOC_199/A -0.00fF
C8511 INVX1_LOC_272/Y INVX1_LOC_601/Y 0.00fF
C8512 INVX1_LOC_292/A INVX1_LOC_79/A 0.01fF
C8513 NAND2X1_LOC_673/B INVX1_LOC_531/A 0.00fF
C8514 INVX1_LOC_187/A INVX1_LOC_32/Y 0.32fF
C8515 INVX1_LOC_282/A NAND2X1_LOC_260/Y 0.59fF
C8516 INVX1_LOC_266/Y INVX1_LOC_44/Y 0.09fF
C8517 INVX1_LOC_312/Y INVX1_LOC_230/Y 0.91fF
C8518 NAND2X1_LOC_318/A INVX1_LOC_58/Y 0.06fF
C8519 INVX1_LOC_370/Y INVX1_LOC_665/Y 0.02fF
C8520 INVX1_LOC_407/Y INVX1_LOC_98/Y 0.02fF
C8521 INVX1_LOC_53/Y INVX1_LOC_611/Y 0.01fF
C8522 INVX1_LOC_20/Y NAND2X1_LOC_334/A 0.05fF
C8523 INVX1_LOC_352/Y INVX1_LOC_252/Y 0.10fF
C8524 INVX1_LOC_7/Y INVX1_LOC_327/Y 0.05fF
C8525 INVX1_LOC_202/Y NAND2X1_LOC_76/A 0.03fF
C8526 INVX1_LOC_53/Y INVX1_LOC_257/A 0.07fF
C8527 NAND2X1_LOC_318/B INVX1_LOC_87/A 0.05fF
C8528 INVX1_LOC_48/Y INVX1_LOC_230/A 0.08fF
C8529 INVX1_LOC_649/Y INVX1_LOC_199/Y 0.00fF
C8530 INVX1_LOC_49/Y INVX1_LOC_658/A 0.01fF
C8531 NAND2X1_LOC_152/Y INVX1_LOC_662/A 0.04fF
C8532 INVX1_LOC_287/Y INVX1_LOC_245/A 0.03fF
C8533 INVX1_LOC_655/A INVX1_LOC_242/A 0.09fF
C8534 INVX1_LOC_270/A INVX1_LOC_245/A 0.00fF
C8535 INVX1_LOC_188/Y INVX1_LOC_496/A 0.09fF
C8536 NAND2X1_LOC_320/Y INVX1_LOC_89/Y 0.03fF
C8537 INVX1_LOC_84/A NAND2X1_LOC_845/B 0.02fF
C8538 INVX1_LOC_197/A INVX1_LOC_196/Y 0.15fF
C8539 INVX1_LOC_617/Y INVX1_LOC_128/A 0.01fF
C8540 INVX1_LOC_312/A INVX1_LOC_328/Y 0.01fF
C8541 INVX1_LOC_662/Y INVX1_LOC_283/A 0.03fF
C8542 INVX1_LOC_17/Y INVX1_LOC_6/Y 0.31fF
C8543 NAND2X1_LOC_652/a_36_24# INVX1_LOC_50/Y 0.00fF
C8544 INPUT_5 INVX1_LOC_29/Y 0.47fF
C8545 INVX1_LOC_43/A INVX1_LOC_54/Y 0.01fF
C8546 INVX1_LOC_556/Y INVX1_LOC_568/A -0.00fF
C8547 NAND2X1_LOC_307/A INVX1_LOC_557/Y 0.01fF
C8548 INVX1_LOC_145/Y INVX1_LOC_139/Y 0.02fF
C8549 INVX1_LOC_669/Y INVX1_LOC_646/Y 0.00fF
C8550 INPUT_0 INVX1_LOC_462/Y 0.12fF
C8551 NAND2X1_LOC_398/a_36_24# INVX1_LOC_63/Y 0.00fF
C8552 INVX1_LOC_300/A NAND2X1_LOC_334/A 0.02fF
C8553 INVX1_LOC_117/Y INVX1_LOC_108/A 0.01fF
C8554 INVX1_LOC_80/A NAND2X1_LOC_274/B 0.07fF
C8555 NAND2X1_LOC_403/A INVX1_LOC_63/Y 0.01fF
C8556 INVX1_LOC_169/A NAND2X1_LOC_488/Y 0.01fF
C8557 INVX1_LOC_49/Y INVX1_LOC_178/A 0.07fF
C8558 INVX1_LOC_419/A INVX1_LOC_159/Y 0.03fF
C8559 NAND2X1_LOC_517/Y INVX1_LOC_502/A 0.18fF
C8560 INVX1_LOC_6/Y INVX1_LOC_650/Y 0.01fF
C8561 INVX1_LOC_63/Y INVX1_LOC_453/Y 0.04fF
C8562 INVX1_LOC_202/Y INVX1_LOC_58/Y 0.16fF
C8563 INVX1_LOC_339/Y NAND2X1_LOC_415/B 0.16fF
C8564 NAND2X1_LOC_638/A INVX1_LOC_26/Y 0.05fF
C8565 INVX1_LOC_387/Y INVX1_LOC_608/A 0.23fF
C8566 INVX1_LOC_204/Y INVX1_LOC_623/Y 0.03fF
C8567 INVX1_LOC_99/Y NAND2X1_LOC_420/Y 0.19fF
C8568 INVX1_LOC_625/A INVX1_LOC_9/Y 0.06fF
C8569 INVX1_LOC_575/Y INVX1_LOC_476/A 1.13fF
C8570 NAND2X1_LOC_388/A INVX1_LOC_32/Y 0.03fF
C8571 INVX1_LOC_642/Y INVX1_LOC_178/A 0.02fF
C8572 NAND2X1_LOC_231/A INVX1_LOC_91/Y 0.00fF
C8573 INVX1_LOC_578/Y INVX1_LOC_532/Y 0.01fF
C8574 INVX1_LOC_6/Y INVX1_LOC_601/Y 0.01fF
C8575 INVX1_LOC_99/A INVX1_LOC_100/Y 0.05fF
C8576 INVX1_LOC_211/Y INVX1_LOC_245/A 1.77fF
C8577 INVX1_LOC_681/A INVX1_LOC_79/A 0.00fF
C8578 NAND2X1_LOC_307/B INVX1_LOC_6/Y 0.16fF
C8579 INVX1_LOC_506/Y INVX1_LOC_114/A 0.15fF
C8580 INVX1_LOC_89/Y INVX1_LOC_199/Y 1.55fF
C8581 INVX1_LOC_11/Y NAND2X1_LOC_274/B 0.07fF
C8582 INVX1_LOC_674/A NAND2X1_LOC_334/B 0.01fF
C8583 INVX1_LOC_242/Y INVX1_LOC_432/A 0.01fF
C8584 INVX1_LOC_387/Y INVX1_LOC_58/Y 0.03fF
C8585 NAND2X1_LOC_646/A INVX1_LOC_114/A 0.04fF
C8586 INVX1_LOC_520/A INVX1_LOC_9/Y 0.00fF
C8587 INVX1_LOC_402/Y INVX1_LOC_479/A 0.03fF
C8588 INVX1_LOC_671/A INVX1_LOC_664/Y 0.15fF
C8589 INVX1_LOC_386/A NAND2X1_LOC_252/Y 0.05fF
C8590 INVX1_LOC_63/Y INVX1_LOC_204/Y 0.01fF
C8591 INVX1_LOC_46/Y INVX1_LOC_245/A 0.13fF
C8592 INVX1_LOC_435/A NAND2X1_LOC_528/Y 0.02fF
C8593 INVX1_LOC_49/Y INVX1_LOC_58/Y 2.61fF
C8594 INVX1_LOC_656/A INVX1_LOC_657/A 0.07fF
C8595 INVX1_LOC_380/A VDD 0.00fF
C8596 INVX1_LOC_137/Y INVX1_LOC_74/Y 0.00fF
C8597 VDD INVX1_LOC_627/A -0.00fF
C8598 INVX1_LOC_642/Y INVX1_LOC_58/Y 0.01fF
C8599 INVX1_LOC_681/Y INVX1_LOC_75/Y 0.09fF
C8600 VDD INVX1_LOC_133/Y 0.21fF
C8601 INVX1_LOC_75/Y INPUT_1 0.07fF
C8602 INVX1_LOC_491/A INVX1_LOC_496/A 0.20fF
C8603 NAND2X1_LOC_136/Y NAND2X1_LOC_284/A 0.02fF
C8604 INVX1_LOC_355/Y INVX1_LOC_74/Y 0.00fF
C8605 INVX1_LOC_63/Y INVX1_LOC_114/A 3.71fF
C8606 VDD INVX1_LOC_239/Y 0.24fF
C8607 VDD NAND2X1_LOC_759/B 0.01fF
C8608 INVX1_LOC_242/Y INVX1_LOC_376/Y 0.01fF
C8609 INVX1_LOC_519/Y INVX1_LOC_9/Y 0.03fF
C8610 INVX1_LOC_492/A INVX1_LOC_92/A 0.05fF
C8611 INVX1_LOC_206/Y NAND2X1_LOC_373/Y 0.04fF
C8612 VDD INVX1_LOC_307/Y 0.21fF
C8613 INVX1_LOC_199/Y NAND2X1_LOC_544/B 0.03fF
C8614 INVX1_LOC_58/Y INVX1_LOC_92/Y 0.00fF
C8615 VDD NAND2X1_LOC_271/B 0.02fF
C8616 NAND2X1_LOC_543/B INVX1_LOC_560/A 0.03fF
C8617 VDD NAND2X1_LOC_317/B 0.01fF
C8618 INVX1_LOC_498/A INVX1_LOC_462/Y 0.08fF
C8619 VDD INVX1_LOC_97/A -0.00fF
C8620 INVX1_LOC_409/Y INVX1_LOC_255/Y 0.05fF
C8621 NAND2X1_LOC_573/a_36_24# NAND2X1_LOC_457/A 0.00fF
C8622 INVX1_LOC_438/Y INVX1_LOC_445/A 0.03fF
C8623 INVX1_LOC_622/Y INVX1_LOC_621/Y 0.05fF
C8624 INVX1_LOC_75/A INVX1_LOC_245/A 0.01fF
C8625 INVX1_LOC_395/A INVX1_LOC_553/Y 0.00fF
C8626 NAND2X1_LOC_637/A NAND2X1_LOC_122/Y 0.24fF
C8627 INVX1_LOC_447/A INVX1_LOC_45/Y 0.03fF
C8628 INVX1_LOC_395/A INVX1_LOC_410/Y 0.03fF
C8629 VDD INVX1_LOC_630/Y 0.14fF
C8630 INVX1_LOC_395/A INVX1_LOC_375/A 0.05fF
C8631 VDD NAND2X1_LOC_613/Y 0.01fF
C8632 INVX1_LOC_614/A INVX1_LOC_133/Y 0.00fF
C8633 INVX1_LOC_395/A INVX1_LOC_546/A 0.01fF
C8634 INVX1_LOC_617/A NAND2X1_LOC_249/Y 0.03fF
C8635 INVX1_LOC_412/Y INVX1_LOC_51/Y 0.65fF
C8636 INVX1_LOC_602/A NAND2X1_LOC_770/A 0.01fF
C8637 VDD INVX1_LOC_169/A 0.00fF
C8638 NAND2X1_LOC_475/A NAND2X1_LOC_491/a_36_24# 0.00fF
C8639 INVX1_LOC_510/Y NAND2X1_LOC_317/B 0.01fF
C8640 NAND2X1_LOC_373/Y INVX1_LOC_686/A 0.04fF
C8641 VDD INVX1_LOC_337/Y 0.43fF
C8642 VDD INVX1_LOC_495/A -0.00fF
C8643 NAND2X1_LOC_13/a_36_24# NAND2X1_LOC_475/A 0.01fF
C8644 INVX1_LOC_266/A INVX1_LOC_412/Y 0.03fF
C8645 INVX1_LOC_301/A NAND2X1_LOC_542/a_36_24# 0.01fF
C8646 VDD INVX1_LOC_633/Y 0.46fF
C8647 INVX1_LOC_117/Y INVX1_LOC_192/A 0.05fF
C8648 INVX1_LOC_410/Y INVX1_LOC_683/Y 0.02fF
C8649 INVX1_LOC_586/A NAND2X1_LOC_682/a_36_24# 0.01fF
C8650 INVX1_LOC_185/Y INVX1_LOC_522/Y 0.06fF
C8651 NAND2X1_LOC_770/A INVX1_LOC_117/Y 0.08fF
C8652 NAND2X1_LOC_790/B INVX1_LOC_153/A 0.01fF
C8653 NAND2X1_LOC_572/a_36_24# INVX1_LOC_51/Y 0.00fF
C8654 INPUT_0 INVX1_LOC_379/A 0.07fF
C8655 NAND2X1_LOC_69/B INVX1_LOC_100/A 0.14fF
C8656 INPUT_0 INVX1_LOC_35/Y 0.06fF
C8657 INVX1_LOC_607/A INVX1_LOC_679/Y 0.05fF
C8658 INPUT_0 INVX1_LOC_304/A 0.03fF
C8659 NAND2X1_LOC_526/Y INVX1_LOC_145/Y 0.08fF
C8660 VDD INVX1_LOC_317/A 0.00fF
C8661 NAND2X1_LOC_520/B NAND2X1_LOC_275/Y 0.03fF
C8662 INPUT_0 NAND2X1_LOC_634/a_36_24# 0.00fF
C8663 NAND2X1_LOC_597/a_36_24# INVX1_LOC_513/A 0.00fF
C8664 NAND2X1_LOC_24/Y INVX1_LOC_84/A 0.00fF
C8665 INVX1_LOC_590/Y INVX1_LOC_35/Y 0.01fF
C8666 INVX1_LOC_301/A NAND2X1_LOC_542/A 0.02fF
C8667 INVX1_LOC_118/Y INVX1_LOC_105/Y 0.34fF
C8668 INVX1_LOC_312/A NAND2X1_LOC_381/a_36_24# 0.02fF
C8669 INVX1_LOC_197/Y INVX1_LOC_94/A 0.07fF
C8670 INVX1_LOC_515/A NAND2X1_LOC_679/B 0.22fF
C8671 INVX1_LOC_410/Y INVX1_LOC_31/Y 0.00fF
C8672 INVX1_LOC_614/A INVX1_LOC_581/A 0.03fF
C8673 INVX1_LOC_510/Y NAND2X1_LOC_308/a_36_24# 0.00fF
C8674 INVX1_LOC_76/Y NAND2X1_LOC_76/A 0.02fF
C8675 INVX1_LOC_53/Y NAND2X1_LOC_677/Y 0.33fF
C8676 INVX1_LOC_366/A INVX1_LOC_198/A 1.77fF
C8677 INVX1_LOC_370/Y INVX1_LOC_134/Y 0.02fF
C8678 INVX1_LOC_80/Y INVX1_LOC_600/Y 0.00fF
C8679 NAND2X1_LOC_231/A NAND2X1_LOC_333/B 0.07fF
C8680 INVX1_LOC_20/Y INVX1_LOC_432/A 0.03fF
C8681 INVX1_LOC_395/A INVX1_LOC_646/Y 0.03fF
C8682 INVX1_LOC_455/Y INVX1_LOC_316/Y 0.15fF
C8683 INVX1_LOC_522/A NAND2X1_LOC_654/a_36_24# 0.01fF
C8684 INVX1_LOC_435/A INVX1_LOC_12/Y 0.07fF
C8685 INVX1_LOC_556/Y INVX1_LOC_136/Y 0.18fF
C8686 INVX1_LOC_547/Y INVX1_LOC_63/Y 0.03fF
C8687 INVX1_LOC_418/Y INVX1_LOC_80/A 0.01fF
C8688 INVX1_LOC_185/Y INVX1_LOC_508/A 0.02fF
C8689 INVX1_LOC_117/Y INVX1_LOC_12/A 0.01fF
C8690 INVX1_LOC_340/Y INVX1_LOC_638/Y 0.08fF
C8691 NAND2X1_LOC_418/Y INVX1_LOC_352/A 0.02fF
C8692 INVX1_LOC_406/Y INVX1_LOC_31/Y 0.01fF
C8693 INVX1_LOC_97/A NAND2X1_LOC_786/B 0.17fF
C8694 INVX1_LOC_59/Y NAND2X1_LOC_72/Y 0.01fF
C8695 INVX1_LOC_98/A INVX1_LOC_58/Y 0.02fF
C8696 INVX1_LOC_41/Y NAND2X1_LOC_75/a_36_24# 0.01fF
C8697 INPUT_0 INVX1_LOC_518/Y 0.01fF
C8698 INVX1_LOC_486/Y INVX1_LOC_230/Y 0.05fF
C8699 INVX1_LOC_607/Y INVX1_LOC_35/Y 0.11fF
C8700 INVX1_LOC_20/Y NAND2X1_LOC_542/A 0.03fF
C8701 NAND2X1_LOC_635/B INVX1_LOC_677/A 0.00fF
C8702 INVX1_LOC_76/Y INVX1_LOC_58/Y 0.15fF
C8703 INVX1_LOC_65/Y INVX1_LOC_9/Y 0.46fF
C8704 INVX1_LOC_298/Y INVX1_LOC_678/A 0.01fF
C8705 INVX1_LOC_63/Y INVX1_LOC_378/A 0.03fF
C8706 INVX1_LOC_300/A INVX1_LOC_432/A 0.00fF
C8707 INVX1_LOC_32/Y INVX1_LOC_104/Y 0.02fF
C8708 INVX1_LOC_374/A INVX1_LOC_114/A 0.26fF
C8709 INVX1_LOC_53/Y INVX1_LOC_89/Y 4.07fF
C8710 INPUT_0 INVX1_LOC_79/Y 0.02fF
C8711 INVX1_LOC_117/Y INVX1_LOC_7/Y 0.26fF
C8712 INVX1_LOC_681/A INVX1_LOC_48/Y 0.00fF
C8713 INVX1_LOC_254/Y INVX1_LOC_400/A 0.02fF
C8714 INVX1_LOC_11/Y INVX1_LOC_159/Y 0.13fF
C8715 INVX1_LOC_69/Y INVX1_LOC_519/A 0.02fF
C8716 NAND2X1_LOC_673/A INVX1_LOC_48/Y 0.02fF
C8717 NAND2X1_LOC_165/a_36_24# NAND2X1_LOC_165/Y 0.02fF
C8718 NAND2X1_LOC_318/A INVX1_LOC_245/A 0.06fF
C8719 INVX1_LOC_268/Y INVX1_LOC_245/A 0.02fF
C8720 NAND2X1_LOC_775/B INVX1_LOC_105/A 0.03fF
C8721 INVX1_LOC_282/A INVX1_LOC_663/Y 0.01fF
C8722 INVX1_LOC_492/A INPUT_1 0.03fF
C8723 INVX1_LOC_285/A INVX1_LOC_44/Y 0.02fF
C8724 INVX1_LOC_298/A INVX1_LOC_35/Y 0.04fF
C8725 INVX1_LOC_565/A INVX1_LOC_47/Y 0.01fF
C8726 NAND2X1_LOC_119/a_36_24# INVX1_LOC_509/A 0.00fF
C8727 NAND2X1_LOC_108/Y NAND2X1_LOC_248/B 0.07fF
C8728 INVX1_LOC_65/Y INVX1_LOC_62/Y 0.01fF
C8729 INVX1_LOC_53/Y INVX1_LOC_501/A 0.03fF
C8730 INVX1_LOC_166/A INVX1_LOC_371/A 0.00fF
C8731 INVX1_LOC_297/A INVX1_LOC_328/Y 0.03fF
C8732 NAND2X1_LOC_849/a_36_24# INVX1_LOC_371/A 0.01fF
C8733 INVX1_LOC_117/Y INVX1_LOC_345/Y 0.03fF
C8734 NAND2X1_LOC_27/Y INVX1_LOC_46/Y 0.01fF
C8735 INVX1_LOC_527/Y NAND2X1_LOC_448/B 0.12fF
C8736 INVX1_LOC_254/Y INVX1_LOC_93/Y 0.01fF
C8737 INVX1_LOC_47/Y NAND2X1_LOC_307/a_36_24# 0.01fF
C8738 NAND2X1_LOC_184/Y INVX1_LOC_50/Y 0.17fF
C8739 INVX1_LOC_31/Y INVX1_LOC_674/A 0.07fF
C8740 INVX1_LOC_555/A NAND2X1_LOC_708/A 0.17fF
C8741 INVX1_LOC_207/A NAND2X1_LOC_234/Y 0.00fF
C8742 NAND2X1_LOC_679/B INVX1_LOC_168/Y 0.00fF
C8743 INVX1_LOC_117/Y INVX1_LOC_32/Y 0.78fF
C8744 INVX1_LOC_59/Y INVX1_LOC_351/Y 0.03fF
C8745 INVX1_LOC_224/Y INVX1_LOC_92/A 0.07fF
C8746 INVX1_LOC_469/Y INVX1_LOC_355/Y 0.03fF
C8747 INVX1_LOC_6/Y INVX1_LOC_198/A 0.01fF
C8748 INVX1_LOC_199/Y INVX1_LOC_194/Y 0.10fF
C8749 INVX1_LOC_127/Y INVX1_LOC_670/A 0.02fF
C8750 INVX1_LOC_366/A INVX1_LOC_598/Y 0.00fF
C8751 NAND2X1_LOC_605/B INVX1_LOC_469/A 0.01fF
C8752 INVX1_LOC_26/Y INVX1_LOC_600/A 0.26fF
C8753 NAND2X1_LOC_333/A INVX1_LOC_267/A 0.06fF
C8754 INVX1_LOC_284/A INVX1_LOC_273/Y 0.17fF
C8755 INVX1_LOC_592/Y INVX1_LOC_93/Y 0.09fF
C8756 INVX1_LOC_578/A INVX1_LOC_92/A 0.08fF
C8757 INVX1_LOC_202/Y INVX1_LOC_245/A 0.03fF
C8758 INVX1_LOC_21/Y INVX1_LOC_369/Y 0.45fF
C8759 INVX1_LOC_168/Y INVX1_LOC_48/Y 0.09fF
C8760 INVX1_LOC_367/A INVX1_LOC_479/A 0.42fF
C8761 NAND2X1_LOC_274/B INVX1_LOC_367/Y 0.03fF
C8762 INVX1_LOC_523/Y GATE_662 0.09fF
C8763 INVX1_LOC_272/Y INVX1_LOC_598/Y 0.00fF
C8764 INVX1_LOC_520/Y INVX1_LOC_46/Y 0.02fF
C8765 NAND2X1_LOC_307/a_36_24# INVX1_LOC_119/Y 0.00fF
C8766 INVX1_LOC_430/A INVX1_LOC_453/Y 0.52fF
C8767 INVX1_LOC_53/Y NAND2X1_LOC_544/B 0.01fF
C8768 NAND2X1_LOC_308/A INVX1_LOC_338/Y 0.35fF
C8769 INVX1_LOC_137/Y INVX1_LOC_79/A 0.04fF
C8770 INVX1_LOC_204/Y NAND2X1_LOC_836/B 0.39fF
C8771 INVX1_LOC_419/Y INVX1_LOC_100/Y 0.07fF
C8772 INVX1_LOC_349/A NAND2X1_LOC_545/A 0.00fF
C8773 INVX1_LOC_69/Y INVX1_LOC_659/A 0.21fF
C8774 NAND2X1_LOC_165/Y INVX1_LOC_90/Y 0.04fF
C8775 INVX1_LOC_454/Y INVX1_LOC_259/Y 0.02fF
C8776 INVX1_LOC_479/A INVX1_LOC_669/Y 0.02fF
C8777 NAND2X1_LOC_274/B INVX1_LOC_374/Y 0.01fF
C8778 INVX1_LOC_44/Y INVX1_LOC_199/Y 0.09fF
C8779 INVX1_LOC_79/A INVX1_LOC_355/Y 0.00fF
C8780 NAND2X1_LOC_441/a_36_24# INPUT_1 0.00fF
C8781 INVX1_LOC_400/A INVX1_LOC_479/A 0.02fF
C8782 INVX1_LOC_118/Y INVX1_LOC_109/Y 0.03fF
C8783 INVX1_LOC_35/Y INVX1_LOC_211/A 0.10fF
C8784 INVX1_LOC_49/Y INVX1_LOC_245/A 0.06fF
C8785 INVX1_LOC_75/Y INVX1_LOC_50/Y 0.07fF
C8786 INVX1_LOC_119/Y NAND2X1_LOC_586/Y 0.03fF
C8787 NAND2X1_LOC_846/A INVX1_LOC_667/A 0.09fF
C8788 INVX1_LOC_93/Y INVX1_LOC_479/A 0.67fF
C8789 INVX1_LOC_568/Y INVX1_LOC_92/A 0.02fF
C8790 NAND2X1_LOC_281/a_36_24# NAND2X1_LOC_248/B 0.00fF
C8791 INVX1_LOC_17/Y INVX1_LOC_636/A 0.07fF
C8792 INVX1_LOC_226/Y INVX1_LOC_224/A 0.19fF
C8793 INVX1_LOC_446/A NAND2X1_LOC_457/A 0.17fF
C8794 INVX1_LOC_468/Y INVX1_LOC_92/A 0.12fF
C8795 INVX1_LOC_82/Y INVX1_LOC_81/A 0.00fF
C8796 NAND2X1_LOC_69/B INVX1_LOC_308/Y 0.01fF
C8797 INVX1_LOC_6/Y INVX1_LOC_598/Y 0.00fF
C8798 INVX1_LOC_217/A INVX1_LOC_217/Y 0.04fF
C8799 INVX1_LOC_376/A INVX1_LOC_74/Y 0.02fF
C8800 INVX1_LOC_92/Y INVX1_LOC_245/A 0.04fF
C8801 INVX1_LOC_62/Y NAND2X1_LOC_633/a_36_24# 0.00fF
C8802 NAND2X1_LOC_391/A INVX1_LOC_109/Y 0.03fF
C8803 VDD INVX1_LOC_317/Y 0.24fF
C8804 INVX1_LOC_150/A INVX1_LOC_586/A 0.17fF
C8805 INVX1_LOC_166/Y INVX1_LOC_588/A 0.02fF
C8806 INVX1_LOC_540/Y INVX1_LOC_45/Y 0.01fF
C8807 INVX1_LOC_553/Y INVX1_LOC_51/Y 0.10fF
C8808 INVX1_LOC_62/Y INVX1_LOC_588/A 0.19fF
C8809 INVX1_LOC_20/Y INVX1_LOC_121/Y 0.20fF
C8810 INVX1_LOC_375/A NAND2X1_LOC_794/a_36_24# 0.00fF
C8811 NAND2X1_LOC_231/B INVX1_LOC_203/A 0.05fF
C8812 INVX1_LOC_271/A INVX1_LOC_45/Y 0.39fF
C8813 VDD INVX1_LOC_249/A -0.00fF
C8814 INVX1_LOC_173/A INVX1_LOC_45/Y 0.01fF
C8815 INVX1_LOC_409/A INVX1_LOC_80/A 0.01fF
C8816 NAND2X1_LOC_780/B INVX1_LOC_53/Y 0.06fF
C8817 NAND2X1_LOC_843/B NAND2X1_LOC_245/a_36_24# 0.00fF
C8818 VDD INVX1_LOC_106/A -0.00fF
C8819 INVX1_LOC_68/Y NAND2X1_LOC_97/a_36_24# 0.00fF
C8820 INVX1_LOC_20/Y NAND2X1_LOC_142/Y 0.02fF
C8821 NAND2X1_LOC_13/Y INVX1_LOC_321/A 0.01fF
C8822 INVX1_LOC_449/Y VDD 0.17fF
C8823 INVX1_LOC_20/Y NAND2X1_LOC_845/a_36_24# 0.00fF
C8824 INVX1_LOC_53/Y INVX1_LOC_137/A 0.21fF
C8825 INPUT_0 INVX1_LOC_338/A 0.00fF
C8826 NAND2X1_LOC_321/a_36_24# INVX1_LOC_374/A 0.00fF
C8827 VDD INVX1_LOC_588/Y 0.32fF
C8828 NAND2X1_LOC_554/a_36_24# NAND2X1_LOC_706/B -0.01fF
C8829 INVX1_LOC_21/Y INVX1_LOC_428/A 0.00fF
C8830 INVX1_LOC_547/Y NAND2X1_LOC_499/a_36_24# 0.00fF
C8831 INVX1_LOC_586/A INVX1_LOC_519/A 0.01fF
C8832 INVX1_LOC_45/Y NAND2X1_LOC_496/Y 0.01fF
C8833 INVX1_LOC_448/Y INVX1_LOC_32/Y 0.01fF
C8834 INVX1_LOC_224/Y INVX1_LOC_681/Y 0.02fF
C8835 NAND2X1_LOC_267/A NAND2X1_LOC_75/a_36_24# 0.01fF
C8836 INVX1_LOC_224/Y INPUT_1 0.07fF
C8837 INVX1_LOC_433/Y NAND2X1_LOC_294/Y 0.11fF
C8838 VDD INVX1_LOC_239/A 0.01fF
C8839 INVX1_LOC_20/Y NAND2X1_LOC_603/Y 0.16fF
C8840 INVX1_LOC_72/Y NAND2X1_LOC_378/Y 0.02fF
C8841 INVX1_LOC_245/A INVX1_LOC_297/Y 1.24fF
C8842 INVX1_LOC_578/A INVX1_LOC_681/Y 0.00fF
C8843 VDD NAND2X1_LOC_111/Y 0.04fF
C8844 INVX1_LOC_206/Y NAND2X1_LOC_106/Y 0.07fF
C8845 INVX1_LOC_20/Y INVX1_LOC_296/Y 0.07fF
C8846 INVX1_LOC_312/Y INVX1_LOC_519/A 0.03fF
C8847 INVX1_LOC_578/A INPUT_1 0.38fF
C8848 INVX1_LOC_246/Y NAND2X1_LOC_296/Y 0.00fF
C8849 INVX1_LOC_434/A NAND2X1_LOC_344/B 2.49fF
C8850 INVX1_LOC_384/A INVX1_LOC_35/Y 0.07fF
C8851 INVX1_LOC_51/Y INVX1_LOC_61/A 0.04fF
C8852 INPUT_3 NAND2X1_LOC_397/Y 0.00fF
C8853 INVX1_LOC_85/Y INVX1_LOC_195/Y 0.21fF
C8854 INPUT_3 NAND2X1_LOC_415/B 0.35fF
C8855 NAND2X1_LOC_706/B INVX1_LOC_45/Y 0.59fF
C8856 INVX1_LOC_409/Y NAND2X1_LOC_605/B 0.05fF
C8857 INVX1_LOC_592/Y INVX1_LOC_395/A 0.02fF
C8858 NAND2X1_LOC_45/Y INVX1_LOC_183/A 0.13fF
C8859 INVX1_LOC_137/Y INVX1_LOC_610/Y 0.01fF
C8860 INVX1_LOC_184/A INVX1_LOC_42/Y 0.03fF
C8861 INVX1_LOC_166/A INVX1_LOC_510/Y 1.40fF
C8862 INVX1_LOC_139/A INVX1_LOC_58/Y 0.00fF
C8863 VDD INVX1_LOC_153/Y 0.29fF
C8864 INVX1_LOC_417/Y INVX1_LOC_99/A 0.00fF
C8865 INVX1_LOC_134/Y INVX1_LOC_98/Y 0.12fF
C8866 VDD NAND2X1_LOC_136/Y 0.02fF
C8867 INVX1_LOC_395/A INVX1_LOC_309/Y 0.03fF
C8868 INVX1_LOC_360/Y INVX1_LOC_633/Y 0.06fF
C8869 INVX1_LOC_596/A INVX1_LOC_665/Y 0.03fF
C8870 INVX1_LOC_80/A INVX1_LOC_352/Y 0.01fF
C8871 INVX1_LOC_296/Y INVX1_LOC_300/A 0.02fF
C8872 INVX1_LOC_28/Y NAND2X1_LOC_84/B 0.03fF
C8873 NAND2X1_LOC_383/Y INVX1_LOC_89/Y 0.02fF
C8874 INVX1_LOC_400/A INVX1_LOC_12/Y 0.07fF
C8875 INVX1_LOC_448/A INVX1_LOC_35/Y 0.19fF
C8876 INVX1_LOC_414/Y INVX1_LOC_63/Y 0.10fF
C8877 VDD INVX1_LOC_531/Y 2.64fF
C8878 INVX1_LOC_35/Y NAND2X1_LOC_612/A 0.01fF
C8879 INVX1_LOC_167/A INVX1_LOC_197/A 0.02fF
C8880 NAND2X1_LOC_516/B INVX1_LOC_66/A 0.01fF
C8881 INVX1_LOC_80/A INVX1_LOC_345/A 0.00fF
C8882 INVX1_LOC_7/Y INVX1_LOC_178/A 0.05fF
C8883 INVX1_LOC_393/Y NAND2X1_LOC_274/B 0.00fF
C8884 INVX1_LOC_352/A INVX1_LOC_252/Y 0.00fF
C8885 INVX1_LOC_228/A INVX1_LOC_178/A 0.03fF
C8886 INVX1_LOC_137/Y NAND2X1_LOC_679/B 0.96fF
C8887 INVX1_LOC_11/Y NAND2X1_LOC_595/Y 0.03fF
C8888 INVX1_LOC_35/Y INVX1_LOC_145/Y 0.49fF
C8889 INVX1_LOC_612/Y INVX1_LOC_609/Y 0.01fF
C8890 NAND2X1_LOC_335/a_36_24# INVX1_LOC_9/Y 0.00fF
C8891 INVX1_LOC_420/Y INVX1_LOC_41/Y 0.03fF
C8892 VDD INVX1_LOC_528/Y 0.21fF
C8893 INVX1_LOC_93/Y INVX1_LOC_12/Y 0.07fF
C8894 INVX1_LOC_228/Y INVX1_LOC_531/Y 0.04fF
C8895 NAND2X1_LOC_796/a_36_24# INVX1_LOC_54/Y 0.00fF
C8896 NAND2X1_LOC_142/Y INVX1_LOC_655/A 0.04fF
C8897 INVX1_LOC_51/A INVX1_LOC_41/Y 0.00fF
C8898 INVX1_LOC_484/A INVX1_LOC_369/A 0.02fF
C8899 INVX1_LOC_438/A INVX1_LOC_75/Y 0.03fF
C8900 NAND2X1_LOC_147/B NAND2X1_LOC_148/B 0.02fF
C8901 INVX1_LOC_11/Y INVX1_LOC_352/Y 0.03fF
C8902 INVX1_LOC_468/Y INPUT_1 0.03fF
C8903 INPUT_4 NAND2X1_LOC_64/a_36_24# 0.00fF
C8904 INVX1_LOC_32/Y INVX1_LOC_281/Y 0.03fF
C8905 INVX1_LOC_76/Y INVX1_LOC_245/A 0.06fF
C8906 NAND2X1_LOC_191/a_36_24# INVX1_LOC_99/Y 0.00fF
C8907 INVX1_LOC_395/A NAND2X1_LOC_528/Y 0.16fF
C8908 NAND2X1_LOC_542/A INVX1_LOC_375/Y 0.03fF
C8909 INVX1_LOC_206/Y NAND2X1_LOC_428/Y 0.02fF
C8910 INVX1_LOC_372/Y INVX1_LOC_675/A 0.02fF
C8911 VDD INVX1_LOC_363/A -0.00fF
C8912 NAND2X1_LOC_45/Y INVX1_LOC_109/A 0.02fF
C8913 INVX1_LOC_134/Y INVX1_LOC_338/Y 0.10fF
C8914 INVX1_LOC_395/A INVX1_LOC_479/A 1.86fF
C8915 INVX1_LOC_402/Y INVX1_LOC_66/A 0.93fF
C8916 INVX1_LOC_166/A INVX1_LOC_509/A 0.02fF
C8917 INVX1_LOC_206/Y NAND2X1_LOC_263/a_36_24# 0.01fF
C8918 INVX1_LOC_298/A NAND2X1_LOC_837/B 0.02fF
C8919 INVX1_LOC_53/Y INVX1_LOC_44/Y 3.81fF
C8920 INVX1_LOC_145/Y INVX1_LOC_620/A 0.00fF
C8921 NAND2X1_LOC_755/B NAND2X1_LOC_753/Y 0.04fF
C8922 VDD INVX1_LOC_613/A 0.20fF
C8923 INVX1_LOC_237/Y NAND2X1_LOC_843/B 0.01fF
C8924 INVX1_LOC_145/Y NAND2X1_LOC_253/Y 0.73fF
C8925 INVX1_LOC_17/Y NAND2X1_LOC_200/a_36_24# 0.00fF
C8926 INVX1_LOC_32/Y NAND2X1_LOC_76/A 0.08fF
C8927 INVX1_LOC_206/Y INVX1_LOC_270/Y 0.06fF
C8928 INVX1_LOC_276/A NAND2X1_LOC_342/B 0.01fF
C8929 INVX1_LOC_662/A INVX1_LOC_649/Y 0.05fF
C8930 INVX1_LOC_392/A NAND2X1_LOC_521/Y 0.17fF
C8931 INPUT_0 INVX1_LOC_488/Y 0.00fF
C8932 NAND2X1_LOC_260/Y INVX1_LOC_654/Y 0.01fF
C8933 NAND2X1_LOC_106/Y NAND2X1_LOC_706/a_36_24# 0.00fF
C8934 INVX1_LOC_376/Y INVX1_LOC_375/Y 0.26fF
C8935 INVX1_LOC_175/A INVX1_LOC_100/Y 0.04fF
C8936 INVX1_LOC_254/Y INVX1_LOC_31/Y 0.03fF
C8937 INVX1_LOC_58/Y INVX1_LOC_7/Y 0.00fF
C8938 INVX1_LOC_297/A INVX1_LOC_224/A 0.00fF
C8939 INVX1_LOC_438/A NAND2X1_LOC_271/A 0.00fF
C8940 INVX1_LOC_318/Y INVX1_LOC_90/Y 0.01fF
C8941 INVX1_LOC_435/A INVX1_LOC_296/A 0.08fF
C8942 INVX1_LOC_47/Y INVX1_LOC_304/Y 0.03fF
C8943 INVX1_LOC_670/Y INVX1_LOC_9/Y 0.31fF
C8944 INVX1_LOC_65/A INVX1_LOC_98/Y 0.46fF
C8945 INVX1_LOC_145/Y INVX1_LOC_621/Y 0.01fF
C8946 NAND2X1_LOC_307/A INVX1_LOC_79/A 0.05fF
C8947 INVX1_LOC_206/Y INVX1_LOC_92/A 0.10fF
C8948 INVX1_LOC_671/A INVX1_LOC_671/Y 0.21fF
C8949 INVX1_LOC_545/Y INVX1_LOC_79/A 0.00fF
C8950 INVX1_LOC_686/A NAND2X1_LOC_123/B 0.02fF
C8951 INVX1_LOC_321/Y INVX1_LOC_482/Y 0.01fF
C8952 NAND2X1_LOC_333/A INVX1_LOC_93/Y 0.03fF
C8953 INVX1_LOC_367/A INVX1_LOC_680/A -0.02fF
C8954 INVX1_LOC_8/Y INVX1_LOC_63/Y 0.05fF
C8955 INVX1_LOC_32/Y INVX1_LOC_157/A 0.00fF
C8956 NAND2X1_LOC_111/Y INVX1_LOC_103/Y 0.11fF
C8957 INVX1_LOC_449/A INVX1_LOC_665/A 0.04fF
C8958 INVX1_LOC_80/A INVX1_LOC_203/A 0.01fF
C8959 INVX1_LOC_80/A NAND2X1_LOC_372/Y 0.03fF
C8960 INVX1_LOC_32/Y INVX1_LOC_58/Y 0.12fF
C8961 NAND2X1_LOC_835/A INVX1_LOC_659/A 0.02fF
C8962 INVX1_LOC_523/Y INVX1_LOC_199/Y 0.87fF
C8963 INVX1_LOC_17/Y INVX1_LOC_100/Y 0.20fF
C8964 NAND2X1_LOC_301/B INVX1_LOC_440/Y 0.42fF
C8965 NAND2X1_LOC_433/Y INVX1_LOC_345/A 0.05fF
C8966 NAND2X1_LOC_137/A NAND2X1_LOC_768/B 0.17fF
C8967 INVX1_LOC_361/Y NAND2X1_LOC_274/B 0.61fF
C8968 NAND2X1_LOC_814/Y NAND2X1_LOC_846/B 0.16fF
C8969 INVX1_LOC_17/Y INVX1_LOC_74/Y 0.21fF
C8970 INVX1_LOC_54/Y NAND2X1_LOC_545/A 0.10fF
C8971 NAND2X1_LOC_286/A INVX1_LOC_58/Y 0.01fF
C8972 INVX1_LOC_41/Y INVX1_LOC_371/A 0.00fF
C8973 INVX1_LOC_183/A INVX1_LOC_47/Y 0.14fF
C8974 INVX1_LOC_298/A INVX1_LOC_657/A 0.04fF
C8975 INVX1_LOC_11/Y NAND2X1_LOC_372/Y 0.00fF
C8976 INVX1_LOC_548/A INVX1_LOC_479/A 0.02fF
C8977 INVX1_LOC_62/Y NAND2X1_LOC_646/A 0.02fF
C8978 INVX1_LOC_686/A INVX1_LOC_92/A 0.01fF
C8979 INVX1_LOC_285/Y INVX1_LOC_63/Y 0.01fF
C8980 INVX1_LOC_477/Y INVX1_LOC_655/A 0.02fF
C8981 INVX1_LOC_54/Y INVX1_LOC_653/Y 0.08fF
C8982 INVX1_LOC_63/Y INVX1_LOC_9/Y 0.71fF
C8983 INVX1_LOC_531/Y INVX1_LOC_68/A 0.06fF
C8984 INVX1_LOC_588/Y INVX1_LOC_635/Y 0.03fF
C8985 INVX1_LOC_328/Y NAND2X1_LOC_236/a_36_24# 0.00fF
C8986 INVX1_LOC_451/A NAND2X1_LOC_416/B 0.04fF
C8987 NAND2X1_LOC_647/A INVX1_LOC_614/Y 0.13fF
C8988 INVX1_LOC_31/Y INVX1_LOC_479/A 0.05fF
C8989 INVX1_LOC_376/A INVX1_LOC_79/A 0.60fF
C8990 INVX1_LOC_183/Y INVX1_LOC_26/Y 0.34fF
C8991 INVX1_LOC_618/A INVX1_LOC_375/A 0.01fF
C8992 NAND2X1_LOC_420/Y INVX1_LOC_353/A 0.11fF
C8993 INVX1_LOC_351/A INVX1_LOC_90/Y 0.01fF
C8994 INVX1_LOC_425/A INVX1_LOC_109/Y 0.05fF
C8995 INVX1_LOC_241/A INVX1_LOC_66/A 0.01fF
C8996 NAND2X1_LOC_843/B INVX1_LOC_212/Y 0.05fF
C8997 INVX1_LOC_103/Y INVX1_LOC_363/A 0.01fF
C8998 INVX1_LOC_50/Y NAND2X1_LOC_98/B 0.23fF
C8999 INVX1_LOC_63/Y INVX1_LOC_62/Y 2.31fF
C9000 INVX1_LOC_204/A INVX1_LOC_273/Y 0.01fF
C9001 INVX1_LOC_369/Y INVX1_LOC_26/Y 0.46fF
C9002 INVX1_LOC_121/Y INVX1_LOC_553/A 0.02fF
C9003 INVX1_LOC_68/Y NAND2X1_LOC_790/B 0.08fF
C9004 INPUT_6 INVX1_LOC_33/A 0.13fF
C9005 NAND2X1_LOC_457/A NAND2X1_LOC_368/a_36_24# 0.02fF
C9006 VDD INVX1_LOC_302/A -0.00fF
C9007 NAND2X1_LOC_480/a_36_24# INVX1_LOC_443/A 0.05fF
C9008 VDD INVX1_LOC_580/A -0.00fF
C9009 INVX1_LOC_44/Y NAND2X1_LOC_60/Y 0.06fF
C9010 NAND2X1_LOC_271/B INVX1_LOC_45/Y 0.11fF
C9011 INVX1_LOC_41/Y INVX1_LOC_441/A 0.00fF
C9012 VDD NAND2X1_LOC_467/A 0.17fF
C9013 INVX1_LOC_190/Y INVX1_LOC_366/A 0.05fF
C9014 NAND2X1_LOC_208/a_36_24# INVX1_LOC_190/Y 0.00fF
C9015 INVX1_LOC_578/A INVX1_LOC_134/A 0.05fF
C9016 NAND2X1_LOC_13/Y INVX1_LOC_410/Y 0.03fF
C9017 INVX1_LOC_257/Y INVX1_LOC_256/Y 0.06fF
C9018 NAND2X1_LOC_385/a_36_24# INVX1_LOC_600/A 0.01fF
C9019 NAND2X1_LOC_374/a_36_24# NAND2X1_LOC_325/B 0.01fF
C9020 INVX1_LOC_499/Y INVX1_LOC_512/A 0.00fF
C9021 INVX1_LOC_6/Y INVX1_LOC_423/A 0.09fF
C9022 VDD INVX1_LOC_640/A -0.00fF
C9023 INVX1_LOC_206/Y INVX1_LOC_679/Y 0.09fF
C9024 INVX1_LOC_288/A NAND2X1_LOC_120/a_36_24# 0.00fF
C9025 INVX1_LOC_45/Y INVX1_LOC_169/A 0.00fF
C9026 INVX1_LOC_122/Y NAND2X1_LOC_130/Y 0.19fF
C9027 NAND2X1_LOC_750/Y INVX1_LOC_21/Y 0.04fF
C9028 INVX1_LOC_435/Y INVX1_LOC_134/Y 0.10fF
C9029 INVX1_LOC_21/Y INVX1_LOC_51/A 0.03fF
C9030 INVX1_LOC_395/A INVX1_LOC_12/Y 0.14fF
C9031 INVX1_LOC_629/A INVX1_LOC_17/Y 0.01fF
C9032 INVX1_LOC_563/Y NAND2X1_LOC_755/B 0.02fF
C9033 INVX1_LOC_596/A INVX1_LOC_364/Y 0.01fF
C9034 INVX1_LOC_185/Y INVX1_LOC_633/Y 0.03fF
C9035 INVX1_LOC_45/Y INVX1_LOC_633/Y 0.08fF
C9036 NAND2X1_LOC_711/a_36_24# INVX1_LOC_6/Y 0.00fF
C9037 INVX1_LOC_413/Y INVX1_LOC_99/Y 0.22fF
C9038 INVX1_LOC_257/Y INVX1_LOC_360/A 0.01fF
C9039 INVX1_LOC_224/Y INVX1_LOC_50/Y 1.61fF
C9040 INVX1_LOC_409/A INVX1_LOC_374/Y 0.02fF
C9041 INVX1_LOC_206/Y INPUT_1 0.10fF
C9042 INVX1_LOC_454/A INVX1_LOC_340/A 0.27fF
C9043 INVX1_LOC_490/Y INVX1_LOC_54/Y 0.03fF
C9044 INVX1_LOC_662/Y NAND2X1_LOC_108/Y 0.04fF
C9045 INVX1_LOC_412/Y INVX1_LOC_359/A 0.04fF
C9046 NAND2X1_LOC_475/A NAND2X1_LOC_422/a_36_24# 0.00fF
C9047 INVX1_LOC_596/A INVX1_LOC_134/Y 0.07fF
C9048 INVX1_LOC_395/A INVX1_LOC_138/Y 0.01fF
C9049 INVX1_LOC_578/A INVX1_LOC_50/Y 0.07fF
C9050 INVX1_LOC_293/Y NAND2X1_LOC_496/Y 0.08fF
C9051 INVX1_LOC_412/Y NAND2X1_LOC_466/a_36_24# 0.00fF
C9052 INVX1_LOC_206/Y INVX1_LOC_292/Y 1.95fF
C9053 VDD INVX1_LOC_411/Y 0.55fF
C9054 NAND2X1_LOC_332/B INVX1_LOC_35/Y 0.06fF
C9055 NAND2X1_LOC_745/a_36_24# INVX1_LOC_53/Y 0.00fF
C9056 INVX1_LOC_54/Y NAND2X1_LOC_16/Y -0.08fF
C9057 INVX1_LOC_255/Y INVX1_LOC_359/Y 0.01fF
C9058 NAND2X1_LOC_271/B NAND2X1_LOC_276/A 0.02fF
C9059 INVX1_LOC_312/Y NAND2X1_LOC_147/B 0.03fF
C9060 INVX1_LOC_80/A INVX1_LOC_67/Y 0.28fF
C9061 VDD INVX1_LOC_301/Y 0.46fF
C9062 INVX1_LOC_84/A INVX1_LOC_194/A 0.01fF
C9063 INVX1_LOC_45/Y INVX1_LOC_490/A 0.03fF
C9064 INVX1_LOC_125/Y INVX1_LOC_35/Y 0.10fF
C9065 NAND2X1_LOC_710/a_36_24# INVX1_LOC_47/Y 0.01fF
C9066 INVX1_LOC_504/A INVX1_LOC_134/Y 0.07fF
C9067 NAND2X1_LOC_521/Y INVX1_LOC_362/Y 0.01fF
C9068 INPUT_1 INVX1_LOC_242/A 0.00fF
C9069 INVX1_LOC_274/A INVX1_LOC_80/A 0.18fF
C9070 INVX1_LOC_229/Y INVX1_LOC_178/A 0.02fF
C9071 INVX1_LOC_446/A INVX1_LOC_62/Y 0.07fF
C9072 INVX1_LOC_288/Y INVX1_LOC_676/Y 0.00fF
C9073 INVX1_LOC_72/Y INVX1_LOC_6/Y 0.03fF
C9074 INVX1_LOC_192/Y INVX1_LOC_390/A 0.01fF
C9075 INVX1_LOC_54/Y NAND2X1_LOC_783/a_36_24# 0.00fF
C9076 INVX1_LOC_209/A INVX1_LOC_80/A 0.03fF
C9077 INPUT_0 INVX1_LOC_223/Y 0.24fF
C9078 NAND2X1_LOC_460/A INVX1_LOC_35/Y 0.14fF
C9079 INVX1_LOC_531/A INVX1_LOC_145/Y 0.03fF
C9080 INVX1_LOC_385/Y INVX1_LOC_451/Y 0.02fF
C9081 INVX1_LOC_628/A INVX1_LOC_17/Y 0.00fF
C9082 INVX1_LOC_449/A INVX1_LOC_11/Y 0.07fF
C9083 INVX1_LOC_492/A NAND2X1_LOC_513/A 0.03fF
C9084 INVX1_LOC_686/A INPUT_1 0.11fF
C9085 NAND2X1_LOC_307/A INVX1_LOC_48/Y 0.01fF
C9086 INVX1_LOC_412/Y NAND2X1_LOC_301/B 0.03fF
C9087 VDD INVX1_LOC_41/Y 1.68fF
C9088 INVX1_LOC_416/A INVX1_LOC_417/Y 0.03fF
C9089 NAND2X1_LOC_685/A INVX1_LOC_496/Y 0.00fF
C9090 INVX1_LOC_419/Y INVX1_LOC_417/Y 0.41fF
C9091 INVX1_LOC_268/Y NAND2X1_LOC_753/Y 0.02fF
C9092 INVX1_LOC_587/A INVX1_LOC_659/A 0.01fF
C9093 INVX1_LOC_214/Y INVX1_LOC_145/Y 0.03fF
C9094 INVX1_LOC_372/Y INVX1_LOC_31/Y 0.38fF
C9095 INVX1_LOC_160/A NAND2X1_LOC_775/B 0.00fF
C9096 NAND2X1_LOC_710/a_36_24# INVX1_LOC_119/Y 0.00fF
C9097 INVX1_LOC_145/Y NAND2X1_LOC_837/B 0.42fF
C9098 INVX1_LOC_547/A INVX1_LOC_63/Y 0.00fF
C9099 INVX1_LOC_428/A INVX1_LOC_26/Y 0.01fF
C9100 NAND2X1_LOC_596/Y INVX1_LOC_41/Y 0.58fF
C9101 INVX1_LOC_367/A INVX1_LOC_66/A 0.01fF
C9102 INVX1_LOC_12/Y INVX1_LOC_31/Y 5.36fF
C9103 NAND2X1_LOC_720/a_36_24# INVX1_LOC_298/A 0.00fF
C9104 INPUT_1 INVX1_LOC_14/A 0.04fF
C9105 INVX1_LOC_228/Y INVX1_LOC_41/Y 0.01fF
C9106 INVX1_LOC_277/A INVX1_LOC_679/A 0.13fF
C9107 INVX1_LOC_116/Y NAND2X1_LOC_603/a_36_24# 0.00fF
C9108 INVX1_LOC_229/Y INVX1_LOC_58/Y 0.02fF
C9109 INVX1_LOC_400/A NAND2X1_LOC_615/B 0.02fF
C9110 NAND2X1_LOC_416/Y INVX1_LOC_46/Y 0.03fF
C9111 INVX1_LOC_42/Y INVX1_LOC_86/Y 0.09fF
C9112 INVX1_LOC_402/A INVX1_LOC_89/Y 0.03fF
C9113 NAND2X1_LOC_331/A INVX1_LOC_588/A 0.18fF
C9114 INVX1_LOC_17/Y INVX1_LOC_469/Y 0.05fF
C9115 INVX1_LOC_17/Y INVX1_LOC_350/Y -0.00fF
C9116 INVX1_LOC_323/Y INVX1_LOC_6/Y 0.04fF
C9117 INVX1_LOC_337/Y INVX1_LOC_89/A 0.01fF
C9118 NAND2X1_LOC_93/Y NAND2X1_LOC_98/B 0.02fF
C9119 GATE_865 INVX1_LOC_259/Y 0.03fF
C9120 INVX1_LOC_374/A INVX1_LOC_62/Y 0.03fF
C9121 INVX1_LOC_361/Y INVX1_LOC_159/Y 0.07fF
C9122 INVX1_LOC_516/A INVX1_LOC_66/A 0.02fF
C9123 INVX1_LOC_16/Y INVX1_LOC_338/Y 0.07fF
C9124 INVX1_LOC_669/Y INVX1_LOC_66/A 0.00fF
C9125 INVX1_LOC_352/Y INVX1_LOC_374/Y 0.42fF
C9126 INVX1_LOC_17/Y NAND2X1_LOC_181/A 0.02fF
C9127 INVX1_LOC_51/Y NAND2X1_LOC_528/Y 0.00fF
C9128 NAND2X1_LOC_789/A INVX1_LOC_198/A 0.10fF
C9129 INVX1_LOC_444/Y NAND2X1_LOC_531/Y 0.03fF
C9130 INVX1_LOC_166/A INVX1_LOC_105/A 0.01fF
C9131 INVX1_LOC_395/A INVX1_LOC_212/A 0.05fF
C9132 INVX1_LOC_51/Y INVX1_LOC_479/A 0.15fF
C9133 INVX1_LOC_530/Y INVX1_LOC_483/A -0.03fF
C9134 INVX1_LOC_87/A INVX1_LOC_86/Y 0.17fF
C9135 INVX1_LOC_50/Y INVX1_LOC_93/A 0.09fF
C9136 INVX1_LOC_42/Y INVX1_LOC_63/Y 0.00fF
C9137 INVX1_LOC_7/Y INVX1_LOC_245/A 0.06fF
C9138 NAND2X1_LOC_111/Y INVX1_LOC_105/A 0.03fF
C9139 INVX1_LOC_93/Y INVX1_LOC_66/A 0.03fF
C9140 INVX1_LOC_100/Y NAND2X1_LOC_616/Y 0.05fF
C9141 INVX1_LOC_266/A INVX1_LOC_479/A 0.08fF
C9142 INVX1_LOC_376/A INVX1_LOC_48/Y 0.07fF
C9143 INVX1_LOC_336/Y NAND2X1_LOC_410/Y 0.02fF
C9144 INVX1_LOC_11/Y INVX1_LOC_328/Y 0.03fF
C9145 INVX1_LOC_35/Y INVX1_LOC_242/Y 0.11fF
C9146 INVX1_LOC_11/Y INVX1_LOC_518/A 0.07fF
C9147 INVX1_LOC_170/A INVX1_LOC_31/Y 0.08fF
C9148 INVX1_LOC_90/Y INVX1_LOC_98/Y 0.12fF
C9149 INVX1_LOC_17/Y INVX1_LOC_79/A 0.22fF
C9150 INVX1_LOC_6/Y NAND2X1_LOC_846/A 0.17fF
C9151 INVX1_LOC_345/Y NAND2X1_LOC_440/A 0.01fF
C9152 NAND2X1_LOC_814/Y INVX1_LOC_199/Y 0.00fF
C9153 INVX1_LOC_356/Y INVX1_LOC_463/Y 0.01fF
C9154 INVX1_LOC_103/Y INVX1_LOC_301/Y 0.46fF
C9155 INVX1_LOC_41/Y INVX1_LOC_116/A 0.01fF
C9156 INVX1_LOC_17/Y INVX1_LOC_460/A 0.01fF
C9157 INVX1_LOC_49/Y NAND2X1_LOC_753/Y 0.65fF
C9158 INVX1_LOC_367/Y INVX1_LOC_280/A 4.20fF
C9159 INVX1_LOC_371/Y INVX1_LOC_666/Y 0.27fF
C9160 INVX1_LOC_35/Y INVX1_LOC_487/A 0.01fF
C9161 INVX1_LOC_502/A INVX1_LOC_48/Y 0.07fF
C9162 INVX1_LOC_32/Y INVX1_LOC_245/A 0.55fF
C9163 INVX1_LOC_63/Y INVX1_LOC_624/Y 0.01fF
C9164 INVX1_LOC_42/Y NAND2X1_LOC_214/a_36_24# 0.00fF
C9165 INVX1_LOC_145/Y INVX1_LOC_364/A 0.01fF
C9166 NAND2X1_LOC_432/a_36_24# INVX1_LOC_345/A 0.01fF
C9167 INVX1_LOC_274/A NAND2X1_LOC_244/a_36_24# 0.02fF
C9168 INVX1_LOC_361/Y INVX1_LOC_468/A 0.01fF
C9169 INVX1_LOC_103/Y INVX1_LOC_41/Y 0.76fF
C9170 NAND2X1_LOC_157/a_36_24# NAND2X1_LOC_836/B 0.00fF
C9171 INVX1_LOC_485/Y INVX1_LOC_486/A 0.12fF
C9172 INVX1_LOC_74/Y INVX1_LOC_497/Y 0.03fF
C9173 INVX1_LOC_89/Y NAND2X1_LOC_545/A 0.10fF
C9174 INVX1_LOC_444/Y INVX1_LOC_443/A 0.05fF
C9175 INVX1_LOC_117/Y INVX1_LOC_75/Y 0.22fF
C9176 NAND2X1_LOC_186/a_36_24# INVX1_LOC_588/A 0.01fF
C9177 INVX1_LOC_81/A INVX1_LOC_9/Y 0.01fF
C9178 INVX1_LOC_89/Y INVX1_LOC_666/Y 0.07fF
C9179 INVX1_LOC_555/A INVX1_LOC_645/Y 0.00fF
C9180 INVX1_LOC_49/Y INVX1_LOC_652/Y 0.01fF
C9181 NAND2X1_LOC_406/a_36_24# INVX1_LOC_636/A -0.01fF
C9182 INVX1_LOC_9/Y INVX1_LOC_669/A 0.01fF
C9183 INVX1_LOC_224/Y INVX1_LOC_438/A 0.17fF
C9184 INVX1_LOC_41/Y NAND2X1_LOC_786/B 0.10fF
C9185 VDD INVX1_LOC_160/Y 0.21fF
C9186 INVX1_LOC_63/Y NAND2X1_LOC_224/a_36_24# 0.00fF
C9187 INVX1_LOC_438/A INVX1_LOC_578/A 0.05fF
C9188 INVX1_LOC_192/Y INVX1_LOC_395/A 0.00fF
C9189 VDD INVX1_LOC_315/Y 0.31fF
C9190 NAND2X1_LOC_542/A INVX1_LOC_92/A -0.00fF
C9191 INVX1_LOC_604/A INVX1_LOC_395/A 0.01fF
C9192 INVX1_LOC_41/Y INVX1_LOC_635/Y 0.05fF
C9193 INVX1_LOC_328/Y INVX1_LOC_231/Y 0.05fF
C9194 INVX1_LOC_26/Y NAND2X1_LOC_832/A 0.05fF
C9195 INVX1_LOC_206/Y INVX1_LOC_134/A 0.01fF
C9196 INVX1_LOC_434/A INVX1_LOC_384/A 0.07fF
C9197 INVX1_LOC_578/A INVX1_LOC_441/Y 0.01fF
C9198 INVX1_LOC_376/Y INVX1_LOC_92/A 0.07fF
C9199 INPUT_6 INVX1_LOC_333/A 0.01fF
C9200 INVX1_LOC_426/A INVX1_LOC_12/Y 0.19fF
C9201 INVX1_LOC_203/A INVX1_LOC_91/Y 0.01fF
C9202 VDD INVX1_LOC_358/Y 0.57fF
C9203 INVX1_LOC_255/Y NAND2X1_LOC_173/Y 0.01fF
C9204 VDD INVX1_LOC_21/Y 3.35fF
C9205 INVX1_LOC_335/Y VDD 0.54fF
C9206 NAND2X1_LOC_294/Y INVX1_LOC_423/A 0.03fF
C9207 INVX1_LOC_424/A NAND2X1_LOC_416/Y 0.00fF
C9208 INVX1_LOC_301/A INVX1_LOC_35/Y 0.07fF
C9209 NAND2X1_LOC_475/A INVX1_LOC_154/Y 0.00fF
C9210 INVX1_LOC_301/A INVX1_LOC_304/A 0.00fF
C9211 NAND2X1_LOC_173/Y INVX1_LOC_577/Y 0.09fF
C9212 INVX1_LOC_335/Y NAND2X1_LOC_596/Y 0.77fF
C9213 INVX1_LOC_454/A INVX1_LOC_455/A 0.94fF
C9214 INVX1_LOC_48/Y INVX1_LOC_388/Y 0.00fF
C9215 INVX1_LOC_134/A INVX1_LOC_686/A 0.01fF
C9216 INVX1_LOC_290/Y INVX1_LOC_602/Y 0.05fF
C9217 INVX1_LOC_410/Y NAND2X1_LOC_102/a_36_24# 0.00fF
C9218 NAND2X1_LOC_543/B NAND2X1_LOC_444/A 0.03fF
C9219 INVX1_LOC_80/A INVX1_LOC_266/Y 0.04fF
C9220 INVX1_LOC_556/A INVX1_LOC_99/Y 0.07fF
C9221 INVX1_LOC_257/Y INVX1_LOC_350/A 0.01fF
C9222 INVX1_LOC_617/Y INVX1_LOC_551/Y 0.10fF
C9223 INVX1_LOC_11/Y NAND2X1_LOC_317/A 0.18fF
C9224 VDD NAND2X1_LOC_267/A 0.08fF
C9225 INPUT_0 NAND2X1_LOC_606/Y 0.01fF
C9226 NAND2X1_LOC_98/a_36_24# NAND2X1_LOC_333/B 0.00fF
C9227 INVX1_LOC_206/Y INVX1_LOC_50/Y 0.37fF
C9228 INVX1_LOC_54/A INVX1_LOC_54/Y 0.02fF
C9229 NAND2X1_LOC_331/A NAND2X1_LOC_646/A 0.00fF
C9230 INVX1_LOC_238/Y INVX1_LOC_520/A 0.09fF
C9231 INVX1_LOC_21/Y INVX1_LOC_510/Y 0.15fF
C9232 INVX1_LOC_547/A INVX1_LOC_387/A 0.06fF
C9233 INVX1_LOC_11/Y INVX1_LOC_165/Y 0.03fF
C9234 VDD INVX1_LOC_181/Y 0.21fF
C9235 INVX1_LOC_603/Y NAND2X1_LOC_508/a_36_24# 0.01fF
C9236 INVX1_LOC_417/A INVX1_LOC_270/A 0.03fF
C9237 INVX1_LOC_224/Y NAND2X1_LOC_388/A 0.04fF
C9238 VDD INVX1_LOC_107/Y 0.38fF
C9239 INVX1_LOC_286/Y INVX1_LOC_59/Y 0.02fF
C9240 INVX1_LOC_285/A INVX1_LOC_599/Y 0.20fF
C9241 INVX1_LOC_533/Y NAND2X1_LOC_448/B 0.41fF
C9242 INVX1_LOC_395/A INVX1_LOC_66/A 0.16fF
C9243 INVX1_LOC_20/Y INVX1_LOC_35/Y 2.65fF
C9244 INVX1_LOC_442/A INVX1_LOC_93/Y 0.07fF
C9245 INVX1_LOC_166/A INVX1_LOC_45/Y 0.04fF
C9246 INVX1_LOC_197/A INVX1_LOC_115/A 0.15fF
C9247 INVX1_LOC_578/A NAND2X1_LOC_388/A 0.03fF
C9248 INVX1_LOC_26/Y INVX1_LOC_180/Y 0.01fF
C9249 NAND2X1_LOC_673/B INVX1_LOC_169/A 0.00fF
C9250 INVX1_LOC_379/A NAND2X1_LOC_473/a_36_24# 0.01fF
C9251 INVX1_LOC_254/Y NAND2X1_LOC_13/Y 0.03fF
C9252 INVX1_LOC_286/Y INVX1_LOC_48/Y 0.01fF
C9253 INVX1_LOC_395/A INVX1_LOC_296/A 0.01fF
C9254 INVX1_LOC_404/Y INVX1_LOC_63/Y 0.06fF
C9255 INVX1_LOC_416/A NAND2X1_LOC_129/a_36_24# 0.00fF
C9256 NAND2X1_LOC_333/A INVX1_LOC_51/Y 0.05fF
C9257 NAND2X1_LOC_331/A INVX1_LOC_63/Y 0.00fF
C9258 INVX1_LOC_544/A INVX1_LOC_367/A 0.04fF
C9259 INVX1_LOC_80/A INVX1_LOC_352/A 0.01fF
C9260 INVX1_LOC_50/Y INVX1_LOC_242/A 0.03fF
C9261 INVX1_LOC_267/Y NAND2X1_LOC_755/B 0.21fF
C9262 INVX1_LOC_188/Y INVX1_LOC_99/Y 0.03fF
C9263 INVX1_LOC_454/A NAND2X1_LOC_823/Y 0.02fF
C9264 INVX1_LOC_362/Y INVX1_LOC_66/A 0.07fF
C9265 INVX1_LOC_191/A INVX1_LOC_86/Y 0.01fF
C9266 INVX1_LOC_449/A INVX1_LOC_367/Y 0.07fF
C9267 INVX1_LOC_603/Y INVX1_LOC_99/Y 0.03fF
C9268 INVX1_LOC_17/Y INVX1_LOC_632/A 0.07fF
C9269 INVX1_LOC_686/A INVX1_LOC_50/Y 0.07fF
C9270 INVX1_LOC_393/A INVX1_LOC_49/Y 0.04fF
C9271 NAND2X1_LOC_750/Y INVX1_LOC_26/Y 0.00fF
C9272 INVX1_LOC_20/Y NAND2X1_LOC_448/B 0.42fF
C9273 INVX1_LOC_51/Y INVX1_LOC_188/A 0.00fF
C9274 INVX1_LOC_20/Y INVX1_LOC_620/A 0.03fF
C9275 INVX1_LOC_21/Y INVX1_LOC_509/A 0.01fF
C9276 INVX1_LOC_353/Y INVX1_LOC_89/Y 0.01fF
C9277 NAND2X1_LOC_241/B INVX1_LOC_26/Y 0.01fF
C9278 INVX1_LOC_395/A INVX1_LOC_178/Y 0.03fF
C9279 INVX1_LOC_170/A INVX1_LOC_51/Y 0.05fF
C9280 INPUT_4 INVX1_LOC_59/A 0.03fF
C9281 INVX1_LOC_544/A INVX1_LOC_669/Y 0.20fF
C9282 INVX1_LOC_463/A INVX1_LOC_479/A 0.08fF
C9283 NAND2X1_LOC_471/a_36_24# INVX1_LOC_510/A 0.00fF
C9284 INVX1_LOC_397/Y INVX1_LOC_398/A 0.07fF
C9285 INVX1_LOC_17/Y INVX1_LOC_59/Y 0.05fF
C9286 INVX1_LOC_300/A INVX1_LOC_35/Y 0.07fF
C9287 INVX1_LOC_353/Y INVX1_LOC_154/A 0.01fF
C9288 NAND2X1_LOC_39/Y INVX1_LOC_6/Y 0.19fF
C9289 INVX1_LOC_35/Y INVX1_LOC_197/Y 0.03fF
C9290 INVX1_LOC_11/Y INVX1_LOC_352/A 0.00fF
C9291 INVX1_LOC_683/Y INVX1_LOC_66/A 0.03fF
C9292 INVX1_LOC_165/Y NAND2X1_LOC_433/Y 0.19fF
C9293 INVX1_LOC_361/Y INVX1_LOC_377/A 0.00fF
C9294 NAND2X1_LOC_643/a_36_24# INVX1_LOC_510/A 0.00fF
C9295 INVX1_LOC_12/Y INVX1_LOC_254/A 0.00fF
C9296 INVX1_LOC_574/Y INVX1_LOC_6/Y 0.01fF
C9297 INVX1_LOC_406/A NAND2X1_LOC_541/B 0.01fF
C9298 NAND2X1_LOC_370/A INVX1_LOC_100/Y 0.03fF
C9299 INVX1_LOC_614/A INVX1_LOC_555/A 0.08fF
C9300 NAND2X1_LOC_274/B INVX1_LOC_618/Y 0.01fF
C9301 INVX1_LOC_21/Y INVX1_LOC_103/Y 0.28fF
C9302 INVX1_LOC_17/Y INVX1_LOC_48/Y 0.34fF
C9303 INVX1_LOC_603/Y INVX1_LOC_589/Y 0.05fF
C9304 INVX1_LOC_208/Y NAND2X1_LOC_241/a_36_24# 0.00fF
C9305 NAND2X1_LOC_387/Y INVX1_LOC_99/Y 0.13fF
C9306 INVX1_LOC_47/Y INVX1_LOC_188/Y 0.07fF
C9307 INVX1_LOC_197/A INVX1_LOC_49/Y 0.03fF
C9308 NAND2X1_LOC_331/B INVX1_LOC_495/Y 0.09fF
C9309 INVX1_LOC_11/Y INVX1_LOC_172/A 0.02fF
C9310 INVX1_LOC_531/Y NAND2X1_LOC_506/B 0.08fF
C9311 INVX1_LOC_444/Y INVX1_LOC_382/A 0.03fF
C9312 INVX1_LOC_525/Y NAND2X1_LOC_755/B 0.01fF
C9313 INVX1_LOC_300/A NAND2X1_LOC_448/B 0.05fF
C9314 INVX1_LOC_93/Y INVX1_LOC_116/Y 0.10fF
C9315 NAND2X1_LOC_173/Y INVX1_LOC_26/Y 0.06fF
C9316 INVX1_LOC_51/Y INVX1_LOC_680/A 0.01fF
C9317 INVX1_LOC_84/A INVX1_LOC_9/Y 0.17fF
C9318 INVX1_LOC_45/Y INVX1_LOC_531/Y 0.05fF
C9319 NAND2X1_LOC_370/A INVX1_LOC_74/Y 0.03fF
C9320 INVX1_LOC_11/Y INVX1_LOC_105/Y 0.00fF
C9321 INVX1_LOC_206/Y INVX1_LOC_658/Y 0.14fF
C9322 INVX1_LOC_355/A INVX1_LOC_479/A 0.00fF
C9323 INVX1_LOC_249/Y INVX1_LOC_74/Y 0.01fF
C9324 INVX1_LOC_412/Y INVX1_LOC_634/Y 0.08fF
C9325 NAND2X1_LOC_410/a_36_24# INVX1_LOC_9/Y -0.02fF
C9326 INVX1_LOC_255/Y INVX1_LOC_354/A 0.00fF
C9327 NAND2X1_LOC_700/a_36_24# NAND2X1_LOC_274/B 0.00fF
C9328 NAND2X1_LOC_122/Y INVX1_LOC_74/Y 0.80fF
C9329 INVX1_LOC_442/A NAND2X1_LOC_62/a_36_24# 0.01fF
C9330 INVX1_LOC_49/Y NAND2X1_LOC_416/Y 0.03fF
C9331 INVX1_LOC_48/Y INVX1_LOC_601/Y 0.03fF
C9332 INVX1_LOC_582/Y INVX1_LOC_62/Y 0.01fF
C9333 NAND2X1_LOC_707/A INVX1_LOC_148/Y 0.00fF
C9334 INVX1_LOC_31/Y NAND2X1_LOC_615/B 0.03fF
C9335 INVX1_LOC_137/Y INVX1_LOC_633/A 0.02fF
C9336 INVX1_LOC_507/Y NAND2X1_LOC_612/A 0.01fF
C9337 INVX1_LOC_45/Y INVX1_LOC_528/Y 0.00fF
C9338 NAND2X1_LOC_620/a_36_24# INVX1_LOC_62/Y 0.01fF
C9339 INVX1_LOC_399/Y NAND2X1_LOC_237/Y 0.02fF
C9340 INVX1_LOC_338/Y INVX1_LOC_98/Y 0.33fF
C9341 NAND2X1_LOC_128/B INVX1_LOC_118/A 0.05fF
C9342 NAND2X1_LOC_427/Y INVX1_LOC_505/Y 0.13fF
C9343 NAND2X1_LOC_387/Y INVX1_LOC_589/Y 0.01fF
C9344 INVX1_LOC_588/Y NAND2X1_LOC_837/A 0.01fF
C9345 INVX1_LOC_188/Y INVX1_LOC_119/Y 0.11fF
C9346 INVX1_LOC_84/A INVX1_LOC_62/Y 0.08fF
C9347 NAND2X1_LOC_845/B INVX1_LOC_99/Y 0.02fF
C9348 NAND2X1_LOC_13/Y INVX1_LOC_479/A 0.04fF
C9349 INVX1_LOC_21/Y NAND2X1_LOC_786/B 0.56fF
C9350 NAND2X1_LOC_542/A INPUT_1 0.03fF
C9351 INVX1_LOC_344/Y INVX1_LOC_114/A 0.03fF
C9352 INVX1_LOC_86/Y INVX1_LOC_182/Y 0.01fF
C9353 NAND2X1_LOC_387/Y INVX1_LOC_47/Y 0.00fF
C9354 INVX1_LOC_17/Y NAND2X1_LOC_434/B 0.01fF
C9355 INVX1_LOC_400/A INVX1_LOC_179/A 0.02fF
C9356 NAND2X1_LOC_334/A INVX1_LOC_50/Y 0.03fF
C9357 INVX1_LOC_44/A INVX1_LOC_26/Y 0.37fF
C9358 INVX1_LOC_84/A INVX1_LOC_13/Y 0.01fF
C9359 INVX1_LOC_100/Y NAND2X1_LOC_393/Y 0.02fF
C9360 INVX1_LOC_42/Y INVX1_LOC_81/A 0.01fF
C9361 INVX1_LOC_183/Y INVX1_LOC_81/Y 0.02fF
C9362 INVX1_LOC_93/Y INVX1_LOC_255/A 0.01fF
C9363 NAND2X1_LOC_184/Y INVX1_LOC_58/Y 0.17fF
C9364 INVX1_LOC_267/A INVX1_LOC_69/Y 0.01fF
C9365 NAND2X1_LOC_521/a_36_24# INVX1_LOC_26/Y 0.01fF
C9366 INPUT_1 INVX1_LOC_376/Y 0.07fF
C9367 INVX1_LOC_335/Y INVX1_LOC_635/Y 0.03fF
C9368 NAND2X1_LOC_520/A INVX1_LOC_69/Y 0.16fF
C9369 INVX1_LOC_17/Y NAND2X1_LOC_629/a_36_24# 0.00fF
C9370 INVX1_LOC_417/A INVX1_LOC_75/A 0.04fF
C9371 INVX1_LOC_360/Y INVX1_LOC_41/Y 0.07fF
C9372 INVX1_LOC_47/Y NAND2X1_LOC_684/a_36_24# 0.01fF
C9373 INVX1_LOC_183/A INVX1_LOC_326/Y 0.00fF
C9374 INVX1_LOC_682/Y INVX1_LOC_66/A 0.07fF
C9375 INVX1_LOC_127/Y INVX1_LOC_128/A 0.14fF
C9376 INVX1_LOC_442/Y INVX1_LOC_450/Y 0.04fF
C9377 INVX1_LOC_58/Y INVX1_LOC_498/Y 0.18fF
C9378 INVX1_LOC_116/Y NAND2X1_LOC_62/a_36_24# 0.01fF
C9379 INVX1_LOC_551/A INVX1_LOC_58/Y 0.00fF
C9380 INVX1_LOC_105/A INVX1_LOC_41/Y 0.04fF
C9381 INVX1_LOC_47/Y NAND2X1_LOC_845/B 0.02fF
C9382 INVX1_LOC_79/A INVX1_LOC_230/Y 0.04fF
C9383 INVX1_LOC_50/Y NAND2X1_LOC_609/B 0.06fF
C9384 INVX1_LOC_203/A NAND2X1_LOC_333/B 0.05fF
C9385 INVX1_LOC_641/Y INVX1_LOC_454/Y 0.04fF
C9386 INVX1_LOC_281/A INVX1_LOC_280/A 0.10fF
C9387 INVX1_LOC_194/Y INVX1_LOC_666/Y 0.09fF
C9388 INVX1_LOC_63/Y NAND2X1_LOC_833/B 0.02fF
C9389 INVX1_LOC_145/A INVX1_LOC_41/Y 0.13fF
C9390 INVX1_LOC_31/Y NAND2X1_LOC_621/B 0.05fF
C9391 INVX1_LOC_117/Y NAND2X1_LOC_619/a_36_24# 0.01fF
C9392 INVX1_LOC_62/Y INVX1_LOC_496/A 0.66fF
C9393 INVX1_LOC_75/Y INVX1_LOC_58/Y 0.00fF
C9394 INVX1_LOC_479/A INVX1_LOC_361/A 0.03fF
C9395 VDD NAND2X1_LOC_710/B 0.04fF
C9396 INVX1_LOC_69/Y NAND2X1_LOC_227/A 0.01fF
C9397 INVX1_LOC_438/A INVX1_LOC_206/Y 0.01fF
C9398 INVX1_LOC_80/A INVX1_LOC_109/Y 0.03fF
C9399 VDD INVX1_LOC_255/Y 0.44fF
C9400 NAND2X1_LOC_122/Y NAND2X1_LOC_591/B 0.00fF
C9401 INVX1_LOC_477/Y INVX1_LOC_92/A 0.01fF
C9402 NAND2X1_LOC_847/A NAND2X1_LOC_245/a_36_24# 0.00fF
C9403 INPUT_0 NAND2X1_LOC_154/a_36_24# 0.00fF
C9404 VDD INVX1_LOC_577/Y 0.25fF
C9405 INPUT_0 NAND2X1_LOC_690/Y 0.01fF
C9406 INVX1_LOC_629/A NAND2X1_LOC_122/Y 0.03fF
C9407 NAND2X1_LOC_242/A INVX1_LOC_273/A 0.01fF
C9408 INVX1_LOC_395/A INVX1_LOC_442/A 0.17fF
C9409 NAND2X1_LOC_710/B INVX1_LOC_510/Y 0.10fF
C9410 NAND2X1_LOC_317/A NAND2X1_LOC_704/B 0.07fF
C9411 INVX1_LOC_11/Y INVX1_LOC_109/Y 0.07fF
C9412 NAND2X1_LOC_721/a_36_24# INVX1_LOC_586/A 0.00fF
C9413 INVX1_LOC_551/Y INVX1_LOC_553/Y 0.04fF
C9414 NAND2X1_LOC_24/Y NAND2X1_LOC_45/Y 0.19fF
C9415 VDD INVX1_LOC_474/Y 0.21fF
C9416 INVX1_LOC_551/Y INVX1_LOC_375/A 0.03fF
C9417 INVX1_LOC_185/A INVX1_LOC_492/A 0.00fF
C9418 INVX1_LOC_449/A NAND2X1_LOC_541/a_36_24# 0.00fF
C9419 INVX1_LOC_603/Y NAND2X1_LOC_475/A 0.01fF
C9420 INVX1_LOC_434/A NAND2X1_LOC_260/Y 0.07fF
C9421 INVX1_LOC_372/Y INVX1_LOC_355/A 0.02fF
C9422 NAND2X1_LOC_373/Y INVX1_LOC_304/A 0.01fF
C9423 NAND2X1_LOC_373/Y INVX1_LOC_35/Y 0.12fF
C9424 INVX1_LOC_395/Y INVX1_LOC_615/A 0.04fF
C9425 VDD INVX1_LOC_444/Y 0.46fF
C9426 VDD INVX1_LOC_481/Y 0.21fF
C9427 INVX1_LOC_447/A INVX1_LOC_145/Y 0.04fF
C9428 INVX1_LOC_449/A INVX1_LOC_393/Y 0.00fF
C9429 NAND2X1_LOC_636/A INVX1_LOC_54/Y 0.15fF
C9430 INPUT_0 NAND2X1_LOC_266/a_36_24# 0.00fF
C9431 INVX1_LOC_20/Y INVX1_LOC_291/A 0.15fF
C9432 INVX1_LOC_679/Y NAND2X1_LOC_142/Y 0.01fF
C9433 INVX1_LOC_191/Y INVX1_LOC_198/A 0.02fF
C9434 INVX1_LOC_395/A INVX1_LOC_116/Y 0.07fF
C9435 INVX1_LOC_76/Y INVX1_LOC_197/A 0.01fF
C9436 NAND2X1_LOC_336/B NAND2X1_LOC_538/B 0.01fF
C9437 NAND2X1_LOC_498/Y INVX1_LOC_504/Y 0.21fF
C9438 NAND2X1_LOC_788/A INVX1_LOC_31/Y 0.03fF
C9439 INVX1_LOC_628/A NAND2X1_LOC_122/Y 0.03fF
C9440 INVX1_LOC_584/A INVX1_LOC_259/Y 0.01fF
C9441 INVX1_LOC_224/Y INVX1_LOC_117/Y 1.54fF
C9442 INVX1_LOC_402/Y INVX1_LOC_586/A 0.03fF
C9443 INVX1_LOC_236/A INVX1_LOC_521/Y 0.20fF
C9444 INVX1_LOC_418/Y INVX1_LOC_412/A 0.02fF
C9445 NAND2X1_LOC_363/a_36_24# INVX1_LOC_381/A 0.00fF
C9446 INVX1_LOC_412/A INVX1_LOC_159/Y 0.00fF
C9447 NAND2X1_LOC_13/Y INVX1_LOC_12/Y 0.02fF
C9448 INVX1_LOC_412/Y INVX1_LOC_46/Y 0.03fF
C9449 INVX1_LOC_45/A INVX1_LOC_29/Y 0.01fF
C9450 NAND2X1_LOC_394/a_36_24# INVX1_LOC_183/A 0.00fF
C9451 INVX1_LOC_211/Y INVX1_LOC_321/A 0.00fF
C9452 INVX1_LOC_364/Y INVX1_LOC_370/A 0.16fF
C9453 INVX1_LOC_578/A INVX1_LOC_117/Y 0.07fF
C9454 NAND2X1_LOC_615/Y INVX1_LOC_388/Y 0.01fF
C9455 INVX1_LOC_206/Y NAND2X1_LOC_388/A 0.11fF
C9456 INVX1_LOC_51/Y INVX1_LOC_159/A 0.04fF
C9457 INVX1_LOC_522/Y NAND2X1_LOC_612/A 0.02fF
C9458 INVX1_LOC_53/Y NAND2X1_LOC_527/a_36_24# 0.01fF
C9459 INVX1_LOC_570/Y INVX1_LOC_569/Y 0.13fF
C9460 INVX1_LOC_180/A INVX1_LOC_198/A 0.05fF
C9461 NAND2X1_LOC_341/a_36_24# INVX1_LOC_94/A 0.00fF
C9462 INVX1_LOC_522/Y INVX1_LOC_145/Y 0.12fF
C9463 INVX1_LOC_683/Y INVX1_LOC_116/Y 0.00fF
C9464 INVX1_LOC_544/A INVX1_LOC_683/Y 0.01fF
C9465 INVX1_LOC_442/A INVX1_LOC_31/Y 0.08fF
C9466 INVX1_LOC_84/A INVX1_LOC_42/Y 0.84fF
C9467 INVX1_LOC_196/A INVX1_LOC_189/Y 0.00fF
C9468 INVX1_LOC_321/A INVX1_LOC_46/Y 0.03fF
C9469 NAND2X1_LOC_513/Y NAND2X1_LOC_307/B 0.12fF
C9470 INVX1_LOC_542/A INVX1_LOC_496/Y 0.01fF
C9471 NAND2X1_LOC_320/Y INVX1_LOC_80/A 0.00fF
C9472 INVX1_LOC_20/Y INVX1_LOC_360/A 0.00fF
C9473 INVX1_LOC_435/A INVX1_LOC_312/Y 0.19fF
C9474 NAND2X1_LOC_513/A INVX1_LOC_14/A 0.24fF
C9475 INVX1_LOC_11/Y INVX1_LOC_126/Y 0.06fF
C9476 VDD INVX1_LOC_128/Y 0.30fF
C9477 VDD INVX1_LOC_26/Y 1.67fF
C9478 INVX1_LOC_566/A NAND2X1_LOC_406/a_36_24# -0.02fF
C9479 INVX1_LOC_51/Y INVX1_LOC_66/A 0.17fF
C9480 INVX1_LOC_134/Y INVX1_LOC_370/A 0.01fF
C9481 NAND2X1_LOC_61/A INVX1_LOC_41/Y 0.07fF
C9482 INVX1_LOC_90/Y NAND2X1_LOC_76/B 0.01fF
C9483 INPUT_0 NAND2X1_LOC_467/a_36_24# 0.00fF
C9484 NAND2X1_LOC_97/B INVX1_LOC_202/Y 0.02fF
C9485 NAND2X1_LOC_336/B INVX1_LOC_159/Y 0.52fF
C9486 INVX1_LOC_417/Y INVX1_LOC_545/A 0.02fF
C9487 INVX1_LOC_607/A INVX1_LOC_58/Y 0.02fF
C9488 INVX1_LOC_395/A INVX1_LOC_179/A 0.03fF
C9489 INVX1_LOC_386/Y NAND2X1_LOC_416/Y 0.03fF
C9490 NAND2X1_LOC_520/A INVX1_LOC_586/A 0.02fF
C9491 INVX1_LOC_119/A INVX1_LOC_46/Y 0.04fF
C9492 INVX1_LOC_617/Y INVX1_LOC_46/Y 0.03fF
C9493 NAND2X1_LOC_140/B INVX1_LOC_35/Y 0.16fF
C9494 INVX1_LOC_12/Y NAND2X1_LOC_670/a_36_24# 0.01fF
C9495 INVX1_LOC_584/A INVX1_LOC_114/A 0.02fF
C9496 INVX1_LOC_84/A INVX1_LOC_87/A 0.00fF
C9497 INVX1_LOC_11/Y NAND2X1_LOC_320/Y 0.00fF
C9498 INVX1_LOC_232/Y INVX1_LOC_48/Y 0.02fF
C9499 INVX1_LOC_632/A INVX1_LOC_497/Y 0.02fF
C9500 INVX1_LOC_288/Y INVX1_LOC_505/A 0.00fF
C9501 INVX1_LOC_602/A INVX1_LOC_93/A 0.02fF
C9502 NAND2X1_LOC_378/a_36_24# INVX1_LOC_41/Y 0.00fF
C9503 INVX1_LOC_183/A NAND2X1_LOC_6/a_36_24# 0.00fF
C9504 INVX1_LOC_69/Y INVX1_LOC_59/A 0.04fF
C9505 INVX1_LOC_535/Y NAND2X1_LOC_677/Y 0.01fF
C9506 NAND2X1_LOC_370/A INVX1_LOC_79/A 0.00fF
C9507 INVX1_LOC_383/A INVX1_LOC_128/Y 0.01fF
C9508 NAND2X1_LOC_24/Y INVX1_LOC_47/Y 0.03fF
C9509 INVX1_LOC_543/Y INVX1_LOC_7/Y 0.09fF
C9510 INVX1_LOC_54/Y INVX1_LOC_230/A 0.47fF
C9511 INVX1_LOC_268/A INVX1_LOC_31/Y 0.05fF
C9512 INVX1_LOC_53/Y INVX1_LOC_234/Y 0.01fF
C9513 INVX1_LOC_80/A INVX1_LOC_199/Y 0.09fF
C9514 NAND2X1_LOC_122/Y INVX1_LOC_79/A 0.03fF
C9515 INVX1_LOC_352/A INVX1_LOC_374/Y 0.00fF
C9516 INVX1_LOC_619/A INVX1_LOC_181/Y 0.04fF
C9517 INVX1_LOC_273/A INVX1_LOC_79/A 0.14fF
C9518 NAND2X1_LOC_442/a_36_24# INVX1_LOC_98/Y 0.06fF
C9519 INVX1_LOC_267/Y INVX1_LOC_49/Y 0.03fF
C9520 INVX1_LOC_89/Y NAND2X1_LOC_284/a_36_24# -0.00fF
C9521 INVX1_LOC_31/Y INVX1_LOC_116/Y 0.03fF
C9522 INVX1_LOC_45/Y INVX1_LOC_41/Y 6.00fF
C9523 INVX1_LOC_12/Y INVX1_LOC_361/A 0.04fF
C9524 INVX1_LOC_48/Y INVX1_LOC_189/A 0.07fF
C9525 INVX1_LOC_97/Y INVX1_LOC_44/Y 0.04fF
C9526 INVX1_LOC_254/A NAND2X1_LOC_615/B 0.00fF
C9527 INVX1_LOC_31/Y NAND2X1_LOC_432/Y -0.07fF
C9528 INVX1_LOC_48/Y INVX1_LOC_230/Y 0.05fF
C9529 INVX1_LOC_400/A INVX1_LOC_69/Y 0.07fF
C9530 NAND2X1_LOC_387/Y INVX1_LOC_153/A 0.02fF
C9531 INVX1_LOC_186/A INVX1_LOC_168/Y 0.03fF
C9532 INVX1_LOC_556/Y NAND2X1_LOC_284/A 0.01fF
C9533 INVX1_LOC_42/A INVX1_LOC_26/Y 0.02fF
C9534 NAND2X1_LOC_756/Y INVX1_LOC_531/Y 0.11fF
C9535 INVX1_LOC_11/Y INVX1_LOC_199/Y 0.14fF
C9536 INVX1_LOC_330/A INVX1_LOC_331/Y 0.00fF
C9537 INVX1_LOC_651/Y NAND2X1_LOC_843/B 0.73fF
C9538 INVX1_LOC_451/A INVX1_LOC_63/Y 0.03fF
C9539 INVX1_LOC_49/Y INVX1_LOC_510/A 0.02fF
C9540 INVX1_LOC_492/A INVX1_LOC_58/Y 0.04fF
C9541 INVX1_LOC_356/A INVX1_LOC_74/Y 0.14fF
C9542 INVX1_LOC_100/Y INVX1_LOC_519/A 0.03fF
C9543 NAND2X1_LOC_542/A INVX1_LOC_50/Y 0.03fF
C9544 NAND2X1_LOC_700/a_36_24# INVX1_LOC_468/A 0.00fF
C9545 INVX1_LOC_444/Y INVX1_LOC_339/Y 0.10fF
C9546 INVX1_LOC_682/Y INVX1_LOC_116/Y 0.18fF
C9547 INVX1_LOC_53/Y INVX1_LOC_665/A 0.03fF
C9548 NAND2X1_LOC_320/Y NAND2X1_LOC_433/Y 0.00fF
C9549 INVX1_LOC_602/A INVX1_LOC_621/A 0.21fF
C9550 NAND2X1_LOC_387/Y INVX1_LOC_96/A 0.01fF
C9551 INVX1_LOC_435/A INVX1_LOC_225/Y 0.02fF
C9552 INVX1_LOC_556/Y NAND2X1_LOC_768/B 0.01fF
C9553 INVX1_LOC_323/Y INVX1_LOC_100/Y 0.05fF
C9554 INVX1_LOC_20/Y NAND2X1_LOC_71/a_36_24# 0.00fF
C9555 GATE_579 INVX1_LOC_443/A 0.19fF
C9556 INVX1_LOC_93/Y INVX1_LOC_69/Y 0.58fF
C9557 INVX1_LOC_467/Y INVX1_LOC_58/Y 0.01fF
C9558 INVX1_LOC_625/A INVX1_LOC_90/Y 0.02fF
C9559 NAND2X1_LOC_586/a_36_24# NAND2X1_LOC_586/Y 0.02fF
C9560 INVX1_LOC_369/A NAND2X1_LOC_488/Y 0.01fF
C9561 INVX1_LOC_117/Y INVX1_LOC_120/Y 0.02fF
C9562 INVX1_LOC_31/Y INVX1_LOC_255/A 0.07fF
C9563 INVX1_LOC_134/Y INVX1_LOC_588/A 0.09fF
C9564 INVX1_LOC_376/Y INVX1_LOC_50/Y 0.07fF
C9565 INVX1_LOC_79/Y INVX1_LOC_600/Y 0.01fF
C9566 INVX1_LOC_525/Y INVX1_LOC_49/Y 0.23fF
C9567 INVX1_LOC_306/Y NAND2X1_LOC_376/B 0.27fF
C9568 INVX1_LOC_41/Y NAND2X1_LOC_376/Y 0.02fF
C9569 INVX1_LOC_361/Y INVX1_LOC_518/A 0.07fF
C9570 INVX1_LOC_442/Y INVX1_LOC_280/A 0.02fF
C9571 INVX1_LOC_294/A INVX1_LOC_90/Y 0.01fF
C9572 INVX1_LOC_442/Y NAND2X1_LOC_372/Y 0.07fF
C9573 INVX1_LOC_573/Y INVX1_LOC_582/A 0.02fF
C9574 NAND2X1_LOC_847/A INVX1_LOC_212/Y 0.04fF
C9575 INVX1_LOC_26/Y NAND2X1_LOC_243/A 0.66fF
C9576 INVX1_LOC_103/Y INVX1_LOC_26/Y 0.00fF
C9577 INVX1_LOC_241/A INVX1_LOC_241/Y 0.01fF
C9578 INVX1_LOC_649/A INVX1_LOC_655/A 0.04fF
C9579 INVX1_LOC_103/Y INVX1_LOC_128/Y 0.18fF
C9580 INVX1_LOC_513/Y INVX1_LOC_58/Y 0.03fF
C9581 INVX1_LOC_258/Y INVX1_LOC_347/Y 0.01fF
C9582 INVX1_LOC_662/A NAND2X1_LOC_814/Y 0.03fF
C9583 INVX1_LOC_69/Y NAND2X1_LOC_334/B 0.02fF
C9584 INVX1_LOC_62/A INVX1_LOC_62/Y 0.01fF
C9585 INVX1_LOC_117/Y INVX1_LOC_621/A 0.06fF
C9586 INVX1_LOC_48/Y INVX1_LOC_598/Y 0.00fF
C9587 INVX1_LOC_100/Y NAND2X1_LOC_846/A 0.01fF
C9588 NAND2X1_LOC_635/B NAND2X1_LOC_428/Y 0.00fF
C9589 INVX1_LOC_153/A INVX1_LOC_91/A 0.02fF
C9590 INVX1_LOC_90/Y NAND2X1_LOC_52/Y 0.01fF
C9591 VDD INVX1_LOC_426/Y 0.23fF
C9592 INVX1_LOC_665/A NAND2X1_LOC_274/Y 0.01fF
C9593 NAND2X1_LOC_532/Y INVX1_LOC_62/Y 0.05fF
C9594 NAND2X1_LOC_276/A INVX1_LOC_41/Y 0.02fF
C9595 GATE_662 NAND2X1_LOC_843/B 0.03fF
C9596 VDD NAND2X1_LOC_249/Y 0.47fF
C9597 INVX1_LOC_404/Y INVX1_LOC_405/A 0.04fF
C9598 VDD INVX1_LOC_238/A -0.00fF
C9599 INVX1_LOC_479/A NAND2X1_LOC_449/B 0.01fF
C9600 INVX1_LOC_26/Y NAND2X1_LOC_786/B 0.00fF
C9601 INVX1_LOC_659/A INVX1_LOC_74/Y 0.08fF
C9602 INVX1_LOC_659/A INVX1_LOC_660/A 0.07fF
C9603 NAND2X1_LOC_107/a_36_24# NAND2X1_LOC_248/B 0.00fF
C9604 NAND2X1_LOC_393/a_36_24# INVX1_LOC_206/Y 0.00fF
C9605 NAND2X1_LOC_157/a_36_24# NAND2X1_LOC_409/Y 0.02fF
C9606 INVX1_LOC_275/A INVX1_LOC_94/A 0.06fF
C9607 VDD INVX1_LOC_564/Y 0.14fF
C9608 INVX1_LOC_75/Y INVX1_LOC_245/A 0.11fF
C9609 INPUT_0 INVX1_LOC_97/A 0.37fF
C9610 INVX1_LOC_26/Y INVX1_LOC_635/Y 0.03fF
C9611 INVX1_LOC_279/A INVX1_LOC_220/Y 0.00fF
C9612 NAND2X1_LOC_544/a_36_24# NAND2X1_LOC_373/Y 0.00fF
C9613 INVX1_LOC_445/Y INVX1_LOC_278/A 0.00fF
C9614 NAND2X1_LOC_543/B NAND2X1_LOC_180/B 0.05fF
C9615 NAND2X1_LOC_516/Y NAND2X1_LOC_317/B 0.01fF
C9616 INVX1_LOC_366/A INVX1_LOC_616/Y 0.03fF
C9617 NAND2X1_LOC_475/A INVX1_LOC_269/A 0.03fF
C9618 INVX1_LOC_168/Y INVX1_LOC_611/A 0.02fF
C9619 INVX1_LOC_62/Y INVX1_LOC_135/Y 0.02fF
C9620 INVX1_LOC_76/A INVX1_LOC_9/Y 0.06fF
C9621 INPUT_0 INVX1_LOC_169/A 0.01fF
C9622 INVX1_LOC_160/Y INVX1_LOC_45/Y 0.03fF
C9623 INVX1_LOC_442/A INVX1_LOC_51/Y 0.01fF
C9624 VDD INVX1_LOC_369/A 0.06fF
C9625 NAND2X1_LOC_585/a_36_24# INVX1_LOC_632/A 0.01fF
C9626 INVX1_LOC_315/Y INVX1_LOC_45/Y 1.49fF
C9627 INVX1_LOC_600/A NAND2X1_LOC_772/a_36_24# 0.02fF
C9628 INVX1_LOC_20/Y NAND2X1_LOC_589/a_36_24# 0.00fF
C9629 INVX1_LOC_629/A INVX1_LOC_579/A 0.02fF
C9630 INPUT_0 INVX1_LOC_633/Y 0.03fF
C9631 INVX1_LOC_62/Y INVX1_LOC_76/A 0.09fF
C9632 INVX1_LOC_266/A INVX1_LOC_442/A 1.30fF
C9633 VDD NAND2X1_LOC_275/Y 0.12fF
C9634 NAND2X1_LOC_76/B INVX1_LOC_98/Y 0.20fF
C9635 INVX1_LOC_412/Y INVX1_LOC_115/A 0.01fF
C9636 INVX1_LOC_68/Y NAND2X1_LOC_357/a_36_24# 0.00fF
C9637 INVX1_LOC_618/A INVX1_LOC_66/A 0.07fF
C9638 VDD INVX1_LOC_58/A -0.00fF
C9639 INVX1_LOC_20/Y NAND2X1_LOC_315/a_36_24# 0.00fF
C9640 INVX1_LOC_586/A INVX1_LOC_367/A 0.00fF
C9641 INVX1_LOC_201/A INVX1_LOC_97/A 0.01fF
C9642 INVX1_LOC_133/Y INVX1_LOC_476/Y 0.03fF
C9643 NAND2X1_LOC_152/Y INVX1_LOC_569/A 0.06fF
C9644 INVX1_LOC_33/Y INVX1_LOC_310/Y 0.08fF
C9645 INVX1_LOC_45/Y INVX1_LOC_358/Y 0.00fF
C9646 NAND2X1_LOC_122/Y INVX1_LOC_632/A 0.03fF
C9647 INVX1_LOC_158/Y INVX1_LOC_560/A 0.06fF
C9648 INVX1_LOC_445/Y INVX1_LOC_453/Y 0.80fF
C9649 INVX1_LOC_335/Y INVX1_LOC_45/Y 0.06fF
C9650 INVX1_LOC_44/Y INVX1_LOC_615/A 0.03fF
C9651 NAND2X1_LOC_548/B INVX1_LOC_171/Y 0.12fF
C9652 INVX1_LOC_21/Y INVX1_LOC_45/Y 0.32fF
C9653 INVX1_LOC_578/A NAND2X1_LOC_143/a_36_24# 0.01fF
C9654 INVX1_LOC_121/Y INVX1_LOC_50/Y 0.34fF
C9655 NAND2X1_LOC_97/B INVX1_LOC_76/Y 0.02fF
C9656 NAND2X1_LOC_543/a_36_24# INVX1_LOC_270/A 0.01fF
C9657 INVX1_LOC_686/A INVX1_LOC_111/A 0.00fF
C9658 INVX1_LOC_206/Y INVX1_LOC_117/Y 0.35fF
C9659 INVX1_LOC_557/A INVX1_LOC_251/Y 0.05fF
C9660 INVX1_LOC_255/Y INVX1_LOC_360/Y 0.09fF
C9661 INVX1_LOC_173/A INVX1_LOC_145/Y 0.03fF
C9662 INVX1_LOC_459/A INVX1_LOC_501/A 0.01fF
C9663 INVX1_LOC_6/Y INVX1_LOC_616/Y 0.01fF
C9664 INVX1_LOC_51/Y INVX1_LOC_116/Y 0.09fF
C9665 INVX1_LOC_312/Y INVX1_LOC_367/A 0.07fF
C9666 INVX1_LOC_544/A INVX1_LOC_51/Y 0.03fF
C9667 INVX1_LOC_421/A NAND2X1_LOC_457/A 0.03fF
C9668 NAND2X1_LOC_370/A INVX1_LOC_48/Y 0.03fF
C9669 INVX1_LOC_286/Y INVX1_LOC_155/Y 0.01fF
C9670 INVX1_LOC_410/Y INVX1_LOC_46/Y 0.03fF
C9671 INVX1_LOC_276/A NAND2X1_LOC_285/B 0.00fF
C9672 INVX1_LOC_53/Y INVX1_LOC_80/A 0.30fF
C9673 INVX1_LOC_21/Y INPUT_3 0.12fF
C9674 INVX1_LOC_375/A INVX1_LOC_46/Y 0.03fF
C9675 INVX1_LOC_53/Y NAND2X1_LOC_768/A 0.18fF
C9676 NAND2X1_LOC_122/Y INVX1_LOC_48/Y 0.03fF
C9677 INVX1_LOC_546/A INVX1_LOC_46/Y 0.02fF
C9678 INVX1_LOC_53/Y INVX1_LOC_579/Y 0.14fF
C9679 INVX1_LOC_276/A NAND2X1_LOC_106/B 0.01fF
C9680 INVX1_LOC_266/A INVX1_LOC_116/Y 0.26fF
C9681 INVX1_LOC_114/Y INVX1_LOC_259/Y 0.00fF
C9682 INVX1_LOC_45/Y NAND2X1_LOC_267/A 0.07fF
C9683 INVX1_LOC_224/Y INVX1_LOC_58/Y 0.07fF
C9684 INVX1_LOC_393/A INVX1_LOC_32/Y 0.01fF
C9685 INVX1_LOC_628/A INVX1_LOC_579/A 0.02fF
C9686 INVX1_LOC_273/A INVX1_LOC_48/Y 0.00fF
C9687 NAND2X1_LOC_123/A INVX1_LOC_633/Y 0.04fF
C9688 INVX1_LOC_17/Y INVX1_LOC_634/A 0.01fF
C9689 INVX1_LOC_93/Y NAND2X1_LOC_419/a_36_24# 0.01fF
C9690 VDD NAND2X1_LOC_605/B 0.04fF
C9691 INVX1_LOC_395/A INVX1_LOC_69/Y 0.37fF
C9692 INVX1_LOC_435/A INVX1_LOC_486/Y 0.07fF
C9693 NAND2X1_LOC_331/A INVX1_LOC_496/A 0.09fF
C9694 INVX1_LOC_93/Y INVX1_LOC_586/A 0.72fF
C9695 INVX1_LOC_435/A INVX1_LOC_294/Y 0.01fF
C9696 INVX1_LOC_117/Y INVX1_LOC_242/A 0.07fF
C9697 INVX1_LOC_555/A INVX1_LOC_185/Y 0.03fF
C9698 INVX1_LOC_256/A INVX1_LOC_197/A 0.02fF
C9699 INVX1_LOC_288/Y INVX1_LOC_675/Y 0.01fF
C9700 INVX1_LOC_174/Y INVX1_LOC_87/A 0.01fF
C9701 INVX1_LOC_84/A INVX1_LOC_480/Y 0.05fF
C9702 NAND2X1_LOC_673/a_36_24# INVX1_LOC_600/A 0.00fF
C9703 INVX1_LOC_254/Y INVX1_LOC_551/Y 1.24fF
C9704 NAND2X1_LOC_13/Y NAND2X1_LOC_615/B 0.27fF
C9705 INVX1_LOC_89/Y INVX1_LOC_624/A 0.01fF
C9706 VDD INVX1_LOC_632/Y 0.31fF
C9707 INVX1_LOC_578/A INVX1_LOC_58/Y 0.07fF
C9708 INVX1_LOC_21/Y NAND2X1_LOC_376/Y 0.02fF
C9709 INVX1_LOC_362/Y INVX1_LOC_69/Y 0.03fF
C9710 INVX1_LOC_11/Y INVX1_LOC_53/Y 10.44fF
C9711 NAND2X1_LOC_416/Y INVX1_LOC_7/Y 0.13fF
C9712 INVX1_LOC_406/Y INVX1_LOC_46/Y 0.03fF
C9713 INVX1_LOC_117/Y INVX1_LOC_686/A 0.07fF
C9714 INVX1_LOC_51/Y INVX1_LOC_255/A 0.03fF
C9715 INVX1_LOC_567/Y INVX1_LOC_35/Y 0.34fF
C9716 NAND2X1_LOC_516/B INVX1_LOC_6/Y 0.02fF
C9717 INVX1_LOC_84/A INVX1_LOC_169/Y 0.10fF
C9718 NAND2X1_LOC_835/A INVX1_LOC_59/A 0.01fF
C9719 INVX1_LOC_625/A INVX1_LOC_98/Y 0.02fF
C9720 INVX1_LOC_312/Y INVX1_LOC_93/Y 0.03fF
C9721 NAND2X1_LOC_704/B INVX1_LOC_199/Y 0.75fF
C9722 INVX1_LOC_372/Y INVX1_LOC_359/A 0.16fF
C9723 INVX1_LOC_65/Y INVX1_LOC_351/A 0.01fF
C9724 NAND2X1_LOC_781/A INVX1_LOC_93/Y 0.01fF
C9725 INVX1_LOC_100/Y INVX1_LOC_445/A 0.45fF
C9726 INVX1_LOC_201/Y NAND2X1_LOC_226/Y 0.15fF
C9727 INVX1_LOC_451/A NAND2X1_LOC_414/a_36_24# 0.06fF
C9728 INVX1_LOC_586/A INVX1_LOC_390/A 0.03fF
C9729 NAND2X1_LOC_598/a_36_24# INVX1_LOC_588/A 0.01fF
C9730 INVX1_LOC_44/A INVX1_LOC_81/Y 0.01fF
C9731 INVX1_LOC_266/A INVX1_LOC_255/A 0.10fF
C9732 INVX1_LOC_99/Y INVX1_LOC_259/Y 0.04fF
C9733 INVX1_LOC_54/Y NAND2X1_LOC_72/Y 0.72fF
C9734 INVX1_LOC_20/Y NAND2X1_LOC_686/B 0.01fF
C9735 NAND2X1_LOC_498/Y INVX1_LOC_114/A 0.41fF
C9736 INVX1_LOC_683/Y INVX1_LOC_69/Y 0.00fF
C9737 INVX1_LOC_586/A NAND2X1_LOC_334/B 0.15fF
C9738 INVX1_LOC_674/A NAND2X1_LOC_755/B 0.02fF
C9739 INVX1_LOC_617/Y INVX1_LOC_49/Y 0.07fF
C9740 NAND2X1_LOC_181/A INVX1_LOC_519/A 0.61fF
C9741 INVX1_LOC_65/Y INVX1_LOC_90/Y 0.07fF
C9742 INVX1_LOC_587/A NAND2X1_LOC_822/a_36_24# 0.00fF
C9743 INVX1_LOC_581/A INVX1_LOC_476/Y 0.08fF
C9744 INVX1_LOC_296/Y INVX1_LOC_431/Y 0.01fF
C9745 INVX1_LOC_402/Y INVX1_LOC_6/Y 0.09fF
C9746 NAND2X1_LOC_325/B INVX1_LOC_257/A 0.02fF
C9747 INVX1_LOC_97/A INVX1_LOC_211/A 0.65fF
C9748 INVX1_LOC_63/Y INVX1_LOC_134/Y 0.20fF
C9749 INVX1_LOC_47/Y NAND2X1_LOC_423/a_36_24# 0.01fF
C9750 NAND2X1_LOC_32/a_36_24# INVX1_LOC_41/Y 0.00fF
C9751 NAND2X1_LOC_48/Y INVX1_LOC_63/Y 0.00fF
C9752 INVX1_LOC_284/A INVX1_LOC_69/Y 0.00fF
C9753 INVX1_LOC_89/Y INVX1_LOC_230/A 0.07fF
C9754 INVX1_LOC_17/Y NAND2X1_LOC_486/A 0.19fF
C9755 NAND2X1_LOC_174/B INVX1_LOC_32/Y 4.03fF
C9756 INVX1_LOC_468/Y INVX1_LOC_58/Y 0.03fF
C9757 GATE_865 INVX1_LOC_631/Y 0.01fF
C9758 NAND2X1_LOC_591/Y INVX1_LOC_32/Y 0.13fF
C9759 INVX1_LOC_47/Y INVX1_LOC_259/Y 0.03fF
C9760 INVX1_LOC_425/A INVX1_LOC_666/Y 0.07fF
C9761 INPUT_1 NAND2X1_LOC_443/a_36_24# 0.00fF
C9762 INVX1_LOC_619/A INVX1_LOC_26/Y 0.38fF
C9763 INVX1_LOC_173/Y INVX1_LOC_32/Y 0.02fF
C9764 INVX1_LOC_293/Y INVX1_LOC_41/Y 0.10fF
C9765 INVX1_LOC_84/A NAND2X1_LOC_615/a_36_24# 0.01fF
C9766 INVX1_LOC_145/Y NAND2X1_LOC_467/a_36_24# 0.01fF
C9767 INVX1_LOC_116/A NAND2X1_LOC_605/B 0.06fF
C9768 INVX1_LOC_169/A INVX1_LOC_211/A 0.32fF
C9769 INVX1_LOC_551/Y INVX1_LOC_479/A 0.16fF
C9770 NAND2X1_LOC_615/B INVX1_LOC_361/A 0.01fF
C9771 INVX1_LOC_376/Y NAND2X1_LOC_648/a_36_24# 0.00fF
C9772 INVX1_LOC_479/Y INVX1_LOC_351/A 0.03fF
C9773 INVX1_LOC_99/Y INVX1_LOC_114/A 0.06fF
C9774 INVX1_LOC_47/Y NAND2X1_LOC_707/B 0.03fF
C9775 NAND2X1_LOC_521/Y NAND2X1_LOC_523/a_36_24# 0.01fF
C9776 NAND2X1_LOC_334/a_36_24# INVX1_LOC_79/A 0.00fF
C9777 INVX1_LOC_31/Y INVX1_LOC_69/Y 0.23fF
C9778 INVX1_LOC_578/Y INVX1_LOC_347/Y 0.00fF
C9779 NAND2X1_LOC_818/a_36_24# NAND2X1_LOC_843/B 0.00fF
C9780 NAND2X1_LOC_186/a_36_24# INVX1_LOC_496/A 0.00fF
C9781 INVX1_LOC_160/A INVX1_LOC_41/Y 0.03fF
C9782 INVX1_LOC_411/A INVX1_LOC_242/Y 0.04fF
C9783 INVX1_LOC_479/Y INVX1_LOC_90/Y 0.01fF
C9784 INVX1_LOC_16/Y INVX1_LOC_588/A 0.01fF
C9785 INVX1_LOC_641/A INVX1_LOC_69/Y 0.06fF
C9786 INVX1_LOC_105/A INVX1_LOC_128/Y 0.02fF
C9787 INVX1_LOC_685/Y INVX1_LOC_454/Y 0.00fF
C9788 INVX1_LOC_394/Y INVX1_LOC_615/A 0.09fF
C9789 NAND2X1_LOC_387/Y INVX1_LOC_353/A 0.02fF
C9790 INVX1_LOC_532/Y INVX1_LOC_347/Y 0.00fF
C9791 VDD INVX1_LOC_41/A 0.00fF
C9792 INVX1_LOC_318/A INVX1_LOC_90/Y 0.01fF
C9793 INVX1_LOC_69/Y INVX1_LOC_682/Y 0.01fF
C9794 INVX1_LOC_413/A INVX1_LOC_62/Y 0.02fF
C9795 INVX1_LOC_600/A NAND2X1_LOC_237/a_36_24# 0.01fF
C9796 INVX1_LOC_504/A INVX1_LOC_346/Y 0.05fF
C9797 INVX1_LOC_117/Y NAND2X1_LOC_609/B 0.09fF
C9798 INVX1_LOC_47/Y INVX1_LOC_114/A 0.14fF
C9799 VDD NAND2X1_LOC_790/B 0.73fF
C9800 INVX1_LOC_95/A INVX1_LOC_90/Y 0.01fF
C9801 INVX1_LOC_319/A INVX1_LOC_199/Y 0.03fF
C9802 INVX1_LOC_35/Y INVX1_LOC_485/A 0.02fF
C9803 INVX1_LOC_329/Y NAND2X1_LOC_448/B 0.34fF
C9804 INVX1_LOC_314/Y INVX1_LOC_90/Y 0.05fF
C9805 INVX1_LOC_132/A INVX1_LOC_669/A 0.01fF
C9806 INVX1_LOC_137/Y INVX1_LOC_611/A 0.03fF
C9807 INVX1_LOC_35/Y INVX1_LOC_92/A 0.11fF
C9808 INVX1_LOC_199/Y NAND2X1_LOC_843/B 0.01fF
C9809 INVX1_LOC_304/A INVX1_LOC_92/A 0.00fF
C9810 INVX1_LOC_667/Y INVX1_LOC_655/A 0.00fF
C9811 INVX1_LOC_26/Y NAND2X1_LOC_80/a_36_24# 0.00fF
C9812 VDD INVX1_LOC_122/Y 0.26fF
C9813 INVX1_LOC_321/A INVX1_LOC_297/Y 0.01fF
C9814 NAND2X1_LOC_54/a_36_24# NAND2X1_LOC_513/Y 0.00fF
C9815 INVX1_LOC_119/Y INVX1_LOC_114/A 0.09fF
C9816 VDD INVX1_LOC_373/A 0.00fF
C9817 VDD INVX1_LOC_103/A -0.00fF
C9818 NAND2X1_LOC_45/Y NAND2X1_LOC_457/A 0.01fF
C9819 INVX1_LOC_446/Y NAND2X1_LOC_271/B 0.04fF
C9820 NAND2X1_LOC_475/A NAND2X1_LOC_337/a_36_24# 0.00fF
C9821 INVX1_LOC_272/A INVX1_LOC_91/Y 0.01fF
C9822 NAND2X1_LOC_184/a_36_24# INVX1_LOC_384/A -0.01fF
C9823 INVX1_LOC_613/Y INVX1_LOC_627/A 0.22fF
C9824 INVX1_LOC_613/Y INVX1_LOC_133/Y 0.17fF
C9825 INVX1_LOC_424/A INVX1_LOC_406/Y 0.01fF
C9826 VDD INVX1_LOC_235/Y 0.86fF
C9827 INVX1_LOC_561/Y NAND2X1_LOC_122/Y 0.01fF
C9828 INVX1_LOC_412/Y INVX1_LOC_76/Y 0.03fF
C9829 VDD NAND2X1_LOC_820/Y 0.03fF
C9830 INVX1_LOC_3/Y INVX1_LOC_45/A 0.00fF
C9831 INVX1_LOC_133/Y NAND2X1_LOC_612/A 0.06fF
C9832 INVX1_LOC_395/A INVX1_LOC_586/A 1.63fF
C9833 NAND2X1_LOC_69/B NAND2X1_LOC_616/Y 0.12fF
C9834 INVX1_LOC_255/Y INVX1_LOC_45/Y 0.03fF
C9835 INVX1_LOC_162/Y INVX1_LOC_586/A 0.01fF
C9836 INVX1_LOC_206/Y NAND2X1_LOC_7/a_36_24# 0.00fF
C9837 INVX1_LOC_584/Y NAND2X1_LOC_707/A 0.02fF
C9838 INVX1_LOC_362/Y INVX1_LOC_586/A 0.03fF
C9839 INVX1_LOC_505/A NAND2X1_LOC_801/A 0.01fF
C9840 NAND2X1_LOC_593/a_36_24# INVX1_LOC_288/A 0.00fF
C9841 INVX1_LOC_257/Y INVX1_LOC_633/Y 0.01fF
C9842 INVX1_LOC_321/A INVX1_LOC_76/Y 0.03fF
C9843 INVX1_LOC_312/Y INVX1_LOC_395/A 0.72fF
C9844 NAND2X1_LOC_67/a_36_24# INVX1_LOC_93/Y 0.00fF
C9845 INVX1_LOC_206/Y INVX1_LOC_281/Y 0.03fF
C9846 VDD INVX1_LOC_556/Y 0.89fF
C9847 VDD INVX1_LOC_81/Y 0.46fF
C9848 INVX1_LOC_193/Y INVX1_LOC_99/A 0.01fF
C9849 INVX1_LOC_374/A INVX1_LOC_134/Y 0.03fF
C9850 INVX1_LOC_587/A INVX1_LOC_59/A 0.83fF
C9851 NAND2X1_LOC_271/B INVX1_LOC_145/Y 0.01fF
C9852 INVX1_LOC_312/Y INVX1_LOC_362/Y 0.07fF
C9853 INVX1_LOC_206/Y INVX1_LOC_178/A 0.34fF
C9854 NAND2X1_LOC_595/Y INVX1_LOC_215/Y 0.20fF
C9855 INVX1_LOC_20/Y INVX1_LOC_522/Y 0.07fF
C9856 INVX1_LOC_185/Y INVX1_LOC_474/Y 0.01fF
C9857 INVX1_LOC_395/A NAND2X1_LOC_378/Y 0.03fF
C9858 INVX1_LOC_206/Y NAND2X1_LOC_76/A 0.01fF
C9859 VDD INVX1_LOC_506/A 0.00fF
C9860 NAND2X1_LOC_391/B INVX1_LOC_320/A 0.13fF
C9861 INVX1_LOC_68/Y INVX1_LOC_603/Y 0.03fF
C9862 INVX1_LOC_53/Y NAND2X1_LOC_704/B 0.95fF
C9863 INVX1_LOC_26/Y NAND2X1_LOC_227/a_36_24# 0.00fF
C9864 INVX1_LOC_54/Y NAND2X1_LOC_749/Y 0.03fF
C9865 INVX1_LOC_65/Y INVX1_LOC_98/Y 0.07fF
C9866 INVX1_LOC_444/Y INVX1_LOC_45/Y 0.03fF
C9867 INVX1_LOC_45/Y INVX1_LOC_481/Y 0.01fF
C9868 INVX1_LOC_551/Y INVX1_LOC_12/Y 0.03fF
C9869 INVX1_LOC_390/Y INVX1_LOC_117/Y 0.02fF
C9870 INPUT_0 INVX1_LOC_166/A 0.07fF
C9871 INVX1_LOC_103/A INVX1_LOC_103/Y 0.02fF
C9872 INVX1_LOC_595/Y INVX1_LOC_33/Y 0.14fF
C9873 INVX1_LOC_378/A INVX1_LOC_99/Y 0.03fF
C9874 INVX1_LOC_465/Y INVX1_LOC_501/A 0.01fF
C9875 NAND2X1_LOC_525/Y INVX1_LOC_54/Y 0.29fF
C9876 NAND2X1_LOC_324/B INVX1_LOC_197/A 0.07fF
C9877 INVX1_LOC_20/Y NAND2X1_LOC_448/A 0.02fF
C9878 INVX1_LOC_676/Y NAND2X1_LOC_635/a_36_24# 0.01fF
C9879 INVX1_LOC_169/A INVX1_LOC_145/Y 0.03fF
C9880 INVX1_LOC_68/Y INVX1_LOC_478/Y 0.00fF
C9881 INVX1_LOC_80/A NAND2X1_LOC_148/A 0.04fF
C9882 INVX1_LOC_449/A NAND2X1_LOC_272/a_36_24# 0.00fF
C9883 INVX1_LOC_21/Y INVX1_LOC_293/Y 0.01fF
C9884 NAND2X1_LOC_516/Y INVX1_LOC_166/A 0.03fF
C9885 INVX1_LOC_11/Y NAND2X1_LOC_383/Y 0.10fF
C9886 INVX1_LOC_80/A NAND2X1_LOC_107/Y 1.29fF
C9887 NAND2X1_LOC_775/B NAND2X1_LOC_332/B 0.01fF
C9888 INVX1_LOC_579/A INVX1_LOC_632/A 0.31fF
C9889 INVX1_LOC_397/A INVX1_LOC_117/Y 0.02fF
C9890 INVX1_LOC_353/Y INVX1_LOC_252/Y 0.01fF
C9891 INPUT_0 NAND2X1_LOC_111/Y 0.07fF
C9892 INVX1_LOC_613/Y INVX1_LOC_581/A 0.03fF
C9893 NAND2X1_LOC_314/a_36_24# INVX1_LOC_47/Y 0.01fF
C9894 NAND2X1_LOC_768/A NAND2X1_LOC_107/Y 0.18fF
C9895 NAND2X1_LOC_574/a_36_24# INVX1_LOC_670/A 0.01fF
C9896 INVX1_LOC_206/Y INVX1_LOC_58/Y 0.24fF
C9897 INVX1_LOC_249/Y INVX1_LOC_559/Y 0.00fF
C9898 INPUT_3 INVX1_LOC_444/Y 3.02fF
C9899 INVX1_LOC_553/Y INVX1_LOC_49/Y 0.44fF
C9900 INVX1_LOC_340/Y INVX1_LOC_497/Y 0.06fF
C9901 INVX1_LOC_249/A NAND2X1_LOC_123/A 0.03fF
C9902 INVX1_LOC_581/A NAND2X1_LOC_612/A 0.02fF
C9903 NAND2X1_LOC_143/a_36_24# INVX1_LOC_686/A 0.05fF
C9904 INVX1_LOC_68/Y NAND2X1_LOC_387/Y 0.02fF
C9905 VDD NAND2X1_LOC_420/Y 0.01fF
C9906 INVX1_LOC_410/Y INVX1_LOC_49/Y 0.09fF
C9907 INVX1_LOC_603/Y INVX1_LOC_600/A 0.00fF
C9908 INVX1_LOC_671/A INVX1_LOC_651/Y 0.00fF
C9909 INVX1_LOC_167/Y INVX1_LOC_54/Y 0.00fF
C9910 INVX1_LOC_31/Y INVX1_LOC_586/A 0.55fF
C9911 INVX1_LOC_268/Y INVX1_LOC_674/A 0.08fF
C9912 INVX1_LOC_20/Y INVX1_LOC_295/Y 0.03fF
C9913 INVX1_LOC_53/Y INVX1_LOC_367/Y 0.03fF
C9914 INVX1_LOC_236/A INVX1_LOC_53/Y 0.04fF
C9915 INVX1_LOC_648/Y INVX1_LOC_58/Y 0.01fF
C9916 INVX1_LOC_375/A INVX1_LOC_49/Y 0.06fF
C9917 INVX1_LOC_21/Y INVX1_LOC_160/A 0.03fF
C9918 INVX1_LOC_53/Y NAND2X1_LOC_282/a_36_24# 0.00fF
C9919 INVX1_LOC_168/A INVX1_LOC_50/Y 0.01fF
C9920 INVX1_LOC_546/A INVX1_LOC_49/Y 0.01fF
C9921 INVX1_LOC_392/Y INVX1_LOC_6/Y 0.01fF
C9922 INVX1_LOC_224/Y INVX1_LOC_245/A 0.01fF
C9923 INVX1_LOC_614/A INVX1_LOC_556/Y 0.01fF
C9924 INVX1_LOC_17/Y NAND2X1_LOC_197/a_36_24# 0.00fF
C9925 INVX1_LOC_361/Y INVX1_LOC_126/Y 0.02fF
C9926 INVX1_LOC_51/Y INVX1_LOC_69/Y 0.10fF
C9927 INVX1_LOC_607/Y INVX1_LOC_106/A 0.03fF
C9928 INVX1_LOC_213/Y INVX1_LOC_80/A 0.07fF
C9929 INVX1_LOC_586/A INVX1_LOC_641/A 0.03fF
C9930 NAND2X1_LOC_185/a_36_24# INVX1_LOC_496/A 0.00fF
C9931 INVX1_LOC_400/Y INVX1_LOC_9/Y 0.07fF
C9932 INPUT_0 NAND2X1_LOC_136/Y 0.01fF
C9933 NAND2X1_LOC_314/a_36_24# INVX1_LOC_119/Y 0.00fF
C9934 INVX1_LOC_272/Y INVX1_LOC_93/Y 0.01fF
C9935 INVX1_LOC_194/A INVX1_LOC_99/Y 0.00fF
C9936 INVX1_LOC_21/Y NAND2X1_LOC_673/B 0.01fF
C9937 INVX1_LOC_6/Y INVX1_LOC_59/A 0.03fF
C9938 INVX1_LOC_661/A INVX1_LOC_671/Y 0.21fF
C9939 INVX1_LOC_58/Y INVX1_LOC_242/A 0.03fF
C9940 INVX1_LOC_266/A INVX1_LOC_69/Y 0.12fF
C9941 INVX1_LOC_27/Y NAND2X1_LOC_84/B 0.03fF
C9942 INPUT_0 INVX1_LOC_531/Y 0.03fF
C9943 INVX1_LOC_259/A INVX1_LOC_242/Y 0.01fF
C9944 NAND2X1_LOC_387/Y INVX1_LOC_600/A 0.07fF
C9945 INVX1_LOC_367/A INVX1_LOC_6/Y 0.78fF
C9946 NAND2X1_LOC_662/a_36_24# INVX1_LOC_476/A 0.00fF
C9947 INVX1_LOC_49/Y NAND2X1_LOC_644/a_36_24# 0.01fF
C9948 INVX1_LOC_406/Y INVX1_LOC_49/Y 0.04fF
C9949 INVX1_LOC_35/Y INVX1_LOC_681/Y 0.03fF
C9950 INVX1_LOC_45/Y INVX1_LOC_26/Y 1.15fF
C9951 INVX1_LOC_160/A NAND2X1_LOC_267/A 0.05fF
C9952 INVX1_LOC_51/Y INVX1_LOC_247/Y 0.01fF
C9953 INVX1_LOC_379/A INPUT_1 0.07fF
C9954 INVX1_LOC_686/A INVX1_LOC_58/Y 0.07fF
C9955 INVX1_LOC_366/A INVX1_LOC_543/A 0.03fF
C9956 INVX1_LOC_11/Y INVX1_LOC_213/Y 1.43fF
C9957 INVX1_LOC_537/A INVX1_LOC_539/Y 0.03fF
C9958 NAND2X1_LOC_677/Y NAND2X1_LOC_647/A 0.01fF
C9959 INVX1_LOC_35/Y INPUT_1 0.20fF
C9960 NAND2X1_LOC_325/B INVX1_LOC_89/Y 0.14fF
C9961 INVX1_LOC_590/Y INVX1_LOC_531/Y 0.05fF
C9962 INVX1_LOC_400/Y INVX1_LOC_62/Y 5.09fF
C9963 INVX1_LOC_63/Y INVX1_LOC_318/Y 0.11fF
C9964 INVX1_LOC_248/Y INVX1_LOC_559/Y 0.09fF
C9965 INVX1_LOC_54/Y INVX1_LOC_137/Y 2.30fF
C9966 NAND2X1_LOC_842/a_36_24# INVX1_LOC_664/A 0.01fF
C9967 NAND2X1_LOC_190/A INVX1_LOC_413/A 0.01fF
C9968 INVX1_LOC_544/Y INVX1_LOC_80/A 0.04fF
C9969 INVX1_LOC_31/A INVX1_LOC_26/Y 0.04fF
C9970 INVX1_LOC_12/Y INVX1_LOC_486/A 0.01fF
C9971 INVX1_LOC_117/Y INVX1_LOC_432/A 0.00fF
C9972 INVX1_LOC_312/Y INVX1_LOC_682/Y 0.07fF
C9973 INVX1_LOC_44/Y INVX1_LOC_635/A 0.02fF
C9974 INVX1_LOC_669/Y INVX1_LOC_6/Y 0.02fF
C9975 INVX1_LOC_32/Y INVX1_LOC_510/A 0.12fF
C9976 INPUT_3 INVX1_LOC_26/Y 0.03fF
C9977 INVX1_LOC_44/Y NAND2X1_LOC_237/Y 0.05fF
C9978 INVX1_LOC_137/Y INVX1_LOC_611/Y 0.01fF
C9979 INVX1_LOC_80/A INVX1_LOC_662/A 0.19fF
C9980 NAND2X1_LOC_677/Y INVX1_LOC_168/Y 0.02fF
C9981 INVX1_LOC_407/Y NAND2X1_LOC_532/Y 0.05fF
C9982 INVX1_LOC_418/A INVX1_LOC_479/A 0.00fF
C9983 INVX1_LOC_316/Y NAND2X1_LOC_836/B 0.01fF
C9984 INVX1_LOC_35/Y INVX1_LOC_292/Y 0.00fF
C9985 INVX1_LOC_254/Y INVX1_LOC_46/Y 0.02fF
C9986 INVX1_LOC_367/Y NAND2X1_LOC_274/Y 0.03fF
C9987 INVX1_LOC_558/A INVX1_LOC_479/A 0.07fF
C9988 INVX1_LOC_392/A INVX1_LOC_6/Y 0.03fF
C9989 NAND2X1_LOC_39/Y INVX1_LOC_79/A 0.01fF
C9990 INVX1_LOC_68/Y INVX1_LOC_91/A 0.54fF
C9991 INVX1_LOC_276/A NAND2X1_LOC_248/B 0.00fF
C9992 NAND2X1_LOC_106/Y INVX1_LOC_118/A 0.03fF
C9993 INVX1_LOC_69/Y INVX1_LOC_40/Y 0.00fF
C9994 INVX1_LOC_366/A INVX1_LOC_86/A 0.06fF
C9995 INVX1_LOC_504/A NAND2X1_LOC_686/A 0.03fF
C9996 INVX1_LOC_93/Y INVX1_LOC_6/Y 0.19fF
C9997 INVX1_LOC_674/A INVX1_LOC_49/Y 0.07fF
C9998 INVX1_LOC_521/A INVX1_LOC_137/Y 0.03fF
C9999 INVX1_LOC_117/Y NAND2X1_LOC_542/A 0.07fF
C10000 INVX1_LOC_199/Y NAND2X1_LOC_333/B 0.01fF
C10001 INVX1_LOC_368/A INVX1_LOC_379/A 0.03fF
C10002 NAND2X1_LOC_804/a_36_24# INVX1_LOC_347/A 0.00fF
C10003 NAND2X1_LOC_184/Y INVX1_LOC_293/A 0.03fF
C10004 INVX1_LOC_58/Y INVX1_LOC_342/A 0.03fF
C10005 INVX1_LOC_53/Y NAND2X1_LOC_843/B 0.92fF
C10006 INVX1_LOC_333/Y NAND2X1_LOC_409/Y 0.04fF
C10007 NAND2X1_LOC_775/B INVX1_LOC_242/Y 0.16fF
C10008 INVX1_LOC_11/Y INVX1_LOC_653/A 0.02fF
C10009 INVX1_LOC_309/Y INVX1_LOC_46/Y 0.01fF
C10010 NAND2X1_LOC_844/a_36_24# INVX1_LOC_367/Y 0.01fF
C10011 INVX1_LOC_227/Y INVX1_LOC_245/A 0.01fF
C10012 INVX1_LOC_537/A INVX1_LOC_62/Y 0.07fF
C10013 INVX1_LOC_292/Y INVX1_LOC_621/Y 0.00fF
C10014 INVX1_LOC_513/A INVX1_LOC_79/A 0.03fF
C10015 INVX1_LOC_84/Y INVX1_LOC_9/Y 0.16fF
C10016 INVX1_LOC_53/Y INVX1_LOC_91/Y 0.05fF
C10017 NAND2X1_LOC_334/B INVX1_LOC_6/Y 0.03fF
C10018 INVX1_LOC_643/Y INVX1_LOC_6/Y 0.01fF
C10019 INVX1_LOC_298/A INVX1_LOC_531/Y 0.01fF
C10020 INVX1_LOC_179/A INVX1_LOC_361/A 0.02fF
C10021 INVX1_LOC_6/Y NAND2X1_LOC_624/a_36_24# 0.00fF
C10022 INVX1_LOC_254/Y INVX1_LOC_75/A 0.05fF
C10023 INVX1_LOC_508/A INVX1_LOC_655/A 0.11fF
C10024 INVX1_LOC_62/Y INVX1_LOC_496/Y 0.03fF
C10025 INVX1_LOC_63/Y INVX1_LOC_90/Y 0.08fF
C10026 NAND2X1_LOC_294/Y NAND2X1_LOC_401/a_36_24# 0.01fF
C10027 INVX1_LOC_298/A INVX1_LOC_528/Y 0.01fF
C10028 INVX1_LOC_479/A INVX1_LOC_46/Y 0.36fF
C10029 INVX1_LOC_58/Y NAND2X1_LOC_609/B 0.03fF
C10030 NAND2X1_LOC_433/Y INVX1_LOC_653/A 0.09fF
C10031 INVX1_LOC_338/Y INVX1_LOC_588/A 0.51fF
C10032 NAND2X1_LOC_274/B INVX1_LOC_468/A 0.01fF
C10033 INVX1_LOC_426/A INVX1_LOC_586/A 0.01fF
C10034 INVX1_LOC_112/Y INVX1_LOC_41/Y 0.03fF
C10035 NAND2X1_LOC_249/Y INVX1_LOC_45/Y 0.03fF
C10036 INVX1_LOC_20/Y NAND2X1_LOC_99/a_36_24# 0.00fF
C10037 NAND2X1_LOC_335/B INVX1_LOC_269/A 0.09fF
C10038 VDD GATE_741 0.15fF
C10039 INVX1_LOC_442/Y INVX1_LOC_109/Y 0.07fF
C10040 INVX1_LOC_195/A INVX1_LOC_85/Y 0.01fF
C10041 INVX1_LOC_531/Y INVX1_LOC_211/A 0.07fF
C10042 INVX1_LOC_426/A INVX1_LOC_312/Y 0.46fF
C10043 NAND2X1_LOC_475/A INVX1_LOC_482/A 0.02fF
C10044 INVX1_LOC_410/Y INVX1_LOC_76/Y 0.14fF
C10045 INVX1_LOC_479/A INVX1_LOC_75/A 0.04fF
C10046 INPUT_0 NAND2X1_LOC_467/A 0.22fF
C10047 INVX1_LOC_12/Y INVX1_LOC_596/Y 0.00fF
C10048 INVX1_LOC_7/A INVX1_LOC_7/Y 0.01fF
C10049 INVX1_LOC_405/A INVX1_LOC_235/A 0.01fF
C10050 NAND2X1_LOC_331/B INVX1_LOC_495/A 0.50fF
C10051 VDD INVX1_LOC_310/Y 0.36fF
C10052 VDD INVX1_LOC_565/A 0.00fF
C10053 INVX1_LOC_20/Y INVX1_LOC_271/A 0.28fF
C10054 INVX1_LOC_51/Y INVX1_LOC_586/A 0.40fF
C10055 INVX1_LOC_272/Y INVX1_LOC_395/A 0.02fF
C10056 INVX1_LOC_395/A NAND2X1_LOC_820/A 0.03fF
C10057 INVX1_LOC_74/Y NAND2X1_LOC_418/a_36_24# 0.00fF
C10058 NAND2X1_LOC_234/Y INVX1_LOC_619/Y 0.00fF
C10059 INVX1_LOC_20/Y INVX1_LOC_173/A 0.30fF
C10060 INVX1_LOC_145/A INVX1_LOC_41/A 0.02fF
C10061 INVX1_LOC_301/A NAND2X1_LOC_775/B 0.49fF
C10062 INVX1_LOC_266/A INVX1_LOC_586/A 0.11fF
C10063 INVX1_LOC_137/A INVX1_LOC_492/Y 0.00fF
C10064 NAND2X1_LOC_836/B NAND2X1_LOC_31/a_36_24# 0.01fF
C10065 NAND2X1_LOC_475/A INVX1_LOC_194/A 0.02fF
C10066 INVX1_LOC_416/Y INVX1_LOC_12/Y 0.02fF
C10067 INVX1_LOC_312/Y INVX1_LOC_51/Y 0.07fF
C10068 INVX1_LOC_45/Y INVX1_LOC_369/A 0.03fF
C10069 INVX1_LOC_395/A INVX1_LOC_252/A 0.01fF
C10070 INVX1_LOC_65/Y NAND2X1_LOC_318/B 0.02fF
C10071 INVX1_LOC_206/Y NAND2X1_LOC_672/a_36_24# 0.00fF
C10072 INVX1_LOC_300/A INVX1_LOC_271/A 0.03fF
C10073 INVX1_LOC_122/Y INVX1_LOC_105/A 0.01fF
C10074 INVX1_LOC_585/Y NAND2X1_LOC_749/Y 0.00fF
C10075 INVX1_LOC_271/A INVX1_LOC_197/Y 0.07fF
C10076 NAND2X1_LOC_176/a_36_24# NAND2X1_LOC_307/A 0.01fF
C10077 NAND2X1_LOC_45/Y NAND2X1_LOC_190/a_36_24# 0.01fF
C10078 INVX1_LOC_45/Y NAND2X1_LOC_275/Y 1.47fF
C10079 NAND2X1_LOC_498/Y INVX1_LOC_303/Y 0.10fF
C10080 INVX1_LOC_412/Y INVX1_LOC_32/Y 0.06fF
C10081 INVX1_LOC_65/Y INVX1_LOC_177/A 0.11fF
C10082 VDD NAND2X1_LOC_586/Y 0.01fF
C10083 INVX1_LOC_84/A NAND2X1_LOC_48/Y 0.02fF
C10084 NAND2X1_LOC_97/A INVX1_LOC_59/Y 0.01fF
C10085 INVX1_LOC_432/Y NAND2X1_LOC_383/Y 0.33fF
C10086 INVX1_LOC_150/Y INVX1_LOC_137/Y 0.05fF
C10087 NAND2X1_LOC_299/Y INVX1_LOC_197/A 0.07fF
C10088 INVX1_LOC_510/Y NAND2X1_LOC_307/a_36_24# 0.00fF
C10089 INVX1_LOC_80/A NAND2X1_LOC_147/a_36_24# 0.00fF
C10090 INVX1_LOC_500/Y INVX1_LOC_586/A 0.01fF
C10091 INVX1_LOC_84/A INVX1_LOC_47/A 0.03fF
C10092 INVX1_LOC_406/Y INVX1_LOC_386/Y 0.03fF
C10093 INVX1_LOC_588/Y INVX1_LOC_288/A 0.07fF
C10094 INVX1_LOC_273/A NAND2X1_LOC_226/a_36_24# 0.00fF
C10095 INVX1_LOC_37/Y INVX1_LOC_6/Y 0.01fF
C10096 INVX1_LOC_313/Y NAND2X1_LOC_383/Y 0.09fF
C10097 INVX1_LOC_570/Y NAND2X1_LOC_846/B 0.10fF
C10098 INVX1_LOC_449/Y INVX1_LOC_384/A 0.02fF
C10099 INVX1_LOC_366/A NAND2X1_LOC_223/a_36_24# 0.00fF
C10100 INVX1_LOC_395/A INVX1_LOC_6/Y 0.37fF
C10101 NAND2X1_LOC_780/B INVX1_LOC_168/Y 0.02fF
C10102 INVX1_LOC_54/Y NAND2X1_LOC_29/a_36_24# 0.00fF
C10103 NAND2X1_LOC_543/B INVX1_LOC_114/A 0.03fF
C10104 INVX1_LOC_365/Y NAND2X1_LOC_378/Y 0.01fF
C10105 INVX1_LOC_137/A NAND2X1_LOC_647/A 0.17fF
C10106 INVX1_LOC_206/Y NAND2X1_LOC_440/A 0.05fF
C10107 INPUT_2 NAND2X1_LOC_84/B 0.01fF
C10108 INVX1_LOC_292/A INVX1_LOC_44/Y 0.06fF
C10109 NAND2X1_LOC_391/A INVX1_LOC_230/A 0.08fF
C10110 INVX1_LOC_596/A INVX1_LOC_370/A 0.12fF
C10111 INVX1_LOC_551/Y NAND2X1_LOC_615/B 0.01fF
C10112 INVX1_LOC_362/Y INVX1_LOC_6/Y 0.07fF
C10113 NAND2X1_LOC_108/Y INVX1_LOC_69/Y 0.01fF
C10114 INVX1_LOC_237/Y INVX1_LOC_212/Y 0.01fF
C10115 INVX1_LOC_409/A NAND2X1_LOC_274/B 0.01fF
C10116 INVX1_LOC_384/A NAND2X1_LOC_849/a_36_24# 0.01fF
C10117 NAND2X1_LOC_177/a_36_24# NAND2X1_LOC_444/A 0.00fF
C10118 INVX1_LOC_206/Y INVX1_LOC_245/A 0.21fF
C10119 INVX1_LOC_106/A INVX1_LOC_145/Y 0.01fF
C10120 INVX1_LOC_214/Y INVX1_LOC_679/Y 0.02fF
C10121 INVX1_LOC_211/Y INVX1_LOC_12/Y 0.07fF
C10122 INVX1_LOC_248/Y INVX1_LOC_155/Y 0.00fF
C10123 NAND2X1_LOC_136/a_36_24# INVX1_LOC_6/Y 0.00fF
C10124 INVX1_LOC_617/Y INVX1_LOC_32/Y 0.03fF
C10125 INVX1_LOC_176/Y INVX1_LOC_32/Y 0.02fF
C10126 NAND2X1_LOC_396/a_36_24# INVX1_LOC_245/A 0.01fF
C10127 INVX1_LOC_295/A INVX1_LOC_117/Y 0.03fF
C10128 INVX1_LOC_54/Y NAND2X1_LOC_307/A 0.25fF
C10129 INVX1_LOC_137/Y NAND2X1_LOC_677/Y 0.59fF
C10130 INVX1_LOC_210/Y INVX1_LOC_21/Y 0.00fF
C10131 INVX1_LOC_58/Y INVX1_LOC_94/A 0.05fF
C10132 NAND2X1_LOC_498/Y INVX1_LOC_9/Y 0.07fF
C10133 NAND2X1_LOC_638/A INVX1_LOC_259/Y 0.03fF
C10134 INVX1_LOC_53/Y INVX1_LOC_361/Y 0.03fF
C10135 INVX1_LOC_570/A INVX1_LOC_9/Y 0.06fF
C10136 INVX1_LOC_551/Y INVX1_LOC_66/A 0.03fF
C10137 INVX1_LOC_291/A INVX1_LOC_292/Y 0.00fF
C10138 INVX1_LOC_17/Y INVX1_LOC_176/A 1.23fF
C10139 INVX1_LOC_133/A NAND2X1_LOC_286/A 0.03fF
C10140 INVX1_LOC_683/Y INVX1_LOC_6/Y 0.01fF
C10141 NAND2X1_LOC_45/Y INVX1_LOC_62/Y 2.06fF
C10142 INPUT_0 INVX1_LOC_41/Y 1.22fF
C10143 NAND2X1_LOC_327/a_36_24# INVX1_LOC_353/A 0.01fF
C10144 INVX1_LOC_12/Y INVX1_LOC_46/Y 0.20fF
C10145 INVX1_LOC_318/A NAND2X1_LOC_318/B 0.24fF
C10146 INVX1_LOC_561/A INVX1_LOC_579/Y 0.00fF
C10147 INVX1_LOC_35/Y NAND2X1_LOC_465/a_36_24# 0.00fF
C10148 NAND2X1_LOC_545/B INVX1_LOC_253/Y 0.03fF
C10149 INVX1_LOC_587/Y INVX1_LOC_99/Y 0.48fF
C10150 INVX1_LOC_53/Y INVX1_LOC_261/Y 0.03fF
C10151 INVX1_LOC_338/A INPUT_1 0.05fF
C10152 INVX1_LOC_448/A NAND2X1_LOC_849/a_36_24# 0.00fF
C10153 INVX1_LOC_257/A INVX1_LOC_545/Y -0.05fF
C10154 INVX1_LOC_254/Y INVX1_LOC_202/Y 0.02fF
C10155 INVX1_LOC_379/A INVX1_LOC_50/Y 0.07fF
C10156 NAND2X1_LOC_538/a_36_24# INVX1_LOC_98/Y 0.00fF
C10157 INVX1_LOC_418/Y INVX1_LOC_159/Y 0.01fF
C10158 INVX1_LOC_140/Y INVX1_LOC_473/Y 0.29fF
C10159 GATE_865 INVX1_LOC_685/Y 0.14fF
C10160 INVX1_LOC_45/Y NAND2X1_LOC_626/Y 0.04fF
C10161 INVX1_LOC_17/Y INVX1_LOC_354/Y 0.01fF
C10162 NAND2X1_LOC_516/Y INVX1_LOC_41/Y 0.03fF
C10163 INVX1_LOC_35/Y INVX1_LOC_50/Y 0.21fF
C10164 NAND2X1_LOC_333/A NAND2X1_LOC_755/B 0.00fF
C10165 INVX1_LOC_548/Y INVX1_LOC_479/A 0.05fF
C10166 INVX1_LOC_455/Y NAND2X1_LOC_836/B 0.01fF
C10167 INVX1_LOC_134/Y INVX1_LOC_496/A 0.13fF
C10168 INVX1_LOC_419/Y INVX1_LOC_54/Y 0.00fF
C10169 INVX1_LOC_570/A INVX1_LOC_62/Y 0.03fF
C10170 NAND2X1_LOC_184/Y NAND2X1_LOC_106/B 0.06fF
C10171 NAND2X1_LOC_391/B INVX1_LOC_79/A 0.00fF
C10172 INVX1_LOC_6/A INVX1_LOC_18/Y 0.00fF
C10173 NAND2X1_LOC_389/a_36_24# INVX1_LOC_35/Y 0.00fF
C10174 INVX1_LOC_686/A INVX1_LOC_245/A 0.07fF
C10175 INVX1_LOC_293/Y INVX1_LOC_26/Y 0.06fF
C10176 NAND2X1_LOC_516/B INVX1_LOC_100/Y 0.05fF
C10177 INVX1_LOC_131/A INVX1_LOC_662/A 0.03fF
C10178 INVX1_LOC_54/Y NAND2X1_LOC_747/a_36_24# 0.00fF
C10179 NAND2X1_LOC_56/Y NAND2X1_LOC_845/B 0.00fF
C10180 INVX1_LOC_548/A INVX1_LOC_6/Y 0.58fF
C10181 INVX1_LOC_89/Y INVX1_LOC_137/Y 0.06fF
C10182 INVX1_LOC_17/Y INVX1_LOC_410/A 0.03fF
C10183 INVX1_LOC_551/Y NAND2X1_LOC_601/Y 0.47fF
C10184 INVX1_LOC_267/A NAND2X1_LOC_720/A 0.04fF
C10185 INVX1_LOC_138/Y INVX1_LOC_46/Y 0.01fF
C10186 INVX1_LOC_17/Y INVX1_LOC_170/Y 0.01fF
C10187 INVX1_LOC_63/Y INVX1_LOC_98/Y 0.07fF
C10188 NAND2X1_LOC_260/a_36_24# INVX1_LOC_283/A 0.00fF
C10189 INVX1_LOC_38/A INVX1_LOC_39/Y 0.18fF
C10190 INVX1_LOC_50/Y INVX1_LOC_620/A 0.10fF
C10191 INVX1_LOC_11/Y NAND2X1_LOC_258/Y 0.01fF
C10192 INVX1_LOC_183/A NAND2X1_LOC_621/a_36_24# 0.01fF
C10193 NAND2X1_LOC_318/A INVX1_LOC_479/A 0.03fF
C10194 INVX1_LOC_99/Y INVX1_LOC_9/Y 0.17fF
C10195 NAND2X1_LOC_274/B INVX1_LOC_377/A 0.01fF
C10196 INVX1_LOC_338/Y NAND2X1_LOC_646/A 0.03fF
C10197 INVX1_LOC_47/Y INVX1_LOC_539/Y 0.04fF
C10198 NAND2X1_LOC_274/B NAND2X1_LOC_595/Y 0.02fF
C10199 INVX1_LOC_31/Y INVX1_LOC_6/Y 0.30fF
C10200 INVX1_LOC_402/Y INVX1_LOC_100/Y 0.03fF
C10201 NAND2X1_LOC_532/Y NAND2X1_LOC_308/A 0.73fF
C10202 NAND2X1_LOC_301/B INVX1_LOC_116/Y 0.03fF
C10203 NAND2X1_LOC_148/A NAND2X1_LOC_843/B 0.45fF
C10204 INVX1_LOC_166/Y INVX1_LOC_99/Y 0.00fF
C10205 NAND2X1_LOC_274/B INVX1_LOC_352/Y 0.01fF
C10206 NAND2X1_LOC_107/Y NAND2X1_LOC_843/B 0.10fF
C10207 NAND2X1_LOC_673/B INVX1_LOC_26/Y 0.01fF
C10208 INVX1_LOC_80/A INVX1_LOC_666/Y 0.10fF
C10209 INVX1_LOC_501/A INVX1_LOC_355/Y 0.12fF
C10210 INVX1_LOC_531/Y INVX1_LOC_145/Y 0.12fF
C10211 INVX1_LOC_257/A NAND2X1_LOC_325/a_36_24# 0.00fF
C10212 INVX1_LOC_668/Y INVX1_LOC_669/A 0.14fF
C10213 INVX1_LOC_62/Y INVX1_LOC_99/Y 0.19fF
C10214 GATE_662 NAND2X1_LOC_847/A 0.06fF
C10215 INVX1_LOC_123/A INVX1_LOC_9/Y 0.04fF
C10216 INVX1_LOC_69/Y INVX1_LOC_361/A 0.03fF
C10217 INVX1_LOC_54/Y INVX1_LOC_502/A 0.10fF
C10218 NAND2X1_LOC_315/a_36_24# INVX1_LOC_92/A 0.00fF
C10219 INVX1_LOC_568/A INVX1_LOC_9/Y 0.01fF
C10220 INVX1_LOC_504/A INVX1_LOC_588/A 0.32fF
C10221 INVX1_LOC_99/Y NAND2X1_LOC_844/A 0.05fF
C10222 INVX1_LOC_6/Y NAND2X1_LOC_623/a_36_24# 0.00fF
C10223 INVX1_LOC_317/A INVX1_LOC_242/Y 0.04fF
C10224 INVX1_LOC_63/Y INVX1_LOC_338/Y 0.07fF
C10225 INVX1_LOC_309/Y INVX1_LOC_49/Y 0.05fF
C10226 INVX1_LOC_11/Y INVX1_LOC_653/Y 0.08fF
C10227 INVX1_LOC_47/Y INVX1_LOC_9/Y 3.82fF
C10228 INVX1_LOC_202/Y INVX1_LOC_479/A 0.16fF
C10229 NAND2X1_LOC_557/B INVX1_LOC_9/Y 0.78fF
C10230 INVX1_LOC_573/Y NAND2X1_LOC_679/A 0.09fF
C10231 INVX1_LOC_213/Y NAND2X1_LOC_843/B 0.02fF
C10232 INVX1_LOC_298/A INVX1_LOC_41/Y 0.03fF
C10233 INVX1_LOC_58/Y INVX1_LOC_376/Y 0.07fF
C10234 NAND2X1_LOC_334/A INVX1_LOC_245/A 0.03fF
C10235 INVX1_LOC_41/Y INVX1_LOC_498/A 5.38fF
C10236 INVX1_LOC_681/Y INVX1_LOC_364/A 0.05fF
C10237 INVX1_LOC_133/Y INVX1_LOC_626/Y 0.01fF
C10238 INVX1_LOC_47/Y INVX1_LOC_166/Y 0.02fF
C10239 INVX1_LOC_47/Y INVX1_LOC_62/Y 0.22fF
C10240 NAND2X1_LOC_410/Y INVX1_LOC_66/A 0.01fF
C10241 INPUT_1 INVX1_LOC_488/Y 0.01fF
C10242 INVX1_LOC_261/Y NAND2X1_LOC_451/B 0.03fF
C10243 NAND2X1_LOC_66/Y INVX1_LOC_9/Y 0.07fF
C10244 INVX1_LOC_46/Y INVX1_LOC_212/A 0.01fF
C10245 INVX1_LOC_49/Y INVX1_LOC_479/A 0.46fF
C10246 INVX1_LOC_166/Y INVX1_LOC_119/Y 0.01fF
C10247 NAND2X1_LOC_69/B INVX1_LOC_72/Y 0.22fF
C10248 NAND2X1_LOC_790/B INVX1_LOC_45/Y 0.09fF
C10249 INVX1_LOC_380/A INVX1_LOC_20/Y 0.01fF
C10250 INVX1_LOC_93/Y INVX1_LOC_636/A 0.08fF
C10251 NAND2X1_LOC_336/B INVX1_LOC_109/Y 0.00fF
C10252 INVX1_LOC_567/A INVX1_LOC_51/Y 0.00fF
C10253 INVX1_LOC_62/Y INVX1_LOC_119/Y 0.07fF
C10254 NAND2X1_LOC_274/B NAND2X1_LOC_372/Y 0.03fF
C10255 NAND2X1_LOC_433/Y INVX1_LOC_653/Y 0.00fF
C10256 NAND2X1_LOC_7/Y INVX1_LOC_169/A 0.00fF
C10257 INVX1_LOC_239/Y INVX1_LOC_132/Y 0.03fF
C10258 NAND2X1_LOC_537/A INVX1_LOC_586/A 0.01fF
C10259 NAND2X1_LOC_206/a_36_24# INVX1_LOC_395/A 0.00fF
C10260 INVX1_LOC_41/Y INVX1_LOC_211/A 0.07fF
C10261 INVX1_LOC_103/A INVX1_LOC_45/Y 0.03fF
C10262 NAND2X1_LOC_249/Y INVX1_LOC_293/Y 0.00fF
C10263 INVX1_LOC_41/Y INVX1_LOC_64/Y 0.65fF
C10264 INVX1_LOC_344/Y INVX1_LOC_638/A -0.05fF
C10265 INVX1_LOC_79/A NAND2X1_LOC_418/a_36_24# 0.01fF
C10266 INVX1_LOC_160/Y INVX1_LOC_286/A 0.01fF
C10267 INVX1_LOC_35/Y INVX1_LOC_275/A 0.02fF
C10268 INVX1_LOC_626/Y INVX1_LOC_581/A 0.01fF
C10269 INVX1_LOC_51/Y INVX1_LOC_366/A 0.00fF
C10270 INVX1_LOC_442/A INVX1_LOC_551/Y 0.03fF
C10271 INVX1_LOC_523/A INVX1_LOC_508/Y 0.02fF
C10272 INVX1_LOC_45/Y INVX1_LOC_235/Y 0.07fF
C10273 NAND2X1_LOC_13/Y INVX1_LOC_586/A 0.03fF
C10274 INPUT_0 INVX1_LOC_358/Y 0.04fF
C10275 INVX1_LOC_312/Y INVX1_LOC_216/Y 0.01fF
C10276 INVX1_LOC_335/Y INPUT_0 0.12fF
C10277 NAND2X1_LOC_373/Y NAND2X1_LOC_775/B 0.04fF
C10278 NAND2X1_LOC_93/Y INVX1_LOC_35/Y 0.08fF
C10279 INVX1_LOC_438/A INVX1_LOC_379/A 1.21fF
C10280 INVX1_LOC_435/Y INVX1_LOC_434/Y 0.05fF
C10281 INVX1_LOC_628/Y INVX1_LOC_629/Y 0.13fF
C10282 INPUT_0 INVX1_LOC_21/Y 2.48fF
C10283 VDD INVX1_LOC_595/Y 0.29fF
C10284 INVX1_LOC_300/A INVX1_LOC_562/A 0.03fF
C10285 VDD INVX1_LOC_304/Y 0.70fF
C10286 INVX1_LOC_272/Y INVX1_LOC_51/Y 3.79fF
C10287 NAND2X1_LOC_791/B INVX1_LOC_51/Y 0.07fF
C10288 NAND2X1_LOC_744/a_36_24# INVX1_LOC_549/Y 0.00fF
C10289 INVX1_LOC_438/A INVX1_LOC_35/Y 0.07fF
C10290 INVX1_LOC_560/A INVX1_LOC_160/A 0.15fF
C10291 INVX1_LOC_51/Y INVX1_LOC_486/Y 0.01fF
C10292 NAND2X1_LOC_780/B INVX1_LOC_137/Y 0.06fF
C10293 INVX1_LOC_619/Y INVX1_LOC_623/A 0.00fF
C10294 INVX1_LOC_530/Y INVX1_LOC_12/Y 0.15fF
C10295 INVX1_LOC_162/Y INVX1_LOC_161/A 0.00fF
C10296 INVX1_LOC_160/Y NAND2X1_LOC_123/A 0.03fF
C10297 INVX1_LOC_52/Y INPUT_1 0.01fF
C10298 INVX1_LOC_11/Y INVX1_LOC_490/Y 0.23fF
C10299 INVX1_LOC_20/Y INVX1_LOC_581/A 0.15fF
C10300 NAND2X1_LOC_318/A INVX1_LOC_12/Y 0.01fF
C10301 NAND2X1_LOC_93/Y INVX1_LOC_620/A 0.01fF
C10302 INVX1_LOC_435/Y NAND2X1_LOC_250/Y 0.05fF
C10303 INVX1_LOC_580/Y INVX1_LOC_99/Y 0.09fF
C10304 INVX1_LOC_580/A INVX1_LOC_145/Y 0.09fF
C10305 INVX1_LOC_312/Y NAND2X1_LOC_768/a_36_24# 0.01fF
C10306 NAND2X1_LOC_32/Y INVX1_LOC_395/A -0.07fF
C10307 INVX1_LOC_11/Y NAND2X1_LOC_16/Y 0.03fF
C10308 INVX1_LOC_137/A INVX1_LOC_137/Y 0.14fF
C10309 INVX1_LOC_607/A NAND2X1_LOC_106/B 0.02fF
C10310 INVX1_LOC_556/Y INVX1_LOC_45/Y 0.03fF
C10311 INPUT_3 NAND2X1_LOC_19/a_36_24# 0.00fF
C10312 NAND2X1_LOC_475/A INVX1_LOC_155/A 0.01fF
C10313 INVX1_LOC_21/Y INVX1_LOC_586/Y 0.01fF
C10314 INVX1_LOC_133/Y INVX1_LOC_655/A 0.01fF
C10315 INVX1_LOC_406/Y INVX1_LOC_7/Y 0.00fF
C10316 INVX1_LOC_551/Y INVX1_LOC_116/Y 0.10fF
C10317 INVX1_LOC_519/A INVX1_LOC_383/Y 0.02fF
C10318 INVX1_LOC_502/Y INVX1_LOC_303/Y 0.01fF
C10319 VDD INVX1_LOC_183/A 0.06fF
C10320 INVX1_LOC_276/A INVX1_LOC_662/Y 0.10fF
C10321 INVX1_LOC_17/Y NAND2X1_LOC_176/a_36_24# 0.01fF
C10322 INVX1_LOC_254/Y INVX1_LOC_76/Y 0.03fF
C10323 INVX1_LOC_286/A NAND2X1_LOC_267/A 0.13fF
C10324 INVX1_LOC_239/Y INVX1_LOC_655/A 0.02fF
C10325 INVX1_LOC_409/Y INVX1_LOC_114/A 0.05fF
C10326 INVX1_LOC_298/A INVX1_LOC_315/Y 0.01fF
C10327 NAND2X1_LOC_391/B INVX1_LOC_48/Y 0.01fF
C10328 INVX1_LOC_442/Y INVX1_LOC_53/Y 0.07fF
C10329 INVX1_LOC_412/A INVX1_LOC_199/Y 0.91fF
C10330 VDD INVX1_LOC_389/Y 0.21fF
C10331 INVX1_LOC_605/A NAND2X1_LOC_307/B 0.00fF
C10332 NAND2X1_LOC_150/a_36_24# INVX1_LOC_46/Y 0.01fF
C10333 INVX1_LOC_44/Y NAND2X1_LOC_749/Y 2.52fF
C10334 NAND2X1_LOC_475/A INVX1_LOC_9/Y 0.05fF
C10335 INVX1_LOC_166/A NAND2X1_LOC_332/B 0.07fF
C10336 INVX1_LOC_291/A INVX1_LOC_50/Y 0.17fF
C10337 INVX1_LOC_558/A INVX1_LOC_66/A 0.01fF
C10338 NAND2X1_LOC_635/a_36_24# INVX1_LOC_505/A 0.00fF
C10339 INVX1_LOC_512/Y NAND2X1_LOC_829/B 0.16fF
C10340 NAND2X1_LOC_498/Y INVX1_LOC_624/Y 0.02fF
C10341 INVX1_LOC_51/Y INVX1_LOC_6/Y 0.07fF
C10342 INVX1_LOC_435/Y INVX1_LOC_63/Y 0.05fF
C10343 INVX1_LOC_381/A INVX1_LOC_93/Y 0.07fF
C10344 INVX1_LOC_35/Y NAND2X1_LOC_513/A 0.03fF
C10345 INVX1_LOC_626/A NAND2X1_LOC_796/a_36_24# 0.00fF
C10346 INVX1_LOC_168/A INVX1_LOC_117/Y 0.03fF
C10347 INVX1_LOC_570/A INVX1_LOC_624/Y 0.00fF
C10348 NAND2X1_LOC_673/B INVX1_LOC_369/A 0.07fF
C10349 NAND2X1_LOC_142/Y INVX1_LOC_58/Y 0.01fF
C10350 INVX1_LOC_21/Y INVX1_LOC_201/A 0.00fF
C10351 INVX1_LOC_202/Y INVX1_LOC_12/Y 1.30fF
C10352 NAND2X1_LOC_333/A INVX1_LOC_268/Y 0.16fF
C10353 INVX1_LOC_580/Y INVX1_LOC_47/Y 0.03fF
C10354 INVX1_LOC_266/Y INVX1_LOC_77/Y 0.26fF
C10355 INVX1_LOC_20/Y INVX1_LOC_317/A 0.03fF
C10356 INVX1_LOC_395/A INVX1_LOC_557/Y 0.01fF
C10357 NAND2X1_LOC_111/Y NAND2X1_LOC_332/B 0.10fF
C10358 INVX1_LOC_193/A INVX1_LOC_134/Y 0.02fF
C10359 INVX1_LOC_447/Y INVX1_LOC_17/Y 0.01fF
C10360 INVX1_LOC_586/A NAND2X1_LOC_668/Y 0.01fF
C10361 NAND2X1_LOC_475/A INVX1_LOC_62/Y 0.06fF
C10362 INVX1_LOC_520/Y INVX1_LOC_242/A 0.01fF
C10363 INVX1_LOC_672/Y INVX1_LOC_679/A 0.14fF
C10364 INVX1_LOC_257/Y INVX1_LOC_41/Y 0.07fF
C10365 INVX1_LOC_551/Y INVX1_LOC_255/A 0.12fF
C10366 INVX1_LOC_45/Y NAND2X1_LOC_420/Y 0.02fF
C10367 INVX1_LOC_160/A INVX1_LOC_603/A 0.40fF
C10368 INVX1_LOC_206/Y NAND2X1_LOC_597/Y 0.05fF
C10369 INVX1_LOC_358/Y INVX1_LOC_498/A 0.03fF
C10370 INVX1_LOC_335/Y INVX1_LOC_298/A 0.03fF
C10371 INVX1_LOC_545/Y INVX1_LOC_89/Y 0.02fF
C10372 GATE_865 INVX1_LOC_631/A 0.05fF
C10373 NAND2X1_LOC_530/a_36_24# INVX1_LOC_6/Y 0.00fF
C10374 NAND2X1_LOC_307/A INVX1_LOC_89/Y 0.14fF
C10375 NAND2X1_LOC_123/A NAND2X1_LOC_267/A 0.07fF
C10376 INVX1_LOC_604/Y INVX1_LOC_208/Y 0.04fF
C10377 NAND2X1_LOC_664/a_36_24# INVX1_LOC_50/Y 0.00fF
C10378 INVX1_LOC_384/A INVX1_LOC_301/Y 0.07fF
C10379 NAND2X1_LOC_336/B INVX1_LOC_199/Y 0.03fF
C10380 INVX1_LOC_338/A INVX1_LOC_50/Y 0.01fF
C10381 NAND2X1_LOC_532/Y INVX1_LOC_134/Y 0.05fF
C10382 INVX1_LOC_17/Y INVX1_LOC_54/Y 1.93fF
C10383 INVX1_LOC_549/Y INVX1_LOC_186/Y 0.02fF
C10384 INVX1_LOC_372/Y INVX1_LOC_49/Y 0.00fF
C10385 INPUT_0 INVX1_LOC_209/Y 0.07fF
C10386 INVX1_LOC_446/Y INVX1_LOC_41/Y 0.02fF
C10387 NAND2X1_LOC_142/Y NAND2X1_LOC_342/B 0.34fF
C10388 INVX1_LOC_596/A INVX1_LOC_63/Y 0.01fF
C10389 INVX1_LOC_392/Y INVX1_LOC_100/Y 0.01fF
C10390 INVX1_LOC_21/Y INVX1_LOC_83/A 0.00fF
C10391 INPUT_1 INVX1_LOC_350/A 0.01fF
C10392 NAND2X1_LOC_837/B INVX1_LOC_50/Y 0.10fF
C10393 INVX1_LOC_300/A INVX1_LOC_317/A 0.03fF
C10394 INVX1_LOC_288/A INVX1_LOC_41/Y 0.07fF
C10395 NAND2X1_LOC_409/a_36_24# INVX1_LOC_93/A 0.00fF
C10396 INVX1_LOC_442/Y NAND2X1_LOC_346/B 0.07fF
C10397 INVX1_LOC_12/Y INVX1_LOC_49/Y 0.22fF
C10398 INVX1_LOC_319/Y INVX1_LOC_666/Y 0.01fF
C10399 INVX1_LOC_58/Y INVX1_LOC_676/A 0.01fF
C10400 INVX1_LOC_35/Y NAND2X1_LOC_63/a_36_24# 0.00fF
C10401 NAND2X1_LOC_318/B INVX1_LOC_63/Y 0.02fF
C10402 NAND2X1_LOC_137/A NAND2X1_LOC_859/a_36_24# 0.00fF
C10403 NAND2X1_LOC_498/B INVX1_LOC_479/A 0.01fF
C10404 INVX1_LOC_442/Y NAND2X1_LOC_274/Y 0.01fF
C10405 INVX1_LOC_93/Y NAND2X1_LOC_720/A 0.07fF
C10406 INVX1_LOC_84/A INVX1_LOC_90/Y 0.08fF
C10407 NAND2X1_LOC_388/A INVX1_LOC_35/Y 0.00fF
C10408 INVX1_LOC_674/A INVX1_LOC_32/Y 0.12fF
C10409 INVX1_LOC_416/A INVX1_LOC_89/Y 0.03fF
C10410 INVX1_LOC_136/Y INVX1_LOC_9/Y 0.06fF
C10411 INVX1_LOC_384/A INVX1_LOC_41/Y 0.61fF
C10412 INVX1_LOC_12/Y INVX1_LOC_642/Y 0.01fF
C10413 NAND2X1_LOC_615/B INVX1_LOC_46/Y 0.05fF
C10414 INVX1_LOC_448/A INVX1_LOC_301/Y 0.07fF
C10415 INVX1_LOC_504/A INVX1_LOC_63/Y 0.08fF
C10416 INVX1_LOC_444/Y NAND2X1_LOC_344/B 0.00fF
C10417 NAND2X1_LOC_172/a_36_24# INVX1_LOC_561/A 0.00fF
C10418 INVX1_LOC_117/Y NAND2X1_LOC_619/Y 0.07fF
C10419 INVX1_LOC_211/Y INVX1_LOC_296/A 0.00fF
C10420 INVX1_LOC_367/A INVX1_LOC_100/Y 0.07fF
C10421 INVX1_LOC_581/A INVX1_LOC_655/A -0.03fF
C10422 INVX1_LOC_607/Y INVX1_LOC_107/Y 0.04fF
C10423 INVX1_LOC_490/Y INVX1_LOC_231/Y 0.00fF
C10424 INVX1_LOC_449/A NAND2X1_LOC_274/B 0.03fF
C10425 INVX1_LOC_76/Y INVX1_LOC_479/A 0.15fF
C10426 NAND2X1_LOC_152/a_36_24# INVX1_LOC_655/A 0.01fF
C10427 INVX1_LOC_442/A INVX1_LOC_634/Y 0.49fF
C10428 INVX1_LOC_177/A INVX1_LOC_63/Y 0.01fF
C10429 INVX1_LOC_556/Y INVX1_LOC_89/A 0.01fF
C10430 INVX1_LOC_93/Y NAND2X1_LOC_200/a_36_24# 0.00fF
C10431 INVX1_LOC_660/A INVX1_LOC_59/A 0.01fF
C10432 NAND2X1_LOC_43/Y INVX1_LOC_9/Y 0.01fF
C10433 INVX1_LOC_46/Y INVX1_LOC_66/A 0.08fF
C10434 NAND2X1_LOC_106/Y NAND2X1_LOC_115/a_36_24# 0.00fF
C10435 NAND2X1_LOC_521/Y INVX1_LOC_387/Y 0.01fF
C10436 INVX1_LOC_74/Y INVX1_LOC_59/A 0.03fF
C10437 NAND2X1_LOC_333/B NAND2X1_LOC_790/a_36_24# 0.00fF
C10438 INVX1_LOC_364/Y NAND2X1_LOC_457/a_36_24# 0.00fF
C10439 INVX1_LOC_62/Y INVX1_LOC_136/Y 0.01fF
C10440 INVX1_LOC_448/A INVX1_LOC_41/Y 0.07fF
C10441 INVX1_LOC_432/A INVX1_LOC_245/A 0.00fF
C10442 NAND2X1_LOC_307/A NAND2X1_LOC_544/B 0.03fF
C10443 INVX1_LOC_545/Y NAND2X1_LOC_544/B 0.02fF
C10444 NAND2X1_LOC_333/A INVX1_LOC_49/Y 0.01fF
C10445 INVX1_LOC_435/A INVX1_LOC_79/A 0.07fF
C10446 INVX1_LOC_400/A INVX1_LOC_100/Y 0.16fF
C10447 INVX1_LOC_477/Y INVX1_LOC_58/Y 0.04fF
C10448 INVX1_LOC_347/Y INVX1_LOC_372/A 0.02fF
C10449 INVX1_LOC_145/Y INVX1_LOC_41/Y 0.16fF
C10450 NAND2X1_LOC_766/a_36_24# INVX1_LOC_26/Y 0.00fF
C10451 INVX1_LOC_516/A INVX1_LOC_74/Y 0.01fF
C10452 INVX1_LOC_50/A INVX1_LOC_18/Y 0.01fF
C10453 INVX1_LOC_21/Y INVX1_LOC_211/A 0.04fF
C10454 INVX1_LOC_170/A INVX1_LOC_49/Y 0.01fF
C10455 INVX1_LOC_17/Y INVX1_LOC_388/A 0.04fF
C10456 INVX1_LOC_188/Y NAND2X1_LOC_832/A 0.03fF
C10457 INVX1_LOC_199/Y NAND2X1_LOC_847/A 0.02fF
C10458 INVX1_LOC_58/Y INVX1_LOC_139/Y 0.01fF
C10459 INVX1_LOC_679/A NAND2X1_LOC_843/B 0.01fF
C10460 INVX1_LOC_400/A INVX1_LOC_74/Y 0.11fF
C10461 INVX1_LOC_93/Y INVX1_LOC_100/Y 0.35fF
C10462 INVX1_LOC_159/Y NAND2X1_LOC_372/Y 0.00fF
C10463 INVX1_LOC_376/A INVX1_LOC_501/A 0.08fF
C10464 INVX1_LOC_248/A INVX1_LOC_41/Y 0.08fF
C10465 INVX1_LOC_496/A NAND2X1_LOC_221/a_36_24# 0.00fF
C10466 INVX1_LOC_116/Y INVX1_LOC_634/Y 0.14fF
C10467 NAND2X1_LOC_301/B INVX1_LOC_69/Y 0.03fF
C10468 NAND2X1_LOC_837/B INVX1_LOC_658/Y 0.33fF
C10469 INVX1_LOC_49/Y INVX1_LOC_488/A 0.07fF
C10470 INVX1_LOC_93/Y INVX1_LOC_74/Y 0.18fF
C10471 INVX1_LOC_108/A INVX1_LOC_479/A 0.00fF
C10472 INVX1_LOC_93/Y INVX1_LOC_483/Y 0.00fF
C10473 INVX1_LOC_141/Y INVX1_LOC_41/Y 0.00fF
C10474 INVX1_LOC_50/Y INVX1_LOC_488/Y 0.08fF
C10475 NAND2X1_LOC_490/a_36_24# INVX1_LOC_41/Y 0.00fF
C10476 INVX1_LOC_584/A INVX1_LOC_638/A 0.02fF
C10477 INVX1_LOC_117/A INVX1_LOC_26/Y 0.02fF
C10478 NAND2X1_LOC_274/B INVX1_LOC_518/A 0.04fF
C10479 INVX1_LOC_166/Y INVX1_LOC_15/Y 0.04fF
C10480 NAND2X1_LOC_334/A NAND2X1_LOC_597/Y 0.01fF
C10481 INVX1_LOC_100/Y INVX1_LOC_643/Y 0.01fF
C10482 INVX1_LOC_675/A INVX1_LOC_74/Y 0.16fF
C10483 INVX1_LOC_446/A INVX1_LOC_435/Y 0.01fF
C10484 INVX1_LOC_62/Y INVX1_LOC_15/Y 0.01fF
C10485 INVX1_LOC_601/Y INVX1_LOC_619/Y 0.01fF
C10486 VDD INVX1_LOC_200/Y 0.21fF
C10487 INVX1_LOC_424/A INVX1_LOC_421/Y 0.01fF
C10488 INVX1_LOC_31/Y INVX1_LOC_636/A 0.07fF
C10489 INVX1_LOC_255/A INVX1_LOC_634/Y 0.02fF
C10490 INVX1_LOC_317/Y INVX1_LOC_301/A 0.00fF
C10491 VDD INVX1_LOC_413/Y 0.53fF
C10492 NAND2X1_LOC_392/a_36_24# NAND2X1_LOC_475/A 0.00fF
C10493 INVX1_LOC_80/A INVX1_LOC_615/A 0.10fF
C10494 INVX1_LOC_12/Y INVX1_LOC_297/Y 0.03fF
C10495 INVX1_LOC_319/A INVX1_LOC_666/Y 0.00fF
C10496 NAND2X1_LOC_93/Y INVX1_LOC_291/A 0.04fF
C10497 INVX1_LOC_618/A INVX1_LOC_252/A 0.27fF
C10498 NAND2X1_LOC_710/a_36_24# INVX1_LOC_510/Y 0.01fF
C10499 INVX1_LOC_418/A INVX1_LOC_442/A 0.15fF
C10500 NAND2X1_LOC_791/B NAND2X1_LOC_358/a_36_24# 0.00fF
C10501 INPUT_3 INVX1_LOC_49/A 0.01fF
C10502 INVX1_LOC_412/Y NAND2X1_LOC_299/Y 0.16fF
C10503 VDD INVX1_LOC_154/Y 0.29fF
C10504 VDD INVX1_LOC_288/Y 0.21fF
C10505 NAND2X1_LOC_384/a_36_24# INVX1_LOC_321/A 0.00fF
C10506 INVX1_LOC_20/Y INVX1_LOC_317/Y 0.19fF
C10507 INVX1_LOC_395/A INVX1_LOC_320/A 0.01fF
C10508 INVX1_LOC_21/Y INVX1_LOC_257/Y 0.07fF
C10509 INVX1_LOC_53/Y INVX1_LOC_412/A 0.01fF
C10510 INVX1_LOC_578/A INVX1_LOC_197/A 0.07fF
C10511 INVX1_LOC_404/Y INVX1_LOC_99/Y 0.03fF
C10512 INVX1_LOC_133/Y INVX1_LOC_627/Y 0.00fF
C10513 INVX1_LOC_53/Y INVX1_LOC_618/Y 0.01fF
C10514 INVX1_LOC_409/A INVX1_LOC_352/Y 0.01fF
C10515 NAND2X1_LOC_331/A INVX1_LOC_99/Y 0.03fF
C10516 INVX1_LOC_171/Y INVX1_LOC_175/A 0.00fF
C10517 INVX1_LOC_198/A NAND2X1_LOC_205/a_36_24# 0.00fF
C10518 NAND2X1_LOC_45/Y INVX1_LOC_480/Y 0.01fF
C10519 INVX1_LOC_255/Y NAND2X1_LOC_123/A 0.10fF
C10520 INVX1_LOC_447/A INPUT_1 0.06fF
C10521 INVX1_LOC_335/Y INVX1_LOC_288/A 0.07fF
C10522 INVX1_LOC_463/A NAND2X1_LOC_688/a_36_24# 0.00fF
C10523 INVX1_LOC_293/Y INVX1_LOC_235/Y 0.02fF
C10524 INVX1_LOC_374/A INVX1_LOC_504/A 0.25fF
C10525 INVX1_LOC_12/Y INVX1_LOC_76/Y 0.08fF
C10526 INVX1_LOC_317/Y INVX1_LOC_300/A 0.20fF
C10527 NAND2X1_LOC_45/Y INVX1_LOC_169/Y 0.10fF
C10528 INVX1_LOC_418/A INVX1_LOC_116/Y 0.01fF
C10529 INVX1_LOC_625/A NAND2X1_LOC_335/a_36_24# 0.01fF
C10530 INVX1_LOC_224/Y INVX1_LOC_260/Y 0.01fF
C10531 INVX1_LOC_301/A NAND2X1_LOC_111/Y 0.09fF
C10532 INVX1_LOC_21/Y INVX1_LOC_384/A 0.10fF
C10533 INVX1_LOC_407/Y INVX1_LOC_570/A 0.25fF
C10534 INVX1_LOC_395/A NAND2X1_LOC_720/A 0.01fF
C10535 INVX1_LOC_315/Y INVX1_LOC_145/Y 0.02fF
C10536 NAND2X1_LOC_121/a_36_24# INVX1_LOC_632/A 0.01fF
C10537 INVX1_LOC_20/Y INVX1_LOC_106/A 0.05fF
C10538 INVX1_LOC_63/Y NAND2X1_LOC_76/B 0.18fF
C10539 INVX1_LOC_408/Y INVX1_LOC_46/Y 0.01fF
C10540 INVX1_LOC_629/Y INVX1_LOC_261/Y 0.15fF
C10541 INVX1_LOC_340/Y INVX1_LOC_513/A 0.00fF
C10542 INVX1_LOC_442/A INVX1_LOC_46/Y 0.07fF
C10543 INVX1_LOC_17/Y INVX1_LOC_655/Y 0.01fF
C10544 INVX1_LOC_384/A NAND2X1_LOC_274/a_36_24# 0.00fF
C10545 INVX1_LOC_629/A INVX1_LOC_675/A 0.03fF
C10546 NAND2X1_LOC_318/A NAND2X1_LOC_615/B 0.28fF
C10547 INVX1_LOC_602/A INVX1_LOC_35/Y 0.07fF
C10548 INVX1_LOC_258/A INVX1_LOC_504/Y 0.01fF
C10549 NAND2X1_LOC_513/A INVX1_LOC_338/A 0.08fF
C10550 NAND2X1_LOC_411/Y NAND2X1_LOC_413/Y 0.01fF
C10551 INVX1_LOC_358/Y INVX1_LOC_145/Y 0.04fF
C10552 INVX1_LOC_392/Y NAND2X1_LOC_181/A 0.14fF
C10553 INVX1_LOC_522/Y INPUT_1 0.17fF
C10554 NAND2X1_LOC_571/a_36_24# INVX1_LOC_17/Y 0.00fF
C10555 INVX1_LOC_20/Y INVX1_LOC_166/A 0.39fF
C10556 INVX1_LOC_87/Y INVX1_LOC_88/Y 0.01fF
C10557 INVX1_LOC_381/A INVX1_LOC_31/Y 0.07fF
C10558 NAND2X1_LOC_543/B INVX1_LOC_62/Y 0.55fF
C10559 INVX1_LOC_21/Y INVX1_LOC_145/Y 0.87fF
C10560 INVX1_LOC_43/Y INVX1_LOC_44/A 0.01fF
C10561 INVX1_LOC_93/Y INVX1_LOC_566/A 0.14fF
C10562 INVX1_LOC_20/Y NAND2X1_LOC_849/a_36_24# 0.01fF
C10563 INPUT_0 INVX1_LOC_26/Y 0.33fF
C10564 INPUT_0 INVX1_LOC_128/Y 0.03fF
C10565 INVX1_LOC_20/Y INVX1_LOC_239/A 0.01fF
C10566 NAND2X1_LOC_13/Y INVX1_LOC_6/Y 0.00fF
C10567 INVX1_LOC_482/A NAND2X1_LOC_613/a_36_24# 0.00fF
C10568 INVX1_LOC_407/Y INVX1_LOC_99/Y 0.09fF
C10569 INVX1_LOC_551/Y INVX1_LOC_69/Y 0.05fF
C10570 INVX1_LOC_137/Y INVX1_LOC_610/A -0.00fF
C10571 INVX1_LOC_391/Y INVX1_LOC_367/Y 0.02fF
C10572 INVX1_LOC_170/A INVX1_LOC_76/Y 0.00fF
C10573 INVX1_LOC_251/A INVX1_LOC_251/Y 0.03fF
C10574 INVX1_LOC_395/A INVX1_LOC_100/Y 3.59fF
C10575 NAND2X1_LOC_516/Y INVX1_LOC_128/Y 0.44fF
C10576 INVX1_LOC_99/Y INVX1_LOC_480/Y 0.03fF
C10577 INVX1_LOC_384/Y GATE_479 0.04fF
C10578 INVX1_LOC_670/Y INVX1_LOC_520/A 0.00fF
C10579 NAND2X1_LOC_861/a_36_24# INVX1_LOC_51/Y 0.01fF
C10580 INVX1_LOC_581/A INVX1_LOC_627/Y 0.02fF
C10581 INVX1_LOC_168/A INVX1_LOC_58/Y 0.01fF
C10582 INVX1_LOC_557/Y INVX1_LOC_51/Y 0.04fF
C10583 INVX1_LOC_546/Y INVX1_LOC_79/A 0.01fF
C10584 NAND2X1_LOC_37/a_36_24# INVX1_LOC_451/A 0.09fF
C10585 INVX1_LOC_588/Y INVX1_LOC_300/A 0.07fF
C10586 INPUT_0 NAND2X1_LOC_608/a_36_24# 0.00fF
C10587 INVX1_LOC_683/A INVX1_LOC_105/Y 0.01fF
C10588 INVX1_LOC_273/A INVX1_LOC_399/Y -0.00fF
C10589 INVX1_LOC_305/Y INVX1_LOC_46/Y 0.01fF
C10590 INVX1_LOC_628/A INVX1_LOC_93/Y 0.00fF
C10591 NAND2X1_LOC_192/a_36_24# INVX1_LOC_496/A 0.00fF
C10592 NAND2X1_LOC_106/Y NAND2X1_LOC_496/Y 0.04fF
C10593 INVX1_LOC_435/A INVX1_LOC_48/Y 0.02fF
C10594 INVX1_LOC_545/A INVX1_LOC_54/Y 0.00fF
C10595 INVX1_LOC_206/Y INVX1_LOC_483/A 0.00fF
C10596 INVX1_LOC_202/Y NAND2X1_LOC_615/B 0.04fF
C10597 INVX1_LOC_117/Y INVX1_LOC_379/A 0.09fF
C10598 INVX1_LOC_586/A NAND2X1_LOC_301/B 0.05fF
C10599 INVX1_LOC_362/Y INVX1_LOC_100/Y 0.07fF
C10600 INVX1_LOC_617/A INVX1_LOC_9/Y 0.03fF
C10601 INVX1_LOC_602/A INVX1_LOC_621/Y 0.01fF
C10602 INVX1_LOC_99/Y INVX1_LOC_169/Y 0.01fF
C10603 INVX1_LOC_17/Y NAND2X1_LOC_507/A 0.18fF
C10604 INVX1_LOC_395/A INVX1_LOC_74/Y 0.00fF
C10605 INVX1_LOC_117/Y INVX1_LOC_35/Y 0.39fF
C10606 INVX1_LOC_566/A NAND2X1_LOC_334/B 0.00fF
C10607 INVX1_LOC_139/A INVX1_LOC_479/A 0.03fF
C10608 INVX1_LOC_116/Y INVX1_LOC_46/Y 0.07fF
C10609 INVX1_LOC_555/A NAND2X1_LOC_612/A 0.03fF
C10610 INVX1_LOC_78/A NAND2X1_LOC_308/A 0.01fF
C10611 INVX1_LOC_438/A INVX1_LOC_488/Y 0.02fF
C10612 INVX1_LOC_555/A INVX1_LOC_145/Y 0.03fF
C10613 INVX1_LOC_53/Y NAND2X1_LOC_847/A 0.01fF
C10614 INVX1_LOC_76/Y INVX1_LOC_488/A 0.01fF
C10615 INVX1_LOC_267/A INVX1_LOC_59/Y 0.01fF
C10616 INVX1_LOC_20/Y INVX1_LOC_153/Y 0.20fF
C10617 INVX1_LOC_575/A INVX1_LOC_568/A 0.02fF
C10618 INVX1_LOC_607/A NAND2X1_LOC_248/B 0.31fF
C10619 INVX1_LOC_530/A INVX1_LOC_63/Y 0.03fF
C10620 INVX1_LOC_17/Y INVX1_LOC_89/Y 0.04fF
C10621 INVX1_LOC_145/Y INVX1_LOC_181/Y 0.01fF
C10622 INVX1_LOC_331/Y NAND2X1_LOC_679/B 0.01fF
C10623 INVX1_LOC_437/A INVX1_LOC_387/Y 0.01fF
C10624 INVX1_LOC_628/A INVX1_LOC_675/A 0.02fF
C10625 NAND2X1_LOC_332/B INVX1_LOC_41/Y 0.05fF
C10626 INVX1_LOC_545/A INVX1_LOC_257/A 0.04fF
C10627 INVX1_LOC_530/Y NAND2X1_LOC_621/B 0.04fF
C10628 INVX1_LOC_392/A NAND2X1_LOC_181/A 0.42fF
C10629 INVX1_LOC_683/Y INVX1_LOC_100/Y 0.03fF
C10630 INVX1_LOC_20/Y INVX1_LOC_531/Y 0.11fF
C10631 INVX1_LOC_625/A INVX1_LOC_63/Y 0.04fF
C10632 INVX1_LOC_309/Y INVX1_LOC_7/Y 0.04fF
C10633 INVX1_LOC_425/Y INVX1_LOC_47/Y 0.11fF
C10634 INVX1_LOC_469/Y INVX1_LOC_93/Y 0.03fF
C10635 INVX1_LOC_107/Y INVX1_LOC_145/Y 0.00fF
C10636 INVX1_LOC_46/Y INVX1_LOC_328/A 0.00fF
C10637 NAND2X1_LOC_106/Y NAND2X1_LOC_706/B 0.36fF
C10638 INVX1_LOC_296/Y INVX1_LOC_245/A 0.01fF
C10639 INVX1_LOC_17/Y INVX1_LOC_501/A 0.03fF
C10640 INVX1_LOC_271/A INVX1_LOC_270/Y 0.01fF
C10641 NAND2X1_LOC_755/B NAND2X1_LOC_719/A 0.06fF
C10642 INVX1_LOC_519/Y INVX1_LOC_670/Y 0.03fF
C10643 INVX1_LOC_119/A INVX1_LOC_75/Y 0.02fF
C10644 INVX1_LOC_106/A INVX1_LOC_655/A 0.03fF
C10645 INVX1_LOC_93/Y NAND2X1_LOC_181/A 0.01fF
C10646 INVX1_LOC_586/A INVX1_LOC_291/Y 0.03fF
C10647 INVX1_LOC_508/A INPUT_1 0.03fF
C10648 NAND2X1_LOC_274/B INVX1_LOC_352/A 0.03fF
C10649 INVX1_LOC_561/A INVX1_LOC_261/Y 0.00fF
C10650 INVX1_LOC_201/A INVX1_LOC_26/Y 0.03fF
C10651 INVX1_LOC_300/A INVX1_LOC_153/Y 0.08fF
C10652 INVX1_LOC_516/A INVX1_LOC_79/A 0.01fF
C10653 INVX1_LOC_80/A INVX1_LOC_274/Y 0.01fF
C10654 INVX1_LOC_255/A INVX1_LOC_46/Y 0.16fF
C10655 INVX1_LOC_117/Y INVX1_LOC_621/Y 0.04fF
C10656 INVX1_LOC_507/Y INVX1_LOC_50/Y 0.01fF
C10657 INVX1_LOC_400/A INVX1_LOC_77/A 0.01fF
C10658 INVX1_LOC_89/Y NAND2X1_LOC_307/B 0.17fF
C10659 INVX1_LOC_469/Y INVX1_LOC_675/A 0.08fF
C10660 INVX1_LOC_208/Y INVX1_LOC_63/Y 0.03fF
C10661 INVX1_LOC_455/A NAND2X1_LOC_823/Y 0.05fF
C10662 INVX1_LOC_223/Y INVX1_LOC_50/Y 0.01fF
C10663 INVX1_LOC_51/Y INVX1_LOC_636/A 0.22fF
C10664 INVX1_LOC_6/Y NAND2X1_LOC_668/Y 0.01fF
C10665 INVX1_LOC_49/Y INVX1_LOC_66/A 0.16fF
C10666 INVX1_LOC_548/A INVX1_LOC_100/Y 0.51fF
C10667 INVX1_LOC_531/Y INVX1_LOC_197/Y 0.07fF
C10668 INVX1_LOC_508/A NAND2X1_LOC_277/a_36_24# 0.01fF
C10669 INVX1_LOC_480/Y NAND2X1_LOC_66/Y 0.03fF
C10670 INVX1_LOC_199/Y INVX1_LOC_77/Y 0.04fF
C10671 NAND2X1_LOC_184/Y INVX1_LOC_664/A 0.21fF
C10672 INVX1_LOC_298/A INVX1_LOC_26/Y 0.03fF
C10673 INVX1_LOC_69/Y NAND2X1_LOC_759/Y 0.01fF
C10674 INVX1_LOC_326/Y INVX1_LOC_9/Y 0.07fF
C10675 INVX1_LOC_496/A INVX1_LOC_338/Y 0.00fF
C10676 INVX1_LOC_479/A NAND2X1_LOC_259/A 0.04fF
C10677 INVX1_LOC_17/Y NAND2X1_LOC_544/B 0.52fF
C10678 INVX1_LOC_93/Y INVX1_LOC_79/A 12.60fF
C10679 NAND2X1_LOC_66/Y INVX1_LOC_169/Y 0.01fF
C10680 INVX1_LOC_31/Y INVX1_LOC_100/Y 0.39fF
C10681 INVX1_LOC_239/A INVX1_LOC_655/A 0.01fF
C10682 INVX1_LOC_32/Y NAND2X1_LOC_528/Y 0.46fF
C10683 INVX1_LOC_242/Y INVX1_LOC_411/Y 0.10fF
C10684 INVX1_LOC_17/A INVX1_LOC_66/A 0.04fF
C10685 INVX1_LOC_361/Y INVX1_LOC_666/Y 0.00fF
C10686 INVX1_LOC_31/Y INVX1_LOC_74/Y 0.44fF
C10687 INVX1_LOC_32/Y INVX1_LOC_479/A 0.10fF
C10688 INVX1_LOC_675/A INVX1_LOC_79/A 0.07fF
C10689 INVX1_LOC_183/Y INVX1_LOC_82/Y 0.02fF
C10690 INVX1_LOC_49/Y NAND2X1_LOC_601/Y 0.02fF
C10691 INVX1_LOC_390/A INVX1_LOC_79/A 0.00fF
C10692 INVX1_LOC_100/Y INVX1_LOC_682/Y 0.05fF
C10693 INVX1_LOC_675/A INVX1_LOC_460/A 0.04fF
C10694 INVX1_LOC_454/A NAND2X1_LOC_581/a_36_24# 0.02fF
C10695 NAND2X1_LOC_334/B INVX1_LOC_79/A 0.00fF
C10696 NAND2X1_LOC_775/B INVX1_LOC_92/A 0.07fF
C10697 INVX1_LOC_523/Y INVX1_LOC_647/Y 0.03fF
C10698 INVX1_LOC_41/Y INVX1_LOC_242/Y 0.19fF
C10699 INVX1_LOC_69/Y INVX1_LOC_634/Y 0.06fF
C10700 INVX1_LOC_563/Y INVX1_LOC_206/Y 0.03fF
C10701 INVX1_LOC_114/Y INVX1_LOC_638/A 0.05fF
C10702 NAND2X1_LOC_242/A INVX1_LOC_395/A 0.08fF
C10703 INPUT_0 INVX1_LOC_560/A 0.42fF
C10704 INVX1_LOC_26/Y INVX1_LOC_211/A 0.97fF
C10705 INVX1_LOC_683/A INVX1_LOC_109/Y 0.01fF
C10706 INVX1_LOC_257/Y INVX1_LOC_255/Y 0.04fF
C10707 NAND2X1_LOC_475/A INVX1_LOC_271/Y 0.01fF
C10708 INVX1_LOC_393/Y INVX1_LOC_490/Y 0.11fF
C10709 VDD NAND2X1_LOC_180/B 0.26fF
C10710 INVX1_LOC_348/Y INVX1_LOC_114/A 0.01fF
C10711 INVX1_LOC_203/Y INVX1_LOC_286/Y 0.27fF
C10712 INVX1_LOC_454/A INVX1_LOC_55/Y 0.03fF
C10713 VDD NAND2X1_LOC_728/B 0.03fF
C10714 VDD INVX1_LOC_311/Y 0.26fF
C10715 INVX1_LOC_255/Y INVX1_LOC_288/A 0.02fF
C10716 NAND2X1_LOC_776/a_36_24# INVX1_LOC_273/A 0.01fF
C10717 VDD INVX1_LOC_324/Y 0.28fF
C10718 NAND2X1_LOC_176/Y NAND2X1_LOC_307/A 0.28fF
C10719 INVX1_LOC_99/Y INVX1_LOC_638/A 0.07fF
C10720 VDD INVX1_LOC_188/Y 0.36fF
C10721 VDD INVX1_LOC_603/Y 0.38fF
C10722 NAND2X1_LOC_516/B NAND2X1_LOC_513/Y 0.05fF
C10723 VDD NAND2X1_LOC_411/Y 0.00fF
C10724 INVX1_LOC_185/A INVX1_LOC_35/Y 0.00fF
C10725 VDD INVX1_LOC_43/Y 0.39fF
C10726 INVX1_LOC_224/Y NAND2X1_LOC_97/B 0.02fF
C10727 INVX1_LOC_612/Y INVX1_LOC_627/A 0.00fF
C10728 INVX1_LOC_607/Y NAND2X1_LOC_249/Y 0.09fF
C10729 INPUT_0 INVX1_LOC_369/A 0.00fF
C10730 INVX1_LOC_224/Y INVX1_LOC_417/A 0.02fF
C10731 INVX1_LOC_381/A INVX1_LOC_51/Y 0.07fF
C10732 INVX1_LOC_144/Y INVX1_LOC_142/A 0.20fF
C10733 INVX1_LOC_551/Y INVX1_LOC_586/A 0.46fF
C10734 INVX1_LOC_400/Y INVX1_LOC_134/Y 0.07fF
C10735 NAND2X1_LOC_97/B INVX1_LOC_578/A 0.02fF
C10736 VDD INVX1_LOC_478/Y 0.21fF
C10737 INVX1_LOC_385/Y INVX1_LOC_445/A 0.03fF
C10738 VDD INVX1_LOC_403/Y 0.21fF
C10739 INVX1_LOC_20/Y NAND2X1_LOC_467/A 0.08fF
C10740 VDD INVX1_LOC_382/Y 0.20fF
C10741 INVX1_LOC_402/Y NAND2X1_LOC_513/Y 0.00fF
C10742 INVX1_LOC_31/Y NAND2X1_LOC_591/B 0.76fF
C10743 INVX1_LOC_60/Y INVX1_LOC_55/Y 0.01fF
C10744 INVX1_LOC_447/A INVX1_LOC_50/Y 0.03fF
C10745 NAND2X1_LOC_45/Y INVX1_LOC_665/Y 0.04fF
C10746 VDD NAND2X1_LOC_387/Y 0.03fF
C10747 INVX1_LOC_224/Y INVX1_LOC_440/Y 0.01fF
C10748 INVX1_LOC_47/Y INVX1_LOC_638/A 0.09fF
C10749 NAND2X1_LOC_274/B INVX1_LOC_109/Y 0.03fF
C10750 INVX1_LOC_446/Y INVX1_LOC_444/Y 0.07fF
C10751 INVX1_LOC_445/Y INVX1_LOC_451/A 0.03fF
C10752 INVX1_LOC_454/A INVX1_LOC_18/Y 0.04fF
C10753 NAND2X1_LOC_526/a_36_24# INVX1_LOC_145/Y 0.01fF
C10754 NAND2X1_LOC_475/A NAND2X1_LOC_265/a_36_24# 0.00fF
C10755 NAND2X1_LOC_703/a_36_24# INVX1_LOC_442/A 0.00fF
C10756 INVX1_LOC_425/A INVX1_LOC_99/A 0.24fF
C10757 INVX1_LOC_217/A NAND2X1_LOC_252/Y 0.00fF
C10758 INVX1_LOC_166/A INVX1_LOC_553/A 0.01fF
C10759 INVX1_LOC_578/A INVX1_LOC_440/Y 0.02fF
C10760 INVX1_LOC_197/A INVX1_LOC_686/A 0.07fF
C10761 INVX1_LOC_577/A INVX1_LOC_93/Y 0.11fF
C10762 NAND2X1_LOC_498/Y INVX1_LOC_665/Y 0.03fF
C10763 INVX1_LOC_301/A INVX1_LOC_411/Y 0.00fF
C10764 INVX1_LOC_228/Y NAND2X1_LOC_387/Y 0.00fF
C10765 NAND2X1_LOC_561/a_36_24# INVX1_LOC_321/A 0.00fF
C10766 INVX1_LOC_577/Y INVX1_LOC_145/Y 0.02fF
C10767 NAND2X1_LOC_788/A INVX1_LOC_49/Y 0.05fF
C10768 INVX1_LOC_570/A INVX1_LOC_575/Y 0.06fF
C10769 INVX1_LOC_444/Y INVX1_LOC_384/A 0.00fF
C10770 INVX1_LOC_398/A INVX1_LOC_99/Y 0.01fF
C10771 INVX1_LOC_438/A INVX1_LOC_378/Y 0.03fF
C10772 INVX1_LOC_392/Y INVX1_LOC_48/Y 0.03fF
C10773 INVX1_LOC_428/A NAND2X1_LOC_693/a_36_24# 0.00fF
C10774 INVX1_LOC_452/A INVX1_LOC_384/Y 0.31fF
C10775 INVX1_LOC_51/Y NAND2X1_LOC_720/A 0.15fF
C10776 NAND2X1_LOC_701/a_36_24# INVX1_LOC_47/Y 0.01fF
C10777 NAND2X1_LOC_88/B INVX1_LOC_21/Y 0.03fF
C10778 INVX1_LOC_301/A INVX1_LOC_301/Y 0.05fF
C10779 INVX1_LOC_586/A INVX1_LOC_493/A 0.00fF
C10780 INVX1_LOC_524/Y INVX1_LOC_59/Y 0.01fF
C10781 INVX1_LOC_570/Y INVX1_LOC_662/A 0.02fF
C10782 NAND2X1_LOC_88/Y INVX1_LOC_179/Y 0.00fF
C10783 VDD NAND2X1_LOC_845/B 0.32fF
C10784 NAND2X1_LOC_335/B INVX1_LOC_9/Y 0.01fF
C10785 NAND2X1_LOC_666/Y INVX1_LOC_562/A 0.44fF
C10786 INVX1_LOC_76/Y NAND2X1_LOC_615/B 0.04fF
C10787 INVX1_LOC_570/A NAND2X1_LOC_308/A 0.07fF
C10788 NAND2X1_LOC_164/Y INVX1_LOC_63/Y 0.04fF
C10789 INVX1_LOC_35/Y INVX1_LOC_658/A 0.08fF
C10790 INVX1_LOC_12/Y INVX1_LOC_7/Y 0.03fF
C10791 INVX1_LOC_191/Y INVX1_LOC_543/A 0.03fF
C10792 INVX1_LOC_524/Y INVX1_LOC_48/Y 0.03fF
C10793 INVX1_LOC_575/A INVX1_LOC_136/Y 0.01fF
C10794 INVX1_LOC_12/Y INVX1_LOC_228/A 0.05fF
C10795 INVX1_LOC_133/A INVX1_LOC_240/A 0.24fF
C10796 NAND2X1_LOC_137/A NAND2X1_LOC_332/B 0.07fF
C10797 INVX1_LOC_509/Y INVX1_LOC_516/A 0.00fF
C10798 INVX1_LOC_362/Y NAND2X1_LOC_181/A 0.07fF
C10799 INVX1_LOC_418/A INVX1_LOC_69/Y 0.01fF
C10800 INVX1_LOC_33/Y INVX1_LOC_204/Y 0.01fF
C10801 INVX1_LOC_522/Y INVX1_LOC_50/Y 0.05fF
C10802 INVX1_LOC_407/Y INVX1_LOC_136/Y 0.01fF
C10803 NAND2X1_LOC_174/B INVX1_LOC_686/A 0.03fF
C10804 INVX1_LOC_409/Y INVX1_LOC_62/Y 0.03fF
C10805 NAND2X1_LOC_592/B INVX1_LOC_501/A 0.01fF
C10806 NAND2X1_LOC_427/Y INVX1_LOC_463/Y 0.03fF
C10807 INVX1_LOC_406/Y NAND2X1_LOC_184/Y 0.00fF
C10808 INVX1_LOC_301/A INVX1_LOC_41/Y 0.22fF
C10809 INVX1_LOC_323/Y INVX1_LOC_176/A 0.00fF
C10810 INVX1_LOC_184/A INVX1_LOC_86/Y 0.11fF
C10811 INVX1_LOC_333/Y INVX1_LOC_25/Y 0.24fF
C10812 INVX1_LOC_566/A INVX1_LOC_31/Y 0.15fF
C10813 INVX1_LOC_372/Y INVX1_LOC_345/Y -0.00fF
C10814 INVX1_LOC_40/Y INVX1_LOC_29/Y 0.37fF
C10815 NAND2X1_LOC_591/Y INVX1_LOC_686/A 0.02fF
C10816 INVX1_LOC_65/Y INVX1_LOC_63/Y 0.28fF
C10817 INVX1_LOC_589/Y INVX1_LOC_398/A 0.35fF
C10818 INVX1_LOC_395/A NAND2X1_LOC_558/B 0.00fF
C10819 INVX1_LOC_612/Y INVX1_LOC_581/A 0.02fF
C10820 INVX1_LOC_324/A INVX1_LOC_327/Y 0.15fF
C10821 INVX1_LOC_363/Y INVX1_LOC_116/Y 0.01fF
C10822 INVX1_LOC_444/Y INVX1_LOC_145/Y 0.03fF
C10823 NAND2X1_LOC_137/A INVX1_LOC_125/Y 0.05fF
C10824 NAND2X1_LOC_701/a_36_24# INVX1_LOC_119/Y 0.00fF
C10825 INVX1_LOC_76/Y INVX1_LOC_296/A 0.02fF
C10826 INVX1_LOC_573/Y INVX1_LOC_515/A 0.00fF
C10827 NAND2X1_LOC_739/a_36_24# INVX1_LOC_62/Y 0.00fF
C10828 NAND2X1_LOC_697/Y INVX1_LOC_609/A 0.13fF
C10829 NAND2X1_LOC_726/a_36_24# INVX1_LOC_6/Y 0.00fF
C10830 INVX1_LOC_437/A INVX1_LOC_386/Y 0.08fF
C10831 INVX1_LOC_270/A INVX1_LOC_69/Y 0.72fF
C10832 INVX1_LOC_35/Y INVX1_LOC_178/A 0.00fF
C10833 INVX1_LOC_395/A INVX1_LOC_79/A 2.51fF
C10834 INVX1_LOC_400/A INVX1_LOC_59/Y 0.00fF
C10835 INVX1_LOC_421/A INVX1_LOC_134/Y 0.00fF
C10836 INVX1_LOC_17/Y INVX1_LOC_194/Y 0.10fF
C10837 NAND2X1_LOC_152/B INVX1_LOC_6/Y 0.03fF
C10838 INVX1_LOC_293/A INVX1_LOC_654/A 0.15fF
C10839 INVX1_LOC_12/Y INVX1_LOC_32/Y 0.07fF
C10840 INVX1_LOC_11/Y INVX1_LOC_230/A 0.19fF
C10841 INVX1_LOC_511/Y INVX1_LOC_514/A 0.00fF
C10842 INVX1_LOC_417/Y INVX1_LOC_93/Y 0.43fF
C10843 INVX1_LOC_288/A INVX1_LOC_26/Y 0.03fF
C10844 INVX1_LOC_93/Y INVX1_LOC_509/Y 0.01fF
C10845 NAND2X1_LOC_505/Y INVX1_LOC_100/Y 0.01fF
C10846 NAND2X1_LOC_318/A INVX1_LOC_179/A 0.07fF
C10847 INVX1_LOC_586/A INVX1_LOC_500/A 0.01fF
C10848 INVX1_LOC_62/A INVX1_LOC_98/Y 0.03fF
C10849 INVX1_LOC_166/A NAND2X1_LOC_140/B 0.04fF
C10850 INVX1_LOC_400/A INVX1_LOC_48/Y 0.07fF
C10851 INVX1_LOC_133/Y INVX1_LOC_92/A 0.00fF
C10852 INVX1_LOC_117/Y INVX1_LOC_338/A 0.02fF
C10853 INVX1_LOC_20/Y INVX1_LOC_301/Y 0.03fF
C10854 INVX1_LOC_410/Y INVX1_LOC_75/Y 0.08fF
C10855 INPUT_3 INVX1_LOC_183/A 0.03fF
C10856 INVX1_LOC_51/Y INVX1_LOC_100/Y 0.26fF
C10857 INVX1_LOC_384/A INVX1_LOC_26/Y 0.07fF
C10858 INVX1_LOC_50/Y NAND2X1_LOC_606/Y 0.04fF
C10859 INVX1_LOC_93/Y INVX1_LOC_59/Y 0.03fF
C10860 NAND2X1_LOC_775/B INPUT_1 0.44fF
C10861 NAND2X1_LOC_308/A INVX1_LOC_99/Y 0.00fF
C10862 NAND2X1_LOC_148/A NAND2X1_LOC_847/A 0.12fF
C10863 INVX1_LOC_662/A INVX1_LOC_517/A 0.14fF
C10864 NAND2X1_LOC_446/a_36_24# INVX1_LOC_66/A 0.01fF
C10865 INVX1_LOC_69/Y NAND2X1_LOC_755/B 0.07fF
C10866 INVX1_LOC_268/A INVX1_LOC_49/Y 0.08fF
C10867 INVX1_LOC_369/Y INVX1_LOC_378/A 0.01fF
C10868 NAND2X1_LOC_532/Y INVX1_LOC_98/Y 0.02fF
C10869 INVX1_LOC_117/Y INVX1_LOC_118/A 0.00fF
C10870 INVX1_LOC_266/A INVX1_LOC_100/Y 0.05fF
C10871 INVX1_LOC_604/Y INVX1_LOC_63/Y 0.08fF
C10872 INVX1_LOC_51/Y INVX1_LOC_74/Y 0.10fF
C10873 INVX1_LOC_93/Y INVX1_LOC_48/Y 0.29fF
C10874 INVX1_LOC_600/A INVX1_LOC_9/Y 0.03fF
C10875 NAND2X1_LOC_703/a_36_24# INVX1_LOC_255/A 0.00fF
C10876 INVX1_LOC_20/Y INVX1_LOC_41/Y 2.16fF
C10877 NAND2X1_LOC_130/Y INVX1_LOC_9/Y 0.03fF
C10878 NAND2X1_LOC_156/Y INVX1_LOC_168/Y 0.04fF
C10879 INVX1_LOC_62/Y INVX1_LOC_147/Y 0.17fF
C10880 INVX1_LOC_258/A INVX1_LOC_114/A 0.01fF
C10881 INVX1_LOC_255/A INVX1_LOC_349/Y -0.02fF
C10882 NAND2X1_LOC_387/Y INVX1_LOC_68/A 0.04fF
C10883 INVX1_LOC_47/Y INVX1_LOC_665/Y 0.03fF
C10884 INVX1_LOC_31/Y INVX1_LOC_350/Y 0.00fF
C10885 INVX1_LOC_183/A NAND2X1_LOC_376/Y 0.08fF
C10886 INVX1_LOC_35/Y INVX1_LOC_58/Y 2.16fF
C10887 INVX1_LOC_211/A NAND2X1_LOC_97/a_36_24# 0.01fF
C10888 INVX1_LOC_45/Y INVX1_LOC_109/A 0.00fF
C10889 NAND2X1_LOC_333/A INVX1_LOC_32/Y 0.04fF
C10890 INVX1_LOC_21/Y INVX1_LOC_242/Y 0.07fF
C10891 INVX1_LOC_511/Y INVX1_LOC_534/Y 0.26fF
C10892 NAND2X1_LOC_73/a_36_24# INVX1_LOC_9/Y 0.00fF
C10893 INVX1_LOC_452/A NAND2X1_LOC_555/B 3.32fF
C10894 INVX1_LOC_49/Y NAND2X1_LOC_432/Y 0.01fF
C10895 INVX1_LOC_448/A INVX1_LOC_128/Y 0.02fF
C10896 NAND2X1_LOC_123/B INVX1_LOC_633/Y 0.16fF
C10897 NAND2X1_LOC_334/B INVX1_LOC_59/Y 0.31fF
C10898 INVX1_LOC_202/Y INVX1_LOC_179/A 0.00fF
C10899 INVX1_LOC_675/A INVX1_LOC_48/Y 0.07fF
C10900 INVX1_LOC_76/Y NAND2X1_LOC_646/B 0.01fF
C10901 NAND2X1_LOC_791/A INVX1_LOC_26/Y 0.07fF
C10902 INVX1_LOC_284/A INVX1_LOC_79/A 0.09fF
C10903 INVX1_LOC_145/Y INVX1_LOC_26/Y 3.17fF
C10904 INVX1_LOC_69/Y INVX1_LOC_46/Y 1.01fF
C10905 INVX1_LOC_488/A INVX1_LOC_7/Y 0.01fF
C10906 INVX1_LOC_32/Y INVX1_LOC_188/A 0.01fF
C10907 NAND2X1_LOC_428/Y INVX1_LOC_495/A 0.05fF
C10908 INVX1_LOC_62/Y NAND2X1_LOC_302/A 0.04fF
C10909 INVX1_LOC_170/A INVX1_LOC_32/Y 0.09fF
C10910 INVX1_LOC_390/A INVX1_LOC_48/Y 0.01fF
C10911 NAND2X1_LOC_308/A INVX1_LOC_47/Y 0.03fF
C10912 INVX1_LOC_449/A NAND2X1_LOC_372/Y 0.45fF
C10913 GATE_662 INVX1_LOC_212/Y 0.01fF
C10914 INVX1_LOC_179/Y INVX1_LOC_198/A 0.01fF
C10915 INVX1_LOC_261/Y NAND2X1_LOC_355/A 0.02fF
C10916 INVX1_LOC_451/A NAND2X1_LOC_66/Y 0.03fF
C10917 INVX1_LOC_572/Y INVX1_LOC_58/Y 0.52fF
C10918 INVX1_LOC_300/A INVX1_LOC_41/Y 0.58fF
C10919 NAND2X1_LOC_532/Y INVX1_LOC_338/Y 0.07fF
C10920 INVX1_LOC_62/Y NAND2X1_LOC_73/a_36_24# 0.01fF
C10921 INVX1_LOC_41/Y INVX1_LOC_197/Y 0.01fF
C10922 INVX1_LOC_17/Y INVX1_LOC_347/A 0.01fF
C10923 INVX1_LOC_44/A INVX1_LOC_190/A 0.34fF
C10924 INVX1_LOC_545/A NAND2X1_LOC_544/B 0.00fF
C10925 INVX1_LOC_254/A INVX1_LOC_100/Y 0.03fF
C10926 NAND2X1_LOC_286/a_36_24# INVX1_LOC_655/A 0.00fF
C10927 INVX1_LOC_31/Y INVX1_LOC_79/A 0.87fF
C10928 INVX1_LOC_74/Y INVX1_LOC_40/Y 0.01fF
C10929 NAND2X1_LOC_300/a_36_24# INVX1_LOC_114/A 0.00fF
C10930 INVX1_LOC_569/Y NAND2X1_LOC_846/B 0.05fF
C10931 NAND2X1_LOC_308/A INVX1_LOC_119/Y 0.01fF
C10932 NAND2X1_LOC_646/A INVX1_LOC_588/A 0.01fF
C10933 NAND2X1_LOC_274/B INVX1_LOC_199/Y 0.03fF
C10934 INVX1_LOC_662/A NAND2X1_LOC_847/A 0.09fF
C10935 INVX1_LOC_63/Y NAND2X1_LOC_813/a_36_24# 0.00fF
C10936 INVX1_LOC_675/A NAND2X1_LOC_434/B 0.05fF
C10937 INVX1_LOC_254/A INVX1_LOC_74/Y 0.03fF
C10938 INVX1_LOC_110/A INVX1_LOC_479/A 0.04fF
C10939 INVX1_LOC_76/A INVX1_LOC_98/Y 0.05fF
C10940 INVX1_LOC_560/Y NAND2X1_LOC_76/B 0.03fF
C10941 INVX1_LOC_69/Y INVX1_LOC_75/A 0.08fF
C10942 INVX1_LOC_63/Y INVX1_LOC_588/A 0.03fF
C10943 NAND2X1_LOC_286/A INVX1_LOC_212/A 0.11fF
C10944 INVX1_LOC_317/A INVX1_LOC_92/A 0.02fF
C10945 VDD INVX1_LOC_269/A 0.00fF
C10946 INPUT_0 INVX1_LOC_373/A 0.76fF
C10947 INVX1_LOC_404/Y NAND2X1_LOC_520/B 0.02fF
C10948 NAND2X1_LOC_373/Y NAND2X1_LOC_322/a_36_24# 0.00fF
C10949 INVX1_LOC_114/A NAND2X1_LOC_832/A 0.03fF
C10950 INVX1_LOC_65/Y INVX1_LOC_552/Y 0.02fF
C10951 INVX1_LOC_159/Y INVX1_LOC_109/Y 0.03fF
C10952 INVX1_LOC_278/A NAND2X1_LOC_261/Y 0.01fF
C10953 INVX1_LOC_605/Y VDD 0.21fF
C10954 INVX1_LOC_416/Y INVX1_LOC_586/A 0.01fF
C10955 VDD NAND2X1_LOC_24/Y 0.13fF
C10956 INVX1_LOC_408/Y INVX1_LOC_76/Y 0.01fF
C10957 INPUT_0 INVX1_LOC_235/Y 0.07fF
C10958 VDD INVX1_LOC_22/Y 0.21fF
C10959 INVX1_LOC_438/A INVX1_LOC_489/A 0.03fF
C10960 INVX1_LOC_558/A INVX1_LOC_586/A 0.07fF
C10961 NAND2X1_LOC_45/Y INVX1_LOC_134/Y 0.12fF
C10962 INVX1_LOC_426/Y INVX1_LOC_145/Y 0.01fF
C10963 NAND2X1_LOC_88/Y INVX1_LOC_205/Y 0.09fF
C10964 INVX1_LOC_578/A INVX1_LOC_119/A 0.08fF
C10965 INVX1_LOC_617/Y INVX1_LOC_557/A 0.39fF
C10966 INVX1_LOC_20/Y INVX1_LOC_160/Y 0.96fF
C10967 NAND2X1_LOC_249/Y INVX1_LOC_145/Y 0.25fF
C10968 INVX1_LOC_625/A INVX1_LOC_560/Y 0.14fF
C10969 NAND2X1_LOC_572/a_36_24# INVX1_LOC_578/A 0.00fF
C10970 VDD INVX1_LOC_504/Y 0.01fF
C10971 INVX1_LOC_564/A INVX1_LOC_635/A 0.36fF
C10972 NAND2X1_LOC_357/a_36_24# INVX1_LOC_45/Y 0.01fF
C10973 NAND2X1_LOC_99/a_36_24# INVX1_LOC_50/Y 0.01fF
C10974 INVX1_LOC_17/Y NAND2X1_LOC_176/Y 0.07fF
C10975 INVX1_LOC_80/A INVX1_LOC_107/A 0.03fF
C10976 INVX1_LOC_566/A INVX1_LOC_51/Y 0.09fF
C10977 INVX1_LOC_573/A INVX1_LOC_571/A 0.08fF
C10978 NAND2X1_LOC_768/A INVX1_LOC_107/A 0.03fF
C10979 NAND2X1_LOC_498/Y INVX1_LOC_134/Y 0.11fF
C10980 INVX1_LOC_417/Y INVX1_LOC_395/A 0.04fF
C10981 INVX1_LOC_570/A INVX1_LOC_134/Y 0.07fF
C10982 INVX1_LOC_239/Y INPUT_1 0.07fF
C10983 NAND2X1_LOC_503/B INVX1_LOC_395/Y 0.20fF
C10984 INVX1_LOC_76/Y INVX1_LOC_196/A 0.01fF
C10985 NAND2X1_LOC_163/a_36_24# INVX1_LOC_147/Y 0.00fF
C10986 INVX1_LOC_206/Y INVX1_LOC_510/A 0.72fF
C10987 INVX1_LOC_661/A INVX1_LOC_651/Y 0.02fF
C10988 INPUT_0 INVX1_LOC_556/Y 0.00fF
C10989 NAND2X1_LOC_513/Y INVX1_LOC_516/A 0.42fF
C10990 INVX1_LOC_446/Y NAND2X1_LOC_275/Y 0.17fF
C10991 NAND2X1_LOC_16/a_36_24# INVX1_LOC_53/Y 0.01fF
C10992 NAND2X1_LOC_13/Y INVX1_LOC_320/A 0.00fF
C10993 INVX1_LOC_378/A INVX1_LOC_489/Y 0.15fF
C10994 INVX1_LOC_160/Y INVX1_LOC_300/A 0.47fF
C10995 INVX1_LOC_160/Y INVX1_LOC_197/Y 0.03fF
C10996 INVX1_LOC_586/A NAND2X1_LOC_755/B 0.15fF
C10997 INVX1_LOC_395/A INVX1_LOC_48/Y 0.20fF
C10998 INVX1_LOC_20/Y INVX1_LOC_358/Y 0.03fF
C10999 INVX1_LOC_522/Y NAND2X1_LOC_513/A 0.51fF
C11000 INVX1_LOC_454/A INVX1_LOC_638/Y 0.01fF
C11001 INVX1_LOC_20/Y INVX1_LOC_21/Y 0.07fF
C11002 NAND2X1_LOC_24/Y INVX1_LOC_42/A 0.00fF
C11003 NAND2X1_LOC_589/a_36_24# INVX1_LOC_117/Y 0.01fF
C11004 INVX1_LOC_134/A NAND2X1_LOC_775/B 0.02fF
C11005 INVX1_LOC_229/Y INVX1_LOC_12/Y 0.03fF
C11006 NAND2X1_LOC_261/Y INVX1_LOC_453/Y 0.03fF
C11007 INVX1_LOC_362/Y INVX1_LOC_48/Y 0.08fF
C11008 INVX1_LOC_425/A INVX1_LOC_416/A 0.53fF
C11009 INVX1_LOC_617/Y INVX1_LOC_468/Y 0.23fF
C11010 INVX1_LOC_425/A INVX1_LOC_419/Y 0.13fF
C11011 INVX1_LOC_54/Y INVX1_LOC_72/Y 0.00fF
C11012 NAND2X1_LOC_325/B INVX1_LOC_80/A 0.09fF
C11013 INVX1_LOC_322/Y INVX1_LOC_50/Y 0.02fF
C11014 NAND2X1_LOC_173/Y INVX1_LOC_259/Y 0.03fF
C11015 INVX1_LOC_502/Y INVX1_LOC_665/Y 0.72fF
C11016 INVX1_LOC_384/Y INVX1_LOC_282/A 0.03fF
C11017 INVX1_LOC_469/Y INVX1_LOC_51/Y 0.03fF
C11018 INVX1_LOC_412/Y NAND2X1_LOC_854/a_36_24# 0.00fF
C11019 INVX1_LOC_312/A INVX1_LOC_17/Y 0.02fF
C11020 NAND2X1_LOC_370/A INVX1_LOC_89/Y 0.01fF
C11021 INVX1_LOC_134/Y INVX1_LOC_99/Y 0.06fF
C11022 INVX1_LOC_447/Y INVX1_LOC_519/A 0.02fF
C11023 INVX1_LOC_249/Y INVX1_LOC_89/Y 0.01fF
C11024 INVX1_LOC_73/Y INVX1_LOC_41/Y 0.01fF
C11025 INVX1_LOC_586/A INVX1_LOC_46/Y 2.27fF
C11026 INVX1_LOC_369/A INVX1_LOC_145/Y 0.03fF
C11027 INVX1_LOC_53/Y INVX1_LOC_549/Y 0.00fF
C11028 INVX1_LOC_516/Y INVX1_LOC_46/Y 0.01fF
C11029 NAND2X1_LOC_537/A INVX1_LOC_100/Y 0.11fF
C11030 INVX1_LOC_658/A NAND2X1_LOC_837/B 0.01fF
C11031 INVX1_LOC_237/Y INVX1_LOC_199/Y 0.03fF
C11032 INVX1_LOC_89/Y NAND2X1_LOC_122/Y 0.01fF
C11033 INVX1_LOC_97/A INVX1_LOC_399/A 0.04fF
C11034 INVX1_LOC_47/A INVX1_LOC_99/Y 0.01fF
C11035 INVX1_LOC_20/Y NAND2X1_LOC_267/A 0.69fF
C11036 INVX1_LOC_21/Y INVX1_LOC_300/A 0.07fF
C11037 INVX1_LOC_335/Y INVX1_LOC_300/A 0.07fF
C11038 INVX1_LOC_257/Y NAND2X1_LOC_605/B 0.02fF
C11039 INVX1_LOC_20/Y NAND2X1_LOC_137/A 0.03fF
C11040 NAND2X1_LOC_373/Y INVX1_LOC_41/Y 0.23fF
C11041 INVX1_LOC_21/Y INVX1_LOC_197/Y 0.03fF
C11042 INVX1_LOC_261/Y INVX1_LOC_677/Y 0.02fF
C11043 NAND2X1_LOC_41/Y INVX1_LOC_99/Y 0.01fF
C11044 NAND2X1_LOC_790/B INVX1_LOC_211/A 0.01fF
C11045 INVX1_LOC_551/Y INVX1_LOC_6/Y 0.00fF
C11046 NAND2X1_LOC_318/A INVX1_LOC_69/Y 0.08fF
C11047 INVX1_LOC_145/Y NAND2X1_LOC_275/Y 0.12fF
C11048 INVX1_LOC_268/Y INVX1_LOC_69/Y 0.03fF
C11049 INVX1_LOC_381/A INVX1_LOC_380/Y 0.06fF
C11050 NAND2X1_LOC_122/Y INVX1_LOC_501/A 0.03fF
C11051 INVX1_LOC_547/Y NAND2X1_LOC_106/a_36_24# 0.00fF
C11052 INVX1_LOC_35/Y INVX1_LOC_1/Y 0.91fF
C11053 INVX1_LOC_504/Y INVX1_LOC_509/A 0.03fF
C11054 INVX1_LOC_205/Y INVX1_LOC_198/A 0.02fF
C11055 INVX1_LOC_11/Y INVX1_LOC_681/A 0.03fF
C11056 INVX1_LOC_80/A NAND2X1_LOC_285/A 0.39fF
C11057 INVX1_LOC_400/Y INVX1_LOC_90/Y 0.08fF
C11058 NAND2X1_LOC_768/A NAND2X1_LOC_285/A 0.01fF
C11059 INVX1_LOC_31/Y INVX1_LOC_632/A 0.09fF
C11060 INVX1_LOC_206/Y NAND2X1_LOC_248/B 0.00fF
C11061 NAND2X1_LOC_108/Y INVX1_LOC_100/Y 0.15fF
C11062 INVX1_LOC_31/Y INVX1_LOC_509/Y 0.01fF
C11063 INVX1_LOC_84/A NAND2X1_LOC_52/Y 0.00fF
C11064 NAND2X1_LOC_165/Y INVX1_LOC_99/Y 0.03fF
C11065 INVX1_LOC_486/Y INVX1_LOC_486/A 0.09fF
C11066 INVX1_LOC_417/Y INVX1_LOC_31/Y 0.10fF
C11067 INVX1_LOC_189/Y INVX1_LOC_48/Y 0.00fF
C11068 INVX1_LOC_47/Y INVX1_LOC_134/Y 0.22fF
C11069 NAND2X1_LOC_791/B NAND2X1_LOC_759/Y 0.02fF
C11070 INVX1_LOC_300/A NAND2X1_LOC_267/A 0.43fF
C11071 INVX1_LOC_79/A NAND2X1_LOC_794/a_36_24# 0.00fF
C11072 INVX1_LOC_272/Y NAND2X1_LOC_759/Y 0.03fF
C11073 NAND2X1_LOC_267/A INVX1_LOC_197/Y 0.07fF
C11074 INVX1_LOC_51/Y INVX1_LOC_79/A 0.28fF
C11075 NAND2X1_LOC_332/B INVX1_LOC_128/Y 0.03fF
C11076 NAND2X1_LOC_48/Y INVX1_LOC_47/Y 0.04fF
C11077 NAND2X1_LOC_529/Y INVX1_LOC_46/Y 0.09fF
C11078 INVX1_LOC_46/Y NAND2X1_LOC_378/Y 0.04fF
C11079 INVX1_LOC_47/A INVX1_LOC_47/Y 0.01fF
C11080 NAND2X1_LOC_513/A INVX1_LOC_508/A 0.12fF
C11081 NAND2X1_LOC_775/B INVX1_LOC_50/Y 0.02fF
C11082 INVX1_LOC_31/Y INVX1_LOC_59/Y 0.18fF
C11083 INVX1_LOC_412/A INVX1_LOC_666/Y 0.03fF
C11084 INVX1_LOC_29/A INPUT_4 0.24fF
C11085 INVX1_LOC_11/Y NAND2X1_LOC_482/Y 0.35fF
C11086 INVX1_LOC_51/Y INVX1_LOC_460/A 0.08fF
C11087 INVX1_LOC_342/Y INVX1_LOC_340/A 0.94fF
C11088 INVX1_LOC_69/Y INVX1_LOC_115/A 0.03fF
C11089 NAND2X1_LOC_755/B NAND2X1_LOC_825/a_36_24# 0.00fF
C11090 NAND2X1_LOC_492/a_36_24# INVX1_LOC_319/A 0.00fF
C11091 INVX1_LOC_248/Y INVX1_LOC_154/A 0.01fF
C11092 NAND2X1_LOC_13/Y INVX1_LOC_100/Y 1.76fF
C11093 INVX1_LOC_266/A INVX1_LOC_79/A 0.03fF
C11094 INVX1_LOC_69/Y INVX1_LOC_363/Y 0.01fF
C11095 INVX1_LOC_32/Y NAND2X1_LOC_615/B 0.46fF
C11096 INVX1_LOC_575/A NAND2X1_LOC_611/a_36_24# 0.02fF
C11097 INVX1_LOC_31/Y INVX1_LOC_48/Y 0.76fF
C11098 INVX1_LOC_202/Y INVX1_LOC_69/Y 0.03fF
C11099 INVX1_LOC_338/A INVX1_LOC_58/Y 0.01fF
C11100 INVX1_LOC_69/Y INVX1_LOC_349/Y 0.01fF
C11101 INVX1_LOC_53/Y NAND2X1_LOC_274/B 0.07fF
C11102 INVX1_LOC_214/Y INVX1_LOC_58/Y 0.14fF
C11103 INVX1_LOC_63/Y INVX1_LOC_506/Y 0.04fF
C11104 INVX1_LOC_134/Y INVX1_LOC_119/Y 0.13fF
C11105 GATE_811 INVX1_LOC_641/Y 0.01fF
C11106 INVX1_LOC_159/Y INVX1_LOC_199/Y 0.07fF
C11107 INVX1_LOC_573/Y INVX1_LOC_137/Y 0.01fF
C11108 NAND2X1_LOC_675/B INVX1_LOC_48/Y 0.07fF
C11109 INVX1_LOC_32/Y INVX1_LOC_66/A 0.03fF
C11110 INVX1_LOC_63/Y NAND2X1_LOC_646/A 0.27fF
C11111 INVX1_LOC_686/A INVX1_LOC_66/Y 0.01fF
C11112 INVX1_LOC_17/Y INVX1_LOC_226/Y 0.01fF
C11113 INVX1_LOC_183/A NAND2X1_LOC_673/B 0.02fF
C11114 INVX1_LOC_35/Y INVX1_LOC_245/A 0.10fF
C11115 INVX1_LOC_21/Y NAND2X1_LOC_269/B 0.01fF
C11116 NAND2X1_LOC_307/B INVX1_LOC_523/Y 0.01fF
C11117 INVX1_LOC_387/Y INVX1_LOC_69/Y 0.03fF
C11118 INVX1_LOC_117/Y INVX1_LOC_507/Y 0.01fF
C11119 INVX1_LOC_356/A NAND2X1_LOC_428/a_36_24# 0.01fF
C11120 INVX1_LOC_366/A NAND2X1_LOC_793/a_36_24# 0.00fF
C11121 INVX1_LOC_317/Y INVX1_LOC_92/A 0.07fF
C11122 NAND2X1_LOC_336/B INVX1_LOC_666/Y 0.03fF
C11123 NAND2X1_LOC_140/B INVX1_LOC_41/Y 0.54fF
C11124 NAND2X1_LOC_41/Y NAND2X1_LOC_66/Y 0.03fF
C11125 INVX1_LOC_261/Y INVX1_LOC_638/Y 0.01fF
C11126 INVX1_LOC_6/Y INVX1_LOC_486/A 0.02fF
C11127 INVX1_LOC_319/A INVX1_LOC_230/A 0.09fF
C11128 INVX1_LOC_199/Y INVX1_LOC_212/Y 0.07fF
C11129 INVX1_LOC_598/A INVX1_LOC_26/Y 0.06fF
C11130 INVX1_LOC_253/Y INVX1_LOC_63/Y 0.01fF
C11131 INVX1_LOC_49/Y INVX1_LOC_69/Y 1.39fF
C11132 INVX1_LOC_635/A INVX1_LOC_91/Y 0.00fF
C11133 NAND2X1_LOC_725/a_36_24# INVX1_LOC_92/A 0.00fF
C11134 NAND2X1_LOC_448/B INVX1_LOC_245/A 0.01fF
C11135 INVX1_LOC_368/A INVX1_LOC_490/A 0.01fF
C11136 INVX1_LOC_53/Y NAND2X1_LOC_245/a_36_24# 0.00fF
C11137 INVX1_LOC_555/A INVX1_LOC_655/A 0.87fF
C11138 INVX1_LOC_354/A INVX1_LOC_259/Y 0.01fF
C11139 NAND2X1_LOC_274/B NAND2X1_LOC_274/Y 0.06fF
C11140 NAND2X1_LOC_531/Y INVX1_LOC_422/A 0.35fF
C11141 INVX1_LOC_373/Y INVX1_LOC_338/Y 0.01fF
C11142 NAND2X1_LOC_184/Y INVX1_LOC_479/A 3.03fF
C11143 INVX1_LOC_183/Y INVX1_LOC_9/Y 0.19fF
C11144 INVX1_LOC_446/A NAND2X1_LOC_573/a_36_24# 0.00fF
C11145 INVX1_LOC_6/Y NAND2X1_LOC_410/Y 0.02fF
C11146 INVX1_LOC_199/Y INVX1_LOC_468/A 0.01fF
C11147 NAND2X1_LOC_249/Y NAND2X1_LOC_595/a_36_24# 0.00fF
C11148 INVX1_LOC_26/Y INVX1_LOC_242/Y 0.06fF
C11149 INVX1_LOC_41/Y INVX1_LOC_494/Y 0.01fF
C11150 NAND2X1_LOC_691/A INVX1_LOC_338/Y 0.01fF
C11151 INVX1_LOC_612/Y INVX1_LOC_613/A 0.44fF
C11152 INVX1_LOC_74/Y INVX1_LOC_361/A 0.01fF
C11153 VDD INVX1_LOC_278/A 0.06fF
C11154 INVX1_LOC_479/A INVX1_LOC_498/Y 0.07fF
C11155 NAND2X1_LOC_274/B NAND2X1_LOC_844/a_36_24# 0.00fF
C11156 INVX1_LOC_166/A INVX1_LOC_92/A 0.03fF
C11157 INVX1_LOC_224/Y INVX1_LOC_410/Y 0.07fF
C11158 INVX1_LOC_223/A INVX1_LOC_9/Y 0.05fF
C11159 VDD INVX1_LOC_542/A -0.00fF
C11160 INVX1_LOC_377/A INVX1_LOC_109/Y 0.06fF
C11161 INPUT_6 INVX1_LOC_4/Y 0.01fF
C11162 INVX1_LOC_578/A INVX1_LOC_410/Y 0.45fF
C11163 NAND2X1_LOC_528/Y INVX1_LOC_75/Y 0.06fF
C11164 INVX1_LOC_557/A INVX1_LOC_375/A 0.04fF
C11165 INVX1_LOC_577/A INVX1_LOC_51/Y 0.00fF
C11166 INVX1_LOC_21/Y INVX1_LOC_73/Y 0.01fF
C11167 INVX1_LOC_426/A INVX1_LOC_417/Y 0.10fF
C11168 INVX1_LOC_20/Y NAND2X1_LOC_710/B 0.10fF
C11169 INVX1_LOC_617/Y INVX1_LOC_206/Y 0.07fF
C11170 NAND2X1_LOC_331/A INVX1_LOC_147/Y 0.01fF
C11171 INVX1_LOC_412/Y INVX1_LOC_686/A 0.07fF
C11172 INVX1_LOC_287/A INVX1_LOC_560/Y 0.21fF
C11173 NAND2X1_LOC_596/a_36_24# NAND2X1_LOC_596/Y 0.00fF
C11174 INVX1_LOC_20/Y INVX1_LOC_255/Y 0.04fF
C11175 INVX1_LOC_446/Y INVX1_LOC_235/Y 0.02fF
C11176 INVX1_LOC_268/Y INVX1_LOC_586/A 0.04fF
C11177 VDD INVX1_LOC_453/Y 1.85fF
C11178 INVX1_LOC_84/A INVX1_LOC_65/Y 0.44fF
C11179 INPUT_6 INVX1_LOC_56/Y 0.01fF
C11180 INVX1_LOC_438/Y INVX1_LOC_7/Y 0.05fF
C11181 NAND2X1_LOC_685/A INVX1_LOC_45/Y 0.03fF
C11182 INVX1_LOC_133/A INVX1_LOC_242/A 0.21fF
C11183 INVX1_LOC_429/A INVX1_LOC_386/Y 0.08fF
C11184 VDD INVX1_LOC_259/Y 1.08fF
C11185 NAND2X1_LOC_331/A INVX1_LOC_511/Y 0.03fF
C11186 INVX1_LOC_617/Y INVX1_LOC_242/A 0.01fF
C11187 INVX1_LOC_567/A INVX1_LOC_46/Y 0.00fF
C11188 INVX1_LOC_202/A INVX1_LOC_31/Y 0.01fF
C11189 INVX1_LOC_45/Y INVX1_LOC_188/Y 0.03fF
C11190 INVX1_LOC_373/A INVX1_LOC_145/Y 0.06fF
C11191 NAND2X1_LOC_498/Y INVX1_LOC_370/Y 0.01fF
C11192 NAND2X1_LOC_184/a_36_24# INVX1_LOC_50/Y 0.01fF
C11193 INVX1_LOC_603/Y INVX1_LOC_45/Y 0.03fF
C11194 INVX1_LOC_468/Y INVX1_LOC_375/A 0.02fF
C11195 INVX1_LOC_502/Y INVX1_LOC_134/Y 0.00fF
C11196 INVX1_LOC_51/Y INVX1_LOC_632/A 0.47fF
C11197 INVX1_LOC_468/Y INVX1_LOC_546/A 0.00fF
C11198 INVX1_LOC_563/A INVX1_LOC_586/A 0.02fF
C11199 NAND2X1_LOC_310/a_36_24# NAND2X1_LOC_267/A 0.01fF
C11200 INVX1_LOC_686/A INVX1_LOC_119/A 0.04fF
C11201 VDD NAND2X1_LOC_707/B 0.14fF
C11202 INVX1_LOC_6/Y INVX1_LOC_596/Y 0.00fF
C11203 NAND2X1_LOC_142/Y NAND2X1_LOC_285/B 0.02fF
C11204 NAND2X1_LOC_249/Y NAND2X1_LOC_128/B 0.05fF
C11205 INVX1_LOC_374/A INVX1_LOC_506/Y 0.01fF
C11206 NAND2X1_LOC_598/a_36_24# INVX1_LOC_47/Y 0.01fF
C11207 VDD INVX1_LOC_204/Y 0.53fF
C11208 NAND2X1_LOC_503/B INVX1_LOC_44/Y 0.02fF
C11209 INVX1_LOC_587/A NAND2X1_LOC_755/B 0.03fF
C11210 NAND2X1_LOC_637/A INVX1_LOC_49/Y 0.03fF
C11211 INVX1_LOC_51/Y INVX1_LOC_59/Y 0.03fF
C11212 NAND2X1_LOC_142/Y NAND2X1_LOC_106/B 0.01fF
C11213 INVX1_LOC_202/Y INVX1_LOC_586/A 0.07fF
C11214 INVX1_LOC_435/Y INVX1_LOC_221/Y 0.07fF
C11215 INVX1_LOC_561/Y INVX1_LOC_31/Y 0.28fF
C11216 NAND2X1_LOC_505/Y INVX1_LOC_48/Y 0.03fF
C11217 INVX1_LOC_677/Y INVX1_LOC_290/A 0.23fF
C11218 NAND2X1_LOC_331/A INVX1_LOC_538/A 0.09fF
C11219 INVX1_LOC_586/A INVX1_LOC_349/Y 0.01fF
C11220 INVX1_LOC_134/Y INVX1_LOC_136/Y 0.01fF
C11221 INVX1_LOC_618/A INVX1_LOC_79/A 0.24fF
C11222 INVX1_LOC_51/Y INVX1_LOC_48/Y 0.12fF
C11223 NAND2X1_LOC_791/B NAND2X1_LOC_755/B 0.01fF
C11224 NAND2X1_LOC_387/Y NAND2X1_LOC_506/B 0.03fF
C11225 INVX1_LOC_524/Y NAND2X1_LOC_93/a_36_24# 0.00fF
C11226 INVX1_LOC_235/Y INVX1_LOC_145/Y 0.11fF
C11227 INVX1_LOC_272/Y NAND2X1_LOC_755/B 0.15fF
C11228 INVX1_LOC_442/A INVX1_LOC_32/Y 0.14fF
C11229 NAND2X1_LOC_387/Y INVX1_LOC_45/Y 0.68fF
C11230 INVX1_LOC_312/Y INVX1_LOC_363/Y 0.05fF
C11231 VDD INVX1_LOC_82/Y 0.04fF
C11232 INVX1_LOC_106/A INVX1_LOC_679/Y 0.01fF
C11233 INVX1_LOC_617/A INVX1_LOC_665/Y 0.00fF
C11234 INVX1_LOC_211/Y INVX1_LOC_486/Y 0.02fF
C11235 INVX1_LOC_570/A INVX1_LOC_476/A 0.05fF
C11236 INVX1_LOC_117/Y INVX1_LOC_163/Y 0.01fF
C11237 INVX1_LOC_99/Y INVX1_LOC_16/Y 0.01fF
C11238 INVX1_LOC_558/A INVX1_LOC_6/Y 0.57fF
C11239 VDD INVX1_LOC_114/A 1.72fF
C11240 INVX1_LOC_21/Y INVX1_LOC_600/Y 0.05fF
C11241 INVX1_LOC_552/Y INVX1_LOC_63/Y 0.01fF
C11242 INVX1_LOC_305/Y INVX1_LOC_7/Y 0.03fF
C11243 INVX1_LOC_266/A INVX1_LOC_48/Y 0.05fF
C11244 INVX1_LOC_387/Y INVX1_LOC_586/A 0.00fF
C11245 INVX1_LOC_382/A INVX1_LOC_378/A 0.03fF
C11246 NAND2X1_LOC_45/Y INVX1_LOC_90/Y 0.05fF
C11247 INVX1_LOC_117/Y INVX1_LOC_522/Y 0.14fF
C11248 INVX1_LOC_344/Y INVX1_LOC_504/A 0.02fF
C11249 INVX1_LOC_337/Y INVX1_LOC_50/Y 0.01fF
C11250 INVX1_LOC_374/A INVX1_LOC_63/Y 0.04fF
C11251 INVX1_LOC_53/Y INVX1_LOC_159/Y 0.01fF
C11252 NAND2X1_LOC_596/Y INVX1_LOC_114/A 0.01fF
C11253 INVX1_LOC_586/A INVX1_LOC_49/Y 0.30fF
C11254 INVX1_LOC_316/Y INVX1_LOC_25/Y 0.01fF
C11255 INVX1_LOC_560/A INVX1_LOC_242/Y 0.02fF
C11256 INVX1_LOC_50/Y INVX1_LOC_633/Y 0.03fF
C11257 INVX1_LOC_76/Y INVX1_LOC_69/Y 0.10fF
C11258 INVX1_LOC_340/Y INVX1_LOC_675/A 0.07fF
C11259 NAND2X1_LOC_782/A INVX1_LOC_53/Y 0.16fF
C11260 INVX1_LOC_123/A INVX1_LOC_318/Y 0.02fF
C11261 INVX1_LOC_268/Y INVX1_LOC_157/Y 0.08fF
C11262 INVX1_LOC_17/Y INVX1_LOC_252/Y 0.03fF
C11263 NAND2X1_LOC_478/a_36_24# INVX1_LOC_510/A 0.01fF
C11264 INVX1_LOC_312/A INVX1_LOC_230/Y 0.01fF
C11265 NAND2X1_LOC_820/A INVX1_LOC_46/Y 0.01fF
C11266 INVX1_LOC_273/A INVX1_LOC_44/Y 0.03fF
C11267 INVX1_LOC_80/A INVX1_LOC_355/Y 0.01fF
C11268 INVX1_LOC_81/Y INVX1_LOC_145/Y 0.00fF
C11269 NAND2X1_LOC_41/Y NAND2X1_LOC_43/Y 0.08fF
C11270 INVX1_LOC_45/Y NAND2X1_LOC_845/B 0.00fF
C11271 INVX1_LOC_36/A INVX1_LOC_90/Y 0.01fF
C11272 INVX1_LOC_533/Y INVX1_LOC_26/Y 0.00fF
C11273 NAND2X1_LOC_556/a_36_24# INVX1_LOC_453/Y 0.06fF
C11274 NAND2X1_LOC_399/B INVX1_LOC_328/A 0.04fF
C11275 INVX1_LOC_100/A INVX1_LOC_307/A 0.12fF
C11276 INVX1_LOC_355/A INVX1_LOC_79/A 0.01fF
C11277 INVX1_LOC_579/A INVX1_LOC_89/Y 0.01fF
C11278 INVX1_LOC_117/Y NAND2X1_LOC_448/A 0.02fF
C11279 INVX1_LOC_11/Y INVX1_LOC_137/Y 0.02fF
C11280 INVX1_LOC_7/Y INVX1_LOC_328/A 0.02fF
C11281 INVX1_LOC_93/Y INVX1_LOC_155/Y 0.03fF
C11282 INVX1_LOC_649/Y NAND2X1_LOC_846/A 0.01fF
C11283 INVX1_LOC_312/Y INVX1_LOC_49/Y 0.07fF
C11284 NAND2X1_LOC_13/Y NAND2X1_LOC_558/B 0.01fF
C11285 INVX1_LOC_254/A INVX1_LOC_59/Y 0.00fF
C11286 NAND2X1_LOC_313/a_36_24# INVX1_LOC_251/Y 0.00fF
C11287 INVX1_LOC_32/Y INVX1_LOC_116/Y 0.07fF
C11288 NAND2X1_LOC_834/a_36_24# INVX1_LOC_6/Y -0.00fF
C11289 INVX1_LOC_107/A NAND2X1_LOC_843/B 0.01fF
C11290 INVX1_LOC_428/A INVX1_LOC_62/Y 0.03fF
C11291 INVX1_LOC_20/Y NAND2X1_LOC_420/a_36_24# 0.00fF
C11292 INVX1_LOC_536/A INVX1_LOC_58/Y 0.03fF
C11293 INVX1_LOC_370/Y INVX1_LOC_47/Y 0.06fF
C11294 INVX1_LOC_20/Y INVX1_LOC_26/Y 0.18fF
C11295 NAND2X1_LOC_755/B INVX1_LOC_6/Y 0.03fF
C11296 INVX1_LOC_586/A INVX1_LOC_17/A 0.01fF
C11297 INVX1_LOC_551/A INVX1_LOC_12/Y 0.00fF
C11298 NAND2X1_LOC_13/Y INVX1_LOC_79/A 0.00fF
C11299 INVX1_LOC_672/A INVX1_LOC_283/A 0.17fF
C11300 INVX1_LOC_607/A INVX1_LOC_479/A 0.04fF
C11301 INVX1_LOC_117/Y INVX1_LOC_295/Y 0.04fF
C11302 INVX1_LOC_484/A INVX1_LOC_480/Y 0.17fF
C11303 INVX1_LOC_211/Y INVX1_LOC_6/Y 0.01fF
C11304 INVX1_LOC_562/Y INVX1_LOC_41/Y 0.01fF
C11305 INVX1_LOC_20/Y NAND2X1_LOC_210/a_36_24# 0.01fF
C11306 INVX1_LOC_78/A INVX1_LOC_338/Y 0.05fF
C11307 INVX1_LOC_166/A INPUT_1 0.11fF
C11308 INVX1_LOC_369/A INVX1_LOC_484/Y 0.01fF
C11309 NAND2X1_LOC_165/Y INVX1_LOC_153/A 0.10fF
C11310 NAND2X1_LOC_775/B NAND2X1_LOC_388/A 0.03fF
C11311 INVX1_LOC_576/A INVX1_LOC_26/Y 0.00fF
C11312 INVX1_LOC_32/Y INVX1_LOC_328/A 0.02fF
C11313 NAND2X1_LOC_542/A INVX1_LOC_510/A 0.07fF
C11314 INVX1_LOC_419/Y INVX1_LOC_419/A 0.01fF
C11315 NAND2X1_LOC_616/Y NAND2X1_LOC_616/a_36_24# 0.01fF
C11316 NAND2X1_LOC_399/a_36_24# INVX1_LOC_63/Y 0.00fF
C11317 NAND2X1_LOC_531/Y INVX1_LOC_8/Y 0.00fF
C11318 INVX1_LOC_300/A NAND2X1_LOC_290/a_36_24# 0.00fF
C11319 INVX1_LOC_520/Y INVX1_LOC_35/Y 0.01fF
C11320 NAND2X1_LOC_486/B INVX1_LOC_479/A 0.33fF
C11321 NAND2X1_LOC_517/Y NAND2X1_LOC_642/a_36_24# 0.00fF
C11322 NAND2X1_LOC_184/Y NAND2X1_LOC_521/Y 0.22fF
C11323 INVX1_LOC_99/Y INVX1_LOC_351/A 0.01fF
C11324 INVX1_LOC_484/A INVX1_LOC_169/Y 0.09fF
C11325 INVX1_LOC_223/Y INVX1_LOC_178/A 0.19fF
C11326 INVX1_LOC_6/Y INVX1_LOC_46/Y 0.13fF
C11327 INVX1_LOC_183/Y INVX1_LOC_42/Y 0.01fF
C11328 INVX1_LOC_93/Y INVX1_LOC_633/A 0.00fF
C11329 NAND2X1_LOC_503/Y INVX1_LOC_69/Y 0.31fF
C11330 INVX1_LOC_300/A INVX1_LOC_26/Y 0.07fF
C11331 INVX1_LOC_53/Y INVX1_LOC_468/A 0.45fF
C11332 INVX1_LOC_376/Y INVX1_LOC_510/A 0.14fF
C11333 INVX1_LOC_255/A INVX1_LOC_32/Y 0.07fF
C11334 INVX1_LOC_99/Y INVX1_LOC_90/Y 0.12fF
C11335 INVX1_LOC_26/Y INVX1_LOC_197/Y 0.03fF
C11336 NAND2X1_LOC_433/Y INVX1_LOC_137/Y 0.25fF
C11337 INVX1_LOC_172/A INVX1_LOC_328/Y 0.04fF
C11338 INVX1_LOC_509/A INVX1_LOC_114/A 0.00fF
C11339 INVX1_LOC_338/Y INVX1_LOC_496/Y 0.01fF
C11340 INVX1_LOC_12/Y INVX1_LOC_75/Y 0.24fF
C11341 INVX1_LOC_31/Y NAND2X1_LOC_615/Y 0.22fF
C11342 INVX1_LOC_242/Y INVX1_LOC_603/A 0.02fF
C11343 INVX1_LOC_32/Y INVX1_LOC_179/A 0.07fF
C11344 INVX1_LOC_209/Y INVX1_LOC_600/Y 0.01fF
C11345 INVX1_LOC_63/Y NAND2X1_LOC_836/B 0.05fF
C11346 INVX1_LOC_293/A INVX1_LOC_654/Y 0.00fF
C11347 NAND2X1_LOC_148/A NAND2X1_LOC_245/a_36_24# 0.00fF
C11348 INVX1_LOC_53/Y INVX1_LOC_620/Y 0.08fF
C11349 INVX1_LOC_394/Y NAND2X1_LOC_503/B 0.00fF
C11350 INVX1_LOC_507/Y INVX1_LOC_58/Y 0.01fF
C11351 INVX1_LOC_409/Y INVX1_LOC_638/A 0.01fF
C11352 INVX1_LOC_223/Y INVX1_LOC_58/Y 0.01fF
C11353 INVX1_LOC_47/Y INVX1_LOC_90/Y 0.10fF
C11354 INVX1_LOC_346/A INVX1_LOC_114/A 0.01fF
C11355 NAND2X1_LOC_633/a_36_24# INVX1_LOC_496/A 0.00fF
C11356 NAND2X1_LOC_136/Y NAND2X1_LOC_279/a_36_24# 0.00fF
C11357 INVX1_LOC_531/Y INVX1_LOC_292/Y 0.14fF
C11358 INVX1_LOC_359/A INVX1_LOC_74/Y 0.01fF
C11359 INVX1_LOC_79/A INVX1_LOC_361/A 0.00fF
C11360 NAND2X1_LOC_285/A NAND2X1_LOC_843/B 0.02fF
C11361 INVX1_LOC_328/Y INVX1_LOC_224/A 0.00fF
C11362 NAND2X1_LOC_451/B INVX1_LOC_340/A 0.03fF
C11363 NAND2X1_LOC_69/B INVX1_LOC_395/A 0.03fF
C11364 VDD INVX1_LOC_554/Y 0.24fF
C11365 INVX1_LOC_496/A INVX1_LOC_588/A 0.08fF
C11366 INVX1_LOC_301/A INVX1_LOC_560/A 0.03fF
C11367 INVX1_LOC_513/Y INVX1_LOC_479/A 0.01fF
C11368 INVX1_LOC_483/Y INVX1_LOC_480/A 0.01fF
C11369 NAND2X1_LOC_710/B INVX1_LOC_553/A 0.01fF
C11370 VDD INVX1_LOC_547/Y 0.35fF
C11371 INVX1_LOC_206/Y INVX1_LOC_410/Y 0.01fF
C11372 NAND2X1_LOC_176/Y NAND2X1_LOC_370/A 0.00fF
C11373 INVX1_LOC_206/Y INVX1_LOC_375/A 0.03fF
C11374 NAND2X1_LOC_123/B INVX1_LOC_41/Y 0.03fF
C11375 VDD INVX1_LOC_499/Y 0.05fF
C11376 INVX1_LOC_554/A NAND2X1_LOC_159/a_36_24# 0.01fF
C11377 NAND2X1_LOC_183/a_36_24# INVX1_LOC_362/Y 0.00fF
C11378 INVX1_LOC_245/A INVX1_LOC_488/Y 0.02fF
C11379 INVX1_LOC_627/A NAND2X1_LOC_513/A 0.01fF
C11380 INVX1_LOC_92/A INVX1_LOC_411/Y 0.31fF
C11381 INVX1_LOC_133/Y NAND2X1_LOC_513/A 1.17fF
C11382 INVX1_LOC_266/A NAND2X1_LOC_370/a_36_24# 0.07fF
C11383 INVX1_LOC_438/A NAND2X1_LOC_613/Y 0.02fF
C11384 INVX1_LOC_510/Y NAND2X1_LOC_314/a_36_24# 0.00fF
C11385 NAND2X1_LOC_331/Y NAND2X1_LOC_801/A 0.00fF
C11386 VDD INVX1_LOC_439/A -0.00fF
C11387 NAND2X1_LOC_513/Y INVX1_LOC_51/Y 0.01fF
C11388 INVX1_LOC_438/Y INVX1_LOC_424/Y 0.11fF
C11389 INVX1_LOC_41/Y INVX1_LOC_270/Y 0.12fF
C11390 NAND2X1_LOC_475/A INVX1_LOC_318/Y 0.00fF
C11391 INVX1_LOC_375/A INVX1_LOC_242/A 0.12fF
C11392 INVX1_LOC_98/A INVX1_LOC_586/A 1.11fF
C11393 INVX1_LOC_428/A INVX1_LOC_547/A 0.03fF
C11394 NAND2X1_LOC_710/A INVX1_LOC_395/A 0.01fF
C11395 INVX1_LOC_410/Y INVX1_LOC_686/A 0.42fF
C11396 INVX1_LOC_395/A INVX1_LOC_508/Y 0.02fF
C11397 INVX1_LOC_41/Y INVX1_LOC_92/A 0.03fF
C11398 INVX1_LOC_76/Y INVX1_LOC_586/A 0.19fF
C11399 INVX1_LOC_308/Y INVX1_LOC_307/A 0.21fF
C11400 INVX1_LOC_76/Y INVX1_LOC_516/Y 0.01fF
C11401 INVX1_LOC_174/Y INVX1_LOC_184/A 0.06fF
C11402 NAND2X1_LOC_69/B INVX1_LOC_31/Y 0.01fF
C11403 INVX1_LOC_121/Y INVX1_LOC_510/A 0.03fF
C11404 NAND2X1_LOC_704/a_36_24# INVX1_LOC_251/Y 0.00fF
C11405 INVX1_LOC_254/Y INVX1_LOC_224/Y 0.07fF
C11406 VDD INVX1_LOC_87/Y 0.26fF
C11407 INVX1_LOC_206/Y INVX1_LOC_674/A 0.07fF
C11408 NAND2X1_LOC_525/Y INVX1_LOC_367/Y 0.68fF
C11409 NAND2X1_LOC_498/Y INVX1_LOC_98/Y 0.10fF
C11410 INVX1_LOC_405/A INVX1_LOC_63/Y 0.03fF
C11411 INVX1_LOC_570/A INVX1_LOC_98/Y 0.07fF
C11412 INVX1_LOC_185/A INVX1_LOC_508/A 0.27fF
C11413 INVX1_LOC_335/Y INVX1_LOC_562/Y 0.03fF
C11414 NAND2X1_LOC_519/a_36_24# NAND2X1_LOC_275/Y 0.00fF
C11415 INVX1_LOC_45/Y INVX1_LOC_504/Y 0.07fF
C11416 NAND2X1_LOC_457/A INVX1_LOC_103/Y 0.03fF
C11417 INVX1_LOC_438/A INVX1_LOC_490/A 0.09fF
C11418 INPUT_0 NAND2X1_LOC_191/a_36_24# 0.00fF
C11419 INVX1_LOC_32/A INVX1_LOC_6/Y 0.01fF
C11420 INVX1_LOC_398/A INVX1_LOC_600/A 0.03fF
C11421 NAND2X1_LOC_307/A INVX1_LOC_80/A 0.03fF
C11422 INVX1_LOC_560/Y INVX1_LOC_63/Y 0.03fF
C11423 INVX1_LOC_80/A INVX1_LOC_545/Y 0.09fF
C11424 INVX1_LOC_321/A INVX1_LOC_432/A 0.02fF
C11425 INVX1_LOC_556/Y NAND2X1_LOC_332/B 0.01fF
C11426 INVX1_LOC_435/Y INVX1_LOC_421/A 0.10fF
C11427 INVX1_LOC_581/A NAND2X1_LOC_513/A 0.03fF
C11428 INVX1_LOC_395/A INVX1_LOC_633/A 0.02fF
C11429 NAND2X1_LOC_523/B INVX1_LOC_99/Y 0.01fF
C11430 INVX1_LOC_406/Y INVX1_LOC_452/A 0.03fF
C11431 INVX1_LOC_366/A NAND2X1_LOC_222/a_36_24# 0.01fF
C11432 INVX1_LOC_556/Y INVX1_LOC_125/Y 0.01fF
C11433 INVX1_LOC_190/Y INVX1_LOC_44/Y 0.09fF
C11434 NAND2X1_LOC_13/Y INVX1_LOC_48/Y 0.04fF
C11435 NAND2X1_LOC_545/B INVX1_LOC_99/Y 0.02fF
C11436 INVX1_LOC_51/Y INVX1_LOC_559/Y 0.01fF
C11437 INVX1_LOC_288/A NAND2X1_LOC_453/a_36_24# 0.00fF
C11438 INVX1_LOC_20/Y INVX1_LOC_603/A 0.03fF
C11439 NAND2X1_LOC_786/a_36_24# NAND2X1_LOC_243/A -0.00fF
C11440 INVX1_LOC_455/Y INVX1_LOC_25/Y 0.19fF
C11441 VDD INVX1_LOC_422/A -0.00fF
C11442 NAND2X1_LOC_322/a_36_24# INPUT_1 0.01fF
C11443 INVX1_LOC_11/Y NAND2X1_LOC_307/A 0.02fF
C11444 INVX1_LOC_310/Y INVX1_LOC_145/Y 0.03fF
C11445 NAND2X1_LOC_486/B INVX1_LOC_391/A 0.10fF
C11446 INVX1_LOC_288/A NAND2X1_LOC_586/Y 0.03fF
C11447 NAND2X1_LOC_756/Y NAND2X1_LOC_387/Y 0.09fF
C11448 INVX1_LOC_570/A INVX1_LOC_338/Y 0.07fF
C11449 NAND2X1_LOC_475/A INVX1_LOC_90/Y 0.00fF
C11450 NAND2X1_LOC_231/A INVX1_LOC_94/Y 0.14fF
C11451 INVX1_LOC_340/Y INVX1_LOC_641/A 0.32fF
C11452 INVX1_LOC_20/Y NAND2X1_LOC_309/a_36_24# 0.00fF
C11453 INVX1_LOC_99/Y INVX1_LOC_98/Y 0.09fF
C11454 INVX1_LOC_114/Y INVX1_LOC_497/A 0.02fF
C11455 INVX1_LOC_31/Y INVX1_LOC_634/A 0.02fF
C11456 INVX1_LOC_31/Y NAND2X1_LOC_541/B 0.31fF
C11457 INVX1_LOC_300/A NAND2X1_LOC_211/a_36_24# 0.00fF
C11458 INVX1_LOC_163/Y INVX1_LOC_58/Y 0.15fF
C11459 INVX1_LOC_617/Y NAND2X1_LOC_542/A 0.07fF
C11460 INVX1_LOC_558/A INVX1_LOC_557/Y 0.03fF
C11461 INVX1_LOC_224/Y NAND2X1_LOC_528/Y 0.15fF
C11462 INVX1_LOC_142/Y INVX1_LOC_168/Y 0.04fF
C11463 NAND2X1_LOC_13/Y NAND2X1_LOC_491/Y 0.01fF
C11464 INVX1_LOC_300/A INVX1_LOC_603/A 0.02fF
C11465 INVX1_LOC_224/Y INVX1_LOC_479/A 0.07fF
C11466 INVX1_LOC_51/A INVX1_LOC_62/Y 0.00fF
C11467 INVX1_LOC_599/Y INVX1_LOC_601/Y 0.03fF
C11468 INVX1_LOC_84/A INVX1_LOC_63/Y 0.24fF
C11469 INVX1_LOC_80/A NAND2X1_LOC_342/A 0.00fF
C11470 INVX1_LOC_21/Y NAND2X1_LOC_106/Y 0.00fF
C11471 INVX1_LOC_591/Y INVX1_LOC_63/Y 0.01fF
C11472 NAND2X1_LOC_670/a_36_24# INVX1_LOC_48/Y 0.00fF
C11473 INVX1_LOC_617/Y INVX1_LOC_376/Y 0.02fF
C11474 INVX1_LOC_20/Y NAND2X1_LOC_605/B 0.02fF
C11475 NAND2X1_LOC_775/B NAND2X1_LOC_112/a_36_24# 0.01fF
C11476 INVX1_LOC_654/A INVX1_LOC_664/A 0.03fF
C11477 INVX1_LOC_578/A INVX1_LOC_479/A 0.07fF
C11478 INVX1_LOC_492/A INVX1_LOC_138/Y 0.00fF
C11479 INVX1_LOC_80/A INVX1_LOC_376/A 0.07fF
C11480 NAND2X1_LOC_142/Y NAND2X1_LOC_248/B 0.15fF
C11481 INVX1_LOC_557/A INVX1_LOC_479/A 0.01fF
C11482 INVX1_LOC_366/A INVX1_LOC_210/A 0.04fF
C11483 INVX1_LOC_588/Y INVX1_LOC_50/Y 0.01fF
C11484 INVX1_LOC_551/Y INVX1_LOC_100/Y 2.35fF
C11485 INVX1_LOC_47/Y INVX1_LOC_98/Y 0.10fF
C11486 INVX1_LOC_415/Y INVX1_LOC_46/Y 0.28fF
C11487 INVX1_LOC_145/Y NAND2X1_LOC_586/Y 0.15fF
C11488 INVX1_LOC_35/Y NAND2X1_LOC_753/Y 0.17fF
C11489 INVX1_LOC_99/Y INVX1_LOC_338/Y 0.03fF
C11490 INVX1_LOC_166/A INVX1_LOC_50/Y 0.07fF
C11491 INVX1_LOC_555/A NAND2X1_LOC_696/a_36_24# 0.00fF
C11492 INVX1_LOC_49/Y INVX1_LOC_252/A 0.02fF
C11493 INVX1_LOC_6/Y INVX1_LOC_381/Y 0.03fF
C11494 INVX1_LOC_63/Y NAND2X1_LOC_67/Y 0.00fF
C11495 INVX1_LOC_59/Y INVX1_LOC_361/A 0.01fF
C11496 INVX1_LOC_128/A INVX1_LOC_383/Y 0.00fF
C11497 INVX1_LOC_128/Y INVX1_LOC_375/Y 0.06fF
C11498 INVX1_LOC_550/A INVX1_LOC_6/Y 0.01fF
C11499 INVX1_LOC_469/Y INVX1_LOC_359/A 0.01fF
C11500 INVX1_LOC_80/A INVX1_LOC_502/A 0.07fF
C11501 INVX1_LOC_298/Y INVX1_LOC_300/Y 0.39fF
C11502 INVX1_LOC_551/Y INVX1_LOC_74/Y 0.01fF
C11503 INVX1_LOC_160/Y INVX1_LOC_270/Y 0.01fF
C11504 INVX1_LOC_496/A NAND2X1_LOC_646/A 0.03fF
C11505 INVX1_LOC_361/A INVX1_LOC_48/Y 0.03fF
C11506 INVX1_LOC_32/Y INVX1_LOC_69/Y 5.81fF
C11507 INVX1_LOC_551/A NAND2X1_LOC_615/B 0.00fF
C11508 INVX1_LOC_674/A NAND2X1_LOC_334/A 0.07fF
C11509 NAND2X1_LOC_388/A INVX1_LOC_317/A 0.00fF
C11510 INVX1_LOC_387/Y INVX1_LOC_6/Y 0.03fF
C11511 INVX1_LOC_371/A INVX1_LOC_9/Y 0.07fF
C11512 INVX1_LOC_513/A INVX1_LOC_501/A 0.00fF
C11513 INVX1_LOC_119/Y INVX1_LOC_98/Y 0.03fF
C11514 INVX1_LOC_282/A INVX1_LOC_664/A 0.00fF
C11515 INVX1_LOC_360/Y INVX1_LOC_114/A 0.01fF
C11516 INVX1_LOC_301/Y INPUT_1 0.03fF
C11517 INVX1_LOC_358/A INVX1_LOC_479/A 0.03fF
C11518 INVX1_LOC_49/Y INVX1_LOC_6/Y 0.23fF
C11519 INVX1_LOC_11/Y INVX1_LOC_502/A 0.08fF
C11520 INVX1_LOC_204/Y NAND2X1_LOC_824/a_36_24# 0.01fF
C11521 INVX1_LOC_382/A INVX1_LOC_9/Y 0.02fF
C11522 INVX1_LOC_557/Y INVX1_LOC_46/Y 0.05fF
C11523 NAND2X1_LOC_136/Y INVX1_LOC_50/Y 0.22fF
C11524 INVX1_LOC_17/Y INVX1_LOC_505/Y 0.02fF
C11525 INVX1_LOC_298/Y INVX1_LOC_660/A 0.09fF
C11526 INVX1_LOC_63/Y INVX1_LOC_496/A 0.09fF
C11527 INVX1_LOC_153/A INVX1_LOC_90/Y 0.02fF
C11528 INVX1_LOC_531/Y INVX1_LOC_50/Y 0.07fF
C11529 INVX1_LOC_159/A INVX1_LOC_75/Y 0.02fF
C11530 INVX1_LOC_41/Y INPUT_1 0.22fF
C11531 INVX1_LOC_21/Y INVX1_LOC_270/Y 0.02fF
C11532 NAND2X1_LOC_686/B INVX1_LOC_245/A 0.02fF
C11533 NAND2X1_LOC_178/a_36_24# NAND2X1_LOC_274/B 0.00fF
C11534 INVX1_LOC_75/Y NAND2X1_LOC_615/B 0.02fF
C11535 INVX1_LOC_569/Y INVX1_LOC_662/A 0.03fF
C11536 INVX1_LOC_6/Y INVX1_LOC_210/A 0.01fF
C11537 INVX1_LOC_21/Y INVX1_LOC_92/A 0.03fF
C11538 NAND2X1_LOC_346/B INVX1_LOC_280/A 0.16fF
C11539 NAND2X1_LOC_666/a_36_24# INVX1_LOC_636/A 0.01fF
C11540 INVX1_LOC_75/Y INVX1_LOC_66/A 0.16fF
C11541 NAND2X1_LOC_373/a_36_24# NAND2X1_LOC_373/Y 0.02fF
C11542 NAND2X1_LOC_267/A INVX1_LOC_270/Y 0.02fF
C11543 NAND2X1_LOC_267/A INVX1_LOC_92/A 0.20fF
C11544 INVX1_LOC_555/A INVX1_LOC_92/A 0.11fF
C11545 INVX1_LOC_414/Y VDD 0.21fF
C11546 INVX1_LOC_486/Y INVX1_LOC_297/Y 0.16fF
C11547 NAND2X1_LOC_116/a_36_24# INVX1_LOC_109/A 0.02fF
C11548 INVX1_LOC_390/Y INVX1_LOC_410/Y 0.10fF
C11549 INVX1_LOC_20/Y NAND2X1_LOC_790/B 0.07fF
C11550 NAND2X1_LOC_274/B INVX1_LOC_666/Y 0.00fF
C11551 INVX1_LOC_100/Y NAND2X1_LOC_410/Y 0.05fF
C11552 INVX1_LOC_150/A NAND2X1_LOC_685/B 0.10fF
C11553 NAND2X1_LOC_161/a_36_24# INVX1_LOC_586/A 0.01fF
C11554 INVX1_LOC_62/Y INVX1_LOC_441/A 0.00fF
C11555 INVX1_LOC_20/Y NAND2X1_LOC_385/a_36_24# 0.00fF
C11556 INVX1_LOC_62/Y INVX1_LOC_645/Y 0.01fF
C11557 NAND2X1_LOC_764/Y INVX1_LOC_366/A 0.01fF
C11558 INVX1_LOC_266/A NAND2X1_LOC_374/a_36_24# 0.00fF
C11559 INVX1_LOC_549/A NAND2X1_LOC_707/A 0.10fF
C11560 INVX1_LOC_177/Y INVX1_LOC_65/Y 0.02fF
C11561 INVX1_LOC_139/A INVX1_LOC_586/A 0.00fF
C11562 NAND2X1_LOC_322/Y INVX1_LOC_134/Y 0.02fF
C11563 INVX1_LOC_20/Y INVX1_LOC_122/Y 0.01fF
C11564 INVX1_LOC_424/A NAND2X1_LOC_517/Y 0.01fF
C11565 INVX1_LOC_647/Y NAND2X1_LOC_843/B 0.01fF
C11566 INVX1_LOC_542/A INVX1_LOC_45/Y 0.03fF
C11567 INVX1_LOC_140/Y INVX1_LOC_76/Y 0.00fF
C11568 INVX1_LOC_618/Y INVX1_LOC_624/A 0.00fF
C11569 INVX1_LOC_105/Y INVX1_LOC_109/Y 0.01fF
C11570 INVX1_LOC_74/Y INVX1_LOC_634/Y 0.07fF
C11571 NAND2X1_LOC_790/B INVX1_LOC_197/Y 0.07fF
C11572 NAND2X1_LOC_744/a_36_24# INVX1_LOC_53/Y 0.00fF
C11573 INVX1_LOC_617/Y INVX1_LOC_253/A 0.02fF
C11574 INVX1_LOC_224/Y INVX1_LOC_12/Y 0.07fF
C11575 INVX1_LOC_412/Y NAND2X1_LOC_603/Y 0.01fF
C11576 INPUT_0 INVX1_LOC_174/A 0.20fF
C11577 NAND2X1_LOC_542/a_36_24# INVX1_LOC_410/Y 0.00fF
C11578 NAND2X1_LOC_498/Y INVX1_LOC_596/A 0.07fF
C11579 NAND2X1_LOC_764/Y INVX1_LOC_597/A 0.13fF
C11580 INVX1_LOC_20/Y NAND2X1_LOC_491/a_36_24# 0.00fF
C11581 NAND2X1_LOC_756/Y NAND2X1_LOC_101/a_36_24# 0.01fF
C11582 VDD INVX1_LOC_8/Y 0.26fF
C11583 NAND2X1_LOC_475/A INVX1_LOC_98/Y 0.10fF
C11584 VDD INVX1_LOC_303/Y 0.21fF
C11585 NAND2X1_LOC_586/a_36_24# INVX1_LOC_638/A 0.00fF
C11586 INVX1_LOC_578/A INVX1_LOC_12/Y 0.13fF
C11587 INPUT_0 INVX1_LOC_288/Y 0.10fF
C11588 VDD INVX1_LOC_514/A -0.00fF
C11589 INVX1_LOC_434/A INVX1_LOC_218/Y 0.11fF
C11590 INVX1_LOC_325/Y INPUT_2 0.02fF
C11591 VDD INVX1_LOC_587/Y 0.26fF
C11592 INVX1_LOC_20/Y NAND2X1_LOC_13/a_36_24# 0.00fF
C11593 INVX1_LOC_233/Y INVX1_LOC_134/Y 0.16fF
C11594 INVX1_LOC_563/Y INVX1_LOC_35/Y 0.01fF
C11595 INVX1_LOC_76/Y INVX1_LOC_486/Y 0.04fF
C11596 INVX1_LOC_435/Y INVX1_LOC_99/Y 0.11fF
C11597 VDD INVX1_LOC_539/Y 0.21fF
C11598 NAND2X1_LOC_507/a_36_24# INVX1_LOC_600/A 0.01fF
C11599 NAND2X1_LOC_704/B NAND2X1_LOC_307/A 0.00fF
C11600 INVX1_LOC_254/Y INVX1_LOC_206/Y 0.15fF
C11601 INVX1_LOC_286/Y INVX1_LOC_80/A 0.02fF
C11602 INVX1_LOC_296/Y INVX1_LOC_321/A 0.01fF
C11603 INVX1_LOC_51/Y INVX1_LOC_155/Y 0.03fF
C11604 INVX1_LOC_428/A NAND2X1_LOC_485/a_36_24# 0.00fF
C11605 NAND2X1_LOC_750/Y INVX1_LOC_87/A 0.01fF
C11606 VDD INVX1_LOC_306/Y 0.26fF
C11607 INVX1_LOC_554/A NAND2X1_LOC_846/B 0.01fF
C11608 NAND2X1_LOC_537/B INVX1_LOC_32/Y 0.01fF
C11609 INVX1_LOC_395/A INVX1_LOC_315/A 0.20fF
C11610 INVX1_LOC_386/A INVX1_LOC_220/A 0.02fF
C11611 INVX1_LOC_29/Y INVX1_LOC_333/A 0.04fF
C11612 NAND2X1_LOC_764/Y INVX1_LOC_6/Y 0.02fF
C11613 INVX1_LOC_206/Y INVX1_LOC_592/Y 0.02fF
C11614 NAND2X1_LOC_636/B INVX1_LOC_633/Y 0.06fF
C11615 NAND2X1_LOC_669/Y INVX1_LOC_53/Y 0.02fF
C11616 INVX1_LOC_449/A INVX1_LOC_53/Y 0.07fF
C11617 INVX1_LOC_85/Y INVX1_LOC_198/A 0.12fF
C11618 INVX1_LOC_224/Y INVX1_LOC_188/A 0.06fF
C11619 INVX1_LOC_680/Y INVX1_LOC_367/A 0.02fF
C11620 INVX1_LOC_413/Y INVX1_LOC_362/A 0.05fF
C11621 VDD INVX1_LOC_285/Y 0.21fF
C11622 INVX1_LOC_20/Y INVX1_LOC_556/Y 0.03fF
C11623 NAND2X1_LOC_460/A INVX1_LOC_310/Y 0.16fF
C11624 INVX1_LOC_211/Y INVX1_LOC_381/A 0.02fF
C11625 VDD INVX1_LOC_534/Y 0.35fF
C11626 INVX1_LOC_174/Y INVX1_LOC_86/Y 0.02fF
C11627 VDD INVX1_LOC_9/Y 1.47fF
C11628 INVX1_LOC_68/Y NAND2X1_LOC_165/Y 0.02fF
C11629 INVX1_LOC_410/Y NAND2X1_LOC_542/A 0.25fF
C11630 VDD NAND2X1_LOC_800/B 0.01fF
C11631 INVX1_LOC_531/Y INVX1_LOC_275/A 0.12fF
C11632 INVX1_LOC_608/Y INVX1_LOC_80/A 0.03fF
C11633 INVX1_LOC_45/Y NAND2X1_LOC_707/B 0.01fF
C11634 INVX1_LOC_586/A INVX1_LOC_32/Y 0.35fF
C11635 INVX1_LOC_47/A INVX1_LOC_600/A 0.01fF
C11636 INVX1_LOC_17/Y NAND2X1_LOC_528/a_36_24# 0.00fF
C11637 INVX1_LOC_117/Y NAND2X1_LOC_613/Y 0.03fF
C11638 INVX1_LOC_17/Y INVX1_LOC_80/A 1.02fF
C11639 INVX1_LOC_317/Y NAND2X1_LOC_388/A 0.00fF
C11640 INVX1_LOC_136/Y INVX1_LOC_98/Y 0.03fF
C11641 NAND2X1_LOC_318/B INVX1_LOC_99/Y 0.04fF
C11642 INVX1_LOC_45/Y INVX1_LOC_204/Y 0.00fF
C11643 INVX1_LOC_381/A INVX1_LOC_46/Y 0.07fF
C11644 INVX1_LOC_228/Y INVX1_LOC_9/Y -0.03fF
C11645 VDD INVX1_LOC_166/Y 0.39fF
C11646 INVX1_LOC_504/A INVX1_LOC_99/Y 0.07fF
C11647 INVX1_LOC_117/Y INVX1_LOC_337/Y 0.06fF
C11648 INVX1_LOC_375/A INVX1_LOC_376/Y 0.17fF
C11649 INVX1_LOC_76/Y INVX1_LOC_6/Y 0.00fF
C11650 INVX1_LOC_379/A NAND2X1_LOC_416/Y 0.01fF
C11651 INVX1_LOC_266/Y INVX1_LOC_199/Y 0.02fF
C11652 INVX1_LOC_546/A INVX1_LOC_376/Y 0.01fF
C11653 INVX1_LOC_7/Y NAND2X1_LOC_378/Y 0.03fF
C11654 INVX1_LOC_53/Y INVX1_LOC_186/Y 0.07fF
C11655 INVX1_LOC_31/A INVX1_LOC_204/Y 0.05fF
C11656 VDD INVX1_LOC_62/Y 1.44fF
C11657 INVX1_LOC_248/Y INVX1_LOC_252/Y 0.01fF
C11658 INVX1_LOC_117/Y INVX1_LOC_633/Y 0.07fF
C11659 NAND2X1_LOC_266/a_36_24# INVX1_LOC_178/A 0.01fF
C11660 INVX1_LOC_291/A NAND2X1_LOC_753/Y 0.02fF
C11661 NAND2X1_LOC_331/Y INVX1_LOC_259/Y 0.00fF
C11662 INVX1_LOC_320/A INVX1_LOC_46/Y 0.02fF
C11663 INVX1_LOC_53/Y NAND2X1_LOC_146/a_36_24# 0.00fF
C11664 INVX1_LOC_608/Y INVX1_LOC_11/Y 0.02fF
C11665 INVX1_LOC_541/Y INVX1_LOC_496/Y 0.01fF
C11666 VDD INVX1_LOC_13/Y 0.38fF
C11667 INVX1_LOC_304/Y INVX1_LOC_145/Y 0.05fF
C11668 INVX1_LOC_608/A NAND2X1_LOC_496/Y 0.06fF
C11669 INVX1_LOC_11/Y INVX1_LOC_17/Y 5.26fF
C11670 NAND2X1_LOC_697/Y NAND2X1_LOC_708/A 0.10fF
C11671 INVX1_LOC_371/Y INVX1_LOC_670/A 0.20fF
C11672 INVX1_LOC_21/Y INPUT_1 0.12fF
C11673 VDD INVX1_LOC_529/Y 0.26fF
C11674 NAND2X1_LOC_755/B NAND2X1_LOC_720/A 0.31fF
C11675 INVX1_LOC_206/Y NAND2X1_LOC_528/Y 0.02fF
C11676 NAND2X1_LOC_596/Y INVX1_LOC_62/Y 0.07fF
C11677 NAND2X1_LOC_829/Y INVX1_LOC_463/Y 0.01fF
C11678 INVX1_LOC_131/A NAND2X1_LOC_342/A 0.21fF
C11679 INVX1_LOC_45/Y INVX1_LOC_114/A 0.07fF
C11680 INVX1_LOC_418/A INVX1_LOC_100/Y 0.14fF
C11681 INVX1_LOC_206/Y INVX1_LOC_479/A 0.26fF
C11682 INVX1_LOC_93/Y INVX1_LOC_186/A 0.01fF
C11683 INVX1_LOC_558/A INVX1_LOC_100/Y 0.09fF
C11684 INVX1_LOC_255/Y NAND2X1_LOC_123/B 0.07fF
C11685 NAND2X1_LOC_324/B INVX1_LOC_69/Y 0.13fF
C11686 INPUT_5 INVX1_LOC_60/Y 0.01fF
C11687 INVX1_LOC_435/A INVX1_LOC_54/Y 0.18fF
C11688 INVX1_LOC_678/A INVX1_LOC_673/Y 0.09fF
C11689 INVX1_LOC_288/Y INVX1_LOC_498/A 0.15fF
C11690 INVX1_LOC_562/Y INVX1_LOC_26/Y 0.01fF
C11691 INVX1_LOC_449/A NAND2X1_LOC_274/Y 0.01fF
C11692 INVX1_LOC_93/Y INVX1_LOC_176/A 0.21fF
C11693 INVX1_LOC_20/Y NAND2X1_LOC_420/Y -0.00fF
C11694 INVX1_LOC_581/Y NAND2X1_LOC_679/B 0.05fF
C11695 NAND2X1_LOC_318/B INVX1_LOC_47/Y 0.02fF
C11696 INVX1_LOC_386/Y INVX1_LOC_6/Y 0.03fF
C11697 INVX1_LOC_58/Y NAND2X1_LOC_496/Y 0.19fF
C11698 INVX1_LOC_134/A INVX1_LOC_41/Y 0.01fF
C11699 INVX1_LOC_173/Y INVX1_LOC_35/Y 0.00fF
C11700 INVX1_LOC_298/A NAND2X1_LOC_826/a_36_24# 0.00fF
C11701 INVX1_LOC_12/Y INVX1_LOC_120/Y 0.03fF
C11702 INVX1_LOC_32/Y NAND2X1_LOC_74/a_36_24# 0.01fF
C11703 INVX1_LOC_614/A INVX1_LOC_9/Y 0.15fF
C11704 NAND2X1_LOC_820/Y INVX1_LOC_655/A 0.04fF
C11705 INVX1_LOC_679/Y INVX1_LOC_107/Y 0.01fF
C11706 INVX1_LOC_551/Y INVX1_LOC_79/A 0.07fF
C11707 INVX1_LOC_348/A INVX1_LOC_114/A 0.01fF
C11708 INVX1_LOC_53/Y INVX1_LOC_328/Y 0.03fF
C11709 INVX1_LOC_366/A INVX1_LOC_184/Y 0.03fF
C11710 INVX1_LOC_93/Y INVX1_LOC_349/A 0.02fF
C11711 INVX1_LOC_270/A INVX1_LOC_100/Y 0.03fF
C11712 NAND2X1_LOC_121/Y INVX1_LOC_632/A 0.02fF
C11713 INVX1_LOC_42/A INVX1_LOC_9/Y 0.01fF
C11714 NAND2X1_LOC_294/Y INVX1_LOC_381/Y 0.03fF
C11715 NAND2X1_LOC_706/B INVX1_LOC_608/A 0.21fF
C11716 INVX1_LOC_69/Y NAND2X1_LOC_226/Y 0.18fF
C11717 INVX1_LOC_235/Y NAND2X1_LOC_269/B 0.01fF
C11718 INVX1_LOC_53/Y INVX1_LOC_518/A 0.04fF
C11719 NAND2X1_LOC_137/A INPUT_1 0.03fF
C11720 INVX1_LOC_17/Y NAND2X1_LOC_359/a_36_24# 0.00fF
C11721 INVX1_LOC_11/Y NAND2X1_LOC_307/B 0.02fF
C11722 INVX1_LOC_659/A INVX1_LOC_656/Y 0.03fF
C11723 INVX1_LOC_555/A INPUT_1 0.02fF
C11724 INVX1_LOC_183/A INVX1_LOC_145/Y 0.02fF
C11725 NAND2X1_LOC_333/a_36_24# INVX1_LOC_50/Y 0.00fF
C11726 INVX1_LOC_479/A INVX1_LOC_242/A 0.03fF
C11727 NAND2X1_LOC_686/A INVX1_LOC_537/A 0.04fF
C11728 INVX1_LOC_270/A INVX1_LOC_74/Y 0.03fF
C11729 INVX1_LOC_124/A INVX1_LOC_669/Y 0.14fF
C11730 INVX1_LOC_108/A INVX1_LOC_6/Y 0.01fF
C11731 INVX1_LOC_326/A INVX1_LOC_326/Y 0.01fF
C11732 INVX1_LOC_32/Y INVX1_LOC_157/Y 0.01fF
C11733 INVX1_LOC_614/A INVX1_LOC_62/Y 0.02fF
C11734 INVX1_LOC_449/A NAND2X1_LOC_844/a_36_24# 0.00fF
C11735 INVX1_LOC_48/Y INVX1_LOC_480/A 0.01fF
C11736 INVX1_LOC_400/A INVX1_LOC_399/Y 0.03fF
C11737 INVX1_LOC_686/A INVX1_LOC_479/A 0.07fF
C11738 INVX1_LOC_74/Y INVX1_LOC_333/A 0.14fF
C11739 INVX1_LOC_555/A NAND2X1_LOC_277/a_36_24# 0.01fF
C11740 INVX1_LOC_504/A INVX1_LOC_119/Y 0.08fF
C11741 INVX1_LOC_675/A INVX1_LOC_354/Y 0.05fF
C11742 INVX1_LOC_502/A INVX1_LOC_367/Y 0.07fF
C11743 NAND2X1_LOC_27/Y INVX1_LOC_223/Y 0.02fF
C11744 INVX1_LOC_93/Y INVX1_LOC_170/Y 0.00fF
C11745 INVX1_LOC_301/Y INVX1_LOC_50/Y 0.03fF
C11746 GATE_662 INVX1_LOC_199/Y 0.00fF
C11747 INVX1_LOC_277/Y INVX1_LOC_283/A 0.16fF
C11748 INVX1_LOC_103/Y INVX1_LOC_9/Y 0.06fF
C11749 INVX1_LOC_62/Y INVX1_LOC_116/A 0.01fF
C11750 INVX1_LOC_93/Y INVX1_LOC_124/A 0.01fF
C11751 INVX1_LOC_344/Y INVX1_LOC_588/A 0.06fF
C11752 INVX1_LOC_599/Y INVX1_LOC_598/Y 0.00fF
C11753 NAND2X1_LOC_545/A INVX1_LOC_159/Y 0.05fF
C11754 NAND2X1_LOC_679/A INVX1_LOC_463/Y 0.04fF
C11755 INVX1_LOC_513/A INVX1_LOC_461/Y 0.01fF
C11756 INVX1_LOC_167/A INVX1_LOC_79/A 0.01fF
C11757 INVX1_LOC_199/Y NAND2X1_LOC_846/B 0.01fF
C11758 NAND2X1_LOC_666/a_36_24# INVX1_LOC_74/Y 0.01fF
C11759 INVX1_LOC_75/Y INVX1_LOC_116/Y 0.02fF
C11760 INVX1_LOC_133/Y INVX1_LOC_185/A 0.01fF
C11761 INVX1_LOC_298/A NAND2X1_LOC_836/a_36_24# 0.00fF
C11762 NAND2X1_LOC_106/Y INVX1_LOC_26/Y 0.03fF
C11763 INVX1_LOC_41/Y INVX1_LOC_50/Y 3.15fF
C11764 INVX1_LOC_100/Y INVX1_LOC_46/Y 0.32fF
C11765 INVX1_LOC_99/Y INVX1_LOC_346/Y 0.07fF
C11766 NAND2X1_LOC_513/A INVX1_LOC_613/A 0.08fF
C11767 NAND2X1_LOC_847/A NAND2X1_LOC_817/a_36_24# 0.00fF
C11768 INVX1_LOC_15/Y INVX1_LOC_338/Y 0.04fF
C11769 INVX1_LOC_159/Y INVX1_LOC_666/Y 0.46fF
C11770 INVX1_LOC_103/Y INVX1_LOC_62/Y 0.03fF
C11771 INVX1_LOC_587/Y INVX1_LOC_635/Y 0.02fF
C11772 INVX1_LOC_79/A NAND2X1_LOC_759/Y 0.01fF
C11773 NAND2X1_LOC_843/B NAND2X1_LOC_342/A 0.03fF
C11774 NAND2X1_LOC_287/a_36_24# INVX1_LOC_66/A 0.00fF
C11775 INVX1_LOC_152/Y INVX1_LOC_150/A 0.20fF
C11776 INVX1_LOC_469/Y INVX1_LOC_634/Y 0.01fF
C11777 INVX1_LOC_353/A INVX1_LOC_90/Y 0.03fF
C11778 NAND2X1_LOC_334/A INVX1_LOC_479/A 0.07fF
C11779 INVX1_LOC_93/Y INVX1_LOC_611/A 0.01fF
C11780 INVX1_LOC_121/Y INVX1_LOC_553/Y 0.01fF
C11781 INVX1_LOC_192/Y INVX1_LOC_224/Y 0.03fF
C11782 INVX1_LOC_434/A INVX1_LOC_429/Y 0.11fF
C11783 INVX1_LOC_3/Y INVX1_LOC_33/A 0.32fF
C11784 INPUT_6 NAND2X1_LOC_25/a_36_24# 0.00fF
C11785 INVX1_LOC_329/Y INVX1_LOC_26/Y 0.01fF
C11786 INVX1_LOC_373/Y INVX1_LOC_588/A 0.98fF
C11787 VDD INVX1_LOC_580/Y 0.35fF
C11788 INVX1_LOC_49/Y INVX1_LOC_636/A 0.07fF
C11789 NAND2X1_LOC_46/a_36_24# INVX1_LOC_578/A 0.00fF
C11790 NAND2X1_LOC_770/A NAND2X1_LOC_791/B 0.02fF
C11791 NAND2X1_LOC_770/A INVX1_LOC_272/Y 0.00fF
C11792 INVX1_LOC_62/Y INVX1_LOC_635/Y 0.03fF
C11793 INVX1_LOC_119/Y INVX1_LOC_346/Y 0.01fF
C11794 INVX1_LOC_375/A INVX1_LOC_253/A 0.03fF
C11795 NAND2X1_LOC_750/Y INVX1_LOC_191/A 0.00fF
C11796 INVX1_LOC_578/A NAND2X1_LOC_150/a_36_24# 0.00fF
C11797 NAND2X1_LOC_475/A INVX1_LOC_596/A 0.02fF
C11798 INVX1_LOC_206/Y INVX1_LOC_372/Y 0.03fF
C11799 VDD INVX1_LOC_344/A -0.00fF
C11800 NAND2X1_LOC_317/A INVX1_LOC_53/Y 0.03fF
C11801 NAND2X1_LOC_45/Y INVX1_LOC_530/A 0.04fF
C11802 NAND2X1_LOC_754/a_36_24# INVX1_LOC_98/Y 0.00fF
C11803 NAND2X1_LOC_543/B INVX1_LOC_98/Y 0.10fF
C11804 INVX1_LOC_206/Y INVX1_LOC_12/Y 4.60fF
C11805 INPUT_0 INVX1_LOC_188/Y 0.03fF
C11806 VDD INVX1_LOC_42/Y 0.21fF
C11807 INVX1_LOC_436/Y VDD 0.16fF
C11808 INPUT_0 NAND2X1_LOC_411/Y 0.01fF
C11809 INVX1_LOC_53/Y INVX1_LOC_521/Y 0.30fF
C11810 INVX1_LOC_359/Y INVX1_LOC_638/A 0.03fF
C11811 VDD NAND2X1_LOC_190/A 0.08fF
C11812 NAND2X1_LOC_79/a_36_24# INVX1_LOC_366/A 0.01fF
C11813 INPUT_3 INVX1_LOC_378/A 0.01fF
C11814 VDD INVX1_LOC_593/Y 0.54fF
C11815 VDD INVX1_LOC_87/A 0.31fF
C11816 VDD INVX1_LOC_641/Y 0.22fF
C11817 INVX1_LOC_413/Y INVX1_LOC_145/Y 0.07fF
C11818 NAND2X1_LOC_249/Y NAND2X1_LOC_106/Y 0.03fF
C11819 INVX1_LOC_554/A INVX1_LOC_199/Y 0.03fF
C11820 INVX1_LOC_130/Y INVX1_LOC_586/A 0.01fF
C11821 NAND2X1_LOC_788/A NAND2X1_LOC_469/a_36_24# 0.00fF
C11822 INVX1_LOC_578/A INVX1_LOC_159/A 0.01fF
C11823 INVX1_LOC_372/Y INVX1_LOC_686/A 0.00fF
C11824 VDD INVX1_LOC_631/Y 0.21fF
C11825 INVX1_LOC_366/A INVX1_LOC_7/Y 0.01fF
C11826 NAND2X1_LOC_193/a_36_24# INVX1_LOC_6/Y 0.00fF
C11827 INVX1_LOC_68/Y NAND2X1_LOC_165/a_36_24# 0.00fF
C11828 INVX1_LOC_417/Y INVX1_LOC_551/Y 0.25fF
C11829 INVX1_LOC_662/Y NAND2X1_LOC_142/Y 0.32fF
C11830 INVX1_LOC_540/Y NAND2X1_LOC_689/B 0.06fF
C11831 INVX1_LOC_193/Y INVX1_LOC_93/Y 0.01fF
C11832 VDD INVX1_LOC_624/Y 0.27fF
C11833 INVX1_LOC_12/Y INVX1_LOC_686/A 0.02fF
C11834 INVX1_LOC_680/Y INVX1_LOC_683/Y 0.97fF
C11835 INVX1_LOC_590/Y NAND2X1_LOC_387/Y 0.03fF
C11836 INVX1_LOC_224/Y INVX1_LOC_296/A 0.00fF
C11837 INVX1_LOC_551/Y INVX1_LOC_59/Y 0.01fF
C11838 INVX1_LOC_315/Y INVX1_LOC_50/Y 0.03fF
C11839 INVX1_LOC_84/A NAND2X1_LOC_67/Y 0.03fF
C11840 INVX1_LOC_386/Y NAND2X1_LOC_517/Y 0.03fF
C11841 INVX1_LOC_578/A INVX1_LOC_66/A 0.07fF
C11842 INVX1_LOC_551/Y INVX1_LOC_48/Y 0.03fF
C11843 INVX1_LOC_545/A INVX1_LOC_80/A 0.00fF
C11844 INVX1_LOC_373/A INVX1_LOC_494/Y 0.01fF
C11845 INVX1_LOC_193/Y INVX1_LOC_390/A 0.00fF
C11846 INVX1_LOC_561/Y NAND2X1_LOC_121/Y 0.00fF
C11847 INVX1_LOC_288/Y INVX1_LOC_677/A 0.01fF
C11848 INVX1_LOC_300/A INVX1_LOC_565/A 0.06fF
C11849 INVX1_LOC_540/Y INVX1_LOC_245/A 0.02fF
C11850 INPUT_0 NAND2X1_LOC_845/B 0.01fF
C11851 INVX1_LOC_595/Y NAND2X1_LOC_460/A 0.01fF
C11852 INVX1_LOC_417/A INVX1_LOC_35/Y 0.01fF
C11853 INVX1_LOC_54/Y INVX1_LOC_367/A 0.10fF
C11854 INVX1_LOC_625/A INVX1_LOC_99/Y 0.02fF
C11855 INVX1_LOC_362/Y INVX1_LOC_420/A 0.02fF
C11856 INVX1_LOC_53/Y INVX1_LOC_172/A 0.02fF
C11857 INVX1_LOC_361/Y INVX1_LOC_545/Y 0.03fF
C11858 NAND2X1_LOC_516/B INVX1_LOC_89/Y 0.00fF
C11859 INVX1_LOC_340/A INVX1_LOC_55/Y 0.01fF
C11860 INVX1_LOC_294/Y INVX1_LOC_32/Y 0.01fF
C11861 INVX1_LOC_206/Y INVX1_LOC_680/A 0.01fF
C11862 INVX1_LOC_17/Y INVX1_LOC_367/Y 0.16fF
C11863 NAND2X1_LOC_498/B NAND2X1_LOC_192/A 0.03fF
C11864 INVX1_LOC_271/A INVX1_LOC_245/A 0.01fF
C11865 INVX1_LOC_393/Y INVX1_LOC_502/A 0.01fF
C11866 INVX1_LOC_68/Y INVX1_LOC_351/A 0.05fF
C11867 INVX1_LOC_21/Y INVX1_LOC_50/Y 0.10fF
C11868 INVX1_LOC_381/A INVX1_LOC_49/Y 0.00fF
C11869 INVX1_LOC_415/Y INVX1_LOC_386/Y 0.15fF
C11870 INVX1_LOC_214/Y NAND2X1_LOC_106/B 0.02fF
C11871 NAND2X1_LOC_192/A INVX1_LOC_76/Y 0.00fF
C11872 INVX1_LOC_493/A INVX1_LOC_491/Y 0.02fF
C11873 INVX1_LOC_243/A INVX1_LOC_46/Y 0.01fF
C11874 INVX1_LOC_58/Y INVX1_LOC_337/Y 0.08fF
C11875 INVX1_LOC_58/Y INVX1_LOC_495/A 0.06fF
C11876 NAND2X1_LOC_299/Y INVX1_LOC_69/Y 0.07fF
C11877 INVX1_LOC_530/Y INVX1_LOC_100/Y 0.07fF
C11878 INVX1_LOC_400/A INVX1_LOC_54/Y 0.07fF
C11879 INVX1_LOC_68/Y INVX1_LOC_90/Y 0.03fF
C11880 INVX1_LOC_402/Y INVX1_LOC_89/Y 0.00fF
C11881 INVX1_LOC_54/Y INVX1_LOC_392/A 0.03fF
C11882 INVX1_LOC_441/Y INVX1_LOC_41/Y 0.02fF
C11883 INVX1_LOC_47/Y INVX1_LOC_530/A 0.01fF
C11884 INVX1_LOC_58/Y INVX1_LOC_633/Y 0.03fF
C11885 INVX1_LOC_386/Y NAND2X1_LOC_294/Y 0.03fF
C11886 GATE_865 INVX1_LOC_263/Y 0.01fF
C11887 INVX1_LOC_31/Y INVX1_LOC_176/A 0.17fF
C11888 INVX1_LOC_684/A INVX1_LOC_641/Y 0.01fF
C11889 INVX1_LOC_419/Y INVX1_LOC_361/Y 0.07fF
C11890 INVX1_LOC_6/Y INVX1_LOC_7/Y 0.22fF
C11891 INVX1_LOC_53/Y NAND2X1_LOC_846/B 0.05fF
C11892 NAND2X1_LOC_318/A INVX1_LOC_100/Y 0.18fF
C11893 INVX1_LOC_525/Y INVX1_LOC_35/Y 0.03fF
C11894 INVX1_LOC_468/Y INVX1_LOC_66/A 0.04fF
C11895 INVX1_LOC_11/Y INVX1_LOC_230/Y 0.07fF
C11896 INVX1_LOC_435/A INVX1_LOC_89/Y 0.94fF
C11897 INVX1_LOC_288/A NAND2X1_LOC_434/a_36_24# 0.00fF
C11898 INPUT_3 INVX1_LOC_422/A 0.03fF
C11899 INVX1_LOC_270/A INVX1_LOC_79/A 0.01fF
C11900 INVX1_LOC_451/A NAND2X1_LOC_531/Y 0.05fF
C11901 NAND2X1_LOC_748/a_36_24# INVX1_LOC_198/A 0.00fF
C11902 INVX1_LOC_99/Y NAND2X1_LOC_52/Y 0.01fF
C11903 INVX1_LOC_54/Y INVX1_LOC_93/Y 0.58fF
C11904 INVX1_LOC_166/A INVX1_LOC_117/Y 0.03fF
C11905 INVX1_LOC_530/Y INVX1_LOC_483/Y 0.01fF
C11906 INVX1_LOC_351/A INVX1_LOC_600/A 0.02fF
C11907 INVX1_LOC_298/A NAND2X1_LOC_387/Y 0.01fF
C11908 NAND2X1_LOC_318/A INVX1_LOC_74/Y 0.06fF
C11909 NAND2X1_LOC_111/Y NAND2X1_LOC_112/a_36_24# 0.00fF
C11910 INVX1_LOC_560/A INVX1_LOC_92/A 0.07fF
C11911 INVX1_LOC_32/Y INVX1_LOC_6/Y 0.68fF
C11912 NAND2X1_LOC_415/B INVX1_LOC_245/A 0.32fF
C11913 INVX1_LOC_600/A INVX1_LOC_90/Y 0.01fF
C11914 INVX1_LOC_49/Y NAND2X1_LOC_720/A 0.02fF
C11915 INVX1_LOC_525/Y INVX1_LOC_620/A 0.18fF
C11916 NAND2X1_LOC_184/Y INVX1_LOC_69/Y 0.06fF
C11917 NAND2X1_LOC_770/B INVX1_LOC_63/Y 0.02fF
C11918 NAND2X1_LOC_755/B INVX1_LOC_79/A 0.03fF
C11919 INVX1_LOC_410/A INVX1_LOC_31/Y 0.00fF
C11920 INVX1_LOC_286/Y INVX1_LOC_91/Y 0.02fF
C11921 INVX1_LOC_100/Y INVX1_LOC_363/Y 0.01fF
C11922 INVX1_LOC_31/Y INVX1_LOC_420/A 0.00fF
C11923 INVX1_LOC_170/Y INVX1_LOC_31/Y 0.03fF
C11924 INVX1_LOC_304/Y INVX1_LOC_242/Y 0.02fF
C11925 INVX1_LOC_6/Y NAND2X1_LOC_815/a_36_24# 0.00fF
C11926 INVX1_LOC_202/Y INVX1_LOC_100/Y 0.10fF
C11927 INVX1_LOC_357/Y INVX1_LOC_463/Y 0.01fF
C11928 INVX1_LOC_513/A NAND2X1_LOC_436/a_36_24# 0.00fF
C11929 INVX1_LOC_47/Y NAND2X1_LOC_52/Y 0.01fF
C11930 INPUT_1 INVX1_LOC_26/Y 0.03fF
C11931 INVX1_LOC_377/A INVX1_LOC_666/Y 0.05fF
C11932 INVX1_LOC_115/A INVX1_LOC_74/Y 0.00fF
C11933 NAND2X1_LOC_827/Y INVX1_LOC_659/A 0.01fF
C11934 INVX1_LOC_360/Y INVX1_LOC_62/Y 0.07fF
C11935 INPUT_1 INVX1_LOC_128/Y 0.78fF
C11936 INVX1_LOC_117/Y NAND2X1_LOC_136/Y 0.10fF
C11937 GATE_865 INVX1_LOC_454/Y 0.00fF
C11938 INVX1_LOC_376/A INVX1_LOC_258/Y 0.02fF
C11939 INVX1_LOC_202/Y INVX1_LOC_74/Y 0.07fF
C11940 INVX1_LOC_79/A INVX1_LOC_46/Y 0.06fF
C11941 INVX1_LOC_47/Y NAND2X1_LOC_686/A 0.02fF
C11942 INVX1_LOC_369/A INVX1_LOC_485/A 0.01fF
C11943 NAND2X1_LOC_157/a_36_24# INVX1_LOC_145/A 0.00fF
C11944 INVX1_LOC_117/Y INVX1_LOC_531/Y 0.23fF
C11945 INVX1_LOC_26/Y INVX1_LOC_292/Y 0.09fF
C11946 INVX1_LOC_484/A INVX1_LOC_90/Y 0.00fF
C11947 INVX1_LOC_387/Y INVX1_LOC_100/Y 0.03fF
C11948 INVX1_LOC_17/Y INVX1_LOC_625/Y 0.00fF
C11949 NAND2X1_LOC_631/B INVX1_LOC_46/Y 0.02fF
C11950 INVX1_LOC_478/Y INVX1_LOC_211/A 0.01fF
C11951 NAND2X1_LOC_416/Y INVX1_LOC_488/Y 0.16fF
C11952 INVX1_LOC_47/Y INVX1_LOC_519/Y 0.01fF
C11953 INVX1_LOC_664/A INVX1_LOC_654/Y 0.03fF
C11954 INVX1_LOC_26/Y INVX1_LOC_284/Y 0.14fF
C11955 INVX1_LOC_451/A INVX1_LOC_443/A 0.19fF
C11956 NAND2X1_LOC_388/A INVX1_LOC_41/Y 0.00fF
C11957 NAND2X1_LOC_387/Y INVX1_LOC_211/A 0.07fF
C11958 INVX1_LOC_49/Y INVX1_LOC_100/Y 0.40fF
C11959 INVX1_LOC_255/A NAND2X1_LOC_441/a_36_24# 0.01fF
C11960 INVX1_LOC_399/A INVX1_LOC_26/Y 0.04fF
C11961 NAND2X1_LOC_409/Y NAND2X1_LOC_836/B 0.12fF
C11962 NAND2X1_LOC_686/A INVX1_LOC_119/Y 0.01fF
C11963 INVX1_LOC_270/Y INVX1_LOC_603/A 0.00fF
C11964 NAND2X1_LOC_174/a_36_24# INVX1_LOC_636/A 0.01fF
C11965 INVX1_LOC_69/Y INVX1_LOC_75/Y 0.03fF
C11966 NAND2X1_LOC_542/A INVX1_LOC_479/A 0.00fF
C11967 NAND2X1_LOC_475/A NAND2X1_LOC_76/B 0.04fF
C11968 INVX1_LOC_49/Y INVX1_LOC_74/Y 0.17fF
C11969 INVX1_LOC_519/Y INVX1_LOC_119/Y 0.00fF
C11970 INVX1_LOC_49/Y INVX1_LOC_483/Y 0.02fF
C11971 INVX1_LOC_603/A INVX1_LOC_92/A 0.02fF
C11972 VDD INVX1_LOC_404/Y 0.80fF
C11973 VDD NAND2X1_LOC_331/A 0.88fF
C11974 INVX1_LOC_479/A INVX1_LOC_376/Y 0.07fF
C11975 INVX1_LOC_381/A INVX1_LOC_297/Y 0.02fF
C11976 INVX1_LOC_424/A INVX1_LOC_450/A 0.18fF
C11977 NAND2X1_LOC_173/Y INVX1_LOC_638/A 0.20fF
C11978 NAND2X1_LOC_309/a_36_24# INVX1_LOC_92/A 0.00fF
C11979 VDD INVX1_LOC_271/Y 0.21fF
C11980 INVX1_LOC_69/Y NAND2X1_LOC_271/A 0.17fF
C11981 INVX1_LOC_193/Y INVX1_LOC_395/A 0.02fF
C11982 INVX1_LOC_79/A INVX1_LOC_75/A 0.00fF
C11983 INVX1_LOC_605/A INVX1_LOC_395/A 0.05fF
C11984 VDD INVX1_LOC_191/A -0.00fF
C11985 INVX1_LOC_85/Y INVX1_LOC_190/Y 0.41fF
C11986 NAND2X1_LOC_503/B INVX1_LOC_80/A 0.00fF
C11987 INVX1_LOC_554/A INVX1_LOC_53/Y 0.04fF
C11988 INVX1_LOC_578/A INVX1_LOC_442/A 0.31fF
C11989 INVX1_LOC_257/Y NAND2X1_LOC_180/B 0.01fF
C11990 INVX1_LOC_445/Y INVX1_LOC_220/Y 0.15fF
C11991 INVX1_LOC_21/Y INVX1_LOC_275/A 0.00fF
C11992 INVX1_LOC_3/Y INVX1_LOC_333/A 0.00fF
C11993 INVX1_LOC_293/Y NAND2X1_LOC_457/A 0.03fF
C11994 NAND2X1_LOC_249/Y INVX1_LOC_679/Y 0.16fF
C11995 INVX1_LOC_333/Y VDD 0.23fF
C11996 INVX1_LOC_21/Y INVX1_LOC_438/A 0.07fF
C11997 INVX1_LOC_616/A INVX1_LOC_366/A 0.06fF
C11998 INVX1_LOC_293/Y INVX1_LOC_547/Y 0.05fF
C11999 NAND2X1_LOC_788/A INVX1_LOC_468/Y 0.01fF
C12000 NAND2X1_LOC_24/Y NAND2X1_LOC_24/a_36_24# 0.03fF
C12001 INVX1_LOC_156/Y INVX1_LOC_577/Y 0.01fF
C12002 INVX1_LOC_301/A INVX1_LOC_304/Y 0.00fF
C12003 INVX1_LOC_625/A NAND2X1_LOC_475/A 0.09fF
C12004 VDD INVX1_LOC_407/Y -0.00fF
C12005 INVX1_LOC_21/Y INVX1_LOC_24/A 0.00fF
C12006 VDD INVX1_LOC_425/Y 0.21fF
C12007 INVX1_LOC_139/A INVX1_LOC_161/A 0.20fF
C12008 NAND2X1_LOC_551/a_36_24# INVX1_LOC_301/A 0.00fF
C12009 VDD INVX1_LOC_480/Y 0.39fF
C12010 INVX1_LOC_381/A INVX1_LOC_76/Y 0.08fF
C12011 NAND2X1_LOC_164/Y INVX1_LOC_99/Y 0.06fF
C12012 INVX1_LOC_412/A INVX1_LOC_99/A 0.39fF
C12013 INVX1_LOC_288/A INVX1_LOC_188/Y 0.03fF
C12014 INVX1_LOC_17/Y INVX1_LOC_393/Y 0.22fF
C12015 INVX1_LOC_80/A INVX1_LOC_273/A 0.07fF
C12016 NAND2X1_LOC_122/Y INVX1_LOC_579/Y 0.01fF
C12017 VDD INVX1_LOC_169/Y 0.21fF
C12018 INVX1_LOC_320/A INVX1_LOC_76/Y 0.02fF
C12019 INVX1_LOC_578/A INVX1_LOC_116/Y 0.57fF
C12020 INVX1_LOC_11/Y INVX1_LOC_127/A 0.13fF
C12021 INVX1_LOC_206/Y NAND2X1_LOC_615/B 0.47fF
C12022 INVX1_LOC_680/Y INVX1_LOC_51/Y 0.03fF
C12023 INVX1_LOC_65/Y INVX1_LOC_99/Y 0.06fF
C12024 NAND2X1_LOC_511/a_36_24# INVX1_LOC_14/A 0.00fF
C12025 NAND2X1_LOC_710/B INVX1_LOC_50/Y 0.04fF
C12026 INVX1_LOC_380/A INVX1_LOC_245/A 0.01fF
C12027 INVX1_LOC_293/Y INVX1_LOC_651/A 0.00fF
C12028 NAND2X1_LOC_705/a_36_24# INVX1_LOC_387/A 0.00fF
C12029 INVX1_LOC_414/A INVX1_LOC_46/Y 0.01fF
C12030 VDD INVX1_LOC_3/A -0.00fF
C12031 INVX1_LOC_51/Y INVX1_LOC_176/A 0.07fF
C12032 INVX1_LOC_118/Y INVX1_LOC_670/A 0.00fF
C12033 INVX1_LOC_54/Y INVX1_LOC_395/A 0.20fF
C12034 VDD INVX1_LOC_182/Y 0.21fF
C12035 INVX1_LOC_68/Y INVX1_LOC_98/Y 0.00fF
C12036 INVX1_LOC_457/Y INVX1_LOC_31/Y 0.01fF
C12037 INVX1_LOC_285/A INVX1_LOC_53/Y 0.02fF
C12038 INVX1_LOC_28/Y INVX1_LOC_27/A 0.03fF
C12039 INVX1_LOC_206/Y INVX1_LOC_66/A 0.02fF
C12040 INVX1_LOC_287/Y INVX1_LOC_59/Y 0.02fF
C12041 INVX1_LOC_54/Y INVX1_LOC_362/Y 0.03fF
C12042 INVX1_LOC_213/Y INVX1_LOC_651/Y 0.18fF
C12043 INVX1_LOC_57/Y INVX1_LOC_55/Y 1.02fF
C12044 INVX1_LOC_395/A INVX1_LOC_257/A 0.51fF
C12045 INVX1_LOC_617/Y INVX1_LOC_35/Y 0.39fF
C12046 INVX1_LOC_20/Y INVX1_LOC_304/Y 0.03fF
C12047 INVX1_LOC_438/Y GATE_479 0.10fF
C12048 INVX1_LOC_648/Y INVX1_LOC_66/A 0.04fF
C12049 INVX1_LOC_45/Y INVX1_LOC_539/Y 0.02fF
C12050 NAND2X1_LOC_299/Y NAND2X1_LOC_808/a_36_24# 0.01fF
C12051 INVX1_LOC_119/A INVX1_LOC_304/A 0.05fF
C12052 INVX1_LOC_605/Y INVX1_LOC_607/Y 0.06fF
C12053 INVX1_LOC_21/Y NAND2X1_LOC_513/A 0.00fF
C12054 INVX1_LOC_546/Y INVX1_LOC_89/Y 0.02fF
C12055 NAND2X1_LOC_184/Y INVX1_LOC_586/A 0.03fF
C12056 INVX1_LOC_26/Y INVX1_LOC_181/A 0.15fF
C12057 INVX1_LOC_455/A INVX1_LOC_55/Y 0.67fF
C12058 INVX1_LOC_176/Y INVX1_LOC_35/Y 0.00fF
C12059 INVX1_LOC_614/A INVX1_LOC_575/A 0.02fF
C12060 INVX1_LOC_287/Y INVX1_LOC_48/Y 0.01fF
C12061 INVX1_LOC_270/A INVX1_LOC_48/Y 0.03fF
C12062 VDD NAND2X1_LOC_833/B 0.03fF
C12063 INVX1_LOC_578/A INVX1_LOC_255/A 1.07fF
C12064 INVX1_LOC_286/Y NAND2X1_LOC_333/B 0.07fF
C12065 INVX1_LOC_607/A INVX1_LOC_69/Y 0.02fF
C12066 INVX1_LOC_65/Y INVX1_LOC_47/Y 0.03fF
C12067 INVX1_LOC_400/Y INVX1_LOC_63/Y 0.05fF
C12068 INVX1_LOC_616/A INVX1_LOC_6/Y 0.01fF
C12069 NAND2X1_LOC_789/B INVX1_LOC_26/Y 0.01fF
C12070 INVX1_LOC_11/Y NAND2X1_LOC_382/a_36_24# -0.00fF
C12071 INVX1_LOC_354/A INVX1_LOC_638/A 0.01fF
C12072 INVX1_LOC_66/A INVX1_LOC_242/A 0.06fF
C12073 INVX1_LOC_291/A INVX1_LOC_525/Y 0.11fF
C12074 INVX1_LOC_321/Y INVX1_LOC_681/A 0.04fF
C12075 NAND2X1_LOC_486/B INVX1_LOC_69/Y 0.03fF
C12076 INVX1_LOC_567/Y INVX1_LOC_556/Y 0.05fF
C12077 NAND2X1_LOC_755/B INVX1_LOC_59/Y 0.01fF
C12078 INPUT_4 NAND2X1_LOC_53/a_36_24# 0.00fF
C12079 INVX1_LOC_369/A INPUT_1 0.01fF
C12080 INVX1_LOC_424/Y INVX1_LOC_6/Y 0.03fF
C12081 INVX1_LOC_586/A INVX1_LOC_498/Y 0.46fF
C12082 INVX1_LOC_113/Y INVX1_LOC_675/A 0.07fF
C12083 INVX1_LOC_45/Y INVX1_LOC_9/Y 0.06fF
C12084 NAND2X1_LOC_679/B NAND2X1_LOC_728/A 0.05fF
C12085 INVX1_LOC_367/A INVX1_LOC_199/A 0.00fF
C12086 VDD INVX1_LOC_74/A -0.00fF
C12087 INVX1_LOC_686/A INVX1_LOC_66/A 0.01fF
C12088 INVX1_LOC_594/Y INVX1_LOC_479/A 0.03fF
C12089 INVX1_LOC_21/Y INVX1_LOC_327/Y 0.28fF
C12090 INVX1_LOC_93/Y NAND2X1_LOC_677/Y 0.01fF
C12091 INVX1_LOC_121/Y INVX1_LOC_479/A 0.01fF
C12092 NAND2X1_LOC_274/B INVX1_LOC_624/A 0.01fF
C12093 INVX1_LOC_417/Y INVX1_LOC_46/Y 0.20fF
C12094 INVX1_LOC_555/A NAND2X1_LOC_513/A 0.03fF
C12095 INVX1_LOC_469/Y INVX1_LOC_115/A 0.00fF
C12096 INVX1_LOC_206/Y NAND2X1_LOC_621/B 0.01fF
C12097 INVX1_LOC_211/Y INVX1_LOC_48/Y 0.08fF
C12098 INVX1_LOC_175/Y INVX1_LOC_183/A 0.00fF
C12099 NAND2X1_LOC_387/Y INVX1_LOC_145/Y 0.04fF
C12100 INVX1_LOC_318/A INVX1_LOC_99/Y 0.01fF
C12101 INVX1_LOC_53/Y INVX1_LOC_199/Y 4.03fF
C12102 INVX1_LOC_54/Y INVX1_LOC_548/A 0.10fF
C12103 INVX1_LOC_449/A NAND2X1_LOC_178/a_36_24# 0.00fF
C12104 NAND2X1_LOC_294/Y INVX1_LOC_7/Y 0.00fF
C12105 INVX1_LOC_360/A INVX1_LOC_440/Y 0.04fF
C12106 INVX1_LOC_21/Y NAND2X1_LOC_388/A 0.13fF
C12107 NAND2X1_LOC_318/A INVX1_LOC_77/A 0.02fF
C12108 INVX1_LOC_451/A INVX1_LOC_382/A 0.03fF
C12109 INVX1_LOC_45/Y INVX1_LOC_166/Y 0.01fF
C12110 INPUT_3 INVX1_LOC_9/Y 0.25fF
C12111 INVX1_LOC_300/A NAND2X1_LOC_422/a_36_24# 0.00fF
C12112 INVX1_LOC_156/Y INVX1_LOC_26/Y 0.01fF
C12113 INVX1_LOC_12/Y NAND2X1_LOC_542/A 0.34fF
C12114 INVX1_LOC_206/Y NAND2X1_LOC_646/B 0.02fF
C12115 INVX1_LOC_89/Y INVX1_LOC_516/A 0.00fF
C12116 INVX1_LOC_166/A INVX1_LOC_251/Y 0.01fF
C12117 INVX1_LOC_76/Y INVX1_LOC_100/Y 0.14fF
C12118 INVX1_LOC_479/A INVX1_LOC_253/A 0.03fF
C12119 INVX1_LOC_397/Y INVX1_LOC_99/Y 0.04fF
C12120 NAND2X1_LOC_318/A INVX1_LOC_79/A 0.00fF
C12121 INVX1_LOC_455/A INVX1_LOC_18/Y 0.05fF
C12122 INVX1_LOC_45/Y INVX1_LOC_62/Y 8.35fF
C12123 INVX1_LOC_268/Y INVX1_LOC_79/A 0.00fF
C12124 INVX1_LOC_17/Y INVX1_LOC_261/Y 0.03fF
C12125 INVX1_LOC_106/A INVX1_LOC_58/Y 0.01fF
C12126 NAND2X1_LOC_498/B INVX1_LOC_74/Y 0.00fF
C12127 INVX1_LOC_378/Y NAND2X1_LOC_416/Y 0.01fF
C12128 INVX1_LOC_46/Y INVX1_LOC_48/Y 0.03fF
C12129 INVX1_LOC_649/Y INVX1_LOC_643/Y 0.05fF
C12130 INVX1_LOC_277/A INVX1_LOC_283/A 0.03fF
C12131 INVX1_LOC_586/A INVX1_LOC_75/Y 0.03fF
C12132 INVX1_LOC_17/Y INVX1_LOC_258/Y 0.04fF
C12133 INVX1_LOC_54/Y INVX1_LOC_31/Y 0.28fF
C12134 INVX1_LOC_95/A INVX1_LOC_99/Y 0.00fF
C12135 INVX1_LOC_137/Y NAND2X1_LOC_803/a_36_24# 0.00fF
C12136 NAND2X1_LOC_187/a_36_24# INVX1_LOC_48/Y 0.01fF
C12137 INVX1_LOC_166/A INVX1_LOC_608/A 0.01fF
C12138 INVX1_LOC_45/Y INVX1_LOC_529/Y 0.01fF
C12139 NAND2X1_LOC_344/B INVX1_LOC_453/Y 0.16fF
C12140 NAND2X1_LOC_56/Y INVX1_LOC_90/Y 0.01fF
C12141 INVX1_LOC_76/Y INVX1_LOC_74/Y 6.36fF
C12142 INVX1_LOC_356/A INVX1_LOC_505/Y 0.14fF
C12143 INVX1_LOC_587/Y NAND2X1_LOC_837/A 0.11fF
C12144 INVX1_LOC_602/A INVX1_LOC_41/Y 0.07fF
C12145 INVX1_LOC_93/Y INVX1_LOC_199/A 0.01fF
C12146 INVX1_LOC_361/Y NAND2X1_LOC_307/B 0.01fF
C12147 NAND2X1_LOC_845/B INVX1_LOC_145/Y 0.01fF
C12148 INVX1_LOC_93/Y INVX1_LOC_89/Y 0.97fF
C12149 NAND2X1_LOC_785/a_36_24# INVX1_LOC_26/Y 0.00fF
C12150 INVX1_LOC_318/A INVX1_LOC_47/Y 0.01fF
C12151 INVX1_LOC_589/Y INVX1_LOC_397/Y 0.11fF
C12152 INVX1_LOC_312/Y INVX1_LOC_75/Y 0.07fF
C12153 NAND2X1_LOC_181/A INVX1_LOC_387/Y 0.00fF
C12154 INVX1_LOC_49/Y INVX1_LOC_350/Y 0.03fF
C12155 INVX1_LOC_442/Y INVX1_LOC_502/A 0.01fF
C12156 INVX1_LOC_53/A INVX1_LOC_26/Y 0.39fF
C12157 INVX1_LOC_42/Y NAND2X1_LOC_80/a_36_24# 0.00fF
C12158 INVX1_LOC_202/Y INVX1_LOC_77/A 0.01fF
C12159 INVX1_LOC_544/Y INVX1_LOC_105/Y 0.15fF
C12160 INVX1_LOC_166/A INVX1_LOC_58/Y 0.03fF
C12161 INVX1_LOC_586/A NAND2X1_LOC_271/A 0.09fF
C12162 INVX1_LOC_93/Y INVX1_LOC_501/A 0.03fF
C12163 NAND2X1_LOC_181/A INVX1_LOC_49/Y 0.02fF
C12164 INVX1_LOC_32/Y INVX1_LOC_206/A 0.03fF
C12165 INVX1_LOC_128/Y INVX1_LOC_50/Y 0.03fF
C12166 INVX1_LOC_26/Y INVX1_LOC_50/Y 0.17fF
C12167 INVX1_LOC_173/Y INVX1_LOC_223/Y 0.00fF
C12168 INVX1_LOC_77/Y INVX1_LOC_351/Y 0.05fF
C12169 INVX1_LOC_417/Y INVX1_LOC_75/A 0.01fF
C12170 INVX1_LOC_99/Y INVX1_LOC_588/A 0.09fF
C12171 INVX1_LOC_134/Y NAND2X1_LOC_832/A 0.11fF
C12172 INVX1_LOC_497/A NAND2X1_LOC_637/a_36_24# 0.02fF
C12173 INVX1_LOC_317/A INVX1_LOC_245/A 0.00fF
C12174 INVX1_LOC_74/Y NAND2X1_LOC_446/a_36_24# 0.00fF
C12175 INVX1_LOC_456/Y INVX1_LOC_74/A 0.10fF
C12176 NAND2X1_LOC_631/B INVX1_LOC_381/Y 0.11fF
C12177 INVX1_LOC_662/A GATE_662 0.03fF
C12178 INVX1_LOC_214/Y NAND2X1_LOC_248/B 0.09fF
C12179 INVX1_LOC_342/Y NAND2X1_LOC_451/B 0.03fF
C12180 INVX1_LOC_675/A INVX1_LOC_501/A 0.07fF
C12181 INVX1_LOC_117/Y INVX1_LOC_41/Y 2.38fF
C12182 NAND2X1_LOC_603/a_36_24# INVX1_LOC_347/A 0.00fF
C12183 INVX1_LOC_239/A NAND2X1_LOC_342/B 0.03fF
C12184 INVX1_LOC_662/A NAND2X1_LOC_846/B 0.28fF
C12185 INVX1_LOC_89/A INVX1_LOC_9/Y 0.04fF
C12186 INVX1_LOC_48/Y INVX1_LOC_75/A 0.01fF
C12187 INVX1_LOC_153/Y INVX1_LOC_58/Y 0.01fF
C12188 INVX1_LOC_49/Y INVX1_LOC_79/A 10.98fF
C12189 INVX1_LOC_531/Y INVX1_LOC_58/Y 0.18fF
C12190 INVX1_LOC_556/Y INVX1_LOC_92/A 2.82fF
C12191 INVX1_LOC_47/Y INVX1_LOC_588/A 0.07fF
C12192 INVX1_LOC_112/Y INVX1_LOC_114/A 0.06fF
C12193 INVX1_LOC_369/Y INVX1_LOC_90/Y 0.05fF
C12194 INVX1_LOC_32/Y INVX1_LOC_636/A 0.07fF
C12195 INVX1_LOC_204/Y INVX1_LOC_622/Y 0.01fF
C12196 INVX1_LOC_44/Y NAND2X1_LOC_227/A 0.05fF
C12197 INVX1_LOC_119/Y INVX1_LOC_588/A 0.01fF
C12198 NAND2X1_LOC_475/A INVX1_LOC_65/Y 0.08fF
C12199 INVX1_LOC_206/Y INVX1_LOC_442/A 0.07fF
C12200 VDD INVX1_LOC_144/Y 0.26fF
C12201 INVX1_LOC_26/Y INVX1_LOC_658/Y 0.03fF
C12202 INPUT_0 INVX1_LOC_542/A 0.34fF
C12203 VDD INVX1_LOC_398/A 0.00fF
C12204 NAND2X1_LOC_370/a_36_24# INVX1_LOC_270/A 0.00fF
C12205 VDD INVX1_LOC_101/Y 0.21fF
C12206 NAND2X1_LOC_609/B NAND2X1_LOC_646/B 0.02fF
C12207 INVX1_LOC_558/A NAND2X1_LOC_513/Y 0.11fF
C12208 VDD INVX1_LOC_10/Y 0.21fF
C12209 INVX1_LOC_420/Y INVX1_LOC_134/Y 0.00fF
C12210 INVX1_LOC_21/Y NAND2X1_LOC_393/a_36_24# 0.01fF
C12211 INVX1_LOC_287/A NAND2X1_LOC_475/A 0.12fF
C12212 INVX1_LOC_547/A INVX1_LOC_45/Y 0.01fF
C12213 VDD NAND2X1_LOC_697/Y 0.03fF
C12214 NAND2X1_LOC_56/a_36_24# INVX1_LOC_206/Y 0.00fF
C12215 VDD INVX1_LOC_451/A 2.60fF
C12216 VDD INVX1_LOC_685/Y 0.27fF
C12217 INVX1_LOC_442/A INVX1_LOC_686/A 1.01fF
C12218 INVX1_LOC_438/A INVX1_LOC_444/Y 0.07fF
C12219 NAND2X1_LOC_307/A INVX1_LOC_618/Y 0.00fF
C12220 INVX1_LOC_446/A INVX1_LOC_421/A 0.05fF
C12221 INVX1_LOC_206/Y INVX1_LOC_116/Y 0.07fF
C12222 INVX1_LOC_438/Y INVX1_LOC_452/A 0.07fF
C12223 INVX1_LOC_206/Y INVX1_LOC_544/A 0.01fF
C12224 INVX1_LOC_257/Y INVX1_LOC_504/Y 0.01fF
C12225 VDD INVX1_LOC_665/Y 0.57fF
C12226 INVX1_LOC_273/A NAND2X1_LOC_238/a_36_24# 0.01fF
C12227 VDD INVX1_LOC_575/Y 0.22fF
C12228 INVX1_LOC_32/A INVX1_LOC_48/Y 0.06fF
C12229 INVX1_LOC_412/Y INVX1_LOC_360/A 0.02fF
C12230 INVX1_LOC_410/Y INVX1_LOC_304/A 0.12fF
C12231 NAND2X1_LOC_173/Y INVX1_LOC_134/Y 0.05fF
C12232 NAND2X1_LOC_534/Y INVX1_LOC_31/Y 0.01fF
C12233 INVX1_LOC_628/Y NAND2X1_LOC_122/Y 0.15fF
C12234 INVX1_LOC_419/Y INVX1_LOC_412/A 0.18fF
C12235 NAND2X1_LOC_780/B INVX1_LOC_93/Y 0.01fF
C12236 NAND2X1_LOC_498/Y INVX1_LOC_506/Y 0.02fF
C12237 VDD NAND2X1_LOC_308/A 0.14fF
C12238 INVX1_LOC_447/Y INVX1_LOC_51/Y 0.05fF
C12239 INVX1_LOC_619/A INVX1_LOC_191/A 0.03fF
C12240 INVX1_LOC_562/Y INVX1_LOC_565/A 0.15fF
C12241 NAND2X1_LOC_460/A INVX1_LOC_311/Y 0.01fF
C12242 INVX1_LOC_20/Y INVX1_LOC_154/Y 0.00fF
C12243 VDD INVX1_LOC_132/A -0.00fF
C12244 INPUT_0 NAND2X1_LOC_707/B 0.00fF
C12245 INVX1_LOC_414/A INVX1_LOC_387/Y 0.00fF
C12246 INVX1_LOC_683/Y INVX1_LOC_371/Y 0.02fF
C12247 INVX1_LOC_564/Y INVX1_LOC_50/Y 0.01fF
C12248 INVX1_LOC_381/A INVX1_LOC_7/Y 0.19fF
C12249 NAND2X1_LOC_190/A INVX1_LOC_45/Y 0.05fF
C12250 INVX1_LOC_335/Y INVX1_LOC_111/A 0.09fF
C12251 INVX1_LOC_80/A INVX1_LOC_519/A 0.03fF
C12252 NAND2X1_LOC_318/A INVX1_LOC_59/Y 0.25fF
C12253 INVX1_LOC_554/A INVX1_LOC_662/A 0.05fF
C12254 INVX1_LOC_26/A INVX1_LOC_18/Y 0.01fF
C12255 NAND2X1_LOC_615/Y INVX1_LOC_596/Y 0.07fF
C12256 INVX1_LOC_482/Y INVX1_LOC_388/Y 0.01fF
C12257 INVX1_LOC_26/Y INVX1_LOC_275/A 0.03fF
C12258 INVX1_LOC_651/Y INVX1_LOC_679/A 0.02fF
C12259 INVX1_LOC_459/Y INVX1_LOC_460/Y 0.17fF
C12260 INVX1_LOC_335/Y INVX1_LOC_602/A 0.08fF
C12261 INVX1_LOC_268/Y INVX1_LOC_59/Y 0.54fF
C12262 NAND2X1_LOC_538/B INVX1_LOC_230/A 0.05fF
C12263 INVX1_LOC_224/Y INVX1_LOC_69/Y 0.14fF
C12264 NAND2X1_LOC_513/Y INVX1_LOC_46/Y 0.12fF
C12265 INVX1_LOC_206/Y INVX1_LOC_255/A 0.01fF
C12266 INVX1_LOC_395/A INVX1_LOC_89/Y 1.46fF
C12267 INVX1_LOC_54/Y INVX1_LOC_51/Y 0.23fF
C12268 NAND2X1_LOC_45/Y INVX1_LOC_63/Y 0.20fF
C12269 INVX1_LOC_269/Y INVX1_LOC_32/Y 0.04fF
C12270 INVX1_LOC_556/A NAND2X1_LOC_128/B 0.03fF
C12271 NAND2X1_LOC_174/a_36_24# INVX1_LOC_566/A 0.00fF
C12272 NAND2X1_LOC_863/a_36_24# INVX1_LOC_684/A 0.02fF
C12273 INVX1_LOC_542/A INVX1_LOC_498/A 0.03fF
C12274 NAND2X1_LOC_318/A INVX1_LOC_48/Y 3.33fF
C12275 INVX1_LOC_315/Y INVX1_LOC_117/Y 0.05fF
C12276 INVX1_LOC_489/A NAND2X1_LOC_416/Y 0.01fF
C12277 INVX1_LOC_686/A INVX1_LOC_116/Y 0.50fF
C12278 NAND2X1_LOC_498/Y INVX1_LOC_253/Y 0.00fF
C12279 INVX1_LOC_578/A INVX1_LOC_69/Y 0.16fF
C12280 NAND2X1_LOC_318/B INVX1_LOC_600/A 0.01fF
C12281 INVX1_LOC_435/A INVX1_LOC_312/A 0.03fF
C12282 INVX1_LOC_235/Y INVX1_LOC_681/Y 0.01fF
C12283 INVX1_LOC_206/Y INVX1_LOC_179/A 0.18fF
C12284 INVX1_LOC_435/A NAND2X1_LOC_391/A 0.01fF
C12285 NAND2X1_LOC_457/A INVX1_LOC_682/A 0.03fF
C12286 INVX1_LOC_266/A INVX1_LOC_54/Y 0.01fF
C12287 INVX1_LOC_469/Y INVX1_LOC_76/Y 0.04fF
C12288 INVX1_LOC_416/A NAND2X1_LOC_336/B 0.02fF
C12289 INVX1_LOC_235/Y INPUT_1 0.07fF
C12290 INVX1_LOC_510/Y NAND2X1_LOC_308/A 0.02fF
C12291 INVX1_LOC_419/Y NAND2X1_LOC_336/B 0.01fF
C12292 INVX1_LOC_438/A INVX1_LOC_26/Y 0.07fF
C12293 INVX1_LOC_381/A INVX1_LOC_32/Y 0.07fF
C12294 INVX1_LOC_515/A INVX1_LOC_463/Y 0.01fF
C12295 NAND2X1_LOC_498/Y INVX1_LOC_63/Y 0.12fF
C12296 INVX1_LOC_224/Y INVX1_LOC_247/Y 0.16fF
C12297 INVX1_LOC_300/A INVX1_LOC_154/Y 0.01fF
C12298 INVX1_LOC_490/Y INVX1_LOC_328/Y 0.03fF
C12299 INVX1_LOC_570/A INVX1_LOC_63/Y 0.13fF
C12300 INVX1_LOC_11/Y INVX1_LOC_519/A 0.01fF
C12301 INVX1_LOC_556/Y INVX1_LOC_679/Y 0.03fF
C12302 INVX1_LOC_395/A INVX1_LOC_179/Y 0.02fF
C12303 INVX1_LOC_158/A INVX1_LOC_79/A 0.01fF
C12304 INVX1_LOC_53/Y INVX1_LOC_460/Y 0.06fF
C12305 INVX1_LOC_54/Y INVX1_LOC_365/Y 0.02fF
C12306 INVX1_LOC_17/Y INVX1_LOC_442/Y 0.07fF
C12307 INPUT_0 INVX1_LOC_114/A 0.00fF
C12308 INVX1_LOC_11/Y INVX1_LOC_323/Y 0.58fF
C12309 INVX1_LOC_513/Y INVX1_LOC_586/A 0.03fF
C12310 INVX1_LOC_424/Y NAND2X1_LOC_294/Y 0.03fF
C12311 INVX1_LOC_369/A INVX1_LOC_50/Y 0.03fF
C12312 INVX1_LOC_266/A INVX1_LOC_257/A 0.45fF
C12313 INVX1_LOC_202/Y INVX1_LOC_59/Y 0.64fF
C12314 INVX1_LOC_317/Y INVX1_LOC_245/A 0.21fF
C12315 INVX1_LOC_115/Y INVX1_LOC_440/Y 0.09fF
C12316 INVX1_LOC_99/Y NAND2X1_LOC_646/A 0.01fF
C12317 NAND2X1_LOC_467/A INVX1_LOC_58/Y 0.01fF
C12318 INVX1_LOC_21/Y INVX1_LOC_117/Y 0.04fF
C12319 NAND2X1_LOC_538/a_36_24# INVX1_LOC_99/Y 0.01fF
C12320 NAND2X1_LOC_451/a_36_24# INVX1_LOC_505/A 0.00fF
C12321 INVX1_LOC_255/A INVX1_LOC_686/A 0.02fF
C12322 INVX1_LOC_202/Y INVX1_LOC_48/Y 0.22fF
C12323 INVX1_LOC_17/Y INVX1_LOC_671/A 0.82fF
C12324 NAND2X1_LOC_498/B INVX1_LOC_79/A 0.02fF
C12325 INVX1_LOC_545/A INVX1_LOC_361/Y 0.10fF
C12326 INVX1_LOC_316/Y INVX1_LOC_341/Y 0.18fF
C12327 INVX1_LOC_76/Y NAND2X1_LOC_558/B 0.02fF
C12328 INVX1_LOC_556/Y INPUT_1 0.03fF
C12329 INVX1_LOC_550/Y INVX1_LOC_48/Y 0.01fF
C12330 INVX1_LOC_47/Y INVX1_LOC_670/Y 0.01fF
C12331 INVX1_LOC_619/A INVX1_LOC_182/Y 0.03fF
C12332 NAND2X1_LOC_180/B INVX1_LOC_242/Y 0.05fF
C12333 INVX1_LOC_49/Y INVX1_LOC_632/A 0.07fF
C12334 INVX1_LOC_76/Y INVX1_LOC_79/A 0.07fF
C12335 INVX1_LOC_368/A INVX1_LOC_235/Y 0.02fF
C12336 INVX1_LOC_276/A INVX1_LOC_100/Y 0.00fF
C12337 INVX1_LOC_550/A INVX1_LOC_48/Y 0.03fF
C12338 INVX1_LOC_48/Y NAND2X1_LOC_213/a_36_24# 0.00fF
C12339 NAND2X1_LOC_526/Y INVX1_LOC_479/A 0.00fF
C12340 INVX1_LOC_49/Y INVX1_LOC_509/Y 0.05fF
C12341 INVX1_LOC_54/Y INVX1_LOC_254/A 0.01fF
C12342 INVX1_LOC_498/A INVX1_LOC_259/Y 0.01fF
C12343 NAND2X1_LOC_274/B NAND2X1_LOC_273/a_36_24# 0.02fF
C12344 INVX1_LOC_117/Y NAND2X1_LOC_267/A 0.01fF
C12345 INVX1_LOC_63/Y INVX1_LOC_99/Y 0.83fF
C12346 INVX1_LOC_387/Y INVX1_LOC_48/Y 0.00fF
C12347 INVX1_LOC_49/Y INVX1_LOC_59/Y 0.00fF
C12348 NAND2X1_LOC_137/A INVX1_LOC_117/Y 0.03fF
C12349 NAND2X1_LOC_33/a_36_24# INVX1_LOC_26/Y 0.00fF
C12350 INVX1_LOC_188/Y INVX1_LOC_242/Y 0.01fF
C12351 INVX1_LOC_549/Y INVX1_LOC_168/Y 0.05fF
C12352 INVX1_LOC_293/Y INVX1_LOC_62/Y 9.19fF
C12353 NAND2X1_LOC_184/Y INVX1_LOC_6/Y 0.48fF
C12354 INVX1_LOC_261/Y INVX1_LOC_497/Y 0.23fF
C12355 INVX1_LOC_211/Y NAND2X1_LOC_615/Y 0.11fF
C12356 INVX1_LOC_670/Y INVX1_LOC_119/Y 0.01fF
C12357 NAND2X1_LOC_527/Y INVX1_LOC_69/Y 0.01fF
C12358 NAND2X1_LOC_557/B INVX1_LOC_86/Y 0.03fF
C12359 INVX1_LOC_49/Y INVX1_LOC_48/Y 7.49fF
C12360 INVX1_LOC_298/A INVX1_LOC_204/Y 0.00fF
C12361 INVX1_LOC_89/Y INVX1_LOC_31/Y 0.24fF
C12362 NAND2X1_LOC_399/B INVX1_LOC_100/Y 0.19fF
C12363 INVX1_LOC_435/A INVX1_LOC_226/Y 0.04fF
C12364 INVX1_LOC_390/A INVX1_LOC_194/Y 0.01fF
C12365 INVX1_LOC_75/Y INVX1_LOC_486/Y 0.09fF
C12366 NAND2X1_LOC_673/B INVX1_LOC_9/Y 1.68fF
C12367 INVX1_LOC_100/Y INVX1_LOC_7/Y 0.07fF
C12368 INVX1_LOC_466/A INVX1_LOC_58/Y 0.25fF
C12369 INVX1_LOC_117/Y INVX1_LOC_107/Y 0.02fF
C12370 INVX1_LOC_93/Y INVX1_LOC_44/Y 0.03fF
C12371 NAND2X1_LOC_542/A INVX1_LOC_66/A 0.04fF
C12372 INVX1_LOC_134/Y INVX1_LOC_354/A 0.02fF
C12373 INVX1_LOC_123/A INVX1_LOC_63/Y 0.01fF
C12374 INVX1_LOC_386/Y NAND2X1_LOC_631/B 0.05fF
C12375 INVX1_LOC_588/Y INVX1_LOC_245/A 0.03fF
C12376 INVX1_LOC_589/Y INVX1_LOC_63/Y 0.03fF
C12377 INVX1_LOC_89/Y NAND2X1_LOC_675/B 0.23fF
C12378 NAND2X1_LOC_615/Y INVX1_LOC_46/Y 0.02fF
C12379 INVX1_LOC_31/Y INVX1_LOC_501/A 0.07fF
C12380 INVX1_LOC_634/A INVX1_LOC_634/Y 0.01fF
C12381 INVX1_LOC_41/Y INVX1_LOC_178/A 0.07fF
C12382 INVX1_LOC_47/Y INVX1_LOC_63/Y 0.31fF
C12383 NAND2X1_LOC_698/Y INVX1_LOC_199/Y 0.06fF
C12384 NAND2X1_LOC_557/B INVX1_LOC_63/Y 0.12fF
C12385 INVX1_LOC_376/Y INVX1_LOC_66/A 0.07fF
C12386 NAND2X1_LOC_819/a_36_24# INVX1_LOC_655/A 0.01fF
C12387 NAND2X1_LOC_847/A NAND2X1_LOC_342/A 0.05fF
C12388 INVX1_LOC_41/Y NAND2X1_LOC_76/A 0.01fF
C12389 INVX1_LOC_59/Y INVX1_LOC_92/Y 0.02fF
C12390 INVX1_LOC_251/A INVX1_LOC_479/A 0.04fF
C12391 INVX1_LOC_32/Y INVX1_LOC_100/Y 1.25fF
C12392 INVX1_LOC_620/A INVX1_LOC_273/Y 0.00fF
C12393 INVX1_LOC_662/A INVX1_LOC_199/Y 0.02fF
C12394 INVX1_LOC_608/A INVX1_LOC_41/Y 0.01fF
C12395 INVX1_LOC_48/Y INVX1_LOC_92/Y 0.01fF
C12396 INVX1_LOC_513/A INVX1_LOC_505/Y 0.00fF
C12397 INVX1_LOC_187/Y INVX1_LOC_90/Y 0.00fF
C12398 INVX1_LOC_49/Y NAND2X1_LOC_434/B 0.01fF
C12399 INVX1_LOC_100/Y NAND2X1_LOC_815/a_36_24# 0.00fF
C12400 INVX1_LOC_32/Y INVX1_LOC_74/Y 2.91fF
C12401 INVX1_LOC_63/Y INVX1_LOC_119/Y 0.07fF
C12402 INVX1_LOC_446/A NAND2X1_LOC_45/Y 0.10fF
C12403 INVX1_LOC_63/Y NAND2X1_LOC_66/Y 0.07fF
C12404 INVX1_LOC_32/Y INVX1_LOC_483/Y 0.02fF
C12405 NAND2X1_LOC_271/a_36_24# INVX1_LOC_41/Y 0.00fF
C12406 NAND2X1_LOC_663/a_36_24# NAND2X1_LOC_843/B 0.00fF
C12407 INVX1_LOC_6/Y INVX1_LOC_75/Y 0.00fF
C12408 INVX1_LOC_426/Y INVX1_LOC_438/A 0.04fF
C12409 INVX1_LOC_41/Y INVX1_LOC_58/Y 1.48fF
C12410 NAND2X1_LOC_335/B NAND2X1_LOC_76/B 0.03fF
C12411 NAND2X1_LOC_707/B INVX1_LOC_464/Y 0.12fF
C12412 INVX1_LOC_153/Y INVX1_LOC_245/A 0.03fF
C12413 VDD INVX1_LOC_238/Y 0.14fF
C12414 NAND2X1_LOC_601/Y INVX1_LOC_376/Y 0.02fF
C12415 VDD INVX1_LOC_264/Y 0.21fF
C12416 NAND2X1_LOC_628/Y INVX1_LOC_90/Y 0.02fF
C12417 INVX1_LOC_15/Y INVX1_LOC_588/A 0.01fF
C12418 NAND2X1_LOC_543/B INVX1_LOC_65/Y 0.04fF
C12419 INPUT_0 NAND2X1_LOC_457/A 0.03fF
C12420 INVX1_LOC_279/A NAND2X1_LOC_261/Y 0.01fF
C12421 VDD INVX1_LOC_364/Y 0.22fF
C12422 INVX1_LOC_652/A INVX1_LOC_479/A 0.01fF
C12423 INVX1_LOC_68/Y NAND2X1_LOC_76/B 0.00fF
C12424 NAND2X1_LOC_475/A NAND2X1_LOC_335/a_36_24# 0.00fF
C12425 VDD INVX1_LOC_5/Y 0.23fF
C12426 INVX1_LOC_224/Y INVX1_LOC_586/A 0.13fF
C12427 INVX1_LOC_404/Y INVX1_LOC_45/Y 1.00fF
C12428 INVX1_LOC_395/A INVX1_LOC_137/A 0.02fF
C12429 NAND2X1_LOC_498/Y INVX1_LOC_374/A 0.08fF
C12430 NAND2X1_LOC_405/a_36_24# INVX1_LOC_636/A 0.01fF
C12431 INVX1_LOC_274/A INVX1_LOC_615/A 0.29fF
C12432 VDD NAND2X1_LOC_379/Y 0.02fF
C12433 INVX1_LOC_578/A INVX1_LOC_586/A 0.12fF
C12434 VDD INVX1_LOC_134/Y 3.64fF
C12435 INVX1_LOC_271/Y INVX1_LOC_45/Y 0.09fF
C12436 VDD NAND2X1_LOC_48/Y 0.01fF
C12437 VDD INVX1_LOC_47/A 0.00fF
C12438 INVX1_LOC_224/Y INVX1_LOC_312/Y 0.12fF
C12439 INVX1_LOC_118/Y INVX1_LOC_367/A 0.01fF
C12440 INVX1_LOC_360/Y INVX1_LOC_638/A 0.03fF
C12441 INVX1_LOC_400/Y INVX1_LOC_84/A 0.07fF
C12442 VDD INVX1_LOC_316/Y 0.21fF
C12443 INVX1_LOC_447/A NAND2X1_LOC_179/Y 0.01fF
C12444 INVX1_LOC_625/A NAND2X1_LOC_335/B 0.03fF
C12445 INVX1_LOC_312/Y INVX1_LOC_578/A 0.07fF
C12446 INVX1_LOC_564/Y INVX1_LOC_187/A 0.00fF
C12447 NAND2X1_LOC_790/B INVX1_LOC_50/Y 0.00fF
C12448 NAND2X1_LOC_69/B INVX1_LOC_46/Y 0.00fF
C12449 INVX1_LOC_205/Y INVX1_LOC_395/A 0.02fF
C12450 INVX1_LOC_54/Y NAND2X1_LOC_537/A 0.11fF
C12451 INVX1_LOC_32/Y NAND2X1_LOC_591/B 0.01fF
C12452 INVX1_LOC_201/Y INVX1_LOC_97/A 0.03fF
C12453 INVX1_LOC_552/Y INVX1_LOC_99/Y 0.01fF
C12454 INVX1_LOC_510/Y INVX1_LOC_134/Y 0.09fF
C12455 INVX1_LOC_412/Y INVX1_LOC_350/A 0.02fF
C12456 INVX1_LOC_438/Y INVX1_LOC_282/A 0.03fF
C12457 INVX1_LOC_450/A INVX1_LOC_7/Y 0.03fF
C12458 INVX1_LOC_185/A INVX1_LOC_555/A 0.02fF
C12459 NAND2X1_LOC_97/A INVX1_LOC_80/A 0.02fF
C12460 VDD NAND2X1_LOC_165/Y 0.01fF
C12461 INVX1_LOC_400/Y INVX1_LOC_129/A 0.07fF
C12462 INVX1_LOC_158/A INVX1_LOC_48/Y 0.01fF
C12463 INVX1_LOC_426/A INVX1_LOC_89/Y 0.40fF
C12464 INVX1_LOC_555/Y INVX1_LOC_53/Y 0.01fF
C12465 INVX1_LOC_586/A INVX1_LOC_358/A 0.13fF
C12466 INVX1_LOC_374/A INVX1_LOC_99/Y 0.06fF
C12467 NAND2X1_LOC_122/Y NAND2X1_LOC_802/a_36_24# 0.00fF
C12468 NAND2X1_LOC_764/Y INVX1_LOC_48/Y 0.01fF
C12469 INVX1_LOC_236/A INVX1_LOC_523/A 0.05fF
C12470 INVX1_LOC_395/A INVX1_LOC_194/Y 0.10fF
C12471 NAND2X1_LOC_242/A INVX1_LOC_32/Y 0.01fF
C12472 NAND2X1_LOC_837/a_36_24# INVX1_LOC_59/A 0.00fF
C12473 INVX1_LOC_79/A INVX1_LOC_192/A 0.01fF
C12474 INVX1_LOC_68/Y INVX1_LOC_625/A 0.02fF
C12475 INVX1_LOC_118/Y INVX1_LOC_93/Y 0.07fF
C12476 INVX1_LOC_127/A INVX1_LOC_361/Y 0.09fF
C12477 INVX1_LOC_98/A INVX1_LOC_59/Y 0.00fF
C12478 INVX1_LOC_20/Y INVX1_LOC_603/Y 0.01fF
C12479 INVX1_LOC_150/Y INVX1_LOC_500/Y 0.05fF
C12480 VDD INVX1_LOC_65/A 0.00fF
C12481 INVX1_LOC_287/Y INVX1_LOC_155/Y 0.05fF
C12482 INVX1_LOC_45/Y INVX1_LOC_480/Y 0.01fF
C12483 INVX1_LOC_255/Y INVX1_LOC_117/Y 0.01fF
C12484 INVX1_LOC_76/Y INVX1_LOC_59/Y 2.35fF
C12485 INVX1_LOC_384/A INVX1_LOC_453/Y 0.07fF
C12486 INVX1_LOC_53/Y NAND2X1_LOC_148/A 0.01fF
C12487 INVX1_LOC_206/Y INVX1_LOC_69/Y 0.42fF
C12488 NAND2X1_LOC_475/A INVX1_LOC_63/Y 0.08fF
C12489 INVX1_LOC_560/A NAND2X1_LOC_388/A 0.06fF
C12490 INVX1_LOC_259/A INVX1_LOC_260/Y 0.00fF
C12491 INVX1_LOC_404/Y NAND2X1_LOC_276/A 0.01fF
C12492 INVX1_LOC_666/Y INVX1_LOC_109/Y 0.03fF
C12493 NAND2X1_LOC_147/B INVX1_LOC_80/A 0.02fF
C12494 NAND2X1_LOC_788/A INVX1_LOC_376/Y 0.08fF
C12495 INVX1_LOC_552/Y INVX1_LOC_47/Y 0.02fF
C12496 NAND2X1_LOC_527/Y INVX1_LOC_586/A 0.00fF
C12497 NAND2X1_LOC_526/Y NAND2X1_LOC_521/Y 0.01fF
C12498 INVX1_LOC_103/Y INVX1_LOC_364/Y 0.03fF
C12499 INVX1_LOC_628/Y INVX1_LOC_579/A 0.01fF
C12500 INVX1_LOC_45/Y INVX1_LOC_169/Y 0.11fF
C12501 INVX1_LOC_656/Y INVX1_LOC_59/A 0.01fF
C12502 INVX1_LOC_76/Y INVX1_LOC_48/Y 0.26fF
C12503 INVX1_LOC_561/Y INVX1_LOC_49/Y 0.03fF
C12504 INVX1_LOC_607/Y INVX1_LOC_651/A 0.01fF
C12505 NAND2X1_LOC_770/A INVX1_LOC_79/A 0.01fF
C12506 NAND2X1_LOC_13/Y INVX1_LOC_54/Y 0.03fF
C12507 INVX1_LOC_51/Y INVX1_LOC_199/A 0.01fF
C12508 NAND2X1_LOC_307/A NAND2X1_LOC_317/a_36_24# 0.00fF
C12509 INVX1_LOC_435/A INVX1_LOC_297/A 0.00fF
C12510 NAND2X1_LOC_190/A INVX1_LOC_293/Y 0.04fF
C12511 INVX1_LOC_224/Y INVX1_LOC_225/Y 0.01fF
C12512 INVX1_LOC_442/A NAND2X1_LOC_542/A 0.02fF
C12513 INVX1_LOC_625/A INVX1_LOC_600/A 0.02fF
C12514 INVX1_LOC_134/Y INVX1_LOC_509/A 0.02fF
C12515 INVX1_LOC_442/Y INVX1_LOC_232/Y 0.03fF
C12516 INVX1_LOC_395/A INVX1_LOC_44/Y 0.23fF
C12517 INVX1_LOC_20/Y NAND2X1_LOC_387/Y 0.08fF
C12518 INVX1_LOC_21/Y INVX1_LOC_281/Y 0.10fF
C12519 INVX1_LOC_603/Y INVX1_LOC_300/A 0.02fF
C12520 INVX1_LOC_89/Y INVX1_LOC_51/Y 0.28fF
C12521 INVX1_LOC_235/Y INVX1_LOC_50/Y 0.08fF
C12522 NAND2X1_LOC_122/Y INVX1_LOC_261/Y 0.01fF
C12523 INVX1_LOC_367/Y NAND2X1_LOC_296/Y 0.01fF
C12524 INVX1_LOC_566/A INVX1_LOC_32/Y 0.07fF
C12525 INVX1_LOC_213/Y INVX1_LOC_53/Y 0.99fF
C12526 INVX1_LOC_21/Y INVX1_LOC_178/A 0.04fF
C12527 NAND2X1_LOC_106/B NAND2X1_LOC_496/Y 0.16fF
C12528 NAND2X1_LOC_467/A NAND2X1_LOC_689/B 0.00fF
C12529 INVX1_LOC_257/Y INVX1_LOC_114/A 0.10fF
C12530 INPUT_3 INVX1_LOC_169/Y 0.19fF
C12531 INVX1_LOC_586/A INVX1_LOC_120/Y 0.02fF
C12532 INVX1_LOC_508/Y INVX1_LOC_46/Y 0.02fF
C12533 INVX1_LOC_266/A INVX1_LOC_89/Y 0.18fF
C12534 NAND2X1_LOC_541/B INVX1_LOC_46/Y 0.16fF
C12535 INVX1_LOC_103/Y INVX1_LOC_134/Y 0.14fF
C12536 INVX1_LOC_51/Y INVX1_LOC_501/A 0.03fF
C12537 INVX1_LOC_76/Y NAND2X1_LOC_491/Y 0.04fF
C12538 INVX1_LOC_300/A INVX1_LOC_637/A 0.06fF
C12539 INVX1_LOC_145/Y INVX1_LOC_259/Y 0.03fF
C12540 INVX1_LOC_686/A INVX1_LOC_69/Y 0.24fF
C12541 INVX1_LOC_21/Y INVX1_LOC_608/A 0.00fF
C12542 INVX1_LOC_20/Y NAND2X1_LOC_684/a_36_24# 0.00fF
C12543 INVX1_LOC_374/A INVX1_LOC_119/Y 0.04fF
C12544 INVX1_LOC_254/Y INVX1_LOC_35/Y 1.97fF
C12545 INVX1_LOC_45/Y NAND2X1_LOC_833/B 0.01fF
C12546 INVX1_LOC_288/A INVX1_LOC_114/A 0.06fF
C12547 NAND2X1_LOC_387/Y INVX1_LOC_197/Y 0.07fF
C12548 INVX1_LOC_556/Y INVX1_LOC_50/Y 0.00fF
C12549 INVX1_LOC_20/Y NAND2X1_LOC_845/B 0.00fF
C12550 NAND2X1_LOC_312/a_36_24# INVX1_LOC_75/A 0.00fF
C12551 INVX1_LOC_600/A NAND2X1_LOC_52/Y 0.18fF
C12552 INVX1_LOC_21/Y INVX1_LOC_58/Y 14.10fF
C12553 INVX1_LOC_31/Y INVX1_LOC_194/Y 0.03fF
C12554 INVX1_LOC_204/Y INVX1_LOC_145/Y 0.01fF
C12555 NAND2X1_LOC_542/A INVX1_LOC_116/Y 0.02fF
C12556 INVX1_LOC_53/Y INVX1_LOC_662/A 0.16fF
C12557 INVX1_LOC_45/Y INVX1_LOC_74/A 0.09fF
C12558 INVX1_LOC_602/A INVX1_LOC_26/Y 0.09fF
C12559 INVX1_LOC_592/Y INVX1_LOC_35/Y 0.01fF
C12560 INVX1_LOC_492/A INVX1_LOC_6/Y 0.03fF
C12561 INVX1_LOC_284/A INVX1_LOC_44/Y 0.02fF
C12562 INVX1_LOC_354/Y INVX1_LOC_359/A 0.00fF
C12563 NAND2X1_LOC_383/a_36_24# INVX1_LOC_6/Y -0.00fF
C12564 NAND2X1_LOC_388/A INVX1_LOC_603/A 0.00fF
C12565 INVX1_LOC_287/A INVX1_LOC_353/A 0.15fF
C12566 INVX1_LOC_104/Y INVX1_LOC_26/Y 0.01fF
C12567 INVX1_LOC_183/Y INVX1_LOC_366/Y 0.02fF
C12568 NAND2X1_LOC_130/Y INVX1_LOC_519/Y 0.59fF
C12569 INVX1_LOC_463/Y NAND2X1_LOC_829/B 0.01fF
C12570 NAND2X1_LOC_181/A INVX1_LOC_32/Y 0.01fF
C12571 INVX1_LOC_116/A NAND2X1_LOC_604/a_36_24# 0.00fF
C12572 INVX1_LOC_266/A NAND2X1_LOC_544/B 0.05fF
C12573 INVX1_LOC_130/Y INVX1_LOC_100/Y 0.03fF
C12574 INVX1_LOC_500/Y INVX1_LOC_501/A 0.14fF
C12575 INVX1_LOC_145/Y INVX1_LOC_114/A 0.03fF
C12576 INVX1_LOC_79/A INVX1_LOC_7/Y 0.03fF
C12577 NAND2X1_LOC_123/a_36_24# INVX1_LOC_347/Y 0.00fF
C12578 INVX1_LOC_58/Y NAND2X1_LOC_267/A 0.08fF
C12579 INVX1_LOC_47/Y NAND2X1_LOC_695/a_36_24# 0.01fF
C12580 NAND2X1_LOC_631/B INVX1_LOC_7/Y 0.03fF
C12581 NAND2X1_LOC_274/B INVX1_LOC_137/Y 0.04fF
C12582 INVX1_LOC_31/Y INVX1_LOC_44/Y 0.09fF
C12583 INVX1_LOC_555/A INVX1_LOC_58/Y 0.00fF
C12584 INVX1_LOC_41/Y INVX1_LOC_1/Y 0.01fF
C12585 INVX1_LOC_379/A NAND2X1_LOC_528/Y 0.05fF
C12586 INVX1_LOC_207/Y GATE_222 0.04fF
C12587 INVX1_LOC_117/Y INVX1_LOC_26/Y 1.72fF
C12588 INVX1_LOC_345/Y INVX1_LOC_79/A 0.02fF
C12589 NAND2X1_LOC_27/Y INVX1_LOC_531/Y 0.00fF
C12590 INVX1_LOC_35/Y INVX1_LOC_479/A 0.10fF
C12591 INVX1_LOC_107/Y INVX1_LOC_58/Y 0.00fF
C12592 INVX1_LOC_32/Y INVX1_LOC_79/A 0.39fF
C12593 INVX1_LOC_209/A INVX1_LOC_274/Y 0.00fF
C12594 NAND2X1_LOC_790/B INVX1_LOC_275/A 0.02fF
C12595 NAND2X1_LOC_191/a_36_24# NAND2X1_LOC_123/B 0.01fF
C12596 INVX1_LOC_500/A INVX1_LOC_493/Y 0.05fF
C12597 INVX1_LOC_504/A INVX1_LOC_348/Y 0.02fF
C12598 INVX1_LOC_32/Y NAND2X1_LOC_396/Y 0.02fF
C12599 NAND2X1_LOC_689/B INVX1_LOC_41/Y 0.00fF
C12600 INVX1_LOC_110/A INVX1_LOC_74/Y 0.06fF
C12601 VDD INVX1_LOC_279/A -0.00fF
C12602 INVX1_LOC_31/Y INVX1_LOC_347/A 0.34fF
C12603 NAND2X1_LOC_93/Y NAND2X1_LOC_790/B 0.01fF
C12604 INVX1_LOC_520/Y NAND2X1_LOC_136/Y 0.00fF
C12605 INVX1_LOC_117/A INVX1_LOC_9/Y 0.01fF
C12606 INVX1_LOC_479/A NAND2X1_LOC_253/Y 0.02fF
C12607 NAND2X1_LOC_637/A INVX1_LOC_206/Y 0.01fF
C12608 NAND2X1_LOC_106/Y INVX1_LOC_109/A 0.23fF
C12609 INVX1_LOC_476/A INVX1_LOC_645/Y 0.00fF
C12610 INVX1_LOC_41/Y INVX1_LOC_245/A 0.06fF
C12611 INVX1_LOC_45/Y INVX1_LOC_638/A 0.01fF
C12612 INVX1_LOC_85/Y INVX1_LOC_616/Y 0.01fF
C12613 INVX1_LOC_446/Y NAND2X1_LOC_457/A 0.06fF
C12614 INVX1_LOC_442/A NAND2X1_LOC_332/a_36_24# 0.02fF
C12615 INVX1_LOC_118/Y INVX1_LOC_362/Y 0.00fF
C12616 INVX1_LOC_206/Y INVX1_LOC_586/A 0.11fF
C12617 NAND2X1_LOC_219/a_36_24# INVX1_LOC_366/A 0.01fF
C12618 INVX1_LOC_435/Y INVX1_LOC_428/A 0.05fF
C12619 VDD INVX1_LOC_668/A -0.00fF
C12620 INVX1_LOC_434/A INVX1_LOC_406/Y 0.06fF
C12621 VDD INVX1_LOC_318/Y 0.49fF
C12622 VDD INVX1_LOC_565/Y 0.21fF
C12623 INVX1_LOC_438/A INVX1_LOC_235/Y 0.06fF
C12624 NAND2X1_LOC_45/Y INVX1_LOC_84/A 0.03fF
C12625 INVX1_LOC_405/A INVX1_LOC_99/Y 0.03fF
C12626 VDD INVX1_LOC_455/Y 0.22fF
C12627 INVX1_LOC_224/Y INVX1_LOC_486/Y 0.03fF
C12628 INVX1_LOC_118/Y INVX1_LOC_683/Y 0.02fF
C12629 INVX1_LOC_312/Y INVX1_LOC_206/Y 0.03fF
C12630 VDD INVX1_LOC_16/Y 0.26fF
C12631 VDD INVX1_LOC_370/Y 0.51fF
C12632 INVX1_LOC_228/Y INVX1_LOC_318/Y 0.90fF
C12633 INVX1_LOC_396/Y INVX1_LOC_586/A 0.11fF
C12634 INVX1_LOC_20/Y INVX1_LOC_269/A 0.32fF
C12635 INVX1_LOC_450/A INVX1_LOC_424/Y 0.02fF
C12636 INVX1_LOC_393/Y INVX1_LOC_519/A 0.26fF
C12637 INVX1_LOC_346/Y INVX1_LOC_348/Y 0.01fF
C12638 INVX1_LOC_191/Y INVX1_LOC_7/Y 0.50fF
C12639 INVX1_LOC_398/A INVX1_LOC_45/Y 0.01fF
C12640 NAND2X1_LOC_231/A INVX1_LOC_286/Y 0.03fF
C12641 NAND2X1_LOC_391/A INVX1_LOC_395/A 0.03fF
C12642 INVX1_LOC_578/A INVX1_LOC_486/Y 0.02fF
C12643 VDD INVX1_LOC_668/Y 0.21fF
C12644 NAND2X1_LOC_332/a_36_24# INVX1_LOC_116/Y 0.00fF
C12645 INVX1_LOC_278/A NAND2X1_LOC_260/Y 0.27fF
C12646 INVX1_LOC_586/A INVX1_LOC_686/A 0.10fF
C12647 NAND2X1_LOC_457/A INVX1_LOC_145/Y 0.04fF
C12648 NAND2X1_LOC_416/B NAND2X1_LOC_415/a_36_24# 0.02fF
C12649 INVX1_LOC_450/A NAND2X1_LOC_559/a_36_24# 0.01fF
C12650 INVX1_LOC_139/A INVX1_LOC_491/Y 0.22fF
C12651 INVX1_LOC_395/A NAND2X1_LOC_418/Y 0.32fF
C12652 INVX1_LOC_442/A NAND2X1_LOC_603/Y 0.01fF
C12653 INVX1_LOC_206/Y NAND2X1_LOC_202/a_36_24# 0.00fF
C12654 NAND2X1_LOC_99/a_36_24# INVX1_LOC_525/Y 0.00fF
C12655 NAND2X1_LOC_249/Y INVX1_LOC_117/Y 0.07fF
C12656 INVX1_LOC_118/Y INVX1_LOC_548/A 0.00fF
C12657 INVX1_LOC_65/Y INVX1_LOC_600/A 0.08fF
C12658 INVX1_LOC_206/Y NAND2X1_LOC_74/a_36_24# 0.00fF
C12659 INVX1_LOC_545/A INVX1_LOC_412/A 0.28fF
C12660 INVX1_LOC_395/A INVX1_LOC_365/A 0.04fF
C12661 INPUT_0 INVX1_LOC_8/Y 0.09fF
C12662 INVX1_LOC_442/A NAND2X1_LOC_323/a_36_24# 0.00fF
C12663 INVX1_LOC_238/A INVX1_LOC_117/Y 0.04fF
C12664 INVX1_LOC_547/Y INVX1_LOC_145/Y 0.54fF
C12665 INVX1_LOC_65/Y INVX1_LOC_64/A 0.03fF
C12666 NAND2X1_LOC_176/Y INVX1_LOC_31/Y 0.01fF
C12667 INVX1_LOC_581/A NAND2X1_LOC_155/a_36_24# 0.00fF
C12668 INVX1_LOC_367/A INVX1_LOC_126/A 0.03fF
C12669 VDD INVX1_LOC_326/A 0.00fF
C12670 INVX1_LOC_300/A INVX1_LOC_269/A 0.04fF
C12671 INPUT_3 INVX1_LOC_10/Y 0.01fF
C12672 INVX1_LOC_451/A INVX1_LOC_45/Y 0.12fF
C12673 INVX1_LOC_50/Y INVX1_LOC_49/A 0.01fF
C12674 INVX1_LOC_577/A INVX1_LOC_32/Y 0.01fF
C12675 NAND2X1_LOC_637/A NAND2X1_LOC_334/A 0.05fF
C12676 INVX1_LOC_560/A INVX1_LOC_117/Y 0.08fF
C12677 INVX1_LOC_454/A INVX1_LOC_659/A 0.07fF
C12678 INVX1_LOC_241/Y INVX1_LOC_242/A 0.01fF
C12679 INVX1_LOC_463/A INVX1_LOC_501/A 0.01fF
C12680 INVX1_LOC_21/A INVX1_LOC_22/Y 0.00fF
C12681 INVX1_LOC_45/Y INVX1_LOC_665/Y 0.03fF
C12682 INVX1_LOC_68/Y INVX1_LOC_479/Y 0.01fF
C12683 INVX1_LOC_249/Y INVX1_LOC_578/Y 1.01fF
C12684 INVX1_LOC_395/A INVX1_LOC_523/Y 0.54fF
C12685 INVX1_LOC_84/A INVX1_LOC_99/Y 0.35fF
C12686 INVX1_LOC_287/A INVX1_LOC_250/Y 0.45fF
C12687 NAND2X1_LOC_147/B INVX1_LOC_131/A 0.02fF
C12688 INVX1_LOC_579/A NAND2X1_LOC_802/a_36_24# 0.00fF
C12689 INVX1_LOC_11/Y NAND2X1_LOC_391/B 0.01fF
C12690 INVX1_LOC_402/A INVX1_LOC_53/Y 0.00fF
C12691 INVX1_LOC_578/Y NAND2X1_LOC_122/Y 0.01fF
C12692 INPUT_3 INVX1_LOC_451/A 2.87fF
C12693 INVX1_LOC_250/A INVX1_LOC_559/Y 0.10fF
C12694 INVX1_LOC_145/Y INVX1_LOC_651/A 0.00fF
C12695 NAND2X1_LOC_336/B INVX1_LOC_545/A 0.03fF
C12696 INVX1_LOC_604/Y INVX1_LOC_600/A 0.14fF
C12697 INVX1_LOC_425/A INVX1_LOC_93/Y 0.09fF
C12698 VDD INVX1_LOC_90/Y 2.42fF
C12699 INVX1_LOC_116/Y NAND2X1_LOC_603/Y 0.01fF
C12700 NAND2X1_LOC_779/a_36_24# INVX1_LOC_581/A -0.02fF
C12701 INPUT_0 INVX1_LOC_9/Y 1.18fF
C12702 NAND2X1_LOC_122/Y INVX1_LOC_532/Y 0.01fF
C12703 INVX1_LOC_12/Y INVX1_LOC_35/Y 0.18fF
C12704 INVX1_LOC_577/Y INVX1_LOC_157/A 0.02fF
C12705 INVX1_LOC_93/Y INVX1_LOC_126/A 0.01fF
C12706 INVX1_LOC_12/Y INVX1_LOC_304/A 1.03fF
C12707 NAND2X1_LOC_323/a_36_24# INVX1_LOC_116/Y 0.01fF
C12708 INVX1_LOC_355/A INVX1_LOC_501/A 0.03fF
C12709 INVX1_LOC_105/A INVX1_LOC_134/Y 0.02fF
C12710 INVX1_LOC_99/Y NAND2X1_LOC_67/Y 0.01fF
C12711 NAND2X1_LOC_260/Y INVX1_LOC_453/Y 0.25fF
C12712 NAND2X1_LOC_413/Y INVX1_LOC_98/Y 0.04fF
C12713 INVX1_LOC_84/A INVX1_LOC_123/A 0.03fF
C12714 INVX1_LOC_202/Y INVX1_LOC_155/Y 0.30fF
C12715 NAND2X1_LOC_108/Y NAND2X1_LOC_108/a_36_24# 0.02fF
C12716 INVX1_LOC_361/Y INVX1_LOC_519/A 0.06fF
C12717 INVX1_LOC_468/Y INVX1_LOC_252/A 0.00fF
C12718 INVX1_LOC_418/Y INVX1_LOC_99/A 0.06fF
C12719 INVX1_LOC_586/A NAND2X1_LOC_334/A 0.01fF
C12720 INVX1_LOC_117/Y INVX1_LOC_369/A 0.03fF
C12721 INVX1_LOC_51/Y INVX1_LOC_44/Y 0.07fF
C12722 INVX1_LOC_228/Y INVX1_LOC_90/Y 0.07fF
C12723 INVX1_LOC_99/A INVX1_LOC_159/Y 0.01fF
C12724 INVX1_LOC_80/A INVX1_LOC_670/A 0.03fF
C12725 INPUT_0 INVX1_LOC_166/Y 0.03fF
C12726 INVX1_LOC_160/Y INVX1_LOC_245/A 0.01fF
C12727 INVX1_LOC_586/A NAND2X1_LOC_452/a_36_24# 0.01fF
C12728 INVX1_LOC_53/Y INVX1_LOC_561/A 0.08fF
C12729 INVX1_LOC_84/A INVX1_LOC_47/Y 1.62fF
C12730 INVX1_LOC_7/Y INVX1_LOC_48/Y 0.07fF
C12731 NAND2X1_LOC_827/Y INVX1_LOC_59/A 0.01fF
C12732 INVX1_LOC_32/Y INVX1_LOC_632/A 0.07fF
C12733 INVX1_LOC_84/A NAND2X1_LOC_557/B 0.12fF
C12734 INVX1_LOC_318/A INVX1_LOC_600/A 0.03fF
C12735 INPUT_0 INVX1_LOC_62/Y 0.16fF
C12736 INVX1_LOC_370/Y INVX1_LOC_103/Y 0.01fF
C12737 INVX1_LOC_358/Y NAND2X1_LOC_689/B 0.02fF
C12738 NAND2X1_LOC_710/A INVX1_LOC_49/Y 0.01fF
C12739 INVX1_LOC_579/A INVX1_LOC_261/Y 0.01fF
C12740 NAND2X1_LOC_41/Y INVX1_LOC_171/A 0.09fF
C12741 INVX1_LOC_614/A INVX1_LOC_476/A 0.03fF
C12742 INVX1_LOC_304/Y INVX1_LOC_681/Y 0.02fF
C12743 INVX1_LOC_31/Y NAND2X1_LOC_418/Y 0.22fF
C12744 INVX1_LOC_49/Y NAND2X1_LOC_541/B 0.29fF
C12745 INVX1_LOC_366/A NAND2X1_LOC_699/a_36_24# 0.01fF
C12746 INVX1_LOC_398/Y INVX1_LOC_32/Y 0.01fF
C12747 INVX1_LOC_490/A NAND2X1_LOC_416/Y 0.04fF
C12748 INVX1_LOC_93/Y INVX1_LOC_252/Y 0.07fF
C12749 NAND2X1_LOC_782/A INVX1_LOC_137/Y 0.02fF
C12750 INVX1_LOC_35/Y INVX1_LOC_138/Y 0.01fF
C12751 NAND2X1_LOC_56/Y NAND2X1_LOC_52/Y 0.30fF
C12752 INVX1_LOC_32/Y INVX1_LOC_59/Y 0.15fF
C12753 INVX1_LOC_566/A NAND2X1_LOC_405/a_36_24# 0.00fF
C12754 INVX1_LOC_17/Y INVX1_LOC_671/Y 0.13fF
C12755 INVX1_LOC_596/A NAND2X1_LOC_768/B 0.03fF
C12756 INVX1_LOC_49/Y INVX1_LOC_383/Y 0.05fF
C12757 INVX1_LOC_11/Y INVX1_LOC_670/A 0.01fF
C12758 INVX1_LOC_47/Y NAND2X1_LOC_67/Y 0.02fF
C12759 INVX1_LOC_51/Y INVX1_LOC_347/A 0.16fF
C12760 NAND2X1_LOC_413/Y INVX1_LOC_338/Y 0.21fF
C12761 NAND2X1_LOC_444/A INPUT_1 0.29fF
C12762 INVX1_LOC_32/Y INVX1_LOC_48/Y 3.37fF
C12763 INVX1_LOC_25/Y NAND2X1_LOC_836/B 0.43fF
C12764 INVX1_LOC_17/Y INVX1_LOC_77/Y 0.13fF
C12765 NAND2X1_LOC_148/A INVX1_LOC_662/A 0.05fF
C12766 INVX1_LOC_84/A NAND2X1_LOC_66/Y 1.39fF
C12767 NAND2X1_LOC_307/A NAND2X1_LOC_274/B 0.03fF
C12768 INVX1_LOC_545/Y NAND2X1_LOC_274/B 0.00fF
C12769 INVX1_LOC_183/A NAND2X1_LOC_671/a_36_24# 0.00fF
C12770 INVX1_LOC_68/Y NAND2X1_LOC_94/a_36_24# 0.00fF
C12771 INVX1_LOC_261/A INVX1_LOC_659/Y 0.01fF
C12772 INVX1_LOC_170/A INVX1_LOC_35/Y 0.00fF
C12773 INVX1_LOC_21/Y INVX1_LOC_245/A 0.36fF
C12774 INPUT_0 NAND2X1_LOC_269/a_36_24# 0.01fF
C12775 INVX1_LOC_598/A INVX1_LOC_204/Y 0.00fF
C12776 NAND2X1_LOC_791/B INVX1_LOC_621/A 0.02fF
C12777 INVX1_LOC_607/Y INVX1_LOC_9/Y 0.09fF
C12778 NAND2X1_LOC_467/A NAND2X1_LOC_689/a_36_24# 0.00fF
C12779 INVX1_LOC_366/A NAND2X1_LOC_85/a_36_24# 0.00fF
C12780 INVX1_LOC_26/Y INVX1_LOC_281/Y 0.05fF
C12781 NAND2X1_LOC_586/Y INVX1_LOC_50/Y 0.02fF
C12782 INVX1_LOC_117/A INVX1_LOC_42/Y 0.01fF
C12783 NAND2X1_LOC_299/Y INVX1_LOC_74/Y 0.03fF
C12784 INVX1_LOC_26/Y INVX1_LOC_178/A 0.32fF
C12785 NAND2X1_LOC_91/a_36_24# NAND2X1_LOC_267/A 0.01fF
C12786 NAND2X1_LOC_167/a_36_24# INPUT_1 0.00fF
C12787 NAND2X1_LOC_66/Y NAND2X1_LOC_67/Y 0.00fF
C12788 NAND2X1_LOC_274/B NAND2X1_LOC_600/a_36_24# 0.00fF
C12789 INVX1_LOC_242/Y INVX1_LOC_259/Y 0.11fF
C12790 INVX1_LOC_69/Y NAND2X1_LOC_542/A 0.02fF
C12791 NAND2X1_LOC_147/B NAND2X1_LOC_843/B 0.02fF
C12792 NAND2X1_LOC_267/A INVX1_LOC_245/A 0.02fF
C12793 INVX1_LOC_261/Y INVX1_LOC_659/A 0.03fF
C12794 INVX1_LOC_573/Y INVX1_LOC_331/Y 0.01fF
C12795 INPUT_5 INVX1_LOC_340/A 0.01fF
C12796 INVX1_LOC_294/A INVX1_LOC_369/Y 0.01fF
C12797 INVX1_LOC_608/A INVX1_LOC_26/Y 0.45fF
C12798 INVX1_LOC_54/Y NAND2X1_LOC_301/B 0.01fF
C12799 INVX1_LOC_83/A INVX1_LOC_9/Y 0.01fF
C12800 INVX1_LOC_110/A INVX1_LOC_79/A 0.07fF
C12801 NAND2X1_LOC_184/Y INVX1_LOC_100/Y 0.92fF
C12802 INVX1_LOC_214/Y INVX1_LOC_479/A 0.00fF
C12803 NAND2X1_LOC_27/Y INVX1_LOC_41/Y 0.02fF
C12804 INVX1_LOC_69/Y INVX1_LOC_376/Y 0.07fF
C12805 INVX1_LOC_643/Y NAND2X1_LOC_814/Y 0.00fF
C12806 INVX1_LOC_644/Y INVX1_LOC_6/Y 0.01fF
C12807 INVX1_LOC_157/A INVX1_LOC_26/Y 0.01fF
C12808 INVX1_LOC_179/A NAND2X1_LOC_455/a_36_24# 0.01fF
C12809 INVX1_LOC_298/A INVX1_LOC_62/Y 0.03fF
C12810 INVX1_LOC_479/A INVX1_LOC_118/A 0.01fF
C12811 INVX1_LOC_35/Y INVX1_LOC_212/A 0.04fF
C12812 INVX1_LOC_58/Y INVX1_LOC_26/Y 0.04fF
C12813 INVX1_LOC_166/A INVX1_LOC_652/Y 0.00fF
C12814 INVX1_LOC_298/A INVX1_LOC_529/Y 0.01fF
C12815 INVX1_LOC_551/A INVX1_LOC_100/Y 0.03fF
C12816 INVX1_LOC_551/A INVX1_LOC_74/Y 0.03fF
C12817 INVX1_LOC_647/Y INVX1_LOC_212/Y 0.01fF
C12818 INVX1_LOC_366/A NAND2X1_LOC_86/Y 0.02fF
C12819 NAND2X1_LOC_274/B NAND2X1_LOC_602/a_36_24# 0.00fF
C12820 INVX1_LOC_206/Y INVX1_LOC_140/Y 0.03fF
C12821 INVX1_LOC_100/Y INVX1_LOC_75/Y 0.15fF
C12822 NAND2X1_LOC_310/a_36_24# INVX1_LOC_269/A 0.01fF
C12823 NAND2X1_LOC_704/a_36_24# INVX1_LOC_546/A 0.02fF
C12824 INVX1_LOC_118/Y INVX1_LOC_51/Y 0.07fF
C12825 INVX1_LOC_426/A NAND2X1_LOC_391/A 0.01fF
C12826 INVX1_LOC_266/A NAND2X1_LOC_176/Y 0.03fF
C12827 INVX1_LOC_206/Y NAND2X1_LOC_426/Y 0.01fF
C12828 INVX1_LOC_62/Y INVX1_LOC_211/A 0.02fF
C12829 VDD NAND2X1_LOC_523/B 0.01fF
C12830 INVX1_LOC_84/A NAND2X1_LOC_475/A 0.04fF
C12831 INVX1_LOC_425/A INVX1_LOC_395/A 0.67fF
C12832 VDD NAND2X1_LOC_545/B 0.04fF
C12833 INVX1_LOC_206/Y NAND2X1_LOC_791/B 0.03fF
C12834 INVX1_LOC_206/Y INVX1_LOC_272/Y 0.02fF
C12835 INVX1_LOC_206/Y INVX1_LOC_294/Y 0.05fF
C12836 INVX1_LOC_405/A NAND2X1_LOC_276/a_36_24# 0.00fF
C12837 NAND2X1_LOC_330/a_36_24# INVX1_LOC_495/A 0.00fF
C12838 INVX1_LOC_586/A INVX1_LOC_94/A 0.24fF
C12839 INVX1_LOC_20/Y NAND2X1_LOC_337/a_36_24# 0.00fF
C12840 INVX1_LOC_38/A NAND2X1_LOC_29/a_36_24# 0.00fF
C12841 NAND2X1_LOC_750/Y NAND2X1_LOC_318/B 0.02fF
C12842 NAND2X1_LOC_562/a_36_24# INVX1_LOC_384/Y 0.01fF
C12843 INVX1_LOC_490/Y INVX1_LOC_53/Y 0.03fF
C12844 INVX1_LOC_648/Y NAND2X1_LOC_820/A 0.19fF
C12845 INVX1_LOC_103/A INVX1_LOC_104/Y 0.00fF
C12846 VDD INVX1_LOC_98/Y 2.74fF
C12847 INVX1_LOC_145/A NAND2X1_LOC_31/a_36_24# 0.00fF
C12848 NAND2X1_LOC_537/A INVX1_LOC_194/Y 0.05fF
C12849 NAND2X1_LOC_16/Y INVX1_LOC_53/Y 0.38fF
C12850 INVX1_LOC_6/Y NAND2X1_LOC_86/Y 0.01fF
C12851 INVX1_LOC_45/Y INVX1_LOC_134/Y 0.16fF
C12852 INVX1_LOC_72/Y INVX1_LOC_307/A 0.06fF
C12853 INVX1_LOC_76/Y INVX1_LOC_508/Y 0.02fF
C12854 INVX1_LOC_182/A INVX1_LOC_21/Y 0.01fF
C12855 INVX1_LOC_412/Y NAND2X1_LOC_775/B 0.19fF
C12856 NAND2X1_LOC_533/a_36_24# INVX1_LOC_31/Y 0.00fF
C12857 NAND2X1_LOC_377/a_36_24# INVX1_LOC_178/A 0.00fF
C12858 INVX1_LOC_47/A INVX1_LOC_45/Y 0.01fF
C12859 INVX1_LOC_316/Y INVX1_LOC_45/Y 0.14fF
C12860 INVX1_LOC_435/Y NAND2X1_LOC_521/a_36_24# 0.06fF
C12861 NAND2X1_LOC_41/Y INVX1_LOC_45/Y 0.01fF
C12862 INVX1_LOC_409/Y INVX1_LOC_63/Y 0.06fF
C12863 INVX1_LOC_533/Y INVX1_LOC_259/Y 0.07fF
C12864 INVX1_LOC_594/Y INVX1_LOC_69/Y 0.03fF
C12865 INVX1_LOC_510/Y INVX1_LOC_98/Y 0.10fF
C12866 NAND2X1_LOC_249/Y INVX1_LOC_58/Y 0.16fF
C12867 VDD INVX1_LOC_497/A -0.00fF
C12868 INVX1_LOC_432/Y NAND2X1_LOC_391/B 0.01fF
C12869 INVX1_LOC_206/Y INVX1_LOC_6/Y 1.31fF
C12870 VDD INVX1_LOC_338/Y 1.46fF
C12871 NAND2X1_LOC_335/B INVX1_LOC_63/Y 0.01fF
C12872 INPUT_7 INVX1_LOC_69/A 0.38fF
C12873 NAND2X1_LOC_148/B NAND2X1_LOC_142/Y 0.00fF
C12874 INVX1_LOC_384/A INVX1_LOC_303/Y 0.05fF
C12875 NAND2X1_LOC_165/Y INVX1_LOC_45/Y 0.02fF
C12876 NAND2X1_LOC_13/Y INVX1_LOC_194/Y 0.01fF
C12877 NAND2X1_LOC_97/A NAND2X1_LOC_333/B 0.03fF
C12878 INVX1_LOC_20/Y INVX1_LOC_259/Y 0.03fF
C12879 NAND2X1_LOC_44/a_36_24# INVX1_LOC_93/A 0.00fF
C12880 INVX1_LOC_442/Y INVX1_LOC_519/A 0.03fF
C12881 INVX1_LOC_435/A NAND2X1_LOC_528/a_36_24# 0.00fF
C12882 INVX1_LOC_417/Y INVX1_LOC_130/Y 0.32fF
C12883 INVX1_LOC_596/A NAND2X1_LOC_464/a_36_24# 0.01fF
C12884 INVX1_LOC_54/Y INVX1_LOC_551/Y 1.73fF
C12885 NAND2X1_LOC_516/a_36_24# INVX1_LOC_6/Y 0.01fF
C12886 INVX1_LOC_435/A INVX1_LOC_80/A 0.02fF
C12887 INVX1_LOC_293/Y INVX1_LOC_665/Y 0.03fF
C12888 INVX1_LOC_369/A INVX1_LOC_178/A 0.07fF
C12889 NAND2X1_LOC_142/Y INVX1_LOC_69/Y 0.04fF
C12890 NAND2X1_LOC_535/a_36_24# NAND2X1_LOC_274/B 0.00fF
C12891 INVX1_LOC_117/Y INVX1_LOC_235/Y 0.23fF
C12892 NAND2X1_LOC_759/a_36_24# INVX1_LOC_53/Y 0.00fF
C12893 INVX1_LOC_584/Y INVX1_LOC_168/Y 0.04fF
C12894 INVX1_LOC_20/Y NAND2X1_LOC_707/B 0.01fF
C12895 INVX1_LOC_586/A NAND2X1_LOC_542/A 0.00fF
C12896 INVX1_LOC_6/Y INVX1_LOC_242/A 0.03fF
C12897 INVX1_LOC_586/Y INVX1_LOC_87/A 0.01fF
C12898 INVX1_LOC_625/A NAND2X1_LOC_795/a_36_24# 0.02fF
C12899 INVX1_LOC_578/A NAND2X1_LOC_861/a_36_24# 0.00fF
C12900 INVX1_LOC_579/A INVX1_LOC_578/Y 0.02fF
C12901 INVX1_LOC_68/Y INVX1_LOC_63/Y 0.04fF
C12902 NAND2X1_LOC_88/B INVX1_LOC_87/Y 0.01fF
C12903 INVX1_LOC_166/A INVX1_LOC_197/A 0.03fF
C12904 INVX1_LOC_551/Y INVX1_LOC_257/A 0.10fF
C12905 INVX1_LOC_469/Y NAND2X1_LOC_299/Y 0.00fF
C12906 INVX1_LOC_20/Y INVX1_LOC_204/Y 0.05fF
C12907 INVX1_LOC_21/Y NAND2X1_LOC_27/Y 0.00fF
C12908 NAND2X1_LOC_45/a_36_24# INVX1_LOC_62/Y 0.01fF
C12909 INVX1_LOC_586/A INVX1_LOC_376/Y 0.10fF
C12910 INVX1_LOC_53/Y INVX1_LOC_18/Y 0.03fF
C12911 INVX1_LOC_257/Y INVX1_LOC_62/Y 0.07fF
C12912 INVX1_LOC_435/A INVX1_LOC_11/Y 0.02fF
C12913 INVX1_LOC_85/Y INVX1_LOC_543/A 0.01fF
C12914 INVX1_LOC_156/A INVX1_LOC_99/Y 0.15fF
C12915 INVX1_LOC_577/Y INVX1_LOC_245/A 0.03fF
C12916 INVX1_LOC_384/A INVX1_LOC_9/Y 0.07fF
C12917 INVX1_LOC_418/Y INVX1_LOC_419/Y 0.01fF
C12918 INVX1_LOC_587/Y INVX1_LOC_145/Y 0.03fF
C12919 NAND2X1_LOC_822/Y INVX1_LOC_99/Y 0.01fF
C12920 INVX1_LOC_607/A INVX1_LOC_100/Y 0.28fF
C12921 INVX1_LOC_416/A INVX1_LOC_159/Y 0.01fF
C12922 INVX1_LOC_35/Y NAND2X1_LOC_615/B 0.03fF
C12923 INVX1_LOC_93/Y NAND2X1_LOC_156/Y 0.15fF
C12924 INVX1_LOC_609/Y INVX1_LOC_6/Y 0.01fF
C12925 INVX1_LOC_140/Y NAND2X1_LOC_609/B 0.00fF
C12926 INVX1_LOC_419/Y INVX1_LOC_159/Y 0.02fF
C12927 INVX1_LOC_556/Y INVX1_LOC_117/Y 0.19fF
C12928 INVX1_LOC_369/A INVX1_LOC_58/Y 0.03fF
C12929 INVX1_LOC_31/Y INVX1_LOC_252/Y 0.03fF
C12930 INVX1_LOC_588/Y NAND2X1_LOC_174/B 0.03fF
C12931 INVX1_LOC_17/Y INVX1_LOC_372/A 0.01fF
C12932 NAND2X1_LOC_532/Y INVX1_LOC_99/Y 0.03fF
C12933 INVX1_LOC_288/A INVX1_LOC_62/Y 0.07fF
C12934 INVX1_LOC_20/Y INVX1_LOC_114/A 0.03fF
C12935 INVX1_LOC_261/A INVX1_LOC_55/Y 0.03fF
C12936 INVX1_LOC_63/Y INVX1_LOC_600/A 0.02fF
C12937 NAND2X1_LOC_285/B INVX1_LOC_239/A 0.14fF
C12938 INVX1_LOC_35/Y INVX1_LOC_66/A 0.68fF
C12939 NAND2X1_LOC_147/a_36_24# INVX1_LOC_662/A 0.01fF
C12940 INVX1_LOC_396/A INVX1_LOC_32/Y 0.01fF
C12941 INVX1_LOC_452/A INVX1_LOC_6/Y 0.56fF
C12942 INPUT_0 NAND2X1_LOC_224/a_36_24# 0.01fF
C12943 INVX1_LOC_63/Y INVX1_LOC_64/A 0.01fF
C12944 INVX1_LOC_9/A INVX1_LOC_9/Y 0.00fF
C12945 INVX1_LOC_17/Y NAND2X1_LOC_537/a_36_24# 0.00fF
C12946 INVX1_LOC_384/A INVX1_LOC_62/Y 0.08fF
C12947 INVX1_LOC_448/A INVX1_LOC_9/Y 0.07fF
C12948 INVX1_LOC_213/Y NAND2X1_LOC_258/Y 0.01fF
C12949 INVX1_LOC_85/Y INVX1_LOC_86/A 0.06fF
C12950 INVX1_LOC_384/A NAND2X1_LOC_844/A 0.04fF
C12951 INVX1_LOC_47/Y INVX1_LOC_156/A 0.04fF
C12952 INVX1_LOC_145/Y INVX1_LOC_9/Y 0.07fF
C12953 NAND2X1_LOC_184/Y NAND2X1_LOC_181/A 0.00fF
C12954 INVX1_LOC_58/Y INVX1_LOC_603/A 0.03fF
C12955 INVX1_LOC_444/Y INVX1_LOC_245/A 0.03fF
C12956 NAND2X1_LOC_274/B INVX1_LOC_503/A 0.01fF
C12957 INVX1_LOC_545/Y INVX1_LOC_468/A 0.00fF
C12958 INVX1_LOC_419/A INVX1_LOC_93/Y 0.03fF
C12959 INVX1_LOC_340/A NAND2X1_LOC_425/a_36_24# 0.02fF
C12960 INVX1_LOC_93/Y INVX1_LOC_234/Y 0.10fF
C12961 INVX1_LOC_17/Y NAND2X1_LOC_274/B 0.03fF
C12962 INVX1_LOC_194/A INVX1_LOC_242/Y 0.01fF
C12963 INVX1_LOC_168/Y INVX1_LOC_186/Y 0.04fF
C12964 INVX1_LOC_26/Y INVX1_LOC_1/Y 0.02fF
C12965 INVX1_LOC_183/A INVX1_LOC_50/Y 0.14fF
C12966 NAND2X1_LOC_145/a_36_24# NAND2X1_LOC_843/B 0.00fF
C12967 INVX1_LOC_255/A NAND2X1_LOC_443/a_36_24# 0.01fF
C12968 INVX1_LOC_212/Y NAND2X1_LOC_342/A 0.21fF
C12969 INVX1_LOC_501/A INVX1_LOC_359/A 0.07fF
C12970 NAND2X1_LOC_334/A INVX1_LOC_6/Y 0.02fF
C12971 INVX1_LOC_502/A INVX1_LOC_159/Y 0.07fF
C12972 INVX1_LOC_62/Y INVX1_LOC_145/Y 5.89fF
C12973 NAND2X1_LOC_84/B INVX1_LOC_85/A 0.10fF
C12974 NAND2X1_LOC_133/a_36_24# INVX1_LOC_9/Y 0.00fF
C12975 INVX1_LOC_145/Y NAND2X1_LOC_844/A 0.01fF
C12976 INVX1_LOC_99/Y NAND2X1_LOC_497/a_36_24# 0.01fF
C12977 INVX1_LOC_501/A NAND2X1_LOC_449/B 0.04fF
C12978 INVX1_LOC_603/Y INVX1_LOC_270/Y 0.02fF
C12979 INVX1_LOC_93/Y INVX1_LOC_665/A 0.09fF
C12980 INVX1_LOC_89/Y NAND2X1_LOC_301/B 0.07fF
C12981 INVX1_LOC_543/Y INVX1_LOC_41/Y 0.00fF
C12982 INVX1_LOC_518/Y INVX1_LOC_66/A 0.01fF
C12983 INVX1_LOC_173/Y INVX1_LOC_531/Y 0.02fF
C12984 INVX1_LOC_154/A NAND2X1_LOC_301/B 0.00fF
C12985 INVX1_LOC_603/Y INVX1_LOC_92/A 0.09fF
C12986 INVX1_LOC_58/Y INVX1_LOC_632/Y 0.03fF
C12987 NAND2X1_LOC_691/A INVX1_LOC_496/Y 0.01fF
C12988 INVX1_LOC_435/A INVX1_LOC_231/Y 0.05fF
C12989 INVX1_LOC_54/Y INVX1_LOC_634/Y 0.01fF
C12990 INVX1_LOC_26/Y INVX1_LOC_245/A 0.06fF
C12991 INVX1_LOC_382/A NAND2X1_LOC_416/B 0.03fF
C12992 NAND2X1_LOC_686/B INVX1_LOC_479/A 0.01fF
C12993 INVX1_LOC_405/Y INVX1_LOC_502/A 0.00fF
C12994 INVX1_LOC_405/A NAND2X1_LOC_520/B 0.11fF
C12995 NAND2X1_LOC_123/B INVX1_LOC_491/A 0.23fF
C12996 INVX1_LOC_89/Y INVX1_LOC_291/Y 0.01fF
C12997 INVX1_LOC_662/A INVX1_LOC_653/Y 0.03fF
C12998 INVX1_LOC_409/Y INVX1_LOC_374/A 0.00fF
C12999 INVX1_LOC_435/Y VDD 3.23fF
C13000 INVX1_LOC_425/A INVX1_LOC_426/A 0.02fF
C13001 INPUT_0 NAND2X1_LOC_331/A 0.03fF
C13002 INVX1_LOC_239/Y INVX1_LOC_133/A 0.00fF
C13003 INVX1_LOC_79/A INVX1_LOC_75/Y 0.04fF
C13004 INVX1_LOC_118/Y INVX1_LOC_216/Y 0.01fF
C13005 INVX1_LOC_594/Y INVX1_LOC_586/A 0.03fF
C13006 INVX1_LOC_230/A INVX1_LOC_109/Y 0.02fF
C13007 INVX1_LOC_488/A INVX1_LOC_488/Y 0.01fF
C13008 NAND2X1_LOC_110/a_36_24# INVX1_LOC_45/Y 0.00fF
C13009 INVX1_LOC_224/Y INVX1_LOC_381/A 0.02fF
C13010 VDD INVX1_LOC_596/A 0.37fF
C13011 INVX1_LOC_79/A NAND2X1_LOC_271/A 0.03fF
C13012 NAND2X1_LOC_69/B INVX1_LOC_7/Y 0.03fF
C13013 INVX1_LOC_1/A INVX1_LOC_4/Y 0.01fF
C13014 INVX1_LOC_425/A NAND2X1_LOC_539/a_36_24# 0.00fF
C13015 INVX1_LOC_271/Y INVX1_LOC_286/A 0.14fF
C13016 INVX1_LOC_54/A INVX1_LOC_53/Y 0.03fF
C13017 VDD NAND2X1_LOC_318/B 0.05fF
C13018 INVX1_LOC_224/Y INVX1_LOC_320/A 0.02fF
C13019 INVX1_LOC_412/Y INVX1_LOC_633/Y 0.00fF
C13020 VDD INVX1_LOC_366/Y 0.22fF
C13021 VDD INVX1_LOC_504/A 0.00fF
C13022 INVX1_LOC_218/A INVX1_LOC_384/A 0.16fF
C13023 INVX1_LOC_51/Y INVX1_LOC_126/A 0.01fF
C13024 INVX1_LOC_32/A INVX1_LOC_176/A 0.03fF
C13025 INVX1_LOC_228/Y NAND2X1_LOC_318/B 0.88fF
C13026 INVX1_LOC_425/A INVX1_LOC_266/A 0.03fF
C13027 INVX1_LOC_552/Y INVX1_LOC_600/A -0.01fF
C13028 INVX1_LOC_20/Y INVX1_LOC_482/A 0.00fF
C13029 INVX1_LOC_300/A NAND2X1_LOC_719/a_36_24# 0.00fF
C13030 INVX1_LOC_584/A INVX1_LOC_537/A 0.01fF
C13031 INVX1_LOC_552/Y INVX1_LOC_64/A 0.04fF
C13032 INVX1_LOC_438/A INVX1_LOC_304/Y 0.03fF
C13033 INVX1_LOC_620/Y INVX1_LOC_623/A 0.00fF
C13034 INVX1_LOC_455/Y INVX1_LOC_45/Y 0.07fF
C13035 INVX1_LOC_222/Y INVX1_LOC_671/Y 0.02fF
C13036 NAND2X1_LOC_176/a_36_24# INVX1_LOC_270/A 0.01fF
C13037 INVX1_LOC_317/Y INVX1_LOC_417/A 0.01fF
C13038 INVX1_LOC_288/A INVX1_LOC_344/A 0.13fF
C13039 INVX1_LOC_20/Y INVX1_LOC_651/A 0.01fF
C13040 NAND2X1_LOC_790/B INVX1_LOC_58/Y 0.04fF
C13041 INVX1_LOC_442/A INVX1_LOC_35/Y 0.03fF
C13042 INVX1_LOC_558/A NAND2X1_LOC_461/a_36_24# 0.01fF
C13043 INVX1_LOC_428/Y INVX1_LOC_413/Y 0.13fF
C13044 INVX1_LOC_80/A INVX1_LOC_524/Y 0.15fF
C13045 INVX1_LOC_293/Y INVX1_LOC_134/Y 0.07fF
C13046 INVX1_LOC_671/A INVX1_LOC_445/A 0.08fF
C13047 INVX1_LOC_312/Y INVX1_LOC_295/A 0.13fF
C13048 INVX1_LOC_442/A INVX1_LOC_304/A 0.04fF
C13049 INVX1_LOC_51/Y INVX1_LOC_252/Y 0.20fF
C13050 INVX1_LOC_80/A INVX1_LOC_367/A 0.07fF
C13051 INVX1_LOC_218/A INVX1_LOC_145/Y 0.00fF
C13052 INVX1_LOC_55/Y INVX1_LOC_69/A 0.01fF
C13053 NAND2X1_LOC_241/B INVX1_LOC_208/Y 0.18fF
C13054 INVX1_LOC_193/Y INVX1_LOC_46/Y 0.01fF
C13055 INVX1_LOC_547/A INVX1_LOC_145/Y 0.11fF
C13056 INVX1_LOC_413/Y INVX1_LOC_50/Y 0.10fF
C13057 INVX1_LOC_605/A INVX1_LOC_46/Y 0.01fF
C13058 INVX1_LOC_20/Y INVX1_LOC_194/A 0.03fF
C13059 INVX1_LOC_257/Y INVX1_LOC_624/Y 0.01fF
C13060 NAND2X1_LOC_595/a_36_24# INVX1_LOC_9/Y 0.00fF
C13061 INVX1_LOC_112/Y INVX1_LOC_638/A 0.05fF
C13062 NAND2X1_LOC_352/a_36_24# NAND2X1_LOC_267/A 0.00fF
C13063 INVX1_LOC_139/A INVX1_LOC_149/Y 0.09fF
C13064 INVX1_LOC_560/Y INVX1_LOC_353/A 0.09fF
C13065 INVX1_LOC_80/A INVX1_LOC_669/Y 0.03fF
C13066 NAND2X1_LOC_180/B INPUT_1 0.01fF
C13067 INVX1_LOC_11/Y INVX1_LOC_367/A 0.07fF
C13068 INVX1_LOC_185/Y INVX1_LOC_476/A 0.00fF
C13069 NAND2X1_LOC_526/Y INVX1_LOC_69/Y 0.08fF
C13070 INVX1_LOC_418/A INVX1_LOC_257/A 0.03fF
C13071 INVX1_LOC_400/A INVX1_LOC_80/A 0.02fF
C13072 INVX1_LOC_54/Y INVX1_LOC_270/A 0.13fF
C13073 NAND2X1_LOC_756/Y NAND2X1_LOC_165/Y 0.04fF
C13074 INVX1_LOC_344/Y INVX1_LOC_99/Y 0.08fF
C13075 INVX1_LOC_21/Y INVX1_LOC_201/Y 0.01fF
C13076 INVX1_LOC_268/A INVX1_LOC_35/Y 0.01fF
C13077 INVX1_LOC_224/Y INVX1_LOC_100/Y 0.14fF
C13078 INVX1_LOC_596/A INVX1_LOC_103/Y 0.03fF
C13079 INVX1_LOC_554/Y INVX1_LOC_655/A 0.04fF
C13080 INVX1_LOC_586/A INVX1_LOC_139/Y 0.01fF
C13081 INVX1_LOC_551/Y INVX1_LOC_89/Y 0.01fF
C13082 INVX1_LOC_664/Y INVX1_LOC_445/A 0.01fF
C13083 INPUT_3 INVX1_LOC_326/A 0.01fF
C13084 INVX1_LOC_564/Y INVX1_LOC_245/A 0.02fF
C13085 INVX1_LOC_432/Y INVX1_LOC_435/A 0.00fF
C13086 INVX1_LOC_300/A INVX1_LOC_194/A 0.00fF
C13087 INVX1_LOC_35/Y INVX1_LOC_116/Y 0.12fF
C13088 INVX1_LOC_45/Y INVX1_LOC_351/A 0.01fF
C13089 INVX1_LOC_11/Y INVX1_LOC_516/A 0.00fF
C13090 INVX1_LOC_93/Y INVX1_LOC_80/A 0.29fF
C13091 INVX1_LOC_182/A INVX1_LOC_26/Y 0.02fF
C13092 INVX1_LOC_304/A INVX1_LOC_116/Y 0.03fF
C13093 INVX1_LOC_93/Y NAND2X1_LOC_768/A 0.02fF
C13094 NAND2X1_LOC_59/a_36_24# INVX1_LOC_204/Y 0.00fF
C13095 INVX1_LOC_330/A INVX1_LOC_332/Y 0.08fF
C13096 INVX1_LOC_578/A INVX1_LOC_100/Y 0.09fF
C13097 INVX1_LOC_17/Y INVX1_LOC_159/Y 0.12fF
C13098 INVX1_LOC_224/Y INVX1_LOC_74/Y 2.30fF
C13099 INVX1_LOC_21/Y INVX1_LOC_543/Y 0.03fF
C13100 INVX1_LOC_150/Y INVX1_LOC_500/A 0.01fF
C13101 NAND2X1_LOC_570/a_36_24# INVX1_LOC_452/A 0.01fF
C13102 INVX1_LOC_218/Y INVX1_LOC_444/Y 0.01fF
C13103 NAND2X1_LOC_332/B INVX1_LOC_9/Y 7.25fF
C13104 INVX1_LOC_11/Y INVX1_LOC_392/A 0.17fF
C13105 INVX1_LOC_18/Y INVX1_LOC_69/A 0.20fF
C13106 NAND2X1_LOC_117/a_36_24# NAND2X1_LOC_267/A 0.00fF
C13107 INVX1_LOC_449/A INVX1_LOC_406/A 0.03fF
C13108 VDD INVX1_LOC_346/Y 0.39fF
C13109 INVX1_LOC_45/Y INVX1_LOC_90/Y 0.08fF
C13110 INVX1_LOC_32/Y INVX1_LOC_155/Y 0.03fF
C13111 INVX1_LOC_511/A INVX1_LOC_498/Y 0.12fF
C13112 INVX1_LOC_145/Y INVX1_LOC_87/A 0.07fF
C13113 INVX1_LOC_320/A INVX1_LOC_120/Y 0.14fF
C13114 VDD NAND2X1_LOC_416/B 0.03fF
C13115 INVX1_LOC_199/Y NAND2X1_LOC_237/Y 0.03fF
C13116 INVX1_LOC_578/A INVX1_LOC_74/Y 0.17fF
C13117 INPUT_1 NAND2X1_LOC_444/a_36_24# 0.00fF
C13118 INVX1_LOC_11/Y INVX1_LOC_93/Y 0.84fF
C13119 INVX1_LOC_166/A INVX1_LOC_510/A 0.01fF
C13120 INVX1_LOC_452/A NAND2X1_LOC_294/Y 0.02fF
C13121 INVX1_LOC_522/A INVX1_LOC_514/A 0.00fF
C13122 NAND2X1_LOC_849/a_36_24# INVX1_LOC_510/A 0.00fF
C13123 NAND2X1_LOC_486/A NAND2X1_LOC_259/A 0.01fF
C13124 NAND2X1_LOC_184/Y INVX1_LOC_48/Y 0.16fF
C13125 INVX1_LOC_504/A INVX1_LOC_346/A 0.13fF
C13126 INPUT_3 INVX1_LOC_90/Y 0.48fF
C13127 INVX1_LOC_361/Y INVX1_LOC_670/A 0.23fF
C13128 INVX1_LOC_526/A INVX1_LOC_41/Y 0.01fF
C13129 INVX1_LOC_12/Y INVX1_LOC_223/Y 0.67fF
C13130 INVX1_LOC_54/Y NAND2X1_LOC_196/a_36_24# 0.01fF
C13131 INVX1_LOC_54/Y INVX1_LOC_46/Y 0.04fF
C13132 INVX1_LOC_651/A INVX1_LOC_655/A 0.06fF
C13133 INVX1_LOC_635/A INVX1_LOC_272/A 0.06fF
C13134 INVX1_LOC_206/Y INVX1_LOC_636/A 0.07fF
C13135 INVX1_LOC_176/A INVX1_LOC_49/Y 0.09fF
C13136 INVX1_LOC_551/A INVX1_LOC_59/Y 0.00fF
C13137 INVX1_LOC_556/Y INVX1_LOC_58/Y 0.02fF
C13138 INVX1_LOC_677/Y NAND2X1_LOC_451/B 0.03fF
C13139 NAND2X1_LOC_318/B NAND2X1_LOC_786/B 0.02fF
C13140 INVX1_LOC_376/Y INVX1_LOC_252/A 0.03fF
C13141 NAND2X1_LOC_635/B INVX1_LOC_69/Y 0.04fF
C13142 NAND2X1_LOC_387/Y INVX1_LOC_292/Y 0.06fF
C13143 INVX1_LOC_551/Y NAND2X1_LOC_544/B 0.03fF
C13144 NAND2X1_LOC_839/a_36_24# INVX1_LOC_59/A 0.00fF
C13145 INVX1_LOC_269/A INVX1_LOC_270/Y 0.00fF
C13146 INVX1_LOC_35/Y INVX1_LOC_179/A 0.03fF
C13147 INVX1_LOC_522/Y INVX1_LOC_479/A 0.14fF
C13148 INVX1_LOC_344/Y INVX1_LOC_119/Y 0.02fF
C13149 INVX1_LOC_197/A INVX1_LOC_41/Y 0.20fF
C13150 INVX1_LOC_220/Y INVX1_LOC_443/A 0.05fF
C13151 INVX1_LOC_376/A INVX1_LOC_345/A 0.06fF
C13152 NAND2X1_LOC_542/A INVX1_LOC_6/Y 0.41fF
C13153 INVX1_LOC_347/Y INVX1_LOC_355/Y 0.02fF
C13154 INVX1_LOC_177/A NAND2X1_LOC_786/B 0.02fF
C13155 INVX1_LOC_183/A INVX1_LOC_327/Y 0.01fF
C13156 INVX1_LOC_269/A INVX1_LOC_92/A 0.07fF
C13157 INVX1_LOC_387/Y INVX1_LOC_420/A 0.01fF
C13158 INVX1_LOC_245/A INVX1_LOC_603/A 0.00fF
C13159 INVX1_LOC_522/A INVX1_LOC_534/Y 0.01fF
C13160 INVX1_LOC_521/A INVX1_LOC_46/Y 0.01fF
C13161 INVX1_LOC_106/A NAND2X1_LOC_248/B 0.02fF
C13162 INVX1_LOC_21/Y INVX1_LOC_652/Y 0.01fF
C13163 NAND2X1_LOC_123/B INVX1_LOC_504/Y 0.08fF
C13164 INVX1_LOC_25/Y NAND2X1_LOC_409/Y 0.51fF
C13165 INVX1_LOC_417/Y INVX1_LOC_75/Y 0.81fF
C13166 INVX1_LOC_468/Y INVX1_LOC_74/Y 0.06fF
C13167 INVX1_LOC_93/Y NAND2X1_LOC_433/Y 0.07fF
C13168 INVX1_LOC_49/Y INVX1_LOC_420/A 0.01fF
C13169 INVX1_LOC_170/Y INVX1_LOC_49/Y 0.05fF
C13170 INVX1_LOC_17/Y NAND2X1_LOC_489/a_36_24# 0.00fF
C13171 INVX1_LOC_75/Y INVX1_LOC_59/Y 0.02fF
C13172 INVX1_LOC_79/A NAND2X1_LOC_469/a_36_24# 0.01fF
C13173 INVX1_LOC_75/Y INVX1_LOC_48/Y 0.06fF
C13174 INVX1_LOC_31/Y INVX1_LOC_665/A 0.18fF
C13175 INVX1_LOC_183/Y INVX1_LOC_63/Y 0.01fF
C13176 INVX1_LOC_47/Y INVX1_LOC_373/Y 0.00fF
C13177 INVX1_LOC_54/Y INVX1_LOC_75/A 0.03fF
C13178 NAND2X1_LOC_826/a_36_24# INVX1_LOC_658/Y 0.00fF
C13179 INVX1_LOC_49/Y NAND2X1_LOC_630/a_36_24# 0.01fF
C13180 INVX1_LOC_74/Y INVX1_LOC_93/A 0.00fF
C13181 INVX1_LOC_242/Y INVX1_LOC_9/Y 0.06fF
C13182 INVX1_LOC_89/Y NAND2X1_LOC_410/Y 0.17fF
C13183 VDD NAND2X1_LOC_76/B 0.17fF
C13184 NAND2X1_LOC_126/a_36_24# INVX1_LOC_26/Y 0.00fF
C13185 NAND2X1_LOC_274/B NAND2X1_LOC_657/a_36_24# 0.00fF
C13186 INVX1_LOC_267/A INVX1_LOC_91/Y 0.01fF
C13187 INVX1_LOC_48/Y NAND2X1_LOC_271/A 0.07fF
C13188 INVX1_LOC_100/Y INVX1_LOC_644/Y 0.01fF
C13189 NAND2X1_LOC_491/Y INVX1_LOC_75/Y 0.11fF
C13190 INVX1_LOC_93/Y INVX1_LOC_231/Y 0.05fF
C13191 INVX1_LOC_601/Y INVX1_LOC_620/Y 0.02fF
C13192 INVX1_LOC_63/Y INVX1_LOC_223/A 0.24fF
C13193 INVX1_LOC_62/Y INVX1_LOC_242/Y 0.08fF
C13194 INVX1_LOC_502/A INVX1_LOC_280/A 0.07fF
C13195 NAND2X1_LOC_301/B INVX1_LOC_347/A 0.07fF
C13196 NAND2X1_LOC_164/Y NAND2X1_LOC_241/B 0.05fF
C13197 INVX1_LOC_68/Y INVX1_LOC_560/Y 0.00fF
C13198 INVX1_LOC_404/Y INVX1_LOC_446/Y 0.17fF
C13199 NAND2X1_LOC_750/Y INVX1_LOC_65/Y 0.00fF
C13200 NAND2X1_LOC_334/A INVX1_LOC_636/A 0.02fF
C13201 INVX1_LOC_681/A INVX1_LOC_109/Y 0.01fF
C13202 INVX1_LOC_1/Y INVX1_LOC_41/A 0.01fF
C13203 INVX1_LOC_400/Y NAND2X1_LOC_498/Y 0.05fF
C13204 INVX1_LOC_406/Y INVX1_LOC_453/A 0.01fF
C13205 INVX1_LOC_563/Y INVX1_LOC_315/Y 0.07fF
C13206 INVX1_LOC_244/Y INVX1_LOC_443/A 0.10fF
C13207 NAND2X1_LOC_615/a_36_24# INVX1_LOC_211/A 0.00fF
C13208 NAND2X1_LOC_843/B INVX1_LOC_241/A 0.08fF
C13209 INVX1_LOC_206/Y INVX1_LOC_381/A 0.07fF
C13210 VDD INVX1_LOC_541/Y 0.21fF
C13211 INVX1_LOC_406/Y NAND2X1_LOC_271/B 0.01fF
C13212 NAND2X1_LOC_123/A INVX1_LOC_638/A 0.15fF
C13213 INVX1_LOC_224/Y INVX1_LOC_566/A 0.07fF
C13214 INVX1_LOC_618/A INVX1_LOC_252/Y 0.15fF
C13215 INVX1_LOC_560/Y INVX1_LOC_250/Y 0.07fF
C13216 NAND2X1_LOC_526/Y INVX1_LOC_586/A 0.21fF
C13217 INVX1_LOC_285/A INVX1_LOC_292/A 0.21fF
C13218 NAND2X1_LOC_756/a_36_24# INVX1_LOC_396/Y 0.00fF
C13219 INVX1_LOC_53/Y INVX1_LOC_549/A 0.07fF
C13220 INVX1_LOC_625/A VDD 0.19fF
C13221 INVX1_LOC_220/Y NAND2X1_LOC_261/Y 0.01fF
C13222 INVX1_LOC_395/A INVX1_LOC_80/A 0.23fF
C13223 INVX1_LOC_604/Y NAND2X1_LOC_241/B 0.03fF
C13224 INVX1_LOC_498/A INVX1_LOC_638/A 0.07fF
C13225 VDD INVX1_LOC_294/A 0.00fF
C13226 INVX1_LOC_434/A INVX1_LOC_437/A 0.03fF
C13227 INVX1_LOC_404/Y INVX1_LOC_145/Y 0.03fF
C13228 NAND2X1_LOC_331/A INVX1_LOC_145/Y 0.03fF
C13229 INVX1_LOC_53/Y INVX1_LOC_624/A 0.02fF
C13230 INVX1_LOC_172/Y INVX1_LOC_175/A 0.14fF
C13231 INVX1_LOC_400/Y INVX1_LOC_99/Y 0.03fF
C13232 INVX1_LOC_278/Y INVX1_LOC_445/A 0.01fF
C13233 VDD INVX1_LOC_208/Y 0.22fF
C13234 INVX1_LOC_206/Y NAND2X1_LOC_720/A 0.01fF
C13235 INVX1_LOC_562/A INVX1_LOC_674/A 0.05fF
C13236 INVX1_LOC_90/A INVX1_LOC_76/Y 0.01fF
C13237 INVX1_LOC_11/Y INVX1_LOC_395/A 0.66fF
C13238 NAND2X1_LOC_780/A INVX1_LOC_581/A 0.05fF
C13239 INPUT_7 INVX1_LOC_55/Y 0.06fF
C13240 INVX1_LOC_27/A INPUT_2 0.01fF
C13241 INVX1_LOC_335/Y INVX1_LOC_526/A 0.05fF
C13242 INVX1_LOC_521/Y INVX1_LOC_137/Y 0.02fF
C13243 NAND2X1_LOC_544/a_36_24# INVX1_LOC_116/Y 0.00fF
C13244 INVX1_LOC_165/Y INVX1_LOC_137/Y 0.15fF
C13245 INVX1_LOC_80/A INVX1_LOC_683/Y 0.02fF
C13246 INVX1_LOC_45/Y INVX1_LOC_98/Y 0.02fF
C13247 INVX1_LOC_11/Y INVX1_LOC_362/Y 0.15fF
C13248 INVX1_LOC_84/A INVX1_LOC_600/A 0.03fF
C13249 VDD NAND2X1_LOC_52/Y 0.01fF
C13250 INVX1_LOC_564/A INVX1_LOC_93/Y 0.03fF
C13251 INVX1_LOC_53/Y INVX1_LOC_635/A 0.02fF
C13252 INPUT_0 NAND2X1_LOC_308/A 0.15fF
C13253 INVX1_LOC_191/A INVX1_LOC_145/Y 0.01fF
C13254 INVX1_LOC_301/A INVX1_LOC_9/Y 0.03fF
C13255 INVX1_LOC_584/A INVX1_LOC_47/Y 0.02fF
C13256 NAND2X1_LOC_635/B INVX1_LOC_586/A 0.01fF
C13257 NAND2X1_LOC_707/A INVX1_LOC_513/A 0.02fF
C13258 INVX1_LOC_44/A INVX1_LOC_184/A 0.01fF
C13259 INVX1_LOC_17/Y INVX1_LOC_661/A 0.08fF
C13260 INVX1_LOC_54/Y NAND2X1_LOC_318/A 0.13fF
C13261 NAND2X1_LOC_318/A NAND2X1_LOC_614/a_36_24# 0.01fF
C13262 INVX1_LOC_11/Y INVX1_LOC_683/Y 0.02fF
C13263 INVX1_LOC_558/A INVX1_LOC_199/A 0.01fF
C13264 INVX1_LOC_418/A INVX1_LOC_89/Y 0.02fF
C13265 INVX1_LOC_558/A INVX1_LOC_89/Y 0.24fF
C13266 VDD INVX1_LOC_519/Y 0.41fF
C13267 INVX1_LOC_676/Y INVX1_LOC_537/A 0.02fF
C13268 NAND2X1_LOC_338/a_36_24# INVX1_LOC_50/Y 0.00fF
C13269 INVX1_LOC_171/Y INVX1_LOC_46/Y 0.03fF
C13270 INVX1_LOC_548/A INVX1_LOC_80/A 0.15fF
C13271 INVX1_LOC_224/Y NAND2X1_LOC_558/B 0.05fF
C13272 INVX1_LOC_522/Y INVX1_LOC_138/Y 0.01fF
C13273 NAND2X1_LOC_595/Y INVX1_LOC_503/A 0.10fF
C13274 INVX1_LOC_301/A INVX1_LOC_62/Y 0.02fF
C13275 INVX1_LOC_206/Y INVX1_LOC_100/Y 0.55fF
C13276 INVX1_LOC_666/A INVX1_LOC_199/Y 0.03fF
C13277 INVX1_LOC_20/Y INVX1_LOC_155/A 0.02fF
C13278 INVX1_LOC_224/Y INVX1_LOC_79/A 0.06fF
C13279 INVX1_LOC_584/A INVX1_LOC_119/Y 0.02fF
C13280 INVX1_LOC_84/A INVX1_LOC_484/A 0.01fF
C13281 INVX1_LOC_270/A INVX1_LOC_89/Y 0.00fF
C13282 INVX1_LOC_188/Y INVX1_LOC_50/Y 0.00fF
C13283 INPUT_7 INVX1_LOC_18/Y 0.44fF
C13284 NAND2X1_LOC_111/Y INVX1_LOC_119/A 0.07fF
C13285 INVX1_LOC_17/Y INVX1_LOC_352/Y 0.03fF
C13286 INVX1_LOC_392/A INVX1_LOC_367/Y 0.00fF
C13287 INVX1_LOC_80/A INVX1_LOC_31/Y 0.23fF
C13288 INVX1_LOC_343/Y INVX1_LOC_69/A 0.02fF
C13289 INVX1_LOC_578/A INVX1_LOC_79/A 0.07fF
C13290 INVX1_LOC_545/A INVX1_LOC_159/Y 0.01fF
C13291 INVX1_LOC_579/Y INVX1_LOC_31/Y 0.05fF
C13292 INVX1_LOC_370/A NAND2X1_LOC_464/a_36_24# 0.02fF
C13293 INVX1_LOC_542/Y NAND2X1_LOC_829/Y 0.09fF
C13294 INVX1_LOC_557/A INVX1_LOC_79/A 0.05fF
C13295 INVX1_LOC_116/Y INVX1_LOC_360/A 0.39fF
C13296 INVX1_LOC_206/Y INVX1_LOC_74/Y 1.77fF
C13297 INVX1_LOC_335/A INVX1_LOC_137/Y 5.09fF
C13298 INVX1_LOC_569/A NAND2X1_LOC_846/B 0.04fF
C13299 INVX1_LOC_540/Y INVX1_LOC_479/A 0.04fF
C13300 INVX1_LOC_628/Y INVX1_LOC_93/Y 0.01fF
C13301 INVX1_LOC_54/Y INVX1_LOC_202/Y 0.03fF
C13302 INVX1_LOC_206/Y INVX1_LOC_483/Y 0.01fF
C13303 INVX1_LOC_468/Y INVX1_LOC_469/Y 0.02fF
C13304 INVX1_LOC_468/Y INVX1_LOC_350/Y 0.02fF
C13305 INVX1_LOC_17/Y NAND2X1_LOC_504/a_36_24# 0.00fF
C13306 INVX1_LOC_20/Y INVX1_LOC_9/Y 0.83fF
C13307 INVX1_LOC_258/A INVX1_LOC_63/Y 0.01fF
C13308 INVX1_LOC_555/A NAND2X1_LOC_610/a_36_24# -0.02fF
C13309 INVX1_LOC_672/Y INVX1_LOC_283/A 0.01fF
C13310 INVX1_LOC_595/Y INVX1_LOC_117/Y 0.25fF
C13311 INVX1_LOC_566/Y NAND2X1_LOC_334/B 0.14fF
C13312 INVX1_LOC_117/Y INVX1_LOC_304/Y 0.02fF
C13313 INVX1_LOC_89/Y NAND2X1_LOC_755/B 0.03fF
C13314 INVX1_LOC_63/Y INVX1_LOC_489/Y 0.03fF
C13315 INVX1_LOC_155/A INVX1_LOC_300/A 0.01fF
C13316 INVX1_LOC_53/Y NAND2X1_LOC_817/a_36_24# 0.00fF
C13317 INVX1_LOC_54/Y INVX1_LOC_550/A 0.03fF
C13318 INVX1_LOC_583/A INVX1_LOC_168/Y 0.02fF
C13319 INVX1_LOC_47/Y INVX1_LOC_537/A 0.03fF
C13320 INVX1_LOC_439/Y INVX1_LOC_444/A -0.04fF
C13321 INVX1_LOC_682/A INVX1_LOC_134/Y 0.01fF
C13322 INVX1_LOC_21/A INVX1_LOC_9/Y 0.09fF
C13323 INVX1_LOC_11/Y INVX1_LOC_31/Y 1.93fF
C13324 INVX1_LOC_155/A INVX1_LOC_197/Y 0.01fF
C13325 INVX1_LOC_607/A NAND2X1_LOC_247/a_36_24# 0.00fF
C13326 INVX1_LOC_345/A NAND2X1_LOC_435/a_36_24# 0.02fF
C13327 INVX1_LOC_80/A INVX1_LOC_682/Y 0.01fF
C13328 INVX1_LOC_159/Y INVX1_LOC_230/Y 0.09fF
C13329 NAND2X1_LOC_387/Y INVX1_LOC_50/Y 0.07fF
C13330 INVX1_LOC_418/A NAND2X1_LOC_544/B 0.03fF
C13331 INVX1_LOC_145/Y INVX1_LOC_182/Y 0.02fF
C13332 INVX1_LOC_211/Y INVX1_LOC_89/Y 0.11fF
C13333 INVX1_LOC_385/A NAND2X1_LOC_479/a_36_24# 0.02fF
C13334 INVX1_LOC_447/Y INVX1_LOC_49/Y 0.02fF
C13335 INVX1_LOC_293/Y INVX1_LOC_90/Y 0.00fF
C13336 INVX1_LOC_69/Y INVX1_LOC_304/A 0.01fF
C13337 INVX1_LOC_686/A INVX1_LOC_100/Y 0.04fF
C13338 INVX1_LOC_69/Y INVX1_LOC_35/Y 2.61fF
C13339 NAND2X1_LOC_673/A INVX1_LOC_199/Y 0.23fF
C13340 INVX1_LOC_20/Y INVX1_LOC_62/Y 10.46fF
C13341 INVX1_LOC_54/Y INVX1_LOC_387/Y 0.03fF
C13342 INVX1_LOC_267/A NAND2X1_LOC_333/B 0.02fF
C13343 NAND2X1_LOC_106/Y NAND2X1_LOC_693/a_36_24# 0.00fF
C13344 INVX1_LOC_374/A INVX1_LOC_348/Y 0.02fF
C13345 INVX1_LOC_49/Y NAND2X1_LOC_602/A 0.06fF
C13346 INVX1_LOC_273/A NAND2X1_LOC_242/a_36_24# 0.01fF
C13347 INVX1_LOC_300/A INVX1_LOC_9/Y 1.10fF
C13348 INVX1_LOC_89/Y INVX1_LOC_46/Y 0.06fF
C13349 INVX1_LOC_54/Y INVX1_LOC_49/Y 0.26fF
C13350 INVX1_LOC_576/A INVX1_LOC_62/Y 0.11fF
C13351 INVX1_LOC_398/A INVX1_LOC_211/A 0.03fF
C13352 INVX1_LOC_686/A INVX1_LOC_74/Y 0.62fF
C13353 INVX1_LOC_379/A INVX1_LOC_247/Y 0.01fF
C13354 INVX1_LOC_508/A INVX1_LOC_138/Y 0.01fF
C13355 NAND2X1_LOC_833/B INVX1_LOC_145/Y 0.03fF
C13356 NAND2X1_LOC_97/B INVX1_LOC_41/Y 0.04fF
C13357 INVX1_LOC_201/Y INVX1_LOC_26/Y 0.22fF
C13358 INVX1_LOC_69/Y INVX1_LOC_620/A 0.03fF
C13359 INVX1_LOC_468/Y INVX1_LOC_79/A 0.04fF
C13360 INVX1_LOC_6/Y NAND2X1_LOC_612/a_36_24# 0.00fF
C13361 INVX1_LOC_89/Y NAND2X1_LOC_305/a_36_24# 0.00fF
C13362 INVX1_LOC_11/Y INVX1_LOC_128/A 0.02fF
C13363 INVX1_LOC_183/A INVX1_LOC_117/Y 0.16fF
C13364 INVX1_LOC_69/Y NAND2X1_LOC_253/Y 0.02fF
C13365 INVX1_LOC_524/Y INVX1_LOC_91/Y 0.28fF
C13366 INVX1_LOC_479/A NAND2X1_LOC_496/Y 0.02fF
C13367 NAND2X1_LOC_706/a_36_24# INVX1_LOC_100/Y 0.01fF
C13368 INVX1_LOC_300/A INVX1_LOC_62/Y 0.14fF
C13369 INVX1_LOC_491/A INVX1_LOC_50/Y 0.08fF
C13370 NAND2X1_LOC_531/Y INVX1_LOC_63/Y 0.03fF
C13371 INVX1_LOC_449/A NAND2X1_LOC_255/a_36_24# 0.00fF
C13372 INVX1_LOC_17/Y NAND2X1_LOC_372/Y 0.03fF
C13373 INVX1_LOC_62/Y INVX1_LOC_197/Y 0.01fF
C13374 INVX1_LOC_543/Y INVX1_LOC_26/Y 0.01fF
C13375 INVX1_LOC_41/Y INVX1_LOC_510/A 0.07fF
C13376 INVX1_LOC_669/Y NAND2X1_LOC_843/B 0.01fF
C13377 INVX1_LOC_31/Y NAND2X1_LOC_433/Y 0.18fF
C13378 INVX1_LOC_41/Y INVX1_LOC_440/Y 0.03fF
C13379 INVX1_LOC_116/Y INVX1_LOC_364/A 0.02fF
C13380 INVX1_LOC_44/Y NAND2X1_LOC_759/Y 0.04fF
C13381 NAND2X1_LOC_775/B INVX1_LOC_479/A 0.46fF
C13382 NAND2X1_LOC_768/B INVX1_LOC_63/Y 0.04fF
C13383 INVX1_LOC_632/Y INVX1_LOC_639/A 0.01fF
C13384 INVX1_LOC_59/Y NAND2X1_LOC_98/B 0.01fF
C13385 INVX1_LOC_660/A INVX1_LOC_342/A 0.03fF
C13386 INVX1_LOC_120/Y INVX1_LOC_79/A 0.03fF
C13387 INVX1_LOC_46/Y NAND2X1_LOC_544/B 0.03fF
C13388 INVX1_LOC_438/Y INVX1_LOC_220/A 0.06fF
C13389 INVX1_LOC_183/Y INVX1_LOC_81/A 0.05fF
C13390 INVX1_LOC_117/Y INVX1_LOC_109/A -0.00fF
C13391 INVX1_LOC_257/Y INVX1_LOC_638/A 0.01fF
C13392 INVX1_LOC_211/A NAND2X1_LOC_203/a_36_24# 0.00fF
C13393 INVX1_LOC_93/Y INVX1_LOC_625/Y 0.02fF
C13394 INVX1_LOC_390/A INVX1_LOC_319/A 0.11fF
C13395 INVX1_LOC_502/A INVX1_LOC_328/Y 0.01fF
C13396 INVX1_LOC_93/Y INVX1_LOC_91/Y 0.09fF
C13397 NAND2X1_LOC_334/A INVX1_LOC_74/Y 0.03fF
C13398 INVX1_LOC_49/Y INVX1_LOC_388/A 0.00fF
C13399 INVX1_LOC_434/A INVX1_LOC_438/Y 0.03fF
C13400 VDD NAND2X1_LOC_164/Y 0.10fF
C13401 INVX1_LOC_288/A INVX1_LOC_638/A 1.41fF
C13402 NAND2X1_LOC_242/A INVX1_LOC_206/Y 0.01fF
C13403 NAND2X1_LOC_123/B INVX1_LOC_114/A 0.03fF
C13404 INVX1_LOC_63/Y NAND2X1_LOC_832/A 0.03fF
C13405 INVX1_LOC_63/Y INVX1_LOC_443/A 0.03fF
C13406 INVX1_LOC_577/Y INVX1_LOC_458/Y 0.01fF
C13407 INVX1_LOC_62/Y NAND2X1_LOC_269/B 0.02fF
C13408 INVX1_LOC_400/Y NAND2X1_LOC_475/A 0.03fF
C13409 VDD INVX1_LOC_65/Y 0.59fF
C13410 VDD INVX1_LOC_220/Y 0.21fF
C13411 INVX1_LOC_564/A INVX1_LOC_395/A 0.00fF
C13412 INVX1_LOC_228/Y INVX1_LOC_65/Y 0.02fF
C13413 VDD INVX1_LOC_501/Y 0.25fF
C13414 INVX1_LOC_393/Y INVX1_LOC_392/Y 0.05fF
C13415 INVX1_LOC_203/Y INVX1_LOC_287/Y 0.02fF
C13416 INVX1_LOC_454/A INVX1_LOC_59/A 0.03fF
C13417 NAND2X1_LOC_498/Y INVX1_LOC_570/A 0.08fF
C13418 VDD INVX1_LOC_184/A 0.02fF
C13419 INVX1_LOC_435/Y INVX1_LOC_45/Y 0.06fF
C13420 INVX1_LOC_395/A NAND2X1_LOC_704/B 0.45fF
C13421 NAND2X1_LOC_61/A NAND2X1_LOC_318/B 0.28fF
C13422 INVX1_LOC_145/Y INVX1_LOC_638/A 0.07fF
C13423 INVX1_LOC_629/A INVX1_LOC_686/A 0.02fF
C13424 INVX1_LOC_634/Y INVX1_LOC_347/A 0.09fF
C13425 NAND2X1_LOC_269/B NAND2X1_LOC_269/a_36_24# 0.01fF
C13426 NAND2X1_LOC_317/A NAND2X1_LOC_307/A 0.43fF
C13427 VDD INVX1_LOC_604/Y 0.50fF
C13428 NAND2X1_LOC_515/a_36_24# NAND2X1_LOC_513/Y 0.00fF
C13429 INPUT_0 INVX1_LOC_134/Y 0.17fF
C13430 INVX1_LOC_53/Y INVX1_LOC_292/A 0.01fF
C13431 INVX1_LOC_20/Y NAND2X1_LOC_392/a_36_24# 0.00fF
C13432 NAND2X1_LOC_498/Y INVX1_LOC_377/Y 0.01fF
C13433 INVX1_LOC_390/Y INVX1_LOC_320/A 0.00fF
C13434 VDD INVX1_LOC_427/Y 0.21fF
C13435 INVX1_LOC_224/Y INVX1_LOC_417/Y 0.03fF
C13436 NAND2X1_LOC_45/Y INVX1_LOC_99/Y 0.22fF
C13437 INVX1_LOC_255/Y INVX1_LOC_197/A 0.03fF
C13438 INVX1_LOC_607/Y INVX1_LOC_238/Y 0.05fF
C13439 INVX1_LOC_374/A INVX1_LOC_258/A 0.01fF
C13440 INVX1_LOC_317/Y NAND2X1_LOC_543/a_36_24# 0.00fF
C13441 INVX1_LOC_596/A INVX1_LOC_45/Y 0.05fF
C13442 VDD INVX1_LOC_479/Y 0.24fF
C13443 INVX1_LOC_447/A INVX1_LOC_159/A 0.04fF
C13444 INVX1_LOC_428/A INVX1_LOC_387/A 0.27fF
C13445 INVX1_LOC_86/Y INVX1_LOC_180/Y 0.64fF
C13446 INVX1_LOC_434/A INVX1_LOC_219/Y 0.00fF
C13447 INVX1_LOC_80/A INVX1_LOC_51/Y 0.18fF
C13448 NAND2X1_LOC_537/B INVX1_LOC_35/Y 0.05fF
C13449 INVX1_LOC_236/A INVX1_LOC_395/A 0.01fF
C13450 NAND2X1_LOC_12/a_36_24# INVX1_LOC_53/Y 0.00fF
C13451 NAND2X1_LOC_318/B INVX1_LOC_45/Y 0.04fF
C13452 INVX1_LOC_224/Y INVX1_LOC_48/Y 0.69fF
C13453 INVX1_LOC_446/Y INVX1_LOC_451/A 0.10fF
C13454 NAND2X1_LOC_750/Y INVX1_LOC_86/Y 0.11fF
C13455 INVX1_LOC_592/Y NAND2X1_LOC_759/B 0.21fF
C13456 INVX1_LOC_266/A INVX1_LOC_80/A 0.01fF
C13457 VDD INVX1_LOC_397/Y 0.28fF
C13458 INVX1_LOC_362/Y INVX1_LOC_367/Y 0.03fF
C13459 INVX1_LOC_586/A INVX1_LOC_379/A 0.10fF
C13460 NAND2X1_LOC_331/A INVX1_LOC_522/A 0.00fF
C13461 INVX1_LOC_166/A INVX1_LOC_553/Y 0.00fF
C13462 INVX1_LOC_84/A NAND2X1_LOC_56/Y 0.00fF
C13463 INVX1_LOC_425/A NAND2X1_LOC_102/a_36_24# 0.00fF
C13464 INVX1_LOC_578/A INVX1_LOC_48/Y 0.04fF
C13465 INVX1_LOC_442/A INVX1_LOC_350/A 0.01fF
C13466 INVX1_LOC_53/Y INVX1_LOC_492/Y 0.09fF
C13467 INVX1_LOC_228/Y INVX1_LOC_318/A 0.16fF
C13468 NAND2X1_LOC_45/Y INVX1_LOC_47/Y 0.11fF
C13469 INVX1_LOC_586/A INVX1_LOC_35/Y 1.96fF
C13470 INVX1_LOC_586/A INVX1_LOC_304/A 0.00fF
C13471 INVX1_LOC_11/Y INVX1_LOC_51/Y 8.70fF
C13472 INVX1_LOC_424/Y INVX1_LOC_385/Y 0.12fF
C13473 NAND2X1_LOC_534/Y INVX1_LOC_49/Y 0.04fF
C13474 INVX1_LOC_628/A INVX1_LOC_686/A 0.02fF
C13475 INVX1_LOC_444/Y INVX1_LOC_384/Y 0.00fF
C13476 INVX1_LOC_504/A INVX1_LOC_348/A 0.03fF
C13477 INVX1_LOC_166/A INVX1_LOC_546/A 0.03fF
C13478 INVX1_LOC_52/Y INVX1_LOC_255/A 0.04fF
C13479 VDD INVX1_LOC_314/Y 0.26fF
C13480 INVX1_LOC_10/Y INVX1_LOC_9/A 0.00fF
C13481 NAND2X1_LOC_111/Y INVX1_LOC_410/Y 0.07fF
C13482 NAND2X1_LOC_750/Y INVX1_LOC_63/Y 0.00fF
C13483 INVX1_LOC_246/Y INVX1_LOC_379/A 0.05fF
C13484 NAND2X1_LOC_174/B INVX1_LOC_577/Y 0.00fF
C13485 INVX1_LOC_26/Y INVX1_LOC_458/Y 0.01fF
C13486 INVX1_LOC_137/A INVX1_LOC_46/Y 0.01fF
C13487 NAND2X1_LOC_106/Y INVX1_LOC_547/Y 0.04fF
C13488 INVX1_LOC_384/A INVX1_LOC_665/Y 0.04fF
C13489 INVX1_LOC_449/Y INVX1_LOC_406/Y 0.02fF
C13490 INVX1_LOC_65/Y INVX1_LOC_68/A 0.02fF
C13491 INVX1_LOC_21/Y NAND2X1_LOC_97/B 0.07fF
C13492 INVX1_LOC_564/Y NAND2X1_LOC_753/Y 0.00fF
C13493 INVX1_LOC_312/Y INVX1_LOC_379/A 0.14fF
C13494 INVX1_LOC_54/Y INVX1_LOC_76/Y 0.16fF
C13495 INVX1_LOC_570/A INVX1_LOC_568/A -0.00fF
C13496 NAND2X1_LOC_300/a_36_24# INVX1_LOC_374/A 0.00fF
C13497 NAND2X1_LOC_79/B INVX1_LOC_198/Y 0.01fF
C13498 NAND2X1_LOC_498/Y INVX1_LOC_47/Y 0.14fF
C13499 NAND2X1_LOC_241/B INVX1_LOC_63/Y 0.60fF
C13500 INVX1_LOC_570/A INVX1_LOC_47/Y 0.07fF
C13501 INVX1_LOC_312/Y INVX1_LOC_35/Y 0.06fF
C13502 NAND2X1_LOC_781/A INVX1_LOC_35/Y 0.02fF
C13503 NAND2X1_LOC_507/A NAND2X1_LOC_318/A 0.04fF
C13504 INVX1_LOC_449/A INVX1_LOC_17/Y 0.07fF
C13505 INVX1_LOC_586/A INVX1_LOC_620/A 0.07fF
C13506 INVX1_LOC_93/Y INVX1_LOC_142/Y 0.01fF
C13507 INVX1_LOC_402/A NAND2X1_LOC_284/a_36_24# 0.01fF
C13508 NAND2X1_LOC_574/a_36_24# NAND2X1_LOC_542/A 0.01fF
C13509 INVX1_LOC_12/Y NAND2X1_LOC_266/a_36_24# 0.01fF
C13510 VDD INVX1_LOC_244/Y 1.29fF
C13511 INVX1_LOC_290/Y INVX1_LOC_300/Y 0.00fF
C13512 INVX1_LOC_133/A NAND2X1_LOC_286/a_36_24# 0.00fF
C13513 INVX1_LOC_259/A INVX1_LOC_188/A 0.35fF
C13514 NAND2X1_LOC_132/a_36_24# NAND2X1_LOC_332/B 0.00fF
C13515 INVX1_LOC_17/Y INVX1_LOC_67/Y 0.13fF
C13516 INVX1_LOC_33/Y NAND2X1_LOC_836/B 0.02fF
C13517 INVX1_LOC_206/Y INVX1_LOC_77/A 0.01fF
C13518 INVX1_LOC_524/Y NAND2X1_LOC_333/B 0.12fF
C13519 INVX1_LOC_320/A INVX1_LOC_432/A 0.57fF
C13520 INVX1_LOC_583/A INVX1_LOC_137/Y 0.01fF
C13521 INVX1_LOC_20/Y INVX1_LOC_87/A 0.12fF
C13522 NAND2X1_LOC_45/Y NAND2X1_LOC_66/Y 0.03fF
C13523 INVX1_LOC_356/A INVX1_LOC_463/Y 0.02fF
C13524 INVX1_LOC_245/A INVX1_LOC_49/A 0.01fF
C13525 INVX1_LOC_553/Y NAND2X1_LOC_136/Y 0.12fF
C13526 INVX1_LOC_469/Y INVX1_LOC_686/A 0.03fF
C13527 INVX1_LOC_686/A INVX1_LOC_350/Y -0.00fF
C13528 INVX1_LOC_18/Y INVX1_LOC_55/Y 0.14fF
C13529 NAND2X1_LOC_24/Y INVX1_LOC_50/Y 0.01fF
C13530 INVX1_LOC_206/Y INVX1_LOC_79/A 1.01fF
C13531 INVX1_LOC_176/A INVX1_LOC_7/Y 0.43fF
C13532 INVX1_LOC_589/Y NAND2X1_LOC_508/a_36_24# 0.01fF
C13533 NAND2X1_LOC_180/B NAND2X1_LOC_388/A 0.02fF
C13534 INVX1_LOC_444/Y NAND2X1_LOC_416/Y 0.03fF
C13535 NAND2X1_LOC_697/Y INVX1_LOC_145/Y 0.01fF
C13536 INPUT_7 INVX1_LOC_343/Y 0.01fF
C13537 INVX1_LOC_324/Y INVX1_LOC_327/Y 0.21fF
C13538 INVX1_LOC_106/A INVX1_LOC_662/Y 0.02fF
C13539 INVX1_LOC_451/A INVX1_LOC_145/Y 0.03fF
C13540 NAND2X1_LOC_574/a_36_24# INVX1_LOC_376/Y 0.00fF
C13541 INVX1_LOC_448/A INVX1_LOC_665/Y 0.02fF
C13542 NAND2X1_LOC_529/Y INVX1_LOC_35/Y 0.01fF
C13543 NAND2X1_LOC_97/B NAND2X1_LOC_267/A 0.02fF
C13544 INVX1_LOC_550/A NAND2X1_LOC_677/Y 0.01fF
C13545 INVX1_LOC_147/A INVX1_LOC_493/A 0.19fF
C13546 VDD INVX1_LOC_588/A 0.56fF
C13547 INVX1_LOC_412/Y INVX1_LOC_41/Y 0.14fF
C13548 INVX1_LOC_261/Y INVX1_LOC_59/A 0.05fF
C13549 INVX1_LOC_116/Y INVX1_LOC_350/A 0.02fF
C13550 INVX1_LOC_53/Y NAND2X1_LOC_285/A 0.46fF
C13551 INVX1_LOC_76/Y INVX1_LOC_521/A 0.01fF
C13552 NAND2X1_LOC_498/Y INVX1_LOC_119/Y 0.09fF
C13553 INVX1_LOC_439/Y INVX1_LOC_451/Y 0.04fF
C13554 NAND2X1_LOC_505/a_36_24# INVX1_LOC_100/Y 0.00fF
C13555 INVX1_LOC_21/Y INVX1_LOC_280/Y 0.04fF
C13556 INVX1_LOC_570/A INVX1_LOC_119/Y 0.03fF
C13557 INVX1_LOC_145/Y INVX1_LOC_665/Y 0.04fF
C13558 INVX1_LOC_65/Y NAND2X1_LOC_786/B 0.83fF
C13559 INVX1_LOC_53/Y NAND2X1_LOC_647/A 0.00fF
C13560 NAND2X1_LOC_396/a_36_24# NAND2X1_LOC_396/Y 0.02fF
C13561 INVX1_LOC_44/A INVX1_LOC_86/Y 0.01fF
C13562 INVX1_LOC_397/A INVX1_LOC_100/Y 0.37fF
C13563 NAND2X1_LOC_317/B INVX1_LOC_479/A 0.14fF
C13564 INVX1_LOC_316/Y INVX1_LOC_298/A 0.02fF
C13565 INVX1_LOC_617/Y INVX1_LOC_301/Y 0.46fF
C13566 INVX1_LOC_395/A NAND2X1_LOC_843/B 0.13fF
C13567 INVX1_LOC_103/Y INVX1_LOC_370/A 0.01fF
C13568 INVX1_LOC_176/A INVX1_LOC_32/Y 0.01fF
C13569 INVX1_LOC_31/Y INVX1_LOC_367/Y 0.03fF
C13570 INVX1_LOC_84/A INVX1_LOC_183/Y 0.02fF
C13571 INVX1_LOC_589/Y INVX1_LOC_99/Y 0.01fF
C13572 INVX1_LOC_662/A NAND2X1_LOC_846/a_36_24# 0.01fF
C13573 INVX1_LOC_89/Y INVX1_LOC_115/A 0.01fF
C13574 INVX1_LOC_53/Y INVX1_LOC_168/Y 0.07fF
C13575 INVX1_LOC_588/Y INVX1_LOC_674/A 0.19fF
C13576 INVX1_LOC_49/Y INVX1_LOC_371/Y 0.04fF
C13577 NAND2X1_LOC_145/a_36_24# NAND2X1_LOC_847/A 0.00fF
C13578 NAND2X1_LOC_527/Y INVX1_LOC_48/Y 0.01fF
C13579 INVX1_LOC_47/Y INVX1_LOC_99/Y 1.30fF
C13580 INVX1_LOC_313/Y INVX1_LOC_31/Y 0.01fF
C13581 INVX1_LOC_227/Y INVX1_LOC_48/Y 0.02fF
C13582 INVX1_LOC_417/Y INVX1_LOC_120/Y 0.04fF
C13583 NAND2X1_LOC_557/B INVX1_LOC_99/Y 0.31fF
C13584 INVX1_LOC_451/A INVX1_LOC_433/A 0.09fF
C13585 INVX1_LOC_654/A INVX1_LOC_100/Y 0.02fF
C13586 NAND2X1_LOC_829/Y NAND2X1_LOC_679/A 0.02fF
C13587 INVX1_LOC_377/Y INVX1_LOC_119/Y 0.09fF
C13588 INVX1_LOC_69/Y INVX1_LOC_357/A 0.01fF
C13589 INVX1_LOC_361/Y INVX1_LOC_93/Y 0.14fF
C13590 INVX1_LOC_686/A INVX1_LOC_79/A 0.14fF
C13591 INVX1_LOC_662/Y INVX1_LOC_239/A 0.38fF
C13592 INVX1_LOC_214/Y INVX1_LOC_69/Y 0.53fF
C13593 INVX1_LOC_63/Y NAND2X1_LOC_621/a_36_24# 0.00fF
C13594 INVX1_LOC_93/Y NAND2X1_LOC_333/B 0.10fF
C13595 NAND2X1_LOC_274/B INVX1_LOC_519/A 0.02fF
C13596 NAND2X1_LOC_755/B INVX1_LOC_44/Y 0.09fF
C13597 INVX1_LOC_84/A INVX1_LOC_369/Y 0.91fF
C13598 INVX1_LOC_69/Y NAND2X1_LOC_837/B 0.32fF
C13599 INVX1_LOC_617/Y INVX1_LOC_41/Y 0.15fF
C13600 NAND2X1_LOC_140/B INVX1_LOC_9/Y 0.09fF
C13601 INVX1_LOC_17/Y INVX1_LOC_347/Y 0.67fF
C13602 INVX1_LOC_119/A INVX1_LOC_41/Y 0.06fF
C13603 INVX1_LOC_255/A INVX1_LOC_350/A 0.05fF
C13604 INVX1_LOC_31/Y INVX1_LOC_374/Y 0.03fF
C13605 INVX1_LOC_520/Y INVX1_LOC_556/Y 0.01fF
C13606 INVX1_LOC_147/A INVX1_LOC_500/A 0.23fF
C13607 INVX1_LOC_686/A INVX1_LOC_460/A 0.01fF
C13608 INVX1_LOC_444/Y NAND2X1_LOC_555/B 0.00fF
C13609 INVX1_LOC_69/Y INVX1_LOC_360/A 0.01fF
C13610 INVX1_LOC_452/A NAND2X1_LOC_481/a_36_24# 0.01fF
C13611 INVX1_LOC_379/A INVX1_LOC_225/Y 0.04fF
C13612 INVX1_LOC_17/Y INVX1_LOC_328/Y 0.08fF
C13613 INVX1_LOC_295/Y INVX1_LOC_296/A 0.22fF
C13614 INVX1_LOC_208/A INVX1_LOC_69/Y 0.15fF
C13615 INVX1_LOC_93/Y INVX1_LOC_261/Y 0.00fF
C13616 INVX1_LOC_99/Y INVX1_LOC_119/Y 0.03fF
C13617 NAND2X1_LOC_755/a_36_24# INVX1_LOC_26/Y 0.00fF
C13618 INVX1_LOC_410/A INVX1_LOC_32/Y 0.00fF
C13619 INVX1_LOC_79/A INVX1_LOC_14/A 0.01fF
C13620 INVX1_LOC_50/A INVX1_LOC_40/Y 0.03fF
C13621 NAND2X1_LOC_630/a_36_24# INVX1_LOC_7/Y 0.00fF
C13622 INVX1_LOC_382/A INVX1_LOC_63/Y 0.03fF
C13623 NAND2X1_LOC_426/Y INVX1_LOC_462/Y 0.01fF
C13624 INVX1_LOC_170/Y INVX1_LOC_32/Y 0.06fF
C13625 INVX1_LOC_99/Y NAND2X1_LOC_66/Y 1.64fF
C13626 INVX1_LOC_479/A INVX1_LOC_633/Y 0.07fF
C13627 NAND2X1_LOC_306/a_36_24# INVX1_LOC_47/Y 0.01fF
C13628 NAND2X1_LOC_301/B INVX1_LOC_252/Y 0.02fF
C13629 INVX1_LOC_232/Y INVX1_LOC_280/A 0.04fF
C13630 INVX1_LOC_47/Y NAND2X1_LOC_557/B 0.94fF
C13631 INVX1_LOC_89/Y INVX1_LOC_49/Y 1.02fF
C13632 NAND2X1_LOC_174/B INVX1_LOC_26/Y 0.00fF
C13633 INPUT_3 NAND2X1_LOC_416/B 0.01fF
C13634 INVX1_LOC_282/A INVX1_LOC_100/Y 0.00fF
C13635 INVX1_LOC_105/A INVX1_LOC_519/Y 0.00fF
C13636 INVX1_LOC_261/Y INVX1_LOC_675/A 0.02fF
C13637 INVX1_LOC_399/Y INVX1_LOC_32/Y 0.02fF
C13638 INVX1_LOC_386/A NAND2X1_LOC_483/a_36_24# 0.02fF
C13639 INVX1_LOC_89/Y INVX1_LOC_533/A 0.01fF
C13640 NAND2X1_LOC_35/a_36_24# INVX1_LOC_190/A 0.01fF
C13641 INVX1_LOC_258/Y INVX1_LOC_675/A 0.32fF
C13642 NAND2X1_LOC_318/a_36_24# INVX1_LOC_100/Y 0.00fF
C13643 INVX1_LOC_582/A INVX1_LOC_168/Y 0.09fF
C13644 INVX1_LOC_49/Y INVX1_LOC_501/A 0.03fF
C13645 INVX1_LOC_183/A INVX1_LOC_58/Y 0.00fF
C13646 INVX1_LOC_31/Y INVX1_LOC_319/A 0.01fF
C13647 INVX1_LOC_31/Y NAND2X1_LOC_432/a_36_24# 0.00fF
C13648 NAND2X1_LOC_306/a_36_24# INVX1_LOC_119/Y 0.00fF
C13649 INVX1_LOC_501/A INVX1_LOC_533/A 0.05fF
C13650 INVX1_LOC_47/Y INVX1_LOC_119/Y 0.48fF
C13651 NAND2X1_LOC_542/A INVX1_LOC_100/Y 0.02fF
C13652 INVX1_LOC_69/Y INVX1_LOC_657/A 0.00fF
C13653 NAND2X1_LOC_334/A INVX1_LOC_79/A 0.02fF
C13654 INVX1_LOC_601/Y INVX1_LOC_597/Y 0.00fF
C13655 INVX1_LOC_317/A INVX1_LOC_479/A 0.01fF
C13656 INVX1_LOC_100/Y INVX1_LOC_376/Y 0.07fF
C13657 INVX1_LOC_31/Y INVX1_LOC_625/Y 0.03fF
C13658 NAND2X1_LOC_762/a_36_24# INVX1_LOC_33/A 0.00fF
C13659 INVX1_LOC_69/Y INVX1_LOC_495/Y 0.05fF
C13660 INVX1_LOC_69/Y INVX1_LOC_364/A 0.00fF
C13661 INVX1_LOC_107/Y NAND2X1_LOC_248/B 0.01fF
C13662 INVX1_LOC_199/Y INVX1_LOC_647/Y 0.03fF
C13663 INVX1_LOC_434/A INVX1_LOC_429/A 0.03fF
C13664 INVX1_LOC_376/Y INVX1_LOC_74/Y 0.10fF
C13665 NAND2X1_LOC_750/Y INVX1_LOC_552/Y 0.00fF
C13666 NAND2X1_LOC_283/a_36_24# INVX1_LOC_212/A 0.00fF
C13667 INVX1_LOC_97/Y INVX1_LOC_615/A 0.14fF
C13668 NAND2X1_LOC_176/Y INVX1_LOC_270/A 0.00fF
C13669 INVX1_LOC_612/A INVX1_LOC_611/A 0.16fF
C13670 INVX1_LOC_20/Y NAND2X1_LOC_331/A 0.03fF
C13671 VDD INVX1_LOC_434/Y 0.21fF
C13672 NAND2X1_LOC_498/Y INVX1_LOC_502/Y 0.02fF
C13673 VDD INVX1_LOC_670/Y 0.59fF
C13674 INVX1_LOC_257/Y INVX1_LOC_134/Y 1.00fF
C13675 INVX1_LOC_206/Y INVX1_LOC_632/A 0.07fF
C13676 INVX1_LOC_435/Y INVX1_LOC_293/Y 0.05fF
C13677 NAND2X1_LOC_704/B INVX1_LOC_51/Y 0.17fF
C13678 INVX1_LOC_20/Y INVX1_LOC_271/Y 0.02fF
C13679 INVX1_LOC_417/Y INVX1_LOC_206/Y 0.14fF
C13680 INVX1_LOC_21/Y INVX1_LOC_412/Y 0.03fF
C13681 INPUT_0 INVX1_LOC_16/Y 0.01fF
C13682 VDD INVX1_LOC_506/Y 0.29fF
C13683 INVX1_LOC_416/Y NAND2X1_LOC_391/A 0.00fF
C13684 NAND2X1_LOC_249/Y NAND2X1_LOC_106/B 0.02fF
C13685 INVX1_LOC_291/A INVX1_LOC_586/A 0.03fF
C13686 NAND2X1_LOC_475/A INVX1_LOC_99/Y 0.10fF
C13687 NAND2X1_LOC_525/Y INVX1_LOC_53/Y 0.07fF
C13688 INVX1_LOC_80/A NAND2X1_LOC_114/a_36_24# 0.00fF
C13689 INVX1_LOC_80/A INVX1_LOC_355/A 0.04fF
C13690 INVX1_LOC_80/A NAND2X1_LOC_108/Y 0.00fF
C13691 INVX1_LOC_206/Y INVX1_LOC_398/Y 0.03fF
C13692 INVX1_LOC_203/Y INVX1_LOC_202/Y 0.09fF
C13693 INVX1_LOC_570/A INVX1_LOC_136/Y 0.03fF
C13694 INVX1_LOC_542/A NAND2X1_LOC_681/a_36_24# -0.00fF
C13695 VDD NAND2X1_LOC_646/A -0.00fF
C13696 INVX1_LOC_206/Y INVX1_LOC_59/Y 0.03fF
C13697 INVX1_LOC_288/A INVX1_LOC_134/Y 0.00fF
C13698 VDD INVX1_LOC_623/Y 0.24fF
C13699 INVX1_LOC_17/Y NAND2X1_LOC_536/a_36_24# 0.00fF
C13700 INVX1_LOC_580/A INVX1_LOC_576/Y 0.00fF
C13701 NAND2X1_LOC_710/B INVX1_LOC_510/A 0.01fF
C13702 VDD INVX1_LOC_86/Y 0.64fF
C13703 NAND2X1_LOC_457/A INVX1_LOC_681/Y 0.00fF
C13704 INVX1_LOC_510/Y INVX1_LOC_670/Y 0.10fF
C13705 INVX1_LOC_206/Y INVX1_LOC_48/Y 0.40fF
C13706 INVX1_LOC_446/Y INVX1_LOC_235/A 0.03fF
C13707 NAND2X1_LOC_69/a_36_24# INVX1_LOC_178/A 0.00fF
C13708 NAND2X1_LOC_457/A INPUT_1 0.03fF
C13709 INVX1_LOC_625/A INVX1_LOC_45/Y 0.02fF
C13710 INVX1_LOC_271/Y INVX1_LOC_300/A 0.01fF
C13711 INVX1_LOC_11/Y INVX1_LOC_216/Y 0.01fF
C13712 INVX1_LOC_12/Y INVX1_LOC_169/A 0.04fF
C13713 NAND2X1_LOC_475/A INVX1_LOC_123/A 0.02fF
C13714 VDD INVX1_LOC_253/Y 0.29fF
C13715 INVX1_LOC_224/Y INVX1_LOC_559/Y 0.04fF
C13716 INVX1_LOC_17/Y INVX1_LOC_266/Y 2.46fF
C13717 INVX1_LOC_395/A INVX1_LOC_361/Y 0.10fF
C13718 INVX1_LOC_158/A INVX1_LOC_89/Y 0.05fF
C13719 INVX1_LOC_556/A INVX1_LOC_117/Y 0.22fF
C13720 INPUT_3 INVX1_LOC_530/A 0.08fF
C13721 INVX1_LOC_454/A INVX1_LOC_641/A 0.01fF
C13722 INVX1_LOC_17/Y INVX1_LOC_651/Y 0.07fF
C13723 NAND2X1_LOC_475/A INVX1_LOC_47/Y 0.03fF
C13724 INVX1_LOC_686/A INVX1_LOC_632/A 0.14fF
C13725 VDD INVX1_LOC_63/Y 2.15fF
C13726 INVX1_LOC_35/Y INVX1_LOC_366/A 0.00fF
C13727 INVX1_LOC_679/Y INVX1_LOC_651/A 0.00fF
C13728 NAND2X1_LOC_150/a_36_24# NAND2X1_LOC_775/B 0.00fF
C13729 INVX1_LOC_52/Y INVX1_LOC_69/Y 0.01fF
C13730 INVX1_LOC_586/A INVX1_LOC_360/A 0.01fF
C13731 INVX1_LOC_257/Y INVX1_LOC_65/A 0.03fF
C13732 INVX1_LOC_482/A INVX1_LOC_681/Y 0.01fF
C13733 INVX1_LOC_11/Y NAND2X1_LOC_13/Y 0.03fF
C13734 INVX1_LOC_379/A INVX1_LOC_486/Y 0.17fF
C13735 NAND2X1_LOC_755/B NAND2X1_LOC_837/a_36_24# 0.00fF
C13736 INVX1_LOC_272/Y INVX1_LOC_35/Y 0.01fF
C13737 INVX1_LOC_134/Y INVX1_LOC_145/Y 0.07fF
C13738 INVX1_LOC_136/Y INVX1_LOC_99/Y 0.08fF
C13739 NAND2X1_LOC_692/Y INVX1_LOC_367/A 0.05fF
C13740 INVX1_LOC_228/Y INVX1_LOC_63/Y 0.28fF
C13741 INVX1_LOC_35/Y NAND2X1_LOC_820/A 0.01fF
C13742 NAND2X1_LOC_498/B INVX1_LOC_89/Y 0.08fF
C13743 INVX1_LOC_175/A INVX1_LOC_172/A 0.18fF
C13744 INVX1_LOC_312/A INVX1_LOC_211/Y 0.01fF
C13745 INPUT_3 INVX1_LOC_294/A 0.01fF
C13746 INVX1_LOC_492/A INVX1_LOC_508/Y 0.02fF
C13747 INVX1_LOC_206/Y NAND2X1_LOC_434/B 0.02fF
C13748 INVX1_LOC_174/A INVX1_LOC_178/A 0.11fF
C13749 INVX1_LOC_47/A INVX1_LOC_145/Y 0.03fF
C13750 INVX1_LOC_686/A INVX1_LOC_48/Y 0.07fF
C13751 INVX1_LOC_53/Y INVX1_LOC_137/Y 0.38fF
C13752 INVX1_LOC_54/Y INVX1_LOC_12/A 0.01fF
C13753 INVX1_LOC_343/Y INVX1_LOC_55/Y 0.01fF
C13754 INVX1_LOC_361/Y INVX1_LOC_683/Y 0.13fF
C13755 NAND2X1_LOC_636/A INVX1_LOC_653/Y 0.02fF
C13756 INVX1_LOC_89/Y INVX1_LOC_76/Y 0.17fF
C13757 INVX1_LOC_45/Y NAND2X1_LOC_52/Y 0.00fF
C13758 INVX1_LOC_390/Y NAND2X1_LOC_558/B 0.42fF
C13759 INPUT_0 INVX1_LOC_90/Y 0.19fF
C13760 NAND2X1_LOC_210/A INVX1_LOC_186/A 0.02fF
C13761 NAND2X1_LOC_43/Y INVX1_LOC_99/Y 0.26fF
C13762 INVX1_LOC_145/Y INVX1_LOC_235/A 0.01fF
C13763 NAND2X1_LOC_791/B INVX1_LOC_620/A 0.68fF
C13764 INVX1_LOC_390/Y INVX1_LOC_79/A 0.01fF
C13765 INVX1_LOC_117/Y INVX1_LOC_188/Y 0.17fF
C13766 INVX1_LOC_45/Y NAND2X1_LOC_686/A 0.03fF
C13767 INVX1_LOC_455/Y INVX1_LOC_298/A 0.01fF
C13768 INVX1_LOC_506/Y INVX1_LOC_509/A 0.01fF
C13769 INVX1_LOC_50/Y NAND2X1_LOC_297/a_36_24# 0.00fF
C13770 INVX1_LOC_410/Y INVX1_LOC_41/Y 3.56fF
C13771 INVX1_LOC_268/Y INVX1_LOC_44/Y 0.03fF
C13772 INVX1_LOC_54/Y INVX1_LOC_7/Y 0.55fF
C13773 INVX1_LOC_202/Y INVX1_LOC_194/Y 0.40fF
C13774 NAND2X1_LOC_768/A NAND2X1_LOC_281/a_36_24# 0.00fF
C13775 NAND2X1_LOC_250/Y NAND2X1_LOC_843/A 0.00fF
C13776 NAND2X1_LOC_108/Y INVX1_LOC_102/Y 0.01fF
C13777 INVX1_LOC_568/A INVX1_LOC_136/Y 0.01fF
C13778 NAND2X1_LOC_142/Y INVX1_LOC_100/Y 0.01fF
C13779 INVX1_LOC_503/Y INVX1_LOC_665/Y 0.01fF
C13780 NAND2X1_LOC_403/A INVX1_LOC_50/Y 0.01fF
C13781 INVX1_LOC_545/Y INVX1_LOC_199/Y 0.03fF
C13782 INVX1_LOC_375/A INVX1_LOC_41/Y 0.00fF
C13783 INVX1_LOC_153/A INVX1_LOC_99/Y 0.01fF
C13784 NAND2X1_LOC_307/A INVX1_LOC_199/Y 0.04fF
C13785 INVX1_LOC_300/A NAND2X1_LOC_265/a_36_24# 0.02fF
C13786 INVX1_LOC_442/Y INVX1_LOC_93/Y 0.07fF
C13787 INVX1_LOC_168/A NAND2X1_LOC_192/A 0.02fF
C13788 INVX1_LOC_447/Y INVX1_LOC_32/Y 0.19fF
C13789 INVX1_LOC_272/Y INVX1_LOC_621/Y 0.05fF
C13790 INVX1_LOC_69/Y INVX1_LOC_536/A 0.03fF
C13791 INVX1_LOC_382/A NAND2X1_LOC_414/a_36_24# 0.00fF
C13792 INVX1_LOC_195/Y INVX1_LOC_198/A 0.12fF
C13793 NAND2X1_LOC_646/A NAND2X1_LOC_607/a_36_24# 0.02fF
C13794 INVX1_LOC_46/Y INVX1_LOC_365/A 0.01fF
C13795 INVX1_LOC_174/A INVX1_LOC_58/Y 0.01fF
C13796 INVX1_LOC_50/Y INVX1_LOC_259/Y 0.03fF
C13797 NAND2X1_LOC_334/A INVX1_LOC_632/A 0.07fF
C13798 INVX1_LOC_686/A NAND2X1_LOC_434/B 0.01fF
C13799 INVX1_LOC_96/A INVX1_LOC_99/Y 0.01fF
C13800 INVX1_LOC_403/Y INVX1_LOC_117/Y 0.04fF
C13801 INVX1_LOC_213/Y NAND2X1_LOC_482/Y 0.25fF
C13802 INVX1_LOC_69/Y INVX1_LOC_115/Y 0.01fF
C13803 INVX1_LOC_186/Y INVX1_LOC_189/A 0.03fF
C13804 INVX1_LOC_35/Y INVX1_LOC_6/Y 4.82fF
C13805 NAND2X1_LOC_65/Y INVX1_LOC_41/Y 0.01fF
C13806 INVX1_LOC_317/Y INVX1_LOC_479/A 0.14fF
C13807 INVX1_LOC_53/A INVX1_LOC_204/Y 0.16fF
C13808 INVX1_LOC_548/A NAND2X1_LOC_125/a_36_24# 0.00fF
C13809 NAND2X1_LOC_534/a_36_24# NAND2X1_LOC_274/B 0.00fF
C13810 INVX1_LOC_86/Y NAND2X1_LOC_243/A 0.02fF
C13811 INVX1_LOC_54/Y INVX1_LOC_32/Y 0.20fF
C13812 NAND2X1_LOC_387/Y INVX1_LOC_117/Y 0.61fF
C13813 INVX1_LOC_93/Y INVX1_LOC_578/Y 0.01fF
C13814 NAND2X1_LOC_320/Y INVX1_LOC_376/A 0.01fF
C13815 INVX1_LOC_69/Y INVX1_LOC_350/A 0.01fF
C13816 INVX1_LOC_586/A INVX1_LOC_364/A 0.01fF
C13817 INVX1_LOC_361/Y INVX1_LOC_31/Y 0.01fF
C13818 INVX1_LOC_567/Y INVX1_LOC_9/Y 0.12fF
C13819 INVX1_LOC_406/Y INVX1_LOC_41/Y 0.16fF
C13820 INVX1_LOC_281/A INVX1_LOC_31/Y 0.03fF
C13821 INVX1_LOC_99/Y INVX1_LOC_15/Y 0.06fF
C13822 INVX1_LOC_419/Y INVX1_LOC_199/Y 0.84fF
C13823 INVX1_LOC_582/A INVX1_LOC_137/Y 0.01fF
C13824 INVX1_LOC_63/Y INVX1_LOC_509/A 0.01fF
C13825 INVX1_LOC_51/Y INVX1_LOC_91/Y 0.03fF
C13826 INVX1_LOC_51/Y INVX1_LOC_625/Y 0.10fF
C13827 INVX1_LOC_523/Y INVX1_LOC_46/Y 0.18fF
C13828 INVX1_LOC_557/Y INVX1_LOC_251/A 0.11fF
C13829 INVX1_LOC_31/Y INVX1_LOC_261/Y 0.05fF
C13830 INVX1_LOC_399/Y NAND2X1_LOC_226/Y 0.21fF
C13831 INVX1_LOC_17/Y INVX1_LOC_224/A 0.03fF
C13832 INVX1_LOC_93/Y INVX1_LOC_532/Y 0.01fF
C13833 INVX1_LOC_183/A NAND2X1_LOC_672/a_36_24# 0.01fF
C13834 INVX1_LOC_575/A INVX1_LOC_655/A 0.17fF
C13835 NAND2X1_LOC_846/B INVX1_LOC_650/Y 0.08fF
C13836 INVX1_LOC_99/Y NAND2X1_LOC_627/Y 0.01fF
C13837 INVX1_LOC_318/Y INVX1_LOC_211/A 0.00fF
C13838 INVX1_LOC_298/A NAND2X1_LOC_669/a_36_24# 0.00fF
C13839 INVX1_LOC_659/A INVX1_LOC_340/A 0.07fF
C13840 INVX1_LOC_128/Y INVX1_LOC_510/A 0.01fF
C13841 INVX1_LOC_476/A INVX1_LOC_476/Y 0.04fF
C13842 INVX1_LOC_567/Y INVX1_LOC_62/Y 0.44fF
C13843 NAND2X1_LOC_43/Y NAND2X1_LOC_66/Y 0.03fF
C13844 INVX1_LOC_376/Y INVX1_LOC_350/Y 0.01fF
C13845 INVX1_LOC_527/Y INVX1_LOC_90/Y 0.47fF
C13846 INVX1_LOC_319/A NAND2X1_LOC_267/a_36_24# 0.00fF
C13847 INVX1_LOC_199/Y NAND2X1_LOC_342/A 0.02fF
C13848 INVX1_LOC_361/Y INVX1_LOC_128/A 0.04fF
C13849 INVX1_LOC_79/A INVX1_LOC_432/A 0.01fF
C13850 INVX1_LOC_54/Y INVX1_LOC_612/A 0.01fF
C13851 INVX1_LOC_117/Y INVX1_LOC_491/A 0.93fF
C13852 INVX1_LOC_50/Y INVX1_LOC_114/A 0.03fF
C13853 INVX1_LOC_207/Y INVX1_LOC_198/A 0.01fF
C13854 INVX1_LOC_298/A INVX1_LOC_90/Y 0.17fF
C13855 INVX1_LOC_525/Y NAND2X1_LOC_420/a_36_24# 0.00fF
C13856 INVX1_LOC_666/Y INVX1_LOC_230/A 0.07fF
C13857 INVX1_LOC_49/Y INVX1_LOC_44/Y 0.07fF
C13858 INVX1_LOC_611/Y INVX1_LOC_612/A 0.14fF
C13859 INVX1_LOC_674/A INVX1_LOC_41/Y 0.07fF
C13860 INVX1_LOC_53/Y NAND2X1_LOC_781/a_36_24# 0.00fF
C13861 INVX1_LOC_518/Y INVX1_LOC_6/Y 0.06fF
C13862 INVX1_LOC_642/Y INVX1_LOC_44/Y 0.11fF
C13863 INVX1_LOC_634/Y INVX1_LOC_252/Y 0.95fF
C13864 NAND2X1_LOC_334/A NAND2X1_LOC_434/B 0.07fF
C13865 INVX1_LOC_217/A INVX1_LOC_220/A 0.03fF
C13866 INVX1_LOC_63/Y NAND2X1_LOC_786/B 0.23fF
C13867 INVX1_LOC_32/Y INVX1_LOC_388/A 0.00fF
C13868 NAND2X1_LOC_106/Y INVX1_LOC_62/Y 0.04fF
C13869 INVX1_LOC_166/A INVX1_LOC_479/A 0.04fF
C13870 INVX1_LOC_592/Y INVX1_LOC_531/Y 0.03fF
C13871 INPUT_5 INVX1_LOC_261/A 0.04fF
C13872 INVX1_LOC_202/A INVX1_LOC_206/Y 0.01fF
C13873 NAND2X1_LOC_10/a_36_24# INVX1_LOC_578/A 0.00fF
C13874 INVX1_LOC_79/A INVX1_LOC_376/Y 0.24fF
C13875 INVX1_LOC_289/Y NAND2X1_LOC_801/A 0.01fF
C13876 NAND2X1_LOC_498/a_36_24# INVX1_LOC_74/Y 0.00fF
C13877 NAND2X1_LOC_370/a_36_24# INVX1_LOC_206/Y 0.00fF
C13878 INVX1_LOC_279/Y INVX1_LOC_445/Y 0.20fF
C13879 INVX1_LOC_74/Y NAND2X1_LOC_455/a_36_24# 0.00fF
C13880 NAND2X1_LOC_847/A INVX1_LOC_241/A 0.06fF
C13881 INVX1_LOC_400/Y NAND2X1_LOC_322/Y 0.06fF
C13882 VDD INVX1_LOC_552/Y 0.59fF
C13883 NAND2X1_LOC_61/A INVX1_LOC_65/Y 0.06fF
C13884 NAND2X1_LOC_66/Y NAND2X1_LOC_627/Y 0.01fF
C13885 INVX1_LOC_206/Y INVX1_LOC_561/Y 0.03fF
C13886 INVX1_LOC_351/A INVX1_LOC_211/A 0.02fF
C13887 INVX1_LOC_166/Y NAND2X1_LOC_123/B 0.01fF
C13888 NAND2X1_LOC_136/Y INVX1_LOC_479/A 0.04fF
C13889 INVX1_LOC_20/Y INVX1_LOC_638/A 0.14fF
C13890 NAND2X1_LOC_123/B INVX1_LOC_62/Y 0.09fF
C13891 INVX1_LOC_412/Y INVX1_LOC_255/Y 1.07fF
C13892 INVX1_LOC_211/A INVX1_LOC_90/Y 0.01fF
C13893 INVX1_LOC_270/Y INVX1_LOC_9/Y 0.02fF
C13894 INVX1_LOC_17/Y INVX1_LOC_109/Y 0.07fF
C13895 INVX1_LOC_52/Y INVX1_LOC_586/A 0.01fF
C13896 NAND2X1_LOC_164/Y INVX1_LOC_45/Y 0.03fF
C13897 INVX1_LOC_203/Y INVX1_LOC_76/Y 0.01fF
C13898 VDD INVX1_LOC_20/A -0.00fF
C13899 INVX1_LOC_436/A VDD 0.00fF
C13900 INVX1_LOC_393/Y INVX1_LOC_51/Y 0.02fF
C13901 INVX1_LOC_9/Y INVX1_LOC_92/A 0.13fF
C13902 NAND2X1_LOC_750/Y INVX1_LOC_84/A 0.12fF
C13903 INVX1_LOC_425/A INVX1_LOC_416/Y 0.09fF
C13904 INVX1_LOC_65/Y INVX1_LOC_45/Y 0.03fF
C13905 INVX1_LOC_414/Y INVX1_LOC_427/A 0.14fF
C13906 NAND2X1_LOC_503/B INVX1_LOC_274/A 0.06fF
C13907 NAND2X1_LOC_13/Y INVX1_LOC_319/Y 0.01fF
C13908 INVX1_LOC_405/A NAND2X1_LOC_520/a_36_24# 0.00fF
C13909 INVX1_LOC_617/A NAND2X1_LOC_498/Y 0.01fF
C13910 INVX1_LOC_160/A NAND2X1_LOC_76/B 0.02fF
C13911 INVX1_LOC_594/Y NAND2X1_LOC_856/a_36_24# 0.00fF
C13912 INVX1_LOC_62/Y INVX1_LOC_92/A 0.20fF
C13913 GATE_579 INVX1_LOC_384/Y 0.14fF
C13914 INVX1_LOC_558/A INVX1_LOC_126/A 0.10fF
C13915 NAND2X1_LOC_97/B INVX1_LOC_560/A 0.23fF
C13916 INVX1_LOC_224/Y INVX1_LOC_155/Y 0.01fF
C13917 INVX1_LOC_395/A INVX1_LOC_307/A 0.03fF
C13918 INVX1_LOC_267/Y INVX1_LOC_564/Y 0.92fF
C13919 INVX1_LOC_417/A INVX1_LOC_560/A 0.01fF
C13920 INVX1_LOC_454/A INVX1_LOC_40/Y 0.19fF
C13921 VDD INVX1_LOC_263/Y 0.21fF
C13922 INPUT_0 INVX1_LOC_98/Y 0.05fF
C13923 INVX1_LOC_20/Y INVX1_LOC_101/Y 0.01fF
C13924 NAND2X1_LOC_332/B INVX1_LOC_134/Y 0.02fF
C13925 INVX1_LOC_51/Y NAND2X1_LOC_802/a_36_24# 0.01fF
C13926 INVX1_LOC_206/Y INVX1_LOC_396/A 0.01fF
C13927 NAND2X1_LOC_249/Y NAND2X1_LOC_128/A 0.39fF
C13928 INVX1_LOC_554/A NAND2X1_LOC_307/B 0.31fF
C13929 NAND2X1_LOC_720/a_36_24# INVX1_LOC_586/A 0.00fF
C13930 INVX1_LOC_398/Y INVX1_LOC_397/A 0.01fF
C13931 INVX1_LOC_686/A NAND2X1_LOC_129/a_36_24# 0.00fF
C13932 NAND2X1_LOC_457/A INVX1_LOC_50/Y 0.03fF
C13933 INVX1_LOC_374/A INVX1_LOC_509/A 0.03fF
C13934 INVX1_LOC_33/A INVX1_LOC_6/A 0.37fF
C13935 INVX1_LOC_572/A INVX1_LOC_542/Y 0.00fF
C13936 INVX1_LOC_370/Y INVX1_LOC_384/A 0.01fF
C13937 INVX1_LOC_59/Y INVX1_LOC_94/A 0.01fF
C13938 INVX1_LOC_447/A INVX1_LOC_69/Y 0.00fF
C13939 INVX1_LOC_442/A NAND2X1_LOC_775/B 1.09fF
C13940 VDD NAND2X1_LOC_836/B 0.15fF
C13941 INVX1_LOC_21/A INVX1_LOC_10/Y 0.01fF
C13942 INVX1_LOC_53/Y NAND2X1_LOC_307/A 1.79fF
C13943 INVX1_LOC_397/A INVX1_LOC_48/Y 0.07fF
C13944 NAND2X1_LOC_331/A NAND2X1_LOC_687/a_36_24# 0.01fF
C13945 INVX1_LOC_118/Y INVX1_LOC_387/Y 0.29fF
C13946 INVX1_LOC_53/Y INVX1_LOC_545/Y 0.03fF
C13947 INVX1_LOC_93/Y INVX1_LOC_412/A 0.02fF
C13948 INVX1_LOC_586/A INVX1_LOC_350/A 0.01fF
C13949 INVX1_LOC_209/A INVX1_LOC_273/A 0.04fF
C13950 NAND2X1_LOC_379/Y NAND2X1_LOC_460/A 0.02fF
C13951 INVX1_LOC_432/Y NAND2X1_LOC_13/Y 0.01fF
C13952 NAND2X1_LOC_391/a_36_24# INVX1_LOC_11/Y 0.01fF
C13953 INVX1_LOC_17/Y NAND2X1_LOC_698/a_36_24# 0.00fF
C13954 NAND2X1_LOC_130/a_36_24# INVX1_LOC_47/Y 0.01fF
C13955 INVX1_LOC_442/Y INVX1_LOC_683/Y 0.23fF
C13956 INVX1_LOC_76/Y INVX1_LOC_194/Y 0.17fF
C13957 INVX1_LOC_97/Y NAND2X1_LOC_237/Y 0.63fF
C13958 INVX1_LOC_322/Y INVX1_LOC_328/A 0.01fF
C13959 INVX1_LOC_318/A INVX1_LOC_45/Y 0.00fF
C13960 INVX1_LOC_51/Y NAND2X1_LOC_333/B 1.25fF
C13961 INVX1_LOC_281/A INVX1_LOC_51/Y 0.03fF
C13962 NAND2X1_LOC_550/a_36_24# NAND2X1_LOC_346/B 0.00fF
C13963 INVX1_LOC_561/Y NAND2X1_LOC_334/A 0.03fF
C13964 INPUT_0 INVX1_LOC_338/Y 0.14fF
C13965 INVX1_LOC_206/Y NAND2X1_LOC_615/Y 0.03fF
C13966 VDD INVX1_LOC_81/A -0.00fF
C13967 INVX1_LOC_169/A NAND2X1_LOC_615/B 0.01fF
C13968 INVX1_LOC_378/A INVX1_LOC_50/Y 0.01fF
C13969 INVX1_LOC_233/Y INVX1_LOC_421/A 0.06fF
C13970 NAND2X1_LOC_638/A INVX1_LOC_99/Y 0.03fF
C13971 INVX1_LOC_448/A INVX1_LOC_370/Y 0.02fF
C13972 INVX1_LOC_425/A INVX1_LOC_46/Y 0.01fF
C13973 VDD INVX1_LOC_430/A -0.00fF
C13974 INVX1_LOC_397/Y INVX1_LOC_45/Y 0.01fF
C13975 INVX1_LOC_211/Y INVX1_LOC_297/A 0.04fF
C13976 INVX1_LOC_266/A INVX1_LOC_361/Y 0.07fF
C13977 NAND2X1_LOC_715/a_36_24# INVX1_LOC_6/Y 0.00fF
C13978 INVX1_LOC_171/Y INVX1_LOC_32/Y 0.05fF
C13979 INVX1_LOC_51/Y INVX1_LOC_261/Y 0.03fF
C13980 INVX1_LOC_412/Y INVX1_LOC_26/Y 0.03fF
C13981 INVX1_LOC_419/Y INVX1_LOC_53/Y 0.01fF
C13982 INPUT_2 INVX1_LOC_46/Y 0.06fF
C13983 INVX1_LOC_95/A NAND2X1_LOC_506/B 0.18fF
C13984 INVX1_LOC_625/A INVX1_LOC_160/A 0.03fF
C13985 VDD INVX1_LOC_454/Y 0.50fF
C13986 INVX1_LOC_676/Y INVX1_LOC_505/A 0.02fF
C13987 NAND2X1_LOC_523/B INVX1_LOC_362/A 0.25fF
C13988 INVX1_LOC_45/Y INVX1_LOC_95/A 0.00fF
C13989 NAND2X1_LOC_24/Y INVX1_LOC_117/Y 0.03fF
C13990 NAND2X1_LOC_97/B INVX1_LOC_603/A 0.21fF
C13991 NAND2X1_LOC_249/Y NAND2X1_LOC_248/B 0.00fF
C13992 INVX1_LOC_556/Y INVX1_LOC_124/Y 0.01fF
C13993 INVX1_LOC_459/Y INVX1_LOC_376/A 0.00fF
C13994 NAND2X1_LOC_130/a_36_24# INVX1_LOC_119/Y 0.00fF
C13995 NAND2X1_LOC_122/Y INVX1_LOC_347/Y 0.02fF
C13996 INVX1_LOC_552/Y NAND2X1_LOC_786/B 0.02fF
C13997 INVX1_LOC_619/A INVX1_LOC_86/Y 0.02fF
C13998 NAND2X1_LOC_336/B INVX1_LOC_93/Y 0.02fF
C13999 INVX1_LOC_335/Y INVX1_LOC_674/A 0.07fF
C14000 INVX1_LOC_282/A NAND2X1_LOC_261/a_36_24# 0.00fF
C14001 INVX1_LOC_337/Y INVX1_LOC_66/A 0.22fF
C14002 INVX1_LOC_586/A INVX1_LOC_223/Y 1.27fF
C14003 NAND2X1_LOC_692/Y INVX1_LOC_548/A 0.09fF
C14004 NAND2X1_LOC_775/B INVX1_LOC_116/Y 0.09fF
C14005 INVX1_LOC_79/A INVX1_LOC_253/A 0.03fF
C14006 INVX1_LOC_31/Y INVX1_LOC_307/A 0.02fF
C14007 NAND2X1_LOC_493/B INVX1_LOC_390/A 0.27fF
C14008 INVX1_LOC_227/Y INVX1_LOC_155/Y 0.02fF
C14009 NAND2X1_LOC_403/A INVX1_LOC_327/Y 0.00fF
C14010 INVX1_LOC_80/A NAND2X1_LOC_449/B 0.25fF
C14011 INVX1_LOC_442/Y INVX1_LOC_31/Y 0.07fF
C14012 NAND2X1_LOC_638/A INVX1_LOC_47/Y 1.94fF
C14013 INVX1_LOC_48/Y INVX1_LOC_432/A 0.00fF
C14014 INVX1_LOC_569/A INVX1_LOC_662/A 0.16fF
C14015 INVX1_LOC_587/A INVX1_LOC_657/A 0.04fF
C14016 INVX1_LOC_188/Y INVX1_LOC_58/Y 0.09fF
C14017 INVX1_LOC_303/Y INPUT_1 0.01fF
C14018 INVX1_LOC_33/Y NAND2X1_LOC_409/Y 0.04fF
C14019 INVX1_LOC_417/Y NAND2X1_LOC_542/A 0.02fF
C14020 NAND2X1_LOC_336/B INVX1_LOC_390/A 0.00fF
C14021 INVX1_LOC_603/Y INVX1_LOC_58/Y 0.03fF
C14022 NAND2X1_LOC_108/Y NAND2X1_LOC_843/B 0.02fF
C14023 INVX1_LOC_617/Y INVX1_LOC_128/Y 0.04fF
C14024 NAND2X1_LOC_755/B NAND2X1_LOC_827/Y 0.00fF
C14025 NAND2X1_LOC_851/a_36_24# INVX1_LOC_283/A -0.00fF
C14026 INVX1_LOC_54/Y INVX1_LOC_110/A 0.01fF
C14027 NAND2X1_LOC_13/Y INVX1_LOC_319/A 0.23fF
C14028 INVX1_LOC_101/Y INVX1_LOC_655/A 0.03fF
C14029 INVX1_LOC_45/Y INVX1_LOC_588/A 0.03fF
C14030 INPUT_5 INVX1_LOC_69/A 0.01fF
C14031 INVX1_LOC_17/Y INVX1_LOC_199/Y 0.19fF
C14032 INVX1_LOC_134/Y INVX1_LOC_242/Y 0.02fF
C14033 INVX1_LOC_369/A INVX1_LOC_485/Y 0.01fF
C14034 NAND2X1_LOC_507/A INVX1_LOC_32/Y 0.05fF
C14035 INVX1_LOC_295/A INVX1_LOC_79/A 0.01fF
C14036 INVX1_LOC_669/Y NAND2X1_LOC_847/A 0.01fF
C14037 INVX1_LOC_328/Y NAND2X1_LOC_393/Y 0.02fF
C14038 INVX1_LOC_53/Y INVX1_LOC_502/A 0.07fF
C14039 NAND2X1_LOC_775/B INVX1_LOC_255/A 0.59fF
C14040 INVX1_LOC_6/Y INVX1_LOC_118/A 0.01fF
C14041 INVX1_LOC_80/A NAND2X1_LOC_301/B 0.01fF
C14042 INVX1_LOC_154/Y INVX1_LOC_245/A 0.01fF
C14043 INVX1_LOC_442/Y INVX1_LOC_682/Y 0.01fF
C14044 INVX1_LOC_84/A NAND2X1_LOC_488/Y 0.01fF
C14045 INVX1_LOC_58/Y INVX1_LOC_478/Y 0.02fF
C14046 NAND2X1_LOC_677/Y INVX1_LOC_612/A 0.23fF
C14047 INVX1_LOC_6/Y INVX1_LOC_649/A 0.18fF
C14048 INVX1_LOC_21/Y INVX1_LOC_273/Y 0.01fF
C14049 INVX1_LOC_89/Y INVX1_LOC_32/Y 4.63fF
C14050 INVX1_LOC_171/A INVX1_LOC_63/Y 0.03fF
C14051 NAND2X1_LOC_622/a_36_24# INVX1_LOC_169/Y 0.00fF
C14052 INVX1_LOC_99/Y INVX1_LOC_353/A 0.01fF
C14053 INVX1_LOC_578/Y NAND2X1_LOC_675/B 0.01fF
C14054 NAND2X1_LOC_845/B INVX1_LOC_178/A 0.02fF
C14055 INVX1_LOC_154/A INVX1_LOC_32/Y 0.00fF
C14056 INVX1_LOC_12/Y INVX1_LOC_531/Y 0.02fF
C14057 INVX1_LOC_145/Y INVX1_LOC_90/Y 0.03fF
C14058 NAND2X1_LOC_184/Y INVX1_LOC_420/A 0.01fF
C14059 INVX1_LOC_26/Y NAND2X1_LOC_81/a_36_24# 0.00fF
C14060 NAND2X1_LOC_387/Y INVX1_LOC_58/Y 0.02fF
C14061 INVX1_LOC_519/A NAND2X1_LOC_372/Y 0.03fF
C14062 NAND2X1_LOC_164/a_36_24# INVX1_LOC_26/Y 0.00fF
C14063 INVX1_LOC_345/Y INVX1_LOC_501/A 0.03fF
C14064 NAND2X1_LOC_605/B INVX1_LOC_440/Y 0.03fF
C14065 NAND2X1_LOC_503/Y INVX1_LOC_44/Y 0.06fF
C14066 INVX1_LOC_275/Y INVX1_LOC_274/Y 0.24fF
C14067 INPUT_1 INVX1_LOC_9/Y 5.97fF
C14068 INVX1_LOC_32/Y INVX1_LOC_501/A 0.03fF
C14069 NAND2X1_LOC_307/B INVX1_LOC_199/Y 1.19fF
C14070 INVX1_LOC_637/Y INVX1_LOC_641/A 0.00fF
C14071 INVX1_LOC_532/Y NAND2X1_LOC_675/B 0.17fF
C14072 NAND2X1_LOC_325/B INVX1_LOC_666/Y 0.07fF
C14073 INVX1_LOC_575/Y INVX1_LOC_655/A 0.14fF
C14074 NAND2X1_LOC_274/B INVX1_LOC_670/A 0.39fF
C14075 INVX1_LOC_254/Y INVX1_LOC_41/Y 0.03fF
C14076 INVX1_LOC_62/Y INVX1_LOC_681/Y 0.01fF
C14077 INVX1_LOC_211/A INVX1_LOC_98/Y 0.01fF
C14078 INVX1_LOC_62/Y INPUT_1 0.07fF
C14079 NAND2X1_LOC_845/B INVX1_LOC_58/Y 0.03fF
C14080 INVX1_LOC_491/A INVX1_LOC_58/Y 0.04fF
C14081 VDD INVX1_LOC_405/A 0.00fF
C14082 INVX1_LOC_132/A INVX1_LOC_655/A 0.02fF
C14083 INVX1_LOC_574/A INVX1_LOC_133/Y 0.01fF
C14084 INVX1_LOC_100/Y INVX1_LOC_654/Y 0.29fF
C14085 INVX1_LOC_32/Y NAND2X1_LOC_544/B 0.02fF
C14086 NAND2X1_LOC_69/B INVX1_LOC_206/Y 0.02fF
C14087 VDD INVX1_LOC_560/Y 0.22fF
C14088 INVX1_LOC_309/Y INVX1_LOC_41/Y 0.01fF
C14089 NAND2X1_LOC_68/a_36_24# INVX1_LOC_395/A 0.00fF
C14090 INVX1_LOC_206/Y NAND2X1_LOC_374/a_36_24# 0.01fF
C14091 INVX1_LOC_58/Y INVX1_LOC_91/A 0.24fF
C14092 INVX1_LOC_409/Y NAND2X1_LOC_498/Y 0.03fF
C14093 INVX1_LOC_471/Y INVX1_LOC_473/Y 0.98fF
C14094 NAND2X1_LOC_448/B INVX1_LOC_636/A 0.04fF
C14095 NAND2X1_LOC_710/B INVX1_LOC_553/Y 0.06fF
C14096 INVX1_LOC_11/A INVX1_LOC_100/Y 0.02fF
C14097 INVX1_LOC_312/A INVX1_LOC_297/Y 0.00fF
C14098 INVX1_LOC_652/A INVX1_LOC_74/Y 0.04fF
C14099 INVX1_LOC_560/A NAND2X1_LOC_558/a_36_24# 0.00fF
C14100 VDD INVX1_LOC_512/A -0.00fF
C14101 INVX1_LOC_447/A INVX1_LOC_586/A 0.01fF
C14102 INVX1_LOC_582/Y VDD 0.21fF
C14103 INVX1_LOC_395/A INVX1_LOC_412/A 0.30fF
C14104 INVX1_LOC_479/A INVX1_LOC_41/Y 0.29fF
C14105 INVX1_LOC_206/Y INVX1_LOC_340/Y 0.53fF
C14106 NAND2X1_LOC_567/a_36_24# INVX1_LOC_51/Y 0.00fF
C14107 INVX1_LOC_438/A INVX1_LOC_378/A 0.01fF
C14108 VDD INVX1_LOC_84/A 1.40fF
C14109 NAND2X1_LOC_97/B NAND2X1_LOC_790/B 0.05fF
C14110 VDD INVX1_LOC_591/Y 0.21fF
C14111 INVX1_LOC_301/A INVX1_LOC_134/Y 0.03fF
C14112 INVX1_LOC_409/A NAND2X1_LOC_534/a_36_24# 0.00fF
C14113 NAND2X1_LOC_164/Y NAND2X1_LOC_756/Y 0.02fF
C14114 INVX1_LOC_230/Y INVX1_LOC_109/Y 0.09fF
C14115 INVX1_LOC_74/Y INVX1_LOC_462/Y 0.09fF
C14116 INVX1_LOC_428/A NAND2X1_LOC_705/a_36_24# 0.00fF
C14117 INVX1_LOC_266/Y INVX1_LOC_273/A 0.05fF
C14118 VDD INVX1_LOC_129/A 0.00fF
C14119 NAND2X1_LOC_336/B INVX1_LOC_395/A 0.44fF
C14120 VDD NAND2X1_LOC_67/Y 0.21fF
C14121 INPUT_0 NAND2X1_LOC_318/B 0.02fF
C14122 INVX1_LOC_400/Y NAND2X1_LOC_56/Y 0.01fF
C14123 INVX1_LOC_562/A INVX1_LOC_526/Y 0.02fF
C14124 INVX1_LOC_617/A INVX1_LOC_502/Y 0.00fF
C14125 INVX1_LOC_586/A INVX1_LOC_522/Y 0.05fF
C14126 INVX1_LOC_340/Y INVX1_LOC_686/A 0.07fF
C14127 INVX1_LOC_63/Y NAND2X1_LOC_227/a_36_24# 0.00fF
C14128 INVX1_LOC_257/Y INVX1_LOC_98/Y 0.10fF
C14129 NAND2X1_LOC_765/a_36_24# INVX1_LOC_117/Y 0.01fF
C14130 NAND2X1_LOC_523/B INVX1_LOC_384/A 0.07fF
C14131 NAND2X1_LOC_790/B INVX1_LOC_525/Y 0.02fF
C14132 INPUT_0 INVX1_LOC_177/A 0.03fF
C14133 INVX1_LOC_312/A INVX1_LOC_76/Y 0.01fF
C14134 INVX1_LOC_58/Y NAND2X1_LOC_801/A 0.03fF
C14135 NAND2X1_LOC_829/Y INVX1_LOC_515/A 0.02fF
C14136 INVX1_LOC_203/Y INVX1_LOC_32/Y 0.02fF
C14137 INVX1_LOC_20/Y INVX1_LOC_134/Y 0.07fF
C14138 INVX1_LOC_686/A INVX1_LOC_634/A 0.01fF
C14139 INVX1_LOC_442/Y INVX1_LOC_51/Y 0.07fF
C14140 NAND2X1_LOC_781/A INVX1_LOC_522/Y 0.05fF
C14141 INVX1_LOC_551/Y INVX1_LOC_80/A 0.19fF
C14142 INVX1_LOC_301/A INVX1_LOC_65/A 0.35fF
C14143 NAND2X1_LOC_843/a_36_24# NAND2X1_LOC_260/Y 0.00fF
C14144 INVX1_LOC_414/Y INVX1_LOC_428/Y 0.02fF
C14145 INVX1_LOC_459/Y INVX1_LOC_17/Y 0.06fF
C14146 NAND2X1_LOC_61/A INVX1_LOC_63/Y 0.01fF
C14147 INVX1_LOC_174/Y INVX1_LOC_44/A 0.00fF
C14148 INVX1_LOC_68/Y INVX1_LOC_99/Y 0.01fF
C14149 INVX1_LOC_289/Y INVX1_LOC_259/Y 0.01fF
C14150 INVX1_LOC_42/A INVX1_LOC_84/A 0.01fF
C14151 NAND2X1_LOC_45/Y INVX1_LOC_484/A -0.02fF
C14152 INVX1_LOC_434/A INVX1_LOC_6/Y 0.06fF
C14153 INVX1_LOC_118/Y INVX1_LOC_108/A 0.14fF
C14154 NAND2X1_LOC_770/A INVX1_LOC_44/Y 0.05fF
C14155 VDD INVX1_LOC_496/A 0.00fF
C14156 VDD INVX1_LOC_674/Y 0.35fF
C14157 NAND2X1_LOC_328/a_36_24# INPUT_4 0.00fF
C14158 INVX1_LOC_406/Y INVX1_LOC_444/Y 0.03fF
C14159 NAND2X1_LOC_523/B INVX1_LOC_145/Y 0.01fF
C14160 INVX1_LOC_11/Y INVX1_LOC_551/Y 0.10fF
C14161 INVX1_LOC_608/Y INVX1_LOC_53/Y 0.03fF
C14162 INVX1_LOC_435/Y INVX1_LOC_283/Y 0.16fF
C14163 INVX1_LOC_556/Y INVX1_LOC_336/Y 0.01fF
C14164 INVX1_LOC_17/Y INVX1_LOC_53/Y 0.30fF
C14165 NAND2X1_LOC_79/Y INVX1_LOC_198/A 0.06fF
C14166 INVX1_LOC_562/A NAND2X1_LOC_719/A 0.09fF
C14167 INVX1_LOC_111/A INVX1_LOC_259/Y 0.00fF
C14168 INVX1_LOC_395/A NAND2X1_LOC_847/A 0.01fF
C14169 NAND2X1_LOC_475/A INVX1_LOC_353/A 0.03fF
C14170 INVX1_LOC_99/Y INVX1_LOC_600/A 0.24fF
C14171 INVX1_LOC_412/Y NAND2X1_LOC_605/B 0.02fF
C14172 INVX1_LOC_295/A INVX1_LOC_48/Y 0.01fF
C14173 INVX1_LOC_312/Y INVX1_LOC_295/Y 0.01fF
C14174 INVX1_LOC_269/A INVX1_LOC_58/Y 0.11fF
C14175 INVX1_LOC_45/Y INVX1_LOC_63/Y 0.16fF
C14176 INVX1_LOC_340/Y NAND2X1_LOC_811/a_36_24# 0.00fF
C14177 INVX1_LOC_53/Y INVX1_LOC_650/Y 0.01fF
C14178 INVX1_LOC_370/Y INVX1_LOC_503/Y 0.08fF
C14179 NAND2X1_LOC_679/B INVX1_LOC_332/Y 0.01fF
C14180 INVX1_LOC_375/A INVX1_LOC_128/Y 0.01fF
C14181 INVX1_LOC_7/Y INVX1_LOC_194/Y 0.02fF
C14182 NAND2X1_LOC_336/B INVX1_LOC_31/Y 0.03fF
C14183 INVX1_LOC_228/A INVX1_LOC_194/Y 0.46fF
C14184 INVX1_LOC_172/A NAND2X1_LOC_393/Y 0.06fF
C14185 INVX1_LOC_602/A INVX1_LOC_204/Y 0.04fF
C14186 INVX1_LOC_17/Y INVX1_LOC_460/Y 0.03fF
C14187 INPUT_3 INVX1_LOC_63/Y 0.10fF
C14188 INVX1_LOC_53/Y NAND2X1_LOC_307/B 0.03fF
C14189 INVX1_LOC_35/Y NAND2X1_LOC_720/A 0.03fF
C14190 NAND2X1_LOC_24/Y INVX1_LOC_58/Y 0.01fF
C14191 INVX1_LOC_602/Y INVX1_LOC_641/Y 0.34fF
C14192 INVX1_LOC_193/Y INVX1_LOC_75/Y 0.00fF
C14193 NAND2X1_LOC_148/A NAND2X1_LOC_342/A 0.03fF
C14194 INVX1_LOC_69/Y NAND2X1_LOC_496/Y 0.21fF
C14195 NAND2X1_LOC_130/Y INVX1_LOC_47/Y 0.02fF
C14196 INVX1_LOC_47/Y INVX1_LOC_600/A 0.04fF
C14197 INVX1_LOC_303/Y INVX1_LOC_50/Y 0.01fF
C14198 INVX1_LOC_484/A INVX1_LOC_99/Y 0.01fF
C14199 NAND2X1_LOC_557/B INVX1_LOC_600/A 0.02fF
C14200 INVX1_LOC_117/Y INVX1_LOC_259/Y 0.03fF
C14201 INVX1_LOC_12/Y INVX1_LOC_411/Y 0.24fF
C14202 INPUT_5 INPUT_7 0.26fF
C14203 NAND2X1_LOC_106/Y NAND2X1_LOC_485/a_36_24# 0.00fF
C14204 INVX1_LOC_32/Y INVX1_LOC_194/Y 0.05fF
C14205 INVX1_LOC_134/A INVX1_LOC_62/Y 0.01fF
C14206 INVX1_LOC_366/A NAND2X1_LOC_243/a_36_24# 0.01fF
C14207 INVX1_LOC_587/Y INVX1_LOC_50/Y 0.03fF
C14208 NAND2X1_LOC_184/Y INVX1_LOC_54/Y 0.54fF
C14209 INVX1_LOC_385/Y GATE_479 0.05fF
C14210 INVX1_LOC_436/A INVX1_LOC_430/Y 0.01fF
C14211 INVX1_LOC_21/Y INVX1_LOC_309/Y 0.01fF
C14212 INPUT_7 INVX1_LOC_2/Y 0.02fF
C14213 INVX1_LOC_491/Y INVX1_LOC_139/Y 0.00fF
C14214 INVX1_LOC_145/Y INVX1_LOC_497/A 0.04fF
C14215 INVX1_LOC_145/Y INVX1_LOC_338/Y 0.03fF
C14216 INVX1_LOC_49/Y INVX1_LOC_252/Y 0.09fF
C14217 INVX1_LOC_20/Y NAND2X1_LOC_791/a_36_24# 0.01fF
C14218 INVX1_LOC_44/Y INVX1_LOC_7/Y 0.01fF
C14219 INVX1_LOC_44/Y INVX1_LOC_228/A 0.06fF
C14220 INVX1_LOC_400/A INVX1_LOC_77/Y 0.43fF
C14221 NAND2X1_LOC_775/B INVX1_LOC_69/Y 0.11fF
C14222 INVX1_LOC_63/Y NAND2X1_LOC_69/Y 0.01fF
C14223 INVX1_LOC_603/Y INVX1_LOC_245/A 0.03fF
C14224 INVX1_LOC_576/Y INVX1_LOC_26/Y 0.02fF
C14225 INVX1_LOC_166/A INVX1_LOC_127/Y 0.03fF
C14226 INVX1_LOC_684/A INVX1_LOC_674/Y 0.00fF
C14227 INVX1_LOC_573/Y NAND2X1_LOC_728/A 0.10fF
C14228 INVX1_LOC_89/Y INVX1_LOC_110/A 0.01fF
C14229 INVX1_LOC_366/A NAND2X1_LOC_771/a_36_24# 0.00fF
C14230 INVX1_LOC_671/Y INVX1_LOC_283/A 0.12fF
C14231 INVX1_LOC_166/A INVX1_LOC_66/A 0.06fF
C14232 INVX1_LOC_117/Y INVX1_LOC_204/Y 0.05fF
C14233 NAND2X1_LOC_130/Y INVX1_LOC_119/Y 0.01fF
C14234 INVX1_LOC_419/A INVX1_LOC_46/Y 0.01fF
C14235 INVX1_LOC_54/Y INVX1_LOC_551/A 0.04fF
C14236 INVX1_LOC_674/A NAND2X1_LOC_290/a_36_24# 0.00fF
C14237 INVX1_LOC_12/Y INVX1_LOC_41/Y 0.06fF
C14238 GATE_662 NAND2X1_LOC_663/a_36_24# 0.02fF
C14239 NAND2X1_LOC_465/a_36_24# INVX1_LOC_9/Y 0.00fF
C14240 INVX1_LOC_251/A INVX1_LOC_79/A 0.15fF
C14241 INVX1_LOC_32/Y INVX1_LOC_44/Y 0.47fF
C14242 INVX1_LOC_21/Y NAND2X1_LOC_528/Y 0.07fF
C14243 INVX1_LOC_50/Y INVX1_LOC_9/Y 7.51fF
C14244 INVX1_LOC_35/Y INVX1_LOC_100/Y 1.93fF
C14245 INVX1_LOC_358/Y INVX1_LOC_479/A 0.79fF
C14246 INVX1_LOC_304/A INVX1_LOC_100/Y 0.00fF
C14247 INVX1_LOC_145/A NAND2X1_LOC_836/B 0.05fF
C14248 INVX1_LOC_335/Y INVX1_LOC_479/A 0.03fF
C14249 INVX1_LOC_674/A INVX1_LOC_26/Y 0.07fF
C14250 INVX1_LOC_21/Y INVX1_LOC_479/A 0.25fF
C14251 NAND2X1_LOC_836/B NAND2X1_LOC_824/a_36_24# 0.00fF
C14252 INVX1_LOC_141/Y INVX1_LOC_338/Y 0.01fF
C14253 INVX1_LOC_117/Y INVX1_LOC_114/A 0.03fF
C14254 INVX1_LOC_99/A INVX1_LOC_666/Y 0.03fF
C14255 INVX1_LOC_80/A INVX1_LOC_634/Y 0.17fF
C14256 INVX1_LOC_525/Y NAND2X1_LOC_420/Y 0.04fF
C14257 INVX1_LOC_35/Y INVX1_LOC_74/Y 0.05fF
C14258 INVX1_LOC_137/Y INVX1_LOC_653/Y 0.53fF
C14259 INVX1_LOC_662/A NAND2X1_LOC_342/A 0.07fF
C14260 INVX1_LOC_35/Y INVX1_LOC_483/Y 0.00fF
C14261 NAND2X1_LOC_136/Y INVX1_LOC_66/A 0.01fF
C14262 INVX1_LOC_484/A NAND2X1_LOC_66/Y 0.01fF
C14263 INVX1_LOC_62/Y INVX1_LOC_50/Y 16.25fF
C14264 INVX1_LOC_54/Y INVX1_LOC_75/Y 0.10fF
C14265 INVX1_LOC_177/A INVX1_LOC_64/Y 0.01fF
C14266 NAND2X1_LOC_684/a_36_24# INVX1_LOC_245/A 0.00fF
C14267 NAND2X1_LOC_521/Y INVX1_LOC_41/Y 0.83fF
C14268 INVX1_LOC_479/A NAND2X1_LOC_267/A 0.04fF
C14269 INVX1_LOC_11/Y INVX1_LOC_634/Y 0.07fF
C14270 NAND2X1_LOC_137/A INVX1_LOC_479/A 0.01fF
C14271 INVX1_LOC_587/Y INVX1_LOC_658/Y 0.16fF
C14272 INVX1_LOC_575/A INVX1_LOC_92/A 0.44fF
C14273 INVX1_LOC_484/Y INVX1_LOC_90/Y 0.01fF
C14274 INVX1_LOC_517/Y INVX1_LOC_62/Y 0.01fF
C14275 NAND2X1_LOC_61/A INVX1_LOC_552/Y 0.15fF
C14276 NAND2X1_LOC_475/A NAND2X1_LOC_335/B 0.01fF
C14277 INVX1_LOC_54/Y NAND2X1_LOC_271/A 0.25fF
C14278 INVX1_LOC_107/Y INVX1_LOC_479/A 0.02fF
C14279 INVX1_LOC_363/A INVX1_LOC_66/A 0.01fF
C14280 INVX1_LOC_652/A INVX1_LOC_79/A 0.01fF
C14281 INVX1_LOC_183/A INVX1_LOC_483/A -0.02fF
C14282 NAND2X1_LOC_99/a_36_24# INVX1_LOC_586/A 0.00fF
C14283 INVX1_LOC_560/A INVX1_LOC_410/Y 0.46fF
C14284 VDD INVX1_LOC_174/Y 0.35fF
C14285 VDD NAND2X1_LOC_79/B 0.38fF
C14286 NAND2X1_LOC_537/B INVX1_LOC_173/A 0.03fF
C14287 INVX1_LOC_68/Y NAND2X1_LOC_475/A 0.02fF
C14288 INVX1_LOC_20/Y NAND2X1_LOC_598/a_36_24# 0.00fF
C14289 INVX1_LOC_435/Y INVX1_LOC_446/Y 0.00fF
C14290 INVX1_LOC_521/Y INVX1_LOC_523/A 0.00fF
C14291 INVX1_LOC_552/Y INVX1_LOC_45/Y 0.00fF
C14292 INVX1_LOC_362/Y INVX1_LOC_215/Y 0.03fF
C14293 NAND2X1_LOC_231/A INVX1_LOC_395/A 0.02fF
C14294 INVX1_LOC_374/A INVX1_LOC_45/Y 0.03fF
C14295 NAND2X1_LOC_373/Y INVX1_LOC_134/Y 0.04fF
C14296 INVX1_LOC_62/Y INVX1_LOC_658/Y 0.03fF
C14297 INVX1_LOC_447/A INVX1_LOC_486/Y 0.03fF
C14298 INVX1_LOC_173/A INVX1_LOC_586/A 0.03fF
C14299 INVX1_LOC_435/Y INVX1_LOC_384/A 0.10fF
C14300 INVX1_LOC_266/A INVX1_LOC_412/A 0.03fF
C14301 INVX1_LOC_529/Y INVX1_LOC_658/Y 0.01fF
C14302 INPUT_0 INVX1_LOC_541/Y 0.01fF
C14303 INVX1_LOC_374/A INVX1_LOC_348/A 0.01fF
C14304 INVX1_LOC_20/Y NAND2X1_LOC_830/a_36_24# -0.00fF
C14305 NAND2X1_LOC_320/a_36_24# NAND2X1_LOC_320/Y 0.02fF
C14306 INVX1_LOC_239/Y NAND2X1_LOC_148/B 0.08fF
C14307 VDD INVX1_LOC_62/A -0.00fF
C14308 INVX1_LOC_418/A INVX1_LOC_80/A 0.01fF
C14309 INVX1_LOC_625/A INPUT_0 0.01fF
C14310 NAND2X1_LOC_242/A INVX1_LOC_35/Y 0.02fF
C14311 INVX1_LOC_558/A INVX1_LOC_80/A 0.07fF
C14312 VDD INVX1_LOC_156/A -0.00fF
C14313 INVX1_LOC_45/Y INVX1_LOC_387/A 0.01fF
C14314 INVX1_LOC_596/A INVX1_LOC_384/A 0.07fF
C14315 VDD NAND2X1_LOC_822/Y 0.03fF
C14316 NAND2X1_LOC_388/a_36_24# INVX1_LOC_270/A 0.00fF
C14317 INVX1_LOC_435/Y INVX1_LOC_145/Y 0.18fF
C14318 NAND2X1_LOC_788/A INVX1_LOC_166/A 0.02fF
C14319 NAND2X1_LOC_176/Y INVX1_LOC_32/Y 0.03fF
C14320 INVX1_LOC_435/Y INVX1_LOC_661/Y 0.06fF
C14321 INVX1_LOC_206/Y INVX1_LOC_315/A 0.04fF
C14322 INVX1_LOC_287/Y INVX1_LOC_80/A 0.04fF
C14323 NAND2X1_LOC_457/A INVX1_LOC_117/Y 0.03fF
C14324 INVX1_LOC_140/Y NAND2X1_LOC_606/Y 0.21fF
C14325 NAND2X1_LOC_525/Y INVX1_LOC_391/Y 0.01fF
C14326 NAND2X1_LOC_759/B INVX1_LOC_69/Y 0.01fF
C14327 INVX1_LOC_434/A NAND2X1_LOC_294/Y 0.06fF
C14328 INVX1_LOC_492/A INVX1_LOC_605/A 0.01fF
C14329 VDD NAND2X1_LOC_532/Y 0.24fF
C14330 INVX1_LOC_578/A INVX1_LOC_349/A 0.04fF
C14331 INPUT_0 INVX1_LOC_520/A 0.00fF
C14332 INVX1_LOC_118/Y INVX1_LOC_32/Y 0.00fF
C14333 VDD NAND2X1_LOC_376/B 0.04fF
C14334 NAND2X1_LOC_775/B INVX1_LOC_586/A 0.13fF
C14335 INVX1_LOC_448/A INVX1_LOC_596/A 0.07fF
C14336 NAND2X1_LOC_156/a_36_24# INVX1_LOC_186/A 0.00fF
C14337 NAND2X1_LOC_271/B INVX1_LOC_69/Y 0.28fF
C14338 INVX1_LOC_683/A INVX1_LOC_367/A 0.04fF
C14339 NAND2X1_LOC_317/B INVX1_LOC_69/Y 0.02fF
C14340 INVX1_LOC_85/Y NAND2X1_LOC_222/a_36_24# 0.00fF
C14341 INVX1_LOC_97/A INVX1_LOC_69/Y 0.00fF
C14342 INVX1_LOC_96/Y INVX1_LOC_32/Y 0.40fF
C14343 NAND2X1_LOC_7/Y INVX1_LOC_90/Y -0.01fF
C14344 INVX1_LOC_452/Y INVX1_LOC_671/A 0.14fF
C14345 INVX1_LOC_300/A INVX1_LOC_318/Y 0.01fF
C14346 INVX1_LOC_565/Y INVX1_LOC_300/A 0.05fF
C14347 INVX1_LOC_596/A INVX1_LOC_145/Y 0.02fF
C14348 INVX1_LOC_133/Y INVX1_LOC_667/A 0.01fF
C14349 INVX1_LOC_137/Y NAND2X1_LOC_783/a_36_24# 0.00fF
C14350 INVX1_LOC_21/Y INVX1_LOC_12/Y 0.01fF
C14351 NAND2X1_LOC_56/Y INVX1_LOC_99/Y 0.00fF
C14352 INVX1_LOC_68/Y INVX1_LOC_153/A 0.02fF
C14353 INVX1_LOC_293/Y NAND2X1_LOC_250/Y 0.01fF
C14354 NAND2X1_LOC_123/B INVX1_LOC_638/A 0.01fF
C14355 NAND2X1_LOC_38/a_36_24# INVX1_LOC_600/A 0.00fF
C14356 INVX1_LOC_117/Y INVX1_LOC_482/A 0.03fF
C14357 VDD INVX1_LOC_106/Y 0.21fF
C14358 NAND2X1_LOC_79/B NAND2X1_LOC_243/A 0.01fF
C14359 NAND2X1_LOC_370/A INVX1_LOC_199/Y 0.05fF
C14360 INVX1_LOC_229/Y INVX1_LOC_194/Y 0.03fF
C14361 INVX1_LOC_27/Y INVX1_LOC_7/Y 0.15fF
C14362 INVX1_LOC_442/A NAND2X1_LOC_111/Y 0.49fF
C14363 INVX1_LOC_53/Y INVX1_LOC_108/Y 0.01fF
C14364 NAND2X1_LOC_532/Y INVX1_LOC_510/Y 0.00fF
C14365 NAND2X1_LOC_318/B INVX1_LOC_145/Y 0.01fF
C14366 INVX1_LOC_45/Y NAND2X1_LOC_836/B 0.02fF
C14367 INVX1_LOC_523/A NAND2X1_LOC_846/B 0.03fF
C14368 NAND2X1_LOC_184/Y INVX1_LOC_655/Y 0.01fF
C14369 INVX1_LOC_542/A INVX1_LOC_58/Y 0.03fF
C14370 INVX1_LOC_273/A INVX1_LOC_199/Y 0.00fF
C14371 VDD NAND2X1_LOC_409/Y 0.36fF
C14372 INVX1_LOC_269/A NAND2X1_LOC_91/a_36_24# 0.00fF
C14373 INVX1_LOC_452/A INVX1_LOC_385/Y 0.23fF
C14374 INVX1_LOC_7/Y INVX1_LOC_365/A 0.03fF
C14375 INVX1_LOC_53/Y INVX1_LOC_189/A 0.01fF
C14376 VDD INVX1_LOC_135/Y 0.21fF
C14377 INVX1_LOC_150/Y INVX1_LOC_498/Y 0.07fF
C14378 INPUT_0 INVX1_LOC_519/Y 0.03fF
C14379 NAND2X1_LOC_191/a_36_24# INVX1_LOC_197/A 0.00fF
C14380 INVX1_LOC_401/A NAND2X1_LOC_308/A 0.02fF
C14381 NAND2X1_LOC_635/B INVX1_LOC_632/A 0.11fF
C14382 INVX1_LOC_31/A NAND2X1_LOC_836/B 0.06fF
C14383 INVX1_LOC_323/Y INVX1_LOC_172/A 0.02fF
C14384 INVX1_LOC_53/Y NAND2X1_LOC_770/a_36_24# 0.00fF
C14385 INVX1_LOC_80/A INVX1_LOC_46/Y 0.03fF
C14386 INVX1_LOC_608/Y INVX1_LOC_213/Y 0.00fF
C14387 INVX1_LOC_546/Y NAND2X1_LOC_274/B 0.01fF
C14388 INVX1_LOC_438/A INVX1_LOC_62/Y 0.36fF
C14389 INVX1_LOC_269/A INVX1_LOC_245/A 0.01fF
C14390 INVX1_LOC_69/Y INVX1_LOC_495/A 0.94fF
C14391 INVX1_LOC_609/A NAND2X1_LOC_708/A 0.33fF
C14392 INVX1_LOC_213/Y INVX1_LOC_17/Y 0.72fF
C14393 INVX1_LOC_377/A INVX1_LOC_670/A 0.02fF
C14394 INVX1_LOC_211/A NAND2X1_LOC_76/B 0.00fF
C14395 NAND2X1_LOC_755/B NAND2X1_LOC_667/a_36_24# 0.00fF
C14396 NAND2X1_LOC_299/Y INVX1_LOC_89/Y 0.12fF
C14397 NAND2X1_LOC_756/Y INVX1_LOC_63/Y 0.09fF
C14398 INVX1_LOC_612/Y NAND2X1_LOC_697/Y 0.22fF
C14399 NAND2X1_LOC_830/a_36_24# INVX1_LOC_655/A -0.02fF
C14400 INVX1_LOC_392/Y NAND2X1_LOC_274/B 0.01fF
C14401 NAND2X1_LOC_56/Y INVX1_LOC_47/Y 0.00fF
C14402 INVX1_LOC_293/Y INVX1_LOC_63/Y 0.03fF
C14403 NAND2X1_LOC_710/B INVX1_LOC_479/A 0.00fF
C14404 INVX1_LOC_69/Y INVX1_LOC_633/Y 0.04fF
C14405 INPUT_5 INVX1_LOC_55/Y 0.13fF
C14406 INVX1_LOC_194/A INVX1_LOC_117/Y 0.02fF
C14407 INVX1_LOC_93/Y INVX1_LOC_549/Y 0.02fF
C14408 INVX1_LOC_492/A INVX1_LOC_54/Y 0.08fF
C14409 INVX1_LOC_229/Y INVX1_LOC_44/Y 0.06fF
C14410 NAND2X1_LOC_710/A INVX1_LOC_376/Y 0.03fF
C14411 INVX1_LOC_441/Y INVX1_LOC_62/Y 0.01fF
C14412 INVX1_LOC_20/Y INVX1_LOC_90/Y 0.33fF
C14413 INVX1_LOC_11/Y INVX1_LOC_46/Y 0.13fF
C14414 INVX1_LOC_193/A INVX1_LOC_103/Y 0.01fF
C14415 INVX1_LOC_668/A INVX1_LOC_655/A 0.04fF
C14416 VDD INVX1_LOC_76/A -0.00fF
C14417 INVX1_LOC_160/A INVX1_LOC_63/Y 0.03fF
C14418 INVX1_LOC_551/Y INVX1_LOC_319/A 0.04fF
C14419 INVX1_LOC_662/A NAND2X1_LOC_820/a_36_24# 0.01fF
C14420 NAND2X1_LOC_500/a_36_24# NAND2X1_LOC_521/Y 0.01fF
C14421 NAND2X1_LOC_619/Y INVX1_LOC_48/Y 0.01fF
C14422 NAND2X1_LOC_111/Y INVX1_LOC_116/Y 0.10fF
C14423 NAND2X1_LOC_693/a_36_24# INVX1_LOC_608/A 0.00fF
C14424 INVX1_LOC_17/Y NAND2X1_LOC_698/Y 0.04fF
C14425 NAND2X1_LOC_307/A NAND2X1_LOC_545/A 0.03fF
C14426 INVX1_LOC_145/Y INVX1_LOC_622/A 0.01fF
C14427 INVX1_LOC_44/Y NAND2X1_LOC_226/Y 0.05fF
C14428 INVX1_LOC_555/A INVX1_LOC_138/Y -0.01fF
C14429 INVX1_LOC_58/Y INVX1_LOC_259/Y 0.03fF
C14430 NAND2X1_LOC_673/B INVX1_LOC_63/Y 0.01fF
C14431 NAND2X1_LOC_115/a_36_24# INVX1_LOC_6/Y 0.00fF
C14432 INVX1_LOC_531/A INVX1_LOC_100/Y 0.03fF
C14433 NAND2X1_LOC_267/A INVX1_LOC_188/A 0.04fF
C14434 INVX1_LOC_614/A INVX1_LOC_135/Y 0.03fF
C14435 INVX1_LOC_300/A INVX1_LOC_90/Y 0.00fF
C14436 INVX1_LOC_242/Y INVX1_LOC_98/Y 0.10fF
C14437 NAND2X1_LOC_513/A INVX1_LOC_62/Y 0.17fF
C14438 INVX1_LOC_300/Y INVX1_LOC_673/Y 0.02fF
C14439 INVX1_LOC_379/A INVX1_LOC_79/A 0.08fF
C14440 INVX1_LOC_197/Y INVX1_LOC_90/Y 0.07fF
C14441 INVX1_LOC_655/A INVX1_LOC_668/Y 0.04fF
C14442 INVX1_LOC_392/A NAND2X1_LOC_274/B 0.03fF
C14443 INVX1_LOC_662/A INVX1_LOC_650/Y 0.02fF
C14444 INVX1_LOC_214/Y INVX1_LOC_100/Y 0.00fF
C14445 INVX1_LOC_327/Y INVX1_LOC_9/Y 0.06fF
C14446 INVX1_LOC_35/Y INVX1_LOC_79/A 0.13fF
C14447 INVX1_LOC_675/A INVX1_LOC_372/A 0.05fF
C14448 INVX1_LOC_35/Y NAND2X1_LOC_631/B 1.24fF
C14449 NAND2X1_LOC_846/A NAND2X1_LOC_846/B 0.05fF
C14450 INVX1_LOC_301/Y INVX1_LOC_66/A 4.16fF
C14451 INVX1_LOC_357/A INVX1_LOC_74/Y 0.03fF
C14452 INVX1_LOC_32/Y NAND2X1_LOC_436/a_36_24# 0.01fF
C14453 INVX1_LOC_93/Y NAND2X1_LOC_274/B 0.07fF
C14454 NAND2X1_LOC_121/Y INVX1_LOC_261/Y 0.15fF
C14455 INVX1_LOC_490/A INVX1_LOC_247/Y 0.01fF
C14456 INVX1_LOC_625/A INVX1_LOC_211/A 0.02fF
C14457 INVX1_LOC_41/Y NAND2X1_LOC_615/B 0.30fF
C14458 INVX1_LOC_592/Y INVX1_LOC_26/Y 0.00fF
C14459 INVX1_LOC_79/A INVX1_LOC_620/A 0.03fF
C14460 INVX1_LOC_554/A NAND2X1_LOC_711/a_36_24# 0.02fF
C14461 INVX1_LOC_99/Y INVX1_LOC_348/Y 0.05fF
C14462 INVX1_LOC_476/A INVX1_LOC_655/A 0.14fF
C14463 NAND2X1_LOC_137/A INVX1_LOC_680/A -0.00fF
C14464 INVX1_LOC_202/Y NAND2X1_LOC_231/B 0.04fF
C14465 INVX1_LOC_116/Y INVX1_LOC_363/A 0.01fF
C14466 NAND2X1_LOC_822/Y INVX1_LOC_635/Y 0.01fF
C14467 INVX1_LOC_58/Y INVX1_LOC_114/A 0.07fF
C14468 INVX1_LOC_41/Y INVX1_LOC_66/A 0.03fF
C14469 NAND2X1_LOC_388/A INVX1_LOC_62/Y 0.15fF
C14470 INVX1_LOC_49/Y INVX1_LOC_665/A 0.01fF
C14471 INVX1_LOC_89/Y INVX1_LOC_75/Y 0.07fF
C14472 NAND2X1_LOC_843/B NAND2X1_LOC_246/a_36_24# 0.00fF
C14473 INVX1_LOC_241/A INVX1_LOC_212/Y 0.01fF
C14474 INVX1_LOC_49/Y INVX1_LOC_505/Y 0.04fF
C14475 INVX1_LOC_50/Y NAND2X1_LOC_96/a_36_24# 0.00fF
C14476 INVX1_LOC_531/Y INVX1_LOC_179/A 0.07fF
C14477 INVX1_LOC_554/A INVX1_LOC_523/A 0.02fF
C14478 INVX1_LOC_47/Y INVX1_LOC_223/A 0.01fF
C14479 INVX1_LOC_211/A NAND2X1_LOC_52/Y 0.08fF
C14480 INVX1_LOC_405/A INVX1_LOC_45/Y 0.23fF
C14481 INVX1_LOC_177/Y VDD 0.21fF
C14482 NAND2X1_LOC_528/Y INVX1_LOC_26/Y 0.07fF
C14483 INVX1_LOC_519/A INVX1_LOC_109/Y 0.03fF
C14484 INVX1_LOC_193/Y INVX1_LOC_224/Y 0.03fF
C14485 INVX1_LOC_68/Y NAND2X1_LOC_754/a_36_24# 0.00fF
C14486 INVX1_LOC_463/A NAND2X1_LOC_707/A 0.07fF
C14487 INVX1_LOC_479/A INVX1_LOC_26/Y 0.10fF
C14488 INVX1_LOC_560/Y INVX1_LOC_45/Y 0.07fF
C14489 NAND2X1_LOC_45/Y INVX1_LOC_428/A 0.08fF
C14490 INVX1_LOC_446/A INVX1_LOC_293/Y 0.07fF
C14491 INVX1_LOC_100/Y INVX1_LOC_364/A 0.00fF
C14492 INVX1_LOC_193/Y INVX1_LOC_578/A 0.01fF
C14493 INVX1_LOC_562/A INVX1_LOC_586/A 0.01fF
C14494 INPUT_0 INVX1_LOC_65/Y 0.03fF
C14495 NAND2X1_LOC_271/B INVX1_LOC_586/A 0.05fF
C14496 NAND2X1_LOC_317/B INVX1_LOC_586/A 0.03fF
C14497 INVX1_LOC_119/Y INVX1_LOC_348/Y 0.52fF
C14498 INVX1_LOC_301/A NAND2X1_LOC_545/B 0.01fF
C14499 NAND2X1_LOC_789/B INVX1_LOC_191/A 0.01fF
C14500 NAND2X1_LOC_710/A INVX1_LOC_121/Y 0.24fF
C14501 INVX1_LOC_409/Y INVX1_LOC_469/A 0.01fF
C14502 NAND2X1_LOC_543/B NAND2X1_LOC_369/a_36_24# 0.02fF
C14503 VDD INVX1_LOC_344/Y 0.36fF
C14504 INVX1_LOC_558/A NAND2X1_LOC_704/B 0.17fF
C14505 INVX1_LOC_442/A NAND2X1_LOC_322/a_36_24# 0.00fF
C14506 INVX1_LOC_301/A INVX1_LOC_98/Y 0.03fF
C14507 INVX1_LOC_548/Y INVX1_LOC_80/A 0.03fF
C14508 INVX1_LOC_634/Y INVX1_LOC_625/Y 0.08fF
C14509 INVX1_LOC_206/Y INVX1_LOC_680/Y 0.15fF
C14510 INVX1_LOC_255/Y INVX1_LOC_372/Y 0.01fF
C14511 INVX1_LOC_437/Y VDD 0.20fF
C14512 INVX1_LOC_84/A INVX1_LOC_45/Y 0.10fF
C14513 INVX1_LOC_586/A INVX1_LOC_495/A 0.07fF
C14514 INVX1_LOC_307/Y NAND2X1_LOC_378/Y 0.14fF
C14515 NAND2X1_LOC_13/Y NAND2X1_LOC_493/B 0.02fF
C14516 NAND2X1_LOC_427/Y INVX1_LOC_356/A 0.13fF
C14517 INVX1_LOC_32/A INVX1_LOC_11/Y 0.02fF
C14518 VDD INVX1_LOC_221/Y 0.21fF
C14519 VDD NAND2X1_LOC_770/B 0.01fF
C14520 INVX1_LOC_564/A NAND2X1_LOC_755/B 0.05fF
C14521 INVX1_LOC_53/Y NAND2X1_LOC_122/Y 0.03fF
C14522 INVX1_LOC_435/Y NAND2X1_LOC_260/Y 0.03fF
C14523 INVX1_LOC_596/A NAND2X1_LOC_332/B 0.01fF
C14524 INVX1_LOC_312/Y NAND2X1_LOC_613/Y 0.01fF
C14525 INVX1_LOC_405/A NAND2X1_LOC_276/A 0.01fF
C14526 NAND2X1_LOC_318/A INVX1_LOC_80/A 0.06fF
C14527 INVX1_LOC_428/A INVX1_LOC_99/Y 0.03fF
C14528 INPUT_3 INVX1_LOC_84/A 0.30fF
C14529 NAND2X1_LOC_13/Y NAND2X1_LOC_336/B 0.00fF
C14530 INVX1_LOC_224/Y INVX1_LOC_54/Y 0.10fF
C14531 INVX1_LOC_11/Y INVX1_LOC_548/Y 0.01fF
C14532 INVX1_LOC_254/Y INVX1_LOC_560/A 0.07fF
C14533 NAND2X1_LOC_79/B INVX1_LOC_619/A 0.03fF
C14534 INVX1_LOC_45/Y NAND2X1_LOC_67/Y 0.01fF
C14535 NAND2X1_LOC_331/A INVX1_LOC_50/Y 0.67fF
C14536 INVX1_LOC_161/A INVX1_LOC_163/Y 0.03fF
C14537 INVX1_LOC_420/Y INVX1_LOC_421/A 0.00fF
C14538 INVX1_LOC_412/Y NAND2X1_LOC_453/a_36_24# 0.00fF
C14539 INVX1_LOC_578/A INVX1_LOC_54/Y 0.06fF
C14540 INPUT_2 INVX1_LOC_7/Y 0.08fF
C14541 NAND2X1_LOC_863/a_36_24# INVX1_LOC_602/Y 0.00fF
C14542 INVX1_LOC_20/Y INVX1_LOC_98/Y 0.01fF
C14543 NAND2X1_LOC_322/a_36_24# INVX1_LOC_116/Y 0.00fF
C14544 INVX1_LOC_206/Y INVX1_LOC_410/A 0.02fF
C14545 NAND2X1_LOC_521/Y NAND2X1_LOC_526/a_36_24# 0.00fF
C14546 INVX1_LOC_542/A NAND2X1_LOC_689/B 0.04fF
C14547 INVX1_LOC_80/A INVX1_LOC_363/Y 0.01fF
C14548 INVX1_LOC_596/A INVX1_LOC_503/Y 0.03fF
C14549 INVX1_LOC_99/Y INVX1_LOC_489/Y 0.03fF
C14550 VDD INVX1_LOC_373/Y 0.19fF
C14551 NAND2X1_LOC_88/B INVX1_LOC_177/A 0.03fF
C14552 INPUT_0 INVX1_LOC_314/Y 0.01fF
C14553 NAND2X1_LOC_362/a_36_24# INVX1_LOC_296/A 0.02fF
C14554 NAND2X1_LOC_333/A INVX1_LOC_577/Y 0.02fF
C14555 NAND2X1_LOC_704/B INVX1_LOC_46/Y 0.78fF
C14556 INVX1_LOC_551/Y INVX1_LOC_361/Y 0.10fF
C14557 INVX1_LOC_206/Y INVX1_LOC_399/Y 0.16fF
C14558 INVX1_LOC_202/Y INVX1_LOC_80/A 0.76fF
C14559 INVX1_LOC_547/Y INVX1_LOC_58/Y 0.07fF
C14560 NAND2X1_LOC_106/Y NAND2X1_LOC_692/a_36_24# 0.00fF
C14561 INVX1_LOC_317/Y INVX1_LOC_69/Y 0.04fF
C14562 INPUT_0 NAND2X1_LOC_813/a_36_24# 0.00fF
C14563 INVX1_LOC_434/A INVX1_LOC_100/Y 0.03fF
C14564 INVX1_LOC_501/Y INVX1_LOC_498/A 0.02fF
C14565 INVX1_LOC_686/A INVX1_LOC_354/Y 0.03fF
C14566 INVX1_LOC_417/Y INVX1_LOC_35/Y 0.05fF
C14567 INVX1_LOC_417/Y INVX1_LOC_304/A 0.04fF
C14568 INVX1_LOC_150/Y INVX1_LOC_513/Y 0.03fF
C14569 INVX1_LOC_499/Y INVX1_LOC_58/Y 0.21fF
C14570 INVX1_LOC_246/Y INVX1_LOC_490/A 0.02fF
C14571 INVX1_LOC_300/A INVX1_LOC_98/Y 0.01fF
C14572 NAND2X1_LOC_515/a_36_24# INVX1_LOC_89/Y 0.00fF
C14573 INVX1_LOC_340/A INVX1_LOC_59/A 0.06fF
C14574 INVX1_LOC_395/A NAND2X1_LOC_274/B 0.05fF
C14575 INVX1_LOC_297/A INVX1_LOC_32/Y 0.03fF
C14576 INVX1_LOC_398/Y INVX1_LOC_35/Y 0.01fF
C14577 INVX1_LOC_442/A INVX1_LOC_301/Y 0.29fF
C14578 INVX1_LOC_385/Y INVX1_LOC_282/A 0.03fF
C14579 NAND2X1_LOC_249/Y INVX1_LOC_479/A 0.03fF
C14580 INVX1_LOC_432/Y INVX1_LOC_211/Y 0.07fF
C14581 INVX1_LOC_490/Y INVX1_LOC_502/A 0.01fF
C14582 INVX1_LOC_35/Y INVX1_LOC_59/Y 0.03fF
C14583 INVX1_LOC_20/Y INVX1_LOC_338/Y 0.03fF
C14584 INVX1_LOC_238/A INVX1_LOC_479/A 0.01fF
C14585 INVX1_LOC_173/Y INVX1_LOC_174/A 0.01fF
C14586 INVX1_LOC_379/A INVX1_LOC_48/Y 0.07fF
C14587 NAND2X1_LOC_373/a_36_24# INVX1_LOC_479/A 0.01fF
C14588 INVX1_LOC_11/Y INVX1_LOC_202/Y 0.07fF
C14589 INVX1_LOC_362/Y NAND2X1_LOC_274/B 0.75fF
C14590 INVX1_LOC_468/Y INVX1_LOC_54/Y 0.03fF
C14591 INVX1_LOC_68/Y INVX1_LOC_353/A 0.13fF
C14592 INVX1_LOC_35/Y INVX1_LOC_48/Y 2.01fF
C14593 INVX1_LOC_72/Y INVX1_LOC_85/A 0.01fF
C14594 INVX1_LOC_58/Y INVX1_LOC_651/A 0.00fF
C14595 INVX1_LOC_432/Y INVX1_LOC_46/Y 0.05fF
C14596 INVX1_LOC_407/Y INVX1_LOC_50/Y 0.02fF
C14597 INPUT_0 INVX1_LOC_588/A 0.08fF
C14598 NAND2X1_LOC_400/B NAND2X1_LOC_393/Y 0.00fF
C14599 NAND2X1_LOC_336/B INVX1_LOC_361/A 0.25fF
C14600 INVX1_LOC_421/A NAND2X1_LOC_270/a_36_24# 0.00fF
C14601 INVX1_LOC_560/A INVX1_LOC_479/A 0.07fF
C14602 INVX1_LOC_21/Y INVX1_LOC_66/A 0.08fF
C14603 INVX1_LOC_80/A INVX1_LOC_49/Y 0.52fF
C14604 INVX1_LOC_352/Y NAND2X1_LOC_603/a_36_24# 0.01fF
C14605 INVX1_LOC_17/Y INVX1_LOC_561/A 0.01fF
C14606 INVX1_LOC_87/Y INVX1_LOC_178/A 0.11fF
C14607 INVX1_LOC_6/Y NAND2X1_LOC_397/Y 0.14fF
C14608 NAND2X1_LOC_517/a_36_24# INVX1_LOC_502/A 0.02fF
C14609 INVX1_LOC_442/A INVX1_LOC_41/Y 0.11fF
C14610 INVX1_LOC_117/Y INVX1_LOC_303/Y 0.03fF
C14611 INVX1_LOC_535/Y INVX1_LOC_137/Y 0.01fF
C14612 INPUT_1 INVX1_LOC_665/Y 0.06fF
C14613 INVX1_LOC_59/Y INVX1_LOC_620/A 0.01fF
C14614 INVX1_LOC_418/Y INVX1_LOC_93/Y 0.01fF
C14615 INVX1_LOC_93/Y INVX1_LOC_159/Y 1.00fF
C14616 INVX1_LOC_85/Y INVX1_LOC_184/Y 0.01fF
C14617 NAND2X1_LOC_531/Y INVX1_LOC_99/Y 0.09fF
C14618 NAND2X1_LOC_315/a_36_24# INVX1_LOC_100/Y 0.01fF
C14619 INVX1_LOC_54/Y NAND2X1_LOC_527/Y 0.08fF
C14620 INVX1_LOC_298/Y INVX1_LOC_261/Y 0.02fF
C14621 NAND2X1_LOC_274/B INVX1_LOC_683/Y 0.02fF
C14622 INVX1_LOC_469/Y INVX1_LOC_360/A 0.09fF
C14623 INVX1_LOC_204/Y INVX1_LOC_1/Y 0.06fF
C14624 INVX1_LOC_372/Y INVX1_LOC_26/Y 0.28fF
C14625 INVX1_LOC_11/Y INVX1_LOC_387/Y 0.04fF
C14626 INVX1_LOC_17/Y NAND2X1_LOC_258/Y 0.06fF
C14627 INVX1_LOC_270/A INVX1_LOC_319/A 0.03fF
C14628 INVX1_LOC_250/Y INVX1_LOC_353/A 0.12fF
C14629 NAND2X1_LOC_448/B INVX1_LOC_48/Y 0.01fF
C14630 INVX1_LOC_445/Y INVX1_LOC_443/A 0.03fF
C14631 INVX1_LOC_65/Y INVX1_LOC_211/A 0.07fF
C14632 INVX1_LOC_145/Y NAND2X1_LOC_52/Y 0.01fF
C14633 NAND2X1_LOC_445/a_36_24# INVX1_LOC_600/A 0.01fF
C14634 INVX1_LOC_65/Y INVX1_LOC_64/Y 0.08fF
C14635 INVX1_LOC_620/A INVX1_LOC_48/Y 0.51fF
C14636 INVX1_LOC_342/Y INVX1_LOC_659/A 0.03fF
C14637 NAND2X1_LOC_706/B INVX1_LOC_6/Y 0.19fF
C14638 NAND2X1_LOC_308/A INPUT_1 0.79fF
C14639 INVX1_LOC_98/A NAND2X1_LOC_231/B 0.10fF
C14640 NAND2X1_LOC_141/a_36_24# INVX1_LOC_361/Y 0.00fF
C14641 INVX1_LOC_21/Y INVX1_LOC_178/Y 0.01fF
C14642 INVX1_LOC_11/Y INVX1_LOC_49/Y 0.32fF
C14643 INVX1_LOC_588/Y INVX1_LOC_69/Y 0.06fF
C14644 NAND2X1_LOC_148/B INVX1_LOC_239/A 0.00fF
C14645 INVX1_LOC_301/Y INVX1_LOC_116/Y 0.01fF
C14646 NAND2X1_LOC_123/B INVX1_LOC_134/Y 0.07fF
C14647 INVX1_LOC_306/Y INVX1_LOC_117/Y 0.02fF
C14648 INVX1_LOC_76/Y NAND2X1_LOC_231/B 0.14fF
C14649 INVX1_LOC_166/A INVX1_LOC_69/Y 0.07fF
C14650 NAND2X1_LOC_636/B INVX1_LOC_62/Y 0.21fF
C14651 INVX1_LOC_598/A INVX1_LOC_622/A 0.02fF
C14652 INVX1_LOC_80/A INVX1_LOC_92/Y 0.01fF
C14653 INVX1_LOC_287/Y INVX1_LOC_91/Y 0.00fF
C14654 INVX1_LOC_338/A INVX1_LOC_79/A 0.00fF
C14655 INVX1_LOC_305/Y INVX1_LOC_41/Y 0.04fF
C14656 INVX1_LOC_17/Y NAND2X1_LOC_545/A 0.03fF
C14657 INVX1_LOC_245/A INVX1_LOC_259/Y 0.03fF
C14658 NAND2X1_LOC_111/Y INVX1_LOC_69/Y 0.03fF
C14659 INVX1_LOC_117/Y INVX1_LOC_9/Y 0.50fF
C14660 NAND2X1_LOC_846/A INVX1_LOC_199/Y 0.04fF
C14661 INVX1_LOC_41/Y INVX1_LOC_116/Y 0.11fF
C14662 INVX1_LOC_670/A INVX1_LOC_518/A 0.07fF
C14663 INVX1_LOC_115/Y INVX1_LOC_74/Y 0.13fF
C14664 INVX1_LOC_604/Y INVX1_LOC_211/A 0.65fF
C14665 INVX1_LOC_149/Y INVX1_LOC_139/Y 0.01fF
C14666 INVX1_LOC_31/Y NAND2X1_LOC_274/B 0.08fF
C14667 NAND2X1_LOC_333/A INVX1_LOC_26/Y 0.03fF
C14668 NAND2X1_LOC_521/Y INVX1_LOC_26/Y 0.33fF
C14669 INVX1_LOC_11/Y INVX1_LOC_92/Y 0.05fF
C14670 INVX1_LOC_513/Y INVX1_LOC_501/A 0.80fF
C14671 NAND2X1_LOC_755/B INVX1_LOC_91/Y 0.01fF
C14672 INVX1_LOC_134/Y INVX1_LOC_92/A 0.07fF
C14673 INVX1_LOC_117/Y INVX1_LOC_62/Y 4.13fF
C14674 INVX1_LOC_479/Y INVX1_LOC_211/A 0.01fF
C14675 INVX1_LOC_26/Y INVX1_LOC_188/A 0.15fF
C14676 NAND2X1_LOC_433/Y INVX1_LOC_49/Y 0.22fF
C14677 INVX1_LOC_89/Y NAND2X1_LOC_441/a_36_24# 0.01fF
C14678 INVX1_LOC_117/Y INVX1_LOC_13/Y 0.22fF
C14679 INVX1_LOC_451/A INVX1_LOC_443/Y 0.00fF
C14680 NAND2X1_LOC_843/B INVX1_LOC_46/Y 0.01fF
C14681 INVX1_LOC_499/A NAND2X1_LOC_639/a_36_24# 0.02fF
C14682 INVX1_LOC_69/Y INVX1_LOC_531/Y 0.16fF
C14683 NAND2X1_LOC_409/Y INVX1_LOC_145/A 0.18fF
C14684 INVX1_LOC_318/A INVX1_LOC_211/A 0.00fF
C14685 INVX1_LOC_255/A INVX1_LOC_41/Y 0.03fF
C14686 NAND2X1_LOC_440/A INVX1_LOC_114/A 0.03fF
C14687 NAND2X1_LOC_274/B INVX1_LOC_128/A 0.22fF
C14688 INVX1_LOC_114/A INVX1_LOC_245/A 0.03fF
C14689 INVX1_LOC_397/Y INVX1_LOC_211/A 0.03fF
C14690 INVX1_LOC_100/Y INVX1_LOC_667/Y -0.00fF
C14691 INVX1_LOC_30/Y VDD 0.26fF
C14692 NAND2X1_LOC_475/A NAND2X1_LOC_75/a_36_24# 0.00fF
C14693 INVX1_LOC_179/A INVX1_LOC_41/Y 0.03fF
C14694 VDD INVX1_LOC_584/A 0.15fF
C14695 INVX1_LOC_31/Y NAND2X1_LOC_449/a_36_24# 0.00fF
C14696 INVX1_LOC_47/Y NAND2X1_LOC_832/A 0.10fF
C14697 INVX1_LOC_69/Y INVX1_LOC_363/A 0.01fF
C14698 INVX1_LOC_404/Y INVX1_LOC_438/A 0.02fF
C14699 NAND2X1_LOC_67/a_36_24# INVX1_LOC_169/A 0.00fF
C14700 VDD INVX1_LOC_400/Y 0.44fF
C14701 NAND2X1_LOC_636/A INVX1_LOC_167/Y 0.02fF
C14702 INVX1_LOC_65/A INVX1_LOC_92/A 0.09fF
C14703 INVX1_LOC_133/Y NAND2X1_LOC_820/A 0.00fF
C14704 INVX1_LOC_237/Y INVX1_LOC_395/A 0.05fF
C14705 INVX1_LOC_119/Y NAND2X1_LOC_832/A 0.09fF
C14706 NAND2X1_LOC_791/B NAND2X1_LOC_759/B 0.03fF
C14707 NAND2X1_LOC_66/Y INVX1_LOC_443/A 0.05fF
C14708 INVX1_LOC_38/A INVX1_LOC_395/A 0.08fF
C14709 NAND2X1_LOC_98/a_36_24# INVX1_LOC_524/Y 0.00fF
C14710 INVX1_LOC_426/Y INVX1_LOC_12/Y 0.09fF
C14711 INVX1_LOC_445/Y NAND2X1_LOC_261/Y 0.23fF
C14712 INVX1_LOC_206/Y NAND2X1_LOC_176/a_36_24# 0.00fF
C14713 VDD INVX1_LOC_514/Y 0.21fF
C14714 INVX1_LOC_193/Y INVX1_LOC_686/A 0.00fF
C14715 NAND2X1_LOC_788/A INVX1_LOC_21/Y 0.01fF
C14716 INVX1_LOC_560/Y INVX1_LOC_160/A 0.65fF
C14717 NAND2X1_LOC_636/A INVX1_LOC_137/Y 0.05fF
C14718 NAND2X1_LOC_534/Y INVX1_LOC_468/Y 0.01fF
C14719 VDD INVX1_LOC_55/A -0.00fF
C14720 INVX1_LOC_50/Y INVX1_LOC_638/A 0.07fF
C14721 INPUT_0 INVX1_LOC_670/Y 0.07fF
C14722 VDD INVX1_LOC_125/A -0.00fF
C14723 INVX1_LOC_53/Y INVX1_LOC_523/A 0.23fF
C14724 INVX1_LOC_627/A INVX1_LOC_6/Y 0.07fF
C14725 INVX1_LOC_420/Y INVX1_LOC_99/Y 0.04fF
C14726 INVX1_LOC_133/Y INVX1_LOC_6/Y 0.09fF
C14727 INVX1_LOC_68/Y INVX1_LOC_250/Y 0.10fF
C14728 INVX1_LOC_80/A INVX1_LOC_98/A 0.00fF
C14729 INVX1_LOC_17/Y INVX1_LOC_490/Y 0.28fF
C14730 INVX1_LOC_21/Y INVX1_LOC_442/A 0.07fF
C14731 INVX1_LOC_80/A INVX1_LOC_76/Y 1.29fF
C14732 INVX1_LOC_20/Y INVX1_LOC_596/A 0.00fF
C14733 INVX1_LOC_206/Y INVX1_LOC_54/Y 0.24fF
C14734 INPUT_0 NAND2X1_LOC_646/A 0.03fF
C14735 VDD INVX1_LOC_496/Y 0.45fF
C14736 INVX1_LOC_206/Y NAND2X1_LOC_614/a_36_24# 0.00fF
C14737 INVX1_LOC_68/Y INVX1_LOC_600/A 0.01fF
C14738 INVX1_LOC_418/Y INVX1_LOC_395/A 0.40fF
C14739 INVX1_LOC_683/A INVX1_LOC_51/Y 0.01fF
C14740 VDD INVX1_LOC_84/Y 0.12fF
C14741 INVX1_LOC_85/Y INVX1_LOC_7/Y 0.00fF
C14742 INVX1_LOC_65/Y INVX1_LOC_145/Y 0.15fF
C14743 INVX1_LOC_395/A INVX1_LOC_159/Y 0.13fF
C14744 INVX1_LOC_425/A INVX1_LOC_130/Y 0.06fF
C14745 INPUT_0 INVX1_LOC_86/Y 0.17fF
C14746 NAND2X1_LOC_498/Y INVX1_LOC_371/A 0.01fF
C14747 NAND2X1_LOC_184/a_36_24# INVX1_LOC_6/Y -0.00fF
C14748 INVX1_LOC_492/A INVX1_LOC_137/A 0.01fF
C14749 INVX1_LOC_11/Y NAND2X1_LOC_498/B 0.16fF
C14750 INVX1_LOC_307/Y INVX1_LOC_6/Y 0.01fF
C14751 NAND2X1_LOC_173/Y INVX1_LOC_99/Y 0.00fF
C14752 INVX1_LOC_11/Y INVX1_LOC_98/A 0.02fF
C14753 NAND2X1_LOC_475/A INVX1_LOC_187/Y 0.01fF
C14754 INVX1_LOC_224/Y INVX1_LOC_89/Y 0.82fF
C14755 NAND2X1_LOC_750/Y INVX1_LOC_47/Y 0.00fF
C14756 INVX1_LOC_20/Y INVX1_LOC_504/A 0.07fF
C14757 INVX1_LOC_224/Y INVX1_LOC_154/A 0.01fF
C14758 NAND2X1_LOC_333/A INVX1_LOC_564/Y 0.01fF
C14759 INVX1_LOC_588/Y INVX1_LOC_586/A 0.03fF
C14760 INVX1_LOC_107/A NAND2X1_LOC_285/A 0.30fF
C14761 INVX1_LOC_12/Y INVX1_LOC_369/A 0.03fF
C14762 INVX1_LOC_11/Y INVX1_LOC_76/Y 0.31fF
C14763 INVX1_LOC_291/A INVX1_LOC_59/Y 0.01fF
C14764 INVX1_LOC_54/Y INVX1_LOC_143/Y 0.04fF
C14765 INVX1_LOC_526/A INVX1_LOC_637/A 0.15fF
C14766 INVX1_LOC_395/A INVX1_LOC_212/Y 0.29fF
C14767 INVX1_LOC_578/A INVX1_LOC_89/Y 0.14fF
C14768 INVX1_LOC_557/A INVX1_LOC_89/Y 0.21fF
C14769 INVX1_LOC_166/A INVX1_LOC_586/A 0.01fF
C14770 INPUT_0 INVX1_LOC_63/Y 2.53fF
C14771 INVX1_LOC_564/A INVX1_LOC_49/Y 0.01fF
C14772 INVX1_LOC_224/Y INVX1_LOC_501/A -0.00fF
C14773 INVX1_LOC_242/Y NAND2X1_LOC_76/B 0.02fF
C14774 INVX1_LOC_291/A INVX1_LOC_48/Y 0.07fF
C14775 INVX1_LOC_21/Y INVX1_LOC_305/Y 0.01fF
C14776 INVX1_LOC_84/A NAND2X1_LOC_673/B 0.03fF
C14777 NAND2X1_LOC_702/a_36_24# INVX1_LOC_367/A 0.00fF
C14778 INVX1_LOC_578/A NAND2X1_LOC_319/a_36_24# 0.00fF
C14779 INVX1_LOC_287/Y NAND2X1_LOC_333/B 0.02fF
C14780 INVX1_LOC_278/A INVX1_LOC_386/A 0.30fF
C14781 NAND2X1_LOC_24/a_36_24# INVX1_LOC_63/Y 0.00fF
C14782 INVX1_LOC_361/Y INVX1_LOC_270/A 0.12fF
C14783 INVX1_LOC_54/Y INVX1_LOC_686/A 0.09fF
C14784 INVX1_LOC_447/A INVX1_LOC_100/Y 0.00fF
C14785 NAND2X1_LOC_538/B INVX1_LOC_31/Y 0.06fF
C14786 INVX1_LOC_21/Y INVX1_LOC_116/Y 0.03fF
C14787 INVX1_LOC_587/Y INVX1_LOC_658/A 0.01fF
C14788 INVX1_LOC_169/A INVX1_LOC_6/Y 0.05fF
C14789 INVX1_LOC_661/A INVX1_LOC_283/A 0.32fF
C14790 INVX1_LOC_134/Y INPUT_1 2.00fF
C14791 INVX1_LOC_312/Y INVX1_LOC_166/A 0.03fF
C14792 INVX1_LOC_604/A INVX1_LOC_26/Y 0.01fF
C14793 INVX1_LOC_609/Y INVX1_LOC_54/Y 0.01fF
C14794 INVX1_LOC_412/Y NAND2X1_LOC_109/a_36_24# 0.00fF
C14795 INVX1_LOC_397/A INVX1_LOC_399/Y 0.00fF
C14796 INVX1_LOC_435/Y INVX1_LOC_655/A 0.10fF
C14797 INVX1_LOC_6/Y INVX1_LOC_337/Y 0.03fF
C14798 NAND2X1_LOC_685/B INVX1_LOC_498/Y 0.04fF
C14799 NAND2X1_LOC_134/a_36_24# INVX1_LOC_124/A 0.00fF
C14800 INVX1_LOC_17/Y INVX1_LOC_391/Y 0.02fF
C14801 INVX1_LOC_531/A INVX1_LOC_48/Y 0.02fF
C14802 INVX1_LOC_565/A INVX1_LOC_674/A 0.04fF
C14803 INVX1_LOC_367/A NAND2X1_LOC_225/a_36_24# -0.02fF
C14804 NAND2X1_LOC_673/B NAND2X1_LOC_67/Y 0.05fF
C14805 NAND2X1_LOC_498/B NAND2X1_LOC_433/Y 0.10fF
C14806 NAND2X1_LOC_308/a_36_24# INVX1_LOC_252/A 0.02fF
C14807 INVX1_LOC_257/A INVX1_LOC_686/A 0.10fF
C14808 INVX1_LOC_566/Y INVX1_LOC_49/Y 0.03fF
C14809 INVX1_LOC_581/A INVX1_LOC_6/Y 0.42fF
C14810 INVX1_LOC_54/Y INVX1_LOC_14/A 0.01fF
C14811 INVX1_LOC_17/Y INVX1_LOC_431/A 0.05fF
C14812 NAND2X1_LOC_274/B NAND2X1_LOC_794/a_36_24# 0.00fF
C14813 INVX1_LOC_218/Y INVX1_LOC_453/Y 0.04fF
C14814 NAND2X1_LOC_755/B NAND2X1_LOC_333/B 0.03fF
C14815 INVX1_LOC_51/Y NAND2X1_LOC_274/B 0.03fF
C14816 INVX1_LOC_396/A INVX1_LOC_35/Y 0.01fF
C14817 NAND2X1_LOC_152/a_36_24# INVX1_LOC_6/Y 0.00fF
C14818 INVX1_LOC_378/A INVX1_LOC_245/A 0.01fF
C14819 INVX1_LOC_482/A INVX1_LOC_245/A 0.00fF
C14820 INVX1_LOC_76/Y NAND2X1_LOC_433/Y 0.69fF
C14821 INVX1_LOC_117/Y INVX1_LOC_42/Y 0.00fF
C14822 INVX1_LOC_318/A INVX1_LOC_145/Y 0.00fF
C14823 INVX1_LOC_373/A INVX1_LOC_479/A 0.03fF
C14824 INVX1_LOC_492/Y INVX1_LOC_168/Y 0.00fF
C14825 NAND2X1_LOC_454/a_36_24# INVX1_LOC_440/Y 0.00fF
C14826 INVX1_LOC_544/A NAND2X1_LOC_137/A 0.00fF
C14827 INVX1_LOC_50/Y INVX1_LOC_665/Y 0.06fF
C14828 INVX1_LOC_395/A INVX1_LOC_39/Y 0.03fF
C14829 INVX1_LOC_387/Y INVX1_LOC_367/Y 0.47fF
C14830 INVX1_LOC_21/Y INVX1_LOC_255/A 0.07fF
C14831 INVX1_LOC_468/Y INVX1_LOC_89/Y 0.04fF
C14832 INVX1_LOC_608/A INVX1_LOC_303/Y 0.10fF
C14833 INVX1_LOC_586/A INVX1_LOC_531/Y 0.06fF
C14834 INVX1_LOC_93/Y INVX1_LOC_352/Y 0.02fF
C14835 INVX1_LOC_31/Y INVX1_LOC_159/Y 0.07fF
C14836 NAND2X1_LOC_567/a_36_24# INVX1_LOC_634/Y 0.00fF
C14837 NAND2X1_LOC_376/B NAND2X1_LOC_376/Y 0.00fF
C14838 NAND2X1_LOC_188/a_36_24# INVX1_LOC_74/Y 0.00fF
C14839 INVX1_LOC_649/Y INVX1_LOC_644/Y 0.02fF
C14840 INVX1_LOC_197/A INVX1_LOC_491/A 0.14fF
C14841 INVX1_LOC_31/A NAND2X1_LOC_409/Y 0.01fF
C14842 INVX1_LOC_361/Y INVX1_LOC_46/Y 0.03fF
C14843 INVX1_LOC_49/Y INVX1_LOC_367/Y 0.07fF
C14844 INVX1_LOC_335/Y NAND2X1_LOC_719/A 0.00fF
C14845 INVX1_LOC_607/Y INVX1_LOC_63/Y 0.11fF
C14846 INVX1_LOC_105/Y INVX1_LOC_670/A 0.00fF
C14847 INVX1_LOC_47/Y INVX1_LOC_371/A 0.11fF
C14848 INVX1_LOC_201/A INVX1_LOC_63/Y 0.01fF
C14849 INVX1_LOC_21/Y INVX1_LOC_179/A 0.00fF
C14850 NAND2X1_LOC_528/Y INVX1_LOC_235/Y 0.27fF
C14851 NAND2X1_LOC_57/Y INVX1_LOC_223/Y 0.01fF
C14852 INVX1_LOC_586/A NAND2X1_LOC_626/a_36_24# 0.00fF
C14853 INVX1_LOC_435/A INVX1_LOC_328/Y 0.03fF
C14854 INVX1_LOC_466/A INVX1_LOC_69/Y 0.00fF
C14855 INVX1_LOC_65/A INPUT_1 0.28fF
C14856 INVX1_LOC_178/A INVX1_LOC_9/Y 0.07fF
C14857 INVX1_LOC_625/A INVX1_LOC_242/Y 0.02fF
C14858 INVX1_LOC_662/A NAND2X1_LOC_288/a_36_24# 0.01fF
C14859 INVX1_LOC_194/A INVX1_LOC_245/A 0.00fF
C14860 INVX1_LOC_340/Y INVX1_LOC_462/Y 0.01fF
C14861 INVX1_LOC_268/Y INVX1_LOC_91/Y 0.23fF
C14862 INVX1_LOC_49/Y INVX1_LOC_374/Y 0.01fF
C14863 INVX1_LOC_17/Y NAND2X1_LOC_489/A -0.06fF
C14864 INVX1_LOC_641/A INVX1_LOC_340/A 0.23fF
C14865 INVX1_LOC_99/Y NAND2X1_LOC_488/Y 0.01fF
C14866 INVX1_LOC_411/A INVX1_LOC_100/Y 0.03fF
C14867 INVX1_LOC_25/Y INVX1_LOC_25/A 0.01fF
C14868 INVX1_LOC_77/Y INVX1_LOC_361/A 0.06fF
C14869 INVX1_LOC_592/Y NAND2X1_LOC_420/Y 0.05fF
C14870 INVX1_LOC_556/Y INVX1_LOC_479/A 2.43fF
C14871 INVX1_LOC_338/Y INVX1_LOC_494/Y 0.02fF
C14872 INVX1_LOC_301/Y INVX1_LOC_69/Y 0.04fF
C14873 INVX1_LOC_58/Y INVX1_LOC_9/Y 0.29fF
C14874 INVX1_LOC_608/A INVX1_LOC_62/Y 0.03fF
C14875 INVX1_LOC_261/A INVX1_LOC_659/A 0.21fF
C14876 INVX1_LOC_202/Y INVX1_LOC_91/Y 0.26fF
C14877 NAND2X1_LOC_90/a_36_24# INVX1_LOC_9/Y 0.00fF
C14878 INVX1_LOC_430/A NAND2X1_LOC_344/B 0.11fF
C14879 INVX1_LOC_361/Y INVX1_LOC_75/A 0.01fF
C14880 INVX1_LOC_170/A NAND2X1_LOC_626/Y 0.02fF
C14881 INVX1_LOC_352/A NAND2X1_LOC_418/a_36_24# 0.00fF
C14882 INVX1_LOC_69/Y INVX1_LOC_41/Y 11.59fF
C14883 INVX1_LOC_48/Y INVX1_LOC_488/Y 0.11fF
C14884 NAND2X1_LOC_557/B NAND2X1_LOC_488/Y 0.08fF
C14885 INVX1_LOC_32/Y NAND2X1_LOC_231/B 0.15fF
C14886 INVX1_LOC_446/A INPUT_0 0.07fF
C14887 VDD INVX1_LOC_19/Y 0.21fF
C14888 INVX1_LOC_62/Y INVX1_LOC_58/Y 0.17fF
C14889 VDD NAND2X1_LOC_45/Y 2.03fF
C14890 NAND2X1_LOC_391/B INVX1_LOC_109/Y 0.03fF
C14891 INVX1_LOC_141/Y INVX1_LOC_588/A 0.02fF
C14892 INVX1_LOC_62/Y NAND2X1_LOC_636/a_36_24# 0.00fF
C14893 INVX1_LOC_224/Y INVX1_LOC_203/Y 0.01fF
C14894 INVX1_LOC_63/Y INVX1_LOC_211/A 0.03fF
C14895 VDD INVX1_LOC_445/Y 0.28fF
C14896 INVX1_LOC_63/Y INVX1_LOC_64/Y 0.18fF
C14897 VDD INVX1_LOC_36/A -0.00fF
C14898 INVX1_LOC_49/Y INVX1_LOC_91/Y 0.01fF
C14899 VDD INVX1_LOC_570/A 0.13fF
C14900 NAND2X1_LOC_597/Y INVX1_LOC_114/A 0.01fF
C14901 INVX1_LOC_193/Y INVX1_LOC_390/Y 0.04fF
C14902 INVX1_LOC_192/Y INVX1_LOC_560/A 0.06fF
C14903 INPUT_0 INVX1_LOC_552/Y 0.01fF
C14904 INVX1_LOC_476/A INVX1_LOC_92/A 0.18fF
C14905 INPUT_0 NAND2X1_LOC_691/a_36_24# 0.00fF
C14906 INVX1_LOC_20/Y NAND2X1_LOC_76/B 0.40fF
C14907 INVX1_LOC_629/Y NAND2X1_LOC_122/Y 0.01fF
C14908 VDD INVX1_LOC_377/Y 0.41fF
C14909 INVX1_LOC_442/A INVX1_LOC_255/Y 0.01fF
C14910 INVX1_LOC_485/A INVX1_LOC_90/Y 0.01fF
C14911 NAND2X1_LOC_498/Y INVX1_LOC_383/A 0.01fF
C14912 INVX1_LOC_73/Y INVX1_LOC_366/Y 0.06fF
C14913 INVX1_LOC_319/Y INVX1_LOC_76/Y 0.03fF
C14914 INVX1_LOC_570/A INVX1_LOC_510/Y 0.07fF
C14915 INVX1_LOC_555/Y INVX1_LOC_523/A 0.04fF
C14916 INVX1_LOC_551/Y INVX1_LOC_412/A 0.10fF
C14917 VDD INVX1_LOC_676/Y 0.58fF
C14918 INVX1_LOC_85/Y INVX1_LOC_616/A 0.01fF
C14919 VDD INVX1_LOC_99/Y 2.61fF
C14920 INVX1_LOC_300/A NAND2X1_LOC_76/B 0.46fF
C14921 INVX1_LOC_426/A INVX1_LOC_159/Y 0.01fF
C14922 VDD INVX1_LOC_609/A 0.01fF
C14923 NAND2X1_LOC_467/A INVX1_LOC_586/A 0.01fF
C14924 INVX1_LOC_383/A INVX1_LOC_377/Y 0.01fF
C14925 NAND2X1_LOC_88/B INVX1_LOC_65/Y 0.31fF
C14926 INVX1_LOC_438/A INVX1_LOC_451/A 0.10fF
C14927 INVX1_LOC_614/A INVX1_LOC_570/A 0.39fF
C14928 INVX1_LOC_438/Y INVX1_LOC_444/Y 0.03fF
C14929 NAND2X1_LOC_583/a_36_24# INVX1_LOC_54/Y 0.01fF
C14930 INVX1_LOC_113/Y INVX1_LOC_686/A 0.03fF
C14931 NAND2X1_LOC_307/A INVX1_LOC_624/A 0.07fF
C14932 NAND2X1_LOC_79/B NAND2X1_LOC_773/A 0.02fF
C14933 INVX1_LOC_228/Y INVX1_LOC_99/Y 0.02fF
C14934 INVX1_LOC_449/A INVX1_LOC_392/Y 0.00fF
C14935 INVX1_LOC_167/Y INVX1_LOC_492/Y 0.09fF
C14936 INVX1_LOC_203/Y INVX1_LOC_227/Y 0.01fF
C14937 NAND2X1_LOC_218/a_36_24# INVX1_LOC_230/A 0.00fF
C14938 VDD INVX1_LOC_123/A 0.00fF
C14939 INVX1_LOC_143/Y NAND2X1_LOC_677/Y 0.01fF
C14940 INVX1_LOC_276/A INVX1_LOC_80/A 0.01fF
C14941 INVX1_LOC_255/Y INVX1_LOC_116/Y 0.00fF
C14942 NAND2X1_LOC_45/Y INVX1_LOC_103/Y 0.03fF
C14943 INVX1_LOC_429/Y INVX1_LOC_453/Y 0.44fF
C14944 INVX1_LOC_362/Y NAND2X1_LOC_595/Y 0.06fF
C14945 INVX1_LOC_453/A NAND2X1_LOC_294/Y 0.01fF
C14946 VDD INVX1_LOC_589/Y 0.21fF
C14947 NAND2X1_LOC_336/B INVX1_LOC_551/Y 0.06fF
C14948 NAND2X1_LOC_249/Y INVX1_LOC_66/A 0.03fF
C14949 VDD INVX1_LOC_568/A 0.00fF
C14950 INVX1_LOC_459/A INVX1_LOC_376/A 0.01fF
C14951 NAND2X1_LOC_498/Y INVX1_LOC_509/A 0.01fF
C14952 INVX1_LOC_409/A INVX1_LOC_31/Y 0.07fF
C14953 NAND2X1_LOC_331/A INVX1_LOC_117/Y 0.12fF
C14954 VDD INVX1_LOC_47/Y 2.32fF
C14955 NAND2X1_LOC_789/a_36_24# INVX1_LOC_191/A 0.00fF
C14956 NAND2X1_LOC_39/Y INVX1_LOC_53/Y 0.03fF
C14957 INVX1_LOC_12/Y INVX1_LOC_235/Y 0.03fF
C14958 INVX1_LOC_179/Y NAND2X1_LOC_86/Y 0.00fF
C14959 VDD NAND2X1_LOC_557/B 1.12fF
C14960 INVX1_LOC_206/Y INVX1_LOC_199/A 0.01fF
C14961 INVX1_LOC_618/A NAND2X1_LOC_274/B 0.21fF
C14962 INVX1_LOC_206/Y INVX1_LOC_89/Y 0.09fF
C14963 INVX1_LOC_432/Y INVX1_LOC_76/Y 0.04fF
C14964 INVX1_LOC_228/Y INVX1_LOC_123/A 0.04fF
C14965 INVX1_LOC_683/Y INVX1_LOC_377/A 0.41fF
C14966 INVX1_LOC_381/A NAND2X1_LOC_415/B 0.08fF
C14967 INVX1_LOC_76/Y INVX1_LOC_367/Y 0.12fF
C14968 INVX1_LOC_20/Y INVX1_LOC_625/A 0.02fF
C14969 INVX1_LOC_51/Y INVX1_LOC_159/Y 0.00fF
C14970 INVX1_LOC_584/Y INVX1_LOC_93/Y 0.00fF
C14971 INVX1_LOC_556/A NAND2X1_LOC_128/A 0.01fF
C14972 NAND2X1_LOC_596/Y INVX1_LOC_47/Y 0.02fF
C14973 INVX1_LOC_333/Y INVX1_LOC_602/A 0.04fF
C14974 NAND2X1_LOC_56/Y INVX1_LOC_600/A 0.01fF
C14975 NAND2X1_LOC_311/a_36_24# INVX1_LOC_230/A 0.01fF
C14976 INVX1_LOC_228/Y INVX1_LOC_47/Y 0.02fF
C14977 NAND2X1_LOC_707/A INVX1_LOC_493/A 0.03fF
C14978 INVX1_LOC_193/Y NAND2X1_LOC_542/A 0.01fF
C14979 INVX1_LOC_53/Y NAND2X1_LOC_147/B 0.01fF
C14980 INVX1_LOC_257/Y INVX1_LOC_63/Y 0.07fF
C14981 INVX1_LOC_609/Y NAND2X1_LOC_677/Y 0.01fF
C14982 INVX1_LOC_266/A INVX1_LOC_418/Y 0.02fF
C14983 NAND2X1_LOC_865/a_36_24# INVX1_LOC_116/Y 0.00fF
C14984 INVX1_LOC_266/A INVX1_LOC_159/Y 0.10fF
C14985 INVX1_LOC_206/Y INVX1_LOC_501/A 3.53fF
C14986 INVX1_LOC_35/Y INVX1_LOC_508/Y 0.01fF
C14987 INVX1_LOC_393/Y INVX1_LOC_49/Y 0.02fF
C14988 INVX1_LOC_197/A INVX1_LOC_504/Y 0.07fF
C14989 INVX1_LOC_256/A INVX1_LOC_80/A 0.01fF
C14990 INVX1_LOC_561/A NAND2X1_LOC_122/Y 0.03fF
C14991 INVX1_LOC_137/Y INVX1_LOC_492/Y 0.05fF
C14992 INVX1_LOC_446/Y INVX1_LOC_63/Y 0.07fF
C14993 VDD INVX1_LOC_119/Y 0.75fF
C14994 INVX1_LOC_628/A NAND2X1_LOC_448/A 0.04fF
C14995 INVX1_LOC_510/Y NAND2X1_LOC_306/a_36_24# 0.00fF
C14996 VDD NAND2X1_LOC_66/Y 0.70fF
C14997 INVX1_LOC_515/A NAND2X1_LOC_829/B 0.01fF
C14998 INVX1_LOC_510/Y INVX1_LOC_47/Y 1.39fF
C14999 INVX1_LOC_449/A INVX1_LOC_392/A 0.01fF
C15000 INVX1_LOC_89/Y INVX1_LOC_242/A 0.03fF
C15001 INVX1_LOC_126/Y INVX1_LOC_670/A 0.02fF
C15002 INVX1_LOC_287/A INVX1_LOC_440/A 0.01fF
C15003 INVX1_LOC_625/A INVX1_LOC_300/A 0.04fF
C15004 INVX1_LOC_53/Y INVX1_LOC_513/A 0.06fF
C15005 INVX1_LOC_523/A INVX1_LOC_662/A 0.07fF
C15006 INVX1_LOC_583/Y INVX1_LOC_168/Y 0.04fF
C15007 INVX1_LOC_80/A INVX1_LOC_345/Y 0.00fF
C15008 NAND2X1_LOC_131/a_36_24# INVX1_LOC_35/Y 0.00fF
C15009 NAND2X1_LOC_596/Y INVX1_LOC_119/Y 0.00fF
C15010 INVX1_LOC_134/Y INVX1_LOC_50/Y 3.54fF
C15011 INVX1_LOC_586/A INVX1_LOC_411/Y 0.02fF
C15012 INVX1_LOC_11/Y NAND2X1_LOC_399/B 0.12fF
C15013 NAND2X1_LOC_111/a_36_24# INVX1_LOC_686/A 0.01fF
C15014 NAND2X1_LOC_48/Y INVX1_LOC_50/Y 0.02fF
C15015 INVX1_LOC_11/Y INVX1_LOC_7/Y 1.61fF
C15016 INVX1_LOC_89/Y INVX1_LOC_686/A 0.25fF
C15017 INVX1_LOC_384/A INVX1_LOC_63/Y 0.07fF
C15018 NAND2X1_LOC_250/Y INVX1_LOC_145/Y 0.01fF
C15019 INVX1_LOC_80/A INVX1_LOC_32/Y 0.10fF
C15020 INVX1_LOC_579/Y INVX1_LOC_32/Y 0.03fF
C15021 INVX1_LOC_449/A INVX1_LOC_93/Y 0.07fF
C15022 INVX1_LOC_20/Y NAND2X1_LOC_52/Y 0.33fF
C15023 NAND2X1_LOC_669/Y INVX1_LOC_93/Y 0.01fF
C15024 INVX1_LOC_65/Y INVX1_LOC_242/Y 0.15fF
C15025 INVX1_LOC_99/Y NAND2X1_LOC_607/a_36_24# 0.00fF
C15026 INVX1_LOC_11/Y NAND2X1_LOC_259/A 0.02fF
C15027 INVX1_LOC_370/Y INPUT_1 0.02fF
C15028 INVX1_LOC_444/Y INVX1_LOC_219/Y 0.02fF
C15029 INVX1_LOC_307/A INVX1_LOC_46/Y 0.39fF
C15030 INVX1_LOC_614/A INVX1_LOC_568/A 0.01fF
C15031 INVX1_LOC_167/Y INVX1_LOC_168/Y 0.96fF
C15032 NAND2X1_LOC_390/a_36_24# INVX1_LOC_9/Y 0.00fF
C15033 INVX1_LOC_442/A INVX1_LOC_128/Y 0.02fF
C15034 INVX1_LOC_145/Y INVX1_LOC_623/Y 0.02fF
C15035 INVX1_LOC_401/A INVX1_LOC_338/Y 0.01fF
C15036 INVX1_LOC_45/Y INVX1_LOC_373/Y 0.00fF
C15037 INVX1_LOC_145/Y INVX1_LOC_86/Y 1.45fF
C15038 INVX1_LOC_383/A INVX1_LOC_119/Y 0.01fF
C15039 INVX1_LOC_173/A INVX1_LOC_100/Y 0.03fF
C15040 NAND2X1_LOC_448/B INVX1_LOC_155/Y 0.01fF
C15041 INVX1_LOC_442/Y INVX1_LOC_46/Y 0.07fF
C15042 INVX1_LOC_20/Y NAND2X1_LOC_686/A 0.02fF
C15043 INVX1_LOC_510/Y INVX1_LOC_119/Y 0.08fF
C15044 NAND2X1_LOC_703/a_36_24# INVX1_LOC_361/Y 0.01fF
C15045 INVX1_LOC_322/Y INVX1_LOC_100/Y 0.05fF
C15046 INVX1_LOC_99/Y INVX1_LOC_68/A 0.01fF
C15047 INVX1_LOC_686/A INVX1_LOC_501/A 0.07fF
C15048 INVX1_LOC_407/Y INVX1_LOC_117/Y 0.64fF
C15049 INVX1_LOC_166/A INVX1_LOC_252/A 0.02fF
C15050 INVX1_LOC_202/Y NAND2X1_LOC_333/B 0.19fF
C15051 INVX1_LOC_335/Y INVX1_LOC_69/Y 0.03fF
C15052 INVX1_LOC_87/A INVX1_LOC_178/A 0.05fF
C15053 INVX1_LOC_460/Y INVX1_LOC_513/A 0.01fF
C15054 INVX1_LOC_21/Y INVX1_LOC_69/Y 0.25fF
C15055 INVX1_LOC_117/Y INVX1_LOC_480/Y 0.01fF
C15056 INVX1_LOC_312/Y INVX1_LOC_301/Y 0.98fF
C15057 INVX1_LOC_20/Y INVX1_LOC_519/Y 0.01fF
C15058 INVX1_LOC_11/Y INVX1_LOC_32/Y 0.13fF
C15059 INVX1_LOC_84/A INVX1_LOC_117/A 0.01fF
C15060 INVX1_LOC_31/Y INVX1_LOC_352/Y 0.03fF
C15061 INVX1_LOC_276/A INVX1_LOC_102/Y 0.01fF
C15062 INVX1_LOC_586/A INVX1_LOC_41/Y 6.59fF
C15063 INVX1_LOC_76/Y INVX1_LOC_319/A 0.03fF
C15064 NAND2X1_LOC_192/A INVX1_LOC_633/Y 0.00fF
C15065 INVX1_LOC_362/Y NAND2X1_LOC_372/Y 0.23fF
C15066 INVX1_LOC_46/Y INVX1_LOC_83/Y 0.72fF
C15067 INVX1_LOC_686/Y INVX1_LOC_259/Y 0.01fF
C15068 INVX1_LOC_35/Y INVX1_LOC_633/A 0.00fF
C15069 INVX1_LOC_367/A INVX1_LOC_518/A 0.03fF
C15070 INVX1_LOC_186/A INVX1_LOC_139/Y 0.00fF
C15071 INVX1_LOC_93/Y INVX1_LOC_186/Y 0.10fF
C15072 INVX1_LOC_492/A INVX1_LOC_523/Y 0.01fF
C15073 INVX1_LOC_47/Y INVX1_LOC_509/A 0.02fF
C15074 INVX1_LOC_449/Y INVX1_LOC_6/Y 0.01fF
C15075 NAND2X1_LOC_822/Y INVX1_LOC_656/A 0.09fF
C15076 INVX1_LOC_31/Y INVX1_LOC_345/A 0.03fF
C15077 INVX1_LOC_117/Y INVX1_LOC_169/Y 0.19fF
C15078 INVX1_LOC_63/Y INVX1_LOC_145/Y 1.10fF
C15079 INVX1_LOC_562/A INVX1_LOC_636/A 0.08fF
C15080 INVX1_LOC_425/A INVX1_LOC_75/Y 0.04fF
C15081 INVX1_LOC_539/Y NAND2X1_LOC_689/B 0.00fF
C15082 INVX1_LOC_272/Y INVX1_LOC_531/Y 0.00fF
C15083 INVX1_LOC_287/A INVX1_LOC_242/Y 0.02fF
C15084 INVX1_LOC_69/Y NAND2X1_LOC_274/a_36_24# 0.01fF
C15085 INVX1_LOC_489/A NAND2X1_LOC_631/B 0.00fF
C15086 INVX1_LOC_103/Y INVX1_LOC_47/Y 0.03fF
C15087 INVX1_LOC_312/Y INVX1_LOC_41/Y 0.03fF
C15088 INVX1_LOC_137/Y INVX1_LOC_168/Y 0.08fF
C15089 NAND2X1_LOC_450/a_36_24# INVX1_LOC_74/Y 0.02fF
C15090 INVX1_LOC_355/A NAND2X1_LOC_449/a_36_24# 0.02fF
C15091 INVX1_LOC_166/A INVX1_LOC_6/Y 0.02fF
C15092 INVX1_LOC_211/Y INVX1_LOC_482/Y 0.05fF
C15093 INVX1_LOC_69/Y NAND2X1_LOC_267/A 0.19fF
C15094 INVX1_LOC_361/Y INVX1_LOC_49/Y 0.14fF
C15095 NAND2X1_LOC_602/A INVX1_LOC_376/Y 0.05fF
C15096 INVX1_LOC_298/A NAND2X1_LOC_836/B 0.00fF
C15097 INVX1_LOC_435/A INVX1_LOC_224/A 0.05fF
C15098 INVX1_LOC_507/Y INVX1_LOC_48/Y 0.08fF
C15099 INVX1_LOC_686/A NAND2X1_LOC_544/B 0.31fF
C15100 INVX1_LOC_602/A INVX1_LOC_74/A 0.02fF
C15101 INVX1_LOC_76/Y INVX1_LOC_91/Y 0.03fF
C15102 INVX1_LOC_49/Y NAND2X1_LOC_333/B 0.70fF
C15103 INVX1_LOC_116/Y INVX1_LOC_128/Y 0.01fF
C15104 INVX1_LOC_54/Y INVX1_LOC_376/Y 0.07fF
C15105 INVX1_LOC_58/Y INVX1_LOC_641/Y 0.03fF
C15106 INVX1_LOC_93/Y INVX1_LOC_347/Y 0.03fF
C15107 INVX1_LOC_476/A NAND2X1_LOC_277/a_36_24# 0.00fF
C15108 INVX1_LOC_119/Y INVX1_LOC_509/A 0.04fF
C15109 INVX1_LOC_607/Y INVX1_LOC_669/A 0.02fF
C15110 INVX1_LOC_26/Y NAND2X1_LOC_432/Y 0.15fF
C15111 INVX1_LOC_93/Y INVX1_LOC_328/Y 0.03fF
C15112 INVX1_LOC_261/Y INVX1_LOC_49/Y 0.03fF
C15113 NAND2X1_LOC_775/B INVX1_LOC_100/Y 0.47fF
C15114 INVX1_LOC_41/Y NAND2X1_LOC_378/Y 0.01fF
C15115 INVX1_LOC_411/A INVX1_LOC_79/A 0.01fF
C15116 INVX1_LOC_99/Y INVX1_LOC_635/Y 0.61fF
C15117 INPUT_1 INVX1_LOC_90/Y 0.07fF
C15118 INVX1_LOC_79/A INVX1_LOC_295/Y 0.01fF
C15119 NAND2X1_LOC_847/A NAND2X1_LOC_246/a_36_24# 0.01fF
C15120 NAND2X1_LOC_706/B INVX1_LOC_100/Y 0.17fF
C15121 INVX1_LOC_103/Y INVX1_LOC_119/Y 0.00fF
C15122 INVX1_LOC_155/A INVX1_LOC_245/A 0.01fF
C15123 INVX1_LOC_675/A INVX1_LOC_347/Y 0.07fF
C15124 INVX1_LOC_501/A NAND2X1_LOC_334/A 0.03fF
C15125 NAND2X1_LOC_775/B INVX1_LOC_74/Y 0.07fF
C15126 INVX1_LOC_662/A NAND2X1_LOC_846/A 0.03fF
C15127 NAND2X1_LOC_136/Y INVX1_LOC_6/Y 0.01fF
C15128 NAND2X1_LOC_545/B INVX1_LOC_92/A 0.03fF
C15129 INVX1_LOC_47/Y NAND2X1_LOC_786/B 0.01fF
C15130 INVX1_LOC_292/Y INVX1_LOC_90/Y 0.00fF
C15131 NAND2X1_LOC_333/B INVX1_LOC_92/Y 0.01fF
C15132 INVX1_LOC_346/A INVX1_LOC_119/Y 0.01fF
C15133 INVX1_LOC_31/Y INVX1_LOC_280/A 5.38fF
C15134 INVX1_LOC_245/A INVX1_LOC_9/Y 0.07fF
C15135 NAND2X1_LOC_123/B INVX1_LOC_338/Y 0.07fF
C15136 INVX1_LOC_92/A INVX1_LOC_98/Y 0.11fF
C15137 NAND2X1_LOC_695/a_36_24# INVX1_LOC_464/Y 0.00fF
C15138 INVX1_LOC_51/A NAND2X1_LOC_543/B 0.04fF
C15139 INVX1_LOC_446/A INVX1_LOC_446/Y 0.09fF
C15140 INVX1_LOC_44/Y INVX1_LOC_621/A 0.04fF
C15141 INVX1_LOC_224/Y NAND2X1_LOC_176/Y 0.03fF
C15142 VDD INVX1_LOC_265/Y 0.26fF
C15143 INVX1_LOC_62/Y INVX1_LOC_245/A 0.10fF
C15144 INVX1_LOC_682/Y NAND2X1_LOC_372/Y 0.25fF
C15145 INVX1_LOC_6/Y INVX1_LOC_613/A 0.04fF
C15146 NAND2X1_LOC_475/A INVX1_LOC_228/Y -0.03fF
C15147 NAND2X1_LOC_373/a_36_24# INVX1_LOC_442/A 0.00fF
C15148 INVX1_LOC_257/Y INVX1_LOC_374/A 0.00fF
C15149 VDD INVX1_LOC_502/Y 0.46fF
C15150 INVX1_LOC_111/A INVX1_LOC_638/A 0.05fF
C15151 INVX1_LOC_338/Y INVX1_LOC_92/A 0.07fF
C15152 INVX1_LOC_584/A INVX1_LOC_45/Y 0.00fF
C15153 INVX1_LOC_435/A INVX1_LOC_109/Y 0.00fF
C15154 INVX1_LOC_412/Y NAND2X1_LOC_180/B 0.02fF
C15155 INVX1_LOC_205/Y NAND2X1_LOC_86/Y 0.09fF
C15156 INVX1_LOC_274/A INVX1_LOC_615/Y 0.00fF
C15157 INVX1_LOC_402/Y INVX1_LOC_554/A 0.01fF
C15158 VDD INVX1_LOC_136/Y 0.43fF
C15159 INVX1_LOC_446/A INVX1_LOC_145/Y 0.08fF
C15160 INPUT_0 INVX1_LOC_84/A 0.17fF
C15161 INVX1_LOC_224/Y INVX1_LOC_312/A 0.02fF
C15162 INVX1_LOC_224/Y NAND2X1_LOC_391/A 0.04fF
C15163 INVX1_LOC_315/Y INVX1_LOC_586/A 0.01fF
C15164 INVX1_LOC_560/Y NAND2X1_LOC_123/A 0.07fF
C15165 INVX1_LOC_573/A NAND2X1_LOC_728/A 0.10fF
C15166 INVX1_LOC_412/Y INVX1_LOC_188/Y 0.03fF
C15167 INVX1_LOC_424/A INVX1_LOC_442/Y 0.03fF
C15168 INVX1_LOC_629/Y INVX1_LOC_579/A 0.01fF
C15169 INVX1_LOC_566/A INVX1_LOC_259/A 0.03fF
C15170 VDD INVX1_LOC_25/Y 0.86fF
C15171 INVX1_LOC_20/Y INVX1_LOC_65/Y 0.10fF
C15172 INVX1_LOC_625/A NAND2X1_LOC_310/a_36_24# 0.00fF
C15173 VDD NAND2X1_LOC_43/Y 0.03fF
C15174 NAND2X1_LOC_669/Y INVX1_LOC_395/A 0.03fF
C15175 NAND2X1_LOC_790/B NAND2X1_LOC_615/B 0.18fF
C15176 INVX1_LOC_117/Y INVX1_LOC_638/A 0.07fF
C15177 NAND2X1_LOC_373/a_36_24# INVX1_LOC_116/Y 0.00fF
C15178 NAND2X1_LOC_164/Y INVX1_LOC_197/Y 0.03fF
C15179 INVX1_LOC_274/A INVX1_LOC_395/A 0.52fF
C15180 INVX1_LOC_552/Y INVX1_LOC_145/Y 0.03fF
C15181 NAND2X1_LOC_97/B INVX1_LOC_269/A 0.01fF
C15182 INVX1_LOC_206/Y INVX1_LOC_194/Y 0.03fF
C15183 INVX1_LOC_273/A INVX1_LOC_97/Y 0.01fF
C15184 INVX1_LOC_335/Y INVX1_LOC_586/A 0.03fF
C15185 INVX1_LOC_395/A INVX1_LOC_209/A 0.02fF
C15186 NAND2X1_LOC_332/B INVX1_LOC_670/Y 0.19fF
C15187 INVX1_LOC_511/A INVX1_LOC_522/Y 0.19fF
C15188 INVX1_LOC_21/Y INVX1_LOC_586/A 0.74fF
C15189 NAND2X1_LOC_336/B INVX1_LOC_270/A 0.04fF
C15190 INVX1_LOC_439/Y INVX1_LOC_445/A 0.05fF
C15191 INVX1_LOC_45/Y INVX1_LOC_537/A 0.39fF
C15192 INVX1_LOC_65/Y INVX1_LOC_300/A 0.08fF
C15193 INVX1_LOC_20/Y INVX1_LOC_287/A 0.12fF
C15194 INVX1_LOC_395/A INVX1_LOC_186/Y 0.41fF
C15195 NAND2X1_LOC_498/Y INVX1_LOC_105/A 0.07fF
C15196 INVX1_LOC_400/A INVX1_LOC_266/Y 0.07fF
C15197 NAND2X1_LOC_547/a_36_24# NAND2X1_LOC_457/A 0.00fF
C15198 INVX1_LOC_51/Y INVX1_LOC_352/Y 0.03fF
C15199 NAND2X1_LOC_324/B INVX1_LOC_80/A 0.03fF
C15200 INVX1_LOC_248/Y INVX1_LOC_353/Y 0.92fF
C15201 INVX1_LOC_614/A INVX1_LOC_136/Y 0.01fF
C15202 INVX1_LOC_291/A NAND2X1_LOC_93/a_36_24# -0.01fF
C15203 INVX1_LOC_412/A INVX1_LOC_46/Y 0.01fF
C15204 INVX1_LOC_53/Y NAND2X1_LOC_145/a_36_24# 0.00fF
C15205 NAND2X1_LOC_507/A INVX1_LOC_397/A 0.09fF
C15206 INVX1_LOC_133/Y INVX1_LOC_100/Y 0.00fF
C15207 NAND2X1_LOC_185/a_36_24# INVX1_LOC_117/Y 0.00fF
C15208 INVX1_LOC_93/Y INVX1_LOC_165/Y 0.07fF
C15209 VDD INVX1_LOC_15/Y 0.21fF
C15210 INVX1_LOC_210/Y NAND2X1_LOC_79/B 0.11fF
C15211 INVX1_LOC_435/Y NAND2X1_LOC_106/Y 0.05fF
C15212 INVX1_LOC_98/A NAND2X1_LOC_333/B 0.83fF
C15213 INVX1_LOC_586/A NAND2X1_LOC_267/A 0.07fF
C15214 INVX1_LOC_167/Y INVX1_LOC_137/Y 0.13fF
C15215 INVX1_LOC_526/A INVX1_LOC_259/Y 0.28fF
C15216 INPUT_0 INVX1_LOC_496/A 0.05fF
C15217 NAND2X1_LOC_534/Y INVX1_LOC_376/Y 0.02fF
C15218 INVX1_LOC_206/Y INVX1_LOC_44/Y 0.16fF
C15219 INVX1_LOC_421/A INVX1_LOC_45/Y 0.21fF
C15220 INVX1_LOC_45/Y INVX1_LOC_496/Y 0.03fF
C15221 NAND2X1_LOC_331/A INVX1_LOC_58/Y 0.06fF
C15222 INVX1_LOC_164/Y INVX1_LOC_76/Y 0.17fF
C15223 INPUT_3 NAND2X1_LOC_37/a_36_24# 0.01fF
C15224 VDD INVX1_LOC_663/A 0.00fF
C15225 INVX1_LOC_103/Y INVX1_LOC_502/Y 0.01fF
C15226 INVX1_LOC_76/Y NAND2X1_LOC_333/B 0.05fF
C15227 INVX1_LOC_255/Y INVX1_LOC_69/Y 0.05fF
C15228 INVX1_LOC_145/Y INVX1_LOC_387/A 0.09fF
C15229 INVX1_LOC_522/Y INVX1_LOC_48/Y 0.08fF
C15230 INVX1_LOC_413/A INVX1_LOC_293/Y 0.08fF
C15231 INVX1_LOC_287/A INVX1_LOC_300/A 0.01fF
C15232 INVX1_LOC_224/Y INVX1_LOC_226/Y 0.01fF
C15233 INVX1_LOC_37/Y INVX1_LOC_328/Y 0.01fF
C15234 INVX1_LOC_287/A INVX1_LOC_197/Y 1.46fF
C15235 NAND2X1_LOC_526/Y INVX1_LOC_420/A 0.17fF
C15236 VDD NAND2X1_LOC_627/Y 0.01fF
C15237 INVX1_LOC_395/A INVX1_LOC_328/Y 0.03fF
C15238 INVX1_LOC_21/Y NAND2X1_LOC_378/Y 0.82fF
C15239 VDD INVX1_LOC_475/Y 0.26fF
C15240 INVX1_LOC_442/Y INVX1_LOC_363/Y 0.03fF
C15241 INVX1_LOC_577/Y INVX1_LOC_69/Y 0.03fF
C15242 INVX1_LOC_206/Y INVX1_LOC_461/Y 0.26fF
C15243 INVX1_LOC_105/Y INVX1_LOC_367/A 0.01fF
C15244 NAND2X1_LOC_545/B INPUT_1 0.59fF
C15245 NAND2X1_LOC_821/a_36_24# INVX1_LOC_59/A 0.00fF
C15246 NAND2X1_LOC_317/B INVX1_LOC_100/Y 0.03fF
C15247 INPUT_3 INVX1_LOC_84/Y 0.03fF
C15248 INVX1_LOC_517/A INVX1_LOC_46/Y 0.01fF
C15249 NAND2X1_LOC_332/B INVX1_LOC_63/Y 0.01fF
C15250 NAND2X1_LOC_516/B INVX1_LOC_199/Y 0.18fF
C15251 NAND2X1_LOC_336/B INVX1_LOC_46/Y 0.04fF
C15252 INVX1_LOC_445/Y INVX1_LOC_430/Y 0.18fF
C15253 INVX1_LOC_370/Y INVX1_LOC_50/Y 0.02fF
C15254 INVX1_LOC_449/A INVX1_LOC_31/Y 0.02fF
C15255 INVX1_LOC_171/A INVX1_LOC_99/Y 0.01fF
C15256 INVX1_LOC_300/A NAND2X1_LOC_807/a_36_24# 0.00fF
C15257 INVX1_LOC_20/Y INVX1_LOC_95/A 0.03fF
C15258 INVX1_LOC_562/A INVX1_LOC_74/Y 0.16fF
C15259 INVX1_LOC_455/A INVX1_LOC_40/Y 0.01fF
C15260 INVX1_LOC_335/Y NAND2X1_LOC_835/A 0.08fF
C15261 INPUT_1 INVX1_LOC_98/Y 0.03fF
C15262 INVX1_LOC_189/Y INVX1_LOC_186/Y 0.12fF
C15263 INVX1_LOC_140/Y INVX1_LOC_41/Y 0.04fF
C15264 INVX1_LOC_105/Y INVX1_LOC_669/Y 0.00fF
C15265 INVX1_LOC_449/Y INVX1_LOC_415/Y 0.92fF
C15266 INVX1_LOC_659/Y INVX1_LOC_659/A 0.10fF
C15267 NAND2X1_LOC_174/B INVX1_LOC_259/Y 0.03fF
C15268 INVX1_LOC_11/Y INVX1_LOC_110/A 0.03fF
C15269 INVX1_LOC_402/Y INVX1_LOC_199/Y 0.06fF
C15270 INVX1_LOC_48/Y INVX1_LOC_295/Y 0.03fF
C15271 INVX1_LOC_117/Y INVX1_LOC_665/Y 0.03fF
C15272 NAND2X1_LOC_591/Y INVX1_LOC_259/Y 0.01fF
C15273 INVX1_LOC_51/Y INVX1_LOC_280/A 0.12fF
C15274 NAND2X1_LOC_48/a_36_24# INVX1_LOC_63/Y 0.00fF
C15275 INVX1_LOC_600/A NAND2X1_LOC_52/a_36_24# 0.01fF
C15276 INVX1_LOC_51/Y NAND2X1_LOC_372/Y 0.07fF
C15277 NAND2X1_LOC_426/Y INVX1_LOC_41/Y 0.02fF
C15278 INVX1_LOC_449/Y NAND2X1_LOC_294/Y 0.06fF
C15279 NAND2X1_LOC_836/B INVX1_LOC_145/Y 0.06fF
C15280 INVX1_LOC_442/Y INVX1_LOC_49/Y 0.07fF
C15281 INVX1_LOC_556/Y INVX1_LOC_66/A 0.03fF
C15282 INVX1_LOC_197/A INVX1_LOC_114/A 0.03fF
C15283 INVX1_LOC_344/A INVX1_LOC_245/A 0.03fF
C15284 INVX1_LOC_543/Y INVX1_LOC_87/Y 0.15fF
C15285 NAND2X1_LOC_147/B INVX1_LOC_662/A 0.35fF
C15286 INVX1_LOC_407/Y INVX1_LOC_58/Y 0.21fF
C15287 INVX1_LOC_105/A INVX1_LOC_47/Y 0.09fF
C15288 INVX1_LOC_20/Y INVX1_LOC_588/A 0.03fF
C15289 INVX1_LOC_359/A INVX1_LOC_372/A 0.17fF
C15290 NAND2X1_LOC_140/B INVX1_LOC_519/Y 0.08fF
C15291 INVX1_LOC_495/A INVX1_LOC_74/Y 0.02fF
C15292 INVX1_LOC_686/A INVX1_LOC_347/A 0.04fF
C15293 INVX1_LOC_266/A NAND2X1_LOC_438/a_36_24# 0.00fF
C15294 INVX1_LOC_116/Y NAND2X1_LOC_605/B 0.00fF
C15295 INVX1_LOC_598/A INVX1_LOC_63/Y 0.01fF
C15296 INVX1_LOC_6/Y NAND2X1_LOC_627/a_36_24# 0.00fF
C15297 INPUT_1 INVX1_LOC_338/Y 0.53fF
C15298 INVX1_LOC_84/A INVX1_LOC_211/A 0.03fF
C15299 NAND2X1_LOC_27/Y INVX1_LOC_9/Y 0.05fF
C15300 INVX1_LOC_578/Y INVX1_LOC_533/A 0.01fF
C15301 INVX1_LOC_89/Y NAND2X1_LOC_542/A 0.04fF
C15302 NAND2X1_LOC_336/B INVX1_LOC_75/A 0.26fF
C15303 NAND2X1_LOC_847/A INVX1_LOC_46/Y 0.00fF
C15304 INVX1_LOC_519/A INVX1_LOC_666/Y 0.02fF
C15305 INVX1_LOC_504/A NAND2X1_LOC_123/B 0.17fF
C15306 NAND2X1_LOC_775/B INVX1_LOC_79/A 0.11fF
C15307 NAND2X1_LOC_128/B INVX1_LOC_63/Y 0.05fF
C15308 INVX1_LOC_31/Y INVX1_LOC_328/Y 0.07fF
C15309 INVX1_LOC_166/A INVX1_LOC_557/Y 0.00fF
C15310 INVX1_LOC_105/A INVX1_LOC_119/Y 1.67fF
C15311 NAND2X1_LOC_503/B INVX1_LOC_615/A 0.08fF
C15312 INVX1_LOC_171/A NAND2X1_LOC_66/Y 0.01fF
C15313 INVX1_LOC_50/Y INVX1_LOC_90/Y 0.03fF
C15314 INVX1_LOC_89/Y INVX1_LOC_376/Y 0.07fF
C15315 INVX1_LOC_532/Y INVX1_LOC_533/A 0.19fF
C15316 NAND2X1_LOC_675/B INVX1_LOC_347/Y 0.17fF
C15317 NAND2X1_LOC_308/a_36_24# INVX1_LOC_74/Y 0.00fF
C15318 NAND2X1_LOC_184/Y INVX1_LOC_665/A 0.06fF
C15319 INVX1_LOC_431/Y INVX1_LOC_90/Y 0.02fF
C15320 INVX1_LOC_69/Y INVX1_LOC_128/Y 0.00fF
C15321 INVX1_LOC_69/Y INVX1_LOC_26/Y 0.33fF
C15322 INVX1_LOC_63/Y INVX1_LOC_242/Y 0.07fF
C15323 INVX1_LOC_643/Y NAND2X1_LOC_846/B 0.05fF
C15324 VDD INVX1_LOC_279/Y 0.18fF
C15325 NAND2X1_LOC_119/a_36_24# INVX1_LOC_74/Y 0.00fF
C15326 INVX1_LOC_6/Y INVX1_LOC_41/Y 1.39fF
C15327 VDD NAND2X1_LOC_543/B 0.37fF
C15328 INVX1_LOC_75/Y INVX1_LOC_234/Y 0.02fF
C15329 INVX1_LOC_459/A NAND2X1_LOC_592/B 0.12fF
C15330 INVX1_LOC_405/A INVX1_LOC_446/Y 0.04fF
C15331 INVX1_LOC_199/Y INVX1_LOC_241/A 0.00fF
C15332 NAND2X1_LOC_286/A NAND2X1_LOC_843/B 0.03fF
C15333 INVX1_LOC_588/Y INVX1_LOC_636/A 0.02fF
C15334 INVX1_LOC_206/Y NAND2X1_LOC_176/Y 0.01fF
C15335 INVX1_LOC_386/A INVX1_LOC_62/Y 0.01fF
C15336 INVX1_LOC_273/A INVX1_LOC_615/A 0.33fF
C15337 INVX1_LOC_367/A INVX1_LOC_109/Y 0.02fF
C15338 INVX1_LOC_450/A INVX1_LOC_453/A 0.27fF
C15339 VDD NAND2X1_LOC_520/B 0.01fF
C15340 NAND2X1_LOC_317/A INVX1_LOC_395/A 0.02fF
C15341 VDD INVX1_LOC_131/Y 0.21fF
C15342 NAND2X1_LOC_45/Y INVX1_LOC_45/Y 0.18fF
C15343 NAND2X1_LOC_798/a_36_24# INVX1_LOC_638/A 0.00fF
C15344 INVX1_LOC_206/Y INVX1_LOC_96/Y 0.03fF
C15345 INVX1_LOC_203/Y INVX1_LOC_94/A 0.03fF
C15346 INVX1_LOC_665/A INVX1_LOC_75/Y 0.04fF
C15347 INVX1_LOC_395/A INVX1_LOC_521/Y 0.01fF
C15348 GATE_579 INVX1_LOC_438/Y 0.35fF
C15349 INVX1_LOC_554/A INVX1_LOC_367/A 0.06fF
C15350 INVX1_LOC_233/Y INVX1_LOC_420/Y 0.01fF
C15351 VDD INVX1_LOC_23/Y 0.24fF
C15352 NAND2X1_LOC_45/Y INPUT_3 0.12fF
C15353 NAND2X1_LOC_498/Y INVX1_LOC_45/Y 0.01fF
C15354 INPUT_0 NAND2X1_LOC_79/B 0.01fF
C15355 INVX1_LOC_405/A INVX1_LOC_145/Y 0.01fF
C15356 INVX1_LOC_425/A INVX1_LOC_578/A 0.79fF
C15357 INVX1_LOC_479/A INVX1_LOC_109/A 0.00fF
C15358 VDD NAND2X1_LOC_638/A 0.20fF
C15359 INVX1_LOC_96/Y INVX1_LOC_396/Y 0.06fF
C15360 INVX1_LOC_224/Y INVX1_LOC_297/A 0.09fF
C15361 VDD INVX1_LOC_469/A -0.00fF
C15362 NAND2X1_LOC_554/a_36_24# INVX1_LOC_99/Y 0.01fF
C15363 INVX1_LOC_321/Y INVX1_LOC_596/Y 0.92fF
C15364 NAND2X1_LOC_383/Y NAND2X1_LOC_391/B 0.27fF
C15365 INVX1_LOC_20/Y NAND2X1_LOC_335/a_36_24# 0.00fF
C15366 INVX1_LOC_95/Y INVX1_LOC_93/Y 0.06fF
C15367 NAND2X1_LOC_750/Y INVX1_LOC_64/A -0.00fF
C15368 NAND2X1_LOC_231/A INVX1_LOC_287/Y 0.00fF
C15369 INVX1_LOC_490/Y INVX1_LOC_519/A 0.03fF
C15370 INVX1_LOC_185/A INVX1_LOC_575/Y 0.02fF
C15371 VDD INVX1_LOC_505/A 0.38fF
C15372 INVX1_LOC_448/Y INVX1_LOC_665/Y 0.01fF
C15373 INVX1_LOC_435/Y INVX1_LOC_679/Y 0.44fF
C15374 INVX1_LOC_272/Y INVX1_LOC_315/Y 0.01fF
C15375 INVX1_LOC_224/Y INVX1_LOC_252/Y 0.61fF
C15376 INVX1_LOC_390/A INVX1_LOC_109/Y 0.00fF
C15377 INVX1_LOC_395/A INVX1_LOC_352/A 0.01fF
C15378 INVX1_LOC_45/Y INVX1_LOC_676/Y 0.02fF
C15379 INVX1_LOC_449/A INVX1_LOC_51/Y 0.46fF
C15380 INVX1_LOC_560/Y INVX1_LOC_248/A 0.01fF
C15381 NAND2X1_LOC_703/a_36_24# INVX1_LOC_412/A 0.00fF
C15382 INVX1_LOC_395/A NAND2X1_LOC_459/a_36_24# 0.00fF
C15383 INVX1_LOC_578/A INVX1_LOC_252/Y 0.07fF
C15384 INVX1_LOC_238/Y INVX1_LOC_117/Y 0.03fF
C15385 INVX1_LOC_99/Y NAND2X1_LOC_506/B 0.40fF
C15386 INVX1_LOC_482/Y INVX1_LOC_297/Y 0.38fF
C15387 INVX1_LOC_193/A INPUT_0 0.06fF
C15388 INVX1_LOC_53/Y NAND2X1_LOC_516/B 0.01fF
C15389 INVX1_LOC_301/A INVX1_LOC_253/Y 0.08fF
C15390 INVX1_LOC_335/Y INVX1_LOC_587/A 0.03fF
C15391 INVX1_LOC_367/A INVX1_LOC_126/Y 0.02fF
C15392 VDD INVX1_LOC_326/Y 0.36fF
C15393 INVX1_LOC_21/Y INVX1_LOC_366/A 0.01fF
C15394 INVX1_LOC_45/Y INVX1_LOC_99/Y 6.68fF
C15395 NAND2X1_LOC_249/Y INVX1_LOC_69/Y 0.14fF
C15396 INVX1_LOC_547/Y NAND2X1_LOC_106/B 0.00fF
C15397 INVX1_LOC_20/Y INVX1_LOC_670/Y 0.16fF
C15398 INVX1_LOC_54/Y NAND2X1_LOC_750/a_36_24# 0.00fF
C15399 INVX1_LOC_266/A INVX1_LOC_67/Y 0.00fF
C15400 INVX1_LOC_17/Y INVX1_LOC_666/A 0.03fF
C15401 INVX1_LOC_271/A INVX1_LOC_48/Y 0.01fF
C15402 INVX1_LOC_378/A NAND2X1_LOC_416/Y 0.00fF
C15403 INVX1_LOC_393/Y INVX1_LOC_32/Y 0.02fF
C15404 INVX1_LOC_596/A INVX1_LOC_679/Y 0.48fF
C15405 INPUT_0 NAND2X1_LOC_532/Y 0.03fF
C15406 INVX1_LOC_134/Y INVX1_LOC_104/Y 0.04fF
C15407 NAND2X1_LOC_148/A NAND2X1_LOC_145/a_36_24# 0.02fF
C15408 INPUT_3 INVX1_LOC_99/Y 0.05fF
C15409 INVX1_LOC_21/Y INVX1_LOC_294/Y 0.10fF
C15410 INVX1_LOC_90/Y INVX1_LOC_275/A 0.04fF
C15411 INVX1_LOC_395/A GATE_662 0.05fF
C15412 INVX1_LOC_648/Y INVX1_LOC_523/Y 0.03fF
C15413 INVX1_LOC_165/Y INVX1_LOC_31/Y 0.03fF
C15414 INVX1_LOC_218/Y INVX1_LOC_218/A 0.15fF
C15415 INVX1_LOC_84/A INVX1_LOC_145/Y 0.13fF
C15416 INVX1_LOC_602/A INVX1_LOC_316/Y 0.03fF
C15417 INVX1_LOC_402/Y INVX1_LOC_53/Y 0.01fF
C15418 INVX1_LOC_89/Y INVX1_LOC_253/A 0.00fF
C15419 INVX1_LOC_342/Y INVX1_LOC_59/A 0.01fF
C15420 NAND2X1_LOC_303/a_36_24# INVX1_LOC_559/Y 0.00fF
C15421 INVX1_LOC_560/A INVX1_LOC_69/Y 0.08fF
C15422 INVX1_LOC_428/Y NAND2X1_LOC_523/B 0.06fF
C15423 VDD INVX1_LOC_353/A 0.09fF
C15424 NAND2X1_LOC_759/B INVX1_LOC_79/A 0.01fF
C15425 INVX1_LOC_589/Y INVX1_LOC_45/Y 0.01fF
C15426 INVX1_LOC_564/Y INVX1_LOC_69/Y 0.01fF
C15427 INVX1_LOC_451/A INVX1_LOC_46/A 0.37fF
C15428 INVX1_LOC_671/A NAND2X1_LOC_842/a_36_24# 0.01fF
C15429 NAND2X1_LOC_106/B INVX1_LOC_651/A 0.00fF
C15430 INVX1_LOC_168/A INVX1_LOC_54/Y 0.07fF
C15431 NAND2X1_LOC_93/Y INVX1_LOC_90/Y 0.01fF
C15432 NAND2X1_LOC_181/a_36_24# INVX1_LOC_519/A 0.01fF
C15433 INVX1_LOC_315/Y INVX1_LOC_6/Y 0.03fF
C15434 INVX1_LOC_395/A NAND2X1_LOC_846/B 0.03fF
C15435 INVX1_LOC_206/Y NAND2X1_LOC_616/a_36_24# 0.00fF
C15436 INVX1_LOC_47/Y INVX1_LOC_45/Y 0.25fF
C15437 INVX1_LOC_45/Y NAND2X1_LOC_557/B 0.00fF
C15438 INVX1_LOC_49/Y INVX1_LOC_618/Y 0.03fF
C15439 INVX1_LOC_386/Y INVX1_LOC_442/Y 0.07fF
C15440 INVX1_LOC_596/A INPUT_1 0.03fF
C15441 INVX1_LOC_523/Y INVX1_LOC_242/A 0.65fF
C15442 INVX1_LOC_105/Y INVX1_LOC_683/Y 0.01fF
C15443 INVX1_LOC_366/A INVX1_LOC_181/Y 0.03fF
C15444 INVX1_LOC_12/Y INVX1_LOC_304/Y 0.04fF
C15445 INVX1_LOC_93/Y INVX1_LOC_126/Y 0.08fF
C15446 INVX1_LOC_293/Y INVX1_LOC_421/A 0.65fF
C15447 NAND2X1_LOC_317/B INVX1_LOC_79/A 0.02fF
C15448 INVX1_LOC_409/Y INVX1_LOC_441/A 0.01fF
C15449 INVX1_LOC_145/Y NAND2X1_LOC_67/Y 0.18fF
C15450 INVX1_LOC_45/A INVX1_LOC_18/Y 0.00fF
C15451 INVX1_LOC_117/Y INVX1_LOC_134/Y 3.44fF
C15452 INVX1_LOC_468/Y INVX1_LOC_252/Y 0.83fF
C15453 INVX1_LOC_419/Y INVX1_LOC_99/A 0.01fF
C15454 INVX1_LOC_211/Y INVX1_LOC_321/Y 0.05fF
C15455 INVX1_LOC_425/A INVX1_LOC_120/Y 0.01fF
C15456 NAND2X1_LOC_184/Y INVX1_LOC_80/A 0.19fF
C15457 INVX1_LOC_469/Y INVX1_LOC_633/Y 0.02fF
C15458 INVX1_LOC_176/A INVX1_LOC_35/Y 0.01fF
C15459 INVX1_LOC_17/Y NAND2X1_LOC_673/A 0.02fF
C15460 INPUT_3 INVX1_LOC_47/Y 0.07fF
C15461 INVX1_LOC_583/A INVX1_LOC_93/Y 0.00fF
C15462 INVX1_LOC_51/Y INVX1_LOC_328/Y 0.09fF
C15463 INVX1_LOC_271/Y INVX1_LOC_245/A 0.01fF
C15464 INVX1_LOC_53/Y NAND2X1_LOC_718/a_36_24# 0.01fF
C15465 INVX1_LOC_20/Y INVX1_LOC_63/Y 0.81fF
C15466 INVX1_LOC_76/Y INVX1_LOC_482/Y 0.02fF
C15467 INVX1_LOC_51/Y INVX1_LOC_518/A 0.16fF
C15468 INVX1_LOC_175/Y INVX1_LOC_63/Y 0.01fF
C15469 INVX1_LOC_586/A NAND2X1_LOC_420/a_36_24# 0.00fF
C15470 NAND2X1_LOC_863/a_36_24# INVX1_LOC_58/Y 0.01fF
C15471 INVX1_LOC_367/A INVX1_LOC_199/Y 0.02fF
C15472 INVX1_LOC_586/A INVX1_LOC_26/Y 0.13fF
C15473 INVX1_LOC_45/Y INVX1_LOC_119/Y 0.53fF
C15474 NAND2X1_LOC_43/Y INVX1_LOC_171/A 0.02fF
C15475 INVX1_LOC_317/Y INVX1_LOC_100/Y 0.11fF
C15476 INVX1_LOC_50/Y INVX1_LOC_98/Y 0.07fF
C15477 NAND2X1_LOC_320/Y INVX1_LOC_93/Y 0.01fF
C15478 INVX1_LOC_76/Y INVX1_LOC_471/Y 0.00fF
C15479 INVX1_LOC_45/Y NAND2X1_LOC_66/Y 0.08fF
C15480 INVX1_LOC_335/Y INVX1_LOC_6/Y 0.05fF
C15481 INVX1_LOC_31/Y INVX1_LOC_352/A 0.01fF
C15482 INVX1_LOC_21/Y INVX1_LOC_6/Y 3.11fF
C15483 NAND2X1_LOC_775/B INVX1_LOC_48/Y 0.07fF
C15484 INVX1_LOC_270/Y NAND2X1_LOC_76/B 0.04fF
C15485 INVX1_LOC_674/A INVX1_LOC_637/A 0.07fF
C15486 NAND2X1_LOC_747/a_36_24# INVX1_LOC_137/Y 0.00fF
C15487 NAND2X1_LOC_613/Y INVX1_LOC_79/A 0.01fF
C15488 INVX1_LOC_551/Y NAND2X1_LOC_274/B 0.03fF
C15489 INVX1_LOC_11/Y NAND2X1_LOC_184/Y 0.07fF
C15490 INVX1_LOC_99/Y NAND2X1_LOC_276/A 0.09fF
C15491 INVX1_LOC_183/A INVX1_LOC_12/Y 0.72fF
C15492 INVX1_LOC_25/Y INVX1_LOC_145/A 0.21fF
C15493 INVX1_LOC_47/Y NAND2X1_LOC_69/Y 0.03fF
C15494 INVX1_LOC_92/A NAND2X1_LOC_76/B 0.00fF
C15495 INVX1_LOC_69/Y NAND2X1_LOC_275/Y 0.01fF
C15496 NAND2X1_LOC_662/a_36_24# INVX1_LOC_655/A 0.00fF
C15497 INPUT_3 NAND2X1_LOC_66/Y 1.22fF
C15498 INVX1_LOC_32/Y NAND2X1_LOC_333/B 0.07fF
C15499 NAND2X1_LOC_442/a_36_24# INPUT_1 0.00fF
C15500 INVX1_LOC_6/Y NAND2X1_LOC_274/a_36_24# 0.00fF
C15501 INVX1_LOC_410/A INVX1_LOC_35/Y 0.01fF
C15502 INVX1_LOC_400/A INVX1_LOC_199/Y 0.82fF
C15503 INVX1_LOC_300/A INVX1_LOC_63/Y 0.29fF
C15504 INVX1_LOC_63/Y INVX1_LOC_197/Y 0.03fF
C15505 INVX1_LOC_170/Y INVX1_LOC_35/Y 0.01fF
C15506 INVX1_LOC_79/A INVX1_LOC_633/Y 0.03fF
C15507 INVX1_LOC_587/Y NAND2X1_LOC_753/Y 0.05fF
C15508 INVX1_LOC_261/Y INVX1_LOC_32/Y 0.03fF
C15509 INVX1_LOC_504/A NAND2X1_LOC_683/a_36_24# 0.00fF
C15510 INVX1_LOC_497/A INVX1_LOC_50/Y 0.03fF
C15511 INVX1_LOC_399/Y INVX1_LOC_35/Y 0.00fF
C15512 INVX1_LOC_50/Y INVX1_LOC_338/Y 0.03fF
C15513 INVX1_LOC_93/Y INVX1_LOC_199/Y 1.49fF
C15514 INVX1_LOC_26/Y NAND2X1_LOC_378/Y 0.03fF
C15515 NAND2X1_LOC_126/a_36_24# INVX1_LOC_42/Y 0.00fF
C15516 INVX1_LOC_80/A INVX1_LOC_75/Y 0.07fF
C15517 INVX1_LOC_249/A INVX1_LOC_74/Y 0.15fF
C15518 INVX1_LOC_161/A INVX1_LOC_41/Y 0.00fF
C15519 INVX1_LOC_6/Y INVX1_LOC_181/Y 0.01fF
C15520 NAND2X1_LOC_488/Y INVX1_LOC_600/A 0.01fF
C15521 INVX1_LOC_580/A INVX1_LOC_636/A 0.05fF
C15522 NAND2X1_LOC_638/A INVX1_LOC_635/Y 0.03fF
C15523 INVX1_LOC_376/A INVX1_LOC_355/Y 0.02fF
C15524 INVX1_LOC_507/Y INVX1_LOC_633/A 0.01fF
C15525 INVX1_LOC_292/Y INVX1_LOC_622/A 0.01fF
C15526 INPUT_5 NAND2X1_LOC_425/a_36_24# 0.00fF
C15527 INVX1_LOC_288/Y INVX1_LOC_479/A 0.03fF
C15528 INVX1_LOC_54/Y INVX1_LOC_652/A 0.12fF
C15529 INVX1_LOC_93/Y INVX1_LOC_272/A 0.00fF
C15530 INVX1_LOC_166/A INVX1_LOC_100/Y 0.06fF
C15531 NAND2X1_LOC_32/Y INVX1_LOC_41/Y 0.00fF
C15532 INVX1_LOC_11/Y INVX1_LOC_75/Y 0.81fF
C15533 INVX1_LOC_644/Y NAND2X1_LOC_814/Y 0.23fF
C15534 INVX1_LOC_69/Y NAND2X1_LOC_605/B 0.01fF
C15535 INVX1_LOC_317/A INVX1_LOC_79/A 0.01fF
C15536 INVX1_LOC_588/Y INVX1_LOC_74/Y 0.03fF
C15537 INVX1_LOC_395/A INVX1_LOC_109/Y 0.20fF
C15538 INVX1_LOC_625/A INVX1_LOC_270/Y 0.02fF
C15539 NAND2X1_LOC_111/Y INVX1_LOC_100/Y 0.06fF
C15540 INVX1_LOC_166/A INVX1_LOC_74/Y 0.15fF
C15541 VDD NAND2X1_LOC_781/B 0.01fF
C15542 VDD INVX1_LOC_409/Y 0.44fF
C15543 INVX1_LOC_662/A NAND2X1_LOC_841/a_36_24# 0.02fF
C15544 INVX1_LOC_362/Y INVX1_LOC_109/Y 0.05fF
C15545 INVX1_LOC_625/A INVX1_LOC_92/A 0.38fF
C15546 INVX1_LOC_35/Y INVX1_LOC_611/A 0.01fF
C15547 NAND2X1_LOC_709/a_36_24# INVX1_LOC_100/Y 0.00fF
C15548 INVX1_LOC_95/Y INVX1_LOC_395/A 0.01fF
C15549 INVX1_LOC_26/Y INVX1_LOC_225/Y 0.09fF
C15550 VDD NAND2X1_LOC_335/B 0.03fF
C15551 INVX1_LOC_11/Y NAND2X1_LOC_271/A 0.17fF
C15552 NAND2X1_LOC_192/A INVX1_LOC_41/Y 0.01fF
C15553 INVX1_LOC_683/Y INVX1_LOC_109/Y 0.13fF
C15554 INVX1_LOC_463/A INVX1_LOC_584/Y 0.00fF
C15555 INVX1_LOC_366/A NAND2X1_LOC_86/a_36_24# 0.01fF
C15556 INVX1_LOC_531/Y INVX1_LOC_100/Y 0.05fF
C15557 INVX1_LOC_426/Y INVX1_LOC_586/A 0.01fF
C15558 INVX1_LOC_68/Y VDD 0.67fF
C15559 VDD INVX1_LOC_233/Y 0.30fF
C15560 NAND2X1_LOC_475/A INVX1_LOC_45/Y 0.03fF
C15561 VDD INVX1_LOC_88/Y 0.26fF
C15562 VDD INVX1_LOC_147/Y 0.21fF
C15563 NAND2X1_LOC_219/a_36_24# INVX1_LOC_85/Y 0.00fF
C15564 INVX1_LOC_425/A INVX1_LOC_206/Y 0.08fF
C15565 INVX1_LOC_100/Y INVX1_LOC_363/A 0.01fF
C15566 INVX1_LOC_426/Y INVX1_LOC_312/Y 0.01fF
C15567 INVX1_LOC_560/A INVX1_LOC_586/A 0.07fF
C15568 NAND2X1_LOC_249/Y INVX1_LOC_312/Y 0.13fF
C15569 INVX1_LOC_34/Y INVX1_LOC_33/A 0.02fF
C15570 INVX1_LOC_206/Y INVX1_LOC_126/A 0.00fF
C15571 VDD INVX1_LOC_250/Y 0.22fF
C15572 INVX1_LOC_96/Y INVX1_LOC_94/A 0.05fF
C15573 VDD INVX1_LOC_675/Y 0.21fF
C15574 VDD NAND2X1_LOC_130/Y 0.06fF
C15575 VDD INVX1_LOC_600/A 0.12fF
C15576 INVX1_LOC_206/Y INVX1_LOC_297/A 0.12fF
C15577 INVX1_LOC_182/A INVX1_LOC_191/A 0.04fF
C15578 INVX1_LOC_502/Y INVX1_LOC_45/Y 0.01fF
C15579 INVX1_LOC_41/Y INVX1_LOC_636/A 0.07fF
C15580 VDD INVX1_LOC_64/A -0.00fF
C15581 INVX1_LOC_20/Y INVX1_LOC_374/A 0.03fF
C15582 VDD INVX1_LOC_511/Y 0.11fF
C15583 INVX1_LOC_434/A INVX1_LOC_385/Y 0.03fF
C15584 NAND2X1_LOC_39/Y NAND2X1_LOC_16/Y 0.17fF
C15585 INVX1_LOC_76/Y NAND2X1_LOC_493/B 0.01fF
C15586 INVX1_LOC_266/A INVX1_LOC_266/Y 0.01fF
C15587 INVX1_LOC_588/Y NAND2X1_LOC_591/B 0.03fF
C15588 INVX1_LOC_546/Y INVX1_LOC_53/Y 0.01fF
C15589 INVX1_LOC_560/Y INVX1_LOC_440/A 0.01fF
C15590 INVX1_LOC_607/A INVX1_LOC_80/A 0.02fF
C15591 VDD INVX1_LOC_198/Y 0.22fF
C15592 INVX1_LOC_425/A INVX1_LOC_686/A 0.06fF
C15593 INVX1_LOC_76/Y INVX1_LOC_517/A 0.01fF
C15594 INVX1_LOC_193/Y INVX1_LOC_304/A 0.01fF
C15595 INVX1_LOC_231/Y NAND2X1_LOC_271/A 0.20fF
C15596 NAND2X1_LOC_525/Y INVX1_LOC_17/Y 0.08fF
C15597 NAND2X1_LOC_271/B INVX1_LOC_48/Y 0.04fF
C15598 INVX1_LOC_273/A NAND2X1_LOC_237/Y 0.01fF
C15599 INVX1_LOC_581/A INVX1_LOC_610/Y 0.02fF
C15600 INVX1_LOC_605/A INVX1_LOC_35/Y 0.01fF
C15601 NAND2X1_LOC_373/Y INVX1_LOC_253/Y 0.41fF
C15602 INVX1_LOC_25/Y INVX1_LOC_45/Y 0.02fF
C15603 INVX1_LOC_586/A NAND2X1_LOC_275/Y 0.23fF
C15604 NAND2X1_LOC_43/Y INVX1_LOC_45/Y 0.26fF
C15605 INVX1_LOC_11/Y INVX1_LOC_607/A 0.01fF
C15606 INVX1_LOC_53/Y INVX1_LOC_367/A 0.09fF
C15607 INVX1_LOC_245/A INVX1_LOC_638/A 0.07fF
C15608 NAND2X1_LOC_79/B INVX1_LOC_145/Y 0.70fF
C15609 NAND2X1_LOC_756/Y INVX1_LOC_99/Y 0.04fF
C15610 INVX1_LOC_238/Y INVX1_LOC_58/Y 0.00fF
C15611 INVX1_LOC_172/A INVX1_LOC_51/Y 0.03fF
C15612 INVX1_LOC_293/Y INVX1_LOC_99/Y 0.03fF
C15613 INVX1_LOC_556/Y INVX1_LOC_146/A 0.01fF
C15614 INVX1_LOC_12/Y INVX1_LOC_174/A 0.03fF
C15615 INVX1_LOC_103/A INVX1_LOC_69/Y 0.01fF
C15616 INVX1_LOC_153/A INVX1_LOC_45/Y 0.01fF
C15617 INVX1_LOC_686/A INVX1_LOC_252/Y 0.07fF
C15618 INVX1_LOC_51/Y INVX1_LOC_105/Y 0.06fF
C15619 INVX1_LOC_413/Y NAND2X1_LOC_521/Y 0.25fF
C15620 INVX1_LOC_551/Y INVX1_LOC_159/Y 0.10fF
C15621 INVX1_LOC_581/A NAND2X1_LOC_679/B 0.10fF
C15622 INVX1_LOC_395/A INVX1_LOC_199/Y 1.16fF
C15623 INVX1_LOC_24/A INVX1_LOC_338/Y 0.03fF
C15624 INVX1_LOC_578/A INVX1_LOC_419/A 0.13fF
C15625 INVX1_LOC_169/A INVX1_LOC_48/Y 0.04fF
C15626 INVX1_LOC_53/Y INVX1_LOC_669/Y 0.01fF
C15627 INVX1_LOC_307/A INVX1_LOC_7/Y 0.01fF
C15628 INVX1_LOC_560/Y INVX1_LOC_242/Y 0.02fF
C15629 INVX1_LOC_588/Y INVX1_LOC_566/A 0.04fF
C15630 INVX1_LOC_369/A NAND2X1_LOC_378/Y 0.01fF
C15631 INVX1_LOC_96/A NAND2X1_LOC_506/B 0.01fF
C15632 NAND2X1_LOC_382/a_36_24# INVX1_LOC_230/A -0.00fF
C15633 INVX1_LOC_134/Y INVX1_LOC_251/Y 0.81fF
C15634 INVX1_LOC_45/Y INVX1_LOC_96/A 0.04fF
C15635 INVX1_LOC_392/A INVX1_LOC_53/Y 0.03fF
C15636 INVX1_LOC_442/Y INVX1_LOC_7/Y 0.02fF
C15637 INVX1_LOC_596/A INVX1_LOC_50/Y 0.03fF
C15638 INVX1_LOC_117/Y INVX1_LOC_318/Y 0.34fF
C15639 INVX1_LOC_278/A INVX1_LOC_664/A 0.08fF
C15640 INVX1_LOC_412/Y INVX1_LOC_114/A 0.00fF
C15641 INVX1_LOC_20/Y NAND2X1_LOC_695/a_36_24# 0.00fF
C15642 INPUT_0 INVX1_LOC_373/Y 0.01fF
C15643 INVX1_LOC_459/Y INVX1_LOC_675/A 0.18fF
C15644 INVX1_LOC_395/A INVX1_LOC_272/A 0.01fF
C15645 NAND2X1_LOC_318/A INVX1_LOC_77/Y 0.23fF
C15646 INVX1_LOC_140/Y INVX1_LOC_26/Y 0.03fF
C15647 NAND2X1_LOC_242/A INVX1_LOC_531/Y 0.03fF
C15648 INVX1_LOC_522/Y INVX1_LOC_633/A 0.02fF
C15649 INVX1_LOC_20/Y NAND2X1_LOC_836/B 0.02fF
C15650 INVX1_LOC_21/Y NAND2X1_LOC_32/Y 0.01fF
C15651 NAND2X1_LOC_673/B INVX1_LOC_99/Y 0.06fF
C15652 INVX1_LOC_53/Y INVX1_LOC_93/Y 1.08fF
C15653 INVX1_LOC_54/Y INVX1_LOC_379/A 0.10fF
C15654 INPUT_0 NAND2X1_LOC_691/A 0.01fF
C15655 NAND2X1_LOC_545/B NAND2X1_LOC_388/A 0.03fF
C15656 INVX1_LOC_600/A INVX1_LOC_68/A 0.03fF
C15657 INVX1_LOC_504/A INVX1_LOC_50/Y 0.34fF
C15658 INVX1_LOC_85/Y NAND2X1_LOC_699/a_36_24# 0.00fF
C15659 INVX1_LOC_68/Y NAND2X1_LOC_786/B 0.04fF
C15660 INVX1_LOC_366/A INVX1_LOC_26/Y 0.13fF
C15661 INVX1_LOC_656/A INVX1_LOC_99/Y 0.01fF
C15662 NAND2X1_LOC_184/Y INVX1_LOC_367/Y 3.11fF
C15663 INVX1_LOC_442/Y INVX1_LOC_32/Y 0.07fF
C15664 NAND2X1_LOC_320/Y INVX1_LOC_31/Y 0.03fF
C15665 INVX1_LOC_54/Y INVX1_LOC_35/Y 0.27fF
C15666 INVX1_LOC_45/Y NAND2X1_LOC_627/Y 0.01fF
C15667 INVX1_LOC_586/A NAND2X1_LOC_626/Y 0.18fF
C15668 INVX1_LOC_681/A INVX1_LOC_230/Y 0.01fF
C15669 INVX1_LOC_269/Y INVX1_LOC_41/Y 0.03fF
C15670 INVX1_LOC_185/Y INVX1_LOC_475/Y 0.01fF
C15671 INVX1_LOC_134/Y INVX1_LOC_58/Y 0.10fF
C15672 INVX1_LOC_17/Y INVX1_LOC_355/Y 0.02fF
C15673 INVX1_LOC_53/Y INVX1_LOC_675/A 0.07fF
C15674 INVX1_LOC_556/A INVX1_LOC_479/A 0.03fF
C15675 NAND2X1_LOC_513/A INVX1_LOC_338/Y 0.01fF
C15676 INVX1_LOC_235/Y INVX1_LOC_247/Y 0.04fF
C15677 INVX1_LOC_678/A INVX1_LOC_641/Y 0.00fF
C15678 INVX1_LOC_261/A INVX1_LOC_59/A 0.10fF
C15679 NAND2X1_LOC_184/Y NAND2X1_LOC_251/a_36_24# 0.00fF
C15680 INVX1_LOC_84/A INVX1_LOC_242/Y 0.00fF
C15681 NAND2X1_LOC_388/A INVX1_LOC_98/Y 0.05fF
C15682 INVX1_LOC_89/Y INVX1_LOC_251/A 0.01fF
C15683 INVX1_LOC_444/Y INVX1_LOC_6/Y 0.07fF
C15684 NAND2X1_LOC_791/B INVX1_LOC_26/Y 0.81fF
C15685 INVX1_LOC_272/Y INVX1_LOC_26/Y 0.07fF
C15686 INVX1_LOC_132/Y INVX1_LOC_669/A 0.01fF
C15687 NAND2X1_LOC_376/B INVX1_LOC_145/Y 0.03fF
C15688 INVX1_LOC_490/A INVX1_LOC_48/Y 0.03fF
C15689 INVX1_LOC_257/A INVX1_LOC_35/Y 0.08fF
C15690 INVX1_LOC_63/Y NAND2X1_LOC_61/a_36_24# 0.00fF
C15691 INVX1_LOC_316/Y INVX1_LOC_58/Y 0.46fF
C15692 INVX1_LOC_317/A INVX1_LOC_48/Y 0.05fF
C15693 INVX1_LOC_202/Y INVX1_LOC_77/Y 0.01fF
C15694 INVX1_LOC_551/Y INVX1_LOC_468/A 0.09fF
C15695 INVX1_LOC_47/Y NAND2X1_LOC_673/B 0.00fF
C15696 NAND2X1_LOC_333/a_36_24# NAND2X1_LOC_720/A 0.00fF
C15697 INVX1_LOC_565/A NAND2X1_LOC_719/A 0.04fF
C15698 INVX1_LOC_304/Y INVX1_LOC_296/A 0.00fF
C15699 NAND2X1_LOC_557/B NAND2X1_LOC_673/B 0.09fF
C15700 INVX1_LOC_625/A INVX1_LOC_399/A 0.02fF
C15701 INVX1_LOC_85/Y NAND2X1_LOC_85/a_36_24# 0.00fF
C15702 INVX1_LOC_197/A INVX1_LOC_166/Y 0.00fF
C15703 INVX1_LOC_11/Y NAND2X1_LOC_259/a_36_24# 0.00fF
C15704 INVX1_LOC_384/A NAND2X1_LOC_497/a_36_24# 0.01fF
C15705 NAND2X1_LOC_274/B NAND2X1_LOC_471/a_36_24# 0.00fF
C15706 INVX1_LOC_592/Y NAND2X1_LOC_387/Y 0.02fF
C15707 NAND2X1_LOC_527/Y INVX1_LOC_234/Y 0.22fF
C15708 NAND2X1_LOC_786/B INVX1_LOC_64/A -0.01fF
C15709 NAND2X1_LOC_685/A INVX1_LOC_479/A 0.23fF
C15710 INVX1_LOC_675/A INVX1_LOC_460/Y 0.14fF
C15711 INVX1_LOC_197/A INVX1_LOC_62/Y 10.83fF
C15712 INVX1_LOC_451/A INVX1_LOC_245/A 0.03fF
C15713 INVX1_LOC_651/A NAND2X1_LOC_248/B 0.39fF
C15714 NAND2X1_LOC_274/B NAND2X1_LOC_643/a_36_24# 0.00fF
C15715 INVX1_LOC_41/Y INVX1_LOC_29/Y 0.01fF
C15716 NAND2X1_LOC_165/Y INVX1_LOC_58/Y 0.01fF
C15717 INVX1_LOC_31/Y INVX1_LOC_199/Y 0.12fF
C15718 INVX1_LOC_168/Y INVX1_LOC_189/A 0.04fF
C15719 NAND2X1_LOC_603/Y INVX1_LOC_347/A 0.02fF
C15720 INVX1_LOC_65/Y INVX1_LOC_92/A 0.01fF
C15721 INVX1_LOC_426/A INVX1_LOC_109/Y 0.07fF
C15722 INVX1_LOC_117/Y INVX1_LOC_351/A 0.00fF
C15723 INVX1_LOC_188/Y INVX1_LOC_479/A 0.07fF
C15724 NAND2X1_LOC_301/B INVX1_LOC_352/Y 4.37fF
C15725 NAND2X1_LOC_57/Y INVX1_LOC_531/Y 0.01fF
C15726 NAND2X1_LOC_409/Y INVX1_LOC_145/Y 0.72fF
C15727 INVX1_LOC_588/Y INVX1_LOC_79/A 0.04fF
C15728 INVX1_LOC_117/Y INVX1_LOC_90/Y 0.10fF
C15729 NAND2X1_LOC_274/B INVX1_LOC_46/Y 0.03fF
C15730 INVX1_LOC_62/Y NAND2X1_LOC_106/B 0.02fF
C15731 INVX1_LOC_35/Y INVX1_LOC_388/A 0.01fF
C15732 INVX1_LOC_166/A INVX1_LOC_79/A 0.06fF
C15733 INVX1_LOC_328/Y INVX1_LOC_380/Y 0.05fF
C15734 INVX1_LOC_6/Y INVX1_LOC_26/Y 1.69fF
C15735 INVX1_LOC_89/Y INVX1_LOC_652/A 0.01fF
C15736 INVX1_LOC_403/Y INVX1_LOC_479/A 0.01fF
C15737 INVX1_LOC_335/Y INVX1_LOC_636/A 0.07fF
C15738 NAND2X1_LOC_184/Y NAND2X1_LOC_843/B 0.07fF
C15739 INVX1_LOC_466/A INVX1_LOC_74/Y 0.07fF
C15740 INVX1_LOC_41/Y INVX1_LOC_470/Y 0.02fF
C15741 INVX1_LOC_367/Y NAND2X1_LOC_271/A 0.07fF
C15742 INVX1_LOC_51/Y INVX1_LOC_109/Y 0.02fF
C15743 INVX1_LOC_50/Y INVX1_LOC_346/Y 0.01fF
C15744 NAND2X1_LOC_234/Y INVX1_LOC_601/Y 0.20fF
C15745 INVX1_LOC_301/Y INVX1_LOC_100/Y 0.15fF
C15746 INVX1_LOC_26/Y NAND2X1_LOC_81/Y 0.01fF
C15747 INVX1_LOC_382/A NAND2X1_LOC_415/a_36_24# 0.00fF
C15748 INVX1_LOC_85/Y NAND2X1_LOC_86/Y 0.01fF
C15749 NAND2X1_LOC_531/Y INVX1_LOC_443/A 0.05fF
C15750 INVX1_LOC_655/A INVX1_LOC_669/A 0.20fF
C15751 INVX1_LOC_183/A NAND2X1_LOC_621/B 0.18fF
C15752 NAND2X1_LOC_790/B INVX1_LOC_586/A 0.07fF
C15753 INVX1_LOC_554/A INVX1_LOC_51/Y 0.02fF
C15754 INVX1_LOC_531/Y INVX1_LOC_79/A 0.06fF
C15755 INVX1_LOC_662/A INVX1_LOC_241/A 0.02fF
C15756 INVX1_LOC_100/Y INVX1_LOC_41/Y 2.51fF
C15757 NAND2X1_LOC_336/B INVX1_LOC_192/A 0.01fF
C15758 INVX1_LOC_435/Y INVX1_LOC_438/A 0.00fF
C15759 INVX1_LOC_75/Y INVX1_LOC_319/A 0.01fF
C15760 NAND2X1_LOC_123/B INVX1_LOC_588/A 0.03fF
C15761 INVX1_LOC_373/Y INVX1_LOC_464/Y 0.01fF
C15762 INVX1_LOC_41/Y INVX1_LOC_74/Y 0.34fF
C15763 INVX1_LOC_20/Y INVX1_LOC_560/Y 0.07fF
C15764 INVX1_LOC_400/Y NAND2X1_LOC_516/Y 0.04fF
C15765 INVX1_LOC_321/Y INVX1_LOC_297/Y 0.01fF
C15766 INVX1_LOC_139/A NAND2X1_LOC_707/A 0.00fF
C15767 INVX1_LOC_269/Y INVX1_LOC_160/Y 0.17fF
C15768 VDD NAND2X1_LOC_56/Y 0.04fF
C15769 NAND2X1_LOC_520/B INVX1_LOC_45/Y 0.02fF
C15770 INVX1_LOC_438/A INVX1_LOC_596/A 0.12fF
C15771 NAND2X1_LOC_572/a_36_24# NAND2X1_LOC_457/A 0.00fF
C15772 INVX1_LOC_301/A INVX1_LOC_129/A 0.02fF
C15773 INVX1_LOC_224/Y INVX1_LOC_80/A 0.14fF
C15774 INVX1_LOC_409/Y INVX1_LOC_360/Y 0.13fF
C15775 NAND2X1_LOC_231/A INVX1_LOC_76/Y 0.05fF
C15776 INVX1_LOC_560/Y INVX1_LOC_197/Y 0.07fF
C15777 INVX1_LOC_395/A INVX1_LOC_53/Y 0.30fF
C15778 INVX1_LOC_375/A NAND2X1_LOC_601/a_36_24# 0.00fF
C15779 NAND2X1_LOC_475/A INVX1_LOC_160/A 0.05fF
C15780 INVX1_LOC_578/A INVX1_LOC_80/A 0.14fF
C15781 INVX1_LOC_586/A INVX1_LOC_235/Y 0.10fF
C15782 INVX1_LOC_51/Y INVX1_LOC_126/Y 0.02fF
C15783 INPUT_0 INVX1_LOC_78/A 0.01fF
C15784 INPUT_0 INVX1_LOC_537/A 0.07fF
C15785 INVX1_LOC_53/Y INVX1_LOC_362/Y 0.03fF
C15786 INPUT_0 INVX1_LOC_125/A 0.06fF
C15787 NAND2X1_LOC_638/A INVX1_LOC_45/Y 0.01fF
C15788 INVX1_LOC_224/Y INVX1_LOC_11/Y 0.12fF
C15789 INVX1_LOC_20/Y INVX1_LOC_84/A 0.37fF
C15790 INVX1_LOC_317/Y INVX1_LOC_417/Y 0.00fF
C15791 INVX1_LOC_271/A INVX1_LOC_155/Y 0.02fF
C15792 INVX1_LOC_288/A INVX1_LOC_344/Y -0.00fF
C15793 INVX1_LOC_246/Y INVX1_LOC_235/Y 0.06fF
C15794 INVX1_LOC_185/A INVX1_LOC_476/A 0.02fF
C15795 INVX1_LOC_425/A NAND2X1_LOC_542/a_36_24# 0.00fF
C15796 INPUT_3 INVX1_LOC_23/Y 0.06fF
C15797 NAND2X1_LOC_249/Y INVX1_LOC_6/Y 0.03fF
C15798 INVX1_LOC_312/Y INVX1_LOC_235/Y 0.10fF
C15799 INVX1_LOC_11/Y INVX1_LOC_578/A 0.85fF
C15800 INVX1_LOC_416/Y INVX1_LOC_159/Y 0.01fF
C15801 INVX1_LOC_11/Y INVX1_LOC_557/A 0.08fF
C15802 INVX1_LOC_312/Y NAND2X1_LOC_361/a_36_24# 0.00fF
C15803 INVX1_LOC_21/Y INVX1_LOC_381/A 0.07fF
C15804 INVX1_LOC_418/Y INVX1_LOC_418/A 0.23fF
C15805 INVX1_LOC_43/A INVX1_LOC_395/A 0.09fF
C15806 INPUT_0 INVX1_LOC_421/A 0.35fF
C15807 INVX1_LOC_369/A INVX1_LOC_486/Y 0.01fF
C15808 INVX1_LOC_321/Y INVX1_LOC_76/Y 0.01fF
C15809 NAND2X1_LOC_564/a_36_24# INVX1_LOC_578/A 0.00fF
C15810 INVX1_LOC_556/Y INVX1_LOC_586/A 0.01fF
C15811 INPUT_0 INVX1_LOC_496/Y 0.04fF
C15812 INVX1_LOC_372/Y INVX1_LOC_188/Y 0.12fF
C15813 INVX1_LOC_317/Y INVX1_LOC_48/Y 0.07fF
C15814 INVX1_LOC_206/Y INVX1_LOC_419/A 0.02fF
C15815 INVX1_LOC_200/Y INVX1_LOC_66/A 0.01fF
C15816 INVX1_LOC_269/Y NAND2X1_LOC_267/A 0.04fF
C15817 INVX1_LOC_65/Y INPUT_1 0.01fF
C15818 INVX1_LOC_171/Y INVX1_LOC_35/Y 0.01fF
C15819 INVX1_LOC_315/Y NAND2X1_LOC_720/A 0.00fF
C15820 INVX1_LOC_84/A INVX1_LOC_300/A 0.04fF
C15821 INVX1_LOC_237/Y INVX1_LOC_46/Y 0.01fF
C15822 INVX1_LOC_193/A NAND2X1_LOC_332/B 0.02fF
C15823 INVX1_LOC_406/Y INVX1_LOC_453/Y 0.03fF
C15824 VDD INVX1_LOC_183/Y 0.21fF
C15825 INVX1_LOC_133/Y INVX1_LOC_614/Y 0.01fF
C15826 INVX1_LOC_459/Y INVX1_LOC_31/Y 0.06fF
C15827 NAND2X1_LOC_707/A INVX1_LOC_32/Y 0.16fF
C15828 INVX1_LOC_445/Y NAND2X1_LOC_344/B 0.42fF
C15829 INVX1_LOC_298/A NAND2X1_LOC_387/a_36_24# 0.00fF
C15830 INVX1_LOC_17/Y NAND2X1_LOC_307/A 4.20fF
C15831 NAND2X1_LOC_148/A INVX1_LOC_669/Y 0.01fF
C15832 INVX1_LOC_558/Y NAND2X1_LOC_413/Y 0.03fF
C15833 INVX1_LOC_468/Y INVX1_LOC_80/A 0.05fF
C15834 INVX1_LOC_444/Y NAND2X1_LOC_517/Y 0.06fF
C15835 INVX1_LOC_312/Y INVX1_LOC_556/Y 0.03fF
C15836 INVX1_LOC_53/Y INVX1_LOC_189/Y 0.01fF
C15837 NAND2X1_LOC_544/a_36_24# INVX1_LOC_257/A 0.00fF
C15838 INVX1_LOC_54/Y NAND2X1_LOC_336/a_36_24# 0.01fF
C15839 INVX1_LOC_548/A INVX1_LOC_53/Y 0.15fF
C15840 VDD INVX1_LOC_369/Y 0.49fF
C15841 NAND2X1_LOC_756/Y INVX1_LOC_153/A 0.07fF
C15842 INVX1_LOC_51/Y INVX1_LOC_199/Y 0.11fF
C15843 INVX1_LOC_425/A NAND2X1_LOC_542/A 0.08fF
C15844 INVX1_LOC_619/A INVX1_LOC_198/Y 0.15fF
C15845 INVX1_LOC_588/Y INVX1_LOC_632/A 0.07fF
C15846 NAND2X1_LOC_174/B INVX1_LOC_344/A 0.09fF
C15847 INPUT_3 INVX1_LOC_326/Y 0.04fF
C15848 NAND2X1_LOC_130/Y INVX1_LOC_105/A 0.00fF
C15849 INVX1_LOC_530/A INVX1_LOC_50/Y 0.00fF
C15850 NAND2X1_LOC_756/Y INVX1_LOC_96/A 0.10fF
C15851 INVX1_LOC_11/Y INVX1_LOC_468/Y 0.03fF
C15852 INVX1_LOC_53/Y INVX1_LOC_31/Y 0.13fF
C15853 NAND2X1_LOC_387/Y INVX1_LOC_12/Y 0.03fF
C15854 INVX1_LOC_266/A INVX1_LOC_199/Y 0.08fF
C15855 INVX1_LOC_382/A INVX1_LOC_489/Y 0.01fF
C15856 NAND2X1_LOC_59/a_36_24# NAND2X1_LOC_836/B 0.01fF
C15857 INVX1_LOC_236/A INVX1_LOC_492/A 0.01fF
C15858 INVX1_LOC_586/A NAND2X1_LOC_420/Y -0.07fF
C15859 INVX1_LOC_45/Y INVX1_LOC_353/A 0.08fF
C15860 INVX1_LOC_524/Y NAND2X1_LOC_790/a_36_24# 0.00fF
C15861 GATE_366 INVX1_LOC_300/Y 0.00fF
C15862 INVX1_LOC_206/Y INVX1_LOC_505/Y 0.41fF
C15863 INVX1_LOC_166/A INVX1_LOC_509/Y 0.01fF
C15864 INVX1_LOC_369/A INVX1_LOC_6/Y 1.06fF
C15865 INVX1_LOC_169/A NAND2X1_LOC_615/Y 0.02fF
C15866 NAND2X1_LOC_163/B INVX1_LOC_500/A 0.05fF
C15867 INVX1_LOC_54/Y INVX1_LOC_338/A 0.00fF
C15868 INVX1_LOC_588/Y INVX1_LOC_59/Y 0.12fF
C15869 INVX1_LOC_221/Y INVX1_LOC_661/Y 0.03fF
C15870 INVX1_LOC_318/Y INVX1_LOC_58/Y 0.01fF
C15871 INVX1_LOC_537/A INVX1_LOC_498/A 0.07fF
C15872 VDD INVX1_LOC_348/Y 0.34fF
C15873 INVX1_LOC_117/Y INVX1_LOC_98/Y 1.28fF
C15874 INVX1_LOC_544/Y INVX1_LOC_367/A 0.02fF
C15875 INVX1_LOC_442/A NAND2X1_LOC_109/a_36_24# 0.02fF
C15876 NAND2X1_LOC_507/A INVX1_LOC_35/Y 0.02fF
C15877 INVX1_LOC_393/Y INVX1_LOC_75/Y 0.04fF
C15878 INVX1_LOC_235/Y INVX1_LOC_225/Y 0.02fF
C15879 INVX1_LOC_294/A INVX1_LOC_50/Y 0.02fF
C15880 INVX1_LOC_11/Y NAND2X1_LOC_527/Y 0.00fF
C15881 INVX1_LOC_444/Y NAND2X1_LOC_294/Y 0.07fF
C15882 INVX1_LOC_114/Y INVX1_LOC_112/Y 0.92fF
C15883 VDD INVX1_LOC_240/Y 0.21fF
C15884 INVX1_LOC_336/Y INVX1_LOC_9/Y 0.05fF
C15885 INVX1_LOC_438/A NAND2X1_LOC_416/B 0.08fF
C15886 INVX1_LOC_418/Y INVX1_LOC_46/Y 0.00fF
C15887 INVX1_LOC_607/A NAND2X1_LOC_843/B 0.02fF
C15888 INVX1_LOC_134/Y NAND2X1_LOC_440/A 0.03fF
C15889 INVX1_LOC_400/Y INVX1_LOC_211/A 0.01fF
C15890 INVX1_LOC_160/Y INVX1_LOC_74/Y 0.14fF
C15891 INVX1_LOC_159/Y INVX1_LOC_46/Y 0.04fF
C15892 INVX1_LOC_89/Y INVX1_LOC_35/Y 0.06fF
C15893 NAND2X1_LOC_486/A NAND2X1_LOC_257/a_36_24# 0.00fF
C15894 INVX1_LOC_89/Y INVX1_LOC_304/A 0.02fF
C15895 INVX1_LOC_224/Y INVX1_LOC_231/Y 0.01fF
C15896 INVX1_LOC_31/Y INVX1_LOC_460/Y 0.36fF
C15897 INVX1_LOC_12/Y NAND2X1_LOC_845/B 0.01fF
C15898 INVX1_LOC_300/A INVX1_LOC_674/Y 0.10fF
C15899 INVX1_LOC_17/Y INVX1_LOC_376/A 0.05fF
C15900 INVX1_LOC_498/A INVX1_LOC_496/Y 0.03fF
C15901 NAND2X1_LOC_538/B INVX1_LOC_75/A 0.17fF
C15902 INVX1_LOC_376/Y INVX1_LOC_252/Y 0.03fF
C15903 INVX1_LOC_254/A INVX1_LOC_199/Y 0.02fF
C15904 INVX1_LOC_89/Y NAND2X1_LOC_448/B 0.06fF
C15905 INVX1_LOC_581/A INVX1_LOC_614/Y 0.02fF
C15906 INVX1_LOC_84/Y INVX1_LOC_83/A 0.06fF
C15907 INVX1_LOC_21/Y INVX1_LOC_100/Y 0.07fF
C15908 INVX1_LOC_281/Y INVX1_LOC_90/Y 0.04fF
C15909 INVX1_LOC_510/A INVX1_LOC_9/Y 0.07fF
C15910 INVX1_LOC_46/Y INVX1_LOC_212/Y 0.04fF
C15911 INVX1_LOC_255/A NAND2X1_LOC_444/A 0.15fF
C15912 NAND2X1_LOC_261/Y INVX1_LOC_443/A 0.03fF
C15913 INVX1_LOC_117/Y INVX1_LOC_338/Y 0.03fF
C15914 NAND2X1_LOC_97/B INVX1_LOC_62/Y 0.02fF
C15915 INVX1_LOC_17/Y INVX1_LOC_502/A 0.00fF
C15916 INVX1_LOC_153/Y INVX1_LOC_59/Y 0.15fF
C15917 INVX1_LOC_31/Y NAND2X1_LOC_274/Y 0.25fF
C15918 INVX1_LOC_183/A INVX1_LOC_328/A 0.02fF
C15919 NAND2X1_LOC_335/a_36_24# INVX1_LOC_92/A 0.00fF
C15920 NAND2X1_LOC_106/Y INVX1_LOC_63/Y 0.01fF
C15921 NAND2X1_LOC_280/a_36_24# INVX1_LOC_6/Y 0.00fF
C15922 NAND2X1_LOC_686/A INVX1_LOC_50/Y 0.01fF
C15923 INVX1_LOC_347/Y INVX1_LOC_359/A 0.02fF
C15924 INVX1_LOC_398/Y INVX1_LOC_531/Y 0.05fF
C15925 INVX1_LOC_90/Y NAND2X1_LOC_76/A 0.02fF
C15926 NAND2X1_LOC_109/a_36_24# INVX1_LOC_116/Y 0.00fF
C15927 INVX1_LOC_335/Y INVX1_LOC_74/Y 0.04fF
C15928 INVX1_LOC_577/Y INVX1_LOC_636/A 0.03fF
C15929 INVX1_LOC_21/Y INVX1_LOC_74/Y 0.03fF
C15930 NAND2X1_LOC_510/a_36_24# INVX1_LOC_100/Y 0.00fF
C15931 NAND2X1_LOC_179/Y INVX1_LOC_62/Y 0.01fF
C15932 INVX1_LOC_613/A INVX1_LOC_610/Y 0.12fF
C15933 INVX1_LOC_476/A INVX1_LOC_58/Y 0.00fF
C15934 NAND2X1_LOC_113/a_36_24# NAND2X1_LOC_248/B 0.00fF
C15935 INVX1_LOC_347/Y NAND2X1_LOC_466/a_36_24# 0.00fF
C15936 INVX1_LOC_153/Y INVX1_LOC_48/Y 0.03fF
C15937 INVX1_LOC_93/Y INVX1_LOC_653/A 0.03fF
C15938 NAND2X1_LOC_655/a_36_24# INVX1_LOC_74/Y 0.00fF
C15939 INVX1_LOC_50/A INVX1_LOC_93/A 0.00fF
C15940 INVX1_LOC_100/Y NAND2X1_LOC_267/A 0.07fF
C15941 NAND2X1_LOC_286/A NAND2X1_LOC_847/A 0.05fF
C15942 INVX1_LOC_62/Y INVX1_LOC_440/Y 0.12fF
C15943 NAND2X1_LOC_167/a_36_24# INVX1_LOC_255/A 0.01fF
C15944 INVX1_LOC_531/Y INVX1_LOC_48/Y 0.17fF
C15945 INVX1_LOC_492/A NAND2X1_LOC_843/B 0.02fF
C15946 INVX1_LOC_35/Y NAND2X1_LOC_544/B 0.00fF
C15947 INVX1_LOC_79/A NAND2X1_LOC_627/a_36_24# 0.01fF
C15948 INVX1_LOC_58/Y INVX1_LOC_351/A 0.00fF
C15949 INVX1_LOC_469/Y INVX1_LOC_41/Y 0.03fF
C15950 INVX1_LOC_204/Y INVX1_LOC_273/Y 0.05fF
C15951 INVX1_LOC_6/Y NAND2X1_LOC_626/Y 0.50fF
C15952 INVX1_LOC_141/Y INVX1_LOC_373/Y 0.24fF
C15953 NAND2X1_LOC_301/a_36_24# INVX1_LOC_41/Y 0.01fF
C15954 INVX1_LOC_74/Y NAND2X1_LOC_267/A 0.14fF
C15955 NAND2X1_LOC_274/B INVX1_LOC_49/Y 0.08fF
C15956 INPUT_1 INVX1_LOC_588/A 0.03fF
C15957 INVX1_LOC_352/Y INVX1_LOC_634/Y 0.07fF
C15958 INVX1_LOC_58/Y INVX1_LOC_90/Y 0.04fF
C15959 NAND2X1_LOC_181/A INVX1_LOC_41/Y 0.03fF
C15960 INVX1_LOC_79/A INVX1_LOC_411/Y 0.03fF
C15961 INVX1_LOC_662/A INVX1_LOC_643/Y 0.03fF
C15962 NAND2X1_LOC_123/B INVX1_LOC_63/Y 0.40fF
C15963 NAND2X1_LOC_346/a_36_24# INVX1_LOC_280/A 0.02fF
C15964 INVX1_LOC_641/A NAND2X1_LOC_451/B 0.03fF
C15965 INVX1_LOC_382/A INVX1_LOC_443/A 0.19fF
C15966 NAND2X1_LOC_334/A INVX1_LOC_505/Y 0.03fF
C15967 INVX1_LOC_601/Y INVX1_LOC_623/A 0.01fF
C15968 INVX1_LOC_77/A INVX1_LOC_41/Y 0.03fF
C15969 INPUT_0 NAND2X1_LOC_45/Y 0.03fF
C15970 INVX1_LOC_346/A INVX1_LOC_348/Y 0.01fF
C15971 INVX1_LOC_62/Y INVX1_LOC_485/Y 0.10fF
C15972 INVX1_LOC_409/Y INVX1_LOC_45/Y 0.03fF
C15973 INVX1_LOC_63/Y NAND2X1_LOC_263/a_36_24# 0.00fF
C15974 VDD INVX1_LOC_428/A 0.00fF
C15975 INVX1_LOC_79/A INVX1_LOC_41/Y 0.09fF
C15976 NAND2X1_LOC_45/Y NAND2X1_LOC_24/a_36_24# 0.00fF
C15977 INVX1_LOC_317/Y NAND2X1_LOC_370/a_36_24# 0.00fF
C15978 VDD INVX1_LOC_33/Y 0.77fF
C15979 INVX1_LOC_63/Y INVX1_LOC_270/Y 0.07fF
C15980 INVX1_LOC_253/Y INVX1_LOC_92/A 0.01fF
C15981 INPUT_0 INVX1_LOC_36/A 0.01fF
C15982 INPUT_0 NAND2X1_LOC_498/Y 0.07fF
C15983 INPUT_0 INVX1_LOC_570/A 0.03fF
C15984 INVX1_LOC_562/A INVX1_LOC_340/Y 0.05fF
C15985 INVX1_LOC_63/Y INVX1_LOC_92/A 0.07fF
C15986 INVX1_LOC_584/A INVX1_LOC_288/A 0.02fF
C15987 NAND2X1_LOC_516/Y NAND2X1_LOC_498/Y 0.08fF
C15988 NAND2X1_LOC_843/B NAND2X1_LOC_287/a_36_24# 0.00fF
C15989 INVX1_LOC_555/Y INVX1_LOC_395/A 0.04fF
C15990 INVX1_LOC_74/A NAND2X1_LOC_70/a_36_24# 0.02fF
C15991 INVX1_LOC_206/Y NAND2X1_LOC_388/a_36_24# 0.00fF
C15992 INVX1_LOC_26/Y INVX1_LOC_636/A 0.24fF
C15993 VDD INVX1_LOC_489/Y 0.22fF
C15994 VDD INVX1_LOC_558/Y 0.29fF
C15995 INPUT_0 INVX1_LOC_377/Y 0.70fF
C15996 INVX1_LOC_65/Y INVX1_LOC_134/A 0.14fF
C15997 INVX1_LOC_459/Y INVX1_LOC_51/Y 0.92fF
C15998 INVX1_LOC_68/Y INVX1_LOC_45/Y 0.06fF
C15999 INVX1_LOC_233/Y INVX1_LOC_45/Y 0.01fF
C16000 INVX1_LOC_206/Y INVX1_LOC_80/A 3.05fF
C16001 INVX1_LOC_206/Y NAND2X1_LOC_768/A 0.00fF
C16002 INVX1_LOC_17/Y INVX1_LOC_388/Y 0.05fF
C16003 INVX1_LOC_567/A INVX1_LOC_556/Y 0.00fF
C16004 NAND2X1_LOC_88/B INVX1_LOC_177/Y 0.01fF
C16005 INVX1_LOC_7/A INVX1_LOC_8/Y 0.05fF
C16006 INVX1_LOC_395/A NAND2X1_LOC_148/A 0.03fF
C16007 INVX1_LOC_91/Y NAND2X1_LOC_98/B 0.04fF
C16008 INVX1_LOC_193/A INVX1_LOC_301/A 0.00fF
C16009 INVX1_LOC_404/Y NAND2X1_LOC_416/Y 0.04fF
C16010 NAND2X1_LOC_780/B INVX1_LOC_35/Y 0.01fF
C16011 INPUT_0 INVX1_LOC_99/Y 7.09fF
C16012 INVX1_LOC_224/Y INVX1_LOC_367/Y 0.00fF
C16013 INVX1_LOC_130/Y INVX1_LOC_412/A 0.01fF
C16014 INVX1_LOC_584/A INVX1_LOC_145/Y 0.03fF
C16015 INVX1_LOC_250/Y INVX1_LOC_45/Y 0.03fF
C16016 INVX1_LOC_133/Y INVX1_LOC_633/A 0.00fF
C16017 INVX1_LOC_53/Y NAND2X1_LOC_794/a_36_24# 0.01fF
C16018 INVX1_LOC_53/Y INVX1_LOC_51/Y 0.23fF
C16019 INVX1_LOC_45/Y NAND2X1_LOC_302/A 0.08fF
C16020 VDD INVX1_LOC_359/Y 0.21fF
C16021 INVX1_LOC_11/Y INVX1_LOC_206/Y 0.12fF
C16022 INVX1_LOC_45/Y INVX1_LOC_600/A 0.03fF
C16023 INVX1_LOC_435/A INVX1_LOC_490/Y 0.44fF
C16024 INVX1_LOC_590/Y INVX1_LOC_99/Y 0.02fF
C16025 INVX1_LOC_235/Y INVX1_LOC_486/Y 0.16fF
C16026 INVX1_LOC_565/A INVX1_LOC_586/A 0.00fF
C16027 NAND2X1_LOC_719/a_36_24# INVX1_LOC_674/A 0.00fF
C16028 INVX1_LOC_588/Y INVX1_LOC_561/Y 0.20fF
C16029 INVX1_LOC_266/A INVX1_LOC_53/Y 0.78fF
C16030 NAND2X1_LOC_820/Y NAND2X1_LOC_820/A 0.01fF
C16031 INVX1_LOC_137/A INVX1_LOC_35/Y 0.01fF
C16032 INVX1_LOC_217/Y NAND2X1_LOC_482/Y 0.12fF
C16033 NAND2X1_LOC_537/A INVX1_LOC_199/Y 0.06fF
C16034 VDD INVX1_LOC_187/Y 0.22fF
C16035 VDD NAND2X1_LOC_284/A -0.00fF
C16036 INVX1_LOC_80/A INVX1_LOC_686/A 0.39fF
C16037 INVX1_LOC_76/Y INVX1_LOC_549/Y 0.35fF
C16038 NAND2X1_LOC_24/Y INVX1_LOC_12/Y 0.03fF
C16039 INVX1_LOC_80/Y INVX1_LOC_80/A 0.01fF
C16040 INVX1_LOC_81/Y INVX1_LOC_366/A 0.00fF
C16041 INVX1_LOC_444/Y INVX1_LOC_381/A 0.07fF
C16042 INVX1_LOC_51/Y INVX1_LOC_460/Y 0.03fF
C16043 INVX1_LOC_186/A INVX1_LOC_522/Y 0.02fF
C16044 INVX1_LOC_402/A INVX1_LOC_367/A 0.01fF
C16045 INVX1_LOC_238/Y INVX1_LOC_520/Y 1.59fF
C16046 INPUT_0 INVX1_LOC_47/Y 0.15fF
C16047 INVX1_LOC_11/Y INVX1_LOC_242/A 0.07fF
C16048 VDD NAND2X1_LOC_768/B 0.02fF
C16049 NAND2X1_LOC_694/a_36_24# INVX1_LOC_513/A 0.00fF
C16050 INVX1_LOC_17/Y NAND2X1_LOC_840/a_36_24# 0.01fF
C16051 NAND2X1_LOC_516/Y INVX1_LOC_47/Y 0.07fF
C16052 INVX1_LOC_558/A NAND2X1_LOC_225/a_36_24# 0.00fF
C16053 INVX1_LOC_45/Y INVX1_LOC_484/A 0.01fF
C16054 INVX1_LOC_11/Y INVX1_LOC_686/A 0.07fF
C16055 NAND2X1_LOC_383/Y INVX1_LOC_31/Y 0.58fF
C16056 INVX1_LOC_424/A INVX1_LOC_405/Y 0.01fF
C16057 INVX1_LOC_662/Y INVX1_LOC_651/A 0.03fF
C16058 INVX1_LOC_172/Y INVX1_LOC_46/Y 0.02fF
C16059 INVX1_LOC_395/A INVX1_LOC_662/A 0.08fF
C16060 NAND2X1_LOC_250/Y INVX1_LOC_679/Y 0.15fF
C16061 INVX1_LOC_537/A INVX1_LOC_145/Y 0.07fF
C16062 NAND2X1_LOC_180/B INVX1_LOC_66/A 0.14fF
C16063 INVX1_LOC_596/A INVX1_LOC_117/Y 0.00fF
C16064 INVX1_LOC_607/Y INVX1_LOC_99/Y 0.13fF
C16065 INVX1_LOC_427/A INVX1_LOC_63/Y 0.03fF
C16066 INPUT_0 INVX1_LOC_119/Y 0.03fF
C16067 INVX1_LOC_20/Y NAND2X1_LOC_285/a_36_24# 0.00fF
C16068 INVX1_LOC_11/Y INVX1_LOC_14/A 0.03fF
C16069 INVX1_LOC_427/Y INVX1_LOC_428/Y 0.09fF
C16070 NAND2X1_LOC_13/Y INVX1_LOC_199/Y 0.04fF
C16071 INVX1_LOC_584/Y INVX1_LOC_500/A 0.49fF
C16072 INVX1_LOC_670/Y INPUT_1 0.08fF
C16073 INVX1_LOC_251/Y INVX1_LOC_98/Y 0.04fF
C16074 INVX1_LOC_51/Y NAND2X1_LOC_406/B 0.08fF
C16075 INVX1_LOC_412/Y INVX1_LOC_62/Y 0.03fF
C16076 INVX1_LOC_419/Y INVX1_LOC_545/A 0.00fF
C16077 INVX1_LOC_321/A INVX1_LOC_9/Y 0.06fF
C16078 NAND2X1_LOC_516/Y INVX1_LOC_119/Y 0.08fF
C16079 NAND2X1_LOC_76/A INVX1_LOC_98/Y 0.04fF
C16080 INVX1_LOC_35/Y INVX1_LOC_194/Y 0.01fF
C16081 INVX1_LOC_581/A INVX1_LOC_633/A 0.03fF
C16082 INVX1_LOC_159/Y INVX1_LOC_349/Y 0.00fF
C16083 INVX1_LOC_117/Y INVX1_LOC_504/A 0.07fF
C16084 VDD NAND2X1_LOC_832/A -0.00fF
C16085 INVX1_LOC_315/Y INVX1_LOC_79/A 0.03fF
C16086 NAND2X1_LOC_411/Y INVX1_LOC_66/A 0.01fF
C16087 INVX1_LOC_374/A NAND2X1_LOC_123/B 0.40fF
C16088 INVX1_LOC_468/Y INVX1_LOC_374/Y 0.01fF
C16089 INVX1_LOC_54/Y INVX1_LOC_350/A 0.00fF
C16090 VDD INVX1_LOC_443/A 5.78fF
C16091 INVX1_LOC_478/Y NAND2X1_LOC_615/B 0.06fF
C16092 INVX1_LOC_421/A INVX1_LOC_145/Y 0.01fF
C16093 INVX1_LOC_617/Y INVX1_LOC_9/Y 0.07fF
C16094 NAND2X1_LOC_152/B NAND2X1_LOC_846/B 0.18fF
C16095 INVX1_LOC_21/Y NAND2X1_LOC_181/A 0.64fF
C16096 INVX1_LOC_602/A INVX1_LOC_622/A 0.01fF
C16097 INVX1_LOC_145/Y INVX1_LOC_496/Y 0.03fF
C16098 INVX1_LOC_679/A INVX1_LOC_283/A 0.01fF
C16099 INVX1_LOC_224/Y INVX1_LOC_625/Y 0.00fF
C16100 INVX1_LOC_381/A INVX1_LOC_26/Y 0.07fF
C16101 INVX1_LOC_20/Y INVX1_LOC_106/Y 0.01fF
C16102 INVX1_LOC_255/Y INVX1_LOC_74/Y 1.06fF
C16103 NAND2X1_LOC_770/B INVX1_LOC_598/A 0.11fF
C16104 INVX1_LOC_625/A NAND2X1_LOC_388/A 0.00fF
C16105 INVX1_LOC_679/Y INVX1_LOC_63/Y 0.05fF
C16106 INVX1_LOC_318/Y INVX1_LOC_245/A 0.21fF
C16107 INVX1_LOC_417/Y INVX1_LOC_411/Y 0.24fF
C16108 INVX1_LOC_47/Y NAND2X1_LOC_686/a_36_24# 0.00fF
C16109 INVX1_LOC_206/Y INVX1_LOC_231/Y 0.08fF
C16110 INVX1_LOC_542/A INVX1_LOC_479/A 0.11fF
C16111 INVX1_LOC_556/Y INVX1_LOC_6/Y 0.18fF
C16112 INVX1_LOC_578/A INVX1_LOC_625/Y 0.07fF
C16113 NAND2X1_LOC_184/Y INVX1_LOC_671/A 0.00fF
C16114 INVX1_LOC_81/Y INVX1_LOC_6/Y 0.00fF
C16115 INVX1_LOC_530/Y NAND2X1_LOC_617/a_36_24# 0.01fF
C16116 INVX1_LOC_287/Y INVX1_LOC_203/A 0.04fF
C16117 INVX1_LOC_89/Y INVX1_LOC_360/A 0.02fF
C16118 INVX1_LOC_58/Y INVX1_LOC_98/Y 0.59fF
C16119 INVX1_LOC_318/A NAND2X1_LOC_389/a_36_24# 0.02fF
C16120 NAND2X1_LOC_173/Y INVX1_LOC_354/A 0.06fF
C16121 INVX1_LOC_35/Y INVX1_LOC_44/Y 2.23fF
C16122 INVX1_LOC_253/Y INPUT_1 0.02fF
C16123 NAND2X1_LOC_231/B INVX1_LOC_94/A 0.39fF
C16124 INVX1_LOC_69/Y NAND2X1_LOC_444/A 0.01fF
C16125 INVX1_LOC_21/Y INVX1_LOC_79/A 0.24fF
C16126 INVX1_LOC_63/Y INPUT_1 0.06fF
C16127 INVX1_LOC_632/A INVX1_LOC_41/Y 0.07fF
C16128 INVX1_LOC_95/A INVX1_LOC_50/Y 0.01fF
C16129 INVX1_LOC_54/Y INVX1_LOC_507/Y 0.19fF
C16130 INVX1_LOC_444/Y INVX1_LOC_100/Y 0.07fF
C16131 INVX1_LOC_561/A INVX1_LOC_675/A 0.02fF
C16132 INVX1_LOC_44/Y INVX1_LOC_620/A 0.07fF
C16133 INVX1_LOC_63/Y INVX1_LOC_292/Y 0.04fF
C16134 INVX1_LOC_41/Y INVX1_LOC_59/Y 0.15fF
C16135 INVX1_LOC_199/Y INVX1_LOC_361/A 0.08fF
C16136 INVX1_LOC_442/Y INVX1_LOC_75/Y 0.07fF
C16137 INVX1_LOC_522/Y INVX1_LOC_611/A 0.03fF
C16138 INVX1_LOC_159/Y INVX1_LOC_17/A 0.00fF
C16139 NAND2X1_LOC_789/A INVX1_LOC_26/Y 0.07fF
C16140 INVX1_LOC_58/Y INVX1_LOC_338/Y 0.07fF
C16141 INVX1_LOC_99/Y INVX1_LOC_211/A 0.10fF
C16142 INVX1_LOC_31/Y INVX1_LOC_653/A 0.09fF
C16143 INVX1_LOC_396/A INVX1_LOC_531/Y 0.04fF
C16144 INVX1_LOC_63/Y INVX1_LOC_284/Y 0.01fF
C16145 INVX1_LOC_41/Y INVX1_LOC_48/Y 7.29fF
C16146 INVX1_LOC_93/Y NAND2X1_LOC_545/A 0.04fF
C16147 INVX1_LOC_615/A INVX1_LOC_616/Y 0.00fF
C16148 INVX1_LOC_399/A INVX1_LOC_63/Y 0.16fF
C16149 INVX1_LOC_479/A INVX1_LOC_259/Y 0.00fF
C16150 NAND2X1_LOC_285/a_36_24# INVX1_LOC_655/A 0.01fF
C16151 INVX1_LOC_93/Y INVX1_LOC_653/Y 0.24fF
C16152 INVX1_LOC_50/Y INVX1_LOC_588/A 4.32fF
C16153 INVX1_LOC_261/Y INVX1_LOC_660/Y 0.91fF
C16154 VDD INVX1_LOC_180/Y 0.34fF
C16155 INVX1_LOC_93/Y INVX1_LOC_666/Y 0.14fF
C16156 NAND2X1_LOC_707/B INVX1_LOC_479/A 0.02fF
C16157 NAND2X1_LOC_164/Y INVX1_LOC_275/A 2.80fF
C16158 INVX1_LOC_183/Y NAND2X1_LOC_80/a_36_24# 0.00fF
C16159 INVX1_LOC_49/Y INVX1_LOC_468/A 0.04fF
C16160 INVX1_LOC_589/Y INVX1_LOC_211/A 0.09fF
C16161 INVX1_LOC_90/Y INVX1_LOC_245/A 0.04fF
C16162 NAND2X1_LOC_333/B NAND2X1_LOC_98/B 0.02fF
C16163 NAND2X1_LOC_493/a_36_24# INVX1_LOC_319/A 0.01fF
C16164 INVX1_LOC_106/Y INVX1_LOC_655/A 0.02fF
C16165 NAND2X1_LOC_750/Y VDD 0.14fF
C16166 INVX1_LOC_47/Y INVX1_LOC_211/A 0.15fF
C16167 INVX1_LOC_47/Y INVX1_LOC_464/Y 0.11fF
C16168 INVX1_LOC_100/Y INVX1_LOC_128/Y 0.01fF
C16169 VDD INVX1_LOC_420/Y 0.45fF
C16170 INVX1_LOC_100/Y INVX1_LOC_26/Y 0.07fF
C16171 INVX1_LOC_47/Y INVX1_LOC_64/Y 0.15fF
C16172 VDD NAND2X1_LOC_241/B 0.05fF
C16173 VDD INVX1_LOC_606/Y 0.21fF
C16174 INPUT_0 NAND2X1_LOC_475/A 0.03fF
C16175 INVX1_LOC_390/A INVX1_LOC_666/Y 0.03fF
C16176 NAND2X1_LOC_750/Y INVX1_LOC_228/Y 0.00fF
C16177 INVX1_LOC_26/Y INVX1_LOC_74/Y 0.13fF
C16178 INVX1_LOC_347/Y INVX1_LOC_634/Y 0.09fF
C16179 INVX1_LOC_41/Y INVX1_LOC_472/Y 0.02fF
C16180 INVX1_LOC_577/Y NAND2X1_LOC_591/B 0.00fF
C16181 INVX1_LOC_479/A INVX1_LOC_114/A 0.08fF
C16182 INVX1_LOC_629/A INVX1_LOC_255/Y 0.14fF
C16183 INVX1_LOC_491/A NAND2X1_LOC_646/B 0.06fF
C16184 VDD NAND2X1_LOC_261/Y 0.20fF
C16185 NAND2X1_LOC_475/A INVX1_LOC_286/A 0.15fF
C16186 INVX1_LOC_445/Y INVX1_LOC_446/Y 0.02fF
C16187 VDD NAND2X1_LOC_173/Y 0.11fF
C16188 INVX1_LOC_393/Y INVX1_LOC_578/A 0.09fF
C16189 INVX1_LOC_317/Y NAND2X1_LOC_312/a_36_24# 0.00fF
C16190 INVX1_LOC_554/A NAND2X1_LOC_152/B 0.00fF
C16191 INVX1_LOC_197/A INVX1_LOC_638/A 0.03fF
C16192 NAND2X1_LOC_45/Y INVX1_LOC_384/A 0.16fF
C16193 INVX1_LOC_445/Y INVX1_LOC_384/A 0.13fF
C16194 INVX1_LOC_206/Y INVX1_LOC_566/Y 0.03fF
C16195 NAND2X1_LOC_498/Y INVX1_LOC_384/A 0.03fF
C16196 INVX1_LOC_288/A INVX1_LOC_114/Y 0.03fF
C16197 INVX1_LOC_442/A NAND2X1_LOC_180/B 0.02fF
C16198 NAND2X1_LOC_571/a_36_24# INVX1_LOC_434/A 0.00fF
C16199 VDD NAND2X1_LOC_413/Y 0.28fF
C16200 INVX1_LOC_21/Y INVX1_LOC_191/Y 0.02fF
C16201 VDD INVX1_LOC_44/A -0.00fF
C16202 NAND2X1_LOC_174/B INVX1_LOC_638/A 0.11fF
C16203 INVX1_LOC_560/A INVX1_LOC_320/A 0.15fF
C16204 NAND2X1_LOC_475/A NAND2X1_LOC_123/A 0.02fF
C16205 INVX1_LOC_446/A INPUT_1 0.46fF
C16206 NAND2X1_LOC_45/Y INVX1_LOC_145/Y 0.04fF
C16207 NAND2X1_LOC_591/Y INVX1_LOC_638/A 0.07fF
C16208 INVX1_LOC_577/Y INVX1_LOC_566/A 0.05fF
C16209 INVX1_LOC_428/A NAND2X1_LOC_486/a_36_24# 0.00fF
C16210 INVX1_LOC_86/Y INVX1_LOC_181/A 0.01fF
C16211 NAND2X1_LOC_243/A INVX1_LOC_180/Y 0.03fF
C16212 NAND2X1_LOC_56/Y INVX1_LOC_45/Y 0.02fF
C16213 INVX1_LOC_448/A NAND2X1_LOC_498/Y 0.75fF
C16214 INVX1_LOC_384/A INVX1_LOC_377/Y 0.13fF
C16215 INVX1_LOC_118/Y INVX1_LOC_35/Y 0.01fF
C16216 INVX1_LOC_628/A INVX1_LOC_255/Y 0.00fF
C16217 INVX1_LOC_206/Y INVX1_LOC_313/Y 0.01fF
C16218 INVX1_LOC_80/A INVX1_LOC_94/A 0.08fF
C16219 NAND2X1_LOC_475/A INVX1_LOC_527/Y 0.00fF
C16220 INVX1_LOC_446/Y INVX1_LOC_99/Y 0.07fF
C16221 VDD INVX1_LOC_341/Y 0.21fF
C16222 INVX1_LOC_55/Y INVX1_LOC_59/A 0.04fF
C16223 INVX1_LOC_310/Y INVX1_LOC_366/A 0.00fF
C16224 INVX1_LOC_288/A INVX1_LOC_99/Y 0.07fF
C16225 NAND2X1_LOC_789/B INVX1_LOC_86/Y 0.01fF
C16226 INVX1_LOC_224/Y INVX1_LOC_361/Y 0.03fF
C16227 INPUT_6 INVX1_LOC_3/A 0.02fF
C16228 INVX1_LOC_96/Y INVX1_LOC_35/Y 0.39fF
C16229 NAND2X1_LOC_79/B INVX1_LOC_600/Y 0.02fF
C16230 INVX1_LOC_564/Y NAND2X1_LOC_720/A 0.01fF
C16231 INVX1_LOC_142/A INVX1_LOC_145/Y 0.00fF
C16232 INVX1_LOC_384/A INVX1_LOC_99/Y 0.09fF
C16233 INVX1_LOC_578/A INVX1_LOC_361/Y 0.07fF
C16234 INVX1_LOC_490/Y INVX1_LOC_93/Y 0.03fF
C16235 INVX1_LOC_448/A INVX1_LOC_377/Y 0.02fF
C16236 INVX1_LOC_393/A INVX1_LOC_665/Y 0.01fF
C16237 INVX1_LOC_52/Y INVX1_LOC_89/Y 0.01fF
C16238 NAND2X1_LOC_332/B INVX1_LOC_125/A 0.34fF
C16239 NAND2X1_LOC_180/B INVX1_LOC_116/Y 0.05fF
C16240 INVX1_LOC_11/Y INVX1_LOC_94/A 0.01fF
C16241 NAND2X1_LOC_93/Y INVX1_LOC_95/A 0.01fF
C16242 NAND2X1_LOC_391/B INVX1_LOC_230/A 0.00fF
C16243 INVX1_LOC_160/Y INVX1_LOC_48/Y 0.24fF
C16244 INVX1_LOC_586/A INVX1_LOC_304/Y 0.05fF
C16245 INVX1_LOC_409/A INVX1_LOC_49/Y 0.19fF
C16246 INVX1_LOC_255/Y INVX1_LOC_469/Y 1.01fF
C16247 INVX1_LOC_412/Y INVX1_LOC_624/Y 0.00fF
C16248 INVX1_LOC_445/Y INVX1_LOC_433/A 0.02fF
C16249 INVX1_LOC_26/Y NAND2X1_LOC_591/B 0.01fF
C16250 NAND2X1_LOC_786/B INVX1_LOC_180/Y 0.05fF
C16251 INVX1_LOC_312/A INVX1_LOC_379/A 0.01fF
C16252 INVX1_LOC_335/Y INVX1_LOC_632/A 0.07fF
C16253 INVX1_LOC_11/Y INVX1_LOC_654/A 0.01fF
C16254 INVX1_LOC_676/Y INVX1_LOC_677/A 0.00fF
C16255 INVX1_LOC_586/A NAND2X1_LOC_444/A 0.01fF
C16256 INVX1_LOC_65/Y NAND2X1_LOC_388/A 0.02fF
C16257 INVX1_LOC_21/Y INVX1_LOC_509/Y 0.01fF
C16258 NAND2X1_LOC_773/A INVX1_LOC_198/Y 0.02fF
C16259 INVX1_LOC_101/Y NAND2X1_LOC_106/B 0.00fF
C16260 NAND2X1_LOC_504/a_36_24# NAND2X1_LOC_318/A 0.01fF
C16261 INVX1_LOC_35/Y NAND2X1_LOC_837/a_36_24# 0.01fF
C16262 INVX1_LOC_413/Y INVX1_LOC_69/Y 0.07fF
C16263 INVX1_LOC_435/Y INVX1_LOC_58/Y 0.03fF
C16264 INVX1_LOC_553/Y INVX1_LOC_9/Y 0.14fF
C16265 NAND2X1_LOC_249/Y INVX1_LOC_100/Y 0.07fF
C16266 INPUT_0 INVX1_LOC_15/Y 0.11fF
C16267 INVX1_LOC_288/A INVX1_LOC_47/Y 0.45fF
C16268 INVX1_LOC_312/Y INVX1_LOC_304/Y 0.03fF
C16269 NAND2X1_LOC_391/A INVX1_LOC_304/A 0.00fF
C16270 INVX1_LOC_54/Y INVX1_LOC_522/Y 0.07fF
C16271 NAND2X1_LOC_242/A INVX1_LOC_26/Y 0.20fF
C16272 VDD INVX1_LOC_245/Y 0.24fF
C16273 INVX1_LOC_410/A INVX1_LOC_173/A 0.12fF
C16274 INVX1_LOC_93/Y INVX1_LOC_353/Y 0.05fF
C16275 INVX1_LOC_410/Y INVX1_LOC_9/Y 0.10fF
C16276 NAND2X1_LOC_26/a_36_24# INVX1_LOC_204/Y 0.00fF
C16277 NAND2X1_LOC_750/Y NAND2X1_LOC_786/B 0.00fF
C16278 NAND2X1_LOC_318/B INVX1_LOC_178/A 0.02fF
C16279 INVX1_LOC_21/Y INVX1_LOC_59/Y 0.02fF
C16280 NAND2X1_LOC_710/A INVX1_LOC_166/A 0.02fF
C16281 INVX1_LOC_99/Y INVX1_LOC_145/Y 2.54fF
C16282 INVX1_LOC_384/A INVX1_LOC_47/Y 0.07fF
C16283 INVX1_LOC_188/Y NAND2X1_LOC_432/Y 0.08fF
C16284 INVX1_LOC_40/Y INVX1_LOC_69/A 0.02fF
C16285 VDD NAND2X1_LOC_488/Y 0.04fF
C16286 NAND2X1_LOC_673/B INVX1_LOC_600/A 0.00fF
C16287 INVX1_LOC_544/Y INVX1_LOC_51/Y 0.01fF
C16288 NAND2X1_LOC_591/a_36_24# NAND2X1_LOC_591/Y 0.02fF
C16289 INVX1_LOC_451/A NAND2X1_LOC_416/Y 0.54fF
C16290 INVX1_LOC_400/Y INVX1_LOC_242/Y 0.03fF
C16291 NAND2X1_LOC_180/B INVX1_LOC_255/A 0.04fF
C16292 INVX1_LOC_324/Y INVX1_LOC_328/A 0.12fF
C16293 INVX1_LOC_42/Y NAND2X1_LOC_81/a_36_24# 0.00fF
C16294 INVX1_LOC_670/Y INVX1_LOC_50/Y 0.01fF
C16295 INVX1_LOC_560/A INVX1_LOC_100/Y 0.14fF
C16296 INVX1_LOC_522/A INVX1_LOC_514/Y 0.00fF
C16297 NAND2X1_LOC_563/a_36_24# INVX1_LOC_386/Y 0.01fF
C16298 VDD INVX1_LOC_441/A 0.00fF
C16299 INVX1_LOC_117/Y INVX1_LOC_530/A 0.01fF
C16300 INVX1_LOC_21/Y INVX1_LOC_48/Y 3.23fF
C16301 VDD INVX1_LOC_645/Y 0.15fF
C16302 INVX1_LOC_51/Y INVX1_LOC_662/A 0.03fF
C16303 INVX1_LOC_449/A INVX1_LOC_46/Y 0.01fF
C16304 INVX1_LOC_558/A INVX1_LOC_518/A 0.01fF
C16305 NAND2X1_LOC_457/A NAND2X1_LOC_528/Y 0.00fF
C16306 INVX1_LOC_206/Y NAND2X1_LOC_843/B 0.01fF
C16307 INVX1_LOC_566/Y NAND2X1_LOC_334/A 0.05fF
C16308 INVX1_LOC_410/Y INVX1_LOC_62/Y 0.03fF
C16309 INVX1_LOC_581/Y INVX1_LOC_583/A 0.02fF
C16310 INVX1_LOC_288/A INVX1_LOC_119/Y 0.00fF
C16311 INVX1_LOC_80/A NAND2X1_LOC_542/A 0.02fF
C16312 INVX1_LOC_139/A INVX1_LOC_148/Y 0.37fF
C16313 NAND2X1_LOC_314/a_36_24# INVX1_LOC_479/A 0.01fF
C16314 INVX1_LOC_310/Y INVX1_LOC_6/Y 0.02fF
C16315 INVX1_LOC_25/Y INVX1_LOC_298/A 0.00fF
C16316 NAND2X1_LOC_775/B INVX1_LOC_349/A 0.10fF
C16317 INVX1_LOC_560/A INVX1_LOC_74/Y 0.07fF
C16318 INVX1_LOC_45/Y INVX1_LOC_369/Y 0.21fF
C16319 INVX1_LOC_59/Y NAND2X1_LOC_267/A 0.02fF
C16320 INVX1_LOC_565/A INVX1_LOC_6/Y 0.00fF
C16321 INVX1_LOC_448/A INVX1_LOC_47/Y 0.07fF
C16322 INVX1_LOC_17/Y INVX1_LOC_230/Y 0.07fF
C16323 INVX1_LOC_648/Y NAND2X1_LOC_843/B 0.01fF
C16324 INVX1_LOC_387/Y NAND2X1_LOC_595/Y 0.13fF
C16325 INVX1_LOC_412/A INVX1_LOC_75/Y 0.02fF
C16326 INVX1_LOC_577/Y INVX1_LOC_79/A 0.03fF
C16327 INVX1_LOC_137/A NAND2X1_LOC_647/a_36_24# 0.00fF
C16328 INVX1_LOC_384/A INVX1_LOC_119/Y 0.02fF
C16329 INVX1_LOC_50/Y NAND2X1_LOC_646/A 0.00fF
C16330 INVX1_LOC_89/Y INVX1_LOC_115/Y 0.03fF
C16331 INVX1_LOC_395/A INVX1_LOC_666/Y 0.18fF
C16332 INVX1_LOC_566/A INVX1_LOC_26/Y 0.23fF
C16333 INVX1_LOC_547/Y INVX1_LOC_479/A 0.09fF
C16334 INVX1_LOC_20/Y INVX1_LOC_373/Y 0.00fF
C16335 INVX1_LOC_49/Y INVX1_LOC_377/A 0.04fF
C16336 INVX1_LOC_523/Y INVX1_LOC_35/Y 0.21fF
C16337 INVX1_LOC_196/A INVX1_LOC_491/A 0.06fF
C16338 INVX1_LOC_47/Y INVX1_LOC_145/Y 0.78fF
C16339 NAND2X1_LOC_267/A INVX1_LOC_48/Y 0.86fF
C16340 INVX1_LOC_288/Y INVX1_LOC_69/Y 0.03fF
C16341 INVX1_LOC_80/A INVX1_LOC_376/Y 0.08fF
C16342 INVX1_LOC_49/Y NAND2X1_LOC_595/Y 0.05fF
C16343 NAND2X1_LOC_557/B INVX1_LOC_145/Y 0.21fF
C16344 INVX1_LOC_372/Y INVX1_LOC_114/A 0.05fF
C16345 INVX1_LOC_649/Y INVX1_LOC_667/Y 0.01fF
C16346 INVX1_LOC_117/Y INVX1_LOC_520/A 0.02fF
C16347 NAND2X1_LOC_785/a_36_24# INVX1_LOC_63/Y 0.00fF
C16348 INPUT_3 INVX1_LOC_369/Y 0.00fF
C16349 INVX1_LOC_573/Y INVX1_LOC_332/Y 0.02fF
C16350 INVX1_LOC_555/A INVX1_LOC_48/Y 0.03fF
C16351 NAND2X1_LOC_843/B INVX1_LOC_242/A 0.03fF
C16352 INVX1_LOC_11/Y NAND2X1_LOC_542/A 0.07fF
C16353 INVX1_LOC_255/A NAND2X1_LOC_444/a_36_24# 0.01fF
C16354 INVX1_LOC_428/Y INVX1_LOC_63/Y 0.03fF
C16355 INVX1_LOC_49/Y INVX1_LOC_352/Y 0.02fF
C16356 INVX1_LOC_93/Y INVX1_LOC_18/Y 0.01fF
C16357 INVX1_LOC_188/A INVX1_LOC_259/Y 0.09fF
C16358 INVX1_LOC_100/Y INVX1_LOC_369/A 0.03fF
C16359 INVX1_LOC_123/A NAND2X1_LOC_133/a_36_24# 0.00fF
C16360 INVX1_LOC_147/A NAND2X1_LOC_640/a_36_24# 0.00fF
C16361 INVX1_LOC_448/A INVX1_LOC_119/Y 0.03fF
C16362 INVX1_LOC_379/A INVX1_LOC_226/Y 0.03fF
C16363 INVX1_LOC_49/Y INVX1_LOC_345/A 0.01fF
C16364 INVX1_LOC_211/Y INVX1_LOC_328/Y 0.67fF
C16365 INVX1_LOC_245/A INVX1_LOC_98/Y 0.03fF
C16366 INVX1_LOC_179/A INVX1_LOC_478/Y 0.01fF
C16367 INVX1_LOC_386/Y INVX1_LOC_405/Y 0.11fF
C16368 INVX1_LOC_11/Y INVX1_LOC_376/Y 0.07fF
C16369 NAND2X1_LOC_350/a_36_24# INVX1_LOC_79/A 0.01fF
C16370 INVX1_LOC_63/Y INVX1_LOC_50/Y 0.11fF
C16371 INVX1_LOC_576/Y INVX1_LOC_62/Y 0.11fF
C16372 NAND2X1_LOC_336/B INVX1_LOC_75/Y 0.11fF
C16373 INVX1_LOC_134/Y INVX1_LOC_652/Y 0.06fF
C16374 INVX1_LOC_145/Y INVX1_LOC_119/Y 0.04fF
C16375 INVX1_LOC_585/Y INVX1_LOC_223/Y 0.01fF
C16376 NAND2X1_LOC_24/Y NAND2X1_LOC_621/B 0.02fF
C16377 INVX1_LOC_208/A INVX1_LOC_44/Y 0.06fF
C16378 INVX1_LOC_614/A INVX1_LOC_645/Y 0.02fF
C16379 NAND2X1_LOC_689/B INVX1_LOC_338/Y 0.04fF
C16380 NAND2X1_LOC_513/A INVX1_LOC_588/A 0.75fF
C16381 INVX1_LOC_686/A INVX1_LOC_625/Y 0.08fF
C16382 NAND2X1_LOC_387/Y INVX1_LOC_179/A 0.07fF
C16383 INVX1_LOC_47/Y INVX1_LOC_141/Y 0.02fF
C16384 INVX1_LOC_382/A INVX1_LOC_339/Y 0.01fF
C16385 INVX1_LOC_444/Y NAND2X1_LOC_631/B 0.06fF
C16386 INVX1_LOC_221/Y INVX1_LOC_655/A 0.03fF
C16387 NAND2X1_LOC_557/B NAND2X1_LOC_490/a_36_24# 0.02fF
C16388 NAND2X1_LOC_196/a_36_24# INVX1_LOC_328/Y 0.00fF
C16389 INVX1_LOC_202/Y INVX1_LOC_203/A 0.04fF
C16390 INVX1_LOC_469/Y INVX1_LOC_26/Y 0.03fF
C16391 NAND2X1_LOC_274/B INVX1_LOC_32/Y 0.02fF
C16392 INVX1_LOC_386/Y INVX1_LOC_450/Y 0.01fF
C16393 INVX1_LOC_93/Y NAND2X1_LOC_489/A 0.05fF
C16394 INVX1_LOC_31/Y NAND2X1_LOC_545/A 0.15fF
C16395 INVX1_LOC_674/A INVX1_LOC_62/Y 0.07fF
C16396 NAND2X1_LOC_686/B INVX1_LOC_501/A 0.01fF
C16397 NAND2X1_LOC_181/A INVX1_LOC_26/Y 0.03fF
C16398 INVX1_LOC_360/A INVX1_LOC_347/A 0.07fF
C16399 INVX1_LOC_31/Y INVX1_LOC_653/Y 0.02fF
C16400 INVX1_LOC_387/Y NAND2X1_LOC_372/Y 0.01fF
C16401 NAND2X1_LOC_290/a_36_24# INVX1_LOC_79/A 0.00fF
C16402 INVX1_LOC_31/Y INVX1_LOC_666/Y 0.01fF
C16403 INVX1_LOC_129/A INVX1_LOC_92/A 0.01fF
C16404 NAND2X1_LOC_123/B INVX1_LOC_496/A 0.14fF
C16405 INVX1_LOC_601/Y INVX1_LOC_598/Y 0.27fF
C16406 INVX1_LOC_49/Y INVX1_LOC_280/A 0.13fF
C16407 INVX1_LOC_49/Y NAND2X1_LOC_372/Y 0.07fF
C16408 VDD NAND2X1_LOC_596/Y 0.01fF
C16409 INVX1_LOC_79/A INVX1_LOC_26/Y 4.91fF
C16410 INVX1_LOC_454/A INVX1_LOC_206/Y 0.05fF
C16411 VDD INVX1_LOC_228/Y 0.59fF
C16412 INVX1_LOC_301/A INVX1_LOC_400/Y 0.07fF
C16413 INVX1_LOC_133/Y NAND2X1_LOC_152/Y 0.79fF
C16414 INVX1_LOC_29/Y INVX1_LOC_41/A 0.01fF
C16415 INVX1_LOC_128/A INVX1_LOC_666/Y 0.01fF
C16416 VDD INVX1_LOC_383/A 0.00fF
C16417 INVX1_LOC_554/A INVX1_LOC_551/Y 0.02fF
C16418 VDD INVX1_LOC_510/Y 0.33fF
C16419 INVX1_LOC_629/Y INVX1_LOC_51/Y 0.04fF
C16420 INVX1_LOC_430/Y INVX1_LOC_443/A 0.03fF
C16421 INVX1_LOC_577/A INVX1_LOC_577/Y 0.04fF
C16422 INVX1_LOC_428/A INVX1_LOC_45/Y 0.07fF
C16423 INVX1_LOC_619/A INVX1_LOC_180/Y 0.03fF
C16424 INVX1_LOC_614/A VDD 0.01fF
C16425 INVX1_LOC_20/Y INVX1_LOC_584/A 0.03fF
C16426 VDD INVX1_LOC_42/A -0.00fF
C16427 INVX1_LOC_413/Y INVX1_LOC_586/A 0.15fF
C16428 NAND2X1_LOC_498/Y NAND2X1_LOC_332/B 0.07fF
C16429 INVX1_LOC_20/Y INVX1_LOC_400/Y 0.03fF
C16430 INVX1_LOC_31/A INVX1_LOC_33/Y 0.01fF
C16431 NAND2X1_LOC_750/Y INVX1_LOC_619/A 0.01fF
C16432 VDD INVX1_LOC_116/A 0.00fF
C16433 VDD INVX1_LOC_456/Y 0.21fF
C16434 INVX1_LOC_384/A INVX1_LOC_502/Y 0.02fF
C16435 VDD INVX1_LOC_684/A 0.00fF
C16436 VDD INVX1_LOC_158/Y 0.21fF
C16437 INVX1_LOC_446/A INVX1_LOC_50/Y 0.07fF
C16438 INVX1_LOC_395/A INVX1_LOC_97/Y 0.00fF
C16439 NAND2X1_LOC_721/a_36_24# INVX1_LOC_635/A 0.01fF
C16440 NAND2X1_LOC_475/A INVX1_LOC_145/Y 0.03fF
C16441 NAND2X1_LOC_13/Y NAND2X1_LOC_383/Y 0.12fF
C16442 VDD NAND2X1_LOC_843/A 0.05fF
C16443 INVX1_LOC_573/A NAND2X1_LOC_728/a_36_24# 0.00fF
C16444 INVX1_LOC_80/A NAND2X1_LOC_142/Y 0.01fF
C16445 INVX1_LOC_21/Y NAND2X1_LOC_513/Y 0.02fF
C16446 INVX1_LOC_11/Y INVX1_LOC_121/Y 0.38fF
C16447 VDD INVX1_LOC_103/Y 0.41fF
C16448 INVX1_LOC_400/Y INVX1_LOC_300/A 0.19fF
C16449 INVX1_LOC_402/A INVX1_LOC_51/Y 0.02fF
C16450 INVX1_LOC_206/Y INVX1_LOC_361/Y 0.14fF
C16451 INVX1_LOC_12/Y INVX1_LOC_482/A 0.03fF
C16452 INVX1_LOC_63/Y INVX1_LOC_275/A 0.03fF
C16453 INVX1_LOC_118/Y INVX1_LOC_118/A 0.00fF
C16454 NAND2X1_LOC_498/Y INVX1_LOC_503/Y 0.03fF
C16455 INVX1_LOC_448/A INVX1_LOC_502/Y 0.02fF
C16456 INVX1_LOC_288/Y INVX1_LOC_586/A 0.03fF
C16457 INVX1_LOC_11/Y INVX1_LOC_253/A 0.01fF
C16458 NAND2X1_LOC_475/A NAND2X1_LOC_133/a_36_24# 0.01fF
C16459 NAND2X1_LOC_317/A INVX1_LOC_46/Y 0.03fF
C16460 VDD INVX1_LOC_346/A 0.00fF
C16461 INVX1_LOC_391/Y INVX1_LOC_362/Y 0.00fF
C16462 INVX1_LOC_255/Y INVX1_LOC_48/Y 0.03fF
C16463 NAND2X1_LOC_152/B INVX1_LOC_53/Y 0.12fF
C16464 INVX1_LOC_197/A INVX1_LOC_134/Y 0.07fF
C16465 INVX1_LOC_522/Y NAND2X1_LOC_677/Y 0.03fF
C16466 INVX1_LOC_454/A NAND2X1_LOC_811/a_36_24# 0.01fF
C16467 INVX1_LOC_206/Y INVX1_LOC_261/Y 0.03fF
C16468 INVX1_LOC_20/Y INVX1_LOC_537/A 0.10fF
C16469 INVX1_LOC_58/Y NAND2X1_LOC_76/B 0.19fF
C16470 INVX1_LOC_425/A INVX1_LOC_304/A 0.04fF
C16471 INVX1_LOC_374/A INVX1_LOC_50/Y 0.49fF
C16472 INVX1_LOC_595/Y INVX1_LOC_366/A 0.01fF
C16473 INVX1_LOC_521/Y INVX1_LOC_46/Y 0.52fF
C16474 NAND2X1_LOC_24/Y INVX1_LOC_305/Y 0.10fF
C16475 INVX1_LOC_438/A INVX1_LOC_63/Y 0.07fF
C16476 INVX1_LOC_65/Y INVX1_LOC_117/Y 0.08fF
C16477 VDD INVX1_LOC_339/Y 0.21fF
C16478 NAND2X1_LOC_16/Y INVX1_LOC_31/Y 0.03fF
C16479 INVX1_LOC_35/Y INPUT_2 0.03fF
C16480 NAND2X1_LOC_669/Y INVX1_LOC_563/A 0.06fF
C16481 INVX1_LOC_391/A INVX1_LOC_547/Y 0.06fF
C16482 INVX1_LOC_395/A INVX1_LOC_94/Y 0.03fF
C16483 INVX1_LOC_361/Y INVX1_LOC_242/A 0.07fF
C16484 INVX1_LOC_375/A INVX1_LOC_624/Y 0.02fF
C16485 VDD NAND2X1_LOC_786/B 0.30fF
C16486 NAND2X1_LOC_69/B INVX1_LOC_41/Y 0.03fF
C16487 INVX1_LOC_191/Y INVX1_LOC_26/Y 0.09fF
C16488 INVX1_LOC_11/Y INVX1_LOC_295/A 0.18fF
C16489 INPUT_7 INVX1_LOC_40/Y 0.44fF
C16490 NAND2X1_LOC_385/a_36_24# INVX1_LOC_100/Y 0.00fF
C16491 INVX1_LOC_84/A INPUT_1 0.01fF
C16492 INVX1_LOC_361/Y INVX1_LOC_686/A 0.07fF
C16493 NAND2X1_LOC_332/B INVX1_LOC_47/Y 0.07fF
C16494 INVX1_LOC_20/Y INVX1_LOC_496/Y 0.03fF
C16495 INVX1_LOC_554/A NAND2X1_LOC_410/Y 0.00fF
C16496 INVX1_LOC_560/A NAND2X1_LOC_558/B 0.21fF
C16497 INVX1_LOC_577/A INVX1_LOC_26/Y 0.00fF
C16498 INVX1_LOC_25/Y INVX1_LOC_145/Y 0.03fF
C16499 INVX1_LOC_137/A INVX1_LOC_507/Y 0.00fF
C16500 INVX1_LOC_228/Y NAND2X1_LOC_786/B 0.02fF
C16501 NAND2X1_LOC_158/a_36_24# INVX1_LOC_186/A 0.00fF
C16502 INVX1_LOC_474/Y INVX1_LOC_48/Y 0.10fF
C16503 NAND2X1_LOC_180/B INVX1_LOC_69/Y 0.03fF
C16504 NAND2X1_LOC_754/a_36_24# INVX1_LOC_211/A 0.00fF
C16505 VDD INVX1_LOC_635/Y 0.64fF
C16506 INVX1_LOC_530/Y INVX1_LOC_328/Y 0.05fF
C16507 NAND2X1_LOC_768/B INVX1_LOC_45/Y 0.01fF
C16508 NAND2X1_LOC_498/Y INVX1_LOC_242/Y 0.03fF
C16509 INVX1_LOC_294/A INVX1_LOC_281/Y 0.00fF
C16510 INVX1_LOC_435/A INVX1_LOC_230/A 0.14fF
C16511 INVX1_LOC_560/A INVX1_LOC_79/A 0.01fF
C16512 NAND2X1_LOC_532/Y INVX1_LOC_401/A 0.18fF
C16513 INPUT_3 NAND2X1_LOC_531/Y 0.05fF
C16514 NAND2X1_LOC_638/A INVX1_LOC_298/A 0.11fF
C16515 INVX1_LOC_261/Y INVX1_LOC_686/A 0.02fF
C16516 INVX1_LOC_437/A INVX1_LOC_453/Y 0.08fF
C16517 NAND2X1_LOC_638/A INVX1_LOC_498/A 0.01fF
C16518 INVX1_LOC_564/Y INVX1_LOC_79/A 0.00fF
C16519 INVX1_LOC_258/Y INVX1_LOC_686/A 0.07fF
C16520 INVX1_LOC_442/Y NAND2X1_LOC_527/Y 0.00fF
C16521 INVX1_LOC_180/A INVX1_LOC_26/Y 0.01fF
C16522 INVX1_LOC_481/Y INVX1_LOC_48/Y 0.01fF
C16523 NAND2X1_LOC_142/Y INVX1_LOC_102/Y 0.01fF
C16524 INVX1_LOC_510/A INVX1_LOC_665/Y 0.01fF
C16525 INVX1_LOC_54/Y NAND2X1_LOC_775/B 0.02fF
C16526 INVX1_LOC_550/Y INVX1_LOC_186/Y 0.04fF
C16527 INVX1_LOC_449/A INVX1_LOC_49/Y 0.03fF
C16528 NAND2X1_LOC_332/B INVX1_LOC_119/Y 0.10fF
C16529 INVX1_LOC_89/Y NAND2X1_LOC_448/A 0.18fF
C16530 INVX1_LOC_195/Y NAND2X1_LOC_222/a_36_24# 0.00fF
C16531 INVX1_LOC_603/Y INVX1_LOC_69/Y 0.37fF
C16532 INVX1_LOC_32/Y INVX1_LOC_159/Y 0.07fF
C16533 INVX1_LOC_358/A INVX1_LOC_356/Y 0.01fF
C16534 INVX1_LOC_340/Y INVX1_LOC_41/Y 0.03fF
C16535 INVX1_LOC_596/A INVX1_LOC_245/A 0.00fF
C16536 INVX1_LOC_54/Y NAND2X1_LOC_706/B 0.10fF
C16537 INVX1_LOC_550/A INVX1_LOC_186/Y 0.01fF
C16538 INVX1_LOC_266/A NAND2X1_LOC_545/A 0.05fF
C16539 INVX1_LOC_51/Y INVX1_LOC_653/Y 0.46fF
C16540 INVX1_LOC_347/Y INVX1_LOC_115/A 0.48fF
C16541 INVX1_LOC_595/Y INVX1_LOC_6/Y 0.04fF
C16542 INVX1_LOC_76/Y INVX1_LOC_203/A 0.01fF
C16543 INVX1_LOC_602/Y INVX1_LOC_674/Y 0.02fF
C16544 INVX1_LOC_53/A NAND2X1_LOC_836/B 0.07fF
C16545 INVX1_LOC_625/A INVX1_LOC_58/Y 1.27fF
C16546 INVX1_LOC_257/A NAND2X1_LOC_775/B 0.20fF
C16547 INVX1_LOC_69/Y INVX1_LOC_478/Y 0.09fF
C16548 INVX1_LOC_293/Y INVX1_LOC_369/Y 0.01fF
C16549 INVX1_LOC_89/Y INVX1_LOC_295/Y 0.01fF
C16550 INVX1_LOC_504/A NAND2X1_LOC_440/A 0.03fF
C16551 INVX1_LOC_502/A INVX1_LOC_519/A 0.03fF
C16552 INVX1_LOC_31/Y INVX1_LOC_18/Y 0.00fF
C16553 INVX1_LOC_45/Y NAND2X1_LOC_832/A 0.83fF
C16554 INVX1_LOC_41/Y NAND2X1_LOC_541/B 0.22fF
C16555 INVX1_LOC_45/Y INVX1_LOC_443/A 0.03fF
C16556 INVX1_LOC_91/Y INVX1_LOC_94/A 0.03fF
C16557 INVX1_LOC_504/A INVX1_LOC_245/A 0.03fF
C16558 GATE_662 INVX1_LOC_46/Y 0.01fF
C16559 INVX1_LOC_266/A INVX1_LOC_666/Y 0.07fF
C16560 NAND2X1_LOC_387/Y INVX1_LOC_69/Y 0.25fF
C16561 INVX1_LOC_99/Y INVX1_LOC_242/Y 0.13fF
C16562 INVX1_LOC_405/Y INVX1_LOC_7/Y 0.05fF
C16563 INVX1_LOC_211/Y INVX1_LOC_224/A 0.06fF
C16564 INVX1_LOC_41/Y INVX1_LOC_383/Y 0.05fF
C16565 INVX1_LOC_254/Y INVX1_LOC_9/Y 0.07fF
C16566 NAND2X1_LOC_612/A INVX1_LOC_475/Y 0.19fF
C16567 INVX1_LOC_99/Y INVX1_LOC_487/A 0.01fF
C16568 INVX1_LOC_657/A INVX1_LOC_656/Y 0.15fF
C16569 INVX1_LOC_79/A NAND2X1_LOC_211/a_36_24# 0.00fF
C16570 INVX1_LOC_556/Y INVX1_LOC_100/Y 0.03fF
C16571 INVX1_LOC_567/Y INVX1_LOC_135/Y 0.01fF
C16572 INVX1_LOC_615/A INVX1_LOC_615/Y 0.02fF
C16573 NAND2X1_LOC_388/A INVX1_LOC_63/Y 0.03fF
C16574 INVX1_LOC_26/Y INVX1_LOC_48/Y 0.22fF
C16575 INVX1_LOC_261/Y NAND2X1_LOC_334/A 0.03fF
C16576 INVX1_LOC_376/Y INVX1_LOC_374/Y 0.02fF
C16577 NAND2X1_LOC_782/A INVX1_LOC_612/A 0.09fF
C16578 INVX1_LOC_469/Y NAND2X1_LOC_605/B 0.24fF
C16579 INVX1_LOC_79/A INVX1_LOC_603/A 0.01fF
C16580 INVX1_LOC_183/A INVX1_LOC_6/Y 0.07fF
C16581 INVX1_LOC_58/Y NAND2X1_LOC_52/Y 0.07fF
C16582 INVX1_LOC_350/A INVX1_LOC_347/A 0.13fF
C16583 NAND2X1_LOC_364/a_36_24# INVX1_LOC_90/Y 0.00fF
C16584 INVX1_LOC_254/Y INVX1_LOC_62/Y 0.03fF
C16585 INVX1_LOC_389/Y INVX1_LOC_6/Y 0.02fF
C16586 INVX1_LOC_581/A INVX1_LOC_611/A 0.01fF
C16587 INVX1_LOC_49/Y INVX1_LOC_328/Y 0.07fF
C16588 INVX1_LOC_47/Y INVX1_LOC_242/Y 0.04fF
C16589 NAND2X1_LOC_753/Y INVX1_LOC_90/Y 0.09fF
C16590 INVX1_LOC_514/A INVX1_LOC_479/A 0.00fF
C16591 INVX1_LOC_49/Y INVX1_LOC_518/A 0.03fF
C16592 INVX1_LOC_223/Y INVX1_LOC_44/Y 0.09fF
C16593 NAND2X1_LOC_334/A NAND2X1_LOC_431/a_36_24# 0.01fF
C16594 NAND2X1_LOC_673/B INVX1_LOC_223/A 0.02fF
C16595 INVX1_LOC_565/A INVX1_LOC_636/A 0.05fF
C16596 INVX1_LOC_117/Y INVX1_LOC_588/A 0.14fF
C16597 INVX1_LOC_539/Y INVX1_LOC_479/A 0.01fF
C16598 INVX1_LOC_506/A INVX1_LOC_74/Y 0.02fF
C16599 INVX1_LOC_412/Y INVX1_LOC_638/A 0.44fF
C16600 INVX1_LOC_395/A INVX1_LOC_615/A 0.85fF
C16601 NAND2X1_LOC_750/Y NAND2X1_LOC_61/A 0.01fF
C16602 NAND2X1_LOC_228/a_36_24# INVX1_LOC_206/Y 0.00fF
C16603 INVX1_LOC_257/Y NAND2X1_LOC_543/B 0.00fF
C16604 NAND2X1_LOC_814/a_36_24# INVX1_LOC_655/A 0.01fF
C16605 INVX1_LOC_6/Y INVX1_LOC_109/A 0.03fF
C16606 INVX1_LOC_193/A INVX1_LOC_92/A 0.00fF
C16607 INVX1_LOC_62/A INVX1_LOC_92/A 0.08fF
C16608 INVX1_LOC_26/Y INVX1_LOC_472/Y 0.07fF
C16609 NAND2X1_LOC_847/A NAND2X1_LOC_287/a_36_24# 0.00fF
C16610 INVX1_LOC_400/Y NAND2X1_LOC_373/Y 0.03fF
C16611 INVX1_LOC_554/A INVX1_LOC_558/A 0.04fF
C16612 INVX1_LOC_534/Y INVX1_LOC_479/A 0.04fF
C16613 NAND2X1_LOC_66/Y INVX1_LOC_487/A 0.02fF
C16614 INVX1_LOC_479/A INVX1_LOC_9/Y 0.11fF
C16615 INVX1_LOC_438/Y INVX1_LOC_278/A 0.03fF
C16616 INVX1_LOC_207/Y INVX1_LOC_210/A 0.00fF
C16617 INVX1_LOC_265/Y NAND2X1_LOC_331/B 0.19fF
C16618 INVX1_LOC_279/A INVX1_LOC_384/Y 0.09fF
C16619 NAND2X1_LOC_471/a_36_24# INVX1_LOC_109/Y 0.01fF
C16620 INVX1_LOC_166/Y INVX1_LOC_479/A 0.02fF
C16621 INPUT_6 INVX1_LOC_5/Y 0.01fF
C16622 NAND2X1_LOC_528/Y INVX1_LOC_62/Y 0.11fF
C16623 INVX1_LOC_578/A INVX1_LOC_412/A 0.53fF
C16624 INVX1_LOC_420/Y INVX1_LOC_45/Y 0.00fF
C16625 NAND2X1_LOC_416/B INVX1_LOC_245/A 0.22fF
C16626 INVX1_LOC_62/Y INVX1_LOC_479/A 0.39fF
C16627 INVX1_LOC_68/Y INPUT_0 0.00fF
C16628 INVX1_LOC_446/Y NAND2X1_LOC_520/B 0.03fF
C16629 NAND2X1_LOC_714/a_36_24# INVX1_LOC_375/A 0.00fF
C16630 INVX1_LOC_490/Y INVX1_LOC_51/Y 0.00fF
C16631 NAND2X1_LOC_780/B INVX1_LOC_522/Y 0.03fF
C16632 INVX1_LOC_21/Y NAND2X1_LOC_69/B 0.04fF
C16633 NAND2X1_LOC_16/Y INVX1_LOC_51/Y 0.03fF
C16634 NAND2X1_LOC_7/Y INVX1_LOC_99/Y 0.08fF
C16635 INVX1_LOC_381/A INVX1_LOC_49/A 0.03fF
C16636 INVX1_LOC_409/Y NAND2X1_LOC_123/A 0.01fF
C16637 INVX1_LOC_46/Y INVX1_LOC_109/Y 0.03fF
C16638 NAND2X1_LOC_502/a_36_24# INVX1_LOC_274/A 0.00fF
C16639 NAND2X1_LOC_13/Y INVX1_LOC_320/Y 0.01fF
C16640 INVX1_LOC_224/Y NAND2X1_LOC_336/B 0.10fF
C16641 INVX1_LOC_20/Y NAND2X1_LOC_498/Y 0.07fF
C16642 INVX1_LOC_505/Y INVX1_LOC_462/Y 0.07fF
C16643 INVX1_LOC_301/A INVX1_LOC_99/Y 0.01fF
C16644 INVX1_LOC_627/A INVX1_LOC_54/Y 0.01fF
C16645 INVX1_LOC_133/Y INVX1_LOC_54/Y 0.00fF
C16646 INVX1_LOC_206/Y INVX1_LOC_307/A 0.20fF
C16647 NAND2X1_LOC_318/A INVX1_LOC_266/Y 0.07fF
C16648 NAND2X1_LOC_180/B INVX1_LOC_586/A 0.03fF
C16649 INVX1_LOC_428/A INVX1_LOC_293/Y 0.03fF
C16650 INVX1_LOC_137/A INVX1_LOC_522/Y 0.02fF
C16651 INVX1_LOC_353/Y INVX1_LOC_51/Y 0.03fF
C16652 NAND2X1_LOC_336/B INVX1_LOC_578/A 0.01fF
C16653 INVX1_LOC_257/Y INVX1_LOC_469/A 0.04fF
C16654 VDD INVX1_LOC_360/Y 0.26fF
C16655 INPUT_0 INVX1_LOC_600/A 0.08fF
C16656 INPUT_0 NAND2X1_LOC_130/Y 0.03fF
C16657 INVX1_LOC_558/A INVX1_LOC_126/Y 0.01fF
C16658 INVX1_LOC_400/Y INVX1_LOC_375/Y 0.17fF
C16659 INVX1_LOC_617/A INVX1_LOC_384/A 0.04fF
C16660 INPUT_0 INVX1_LOC_64/A 0.00fF
C16661 INVX1_LOC_417/Y INVX1_LOC_560/A 0.02fF
C16662 NAND2X1_LOC_685/A INVX1_LOC_586/A 0.10fF
C16663 INVX1_LOC_438/Y INVX1_LOC_453/Y 1.42fF
C16664 INVX1_LOC_554/A INVX1_LOC_46/Y 0.02fF
C16665 VDD INVX1_LOC_105/A 0.15fF
C16666 INVX1_LOC_192/Y INVX1_LOC_194/A 0.00fF
C16667 INVX1_LOC_54/Y NAND2X1_LOC_184/a_36_24# 0.04fF
C16668 NAND2X1_LOC_457/A INVX1_LOC_159/A 0.02fF
C16669 NAND2X1_LOC_685/B INVX1_LOC_536/A 0.12fF
C16670 INVX1_LOC_54/Y INVX1_LOC_307/Y 0.01fF
C16671 INVX1_LOC_160/Y INVX1_LOC_155/Y 0.01fF
C16672 INVX1_LOC_533/Y INVX1_LOC_99/Y 0.00fF
C16673 INVX1_LOC_335/Y INVX1_LOC_340/Y 0.03fF
C16674 INVX1_LOC_564/Y INVX1_LOC_59/Y 0.01fF
C16675 INVX1_LOC_68/Y NAND2X1_LOC_123/A 0.44fF
C16676 INVX1_LOC_586/A NAND2X1_LOC_411/Y 0.01fF
C16677 INVX1_LOC_328/Y INVX1_LOC_297/Y 0.01fF
C16678 NAND2X1_LOC_520/B INVX1_LOC_145/Y 0.15fF
C16679 INVX1_LOC_551/Y INVX1_LOC_53/Y 0.07fF
C16680 INVX1_LOC_468/Y INVX1_LOC_618/Y 0.01fF
C16681 INVX1_LOC_45/Y NAND2X1_LOC_270/a_36_24# 0.00fF
C16682 INVX1_LOC_6/Y NAND2X1_LOC_772/a_36_24# 0.00fF
C16683 INVX1_LOC_560/A INVX1_LOC_48/Y 0.07fF
C16684 INVX1_LOC_76/A INVX1_LOC_92/A 0.03fF
C16685 INVX1_LOC_374/A NAND2X1_LOC_648/a_36_24# 0.00fF
C16686 INVX1_LOC_65/Y INVX1_LOC_178/A 0.00fF
C16687 NAND2X1_LOC_25/a_36_24# INVX1_LOC_6/A 0.00fF
C16688 INVX1_LOC_617/A INVX1_LOC_448/A 0.31fF
C16689 INVX1_LOC_564/Y INVX1_LOC_48/Y 0.03fF
C16690 NAND2X1_LOC_520/a_36_24# INVX1_LOC_45/Y 0.00fF
C16691 INVX1_LOC_202/Y INVX1_LOC_266/Y 0.03fF
C16692 INVX1_LOC_20/Y INVX1_LOC_99/Y 0.21fF
C16693 INPUT_0 INVX1_LOC_484/A 0.00fF
C16694 INVX1_LOC_200/Y INVX1_LOC_6/Y 0.01fF
C16695 INVX1_LOC_54/Y NAND2X1_LOC_831/a_36_24# 0.01fF
C16696 INVX1_LOC_586/A INVX1_LOC_637/A 0.01fF
C16697 NAND2X1_LOC_393/a_36_24# INVX1_LOC_63/Y 0.00fF
C16698 INVX1_LOC_290/Y INVX1_LOC_261/Y 3.93fF
C16699 NAND2X1_LOC_333/B INVX1_LOC_94/A 0.02fF
C16700 INVX1_LOC_442/Y INVX1_LOC_686/A 0.17fF
C16701 NAND2X1_LOC_164/Y INVX1_LOC_58/Y 0.06fF
C16702 NAND2X1_LOC_387/Y INVX1_LOC_586/A 0.04fF
C16703 INVX1_LOC_245/A NAND2X1_LOC_76/B 0.04fF
C16704 INVX1_LOC_76/Y INVX1_LOC_186/Y 0.02fF
C16705 NAND2X1_LOC_179/Y INVX1_LOC_134/Y 0.06fF
C16706 INVX1_LOC_40/Y INVX1_LOC_55/Y 0.22fF
C16707 INVX1_LOC_540/Y INVX1_LOC_501/A 0.01fF
C16708 NAND2X1_LOC_472/a_36_24# INVX1_LOC_50/Y 0.00fF
C16709 INVX1_LOC_271/A INVX1_LOC_154/A 0.10fF
C16710 INVX1_LOC_17/Y INVX1_LOC_519/A 0.02fF
C16711 INVX1_LOC_617/Y INVX1_LOC_665/Y 0.02fF
C16712 INVX1_LOC_275/Y INVX1_LOC_284/A 0.02fF
C16713 VDD INVX1_LOC_430/Y 0.38fF
C16714 INVX1_LOC_137/A INVX1_LOC_508/A 0.02fF
C16715 INVX1_LOC_558/A INVX1_LOC_199/Y 0.12fF
C16716 INVX1_LOC_165/Y INVX1_LOC_49/Y 0.01fF
C16717 INVX1_LOC_84/A INVX1_LOC_50/Y 0.03fF
C16718 INVX1_LOC_172/Y INVX1_LOC_32/Y 0.04fF
C16719 INVX1_LOC_602/A INVX1_LOC_623/Y 0.00fF
C16720 INVX1_LOC_65/Y INVX1_LOC_58/Y 0.03fF
C16721 INVX1_LOC_400/A NAND2X1_LOC_237/Y 0.01fF
C16722 INVX1_LOC_20/Y INVX1_LOC_123/A 0.06fF
C16723 INPUT_3 INVX1_LOC_382/A 0.00fF
C16724 INVX1_LOC_300/A INVX1_LOC_99/Y 0.22fF
C16725 INVX1_LOC_369/A INVX1_LOC_48/Y 0.03fF
C16726 INVX1_LOC_259/A INVX1_LOC_501/A 0.04fF
C16727 INVX1_LOC_561/Y INVX1_LOC_26/Y 0.04fF
C16728 INVX1_LOC_99/Y INVX1_LOC_197/Y 0.03fF
C16729 INVX1_LOC_54/Y INVX1_LOC_633/Y 0.06fF
C16730 INVX1_LOC_54/Y INVX1_LOC_581/A 0.03fF
C16731 INVX1_LOC_418/Y INVX1_LOC_130/Y 0.03fF
C16732 INVX1_LOC_20/Y INVX1_LOC_47/Y 0.47fF
C16733 INVX1_LOC_435/A INVX1_LOC_681/A 0.01fF
C16734 INVX1_LOC_130/Y INVX1_LOC_159/Y 0.02fF
C16735 INVX1_LOC_133/A INVX1_LOC_132/A 0.01fF
C16736 INVX1_LOC_93/Y INVX1_LOC_635/A 0.08fF
C16737 INVX1_LOC_619/A NAND2X1_LOC_243/A 0.09fF
C16738 INVX1_LOC_555/A INVX1_LOC_508/Y -0.01fF
C16739 INVX1_LOC_76/Y INVX1_LOC_347/Y 0.14fF
C16740 INVX1_LOC_270/A INVX1_LOC_199/Y 0.04fF
C16741 INVX1_LOC_570/A INVX1_LOC_655/A 0.07fF
C16742 INVX1_LOC_581/A INVX1_LOC_611/Y 0.02fF
C16743 INVX1_LOC_11/Y INVX1_LOC_251/A 0.08fF
C16744 INVX1_LOC_501/Y INVX1_LOC_58/Y 0.01fF
C16745 INVX1_LOC_361/Y NAND2X1_LOC_478/a_36_24# 0.00fF
C16746 NAND2X1_LOC_267/A INVX1_LOC_155/Y 0.03fF
C16747 INVX1_LOC_586/A INVX1_LOC_491/A 0.00fF
C16748 INVX1_LOC_50/Y NAND2X1_LOC_67/Y 0.02fF
C16749 INVX1_LOC_76/Y INVX1_LOC_328/Y 0.04fF
C16750 INVX1_LOC_576/A INVX1_LOC_47/Y 0.00fF
C16751 NAND2X1_LOC_275/Y INVX1_LOC_48/Y 0.07fF
C16752 INVX1_LOC_32/Y NAND2X1_LOC_595/Y 0.61fF
C16753 INVX1_LOC_174/A INVX1_LOC_6/Y 0.09fF
C16754 INVX1_LOC_602/A INVX1_LOC_63/Y 0.12fF
C16755 INVX1_LOC_452/A INVX1_LOC_671/A 0.53fF
C16756 INVX1_LOC_300/A INVX1_LOC_123/A 0.03fF
C16757 NAND2X1_LOC_726/a_36_24# INVX1_LOC_662/A 0.00fF
C16758 INVX1_LOC_53/Y NAND2X1_LOC_759/Y 0.02fF
C16759 INVX1_LOC_48/Y INVX1_LOC_603/A 0.01fF
C16760 NAND2X1_LOC_147/B NAND2X1_LOC_342/A 0.02fF
C16761 INVX1_LOC_117/Y NAND2X1_LOC_646/A 0.06fF
C16762 INVX1_LOC_45/Y NAND2X1_LOC_488/Y 0.06fF
C16763 INVX1_LOC_300/A INVX1_LOC_47/Y 0.03fF
C16764 NAND2X1_LOC_152/B INVX1_LOC_662/A 0.07fF
C16765 NAND2X1_LOC_142/Y NAND2X1_LOC_843/B 0.02fF
C16766 INVX1_LOC_20/Y INVX1_LOC_119/Y 0.04fF
C16767 INVX1_LOC_197/A NAND2X1_LOC_221/a_36_24# 0.02fF
C16768 INVX1_LOC_40/Y INVX1_LOC_18/Y 0.22fF
C16769 INVX1_LOC_117/Y INVX1_LOC_623/Y 0.00fF
C16770 INVX1_LOC_69/Y INVX1_LOC_504/Y 0.08fF
C16771 INVX1_LOC_235/Y INVX1_LOC_79/A 0.19fF
C16772 INVX1_LOC_185/Y INVX1_LOC_645/Y 0.13fF
C16773 INVX1_LOC_49/Y INVX1_LOC_352/A 0.01fF
C16774 NAND2X1_LOC_722/a_36_24# INVX1_LOC_41/Y 0.01fF
C16775 NAND2X1_LOC_775/B INVX1_LOC_89/Y 0.10fF
C16776 INVX1_LOC_586/A INVX1_LOC_91/A 0.03fF
C16777 INVX1_LOC_12/Y INVX1_LOC_9/Y 0.16fF
C16778 INVX1_LOC_17/Y INVX1_LOC_659/A 0.01fF
C16779 INVX1_LOC_671/A NAND2X1_LOC_850/a_36_24# 0.01fF
C16780 INVX1_LOC_469/Y INVX1_LOC_506/A 0.00fF
C16781 NAND2X1_LOC_837/B NAND2X1_LOC_827/Y 0.06fF
C16782 INVX1_LOC_625/A NAND2X1_LOC_91/a_36_24# 0.00fF
C16783 INVX1_LOC_68/Y INVX1_LOC_211/A 0.15fF
C16784 NAND2X1_LOC_531/Y NAND2X1_LOC_4/a_36_24# 0.00fF
C16785 INVX1_LOC_619/A NAND2X1_LOC_786/B 0.01fF
C16786 INVX1_LOC_169/A INVX1_LOC_388/A 0.02fF
C16787 NAND2X1_LOC_532/Y INPUT_1 0.03fF
C16788 INVX1_LOC_547/A INVX1_LOC_479/A 0.01fF
C16789 INVX1_LOC_80/A INVX1_LOC_652/A 0.01fF
C16790 INVX1_LOC_68/Y INVX1_LOC_64/Y 0.27fF
C16791 NAND2X1_LOC_260/Y INVX1_LOC_663/A 0.01fF
C16792 INVX1_LOC_31/Y INVX1_LOC_100/A 0.21fF
C16793 INVX1_LOC_58/Y INVX1_LOC_479/Y 0.01fF
C16794 INVX1_LOC_390/A INVX1_LOC_230/A 0.04fF
C16795 INVX1_LOC_625/A INVX1_LOC_245/A 0.02fF
C16796 NAND2X1_LOC_13/Y INVX1_LOC_666/Y 0.16fF
C16797 INVX1_LOC_361/Y NAND2X1_LOC_542/A 0.07fF
C16798 INVX1_LOC_6/Y NAND2X1_LOC_819/a_36_24# 0.00fF
C16799 NAND2X1_LOC_755/B INVX1_LOC_272/A 0.02fF
C16800 INVX1_LOC_100/A NAND2X1_LOC_104/a_36_24# 0.01fF
C16801 INVX1_LOC_496/A INVX1_LOC_50/Y 0.08fF
C16802 NAND2X1_LOC_813/a_36_24# INVX1_LOC_178/A 0.01fF
C16803 INVX1_LOC_199/Y INVX1_LOC_46/Y 0.37fF
C16804 INVX1_LOC_555/A INVX1_LOC_633/A 0.05fF
C16805 INVX1_LOC_11/Y NAND2X1_LOC_258/a_36_24# 0.00fF
C16806 INVX1_LOC_117/Y INVX1_LOC_63/Y 0.80fF
C16807 INVX1_LOC_318/A INVX1_LOC_58/Y 0.00fF
C16808 INVX1_LOC_53/Y NAND2X1_LOC_410/Y 0.02fF
C16809 INVX1_LOC_116/Y INVX1_LOC_114/A 0.00fF
C16810 INVX1_LOC_294/A INVX1_LOC_245/A 0.01fF
C16811 INVX1_LOC_12/Y INVX1_LOC_62/Y 0.10fF
C16812 INVX1_LOC_361/Y INVX1_LOC_376/Y 0.07fF
C16813 INVX1_LOC_11/Y INVX1_LOC_652/A 0.04fF
C16814 INVX1_LOC_638/Y INVX1_LOC_641/A 0.01fF
C16815 INVX1_LOC_504/A NAND2X1_LOC_597/Y 0.09fF
C16816 INVX1_LOC_211/A INVX1_LOC_600/A 0.13fF
C16817 NAND2X1_LOC_184/Y NAND2X1_LOC_274/B 0.46fF
C16818 INVX1_LOC_48/Y NAND2X1_LOC_626/Y 0.01fF
C16819 INVX1_LOC_178/Y INVX1_LOC_87/Y 0.46fF
C16820 INVX1_LOC_11/Y INVX1_LOC_11/A 0.01fF
C16821 INVX1_LOC_315/A INVX1_LOC_41/Y 0.05fF
C16822 NAND2X1_LOC_775/B NAND2X1_LOC_544/B 0.02fF
C16823 INVX1_LOC_176/A NAND2X1_LOC_626/a_36_24# 0.00fF
C16824 INVX1_LOC_32/Y NAND2X1_LOC_372/Y 0.03fF
C16825 VDD NAND2X1_LOC_61/A -0.00fF
C16826 INVX1_LOC_391/A INVX1_LOC_62/Y 0.01fF
C16827 NAND2X1_LOC_686/A INVX1_LOC_245/A 0.08fF
C16828 NAND2X1_LOC_521/Y NAND2X1_LOC_844/A 0.04fF
C16829 INVX1_LOC_257/Y INVX1_LOC_409/Y 0.03fF
C16830 INVX1_LOC_74/Y NAND2X1_LOC_586/Y 0.01fF
C16831 INVX1_LOC_65/A INVX1_LOC_66/Y 0.00fF
C16832 NAND2X1_LOC_61/A INVX1_LOC_228/Y 0.04fF
C16833 INVX1_LOC_652/Y INVX1_LOC_338/Y 0.02fF
C16834 INVX1_LOC_199/Y INVX1_LOC_75/A 0.04fF
C16835 INVX1_LOC_58/Y INVX1_LOC_588/A 0.04fF
C16836 INVX1_LOC_399/Y INVX1_LOC_531/Y 0.04fF
C16837 NAND2X1_LOC_503/B INVX1_LOC_273/A 0.08fF
C16838 VDD NAND2X1_LOC_506/B 0.11fF
C16839 NAND2X1_LOC_627/Y INVX1_LOC_487/A 0.00fF
C16840 INVX1_LOC_206/Y INVX1_LOC_412/A 0.03fF
C16841 VDD INVX1_LOC_185/Y 0.26fF
C16842 NAND2X1_LOC_274/B INVX1_LOC_75/Y 0.01fF
C16843 INVX1_LOC_203/Y INVX1_LOC_271/A 0.00fF
C16844 VDD INVX1_LOC_45/Y 1.85fF
C16845 NAND2X1_LOC_585/a_36_24# NAND2X1_LOC_122/Y 0.00fF
C16846 INVX1_LOC_133/Y INVX1_LOC_649/Y 0.01fF
C16847 INVX1_LOC_162/Y INVX1_LOC_549/A 0.07fF
C16848 INVX1_LOC_627/A NAND2X1_LOC_677/Y 0.01fF
C16849 INVX1_LOC_206/Y NAND2X1_LOC_707/A 0.01fF
C16850 INVX1_LOC_228/Y INVX1_LOC_45/Y 0.02fF
C16851 INVX1_LOC_133/Y NAND2X1_LOC_677/Y 1.03fF
C16852 INVX1_LOC_151/Y NAND2X1_LOC_685/A 0.02fF
C16853 VDD INPUT_3 0.87fF
C16854 INVX1_LOC_20/Y NAND2X1_LOC_475/A 0.09fF
C16855 INVX1_LOC_289/A NAND2X1_LOC_801/A 0.15fF
C16856 INVX1_LOC_165/Y NAND2X1_LOC_498/B 0.01fF
C16857 INVX1_LOC_249/Y NAND2X1_LOC_122/Y 0.01fF
C16858 INVX1_LOC_521/Y INVX1_LOC_76/Y 0.01fF
C16859 INVX1_LOC_165/Y INVX1_LOC_76/Y 0.01fF
C16860 NAND2X1_LOC_781/B INVX1_LOC_145/Y 0.03fF
C16861 NAND2X1_LOC_790/B INVX1_LOC_59/Y 0.27fF
C16862 INVX1_LOC_206/Y NAND2X1_LOC_336/B 0.02fF
C16863 VDD NAND2X1_LOC_331/Y 0.13fF
C16864 INVX1_LOC_412/Y INVX1_LOC_134/Y 0.01fF
C16865 NAND2X1_LOC_101/a_36_24# INVX1_LOC_586/A 0.00fF
C16866 INVX1_LOC_412/A INVX1_LOC_686/A 0.04fF
C16867 VDD NAND2X1_LOC_376/Y 0.00fF
C16868 INVX1_LOC_266/Y INVX1_LOC_76/Y 0.07fF
C16869 VDD NAND2X1_LOC_69/Y 0.01fF
C16870 NAND2X1_LOC_790/B INVX1_LOC_48/Y 0.44fF
C16871 INVX1_LOC_317/Y NAND2X1_LOC_176/a_36_24# 0.00fF
C16872 INVX1_LOC_224/Y NAND2X1_LOC_169/A 0.01fF
C16873 INVX1_LOC_49/Y INVX1_LOC_109/Y 0.07fF
C16874 NAND2X1_LOC_475/A INVX1_LOC_300/A 0.04fF
C16875 INVX1_LOC_446/A INVX1_LOC_117/Y 0.46fF
C16876 INVX1_LOC_140/Y INVX1_LOC_188/Y 0.03fF
C16877 NAND2X1_LOC_498/Y INVX1_LOC_375/Y 0.16fF
C16878 INVX1_LOC_395/A NAND2X1_LOC_237/Y 0.05fF
C16879 NAND2X1_LOC_475/A INVX1_LOC_197/Y 0.03fF
C16880 INVX1_LOC_459/A INVX1_LOC_31/Y 0.02fF
C16881 INVX1_LOC_614/A INVX1_LOC_185/Y 0.03fF
C16882 INVX1_LOC_418/A INVX1_LOC_53/Y 0.30fF
C16883 INVX1_LOC_191/Y INVX1_LOC_81/Y 0.00fF
C16884 INVX1_LOC_311/Y INVX1_LOC_366/A 0.01fF
C16885 NAND2X1_LOC_457/A INVX1_LOC_116/Y 0.04fF
C16886 INVX1_LOC_558/A INVX1_LOC_53/Y 0.21fF
C16887 INVX1_LOC_17/Y INVX1_LOC_445/A 0.06fF
C16888 INVX1_LOC_429/A INVX1_LOC_453/Y 0.03fF
C16889 INVX1_LOC_95/Y INVX1_LOC_49/Y 0.15fF
C16890 INVX1_LOC_395/A INVX1_LOC_230/A 0.00fF
C16891 INVX1_LOC_602/A INVX1_LOC_20/A 0.04fF
C16892 INVX1_LOC_557/A NAND2X1_LOC_317/a_36_24# 0.01fF
C16893 INVX1_LOC_121/Y INVX1_LOC_361/Y 0.13fF
C16894 INVX1_LOC_457/Y INVX1_LOC_588/Y 0.35fF
C16895 INVX1_LOC_410/Y INVX1_LOC_665/Y 0.01fF
C16896 INVX1_LOC_103/A INVX1_LOC_48/Y 0.01fF
C16897 INVX1_LOC_617/Y INVX1_LOC_134/Y 0.68fF
C16898 INVX1_LOC_119/A INVX1_LOC_134/Y 0.01fF
C16899 INVX1_LOC_43/Y INVX1_LOC_366/A 0.01fF
C16900 INVX1_LOC_560/Y NAND2X1_LOC_388/A 0.01fF
C16901 INVX1_LOC_68/Y INVX1_LOC_145/Y 0.09fF
C16902 NAND2X1_LOC_336/B INVX1_LOC_686/A 0.00fF
C16903 INVX1_LOC_45/Y INVX1_LOC_509/A 0.13fF
C16904 INVX1_LOC_377/Y INVX1_LOC_375/Y 0.01fF
C16905 NAND2X1_LOC_33/a_36_24# INVX1_LOC_84/A 0.00fF
C16906 INVX1_LOC_395/Y INVX1_LOC_97/A 0.03fF
C16907 INVX1_LOC_308/Y INVX1_LOC_31/Y 0.03fF
C16908 NAND2X1_LOC_23/a_36_24# INVX1_LOC_6/Y 0.00fF
C16909 NAND2X1_LOC_467/A INVX1_LOC_186/A 0.00fF
C16910 INVX1_LOC_553/A INVX1_LOC_47/Y 0.03fF
C16911 INVX1_LOC_374/A INVX1_LOC_117/Y 0.03fF
C16912 NAND2X1_LOC_69/B INVX1_LOC_26/Y 0.00fF
C16913 INVX1_LOC_412/Y INVX1_LOC_65/A 0.02fF
C16914 INVX1_LOC_581/A NAND2X1_LOC_677/Y 0.02fF
C16915 INVX1_LOC_556/A INVX1_LOC_6/Y 1.01fF
C16916 INVX1_LOC_677/A INVX1_LOC_675/Y 0.00fF
C16917 INVX1_LOC_406/Y INVX1_LOC_451/A 0.00fF
C16918 NAND2X1_LOC_61/A NAND2X1_LOC_786/B 0.02fF
C16919 NAND2X1_LOC_543/B INVX1_LOC_242/Y 0.29fF
C16920 INVX1_LOC_103/Y INVX1_LOC_45/Y 0.37fF
C16921 INVX1_LOC_45/Y INVX1_LOC_68/A 0.01fF
C16922 NAND2X1_LOC_528/a_36_24# INVX1_LOC_379/A 0.00fF
C16923 INVX1_LOC_53/Y NAND2X1_LOC_755/B 0.03fF
C16924 INVX1_LOC_80/A INVX1_LOC_379/A 0.06fF
C16925 INVX1_LOC_435/Y INVX1_LOC_293/A 0.03fF
C16926 INVX1_LOC_235/Y INVX1_LOC_48/Y 0.01fF
C16927 INVX1_LOC_662/Y INVX1_LOC_101/Y 0.05fF
C16928 INVX1_LOC_80/A INVX1_LOC_35/Y 0.10fF
C16929 INVX1_LOC_671/A INVX1_LOC_654/A 0.02fF
C16930 INVX1_LOC_542/A INVX1_LOC_69/Y 0.07fF
C16931 INVX1_LOC_80/A INVX1_LOC_304/A 0.01fF
C16932 INVX1_LOC_97/A INVX1_LOC_179/Y 0.02fF
C16933 INVX1_LOC_145/Y INVX1_LOC_600/A 0.07fF
C16934 INVX1_LOC_320/A INVX1_LOC_304/Y 0.04fF
C16935 INVX1_LOC_553/A INVX1_LOC_119/Y 0.01fF
C16936 INVX1_LOC_272/Y NAND2X1_LOC_387/Y 0.01fF
C16937 NAND2X1_LOC_391/A INVX1_LOC_295/Y 0.00fF
C16938 INVX1_LOC_93/Y INVX1_LOC_492/Y 0.07fF
C16939 INVX1_LOC_370/Y INVX1_LOC_510/A 0.00fF
C16940 INVX1_LOC_400/A NAND2X1_LOC_72/Y 0.38fF
C16941 NAND2X1_LOC_707/A NAND2X1_LOC_334/A 0.16fF
C16942 NAND2X1_LOC_318/A INVX1_LOC_199/Y 0.34fF
C16943 INVX1_LOC_20/Y INVX1_LOC_96/A 0.25fF
C16944 INVX1_LOC_526/A INVX1_LOC_497/A 0.01fF
C16945 INVX1_LOC_31/Y NAND2X1_LOC_804/a_36_24# 0.00fF
C16946 INPUT_0 INVX1_LOC_369/Y 0.08fF
C16947 INVX1_LOC_89/Y INVX1_LOC_337/Y 0.05fF
C16948 INVX1_LOC_311/Y INVX1_LOC_6/Y 0.01fF
C16949 INVX1_LOC_53/Y INVX1_LOC_46/Y 0.69fF
C16950 INVX1_LOC_335/Y INVX1_LOC_315/A 0.03fF
C16951 INVX1_LOC_449/A INVX1_LOC_32/Y 0.10fF
C16952 NAND2X1_LOC_266/a_36_24# INVX1_LOC_194/Y 0.06fF
C16953 INVX1_LOC_7/Y INVX1_LOC_195/Y 0.03fF
C16954 INVX1_LOC_65/Y INVX1_LOC_245/A 0.18fF
C16955 INVX1_LOC_11/Y INVX1_LOC_379/A 0.19fF
C16956 NAND2X1_LOC_847/A INVX1_LOC_242/A 0.68fF
C16957 INVX1_LOC_32/Y INVX1_LOC_67/Y 0.16fF
C16958 INVX1_LOC_12/Y INVX1_LOC_87/A 0.00fF
C16959 INVX1_LOC_198/Y INVX1_LOC_145/Y 0.03fF
C16960 INVX1_LOC_11/Y INVX1_LOC_35/Y 1.37fF
C16961 INVX1_LOC_192/Y INVX1_LOC_62/Y 0.01fF
C16962 NAND2X1_LOC_325/B INVX1_LOC_93/Y 0.17fF
C16963 INVX1_LOC_602/A NAND2X1_LOC_836/B 0.25fF
C16964 INVX1_LOC_89/Y INVX1_LOC_633/Y 0.03fF
C16965 INVX1_LOC_80/A NAND2X1_LOC_253/Y 0.38fF
C16966 INVX1_LOC_17/Y INVX1_LOC_513/A 0.00fF
C16967 NAND2X1_LOC_331/A INVX1_LOC_479/A 0.05fF
C16968 INVX1_LOC_474/Y INVX1_LOC_633/A 0.16fF
C16969 INVX1_LOC_197/A INVX1_LOC_338/Y 0.07fF
C16970 NAND2X1_LOC_411/Y INVX1_LOC_6/Y 0.02fF
C16971 INPUT_3 INVX1_LOC_339/Y 0.01fF
C16972 INVX1_LOC_31/Y INVX1_LOC_230/A 0.07fF
C16973 INVX1_LOC_43/Y INVX1_LOC_6/Y 0.01fF
C16974 INVX1_LOC_268/Y INVX1_LOC_272/A 0.03fF
C16975 NAND2X1_LOC_140/B INVX1_LOC_47/Y 0.60fF
C16976 INVX1_LOC_40/Y INVX1_LOC_343/Y 0.01fF
C16977 INVX1_LOC_176/A NAND2X1_LOC_627/a_36_24# -0.01fF
C16978 INVX1_LOC_282/A INVX1_LOC_671/A 0.14fF
C16979 INVX1_LOC_369/A NAND2X1_LOC_615/Y 0.00fF
C16980 INVX1_LOC_62/A INVX1_LOC_50/Y 0.01fF
C16981 NAND2X1_LOC_320/Y INVX1_LOC_49/Y 0.01fF
C16982 INVX1_LOC_166/A INVX1_LOC_54/Y 0.30fF
C16983 INVX1_LOC_385/Y NAND2X1_LOC_480/a_36_24# 0.01fF
C16984 INVX1_LOC_11/Y NAND2X1_LOC_253/Y 0.01fF
C16985 INVX1_LOC_202/Y INVX1_LOC_199/Y 0.12fF
C16986 NAND2X1_LOC_308/A INVX1_LOC_61/A 0.00fF
C16987 INVX1_LOC_105/Y INVX1_LOC_108/A 0.01fF
C16988 INVX1_LOC_467/Y INVX1_LOC_463/Y 0.02fF
C16989 NAND2X1_LOC_399/B INVX1_LOC_328/Y 0.06fF
C16990 INVX1_LOC_400/A INVX1_LOC_351/Y 0.03fF
C16991 INVX1_LOC_287/A INVX1_LOC_245/A 0.00fF
C16992 INVX1_LOC_331/Y INVX1_LOC_137/Y 0.06fF
C16993 NAND2X1_LOC_250/Y INVX1_LOC_58/Y 0.01fF
C16994 INVX1_LOC_119/Y INVX1_LOC_375/Y 0.03fF
C16995 INVX1_LOC_63/Y INVX1_LOC_178/A 0.05fF
C16996 NAND2X1_LOC_97/B INVX1_LOC_90/Y 0.02fF
C16997 INVX1_LOC_6/Y INVX1_LOC_382/Y 0.01fF
C16998 INVX1_LOC_69/Y INVX1_LOC_259/Y 0.07fF
C16999 NAND2X1_LOC_532/Y INVX1_LOC_50/Y 0.01fF
C17000 INVX1_LOC_128/Y INVX1_LOC_383/Y 0.92fF
C17001 NAND2X1_LOC_538/B INVX1_LOC_75/Y 0.17fF
C17002 NAND2X1_LOC_708/a_36_24# INVX1_LOC_6/Y 0.00fF
C17003 NAND2X1_LOC_400/B INVX1_LOC_46/Y 0.01fF
C17004 INVX1_LOC_58/Y NAND2X1_LOC_646/A 0.00fF
C17005 NAND2X1_LOC_346/B INVX1_LOC_46/Y 0.03fF
C17006 INVX1_LOC_400/Y INVX1_LOC_92/A 0.03fF
C17007 INVX1_LOC_89/Y INVX1_LOC_317/A 0.02fF
C17008 INVX1_LOC_345/Y INVX1_LOC_347/Y 0.02fF
C17009 INVX1_LOC_80/A INVX1_LOC_79/Y 0.01fF
C17010 INVX1_LOC_520/Y INVX1_LOC_520/A 0.02fF
C17011 INVX1_LOC_463/Y NAND2X1_LOC_427/a_36_24# 0.00fF
C17012 INVX1_LOC_26/Y NAND2X1_LOC_226/a_36_24# 0.00fF
C17013 NAND2X1_LOC_628/a_36_24# INVX1_LOC_7/Y 0.00fF
C17014 INVX1_LOC_440/A INVX1_LOC_353/A 0.06fF
C17015 INVX1_LOC_93/Y INVX1_LOC_168/Y 0.05fF
C17016 INVX1_LOC_282/A INVX1_LOC_664/Y 0.01fF
C17017 NAND2X1_LOC_56/Y INVX1_LOC_211/A 0.05fF
C17018 INVX1_LOC_32/Y INVX1_LOC_328/Y 0.10fF
C17019 INVX1_LOC_53/A NAND2X1_LOC_409/Y 0.01fF
C17020 INVX1_LOC_49/Y INVX1_LOC_199/Y 0.60fF
C17021 INVX1_LOC_66/A INVX1_LOC_9/Y 0.90fF
C17022 INVX1_LOC_349/A INVX1_LOC_41/Y 0.01fF
C17023 INVX1_LOC_63/Y INVX1_LOC_58/Y 0.26fF
C17024 INVX1_LOC_62/Y INVX1_LOC_159/A 0.06fF
C17025 NAND2X1_LOC_274/B NAND2X1_LOC_469/a_36_24# 0.00fF
C17026 INVX1_LOC_54/Y INVX1_LOC_531/Y 0.07fF
C17027 NAND2X1_LOC_486/A INVX1_LOC_26/Y 0.16fF
C17028 INVX1_LOC_418/Y INVX1_LOC_75/Y 0.01fF
C17029 INVX1_LOC_62/Y NAND2X1_LOC_615/B 0.30fF
C17030 INVX1_LOC_525/Y INVX1_LOC_90/Y 0.01fF
C17031 INVX1_LOC_159/Y INVX1_LOC_75/Y 0.09fF
C17032 NAND2X1_LOC_846/B NAND2X1_LOC_816/a_36_24# 0.02fF
C17033 INVX1_LOC_69/Y INVX1_LOC_114/A 0.05fF
C17034 INVX1_LOC_49/Y INVX1_LOC_272/A 0.02fF
C17035 NAND2X1_LOC_444/A INVX1_LOC_74/Y 0.08fF
C17036 INVX1_LOC_379/A INVX1_LOC_231/Y 0.07fF
C17037 NAND2X1_LOC_543/B INVX1_LOC_301/A 0.07fF
C17038 INVX1_LOC_62/Y INVX1_LOC_66/A 0.39fF
C17039 INVX1_LOC_78/A INVX1_LOC_92/A 0.16fF
C17040 INVX1_LOC_54/Y NAND2X1_LOC_626/a_36_24# 0.01fF
C17041 INVX1_LOC_41/Y INVX1_LOC_420/A 0.01fF
C17042 INVX1_LOC_183/A INVX1_LOC_100/Y 0.03fF
C17043 NAND2X1_LOC_837/A INVX1_LOC_635/Y 0.13fF
C17044 INVX1_LOC_62/Y INVX1_LOC_296/A 0.01fF
C17045 INVX1_LOC_242/Y INVX1_LOC_353/A 0.01fF
C17046 INVX1_LOC_485/Y INVX1_LOC_90/Y 0.01fF
C17047 INVX1_LOC_54/Y INVX1_LOC_613/A 0.01fF
C17048 INVX1_LOC_133/Y INVX1_LOC_137/A 0.00fF
C17049 NAND2X1_LOC_475/A NAND2X1_LOC_310/a_36_24# 0.01fF
C17050 INVX1_LOC_50/Y INVX1_LOC_76/A 0.01fF
C17051 INVX1_LOC_183/A INVX1_LOC_483/Y 0.04fF
C17052 INVX1_LOC_554/A INVX1_LOC_76/Y 0.26fF
C17053 INVX1_LOC_549/A NAND2X1_LOC_707/a_36_24# 0.01fF
C17054 NAND2X1_LOC_833/B INVX1_LOC_479/A 0.12fF
C17055 INVX1_LOC_150/A NAND2X1_LOC_682/a_36_24# 0.01fF
C17056 VDD NAND2X1_LOC_773/A -0.00fF
C17057 NAND2X1_LOC_231/A INVX1_LOC_206/Y 0.01fF
C17058 NAND2X1_LOC_69/B INVX1_LOC_369/A 0.03fF
C17059 VDD NAND2X1_LOC_756/Y 0.07fF
C17060 NAND2X1_LOC_769/a_36_24# INVX1_LOC_366/A 0.00fF
C17061 VDD INVX1_LOC_293/Y 0.56fF
C17062 INVX1_LOC_62/Y NAND2X1_LOC_646/B 0.01fF
C17063 NAND2X1_LOC_780/B INVX1_LOC_581/A 0.07fF
C17064 INVX1_LOC_542/A INVX1_LOC_586/A 0.03fF
C17065 INVX1_LOC_395/A INVX1_LOC_492/Y 0.03fF
C17066 NAND2X1_LOC_336/B INVX1_LOC_390/Y 0.01fF
C17067 INVX1_LOC_410/Y INVX1_LOC_134/Y 0.07fF
C17068 INVX1_LOC_548/Y INVX1_LOC_53/Y 0.01fF
C17069 INVX1_LOC_127/A INVX1_LOC_519/A 0.21fF
C17070 INVX1_LOC_375/A INVX1_LOC_134/Y 0.03fF
C17071 INPUT_0 INVX1_LOC_558/Y 0.01fF
C17072 INVX1_LOC_546/A INVX1_LOC_134/Y 0.03fF
C17073 INVX1_LOC_205/Y INVX1_LOC_97/A 0.08fF
C17074 NAND2X1_LOC_637/A INVX1_LOC_259/Y 0.01fF
C17075 VDD NAND2X1_LOC_673/B 0.58fF
C17076 INVX1_LOC_581/A INVX1_LOC_137/A 0.03fF
C17077 NAND2X1_LOC_505/Y NAND2X1_LOC_237/Y 0.05fF
C17078 NAND2X1_LOC_715/a_36_24# INVX1_LOC_80/A 0.01fF
C17079 INVX1_LOC_579/A NAND2X1_LOC_122/Y 0.97fF
C17080 INVX1_LOC_51/Y INVX1_LOC_635/A 0.10fF
C17081 INVX1_LOC_564/Y INVX1_LOC_155/Y 0.16fF
C17082 INVX1_LOC_395/A INVX1_LOC_681/A 0.00fF
C17083 NAND2X1_LOC_88/B INVX1_LOC_88/Y 0.18fF
C17084 INVX1_LOC_552/Y INVX1_LOC_178/A 0.03fF
C17085 INVX1_LOC_564/A INVX1_LOC_35/Y 0.00fF
C17086 INVX1_LOC_53/Y INVX1_LOC_268/Y 0.03fF
C17087 NAND2X1_LOC_320/Y NAND2X1_LOC_498/B 0.01fF
C17088 INVX1_LOC_584/Y NAND2X1_LOC_210/A 0.00fF
C17089 NAND2X1_LOC_130/Y NAND2X1_LOC_332/B 0.05fF
C17090 INVX1_LOC_291/A INVX1_LOC_80/A 0.01fF
C17091 INVX1_LOC_435/Y NAND2X1_LOC_106/B 0.34fF
C17092 INVX1_LOC_118/Y NAND2X1_LOC_706/B 0.01fF
C17093 NAND2X1_LOC_525/Y INVX1_LOC_392/A 0.04fF
C17094 INVX1_LOC_406/Y INVX1_LOC_134/Y 0.00fF
C17095 INVX1_LOC_424/A NAND2X1_LOC_346/B 0.03fF
C17096 NAND2X1_LOC_45/Y NAND2X1_LOC_106/Y 0.04fF
C17097 INVX1_LOC_23/Y INVX1_LOC_21/A 0.19fF
C17098 INVX1_LOC_360/Y INVX1_LOC_45/Y 0.07fF
C17099 INVX1_LOC_256/Y INVX1_LOC_80/A 0.01fF
C17100 NAND2X1_LOC_548/B NAND2X1_LOC_530/a_36_24# 0.02fF
C17101 INVX1_LOC_20/Y INVX1_LOC_469/A 0.01fF
C17102 INVX1_LOC_400/Y INPUT_1 0.04fF
C17103 NAND2X1_LOC_759/B INVX1_LOC_44/Y 0.06fF
C17104 INVX1_LOC_617/Y INVX1_LOC_370/Y 0.01fF
C17105 VDD NAND2X1_LOC_240/A -0.00fF
C17106 INVX1_LOC_171/A INVX1_LOC_45/Y 0.01fF
C17107 INVX1_LOC_211/Y NAND2X1_LOC_383/Y 0.00fF
C17108 INVX1_LOC_586/A INVX1_LOC_259/Y 0.03fF
C17109 INVX1_LOC_401/A INVX1_LOC_99/Y 0.35fF
C17110 NAND2X1_LOC_457/A INVX1_LOC_69/Y 0.00fF
C17111 INVX1_LOC_563/A INVX1_LOC_53/Y 0.08fF
C17112 INPUT_0 NAND2X1_LOC_531/Y 0.22fF
C17113 INVX1_LOC_206/Y INVX1_LOC_77/Y 0.01fF
C17114 INVX1_LOC_395/A NAND2X1_LOC_647/A 0.02fF
C17115 INVX1_LOC_224/Y NAND2X1_LOC_212/a_36_24# 0.00fF
C17116 INVX1_LOC_583/Y INVX1_LOC_93/Y 0.01fF
C17117 NAND2X1_LOC_862/a_36_24# INVX1_LOC_367/A 0.00fF
C17118 NAND2X1_LOC_322/Y INVX1_LOC_242/Y 0.03fF
C17119 NAND2X1_LOC_586/a_36_24# INVX1_LOC_288/A 0.00fF
C17120 INVX1_LOC_566/Y INVX1_LOC_35/Y 0.03fF
C17121 INVX1_LOC_266/Y INVX1_LOC_32/Y 0.36fF
C17122 INVX1_LOC_97/A INVX1_LOC_44/Y 0.02fF
C17123 NAND2X1_LOC_56/Y INVX1_LOC_145/Y 0.01fF
C17124 INVX1_LOC_293/Y NAND2X1_LOC_843/A 0.02fF
C17125 INVX1_LOC_547/Y INVX1_LOC_69/Y 0.02fF
C17126 INVX1_LOC_31/Y INVX1_LOC_666/A 0.00fF
C17127 NAND2X1_LOC_383/Y INVX1_LOC_46/Y 0.19fF
C17128 INVX1_LOC_317/Y INVX1_LOC_89/Y 0.00fF
C17129 NAND2X1_LOC_638/A INVX1_LOC_300/A 0.07fF
C17130 INVX1_LOC_214/Y INVX1_LOC_80/A 0.00fF
C17131 INVX1_LOC_395/A INVX1_LOC_168/Y 0.00fF
C17132 INVX1_LOC_250/Y INVX1_LOC_440/A 0.05fF
C17133 NAND2X1_LOC_336/B INVX1_LOC_432/A 0.00fF
C17134 INVX1_LOC_550/Y INVX1_LOC_53/Y 0.01fF
C17135 INVX1_LOC_417/A INVX1_LOC_98/Y 0.07fF
C17136 INVX1_LOC_84/A INVX1_LOC_117/Y 0.54fF
C17137 INVX1_LOC_21/Y INVX1_LOC_176/A 0.08fF
C17138 INVX1_LOC_293/Y INVX1_LOC_103/Y 0.03fF
C17139 INVX1_LOC_61/A INVX1_LOC_134/Y 0.12fF
C17140 INVX1_LOC_425/Y INVX1_LOC_12/Y 0.02fF
C17141 INVX1_LOC_444/Y INVX1_LOC_385/Y 0.03fF
C17142 INVX1_LOC_12/Y INVX1_LOC_480/Y 0.01fF
C17143 NAND2X1_LOC_184/Y INVX1_LOC_661/A 0.01fF
C17144 INVX1_LOC_558/A INVX1_LOC_544/Y 0.01fF
C17145 INVX1_LOC_27/A NAND2X1_LOC_84/B 0.09fF
C17146 INPUT_0 NAND2X1_LOC_628/Y 0.16fF
C17147 INVX1_LOC_158/Y INVX1_LOC_160/A 0.00fF
C17148 INVX1_LOC_562/Y INVX1_LOC_47/Y 0.01fF
C17149 INVX1_LOC_53/Y INVX1_LOC_550/A 0.02fF
C17150 INVX1_LOC_80/A INVX1_LOC_118/A 0.00fF
C17151 NAND2X1_LOC_578/a_36_24# INVX1_LOC_385/Y 0.01fF
C17152 INVX1_LOC_625/A INVX1_LOC_201/Y 0.02fF
C17153 INVX1_LOC_31/Y NAND2X1_LOC_273/a_36_24# 0.00fF
C17154 INVX1_LOC_76/Y INVX1_LOC_199/Y 0.13fF
C17155 INVX1_LOC_442/A INVX1_LOC_9/Y 0.07fF
C17156 INVX1_LOC_53/Y NAND2X1_LOC_213/a_36_24# 0.00fF
C17157 INVX1_LOC_376/Y INVX1_LOC_618/Y 0.00fF
C17158 NAND2X1_LOC_322/a_36_24# INVX1_LOC_257/A 0.00fF
C17159 NAND2X1_LOC_22/a_36_24# NAND2X1_LOC_836/B 0.00fF
C17160 INVX1_LOC_310/Y INVX1_LOC_48/Y 0.03fF
C17161 INVX1_LOC_236/A INVX1_LOC_35/Y 0.01fF
C17162 NAND2X1_LOC_399/B INVX1_LOC_172/A 0.09fF
C17163 INVX1_LOC_230/A NAND2X1_LOC_267/a_36_24# 0.02fF
C17164 NAND2X1_LOC_148/A INVX1_LOC_46/Y 0.00fF
C17165 INVX1_LOC_344/Y INVX1_LOC_50/Y 0.00fF
C17166 INVX1_LOC_557/A NAND2X1_LOC_274/B 0.04fF
C17167 INVX1_LOC_289/A INVX1_LOC_259/Y 0.20fF
C17168 INVX1_LOC_172/A INVX1_LOC_7/Y 0.07fF
C17169 INVX1_LOC_53/Y INVX1_LOC_387/Y 0.03fF
C17170 INVX1_LOC_12/Y INVX1_LOC_169/Y 0.07fF
C17171 INVX1_LOC_11/Y INVX1_LOC_214/Y 0.01fF
C17172 INVX1_LOC_511/Y INVX1_LOC_522/A 0.01fF
C17173 INVX1_LOC_69/Y INVX1_LOC_651/A 0.00fF
C17174 INVX1_LOC_358/A INVX1_LOC_463/Y 0.26fF
C17175 INVX1_LOC_249/A INVX1_LOC_89/Y 0.01fF
C17176 INVX1_LOC_278/Y INVX1_LOC_282/A 0.01fF
C17177 INVX1_LOC_93/Y INVX1_LOC_99/A 0.04fF
C17178 INVX1_LOC_68/Y INVX1_LOC_242/Y 0.00fF
C17179 NAND2X1_LOC_336/B NAND2X1_LOC_542/A 0.00fF
C17180 INVX1_LOC_612/Y INVX1_LOC_609/A 0.13fF
C17181 INVX1_LOC_408/Y INVX1_LOC_62/Y 0.01fF
C17182 NAND2X1_LOC_137/A INVX1_LOC_680/Y 0.01fF
C17183 INVX1_LOC_31/Y NAND2X1_LOC_72/Y 0.08fF
C17184 INVX1_LOC_131/Y INVX1_LOC_655/A 0.01fF
C17185 INVX1_LOC_401/Y INVX1_LOC_338/Y 0.05fF
C17186 INVX1_LOC_361/Y INVX1_LOC_251/A 0.01fF
C17187 INPUT_5 INVX1_LOC_59/A 0.01fF
C17188 NAND2X1_LOC_321/a_36_24# INVX1_LOC_69/Y 0.01fF
C17189 INVX1_LOC_53/Y INVX1_LOC_49/Y 0.36fF
C17190 NAND2X1_LOC_586/a_36_24# INVX1_LOC_145/Y 0.01fF
C17191 NAND2X1_LOC_636/B INVX1_LOC_496/A 0.05fF
C17192 NAND2X1_LOC_106/Y INVX1_LOC_99/Y 0.04fF
C17193 NAND2X1_LOC_700/a_36_24# INVX1_LOC_376/Y 0.00fF
C17194 INVX1_LOC_442/A INVX1_LOC_62/Y 0.01fF
C17195 INVX1_LOC_20/Y INVX1_LOC_353/A 0.08fF
C17196 INVX1_LOC_93/Y INVX1_LOC_137/Y 2.57fF
C17197 INVX1_LOC_31/Y NAND2X1_LOC_673/A 0.02fF
C17198 INVX1_LOC_172/A INVX1_LOC_32/Y 0.59fF
C17199 INVX1_LOC_366/A INVX1_LOC_190/A 0.29fF
C17200 INVX1_LOC_250/Y INVX1_LOC_242/Y 0.05fF
C17201 INVX1_LOC_492/A INVX1_LOC_212/Y 0.26fF
C17202 NAND2X1_LOC_294/Y INVX1_LOC_382/Y 0.01fF
C17203 INVX1_LOC_527/Y INVX1_LOC_187/Y 0.01fF
C17204 INVX1_LOC_109/Y INVX1_LOC_192/A 0.00fF
C17205 INVX1_LOC_189/Y INVX1_LOC_168/Y 0.04fF
C17206 INVX1_LOC_161/A INVX1_LOC_491/A 0.03fF
C17207 NAND2X1_LOC_635/B INVX1_LOC_261/Y 0.01fF
C17208 INVX1_LOC_196/A INVX1_LOC_62/Y 0.01fF
C17209 INVX1_LOC_116/Y INVX1_LOC_9/Y 0.03fF
C17210 INVX1_LOC_166/A INVX1_LOC_89/Y 0.04fF
C17211 NAND2X1_LOC_274/a_36_24# INVX1_LOC_420/A 0.01fF
C17212 NAND2X1_LOC_672/a_36_24# INVX1_LOC_63/Y 0.00fF
C17213 INVX1_LOC_300/A INVX1_LOC_353/A 0.07fF
C17214 INVX1_LOC_58/Y INVX1_LOC_263/Y 0.05fF
C17215 NAND2X1_LOC_498/Y INVX1_LOC_92/A 0.07fF
C17216 INVX1_LOC_117/Y INVX1_LOC_496/A 0.08fF
C17217 INVX1_LOC_468/Y NAND2X1_LOC_274/B 0.01fF
C17218 INVX1_LOC_353/A INVX1_LOC_197/Y 0.07fF
C17219 NAND2X1_LOC_111/Y NAND2X1_LOC_111/a_36_24# 0.02fF
C17220 INVX1_LOC_570/A INVX1_LOC_92/A 0.01fF
C17221 INVX1_LOC_304/Y NAND2X1_LOC_558/B 0.35fF
C17222 INVX1_LOC_675/A INVX1_LOC_355/Y 0.07fF
C17223 NAND2X1_LOC_111/Y INVX1_LOC_89/Y 0.05fF
C17224 NAND2X1_LOC_123/B INVX1_LOC_99/Y 0.03fF
C17225 INVX1_LOC_137/Y NAND2X1_LOC_9/a_36_24# 0.01fF
C17226 INVX1_LOC_80/A INVX1_LOC_364/A 0.00fF
C17227 INVX1_LOC_66/A INVX1_LOC_624/Y 0.03fF
C17228 INVX1_LOC_328/A INVX1_LOC_9/Y 0.13fF
C17229 INVX1_LOC_35/Y INVX1_LOC_319/A 0.01fF
C17230 INVX1_LOC_304/Y INVX1_LOC_79/A 1.38fF
C17231 INVX1_LOC_49/Y NAND2X1_LOC_346/B 0.01fF
C17232 INVX1_LOC_662/A INVX1_LOC_46/Y 0.03fF
C17233 INVX1_LOC_676/Y NAND2X1_LOC_428/Y 0.10fF
C17234 INVX1_LOC_62/Y INVX1_LOC_116/Y 0.00fF
C17235 INVX1_LOC_49/Y NAND2X1_LOC_274/Y 0.00fF
C17236 INVX1_LOC_288/Y INVX1_LOC_74/Y 0.01fF
C17237 INVX1_LOC_329/Y INVX1_LOC_99/Y 0.01fF
C17238 NAND2X1_LOC_137/A INVX1_LOC_124/A 0.06fF
C17239 INVX1_LOC_35/Y NAND2X1_LOC_843/B 0.04fF
C17240 NAND2X1_LOC_187/Y INVX1_LOC_41/Y 0.29fF
C17241 INVX1_LOC_585/Y INVX1_LOC_531/Y 0.01fF
C17242 INVX1_LOC_479/A INVX1_LOC_685/Y 0.31fF
C17243 INVX1_LOC_54/Y INVX1_LOC_41/Y 3.40fF
C17244 INVX1_LOC_63/Y NAND2X1_LOC_440/A 0.03fF
C17245 NAND2X1_LOC_507/A INVX1_LOC_531/Y 0.06fF
C17246 INVX1_LOC_89/Y NAND2X1_LOC_136/Y 0.61fF
C17247 NAND2X1_LOC_677/Y INVX1_LOC_613/A 0.31fF
C17248 INVX1_LOC_154/A INVX1_LOC_153/Y 0.04fF
C17249 INVX1_LOC_17/Y INVX1_LOC_282/Y 0.01fF
C17250 INVX1_LOC_63/Y INVX1_LOC_245/A 0.10fF
C17251 INVX1_LOC_35/Y INVX1_LOC_91/Y 0.00fF
C17252 NAND2X1_LOC_416/Y NAND2X1_LOC_416/B 0.00fF
C17253 INVX1_LOC_656/A INVX1_LOC_635/Y 0.01fF
C17254 NAND2X1_LOC_520/A INVX1_LOC_502/A -0.02fF
C17255 INVX1_LOC_89/Y INVX1_LOC_531/Y 0.02fF
C17256 INVX1_LOC_47/Y NAND2X1_LOC_123/B 0.07fF
C17257 NAND2X1_LOC_292/Y INVX1_LOC_41/Y 0.02fF
C17258 INVX1_LOC_257/A INVX1_LOC_41/Y 0.16fF
C17259 INVX1_LOC_99/Y INVX1_LOC_92/A 0.03fF
C17260 INVX1_LOC_58/Y INVX1_LOC_669/A 0.00fF
C17261 NAND2X1_LOC_308/A INVX1_LOC_479/A 0.11fF
C17262 INPUT_0 INVX1_LOC_180/Y 0.08fF
C17263 INVX1_LOC_620/A INVX1_LOC_91/Y 0.01fF
C17264 NAND2X1_LOC_123/B INVX1_LOC_119/Y 0.07fF
C17265 NAND2X1_LOC_750/Y INPUT_0 1.14fF
C17266 INVX1_LOC_261/Y INVX1_LOC_462/Y 0.03fF
C17267 INVX1_LOC_568/A INVX1_LOC_92/A 0.01fF
C17268 INVX1_LOC_151/Y INVX1_LOC_542/A 0.01fF
C17269 INVX1_LOC_395/A NAND2X1_LOC_749/Y 0.07fF
C17270 INVX1_LOC_47/Y INVX1_LOC_92/A 0.07fF
C17271 INVX1_LOC_601/A NAND2X1_LOC_79/B 0.04fF
C17272 NAND2X1_LOC_76/a_36_24# INVX1_LOC_206/Y 0.00fF
C17273 INVX1_LOC_20/Y INVX1_LOC_409/Y 0.01fF
C17274 INVX1_LOC_372/Y INVX1_LOC_638/A 0.01fF
C17275 NAND2X1_LOC_457/A INVX1_LOC_586/A 0.03fF
C17276 INVX1_LOC_20/Y NAND2X1_LOC_335/B 0.01fF
C17277 INVX1_LOC_75/Y NAND2X1_LOC_372/Y 0.02fF
C17278 INVX1_LOC_100/Y NAND2X1_LOC_237/a_36_24# 0.00fF
C17279 INVX1_LOC_224/Y NAND2X1_LOC_538/B 0.07fF
C17280 NAND2X1_LOC_525/Y INVX1_LOC_362/Y 0.01fF
C17281 NAND2X1_LOC_751/a_36_24# INVX1_LOC_191/A 0.00fF
C17282 INVX1_LOC_45/Y NAND2X1_LOC_506/B 0.09fF
C17283 INVX1_LOC_429/Y INVX1_LOC_220/Y 0.18fF
C17284 INVX1_LOC_119/Y INVX1_LOC_92/A 0.03fF
C17285 INVX1_LOC_257/Y INVX1_LOC_258/A 0.01fF
C17286 NAND2X1_LOC_231/A INVX1_LOC_94/A 0.02fF
C17287 INVX1_LOC_280/A NAND2X1_LOC_271/A 0.07fF
C17288 INVX1_LOC_11/Y INVX1_LOC_220/A 0.02fF
C17289 NAND2X1_LOC_335/B INVX1_LOC_300/A 0.03fF
C17290 INVX1_LOC_20/Y INVX1_LOC_68/Y 0.03fF
C17291 INVX1_LOC_206/Y INVX1_LOC_683/A 0.01fF
C17292 INVX1_LOC_210/Y VDD 0.49fF
C17293 INPUT_3 INVX1_LOC_45/Y 0.60fF
C17294 INVX1_LOC_561/Y INVX1_LOC_565/A 0.00fF
C17295 INVX1_LOC_3/Y INVX1_LOC_595/Y 0.01fF
C17296 INPUT_0 NAND2X1_LOC_413/Y 0.34fF
C17297 INVX1_LOC_370/Y INVX1_LOC_410/Y 0.03fF
C17298 INVX1_LOC_586/A NAND2X1_LOC_635/a_36_24# 0.01fF
C17299 INVX1_LOC_395/A INVX1_LOC_99/A 0.17fF
C17300 INVX1_LOC_412/Y INVX1_LOC_98/Y 0.03fF
C17301 INVX1_LOC_607/Y INVX1_LOC_606/Y 0.06fF
C17302 NAND2X1_LOC_516/Y NAND2X1_LOC_413/Y 0.02fF
C17303 INVX1_LOC_312/Y INVX1_LOC_482/A 0.33fF
C17304 INVX1_LOC_224/Y INVX1_LOC_159/Y 0.03fF
C17305 INVX1_LOC_402/A INVX1_LOC_558/A 0.04fF
C17306 INVX1_LOC_405/A NAND2X1_LOC_271/a_36_24# 0.00fF
C17307 NAND2X1_LOC_45/Y INPUT_1 0.05fF
C17308 INVX1_LOC_428/A INVX1_LOC_145/Y 0.03fF
C17309 INVX1_LOC_53/Y INVX1_LOC_76/Y 0.04fF
C17310 INVX1_LOC_395/A INVX1_LOC_137/Y 0.07fF
C17311 INVX1_LOC_20/Y INVX1_LOC_250/Y 0.03fF
C17312 NAND2X1_LOC_176/Y INVX1_LOC_317/A 0.01fF
C17313 INVX1_LOC_418/Y INVX1_LOC_578/A 0.02fF
C17314 INVX1_LOC_33/Y INVX1_LOC_145/Y 0.05fF
C17315 INVX1_LOC_584/A INVX1_LOC_50/Y 0.02fF
C17316 NAND2X1_LOC_773/A INVX1_LOC_619/A 0.04fF
C17317 INVX1_LOC_68/Y INVX1_LOC_300/A 0.08fF
C17318 INVX1_LOC_578/A INVX1_LOC_159/Y 0.00fF
C17319 INVX1_LOC_20/Y NAND2X1_LOC_130/Y 0.93fF
C17320 INVX1_LOC_20/Y INVX1_LOC_600/A 0.24fF
C17321 INVX1_LOC_68/Y INVX1_LOC_197/Y 0.03fF
C17322 INVX1_LOC_36/A INPUT_1 0.01fF
C17323 INVX1_LOC_194/A INVX1_LOC_586/A 0.02fF
C17324 INVX1_LOC_266/A NAND2X1_LOC_325/B 0.06fF
C17325 VDD NAND2X1_LOC_344/B 0.20fF
C17326 INVX1_LOC_400/Y INVX1_LOC_50/Y 0.29fF
C17327 INVX1_LOC_560/Y INVX1_LOC_58/Y 0.05fF
C17328 NAND2X1_LOC_788/A INVX1_LOC_624/Y 0.00fF
C17329 NAND2X1_LOC_498/Y INPUT_1 0.17fF
C17330 INVX1_LOC_182/A INVX1_LOC_86/Y 0.02fF
C17331 INVX1_LOC_255/Y INVX1_LOC_354/Y 0.02fF
C17332 NAND2X1_LOC_13/Y INVX1_LOC_230/A 0.07fF
C17333 NAND2X1_LOC_156/Y INVX1_LOC_522/Y 0.05fF
C17334 INVX1_LOC_288/A INVX1_LOC_359/Y 0.01fF
C17335 INVX1_LOC_543/Y INVX1_LOC_65/Y 0.01fF
C17336 VDD INVX1_LOC_262/Y 0.21fF
C17337 INVX1_LOC_561/Y NAND2X1_LOC_586/Y 0.00fF
C17338 INVX1_LOC_84/A INVX1_LOC_178/A 0.07fF
C17339 INVX1_LOC_567/Y INVX1_LOC_136/Y 0.01fF
C17340 INVX1_LOC_581/A INVX1_LOC_610/A -0.02fF
C17341 VDD INVX1_LOC_117/A -0.00fF
C17342 INVX1_LOC_596/A INVX1_LOC_510/A 0.03fF
C17343 NAND2X1_LOC_57/Y INVX1_LOC_174/A 0.00fF
C17344 NAND2X1_LOC_338/a_36_24# NAND2X1_LOC_720/A 0.00fF
C17345 INVX1_LOC_250/Y INVX1_LOC_197/Y 0.05fF
C17346 INVX1_LOC_679/Y INVX1_LOC_99/Y 0.09fF
C17347 INVX1_LOC_406/A INVX1_LOC_362/Y 0.14fF
C17348 INVX1_LOC_80/A INVX1_LOC_350/A 0.00fF
C17349 INVX1_LOC_377/Y INPUT_1 0.32fF
C17350 INVX1_LOC_442/A INVX1_LOC_624/Y 0.01fF
C17351 NAND2X1_LOC_218/a_36_24# INVX1_LOC_390/A 0.00fF
C17352 INVX1_LOC_206/Y NAND2X1_LOC_274/B 0.03fF
C17353 INVX1_LOC_288/Y NAND2X1_LOC_856/a_36_24# 0.00fF
C17354 INVX1_LOC_565/Y INVX1_LOC_674/A 0.05fF
C17355 INVX1_LOC_417/Y INVX1_LOC_304/Y 0.09fF
C17356 INVX1_LOC_512/A INVX1_LOC_58/Y 0.01fF
C17357 NAND2X1_LOC_516/B NAND2X1_LOC_307/B 0.04fF
C17358 INVX1_LOC_374/A NAND2X1_LOC_440/A 0.01fF
C17359 INVX1_LOC_599/A INVX1_LOC_623/Y 0.01fF
C17360 NAND2X1_LOC_67/Y INVX1_LOC_178/A 0.01fF
C17361 INVX1_LOC_410/Y INVX1_LOC_90/Y 0.03fF
C17362 INVX1_LOC_93/Y NAND2X1_LOC_307/A 0.12fF
C17363 INVX1_LOC_435/A INVX1_LOC_17/Y 0.07fF
C17364 INVX1_LOC_686/A INVX1_LOC_372/A 0.03fF
C17365 NAND2X1_LOC_698/Y NAND2X1_LOC_318/A 0.03fF
C17366 INVX1_LOC_556/A INVX1_LOC_100/Y 0.08fF
C17367 INVX1_LOC_53/Y INVX1_LOC_108/A 0.00fF
C17368 INVX1_LOC_140/Y INVX1_LOC_114/A 0.02fF
C17369 INVX1_LOC_449/A NAND2X1_LOC_184/Y -0.04fF
C17370 INVX1_LOC_21/Y INVX1_LOC_54/Y 2.20fF
C17371 NAND2X1_LOC_775/B INVX1_LOC_252/Y 3.04fF
C17372 INVX1_LOC_238/Y INVX1_LOC_479/A 0.01fF
C17373 INVX1_LOC_272/Y INVX1_LOC_204/Y 0.00fF
C17374 INVX1_LOC_254/A NAND2X1_LOC_72/Y 0.01fF
C17375 INVX1_LOC_99/Y INPUT_1 0.11fF
C17376 INVX1_LOC_84/A INVX1_LOC_58/Y 0.03fF
C17377 INVX1_LOC_146/A INVX1_LOC_9/Y 0.07fF
C17378 VDD INVX1_LOC_622/Y 0.21fF
C17379 INVX1_LOC_304/Y INVX1_LOC_48/Y 0.00fF
C17380 NAND2X1_LOC_750/Y INVX1_LOC_64/Y 0.00fF
C17381 INVX1_LOC_595/Y INVX1_LOC_48/Y 0.01fF
C17382 INVX1_LOC_35/Y NAND2X1_LOC_333/B 0.02fF
C17383 INVX1_LOC_361/Y INVX1_LOC_35/Y 0.30fF
C17384 NAND2X1_LOC_274/B INVX1_LOC_242/A 0.03fF
C17385 NAND2X1_LOC_299/Y INVX1_LOC_347/Y 0.15fF
C17386 INVX1_LOC_210/Y NAND2X1_LOC_243/A 0.00fF
C17387 INVX1_LOC_402/Y NAND2X1_LOC_307/B 0.03fF
C17388 NAND2X1_LOC_27/Y INVX1_LOC_86/Y 0.00fF
C17389 INVX1_LOC_619/A NAND2X1_LOC_240/A 0.07fF
C17390 NAND2X1_LOC_98/a_36_24# NAND2X1_LOC_98/B 0.00fF
C17391 INVX1_LOC_571/A NAND2X1_LOC_728/A 0.00fF
C17392 NAND2X1_LOC_107/Y NAND2X1_LOC_107/a_36_24# 0.02fF
C17393 NAND2X1_LOC_331/A NAND2X1_LOC_646/B 0.01fF
C17394 INVX1_LOC_31/Y INVX1_LOC_137/Y 0.00fF
C17395 NAND2X1_LOC_475/A INVX1_LOC_270/Y 0.01fF
C17396 INVX1_LOC_419/Y INVX1_LOC_93/Y 0.01fF
C17397 INVX1_LOC_53/Y NAND2X1_LOC_816/a_36_24# 0.00fF
C17398 INVX1_LOC_395/A INVX1_LOC_647/Y 0.05fF
C17399 INVX1_LOC_62/A INVX1_LOC_117/Y 0.03fF
C17400 INVX1_LOC_6/Y INVX1_LOC_453/Y 0.06fF
C17401 INVX1_LOC_206/Y NAND2X1_LOC_449/a_36_24# 0.01fF
C17402 INVX1_LOC_116/Y INVX1_LOC_624/Y 0.00fF
C17403 NAND2X1_LOC_836/B INVX1_LOC_1/Y 0.11fF
C17404 INVX1_LOC_58/Y NAND2X1_LOC_67/Y 0.02fF
C17405 INVX1_LOC_298/A INVX1_LOC_341/Y 0.00fF
C17406 INVX1_LOC_76/Y INVX1_LOC_368/Y 0.01fF
C17407 NAND2X1_LOC_475/A INVX1_LOC_92/A 0.09fF
C17408 INVX1_LOC_446/Y INVX1_LOC_443/A 0.41fF
C17409 INVX1_LOC_54/Y INVX1_LOC_555/A 0.07fF
C17410 INVX1_LOC_620/A NAND2X1_LOC_333/B 0.03fF
C17411 NAND2X1_LOC_180/B INVX1_LOC_74/Y 0.28fF
C17412 NAND2X1_LOC_532/Y INVX1_LOC_117/Y 0.04fF
C17413 NAND2X1_LOC_759/a_36_24# NAND2X1_LOC_759/Y 0.02fF
C17414 INVX1_LOC_602/A NAND2X1_LOC_409/Y 0.02fF
C17415 INVX1_LOC_98/A NAND2X1_LOC_230/a_36_24# 0.00fF
C17416 INVX1_LOC_47/Y INPUT_1 0.21fF
C17417 INVX1_LOC_120/Y INVX1_LOC_159/Y 0.02fF
C17418 INVX1_LOC_587/Y INVX1_LOC_69/Y 0.01fF
C17419 NAND2X1_LOC_27/Y INVX1_LOC_63/Y 0.01fF
C17420 NAND2X1_LOC_376/B INVX1_LOC_117/Y 0.06fF
C17421 NAND2X1_LOC_411/Y INVX1_LOC_100/Y 0.08fF
C17422 INVX1_LOC_406/A INVX1_LOC_31/Y 0.00fF
C17423 INVX1_LOC_671/A INVX1_LOC_654/Y 0.02fF
C17424 INVX1_LOC_11/Y INVX1_LOC_223/Y 0.09fF
C17425 INVX1_LOC_32/Y INVX1_LOC_199/Y 0.11fF
C17426 NAND2X1_LOC_584/a_36_24# INVX1_LOC_62/Y 0.00fF
C17427 INVX1_LOC_384/A INVX1_LOC_443/A 0.31fF
C17428 NAND2X1_LOC_529/Y INVX1_LOC_422/A 0.14fF
C17429 INVX1_LOC_134/Y INVX1_LOC_479/A 0.21fF
C17430 INVX1_LOC_598/A NAND2X1_LOC_792/a_36_24# 0.00fF
C17431 INVX1_LOC_291/A INVX1_LOC_91/Y 0.01fF
C17432 INVX1_LOC_188/Y INVX1_LOC_74/Y 0.03fF
C17433 INVX1_LOC_93/Y INVX1_LOC_376/A 0.07fF
C17434 INVX1_LOC_186/A NAND2X1_LOC_210/a_36_24# 0.00fF
C17435 INVX1_LOC_449/A INVX1_LOC_75/Y 0.01fF
C17436 INVX1_LOC_103/Y INVX1_LOC_682/A 0.00fF
C17437 INVX1_LOC_468/Y INVX1_LOC_468/A 0.09fF
C17438 NAND2X1_LOC_452/a_36_24# INVX1_LOC_463/Y 0.00fF
C17439 INVX1_LOC_531/Y INVX1_LOC_194/Y 0.05fF
C17440 NAND2X1_LOC_645/a_36_24# INVX1_LOC_74/Y 0.00fF
C17441 INPUT_1 INVX1_LOC_119/Y 0.06fF
C17442 INVX1_LOC_670/A NAND2X1_LOC_657/a_36_24# 0.01fF
C17443 INVX1_LOC_58/Y INVX1_LOC_496/A 0.01fF
C17444 NAND2X1_LOC_297/Y INVX1_LOC_369/Y 0.06fF
C17445 INVX1_LOC_58/Y INVX1_LOC_674/Y 0.03fF
C17446 INVX1_LOC_214/Y NAND2X1_LOC_843/B 0.01fF
C17447 INVX1_LOC_285/Y INVX1_LOC_69/Y 0.01fF
C17448 NAND2X1_LOC_387/Y INVX1_LOC_100/Y 0.01fF
C17449 INVX1_LOC_93/Y INVX1_LOC_502/A 0.07fF
C17450 INVX1_LOC_69/Y INVX1_LOC_9/Y 0.10fF
C17451 INVX1_LOC_11/A INVX1_LOC_83/Y 0.04fF
C17452 INVX1_LOC_585/Y INVX1_LOC_41/Y 0.02fF
C17453 INVX1_LOC_478/Y INVX1_LOC_74/Y 0.01fF
C17454 INVX1_LOC_534/Y INVX1_LOC_69/Y 0.60fF
C17455 NAND2X1_LOC_545/A INVX1_LOC_46/Y 0.22fF
C17456 INVX1_LOC_386/A INVX1_LOC_63/Y 0.01fF
C17457 INVX1_LOC_136/Y INVX1_LOC_92/A 0.06fF
C17458 INVX1_LOC_465/Y INVX1_LOC_463/A 0.02fF
C17459 INVX1_LOC_653/A INVX1_LOC_49/Y 0.01fF
C17460 INVX1_LOC_26/Y INVX1_LOC_420/A 0.01fF
C17461 INVX1_LOC_89/Y INVX1_LOC_41/Y 0.29fF
C17462 NAND2X1_LOC_322/Y NAND2X1_LOC_373/Y 0.29fF
C17463 INVX1_LOC_166/Y INVX1_LOC_69/Y 0.01fF
C17464 INVX1_LOC_154/A INVX1_LOC_41/Y 0.03fF
C17465 INVX1_LOC_327/A INVX1_LOC_46/Y 0.01fF
C17466 INVX1_LOC_46/Y INVX1_LOC_666/Y 0.03fF
C17467 INVX1_LOC_69/Y INVX1_LOC_62/Y 0.15fF
C17468 INVX1_LOC_399/Y INVX1_LOC_26/Y -0.00fF
C17469 INVX1_LOC_100/Y NAND2X1_LOC_845/B 0.02fF
C17470 INVX1_LOC_501/A INVX1_LOC_41/Y 0.02fF
C17471 INPUT_0 VDD 0.60fF
C17472 INVX1_LOC_443/A INVX1_LOC_433/A 0.05fF
C17473 INVX1_LOC_117/Y INVX1_LOC_76/A 0.01fF
C17474 INVX1_LOC_328/Y INVX1_LOC_75/Y 0.09fF
C17475 VDD NAND2X1_LOC_516/Y 0.44fF
C17476 INVX1_LOC_257/Y INVX1_LOC_51/A 0.01fF
C17477 VDD INVX1_LOC_590/Y 0.26fF
C17478 INPUT_0 INVX1_LOC_228/Y 0.01fF
C17479 INVX1_LOC_317/Y NAND2X1_LOC_176/Y 0.01fF
C17480 NAND2X1_LOC_537/A INVX1_LOC_666/A 0.02fF
C17481 INVX1_LOC_414/A INVX1_LOC_413/Y 0.07fF
C17482 INVX1_LOC_107/A NAND2X1_LOC_114/a_36_24# 0.02fF
C17483 INVX1_LOC_41/Y NAND2X1_LOC_544/B 0.01fF
C17484 INPUT_0 INVX1_LOC_383/A 0.02fF
C17485 VDD INVX1_LOC_586/Y 0.21fF
C17486 INVX1_LOC_328/Y NAND2X1_LOC_271/A 0.02fF
C17487 INVX1_LOC_107/A NAND2X1_LOC_108/Y 0.01fF
C17488 NAND2X1_LOC_770/A INVX1_LOC_53/Y 0.01fF
C17489 INVX1_LOC_457/Y INVX1_LOC_577/Y -0.00fF
C17490 INVX1_LOC_420/Y INVX1_LOC_384/A 0.01fF
C17491 INVX1_LOC_578/A NAND2X1_LOC_568/a_36_24# 0.00fF
C17492 NAND2X1_LOC_29/a_36_24# INVX1_LOC_395/A 0.00fF
C17493 NAND2X1_LOC_516/Y INVX1_LOC_510/Y 0.07fF
C17494 INVX1_LOC_447/A INVX1_LOC_80/A 0.03fF
C17495 NAND2X1_LOC_97/B NAND2X1_LOC_76/B 0.01fF
C17496 VDD INVX1_LOC_515/Y 0.21fF
C17497 NAND2X1_LOC_331/A INVX1_LOC_196/A 0.06fF
C17498 NAND2X1_LOC_457/A INVX1_LOC_486/Y 0.01fF
C17499 NAND2X1_LOC_534/Y INVX1_LOC_21/Y 0.01fF
C17500 INVX1_LOC_288/A NAND2X1_LOC_173/Y 0.09fF
C17501 INVX1_LOC_145/Y INVX1_LOC_180/Y 0.04fF
C17502 VDD NAND2X1_LOC_123/A 0.06fF
C17503 NAND2X1_LOC_756/Y NAND2X1_LOC_506/B 0.01fF
C17504 VDD INVX1_LOC_607/Y 1.96fF
C17505 INVX1_LOC_53/Y INVX1_LOC_139/A 0.03fF
C17506 INVX1_LOC_395/A NAND2X1_LOC_307/A 0.02fF
C17507 NAND2X1_LOC_786/a_36_24# INVX1_LOC_366/A -0.00fF
C17508 NAND2X1_LOC_756/Y INVX1_LOC_45/Y 1.02fF
C17509 NAND2X1_LOC_383/Y INVX1_LOC_76/Y 0.13fF
C17510 INVX1_LOC_409/A INVX1_LOC_468/Y 0.01fF
C17511 INVX1_LOC_293/Y INVX1_LOC_45/Y 0.06fF
C17512 NAND2X1_LOC_750/Y INVX1_LOC_145/Y 0.06fF
C17513 NAND2X1_LOC_175/a_36_24# INVX1_LOC_577/Y 0.00fF
C17514 VDD INVX1_LOC_527/Y 0.39fF
C17515 INVX1_LOC_11/Y INVX1_LOC_447/A 0.04fF
C17516 NAND2X1_LOC_797/a_36_24# INVX1_LOC_6/Y 0.00fF
C17517 INVX1_LOC_420/Y INVX1_LOC_145/Y 0.06fF
C17518 INVX1_LOC_198/A INVX1_LOC_616/Y 0.02fF
C17519 INVX1_LOC_133/Y NAND2X1_LOC_814/Y 0.21fF
C17520 NAND2X1_LOC_539/a_36_24# INVX1_LOC_99/A 0.00fF
C17521 INVX1_LOC_286/Y INVX1_LOC_524/Y 0.00fF
C17522 INVX1_LOC_418/Y INVX1_LOC_206/Y 0.00fF
C17523 INVX1_LOC_206/Y INVX1_LOC_159/Y 0.87fF
C17524 VDD INVX1_LOC_362/A -0.00fF
C17525 VDD INVX1_LOC_498/A 0.12fF
C17526 NAND2X1_LOC_45/Y INVX1_LOC_50/Y 1.85fF
C17527 INVX1_LOC_375/A INVX1_LOC_98/Y 0.03fF
C17528 INVX1_LOC_276/A INVX1_LOC_53/Y 0.00fF
C17529 INVX1_LOC_407/Y INVX1_LOC_408/Y 0.02fF
C17530 INPUT_3 INVX1_LOC_293/Y 0.00fF
C17531 INVX1_LOC_617/Y INVX1_LOC_596/A 0.07fF
C17532 INPUT_0 NAND2X1_LOC_607/a_36_24# 0.00fF
C17533 INVX1_LOC_335/Y INVX1_LOC_113/Y 0.02fF
C17534 INVX1_LOC_20/Y NAND2X1_LOC_56/Y 0.02fF
C17535 NAND2X1_LOC_242/A NAND2X1_LOC_387/Y 0.01fF
C17536 INVX1_LOC_419/Y INVX1_LOC_395/A 0.07fF
C17537 GATE_579 INVX1_LOC_385/Y 0.07fF
C17538 INVX1_LOC_578/A INVX1_LOC_352/Y 0.09fF
C17539 VDD INVX1_LOC_83/A -0.00fF
C17540 INVX1_LOC_566/A INVX1_LOC_188/Y 0.06fF
C17541 VDD INVX1_LOC_476/Y 0.22fF
C17542 INVX1_LOC_166/A INVX1_LOC_118/Y 0.01fF
C17543 INPUT_0 INVX1_LOC_103/Y 0.01fF
C17544 VDD INVX1_LOC_283/Y 0.05fF
C17545 INVX1_LOC_372/Y INVX1_LOC_134/Y 0.03fF
C17546 NAND2X1_LOC_391/a_36_24# INVX1_LOC_230/A 0.01fF
C17547 INVX1_LOC_127/A INVX1_LOC_670/A 0.01fF
C17548 INVX1_LOC_45/Y NAND2X1_LOC_673/B 0.03fF
C17549 INVX1_LOC_156/Y INVX1_LOC_99/Y 0.01fF
C17550 INVX1_LOC_51/Y INVX1_LOC_137/Y 0.07fF
C17551 NAND2X1_LOC_498/Y INVX1_LOC_50/Y 0.07fF
C17552 INVX1_LOC_54/Y INVX1_LOC_255/Y 0.13fF
C17553 INVX1_LOC_570/A INVX1_LOC_50/Y 0.05fF
C17554 INVX1_LOC_554/Y INVX1_LOC_6/Y 0.01fF
C17555 INVX1_LOC_90/A INVX1_LOC_369/A 0.00fF
C17556 NAND2X1_LOC_114/a_36_24# NAND2X1_LOC_285/A 0.00fF
C17557 INVX1_LOC_384/A INVX1_LOC_371/A 0.01fF
C17558 INVX1_LOC_459/Y INVX1_LOC_345/Y 0.03fF
C17559 INVX1_LOC_17/Y INVX1_LOC_59/A 0.00fF
C17560 NAND2X1_LOC_108/Y NAND2X1_LOC_285/A 0.00fF
C17561 INVX1_LOC_608/Y INVX1_LOC_367/A 0.12fF
C17562 INVX1_LOC_587/Y INVX1_LOC_586/A 0.05fF
C17563 INVX1_LOC_114/Y INVX1_LOC_50/Y 0.15fF
C17564 INVX1_LOC_395/A NAND2X1_LOC_342/A 0.03fF
C17565 INVX1_LOC_648/Y INVX1_LOC_212/Y 0.01fF
C17566 NAND2X1_LOC_324/B NAND2X1_LOC_320/Y 0.17fF
C17567 INVX1_LOC_53/Y INVX1_LOC_7/Y 0.18fF
C17568 NAND2X1_LOC_362/a_36_24# INVX1_LOC_89/Y 0.01fF
C17569 INVX1_LOC_502/Y INPUT_1 0.87fF
C17570 INVX1_LOC_614/A INVX1_LOC_607/Y 0.48fF
C17571 NAND2X1_LOC_543/a_36_24# INVX1_LOC_98/Y 0.00fF
C17572 INVX1_LOC_224/Y NAND2X1_LOC_641/a_36_24# 0.00fF
C17573 NAND2X1_LOC_184/Y INVX1_LOC_651/Y 0.09fF
C17574 NAND2X1_LOC_130/Y NAND2X1_LOC_140/B 0.07fF
C17575 INVX1_LOC_418/Y INVX1_LOC_686/A 0.02fF
C17576 INVX1_LOC_625/A NAND2X1_LOC_97/B 0.31fF
C17577 INVX1_LOC_160/Y INVX1_LOC_154/A 0.00fF
C17578 INVX1_LOC_454/A INVX1_LOC_657/A 0.01fF
C17579 INVX1_LOC_291/A NAND2X1_LOC_333/B 0.36fF
C17580 INVX1_LOC_254/Y INVX1_LOC_318/Y 0.02fF
C17581 INVX1_LOC_377/Y INVX1_LOC_50/Y 0.13fF
C17582 NAND2X1_LOC_72/Y NAND2X1_LOC_72/a_36_24# 0.01fF
C17583 INVX1_LOC_210/Y INVX1_LOC_619/A 0.03fF
C17584 NAND2X1_LOC_311/a_36_24# INVX1_LOC_31/Y 0.01fF
C17585 INVX1_LOC_457/Y INVX1_LOC_26/Y 0.01fF
C17586 INPUT_0 NAND2X1_LOC_786/B 0.10fF
C17587 INVX1_LOC_448/A INVX1_LOC_371/A 0.07fF
C17588 INVX1_LOC_160/Y INVX1_LOC_501/A 0.08fF
C17589 INVX1_LOC_212/Y INVX1_LOC_242/A 0.03fF
C17590 INVX1_LOC_53/Y INVX1_LOC_345/Y 0.03fF
C17591 INVX1_LOC_442/Y INVX1_LOC_35/Y 0.07fF
C17592 INVX1_LOC_217/A INVX1_LOC_62/Y 0.01fF
C17593 INVX1_LOC_681/A NAND2X1_LOC_860/a_36_24# 0.02fF
C17594 INVX1_LOC_547/A INVX1_LOC_69/Y 0.37fF
C17595 NAND2X1_LOC_776/a_36_24# INVX1_LOC_26/Y 0.00fF
C17596 INVX1_LOC_18/Y INVX1_LOC_333/A 0.00fF
C17597 NAND2X1_LOC_307/A INVX1_LOC_31/Y 0.02fF
C17598 INVX1_LOC_53/Y INVX1_LOC_32/Y 0.06fF
C17599 INVX1_LOC_17/Y INVX1_LOC_400/A 0.07fF
C17600 INVX1_LOC_198/Y INVX1_LOC_600/Y 0.16fF
C17601 INVX1_LOC_154/Y INVX1_LOC_48/Y 0.18fF
C17602 INVX1_LOC_469/Y INVX1_LOC_188/Y 0.03fF
C17603 INVX1_LOC_224/Y INVX1_LOC_280/A 0.03fF
C17604 INVX1_LOC_220/Y NAND2X1_LOC_555/B 0.00fF
C17605 INVX1_LOC_17/Y INVX1_LOC_392/A 0.34fF
C17606 INVX1_LOC_468/Y INVX1_LOC_352/Y 0.74fF
C17607 NAND2X1_LOC_673/a_36_24# INVX1_LOC_48/Y 0.00fF
C17608 INVX1_LOC_586/A INVX1_LOC_9/Y 0.11fF
C17609 NAND2X1_LOC_673/B NAND2X1_LOC_69/Y 0.04fF
C17610 VDD INVX1_LOC_211/A 0.01fF
C17611 NAND2X1_LOC_332/B NAND2X1_LOC_768/B 0.23fF
C17612 INVX1_LOC_99/Y INVX1_LOC_50/Y 0.26fF
C17613 VDD INVX1_LOC_464/Y 0.21fF
C17614 VDD INVX1_LOC_64/Y 0.21fF
C17615 INVX1_LOC_17/Y NAND2X1_LOC_557/a_36_24# 0.00fF
C17616 NAND2X1_LOC_738/a_36_24# INVX1_LOC_6/Y 0.00fF
C17617 INVX1_LOC_21/Y INVX1_LOC_395/Y 0.01fF
C17618 NAND2X1_LOC_664/a_36_24# NAND2X1_LOC_333/B 0.00fF
C17619 INVX1_LOC_76/Y INVX1_LOC_662/A 0.03fF
C17620 INVX1_LOC_614/A INVX1_LOC_476/Y 0.05fF
C17621 INVX1_LOC_166/A NAND2X1_LOC_418/Y 0.01fF
C17622 INVX1_LOC_257/Y INVX1_LOC_441/A 0.02fF
C17623 INVX1_LOC_330/A INVX1_LOC_514/A 0.02fF
C17624 INVX1_LOC_206/Y NAND2X1_LOC_617/a_36_24# 0.00fF
C17625 INVX1_LOC_96/Y INVX1_LOC_531/Y 0.05fF
C17626 INVX1_LOC_17/Y INVX1_LOC_93/Y 0.36fF
C17627 INVX1_LOC_21/Y INVX1_LOC_89/Y 5.35fF
C17628 INVX1_LOC_53/Y NAND2X1_LOC_286/A 0.01fF
C17629 NAND2X1_LOC_400/B INVX1_LOC_7/Y 0.04fF
C17630 INVX1_LOC_11/Y INVX1_LOC_295/Y 0.03fF
C17631 INVX1_LOC_578/A NAND2X1_LOC_372/Y 0.09fF
C17632 INVX1_LOC_228/Y INVX1_LOC_211/A 0.07fF
C17633 INVX1_LOC_52/Y INVX1_LOC_625/Y 0.02fF
C17634 INVX1_LOC_435/A INVX1_LOC_230/Y 0.02fF
C17635 NAND2X1_LOC_543/B INVX1_LOC_92/A 1.51fF
C17636 INVX1_LOC_84/A INVX1_LOC_245/A 0.03fF
C17637 NAND2X1_LOC_566/a_36_24# INVX1_LOC_353/A 0.01fF
C17638 INVX1_LOC_312/Y INVX1_LOC_9/Y 0.07fF
C17639 INVX1_LOC_384/Y INVX1_LOC_244/Y 0.03fF
C17640 INVX1_LOC_345/Y INVX1_LOC_460/Y 0.17fF
C17641 NAND2X1_LOC_294/Y INVX1_LOC_453/Y 0.01fF
C17642 NAND2X1_LOC_180/B INVX1_LOC_79/A 0.02fF
C17643 INVX1_LOC_586/A INVX1_LOC_62/Y 0.20fF
C17644 INVX1_LOC_358/Y INVX1_LOC_501/A 0.02fF
C17645 INVX1_LOC_516/Y INVX1_LOC_62/Y 0.41fF
C17646 INVX1_LOC_288/A INVX1_LOC_354/A 0.04fF
C17647 INVX1_LOC_543/Y INVX1_LOC_86/Y 0.23fF
C17648 INVX1_LOC_335/Y INVX1_LOC_501/A 0.05fF
C17649 INVX1_LOC_199/Y NAND2X1_LOC_226/Y 0.07fF
C17650 INVX1_LOC_419/A NAND2X1_LOC_775/B 0.01fF
C17651 INVX1_LOC_665/Y INVX1_LOC_66/A 0.03fF
C17652 INVX1_LOC_53/Y INVX1_LOC_612/A 0.34fF
C17653 NAND2X1_LOC_740/a_36_24# INVX1_LOC_62/Y 0.00fF
C17654 INVX1_LOC_47/Y NAND2X1_LOC_465/a_36_24# 0.00fF
C17655 INVX1_LOC_17/Y INVX1_LOC_675/A 0.12fF
C17656 INVX1_LOC_201/Y INVX1_LOC_63/Y 0.34fF
C17657 INVX1_LOC_21/Y INVX1_LOC_179/Y 0.01fF
C17658 NAND2X1_LOC_24/Y INVX1_LOC_100/Y 0.04fF
C17659 INVX1_LOC_261/Y INVX1_LOC_673/Y 0.14fF
C17660 INVX1_LOC_188/Y INVX1_LOC_79/A 0.07fF
C17661 INVX1_LOC_47/Y INVX1_LOC_50/Y 0.77fF
C17662 INVX1_LOC_89/Y NAND2X1_LOC_267/A 0.07fF
C17663 NAND2X1_LOC_57/a_36_24# INVX1_LOC_223/Y 0.00fF
C17664 INVX1_LOC_35/Y INVX1_LOC_482/Y 0.07fF
C17665 GATE_865 INVX1_LOC_58/Y 0.03fF
C17666 NAND2X1_LOC_557/B INVX1_LOC_50/Y 0.01fF
C17667 INVX1_LOC_62/A INVX1_LOC_58/Y 0.01fF
C17668 INVX1_LOC_61/A INVX1_LOC_338/Y 0.04fF
C17669 NAND2X1_LOC_274/B NAND2X1_LOC_478/a_36_24# 0.00fF
C17670 INVX1_LOC_87/Y INVX1_LOC_6/Y 0.04fF
C17671 INVX1_LOC_312/Y INVX1_LOC_62/Y 0.07fF
C17672 INVX1_LOC_154/A NAND2X1_LOC_267/A 0.01fF
C17673 INVX1_LOC_335/A INVX1_LOC_498/Y 0.07fF
C17674 INPUT_5 INVX1_LOC_40/Y 0.01fF
C17675 INVX1_LOC_484/A NAND2X1_LOC_622/a_36_24# 0.02fF
C17676 INVX1_LOC_455/A NAND2X1_LOC_823/a_36_24# 0.00fF
C17677 NAND2X1_LOC_679/A NAND2X1_LOC_728/A 0.08fF
C17678 NAND2X1_LOC_148/a_36_24# INVX1_LOC_655/A 0.01fF
C17679 NAND2X1_LOC_308/A INVX1_LOC_66/A 0.07fF
C17680 INVX1_LOC_201/A NAND2X1_LOC_786/B 0.00fF
C17681 INVX1_LOC_479/A INVX1_LOC_318/Y 0.05fF
C17682 INVX1_LOC_543/Y INVX1_LOC_63/Y 0.03fF
C17683 INVX1_LOC_197/A INVX1_LOC_588/A 0.03fF
C17684 INVX1_LOC_17/Y NAND2X1_LOC_487/a_36_24# 0.00fF
C17685 INVX1_LOC_176/A NAND2X1_LOC_626/Y 0.14fF
C17686 INVX1_LOC_501/A NAND2X1_LOC_267/A 0.02fF
C17687 INVX1_LOC_376/A INVX1_LOC_31/Y 0.07fF
C17688 NAND2X1_LOC_545/A INVX1_LOC_349/Y 0.01fF
C17689 NAND2X1_LOC_532/Y INVX1_LOC_58/Y 0.04fF
C17690 INVX1_LOC_145/Y NAND2X1_LOC_488/Y 0.06fF
C17691 INVX1_LOC_54/Y INVX1_LOC_26/Y 0.40fF
C17692 INVX1_LOC_254/Y INVX1_LOC_90/Y 0.03fF
C17693 INVX1_LOC_119/Y INVX1_LOC_50/Y 2.49fF
C17694 INVX1_LOC_351/Y INVX1_LOC_361/A 0.12fF
C17695 INVX1_LOC_74/Y INVX1_LOC_504/Y 0.07fF
C17696 INVX1_LOC_41/Y INVX1_LOC_194/Y 0.01fF
C17697 NAND2X1_LOC_66/Y INVX1_LOC_50/Y 0.07fF
C17698 INVX1_LOC_31/Y INVX1_LOC_502/A 0.07fF
C17699 INVX1_LOC_202/Y INVX1_LOC_666/Y 1.07fF
C17700 INVX1_LOC_99/Y INVX1_LOC_658/Y 0.01fF
C17701 NAND2X1_LOC_274/B NAND2X1_LOC_542/A 0.03fF
C17702 NAND2X1_LOC_428/Y INVX1_LOC_505/A 0.16fF
C17703 INVX1_LOC_170/Y NAND2X1_LOC_626/Y 0.16fF
C17704 NAND2X1_LOC_274/B INVX1_LOC_376/Y 0.01fF
C17705 INVX1_LOC_520/Y INVX1_LOC_669/A 0.01fF
C17706 INVX1_LOC_44/Y INVX1_LOC_41/Y 0.12fF
C17707 INVX1_LOC_49/Y INVX1_LOC_653/Y 0.01fF
C17708 INVX1_LOC_636/A INVX1_LOC_259/Y 0.00fF
C17709 VDD INVX1_LOC_257/Y 0.97fF
C17710 NAND2X1_LOC_45/Y INVX1_LOC_438/A 0.10fF
C17711 INVX1_LOC_49/Y INVX1_LOC_666/Y 0.70fF
C17712 INVX1_LOC_63/Y INVX1_LOC_483/A 0.06fF
C17713 INVX1_LOC_62/Y INVX1_LOC_225/Y 0.01fF
C17714 NAND2X1_LOC_628/Y INVX1_LOC_487/A 0.17fF
C17715 INVX1_LOC_479/A INVX1_LOC_351/A 0.03fF
C17716 INVX1_LOC_369/Y NAND2X1_LOC_269/B 0.02fF
C17717 VDD INVX1_LOC_446/Y 0.96fF
C17718 INVX1_LOC_41/Y INVX1_LOC_461/Y 0.15fF
C17719 NAND2X1_LOC_637/A INVX1_LOC_580/Y 0.00fF
C17720 INVX1_LOC_479/A INVX1_LOC_90/Y 0.01fF
C17721 INVX1_LOC_203/Y INVX1_LOC_160/Y 0.06fF
C17722 INVX1_LOC_193/Y INVX1_LOC_560/A 0.02fF
C17723 NAND2X1_LOC_611/a_36_24# INVX1_LOC_92/A 0.00fF
C17724 NAND2X1_LOC_786/B INVX1_LOC_64/Y 0.03fF
C17725 INVX1_LOC_424/A NAND2X1_LOC_517/a_36_24# 0.00fF
C17726 INVX1_LOC_58/Y INVX1_LOC_76/A 0.01fF
C17727 INVX1_LOC_20/Y NAND2X1_LOC_75/a_36_24# 0.00fF
C17728 INVX1_LOC_655/A INVX1_LOC_240/Y 0.02fF
C17729 INVX1_LOC_99/Y INVX1_LOC_275/A 0.08fF
C17730 INVX1_LOC_320/Y INVX1_LOC_76/Y 0.02fF
C17731 NAND2X1_LOC_88/B NAND2X1_LOC_750/Y 0.03fF
C17732 VDD INVX1_LOC_9/A -0.00fF
C17733 VDD INVX1_LOC_613/Y 0.33fF
C17734 VDD INVX1_LOC_677/A -0.00fF
C17735 INVX1_LOC_607/A INVX1_LOC_651/Y 0.02fF
C17736 INVX1_LOC_426/A INVX1_LOC_416/A 0.02fF
C17737 VDD INVX1_LOC_145/Y 3.12fF
C17738 VDD NAND2X1_LOC_791/A -0.00fF
C17739 NAND2X1_LOC_93/Y INVX1_LOC_99/Y 0.12fF
C17740 INPUT_0 INVX1_LOC_619/A 0.03fF
C17741 VDD INVX1_LOC_661/Y 0.21fF
C17742 INVX1_LOC_438/A INVX1_LOC_99/Y 0.07fF
C17743 NAND2X1_LOC_543/B INPUT_1 0.02fF
C17744 INVX1_LOC_24/A INVX1_LOC_99/Y 0.02fF
C17745 NAND2X1_LOC_596/Y INVX1_LOC_145/Y 0.24fF
C17746 INVX1_LOC_438/Y INVX1_LOC_451/A 0.07fF
C17747 NAND2X1_LOC_249/Y INVX1_LOC_54/Y 0.08fF
C17748 INVX1_LOC_446/A NAND2X1_LOC_547/a_36_24# 0.00fF
C17749 INVX1_LOC_228/Y INVX1_LOC_145/Y 0.02fF
C17750 INVX1_LOC_206/Y INVX1_LOC_455/A 0.06fF
C17751 INVX1_LOC_17/Y INVX1_LOC_395/A 0.24fF
C17752 INVX1_LOC_166/A NAND2X1_LOC_533/a_36_24# 0.00fF
C17753 INVX1_LOC_417/A INVX1_LOC_65/Y 0.07fF
C17754 VDD INVX1_LOC_248/A -0.00fF
C17755 INVX1_LOC_412/A INVX1_LOC_35/Y 0.07fF
C17756 INVX1_LOC_574/A INVX1_LOC_575/Y 0.26fF
C17757 INVX1_LOC_448/A INVX1_LOC_383/A 0.01fF
C17758 INVX1_LOC_203/Y NAND2X1_LOC_267/A 0.01fF
C17759 INVX1_LOC_412/A INVX1_LOC_304/A 0.03fF
C17760 INVX1_LOC_266/A NAND2X1_LOC_307/A 0.07fF
C17761 INPUT_0 INVX1_LOC_105/A 0.03fF
C17762 VDD INVX1_LOC_433/A 0.00fF
C17763 NAND2X1_LOC_535/a_36_24# INVX1_LOC_31/Y 0.01fF
C17764 INVX1_LOC_266/A INVX1_LOC_545/Y -0.01fF
C17765 NAND2X1_LOC_566/a_36_24# INVX1_LOC_250/Y 0.00fF
C17766 INVX1_LOC_54/Y INVX1_LOC_560/A 0.07fF
C17767 NAND2X1_LOC_261/Y NAND2X1_LOC_260/Y 0.04fF
C17768 INVX1_LOC_492/A INVX1_LOC_521/Y 0.02fF
C17769 INVX1_LOC_17/Y INVX1_LOC_362/Y 0.09fF
C17770 INVX1_LOC_54/A INVX1_LOC_46/Y 0.01fF
C17771 NAND2X1_LOC_722/a_36_24# INVX1_LOC_565/A 0.02fF
C17772 NAND2X1_LOC_475/A INVX1_LOC_431/Y 0.00fF
C17773 VDD INVX1_LOC_141/Y 0.39fF
C17774 NAND2X1_LOC_516/Y INVX1_LOC_105/A 0.42fF
C17775 INVX1_LOC_238/Y INVX1_LOC_66/A 0.00fF
C17776 INVX1_LOC_381/A NAND2X1_LOC_297/a_36_24# 0.00fF
C17777 INVX1_LOC_400/Y INVX1_LOC_117/Y 0.07fF
C17778 NAND2X1_LOC_373/a_36_24# INVX1_LOC_257/A 0.00fF
C17779 INVX1_LOC_12/Y INVX1_LOC_318/Y 0.31fF
C17780 INVX1_LOC_567/A INVX1_LOC_9/Y 0.04fF
C17781 INVX1_LOC_444/Y INVX1_LOC_171/Y 0.03fF
C17782 NAND2X1_LOC_65/Y INVX1_LOC_177/A 0.11fF
C17783 INVX1_LOC_75/Y INVX1_LOC_109/Y 0.07fF
C17784 NAND2X1_LOC_332/B INVX1_LOC_371/A 0.03fF
C17785 INVX1_LOC_80/A NAND2X1_LOC_496/Y 0.34fF
C17786 INVX1_LOC_551/Y INVX1_LOC_230/A 0.11fF
C17787 INVX1_LOC_404/Y INVX1_LOC_69/Y 0.00fF
C17788 NAND2X1_LOC_331/A INVX1_LOC_69/Y 0.02fF
C17789 INVX1_LOC_131/Y INPUT_1 0.01fF
C17790 INVX1_LOC_395/A NAND2X1_LOC_307/B 0.07fF
C17791 INVX1_LOC_502/Y INVX1_LOC_50/Y 0.02fF
C17792 NAND2X1_LOC_180/B INVX1_LOC_48/Y 0.03fF
C17793 INVX1_LOC_137/A INVX1_LOC_555/A 0.14fF
C17794 INVX1_LOC_686/A INVX1_LOC_352/Y 0.07fF
C17795 NAND2X1_LOC_513/A INVX1_LOC_99/Y 0.73fF
C17796 INVX1_LOC_586/A INVX1_LOC_87/A 0.00fF
C17797 INVX1_LOC_224/Y INVX1_LOC_328/Y 0.04fF
C17798 NAND2X1_LOC_336/B INVX1_LOC_35/Y 0.31fF
C17799 INVX1_LOC_409/Y NAND2X1_LOC_123/B 0.23fF
C17800 INVX1_LOC_617/A INPUT_1 0.00fF
C17801 INVX1_LOC_21/Y INVX1_LOC_205/Y 0.01fF
C17802 NAND2X1_LOC_336/B INVX1_LOC_304/A 0.00fF
C17803 INVX1_LOC_364/Y INVX1_LOC_66/A 0.03fF
C17804 INVX1_LOC_118/Y INVX1_LOC_301/Y 0.00fF
C17805 INVX1_LOC_435/A NAND2X1_LOC_382/a_36_24# -0.01fF
C17806 NAND2X1_LOC_457/A NAND2X1_LOC_861/a_36_24# 0.00fF
C17807 INVX1_LOC_578/A INVX1_LOC_347/Y 0.09fF
C17808 INVX1_LOC_134/Y INVX1_LOC_159/A 0.05fF
C17809 INVX1_LOC_311/Y INVX1_LOC_48/Y 0.01fF
C17810 INVX1_LOC_603/Y INVX1_LOC_59/Y 0.02fF
C17811 INVX1_LOC_80/A NAND2X1_LOC_775/B 0.03fF
C17812 INVX1_LOC_206/Y NAND2X1_LOC_823/Y 0.18fF
C17813 INVX1_LOC_254/Y NAND2X1_LOC_545/B 0.00fF
C17814 INVX1_LOC_404/Y INVX1_LOC_247/Y 0.13fF
C17815 INVX1_LOC_255/Y INVX1_LOC_501/A 0.03fF
C17816 INVX1_LOC_11/Y NAND2X1_LOC_496/Y 0.02fF
C17817 INVX1_LOC_360/Y NAND2X1_LOC_123/A 0.17fF
C17818 INVX1_LOC_54/Y INVX1_LOC_369/A 0.05fF
C17819 INVX1_LOC_287/A INVX1_LOC_440/Y 0.01fF
C17820 INVX1_LOC_136/Y INVX1_LOC_50/Y 0.01fF
C17821 INVX1_LOC_315/Y INVX1_LOC_44/Y 0.03fF
C17822 INVX1_LOC_21/Y INVX1_LOC_194/Y 0.05fF
C17823 INVX1_LOC_278/A INVX1_LOC_100/Y 0.40fF
C17824 INVX1_LOC_53/A INVX1_LOC_25/Y 0.00fF
C17825 INVX1_LOC_603/Y INVX1_LOC_48/Y 0.01fF
C17826 INVX1_LOC_20/Y INVX1_LOC_187/Y 0.16fF
C17827 NAND2X1_LOC_317/a_36_24# INVX1_LOC_251/A 0.00fF
C17828 INVX1_LOC_670/A INVX1_LOC_519/A 0.03fF
C17829 INVX1_LOC_439/A NAND2X1_LOC_294/Y 0.01fF
C17830 NAND2X1_LOC_843/A INVX1_LOC_145/Y 0.46fF
C17831 NAND2X1_LOC_274/B INVX1_LOC_253/A 0.02fF
C17832 INVX1_LOC_266/A NAND2X1_LOC_325/a_36_24# -0.00fF
C17833 INVX1_LOC_118/Y INVX1_LOC_41/Y 0.03fF
C17834 INVX1_LOC_478/Y INVX1_LOC_59/Y 0.01fF
C17835 INVX1_LOC_366/A INVX1_LOC_9/Y 0.00fF
C17836 INVX1_LOC_20/Y NAND2X1_LOC_52/a_36_24# 0.00fF
C17837 INVX1_LOC_134/Y INVX1_LOC_66/A 0.17fF
C17838 NAND2X1_LOC_250/Y NAND2X1_LOC_106/B 0.00fF
C17839 INVX1_LOC_213/Y NAND2X1_LOC_259/A 0.02fF
C17840 INVX1_LOC_451/A INVX1_LOC_219/Y 0.02fF
C17841 INVX1_LOC_254/Y INVX1_LOC_98/Y 0.07fF
C17842 INVX1_LOC_25/Y INVX1_LOC_50/Y 0.01fF
C17843 INVX1_LOC_145/Y NAND2X1_LOC_243/A 0.01fF
C17844 INVX1_LOC_398/Y NAND2X1_LOC_387/Y 0.03fF
C17845 INVX1_LOC_103/Y INVX1_LOC_145/Y 0.03fF
C17846 NAND2X1_LOC_43/Y INVX1_LOC_50/Y 0.00fF
C17847 NAND2X1_LOC_692/Y INVX1_LOC_118/A 0.04fF
C17848 INVX1_LOC_204/Y INVX1_LOC_29/Y 0.00fF
C17849 INVX1_LOC_51/Y INVX1_LOC_502/A 0.02fF
C17850 INVX1_LOC_117/Y INVX1_LOC_125/A 0.01fF
C17851 INVX1_LOC_469/Y INVX1_LOC_504/Y 0.01fF
C17852 INVX1_LOC_197/A INVX1_LOC_63/Y 0.03fF
C17853 NAND2X1_LOC_791/B INVX1_LOC_285/Y 0.01fF
C17854 INVX1_LOC_17/Y INVX1_LOC_31/Y 0.39fF
C17855 INVX1_LOC_145/Y INVX1_LOC_68/A 0.01fF
C17856 INVX1_LOC_545/A INVX1_LOC_93/Y 0.01fF
C17857 NAND2X1_LOC_335/B INVX1_LOC_270/Y 0.01fF
C17858 INVX1_LOC_93/Y INVX1_LOC_108/Y 0.01fF
C17859 GATE_865 NAND2X1_LOC_866/a_36_24# 0.02fF
C17860 INVX1_LOC_84/A NAND2X1_LOC_126/a_36_24# 0.00fF
C17861 NAND2X1_LOC_387/Y INVX1_LOC_48/Y 0.15fF
C17862 NAND2X1_LOC_820/A INVX1_LOC_9/Y 0.02fF
C17863 NAND2X1_LOC_498/B INVX1_LOC_653/Y 0.29fF
C17864 INVX1_LOC_300/A INVX1_LOC_187/Y 0.02fF
C17865 INVX1_LOC_391/Y INVX1_LOC_387/Y 1.26fF
C17866 INVX1_LOC_21/Y INVX1_LOC_44/Y 0.10fF
C17867 INVX1_LOC_46/Y NAND2X1_LOC_84/B 0.02fF
C17868 NAND2X1_LOC_335/B INVX1_LOC_92/A 0.01fF
C17869 INVX1_LOC_63/Y NAND2X1_LOC_416/Y 0.03fF
C17870 INVX1_LOC_93/Y INVX1_LOC_189/A 0.01fF
C17871 INVX1_LOC_31/Y NAND2X1_LOC_435/a_36_24# 0.00fF
C17872 INVX1_LOC_76/Y INVX1_LOC_653/Y 0.07fF
C17873 INVX1_LOC_236/A INVX1_LOC_508/A 0.02fF
C17874 NAND2X1_LOC_542/A INVX1_LOC_159/Y 0.00fF
C17875 INVX1_LOC_587/Y INVX1_LOC_6/Y 0.03fF
C17876 INVX1_LOC_100/Y NAND2X1_LOC_601/a_36_24# 0.01fF
C17877 INVX1_LOC_76/Y INVX1_LOC_666/Y 0.02fF
C17878 INVX1_LOC_35/Y NAND2X1_LOC_847/A 0.02fF
C17879 INVX1_LOC_63/Y NAND2X1_LOC_106/B 0.05fF
C17880 INVX1_LOC_17/Y INVX1_LOC_682/Y 0.19fF
C17881 INVX1_LOC_100/A INVX1_LOC_46/Y 0.83fF
C17882 INVX1_LOC_96/A INVX1_LOC_50/Y 0.12fF
C17883 INVX1_LOC_12/Y INVX1_LOC_90/Y 0.56fF
C17884 INVX1_LOC_273/A NAND2X1_LOC_227/A 0.01fF
C17885 INVX1_LOC_431/A INVX1_LOC_49/Y 0.02fF
C17886 INVX1_LOC_62/Y INVX1_LOC_486/Y 0.17fF
C17887 INVX1_LOC_492/A NAND2X1_LOC_846/B 0.00fF
C17888 INVX1_LOC_188/Y INVX1_LOC_472/Y 0.01fF
C17889 INVX1_LOC_413/A INVX1_LOC_58/Y 0.01fF
C17890 INVX1_LOC_63/A INVX1_LOC_621/A 0.00fF
C17891 INVX1_LOC_145/Y NAND2X1_LOC_786/B 0.10fF
C17892 INVX1_LOC_556/Y INVX1_LOC_124/A 0.01fF
C17893 INVX1_LOC_17/Y NAND2X1_LOC_488/a_36_24# 0.00fF
C17894 NAND2X1_LOC_403/A INVX1_LOC_100/Y 0.01fF
C17895 NAND2X1_LOC_698/Y INVX1_LOC_32/Y 0.04fF
C17896 INVX1_LOC_20/Y NAND2X1_LOC_832/A 0.05fF
C17897 NAND2X1_LOC_545/B INVX1_LOC_479/A 0.04fF
C17898 INVX1_LOC_369/A INVX1_LOC_388/A 0.12fF
C17899 NAND2X1_LOC_346/B NAND2X1_LOC_295/a_36_24# 0.02fF
C17900 INVX1_LOC_173/Y INVX1_LOC_63/Y 0.00fF
C17901 INVX1_LOC_100/Y INVX1_LOC_453/Y 0.03fF
C17902 INVX1_LOC_491/A INVX1_LOC_48/Y 0.07fF
C17903 INVX1_LOC_21/Y INVX1_LOC_347/A 0.07fF
C17904 INVX1_LOC_543/A INVX1_LOC_198/A 0.09fF
C17905 INVX1_LOC_525/Y INVX1_LOC_95/A 0.02fF
C17906 INVX1_LOC_41/Y INVX1_LOC_365/A 0.02fF
C17907 NAND2X1_LOC_409/Y INVX1_LOC_1/Y 1.07fF
C17908 INVX1_LOC_179/A NAND2X1_LOC_203/a_36_24# 0.03fF
C17909 INVX1_LOC_145/Y INVX1_LOC_635/Y 0.02fF
C17910 INVX1_LOC_54/Y NAND2X1_LOC_626/Y 0.12fF
C17911 INVX1_LOC_551/A INVX1_LOC_199/Y 0.02fF
C17912 INVX1_LOC_6/Y INVX1_LOC_9/Y 0.17fF
C17913 INVX1_LOC_442/Y INVX1_LOC_364/A 0.01fF
C17914 INVX1_LOC_479/A INVX1_LOC_98/Y 0.38fF
C17915 INVX1_LOC_59/Y INVX1_LOC_91/A 0.01fF
C17916 NAND2X1_LOC_854/a_36_24# INVX1_LOC_347/Y 0.00fF
C17917 INVX1_LOC_662/A NAND2X1_LOC_815/a_36_24# 0.01fF
C17918 INVX1_LOC_89/Y INVX1_LOC_128/Y 0.03fF
C17919 INVX1_LOC_89/Y INVX1_LOC_26/Y 0.06fF
C17920 INVX1_LOC_74/Y INVX1_LOC_259/Y 0.03fF
C17921 INVX1_LOC_662/A NAND2X1_LOC_286/A 0.02fF
C17922 INVX1_LOC_69/Y NAND2X1_LOC_833/B 0.02fF
C17923 INVX1_LOC_49/Y NAND2X1_LOC_489/A 0.03fF
C17924 INVX1_LOC_170/A INVX1_LOC_90/Y 0.01fF
C17925 INVX1_LOC_501/A INVX1_LOC_26/Y 0.03fF
C17926 INVX1_LOC_62/Y INVX1_LOC_6/Y 0.10fF
C17927 NAND2X1_LOC_81/Y INVX1_LOC_9/Y 0.01fF
C17928 INVX1_LOC_179/Y INVX1_LOC_26/Y 0.03fF
C17929 INVX1_LOC_6/Y NAND2X1_LOC_844/A 0.04fF
C17930 INPUT_0 NAND2X1_LOC_61/A 0.01fF
C17931 INVX1_LOC_148/Y INVX1_LOC_139/Y 0.17fF
C17932 INVX1_LOC_479/A INVX1_LOC_338/Y 0.03fF
C17933 VDD NAND2X1_LOC_331/B 0.03fF
C17934 INVX1_LOC_468/A INVX1_LOC_376/Y 0.12fF
C17935 NAND2X1_LOC_88/Y INVX1_LOC_395/A 0.05fF
C17936 INVX1_LOC_447/A INVX1_LOC_393/Y 0.18fF
C17937 INVX1_LOC_74/Y INVX1_LOC_114/A 0.08fF
C17938 INVX1_LOC_557/A NAND2X1_LOC_317/A 0.15fF
C17939 NAND2X1_LOC_843/B NAND2X1_LOC_278/a_36_24# 0.02fF
C17940 VDD NAND2X1_LOC_332/B 0.22fF
C17941 INPUT_0 INVX1_LOC_45/Y 0.26fF
C17942 INVX1_LOC_404/Y INVX1_LOC_586/A 0.18fF
C17943 NAND2X1_LOC_331/A INVX1_LOC_586/A 0.02fF
C17944 VDD INVX1_LOC_125/Y 0.22fF
C17945 INVX1_LOC_20/Y NAND2X1_LOC_750/Y 0.03fF
C17946 INVX1_LOC_239/Y INVX1_LOC_80/A 0.01fF
C17947 INVX1_LOC_394/Y INVX1_LOC_21/Y 0.01fF
C17948 NAND2X1_LOC_88/B VDD 0.00fF
C17949 INVX1_LOC_590/Y INVX1_LOC_45/Y 0.01fF
C17950 NAND2X1_LOC_788/A INVX1_LOC_134/Y 0.04fF
C17951 VDD NAND2X1_LOC_460/A -0.00fF
C17952 INPUT_0 INPUT_3 0.03fF
C17953 NAND2X1_LOC_475/A INVX1_LOC_187/A 0.18fF
C17954 NAND2X1_LOC_16/Y INVX1_LOC_76/Y 0.01fF
C17955 VDD NAND2X1_LOC_260/Y 0.01fF
C17956 NAND2X1_LOC_669/Y INVX1_LOC_206/Y 0.03fF
C17957 INVX1_LOC_492/A INVX1_LOC_554/A 0.02fF
C17958 INVX1_LOC_566/A NAND2X1_LOC_327/a_36_24# 0.00fF
C17959 INVX1_LOC_408/Y INVX1_LOC_134/Y 0.08fF
C17960 INVX1_LOC_434/A INVX1_LOC_442/Y 0.19fF
C17961 VDD INVX1_LOC_503/Y 0.28fF
C17962 INVX1_LOC_259/Y NAND2X1_LOC_591/B 0.02fF
C17963 INVX1_LOC_395/A NAND2X1_LOC_616/Y 0.07fF
C17964 INVX1_LOC_21/Y INVX1_LOC_118/Y 0.42fF
C17965 VDD INVX1_LOC_440/A -0.00fF
C17966 INVX1_LOC_374/A INVX1_LOC_197/A 0.03fF
C17967 INVX1_LOC_20/Y NAND2X1_LOC_173/Y 0.03fF
C17968 INVX1_LOC_442/A INVX1_LOC_134/Y 0.03fF
C17969 INVX1_LOC_381/A INVX1_LOC_378/A 0.03fF
C17970 INVX1_LOC_222/Y INVX1_LOC_283/A 0.02fF
C17971 NAND2X1_LOC_249/Y INVX1_LOC_277/A 0.00fF
C17972 NAND2X1_LOC_322/Y INPUT_1 0.11fF
C17973 INVX1_LOC_257/Y INVX1_LOC_360/Y 0.16fF
C17974 INVX1_LOC_142/Y INVX1_LOC_522/Y 0.05fF
C17975 INVX1_LOC_436/A INVX1_LOC_384/Y 0.09fF
C17976 NAND2X1_LOC_164/Y NAND2X1_LOC_164/a_36_24# 0.02fF
C17977 NAND2X1_LOC_241/B INVX1_LOC_197/Y 0.12fF
C17978 NAND2X1_LOC_340/a_36_24# INVX1_LOC_395/A 0.00fF
C17979 INVX1_LOC_98/A INVX1_LOC_97/Y 0.00fF
C17980 NAND2X1_LOC_331/A INVX1_LOC_330/A 0.00fF
C17981 INVX1_LOC_569/A NAND2X1_LOC_726/a_36_24# 0.02fF
C17982 INVX1_LOC_11/Y NAND2X1_LOC_317/B 0.15fF
C17983 INVX1_LOC_629/A INVX1_LOC_259/Y 0.00fF
C17984 INVX1_LOC_434/A INVX1_LOC_671/A 0.14fF
C17985 INVX1_LOC_35/Y INVX1_LOC_215/Y 0.01fF
C17986 INVX1_LOC_69/Y INVX1_LOC_638/A 0.08fF
C17987 INVX1_LOC_400/Y NAND2X1_LOC_143/a_36_24# 0.01fF
C17988 NAND2X1_LOC_45/Y INVX1_LOC_117/Y 0.07fF
C17989 INVX1_LOC_206/Y INVX1_LOC_186/Y 0.03fF
C17990 INVX1_LOC_607/Y INVX1_LOC_45/Y 0.09fF
C17991 VDD NAND2X1_LOC_128/B 0.10fF
C17992 GATE_741 INVX1_LOC_186/A 0.02fF
C17993 INVX1_LOC_238/A INVX1_LOC_89/Y 0.01fF
C17994 INVX1_LOC_17/Y INVX1_LOC_51/Y 0.17fF
C17995 INVX1_LOC_288/A INVX1_LOC_360/Y 0.02fF
C17996 INVX1_LOC_364/Y INVX1_LOC_116/Y 0.37fF
C17997 INVX1_LOC_395/A INVX1_LOC_189/A 0.05fF
C17998 INVX1_LOC_42/Y INVX1_LOC_366/A 0.11fF
C17999 NAND2X1_LOC_231/A INVX1_LOC_35/Y 0.01fF
C18000 INVX1_LOC_20/Y NAND2X1_LOC_413/Y 0.04fF
C18001 INVX1_LOC_551/Y NAND2X1_LOC_72/Y 0.02fF
C18002 INVX1_LOC_80/A INVX1_LOC_633/Y 0.02fF
C18003 NAND2X1_LOC_498/Y INVX1_LOC_117/Y 0.44fF
C18004 INVX1_LOC_686/A INVX1_LOC_67/Y 0.03fF
C18005 INVX1_LOC_269/A INVX1_LOC_48/Y 0.46fF
C18006 INVX1_LOC_425/Y INVX1_LOC_586/A 0.01fF
C18007 INVX1_LOC_395/A INVX1_LOC_230/Y 0.18fF
C18008 INVX1_LOC_570/A INVX1_LOC_117/Y 0.07fF
C18009 NAND2X1_LOC_592/B INVX1_LOC_31/Y 0.01fF
C18010 INVX1_LOC_266/A INVX1_LOC_17/Y 0.07fF
C18011 INVX1_LOC_11/Y NAND2X1_LOC_613/Y -0.00fF
C18012 INVX1_LOC_270/A INVX1_LOC_230/A 0.23fF
C18013 INVX1_LOC_560/A INVX1_LOC_89/Y 0.69fF
C18014 INVX1_LOC_93/Y INVX1_LOC_249/Y 0.22fF
C18015 INVX1_LOC_29/A INVX1_LOC_55/Y 0.00fF
C18016 INVX1_LOC_298/A INVX1_LOC_45/Y 0.01fF
C18017 INVX1_LOC_11/Y INVX1_LOC_169/A 0.04fF
C18018 INVX1_LOC_45/Y INVX1_LOC_498/A 0.03fF
C18019 INVX1_LOC_20/Y INVX1_LOC_371/A 0.15fF
C18020 INVX1_LOC_206/Y INVX1_LOC_347/Y 0.02fF
C18021 INVX1_LOC_409/A INVX1_LOC_376/Y 0.15fF
C18022 NAND2X1_LOC_755/B INVX1_LOC_635/A 0.10fF
C18023 VDD INVX1_LOC_484/Y 0.21fF
C18024 INVX1_LOC_93/Y NAND2X1_LOC_122/Y 0.05fF
C18025 INVX1_LOC_103/Y NAND2X1_LOC_332/B 0.15fF
C18026 INVX1_LOC_566/A INVX1_LOC_259/Y 0.01fF
C18027 VDD INVX1_LOC_242/Y 2.13fF
C18028 INVX1_LOC_134/Y INVX1_LOC_116/Y 0.01fF
C18029 INVX1_LOC_617/A INVX1_LOC_50/Y 0.00fF
C18030 INVX1_LOC_206/Y INVX1_LOC_328/Y 3.65fF
C18031 INVX1_LOC_619/A INVX1_LOC_145/Y 0.10fF
C18032 INVX1_LOC_439/Y INVX1_LOC_424/Y 0.03fF
C18033 INVX1_LOC_54/Y INVX1_LOC_235/Y 0.10fF
C18034 INVX1_LOC_145/Y NAND2X1_LOC_486/a_36_24# 0.01fF
C18035 INVX1_LOC_21/Y NAND2X1_LOC_418/Y 0.01fF
C18036 INVX1_LOC_400/Y INVX1_LOC_58/Y 0.13fF
C18037 INVX1_LOC_435/A NAND2X1_LOC_363/a_36_24# 0.00fF
C18038 INVX1_LOC_224/Y INVX1_LOC_224/A 0.01fF
C18039 INVX1_LOC_99/A NAND2X1_LOC_102/a_36_24# 0.02fF
C18040 INVX1_LOC_206/Y INVX1_LOC_518/A 0.02fF
C18041 INVX1_LOC_442/A INVX1_LOC_65/A 0.05fF
C18042 INVX1_LOC_5/Y INPUT_4 0.15fF
C18043 INVX1_LOC_11/Y INVX1_LOC_633/Y 0.07fF
C18044 NAND2X1_LOC_307/B INVX1_LOC_51/Y 0.07fF
C18045 INVX1_LOC_318/Y NAND2X1_LOC_615/B 0.01fF
C18046 INVX1_LOC_167/A INVX1_LOC_492/Y 0.02fF
C18047 INVX1_LOC_376/A INVX1_LOC_355/A 0.06fF
C18048 INVX1_LOC_218/A INVX1_LOC_6/Y 0.33fF
C18049 INVX1_LOC_21/Y INVX1_LOC_365/A 0.01fF
C18050 INVX1_LOC_134/Y NAND2X1_LOC_432/Y 0.05fF
C18051 INVX1_LOC_468/Y INVX1_LOC_352/A 0.00fF
C18052 NAND2X1_LOC_843/A NAND2X1_LOC_260/Y 0.00fF
C18053 NAND2X1_LOC_427/Y NAND2X1_LOC_427/a_36_24# 0.02fF
C18054 NAND2X1_LOC_457/A INVX1_LOC_100/Y 0.00fF
C18055 NAND2X1_LOC_184/Y INVX1_LOC_53/Y 0.10fF
C18056 NAND2X1_LOC_523/B NAND2X1_LOC_521/Y 0.01fF
C18057 INVX1_LOC_425/A INVX1_LOC_411/Y 0.01fF
C18058 INPUT_3 INVX1_LOC_83/A -0.02fF
C18059 INVX1_LOC_628/A INVX1_LOC_259/Y 0.00fF
C18060 INVX1_LOC_448/A INVX1_LOC_105/A 0.06fF
C18061 NAND2X1_LOC_503/Y INVX1_LOC_97/Y 0.05fF
C18062 NAND2X1_LOC_130/Y INPUT_1 0.03fF
C18063 INVX1_LOC_47/Y INVX1_LOC_111/A 0.04fF
C18064 INVX1_LOC_31/Y NAND2X1_LOC_616/Y 0.54fF
C18065 INVX1_LOC_117/Y INVX1_LOC_99/Y 0.39fF
C18066 NAND2X1_LOC_719/a_36_24# INVX1_LOC_74/Y 0.01fF
C18067 INVX1_LOC_436/A NAND2X1_LOC_555/B 0.01fF
C18068 INVX1_LOC_686/A INVX1_LOC_347/Y 0.09fF
C18069 INVX1_LOC_17/Y INVX1_LOC_254/A 0.03fF
C18070 INVX1_LOC_518/A INVX1_LOC_242/A 4.35fF
C18071 INVX1_LOC_189/Y INVX1_LOC_189/A 0.16fF
C18072 NAND2X1_LOC_708/A NAND2X1_LOC_696/a_36_24# 0.02fF
C18073 INVX1_LOC_468/A INVX1_LOC_253/A 0.17fF
C18074 INVX1_LOC_54/Y INVX1_LOC_81/Y 0.00fF
C18075 INVX1_LOC_46/Y INVX1_LOC_230/A 0.07fF
C18076 INVX1_LOC_612/Y NAND2X1_LOC_708/A 0.00fF
C18077 INVX1_LOC_255/Y INVX1_LOC_347/A 0.01fF
C18078 NAND2X1_LOC_97/B INVX1_LOC_63/Y 0.01fF
C18079 INVX1_LOC_435/Y INVX1_LOC_479/A 0.10fF
C18080 INVX1_LOC_203/A INVX1_LOC_94/A 0.06fF
C18081 NAND2X1_LOC_387/Y INVX1_LOC_396/A 0.01fF
C18082 INVX1_LOC_581/Y INVX1_LOC_137/Y 0.02fF
C18083 INVX1_LOC_537/A INVX1_LOC_58/Y 0.46fF
C18084 NAND2X1_LOC_259/A NAND2X1_LOC_258/Y 0.00fF
C18085 INVX1_LOC_624/Y INVX1_LOC_252/A 0.00fF
C18086 INVX1_LOC_65/A INVX1_LOC_116/Y 0.01fF
C18087 NAND2X1_LOC_433/Y INVX1_LOC_633/Y 0.07fF
C18088 INVX1_LOC_69/Y INVX1_LOC_685/Y 0.03fF
C18089 INVX1_LOC_399/A INVX1_LOC_600/A 0.01fF
C18090 INVX1_LOC_45/Y INVX1_LOC_211/A 0.04fF
C18091 INVX1_LOC_100/Y INVX1_LOC_651/A 0.00fF
C18092 INVX1_LOC_123/A INVX1_LOC_117/Y 0.03fF
C18093 INVX1_LOC_89/Y INVX1_LOC_603/A 0.06fF
C18094 INVX1_LOC_492/A INVX1_LOC_199/Y 0.06fF
C18095 INVX1_LOC_45/Y INVX1_LOC_464/Y 0.04fF
C18096 INVX1_LOC_561/A INVX1_LOC_32/Y 0.03fF
C18097 INVX1_LOC_355/Y INVX1_LOC_359/A 0.01fF
C18098 GATE_865 INVX1_LOC_639/A 0.15fF
C18099 INVX1_LOC_678/A INVX1_LOC_674/Y 0.03fF
C18100 NAND2X1_LOC_482/Y NAND2X1_LOC_252/Y 0.01fF
C18101 INVX1_LOC_205/Y INVX1_LOC_26/Y 0.03fF
C18102 INVX1_LOC_117/Y INVX1_LOC_47/Y 0.24fF
C18103 INVX1_LOC_6/Y INVX1_LOC_87/A 0.06fF
C18104 NAND2X1_LOC_148/B INVX1_LOC_132/A -0.00fF
C18105 NAND2X1_LOC_635/a_36_24# INVX1_LOC_74/Y 0.00fF
C18106 INVX1_LOC_352/Y INVX1_LOC_376/Y 0.03fF
C18107 INVX1_LOC_596/A INVX1_LOC_479/A 0.01fF
C18108 INVX1_LOC_42/Y NAND2X1_LOC_81/Y -0.00fF
C18109 INVX1_LOC_158/Y INVX1_LOC_242/Y 0.04fF
C18110 INVX1_LOC_167/A INVX1_LOC_168/Y 0.15fF
C18111 INVX1_LOC_53/Y INVX1_LOC_75/Y 0.08fF
C18112 INVX1_LOC_406/A NAND2X1_LOC_523/a_36_24# 0.02fF
C18113 NAND2X1_LOC_615/B INVX1_LOC_351/A 0.03fF
C18114 INVX1_LOC_58/Y INVX1_LOC_496/Y 0.06fF
C18115 INVX1_LOC_100/A INVX1_LOC_49/Y 0.23fF
C18116 NAND2X1_LOC_128/A INVX1_LOC_63/Y 0.01fF
C18117 INVX1_LOC_161/A INVX1_LOC_62/Y 0.03fF
C18118 INVX1_LOC_26/Y INVX1_LOC_194/Y 0.03fF
C18119 INVX1_LOC_504/A NAND2X1_LOC_118/a_36_24# 0.01fF
C18120 INVX1_LOC_50/Y INVX1_LOC_353/A 0.06fF
C18121 INVX1_LOC_41/Y INVX1_LOC_252/Y 0.06fF
C18122 INVX1_LOC_79/A INVX1_LOC_259/Y 0.03fF
C18123 INVX1_LOC_255/A INVX1_LOC_65/A 0.08fF
C18124 NAND2X1_LOC_615/B INVX1_LOC_90/Y 0.03fF
C18125 NAND2X1_LOC_502/a_36_24# INVX1_LOC_615/A 0.00fF
C18126 INVX1_LOC_7/Y INVX1_LOC_327/A 0.05fF
C18127 INVX1_LOC_117/Y INVX1_LOC_119/Y 3.56fF
C18128 INVX1_LOC_117/Y NAND2X1_LOC_66/Y 0.03fF
C18129 INVX1_LOC_469/Y INVX1_LOC_114/A 2.77fF
C18130 INVX1_LOC_89/Y NAND2X1_LOC_605/B 0.02fF
C18131 INVX1_LOC_224/Y INVX1_LOC_109/Y 0.67fF
C18132 INVX1_LOC_32/Y NAND2X1_LOC_545/A 0.06fF
C18133 INVX1_LOC_75/A INVX1_LOC_230/A 0.13fF
C18134 INVX1_LOC_53/Y NAND2X1_LOC_271/A 0.19fF
C18135 NAND2X1_LOC_184/Y NAND2X1_LOC_844/a_36_24# 0.00fF
C18136 INVX1_LOC_578/A INVX1_LOC_109/Y 0.07fF
C18137 INVX1_LOC_504/A NAND2X1_LOC_468/a_36_24# 0.00fF
C18138 NAND2X1_LOC_7/Y VDD -0.00fF
C18139 NAND2X1_LOC_689/B NAND2X1_LOC_691/A 0.01fF
C18140 INVX1_LOC_644/Y NAND2X1_LOC_846/B 0.04fF
C18141 INVX1_LOC_44/Y INVX1_LOC_26/Y 0.13fF
C18142 VDD INVX1_LOC_301/A 0.15fF
C18143 NAND2X1_LOC_503/B INVX1_LOC_395/A 0.32fF
C18144 VDD INVX1_LOC_626/Y 0.21fF
C18145 NAND2X1_LOC_283/a_36_24# NAND2X1_LOC_843/B 0.00fF
C18146 INVX1_LOC_63/Y NAND2X1_LOC_248/B 0.00fF
C18147 NAND2X1_LOC_274/B INVX1_LOC_652/A 0.57fF
C18148 NAND2X1_LOC_192/A INVX1_LOC_62/Y 0.38fF
C18149 INVX1_LOC_79/A INVX1_LOC_114/A 0.11fF
C18150 INVX1_LOC_448/Y NAND2X1_LOC_498/Y 0.03fF
C18151 VDD INVX1_LOC_533/Y 0.47fF
C18152 NAND2X1_LOC_331/A INVX1_LOC_140/Y 0.00fF
C18153 VDD INVX1_LOC_132/Y 0.21fF
C18154 INVX1_LOC_153/Y NAND2X1_LOC_231/B 0.02fF
C18155 INVX1_LOC_257/Y INVX1_LOC_45/Y 0.07fF
C18156 INVX1_LOC_206/Y INVX1_LOC_266/Y 0.03fF
C18157 INVX1_LOC_20/Y VDD 1.69fF
C18158 INVX1_LOC_177/Y INVX1_LOC_182/A 0.02fF
C18159 NAND2X1_LOC_711/a_36_24# INVX1_LOC_367/A 0.00fF
C18160 INVX1_LOC_239/Y INVX1_LOC_131/A 0.10fF
C18161 VDD INVX1_LOC_175/Y 0.21fF
C18162 INVX1_LOC_446/Y INVX1_LOC_45/Y 0.07fF
C18163 INVX1_LOC_626/A INVX1_LOC_133/Y 0.01fF
C18164 INVX1_LOC_395/A INVX1_LOC_273/A 0.05fF
C18165 NAND2X1_LOC_808/a_36_24# INVX1_LOC_638/A 0.00fF
C18166 INVX1_LOC_405/A NAND2X1_LOC_416/Y 0.00fF
C18167 INVX1_LOC_20/Y INVX1_LOC_228/Y -0.00fF
C18168 INVX1_LOC_568/Y INVX1_LOC_554/A 0.34fF
C18169 NAND2X1_LOC_61/A INVX1_LOC_145/Y 0.01fF
C18170 NAND2X1_LOC_65/Y INVX1_LOC_65/Y 0.01fF
C18171 INVX1_LOC_223/A NAND2X1_LOC_263/a_36_24# 0.00fF
C18172 INVX1_LOC_384/A INVX1_LOC_45/Y 0.07fF
C18173 INVX1_LOC_62/Y INVX1_LOC_636/A 0.07fF
C18174 NAND2X1_LOC_503/Y INVX1_LOC_615/A 0.05fF
C18175 INVX1_LOC_17/Y NAND2X1_LOC_537/A 0.03fF
C18176 INVX1_LOC_590/Y NAND2X1_LOC_756/Y 0.23fF
C18177 INVX1_LOC_447/A INVX1_LOC_442/Y 0.01fF
C18178 VDD INVX1_LOC_197/Y 0.49fF
C18179 INVX1_LOC_195/A INVX1_LOC_7/Y 0.01fF
C18180 INVX1_LOC_317/Y NAND2X1_LOC_388/a_36_24# 0.00fF
C18181 INVX1_LOC_20/Y INVX1_LOC_510/Y 0.12fF
C18182 NAND2X1_LOC_750/Y NAND2X1_LOC_61/a_36_24# 0.00fF
C18183 INVX1_LOC_191/A INVX1_LOC_366/A 0.03fF
C18184 NAND2X1_LOC_231/A INVX1_LOC_291/A 0.16fF
C18185 INVX1_LOC_120/Y INVX1_LOC_109/Y 0.01fF
C18186 NAND2X1_LOC_209/a_36_24# INVX1_LOC_575/Y 0.00fF
C18187 NAND2X1_LOC_543/a_36_24# INVX1_LOC_65/Y 0.01fF
C18188 NAND2X1_LOC_271/B INVX1_LOC_367/Y 0.03fF
C18189 INVX1_LOC_607/A INVX1_LOC_53/Y 0.01fF
C18190 INVX1_LOC_278/A NAND2X1_LOC_261/a_36_24# 0.00fF
C18191 VDD INVX1_LOC_663/Y 0.21fF
C18192 NAND2X1_LOC_322/Y INVX1_LOC_50/Y 0.00fF
C18193 INVX1_LOC_301/A INVX1_LOC_103/Y 0.00fF
C18194 INVX1_LOC_228/Y INVX1_LOC_300/A 0.01fF
C18195 INVX1_LOC_185/Y NAND2X1_LOC_612/A 0.01fF
C18196 NAND2X1_LOC_486/B INVX1_LOC_53/Y 0.09fF
C18197 INVX1_LOC_206/Y INVX1_LOC_172/A 0.02fF
C18198 NAND2X1_LOC_543/B NAND2X1_LOC_388/A 0.27fF
C18199 INVX1_LOC_459/A INVX1_LOC_49/Y 0.01fF
C18200 NAND2X1_LOC_475/A INVX1_LOC_117/Y 0.12fF
C18201 NAND2X1_LOC_45/Y INVX1_LOC_608/A 0.07fF
C18202 INVX1_LOC_268/Y INVX1_LOC_635/A 0.00fF
C18203 INVX1_LOC_206/Y INVX1_LOC_105/Y 1.05fF
C18204 INVX1_LOC_284/A INVX1_LOC_273/A 0.25fF
C18205 INVX1_LOC_45/Y INVX1_LOC_145/Y 0.42fF
C18206 INVX1_LOC_452/Y INVX1_LOC_17/Y 0.01fF
C18207 INPUT_6 NAND2X1_LOC_836/B 0.02fF
C18208 NAND2X1_LOC_320/a_36_24# INVX1_LOC_31/Y 0.00fF
C18209 INPUT_3 INVX1_LOC_9/A 0.07fF
C18210 INVX1_LOC_21/Y INPUT_2 0.04fF
C18211 INVX1_LOC_490/Y INVX1_LOC_32/Y 0.03fF
C18212 INVX1_LOC_586/A INVX1_LOC_685/Y 0.03fF
C18213 INVX1_LOC_31/A INVX1_LOC_145/Y 0.01fF
C18214 INVX1_LOC_596/A INVX1_LOC_12/Y 0.02fF
C18215 INVX1_LOC_394/Y INVX1_LOC_26/Y 0.10fF
C18216 NAND2X1_LOC_7/a_36_24# INVX1_LOC_99/Y 0.01fF
C18217 INVX1_LOC_340/Y INVX1_LOC_637/A 0.03fF
C18218 NAND2X1_LOC_45/Y INVX1_LOC_58/Y 0.03fF
C18219 INVX1_LOC_224/Y INVX1_LOC_199/Y 0.07fF
C18220 INVX1_LOC_264/Y INVX1_LOC_69/Y 0.03fF
C18221 INVX1_LOC_435/Y NAND2X1_LOC_521/Y 0.42fF
C18222 INVX1_LOC_266/A INVX1_LOC_545/A 0.01fF
C18223 INVX1_LOC_68/Y NAND2X1_LOC_341/a_36_24# 0.00fF
C18224 INVX1_LOC_563/A INVX1_LOC_635/A 0.00fF
C18225 INVX1_LOC_21/Y INVX1_LOC_297/A 0.04fF
C18226 NAND2X1_LOC_370/A INVX1_LOC_31/Y 0.07fF
C18227 INVX1_LOC_68/Y INVX1_LOC_50/Y 0.71fF
C18228 INVX1_LOC_515/A NAND2X1_LOC_728/A 0.04fF
C18229 INVX1_LOC_415/Y INVX1_LOC_218/A 0.01fF
C18230 INVX1_LOC_99/Y INVX1_LOC_658/A 0.00fF
C18231 INVX1_LOC_412/Y INVX1_LOC_63/Y 0.03fF
C18232 INVX1_LOC_372/Y INVX1_LOC_504/A 0.05fF
C18233 INVX1_LOC_80/A INVX1_LOC_106/A 0.50fF
C18234 INVX1_LOC_428/A NAND2X1_LOC_106/Y 0.70fF
C18235 INVX1_LOC_105/A NAND2X1_LOC_332/B 0.01fF
C18236 INVX1_LOC_602/A INVX1_LOC_25/Y 0.20fF
C18237 INVX1_LOC_626/A INVX1_LOC_581/A 0.06fF
C18238 NAND2X1_LOC_768/A INVX1_LOC_106/A 0.01fF
C18239 INVX1_LOC_1/A INVX1_LOC_3/A 0.01fF
C18240 INVX1_LOC_117/Y INVX1_LOC_502/Y 0.03fF
C18241 NAND2X1_LOC_93/Y INVX1_LOC_353/A 0.03fF
C18242 NAND2X1_LOC_122/Y INVX1_LOC_31/Y 0.03fF
C18243 INVX1_LOC_446/Y NAND2X1_LOC_276/A 0.04fF
C18244 INVX1_LOC_51/Y INVX1_LOC_230/Y 0.00fF
C18245 INVX1_LOC_578/A INVX1_LOC_199/Y 0.07fF
C18246 INVX1_LOC_557/A INVX1_LOC_199/Y 2.72fF
C18247 NAND2X1_LOC_785/a_36_24# INVX1_LOC_600/A 0.00fF
C18248 NAND2X1_LOC_498/Y INVX1_LOC_58/Y 0.07fF
C18249 INVX1_LOC_20/Y INVX1_LOC_103/Y 0.03fF
C18250 INVX1_LOC_141/Y INVX1_LOC_45/Y 0.01fF
C18251 VDD NAND2X1_LOC_269/B 0.01fF
C18252 INVX1_LOC_312/Y INVX1_LOC_665/Y 0.03fF
C18253 INVX1_LOC_570/A INVX1_LOC_58/Y 0.06fF
C18254 INVX1_LOC_492/A INVX1_LOC_53/Y 0.06fF
C18255 INVX1_LOC_584/A INVX1_LOC_245/A 0.28fF
C18256 INVX1_LOC_21/Y INVX1_LOC_252/Y 0.03fF
C18257 INVX1_LOC_364/Y INVX1_LOC_69/Y 0.03fF
C18258 INVX1_LOC_370/Y INVX1_LOC_116/Y 0.00fF
C18259 INVX1_LOC_118/Y INVX1_LOC_26/Y 0.01fF
C18260 INVX1_LOC_49/Y INVX1_LOC_624/A 0.02fF
C18261 INVX1_LOC_127/A INVX1_LOC_128/A 0.00fF
C18262 NAND2X1_LOC_122/Y NAND2X1_LOC_675/B 0.23fF
C18263 INVX1_LOC_352/Y NAND2X1_LOC_603/Y 0.08fF
C18264 INVX1_LOC_145/Y NAND2X1_LOC_376/Y 0.04fF
C18265 INVX1_LOC_366/A INVX1_LOC_182/Y 0.03fF
C18266 NAND2X1_LOC_137/A INVX1_LOC_126/A 0.44fF
C18267 INVX1_LOC_191/A INVX1_LOC_6/Y 0.01fF
C18268 INVX1_LOC_84/A INVX1_LOC_173/Y 0.03fF
C18269 INVX1_LOC_632/A INVX1_LOC_259/Y 0.01fF
C18270 INVX1_LOC_400/Y INVX1_LOC_245/A 0.03fF
C18271 NAND2X1_LOC_140/B INVX1_LOC_371/A 0.10fF
C18272 INVX1_LOC_145/Y NAND2X1_LOC_69/Y 0.01fF
C18273 INVX1_LOC_116/A INVX1_LOC_197/Y 0.02fF
C18274 INVX1_LOC_588/Y INVX1_LOC_579/Y 0.03fF
C18275 INVX1_LOC_451/A NAND2X1_LOC_529/Y 0.02fF
C18276 INVX1_LOC_166/A INVX1_LOC_80/A 0.10fF
C18277 INVX1_LOC_117/Y INVX1_LOC_136/Y 0.04fF
C18278 INVX1_LOC_617/Y INVX1_LOC_253/Y 0.02fF
C18279 INVX1_LOC_211/Y INVX1_LOC_681/A 0.01fF
C18280 INVX1_LOC_579/A INVX1_LOC_93/Y 0.00fF
C18281 INVX1_LOC_549/Y INVX1_LOC_35/Y 0.05fF
C18282 INVX1_LOC_479/A NAND2X1_LOC_76/B 0.09fF
C18283 INVX1_LOC_537/Y INVX1_LOC_536/Y 0.01fF
C18284 INVX1_LOC_17/Y NAND2X1_LOC_670/a_36_24# 0.00fF
C18285 INVX1_LOC_32/Y INVX1_LOC_97/Y 0.04fF
C18286 INVX1_LOC_80/A INVX1_LOC_239/A 0.01fF
C18287 INVX1_LOC_659/A INVX1_LOC_59/A 0.00fF
C18288 INVX1_LOC_617/Y INVX1_LOC_63/Y 0.03fF
C18289 INVX1_LOC_176/Y INVX1_LOC_63/Y 0.00fF
C18290 NAND2X1_LOC_389/a_36_24# INVX1_LOC_600/A 0.00fF
C18291 INVX1_LOC_608/A INVX1_LOC_99/Y 0.03fF
C18292 NAND2X1_LOC_111/Y INVX1_LOC_80/A 0.01fF
C18293 INVX1_LOC_600/A INVX1_LOC_431/Y 0.12fF
C18294 NAND2X1_LOC_615/B INVX1_LOC_98/Y 0.03fF
C18295 INVX1_LOC_69/Y INVX1_LOC_134/Y 0.18fF
C18296 INVX1_LOC_197/A INVX1_LOC_496/A 0.17fF
C18297 INVX1_LOC_537/A NAND2X1_LOC_689/B 0.02fF
C18298 INVX1_LOC_49/Y INVX1_LOC_635/A 0.01fF
C18299 INVX1_LOC_361/Y NAND2X1_LOC_775/B 0.03fF
C18300 INVX1_LOC_167/A INVX1_LOC_137/Y 0.02fF
C18301 INVX1_LOC_674/A NAND2X1_LOC_807/a_36_24# 0.01fF
C18302 INVX1_LOC_490/A INVX1_LOC_367/Y 0.00fF
C18303 INVX1_LOC_20/Y NAND2X1_LOC_786/B 0.72fF
C18304 INVX1_LOC_157/A INVX1_LOC_99/Y 0.03fF
C18305 INVX1_LOC_482/A INVX1_LOC_79/A 0.01fF
C18306 INVX1_LOC_213/Y NAND2X1_LOC_184/Y 0.03fF
C18307 INVX1_LOC_676/Y INVX1_LOC_58/Y 0.03fF
C18308 INVX1_LOC_11/Y INVX1_LOC_166/A 0.91fF
C18309 INVX1_LOC_575/A INVX1_LOC_6/Y 0.03fF
C18310 INVX1_LOC_66/A INVX1_LOC_98/Y 0.05fF
C18311 INVX1_LOC_316/Y INVX1_LOC_69/Y 0.03fF
C18312 INVX1_LOC_431/A INVX1_LOC_32/Y 0.00fF
C18313 INVX1_LOC_320/A INVX1_LOC_9/Y 0.01fF
C18314 INVX1_LOC_145/Y NAND2X1_LOC_276/A 0.01fF
C18315 INVX1_LOC_99/Y NAND2X1_LOC_271/a_36_24# 0.01fF
C18316 INVX1_LOC_556/Y INVX1_LOC_89/Y 0.01fF
C18317 GATE_865 INVX1_LOC_686/Y 0.14fF
C18318 INVX1_LOC_47/Y INVX1_LOC_178/A 0.02fF
C18319 NAND2X1_LOC_557/B INVX1_LOC_178/A 0.02fF
C18320 INVX1_LOC_47/Y INVX1_LOC_251/Y 0.29fF
C18321 NAND2X1_LOC_32/Y INVX1_LOC_87/A 0.11fF
C18322 INVX1_LOC_99/Y INVX1_LOC_58/Y 0.60fF
C18323 INVX1_LOC_614/A INVX1_LOC_655/A 0.04fF
C18324 INVX1_LOC_80/A INVX1_LOC_153/Y 0.01fF
C18325 NAND2X1_LOC_697/a_36_24# INVX1_LOC_48/Y 0.00fF
C18326 INVX1_LOC_261/A INVX1_LOC_673/A 0.07fF
C18327 INVX1_LOC_204/Y INVX1_LOC_48/Y 0.03fF
C18328 INVX1_LOC_258/A NAND2X1_LOC_123/B 0.10fF
C18329 INVX1_LOC_80/A INVX1_LOC_531/Y 0.07fF
C18330 NAND2X1_LOC_689/B INVX1_LOC_496/Y 0.02fF
C18331 INVX1_LOC_537/A INVX1_LOC_245/A 0.03fF
C18332 INVX1_LOC_94/Y INVX1_LOC_32/Y 0.18fF
C18333 INVX1_LOC_320/A INVX1_LOC_62/Y 0.01fF
C18334 NAND2X1_LOC_274/B INVX1_LOC_35/Y 0.03fF
C18335 INVX1_LOC_471/Y NAND2X1_LOC_606/Y 0.38fF
C18336 INVX1_LOC_119/Y INVX1_LOC_251/Y 0.01fF
C18337 INVX1_LOC_6/Y INVX1_LOC_182/Y 0.05fF
C18338 NAND2X1_LOC_843/A INVX1_LOC_655/A 0.00fF
C18339 INVX1_LOC_580/Y INVX1_LOC_636/A 0.01fF
C18340 INVX1_LOC_194/A INVX1_LOC_79/A 0.01fF
C18341 INVX1_LOC_338/Y INVX1_LOC_66/A 0.03fF
C18342 NAND2X1_LOC_409/a_36_24# NAND2X1_LOC_409/Y 0.02fF
C18343 INVX1_LOC_303/Y INVX1_LOC_100/Y 0.03fF
C18344 INVX1_LOC_48/Y INVX1_LOC_114/A 0.03fF
C18345 INVX1_LOC_69/Y INVX1_LOC_65/A 0.00fF
C18346 INVX1_LOC_47/Y INVX1_LOC_58/Y 0.15fF
C18347 NAND2X1_LOC_557/B INVX1_LOC_58/Y 0.03fF
C18348 INVX1_LOC_300/A INVX1_LOC_635/Y 0.02fF
C18349 INVX1_LOC_166/A NAND2X1_LOC_433/Y 0.01fF
C18350 INVX1_LOC_80/A INVX1_LOC_363/A 0.01fF
C18351 INVX1_LOC_11/Y INVX1_LOC_531/Y 0.03fF
C18352 INVX1_LOC_292/Y NAND2X1_LOC_792/a_36_24# 0.00fF
C18353 NAND2X1_LOC_106/Y NAND2X1_LOC_106/a_36_24# 0.02fF
C18354 INVX1_LOC_369/Y INPUT_1 0.01fF
C18355 INVX1_LOC_32/Y NAND2X1_LOC_489/A 0.09fF
C18356 INVX1_LOC_206/Y INVX1_LOC_109/Y 0.01fF
C18357 NAND2X1_LOC_542/A INVX1_LOC_518/A 0.04fF
C18358 VDD INVX1_LOC_73/Y 0.26fF
C18359 INVX1_LOC_558/Y INVX1_LOC_92/A 0.05fF
C18360 INVX1_LOC_179/A INVX1_LOC_351/A 0.01fF
C18361 INVX1_LOC_95/Y INVX1_LOC_206/Y 0.01fF
C18362 INVX1_LOC_479/A INVX1_LOC_520/A 0.00fF
C18363 INVX1_LOC_58/Y INVX1_LOC_119/Y 0.03fF
C18364 NAND2X1_LOC_790/B INVX1_LOC_203/Y 0.03fF
C18365 INVX1_LOC_518/A INVX1_LOC_376/Y 0.12fF
C18366 INVX1_LOC_6/Y NAND2X1_LOC_615/a_36_24# 0.00fF
C18367 VDD NAND2X1_LOC_373/Y 0.09fF
C18368 INVX1_LOC_179/A INVX1_LOC_90/Y 0.03fF
C18369 INVX1_LOC_100/Y INVX1_LOC_9/Y 0.79fF
C18370 VDD INVX1_LOC_553/A -0.00fF
C18371 NAND2X1_LOC_249/Y INVX1_LOC_118/Y 0.04fF
C18372 INVX1_LOC_368/A INVX1_LOC_369/Y 0.00fF
C18373 INVX1_LOC_261/A INVX1_LOC_660/Y 0.27fF
C18374 NAND2X1_LOC_176/Y INVX1_LOC_560/A 0.09fF
C18375 INVX1_LOC_686/A INVX1_LOC_109/Y 0.07fF
C18376 NAND2X1_LOC_605/B INVX1_LOC_347/A 0.03fF
C18377 INVX1_LOC_74/Y INVX1_LOC_9/Y 0.07fF
C18378 NAND2X1_LOC_631/B INVX1_LOC_422/A 0.05fF
C18379 INVX1_LOC_68/Y INVX1_LOC_275/A 0.02fF
C18380 NAND2X1_LOC_686/A INVX1_LOC_479/A 0.01fF
C18381 INVX1_LOC_100/Y INVX1_LOC_62/Y 0.14fF
C18382 NAND2X1_LOC_636/A INVX1_LOC_76/Y 0.00fF
C18383 INVX1_LOC_448/Y INVX1_LOC_502/Y 0.01fF
C18384 INVX1_LOC_395/A INVX1_LOC_523/A 0.04fF
C18385 INVX1_LOC_505/Y INVX1_LOC_41/Y 0.11fF
C18386 INVX1_LOC_553/A INVX1_LOC_510/Y 0.02fF
C18387 INVX1_LOC_62/Y INVX1_LOC_74/Y 0.13fF
C18388 INVX1_LOC_395/A INVX1_LOC_72/Y 0.01fF
C18389 INVX1_LOC_206/Y NAND2X1_LOC_427/Y 0.03fF
C18390 INVX1_LOC_41/Y NAND2X1_LOC_231/B 0.02fF
C18391 INVX1_LOC_206/Y INVX1_LOC_126/Y 0.01fF
C18392 VDD INVX1_LOC_375/Y 0.21fF
C18393 NAND2X1_LOC_582/a_36_24# INVX1_LOC_685/Y 0.00fF
C18394 INVX1_LOC_249/Y INVX1_LOC_51/Y 0.02fF
C18395 NAND2X1_LOC_97/B INVX1_LOC_560/Y 0.01fF
C18396 NAND2X1_LOC_122/Y INVX1_LOC_51/Y 0.03fF
C18397 VDD INVX1_LOC_600/Y 0.46fF
C18398 INVX1_LOC_224/Y INVX1_LOC_53/Y 0.03fF
C18399 NAND2X1_LOC_332/B INVX1_LOC_45/Y 0.06fF
C18400 VDD NAND2X1_LOC_140/B 0.01fF
C18401 INVX1_LOC_404/Y NAND2X1_LOC_517/Y 0.08fF
C18402 INVX1_LOC_553/Y INVX1_LOC_670/Y 1.48fF
C18403 INVX1_LOC_54/A INVX1_LOC_7/Y 0.02fF
C18404 INVX1_LOC_578/A INVX1_LOC_53/Y 0.01fF
C18405 NAND2X1_LOC_331/A INVX1_LOC_161/A 0.01fF
C18406 INVX1_LOC_557/A INVX1_LOC_53/Y 0.04fF
C18407 INVX1_LOC_651/Y INVX1_LOC_654/A 0.05fF
C18408 INVX1_LOC_442/A NAND2X1_LOC_545/B 0.02fF
C18409 INVX1_LOC_560/Y INVX1_LOC_440/Y 0.02fF
C18410 INVX1_LOC_293/Y INVX1_LOC_384/A 0.07fF
C18411 INVX1_LOC_383/A INVX1_LOC_375/Y 0.01fF
C18412 INVX1_LOC_586/A INVX1_LOC_134/Y 0.17fF
C18413 INVX1_LOC_210/Y INPUT_0 0.00fF
C18414 INVX1_LOC_408/Y INVX1_LOC_98/Y 0.12fF
C18415 INVX1_LOC_418/A INVX1_LOC_99/A 0.00fF
C18416 GATE_741 NAND2X1_LOC_677/Y 0.02fF
C18417 INVX1_LOC_21/Y INVX1_LOC_85/Y 0.00fF
C18418 INVX1_LOC_561/Y INVX1_LOC_259/Y 0.72fF
C18419 VDD INVX1_LOC_627/Y 0.21fF
C18420 INVX1_LOC_361/Y NAND2X1_LOC_317/B 0.30fF
C18421 INVX1_LOC_442/A INVX1_LOC_98/Y 0.10fF
C18422 INVX1_LOC_237/Y INVX1_LOC_35/Y 0.02fF
C18423 INVX1_LOC_465/Y INVX1_LOC_49/Y 0.32fF
C18424 INVX1_LOC_248/Y INVX1_LOC_51/Y 0.04fF
C18425 INVX1_LOC_683/Y INVX1_LOC_519/A 0.03fF
C18426 INVX1_LOC_213/Y INVX1_LOC_607/A 0.74fF
C18427 INVX1_LOC_11/Y NAND2X1_LOC_778/a_36_24# 0.00fF
C18428 INVX1_LOC_11/Y INVX1_LOC_302/A 0.03fF
C18429 NAND2X1_LOC_638/A INVX1_LOC_111/A 0.00fF
C18430 INVX1_LOC_312/Y INVX1_LOC_134/Y 0.07fF
C18431 NAND2X1_LOC_307/A NAND2X1_LOC_304/a_36_24# 0.02fF
C18432 INVX1_LOC_202/Y INVX1_LOC_666/A 0.00fF
C18433 INVX1_LOC_76/Y INVX1_LOC_230/A -0.01fF
C18434 NAND2X1_LOC_773/A INVX1_LOC_145/Y 0.01fF
C18435 INVX1_LOC_492/A INVX1_LOC_555/Y 0.01fF
C18436 VDD INVX1_LOC_494/Y 0.26fF
C18437 NAND2X1_LOC_297/Y INVX1_LOC_45/Y 0.02fF
C18438 INVX1_LOC_206/Y INVX1_LOC_199/Y 0.25fF
C18439 INVX1_LOC_20/Y INVX1_LOC_360/Y 0.21fF
C18440 INVX1_LOC_444/Y INPUT_2 0.18fF
C18441 NAND2X1_LOC_475/A INVX1_LOC_58/Y 0.09fF
C18442 NAND2X1_LOC_538/B INVX1_LOC_35/Y 0.25fF
C18443 INVX1_LOC_293/Y INVX1_LOC_145/Y 0.10fF
C18444 INVX1_LOC_282/A INVX1_LOC_651/Y 0.00fF
C18445 INVX1_LOC_375/A INVX1_LOC_253/Y 0.01fF
C18446 NAND2X1_LOC_165/Y INVX1_LOC_586/A 0.03fF
C18447 INVX1_LOC_482/A INVX1_LOC_48/Y 0.00fF
C18448 INVX1_LOC_419/Y INVX1_LOC_551/Y 0.10fF
C18449 INVX1_LOC_378/A INVX1_LOC_48/Y 0.03fF
C18450 INVX1_LOC_581/A NAND2X1_LOC_678/a_36_24# 0.00fF
C18451 INVX1_LOC_648/Y INVX1_LOC_199/Y 0.03fF
C18452 INVX1_LOC_578/A NAND2X1_LOC_545/a_36_24# 0.00fF
C18453 INVX1_LOC_20/Y INVX1_LOC_105/A 0.00fF
C18454 INVX1_LOC_468/Y INVX1_LOC_53/Y 0.01fF
C18455 NAND2X1_LOC_45/Y INVX1_LOC_245/A 0.05fF
C18456 INVX1_LOC_166/A NAND2X1_LOC_704/B 0.00fF
C18457 INVX1_LOC_375/A INVX1_LOC_63/Y 0.01fF
C18458 INVX1_LOC_121/Y INVX1_LOC_518/A 0.03fF
C18459 INVX1_LOC_546/A INVX1_LOC_63/Y 0.00fF
C18460 INVX1_LOC_619/A INVX1_LOC_197/Y 0.07fF
C18461 INPUT_3 NAND2X1_LOC_297/Y 0.01fF
C18462 INVX1_LOC_413/Y INVX1_LOC_420/A 0.03fF
C18463 INVX1_LOC_85/Y INVX1_LOC_181/Y 0.01fF
C18464 INVX1_LOC_206/Y INVX1_LOC_272/A 0.01fF
C18465 NAND2X1_LOC_336/B INVX1_LOC_411/A 0.01fF
C18466 INVX1_LOC_409/A INVX1_LOC_652/A 0.13fF
C18467 NAND2X1_LOC_152/B INVX1_LOC_650/Y 0.04fF
C18468 INVX1_LOC_412/Y NAND2X1_LOC_299/a_36_24# 0.00fF
C18469 INVX1_LOC_586/A INVX1_LOC_65/A 0.00fF
C18470 INVX1_LOC_202/Y NAND2X1_LOC_72/Y 0.01fF
C18471 NAND2X1_LOC_527/Y INVX1_LOC_53/Y 0.08fF
C18472 INVX1_LOC_199/Y INVX1_LOC_242/A 0.07fF
C18473 INVX1_LOC_116/Y INVX1_LOC_98/Y 0.10fF
C18474 NAND2X1_LOC_65/Y INVX1_LOC_63/Y 0.01fF
C18475 NAND2X1_LOC_397/Y INVX1_LOC_83/Y 0.00fF
C18476 NAND2X1_LOC_148/A INVX1_LOC_240/A 0.04fF
C18477 INVX1_LOC_596/A INVX1_LOC_66/A 0.03fF
C18478 INVX1_LOC_7/Y NAND2X1_LOC_84/B 0.19fF
C18479 NAND2X1_LOC_673/B INVX1_LOC_145/Y 0.08fF
C18480 INVX1_LOC_131/A INVX1_LOC_239/A 0.17fF
C18481 INVX1_LOC_45/Y INVX1_LOC_242/Y 0.07fF
C18482 INVX1_LOC_686/A INVX1_LOC_199/Y 0.07fF
C18483 INVX1_LOC_584/A NAND2X1_LOC_597/Y 0.06fF
C18484 INVX1_LOC_406/Y INVX1_LOC_63/Y 0.03fF
C18485 INVX1_LOC_248/A INVX1_LOC_160/A 0.03fF
C18486 INVX1_LOC_35/Y INVX1_LOC_159/Y 0.10fF
C18487 INVX1_LOC_304/A INVX1_LOC_159/Y 0.00fF
C18488 INVX1_LOC_600/A NAND2X1_LOC_63/a_36_24# 0.01fF
C18489 INVX1_LOC_194/A INVX1_LOC_48/Y 0.00fF
C18490 INVX1_LOC_99/A INVX1_LOC_46/Y 0.00fF
C18491 INVX1_LOC_81/Y INVX1_LOC_194/Y 0.17fF
C18492 INVX1_LOC_100/A INVX1_LOC_7/Y 0.04fF
C18493 NAND2X1_LOC_545/B INVX1_LOC_255/A 0.01fF
C18494 INVX1_LOC_136/Y INVX1_LOC_58/Y 0.01fF
C18495 INVX1_LOC_17/Y INVX1_LOC_359/A 0.01fF
C18496 INVX1_LOC_45/Y INVX1_LOC_487/A 0.01fF
C18497 INVX1_LOC_357/A INVX1_LOC_463/Y 0.05fF
C18498 INVX1_LOC_12/Y NAND2X1_LOC_52/Y 0.00fF
C18499 NAND2X1_LOC_174/B INVX1_LOC_156/A 0.00fF
C18500 NAND2X1_LOC_697/Y INVX1_LOC_6/Y 0.03fF
C18501 INVX1_LOC_370/Y INVX1_LOC_69/Y 0.01fF
C18502 INVX1_LOC_137/Y INVX1_LOC_46/Y 0.18fF
C18503 INVX1_LOC_451/A INVX1_LOC_6/Y 0.06fF
C18504 NAND2X1_LOC_285/B NAND2X1_LOC_285/a_36_24# 0.00fF
C18505 INVX1_LOC_80/A INVX1_LOC_301/Y 0.09fF
C18506 INVX1_LOC_682/Y INVX1_LOC_519/A 0.01fF
C18507 INVX1_LOC_11/Y NAND2X1_LOC_627/a_36_24# 0.00fF
C18508 NAND2X1_LOC_757/a_36_24# INVX1_LOC_26/Y -0.02fF
C18509 INVX1_LOC_65/Y INVX1_LOC_479/A 0.06fF
C18510 INVX1_LOC_54/Y NAND2X1_LOC_444/A 0.07fF
C18511 INVX1_LOC_35/Y INVX1_LOC_212/Y 0.03fF
C18512 INVX1_LOC_128/A INVX1_LOC_519/A 0.35fF
C18513 INVX1_LOC_297/A INVX1_LOC_26/Y 0.03fF
C18514 INVX1_LOC_255/A INVX1_LOC_98/Y 0.10fF
C18515 INVX1_LOC_25/Y INVX1_LOC_58/Y 0.01fF
C18516 INVX1_LOC_6/Y INVX1_LOC_665/Y 0.01fF
C18517 INVX1_LOC_145/Y NAND2X1_LOC_240/A 0.02fF
C18518 INVX1_LOC_17/Y INVX1_LOC_480/A 0.05fF
C18519 INVX1_LOC_202/Y INVX1_LOC_351/Y 0.01fF
C18520 INVX1_LOC_243/A INVX1_LOC_9/Y 0.01fF
C18521 INVX1_LOC_575/Y INVX1_LOC_6/Y 0.03fF
C18522 NAND2X1_LOC_673/A INVX1_LOC_49/Y 0.02fF
C18523 INVX1_LOC_376/Y INVX1_LOC_352/A 0.07fF
C18524 INVX1_LOC_17/Y NAND2X1_LOC_121/Y 0.02fF
C18525 INVX1_LOC_213/Y NAND2X1_LOC_259/a_36_24# 0.00fF
C18526 INVX1_LOC_99/Y INVX1_LOC_245/A 0.36fF
C18527 NAND2X1_LOC_531/Y INPUT_1 0.15fF
C18528 INVX1_LOC_550/Y INVX1_LOC_168/Y 0.04fF
C18529 INVX1_LOC_81/Y INVX1_LOC_44/Y 0.03fF
C18530 NAND2X1_LOC_786/B NAND2X1_LOC_61/a_36_24# 0.00fF
C18531 INVX1_LOC_80/A INVX1_LOC_41/Y 6.60fF
C18532 INVX1_LOC_11/Y INVX1_LOC_301/Y 0.01fF
C18533 INVX1_LOC_47/Y NAND2X1_LOC_689/B 0.03fF
C18534 INVX1_LOC_53/Y INVX1_LOC_621/A 0.28fF
C18535 INVX1_LOC_492/A INVX1_LOC_662/A 0.03fF
C18536 INVX1_LOC_153/A INVX1_LOC_58/Y 0.08fF
C18537 INVX1_LOC_17/Y NAND2X1_LOC_301/B 0.03fF
C18538 INVX1_LOC_550/A INVX1_LOC_168/Y 0.02fF
C18539 INVX1_LOC_54/Y INVX1_LOC_183/A 0.07fF
C18540 INVX1_LOC_335/Y INVX1_LOC_505/Y 0.07fF
C18541 INVX1_LOC_344/A INVX1_LOC_74/Y 0.01fF
C18542 NAND2X1_LOC_531/Y INVX1_LOC_422/Y 0.09fF
C18543 INVX1_LOC_106/A NAND2X1_LOC_843/B 0.00fF
C18544 INVX1_LOC_652/A INVX1_LOC_352/Y 0.01fF
C18545 INVX1_LOC_54/Y INVX1_LOC_389/Y 0.01fF
C18546 INVX1_LOC_662/A INVX1_LOC_240/A 0.15fF
C18547 INVX1_LOC_501/A NAND2X1_LOC_453/a_36_24# 0.01fF
C18548 NAND2X1_LOC_628/Y INPUT_1 0.01fF
C18549 INVX1_LOC_123/A INVX1_LOC_245/A 0.01fF
C18550 INVX1_LOC_11/Y INVX1_LOC_41/Y 0.56fF
C18551 INVX1_LOC_369/Y INVX1_LOC_50/Y 0.00fF
C18552 INVX1_LOC_69/Y INVX1_LOC_351/A 0.01fF
C18553 INVX1_LOC_47/Y INVX1_LOC_245/A 0.25fF
C18554 INVX1_LOC_390/Y INVX1_LOC_109/Y 0.04fF
C18555 INVX1_LOC_69/Y INVX1_LOC_90/Y 0.10fF
C18556 INVX1_LOC_469/Y INVX1_LOC_62/Y 0.03fF
C18557 INVX1_LOC_257/A NAND2X1_LOC_109/a_36_24# 0.00fF
C18558 NAND2X1_LOC_413/Y INVX1_LOC_92/A 0.07fF
C18559 NAND2X1_LOC_181/A INVX1_LOC_62/Y 0.01fF
C18560 INVX1_LOC_223/A INVX1_LOC_50/Y 0.15fF
C18561 NAND2X1_LOC_558/B INVX1_LOC_9/Y 0.06fF
C18562 INVX1_LOC_50/Y INVX1_LOC_348/Y 0.01fF
C18563 INVX1_LOC_285/Y INVX1_LOC_79/A 0.01fF
C18564 INVX1_LOC_647/Y INVX1_LOC_46/Y 0.01fF
C18565 INVX1_LOC_79/A INVX1_LOC_9/Y 0.10fF
C18566 INVX1_LOC_119/Y INVX1_LOC_245/A 0.03fF
C18567 INVX1_LOC_74/Y INVX1_LOC_624/Y 0.03fF
C18568 NAND2X1_LOC_66/Y INVX1_LOC_245/A 0.04fF
C18569 NAND2X1_LOC_628/Y INVX1_LOC_487/Y 0.18fF
C18570 NAND2X1_LOC_433/Y INVX1_LOC_41/Y 0.07fF
C18571 INVX1_LOC_85/Y NAND2X1_LOC_86/a_36_24# 0.00fF
C18572 NAND2X1_LOC_558/B INVX1_LOC_62/Y 0.02fF
C18573 INVX1_LOC_166/Y INVX1_LOC_79/A 0.02fF
C18574 INVX1_LOC_422/Y INVX1_LOC_443/A 0.49fF
C18575 INVX1_LOC_62/Y INVX1_LOC_79/A 0.15fF
C18576 INVX1_LOC_549/A INVX1_LOC_139/A 0.04fF
C18577 NAND2X1_LOC_170/a_36_24# INVX1_LOC_76/Y 0.01fF
C18578 INPUT_0 NAND2X1_LOC_516/Y 0.01fF
C18579 INVX1_LOC_414/Y INVX1_LOC_414/A 0.01fF
C18580 VDD INVX1_LOC_562/Y 0.21fF
C18581 INVX1_LOC_459/Y INVX1_LOC_206/Y 0.02fF
C18582 INVX1_LOC_153/Y INVX1_LOC_91/Y 0.02fF
C18583 NAND2X1_LOC_390/a_36_24# NAND2X1_LOC_475/A 0.00fF
C18584 INVX1_LOC_230/A INVX1_LOC_192/A 0.05fF
C18585 INVX1_LOC_540/Y NAND2X1_LOC_707/A 0.01fF
C18586 VDD INVX1_LOC_401/A 0.00fF
C18587 NAND2X1_LOC_770/A INVX1_LOC_635/A 0.06fF
C18588 INVX1_LOC_432/A INVX1_LOC_109/Y 0.01fF
C18589 INVX1_LOC_681/A INVX1_LOC_297/Y 0.00fF
C18590 INVX1_LOC_75/Y INVX1_LOC_666/Y 0.07fF
C18591 INVX1_LOC_479/A INVX1_LOC_588/A 1.55fF
C18592 VDD INVX1_LOC_595/A -0.00fF
C18593 INVX1_LOC_1/A INVX1_LOC_5/Y 0.01fF
C18594 VDD INVX1_LOC_567/Y 0.36fF
C18595 INVX1_LOC_206/Y INVX1_LOC_53/Y 0.24fF
C18596 INVX1_LOC_20/Y NAND2X1_LOC_506/B 0.17fF
C18597 INVX1_LOC_442/Y INVX1_LOC_453/A 0.05fF
C18598 INVX1_LOC_20/Y INVX1_LOC_45/Y 1.72fF
C18599 INVX1_LOC_459/A INVX1_LOC_345/Y 0.00fF
C18600 INVX1_LOC_140/Y INVX1_LOC_134/Y 0.03fF
C18601 INVX1_LOC_601/A INVX1_LOC_198/Y 0.10fF
C18602 INVX1_LOC_312/Y NAND2X1_LOC_249/a_36_24# 0.01fF
C18603 INVX1_LOC_459/Y INVX1_LOC_686/A 0.01fF
C18604 INVX1_LOC_442/Y NAND2X1_LOC_271/B 0.01fF
C18605 INVX1_LOC_84/A INVX1_LOC_321/A 0.05fF
C18606 NAND2X1_LOC_23/a_36_24# INVX1_LOC_176/A 0.01fF
C18607 INVX1_LOC_565/Y INVX1_LOC_586/A 0.01fF
C18608 INPUT_0 INVX1_LOC_201/A 0.00fF
C18609 NAND2X1_LOC_615/B NAND2X1_LOC_76/B 0.02fF
C18610 INVX1_LOC_579/A INVX1_LOC_51/Y 0.68fF
C18611 VDD INVX1_LOC_612/Y 0.42fF
C18612 INVX1_LOC_20/Y INVX1_LOC_348/A 0.02fF
C18613 INVX1_LOC_51/Y INVX1_LOC_519/A 0.05fF
C18614 INVX1_LOC_76/Y INVX1_LOC_492/Y 0.02fF
C18615 NAND2X1_LOC_379/Y INVX1_LOC_366/A 0.01fF
C18616 INVX1_LOC_65/Y INVX1_LOC_12/Y 0.16fF
C18617 INVX1_LOC_560/A INVX1_LOC_252/Y 0.00fF
C18618 NAND2X1_LOC_185/a_36_24# INVX1_LOC_161/A 0.02fF
C18619 INVX1_LOC_206/Y INVX1_LOC_460/Y 0.10fF
C18620 INVX1_LOC_53/Y INVX1_LOC_242/A 0.03fF
C18621 INVX1_LOC_412/A NAND2X1_LOC_775/B 0.06fF
C18622 INVX1_LOC_312/A INVX1_LOC_235/Y 0.01fF
C18623 INVX1_LOC_416/A INVX1_LOC_416/Y 0.04fF
C18624 INVX1_LOC_300/A INVX1_LOC_45/Y 0.07fF
C18625 INVX1_LOC_218/Y INVX1_LOC_445/Y 0.02fF
C18626 INPUT_3 INVX1_LOC_21/A 0.10fF
C18627 INVX1_LOC_197/Y NAND2X1_LOC_506/B 0.01fF
C18628 INVX1_LOC_51/A INPUT_1 0.01fF
C18629 INVX1_LOC_45/Y INVX1_LOC_197/Y 0.03fF
C18630 INVX1_LOC_11/Y NAND2X1_LOC_362/a_36_24# 0.00fF
C18631 INVX1_LOC_53/Y INVX1_LOC_686/A 0.14fF
C18632 NAND2X1_LOC_543/B INVX1_LOC_58/Y 0.02fF
C18633 NAND2X1_LOC_98/a_36_24# INVX1_LOC_620/A 0.00fF
C18634 INVX1_LOC_587/A INVX1_LOC_316/Y 0.01fF
C18635 INPUT_0 INVX1_LOC_498/A 0.39fF
C18636 INVX1_LOC_549/A INVX1_LOC_32/Y 0.02fF
C18637 INVX1_LOC_402/Y NAND2X1_LOC_516/B 0.26fF
C18638 INVX1_LOC_681/A INVX1_LOC_76/Y 0.01fF
C18639 INVX1_LOC_428/A INVX1_LOC_50/Y 0.03fF
C18640 INVX1_LOC_413/Y INVX1_LOC_54/Y 0.27fF
C18641 INVX1_LOC_293/Y NAND2X1_LOC_260/Y 0.01fF
C18642 VDD NAND2X1_LOC_666/Y 0.01fF
C18643 INVX1_LOC_340/Y INVX1_LOC_259/Y 0.03fF
C18644 INVX1_LOC_437/Y INVX1_LOC_384/Y 0.13fF
C18645 INVX1_LOC_659/Y INVX1_LOC_673/A 0.10fF
C18646 INVX1_LOC_84/A NAND2X1_LOC_81/a_36_24# 0.00fF
C18647 NAND2X1_LOC_548/B INVX1_LOC_7/Y 0.08fF
C18648 NAND2X1_LOC_475/A NAND2X1_LOC_91/a_36_24# 0.00fF
C18649 INVX1_LOC_614/A INVX1_LOC_567/Y 0.12fF
C18650 NAND2X1_LOC_525/Y INVX1_LOC_387/Y 0.01fF
C18651 INVX1_LOC_21/Y INVX1_LOC_80/A 0.18fF
C18652 INVX1_LOC_68/Y INVX1_LOC_117/Y 0.00fF
C18653 INVX1_LOC_596/A INVX1_LOC_116/Y 0.12fF
C18654 INVX1_LOC_619/A INVX1_LOC_600/Y 0.01fF
C18655 INVX1_LOC_544/A INVX1_LOC_596/A 0.03fF
C18656 INVX1_LOC_134/Y INVX1_LOC_252/A 0.04fF
C18657 INVX1_LOC_45/A INVX1_LOC_40/Y 0.00fF
C18658 INVX1_LOC_17/Y NAND2X1_LOC_304/a_36_24# 0.01fF
C18659 INVX1_LOC_445/Y NAND2X1_LOC_256/a_36_24# 0.01fF
C18660 NAND2X1_LOC_475/A INVX1_LOC_245/A 0.01fF
C18661 INVX1_LOC_397/A INVX1_LOC_199/Y 0.15fF
C18662 NAND2X1_LOC_177/a_36_24# INPUT_1 0.00fF
C18663 INVX1_LOC_642/Y NAND2X1_LOC_749/Y 0.02fF
C18664 INVX1_LOC_686/A INVX1_LOC_460/Y 0.03fF
C18665 NAND2X1_LOC_789/A INVX1_LOC_191/A 0.07fF
C18666 INVX1_LOC_511/A INVX1_LOC_514/A 0.00fF
C18667 VDD NAND2X1_LOC_123/B 0.09fF
C18668 NAND2X1_LOC_708/A NAND2X1_LOC_513/A 0.05fF
C18669 INVX1_LOC_105/A INVX1_LOC_375/Y 0.12fF
C18670 NAND2X1_LOC_39/Y INVX1_LOC_31/Y 0.05fF
C18671 INVX1_LOC_35/Y NAND2X1_LOC_595/Y 0.03fF
C18672 INVX1_LOC_80/A NAND2X1_LOC_267/A 0.07fF
C18673 INVX1_LOC_21/Y INVX1_LOC_11/Y 1.61fF
C18674 INVX1_LOC_25/Y INVX1_LOC_1/Y 0.02fF
C18675 INVX1_LOC_54/Y INVX1_LOC_174/A 0.12fF
C18676 NAND2X1_LOC_307/A INVX1_LOC_46/Y 0.03fF
C18677 INVX1_LOC_384/A NAND2X1_LOC_344/B 0.05fF
C18678 INVX1_LOC_210/Y INVX1_LOC_145/Y 0.01fF
C18679 INVX1_LOC_586/A NAND2X1_LOC_669/a_36_24# 0.01fF
C18680 NAND2X1_LOC_140/B INVX1_LOC_105/A 0.11fF
C18681 NAND2X1_LOC_174/B INVX1_LOC_344/Y 0.15fF
C18682 VDD INVX1_LOC_329/Y 0.21fF
C18683 NAND2X1_LOC_137/A INVX1_LOC_80/A 0.03fF
C18684 INVX1_LOC_117/Y INVX1_LOC_600/A 0.08fF
C18685 INVX1_LOC_318/A INVX1_LOC_12/Y 0.00fF
C18686 INVX1_LOC_514/A NAND2X1_LOC_679/B 0.03fF
C18687 INVX1_LOC_76/Y INVX1_LOC_168/Y 0.11fF
C18688 VDD NAND2X1_LOC_428/Y -0.00fF
C18689 INVX1_LOC_32/Y NAND2X1_LOC_237/Y 0.13fF
C18690 NAND2X1_LOC_379/Y INVX1_LOC_6/Y 0.26fF
C18691 INVX1_LOC_330/A NAND2X1_LOC_407/a_36_24# 0.02fF
C18692 INVX1_LOC_185/Y INVX1_LOC_655/A 0.02fF
C18693 INVX1_LOC_603/A INVX1_LOC_252/Y 0.04fF
C18694 INVX1_LOC_85/Y INVX1_LOC_26/Y 0.51fF
C18695 NAND2X1_LOC_545/B INVX1_LOC_69/Y 0.47fF
C18696 INVX1_LOC_587/Y INVX1_LOC_59/Y 0.01fF
C18697 INVX1_LOC_340/Y INVX1_LOC_114/A 0.02fF
C18698 INVX1_LOC_288/A INVX1_LOC_112/Y 0.05fF
C18699 INVX1_LOC_586/A INVX1_LOC_90/Y 0.21fF
C18700 VDD INVX1_LOC_270/Y 0.65fF
C18701 INVX1_LOC_490/Y INVX1_LOC_75/Y 0.10fF
C18702 INVX1_LOC_550/A INVX1_LOC_137/Y 0.02fF
C18703 NAND2X1_LOC_184/Y INVX1_LOC_391/Y 0.05fF
C18704 INPUT_1 INVX1_LOC_371/A 0.00fF
C18705 INPUT_0 INVX1_LOC_211/A 0.08fF
C18706 NAND2X1_LOC_504/a_36_24# INVX1_LOC_35/Y 0.00fF
C18707 VDD INVX1_LOC_485/A -0.00fF
C18708 INVX1_LOC_235/Y INVX1_LOC_226/Y 0.02fF
C18709 INVX1_LOC_11/Y NAND2X1_LOC_267/A 0.07fF
C18710 INPUT_0 INVX1_LOC_64/Y 0.01fF
C18711 NAND2X1_LOC_768/A INVX1_LOC_107/Y 0.15fF
C18712 INVX1_LOC_416/A INVX1_LOC_46/Y 0.01fF
C18713 NAND2X1_LOC_41/Y INVX1_LOC_6/Y 0.01fF
C18714 INVX1_LOC_419/Y INVX1_LOC_46/Y 0.01fF
C18715 INVX1_LOC_451/A NAND2X1_LOC_294/Y 0.05fF
C18716 INVX1_LOC_12/Y INVX1_LOC_314/Y 0.03fF
C18717 VDD INVX1_LOC_92/A 1.63fF
C18718 INVX1_LOC_89/Y INVX1_LOC_304/Y 0.03fF
C18719 INVX1_LOC_31/Y INVX1_LOC_513/A 0.01fF
C18720 INPUT_3 NAND2X1_LOC_269/B 0.01fF
C18721 INVX1_LOC_69/Y INVX1_LOC_98/Y 0.12fF
C18722 INVX1_LOC_166/A INVX1_LOC_361/Y 0.11fF
C18723 INVX1_LOC_417/Y INVX1_LOC_9/Y 0.42fF
C18724 INVX1_LOC_361/Y NAND2X1_LOC_849/a_36_24# 0.00fF
C18725 NAND2X1_LOC_190/A NAND2X1_LOC_181/A 0.00fF
C18726 INVX1_LOC_155/A INVX1_LOC_48/Y 0.01fF
C18727 INVX1_LOC_93/Y INVX1_LOC_670/A 0.38fF
C18728 INVX1_LOC_254/Y INVX1_LOC_253/Y 0.00fF
C18729 NAND2X1_LOC_527/a_36_24# INVX1_LOC_26/Y 0.00fF
C18730 INVX1_LOC_117/Y INVX1_LOC_484/A 0.03fF
C18731 INVX1_LOC_588/Y INVX1_LOC_261/Y 0.03fF
C18732 INVX1_LOC_49/Y INVX1_LOC_137/Y 0.08fF
C18733 NAND2X1_LOC_27/Y NAND2X1_LOC_557/B 0.44fF
C18734 INVX1_LOC_490/Y NAND2X1_LOC_271/A 0.00fF
C18735 INVX1_LOC_682/A INVX1_LOC_145/Y 0.01fF
C18736 INVX1_LOC_437/Y NAND2X1_LOC_555/B 0.02fF
C18737 INVX1_LOC_160/A INVX1_LOC_242/Y 0.04fF
C18738 INVX1_LOC_50/Y NAND2X1_LOC_284/A 0.02fF
C18739 INVX1_LOC_520/A INVX1_LOC_66/A 0.01fF
C18740 INVX1_LOC_59/Y INVX1_LOC_9/Y 0.01fF
C18741 INVX1_LOC_254/Y INVX1_LOC_63/Y 0.05fF
C18742 INVX1_LOC_344/A INVX1_LOC_79/A 0.02fF
C18743 INVX1_LOC_659/Y INVX1_LOC_660/Y 0.01fF
C18744 NAND2X1_LOC_615/B NAND2X1_LOC_52/Y 0.00fF
C18745 INVX1_LOC_439/Y GATE_479 0.25fF
C18746 INVX1_LOC_177/A INVX1_LOC_179/A 0.34fF
C18747 INVX1_LOC_46/Y NAND2X1_LOC_342/A 0.01fF
C18748 INVX1_LOC_406/A INVX1_LOC_387/Y 0.01fF
C18749 INVX1_LOC_350/Y INVX1_LOC_624/Y 0.34fF
C18750 INVX1_LOC_255/A NAND2X1_LOC_442/a_36_24# 0.01fF
C18751 INVX1_LOC_62/Y INVX1_LOC_632/A 0.07fF
C18752 INVX1_LOC_417/Y INVX1_LOC_62/Y 0.03fF
C18753 INVX1_LOC_80/A INVX1_LOC_209/Y 0.01fF
C18754 INVX1_LOC_48/Y INVX1_LOC_9/Y 9.67fF
C18755 INVX1_LOC_74/A INVX1_LOC_29/Y 0.01fF
C18756 INVX1_LOC_183/A NAND2X1_LOC_404/a_36_24# 0.00fF
C18757 INVX1_LOC_510/Y INVX1_LOC_92/A 0.07fF
C18758 INVX1_LOC_62/Y NAND2X1_LOC_679/B 0.01fF
C18759 INVX1_LOC_537/Y INVX1_LOC_495/Y 0.58fF
C18760 INVX1_LOC_670/Y INVX1_LOC_479/A 0.49fF
C18761 INVX1_LOC_406/A INVX1_LOC_49/Y 0.01fF
C18762 NAND2X1_LOC_387/Y INVX1_LOC_399/Y 0.01fF
C18763 INVX1_LOC_367/Y INVX1_LOC_41/Y 0.03fF
C18764 INVX1_LOC_379/A INVX1_LOC_280/A 0.07fF
C18765 INVX1_LOC_62/Y INVX1_LOC_491/Y 0.63fF
C18766 INVX1_LOC_592/Y INVX1_LOC_63/Y 0.00fF
C18767 INVX1_LOC_153/Y NAND2X1_LOC_333/B 0.03fF
C18768 INVX1_LOC_502/A INVX1_LOC_46/Y 0.07fF
C18769 INVX1_LOC_199/Y INVX1_LOC_376/Y 0.07fF
C18770 NAND2X1_LOC_283/a_36_24# NAND2X1_LOC_847/A 0.01fF
C18771 INVX1_LOC_127/Y INVX1_LOC_519/Y 0.01fF
C18772 INVX1_LOC_62/Y INVX1_LOC_48/Y 1.08fF
C18773 INVX1_LOC_614/A INVX1_LOC_92/A 0.09fF
C18774 INVX1_LOC_519/Y INVX1_LOC_66/A 0.23fF
C18775 INVX1_LOC_480/Y INVX1_LOC_483/Y 0.24fF
C18776 NAND2X1_LOC_491/Y INVX1_LOC_9/Y 0.04fF
C18777 INVX1_LOC_159/Y INVX1_LOC_364/A 0.00fF
C18778 INVX1_LOC_26/Y INVX1_LOC_234/Y 0.02fF
C18779 INVX1_LOC_133/Y INVX1_LOC_570/Y 0.01fF
C18780 INVX1_LOC_17/Y INVX1_LOC_634/Y 0.19fF
C18781 INVX1_LOC_145/Y INVX1_LOC_622/Y 0.01fF
C18782 INVX1_LOC_47/Y NAND2X1_LOC_470/a_36_24# 0.00fF
C18783 INPUT_1 INVX1_LOC_441/A 0.18fF
C18784 INVX1_LOC_180/Y INVX1_LOC_181/A 0.02fF
C18785 INVX1_LOC_79/A INVX1_LOC_624/Y 0.09fF
C18786 INVX1_LOC_662/A INVX1_LOC_644/Y 0.03fF
C18787 INVX1_LOC_50/Y NAND2X1_LOC_832/A 0.27fF
C18788 INVX1_LOC_253/Y INVX1_LOC_479/A 0.11fF
C18789 INVX1_LOC_11/A INVX1_LOC_328/Y 0.15fF
C18790 INVX1_LOC_63/Y INVX1_LOC_479/A 2.58fF
C18791 INVX1_LOC_665/A INVX1_LOC_26/Y 0.03fF
C18792 NAND2X1_LOC_750/Y NAND2X1_LOC_789/B 0.14fF
C18793 INVX1_LOC_295/A INVX1_LOC_109/Y 0.03fF
C18794 NAND2X1_LOC_597/Y INVX1_LOC_119/Y 0.01fF
C18795 INVX1_LOC_41/Y INVX1_LOC_319/A 0.04fF
C18796 INVX1_LOC_429/Y INVX1_LOC_445/Y 0.03fF
C18797 INPUT_0 INVX1_LOC_288/A 0.05fF
C18798 INVX1_LOC_206/Y NAND2X1_LOC_383/Y 0.01fF
C18799 NAND2X1_LOC_98/a_36_24# INVX1_LOC_291/A 0.00fF
C18800 INVX1_LOC_564/A INVX1_LOC_315/Y 0.00fF
C18801 INVX1_LOC_41/Y INVX1_LOC_625/Y 0.02fF
C18802 NAND2X1_LOC_391/B INVX1_LOC_395/A 0.00fF
C18803 INVX1_LOC_276/A INVX1_LOC_107/A 0.01fF
C18804 VDD INVX1_LOC_679/Y 0.98fF
C18805 INVX1_LOC_84/A INVX1_LOC_410/Y 0.07fF
C18806 INVX1_LOC_438/A INVX1_LOC_489/Y 0.16fF
C18807 VDD INVX1_LOC_602/Y 0.51fF
C18808 INVX1_LOC_257/Y NAND2X1_LOC_123/A 0.01fF
C18809 INPUT_0 INVX1_LOC_448/A 0.03fF
C18810 INVX1_LOC_167/Y INVX1_LOC_76/Y 0.09fF
C18811 NAND2X1_LOC_39/Y INVX1_LOC_51/Y 0.06fF
C18812 VDD INVX1_LOC_681/Y 0.29fF
C18813 NAND2X1_LOC_317/A INVX1_LOC_251/A 0.13fF
C18814 INPUT_0 INVX1_LOC_145/Y 0.31fF
C18815 INVX1_LOC_20/Y NAND2X1_LOC_756/Y 0.39fF
C18816 INVX1_LOC_448/A NAND2X1_LOC_516/Y 0.00fF
C18817 VDD INPUT_1 1.66fF
C18818 NAND2X1_LOC_545/B INVX1_LOC_586/A 0.02fF
C18819 INVX1_LOC_45/Y NAND2X1_LOC_298/a_36_24# 0.01fF
C18820 INVX1_LOC_11/Y NAND2X1_LOC_710/B 0.03fF
C18821 INVX1_LOC_580/Y INVX1_LOC_632/A 0.01fF
C18822 NAND2X1_LOC_318/A NAND2X1_LOC_307/A 0.01fF
C18823 INVX1_LOC_133/Y NAND2X1_LOC_847/A 0.18fF
C18824 INVX1_LOC_668/A NAND2X1_LOC_820/A 0.06fF
C18825 VDD INVX1_LOC_292/Y 0.37fF
C18826 NAND2X1_LOC_743/a_36_24# INVX1_LOC_581/A 0.00fF
C18827 INVX1_LOC_21/Y NAND2X1_LOC_704/B 0.00fF
C18828 INVX1_LOC_11/Y INVX1_LOC_255/Y 0.13fF
C18829 INVX1_LOC_556/A INVX1_LOC_54/Y 0.10fF
C18830 VDD INVX1_LOC_422/Y 0.26fF
C18831 INVX1_LOC_586/A INVX1_LOC_98/Y 0.03fF
C18832 NAND2X1_LOC_498/B INVX1_LOC_137/Y 0.06fF
C18833 VDD INVX1_LOC_284/Y 0.21fF
C18834 INVX1_LOC_20/Y INVX1_LOC_160/A 0.03fF
C18835 INVX1_LOC_516/Y INVX1_LOC_98/Y 0.10fF
C18836 INVX1_LOC_65/Y NAND2X1_LOC_615/B 0.03fF
C18837 INVX1_LOC_163/Y INVX1_LOC_549/Y 0.96fF
C18838 INVX1_LOC_391/Y NAND2X1_LOC_486/B 0.05fF
C18839 INVX1_LOC_68/Y NAND2X1_LOC_76/A 0.01fF
C18840 NAND2X1_LOC_721/a_36_24# INVX1_LOC_93/Y 0.01fF
C18841 NAND2X1_LOC_335/B INVX1_LOC_58/Y 0.01fF
C18842 INVX1_LOC_76/Y INVX1_LOC_137/Y 0.10fF
C18843 INVX1_LOC_451/A INVX1_LOC_381/A 0.10fF
C18844 INVX1_LOC_402/Y INVX1_LOC_367/A 0.04fF
C18845 INVX1_LOC_17/Y INVX1_LOC_270/A 0.07fF
C18846 NAND2X1_LOC_756/Y INVX1_LOC_197/Y 0.07fF
C18847 INPUT_0 INVX1_LOC_141/Y 0.00fF
C18848 INVX1_LOC_383/A INPUT_1 0.01fF
C18849 INVX1_LOC_510/Y INPUT_1 0.07fF
C18850 INVX1_LOC_549/Y INVX1_LOC_522/Y 0.06fF
C18851 INVX1_LOC_537/Y INVX1_LOC_536/A 0.00fF
C18852 INVX1_LOC_206/Y INVX1_LOC_544/Y 0.01fF
C18853 INVX1_LOC_556/Y INVX1_LOC_126/A 0.01fF
C18854 INVX1_LOC_54/Y NAND2X1_LOC_180/B 0.00fF
C18855 INVX1_LOC_435/Y INVX1_LOC_69/Y 0.12fF
C18856 INVX1_LOC_63/A INVX1_LOC_35/Y 0.21fF
C18857 INVX1_LOC_32/Y INVX1_LOC_666/A 0.00fF
C18858 INVX1_LOC_199/Y INVX1_LOC_253/A 0.03fF
C18859 VDD INVX1_LOC_487/Y 0.22fF
C18860 INVX1_LOC_424/A INVX1_LOC_502/A 0.00fF
C18861 INVX1_LOC_446/A NAND2X1_LOC_528/Y 0.01fF
C18862 INVX1_LOC_558/A NAND2X1_LOC_307/B 0.07fF
C18863 NAND2X1_LOC_669/Y INVX1_LOC_35/Y 0.01fF
C18864 INVX1_LOC_276/A NAND2X1_LOC_285/A 0.00fF
C18865 INVX1_LOC_74/Y INVX1_LOC_638/A 0.14fF
C18866 INVX1_LOC_175/A INVX1_LOC_46/Y 0.09fF
C18867 INVX1_LOC_300/A INVX1_LOC_160/A 0.01fF
C18868 INVX1_LOC_607/Y INVX1_LOC_145/Y 0.02fF
C18869 INVX1_LOC_503/A NAND2X1_LOC_643/a_36_24# 0.00fF
C18870 INVX1_LOC_585/Y INVX1_LOC_174/A 0.03fF
C18871 INVX1_LOC_17/Y NAND2X1_LOC_755/B 2.83fF
C18872 INVX1_LOC_602/Y INVX1_LOC_684/A -0.00fF
C18873 INVX1_LOC_614/A INPUT_1 0.14fF
C18874 NAND2X1_LOC_299/Y NAND2X1_LOC_123/a_36_24# 0.00fF
C18875 INVX1_LOC_68/Y INVX1_LOC_58/Y 0.02fF
C18876 INVX1_LOC_249/A INVX1_LOC_578/Y 0.01fF
C18877 NAND2X1_LOC_331/A INVX1_LOC_79/A 0.19fF
C18878 INVX1_LOC_17/Y INVX1_LOC_211/Y 0.03fF
C18879 INVX1_LOC_651/Y INVX1_LOC_654/Y 0.05fF
C18880 INVX1_LOC_427/Y INVX1_LOC_437/A 0.18fF
C18881 INVX1_LOC_449/Y INVX1_LOC_442/Y 0.05fF
C18882 NAND2X1_LOC_121/Y NAND2X1_LOC_122/Y 0.06fF
C18883 INVX1_LOC_147/Y INVX1_LOC_58/Y 0.10fF
C18884 INVX1_LOC_584/Y NAND2X1_LOC_640/a_36_24# 0.01fF
C18885 INVX1_LOC_565/Y INVX1_LOC_6/Y 0.02fF
C18886 INVX1_LOC_578/A NAND2X1_LOC_545/A 0.06fF
C18887 INVX1_LOC_43/Y INVX1_LOC_54/Y 0.01fF
C18888 INVX1_LOC_187/A INVX1_LOC_187/Y 0.10fF
C18889 INVX1_LOC_342/A INVX1_LOC_69/A 0.05fF
C18890 NAND2X1_LOC_74/a_36_24# INVX1_LOC_98/Y 0.00fF
C18891 INVX1_LOC_596/A INVX1_LOC_69/Y 0.03fF
C18892 INVX1_LOC_21/Y INVX1_LOC_374/Y 0.03fF
C18893 INVX1_LOC_561/Y INVX1_LOC_62/Y 0.03fF
C18894 NAND2X1_LOC_45/Y INVX1_LOC_483/A 0.02fF
C18895 NAND2X1_LOC_714/a_36_24# INVX1_LOC_79/A 0.00fF
C18896 INVX1_LOC_159/Y INVX1_LOC_350/A 0.02fF
C18897 INVX1_LOC_439/Y INVX1_LOC_452/A 0.14fF
C18898 INVX1_LOC_224/Y INVX1_LOC_666/Y 0.07fF
C18899 INVX1_LOC_581/A NAND2X1_LOC_803/a_36_24# 0.00fF
C18900 INVX1_LOC_662/A INVX1_LOC_242/A 0.18fF
C18901 INVX1_LOC_53/Y NAND2X1_LOC_542/A 0.69fF
C18902 INVX1_LOC_371/A NAND2X1_LOC_465/a_36_24# 0.02fF
C18903 INVX1_LOC_298/A INVX1_LOC_145/Y 0.02fF
C18904 NAND2X1_LOC_307/A INVX1_LOC_49/Y 0.08fF
C18905 INVX1_LOC_35/Y INVX1_LOC_186/Y 0.03fF
C18906 INVX1_LOC_372/Y INVX1_LOC_63/Y 0.05fF
C18907 INVX1_LOC_374/A NAND2X1_LOC_118/a_36_24# 0.00fF
C18908 INPUT_1 INVX1_LOC_509/A 0.01fF
C18909 INVX1_LOC_545/Y INVX1_LOC_49/Y 0.02fF
C18910 VDD INVX1_LOC_443/Y 0.21fF
C18911 INVX1_LOC_479/Y NAND2X1_LOC_615/B 0.19fF
C18912 INVX1_LOC_435/A INVX1_LOC_93/Y 0.03fF
C18913 INVX1_LOC_17/Y INVX1_LOC_46/Y 0.07fF
C18914 INVX1_LOC_371/A INVX1_LOC_50/Y 0.00fF
C18915 NAND2X1_LOC_190/A INVX1_LOC_48/Y 0.06fF
C18916 INVX1_LOC_602/A NAND2X1_LOC_792/a_36_24# 0.00fF
C18917 NAND2X1_LOC_673/A INVX1_LOC_32/Y 0.01fF
C18918 INVX1_LOC_99/Y NAND2X1_LOC_753/Y 0.19fF
C18919 NAND2X1_LOC_822/a_36_24# INVX1_LOC_59/A 0.00fF
C18920 INVX1_LOC_578/A INVX1_LOC_666/Y 0.07fF
C18921 INVX1_LOC_12/Y INVX1_LOC_63/Y 0.09fF
C18922 INVX1_LOC_58/Y INVX1_LOC_600/A 0.08fF
C18923 INVX1_LOC_53/Y INVX1_LOC_376/Y 0.07fF
C18924 INVX1_LOC_236/A INVX1_LOC_555/A 0.02fF
C18925 INVX1_LOC_398/A INVX1_LOC_100/Y 0.30fF
C18926 INVX1_LOC_54/Y NAND2X1_LOC_708/a_36_24# 0.00fF
C18927 INVX1_LOC_293/Y INVX1_LOC_655/A 0.00fF
C18928 INVX1_LOC_54/Y NAND2X1_LOC_387/Y 0.66fF
C18929 INVX1_LOC_318/A NAND2X1_LOC_615/B 0.00fF
C18930 INVX1_LOC_103/Y INPUT_1 0.03fF
C18931 NAND2X1_LOC_511/a_36_24# INVX1_LOC_588/A 0.01fF
C18932 INVX1_LOC_293/Y NAND2X1_LOC_269/B 0.13fF
C18933 INVX1_LOC_486/Y INVX1_LOC_90/Y 0.03fF
C18934 INVX1_LOC_294/Y INVX1_LOC_90/Y 0.22fF
C18935 INVX1_LOC_80/A INVX1_LOC_26/Y 0.09fF
C18936 INVX1_LOC_80/A INVX1_LOC_128/Y 0.02fF
C18937 INVX1_LOC_344/A NAND2X1_LOC_434/B 0.00fF
C18938 NAND2X1_LOC_333/a_36_24# NAND2X1_LOC_333/B 0.00fF
C18939 INVX1_LOC_379/A INVX1_LOC_328/Y 0.07fF
C18940 NAND2X1_LOC_230/a_36_24# INVX1_LOC_94/A 0.01fF
C18941 INPUT_5 INVX1_LOC_29/A 0.19fF
C18942 INVX1_LOC_35/Y INVX1_LOC_328/Y 0.08fF
C18943 NAND2X1_LOC_307/B INVX1_LOC_46/Y 0.03fF
C18944 INVX1_LOC_680/A INVX1_LOC_670/Y 0.01fF
C18945 NAND2X1_LOC_733/a_36_24# INVX1_LOC_62/Y 0.01fF
C18946 INVX1_LOC_476/A INVX1_LOC_6/Y 0.03fF
C18947 INVX1_LOC_595/Y INVX1_LOC_48/A 0.01fF
C18948 INVX1_LOC_451/A INVX1_LOC_100/Y 0.10fF
C18949 INVX1_LOC_11/Y INVX1_LOC_26/Y 0.25fF
C18950 INVX1_LOC_479/A INVX1_LOC_387/A 0.06fF
C18951 INVX1_LOC_455/A INVX1_LOC_657/A -0.00fF
C18952 INVX1_LOC_391/A INVX1_LOC_63/Y 0.01fF
C18953 INVX1_LOC_360/Y NAND2X1_LOC_123/B 0.01fF
C18954 INVX1_LOC_100/Y INVX1_LOC_665/Y 0.03fF
C18955 INVX1_LOC_99/Y INVX1_LOC_652/Y 0.00fF
C18956 INVX1_LOC_670/A INVX1_LOC_128/A 0.12fF
C18957 INVX1_LOC_421/A NAND2X1_LOC_292/a_36_24# 0.00fF
C18958 INVX1_LOC_21/Y INVX1_LOC_625/Y 0.45fF
C18959 INVX1_LOC_376/A INVX1_LOC_49/Y 0.01fF
C18960 INVX1_LOC_31/Y NAND2X1_LOC_832/a_36_24# 0.00fF
C18961 INVX1_LOC_319/A NAND2X1_LOC_267/A 0.13fF
C18962 INVX1_LOC_172/A INVX1_LOC_11/A 0.02fF
C18963 INVX1_LOC_361/Y INVX1_LOC_41/Y 0.09fF
C18964 INVX1_LOC_41/Y NAND2X1_LOC_333/B 0.01fF
C18965 INVX1_LOC_442/Y INVX1_LOC_363/A 0.01fF
C18966 INVX1_LOC_6/Y INVX1_LOC_90/Y 0.02fF
C18967 NAND2X1_LOC_615/Y INVX1_LOC_9/Y 0.03fF
C18968 INVX1_LOC_50/Y INVX1_LOC_645/Y 0.01fF
C18969 INVX1_LOC_49/Y INVX1_LOC_502/A 0.07fF
C18970 INVX1_LOC_74/Y NAND2X1_LOC_203/a_36_24# 0.00fF
C18971 INVX1_LOC_261/Y INVX1_LOC_41/Y 0.03fF
C18972 VDD INVX1_LOC_181/A -0.00fF
C18973 NAND2X1_LOC_308/A INVX1_LOC_74/Y 0.29fF
C18974 INVX1_LOC_629/A INVX1_LOC_638/A 0.04fF
C18975 INVX1_LOC_598/A INVX1_LOC_622/Y 0.01fF
C18976 INVX1_LOC_353/A INVX1_LOC_245/A 0.03fF
C18977 INVX1_LOC_117/Y INVX1_LOC_348/Y 0.05fF
C18978 INVX1_LOC_47/Y INVX1_LOC_652/Y 0.02fF
C18979 NAND2X1_LOC_241/B INVX1_LOC_275/A 0.05fF
C18980 INVX1_LOC_47/Y INVX1_LOC_483/A 0.03fF
C18981 INVX1_LOC_518/Y INVX1_LOC_518/A 0.15fF
C18982 NAND2X1_LOC_789/B VDD 0.01fF
C18983 NAND2X1_LOC_823/Y INVX1_LOC_657/A 0.07fF
C18984 INVX1_LOC_107/Y NAND2X1_LOC_843/B -0.00fF
C18985 INVX1_LOC_31/Y NAND2X1_LOC_418/a_36_24# 0.00fF
C18986 INVX1_LOC_395/A INVX1_LOC_616/Y 0.00fF
C18987 NAND2X1_LOC_354/a_36_24# INVX1_LOC_638/A 0.02fF
C18988 INVX1_LOC_224/Y INVX1_LOC_490/Y 0.03fF
C18989 INVX1_LOC_119/Y INVX1_LOC_652/Y 0.01fF
C18990 INVX1_LOC_577/Y NAND2X1_LOC_590/a_36_24# 0.00fF
C18991 INVX1_LOC_491/A NAND2X1_LOC_609/a_36_24# 0.00fF
C18992 INVX1_LOC_490/Y INVX1_LOC_578/A 0.14fF
C18993 INVX1_LOC_393/Y NAND2X1_LOC_735/a_36_24# 0.00fF
C18994 NAND2X1_LOC_475/A NAND2X1_LOC_352/a_36_24# 0.00fF
C18995 VDD INVX1_LOC_156/Y 0.21fF
C18996 INVX1_LOC_380/A INVX1_LOC_321/Y 0.04fF
C18997 NAND2X1_LOC_45/a_36_24# INVX1_LOC_384/A 0.01fF
C18998 INVX1_LOC_580/Y INVX1_LOC_561/Y 0.02fF
C18999 INPUT_0 NAND2X1_LOC_332/B 0.03fF
C19000 INVX1_LOC_224/Y INVX1_LOC_353/Y 0.01fF
C19001 INVX1_LOC_628/A INVX1_LOC_638/A 0.02fF
C19002 INVX1_LOC_435/Y INVX1_LOC_586/A 0.03fF
C19003 NAND2X1_LOC_249/Y INVX1_LOC_80/A 2.80fF
C19004 INVX1_LOC_445/Y INVX1_LOC_384/Y 0.03fF
C19005 INVX1_LOC_99/Y INVX1_LOC_458/Y 0.01fF
C19006 INVX1_LOC_578/A INVX1_LOC_353/Y 0.02fF
C19007 NAND2X1_LOC_331/A INVX1_LOC_511/A 0.02fF
C19008 INPUT_6 INVX1_LOC_55/A 0.02fF
C19009 NAND2X1_LOC_152/B INVX1_LOC_523/A 0.04fF
C19010 VDD INVX1_LOC_428/Y 0.38fF
C19011 VDD INVX1_LOC_53/A -0.00fF
C19012 NAND2X1_LOC_717/a_36_24# INVX1_LOC_320/A 0.00fF
C19013 NAND2X1_LOC_475/A NAND2X1_LOC_117/a_36_24# 0.00fF
C19014 INVX1_LOC_372/Y INVX1_LOC_374/A 0.98fF
C19015 INVX1_LOC_32/A INVX1_LOC_17/Y 0.05fF
C19016 INVX1_LOC_142/A NAND2X1_LOC_155/a_36_24# 0.02fF
C19017 INVX1_LOC_11/Y NAND2X1_LOC_249/Y 0.10fF
C19018 INVX1_LOC_53/Y INVX1_LOC_253/A 0.00fF
C19019 INVX1_LOC_463/A INVX1_LOC_513/A 0.05fF
C19020 INVX1_LOC_469/Y INVX1_LOC_638/A 0.01fF
C19021 INVX1_LOC_317/Y NAND2X1_LOC_336/B 0.01fF
C19022 INVX1_LOC_21/Y INVX1_LOC_393/Y 0.05fF
C19023 INVX1_LOC_596/A INVX1_LOC_586/A 0.02fF
C19024 INVX1_LOC_402/Y INVX1_LOC_395/A 0.03fF
C19025 INVX1_LOC_53/Y NAND2X1_LOC_142/Y 0.00fF
C19026 INVX1_LOC_374/A NAND2X1_LOC_326/a_36_24# 0.00fF
C19027 INVX1_LOC_447/A INVX1_LOC_159/Y 0.12fF
C19028 NAND2X1_LOC_331/A INVX1_LOC_491/Y 0.01fF
C19029 VDD INVX1_LOC_50/Y 1.98fF
C19030 INVX1_LOC_435/A INVX1_LOC_395/A 0.07fF
C19031 INVX1_LOC_446/Y INVX1_LOC_145/Y 0.17fF
C19032 NAND2X1_LOC_307/A INVX1_LOC_76/Y -0.01fF
C19033 NAND2X1_LOC_106/Y NAND2X1_LOC_554/a_36_24# 0.00fF
C19034 INVX1_LOC_47/Y INVX1_LOC_458/Y 0.01fF
C19035 INVX1_LOC_404/Y INVX1_LOC_48/Y 0.03fF
C19036 INVX1_LOC_288/A INVX1_LOC_145/Y 0.07fF
C19037 INVX1_LOC_450/A INVX1_LOC_451/A 0.03fF
C19038 INVX1_LOC_521/Y INVX1_LOC_35/Y 0.17fF
C19039 NAND2X1_LOC_331/A INVX1_LOC_48/Y 0.01fF
C19040 NAND2X1_LOC_596/Y INVX1_LOC_50/Y 0.09fF
C19041 INVX1_LOC_400/Y INVX1_LOC_510/A 0.03fF
C19042 VDD INVX1_LOC_431/Y 0.45fF
C19043 INVX1_LOC_438/A INVX1_LOC_382/A 0.02fF
C19044 INVX1_LOC_193/A INVX1_LOC_410/Y 0.01fF
C19045 INVX1_LOC_448/A INVX1_LOC_384/A 0.91fF
C19046 INVX1_LOC_402/A INVX1_LOC_242/A 0.07fF
C19047 INVX1_LOC_312/Y INVX1_LOC_596/A 10.79fF
C19048 INVX1_LOC_49/Y INVX1_LOC_388/Y 0.01fF
C19049 INVX1_LOC_266/Y INVX1_LOC_35/Y 0.03fF
C19050 INVX1_LOC_392/A INVX1_LOC_392/Y 0.01fF
C19051 INVX1_LOC_384/A INVX1_LOC_145/Y 0.08fF
C19052 INVX1_LOC_85/Y INVX1_LOC_81/Y 0.01fF
C19053 INVX1_LOC_228/Y NAND2X1_LOC_389/a_36_24# 0.00fF
C19054 INVX1_LOC_17/Y NAND2X1_LOC_318/A 7.06fF
C19055 VDD INVX1_LOC_517/Y 0.25fF
C19056 INVX1_LOC_271/Y INVX1_LOC_48/Y 0.02fF
C19057 INVX1_LOC_383/A INVX1_LOC_50/Y 0.01fF
C19058 INVX1_LOC_504/A NAND2X1_LOC_440/a_36_24# 0.01fF
C19059 INVX1_LOC_446/Y INVX1_LOC_433/A 0.04fF
C19060 INVX1_LOC_79/A INVX1_LOC_638/A 0.07fF
C19061 INVX1_LOC_510/Y INVX1_LOC_50/Y 1.55fF
C19062 INVX1_LOC_197/A INVX1_LOC_99/Y 0.03fF
C19063 INVX1_LOC_367/A INVX1_LOC_669/Y 0.02fF
C19064 INVX1_LOC_392/Y INVX1_LOC_93/Y 0.01fF
C19065 NAND2X1_LOC_538/B INVX1_LOC_411/A 0.00fF
C19066 INVX1_LOC_213/Y INVX1_LOC_654/A 0.00fF
C19067 INVX1_LOC_11/Y NAND2X1_LOC_833/a_36_24# 0.01fF
C19068 NAND2X1_LOC_335/B INVX1_LOC_245/A 0.01fF
C19069 NAND2X1_LOC_106/Y INVX1_LOC_45/Y 0.01fF
C19070 INVX1_LOC_613/Y NAND2X1_LOC_612/A 0.05fF
C19071 NAND2X1_LOC_513/a_36_24# INVX1_LOC_516/A 0.01fF
C19072 INVX1_LOC_460/A INVX1_LOC_638/A 0.03fF
C19073 INVX1_LOC_140/Y INVX1_LOC_338/Y 0.47fF
C19074 INVX1_LOC_604/A INVX1_LOC_63/Y 0.01fF
C19075 NAND2X1_LOC_391/A INVX1_LOC_304/Y 0.28fF
C19076 INVX1_LOC_445/Y NAND2X1_LOC_555/B 0.03fF
C19077 INVX1_LOC_65/Y INVX1_LOC_255/A 0.02fF
C19078 INVX1_LOC_299/A INVX1_LOC_300/Y 0.01fF
C19079 NAND2X1_LOC_26/a_36_24# NAND2X1_LOC_836/B 0.01fF
C19080 NAND2X1_LOC_537/a_36_24# INVX1_LOC_173/A 0.00fF
C19081 INPUT_0 INVX1_LOC_484/Y 0.01fF
C19082 NAND2X1_LOC_416/Y INVX1_LOC_99/Y 0.03fF
C19083 INPUT_0 INVX1_LOC_242/Y 0.03fF
C19084 NAND2X1_LOC_24/Y INVX1_LOC_54/Y 0.03fF
C19085 INVX1_LOC_93/Y INVX1_LOC_524/Y 0.05fF
C19086 INVX1_LOC_80/A INVX1_LOC_603/A 0.03fF
C19087 INVX1_LOC_438/Y INVX1_LOC_244/Y 0.03fF
C19088 INVX1_LOC_17/Y INVX1_LOC_115/A 0.01fF
C19089 INVX1_LOC_366/Y NAND2X1_LOC_378/Y 0.45fF
C19090 NAND2X1_LOC_180/B INVX1_LOC_89/Y 0.02fF
C19091 INVX1_LOC_526/A INVX1_LOC_47/Y 0.03fF
C19092 INVX1_LOC_99/Y NAND2X1_LOC_285/B 0.01fF
C19093 INVX1_LOC_93/A INVX1_LOC_55/Y 0.00fF
C19094 INVX1_LOC_206/Y NAND2X1_LOC_545/A 0.00fF
C19095 INVX1_LOC_93/Y INVX1_LOC_367/A 0.14fF
C19096 INVX1_LOC_145/Y INVX1_LOC_661/Y 0.19fF
C19097 INVX1_LOC_561/A INVX1_LOC_686/A 0.00fF
C19098 INVX1_LOC_252/A INVX1_LOC_98/Y 0.65fF
C19099 INPUT_7 INVX1_LOC_342/A 0.01fF
C19100 INVX1_LOC_65/Y INVX1_LOC_179/A 0.12fF
C19101 NAND2X1_LOC_790/B NAND2X1_LOC_231/B 0.03fF
C19102 INVX1_LOC_17/Y INVX1_LOC_202/Y 0.05fF
C19103 INVX1_LOC_99/Y NAND2X1_LOC_106/B 0.07fF
C19104 NAND2X1_LOC_523/B INVX1_LOC_6/Y 0.01fF
C19105 NAND2X1_LOC_516/Y INVX1_LOC_242/Y 0.02fF
C19106 INVX1_LOC_370/A INVX1_LOC_116/Y 0.15fF
C19107 INVX1_LOC_522/A INVX1_LOC_515/Y 0.15fF
C19108 INPUT_0 INVX1_LOC_487/A 0.01fF
C19109 INVX1_LOC_594/Y NAND2X1_LOC_451/B 0.03fF
C19110 INVX1_LOC_21/Y NAND2X1_LOC_333/B 0.03fF
C19111 NAND2X1_LOC_174/B INVX1_LOC_99/Y 4.12fF
C19112 INVX1_LOC_53/Y INVX1_LOC_477/Y 0.01fF
C19113 INVX1_LOC_21/Y INVX1_LOC_281/A 0.09fF
C19114 INVX1_LOC_68/Y INVX1_LOC_245/A 0.03fF
C19115 INVX1_LOC_89/Y INVX1_LOC_188/Y 0.03fF
C19116 INVX1_LOC_47/Y INVX1_LOC_197/A 0.07fF
C19117 INVX1_LOC_264/Y INVX1_LOC_74/Y 0.05fF
C19118 NAND2X1_LOC_591/Y INVX1_LOC_99/Y 0.01fF
C19119 VDD INVX1_LOC_658/Y 0.22fF
C19120 INVX1_LOC_172/A INVX1_LOC_35/Y 0.01fF
C19121 INVX1_LOC_93/Y INVX1_LOC_516/A 0.01fF
C19122 INVX1_LOC_670/Y INVX1_LOC_66/A 0.02fF
C19123 INVX1_LOC_206/Y INVX1_LOC_666/Y 0.01fF
C19124 NAND2X1_LOC_507/a_36_24# INVX1_LOC_100/Y 0.00fF
C19125 INVX1_LOC_93/Y INVX1_LOC_669/Y 0.02fF
C19126 INVX1_LOC_364/Y INVX1_LOC_100/Y 0.04fF
C19127 INVX1_LOC_480/Y INVX1_LOC_48/Y 0.04fF
C19128 INVX1_LOC_173/Y INVX1_LOC_99/Y 0.09fF
C19129 INVX1_LOC_335/Y INVX1_LOC_261/Y 0.03fF
C19130 INVX1_LOC_439/Y INVX1_LOC_282/A 0.53fF
C19131 INVX1_LOC_105/Y INVX1_LOC_35/Y 0.01fF
C19132 INVX1_LOC_45/Y NAND2X1_LOC_123/B 0.09fF
C19133 INVX1_LOC_208/A INVX1_LOC_209/A 0.14fF
C19134 NAND2X1_LOC_334/B INVX1_LOC_59/A 0.15fF
C19135 INVX1_LOC_545/A INVX1_LOC_46/Y 0.01fF
C19136 INVX1_LOC_395/A INVX1_LOC_241/A 0.02fF
C19137 INVX1_LOC_145/Y INVX1_LOC_433/A 0.00fF
C19138 INVX1_LOC_76/Y INVX1_LOC_502/A 0.01fF
C19139 INVX1_LOC_17/Y INVX1_LOC_387/Y 0.05fF
C19140 INVX1_LOC_392/A INVX1_LOC_93/Y 0.00fF
C19141 INVX1_LOC_566/Y INVX1_LOC_26/Y 0.03fF
C19142 INVX1_LOC_105/A INPUT_1 0.07fF
C19143 INVX1_LOC_103/Y INVX1_LOC_50/Y 0.09fF
C19144 INVX1_LOC_625/A INVX1_LOC_69/Y 0.02fF
C19145 GATE_662 INVX1_LOC_35/Y 0.01fF
C19146 INVX1_LOC_49/Y INVX1_LOC_503/A 0.04fF
C19147 INVX1_LOC_26/Y NAND2X1_LOC_238/a_36_24# 0.00fF
C19148 INVX1_LOC_169/Y INVX1_LOC_48/Y 0.01fF
C19149 NAND2X1_LOC_507/A NAND2X1_LOC_387/Y 0.04fF
C19150 INVX1_LOC_251/A INVX1_LOC_199/Y 0.03fF
C19151 INVX1_LOC_345/Y INVX1_LOC_355/Y 0.98fF
C19152 INVX1_LOC_17/Y INVX1_LOC_49/Y 0.17fF
C19153 INVX1_LOC_197/A INVX1_LOC_119/Y 0.07fF
C19154 NAND2X1_LOC_181/A INVX1_LOC_665/Y 0.02fF
C19155 INVX1_LOC_403/Y INVX1_LOC_89/Y 0.01fF
C19156 NAND2X1_LOC_174/B INVX1_LOC_47/Y 0.38fF
C19157 NAND2X1_LOC_131/a_36_24# INVX1_LOC_9/Y 0.00fF
C19158 INVX1_LOC_100/Y INVX1_LOC_134/Y 0.17fF
C19159 INVX1_LOC_442/Y INVX1_LOC_301/Y 0.28fF
C19160 NAND2X1_LOC_387/Y INVX1_LOC_89/Y 0.07fF
C19161 NAND2X1_LOC_123/A INVX1_LOC_242/Y 0.42fF
C19162 INVX1_LOC_35/Y NAND2X1_LOC_846/B 0.01fF
C19163 NAND2X1_LOC_210/A INVX1_LOC_168/Y 0.04fF
C19164 NAND2X1_LOC_180/B NAND2X1_LOC_544/B 0.02fF
C19165 INVX1_LOC_62/Y INVX1_LOC_508/Y 0.00fF
C19166 INVX1_LOC_346/A INVX1_LOC_50/Y 0.30fF
C19167 NAND2X1_LOC_48/Y INVX1_LOC_100/Y 0.03fF
C19168 INVX1_LOC_18/Y INVX1_LOC_93/A 0.01fF
C19169 INVX1_LOC_47/A INVX1_LOC_100/Y 0.05fF
C19170 INVX1_LOC_379/A INVX1_LOC_224/A 0.06fF
C19171 INVX1_LOC_117/Y NAND2X1_LOC_284/A 0.05fF
C19172 INVX1_LOC_208/Y INVX1_LOC_69/Y 0.03fF
C19173 INVX1_LOC_307/A INVX1_LOC_41/Y 0.03fF
C19174 INVX1_LOC_173/Y INVX1_LOC_47/Y 0.01fF
C19175 INVX1_LOC_367/Y INVX1_LOC_26/Y 0.09fF
C19176 INVX1_LOC_686/A INVX1_LOC_666/Y 0.42fF
C19177 INVX1_LOC_134/Y INVX1_LOC_74/Y 0.14fF
C19178 INVX1_LOC_369/Y INVX1_LOC_281/Y 0.11fF
C19179 INVX1_LOC_93/Y INVX1_LOC_675/A 0.40fF
C19180 NAND2X1_LOC_427/Y INVX1_LOC_462/Y 0.14fF
C19181 INVX1_LOC_662/Y INVX1_LOC_106/Y 0.07fF
C19182 INVX1_LOC_137/Y INVX1_LOC_612/A 0.13fF
C19183 INVX1_LOC_117/Y NAND2X1_LOC_768/B 0.07fF
C19184 INVX1_LOC_442/Y INVX1_LOC_41/Y 0.07fF
C19185 INVX1_LOC_451/A NAND2X1_LOC_631/B 0.01fF
C19186 INVX1_LOC_63/Y INVX1_LOC_66/A 0.03fF
C19187 INVX1_LOC_11/Y NAND2X1_LOC_626/Y 0.05fF
C19188 INVX1_LOC_93/Y NAND2X1_LOC_334/B 0.01fF
C19189 INVX1_LOC_14/A INVX1_LOC_653/Y 0.02fF
C19190 INVX1_LOC_316/Y INVX1_LOC_74/Y 0.00fF
C19191 INVX1_LOC_382/A NAND2X1_LOC_293/a_36_24# 0.01fF
C19192 INVX1_LOC_75/Y INVX1_LOC_230/A 0.13fF
C19193 INVX1_LOC_93/Y NAND2X1_LOC_487/a_36_24# 0.00fF
C19194 INVX1_LOC_6/Y NAND2X1_LOC_41/a_36_24# 0.00fF
C19195 INVX1_LOC_223/A INVX1_LOC_178/A 0.04fF
C19196 INVX1_LOC_50/Y INVX1_LOC_635/Y 0.04fF
C19197 VDD INVX1_LOC_275/A 0.10fF
C19198 NAND2X1_LOC_679/A NAND2X1_LOC_676/a_36_24# 0.02fF
C19199 NAND2X1_LOC_646/A NAND2X1_LOC_646/B 0.01fF
C19200 NAND2X1_LOC_7/Y INPUT_0 0.03fF
C19201 NAND2X1_LOC_93/Y VDD -0.00fF
C19202 INVX1_LOC_62/Y INVX1_LOC_149/Y 0.01fF
C19203 INVX1_LOC_63/Y NAND2X1_LOC_601/Y 0.31fF
C19204 INVX1_LOC_65/A INVX1_LOC_74/Y 0.01fF
C19205 VDD INVX1_LOC_438/A 0.08fF
C19206 INPUT_0 INVX1_LOC_301/A 0.07fF
C19207 INVX1_LOC_479/A INVX1_LOC_496/A 0.07fF
C19208 INVX1_LOC_63/Y NAND2X1_LOC_621/B 0.01fF
C19209 INVX1_LOC_41/Y INVX1_LOC_471/Y 0.15fF
C19210 INVX1_LOC_58/Y INVX1_LOC_223/A 0.01fF
C19211 INVX1_LOC_63/Y NAND2X1_LOC_646/B 0.01fF
C19212 VDD INVX1_LOC_441/Y 0.21fF
C19213 INVX1_LOC_206/Y INVX1_LOC_490/Y 0.03fF
C19214 INVX1_LOC_586/A NAND2X1_LOC_76/B 0.09fF
C19215 INVX1_LOC_379/A INVX1_LOC_109/Y 0.10fF
C19216 INVX1_LOC_35/Y INVX1_LOC_109/Y 0.10fF
C19217 INVX1_LOC_89/A INVX1_LOC_92/A 0.13fF
C19218 NAND2X1_LOC_790/B INVX1_LOC_80/A 0.14fF
C19219 INVX1_LOC_632/A INVX1_LOC_638/A 0.09fF
C19220 INVX1_LOC_17/Y INVX1_LOC_297/Y 0.03fF
C19221 VDD INVX1_LOC_187/A -0.00fF
C19222 NAND2X1_LOC_152/Y INVX1_LOC_554/Y 0.18fF
C19223 INVX1_LOC_212/A INVX1_LOC_669/A -0.01fF
C19224 INVX1_LOC_20/Y INPUT_0 0.22fF
C19225 INVX1_LOC_619/A INVX1_LOC_181/A 0.03fF
C19226 INVX1_LOC_635/Y INVX1_LOC_658/Y 0.01fF
C19227 VDD NAND2X1_LOC_513/A 0.05fF
C19228 INVX1_LOC_95/Y INVX1_LOC_35/Y 0.01fF
C19229 INVX1_LOC_393/A INVX1_LOC_502/Y 0.01fF
C19230 INVX1_LOC_20/Y NAND2X1_LOC_516/Y 0.06fF
C19231 INVX1_LOC_554/A INVX1_LOC_35/Y 0.02fF
C19232 INVX1_LOC_617/Y INVX1_LOC_400/Y 0.09fF
C19233 NAND2X1_LOC_370/A INVX1_LOC_270/A 0.04fF
C19234 INVX1_LOC_446/A INVX1_LOC_159/A 0.03fF
C19235 NAND2X1_LOC_789/B INVX1_LOC_619/A 0.11fF
C19236 INVX1_LOC_206/Y INVX1_LOC_97/Y 0.02fF
C19237 INVX1_LOC_11/Y NAND2X1_LOC_790/B 0.09fF
C19238 INVX1_LOC_395/A INVX1_LOC_367/A 0.01fF
C19239 INVX1_LOC_48/Y INVX1_LOC_638/A 0.07fF
C19240 NAND2X1_LOC_516/B INVX1_LOC_51/Y 0.12fF
C19241 INVX1_LOC_384/A NAND2X1_LOC_332/B 0.07fF
C19242 INVX1_LOC_20/Y INVX1_LOC_286/A 0.16fF
C19243 NAND2X1_LOC_45/Y NAND2X1_LOC_179/Y 0.07fF
C19244 NAND2X1_LOC_467/A NAND2X1_LOC_707/A 0.02fF
C19245 INVX1_LOC_286/Y INVX1_LOC_76/Y 0.35fF
C19246 INVX1_LOC_95/Y INVX1_LOC_620/A 0.10fF
C19247 INPUT_0 INVX1_LOC_300/A 0.03fF
C19248 INPUT_0 INVX1_LOC_197/Y 0.03fF
C19249 INVX1_LOC_395/A INVX1_LOC_669/Y 0.03fF
C19250 INPUT_7 INVX1_LOC_4/Y 0.09fF
C19251 VDD INVX1_LOC_327/Y 0.26fF
C19252 NAND2X1_LOC_136/a_36_24# INVX1_LOC_367/A 0.00fF
C19253 INVX1_LOC_679/Y INVX1_LOC_45/Y 0.00fF
C19254 INVX1_LOC_11/Y INVX1_LOC_122/Y 0.05fF
C19255 INVX1_LOC_530/Y NAND2X1_LOC_616/Y 0.46fF
C19256 INVX1_LOC_206/Y INVX1_LOC_431/A 0.30fF
C19257 INVX1_LOC_11/Y INVX1_LOC_103/A 0.02fF
C19258 INVX1_LOC_402/Y INVX1_LOC_51/Y 0.03fF
C19259 INVX1_LOC_396/Y INVX1_LOC_97/Y 0.01fF
C19260 INVX1_LOC_448/A NAND2X1_LOC_332/B 0.07fF
C19261 NAND2X1_LOC_710/B INVX1_LOC_361/Y 0.02fF
C19262 INVX1_LOC_367/A INVX1_LOC_683/Y 0.02fF
C19263 NAND2X1_LOC_498/Y INVX1_LOC_510/A 0.00fF
C19264 INVX1_LOC_80/A INVX1_LOC_235/Y 0.08fF
C19265 VDD NAND2X1_LOC_388/A 0.61fF
C19266 INVX1_LOC_286/A INVX1_LOC_300/A 0.01fF
C19267 INVX1_LOC_84/A INVX1_LOC_12/Y 0.13fF
C19268 INVX1_LOC_392/A INVX1_LOC_362/Y 0.42fF
C19269 INVX1_LOC_166/A INVX1_LOC_215/Y 0.01fF
C19270 INVX1_LOC_395/A INVX1_LOC_93/Y 0.43fF
C19271 INVX1_LOC_17/Y INVX1_LOC_76/Y 0.21fF
C19272 INVX1_LOC_20/Y INVX1_LOC_607/Y 0.07fF
C19273 NAND2X1_LOC_788/A INVX1_LOC_63/Y 0.01fF
C19274 NAND2X1_LOC_434/B INVX1_LOC_638/A 0.05fF
C19275 INPUT_3 NAND2X1_LOC_671/a_36_24# 0.01fF
C19276 INVX1_LOC_614/A NAND2X1_LOC_513/A 0.07fF
C19277 INVX1_LOC_214/Y INVX1_LOC_651/Y 0.01fF
C19278 INVX1_LOC_428/A INVX1_LOC_608/A 0.44fF
C19279 INVX1_LOC_20/Y NAND2X1_LOC_686/a_36_24# 0.00fF
C19280 INVX1_LOC_384/A INVX1_LOC_503/Y 0.02fF
C19281 NAND2X1_LOC_591/a_36_24# INVX1_LOC_632/A 0.00fF
C19282 INVX1_LOC_206/Y INVX1_LOC_94/Y 0.04fF
C19283 INVX1_LOC_425/A INVX1_LOC_304/Y 0.01fF
C19284 INVX1_LOC_185/Y INPUT_1 0.03fF
C19285 INVX1_LOC_45/Y INPUT_1 0.09fF
C19286 INVX1_LOC_51/Y NAND2X1_LOC_603/a_36_24# 0.00fF
C19287 NAND2X1_LOC_164/Y INVX1_LOC_69/Y 0.27fF
C19288 INVX1_LOC_35/Y NAND2X1_LOC_698/a_36_24# 0.00fF
C19289 INVX1_LOC_401/Y INVX1_LOC_99/Y 0.01fF
C19290 INVX1_LOC_425/A NAND2X1_LOC_551/a_36_24# 0.03fF
C19291 INVX1_LOC_93/Y INVX1_LOC_362/Y 0.07fF
C19292 INVX1_LOC_35/Y INVX1_LOC_126/Y 0.03fF
C19293 INVX1_LOC_435/Y INVX1_LOC_6/Y 0.01fF
C19294 INVX1_LOC_20/Y NAND2X1_LOC_859/a_36_24# 0.01fF
C19295 INVX1_LOC_377/Y INVX1_LOC_510/A 0.01fF
C19296 INVX1_LOC_21/Y INVX1_LOC_307/A 0.00fF
C19297 NAND2X1_LOC_531/Y NAND2X1_LOC_529/a_36_24# 0.00fF
C19298 INVX1_LOC_11/Y INVX1_LOC_235/Y 0.08fF
C19299 NAND2X1_LOC_173/Y INVX1_LOC_117/Y 0.03fF
C19300 INVX1_LOC_267/A INVX1_LOC_51/Y 0.07fF
C19301 INVX1_LOC_269/A INVX1_LOC_89/Y 0.52fF
C19302 INVX1_LOC_442/A INVX1_LOC_253/Y 0.55fF
C19303 INVX1_LOC_412/A INVX1_LOC_411/Y 0.01fF
C19304 INVX1_LOC_548/A INVX1_LOC_367/A 0.04fF
C19305 NAND2X1_LOC_592/B INVX1_LOC_49/Y 0.01fF
C19306 NAND2X1_LOC_184/a_36_24# NAND2X1_LOC_274/B -0.00fF
C19307 INVX1_LOC_129/A INVX1_LOC_12/Y 0.00fF
C19308 INVX1_LOC_130/Y INVX1_LOC_99/A 0.14fF
C19309 NAND2X1_LOC_68/a_36_24# INVX1_LOC_41/Y 0.00fF
C19310 INVX1_LOC_45/Y INVX1_LOC_292/Y 0.00fF
C19311 INVX1_LOC_80/A INVX1_LOC_556/Y 0.03fF
C19312 INVX1_LOC_255/Y INVX1_LOC_258/Y 0.37fF
C19313 INVX1_LOC_65/Y INVX1_LOC_69/Y 11.29fF
C19314 INVX1_LOC_20/Y INVX1_LOC_298/A 0.07fF
C19315 INVX1_LOC_11/Y NAND2X1_LOC_361/a_36_24# 0.00fF
C19316 INVX1_LOC_428/A INVX1_LOC_58/Y 0.03fF
C19317 INVX1_LOC_544/A INVX1_LOC_670/Y 0.02fF
C19318 INVX1_LOC_21/Y INVX1_LOC_442/Y 0.08fF
C19319 INPUT_3 INPUT_1 0.06fF
C19320 INVX1_LOC_395/A INVX1_LOC_390/A 0.00fF
C19321 INVX1_LOC_145/Y NAND2X1_LOC_260/Y 0.03fF
C19322 INVX1_LOC_556/Y NAND2X1_LOC_768/A 0.02fF
C19323 INVX1_LOC_300/A NAND2X1_LOC_123/A 0.02fF
C19324 INVX1_LOC_442/A INVX1_LOC_63/Y 0.07fF
C19325 INVX1_LOC_448/A INVX1_LOC_503/Y 0.03fF
C19326 INVX1_LOC_632/A INVX1_LOC_685/Y 0.14fF
C19327 INVX1_LOC_325/Y INVX1_LOC_46/Y 0.04fF
C19328 INVX1_LOC_342/A INVX1_LOC_55/Y 0.07fF
C19329 INVX1_LOC_395/A NAND2X1_LOC_334/B 0.00fF
C19330 NAND2X1_LOC_260/Y INVX1_LOC_661/Y 0.02fF
C19331 INVX1_LOC_210/Y INVX1_LOC_600/Y 0.24fF
C19332 NAND2X1_LOC_7/Y INVX1_LOC_211/A 0.06fF
C19333 INVX1_LOC_586/A NAND2X1_LOC_52/Y 0.01fF
C19334 NAND2X1_LOC_717/a_36_24# NAND2X1_LOC_558/B 0.00fF
C19335 INVX1_LOC_393/Y INVX1_LOC_26/Y 0.07fF
C19336 INVX1_LOC_367/Y NAND2X1_LOC_275/Y 1.97fF
C19337 NAND2X1_LOC_249/Y NAND2X1_LOC_843/B 0.01fF
C19338 NAND2X1_LOC_106/Y INVX1_LOC_293/Y 0.03fF
C19339 INVX1_LOC_545/A NAND2X1_LOC_703/a_36_24# 0.02fF
C19340 INVX1_LOC_21/Y INVX1_LOC_83/Y 0.02fF
C19341 INPUT_0 NAND2X1_LOC_269/B 0.05fF
C19342 INVX1_LOC_662/A NAND2X1_LOC_142/Y 0.07fF
C19343 INVX1_LOC_80/A INVX1_LOC_506/A 0.01fF
C19344 INVX1_LOC_469/Y INVX1_LOC_134/Y 0.03fF
C19345 INVX1_LOC_395/A NAND2X1_LOC_624/a_36_24# 0.01fF
C19346 INVX1_LOC_596/A INVX1_LOC_6/Y 0.03fF
C19347 INVX1_LOC_285/A INVX1_LOC_620/A 0.08fF
C19348 NAND2X1_LOC_588/a_36_24# INVX1_LOC_298/A 0.00fF
C19349 INVX1_LOC_300/A INVX1_LOC_527/Y 0.03fF
C19350 NAND2X1_LOC_697/Y INVX1_LOC_48/Y 0.01fF
C19351 INVX1_LOC_84/A INVX1_LOC_170/A 0.00fF
C19352 INVX1_LOC_598/A INVX1_LOC_145/Y 0.00fF
C19353 INVX1_LOC_412/A INVX1_LOC_41/Y 0.00fF
C19354 NAND2X1_LOC_181/A INVX1_LOC_134/Y 0.01fF
C19355 NAND2X1_LOC_393/Y INVX1_LOC_46/Y 0.00fF
C19356 INVX1_LOC_183/A INPUT_2 0.01fF
C19357 NAND2X1_LOC_775/B INVX1_LOC_159/Y 1.48fF
C19358 INVX1_LOC_31/Y INVX1_LOC_516/A 0.03fF
C19359 NAND2X1_LOC_318/B INVX1_LOC_6/Y 0.01fF
C19360 NAND2X1_LOC_336/B INVX1_LOC_411/Y 0.02fF
C19361 INVX1_LOC_662/Y INVX1_LOC_221/Y 0.03fF
C19362 INVX1_LOC_93/Y INVX1_LOC_189/Y 0.01fF
C19363 NAND2X1_LOC_192/a_36_24# NAND2X1_LOC_192/A 0.00fF
C19364 NAND2X1_LOC_128/A INVX1_LOC_99/Y 0.08fF
C19365 INVX1_LOC_166/A NAND2X1_LOC_317/a_36_24# 0.00fF
C19366 INVX1_LOC_272/Y INVX1_LOC_622/A 0.01fF
C19367 INVX1_LOC_525/Y INVX1_LOC_99/Y 1.24fF
C19368 INVX1_LOC_665/Y INVX1_LOC_48/Y 0.03fF
C19369 INVX1_LOC_402/A NAND2X1_LOC_542/A 0.56fF
C19370 INVX1_LOC_604/Y INVX1_LOC_69/Y 0.11fF
C19371 INVX1_LOC_548/A INVX1_LOC_93/Y 0.28fF
C19372 INVX1_LOC_400/A INVX1_LOC_31/Y 0.03fF
C19373 INVX1_LOC_105/A INVX1_LOC_50/Y 0.02fF
C19374 INVX1_LOC_197/A INVX1_LOC_15/Y 0.01fF
C19375 INVX1_LOC_28/Y INVX1_LOC_9/Y 0.01fF
C19376 NAND2X1_LOC_231/A INVX1_LOC_531/Y 0.02fF
C19377 INPUT_3 INVX1_LOC_368/A 0.00fF
C19378 INVX1_LOC_253/Y INVX1_LOC_116/Y 0.02fF
C19379 NAND2X1_LOC_707/A INVX1_LOC_41/Y 0.36fF
C19380 INVX1_LOC_158/Y NAND2X1_LOC_388/A 0.01fF
C19381 INVX1_LOC_161/A INVX1_LOC_338/Y 0.00fF
C19382 INVX1_LOC_358/A INVX1_LOC_357/Y 0.12fF
C19383 INVX1_LOC_603/Y INVX1_LOC_44/Y 0.09fF
C19384 INVX1_LOC_177/A INVX1_LOC_6/Y 0.03fF
C19385 INVX1_LOC_551/A NAND2X1_LOC_72/Y 0.01fF
C19386 INVX1_LOC_69/Y INVX1_LOC_370/A 0.01fF
C19387 INVX1_LOC_47/Y INVX1_LOC_510/A 0.04fF
C19388 NAND2X1_LOC_47/a_36_24# NAND2X1_LOC_836/B 0.00fF
C19389 INVX1_LOC_35/Y INVX1_LOC_199/Y 0.15fF
C19390 INVX1_LOC_564/Y INVX1_LOC_91/Y 0.01fF
C19391 INVX1_LOC_298/Y INVX1_LOC_659/A 0.02fF
C19392 INVX1_LOC_684/Y INVX1_LOC_674/Y 0.01fF
C19393 INVX1_LOC_63/Y INVX1_LOC_116/Y 0.03fF
C19394 NAND2X1_LOC_180/B INVX1_LOC_347/A 0.04fF
C19395 INVX1_LOC_256/A INVX1_LOC_376/A 0.05fF
C19396 INVX1_LOC_93/Y INVX1_LOC_31/Y 0.19fF
C19397 INVX1_LOC_134/Y INVX1_LOC_79/A 0.27fF
C19398 INVX1_LOC_504/A NAND2X1_LOC_437/a_36_24# 0.01fF
C19399 INVX1_LOC_20/Y INVX1_LOC_211/A 0.07fF
C19400 NAND2X1_LOC_594/Y INVX1_LOC_168/Y 0.04fF
C19401 INVX1_LOC_20/Y INVX1_LOC_464/Y 0.03fF
C19402 INVX1_LOC_370/Y INVX1_LOC_100/Y 0.01fF
C19403 INVX1_LOC_318/Y INVX1_LOC_74/Y 0.01fF
C19404 INVX1_LOC_17/Y NAND2X1_LOC_264/a_36_24# 0.00fF
C19405 INVX1_LOC_63/Y INVX1_LOC_328/A 0.03fF
C19406 INVX1_LOC_35/Y INVX1_LOC_272/A 0.00fF
C19407 INVX1_LOC_93/Y NAND2X1_LOC_675/B 0.01fF
C19408 INVX1_LOC_507/Y INVX1_LOC_186/Y 0.16fF
C19409 INVX1_LOC_376/A INVX1_LOC_345/Y 0.01fF
C19410 INVX1_LOC_455/Y INVX1_LOC_74/Y 0.04fF
C19411 INVX1_LOC_31/Y INVX1_LOC_675/A 0.07fF
C19412 NAND2X1_LOC_846/B INVX1_LOC_649/A 0.05fF
C19413 INVX1_LOC_119/Y INVX1_LOC_510/A 0.18fF
C19414 INVX1_LOC_437/A INVX1_LOC_430/A 0.01fF
C19415 INVX1_LOC_253/Y INVX1_LOC_255/A 0.07fF
C19416 INVX1_LOC_235/Y INVX1_LOC_231/Y 0.02fF
C19417 INVX1_LOC_31/Y NAND2X1_LOC_334/B 0.14fF
C19418 INVX1_LOC_75/Y NAND2X1_LOC_72/Y 0.01fF
C19419 NAND2X1_LOC_720/A INVX1_LOC_90/Y 0.07fF
C19420 INVX1_LOC_248/A INVX1_LOC_242/Y 0.04fF
C19421 NAND2X1_LOC_286/A NAND2X1_LOC_342/A 0.03fF
C19422 INVX1_LOC_99/Y NAND2X1_LOC_248/B 0.00fF
C19423 INVX1_LOC_54/Y INVX1_LOC_114/A 0.05fF
C19424 INVX1_LOC_255/A INVX1_LOC_63/Y 0.07fF
C19425 INVX1_LOC_210/A INVX1_LOC_198/A 0.24fF
C19426 INVX1_LOC_58/Y NAND2X1_LOC_52/a_36_24# 0.01fF
C19427 INVX1_LOC_32/Y INVX1_LOC_502/A 0.07fF
C19428 INVX1_LOC_54/Y NAND2X1_LOC_782/a_36_24# 0.00fF
C19429 INVX1_LOC_353/A NAND2X1_LOC_753/Y 0.17fF
C19430 INVX1_LOC_63/Y INVX1_LOC_179/A 0.03fF
C19431 NAND2X1_LOC_192/A INVX1_LOC_338/Y 0.02fF
C19432 INVX1_LOC_655/A INVX1_LOC_476/Y 0.06fF
C19433 GATE_865 INVX1_LOC_479/A 0.07fF
C19434 INVX1_LOC_160/A INVX1_LOC_270/Y 0.00fF
C19435 NAND2X1_LOC_635/B NAND2X1_LOC_451/B 0.16fF
C19436 INVX1_LOC_66/A INVX1_LOC_669/A 0.29fF
C19437 INVX1_LOC_117/Y INVX1_LOC_645/Y 0.03fF
C19438 INVX1_LOC_63/Y NAND2X1_LOC_262/a_36_24# 0.00fF
C19439 INVX1_LOC_625/Y INVX1_LOC_603/A 0.01fF
C19440 INVX1_LOC_395/A INVX1_LOC_615/Y 0.03fF
C19441 INVX1_LOC_62/Y INVX1_LOC_493/Y 0.01fF
C19442 NAND2X1_LOC_532/Y INVX1_LOC_479/A 0.02fF
C19443 INVX1_LOC_100/Y INVX1_LOC_351/A 0.03fF
C19444 INVX1_LOC_6/Y NAND2X1_LOC_411/a_36_24# 0.00fF
C19445 INVX1_LOC_257/Y INVX1_LOC_301/A 0.03fF
C19446 NAND2X1_LOC_542/A INVX1_LOC_666/Y 0.07fF
C19447 INVX1_LOC_369/Y INVX1_LOC_245/A 0.05fF
C19448 INVX1_LOC_100/Y INVX1_LOC_90/Y 0.14fF
C19449 INVX1_LOC_74/Y INVX1_LOC_351/A 0.03fF
C19450 NAND2X1_LOC_711/a_36_24# INVX1_LOC_558/A 0.00fF
C19451 VDD INVX1_LOC_289/Y 0.21fF
C19452 INVX1_LOC_376/Y INVX1_LOC_666/Y 0.02fF
C19453 INVX1_LOC_74/Y INVX1_LOC_90/Y 0.08fF
C19454 INVX1_LOC_400/Y INVX1_LOC_375/A 0.01fF
C19455 NAND2X1_LOC_415/a_36_24# INVX1_LOC_245/A 0.00fF
C19456 VDD INVX1_LOC_111/A 0.00fF
C19457 NAND2X1_LOC_164/Y INVX1_LOC_586/A 0.18fF
C19458 VDD INVX1_LOC_602/A 0.11fF
C19459 INVX1_LOC_20/Y INVX1_LOC_257/Y 0.03fF
C19460 VDD NAND2X1_LOC_636/B 0.01fF
C19461 VDD INVX1_LOC_104/Y 0.21fF
C19462 INVX1_LOC_381/A NAND2X1_LOC_42/a_36_24# 0.00fF
C19463 INVX1_LOC_65/Y INVX1_LOC_586/A 0.03fF
C19464 NAND2X1_LOC_370/A NAND2X1_LOC_318/A 0.00fF
C19465 NAND2X1_LOC_97/B NAND2X1_LOC_475/A 0.01fF
C19466 INVX1_LOC_617/Y NAND2X1_LOC_498/Y 0.01fF
C19467 INVX1_LOC_20/Y INVX1_LOC_288/A 0.07fF
C19468 INPUT_0 INVX1_LOC_375/Y 0.03fF
C19469 INVX1_LOC_613/Y INVX1_LOC_626/Y 0.09fF
C19470 INVX1_LOC_584/Y INVX1_LOC_522/Y 0.13fF
C19471 NAND2X1_LOC_797/a_36_24# INVX1_LOC_54/Y 0.00fF
C19472 INPUT_6 INVX1_LOC_25/Y 0.62fF
C19473 INVX1_LOC_626/Y NAND2X1_LOC_612/A 0.16fF
C19474 INVX1_LOC_501/Y INVX1_LOC_586/A 0.07fF
C19475 INVX1_LOC_362/Y INVX1_LOC_683/Y 0.07fF
C19476 INPUT_0 INVX1_LOC_600/Y 0.01fF
C19477 INVX1_LOC_20/Y INVX1_LOC_384/A 0.07fF
C19478 NAND2X1_LOC_516/Y INVX1_LOC_375/Y 0.01fF
C19479 INPUT_0 NAND2X1_LOC_61/a_36_24# 0.00fF
C19480 INPUT_6 NAND2X1_LOC_50/a_36_24# 0.00fF
C19481 NAND2X1_LOC_750/Y INVX1_LOC_178/A 0.08fF
C19482 INVX1_LOC_224/Y INVX1_LOC_230/A 0.02fF
C19483 NAND2X1_LOC_332/B INVX1_LOC_125/Y 0.01fF
C19484 INVX1_LOC_51/Y INVX1_LOC_367/A 0.02fF
C19485 NAND2X1_LOC_798/a_36_24# NAND2X1_LOC_173/Y 0.00fF
C19486 VDD INVX1_LOC_117/Y 4.47fF
C19487 INVX1_LOC_32/Y INVX1_LOC_388/Y 0.00fF
C19488 INVX1_LOC_193/Y INVX1_LOC_194/A 0.03fF
C19489 INVX1_LOC_395/A INVX1_LOC_189/Y 0.07fF
C19490 INVX1_LOC_617/Y INVX1_LOC_377/Y 0.22fF
C19491 INVX1_LOC_271/Y INVX1_LOC_155/Y 0.01fF
C19492 NAND2X1_LOC_707/A INVX1_LOC_358/Y 0.05fF
C19493 INVX1_LOC_54/Y NAND2X1_LOC_457/A 0.03fF
C19494 INVX1_LOC_133/Y INVX1_LOC_569/Y 0.15fF
C19495 NAND2X1_LOC_638/A INVX1_LOC_526/A 0.14fF
C19496 INVX1_LOC_51/Y INVX1_LOC_516/A 0.02fF
C19497 INVX1_LOC_468/Y INVX1_LOC_624/A 0.01fF
C19498 NAND2X1_LOC_122/Y INVX1_LOC_115/A 0.00fF
C19499 INVX1_LOC_45/A INVX1_LOC_333/A 0.02fF
C19500 INVX1_LOC_321/A INVX1_LOC_99/Y 0.01fF
C19501 INVX1_LOC_51/Y INVX1_LOC_669/Y 0.01fF
C19502 INVX1_LOC_33/Y INVX1_LOC_1/Y 0.10fF
C19503 INVX1_LOC_228/Y INVX1_LOC_117/Y 0.01fF
C19504 INVX1_LOC_560/A INVX1_LOC_361/Y 0.02fF
C19505 INVX1_LOC_20/Y INVX1_LOC_448/A 0.07fF
C19506 NAND2X1_LOC_284/a_36_24# INVX1_LOC_242/A 0.01fF
C19507 NAND2X1_LOC_179/Y INVX1_LOC_502/Y 0.02fF
C19508 INVX1_LOC_206/Y INVX1_LOC_100/A 0.33fF
C19509 INVX1_LOC_293/Y INVX1_LOC_679/Y 0.42fF
C19510 INVX1_LOC_537/Y INVX1_LOC_495/A 0.12fF
C19511 INVX1_LOC_50/Y NAND2X1_LOC_506/B 0.03fF
C19512 INVX1_LOC_395/A INVX1_LOC_31/Y 0.14fF
C19513 INVX1_LOC_21/A INVX1_LOC_9/A 0.01fF
C19514 INVX1_LOC_20/Y NAND2X1_LOC_791/A 0.02fF
C19515 INVX1_LOC_523/A INVX1_LOC_46/Y 0.02fF
C19516 NAND2X1_LOC_525/Y NAND2X1_LOC_184/Y 0.32fF
C19517 INVX1_LOC_31/A INVX1_LOC_53/A 0.02fF
C19518 INVX1_LOC_20/Y INVX1_LOC_145/Y 8.57fF
C19519 INVX1_LOC_45/Y INVX1_LOC_50/Y 0.79fF
C19520 INVX1_LOC_176/Y INVX1_LOC_99/Y 0.00fF
C19521 NAND2X1_LOC_387/Y INVX1_LOC_96/Y 0.31fF
C19522 INVX1_LOC_235/Y INVX1_LOC_367/Y 0.07fF
C19523 INVX1_LOC_290/Y NAND2X1_LOC_355/A 0.01fF
C19524 INVX1_LOC_134/Y INVX1_LOC_509/Y 0.06fF
C19525 INVX1_LOC_602/A INVX1_LOC_456/Y 0.05fF
C19526 NAND2X1_LOC_331/A INVX1_LOC_149/Y 0.01fF
C19527 NAND2X1_LOC_513/Y NAND2X1_LOC_308/A 0.00fF
C19528 INVX1_LOC_428/A NAND2X1_LOC_496/a_36_24# 0.00fF
C19529 INVX1_LOC_71/Y NAND2X1_LOC_66/Y 0.21fF
C19530 INVX1_LOC_51/A INVX1_LOC_58/Y 0.02fF
C19531 INVX1_LOC_72/Y INVX1_LOC_46/Y 0.02fF
C19532 INVX1_LOC_93/Y INVX1_LOC_51/Y 0.26fF
C19533 INVX1_LOC_53/Y INVX1_LOC_379/A 0.07fF
C19534 NAND2X1_LOC_241/B INVX1_LOC_58/Y 0.08fF
C19535 INVX1_LOC_312/Y INVX1_LOC_370/A 0.03fF
C19536 INVX1_LOC_606/Y INVX1_LOC_58/Y 0.01fF
C19537 INPUT_0 INVX1_LOC_494/Y 0.01fF
C19538 INVX1_LOC_348/A INVX1_LOC_50/Y 0.03fF
C19539 NAND2X1_LOC_534/Y INVX1_LOC_114/A 0.00fF
C19540 INVX1_LOC_53/Y INVX1_LOC_35/Y 2.35fF
C19541 INVX1_LOC_84/A NAND2X1_LOC_615/B 0.01fF
C19542 INVX1_LOC_286/Y INVX1_LOC_32/Y 0.01fF
C19543 INVX1_LOC_321/A INVX1_LOC_47/Y 0.03fF
C19544 INVX1_LOC_522/Y INVX1_LOC_186/Y 0.95fF
C19545 INPUT_3 INVX1_LOC_50/Y 0.15fF
C19546 INVX1_LOC_266/A INVX1_LOC_93/Y 0.10fF
C19547 INVX1_LOC_175/A INVX1_LOC_32/Y 0.04fF
C19548 INVX1_LOC_201/Y INVX1_LOC_600/A 0.00fF
C19549 NAND2X1_LOC_153/a_36_24# INVX1_LOC_508/A 0.00fF
C19550 INVX1_LOC_54/Y INVX1_LOC_651/A 0.00fF
C19551 INVX1_LOC_438/Y INVX1_LOC_430/A 0.06fF
C19552 INVX1_LOC_406/Y INVX1_LOC_421/A 0.00fF
C19553 NAND2X1_LOC_379/Y INVX1_LOC_48/Y 0.01fF
C19554 INVX1_LOC_20/Y NAND2X1_LOC_133/a_36_24# 0.00fF
C19555 INVX1_LOC_300/A INVX1_LOC_145/Y 0.07fF
C19556 NAND2X1_LOC_122/Y INVX1_LOC_49/Y 0.03fF
C19557 INVX1_LOC_134/Y INVX1_LOC_48/Y 0.22fF
C19558 INVX1_LOC_17/Y INVX1_LOC_7/Y 0.01fF
C19559 INVX1_LOC_444/Y INVX1_LOC_442/Y 0.07fF
C19560 INVX1_LOC_185/A INVX1_LOC_645/Y 0.00fF
C19561 INVX1_LOC_51/Y INVX1_LOC_675/A 0.07fF
C19562 INVX1_LOC_542/A INVX1_LOC_501/A 0.02fF
C19563 NAND2X1_LOC_782/A INVX1_LOC_581/A 0.04fF
C19564 INVX1_LOC_586/A INVX1_LOC_95/A 0.03fF
C19565 INVX1_LOC_193/A INVX1_LOC_12/Y 0.03fF
C19566 INVX1_LOC_419/Y INVX1_LOC_130/Y 0.23fF
C19567 INVX1_LOC_17/Y NAND2X1_LOC_259/A 0.03fF
C19568 INVX1_LOC_145/Y INVX1_LOC_197/Y 0.16fF
C19569 INVX1_LOC_202/Y INVX1_LOC_248/Y 0.03fF
C19570 INVX1_LOC_617/Y INVX1_LOC_47/Y 0.07fF
C19571 INVX1_LOC_20/Y INVX1_LOC_141/Y 0.01fF
C19572 NAND2X1_LOC_122/Y INVX1_LOC_533/A 0.24fF
C19573 INVX1_LOC_76/Y INVX1_LOC_507/A 0.01fF
C19574 INVX1_LOC_103/Y INVX1_LOC_104/Y 0.01fF
C19575 NAND2X1_LOC_790/B INVX1_LOC_91/Y 0.14fF
C19576 INVX1_LOC_453/A INVX1_LOC_450/Y 0.14fF
C19577 INVX1_LOC_78/A INVX1_LOC_61/A 0.27fF
C19578 INVX1_LOC_53/Y INVX1_LOC_620/A 0.03fF
C19579 NAND2X1_LOC_756/Y INVX1_LOC_284/Y 0.14fF
C19580 INVX1_LOC_595/Y INVX1_LOC_6/A 0.01fF
C19581 INVX1_LOC_84/A INVX1_LOC_296/A 0.03fF
C19582 INVX1_LOC_686/A INVX1_LOC_638/Y 0.09fF
C19583 INVX1_LOC_41/Y INVX1_LOC_215/Y 0.01fF
C19584 NAND2X1_LOC_41/Y INVX1_LOC_48/Y 0.04fF
C19585 INVX1_LOC_235/A INVX1_LOC_48/Y 0.02fF
C19586 INVX1_LOC_542/Y INVX1_LOC_676/A 0.19fF
C19587 INVX1_LOC_50/Y NAND2X1_LOC_69/Y 0.02fF
C19588 INVX1_LOC_452/A INVX1_LOC_444/A 0.14fF
C19589 NAND2X1_LOC_165/Y INVX1_LOC_59/Y 0.01fF
C19590 INVX1_LOC_17/Y INVX1_LOC_32/Y 8.47fF
C19591 INVX1_LOC_400/A INVX1_LOC_254/A 0.05fF
C19592 NAND2X1_LOC_491/a_36_24# INVX1_LOC_319/A 0.00fF
C19593 NAND2X1_LOC_324/B INVX1_LOC_376/A 0.17fF
C19594 INVX1_LOC_531/A INVX1_LOC_199/Y 0.04fF
C19595 NAND2X1_LOC_400/B INVX1_LOC_35/Y 0.12fF
C19596 INVX1_LOC_617/Y INVX1_LOC_119/Y 0.07fF
C19597 NAND2X1_LOC_755/B INVX1_LOC_659/A 0.07fF
C19598 INVX1_LOC_103/Y INVX1_LOC_117/Y 0.03fF
C19599 INVX1_LOC_492/A NAND2X1_LOC_647/A 0.00fF
C19600 INVX1_LOC_54/Y INVX1_LOC_87/Y 0.01fF
C19601 INVX1_LOC_176/Y NAND2X1_LOC_66/Y -0.01fF
C19602 NAND2X1_LOC_333/A INVX1_LOC_156/A 0.13fF
C19603 INVX1_LOC_343/Y INVX1_LOC_342/A 0.00fF
C19604 INVX1_LOC_89/Y INVX1_LOC_259/Y 0.06fF
C19605 INVX1_LOC_117/Y INVX1_LOC_68/A 0.03fF
C19606 INVX1_LOC_120/Y INVX1_LOC_230/A 0.01fF
C19607 INVX1_LOC_53/Y INVX1_LOC_518/Y 0.03fF
C19608 INVX1_LOC_169/A NAND2X1_LOC_489/a_36_24# 0.00fF
C19609 NAND2X1_LOC_837/A INVX1_LOC_50/Y 0.32fF
C19610 INVX1_LOC_6/Y INVX1_LOC_520/A 0.01fF
C19611 NAND2X1_LOC_184/Y INVX1_LOC_406/A 0.01fF
C19612 INVX1_LOC_65/A INVX1_LOC_48/Y 0.00fF
C19613 INVX1_LOC_137/Y INVX1_LOC_498/Y 0.46fF
C19614 INVX1_LOC_176/A INVX1_LOC_9/Y 0.07fF
C19615 INVX1_LOC_79/A INVX1_LOC_16/Y 0.01fF
C19616 INVX1_LOC_442/Y INVX1_LOC_26/Y 0.08fF
C19617 INVX1_LOC_501/A INVX1_LOC_259/Y 0.09fF
C19618 INVX1_LOC_145/Y INVX1_LOC_655/A 0.39fF
C19619 NAND2X1_LOC_692/Y INVX1_LOC_26/Y 0.16fF
C19620 INVX1_LOC_525/Y INVX1_LOC_96/A 0.07fF
C19621 INVX1_LOC_661/Y INVX1_LOC_655/A 0.18fF
C19622 INVX1_LOC_89/A INVX1_LOC_50/Y 0.01fF
C19623 INVX1_LOC_213/Y NAND2X1_LOC_258/a_36_24# 0.00fF
C19624 INVX1_LOC_80/Y INVX1_LOC_274/Y 0.02fF
C19625 INVX1_LOC_58/Y INVX1_LOC_341/Y 0.08fF
C19626 INVX1_LOC_242/Y INVX1_LOC_440/A 0.02fF
C19627 INVX1_LOC_100/Y INVX1_LOC_98/Y 0.19fF
C19628 INVX1_LOC_253/Y INVX1_LOC_69/Y 0.06fF
C19629 INVX1_LOC_338/Y INVX1_LOC_470/Y 0.01fF
C19630 INVX1_LOC_186/A INVX1_LOC_62/Y 0.02fF
C19631 NAND2X1_LOC_707/B INVX1_LOC_501/A 0.03fF
C19632 INVX1_LOC_578/Y INVX1_LOC_26/Y 0.03fF
C19633 INVX1_LOC_99/A INVX1_LOC_75/Y 0.03fF
C19634 INVX1_LOC_69/Y INVX1_LOC_63/Y 3.75fF
C19635 INVX1_LOC_211/A INVX1_LOC_600/Y 0.15fF
C19636 INVX1_LOC_25/A INVX1_LOC_1/Y 0.14fF
C19637 INVX1_LOC_353/A INVX1_LOC_260/Y 0.04fF
C19638 INVX1_LOC_166/A NAND2X1_LOC_274/B 2.88fF
C19639 INVX1_LOC_74/Y INVX1_LOC_98/Y 0.21fF
C19640 NAND2X1_LOC_274/B NAND2X1_LOC_849/a_36_24# 0.00fF
C19641 INVX1_LOC_349/A INVX1_LOC_62/Y 0.01fF
C19642 NAND2X1_LOC_531/Y INVX1_LOC_245/A 0.03fF
C19643 INVX1_LOC_513/Y INVX1_LOC_168/Y 0.14fF
C19644 INVX1_LOC_187/Y INVX1_LOC_245/A 0.01fF
C19645 NAND2X1_LOC_503/B NAND2X1_LOC_502/a_36_24# 0.02fF
C19646 INVX1_LOC_89/Y INVX1_LOC_114/A 0.01fF
C19647 INVX1_LOC_532/Y INVX1_LOC_26/Y 0.03fF
C19648 INVX1_LOC_261/Y INVX1_LOC_632/Y 0.03fF
C19649 INVX1_LOC_459/A INVX1_LOC_206/Y 0.02fF
C19650 VDD INVX1_LOC_448/Y 0.21fF
C19651 INVX1_LOC_77/A INVX1_LOC_351/A 0.01fF
C19652 INVX1_LOC_501/A INVX1_LOC_114/A 0.09fF
C19653 INVX1_LOC_77/A INVX1_LOC_90/Y 0.03fF
C19654 INVX1_LOC_58/Y INVX1_LOC_645/Y 0.01fF
C19655 INVX1_LOC_79/A INVX1_LOC_90/Y 0.09fF
C19656 INVX1_LOC_45/Y INVX1_LOC_275/A 0.02fF
C19657 INVX1_LOC_496/A NAND2X1_LOC_646/B 0.03fF
C19658 INVX1_LOC_340/Y INVX1_LOC_638/A 0.07fF
C19659 INVX1_LOC_206/Y INVX1_LOC_308/Y 0.01fF
C19660 INVX1_LOC_373/Y INVX1_LOC_479/A 0.02fF
C19661 INVX1_LOC_438/A INVX1_LOC_45/Y 0.07fF
C19662 NAND2X1_LOC_498/Y INVX1_LOC_410/Y 0.18fF
C19663 INVX1_LOC_443/A INVX1_LOC_245/A 2.82fF
C19664 NAND2X1_LOC_475/A INVX1_LOC_321/A 1.09fF
C19665 NAND2X1_LOC_498/Y INVX1_LOC_375/A 0.19fF
C19666 INVX1_LOC_614/A INVX1_LOC_185/A 0.02fF
C19667 INVX1_LOC_570/A INVX1_LOC_375/A 0.04fF
C19668 NAND2X1_LOC_498/Y INVX1_LOC_546/A 0.01fF
C19669 INVX1_LOC_409/Y INVX1_LOC_197/A 0.03fF
C19670 INVX1_LOC_395/A INVX1_LOC_51/Y 0.17fF
C19671 INVX1_LOC_152/Y NAND2X1_LOC_685/A 0.01fF
C19672 VDD INVX1_LOC_46/A 0.00fF
C19673 INVX1_LOC_601/A INVX1_LOC_619/A 0.37fF
C19674 VDD INVX1_LOC_658/A -0.00fF
C19675 INVX1_LOC_249/Y INVX1_LOC_250/A 0.01fF
C19676 NAND2X1_LOC_97/B NAND2X1_LOC_543/B 0.25fF
C19677 INVX1_LOC_417/A NAND2X1_LOC_543/B 0.01fF
C19678 INPUT_0 INVX1_LOC_401/A 0.01fF
C19679 INVX1_LOC_406/Y INVX1_LOC_445/Y 0.02fF
C19680 INVX1_LOC_362/Y INVX1_LOC_51/Y 0.07fF
C19681 INVX1_LOC_410/Y INVX1_LOC_377/Y 0.43fF
C19682 INVX1_LOC_266/A INVX1_LOC_395/A 0.05fF
C19683 VDD INVX1_LOC_281/Y 0.33fF
C19684 INVX1_LOC_521/Y INVX1_LOC_522/Y 0.05fF
C19685 INVX1_LOC_395/A INVX1_LOC_365/Y 0.03fF
C19686 INVX1_LOC_206/Y NAND2X1_LOC_237/Y 0.11fF
C19687 NAND2X1_LOC_249/Y NAND2X1_LOC_692/Y 0.09fF
C19688 VDD INVX1_LOC_251/Y 0.22fF
C19689 NAND2X1_LOC_377/a_36_24# INVX1_LOC_307/A 0.04fF
C19690 NAND2X1_LOC_513/Y INVX1_LOC_134/Y 0.46fF
C19691 INVX1_LOC_20/Y NAND2X1_LOC_332/B 0.06fF
C19692 NAND2X1_LOC_790/B NAND2X1_LOC_333/B 0.01fF
C19693 NAND2X1_LOC_475/A NAND2X1_LOC_366/a_36_24# 0.00fF
C19694 INVX1_LOC_51/Y INVX1_LOC_683/Y 0.02fF
C19695 NAND2X1_LOC_503/B NAND2X1_LOC_503/Y 0.02fF
C19696 VDD NAND2X1_LOC_76/A -0.00fF
C19697 INVX1_LOC_224/Y INVX1_LOC_681/A 0.01fF
C19698 NAND2X1_LOC_592/a_36_24# INVX1_LOC_31/Y 0.00fF
C19699 INVX1_LOC_617/Y INVX1_LOC_502/Y 0.24fF
C19700 INVX1_LOC_184/A INVX1_LOC_366/A 0.03fF
C19701 INVX1_LOC_410/Y INVX1_LOC_99/Y 0.03fF
C19702 NAND2X1_LOC_544/a_36_24# INVX1_LOC_53/Y 0.01fF
C19703 INVX1_LOC_185/Y NAND2X1_LOC_513/A 0.03fF
C19704 VDD INVX1_LOC_608/A 0.31fF
C19705 INVX1_LOC_228/Y INVX1_LOC_178/A 0.02fF
C19706 INVX1_LOC_122/Y INVX1_LOC_361/Y 0.03fF
C19707 INVX1_LOC_396/Y NAND2X1_LOC_237/Y 0.00fF
C19708 VDD INVX1_LOC_157/A 0.00fF
C19709 INVX1_LOC_248/Y INVX1_LOC_76/Y 0.03fF
C19710 INVX1_LOC_217/Y INVX1_LOC_387/Y 0.22fF
C19711 INVX1_LOC_510/Y INVX1_LOC_251/Y 0.01fF
C19712 NAND2X1_LOC_356/a_36_24# INVX1_LOC_259/Y 0.00fF
C19713 INVX1_LOC_570/A INVX1_LOC_61/A 0.03fF
C19714 VDD INVX1_LOC_58/Y 2.77fF
C19715 INVX1_LOC_555/Y INVX1_LOC_35/Y 0.02fF
C19716 INVX1_LOC_217/A INVX1_LOC_63/Y 0.01fF
C19717 INVX1_LOC_406/Y INVX1_LOC_99/Y 0.06fF
C19718 INVX1_LOC_197/A NAND2X1_LOC_302/A 0.01fF
C19719 INVX1_LOC_553/Y INVX1_LOC_47/Y 0.01fF
C19720 INVX1_LOC_410/Y INVX1_LOC_47/Y 0.03fF
C19721 INVX1_LOC_448/A INVX1_LOC_375/Y 0.03fF
C19722 NAND2X1_LOC_331/A INVX1_LOC_493/Y 0.15fF
C19723 INVX1_LOC_301/A INVX1_LOC_242/Y 0.08fF
C19724 NAND2X1_LOC_503/Y INVX1_LOC_273/A 0.02fF
C19725 INVX1_LOC_318/Y INVX1_LOC_59/Y 0.01fF
C19726 INVX1_LOC_228/Y INVX1_LOC_58/Y 0.03fF
C19727 INVX1_LOC_31/Y INVX1_LOC_51/Y 9.18fF
C19728 INVX1_LOC_546/A INVX1_LOC_47/Y 0.03fF
C19729 INVX1_LOC_363/Y INVX1_LOC_519/A 0.01fF
C19730 INVX1_LOC_65/Y INVX1_LOC_6/Y 0.00fF
C19731 INVX1_LOC_20/Y INVX1_LOC_598/A 0.08fF
C19732 INVX1_LOC_374/A INVX1_LOC_69/Y 0.03fF
C19733 NAND2X1_LOC_79/a_36_24# INVX1_LOC_198/A 0.00fF
C19734 INVX1_LOC_521/Y INVX1_LOC_508/A 0.00fF
C19735 INVX1_LOC_214/Y INVX1_LOC_53/Y 0.01fF
C19736 NAND2X1_LOC_148/A INVX1_LOC_35/Y 0.00fF
C19737 INVX1_LOC_586/A INVX1_LOC_253/Y 0.17fF
C19738 VDD NAND2X1_LOC_342/B 0.01fF
C19739 INVX1_LOC_145/Y INVX1_LOC_600/Y 0.03fF
C19740 INVX1_LOC_293/Y INVX1_LOC_50/Y 0.05fF
C19741 INVX1_LOC_318/Y INVX1_LOC_48/Y 0.00fF
C19742 INVX1_LOC_266/A INVX1_LOC_31/Y 0.01fF
C19743 INVX1_LOC_553/Y INVX1_LOC_119/Y 0.01fF
C19744 INVX1_LOC_442/Y NAND2X1_LOC_275/Y 0.00fF
C19745 INVX1_LOC_248/Y INVX1_LOC_559/A 0.01fF
C19746 INVX1_LOC_53/Y INVX1_LOC_118/A 0.01fF
C19747 INVX1_LOC_584/Y NAND2X1_LOC_467/a_36_24# 0.01fF
C19748 INVX1_LOC_510/Y INVX1_LOC_58/Y 0.06fF
C19749 INVX1_LOC_400/A NAND2X1_LOC_72/a_36_24# 0.00fF
C19750 INVX1_LOC_586/A INVX1_LOC_63/Y 0.15fF
C19751 INVX1_LOC_53/Y INVX1_LOC_649/A 0.04fF
C19752 INVX1_LOC_410/Y INVX1_LOC_119/Y 0.14fF
C19753 NAND2X1_LOC_679/B NAND2X1_LOC_407/a_36_24# 0.00fF
C19754 INPUT_0 NAND2X1_LOC_123/B 0.03fF
C19755 INVX1_LOC_605/Y INVX1_LOC_523/Y 0.04fF
C19756 INVX1_LOC_663/Y NAND2X1_LOC_260/Y 0.01fF
C19757 INVX1_LOC_447/Y INVX1_LOC_303/Y 0.17fF
C19758 INVX1_LOC_322/Y INVX1_LOC_328/Y 0.19fF
C19759 INVX1_LOC_61/A INVX1_LOC_99/Y 0.10fF
C19760 INVX1_LOC_546/A INVX1_LOC_119/Y 0.03fF
C19761 INVX1_LOC_7/Y INVX1_LOC_198/A 0.03fF
C19762 NAND2X1_LOC_271/B INVX1_LOC_280/A 0.06fF
C19763 INVX1_LOC_435/Y INVX1_LOC_100/Y 0.05fF
C19764 INVX1_LOC_440/A INVX1_LOC_197/Y 0.08fF
C19765 INVX1_LOC_674/A INVX1_LOC_99/Y 0.07fF
C19766 INVX1_LOC_193/Y INVX1_LOC_62/Y 0.00fF
C19767 INVX1_LOC_196/A INVX1_LOC_496/A 0.04fF
C19768 INVX1_LOC_173/Y INVX1_LOC_600/A 0.02fF
C19769 NAND2X1_LOC_13/Y INVX1_LOC_390/A 0.07fF
C19770 INVX1_LOC_613/Y INVX1_LOC_627/Y 0.03fF
C19771 INVX1_LOC_576/Y INVX1_LOC_47/Y 0.01fF
C19772 INVX1_LOC_584/A INVX1_LOC_479/A 0.02fF
C19773 INVX1_LOC_69/Y INVX1_LOC_387/A 0.03fF
C19774 INVX1_LOC_312/Y INVX1_LOC_63/Y 0.09fF
C19775 NAND2X1_LOC_76/a_36_24# INVX1_LOC_41/Y 0.01fF
C19776 INVX1_LOC_685/A INVX1_LOC_641/Y 0.14fF
C19777 INVX1_LOC_49/Y INVX1_LOC_519/A 0.03fF
C19778 INVX1_LOC_614/A INVX1_LOC_58/Y 0.05fF
C19779 INVX1_LOC_20/Y INVX1_LOC_242/Y 0.07fF
C19780 NAND2X1_LOC_673/B INVX1_LOC_50/Y 0.01fF
C19781 INVX1_LOC_140/Y INVX1_LOC_588/A 0.04fF
C19782 NAND2X1_LOC_372/a_36_24# INVX1_LOC_100/Y 0.01fF
C19783 INVX1_LOC_369/A INVX1_LOC_482/Y 0.00fF
C19784 INVX1_LOC_536/A INVX1_LOC_499/A -0.00fF
C19785 NAND2X1_LOC_334/a_36_24# INVX1_LOC_49/Y 0.01fF
C19786 INVX1_LOC_213/Y NAND2X1_LOC_253/Y 0.09fF
C19787 INPUT_0 INVX1_LOC_485/A 0.01fF
C19788 INVX1_LOC_596/A INVX1_LOC_100/Y 0.03fF
C19789 INVX1_LOC_63/Y NAND2X1_LOC_378/Y 0.03fF
C19790 NAND2X1_LOC_698/Y INVX1_LOC_35/Y 0.02fF
C19791 INVX1_LOC_58/Y INVX1_LOC_684/A 0.13fF
C19792 INVX1_LOC_400/A INVX1_LOC_361/A 0.02fF
C19793 INVX1_LOC_466/A INVX1_LOC_463/Y 0.12fF
C19794 INVX1_LOC_63/Y NAND2X1_LOC_202/a_36_24# 0.00fF
C19795 INVX1_LOC_6/Y INVX1_LOC_385/A 0.05fF
C19796 NAND2X1_LOC_843/A INVX1_LOC_58/Y 0.32fF
C19797 INPUT_0 INVX1_LOC_92/A 0.07fF
C19798 INVX1_LOC_54/Y INVX1_LOC_306/Y 0.01fF
C19799 NAND2X1_LOC_311/a_36_24# INVX1_LOC_75/Y 0.00fF
C19800 INVX1_LOC_59/Y INVX1_LOC_351/A 0.00fF
C19801 NAND2X1_LOC_260/Y INVX1_LOC_655/A 0.22fF
C19802 NAND2X1_LOC_141/a_36_24# INVX1_LOC_670/A 0.00fF
C19803 INVX1_LOC_662/A INVX1_LOC_35/Y 0.03fF
C19804 NAND2X1_LOC_318/B INVX1_LOC_100/Y 0.00fF
C19805 INVX1_LOC_658/A INVX1_LOC_635/Y 0.01fF
C19806 INVX1_LOC_290/A INVX1_LOC_632/Y 0.00fF
C19807 INVX1_LOC_242/Y INVX1_LOC_197/Y 0.07fF
C19808 INVX1_LOC_77/A INVX1_LOC_98/Y 0.03fF
C19809 INVX1_LOC_682/A INVX1_LOC_681/Y 0.00fF
C19810 INVX1_LOC_276/Y INVX1_LOC_221/Y 0.29fF
C19811 NAND2X1_LOC_786/B INVX1_LOC_178/A 0.23fF
C19812 INVX1_LOC_351/A INVX1_LOC_48/Y 0.08fF
C19813 INVX1_LOC_93/Y NAND2X1_LOC_668/Y 0.01fF
C19814 NAND2X1_LOC_532/Y INVX1_LOC_66/A 0.11fF
C19815 NAND2X1_LOC_123/A NAND2X1_LOC_123/B 0.00fF
C19816 INVX1_LOC_59/Y INVX1_LOC_90/Y 1.65fF
C19817 INVX1_LOC_54/Y INVX1_LOC_9/Y 0.10fF
C19818 INVX1_LOC_620/A NAND2X1_LOC_790/a_36_24# 0.03fF
C19819 INVX1_LOC_440/Y INVX1_LOC_353/A 0.03fF
C19820 INVX1_LOC_79/A INVX1_LOC_98/Y 0.08fF
C19821 INVX1_LOC_381/A NAND2X1_LOC_416/B 0.01fF
C19822 INVX1_LOC_261/A INVX1_LOC_673/Y 0.01fF
C19823 INVX1_LOC_48/Y INVX1_LOC_90/Y 0.20fF
C19824 INVX1_LOC_314/Y INVX1_LOC_6/Y 0.01fF
C19825 INVX1_LOC_382/A INVX1_LOC_245/A 0.26fF
C19826 INVX1_LOC_537/A INVX1_LOC_479/A 0.17fF
C19827 INVX1_LOC_504/A INVX1_LOC_74/Y 0.01fF
C19828 INVX1_LOC_125/A INVX1_LOC_479/A 0.01fF
C19829 INVX1_LOC_357/A NAND2X1_LOC_451/B 0.04fF
C19830 INVX1_LOC_525/Y INVX1_LOC_353/A 0.05fF
C19831 INVX1_LOC_416/A INVX1_LOC_75/Y 0.05fF
C19832 INVX1_LOC_419/Y INVX1_LOC_75/Y 0.02fF
C19833 INVX1_LOC_54/Y INVX1_LOC_62/Y 0.21fF
C19834 NAND2X1_LOC_334/B NAND2X1_LOC_668/Y 0.10fF
C19835 INVX1_LOC_6/Y INVX1_LOC_244/Y 0.14fF
C19836 NAND2X1_LOC_636/A NAND2X1_LOC_583/a_36_24# 0.02fF
C19837 INVX1_LOC_54/Y INVX1_LOC_13/Y 0.00fF
C19838 INVX1_LOC_490/A INVX1_LOC_280/A 0.12fF
C19839 INVX1_LOC_41/Y INVX1_LOC_463/Y 0.03fF
C19840 INVX1_LOC_69/Y INVX1_LOC_454/Y 0.06fF
C19841 INVX1_LOC_79/A INVX1_LOC_338/Y 0.08fF
C19842 INVX1_LOC_479/A INVX1_LOC_496/Y 0.02fF
C19843 INVX1_LOC_301/Y NAND2X1_LOC_274/B 0.12fF
C19844 INVX1_LOC_663/A INVX1_LOC_664/A 0.04fF
C19845 NAND2X1_LOC_543/B INVX1_LOC_412/Y 0.03fF
C19846 INVX1_LOC_521/A INVX1_LOC_62/Y 0.01fF
C19847 INVX1_LOC_461/Y INVX1_LOC_114/A 0.01fF
C19848 NAND2X1_LOC_274/B INVX1_LOC_41/Y 0.03fF
C19849 INVX1_LOC_446/A INVX1_LOC_586/A 0.01fF
C19850 NAND2X1_LOC_475/A INVX1_LOC_410/Y 0.03fF
C19851 INVX1_LOC_114/A INVX1_LOC_347/A 0.00fF
C19852 INVX1_LOC_269/Y NAND2X1_LOC_76/B 0.15fF
C19853 INVX1_LOC_502/A INVX1_LOC_75/Y 0.07fF
C19854 INVX1_LOC_20/Y NAND2X1_LOC_7/Y 0.01fF
C19855 INVX1_LOC_182/A NAND2X1_LOC_750/Y 0.02fF
C19856 NAND2X1_LOC_373/Y NAND2X1_LOC_332/B 0.15fF
C19857 NAND2X1_LOC_249/Y NAND2X1_LOC_128/a_36_24# 0.01fF
C19858 INVX1_LOC_148/Y INVX1_LOC_41/Y 0.00fF
C19859 INVX1_LOC_100/Y NAND2X1_LOC_411/a_36_24# 0.01fF
C19860 INVX1_LOC_594/Y INVX1_LOC_677/Y 0.11fF
C19861 INVX1_LOC_206/Y INVX1_LOC_666/A 0.02fF
C19862 INVX1_LOC_433/Y INVX1_LOC_424/Y 0.01fF
C19863 INVX1_LOC_362/Y INVX1_LOC_216/Y 0.07fF
C19864 INVX1_LOC_295/Y INVX1_LOC_109/Y 0.05fF
C19865 INVX1_LOC_438/A INVX1_LOC_293/Y 0.02fF
C19866 INVX1_LOC_62/Y NAND2X1_LOC_609/a_36_24# 0.00fF
C19867 INVX1_LOC_502/A NAND2X1_LOC_271/A 0.19fF
C19868 INVX1_LOC_414/A NAND2X1_LOC_523/B 0.47fF
C19869 INVX1_LOC_74/Y INVX1_LOC_346/Y 0.00fF
C19870 NAND2X1_LOC_97/B NAND2X1_LOC_335/B 0.02fF
C19871 INVX1_LOC_449/A NAND2X1_LOC_184/a_36_24# -0.02fF
C19872 INVX1_LOC_542/A NAND2X1_LOC_685/B 0.02fF
C19873 INVX1_LOC_512/Y INVX1_LOC_499/Y 0.96fF
C19874 NAND2X1_LOC_336/B INVX1_LOC_560/A 0.06fF
C19875 INVX1_LOC_206/Y NAND2X1_LOC_325/B 0.07fF
C19876 INVX1_LOC_131/Y INVX1_LOC_133/A 0.00fF
C19877 INVX1_LOC_374/A NAND2X1_LOC_440/a_36_24# 0.00fF
C19878 VDD INVX1_LOC_1/Y 0.61fF
C19879 INVX1_LOC_412/Y INVX1_LOC_469/A 0.01fF
C19880 INVX1_LOC_206/Y NAND2X1_LOC_72/Y 0.09fF
C19881 INVX1_LOC_602/A INVX1_LOC_45/Y 0.03fF
C19882 INVX1_LOC_400/Y INVX1_LOC_12/Y 0.05fF
C19883 INVX1_LOC_442/Y INVX1_LOC_103/A 0.01fF
C19884 INVX1_LOC_274/A INVX1_LOC_97/A 0.09fF
C19885 INVX1_LOC_578/A INVX1_LOC_99/A 0.10fF
C19886 INVX1_LOC_617/A INVX1_LOC_617/Y 0.01fF
C19887 INVX1_LOC_397/A NAND2X1_LOC_237/Y 0.05fF
C19888 INVX1_LOC_390/Y INVX1_LOC_230/A 0.05fF
C19889 INVX1_LOC_45/Y INVX1_LOC_104/Y 0.01fF
C19890 NAND2X1_LOC_736/a_36_24# NAND2X1_LOC_122/Y 0.00fF
C19891 INVX1_LOC_31/A INVX1_LOC_602/A 0.02fF
C19892 INVX1_LOC_68/Y NAND2X1_LOC_97/B 0.00fF
C19893 INVX1_LOC_405/A INVX1_LOC_69/Y 0.05fF
C19894 VDD NAND2X1_LOC_689/B 0.18fF
C19895 INVX1_LOC_380/A INVX1_LOC_328/Y 0.00fF
C19896 INVX1_LOC_85/Y INVX1_LOC_43/Y 0.00fF
C19897 INVX1_LOC_11/Y NAND2X1_LOC_710/a_36_24# 0.00fF
C19898 INVX1_LOC_22/Y INPUT_2 0.01fF
C19899 NAND2X1_LOC_140/B NAND2X1_LOC_332/B 0.57fF
C19900 INPUT_0 INPUT_1 1.55fF
C19901 INVX1_LOC_465/Y NAND2X1_LOC_334/A 0.03fF
C19902 INVX1_LOC_140/Y NAND2X1_LOC_646/A 0.01fF
C19903 NAND2X1_LOC_788/A NAND2X1_LOC_532/Y 0.03fF
C19904 INVX1_LOC_583/A INVX1_LOC_522/Y 0.02fF
C19905 INVX1_LOC_402/Y INVX1_LOC_551/Y 0.17fF
C19906 NAND2X1_LOC_97/A INVX1_LOC_202/Y 0.02fF
C19907 INVX1_LOC_193/A INVX1_LOC_442/A 0.32fF
C19908 NAND2X1_LOC_516/Y INPUT_1 0.05fF
C19909 INVX1_LOC_20/Y INVX1_LOC_300/A 1.10fF
C19910 INVX1_LOC_575/A NAND2X1_LOC_152/Y 0.00fF
C19911 INVX1_LOC_172/A INVX1_LOC_322/Y 0.35fF
C19912 INVX1_LOC_31/Y INVX1_LOC_355/A 0.01fF
C19913 INVX1_LOC_417/Y NAND2X1_LOC_545/B 0.12fF
C19914 INVX1_LOC_117/Y INVX1_LOC_45/Y 0.31fF
C19915 INVX1_LOC_206/Y INVX1_LOC_351/Y 0.01fF
C19916 NAND2X1_LOC_720/a_36_24# INVX1_LOC_53/Y 0.01fF
C19917 INVX1_LOC_20/Y INVX1_LOC_197/Y 0.17fF
C19918 INVX1_LOC_408/Y NAND2X1_LOC_532/Y 0.03fF
C19919 INVX1_LOC_366/A INVX1_LOC_623/Y 0.01fF
C19920 INVX1_LOC_616/A INVX1_LOC_198/A 0.02fF
C19921 INVX1_LOC_202/A INVX1_LOC_90/Y 0.02fF
C19922 INVX1_LOC_395/A INVX1_LOC_380/Y 0.05fF
C19923 INVX1_LOC_366/A INVX1_LOC_86/Y 0.04fF
C19924 GATE_579 INVX1_LOC_671/A 0.45fF
C19925 NAND2X1_LOC_122/Y INVX1_LOC_32/Y 0.03fF
C19926 NAND2X1_LOC_373/Y INVX1_LOC_242/Y 0.02fF
C19927 INVX1_LOC_206/Y INVX1_LOC_168/Y 0.09fF
C19928 VDD INVX1_LOC_245/A 1.75fF
C19929 INVX1_LOC_294/A INVX1_LOC_381/A 0.04fF
C19930 INVX1_LOC_576/A INVX1_LOC_300/A 0.03fF
C19931 INVX1_LOC_273/A INVX1_LOC_32/Y 0.01fF
C19932 INVX1_LOC_395/A NAND2X1_LOC_668/Y 0.04fF
C19933 INVX1_LOC_17/Y NAND2X1_LOC_299/Y 0.01fF
C19934 INVX1_LOC_140/Y INVX1_LOC_63/Y 0.03fF
C19935 INVX1_LOC_607/Y INVX1_LOC_679/Y 0.60fF
C19936 INVX1_LOC_68/Y INVX1_LOC_525/Y 0.20fF
C19937 NAND2X1_LOC_391/B INVX1_LOC_46/Y 0.02fF
C19938 INVX1_LOC_100/Y NAND2X1_LOC_76/B 2.01fF
C19939 NAND2X1_LOC_393/Y INVX1_LOC_7/Y 0.07fF
C19940 INPUT_3 INVX1_LOC_117/Y 0.03fF
C19941 INVX1_LOC_272/Y INVX1_LOC_623/Y 0.00fF
C19942 NAND2X1_LOC_13/Y INVX1_LOC_31/Y 0.03fF
C19943 INVX1_LOC_250/Y INVX1_LOC_440/Y 0.09fF
C19944 INVX1_LOC_228/Y INVX1_LOC_245/A 0.29fF
C19945 INVX1_LOC_417/Y INVX1_LOC_98/Y 0.03fF
C19946 INVX1_LOC_523/A NAND2X1_LOC_816/a_36_24# 0.00fF
C19947 INVX1_LOC_451/A INVX1_LOC_385/Y 0.15fF
C19948 NAND2X1_LOC_184/Y NAND2X1_LOC_840/a_36_24# 0.00fF
C19949 INPUT_0 INVX1_LOC_487/Y 0.02fF
C19950 INVX1_LOC_300/A INVX1_LOC_197/Y 0.07fF
C19951 INVX1_LOC_74/Y NAND2X1_LOC_76/B 0.07fF
C19952 INVX1_LOC_613/Y INVX1_LOC_612/Y 0.19fF
C19953 INVX1_LOC_257/Y NAND2X1_LOC_123/B 0.14fF
C19954 INVX1_LOC_59/Y INVX1_LOC_98/Y 0.02fF
C19955 NAND2X1_LOC_45/Y NAND2X1_LOC_528/Y 0.10fF
C19956 INVX1_LOC_376/Y INVX1_LOC_624/A 0.01fF
C19957 INVX1_LOC_597/A INVX1_LOC_623/Y 0.01fF
C19958 NAND2X1_LOC_355/a_36_24# INVX1_LOC_259/Y 0.00fF
C19959 NAND2X1_LOC_400/B INVX1_LOC_324/A 0.02fF
C19960 INVX1_LOC_291/A NAND2X1_LOC_790/a_36_24# 0.00fF
C19961 INVX1_LOC_435/Y INVX1_LOC_79/A 0.12fF
C19962 INVX1_LOC_230/A INVX1_LOC_432/A 0.04fF
C19963 INVX1_LOC_591/Y INVX1_LOC_69/Y 0.02fF
C19964 INVX1_LOC_193/A INVX1_LOC_116/Y 0.02fF
C19965 NAND2X1_LOC_779/a_36_24# NAND2X1_LOC_708/A 0.01fF
C19966 INVX1_LOC_213/Y INVX1_LOC_214/Y 0.02fF
C19967 INVX1_LOC_358/Y INVX1_LOC_463/Y -0.00fF
C19968 INVX1_LOC_32/Y NAND2X1_LOC_393/Y 0.00fF
C19969 INVX1_LOC_48/Y INVX1_LOC_98/Y 1.70fF
C19970 INVX1_LOC_607/Y INPUT_1 0.09fF
C19971 INVX1_LOC_166/A NAND2X1_LOC_595/Y 0.34fF
C19972 NAND2X1_LOC_534/a_36_24# INVX1_LOC_49/Y 0.01fF
C19973 NAND2X1_LOC_791/B INVX1_LOC_63/Y 0.04fF
C19974 INVX1_LOC_272/Y INVX1_LOC_63/Y 0.03fF
C19975 INVX1_LOC_17/Y NAND2X1_LOC_184/Y 0.19fF
C19976 INVX1_LOC_361/Y NAND2X1_LOC_307/a_36_24# 0.00fF
C19977 INVX1_LOC_132/Y INVX1_LOC_655/A 0.01fF
C19978 INPUT_5 NAND2X1_LOC_53/a_36_24# 0.00fF
C19979 NAND2X1_LOC_190/A INVX1_LOC_54/Y 0.02fF
C19980 INVX1_LOC_160/A NAND2X1_LOC_388/A 0.00fF
C19981 INVX1_LOC_632/A INVX1_LOC_497/A 0.14fF
C19982 INVX1_LOC_629/A INVX1_LOC_346/Y 0.00fF
C19983 INVX1_LOC_347/Y INVX1_LOC_633/Y 0.00fF
C19984 INVX1_LOC_20/Y NAND2X1_LOC_447/a_36_24# 0.00fF
C19985 INVX1_LOC_53/Y INVX1_LOC_507/Y 0.17fF
C19986 INVX1_LOC_20/Y INVX1_LOC_655/A 0.09fF
C19987 NAND2X1_LOC_498/Y INVX1_LOC_479/A 0.09fF
C19988 INVX1_LOC_570/A INVX1_LOC_479/A 0.07fF
C19989 INVX1_LOC_254/Y INVX1_LOC_123/A 0.02fF
C19990 NAND2X1_LOC_847/a_36_24# INVX1_LOC_655/A 0.01fF
C19991 INVX1_LOC_54/Y INVX1_LOC_87/A 0.05fF
C19992 INVX1_LOC_366/A NAND2X1_LOC_214/a_36_24# 0.01fF
C19993 INVX1_LOC_596/A INVX1_LOC_79/A 0.02fF
C19994 INVX1_LOC_63/Y INVX1_LOC_252/A 0.00fF
C19995 INVX1_LOC_429/Y INVX1_LOC_443/A 0.09fF
C19996 INVX1_LOC_257/Y INVX1_LOC_92/A 0.01fF
C19997 INVX1_LOC_6/Y INVX1_LOC_623/Y 0.01fF
C19998 INVX1_LOC_17/Y INVX1_LOC_551/A -0.06fF
C19999 NAND2X1_LOC_294/Y INVX1_LOC_385/A 0.16fF
C20000 INVX1_LOC_6/Y INVX1_LOC_86/Y 0.03fF
C20001 INVX1_LOC_418/Y INVX1_LOC_411/Y 0.00fF
C20002 INVX1_LOC_21/Y NAND2X1_LOC_274/B 0.09fF
C20003 INVX1_LOC_201/A INVX1_LOC_399/A 0.09fF
C20004 INVX1_LOC_298/A INVX1_LOC_292/Y 0.01fF
C20005 INVX1_LOC_159/Y INVX1_LOC_411/Y 0.00fF
C20006 INVX1_LOC_530/A INVX1_LOC_100/Y 0.02fF
C20007 INVX1_LOC_402/A INVX1_LOC_518/Y 0.04fF
C20008 INVX1_LOC_49/Y INVX1_LOC_513/A 0.03fF
C20009 INVX1_LOC_572/Y INVX1_LOC_542/Y 0.09fF
C20010 INVX1_LOC_338/Y INVX1_LOC_48/Y 0.12fF
C20011 INVX1_LOC_54/Y INVX1_LOC_624/Y 0.02fF
C20012 INVX1_LOC_240/A NAND2X1_LOC_342/A 0.01fF
C20013 INVX1_LOC_504/A INVX1_LOC_79/A 0.46fF
C20014 INVX1_LOC_625/A INVX1_LOC_100/Y 0.02fF
C20015 INVX1_LOC_31/Y NAND2X1_LOC_668/Y 0.01fF
C20016 INVX1_LOC_7/Y NAND2X1_LOC_416/a_36_24# 0.01fF
C20017 NAND2X1_LOC_677/Y INVX1_LOC_62/Y 0.00fF
C20018 INVX1_LOC_117/Y INVX1_LOC_89/A 0.02fF
C20019 INVX1_LOC_93/Y INVX1_LOC_480/A 0.02fF
C20020 INVX1_LOC_31/Y INVX1_LOC_361/A 0.00fF
C20021 NAND2X1_LOC_253/Y NAND2X1_LOC_258/Y 0.45fF
C20022 INVX1_LOC_501/A INVX1_LOC_539/Y 0.01fF
C20023 INVX1_LOC_675/A INVX1_LOC_359/A 0.04fF
C20024 INVX1_LOC_261/Y NAND2X1_LOC_586/Y 0.00fF
C20025 INVX1_LOC_662/A INVX1_LOC_649/A 0.15fF
C20026 NAND2X1_LOC_274/B NAND2X1_LOC_274/a_36_24# 0.00fF
C20027 INVX1_LOC_63/Y INVX1_LOC_6/Y 4.46fF
C20028 NAND2X1_LOC_404/a_36_24# INVX1_LOC_9/Y 0.01fF
C20029 INVX1_LOC_48/Y NAND2X1_LOC_41/a_36_24# 0.01fF
C20030 INVX1_LOC_161/A INVX1_LOC_588/A 0.00fF
C20031 INVX1_LOC_402/Y NAND2X1_LOC_410/Y 0.00fF
C20032 INVX1_LOC_69/Y INVX1_LOC_674/Y 0.03fF
C20033 INVX1_LOC_199/A INVX1_LOC_9/Y 0.01fF
C20034 INVX1_LOC_35/Y NAND2X1_LOC_625/a_36_24# 0.01fF
C20035 INVX1_LOC_479/A INVX1_LOC_99/Y 0.09fF
C20036 INVX1_LOC_89/Y INVX1_LOC_9/Y 10.14fF
C20037 INVX1_LOC_418/Y INVX1_LOC_41/Y 0.08fF
C20038 INVX1_LOC_17/Y INVX1_LOC_75/Y 0.09fF
C20039 INVX1_LOC_93/Y NAND2X1_LOC_301/B 0.12fF
C20040 NAND2X1_LOC_451/a_36_24# INVX1_LOC_74/Y 0.00fF
C20041 INVX1_LOC_628/A INVX1_LOC_346/Y 0.03fF
C20042 INVX1_LOC_304/A INVX1_LOC_666/Y 0.03fF
C20043 INVX1_LOC_244/Y NAND2X1_LOC_294/Y 0.00fF
C20044 INVX1_LOC_63/Y NAND2X1_LOC_437/a_36_24# 0.01fF
C20045 INVX1_LOC_166/A NAND2X1_LOC_372/Y 0.05fF
C20046 INVX1_LOC_63/Y NAND2X1_LOC_81/Y 0.17fF
C20047 INVX1_LOC_116/Y NAND2X1_LOC_457/a_36_24# -0.00fF
C20048 INVX1_LOC_100/Y NAND2X1_LOC_52/Y 0.01fF
C20049 INVX1_LOC_339/Y INVX1_LOC_245/A 0.04fF
C20050 INVX1_LOC_89/Y INVX1_LOC_62/Y 0.39fF
C20051 INVX1_LOC_338/Y INVX1_LOC_472/Y 0.04fF
C20052 NAND2X1_LOC_615/Y INVX1_LOC_90/Y 0.02fF
C20053 NAND2X1_LOC_603/a_36_24# INVX1_LOC_634/Y 0.00fF
C20054 INVX1_LOC_469/Y INVX1_LOC_346/Y 0.22fF
C20055 INVX1_LOC_409/Y INVX1_LOC_412/Y 0.26fF
C20056 INVX1_LOC_47/Y INVX1_LOC_479/A 0.16fF
C20057 INVX1_LOC_93/Y INVX1_LOC_291/Y 0.01fF
C20058 INVX1_LOC_150/A NAND2X1_LOC_161/a_36_24# 0.02fF
C20059 INVX1_LOC_501/A INVX1_LOC_62/Y 0.03fF
C20060 NAND2X1_LOC_249/Y INVX1_LOC_215/Y 0.01fF
C20061 NAND2X1_LOC_192/A INVX1_LOC_588/A 0.01fF
C20062 INVX1_LOC_405/A INVX1_LOC_586/A 0.04fF
C20063 INVX1_LOC_182/A VDD 0.19fF
C20064 INVX1_LOC_152/Y INVX1_LOC_542/A 0.01fF
C20065 INVX1_LOC_479/A INVX1_LOC_119/Y 0.05fF
C20066 INVX1_LOC_560/Y INVX1_LOC_586/A 0.03fF
C20067 INVX1_LOC_601/A NAND2X1_LOC_773/A 0.00fF
C20068 INVX1_LOC_446/A INVX1_LOC_486/Y 0.07fF
C20069 INVX1_LOC_79/A INVX1_LOC_346/Y 0.07fF
C20070 INVX1_LOC_20/Y NAND2X1_LOC_310/a_36_24# 0.00fF
C20071 INVX1_LOC_373/A NAND2X1_LOC_707/A 0.02fF
C20072 INVX1_LOC_20/Y INVX1_LOC_553/A 0.01fF
C20073 INVX1_LOC_460/A INVX1_LOC_346/Y 0.00fF
C20074 INVX1_LOC_301/A NAND2X1_LOC_524/a_36_24# 0.00fF
C20075 NAND2X1_LOC_631/B NAND2X1_LOC_416/B 0.18fF
C20076 VDD INVX1_LOC_599/A -0.00fF
C20077 INVX1_LOC_84/A NAND2X1_LOC_537/B 0.01fF
C20078 NAND2X1_LOC_231/B INVX1_LOC_91/A 0.18fF
C20079 INVX1_LOC_224/Y NAND2X1_LOC_307/A 0.02fF
C20080 NAND2X1_LOC_97/A INVX1_LOC_98/A 0.23fF
C20081 NAND2X1_LOC_685/B INVX1_LOC_499/Y 0.00fF
C20082 NAND2X1_LOC_61/A INVX1_LOC_178/A 0.02fF
C20083 NAND2X1_LOC_45/Y INVX1_LOC_12/Y 1.83fF
C20084 INVX1_LOC_395/A NAND2X1_LOC_152/B 0.02fF
C20085 INVX1_LOC_213/Y INVX1_LOC_220/A 0.02fF
C20086 NAND2X1_LOC_704/a_36_24# INVX1_LOC_53/Y 0.01fF
C20087 INVX1_LOC_558/A NAND2X1_LOC_516/B 0.05fF
C20088 NAND2X1_LOC_97/A INVX1_LOC_76/Y 0.01fF
C20089 NAND2X1_LOC_370/a_36_24# INVX1_LOC_98/Y 0.00fF
C20090 INVX1_LOC_578/A NAND2X1_LOC_307/A 0.07fF
C20091 INVX1_LOC_556/A INVX1_LOC_80/A 0.76fF
C20092 NAND2X1_LOC_163/B NAND2X1_LOC_467/A 0.03fF
C20093 INVX1_LOC_206/Y INVX1_LOC_99/A 0.05fF
C20094 INVX1_LOC_557/A NAND2X1_LOC_307/A 0.06fF
C20095 INVX1_LOC_412/Y NAND2X1_LOC_369/a_36_24# 0.00fF
C20096 INVX1_LOC_557/A INVX1_LOC_545/Y 0.22fF
C20097 INVX1_LOC_354/Y INVX1_LOC_638/A 0.03fF
C20098 INVX1_LOC_84/A INVX1_LOC_586/A 0.11fF
C20099 INVX1_LOC_190/Y INVX1_LOC_7/Y 0.01fF
C20100 INVX1_LOC_165/Y INVX1_LOC_633/Y 0.10fF
C20101 VDD INVX1_LOC_218/Y 0.21fF
C20102 INVX1_LOC_31/A NAND2X1_LOC_22/a_36_24# 0.02fF
C20103 INVX1_LOC_133/Y GATE_662 0.38fF
C20104 NAND2X1_LOC_39/Y INVX1_LOC_76/Y 0.01fF
C20105 NAND2X1_LOC_554/a_36_24# INVX1_LOC_608/A -0.00fF
C20106 NAND2X1_LOC_23/a_36_24# INVX1_LOC_11/Y 0.00fF
C20107 INVX1_LOC_490/Y INVX1_LOC_379/A 0.03fF
C20108 INVX1_LOC_254/Y NAND2X1_LOC_475/A 0.07fF
C20109 INVX1_LOC_434/A INVX1_LOC_439/Y 0.03fF
C20110 INVX1_LOC_312/Y NAND2X1_LOC_620/a_36_24# 0.00fF
C20111 NAND2X1_LOC_513/Y INVX1_LOC_98/Y 0.10fF
C20112 INVX1_LOC_608/Y INVX1_LOC_607/A 0.01fF
C20113 INVX1_LOC_402/Y INVX1_LOC_558/A 0.03fF
C20114 INVX1_LOC_551/Y INVX1_LOC_367/A 0.03fF
C20115 NAND2X1_LOC_180/B INVX1_LOC_80/A 0.00fF
C20116 INVX1_LOC_45/Y INVX1_LOC_281/Y 0.09fF
C20117 INVX1_LOC_257/Y INPUT_1 0.07fF
C20118 NAND2X1_LOC_331/A NAND2X1_LOC_187/Y 0.10fF
C20119 INVX1_LOC_413/Y INVX1_LOC_367/Y 0.08fF
C20120 INVX1_LOC_72/Y INVX1_LOC_7/Y 0.05fF
C20121 INVX1_LOC_133/Y NAND2X1_LOC_846/B 0.18fF
C20122 INVX1_LOC_11/Y INVX1_LOC_556/A 0.00fF
C20123 NAND2X1_LOC_750/Y INVX1_LOC_543/Y 0.05fF
C20124 INVX1_LOC_21/Y INVX1_LOC_38/A 0.01fF
C20125 INPUT_3 INVX1_LOC_46/A 0.07fF
C20126 INVX1_LOC_416/A INVX1_LOC_578/A 0.05fF
C20127 INPUT_0 INVX1_LOC_50/Y 0.20fF
C20128 INVX1_LOC_419/Y INVX1_LOC_578/A 0.59fF
C20129 INVX1_LOC_129/A INVX1_LOC_586/A 0.01fF
C20130 INVX1_LOC_53/Y INVX1_LOC_522/Y 0.34fF
C20131 INVX1_LOC_45/Y INVX1_LOC_178/A 0.00fF
C20132 INVX1_LOC_601/A NAND2X1_LOC_240/A 0.04fF
C20133 INVX1_LOC_203/Y INVX1_LOC_155/A 0.00fF
C20134 VDD INVX1_LOC_639/A 0.00fF
C20135 INVX1_LOC_435/Y INVX1_LOC_48/Y 0.03fF
C20136 INVX1_LOC_20/Y NAND2X1_LOC_140/B 0.56fF
C20137 INVX1_LOC_273/A NAND2X1_LOC_226/Y 0.01fF
C20138 INVX1_LOC_400/Y NAND2X1_LOC_615/B 0.08fF
C20139 INVX1_LOC_293/Y INVX1_LOC_104/Y 0.10fF
C20140 VDD INVX1_LOC_520/Y 0.08fF
C20141 INVX1_LOC_17/Y NAND2X1_LOC_486/B 0.17fF
C20142 NAND2X1_LOC_516/Y INVX1_LOC_50/Y 0.05fF
C20143 INVX1_LOC_143/Y INVX1_LOC_137/Y 0.01fF
C20144 INPUT_0 INVX1_LOC_431/Y 0.01fF
C20145 INVX1_LOC_579/A NAND2X1_LOC_736/a_36_24# 0.02fF
C20146 INPUT_3 INVX1_LOC_281/Y 0.01fF
C20147 INVX1_LOC_80/A INVX1_LOC_188/Y 0.03fF
C20148 NAND2X1_LOC_13/Y NAND2X1_LOC_267/a_36_24# 0.00fF
C20149 INVX1_LOC_99/A INVX1_LOC_686/A 0.57fF
C20150 VDD INVX1_LOC_386/A 0.00fF
C20151 INVX1_LOC_603/Y INVX1_LOC_80/A 0.56fF
C20152 INVX1_LOC_45/Y INVX1_LOC_608/A 0.04fF
C20153 INVX1_LOC_372/Y INVX1_LOC_99/Y 0.07fF
C20154 INVX1_LOC_298/Y INVX1_LOC_59/A 0.01fF
C20155 INVX1_LOC_400/A INVX1_LOC_551/Y 0.02fF
C20156 INVX1_LOC_255/Y INVX1_LOC_372/A 0.08fF
C20157 INVX1_LOC_561/Y INVX1_LOC_497/A 0.00fF
C20158 INVX1_LOC_468/Y NAND2X1_LOC_307/A 0.03fF
C20159 INVX1_LOC_384/A INPUT_1 0.10fF
C20160 INVX1_LOC_468/Y INVX1_LOC_545/Y 0.18fF
C20161 NAND2X1_LOC_635/B INVX1_LOC_677/Y 0.20fF
C20162 INVX1_LOC_323/Y NAND2X1_LOC_399/B 0.10fF
C20163 INVX1_LOC_77/A NAND2X1_LOC_76/B 0.01fF
C20164 NAND2X1_LOC_416/Y INVX1_LOC_489/Y 0.01fF
C20165 NAND2X1_LOC_152/Y INVX1_LOC_575/Y 0.01fF
C20166 INVX1_LOC_12/Y INVX1_LOC_99/Y 0.11fF
C20167 INVX1_LOC_323/Y INVX1_LOC_7/Y 0.03fF
C20168 INVX1_LOC_679/Y INVX1_LOC_145/Y 0.32fF
C20169 NAND2X1_LOC_513/Y INVX1_LOC_338/Y 0.01fF
C20170 NAND2X1_LOC_523/a_36_24# INVX1_LOC_362/Y 0.00fF
C20171 INVX1_LOC_173/A INVX1_LOC_199/Y 0.05fF
C20172 INVX1_LOC_80/A INVX1_LOC_478/Y 0.06fF
C20173 INVX1_LOC_35/Y INVX1_LOC_97/Y 0.00fF
C20174 INVX1_LOC_551/Y INVX1_LOC_93/Y 0.10fF
C20175 INVX1_LOC_596/A INVX1_LOC_48/Y 0.02fF
C20176 INVX1_LOC_609/Y INVX1_LOC_137/Y 0.01fF
C20177 INVX1_LOC_45/Y INVX1_LOC_58/Y 0.43fF
C20178 INVX1_LOC_659/Y INVX1_LOC_673/Y 0.96fF
C20179 INVX1_LOC_686/A INVX1_LOC_355/Y 0.01fF
C20180 NAND2X1_LOC_387/Y INVX1_LOC_80/A 0.07fF
C20181 NAND2X1_LOC_638/A INVX1_LOC_674/A 0.07fF
C20182 INVX1_LOC_374/A NAND2X1_LOC_437/a_36_24# 0.00fF
C20183 INVX1_LOC_586/A INVX1_LOC_674/Y 0.01fF
C20184 INVX1_LOC_137/Y INVX1_LOC_14/A 0.07fF
C20185 NAND2X1_LOC_69/Y INVX1_LOC_178/A 0.12fF
C20186 INVX1_LOC_435/A INVX1_LOC_211/Y 0.01fF
C20187 INVX1_LOC_448/A INPUT_1 0.08fF
C20188 INVX1_LOC_578/A INVX1_LOC_502/A 0.22fF
C20189 INVX1_LOC_681/Y INVX1_LOC_145/Y 0.02fF
C20190 INVX1_LOC_476/A INVX1_LOC_508/Y 0.00fF
C20191 INVX1_LOC_534/Y INVX1_LOC_512/Y 0.02fF
C20192 NAND2X1_LOC_596/Y NAND2X1_LOC_597/Y 0.04fF
C20193 INVX1_LOC_372/Y INVX1_LOC_47/Y 0.04fF
C20194 INVX1_LOC_504/A INVX1_LOC_48/Y 0.44fF
C20195 INVX1_LOC_323/Y INVX1_LOC_32/Y 0.02fF
C20196 INVX1_LOC_123/A INVX1_LOC_12/Y 0.03fF
C20197 NAND2X1_LOC_475/A INVX1_LOC_479/A 0.08fF
C20198 INVX1_LOC_431/A INVX1_LOC_35/Y 0.01fF
C20199 INVX1_LOC_145/Y INPUT_1 0.03fF
C20200 INVX1_LOC_65/Y INVX1_LOC_100/Y 0.03fF
C20201 INVX1_LOC_12/Y INVX1_LOC_47/Y 0.39fF
C20202 INVX1_LOC_267/A NAND2X1_LOC_755/B 0.01fF
C20203 NAND2X1_LOC_333/A INVX1_LOC_99/Y 0.03fF
C20204 NAND2X1_LOC_521/Y INVX1_LOC_99/Y 0.00fF
C20205 INVX1_LOC_53/Y INVX1_LOC_508/A 0.39fF
C20206 NAND2X1_LOC_517/Y INVX1_LOC_63/Y 0.06fF
C20207 NAND2X1_LOC_325/B NAND2X1_LOC_542/A 0.03fF
C20208 INVX1_LOC_12/Y NAND2X1_LOC_557/B 0.13fF
C20209 INVX1_LOC_527/Y INVX1_LOC_50/Y 0.00fF
C20210 INVX1_LOC_78/A INVX1_LOC_66/A 0.01fF
C20211 INVX1_LOC_117/Y NAND2X1_LOC_673/B 0.23fF
C20212 INVX1_LOC_35/Y INVX1_LOC_18/Y 0.20fF
C20213 INVX1_LOC_302/A NAND2X1_LOC_372/Y 0.04fF
C20214 NAND2X1_LOC_32/Y INVX1_LOC_86/Y 0.04fF
C20215 INVX1_LOC_99/Y INVX1_LOC_188/A 0.16fF
C20216 INVX1_LOC_65/Y INVX1_LOC_74/Y 0.03fF
C20217 INVX1_LOC_85/Y INVX1_LOC_190/A 0.10fF
C20218 INVX1_LOC_298/A INVX1_LOC_50/Y 0.03fF
C20219 INVX1_LOC_145/A INVX1_LOC_1/Y 0.01fF
C20220 INVX1_LOC_170/A INVX1_LOC_99/Y 0.00fF
C20221 INVX1_LOC_395/A INVX1_LOC_291/Y 0.03fF
C20222 INVX1_LOC_372/Y INVX1_LOC_119/Y 0.03fF
C20223 INVX1_LOC_167/A INVX1_LOC_93/Y 0.05fF
C20224 INVX1_LOC_94/Y INVX1_LOC_35/Y 0.04fF
C20225 INVX1_LOC_492/A NAND2X1_LOC_307/B 0.28fF
C20226 INVX1_LOC_58/Y NAND2X1_LOC_69/Y 0.01fF
C20227 NAND2X1_LOC_775/B INVX1_LOC_199/Y 0.03fF
C20228 GATE_865 INVX1_LOC_69/Y 0.03fF
C20229 INVX1_LOC_301/Y NAND2X1_LOC_595/Y 0.00fF
C20230 INVX1_LOC_416/A INVX1_LOC_120/Y 0.00fF
C20231 INVX1_LOC_193/A INVX1_LOC_69/Y 0.00fF
C20232 INVX1_LOC_69/Y INVX1_LOC_156/A 0.03fF
C20233 INVX1_LOC_12/Y NAND2X1_LOC_66/Y 0.03fF
C20234 NAND2X1_LOC_820/A INVX1_LOC_669/A 0.04fF
C20235 INVX1_LOC_415/Y INVX1_LOC_63/Y 0.03fF
C20236 INVX1_LOC_69/Y NAND2X1_LOC_822/Y 0.02fF
C20237 INVX1_LOC_155/Y INVX1_LOC_90/Y 0.02fF
C20238 INVX1_LOC_31/Y NAND2X1_LOC_449/B 0.01fF
C20239 INVX1_LOC_49/Y INVX1_LOC_670/A 0.02fF
C20240 INVX1_LOC_194/Y INVX1_LOC_9/Y 0.00fF
C20241 INVX1_LOC_625/A INVX1_LOC_79/A 0.00fF
C20242 INVX1_LOC_384/Y INVX1_LOC_443/A 0.21fF
C20243 INVX1_LOC_80/A INVX1_LOC_91/A 0.01fF
C20244 NAND2X1_LOC_836/B INVX1_LOC_6/Y 0.07fF
C20245 NAND2X1_LOC_595/Y INVX1_LOC_41/Y 0.03fF
C20246 INVX1_LOC_100/Y INVX1_LOC_370/A 0.01fF
C20247 INVX1_LOC_171/A INVX1_LOC_245/A 0.18fF
C20248 INVX1_LOC_35/Y NAND2X1_LOC_489/A 0.04fF
C20249 INPUT_5 INVX1_LOC_342/A 0.03fF
C20250 INVX1_LOC_89/Y INVX1_LOC_624/Y 0.10fF
C20251 INVX1_LOC_21/Y INVX1_LOC_39/Y 0.01fF
C20252 INVX1_LOC_145/Y NAND2X1_LOC_827/a_36_24# 0.00fF
C20253 INVX1_LOC_166/A INVX1_LOC_518/A 0.07fF
C20254 INVX1_LOC_338/A INVX1_LOC_653/Y 0.01fF
C20255 INVX1_LOC_41/Y INVX1_LOC_352/Y 0.00fF
C20256 NAND2X1_LOC_527/Y INVX1_LOC_502/A 0.02fF
C20257 INVX1_LOC_62/Y INVX1_LOC_194/Y 0.03fF
C20258 INVX1_LOC_133/Y INVX1_LOC_554/A 0.00fF
C20259 INVX1_LOC_208/Y INVX1_LOC_79/A 0.07fF
C20260 INVX1_LOC_318/A INVX1_LOC_100/Y 0.03fF
C20261 INVX1_LOC_280/Y INVX1_LOC_369/Y 0.04fF
C20262 INVX1_LOC_58/Y INVX1_LOC_89/A 0.16fF
C20263 INVX1_LOC_26/Y INVX1_LOC_372/A 0.01fF
C20264 INVX1_LOC_479/Y INVX1_LOC_74/Y 0.01fF
C20265 INVX1_LOC_63/Y INVX1_LOC_206/A 0.02fF
C20266 INVX1_LOC_11/Y INVX1_LOC_91/A 0.00fF
C20267 INVX1_LOC_285/Y INVX1_LOC_44/Y 0.06fF
C20268 INVX1_LOC_17/Y NAND2X1_LOC_619/a_36_24# 0.00fF
C20269 INVX1_LOC_89/A NAND2X1_LOC_90/a_36_24# 0.02fF
C20270 INVX1_LOC_397/Y INVX1_LOC_100/Y 0.09fF
C20271 INVX1_LOC_318/A INVX1_LOC_74/Y 0.08fF
C20272 INVX1_LOC_170/A NAND2X1_LOC_66/Y 0.00fF
C20273 INVX1_LOC_75/Y INVX1_LOC_230/Y 0.15fF
C20274 INVX1_LOC_241/A INVX1_LOC_46/Y 0.00fF
C20275 INVX1_LOC_662/A INVX1_LOC_667/Y -0.03fF
C20276 INVX1_LOC_298/A INVX1_LOC_658/Y 0.35fF
C20277 INVX1_LOC_470/Y INVX1_LOC_588/A 0.01fF
C20278 INPUT_0 INVX1_LOC_275/A 0.09fF
C20279 NAND2X1_LOC_686/A INVX1_LOC_79/A 0.01fF
C20280 NAND2X1_LOC_613/Y INVX1_LOC_109/Y 0.04fF
C20281 NAND2X1_LOC_274/B INVX1_LOC_26/Y 0.03fF
C20282 NAND2X1_LOC_274/B INVX1_LOC_128/Y 0.01fF
C20283 INPUT_0 INVX1_LOC_438/A 0.07fF
C20284 NAND2X1_LOC_242/A NAND2X1_LOC_164/Y 0.01fF
C20285 VDD INVX1_LOC_429/Y 0.21fF
C20286 NAND2X1_LOC_231/A NAND2X1_LOC_790/B 0.01fF
C20287 INPUT_0 INVX1_LOC_24/A 0.01fF
C20288 INVX1_LOC_62/Y INVX1_LOC_461/Y 0.15fF
C20289 NAND2X1_LOC_555/B INVX1_LOC_443/A 0.03fF
C20290 INVX1_LOC_41/Y INVX1_LOC_280/A 0.03fF
C20291 NAND2X1_LOC_636/A INVX1_LOC_168/A 0.06fF
C20292 INVX1_LOC_41/Y NAND2X1_LOC_372/Y 0.02fF
C20293 INVX1_LOC_26/Y NAND2X1_LOC_242/a_36_24# 0.00fF
C20294 INVX1_LOC_554/A INVX1_LOC_337/Y 0.01fF
C20295 INVX1_LOC_257/Y INVX1_LOC_134/A 0.00fF
C20296 NAND2X1_LOC_331/A INVX1_LOC_150/Y 0.15fF
C20297 INVX1_LOC_400/Y INVX1_LOC_442/A 0.07fF
C20298 INVX1_LOC_107/A NAND2X1_LOC_142/Y 0.01fF
C20299 INVX1_LOC_74/Y INVX1_LOC_588/A -0.00fF
C20300 INVX1_LOC_242/Y INVX1_LOC_92/A 0.22fF
C20301 INVX1_LOC_317/Y INVX1_LOC_266/Y 0.10fF
C20302 INVX1_LOC_395/A INVX1_LOC_551/Y 0.10fF
C20303 INVX1_LOC_206/Y NAND2X1_LOC_307/A 0.43fF
C20304 INVX1_LOC_174/Y INVX1_LOC_586/A 0.08fF
C20305 INVX1_LOC_584/Y NAND2X1_LOC_467/A 0.60fF
C20306 NAND2X1_LOC_332/a_36_24# NAND2X1_LOC_325/B 0.01fF
C20307 INVX1_LOC_145/Y INVX1_LOC_181/A 0.01fF
C20308 NAND2X1_LOC_475/A INVX1_LOC_12/Y 0.05fF
C20309 INVX1_LOC_409/A INVX1_LOC_21/Y 0.06fF
C20310 INPUT_0 NAND2X1_LOC_513/A 0.71fF
C20311 NAND2X1_LOC_242/A INVX1_LOC_604/Y 0.10fF
C20312 VDD INVX1_LOC_201/Y 0.21fF
C20313 INVX1_LOC_666/A NAND2X1_LOC_845/a_36_24# 0.02fF
C20314 NAND2X1_LOC_391/B INVX1_LOC_76/Y 0.01fF
C20315 INVX1_LOC_59/Y NAND2X1_LOC_76/B 0.11fF
C20316 NAND2X1_LOC_261/Y INVX1_LOC_384/Y 0.05fF
C20317 INVX1_LOC_233/Y INVX1_LOC_406/Y 0.01fF
C20318 INVX1_LOC_558/A INVX1_LOC_367/A 0.52fF
C20319 NAND2X1_LOC_789/B INVX1_LOC_145/Y 0.02fF
C20320 INVX1_LOC_224/Y INVX1_LOC_17/Y 0.21fF
C20321 INVX1_LOC_269/A INVX1_LOC_80/A 0.07fF
C20322 NAND2X1_LOC_173/a_36_24# INVX1_LOC_638/A 0.00fF
C20323 INVX1_LOC_182/A INVX1_LOC_619/A 0.02fF
C20324 NAND2X1_LOC_56/a_36_24# INVX1_LOC_400/Y -0.00fF
C20325 NAND2X1_LOC_45/Y INVX1_LOC_159/A 0.11fF
C20326 INVX1_LOC_48/Y NAND2X1_LOC_76/B 2.08fF
C20327 NAND2X1_LOC_312/a_36_24# INVX1_LOC_98/Y 0.00fF
C20328 INVX1_LOC_421/Y INVX1_LOC_99/Y 0.14fF
C20329 NAND2X1_LOC_299/Y NAND2X1_LOC_122/Y 0.03fF
C20330 INVX1_LOC_133/Y INVX1_LOC_199/Y 0.00fF
C20331 INVX1_LOC_419/Y INVX1_LOC_206/Y 0.01fF
C20332 VDD INVX1_LOC_543/Y 0.28fF
C20333 INVX1_LOC_400/Y INVX1_LOC_116/Y 0.07fF
C20334 VDD INVX1_LOC_686/Y 0.21fF
C20335 INVX1_LOC_17/Y INVX1_LOC_578/A 0.16fF
C20336 INVX1_LOC_437/A INVX1_LOC_445/Y 0.03fF
C20337 NAND2X1_LOC_258/Y INVX1_LOC_220/A 0.08fF
C20338 NAND2X1_LOC_332/B INVX1_LOC_679/Y 0.33fF
C20339 NAND2X1_LOC_511/a_36_24# INVX1_LOC_99/Y 0.00fF
C20340 INVX1_LOC_591/Y NAND2X1_LOC_791/B 0.04fF
C20341 INVX1_LOC_166/A NAND2X1_LOC_317/A 0.01fF
C20342 NAND2X1_LOC_523/B NAND2X1_LOC_541/B 0.01fF
C20343 NAND2X1_LOC_307/A INVX1_LOC_686/A 0.07fF
C20344 INVX1_LOC_545/Y INVX1_LOC_686/A -0.00fF
C20345 INVX1_LOC_30/Y INPUT_4 0.01fF
C20346 NAND2X1_LOC_45/Y INVX1_LOC_66/A 0.00fF
C20347 NAND2X1_LOC_710/a_36_24# INVX1_LOC_361/Y 0.00fF
C20348 NAND2X1_LOC_148/a_36_24# INVX1_LOC_133/A 0.00fF
C20349 NAND2X1_LOC_140/a_36_24# INVX1_LOC_670/A 0.00fF
C20350 INVX1_LOC_31/A INVX1_LOC_1/Y 0.01fF
C20351 NAND2X1_LOC_475/A INVX1_LOC_188/A 0.02fF
C20352 INVX1_LOC_288/A INVX1_LOC_50/Y 0.07fF
C20353 INVX1_LOC_586/A GATE_865 0.03fF
C20354 NAND2X1_LOC_755/B INVX1_LOC_59/A 0.84fF
C20355 INVX1_LOC_293/Y INVX1_LOC_281/Y 0.00fF
C20356 INVX1_LOC_524/Y NAND2X1_LOC_755/B 0.00fF
C20357 INVX1_LOC_53/Y NAND2X1_LOC_496/Y 0.35fF
C20358 NAND2X1_LOC_317/B INVX1_LOC_199/Y 0.42fF
C20359 INVX1_LOC_166/A INVX1_LOC_165/Y 0.01fF
C20360 INVX1_LOC_193/A INVX1_LOC_586/A 0.00fF
C20361 NAND2X1_LOC_566/a_36_24# INVX1_LOC_197/Y 0.01fF
C20362 INVX1_LOC_295/A INVX1_LOC_681/A 0.04fF
C20363 INVX1_LOC_558/A INVX1_LOC_93/Y 0.15fF
C20364 NAND2X1_LOC_498/Y INVX1_LOC_66/A 0.14fF
C20365 NAND2X1_LOC_332/B INPUT_1 0.06fF
C20366 INVX1_LOC_206/Y INVX1_LOC_376/A 0.07fF
C20367 NAND2X1_LOC_142/Y NAND2X1_LOC_285/A 0.00fF
C20368 INVX1_LOC_395/A INVX1_LOC_486/A 0.09fF
C20369 INVX1_LOC_45/Y NAND2X1_LOC_689/B 0.01fF
C20370 NAND2X1_LOC_320/Y INVX1_LOC_633/Y 0.02fF
C20371 INVX1_LOC_384/A INVX1_LOC_50/Y 0.09fF
C20372 INVX1_LOC_570/A INVX1_LOC_66/A 0.03fF
C20373 NAND2X1_LOC_714/a_36_24# INVX1_LOC_89/Y 0.01fF
C20374 INVX1_LOC_416/A INVX1_LOC_686/A 0.20fF
C20375 INVX1_LOC_80/A INVX1_LOC_504/Y 0.35fF
C20376 INVX1_LOC_419/Y INVX1_LOC_686/A 0.00fF
C20377 NAND2X1_LOC_325/B NAND2X1_LOC_323/a_36_24# 0.02fF
C20378 INVX1_LOC_118/Y INVX1_LOC_9/Y 0.03fF
C20379 INVX1_LOC_53/Y NAND2X1_LOC_775/B 0.07fF
C20380 INVX1_LOC_551/Y INVX1_LOC_31/Y 0.03fF
C20381 INVX1_LOC_125/Y INPUT_1 0.02fF
C20382 INVX1_LOC_269/Y INVX1_LOC_63/Y 0.18fF
C20383 INVX1_LOC_293/Y INVX1_LOC_608/A 0.03fF
C20384 INPUT_6 INVX1_LOC_25/A 0.34fF
C20385 INVX1_LOC_625/A INVX1_LOC_398/Y 0.04fF
C20386 INVX1_LOC_21/Y INVX1_LOC_352/Y 0.03fF
C20387 INVX1_LOC_625/A INVX1_LOC_59/Y 0.02fF
C20388 VDD INVX1_LOC_657/Y 0.26fF
C20389 INVX1_LOC_53/A INVX1_LOC_145/Y 0.13fF
C20390 NAND2X1_LOC_164/Y INVX1_LOC_79/A 0.09fF
C20391 INVX1_LOC_455/Y INVX1_LOC_315/A 0.06fF
C20392 NAND2X1_LOC_705/a_36_24# INVX1_LOC_69/Y 0.00fF
C20393 VDD INVX1_LOC_652/Y 0.36fF
C20394 INVX1_LOC_84/A INVX1_LOC_6/Y 0.16fF
C20395 NAND2X1_LOC_41/Y INVX1_LOC_176/A 0.03fF
C20396 INVX1_LOC_169/A INVX1_LOC_199/Y 0.00fF
C20397 INVX1_LOC_448/A INVX1_LOC_50/Y 0.01fF
C20398 VDD INVX1_LOC_483/A -0.00fF
C20399 INVX1_LOC_678/A INVX1_LOC_684/A 0.04fF
C20400 NAND2X1_LOC_682/a_36_24# INVX1_LOC_498/Y 0.00fF
C20401 INVX1_LOC_45/Y INVX1_LOC_245/A 0.61fF
C20402 NAND2X1_LOC_13/Y INVX1_LOC_361/A 0.06fF
C20403 INVX1_LOC_381/A INVX1_LOC_63/Y 0.07fF
C20404 INVX1_LOC_447/Y INVX1_LOC_665/Y 0.02fF
C20405 INVX1_LOC_99/Y NAND2X1_LOC_615/B 0.03fF
C20406 INVX1_LOC_199/Y INVX1_LOC_337/Y 0.00fF
C20407 NAND2X1_LOC_673/B INVX1_LOC_178/A 0.04fF
C20408 NAND2X1_LOC_756/Y INVX1_LOC_58/Y 0.02fF
C20409 INVX1_LOC_625/A INVX1_LOC_48/Y 0.01fF
C20410 NAND2X1_LOC_697/Y INVX1_LOC_54/Y 0.02fF
C20411 NAND2X1_LOC_45/Y NAND2X1_LOC_621/B 0.14fF
C20412 INVX1_LOC_145/Y INVX1_LOC_50/Y 14.02fF
C20413 INVX1_LOC_65/Y INVX1_LOC_79/A 0.16fF
C20414 INVX1_LOC_293/Y INVX1_LOC_58/Y 0.03fF
C20415 INVX1_LOC_35/Y NAND2X1_LOC_84/B 0.85fF
C20416 INVX1_LOC_93/Y NAND2X1_LOC_755/B 2.01fF
C20417 NAND2X1_LOC_498/Y NAND2X1_LOC_601/Y 0.02fF
C20418 INVX1_LOC_382/A NAND2X1_LOC_416/Y 0.01fF
C20419 INVX1_LOC_51/Y NAND2X1_LOC_301/B 0.08fF
C20420 INVX1_LOC_584/Y INVX1_LOC_41/Y 0.02fF
C20421 NAND2X1_LOC_513/A INVX1_LOC_476/Y 0.17fF
C20422 INVX1_LOC_516/A INVX1_LOC_46/Y 0.00fF
C20423 INVX1_LOC_166/A INVX1_LOC_352/A 0.02fF
C20424 INPUT_1 INVX1_LOC_503/Y 0.01fF
C20425 NAND2X1_LOC_712/a_36_24# INVX1_LOC_48/Y 0.00fF
C20426 INVX1_LOC_53/Y NAND2X1_LOC_283/a_36_24# 0.00fF
C20427 INVX1_LOC_599/Y INVX1_LOC_204/Y 0.16fF
C20428 INVX1_LOC_99/Y INVX1_LOC_66/A 0.01fF
C20429 INVX1_LOC_145/Y INVX1_LOC_431/Y 0.09fF
C20430 INPUT_3 INVX1_LOC_245/A 0.07fF
C20431 INVX1_LOC_266/Y INVX1_LOC_531/Y 0.07fF
C20432 INVX1_LOC_99/A NAND2X1_LOC_542/A 0.27fF
C20433 INVX1_LOC_301/A INVX1_LOC_92/A 0.47fF
C20434 INVX1_LOC_345/Y INVX1_LOC_513/A 0.01fF
C20435 INVX1_LOC_288/Y INVX1_LOC_261/Y 0.25fF
C20436 INVX1_LOC_84/A NAND2X1_LOC_81/Y 0.05fF
C20437 NAND2X1_LOC_391/A INVX1_LOC_9/Y 0.03fF
C20438 INVX1_LOC_402/Y INVX1_LOC_49/Y 0.02fF
C20439 INVX1_LOC_160/A INVX1_LOC_58/Y 0.03fF
C20440 INVX1_LOC_87/A INVX1_LOC_194/Y 0.05fF
C20441 INVX1_LOC_32/Y INVX1_LOC_513/A 0.03fF
C20442 NAND2X1_LOC_789/A INVX1_LOC_86/Y 0.01fF
C20443 INVX1_LOC_166/A INVX1_LOC_105/Y 0.00fF
C20444 INVX1_LOC_300/A NAND2X1_LOC_666/Y 0.03fF
C20445 INVX1_LOC_17/Y GATE_479 0.04fF
C20446 NAND2X1_LOC_545/a_36_24# NAND2X1_LOC_775/B 0.01fF
C20447 INVX1_LOC_27/Y INVX1_LOC_9/Y 0.18fF
C20448 INVX1_LOC_598/A INVX1_LOC_292/Y 0.00fF
C20449 INVX1_LOC_93/Y INVX1_LOC_46/Y 0.25fF
C20450 NAND2X1_LOC_755/B NAND2X1_LOC_334/B 0.02fF
C20451 NAND2X1_LOC_673/B INVX1_LOC_58/Y 0.10fF
C20452 NAND2X1_LOC_770/B INVX1_LOC_69/Y 0.02fF
C20453 INVX1_LOC_20/Y INVX1_LOC_329/Y 0.01fF
C20454 INVX1_LOC_183/Y NAND2X1_LOC_81/a_36_24# 0.00fF
C20455 INVX1_LOC_604/Y INVX1_LOC_79/A 0.19fF
C20456 INVX1_LOC_312/A INVX1_LOC_62/Y 0.00fF
C20457 INVX1_LOC_188/Y NAND2X1_LOC_432/a_36_24# 0.01fF
C20458 INVX1_LOC_127/Y INVX1_LOC_47/Y 0.02fF
C20459 NAND2X1_LOC_391/A INVX1_LOC_62/Y 0.03fF
C20460 INVX1_LOC_449/A INVX1_LOC_41/Y 0.08fF
C20461 INVX1_LOC_183/A INVX1_LOC_83/Y 0.00fF
C20462 INVX1_LOC_201/Y NAND2X1_LOC_786/B 0.02fF
C20463 INVX1_LOC_444/Y INVX1_LOC_405/Y 0.05fF
C20464 INVX1_LOC_317/A INVX1_LOC_199/Y 0.01fF
C20465 INVX1_LOC_47/Y INVX1_LOC_66/A 0.07fF
C20466 NAND2X1_LOC_647/A NAND2X1_LOC_612/a_36_24# 0.02fF
C20467 INVX1_LOC_147/A INVX1_LOC_62/Y 0.37fF
C20468 INVX1_LOC_324/A INVX1_LOC_327/A 0.01fF
C20469 INVX1_LOC_267/A INVX1_LOC_49/Y 0.01fF
C20470 INVX1_LOC_21/Y INVX1_LOC_280/A 0.02fF
C20471 INVX1_LOC_20/Y INVX1_LOC_270/Y 0.01fF
C20472 INVX1_LOC_44/Y INVX1_LOC_87/A 0.03fF
C20473 INVX1_LOC_47/Y INVX1_LOC_296/A 0.01fF
C20474 INVX1_LOC_133/A INVX1_LOC_240/Y 0.01fF
C20475 NAND2X1_LOC_250/Y INVX1_LOC_100/Y 0.34fF
C20476 NAND2X1_LOC_545/A INVX1_LOC_350/A 0.04fF
C20477 INPUT_1 INVX1_LOC_242/Y 0.01fF
C20478 INVX1_LOC_602/A INVX1_LOC_622/Y 0.01fF
C20479 INVX1_LOC_117/Y INVX1_LOC_117/A 0.01fF
C20480 INVX1_LOC_13/Y INVX1_LOC_27/Y 0.13fF
C20481 INVX1_LOC_523/Y INVX1_LOC_9/Y 0.08fF
C20482 INVX1_LOC_543/Y NAND2X1_LOC_786/B 0.03fF
C20483 NAND2X1_LOC_198/a_36_24# INVX1_LOC_223/Y 0.00fF
C20484 INVX1_LOC_20/Y INVX1_LOC_92/A 1.22fF
C20485 INVX1_LOC_139/Y INVX1_LOC_168/Y 0.05fF
C20486 INVX1_LOC_652/Y INVX1_LOC_509/A 0.11fF
C20487 INVX1_LOC_444/Y INVX1_LOC_450/Y 0.11fF
C20488 INPUT_1 INVX1_LOC_487/A 0.00fF
C20489 INVX1_LOC_479/A INVX1_LOC_505/A 0.03fF
C20490 INVX1_LOC_119/Y INVX1_LOC_66/A 0.03fF
C20491 INVX1_LOC_145/Y INVX1_LOC_658/Y 0.02fF
C20492 INVX1_LOC_253/Y INVX1_LOC_100/Y 0.05fF
C20493 INVX1_LOC_300/A INVX1_LOC_270/Y 0.02fF
C20494 VDD INVX1_LOC_458/Y 0.26fF
C20495 INVX1_LOC_63/Y INVX1_LOC_100/Y 0.57fF
C20496 INVX1_LOC_300/A INVX1_LOC_92/A 0.02fF
C20497 INVX1_LOC_46/Y INVX1_LOC_86/A 0.02fF
C20498 NAND2X1_LOC_753/Y INVX1_LOC_635/Y 0.05fF
C20499 INVX1_LOC_347/Y INVX1_LOC_41/Y 0.05fF
C20500 INVX1_LOC_624/Y INVX1_LOC_347/A 0.01fF
C20501 INVX1_LOC_47/Y NAND2X1_LOC_621/B 0.03fF
C20502 INVX1_LOC_31/Y INVX1_LOC_634/Y 0.44fF
C20503 INPUT_5 INVX1_LOC_40/A 0.03fF
C20504 INVX1_LOC_63/Y INVX1_LOC_74/Y 0.12fF
C20505 VDD INVX1_LOC_563/Y 0.25fF
C20506 INVX1_LOC_63/Y INVX1_LOC_483/Y 0.00fF
C20507 INVX1_LOC_62/Y INVX1_LOC_226/Y 0.08fF
C20508 INVX1_LOC_113/Y INVX1_LOC_638/A 0.04fF
C20509 NAND2X1_LOC_788/A NAND2X1_LOC_498/Y 0.05fF
C20510 INVX1_LOC_438/Y INVX1_LOC_445/Y 8.31fF
C20511 NAND2X1_LOC_788/A INVX1_LOC_570/A 0.04fF
C20512 VDD INVX1_LOC_393/A 0.00fF
C20513 INVX1_LOC_505/Y INVX1_LOC_114/A 0.03fF
C20514 INVX1_LOC_79/A INVX1_LOC_588/A 1.49fF
C20515 INVX1_LOC_203/Y INVX1_LOC_271/Y 0.01fF
C20516 INVX1_LOC_133/Y INVX1_LOC_53/Y 0.53fF
C20517 VDD INVX1_LOC_384/Y 0.29fF
C20518 VDD INVX1_LOC_526/A 0.59fF
C20519 INVX1_LOC_405/A NAND2X1_LOC_517/Y 0.29fF
C20520 INVX1_LOC_79/Y INVX1_LOC_274/Y 0.01fF
C20521 INVX1_LOC_418/A INVX1_LOC_395/A 0.22fF
C20522 INVX1_LOC_558/A INVX1_LOC_395/A 0.10fF
C20523 NAND2X1_LOC_331/A INVX1_LOC_512/Y 0.03fF
C20524 NAND2X1_LOC_759/B INVX1_LOC_53/Y -0.00fF
C20525 VDD INVX1_LOC_197/A 0.17fF
C20526 INVX1_LOC_655/A INVX1_LOC_92/A 0.21fF
C20527 NAND2X1_LOC_69/B INVX1_LOC_366/Y 0.01fF
C20528 INVX1_LOC_166/A INVX1_LOC_109/Y 0.03fF
C20529 INVX1_LOC_560/A NAND2X1_LOC_538/B 0.04fF
C20530 NAND2X1_LOC_582/a_36_24# GATE_865 0.00fF
C20531 VDD INVX1_LOC_124/Y 0.21fF
C20532 INVX1_LOC_174/Y INVX1_LOC_366/A 0.01fF
C20533 INVX1_LOC_558/A NAND2X1_LOC_136/a_36_24# 0.01fF
C20534 VDD NAND2X1_LOC_416/Y 0.40fF
C20535 VDD NAND2X1_LOC_285/B 0.01fF
C20536 INVX1_LOC_551/Y INVX1_LOC_51/Y 0.18fF
C20537 NAND2X1_LOC_79/B INVX1_LOC_366/A 0.01fF
C20538 INVX1_LOC_426/Y INVX1_LOC_159/Y 0.01fF
C20539 INVX1_LOC_438/A INVX1_LOC_145/Y 0.34fF
C20540 VDD NAND2X1_LOC_106/B 0.54fF
C20541 NAND2X1_LOC_45/Y INVX1_LOC_544/A 0.10fF
C20542 INVX1_LOC_17/Y INVX1_LOC_206/Y 0.48fF
C20543 NAND2X1_LOC_15/a_36_24# INVX1_LOC_99/Y 0.00fF
C20544 INVX1_LOC_301/A INPUT_1 0.09fF
C20545 INVX1_LOC_395/A NAND2X1_LOC_755/B 0.07fF
C20546 INVX1_LOC_584/Y INVX1_LOC_358/Y 0.18fF
C20547 VDD NAND2X1_LOC_174/B 0.14fF
C20548 INVX1_LOC_266/A INVX1_LOC_551/Y 0.10fF
C20549 NAND2X1_LOC_669/Y INVX1_LOC_315/Y 0.07fF
C20550 VDD INVX1_LOC_260/Y 0.21fF
C20551 INVX1_LOC_211/Y INVX1_LOC_395/A 0.03fF
C20552 INVX1_LOC_578/A INVX1_LOC_545/A 0.02fF
C20553 INVX1_LOC_501/Y INVX1_LOC_511/A 0.06fF
C20554 VDD INVX1_LOC_173/Y 0.39fF
C20555 INVX1_LOC_7/A NAND2X1_LOC_531/Y 0.01fF
C20556 NAND2X1_LOC_39/Y NAND2X1_LOC_39/a_36_24# 0.00fF
C20557 INVX1_LOC_144/Y NAND2X1_LOC_677/Y 0.01fF
C20558 INVX1_LOC_19/Y INPUT_4 0.02fF
C20559 INVX1_LOC_560/A INVX1_LOC_159/Y 0.02fF
C20560 INVX1_LOC_445/Y INVX1_LOC_219/Y 0.93fF
C20561 INVX1_LOC_255/Y INVX1_LOC_352/Y 0.03fF
C20562 INVX1_LOC_65/Y INVX1_LOC_59/Y 0.03fF
C20563 INVX1_LOC_412/Y INVX1_LOC_359/Y 0.01fF
C20564 INVX1_LOC_202/A NAND2X1_LOC_52/Y 0.02fF
C20565 INVX1_LOC_435/Y INVX1_LOC_672/A 0.18fF
C20566 NAND2X1_LOC_551/a_36_24# INVX1_LOC_412/A 0.00fF
C20567 INPUT_0 INVX1_LOC_117/Y 0.16fF
C20568 INVX1_LOC_224/Y INVX1_LOC_230/Y 0.17fF
C20569 INVX1_LOC_501/A INVX1_LOC_638/A 0.07fF
C20570 NAND2X1_LOC_788/A INVX1_LOC_47/Y 0.04fF
C20571 INVX1_LOC_395/A INVX1_LOC_46/Y 0.49fF
C20572 INVX1_LOC_581/A INVX1_LOC_53/Y 0.08fF
C20573 INVX1_LOC_53/Y INVX1_LOC_633/Y 0.01fF
C20574 INVX1_LOC_683/Y NAND2X1_LOC_471/a_36_24# 0.01fF
C20575 INVX1_LOC_435/A INVX1_LOC_76/Y 0.01fF
C20576 NAND2X1_LOC_475/A INVX1_LOC_296/A 0.02fF
C20577 INVX1_LOC_65/Y INVX1_LOC_48/Y 0.03fF
C20578 INVX1_LOC_400/A NAND2X1_LOC_318/A 0.14fF
C20579 INVX1_LOC_451/A INVX1_LOC_171/Y 0.03fF
C20580 VDD NAND2X1_LOC_555/B 0.17fF
C20581 INVX1_LOC_444/Y INVX1_LOC_172/Y 0.05fF
C20582 INVX1_LOC_381/A NAND2X1_LOC_414/a_36_24# 0.00fF
C20583 INVX1_LOC_150/A INVX1_LOC_498/Y 0.06fF
C20584 NAND2X1_LOC_242/A INVX1_LOC_63/Y 0.03fF
C20585 INVX1_LOC_613/Y NAND2X1_LOC_513/A 0.02fF
C20586 INVX1_LOC_17/Y INVX1_LOC_686/A 0.15fF
C20587 INVX1_LOC_95/Y INVX1_LOC_531/Y 0.04fF
C20588 NAND2X1_LOC_332/B INVX1_LOC_50/Y 0.03fF
C20589 INVX1_LOC_21/Y INVX1_LOC_449/A 0.10fF
C20590 NAND2X1_LOC_513/A NAND2X1_LOC_612/A 0.07fF
C20591 INVX1_LOC_447/Y INVX1_LOC_134/Y 0.00fF
C20592 INVX1_LOC_587/A NAND2X1_LOC_822/Y 0.01fF
C20593 INVX1_LOC_400/Y INVX1_LOC_69/Y 0.03fF
C20594 NAND2X1_LOC_153/a_36_24# INVX1_LOC_555/A 0.00fF
C20595 NAND2X1_LOC_548/B INVX1_LOC_35/Y 0.01fF
C20596 NAND2X1_LOC_336/B INVX1_LOC_304/Y 0.10fF
C20597 INVX1_LOC_20/Y INPUT_1 0.06fF
C20598 INVX1_LOC_355/A NAND2X1_LOC_449/B 0.05fF
C20599 NAND2X1_LOC_788/A INVX1_LOC_119/Y 0.03fF
C20600 INVX1_LOC_546/Y INVX1_LOC_49/Y 0.01fF
C20601 INVX1_LOC_35/Y INVX1_LOC_635/A 0.02fF
C20602 NAND2X1_LOC_697/Y NAND2X1_LOC_677/Y 0.22fF
C20603 NAND2X1_LOC_516/a_36_24# NAND2X1_LOC_307/B 0.01fF
C20604 INVX1_LOC_174/Y INVX1_LOC_6/Y 0.01fF
C20605 INVX1_LOC_317/Y INVX1_LOC_199/Y 0.03fF
C20606 INVX1_LOC_21/Y INVX1_LOC_274/A 0.08fF
C20607 INVX1_LOC_416/A NAND2X1_LOC_542/a_36_24# 0.02fF
C20608 INVX1_LOC_35/Y NAND2X1_LOC_237/Y 0.34fF
C20609 INVX1_LOC_288/Y INVX1_LOC_290/A 0.14fF
C20610 INVX1_LOC_166/A INVX1_LOC_126/Y 0.01fF
C20611 INVX1_LOC_392/Y INVX1_LOC_49/Y 0.02fF
C20612 INVX1_LOC_270/A INVX1_LOC_31/Y 0.01fF
C20613 INVX1_LOC_602/A INVX1_LOC_298/A 0.03fF
C20614 NAND2X1_LOC_79/B INVX1_LOC_6/Y 0.01fF
C20615 INVX1_LOC_579/Y INVX1_LOC_259/Y 0.54fF
C20616 INVX1_LOC_54/Y INVX1_LOC_134/Y 0.17fF
C20617 INVX1_LOC_213/Y NAND2X1_LOC_496/Y 0.07fF
C20618 INVX1_LOC_449/A NAND2X1_LOC_274/a_36_24# 0.00fF
C20619 INVX1_LOC_21/Y INVX1_LOC_209/A 0.00fF
C20620 INVX1_LOC_20/Y INVX1_LOC_292/Y 0.06fF
C20621 INVX1_LOC_293/Y NAND2X1_LOC_496/a_36_24# 0.01fF
C20622 INVX1_LOC_371/Y INVX1_LOC_665/Y 0.16fF
C20623 INVX1_LOC_287/A INVX1_LOC_48/Y 0.00fF
C20624 INVX1_LOC_21/Y INVX1_LOC_195/Y 0.23fF
C20625 INVX1_LOC_17/Y INVX1_LOC_452/A 0.11fF
C20626 NAND2X1_LOC_48/Y INVX1_LOC_54/Y 0.01fF
C20627 INVX1_LOC_261/A NAND2X1_LOC_328/a_36_24# 0.02fF
C20628 INVX1_LOC_552/Y INVX1_LOC_100/Y 0.00fF
C20629 INVX1_LOC_35/Y INVX1_LOC_230/A 0.09fF
C20630 INVX1_LOC_603/Y NAND2X1_LOC_333/B 0.07fF
C20631 INVX1_LOC_400/A INVX1_LOC_202/Y 0.00fF
C20632 INVX1_LOC_563/A INVX1_LOC_93/Y 0.01fF
C20633 INVX1_LOC_479/Y INVX1_LOC_59/Y 0.05fF
C20634 INVX1_LOC_425/A INVX1_LOC_9/Y 0.03fF
C20635 INVX1_LOC_137/Y INVX1_LOC_332/Y 0.02fF
C20636 INVX1_LOC_429/Y INVX1_LOC_430/Y 0.00fF
C20637 INVX1_LOC_524/Y INVX1_LOC_49/Y 0.07fF
C20638 INVX1_LOC_371/A INVX1_LOC_510/A 0.00fF
C20639 NAND2X1_LOC_122/a_36_24# INVX1_LOC_62/Y 0.01fF
C20640 INVX1_LOC_49/Y INVX1_LOC_59/A 0.01fF
C20641 INVX1_LOC_442/A INVX1_LOC_119/Y 0.02fF
C20642 INVX1_LOC_607/Y INVX1_LOC_117/Y 0.09fF
C20643 NAND2X1_LOC_843/A NAND2X1_LOC_106/B 0.08fF
C20644 INVX1_LOC_257/A INVX1_LOC_134/Y 0.03fF
C20645 INVX1_LOC_268/Y NAND2X1_LOC_334/B 0.04fF
C20646 INVX1_LOC_373/A INVX1_LOC_148/Y 0.00fF
C20647 INVX1_LOC_367/A INVX1_LOC_49/Y 0.00fF
C20648 INVX1_LOC_166/A NAND2X1_LOC_320/Y 0.02fF
C20649 INVX1_LOC_93/Y INVX1_LOC_115/A 0.02fF
C20650 INVX1_LOC_31/Y NAND2X1_LOC_755/B 0.03fF
C20651 INVX1_LOC_50/Y INVX1_LOC_503/Y 0.21fF
C20652 INPUT_2 INVX1_LOC_9/Y 0.04fF
C20653 INVX1_LOC_126/A INVX1_LOC_9/Y 0.00fF
C20654 NAND2X1_LOC_836/B INVX1_LOC_29/Y 0.01fF
C20655 INVX1_LOC_84/A INVX1_LOC_206/A 0.00fF
C20656 INVX1_LOC_318/A INVX1_LOC_59/Y 0.00fF
C20657 INVX1_LOC_635/A INVX1_LOC_621/Y 0.14fF
C20658 INVX1_LOC_93/Y INVX1_LOC_349/Y -0.03fF
C20659 INVX1_LOC_293/Y INVX1_LOC_245/A 0.00fF
C20660 INVX1_LOC_211/Y INVX1_LOC_31/Y 0.01fF
C20661 NAND2X1_LOC_307/A INVX1_LOC_376/Y 0.07fF
C20662 INVX1_LOC_550/Y INVX1_LOC_93/Y 0.01fF
C20663 INVX1_LOC_374/A INVX1_LOC_74/Y 0.12fF
C20664 INVX1_LOC_266/Y INVX1_LOC_41/Y 0.01fF
C20665 NAND2X1_LOC_297/Y INVX1_LOC_50/Y 0.02fF
C20666 INVX1_LOC_161/A INVX1_LOC_496/A 0.06fF
C20667 INVX1_LOC_69/Y INVX1_LOC_537/A 0.44fF
C20668 INVX1_LOC_545/Y INVX1_LOC_376/Y 0.01fF
C20669 NAND2X1_LOC_409/Y INVX1_LOC_366/A 0.02fF
C20670 INVX1_LOC_243/A INVX1_LOC_63/Y 0.01fF
C20671 INVX1_LOC_47/Y INVX1_LOC_116/Y 0.03fF
C20672 INVX1_LOC_392/A INVX1_LOC_387/Y 0.05fF
C20673 INVX1_LOC_298/A INVX1_LOC_117/Y 0.03fF
C20674 INVX1_LOC_51/Y NAND2X1_LOC_410/Y 0.02fF
C20675 NAND2X1_LOC_310/a_36_24# INVX1_LOC_92/A 0.00fF
C20676 INVX1_LOC_550/A INVX1_LOC_93/Y 0.00fF
C20677 NAND2X1_LOC_57/Y INVX1_LOC_63/Y 0.02fF
C20678 INVX1_LOC_68/Y INVX1_LOC_479/A 0.00fF
C20679 INVX1_LOC_17/Y NAND2X1_LOC_334/A 0.03fF
C20680 INVX1_LOC_416/A NAND2X1_LOC_542/A 0.10fF
C20681 INVX1_LOC_21/Y INVX1_LOC_328/Y 0.13fF
C20682 INVX1_LOC_555/A INVX1_LOC_186/Y 0.04fF
C20683 INVX1_LOC_47/Y NAND2X1_LOC_432/Y -0.00fF
C20684 INVX1_LOC_392/A INVX1_LOC_49/Y 0.01fF
C20685 INVX1_LOC_80/A INVX1_LOC_114/A 0.04fF
C20686 INVX1_LOC_90/A INVX1_LOC_90/Y 0.01fF
C20687 INVX1_LOC_95/A INVX1_LOC_59/Y 0.01fF
C20688 INVX1_LOC_179/A INVX1_LOC_99/Y 0.03fF
C20689 INVX1_LOC_31/Y INVX1_LOC_46/Y 0.26fF
C20690 INVX1_LOC_160/A INVX1_LOC_245/A 0.00fF
C20691 INVX1_LOC_93/Y INVX1_LOC_387/Y 0.03fF
C20692 INVX1_LOC_51/Y INVX1_LOC_634/Y 0.08fF
C20693 INPUT_2 INVX1_LOC_13/Y 0.64fF
C20694 INVX1_LOC_587/Y NAND2X1_LOC_827/Y 0.01fF
C20695 INVX1_LOC_54/Y INVX1_LOC_65/A 0.01fF
C20696 INVX1_LOC_166/A INVX1_LOC_199/Y 0.03fF
C20697 INVX1_LOC_89/Y NAND2X1_LOC_308/A 0.11fF
C20698 NAND2X1_LOC_451/B INVX1_LOC_495/A 0.00fF
C20699 INVX1_LOC_421/A INVX1_LOC_69/Y 0.08fF
C20700 NAND2X1_LOC_600/a_36_24# INVX1_LOC_376/Y 0.00fF
C20701 INVX1_LOC_435/A NAND2X1_LOC_264/a_36_24# 0.01fF
C20702 INVX1_LOC_469/Y INVX1_LOC_63/Y 0.00fF
C20703 INVX1_LOC_63/Y INVX1_LOC_350/Y 0.04fF
C20704 INVX1_LOC_93/Y INVX1_LOC_49/Y 2.64fF
C20705 INVX1_LOC_116/Y INVX1_LOC_119/Y 0.09fF
C20706 INVX1_LOC_479/A INVX1_LOC_675/Y 0.01fF
C20707 INVX1_LOC_369/A NAND2X1_LOC_489/a_36_24# 0.01fF
C20708 INVX1_LOC_75/Y INVX1_LOC_519/A 0.02fF
C20709 INVX1_LOC_11/Y INVX1_LOC_114/A 0.04fF
C20710 INVX1_LOC_93/Y INVX1_LOC_533/A 0.01fF
C20711 NAND2X1_LOC_699/a_36_24# INVX1_LOC_198/A 0.00fF
C20712 INVX1_LOC_164/Y INVX1_LOC_491/A 0.12fF
C20713 INVX1_LOC_119/Y NAND2X1_LOC_432/Y 0.03fF
C20714 INVX1_LOC_26/Y INVX1_LOC_345/A 0.48fF
C20715 INVX1_LOC_242/Y INVX1_LOC_50/Y 0.01fF
C20716 INVX1_LOC_62/Y INVX1_LOC_252/Y 0.03fF
C20717 INPUT_1 INVX1_LOC_655/A 0.09fF
C20718 INVX1_LOC_41/Y NAND2X1_LOC_459/a_36_24# 0.00fF
C20719 INVX1_LOC_511/Y INVX1_LOC_479/A 0.02fF
C20720 INVX1_LOC_274/A INVX1_LOC_209/Y 0.07fF
C20721 INVX1_LOC_675/A INVX1_LOC_49/Y 0.07fF
C20722 INVX1_LOC_335/A INVX1_LOC_41/Y 0.09fF
C20723 NAND2X1_LOC_192/A INVX1_LOC_496/A 0.02fF
C20724 NAND2X1_LOC_277/a_36_24# INVX1_LOC_655/A 0.01fF
C20725 INVX1_LOC_105/Y INVX1_LOC_41/Y 0.01fF
C20726 INVX1_LOC_49/Y NAND2X1_LOC_334/B 0.02fF
C20727 INVX1_LOC_376/A INVX1_LOC_376/Y 0.08fF
C20728 INVX1_LOC_253/Y INVX1_LOC_79/A 0.09fF
C20729 NAND2X1_LOC_88/Y NAND2X1_LOC_86/Y 0.15fF
C20730 INVX1_LOC_48/Y INVX1_LOC_588/A 0.05fF
C20731 NAND2X1_LOC_136/Y INVX1_LOC_199/Y 0.03fF
C20732 INVX1_LOC_410/A INVX1_LOC_90/Y 0.01fF
C20733 NAND2X1_LOC_333/B INVX1_LOC_91/A 0.04fF
C20734 NAND2X1_LOC_409/Y INVX1_LOC_6/Y 0.03fF
C20735 INVX1_LOC_117/Y INVX1_LOC_211/A 0.07fF
C20736 INVX1_LOC_63/Y INVX1_LOC_79/A 0.37fF
C20737 INVX1_LOC_531/Y INVX1_LOC_199/Y 0.15fF
C20738 INPUT_6 VDD 0.27fF
C20739 INVX1_LOC_31/Y INVX1_LOC_75/A 0.00fF
C20740 INVX1_LOC_62/Y NAND2X1_LOC_827/Y 0.01fF
C20741 NAND2X1_LOC_836/B INVX1_LOC_74/Y 0.02fF
C20742 INVX1_LOC_6/Y NAND2X1_LOC_497/a_36_24# 0.00fF
C20743 INVX1_LOC_63/Y NAND2X1_LOC_396/Y 0.01fF
C20744 INVX1_LOC_584/A NAND2X1_LOC_637/A 0.05fF
C20745 INVX1_LOC_426/A INVX1_LOC_416/Y 0.03fF
C20746 NAND2X1_LOC_602/a_36_24# INVX1_LOC_376/Y 0.00fF
C20747 NAND2X1_LOC_88/a_36_24# INVX1_LOC_395/A 0.00fF
C20748 INVX1_LOC_26/Y INVX1_LOC_280/A 0.14fF
C20749 INVX1_LOC_447/A INVX1_LOC_490/Y 0.01fF
C20750 INVX1_LOC_51/A INVX1_LOC_412/Y 0.02fF
C20751 INVX1_LOC_301/A INVX1_LOC_134/A 0.02fF
C20752 NAND2X1_LOC_749/Y NAND2X1_LOC_750/a_36_24# 0.01fF
C20753 INVX1_LOC_224/Y NAND2X1_LOC_370/A 0.02fF
C20754 INVX1_LOC_224/Y INVX1_LOC_249/Y 0.03fF
C20755 INVX1_LOC_472/Y INVX1_LOC_588/A 0.01fF
C20756 INVX1_LOC_412/Y NAND2X1_LOC_173/Y 0.10fF
C20757 INVX1_LOC_578/A INVX1_LOC_249/Y 0.00fF
C20758 INVX1_LOC_239/Y NAND2X1_LOC_148/A 0.03fF
C20759 VDD INVX1_LOC_336/Y 0.21fF
C20760 INVX1_LOC_401/Y VDD 0.33fF
C20761 INVX1_LOC_578/A NAND2X1_LOC_122/Y 0.03fF
C20762 INVX1_LOC_400/Y INVX1_LOC_586/A 0.03fF
C20763 VDD NAND2X1_LOC_97/B 0.43fF
C20764 INVX1_LOC_558/A INVX1_LOC_51/Y 0.02fF
C20765 VDD INVX1_LOC_417/A -0.00fF
C20766 INVX1_LOC_601/A INVX1_LOC_145/Y 0.00fF
C20767 NAND2X1_LOC_249/Y NAND2X1_LOC_595/Y 0.06fF
C20768 NAND2X1_LOC_457/A INVX1_LOC_80/A 0.03fF
C20769 INVX1_LOC_198/A NAND2X1_LOC_86/Y 0.06fF
C20770 NAND2X1_LOC_387/a_36_24# INVX1_LOC_586/A 0.01fF
C20771 VDD NAND2X1_LOC_179/Y 0.09fF
C20772 INVX1_LOC_266/A INVX1_LOC_418/A 0.31fF
C20773 INVX1_LOC_206/Y NAND2X1_LOC_616/Y 0.01fF
C20774 INVX1_LOC_288/A INVX1_LOC_111/A 0.03fF
C20775 NAND2X1_LOC_331/A INVX1_LOC_147/A 0.01fF
C20776 NAND2X1_LOC_307/A INVX1_LOC_253/A 0.01fF
C20777 INVX1_LOC_545/Y INVX1_LOC_253/A 0.00fF
C20778 INVX1_LOC_80/A INVX1_LOC_547/Y 0.43fF
C20779 INVX1_LOC_563/A INVX1_LOC_395/A 0.01fF
C20780 INVX1_LOC_224/Y INVX1_LOC_248/Y 0.96fF
C20781 INPUT_0 INVX1_LOC_281/Y 0.03fF
C20782 VDD INVX1_LOC_440/Y 0.29fF
C20783 NAND2X1_LOC_61/A INVX1_LOC_543/Y 0.11fF
C20784 INVX1_LOC_381/A NAND2X1_LOC_472/a_36_24# 0.00fF
C20785 INVX1_LOC_206/Y INVX1_LOC_545/A 0.01fF
C20786 NAND2X1_LOC_13/Y INVX1_LOC_551/Y 0.03fF
C20787 INVX1_LOC_524/Y INVX1_LOC_76/Y 0.04fF
C20788 NAND2X1_LOC_373/Y INPUT_1 0.10fF
C20789 INVX1_LOC_301/Y INVX1_LOC_109/Y 0.03fF
C20790 INVX1_LOC_206/Y INVX1_LOC_108/Y 0.01fF
C20791 INVX1_LOC_167/Y INVX1_LOC_168/A 0.00fF
C20792 INPUT_0 INVX1_LOC_178/A 0.11fF
C20793 INVX1_LOC_266/A INVX1_LOC_270/A 0.03fF
C20794 VDD INVX1_LOC_280/Y 0.23fF
C20795 INVX1_LOC_191/Y INVX1_LOC_86/Y 0.32fF
C20796 INVX1_LOC_11/Y NAND2X1_LOC_457/A 0.03fF
C20797 INVX1_LOC_548/Y INVX1_LOC_548/A 0.02fF
C20798 NAND2X1_LOC_164/Y INVX1_LOC_396/A 0.23fF
C20799 INVX1_LOC_32/A INVX1_LOC_31/Y 0.03fF
C20800 VDD INVX1_LOC_525/Y 0.22fF
C20801 INVX1_LOC_51/Y NAND2X1_LOC_755/B 0.03fF
C20802 INVX1_LOC_492/A INVX1_LOC_523/A 0.03fF
C20803 INVX1_LOC_586/A INVX1_LOC_537/A 0.07fF
C20804 INVX1_LOC_11/Y INVX1_LOC_547/Y 0.15fF
C20805 INVX1_LOC_84/A INVX1_LOC_320/A 0.17fF
C20806 INVX1_LOC_133/Y INVX1_LOC_662/A 0.02fF
C20807 INVX1_LOC_41/Y INVX1_LOC_109/Y 0.03fF
C20808 INVX1_LOC_76/Y INVX1_LOC_516/A 0.00fF
C20809 INVX1_LOC_238/Y INVX1_LOC_89/Y 0.00fF
C20810 INVX1_LOC_383/A INVX1_LOC_510/A 0.02fF
C20811 NAND2X1_LOC_45/Y INVX1_LOC_69/Y 0.01fF
C20812 INVX1_LOC_292/A INVX1_LOC_620/A 0.05fF
C20813 INVX1_LOC_35/Y INVX1_LOC_666/A 0.01fF
C20814 NAND2X1_LOC_12/a_36_24# INVX1_LOC_35/Y 0.01fF
C20815 INVX1_LOC_239/Y INVX1_LOC_662/A 0.02fF
C20816 INVX1_LOC_400/A INVX1_LOC_76/Y 0.01fF
C20817 INVX1_LOC_288/A INVX1_LOC_117/Y 0.07fF
C20818 INVX1_LOC_469/Y INVX1_LOC_374/A 0.00fF
C20819 INVX1_LOC_11/Y INVX1_LOC_482/A 0.32fF
C20820 NAND2X1_LOC_336/a_36_24# INVX1_LOC_230/A 0.00fF
C20821 INVX1_LOC_270/A NAND2X1_LOC_267/a_36_24# 0.00fF
C20822 INVX1_LOC_414/A INVX1_LOC_63/Y 0.03fF
C20823 INVX1_LOC_206/Y INVX1_LOC_507/A 0.08fF
C20824 INVX1_LOC_93/Y NAND2X1_LOC_498/B 0.01fF
C20825 INVX1_LOC_177/Y INVX1_LOC_6/Y 0.02fF
C20826 INVX1_LOC_602/A INVX1_LOC_145/Y 0.08fF
C20827 INVX1_LOC_602/A NAND2X1_LOC_791/A 0.04fF
C20828 INVX1_LOC_266/Y NAND2X1_LOC_267/A 0.02fF
C20829 INVX1_LOC_521/Y INVX1_LOC_555/A 0.00fF
C20830 INVX1_LOC_168/A INVX1_LOC_137/Y 0.03fF
C20831 INVX1_LOC_545/A INVX1_LOC_686/A 0.01fF
C20832 INVX1_LOC_530/Y INVX1_LOC_31/Y 0.19fF
C20833 INPUT_0 INVX1_LOC_58/Y 0.07fF
C20834 INVX1_LOC_12/Y INVX1_LOC_600/A 0.06fF
C20835 INVX1_LOC_51/Y INVX1_LOC_46/Y 0.07fF
C20836 INVX1_LOC_617/Y INVX1_LOC_371/A 0.01fF
C20837 VDD INVX1_LOC_485/Y 0.21fF
C20838 INVX1_LOC_384/A INVX1_LOC_117/Y 0.07fF
C20839 INVX1_LOC_35/Y INVX1_LOC_492/Y 0.01fF
C20840 NAND2X1_LOC_535/a_36_24# INVX1_LOC_376/Y 0.00fF
C20841 INVX1_LOC_395/A INVX1_LOC_49/Y 0.29fF
C20842 INVX1_LOC_421/A INVX1_LOC_586/A 0.08fF
C20843 INVX1_LOC_360/Y INVX1_LOC_197/A 0.07fF
C20844 NAND2X1_LOC_498/Y INVX1_LOC_69/Y 0.07fF
C20845 INVX1_LOC_586/A INVX1_LOC_496/Y 0.03fF
C20846 INVX1_LOC_20/Y INVX1_LOC_50/Y 2.01fF
C20847 INVX1_LOC_362/Y INVX1_LOC_387/Y 0.01fF
C20848 NAND2X1_LOC_546/a_36_24# NAND2X1_LOC_521/Y 0.00fF
C20849 INVX1_LOC_93/Y INVX1_LOC_76/Y 0.19fF
C20850 NAND2X1_LOC_142/Y NAND2X1_LOC_342/A 0.18fF
C20851 INVX1_LOC_40/Y INVX1_LOC_333/A 0.00fF
C20852 NAND2X1_LOC_318/A INVX1_LOC_31/Y 0.00fF
C20853 NAND2X1_LOC_710/B INVX1_LOC_518/A 0.01fF
C20854 INVX1_LOC_21/Y INVX1_LOC_352/A 0.01fF
C20855 INVX1_LOC_255/Y INVX1_LOC_347/Y 0.04fF
C20856 NAND2X1_LOC_770/B NAND2X1_LOC_791/B 0.04fF
C20857 INVX1_LOC_54/Y INVX1_LOC_318/Y 0.07fF
C20858 INVX1_LOC_266/A INVX1_LOC_46/Y 0.07fF
C20859 NAND2X1_LOC_325/B INVX1_LOC_304/A 0.07fF
C20860 INVX1_LOC_20/Y INVX1_LOC_431/Y 0.44fF
C20861 INVX1_LOC_576/A INVX1_LOC_50/Y 0.02fF
C20862 INVX1_LOC_35/Y NAND2X1_LOC_72/Y 0.19fF
C20863 INVX1_LOC_335/A INVX1_LOC_358/Y 0.00fF
C20864 NAND2X1_LOC_249/Y NAND2X1_LOC_372/Y 0.33fF
C20865 VDD INVX1_LOC_66/Y 0.21fF
C20866 INPUT_1 INVX1_LOC_375/Y 0.01fF
C20867 INVX1_LOC_26/A INVX1_LOC_26/Y 0.02fF
C20868 INVX1_LOC_578/Y INVX1_LOC_188/Y 0.03fF
C20869 VDD NAND2X1_LOC_248/B 0.02fF
C20870 INVX1_LOC_108/A INVX1_LOC_367/A 0.03fF
C20871 NAND2X1_LOC_524/a_36_24# INPUT_1 0.00fF
C20872 INVX1_LOC_365/Y INVX1_LOC_46/Y 0.01fF
C20873 INVX1_LOC_166/A INVX1_LOC_53/Y 0.03fF
C20874 INVX1_LOC_21/Y INVX1_LOC_172/A 0.05fF
C20875 INVX1_LOC_54/Y INVX1_LOC_16/Y 0.02fF
C20876 INVX1_LOC_116/A INVX1_LOC_440/Y 0.02fF
C20877 INVX1_LOC_625/A NAND2X1_LOC_226/a_36_24# 0.01fF
C20878 INPUT_3 NAND2X1_LOC_82/a_36_24# 0.00fF
C20879 INVX1_LOC_560/Y INVX1_LOC_74/Y 0.08fF
C20880 INVX1_LOC_628/Y INVX1_LOC_259/Y 0.01fF
C20881 INVX1_LOC_208/A NAND2X1_LOC_237/Y 0.00fF
C20882 INVX1_LOC_85/Y INVX1_LOC_9/Y 0.01fF
C20883 NAND2X1_LOC_140/B INPUT_1 0.17fF
C20884 NAND2X1_LOC_673/A INVX1_LOC_35/Y 0.02fF
C20885 INVX1_LOC_17/Y INVX1_LOC_282/A 0.02fF
C20886 INVX1_LOC_76/Y INVX1_LOC_390/A 0.01fF
C20887 INVX1_LOC_683/Y INVX1_LOC_49/Y 0.02fF
C20888 INVX1_LOC_300/A INVX1_LOC_50/Y 0.07fF
C20889 INVX1_LOC_89/Y INVX1_LOC_134/Y 1.11fF
C20890 INVX1_LOC_374/A INVX1_LOC_79/A 0.06fF
C20891 INVX1_LOC_412/Y INVX1_LOC_441/A 0.14fF
C20892 INVX1_LOC_12/Y INVX1_LOC_484/A 0.02fF
C20893 NAND2X1_LOC_261/Y INVX1_LOC_664/A 0.04fF
C20894 NAND2X1_LOC_179/Y INVX1_LOC_103/Y 0.11fF
C20895 INVX1_LOC_412/Y INVX1_LOC_354/A 0.05fF
C20896 NAND2X1_LOC_587/a_36_24# INVX1_LOC_40/Y 0.00fF
C20897 INVX1_LOC_117/Y INVX1_LOC_145/Y 0.24fF
C20898 INVX1_LOC_335/Y NAND2X1_LOC_821/a_36_24# 0.01fF
C20899 INVX1_LOC_17/Y NAND2X1_LOC_318/a_36_24# 0.00fF
C20900 INVX1_LOC_188/Y INVX1_LOC_532/Y 0.14fF
C20901 INVX1_LOC_417/Y INVX1_LOC_253/Y 0.03fF
C20902 INVX1_LOC_435/A INVX1_LOC_32/Y 0.03fF
C20903 INVX1_LOC_69/Y INVX1_LOC_676/Y 0.03fF
C20904 INVX1_LOC_300/A INVX1_LOC_431/Y 0.04fF
C20905 INVX1_LOC_31/Y INVX1_LOC_349/Y 0.01fF
C20906 INVX1_LOC_48/Y INVX1_LOC_623/Y 0.03fF
C20907 INVX1_LOC_202/Y INVX1_LOC_31/Y 0.04fF
C20908 INVX1_LOC_501/A INVX1_LOC_134/Y 0.20fF
C20909 INVX1_LOC_384/Y INVX1_LOC_430/Y 0.05fF
C20910 INVX1_LOC_69/Y INVX1_LOC_99/Y 0.24fF
C20911 NAND2X1_LOC_231/a_36_24# INVX1_LOC_94/A 0.01fF
C20912 INVX1_LOC_35/Y NAND2X1_LOC_647/A 0.03fF
C20913 INVX1_LOC_607/Y INVX1_LOC_58/Y 0.04fF
C20914 NAND2X1_LOC_427/Y INVX1_LOC_41/Y 0.04fF
C20915 INVX1_LOC_258/Y INVX1_LOC_504/Y 0.94fF
C20916 INVX1_LOC_84/A INVX1_LOC_100/Y 0.39fF
C20917 NAND2X1_LOC_152/a_36_24# INVX1_LOC_662/A 0.01fF
C20918 INVX1_LOC_624/Y INVX1_LOC_252/Y 0.01fF
C20919 NAND2X1_LOC_243/A NAND2X1_LOC_204/a_36_24# 0.00fF
C20920 INVX1_LOC_63/Y INVX1_LOC_59/Y 0.06fF
C20921 INVX1_LOC_449/A INVX1_LOC_26/Y 0.07fF
C20922 INVX1_LOC_93/Y INVX1_LOC_108/A 0.00fF
C20923 INVX1_LOC_53/Y NAND2X1_LOC_136/Y 0.04fF
C20924 NAND2X1_LOC_137/A INVX1_LOC_105/Y 0.00fF
C20925 INVX1_LOC_682/Y INVX1_LOC_363/Y 0.03fF
C20926 INVX1_LOC_35/Y INVX1_LOC_168/Y 0.04fF
C20927 INVX1_LOC_573/Y INVX1_LOC_514/A 0.00fF
C20928 NAND2X1_LOC_482/Y NAND2X1_LOC_253/Y 0.07fF
C20929 INVX1_LOC_274/A INVX1_LOC_26/Y 0.07fF
C20930 INVX1_LOC_63/Y NAND2X1_LOC_60/a_36_24# 0.00fF
C20931 INVX1_LOC_63/Y INVX1_LOC_48/Y 4.24fF
C20932 INVX1_LOC_84/A INVX1_LOC_483/Y 0.35fF
C20933 NAND2X1_LOC_7/a_36_24# INVX1_LOC_211/A 0.00fF
C20934 INVX1_LOC_176/A NAND2X1_LOC_41/a_36_24# 0.01fF
C20935 INVX1_LOC_298/A INVX1_LOC_58/Y 0.00fF
C20936 INVX1_LOC_58/Y INVX1_LOC_498/A 0.00fF
C20937 INVX1_LOC_100/Y NAND2X1_LOC_67/Y 0.02fF
C20938 INVX1_LOC_209/A INVX1_LOC_26/Y 0.03fF
C20939 INVX1_LOC_31/Y INVX1_LOC_49/Y 5.67fF
C20940 NAND2X1_LOC_614/a_36_24# INVX1_LOC_351/A 0.00fF
C20941 NAND2X1_LOC_837/A NAND2X1_LOC_753/Y 0.08fF
C20942 INVX1_LOC_134/Y NAND2X1_LOC_544/B 0.11fF
C20943 INVX1_LOC_406/Y INVX1_LOC_443/A 0.05fF
C20944 INVX1_LOC_89/Y INVX1_LOC_65/A 0.03fF
C20945 NAND2X1_LOC_320/Y INVX1_LOC_41/Y 0.11fF
C20946 INVX1_LOC_47/Y INVX1_LOC_69/Y 0.58fF
C20947 NAND2X1_LOC_104/a_36_24# INVX1_LOC_49/Y 0.01fF
C20948 INVX1_LOC_26/Y INVX1_LOC_195/Y 0.23fF
C20949 NAND2X1_LOC_775/B NAND2X1_LOC_545/A 0.18fF
C20950 INVX1_LOC_555/A NAND2X1_LOC_846/B 0.03fF
C20951 INVX1_LOC_280/A NAND2X1_LOC_275/Y 0.06fF
C20952 INVX1_LOC_54/Y INVX1_LOC_90/Y 0.10fF
C20953 INVX1_LOC_50/Y NAND2X1_LOC_269/B 0.01fF
C20954 INVX1_LOC_374/Y INVX1_LOC_114/A 0.00fF
C20955 NAND2X1_LOC_675/B INVX1_LOC_533/A 0.01fF
C20956 NAND2X1_LOC_491/Y INVX1_LOC_63/Y 0.06fF
C20957 NAND2X1_LOC_388/A INVX1_LOC_242/Y 0.07fF
C20958 INVX1_LOC_300/Y INVX1_LOC_674/Y 0.56fF
C20959 INVX1_LOC_314/Y NAND2X1_LOC_615/Y 0.07fF
C20960 NAND2X1_LOC_775/B INVX1_LOC_666/Y 0.07fF
C20961 INVX1_LOC_211/A NAND2X1_LOC_76/A 0.02fF
C20962 INVX1_LOC_49/Y INVX1_LOC_128/A 0.02fF
C20963 INVX1_LOC_69/Y INVX1_LOC_119/Y 0.21fF
C20964 INVX1_LOC_347/Y INVX1_LOC_26/Y 1.72fF
C20965 VDD INVX1_LOC_71/Y 0.24fF
C20966 VDD INVX1_LOC_7/A -0.00fF
C20967 INVX1_LOC_567/Y INVX1_LOC_92/A 0.02fF
C20968 INVX1_LOC_395/A INVX1_LOC_297/Y 0.03fF
C20969 INVX1_LOC_328/Y INVX1_LOC_26/Y 0.03fF
C20970 INVX1_LOC_419/A INVX1_LOC_62/Y 0.01fF
C20971 INVX1_LOC_660/Y INVX1_LOC_659/A 0.03fF
C20972 INVX1_LOC_41/Y INVX1_LOC_199/Y 0.12fF
C20973 NAND2X1_LOC_555/B INVX1_LOC_430/Y 0.02fF
C20974 INVX1_LOC_573/Y INVX1_LOC_62/Y 0.00fF
C20975 INVX1_LOC_518/A INVX1_LOC_128/Y 0.09fF
C20976 INVX1_LOC_459/A NAND2X1_LOC_589/a_36_24# 0.00fF
C20977 VDD INVX1_LOC_412/Y 0.22fF
C20978 INVX1_LOC_65/A NAND2X1_LOC_544/B 0.04fF
C20979 INVX1_LOC_156/A INVX1_LOC_636/A 0.03fF
C20980 NAND2X1_LOC_189/a_36_24# INVX1_LOC_62/Y 0.01fF
C20981 INVX1_LOC_58/Y INVX1_LOC_211/A 0.07fF
C20982 NAND2X1_LOC_543/B INVX1_LOC_442/A 0.03fF
C20983 INVX1_LOC_388/A INVX1_LOC_90/Y 0.00fF
C20984 INVX1_LOC_573/A NAND2X1_LOC_728/B 0.08fF
C20985 VDD INVX1_LOC_321/A 0.00fF
C20986 INVX1_LOC_206/Y NAND2X1_LOC_370/A 0.05fF
C20987 INVX1_LOC_448/Y INVX1_LOC_384/A 0.04fF
C20988 NAND2X1_LOC_45/Y INVX1_LOC_586/A 0.03fF
C20989 INVX1_LOC_206/Y NAND2X1_LOC_122/Y 0.03fF
C20990 INVX1_LOC_62/Y INVX1_LOC_505/Y 0.07fF
C20991 INVX1_LOC_665/A NAND2X1_LOC_844/A 0.17fF
C20992 INVX1_LOC_114/A INVX1_LOC_625/Y 0.03fF
C20993 INVX1_LOC_563/Y INVX1_LOC_45/Y 0.01fF
C20994 INVX1_LOC_617/Y VDD 1.32fF
C20995 INVX1_LOC_560/Y INVX1_LOC_566/A 0.03fF
C20996 VDD INVX1_LOC_176/Y 0.14fF
C20997 INVX1_LOC_37/Y INVX1_LOC_76/Y 0.01fF
C20998 INVX1_LOC_290/A NAND2X1_LOC_801/A 0.01fF
C20999 NAND2X1_LOC_753/a_36_24# NAND2X1_LOC_755/B 0.00fF
C21000 NAND2X1_LOC_498/Y INVX1_LOC_586/A 0.10fF
C21001 INVX1_LOC_395/A INVX1_LOC_76/Y 0.07fF
C21002 INVX1_LOC_420/Y INVX1_LOC_406/Y 0.61fF
C21003 INVX1_LOC_448/A INVX1_LOC_448/Y 0.01fF
C21004 INVX1_LOC_197/Y INVX1_LOC_275/A 4.02fF
C21005 NAND2X1_LOC_505/Y NAND2X1_LOC_318/A 0.16fF
C21006 NAND2X1_LOC_543/B INVX1_LOC_116/Y 0.02fF
C21007 INVX1_LOC_626/Y NAND2X1_LOC_513/A 0.06fF
C21008 INVX1_LOC_434/A INVX1_LOC_451/Y 0.01fF
C21009 INVX1_LOC_206/Y NAND2X1_LOC_393/Y 0.21fF
C21010 INVX1_LOC_312/Y NAND2X1_LOC_498/Y 0.07fF
C21011 INVX1_LOC_617/Y INVX1_LOC_383/A 0.01fF
C21012 NAND2X1_LOC_798/a_36_24# INVX1_LOC_288/A 0.00fF
C21013 NAND2X1_LOC_391/B NAND2X1_LOC_384/a_36_24# 0.02fF
C21014 INVX1_LOC_578/A INVX1_LOC_519/A 0.01fF
C21015 INVX1_LOC_553/Y NAND2X1_LOC_413/Y 0.15fF
C21016 NAND2X1_LOC_231/A NAND2X1_LOC_357/a_36_24# 0.00fF
C21017 NAND2X1_LOC_537/B INVX1_LOC_99/Y 0.05fF
C21018 INVX1_LOC_45/Y INVX1_LOC_197/A 0.06fF
C21019 NAND2X1_LOC_373/Y INVX1_LOC_50/Y 0.03fF
C21020 NAND2X1_LOC_13/Y INVX1_LOC_270/A 0.37fF
C21021 INVX1_LOC_390/A INVX1_LOC_192/A 0.02fF
C21022 INVX1_LOC_568/Y INVX1_LOC_523/A 0.00fF
C21023 INVX1_LOC_586/A INVX1_LOC_676/Y 0.09fF
C21024 INVX1_LOC_319/Y INVX1_LOC_194/A 0.06fF
C21025 INVX1_LOC_410/Y INVX1_LOC_371/A 0.20fF
C21026 INVX1_LOC_270/Y INVX1_LOC_92/A 0.01fF
C21027 INVX1_LOC_151/Y INVX1_LOC_496/Y 0.01fF
C21028 INVX1_LOC_301/A NAND2X1_LOC_388/A 0.02fF
C21029 NAND2X1_LOC_543/B INVX1_LOC_255/A 0.02fF
C21030 INVX1_LOC_158/A INVX1_LOC_31/Y 0.01fF
C21031 INVX1_LOC_649/Y INVX1_LOC_668/A 0.00fF
C21032 INVX1_LOC_358/A INVX1_LOC_356/A 0.18fF
C21033 INVX1_LOC_358/Y NAND2X1_LOC_427/Y 0.12fF
C21034 INVX1_LOC_586/A INVX1_LOC_99/Y 0.45fF
C21035 INVX1_LOC_85/Y INVX1_LOC_42/Y 0.67fF
C21036 INVX1_LOC_3/Y NAND2X1_LOC_836/B 0.02fF
C21037 INVX1_LOC_202/Y INVX1_LOC_51/Y 0.00fF
C21038 INVX1_LOC_395/A NAND2X1_LOC_503/Y 0.08fF
C21039 INVX1_LOC_374/A INVX1_LOC_48/Y 0.03fF
C21040 INPUT_0 NAND2X1_LOC_689/B 0.00fF
C21041 INVX1_LOC_17/Y NAND2X1_LOC_845/a_36_24# 0.00fF
C21042 NAND2X1_LOC_475/A INVX1_LOC_69/Y 0.07fF
C21043 INVX1_LOC_76/Y INVX1_LOC_189/Y 0.02fF
C21044 INVX1_LOC_596/A INVX1_LOC_680/Y 0.00fF
C21045 NAND2X1_LOC_537/B INVX1_LOC_47/Y 0.01fF
C21046 NAND2X1_LOC_56/Y INVX1_LOC_12/Y 0.01fF
C21047 INVX1_LOC_265/Y INVX1_LOC_69/Y 0.01fF
C21048 INVX1_LOC_68/Y NAND2X1_LOC_615/B 0.01fF
C21049 INVX1_LOC_257/Y INVX1_LOC_58/Y 0.07fF
C21050 NAND2X1_LOC_176/a_36_24# INVX1_LOC_98/Y 0.00fF
C21051 INVX1_LOC_80/A NAND2X1_LOC_113/a_36_24# 0.01fF
C21052 NAND2X1_LOC_498/B INVX1_LOC_31/Y -0.05fF
C21053 INVX1_LOC_392/Y INVX1_LOC_32/Y 0.01fF
C21054 INVX1_LOC_300/A INVX1_LOC_187/A 0.10fF
C21055 NAND2X1_LOC_796/a_36_24# INVX1_LOC_581/A 0.00fF
C21056 NAND2X1_LOC_768/A NAND2X1_LOC_113/a_36_24# 0.00fF
C21057 NAND2X1_LOC_107/Y INVX1_LOC_106/A 0.07fF
C21058 VDD INVX1_LOC_664/A 0.00fF
C21059 NAND2X1_LOC_332/B INVX1_LOC_117/Y 0.03fF
C21060 INVX1_LOC_173/Y INVX1_LOC_45/Y 0.01fF
C21061 INVX1_LOC_649/Y INVX1_LOC_668/Y 0.01fF
C21062 NAND2X1_LOC_307/A INVX1_LOC_251/A 0.28fF
C21063 INVX1_LOC_287/A INVX1_LOC_155/Y 0.20fF
C21064 INVX1_LOC_387/Y INVX1_LOC_51/Y 0.03fF
C21065 NAND2X1_LOC_790/B INVX1_LOC_203/A 0.03fF
C21066 INVX1_LOC_31/Y INVX1_LOC_76/Y 0.17fF
C21067 INVX1_LOC_17/Y NAND2X1_LOC_603/Y 0.01fF
C21068 INVX1_LOC_560/Y INVX1_LOC_79/A 0.04fF
C21069 NAND2X1_LOC_192/a_36_24# INVX1_LOC_54/Y 0.01fF
C21070 INVX1_LOC_401/A INPUT_1 0.01fF
C21071 INVX1_LOC_103/Y INVX1_LOC_119/A 0.00fF
C21072 NAND2X1_LOC_20/Y NAND2X1_LOC_84/B 0.04fF
C21073 INVX1_LOC_47/Y INVX1_LOC_586/A 0.16fF
C21074 INPUT_0 INVX1_LOC_245/A 0.06fF
C21075 INVX1_LOC_117/Y INVX1_LOC_125/Y 0.06fF
C21076 INVX1_LOC_602/A INVX1_LOC_598/A 0.39fF
C21077 INVX1_LOC_116/Y INVX1_LOC_469/A 0.01fF
C21078 INVX1_LOC_51/Y INVX1_LOC_49/Y 0.29fF
C21079 INVX1_LOC_502/Y INVX1_LOC_69/Y 0.01fF
C21080 NAND2X1_LOC_122/Y NAND2X1_LOC_674/a_36_24# 0.00fF
C21081 INVX1_LOC_438/A NAND2X1_LOC_269/B 0.01fF
C21082 NAND2X1_LOC_122/Y NAND2X1_LOC_334/A 0.03fF
C21083 INVX1_LOC_54/Y NAND2X1_LOC_545/B 0.00fF
C21084 INVX1_LOC_99/A INVX1_LOC_304/A 0.02fF
C21085 NAND2X1_LOC_132/a_36_24# INVX1_LOC_126/A 0.00fF
C21086 INVX1_LOC_50/Y INVX1_LOC_375/Y 0.01fF
C21087 INVX1_LOC_145/Y INVX1_LOC_178/A 0.08fF
C21088 INVX1_LOC_45/A INVX1_LOC_93/A 0.10fF
C21089 INVX1_LOC_137/Y INVX1_LOC_35/Y 0.03fF
C21090 INVX1_LOC_270/A INVX1_LOC_361/A 0.03fF
C21091 INVX1_LOC_286/A INVX1_LOC_245/A 0.01fF
C21092 INVX1_LOC_127/Y NAND2X1_LOC_130/Y 0.02fF
C21093 NAND2X1_LOC_838/a_36_24# INVX1_LOC_59/A 0.00fF
C21094 INVX1_LOC_312/Y INVX1_LOC_47/Y 0.01fF
C21095 INVX1_LOC_444/Y INVX1_LOC_172/A 0.19fF
C21096 INVX1_LOC_315/Y INVX1_LOC_272/A 0.00fF
C21097 INVX1_LOC_54/Y INVX1_LOC_98/Y 0.10fF
C21098 INVX1_LOC_11/Y INVX1_LOC_303/Y 0.03fF
C21099 INVX1_LOC_586/A INVX1_LOC_119/Y 0.01fF
C21100 INVX1_LOC_105/A INVX1_LOC_510/A 0.07fF
C21101 NAND2X1_LOC_835/A INVX1_LOC_99/Y 0.01fF
C21102 INVX1_LOC_256/A INVX1_LOC_93/Y 0.01fF
C21103 INVX1_LOC_586/A NAND2X1_LOC_66/Y 0.00fF
C21104 INVX1_LOC_178/Y INVX1_LOC_88/Y 0.00fF
C21105 INVX1_LOC_202/Y INVX1_LOC_254/A 0.00fF
C21106 NAND2X1_LOC_308/A NAND2X1_LOC_418/Y 0.36fF
C21107 INVX1_LOC_400/A INVX1_LOC_32/Y 0.08fF
C21108 INVX1_LOC_392/A INVX1_LOC_32/Y 0.00fF
C21109 NAND2X1_LOC_197/a_36_24# NAND2X1_LOC_52/Y 0.01fF
C21110 INVX1_LOC_84/A NAND2X1_LOC_558/B 0.02fF
C21111 INVX1_LOC_428/A INVX1_LOC_479/A 0.03fF
C21112 INVX1_LOC_80/A INVX1_LOC_9/Y 0.06fF
C21113 INVX1_LOC_25/Y INVX1_LOC_69/Y 0.12fF
C21114 INVX1_LOC_84/A INVX1_LOC_79/A 0.01fF
C21115 INVX1_LOC_145/Y INVX1_LOC_58/Y 0.18fF
C21116 INVX1_LOC_211/Y INVX1_LOC_380/Y 0.01fF
C21117 NAND2X1_LOC_638/A NAND2X1_LOC_719/A 0.02fF
C21118 INVX1_LOC_591/Y INVX1_LOC_79/A 0.01fF
C21119 INVX1_LOC_93/Y INVX1_LOC_32/Y 0.61fF
C21120 INVX1_LOC_261/Y INVX1_LOC_259/Y 0.02fF
C21121 INVX1_LOC_235/Y INVX1_LOC_280/A 0.07fF
C21122 NAND2X1_LOC_513/A INVX1_LOC_655/A 0.29fF
C21123 NAND2X1_LOC_123/A INVX1_LOC_245/A 0.01fF
C21124 INVX1_LOC_117/Y NAND2X1_LOC_128/B 0.28fF
C21125 INVX1_LOC_218/Y NAND2X1_LOC_344/B 0.14fF
C21126 INVX1_LOC_543/A INVX1_LOC_7/Y 0.01fF
C21127 NAND2X1_LOC_187/Y INVX1_LOC_338/Y 0.04fF
C21128 NAND2X1_LOC_686/a_36_24# INVX1_LOC_245/A 0.01fF
C21129 INVX1_LOC_53/Y INVX1_LOC_41/Y 0.10fF
C21130 INVX1_LOC_199/Y NAND2X1_LOC_267/A 0.04fF
C21131 INVX1_LOC_54/Y INVX1_LOC_338/Y 0.18fF
C21132 INVX1_LOC_632/A INVX1_LOC_454/Y 0.00fF
C21133 INVX1_LOC_651/A NAND2X1_LOC_843/B 0.01fF
C21134 NAND2X1_LOC_409/Y INVX1_LOC_29/Y 0.04fF
C21135 INVX1_LOC_80/A INVX1_LOC_62/Y 5.22fF
C21136 INVX1_LOC_11/Y INVX1_LOC_9/Y 0.88fF
C21137 INVX1_LOC_653/Y INVX1_LOC_633/Y 0.07fF
C21138 INVX1_LOC_675/A INVX1_LOC_32/Y 0.07fF
C21139 INVX1_LOC_527/Y INVX1_LOC_245/A 0.03fF
C21140 INVX1_LOC_372/Y INVX1_LOC_348/Y 0.00fF
C21141 INVX1_LOC_117/Y INVX1_LOC_242/Y 0.23fF
C21142 INVX1_LOC_11/Y INVX1_LOC_166/Y 0.03fF
C21143 INVX1_LOC_193/A INVX1_LOC_100/Y 0.02fF
C21144 INVX1_LOC_12/Y INVX1_LOC_223/A 0.01fF
C21145 INVX1_LOC_166/A INVX1_LOC_653/A 0.36fF
C21146 INVX1_LOC_662/A INVX1_LOC_239/A 0.02fF
C21147 INVX1_LOC_11/Y INVX1_LOC_62/Y 0.93fF
C21148 INVX1_LOC_7/Y INVX1_LOC_86/A 0.01fF
C21149 INVX1_LOC_386/A NAND2X1_LOC_344/B 0.00fF
C21150 INVX1_LOC_43/A INVX1_LOC_41/Y 0.09fF
C21151 NAND2X1_LOC_814/a_36_24# INVX1_LOC_6/Y 0.00fF
C21152 INVX1_LOC_89/Y INVX1_LOC_90/Y 2.91fF
C21153 INVX1_LOC_35/Y INVX1_LOC_647/Y 0.02fF
C21154 INVX1_LOC_258/Y INVX1_LOC_114/A 0.02fF
C21155 NAND2X1_LOC_647/A NAND2X1_LOC_647/a_36_24# 0.00fF
C21156 NAND2X1_LOC_657/a_36_24# INVX1_LOC_376/Y 0.00fF
C21157 NAND2X1_LOC_532/Y INVX1_LOC_74/Y 0.00fF
C21158 NAND2X1_LOC_698/Y INVX1_LOC_531/Y 0.02fF
C21159 INVX1_LOC_479/A NAND2X1_LOC_284/A 0.04fF
C21160 VDD INVX1_LOC_553/Y 0.07fF
C21161 NAND2X1_LOC_433/Y INVX1_LOC_166/Y 0.10fF
C21162 VDD INVX1_LOC_410/Y 0.32fF
C21163 INVX1_LOC_361/A INVX1_LOC_75/A 0.06fF
C21164 INPUT_1 INVX1_LOC_92/A 0.05fF
C21165 NAND2X1_LOC_768/B INVX1_LOC_479/A 0.02fF
C21166 NAND2X1_LOC_865/a_36_24# INVX1_LOC_109/Y 0.01fF
C21167 NAND2X1_LOC_433/Y INVX1_LOC_62/Y 0.07fF
C21168 VDD INVX1_LOC_375/A 0.00fF
C21169 INVX1_LOC_409/Y INVX1_LOC_442/A 0.01fF
C21170 NAND2X1_LOC_322/Y INVX1_LOC_442/A 0.26fF
C21171 INVX1_LOC_393/Y NAND2X1_LOC_457/A 0.17fF
C21172 NAND2X1_LOC_249/Y INVX1_LOC_651/Y 0.42fF
C21173 NAND2X1_LOC_65/Y VDD 0.01fF
C21174 NAND2X1_LOC_475/A INVX1_LOC_586/A 0.10fF
C21175 INVX1_LOC_584/Y INVX1_LOC_373/A 0.32fF
C21176 NAND2X1_LOC_301/B INVX1_LOC_634/Y 0.07fF
C21177 VDD NAND2X1_LOC_780/A -0.00fF
C21178 INVX1_LOC_553/Y INVX1_LOC_510/Y 0.00fF
C21179 VDD INVX1_LOC_406/Y 0.71fF
C21180 INVX1_LOC_206/Y INVX1_LOC_356/A 0.02fF
C21181 INVX1_LOC_549/A INVX1_LOC_163/Y 0.02fF
C21182 INVX1_LOC_510/Y INVX1_LOC_546/A 0.01fF
C21183 VDD INVX1_LOC_576/Y 0.21fF
C21184 INVX1_LOC_312/Y NAND2X1_LOC_475/A 0.64fF
C21185 INVX1_LOC_250/A INVX1_LOC_51/Y 0.01fF
C21186 NAND2X1_LOC_45/Y INVX1_LOC_486/Y 0.23fF
C21187 INVX1_LOC_479/A NAND2X1_LOC_832/A 0.04fF
C21188 INVX1_LOC_62/Y INVX1_LOC_231/Y 0.20fF
C21189 INVX1_LOC_41/Y NAND2X1_LOC_60/Y 0.01fF
C21190 INVX1_LOC_409/Y INVX1_LOC_116/Y 0.00fF
C21191 INVX1_LOC_601/A INVX1_LOC_197/Y 0.00fF
C21192 INVX1_LOC_206/Y NAND2X1_LOC_363/a_36_24# 0.01fF
C21193 NAND2X1_LOC_322/Y INVX1_LOC_116/Y 0.02fF
C21194 INVX1_LOC_405/A INVX1_LOC_48/Y 0.03fF
C21195 INVX1_LOC_51/Y INVX1_LOC_76/Y 0.06fF
C21196 INVX1_LOC_85/Y INVX1_LOC_191/A 0.54fF
C21197 VDD INVX1_LOC_662/Y 0.86fF
C21198 NAND2X1_LOC_482/Y INVX1_LOC_220/A 0.18fF
C21199 INVX1_LOC_266/A INVX1_LOC_76/Y 0.00fF
C21200 INVX1_LOC_412/Y INVX1_LOC_360/Y -0.00fF
C21201 INVX1_LOC_395/A INVX1_LOC_7/Y 0.73fF
C21202 INVX1_LOC_560/Y INVX1_LOC_48/Y 0.46fF
C21203 INVX1_LOC_315/Y INVX1_LOC_53/Y 0.03fF
C21204 INVX1_LOC_140/Y INVX1_LOC_99/Y 0.36fF
C21205 INVX1_LOC_618/A INVX1_LOC_49/Y 0.04fF
C21206 INVX1_LOC_20/Y INVX1_LOC_602/A 0.06fF
C21207 NAND2X1_LOC_498/Y INVX1_LOC_252/A 0.01fF
C21208 INVX1_LOC_442/A NAND2X1_LOC_369/a_36_24# 0.00fF
C21209 INVX1_LOC_231/Y NAND2X1_LOC_269/a_36_24# 0.00fF
C21210 INVX1_LOC_547/A INVX1_LOC_80/A 0.07fF
C21211 NAND2X1_LOC_526/Y INVX1_LOC_17/Y 0.01fF
C21212 NAND2X1_LOC_543/B INVX1_LOC_69/Y 0.15fF
C21213 NAND2X1_LOC_179/Y INVX1_LOC_45/Y 0.01fF
C21214 INVX1_LOC_409/Y INVX1_LOC_255/A 0.03fF
C21215 NAND2X1_LOC_69/B INVX1_LOC_63/Y 0.02fF
C21216 INVX1_LOC_10/Y INPUT_2 0.01fF
C21217 INVX1_LOC_581/A NAND2X1_LOC_783/a_36_24# 0.00fF
C21218 INVX1_LOC_278/A INVX1_LOC_671/A 0.09fF
C21219 INVX1_LOC_220/Y INVX1_LOC_385/Y 0.01fF
C21220 INVX1_LOC_361/Y NAND2X1_LOC_314/a_36_24# 0.00fF
C21221 INVX1_LOC_559/A INVX1_LOC_51/Y 0.01fF
C21222 INVX1_LOC_582/Y NAND2X1_LOC_679/B 0.01fF
C21223 INVX1_LOC_465/Y NAND2X1_LOC_686/B 0.02fF
C21224 INVX1_LOC_463/A INVX1_LOC_49/Y 0.08fF
C21225 INVX1_LOC_587/A INVX1_LOC_99/Y 0.00fF
C21226 INVX1_LOC_410/Y INVX1_LOC_103/Y 0.03fF
C21227 NAND2X1_LOC_45/Y INVX1_LOC_6/Y 5.09fF
C21228 INVX1_LOC_686/A INVX1_LOC_519/A 0.00fF
C21229 INVX1_LOC_435/Y INVX1_LOC_54/Y 0.72fF
C21230 VDD INVX1_LOC_646/Y 0.21fF
C21231 INVX1_LOC_395/A INVX1_LOC_32/Y 0.11fF
C21232 INVX1_LOC_96/Y NAND2X1_LOC_165/Y 0.19fF
C21233 INVX1_LOC_445/Y INVX1_LOC_6/Y 0.02fF
C21234 INVX1_LOC_451/A INPUT_2 0.17fF
C21235 INVX1_LOC_280/Y INVX1_LOC_45/Y 0.01fF
C21236 INVX1_LOC_11/Y INVX1_LOC_547/A 0.02fF
C21237 INVX1_LOC_21/Y INVX1_LOC_53/Y 0.49fF
C21238 INVX1_LOC_36/A INVX1_LOC_6/Y 0.02fF
C21239 INVX1_LOC_428/A INVX1_LOC_391/A 0.02fF
C21240 INVX1_LOC_362/Y INVX1_LOC_32/Y 0.05fF
C21241 NAND2X1_LOC_231/A NAND2X1_LOC_387/Y 0.01fF
C21242 INVX1_LOC_525/Y NAND2X1_LOC_506/B 0.07fF
C21243 INVX1_LOC_134/Y NAND2X1_LOC_418/Y 0.08fF
C21244 INVX1_LOC_431/A INVX1_LOC_169/A 0.02fF
C21245 INVX1_LOC_153/A INVX1_LOC_586/A 0.05fF
C21246 INVX1_LOC_570/A INVX1_LOC_6/Y 0.06fF
C21247 INVX1_LOC_395/A NAND2X1_LOC_286/A 0.03fF
C21248 NAND2X1_LOC_148/B INVX1_LOC_131/Y 0.01fF
C21249 INVX1_LOC_293/Y NAND2X1_LOC_106/B 0.81fF
C21250 INVX1_LOC_51/Y INVX1_LOC_108/A 0.03fF
C21251 INVX1_LOC_525/Y INVX1_LOC_45/Y 0.02fF
C21252 VDD INVX1_LOC_273/Y 0.36fF
C21253 NAND2X1_LOC_307/A INVX1_LOC_35/Y 0.04fF
C21254 INVX1_LOC_429/Y NAND2X1_LOC_344/B 0.01fF
C21255 INVX1_LOC_176/Y INVX1_LOC_171/A 0.00fF
C21256 INVX1_LOC_566/A INVX1_LOC_156/A 0.11fF
C21257 NAND2X1_LOC_520/B INVX1_LOC_69/Y 0.01fF
C21258 INVX1_LOC_355/A INVX1_LOC_49/Y 0.00fF
C21259 INVX1_LOC_84/A INVX1_LOC_48/Y 0.25fF
C21260 INVX1_LOC_20/Y INVX1_LOC_117/Y 0.25fF
C21261 INVX1_LOC_417/Y INVX1_LOC_129/A 0.01fF
C21262 INVX1_LOC_203/Y INVX1_LOC_90/Y 0.08fF
C21263 INPUT_3 INVX1_LOC_280/Y 0.01fF
C21264 INVX1_LOC_85/Y INVX1_LOC_182/Y 0.01fF
C21265 INVX1_LOC_586/A INVX1_LOC_96/A 0.05fF
C21266 INVX1_LOC_319/Y INVX1_LOC_9/Y 0.03fF
C21267 NAND2X1_LOC_369/a_36_24# INVX1_LOC_116/Y 0.00fF
C21268 NAND2X1_LOC_56/Y NAND2X1_LOC_615/B 0.04fF
C21269 INVX1_LOC_278/A INVX1_LOC_664/Y 0.01fF
C21270 INVX1_LOC_372/Y INVX1_LOC_359/Y 0.04fF
C21271 INVX1_LOC_145/Y INVX1_LOC_1/Y 0.01fF
C21272 INVX1_LOC_295/A INVX1_LOC_230/Y 0.11fF
C21273 INVX1_LOC_442/Y INVX1_LOC_453/Y 0.03fF
C21274 INVX1_LOC_137/Y INVX1_LOC_338/A 0.00fF
C21275 NAND2X1_LOC_65/a_36_24# INVX1_LOC_63/Y 0.00fF
C21276 INVX1_LOC_54/Y NAND2X1_LOC_318/B 1.35fF
C21277 INVX1_LOC_288/A INVX1_LOC_245/A 0.07fF
C21278 INVX1_LOC_567/Y INVX1_LOC_50/Y 0.01fF
C21279 INVX1_LOC_290/A INVX1_LOC_259/Y 0.03fF
C21280 INVX1_LOC_21/Y INVX1_LOC_43/A 0.01fF
C21281 INVX1_LOC_68/Y INVX1_LOC_179/A 0.19fF
C21282 INVX1_LOC_54/Y INVX1_LOC_366/Y 0.01fF
C21283 INVX1_LOC_411/A INVX1_LOC_230/A 0.05fF
C21284 INVX1_LOC_416/A INVX1_LOC_304/A 0.01fF
C21285 INVX1_LOC_419/Y INVX1_LOC_35/Y 0.07fF
C21286 INVX1_LOC_53/Y INVX1_LOC_555/A 0.15fF
C21287 INVX1_LOC_48/Y NAND2X1_LOC_67/Y 0.01fF
C21288 INVX1_LOC_93/Y INVX1_LOC_130/Y 0.01fF
C21289 NAND2X1_LOC_513/A INVX1_LOC_627/Y 0.01fF
C21290 INPUT_0 NAND2X1_LOC_689/a_36_24# 0.00fF
C21291 INVX1_LOC_11/Y NAND2X1_LOC_190/A 0.06fF
C21292 NAND2X1_LOC_710/A INVX1_LOC_63/Y 0.01fF
C21293 INVX1_LOC_230/A INVX1_LOC_295/Y 0.11fF
C21294 INVX1_LOC_300/A INVX1_LOC_117/Y 0.15fF
C21295 INVX1_LOC_84/A NAND2X1_LOC_491/Y 0.03fF
C21296 INVX1_LOC_304/Y INVX1_LOC_159/Y 1.40fF
C21297 INVX1_LOC_21/Y NAND2X1_LOC_400/B 0.29fF
C21298 INVX1_LOC_81/Y INVX1_LOC_195/Y 0.01fF
C21299 INVX1_LOC_31/Y INVX1_LOC_7/Y 0.01fF
C21300 INVX1_LOC_235/Y INVX1_LOC_328/Y 0.07fF
C21301 INVX1_LOC_80/A INVX1_LOC_624/Y 0.05fF
C21302 NAND2X1_LOC_65/Y NAND2X1_LOC_786/B 0.03fF
C21303 NAND2X1_LOC_638/A INVX1_LOC_69/Y 0.03fF
C21304 INVX1_LOC_507/Y INVX1_LOC_492/Y 0.03fF
C21305 INVX1_LOC_17/Y NAND2X1_LOC_619/Y 0.02fF
C21306 INVX1_LOC_93/Y NAND2X1_LOC_210/A 0.01fF
C21307 INVX1_LOC_53/Y INVX1_LOC_107/Y 0.03fF
C21308 INVX1_LOC_99/Y INVX1_LOC_6/Y 2.22fF
C21309 NAND2X1_LOC_79/Y INVX1_LOC_26/Y 0.16fF
C21310 INVX1_LOC_578/Y INVX1_LOC_259/Y 0.17fF
C21311 INVX1_LOC_169/A NAND2X1_LOC_489/A -0.00fF
C21312 INVX1_LOC_159/Y NAND2X1_LOC_444/A 0.03fF
C21313 INVX1_LOC_609/A INVX1_LOC_6/Y 0.17fF
C21314 INVX1_LOC_89/Y INVX1_LOC_98/Y 0.33fF
C21315 INVX1_LOC_47/Y INVX1_LOC_252/A 0.04fF
C21316 INVX1_LOC_607/Y INVX1_LOC_520/Y 0.05fF
C21317 INVX1_LOC_491/Y INVX1_LOC_496/A 0.07fF
C21318 INVX1_LOC_285/A INVX1_LOC_26/Y 0.03fF
C21319 INVX1_LOC_179/A INVX1_LOC_600/A 0.07fF
C21320 INVX1_LOC_35/Y NAND2X1_LOC_342/A 0.01fF
C21321 INVX1_LOC_93/Y INVX1_LOC_110/A 0.01fF
C21322 INVX1_LOC_31/Y INVX1_LOC_345/Y 0.03fF
C21323 NAND2X1_LOC_106/Y INVX1_LOC_50/Y 0.00fF
C21324 INVX1_LOC_69/Y INVX1_LOC_505/A 1.29fF
C21325 INVX1_LOC_532/Y INVX1_LOC_259/Y 0.09fF
C21326 INVX1_LOC_31/Y INVX1_LOC_32/Y 1.65fF
C21327 INVX1_LOC_17/Y NAND2X1_LOC_618/a_36_24# 0.00fF
C21328 INVX1_LOC_478/Y INVX1_LOC_77/Y 0.01fF
C21329 INVX1_LOC_202/Y INVX1_LOC_361/A 0.02fF
C21330 INVX1_LOC_566/Y INVX1_LOC_62/Y 0.01fF
C21331 INVX1_LOC_63/Y NAND2X1_LOC_226/a_36_24# 0.00fF
C21332 INVX1_LOC_432/Y INVX1_LOC_9/Y 0.03fF
C21333 INVX1_LOC_551/Y NAND2X1_LOC_410/Y 0.14fF
C21334 INVX1_LOC_496/A INVX1_LOC_48/Y 0.07fF
C21335 INVX1_LOC_145/Y INVX1_LOC_245/A 0.06fF
C21336 INVX1_LOC_402/A NAND2X1_LOC_136/Y 0.42fF
C21337 INVX1_LOC_385/Y INVX1_LOC_244/Y 0.03fF
C21338 INVX1_LOC_47/Y NAND2X1_LOC_688/a_36_24# 0.01fF
C21339 INVX1_LOC_119/Y INVX1_LOC_252/A 0.03fF
C21340 INVX1_LOC_659/A INVX1_LOC_342/A 0.09fF
C21341 INVX1_LOC_47/Y INVX1_LOC_6/Y 0.13fF
C21342 NAND2X1_LOC_557/B INVX1_LOC_6/Y 0.25fF
C21343 INVX1_LOC_134/A INVX1_LOC_92/A 0.16fF
C21344 INVX1_LOC_194/Y INVX1_LOC_90/Y 0.07fF
C21345 INVX1_LOC_187/Y INVX1_LOC_188/A 0.03fF
C21346 INVX1_LOC_344/Y INVX1_LOC_74/Y 0.00fF
C21347 INVX1_LOC_507/Y NAND2X1_LOC_647/A 0.00fF
C21348 INVX1_LOC_662/A NAND2X1_LOC_286/a_36_24# 0.01fF
C21349 INVX1_LOC_487/Y INPUT_1 0.18fF
C21350 NAND2X1_LOC_544/B INVX1_LOC_98/Y 0.10fF
C21351 NAND2X1_LOC_123/B INVX1_LOC_50/Y 0.00fF
C21352 INVX1_LOC_367/Y NAND2X1_LOC_844/A 0.03fF
C21353 INVX1_LOC_507/Y INVX1_LOC_168/Y 0.14fF
C21354 INVX1_LOC_674/A INVX1_LOC_635/Y 0.02fF
C21355 INVX1_LOC_560/A INVX1_LOC_109/Y 0.02fF
C21356 NAND2X1_LOC_532/Y INVX1_LOC_79/A 0.00fF
C21357 INVX1_LOC_199/Y INVX1_LOC_26/Y 0.00fF
C21358 INVX1_LOC_6/Y NAND2X1_LOC_66/Y 0.52fF
C21359 INVX1_LOC_58/Y INVX1_LOC_242/Y 0.07fF
C21360 INVX1_LOC_166/A INVX1_LOC_653/Y 0.00fF
C21361 INVX1_LOC_97/A INVX1_LOC_615/A 0.04fF
C21362 NAND2X1_LOC_494/a_36_24# INVX1_LOC_9/Y 0.00fF
C21363 INVX1_LOC_471/Y INVX1_LOC_114/A 0.04fF
C21364 INVX1_LOC_319/A INVX1_LOC_9/Y 0.07fF
C21365 INVX1_LOC_26/Y INVX1_LOC_85/A 0.56fF
C21366 INVX1_LOC_50/Y INVX1_LOC_92/A 0.06fF
C21367 NAND2X1_LOC_843/B INVX1_LOC_9/Y 0.26fF
C21368 INVX1_LOC_183/A NAND2X1_LOC_617/a_36_24# 0.00fF
C21369 NAND2X1_LOC_770/A INVX1_LOC_51/Y 0.01fF
C21370 NAND2X1_LOC_543/B INVX1_LOC_586/A 0.91fF
C21371 INVX1_LOC_62/Y INVX1_LOC_319/A 0.03fF
C21372 NAND2X1_LOC_520/A NAND2X1_LOC_271/A 0.04fF
C21373 NAND2X1_LOC_707/a_36_24# INVX1_LOC_139/A 0.00fF
C21374 INVX1_LOC_412/Y INVX1_LOC_45/Y 0.03fF
C21375 INVX1_LOC_230/A NAND2X1_LOC_216/a_36_24# 0.01fF
C21376 INVX1_LOC_224/Y NAND2X1_LOC_391/B 0.03fF
C21377 INVX1_LOC_62/Y INVX1_LOC_625/Y 0.02fF
C21378 INVX1_LOC_601/A INVX1_LOC_600/Y 0.01fF
C21379 NAND2X1_LOC_520/B INVX1_LOC_586/A 0.01fF
C21380 INVX1_LOC_286/A NAND2X1_LOC_352/a_36_24# 0.02fF
C21381 NAND2X1_LOC_750/Y INVX1_LOC_12/Y 0.06fF
C21382 INVX1_LOC_301/A NAND2X1_LOC_143/a_36_24# 0.00fF
C21383 VDD INVX1_LOC_70/Y 0.21fF
C21384 INVX1_LOC_35/Y INVX1_LOC_388/Y 0.03fF
C21385 INVX1_LOC_558/A INVX1_LOC_551/Y 0.01fF
C21386 INVX1_LOC_176/Y INVX1_LOC_45/Y 0.00fF
C21387 INVX1_LOC_442/Y NAND2X1_LOC_457/A 0.01fF
C21388 NAND2X1_LOC_13/Y INVX1_LOC_76/Y 0.06fF
C21389 INVX1_LOC_380/Y INVX1_LOC_297/Y 0.01fF
C21390 INVX1_LOC_395/A INVX1_LOC_130/Y 0.04fF
C21391 INVX1_LOC_254/Y VDD 0.36fF
C21392 INPUT_0 INVX1_LOC_201/Y 0.01fF
C21393 INVX1_LOC_551/Y INVX1_LOC_270/A 0.47fF
C21394 INVX1_LOC_452/A INVX1_LOC_445/A 0.40fF
C21395 NAND2X1_LOC_638/A INVX1_LOC_586/A 0.03fF
C21396 INVX1_LOC_53/Y INVX1_LOC_577/Y 0.03fF
C21397 INVX1_LOC_206/Y INVX1_LOC_513/A 0.02fF
C21398 INVX1_LOC_182/A INVX1_LOC_145/Y 0.02fF
C21399 INVX1_LOC_560/Y INVX1_LOC_559/Y 0.19fF
C21400 INVX1_LOC_409/Y INVX1_LOC_69/Y 0.12fF
C21401 INVX1_LOC_522/Y INVX1_LOC_492/Y 0.02fF
C21402 INVX1_LOC_254/Y INVX1_LOC_228/Y 0.02fF
C21403 NAND2X1_LOC_322/Y INVX1_LOC_69/Y 0.01fF
C21404 VDD INVX1_LOC_592/Y 0.40fF
C21405 INPUT_0 INVX1_LOC_543/Y 0.02fF
C21406 INVX1_LOC_435/Y INVX1_LOC_277/A 0.05fF
C21407 INVX1_LOC_401/A NAND2X1_LOC_513/A 0.07fF
C21408 INVX1_LOC_428/Y INVX1_LOC_427/A 0.01fF
C21409 INVX1_LOC_587/A INVX1_LOC_25/Y 0.01fF
C21410 INVX1_LOC_255/Y INVX1_LOC_460/Y 0.01fF
C21411 INPUT_0 NAND2X1_LOC_547/a_36_24# 0.01fF
C21412 INVX1_LOC_586/A INVX1_LOC_505/A 0.03fF
C21413 INVX1_LOC_310/Y INVX1_LOC_63/A 0.15fF
C21414 VDD INVX1_LOC_309/Y 0.21fF
C21415 INVX1_LOC_20/Y INVX1_LOC_178/A 0.07fF
C21416 INVX1_LOC_445/Y NAND2X1_LOC_294/Y 0.02fF
C21417 INVX1_LOC_53/Y INVX1_LOC_474/Y 0.21fF
C21418 NAND2X1_LOC_505/Y INVX1_LOC_32/Y 0.13fF
C21419 INVX1_LOC_51/Y INVX1_LOC_345/Y 0.03fF
C21420 INVX1_LOC_185/A INVX1_LOC_655/A 0.02fF
C21421 INVX1_LOC_218/Y INVX1_LOC_384/A 0.04fF
C21422 INVX1_LOC_134/A INPUT_1 0.01fF
C21423 INVX1_LOC_560/A INVX1_LOC_199/Y 0.07fF
C21424 INVX1_LOC_365/Y INVX1_LOC_7/Y 0.04fF
C21425 INVX1_LOC_51/Y INVX1_LOC_32/Y 1.61fF
C21426 NAND2X1_LOC_97/B INVX1_LOC_160/A 0.02fF
C21427 INVX1_LOC_223/Y NAND2X1_LOC_749/Y 0.51fF
C21428 NAND2X1_LOC_123/A NAND2X1_LOC_117/a_36_24# 0.02fF
C21429 INVX1_LOC_266/A INVX1_LOC_32/Y 0.03fF
C21430 INVX1_LOC_551/Y INVX1_LOC_46/Y 0.03fF
C21431 INVX1_LOC_68/Y INVX1_LOC_69/Y 0.05fF
C21432 INVX1_LOC_233/Y INVX1_LOC_69/Y 0.01fF
C21433 INVX1_LOC_76/Y INVX1_LOC_380/Y 0.02fF
C21434 INVX1_LOC_17/Y INVX1_LOC_379/A 0.06fF
C21435 VDD NAND2X1_LOC_528/Y 0.52fF
C21436 NAND2X1_LOC_685/A INVX1_LOC_463/Y 0.03fF
C21437 GATE_865 INVX1_LOC_632/A 0.21fF
C21438 INVX1_LOC_612/Y NAND2X1_LOC_513/A 0.02fF
C21439 INVX1_LOC_201/A INVX1_LOC_201/Y 0.16fF
C21440 INVX1_LOC_76/Y INVX1_LOC_361/A 0.03fF
C21441 INVX1_LOC_581/A INVX1_LOC_535/Y 0.05fF
C21442 INVX1_LOC_522/Y NAND2X1_LOC_647/A 0.01fF
C21443 INVX1_LOC_384/A NAND2X1_LOC_256/a_36_24# 0.01fF
C21444 INVX1_LOC_193/A INVX1_LOC_417/Y 0.01fF
C21445 INVX1_LOC_54/Y INVX1_LOC_530/A 0.19fF
C21446 INVX1_LOC_17/Y INVX1_LOC_35/Y 13.72fF
C21447 VDD INVX1_LOC_479/A 4.50fF
C21448 NAND2X1_LOC_299/Y INVX1_LOC_93/Y 2.03fF
C21449 INVX1_LOC_435/A NAND2X1_LOC_561/a_36_24# 0.00fF
C21450 INVX1_LOC_20/Y INVX1_LOC_58/Y 0.22fF
C21451 INVX1_LOC_400/Y INVX1_LOC_100/Y 0.07fF
C21452 INVX1_LOC_76/Y INVX1_LOC_196/Y 0.01fF
C21453 NAND2X1_LOC_638/A NAND2X1_LOC_835/A 0.02fF
C21454 INVX1_LOC_393/Y INVX1_LOC_62/Y 0.11fF
C21455 INVX1_LOC_586/A INVX1_LOC_353/A 0.03fF
C21456 INVX1_LOC_584/A INVX1_LOC_74/Y 0.16fF
C21457 INPUT_0 INVX1_LOC_652/Y 0.02fF
C21458 INVX1_LOC_522/Y INVX1_LOC_168/Y 0.46fF
C21459 INVX1_LOC_558/Y INVX1_LOC_66/A 0.01fF
C21460 NAND2X1_LOC_596/Y INVX1_LOC_479/A 0.06fF
C21461 INVX1_LOC_256/Y INVX1_LOC_376/A 0.05fF
C21462 INVX1_LOC_84/A NAND2X1_LOC_615/Y 0.08fF
C21463 NAND2X1_LOC_707/A INVX1_LOC_114/A 0.00fF
C21464 INVX1_LOC_228/Y INVX1_LOC_479/A 0.17fF
C21465 NAND2X1_LOC_184/Y INVX1_LOC_392/A 0.03fF
C21466 NAND2X1_LOC_299/Y INVX1_LOC_675/A 0.01fF
C21467 INVX1_LOC_69/Y INVX1_LOC_600/A 0.10fF
C21468 INVX1_LOC_235/Y INVX1_LOC_224/A 0.03fF
C21469 INVX1_LOC_300/A INVX1_LOC_157/A 0.03fF
C21470 NAND2X1_LOC_360/a_36_24# INVX1_LOC_50/Y 0.00fF
C21471 INVX1_LOC_17/Y NAND2X1_LOC_253/Y 0.07fF
C21472 NAND2X1_LOC_43/Y INVX1_LOC_6/Y 0.01fF
C21473 INPUT_1 INVX1_LOC_50/Y 12.26fF
C21474 INVX1_LOC_20/Y NAND2X1_LOC_342/B 0.32fF
C21475 INVX1_LOC_558/A NAND2X1_LOC_410/Y 0.04fF
C21476 NAND2X1_LOC_307/B INVX1_LOC_35/Y 0.00fF
C21477 INVX1_LOC_300/A INVX1_LOC_58/Y 0.27fF
C21478 INVX1_LOC_510/Y INVX1_LOC_479/A 0.28fF
C21479 INVX1_LOC_53/Y INVX1_LOC_26/Y 6.39fF
C21480 INVX1_LOC_254/A INVX1_LOC_32/Y 0.00fF
C21481 INVX1_LOC_80/A NAND2X1_LOC_833/B 0.16fF
C21482 INVX1_LOC_31/Y INVX1_LOC_110/A 0.04fF
C21483 NAND2X1_LOC_184/Y INVX1_LOC_93/Y 0.05fF
C21484 INVX1_LOC_58/Y INVX1_LOC_197/Y 0.01fF
C21485 INVX1_LOC_527/Y NAND2X1_LOC_753/Y 0.02fF
C21486 INVX1_LOC_504/A INVX1_LOC_501/A 0.07fF
C21487 NAND2X1_LOC_192/A INVX1_LOC_99/Y 0.01fF
C21488 INVX1_LOC_400/A INVX1_LOC_551/A 0.01fF
C21489 INVX1_LOC_137/Y INVX1_LOC_507/Y 0.07fF
C21490 NAND2X1_LOC_179/a_36_24# INVX1_LOC_116/Y 0.00fF
C21491 INVX1_LOC_551/Y INVX1_LOC_75/A 0.01fF
C21492 INVX1_LOC_513/A NAND2X1_LOC_334/A 0.03fF
C21493 INVX1_LOC_293/Y NAND2X1_LOC_248/B 0.01fF
C21494 INVX1_LOC_50/Y NAND2X1_LOC_279/a_36_24# 0.01fF
C21495 INVX1_LOC_344/Y INVX1_LOC_79/A 0.07fF
C21496 INVX1_LOC_50/Y INVX1_LOC_284/Y 0.16fF
C21497 INVX1_LOC_549/Y INVX1_LOC_491/A 0.02fF
C21498 INVX1_LOC_97/Y INVX1_LOC_531/Y 0.05fF
C21499 INVX1_LOC_281/Y NAND2X1_LOC_269/B 0.01fF
C21500 INVX1_LOC_31/Y NAND2X1_LOC_275/a_36_24# 0.01fF
C21501 NAND2X1_LOC_137/A INVX1_LOC_544/Y 0.01fF
C21502 INVX1_LOC_11/Y NAND2X1_LOC_833/B 0.72fF
C21503 INVX1_LOC_361/Y INVX1_LOC_9/Y 0.06fF
C21504 INVX1_LOC_508/A NAND2X1_LOC_647/A 0.06fF
C21505 NAND2X1_LOC_683/a_36_24# INVX1_LOC_50/Y 0.00fF
C21506 NAND2X1_LOC_297/Y INVX1_LOC_245/A 0.01fF
C21507 INVX1_LOC_62/Y NAND2X1_LOC_678/a_36_24# 0.00fF
C21508 INVX1_LOC_368/A INVX1_LOC_50/Y 0.04fF
C21509 INVX1_LOC_283/Y INVX1_LOC_293/A 0.03fF
C21510 NAND2X1_LOC_597/Y INVX1_LOC_145/Y 0.02fF
C21511 INVX1_LOC_537/A INVX1_LOC_74/Y 0.03fF
C21512 INVX1_LOC_49/Y NAND2X1_LOC_449/B 0.06fF
C21513 NAND2X1_LOC_770/B INVX1_LOC_79/A 0.01fF
C21514 INVX1_LOC_555/A INVX1_LOC_662/A 0.07fF
C21515 INVX1_LOC_49/Y INVX1_LOC_480/A 0.03fF
C21516 NAND2X1_LOC_555/B NAND2X1_LOC_344/B 0.03fF
C21517 INVX1_LOC_400/A INVX1_LOC_75/Y 0.00fF
C21518 INVX1_LOC_479/A INVX1_LOC_509/A 0.01fF
C21519 INVX1_LOC_557/Y INVX1_LOC_47/Y 0.02fF
C21520 NAND2X1_LOC_409/Y INVX1_LOC_48/Y 0.09fF
C21521 INVX1_LOC_164/Y INVX1_LOC_62/Y 0.21fF
C21522 NAND2X1_LOC_294/Y NAND2X1_LOC_66/Y 0.10fF
C21523 INVX1_LOC_361/Y INVX1_LOC_62/Y 0.19fF
C21524 NAND2X1_LOC_827/a_36_24# INVX1_LOC_50/Y 0.00fF
C21525 INVX1_LOC_26/Y NAND2X1_LOC_274/Y 0.00fF
C21526 INVX1_LOC_6/Y NAND2X1_LOC_627/Y 0.01fF
C21527 INVX1_LOC_58/Y INVX1_LOC_655/A 0.02fF
C21528 INVX1_LOC_93/Y INVX1_LOC_75/Y 0.21fF
C21529 INVX1_LOC_437/A INVX1_LOC_443/A 0.14fF
C21530 INVX1_LOC_94/Y INVX1_LOC_531/Y 0.14fF
C21531 INVX1_LOC_99/Y INVX1_LOC_636/A 0.46fF
C21532 INVX1_LOC_26/Y NAND2X1_LOC_406/B 0.01fF
C21533 INVX1_LOC_261/Y INVX1_LOC_62/Y 0.03fF
C21534 INVX1_LOC_557/Y INVX1_LOC_119/Y 0.00fF
C21535 INVX1_LOC_235/Y INVX1_LOC_109/Y 0.10fF
C21536 INVX1_LOC_666/Y INVX1_LOC_411/Y 0.01fF
C21537 INVX1_LOC_93/Y NAND2X1_LOC_271/A 0.20fF
C21538 INVX1_LOC_100/Y NAND2X1_LOC_814/a_36_24# 0.00fF
C21539 INVX1_LOC_655/A NAND2X1_LOC_342/B 0.03fF
C21540 NAND2X1_LOC_170/a_36_24# INVX1_LOC_271/A 0.00fF
C21541 NAND2X1_LOC_781/B INVX1_LOC_586/A 0.01fF
C21542 NAND2X1_LOC_545/A INVX1_LOC_41/Y 0.09fF
C21543 NAND2X1_LOC_388/A INVX1_LOC_92/A 0.12fF
C21544 INVX1_LOC_420/Y INVX1_LOC_421/Y 0.15fF
C21545 INVX1_LOC_47/Y INVX1_LOC_636/A 0.01fF
C21546 INVX1_LOC_51/A NAND2X1_LOC_46/a_36_24# 0.02fF
C21547 NAND2X1_LOC_241/B INVX1_LOC_604/A 0.01fF
C21548 INVX1_LOC_41/Y INVX1_LOC_653/Y 0.73fF
C21549 NAND2X1_LOC_142/a_36_24# NAND2X1_LOC_142/Y 0.02fF
C21550 INVX1_LOC_41/Y INVX1_LOC_666/Y 0.10fF
C21551 NAND2X1_LOC_781/A NAND2X1_LOC_781/B 0.03fF
C21552 NAND2X1_LOC_45/Y INVX1_LOC_381/A 0.10fF
C21553 NAND2X1_LOC_636/A INVX1_LOC_633/Y 0.03fF
C21554 VDD INVX1_LOC_372/Y 0.44fF
C21555 NAND2X1_LOC_249/Y INVX1_LOC_53/Y 0.03fF
C21556 INVX1_LOC_241/A NAND2X1_LOC_287/a_36_24# 0.02fF
C21557 VDD INVX1_LOC_12/Y 1.29fF
C21558 INVX1_LOC_19/Y INVX1_LOC_29/Y 0.01fF
C21559 INVX1_LOC_276/A NAND2X1_LOC_108/Y 0.01fF
C21560 NAND2X1_LOC_97/A INVX1_LOC_94/A 0.15fF
C21561 INVX1_LOC_68/Y INVX1_LOC_586/A 0.03fF
C21562 INVX1_LOC_233/Y INVX1_LOC_586/A 0.02fF
C21563 INVX1_LOC_554/A INVX1_LOC_556/Y 1.25fF
C21564 INPUT_0 INVX1_LOC_197/A 0.29fF
C21565 INVX1_LOC_560/Y INVX1_LOC_155/Y 0.02fF
C21566 VDD INVX1_LOC_684/Y 0.21fF
C21567 INVX1_LOC_586/A INVX1_LOC_147/Y 0.01fF
C21568 INVX1_LOC_406/Y INVX1_LOC_45/Y 0.00fF
C21569 NAND2X1_LOC_88/B INVX1_LOC_182/A 0.01fF
C21570 NAND2X1_LOC_537/B INVX1_LOC_600/A -0.01fF
C21571 INVX1_LOC_211/Y INVX1_LOC_596/Y 0.01fF
C21572 INVX1_LOC_583/Y INVX1_LOC_522/Y 0.05fF
C21573 INVX1_LOC_228/Y INVX1_LOC_12/Y 0.05fF
C21574 NAND2X1_LOC_176/Y INVX1_LOC_98/Y 0.05fF
C21575 INVX1_LOC_20/Y NAND2X1_LOC_390/a_36_24# 0.00fF
C21576 INVX1_LOC_286/Y INVX1_LOC_291/A 0.00fF
C21577 INVX1_LOC_224/Y INVX1_LOC_435/A 0.12fF
C21578 INVX1_LOC_404/Y INVX1_LOC_367/Y 0.39fF
C21579 INVX1_LOC_438/A INVX1_LOC_681/Y 0.02fF
C21580 VDD INVX1_LOC_138/Y 0.21fF
C21581 NAND2X1_LOC_537/A INVX1_LOC_32/Y 0.01fF
C21582 INVX1_LOC_438/A INPUT_1 0.07fF
C21583 INVX1_LOC_586/A INVX1_LOC_600/A 0.07fF
C21584 INVX1_LOC_587/A NAND2X1_LOC_638/A 0.03fF
C21585 NAND2X1_LOC_790/B INVX1_LOC_199/Y 0.60fF
C21586 VDD NAND2X1_LOC_333/A 0.27fF
C21587 INVX1_LOC_282/A INVX1_LOC_445/A 0.11fF
C21588 VDD INVX1_LOC_391/A 0.00fF
C21589 INVX1_LOC_24/A INPUT_1 0.01fF
C21590 INVX1_LOC_206/Y INVX1_LOC_670/A 0.04fF
C21591 INVX1_LOC_89/Y NAND2X1_LOC_76/B 0.14fF
C21592 INVX1_LOC_563/Y INVX1_LOC_298/A 0.01fF
C21593 INVX1_LOC_154/A NAND2X1_LOC_76/B 0.06fF
C21594 INVX1_LOC_80/A INVX1_LOC_101/Y 0.01fF
C21595 VDD INVX1_LOC_188/A -0.00fF
C21596 INPUT_0 INVX1_LOC_173/Y 0.16fF
C21597 VDD INVX1_LOC_170/A 0.00fF
C21598 INVX1_LOC_381/A INVX1_LOC_99/Y 0.07fF
C21599 INVX1_LOC_355/A INVX1_LOC_345/Y 0.00fF
C21600 INVX1_LOC_54/Y INVX1_LOC_65/Y 0.03fF
C21601 INVX1_LOC_68/Y NAND2X1_LOC_74/a_36_24# 0.00fF
C21602 VDD INVX1_LOC_276/Y 0.21fF
C21603 NAND2X1_LOC_184/Y INVX1_LOC_362/Y 0.05fF
C21604 INVX1_LOC_197/A NAND2X1_LOC_123/A 0.05fF
C21605 INVX1_LOC_202/Y INVX1_LOC_551/Y 0.05fF
C21606 INVX1_LOC_523/A INVX1_LOC_477/Y 0.02fF
C21607 NAND2X1_LOC_180/B INVX1_LOC_159/Y 0.04fF
C21608 NAND2X1_LOC_532/Y NAND2X1_LOC_513/Y 0.03fF
C21609 INVX1_LOC_27/A INVX1_LOC_7/Y 0.31fF
C21610 INVX1_LOC_320/A INVX1_LOC_99/Y 0.00fF
C21611 INVX1_LOC_522/Y INVX1_LOC_137/Y 0.07fF
C21612 NAND2X1_LOC_336/B INVX1_LOC_194/A 0.00fF
C21613 INVX1_LOC_670/A INVX1_LOC_242/A 0.82fF
C21614 NAND2X1_LOC_750/Y INVX1_LOC_178/Y 0.06fF
C21615 VDD INVX1_LOC_488/A -0.00fF
C21616 INVX1_LOC_438/A INVX1_LOC_368/A 0.02fF
C21617 INVX1_LOC_526/A INVX1_LOC_498/A 0.12fF
C21618 INVX1_LOC_424/A NAND2X1_LOC_642/a_36_24# 0.00fF
C21619 VDD INVX1_LOC_680/A 0.00fF
C21620 INVX1_LOC_580/Y INVX1_LOC_261/Y 0.02fF
C21621 INVX1_LOC_17/Y INVX1_LOC_531/A 0.04fF
C21622 NAND2X1_LOC_45/Y INVX1_LOC_100/Y 0.12fF
C21623 NAND2X1_LOC_325/B NAND2X1_LOC_775/B 0.21fF
C21624 INVX1_LOC_614/A INVX1_LOC_138/Y 0.03fF
C21625 INVX1_LOC_607/Y NAND2X1_LOC_285/B 0.02fF
C21626 INVX1_LOC_608/Y INVX1_LOC_214/Y 0.08fF
C21627 NAND2X1_LOC_513/A INPUT_1 4.06fF
C21628 INVX1_LOC_511/Y INVX1_LOC_330/A 0.00fF
C21629 INVX1_LOC_607/Y NAND2X1_LOC_106/B 0.18fF
C21630 INVX1_LOC_378/A INVX1_LOC_379/Y 0.01fF
C21631 INVX1_LOC_51/Y NAND2X1_LOC_405/a_36_24# 0.01fF
C21632 INVX1_LOC_400/Y INVX1_LOC_79/A 0.03fF
C21633 INVX1_LOC_551/Y INVX1_LOC_49/Y 0.10fF
C21634 INVX1_LOC_567/Y INVX1_LOC_117/Y 0.02fF
C21635 INVX1_LOC_20/Y NAND2X1_LOC_91/a_36_24# 0.00fF
C21636 INVX1_LOC_80/A NAND2X1_LOC_308/A 0.42fF
C21637 NAND2X1_LOC_498/Y INVX1_LOC_100/Y 0.08fF
C21638 INVX1_LOC_17/Y INVX1_LOC_360/A 0.00fF
C21639 INVX1_LOC_439/Y INVX1_LOC_444/Y 0.03fF
C21640 NAND2X1_LOC_45/Y INVX1_LOC_483/Y 0.06fF
C21641 INVX1_LOC_312/Y NAND2X1_LOC_613/a_36_24# 0.00fF
C21642 INVX1_LOC_134/Y INVX1_LOC_234/Y 0.04fF
C21643 INVX1_LOC_543/Y INVX1_LOC_145/Y 3.28fF
C21644 INVX1_LOC_11/Y INVX1_LOC_665/Y 0.03fF
C21645 INVX1_LOC_35/Y INVX1_LOC_189/A 0.01fF
C21646 VDD INVX1_LOC_212/A 0.00fF
C21647 INVX1_LOC_379/A INVX1_LOC_230/Y 0.02fF
C21648 INVX1_LOC_20/Y INVX1_LOC_245/A 0.61fF
C21649 INVX1_LOC_395/A INVX1_LOC_75/Y 0.08fF
C21650 INVX1_LOC_99/Y INVX1_LOC_470/Y 0.01fF
C21651 NAND2X1_LOC_413/Y INVX1_LOC_66/A 0.20fF
C21652 INVX1_LOC_35/Y INVX1_LOC_230/Y 0.07fF
C21653 INVX1_LOC_541/Y INVX1_LOC_501/A 0.34fF
C21654 NAND2X1_LOC_498/Y INVX1_LOC_74/Y 0.08fF
C21655 NAND2X1_LOC_534/a_36_24# INVX1_LOC_376/Y 0.00fF
C21656 INVX1_LOC_21/Y NAND2X1_LOC_178/a_36_24# 0.06fF
C21657 INVX1_LOC_570/A INVX1_LOC_74/Y 0.03fF
C21658 NAND2X1_LOC_858/a_36_24# INVX1_LOC_283/A 0.00fF
C21659 INVX1_LOC_438/Y INVX1_LOC_443/A 0.12fF
C21660 INVX1_LOC_293/Y INVX1_LOC_664/A 0.03fF
C21661 INVX1_LOC_625/A INVX1_LOC_89/Y 0.04fF
C21662 NAND2X1_LOC_318/B INVX1_LOC_44/Y 0.02fF
C21663 INVX1_LOC_650/Y INVX1_LOC_649/A 0.19fF
C21664 INVX1_LOC_54/Y INVX1_LOC_318/A 0.02fF
C21665 INVX1_LOC_11/Y NAND2X1_LOC_308/A 0.21fF
C21666 INVX1_LOC_114/Y INVX1_LOC_74/Y 0.01fF
C21667 INVX1_LOC_353/Y INVX1_LOC_41/Y 0.04fF
C21668 NAND2X1_LOC_475/A INVX1_LOC_636/A 0.02fF
C21669 INVX1_LOC_556/Y INVX1_LOC_199/Y 0.06fF
C21670 INVX1_LOC_176/A INVX1_LOC_63/Y 0.06fF
C21671 INVX1_LOC_660/Y INVX1_LOC_59/A 0.28fF
C21672 INVX1_LOC_297/A INVX1_LOC_90/Y 0.00fF
C21673 NAND2X1_LOC_106/Y INVX1_LOC_117/Y 0.03fF
C21674 NAND2X1_LOC_184/Y INVX1_LOC_31/Y 0.00fF
C21675 INVX1_LOC_12/Y NAND2X1_LOC_786/B 0.65fF
C21676 NAND2X1_LOC_388/A INPUT_1 0.02fF
C21677 INVX1_LOC_53/Y NAND2X1_LOC_626/Y 0.05fF
C21678 NAND2X1_LOC_179/Y INVX1_LOC_682/A 0.04fF
C21679 INVX1_LOC_89/Y INVX1_LOC_520/A 0.02fF
C21680 INVX1_LOC_177/A INVX1_LOC_44/Y 0.03fF
C21681 INVX1_LOC_315/A NAND2X1_LOC_836/B 0.04fF
C21682 INVX1_LOC_300/A INVX1_LOC_245/A 0.08fF
C21683 INVX1_LOC_270/A INVX1_LOC_75/A 0.10fF
C21684 INVX1_LOC_197/Y INVX1_LOC_245/A 0.03fF
C21685 INVX1_LOC_261/Y INVX1_LOC_641/Y 0.03fF
C21686 NAND2X1_LOC_136/Y NAND2X1_LOC_284/a_36_24# -0.00fF
C21687 INVX1_LOC_517/Y INVX1_LOC_50/Y 0.07fF
C21688 INVX1_LOC_326/Y INVX1_LOC_6/Y 0.00fF
C21689 INVX1_LOC_83/Y INVX1_LOC_9/Y 0.24fF
C21690 INVX1_LOC_100/Y INVX1_LOC_99/Y 4.76fF
C21691 INVX1_LOC_81/Y INVX1_LOC_85/A 0.06fF
C21692 INVX1_LOC_442/Y INVX1_LOC_62/Y 0.07fF
C21693 INVX1_LOC_21/Y INVX1_LOC_653/Y 0.04fF
C21694 INVX1_LOC_524/Y NAND2X1_LOC_98/B 0.30fF
C21695 INVX1_LOC_455/A NAND2X1_LOC_836/a_36_24# 0.00fF
C21696 INVX1_LOC_21/Y INVX1_LOC_327/A 0.01fF
C21697 INVX1_LOC_99/Y INVX1_LOC_74/Y 0.10fF
C21698 NAND2X1_LOC_346/a_36_24# INVX1_LOC_49/Y 0.01fF
C21699 INVX1_LOC_149/Y INVX1_LOC_496/A 0.03fF
C21700 INVX1_LOC_391/Y INVX1_LOC_41/Y 0.00fF
C21701 INVX1_LOC_99/Y INVX1_LOC_483/Y 0.02fF
C21702 INVX1_LOC_17/Y INVX1_LOC_364/A 0.14fF
C21703 INVX1_LOC_117/Y NAND2X1_LOC_123/B 0.03fF
C21704 NAND2X1_LOC_187/Y INVX1_LOC_588/A 0.01fF
C21705 INVX1_LOC_399/Y INVX1_LOC_63/Y 0.00fF
C21706 INVX1_LOC_41/Y INVX1_LOC_18/Y 0.06fF
C21707 INVX1_LOC_183/A INVX1_LOC_328/Y 1.19fF
C21708 INVX1_LOC_124/A INVX1_LOC_63/Y 0.01fF
C21709 NAND2X1_LOC_192/A INVX1_LOC_15/Y 0.07fF
C21710 NAND2X1_LOC_686/A INVX1_LOC_501/A 0.00fF
C21711 INVX1_LOC_54/Y INVX1_LOC_588/A 0.03fF
C21712 INVX1_LOC_47/Y INVX1_LOC_100/Y 0.50fF
C21713 NAND2X1_LOC_557/B INVX1_LOC_100/Y 1.04fF
C21714 NAND2X1_LOC_333/A INVX1_LOC_635/Y 0.04fF
C21715 INVX1_LOC_31/Y INVX1_LOC_75/Y 4.06fF
C21716 NAND2X1_LOC_432/Y NAND2X1_LOC_832/A 0.00fF
C21717 INVX1_LOC_50/Y INVX1_LOC_658/Y 0.04fF
C21718 NAND2X1_LOC_306/a_36_24# INVX1_LOC_74/Y 0.00fF
C21719 NAND2X1_LOC_165/Y NAND2X1_LOC_231/B 0.06fF
C21720 INVX1_LOC_47/Y INVX1_LOC_74/Y 0.37fF
C21721 INVX1_LOC_93/Y NAND2X1_LOC_619/a_36_24# 0.00fF
C21722 INVX1_LOC_47/Y INVX1_LOC_483/Y 0.02fF
C21723 NAND2X1_LOC_269/B INVX1_LOC_245/A 0.01fF
C21724 INVX1_LOC_93/Y NAND2X1_LOC_98/B 0.06fF
C21725 VDD INVX1_LOC_192/Y 0.21fF
C21726 INVX1_LOC_100/Y INVX1_LOC_119/Y 0.04fF
C21727 VDD INVX1_LOC_421/Y 0.23fF
C21728 INVX1_LOC_31/Y NAND2X1_LOC_271/A 0.07fF
C21729 INVX1_LOC_117/Y INVX1_LOC_92/A 0.29fF
C21730 INVX1_LOC_119/Y INVX1_LOC_74/Y 1.72fF
C21731 INVX1_LOC_269/Y NAND2X1_LOC_475/A 0.01fF
C21732 NAND2X1_LOC_66/Y INVX1_LOC_483/Y 0.02fF
C21733 INVX1_LOC_51/A INVX1_LOC_442/A 0.01fF
C21734 INVX1_LOC_445/Y INVX1_LOC_450/A 0.06fF
C21735 INVX1_LOC_438/Y NAND2X1_LOC_261/Y 0.03fF
C21736 INVX1_LOC_546/Y INVX1_LOC_557/A 0.12fF
C21737 NAND2X1_LOC_249/Y NAND2X1_LOC_107/Y 0.02fF
C21738 INVX1_LOC_17/Y INVX1_LOC_220/A 0.06fF
C21739 NAND2X1_LOC_58/a_36_24# NAND2X1_LOC_318/B 0.01fF
C21740 NAND2X1_LOC_475/A INVX1_LOC_320/A 0.02fF
C21741 INVX1_LOC_99/Y NAND2X1_LOC_591/B 0.04fF
C21742 INVX1_LOC_118/Y INVX1_LOC_596/A 0.03fF
C21743 INVX1_LOC_257/Y INVX1_LOC_197/A 0.07fF
C21744 INVX1_LOC_401/Y INPUT_0 0.01fF
C21745 INVX1_LOC_393/A INVX1_LOC_384/A 0.06fF
C21746 NAND2X1_LOC_704/a_36_24# NAND2X1_LOC_307/A 0.00fF
C21747 INVX1_LOC_299/Y GATE_366 0.26fF
C21748 INVX1_LOC_53/Y INVX1_LOC_373/A 0.05fF
C21749 NAND2X1_LOC_341/a_36_24# INVX1_LOC_275/A 0.02fF
C21750 INVX1_LOC_150/Y INVX1_LOC_501/Y 0.01fF
C21751 INVX1_LOC_584/A INVX1_LOC_632/A 0.05fF
C21752 NAND2X1_LOC_172/a_36_24# INVX1_LOC_638/A 0.01fF
C21753 INVX1_LOC_434/A INVX1_LOC_17/Y 0.56fF
C21754 INVX1_LOC_384/A INVX1_LOC_384/Y 0.05fF
C21755 NAND2X1_LOC_242/A INVX1_LOC_99/Y 0.02fF
C21756 VDD INVX1_LOC_159/A 0.00fF
C21757 INVX1_LOC_213/Y NAND2X1_LOC_249/Y 0.01fF
C21758 INVX1_LOC_21/Y INVX1_LOC_490/Y 0.12fF
C21759 INVX1_LOC_551/Y INVX1_LOC_76/Y 0.17fF
C21760 INVX1_LOC_435/A INVX1_LOC_206/Y 0.03fF
C21761 INVX1_LOC_270/A NAND2X1_LOC_318/A 0.09fF
C21762 INVX1_LOC_417/Y INVX1_LOC_400/Y 0.72fF
C21763 INVX1_LOC_133/Y NAND2X1_LOC_647/A 0.01fF
C21764 INVX1_LOC_51/A INVX1_LOC_116/Y 0.02fF
C21765 INVX1_LOC_595/Y NAND2X1_LOC_763/Y 0.02fF
C21766 VDD NAND2X1_LOC_615/B 0.50fF
C21767 NAND2X1_LOC_56/Y INVX1_LOC_586/A 0.07fF
C21768 INVX1_LOC_80/A INVX1_LOC_364/Y 0.01fF
C21769 NAND2X1_LOC_93/Y INVX1_LOC_50/Y 0.42fF
C21770 NAND2X1_LOC_690/a_36_24# INVX1_LOC_542/A 0.00fF
C21771 INVX1_LOC_446/Y NAND2X1_LOC_416/Y 0.05fF
C21772 INPUT_0 INVX1_LOC_510/A 0.07fF
C21773 NAND2X1_LOC_147/B NAND2X1_LOC_142/Y 0.18fF
C21774 INVX1_LOC_127/A INVX1_LOC_35/Y 0.17fF
C21775 VDD INVX1_LOC_127/Y 0.20fF
C21776 INVX1_LOC_468/Y INVX1_LOC_546/Y 0.01fF
C21777 INVX1_LOC_438/A INVX1_LOC_50/Y 0.08fF
C21778 INVX1_LOC_400/Y INVX1_LOC_59/Y 0.09fF
C21779 INVX1_LOC_59/A NAND2X1_LOC_53/a_36_24# 0.02fF
C21780 INVX1_LOC_492/A INVX1_LOC_395/A 0.11fF
C21781 INVX1_LOC_47/Y NAND2X1_LOC_591/B 0.03fF
C21782 INVX1_LOC_84/A INVX1_LOC_28/Y 0.02fF
C21783 INVX1_LOC_53/Y INVX1_LOC_235/Y 0.07fF
C21784 INVX1_LOC_224/Y INVX1_LOC_93/Y 0.03fF
C21785 INVX1_LOC_228/Y NAND2X1_LOC_615/B 0.03fF
C21786 NAND2X1_LOC_331/A INVX1_LOC_164/Y 0.15fF
C21787 NAND2X1_LOC_516/Y INVX1_LOC_510/A 0.01fF
C21788 VDD INVX1_LOC_66/A 1.26fF
C21789 INVX1_LOC_400/Y INVX1_LOC_48/Y 0.03fF
C21790 INVX1_LOC_492/Y INVX1_LOC_633/Y 0.27fF
C21791 NAND2X1_LOC_45/Y NAND2X1_LOC_181/A 0.03fF
C21792 INVX1_LOC_321/Y INVX1_LOC_482/A 0.00fF
C21793 INVX1_LOC_268/Y NAND2X1_LOC_755/B 0.00fF
C21794 INVX1_LOC_80/A INVX1_LOC_134/Y 0.43fF
C21795 INVX1_LOC_566/A INVX1_LOC_99/Y 0.35fF
C21796 NAND2X1_LOC_498/Y INVX1_LOC_350/Y 0.04fF
C21797 NAND2X1_LOC_174/B INVX1_LOC_288/A 0.14fF
C21798 INVX1_LOC_578/A INVX1_LOC_93/Y 0.14fF
C21799 INVX1_LOC_570/A INVX1_LOC_350/Y 0.01fF
C21800 NAND2X1_LOC_673/A INVX1_LOC_169/A 0.01fF
C21801 INVX1_LOC_602/A INVX1_LOC_602/Y 0.02fF
C21802 INVX1_LOC_288/A NAND2X1_LOC_591/Y 0.07fF
C21803 INVX1_LOC_198/Y INVX1_LOC_366/A 0.04fF
C21804 INVX1_LOC_51/A INVX1_LOC_255/A 0.05fF
C21805 INVX1_LOC_21/Y INVX1_LOC_97/Y 0.03fF
C21806 NAND2X1_LOC_122/a_36_24# INVX1_LOC_497/A 0.00fF
C21807 INVX1_LOC_542/A INVX1_LOC_463/Y 0.03fF
C21808 INVX1_LOC_167/A INVX1_LOC_76/Y 0.00fF
C21809 NAND2X1_LOC_122/Y NAND2X1_LOC_448/B 0.00fF
C21810 VDD INVX1_LOC_178/Y 0.30fF
C21811 INVX1_LOC_224/Y INVX1_LOC_390/A 0.01fF
C21812 INVX1_LOC_213/Y NAND2X1_LOC_833/a_36_24# 0.00fF
C21813 INVX1_LOC_428/A INVX1_LOC_69/Y 0.12fF
C21814 INVX1_LOC_514/Y NAND2X1_LOC_679/B 0.01fF
C21815 INVX1_LOC_25/Y INVX1_LOC_29/Y 0.04fF
C21816 INVX1_LOC_592/Y INVX1_LOC_45/Y 0.01fF
C21817 INVX1_LOC_510/Y INVX1_LOC_66/A 0.07fF
C21818 INVX1_LOC_53/Y INVX1_LOC_556/Y 0.14fF
C21819 INVX1_LOC_447/A INVX1_LOC_502/A 0.15fF
C21820 INVX1_LOC_11/Y INVX1_LOC_134/Y 0.27fF
C21821 NAND2X1_LOC_45/Y INVX1_LOC_79/A 0.01fF
C21822 NAND2X1_LOC_704/B NAND2X1_LOC_308/A 0.27fF
C21823 VDD NAND2X1_LOC_601/Y 0.04fF
C21824 INVX1_LOC_584/A NAND2X1_LOC_434/B 0.28fF
C21825 INPUT_0 INVX1_LOC_485/Y 0.01fF
C21826 INVX1_LOC_426/A INVX1_LOC_75/Y 0.09fF
C21827 NAND2X1_LOC_475/A INVX1_LOC_100/Y 0.10fF
C21828 INVX1_LOC_558/A INVX1_LOC_49/Y 0.00fF
C21829 INVX1_LOC_88/Y INVX1_LOC_6/Y 0.01fF
C21830 NAND2X1_LOC_416/Y INVX1_LOC_145/Y 0.06fF
C21831 INVX1_LOC_145/Y NAND2X1_LOC_285/B 0.03fF
C21832 NAND2X1_LOC_513/A INVX1_LOC_50/Y 0.04fF
C21833 INVX1_LOC_188/Y INVX1_LOC_345/A 0.07fF
C21834 INVX1_LOC_80/A NAND2X1_LOC_165/Y 0.01fF
C21835 INPUT_7 NAND2X1_LOC_429/a_36_24# 0.00fF
C21836 INVX1_LOC_566/A INVX1_LOC_47/Y 0.06fF
C21837 INVX1_LOC_117/Y INVX1_LOC_679/Y 0.07fF
C21838 INVX1_LOC_454/A INVX1_LOC_74/A 0.03fF
C21839 INVX1_LOC_145/Y NAND2X1_LOC_106/B 0.04fF
C21840 INVX1_LOC_17/Y INVX1_LOC_350/A 0.00fF
C21841 NAND2X1_LOC_177/a_36_24# INVX1_LOC_255/A 0.01fF
C21842 INVX1_LOC_65/Y INVX1_LOC_179/Y 0.01fF
C21843 VDD NAND2X1_LOC_621/B 0.01fF
C21844 NAND2X1_LOC_464/a_36_24# INVX1_LOC_116/Y 0.00fF
C21845 INVX1_LOC_602/A INVX1_LOC_292/Y 0.31fF
C21846 INVX1_LOC_437/A NAND2X1_LOC_556/a_36_24# 0.00fF
C21847 INVX1_LOC_11/Y NAND2X1_LOC_41/Y 0.02fF
C21848 NAND2X1_LOC_475/A INVX1_LOC_74/Y 0.10fF
C21849 NAND2X1_LOC_498/Y INVX1_LOC_79/A 0.10fF
C21850 INVX1_LOC_401/A INVX1_LOC_58/Y 0.03fF
C21851 INVX1_LOC_581/A NAND2X1_LOC_647/A 0.03fF
C21852 INVX1_LOC_570/A INVX1_LOC_79/A 0.05fF
C21853 NAND2X1_LOC_493/B INVX1_LOC_9/Y 0.01fF
C21854 VDD NAND2X1_LOC_646/B 0.07fF
C21855 INVX1_LOC_265/Y INVX1_LOC_74/Y 0.01fF
C21856 INVX1_LOC_335/Y INVX1_LOC_18/Y 0.09fF
C21857 INVX1_LOC_469/Y INVX1_LOC_99/Y 0.05fF
C21858 INVX1_LOC_80/A INVX1_LOC_65/A 0.01fF
C21859 INVX1_LOC_6/Y INVX1_LOC_600/A 0.06fF
C21860 INVX1_LOC_173/Y INVX1_LOC_145/Y 0.00fF
C21861 INVX1_LOC_287/A INVX1_LOC_154/A 0.01fF
C21862 INVX1_LOC_586/A INVX1_LOC_369/Y 0.10fF
C21863 INVX1_LOC_502/Y INVX1_LOC_100/Y 0.03fF
C21864 INVX1_LOC_439/Y NAND2X1_LOC_348/a_36_24# 0.08fF
C21865 INVX1_LOC_103/Y INVX1_LOC_159/A 0.00fF
C21866 INVX1_LOC_633/Y INVX1_LOC_168/Y 0.00fF
C21867 INVX1_LOC_117/Y INVX1_LOC_681/Y 0.03fF
C21868 INVX1_LOC_293/A NAND2X1_LOC_260/Y 0.02fF
C21869 INVX1_LOC_567/Y INVX1_LOC_58/Y 0.01fF
C21870 INVX1_LOC_20/Y NAND2X1_LOC_470/a_36_24# 0.00fF
C21871 INVX1_LOC_442/A INVX1_LOC_441/A 0.02fF
C21872 INVX1_LOC_117/Y INPUT_1 0.17fF
C21873 NAND2X1_LOC_707/A INVX1_LOC_62/Y 4.09fF
C21874 INVX1_LOC_45/Y INVX1_LOC_479/A 2.22fF
C21875 INVX1_LOC_49/Y NAND2X1_LOC_755/B 0.02fF
C21876 INVX1_LOC_421/A INVX1_LOC_48/Y 0.29fF
C21877 INVX1_LOC_51/Y INVX1_LOC_75/Y 0.03fF
C21878 NAND2X1_LOC_383/a_36_24# INVX1_LOC_31/Y 0.01fF
C21879 NAND2X1_LOC_493/B INVX1_LOC_62/Y 0.07fF
C21880 INVX1_LOC_525/Y INVX1_LOC_527/Y 0.11fF
C21881 INVX1_LOC_164/Y NAND2X1_LOC_186/a_36_24# 0.00fF
C21882 NAND2X1_LOC_433/Y INVX1_LOC_134/Y 0.07fF
C21883 NAND2X1_LOC_527/Y INVX1_LOC_93/Y 0.03fF
C21884 NAND2X1_LOC_274/B NAND2X1_LOC_601/a_36_24# 0.00fF
C21885 INVX1_LOC_625/A INVX1_LOC_44/Y 0.03fF
C21886 INVX1_LOC_198/Y INVX1_LOC_6/Y 0.61fF
C21887 INVX1_LOC_341/Y INPUT_4 0.07fF
C21888 NAND2X1_LOC_106/Y INVX1_LOC_608/A 0.02fF
C21889 INVX1_LOC_241/A INVX1_LOC_242/A 0.10fF
C21890 INVX1_LOC_103/Y INVX1_LOC_66/A 0.03fF
C21891 INVX1_LOC_531/Y INVX1_LOC_635/A 0.42fF
C21892 INVX1_LOC_62/Y INVX1_LOC_517/A 0.01fF
C21893 NAND2X1_LOC_336/B INVX1_LOC_62/Y 0.02fF
C21894 NAND2X1_LOC_542/A INVX1_LOC_670/A 0.12fF
C21895 INVX1_LOC_504/A NAND2X1_LOC_436/a_36_24# 0.01fF
C21896 INVX1_LOC_54/Y INVX1_LOC_63/Y 0.21fF
C21897 INVX1_LOC_76/Y INVX1_LOC_634/Y 0.07fF
C21898 INVX1_LOC_531/Y NAND2X1_LOC_237/Y 0.06fF
C21899 INVX1_LOC_484/A INVX1_LOC_6/Y 0.03fF
C21900 INVX1_LOC_183/A INVX1_LOC_172/A 0.03fF
C21901 INVX1_LOC_99/Y INVX1_LOC_79/A 0.26fF
C21902 INVX1_LOC_49/Y INVX1_LOC_46/Y 0.11fF
C21903 INVX1_LOC_51/Y NAND2X1_LOC_271/A 0.09fF
C21904 INVX1_LOC_257/A INVX1_LOC_253/Y 0.03fF
C21905 INVX1_LOC_32/Y INVX1_LOC_480/A 0.01fF
C21906 NAND2X1_LOC_106/Y INVX1_LOC_58/Y 0.03fF
C21907 INVX1_LOC_356/A INVX1_LOC_462/Y 0.20fF
C21908 NAND2X1_LOC_24/Y NAND2X1_LOC_617/a_36_24# 0.01fF
C21909 INVX1_LOC_208/Y INVX1_LOC_44/Y 0.06fF
C21910 INVX1_LOC_99/Y INVX1_LOC_460/A 0.01fF
C21911 INVX1_LOC_670/A INVX1_LOC_376/Y 1.07fF
C21912 NAND2X1_LOC_97/B INVX1_LOC_211/A 0.00fF
C21913 INVX1_LOC_607/Y NAND2X1_LOC_248/B 0.00fF
C21914 INVX1_LOC_496/A INVX1_LOC_493/Y 0.03fF
C21915 INVX1_LOC_25/Y INVX1_LOC_74/Y 0.12fF
C21916 INVX1_LOC_116/Y INVX1_LOC_441/A 0.02fF
C21917 INVX1_LOC_6/Y NAND2X1_LOC_780/a_36_24# 0.00fF
C21918 INVX1_LOC_297/Y INVX1_LOC_596/Y 0.02fF
C21919 NAND2X1_LOC_165/a_36_24# NAND2X1_LOC_231/B 0.01fF
C21920 NAND2X1_LOC_638/A INVX1_LOC_636/A 0.07fF
C21921 NAND2X1_LOC_263/a_36_24# INVX1_LOC_178/A 0.01fF
C21922 INVX1_LOC_47/Y INVX1_LOC_79/A 0.33fF
C21923 NAND2X1_LOC_334/B NAND2X1_LOC_291/a_36_24# 0.02fF
C21924 NAND2X1_LOC_123/B INVX1_LOC_58/Y 0.00fF
C21925 INVX1_LOC_89/Y INVX1_LOC_588/A 0.03fF
C21926 INVX1_LOC_105/Y INVX1_LOC_109/A 0.00fF
C21927 INVX1_LOC_251/Y INVX1_LOC_92/A 0.07fF
C21928 INVX1_LOC_255/A INVX1_LOC_441/A 0.10fF
C21929 VDD INVX1_LOC_438/Y 0.39fF
C21930 INVX1_LOC_433/Y INVX1_LOC_434/A 0.08fF
C21931 NAND2X1_LOC_274/B INVX1_LOC_114/A 0.00fF
C21932 INVX1_LOC_100/Y INVX1_LOC_663/A 0.01fF
C21933 INVX1_LOC_79/A INVX1_LOC_119/Y 0.26fF
C21934 INVX1_LOC_501/A INVX1_LOC_588/A 0.03fF
C21935 INVX1_LOC_79/A NAND2X1_LOC_66/Y 0.07fF
C21936 VDD INVX1_LOC_408/Y 0.22fF
C21937 INVX1_LOC_69/Y NAND2X1_LOC_832/A 0.02fF
C21938 NAND2X1_LOC_66/Y NAND2X1_LOC_631/B 0.01fF
C21939 INVX1_LOC_224/Y INVX1_LOC_395/A 0.07fF
C21940 INVX1_LOC_58/Y INVX1_LOC_270/Y 0.02fF
C21941 INVX1_LOC_584/A INVX1_LOC_561/Y 0.00fF
C21942 INVX1_LOC_133/Y INVX1_LOC_569/A 0.01fF
C21943 INPUT_0 NAND2X1_LOC_558/a_36_24# 0.01fF
C21944 NAND2X1_LOC_788/A INVX1_LOC_510/Y 0.03fF
C21945 INVX1_LOC_128/Y INVX1_LOC_666/Y 0.05fF
C21946 INVX1_LOC_76/Y INVX1_LOC_596/Y 0.00fF
C21947 NAND2X1_LOC_231/B INVX1_LOC_90/Y 0.03fF
C21948 INVX1_LOC_58/Y INVX1_LOC_92/A 0.15fF
C21949 INVX1_LOC_578/A INVX1_LOC_395/A 0.14fF
C21950 INVX1_LOC_557/A INVX1_LOC_395/A 0.36fF
C21951 INVX1_LOC_21/Y INVX1_LOC_615/A 0.00fF
C21952 INPUT_0 INVX1_LOC_321/A 0.03fF
C21953 NAND2X1_LOC_90/a_36_24# INVX1_LOC_92/A 0.01fF
C21954 INVX1_LOC_304/Y INVX1_LOC_109/Y 0.05fF
C21955 VDD INVX1_LOC_196/A -0.00fF
C21956 INVX1_LOC_158/A INVX1_LOC_270/A 0.03fF
C21957 NAND2X1_LOC_475/A INVX1_LOC_566/A 0.05fF
C21958 INVX1_LOC_206/Y INVX1_LOC_59/A 0.03fF
C21959 INVX1_LOC_211/Y INVX1_LOC_297/Y 0.03fF
C21960 INVX1_LOC_617/Y INPUT_0 0.07fF
C21961 INVX1_LOC_206/Y INVX1_LOC_367/A 0.07fF
C21962 INVX1_LOC_627/A INVX1_LOC_137/Y 0.01fF
C21963 INVX1_LOC_133/Y INVX1_LOC_137/Y 0.01fF
C21964 INVX1_LOC_86/A NAND2X1_LOC_85/a_36_24# 0.02fF
C21965 INVX1_LOC_287/A INVX1_LOC_203/Y 0.00fF
C21966 VDD INVX1_LOC_268/A 0.00fF
C21967 INVX1_LOC_402/A INVX1_LOC_238/A 0.06fF
C21968 INVX1_LOC_617/Y NAND2X1_LOC_516/Y 0.10fF
C21969 VDD INVX1_LOC_526/Y 0.26fF
C21970 INVX1_LOC_24/A NAND2X1_LOC_513/A 0.01fF
C21971 INVX1_LOC_21/Y INVX1_LOC_54/A 0.01fF
C21972 VDD INVX1_LOC_116/Y 0.21fF
C21973 INVX1_LOC_447/A INVX1_LOC_17/Y 0.00fF
C21974 INVX1_LOC_412/Y NAND2X1_LOC_123/A 0.23fF
C21975 INVX1_LOC_20/Y NAND2X1_LOC_352/a_36_24# 0.01fF
C21976 INVX1_LOC_446/A INVX1_LOC_54/Y 0.25fF
C21977 INVX1_LOC_372/Y INVX1_LOC_45/Y 0.03fF
C21978 INVX1_LOC_287/Y INVX1_LOC_76/Y 0.02fF
C21979 INVX1_LOC_206/Y INVX1_LOC_669/Y 0.00fF
C21980 VDD INVX1_LOC_219/Y 0.36fF
C21981 INVX1_LOC_270/A INVX1_LOC_76/Y 0.00fF
C21982 INVX1_LOC_577/A INVX1_LOC_99/Y 0.03fF
C21983 NAND2X1_LOC_217/a_36_24# NAND2X1_LOC_111/Y 0.00fF
C21984 VDD NAND2X1_LOC_432/Y -0.00fF
C21985 INVX1_LOC_448/Y INPUT_1 0.01fF
C21986 VDD INVX1_LOC_18/A 0.00fF
C21987 INVX1_LOC_206/Y INVX1_LOC_400/A 0.51fF
C21988 INVX1_LOC_568/Y INVX1_LOC_395/A 0.01fF
C21989 INVX1_LOC_78/A NAND2X1_LOC_513/Y 0.18fF
C21990 VDD INVX1_LOC_328/A -0.00fF
C21991 INVX1_LOC_12/Y INVX1_LOC_45/Y 0.07fF
C21992 NAND2X1_LOC_45/Y INVX1_LOC_48/Y 0.04fF
C21993 INVX1_LOC_367/A INVX1_LOC_242/A 0.46fF
C21994 INVX1_LOC_261/Y INVX1_LOC_638/A 1.36fF
C21995 NAND2X1_LOC_704/B INVX1_LOC_134/Y 0.07fF
C21996 INVX1_LOC_372/Y INVX1_LOC_348/A 0.01fF
C21997 INVX1_LOC_114/Y INVX1_LOC_632/A 0.02fF
C21998 VDD INPUT_4 0.56fF
C21999 INVX1_LOC_523/A INVX1_LOC_35/Y 0.09fF
C22000 INVX1_LOC_167/Y INVX1_LOC_633/Y 0.01fF
C22001 INVX1_LOC_258/Y INVX1_LOC_638/A 0.02fF
C22002 INVX1_LOC_393/Y INVX1_LOC_665/Y 0.02fF
C22003 INVX1_LOC_121/Y INVX1_LOC_670/A 0.03fF
C22004 NAND2X1_LOC_701/a_36_24# INVX1_LOC_361/Y 0.00fF
C22005 INVX1_LOC_206/Y INVX1_LOC_93/Y 0.73fF
C22006 INVX1_LOC_224/Y INVX1_LOC_31/Y 0.17fF
C22007 NAND2X1_LOC_332/B INVX1_LOC_124/Y 0.03fF
C22008 INVX1_LOC_65/Y INVX1_LOC_194/Y 0.10fF
C22009 INVX1_LOC_54/Y INVX1_LOC_374/A 0.03fF
C22010 NAND2X1_LOC_151/a_36_24# INVX1_LOC_53/Y 0.01fF
C22011 INVX1_LOC_578/A INVX1_LOC_31/Y 0.07fF
C22012 INVX1_LOC_202/Y NAND2X1_LOC_318/A 0.05fF
C22013 NAND2X1_LOC_534/Y INVX1_LOC_63/Y 0.02fF
C22014 INVX1_LOC_384/A INVX1_LOC_510/A 0.47fF
C22015 NAND2X1_LOC_431/a_36_24# INVX1_LOC_638/A 0.01fF
C22016 INVX1_LOC_32/A INVX1_LOC_49/Y 0.01fF
C22017 INVX1_LOC_211/Y INVX1_LOC_76/Y 0.02fF
C22018 INVX1_LOC_185/Y INVX1_LOC_138/Y 0.01fF
C22019 NAND2X1_LOC_763/a_36_24# INVX1_LOC_366/A 0.00fF
C22020 INVX1_LOC_442/A INVX1_LOC_103/Y 0.01fF
C22021 GATE_579 INVX1_LOC_439/Y 0.10fF
C22022 INVX1_LOC_51/A INVX1_LOC_69/Y 0.00fF
C22023 VDD INVX1_LOC_179/A 0.06fF
C22024 INVX1_LOC_206/Y INVX1_LOC_675/A 0.18fF
C22025 INVX1_LOC_370/Y INVX1_LOC_80/A 0.03fF
C22026 INVX1_LOC_84/A INVX1_LOC_176/A 0.01fF
C22027 NAND2X1_LOC_241/B INVX1_LOC_69/Y 0.01fF
C22028 VDD NAND2X1_LOC_719/A 0.00fF
C22029 INVX1_LOC_208/A INVX1_LOC_273/A 0.03fF
C22030 INVX1_LOC_602/A INVX1_LOC_53/A 0.02fF
C22031 INVX1_LOC_391/A INVX1_LOC_45/Y 0.00fF
C22032 NAND2X1_LOC_164/Y INVX1_LOC_44/Y 0.12fF
C22033 INVX1_LOC_395/A INVX1_LOC_120/Y 0.03fF
C22034 NAND2X1_LOC_543/B INVX1_LOC_100/Y 0.08fF
C22035 INVX1_LOC_367/Y INVX1_LOC_134/Y 0.07fF
C22036 INVX1_LOC_632/A INVX1_LOC_99/Y 0.07fF
C22037 INVX1_LOC_499/Y INVX1_LOC_463/Y 0.01fF
C22038 INVX1_LOC_21/Y INVX1_LOC_275/Y 0.21fF
C22039 INVX1_LOC_206/Y NAND2X1_LOC_334/B 0.00fF
C22040 NAND2X1_LOC_475/A NAND2X1_LOC_558/B 0.02fF
C22041 INVX1_LOC_76/Y INVX1_LOC_46/Y 2.11fF
C22042 NAND2X1_LOC_636/A INVX1_LOC_41/Y 0.01fF
C22043 NAND2X1_LOC_706/a_36_24# INVX1_LOC_367/A 0.00fF
C22044 INVX1_LOC_35/Y INVX1_LOC_519/A 0.06fF
C22045 INVX1_LOC_379/A NAND2X1_LOC_296/Y 0.05fF
C22046 NAND2X1_LOC_307/A NAND2X1_LOC_775/B 0.07fF
C22047 INVX1_LOC_417/Y INVX1_LOC_99/Y 0.01fF
C22048 INVX1_LOC_195/A INVX1_LOC_26/Y 0.01fF
C22049 INVX1_LOC_137/Y INVX1_LOC_633/Y 5.16fF
C22050 INVX1_LOC_581/A INVX1_LOC_137/Y 0.34fF
C22051 INVX1_LOC_624/Y INVX1_LOC_618/Y 0.96fF
C22052 NAND2X1_LOC_775/B INVX1_LOC_545/Y 0.00fF
C22053 INVX1_LOC_20/Y NAND2X1_LOC_364/a_36_24# 0.00fF
C22054 INVX1_LOC_602/A INVX1_LOC_50/Y 0.02fF
C22055 INVX1_LOC_9/Y INVX1_LOC_215/Y 0.01fF
C22056 INVX1_LOC_323/Y INVX1_LOC_35/Y 0.01fF
C22057 INVX1_LOC_170/A INVX1_LOC_45/Y 0.00fF
C22058 INVX1_LOC_398/Y INVX1_LOC_99/Y 0.01fF
C22059 INVX1_LOC_342/A INVX1_LOC_59/A 0.06fF
C22060 INVX1_LOC_93/Y INVX1_LOC_686/A 0.10fF
C22061 INVX1_LOC_11/Y NAND2X1_LOC_253/a_36_24# 0.00fF
C22062 INVX1_LOC_166/A NAND2X1_LOC_273/a_36_24# 0.00fF
C22063 INVX1_LOC_448/A INVX1_LOC_510/A 0.12fF
C22064 INVX1_LOC_65/Y INVX1_LOC_44/Y 0.09fF
C22065 NAND2X1_LOC_543/B INVX1_LOC_74/Y 0.08fF
C22066 INVX1_LOC_99/Y INVX1_LOC_59/Y 0.03fF
C22067 NAND2X1_LOC_636/B INVX1_LOC_50/Y 0.04fF
C22068 INVX1_LOC_20/Y NAND2X1_LOC_753/Y 0.12fF
C22069 INVX1_LOC_490/Y INVX1_LOC_26/Y 0.09fF
C22070 INVX1_LOC_579/A NAND2X1_LOC_448/B 0.00fF
C22071 INVX1_LOC_171/Y INVX1_LOC_63/Y 0.00fF
C22072 INVX1_LOC_268/Y INVX1_LOC_49/Y 0.01fF
C22073 NAND2X1_LOC_532/Y NAND2X1_LOC_512/a_36_24# 0.01fF
C22074 INVX1_LOC_84/A INVX1_LOC_410/A 0.01fF
C22075 INVX1_LOC_99/Y INVX1_LOC_48/Y 6.61fF
C22076 INVX1_LOC_549/A INVX1_LOC_41/Y 0.13fF
C22077 INVX1_LOC_257/Y INVX1_LOC_66/Y 0.03fF
C22078 INVX1_LOC_183/Y INVX1_LOC_366/A 0.11fF
C22079 INVX1_LOC_670/Y INVX1_LOC_199/A 0.01fF
C22080 INVX1_LOC_419/A NAND2X1_LOC_545/B 0.00fF
C22081 INVX1_LOC_84/A INVX1_LOC_170/Y 0.06fF
C22082 NAND2X1_LOC_250/Y INVX1_LOC_277/A 0.22fF
C22083 INVX1_LOC_675/A INVX1_LOC_686/A 2.39fF
C22084 INVX1_LOC_47/Y INVX1_LOC_632/A 0.07fF
C22085 INVX1_LOC_184/A INVX1_LOC_44/Y 0.01fF
C22086 INVX1_LOC_103/Y INVX1_LOC_116/Y -0.02fF
C22087 INVX1_LOC_468/Y INVX1_LOC_31/Y 0.03fF
C22088 INVX1_LOC_672/A INVX1_LOC_221/Y 0.01fF
C22089 INVX1_LOC_662/A NAND2X1_LOC_820/Y 0.06fF
C22090 INVX1_LOC_47/Y INVX1_LOC_509/Y 0.01fF
C22091 NAND2X1_LOC_111/Y NAND2X1_LOC_325/B 0.36fF
C22092 INVX1_LOC_560/A INVX1_LOC_666/Y 0.07fF
C22093 INVX1_LOC_188/Y INVX1_LOC_347/Y 0.03fF
C22094 INVX1_LOC_679/Y INVX1_LOC_58/Y 0.69fF
C22095 INVX1_LOC_312/Y NAND2X1_LOC_768/B 0.01fF
C22096 INVX1_LOC_361/Y INVX1_LOC_665/Y 0.00fF
C22097 INVX1_LOC_531/Y INVX1_LOC_666/A 0.19fF
C22098 INVX1_LOC_80/A INVX1_LOC_351/A 0.03fF
C22099 INVX1_LOC_117/Y INVX1_LOC_50/Y 0.27fF
C22100 NAND2X1_LOC_529/Y NAND2X1_LOC_531/Y 0.02fF
C22101 INVX1_LOC_69/Y NAND2X1_LOC_270/a_36_24# 0.01fF
C22102 INVX1_LOC_602/Y INVX1_LOC_58/Y 1.46fF
C22103 INVX1_LOC_604/Y INVX1_LOC_44/Y 0.11fF
C22104 INVX1_LOC_127/Y INVX1_LOC_105/A 0.01fF
C22105 INVX1_LOC_261/Y INVX1_LOC_685/Y 0.23fF
C22106 INVX1_LOC_123/A INVX1_LOC_48/Y 0.01fF
C22107 NAND2X1_LOC_708/A INVX1_LOC_6/Y 0.18fF
C22108 NAND2X1_LOC_491/Y INVX1_LOC_99/Y 0.04fF
C22109 NAND2X1_LOC_520/a_36_24# INVX1_LOC_69/Y 0.01fF
C22110 INVX1_LOC_685/A INVX1_LOC_674/Y 0.01fF
C22111 INVX1_LOC_230/A INVX1_LOC_411/Y 0.03fF
C22112 INVX1_LOC_97/Y INVX1_LOC_26/Y 0.00fF
C22113 INVX1_LOC_80/A INVX1_LOC_90/Y 0.09fF
C22114 NAND2X1_LOC_324/a_36_24# INVX1_LOC_376/A 0.00fF
C22115 INVX1_LOC_294/Y INVX1_LOC_369/Y 0.01fF
C22116 INVX1_LOC_47/Y INVX1_LOC_48/Y 2.19fF
C22117 NAND2X1_LOC_13/Y INVX1_LOC_75/Y 0.08fF
C22118 INVX1_LOC_76/Y INVX1_LOC_75/A 0.02fF
C22119 INVX1_LOC_500/Y INVX1_LOC_513/Y 0.05fF
C22120 INVX1_LOC_293/Y NAND2X1_LOC_528/Y 0.28fF
C22121 INVX1_LOC_448/A NAND2X1_LOC_477/a_36_24# 0.00fF
C22122 NAND2X1_LOC_557/B INVX1_LOC_48/Y 0.04fF
C22123 INVX1_LOC_502/A NAND2X1_LOC_658/a_36_24# 0.00fF
C22124 NAND2X1_LOC_106/Y NAND2X1_LOC_496/a_36_24# 0.00fF
C22125 INVX1_LOC_509/Y INVX1_LOC_119/Y 0.01fF
C22126 INVX1_LOC_585/Y INVX1_LOC_63/Y 0.01fF
C22127 INVX1_LOC_293/Y INVX1_LOC_479/A 0.07fF
C22128 INPUT_1 INVX1_LOC_58/Y 0.30fF
C22129 NAND2X1_LOC_601/a_36_24# INVX1_LOC_468/A 0.00fF
C22130 INVX1_LOC_117/Y INVX1_LOC_517/Y 0.04fF
C22131 INVX1_LOC_41/Y NAND2X1_LOC_237/Y 0.05fF
C22132 INVX1_LOC_507/Y INVX1_LOC_189/A 0.03fF
C22133 INVX1_LOC_99/Y INVX1_LOC_472/Y 0.01fF
C22134 INVX1_LOC_391/Y INVX1_LOC_26/Y 0.00fF
C22135 INVX1_LOC_89/Y INVX1_LOC_253/Y 0.00fF
C22136 NAND2X1_LOC_759/a_36_24# INVX1_LOC_26/Y 0.00fF
C22137 NAND2X1_LOC_638/A INVX1_LOC_74/Y 9.27fF
C22138 INVX1_LOC_437/A INVX1_LOC_430/Y 0.09fF
C22139 INVX1_LOC_21/Y INVX1_LOC_274/Y 0.03fF
C22140 INVX1_LOC_179/Y INVX1_LOC_86/Y 0.02fF
C22141 INVX1_LOC_11/Y INVX1_LOC_90/Y 0.19fF
C22142 INVX1_LOC_253/Y NAND2X1_LOC_319/a_36_24# 0.00fF
C22143 INVX1_LOC_89/Y INVX1_LOC_63/Y 1.20fF
C22144 INVX1_LOC_41/Y INVX1_LOC_230/A 0.00fF
C22145 INVX1_LOC_119/Y INVX1_LOC_48/Y 0.10fF
C22146 INVX1_LOC_145/Y NAND2X1_LOC_248/B 0.00fF
C22147 NAND2X1_LOC_66/Y INVX1_LOC_48/Y 0.11fF
C22148 INVX1_LOC_31/Y NAND2X1_LOC_291/a_36_24# 0.01fF
C22149 INVX1_LOC_242/Y INVX1_LOC_260/Y 0.01fF
C22150 INVX1_LOC_202/Y INVX1_LOC_92/Y 0.02fF
C22151 INVX1_LOC_675/A NAND2X1_LOC_334/A 0.07fF
C22152 INVX1_LOC_26/Y INVX1_LOC_18/Y 0.78fF
C22153 NAND2X1_LOC_243/a_36_24# INVX1_LOC_198/A 0.00fF
C22154 INVX1_LOC_501/A INVX1_LOC_63/Y 0.06fF
C22155 INVX1_LOC_507/A INVX1_LOC_507/Y 0.00fF
C22156 INVX1_LOC_74/Y INVX1_LOC_505/A 0.23fF
C22157 INVX1_LOC_46/Y INVX1_LOC_184/Y 0.04fF
C22158 INVX1_LOC_369/Y INVX1_LOC_6/Y 0.01fF
C22159 INVX1_LOC_183/Y NAND2X1_LOC_81/Y -0.06fF
C22160 INVX1_LOC_179/A NAND2X1_LOC_786/B 0.07fF
C22161 INVX1_LOC_15/Y INVX1_LOC_79/A 0.01fF
C22162 INVX1_LOC_395/A NAND2X1_LOC_86/Y 0.01fF
C22163 INVX1_LOC_253/Y NAND2X1_LOC_544/B 0.02fF
C22164 INVX1_LOC_513/A INVX1_LOC_462/Y 0.00fF
C22165 INVX1_LOC_100/Y NAND2X1_LOC_445/a_36_24# 0.00fF
C22166 INVX1_LOC_69/Y INVX1_LOC_441/A 0.00fF
C22167 NAND2X1_LOC_786/B NAND2X1_LOC_262/a_36_24# 0.02fF
C22168 INVX1_LOC_426/A INVX1_LOC_578/A 0.47fF
C22169 INVX1_LOC_257/Y INVX1_LOC_412/Y 0.01fF
C22170 INVX1_LOC_79/A NAND2X1_LOC_627/Y 0.08fF
C22171 INVX1_LOC_204/Y INVX1_LOC_620/Y 0.01fF
C22172 INVX1_LOC_74/Y INVX1_LOC_353/A 0.07fF
C22173 INPUT_0 INVX1_LOC_553/Y 0.00fF
C22174 INVX1_LOC_206/Y INVX1_LOC_395/A 0.35fF
C22175 INPUT_0 INVX1_LOC_410/Y 0.07fF
C22176 INVX1_LOC_395/A INVX1_LOC_648/Y 0.06fF
C22177 INVX1_LOC_412/Y INVX1_LOC_288/A 0.92fF
C22178 NAND2X1_LOC_164/Y INVX1_LOC_96/Y 0.55fF
C22179 VDD INVX1_LOC_146/A -0.00fF
C22180 INVX1_LOC_270/Y INVX1_LOC_245/A 1.47fF
C22181 NAND2X1_LOC_91/a_36_24# INVX1_LOC_92/A 0.00fF
C22182 INVX1_LOC_224/Y INVX1_LOC_51/Y 0.03fF
C22183 NAND2X1_LOC_516/Y INVX1_LOC_375/A 0.03fF
C22184 INVX1_LOC_209/Y INVX1_LOC_274/Y 0.98fF
C22185 INVX1_LOC_570/A NAND2X1_LOC_513/Y 0.07fF
C22186 INVX1_LOC_51/A INVX1_LOC_586/A 0.01fF
C22187 NAND2X1_LOC_65/Y INPUT_0 0.01fF
C22188 INVX1_LOC_245/A INVX1_LOC_92/A 0.00fF
C22189 INVX1_LOC_266/A INVX1_LOC_224/Y 0.10fF
C22190 INVX1_LOC_567/A INVX1_LOC_558/Y 0.05fF
C22191 INVX1_LOC_578/A INVX1_LOC_51/Y 0.26fF
C22192 INVX1_LOC_395/A INVX1_LOC_242/A 0.07fF
C22193 INVX1_LOC_206/Y INVX1_LOC_683/Y 0.01fF
C22194 INVX1_LOC_200/Y INVX1_LOC_126/Y 0.01fF
C22195 NAND2X1_LOC_370/A NAND2X1_LOC_315/a_36_24# 0.00fF
C22196 INVX1_LOC_266/A INVX1_LOC_578/A 0.10fF
C22197 NAND2X1_LOC_317/B NAND2X1_LOC_307/A 0.06fF
C22198 INVX1_LOC_395/A INVX1_LOC_686/A 0.24fF
C22199 INVX1_LOC_424/A INVX1_LOC_386/Y 0.03fF
C22200 INVX1_LOC_454/A INVX1_LOC_316/Y 0.03fF
C22201 INVX1_LOC_3/Y INVX1_LOC_25/Y 0.46fF
C22202 INVX1_LOC_252/Y NAND2X1_LOC_76/B 0.00fF
C22203 NAND2X1_LOC_318/A INVX1_LOC_76/Y 0.33fF
C22204 NAND2X1_LOC_475/A INVX1_LOC_59/Y 0.02fF
C22205 INVX1_LOC_617/Y INVX1_LOC_384/A -0.04fF
C22206 INVX1_LOC_448/Y INVX1_LOC_50/Y 0.01fF
C22207 INVX1_LOC_315/Y INVX1_LOC_635/A 0.02fF
C22208 VDD NAND2X1_LOC_148/B 0.02fF
C22209 NAND2X1_LOC_513/Y INVX1_LOC_99/Y 0.39fF
C22210 NAND2X1_LOC_475/A INVX1_LOC_48/Y 0.22fF
C22211 NAND2X1_LOC_457/A INVX1_LOC_159/Y 0.00fF
C22212 INVX1_LOC_438/A INVX1_LOC_117/Y 0.14fF
C22213 INVX1_LOC_20/Y NAND2X1_LOC_105/a_36_24# 0.00fF
C22214 INPUT_0 INVX1_LOC_61/A 0.34fF
C22215 INVX1_LOC_683/Y INVX1_LOC_686/A 0.01fF
C22216 NAND2X1_LOC_362/a_36_24# INVX1_LOC_230/A 0.00fF
C22217 INVX1_LOC_239/Y NAND2X1_LOC_342/A 0.23fF
C22218 INVX1_LOC_586/A NAND2X1_LOC_413/Y 0.15fF
C22219 INVX1_LOC_17/Y INVX1_LOC_173/A 0.06fF
C22220 INVX1_LOC_400/A INVX1_LOC_397/A 0.01fF
C22221 INVX1_LOC_468/Y INVX1_LOC_51/Y 0.03fF
C22222 INVX1_LOC_206/Y INVX1_LOC_31/Y 2.07fF
C22223 INVX1_LOC_76/Y INVX1_LOC_115/A 0.06fF
C22224 NAND2X1_LOC_88/B NAND2X1_LOC_87/a_36_24# 0.00fF
C22225 VDD INVX1_LOC_69/Y 2.25fF
C22226 INVX1_LOC_463/A INVX1_LOC_513/Y 0.09fF
C22227 INVX1_LOC_26/Y INVX1_LOC_615/A 0.08fF
C22228 INVX1_LOC_202/Y INVX1_LOC_98/A 0.00fF
C22229 INVX1_LOC_45/Y INVX1_LOC_159/A 0.01fF
C22230 INVX1_LOC_617/Y INVX1_LOC_448/A 0.02fF
C22231 INVX1_LOC_442/A INVX1_LOC_105/A 0.00fF
C22232 INVX1_LOC_21/A NAND2X1_LOC_5/a_36_24# 0.00fF
C22233 INVX1_LOC_202/Y INVX1_LOC_76/Y 0.52fF
C22234 NAND2X1_LOC_332/B INVX1_LOC_510/A 0.07fF
C22235 INVX1_LOC_20/Y NAND2X1_LOC_285/B 0.02fF
C22236 INVX1_LOC_561/Y INVX1_LOC_47/Y 0.02fF
C22237 NAND2X1_LOC_475/A NAND2X1_LOC_491/Y 0.01fF
C22238 NAND2X1_LOC_527/Y INVX1_LOC_51/Y 0.02fF
C22239 INVX1_LOC_20/Y NAND2X1_LOC_106/B 0.01fF
C22240 NAND2X1_LOC_387/Y INVX1_LOC_266/Y 0.07fF
C22241 INVX1_LOC_21/Y NAND2X1_LOC_237/Y 0.03fF
C22242 INVX1_LOC_435/A INVX1_LOC_295/A 0.03fF
C22243 VDD INVX1_LOC_247/Y 0.26fF
C22244 NAND2X1_LOC_543/B INVX1_LOC_79/A 0.16fF
C22245 INVX1_LOC_435/Y INVX1_LOC_234/Y 0.01fF
C22246 INVX1_LOC_608/Y NAND2X1_LOC_496/Y 0.00fF
C22247 INVX1_LOC_335/A NAND2X1_LOC_685/A 0.12fF
C22248 NAND2X1_LOC_322/Y INVX1_LOC_100/Y 0.14fF
C22249 INVX1_LOC_58/A INVX1_LOC_55/Y 0.03fF
C22250 INVX1_LOC_33/Y INVX1_LOC_6/Y 0.03fF
C22251 INVX1_LOC_80/A INVX1_LOC_98/Y 0.06fF
C22252 INVX1_LOC_17/Y NAND2X1_LOC_496/Y 0.02fF
C22253 INVX1_LOC_84/A INVX1_LOC_54/Y 0.15fF
C22254 INVX1_LOC_409/A INVX1_LOC_114/A 0.00fF
C22255 INVX1_LOC_294/A INVX1_LOC_297/A 0.01fF
C22256 INVX1_LOC_287/Y INVX1_LOC_32/Y 0.01fF
C22257 INVX1_LOC_270/A INVX1_LOC_32/Y 0.46fF
C22258 VDD INVX1_LOC_667/A -0.00fF
C22259 INVX1_LOC_522/Y INVX1_LOC_189/A 0.10fF
C22260 NAND2X1_LOC_498/B INVX1_LOC_49/Y 0.28fF
C22261 INVX1_LOC_510/Y INVX1_LOC_69/Y 0.07fF
C22262 INVX1_LOC_20/Y INVX1_LOC_173/Y 0.01fF
C22263 INVX1_LOC_17/Y NAND2X1_LOC_525/a_36_24# 0.00fF
C22264 INVX1_LOC_10/Y INVX1_LOC_83/Y 0.02fF
C22265 INVX1_LOC_658/A INVX1_LOC_50/Y 0.02fF
C22266 INVX1_LOC_117/Y INVX1_LOC_187/A 0.03fF
C22267 INVX1_LOC_374/A INVX1_LOC_501/A 0.03fF
C22268 INVX1_LOC_409/Y INVX1_LOC_74/Y 0.03fF
C22269 INVX1_LOC_402/A INVX1_LOC_556/Y 0.01fF
C22270 INVX1_LOC_546/Y INVX1_LOC_376/Y 0.00fF
C22271 INPUT_0 INVX1_LOC_273/Y 0.09fF
C22272 INVX1_LOC_12/Y NAND2X1_LOC_673/B 0.14fF
C22273 INVX1_LOC_156/Y INVX1_LOC_157/A 0.14fF
C22274 NAND2X1_LOC_271/B INVX1_LOC_502/A 0.00fF
C22275 INVX1_LOC_164/Y INVX1_LOC_134/Y 0.05fF
C22276 INVX1_LOC_12/A INVX1_LOC_46/Y 0.01fF
C22277 INVX1_LOC_361/Y INVX1_LOC_134/Y 0.07fF
C22278 NAND2X1_LOC_747/a_36_24# INVX1_LOC_581/A 0.00fF
C22279 INVX1_LOC_31/Y INVX1_LOC_686/A 0.15fF
C22280 INVX1_LOC_625/A INVX1_LOC_252/Y 0.00fF
C22281 INVX1_LOC_451/A INVX1_LOC_442/Y 0.00fF
C22282 INVX1_LOC_117/Y NAND2X1_LOC_513/A 0.07fF
C22283 INVX1_LOC_76/Y INVX1_LOC_49/Y 0.08fF
C22284 NAND2X1_LOC_122/Y NAND2X1_LOC_675/a_36_24# 0.00fF
C22285 INVX1_LOC_17/Y NAND2X1_LOC_775/B 0.07fF
C22286 INVX1_LOC_206/Y INVX1_LOC_473/Y 0.46fF
C22287 INVX1_LOC_531/Y NAND2X1_LOC_749/Y 0.03fF
C22288 INVX1_LOC_11/Y INVX1_LOC_98/Y 0.10fF
C22289 NAND2X1_LOC_836/B INVX1_LOC_334/Y 0.04fF
C22290 INVX1_LOC_205/Y INVX1_LOC_86/Y 0.02fF
C22291 INVX1_LOC_396/A INVX1_LOC_99/Y 0.01fF
C22292 INVX1_LOC_503/Y INVX1_LOC_510/A 0.03fF
C22293 INVX1_LOC_50/Y INVX1_LOC_281/Y 0.01fF
C22294 INVX1_LOC_367/A NAND2X1_LOC_542/A 0.09fF
C22295 INVX1_LOC_548/A NAND2X1_LOC_706/a_36_24# 0.00fF
C22296 INVX1_LOC_105/A INVX1_LOC_116/Y 0.01fF
C22297 INVX1_LOC_435/Y INVX1_LOC_665/A 0.03fF
C22298 NAND2X1_LOC_467/A INVX1_LOC_168/Y 0.10fF
C22299 NAND2X1_LOC_43/Y INVX1_LOC_48/Y 0.13fF
C22300 INVX1_LOC_50/Y INVX1_LOC_178/A 0.01fF
C22301 INVX1_LOC_7/Y INVX1_LOC_46/Y 0.84fF
C22302 INVX1_LOC_444/Y INVX1_LOC_444/A 0.00fF
C22303 INVX1_LOC_1/A INVX1_LOC_25/A 0.31fF
C22304 INVX1_LOC_68/Y INVX1_LOC_100/Y 0.06fF
C22305 INVX1_LOC_153/A INVX1_LOC_59/Y 0.00fF
C22306 INVX1_LOC_80/A INVX1_LOC_338/Y 0.02fF
C22307 INVX1_LOC_386/Y INVX1_LOC_387/Y 0.35fF
C22308 INVX1_LOC_194/Y INVX1_LOC_86/Y 0.11fF
C22309 INVX1_LOC_410/Y INVX1_LOC_211/A 0.02fF
C22310 INVX1_LOC_566/A INVX1_LOC_353/A 0.02fF
C22311 INVX1_LOC_166/A INVX1_LOC_137/Y 0.00fF
C22312 INVX1_LOC_53/Y INVX1_LOC_183/A 0.03fF
C22313 INVX1_LOC_69/Y INVX1_LOC_116/A 0.01fF
C22314 INVX1_LOC_98/A INVX1_LOC_92/Y 0.00fF
C22315 NAND2X1_LOC_165/Y NAND2X1_LOC_333/B 0.02fF
C22316 INVX1_LOC_236/A INVX1_LOC_476/A 0.01fF
C22317 INVX1_LOC_40/Y INVX1_LOC_93/A 0.08fF
C22318 NAND2X1_LOC_755/B NAND2X1_LOC_838/a_36_24# 0.00fF
C22319 INVX1_LOC_295/Y INVX1_LOC_230/Y 0.96fF
C22320 INVX1_LOC_68/Y INVX1_LOC_74/Y 0.03fF
C22321 INVX1_LOC_514/A INVX1_LOC_463/Y 0.00fF
C22322 INVX1_LOC_607/Y INVX1_LOC_646/Y 0.06fF
C22323 INVX1_LOC_586/A INVX1_LOC_441/A 0.00fF
C22324 NAND2X1_LOC_97/B INVX1_LOC_242/Y 0.05fF
C22325 NAND2X1_LOC_105/a_36_24# INVX1_LOC_655/A 0.00fF
C22326 INVX1_LOC_76/Y INVX1_LOC_92/Y 0.02fF
C22327 INVX1_LOC_318/Y INVX1_LOC_319/A 0.01fF
C22328 INVX1_LOC_32/Y INVX1_LOC_46/Y 0.09fF
C22329 INVX1_LOC_153/A NAND2X1_LOC_168/a_36_24# 0.02fF
C22330 NAND2X1_LOC_837/B INVX1_LOC_659/A 0.24fF
C22331 INVX1_LOC_417/A INVX1_LOC_242/Y 0.03fF
C22332 INVX1_LOC_11/Y INVX1_LOC_338/Y 1.42fF
C22333 NAND2X1_LOC_65/Y INVX1_LOC_64/Y 0.02fF
C22334 INVX1_LOC_649/Y INVX1_LOC_669/A 0.01fF
C22335 INVX1_LOC_6/Y NAND2X1_LOC_659/a_36_24# 0.00fF
C22336 NAND2X1_LOC_184/Y NAND2X1_LOC_523/a_36_24# 0.00fF
C22337 INVX1_LOC_63/Y INVX1_LOC_194/Y 0.03fF
C22338 INVX1_LOC_103/Y INVX1_LOC_69/Y 2.45fF
C22339 INVX1_LOC_84/A INVX1_LOC_388/A 0.01fF
C22340 INVX1_LOC_100/Y INVX1_LOC_600/A 0.35fF
C22341 INVX1_LOC_93/Y NAND2X1_LOC_542/A 0.03fF
C22342 INVX1_LOC_54/Y INVX1_LOC_496/A 0.03fF
C22343 NAND2X1_LOC_128/A NAND2X1_LOC_128/B 0.09fF
C22344 INVX1_LOC_58/Y INVX1_LOC_50/Y 3.94fF
C22345 INVX1_LOC_69/Y INVX1_LOC_68/A 0.02fF
C22346 NAND2X1_LOC_285/B INVX1_LOC_655/A 0.04fF
C22347 NAND2X1_LOC_286/A INVX1_LOC_46/Y 0.05fF
C22348 NAND2X1_LOC_325/B INVX1_LOC_41/Y 0.13fF
C22349 INVX1_LOC_44/Y INVX1_LOC_86/Y 0.01fF
C22350 INVX1_LOC_74/Y NAND2X1_LOC_302/A 0.02fF
C22351 INVX1_LOC_242/Y INVX1_LOC_440/Y 0.02fF
C22352 NAND2X1_LOC_106/B INVX1_LOC_655/A 0.06fF
C22353 NAND2X1_LOC_274/B INVX1_LOC_303/Y 0.02fF
C22354 INVX1_LOC_519/A INVX1_LOC_364/A 0.00fF
C22355 INVX1_LOC_11/Y NAND2X1_LOC_41/a_36_24# 0.00fF
C22356 INVX1_LOC_352/Y INVX1_LOC_114/A 0.03fF
C22357 INVX1_LOC_313/Y INVX1_LOC_90/Y 0.03fF
C22358 INVX1_LOC_26/Y NAND2X1_LOC_84/B 0.17fF
C22359 INPUT_1 INVX1_LOC_245/A 0.06fF
C22360 INVX1_LOC_53/Y INVX1_LOC_109/A 0.00fF
C22361 NAND2X1_LOC_400/B INVX1_LOC_183/A 0.01fF
C22362 INVX1_LOC_534/Y INVX1_LOC_463/Y 0.04fF
C22363 INVX1_LOC_549/Y INVX1_LOC_62/Y 0.01fF
C22364 INVX1_LOC_89/A INVX1_LOC_66/A 0.29fF
C22365 INVX1_LOC_504/A INVX1_LOC_505/Y 0.07fF
C22366 INVX1_LOC_345/A INVX1_LOC_114/A 0.00fF
C22367 INVX1_LOC_47/Y NAND2X1_LOC_615/Y 0.06fF
C22368 INVX1_LOC_48/Y NAND2X1_LOC_627/Y 0.02fF
C22369 INVX1_LOC_517/Y INVX1_LOC_58/Y 0.01fF
C22370 INVX1_LOC_63/Y INVX1_LOC_44/Y 0.14fF
C22371 INVX1_LOC_69/Y NAND2X1_LOC_786/B 0.01fF
C22372 NAND2X1_LOC_355/A INVX1_LOC_632/Y 0.01fF
C22373 INVX1_LOC_657/A INVX1_LOC_659/A 0.01fF
C22374 NAND2X1_LOC_274/B INVX1_LOC_9/Y 0.03fF
C22375 NAND2X1_LOC_683/a_36_24# INVX1_LOC_245/A 0.01fF
C22376 INVX1_LOC_368/A INVX1_LOC_245/A 0.00fF
C22377 INVX1_LOC_137/Y INVX1_LOC_613/A 0.01fF
C22378 VDD INVX1_LOC_217/A 0.00fF
C22379 INVX1_LOC_484/A INVX1_LOC_483/Y 0.03fF
C22380 INVX1_LOC_69/Y INVX1_LOC_635/Y 0.04fF
C22381 INVX1_LOC_63/Y INVX1_LOC_347/A 0.07fF
C22382 VDD NAND2X1_LOC_537/B 0.04fF
C22383 INVX1_LOC_6/Y INVX1_LOC_443/A 0.09fF
C22384 INVX1_LOC_76/Y INVX1_LOC_297/Y 0.26fF
C22385 INVX1_LOC_496/A NAND2X1_LOC_609/a_36_24# 0.01fF
C22386 NAND2X1_LOC_274/B INVX1_LOC_62/Y 0.03fF
C22387 INVX1_LOC_366/A INVX1_LOC_180/Y 0.04fF
C22388 NAND2X1_LOC_274/B NAND2X1_LOC_844/A 0.03fF
C22389 VDD INVX1_LOC_586/A 4.69fF
C22390 INVX1_LOC_395/A INVX1_LOC_390/Y 0.01fF
C22391 INVX1_LOC_473/Y NAND2X1_LOC_609/B 0.02fF
C22392 VDD INVX1_LOC_516/Y 0.21fF
C22393 INVX1_LOC_169/A INVX1_LOC_388/Y 0.02fF
C22394 INVX1_LOC_62/Y INVX1_LOC_148/Y 0.02fF
C22395 INVX1_LOC_206/Y INVX1_LOC_51/Y 0.40fF
C22396 NAND2X1_LOC_750/Y INVX1_LOC_366/A 0.01fF
C22397 INVX1_LOC_90/Y INVX1_LOC_91/Y 0.07fF
C22398 INVX1_LOC_380/A INVX1_LOC_17/Y 0.03fF
C22399 VDD INVX1_LOC_246/Y 0.21fF
C22400 INVX1_LOC_395/A INVX1_LOC_94/A 0.01fF
C22401 INVX1_LOC_224/Y NAND2X1_LOC_13/Y 0.02fF
C22402 INVX1_LOC_266/A INVX1_LOC_206/Y 0.08fF
C22403 INVX1_LOC_618/A INVX1_LOC_468/Y 0.01fF
C22404 INVX1_LOC_384/A INVX1_LOC_410/Y 0.25fF
C22405 VDD INVX1_LOC_312/Y 0.65fF
C22406 INVX1_LOC_567/A NAND2X1_LOC_413/Y 0.00fF
C22407 INVX1_LOC_490/Y INVX1_LOC_235/Y 0.02fF
C22408 INVX1_LOC_510/Y INVX1_LOC_586/A 0.10fF
C22409 NAND2X1_LOC_498/B INVX1_LOC_76/Y 0.03fF
C22410 INVX1_LOC_424/A INVX1_LOC_7/Y 0.03fF
C22411 VDD INVX1_LOC_289/A -0.00fF
C22412 INVX1_LOC_98/A INVX1_LOC_76/Y 0.00fF
C22413 INVX1_LOC_51/Y INVX1_LOC_242/A 0.07fF
C22414 INVX1_LOC_133/Y INVX1_LOC_650/Y 0.01fF
C22415 VDD INVX1_LOC_241/Y 0.23fF
C22416 NAND2X1_LOC_710/A NAND2X1_LOC_498/Y 0.02fF
C22417 NAND2X1_LOC_539/a_36_24# INVX1_LOC_686/A 0.00fF
C22418 VDD NAND2X1_LOC_529/Y -0.00fF
C22419 VDD NAND2X1_LOC_378/Y 0.05fF
C22420 INVX1_LOC_95/Y NAND2X1_LOC_387/Y 0.01fF
C22421 INVX1_LOC_68/Y INVX1_LOC_566/A 0.24fF
C22422 INVX1_LOC_435/Y INVX1_LOC_80/A 0.10fF
C22423 INVX1_LOC_448/A INVX1_LOC_410/Y 0.01fF
C22424 NAND2X1_LOC_543/B INVX1_LOC_48/Y 0.01fF
C22425 INVX1_LOC_413/Y INVX1_LOC_53/Y 0.01fF
C22426 INVX1_LOC_617/Y NAND2X1_LOC_332/B 0.07fF
C22427 INVX1_LOC_317/Y NAND2X1_LOC_307/A 0.02fF
C22428 INVX1_LOC_51/Y INVX1_LOC_686/A 0.16fF
C22429 NAND2X1_LOC_332/B INVX1_LOC_119/A 0.01fF
C22430 NAND2X1_LOC_498/Y INVX1_LOC_383/Y 0.03fF
C22431 INVX1_LOC_406/Y INVX1_LOC_384/A 0.02fF
C22432 NAND2X1_LOC_170/a_36_24# NAND2X1_LOC_267/A 0.01fF
C22433 INVX1_LOC_409/Y INVX1_LOC_469/Y 0.01fF
C22434 INVX1_LOC_195/A INVX1_LOC_81/Y 0.01fF
C22435 INVX1_LOC_570/Y INVX1_LOC_575/Y 0.00fF
C22436 INVX1_LOC_418/A INVX1_LOC_130/Y 0.00fF
C22437 INVX1_LOC_266/A INVX1_LOC_686/A 0.10fF
C22438 NAND2X1_LOC_522/a_36_24# INVX1_LOC_384/A 0.01fF
C22439 NAND2X1_LOC_69/B INVX1_LOC_47/Y 0.01fF
C22440 VDD NAND2X1_LOC_835/A -0.00fF
C22441 INVX1_LOC_6/Y INVX1_LOC_180/Y 0.01fF
C22442 INVX1_LOC_58/Y INVX1_LOC_275/A 0.96fF
C22443 NAND2X1_LOC_122/Y NAND2X1_LOC_448/A 0.02fF
C22444 INVX1_LOC_206/Y INVX1_LOC_254/A 0.02fF
C22445 INVX1_LOC_395/A INVX1_LOC_432/A 0.01fF
C22446 NAND2X1_LOC_475/A INVX1_LOC_559/Y 0.36fF
C22447 INVX1_LOC_51/Y INVX1_LOC_14/A 0.01fF
C22448 INVX1_LOC_442/Y INVX1_LOC_364/Y 0.03fF
C22449 INVX1_LOC_20/Y NAND2X1_LOC_97/B 0.01fF
C22450 INVX1_LOC_586/A INVX1_LOC_116/A 0.00fF
C22451 INVX1_LOC_435/Y INVX1_LOC_11/Y 0.67fF
C22452 INVX1_LOC_45/Y INVX1_LOC_116/Y 0.00fF
C22453 INVX1_LOC_544/A INVX1_LOC_45/Y 0.04fF
C22454 VDD INVX1_LOC_157/Y 0.26fF
C22455 INVX1_LOC_44/A INVX1_LOC_366/A 0.03fF
C22456 INVX1_LOC_560/Y INVX1_LOC_154/A 0.01fF
C22457 INVX1_LOC_596/A INVX1_LOC_80/A 0.03fF
C22458 NAND2X1_LOC_677/Y NAND2X1_LOC_677/a_36_24# 0.02fF
C22459 INVX1_LOC_377/Y INVX1_LOC_383/Y 0.15fF
C22460 NAND2X1_LOC_208/a_36_24# INVX1_LOC_44/A 0.00fF
C22461 NAND2X1_LOC_58/a_36_24# INVX1_LOC_63/Y 0.00fF
C22462 NAND2X1_LOC_750/Y INVX1_LOC_6/Y 0.04fF
C22463 INVX1_LOC_17/Y NAND2X1_LOC_613/Y 0.02fF
C22464 NAND2X1_LOC_704/B INVX1_LOC_98/Y 0.05fF
C22465 INVX1_LOC_45/Y NAND2X1_LOC_432/Y 0.02fF
C22466 INVX1_LOC_420/Y INVX1_LOC_6/Y 0.01fF
C22467 INVX1_LOC_17/Y INVX1_LOC_169/A 0.06fF
C22468 NAND2X1_LOC_317/B NAND2X1_LOC_307/B 0.00fF
C22469 INVX1_LOC_406/Y INVX1_LOC_145/Y 0.04fF
C22470 INVX1_LOC_594/Y INVX1_LOC_675/A 0.22fF
C22471 INVX1_LOC_197/A NAND2X1_LOC_298/a_36_24# 0.00fF
C22472 INVX1_LOC_606/Y INVX1_LOC_6/Y 0.01fF
C22473 INVX1_LOC_174/Y INVX1_LOC_54/Y 0.01fF
C22474 INVX1_LOC_224/Y INVX1_LOC_361/A 0.02fF
C22475 INVX1_LOC_20/Y INVX1_LOC_510/A 0.07fF
C22476 INVX1_LOC_617/Y INVX1_LOC_503/Y 0.03fF
C22477 INVX1_LOC_99/Y NAND2X1_LOC_541/B 0.17fF
C22478 NAND2X1_LOC_638/A INVX1_LOC_632/A 0.02fF
C22479 INVX1_LOC_530/Y INVX1_LOC_32/Y 0.01fF
C22480 VDD INVX1_LOC_225/Y 0.21fF
C22481 INVX1_LOC_442/Y INVX1_LOC_134/Y 0.80fF
C22482 INVX1_LOC_80/A INVX1_LOC_504/A 0.08fF
C22483 NAND2X1_LOC_548/B INVX1_LOC_444/Y 0.07fF
C22484 INVX1_LOC_17/Y INVX1_LOC_633/Y 0.02fF
C22485 NAND2X1_LOC_97/B INVX1_LOC_300/A 0.01fF
C22486 INVX1_LOC_11/Y INVX1_LOC_596/A 0.09fF
C22487 INVX1_LOC_492/A NAND2X1_LOC_152/B 0.00fF
C22488 INVX1_LOC_552/Y INVX1_LOC_44/Y 0.07fF
C22489 NAND2X1_LOC_318/A INVX1_LOC_32/Y 0.02fF
C22490 INVX1_LOC_99/Y INVX1_LOC_155/Y 0.03fF
C22491 INVX1_LOC_47/Y INVX1_LOC_340/Y 0.03fF
C22492 INVX1_LOC_395/A INVX1_LOC_376/Y 0.10fF
C22493 INVX1_LOC_602/A INVX1_LOC_117/Y 1.72fF
C22494 INVX1_LOC_99/Y NAND2X1_LOC_93/a_36_24# 0.01fF
C22495 INVX1_LOC_312/Y INVX1_LOC_103/Y 0.03fF
C22496 NAND2X1_LOC_382/a_36_24# INVX1_LOC_295/Y -0.00fF
C22497 INVX1_LOC_452/A NAND2X1_LOC_569/a_36_24# 0.01fF
C22498 NAND2X1_LOC_636/B INVX1_LOC_117/Y 0.04fF
C22499 INVX1_LOC_84/A INVX1_LOC_89/Y 0.03fF
C22500 INVX1_LOC_166/A NAND2X1_LOC_307/A 0.03fF
C22501 INVX1_LOC_45/Y INVX1_LOC_179/A 0.03fF
C22502 INVX1_LOC_53/A INVX1_LOC_1/Y 0.01fF
C22503 INVX1_LOC_555/A INVX1_LOC_492/Y 0.01fF
C22504 NAND2X1_LOC_710/A INVX1_LOC_47/Y 0.02fF
C22505 NAND2X1_LOC_307/B INVX1_LOC_337/Y 0.10fF
C22506 INVX1_LOC_89/Y NAND2X1_LOC_410/a_36_24# -0.00fF
C22507 INVX1_LOC_545/A NAND2X1_LOC_775/B 0.03fF
C22508 INVX1_LOC_41/Y NAND2X1_LOC_749/Y 0.10fF
C22509 INVX1_LOC_63/A INVX1_LOC_204/Y 0.30fF
C22510 INVX1_LOC_674/A INVX1_LOC_145/Y 0.07fF
C22511 INPUT_0 NAND2X1_LOC_528/Y 0.01fF
C22512 NAND2X1_LOC_457/A NAND2X1_LOC_372/Y 0.03fF
C22513 INVX1_LOC_20/A INVX1_LOC_44/Y 0.02fF
C22514 INVX1_LOC_68/Y INVX1_LOC_77/A 0.01fF
C22515 INVX1_LOC_130/Y INVX1_LOC_46/Y 0.01fF
C22516 NAND2X1_LOC_13/Y NAND2X1_LOC_493/a_36_24# 0.01fF
C22517 INPUT_0 INVX1_LOC_479/A 0.10fF
C22518 NAND2X1_LOC_525/Y INVX1_LOC_41/Y 0.15fF
C22519 NAND2X1_LOC_413/Y INVX1_LOC_6/Y 0.00fF
C22520 INVX1_LOC_202/Y INVX1_LOC_32/Y 0.22fF
C22521 NAND2X1_LOC_513/A INVX1_LOC_58/Y 0.05fF
C22522 INVX1_LOC_677/Y INVX1_LOC_632/Y 0.02fF
C22523 INVX1_LOC_617/Y INVX1_LOC_242/Y 0.02fF
C22524 NAND2X1_LOC_338/a_36_24# INVX1_LOC_272/A 0.02fF
C22525 NAND2X1_LOC_516/Y INVX1_LOC_479/A 0.03fF
C22526 NAND2X1_LOC_131/a_36_24# INVX1_LOC_47/Y 0.00fF
C22527 INVX1_LOC_40/Y INVX1_LOC_342/A 0.01fF
C22528 INVX1_LOC_49/Y INVX1_LOC_7/Y 0.44fF
C22529 INVX1_LOC_99/A INVX1_LOC_411/Y 0.00fF
C22530 NAND2X1_LOC_710/A INVX1_LOC_119/Y 0.03fF
C22531 INVX1_LOC_586/A INVX1_LOC_635/Y 0.05fF
C22532 INVX1_LOC_360/Y INVX1_LOC_69/Y 0.07fF
C22533 INVX1_LOC_536/A NAND2X1_LOC_639/a_36_24# 0.00fF
C22534 INVX1_LOC_134/Y INVX1_LOC_471/Y 0.01fF
C22535 INVX1_LOC_635/A INVX1_LOC_26/Y 0.02fF
C22536 INVX1_LOC_557/Y INVX1_LOC_558/Y 0.11fF
C22537 NAND2X1_LOC_538/B INVX1_LOC_62/Y 0.01fF
C22538 INVX1_LOC_63/Y INVX1_LOC_365/A 0.01fF
C22539 NAND2X1_LOC_56/Y INVX1_LOC_100/Y 0.01fF
C22540 INVX1_LOC_20/Y NAND2X1_LOC_248/B 0.03fF
C22541 NAND2X1_LOC_260/Y INVX1_LOC_664/A 0.48fF
C22542 INVX1_LOC_26/Y NAND2X1_LOC_237/Y 0.18fF
C22543 INVX1_LOC_105/A INVX1_LOC_69/Y 0.01fF
C22544 INVX1_LOC_119/Y INVX1_LOC_383/Y 0.00fF
C22545 NAND2X1_LOC_403/A INVX1_LOC_328/Y 0.02fF
C22546 INVX1_LOC_403/Y INVX1_LOC_199/Y 0.11fF
C22547 INVX1_LOC_54/Y NAND2X1_LOC_376/B 0.05fF
C22548 NAND2X1_LOC_387/Y INVX1_LOC_199/Y 0.28fF
C22549 INVX1_LOC_59/Y INVX1_LOC_353/A 0.03fF
C22550 INVX1_LOC_145/Y INVX1_LOC_273/Y 0.60fF
C22551 INVX1_LOC_159/Y INVX1_LOC_9/Y 0.03fF
C22552 INVX1_LOC_555/A NAND2X1_LOC_647/A 0.02fF
C22553 INVX1_LOC_277/Y INVX1_LOC_221/Y 0.01fF
C22554 INVX1_LOC_93/Y INVX1_LOC_139/Y 0.02fF
C22555 INVX1_LOC_32/Y INVX1_LOC_49/Y 0.17fF
C22556 INVX1_LOC_50/Y NAND2X1_LOC_440/A 0.00fF
C22557 NAND2X1_LOC_445/a_36_24# INVX1_LOC_48/Y 0.01fF
C22558 INVX1_LOC_239/A NAND2X1_LOC_342/A 0.12fF
C22559 INVX1_LOC_381/A NAND2X1_LOC_415/a_36_24# 0.00fF
C22560 NAND2X1_LOC_388/A INVX1_LOC_58/Y 0.03fF
C22561 INVX1_LOC_353/A INVX1_LOC_48/Y 0.10fF
C22562 INVX1_LOC_50/Y INVX1_LOC_245/A 0.07fF
C22563 INVX1_LOC_31/Y INVX1_LOC_376/Y 0.07fF
C22564 INVX1_LOC_555/A INVX1_LOC_168/Y 0.02fF
C22565 NAND2X1_LOC_299/Y INVX1_LOC_634/Y 0.49fF
C22566 INVX1_LOC_137/Y INVX1_LOC_41/Y 0.03fF
C22567 NAND2X1_LOC_333/B INVX1_LOC_90/Y 0.08fF
C22568 INVX1_LOC_288/Y NAND2X1_LOC_451/B 0.03fF
C22569 INVX1_LOC_431/Y INVX1_LOC_245/A 0.02fF
C22570 INVX1_LOC_212/Y INVX1_LOC_9/Y 0.03fF
C22571 INVX1_LOC_525/Y NAND2X1_LOC_447/a_36_24# 0.01fF
C22572 NAND2X1_LOC_845/B INVX1_LOC_199/Y 0.09fF
C22573 INVX1_LOC_62/Y NAND2X1_LOC_412/a_36_24# 0.00fF
C22574 INVX1_LOC_63/Y NAND2X1_LOC_616/a_36_24# 0.00fF
C22575 NAND2X1_LOC_274/B INVX1_LOC_624/Y 0.00fF
C22576 INVX1_LOC_254/Y INVX1_LOC_211/A 0.02fF
C22577 INVX1_LOC_406/A INVX1_LOC_41/Y 0.00fF
C22578 NAND2X1_LOC_835/A INVX1_LOC_635/Y 0.01fF
C22579 INVX1_LOC_6/Y NAND2X1_LOC_488/Y 0.01fF
C22580 INVX1_LOC_479/A INVX1_LOC_498/A 0.04fF
C22581 INVX1_LOC_347/Y INVX1_LOC_114/A 0.11fF
C22582 VDD INVX1_LOC_151/Y 0.21fF
C22583 INVX1_LOC_301/A INVX1_LOC_412/Y 0.05fF
C22584 NAND2X1_LOC_294/Y INVX1_LOC_443/A 0.05fF
C22585 NAND2X1_LOC_88/Y INVX1_LOC_97/A 0.27fF
C22586 INVX1_LOC_434/A INVX1_LOC_445/A 0.05fF
C22587 VDD INVX1_LOC_140/Y 0.31fF
C22588 INVX1_LOC_655/A NAND2X1_LOC_248/B 0.07fF
C22589 INVX1_LOC_395/A INVX1_LOC_121/Y 0.03fF
C22590 INVX1_LOC_206/Y INVX1_LOC_355/A 0.12fF
C22591 INVX1_LOC_395/A INVX1_LOC_253/A 0.01fF
C22592 INVX1_LOC_301/A INVX1_LOC_119/A 0.02fF
C22593 VDD INVX1_LOC_272/Y 0.32fF
C22594 VDD NAND2X1_LOC_791/B 0.02fF
C22595 INVX1_LOC_410/Y NAND2X1_LOC_332/B 0.04fF
C22596 NAND2X1_LOC_13/Y INVX1_LOC_206/Y 0.00fF
C22597 NAND2X1_LOC_505/Y INVX1_LOC_397/A 0.04fF
C22598 VDD INVX1_LOC_486/Y 0.62fF
C22599 INVX1_LOC_20/Y INVX1_LOC_412/Y 0.09fF
C22600 VDD INVX1_LOC_294/Y 0.25fF
C22601 INVX1_LOC_479/A INVX1_LOC_211/A 0.00fF
C22602 INVX1_LOC_80/A NAND2X1_LOC_76/B 0.21fF
C22603 INVX1_LOC_479/A INVX1_LOC_464/Y 0.03fF
C22604 INVX1_LOC_447/A INVX1_LOC_519/A 0.01fF
C22605 INVX1_LOC_424/A NAND2X1_LOC_559/a_36_24# 0.00fF
C22606 VDD INVX1_LOC_597/A -0.00fF
C22607 INVX1_LOC_523/A INVX1_LOC_522/Y 0.05fF
C22608 INVX1_LOC_295/A INVX1_LOC_395/A 0.01fF
C22609 VDD INVX1_LOC_252/A 0.00fF
C22610 NAND2X1_LOC_271/B INVX1_LOC_232/Y 0.00fF
C22611 NAND2X1_LOC_475/A INVX1_LOC_155/Y 0.02fF
C22612 INVX1_LOC_132/Y INVX1_LOC_133/A 0.16fF
C22613 INVX1_LOC_556/A INVX1_LOC_53/Y 0.24fF
C22614 INVX1_LOC_412/A INVX1_LOC_134/Y 0.01fF
C22615 INPUT_0 INVX1_LOC_12/Y 1.68fF
C22616 INVX1_LOC_20/Y INVX1_LOC_321/A 0.36fF
C22617 NAND2X1_LOC_781/B INVX1_LOC_48/Y 0.14fF
C22618 INVX1_LOC_412/Y NAND2X1_LOC_605/a_36_24# 0.00fF
C22619 INVX1_LOC_21/Y NAND2X1_LOC_749/Y 0.12fF
C22620 INVX1_LOC_206/Y NAND2X1_LOC_72/a_36_24# 0.00fF
C22621 INVX1_LOC_11/Y NAND2X1_LOC_76/B 0.03fF
C22622 INVX1_LOC_85/Y INVX1_LOC_184/A 0.01fF
C22623 INVX1_LOC_445/Y INVX1_LOC_385/Y 8.19fF
C22624 INVX1_LOC_33/Y INVX1_LOC_29/Y 0.34fF
C22625 INVX1_LOC_20/Y INVX1_LOC_617/Y 0.07fF
C22626 NAND2X1_LOC_331/A INVX1_LOC_549/Y 0.01fF
C22627 INVX1_LOC_410/Y INVX1_LOC_503/Y 0.01fF
C22628 INVX1_LOC_560/A INVX1_LOC_230/A 0.02fF
C22629 INVX1_LOC_435/Y INVX1_LOC_367/Y 0.05fF
C22630 INVX1_LOC_435/Y INVX1_LOC_672/Y 0.07fF
C22631 INVX1_LOC_317/Y INVX1_LOC_17/Y 0.03fF
C22632 VDD INVX1_LOC_6/Y 1.37fF
C22633 INVX1_LOC_300/A INVX1_LOC_321/A 0.06fF
C22634 INVX1_LOC_463/A NAND2X1_LOC_334/A 0.07fF
C22635 INVX1_LOC_510/Y INVX1_LOC_252/A 0.03fF
C22636 INVX1_LOC_68/Y INVX1_LOC_59/Y 0.03fF
C22637 INVX1_LOC_452/Y INVX1_LOC_452/A 0.02fF
C22638 INVX1_LOC_670/Y INVX1_LOC_126/A 0.01fF
C22639 INVX1_LOC_76/Y INVX1_LOC_7/Y 0.00fF
C22640 NAND2X1_LOC_331/A INVX1_LOC_463/Y 0.59fF
C22641 INVX1_LOC_335/A INVX1_LOC_542/A 0.03fF
C22642 INVX1_LOC_68/Y INVX1_LOC_48/Y 0.07fF
C22643 INVX1_LOC_511/Y INVX1_LOC_511/A 0.09fF
C22644 INVX1_LOC_395/A INVX1_LOC_477/Y 0.06fF
C22645 INVX1_LOC_233/Y INVX1_LOC_48/Y 0.01fF
C22646 INVX1_LOC_206/Y NAND2X1_LOC_668/Y 0.04fF
C22647 INVX1_LOC_568/Y NAND2X1_LOC_152/B 0.01fF
C22648 INVX1_LOC_238/Y NAND2X1_LOC_847/A 0.01fF
C22649 NAND2X1_LOC_512/a_36_24# INVX1_LOC_99/Y 0.00fF
C22650 INVX1_LOC_53/Y NAND2X1_LOC_411/Y 0.02fF
C22651 INVX1_LOC_206/Y INVX1_LOC_361/A 0.01fF
C22652 INVX1_LOC_579/A NAND2X1_LOC_448/A 0.01fF
C22653 INVX1_LOC_98/A INVX1_LOC_32/Y 0.96fF
C22654 INPUT_0 INVX1_LOC_170/A 0.00fF
C22655 INVX1_LOC_366/A NAND2X1_LOC_243/A 0.13fF
C22656 INVX1_LOC_625/A INVX1_LOC_80/A 0.02fF
C22657 VDD NAND2X1_LOC_81/Y -0.00fF
C22658 INVX1_LOC_38/A INVX1_LOC_87/A 0.01fF
C22659 INVX1_LOC_84/A INVX1_LOC_194/Y 0.00fF
C22660 INVX1_LOC_523/A INVX1_LOC_508/A 0.30fF
C22661 INVX1_LOC_76/Y INVX1_LOC_32/Y 0.62fF
C22662 NAND2X1_LOC_613/Y INVX1_LOC_230/Y -0.04fF
C22663 NAND2X1_LOC_457/A INVX1_LOC_328/Y 0.00fF
C22664 INVX1_LOC_289/Y INVX1_LOC_58/Y 0.01fF
C22665 INVX1_LOC_398/Y INVX1_LOC_600/A 0.03fF
C22666 INVX1_LOC_375/Y INVX1_LOC_510/A 0.04fF
C22667 INVX1_LOC_442/Y INVX1_LOC_370/Y 0.02fF
C22668 INVX1_LOC_45/Y INVX1_LOC_69/Y 1.05fF
C22669 INVX1_LOC_51/Y NAND2X1_LOC_542/A 0.08fF
C22670 INVX1_LOC_292/A INVX1_LOC_26/Y 0.15fF
C22671 INVX1_LOC_410/Y INVX1_LOC_242/Y 0.03fF
C22672 INVX1_LOC_358/Y INVX1_LOC_137/Y 0.03fF
C22673 INVX1_LOC_224/Y NAND2X1_LOC_301/B 0.03fF
C22674 NAND2X1_LOC_140/B INVX1_LOC_510/A 0.05fF
C22675 NAND2X1_LOC_545/B INVX1_LOC_361/Y 0.03fF
C22676 INVX1_LOC_403/Y INVX1_LOC_53/Y 0.01fF
C22677 INVX1_LOC_21/Y INVX1_LOC_137/Y 0.02fF
C22678 NAND2X1_LOC_320/Y INVX1_LOC_504/Y 0.01fF
C22679 INVX1_LOC_602/Y INVX1_LOC_678/A 0.08fF
C22680 INVX1_LOC_375/A INVX1_LOC_242/Y 0.00fF
C22681 INPUT_0 INVX1_LOC_488/A 0.03fF
C22682 INVX1_LOC_435/A INVX1_LOC_379/A 0.07fF
C22683 INVX1_LOC_600/A INVX1_LOC_48/Y 0.53fF
C22684 INVX1_LOC_435/A INVX1_LOC_35/Y 0.07fF
C22685 INVX1_LOC_51/Y INVX1_LOC_376/Y 0.07fF
C22686 INVX1_LOC_376/Y NAND2X1_LOC_794/a_36_24# 0.00fF
C22687 INVX1_LOC_578/A NAND2X1_LOC_301/B 0.07fF
C22688 NAND2X1_LOC_714/a_36_24# NAND2X1_LOC_274/B 0.00fF
C22689 INVX1_LOC_45/Y INVX1_LOC_247/Y 0.05fF
C22690 INVX1_LOC_588/Y INVX1_LOC_17/Y 0.03fF
C22691 INVX1_LOC_614/A INVX1_LOC_6/Y 0.03fF
C22692 NAND2X1_LOC_403/A INVX1_LOC_172/A 0.00fF
C22693 INVX1_LOC_602/A INVX1_LOC_58/Y 0.03fF
C22694 NAND2X1_LOC_331/A INVX1_LOC_148/Y 0.00fF
C22695 INVX1_LOC_84/A INVX1_LOC_44/Y 3.09fF
C22696 INVX1_LOC_366/A NAND2X1_LOC_786/B 0.02fF
C22697 NAND2X1_LOC_333/B INVX1_LOC_98/Y 0.32fF
C22698 INVX1_LOC_361/Y INVX1_LOC_98/Y 0.02fF
C22699 NAND2X1_LOC_12/a_36_24# INVX1_LOC_26/Y 0.00fF
C22700 INVX1_LOC_591/Y INVX1_LOC_44/Y 0.06fF
C22701 INVX1_LOC_133/A INVX1_LOC_655/A 0.04fF
C22702 NAND2X1_LOC_636/B INVX1_LOC_58/Y 0.04fF
C22703 INVX1_LOC_435/Y NAND2X1_LOC_843/B 0.10fF
C22704 INVX1_LOC_413/A INVX1_LOC_54/Y 0.01fF
C22705 NAND2X1_LOC_174/a_36_24# INVX1_LOC_32/Y 0.01fF
C22706 INVX1_LOC_416/Y INVX1_LOC_75/Y 0.05fF
C22707 NAND2X1_LOC_331/Y INVX1_LOC_69/Y 0.03fF
C22708 NAND2X1_LOC_636/B NAND2X1_LOC_636/a_36_24# 0.00fF
C22709 INVX1_LOC_632/A NAND2X1_LOC_637/a_36_24# 0.00fF
C22710 NAND2X1_LOC_27/Y INVX1_LOC_50/Y 0.01fF
C22711 NAND2X1_LOC_106/Y NAND2X1_LOC_106/B 0.03fF
C22712 INVX1_LOC_187/A INVX1_LOC_245/A 0.01fF
C22713 INVX1_LOC_555/A INVX1_LOC_137/Y 0.16fF
C22714 INVX1_LOC_53/Y INVX1_LOC_491/A 0.46fF
C22715 INVX1_LOC_117/Y INVX1_LOC_608/A 0.05fF
C22716 INVX1_LOC_587/A INVX1_LOC_635/Y 0.00fF
C22717 INVX1_LOC_377/A INVX1_LOC_9/Y 0.01fF
C22718 INVX1_LOC_369/A NAND2X1_LOC_92/a_36_24# 0.00fF
C22719 INVX1_LOC_484/A INVX1_LOC_48/Y 0.01fF
C22720 INVX1_LOC_63/Y INVX1_LOC_252/Y 0.06fF
C22721 INVX1_LOC_193/A INVX1_LOC_89/Y 0.02fF
C22722 INVX1_LOC_437/A NAND2X1_LOC_344/B 0.05fF
C22723 INVX1_LOC_93/Y NAND2X1_LOC_619/Y 0.02fF
C22724 INVX1_LOC_17/Y NAND2X1_LOC_709/a_36_24# 0.00fF
C22725 NAND2X1_LOC_294/Y NAND2X1_LOC_479/a_36_24# 0.01fF
C22726 INVX1_LOC_557/Y NAND2X1_LOC_413/Y 0.01fF
C22727 NAND2X1_LOC_595/Y INVX1_LOC_9/Y 0.06fF
C22728 INVX1_LOC_419/Y INVX1_LOC_411/Y 0.04fF
C22729 INVX1_LOC_6/Y NAND2X1_LOC_243/A 0.01fF
C22730 INVX1_LOC_197/A NAND2X1_LOC_123/B 0.09fF
C22731 INVX1_LOC_201/Y INVX1_LOC_399/A 0.44fF
C22732 INVX1_LOC_641/Y INVX1_LOC_340/A 0.04fF
C22733 NAND2X1_LOC_307/A INVX1_LOC_41/Y 0.04fF
C22734 INVX1_LOC_166/A NAND2X1_LOC_307/B 0.00fF
C22735 INVX1_LOC_545/Y INVX1_LOC_41/Y 0.00fF
C22736 INVX1_LOC_117/Y INVX1_LOC_58/Y 0.65fF
C22737 INVX1_LOC_49/Y INVX1_LOC_110/A 0.01fF
C22738 NAND2X1_LOC_532/Y INVX1_LOC_89/Y 0.03fF
C22739 INVX1_LOC_31/Y NAND2X1_LOC_498/a_36_24# 0.00fF
C22740 INVX1_LOC_468/Y NAND2X1_LOC_301/B 0.04fF
C22741 INVX1_LOC_93/Y NAND2X1_LOC_618/a_36_24# 0.00fF
C22742 INVX1_LOC_663/Y INVX1_LOC_664/A 0.05fF
C22743 INVX1_LOC_11/Y INVX1_LOC_519/Y 0.01fF
C22744 INVX1_LOC_7/Y INVX1_LOC_184/Y 0.01fF
C22745 INVX1_LOC_69/Y NAND2X1_LOC_837/A 0.22fF
C22746 INVX1_LOC_261/Y INVX1_LOC_497/A 0.01fF
C22747 INVX1_LOC_17/Y INVX1_LOC_531/Y 0.03fF
C22748 INVX1_LOC_602/Y INVX1_LOC_657/Y 0.08fF
C22749 NAND2X1_LOC_173/Y INVX1_LOC_636/A 0.01fF
C22750 INVX1_LOC_662/A NAND2X1_LOC_819/a_36_24# 0.00fF
C22751 INVX1_LOC_12/Y INVX1_LOC_211/A 0.07fF
C22752 NAND2X1_LOC_528/Y INVX1_LOC_145/Y 0.02fF
C22753 INVX1_LOC_479/A INVX1_LOC_145/Y 0.16fF
C22754 INVX1_LOC_62/Y INVX1_LOC_352/Y 0.00fF
C22755 INVX1_LOC_559/Y INVX1_LOC_353/A 0.10fF
C22756 NAND2X1_LOC_545/A NAND2X1_LOC_444/A 0.08fF
C22757 INVX1_LOC_93/Y INVX1_LOC_652/A 0.00fF
C22758 INVX1_LOC_35/Y INVX1_LOC_241/A 0.01fF
C22759 INVX1_LOC_303/Y NAND2X1_LOC_372/Y 0.19fF
C22760 INVX1_LOC_6/Y NAND2X1_LOC_786/B 0.00fF
C22761 NAND2X1_LOC_597/Y INVX1_LOC_50/Y 0.06fF
C22762 INVX1_LOC_245/Y NAND2X1_LOC_294/Y 0.17fF
C22763 INVX1_LOC_17/Y NAND2X1_LOC_626/a_36_24# 0.00fF
C22764 INVX1_LOC_607/Y INVX1_LOC_212/A 0.06fF
C22765 INPUT_1 INVX1_LOC_652/Y 0.02fF
C22766 INVX1_LOC_89/Y NAND2X1_LOC_138/a_36_24# 0.00fF
C22767 INVX1_LOC_359/Y INVX1_LOC_74/Y 0.01fF
C22768 NAND2X1_LOC_518/a_36_24# INVX1_LOC_502/A 0.01fF
C22769 INVX1_LOC_75/Y INVX1_LOC_46/Y 0.19fF
C22770 INVX1_LOC_6/Y INVX1_LOC_635/Y 0.03fF
C22771 INVX1_LOC_87/A INVX1_LOC_39/Y 0.02fF
C22772 INVX1_LOC_482/Y INVX1_LOC_90/Y 0.39fF
C22773 NAND2X1_LOC_503/B INVX1_LOC_97/A 0.14fF
C22774 NAND2X1_LOC_7/Y INVX1_LOC_410/Y 0.11fF
C22775 INVX1_LOC_376/A INVX1_LOC_41/Y 0.07fF
C22776 INVX1_LOC_141/Y INVX1_LOC_479/A 0.02fF
C22777 INVX1_LOC_301/A INVX1_LOC_410/Y 0.07fF
C22778 INVX1_LOC_637/A INVX1_LOC_636/Y 0.14fF
C22779 INVX1_LOC_369/Y INVX1_LOC_79/A 0.07fF
C22780 INVX1_LOC_46/Y NAND2X1_LOC_271/A 0.07fF
C22781 NAND2X1_LOC_372/Y INVX1_LOC_9/Y 0.11fF
C22782 INVX1_LOC_183/A INVX1_LOC_327/A 0.01fF
C22783 INVX1_LOC_502/A INVX1_LOC_41/Y 0.08fF
C22784 INVX1_LOC_549/A INVX1_LOC_373/A 0.09fF
C22785 INVX1_LOC_675/A INVX1_LOC_462/Y 0.02fF
C22786 INVX1_LOC_395/A NAND2X1_LOC_750/a_36_24# 0.00fF
C22787 INVX1_LOC_62/Y INVX1_LOC_280/A 0.03fF
C22788 NAND2X1_LOC_537/B INVX1_LOC_45/Y 0.03fF
C22789 INVX1_LOC_79/A INVX1_LOC_348/Y 0.11fF
C22790 INVX1_LOC_97/A INVX1_LOC_273/A 0.20fF
C22791 INVX1_LOC_100/Y INVX1_LOC_443/A 0.03fF
C22792 INPUT_6 INVX1_LOC_595/A 0.00fF
C22793 INVX1_LOC_75/Y INVX1_LOC_75/A 0.05fF
C22794 INVX1_LOC_224/Y INVX1_LOC_551/Y 0.10fF
C22795 NAND2X1_LOC_506/B NAND2X1_LOC_419/a_36_24# 0.02fF
C22796 INVX1_LOC_20/Y INVX1_LOC_553/Y 0.00fF
C22797 VDD NAND2X1_LOC_517/Y 0.00fF
C22798 INVX1_LOC_20/Y INVX1_LOC_410/Y 0.06fF
C22799 NAND2X1_LOC_526/Y INVX1_LOC_362/Y 0.01fF
C22800 INVX1_LOC_586/A NAND2X1_LOC_506/B 0.02fF
C22801 NAND2X1_LOC_230/a_36_24# INVX1_LOC_91/A 0.00fF
C22802 INVX1_LOC_45/Y INVX1_LOC_586/A 5.62fF
C22803 INVX1_LOC_578/A INVX1_LOC_551/Y 0.10fF
C22804 NAND2X1_LOC_45/Y INVX1_LOC_90/A -0.01fF
C22805 NAND2X1_LOC_152/Y INVX1_LOC_570/A 0.00fF
C22806 NAND2X1_LOC_89/a_36_24# INVX1_LOC_98/A 0.00fF
C22807 NAND2X1_LOC_685/B INVX1_LOC_512/A 0.01fF
C22808 NAND2X1_LOC_164/Y INVX1_LOC_80/A 4.05fF
C22809 INVX1_LOC_558/A NAND2X1_LOC_515/a_36_24# 0.02fF
C22810 NAND2X1_LOC_331/A INVX1_LOC_537/Y 0.05fF
C22811 INPUT_3 INVX1_LOC_586/A 0.03fF
C22812 INVX1_LOC_288/A INVX1_LOC_372/Y 0.00fF
C22813 INVX1_LOC_312/Y INVX1_LOC_45/Y 4.88fF
C22814 INVX1_LOC_300/A INVX1_LOC_410/Y 0.03fF
C22815 VDD INVX1_LOC_415/Y 0.06fF
C22816 VDD NAND2X1_LOC_32/Y 0.03fF
C22817 INVX1_LOC_356/A NAND2X1_LOC_450/a_36_24# 0.02fF
C22818 INVX1_LOC_372/A INVX1_LOC_638/A 0.03fF
C22819 INVX1_LOC_395/A INVX1_LOC_251/A 0.03fF
C22820 NAND2X1_LOC_638/A INVX1_LOC_340/Y 0.03fF
C22821 INVX1_LOC_51/Y NAND2X1_LOC_603/Y 0.02fF
C22822 INVX1_LOC_619/A INVX1_LOC_366/A 0.11fF
C22823 INVX1_LOC_401/Y INVX1_LOC_401/A 0.01fF
C22824 VDD NAND2X1_LOC_294/Y 0.31fF
C22825 INPUT_0 NAND2X1_LOC_615/B 0.03fF
C22826 INVX1_LOC_11/Y NAND2X1_LOC_713/a_36_24# 0.01fF
C22827 INVX1_LOC_618/A INVX1_LOC_376/Y 0.04fF
C22828 INVX1_LOC_617/Y INVX1_LOC_375/Y 0.01fF
C22829 INVX1_LOC_84/A NAND2X1_LOC_391/A 0.00fF
C22830 INVX1_LOC_142/A INVX1_LOC_186/A 0.04fF
C22831 INVX1_LOC_601/A NAND2X1_LOC_232/a_36_24# 0.00fF
C22832 INPUT_0 INVX1_LOC_127/Y 0.01fF
C22833 INVX1_LOC_139/A INVX1_LOC_32/Y 0.00fF
C22834 INVX1_LOC_576/A INVX1_LOC_576/Y 0.01fF
C22835 INVX1_LOC_84/A INVX1_LOC_27/Y 0.01fF
C22836 INPUT_0 INVX1_LOC_66/A 0.10fF
C22837 INVX1_LOC_393/A INPUT_1 0.01fF
C22838 INVX1_LOC_206/Y NAND2X1_LOC_449/B 0.01fF
C22839 INVX1_LOC_255/Y INVX1_LOC_355/Y 0.00fF
C22840 INVX1_LOC_438/Y NAND2X1_LOC_344/B 2.53fF
C22841 INVX1_LOC_12/A INVX1_LOC_7/Y 0.03fF
C22842 INVX1_LOC_519/A NAND2X1_LOC_658/a_36_24# 0.02fF
C22843 NAND2X1_LOC_102/a_36_24# INVX1_LOC_686/A 0.00fF
C22844 VDD INVX1_LOC_206/A -0.00fF
C22845 INVX1_LOC_85/Y INVX1_LOC_86/Y 0.15fF
C22846 INPUT_3 NAND2X1_LOC_529/Y 0.16fF
C22847 NAND2X1_LOC_370/A INVX1_LOC_317/A 0.26fF
C22848 INVX1_LOC_35/Y INVX1_LOC_59/A 0.03fF
C22849 INVX1_LOC_20/Y INVX1_LOC_662/Y 0.03fF
C22850 VDD INVX1_LOC_557/Y 0.36fF
C22851 NAND2X1_LOC_299/Y INVX1_LOC_115/A 0.05fF
C22852 INVX1_LOC_524/Y INVX1_LOC_35/Y 0.02fF
C22853 NAND2X1_LOC_13/Y INVX1_LOC_432/A 0.00fF
C22854 NAND2X1_LOC_516/Y INVX1_LOC_66/A 0.03fF
C22855 INVX1_LOC_602/A INVX1_LOC_1/Y 0.02fF
C22856 GATE_741 INVX1_LOC_535/Y 0.04fF
C22857 INVX1_LOC_68/Y INVX1_LOC_559/Y 0.14fF
C22858 INVX1_LOC_367/A INVX1_LOC_35/Y 0.07fF
C22859 INVX1_LOC_554/Y NAND2X1_LOC_846/B 0.09fF
C22860 INVX1_LOC_80/A INVX1_LOC_370/A 0.01fF
C22861 INVX1_LOC_12/Y INVX1_LOC_145/Y 0.14fF
C22862 NAND2X1_LOC_331/Y INVX1_LOC_289/A 0.00fF
C22863 INVX1_LOC_586/A NAND2X1_LOC_837/A 0.42fF
C22864 INVX1_LOC_381/A INVX1_LOC_382/A 0.08fF
C22865 INVX1_LOC_80/A INVX1_LOC_479/Y 0.02fF
C22866 INVX1_LOC_449/A INVX1_LOC_303/Y 0.01fF
C22867 INVX1_LOC_576/A INVX1_LOC_674/A 0.05fF
C22868 INVX1_LOC_137/Y INVX1_LOC_474/Y 0.05fF
C22869 INVX1_LOC_679/Y NAND2X1_LOC_106/B 0.16fF
C22870 INVX1_LOC_176/A INVX1_LOC_99/Y 0.08fF
C22871 INVX1_LOC_686/A INVX1_LOC_359/A 0.01fF
C22872 INVX1_LOC_524/Y INVX1_LOC_620/A 0.20fF
C22873 NAND2X1_LOC_307/A NAND2X1_LOC_267/A 0.05fF
C22874 INVX1_LOC_542/A INVX1_LOC_499/A 0.45fF
C22875 INVX1_LOC_599/Y INVX1_LOC_623/Y 0.92fF
C22876 INVX1_LOC_250/Y INVX1_LOC_559/Y 0.28fF
C22877 NAND2X1_LOC_525/Y INVX1_LOC_26/Y 0.35fF
C22878 NAND2X1_LOC_756/Y INVX1_LOC_69/Y 0.00fF
C22879 INVX1_LOC_20/Y INVX1_LOC_646/Y 0.05fF
C22880 INVX1_LOC_551/A NAND2X1_LOC_318/A 0.01fF
C22881 INVX1_LOC_400/A INVX1_LOC_35/Y 0.04fF
C22882 INVX1_LOC_293/Y INVX1_LOC_69/Y 0.05fF
C22883 INVX1_LOC_510/Y INVX1_LOC_557/Y 0.01fF
C22884 NAND2X1_LOC_735/a_36_24# INVX1_LOC_502/A 0.01fF
C22885 INVX1_LOC_300/A INVX1_LOC_674/A 0.88fF
C22886 NAND2X1_LOC_399/B INVX1_LOC_32/Y 0.11fF
C22887 INVX1_LOC_285/A INVX1_LOC_204/Y 0.00fF
C22888 NAND2X1_LOC_198/a_36_24# INVX1_LOC_174/A 0.01fF
C22889 INVX1_LOC_25/Y INVX1_LOC_315/A 0.02fF
C22890 INVX1_LOC_32/Y INVX1_LOC_7/Y 0.07fF
C22891 NAND2X1_LOC_516/Y NAND2X1_LOC_601/Y 0.06fF
C22892 INVX1_LOC_619/A INVX1_LOC_6/Y 0.07fF
C22893 INVX1_LOC_425/Y INVX1_LOC_159/Y 0.01fF
C22894 INVX1_LOC_93/Y INVX1_LOC_379/A 0.07fF
C22895 NAND2X1_LOC_708/A INVX1_LOC_48/Y 0.01fF
C22896 NAND2X1_LOC_159/a_36_24# INVX1_LOC_9/Y 0.00fF
C22897 INVX1_LOC_584/Y INVX1_LOC_62/Y 0.06fF
C22898 NAND2X1_LOC_521/Y INVX1_LOC_145/Y 0.07fF
C22899 INVX1_LOC_17/Y NAND2X1_LOC_627/a_36_24# -0.02fF
C22900 INVX1_LOC_93/Y INVX1_LOC_35/Y 3.63fF
C22901 INVX1_LOC_93/Y INVX1_LOC_304/A 0.03fF
C22902 INVX1_LOC_277/A INVX1_LOC_221/Y 0.00fF
C22903 NAND2X1_LOC_261/Y INVX1_LOC_100/Y 0.01fF
C22904 INVX1_LOC_117/Y NAND2X1_LOC_672/a_36_24# 0.01fF
C22905 INVX1_LOC_492/A INVX1_LOC_46/Y 0.55fF
C22906 INVX1_LOC_607/Y INVX1_LOC_66/A 0.07fF
C22907 INVX1_LOC_147/A INVX1_LOC_496/A 0.02fF
C22908 INVX1_LOC_206/Y INVX1_LOC_291/Y 0.03fF
C22909 NAND2X1_LOC_371/a_36_24# NAND2X1_LOC_372/Y 0.01fF
C22910 VDD INVX1_LOC_636/A 0.00fF
C22911 INVX1_LOC_410/A INVX1_LOC_99/Y 0.01fF
C22912 NAND2X1_LOC_788/a_36_24# INVX1_LOC_66/A 0.01fF
C22913 INVX1_LOC_99/Y INVX1_LOC_420/A 0.00fF
C22914 INVX1_LOC_85/Y NAND2X1_LOC_214/a_36_24# 0.00fF
C22915 NAND2X1_LOC_615/Y INVX1_LOC_600/A 0.04fF
C22916 NAND2X1_LOC_301/B INVX1_LOC_686/A 0.07fF
C22917 INVX1_LOC_54/Y INVX1_LOC_421/A 0.10fF
C22918 INVX1_LOC_345/Y INVX1_LOC_32/Y 0.01fF
C22919 INVX1_LOC_170/Y INVX1_LOC_99/Y 0.03fF
C22920 INVX1_LOC_578/A INVX1_LOC_634/Y 0.74fF
C22921 INVX1_LOC_469/Y INVX1_LOC_359/Y 0.01fF
C22922 NAND2X1_LOC_332/B INVX1_LOC_479/A 0.01fF
C22923 INVX1_LOC_367/A INVX1_LOC_518/Y 0.04fF
C22924 NAND2X1_LOC_173/Y INVX1_LOC_74/Y 0.01fF
C22925 INVX1_LOC_58/Y INVX1_LOC_178/A 0.01fF
C22926 INVX1_LOC_171/A INVX1_LOC_6/Y 0.35fF
C22927 NAND2X1_LOC_353/a_36_24# INVX1_LOC_353/A 0.00fF
C22928 NAND2X1_LOC_770/B INVX1_LOC_89/Y 0.14fF
C22929 INVX1_LOC_450/A INVX1_LOC_443/A 0.55fF
C22930 INVX1_LOC_202/Y INVX1_LOC_551/A 0.00fF
C22931 INVX1_LOC_93/Y NAND2X1_LOC_448/B 0.03fF
C22932 NAND2X1_LOC_184/Y INVX1_LOC_387/Y 0.04fF
C22933 NAND2X1_LOC_177/a_36_24# INVX1_LOC_74/Y 0.01fF
C22934 INVX1_LOC_50/Y NAND2X1_LOC_753/Y 0.08fF
C22935 INVX1_LOC_58/Y NAND2X1_LOC_76/A 0.02fF
C22936 INVX1_LOC_682/A INVX1_LOC_116/Y 0.02fF
C22937 INVX1_LOC_93/Y INVX1_LOC_620/A 0.03fF
C22938 INVX1_LOC_399/Y INVX1_LOC_99/Y 0.03fF
C22939 INVX1_LOC_353/A INVX1_LOC_155/Y 0.06fF
C22940 NAND2X1_LOC_106/Y NAND2X1_LOC_128/A 0.03fF
C22941 INVX1_LOC_421/A NAND2X1_LOC_292/Y 0.02fF
C22942 INVX1_LOC_21/Y INVX1_LOC_502/A 0.07fF
C22943 INVX1_LOC_35/Y NAND2X1_LOC_334/B 0.08fF
C22944 INVX1_LOC_69/Y INVX1_LOC_656/A 0.04fF
C22945 INVX1_LOC_125/Y INVX1_LOC_479/A 0.01fF
C22946 NAND2X1_LOC_320/Y INVX1_LOC_114/A 0.00fF
C22947 NAND2X1_LOC_387/Y NAND2X1_LOC_698/Y 0.04fF
C22948 NAND2X1_LOC_413/Y INVX1_LOC_100/Y 0.33fF
C22949 NAND2X1_LOC_184/Y INVX1_LOC_49/Y -0.00fF
C22950 INVX1_LOC_449/A INVX1_LOC_62/Y 0.08fF
C22951 INVX1_LOC_31/Y NAND2X1_LOC_424/a_36_24# 0.00fF
C22952 INVX1_LOC_176/A NAND2X1_LOC_66/Y 0.02fF
C22953 INVX1_LOC_254/Y INVX1_LOC_242/Y 0.07fF
C22954 INVX1_LOC_662/Y INVX1_LOC_655/A 0.03fF
C22955 INVX1_LOC_35/Y NAND2X1_LOC_487/a_36_24# 0.01fF
C22956 NAND2X1_LOC_837/A NAND2X1_LOC_825/a_36_24# 0.02fF
C22957 NAND2X1_LOC_274/B INVX1_LOC_665/Y 0.01fF
C22958 INVX1_LOC_449/A NAND2X1_LOC_844/A 0.04fF
C22959 INVX1_LOC_410/A INVX1_LOC_47/Y 0.01fF
C22960 NAND2X1_LOC_27/a_36_24# INVX1_LOC_223/Y 0.00fF
C22961 INVX1_LOC_117/Y INVX1_LOC_245/A 0.10fF
C22962 INVX1_LOC_17/Y INVX1_LOC_41/Y 11.81fF
C22963 INVX1_LOC_262/Y INPUT_4 0.01fF
C22964 INVX1_LOC_202/Y INVX1_LOC_75/Y 0.02fF
C22965 NAND2X1_LOC_97/B INVX1_LOC_270/Y 0.02fF
C22966 INVX1_LOC_31/Y INVX1_LOC_652/A 0.04fF
C22967 INVX1_LOC_11/Y INVX1_LOC_588/A 0.06fF
C22968 INVX1_LOC_63/Y NAND2X1_LOC_236/a_36_24# 0.00fF
C22969 NAND2X1_LOC_97/B INVX1_LOC_92/A 0.03fF
C22970 INVX1_LOC_522/A INVX1_LOC_479/A 0.03fF
C22971 INVX1_LOC_471/Y INVX1_LOC_338/Y 0.13fF
C22972 INVX1_LOC_50/Y INVX1_LOC_483/A 0.01fF
C22973 NAND2X1_LOC_615/B INVX1_LOC_211/A 0.01fF
C22974 INVX1_LOC_328/Y INVX1_LOC_9/Y 0.03fF
C22975 NAND2X1_LOC_531/Y NAND2X1_LOC_631/B 0.12fF
C22976 INVX1_LOC_518/A INVX1_LOC_9/Y 0.11fF
C22977 INVX1_LOC_170/Y NAND2X1_LOC_66/Y 0.03fF
C22978 INVX1_LOC_373/Y INVX1_LOC_501/A 0.28fF
C22979 NAND2X1_LOC_128/B INVX1_LOC_479/A 0.19fF
C22980 INVX1_LOC_82/Y INVX1_LOC_85/A 0.05fF
C22981 INVX1_LOC_347/Y INVX1_LOC_62/Y 0.03fF
C22982 INVX1_LOC_482/A INVX1_LOC_109/Y 0.03fF
C22983 INVX1_LOC_49/Y INVX1_LOC_75/Y 0.06fF
C22984 NAND2X1_LOC_628/Y INVX1_LOC_79/A 0.04fF
C22985 INVX1_LOC_62/Y INVX1_LOC_328/Y 0.08fF
C22986 NAND2X1_LOC_242/A NAND2X1_LOC_241/B 0.06fF
C22987 NAND2X1_LOC_239/a_36_24# NAND2X1_LOC_164/Y 0.00fF
C22988 INVX1_LOC_479/A INVX1_LOC_242/Y 0.07fF
C22989 INVX1_LOC_100/Y NAND2X1_LOC_488/Y 0.04fF
C22990 VDD INVX1_LOC_269/Y 0.31fF
C22991 INVX1_LOC_151/Y INVX1_LOC_45/Y 0.01fF
C22992 INVX1_LOC_3/Y INVX1_LOC_33/Y 0.01fF
C22993 INVX1_LOC_49/Y NAND2X1_LOC_271/A 0.07fF
C22994 INVX1_LOC_307/Y INVX1_LOC_72/Y 0.04fF
C22995 INVX1_LOC_75/Y INVX1_LOC_17/A 0.03fF
C22996 INPUT_0 INVX1_LOC_442/A 0.03fF
C22997 INVX1_LOC_416/Y INVX1_LOC_578/A 0.03fF
C22998 INVX1_LOC_194/A INVX1_LOC_109/Y 0.01fF
C22999 INVX1_LOC_79/A NAND2X1_LOC_832/A 0.03fF
C23000 NAND2X1_LOC_331/A NAND2X1_LOC_163/B 0.01fF
C23001 INVX1_LOC_629/A NAND2X1_LOC_173/Y 0.28fF
C23002 INVX1_LOC_74/Y INVX1_LOC_354/A 0.04fF
C23003 NAND2X1_LOC_765/a_36_24# INVX1_LOC_53/Y 0.00fF
C23004 INVX1_LOC_317/Y NAND2X1_LOC_370/A 0.25fF
C23005 NAND2X1_LOC_108/Y NAND2X1_LOC_142/Y 0.70fF
C23006 INVX1_LOC_206/Y INVX1_LOC_551/Y 0.10fF
C23007 INVX1_LOC_224/Y INVX1_LOC_270/A 0.02fF
C23008 NAND2X1_LOC_396/Y INVX1_LOC_443/A 0.59fF
C23009 VDD INVX1_LOC_320/A 0.00fF
C23010 VDD INVX1_LOC_29/Y 0.39fF
C23011 NAND2X1_LOC_164/Y NAND2X1_LOC_238/a_36_24# 0.00fF
C23012 INVX1_LOC_160/Y INVX1_LOC_286/Y 0.04fF
C23013 NAND2X1_LOC_545/B INVX1_LOC_412/A 0.02fF
C23014 INVX1_LOC_560/Y INVX1_LOC_252/Y 0.03fF
C23015 NAND2X1_LOC_756/Y INVX1_LOC_586/A 0.96fF
C23016 INVX1_LOC_272/Y INVX1_LOC_45/Y 0.01fF
C23017 INVX1_LOC_293/Y INVX1_LOC_586/A 0.03fF
C23018 INVX1_LOC_254/Y INVX1_LOC_301/A 0.00fF
C23019 INVX1_LOC_457/Y INVX1_LOC_99/Y -0.00fF
C23020 INVX1_LOC_249/A INVX1_LOC_249/Y 0.01fF
C23021 NAND2X1_LOC_173/Y INVX1_LOC_566/A 0.02fF
C23022 NAND2X1_LOC_715/a_36_24# INVX1_LOC_367/A 0.00fF
C23023 INPUT_0 INVX1_LOC_116/Y 0.07fF
C23024 INVX1_LOC_224/Y INVX1_LOC_211/Y 0.05fF
C23025 INVX1_LOC_395/A INVX1_LOC_379/A 0.65fF
C23026 INVX1_LOC_249/A NAND2X1_LOC_122/Y 0.28fF
C23027 INVX1_LOC_133/Y NAND2X1_LOC_846/A 0.02fF
C23028 INVX1_LOC_84/A INPUT_2 0.03fF
C23029 INVX1_LOC_291/A INVX1_LOC_524/Y 0.12fF
C23030 INVX1_LOC_435/Y INVX1_LOC_442/Y 0.10fF
C23031 NAND2X1_LOC_45/Y INVX1_LOC_54/Y 1.48fF
C23032 INVX1_LOC_447/Y NAND2X1_LOC_498/Y 0.22fF
C23033 INVX1_LOC_551/Y INVX1_LOC_686/A 0.10fF
C23034 INVX1_LOC_395/A INVX1_LOC_35/Y 0.60fF
C23035 INVX1_LOC_395/A INVX1_LOC_304/A 0.01fF
C23036 INVX1_LOC_449/A INVX1_LOC_218/A -0.01fF
C23037 INPUT_3 INVX1_LOC_294/Y 0.01fF
C23038 INPUT_3 INVX1_LOC_486/Y 0.13fF
C23039 INVX1_LOC_160/A INVX1_LOC_586/A 0.03fF
C23040 VDD INVX1_LOC_470/Y 0.21fF
C23041 NAND2X1_LOC_498/Y NAND2X1_LOC_602/A 0.06fF
C23042 INVX1_LOC_68/Y INVX1_LOC_155/Y 0.03fF
C23043 INVX1_LOC_224/Y INVX1_LOC_46/Y 0.07fF
C23044 INVX1_LOC_413/Y INVX1_LOC_391/Y 0.11fF
C23045 INVX1_LOC_628/A NAND2X1_LOC_173/Y 0.03fF
C23046 NAND2X1_LOC_93/Y NAND2X1_LOC_753/Y 0.12fF
C23047 INVX1_LOC_166/A NAND2X1_LOC_320/a_36_24# 0.00fF
C23048 INVX1_LOC_425/A INVX1_LOC_129/A 0.03fF
C23049 INVX1_LOC_362/Y INVX1_LOC_35/Y 0.12fF
C23050 INVX1_LOC_567/A INVX1_LOC_89/A 0.14fF
C23051 INVX1_LOC_166/A INVX1_LOC_127/A 0.03fF
C23052 NAND2X1_LOC_336/B NAND2X1_LOC_545/B 0.00fF
C23053 INVX1_LOC_54/Y NAND2X1_LOC_498/Y 0.07fF
C23054 INVX1_LOC_435/Y INVX1_LOC_671/A 0.01fF
C23055 INVX1_LOC_257/Y INVX1_LOC_66/A 0.02fF
C23056 NAND2X1_LOC_175/a_36_24# INVX1_LOC_99/Y 0.00fF
C23057 INVX1_LOC_393/A INVX1_LOC_50/Y 0.01fF
C23058 INVX1_LOC_578/A INVX1_LOC_46/Y 0.09fF
C23059 INVX1_LOC_395/A INVX1_LOC_620/A 0.07fF
C23060 INVX1_LOC_588/Y NAND2X1_LOC_122/Y 0.03fF
C23061 VDD INVX1_LOC_300/Y 0.35fF
C23062 INVX1_LOC_681/A INVX1_LOC_235/Y 0.00fF
C23063 INVX1_LOC_457/Y INVX1_LOC_47/Y 0.00fF
C23064 INVX1_LOC_80/A INVX1_LOC_670/Y 0.07fF
C23065 INVX1_LOC_442/Y INVX1_LOC_596/A 0.07fF
C23066 INVX1_LOC_429/A NAND2X1_LOC_344/B 0.00fF
C23067 INVX1_LOC_229/Y INVX1_LOC_228/A 0.18fF
C23068 INVX1_LOC_250/Y INVX1_LOC_155/Y 0.04fF
C23069 INVX1_LOC_400/Y INVX1_LOC_89/Y 0.07fF
C23070 INVX1_LOC_683/Y INVX1_LOC_35/Y 0.03fF
C23071 INVX1_LOC_20/Y INVX1_LOC_254/Y 0.03fF
C23072 INVX1_LOC_366/Y INVX1_LOC_307/A 0.00fF
C23073 INVX1_LOC_54/A INVX1_LOC_183/A 0.01fF
C23074 NAND2X1_LOC_837/B INVX1_LOC_59/A 0.11fF
C23075 NAND2X1_LOC_336/B INVX1_LOC_98/Y 0.13fF
C23076 INVX1_LOC_584/A INVX1_LOC_501/A 0.00fF
C23077 NAND2X1_LOC_324/B INVX1_LOC_256/A 0.03fF
C23078 INVX1_LOC_80/A INVX1_LOC_506/Y 0.01fF
C23079 INVX1_LOC_469/Y NAND2X1_LOC_173/Y 0.00fF
C23080 INVX1_LOC_45/Y INVX1_LOC_6/Y 0.23fF
C23081 INVX1_LOC_286/Y NAND2X1_LOC_267/A 0.03fF
C23082 INPUT_0 INVX1_LOC_179/A 0.03fF
C23083 VDD INVX1_LOC_100/Y 2.80fF
C23084 INVX1_LOC_335/Y INVX1_LOC_17/Y 5.29fF
C23085 NAND2X1_LOC_486/B INVX1_LOC_387/Y 0.05fF
C23086 INVX1_LOC_291/A INVX1_LOC_93/Y 0.35fF
C23087 INVX1_LOC_21/Y INVX1_LOC_17/Y 0.28fF
C23088 INVX1_LOC_53/Y INVX1_LOC_259/Y 0.03fF
C23089 INVX1_LOC_571/A NAND2X1_LOC_728/B 0.01fF
C23090 INVX1_LOC_384/A INVX1_LOC_66/A 0.07fF
C23091 INVX1_LOC_401/Y INPUT_1 0.18fF
C23092 INVX1_LOC_367/A INVX1_LOC_118/A 0.07fF
C23093 INVX1_LOC_11/Y INVX1_LOC_670/Y 0.00fF
C23094 INVX1_LOC_31/A INVX1_LOC_6/Y 0.11fF
C23095 INVX1_LOC_197/A INVX1_LOC_50/Y 0.01fF
C23096 INVX1_LOC_301/A INVX1_LOC_479/A 0.07fF
C23097 INPUT_0 NAND2X1_LOC_262/a_36_24# 0.00fF
C23098 INVX1_LOC_3/Y INVX1_LOC_25/A 0.04fF
C23099 INVX1_LOC_20/Y INVX1_LOC_592/Y 0.01fF
C23100 INPUT_3 INVX1_LOC_6/Y 0.03fF
C23101 NAND2X1_LOC_707/A INVX1_LOC_338/Y 0.37fF
C23102 NAND2X1_LOC_800/a_36_24# INVX1_LOC_630/A 0.02fF
C23103 NAND2X1_LOC_97/B INPUT_1 0.00fF
C23104 NAND2X1_LOC_241/B INVX1_LOC_79/A 0.57fF
C23105 VDD INVX1_LOC_74/Y 1.20fF
C23106 NAND2X1_LOC_638/A INVX1_LOC_315/A 0.06fF
C23107 INVX1_LOC_228/Y INVX1_LOC_100/Y 0.16fF
C23108 NAND2X1_LOC_43/Y INVX1_LOC_176/A 0.03fF
C23109 INVX1_LOC_145/Y INVX1_LOC_159/A 0.00fF
C23110 INVX1_LOC_35/Y INVX1_LOC_189/Y 0.01fF
C23111 INVX1_LOC_434/A NAND2X1_LOC_252/a_36_24# 0.01fF
C23112 INVX1_LOC_93/A INVX1_LOC_333/A 0.03fF
C23113 NAND2X1_LOC_187/Y INVX1_LOC_99/Y 0.02fF
C23114 INVX1_LOC_53/Y NAND2X1_LOC_707/B 0.02fF
C23115 VDD INVX1_LOC_483/Y 0.51fF
C23116 INVX1_LOC_266/Y INVX1_LOC_9/Y 0.00fF
C23117 INVX1_LOC_254/Y INVX1_LOC_300/A 0.07fF
C23118 INVX1_LOC_243/A INVX1_LOC_382/A 0.01fF
C23119 INVX1_LOC_54/Y INVX1_LOC_99/Y 2.21fF
C23120 INVX1_LOC_490/A NAND2X1_LOC_296/Y 0.01fF
C23121 NAND2X1_LOC_179/Y INPUT_1 0.01fF
C23122 INVX1_LOC_53/Y NAND2X1_LOC_697/a_36_24# 0.00fF
C23123 INVX1_LOC_80/A INVX1_LOC_253/Y 0.26fF
C23124 INVX1_LOC_609/A INVX1_LOC_54/Y 0.01fF
C23125 INVX1_LOC_459/Y INVX1_LOC_114/A 0.02fF
C23126 INVX1_LOC_53/Y INVX1_LOC_204/Y 0.00fF
C23127 INVX1_LOC_625/A NAND2X1_LOC_333/B 0.32fF
C23128 INVX1_LOC_381/A INVX1_LOC_339/Y 0.03fF
C23129 INVX1_LOC_224/Y INVX1_LOC_75/A 0.02fF
C23130 INVX1_LOC_228/Y INVX1_LOC_74/Y 0.03fF
C23131 NAND2X1_LOC_231/A INVX1_LOC_90/Y 0.00fF
C23132 INVX1_LOC_17/Y NAND2X1_LOC_267/A 0.40fF
C23133 INVX1_LOC_448/A INVX1_LOC_66/A 0.07fF
C23134 INVX1_LOC_31/Y INVX1_LOC_379/A 0.07fF
C23135 INVX1_LOC_468/Y INVX1_LOC_46/Y 0.03fF
C23136 INVX1_LOC_510/Y INVX1_LOC_100/Y 0.07fF
C23137 INVX1_LOC_335/A INVX1_LOC_514/A 0.01fF
C23138 INVX1_LOC_521/Y INVX1_LOC_62/Y 0.01fF
C23139 INPUT_1 INVX1_LOC_510/A 0.08fF
C23140 INVX1_LOC_80/A INVX1_LOC_63/Y 5.86fF
C23141 INVX1_LOC_596/A INVX1_LOC_482/Y 0.08fF
C23142 NAND2X1_LOC_768/A INVX1_LOC_63/Y 0.02fF
C23143 INVX1_LOC_31/Y INVX1_LOC_35/Y 7.63fF
C23144 NAND2X1_LOC_180/B NAND2X1_LOC_545/A 0.01fF
C23145 INVX1_LOC_93/Y NAND2X1_LOC_837/B 0.03fF
C23146 INVX1_LOC_145/Y INVX1_LOC_66/A 0.09fF
C23147 NAND2X1_LOC_102/a_36_24# NAND2X1_LOC_542/A 0.00fF
C23148 INVX1_LOC_89/Y INVX1_LOC_125/A 0.01fF
C23149 INVX1_LOC_359/Y INVX1_LOC_48/Y 0.01fF
C23150 INVX1_LOC_93/Y INVX1_LOC_360/A 0.04fF
C23151 NAND2X1_LOC_173/Y INVX1_LOC_460/A 0.02fF
C23152 INVX1_LOC_657/A INVX1_LOC_59/A 0.03fF
C23153 INVX1_LOC_93/Y INVX1_LOC_118/A 0.01fF
C23154 INVX1_LOC_510/Y INVX1_LOC_74/Y 0.11fF
C23155 NAND2X1_LOC_274/B INVX1_LOC_134/Y 0.07fF
C23156 INVX1_LOC_298/A INPUT_4 0.10fF
C23157 INVX1_LOC_12/Y INVX1_LOC_484/Y 0.01fF
C23158 NAND2X1_LOC_835/A INVX1_LOC_656/A 0.00fF
C23159 INVX1_LOC_76/Y INVX1_LOC_75/Y 0.03fF
C23160 INVX1_LOC_53/Y INVX1_LOC_114/A 0.03fF
C23161 INVX1_LOC_501/A INVX1_LOC_537/A 0.01fF
C23162 INVX1_LOC_412/Y INVX1_LOC_92/A 0.03fF
C23163 INVX1_LOC_608/A NAND2X1_LOC_496/a_36_24# 0.00fF
C23164 INVX1_LOC_49/Y NAND2X1_LOC_462/a_36_24# 0.00fF
C23165 INVX1_LOC_48/Y INVX1_LOC_187/Y 0.04fF
C23166 INVX1_LOC_54/Y INVX1_LOC_47/Y 0.26fF
C23167 INVX1_LOC_281/Y INVX1_LOC_245/A 0.49fF
C23168 INVX1_LOC_300/Y INVX1_LOC_684/A 0.00fF
C23169 INVX1_LOC_54/Y NAND2X1_LOC_557/B 0.03fF
C23170 INVX1_LOC_11/Y INVX1_LOC_63/Y 0.14fF
C23171 INVX1_LOC_20/Y INVX1_LOC_479/A 0.22fF
C23172 INVX1_LOC_35/Y INVX1_LOC_682/Y 0.07fF
C23173 INVX1_LOC_520/Y INVX1_LOC_117/Y 0.03fF
C23174 INVX1_LOC_183/A NAND2X1_LOC_84/B 0.32fF
C23175 NAND2X1_LOC_770/B INVX1_LOC_44/Y 0.06fF
C23176 NAND2X1_LOC_406/B INVX1_LOC_259/Y 0.14fF
C23177 INVX1_LOC_575/Y INVX1_LOC_569/Y 0.01fF
C23178 INVX1_LOC_335/A INVX1_LOC_534/Y 0.09fF
C23179 NAND2X1_LOC_837/A INVX1_LOC_6/Y 0.70fF
C23180 INVX1_LOC_451/A INVX1_LOC_405/Y 0.09fF
C23181 INVX1_LOC_120/Y INVX1_LOC_46/Y 0.08fF
C23182 NAND2X1_LOC_513/A INVX1_LOC_652/Y 0.03fF
C23183 INVX1_LOC_172/A INVX1_LOC_9/Y 0.24fF
C23184 INVX1_LOC_324/Y INVX1_LOC_327/A 0.01fF
C23185 INVX1_LOC_679/Y NAND2X1_LOC_248/B 0.03fF
C23186 NAND2X1_LOC_160/a_36_24# INVX1_LOC_62/Y 0.00fF
C23187 INVX1_LOC_176/A NAND2X1_LOC_627/Y 0.03fF
C23188 INVX1_LOC_76/Y NAND2X1_LOC_271/A 0.02fF
C23189 NAND2X1_LOC_755/B INVX1_LOC_621/A 0.06fF
C23190 INVX1_LOC_501/A INVX1_LOC_496/Y 0.02fF
C23191 NAND2X1_LOC_843/A INVX1_LOC_100/Y 0.04fF
C23192 INVX1_LOC_105/Y INVX1_LOC_9/Y 0.17fF
C23193 INVX1_LOC_686/A INVX1_LOC_634/Y 0.11fF
C23194 INVX1_LOC_460/Y INVX1_LOC_114/A 0.02fF
C23195 INVX1_LOC_545/A INVX1_LOC_41/Y 0.00fF
C23196 INVX1_LOC_54/Y INVX1_LOC_119/Y 0.03fF
C23197 INVX1_LOC_116/A INVX1_LOC_74/Y 0.24fF
C23198 INVX1_LOC_99/Y INVX1_LOC_388/A 0.01fF
C23199 NAND2X1_LOC_56/a_36_24# INVX1_LOC_211/A -0.01fF
C23200 INVX1_LOC_361/Y INVX1_LOC_519/Y 0.04fF
C23201 INVX1_LOC_54/Y NAND2X1_LOC_66/Y 0.03fF
C23202 INVX1_LOC_300/A INVX1_LOC_479/A 0.08fF
C23203 INVX1_LOC_617/Y INVX1_LOC_92/A 0.07fF
C23204 INVX1_LOC_103/Y INVX1_LOC_100/Y 0.56fF
C23205 INVX1_LOC_682/A INVX1_LOC_69/Y 0.00fF
C23206 INVX1_LOC_58/Y NAND2X1_LOC_91/a_36_24# 0.01fF
C23207 INVX1_LOC_74/Y INVX1_LOC_509/A 0.27fF
C23208 INVX1_LOC_77/Y INVX1_LOC_351/A 0.04fF
C23209 INVX1_LOC_157/A INVX1_LOC_245/A 0.00fF
C23210 INVX1_LOC_455/A INVX1_LOC_74/A 0.01fF
C23211 INVX1_LOC_100/Y INVX1_LOC_68/A 0.01fF
C23212 INVX1_LOC_382/A NAND2X1_LOC_631/B 0.03fF
C23213 NAND2X1_LOC_720/A INVX1_LOC_635/Y 0.03fF
C23214 NAND2X1_LOC_451/B INVX1_LOC_259/Y 0.03fF
C23215 INVX1_LOC_242/Y INVX1_LOC_188/A 0.00fF
C23216 INVX1_LOC_58/Y INVX1_LOC_245/A 0.02fF
C23217 INVX1_LOC_77/Y INVX1_LOC_90/Y 0.04fF
C23218 INVX1_LOC_376/A INVX1_LOC_26/Y 0.12fF
C23219 INVX1_LOC_469/Y INVX1_LOC_354/A 0.00fF
C23220 VDD NAND2X1_LOC_591/B 0.05fF
C23221 INVX1_LOC_48/Y NAND2X1_LOC_832/A 0.03fF
C23222 NAND2X1_LOC_301/B INVX1_LOC_376/Y 0.03fF
C23223 NAND2X1_LOC_242/A VDD 0.09fF
C23224 INVX1_LOC_502/A INVX1_LOC_26/Y 0.07fF
C23225 INVX1_LOC_62/Y INVX1_LOC_224/A 0.01fF
C23226 INVX1_LOC_179/A INVX1_LOC_211/A 0.47fF
C23227 INVX1_LOC_95/A INVX1_LOC_91/Y 0.01fF
C23228 INVX1_LOC_179/A INVX1_LOC_64/Y 0.03fF
C23229 NAND2X1_LOC_534/Y NAND2X1_LOC_498/Y 0.01fF
C23230 INVX1_LOC_49/Y NAND2X1_LOC_98/B 0.06fF
C23231 INVX1_LOC_438/Y INVX1_LOC_446/Y 0.03fF
C23232 NAND2X1_LOC_788/A NAND2X1_LOC_727/a_36_24# 0.00fF
C23233 VDD INVX1_LOC_207/A -0.00fF
C23234 INVX1_LOC_133/Y INVX1_LOC_574/Y 0.01fF
C23235 INVX1_LOC_257/Y INVX1_LOC_442/A 0.03fF
C23236 NAND2X1_LOC_331/A INVX1_LOC_584/Y 0.02fF
C23237 INVX1_LOC_206/Y INVX1_LOC_558/A 0.01fF
C23238 INVX1_LOC_446/A INVX1_LOC_80/A 0.07fF
C23239 VDD INVX1_LOC_566/A 0.00fF
C23240 INVX1_LOC_438/Y INVX1_LOC_384/A 0.19fF
C23241 INVX1_LOC_74/Y INVX1_LOC_635/Y 0.03fF
C23242 NAND2X1_LOC_7/Y INVX1_LOC_12/Y 0.01fF
C23243 INVX1_LOC_224/Y NAND2X1_LOC_318/A 0.01fF
C23244 NAND2X1_LOC_758/a_36_24# INVX1_LOC_53/Y 0.00fF
C23245 INVX1_LOC_206/Y INVX1_LOC_270/A 0.60fF
C23246 INVX1_LOC_301/A INVX1_LOC_12/Y 0.01fF
C23247 INVX1_LOC_558/A NAND2X1_LOC_516/a_36_24# 0.01fF
C23248 INVX1_LOC_395/A INVX1_LOC_291/A 0.01fF
C23249 INVX1_LOC_243/A VDD 0.00fF
C23250 NAND2X1_LOC_725/a_36_24# INVX1_LOC_523/A 0.00fF
C23251 INVX1_LOC_21/Y NAND2X1_LOC_88/Y 0.23fF
C23252 INVX1_LOC_53/Y NAND2X1_LOC_457/A 0.03fF
C23253 INVX1_LOC_558/A INVX1_LOC_242/A 0.07fF
C23254 INVX1_LOC_53/Y INVX1_LOC_554/Y 0.01fF
C23255 INVX1_LOC_446/A INVX1_LOC_11/Y 0.07fF
C23256 INVX1_LOC_560/A NAND2X1_LOC_307/A 0.02fF
C23257 VDD NAND2X1_LOC_57/Y -0.00fF
C23258 INVX1_LOC_418/A INVX1_LOC_686/A 0.14fF
C23259 NAND2X1_LOC_773/A INVX1_LOC_366/A 0.01fF
C23260 INVX1_LOC_438/A NAND2X1_LOC_416/Y 0.03fF
C23261 NAND2X1_LOC_543/B INVX1_LOC_349/A 0.01fF
C23262 INVX1_LOC_206/Y NAND2X1_LOC_755/B 0.10fF
C23263 INVX1_LOC_53/Y INVX1_LOC_547/Y 0.26fF
C23264 NAND2X1_LOC_513/Y INVX1_LOC_558/Y 0.01fF
C23265 INVX1_LOC_374/A INVX1_LOC_80/A 0.04fF
C23266 INVX1_LOC_257/Y INVX1_LOC_116/Y 0.01fF
C23267 NAND2X1_LOC_498/Y INVX1_LOC_371/Y 0.01fF
C23268 INVX1_LOC_224/Y INVX1_LOC_202/Y 0.00fF
C23269 INVX1_LOC_211/Y INVX1_LOC_206/Y 0.01fF
C23270 INVX1_LOC_9/Y INVX1_LOC_109/Y 0.10fF
C23271 INVX1_LOC_578/A INVX1_LOC_115/A 0.09fF
C23272 INVX1_LOC_298/Y INVX1_LOC_290/Y 0.00fF
C23273 VDD INVX1_LOC_469/Y 0.81fF
C23274 VDD INVX1_LOC_350/Y 0.39fF
C23275 NAND2X1_LOC_475/A INVX1_LOC_54/Y 0.07fF
C23276 INVX1_LOC_20/Y INVX1_LOC_372/Y 0.05fF
C23277 NAND2X1_LOC_756/Y NAND2X1_LOC_791/B 0.02fF
C23278 NAND2X1_LOC_750/Y NAND2X1_LOC_60/a_36_24# 0.00fF
C23279 INVX1_LOC_17/Y INVX1_LOC_255/Y 1.47fF
C23280 INVX1_LOC_578/A NAND2X1_LOC_703/a_36_24# 0.00fF
C23281 INVX1_LOC_395/A NAND2X1_LOC_837/B 0.01fF
C23282 INVX1_LOC_412/Y INPUT_1 0.03fF
C23283 NAND2X1_LOC_731/a_36_24# INVX1_LOC_575/Y 0.00fF
C23284 INVX1_LOC_420/Y INVX1_LOC_48/Y 0.00fF
C23285 INVX1_LOC_578/A INVX1_LOC_349/Y 0.00fF
C23286 INVX1_LOC_142/A NAND2X1_LOC_677/Y 0.01fF
C23287 NAND2X1_LOC_505/Y INVX1_LOC_35/Y 0.01fF
C23288 INVX1_LOC_293/Y INVX1_LOC_294/Y 0.09fF
C23289 INVX1_LOC_51/Y INVX1_LOC_379/A 0.07fF
C23290 VDD NAND2X1_LOC_181/A 0.15fF
C23291 INVX1_LOC_206/Y NAND2X1_LOC_196/a_36_24# 0.00fF
C23292 INVX1_LOC_400/Y INVX1_LOC_194/Y 0.16fF
C23293 INVX1_LOC_20/Y INVX1_LOC_12/Y 0.10fF
C23294 INVX1_LOC_52/Y INVX1_LOC_93/Y 0.04fF
C23295 NAND2X1_LOC_787/a_36_24# INVX1_LOC_362/Y 0.00fF
C23296 INVX1_LOC_206/Y INVX1_LOC_46/Y 0.79fF
C23297 INVX1_LOC_11/Y INVX1_LOC_374/A 0.03fF
C23298 INVX1_LOC_447/Y INVX1_LOC_502/Y 0.02fF
C23299 INVX1_LOC_395/A INVX1_LOC_208/A 0.05fF
C23300 INVX1_LOC_51/Y INVX1_LOC_35/Y 0.13fF
C23301 INVX1_LOC_438/Y INVX1_LOC_433/A 0.03fF
C23302 INVX1_LOC_574/Y INVX1_LOC_581/A 0.00fF
C23303 INVX1_LOC_554/A INVX1_LOC_9/Y 0.21fF
C23304 INVX1_LOC_238/Y INVX1_LOC_212/Y 0.02fF
C23305 INVX1_LOC_288/Y INVX1_LOC_677/Y 0.42fF
C23306 INVX1_LOC_171/Y INVX1_LOC_99/Y 0.09fF
C23307 INVX1_LOC_62/Y INVX1_LOC_109/Y 1.66fF
C23308 INVX1_LOC_648/Y INVX1_LOC_46/Y 0.02fF
C23309 INVX1_LOC_444/Y INVX1_LOC_175/A 0.03fF
C23310 INVX1_LOC_219/Y INVX1_LOC_384/A 0.02fF
C23311 INVX1_LOC_257/Y INVX1_LOC_255/A 0.01fF
C23312 INVX1_LOC_451/A INVX1_LOC_172/Y 0.04fF
C23313 INPUT_0 INVX1_LOC_69/Y 0.04fF
C23314 INVX1_LOC_266/A INVX1_LOC_35/Y 0.14fF
C23315 INVX1_LOC_193/A INVX1_LOC_425/A 0.01fF
C23316 INVX1_LOC_603/Y INVX1_LOC_97/Y 0.03fF
C23317 INVX1_LOC_266/A INVX1_LOC_304/A 0.21fF
C23318 NAND2X1_LOC_197/a_36_24# INVX1_LOC_600/A 0.00fF
C23319 NAND2X1_LOC_498/Y INVX1_LOC_89/Y 0.11fF
C23320 VDD NAND2X1_LOC_558/B 0.02fF
C23321 INVX1_LOC_51/Y NAND2X1_LOC_448/B 0.54fF
C23322 INVX1_LOC_570/A INVX1_LOC_89/Y 0.07fF
C23323 INVX1_LOC_53/Y NAND2X1_LOC_144/a_36_24# 0.00fF
C23324 INVX1_LOC_587/A INVX1_LOC_656/A 0.09fF
C23325 VDD INVX1_LOC_77/A -0.00fF
C23326 NAND2X1_LOC_516/Y INVX1_LOC_69/Y 0.00fF
C23327 INVX1_LOC_612/Y NAND2X1_LOC_780/A 0.13fF
C23328 INVX1_LOC_300/A INVX1_LOC_12/Y 0.03fF
C23329 VDD INVX1_LOC_79/A 2.00fF
C23330 INVX1_LOC_554/A INVX1_LOC_62/Y 0.03fF
C23331 INVX1_LOC_557/A INVX1_LOC_49/Y 0.15fF
C23332 INVX1_LOC_46/Y INVX1_LOC_242/A 0.03fF
C23333 INVX1_LOC_418/Y INVX1_LOC_134/Y 0.00fF
C23334 INVX1_LOC_617/Y INPUT_1 0.07fF
C23335 INVX1_LOC_609/A NAND2X1_LOC_677/Y 0.24fF
C23336 INVX1_LOC_336/Y INVX1_LOC_50/Y 0.02fF
C23337 NAND2X1_LOC_332/B INVX1_LOC_66/A 0.03fF
C23338 INVX1_LOC_113/Y INVX1_LOC_47/Y 0.03fF
C23339 VDD NAND2X1_LOC_631/B 0.08fF
C23340 INVX1_LOC_20/Y NAND2X1_LOC_333/A 0.14fF
C23341 INVX1_LOC_192/Y INVX1_LOC_242/Y 0.02fF
C23342 VDD INVX1_LOC_460/A -0.00fF
C23343 VDD NAND2X1_LOC_396/Y 0.01fF
C23344 NAND2X1_LOC_773/A INVX1_LOC_6/Y 0.01fF
C23345 INVX1_LOC_11/Y NAND2X1_LOC_499/a_36_24# 0.00fF
C23346 INVX1_LOC_51/Y INVX1_LOC_621/Y 0.05fF
C23347 INVX1_LOC_267/Y INVX1_LOC_50/Y 0.23fF
C23348 INVX1_LOC_145/Y INVX1_LOC_116/Y 0.00fF
C23349 INVX1_LOC_686/A INVX1_LOC_46/Y 0.07fF
C23350 INVX1_LOC_377/A INVX1_LOC_665/Y 0.10fF
C23351 NAND2X1_LOC_373/Y INVX1_LOC_479/A 0.11fF
C23352 INVX1_LOC_366/A NAND2X1_LOC_240/A 0.01fF
C23353 INVX1_LOC_17/Y INVX1_LOC_481/Y 0.01fF
C23354 INVX1_LOC_293/Y INVX1_LOC_6/Y 0.03fF
C23355 GATE_741 INVX1_LOC_168/Y 0.01fF
C23356 INVX1_LOC_166/A INVX1_LOC_519/A 0.01fF
C23357 NAND2X1_LOC_595/Y INVX1_LOC_665/Y 0.00fF
C23358 INVX1_LOC_21/Y INVX1_LOC_198/A 0.02fF
C23359 NAND2X1_LOC_387/Y INVX1_LOC_97/Y 0.01fF
C23360 INVX1_LOC_682/A INVX1_LOC_586/A 0.01fF
C23361 NAND2X1_LOC_320/a_36_24# INVX1_LOC_41/Y 0.01fF
C23362 INVX1_LOC_619/A NAND2X1_LOC_789/A 0.01fF
C23363 INVX1_LOC_304/Y INVX1_LOC_230/A 0.01fF
C23364 INVX1_LOC_127/A INVX1_LOC_41/Y 0.02fF
C23365 NAND2X1_LOC_179/Y INVX1_LOC_50/Y 0.01fF
C23366 INVX1_LOC_20/Y INVX1_LOC_276/Y 0.09fF
C23367 INVX1_LOC_553/A INVX1_LOC_479/A 0.01fF
C23368 NAND2X1_LOC_27/Y INVX1_LOC_178/A 0.03fF
C23369 NAND2X1_LOC_507/A INVX1_LOC_99/Y 0.01fF
C23370 INVX1_LOC_578/A INVX1_LOC_17/A 0.05fF
C23371 INVX1_LOC_435/A INVX1_LOC_295/Y 0.10fF
C23372 INVX1_LOC_607/Y NAND2X1_LOC_148/B 0.04fF
C23373 NAND2X1_LOC_111/Y INVX1_LOC_519/A 0.00fF
C23374 INVX1_LOC_145/A INVX1_LOC_29/Y 0.01fF
C23375 INVX1_LOC_93/Y INVX1_LOC_115/Y 0.03fF
C23376 INVX1_LOC_551/Y INVX1_LOC_376/Y 0.10fF
C23377 INVX1_LOC_51/Y INVX1_LOC_518/Y 0.04fF
C23378 INVX1_LOC_510/Y INVX1_LOC_79/A 0.13fF
C23379 INVX1_LOC_254/A INVX1_LOC_35/Y 0.01fF
C23380 NAND2X1_LOC_370/A INVX1_LOC_41/Y 0.00fF
C23381 INVX1_LOC_50/Y INVX1_LOC_510/A 0.01fF
C23382 NAND2X1_LOC_333/A INVX1_LOC_300/A 0.02fF
C23383 INVX1_LOC_126/Y INVX1_LOC_9/Y 0.01fF
C23384 INVX1_LOC_316/Y INVX1_LOC_340/A 0.01fF
C23385 INVX1_LOC_89/Y INVX1_LOC_99/Y 0.03fF
C23386 INVX1_LOC_93/Y INVX1_LOC_350/A 0.02fF
C23387 NAND2X1_LOC_122/Y INVX1_LOC_41/Y 0.02fF
C23388 INVX1_LOC_273/A INVX1_LOC_41/Y 0.01fF
C23389 INVX1_LOC_171/Y NAND2X1_LOC_66/Y 0.02fF
C23390 INVX1_LOC_607/Y INVX1_LOC_69/Y 0.11fF
C23391 NAND2X1_LOC_88/B INVX1_LOC_178/Y 0.01fF
C23392 INVX1_LOC_280/Y INVX1_LOC_50/Y 0.01fF
C23393 INVX1_LOC_300/A INVX1_LOC_188/A 0.03fF
C23394 NAND2X1_LOC_818/a_36_24# INVX1_LOC_9/Y 0.00fF
C23395 INVX1_LOC_20/Y INVX1_LOC_680/A 0.07fF
C23396 INVX1_LOC_503/Y INVX1_LOC_66/A 0.01fF
C23397 INVX1_LOC_201/A INVX1_LOC_69/Y 0.01fF
C23398 NAND2X1_LOC_673/B INVX1_LOC_6/Y 0.08fF
C23399 INVX1_LOC_468/Y INVX1_LOC_49/Y 0.03fF
C23400 NAND2X1_LOC_57/a_36_24# INVX1_LOC_63/Y 0.00fF
C23401 INVX1_LOC_525/Y INVX1_LOC_50/Y 0.43fF
C23402 INVX1_LOC_501/A INVX1_LOC_99/Y 0.60fF
C23403 INVX1_LOC_198/A INVX1_LOC_181/Y 0.05fF
C23404 INVX1_LOC_179/A INVX1_LOC_145/Y 0.03fF
C23405 INVX1_LOC_555/A INVX1_LOC_189/A 0.04fF
C23406 INVX1_LOC_65/A INVX1_LOC_159/Y 0.01fF
C23407 INVX1_LOC_117/Y NAND2X1_LOC_753/Y 0.07fF
C23408 NAND2X1_LOC_301/B NAND2X1_LOC_603/Y 0.01fF
C23409 INVX1_LOC_103/Y NAND2X1_LOC_181/A 0.10fF
C23410 INVX1_LOC_410/Y INVX1_LOC_92/A 0.00fF
C23411 INVX1_LOC_370/Y NAND2X1_LOC_274/B 0.00fF
C23412 NAND2X1_LOC_27/Y INVX1_LOC_58/Y 0.01fF
C23413 INVX1_LOC_375/A INVX1_LOC_92/A 0.03fF
C23414 INVX1_LOC_298/A INVX1_LOC_69/Y 0.11fF
C23415 NAND2X1_LOC_387/Y INVX1_LOC_94/Y 0.02fF
C23416 INVX1_LOC_546/A INVX1_LOC_92/A 0.01fF
C23417 NAND2X1_LOC_666/Y INVX1_LOC_674/A 0.03fF
C23418 INVX1_LOC_17/Y INVX1_LOC_26/Y 0.27fF
C23419 INVX1_LOC_583/A INVX1_LOC_62/Y 0.17fF
C23420 INVX1_LOC_95/A NAND2X1_LOC_333/B 0.03fF
C23421 INVX1_LOC_54/Y INVX1_LOC_15/Y 0.04fF
C23422 INVX1_LOC_89/Y INVX1_LOC_47/Y 0.15fF
C23423 INVX1_LOC_63/Y INVX1_LOC_374/Y 0.69fF
C23424 INVX1_LOC_502/A NAND2X1_LOC_275/Y 0.07fF
C23425 INVX1_LOC_551/A INVX1_LOC_32/Y -0.00fF
C23426 INVX1_LOC_158/Y INVX1_LOC_79/A 0.01fF
C23427 INVX1_LOC_93/Y INVX1_LOC_507/Y 0.18fF
C23428 INVX1_LOC_79/A INVX1_LOC_509/A 0.08fF
C23429 INVX1_LOC_6/Y NAND2X1_LOC_240/A 0.01fF
C23430 INVX1_LOC_328/Y INVX1_LOC_169/Y 0.37fF
C23431 INVX1_LOC_138/Y INVX1_LOC_655/A 0.04fF
C23432 INVX1_LOC_105/A INVX1_LOC_100/Y 0.02fF
C23433 INVX1_LOC_519/A INVX1_LOC_363/A 0.00fF
C23434 INVX1_LOC_520/Y INVX1_LOC_58/Y 0.05fF
C23435 INVX1_LOC_47/Y INVX1_LOC_501/A 0.08fF
C23436 NAND2X1_LOC_689/B INVX1_LOC_245/A 0.04fF
C23437 INVX1_LOC_360/Y INVX1_LOC_74/Y 1.10fF
C23438 NAND2X1_LOC_250/Y NAND2X1_LOC_843/B 0.01fF
C23439 NAND2X1_LOC_488/Y INVX1_LOC_48/Y 0.04fF
C23440 INVX1_LOC_199/Y INVX1_LOC_9/Y 0.31fF
C23441 INVX1_LOC_665/Y NAND2X1_LOC_372/Y 0.03fF
C23442 INVX1_LOC_89/Y INVX1_LOC_119/Y 0.18fF
C23443 INVX1_LOC_164/Y INVX1_LOC_588/A 0.11fF
C23444 INVX1_LOC_346/A INVX1_LOC_79/A 0.04fF
C23445 INVX1_LOC_32/Y INVX1_LOC_75/Y 0.07fF
C23446 INVX1_LOC_276/Y INVX1_LOC_655/A 0.04fF
C23447 INVX1_LOC_501/A INVX1_LOC_119/Y 0.07fF
C23448 INVX1_LOC_63/Y INVX1_LOC_319/A 0.01fF
C23449 INVX1_LOC_3/Y VDD 0.73fF
C23450 INVX1_LOC_85/A INVX1_LOC_9/Y 0.05fF
C23451 INVX1_LOC_62/Y INVX1_LOC_199/Y 0.04fF
C23452 VDD INVX1_LOC_191/Y 0.23fF
C23453 INVX1_LOC_69/Y INVX1_LOC_211/A 0.10fF
C23454 INVX1_LOC_63/Y NAND2X1_LOC_843/B 0.05fF
C23455 INVX1_LOC_69/Y INVX1_LOC_64/Y 0.26fF
C23456 INVX1_LOC_224/Y INVX1_LOC_158/A 0.03fF
C23457 INVX1_LOC_63/Y INVX1_LOC_625/Y 2.46fF
C23458 INVX1_LOC_682/Y INVX1_LOC_364/A 0.19fF
C23459 INPUT_0 NAND2X1_LOC_537/B 0.01fF
C23460 VDD INVX1_LOC_180/A -0.00fF
C23461 INVX1_LOC_224/Y INVX1_LOC_250/A 0.01fF
C23462 INVX1_LOC_206/Y INVX1_LOC_530/Y 0.15fF
C23463 INVX1_LOC_412/Y INVX1_LOC_134/A 0.02fF
C23464 INVX1_LOC_603/Y INVX1_LOC_615/A 0.13fF
C23465 VDD INVX1_LOC_610/Y 0.21fF
C23466 INPUT_0 INVX1_LOC_586/A 0.60fF
C23467 INVX1_LOC_224/Y INVX1_LOC_76/Y 0.03fF
C23468 INVX1_LOC_206/Y NAND2X1_LOC_318/A 0.67fF
C23469 VDD INVX1_LOC_511/A 0.17fF
C23470 NAND2X1_LOC_503/B INVX1_LOC_21/Y 0.08fF
C23471 NAND2X1_LOC_516/Y INVX1_LOC_586/A 0.03fF
C23472 INVX1_LOC_560/Y INVX1_LOC_80/A 0.03fF
C23473 INVX1_LOC_578/A INVX1_LOC_76/Y 0.07fF
C23474 VDD INVX1_LOC_509/Y 0.21fF
C23475 INVX1_LOC_174/Y INVX1_LOC_85/Y 0.00fF
C23476 VDD INVX1_LOC_417/Y 0.83fF
C23477 INVX1_LOC_442/A NAND2X1_LOC_332/B 0.02fF
C23478 VDD NAND2X1_LOC_679/B 0.01fF
C23479 VDD INVX1_LOC_491/Y 0.21fF
C23480 INVX1_LOC_596/A INVX1_LOC_215/Y 0.01fF
C23481 INVX1_LOC_198/A NAND2X1_LOC_86/a_36_24# 0.00fF
C23482 VDD INVX1_LOC_398/Y 0.21fF
C23483 INVX1_LOC_563/A INVX1_LOC_206/Y 0.01fF
C23484 NAND2X1_LOC_7/Y NAND2X1_LOC_615/B 0.01fF
C23485 INVX1_LOC_381/A INVX1_LOC_45/Y 0.08fF
C23486 INVX1_LOC_266/A NAND2X1_LOC_544/a_36_24# 0.00fF
C23487 NAND2X1_LOC_537/A INVX1_LOC_35/Y 0.19fF
C23488 VDD INVX1_LOC_59/Y 1.08fF
C23489 INVX1_LOC_586/Y INVX1_LOC_586/A 0.02fF
C23490 INVX1_LOC_11/Y INVX1_LOC_560/Y 0.03fF
C23491 NAND2X1_LOC_543/B INVX1_LOC_54/Y 0.05fF
C23492 INVX1_LOC_224/Y INVX1_LOC_559/A 0.01fF
C23493 VDD INVX1_LOC_48/Y 2.23fF
C23494 INVX1_LOC_619/A INVX1_LOC_207/A 0.05fF
C23495 INVX1_LOC_206/Y INVX1_LOC_202/Y 0.08fF
C23496 INVX1_LOC_526/A INVX1_LOC_111/A 0.02fF
C23497 NAND2X1_LOC_355/A NAND2X1_LOC_801/A 0.03fF
C23498 INVX1_LOC_228/Y INVX1_LOC_59/Y 0.03fF
C23499 INVX1_LOC_17/Y INVX1_LOC_560/A 0.07fF
C23500 NAND2X1_LOC_513/Y NAND2X1_LOC_413/Y 0.07fF
C23501 INPUT_3 INVX1_LOC_381/A 0.07fF
C23502 NAND2X1_LOC_331/A INVX1_LOC_335/A 0.04fF
C23503 INVX1_LOC_629/Y INVX1_LOC_259/Y 0.01fF
C23504 INVX1_LOC_35/Y INVX1_LOC_216/Y 0.01fF
C23505 INVX1_LOC_31/A INVX1_LOC_29/Y 0.04fF
C23506 INVX1_LOC_21/Y INVX1_LOC_273/A 0.07fF
C23507 NAND2X1_LOC_76/a_36_24# INVX1_LOC_98/Y 0.00fF
C23508 NAND2X1_LOC_93/Y INVX1_LOC_525/Y 0.06fF
C23509 INVX1_LOC_228/Y INVX1_LOC_48/Y 0.00fF
C23510 INVX1_LOC_347/Y INVX1_LOC_638/A 0.44fF
C23511 INVX1_LOC_410/Y INPUT_1 0.07fF
C23512 INVX1_LOC_213/Y INVX1_LOC_547/Y 0.08fF
C23513 NAND2X1_LOC_475/A INVX1_LOC_89/Y 0.13fF
C23514 INVX1_LOC_375/A INPUT_1 0.02fF
C23515 INVX1_LOC_468/Y INVX1_LOC_76/Y 0.03fF
C23516 INVX1_LOC_544/A NAND2X1_LOC_332/B 0.17fF
C23517 NAND2X1_LOC_332/B INVX1_LOC_116/Y 0.04fF
C23518 INVX1_LOC_401/Y NAND2X1_LOC_513/A 0.05fF
C23519 INVX1_LOC_210/Y INVX1_LOC_366/A -0.02fF
C23520 VDD NAND2X1_LOC_491/Y 0.00fF
C23521 NAND2X1_LOC_370/A NAND2X1_LOC_267/A -0.00fF
C23522 NAND2X1_LOC_475/A INVX1_LOC_154/A 0.02fF
C23523 GATE_741 INVX1_LOC_137/Y 0.02fF
C23524 INVX1_LOC_45/Y NAND2X1_LOC_720/A 0.00fF
C23525 INVX1_LOC_257/Y INVX1_LOC_69/Y 0.12fF
C23526 INVX1_LOC_51/Y INVX1_LOC_360/A 0.07fF
C23527 NAND2X1_LOC_56/Y NAND2X1_LOC_197/a_36_24# 0.00fF
C23528 NAND2X1_LOC_13/Y INVX1_LOC_35/Y 0.03fF
C23529 INVX1_LOC_51/Y INVX1_LOC_118/A 0.02fF
C23530 NAND2X1_LOC_589/a_36_24# INVX1_LOC_31/Y 0.00fF
C23531 INVX1_LOC_686/A INVX1_LOC_115/A 0.02fF
C23532 INVX1_LOC_25/Y INVX1_LOC_334/Y 0.02fF
C23533 INVX1_LOC_435/Y INVX1_LOC_671/Y 0.04fF
C23534 INVX1_LOC_206/Y INVX1_LOC_49/Y 0.35fF
C23535 INVX1_LOC_11/Y NAND2X1_LOC_620/a_36_24# 0.00fF
C23536 INVX1_LOC_596/A INVX1_LOC_321/Y 0.00fF
C23537 INVX1_LOC_180/A NAND2X1_LOC_243/A 0.02fF
C23538 INVX1_LOC_607/Y INVX1_LOC_312/Y 0.09fF
C23539 VDD NAND2X1_LOC_434/B 0.03fF
C23540 INVX1_LOC_298/A INVX1_LOC_586/A 0.05fF
C23541 NAND2X1_LOC_475/A INVX1_LOC_501/A 0.10fF
C23542 INVX1_LOC_586/A INVX1_LOC_498/A 0.00fF
C23543 INVX1_LOC_428/A NAND2X1_LOC_486/A 0.36fF
C23544 INVX1_LOC_446/Y INVX1_LOC_69/Y 0.01fF
C23545 INVX1_LOC_20/Y NAND2X1_LOC_615/B 0.03fF
C23546 INVX1_LOC_11/Y INVX1_LOC_84/A 8.69fF
C23547 INVX1_LOC_17/Y INVX1_LOC_369/A 0.10fF
C23548 INVX1_LOC_21/Y NAND2X1_LOC_393/Y 0.08fF
C23549 INVX1_LOC_321/A INVX1_LOC_431/Y 0.01fF
C23550 INVX1_LOC_395/A INVX1_LOC_507/Y 0.42fF
C23551 NAND2X1_LOC_685/B INVX1_LOC_496/Y 0.16fF
C23552 INVX1_LOC_617/Y INVX1_LOC_50/Y 0.29fF
C23553 INVX1_LOC_554/Y INVX1_LOC_662/A 0.03fF
C23554 INVX1_LOC_558/A NAND2X1_LOC_542/A 0.21fF
C23555 VDD INVX1_LOC_472/Y 0.21fF
C23556 INVX1_LOC_20/Y INVX1_LOC_127/Y 0.01fF
C23557 INVX1_LOC_93/Y INVX1_LOC_522/Y 0.09fF
C23558 INVX1_LOC_449/A INVX1_LOC_665/Y 0.02fF
C23559 INVX1_LOC_384/A INVX1_LOC_69/Y 0.07fF
C23560 INVX1_LOC_117/Y INVX1_LOC_197/A 0.01fF
C23561 INVX1_LOC_20/Y INVX1_LOC_66/A 0.07fF
C23562 INVX1_LOC_134/Y INVX1_LOC_345/A 0.04fF
C23563 INVX1_LOC_442/Y INVX1_LOC_370/A 0.01fF
C23564 NAND2X1_LOC_115/a_36_24# INVX1_LOC_367/A 0.00fF
C23565 INVX1_LOC_455/A INVX1_LOC_316/Y 0.44fF
C23566 INVX1_LOC_20/Y INVX1_LOC_296/A 0.00fF
C23567 INVX1_LOC_361/Y INVX1_LOC_670/Y 0.00fF
C23568 INVX1_LOC_49/Y INVX1_LOC_242/A 0.02fF
C23569 INVX1_LOC_99/Y INVX1_LOC_194/Y 0.04fF
C23570 INVX1_LOC_681/A INVX1_LOC_304/Y 0.00fF
C23571 INVX1_LOC_442/A INVX1_LOC_242/Y 0.19fF
C23572 INVX1_LOC_117/Y INVX1_LOC_124/Y 0.04fF
C23573 NAND2X1_LOC_97/B NAND2X1_LOC_388/A 0.26fF
C23574 INVX1_LOC_686/A INVX1_LOC_49/Y 0.07fF
C23575 NAND2X1_LOC_697/Y INVX1_LOC_186/Y 0.02fF
C23576 INVX1_LOC_158/Y INVX1_LOC_48/Y 0.01fF
C23577 INVX1_LOC_93/Y NAND2X1_LOC_448/A 0.00fF
C23578 INVX1_LOC_45/Y INVX1_LOC_100/Y 0.29fF
C23579 INVX1_LOC_417/A NAND2X1_LOC_388/A 0.01fF
C23580 NAND2X1_LOC_781/B INVX1_LOC_611/A 0.05fF
C23581 NAND2X1_LOC_147/B INVX1_LOC_239/A 0.09fF
C23582 INVX1_LOC_543/Y INVX1_LOC_178/A 0.71fF
C23583 INVX1_LOC_469/Y INVX1_LOC_360/Y 0.01fF
C23584 INVX1_LOC_72/Y INVX1_LOC_41/Y 0.00fF
C23585 INVX1_LOC_410/A INVX1_LOC_600/A 0.04fF
C23586 INVX1_LOC_155/Y INVX1_LOC_187/Y 0.01fF
C23587 INVX1_LOC_682/A INVX1_LOC_486/Y 0.09fF
C23588 INVX1_LOC_588/Y INVX1_LOC_513/A -0.00fF
C23589 INVX1_LOC_31/Y INVX1_LOC_350/A 0.06fF
C23590 NAND2X1_LOC_88/B INVX1_LOC_179/A 0.03fF
C23591 INVX1_LOC_53/Y INVX1_LOC_285/Y 0.00fF
C23592 INVX1_LOC_53/Y INVX1_LOC_9/Y 0.22fF
C23593 INVX1_LOC_45/Y INVX1_LOC_74/Y 0.96fF
C23594 INVX1_LOC_301/Y INVX1_LOC_519/A 0.04fF
C23595 INVX1_LOC_103/Y INVX1_LOC_48/Y 0.09fF
C23596 INVX1_LOC_69/Y INVX1_LOC_145/Y 0.96fF
C23597 INVX1_LOC_300/A INVX1_LOC_296/A 0.00fF
C23598 INVX1_LOC_502/A INVX1_LOC_235/Y 0.02fF
C23599 INVX1_LOC_210/Y INVX1_LOC_6/Y 0.01fF
C23600 INVX1_LOC_561/A INVX1_LOC_259/Y 0.00fF
C23601 INPUT_3 INVX1_LOC_100/Y 0.24fF
C23602 INVX1_LOC_356/A INVX1_LOC_41/Y 0.04fF
C23603 INVX1_LOC_45/Y INVX1_LOC_483/Y 0.00fF
C23604 INVX1_LOC_47/Y INVX1_LOC_194/Y 0.05fF
C23605 INVX1_LOC_586/A INVX1_LOC_211/A 0.07fF
C23606 INVX1_LOC_35/Y NAND2X1_LOC_668/Y 0.04fF
C23607 INVX1_LOC_35/Y INVX1_LOC_361/A 0.07fF
C23608 INVX1_LOC_575/A NAND2X1_LOC_846/B 0.01fF
C23609 NAND2X1_LOC_837/A NAND2X1_LOC_720/A 0.10fF
C23610 INVX1_LOC_507/Y INVX1_LOC_189/Y 0.02fF
C23611 INVX1_LOC_361/Y INVX1_LOC_253/Y 0.14fF
C23612 NAND2X1_LOC_144/a_36_24# INVX1_LOC_662/A 0.00fF
C23613 GATE_865 NAND2X1_LOC_809/a_36_24# 0.00fF
C23614 INVX1_LOC_619/A INVX1_LOC_79/A 0.18fF
C23615 INVX1_LOC_17/Y NAND2X1_LOC_605/B 0.00fF
C23616 INVX1_LOC_316/Y NAND2X1_LOC_823/Y 0.19fF
C23617 INVX1_LOC_116/Y INVX1_LOC_242/Y 0.07fF
C23618 INVX1_LOC_41/Y INVX1_LOC_519/A 0.03fF
C23619 INVX1_LOC_134/Y INVX1_LOC_280/A 0.00fF
C23620 INVX1_LOC_361/Y INVX1_LOC_63/Y 0.03fF
C23621 INVX1_LOC_53/Y INVX1_LOC_62/Y 0.15fF
C23622 INVX1_LOC_63/Y NAND2X1_LOC_333/B 0.08fF
C23623 NAND2X1_LOC_542/A INVX1_LOC_46/Y 0.00fF
C23624 INVX1_LOC_134/Y NAND2X1_LOC_372/Y 0.07fF
C23625 NAND2X1_LOC_274/B INVX1_LOC_98/Y 0.05fF
C23626 NAND2X1_LOC_286/A INVX1_LOC_240/A 0.12fF
C23627 INVX1_LOC_42/Y INVX1_LOC_85/A 0.01fF
C23628 INVX1_LOC_100/Y NAND2X1_LOC_69/Y 0.02fF
C23629 INVX1_LOC_17/Y NAND2X1_LOC_626/Y -0.03fF
C23630 INVX1_LOC_6/Y NAND2X1_LOC_344/B 0.01fF
C23631 NAND2X1_LOC_331/Y INVX1_LOC_74/Y 0.12fF
C23632 INVX1_LOC_272/Y INVX1_LOC_622/Y 0.02fF
C23633 NAND2X1_LOC_786/B INVX1_LOC_48/Y 0.01fF
C23634 INVX1_LOC_26/Y INVX1_LOC_198/A 0.10fF
C23635 INVX1_LOC_130/Y INVX1_LOC_75/Y 0.07fF
C23636 INVX1_LOC_376/Y INVX1_LOC_46/Y 0.07fF
C23637 NAND2X1_LOC_786/B NAND2X1_LOC_60/a_36_24# 0.00fF
C23638 INVX1_LOC_47/Y INVX1_LOC_44/Y 0.05fF
C23639 INVX1_LOC_49/Y NAND2X1_LOC_334/A 11.54fF
C23640 INVX1_LOC_258/Y INVX1_LOC_63/Y 0.01fF
C23641 INVX1_LOC_26/Y NAND2X1_LOC_770/a_36_24# 0.00fF
C23642 INVX1_LOC_59/Y INVX1_LOC_635/Y 0.44fF
C23643 NAND2X1_LOC_603/Y INVX1_LOC_634/Y 0.01fF
C23644 INVX1_LOC_50/Y NAND2X1_LOC_268/a_36_24# 0.00fF
C23645 INVX1_LOC_224/Y INVX1_LOC_192/A 0.04fF
C23646 INVX1_LOC_292/Y INVX1_LOC_273/Y 0.00fF
C23647 INVX1_LOC_211/A NAND2X1_LOC_74/a_36_24# 0.00fF
C23648 INVX1_LOC_202/A VDD -0.00fF
C23649 NAND2X1_LOC_428/a_36_24# INVX1_LOC_505/A 0.00fF
C23650 NAND2X1_LOC_106/Y INVX1_LOC_479/A 0.02fF
C23651 INVX1_LOC_41/Y INVX1_LOC_659/A 0.07fF
C23652 INVX1_LOC_582/A INVX1_LOC_62/Y 0.10fF
C23653 INVX1_LOC_446/A INVX1_LOC_393/Y 0.07fF
C23654 INPUT_0 INVX1_LOC_567/A 0.01fF
C23655 INVX1_LOC_148/Y INVX1_LOC_338/Y 0.12fF
C23656 NAND2X1_LOC_844/A NAND2X1_LOC_274/Y 0.00fF
C23657 INVX1_LOC_254/Y INVX1_LOC_92/A 0.01fF
C23658 INVX1_LOC_58/Y INVX1_LOC_483/A 0.01fF
C23659 INVX1_LOC_203/Y NAND2X1_LOC_475/A 0.00fF
C23660 INVX1_LOC_97/A INVX1_LOC_616/Y 0.01fF
C23661 VDD INVX1_LOC_561/Y 0.47fF
C23662 NAND2X1_LOC_848/a_36_24# INVX1_LOC_655/A 0.01fF
C23663 NAND2X1_LOC_301/B INVX1_LOC_652/A 0.00fF
C23664 INVX1_LOC_206/Y INVX1_LOC_158/A 0.01fF
C23665 NAND2X1_LOC_45/Y INVX1_LOC_118/Y 0.06fF
C23666 VDD NAND2X1_LOC_513/Y 0.00fF
C23667 INVX1_LOC_301/A INVX1_LOC_442/A 0.31fF
C23668 INVX1_LOC_471/Y INVX1_LOC_588/A 0.06fF
C23669 NAND2X1_LOC_790/B INVX1_LOC_286/Y 0.02fF
C23670 INPUT_0 INVX1_LOC_140/Y 0.01fF
C23671 NAND2X1_LOC_123/B INVX1_LOC_479/A 0.07fF
C23672 NAND2X1_LOC_843/B INVX1_LOC_669/A 0.26fF
C23673 NAND2X1_LOC_242/A INVX1_LOC_45/Y 0.01fF
C23674 INPUT_0 INVX1_LOC_366/A 0.02fF
C23675 INVX1_LOC_206/Y INVX1_LOC_76/Y 0.50fF
C23676 INPUT_0 NAND2X1_LOC_426/Y 0.01fF
C23677 INVX1_LOC_479/A NAND2X1_LOC_428/Y 0.03fF
C23678 INVX1_LOC_446/Y INVX1_LOC_586/A 0.31fF
C23679 INVX1_LOC_425/A INVX1_LOC_400/Y 0.07fF
C23680 INVX1_LOC_575/A INVX1_LOC_554/A 0.06fF
C23681 INVX1_LOC_395/A INVX1_LOC_522/Y 1.24fF
C23682 INVX1_LOC_420/Y NAND2X1_LOC_541/B 0.02fF
C23683 INVX1_LOC_397/A NAND2X1_LOC_318/A 0.58fF
C23684 INPUT_0 INVX1_LOC_486/Y 0.01fF
C23685 INVX1_LOC_319/Y INVX1_LOC_84/A 0.03fF
C23686 NAND2X1_LOC_34/a_36_24# INVX1_LOC_54/Y 0.00fF
C23687 INVX1_LOC_98/A INVX1_LOC_396/Y 0.04fF
C23688 INVX1_LOC_301/A INVX1_LOC_116/Y 1.19fF
C23689 INVX1_LOC_20/Y INVX1_LOC_442/A 0.17fF
C23690 INVX1_LOC_384/A INVX1_LOC_586/A 0.07fF
C23691 INVX1_LOC_17/Y NAND2X1_LOC_385/a_36_24# 0.00fF
C23692 INVX1_LOC_479/A INVX1_LOC_92/A 0.23fF
C23693 INVX1_LOC_409/Y INVX1_LOC_54/Y 0.19fF
C23694 INVX1_LOC_118/Y INVX1_LOC_99/Y 0.02fF
C23695 NAND2X1_LOC_537/B INVX1_LOC_145/Y 0.04fF
C23696 VDD INVX1_LOC_396/A -0.00fF
C23697 INVX1_LOC_76/Y INVX1_LOC_686/A 0.07fF
C23698 INVX1_LOC_17/Y INVX1_LOC_103/A 0.04fF
C23699 NAND2X1_LOC_475/A INVX1_LOC_194/Y 0.00fF
C23700 INVX1_LOC_390/A NAND2X1_LOC_216/a_36_24# 0.00fF
C23701 INVX1_LOC_312/Y INVX1_LOC_384/A 0.07fF
C23702 INVX1_LOC_619/A INVX1_LOC_180/A 0.03fF
C23703 INVX1_LOC_269/Y INVX1_LOC_160/A 0.00fF
C23704 INVX1_LOC_293/Y INVX1_LOC_381/A 0.01fF
C23705 INVX1_LOC_570/A NAND2X1_LOC_418/Y 0.19fF
C23706 INVX1_LOC_21/Y INVX1_LOC_72/Y 0.02fF
C23707 NAND2X1_LOC_543/B INVX1_LOC_89/Y 1.80fF
C23708 VDD INVX1_LOC_559/Y 0.21fF
C23709 INVX1_LOC_586/A INVX1_LOC_677/A 0.01fF
C23710 INVX1_LOC_96/Y INVX1_LOC_99/Y 0.01fF
C23711 INVX1_LOC_152/Y INVX1_LOC_496/Y 0.01fF
C23712 NAND2X1_LOC_79/B INVX1_LOC_80/A 0.01fF
C23713 INVX1_LOC_553/Y INVX1_LOC_50/Y 0.16fF
C23714 NAND2X1_LOC_322/Y INVX1_LOC_257/A 0.27fF
C23715 INVX1_LOC_410/Y INVX1_LOC_50/Y 0.03fF
C23716 INVX1_LOC_224/Y INVX1_LOC_32/Y 0.11fF
C23717 INVX1_LOC_301/A INVX1_LOC_255/A 0.03fF
C23718 INVX1_LOC_3/Y INVX1_LOC_145/A 0.02fF
C23719 INVX1_LOC_586/A INVX1_LOC_145/Y 3.45fF
C23720 INVX1_LOC_395/A INVX1_LOC_295/Y 0.01fF
C23721 INVX1_LOC_76/Y INVX1_LOC_14/A 0.03fF
C23722 GATE_579 INVX1_LOC_17/Y 0.06fF
C23723 INVX1_LOC_375/A INVX1_LOC_50/Y 0.03fF
C23724 INVX1_LOC_202/Y INVX1_LOC_94/A 0.03fF
C23725 INVX1_LOC_243/A INPUT_3 0.01fF
C23726 INVX1_LOC_435/A NAND2X1_LOC_613/Y 0.01fF
C23727 INVX1_LOC_578/A INVX1_LOC_32/Y 0.07fF
C23728 INVX1_LOC_367/A NAND2X1_LOC_496/Y 0.01fF
C23729 INPUT_0 INVX1_LOC_6/Y 3.03fF
C23730 INVX1_LOC_20/Y INVX1_LOC_544/A 0.03fF
C23731 INVX1_LOC_448/A INVX1_LOC_312/Y 0.07fF
C23732 INVX1_LOC_118/Y INVX1_LOC_47/Y 0.01fF
C23733 INVX1_LOC_20/Y INVX1_LOC_116/Y 0.03fF
C23734 NAND2X1_LOC_503/B INVX1_LOC_26/Y 0.71fF
C23735 VDD NAND2X1_LOC_615/Y 0.26fF
C23736 NAND2X1_LOC_538/B INVX1_LOC_98/Y 0.13fF
C23737 NAND2X1_LOC_271/B NAND2X1_LOC_520/A 0.02fF
C23738 INVX1_LOC_596/A INVX1_LOC_683/A 0.00fF
C23739 INVX1_LOC_17/Y INVX1_LOC_235/Y 0.13fF
C23740 INVX1_LOC_432/Y INVX1_LOC_84/A 0.06fF
C23741 INVX1_LOC_444/Y INVX1_LOC_325/Y 0.03fF
C23742 NAND2X1_LOC_331/B INVX1_LOC_69/Y 0.01fF
C23743 INVX1_LOC_68/Y NAND2X1_LOC_614/a_36_24# 0.00fF
C23744 INVX1_LOC_469/Y INVX1_LOC_45/Y 0.03fF
C23745 INVX1_LOC_522/Y INVX1_LOC_189/Y 0.02fF
C23746 INVX1_LOC_555/A INVX1_LOC_523/A 0.05fF
C23747 INVX1_LOC_312/Y INVX1_LOC_145/Y 3.57fF
C23748 INVX1_LOC_603/Y NAND2X1_LOC_237/Y 0.03fF
C23749 NAND2X1_LOC_516/Y INVX1_LOC_6/Y 0.03fF
C23750 NAND2X1_LOC_781/A INVX1_LOC_145/Y 0.01fF
C23751 INVX1_LOC_607/Y NAND2X1_LOC_820/A 0.04fF
C23752 NAND2X1_LOC_188/a_36_24# INVX1_LOC_31/Y 0.00fF
C23753 INVX1_LOC_587/A INVX1_LOC_298/A 0.03fF
C23754 INVX1_LOC_395/A INVX1_LOC_508/A 0.04fF
C23755 NAND2X1_LOC_152/B INVX1_LOC_35/Y 0.01fF
C23756 NAND2X1_LOC_107/Y NAND2X1_LOC_113/a_36_24# 0.00fF
C23757 INVX1_LOC_547/Y NAND2X1_LOC_258/Y 0.51fF
C23758 NAND2X1_LOC_181/A INVX1_LOC_45/Y 0.03fF
C23759 NAND2X1_LOC_644/a_36_24# INVX1_LOC_50/Y 0.00fF
C23760 INVX1_LOC_374/A INVX1_LOC_258/Y 0.01fF
C23761 INVX1_LOC_268/A INVX1_LOC_300/A 0.03fF
C23762 INVX1_LOC_233/Y NAND2X1_LOC_292/Y 0.12fF
C23763 NAND2X1_LOC_24/Y NAND2X1_LOC_84/B 0.01fF
C23764 NAND2X1_LOC_545/B INVX1_LOC_159/Y 0.03fF
C23765 INVX1_LOC_549/A INVX1_LOC_491/A 0.77fF
C23766 INVX1_LOC_193/A INVX1_LOC_80/A 0.01fF
C23767 INVX1_LOC_116/Y NAND2X1_LOC_605/a_36_24# 0.00fF
C23768 INVX1_LOC_272/Y INVX1_LOC_298/A 0.00fF
C23769 INVX1_LOC_211/Y INVX1_LOC_296/Y 0.01fF
C23770 VDD INVX1_LOC_614/Y 0.24fF
C23771 INVX1_LOC_117/Y INVX1_LOC_336/Y 0.03fF
C23772 NAND2X1_LOC_706/B INVX1_LOC_367/A 0.25fF
C23773 NAND2X1_LOC_332/B INVX1_LOC_69/Y 0.50fF
C23774 INPUT_2 INVX1_LOC_84/Y 0.15fF
C23775 INVX1_LOC_586/Y INVX1_LOC_6/Y 0.02fF
C23776 INVX1_LOC_366/A NAND2X1_LOC_215/a_36_24# 0.01fF
C23777 INVX1_LOC_576/Y INVX1_LOC_50/Y 0.01fF
C23778 INVX1_LOC_392/A NAND2X1_LOC_525/a_36_24# 0.00fF
C23779 INVX1_LOC_435/Y NAND2X1_LOC_274/B 0.03fF
C23780 INVX1_LOC_444/Y NAND2X1_LOC_548/a_36_24# 0.01fF
C23781 INVX1_LOC_54/Y INVX1_LOC_600/A 0.21fF
C23782 NAND2X1_LOC_551/a_36_24# INVX1_LOC_99/A 0.00fF
C23783 NAND2X1_LOC_387/Y NAND2X1_LOC_237/Y 0.02fF
C23784 INVX1_LOC_159/Y INVX1_LOC_98/Y 0.10fF
C23785 NAND2X1_LOC_383/Y INVX1_LOC_9/Y 0.07fF
C23786 INVX1_LOC_555/Y INVX1_LOC_9/Y 0.01fF
C23787 NAND2X1_LOC_391/A INVX1_LOC_47/Y 0.27fF
C23788 NAND2X1_LOC_122/Y INVX1_LOC_26/Y 0.03fF
C23789 NAND2X1_LOC_179/Y INVX1_LOC_117/Y 0.01fF
C23790 INVX1_LOC_80/A NAND2X1_LOC_285/a_36_24# 0.00fF
C23791 INVX1_LOC_560/Y INVX1_LOC_625/Y 0.05fF
C23792 INVX1_LOC_273/A INVX1_LOC_26/Y 1.22fF
C23793 NAND2X1_LOC_207/a_36_24# INVX1_LOC_63/Y 0.00fF
C23794 INVX1_LOC_45/Y INVX1_LOC_79/A 0.20fF
C23795 INVX1_LOC_410/A NAND2X1_LOC_56/Y 0.04fF
C23796 INVX1_LOC_137/A INVX1_LOC_475/Y 0.01fF
C23797 INVX1_LOC_197/A INVX1_LOC_58/Y 0.01fF
C23798 INVX1_LOC_347/Y INVX1_LOC_134/Y 0.12fF
C23799 INVX1_LOC_45/Y NAND2X1_LOC_631/B 0.01fF
C23800 NAND2X1_LOC_308/A INVX1_LOC_352/A 0.10fF
C23801 INVX1_LOC_173/Y INVX1_LOC_178/A 0.00fF
C23802 INVX1_LOC_607/Y INVX1_LOC_6/Y 0.16fF
C23803 INVX1_LOC_47/Y NAND2X1_LOC_418/Y 0.02fF
C23804 INVX1_LOC_254/Y INPUT_1 0.00fF
C23805 INVX1_LOC_63/Y INVX1_LOC_307/A 0.01fF
C23806 INVX1_LOC_45/Y NAND2X1_LOC_396/Y 0.03fF
C23807 INVX1_LOC_335/Y INVX1_LOC_659/A 0.07fF
C23808 INVX1_LOC_674/A INVX1_LOC_50/Y 0.07fF
C23809 INVX1_LOC_93/Y NAND2X1_LOC_775/B 1.09fF
C23810 NAND2X1_LOC_97/A INVX1_LOC_41/Y 0.01fF
C23811 INVX1_LOC_348/A INVX1_LOC_79/A 0.05fF
C23812 INVX1_LOC_92/Y INVX1_LOC_94/A 0.02fF
C23813 INVX1_LOC_596/A NAND2X1_LOC_274/B 0.03fF
C23814 INPUT_3 INVX1_LOC_79/A 0.03fF
C23815 NAND2X1_LOC_48/Y INVX1_LOC_328/Y 0.00fF
C23816 INVX1_LOC_93/Y NAND2X1_LOC_706/B 0.07fF
C23817 INVX1_LOC_293/Y INVX1_LOC_100/Y 0.01fF
C23818 INVX1_LOC_76/Y NAND2X1_LOC_609/B 0.20fF
C23819 INVX1_LOC_556/Y NAND2X1_LOC_307/B 0.04fF
C23820 NAND2X1_LOC_859/a_36_24# INVX1_LOC_6/Y 0.00fF
C23821 INVX1_LOC_11/Y NAND2X1_LOC_532/Y 0.01fF
C23822 INVX1_LOC_442/Y INVX1_LOC_63/Y 0.09fF
C23823 INVX1_LOC_84/A INVX1_LOC_319/A 0.01fF
C23824 INVX1_LOC_32/Y INVX1_LOC_227/Y 0.01fF
C23825 NAND2X1_LOC_285/B INVX1_LOC_58/Y 0.01fF
C23826 INVX1_LOC_80/A INVX1_LOC_106/Y 0.01fF
C23827 NAND2X1_LOC_707/A INVX1_LOC_588/A 0.00fF
C23828 INVX1_LOC_43/A INVX1_LOC_87/A 0.04fF
C23829 INVX1_LOC_117/Y NAND2X1_LOC_128/A 0.83fF
C23830 INVX1_LOC_166/A INVX1_LOC_670/A 0.04fF
C23831 INVX1_LOC_372/Y NAND2X1_LOC_123/B 0.32fF
C23832 NAND2X1_LOC_355/A INVX1_LOC_259/Y 0.02fF
C23833 INVX1_LOC_261/Y INVX1_LOC_263/Y 0.15fF
C23834 INVX1_LOC_35/Y INVX1_LOC_480/A 0.01fF
C23835 INVX1_LOC_58/Y NAND2X1_LOC_106/B 0.05fF
C23836 INVX1_LOC_298/A INVX1_LOC_6/Y 0.03fF
C23837 INVX1_LOC_300/A NAND2X1_LOC_719/A 0.07fF
C23838 NAND2X1_LOC_326/a_36_24# NAND2X1_LOC_123/B 0.01fF
C23839 NAND2X1_LOC_106/Y INVX1_LOC_391/A 0.02fF
C23840 INVX1_LOC_119/Y NAND2X1_LOC_418/Y 0.01fF
C23841 INVX1_LOC_204/Y INVX1_LOC_18/Y 0.04fF
C23842 INVX1_LOC_508/Y INVX1_LOC_645/Y 0.15fF
C23843 INVX1_LOC_575/Y NAND2X1_LOC_846/B 0.07fF
C23844 INVX1_LOC_6/Y INVX1_LOC_476/Y 0.39fF
C23845 INVX1_LOC_173/Y INVX1_LOC_58/Y 0.02fF
C23846 NAND2X1_LOC_285/B NAND2X1_LOC_342/B 0.37fF
C23847 INVX1_LOC_54/Y NAND2X1_LOC_780/a_36_24# 0.00fF
C23848 INVX1_LOC_679/Y INVX1_LOC_479/A 0.05fF
C23849 NAND2X1_LOC_673/B INVX1_LOC_100/Y 0.24fF
C23850 INVX1_LOC_49/Y NAND2X1_LOC_542/A 0.07fF
C23851 NAND2X1_LOC_606/Y INVX1_LOC_473/Y 0.07fF
C23852 INVX1_LOC_213/Y INVX1_LOC_62/Y 0.04fF
C23853 INVX1_LOC_12/Y INVX1_LOC_485/A 0.01fF
C23854 INVX1_LOC_49/Y INVX1_LOC_376/Y 0.17fF
C23855 INVX1_LOC_385/Y INVX1_LOC_443/A 3.99fF
C23856 INVX1_LOC_154/A INVX1_LOC_353/A 0.19fF
C23857 INVX1_LOC_544/Y INVX1_LOC_9/Y 0.28fF
C23858 NAND2X1_LOC_528/Y INPUT_1 0.35fF
C23859 INVX1_LOC_69/Y INVX1_LOC_242/Y 0.21fF
C23860 INVX1_LOC_479/A INPUT_1 0.28fF
C23861 VDD NAND2X1_LOC_69/B 0.11fF
C23862 INVX1_LOC_35/Y INVX1_LOC_291/Y 0.02fF
C23863 INVX1_LOC_656/A INVX1_LOC_74/Y 0.04fF
C23864 INVX1_LOC_12/Y INVX1_LOC_92/A 0.43fF
C23865 NAND2X1_LOC_184/Y INVX1_LOC_75/Y 0.01fF
C23866 INVX1_LOC_261/Y INVX1_LOC_454/Y 0.00fF
C23867 INVX1_LOC_6/Y INVX1_LOC_211/A 0.05fF
C23868 INVX1_LOC_206/Y NAND2X1_LOC_193/a_36_24# 0.00fF
C23869 INVX1_LOC_662/A INVX1_LOC_62/Y 0.02fF
C23870 INVX1_LOC_653/A INVX1_LOC_166/Y 0.14fF
C23871 INVX1_LOC_166/A NAND2X1_LOC_418/a_36_24# 0.00fF
C23872 NAND2X1_LOC_373/Y INVX1_LOC_442/A 0.15fF
C23873 INVX1_LOC_203/A INVX1_LOC_90/Y 0.07fF
C23874 INVX1_LOC_490/Y NAND2X1_LOC_457/A 0.00fF
C23875 VDD INVX1_LOC_340/Y 0.46fF
C23876 INVX1_LOC_447/A INVX1_LOC_51/Y 0.53fF
C23877 INVX1_LOC_452/Y INVX1_LOC_434/A 0.01fF
C23878 INVX1_LOC_560/A NAND2X1_LOC_370/A 0.06fF
C23879 NAND2X1_LOC_596/Y INVX1_LOC_340/Y 0.02fF
C23880 VDD NAND2X1_LOC_710/A -0.00fF
C23881 NAND2X1_LOC_525/Y INVX1_LOC_413/Y 0.31fF
C23882 VDD INVX1_LOC_634/A -0.00fF
C23883 INVX1_LOC_665/Y INVX1_LOC_109/Y 0.03fF
C23884 VDD INVX1_LOC_508/Y 0.35fF
C23885 VDD NAND2X1_LOC_541/B 0.01fF
C23886 NAND2X1_LOC_242/A NAND2X1_LOC_756/Y 0.03fF
C23887 INVX1_LOC_33/A NAND2X1_LOC_25/a_36_24# 0.02fF
C23888 NAND2X1_LOC_45/Y INVX1_LOC_297/A 0.05fF
C23889 VDD INVX1_LOC_383/Y 0.03fF
C23890 INVX1_LOC_98/A INVX1_LOC_94/A 0.24fF
C23891 NAND2X1_LOC_317/A INVX1_LOC_134/Y 0.09fF
C23892 VDD INVX1_LOC_155/Y 0.41fF
C23893 NAND2X1_LOC_373/Y INVX1_LOC_116/Y 0.03fF
C23894 INVX1_LOC_76/Y INVX1_LOC_94/A 0.00fF
C23895 NAND2X1_LOC_331/A INVX1_LOC_53/Y 0.03fF
C23896 INVX1_LOC_75/Y NAND2X1_LOC_271/A 0.09fF
C23897 INPUT_0 INVX1_LOC_161/A 0.02fF
C23898 INVX1_LOC_165/Y INVX1_LOC_134/Y 0.02fF
C23899 NAND2X1_LOC_710/A INVX1_LOC_510/Y 0.02fF
C23900 INVX1_LOC_442/A NAND2X1_LOC_524/a_36_24# 0.00fF
C23901 INVX1_LOC_578/A INVX1_LOC_130/Y 0.02fF
C23902 INVX1_LOC_312/Y NAND2X1_LOC_332/B 0.03fF
C23903 NAND2X1_LOC_322/Y INVX1_LOC_89/Y 0.03fF
C23904 INVX1_LOC_206/Y INVX1_LOC_345/Y 0.02fF
C23905 NAND2X1_LOC_498/Y INVX1_LOC_252/Y 0.05fF
C23906 NAND2X1_LOC_525/a_36_24# INVX1_LOC_362/Y 0.01fF
C23907 INVX1_LOC_395/A NAND2X1_LOC_775/B 0.14fF
C23908 INVX1_LOC_570/A INVX1_LOC_252/Y 0.14fF
C23909 INVX1_LOC_398/Y INVX1_LOC_45/Y 0.01fF
C23910 NAND2X1_LOC_533/a_36_24# INVX1_LOC_47/Y 0.00fF
C23911 INVX1_LOC_301/A INVX1_LOC_69/Y 0.09fF
C23912 NAND2X1_LOC_261/Y INVX1_LOC_385/Y 0.03fF
C23913 INVX1_LOC_206/Y INVX1_LOC_32/Y 9.24fF
C23914 INVX1_LOC_45/Y INVX1_LOC_59/Y 0.03fF
C23915 NAND2X1_LOC_335/B INVX1_LOC_89/Y 0.02fF
C23916 INVX1_LOC_614/A INVX1_LOC_508/Y 0.03fF
C23917 INVX1_LOC_463/A NAND2X1_LOC_686/B 0.02fF
C23918 INVX1_LOC_366/A INVX1_LOC_145/Y 0.01fF
C23919 INVX1_LOC_133/Y INVX1_LOC_643/Y 0.01fF
C23920 VDD INVX1_LOC_149/Y 0.22fF
C23921 NAND2X1_LOC_45/a_36_24# INVX1_LOC_6/Y 0.00fF
C23922 INVX1_LOC_48/Y NAND2X1_LOC_506/B 0.06fF
C23923 INVX1_LOC_21/Y NAND2X1_LOC_39/Y 0.04fF
C23924 INVX1_LOC_185/Y INVX1_LOC_48/Y 0.01fF
C23925 INVX1_LOC_45/Y INVX1_LOC_48/Y 10.28fF
C23926 INVX1_LOC_245/A INVX1_LOC_458/Y 0.00fF
C23927 INVX1_LOC_121/Y INVX1_LOC_49/Y 0.03fF
C23928 INVX1_LOC_96/Y INVX1_LOC_153/A 0.02fF
C23929 INVX1_LOC_551/Y INVX1_LOC_35/Y 0.01fF
C23930 NAND2X1_LOC_791/A NAND2X1_LOC_791/B 0.04fF
C23931 INVX1_LOC_76/Y INVX1_LOC_432/A 0.02fF
C23932 INVX1_LOC_412/A INVX1_LOC_253/Y 0.01fF
C23933 INVX1_LOC_272/Y INVX1_LOC_145/Y 0.00fF
C23934 NAND2X1_LOC_28/a_36_24# INVX1_LOC_6/Y 0.00fF
C23935 NAND2X1_LOC_370/A NAND2X1_LOC_309/a_36_24# 0.02fF
C23936 INVX1_LOC_282/A NAND2X1_LOC_842/a_36_24# 0.00fF
C23937 INVX1_LOC_213/Y INVX1_LOC_547/A 0.02fF
C23938 INVX1_LOC_677/Y INVX1_LOC_259/Y 0.82fF
C23939 INVX1_LOC_68/Y NAND2X1_LOC_507/A 0.14fF
C23940 INVX1_LOC_145/Y INVX1_LOC_486/Y 0.35fF
C23941 INVX1_LOC_134/Y INVX1_LOC_352/A 0.03fF
C23942 NAND2X1_LOC_557/a_36_24# INVX1_LOC_169/A 0.00fF
C23943 NAND2X1_LOC_148/B INVX1_LOC_132/Y 0.03fF
C23944 INVX1_LOC_413/Y INVX1_LOC_406/A 0.03fF
C23945 NAND2X1_LOC_533/a_36_24# INVX1_LOC_119/Y 0.00fF
C23946 INVX1_LOC_575/A INVX1_LOC_53/Y 0.06fF
C23947 INVX1_LOC_312/Y INVX1_LOC_503/Y 0.05fF
C23948 NAND2X1_LOC_184/Y NAND2X1_LOC_486/B 0.04fF
C23949 INVX1_LOC_396/Y INVX1_LOC_32/Y 0.30fF
C23950 INVX1_LOC_96/Y INVX1_LOC_96/A 0.05fF
C23951 INVX1_LOC_203/Y INVX1_LOC_353/A 0.08fF
C23952 INPUT_0 NAND2X1_LOC_192/A 0.01fF
C23953 INVX1_LOC_53/Y NAND2X1_LOC_485/a_36_24# 0.01fF
C23954 INVX1_LOC_49/Y INVX1_LOC_253/A 0.01fF
C23955 INPUT_3 INVX1_LOC_48/Y 0.05fF
C23956 INVX1_LOC_20/Y NAND2X1_LOC_148/B 0.03fF
C23957 INVX1_LOC_596/A INVX1_LOC_159/Y 0.02fF
C23958 INVX1_LOC_93/Y INVX1_LOC_169/A 0.03fF
C23959 INVX1_LOC_65/Y INVX1_LOC_77/Y 0.07fF
C23960 INPUT_0 INVX1_LOC_557/Y 0.02fF
C23961 INVX1_LOC_17/Y INVX1_LOC_565/A 0.02fF
C23962 INVX1_LOC_602/Y INVX1_LOC_684/Y 0.03fF
C23963 INVX1_LOC_63/Y INVX1_LOC_618/Y 0.19fF
C23964 INVX1_LOC_384/A INVX1_LOC_6/Y 0.19fF
C23965 NAND2X1_LOC_543/B INVX1_LOC_347/A 0.03fF
C23966 INVX1_LOC_190/Y INVX1_LOC_26/Y 0.04fF
C23967 INVX1_LOC_207/A NAND2X1_LOC_240/A 0.02fF
C23968 INVX1_LOC_320/Y INVX1_LOC_9/Y 0.02fF
C23969 INVX1_LOC_235/Y INVX1_LOC_230/Y 0.31fF
C23970 NAND2X1_LOC_572/a_36_24# INVX1_LOC_117/Y 0.01fF
C23971 INVX1_LOC_12/Y INVX1_LOC_681/Y 0.10fF
C23972 INVX1_LOC_686/A INVX1_LOC_32/Y 0.08fF
C23973 NAND2X1_LOC_48/Y INVX1_LOC_172/A 0.26fF
C23974 INVX1_LOC_20/Y INVX1_LOC_69/Y 7.96fF
C23975 INVX1_LOC_335/Y INVX1_LOC_513/A 0.03fF
C23976 INVX1_LOC_93/Y INVX1_LOC_633/Y 0.07fF
C23977 INVX1_LOC_401/A INVX1_LOC_66/A 0.01fF
C23978 INVX1_LOC_12/Y INPUT_1 0.19fF
C23979 NAND2X1_LOC_493/B INVX1_LOC_63/Y 0.01fF
C23980 INVX1_LOC_54/Y NAND2X1_LOC_316/a_36_24# 0.00fF
C23981 NAND2X1_LOC_507/A INVX1_LOC_600/A 0.03fF
C23982 INVX1_LOC_421/A NAND2X1_LOC_527/a_36_24# 0.00fF
C23983 INVX1_LOC_290/A INVX1_LOC_263/Y 0.14fF
C23984 INVX1_LOC_556/Y INVX1_LOC_108/Y 0.01fF
C23985 INVX1_LOC_586/A INVX1_LOC_242/Y 0.13fF
C23986 INVX1_LOC_76/Y INVX1_LOC_376/Y 0.03fF
C23987 INVX1_LOC_72/Y INVX1_LOC_26/Y 0.01fF
C23988 INVX1_LOC_666/A NAND2X1_LOC_845/B 0.03fF
C23989 INVX1_LOC_416/A INVX1_LOC_304/Y 0.01fF
C23990 INVX1_LOC_584/A INVX1_LOC_505/Y 0.02fF
C23991 INVX1_LOC_89/Y NAND2X1_LOC_302/A 0.02fF
C23992 NAND2X1_LOC_301/a_36_24# INVX1_LOC_160/A 0.00fF
C23993 INVX1_LOC_401/Y INVX1_LOC_58/Y 0.05fF
C23994 INVX1_LOC_613/Y INVX1_LOC_6/Y 0.01fF
C23995 INVX1_LOC_81/Y INVX1_LOC_198/A 0.01fF
C23996 INVX1_LOC_522/A INVX1_LOC_330/A 0.03fF
C23997 INVX1_LOC_548/A NAND2X1_LOC_706/B 0.28fF
C23998 NAND2X1_LOC_65/a_36_24# NAND2X1_LOC_786/B 0.00fF
C23999 INVX1_LOC_54/Y NAND2X1_LOC_708/A 0.03fF
C24000 NAND2X1_LOC_612/A INVX1_LOC_6/Y 0.02fF
C24001 INVX1_LOC_567/Y INVX1_LOC_66/A 0.09fF
C24002 INVX1_LOC_573/Y INVX1_LOC_514/Y 0.01fF
C24003 NAND2X1_LOC_97/B INVX1_LOC_58/Y 0.04fF
C24004 INVX1_LOC_145/Y INVX1_LOC_6/Y 8.10fF
C24005 INVX1_LOC_493/A NAND2X1_LOC_634/a_36_24# 0.02fF
C24006 INVX1_LOC_169/A NAND2X1_LOC_487/a_36_24# 0.00fF
C24007 NAND2X1_LOC_775/B INVX1_LOC_31/Y 0.07fF
C24008 INVX1_LOC_300/A INVX1_LOC_69/Y 0.14fF
C24009 INVX1_LOC_99/Y NAND2X1_LOC_827/Y 0.01fF
C24010 INVX1_LOC_491/A INVX1_LOC_492/Y 0.07fF
C24011 NAND2X1_LOC_756/Y INVX1_LOC_79/A 0.12fF
C24012 NAND2X1_LOC_837/A INVX1_LOC_59/Y 0.01fF
C24013 INVX1_LOC_17/Y NAND2X1_LOC_586/Y 0.05fF
C24014 INVX1_LOC_69/Y INVX1_LOC_197/Y 0.04fF
C24015 INVX1_LOC_293/Y INVX1_LOC_79/A 0.05fF
C24016 INVX1_LOC_402/A INVX1_LOC_9/Y 0.00fF
C24017 INVX1_LOC_479/Y INVX1_LOC_77/Y 0.03fF
C24018 INVX1_LOC_638/Y INVX1_LOC_259/Y 0.22fF
C24019 INVX1_LOC_513/Y NAND2X1_LOC_594/Y 0.00fF
C24020 INVX1_LOC_402/Y NAND2X1_LOC_136/Y 0.01fF
C24021 INVX1_LOC_164/Y INVX1_LOC_496/A 0.02fF
C24022 INVX1_LOC_170/A INPUT_1 0.01fF
C24023 INVX1_LOC_160/A INVX1_LOC_79/A 0.03fF
C24024 INVX1_LOC_6/Y INVX1_LOC_433/A 0.05fF
C24025 INVX1_LOC_421/A INVX1_LOC_234/Y 0.02fF
C24026 INVX1_LOC_199/Y NAND2X1_LOC_203/a_36_24# 0.06fF
C24027 NAND2X1_LOC_174/B INVX1_LOC_245/A 0.05fF
C24028 INVX1_LOC_469/A INVX1_LOC_347/A 0.06fF
C24029 NAND2X1_LOC_148/B INVX1_LOC_655/A 0.16fF
C24030 INVX1_LOC_488/A INPUT_1 0.01fF
C24031 INVX1_LOC_54/Y INVX1_LOC_369/Y 0.10fF
C24032 NAND2X1_LOC_528/Y INVX1_LOC_50/Y 0.25fF
C24033 INVX1_LOC_41/Y INVX1_LOC_670/A 0.15fF
C24034 INVX1_LOC_479/A INVX1_LOC_50/Y 4.66fF
C24035 INVX1_LOC_11/A INVX1_LOC_46/Y 0.00fF
C24036 INVX1_LOC_491/A INVX1_LOC_168/Y 0.03fF
C24037 NAND2X1_LOC_768/B INVX1_LOC_124/A 0.04fF
C24038 INVX1_LOC_97/A INVX1_LOC_615/Y 0.03fF
C24039 NAND2X1_LOC_543/B NAND2X1_LOC_176/Y 0.07fF
C24040 INVX1_LOC_328/Y INVX1_LOC_90/Y 0.50fF
C24041 INVX1_LOC_62/Y NAND2X1_LOC_258/Y 0.38fF
C24042 INVX1_LOC_50/Y NAND2X1_LOC_468/a_36_24# 0.00fF
C24043 INVX1_LOC_682/A INVX1_LOC_100/Y 0.00fF
C24044 INVX1_LOC_58/Y NAND2X1_LOC_248/B 0.00fF
C24045 INVX1_LOC_26/Y NAND2X1_LOC_84/a_36_24# 0.00fF
C24046 INVX1_LOC_487/Y INVX1_LOC_488/A 0.05fF
C24047 INVX1_LOC_655/A INVX1_LOC_667/A 0.04fF
C24048 INVX1_LOC_459/Y INVX1_LOC_638/A 0.01fF
C24049 INVX1_LOC_134/Y INVX1_LOC_109/Y 0.07fF
C24050 INVX1_LOC_666/Y INVX1_LOC_9/Y 0.14fF
C24051 INVX1_LOC_395/A INVX1_LOC_307/Y 0.00fF
C24052 INVX1_LOC_62/Y NAND2X1_LOC_545/A 0.01fF
C24053 INVX1_LOC_301/A INVX1_LOC_586/A 0.11fF
C24054 INVX1_LOC_66/A INVX1_LOC_92/A 0.10fF
C24055 INVX1_LOC_395/A NAND2X1_LOC_317/B 0.16fF
C24056 INVX1_LOC_395/A INVX1_LOC_97/A 0.39fF
C24057 INVX1_LOC_112/Y INVX1_LOC_74/Y 0.21fF
C24058 INVX1_LOC_68/Y INVX1_LOC_203/Y 0.04fF
C24059 INVX1_LOC_62/Y INVX1_LOC_653/Y 0.80fF
C24060 INVX1_LOC_53/Y INVX1_LOC_638/A 0.07fF
C24061 INVX1_LOC_62/Y INVX1_LOC_666/Y 0.03fF
C24062 VDD INVX1_LOC_28/Y 0.21fF
C24063 INVX1_LOC_395/A NAND2X1_LOC_613/Y 0.00fF
C24064 INPUT_0 INVX1_LOC_381/A 0.07fF
C24065 INVX1_LOC_617/A INVX1_LOC_118/Y 0.01fF
C24066 INVX1_LOC_20/Y NAND2X1_LOC_537/B 0.03fF
C24067 INVX1_LOC_259/A INVX1_LOC_51/Y 0.01fF
C24068 INVX1_LOC_395/A INVX1_LOC_169/A 0.03fF
C24069 VDD INVX1_LOC_385/Y 0.30fF
C24070 INPUT_0 INVX1_LOC_320/A 0.06fF
C24071 INVX1_LOC_435/Y INVX1_LOC_661/A 0.02fF
C24072 INPUT_6 INVX1_LOC_1/Y 0.01fF
C24073 INVX1_LOC_20/Y NAND2X1_LOC_419/a_36_24# 0.00fF
C24074 INVX1_LOC_460/Y INVX1_LOC_638/A 0.01fF
C24075 INVX1_LOC_446/Y NAND2X1_LOC_517/Y 0.06fF
C24076 INVX1_LOC_206/Y INVX1_LOC_130/Y 0.01fF
C24077 INVX1_LOC_395/A INVX1_LOC_633/Y 0.03fF
C24078 INVX1_LOC_20/Y INVX1_LOC_586/A 4.37fF
C24079 INVX1_LOC_400/Y INVX1_LOC_80/A 0.03fF
C24080 INVX1_LOC_578/A NAND2X1_LOC_299/Y 0.24fF
C24081 INVX1_LOC_576/A INVX1_LOC_586/A 0.01fF
C24082 VDD INVX1_LOC_315/A 0.00fF
C24083 INVX1_LOC_551/Y NAND2X1_LOC_336/a_36_24# 0.06fF
C24084 NAND2X1_LOC_460/A INVX1_LOC_366/A 0.37fF
C24085 INVX1_LOC_51/Y NAND2X1_LOC_658/a_36_24# 0.00fF
C24086 INVX1_LOC_20/Y INVX1_LOC_312/Y 0.19fF
C24087 INVX1_LOC_296/Y INVX1_LOC_76/Y 0.04fF
C24088 NAND2X1_LOC_373/Y INVX1_LOC_69/Y 0.06fF
C24089 INVX1_LOC_418/A INVX1_LOC_35/Y 0.02fF
C24090 INVX1_LOC_312/Y NAND2X1_LOC_473/a_36_24# 0.00fF
C24091 INVX1_LOC_300/A INVX1_LOC_586/A 0.14fF
C24092 INVX1_LOC_558/A INVX1_LOC_35/Y 0.03fF
C24093 INVX1_LOC_410/Y INVX1_LOC_117/Y 0.07fF
C24094 NAND2X1_LOC_46/a_36_24# INPUT_1 0.00fF
C24095 NAND2X1_LOC_271/B INVX1_LOC_31/Y 0.06fF
C24096 INVX1_LOC_586/A INVX1_LOC_197/Y 0.07fF
C24097 INVX1_LOC_142/A NAND2X1_LOC_156/Y 0.06fF
C24098 VDD INVX1_LOC_493/Y 0.29fF
C24099 INVX1_LOC_575/A INVX1_LOC_555/Y 0.03fF
C24100 INVX1_LOC_449/A NAND2X1_LOC_523/B 0.03fF
C24101 INVX1_LOC_396/A NAND2X1_LOC_506/B 0.02fF
C24102 INVX1_LOC_549/A NAND2X1_LOC_707/B 0.05fF
C24103 INVX1_LOC_428/A INVX1_LOC_54/Y 0.31fF
C24104 INVX1_LOC_238/Y INVX1_LOC_199/Y 0.03fF
C24105 INPUT_0 INVX1_LOC_470/Y 0.01fF
C24106 INVX1_LOC_130/Y INVX1_LOC_686/A 0.02fF
C24107 INVX1_LOC_396/A INVX1_LOC_45/Y 0.01fF
C24108 INVX1_LOC_459/A INVX1_LOC_114/A 0.00fF
C24109 INVX1_LOC_412/Y INVX1_LOC_58/Y 0.03fF
C24110 INVX1_LOC_596/A NAND2X1_LOC_595/Y 0.01fF
C24111 INVX1_LOC_397/A INVX1_LOC_32/Y 0.11fF
C24112 INVX1_LOC_270/A INVX1_LOC_35/Y 0.02fF
C24113 INVX1_LOC_415/Y INVX1_LOC_384/A 0.03fF
C24114 NAND2X1_LOC_150/a_36_24# INPUT_1 0.00fF
C24115 INVX1_LOC_420/Y INVX1_LOC_420/A 0.01fF
C24116 NAND2X1_LOC_13/Y INVX1_LOC_411/A 0.11fF
C24117 NAND2X1_LOC_320/Y INVX1_LOC_134/Y 0.01fF
C24118 NAND2X1_LOC_526/Y INVX1_LOC_387/Y 0.03fF
C24119 INVX1_LOC_266/A NAND2X1_LOC_775/B 0.55fF
C24120 INVX1_LOC_32/Y INVX1_LOC_94/A 0.07fF
C24121 NAND2X1_LOC_517/Y INVX1_LOC_145/Y 0.01fF
C24122 NAND2X1_LOC_697/Y INVX1_LOC_53/Y 0.03fF
C24123 INVX1_LOC_521/Y INVX1_LOC_476/A 0.00fF
C24124 NAND2X1_LOC_685/A INVX1_LOC_137/Y 0.14fF
C24125 INVX1_LOC_84/A INVX1_LOC_83/Y 0.00fF
C24126 INVX1_LOC_293/Y INVX1_LOC_48/Y 0.03fF
C24127 NAND2X1_LOC_845/B NAND2X1_LOC_749/Y 0.02fF
C24128 NAND2X1_LOC_791/B INVX1_LOC_598/A 0.01fF
C24129 INVX1_LOC_639/Y INVX1_LOC_640/A 0.00fF
C24130 INVX1_LOC_584/Y INVX1_LOC_338/Y 0.02fF
C24131 INVX1_LOC_272/Y INVX1_LOC_598/A 0.37fF
C24132 INVX1_LOC_31/Y INVX1_LOC_169/A 0.04fF
C24133 NAND2X1_LOC_332/B INVX1_LOC_6/Y 0.05fF
C24134 INVX1_LOC_67/Y INVX1_LOC_98/Y 0.05fF
C24135 INVX1_LOC_372/Y INVX1_LOC_50/Y 0.05fF
C24136 INVX1_LOC_409/Y INVX1_LOC_347/A 0.01fF
C24137 NAND2X1_LOC_756/Y NAND2X1_LOC_168/a_36_24# 0.00fF
C24138 INVX1_LOC_194/Y INVX1_LOC_600/A 0.12fF
C24139 NAND2X1_LOC_708/A NAND2X1_LOC_677/Y 0.15fF
C24140 INVX1_LOC_35/Y NAND2X1_LOC_755/B 0.06fF
C24141 INPUT_0 INVX1_LOC_100/Y 0.28fF
C24142 INVX1_LOC_547/A NAND2X1_LOC_258/Y 0.15fF
C24143 INVX1_LOC_12/Y INVX1_LOC_50/Y 0.11fF
C24144 INVX1_LOC_68/Y INVX1_LOC_44/Y 0.11fF
C24145 INVX1_LOC_438/A NAND2X1_LOC_528/Y 0.03fF
C24146 INVX1_LOC_249/A INVX1_LOC_93/Y 0.12fF
C24147 INVX1_LOC_266/Y INVX1_LOC_351/A 0.01fF
C24148 INVX1_LOC_31/Y INVX1_LOC_633/Y 0.07fF
C24149 INVX1_LOC_160/A INVX1_LOC_48/Y 0.04fF
C24150 INVX1_LOC_17/Y INVX1_LOC_304/Y 0.41fF
C24151 INVX1_LOC_211/Y INVX1_LOC_35/Y 0.03fF
C24152 NAND2X1_LOC_88/B INVX1_LOC_6/Y 0.59fF
C24153 INVX1_LOC_413/A INVX1_LOC_367/Y 0.00fF
C24154 INVX1_LOC_415/Y INVX1_LOC_145/Y 0.22fF
C24155 NAND2X1_LOC_516/Y INVX1_LOC_100/Y 0.05fF
C24156 INVX1_LOC_504/A INVX1_LOC_345/A 0.01fF
C24157 INVX1_LOC_224/Y INVX1_LOC_75/Y 0.09fF
C24158 INVX1_LOC_672/Y INVX1_LOC_221/Y 0.01fF
C24159 NAND2X1_LOC_460/A INVX1_LOC_6/Y 0.01fF
C24160 INVX1_LOC_586/A NAND2X1_LOC_447/a_36_24# 0.00fF
C24161 INVX1_LOC_12/Y INVX1_LOC_431/Y 0.01fF
C24162 INVX1_LOC_298/Y INVX1_LOC_673/Y 0.15fF
C24163 INPUT_0 INVX1_LOC_74/Y 4.84fF
C24164 INVX1_LOC_558/A INVX1_LOC_518/Y 0.03fF
C24165 INVX1_LOC_166/A INVX1_LOC_516/A 0.00fF
C24166 INVX1_LOC_204/Y INVX1_LOC_635/A 0.01fF
C24167 INVX1_LOC_490/Y INVX1_LOC_62/Y 0.05fF
C24168 INVX1_LOC_266/Y INVX1_LOC_90/Y 0.07fF
C24169 INVX1_LOC_134/Y INVX1_LOC_199/Y 0.07fF
C24170 INVX1_LOC_679/Y INVX1_LOC_66/A 0.00fF
C24171 NAND2X1_LOC_260/a_36_24# INVX1_LOC_661/Y 0.00fF
C24172 INVX1_LOC_527/Y NAND2X1_LOC_720/A 0.08fF
C24173 INVX1_LOC_379/A INVX1_LOC_46/Y 0.17fF
C24174 NAND2X1_LOC_299/Y NAND2X1_LOC_854/a_36_24# 0.01fF
C24175 INVX1_LOC_35/Y INVX1_LOC_46/Y 3.58fF
C24176 INVX1_LOC_169/A NAND2X1_LOC_488/a_36_24# 0.00fF
C24177 INVX1_LOC_47/A INVX1_LOC_199/Y 0.03fF
C24178 INVX1_LOC_578/A INVX1_LOC_75/Y 0.02fF
C24179 NAND2X1_LOC_708/a_36_24# INVX1_LOC_137/Y 0.00fF
C24180 INVX1_LOC_304/A INVX1_LOC_46/Y 0.15fF
C24181 INVX1_LOC_300/A INVX1_LOC_157/Y 0.02fF
C24182 INVX1_LOC_11/Y INVX1_LOC_421/A 0.00fF
C24183 INVX1_LOC_298/A NAND2X1_LOC_720/A 0.12fF
C24184 INVX1_LOC_44/Y INVX1_LOC_600/A 0.07fF
C24185 INVX1_LOC_20/Y NAND2X1_LOC_248/a_36_24# 0.00fF
C24186 INVX1_LOC_534/Y NAND2X1_LOC_829/Y 0.17fF
C24187 NAND2X1_LOC_169/A INVX1_LOC_63/Y 0.08fF
C24188 INVX1_LOC_44/Y INVX1_LOC_64/A 0.06fF
C24189 NAND2X1_LOC_97/B INVX1_LOC_245/A 0.03fF
C24190 NAND2X1_LOC_666/Y INVX1_LOC_526/Y 0.19fF
C24191 INVX1_LOC_224/Y NAND2X1_LOC_271/A 0.00fF
C24192 INVX1_LOC_367/A NAND2X1_LOC_136/Y 0.03fF
C24193 NAND2X1_LOC_333/A INVX1_LOC_50/Y 0.00fF
C24194 INVX1_LOC_681/Y INVX1_LOC_66/A 0.20fF
C24195 INVX1_LOC_31/Y NAND2X1_LOC_119/a_36_24# 0.00fF
C24196 INVX1_LOC_166/A INVX1_LOC_93/Y 0.14fF
C24197 INVX1_LOC_261/Y GATE_865 0.01fF
C24198 NAND2X1_LOC_121/a_36_24# INVX1_LOC_41/Y 0.01fF
C24199 INVX1_LOC_353/Y INVX1_LOC_62/Y 0.02fF
C24200 INVX1_LOC_31/Y INVX1_LOC_490/A 0.03fF
C24201 NAND2X1_LOC_189/a_36_24# INVX1_LOC_99/Y 0.00fF
C24202 INPUT_1 INVX1_LOC_66/A 0.16fF
C24203 INVX1_LOC_498/A NAND2X1_LOC_638/a_36_24# 0.02fF
C24204 INVX1_LOC_31/Y INVX1_LOC_317/A 0.01fF
C24205 INVX1_LOC_575/A INVX1_LOC_662/A 0.02fF
C24206 INVX1_LOC_490/Y NAND2X1_LOC_269/a_36_24# 0.00fF
C24207 INVX1_LOC_588/Y INVX1_LOC_675/A 0.07fF
C24208 NAND2X1_LOC_111/Y INVX1_LOC_93/Y 0.14fF
C24209 INVX1_LOC_241/Y INVX1_LOC_655/A 0.03fF
C24210 INVX1_LOC_673/A INVX1_LOC_660/Y 0.11fF
C24211 NAND2X1_LOC_128/B INVX1_LOC_6/Y 0.01fF
C24212 INVX1_LOC_607/Y INVX1_LOC_100/Y 0.15fF
C24213 INVX1_LOC_442/A INVX1_LOC_92/A 0.09fF
C24214 INVX1_LOC_49/Y NAND2X1_LOC_619/Y 0.01fF
C24215 INVX1_LOC_588/Y NAND2X1_LOC_334/B 0.14fF
C24216 INVX1_LOC_665/A INVX1_LOC_99/Y 0.04fF
C24217 INVX1_LOC_213/Y NAND2X1_LOC_833/B 0.01fF
C24218 INVX1_LOC_280/Y INVX1_LOC_245/A 0.01fF
C24219 NAND2X1_LOC_369/a_36_24# INVX1_LOC_347/A 0.00fF
C24220 NAND2X1_LOC_123/A INVX1_LOC_74/Y 0.08fF
C24221 INVX1_LOC_400/A INVX1_LOC_531/Y 0.04fF
C24222 INVX1_LOC_476/A NAND2X1_LOC_846/B 0.02fF
C24223 INVX1_LOC_488/A INVX1_LOC_50/Y 0.01fF
C24224 NAND2X1_LOC_181/a_36_24# INVX1_LOC_62/Y 0.01fF
C24225 INVX1_LOC_93/Y NAND2X1_LOC_136/Y 0.15fF
C24226 INVX1_LOC_6/Y INVX1_LOC_484/Y 0.01fF
C24227 NAND2X1_LOC_451/B INVX1_LOC_685/Y 0.05fF
C24228 INVX1_LOC_391/Y NAND2X1_LOC_844/A 0.00fF
C24229 INVX1_LOC_35/Y INVX1_LOC_75/A 0.00fF
C24230 INVX1_LOC_93/Y INVX1_LOC_531/Y 0.21fF
C24231 INVX1_LOC_298/A INVX1_LOC_74/Y 0.03fF
C24232 INVX1_LOC_298/A INVX1_LOC_660/A 0.00fF
C24233 NAND2X1_LOC_527/Y INVX1_LOC_75/Y 0.02fF
C24234 INVX1_LOC_6/Y INVX1_LOC_487/A 0.03fF
C24235 INVX1_LOC_74/Y INVX1_LOC_498/A 4.95fF
C24236 INVX1_LOC_652/A INVX1_LOC_49/Y 0.00fF
C24237 INVX1_LOC_145/Y INVX1_LOC_636/A 0.07fF
C24238 INVX1_LOC_360/A INVX1_LOC_634/Y 0.05fF
C24239 INVX1_LOC_93/Y INVX1_LOC_528/Y 0.01fF
C24240 NAND2X1_LOC_520/A INVX1_LOC_41/Y 0.02fF
C24241 INVX1_LOC_116/Y INVX1_LOC_92/A 0.07fF
C24242 INVX1_LOC_47/Y INVX1_LOC_505/Y 0.07fF
C24243 NAND2X1_LOC_847/A INVX1_LOC_669/A 0.47fF
C24244 INVX1_LOC_463/A INVX1_LOC_540/Y 0.02fF
C24245 INVX1_LOC_120/Y INVX1_LOC_75/Y 0.01fF
C24246 NAND2X1_LOC_527/Y NAND2X1_LOC_271/A 0.03fF
C24247 INVX1_LOC_655/A NAND2X1_LOC_248/a_36_24# 0.01fF
C24248 NAND2X1_LOC_69/B INVX1_LOC_45/Y 0.02fF
C24249 NAND2X1_LOC_537/A INVX1_LOC_173/A 0.07fF
C24250 INVX1_LOC_505/Y INVX1_LOC_119/Y 0.26fF
C24251 NAND2X1_LOC_373/Y INVX1_LOC_586/A 0.01fF
C24252 INVX1_LOC_255/A INVX1_LOC_92/A 0.07fF
C24253 INVX1_LOC_100/Y INVX1_LOC_211/A 0.14fF
C24254 VDD NAND2X1_LOC_152/Y 0.06fF
C24255 NAND2X1_LOC_271/B INVX1_LOC_51/Y 0.16fF
C24256 NAND2X1_LOC_745/a_36_24# NAND2X1_LOC_781/B 0.01fF
C24257 INVX1_LOC_74/Y INVX1_LOC_211/A 0.00fF
C24258 INVX1_LOC_418/A NAND2X1_LOC_544/a_36_24# 0.02fF
C24259 VDD INVX1_LOC_90/A -0.00fF
C24260 INVX1_LOC_73/Y NAND2X1_LOC_378/Y 0.02fF
C24261 NAND2X1_LOC_69/B NAND2X1_LOC_69/Y 0.15fF
C24262 NAND2X1_LOC_45/Y INVX1_LOC_80/A 1.71fF
C24263 VDD INVX1_LOC_680/Y 0.05fF
C24264 INVX1_LOC_21/Y INVX1_LOC_616/Y 0.00fF
C24265 NAND2X1_LOC_543/B INVX1_LOC_252/Y 0.03fF
C24266 INVX1_LOC_276/A NAND2X1_LOC_142/Y 0.37fF
C24267 NAND2X1_LOC_593/a_36_24# INVX1_LOC_51/Y 0.01fF
C24268 NAND2X1_LOC_97/A NAND2X1_LOC_97/a_36_24# 0.00fF
C24269 NAND2X1_LOC_89/a_36_24# INVX1_LOC_94/A 0.00fF
C24270 INVX1_LOC_438/A INVX1_LOC_12/Y 2.54fF
C24271 VDD INVX1_LOC_186/A -0.00fF
C24272 VDD INVX1_LOC_685/A -0.00fF
C24273 VDD INVX1_LOC_176/A 0.00fF
C24274 INVX1_LOC_118/Y NAND2X1_LOC_130/Y 0.02fF
C24275 NAND2X1_LOC_88/B NAND2X1_LOC_206/a_36_24# 0.00fF
C24276 NAND2X1_LOC_498/Y INVX1_LOC_80/A 0.14fF
C24277 INVX1_LOC_435/Y INVX1_LOC_449/A 0.10fF
C24278 INVX1_LOC_570/A INVX1_LOC_80/A 3.31fF
C24279 VDD INVX1_LOC_349/A 0.00fF
C24280 INVX1_LOC_32/A INVX1_LOC_35/Y 0.01fF
C24281 INVX1_LOC_168/A INVX1_LOC_76/Y 0.01fF
C24282 INVX1_LOC_287/Y INVX1_LOC_291/A 0.02fF
C24283 INVX1_LOC_84/A NAND2X1_LOC_493/B 0.03fF
C24284 NAND2X1_LOC_45/Y INVX1_LOC_11/Y 0.13fF
C24285 NAND2X1_LOC_252/Y INVX1_LOC_220/A 0.20fF
C24286 NAND2X1_LOC_7/Y INVX1_LOC_6/Y 0.08fF
C24287 INVX1_LOC_129/A INVX1_LOC_412/A 0.02fF
C24288 NAND2X1_LOC_788/A INPUT_1 0.03fF
C24289 VDD INVX1_LOC_354/Y 0.21fF
C24290 INVX1_LOC_20/Y NAND2X1_LOC_791/B 0.54fF
C24291 INVX1_LOC_190/Y INVX1_LOC_81/Y 0.01fF
C24292 INVX1_LOC_270/A NAND2X1_LOC_336/a_36_24# 0.02fF
C24293 INVX1_LOC_20/Y INVX1_LOC_272/Y 0.05fF
C24294 INVX1_LOC_45/Y INVX1_LOC_155/Y 0.03fF
C24295 NAND2X1_LOC_750/Y INVX1_LOC_54/Y 0.05fF
C24296 INVX1_LOC_23/Y INPUT_2 0.00fF
C24297 INVX1_LOC_523/A INVX1_LOC_556/Y -0.03fF
C24298 INVX1_LOC_546/A INVX1_LOC_251/Y 0.01fF
C24299 INVX1_LOC_51/A INVX1_LOC_54/Y 0.00fF
C24300 INVX1_LOC_147/A INVX1_LOC_147/Y 0.10fF
C24301 INVX1_LOC_11/Y NAND2X1_LOC_498/Y 0.09fF
C24302 NAND2X1_LOC_710/B INVX1_LOC_670/A 0.01fF
C24303 INVX1_LOC_80/A INVX1_LOC_377/Y 0.14fF
C24304 INVX1_LOC_11/Y INVX1_LOC_570/A 0.07fF
C24305 INVX1_LOC_434/A NAND2X1_LOC_252/Y 0.09fF
C24306 NAND2X1_LOC_299/Y INVX1_LOC_686/A 0.02fF
C24307 INVX1_LOC_278/A NAND2X1_LOC_482/Y 0.01fF
C24308 INVX1_LOC_333/A NAND2X1_LOC_408/a_36_24# 0.02fF
C24309 INVX1_LOC_235/Y NAND2X1_LOC_296/Y 0.04fF
C24310 INVX1_LOC_626/Y INVX1_LOC_6/Y 0.01fF
C24311 VDD INVX1_LOC_420/A 0.00fF
C24312 INVX1_LOC_81/Y INVX1_LOC_72/Y 0.03fF
C24313 INVX1_LOC_366/A INVX1_LOC_197/Y 0.00fF
C24314 INVX1_LOC_65/Y INVX1_LOC_159/Y 0.03fF
C24315 INVX1_LOC_166/A INVX1_LOC_395/A 0.05fF
C24316 VDD INVX1_LOC_170/Y 0.40fF
C24317 NAND2X1_LOC_331/A INVX1_LOC_542/Y 0.03fF
C24318 INVX1_LOC_53/Y INVX1_LOC_134/Y 0.24fF
C24319 INVX1_LOC_291/A NAND2X1_LOC_755/B 0.01fF
C24320 INVX1_LOC_442/A INPUT_1 1.28fF
C24321 INVX1_LOC_420/Y NAND2X1_LOC_292/Y 0.01fF
C24322 INVX1_LOC_7/A INVX1_LOC_245/A 0.01fF
C24323 NAND2X1_LOC_318/A INVX1_LOC_35/Y 0.56fF
C24324 VDD INVX1_LOC_277/Y 0.21fF
C24325 NAND2X1_LOC_48/Y INVX1_LOC_53/Y 0.16fF
C24326 NAND2X1_LOC_78/a_36_24# INVX1_LOC_80/A 0.00fF
C24327 INVX1_LOC_166/A INVX1_LOC_362/Y 0.18fF
C24328 VDD INVX1_LOC_399/Y 0.35fF
C24329 INVX1_LOC_206/Y INVX1_LOC_551/A 0.02fF
C24330 INVX1_LOC_80/A INVX1_LOC_99/Y 0.28fF
C24331 NAND2X1_LOC_768/A INVX1_LOC_99/Y 0.02fF
C24332 INVX1_LOC_51/Y INVX1_LOC_490/A 0.05fF
C24333 INVX1_LOC_579/Y INVX1_LOC_99/Y 0.03fF
C24334 INVX1_LOC_145/Y INVX1_LOC_29/Y 0.01fF
C24335 NAND2X1_LOC_756/Y INVX1_LOC_396/A 0.14fF
C24336 INVX1_LOC_185/Y INVX1_LOC_633/A 0.00fF
C24337 INVX1_LOC_45/Y NAND2X1_LOC_486/A 0.01fF
C24338 INVX1_LOC_544/A INVX1_LOC_679/Y 0.04fF
C24339 NAND2X1_LOC_467/A INVX1_LOC_93/Y 0.00fF
C24340 INVX1_LOC_563/A INVX1_LOC_35/Y 0.01fF
C24341 INPUT_0 NAND2X1_LOC_558/B 0.01fF
C24342 INVX1_LOC_21/Y INVX1_LOC_435/A 0.03fF
C24343 INVX1_LOC_429/Y NAND2X1_LOC_555/B 0.09fF
C24344 NAND2X1_LOC_122/Y NAND2X1_LOC_586/Y 0.06fF
C24345 INVX1_LOC_17/Y NAND2X1_LOC_673/a_36_24# 0.00fF
C24346 INVX1_LOC_166/A INVX1_LOC_683/Y 0.02fF
C24347 NAND2X1_LOC_199/a_36_24# INVX1_LOC_46/Y 0.01fF
C24348 INVX1_LOC_20/Y INVX1_LOC_6/Y 0.21fF
C24349 INVX1_LOC_326/Y INPUT_2 0.16fF
C24350 NAND2X1_LOC_707/A INVX1_LOC_496/A 0.02fF
C24351 INPUT_0 INVX1_LOC_79/A 0.20fF
C24352 INVX1_LOC_395/A NAND2X1_LOC_136/Y 0.03fF
C24353 INVX1_LOC_25/Y INVX1_LOC_6/A 0.01fF
C24354 NAND2X1_LOC_755/B NAND2X1_LOC_837/B 0.02fF
C24355 INVX1_LOC_568/Y INVX1_LOC_492/A 0.00fF
C24356 INVX1_LOC_11/Y INVX1_LOC_99/Y 0.29fF
C24357 INVX1_LOC_194/A INVX1_LOC_230/A 0.07fF
C24358 INVX1_LOC_202/Y INVX1_LOC_35/Y 0.03fF
C24359 INVX1_LOC_53/A NAND2X1_LOC_47/a_36_24# 0.02fF
C24360 INVX1_LOC_428/Y INVX1_LOC_437/A 0.02fF
C24361 GATE_865 INVX1_LOC_290/A 0.02fF
C24362 INVX1_LOC_550/Y INVX1_LOC_35/Y 0.01fF
C24363 NAND2X1_LOC_516/Y INVX1_LOC_79/A 0.00fF
C24364 INVX1_LOC_321/A INVX1_LOC_245/A 0.01fF
C24365 INVX1_LOC_576/A INVX1_LOC_6/Y 0.01fF
C24366 INVX1_LOC_400/Y INVX1_LOC_319/A 0.03fF
C24367 INVX1_LOC_80/A NAND2X1_LOC_306/a_36_24# 0.01fF
C24368 INVX1_LOC_469/Y NAND2X1_LOC_123/A 0.00fF
C24369 INVX1_LOC_257/Y INVX1_LOC_74/Y 0.21fF
C24370 INVX1_LOC_578/A NAND2X1_LOC_441/a_36_24# 0.00fF
C24371 INPUT_7 INVX1_LOC_3/A 0.01fF
C24372 INVX1_LOC_206/Y INVX1_LOC_75/Y 0.14fF
C24373 INVX1_LOC_395/A INVX1_LOC_531/Y 0.08fF
C24374 INVX1_LOC_318/Y INVX1_LOC_199/Y 0.21fF
C24375 INVX1_LOC_439/Y INVX1_LOC_451/A 0.03fF
C24376 INVX1_LOC_116/Y INPUT_1 0.10fF
C24377 INVX1_LOC_80/A INVX1_LOC_47/Y 0.25fF
C24378 INVX1_LOC_550/A INVX1_LOC_35/Y 0.00fF
C24379 INVX1_LOC_134/Y NAND2X1_LOC_274/Y 0.07fF
C24380 NAND2X1_LOC_789/A INVX1_LOC_145/Y 0.01fF
C24381 INVX1_LOC_338/A INVX1_LOC_46/Y 0.01fF
C24382 INVX1_LOC_159/A INVX1_LOC_50/Y 0.02fF
C24383 INVX1_LOC_421/A INVX1_LOC_367/Y 0.07fF
C24384 INVX1_LOC_395/A INVX1_LOC_528/Y 0.05fF
C24385 INVX1_LOC_384/A INVX1_LOC_100/Y 0.07fF
C24386 VDD INVX1_LOC_611/A -0.00fF
C24387 INVX1_LOC_300/A INVX1_LOC_6/Y 0.02fF
C24388 INVX1_LOC_376/A INVX1_LOC_188/Y 0.07fF
C24389 INVX1_LOC_254/Y INVX1_LOC_117/Y 0.02fF
C24390 INVX1_LOC_304/Y INVX1_LOC_230/Y 0.01fF
C24391 INVX1_LOC_387/Y INVX1_LOC_35/Y 0.00fF
C24392 INVX1_LOC_288/A INVX1_LOC_74/Y 0.27fF
C24393 INVX1_LOC_6/Y INVX1_LOC_197/Y 0.02fF
C24394 INVX1_LOC_183/A NAND2X1_LOC_616/Y 0.12fF
C24395 INVX1_LOC_588/Y INVX1_LOC_31/Y 10.31fF
C24396 NAND2X1_LOC_548/B INVX1_LOC_422/A 0.07fF
C24397 INVX1_LOC_379/A INVX1_LOC_49/Y 0.37fF
C24398 NAND2X1_LOC_820/A INVX1_LOC_655/A 0.05fF
C24399 INVX1_LOC_504/A INVX1_LOC_347/Y 0.01fF
C24400 INVX1_LOC_11/Y INVX1_LOC_47/Y 2.83fF
C24401 INVX1_LOC_49/Y INVX1_LOC_35/Y 3.08fF
C24402 INVX1_LOC_41/Y INVX1_LOC_59/A 0.03fF
C24403 INVX1_LOC_166/A INVX1_LOC_31/Y 0.09fF
C24404 INVX1_LOC_80/A INVX1_LOC_119/Y 0.16fF
C24405 INVX1_LOC_11/Y NAND2X1_LOC_557/B 0.22fF
C24406 INVX1_LOC_50/Y INVX1_LOC_66/A 0.17fF
C24407 INVX1_LOC_255/A INPUT_1 0.75fF
C24408 INVX1_LOC_53/Y NAND2X1_LOC_791/a_36_24# 0.00fF
C24409 NAND2X1_LOC_336/a_36_24# INVX1_LOC_75/A 0.00fF
C24410 INVX1_LOC_385/Y INVX1_LOC_430/Y 0.03fF
C24411 INVX1_LOC_353/A INVX1_LOC_252/Y 0.00fF
C24412 INVX1_LOC_89/Y INVX1_LOC_187/Y 0.03fF
C24413 NAND2X1_LOC_106/Y INVX1_LOC_69/Y 0.01fF
C24414 INPUT_7 INVX1_LOC_74/A 0.41fF
C24415 INVX1_LOC_100/Y INVX1_LOC_145/Y 2.44fF
C24416 INVX1_LOC_379/A NAND2X1_LOC_296/a_36_24# 0.00fF
C24417 INVX1_LOC_93/Y INVX1_LOC_411/Y 0.01fF
C24418 NAND2X1_LOC_84/B INVX1_LOC_9/Y 0.09fF
C24419 INVX1_LOC_431/Y INVX1_LOC_296/A 0.03fF
C24420 INVX1_LOC_89/Y NAND2X1_LOC_284/A 0.01fF
C24421 INVX1_LOC_575/Y INVX1_LOC_662/A 0.06fF
C24422 INVX1_LOC_49/Y INVX1_LOC_620/A 0.66fF
C24423 NAND2X1_LOC_788/a_36_24# INVX1_LOC_79/A 0.00fF
C24424 INVX1_LOC_11/Y INVX1_LOC_119/Y 1.19fF
C24425 INVX1_LOC_11/Y NAND2X1_LOC_66/Y 0.08fF
C24426 INVX1_LOC_662/Y NAND2X1_LOC_342/B 0.06fF
C24427 INVX1_LOC_166/A INVX1_LOC_128/A 0.00fF
C24428 INVX1_LOC_400/A INVX1_LOC_41/Y 0.10fF
C24429 INVX1_LOC_145/Y INVX1_LOC_74/Y 0.03fF
C24430 INVX1_LOC_392/A INVX1_LOC_41/Y 0.01fF
C24431 INVX1_LOC_58/Y INVX1_LOC_646/Y 0.15fF
C24432 INVX1_LOC_670/A INVX1_LOC_128/Y 0.01fF
C24433 INVX1_LOC_298/A INVX1_LOC_79/A 0.03fF
C24434 INVX1_LOC_6/Y INVX1_LOC_655/A 0.09fF
C24435 INVX1_LOC_662/A INVX1_LOC_132/A 0.06fF
C24436 INVX1_LOC_47/Y NAND2X1_LOC_433/Y 0.05fF
C24437 INVX1_LOC_253/Y NAND2X1_LOC_274/B 0.00fF
C24438 NAND2X1_LOC_123/a_36_24# INVX1_LOC_62/Y 0.01fF
C24439 INVX1_LOC_31/Y INVX1_LOC_531/Y 0.46fF
C24440 INVX1_LOC_117/Y NAND2X1_LOC_528/Y 0.28fF
C24441 INVX1_LOC_93/Y INVX1_LOC_41/Y 0.36fF
C24442 INVX1_LOC_535/Y INVX1_LOC_62/Y 0.03fF
C24443 NAND2X1_LOC_833/B NAND2X1_LOC_258/Y 0.01fF
C24444 INVX1_LOC_54/Y INVX1_LOC_441/A 0.01fF
C24445 INVX1_LOC_13/Y NAND2X1_LOC_84/B 0.02fF
C24446 INVX1_LOC_108/Y INVX1_LOC_109/A 0.15fF
C24447 INVX1_LOC_50/Y NAND2X1_LOC_621/B 0.03fF
C24448 INVX1_LOC_199/Y INVX1_LOC_90/Y 0.17fF
C24449 NAND2X1_LOC_189/a_36_24# INVX1_LOC_15/Y 0.00fF
C24450 NAND2X1_LOC_274/B INVX1_LOC_63/Y 0.01fF
C24451 INVX1_LOC_117/Y INVX1_LOC_479/A 0.53fF
C24452 INVX1_LOC_69/Y NAND2X1_LOC_123/B 0.13fF
C24453 NAND2X1_LOC_173/a_36_24# INVX1_LOC_354/A 0.01fF
C24454 INVX1_LOC_50/Y NAND2X1_LOC_646/B 0.07fF
C24455 INVX1_LOC_153/A NAND2X1_LOC_231/B 0.03fF
C24456 INVX1_LOC_31/Y NAND2X1_LOC_433/a_36_24# 0.00fF
C24457 INVX1_LOC_675/A INVX1_LOC_41/Y 0.07fF
C24458 INVX1_LOC_46/Y INVX1_LOC_488/Y 0.04fF
C24459 NAND2X1_LOC_433/Y INVX1_LOC_119/Y 0.75fF
C24460 INVX1_LOC_69/Y NAND2X1_LOC_428/Y 0.06fF
C24461 INVX1_LOC_457/Y VDD 0.21fF
C24462 VDD INVX1_LOC_193/Y 0.41fF
C24463 NAND2X1_LOC_97/A NAND2X1_LOC_790/B 0.06fF
C24464 INVX1_LOC_501/A NAND2X1_LOC_832/A 0.04fF
C24465 INVX1_LOC_77/A INVX1_LOC_211/A 0.01fF
C24466 INVX1_LOC_682/Y INVX1_LOC_363/A 0.03fF
C24467 INVX1_LOC_69/Y INVX1_LOC_92/A 0.10fF
C24468 INVX1_LOC_629/A INVX1_LOC_288/A 0.15fF
C24469 NAND2X1_LOC_488/Y INVX1_LOC_388/A 0.03fF
C24470 INVX1_LOC_446/Y INVX1_LOC_450/A 0.09fF
C24471 INVX1_LOC_35/Y INVX1_LOC_297/Y 0.03fF
C24472 INVX1_LOC_302/A INVX1_LOC_362/Y 0.04fF
C24473 INVX1_LOC_134/A INVX1_LOC_442/A 0.05fF
C24474 INVX1_LOC_435/Y INVX1_LOC_651/Y 0.10fF
C24475 NAND2X1_LOC_475/A INVX1_LOC_80/A 0.07fF
C24476 INVX1_LOC_99/Y NAND2X1_LOC_590/a_36_24# 0.00fF
C24477 NAND2X1_LOC_501/a_36_24# INVX1_LOC_384/A 0.01fF
C24478 INVX1_LOC_447/Y VDD 0.36fF
C24479 NAND2X1_LOC_69/B NAND2X1_LOC_673/B 0.12fF
C24480 INVX1_LOC_560/Y NAND2X1_LOC_169/A 0.02fF
C24481 NAND2X1_LOC_331/A NAND2X1_LOC_829/Y 0.01fF
C24482 INVX1_LOC_266/A INVX1_LOC_317/Y 0.17fF
C24483 NAND2X1_LOC_741/a_36_24# INVX1_LOC_632/A 0.01fF
C24484 INPUT_0 INVX1_LOC_417/Y 0.07fF
C24485 NAND2X1_LOC_151/a_36_24# INVX1_LOC_523/A 0.00fF
C24486 NAND2X1_LOC_23/a_36_24# INVX1_LOC_17/Y 0.00fF
C24487 NAND2X1_LOC_69/a_36_24# NAND2X1_LOC_616/Y 0.00fF
C24488 INVX1_LOC_561/A INVX1_LOC_638/A 0.11fF
C24489 INVX1_LOC_11/Y NAND2X1_LOC_475/A 0.10fF
C24490 VDD INVX1_LOC_54/Y 3.94fF
C24491 INVX1_LOC_319/Y INVX1_LOC_99/Y 0.01fF
C24492 NAND2X1_LOC_140/a_36_24# INVX1_LOC_35/Y 0.00fF
C24493 INVX1_LOC_80/A INVX1_LOC_502/Y 0.00fF
C24494 INVX1_LOC_628/A INVX1_LOC_288/A -0.07fF
C24495 INVX1_LOC_21/Y INVX1_LOC_392/Y 0.01fF
C24496 INVX1_LOC_468/Y INVX1_LOC_557/A 0.10fF
C24497 INVX1_LOC_206/Y NAND2X1_LOC_383/a_36_24# 0.00fF
C24498 INVX1_LOC_224/Y INVX1_LOC_227/Y 0.01fF
C24499 VDD INVX1_LOC_611/Y 0.21fF
C24500 INPUT_0 INVX1_LOC_48/Y 0.34fF
C24501 INPUT_0 NAND2X1_LOC_60/a_36_24# 0.00fF
C24502 INVX1_LOC_207/A INVX1_LOC_145/Y 0.00fF
C24503 INVX1_LOC_366/A INVX1_LOC_600/Y 0.00fF
C24504 INPUT_3 INVX1_LOC_28/Y 0.03fF
C24505 VDD NAND2X1_LOC_292/Y -0.00fF
C24506 NAND2X1_LOC_597/a_36_24# INVX1_LOC_50/Y 0.00fF
C24507 INVX1_LOC_257/Y INVX1_LOC_469/Y 0.06fF
C24508 INVX1_LOC_257/Y INVX1_LOC_350/Y -0.00fF
C24509 INVX1_LOC_228/Y INVX1_LOC_54/Y 0.09fF
C24510 INVX1_LOC_408/Y INVX1_LOC_50/Y 0.29fF
C24511 INVX1_LOC_134/A INVX1_LOC_116/Y 0.02fF
C24512 INVX1_LOC_98/A INVX1_LOC_35/Y 0.01fF
C24513 INVX1_LOC_76/Y INVX1_LOC_379/A 0.07fF
C24514 INVX1_LOC_542/A INVX1_LOC_137/Y 0.03fF
C24515 INVX1_LOC_681/A INVX1_LOC_482/A 0.15fF
C24516 INVX1_LOC_335/Y INVX1_LOC_59/A 0.03fF
C24517 INVX1_LOC_17/Y NAND2X1_LOC_180/B 0.00fF
C24518 INVX1_LOC_566/Y INVX1_LOC_99/Y 0.03fF
C24519 INVX1_LOC_76/Y INVX1_LOC_35/Y 0.17fF
C24520 INVX1_LOC_24/A INVX1_LOC_66/A 0.01fF
C24521 INVX1_LOC_51/A INVX1_LOC_89/Y 0.00fF
C24522 INVX1_LOC_442/A INVX1_LOC_50/Y 0.02fF
C24523 VDD INVX1_LOC_521/A -0.00fF
C24524 INVX1_LOC_21/Y INVX1_LOC_367/A 0.01fF
C24525 NAND2X1_LOC_498/Y INVX1_LOC_374/Y 0.05fF
C24526 INVX1_LOC_584/A INVX1_LOC_261/Y 0.01fF
C24527 INVX1_LOC_45/Y INVX1_LOC_315/A 0.01fF
C24528 INVX1_LOC_286/A INVX1_LOC_48/Y 0.01fF
C24529 NAND2X1_LOC_98/a_36_24# INVX1_LOC_95/A 0.02fF
C24530 INVX1_LOC_224/Y INVX1_LOC_120/Y 0.02fF
C24531 INVX1_LOC_288/A INVX1_LOC_469/Y 0.01fF
C24532 NAND2X1_LOC_670/a_36_24# INVX1_LOC_169/A 0.00fF
C24533 INVX1_LOC_450/A INVX1_LOC_433/A 0.32fF
C24534 INVX1_LOC_166/A INVX1_LOC_51/Y 0.06fF
C24535 INVX1_LOC_315/Y INVX1_LOC_93/Y 1.43fF
C24536 INVX1_LOC_26/Y INVX1_LOC_616/Y 0.01fF
C24537 INVX1_LOC_381/A NAND2X1_LOC_297/Y 0.04fF
C24538 INVX1_LOC_395/A INVX1_LOC_411/Y 0.22fF
C24539 INVX1_LOC_17/Y INVX1_LOC_188/Y 0.03fF
C24540 INVX1_LOC_515/Y NAND2X1_LOC_679/B 0.01fF
C24541 INVX1_LOC_578/A INVX1_LOC_120/Y 0.03fF
C24542 NAND2X1_LOC_331/A NAND2X1_LOC_679/A 0.01fF
C24543 NAND2X1_LOC_105/a_36_24# NAND2X1_LOC_106/B 0.02fF
C24544 NAND2X1_LOC_184/Y INVX1_LOC_654/A 0.03fF
C24545 NAND2X1_LOC_636/A INVX1_LOC_62/Y 0.02fF
C24546 INVX1_LOC_21/Y INVX1_LOC_516/A 0.05fF
C24547 INVX1_LOC_677/Y INVX1_LOC_641/Y 0.03fF
C24548 INVX1_LOC_196/A INVX1_LOC_50/Y 0.01fF
C24549 INVX1_LOC_410/Y INVX1_LOC_245/A 0.12fF
C24550 INVX1_LOC_584/A NAND2X1_LOC_431/a_36_24# 0.01fF
C24551 INVX1_LOC_134/A INVX1_LOC_255/A 0.05fF
C24552 INVX1_LOC_372/Y INVX1_LOC_117/Y 0.03fF
C24553 INVX1_LOC_371/Y INVX1_LOC_371/A 0.01fF
C24554 INVX1_LOC_384/A NAND2X1_LOC_181/A 0.02fF
C24555 INVX1_LOC_625/A INVX1_LOC_274/A 0.04fF
C24556 INVX1_LOC_257/Y INVX1_LOC_79/A 0.07fF
C24557 INVX1_LOC_596/A INVX1_LOC_105/Y 0.03fF
C24558 INVX1_LOC_511/A INVX1_LOC_498/A 0.02fF
C24559 INVX1_LOC_367/Y INVX1_LOC_99/Y 0.06fF
C24560 NAND2X1_LOC_704/B INVX1_LOC_47/Y 0.01fF
C24561 VDD INVX1_LOC_388/A -0.00fF
C24562 INVX1_LOC_80/A INVX1_LOC_153/A 0.00fF
C24563 NAND2X1_LOC_666/Y INVX1_LOC_586/A 0.02fF
C24564 INPUT_0 INVX1_LOC_472/Y 0.01fF
C24565 INVX1_LOC_266/A NAND2X1_LOC_111/Y 0.04fF
C24566 INVX1_LOC_324/A INVX1_LOC_46/Y 0.01fF
C24567 INVX1_LOC_362/Y INVX1_LOC_301/Y 0.13fF
C24568 INVX1_LOC_117/Y INVX1_LOC_12/Y 0.17fF
C24569 INVX1_LOC_17/Y INVX1_LOC_478/Y 0.01fF
C24570 NAND2X1_LOC_123/A INVX1_LOC_48/Y 0.01fF
C24571 INVX1_LOC_291/A INVX1_LOC_49/Y 0.07fF
C24572 INVX1_LOC_374/A NAND2X1_LOC_274/B 0.17fF
C24573 NAND2X1_LOC_774/a_36_24# INVX1_LOC_292/Y 0.00fF
C24574 INVX1_LOC_315/Y NAND2X1_LOC_334/B 0.00fF
C24575 INVX1_LOC_522/A NAND2X1_LOC_661/a_36_24# 0.02fF
C24576 INVX1_LOC_632/A INVX1_LOC_498/A 0.07fF
C24577 INVX1_LOC_11/Y NAND2X1_LOC_43/Y 0.05fF
C24578 INVX1_LOC_33/Y INVX1_LOC_48/A -0.00fF
C24579 INVX1_LOC_400/A NAND2X1_LOC_510/a_36_24# 0.02fF
C24580 INVX1_LOC_527/Y INVX1_LOC_59/Y 0.02fF
C24581 INVX1_LOC_384/Y NAND2X1_LOC_555/B 3.33fF
C24582 INVX1_LOC_549/A INVX1_LOC_62/Y 0.06fF
C24583 INVX1_LOC_42/Y NAND2X1_LOC_84/B 0.02fF
C24584 INVX1_LOC_171/A INVX1_LOC_176/A 0.15fF
C24585 INVX1_LOC_21/Y INVX1_LOC_93/Y 0.61fF
C24586 NAND2X1_LOC_727/a_36_24# INVX1_LOC_79/A 0.00fF
C24587 INVX1_LOC_395/A INVX1_LOC_41/Y 1.78fF
C24588 INVX1_LOC_267/Y NAND2X1_LOC_753/Y 0.01fF
C24589 INVX1_LOC_288/A INVX1_LOC_79/A 0.07fF
C24590 INVX1_LOC_53/Y INVX1_LOC_476/A 0.02fF
C24591 NAND2X1_LOC_513/A INVX1_LOC_66/A 0.04fF
C24592 INVX1_LOC_447/Y INVX1_LOC_103/Y 0.01fF
C24593 INVX1_LOC_116/Y INVX1_LOC_50/Y 0.00fF
C24594 INVX1_LOC_333/Y INVX1_LOC_18/Y 0.01fF
C24595 NAND2X1_LOC_492/a_36_24# INVX1_LOC_9/Y 0.00fF
C24596 NAND2X1_LOC_545/B INVX1_LOC_199/Y 0.03fF
C24597 INVX1_LOC_54/Y INVX1_LOC_509/A 0.01fF
C24598 INVX1_LOC_51/Y NAND2X1_LOC_136/Y 0.01fF
C24599 NAND2X1_LOC_331/B INVX1_LOC_74/Y 0.03fF
C24600 INVX1_LOC_436/Y INVX1_LOC_444/A 0.00fF
C24601 NAND2X1_LOC_505/Y INVX1_LOC_531/Y 0.06fF
C24602 INVX1_LOC_17/Y NAND2X1_LOC_387/Y 0.52fF
C24603 VDD INVX1_LOC_619/Y 0.21fF
C24604 INVX1_LOC_6/Y INVX1_LOC_600/Y 0.00fF
C24605 INVX1_LOC_679/Y INVX1_LOC_69/Y 0.03fF
C24606 NAND2X1_LOC_386/a_36_24# INVX1_LOC_298/A 0.00fF
C24607 INVX1_LOC_527/Y INVX1_LOC_48/Y 0.01fF
C24608 INVX1_LOC_89/Y NAND2X1_LOC_413/Y 0.07fF
C24609 NAND2X1_LOC_137/A INVX1_LOC_669/Y 0.02fF
C24610 NAND2X1_LOC_704/B INVX1_LOC_119/Y 0.00fF
C24611 NAND2X1_LOC_332/B INVX1_LOC_100/Y 0.02fF
C24612 INVX1_LOC_288/A INVX1_LOC_460/A 0.07fF
C24613 INVX1_LOC_301/Y INVX1_LOC_683/Y 0.00fF
C24614 INVX1_LOC_51/Y INVX1_LOC_531/Y 0.19fF
C24615 INVX1_LOC_362/Y INVX1_LOC_41/Y 0.09fF
C24616 INVX1_LOC_208/Y INVX1_LOC_209/A 0.44fF
C24617 NAND2X1_LOC_184/Y INVX1_LOC_282/A 0.00fF
C24618 NAND2X1_LOC_181/A INVX1_LOC_145/Y 0.10fF
C24619 INVX1_LOC_602/Y INVX1_LOC_69/Y 0.11fF
C24620 NAND2X1_LOC_174/B NAND2X1_LOC_591/Y 0.02fF
C24621 INVX1_LOC_432/Y INVX1_LOC_47/Y 0.12fF
C24622 INVX1_LOC_335/Y INVX1_LOC_675/A 0.07fF
C24623 INVX1_LOC_54/Y INVX1_LOC_103/Y 0.15fF
C24624 NAND2X1_LOC_148/B INPUT_1 1.46fF
C24625 INVX1_LOC_530/A INVX1_LOC_328/Y 0.04fF
C24626 INVX1_LOC_199/Y INVX1_LOC_98/Y 0.28fF
C24627 INVX1_LOC_320/A INVX1_LOC_242/Y 0.01fF
C24628 INVX1_LOC_183/A NAND2X1_LOC_393/Y 0.02fF
C24629 NAND2X1_LOC_492/a_36_24# INVX1_LOC_62/Y 0.01fF
C24630 NAND2X1_LOC_333/A INVX1_LOC_117/Y 0.03fF
C24631 INVX1_LOC_653/A INVX1_LOC_134/Y 0.05fF
C24632 NAND2X1_LOC_397/a_36_24# INVX1_LOC_183/A 0.00fF
C24633 INVX1_LOC_253/Y INVX1_LOC_159/Y 0.01fF
C24634 INVX1_LOC_586/A NAND2X1_LOC_428/Y 0.03fF
C24635 INVX1_LOC_376/A INVX1_LOC_504/Y 0.03fF
C24636 INVX1_LOC_32/Y NAND2X1_LOC_619/Y 0.01fF
C24637 INVX1_LOC_53/Y INVX1_LOC_90/Y 0.03fF
C24638 INVX1_LOC_683/Y INVX1_LOC_41/Y 0.02fF
C24639 INVX1_LOC_93/Y NAND2X1_LOC_137/A 0.01fF
C24640 INVX1_LOC_49/Y NAND2X1_LOC_837/B 0.15fF
C24641 INVX1_LOC_93/Y INVX1_LOC_555/A 0.01fF
C24642 INVX1_LOC_69/Y INPUT_1 0.10fF
C24643 INVX1_LOC_25/Y INVX1_LOC_50/A 0.01fF
C24644 INVX1_LOC_74/A INVX1_LOC_55/Y 0.02fF
C24645 INVX1_LOC_254/Y INVX1_LOC_58/Y 0.01fF
C24646 INVX1_LOC_230/A INVX1_LOC_9/Y 0.02fF
C24647 INVX1_LOC_62/Y NAND2X1_LOC_656/a_36_24# 0.00fF
C24648 INVX1_LOC_586/A INVX1_LOC_270/Y 0.03fF
C24649 INVX1_LOC_627/Y INVX1_LOC_6/Y 0.01fF
C24650 INVX1_LOC_100/Y NAND2X1_LOC_260/Y 0.02fF
C24651 INVX1_LOC_401/Y INVX1_LOC_652/Y 0.08fF
C24652 INVX1_LOC_379/A NAND2X1_LOC_264/a_36_24# 0.00fF
C24653 INVX1_LOC_533/Y INVX1_LOC_636/A 0.01fF
C24654 INVX1_LOC_435/A INVX1_LOC_26/Y 0.42fF
C24655 INVX1_LOC_525/Y NAND2X1_LOC_753/Y 0.05fF
C24656 INVX1_LOC_294/A INVX1_LOC_328/Y 0.01fF
C24657 INVX1_LOC_145/Y INVX1_LOC_79/A 0.12fF
C24658 INVX1_LOC_99/Y INVX1_LOC_319/A 0.01fF
C24659 INVX1_LOC_93/Y INVX1_LOC_107/Y 0.02fF
C24660 NAND2X1_LOC_399/B INVX1_LOC_11/A 0.31fF
C24661 INVX1_LOC_69/Y INVX1_LOC_292/Y 0.10fF
C24662 NAND2X1_LOC_749/a_36_24# INVX1_LOC_223/Y 0.01fF
C24663 INVX1_LOC_674/A INVX1_LOC_245/A 0.08fF
C24664 INVX1_LOC_145/Y NAND2X1_LOC_631/B 0.03fF
C24665 INVX1_LOC_586/A INVX1_LOC_92/A 0.13fF
C24666 INVX1_LOC_11/A INVX1_LOC_7/Y 0.06fF
C24667 INVX1_LOC_223/Y INVX1_LOC_46/Y 0.01fF
C24668 INVX1_LOC_69/Y INVX1_LOC_284/Y 0.29fF
C24669 INVX1_LOC_20/Y INVX1_LOC_636/A 0.19fF
C24670 INVX1_LOC_99/Y NAND2X1_LOC_843/B 0.48fF
C24671 INVX1_LOC_518/A INVX1_LOC_520/A 0.10fF
C24672 INVX1_LOC_11/Y NAND2X1_LOC_627/Y 0.03fF
C24673 INVX1_LOC_62/Y INVX1_LOC_230/A 0.07fF
C24674 INVX1_LOC_137/Y NAND2X1_LOC_782/a_36_24# 0.00fF
C24675 NAND2X1_LOC_260/a_36_24# INVX1_LOC_655/A 0.01fF
C24676 INVX1_LOC_479/A INVX1_LOC_251/Y 0.01fF
C24677 INVX1_LOC_355/Y INVX1_LOC_114/A 0.02fF
C24678 INVX1_LOC_399/A INVX1_LOC_69/Y 0.04fF
C24679 INVX1_LOC_505/Y INVX1_LOC_505/A 0.00fF
C24680 INVX1_LOC_59/Y INVX1_LOC_211/A 0.02fF
C24681 INVX1_LOC_254/A INVX1_LOC_531/Y 0.02fF
C24682 INVX1_LOC_123/A INVX1_LOC_319/A 0.23fF
C24683 INVX1_LOC_576/A INVX1_LOC_636/A 0.05fF
C24684 INVX1_LOC_99/Y INVX1_LOC_91/Y 0.03fF
C24685 NAND2X1_LOC_128/B INVX1_LOC_100/Y 0.08fF
C24686 INVX1_LOC_32/Y INVX1_LOC_11/A 0.02fF
C24687 INVX1_LOC_31/Y INVX1_LOC_41/Y 0.43fF
C24688 INVX1_LOC_211/A INVX1_LOC_48/Y 0.13fF
C24689 INVX1_LOC_301/Y INVX1_LOC_682/Y 0.12fF
C24690 INVX1_LOC_47/Y NAND2X1_LOC_432/a_36_24# 0.00fF
C24691 INVX1_LOC_253/Y INVX1_LOC_468/A 0.10fF
C24692 INVX1_LOC_74/A INVX1_LOC_18/Y 0.66fF
C24693 INVX1_LOC_300/A INVX1_LOC_636/A 0.15fF
C24694 NAND2X1_LOC_534/Y VDD 0.03fF
C24695 INVX1_LOC_89/Y INVX1_LOC_354/A 0.01fF
C24696 INVX1_LOC_89/Y INVX1_LOC_441/A 0.01fF
C24697 INVX1_LOC_63/Y INVX1_LOC_468/A 0.01fF
C24698 NAND2X1_LOC_542/A INVX1_LOC_75/Y 0.02fF
C24699 INVX1_LOC_519/Y INVX1_LOC_518/A 0.17fF
C24700 INVX1_LOC_100/Y INVX1_LOC_242/Y 0.21fF
C24701 INVX1_LOC_204/Y NAND2X1_LOC_234/Y 0.13fF
C24702 INVX1_LOC_479/A INVX1_LOC_58/Y 0.23fF
C24703 INVX1_LOC_63/Y NAND2X1_LOC_617/a_36_24# 0.00fF
C24704 INVX1_LOC_596/A INVX1_LOC_109/Y 0.03fF
C24705 INVX1_LOC_224/Y INVX1_LOC_206/Y 0.07fF
C24706 NAND2X1_LOC_45/Y INVX1_LOC_393/Y 0.16fF
C24707 INVX1_LOC_49/Y INVX1_LOC_488/Y 0.91fF
C24708 INVX1_LOC_242/Y INVX1_LOC_74/Y 0.10fF
C24709 INVX1_LOC_319/Y NAND2X1_LOC_475/A 0.01fF
C24710 INVX1_LOC_206/Y INVX1_LOC_578/A 0.07fF
C24711 VDD INVX1_LOC_150/Y 0.35fF
C24712 INVX1_LOC_41/Y INVX1_LOC_473/Y 0.01fF
C24713 VDD INVX1_LOC_113/Y 0.26fF
C24714 INVX1_LOC_133/Y NAND2X1_LOC_152/B 0.24fF
C24715 INPUT_0 NAND2X1_LOC_513/Y 0.37fF
C24716 INVX1_LOC_428/A INVX1_LOC_118/Y 0.00fF
C24717 INVX1_LOC_26/Y NAND2X1_LOC_227/A 0.02fF
C24718 VDD INVX1_LOC_171/Y 0.42fF
C24719 INVX1_LOC_21/Y INVX1_LOC_615/Y 0.01fF
C24720 VDD INVX1_LOC_334/Y 0.21fF
C24721 VDD INVX1_LOC_655/Y 0.30fF
C24722 INVX1_LOC_414/A INVX1_LOC_384/A 0.07fF
C24723 NAND2X1_LOC_543/B INVX1_LOC_80/A 0.01fF
C24724 INVX1_LOC_395/A INVX1_LOC_315/Y 0.04fF
C24725 INVX1_LOC_441/Y INVX1_LOC_442/A 0.15fF
C24726 VDD INVX1_LOC_649/Y 0.36fF
C24727 NAND2X1_LOC_245/a_36_24# INVX1_LOC_669/A 0.01fF
C24728 INVX1_LOC_569/A INVX1_LOC_554/Y 0.02fF
C24729 INVX1_LOC_302/A INVX1_LOC_51/Y 0.02fF
C24730 VDD INVX1_LOC_371/Y 0.26fF
C24731 INVX1_LOC_205/Y INVX1_LOC_180/Y 0.02fF
C24732 VDD NAND2X1_LOC_677/Y 0.07fF
C24733 NAND2X1_LOC_797/a_36_24# INVX1_LOC_137/Y 0.00fF
C24734 INVX1_LOC_317/Y NAND2X1_LOC_13/Y 0.06fF
C24735 INVX1_LOC_20/Y INVX1_LOC_269/Y 0.01fF
C24736 INVX1_LOC_578/A INVX1_LOC_686/A 0.06fF
C24737 INVX1_LOC_402/A INVX1_LOC_238/Y 0.01fF
C24738 INVX1_LOC_446/A INVX1_LOC_159/Y 0.20fF
C24739 INVX1_LOC_279/A INVX1_LOC_439/Y 0.06fF
C24740 INVX1_LOC_191/Y INVX1_LOC_145/Y 0.10fF
C24741 INVX1_LOC_432/Y NAND2X1_LOC_475/A 0.01fF
C24742 INVX1_LOC_335/Y INVX1_LOC_395/A 0.12fF
C24743 INVX1_LOC_414/A INVX1_LOC_145/Y 0.01fF
C24744 INVX1_LOC_21/Y INVX1_LOC_395/A 0.35fF
C24745 INVX1_LOC_291/A INVX1_LOC_76/Y 0.01fF
C24746 VDD INVX1_LOC_277/A -0.00fF
C24747 VDD INVX1_LOC_585/Y 0.21fF
C24748 INVX1_LOC_20/Y INVX1_LOC_381/A 0.01fF
C24749 INVX1_LOC_266/A NAND2X1_LOC_322/a_36_24# 0.00fF
C24750 NAND2X1_LOC_750/Y INVX1_LOC_194/Y 0.03fF
C24751 INVX1_LOC_106/A NAND2X1_LOC_108/Y 0.04fF
C24752 INVX1_LOC_80/A INVX1_LOC_131/Y 0.02fF
C24753 NAND2X1_LOC_77/a_36_24# NAND2X1_LOC_513/Y 0.00fF
C24754 INPUT_7 INVX1_LOC_5/Y 0.04fF
C24755 INVX1_LOC_21/Y INVX1_LOC_362/Y 0.10fF
C24756 INVX1_LOC_680/Y INVX1_LOC_45/Y 0.06fF
C24757 VDD INVX1_LOC_395/Y 0.26fF
C24758 INVX1_LOC_269/Y INVX1_LOC_300/A 0.04fF
C24759 INVX1_LOC_20/Y INVX1_LOC_320/A 0.03fF
C24760 VDD INVX1_LOC_89/Y 2.17fF
C24761 INVX1_LOC_180/A INVX1_LOC_145/Y 0.01fF
C24762 INVX1_LOC_398/A INVX1_LOC_97/Y 0.00fF
C24763 INVX1_LOC_45/Y INVX1_LOC_176/A 0.08fF
C24764 INVX1_LOC_192/Y INVX1_LOC_117/Y 0.03fF
C24765 INVX1_LOC_446/Y INVX1_LOC_48/Y 0.07fF
C24766 INVX1_LOC_434/A INVX1_LOC_387/Y 0.01fF
C24767 INVX1_LOC_76/Y INVX1_LOC_338/A 0.01fF
C24768 INVX1_LOC_288/A INVX1_LOC_48/Y 0.03fF
C24769 NAND2X1_LOC_498/Y INVX1_LOC_361/Y 0.07fF
C24770 NAND2X1_LOC_500/a_36_24# INVX1_LOC_362/Y 0.00fF
C24771 NAND2X1_LOC_545/B INVX1_LOC_53/Y 0.08fF
C24772 INVX1_LOC_166/A INVX1_LOC_216/Y 0.01fF
C24773 INVX1_LOC_586/A INVX1_LOC_681/Y 0.02fF
C24774 INVX1_LOC_255/Y INVX1_LOC_93/Y 0.03fF
C24775 INVX1_LOC_409/A INVX1_LOC_63/Y 0.01fF
C24776 VDD INVX1_LOC_501/A 0.48fF
C24777 INVX1_LOC_614/A NAND2X1_LOC_677/Y 0.00fF
C24778 INVX1_LOC_395/A INVX1_LOC_555/A 0.03fF
C24779 INVX1_LOC_384/A NAND2X1_LOC_649/a_36_24# 0.00fF
C24780 NAND2X1_LOC_55/a_36_24# INVX1_LOC_62/Y 0.00fF
C24781 VDD INVX1_LOC_179/Y 0.42fF
C24782 INVX1_LOC_586/A INPUT_1 0.17fF
C24783 INVX1_LOC_384/A INVX1_LOC_48/Y 0.07fF
C24784 INVX1_LOC_617/A INVX1_LOC_11/Y 0.02fF
C24785 NAND2X1_LOC_750/Y INVX1_LOC_44/Y 0.08fF
C24786 INVX1_LOC_551/Y NAND2X1_LOC_775/B 0.23fF
C24787 INVX1_LOC_315/Y INVX1_LOC_31/Y 0.03fF
C24788 INVX1_LOC_20/Y NAND2X1_LOC_720/A 0.03fF
C24789 NAND2X1_LOC_843/A INVX1_LOC_655/Y 0.16fF
C24790 INVX1_LOC_442/A NAND2X1_LOC_388/A 0.00fF
C24791 INVX1_LOC_300/A INVX1_LOC_320/A 0.00fF
C24792 INVX1_LOC_146/A INVX1_LOC_50/Y 0.01fF
C24793 INVX1_LOC_301/A INVX1_LOC_100/Y 0.07fF
C24794 INPUT_0 NAND2X1_LOC_615/Y 0.04fF
C24795 INVX1_LOC_53/Y INVX1_LOC_98/Y 0.70fF
C24796 INVX1_LOC_512/A INVX1_LOC_463/Y 0.11fF
C24797 INVX1_LOC_285/Y INVX1_LOC_292/A 0.16fF
C24798 INVX1_LOC_21/Y INVX1_LOC_284/A 0.01fF
C24799 NAND2X1_LOC_241/B INVX1_LOC_44/Y 0.06fF
C24800 NAND2X1_LOC_333/a_36_24# INVX1_LOC_51/Y 0.01fF
C24801 INVX1_LOC_632/A INVX1_LOC_145/Y 0.07fF
C24802 INVX1_LOC_510/Y INVX1_LOC_89/Y 0.18fF
C24803 INVX1_LOC_441/Y INVX1_LOC_255/A 0.05fF
C24804 NAND2X1_LOC_475/A NAND2X1_LOC_494/a_36_24# 0.00fF
C24805 INVX1_LOC_12/Y INVX1_LOC_178/A 0.08fF
C24806 INVX1_LOC_312/Y INVX1_LOC_681/Y 0.00fF
C24807 INVX1_LOC_361/Y INVX1_LOC_377/Y 0.01fF
C24808 INVX1_LOC_255/Y INVX1_LOC_675/A 0.04fF
C24809 INVX1_LOC_134/A INVX1_LOC_69/Y 0.01fF
C24810 NAND2X1_LOC_537/A INVX1_LOC_531/Y 0.07fF
C24811 INVX1_LOC_410/A INVX1_LOC_45/Y 0.01fF
C24812 INVX1_LOC_317/Y INVX1_LOC_361/A 0.03fF
C24813 INVX1_LOC_114/Y INVX1_LOC_261/Y 0.00fF
C24814 INVX1_LOC_115/A INVX1_LOC_115/Y 0.02fF
C24815 INVX1_LOC_312/Y INPUT_1 0.03fF
C24816 INVX1_LOC_522/Y INVX1_LOC_46/Y 0.03fF
C24817 INVX1_LOC_170/Y INVX1_LOC_45/Y 0.01fF
C24818 INVX1_LOC_448/A NAND2X1_LOC_649/a_36_24# 0.00fF
C24819 INVX1_LOC_301/A INVX1_LOC_74/Y 0.01fF
C24820 INVX1_LOC_604/Y INVX1_LOC_209/A 0.02fF
C24821 NAND2X1_LOC_475/A INVX1_LOC_319/A 0.27fF
C24822 INVX1_LOC_213/Y NAND2X1_LOC_253/a_36_24# 0.00fF
C24823 INVX1_LOC_35/Y INVX1_LOC_7/Y 0.13fF
C24824 INVX1_LOC_202/A INVX1_LOC_211/A 0.04fF
C24825 INVX1_LOC_17/Y INVX1_LOC_504/Y 0.02fF
C24826 VDD NAND2X1_LOC_544/B 0.37fF
C24827 INVX1_LOC_352/Y INVX1_LOC_506/Y 0.05fF
C24828 INVX1_LOC_288/A NAND2X1_LOC_434/B 0.03fF
C24829 INVX1_LOC_399/Y INVX1_LOC_45/Y 0.03fF
C24830 INVX1_LOC_93/Y INVX1_LOC_474/Y 0.01fF
C24831 INVX1_LOC_349/Y INVX1_LOC_350/A 0.14fF
C24832 INVX1_LOC_172/Y INVX1_LOC_63/Y 0.01fF
C24833 INVX1_LOC_145/Y INVX1_LOC_48/Y 3.18fF
C24834 INVX1_LOC_99/Y NAND2X1_LOC_333/B 0.07fF
C24835 INVX1_LOC_51/A INVX1_LOC_347/A 0.06fF
C24836 INVX1_LOC_21/Y INVX1_LOC_31/Y 5.29fF
C24837 INVX1_LOC_559/Y NAND2X1_LOC_123/A 0.52fF
C24838 INVX1_LOC_534/Y INVX1_LOC_515/A 0.01fF
C24839 INVX1_LOC_120/Y INVX1_LOC_686/A 0.00fF
C24840 INVX1_LOC_442/Y INVX1_LOC_421/A 0.02fF
C24841 NAND2X1_LOC_505/Y INVX1_LOC_41/Y 0.05fF
C24842 INVX1_LOC_379/A INVX1_LOC_32/Y 0.07fF
C24843 NAND2X1_LOC_843/A INVX1_LOC_277/A 0.01fF
C24844 NAND2X1_LOC_250/Y NAND2X1_LOC_343/a_36_24# 0.00fF
C24845 INVX1_LOC_53/Y INVX1_LOC_338/Y 0.03fF
C24846 INVX1_LOC_31/Y NAND2X1_LOC_655/a_36_24# 0.00fF
C24847 INVX1_LOC_93/Y INVX1_LOC_481/Y 0.01fF
C24848 NAND2X1_LOC_383/Y INVX1_LOC_90/Y 0.10fF
C24849 INVX1_LOC_567/A INVX1_LOC_92/A 0.10fF
C24850 INVX1_LOC_32/Y INVX1_LOC_35/Y 1.96fF
C24851 INVX1_LOC_662/A INVX1_LOC_668/A 0.06fF
C24852 NAND2X1_LOC_125/a_36_24# INVX1_LOC_99/Y 0.01fF
C24853 INVX1_LOC_89/Y INVX1_LOC_116/A 0.03fF
C24854 INVX1_LOC_12/Y INVX1_LOC_58/Y 0.74fF
C24855 NAND2X1_LOC_318/B INVX1_LOC_199/Y 0.02fF
C24856 INVX1_LOC_566/A INVX1_LOC_242/Y 0.03fF
C24857 INVX1_LOC_261/Y INVX1_LOC_99/Y 0.03fF
C24858 INVX1_LOC_51/Y INVX1_LOC_41/Y 0.10fF
C24859 INVX1_LOC_26/Y INVX1_LOC_59/A 0.03fF
C24860 INVX1_LOC_117/Y NAND2X1_LOC_615/B 0.03fF
C24861 INVX1_LOC_555/A INVX1_LOC_189/Y 0.02fF
C24862 NAND2X1_LOC_253/Y NAND2X1_LOC_259/A 0.01fF
C24863 INVX1_LOC_20/Y INVX1_LOC_100/Y 1.53fF
C24864 INVX1_LOC_158/Y INVX1_LOC_89/Y 0.04fF
C24865 INVX1_LOC_89/Y INVX1_LOC_509/A 0.01fF
C24866 INVX1_LOC_630/A NAND2X1_LOC_800/B 0.45fF
C24867 INVX1_LOC_381/A NAND2X1_LOC_269/B 0.01fF
C24868 INVX1_LOC_367/A INVX1_LOC_26/Y 0.03fF
C24869 NAND2X1_LOC_707/A NAND2X1_LOC_691/A 0.07fF
C24870 INVX1_LOC_358/A NAND2X1_LOC_452/a_36_24# 0.00fF
C24871 INVX1_LOC_175/Y INVX1_LOC_100/Y 0.05fF
C24872 INVX1_LOC_327/Y INVX1_LOC_328/A 0.03fF
C24873 NAND2X1_LOC_520/A NAND2X1_LOC_275/Y 0.01fF
C24874 INVX1_LOC_84/Y INVX1_LOC_83/Y 1.11fF
C24875 INVX1_LOC_549/Y INVX1_LOC_496/A 0.02fF
C24876 INVX1_LOC_537/A INVX1_LOC_356/Y 0.01fF
C24877 INVX1_LOC_44/A INVX1_LOC_44/Y 0.04fF
C24878 INVX1_LOC_31/Y NAND2X1_LOC_267/A 0.08fF
C24879 INVX1_LOC_266/A INVX1_LOC_41/Y 0.13fF
C24880 INVX1_LOC_612/Y INVX1_LOC_6/Y 0.00fF
C24881 INVX1_LOC_35/Y NAND2X1_LOC_286/A 0.01fF
C24882 INVX1_LOC_452/A GATE_479 0.01fF
C24883 INVX1_LOC_297/A INVX1_LOC_369/Y 0.00fF
C24884 INVX1_LOC_32/Y NAND2X1_LOC_448/B 0.01fF
C24885 INVX1_LOC_20/Y INVX1_LOC_74/Y 0.13fF
C24886 INVX1_LOC_117/Y INVX1_LOC_66/A 0.26fF
C24887 INVX1_LOC_63/Y INVX1_LOC_352/Y 0.04fF
C24888 INVX1_LOC_103/Y INVX1_LOC_89/Y 0.23fF
C24889 INVX1_LOC_68/Y NAND2X1_LOC_231/B 0.01fF
C24890 INVX1_LOC_361/Y INVX1_LOC_47/Y 1.09fF
C24891 INVX1_LOC_69/Y INVX1_LOC_50/Y 1.79fF
C24892 INVX1_LOC_62/Y INVX1_LOC_492/Y 0.00fF
C24893 INVX1_LOC_365/Y INVX1_LOC_41/Y 0.01fF
C24894 INVX1_LOC_117/Y INVX1_LOC_296/A 0.02fF
C24895 INVX1_LOC_639/Y INVX1_LOC_632/Y 0.09fF
C24896 INVX1_LOC_662/A INVX1_LOC_668/Y 0.05fF
C24897 NAND2X1_LOC_333/A INVX1_LOC_157/A 0.04fF
C24898 NAND2X1_LOC_106/Y INVX1_LOC_6/Y 0.11fF
C24899 INVX1_LOC_63/Y INVX1_LOC_345/A 0.00fF
C24900 INVX1_LOC_366/Y INVX1_LOC_85/A 0.01fF
C24901 INVX1_LOC_514/A INVX1_LOC_168/Y 0.09fF
C24902 INVX1_LOC_76/Y INVX1_LOC_488/Y 0.02fF
C24903 INVX1_LOC_300/A INVX1_LOC_100/Y 0.10fF
C24904 INVX1_LOC_134/Y INVX1_LOC_653/Y 0.04fF
C24905 INVX1_LOC_508/A INVX1_LOC_46/Y 0.00fF
C24906 INVX1_LOC_254/Y INVX1_LOC_245/A 0.02fF
C24907 INVX1_LOC_47/Y INVX1_LOC_261/Y 0.03fF
C24908 INVX1_LOC_392/A INVX1_LOC_26/Y 0.13fF
C24909 INVX1_LOC_134/Y INVX1_LOC_666/Y 0.07fF
C24910 NAND2X1_LOC_388/A INVX1_LOC_255/A 0.03fF
C24911 INVX1_LOC_681/A INVX1_LOC_62/Y 0.00fF
C24912 INVX1_LOC_663/Y INVX1_LOC_100/Y 0.01fF
C24913 INVX1_LOC_376/Y NAND2X1_LOC_469/a_36_24# 0.00fF
C24914 INVX1_LOC_361/Y INVX1_LOC_119/Y 0.20fF
C24915 INVX1_LOC_598/A INVX1_LOC_79/A 0.01fF
C24916 INVX1_LOC_300/A INVX1_LOC_74/Y 0.13fF
C24917 INVX1_LOC_93/Y INVX1_LOC_128/Y 0.03fF
C24918 INVX1_LOC_41/Y INVX1_LOC_40/Y 0.03fF
C24919 INVX1_LOC_49/Y NAND2X1_LOC_686/B 0.20fF
C24920 INVX1_LOC_93/Y INVX1_LOC_26/Y 1.84fF
C24921 INVX1_LOC_74/Y INVX1_LOC_197/Y 0.01fF
C24922 INVX1_LOC_662/A INVX1_LOC_476/A 0.03fF
C24923 NAND2X1_LOC_106/B NAND2X1_LOC_248/B 0.02fF
C24924 INVX1_LOC_293/A INVX1_LOC_664/A 0.03fF
C24925 INVX1_LOC_340/A INVX1_LOC_454/Y 0.01fF
C24926 NAND2X1_LOC_482/Y INVX1_LOC_62/Y 0.24fF
C24927 INVX1_LOC_507/A INVX1_LOC_491/A 0.05fF
C24928 NAND2X1_LOC_866/a_36_24# INVX1_LOC_479/A 0.01fF
C24929 INVX1_LOC_642/Y INVX1_LOC_223/Y 0.04fF
C24930 INVX1_LOC_675/A INVX1_LOC_26/Y 0.07fF
C24931 INVX1_LOC_65/A NAND2X1_LOC_545/A 0.12fF
C24932 INVX1_LOC_476/Y INVX1_LOC_614/Y 0.09fF
C24933 INVX1_LOC_212/Y INVX1_LOC_669/A 0.03fF
C24934 INVX1_LOC_376/A INVX1_LOC_114/A 0.07fF
C24935 NAND2X1_LOC_689/B INVX1_LOC_479/A 0.03fF
C24936 INVX1_LOC_117/Y NAND2X1_LOC_646/B 0.05fF
C24937 NAND2X1_LOC_558/B INVX1_LOC_242/Y 0.04fF
C24938 NAND2X1_LOC_750/Y NAND2X1_LOC_58/a_36_24# 0.00fF
C24939 INVX1_LOC_543/A INVX1_LOC_26/Y 0.01fF
C24940 VDD INVX1_LOC_203/Y 0.54fF
C24941 VDD NAND2X1_LOC_780/B 0.05fF
C24942 INVX1_LOC_148/Y INVX1_LOC_496/A 0.02fF
C24943 INVX1_LOC_62/Y INVX1_LOC_168/Y 0.15fF
C24944 INVX1_LOC_79/A INVX1_LOC_242/Y 0.34fF
C24945 INVX1_LOC_100/Y INVX1_LOC_655/A 0.18fF
C24946 INVX1_LOC_528/Y NAND2X1_LOC_668/Y 0.11fF
C24947 INVX1_LOC_69/Y INVX1_LOC_658/Y 0.03fF
C24948 INVX1_LOC_6/Y INVX1_LOC_485/A 0.01fF
C24949 NAND2X1_LOC_615/Y INVX1_LOC_211/A 0.01fF
C24950 INVX1_LOC_79/A INVX1_LOC_487/A 0.00fF
C24951 INVX1_LOC_58/Y INVX1_LOC_212/A 0.01fF
C24952 INVX1_LOC_479/A INVX1_LOC_245/A 0.26fF
C24953 INVX1_LOC_224/Y INVX1_LOC_390/Y 0.04fF
C24954 INVX1_LOC_6/Y INVX1_LOC_92/A 0.06fF
C24955 NAND2X1_LOC_331/A INVX1_LOC_549/A 0.00fF
C24956 NAND2X1_LOC_710/B INVX1_LOC_395/A 0.02fF
C24957 INVX1_LOC_409/A INVX1_LOC_374/A 0.27fF
C24958 INVX1_LOC_210/A NAND2X1_LOC_243/a_36_24# 0.00fF
C24959 VDD INVX1_LOC_512/Y 0.14fF
C24960 INVX1_LOC_413/Y INVX1_LOC_217/Y 0.08fF
C24961 INVX1_LOC_26/Y INVX1_LOC_86/A 0.10fF
C24962 INVX1_LOC_400/Y INVX1_LOC_412/A 0.42fF
C24963 INPUT_0 INVX1_LOC_340/Y 2.98fF
C24964 INVX1_LOC_441/A INVX1_LOC_347/A -0.08fF
C24965 INVX1_LOC_206/Y INVX1_LOC_396/Y 0.12fF
C24966 NAND2X1_LOC_249/Y INVX1_LOC_367/A 0.07fF
C24967 INVX1_LOC_409/Y INVX1_LOC_80/A 0.01fF
C24968 NAND2X1_LOC_322/Y INVX1_LOC_80/A 0.01fF
C24969 NAND2X1_LOC_65/a_36_24# INPUT_0 0.00fF
C24970 NAND2X1_LOC_503/B INVX1_LOC_603/Y 0.02fF
C24971 NAND2X1_LOC_735/a_36_24# INVX1_LOC_51/Y 0.00fF
C24972 INVX1_LOC_551/Y NAND2X1_LOC_317/B 0.01fF
C24973 NAND2X1_LOC_526/a_36_24# INVX1_LOC_362/Y 0.00fF
C24974 INVX1_LOC_206/Y INVX1_LOC_686/A 0.54fF
C24975 INVX1_LOC_425/A NAND2X1_LOC_552/a_36_24# 0.00fF
C24976 INVX1_LOC_412/Y INVX1_LOC_197/A 0.03fF
C24977 INVX1_LOC_134/A INVX1_LOC_586/A 0.01fF
C24978 VDD INVX1_LOC_205/Y 0.42fF
C24979 INVX1_LOC_287/Y INVX1_LOC_271/A 0.10fF
C24980 NAND2X1_LOC_710/A NAND2X1_LOC_516/Y 0.02fF
C24981 INVX1_LOC_11/Y INVX1_LOC_409/Y 0.03fF
C24982 INVX1_LOC_454/A INVX1_LOC_25/Y 0.03fF
C24983 INVX1_LOC_400/Y NAND2X1_LOC_336/B 0.03fF
C24984 INVX1_LOC_434/A INVX1_LOC_386/Y 0.03fF
C24985 NAND2X1_LOC_45/Y INVX1_LOC_442/Y 0.10fF
C24986 NAND2X1_LOC_123/a_36_24# INVX1_LOC_638/A 0.01fF
C24987 INVX1_LOC_395/A INVX1_LOC_474/Y 0.05fF
C24988 NAND2X1_LOC_61/A INVX1_LOC_54/Y 0.13fF
C24989 INVX1_LOC_435/Y INVX1_LOC_53/Y 1.39fF
C24990 NAND2X1_LOC_45/Y NAND2X1_LOC_692/Y 0.04fF
C24991 VDD INVX1_LOC_194/Y 1.61fF
C24992 INVX1_LOC_614/A INVX1_LOC_137/A 0.04fF
C24993 INVX1_LOC_561/Y INVX1_LOC_145/Y 0.03fF
C24994 NAND2X1_LOC_554/a_36_24# INVX1_LOC_54/Y 0.06fF
C24995 INVX1_LOC_20/Y INVX1_LOC_566/A 0.12fF
C24996 INVX1_LOC_445/Y INVX1_LOC_442/Y 0.05fF
C24997 NAND2X1_LOC_332/B NAND2X1_LOC_139/a_36_24# 0.00fF
C24998 INVX1_LOC_68/Y INVX1_LOC_80/A 0.04fF
C24999 NAND2X1_LOC_122/Y INVX1_LOC_188/Y 0.03fF
C25000 INVX1_LOC_224/Y INVX1_LOC_432/A 0.00fF
C25001 NAND2X1_LOC_249/Y INVX1_LOC_93/Y 0.03fF
C25002 INVX1_LOC_69/Y INVX1_LOC_275/A 0.03fF
C25003 INVX1_LOC_118/Y INVX1_LOC_371/A 0.01fF
C25004 NAND2X1_LOC_218/a_36_24# INVX1_LOC_194/A 0.02fF
C25005 INVX1_LOC_638/Y INVX1_LOC_638/A 0.03fF
C25006 INVX1_LOC_21/Y INVX1_LOC_51/Y 0.18fF
C25007 INVX1_LOC_603/Y INVX1_LOC_273/A 0.01fF
C25008 INVX1_LOC_54/Y NAND2X1_LOC_378/a_36_24# 0.00fF
C25009 INVX1_LOC_286/A INVX1_LOC_155/Y 0.01fF
C25010 NAND2X1_LOC_520/B INVX1_LOC_367/Y 0.08fF
C25011 INVX1_LOC_447/Y INVX1_LOC_45/Y 0.09fF
C25012 INVX1_LOC_459/Y INVX1_LOC_504/A 0.01fF
C25013 INVX1_LOC_207/A INVX1_LOC_197/Y 0.00fF
C25014 NAND2X1_LOC_707/A INVX1_LOC_537/A 0.07fF
C25015 INVX1_LOC_374/A INVX1_LOC_352/Y 0.00fF
C25016 NAND2X1_LOC_759/B NAND2X1_LOC_759/Y 0.12fF
C25017 INVX1_LOC_76/Y INVX1_LOC_115/Y 0.00fF
C25018 INVX1_LOC_408/Y INVX1_LOC_117/Y 0.04fF
C25019 INVX1_LOC_418/A NAND2X1_LOC_775/B 0.01fF
C25020 INVX1_LOC_199/Y NAND2X1_LOC_76/B 0.31fF
C25021 INVX1_LOC_374/A INVX1_LOC_345/A 0.02fF
C25022 INVX1_LOC_266/Y INVX1_LOC_479/Y 0.05fF
C25023 INVX1_LOC_68/Y INVX1_LOC_11/Y 0.00fF
C25024 INVX1_LOC_54/Y INVX1_LOC_185/Y 0.03fF
C25025 VDD INVX1_LOC_44/Y 3.06fF
C25026 INVX1_LOC_564/Y INVX1_LOC_93/Y 0.13fF
C25027 INVX1_LOC_316/Y INVX1_LOC_55/Y 0.37fF
C25028 INVX1_LOC_300/A INVX1_LOC_566/A 0.01fF
C25029 INVX1_LOC_442/A NAND2X1_LOC_112/a_36_24# 0.00fF
C25030 INVX1_LOC_606/Y INVX1_LOC_523/Y 0.03fF
C25031 INVX1_LOC_54/Y INVX1_LOC_45/Y 0.29fF
C25032 INVX1_LOC_405/A INVX1_LOC_405/Y 0.02fF
C25033 NAND2X1_LOC_526/Y NAND2X1_LOC_184/Y 0.01fF
C25034 INVX1_LOC_80/A INVX1_LOC_600/A 0.18fF
C25035 INVX1_LOC_21/Y INVX1_LOC_365/Y 0.01fF
C25036 INVX1_LOC_677/Y INVX1_LOC_685/Y 0.32fF
C25037 NAND2X1_LOC_130/Y INVX1_LOC_80/A 0.03fF
C25038 INVX1_LOC_586/A INVX1_LOC_50/Y 0.19fF
C25039 INVX1_LOC_435/A INVX1_LOC_235/Y 0.03fF
C25040 INVX1_LOC_206/Y NAND2X1_LOC_334/A 8.84fF
C25041 INVX1_LOC_516/Y INVX1_LOC_50/Y 0.01fF
C25042 INVX1_LOC_53/Y INVX1_LOC_504/A 0.07fF
C25043 INVX1_LOC_550/Y INVX1_LOC_522/Y 0.05fF
C25044 INVX1_LOC_340/Y INVX1_LOC_498/A 0.02fF
C25045 VDD INVX1_LOC_48/A -0.00fF
C25046 INVX1_LOC_435/A NAND2X1_LOC_361/a_36_24# 0.01fF
C25047 INVX1_LOC_578/A NAND2X1_LOC_542/A 0.03fF
C25048 INVX1_LOC_604/A INVX1_LOC_58/Y 0.01fF
C25049 INVX1_LOC_301/A INVX1_LOC_79/A 0.03fF
C25050 INVX1_LOC_577/Y INVX1_LOC_31/Y 0.03fF
C25051 NAND2X1_LOC_707/A INVX1_LOC_496/Y 0.06fF
C25052 NAND2X1_LOC_373/Y INVX1_LOC_100/Y 0.63fF
C25053 INVX1_LOC_441/Y INVX1_LOC_69/Y 0.01fF
C25054 INVX1_LOC_228/Y INVX1_LOC_44/Y 0.07fF
C25055 VDD INVX1_LOC_461/Y 0.21fF
C25056 NAND2X1_LOC_123/A INVX1_LOC_155/Y 0.01fF
C25057 INVX1_LOC_438/A INVX1_LOC_247/Y 0.03fF
C25058 INPUT_3 INVX1_LOC_54/Y 0.06fF
C25059 INVX1_LOC_550/A INVX1_LOC_522/Y 0.02fF
C25060 INVX1_LOC_20/Y INVX1_LOC_469/Y 0.04fF
C25061 INVX1_LOC_266/A NAND2X1_LOC_267/A 0.14fF
C25062 INVX1_LOC_560/A INVX1_LOC_390/A 0.02fF
C25063 NAND2X1_LOC_440/a_36_24# INVX1_LOC_50/Y 0.00fF
C25064 INVX1_LOC_442/Y INVX1_LOC_99/Y 0.07fF
C25065 INVX1_LOC_522/A INVX1_LOC_511/A 0.18fF
C25066 INVX1_LOC_117/Y INVX1_LOC_196/A 0.04fF
C25067 INVX1_LOC_312/Y INVX1_LOC_50/Y 0.03fF
C25068 INPUT_1 INVX1_LOC_486/Y 2.84fF
C25069 INVX1_LOC_11/Y INVX1_LOC_600/A 0.03fF
C25070 INVX1_LOC_11/Y NAND2X1_LOC_130/Y 0.04fF
C25071 NAND2X1_LOC_460/A INVX1_LOC_48/Y 0.40fF
C25072 NAND2X1_LOC_457/A INVX1_LOC_502/A 0.12fF
C25073 INVX1_LOC_167/A INVX1_LOC_633/Y 0.00fF
C25074 NAND2X1_LOC_596/Y INVX1_LOC_461/Y 0.08fF
C25075 INVX1_LOC_557/A INVX1_LOC_376/Y 0.09fF
C25076 INVX1_LOC_395/A INVX1_LOC_26/Y 0.20fF
C25077 INVX1_LOC_335/Y INVX1_LOC_40/Y 0.03fF
C25078 INVX1_LOC_17/Y INVX1_LOC_453/Y 0.03fF
C25079 INVX1_LOC_517/Y INVX1_LOC_516/Y 0.09fF
C25080 INVX1_LOC_527/Y INVX1_LOC_155/Y 0.01fF
C25081 INVX1_LOC_272/Y INVX1_LOC_292/Y 0.00fF
C25082 NAND2X1_LOC_791/B INVX1_LOC_292/Y 0.13fF
C25083 NAND2X1_LOC_775/a_36_24# INVX1_LOC_603/A 0.02fF
C25084 INVX1_LOC_129/A INVX1_LOC_159/Y 0.02fF
C25085 NAND2X1_LOC_520/A INVX1_LOC_235/Y 0.12fF
C25086 INVX1_LOC_206/Y NAND2X1_LOC_609/B 2.23fF
C25087 INVX1_LOC_117/Y INVX1_LOC_305/Y 0.01fF
C25088 INVX1_LOC_85/Y INVX1_LOC_183/Y 0.14fF
C25089 INVX1_LOC_17/Y INVX1_LOC_259/Y 0.03fF
C25090 INVX1_LOC_76/Y INVX1_LOC_507/Y 0.03fF
C25091 INVX1_LOC_504/A INVX1_LOC_460/Y 0.01fF
C25092 NAND2X1_LOC_543/B INVX1_LOC_625/Y 0.01fF
C25093 INVX1_LOC_522/A NAND2X1_LOC_679/B 0.01fF
C25094 INVX1_LOC_362/Y INVX1_LOC_26/Y 0.03fF
C25095 INVX1_LOC_54/Y NAND2X1_LOC_376/Y 0.02fF
C25096 INVX1_LOC_32/Y INVX1_LOC_531/A 0.01fF
C25097 NAND2X1_LOC_791/B INVX1_LOC_284/Y 0.28fF
C25098 INVX1_LOC_686/A NAND2X1_LOC_334/A 0.07fF
C25099 INVX1_LOC_367/A NAND2X1_LOC_280/a_36_24# 0.00fF
C25100 NAND2X1_LOC_112/a_36_24# INVX1_LOC_116/Y 0.01fF
C25101 INVX1_LOC_679/Y INVX1_LOC_6/Y 0.20fF
C25102 INVX1_LOC_41/Y INVX1_LOC_216/Y 0.01fF
C25103 NAND2X1_LOC_397/Y INVX1_LOC_46/Y 0.01fF
C25104 INVX1_LOC_47/Y INVX1_LOC_307/A 0.02fF
C25105 INVX1_LOC_137/Y INVX1_LOC_514/A 0.03fF
C25106 NAND2X1_LOC_615/B NAND2X1_LOC_76/A 0.04fF
C25107 NAND2X1_LOC_415/B INVX1_LOC_46/Y 0.04fF
C25108 INVX1_LOC_20/Y NAND2X1_LOC_558/B 0.01fF
C25109 INVX1_LOC_372/Y NAND2X1_LOC_440/A 0.01fF
C25110 INVX1_LOC_449/A INVX1_LOC_63/Y 0.07fF
C25111 INVX1_LOC_195/Y INVX1_LOC_86/Y 0.01fF
C25112 INVX1_LOC_442/Y INVX1_LOC_47/Y 0.07fF
C25113 NAND2X1_LOC_525/Y NAND2X1_LOC_844/A 0.16fF
C25114 NAND2X1_LOC_321/a_36_24# INVX1_LOC_376/A 0.00fF
C25115 NAND2X1_LOC_775/B INVX1_LOC_46/Y 0.08fF
C25116 INVX1_LOC_20/Y INVX1_LOC_79/A 0.14fF
C25117 INVX1_LOC_625/A INVX1_LOC_199/Y 0.53fF
C25118 INVX1_LOC_45/Y INVX1_LOC_388/A 0.01fF
C25119 INVX1_LOC_519/Y INVX1_LOC_126/Y 0.02fF
C25120 INVX1_LOC_492/A INVX1_LOC_477/Y 0.01fF
C25121 INVX1_LOC_619/A INVX1_LOC_179/Y 0.03fF
C25122 INVX1_LOC_153/A NAND2X1_LOC_333/B 0.02fF
C25123 NAND2X1_LOC_13/Y INVX1_LOC_41/Y 0.01fF
C25124 INVX1_LOC_514/A NAND2X1_LOC_829/B 0.00fF
C25125 INVX1_LOC_221/Y INVX1_LOC_671/Y 0.25fF
C25126 INVX1_LOC_167/Y INVX1_LOC_62/Y 0.01fF
C25127 INVX1_LOC_455/A NAND2X1_LOC_836/B 0.00fF
C25128 INVX1_LOC_12/Y INVX1_LOC_245/A 0.05fF
C25129 INVX1_LOC_11/Y NAND2X1_LOC_613/a_36_24# 0.00fF
C25130 INVX1_LOC_145/Y NAND2X1_LOC_615/Y 0.07fF
C25131 INVX1_LOC_670/Y INVX1_LOC_518/A 0.02fF
C25132 INVX1_LOC_105/A INVX1_LOC_89/Y 0.02fF
C25133 INVX1_LOC_6/Y INPUT_1 0.37fF
C25134 INVX1_LOC_369/A NAND2X1_LOC_624/a_36_24# 0.00fF
C25135 INVX1_LOC_417/Y INVX1_LOC_242/Y 0.83fF
C25136 INVX1_LOC_459/Y INVX1_LOC_346/Y 0.19fF
C25137 INVX1_LOC_209/A INVX1_LOC_63/Y 0.01fF
C25138 NAND2X1_LOC_837/B NAND2X1_LOC_838/a_36_24# 0.00fF
C25139 INVX1_LOC_468/Y INVX1_LOC_376/Y 0.09fF
C25140 INVX1_LOC_284/A INVX1_LOC_26/Y 0.08fF
C25141 INVX1_LOC_21/Y INVX1_LOC_204/A 0.01fF
C25142 INVX1_LOC_99/Y INVX1_LOC_471/Y 0.01fF
C25143 INVX1_LOC_205/Y NAND2X1_LOC_786/B 0.01fF
C25144 NAND2X1_LOC_825/a_36_24# INVX1_LOC_50/Y 0.00fF
C25145 INVX1_LOC_300/A NAND2X1_LOC_558/B 0.01fF
C25146 INVX1_LOC_662/A INVX1_LOC_98/Y 0.45fF
C25147 INVX1_LOC_58/Y NAND2X1_LOC_615/B 0.01fF
C25148 INVX1_LOC_337/Y NAND2X1_LOC_410/Y 0.08fF
C25149 NAND2X1_LOC_128/A NAND2X1_LOC_127/a_36_24# 0.01fF
C25150 INVX1_LOC_204/Y INVX1_LOC_601/Y 0.03fF
C25151 NAND2X1_LOC_184/Y INVX1_LOC_654/Y 0.09fF
C25152 INVX1_LOC_17/Y INVX1_LOC_114/A 0.11fF
C25153 INVX1_LOC_300/A INVX1_LOC_79/A 0.27fF
C25154 INVX1_LOC_548/A INVX1_LOC_26/Y 0.01fF
C25155 INVX1_LOC_79/A INVX1_LOC_197/Y 5.35fF
C25156 NAND2X1_LOC_612/A INVX1_LOC_614/Y 0.03fF
C25157 NAND2X1_LOC_477/a_36_24# INVX1_LOC_510/A 0.01fF
C25158 INVX1_LOC_422/Y INVX1_LOC_6/Y 0.05fF
C25159 NAND2X1_LOC_388/A INVX1_LOC_69/Y 0.09fF
C25160 INVX1_LOC_16/Y INVX1_LOC_653/Y 0.01fF
C25161 INVX1_LOC_117/Y INVX1_LOC_179/A 0.54fF
C25162 INVX1_LOC_562/Y INVX1_LOC_636/A 0.03fF
C25163 INVX1_LOC_242/Y INVX1_LOC_48/Y 0.10fF
C25164 INVX1_LOC_674/Y INVX1_LOC_340/A 0.03fF
C25165 INVX1_LOC_58/Y INVX1_LOC_66/A 0.53fF
C25166 INVX1_LOC_199/Y NAND2X1_LOC_52/Y 0.03fF
C25167 INVX1_LOC_93/Y NAND2X1_LOC_605/B 0.04fF
C25168 INVX1_LOC_120/Y NAND2X1_LOC_542/A 0.15fF
C25169 NAND2X1_LOC_90/a_36_24# INVX1_LOC_66/A 0.00fF
C25170 NAND2X1_LOC_333/A INVX1_LOC_245/A 0.03fF
C25171 INVX1_LOC_534/Y NAND2X1_LOC_829/B 0.01fF
C25172 INVX1_LOC_137/Y INVX1_LOC_62/Y 0.07fF
C25173 INVX1_LOC_31/Y INVX1_LOC_26/Y 0.25fF
C25174 INVX1_LOC_48/Y INVX1_LOC_487/A 0.01fF
C25175 INVX1_LOC_93/Y NAND2X1_LOC_626/Y 0.04fF
C25176 INVX1_LOC_7/Y INVX1_LOC_488/Y 0.01fF
C25177 INVX1_LOC_188/A INVX1_LOC_245/A 0.01fF
C25178 INVX1_LOC_662/A INVX1_LOC_338/Y 0.02fF
C25179 NAND2X1_LOC_799/a_36_24# INVX1_LOC_638/A 0.01fF
C25180 INVX1_LOC_63/Y INVX1_LOC_328/Y 0.04fF
C25181 NAND2X1_LOC_836/B NAND2X1_LOC_823/Y 0.07fF
C25182 INVX1_LOC_394/Y VDD 0.21fF
C25183 NAND2X1_LOC_675/B INVX1_LOC_26/Y 0.06fF
C25184 INVX1_LOC_623/Y INVX1_LOC_597/Y 0.00fF
C25185 INVX1_LOC_44/Y NAND2X1_LOC_786/B 0.06fF
C25186 INVX1_LOC_460/Y INVX1_LOC_346/Y 0.52fF
C25187 INVX1_LOC_574/A INVX1_LOC_185/A 0.12fF
C25188 INVX1_LOC_41/Y INVX1_LOC_361/A 0.03fF
C25189 VDD NAND2X1_LOC_176/Y 0.01fF
C25190 INVX1_LOC_520/Y INVX1_LOC_479/A 0.01fF
C25191 INVX1_LOC_44/Y INVX1_LOC_635/Y 0.03fF
C25192 VDD INVX1_LOC_118/Y 0.71fF
C25193 INVX1_LOC_58/Y NAND2X1_LOC_621/B 0.02fF
C25194 INVX1_LOC_79/A NAND2X1_LOC_269/B 0.00fF
C25195 INVX1_LOC_58/Y NAND2X1_LOC_646/B 0.01fF
C25196 INVX1_LOC_26/Y INVX1_LOC_473/Y 0.10fF
C25197 NAND2X1_LOC_331/A INVX1_LOC_572/A 0.01fF
C25198 VDD INVX1_LOC_96/Y 0.21fF
C25199 NAND2X1_LOC_249/Y INVX1_LOC_362/Y 0.04fF
C25200 INVX1_LOC_647/Y INVX1_LOC_9/Y 0.01fF
C25201 INVX1_LOC_366/A INVX1_LOC_181/A 0.03fF
C25202 NAND2X1_LOC_274/B NAND2X1_LOC_497/a_36_24# 0.00fF
C25203 VDD NAND2X1_LOC_685/B 0.01fF
C25204 INVX1_LOC_666/Y INVX1_LOC_90/Y 0.03fF
C25205 INVX1_LOC_395/A INVX1_LOC_560/A 0.01fF
C25206 INVX1_LOC_206/Y INVX1_LOC_397/A 0.24fF
C25207 NAND2X1_LOC_790/B INVX1_LOC_524/Y 0.02fF
C25208 INVX1_LOC_353/A INVX1_LOC_91/Y 0.03fF
C25209 NAND2X1_LOC_666/Y INVX1_LOC_636/A 0.21fF
C25210 INVX1_LOC_438/A INVX1_LOC_586/A 0.33fF
C25211 INVX1_LOC_206/Y INVX1_LOC_94/A 0.01fF
C25212 NAND2X1_LOC_789/B INVX1_LOC_366/A 0.03fF
C25213 INVX1_LOC_557/A INVX1_LOC_253/A 0.03fF
C25214 NAND2X1_LOC_498/Y INVX1_LOC_618/Y 0.02fF
C25215 INVX1_LOC_150/A NAND2X1_LOC_685/A 0.01fF
C25216 INVX1_LOC_380/A INVX1_LOC_211/Y 0.01fF
C25217 NAND2X1_LOC_331/A INVX1_LOC_515/A 0.01fF
C25218 INVX1_LOC_531/Y INVX1_LOC_291/Y 0.03fF
C25219 INVX1_LOC_438/A INVX1_LOC_246/Y 0.04fF
C25220 VDD NAND2X1_LOC_391/A 0.41fF
C25221 INVX1_LOC_255/Y INVX1_LOC_51/Y 0.04fF
C25222 INVX1_LOC_335/Y INVX1_LOC_463/A 0.07fF
C25223 INVX1_LOC_441/Y INVX1_LOC_586/A 0.01fF
C25224 INVX1_LOC_257/Y INVX1_LOC_634/A 0.01fF
C25225 NAND2X1_LOC_69/B INVX1_LOC_145/Y 0.08fF
C25226 INVX1_LOC_438/A INVX1_LOC_312/Y 0.06fF
C25227 INVX1_LOC_224/Y INVX1_LOC_295/A 0.01fF
C25228 INVX1_LOC_288/A INVX1_LOC_340/Y 0.05fF
C25229 VDD INVX1_LOC_147/A -0.00fF
C25230 NAND2X1_LOC_526/Y NAND2X1_LOC_486/B 0.16fF
C25231 VDD INVX1_LOC_27/Y 0.22fF
C25232 NAND2X1_LOC_790/B INVX1_LOC_400/A 0.02fF
C25233 VDD NAND2X1_LOC_418/Y 0.01fF
C25234 INVX1_LOC_577/Y INVX1_LOC_51/Y 0.01fF
C25235 VDD INVX1_LOC_610/A -0.00fF
C25236 INVX1_LOC_171/Y INVX1_LOC_45/Y 0.43fF
C25237 INVX1_LOC_434/A INVX1_LOC_7/Y 0.23fF
C25238 INVX1_LOC_395/A INVX1_LOC_369/A 0.05fF
C25239 INVX1_LOC_329/Y INVX1_LOC_636/A 0.03fF
C25240 VDD INVX1_LOC_656/Y 0.21fF
C25241 INVX1_LOC_76/Y INVX1_LOC_163/Y 0.04fF
C25242 INVX1_LOC_43/Y INVX1_LOC_190/Y 0.04fF
C25243 INVX1_LOC_567/A INVX1_LOC_50/Y 0.00fF
C25244 INVX1_LOC_301/A INVX1_LOC_48/Y 0.84fF
C25245 NAND2X1_LOC_790/B INVX1_LOC_93/Y 0.01fF
C25246 INVX1_LOC_577/A INVX1_LOC_300/A -0.09fF
C25247 INVX1_LOC_562/A NAND2X1_LOC_666/a_36_24# 0.01fF
C25248 INVX1_LOC_17/Y NAND2X1_LOC_457/A 0.08fF
C25249 INVX1_LOC_76/Y INVX1_LOC_522/Y 0.05fF
C25250 INPUT_3 INVX1_LOC_171/Y 0.03fF
C25251 INVX1_LOC_412/A INVX1_LOC_99/Y 0.02fF
C25252 INVX1_LOC_384/A NAND2X1_LOC_541/B 0.08fF
C25253 INVX1_LOC_608/Y INVX1_LOC_547/Y 0.05fF
C25254 NAND2X1_LOC_763/Y INVX1_LOC_623/Y 0.09fF
C25255 INVX1_LOC_95/Y INVX1_LOC_95/A 0.01fF
C25256 INVX1_LOC_445/Y INVX1_LOC_278/Y 0.01fF
C25257 INVX1_LOC_17/Y INVX1_LOC_547/Y 0.16fF
C25258 INVX1_LOC_6/Y INVX1_LOC_181/A 0.01fF
C25259 INVX1_LOC_384/A INVX1_LOC_383/Y 0.02fF
C25260 INVX1_LOC_202/Y INVX1_LOC_271/A 0.07fF
C25261 VDD INVX1_LOC_523/Y 0.23fF
C25262 NAND2X1_LOC_122/Y NAND2X1_LOC_421/a_36_24# 0.00fF
C25263 INVX1_LOC_510/Y NAND2X1_LOC_418/Y 0.01fF
C25264 NAND2X1_LOC_130/a_36_24# INVX1_LOC_361/Y 0.00fF
C25265 INVX1_LOC_307/Y INVX1_LOC_46/Y 0.10fF
C25266 INVX1_LOC_435/Y INVX1_LOC_213/Y 0.05fF
C25267 INVX1_LOC_33/Y INVX1_LOC_6/A 0.09fF
C25268 INVX1_LOC_398/A NAND2X1_LOC_237/Y 0.01fF
C25269 NAND2X1_LOC_271/B INVX1_LOC_46/Y 0.06fF
C25270 INVX1_LOC_442/Y INVX1_LOC_502/Y 0.00fF
C25271 NAND2X1_LOC_35/a_36_24# INVX1_LOC_366/A -0.01fF
C25272 INVX1_LOC_140/Y INVX1_LOC_50/Y 0.03fF
C25273 INVX1_LOC_87/A NAND2X1_LOC_749/Y 0.09fF
C25274 NAND2X1_LOC_493/B INVX1_LOC_99/Y 0.02fF
C25275 INVX1_LOC_446/A INVX1_LOC_328/Y 0.02fF
C25276 NAND2X1_LOC_542/a_36_24# INVX1_LOC_686/A 0.00fF
C25277 NAND2X1_LOC_789/B INVX1_LOC_6/Y 0.00fF
C25278 INVX1_LOC_17/Y INVX1_LOC_482/A 0.10fF
C25279 INVX1_LOC_560/A INVX1_LOC_31/Y 0.14fF
C25280 NAND2X1_LOC_788/A INVX1_LOC_58/Y 0.01fF
C25281 NAND2X1_LOC_250/Y INVX1_LOC_651/Y -0.00fF
C25282 INVX1_LOC_206/Y NAND2X1_LOC_542/A 0.05fF
C25283 NAND2X1_LOC_32/a_36_24# INVX1_LOC_54/Y 0.00fF
C25284 INVX1_LOC_20/Y INVX1_LOC_59/Y 0.05fF
C25285 NAND2X1_LOC_391/B INVX1_LOC_304/Y 0.00fF
C25286 INVX1_LOC_76/Y NAND2X1_LOC_606/Y 0.05fF
C25287 NAND2X1_LOC_507/A INVX1_LOC_45/Y 0.02fF
C25288 INVX1_LOC_324/A INVX1_LOC_7/Y 0.05fF
C25289 INVX1_LOC_386/Y INVX1_LOC_489/A 0.17fF
C25290 VDD INVX1_LOC_226/Y 0.26fF
C25291 NAND2X1_LOC_336/B INVX1_LOC_99/Y 0.31fF
C25292 INVX1_LOC_581/A NAND2X1_LOC_834/a_36_24# -0.02fF
C25293 INVX1_LOC_448/A INVX1_LOC_383/Y 0.01fF
C25294 INVX1_LOC_617/Y INVX1_LOC_510/A 0.00fF
C25295 INVX1_LOC_145/Y NAND2X1_LOC_541/B 0.11fF
C25296 NAND2X1_LOC_58/a_36_24# NAND2X1_LOC_786/B 0.00fF
C25297 NAND2X1_LOC_475/A INVX1_LOC_482/Y 0.00fF
C25298 INVX1_LOC_619/A INVX1_LOC_205/Y 0.03fF
C25299 INVX1_LOC_408/Y INVX1_LOC_58/Y 0.46fF
C25300 NAND2X1_LOC_509/a_36_24# INVX1_LOC_273/A 0.00fF
C25301 INVX1_LOC_20/Y INVX1_LOC_48/Y 0.64fF
C25302 INVX1_LOC_438/A INVX1_LOC_225/Y 0.03fF
C25303 INVX1_LOC_206/Y INVX1_LOC_376/Y 0.07fF
C25304 NAND2X1_LOC_331/A INVX1_LOC_168/Y 0.07fF
C25305 INVX1_LOC_117/Y INVX1_LOC_146/A 0.03fF
C25306 INVX1_LOC_89/Y INVX1_LOC_45/Y 0.14fF
C25307 NAND2X1_LOC_13/Y NAND2X1_LOC_267/A 0.29fF
C25308 INVX1_LOC_65/Y INVX1_LOC_199/Y 0.08fF
C25309 NAND2X1_LOC_388/A INVX1_LOC_586/A 0.11fF
C25310 INVX1_LOC_54/Y INVX1_LOC_293/Y 0.15fF
C25311 INVX1_LOC_166/A INVX1_LOC_551/Y 0.01fF
C25312 NAND2X1_LOC_791/B INVX1_LOC_50/Y 0.00fF
C25313 INVX1_LOC_169/A INVX1_LOC_46/Y 0.04fF
C25314 INVX1_LOC_93/Y INVX1_LOC_235/Y 0.07fF
C25315 INVX1_LOC_486/Y INVX1_LOC_50/Y 0.03fF
C25316 INVX1_LOC_442/A INVX1_LOC_58/Y 0.07fF
C25317 INVX1_LOC_47/Y NAND2X1_LOC_707/A 0.07fF
C25318 NAND2X1_LOC_712/a_36_24# INVX1_LOC_53/Y 0.00fF
C25319 INVX1_LOC_374/A INVX1_LOC_347/Y 0.00fF
C25320 INVX1_LOC_294/Y INVX1_LOC_50/Y 0.01fF
C25321 INVX1_LOC_270/A INVX1_LOC_317/A 0.01fF
C25322 INVX1_LOC_315/Y NAND2X1_LOC_668/Y 0.06fF
C25323 INVX1_LOC_337/Y INVX1_LOC_46/Y 0.08fF
C25324 NAND2X1_LOC_542/A INVX1_LOC_242/A 0.01fF
C25325 INVX1_LOC_266/Y INVX1_LOC_63/Y 0.10fF
C25326 NAND2X1_LOC_27/Y INVX1_LOC_12/Y 0.02fF
C25327 INVX1_LOC_300/A INVX1_LOC_59/Y 0.05fF
C25328 INVX1_LOC_451/A INVX1_LOC_451/Y 0.01fF
C25329 INVX1_LOC_45/Y INVX1_LOC_501/A 0.03fF
C25330 INVX1_LOC_59/Y INVX1_LOC_197/Y 0.03fF
C25331 INVX1_LOC_53/Y INVX1_LOC_520/A 0.01fF
C25332 INVX1_LOC_556/Y INVX1_LOC_669/Y 0.02fF
C25333 INVX1_LOC_31/Y INVX1_LOC_369/A 0.07fF
C25334 INVX1_LOC_662/Y NAND2X1_LOC_285/B 0.07fF
C25335 INVX1_LOC_105/Y INVX1_LOC_670/Y 0.01fF
C25336 NAND2X1_LOC_505/Y INVX1_LOC_26/Y 0.10fF
C25337 INVX1_LOC_614/A INVX1_LOC_523/Y 0.32fF
C25338 INVX1_LOC_20/Y NAND2X1_LOC_491/Y 0.01fF
C25339 INVX1_LOC_602/A INVX1_LOC_69/Y 2.84fF
C25340 INVX1_LOC_672/A INVX1_LOC_661/Y 0.29fF
C25341 INVX1_LOC_412/Y INVX1_LOC_66/Y 0.01fF
C25342 NAND2X1_LOC_775/B INVX1_LOC_349/Y -0.00fF
C25343 NAND2X1_LOC_16/Y INVX1_LOC_90/Y 0.01fF
C25344 INVX1_LOC_300/A INVX1_LOC_48/Y 1.37fF
C25345 INVX1_LOC_187/A INVX1_LOC_157/Y 0.12fF
C25346 INVX1_LOC_686/A NAND2X1_LOC_542/A 0.02fF
C25347 INVX1_LOC_662/Y NAND2X1_LOC_106/B 0.03fF
C25348 INVX1_LOC_452/A INVX1_LOC_282/A 0.11fF
C25349 INVX1_LOC_196/A INVX1_LOC_58/Y 0.01fF
C25350 INVX1_LOC_63/A NAND2X1_LOC_836/B 0.19fF
C25351 INVX1_LOC_51/Y INVX1_LOC_26/Y 0.19fF
C25352 INVX1_LOC_48/Y INVX1_LOC_197/Y 0.03fF
C25353 INVX1_LOC_376/Y INVX1_LOC_242/A 0.16fF
C25354 INVX1_LOC_613/Y INVX1_LOC_633/A 0.02fF
C25355 INVX1_LOC_69/Y INVX1_LOC_104/Y 0.01fF
C25356 NAND2X1_LOC_638/A INVX1_LOC_261/Y 0.08fF
C25357 INVX1_LOC_193/A INVX1_LOC_159/Y 0.00fF
C25358 INVX1_LOC_31/Y NAND2X1_LOC_275/Y 0.10fF
C25359 INVX1_LOC_93/Y INVX1_LOC_556/Y 0.01fF
C25360 INVX1_LOC_497/Y INVX1_LOC_259/Y 0.21fF
C25361 NAND2X1_LOC_307/A INVX1_LOC_9/Y 0.01fF
C25362 INVX1_LOC_53/A INVX1_LOC_6/Y 0.03fF
C25363 INVX1_LOC_282/A NAND2X1_LOC_850/a_36_24# 0.00fF
C25364 INVX1_LOC_40/Y NAND2X1_LOC_429/a_36_24# 0.00fF
C25365 INVX1_LOC_369/A NAND2X1_LOC_623/a_36_24# 0.00fF
C25366 INVX1_LOC_298/A INVX1_LOC_315/A 0.01fF
C25367 INVX1_LOC_63/Y INVX1_LOC_352/A 0.00fF
C25368 INVX1_LOC_99/Y INVX1_LOC_379/Y 0.11fF
C25369 INVX1_LOC_300/A NAND2X1_LOC_491/Y 0.02fF
C25370 INVX1_LOC_116/Y INVX1_LOC_58/Y 0.03fF
C25371 INVX1_LOC_53/Y INVX1_LOC_519/Y 0.00fF
C25372 INVX1_LOC_6/Y INVX1_LOC_50/Y 0.40fF
C25373 INVX1_LOC_551/A INVX1_LOC_35/Y -0.00fF
C25374 NAND2X1_LOC_599/a_36_24# INVX1_LOC_463/Y 0.00fF
C25375 INVX1_LOC_269/Y INVX1_LOC_270/Y 0.01fF
C25376 NAND2X1_LOC_184/Y NAND2X1_LOC_253/Y 0.08fF
C25377 NAND2X1_LOC_399/a_36_24# INVX1_LOC_328/Y 0.00fF
C25378 INVX1_LOC_117/Y INVX1_LOC_69/Y 0.26fF
C25379 INVX1_LOC_68/Y INVX1_LOC_91/Y 0.10fF
C25380 INVX1_LOC_31/Y NAND2X1_LOC_309/a_36_24# 0.01fF
C25381 INVX1_LOC_79/A INVX1_LOC_600/Y 0.00fF
C25382 NAND2X1_LOC_307/A INVX1_LOC_62/Y 0.12fF
C25383 INVX1_LOC_416/A INVX1_LOC_9/Y 0.03fF
C25384 INVX1_LOC_172/A INVX1_LOC_63/Y 0.56fF
C25385 INVX1_LOC_6/Y INVX1_LOC_431/Y 0.01fF
C25386 INVX1_LOC_318/A INVX1_LOC_199/Y 0.01fF
C25387 INVX1_LOC_361/A NAND2X1_LOC_267/A 0.15fF
C25388 INVX1_LOC_58/Y INPUT_4 0.03fF
C25389 INVX1_LOC_422/Y NAND2X1_LOC_294/Y 0.05fF
C25390 INVX1_LOC_81/Y INVX1_LOC_543/A 0.01fF
C25391 NAND2X1_LOC_545/A INVX1_LOC_98/Y 0.05fF
C25392 INVX1_LOC_431/A INVX1_LOC_90/Y 0.00fF
C25393 INVX1_LOC_11/Y INVX1_LOC_369/Y 0.07fF
C25394 INVX1_LOC_353/A NAND2X1_LOC_333/B 0.07fF
C25395 INVX1_LOC_89/Y INVX1_LOC_89/A 0.10fF
C25396 INVX1_LOC_671/A INVX1_LOC_663/A 0.02fF
C25397 INVX1_LOC_93/Y NAND2X1_LOC_420/Y 0.01fF
C25398 INVX1_LOC_255/A INVX1_LOC_58/Y 0.07fF
C25399 INVX1_LOC_360/Y INVX1_LOC_347/A 0.26fF
C25400 INVX1_LOC_6/A INVX1_LOC_25/A 0.21fF
C25401 INVX1_LOC_559/Y INVX1_LOC_242/Y 0.02fF
C25402 INVX1_LOC_419/Y INVX1_LOC_62/Y 0.10fF
C25403 INVX1_LOC_35/Y INVX1_LOC_75/Y 1.73fF
C25404 INVX1_LOC_304/A INVX1_LOC_75/Y 0.01fF
C25405 NAND2X1_LOC_7/Y INVX1_LOC_202/A 0.00fF
C25406 INVX1_LOC_204/Y INVX1_LOC_35/A 0.01fF
C25407 INVX1_LOC_31/Y NAND2X1_LOC_626/Y 0.03fF
C25408 NAND2X1_LOC_106/Y INVX1_LOC_100/Y 0.03fF
C25409 INVX1_LOC_245/A INVX1_LOC_296/A 0.00fF
C25410 INVX1_LOC_179/A INVX1_LOC_58/Y 0.01fF
C25411 INVX1_LOC_426/A INVX1_LOC_426/Y 0.02fF
C25412 INVX1_LOC_81/Y INVX1_LOC_86/A 0.01fF
C25413 INVX1_LOC_347/Y NAND2X1_LOC_299/a_36_24# 0.00fF
C25414 INVX1_LOC_479/A INVX1_LOC_686/Y 0.01fF
C25415 INVX1_LOC_379/A NAND2X1_LOC_271/A 0.01fF
C25416 VDD INVX1_LOC_152/Y 0.26fF
C25417 INVX1_LOC_204/Y INVX1_LOC_598/Y 0.00fF
C25418 INVX1_LOC_376/A INVX1_LOC_62/Y 0.07fF
C25419 INVX1_LOC_653/Y INVX1_LOC_338/Y 0.05fF
C25420 NAND2X1_LOC_121/Y INVX1_LOC_41/Y 0.09fF
C25421 NAND2X1_LOC_666/Y INVX1_LOC_74/Y 0.10fF
C25422 NAND2X1_LOC_660/a_36_24# INVX1_LOC_62/Y 0.00fF
C25423 NAND2X1_LOC_88/Y NAND2X1_LOC_100/a_36_24# 0.00fF
C25424 INVX1_LOC_206/Y INVX1_LOC_121/Y 0.03fF
C25425 NAND2X1_LOC_301/B INVX1_LOC_41/Y 0.69fF
C25426 INVX1_LOC_502/A INVX1_LOC_62/Y 0.07fF
C25427 INVX1_LOC_85/Y INVX1_LOC_180/Y 0.05fF
C25428 NAND2X1_LOC_249/Y INVX1_LOC_51/Y 3.28fF
C25429 NAND2X1_LOC_533/a_36_24# INVX1_LOC_510/Y 0.00fF
C25430 INVX1_LOC_203/Y INVX1_LOC_45/Y 0.03fF
C25431 NAND2X1_LOC_750/Y INVX1_LOC_85/Y 0.00fF
C25432 INVX1_LOC_459/A INVX1_LOC_134/Y 0.03fF
C25433 INVX1_LOC_301/A NAND2X1_LOC_129/a_36_24# 0.00fF
C25434 VDD INPUT_2 0.75fF
C25435 NAND2X1_LOC_475/A NAND2X1_LOC_493/B 0.01fF
C25436 INVX1_LOC_121/Y INVX1_LOC_242/A 0.03fF
C25437 INVX1_LOC_479/A INVX1_LOC_652/Y 0.02fF
C25438 NAND2X1_LOC_505/a_36_24# INVX1_LOC_397/A 0.00fF
C25439 NAND2X1_LOC_428/Y INVX1_LOC_74/Y 0.04fF
C25440 INVX1_LOC_266/A NAND2X1_LOC_373/a_36_24# 0.00fF
C25441 INVX1_LOC_137/A INVX1_LOC_185/Y 0.01fF
C25442 INVX1_LOC_594/Y INVX1_LOC_686/A 0.10fF
C25443 INVX1_LOC_438/A INVX1_LOC_486/Y 0.07fF
C25444 INVX1_LOC_100/Y INVX1_LOC_92/A 0.10fF
C25445 INVX1_LOC_271/A INVX1_LOC_76/Y 0.07fF
C25446 INVX1_LOC_266/A INVX1_LOC_560/A 0.10fF
C25447 INVX1_LOC_395/A INVX1_LOC_235/Y 0.03fF
C25448 INVX1_LOC_576/A INVX1_LOC_561/Y 0.06fF
C25449 INPUT_0 INVX1_LOC_90/A 0.01fF
C25450 INVX1_LOC_317/Y INVX1_LOC_270/A 0.25fF
C25451 VDD INVX1_LOC_252/Y 0.52fF
C25452 INVX1_LOC_74/Y INVX1_LOC_92/A 0.03fF
C25453 INVX1_LOC_446/Y INVX1_LOC_385/Y 0.70fF
C25454 NAND2X1_LOC_717/a_36_24# INVX1_LOC_230/A 0.01fF
C25455 NAND2X1_LOC_331/A INVX1_LOC_137/Y 0.03fF
C25456 INVX1_LOC_410/Y INVX1_LOC_510/A 0.00fF
C25457 INVX1_LOC_395/A INVX1_LOC_556/Y 0.12fF
C25458 INVX1_LOC_293/Y INVX1_LOC_655/Y 0.01fF
C25459 INVX1_LOC_603/Y NAND2X1_LOC_97/A 0.05fF
C25460 INVX1_LOC_447/A INVX1_LOC_32/Y 0.08fF
C25461 INVX1_LOC_390/Y INVX1_LOC_432/A 0.01fF
C25462 INVX1_LOC_435/Y INVX1_LOC_679/A 0.03fF
C25463 INVX1_LOC_557/A INVX1_LOC_251/A 0.15fF
C25464 INVX1_LOC_375/A INVX1_LOC_510/A 0.12fF
C25465 INVX1_LOC_118/Y INVX1_LOC_105/A 0.01fF
C25466 INVX1_LOC_395/A INVX1_LOC_81/Y 0.00fF
C25467 VDD NAND2X1_LOC_814/Y 0.05fF
C25468 INVX1_LOC_85/Y INVX1_LOC_44/A 0.38fF
C25469 NAND2X1_LOC_231/A INVX1_LOC_99/Y 0.00fF
C25470 INVX1_LOC_11/Y INVX1_LOC_428/A 0.03fF
C25471 NAND2X1_LOC_366/a_36_24# INVX1_LOC_321/A 0.00fF
C25472 INVX1_LOC_51/Y NAND2X1_LOC_275/Y 0.00fF
C25473 INVX1_LOC_384/A INVX1_LOC_385/Y 0.19fF
C25474 NAND2X1_LOC_61/A INVX1_LOC_44/Y 0.05fF
C25475 VDD NAND2X1_LOC_827/Y -0.00fF
C25476 NAND2X1_LOC_457/A INVX1_LOC_230/Y 0.00fF
C25477 INVX1_LOC_45/Y INVX1_LOC_194/Y 0.03fF
C25478 INVX1_LOC_670/Y INVX1_LOC_126/Y 0.02fF
C25479 INVX1_LOC_258/A INVX1_LOC_80/A 0.01fF
C25480 INVX1_LOC_686/A NAND2X1_LOC_603/Y 0.05fF
C25481 INVX1_LOC_576/A NAND2X1_LOC_733/a_36_24# 0.02fF
C25482 NAND2X1_LOC_331/A NAND2X1_LOC_829/B 0.04fF
C25483 NAND2X1_LOC_122/Y INVX1_LOC_259/Y 0.02fF
C25484 INVX1_LOC_575/A INVX1_LOC_569/A 0.05fF
C25485 NAND2X1_LOC_271/B INVX1_LOC_49/Y 0.03fF
C25486 NAND2X1_LOC_20/Y INVX1_LOC_7/Y 0.02fF
C25487 INVX1_LOC_117/Y INVX1_LOC_586/A 0.27fF
C25488 INVX1_LOC_578/A NAND2X1_LOC_443/a_36_24# 0.01fF
C25489 INVX1_LOC_206/Y NAND2X1_LOC_455/a_36_24# 0.00fF
C25490 INVX1_LOC_68/Y NAND2X1_LOC_333/B 0.16fF
C25491 INVX1_LOC_579/A NAND2X1_LOC_421/a_36_24# 0.00fF
C25492 NAND2X1_LOC_786/a_36_24# INVX1_LOC_198/A -0.02fF
C25493 INVX1_LOC_117/Y INVX1_LOC_516/Y 0.10fF
C25494 INVX1_LOC_115/A INVX1_LOC_633/Y 0.29fF
C25495 INVX1_LOC_366/A NAND2X1_LOC_235/a_36_24# 0.01fF
C25496 GATE_741 INVX1_LOC_93/Y 0.01fF
C25497 NAND2X1_LOC_460/A NAND2X1_LOC_379/a_36_24# 0.00fF
C25498 NAND2X1_LOC_360/a_36_24# INVX1_LOC_381/A 0.00fF
C25499 NAND2X1_LOC_733/a_36_24# INVX1_LOC_300/A 0.00fF
C25500 INVX1_LOC_381/A INPUT_1 0.11fF
C25501 INVX1_LOC_482/A INVX1_LOC_230/Y 0.02fF
C25502 INVX1_LOC_293/Y INVX1_LOC_277/A 0.01fF
C25503 NAND2X1_LOC_318/A INVX1_LOC_317/A 0.04fF
C25504 INVX1_LOC_20/Y INVX1_LOC_559/Y 0.04fF
C25505 INVX1_LOC_31/Y INVX1_LOC_235/Y 0.07fF
C25506 INVX1_LOC_395/A NAND2X1_LOC_420/Y -0.01fF
C25507 NAND2X1_LOC_358/a_36_24# INVX1_LOC_26/Y 0.00fF
C25508 INVX1_LOC_312/Y INVX1_LOC_117/Y 0.40fF
C25509 INVX1_LOC_45/Y INVX1_LOC_44/Y 0.03fF
C25510 INVX1_LOC_581/A INVX1_LOC_550/A 0.03fF
C25511 INVX1_LOC_379/A NAND2X1_LOC_462/a_36_24# 0.00fF
C25512 INVX1_LOC_400/Y NAND2X1_LOC_274/B 0.01fF
C25513 NAND2X1_LOC_130/Y INVX1_LOC_361/Y 0.05fF
C25514 INVX1_LOC_49/Y INVX1_LOC_169/A 0.01fF
C25515 INVX1_LOC_588/Y NAND2X1_LOC_755/B 0.00fF
C25516 INVX1_LOC_492/A INVX1_LOC_35/Y 0.03fF
C25517 INVX1_LOC_51/Y NAND2X1_LOC_605/B 0.01fF
C25518 INVX1_LOC_190/Y INVX1_LOC_190/A 0.09fF
C25519 INVX1_LOC_396/A INVX1_LOC_197/Y 0.12fF
C25520 INVX1_LOC_69/Y INVX1_LOC_658/A 0.01fF
C25521 NAND2X1_LOC_513/A INVX1_LOC_6/Y 1.44fF
C25522 INVX1_LOC_558/A NAND2X1_LOC_136/Y 0.04fF
C25523 INVX1_LOC_51/Y NAND2X1_LOC_626/Y 0.03fF
C25524 INVX1_LOC_40/Y INVX1_LOC_58/A 0.01fF
C25525 NAND2X1_LOC_542/a_36_24# NAND2X1_LOC_542/A 0.00fF
C25526 INVX1_LOC_49/Y INVX1_LOC_633/Y 0.03fF
C25527 INVX1_LOC_385/Y INVX1_LOC_433/A 0.03fF
C25528 NAND2X1_LOC_532/a_36_24# INVX1_LOC_62/Y 0.00fF
C25529 INVX1_LOC_537/A INVX1_LOC_463/Y 0.10fF
C25530 INVX1_LOC_285/A INVX1_LOC_63/Y 0.00fF
C25531 INVX1_LOC_670/Y INVX1_LOC_199/Y 0.02fF
C25532 INVX1_LOC_84/A INVX1_LOC_328/Y 0.07fF
C25533 INVX1_LOC_381/A INVX1_LOC_368/A 0.03fF
C25534 INVX1_LOC_160/A INVX1_LOC_89/Y 0.06fF
C25535 NAND2X1_LOC_149/a_36_24# INVX1_LOC_655/A 0.00fF
C25536 NAND2X1_LOC_467/A INVX1_LOC_500/A 0.01fF
C25537 INVX1_LOC_229/Y INVX1_LOC_223/Y 0.05fF
C25538 INVX1_LOC_160/A INVX1_LOC_154/A 0.33fF
C25539 INVX1_LOC_145/Y INVX1_LOC_493/Y 0.05fF
C25540 NAND2X1_LOC_317/a_36_24# INVX1_LOC_47/Y 0.01fF
C25541 INVX1_LOC_317/Y INVX1_LOC_75/A 0.27fF
C25542 NAND2X1_LOC_320/Y INVX1_LOC_63/Y 0.04fF
C25543 INVX1_LOC_326/Y INVX1_LOC_83/Y 0.02fF
C25544 INVX1_LOC_551/Y INVX1_LOC_41/Y 0.03fF
C25545 INVX1_LOC_300/Y INVX1_LOC_602/Y 0.02fF
C25546 INVX1_LOC_166/A INVX1_LOC_46/Y 0.03fF
C25547 NAND2X1_LOC_697/Y INVX1_LOC_168/Y 0.01fF
C25548 INVX1_LOC_268/A INVX1_LOC_245/A 0.03fF
C25549 INVX1_LOC_242/Y INVX1_LOC_155/Y 0.01fF
C25550 INVX1_LOC_463/Y INVX1_LOC_496/Y 0.03fF
C25551 INVX1_LOC_679/Y INVX1_LOC_100/Y 0.08fF
C25552 INVX1_LOC_17/Y INVX1_LOC_9/Y 0.22fF
C25553 INVX1_LOC_566/A INVX1_LOC_329/Y 0.03fF
C25554 NAND2X1_LOC_333/A NAND2X1_LOC_753/Y 0.17fF
C25555 NAND2X1_LOC_148/B INVX1_LOC_58/Y 0.01fF
C25556 INVX1_LOC_65/Y NAND2X1_LOC_60/Y 0.03fF
C25557 INVX1_LOC_380/A INVX1_LOC_297/Y 0.01fF
C25558 INVX1_LOC_197/A INVX1_LOC_479/A 0.07fF
C25559 INVX1_LOC_11/Y NAND2X1_LOC_106/a_36_24# 0.00fF
C25560 INVX1_LOC_468/Y INVX1_LOC_652/A 0.01fF
C25561 INVX1_LOC_53/Y INVX1_LOC_588/A 0.03fF
C25562 NAND2X1_LOC_192/A INVX1_LOC_50/Y 0.00fF
C25563 NAND2X1_LOC_317/a_36_24# INVX1_LOC_119/Y 0.00fF
C25564 INVX1_LOC_50/Y INVX1_LOC_206/A 0.01fF
C25565 INVX1_LOC_49/Y INVX1_LOC_490/A 0.45fF
C25566 INVX1_LOC_520/Y INVX1_LOC_66/A 0.00fF
C25567 INVX1_LOC_608/Y INVX1_LOC_62/Y 0.00fF
C25568 INVX1_LOC_12/Y INVX1_LOC_483/A 0.03fF
C25569 INVX1_LOC_602/Y INVX1_LOC_660/A 0.17fF
C25570 INVX1_LOC_156/Y INVX1_LOC_636/A 0.03fF
C25571 INVX1_LOC_124/Y INVX1_LOC_479/A 0.01fF
C25572 INVX1_LOC_69/Y INVX1_LOC_58/Y 1.08fF
C25573 INVX1_LOC_17/Y INVX1_LOC_62/Y 9.78fF
C25574 INVX1_LOC_80/A NAND2X1_LOC_832/A 0.08fF
C25575 INVX1_LOC_63/Y INVX1_LOC_199/Y 0.12fF
C25576 INVX1_LOC_44/Y NAND2X1_LOC_837/A 0.05fF
C25577 INVX1_LOC_675/A NAND2X1_LOC_586/Y 0.02fF
C25578 INVX1_LOC_100/Y INPUT_1 2.03fF
C25579 NAND2X1_LOC_307/B INVX1_LOC_9/Y 0.13fF
C25580 NAND2X1_LOC_542/A INVX1_LOC_376/Y 0.15fF
C25581 INVX1_LOC_662/Y NAND2X1_LOC_248/B 0.17fF
C25582 INVX1_LOC_493/A INVX1_LOC_41/Y 0.01fF
C25583 INVX1_LOC_479/A NAND2X1_LOC_106/B 0.02fF
C25584 INVX1_LOC_167/A INVX1_LOC_41/Y 0.01fF
C25585 INVX1_LOC_469/Y NAND2X1_LOC_123/B 0.03fF
C25586 INVX1_LOC_531/Y INVX1_LOC_46/Y 0.02fF
C25587 INPUT_1 INVX1_LOC_74/Y 0.15fF
C25588 GATE_662 INVX1_LOC_669/A 0.04fF
C25589 INVX1_LOC_11/Y NAND2X1_LOC_832/A 0.18fF
C25590 INVX1_LOC_63/Y INVX1_LOC_85/A 0.33fF
C25591 NAND2X1_LOC_502/a_36_24# INVX1_LOC_97/A 0.01fF
C25592 NAND2X1_LOC_827/Y INVX1_LOC_635/Y 0.01fF
C25593 INVX1_LOC_410/A INVX1_LOC_211/A 0.05fF
C25594 INVX1_LOC_50/Y INVX1_LOC_636/A 0.07fF
C25595 INVX1_LOC_380/A INVX1_LOC_76/Y 0.01fF
C25596 INVX1_LOC_620/A NAND2X1_LOC_98/B 0.10fF
C25597 NAND2X1_LOC_123/B INVX1_LOC_79/A 0.05fF
C25598 NAND2X1_LOC_249/Y INVX1_LOC_216/Y 0.19fF
C25599 NAND2X1_LOC_249/Y NAND2X1_LOC_108/Y 0.02fF
C25600 INVX1_LOC_601/A INVX1_LOC_366/A 0.35fF
C25601 NAND2X1_LOC_707/a_36_24# INVX1_LOC_373/A 0.00fF
C25602 VDD INVX1_LOC_85/Y 0.27fF
C25603 INVX1_LOC_150/A INVX1_LOC_542/A 0.02fF
C25604 NAND2X1_LOC_433/Y NAND2X1_LOC_832/A 0.03fF
C25605 INVX1_LOC_435/Y INVX1_LOC_490/Y 0.91fF
C25606 INVX1_LOC_118/Y INVX1_LOC_45/Y 0.04fF
C25607 INVX1_LOC_601/A NAND2X1_LOC_240/a_36_24# 0.00fF
C25608 INVX1_LOC_410/Y INVX1_LOC_321/A 0.06fF
C25609 NAND2X1_LOC_271/B INVX1_LOC_76/Y 0.00fF
C25610 INVX1_LOC_40/Y INVX1_LOC_41/A 0.03fF
C25611 INVX1_LOC_3/Y INVX1_LOC_595/A 0.01fF
C25612 INVX1_LOC_96/Y NAND2X1_LOC_506/B 0.11fF
C25613 INVX1_LOC_75/Y INVX1_LOC_364/A 0.03fF
C25614 INVX1_LOC_96/Y INVX1_LOC_45/Y 0.01fF
C25615 NAND2X1_LOC_13/Y INVX1_LOC_560/A 0.06fF
C25616 INVX1_LOC_79/A INVX1_LOC_92/A 0.06fF
C25617 INVX1_LOC_617/Y INVX1_LOC_410/Y 0.08fF
C25618 VDD INVX1_LOC_599/Y 0.04fF
C25619 INVX1_LOC_617/Y INVX1_LOC_375/A 0.01fF
C25620 INVX1_LOC_617/Y INVX1_LOC_546/A 0.03fF
C25621 NAND2X1_LOC_531/a_36_24# INVX1_LOC_7/Y 0.00fF
C25622 INVX1_LOC_317/Y NAND2X1_LOC_318/A 0.28fF
C25623 NAND2X1_LOC_685/B NAND2X1_LOC_651/a_36_24# 0.00fF
C25624 INVX1_LOC_51/A INVX1_LOC_80/A 0.10fF
C25625 INVX1_LOC_386/Y INVX1_LOC_453/A 0.06fF
C25626 NAND2X1_LOC_241/B INVX1_LOC_80/A 0.05fF
C25627 NAND2X1_LOC_475/A INVX1_LOC_321/Y 0.01fF
C25628 INVX1_LOC_51/Y INVX1_LOC_235/Y 0.07fF
C25629 INVX1_LOC_224/Y INVX1_LOC_379/A 0.14fF
C25630 INVX1_LOC_567/A INVX1_LOC_117/Y 0.01fF
C25631 INVX1_LOC_355/Y INVX1_LOC_638/A 0.00fF
C25632 NAND2X1_LOC_498/B INVX1_LOC_633/Y 0.03fF
C25633 INVX1_LOC_224/Y INVX1_LOC_35/Y 0.17fF
C25634 INVX1_LOC_20/Y NAND2X1_LOC_710/A 0.00fF
C25635 INVX1_LOC_218/Y INVX1_LOC_438/Y 0.01fF
C25636 INVX1_LOC_607/Y INVX1_LOC_605/A 0.06fF
C25637 INVX1_LOC_601/A INVX1_LOC_6/Y 0.01fF
C25638 INVX1_LOC_76/Y INVX1_LOC_633/Y 0.28fF
C25639 INPUT_0 NAND2X1_LOC_187/Y 0.01fF
C25640 NAND2X1_LOC_320/Y INVX1_LOC_374/A 0.02fF
C25641 NAND2X1_LOC_399/B INVX1_LOC_322/Y 0.72fF
C25642 NAND2X1_LOC_789/a_36_24# INVX1_LOC_366/A 0.01fF
C25643 INVX1_LOC_578/A INVX1_LOC_35/Y 0.14fF
C25644 INVX1_LOC_428/A INVX1_LOC_367/Y 0.01fF
C25645 INVX1_LOC_578/A INVX1_LOC_304/A 0.06fF
C25646 NAND2X1_LOC_704/B INVX1_LOC_558/Y 0.14fF
C25647 INVX1_LOC_602/A INVX1_LOC_272/Y 0.04fF
C25648 INPUT_0 INVX1_LOC_54/Y 0.35fF
C25649 INVX1_LOC_602/A NAND2X1_LOC_791/B 0.40fF
C25650 INVX1_LOC_214/Y INVX1_LOC_607/A 0.56fF
C25651 NAND2X1_LOC_516/Y NAND2X1_LOC_602/A 0.01fF
C25652 INVX1_LOC_400/Y INVX1_LOC_159/Y 0.07fF
C25653 INVX1_LOC_233/Y INVX1_LOC_442/Y 0.05fF
C25654 VDD INVX1_LOC_419/A 0.00fF
C25655 INVX1_LOC_97/A NAND2X1_LOC_503/Y 0.00fF
C25656 GATE_579 NAND2X1_LOC_569/a_36_24# 0.00fF
C25657 VDD INVX1_LOC_234/Y 0.21fF
C25658 INVX1_LOC_586/A INVX1_LOC_178/A 0.07fF
C25659 VDD INVX1_LOC_573/Y 0.30fF
C25660 INVX1_LOC_117/Y INVX1_LOC_140/Y 0.03fF
C25661 INVX1_LOC_20/Y INVX1_LOC_155/Y 0.06fF
C25662 INPUT_3 INVX1_LOC_27/Y 0.18fF
C25663 INVX1_LOC_17/Y INVX1_LOC_547/A 0.02fF
C25664 INVX1_LOC_144/Y INVX1_LOC_137/Y 0.01fF
C25665 INVX1_LOC_271/A INVX1_LOC_32/Y 0.01fF
C25666 INVX1_LOC_53/Y INVX1_LOC_670/Y 0.01fF
C25667 INVX1_LOC_438/Y NAND2X1_LOC_256/a_36_24# 0.01fF
C25668 INVX1_LOC_255/Y INVX1_LOC_359/A 0.01fF
C25669 NAND2X1_LOC_325/B INVX1_LOC_134/Y 0.01fF
C25670 INVX1_LOC_288/A INVX1_LOC_354/Y 0.01fF
C25671 NAND2X1_LOC_210/A INVX1_LOC_522/Y 0.04fF
C25672 INVX1_LOC_85/Y NAND2X1_LOC_243/A 0.16fF
C25673 INVX1_LOC_173/A INVX1_LOC_32/Y 0.01fF
C25674 NAND2X1_LOC_723/a_36_24# INVX1_LOC_353/A 0.01fF
C25675 INVX1_LOC_322/Y INVX1_LOC_32/Y 0.04fF
C25676 INVX1_LOC_117/Y INVX1_LOC_366/A 0.01fF
C25677 INVX1_LOC_552/Y INVX1_LOC_199/Y 0.03fF
C25678 INVX1_LOC_318/Y INVX1_LOC_230/A 0.04fF
C25679 INVX1_LOC_588/Y INVX1_LOC_268/Y 0.18fF
C25680 INVX1_LOC_560/A INVX1_LOC_361/A 0.02fF
C25681 INVX1_LOC_612/Y INVX1_LOC_610/Y 0.01fF
C25682 INVX1_LOC_54/Y INVX1_LOC_586/Y 0.01fF
C25683 INVX1_LOC_381/A INVX1_LOC_50/Y 0.31fF
C25684 INVX1_LOC_76/Y INVX1_LOC_490/A 0.03fF
C25685 INVX1_LOC_569/A INVX1_LOC_575/Y 0.25fF
C25686 NAND2X1_LOC_45/Y NAND2X1_LOC_274/B 0.40fF
C25687 INVX1_LOC_84/A INVX1_LOC_172/A 0.02fF
C25688 INVX1_LOC_53/A INVX1_LOC_29/Y 0.01fF
C25689 INVX1_LOC_17/Y INVX1_LOC_344/A 0.01fF
C25690 NAND2X1_LOC_397/Y INVX1_LOC_7/Y 0.02fF
C25691 NAND2X1_LOC_231/A INVX1_LOC_96/A 0.03fF
C25692 INVX1_LOC_76/Y INVX1_LOC_317/A 0.00fF
C25693 NAND2X1_LOC_791/B INVX1_LOC_117/Y 0.07fF
C25694 INVX1_LOC_7/Y NAND2X1_LOC_415/B 0.06fF
C25695 INVX1_LOC_300/A INVX1_LOC_155/Y 0.03fF
C25696 INVX1_LOC_579/A INVX1_LOC_259/Y 0.01fF
C25697 INVX1_LOC_272/Y INVX1_LOC_117/Y 3.79fF
C25698 INVX1_LOC_228/A NAND2X1_LOC_266/a_36_24# 0.00fF
C25699 INVX1_LOC_117/Y INVX1_LOC_486/Y 2.82fF
C25700 INVX1_LOC_186/A INVX1_LOC_145/Y 0.00fF
C25701 INVX1_LOC_376/Y INVX1_LOC_253/A 0.03fF
C25702 NAND2X1_LOC_376/Y INVX1_LOC_365/A 0.09fF
C25703 INVX1_LOC_586/A INVX1_LOC_58/Y 2.30fF
C25704 INVX1_LOC_404/Y INVX1_LOC_502/A 0.01fF
C25705 INVX1_LOC_568/Y INVX1_LOC_35/Y 0.01fF
C25706 NAND2X1_LOC_304/a_36_24# NAND2X1_LOC_267/A -0.01fF
C25707 INVX1_LOC_516/Y INVX1_LOC_58/Y 0.01fF
C25708 INVX1_LOC_384/A INVX1_LOC_420/A 0.09fF
C25709 VDD INVX1_LOC_505/Y 0.55fF
C25710 INVX1_LOC_542/A NAND2X1_LOC_639/a_36_24# 0.00fF
C25711 NAND2X1_LOC_259/A NAND2X1_LOC_257/a_36_24# 0.02fF
C25712 INVX1_LOC_602/A INVX1_LOC_6/Y 0.07fF
C25713 NAND2X1_LOC_697/Y INVX1_LOC_137/Y 0.02fF
C25714 NAND2X1_LOC_498/Y NAND2X1_LOC_274/B 0.06fF
C25715 NAND2X1_LOC_383/Y INVX1_LOC_314/Y 0.17fF
C25716 INVX1_LOC_243/A INPUT_1 0.01fF
C25717 INVX1_LOC_570/A NAND2X1_LOC_274/B 0.04fF
C25718 NAND2X1_LOC_190/A INVX1_LOC_17/Y 0.01fF
C25719 INVX1_LOC_597/A INVX1_LOC_117/Y 0.01fF
C25720 INVX1_LOC_255/Y NAND2X1_LOC_301/B 0.03fF
C25721 INVX1_LOC_402/A INVX1_LOC_520/A 0.10fF
C25722 INVX1_LOC_173/Y INVX1_LOC_12/Y 0.06fF
C25723 INVX1_LOC_607/Y INVX1_LOC_54/Y 0.45fF
C25724 INVX1_LOC_676/Y INVX1_LOC_463/Y 0.05fF
C25725 INVX1_LOC_53/Y INVX1_LOC_253/Y 0.44fF
C25726 VDD NAND2X1_LOC_231/B 0.01fF
C25727 INVX1_LOC_300/A NAND2X1_LOC_853/a_36_24# 0.00fF
C25728 INVX1_LOC_11/Y INVX1_LOC_371/A 0.00fF
C25729 NAND2X1_LOC_596/Y INVX1_LOC_505/Y 0.02fF
C25730 INVX1_LOC_85/Y NAND2X1_LOC_786/B 0.02fF
C25731 NAND2X1_LOC_756/Y INVX1_LOC_44/Y 0.09fF
C25732 INPUT_0 INVX1_LOC_388/A 0.00fF
C25733 INVX1_LOC_312/Y INVX1_LOC_58/Y 0.00fF
C25734 NAND2X1_LOC_696/a_36_24# INVX1_LOC_48/Y 0.00fF
C25735 INVX1_LOC_418/A INVX1_LOC_41/Y 0.01fF
C25736 INVX1_LOC_53/Y INVX1_LOC_63/Y 0.22fF
C25737 NAND2X1_LOC_333/a_36_24# NAND2X1_LOC_755/B 0.00fF
C25738 NAND2X1_LOC_720/A INVX1_LOC_50/Y 0.28fF
C25739 INVX1_LOC_439/Y INVX1_LOC_385/A 0.09fF
C25740 NAND2X1_LOC_775/B INVX1_LOC_32/Y 0.07fF
C25741 NAND2X1_LOC_160/a_36_24# INVX1_LOC_496/A 0.01fF
C25742 INVX1_LOC_206/Y INVX1_LOC_462/Y 0.36fF
C25743 INVX1_LOC_377/Y NAND2X1_LOC_274/B 0.01fF
C25744 INVX1_LOC_43/A INVX1_LOC_86/Y 0.01fF
C25745 NAND2X1_LOC_79/B INVX1_LOC_207/Y 0.29fF
C25746 NAND2X1_LOC_318/A INVX1_LOC_531/Y 0.03fF
C25747 INVX1_LOC_410/A INVX1_LOC_145/Y 0.02fF
C25748 INVX1_LOC_508/Y INVX1_LOC_655/A -0.00fF
C25749 INVX1_LOC_482/Y INVX1_LOC_600/A 0.02fF
C25750 INVX1_LOC_145/Y INVX1_LOC_420/A 0.03fF
C25751 INVX1_LOC_17/Y INVX1_LOC_624/Y 0.02fF
C25752 INVX1_LOC_93/Y NAND2X1_LOC_444/A 0.04fF
C25753 INVX1_LOC_270/A INVX1_LOC_41/Y 0.06fF
C25754 INVX1_LOC_120/Y INVX1_LOC_304/A 0.02fF
C25755 INVX1_LOC_117/Y INVX1_LOC_6/Y 0.70fF
C25756 NAND2X1_LOC_576/a_36_24# INVX1_LOC_443/A 0.06fF
C25757 INVX1_LOC_166/A INVX1_LOC_387/Y 0.01fF
C25758 NAND2X1_LOC_818/a_36_24# INVX1_LOC_669/A 0.01fF
C25759 INVX1_LOC_588/Y INVX1_LOC_49/Y 0.03fF
C25760 INVX1_LOC_103/Y INVX1_LOC_234/Y 0.09fF
C25761 NAND2X1_LOC_274/B INVX1_LOC_99/Y 0.03fF
C25762 INVX1_LOC_166/A INVX1_LOC_49/Y 0.07fF
C25763 INVX1_LOC_157/A INVX1_LOC_157/Y 0.00fF
C25764 INVX1_LOC_202/Y INVX1_LOC_153/Y 0.48fF
C25765 INVX1_LOC_46/Y INVX1_LOC_411/Y 0.02fF
C25766 NAND2X1_LOC_755/B INVX1_LOC_41/Y 0.03fF
C25767 INVX1_LOC_672/A INVX1_LOC_655/A 0.03fF
C25768 INVX1_LOC_291/A NAND2X1_LOC_98/B 0.16fF
C25769 INVX1_LOC_367/A INVX1_LOC_109/A 0.03fF
C25770 INVX1_LOC_449/A NAND2X1_LOC_497/a_36_24# 0.00fF
C25771 INVX1_LOC_681/Y INVX1_LOC_79/A 0.03fF
C25772 INVX1_LOC_63/Y NAND2X1_LOC_346/B 0.06fF
C25773 INVX1_LOC_439/Y INVX1_LOC_244/Y 0.03fF
C25774 INVX1_LOC_686/A INVX1_LOC_462/Y 0.02fF
C25775 INVX1_LOC_100/Y INVX1_LOC_50/Y 2.16fF
C25776 INVX1_LOC_79/A INPUT_1 9.59fF
C25777 INVX1_LOC_359/A INVX1_LOC_26/Y 0.01fF
C25778 NAND2X1_LOC_123/B INVX1_LOC_48/Y 0.03fF
C25779 INVX1_LOC_660/Y INVX1_LOC_673/Y 0.00fF
C25780 INVX1_LOC_73/Y NAND2X1_LOC_69/B 0.17fF
C25781 INVX1_LOC_21/Y INVX1_LOC_634/Y 0.07fF
C25782 NAND2X1_LOC_389/a_36_24# INVX1_LOC_100/Y 0.00fF
C25783 INVX1_LOC_281/A INVX1_LOC_369/Y 0.05fF
C25784 INVX1_LOC_69/Y INVX1_LOC_245/A 0.06fF
C25785 INVX1_LOC_47/Y NAND2X1_LOC_274/B 0.07fF
C25786 INVX1_LOC_79/A INVX1_LOC_292/Y 0.04fF
C25787 INVX1_LOC_74/Y INVX1_LOC_50/Y 0.03fF
C25788 INVX1_LOC_41/Y INVX1_LOC_46/Y 0.12fF
C25789 INVX1_LOC_62/Y INVX1_LOC_230/Y 0.29fF
C25790 INVX1_LOC_54/Y INVX1_LOC_211/A 0.07fF
C25791 INVX1_LOC_50/Y INVX1_LOC_483/Y 0.01fF
C25792 INVX1_LOC_417/Y INVX1_LOC_92/A 0.52fF
C25793 INVX1_LOC_145/Y INVX1_LOC_611/A 0.01fF
C25794 INVX1_LOC_79/A INVX1_LOC_284/Y 0.01fF
C25795 NAND2X1_LOC_614/a_36_24# INVX1_LOC_211/A 0.00fF
C25796 INVX1_LOC_199/Y INVX1_LOC_669/A 0.01fF
C25797 NAND2X1_LOC_128/A INVX1_LOC_479/A 0.02fF
C25798 INVX1_LOC_652/Y INVX1_LOC_66/A 0.02fF
C25799 INVX1_LOC_49/Y INVX1_LOC_531/Y 0.02fF
C25800 INVX1_LOC_270/Y INVX1_LOC_48/Y 0.03fF
C25801 INVX1_LOC_93/Y INVX1_LOC_109/A 0.00fF
C25802 INVX1_LOC_507/A INVX1_LOC_62/Y 0.01fF
C25803 INVX1_LOC_81/A INVX1_LOC_85/A 0.06fF
C25804 NAND2X1_LOC_274/B INVX1_LOC_119/Y 0.06fF
C25805 INVX1_LOC_531/Y INVX1_LOC_642/Y 0.01fF
C25806 INVX1_LOC_550/A INVX1_LOC_613/A 0.02fF
C25807 INVX1_LOC_487/Y INVX1_LOC_79/A 0.07fF
C25808 INVX1_LOC_48/Y INVX1_LOC_92/A 2.13fF
C25809 INVX1_LOC_84/A INVX1_LOC_109/Y 0.01fF
C25810 INVX1_LOC_47/Y NAND2X1_LOC_449/a_36_24# 0.00fF
C25811 INVX1_LOC_278/A INVX1_LOC_445/A 0.68fF
C25812 INVX1_LOC_68/Y NAND2X1_LOC_723/a_36_24# 0.00fF
C25813 INVX1_LOC_438/Y INVX1_LOC_429/Y 0.03fF
C25814 INVX1_LOC_63/Y NAND2X1_LOC_60/Y 0.07fF
C25815 NAND2X1_LOC_636/A NAND2X1_LOC_192/a_36_24# 0.01fF
C25816 INVX1_LOC_414/A INVX1_LOC_427/A 0.31fF
C25817 INVX1_LOC_446/A INVX1_LOC_53/Y 0.16fF
C25818 INVX1_LOC_375/A INVX1_LOC_546/A 0.02fF
C25819 INVX1_LOC_41/Y INVX1_LOC_75/A 0.01fF
C25820 NAND2X1_LOC_432/a_36_24# NAND2X1_LOC_832/A 0.00fF
C25821 INVX1_LOC_483/A NAND2X1_LOC_621/B 0.22fF
C25822 INVX1_LOC_459/Y INVX1_LOC_374/A 0.14fF
C25823 VDD INVX1_LOC_80/A 1.47fF
C25824 VDD NAND2X1_LOC_768/A 0.18fF
C25825 VDD INVX1_LOC_579/Y 0.33fF
C25826 NAND2X1_LOC_142/a_36_24# INVX1_LOC_651/A 0.00fF
C25827 INVX1_LOC_200/Y INVX1_LOC_367/A 0.03fF
C25828 INVX1_LOC_317/Y INVX1_LOC_76/Y 0.03fF
C25829 NAND2X1_LOC_457/A INVX1_LOC_519/A 0.03fF
C25830 INVX1_LOC_401/A NAND2X1_LOC_513/Y 0.02fF
C25831 INVX1_LOC_160/Y INVX1_LOC_287/Y 0.01fF
C25832 INVX1_LOC_453/A INVX1_LOC_7/Y 0.10fF
C25833 NAND2X1_LOC_756/Y INVX1_LOC_96/Y 0.05fF
C25834 INVX1_LOC_307/Y INVX1_LOC_7/Y 0.01fF
C25835 NAND2X1_LOC_13/Y NAND2X1_LOC_491/a_36_24# 0.00fF
C25836 VDD INVX1_LOC_11/Y 1.71fF
C25837 INVX1_LOC_206/Y INVX1_LOC_379/A 0.14fF
C25838 INVX1_LOC_156/Y INVX1_LOC_566/A 0.03fF
C25839 INVX1_LOC_206/Y INVX1_LOC_35/Y 0.46fF
C25840 INVX1_LOC_206/Y INVX1_LOC_304/A 0.08fF
C25841 INVX1_LOC_510/Y INVX1_LOC_80/A 0.07fF
C25842 INVX1_LOC_453/Y INVX1_LOC_445/A 0.03fF
C25843 INVX1_LOC_185/A INVX1_LOC_6/Y 0.01fF
C25844 NAND2X1_LOC_302/a_36_24# NAND2X1_LOC_122/Y 0.00fF
C25845 INVX1_LOC_85/Y INVX1_LOC_619/A 0.05fF
C25846 INPUT_3 INPUT_2 0.55fF
C25847 INVX1_LOC_582/Y INVX1_LOC_583/A 0.15fF
C25848 INVX1_LOC_648/Y INVX1_LOC_35/Y 0.01fF
C25849 INVX1_LOC_257/Y INVX1_LOC_54/Y 0.28fF
C25850 INPUT_0 INVX1_LOC_585/Y 0.01fF
C25851 INVX1_LOC_395/A INVX1_LOC_304/Y 0.02fF
C25852 INVX1_LOC_407/Y NAND2X1_LOC_532/a_36_24# 0.00fF
C25853 INVX1_LOC_315/Y NAND2X1_LOC_755/B 0.03fF
C25854 INVX1_LOC_53/Y INVX1_LOC_20/A 0.02fF
C25855 INPUT_3 INVX1_LOC_297/A 0.54fF
C25856 INVX1_LOC_239/Y NAND2X1_LOC_286/A 0.02fF
C25857 INVX1_LOC_567/A INVX1_LOC_58/Y 0.00fF
C25858 NAND2X1_LOC_636/A INVX1_LOC_338/Y 0.02fF
C25859 INVX1_LOC_413/Y INVX1_LOC_392/A 0.00fF
C25860 INVX1_LOC_628/Y NAND2X1_LOC_173/Y 0.05fF
C25861 INVX1_LOC_20/Y NAND2X1_LOC_197/a_36_24# 0.00fF
C25862 NAND2X1_LOC_704/B NAND2X1_LOC_413/Y 0.23fF
C25863 INVX1_LOC_578/A INVX1_LOC_360/A 0.10fF
C25864 INVX1_LOC_447/Y INVX1_LOC_384/A 0.02fF
C25865 INPUT_0 INVX1_LOC_395/Y 0.01fF
C25866 INVX1_LOC_206/Y INVX1_LOC_620/A 0.07fF
C25867 NAND2X1_LOC_21/a_36_24# INPUT_4 0.00fF
C25868 INPUT_0 INVX1_LOC_199/A 0.02fF
C25869 NAND2X1_LOC_538/B INVX1_LOC_99/Y 0.02fF
C25870 INVX1_LOC_11/Y INVX1_LOC_510/Y 0.16fF
C25871 INVX1_LOC_396/Y INVX1_LOC_35/Y 0.28fF
C25872 INPUT_0 INVX1_LOC_89/Y 0.25fF
C25873 INVX1_LOC_35/Y INVX1_LOC_242/A 0.03fF
C25874 INVX1_LOC_375/Y INVX1_LOC_383/Y 0.01fF
C25875 INVX1_LOC_318/Y NAND2X1_LOC_72/Y 0.00fF
C25876 NAND2X1_LOC_475/A NAND2X1_LOC_212/a_36_24# 0.00fF
C25877 INVX1_LOC_294/Y INVX1_LOC_281/Y 0.05fF
C25878 NAND2X1_LOC_637/A INVX1_LOC_245/A 0.07fF
C25879 INVX1_LOC_166/A NAND2X1_LOC_498/B 0.01fF
C25880 VDD INVX1_LOC_50/A -0.00fF
C25881 INVX1_LOC_150/Y INVX1_LOC_498/A 0.09fF
C25882 INVX1_LOC_537/Y INVX1_LOC_676/Y 0.25fF
C25883 INVX1_LOC_288/A NAND2X1_LOC_173/a_36_24# 0.01fF
C25884 INVX1_LOC_54/Y INVX1_LOC_384/A 0.10fF
C25885 INVX1_LOC_549/A INVX1_LOC_338/Y 0.10fF
C25886 INVX1_LOC_558/A NAND2X1_LOC_137/A 0.07fF
C25887 VDD NAND2X1_LOC_433/Y 0.34fF
C25888 INVX1_LOC_302/A INVX1_LOC_387/Y 0.03fF
C25889 INVX1_LOC_686/A INVX1_LOC_35/Y 0.02fF
C25890 INVX1_LOC_686/A INVX1_LOC_304/A 0.04fF
C25891 INPUT_0 INVX1_LOC_501/A 0.16fF
C25892 INVX1_LOC_522/Y NAND2X1_LOC_594/Y 0.04fF
C25893 INVX1_LOC_402/Y NAND2X1_LOC_411/Y 0.01fF
C25894 NAND2X1_LOC_324/B NAND2X1_LOC_324/a_36_24# 0.00fF
C25895 INVX1_LOC_256/A INVX1_LOC_633/Y 0.28fF
C25896 INVX1_LOC_335/Y NAND2X1_LOC_755/B 3.76fF
C25897 INVX1_LOC_166/A INVX1_LOC_76/Y 0.03fF
C25898 INVX1_LOC_287/Y NAND2X1_LOC_267/A 0.03fF
C25899 INVX1_LOC_80/A INVX1_LOC_509/A 0.01fF
C25900 NAND2X1_LOC_140/B NAND2X1_LOC_131/a_36_24# 0.03fF
C25901 INVX1_LOC_32/Y INVX1_LOC_169/A 0.01fF
C25902 INVX1_LOC_270/A NAND2X1_LOC_267/A 0.20fF
C25903 VDD INVX1_LOC_102/Y 0.26fF
C25904 INVX1_LOC_137/Y INVX1_LOC_134/Y 0.13fF
C25905 NAND2X1_LOC_139/a_36_24# INPUT_1 0.01fF
C25906 NAND2X1_LOC_596/a_36_24# INVX1_LOC_513/A 0.00fF
C25907 INVX1_LOC_570/A INVX1_LOC_569/Y 0.14fF
C25908 INVX1_LOC_206/Y INVX1_LOC_518/Y 0.04fF
C25909 NAND2X1_LOC_22/a_36_24# INVX1_LOC_6/Y 0.01fF
C25910 INVX1_LOC_395/A INVX1_LOC_389/Y 0.01fF
C25911 NAND2X1_LOC_370/A INVX1_LOC_9/Y -0.07fF
C25912 NAND2X1_LOC_7/a_36_24# INVX1_LOC_6/Y 0.00fF
C25913 INVX1_LOC_587/A INVX1_LOC_58/Y 0.01fF
C25914 INVX1_LOC_251/Y INVX1_LOC_252/A 0.03fF
C25915 INVX1_LOC_103/Y INVX1_LOC_80/A 0.58fF
C25916 INVX1_LOC_230/A INVX1_LOC_98/Y 0.40fF
C25917 INVX1_LOC_613/Y INVX1_LOC_54/Y 0.01fF
C25918 INVX1_LOC_55/A INVX1_LOC_57/Y 0.00fF
C25919 NAND2X1_LOC_588/a_36_24# INVX1_LOC_315/A 0.00fF
C25920 INVX1_LOC_417/Y INPUT_1 0.00fF
C25921 INVX1_LOC_267/Y NAND2X1_LOC_333/A 0.01fF
C25922 INVX1_LOC_99/Y INVX1_LOC_159/Y 0.03fF
C25923 INVX1_LOC_447/A INVX1_LOC_75/Y 0.02fF
C25924 INVX1_LOC_54/Y NAND2X1_LOC_612/A 0.02fF
C25925 INVX1_LOC_161/A INVX1_LOC_117/Y 0.01fF
C25926 INVX1_LOC_84/A INVX1_LOC_199/Y 0.10fF
C25927 INVX1_LOC_17/Y INVX1_LOC_480/Y 0.02fF
C25928 INVX1_LOC_586/A INVX1_LOC_245/A 0.16fF
C25929 INVX1_LOC_654/A INVX1_LOC_654/Y 0.06fF
C25930 INPUT_5 INVX1_LOC_5/Y 0.04fF
C25931 INVX1_LOC_11/Y INVX1_LOC_509/A 0.11fF
C25932 INVX1_LOC_54/Y INVX1_LOC_145/Y 1.65fF
C25933 NAND2X1_LOC_57/Y INVX1_LOC_50/Y 0.02fF
C25934 NAND2X1_LOC_332/B INVX1_LOC_124/A 0.35fF
C25935 NAND2X1_LOC_45/Y NAND2X1_LOC_617/a_36_24# 0.00fF
C25936 INVX1_LOC_21/Y INVX1_LOC_46/Y 0.05fF
C25937 INVX1_LOC_65/Y NAND2X1_LOC_545/A 0.01fF
C25938 INVX1_LOC_58/Y NAND2X1_LOC_820/A 0.01fF
C25939 INVX1_LOC_502/Y NAND2X1_LOC_274/B 0.00fF
C25940 INVX1_LOC_89/Y NAND2X1_LOC_123/A 0.03fF
C25941 INVX1_LOC_166/A NAND2X1_LOC_446/a_36_24# 0.00fF
C25942 NAND2X1_LOC_498/Y INVX1_LOC_468/A 0.06fF
C25943 INVX1_LOC_17/Y INVX1_LOC_169/Y 0.48fF
C25944 INVX1_LOC_666/A INVX1_LOC_90/Y 0.01fF
C25945 INVX1_LOC_381/A NAND2X1_LOC_293/a_36_24# 0.00fF
C25946 NAND2X1_LOC_677/Y INVX1_LOC_476/Y 0.03fF
C25947 INVX1_LOC_76/Y INVX1_LOC_153/Y 0.01fF
C25948 VDD INVX1_LOC_231/Y 0.21fF
C25949 INVX1_LOC_681/Y INVX1_LOC_48/Y 0.09fF
C25950 INVX1_LOC_98/A INVX1_LOC_531/Y 0.04fF
C25951 INVX1_LOC_11/Y INVX1_LOC_103/Y 0.08fF
C25952 INVX1_LOC_578/A INVX1_LOC_364/A 0.05fF
C25953 INVX1_LOC_544/Y INVX1_LOC_670/Y 0.04fF
C25954 INPUT_1 INVX1_LOC_48/Y 0.04fF
C25955 INVX1_LOC_51/A INVX1_LOC_625/Y 0.24fF
C25956 NAND2X1_LOC_636/B NAND2X1_LOC_192/A 0.19fF
C25957 INVX1_LOC_6/Y INVX1_LOC_178/A 0.31fF
C25958 NAND2X1_LOC_122/Y INVX1_LOC_62/Y 0.11fF
C25959 INVX1_LOC_84/A INVX1_LOC_85/A 0.03fF
C25960 NAND2X1_LOC_318/A INVX1_LOC_41/Y 0.04fF
C25961 INVX1_LOC_89/Y INVX1_LOC_527/Y 0.01fF
C25962 INVX1_LOC_288/Y INVX1_LOC_675/A 0.02fF
C25963 INVX1_LOC_47/Y INVX1_LOC_159/Y 0.03fF
C25964 INVX1_LOC_581/A INVX1_LOC_612/A 0.19fF
C25965 INVX1_LOC_255/Y INVX1_LOC_634/Y 0.01fF
C25966 INVX1_LOC_292/Y INVX1_LOC_48/Y 0.16fF
C25967 INVX1_LOC_12/Y INVX1_LOC_485/Y 0.01fF
C25968 INVX1_LOC_316/Y INPUT_5 0.01fF
C25969 INVX1_LOC_35/Y NAND2X1_LOC_334/A 0.04fF
C25970 NAND2X1_LOC_181/A INVX1_LOC_50/Y 0.01fF
C25971 INVX1_LOC_32/Y INVX1_LOC_317/A 0.01fF
C25972 INVX1_LOC_342/Y INVX1_LOC_674/Y 0.06fF
C25973 INVX1_LOC_608/A INVX1_LOC_6/Y 2.23fF
C25974 INVX1_LOC_301/Y INVX1_LOC_363/Y 0.07fF
C25975 INVX1_LOC_555/A INVX1_LOC_46/Y 0.01fF
C25976 INVX1_LOC_213/Y INVX1_LOC_63/Y 0.04fF
C25977 INVX1_LOC_617/Y INVX1_LOC_479/A 0.07fF
C25978 INVX1_LOC_53/Y INVX1_LOC_669/A 0.03fF
C25979 INVX1_LOC_492/A INVX1_LOC_507/Y 0.18fF
C25980 INVX1_LOC_54/Y NAND2X1_LOC_490/a_36_24# 0.00fF
C25981 NAND2X1_LOC_72/Y INVX1_LOC_90/Y 0.03fF
C25982 NAND2X1_LOC_513/Y INVX1_LOC_92/A 0.09fF
C25983 INVX1_LOC_17/Y NAND2X1_LOC_833/B 0.03fF
C25984 INVX1_LOC_627/Y INVX1_LOC_633/A 0.15fF
C25985 NAND2X1_LOC_192/A INVX1_LOC_117/Y 0.03fF
C25986 INVX1_LOC_115/A INVX1_LOC_41/Y 0.26fF
C25987 INVX1_LOC_183/A INVX1_LOC_31/Y 0.14fF
C25988 INVX1_LOC_6/Y INVX1_LOC_58/Y 0.19fF
C25989 INVX1_LOC_176/A INVX1_LOC_487/A 0.04fF
C25990 INVX1_LOC_132/A NAND2X1_LOC_342/A 0.01fF
C25991 INVX1_LOC_513/A INVX1_LOC_114/A 0.00fF
C25992 INVX1_LOC_487/Y INVX1_LOC_48/Y 0.09fF
C25993 INVX1_LOC_41/Y INVX1_LOC_349/Y 0.02fF
C25994 INVX1_LOC_202/Y INVX1_LOC_41/Y 0.09fF
C25995 INVX1_LOC_387/Y INVX1_LOC_301/Y 0.00fF
C25996 INVX1_LOC_79/A INVX1_LOC_50/Y 0.64fF
C25997 INVX1_LOC_236/A INVX1_LOC_645/Y 0.03fF
C25998 INVX1_LOC_157/Y INVX1_LOC_245/A 0.01fF
C25999 INVX1_LOC_301/Y INVX1_LOC_49/Y 0.07fF
C26000 INVX1_LOC_100/Y NAND2X1_LOC_63/a_36_24# 0.00fF
C26001 INVX1_LOC_411/A INVX1_LOC_75/Y 0.02fF
C26002 NAND2X1_LOC_388/A INVX1_LOC_100/Y 0.08fF
C26003 INVX1_LOC_421/A INVX1_LOC_280/A 0.44fF
C26004 INVX1_LOC_387/Y INVX1_LOC_41/Y 0.01fF
C26005 INVX1_LOC_26/Y NAND2X1_LOC_759/Y 0.06fF
C26006 INVX1_LOC_351/Y INVX1_LOC_90/Y 0.03fF
C26007 NAND2X1_LOC_267/A INVX1_LOC_75/A 0.05fF
C26008 NAND2X1_LOC_242/A INVX1_LOC_275/A 0.25fF
C26009 NAND2X1_LOC_388/A INVX1_LOC_74/Y 0.03fF
C26010 INVX1_LOC_49/Y INVX1_LOC_41/Y 0.38fF
C26011 INVX1_LOC_652/A INVX1_LOC_376/Y 0.11fF
C26012 INVX1_LOC_642/Y INVX1_LOC_41/Y 0.02fF
C26013 INVX1_LOC_117/Y INVX1_LOC_636/A 0.07fF
C26014 VDD INVX1_LOC_564/A -0.00fF
C26015 INVX1_LOC_501/A INVX1_LOC_464/Y 0.01fF
C26016 INVX1_LOC_409/A NAND2X1_LOC_498/Y 0.02fF
C26017 INVX1_LOC_52/Y INVX1_LOC_578/A 0.03fF
C26018 INVX1_LOC_429/Y INVX1_LOC_429/A 0.29fF
C26019 INVX1_LOC_414/Y INVX1_LOC_217/Y 0.02fF
C26020 INVX1_LOC_584/A INVX1_LOC_584/Y 0.00fF
C26021 INVX1_LOC_203/Y INVX1_LOC_286/A 0.01fF
C26022 VDD NAND2X1_LOC_704/B 0.31fF
C26023 INVX1_LOC_41/Y INVX1_LOC_92/Y 0.00fF
C26024 NAND2X1_LOC_451/B INVX1_LOC_454/Y 0.13fF
C26025 VDD INVX1_LOC_566/Y 0.36fF
C26026 INVX1_LOC_653/Y INVX1_LOC_588/A 0.19fF
C26027 INVX1_LOC_438/Y INVX1_LOC_384/Y 0.95fF
C26028 INVX1_LOC_625/A INVX1_LOC_615/A 0.02fF
C26029 VDD INVX1_LOC_131/A -0.00fF
C26030 INVX1_LOC_206/Y INVX1_LOC_291/A 0.01fF
C26031 INVX1_LOC_413/Y INVX1_LOC_362/Y 0.03fF
C26032 INVX1_LOC_459/A INVX1_LOC_504/A 0.01fF
C26033 INVX1_LOC_551/Y INVX1_LOC_560/A 0.10fF
C26034 INVX1_LOC_17/Y INVX1_LOC_638/A 0.10fF
C26035 INVX1_LOC_412/Y INVX1_LOC_372/Y 0.01fF
C26036 INVX1_LOC_288/A INVX1_LOC_113/Y 0.06fF
C26037 INVX1_LOC_580/Y NAND2X1_LOC_122/Y 0.00fF
C26038 INVX1_LOC_68/Y NAND2X1_LOC_231/A 0.02fF
C26039 INVX1_LOC_628/Y VDD 0.21fF
C26040 VDD INVX1_LOC_626/A -0.00fF
C26041 INVX1_LOC_21/Y INVX1_LOC_32/A 0.01fF
C26042 INVX1_LOC_426/A INVX1_LOC_304/Y 0.12fF
C26043 NAND2X1_LOC_704/B INVX1_LOC_510/Y 0.01fF
C26044 VDD INVX1_LOC_432/Y 0.25fF
C26045 INVX1_LOC_203/Y NAND2X1_LOC_123/A 0.00fF
C26046 VDD INVX1_LOC_672/Y 0.21fF
C26047 VDD INVX1_LOC_367/Y 0.53fF
C26048 VDD INVX1_LOC_236/A 0.00fF
C26049 INVX1_LOC_62/A INVX1_LOC_554/A 0.01fF
C26050 INVX1_LOC_395/A INVX1_LOC_174/A 0.17fF
C26051 INPUT_0 INVX1_LOC_205/Y 0.47fF
C26052 VDD INVX1_LOC_313/Y 0.21fF
C26053 INVX1_LOC_414/A INVX1_LOC_428/Y 0.00fF
C26054 NAND2X1_LOC_498/Y INVX1_LOC_377/A 0.03fF
C26055 NAND2X1_LOC_527/a_36_24# INVX1_LOC_45/Y 0.00fF
C26056 INVX1_LOC_206/Y NAND2X1_LOC_837/B 0.04fF
C26057 NAND2X1_LOC_635/B INVX1_LOC_594/Y 0.15fF
C26058 NAND2X1_LOC_498/Y NAND2X1_LOC_595/Y 0.05fF
C26059 INVX1_LOC_578/A INVX1_LOC_115/Y 0.01fF
C26060 INVX1_LOC_584/Y INVX1_LOC_537/A 0.00fF
C26061 VDD INVX1_LOC_374/Y 0.29fF
C26062 INVX1_LOC_563/A INVX1_LOC_315/Y 0.01fF
C26063 NAND2X1_LOC_7/Y INVX1_LOC_410/A 0.06fF
C26064 INPUT_0 INVX1_LOC_194/Y 0.01fF
C26065 INVX1_LOC_34/Y INVX1_LOC_25/Y 0.09fF
C26066 INVX1_LOC_251/A INVX1_LOC_253/A 0.06fF
C26067 NAND2X1_LOC_505/a_36_24# INVX1_LOC_35/Y 0.00fF
C26068 INVX1_LOC_384/A INVX1_LOC_371/Y 0.01fF
C26069 INVX1_LOC_578/A INVX1_LOC_350/A 0.04fF
C26070 NAND2X1_LOC_498/Y INVX1_LOC_352/Y 0.03fF
C26071 INVX1_LOC_397/A INVX1_LOC_35/Y 0.57fF
C26072 INVX1_LOC_160/Y INVX1_LOC_202/Y 0.03fF
C26073 INVX1_LOC_84/A INVX1_LOC_53/Y 4.15fF
C26074 INVX1_LOC_293/Y INVX1_LOC_297/A 0.08fF
C26075 INVX1_LOC_276/A INVX1_LOC_106/A 0.00fF
C26076 INVX1_LOC_12/Y INVX1_LOC_119/A 0.01fF
C26077 INVX1_LOC_591/Y INVX1_LOC_53/Y 0.01fF
C26078 INVX1_LOC_35/Y INVX1_LOC_94/A 0.09fF
C26079 INVX1_LOC_257/Y INVX1_LOC_89/Y 0.07fF
C26080 NAND2X1_LOC_307/A INVX1_LOC_134/Y 0.03fF
C26081 NAND2X1_LOC_513/Y INPUT_1 0.00fF
C26082 INVX1_LOC_377/Y INVX1_LOC_377/A 0.09fF
C26083 INVX1_LOC_545/Y INVX1_LOC_134/Y -0.00fF
C26084 INVX1_LOC_595/Y INVX1_LOC_51/Y 0.02fF
C26085 INVX1_LOC_20/Y INVX1_LOC_186/A 0.13fF
C26086 INVX1_LOC_556/A INVX1_LOC_93/Y 0.36fF
C26087 NAND2X1_LOC_324/B INVX1_LOC_633/Y 0.37fF
C26088 NAND2X1_LOC_756/Y NAND2X1_LOC_506/a_36_24# 0.00fF
C26089 INVX1_LOC_584/Y INVX1_LOC_496/Y 0.02fF
C26090 INVX1_LOC_79/A INVX1_LOC_275/A 0.03fF
C26091 INVX1_LOC_655/Y INVX1_LOC_145/Y 0.15fF
C26092 INVX1_LOC_451/A INVX1_LOC_175/A 0.09fF
C26093 INVX1_LOC_317/Y INVX1_LOC_32/Y 0.12fF
C26094 INVX1_LOC_604/Y INVX1_LOC_97/Y 0.08fF
C26095 INVX1_LOC_613/Y NAND2X1_LOC_677/Y 0.15fF
C26096 INVX1_LOC_402/A INVX1_LOC_670/Y 0.01fF
C26097 INVX1_LOC_438/Y NAND2X1_LOC_555/B 0.05fF
C26098 INVX1_LOC_448/A INVX1_LOC_371/Y 0.00fF
C26099 INPUT_0 INVX1_LOC_44/Y 0.03fF
C26100 NAND2X1_LOC_331/A INVX1_LOC_507/A 0.01fF
C26101 INVX1_LOC_492/A INVX1_LOC_522/Y 0.01fF
C26102 INVX1_LOC_191/A INVX1_LOC_198/A 0.20fF
C26103 INVX1_LOC_587/A NAND2X1_LOC_835/a_36_24# 0.00fF
C26104 NAND2X1_LOC_677/Y NAND2X1_LOC_612/A 0.00fF
C26105 INVX1_LOC_614/A INVX1_LOC_236/A 0.03fF
C26106 INVX1_LOC_436/A INVX1_LOC_439/Y 0.06fF
C26107 NAND2X1_LOC_318/A NAND2X1_LOC_267/A 0.09fF
C26108 INVX1_LOC_381/A INVX1_LOC_117/Y 0.19fF
C26109 NAND2X1_LOC_677/Y INVX1_LOC_145/Y 0.01fF
C26110 INVX1_LOC_686/A INVX1_LOC_360/A 0.02fF
C26111 INVX1_LOC_93/Y NAND2X1_LOC_180/B 0.02fF
C26112 INVX1_LOC_45/Y INVX1_LOC_234/Y 0.06fF
C26113 INVX1_LOC_438/A INVX1_LOC_79/A 0.10fF
C26114 INVX1_LOC_276/A INVX1_LOC_239/A 0.06fF
C26115 INVX1_LOC_68/Y INVX1_LOC_77/Y 0.00fF
C26116 INVX1_LOC_193/Y INVX1_LOC_242/Y 0.02fF
C26117 NAND2X1_LOC_173/Y INVX1_LOC_261/Y 0.03fF
C26118 INVX1_LOC_523/A INVX1_LOC_9/Y 0.01fF
C26119 INVX1_LOC_137/Y INVX1_LOC_16/Y 0.02fF
C26120 INVX1_LOC_338/A INVX1_LOC_14/A 0.02fF
C26121 INVX1_LOC_80/A INVX1_LOC_105/A 0.04fF
C26122 INVX1_LOC_206/Y INVX1_LOC_657/A 0.01fF
C26123 INVX1_LOC_21/Y INVX1_LOC_202/Y 0.02fF
C26124 INVX1_LOC_288/A INVX1_LOC_501/A 0.03fF
C26125 INVX1_LOC_654/A NAND2X1_LOC_253/Y 0.04fF
C26126 INVX1_LOC_24/A INVX1_LOC_79/A 0.00fF
C26127 INVX1_LOC_438/A NAND2X1_LOC_631/B 0.60fF
C26128 INVX1_LOC_320/A INVX1_LOC_117/Y 0.02fF
C26129 VDD NAND2X1_LOC_843/B 0.02fF
C26130 INVX1_LOC_213/Y NAND2X1_LOC_499/a_36_24# 0.00fF
C26131 INVX1_LOC_400/Y INVX1_LOC_518/A 0.05fF
C26132 INVX1_LOC_632/A INVX1_LOC_50/Y 0.08fF
C26133 INVX1_LOC_366/A NAND2X1_LOC_232/a_36_24# 0.00fF
C26134 NAND2X1_LOC_666/Y INVX1_LOC_340/Y 0.01fF
C26135 INVX1_LOC_20/Y INVX1_LOC_410/A 0.01fF
C26136 INVX1_LOC_72/Y INVX1_LOC_9/Y 0.11fF
C26137 INVX1_LOC_228/Y INVX1_LOC_319/A -0.01fF
C26138 INVX1_LOC_93/Y INVX1_LOC_188/Y 0.06fF
C26139 NAND2X1_LOC_250/Y INVX1_LOC_679/A 0.03fF
C26140 INVX1_LOC_336/Y INVX1_LOC_66/A 0.01fF
C26141 INVX1_LOC_401/Y INVX1_LOC_66/A 0.01fF
C26142 INVX1_LOC_503/A INVX1_LOC_665/Y 0.01fF
C26143 INVX1_LOC_17/Y INVX1_LOC_665/Y 0.03fF
C26144 INVX1_LOC_277/A INVX1_LOC_145/Y 0.01fF
C26145 INVX1_LOC_400/A INVX1_LOC_478/Y 0.03fF
C26146 INVX1_LOC_513/Y INVX1_LOC_522/Y 0.30fF
C26147 NAND2X1_LOC_140/a_36_24# INVX1_LOC_41/Y 0.01fF
C26148 VDD INVX1_LOC_625/Y 0.28fF
C26149 INVX1_LOC_553/Y INVX1_LOC_479/A 0.01fF
C26150 INVX1_LOC_257/Y NAND2X1_LOC_544/B 0.61fF
C26151 INVX1_LOC_397/Y INVX1_LOC_97/Y 0.00fF
C26152 INVX1_LOC_59/Y INVX1_LOC_50/Y 0.01fF
C26153 VDD INVX1_LOC_91/Y 0.32fF
C26154 NAND2X1_LOC_307/A INVX1_LOC_65/A 0.00fF
C26155 INVX1_LOC_21/Y INVX1_LOC_387/Y 0.02fF
C26156 INVX1_LOC_11/Y INVX1_LOC_171/A 0.12fF
C26157 INVX1_LOC_369/A INVX1_LOC_486/A 0.01fF
C26158 INVX1_LOC_202/Y NAND2X1_LOC_267/A 0.07fF
C26159 INVX1_LOC_523/A INVX1_LOC_62/Y 0.21fF
C26160 INVX1_LOC_11/Y INVX1_LOC_105/A 0.01fF
C26161 INVX1_LOC_53/Y INVX1_LOC_496/A 0.08fF
C26162 INVX1_LOC_20/Y INVX1_LOC_124/A 0.03fF
C26163 INVX1_LOC_444/Y INVX1_LOC_46/Y 0.06fF
C26164 INVX1_LOC_554/A INVX1_LOC_76/A 0.01fF
C26165 INVX1_LOC_361/Y INVX1_LOC_371/A 0.62fF
C26166 NAND2X1_LOC_318/a_36_24# INVX1_LOC_35/Y 0.00fF
C26167 INVX1_LOC_400/A NAND2X1_LOC_387/Y 0.02fF
C26168 NAND2X1_LOC_171/a_36_24# INVX1_LOC_300/A 0.00fF
C26169 INVX1_LOC_375/A INVX1_LOC_479/A 0.03fF
C26170 NAND2X1_LOC_498/Y NAND2X1_LOC_372/Y 0.07fF
C26171 NAND2X1_LOC_498/B INVX1_LOC_41/Y 0.03fF
C26172 INVX1_LOC_617/A NAND2X1_LOC_274/B 0.03fF
C26173 INVX1_LOC_675/A INVX1_LOC_188/Y 0.07fF
C26174 NAND2X1_LOC_152/Y INVX1_LOC_655/A 0.04fF
C26175 INVX1_LOC_546/A INVX1_LOC_479/A 0.00fF
C26176 INVX1_LOC_376/A INVX1_LOC_134/Y 0.07fF
C26177 INVX1_LOC_25/Y INVX1_LOC_340/A 0.03fF
C26178 INVX1_LOC_98/A INVX1_LOC_41/Y 0.00fF
C26179 INVX1_LOC_117/Y NAND2X1_LOC_720/A 0.19fF
C26180 INVX1_LOC_50/Y INVX1_LOC_48/Y 3.98fF
C26181 INVX1_LOC_486/Y INVX1_LOC_245/A 0.02fF
C26182 INVX1_LOC_6/Y INVX1_LOC_1/Y 0.03fF
C26183 INVX1_LOC_161/A INVX1_LOC_58/Y 0.01fF
C26184 INVX1_LOC_21/Y INVX1_LOC_49/Y 0.66fF
C26185 INVX1_LOC_294/Y INVX1_LOC_245/A 0.01fF
C26186 INVX1_LOC_519/A INVX1_LOC_9/Y 0.03fF
C26187 INVX1_LOC_550/Y INVX1_LOC_555/A 0.16fF
C26188 INVX1_LOC_510/A INVX1_LOC_66/A 0.13fF
C26189 INVX1_LOC_201/Y INVX1_LOC_69/Y 0.00fF
C26190 INVX1_LOC_76/Y INVX1_LOC_41/Y 0.60fF
C26191 INVX1_LOC_110/A NAND2X1_LOC_119/a_36_24# 0.00fF
C26192 INVX1_LOC_266/A NAND2X1_LOC_109/a_36_24# 0.00fF
C26193 NAND2X1_LOC_387/Y INVX1_LOC_93/Y 0.21fF
C26194 INVX1_LOC_304/A NAND2X1_LOC_542/A 0.00fF
C26195 INVX1_LOC_166/A INVX1_LOC_32/Y 0.00fF
C26196 INVX1_LOC_187/A INVX1_LOC_79/A 0.24fF
C26197 INVX1_LOC_501/A INVX1_LOC_145/Y 0.03fF
C26198 INVX1_LOC_550/A INVX1_LOC_555/A 0.05fF
C26199 INVX1_LOC_502/A INVX1_LOC_134/Y 0.01fF
C26200 INVX1_LOC_201/A INVX1_LOC_44/Y 0.04fF
C26201 INVX1_LOC_492/A INVX1_LOC_508/A 0.06fF
C26202 INVX1_LOC_117/Y INVX1_LOC_470/Y 0.01fF
C26203 INVX1_LOC_555/A NAND2X1_LOC_213/a_36_24# 0.01fF
C26204 INVX1_LOC_51/Y INVX1_LOC_109/A 0.01fF
C26205 NAND2X1_LOC_513/A INVX1_LOC_79/A 0.02fF
C26206 INVX1_LOC_47/Y INVX1_LOC_345/A 0.10fF
C26207 INVX1_LOC_198/A INVX1_LOC_182/Y 0.02fF
C26208 INVX1_LOC_179/Y INVX1_LOC_145/Y 0.02fF
C26209 INVX1_LOC_248/A INVX1_LOC_154/A 0.01fF
C26210 INVX1_LOC_111/A INVX1_LOC_74/Y 0.01fF
C26211 NAND2X1_LOC_755/B INVX1_LOC_26/Y 0.03fF
C26212 NAND2X1_LOC_148/A INVX1_LOC_669/A 0.20fF
C26213 INVX1_LOC_602/A INVX1_LOC_74/Y 0.03fF
C26214 NAND2X1_LOC_364/a_36_24# INVX1_LOC_69/Y 0.01fF
C26215 INVX1_LOC_587/Y INVX1_LOC_659/A 0.19fF
C26216 INVX1_LOC_602/A INVX1_LOC_660/A 0.02fF
C26217 INVX1_LOC_557/Y INVX1_LOC_251/Y 0.10fF
C26218 INVX1_LOC_273/A NAND2X1_LOC_224/a_36_24# 0.00fF
C26219 INVX1_LOC_62/Y INVX1_LOC_519/A 0.17fF
C26220 INVX1_LOC_298/A INVX1_LOC_44/Y 0.03fF
C26221 INVX1_LOC_502/A INVX1_LOC_235/A 0.03fF
C26222 INVX1_LOC_69/Y NAND2X1_LOC_753/Y 0.26fF
C26223 INVX1_LOC_21/Y INVX1_LOC_92/Y 0.04fF
C26224 INVX1_LOC_54/Y INVX1_LOC_242/Y 0.07fF
C26225 NAND2X1_LOC_198/a_36_24# INVX1_LOC_63/Y 0.00fF
C26226 INVX1_LOC_119/Y INVX1_LOC_345/A 0.04fF
C26227 INVX1_LOC_63/Y NAND2X1_LOC_258/Y 0.39fF
C26228 INVX1_LOC_141/Y INVX1_LOC_501/A 0.03fF
C26229 INVX1_LOC_26/Y INVX1_LOC_46/Y 0.06fF
C26230 INVX1_LOC_117/Y INVX1_LOC_100/Y 10.77fF
C26231 INVX1_LOC_153/Y INVX1_LOC_32/Y 0.03fF
C26232 INVX1_LOC_6/Y INVX1_LOC_245/A 1.45fF
C26233 NAND2X1_LOC_843/A NAND2X1_LOC_843/B 0.08fF
C26234 NAND2X1_LOC_192/A INVX1_LOC_58/Y 0.00fF
C26235 INVX1_LOC_257/A INVX1_LOC_242/Y 0.47fF
C26236 INVX1_LOC_32/Y INVX1_LOC_531/Y 2.27fF
C26237 INVX1_LOC_442/Y INVX1_LOC_443/A 0.31fF
C26238 NAND2X1_LOC_388/A INVX1_LOC_79/A 1.92fF
C26239 INVX1_LOC_211/A INVX1_LOC_194/Y 0.09fF
C26240 NAND2X1_LOC_267/A INVX1_LOC_92/Y 0.01fF
C26241 INVX1_LOC_117/Y INVX1_LOC_74/Y 0.06fF
C26242 INVX1_LOC_518/Y NAND2X1_LOC_542/A 0.04fF
C26243 INVX1_LOC_277/Y INVX1_LOC_655/A 0.04fF
C26244 INVX1_LOC_394/Y INPUT_0 0.02fF
C26245 INVX1_LOC_454/A VDD 0.17fF
C26246 INVX1_LOC_69/Y INVX1_LOC_657/Y 0.01fF
C26247 INVX1_LOC_62/Y INVX1_LOC_659/A 0.69fF
C26248 INPUT_0 NAND2X1_LOC_58/a_36_24# 0.00fF
C26249 INVX1_LOC_193/Y INVX1_LOC_301/A 0.01fF
C26250 INVX1_LOC_662/A INVX1_LOC_669/A 0.07fF
C26251 NAND2X1_LOC_451/B INVX1_LOC_674/Y 0.01fF
C26252 VDD INVX1_LOC_393/Y 0.35fF
C26253 INVX1_LOC_44/Y INVX1_LOC_211/A 0.07fF
C26254 INVX1_LOC_601/A INVX1_LOC_207/A 0.36fF
C26255 INVX1_LOC_44/Y INVX1_LOC_64/Y 0.08fF
C26256 INVX1_LOC_447/A INVX1_LOC_578/A 0.13fF
C26257 INVX1_LOC_157/A INVX1_LOC_636/A 0.04fF
C26258 VDD INVX1_LOC_142/Y 0.21fF
C26259 NAND2X1_LOC_605/B INVX1_LOC_634/Y 0.03fF
C26260 INVX1_LOC_604/Y INVX1_LOC_615/A 0.00fF
C26261 VDD INVX1_LOC_60/Y 0.21fF
C26262 INVX1_LOC_200/Y INVX1_LOC_51/Y 0.03fF
C26263 NAND2X1_LOC_76/a_36_24# INVX1_LOC_68/Y 0.00fF
C26264 INVX1_LOC_182/A INVX1_LOC_366/A 0.01fF
C26265 INVX1_LOC_635/Y INVX1_LOC_91/Y 0.09fF
C26266 INVX1_LOC_59/Y INVX1_LOC_275/A 0.01fF
C26267 INVX1_LOC_560/A INVX1_LOC_270/A 0.00fF
C26268 INVX1_LOC_160/Y INVX1_LOC_76/Y 0.03fF
C26269 NAND2X1_LOC_45/Y INVX1_LOC_449/A 0.09fF
C26270 INVX1_LOC_577/A INVX1_LOC_187/A 0.01fF
C26271 NAND2X1_LOC_781/B INVX1_LOC_549/Y 0.18fF
C26272 NAND2X1_LOC_543/B INVX1_LOC_159/Y 0.32fF
C26273 INVX1_LOC_424/A INVX1_LOC_444/Y 0.03fF
C26274 INPUT_6 NAND2X1_LOC_17/a_36_24# 0.00fF
C26275 INVX1_LOC_410/Y INVX1_LOC_12/Y 0.07fF
C26276 NAND2X1_LOC_93/Y INVX1_LOC_59/Y 0.00fF
C26277 NAND2X1_LOC_780/B INVX1_LOC_145/Y 0.01fF
C26278 INVX1_LOC_434/A INVX1_LOC_452/A 0.11fF
C26279 INVX1_LOC_603/Y INVX1_LOC_395/A 0.02fF
C26280 INVX1_LOC_301/A INVX1_LOC_54/Y 0.02fF
C26281 INVX1_LOC_449/A NAND2X1_LOC_498/Y 0.14fF
C26282 INVX1_LOC_420/Y INVX1_LOC_442/Y 0.05fF
C26283 INVX1_LOC_84/A NAND2X1_LOC_383/Y 1.02fF
C26284 NAND2X1_LOC_93/Y INVX1_LOC_48/Y 0.03fF
C26285 INVX1_LOC_43/Y INVX1_LOC_395/A 0.01fF
C26286 INVX1_LOC_80/A INVX1_LOC_45/Y 0.20fF
C26287 VDD INVX1_LOC_164/Y 0.21fF
C26288 INVX1_LOC_613/Y INVX1_LOC_137/A 0.01fF
C26289 INVX1_LOC_607/A NAND2X1_LOC_496/Y 0.06fF
C26290 VDD NAND2X1_LOC_333/B 0.03fF
C26291 VDD INVX1_LOC_361/Y 0.30fF
C26292 INVX1_LOC_255/Y INVX1_LOC_115/A 0.01fF
C26293 INVX1_LOC_564/Y NAND2X1_LOC_755/B 0.00fF
C26294 INVX1_LOC_438/A INVX1_LOC_48/Y 0.20fF
C26295 INVX1_LOC_224/Y INVX1_LOC_411/A 0.04fF
C26296 INVX1_LOC_137/A NAND2X1_LOC_612/A 0.35fF
C26297 NAND2X1_LOC_184/Y NAND2X1_LOC_184/a_36_24# 0.02fF
C26298 INPUT_6 INPUT_4 0.03fF
C26299 INVX1_LOC_54/Y INVX1_LOC_626/Y 0.01fF
C26300 INVX1_LOC_195/A INVX1_LOC_86/Y 0.01fF
C26301 INVX1_LOC_599/A INVX1_LOC_366/A 0.01fF
C26302 INVX1_LOC_21/Y INVX1_LOC_98/A 0.14fF
C26303 INVX1_LOC_224/Y INVX1_LOC_295/Y 0.05fF
C26304 INVX1_LOC_556/A INVX1_LOC_548/A 0.00fF
C26305 NAND2X1_LOC_332/B INVX1_LOC_371/Y 0.13fF
C26306 INVX1_LOC_629/A INVX1_LOC_117/Y 0.03fF
C26307 INVX1_LOC_401/A NAND2X1_LOC_512/a_36_24# 0.02fF
C26308 INVX1_LOC_301/A INVX1_LOC_257/A 0.09fF
C26309 INVX1_LOC_290/Y INVX1_LOC_673/Y 0.20fF
C26310 INVX1_LOC_561/Y INVX1_LOC_50/Y 0.03fF
C26311 INVX1_LOC_373/A INVX1_LOC_493/A 0.01fF
C26312 INVX1_LOC_72/Y INVX1_LOC_42/Y 0.00fF
C26313 INVX1_LOC_21/Y INVX1_LOC_76/Y 0.05fF
C26314 VDD INVX1_LOC_261/Y 0.53fF
C26315 INVX1_LOC_17/Y INVX1_LOC_364/Y 0.12fF
C26316 INVX1_LOC_393/Y INVX1_LOC_103/Y 0.48fF
C26317 VDD INVX1_LOC_258/Y 0.20fF
C26318 INVX1_LOC_11/Y INVX1_LOC_45/Y 9.73fF
C26319 INVX1_LOC_395/A NAND2X1_LOC_387/Y 0.91fF
C26320 INVX1_LOC_381/A INVX1_LOC_281/Y 0.00fF
C26321 INVX1_LOC_412/Y INVX1_LOC_66/A 0.00fF
C26322 INVX1_LOC_655/Y NAND2X1_LOC_260/Y 0.01fF
C26323 NAND2X1_LOC_299/Y INVX1_LOC_633/Y 0.02fF
C26324 INVX1_LOC_20/Y NAND2X1_LOC_461/a_36_24# 0.01fF
C26325 NAND2X1_LOC_710/B INVX1_LOC_49/Y 0.02fF
C26326 INVX1_LOC_409/Y NAND2X1_LOC_274/B 0.10fF
C26327 INVX1_LOC_361/Y INVX1_LOC_510/Y 0.15fF
C26328 INVX1_LOC_182/A INVX1_LOC_6/Y 0.82fF
C26329 INVX1_LOC_601/A INVX1_LOC_79/A 0.01fF
C26330 NAND2X1_LOC_364/a_36_24# INVX1_LOC_586/A 0.00fF
C26331 NAND2X1_LOC_475/A NAND2X1_LOC_641/a_36_24# 0.00fF
C26332 INVX1_LOC_11/Y INPUT_3 0.03fF
C26333 INVX1_LOC_428/A NAND2X1_LOC_484/a_36_24# 0.00fF
C26334 INVX1_LOC_584/Y INVX1_LOC_47/Y 0.01fF
C26335 NAND2X1_LOC_45/Y INVX1_LOC_328/Y 0.55fF
C26336 INVX1_LOC_449/A INVX1_LOC_99/Y 0.07fF
C26337 INVX1_LOC_429/A NAND2X1_LOC_555/B 0.02fF
C26338 INVX1_LOC_17/Y INVX1_LOC_134/Y 0.11fF
C26339 INVX1_LOC_686/A INVX1_LOC_350/A 0.01fF
C26340 INVX1_LOC_20/Y INVX1_LOC_54/Y 0.31fF
C26341 INVX1_LOC_76/Y NAND2X1_LOC_267/A 0.09fF
C26342 INVX1_LOC_566/A INVX1_LOC_117/Y 0.07fF
C26343 INVX1_LOC_625/A NAND2X1_LOC_237/Y 0.02fF
C26344 INVX1_LOC_17/Y INVX1_LOC_47/A 0.07fF
C26345 INVX1_LOC_586/A NAND2X1_LOC_753/Y 0.02fF
C26346 NAND2X1_LOC_180/B INVX1_LOC_31/Y 0.02fF
C26347 INVX1_LOC_558/A NAND2X1_LOC_280/a_36_24# 0.00fF
C26348 INVX1_LOC_89/Y NAND2X1_LOC_332/B 0.33fF
C26349 INVX1_LOC_634/A INPUT_1 0.08fF
C26350 INVX1_LOC_205/Y INVX1_LOC_145/Y 0.02fF
C26351 INVX1_LOC_321/A INVX1_LOC_296/A 0.02fF
C26352 INVX1_LOC_187/A INVX1_LOC_48/Y 0.01fF
C26353 INVX1_LOC_394/Y INVX1_LOC_211/A 0.00fF
C26354 INVX1_LOC_53/Y INVX1_LOC_156/A 0.05fF
C26355 NAND2X1_LOC_179/Y INVX1_LOC_116/Y 0.00fF
C26356 INVX1_LOC_577/Y INVX1_LOC_49/Y 0.03fF
C26357 INVX1_LOC_617/Y INVX1_LOC_66/A 0.07fF
C26358 INVX1_LOC_17/Y NAND2X1_LOC_41/Y 0.16fF
C26359 NAND2X1_LOC_498/Y INVX1_LOC_518/A 0.15fF
C26360 INVX1_LOC_162/Y INVX1_LOC_491/A 0.03fF
C26361 INVX1_LOC_89/Y INVX1_LOC_125/Y 0.15fF
C26362 INPUT_1 INVX1_LOC_383/Y 0.01fF
C26363 NAND2X1_LOC_18/a_36_24# INVX1_LOC_26/Y 0.00fF
C26364 INVX1_LOC_455/A INVX1_LOC_25/Y 0.11fF
C26365 NAND2X1_LOC_523/B INVX1_LOC_406/A 0.03fF
C26366 INVX1_LOC_369/A INVX1_LOC_46/Y 0.00fF
C26367 INVX1_LOC_145/Y INVX1_LOC_194/Y 0.10fF
C26368 INVX1_LOC_116/Y INVX1_LOC_440/Y 0.03fF
C26369 INVX1_LOC_21/Y NAND2X1_LOC_503/Y 0.01fF
C26370 INVX1_LOC_31/Y INVX1_LOC_188/Y 0.07fF
C26371 INVX1_LOC_45/Y NAND2X1_LOC_433/Y 0.10fF
C26372 INVX1_LOC_257/Y INVX1_LOC_347/A 0.04fF
C26373 INVX1_LOC_208/Y NAND2X1_LOC_237/Y 0.00fF
C26374 INVX1_LOC_530/Y INVX1_LOC_26/Y 0.07fF
C26375 INVX1_LOC_54/Y INVX1_LOC_300/A 0.07fF
C26376 INVX1_LOC_139/A INVX1_LOC_41/Y 0.01fF
C26377 NAND2X1_LOC_271/B INVX1_LOC_75/Y 0.01fF
C26378 INVX1_LOC_197/A INVX1_LOC_69/Y 0.09fF
C26379 INVX1_LOC_599/A INVX1_LOC_6/Y 0.01fF
C26380 NAND2X1_LOC_567/a_36_24# INVX1_LOC_441/A 0.02fF
C26381 NAND2X1_LOC_97/B INVX1_LOC_255/A 0.02fF
C26382 INVX1_LOC_417/Y NAND2X1_LOC_388/A 0.18fF
C26383 INVX1_LOC_93/Y INVX1_LOC_504/Y 0.07fF
C26384 INVX1_LOC_511/Y INVX1_LOC_463/Y 0.37fF
C26385 INVX1_LOC_560/A INVX1_LOC_75/A 0.01fF
C26386 INVX1_LOC_607/Y INVX1_LOC_523/Y 0.20fF
C26387 INVX1_LOC_97/Y INVX1_LOC_63/Y 0.04fF
C26388 NAND2X1_LOC_537/a_36_24# INVX1_LOC_600/A 0.01fF
C26389 INVX1_LOC_379/Y INVX1_LOC_489/Y 0.01fF
C26390 INVX1_LOC_442/A INVX1_LOC_66/Y 0.03fF
C26391 NAND2X1_LOC_88/B INVX1_LOC_179/Y 0.01fF
C26392 INVX1_LOC_35/Y INVX1_LOC_477/Y 0.01fF
C26393 INVX1_LOC_335/A INVX1_LOC_496/Y 0.00fF
C26394 INVX1_LOC_469/Y INVX1_LOC_117/Y 0.03fF
C26395 INVX1_LOC_17/Y INVX1_LOC_65/A 0.06fF
C26396 INVX1_LOC_502/Y NAND2X1_LOC_372/Y 0.03fF
C26397 INVX1_LOC_602/A INVX1_LOC_79/A 0.09fF
C26398 INVX1_LOC_166/A INVX1_LOC_110/A 0.01fF
C26399 INVX1_LOC_617/Y NAND2X1_LOC_601/Y 0.09fF
C26400 INVX1_LOC_218/Y INVX1_LOC_6/Y 0.02fF
C26401 NAND2X1_LOC_27/Y INVX1_LOC_6/Y 0.04fF
C26402 INVX1_LOC_49/Y INVX1_LOC_481/Y 0.01fF
C26403 NAND2X1_LOC_271/B NAND2X1_LOC_271/A 0.03fF
C26404 INVX1_LOC_44/Y INVX1_LOC_145/Y 0.07fF
C26405 INVX1_LOC_69/Y NAND2X1_LOC_106/B 0.03fF
C26406 NAND2X1_LOC_791/A INVX1_LOC_44/Y 0.06fF
C26407 NAND2X1_LOC_387/Y INVX1_LOC_31/Y 0.01fF
C26408 NAND2X1_LOC_388/A INVX1_LOC_48/Y 0.04fF
C26409 INVX1_LOC_328/Y INVX1_LOC_99/Y 0.03fF
C26410 INVX1_LOC_137/Y INVX1_LOC_338/Y 0.14fF
C26411 INVX1_LOC_276/Y INVX1_LOC_662/Y 0.05fF
C26412 NAND2X1_LOC_591/Y INVX1_LOC_69/Y 0.00fF
C26413 INVX1_LOC_25/Y NAND2X1_LOC_823/Y 0.01fF
C26414 NAND2X1_LOC_286/A NAND2X1_LOC_286/a_36_24# 0.01fF
C26415 INVX1_LOC_42/Y NAND2X1_LOC_84/a_36_24# 0.00fF
C26416 INVX1_LOC_100/Y INVX1_LOC_178/A 0.02fF
C26417 INVX1_LOC_41/Y INVX1_LOC_7/Y 0.07fF
C26418 INVX1_LOC_41/Y INVX1_LOC_228/A 0.01fF
C26419 INVX1_LOC_6/Y NAND2X1_LOC_256/a_36_24# 0.00fF
C26420 INVX1_LOC_301/Y INVX1_LOC_32/Y 0.27fF
C26421 NAND2X1_LOC_615/Y INVX1_LOC_431/Y 0.01fF
C26422 INVX1_LOC_100/Y NAND2X1_LOC_76/A 0.01fF
C26423 INVX1_LOC_117/Y NAND2X1_LOC_558/B 0.02fF
C26424 NAND2X1_LOC_775/B NAND2X1_LOC_441/a_36_24# 0.00fF
C26425 INVX1_LOC_555/A NAND2X1_LOC_816/a_36_24# 0.00fF
C26426 INVX1_LOC_116/Y INVX1_LOC_66/Y 0.01fF
C26427 NAND2X1_LOC_252/a_36_24# INVX1_LOC_453/Y 0.09fF
C26428 INVX1_LOC_117/Y INVX1_LOC_79/A 8.58fF
C26429 INVX1_LOC_74/Y INVX1_LOC_251/Y 0.38fF
C26430 INVX1_LOC_608/A INVX1_LOC_100/Y 2.25fF
C26431 INVX1_LOC_47/Y INVX1_LOC_328/Y 0.07fF
C26432 NAND2X1_LOC_121/Y NAND2X1_LOC_586/Y 0.15fF
C26433 INVX1_LOC_300/Y INVX1_LOC_58/Y 0.03fF
C26434 INVX1_LOC_556/Y NAND2X1_LOC_410/Y -0.00fF
C26435 INVX1_LOC_387/Y INVX1_LOC_26/Y 0.04fF
C26436 INVX1_LOC_74/Y NAND2X1_LOC_76/A 0.01fF
C26437 INVX1_LOC_89/Y INVX1_LOC_242/Y 0.31fF
C26438 INVX1_LOC_513/A INVX1_LOC_62/Y 0.03fF
C26439 INVX1_LOC_47/Y INVX1_LOC_518/A 0.07fF
C26440 INVX1_LOC_154/A INVX1_LOC_242/Y 0.04fF
C26441 GATE_865 NAND2X1_LOC_451/B 0.03fF
C26442 INVX1_LOC_53/Y INVX1_LOC_76/A 0.01fF
C26443 INVX1_LOC_254/Y INVX1_LOC_479/A 4.53fF
C26444 INVX1_LOC_32/Y INVX1_LOC_41/Y 0.89fF
C26445 INVX1_LOC_49/Y INVX1_LOC_26/Y 0.26fF
C26446 INVX1_LOC_400/Y INVX1_LOC_109/Y 0.05fF
C26447 INVX1_LOC_49/Y INVX1_LOC_128/Y 0.09fF
C26448 INVX1_LOC_278/Y INVX1_LOC_443/A 0.45fF
C26449 INVX1_LOC_501/A INVX1_LOC_242/Y 0.03fF
C26450 INVX1_LOC_533/A INVX1_LOC_26/Y 0.06fF
C26451 INVX1_LOC_100/Y INVX1_LOC_58/Y 3.08fF
C26452 INVX1_LOC_328/Y NAND2X1_LOC_66/Y 0.03fF
C26453 INVX1_LOC_518/A INVX1_LOC_119/Y 0.03fF
C26454 INVX1_LOC_446/A INVX1_LOC_490/Y 0.01fF
C26455 INVX1_LOC_58/Y INVX1_LOC_660/A 0.03fF
C26456 INVX1_LOC_58/Y INVX1_LOC_74/Y 1.77fF
C26457 INVX1_LOC_58/Y INVX1_LOC_483/Y 0.08fF
C26458 NAND2X1_LOC_790/B INVX1_LOC_287/Y 0.02fF
C26459 INVX1_LOC_654/A INVX1_LOC_220/A 0.03fF
C26460 INVX1_LOC_224/Y INVX1_LOC_259/A 0.01fF
C26461 INVX1_LOC_412/Y INVX1_LOC_442/A 0.34fF
C26462 NAND2X1_LOC_575/a_36_24# INVX1_LOC_384/A 0.00fF
C26463 NAND2X1_LOC_525/Y INVX1_LOC_435/Y 0.10fF
C26464 INVX1_LOC_564/A INVX1_LOC_45/Y 0.00fF
C26465 INVX1_LOC_563/Y INVX1_LOC_586/A 0.01fF
C26466 INPUT_0 INVX1_LOC_425/A 0.07fF
C26467 INVX1_LOC_245/A INVX1_LOC_636/A 0.07fF
C26468 INVX1_LOC_190/A INVX1_LOC_86/A 0.10fF
C26469 INVX1_LOC_206/Y INVX1_LOC_522/Y 0.15fF
C26470 INVX1_LOC_629/A NAND2X1_LOC_798/a_36_24# 0.00fF
C26471 INVX1_LOC_560/A NAND2X1_LOC_318/A 0.01fF
C26472 VDD INVX1_LOC_307/A 0.00fF
C26473 INVX1_LOC_421/Y INVX1_LOC_406/Y 0.01fF
C26474 INVX1_LOC_255/Y INVX1_LOC_76/Y 0.03fF
C26475 INVX1_LOC_320/Y INVX1_LOC_84/A 0.03fF
C26476 INVX1_LOC_396/A INVX1_LOC_275/A 0.02fF
C26477 INVX1_LOC_626/Y NAND2X1_LOC_677/Y 0.01fF
C26478 INVX1_LOC_605/Y INVX1_LOC_395/A 0.05fF
C26479 VDD INVX1_LOC_442/Y 0.21fF
C26480 INVX1_LOC_442/A INVX1_LOC_119/A 0.05fF
C26481 INVX1_LOC_73/Y INVX1_LOC_54/Y 0.01fF
C26482 INVX1_LOC_206/Y NAND2X1_LOC_646/a_36_24# 0.01fF
C26483 INVX1_LOC_418/Y NAND2X1_LOC_322/Y 0.16fF
C26484 INVX1_LOC_404/Y NAND2X1_LOC_296/Y 0.14fF
C26485 NAND2X1_LOC_592/B INVX1_LOC_134/Y 0.01fF
C26486 NAND2X1_LOC_69/B INVX1_LOC_50/Y 0.02fF
C26487 INVX1_LOC_578/A NAND2X1_LOC_658/a_36_24# 0.00fF
C26488 INVX1_LOC_412/Y INVX1_LOC_116/Y 1.46fF
C26489 VDD INVX1_LOC_83/Y 0.33fF
C26490 NAND2X1_LOC_591/a_36_24# NAND2X1_LOC_122/Y 0.00fF
C26491 INVX1_LOC_239/Y INVX1_LOC_240/A 0.00fF
C26492 INVX1_LOC_434/A INVX1_LOC_282/A 0.18fF
C26493 INVX1_LOC_26/A INVX1_LOC_25/Y 0.00fF
C26494 NAND2X1_LOC_13/a_36_24# INVX1_LOC_270/A 0.00fF
C26495 INVX1_LOC_224/Y NAND2X1_LOC_775/B 0.03fF
C26496 VDD INVX1_LOC_578/Y 0.13fF
C26497 INVX1_LOC_63/Y INVX1_LOC_615/A 0.01fF
C26498 INVX1_LOC_51/Y INVX1_LOC_188/Y 0.01fF
C26499 NAND2X1_LOC_498/Y INVX1_LOC_352/A 0.02fF
C26500 INVX1_LOC_575/A INVX1_LOC_523/A 0.34fF
C26501 INVX1_LOC_449/A INVX1_LOC_502/Y 0.01fF
C26502 INVX1_LOC_570/A INVX1_LOC_352/A 0.01fF
C26503 INVX1_LOC_51/Y NAND2X1_LOC_411/Y 0.04fF
C26504 NAND2X1_LOC_45/Y INVX1_LOC_105/Y 0.02fF
C26505 NAND2X1_LOC_249/Y INVX1_LOC_387/Y 0.04fF
C26506 INVX1_LOC_301/A INVX1_LOC_89/Y 0.80fF
C26507 NAND2X1_LOC_756/Y INVX1_LOC_80/A 0.07fF
C26508 INVX1_LOC_578/A NAND2X1_LOC_775/B 0.10fF
C26509 NAND2X1_LOC_373/Y INVX1_LOC_257/A 0.09fF
C26510 INVX1_LOC_410/Y NAND2X1_LOC_615/B 0.01fF
C26511 INVX1_LOC_266/Y INVX1_LOC_99/Y 0.03fF
C26512 INVX1_LOC_236/A INVX1_LOC_185/Y 0.01fF
C26513 INVX1_LOC_45/Y INVX1_LOC_367/Y 0.07fF
C26514 INVX1_LOC_293/Y INVX1_LOC_80/A 0.07fF
C26515 INVX1_LOC_20/Y INVX1_LOC_371/Y 0.03fF
C26516 INVX1_LOC_20/Y NAND2X1_LOC_677/Y 0.00fF
C26517 NAND2X1_LOC_820/a_36_24# INVX1_LOC_668/A 0.00fF
C26518 INVX1_LOC_301/A NAND2X1_LOC_319/a_36_24# 0.00fF
C26519 VDD INVX1_LOC_532/Y 0.26fF
C26520 VDD INVX1_LOC_637/Y 0.21fF
C26521 NAND2X1_LOC_537/B INVX1_LOC_173/Y 0.21fF
C26522 NAND2X1_LOC_580/a_36_24# INVX1_LOC_17/Y 0.00fF
C26523 INVX1_LOC_111/A INVX1_LOC_632/A 0.05fF
C26524 INVX1_LOC_537/A NAND2X1_LOC_427/Y 0.00fF
C26525 INVX1_LOC_617/A NAND2X1_LOC_595/Y 0.01fF
C26526 INVX1_LOC_628/A NAND2X1_LOC_798/a_36_24# 0.02fF
C26527 INVX1_LOC_465/Y NAND2X1_LOC_686/A 0.00fF
C26528 INVX1_LOC_553/Y INVX1_LOC_66/A 0.02fF
C26529 NAND2X1_LOC_317/A INVX1_LOC_47/Y 0.04fF
C26530 NAND2X1_LOC_299/Y INVX1_LOC_249/A 0.06fF
C26531 INVX1_LOC_21/Y INVX1_LOC_12/A 0.01fF
C26532 INVX1_LOC_435/A INVX1_LOC_482/A 0.03fF
C26533 NAND2X1_LOC_174/a_36_24# INVX1_LOC_577/Y 0.00fF
C26534 VDD INVX1_LOC_356/Y 0.21fF
C26535 NAND2X1_LOC_387/Y NAND2X1_LOC_505/Y 0.04fF
C26536 INVX1_LOC_412/Y INVX1_LOC_255/A 0.16fF
C26537 VDD INVX1_LOC_482/Y 0.41fF
C26538 NAND2X1_LOC_311/a_36_24# INVX1_LOC_98/Y 0.00fF
C26539 INVX1_LOC_119/A INVX1_LOC_116/Y 0.02fF
C26540 INVX1_LOC_596/A NAND2X1_LOC_862/a_36_24# 0.00fF
C26541 INVX1_LOC_232/Y INVX1_LOC_134/Y 0.05fF
C26542 NAND2X1_LOC_242/A INVX1_LOC_58/Y 0.39fF
C26543 INVX1_LOC_160/Y INVX1_LOC_32/Y 1.19fF
C26544 INVX1_LOC_375/A INVX1_LOC_66/A 0.03fF
C26545 INVX1_LOC_451/A INVX1_LOC_325/Y 0.11fF
C26546 NAND2X1_LOC_387/Y INVX1_LOC_51/Y 0.50fF
C26547 INVX1_LOC_160/A INVX1_LOC_80/A 0.03fF
C26548 INVX1_LOC_522/A INVX1_LOC_512/Y 0.02fF
C26549 VDD INVX1_LOC_471/Y 0.04fF
C26550 INVX1_LOC_533/Y INVX1_LOC_89/Y 0.17fF
C26551 INVX1_LOC_543/Y INVX1_LOC_366/A 0.03fF
C26552 INVX1_LOC_604/Y NAND2X1_LOC_237/Y 0.05fF
C26553 INVX1_LOC_90/Y INVX1_LOC_388/Y 0.01fF
C26554 NAND2X1_LOC_752/a_36_24# INVX1_LOC_298/A 0.00fF
C26555 NAND2X1_LOC_475/A INVX1_LOC_328/Y 0.01fF
C26556 NAND2X1_LOC_307/A INVX1_LOC_98/Y 0.02fF
C26557 INVX1_LOC_11/Y INVX1_LOC_293/Y 4.93fF
C26558 VDD INVX1_LOC_664/Y 0.21fF
C26559 INVX1_LOC_165/Y INVX1_LOC_47/Y 0.04fF
C26560 INVX1_LOC_545/A INVX1_LOC_134/Y 0.01fF
C26561 INVX1_LOC_564/Y INVX1_LOC_49/Y 0.00fF
C26562 INVX1_LOC_29/Y INVX1_LOC_1/Y 1.37fF
C26563 INVX1_LOC_21/Y INVX1_LOC_7/Y 0.35fF
C26564 INVX1_LOC_147/A INVX1_LOC_145/Y 0.03fF
C26565 INVX1_LOC_419/Y NAND2X1_LOC_545/B 0.22fF
C26566 INVX1_LOC_508/Y INVX1_LOC_50/Y 0.03fF
C26567 INVX1_LOC_32/A NAND2X1_LOC_626/Y 0.01fF
C26568 INVX1_LOC_570/A NAND2X1_LOC_846/B 0.23fF
C26569 NAND2X1_LOC_636/A INVX1_LOC_588/A 0.01fF
C26570 NAND2X1_LOC_317/A INVX1_LOC_119/Y 0.01fF
C26571 INVX1_LOC_20/A INVX1_LOC_18/Y 0.07fF
C26572 INVX1_LOC_444/Y INVX1_LOC_386/Y 7.13fF
C26573 NAND2X1_LOC_693/a_36_24# INVX1_LOC_367/A 0.00fF
C26574 NAND2X1_LOC_770/B INVX1_LOC_53/Y 0.01fF
C26575 INPUT_2 INVX1_LOC_83/A 0.01fF
C26576 INVX1_LOC_20/Y INVX1_LOC_89/Y 0.41fF
C26577 INVX1_LOC_104/Y INVX1_LOC_48/Y 0.02fF
C26578 NAND2X1_LOC_57/Y INVX1_LOC_178/A 0.02fF
C26579 INVX1_LOC_666/A NAND2X1_LOC_52/Y 0.03fF
C26580 INVX1_LOC_254/Y INVX1_LOC_12/Y 0.64fF
C26581 INVX1_LOC_566/A INVX1_LOC_157/A 0.06fF
C26582 INVX1_LOC_11/Y INVX1_LOC_160/A 0.03fF
C26583 INVX1_LOC_301/A NAND2X1_LOC_544/B 0.05fF
C26584 INVX1_LOC_20/Y INVX1_LOC_154/A 0.03fF
C26585 INVX1_LOC_50/Y INVX1_LOC_383/Y 0.32fF
C26586 NAND2X1_LOC_24/Y INVX1_LOC_31/Y 0.03fF
C26587 INVX1_LOC_269/Y INVX1_LOC_245/A 0.38fF
C26588 INVX1_LOC_537/Y INVX1_LOC_538/A 0.01fF
C26589 INVX1_LOC_165/Y INVX1_LOC_119/Y 0.04fF
C26590 INVX1_LOC_50/Y NAND2X1_LOC_93/a_36_24# -0.00fF
C26591 INVX1_LOC_21/Y INVX1_LOC_32/Y 9.18fF
C26592 INVX1_LOC_117/Y INVX1_LOC_491/Y 0.09fF
C26593 INVX1_LOC_20/Y INVX1_LOC_501/A 0.03fF
C26594 INVX1_LOC_375/A NAND2X1_LOC_601/Y 0.01fF
C26595 NAND2X1_LOC_391/B INVX1_LOC_9/Y 0.03fF
C26596 INVX1_LOC_442/Y INVX1_LOC_103/Y 0.02fF
C26597 INVX1_LOC_117/Y INVX1_LOC_59/Y 0.06fF
C26598 INVX1_LOC_397/Y NAND2X1_LOC_237/Y 0.21fF
C26599 INVX1_LOC_267/Y INVX1_LOC_69/Y 0.04fF
C26600 INVX1_LOC_76/Y INVX1_LOC_26/Y 0.03fF
C26601 INVX1_LOC_549/A INVX1_LOC_588/A 0.01fF
C26602 INVX1_LOC_504/A INVX1_LOC_355/Y 0.01fF
C26603 INVX1_LOC_218/Y INVX1_LOC_415/Y 0.09fF
C26604 NAND2X1_LOC_97/B INVX1_LOC_69/Y 0.30fF
C26605 INVX1_LOC_381/A INVX1_LOC_245/A 0.23fF
C26606 INVX1_LOC_49/Y INVX1_LOC_369/A 0.07fF
C26607 INVX1_LOC_417/A INVX1_LOC_69/Y 0.02fF
C26608 INVX1_LOC_35/Y NAND2X1_LOC_619/Y 0.02fF
C26609 INVX1_LOC_556/Y INVX1_LOC_46/Y 0.17fF
C26610 NAND2X1_LOC_306/a_36_24# INVX1_LOC_352/A 0.00fF
C26611 INVX1_LOC_286/Y INVX1_LOC_90/Y 0.28fF
C26612 INVX1_LOC_300/A INVX1_LOC_89/Y 0.11fF
C26613 INVX1_LOC_361/Y INVX1_LOC_105/A 0.03fF
C26614 INVX1_LOC_47/Y INVX1_LOC_352/A 0.04fF
C26615 INVX1_LOC_89/Y INVX1_LOC_197/Y 0.00fF
C26616 INVX1_LOC_117/Y INVX1_LOC_48/Y 0.29fF
C26617 INVX1_LOC_81/Y INVX1_LOC_46/Y 0.02fF
C26618 INVX1_LOC_300/A INVX1_LOC_154/A 0.01fF
C26619 INVX1_LOC_93/Y INVX1_LOC_259/Y 0.74fF
C26620 INVX1_LOC_130/Y INVX1_LOC_411/Y 0.00fF
C26621 INVX1_LOC_45/Y NAND2X1_LOC_843/B 0.02fF
C26622 NAND2X1_LOC_179/Y INVX1_LOC_69/Y 0.01fF
C26623 NAND2X1_LOC_387/Y INVX1_LOC_254/A 0.03fF
C26624 INVX1_LOC_587/A INVX1_LOC_657/Y 0.01fF
C26625 INVX1_LOC_320/A INVX1_LOC_245/A 0.00fF
C26626 NAND2X1_LOC_57/Y INVX1_LOC_58/Y 0.01fF
C26627 NAND2X1_LOC_391/B INVX1_LOC_62/Y 0.02fF
C26628 INVX1_LOC_649/Y INVX1_LOC_655/A 0.04fF
C26629 INVX1_LOC_32/Y NAND2X1_LOC_267/A 0.26fF
C26630 INVX1_LOC_49/Y NAND2X1_LOC_275/Y 0.01fF
C26631 INVX1_LOC_54/Y INVX1_LOC_627/Y 0.01fF
C26632 INVX1_LOC_61/A INVX1_LOC_66/A 0.01fF
C26633 NAND2X1_LOC_184/Y INVX1_LOC_166/A 0.17fF
C26634 INVX1_LOC_360/Y INVX1_LOC_258/Y 0.34fF
C26635 INVX1_LOC_69/Y INVX1_LOC_440/Y 0.03fF
C26636 INVX1_LOC_300/A INVX1_LOC_501/A -0.07fF
C26637 INVX1_LOC_172/A INVX1_LOC_47/Y 0.12fF
C26638 INVX1_LOC_45/Y INVX1_LOC_91/Y 0.03fF
C26639 INVX1_LOC_543/Y INVX1_LOC_6/Y 0.03fF
C26640 INVX1_LOC_17/Y INVX1_LOC_351/A 0.01fF
C26641 NAND2X1_LOC_677/Y INVX1_LOC_655/A 0.03fF
C26642 INVX1_LOC_372/Y NAND2X1_LOC_118/a_36_24# 0.01fF
C26643 INVX1_LOC_229/Y INVX1_LOC_41/Y 0.01fF
C26644 INVX1_LOC_47/Y INVX1_LOC_105/Y 0.02fF
C26645 NAND2X1_LOC_375/a_36_24# INVX1_LOC_41/Y 0.00fF
C26646 NAND2X1_LOC_324/B INVX1_LOC_41/Y 0.04fF
C26647 INVX1_LOC_45/A INVX1_LOC_74/A 0.03fF
C26648 INVX1_LOC_79/A INVX1_LOC_281/Y 0.03fF
C26649 NAND2X1_LOC_513/A INVX1_LOC_614/Y 0.01fF
C26650 INVX1_LOC_93/Y INVX1_LOC_204/Y 0.02fF
C26651 INVX1_LOC_84/A INVX1_LOC_666/Y 0.07fF
C26652 INVX1_LOC_372/Y INVX1_LOC_479/A 0.01fF
C26653 INVX1_LOC_119/Y INVX1_LOC_352/A 0.10fF
C26654 INVX1_LOC_598/A INVX1_LOC_44/Y 0.03fF
C26655 INVX1_LOC_117/Y NAND2X1_LOC_491/Y 0.03fF
C26656 INVX1_LOC_17/Y INVX1_LOC_90/Y 0.10fF
C26657 NAND2X1_LOC_836/B INVX1_LOC_18/Y 0.13fF
C26658 INVX1_LOC_77/A NAND2X1_LOC_76/A 0.00fF
C26659 INVX1_LOC_382/A INVX1_LOC_379/Y 0.15fF
C26660 INVX1_LOC_100/A INVX1_LOC_63/Y 0.22fF
C26661 INVX1_LOC_670/A INVX1_LOC_9/Y 0.03fF
C26662 INVX1_LOC_277/A INVX1_LOC_655/A 0.05fF
C26663 INVX1_LOC_676/A INVX1_LOC_495/Y 0.00fF
C26664 INVX1_LOC_451/A NAND2X1_LOC_416/a_36_24# 0.09fF
C26665 INVX1_LOC_499/A INVX1_LOC_496/Y 0.03fF
C26666 INVX1_LOC_293/Y INVX1_LOC_231/Y 0.49fF
C26667 NAND2X1_LOC_503/Y INVX1_LOC_26/Y 0.01fF
C26668 NAND2X1_LOC_606/Y NAND2X1_LOC_609/B 0.00fF
C26669 INVX1_LOC_93/Y INVX1_LOC_114/A 0.04fF
C26670 NAND2X1_LOC_45/Y INVX1_LOC_109/Y 0.12fF
C26671 NAND2X1_LOC_334/B INVX1_LOC_204/Y 0.03fF
C26672 INVX1_LOC_157/A INVX1_LOC_79/A 0.03fF
C26673 INVX1_LOC_77/A INVX1_LOC_58/Y 0.01fF
C26674 NAND2X1_LOC_498/Y INVX1_LOC_109/Y 0.07fF
C26675 INVX1_LOC_675/A INVX1_LOC_114/A 0.04fF
C26676 INVX1_LOC_79/A INVX1_LOC_58/Y 0.10fF
C26677 INVX1_LOC_49/Y NAND2X1_LOC_626/Y -0.01fF
C26678 INVX1_LOC_391/A INVX1_LOC_479/A 0.02fF
C26679 VDD INVX1_LOC_570/Y 0.29fF
C26680 INVX1_LOC_69/Y NAND2X1_LOC_248/B 0.01fF
C26681 INVX1_LOC_551/A INVX1_LOC_531/Y -0.05fF
C26682 INVX1_LOC_100/Y INVX1_LOC_245/A 0.21fF
C26683 NAND2X1_LOC_837/A INVX1_LOC_91/Y 0.02fF
C26684 NAND2X1_LOC_788/A INVX1_LOC_375/A 0.04fF
C26685 INVX1_LOC_26/Y INVX1_LOC_184/Y 0.01fF
C26686 INVX1_LOC_74/Y INVX1_LOC_245/A 0.07fF
C26687 INVX1_LOC_158/A INVX1_LOC_560/A 0.05fF
C26688 INVX1_LOC_405/A NAND2X1_LOC_517/a_36_24# 0.00fF
C26689 VDD INVX1_LOC_618/Y 0.06fF
C26690 VDD NAND2X1_LOC_707/A 0.06fF
C26691 INVX1_LOC_626/Y INVX1_LOC_137/A 0.15fF
C26692 INVX1_LOC_557/A NAND2X1_LOC_317/B 0.06fF
C26693 VDD NAND2X1_LOC_493/B 0.01fF
C26694 NAND2X1_LOC_475/A INVX1_LOC_266/Y 0.02fF
C26695 INVX1_LOC_442/A INVX1_LOC_410/Y 0.07fF
C26696 INVX1_LOC_560/Y INVX1_LOC_353/Y 0.01fF
C26697 INPUT_0 INVX1_LOC_85/Y 0.02fF
C26698 INVX1_LOC_393/Y INVX1_LOC_45/Y 0.02fF
C26699 INVX1_LOC_20/Y INVX1_LOC_203/Y 0.03fF
C26700 NAND2X1_LOC_54/a_36_24# INVX1_LOC_134/Y 0.01fF
C26701 NAND2X1_LOC_596/Y NAND2X1_LOC_707/A 0.02fF
C26702 INVX1_LOC_224/Y NAND2X1_LOC_613/Y 0.01fF
C26703 INVX1_LOC_118/Y NAND2X1_LOC_332/B 0.03fF
C26704 INVX1_LOC_438/Y INVX1_LOC_406/Y 0.03fF
C26705 INVX1_LOC_95/Y INVX1_LOC_99/Y 0.06fF
C26706 VDD NAND2X1_LOC_336/B 0.58fF
C26707 NAND2X1_LOC_239/a_36_24# NAND2X1_LOC_756/Y 0.01fF
C26708 INVX1_LOC_563/Y INVX1_LOC_272/Y 0.15fF
C26709 INVX1_LOC_98/A NAND2X1_LOC_97/a_36_24# 0.00fF
C26710 NAND2X1_LOC_790/B INVX1_LOC_202/Y 0.09fF
C26711 INVX1_LOC_47/Y INVX1_LOC_109/Y 8.86fF
C26712 NAND2X1_LOC_163/B INVX1_LOC_147/Y 0.01fF
C26713 INVX1_LOC_409/Y INVX1_LOC_352/Y 0.04fF
C26714 INVX1_LOC_203/Y INVX1_LOC_300/A 0.01fF
C26715 VDD INVX1_LOC_278/Y 0.21fF
C26716 NAND2X1_LOC_39/Y NAND2X1_LOC_194/a_36_24# 0.00fF
C26717 INVX1_LOC_203/Y INVX1_LOC_197/Y 0.03fF
C26718 INVX1_LOC_257/Y INVX1_LOC_252/Y 0.07fF
C26719 INVX1_LOC_410/Y INVX1_LOC_116/Y 0.15fF
C26720 INVX1_LOC_206/Y NAND2X1_LOC_775/B 0.07fF
C26721 VDD INVX1_LOC_538/Y 0.16fF
C26722 NAND2X1_LOC_97/B INVX1_LOC_586/A 0.02fF
C26723 INVX1_LOC_76/Y INVX1_LOC_369/A 0.00fF
C26724 NAND2X1_LOC_373/Y INVX1_LOC_89/Y 0.08fF
C26725 NAND2X1_LOC_790/B INVX1_LOC_49/Y 0.01fF
C26726 INVX1_LOC_273/A NAND2X1_LOC_241/a_36_24# 0.01fF
C26727 NAND2X1_LOC_457/A INVX1_LOC_93/Y 0.03fF
C26728 INVX1_LOC_51/Y INVX1_LOC_504/Y 0.51fF
C26729 INVX1_LOC_9/A INPUT_2 0.01fF
C26730 INVX1_LOC_224/Y INVX1_LOC_490/A 0.07fF
C26731 INVX1_LOC_595/Y INVX1_LOC_33/A 0.09fF
C26732 INVX1_LOC_224/Y INVX1_LOC_317/A 0.02fF
C26733 INVX1_LOC_463/A NAND2X1_LOC_684/a_36_24# 0.00fF
C26734 INVX1_LOC_133/Y INVX1_LOC_644/Y 0.01fF
C26735 INVX1_LOC_46/Y INVX1_LOC_49/A 0.05fF
C26736 INVX1_LOC_76/Y NAND2X1_LOC_275/Y 0.02fF
C26737 VDD INVX1_LOC_379/Y 0.21fF
C26738 INVX1_LOC_586/A INVX1_LOC_440/Y 0.02fF
C26739 INVX1_LOC_412/Y INVX1_LOC_69/Y 0.05fF
C26740 VDD NAND2X1_LOC_847/A -0.00fF
C26741 INVX1_LOC_245/A NAND2X1_LOC_591/B 0.24fF
C26742 INVX1_LOC_45/Y NAND2X1_LOC_333/B 0.07fF
C26743 NAND2X1_LOC_770/A INVX1_LOC_26/Y 0.05fF
C26744 NAND2X1_LOC_537/A NAND2X1_LOC_845/B 0.03fF
C26745 INVX1_LOC_281/A INVX1_LOC_45/Y 0.01fF
C26746 INVX1_LOC_187/A INVX1_LOC_155/Y 0.08fF
C26747 INVX1_LOC_536/A INVX1_LOC_676/A 0.18fF
C26748 INVX1_LOC_395/A INVX1_LOC_204/Y 0.01fF
C26749 INVX1_LOC_308/Y INVX1_LOC_63/Y 0.01fF
C26750 INVX1_LOC_20/Y INVX1_LOC_194/Y 0.02fF
C26751 INVX1_LOC_677/Y INVX1_LOC_263/Y 0.39fF
C26752 INVX1_LOC_393/A INVX1_LOC_6/Y 0.02fF
C26753 INVX1_LOC_406/Y INVX1_LOC_219/Y 0.03fF
C26754 INVX1_LOC_525/Y NAND2X1_LOC_419/a_36_24# 0.00fF
C26755 NAND2X1_LOC_176/Y INVX1_LOC_242/Y 0.03fF
C26756 INVX1_LOC_577/Y INVX1_LOC_32/Y 0.03fF
C26757 INVX1_LOC_312/Y INVX1_LOC_510/A 0.03fF
C26758 NAND2X1_LOC_498/Y INVX1_LOC_199/Y 0.07fF
C26759 NAND2X1_LOC_148/B INVX1_LOC_133/A 0.04fF
C26760 NAND2X1_LOC_775/B INVX1_LOC_686/A 0.31fF
C26761 INVX1_LOC_84/A INVX1_LOC_431/A 0.01fF
C26762 INVX1_LOC_210/Y INVX1_LOC_80/A 0.00fF
C26763 NAND2X1_LOC_790/B INVX1_LOC_92/Y 0.05fF
C26764 INPUT_3 INVX1_LOC_281/A 0.01fF
C26765 INVX1_LOC_602/Y INVX1_LOC_685/A 0.01fF
C26766 INVX1_LOC_519/A INVX1_LOC_665/Y 1.42fF
C26767 INVX1_LOC_63/Y INVX1_LOC_624/A 0.01fF
C26768 INVX1_LOC_384/Y INVX1_LOC_6/Y 0.09fF
C26769 INVX1_LOC_207/A NAND2X1_LOC_232/a_36_24# 0.00fF
C26770 INVX1_LOC_85/Y NAND2X1_LOC_215/a_36_24# 0.00fF
C26771 INVX1_LOC_444/Y INVX1_LOC_7/Y 0.03fF
C26772 INVX1_LOC_465/Y INVX1_LOC_588/A 0.02fF
C26773 INVX1_LOC_17/Y INVX1_LOC_98/Y 0.12fF
C26774 INVX1_LOC_90/A INPUT_1 0.01fF
C26775 NAND2X1_LOC_373/Y NAND2X1_LOC_544/B 0.01fF
C26776 INVX1_LOC_421/A INVX1_LOC_53/Y 0.07fF
C26777 INVX1_LOC_617/Y INVX1_LOC_69/Y 0.07fF
C26778 INVX1_LOC_69/Y INVX1_LOC_119/A 0.00fF
C26779 INVX1_LOC_268/A INVX1_LOC_674/A 0.11fF
C26780 INVX1_LOC_47/Y INVX1_LOC_126/Y 0.01fF
C26781 INVX1_LOC_300/A INVX1_LOC_194/Y 0.00fF
C26782 INVX1_LOC_435/Y INVX1_LOC_502/A 0.10fF
C26783 INVX1_LOC_21/Y INVX1_LOC_110/A 0.00fF
C26784 NAND2X1_LOC_504/a_36_24# INVX1_LOC_600/A 0.01fF
C26785 INVX1_LOC_59/Y NAND2X1_LOC_76/A 0.01fF
C26786 INVX1_LOC_49/Y INVX1_LOC_235/Y 0.02fF
C26787 NAND2X1_LOC_65/Y INVX1_LOC_179/A 0.02fF
C26788 INVX1_LOC_20/Y INVX1_LOC_44/Y 0.20fF
C26789 INVX1_LOC_318/A NAND2X1_LOC_72/Y 0.01fF
C26790 NAND2X1_LOC_538/a_36_24# INVX1_LOC_230/A 0.01fF
C26791 INPUT_0 INVX1_LOC_505/Y 0.07fF
C26792 NAND2X1_LOC_513/A INVX1_LOC_633/A 0.01fF
C26793 NAND2X1_LOC_677/Y INVX1_LOC_627/Y 0.02fF
C26794 INVX1_LOC_511/A INVX1_LOC_58/Y 0.01fF
C26795 INVX1_LOC_437/Y INVX1_LOC_439/Y 0.04fF
C26796 INVX1_LOC_31/Y NAND2X1_LOC_423/a_36_24# 0.00fF
C26797 INVX1_LOC_651/Y INVX1_LOC_663/A 0.02fF
C26798 INVX1_LOC_248/A INVX1_LOC_252/Y 0.01fF
C26799 INVX1_LOC_444/Y INVX1_LOC_32/Y 0.08fF
C26800 INVX1_LOC_32/Y INVX1_LOC_481/Y 0.02fF
C26801 INVX1_LOC_566/A INVX1_LOC_245/A 0.07fF
C26802 INVX1_LOC_63/Y INVX1_LOC_635/A 0.02fF
C26803 NAND2X1_LOC_706/a_36_24# NAND2X1_LOC_706/B 0.01fF
C26804 INVX1_LOC_254/Y NAND2X1_LOC_615/B 0.01fF
C26805 INVX1_LOC_349/A INPUT_1 0.05fF
C26806 INVX1_LOC_573/Y INVX1_LOC_515/Y 0.02fF
C26807 NAND2X1_LOC_320/Y INVX1_LOC_47/Y 0.09fF
C26808 INVX1_LOC_35/Y INVX1_LOC_620/A 0.03fF
C26809 INVX1_LOC_612/Y INVX1_LOC_54/Y 0.01fF
C26810 INVX1_LOC_509/Y INVX1_LOC_58/Y 0.01fF
C26811 INVX1_LOC_80/A INVX1_LOC_682/A 0.00fF
C26812 INVX1_LOC_63/Y NAND2X1_LOC_237/Y 0.05fF
C26813 INVX1_LOC_68/Y INVX1_LOC_203/A 0.01fF
C26814 INVX1_LOC_677/Y INVX1_LOC_454/Y 0.00fF
C26815 INVX1_LOC_12/A INVX1_LOC_26/Y 0.02fF
C26816 INVX1_LOC_99/Y INVX1_LOC_199/Y 0.82fF
C26817 INVX1_LOC_145/Y NAND2X1_LOC_827/Y 0.10fF
C26818 INVX1_LOC_31/Y INVX1_LOC_259/Y 0.05fF
C26819 INVX1_LOC_233/Y INVX1_LOC_280/A 0.01fF
C26820 NAND2X1_LOC_779/a_36_24# INVX1_LOC_6/Y -0.00fF
C26821 INVX1_LOC_84/A NAND2X1_LOC_489/A 0.01fF
C26822 INVX1_LOC_17/Y INVX1_LOC_497/A 0.03fF
C26823 INVX1_LOC_58/Y INVX1_LOC_491/Y 0.01fF
C26824 NAND2X1_LOC_391/A INVX1_LOC_242/Y 0.46fF
C26825 NAND2X1_LOC_106/Y INVX1_LOC_54/Y 0.03fF
C26826 INVX1_LOC_376/A INVX1_LOC_504/A 0.69fF
C26827 INVX1_LOC_58/Y INVX1_LOC_59/Y 0.06fF
C26828 INVX1_LOC_300/A INVX1_LOC_44/Y 0.01fF
C26829 INVX1_LOC_402/Y INVX1_LOC_9/Y 0.01fF
C26830 INVX1_LOC_20/Y INVX1_LOC_347/A 0.10fF
C26831 INVX1_LOC_243/A INVX1_LOC_245/A 0.01fF
C26832 INVX1_LOC_63/Y INVX1_LOC_230/A 0.00fF
C26833 INVX1_LOC_157/A INVX1_LOC_48/Y 0.00fF
C26834 INVX1_LOC_44/Y INVX1_LOC_197/Y 0.07fF
C26835 INVX1_LOC_359/Y INVX1_LOC_372/A 0.09fF
C26836 INVX1_LOC_193/Y INVX1_LOC_92/A 0.01fF
C26837 INVX1_LOC_194/A INVX1_LOC_390/A 0.06fF
C26838 INVX1_LOC_26/Y INVX1_LOC_7/Y 2.07fF
C26839 INVX1_LOC_435/A INVX1_LOC_9/Y 0.16fF
C26840 INVX1_LOC_58/Y INVX1_LOC_48/Y 0.24fF
C26841 INVX1_LOC_421/A NAND2X1_LOC_346/B 0.15fF
C26842 NAND2X1_LOC_299/Y INVX1_LOC_41/Y 0.12fF
C26843 INVX1_LOC_293/Y NAND2X1_LOC_843/B 0.00fF
C26844 NAND2X1_LOC_320/Y INVX1_LOC_119/Y 0.00fF
C26845 INVX1_LOC_31/Y INVX1_LOC_204/Y 0.55fF
C26846 INVX1_LOC_17/Y NAND2X1_LOC_41/a_36_24# 0.00fF
C26847 INVX1_LOC_674/A NAND2X1_LOC_719/A 0.05fF
C26848 INVX1_LOC_47/Y INVX1_LOC_199/Y 0.15fF
C26849 NAND2X1_LOC_605/a_36_24# INVX1_LOC_347/A 0.00fF
C26850 NAND2X1_LOC_557/B INVX1_LOC_199/Y 0.16fF
C26851 INVX1_LOC_435/A INVX1_LOC_62/Y 0.04fF
C26852 INVX1_LOC_32/Y INVX1_LOC_26/Y 0.27fF
C26853 INVX1_LOC_31/Y INVX1_LOC_114/A 0.11fF
C26854 INVX1_LOC_160/A INVX1_LOC_625/Y 0.01fF
C26855 NAND2X1_LOC_184/Y INVX1_LOC_41/Y 0.74fF
C26856 INVX1_LOC_479/A NAND2X1_LOC_615/B 0.02fF
C26857 INVX1_LOC_199/Y INVX1_LOC_119/Y 0.03fF
C26858 INVX1_LOC_560/A INVX1_LOC_192/A 0.04fF
C26859 INVX1_LOC_505/Y INVX1_LOC_498/A 0.23fF
C26860 INVX1_LOC_399/A INVX1_LOC_399/Y -0.00fF
C26861 INVX1_LOC_491/A INVX1_LOC_196/Y 0.03fF
C26862 INVX1_LOC_97/A NAND2X1_LOC_86/Y 0.02fF
C26863 NAND2X1_LOC_558/B INVX1_LOC_245/A 0.01fF
C26864 INVX1_LOC_301/A NAND2X1_LOC_176/Y 0.05fF
C26865 INVX1_LOC_479/A INVX1_LOC_66/A 0.10fF
C26866 INVX1_LOC_79/A NAND2X1_LOC_440/A 0.03fF
C26867 INVX1_LOC_79/A INVX1_LOC_245/A 0.13fF
C26868 INVX1_LOC_75/Y INVX1_LOC_411/Y 0.09fF
C26869 INVX1_LOC_459/A INVX1_LOC_374/A 0.02fF
C26870 NAND2X1_LOC_631/B INVX1_LOC_245/A 0.04fF
C26871 INVX1_LOC_54/Y INVX1_LOC_92/A 0.04fF
C26872 NAND2X1_LOC_396/Y INVX1_LOC_245/A 0.14fF
C26873 VDD INVX1_LOC_215/Y 0.21fF
C26874 INPUT_6 INVX1_LOC_1/A 0.80fF
C26875 NAND2X1_LOC_790/B INVX1_LOC_98/A 0.02fF
C26876 INVX1_LOC_114/A INVX1_LOC_473/Y 0.02fF
C26877 NAND2X1_LOC_790/B INVX1_LOC_76/Y 0.11fF
C26878 INVX1_LOC_395/A NAND2X1_LOC_100/a_36_24# 0.00fF
C26879 INVX1_LOC_479/A NAND2X1_LOC_601/Y 0.05fF
C26880 INVX1_LOC_554/A INVX1_LOC_136/Y 0.02fF
C26881 INVX1_LOC_206/Y INVX1_LOC_169/A 0.06fF
C26882 INVX1_LOC_20/Y INVX1_LOC_118/Y 0.06fF
C26883 INVX1_LOC_84/A INVX1_LOC_54/A 0.09fF
C26884 INVX1_LOC_395/A INVX1_LOC_482/A 0.01fF
C26885 INVX1_LOC_41/Y NAND2X1_LOC_271/A 0.26fF
C26886 INPUT_0 INVX1_LOC_80/A 1.05fF
C26887 VDD INVX1_LOC_321/Y 0.04fF
C26888 INVX1_LOC_3/Y INVX1_LOC_1/Y 0.37fF
C26889 INVX1_LOC_412/Y NAND2X1_LOC_808/a_36_24# 0.00fF
C26890 INVX1_LOC_617/Y INVX1_LOC_586/A 0.10fF
C26891 INVX1_LOC_578/A INVX1_LOC_249/A 0.23fF
C26892 INVX1_LOC_586/A INVX1_LOC_119/A 0.01fF
C26893 NAND2X1_LOC_781/B INVX1_LOC_186/Y 0.02fF
C26894 NAND2X1_LOC_498/Y INVX1_LOC_53/Y 0.24fF
C26895 INVX1_LOC_570/A INVX1_LOC_53/Y 0.03fF
C26896 NAND2X1_LOC_332/B INVX1_LOC_126/A 0.01fF
C26897 NAND2X1_LOC_832/A NAND2X1_LOC_449/a_36_24# 0.00fF
C26898 INVX1_LOC_76/Y INVX1_LOC_235/Y 0.45fF
C26899 INVX1_LOC_95/Y INVX1_LOC_96/A 0.02fF
C26900 INVX1_LOC_581/A INVX1_LOC_143/Y 0.03fF
C26901 INVX1_LOC_364/Y INVX1_LOC_519/A 0.01fF
C26902 NAND2X1_LOC_249/Y INVX1_LOC_32/Y 0.02fF
C26903 INVX1_LOC_395/A INVX1_LOC_194/A 0.01fF
C26904 INVX1_LOC_435/Y INVX1_LOC_17/Y 0.10fF
C26905 INPUT_0 INVX1_LOC_11/Y 0.24fF
C26906 INVX1_LOC_20/Y INVX1_LOC_312/A 0.03fF
C26907 INVX1_LOC_20/Y NAND2X1_LOC_391/A 0.03fF
C26908 INVX1_LOC_617/Y INVX1_LOC_312/Y 0.07fF
C26909 INVX1_LOC_442/Y INVX1_LOC_45/Y 0.10fF
C26910 NAND2X1_LOC_43/a_36_24# INVX1_LOC_6/Y 0.00fF
C26911 INVX1_LOC_96/Y INVX1_LOC_197/Y 0.42fF
C26912 INVX1_LOC_459/Y INVX1_LOC_99/Y 0.58fF
C26913 INVX1_LOC_11/Y NAND2X1_LOC_516/Y 0.49fF
C26914 INVX1_LOC_85/Y INVX1_LOC_145/Y 0.47fF
C26915 NAND2X1_LOC_692/Y INVX1_LOC_45/Y 0.01fF
C26916 INVX1_LOC_20/Y INVX1_LOC_147/A 0.05fF
C26917 INVX1_LOC_686/A INVX1_LOC_633/Y 0.04fF
C26918 INVX1_LOC_409/Y INVX1_LOC_347/Y 0.01fF
C26919 INVX1_LOC_206/Y INVX1_LOC_317/A 0.03fF
C26920 NAND2X1_LOC_457/A INVX1_LOC_31/Y 0.02fF
C26921 INVX1_LOC_133/A INVX1_LOC_241/Y 0.09fF
C26922 INVX1_LOC_510/Y NAND2X1_LOC_317/a_36_24# 0.00fF
C26923 VDD INVX1_LOC_77/Y 0.25fF
C26924 INVX1_LOC_560/A INVX1_LOC_32/Y 0.07fF
C26925 INVX1_LOC_254/Y INVX1_LOC_442/A 0.01fF
C26926 INVX1_LOC_134/Y INVX1_LOC_519/A 0.01fF
C26927 INVX1_LOC_395/A INVX1_LOC_87/Y 0.01fF
C26928 NAND2X1_LOC_475/A INVX1_LOC_199/Y 0.08fF
C26929 INVX1_LOC_51/Y INVX1_LOC_259/Y 0.09fF
C26930 INVX1_LOC_564/Y INVX1_LOC_32/Y 0.00fF
C26931 INVX1_LOC_556/Y INVX1_LOC_76/Y 0.06fF
C26932 INVX1_LOC_166/A INVX1_LOC_557/A 0.03fF
C26933 INVX1_LOC_609/Y INVX1_LOC_581/A 0.03fF
C26934 INVX1_LOC_410/Y INVX1_LOC_69/Y 0.03fF
C26935 INVX1_LOC_596/A INVX1_LOC_503/A 0.12fF
C26936 INVX1_LOC_291/A INVX1_LOC_35/Y 0.06fF
C26937 INVX1_LOC_673/A NAND2X1_LOC_852/a_36_24# 0.00fF
C26938 NAND2X1_LOC_517/Y NAND2X1_LOC_416/Y 0.00fF
C26939 INVX1_LOC_369/A INVX1_LOC_7/Y 0.00fF
C26940 INVX1_LOC_292/A INVX1_LOC_63/Y 0.01fF
C26941 INVX1_LOC_375/A INVX1_LOC_69/Y 0.03fF
C26942 INVX1_LOC_53/Y INVX1_LOC_99/Y 0.32fF
C26943 INVX1_LOC_607/Y INVX1_LOC_80/A 0.18fF
C26944 INVX1_LOC_545/A NAND2X1_LOC_545/B 0.01fF
C26945 INVX1_LOC_366/A NAND2X1_LOC_204/a_36_24# 0.01fF
C26946 INPUT_3 INVX1_LOC_83/Y 0.03fF
C26947 INVX1_LOC_607/Y NAND2X1_LOC_768/A 0.12fF
C26948 INVX1_LOC_76/Y INVX1_LOC_506/A 0.08fF
C26949 NAND2X1_LOC_457/A INVX1_LOC_682/Y 0.01fF
C26950 INVX1_LOC_274/A INVX1_LOC_600/A 0.02fF
C26951 INVX1_LOC_84/A NAND2X1_LOC_84/B 0.15fF
C26952 INVX1_LOC_599/Y INVX1_LOC_145/Y 0.02fF
C26953 INVX1_LOC_587/Y INVX1_LOC_59/A 0.01fF
C26954 INVX1_LOC_51/Y INVX1_LOC_204/Y 0.03fF
C26955 INVX1_LOC_577/A INVX1_LOC_245/A 0.01fF
C26956 INVX1_LOC_295/A INVX1_LOC_295/Y 0.05fF
C26957 INVX1_LOC_574/Y INVX1_LOC_575/Y 0.01fF
C26958 INVX1_LOC_117/Y INVX1_LOC_508/Y 0.01fF
C26959 INVX1_LOC_420/Y NAND2X1_LOC_274/B 0.08fF
C26960 INVX1_LOC_531/A INVX1_LOC_35/Y 0.01fF
C26961 NAND2X1_LOC_156/Y INVX1_LOC_145/Y 0.01fF
C26962 INVX1_LOC_325/Y INVX1_LOC_326/A 0.00fF
C26963 NAND2X1_LOC_65/Y INVX1_LOC_69/Y 0.17fF
C26964 INVX1_LOC_291/A INVX1_LOC_620/A 0.26fF
C26965 INVX1_LOC_45/Y INVX1_LOC_356/Y 0.02fF
C26966 INVX1_LOC_12/Y NAND2X1_LOC_615/B 0.03fF
C26967 INVX1_LOC_54/Y INVX1_LOC_679/Y 0.10fF
C26968 NAND2X1_LOC_866/a_36_24# INVX1_LOC_632/A 0.00fF
C26969 INVX1_LOC_32/Y INVX1_LOC_369/A 0.03fF
C26970 INVX1_LOC_406/Y INVX1_LOC_69/Y 0.03fF
C26971 INVX1_LOC_612/Y NAND2X1_LOC_677/Y 0.06fF
C26972 NAND2X1_LOC_788/A INVX1_LOC_479/A 0.02fF
C26973 NAND2X1_LOC_787/a_36_24# INVX1_LOC_35/Y 0.00fF
C26974 NAND2X1_LOC_302/a_36_24# INVX1_LOC_93/Y 0.01fF
C26975 INVX1_LOC_188/Y INVX1_LOC_359/A 0.01fF
C26976 INVX1_LOC_460/Y INVX1_LOC_99/Y 0.12fF
C26977 INVX1_LOC_35/Y NAND2X1_LOC_837/B 0.01fF
C26978 INVX1_LOC_678/A NAND2X1_LOC_857/a_36_24# 0.02fF
C26979 INVX1_LOC_21/Y NAND2X1_LOC_184/Y 0.03fF
C26980 INVX1_LOC_117/Y INVX1_LOC_155/Y 0.03fF
C26981 INVX1_LOC_522/Y INVX1_LOC_139/Y 0.05fF
C26982 INVX1_LOC_447/Y INPUT_1 0.52fF
C26983 NAND2X1_LOC_638/A NAND2X1_LOC_821/a_36_24# 0.00fF
C26984 INVX1_LOC_176/A INVX1_LOC_50/Y 0.07fF
C26985 INVX1_LOC_53/Y INVX1_LOC_47/Y 0.26fF
C26986 INVX1_LOC_639/Y INVX1_LOC_641/Y 0.00fF
C26987 INVX1_LOC_12/Y INVX1_LOC_66/A 0.65fF
C26988 INVX1_LOC_679/A INVX1_LOC_221/Y 0.01fF
C26989 INVX1_LOC_51/Y INVX1_LOC_114/A 0.22fF
C26990 INVX1_LOC_459/Y INVX1_LOC_119/Y 0.01fF
C26991 INVX1_LOC_425/A INVX1_LOC_242/Y 0.73fF
C26992 INVX1_LOC_616/A INVX1_LOC_26/Y 0.01fF
C26993 NAND2X1_LOC_602/A INPUT_1 0.01fF
C26994 INVX1_LOC_636/A INVX1_LOC_458/Y 0.01fF
C26995 INVX1_LOC_34/Y INVX1_LOC_25/A 0.01fF
C26996 INVX1_LOC_99/Y NAND2X1_LOC_346/B 0.03fF
C26997 NAND2X1_LOC_148/B INVX1_LOC_662/Y 0.00fF
C26998 INVX1_LOC_304/Y INVX1_LOC_46/Y 0.03fF
C26999 INVX1_LOC_367/A INVX1_LOC_9/Y 0.03fF
C27000 INVX1_LOC_556/Y INVX1_LOC_108/A 0.09fF
C27001 INVX1_LOC_392/Y INVX1_LOC_62/Y 0.09fF
C27002 INVX1_LOC_54/Y INPUT_1 0.72fF
C27003 INVX1_LOC_384/A INVX1_LOC_665/A 0.04fF
C27004 INVX1_LOC_99/Y NAND2X1_LOC_274/Y 0.01fF
C27005 INVX1_LOC_442/A INVX1_LOC_479/A 0.09fF
C27006 INPUT_0 INVX1_LOC_231/Y 0.03fF
C27007 INVX1_LOC_467/Y INVX1_LOC_466/A 0.06fF
C27008 INVX1_LOC_632/A INVX1_LOC_245/A 0.08fF
C27009 INVX1_LOC_543/Y NAND2X1_LOC_789/A 0.02fF
C27010 NAND2X1_LOC_775/B NAND2X1_LOC_542/A 0.02fF
C27011 INVX1_LOC_53/Y INVX1_LOC_119/Y 0.06fF
C27012 INVX1_LOC_240/A NAND2X1_LOC_286/a_36_24# 0.00fF
C27013 NAND2X1_LOC_355/A GATE_865 0.03fF
C27014 NAND2X1_LOC_720/A NAND2X1_LOC_753/Y 0.02fF
C27015 INVX1_LOC_99/Y NAND2X1_LOC_406/B 0.01fF
C27016 INVX1_LOC_53/Y NAND2X1_LOC_66/Y 0.03fF
C27017 INVX1_LOC_62/Y INVX1_LOC_59/A 0.03fF
C27018 INVX1_LOC_254/Y INVX1_LOC_255/A 0.00fF
C27019 INVX1_LOC_257/A INPUT_1 0.07fF
C27020 INVX1_LOC_300/Y INVX1_LOC_678/A 0.01fF
C27021 INVX1_LOC_396/A INVX1_LOC_58/Y 0.16fF
C27022 INVX1_LOC_367/A INVX1_LOC_62/Y 0.07fF
C27023 NAND2X1_LOC_570/a_36_24# NAND2X1_LOC_555/B 0.00fF
C27024 INVX1_LOC_59/Y INVX1_LOC_245/A 0.02fF
C27025 NAND2X1_LOC_128/A INVX1_LOC_6/Y 0.35fF
C27026 INVX1_LOC_7/Y NAND2X1_LOC_626/Y 0.46fF
C27027 NAND2X1_LOC_852/a_36_24# INVX1_LOC_660/Y 0.00fF
C27028 INVX1_LOC_242/Y INVX1_LOC_252/Y 0.08fF
C27029 INVX1_LOC_26/Y NAND2X1_LOC_226/Y 0.01fF
C27030 NAND2X1_LOC_127/a_36_24# INVX1_LOC_6/Y 0.00fF
C27031 INVX1_LOC_63/Y NAND2X1_LOC_482/Y 0.92fF
C27032 INVX1_LOC_587/Y NAND2X1_LOC_334/B 0.02fF
C27033 NAND2X1_LOC_274/B INVX1_LOC_371/A 0.16fF
C27034 INVX1_LOC_665/A INVX1_LOC_145/Y 0.01fF
C27035 INVX1_LOC_48/Y INVX1_LOC_245/A 0.14fF
C27036 INVX1_LOC_183/A INVX1_LOC_46/Y 0.03fF
C27037 INVX1_LOC_80/A INVX1_LOC_211/A 0.23fF
C27038 INVX1_LOC_12/Y NAND2X1_LOC_621/B 0.03fF
C27039 INVX1_LOC_21/Y INVX1_LOC_75/Y 0.07fF
C27040 INVX1_LOC_62/Y INVX1_LOC_516/A 0.02fF
C27041 INVX1_LOC_11/Y NAND2X1_LOC_495/a_36_24# 0.00fF
C27042 INVX1_LOC_93/Y INVX1_LOC_9/Y 0.03fF
C27043 INVX1_LOC_460/Y INVX1_LOC_119/Y 0.02fF
C27044 NAND2X1_LOC_555/B NAND2X1_LOC_294/Y 0.09fF
C27045 INVX1_LOC_505/Y INVX1_LOC_145/Y 0.19fF
C27046 INVX1_LOC_198/Y INVX1_LOC_207/Y 0.07fF
C27047 INVX1_LOC_389/Y INVX1_LOC_46/Y 0.01fF
C27048 INVX1_LOC_479/A INVX1_LOC_116/Y 0.07fF
C27049 INVX1_LOC_392/A INVX1_LOC_62/Y 0.05fF
C27050 INVX1_LOC_81/Y INVX1_LOC_184/Y 0.01fF
C27051 INVX1_LOC_32/Y NAND2X1_LOC_626/Y 0.00fF
C27052 INVX1_LOC_6/Y INVX1_LOC_485/Y 0.01fF
C27053 INVX1_LOC_137/Y INVX1_LOC_588/A 0.04fF
C27054 INVX1_LOC_479/A NAND2X1_LOC_432/Y 0.01fF
C27055 INVX1_LOC_17/Y INVX1_LOC_346/Y 0.22fF
C27056 INVX1_LOC_379/A INVX1_LOC_488/Y 0.01fF
C27057 INVX1_LOC_11/Y INVX1_LOC_211/A 0.01fF
C27058 NAND2X1_LOC_409/Y INVX1_LOC_18/Y 0.04fF
C27059 INVX1_LOC_93/Y INVX1_LOC_62/Y 0.40fF
C27060 NAND2X1_LOC_491/Y INVX1_LOC_245/A 0.01fF
C27061 INVX1_LOC_680/A INVX1_LOC_66/A 0.01fF
C27062 NAND2X1_LOC_294/Y NAND2X1_LOC_395/Y 0.09fF
C27063 INVX1_LOC_390/A INVX1_LOC_9/Y 0.02fF
C27064 INVX1_LOC_26/Y NAND2X1_LOC_275/a_36_24# 0.00fF
C27065 INVX1_LOC_293/A INVX1_LOC_100/Y 0.00fF
C27066 INVX1_LOC_181/A NAND2X1_LOC_205/a_36_24# 0.00fF
C27067 INVX1_LOC_93/Y INVX1_LOC_529/Y 0.03fF
C27068 INVX1_LOC_6/Y NAND2X1_LOC_248/B 0.00fF
C27069 INVX1_LOC_513/Y INVX1_LOC_41/Y 0.12fF
C27070 INVX1_LOC_662/A NAND2X1_LOC_814/a_36_24# 0.01fF
C27071 NAND2X1_LOC_387/Y INVX1_LOC_291/Y 0.03fF
C27072 INVX1_LOC_675/A INVX1_LOC_62/Y 0.07fF
C27073 INVX1_LOC_255/A INVX1_LOC_479/A 0.07fF
C27074 NAND2X1_LOC_174/B INVX1_LOC_636/A 0.00fF
C27075 INVX1_LOC_390/A INVX1_LOC_62/Y 0.03fF
C27076 INVX1_LOC_89/Y INVX1_LOC_270/Y 0.00fF
C27077 INVX1_LOC_47/Y NAND2X1_LOC_60/Y 0.06fF
C27078 INVX1_LOC_369/Y INVX1_LOC_280/A 0.02fF
C27079 INVX1_LOC_89/Y INVX1_LOC_92/A 0.27fF
C27080 INVX1_LOC_425/A INVX1_LOC_301/A 0.52fF
C27081 INVX1_LOC_139/A INVX1_LOC_373/A 0.00fF
C27082 INVX1_LOC_100/Y INVX1_LOC_483/A 0.01fF
C27083 INVX1_LOC_317/Y INVX1_LOC_206/Y 0.55fF
C27084 INVX1_LOC_657/Y INVX1_LOC_660/A 0.15fF
C27085 INVX1_LOC_200/Y INVX1_LOC_558/A 0.01fF
C27086 NAND2X1_LOC_457/A INVX1_LOC_51/Y 1.30fF
C27087 INVX1_LOC_74/Y INVX1_LOC_652/Y 0.01fF
C27088 INVX1_LOC_410/Y INVX1_LOC_586/A 0.03fF
C27089 INVX1_LOC_375/A INVX1_LOC_586/A 0.03fF
C27090 INPUT_0 NAND2X1_LOC_704/B 0.12fF
C27091 INVX1_LOC_483/A INVX1_LOC_483/Y 0.18fF
C27092 INVX1_LOC_45/Y NAND2X1_LOC_707/A 0.03fF
C27093 INVX1_LOC_555/Y INVX1_LOC_570/A 0.04fF
C27094 NAND2X1_LOC_69/B INVX1_LOC_178/A 0.00fF
C27095 INVX1_LOC_257/Y INVX1_LOC_80/A 0.28fF
C27096 INVX1_LOC_68/Y INVX1_LOC_266/Y 0.31fF
C27097 INVX1_LOC_312/Y INVX1_LOC_410/Y 0.05fF
C27098 VDD INVX1_LOC_549/Y 0.14fF
C27099 INVX1_LOC_406/Y INVX1_LOC_586/A 0.03fF
C27100 INVX1_LOC_20/Y INVX1_LOC_425/A 0.03fF
C27101 INVX1_LOC_118/Y NAND2X1_LOC_140/B 0.02fF
C27102 INVX1_LOC_255/Y NAND2X1_LOC_299/Y 0.01fF
C27103 NAND2X1_LOC_544/B INVX1_LOC_92/A 0.04fF
C27104 NAND2X1_LOC_536/a_36_24# INVX1_LOC_600/A 0.02fF
C27105 NAND2X1_LOC_790/B INVX1_LOC_32/Y 0.07fF
C27106 INVX1_LOC_65/Y NAND2X1_LOC_307/A 0.51fF
C27107 NAND2X1_LOC_727/a_36_24# INVX1_LOC_80/A 0.01fF
C27108 INVX1_LOC_11/Y INVX1_LOC_257/Y 0.07fF
C27109 NAND2X1_LOC_253/Y INVX1_LOC_220/A 0.20fF
C27110 INVX1_LOC_612/Y NAND2X1_LOC_780/B 0.09fF
C27111 INVX1_LOC_71/Y INVX1_LOC_6/Y 0.01fF
C27112 INPUT_0 INVX1_LOC_313/Y 0.02fF
C27113 INVX1_LOC_384/A INVX1_LOC_80/A 0.07fF
C27114 INVX1_LOC_266/Y INVX1_LOC_600/A 0.07fF
C27115 INVX1_LOC_588/Y INVX1_LOC_206/Y 0.01fF
C27116 INVX1_LOC_21/A INPUT_2 0.22fF
C27117 VDD INVX1_LOC_463/Y 0.51fF
C27118 VDD INVX1_LOC_372/A -0.00fF
C27119 NAND2X1_LOC_370/A INVX1_LOC_98/Y 0.02fF
C27120 NAND2X1_LOC_69/B INVX1_LOC_58/Y 0.68fF
C27121 INVX1_LOC_11/Y INVX1_LOC_446/Y 0.24fF
C27122 INVX1_LOC_439/Y INVX1_LOC_445/Y 0.05fF
C27123 NAND2X1_LOC_636/A INVX1_LOC_496/A 0.03fF
C27124 INVX1_LOC_166/A INVX1_LOC_206/Y 0.08fF
C27125 INVX1_LOC_551/Y NAND2X1_LOC_411/Y 0.22fF
C27126 INVX1_LOC_564/A INVX1_LOC_298/A 0.02fF
C27127 INVX1_LOC_373/A INVX1_LOC_32/Y 0.03fF
C27128 INVX1_LOC_362/Y INVX1_LOC_303/Y 0.05fF
C27129 INVX1_LOC_53/Y INVX1_LOC_136/Y 0.02fF
C27130 INVX1_LOC_291/A NAND2X1_LOC_664/a_36_24# 0.02fF
C27131 INVX1_LOC_293/Y INVX1_LOC_442/Y 0.07fF
C27132 INVX1_LOC_11/Y INVX1_LOC_384/A 0.07fF
C27133 INVX1_LOC_586/A INVX1_LOC_674/A 0.07fF
C27134 INVX1_LOC_54/Y INVX1_LOC_134/A 0.00fF
C27135 INVX1_LOC_404/Y NAND2X1_LOC_520/A 0.01fF
C27136 INVX1_LOC_448/A INVX1_LOC_80/A 0.07fF
C27137 NAND2X1_LOC_184/Y NAND2X1_LOC_526/a_36_24# 0.00fF
C27138 INVX1_LOC_224/Y INVX1_LOC_411/Y 0.03fF
C27139 INVX1_LOC_370/Y INVX1_LOC_519/A 0.02fF
C27140 INVX1_LOC_84/A INVX1_LOC_230/A 0.17fF
C27141 INVX1_LOC_677/Y GATE_865 0.38fF
C27142 INVX1_LOC_549/A INVX1_LOC_496/A 0.09fF
C27143 NAND2X1_LOC_190/a_36_24# INVX1_LOC_362/Y 0.00fF
C27144 INVX1_LOC_63/Y NAND2X1_LOC_749/Y 0.05fF
C27145 INVX1_LOC_12/Y INVX1_LOC_305/Y 0.91fF
C27146 NAND2X1_LOC_475/A NAND2X1_LOC_406/B 0.11fF
C27147 INVX1_LOC_523/A INVX1_LOC_476/A 0.21fF
C27148 INVX1_LOC_80/A INVX1_LOC_145/Y 0.15fF
C27149 VDD NAND2X1_LOC_274/B 0.01fF
C27150 NAND2X1_LOC_107/Y INVX1_LOC_99/Y 0.19fF
C27151 NAND2X1_LOC_768/A INVX1_LOC_145/Y 0.01fF
C27152 INVX1_LOC_166/A INVX1_LOC_242/A 1.24fF
C27153 INVX1_LOC_578/A INVX1_LOC_411/Y 0.02fF
C27154 INVX1_LOC_588/Y INVX1_LOC_686/A 0.07fF
C27155 INVX1_LOC_32/Y INVX1_LOC_235/Y 0.07fF
C27156 INVX1_LOC_395/A INVX1_LOC_9/Y 0.26fF
C27157 INVX1_LOC_293/Y INVX1_LOC_671/A 0.02fF
C27158 INVX1_LOC_561/Y INVX1_LOC_245/A 0.03fF
C27159 NAND2X1_LOC_383/Y INVX1_LOC_47/Y 0.10fF
C27160 NAND2X1_LOC_122/Y INVX1_LOC_497/A 0.18fF
C27161 NAND2X1_LOC_673/B INVX1_LOC_307/A 0.02fF
C27162 INVX1_LOC_599/A INVX1_LOC_48/Y 0.01fF
C27163 NAND2X1_LOC_506/a_36_24# INVX1_LOC_197/Y 0.01fF
C27164 INVX1_LOC_277/A INVX1_LOC_679/Y 0.01fF
C27165 VDD INVX1_LOC_148/Y 0.21fF
C27166 NAND2X1_LOC_831/a_36_24# INVX1_LOC_376/Y 0.00fF
C27167 INVX1_LOC_530/Y INVX1_LOC_183/A 0.28fF
C27168 INVX1_LOC_596/A INVX1_LOC_230/Y 0.29fF
C27169 INVX1_LOC_81/Y INVX1_LOC_7/Y 0.03fF
C27170 INVX1_LOC_570/A INVX1_LOC_662/A 0.14fF
C27171 INVX1_LOC_176/Y INVX1_LOC_6/Y 0.14fF
C27172 INVX1_LOC_206/Y INVX1_LOC_531/Y 1.97fF
C27173 INVX1_LOC_224/Y INVX1_LOC_41/Y 0.03fF
C27174 INVX1_LOC_362/Y INVX1_LOC_9/Y 0.09fF
C27175 INVX1_LOC_371/Y INPUT_1 0.01fF
C27176 INVX1_LOC_511/Y INVX1_LOC_335/A 0.95fF
C27177 INVX1_LOC_11/Y INVX1_LOC_145/Y 2.70fF
C27178 NAND2X1_LOC_130/Y INVX1_LOC_105/Y 0.09fF
C27179 INVX1_LOC_355/A INVX1_LOC_114/A 0.00fF
C27180 NAND2X1_LOC_111/Y INVX1_LOC_686/A 0.01fF
C27181 INVX1_LOC_378/A NAND2X1_LOC_476/a_36_24# 0.00fF
C27182 INVX1_LOC_383/A NAND2X1_LOC_274/B 0.01fF
C27183 INVX1_LOC_447/Y INVX1_LOC_50/Y 0.02fF
C27184 NAND2X1_LOC_190/A INVX1_LOC_392/A 0.00fF
C27185 INVX1_LOC_393/A INVX1_LOC_100/Y 0.08fF
C27186 INVX1_LOC_395/A INVX1_LOC_62/Y 0.25fF
C27187 INVX1_LOC_508/Y INVX1_LOC_58/Y 0.00fF
C27188 INVX1_LOC_578/A INVX1_LOC_41/Y 0.09fF
C27189 INVX1_LOC_206/Y INVX1_LOC_528/Y 0.03fF
C27190 INVX1_LOC_312/Y INVX1_LOC_646/Y 0.11fF
C27191 INVX1_LOC_162/Y INVX1_LOC_62/Y 0.01fF
C27192 NAND2X1_LOC_602/A INVX1_LOC_50/Y 0.09fF
C27193 INVX1_LOC_683/Y INVX1_LOC_9/Y 0.01fF
C27194 NAND2X1_LOC_708/A INVX1_LOC_186/Y 0.03fF
C27195 NAND2X1_LOC_136/Y INVX1_LOC_242/A 0.03fF
C27196 INVX1_LOC_362/Y INVX1_LOC_62/Y 0.07fF
C27197 INVX1_LOC_395/A INVX1_LOC_529/Y 0.04fF
C27198 INVX1_LOC_54/Y INVX1_LOC_50/Y 1.12fF
C27199 INVX1_LOC_513/Y INVX1_LOC_358/Y 0.02fF
C27200 NAND2X1_LOC_190/A INVX1_LOC_93/Y 0.01fF
C27201 INVX1_LOC_400/Y INVX1_LOC_666/Y 0.12fF
C27202 INVX1_LOC_335/Y INVX1_LOC_513/Y 0.02fF
C27203 INVX1_LOC_670/A INVX1_LOC_665/Y 0.09fF
C27204 INVX1_LOC_344/A INVX1_LOC_675/A 0.05fF
C27205 INVX1_LOC_396/Y INVX1_LOC_531/Y 0.17fF
C27206 NAND2X1_LOC_698/Y INVX1_LOC_99/Y 0.01fF
C27207 INVX1_LOC_492/A INVX1_LOC_555/A 0.02fF
C27208 INVX1_LOC_12/Y INVX1_LOC_179/A 0.08fF
C27209 INVX1_LOC_587/Y INVX1_LOC_31/Y 0.03fF
C27210 INVX1_LOC_362/Y NAND2X1_LOC_844/A 0.03fF
C27211 INVX1_LOC_17/Y NAND2X1_LOC_52/Y -0.06fF
C27212 NAND2X1_LOC_79/B INVX1_LOC_274/Y 0.03fF
C27213 INVX1_LOC_526/A INVX1_LOC_74/Y 0.13fF
C27214 INVX1_LOC_89/Y INPUT_1 0.21fF
C27215 INVX1_LOC_297/A NAND2X1_LOC_269/B 0.02fF
C27216 INVX1_LOC_674/A INVX1_LOC_157/Y 0.02fF
C27217 INVX1_LOC_254/Y INVX1_LOC_69/Y 0.15fF
C27218 INVX1_LOC_35/Y INVX1_LOC_507/Y 0.09fF
C27219 INVX1_LOC_662/A INVX1_LOC_99/Y -0.00fF
C27220 INVX1_LOC_257/A INVX1_LOC_50/Y 0.01fF
C27221 INVX1_LOC_53/Y INVX1_LOC_475/Y 0.01fF
C27222 INVX1_LOC_573/Y INVX1_LOC_522/A 0.01fF
C27223 INVX1_LOC_35/Y INVX1_LOC_223/Y 0.00fF
C27224 NAND2X1_LOC_319/a_36_24# INPUT_1 0.00fF
C27225 INVX1_LOC_35/Y NAND2X1_LOC_474/a_36_24# 0.01fF
C27226 INVX1_LOC_89/Y INVX1_LOC_292/Y 0.02fF
C27227 INVX1_LOC_197/A INVX1_LOC_74/Y 0.00fF
C27228 INVX1_LOC_521/A INVX1_LOC_50/Y 0.01fF
C27229 NAND2X1_LOC_274/B INVX1_LOC_509/A 0.08fF
C27230 NAND2X1_LOC_301/B INVX1_LOC_504/Y 0.02fF
C27231 INVX1_LOC_63/Y INVX1_LOC_355/Y 0.01fF
C27232 INVX1_LOC_592/Y INVX1_LOC_69/Y 0.00fF
C27233 INVX1_LOC_89/Y NAND2X1_LOC_279/a_36_24# 0.00fF
C27234 INVX1_LOC_544/A INVX1_LOC_680/A 0.01fF
C27235 INVX1_LOC_100/Y NAND2X1_LOC_106/B 0.03fF
C27236 NAND2X1_LOC_411/Y NAND2X1_LOC_410/Y 0.09fF
C27237 INVX1_LOC_167/A INVX1_LOC_491/A 0.30fF
C27238 NAND2X1_LOC_698/Y INVX1_LOC_47/Y 0.10fF
C27239 INVX1_LOC_204/Y NAND2X1_LOC_668/Y 0.07fF
C27240 INVX1_LOC_524/Y NAND2X1_LOC_96/a_36_24# 0.01fF
C27241 INVX1_LOC_31/Y INVX1_LOC_9/Y 0.18fF
C27242 INVX1_LOC_149/Y INVX1_LOC_58/Y 0.34fF
C27243 INVX1_LOC_607/Y NAND2X1_LOC_843/B 0.04fF
C27244 INVX1_LOC_62/Y INVX1_LOC_189/Y 0.00fF
C27245 NAND2X1_LOC_184/Y INVX1_LOC_26/Y 0.34fF
C27246 INVX1_LOC_517/Y INVX1_LOC_521/A 0.06fF
C27247 INVX1_LOC_173/Y INVX1_LOC_100/Y 0.00fF
C27248 INVX1_LOC_42/Y INVX1_LOC_86/A 0.01fF
C27249 INVX1_LOC_609/Y INVX1_LOC_613/A 0.01fF
C27250 NAND2X1_LOC_814/Y INVX1_LOC_655/A 0.04fF
C27251 INVX1_LOC_31/Y INVX1_LOC_166/Y 0.03fF
C27252 INVX1_LOC_47/Y INVX1_LOC_653/A 0.13fF
C27253 NAND2X1_LOC_174/B INVX1_LOC_74/Y 0.27fF
C27254 INVX1_LOC_79/A NAND2X1_LOC_753/Y 0.07fF
C27255 INVX1_LOC_458/Y NAND2X1_LOC_591/B 0.17fF
C27256 NAND2X1_LOC_591/Y INVX1_LOC_74/Y 0.01fF
C27257 INVX1_LOC_31/Y INVX1_LOC_62/Y 0.24fF
C27258 INVX1_LOC_41/Y INVX1_LOC_93/A 0.05fF
C27259 INVX1_LOC_527/Y INVX1_LOC_91/Y 0.01fF
C27260 INVX1_LOC_31/Y NAND2X1_LOC_844/A 0.22fF
C27261 INVX1_LOC_345/A NAND2X1_LOC_832/A 0.23fF
C27262 INVX1_LOC_369/Y INVX1_LOC_328/Y 0.18fF
C27263 INVX1_LOC_69/Y INVX1_LOC_479/A 7.88fF
C27264 INVX1_LOC_653/A INVX1_LOC_119/Y 0.01fF
C27265 INVX1_LOC_435/Y INVX1_LOC_222/Y 0.08fF
C27266 INVX1_LOC_100/Y NAND2X1_LOC_395/Y 0.01fF
C27267 VDD INVX1_LOC_34/Y 0.24fF
C27268 VDD INVX1_LOC_237/Y 0.21fF
C27269 INVX1_LOC_75/Y INVX1_LOC_26/Y 3.15fF
C27270 INVX1_LOC_79/A INVX1_LOC_652/Y 0.02fF
C27271 VDD INVX1_LOC_38/A 0.00fF
C27272 INVX1_LOC_224/Y INVX1_LOC_160/Y 0.11fF
C27273 INVX1_LOC_566/A INVX1_LOC_458/Y 0.02fF
C27274 INVX1_LOC_206/Y INVX1_LOC_580/A 0.01fF
C27275 VDD NAND2X1_LOC_538/B 0.03fF
C27276 NAND2X1_LOC_475/A NAND2X1_LOC_383/Y 0.00fF
C27277 INVX1_LOC_578/A NAND2X1_LOC_735/a_36_24# 0.01fF
C27278 INPUT_6 INVX1_LOC_29/Y 0.45fF
C27279 NAND2X1_LOC_231/A NAND2X1_LOC_506/B 0.10fF
C27280 NAND2X1_LOC_523/B INVX1_LOC_217/Y 0.00fF
C27281 NAND2X1_LOC_371/a_36_24# INVX1_LOC_362/Y 0.01fF
C27282 VDD INVX1_LOC_537/Y 0.53fF
C27283 NAND2X1_LOC_231/A INVX1_LOC_45/Y 0.04fF
C27284 INVX1_LOC_21/Y INVX1_LOC_224/Y 0.10fF
C27285 NAND2X1_LOC_108/Y INVX1_LOC_651/A 0.36fF
C27286 NAND2X1_LOC_174/B NAND2X1_LOC_591/B 0.06fF
C27287 VDD INVX1_LOC_418/Y 0.21fF
C27288 INVX1_LOC_33/Y INVX1_LOC_63/A 0.02fF
C27289 VDD INVX1_LOC_159/Y 1.38fF
C27290 NAND2X1_LOC_591/Y NAND2X1_LOC_591/B 0.02fF
C27291 INVX1_LOC_84/A INVX1_LOC_666/A 0.02fF
C27292 INVX1_LOC_270/A NAND2X1_LOC_180/B 0.02fF
C27293 INVX1_LOC_438/Y INVX1_LOC_437/A 0.03fF
C27294 NAND2X1_LOC_718/a_36_24# INVX1_LOC_638/A 0.01fF
C27295 INVX1_LOC_21/Y INVX1_LOC_578/A 0.08fF
C27296 INVX1_LOC_71/Y NAND2X1_LOC_294/Y 0.01fF
C27297 INVX1_LOC_320/Y INVX1_LOC_99/Y 0.02fF
C27298 INVX1_LOC_454/A INVX1_LOC_298/A 0.03fF
C27299 INVX1_LOC_375/A INVX1_LOC_252/A 0.00fF
C27300 INVX1_LOC_438/A INVX1_LOC_54/Y 0.10fF
C27301 INVX1_LOC_446/Y INVX1_LOC_367/Y 0.07fF
C27302 INVX1_LOC_558/A NAND2X1_LOC_411/Y 0.05fF
C27303 INVX1_LOC_80/A NAND2X1_LOC_332/B 0.66fF
C27304 INVX1_LOC_191/Y INVX1_LOC_543/Y 0.16fF
C27305 INVX1_LOC_555/Y INVX1_LOC_136/Y 0.00fF
C27306 NAND2X1_LOC_332/B NAND2X1_LOC_768/A 0.00fF
C27307 INVX1_LOC_17/Y INVX1_LOC_65/Y 0.40fF
C27308 INVX1_LOC_24/A INVX1_LOC_54/Y 0.00fF
C27309 VDD INVX1_LOC_340/A 0.09fF
C27310 INVX1_LOC_224/Y NAND2X1_LOC_267/A 0.30fF
C27311 INPUT_0 INVX1_LOC_361/Y 0.07fF
C27312 VDD INVX1_LOC_212/Y 0.48fF
C27313 INVX1_LOC_80/A INVX1_LOC_125/Y 0.06fF
C27314 NAND2X1_LOC_574/a_36_24# INVX1_LOC_510/A 0.01fF
C27315 NAND2X1_LOC_698/a_36_24# INVX1_LOC_600/A 0.01fF
C27316 NAND2X1_LOC_106/Y INVX1_LOC_118/Y 0.01fF
C27317 NAND2X1_LOC_516/Y INVX1_LOC_361/Y 0.07fF
C27318 INVX1_LOC_384/A INVX1_LOC_367/Y 0.07fF
C27319 INVX1_LOC_553/Y INVX1_LOC_6/Y 0.00fF
C27320 NAND2X1_LOC_130/Y INVX1_LOC_126/Y 0.02fF
C27321 NAND2X1_LOC_45/Y NAND2X1_LOC_178/a_36_24# 0.00fF
C27322 NAND2X1_LOC_190/A INVX1_LOC_362/Y 0.05fF
C27323 INVX1_LOC_395/A INVX1_LOC_87/A 0.07fF
C27324 NAND2X1_LOC_338/a_36_24# NAND2X1_LOC_755/B 0.00fF
C27325 INVX1_LOC_160/Y INVX1_LOC_227/Y 0.04fF
C27326 INVX1_LOC_11/Y NAND2X1_LOC_332/B 0.07fF
C27327 VDD INVX1_LOC_569/Y 0.21fF
C27328 INPUT_0 INVX1_LOC_261/Y 0.12fF
C27329 NAND2X1_LOC_172/a_36_24# INVX1_LOC_288/A 0.00fF
C27330 NAND2X1_LOC_13/Y INVX1_LOC_194/A 0.00fF
C27331 INVX1_LOC_410/Y INVX1_LOC_6/Y 0.08fF
C27332 INVX1_LOC_254/Y INVX1_LOC_586/A 0.26fF
C27333 INVX1_LOC_566/Y INVX1_LOC_145/Y 0.22fF
C27334 INVX1_LOC_179/Y INVX1_LOC_181/A 0.00fF
C27335 INVX1_LOC_206/Y INVX1_LOC_411/Y 0.05fF
C27336 INVX1_LOC_374/A INVX1_LOC_355/Y 0.01fF
C27337 INVX1_LOC_55/A INVX1_LOC_55/Y 0.01fF
C27338 INVX1_LOC_358/A INVX1_LOC_358/Y 0.01fF
C27339 INVX1_LOC_522/Y INVX1_LOC_35/Y 0.13fF
C27340 INVX1_LOC_79/A INVX1_LOC_458/Y 0.10fF
C27341 NAND2X1_LOC_576/a_36_24# INVX1_LOC_433/A 0.00fF
C27342 INVX1_LOC_413/Y INVX1_LOC_387/Y 0.01fF
C27343 NAND2X1_LOC_46/a_36_24# INVX1_LOC_255/A 0.00fF
C27344 INVX1_LOC_84/A NAND2X1_LOC_673/A 0.01fF
C27345 NAND2X1_LOC_728/B NAND2X1_LOC_728/A 0.08fF
C27346 INVX1_LOC_442/A INVX1_LOC_66/A 0.01fF
C27347 NAND2X1_LOC_174/B INVX1_LOC_566/A 0.00fF
C27348 INVX1_LOC_613/Y INVX1_LOC_626/A 0.19fF
C27349 VDD INVX1_LOC_405/Y 0.28fF
C27350 INVX1_LOC_381/A INVX1_LOC_280/Y 0.00fF
C27351 INVX1_LOC_626/A NAND2X1_LOC_612/A 0.14fF
C27352 INVX1_LOC_592/Y INVX1_LOC_586/A 0.02fF
C27353 INVX1_LOC_21/Y INVX1_LOC_468/Y 0.03fF
C27354 INVX1_LOC_566/A INVX1_LOC_260/Y 0.01fF
C27355 INVX1_LOC_678/Y INVX1_LOC_641/Y 0.01fF
C27356 NAND2X1_LOC_573/a_36_24# INVX1_LOC_502/A 0.01fF
C27357 NAND2X1_LOC_150/a_36_24# INVX1_LOC_255/A 0.00fF
C27358 INVX1_LOC_68/Y INVX1_LOC_199/Y 0.03fF
C27359 VDD INVX1_LOC_468/A -0.00fF
C27360 INVX1_LOC_377/A INVX1_LOC_371/A 0.20fF
C27361 NAND2X1_LOC_795/a_36_24# INVX1_LOC_274/A 0.00fF
C27362 INVX1_LOC_267/Y NAND2X1_LOC_720/A 0.11fF
C27363 INVX1_LOC_580/A NAND2X1_LOC_334/A 0.08fF
C27364 INVX1_LOC_426/Y INVX1_LOC_75/Y 0.06fF
C27365 NAND2X1_LOC_780/A INVX1_LOC_6/Y 0.15fF
C27366 INVX1_LOC_367/Y INVX1_LOC_145/Y 0.08fF
C27367 NAND2X1_LOC_650/a_36_24# INVX1_LOC_498/A 0.01fF
C27368 INVX1_LOC_54/Y NAND2X1_LOC_513/A 0.01fF
C27369 INVX1_LOC_406/Y INVX1_LOC_6/Y 0.04fF
C27370 INVX1_LOC_469/Y INVX1_LOC_197/A 0.03fF
C27371 INVX1_LOC_672/Y INVX1_LOC_661/Y 0.01fF
C27372 INVX1_LOC_371/Y INVX1_LOC_50/Y 0.21fF
C27373 VDD INVX1_LOC_450/Y 0.21fF
C27374 INVX1_LOC_324/Y INVX1_LOC_46/Y 0.01fF
C27375 INVX1_LOC_206/Y INVX1_LOC_41/Y 0.26fF
C27376 INVX1_LOC_51/Y INVX1_LOC_9/Y 0.08fF
C27377 VDD INVX1_LOC_39/Y 0.26fF
C27378 INVX1_LOC_632/A INVX1_LOC_686/Y 0.03fF
C27379 INVX1_LOC_17/Y INVX1_LOC_479/Y 0.02fF
C27380 INVX1_LOC_612/Y INVX1_LOC_610/A 0.01fF
C27381 NAND2X1_LOC_522/a_36_24# INVX1_LOC_6/Y 0.00fF
C27382 INVX1_LOC_420/Y INVX1_LOC_280/A 0.01fF
C27383 INVX1_LOC_80/A NAND2X1_LOC_128/B 0.07fF
C27384 INVX1_LOC_545/Y INVX1_LOC_253/Y 0.26fF
C27385 INVX1_LOC_31/Y INVX1_LOC_344/A 0.05fF
C27386 INVX1_LOC_134/Y NAND2X1_LOC_606/a_36_24# 0.01fF
C27387 INVX1_LOC_153/Y INVX1_LOC_94/A 0.02fF
C27388 INVX1_LOC_686/A INVX1_LOC_411/Y 0.00fF
C27389 INVX1_LOC_581/A NAND2X1_LOC_612/a_36_24# 0.00fF
C27390 INVX1_LOC_53/Y NAND2X1_LOC_611/a_36_24# 0.00fF
C27391 INVX1_LOC_335/Y INVX1_LOC_93/A 0.03fF
C27392 NAND2X1_LOC_330/a_36_24# INVX1_LOC_74/Y 0.01fF
C27393 INVX1_LOC_17/Y INVX1_LOC_318/A 0.02fF
C27394 NAND2X1_LOC_97/A INVX1_LOC_90/Y 0.03fF
C27395 INVX1_LOC_560/A INVX1_LOC_75/Y 0.07fF
C27396 INVX1_LOC_437/Y INVX1_LOC_444/A 0.14fF
C27397 INVX1_LOC_561/A INVX1_LOC_99/Y 0.08fF
C27398 INVX1_LOC_397/A INVX1_LOC_531/Y 0.06fF
C27399 INVX1_LOC_12/Y INVX1_LOC_69/Y 0.18fF
C27400 NAND2X1_LOC_307/A INVX1_LOC_63/Y 0.04fF
C27401 INVX1_LOC_266/A INVX1_LOC_9/Y 0.03fF
C27402 INVX1_LOC_545/Y INVX1_LOC_63/Y 0.02fF
C27403 VDD INVX1_LOC_620/Y 0.35fF
C27404 INVX1_LOC_257/Y INVX1_LOC_625/Y 0.01fF
C27405 INVX1_LOC_531/Y INVX1_LOC_94/A 0.02fF
C27406 INVX1_LOC_199/Y INVX1_LOC_600/A 0.17fF
C27407 INVX1_LOC_301/Y INVX1_LOC_686/A 0.11fF
C27408 INVX1_LOC_544/A INVX1_LOC_66/A 0.01fF
C27409 INVX1_LOC_258/Y NAND2X1_LOC_123/A 0.03fF
C27410 INVX1_LOC_116/Y INVX1_LOC_66/A 0.05fF
C27411 INVX1_LOC_322/Y INVX1_LOC_11/A 0.00fF
C27412 INVX1_LOC_93/Y INVX1_LOC_480/Y 0.01fF
C27413 INVX1_LOC_51/Y INVX1_LOC_62/Y 0.10fF
C27414 NAND2X1_LOC_498/Y INVX1_LOC_666/Y 0.01fF
C27415 INVX1_LOC_59/Y NAND2X1_LOC_753/Y 0.01fF
C27416 INVX1_LOC_586/A NAND2X1_LOC_528/Y 0.02fF
C27417 NAND2X1_LOC_176/Y INVX1_LOC_92/A 0.03fF
C27418 NAND2X1_LOC_39/Y INVX1_LOC_90/Y 0.01fF
C27419 INVX1_LOC_227/Y NAND2X1_LOC_267/A 0.23fF
C27420 INVX1_LOC_80/A INVX1_LOC_242/Y 0.18fF
C27421 NAND2X1_LOC_591/Y INVX1_LOC_469/Y 0.01fF
C27422 INVX1_LOC_134/A NAND2X1_LOC_544/B 0.00fF
C27423 NAND2X1_LOC_775/B NAND2X1_LOC_443/a_36_24# 0.01fF
C27424 INVX1_LOC_419/Y INVX1_LOC_253/Y 0.01fF
C27425 INVX1_LOC_586/A INVX1_LOC_479/A 1.52fF
C27426 INVX1_LOC_336/Y INVX1_LOC_100/Y 0.01fF
C27427 INVX1_LOC_35/Y INVX1_LOC_508/A 0.65fF
C27428 INVX1_LOC_266/A INVX1_LOC_62/Y 0.03fF
C27429 INVX1_LOC_197/A INVX1_LOC_79/A 0.03fF
C27430 INVX1_LOC_89/Y INVX1_LOC_50/Y 0.22fF
C27431 INVX1_LOC_442/Y INVX1_LOC_682/A 0.01fF
C27432 INVX1_LOC_93/Y INVX1_LOC_169/Y 0.14fF
C27433 INVX1_LOC_674/A INVX1_LOC_6/Y 0.02fF
C27434 INVX1_LOC_54/Y NAND2X1_LOC_388/A 1.04fF
C27435 INVX1_LOC_155/Y INVX1_LOC_245/A 0.01fF
C27436 INVX1_LOC_686/A INVX1_LOC_41/Y 0.18fF
C27437 INVX1_LOC_261/Y INVX1_LOC_498/A 0.71fF
C27438 INVX1_LOC_312/Y NAND2X1_LOC_528/Y 0.01fF
C27439 NAND2X1_LOC_267/a_36_24# INVX1_LOC_9/Y 0.00fF
C27440 INVX1_LOC_166/A NAND2X1_LOC_542/A 0.07fF
C27441 INVX1_LOC_377/Y INVX1_LOC_666/Y 0.17fF
C27442 INVX1_LOC_89/Y INVX1_LOC_431/Y 0.06fF
C27443 NAND2X1_LOC_121/Y INVX1_LOC_259/Y 0.01fF
C27444 NAND2X1_LOC_521/Y INVX1_LOC_69/Y 0.07fF
C27445 INVX1_LOC_312/Y INVX1_LOC_479/A 0.03fF
C27446 NAND2X1_LOC_333/A INVX1_LOC_69/Y 0.74fF
C27447 INVX1_LOC_17/Y INVX1_LOC_244/Y 0.16fF
C27448 INVX1_LOC_391/A INVX1_LOC_69/Y 0.01fF
C27449 INVX1_LOC_501/A INVX1_LOC_50/Y 0.03fF
C27450 NAND2X1_LOC_179/Y INVX1_LOC_100/Y 0.01fF
C27451 INVX1_LOC_347/Y INVX1_LOC_359/Y 0.02fF
C27452 INVX1_LOC_31/Y INVX1_LOC_624/Y 0.00fF
C27453 INVX1_LOC_179/A NAND2X1_LOC_615/B 0.01fF
C27454 INVX1_LOC_11/Y INVX1_LOC_242/Y 0.07fF
C27455 INVX1_LOC_536/A INVX1_LOC_495/Y 0.23fF
C27456 NAND2X1_LOC_416/Y NAND2X1_LOC_631/B 0.01fF
C27457 INVX1_LOC_41/Y INVX1_LOC_14/A 0.01fF
C27458 NAND2X1_LOC_111/Y NAND2X1_LOC_542/A 0.40fF
C27459 INVX1_LOC_105/A NAND2X1_LOC_274/B 0.17fF
C27460 INVX1_LOC_117/Y INVX1_LOC_124/A 0.08fF
C27461 NAND2X1_LOC_270/a_36_24# INVX1_LOC_280/A 0.00fF
C27462 INVX1_LOC_99/Y INVX1_LOC_653/Y 0.00fF
C27463 INVX1_LOC_44/Y INVX1_LOC_292/Y 0.11fF
C27464 INVX1_LOC_145/Y NAND2X1_LOC_843/B 0.08fF
C27465 INVX1_LOC_58/Y INVX1_LOC_493/Y 0.01fF
C27466 INVX1_LOC_11/Y INVX1_LOC_487/A 0.01fF
C27467 INVX1_LOC_99/Y INVX1_LOC_666/Y 0.17fF
C27468 INVX1_LOC_44/Y INVX1_LOC_284/Y 0.04fF
C27469 INVX1_LOC_496/A INVX1_LOC_168/Y 0.02fF
C27470 INVX1_LOC_376/A INVX1_LOC_63/Y 0.18fF
C27471 INVX1_LOC_330/A INVX1_LOC_479/A 0.15fF
C27472 INVX1_LOC_74/Y INVX1_LOC_440/Y 0.22fF
C27473 NAND2X1_LOC_128/A INVX1_LOC_100/Y 0.19fF
C27474 NAND2X1_LOC_451/B INVX1_LOC_505/A 0.12fF
C27475 NAND2X1_LOC_591/Y INVX1_LOC_460/A 0.00fF
C27476 NAND2X1_LOC_133/a_36_24# INVX1_LOC_319/A 0.00fF
C27477 NAND2X1_LOC_231/B INVX1_LOC_197/Y 0.46fF
C27478 INPUT_1 INVX1_LOC_347/A 0.07fF
C27479 NAND2X1_LOC_555/B NAND2X1_LOC_481/a_36_24# 0.02fF
C27480 INVX1_LOC_399/A INVX1_LOC_44/Y 0.06fF
C27481 NAND2X1_LOC_136/Y NAND2X1_LOC_542/A 0.02fF
C27482 NAND2X1_LOC_127/a_36_24# INVX1_LOC_100/Y 0.01fF
C27483 NAND2X1_LOC_449/B INVX1_LOC_114/A 0.09fF
C27484 INVX1_LOC_434/A INVX1_LOC_220/A 0.15fF
C27485 INVX1_LOC_211/A NAND2X1_LOC_333/B 0.01fF
C27486 INVX1_LOC_63/Y INVX1_LOC_502/A 0.68fF
C27487 NAND2X1_LOC_275/Y NAND2X1_LOC_271/A 0.09fF
C27488 INVX1_LOC_47/Y INVX1_LOC_653/Y 0.02fF
C27489 NAND2X1_LOC_334/A INVX1_LOC_41/Y 0.12fF
C27490 NAND2X1_LOC_301/B INVX1_LOC_114/A 0.06fF
C27491 NAND2X1_LOC_528/Y INVX1_LOC_225/Y 0.04fF
C27492 NAND2X1_LOC_370/A NAND2X1_LOC_76/B 0.02fF
C27493 NAND2X1_LOC_249/Y INVX1_LOC_607/A 0.02fF
C27494 NAND2X1_LOC_66/Y NAND2X1_LOC_625/a_36_24# 0.00fF
C27495 INVX1_LOC_320/Y NAND2X1_LOC_475/A 0.01fF
C27496 INVX1_LOC_119/Y INVX1_LOC_653/Y 0.00fF
C27497 NAND2X1_LOC_88/Y INVX1_LOC_65/Y 0.29fF
C27498 INVX1_LOC_100/Y NAND2X1_LOC_248/B 0.04fF
C27499 VDD NAND2X1_LOC_163/B 0.03fF
C27500 INVX1_LOC_119/Y INVX1_LOC_666/Y 0.07fF
C27501 INVX1_LOC_41/Y NAND2X1_LOC_609/B 0.00fF
C27502 INVX1_LOC_548/Y INVX1_LOC_556/A 0.13fF
C27503 NAND2X1_LOC_331/A INVX1_LOC_162/Y 0.01fF
C27504 VDD INVX1_LOC_172/Y 0.21fF
C27505 INVX1_LOC_206/Y INVX1_LOC_315/Y 0.07fF
C27506 INVX1_LOC_74/Y INVX1_LOC_66/Y 0.01fF
C27507 INVX1_LOC_647/Y INVX1_LOC_669/A 0.03fF
C27508 NAND2X1_LOC_781/B INVX1_LOC_53/Y 0.37fF
C27509 NAND2X1_LOC_541/a_36_24# INVX1_LOC_384/A 0.01fF
C27510 INVX1_LOC_19/Y INVX1_LOC_55/Y 0.01fF
C27511 INVX1_LOC_21/Y NAND2X1_LOC_86/Y 0.11fF
C27512 INVX1_LOC_301/A INVX1_LOC_80/A 0.01fF
C27513 INVX1_LOC_393/Y INVX1_LOC_384/A -0.03fF
C27514 NAND2X1_LOC_180/a_36_24# INVX1_LOC_270/A 0.01fF
C27515 NAND2X1_LOC_152/B INVX1_LOC_554/Y 0.18fF
C27516 VDD INVX1_LOC_377/A 0.00fF
C27517 VDD NAND2X1_LOC_595/Y 0.06fF
C27518 NAND2X1_LOC_7/Y INVX1_LOC_11/Y 0.02fF
C27519 INVX1_LOC_420/Y INVX1_LOC_449/A 0.00fF
C27520 NAND2X1_LOC_558/a_36_24# INVX1_LOC_320/A 0.01fF
C27521 INVX1_LOC_335/Y INVX1_LOC_206/Y 0.10fF
C27522 INVX1_LOC_279/Y INVX1_LOC_439/Y 0.04fF
C27523 NAND2X1_LOC_503/a_36_24# INVX1_LOC_273/A 0.01fF
C27524 INVX1_LOC_21/Y INVX1_LOC_206/Y 0.36fF
C27525 VDD INVX1_LOC_57/Y 0.05fF
C27526 VDD INVX1_LOC_455/A 0.16fF
C27527 NAND2X1_LOC_231/A NAND2X1_LOC_756/Y 0.03fF
C27528 VDD INVX1_LOC_352/Y 0.37fF
C27529 INVX1_LOC_93/Y INVX1_LOC_638/A 0.03fF
C27530 NAND2X1_LOC_503/B INVX1_LOC_208/Y 0.11fF
C27531 INPUT_0 INVX1_LOC_442/Y 0.02fF
C27532 INVX1_LOC_463/A INVX1_LOC_539/Y 0.04fF
C27533 NAND2X1_LOC_317/B INVX1_LOC_251/A 0.20fF
C27534 INVX1_LOC_320/A INVX1_LOC_321/A 0.02fF
C27535 INVX1_LOC_393/Y INVX1_LOC_145/Y 0.04fF
C27536 INVX1_LOC_575/A INVX1_LOC_395/A 0.02fF
C27537 NAND2X1_LOC_331/A INVX1_LOC_189/Y 0.01fF
C27538 INVX1_LOC_106/A NAND2X1_LOC_142/Y 0.00fF
C27539 INVX1_LOC_12/Y INVX1_LOC_586/A 0.24fF
C27540 NAND2X1_LOC_241/B INVX1_LOC_209/A 0.01fF
C27541 INVX1_LOC_683/A INVX1_LOC_45/Y 0.03fF
C27542 INVX1_LOC_366/Y INVX1_LOC_72/Y 0.93fF
C27543 INVX1_LOC_206/Y NAND2X1_LOC_267/A 0.09fF
C27544 INVX1_LOC_20/Y INVX1_LOC_80/A 1.27fF
C27545 INVX1_LOC_372/Y NAND2X1_LOC_440/a_36_24# 0.00fF
C27546 INVX1_LOC_551/Y NAND2X1_LOC_601/a_36_24# 0.06fF
C27547 INVX1_LOC_526/A INVX1_LOC_632/A 0.02fF
C27548 INVX1_LOC_442/A INVX1_LOC_116/Y 1.38fF
C27549 INVX1_LOC_118/Y INPUT_1 0.03fF
C27550 INVX1_LOC_168/A INVX1_LOC_633/Y 0.01fF
C27551 INVX1_LOC_166/A INVX1_LOC_121/Y 0.04fF
C27552 INVX1_LOC_675/A INVX1_LOC_638/A 0.00fF
C27553 INVX1_LOC_21/Y INVX1_LOC_396/Y 0.42fF
C27554 INVX1_LOC_173/A INVX1_LOC_35/Y 0.01fF
C27555 INVX1_LOC_76/Y INVX1_LOC_154/Y 0.04fF
C27556 INVX1_LOC_193/Y INVX1_LOC_117/Y 0.02fF
C27557 INVX1_LOC_625/A INVX1_LOC_273/A 0.02fF
C27558 INVX1_LOC_596/A INVX1_LOC_519/A 0.03fF
C27559 INVX1_LOC_142/Y INVX1_LOC_145/Y 0.02fF
C27560 INVX1_LOC_206/Y INVX1_LOC_555/A 0.01fF
C27561 INVX1_LOC_312/Y INVX1_LOC_12/Y 0.06fF
C27562 INVX1_LOC_335/Y INVX1_LOC_686/A 0.07fF
C27563 INVX1_LOC_278/A NAND2X1_LOC_252/Y 0.05fF
C27564 INVX1_LOC_582/A NAND2X1_LOC_739/a_36_24# 0.02fF
C27565 INVX1_LOC_392/Y INVX1_LOC_665/Y 0.01fF
C27566 INVX1_LOC_21/Y INVX1_LOC_686/A 0.07fF
C27567 INVX1_LOC_582/Y INVX1_LOC_137/Y 0.01fF
C27568 INVX1_LOC_166/A INVX1_LOC_253/A 0.02fF
C27569 INVX1_LOC_446/A INVX1_LOC_502/A 0.66fF
C27570 NAND2X1_LOC_513/A NAND2X1_LOC_677/Y 0.20fF
C27571 INVX1_LOC_20/Y INVX1_LOC_11/Y 0.21fF
C27572 INVX1_LOC_21/Y INVX1_LOC_80/Y 0.01fF
C27573 INVX1_LOC_604/A INVX1_LOC_69/Y 0.01fF
C27574 INVX1_LOC_45/Y INVX1_LOC_463/Y 0.04fF
C27575 INVX1_LOC_441/Y INVX1_LOC_89/Y 0.03fF
C27576 INVX1_LOC_300/A INVX1_LOC_80/A 0.07fF
C27577 NAND2X1_LOC_142/Y INVX1_LOC_239/A 0.17fF
C27578 INVX1_LOC_361/Y INVX1_LOC_384/A 0.34fF
C27579 INVX1_LOC_208/Y INVX1_LOC_273/A 0.03fF
C27580 NAND2X1_LOC_194/a_36_24# INVX1_LOC_31/Y 0.01fF
C27581 NAND2X1_LOC_16/Y INVX1_LOC_47/Y 0.04fF
C27582 NAND2X1_LOC_521/Y INVX1_LOC_586/A 0.07fF
C27583 INVX1_LOC_434/Y INVX1_LOC_17/Y 0.01fF
C27584 NAND2X1_LOC_387/Y NAND2X1_LOC_318/A 0.89fF
C27585 INVX1_LOC_97/Y INVX1_LOC_99/Y 0.04fF
C27586 INPUT_0 INVX1_LOC_482/Y 0.00fF
C27587 INVX1_LOC_11/Y NAND2X1_LOC_473/a_36_24# 0.00fF
C27588 INVX1_LOC_80/A INVX1_LOC_197/Y 0.03fF
C27589 NAND2X1_LOC_651/a_36_24# INVX1_LOC_463/Y 0.01fF
C27590 INVX1_LOC_433/Y INVX1_LOC_244/Y 0.04fF
C27591 INVX1_LOC_442/A INVX1_LOC_255/A 0.43fF
C27592 NAND2X1_LOC_169/A INVX1_LOC_160/A 0.02fF
C27593 INVX1_LOC_224/Y INVX1_LOC_26/Y 0.08fF
C27594 INVX1_LOC_129/A INVX1_LOC_99/A 0.01fF
C27595 INVX1_LOC_463/A INVX1_LOC_62/Y 0.07fF
C27596 INVX1_LOC_288/A INVX1_LOC_258/Y 0.01fF
C27597 INPUT_0 INVX1_LOC_471/Y 0.01fF
C27598 INVX1_LOC_374/A INVX1_LOC_376/A 0.21fF
C27599 INVX1_LOC_146/A INVX1_LOC_66/A 0.00fF
C27600 VDD INVX1_LOC_203/A -0.00fF
C27601 INVX1_LOC_9/Y INVX1_LOC_216/Y 0.00fF
C27602 INVX1_LOC_406/Y NAND2X1_LOC_294/Y 3.29fF
C27603 VDD INVX1_LOC_280/A 0.05fF
C27604 NAND2X1_LOC_174/B INVX1_LOC_632/A 0.07fF
C27605 INVX1_LOC_605/Y INVX1_LOC_46/Y 0.01fF
C27606 INVX1_LOC_391/Y INVX1_LOC_99/Y 0.56fF
C27607 INVX1_LOC_127/A INVX1_LOC_519/Y 0.20fF
C27608 VDD NAND2X1_LOC_372/Y 0.04fF
C27609 NAND2X1_LOC_228/a_36_24# INVX1_LOC_211/A 0.00fF
C27610 NAND2X1_LOC_24/Y INVX1_LOC_46/Y 0.06fF
C27611 INVX1_LOC_193/A NAND2X1_LOC_325/B 0.20fF
C27612 INVX1_LOC_578/A INVX1_LOC_26/Y 0.65fF
C27613 INVX1_LOC_11/Y INVX1_LOC_300/A 0.10fF
C27614 INVX1_LOC_106/Y INVX1_LOC_107/A 0.15fF
C27615 NAND2X1_LOC_791/B INVX1_LOC_592/Y 0.01fF
C27616 INVX1_LOC_456/Y INVX1_LOC_455/A 0.00fF
C27617 INVX1_LOC_448/A INVX1_LOC_361/Y 0.18fF
C27618 INVX1_LOC_167/Y INVX1_LOC_496/A 0.02fF
C27619 NAND2X1_LOC_173/Y INVX1_LOC_347/Y 0.01fF
C27620 NAND2X1_LOC_591/Y INVX1_LOC_632/A 0.25fF
C27621 INVX1_LOC_431/A INVX1_LOC_99/Y 0.01fF
C27622 NAND2X1_LOC_416/Y INVX1_LOC_48/Y 0.03fF
C27623 INVX1_LOC_578/Y NAND2X1_LOC_123/A 0.13fF
C27624 INPUT_1 NAND2X1_LOC_418/Y 0.12fF
C27625 NAND2X1_LOC_775/B INVX1_LOC_35/Y 0.01fF
C27626 INVX1_LOC_288/A NAND2X1_LOC_431/a_36_24# 0.00fF
C27627 INVX1_LOC_175/A INVX1_LOC_63/Y 0.24fF
C27628 INVX1_LOC_202/Y INVX1_LOC_478/Y 0.01fF
C27629 INVX1_LOC_45/Y NAND2X1_LOC_274/B 0.03fF
C27630 INVX1_LOC_238/Y INVX1_LOC_241/A 0.03fF
C27631 INVX1_LOC_662/A INVX1_LOC_131/Y 0.03fF
C27632 NAND2X1_LOC_775/B INVX1_LOC_304/A 0.00fF
C27633 INVX1_LOC_412/Y INVX1_LOC_74/Y 0.09fF
C27634 INVX1_LOC_589/Y INVX1_LOC_97/Y 0.02fF
C27635 NAND2X1_LOC_475/A INVX1_LOC_666/Y 0.03fF
C27636 INVX1_LOC_652/A NAND2X1_LOC_831/a_36_24# 0.00fF
C27637 INVX1_LOC_447/Y INVX1_LOC_117/Y 0.12fF
C27638 INVX1_LOC_392/A INVX1_LOC_665/Y 0.00fF
C27639 NAND2X1_LOC_56/Y INVX1_LOC_199/Y 0.08fF
C27640 NAND2X1_LOC_13/Y INVX1_LOC_9/Y 0.08fF
C27641 NAND2X1_LOC_697/Y INVX1_LOC_93/Y 0.01fF
C27642 INVX1_LOC_183/A INVX1_LOC_12/A 0.01fF
C27643 INVX1_LOC_397/A INVX1_LOC_41/Y 0.07fF
C27644 INVX1_LOC_49/Y INVX1_LOC_188/Y 0.03fF
C27645 INVX1_LOC_70/Y INVX1_LOC_6/Y 0.01fF
C27646 INVX1_LOC_381/Y INVX1_LOC_382/Y 0.05fF
C27647 NAND2X1_LOC_111/Y NAND2X1_LOC_323/a_36_24# 0.00fF
C27648 INVX1_LOC_41/Y INVX1_LOC_94/A 0.01fF
C27649 INVX1_LOC_261/Y INVX1_LOC_145/Y 0.03fF
C27650 INVX1_LOC_188/Y INVX1_LOC_533/A 0.03fF
C27651 NAND2X1_LOC_252/Y INVX1_LOC_453/Y 0.50fF
C27652 INVX1_LOC_93/Y INVX1_LOC_665/Y 0.01fF
C27653 INVX1_LOC_54/Y INVX1_LOC_117/Y 0.18fF
C27654 INVX1_LOC_94/Y INVX1_LOC_99/Y 0.03fF
C27655 INVX1_LOC_20/Y INVX1_LOC_102/Y 0.01fF
C27656 INVX1_LOC_617/Y INVX1_LOC_100/Y 0.12fF
C27657 INVX1_LOC_119/A INVX1_LOC_100/Y 0.01fF
C27658 INVX1_LOC_27/A INVX1_LOC_9/Y 0.01fF
C27659 INVX1_LOC_381/A NAND2X1_LOC_268/a_36_24# 0.00fF
C27660 INVX1_LOC_48/Y INVX1_LOC_260/Y 0.10fF
C27661 INVX1_LOC_255/A INVX1_LOC_116/Y 0.05fF
C27662 INVX1_LOC_176/Y INVX1_LOC_100/Y 0.06fF
C27663 NAND2X1_LOC_399/B INVX1_LOC_183/A 0.03fF
C27664 INVX1_LOC_608/Y INVX1_LOC_63/Y 0.00fF
C27665 INVX1_LOC_18/A INPUT_4 0.01fF
C27666 INVX1_LOC_623/Y INVX1_LOC_601/Y 0.32fF
C27667 INVX1_LOC_83/A INVX1_LOC_83/Y 0.01fF
C27668 NAND2X1_LOC_491/a_36_24# INVX1_LOC_75/Y 0.01fF
C27669 INVX1_LOC_69/Y INVX1_LOC_159/A 0.00fF
C27670 INVX1_LOC_17/Y INVX1_LOC_63/Y 0.15fF
C27671 NAND2X1_LOC_13/Y INVX1_LOC_62/Y 0.03fF
C27672 INVX1_LOC_80/A INVX1_LOC_655/A 0.16fF
C27673 INVX1_LOC_537/A INVX1_LOC_357/Y 0.03fF
C27674 INVX1_LOC_183/A INVX1_LOC_7/Y 0.11fF
C27675 INVX1_LOC_452/A NAND2X1_LOC_480/a_36_24# 0.00fF
C27676 INVX1_LOC_137/Y INVX1_LOC_496/A 0.07fF
C27677 INVX1_LOC_431/A NAND2X1_LOC_557/B 0.05fF
C27678 INVX1_LOC_31/Y INVX1_LOC_169/Y 0.01fF
C27679 INVX1_LOC_267/Y INVX1_LOC_79/A 0.13fF
C27680 NAND2X1_LOC_97/B INVX1_LOC_79/A 0.02fF
C27681 INVX1_LOC_69/Y NAND2X1_LOC_615/B 0.03fF
C27682 INVX1_LOC_68/Y NAND2X1_LOC_230/a_36_24# 0.00fF
C27683 NAND2X1_LOC_451/B NAND2X1_LOC_430/a_36_24# 0.02fF
C27684 INVX1_LOC_417/A INVX1_LOC_79/A 0.01fF
C27685 NAND2X1_LOC_528/Y INVX1_LOC_486/Y 0.02fF
C27686 INVX1_LOC_283/Y INVX1_LOC_671/A 0.00fF
C27687 NAND2X1_LOC_333/A INVX1_LOC_157/Y 0.11fF
C27688 NAND2X1_LOC_387/Y INVX1_LOC_49/Y 0.02fF
C27689 INVX1_LOC_166/A NAND2X1_LOC_498/a_36_24# 0.00fF
C27690 INVX1_LOC_44/Y INVX1_LOC_50/Y 0.16fF
C27691 INVX1_LOC_99/Y NAND2X1_LOC_489/A 0.01fF
C27692 INVX1_LOC_99/Y NAND2X1_LOC_806/a_36_24# 0.00fF
C27693 INVX1_LOC_89/Y NAND2X1_LOC_388/A 0.14fF
C27694 INVX1_LOC_117/Y INVX1_LOC_521/A 0.05fF
C27695 NAND2X1_LOC_388/A INVX1_LOC_154/A 0.00fF
C27696 INVX1_LOC_69/Y INVX1_LOC_66/A 0.03fF
C27697 INVX1_LOC_183/A INVX1_LOC_32/Y 0.03fF
C27698 INVX1_LOC_425/A INVX1_LOC_92/A 0.02fF
C27699 NAND2X1_LOC_260/Y NAND2X1_LOC_843/B 0.00fF
C27700 INVX1_LOC_309/Y INVX1_LOC_6/Y 0.02fF
C27701 NAND2X1_LOC_527/Y INVX1_LOC_26/Y 0.03fF
C27702 INVX1_LOC_204/Y NAND2X1_LOC_759/Y 0.00fF
C27703 INVX1_LOC_235/Y NAND2X1_LOC_271/A 0.05fF
C27704 INVX1_LOC_479/A INVX1_LOC_252/A 0.01fF
C27705 INVX1_LOC_106/Y NAND2X1_LOC_285/A 0.00fF
C27706 INVX1_LOC_49/Y NAND2X1_LOC_684/a_36_24# 0.01fF
C27707 INVX1_LOC_202/Y INVX1_LOC_91/A 0.03fF
C27708 INVX1_LOC_361/A INVX1_LOC_9/Y 0.07fF
C27709 INVX1_LOC_576/Y INVX1_LOC_636/A 0.04fF
C27710 INVX1_LOC_103/Y NAND2X1_LOC_372/Y 0.03fF
C27711 NAND2X1_LOC_60/Y INVX1_LOC_64/A 0.00fF
C27712 INVX1_LOC_642/Y NAND2X1_LOC_845/B 0.06fF
C27713 INVX1_LOC_203/Y INVX1_LOC_275/A 0.15fF
C27714 INVX1_LOC_69/Y NAND2X1_LOC_601/Y 0.03fF
C27715 NAND2X1_LOC_542/A INVX1_LOC_41/Y 0.02fF
C27716 NAND2X1_LOC_342/A INVX1_LOC_669/A 0.04fF
C27717 INPUT_6 INVX1_LOC_3/Y 0.84fF
C27718 INVX1_LOC_479/A INVX1_LOC_6/Y 0.09fF
C27719 INVX1_LOC_183/Y INVX1_LOC_85/A 0.71fF
C27720 INVX1_LOC_508/A NAND2X1_LOC_647/a_36_24# 0.00fF
C27721 INVX1_LOC_62/Y INVX1_LOC_361/A 0.14fF
C27722 INVX1_LOC_100/Y INVX1_LOC_664/A 0.33fF
C27723 INVX1_LOC_62/Y INVX1_LOC_196/Y 0.01fF
C27724 INVX1_LOC_41/Y INVX1_LOC_376/Y 0.02fF
C27725 INVX1_LOC_674/A INVX1_LOC_636/A 0.14fF
C27726 INVX1_LOC_102/Y INVX1_LOC_655/A 0.02fF
C27727 INVX1_LOC_15/Y INVX1_LOC_653/Y 0.01fF
C27728 INVX1_LOC_347/Y INVX1_LOC_354/A 0.00fF
C27729 INVX1_LOC_529/Y NAND2X1_LOC_668/Y 0.17fF
C27730 INVX1_LOC_426/Y INVX1_LOC_578/A 0.03fF
C27731 VDD INVX1_LOC_26/A -0.00fF
C27732 INVX1_LOC_438/Y INVX1_LOC_429/A 0.09fF
C27733 INVX1_LOC_206/Y NAND2X1_LOC_710/B 0.10fF
C27734 VDD INVX1_LOC_584/Y 0.42fF
C27735 INVX1_LOC_26/Y INVX1_LOC_621/A 0.07fF
C27736 INVX1_LOC_224/Y INVX1_LOC_560/A 0.01fF
C27737 INVX1_LOC_435/Y INVX1_LOC_445/A 0.02fF
C27738 INVX1_LOC_26/Y NAND2X1_LOC_85/a_36_24# 0.00fF
C27739 INVX1_LOC_242/Y INVX1_LOC_625/Y 0.02fF
C27740 INVX1_LOC_412/Y NAND2X1_LOC_354/a_36_24# 0.00fF
C27741 INVX1_LOC_114/A INVX1_LOC_634/Y 0.01fF
C27742 INVX1_LOC_206/Y INVX1_LOC_577/Y 0.02fF
C27743 INPUT_6 NAND2X1_LOC_2/a_36_24# 0.00fF
C27744 INPUT_0 NAND2X1_LOC_707/A 0.00fF
C27745 NAND2X1_LOC_164/Y INVX1_LOC_273/A 0.03fF
C27746 INVX1_LOC_92/Y INVX1_LOC_91/A 0.06fF
C27747 INVX1_LOC_158/A NAND2X1_LOC_180/B 0.00fF
C27748 NAND2X1_LOC_710/B INVX1_LOC_242/A 0.01fF
C27749 VDD INVX1_LOC_63/A 0.00fF
C27750 INVX1_LOC_380/A INVX1_LOC_35/Y 0.08fF
C27751 NAND2X1_LOC_373/Y INVX1_LOC_80/A 0.60fF
C27752 NAND2X1_LOC_503/B INVX1_LOC_604/Y 0.16fF
C27753 NAND2X1_LOC_269/B INVX1_LOC_231/Y 0.41fF
C27754 VDD NAND2X1_LOC_669/Y 0.07fF
C27755 VDD INVX1_LOC_449/A 0.00fF
C27756 INVX1_LOC_20/Y INVX1_LOC_319/Y 0.01fF
C27757 VDD INVX1_LOC_67/Y 0.22fF
C27758 INPUT_0 NAND2X1_LOC_336/B 0.03fF
C27759 INVX1_LOC_426/A INVX1_LOC_425/Y 0.03fF
C27760 INVX1_LOC_255/Y INVX1_LOC_686/A 0.08fF
C27761 INVX1_LOC_546/Y INVX1_LOC_134/Y 0.09fF
C27762 INVX1_LOC_113/Y INVX1_LOC_111/A 0.19fF
C27763 INVX1_LOC_31/Y INVX1_LOC_638/A 0.07fF
C27764 INVX1_LOC_614/A NAND2X1_LOC_153/a_36_24# 0.01fF
C27765 NAND2X1_LOC_24/Y INVX1_LOC_530/Y 0.56fF
C27766 VDD INVX1_LOC_195/Y 0.22fF
C27767 INVX1_LOC_206/Y INVX1_LOC_481/Y 0.09fF
C27768 INVX1_LOC_137/A NAND2X1_LOC_513/A 0.00fF
C27769 VDD INVX1_LOC_186/Y 0.66fF
C27770 NAND2X1_LOC_692/a_36_24# INVX1_LOC_367/A 0.00fF
C27771 INVX1_LOC_11/Y INVX1_LOC_553/A 0.05fF
C27772 INVX1_LOC_17/Y INVX1_LOC_552/Y -0.03fF
C27773 INVX1_LOC_319/Y INVX1_LOC_300/A 0.07fF
C27774 INVX1_LOC_618/A INVX1_LOC_624/Y 0.01fF
C27775 INVX1_LOC_603/Y INVX1_LOC_98/A 0.07fF
C27776 INVX1_LOC_224/Y INVX1_LOC_603/A 0.02fF
C27777 INVX1_LOC_400/Y INVX1_LOC_230/A 0.07fF
C27778 INVX1_LOC_20/Y INVX1_LOC_131/A 0.06fF
C27779 NAND2X1_LOC_331/A INVX1_LOC_500/Y 0.01fF
C27780 INVX1_LOC_76/Y INVX1_LOC_188/Y 0.00fF
C27781 INVX1_LOC_17/Y INVX1_LOC_374/A 0.00fF
C27782 INVX1_LOC_604/Y INVX1_LOC_273/A 0.02fF
C27783 INVX1_LOC_21/Y INVX1_LOC_94/A 0.18fF
C27784 INVX1_LOC_576/A INVX1_LOC_566/Y 0.03fF
C27785 NAND2X1_LOC_519/a_36_24# INVX1_LOC_367/Y 0.01fF
C27786 INVX1_LOC_603/Y INVX1_LOC_76/Y 0.02fF
C27787 INVX1_LOC_44/Y INVX1_LOC_275/A 0.07fF
C27788 INVX1_LOC_412/Y INVX1_LOC_469/Y 0.01fF
C27789 INVX1_LOC_412/Y INVX1_LOC_350/Y -0.00fF
C27790 NAND2X1_LOC_510/a_36_24# INVX1_LOC_397/A 0.00fF
C27791 INVX1_LOC_76/Y NAND2X1_LOC_645/a_36_24# 0.01fF
C27792 INVX1_LOC_26/Y NAND2X1_LOC_86/Y 0.01fF
C27793 INVX1_LOC_12/Y INVX1_LOC_486/Y 0.01fF
C27794 INVX1_LOC_35/Y NAND2X1_LOC_613/Y 0.01fF
C27795 INVX1_LOC_586/A INVX1_LOC_159/A 0.00fF
C27796 VDD INVX1_LOC_347/Y 0.51fF
C27797 INVX1_LOC_20/Y INVX1_LOC_432/Y 0.41fF
C27798 INVX1_LOC_395/A NAND2X1_LOC_308/A 0.06fF
C27799 INVX1_LOC_35/Y INVX1_LOC_169/A 0.03fF
C27800 INVX1_LOC_25/Y INVX1_LOC_55/Y 0.25fF
C27801 INVX1_LOC_300/A INVX1_LOC_566/Y 0.02fF
C27802 INVX1_LOC_405/A INVX1_LOC_502/A 0.21fF
C27803 INVX1_LOC_586/A NAND2X1_LOC_615/B 0.03fF
C27804 VDD INVX1_LOC_328/Y 0.59fF
C27805 NAND2X1_LOC_140/B INVX1_LOC_80/A 0.07fF
C27806 INVX1_LOC_80/A INVX1_LOC_600/Y 0.01fF
C27807 NAND2X1_LOC_387/Y INVX1_LOC_98/A 0.00fF
C27808 INVX1_LOC_361/Y NAND2X1_LOC_332/B 0.03fF
C27809 INVX1_LOC_134/Y INVX1_LOC_516/A 0.06fF
C27810 VDD INVX1_LOC_518/A 0.11fF
C27811 INVX1_LOC_197/Y NAND2X1_LOC_238/a_36_24# 0.01fF
C27812 NAND2X1_LOC_543/B NAND2X1_LOC_545/A 0.00fF
C27813 INVX1_LOC_595/A INVX1_LOC_6/A 0.01fF
C27814 INVX1_LOC_683/Y INVX1_LOC_665/Y 0.56fF
C27815 INVX1_LOC_17/Y INVX1_LOC_387/A 0.03fF
C27816 INVX1_LOC_442/A INVX1_LOC_69/Y 0.04fF
C27817 INVX1_LOC_307/A INVX1_LOC_145/Y 0.01fF
C27818 NAND2X1_LOC_97/B INVX1_LOC_59/Y 0.02fF
C27819 INVX1_LOC_267/Y INVX1_LOC_59/Y 0.01fF
C27820 INVX1_LOC_287/A INVX1_LOC_248/Y 0.37fF
C27821 INVX1_LOC_35/Y INVX1_LOC_633/Y 0.01fF
C27822 INVX1_LOC_605/A INVX1_LOC_58/Y 0.01fF
C27823 INVX1_LOC_126/A INPUT_1 0.08fF
C27824 INVX1_LOC_586/A INVX1_LOC_66/A 0.04fF
C27825 VDD INVX1_LOC_207/Y 0.33fF
C27826 INVX1_LOC_53/Y NAND2X1_LOC_708/A 0.12fF
C27827 INVX1_LOC_214/Y NAND2X1_LOC_496/Y 0.02fF
C27828 INVX1_LOC_206/Y INVX1_LOC_26/Y 16.08fF
C27829 INVX1_LOC_206/Y INVX1_LOC_128/Y 0.03fF
C27830 INVX1_LOC_412/Y INVX1_LOC_79/A 0.03fF
C27831 INVX1_LOC_442/Y INVX1_LOC_145/Y 0.07fF
C27832 INVX1_LOC_432/Y INVX1_LOC_300/A 0.01fF
C27833 INVX1_LOC_9/A INVX1_LOC_83/Y 0.01fF
C27834 NAND2X1_LOC_837/a_36_24# INVX1_LOC_50/Y 0.00fF
C27835 NAND2X1_LOC_97/B INVX1_LOC_48/Y 0.03fF
C27836 INVX1_LOC_11/Y NAND2X1_LOC_140/B 0.27fF
C27837 INVX1_LOC_578/A NAND2X1_LOC_605/B 0.03fF
C27838 INVX1_LOC_333/Y INVX1_LOC_40/Y 0.21fF
C27839 NAND2X1_LOC_368/a_36_24# INVX1_LOC_502/A 0.00fF
C27840 INVX1_LOC_410/Y INVX1_LOC_100/Y 0.07fF
C27841 INVX1_LOC_577/Y NAND2X1_LOC_334/A 0.03fF
C27842 INVX1_LOC_444/Y INVX1_LOC_452/A 0.02fF
C27843 INVX1_LOC_93/Y INVX1_LOC_134/Y 0.26fF
C27844 INVX1_LOC_193/A INVX1_LOC_99/A 0.06fF
C27845 INVX1_LOC_419/Y INVX1_LOC_129/A 0.07fF
C27846 VDD INVX1_LOC_597/Y 0.21fF
C27847 INVX1_LOC_312/Y INVX1_LOC_66/A 0.03fF
C27848 INVX1_LOC_54/Y INVX1_LOC_281/Y 0.01fF
C27849 INVX1_LOC_375/A INVX1_LOC_100/Y 0.03fF
C27850 INVX1_LOC_603/Y NAND2X1_LOC_503/Y 0.12fF
C27851 NAND2X1_LOC_790/B NAND2X1_LOC_98/B 0.18fF
C27852 INVX1_LOC_321/A NAND2X1_LOC_558/B 0.03fF
C27853 INVX1_LOC_492/A INVX1_LOC_556/Y 0.03fF
C27854 INVX1_LOC_504/A INVX1_LOC_513/A 0.28fF
C27855 INVX1_LOC_154/Y INVX1_LOC_32/Y 0.01fF
C27856 INVX1_LOC_510/A NAND2X1_LOC_649/a_36_24# 0.02fF
C27857 NAND2X1_LOC_757/a_36_24# INVX1_LOC_284/Y -0.00fF
C27858 INPUT_1 INVX1_LOC_252/Y 0.06fF
C27859 INVX1_LOC_54/Y INVX1_LOC_178/A 0.12fF
C27860 INVX1_LOC_12/Y INVX1_LOC_6/Y 0.09fF
C27861 INVX1_LOC_522/Y INVX1_LOC_507/Y 0.56fF
C27862 INVX1_LOC_76/Y INVX1_LOC_491/A 0.04fF
C27863 NAND2X1_LOC_403/A INVX1_LOC_46/Y 0.00fF
C27864 INVX1_LOC_379/A INVX1_LOC_490/A 0.15fF
C27865 INVX1_LOC_375/A INVX1_LOC_74/Y 0.03fF
C27866 INVX1_LOC_128/Y INVX1_LOC_242/A 0.03fF
C27867 INVX1_LOC_558/Y INVX1_LOC_199/Y 0.18fF
C27868 INVX1_LOC_166/A INVX1_LOC_251/A 0.01fF
C27869 INVX1_LOC_25/Y INVX1_LOC_18/Y 0.74fF
C27870 INVX1_LOC_675/A INVX1_LOC_134/Y 0.16fF
C27871 INVX1_LOC_586/A NAND2X1_LOC_601/Y 0.01fF
C27872 INVX1_LOC_372/Y NAND2X1_LOC_437/a_36_24# 0.00fF
C27873 NAND2X1_LOC_698/Y INVX1_LOC_600/A 0.03fF
C27874 INVX1_LOC_525/Y INVX1_LOC_59/Y 0.01fF
C27875 INVX1_LOC_63/Y NAND2X1_LOC_616/Y 0.30fF
C27876 INVX1_LOC_198/A INVX1_LOC_86/Y 0.01fF
C27877 INVX1_LOC_521/Y INVX1_LOC_645/Y 1.21fF
C27878 INVX1_LOC_545/A INVX1_LOC_253/Y 0.00fF
C27879 INVX1_LOC_269/A INVX1_LOC_92/Y 0.12fF
C27880 INVX1_LOC_686/A INVX1_LOC_26/Y 0.07fF
C27881 INVX1_LOC_293/Y NAND2X1_LOC_274/B 0.03fF
C27882 INVX1_LOC_54/Y INVX1_LOC_608/A 0.01fF
C27883 INVX1_LOC_676/Y INVX1_LOC_357/Y 0.05fF
C27884 INVX1_LOC_617/Y INVX1_LOC_79/A 0.02fF
C27885 INVX1_LOC_20/Y INVX1_LOC_319/A 0.43fF
C27886 INVX1_LOC_69/Y INVX1_LOC_116/Y 0.08fF
C27887 NAND2X1_LOC_507/A INVX1_LOC_117/Y 0.03fF
C27888 INVX1_LOC_131/A INVX1_LOC_655/A 0.02fF
C27889 INVX1_LOC_98/A INVX1_LOC_91/A 0.09fF
C27890 INVX1_LOC_525/Y INVX1_LOC_48/Y 0.07fF
C27891 INVX1_LOC_21/Y INVX1_LOC_376/Y 0.07fF
C27892 INVX1_LOC_514/A NAND2X1_LOC_828/a_36_24# 0.00fF
C27893 INVX1_LOC_607/Y NAND2X1_LOC_847/A 0.04fF
C27894 INVX1_LOC_519/Y INVX1_LOC_519/A 0.06fF
C27895 INVX1_LOC_76/Y INVX1_LOC_91/A 0.01fF
C27896 INVX1_LOC_20/Y NAND2X1_LOC_843/B 0.07fF
C27897 INVX1_LOC_89/Y INVX1_LOC_117/Y 0.10fF
C27898 INVX1_LOC_53/Y INVX1_LOC_369/Y 0.07fF
C27899 INVX1_LOC_63/Y INVX1_LOC_108/Y 0.02fF
C27900 INVX1_LOC_459/Y INVX1_LOC_348/Y 0.13fF
C27901 INVX1_LOC_31/Y NAND2X1_LOC_308/A 0.00fF
C27902 INVX1_LOC_54/Y INVX1_LOC_58/Y 0.77fF
C27903 INVX1_LOC_274/A NAND2X1_LOC_786/B 0.01fF
C27904 INVX1_LOC_47/Y INVX1_LOC_100/A 0.01fF
C27905 INVX1_LOC_93/Y INVX1_LOC_65/A 0.01fF
C27906 INVX1_LOC_20/Y INVX1_LOC_91/Y 0.08fF
C27907 INVX1_LOC_236/A INVX1_LOC_655/A 0.03fF
C27908 INVX1_LOC_672/Y INVX1_LOC_655/A 0.02fF
C27909 INVX1_LOC_117/Y INVX1_LOC_501/A 0.03fF
C27910 INVX1_LOC_435/A INVX1_LOC_90/Y 0.00fF
C27911 INVX1_LOC_300/A INVX1_LOC_319/A 0.01fF
C27912 INVX1_LOC_94/Y INVX1_LOC_96/A 0.01fF
C27913 INVX1_LOC_170/A INVX1_LOC_6/Y 0.35fF
C27914 INVX1_LOC_662/Y INVX1_LOC_100/Y 0.02fF
C27915 INVX1_LOC_255/A INVX1_LOC_69/Y 0.02fF
C27916 INVX1_LOC_361/Y INVX1_LOC_242/Y 0.03fF
C27917 INVX1_LOC_50/Y NAND2X1_LOC_436/a_36_24# 0.00fF
C27918 NAND2X1_LOC_334/A NAND2X1_LOC_290/a_36_24# 0.02fF
C27919 INVX1_LOC_507/Y INVX1_LOC_508/A 0.01fF
C27920 INVX1_LOC_521/A INVX1_LOC_58/Y 0.01fF
C27921 INVX1_LOC_166/A INVX1_LOC_652/A 0.02fF
C27922 INVX1_LOC_69/Y INVX1_LOC_179/A 4.41fF
C27923 INVX1_LOC_74/A INVX1_LOC_40/Y 0.29fF
C27924 INVX1_LOC_674/A INVX1_LOC_74/Y 0.07fF
C27925 INVX1_LOC_197/Y INVX1_LOC_91/Y 0.03fF
C27926 INVX1_LOC_680/A INVX1_LOC_6/Y 0.01fF
C27927 INVX1_LOC_623/Y INVX1_LOC_598/Y 0.02fF
C27928 NAND2X1_LOC_334/A INVX1_LOC_26/Y 0.33fF
C27929 INVX1_LOC_581/Y INVX1_LOC_62/Y 0.01fF
C27930 INVX1_LOC_460/Y INVX1_LOC_348/Y 0.04fF
C27931 INVX1_LOC_574/A NAND2X1_LOC_209/a_36_24# 0.00fF
C27932 INVX1_LOC_584/A INVX1_LOC_465/Y 0.00fF
C27933 VDD NAND2X1_LOC_763/Y -0.00fF
C27934 NAND2X1_LOC_121/Y INVX1_LOC_62/Y 0.04fF
C27935 NAND2X1_LOC_846/B INVX1_LOC_645/Y 0.09fF
C27936 INVX1_LOC_51/Y INVX1_LOC_638/A 0.07fF
C27937 INVX1_LOC_26/Y NAND2X1_LOC_609/B 0.01fF
C27938 VDD INVX1_LOC_521/Y 0.04fF
C27939 INVX1_LOC_557/Y INVX1_LOC_479/A 0.02fF
C27940 NAND2X1_LOC_301/B INVX1_LOC_62/Y 0.06fF
C27941 INVX1_LOC_238/Y INVX1_LOC_395/A 0.05fF
C27942 VDD INVX1_LOC_165/Y 0.21fF
C27943 INVX1_LOC_206/Y INVX1_LOC_560/A 0.07fF
C27944 NAND2X1_LOC_843/B INVX1_LOC_655/A 0.02fF
C27945 INVX1_LOC_206/Y NAND2X1_LOC_377/a_36_24# 0.00fF
C27946 INVX1_LOC_419/A INVX1_LOC_92/A 0.03fF
C27947 INVX1_LOC_369/Y INVX1_LOC_368/Y 0.01fF
C27948 VDD INVX1_LOC_266/Y 0.38fF
C27949 VDD INVX1_LOC_651/Y 0.75fF
C27950 NAND2X1_LOC_317/A INVX1_LOC_510/Y 0.02fF
C27951 INVX1_LOC_84/A INVX1_LOC_388/Y 0.00fF
C27952 INVX1_LOC_238/A INVX1_LOC_242/A 0.08fF
C27953 NAND2X1_LOC_248/B NAND2X1_LOC_247/a_36_24# 0.02fF
C27954 INVX1_LOC_371/A INVX1_LOC_109/Y 0.01fF
C27955 NAND2X1_LOC_751/a_36_24# INVX1_LOC_366/A 0.01fF
C27956 NAND2X1_LOC_498/Y INVX1_LOC_624/A 0.01fF
C27957 INVX1_LOC_224/Y INVX1_LOC_235/Y 0.22fF
C27958 INVX1_LOC_400/Y INVX1_LOC_666/A 0.02fF
C27959 INVX1_LOC_438/A INVX1_LOC_312/A 0.01fF
C27960 INVX1_LOC_442/A INVX1_LOC_586/A 0.04fF
C27961 NAND2X1_LOC_636/A INVX1_LOC_99/Y 0.01fF
C27962 INVX1_LOC_190/Y INVX1_LOC_184/A 0.14fF
C27963 INVX1_LOC_465/Y INVX1_LOC_537/A 0.19fF
C27964 INVX1_LOC_206/Y INVX1_LOC_369/A 0.03fF
C27965 INVX1_LOC_406/Y INVX1_LOC_450/A 0.00fF
C27966 INVX1_LOC_526/A INVX1_LOC_340/Y 0.06fF
C27967 INVX1_LOC_454/A INVX1_LOC_300/A 0.19fF
C27968 INVX1_LOC_395/A INVX1_LOC_134/Y 0.16fF
C27969 INVX1_LOC_133/Y INVX1_LOC_649/A 0.01fF
C27970 INVX1_LOC_401/Y NAND2X1_LOC_513/Y 0.05fF
C27971 INVX1_LOC_395/A NAND2X1_LOC_463/a_36_24# 0.00fF
C27972 INVX1_LOC_614/A INVX1_LOC_521/Y 0.12fF
C27973 INVX1_LOC_428/A INVX1_LOC_53/Y 0.03fF
C27974 VDD INVX1_LOC_335/A 0.02fF
C27975 INVX1_LOC_301/A INVX1_LOC_361/Y 1.24fF
C27976 INVX1_LOC_400/Y NAND2X1_LOC_325/B 1.28fF
C27977 NAND2X1_LOC_734/a_36_24# INVX1_LOC_300/A 0.00fF
C27978 INVX1_LOC_429/Y INVX1_LOC_385/Y 0.05fF
C27979 INPUT_3 INVX1_LOC_172/Y 0.01fF
C27980 VDD INVX1_LOC_105/Y 0.68fF
C27981 INVX1_LOC_459/A INVX1_LOC_47/Y 0.05fF
C27982 INVX1_LOC_567/A INVX1_LOC_66/A 0.05fF
C27983 INVX1_LOC_384/A NAND2X1_LOC_272/a_36_24# 0.01fF
C27984 INVX1_LOC_412/Y INVX1_LOC_48/Y 0.03fF
C27985 INVX1_LOC_268/A INVX1_LOC_586/A 0.01fF
C27986 VDD GATE_662 0.04fF
C27987 NAND2X1_LOC_503/B INVX1_LOC_63/Y 0.93fF
C27988 INVX1_LOC_510/Y INVX1_LOC_352/A 0.01fF
C27989 INVX1_LOC_317/Y INVX1_LOC_35/Y 0.00fF
C27990 NAND2X1_LOC_176/Y NAND2X1_LOC_388/A 0.28fF
C27991 NAND2X1_LOC_707/A INVX1_LOC_145/Y 0.07fF
C27992 INVX1_LOC_683/Y INVX1_LOC_134/Y 0.02fF
C27993 INVX1_LOC_531/A INVX1_LOC_169/A 0.01fF
C27994 INVX1_LOC_586/A INVX1_LOC_116/Y 0.10fF
C27995 NAND2X1_LOC_525/Y INVX1_LOC_413/A 0.07fF
C27996 INVX1_LOC_455/A INVX1_LOC_45/Y 0.00fF
C27997 INVX1_LOC_417/Y INVX1_LOC_119/A 0.03fF
C27998 INVX1_LOC_76/Y INVX1_LOC_504/Y 0.07fF
C27999 INVX1_LOC_375/A INVX1_LOC_350/Y 0.12fF
C28000 NAND2X1_LOC_534/Y INVX1_LOC_58/Y 0.00fF
C28001 INVX1_LOC_17/Y NAND2X1_LOC_620/a_36_24# 0.00fF
C28002 INVX1_LOC_51/Y INVX1_LOC_665/Y 0.03fF
C28003 VDD NAND2X1_LOC_846/B 0.66fF
C28004 INVX1_LOC_211/Y INVX1_LOC_482/A 0.06fF
C28005 INVX1_LOC_53/Y INVX1_LOC_558/Y 0.06fF
C28006 INVX1_LOC_45/Y INVX1_LOC_345/A 0.01fF
C28007 INVX1_LOC_459/A INVX1_LOC_119/Y 0.07fF
C28008 INVX1_LOC_308/Y INVX1_LOC_47/Y 0.03fF
C28009 INVX1_LOC_321/A INVX1_LOC_48/Y 0.04fF
C28010 NAND2X1_LOC_843/A INVX1_LOC_651/Y 0.18fF
C28011 NAND2X1_LOC_548/B INVX1_LOC_99/Y 0.03fF
C28012 INVX1_LOC_17/Y INVX1_LOC_84/A 0.11fF
C28013 INVX1_LOC_357/A INVX1_LOC_495/A 0.02fF
C28014 INVX1_LOC_324/Y INVX1_LOC_7/Y 0.05fF
C28015 INVX1_LOC_312/Y INVX1_LOC_116/Y 0.03fF
C28016 INVX1_LOC_606/Y INVX1_LOC_199/Y 0.03fF
C28017 INVX1_LOC_312/Y INVX1_LOC_544/A 0.03fF
C28018 INVX1_LOC_400/A INVX1_LOC_318/Y 0.00fF
C28019 INVX1_LOC_438/A INVX1_LOC_226/Y 0.01fF
C28020 INVX1_LOC_159/A INVX1_LOC_486/Y 0.03fF
C28021 INVX1_LOC_20/Y NAND2X1_LOC_333/B 0.14fF
C28022 NAND2X1_LOC_308/A INVX1_LOC_51/Y 0.21fF
C28023 INVX1_LOC_20/Y INVX1_LOC_361/Y 0.38fF
C28024 INVX1_LOC_99/Y NAND2X1_LOC_237/Y 0.01fF
C28025 INVX1_LOC_566/A INVX1_LOC_674/A 0.01fF
C28026 INVX1_LOC_378/A INVX1_LOC_46/Y 0.03fF
C28027 INVX1_LOC_370/A INVX1_LOC_519/A 0.01fF
C28028 INVX1_LOC_43/Y INVX1_LOC_7/Y 0.00fF
C28029 NAND2X1_LOC_370/A INVX1_LOC_63/Y 0.01fF
C28030 INVX1_LOC_150/Y INVX1_LOC_58/Y 0.01fF
C28031 INVX1_LOC_297/A INVX1_LOC_50/Y 0.58fF
C28032 INVX1_LOC_586/A INVX1_LOC_255/A 0.03fF
C28033 INVX1_LOC_17/Y NAND2X1_LOC_67/Y 0.03fF
C28034 INVX1_LOC_99/Y INVX1_LOC_230/A 0.08fF
C28035 INVX1_LOC_410/Y INVX1_LOC_79/A 0.03fF
C28036 GATE_579 GATE_479 0.04fF
C28037 INVX1_LOC_568/Y INVX1_LOC_556/Y 0.04fF
C28038 INVX1_LOC_273/A INVX1_LOC_63/Y 0.01fF
C28039 INVX1_LOC_160/A INVX1_LOC_159/Y 0.01fF
C28040 INVX1_LOC_31/Y INVX1_LOC_134/Y 0.16fF
C28041 INVX1_LOC_364/Y INVX1_LOC_682/Y 0.15fF
C28042 INVX1_LOC_375/A INVX1_LOC_79/A 1.68fF
C28043 INVX1_LOC_397/A INVX1_LOC_26/Y 0.01fF
C28044 INVX1_LOC_586/A NAND2X1_LOC_719/A 0.02fF
C28045 INVX1_LOC_603/Y INVX1_LOC_32/Y 0.03fF
C28046 INVX1_LOC_45/Y NAND2X1_LOC_823/Y 0.10fF
C28047 NAND2X1_LOC_820/A INVX1_LOC_66/A 0.03fF
C28048 INVX1_LOC_671/A NAND2X1_LOC_260/Y 0.03fF
C28049 NAND2X1_LOC_106/Y INVX1_LOC_80/A 0.01fF
C28050 INVX1_LOC_546/A INVX1_LOC_79/A 0.04fF
C28051 NAND2X1_LOC_121/a_36_24# INVX1_LOC_497/A 0.00fF
C28052 INVX1_LOC_522/Y INVX1_LOC_508/A 0.02fF
C28053 NAND2X1_LOC_775/B INVX1_LOC_350/A 0.03fF
C28054 INVX1_LOC_63/A NAND2X1_LOC_824/a_36_24# 0.00fF
C28055 INVX1_LOC_585/Y INVX1_LOC_178/A 0.01fF
C28056 INVX1_LOC_589/Y NAND2X1_LOC_237/Y 0.01fF
C28057 INVX1_LOC_197/Y NAND2X1_LOC_333/B 0.07fF
C28058 INVX1_LOC_468/Y INVX1_LOC_506/A 0.01fF
C28059 INVX1_LOC_551/Y INVX1_LOC_9/Y 0.11fF
C28060 INVX1_LOC_599/Y INVX1_LOC_292/Y 0.00fF
C28061 NAND2X1_LOC_526/Y INVX1_LOC_41/Y 0.01fF
C28062 INVX1_LOC_166/A INVX1_LOC_35/Y 0.07fF
C28063 INVX1_LOC_614/A NAND2X1_LOC_846/B 0.03fF
C28064 INVX1_LOC_117/Y INVX1_LOC_194/Y 0.00fF
C28065 INVX1_LOC_45/Y INVX1_LOC_280/A 0.28fF
C28066 NAND2X1_LOC_413/Y INVX1_LOC_199/Y 0.37fF
C28067 INVX1_LOC_387/Y INVX1_LOC_453/Y 0.02fF
C28068 INVX1_LOC_686/A NAND2X1_LOC_605/B 0.05fF
C28069 INVX1_LOC_134/Y INVX1_LOC_682/Y 0.01fF
C28070 INVX1_LOC_11/Y NAND2X1_LOC_106/Y 0.06fF
C28071 INVX1_LOC_89/Y INVX1_LOC_251/Y 0.66fF
C28072 INVX1_LOC_63/Y NAND2X1_LOC_393/Y 0.01fF
C28073 INVX1_LOC_524/Y INVX1_LOC_90/Y 0.01fF
C28074 NAND2X1_LOC_304/a_36_24# INVX1_LOC_9/Y -0.02fF
C28075 INVX1_LOC_47/Y INVX1_LOC_230/A 0.10fF
C28076 INVX1_LOC_53/Y NAND2X1_LOC_106/a_36_24# 0.01fF
C28077 NAND2X1_LOC_387/Y INVX1_LOC_32/Y 0.16fF
C28078 INVX1_LOC_435/Y INVX1_LOC_282/Y 0.05fF
C28079 NAND2X1_LOC_548/B NAND2X1_LOC_66/Y 0.07fF
C28080 INVX1_LOC_551/Y INVX1_LOC_62/Y 0.03fF
C28081 INVX1_LOC_360/Y INVX1_LOC_347/Y 0.01fF
C28082 INVX1_LOC_6/Y NAND2X1_LOC_615/B 0.00fF
C28083 INPUT_3 INVX1_LOC_280/A 0.00fF
C28084 INVX1_LOC_419/A INPUT_1 0.02fF
C28085 NAND2X1_LOC_709/a_36_24# INVX1_LOC_35/Y 0.00fF
C28086 INVX1_LOC_49/Y INVX1_LOC_259/Y 0.03fF
C28087 INVX1_LOC_662/A NAND2X1_LOC_148/a_36_24# 0.01fF
C28088 NAND2X1_LOC_260/Y INVX1_LOC_664/Y 0.01fF
C28089 NAND2X1_LOC_827/Y INVX1_LOC_50/Y 0.02fF
C28090 INVX1_LOC_277/A INVX1_LOC_58/Y 0.01fF
C28091 INVX1_LOC_80/A NAND2X1_LOC_123/B 0.04fF
C28092 INVX1_LOC_619/A INVX1_LOC_207/Y 0.05fF
C28093 INVX1_LOC_585/Y INVX1_LOC_58/Y 0.01fF
C28094 INVX1_LOC_400/A INVX1_LOC_351/A 0.01fF
C28095 INVX1_LOC_533/A INVX1_LOC_259/Y 0.17fF
C28096 INVX1_LOC_555/A INVX1_LOC_477/Y 0.02fF
C28097 INVX1_LOC_6/Y INVX1_LOC_66/A 0.57fF
C28098 INVX1_LOC_117/Y INVX1_LOC_44/Y 0.16fF
C28099 INVX1_LOC_283/Y INVX1_LOC_671/Y 0.96fF
C28100 NAND2X1_LOC_707/B INVX1_LOC_49/Y 0.01fF
C28101 NAND2X1_LOC_686/A INVX1_LOC_513/A 0.02fF
C28102 INVX1_LOC_400/A INVX1_LOC_90/Y 0.01fF
C28103 INVX1_LOC_54/Y INVX1_LOC_245/A 0.06fF
C28104 INVX1_LOC_89/Y INVX1_LOC_58/Y 0.42fF
C28105 INVX1_LOC_35/Y INVX1_LOC_531/Y 0.09fF
C28106 INVX1_LOC_32/Y NAND2X1_LOC_845/B 0.02fF
C28107 INVX1_LOC_11/Y NAND2X1_LOC_123/B 0.03fF
C28108 VDD INVX1_LOC_109/Y 0.52fF
C28109 INVX1_LOC_674/A INVX1_LOC_79/A 0.19fF
C28110 INVX1_LOC_80/A INVX1_LOC_270/Y 0.03fF
C28111 NAND2X1_LOC_3/a_36_24# INVX1_LOC_25/A 0.01fF
C28112 INVX1_LOC_46/Y INVX1_LOC_422/A 0.03fF
C28113 INVX1_LOC_93/Y INVX1_LOC_90/Y 0.05fF
C28114 INVX1_LOC_167/A INVX1_LOC_166/Y 0.00fF
C28115 INVX1_LOC_178/Y INVX1_LOC_6/Y 0.01fF
C28116 INVX1_LOC_501/A INVX1_LOC_58/Y 0.00fF
C28117 INVX1_LOC_304/Y INVX1_LOC_75/Y 0.06fF
C28118 INVX1_LOC_62/Y INVX1_LOC_493/A 0.03fF
C28119 INVX1_LOC_35/Y INVX1_LOC_528/Y 0.05fF
C28120 INVX1_LOC_167/A INVX1_LOC_62/Y 0.16fF
C28121 NAND2X1_LOC_836/B INVX1_LOC_35/A 0.03fF
C28122 VDD INVX1_LOC_95/Y 0.26fF
C28123 INVX1_LOC_254/Y INVX1_LOC_74/Y 0.01fF
C28124 INVX1_LOC_80/A INVX1_LOC_92/A 0.05fF
C28125 NAND2X1_LOC_542/A INVX1_LOC_128/Y 0.03fF
C28126 INVX1_LOC_531/Y INVX1_LOC_620/A 0.07fF
C28127 VDD INVX1_LOC_554/A 0.25fF
C28128 INVX1_LOC_49/Y INVX1_LOC_114/A 0.09fF
C28129 INVX1_LOC_32/Y INVX1_LOC_91/A 0.03fF
C28130 INVX1_LOC_62/Y NAND2X1_LOC_252/Y 0.16fF
C28131 INVX1_LOC_11/Y INVX1_LOC_270/Y 0.03fF
C28132 NAND2X1_LOC_790/B INVX1_LOC_206/Y 0.41fF
C28133 INVX1_LOC_128/Y INVX1_LOC_376/Y 0.02fF
C28134 INVX1_LOC_199/Y NAND2X1_LOC_488/Y 0.00fF
C28135 INVX1_LOC_434/A INVX1_LOC_453/A 0.00fF
C28136 INVX1_LOC_11/Y INVX1_LOC_92/A 0.07fF
C28137 INVX1_LOC_490/A INVX1_LOC_488/Y 0.12fF
C28138 INVX1_LOC_77/Y INVX1_LOC_211/A 0.03fF
C28139 NAND2X1_LOC_433/Y NAND2X1_LOC_123/B 0.99fF
C28140 INVX1_LOC_500/A INVX1_LOC_62/Y 0.04fF
C28141 NAND2X1_LOC_410/Y INVX1_LOC_9/Y 0.00fF
C28142 NAND2X1_LOC_710/B INVX1_LOC_121/Y 0.02fF
C28143 NAND2X1_LOC_333/A INVX1_LOC_636/A 0.01fF
C28144 INVX1_LOC_85/Y INVX1_LOC_181/A 0.15fF
C28145 INVX1_LOC_390/Y INVX1_LOC_560/A 0.32fF
C28146 INVX1_LOC_100/Y INVX1_LOC_479/A 6.03fF
C28147 INVX1_LOC_184/Y INVX1_LOC_190/A 0.20fF
C28148 VDD NAND2X1_LOC_427/Y 0.01fF
C28149 NAND2X1_LOC_789/B INVX1_LOC_85/Y 0.01fF
C28150 VDD NAND2X1_LOC_79/Y -0.00fF
C28151 INVX1_LOC_614/A INVX1_LOC_554/A 0.02fF
C28152 INVX1_LOC_662/A INVX1_LOC_240/Y 0.04fF
C28153 NAND2X1_LOC_475/A NAND2X1_LOC_492/a_36_24# 0.00fF
C28154 VDD INVX1_LOC_126/Y 0.43fF
C28155 INVX1_LOC_479/A INVX1_LOC_74/Y 0.13fF
C28156 INVX1_LOC_584/Y INVX1_LOC_45/Y 0.01fF
C28157 INVX1_LOC_206/Y INVX1_LOC_235/Y 0.01fF
C28158 INVX1_LOC_362/Y NAND2X1_LOC_249/a_36_24# 0.00fF
C28159 INVX1_LOC_616/Y VSS 0.13fF
C28160 INVX1_LOC_638/A VSS 1.13fF
C28161 INVX1_LOC_610/Y VSS 0.04fF
C28162 INVX1_LOC_624/A VSS 0.12fF
C28163 INVX1_LOC_618/Y VSS -0.10fF
C28164 NAND2X1_LOC_749/Y VSS 0.20fF
C28165 INVX1_LOC_596/Y VSS 0.14fF
C28166 INVX1_LOC_388/Y VSS 0.58fF
C28167 NAND2X1_LOC_801/A VSS 0.29fF
C28168 NAND2X1_LOC_226/Y VSS 0.08fF
C28169 INVX1_LOC_216/Y VSS 0.06fF
C28170 INVX1_LOC_215/Y VSS 0.25fF
C28171 INVX1_LOC_181/A VSS 0.16fF
C28172 INVX1_LOC_180/Y VSS 0.08fF
C28173 INVX1_LOC_192/A VSS 0.12fF
C28174 INVX1_LOC_109/Y VSS 0.40fF
C28175 INVX1_LOC_98/Y VSS 0.90fF
C28176 INVX1_LOC_333/A VSS 0.25fF
C28177 INVX1_LOC_334/Y VSS 0.25fF
C28178 NAND2X1_LOC_506/B VSS 0.47fF
C28179 NAND2X1_LOC_86/Y VSS 0.06fF
C28180 INVX1_LOC_41/A VSS 0.12fF
C28181 INVX1_LOC_1/Y VSS 0.58fF
C28182 INVX1_LOC_69/A VSS 0.23fF
C28183 INVX1_LOC_29/Y VSS 0.64fF
C28184 INVX1_LOC_59/A VSS 0.39fF
C28185 INVX1_LOC_55/Y VSS 0.41fF
C28186 INVX1_LOC_60/Y VSS 0.25fF
C28187 INVX1_LOC_94/A VSS 0.55fF
C28188 INVX1_LOC_49/A VSS 0.12fF
C28189 NAND2X1_LOC_76/B VSS 0.34fF
C28190 INVX1_LOC_275/A VSS 0.41fF
C28191 INVX1_LOC_297/Y VSS 0.40fF
C28192 INVX1_LOC_242/A VSS 0.08fF
C28193 INVX1_LOC_253/A VSS 0.35fF
C28194 INVX1_LOC_220/A VSS -0.27fF
C28195 INVX1_LOC_423/Y VSS 0.20fF
C28196 INVX1_LOC_423/A VSS 0.02fF
C28197 INVX1_LOC_489/Y VSS 0.23fF
C28198 INVX1_LOC_445/A VSS 0.23fF
C28199 NAND2X1_LOC_591/B VSS 0.07fF
C28200 INVX1_LOC_458/Y VSS 0.06fF
C28201 INVX1_LOC_615/Y VSS 0.25fF
C28202 INVX1_LOC_615/A VSS 0.13fF
C28203 INVX1_LOC_648/Y VSS 0.06fF
C28204 INVX1_LOC_395/A VSS 1.09fF
C28205 INVX1_LOC_626/Y VSS 0.11fF
C28206 INVX1_LOC_623/A VSS 0.12fF
C28207 INVX1_LOC_620/Y VSS 0.34fF
C28208 INVX1_LOC_619/Y VSS 0.25fF
C28209 INVX1_LOC_597/Y VSS 0.23fF
C28210 NAND2X1_LOC_800/B VSS 0.25fF
C28211 INVX1_LOC_182/Y VSS 0.04fF
C28212 INVX1_LOC_181/Y VSS 0.07fF
C28213 NAND2X1_LOC_342/B VSS 0.23fF
C28214 NAND2X1_LOC_258/Y VSS 0.08fF
C28215 INVX1_LOC_342/A VSS 0.15fF
C28216 INVX1_LOC_343/Y VSS 0.23fF
C28217 INVX1_LOC_332/Y VSS 0.19fF
C28218 INVX1_LOC_86/A VSS 0.30fF
C28219 INVX1_LOC_40/A VSS 0.12fF
C28220 NAND2X1_LOC_52/Y VSS 0.31fF
C28221 INVX1_LOC_68/A VSS 0.12fF
C28222 NAND2X1_LOC_76/A VSS 0.19fF
C28223 NAND2X1_LOC_98/B VSS 0.28fF
C28224 INVX1_LOC_91/Y VSS 0.37fF
C28225 INVX1_LOC_274/Y VSS 0.17fF
C28226 INVX1_LOC_296/A VSS 0.47fF
C28227 INVX1_LOC_230/Y VSS 0.35fF
C28228 INVX1_LOC_263/Y VSS 0.14fF
C28229 INVX1_LOC_259/Y VSS -0.36fF
C28230 INVX1_LOC_252/Y VSS 0.21fF
C28231 INVX1_LOC_252/A VSS 0.35fF
C28232 INVX1_LOC_488/Y VSS 0.51fF
C28233 INVX1_LOC_422/A VSS 0.10fF
C28234 INVX1_LOC_411/Y VSS 0.29fF
C28235 INVX1_LOC_433/A VSS -0.07fF
C28236 INVX1_LOC_444/A VSS 0.06fF
C28237 INVX1_LOC_505/A VSS 0.25fF
C28238 INVX1_LOC_92/A VSS -1.86fF
C28239 INVX1_LOC_658/Y VSS 0.19fF
C28240 INVX1_LOC_669/A VSS 0.52fF
C28241 INVX1_LOC_9/Y VSS 1.01fF
C28242 INVX1_LOC_3/A VSS 0.12fF
C28243 INVX1_LOC_603/A VSS 0.42fF
C28244 INVX1_LOC_636/Y VSS 0.04fF
C28245 INVX1_LOC_636/A VSS 0.74fF
C28246 INVX1_LOC_625/Y VSS 0.33fF
C28247 INVX1_LOC_614/Y VSS 0.10fF
C28248 INVX1_LOC_622/A VSS 0.12fF
C28249 INVX1_LOC_621/Y VSS 0.13fF
C28250 NAND2X1_LOC_759/Y VSS 0.28fF
C28251 INVX1_LOC_611/A VSS 0.32fF
C28252 INVX1_LOC_190/A VSS 0.20fF
C28253 INVX1_LOC_184/Y VSS 0.04fF
C28254 INVX1_LOC_206/A VSS 0.12fF
C28255 NAND2X1_LOC_271/A VSS 0.07fF
C28256 INVX1_LOC_231/Y VSS 0.15fF
C28257 NAND2X1_LOC_248/B VSS 0.44fF
C28258 INVX1_LOC_199/A VSS 0.12fF
C28259 INVX1_LOC_347/A VSS -0.49fF
C28260 INVX1_LOC_85/A VSS -1.04fF
C28261 NAND2X1_LOC_81/Y VSS -0.05fF
C28262 INVX1_LOC_93/A VSS 0.02fF
C28263 INVX1_LOC_18/Y VSS 0.60fF
C28264 INVX1_LOC_58/A VSS 0.12fF
C28265 INVX1_LOC_40/Y VSS 0.40fF
C28266 INVX1_LOC_76/A VSS 0.12fF
C28267 INVX1_LOC_66/Y VSS 0.25fF
C28268 INVX1_LOC_273/Y VSS 0.39fF
C28269 INVX1_LOC_284/Y VSS 0.13fF
C28270 INPUT_4 VSS 0.30fF
C28271 INVX1_LOC_295/Y VSS 0.22fF
C28272 INVX1_LOC_251/Y VSS 0.49fF
C28273 INVX1_LOC_240/Y VSS 0.25fF
C28274 NAND2X1_LOC_646/B VSS 0.25fF
C28275 INVX1_LOC_454/Y VSS 0.28fF
C28276 INVX1_LOC_245/A VSS -7.06fF
C28277 INVX1_LOC_498/Y VSS 0.30fF
C28278 INVX1_LOC_476/Y VSS 0.36fF
C28279 INVX1_LOC_432/A VSS 0.16fF
C28280 INVX1_LOC_443/Y VSS 0.25fF
C28281 INVX1_LOC_443/A VSS -9.61fF
C28282 INVX1_LOC_635/Y VSS -0.15fF
C28283 INVX1_LOC_624/Y VSS 0.23fF
C28284 INVX1_LOC_668/Y VSS 0.04fF
C28285 INVX1_LOC_613/A VSS 0.15fF
C28286 NAND2X1_LOC_284/A VSS 0.19fF
C28287 NAND2X1_LOC_243/A VSS 0.43fF
C28288 INVX1_LOC_86/Y VSS 0.53fF
C28289 INVX1_LOC_178/A VSS 0.86fF
C28290 NAND2X1_LOC_69/Y VSS 0.11fF
C28291 NAND2X1_LOC_67/Y VSS 0.25fF
C28292 NAND2X1_LOC_227/A VSS 0.19fF
C28293 NAND2X1_LOC_269/B VSS 0.18fF
C28294 INVX1_LOC_90/Y VSS 0.45fF
C28295 NAND2X1_LOC_342/A VSS 0.15fF
C28296 INVX1_LOC_212/Y VSS 0.32fF
C28297 INVX1_LOC_66/A VSS 0.23fF
C28298 INVX1_LOC_189/A VSS 0.09fF
C28299 INVX1_LOC_186/Y VSS -0.96fF
C28300 NAND2X1_LOC_259/A VSS 0.21fF
C28301 NAND2X1_LOC_832/A VSS 0.38fF
C28302 NAND2X1_LOC_544/B VSS 0.24fF
C28303 NAND2X1_LOC_406/B VSS 0.11fF
C28304 NAND2X1_LOC_84/B VSS 0.44fF
C28305 INVX1_LOC_83/Y VSS 0.27fF
C28306 NAND2X1_LOC_72/Y VSS -0.02fF
C28307 INVX1_LOC_91/A VSS 0.28fF
C28308 INVX1_LOC_92/Y VSS 0.24fF
C28309 INVX1_LOC_272/A VSS 0.29fF
C28310 INVX1_LOC_283/A VSS -0.05fF
C28311 INVX1_LOC_56/Y VSS 0.25fF
C28312 INVX1_LOC_64/A VSS 0.05fF
C28313 NAND2X1_LOC_60/Y VSS 0.14fF
C28314 NAND2X1_LOC_609/B VSS 0.36fF
C28315 INVX1_LOC_473/Y VSS -0.03fF
C28316 INVX1_LOC_486/A VSS 0.14fF
C28317 INVX1_LOC_431/Y VSS 0.26fF
C28318 INVX1_LOC_497/Y VSS 0.21fF
C28319 INVX1_LOC_453/Y VSS 0.59fF
C28320 INVX1_LOC_464/Y VSS 0.26fF
C28321 INVX1_LOC_475/Y VSS -0.31fF
C28322 INVX1_LOC_420/A VSS 0.18fF
C28323 INVX1_LOC_601/Y VSS 0.01fF
C28324 INVX1_LOC_623/Y VSS 0.19fF
C28325 INVX1_LOC_656/Y VSS 0.22fF
C28326 INVX1_LOC_634/Y VSS 0.54fF
C28327 INVX1_LOC_645/Y VSS 0.08fF
C28328 INVX1_LOC_588/A VSS -0.43fF
C28329 INVX1_LOC_667/A VSS 0.12fF
C28330 INVX1_LOC_612/A VSS 0.27fF
C28331 NAND2X1_LOC_753/Y VSS -0.48fF
C28332 NAND2X1_LOC_333/B VSS 0.40fF
C28333 INVX1_LOC_230/A VSS -0.46fF
C28334 INVX1_LOC_212/A VSS 0.26fF
C28335 NAND2X1_LOC_344/B VSS 0.31fF
C28336 GATE_222 VSS -0.01fF
C28337 INVX1_LOC_197/Y VSS 0.30fF
C28338 INVX1_LOC_64/Y VSS 0.36fF
C28339 INVX1_LOC_188/A VSS 0.26fF
C28340 INVX1_LOC_187/Y VSS 0.33fF
C28341 INVX1_LOC_328/A VSS 0.30fF
C28342 INVX1_LOC_327/Y VSS 0.12fF
C28343 INVX1_LOC_365/A VSS 0.12fF
C28344 NAND2X1_LOC_378/Y VSS -0.20fF
C28345 NAND2X1_LOC_376/Y VSS 0.17fF
C28346 NAND2X1_LOC_416/B VSS 0.27fF
C28347 INVX1_LOC_354/A VSS 0.39fF
C28348 INVX1_LOC_114/A VSS 0.47fF
C28349 NAND2X1_LOC_440/A VSS 0.19fF
C28350 INVX1_LOC_83/A VSS 0.12fF
C28351 INVX1_LOC_84/Y VSS 0.11fF
C28352 INVX1_LOC_75/A VSS 0.46fF
C28353 INVX1_LOC_260/Y VSS 0.25fF
C28354 INVX1_LOC_282/Y VSS 0.25fF
C28355 INVX1_LOC_487/A VSS 0.30fF
C28356 NAND2X1_LOC_627/Y VSS 0.07fF
C28357 NAND2X1_LOC_626/Y VSS 0.22fF
C28358 INVX1_LOC_480/A VSS 0.12fF
C28359 NAND2X1_LOC_646/A VSS 0.31fF
C28360 NAND2X1_LOC_606/Y VSS 0.23fF
C28361 INVX1_LOC_485/A VSS 0.05fF
C28362 INVX1_LOC_441/A VSS 0.12fF
C28363 INVX1_LOC_430/Y VSS 0.19fF
C28364 INVX1_LOC_430/A VSS 0.28fF
C28365 INVX1_LOC_496/Y VSS -0.10fF
C28366 INVX1_LOC_48/Y VSS 0.66fF
C28367 INVX1_LOC_600/Y VSS -0.12fF
C28368 INVX1_LOC_600/A VSS -1.53fF
C28369 INVX1_LOC_622/Y VSS 0.25fF
C28370 INVX1_LOC_666/Y VSS 0.11fF
C28371 INVX1_LOC_655/A VSS -3.10fF
C28372 INVX1_LOC_611/Y VSS 0.04fF
C28373 INVX1_LOC_198/A VSS -1.01fF
C28374 INVX1_LOC_195/Y VSS 0.34fF
C28375 INVX1_LOC_194/Y VSS 0.57fF
C28376 INVX1_LOC_228/A VSS 0.17fF
C28377 INVX1_LOC_211/A VSS -1.53fF
C28378 INVX1_LOC_209/Y VSS 0.10fF
C28379 INVX1_LOC_204/A VSS 0.12fF
C28380 INVX1_LOC_46/Y VSS 0.54fF
C28381 INVX1_LOC_241/Y VSS 0.18fF
C28382 INVX1_LOC_169/Y VSS 0.66fF
C28383 INVX1_LOC_155/Y VSS 0.60fF
C28384 INVX1_LOC_327/A VSS 0.12fF
C28385 INVX1_LOC_353/A VSS 0.40fF
C28386 NAND2X1_LOC_420/Y VSS 0.07fF
C28387 INVX1_LOC_340/A VSS 0.37fF
C28388 INVX1_LOC_341/Y VSS 0.12fF
C28389 NAND2X1_LOC_415/B VSS -0.08fF
C28390 INVX1_LOC_7/Y VSS 0.81fF
C28391 INVX1_LOC_364/A VSS 0.23fF
C28392 NAND2X1_LOC_372/Y VSS 0.36fF
C28393 INVX1_LOC_374/Y VSS -0.23fF
C28394 INVX1_LOC_350/Y VSS 0.16fF
C28395 INVX1_LOC_74/A VSS 0.22fF
C28396 INVX1_LOC_292/Y VSS 0.40fF
C28397 INVX1_LOC_18/A VSS 0.12fF
C28398 INVX1_LOC_29/A VSS 0.13fF
C28399 INVX1_LOC_281/Y VSS 0.30fF
C28400 INVX1_LOC_270/Y VSS 0.40fF
C28401 NAND2X1_LOC_621/B VSS 0.17fF
C28402 INVX1_LOC_499/A VSS -0.13fF
C28403 INVX1_LOC_470/Y VSS 0.23fF
C28404 INVX1_LOC_440/Y VSS 0.31fF
C28405 INVX1_LOC_440/A VSS 0.12fF
C28406 INVX1_LOC_451/Y VSS 0.04fF
C28407 INVX1_LOC_462/Y VSS 0.19fF
C28408 INVX1_LOC_495/Y VSS 0.08fF
C28409 INVX1_LOC_639/A VSS 0.09fF
C28410 INVX1_LOC_631/Y VSS 0.25fF
C28411 INVX1_LOC_665/Y VSS 0.07fF
C28412 INVX1_LOC_676/A VSS 0.19fF
C28413 INVX1_LOC_621/A VSS 0.24fF
C28414 INVX1_LOC_632/Y VSS 0.25fF
C28415 INVX1_LOC_654/Y VSS 0.31fF
C28416 INVX1_LOC_610/A VSS -0.05fF
C28417 INVX1_LOC_109/A VSS -0.04fF
C28418 INVX1_LOC_210/A VSS 0.21fF
C28419 INVX1_LOC_207/Y VSS 0.29fF
C28420 NAND2X1_LOC_240/A VSS 0.19fF
C28421 NAND2X1_LOC_267/A VSS 0.44fF
C28422 INVX1_LOC_227/Y VSS 0.06fF
C28423 INVX1_LOC_235/A VSS 0.12fF
C28424 NAND2X1_LOC_275/Y VSS 0.23fF
C28425 NAND2X1_LOC_302/A VSS 0.19fF
C28426 INVX1_LOC_241/A VSS 0.34fF
C28427 NAND2X1_LOC_843/B VSS -1.71fF
C28428 INVX1_LOC_196/Y VSS 0.04fF
C28429 INVX1_LOC_168/Y VSS 0.28fF
C28430 NAND2X1_LOC_253/Y VSS 0.25fF
C28431 NAND2X1_LOC_252/Y VSS 0.27fF
C28432 INVX1_LOC_385/A VSS 0.08fF
C28433 INVX1_LOC_382/Y VSS -0.10fF
C28434 INVX1_LOC_381/Y VSS 0.22fF
C28435 NAND2X1_LOC_397/Y VSS 0.17fF
C28436 INVX1_LOC_363/A VSS 0.12fF
C28437 NAND2X1_LOC_449/B VSS 0.26fF
C28438 INVX1_LOC_345/A VSS 0.08fF
C28439 NAND2X1_LOC_432/Y VSS -0.11fF
C28440 INVX1_LOC_352/A VSS 0.34fF
C28441 NAND2X1_LOC_418/Y VSS 0.24fF
C28442 INVX1_LOC_348/Y VSS 0.32fF
C28443 INVX1_LOC_346/Y VSS 0.40fF
C28444 INVX1_LOC_39/Y VSS -0.01fF
C28445 INVX1_LOC_17/A VSS 0.12fF
C28446 INVX1_LOC_81/A VSS 0.12fF
C28447 INVX1_LOC_82/Y VSS 0.12fF
C28448 INVX1_LOC_498/A VSS -0.09fF
C28449 INVX1_LOC_510/A VSS -2.25fF
C28450 INVX1_LOC_503/Y VSS 0.34fF
C28451 INVX1_LOC_291/Y VSS 0.25fF
C28452 INVX1_LOC_280/A VSS 0.62fF
C28453 INVX1_LOC_469/A VSS 0.12fF
C28454 NAND2X1_LOC_603/Y VSS 0.11fF
C28455 INVX1_LOC_483/Y VSS -0.06fF
C28456 INVX1_LOC_483/A VSS -0.10fF
C28457 INVX1_LOC_472/Y VSS 0.13fF
C28458 INVX1_LOC_494/Y VSS 0.06fF
C28459 INVX1_LOC_338/Y VSS 0.29fF
C28460 INVX1_LOC_649/A VSS 0.24fF
C28461 INVX1_LOC_650/Y VSS 0.06fF
C28462 INVX1_LOC_633/Y VSS 0.29fF
C28463 INVX1_LOC_450/Y VSS 0.04fF
C28464 INVX1_LOC_461/Y VSS 0.04fF
C28465 INVX1_LOC_686/Y VSS 0.04fF
C28466 INVX1_LOC_631/A VSS 0.19fF
C28467 INVX1_LOC_675/Y VSS 0.25fF
C28468 INVX1_LOC_653/Y VSS 0.27fF
C28469 INVX1_LOC_664/Y VSS 0.04fF
C28470 INVX1_LOC_664/A VSS -0.12fF
C28471 INVX1_LOC_620/A VSS 0.18fF
C28472 INVX1_LOC_108/Y VSS -0.06fF
C28473 NAND2X1_LOC_296/Y VSS 0.17fF
C28474 INVX1_LOC_203/A VSS 0.12fF
C28475 INVX1_LOC_224/A VSS -0.17fF
C28476 INVX1_LOC_226/Y VSS 0.06fF
C28477 INVX1_LOC_225/Y VSS 0.25fF
C28478 NAND2X1_LOC_274/Y VSS 0.16fF
C28479 INVX1_LOC_234/Y VSS 0.17fF
C28480 INVX1_LOC_240/A VSS 0.33fF
C28481 INVX1_LOC_189/Y VSS 0.13fF
C28482 INVX1_LOC_388/A VSS 0.42fF
C28483 NAND2X1_LOC_488/Y VSS 0.28fF
C28484 INVX1_LOC_362/A VSS 0.28fF
C28485 INVX1_LOC_383/Y VSS -0.12fF
C28486 INVX1_LOC_375/Y VSS 0.35fF
C28487 INVX1_LOC_325/A VSS 0.12fF
C28488 NAND2X1_LOC_396/Y VSS 0.03fF
C28489 NAND2X1_LOC_395/Y VSS 0.24fF
C28490 INVX1_LOC_351/A VSS 0.32fF
C28491 INVX1_LOC_50/Y VSS -4.03fF
C28492 INVX1_LOC_89/A VSS 0.24fF
C28493 INVX1_LOC_87/A VSS 0.53fF
C28494 INVX1_LOC_290/A VSS 0.15fF
C28495 INVX1_LOC_16/Y VSS 0.06fF
C28496 NAND2X1_LOC_605/B VSS 0.24fF
C28497 INVX1_LOC_497/A VSS 0.20fF
C28498 NAND2X1_LOC_586/Y VSS 0.28fF
C28499 INVX1_LOC_520/A VSS 0.16fF
C28500 INVX1_LOC_509/A VSS 0.26fF
C28501 INVX1_LOC_506/Y VSS -0.40fF
C28502 INVX1_LOC_504/Y VSS 0.27fF
C28503 INVX1_LOC_27/Y VSS 0.22fF
C28504 INVX1_LOC_460/A VSS 0.12fF
C28505 INVX1_LOC_471/Y VSS 0.12fF
C28506 INVX1_LOC_493/Y VSS 0.32fF
C28507 INVX1_LOC_637/A VSS 0.18fF
C28508 NAND2X1_LOC_820/A VSS 0.24fF
C28509 INVX1_LOC_647/Y VSS 0.25fF
C28510 INVX1_LOC_674/Y VSS 0.03fF
C28511 INVX1_LOC_641/Y VSS 0.30fF
C28512 INVX1_LOC_685/Y VSS 0.32fF
C28513 INVX1_LOC_630/A VSS 0.35fF
C28514 INVX1_LOC_652/Y VSS -0.21fF
C28515 INVX1_LOC_663/A VSS 0.12fF
C28516 INVX1_LOC_118/A VSS 0.27fF
C28517 INVX1_LOC_223/A VSS 0.28fF
C28518 INVX1_LOC_247/Y VSS 0.21fF
C28519 INVX1_LOC_239/A VSS -0.08fF
C28520 NAND2X1_LOC_237/Y VSS 0.38fF
C28521 NAND2X1_LOC_231/B VSS 0.24fF
C28522 INVX1_LOC_361/A VSS 0.17fF
C28523 INVX1_LOC_351/Y VSS 0.04fF
C28524 INVX1_LOC_77/Y VSS 0.27fF
C28525 NAND2X1_LOC_448/B VSS 0.19fF
C28526 INVX1_LOC_350/A VSS -0.19fF
C28527 INVX1_LOC_349/Y VSS 0.04fF
C28528 NAND2X1_LOC_496/Y VSS 0.38fF
C28529 INVX1_LOC_74/Y VSS 1.23fF
C28530 INVX1_LOC_376/Y VSS 0.43fF
C28531 INVX1_LOC_372/A VSS 0.14fF
C28532 INVX1_LOC_359/Y VSS 0.25fF
C28533 NAND2X1_LOC_393/Y VSS 0.24fF
C28534 NAND2X1_LOC_410/Y VSS 0.25fF
C28535 INVX1_LOC_48/A VSS 0.05fF
C28536 INVX1_LOC_59/Y VSS 0.29fF
C28537 NAND2X1_LOC_631/B VSS 0.42fF
C28538 NAND2X1_LOC_66/Y VSS 0.23fF
C28539 NAND2X1_LOC_668/Y VSS 0.11fF
C28540 NAND2X1_LOC_615/B VSS 0.16fF
C28541 INVX1_LOC_479/Y VSS -0.14fF
C28542 INVX1_LOC_478/Y VSS 0.18fF
C28543 INVX1_LOC_519/A VSS -0.08fF
C28544 INVX1_LOC_486/Y VSS 0.36fF
C28545 INVX1_LOC_496/A VSS 1.00fF
C28546 INVX1_LOC_481/Y VSS 0.25fF
C28547 INVX1_LOC_492/Y VSS 0.01fF
C28548 INVX1_LOC_660/A VSS -0.08fF
C28549 INVX1_LOC_657/Y VSS 0.31fF
C28550 INVX1_LOC_242/Y VSS 0.45fF
C28551 NAND2X1_LOC_847/A VSS 0.44fF
C28552 INVX1_LOC_646/Y VSS 0.10fF
C28553 NAND2X1_LOC_829/B VSS 0.26fF
C28554 INVX1_LOC_463/Y VSS 0.48fF
C28555 INVX1_LOC_673/Y VSS 0.08fF
C28556 INVX1_LOC_684/A VSS -0.12fF
C28557 INVX1_LOC_651/A VSS 0.13fF
C28558 INVX1_LOC_128/Y VSS -0.11fF
C28559 INVX1_LOC_128/A VSS 0.25fF
C28560 INVX1_LOC_139/Y VSS 0.36fF
C28561 NAND2X1_LOC_786/B VSS 0.33fF
C28562 NAND2X1_LOC_346/B VSS 0.34fF
C28563 NAND2X1_LOC_294/Y VSS -0.84fF
C28564 NAND2X1_LOC_106/B VSS 0.16fF
C28565 NAND2X1_LOC_489/A VSS 0.19fF
C28566 INVX1_LOC_379/Y VSS 0.04fF
C28567 INVX1_LOC_360/A VSS -0.15fF
C28568 INVX1_LOC_352/Y VSS 0.50fF
C28569 NAND2X1_LOC_448/A VSS 0.17fF
C28570 INVX1_LOC_337/Y VSS 0.38fF
C28571 INVX1_LOC_119/Y VSS 0.68fF
C28572 INVX1_LOC_26/Y VSS -2.89fF
C28573 INVX1_LOC_371/A VSS 0.32fF
C28574 INVX1_LOC_25/A VSS -0.12fF
C28575 INVX1_LOC_14/A VSS 0.16fF
C28576 INVX1_LOC_529/Y VSS 0.06fF
C28577 INVX1_LOC_528/Y VSS 0.25fF
C28578 INVX1_LOC_485/Y VSS 0.04fF
C28579 INVX1_LOC_484/Y VSS 0.25fF
C28580 NAND2X1_LOC_728/A VSS 0.16fF
C28581 INVX1_LOC_495/A VSS 0.29fF
C28582 NAND2X1_LOC_428/Y VSS 0.27fF
C28583 INVX1_LOC_468/A VSS 0.38fF
C28584 NAND2X1_LOC_601/Y VSS -0.09fF
C28585 INVX1_LOC_518/A VSS 0.22fF
C28586 INVX1_LOC_659/A VSS -0.72fF
C28587 NAND2X1_LOC_827/Y VSS 0.19fF
C28588 INVX1_LOC_670/A VSS -2.91fF
C28589 INVX1_LOC_480/Y VSS 0.17fF
C28590 INVX1_LOC_491/Y VSS 0.40fF
C28591 INVX1_LOC_635/A VSS 0.11fF
C28592 NAND2X1_LOC_846/B VSS 0.19fF
C28593 INVX1_LOC_58/Y VSS 0.88fF
C28594 INVX1_LOC_661/Y VSS 0.15fF
C28595 INVX1_LOC_149/Y VSS 0.19fF
C28596 INVX1_LOC_138/Y VSS 0.25fF
C28597 INPUT_1 VSS 0.36fF
C28598 INVX1_LOC_116/Y VSS 0.86fF
C28599 INVX1_LOC_116/A VSS 0.17fF
C28600 INVX1_LOC_245/Y VSS -0.14fF
C28601 INVX1_LOC_244/Y VSS 0.12fF
C28602 NAND2X1_LOC_286/A VSS 0.25fF
C28603 INVX1_LOC_199/Y VSS 0.78fF
C28604 NAND2X1_LOC_260/Y VSS 0.21fF
C28605 NAND2X1_LOC_541/B VSS 0.51fF
C28606 INVX1_LOC_319/A VSS 0.47fF
C28607 INVX1_LOC_380/Y VSS 0.32fF
C28608 NAND2X1_LOC_444/A VSS 0.31fF
C28609 INVX1_LOC_370/A VSS 0.24fF
C28610 INVX1_LOC_363/Y VSS 0.12fF
C28611 INVX1_LOC_387/A VSS 0.18fF
C28612 NAND2X1_LOC_844/A VSS 0.57fF
C28613 INVX1_LOC_75/Y VSS 0.30fF
C28614 NAND2X1_LOC_434/B VSS 0.19fF
C28615 INVX1_LOC_359/A VSS 0.09fF
C28616 INVX1_LOC_355/Y VSS 0.14fF
C28617 INVX1_LOC_354/Y VSS 0.25fF
C28618 INVX1_LOC_57/Y VSS 0.10fF
C28619 INVX1_LOC_46/A VSS 0.09fF
C28620 INVX1_LOC_79/Y VSS 0.25fF
C28621 INVX1_LOC_35/A VSS 0.12fF
C28622 NAND2X1_LOC_720/A VSS 0.59fF
C28623 INVX1_LOC_527/Y VSS 0.12fF
C28624 NAND2X1_LOC_679/B VSS 0.26fF
C28625 INVX1_LOC_517/A VSS -0.14fF
C28626 INVX1_LOC_508/Y VSS -0.21fF
C28627 NAND2X1_LOC_691/A VSS 0.19fF
C28628 INVX1_LOC_41/Y VSS 0.94fF
C28629 INVX1_LOC_79/A VSS 0.85fF
C28630 INVX1_LOC_482/Y VSS 0.01fF
C28631 NAND2X1_LOC_615/Y VSS 0.07fF
C28632 NAND2X1_LOC_647/A VSS 0.30fF
C28633 INVX1_LOC_493/A VSS 0.19fF
C28634 INVX1_LOC_13/Y VSS 0.16fF
C28635 INVX1_LOC_15/Y VSS 0.30fF
C28636 NAND2X1_LOC_837/B VSS 0.08fF
C28637 INVX1_LOC_658/A VSS 0.12fF
C28638 INVX1_LOC_667/Y VSS 0.23fF
C28639 NAND2X1_LOC_846/A VSS 0.17fF
C28640 NAND2X1_LOC_814/Y VSS -0.23fF
C28641 INVX1_LOC_6/Y VSS 1.67fF
C28642 INVX1_LOC_669/Y VSS 0.34fF
C28643 INVX1_LOC_634/A VSS 0.12fF
C28644 INVX1_LOC_660/Y VSS 0.24fF
C28645 INVX1_LOC_682/Y VSS 0.43fF
C28646 INVX1_LOC_671/Y VSS 0.40fF
C28647 INVX1_LOC_159/Y VSS 0.16fF
C28648 INVX1_LOC_159/A VSS 0.25fF
C28649 INVX1_LOC_115/Y VSS 0.28fF
C28650 INVX1_LOC_115/A VSS 0.40fF
C28651 INVX1_LOC_104/Y VSS 0.25fF
C28652 INVX1_LOC_126/Y VSS 0.31fF
C28653 INVX1_LOC_126/A VSS 0.22fF
C28654 INVX1_LOC_148/Y VSS 0.34fF
C28655 NAND2X1_LOC_276/A VSS 0.19fF
C28656 INVX1_LOC_221/Y VSS 0.32fF
C28657 NAND2X1_LOC_285/B VSS 0.35fF
C28658 INVX1_LOC_145/Y VSS 0.71fF
C28659 INVX1_LOC_99/Y VSS -4.55fF
C28660 INVX1_LOC_307/A VSS 0.74fF
C28661 INVX1_LOC_318/Y VSS 0.30fF
C28662 INVX1_LOC_329/Y VSS 0.25fF
C28663 INVX1_LOC_328/Y VSS 0.53fF
C28664 INVX1_LOC_369/A VSS 0.35fF
C28665 INVX1_LOC_365/Y VSS 0.12fF
C28666 NAND2X1_LOC_451/B VSS 0.41fF
C28667 NAND2X1_LOC_545/A VSS 0.28fF
C28668 INVX1_LOC_357/Y VSS 0.04fF
C28669 INVX1_LOC_356/Y VSS 0.25fF
C28670 INVX1_LOC_67/Y VSS 0.32fF
C28671 INVX1_LOC_543/A VSS 0.12fF
C28672 INVX1_LOC_484/A VSS 0.26fF
C28673 NAND2X1_LOC_619/Y VSS 0.19fF
C28674 INVX1_LOC_526/Y VSS 0.06fF
C28675 INVX1_LOC_479/A VSS 0.57fF
C28676 INVX1_LOC_491/A VSS -0.29fF
C28677 NAND2X1_LOC_689/B VSS 0.21fF
C28678 INVX1_LOC_539/Y VSS 0.25fF
C28679 INVX1_LOC_516/A VSS 0.21fF
C28680 INVX1_LOC_509/Y VSS 0.25fF
C28681 INVX1_LOC_505/Y VSS -0.56fF
C28682 NAND2X1_LOC_597/Y VSS 0.17fF
C28683 INVX1_LOC_476/A VSS 0.24fF
C28684 INVX1_LOC_477/Y VSS 0.06fF
C28685 NAND2X1_LOC_602/A VSS 0.19fF
C28686 INVX1_LOC_12/A VSS 0.12fF
C28687 INPUT_2 VSS 0.32fF
C28688 INVX1_LOC_657/A VSS 0.19fF
C28689 NAND2X1_LOC_823/Y VSS 0.14fF
C28690 NAND2X1_LOC_837/A VSS 0.23fF
C28691 INVX1_LOC_679/A VSS 0.20fF
C28692 INVX1_LOC_672/Y VSS 0.04fF
C28693 INVX1_LOC_668/A VSS 0.24fF
C28694 NAND2X1_LOC_820/Y VSS 0.13fF
C28695 INVX1_LOC_644/Y VSS 0.06fF
C28696 INVX1_LOC_643/Y VSS 0.07fF
C28697 INVX1_LOC_633/A VSS 0.23fF
C28698 INVX1_LOC_627/Y VSS 0.04fF
C28699 INVX1_LOC_681/Y VSS 0.29fF
C28700 INVX1_LOC_670/Y VSS 0.07fF
C28701 INVX1_LOC_169/A VSS 0.25fF
C28702 INVX1_LOC_125/A VSS 0.21fF
C28703 INVX1_LOC_136/Y VSS 0.18fF
C28704 INVX1_LOC_134/Y VSS -17.39fF
C28705 INVX1_LOC_147/Y VSS 0.26fF
C28706 NAND2X1_LOC_285/A VSS 0.37fF
C28707 INVX1_LOC_232/Y VSS 0.25fF
C28708 INVX1_LOC_339/Y VSS 0.07fF
C28709 INVX1_LOC_317/A VSS 0.32fF
C28710 INVX1_LOC_367/Y VSS 0.26fF
C28711 NAND2X1_LOC_416/Y VSS 0.23fF
C28712 INVX1_LOC_235/Y VSS 0.16fF
C28713 NAND2X1_LOC_833/B VSS 0.25fF
C28714 NAND2X1_LOC_486/A VSS 0.15fF
C28715 INVX1_LOC_357/A VSS 0.30fF
C28716 INVX1_LOC_348/A VSS 0.12fF
C28717 INVX1_LOC_44/Y VSS 0.57fF
C28718 INVX1_LOC_55/A VSS 0.12fF
C28719 INVX1_LOC_88/Y VSS 0.06fF
C28720 INVX1_LOC_77/A VSS 0.12fF
C28721 NAND2X1_LOC_616/Y VSS 0.21fF
C28722 NAND2X1_LOC_719/A VSS 0.17fF
C28723 INVX1_LOC_490/A VSS 0.19fF
C28724 NAND2X1_LOC_612/A VSS -0.05fF
C28725 INVX1_LOC_474/Y VSS 0.22fF
C28726 INVX1_LOC_515/A VSS -0.02fF
C28727 NAND2X1_LOC_679/A VSS 0.37fF
C28728 INVX1_LOC_538/A VSS 0.12fF
C28729 INVX1_LOC_536/Y VSS 0.25fF
C28730 INVX1_LOC_503/A VSS 0.16fF
C28731 NAND2X1_LOC_595/Y VSS 0.39fF
C28732 INVX1_LOC_22/Y VSS 0.25fF
C28733 NAND2X1_LOC_845/B VSS 0.19fF
C28734 INVX1_LOC_223/Y VSS -1.07fF
C28735 INVX1_LOC_642/Y VSS 0.25fF
C28736 NAND2X1_LOC_836/B VSS -0.65fF
C28737 INVX1_LOC_204/Y VSS 0.30fF
C28738 INVX1_LOC_656/A VSS -0.05fF
C28739 NAND2X1_LOC_822/Y VSS 0.13fF
C28740 INVX1_LOC_678/A VSS 0.36fF
C28741 INVX1_LOC_632/A VSS 0.74fF
C28742 INVX1_LOC_680/A VSS 0.10fF
C28743 INVX1_LOC_179/Y VSS 0.41fF
C28744 INVX1_LOC_179/A VSS 0.62fF
C28745 INVX1_LOC_157/Y VSS -0.03fF
C28746 INVX1_LOC_157/A VSS 0.19fF
C28747 INVX1_LOC_124/Y VSS 0.25fF
C28748 INVX1_LOC_135/Y VSS 0.25fF
C28749 INVX1_LOC_62/Y VSS -13.95fF
C28750 INVX1_LOC_102/Y VSS 0.06fF
C28751 INVX1_LOC_100/Y VSS 1.16fF
C28752 NAND2X1_LOC_334/B VSS 0.32fF
C28753 NAND2X1_LOC_542/A VSS -0.48fF
C28754 INVX1_LOC_349/A VSS 0.12fF
C28755 INVX1_LOC_338/A VSS 0.09fF
C28756 INVX1_LOC_305/Y VSS 0.07fF
C28757 INVX1_LOC_378/A VSS 0.30fF
C28758 INVX1_LOC_368/Y VSS 0.14fF
C28759 NAND2X1_LOC_558/B VSS -0.10fF
C28760 NAND2X1_LOC_482/Y VSS 0.41fF
C28761 NAND2X1_LOC_413/Y VSS 0.23fF
C28762 NAND2X1_LOC_411/Y VSS 0.04fF
C28763 INVX1_LOC_356/A VSS 0.23fF
C28764 NAND2X1_LOC_427/Y VSS 0.22fF
C28765 NAND2X1_LOC_426/Y VSS 0.19fF
C28766 INVX1_LOC_519/Y VSS 0.19fF
C28767 INVX1_LOC_508/A VSS 0.24fF
C28768 INVX1_LOC_87/Y VSS 0.25fF
C28769 INVX1_LOC_65/A VSS -0.10fF
C28770 NAND2X1_LOC_755/B VSS 0.33fF
C28771 INVX1_LOC_489/A VSS 0.16fF
C28772 INVX1_LOC_482/A VSS 0.32fF
C28773 NAND2X1_LOC_613/Y VSS 0.07fF
C28774 NAND2X1_LOC_528/Y VSS 0.37fF
C28775 INVX1_LOC_502/A VSS -3.49fF
C28776 INVX1_LOC_405/Y VSS 0.36fF
C28777 INVX1_LOC_533/A VSS 0.13fF
C28778 INVX1_LOC_347/Y VSS 0.39fF
C28779 INVX1_LOC_514/A VSS 0.23fF
C28780 NAND2X1_LOC_594/Y VSS 0.19fF
C28781 INVX1_LOC_537/A VSS -0.90fF
C28782 INVX1_LOC_11/A VSS 0.38fF
C28783 INVX1_LOC_63/Y VSS -4.18fF
C28784 INVX1_LOC_110/A VSS 0.29fF
C28785 INVX1_LOC_677/A VSS 0.12fF
C28786 INVX1_LOC_676/Y VSS 0.24fF
C28787 INVX1_LOC_666/A VSS 0.34fF
C28788 INVX1_LOC_531/Y VSS -2.95fF
C28789 GATE_811 VSS 0.02fF
C28790 INVX1_LOC_640/Y VSS 0.25fF
C28791 NAND2X1_LOC_677/Y VSS 0.24fF
C28792 NAND2X1_LOC_513/A VSS -0.19fF
C28793 INVX1_LOC_630/Y VSS 0.13fF
C28794 INVX1_LOC_178/Y VSS 0.23fF
C28795 INVX1_LOC_145/A VSS 0.18fF
C28796 INVX1_LOC_156/A VSS 0.21fF
C28797 INVX1_LOC_112/Y VSS 0.08fF
C28798 NAND2X1_LOC_334/A VSS 0.72fF
C28799 INVX1_LOC_326/Y VSS 0.40fF
C28800 INVX1_LOC_326/A VSS 0.12fF
C28801 INVX1_LOC_315/A VSS 0.18fF
C28802 INVX1_LOC_304/Y VSS 0.23fF
C28803 INVX1_LOC_304/A VSS 0.20fF
C28804 INVX1_LOC_366/A VSS 0.77fF
C28805 NAND2X1_LOC_409/Y VSS 0.23fF
C28806 INVX1_LOC_390/A VSS 0.27fF
C28807 NAND2X1_LOC_491/Y VSS 0.19fF
C28808 INVX1_LOC_377/A VSS 0.32fF
C28809 INVX1_LOC_371/Y VSS 0.09fF
C28810 INVX1_LOC_518/Y VSS -0.04fF
C28811 INVX1_LOC_507/Y VSS -0.59fF
C28812 INVX1_LOC_507/A VSS 0.08fF
C28813 INVX1_LOC_97/Y VSS 0.19fF
C28814 NAND2X1_LOC_675/B VSS 0.27fF
C28815 INVX1_LOC_532/Y VSS -0.12fF
C28816 NAND2X1_LOC_708/A VSS 0.27fF
C28817 INVX1_LOC_35/Y VSS 1.06fF
C28818 INVX1_LOC_536/A VSS 0.11fF
C28819 INVX1_LOC_20/A VSS 0.12fF
C28820 INVX1_LOC_488/A VSS 0.12fF
C28821 INVX1_LOC_487/Y VSS 0.26fF
C28822 NAND2X1_LOC_628/Y VSS 0.07fF
C28823 INVX1_LOC_501/A VSS -0.30fF
C28824 GATE_662 VSS 0.17fF
C28825 INVX1_LOC_523/Y VSS -0.42fF
C28826 INVX1_LOC_513/A VSS 0.23fF
C28827 INVX1_LOC_460/Y VSS 0.29fF
C28828 INVX1_LOC_42/Y VSS 0.22fF
C28829 INVX1_LOC_9/A VSS 0.12fF
C28830 INVX1_LOC_10/Y VSS 0.25fF
C28831 INVX1_LOC_119/A VSS 0.36fF
C28832 NAND2X1_LOC_123/B VSS 0.32fF
C28833 INVX1_LOC_69/Y VSS 0.85fF
C28834 GATE_865 VSS 0.13fF
C28835 NAND2X1_LOC_829/Y VSS 0.16fF
C28836 INVX1_LOC_654/A VSS 0.36fF
C28837 INVX1_LOC_665/A VSS 0.24fF
C28838 INVX1_LOC_641/A VSS 0.14fF
C28839 INVX1_LOC_638/Y VSS 0.22fF
C28840 INVX1_LOC_637/Y VSS 0.07fF
C28841 INVX1_LOC_177/A VSS 0.19fF
C28842 INVX1_LOC_188/Y VSS -0.51fF
C28843 INVX1_LOC_111/A VSS 0.20fF
C28844 INVX1_LOC_166/Y VSS 0.16fF
C28845 INVX1_LOC_137/Y VSS -1.52fF
C28846 INVX1_LOC_325/Y VSS 0.26fF
C28847 INVX1_LOC_369/Y VSS 0.04fF
C28848 INVX1_LOC_314/Y VSS -0.32fF
C28849 INVX1_LOC_303/Y VSS 0.40fF
C28850 INVX1_LOC_358/Y VSS 0.07fF
C28851 INVX1_LOC_358/A VSS 0.10fF
C28852 INVX1_LOC_336/Y VSS 0.13fF
C28853 NAND2X1_LOC_493/B VSS -0.01fF
C28854 INVX1_LOC_373/Y VSS 0.16fF
C28855 NAND2X1_LOC_555/B VSS 0.33fF
C28856 INVX1_LOC_506/A VSS 0.12fF
C28857 INVX1_LOC_63/A VSS 0.12fF
C28858 INVX1_LOC_96/A VSS 0.32fF
C28859 INVX1_LOC_531/A VSS 0.12fF
C28860 INVX1_LOC_522/Y VSS 0.14fF
C28861 INVX1_LOC_512/A VSS 0.12fF
C28862 INVX1_LOC_499/Y VSS 0.08fF
C28863 INVX1_LOC_500/A VSS 0.17fF
C28864 NAND2X1_LOC_686/B VSS 0.11fF
C28865 INVX1_LOC_49/Y VSS 1.03fF
C28866 NAND2X1_LOC_707/B VSS 0.13fF
C28867 INVX1_LOC_32/Y VSS -4.77fF
C28868 INVX1_LOC_8/Y VSS 0.23fF
C28869 NAND2X1_LOC_123/A VSS 0.37fF
C28870 INVX1_LOC_125/Y VSS 0.33fF
C28871 NAND2X1_LOC_835/A VSS 0.19fF
C28872 INVX1_LOC_640/A VSS 0.12fF
C28873 INVX1_LOC_639/Y VSS 0.13fF
C28874 INVX1_LOC_686/A VSS -4.73fF
C28875 INVX1_LOC_683/Y VSS -0.30fF
C28876 INVX1_LOC_653/A VSS 0.07fF
C28877 NAND2X1_LOC_433/Y VSS 0.37fF
C28878 INVX1_LOC_675/A VSS -1.49fF
C28879 INVX1_LOC_258/Y VSS 0.22fF
C28880 INVX1_LOC_198/Y VSS 0.08fF
C28881 INVX1_LOC_176/A VSS 0.44fF
C28882 INVX1_LOC_154/Y VSS 0.32fF
C28883 INVX1_LOC_187/A VSS 0.18fF
C28884 INVX1_LOC_132/A VSS 0.05fF
C28885 INVX1_LOC_379/A VSS 0.31fF
C28886 INVX1_LOC_324/Y VSS 0.10fF
C28887 INVX1_LOC_324/A VSS 0.19fF
C28888 INVX1_LOC_368/A VSS 0.25fF
C28889 INVX1_LOC_346/A VSS 0.20fF
C28890 INVX1_LOC_608/A VSS 0.29fF
C28891 GATE_479 VSS 0.13fF
C28892 INVX1_LOC_538/Y VSS 0.39fF
C28893 INVX1_LOC_549/Y VSS 0.13fF
C28894 INVX1_LOC_516/Y VSS 0.48fF
C28895 INVX1_LOC_95/A VSS 0.32fF
C28896 NAND2X1_LOC_673/B VSS 0.31fF
C28897 INVX1_LOC_515/Y VSS 0.03fF
C28898 INVX1_LOC_514/Y VSS 0.25fF
C28899 INVX1_LOC_511/A VSS -0.23fF
C28900 NAND2X1_LOC_707/A VSS -0.42fF
C28901 INVX1_LOC_340/Y VSS -0.31fF
C28902 NAND2X1_LOC_686/A VSS 0.24fF
C28903 INVX1_LOC_6/A VSS 0.19fF
C28904 INVX1_LOC_101/Y VSS 0.25fF
C28905 INVX1_LOC_133/A VSS -0.18fF
C28906 INVX1_LOC_132/Y VSS 0.04fF
C28907 INVX1_LOC_131/Y VSS 0.25fF
C28908 NAND2X1_LOC_136/Y VSS 0.41fF
C28909 INVX1_LOC_107/Y VSS 0.17fF
C28910 NAND2X1_LOC_128/B VSS 0.31fF
C28911 INVX1_LOC_674/A VSS 0.63fF
C28912 INVX1_LOC_685/A VSS 0.23fF
C28913 INVX1_LOC_684/Y VSS 0.04fF
C28914 INVX1_LOC_602/Y VSS 0.31fF
C28915 INVX1_LOC_649/Y VSS 0.19fF
C28916 INVX1_LOC_651/Y VSS -0.61fF
C28917 INVX1_LOC_652/A VSS 0.19fF
C28918 NAND2X1_LOC_301/B VSS 0.35fF
C28919 NAND2X1_LOC_274/B VSS 0.86fF
C28920 INVX1_LOC_255/A VSS -0.36fF
C28921 INVX1_LOC_253/Y VSS 0.33fF
C28922 INVX1_LOC_197/A VSS 0.35fF
C28923 INVX1_LOC_153/Y VSS 0.37fF
C28924 INVX1_LOC_120/Y VSS 0.29fF
C28925 INVX1_LOC_186/A VSS 0.21fF
C28926 INVX1_LOC_389/Y VSS 0.25fF
C28927 INVX1_LOC_378/Y VSS 0.25fF
C28928 INVX1_LOC_345/Y VSS 0.19fF
C28929 INVX1_LOC_367/A VSS 0.29fF
C28930 INVX1_LOC_301/Y VSS -0.14fF
C28931 NAND2X1_LOC_557/B VSS 0.32fF
C28932 INVX1_LOC_559/Y VSS 0.41fF
C28933 INVX1_LOC_504/A VSS 0.51fF
C28934 INVX1_LOC_537/Y VSS 0.29fF
C28935 INVX1_LOC_72/Y VSS 0.08fF
C28936 INVX1_LOC_50/A VSS -0.05fF
C28937 INVX1_LOC_94/Y VSS 0.05fF
C28938 INVX1_LOC_61/A VSS 0.10fF
C28939 INVX1_LOC_530/A VSS 0.26fF
C28940 NAND2X1_LOC_685/B VSS 0.12fF
C28941 INVX1_LOC_586/A VSS 1.35fF
C28942 INVX1_LOC_45/Y VSS 1.05fF
C28943 INVX1_LOC_521/A VSS 0.12fF
C28944 INVX1_LOC_517/Y VSS 0.31fF
C28945 NAND2X1_LOC_706/B VSS 0.43fF
C28946 INVX1_LOC_5/Y VSS 0.20fF
C28947 INVX1_LOC_4/Y VSS 0.25fF
C28948 INVX1_LOC_117/A VSS 0.12fF
C28949 INVX1_LOC_100/A VSS 0.19fF
C28950 INVX1_LOC_146/A VSS 0.12fF
C28951 INVX1_LOC_124/A VSS 0.25fF
C28952 NAND2X1_LOC_768/B VSS -0.14fF
C28953 INVX1_LOC_108/A VSS 0.18fF
C28954 INVX1_LOC_105/Y VSS 0.27fF
C28955 INVX1_LOC_673/A VSS 0.16fF
C28956 INVX1_LOC_659/Y VSS 0.10fF
C28957 INVX1_LOC_678/Y VSS 0.04fF
C28958 INVX1_LOC_677/Y VSS -0.21fF
C28959 NAND2X1_LOC_142/Y VSS -0.00fF
C28960 NAND2X1_LOC_108/Y VSS 0.31fF
C28961 INVX1_LOC_662/A VSS -1.60fF
C28962 NAND2X1_LOC_355/A VSS 0.31fF
C28963 INVX1_LOC_261/Y VSS 0.31fF
C28964 INVX1_LOC_254/A VSS 0.18fF
C28965 INVX1_LOC_251/A VSS 0.32fF
C28966 INVX1_LOC_174/A VSS 0.31fF
C28967 INVX1_LOC_196/A VSS 0.12fF
C28968 INVX1_LOC_163/Y VSS 0.10fF
C28969 INVX1_LOC_76/Y VSS -4.23fF
C28970 INVX1_LOC_185/Y VSS 0.26fF
C28971 INVX1_LOC_141/Y VSS 0.12fF
C28972 INVX1_LOC_47/Y VSS -8.20fF
C28973 INVX1_LOC_366/Y VSS 0.04fF
C28974 INVX1_LOC_311/Y VSS 0.06fF
C28975 INVX1_LOC_322/Y VSS -0.23fF
C28976 INVX1_LOC_399/Y VSS -0.24fF
C28977 INVX1_LOC_399/A VSS 0.24fF
C28978 INVX1_LOC_344/Y VSS -0.03fF
C28979 INVX1_LOC_344/A VSS 0.28fF
C28980 INVX1_LOC_377/Y VSS 0.18fF
C28981 INVX1_LOC_355/A VSS 0.30fF
C28982 INVX1_LOC_300/Y VSS 0.39fF
C28983 INVX1_LOC_525/Y VSS 0.57fF
C28984 INVX1_LOC_558/Y VSS 0.14fF
C28985 INVX1_LOC_547/Y VSS 0.29fF
C28986 INVX1_LOC_569/Y VSS -0.22fF
C28987 INVX1_LOC_51/Y VSS -4.89fF
C28988 NAND2X1_LOC_673/A VSS 0.19fF
C28989 NAND2X1_LOC_685/A VSS 0.19fF
C28990 INVX1_LOC_1/A VSS 0.20fF
C28991 INVX1_LOC_2/Y VSS 0.07fF
C28992 INVX1_LOC_154/A VSS 0.11fF
C28993 NAND2X1_LOC_388/A VSS 0.16fF
C28994 NAND2X1_LOC_210/A VSS 0.19fF
C28995 NAND2X1_LOC_156/Y VSS 0.13fF
C28996 INVX1_LOC_131/A VSS 0.15fF
C28997 INVX1_LOC_107/A VSS -0.02fF
C28998 INVX1_LOC_106/Y VSS 0.04fF
C28999 NAND2X1_LOC_128/A VSS 0.50fF
C29000 INVX1_LOC_672/A VSS 0.23fF
C29001 INVX1_LOC_662/Y VSS 0.29fF
C29002 INVX1_LOC_683/A VSS 0.12fF
C29003 INVX1_LOC_680/Y VSS 0.10fF
C29004 INVX1_LOC_679/Y VSS 0.33fF
C29005 INVX1_LOC_661/A VSS -0.05fF
C29006 INVX1_LOC_655/Y VSS 0.33fF
C29007 INVX1_LOC_273/A VSS 0.61fF
C29008 INVX1_LOC_266/Y VSS 0.04fF
C29009 INVX1_LOC_261/A VSS 0.35fF
C29010 INVX1_LOC_262/Y VSS 0.25fF
C29011 NAND2X1_LOC_308/A VSS 0.26fF
C29012 INVX1_LOC_31/Y VSS 0.88fF
C29013 INVX1_LOC_184/A VSS 0.17fF
C29014 INVX1_LOC_173/A VSS 0.26fF
C29015 INVX1_LOC_140/Y VSS 0.42fF
C29016 NAND2X1_LOC_503/Y VSS -0.06fF
C29017 INPUT_7 VSS 0.37fF
C29018 INVX1_LOC_398/A VSS 0.18fF
C29019 INVX1_LOC_321/A VSS 0.19fF
C29020 INVX1_LOC_376/A VSS 0.33fF
C29021 INVX1_LOC_387/Y VSS -0.60fF
C29022 INVX1_LOC_579/Y VSS 0.37fF
C29023 INVX1_LOC_524/Y VSS 0.40fF
C29024 INVX1_LOC_502/Y VSS 0.34fF
C29025 INVX1_LOC_546/A VSS 0.19fF
C29026 INVX1_LOC_557/Y VSS 0.28fF
C29027 INVX1_LOC_513/Y VSS 0.31fF
C29028 INVX1_LOC_568/A VSS 0.12fF
C29029 INVX1_LOC_535/Y VSS 0.14fF
C29030 INVX1_LOC_81/Y VSS 0.19fF
C29031 INVX1_LOC_70/Y VSS 0.25fF
C29032 NAND2X1_LOC_728/B VSS 0.33fF
C29033 INVX1_LOC_542/A VSS 0.20fF
C29034 NAND2X1_LOC_690/Y VSS 0.11fF
C29035 INVX1_LOC_153/A VSS 0.42fF
C29036 NAND2X1_LOC_165/Y VSS 0.28fF
C29037 INVX1_LOC_99/A VSS 0.30fF
C29038 INVX1_LOC_12/Y VSS 0.59fF
C29039 NAND2X1_LOC_122/Y VSS 0.25fF
C29040 NAND2X1_LOC_148/B VSS 0.06fF
C29041 INVX1_LOC_117/Y VSS -8.92fF
C29042 INVX1_LOC_106/A VSS 0.32fF
C29043 NAND2X1_LOC_107/Y VSS 0.31fF
C29044 NAND2X1_LOC_768/A VSS 0.35fF
C29045 NAND2X1_LOC_332/B VSS 0.40fF
C29046 INVX1_LOC_682/A VSS 0.32fF
C29047 INVX1_LOC_671/A VSS -0.06fF
C29048 INVX1_LOC_663/Y VSS 0.09fF
C29049 NAND2X1_LOC_318/B VSS 0.35fF
C29050 INVX1_LOC_268/Y VSS -0.00fF
C29051 INVX1_LOC_259/A VSS 0.11fF
C29052 INVX1_LOC_277/Y VSS 0.04fF
C29053 INVX1_LOC_276/Y VSS 0.22fF
C29054 NAND2X1_LOC_307/B VSS 0.22fF
C29055 INVX1_LOC_89/Y VSS 0.70fF
C29056 INVX1_LOC_172/A VSS -0.49fF
C29057 INVX1_LOC_194/A VSS 0.36fF
C29058 INVX1_LOC_161/A VSS 0.29fF
C29059 INVX1_LOC_396/Y VSS -0.03fF
C29060 NAND2X1_LOC_520/B VSS 0.11fF
C29061 INVX1_LOC_183/Y VSS 0.26fF
C29062 INVX1_LOC_183/A VSS -0.11fF
C29063 INVX1_LOC_397/Y VSS 0.21fF
C29064 INVX1_LOC_342/Y VSS 0.17fF
C29065 INVX1_LOC_320/A VSS 0.38fF
C29066 INVX1_LOC_353/Y VSS 0.08fF
C29067 INVX1_LOC_364/Y VSS 0.37fF
C29068 INVX1_LOC_375/A VSS 0.27fF
C29069 INVX1_LOC_386/A VSS 0.35fF
C29070 INVX1_LOC_331/Y VSS 0.25fF
C29071 INVX1_LOC_589/Y VSS 0.23fF
C29072 INVX1_LOC_578/Y VSS 0.17fF
C29073 INVX1_LOC_556/Y VSS -0.63fF
C29074 INVX1_LOC_567/Y VSS 0.43fF
C29075 INVX1_LOC_545/Y VSS 0.20fF
C29076 INVX1_LOC_501/Y VSS 0.14fF
C29077 INVX1_LOC_512/Y VSS -0.06fF
C29078 INVX1_LOC_523/A VSS 0.47fF
C29079 INVX1_LOC_534/Y VSS 0.39fF
C29080 INVX1_LOC_541/Y VSS 0.25fF
C29081 INVX1_LOC_98/A VSS 0.43fF
C29082 INVX1_LOC_96/Y VSS 0.25fF
C29083 INVX1_LOC_105/A VSS 0.35fF
C29084 NAND2X1_LOC_775/B VSS 0.29fF
C29085 NAND2X1_LOC_148/A VSS 0.44fF
C29086 INVX1_LOC_80/A VSS 0.83fF
C29087 INVX1_LOC_142/Y VSS 0.04fF
C29088 NAND2X1_LOC_192/A VSS 0.32fF
C29089 NAND2X1_LOC_181/A VSS 0.42fF
C29090 INVX1_LOC_681/A VSS 0.35fF
C29091 INVX1_LOC_321/Y VSS 0.18fF
C29092 NAND2X1_LOC_307/A VSS -0.18fF
C29093 NAND2X1_LOC_318/A VSS 0.15fF
C29094 INVX1_LOC_271/A VSS 0.53fF
C29095 INVX1_LOC_293/A VSS 0.29fF
C29096 INVX1_LOC_283/Y VSS 0.10fF
C29097 INVX1_LOC_282/A VSS 0.32fF
C29098 INVX1_LOC_278/Y VSS 0.25fF
C29099 INVX1_LOC_258/A VSS 0.12fF
C29100 INVX1_LOC_256/Y VSS 0.25fF
C29101 INVX1_LOC_171/A VSS 0.16fF
C29102 INVX1_LOC_160/A VSS 0.43fF
C29103 INVX1_LOC_397/A VSS 0.35fF
C29104 NAND2X1_LOC_505/Y VSS 0.27fF
C29105 NAND2X1_LOC_520/A VSS 0.11fF
C29106 INVX1_LOC_396/A VSS 0.19fF
C29107 INVX1_LOC_385/Y VSS 0.28fF
C29108 INVX1_LOC_374/A VSS -0.16fF
C29109 INPUT_5 VSS 0.08fF
C29110 INVX1_LOC_335/A VSS 0.43fF
C29111 INVX1_LOC_330/A VSS 0.29fF
C29112 INVX1_LOC_599/Y VSS 0.18fF
C29113 INVX1_LOC_599/A VSS 0.12fF
C29114 INVX1_LOC_566/Y VSS 0.17fF
C29115 INVX1_LOC_566/A VSS 0.56fF
C29116 INVX1_LOC_577/Y VSS 0.46fF
C29117 INVX1_LOC_533/Y VSS 0.27fF
C29118 INVX1_LOC_544/Y VSS 0.30fF
C29119 INVX1_LOC_555/A VSS 0.84fF
C29120 INVX1_LOC_522/A VSS 0.08fF
C29121 INVX1_LOC_500/Y VSS 0.21fF
C29122 INVX1_LOC_511/Y VSS 0.16fF
C29123 INVX1_LOC_90/A VSS -0.05fF
C29124 INVX1_LOC_175/A VSS 0.13fF
C29125 INVX1_LOC_172/Y VSS 0.04fF
C29126 INVX1_LOC_171/Y VSS 0.20fF
C29127 NAND2X1_LOC_498/B VSS 0.31fF
C29128 INVX1_LOC_165/Y VSS 0.12fF
C29129 INVX1_LOC_97/A VSS -0.15fF
C29130 INVX1_LOC_123/A VSS 0.29fF
C29131 NAND2X1_LOC_169/A VSS 0.09fF
C29132 NAND2X1_LOC_180/B VSS 0.55fF
C29133 NAND2X1_LOC_121/Y VSS 0.17fF
C29134 INVX1_LOC_103/Y VSS -0.04fF
C29135 NAND2X1_LOC_147/B VSS 0.42fF
C29136 INVX1_LOC_142/A VSS 0.35fF
C29137 INVX1_LOC_144/Y VSS 0.06fF
C29138 INVX1_LOC_143/Y VSS 0.25fF
C29139 INVX1_LOC_292/A VSS 0.09fF
C29140 INVX1_LOC_285/Y VSS 0.04fF
C29141 INVX1_LOC_281/A VSS 0.19fF
C29142 INVX1_LOC_280/Y VSS 0.18fF
C29143 NAND2X1_LOC_297/Y VSS 0.19fF
C29144 INVX1_LOC_270/A VSS 0.68fF
C29145 INVX1_LOC_250/A VSS 0.19fF
C29146 INVX1_LOC_249/Y VSS 0.15fF
C29147 NAND2X1_LOC_317/B VSS 0.20fF
C29148 INVX1_LOC_257/A VSS 0.18fF
C29149 INVX1_LOC_412/A VSS -0.12fF
C29150 INVX1_LOC_410/Y VSS 0.57fF
C29151 INVX1_LOC_170/Y VSS 0.17fF
C29152 INVX1_LOC_170/A VSS 0.32fF
C29153 INVX1_LOC_395/Y VSS 0.06fF
C29154 INVX1_LOC_384/Y VSS -0.03fF
C29155 INVX1_LOC_384/A VSS 0.85fF
C29156 INVX1_LOC_362/Y VSS 0.46fF
C29157 INVX1_LOC_373/A VSS 0.17fF
C29158 INVX1_LOC_551/A VSS 0.20fF
C29159 NAND2X1_LOC_698/Y VSS 0.19fF
C29160 INVX1_LOC_598/A VSS 0.34fF
C29161 INVX1_LOC_565/A VSS 0.23fF
C29162 INVX1_LOC_510/Y VSS 0.47fF
C29163 INVX1_LOC_521/Y VSS 0.18fF
C29164 INVX1_LOC_554/Y VSS 0.10fF
C29165 INVX1_LOC_173/Y VSS -0.05fF
C29166 INVX1_LOC_139/A VSS -0.12fF
C29167 INVX1_LOC_129/A VSS 0.12fF
C29168 INVX1_LOC_130/Y VSS 0.11fF
C29169 INVX1_LOC_526/A VSS -0.04fF
C29170 INVX1_LOC_114/Y VSS -0.01fF
C29171 INVX1_LOC_103/A VSS 0.12fF
C29172 NAND2X1_LOC_137/A VSS 0.27fF
C29173 INVX1_LOC_93/Y VSS 0.90fF
C29174 INVX1_LOC_310/Y VSS 0.16fF
C29175 INVX1_LOC_291/A VSS 0.68fF
C29176 INVX1_LOC_287/Y VSS 0.26fF
C29177 INVX1_LOC_286/Y VSS 0.21fF
C29178 INVX1_LOC_269/A VSS 0.52fF
C29179 NAND2X1_LOC_370/A VSS 0.45fF
C29180 NAND2X1_LOC_457/A VSS 0.20fF
C29181 NAND2X1_LOC_271/B VSS 0.40fF
C29182 NAND2X1_LOC_292/Y VSS 0.11fF
C29183 INVX1_LOC_256/A VSS 0.12fF
C29184 NAND2X1_LOC_320/Y VSS 0.28fF
C29185 INVX1_LOC_249/A VSS 0.27fF
C29186 NAND2X1_LOC_299/Y VSS -0.15fF
C29187 INVX1_LOC_191/A VSS 0.21fF
C29188 INVX1_LOC_180/A VSS 0.12fF
C29189 INVX1_LOC_422/Y VSS -0.02fF
C29190 NAND2X1_LOC_531/Y VSS 0.05fF
C29191 INVX1_LOC_411/A VSS 0.27fF
C29192 NAND2X1_LOC_513/Y VSS 0.38fF
C29193 INVX1_LOC_361/Y VSS 0.37fF
C29194 INVX1_LOC_372/Y VSS -0.10fF
C29195 INVX1_LOC_383/A VSS 0.12fF
C29196 INVX1_LOC_562/A VSS 0.34fF
C29197 NAND2X1_LOC_666/Y VSS 0.17fF
C29198 INVX1_LOC_550/A VSS 0.26fF
C29199 INVX1_LOC_597/A VSS 0.18fF
C29200 INVX1_LOC_586/Y VSS 0.25fF
C29201 INVX1_LOC_564/Y VSS -0.04fF
C29202 INVX1_LOC_553/Y VSS 0.17fF
C29203 INVX1_LOC_553/A VSS 0.12fF
C29204 INVX1_LOC_520/Y VSS 0.02fF
C29205 INVX1_LOC_542/Y VSS 0.18fF
C29206 INVX1_LOC_575/Y VSS 0.37fF
C29207 NAND2X1_LOC_56/Y VSS 0.16fF
C29208 INVX1_LOC_156/Y VSS 0.04fF
C29209 NAND2X1_LOC_173/Y VSS 0.44fF
C29210 INVX1_LOC_137/A VSS 0.08fF
C29211 INVX1_LOC_164/Y VSS 0.07fF
C29212 NAND2X1_LOC_140/B VSS 0.36fF
C29213 NAND2X1_LOC_130/Y VSS 0.07fF
C29214 INVX1_LOC_113/Y VSS 0.06fF
C29215 INVX1_LOC_307/Y VSS 0.04fF
C29216 INVX1_LOC_309/Y VSS 0.12fF
C29217 INVX1_LOC_318/A VSS 0.30fF
C29218 NAND2X1_LOC_387/Y VSS 0.40fF
C29219 GATE_366 VSS 0.05fF
C29220 INVX1_LOC_299/Y VSS 0.10fF
C29221 INVX1_LOC_248/A VSS 0.12fF
C29222 NAND2X1_LOC_325/B VSS -0.49fF
C29223 NAND2X1_LOC_261/Y VSS 0.23fF
C29224 INVX1_LOC_220/Y VSS 0.49fF
C29225 INVX1_LOC_289/Y VSS 0.04fF
C29226 INVX1_LOC_190/Y VSS 0.28fF
C29227 INVX1_LOC_410/A VSS 0.33fF
C29228 NAND2X1_LOC_507/A VSS 0.05fF
C29229 NAND2X1_LOC_529/Y VSS 0.17fF
C29230 NAND2X1_LOC_517/Y VSS 0.29fF
C29231 NAND2X1_LOC_516/B VSS 0.22fF
C29232 NAND2X1_LOC_704/B VSS 0.14fF
C29233 INVX1_LOC_572/A VSS 0.12fF
C29234 INVX1_LOC_382/A VSS 0.18fF
C29235 INVX1_LOC_360/Y VSS 0.37fF
C29236 INVX1_LOC_549/A VSS 0.32fF
C29237 INVX1_LOC_561/A VSS 0.10fF
C29238 INVX1_LOC_469/Y VSS 0.27fF
C29239 NAND2X1_LOC_591/Y VSS 0.34fF
C29240 INVX1_LOC_596/A VSS 0.39fF
C29241 INVX1_LOC_530/Y VSS 0.50fF
C29242 INVX1_LOC_552/Y VSS 0.11fF
C29243 INVX1_LOC_53/Y VSS -3.50fF
C29244 NAND2X1_LOC_467/A VSS 0.12fF
C29245 INVX1_LOC_162/Y VSS 0.25fF
C29246 INVX1_LOC_122/Y VSS 0.06fF
C29247 INVX1_LOC_121/Y VSS 0.35fF
C29248 INVX1_LOC_127/Y VSS -0.15fF
C29249 NAND2X1_LOC_403/A VSS -0.18fF
C29250 INVX1_LOC_308/Y VSS 0.06fF
C29251 INVX1_LOC_267/A VSS 0.12fF
C29252 INVX1_LOC_300/A VSS 0.59fF
C29253 INVX1_LOC_296/Y VSS 0.12fF
C29254 NAND2X1_LOC_538/B VSS 0.20fF
C29255 INVX1_LOC_278/A VSS 0.34fF
C29256 INVX1_LOC_217/Y VSS 0.24fF
C29257 INVX1_LOC_289/A VSS 0.21fF
C29258 NAND2X1_LOC_331/Y VSS 0.17fF
C29259 INVX1_LOC_421/A VSS 0.43fF
C29260 NAND2X1_LOC_527/Y VSS 0.27fF
C29261 NAND2X1_LOC_537/B VSS 0.15fF
C29262 INVX1_LOC_403/Y VSS 0.25fF
C29263 INVX1_LOC_381/A VSS 0.36fF
C29264 INVX1_LOC_392/Y VSS 0.15fF
C29265 INVX1_LOC_560/A VSS -1.22fF
C29266 INVX1_LOC_390/Y VSS 0.34fF
C29267 INVX1_LOC_582/A VSS 0.30fF
C29268 INVX1_LOC_573/Y VSS 0.29fF
C29269 INVX1_LOC_571/A VSS 0.12fF
C29270 INVX1_LOC_548/A VSS 0.82fF
C29271 NAND2X1_LOC_692/Y VSS 0.17fF
C29272 INVX1_LOC_370/Y VSS 0.41fF
C29273 INVX1_LOC_595/A VSS 0.12fF
C29274 INVX1_LOC_551/Y VSS 0.29fF
C29275 INVX1_LOC_584/Y VSS -0.15fF
C29276 INVX1_LOC_540/Y VSS -0.01fF
C29277 NAND2X1_LOC_43/Y VSS 0.16fF
C29278 NAND2X1_LOC_41/Y VSS 0.23fF
C29279 NAND2X1_LOC_152/B VSS 0.07fF
C29280 NAND2X1_LOC_163/B VSS 0.13fF
C29281 INVX1_LOC_150/Y VSS 0.19fF
C29282 INVX1_LOC_127/A VSS 0.13fF
C29283 INVX1_LOC_118/Y VSS 0.23fF
C29284 INVX1_LOC_209/A VSS 0.22fF
C29285 NAND2X1_LOC_399/B VSS 0.28fF
C29286 INVX1_LOC_323/Y VSS 0.13fF
C29287 INVX1_LOC_315/Y VSS 0.04fF
C29288 INVX1_LOC_299/A VSS 0.12fF
C29289 INVX1_LOC_290/Y VSS 0.52fF
C29290 NAND2X1_LOC_335/B VSS 0.07fF
C29291 INVX1_LOC_277/A VSS 0.27fF
C29292 NAND2X1_LOC_843/A VSS 0.29fF
C29293 NAND2X1_LOC_250/Y VSS 0.07fF
C29294 NAND2X1_LOC_324/B VSS 0.06fF
C29295 INVX1_LOC_288/A VSS -0.52fF
C29296 INVX1_LOC_255/Y VSS 0.28fF
C29297 NAND2X1_LOC_111/Y VSS 0.67fF
C29298 INVX1_LOC_431/A VSS 0.29fF
C29299 NAND2X1_LOC_545/B VSS 0.22fF
C29300 INVX1_LOC_442/A VSS 0.80fF
C29301 INVX1_LOC_441/Y VSS 0.04fF
C29302 INVX1_LOC_453/A VSS 0.12fF
C29303 INVX1_LOC_449/Y VSS 0.17fF
C29304 INVX1_LOC_401/Y VSS 0.35fF
C29305 NAND2X1_LOC_526/Y VSS 0.27fF
C29306 NAND2X1_LOC_525/Y VSS 0.20fF
C29307 INVX1_LOC_409/A VSS 0.21fF
C29308 NAND2X1_LOC_534/Y VSS 0.07fF
C29309 NAND2X1_LOC_788/A VSS 0.60fF
C29310 NAND2X1_LOC_503/B VSS 0.28fF
C29311 INVX1_LOC_394/Y VSS 0.25fF
C29312 INVX1_LOC_380/A VSS -0.02fF
C29313 INVX1_LOC_391/A VSS 0.19fF
C29314 INVX1_LOC_585/Y VSS 0.25fF
C29315 INVX1_LOC_559/A VSS 0.12fF
C29316 INVX1_LOC_248/Y VSS -0.32fF
C29317 INVX1_LOC_581/A VSS -1.71fF
C29318 INVX1_LOC_574/Y VSS 0.25fF
C29319 INVX1_LOC_547/A VSS 0.37fF
C29320 NAND2X1_LOC_486/B VSS -0.02fF
C29321 INVX1_LOC_570/A VSS -0.15fF
C29322 INVX1_LOC_561/Y VSS 0.15fF
C29323 INVX1_LOC_594/Y VSS 0.25fF
C29324 INVX1_LOC_572/Y VSS 0.36fF
C29325 INVX1_LOC_550/Y VSS 0.04fF
C29326 INVX1_LOC_583/A VSS 0.35fF
C29327 NAND2X1_LOC_16/Y VSS -0.06fF
C29328 NAND2X1_LOC_174/B VSS 0.25fF
C29329 INVX1_LOC_27/A VSS 0.21fF
C29330 INVX1_LOC_28/Y VSS 0.09fF
C29331 INVX1_LOC_134/A VSS 0.18fF
C29332 INVX1_LOC_65/Y VSS 0.47fF
C29333 INVX1_LOC_150/A VSS 0.31fF
C29334 INVX1_LOC_152/Y VSS 0.06fF
C29335 INVX1_LOC_151/Y VSS 0.25fF
C29336 INVX1_LOC_208/Y VSS 0.21fF
C29337 INVX1_LOC_208/A VSS 0.16fF
C29338 INVX1_LOC_219/Y VSS 0.36fF
C29339 NAND2X1_LOC_376/B VSS 0.15fF
C29340 INVX1_LOC_306/Y VSS 0.06fF
C29341 INVX1_LOC_298/A VSS -0.89fF
C29342 INVX1_LOC_25/Y VSS 0.22fF
C29343 INVX1_LOC_316/Y VSS 0.37fF
C29344 INVX1_LOC_250/Y VSS 0.12fF
C29345 INVX1_LOC_419/A VSS 0.12fF
C29346 INVX1_LOC_452/A VSS -0.25fF
C29347 INVX1_LOC_442/Y VSS -1.87fF
C29348 INVX1_LOC_401/A VSS 0.26fF
C29349 NAND2X1_LOC_592/B VSS 0.11fF
C29350 INVX1_LOC_406/A VSS 0.18fF
C29351 NAND2X1_LOC_521/Y VSS 0.34fF
C29352 INVX1_LOC_386/Y VSS 0.35fF
C29353 INVX1_LOC_393/A VSS 0.12fF
C29354 NAND2X1_LOC_498/Y VSS 0.32fF
C29355 INVX1_LOC_412/Y VSS 0.48fF
C29356 NAND2X1_LOC_789/A VSS 0.13fF
C29357 INVX1_LOC_543/Y VSS 0.17fF
C29358 INVX1_LOC_576/Y VSS 0.25fF
C29359 INVX1_LOC_569/A VSS 0.29fF
C29360 NAND2X1_LOC_152/Y VSS 0.16fF
C29361 INVX1_LOC_558/A VSS 0.69fF
C29362 NAND2X1_LOC_317/A VSS 0.11fF
C29363 INVX1_LOC_560/Y VSS 0.42fF
C29364 INVX1_LOC_593/Y VSS 0.38fF
C29365 INVX1_LOC_38/A VSS 0.15fF
C29366 INVX1_LOC_26/A VSS 0.12fF
C29367 NAND2X1_LOC_333/A VSS 0.53fF
C29368 INVX1_LOC_158/Y VSS 0.07fF
C29369 INVX1_LOC_147/A VSS 0.17fF
C29370 INVX1_LOC_229/Y VSS 0.03fF
C29371 INVX1_LOC_218/A VSS 0.16fF
C29372 INVX1_LOC_207/A VSS 0.24fF
C29373 NAND2X1_LOC_537/A VSS 0.43fF
C29374 INVX1_LOC_202/Y VSS 0.29fF
C29375 INVX1_LOC_297/A VSS 0.07fF
C29376 INVX1_LOC_294/Y VSS 0.31fF
C29377 INVX1_LOC_293/Y VSS 0.71fF
C29378 INVX1_LOC_286/A VSS 0.18fF
C29379 INVX1_LOC_271/Y VSS 0.04fF
C29380 INVX1_LOC_160/Y VSS 0.48fF
C29381 NAND2X1_LOC_331/B VSS 0.24fF
C29382 INVX1_LOC_265/Y VSS 0.06fF
C29383 INVX1_LOC_264/Y VSS 0.25fF
C29384 NAND2X1_LOC_373/Y VSS 0.14fF
C29385 NAND2X1_LOC_322/Y VSS 0.31fF
C29386 INVX1_LOC_466/A VSS 0.13fF
C29387 INVX1_LOC_467/Y VSS 0.10fF
C29388 INVX1_LOC_451/A VSS 0.64fF
C29389 INVX1_LOC_444/Y VSS 0.26fF
C29390 NAND2X1_LOC_638/A VSS 0.39fF
C29391 INVX1_LOC_455/Y VSS 0.33fF
C29392 INVX1_LOC_429/A VSS 0.09fF
C29393 NAND2X1_LOC_532/Y VSS 0.25fF
C29394 INVX1_LOC_392/A VSS 0.49fF
C29395 INVX1_LOC_391/Y VSS 0.13fF
C29396 NAND2X1_LOC_523/B VSS 0.22fF
C29397 INVX1_LOC_418/A VSS 0.52fF
C29398 NAND2X1_LOC_764/Y VSS 0.11fF
C29399 NAND2X1_LOC_763/Y VSS 0.19fF
C29400 NAND2X1_LOC_759/B VSS 0.10fF
C29401 INVX1_LOC_592/Y VSS 0.16fF
C29402 NAND2X1_LOC_782/A VSS 0.08fF
C29403 INVX1_LOC_54/Y VSS 0.91fF
C29404 INVX1_LOC_545/A VSS 0.23fF
C29405 INVX1_LOC_579/A VSS 0.27fF
C29406 INVX1_LOC_555/Y VSS 0.25fF
C29407 INVX1_LOC_557/A VSS 0.11fF
C29408 INVX1_LOC_546/Y VSS 0.04fF
C29409 INVX1_LOC_570/Y VSS 0.22fF
C29410 INVX1_LOC_581/Y VSS 0.25fF
C29411 NAND2X1_LOC_39/Y VSS 0.25fF
C29412 INVX1_LOC_36/A VSS 0.12fF
C29413 INVX1_LOC_37/Y VSS 0.25fF
C29414 INVX1_LOC_155/A VSS 0.12fF
C29415 NAND2X1_LOC_179/Y VSS -0.10fF
C29416 INVX1_LOC_168/A VSS 0.12fF
C29417 INVX1_LOC_167/Y VSS -0.23fF
C29418 INVX1_LOC_228/Y VSS 0.01fF
C29419 INVX1_LOC_217/A VSS -0.04fF
C29420 INVX1_LOC_239/Y VSS 0.32fF
C29421 INVX1_LOC_274/A VSS 0.50fF
C29422 INVX1_LOC_285/A VSS 0.29fF
C29423 INVX1_LOC_272/Y VSS 0.04fF
C29424 NAND2X1_LOC_391/B VSS 0.21fF
C29425 NAND2X1_LOC_383/Y VSS 0.38fF
C29426 INVX1_LOC_409/Y VSS -0.01fF
C29427 INVX1_LOC_455/A VSS 0.27fF
C29428 INVX1_LOC_456/Y VSS 0.25fF
C29429 INVX1_LOC_439/A VSS 0.12fF
C29430 INVX1_LOC_424/Y VSS 0.21fF
C29431 INVX1_LOC_450/A VSS 0.29fF
C29432 INVX1_LOC_446/Y VSS -3.14fF
C29433 INVX1_LOC_445/Y VSS 0.42fF
C29434 INVX1_LOC_463/A VSS 0.10fF
C29435 INVX1_LOC_465/Y VSS 0.24fF
C29436 INVX1_LOC_400/A VSS 0.32fF
C29437 INVX1_LOC_398/Y VSS 0.25fF
C29438 INVX1_LOC_408/Y VSS 0.21fF
C29439 NAND2X1_LOC_106/Y VSS 0.23fF
C29440 NAND2X1_LOC_791/B VSS 0.34fF
C29441 NAND2X1_LOC_756/Y VSS -0.83fF
C29442 INVX1_LOC_578/A VSS 1.07fF
C29443 INVX1_LOC_490/Y VSS 0.40fF
C29444 INVX1_LOC_393/Y VSS -0.01fF
C29445 NAND2X1_LOC_781/B VSS 0.33fF
C29446 INVX1_LOC_609/A VSS 0.25fF
C29447 NAND2X1_LOC_697/Y VSS 0.43fF
C29448 INVX1_LOC_556/A VSS -0.11fF
C29449 INVX1_LOC_548/Y VSS 0.04fF
C29450 INVX1_LOC_567/A VSS 0.10fF
C29451 INVX1_LOC_544/A VSS 0.34fF
C29452 INVX1_LOC_591/Y VSS 0.25fF
C29453 INVX1_LOC_580/Y VSS 0.23fF
C29454 INVX1_LOC_580/A VSS 0.12fF
C29455 INVX1_LOC_54/A VSS -0.09fF
C29456 INVX1_LOC_47/A VSS 0.12fF
C29457 INVX1_LOC_158/A VSS 0.12fF
C29458 NAND2X1_LOC_176/Y VSS 0.21fF
C29459 INVX1_LOC_167/A VSS 0.20fF
C29460 NAND2X1_LOC_187/Y VSS 0.16fF
C29461 INVX1_LOC_205/Y VSS 0.39fF
C29462 INVX1_LOC_238/Y VSS 0.13fF
C29463 INVX1_LOC_238/A VSS 0.02fF
C29464 NAND2X1_LOC_400/B VSS 0.21fF
C29465 INVX1_LOC_313/Y VSS 0.25fF
C29466 INVX1_LOC_284/A VSS 0.20fF
C29467 INVX1_LOC_275/Y VSS 0.29fF
C29468 INVX1_LOC_295/A VSS 0.29fF
C29469 INVX1_LOC_425/Y VSS 0.25fF
C29470 NAND2X1_LOC_336/B VSS -0.40fF
C29471 INVX1_LOC_427/A VSS 0.00fF
C29472 INVX1_LOC_413/Y VSS -0.49fF
C29473 NAND2X1_LOC_596/Y VSS 0.32fF
C29474 INVX1_LOC_448/Y VSS 0.04fF
C29475 INVX1_LOC_619/A VSS -5.93fF
C29476 NAND2X1_LOC_773/A VSS 0.19fF
C29477 NAND2X1_LOC_79/B VSS 0.11fF
C29478 INVX1_LOC_590/Y VSS 0.06fF
C29479 INVX1_LOC_577/A VSS 0.41fF
C29480 NAND2X1_LOC_475/A VSS -0.99fF
C29481 NAND2X1_LOC_781/A VSS 0.19fF
C29482 INVX1_LOC_607/A VSS 0.38fF
C29483 NAND2X1_LOC_710/B VSS 0.29fF
C29484 INVX1_LOC_206/Y VSS 1.02fF
C29485 INVX1_LOC_166/A VSS -3.93fF
C29486 NAND2X1_LOC_184/Y VSS -0.69fF
C29487 NAND2X1_LOC_48/Y VSS -0.08fF
C29488 INVX1_LOC_33/Y VSS 0.33fF
C29489 INVX1_LOC_24/A VSS 0.12fF
C29490 INVX1_LOC_237/Y VSS 0.13fF
C29491 INVX1_LOC_294/A VSS 0.12fF
C29492 INVX1_LOC_211/Y VSS 0.18fF
C29493 NAND2X1_LOC_391/A VSS 0.32fF
C29494 INVX1_LOC_312/Y VSS 0.31fF
C29495 INVX1_LOC_84/A VSS 0.55fF
C29496 INVX1_LOC_302/A VSS 0.12fF
C29497 INVX1_LOC_407/Y VSS 0.26fF
C29498 NAND2X1_LOC_548/B VSS 0.32fF
C29499 INVX1_LOC_416/Y VSS 0.14fF
C29500 NAND2X1_LOC_637/A VSS 0.26fF
C29501 INVX1_LOC_437/A VSS 0.20fF
C29502 INVX1_LOC_428/Y VSS 0.21fF
C29503 INVX1_LOC_427/Y VSS 0.10fF
C29504 NAND2X1_LOC_516/Y VSS 0.15fF
C29505 INVX1_LOC_400/Y VSS -0.15fF
C29506 INVX1_LOC_414/A VSS 0.26fF
C29507 NAND2X1_LOC_770/B VSS 0.11fF
C29508 NAND2X1_LOC_791/A VSS 0.19fF
C29509 INVX1_LOC_576/A VSS -0.05fF
C29510 INVX1_LOC_565/Y VSS 0.12fF
C29511 INVX1_LOC_562/Y VSS 0.04fF
C29512 INVX1_LOC_605/A VSS 0.12fF
C29513 INVX1_LOC_606/Y VSS 0.25fF
C29514 NAND2X1_LOC_780/B VSS 0.12fF
C29515 INVX1_LOC_554/A VSS -0.11fF
C29516 INVX1_LOC_468/Y VSS 0.47fF
C29517 NAND2X1_LOC_710/A VSS 0.25fF
C29518 NAND2X1_LOC_61/A VSS 0.19fF
C29519 INVX1_LOC_53/A VSS 0.31fF
C29520 INVX1_LOC_45/A VSS 0.18fF
C29521 INVX1_LOC_269/Y VSS 0.15fF
C29522 INVX1_LOC_492/A VSS 0.35fF
C29523 INVX1_LOC_236/A VSS 0.12fF
C29524 INVX1_LOC_21/A VSS 0.12fF
C29525 INVX1_LOC_23/Y VSS 0.03fF
C29526 INVX1_LOC_33/A VSS 0.16fF
C29527 INVX1_LOC_34/Y VSS 0.30fF
C29528 INVX1_LOC_203/Y VSS 0.30fF
C29529 INVX1_LOC_214/Y VSS 0.33fF
C29530 INVX1_LOC_17/Y VSS 1.15fF
C29531 INVX1_LOC_312/A VSS 0.30fF
C29532 INPUT_3 VSS 0.54fF
C29533 INVX1_LOC_320/Y VSS 0.04fF
C29534 INVX1_LOC_319/Y VSS 0.10fF
C29535 INVX1_LOC_301/A VSS 0.46fF
C29536 NAND2X1_LOC_543/B VSS 0.22fF
C29537 INVX1_LOC_439/Y VSS -5.62fF
C29538 INVX1_LOC_417/Y VSS 0.08fF
C29539 INVX1_LOC_417/A VSS 0.12fF
C29540 INVX1_LOC_406/Y VSS 0.35fF
C29541 INVX1_LOC_428/A VSS 0.13fF
C29542 INVX1_LOC_447/A VSS 0.29fF
C29543 INVX1_LOC_419/Y VSS 0.44fF
C29544 INVX1_LOC_418/Y VSS 0.44fF
C29545 NAND2X1_LOC_636/B VSS 0.28fF
C29546 INVX1_LOC_429/Y VSS 0.11fF
C29547 NAND2X1_LOC_249/Y VSS 0.14fF
C29548 INVX1_LOC_413/A VSS 0.29fF
C29549 NAND2X1_LOC_190/A VSS 0.31fF
C29550 INVX1_LOC_609/Y VSS 0.25fF
C29551 INVX1_LOC_604/A VSS -0.14fF
C29552 NAND2X1_LOC_241/B VSS 0.27fF
C29553 NAND2X1_LOC_164/Y VSS 0.25fF
C29554 NAND2X1_LOC_770/A VSS 0.23fF
C29555 INVX1_LOC_564/A VSS 0.26fF
C29556 INVX1_LOC_563/Y VSS 0.20fF
C29557 NAND2X1_LOC_790/B VSS 0.28fF
C29558 INVX1_LOC_575/A VSS 0.17fF
C29559 INVX1_LOC_568/Y VSS 0.04fF
C29560 NAND2X1_LOC_780/A VSS 0.11fF
C29561 INVX1_LOC_185/A VSS 0.19fF
C29562 INVX1_LOC_133/Y VSS 0.46fF
C29563 INVX1_LOC_44/A VSS 0.25fF
C29564 INVX1_LOC_43/Y VSS 0.26fF
C29565 NAND2X1_LOC_79/Y VSS 0.11fF
C29566 NAND2X1_LOC_69/B VSS 0.27fF
C29567 INVX1_LOC_73/Y VSS 0.06fF
C29568 NAND2X1_LOC_57/Y VSS 0.19fF
C29569 NAND2X1_LOC_13/Y VSS 0.48fF
C29570 INVX1_LOC_51/A VSS 0.23fF
C29571 INVX1_LOC_52/Y VSS 0.25fF
C29572 INVX1_LOC_268/A VSS 0.12fF
C29573 INVX1_LOC_246/Y VSS 0.25fF
C29574 INVX1_LOC_257/Y VSS 0.19fF
C29575 INVX1_LOC_279/Y VSS 0.16fF
C29576 INVX1_LOC_279/A VSS -0.05fF
C29577 INVX1_LOC_213/Y VSS 0.54fF
C29578 INVX1_LOC_11/Y VSS 1.04fF
C29579 NAND2X1_LOC_460/A VSS 0.21fF
C29580 NAND2X1_LOC_379/Y VSS 0.09fF
C29581 INVX1_LOC_438/Y VSS 0.22fF
C29582 INVX1_LOC_438/A VSS -1.52fF
C29583 INVX1_LOC_405/A VSS 0.20fF
C29584 INVX1_LOC_416/A VSS 0.02fF
C29585 INVX1_LOC_449/A VSS 0.34fF
C29586 NAND2X1_LOC_331/A VSS 0.24fF
C29587 NAND2X1_LOC_636/A VSS 0.26fF
C29588 INVX1_LOC_435/A VSS 0.69fF
C29589 INVX1_LOC_432/Y VSS 0.09fF
C29590 INVX1_LOC_421/Y VSS 0.29fF
C29591 INVX1_LOC_608/Y VSS 0.34fF
C29592 INVX1_LOC_616/A VSS 0.12fF
C29593 INVX1_LOC_85/Y VSS 0.49fF
C29594 INVX1_LOC_587/Y VSS 0.08fF
C29595 INVX1_LOC_588/Y VSS -0.48fF
C29596 NAND2X1_LOC_97/B VSS 0.40fF
C29597 GATE_741 VSS -0.05fF
C29598 INVX1_LOC_583/Y VSS 0.25fF
C29599 INVX1_LOC_574/A VSS 0.20fF
C29600 INVX1_LOC_627/A VSS 0.17fF
C29601 INVX1_LOC_612/Y VSS 0.08fF
C29602 INVX1_LOC_563/A VSS 0.12fF
C29603 NAND2X1_LOC_669/Y VSS 0.25fF
C29604 INVX1_LOC_174/Y VSS 0.23fF
C29605 INVX1_LOC_195/A VSS 0.08fF
C29606 INVX1_LOC_191/Y VSS -0.11fF
C29607 INVX1_LOC_43/A VSS 0.26fF
C29608 NAND2X1_LOC_32/Y VSS 0.02fF
C29609 NAND2X1_LOC_27/Y VSS 0.31fF
C29610 INVX1_LOC_80/Y VSS 0.06fF
C29611 INVX1_LOC_32/A VSS 0.12fF
C29612 NAND2X1_LOC_97/A VSS 0.05fF
C29613 NAND2X1_LOC_45/Y VSS 0.47fF
C29614 INVX1_LOC_201/Y VSS 0.23fF
C29615 INVX1_LOC_201/A VSS 0.26fF
C29616 INVX1_LOC_267/Y VSS 0.17fF
C29617 INVX1_LOC_317/Y VSS 0.12fF
C29618 INVX1_LOC_404/Y VSS 0.06fF
C29619 INVX1_LOC_224/Y VSS 0.55fF
C29620 INVX1_LOC_426/Y VSS 0.28fF
C29621 INVX1_LOC_426/A VSS 0.17fF
C29622 INVX1_LOC_415/Y VSS 0.14fF
C29623 INVX1_LOC_218/Y VSS 0.15fF
C29624 INVX1_LOC_448/A VSS 0.36fF
C29625 INVX1_LOC_434/A VSS -0.36fF
C29626 INVX1_LOC_433/Y VSS 0.31fF
C29627 NAND2X1_LOC_635/B VSS 0.23fF
C29628 INVX1_LOC_434/Y VSS 0.25fF
C29629 INVX1_LOC_459/Y VSS 0.25fF
C29630 INVX1_LOC_629/Y VSS 0.31fF
C29631 INVX1_LOC_629/A VSS 0.39fF
C29632 INVX1_LOC_7/A VSS 0.05fF
C29633 INVX1_LOC_618/A VSS 0.12fF
C29634 INVX1_LOC_607/Y VSS -2.46fF
C29635 INVX1_LOC_595/Y VSS 0.19fF
C29636 INVX1_LOC_604/Y VSS 0.29fF
C29637 INVX1_LOC_603/Y VSS -0.31fF
C29638 INVX1_LOC_602/A VSS -1.44fF
C29639 INVX1_LOC_587/A VSS 0.49fF
C29640 INVX1_LOC_584/A VSS 0.28fF
C29641 INVX1_LOC_573/A VSS 0.23fF
C29642 INVX1_LOC_571/Y VSS 0.23fF
C29643 INVX1_LOC_626/A VSS 0.29fF
C29644 INVX1_LOC_613/Y VSS 0.15fF
C29645 INVX1_LOC_176/Y VSS -0.05fF
C29646 INVX1_LOC_175/Y VSS 0.25fF
C29647 NAND2X1_LOC_231/A VSS 0.27fF
C29648 INVX1_LOC_193/Y VSS 0.37fF
C29649 INVX1_LOC_192/Y VSS 0.25fF
C29650 NAND2X1_LOC_88/Y VSS 0.37fF
C29651 INVX1_LOC_95/Y VSS 0.12fF
C29652 INVX1_LOC_288/Y VSS -0.06fF
C29653 INVX1_LOC_42/A VSS 0.12fF
C29654 NAND2X1_LOC_24/Y VSS 0.37fF
C29655 NAND2X1_LOC_20/Y VSS 0.11fF
C29656 INVX1_LOC_31/A VSS 0.47fF
C29657 INVX1_LOC_19/Y VSS 0.23fF
C29658 INVX1_LOC_71/Y VSS -0.09fF
C29659 INVX1_LOC_62/A VSS 0.12fF
C29660 INVX1_LOC_78/A VSS 0.09fF
C29661 INVX1_LOC_21/Y VSS -4.70fF
C29662 INVX1_LOC_266/A VSS 0.63fF
C29663 INVX1_LOC_233/Y VSS 0.08fF
C29664 INVX1_LOC_200/Y VSS 0.13fF
C29665 VDD VSS 2.22fF
C29666 INVX1_LOC_222/Y VSS 0.06fF
C29667 INVX1_LOC_447/Y VSS 0.44fF
C29668 INVX1_LOC_436/A VSS 0.10fF
C29669 INVX1_LOC_425/A VSS -0.25fF
C29670 INVX1_LOC_414/Y VSS 0.04fF
C29671 INPUT_0 VSS 0.75fF
C29672 INVX1_LOC_454/A VSS 0.10fF
C29673 INVX1_LOC_3/Y VSS 0.69fF
C29674 INPUT_6 VSS -0.57fF
C29675 INVX1_LOC_459/A VSS -0.27fF
C29676 INVX1_LOC_437/Y VSS -0.15fF
C29677 INVX1_LOC_436/Y VSS 0.16fF
C29678 INVX1_LOC_628/Y VSS 0.21fF
C29679 INVX1_LOC_628/A VSS 0.15fF
C29680 INVX1_LOC_617/Y VSS 0.47fF
C29681 INVX1_LOC_617/A VSS 0.17fF
C29682 NAND2X1_LOC_789/B VSS 0.11fF
C29683 NAND2X1_LOC_750/Y VSS 0.35fF
C29684 INVX1_LOC_601/A VSS -0.98fF
C29685 INVX1_LOC_625/A VSS -0.00fF
C29686 INVX1_LOC_614/A VSS -1.06fF
C29687 INVX1_LOC_605/Y VSS 0.25fF
C29688 INVX1_LOC_582/Y VSS 0.04fF
C29689 INVX1_LOC_182/A VSS 0.30fF
C29690 INVX1_LOC_177/Y VSS 0.25fF
C29691 NAND2X1_LOC_242/A VSS 0.23fF
C29692 INVX1_LOC_202/A VSS 0.12fF
C29693 NAND2X1_LOC_7/Y VSS 0.33fF
C29694 INVX1_LOC_193/A VSS 0.39fF
C29695 INVX1_LOC_333/Y VSS 0.29fF
C29696 INVX1_LOC_335/Y VSS 0.22fF
C29697 NAND2X1_LOC_88/B VSS 0.11fF
C29698 NAND2X1_LOC_65/Y VSS 0.11fF
C29699 INVX1_LOC_68/Y VSS 0.43fF
C29700 NAND2X1_LOC_93/Y VSS 0.20fF
C29701 INVX1_LOC_254/Y VSS -0.19fF
C29702 INVX1_LOC_298/Y VSS 0.28fF
C29703 INVX1_LOC_287/A VSS 0.27fF
C29704 INVX1_LOC_276/A VSS 0.07fF
C29705 INVX1_LOC_30/Y VSS 0.06fF
C29706 INVX1_LOC_210/Y VSS -0.08fF
C29707 INVX1_LOC_243/A VSS 0.12fF
C29708 INVX1_LOC_20/Y VSS -3.43fF
C29709 INVX1_LOC_435/Y VSS -5.72fF
C29710 INVX1_LOC_457/Y VSS 0.25fF
C29711 INVX1_LOC_424/A VSS 0.31fF
C29712 INVX1_LOC_446/A VSS 0.43fF
C29713 INVX1_LOC_402/Y VSS 0.39fF
C29714 INVX1_LOC_402/A VSS 0.18fF
C29715 GATE_579 VSS 0.10fF
C29716 INVX1_LOC_452/Y VSS 0.25fF
.ends

