magic
tech scmos
magscale 1 2
timestamp 1602073617
<< metal1 >>
rect 7140 8957 7203 8963
rect 7828 8957 7848 8963
rect 1988 8937 2003 8943
rect 3338 8936 3340 8944
rect 5165 8937 5196 8943
rect 7076 8936 7078 8944
rect 8538 8936 8540 8944
rect 2628 8917 2648 8923
rect 3981 8897 3996 8903
rect 5818 8897 5875 8903
rect 11018 8897 11075 8903
rect 5786 8876 5788 8884
rect 6429 8877 6444 8883
rect 9677 8877 9692 8883
rect 10365 8877 10396 8883
rect 10986 8876 10988 8884
rect 1332 8837 1348 8843
rect 676 8757 707 8763
rect 1972 8757 2003 8763
rect 4509 8757 4572 8763
rect 5876 8757 5907 8763
rect 7172 8757 7203 8763
rect 9780 8757 9798 8763
rect 10436 8757 10451 8763
rect 3868 8737 3900 8743
rect 12276 8736 12278 8744
rect 1220 8717 1235 8723
rect 3332 8717 3347 8723
rect 6493 8717 6548 8723
rect 11780 8717 11795 8723
rect 3213 8697 3228 8703
rect 3252 8697 3268 8703
rect 3260 8686 3268 8697
rect 5196 8697 5212 8703
rect 5196 8692 5204 8697
rect 11661 8697 11692 8703
rect 10397 8677 10412 8683
rect 4580 8637 4598 8643
rect 644 8577 707 8583
rect 1332 8577 1348 8583
rect 2596 8577 2648 8583
rect 4509 8577 4540 8583
rect 5818 8577 5836 8583
rect 8468 8577 8499 8583
rect 11661 8577 11676 8583
rect 7796 8557 7848 8563
rect 5197 8537 5219 8543
rect 8538 8536 8540 8544
rect 9748 8537 9763 8543
rect 10324 8536 10328 8544
rect 11044 8537 11062 8543
rect 12228 8537 12278 8543
rect 4596 8516 4598 8524
rect 3868 8497 3923 8503
rect 9828 8496 9830 8504
rect 11780 8497 11795 8503
rect 618 8477 684 8483
rect 7736 8476 7740 8484
rect 7876 8476 7880 8484
rect 11018 8477 11036 8483
rect 3236 8377 3299 8383
rect 5165 8377 5196 8383
rect 7117 8377 7132 8383
rect 9796 8376 9798 8384
rect 676 8357 707 8363
rect 3940 8357 3955 8363
rect 7828 8357 7848 8363
rect 5786 8336 5788 8344
rect 7876 8336 7880 8344
rect 9828 8336 9830 8344
rect 10986 8336 10988 8344
rect 11018 8337 11036 8343
rect 1293 8317 1348 8323
rect 3885 8317 3900 8323
rect 5818 8317 5875 8323
rect 6461 8317 6508 8323
rect 9068 8317 9123 8323
rect 11684 8317 11731 8323
rect 1972 8297 2003 8303
rect 6500 8297 6516 8303
rect 11661 8297 11692 8303
rect 4556 8286 4564 8296
rect 6508 8286 6516 8297
rect 1949 8277 1964 8283
rect 3901 8277 3916 8283
rect 10397 8277 10419 8283
rect 11700 8277 11715 8283
rect 12276 8276 12278 8284
rect 12317 8237 12332 8243
rect 2568 8176 2572 8184
rect 5165 8177 5180 8183
rect 8413 8177 8428 8183
rect 9732 8177 9798 8183
rect 11661 8177 11676 8183
rect 4548 8137 4563 8143
rect 5124 8136 5128 8144
rect 5288 8136 5292 8144
rect 10397 8137 10419 8143
rect 1876 8116 1878 8124
rect 7768 8117 7788 8123
rect 9709 8117 9772 8123
rect 1220 8097 1235 8103
rect 3868 8097 3900 8103
rect 4628 8096 4630 8104
rect 11018 8096 11020 8104
rect 11044 8097 11075 8103
rect 1917 8077 1948 8083
rect 7736 8076 7740 8084
rect 10986 8076 10988 8084
rect 2568 7977 2620 7983
rect 2644 7976 2648 7984
rect 8436 7977 8499 7983
rect 10365 7977 10380 7983
rect 10388 7957 10451 7963
rect 10324 7936 10328 7944
rect 1818 7916 1820 7924
rect 4628 7923 4630 7924
rect 4628 7917 4643 7923
rect 4628 7916 4630 7917
rect 88 7876 92 7884
rect 6500 7877 6515 7883
rect 5818 7836 5820 7844
rect 7188 7837 7203 7843
rect 2644 7776 2648 7784
rect 5236 7777 5251 7783
rect 8413 7777 8428 7783
rect 9709 7777 9740 7783
rect 11018 7776 11020 7784
rect 20 7757 51 7763
rect 88 7736 92 7744
rect 5197 7737 5212 7743
rect 10324 7736 10328 7744
rect 12276 7736 12278 7744
rect 7076 7716 7078 7724
rect 7768 7717 7788 7723
rect 3981 7697 3996 7703
rect 7117 7697 7148 7703
rect 8532 7697 8547 7703
rect 9092 7697 9123 7703
rect 10365 7697 10396 7703
rect 4532 7677 4598 7683
rect 7736 7676 7740 7684
rect 5892 7637 5907 7643
rect 1261 7577 1276 7583
rect 5188 7577 5251 7583
rect 8413 7577 8428 7583
rect 11018 7577 11036 7583
rect 7188 7557 7203 7563
rect 586 7536 588 7544
rect 1917 7537 1980 7543
rect 11629 7537 11644 7543
rect 1380 7517 1395 7523
rect 1940 7517 2003 7523
rect 3981 7517 3996 7523
rect 4628 7523 4630 7524
rect 4628 7517 4643 7523
rect 4628 7516 4630 7517
rect 11661 7517 11731 7523
rect 1300 7497 1316 7503
rect 1308 7486 1316 7497
rect 3252 7497 3268 7503
rect 3260 7486 3268 7497
rect 8538 7496 8540 7504
rect 9709 7497 9740 7503
rect 7149 7477 7164 7483
rect 11700 7477 11715 7483
rect 36 7377 51 7383
rect 4532 7377 4598 7383
rect 9068 7377 9084 7383
rect 4509 7357 4540 7363
rect 9709 7357 9772 7363
rect 5288 7337 5340 7343
rect 7076 7336 7078 7344
rect 10397 7337 10419 7343
rect 12276 7336 12278 7344
rect 5220 7317 5251 7323
rect 7668 7296 7670 7304
rect 11780 7297 11795 7303
rect 3868 7277 3884 7283
rect 5876 7237 5907 7243
rect 11018 7236 11020 7244
rect 4596 7176 4598 7184
rect 7844 7176 7848 7184
rect 9709 7177 9724 7183
rect 1972 7157 2003 7163
rect 5844 7157 5907 7163
rect 4628 7136 4630 7144
rect 7736 7136 7740 7144
rect 9068 7137 9100 7143
rect 9677 7137 9692 7143
rect 10986 7136 10988 7144
rect 11629 7137 11644 7143
rect 1293 7117 1348 7123
rect 2468 7116 2470 7124
rect 6516 7117 6548 7123
rect 7069 7117 7084 7123
rect 9709 7117 9782 7123
rect 11018 7117 11075 7123
rect 11661 7117 11731 7123
rect 3338 7096 3340 7104
rect 5197 7077 5219 7083
rect 11700 7077 11715 7083
rect 12276 7076 12278 7084
rect 2628 7037 2648 7043
rect 10365 7037 10380 7043
rect 12317 7037 12332 7043
rect 3940 6977 3955 6983
rect 5165 6977 5180 6983
rect 6461 6977 6476 6983
rect 7796 6977 7848 6983
rect 10365 6977 10396 6983
rect 11661 6977 11676 6983
rect 11716 6977 11748 6983
rect 7768 6957 7820 6963
rect 2596 6937 2612 6943
rect 3252 6937 3267 6943
rect 6500 6937 6515 6943
rect 10324 6936 10328 6944
rect 2568 6917 2588 6923
rect 7076 6916 7078 6924
rect 1293 6897 1324 6903
rect 4628 6896 4630 6904
rect 9068 6897 9100 6903
rect 11044 6897 11075 6903
rect 88 6876 92 6884
rect 2536 6876 2540 6884
rect 3181 6877 3196 6883
rect 7117 6877 7148 6883
rect 9709 6877 9740 6883
rect 618 6776 620 6784
rect 2568 6776 2572 6784
rect 11018 6777 11036 6783
rect 1917 6737 1948 6743
rect 5933 6737 5948 6743
rect 9068 6737 9100 6743
rect 10986 6736 10988 6744
rect 5165 6717 5222 6723
rect 10365 6717 10396 6723
rect 11044 6717 11075 6723
rect 1876 6696 1878 6704
rect 5124 6696 5128 6704
rect 10324 6696 10328 6704
rect 8452 6677 8467 6683
rect 10404 6677 10419 6683
rect 4532 6577 4598 6583
rect 8468 6577 8499 6583
rect 9140 6557 9155 6563
rect 1949 6537 1964 6543
rect 5197 6537 5219 6543
rect 6500 6537 6515 6543
rect 7844 6536 7848 6544
rect 9101 6537 9116 6543
rect 11076 6517 11107 6523
rect 4509 6497 4572 6503
rect 3213 6477 3244 6483
rect 3868 6477 3900 6483
rect 5818 6477 5852 6483
rect 9828 6476 9830 6484
rect 10456 6476 10460 6484
rect 618 6436 620 6444
rect 692 6437 707 6443
rect 7188 6437 7203 6443
rect 6461 6377 6476 6383
rect 7828 6377 7848 6383
rect 11661 6377 11724 6383
rect 676 6357 707 6363
rect 4532 6337 4598 6343
rect 5786 6336 5788 6344
rect 9677 6337 9692 6343
rect 10986 6336 10988 6344
rect 1818 6316 1820 6324
rect 2746 6316 2748 6324
rect 3981 6317 3996 6323
rect 5818 6317 5875 6323
rect 7768 6317 7820 6323
rect 9709 6317 9782 6323
rect 10365 6317 10422 6323
rect 11018 6317 11075 6323
rect 12269 6317 12284 6323
rect 9748 6297 9764 6303
rect 9756 6286 9764 6297
rect 10404 6297 10420 6303
rect 10412 6292 10420 6297
rect 2516 6277 2531 6283
rect 2596 6277 2612 6283
rect 5197 6277 5219 6283
rect 2568 6236 2572 6244
rect 4509 6237 4524 6243
rect 6484 6237 6548 6243
rect 9092 6177 9155 6183
rect 1972 6157 2003 6163
rect 2628 6157 2648 6163
rect 88 6136 92 6144
rect 692 6137 707 6143
rect 5288 6136 5292 6144
rect 7076 6136 7078 6144
rect 10397 6137 10419 6143
rect 4556 6123 4564 6134
rect 4548 6117 4564 6123
rect 11661 6117 11692 6123
rect 1293 6097 1324 6103
rect 4509 6077 4556 6083
rect 7876 6076 7880 6084
rect 11018 6077 11036 6083
rect 7844 6036 7848 6044
rect 2568 5977 2588 5983
rect 3213 5977 3260 5983
rect 7117 5977 7148 5983
rect 8484 5977 8499 5983
rect 88 5936 92 5944
rect 5786 5936 5788 5944
rect 6429 5937 6444 5943
rect 7736 5936 7740 5944
rect 10986 5936 10988 5944
rect 11629 5937 11644 5943
rect 6500 5917 6531 5923
rect 9085 5917 9139 5923
rect 10365 5917 10396 5923
rect 11661 5917 11731 5923
rect 1261 5897 1324 5903
rect 7768 5897 7788 5903
rect 9748 5897 9764 5903
rect 9756 5886 9764 5897
rect 2596 5877 2612 5883
rect 5197 5877 5219 5883
rect 5844 5877 5862 5883
rect 7796 5877 7812 5883
rect 8538 5877 8556 5883
rect 10324 5876 10328 5884
rect 12276 5876 12278 5884
rect 5818 5836 5820 5844
rect 8452 5837 8499 5843
rect 1332 5777 1348 5783
rect 3284 5777 3299 5783
rect 6461 5777 6476 5783
rect 6500 5777 6548 5783
rect 11661 5777 11692 5783
rect 7188 5757 7203 5763
rect 5236 5737 5251 5743
rect 7149 5737 7164 5743
rect 10324 5736 10328 5744
rect 12349 5737 12364 5743
rect 5196 5723 5204 5728
rect 5196 5717 5212 5723
rect 12269 5697 12284 5703
rect 9709 5677 9740 5683
rect 11018 5677 11052 5683
rect 1988 5637 2003 5643
rect 1332 5577 1348 5583
rect 5188 5577 5251 5583
rect 9068 5577 9084 5583
rect 20 5557 51 5563
rect 2644 5556 2648 5564
rect 12968 5556 12972 5564
rect 5860 5537 5907 5543
rect 10986 5536 10988 5544
rect 3821 5517 3836 5523
rect 4541 5517 4556 5523
rect 7946 5516 7948 5524
rect 8413 5517 8444 5523
rect 12317 5517 12372 5523
rect 7172 5497 7203 5503
rect 11708 5486 11716 5496
rect 3338 5476 3340 5484
rect 10397 5477 10419 5483
rect 9732 5437 9798 5443
rect 618 5376 620 5384
rect 1972 5377 2003 5383
rect 5818 5376 5820 5384
rect 6484 5377 6548 5383
rect 7812 5377 7848 5383
rect 8484 5377 8499 5383
rect 11044 5377 11107 5383
rect 9796 5356 9798 5364
rect 3338 5337 3388 5343
rect 9101 5337 9116 5343
rect 10397 5337 10419 5343
rect 3900 5323 3908 5334
rect 3900 5317 3916 5323
rect 5124 5316 5128 5324
rect 12276 5316 12278 5324
rect 3821 5297 3836 5303
rect 9741 5297 9772 5303
rect 692 5277 707 5283
rect 5818 5277 5836 5283
rect 7736 5276 7740 5284
rect 10986 5276 10988 5284
rect 12317 5277 12348 5283
rect 9124 5257 9155 5263
rect 12968 5236 12972 5244
rect 618 5177 636 5183
rect 3868 5177 3884 5183
rect 644 5157 707 5163
rect 9796 5156 9798 5164
rect 586 5136 588 5144
rect 1997 5137 2012 5143
rect 7117 5137 7148 5143
rect 9828 5136 9830 5144
rect 10986 5136 10988 5144
rect 3213 5117 3228 5123
rect 3981 5117 3996 5123
rect 9741 5117 9772 5123
rect 11661 5117 11724 5123
rect 5876 5097 5907 5103
rect 7076 5096 7078 5104
rect 3252 5077 3267 5083
rect 4548 5077 4563 5083
rect 5124 5076 5128 5084
rect 10397 5077 10419 5083
rect 12349 5077 12364 5083
rect 5818 5037 5836 5043
rect 7768 5036 7772 5044
rect 9124 5037 9155 5043
rect 3268 4977 3299 4983
rect 4596 4976 4598 4984
rect 7117 4977 7132 4983
rect 12968 4976 12972 4984
rect 6461 4957 6476 4963
rect 2644 4936 2648 4944
rect 5197 4937 5219 4943
rect 6500 4937 6515 4943
rect 9748 4937 9763 4943
rect 12884 4937 12931 4943
rect 3900 4923 3908 4934
rect 3900 4917 3916 4923
rect 5818 4897 5852 4903
rect 11661 4897 11692 4903
rect 6429 4877 6444 4883
rect 10365 4877 10396 4883
rect 7140 4837 7203 4843
rect 11018 4836 11020 4844
rect 7188 4777 7203 4783
rect 7844 4776 7848 4784
rect 9796 4776 9798 4784
rect 11684 4777 11748 4783
rect 5204 4757 5251 4763
rect 10436 4757 10451 4763
rect 88 4736 92 4744
rect 1316 4737 1348 4743
rect 2536 4736 2540 4744
rect 7220 4737 7235 4743
rect 9828 4736 9830 4744
rect 4628 4723 4630 4724
rect 4628 4717 4643 4723
rect 4628 4716 4630 4717
rect 8596 4716 8598 4724
rect 10396 4697 10412 4703
rect 10396 4692 10404 4697
rect 11661 4697 11724 4703
rect 12348 4697 12364 4703
rect 12348 4686 12356 4697
rect 5108 4677 5128 4683
rect 7149 4677 7164 4683
rect 9709 4637 9724 4643
rect 5818 4576 5820 4584
rect 5844 4577 5907 4583
rect 7828 4577 7848 4583
rect 9780 4577 9798 4583
rect 11060 4577 11107 4583
rect 20 4557 51 4563
rect 9092 4557 9155 4563
rect 88 4536 92 4544
rect 4548 4537 4563 4543
rect 10397 4537 10419 4543
rect 12349 4537 12364 4543
rect 5212 4523 5220 4528
rect 5204 4517 5220 4523
rect 1220 4497 1235 4503
rect 3868 4497 3923 4503
rect 6580 4497 6595 4503
rect 9741 4497 9772 4503
rect 12269 4497 12284 4503
rect 4477 4477 4492 4483
rect 3213 4437 3228 4443
rect 11018 4436 11020 4444
rect 2628 4377 2648 4383
rect 5892 4377 5907 4383
rect 3892 4357 3955 4363
rect 9140 4357 9155 4363
rect 9828 4336 9830 4344
rect 12317 4337 12348 4343
rect 2468 4316 2470 4324
rect 6420 4317 6435 4323
rect 9085 4317 9100 4323
rect 9741 4317 9798 4323
rect 11661 4317 11708 4323
rect 7768 4297 7788 4303
rect 9100 4297 9116 4303
rect 9100 4286 9108 4297
rect 11700 4297 11716 4303
rect 11708 4286 11716 4297
rect 7076 4276 7078 4284
rect 10397 4277 10419 4283
rect 11044 4277 11062 4283
rect 11018 4236 11020 4244
rect 12968 4236 12972 4244
rect 1972 4177 2003 4183
rect 4532 4177 4598 4183
rect 5818 4176 5820 4184
rect 3252 4137 3267 4143
rect 5197 4137 5219 4143
rect 7076 4136 7078 4144
rect 8452 4137 8467 4143
rect 9748 4137 9763 4143
rect 10324 4136 10328 4144
rect 10488 4136 10492 4144
rect 11684 4137 11748 4143
rect 12349 4137 12364 4143
rect 3332 4097 3347 4103
rect 3868 4097 3923 4103
rect 6644 4096 6648 4104
rect 12269 4097 12284 4103
rect 7768 4077 7788 4083
rect 11661 4077 11724 4083
rect 692 4057 707 4063
rect 618 3976 620 3984
rect 2644 3976 2648 3984
rect 5818 3977 5868 3983
rect 7796 3977 7848 3983
rect 11092 3977 11107 3983
rect 9140 3957 9155 3963
rect 9796 3956 9798 3964
rect 3338 3936 3340 3944
rect 5165 3937 5212 3943
rect 7736 3936 7740 3944
rect 8468 3937 8499 3943
rect 12308 3936 12310 3944
rect 6644 3916 6648 3924
rect 11620 3917 11635 3923
rect 11844 3916 11848 3924
rect 5124 3896 5128 3904
rect 8538 3896 8540 3904
rect 9100 3897 9116 3903
rect 9100 3886 9108 3897
rect 2516 3877 2531 3883
rect 9997 3864 10003 3896
rect 11708 3886 11716 3896
rect 10397 3877 10412 3883
rect 10488 3876 10492 3884
rect 12276 3876 12278 3884
rect 10436 3837 10451 3843
rect 12317 3837 12364 3843
rect 2568 3777 2620 3783
rect 4509 3777 4540 3783
rect 7768 3776 7772 3784
rect 88 3736 92 3744
rect 6500 3737 6515 3743
rect 8452 3737 8467 3743
rect 1380 3697 1395 3703
rect 3908 3697 3939 3703
rect 4628 3703 4630 3704
rect 4628 3697 4643 3703
rect 4628 3696 4630 3697
rect 7946 3696 7948 3704
rect 11018 3697 11075 3703
rect 12269 3697 12284 3703
rect 1229 3677 1244 3683
rect 1917 3677 1948 3683
rect 7076 3676 7078 3684
rect 10986 3676 10988 3684
rect 2596 3657 2648 3663
rect 5204 3637 5251 3643
rect 12388 3637 12403 3643
rect 644 3577 707 3583
rect 2612 3577 2648 3583
rect 5165 3577 5180 3583
rect 5818 3577 5836 3583
rect 2676 3536 2680 3544
rect 5124 3536 5128 3544
rect 10986 3536 10988 3544
rect 3885 3517 3900 3523
rect 5188 3517 5222 3523
rect 6461 3517 6492 3523
rect 6580 3517 6595 3523
rect 7768 3517 7804 3523
rect 8413 3497 8444 3503
rect 4548 3477 4563 3483
rect 6500 3477 6515 3483
rect 9068 3477 9084 3483
rect 10397 3477 10419 3483
rect 12349 3477 12364 3483
rect 7117 3437 7132 3443
rect 9796 3436 9798 3444
rect 3868 3377 3916 3383
rect 3940 3377 3955 3383
rect 5876 3377 5907 3383
rect 10388 3377 10451 3383
rect 12968 3376 12972 3384
rect 9140 3357 9155 3363
rect 88 3336 92 3344
rect 1988 3337 2003 3343
rect 5236 3337 5251 3343
rect 9101 3337 9116 3343
rect 10488 3336 10492 3344
rect 9756 3324 9764 3334
rect 12276 3316 12278 3324
rect 7768 3297 7804 3303
rect 10365 3297 10428 3303
rect 12317 3277 12348 3283
rect 1917 3177 1964 3183
rect 3940 3177 3955 3183
rect 5236 3177 5251 3183
rect 11018 3177 11036 3183
rect 12968 3176 12972 3184
rect 2628 3157 2648 3163
rect 4596 3156 4598 3164
rect 5876 3157 5907 3163
rect 88 3136 92 3144
rect 7117 3137 7148 3143
rect 10986 3136 10988 3144
rect 11629 3137 11644 3143
rect 12317 3137 12348 3143
rect 6580 3117 6595 3123
rect 9068 3117 9123 3123
rect 11780 3117 11795 3123
rect 1300 3097 1316 3103
rect 1308 3086 1316 3097
rect 7076 3096 7078 3104
rect 3338 3077 3356 3083
rect 5197 3077 5212 3083
rect 8413 3077 8444 3083
rect 9837 3077 9852 3083
rect 10397 3077 10419 3083
rect 11661 3077 11692 3083
rect 7768 3037 7788 3043
rect 9796 3036 9798 3044
rect 3213 2977 3276 2983
rect 7844 2976 7848 2984
rect 676 2957 707 2963
rect 2596 2937 2612 2943
rect 5124 2936 5128 2944
rect 11044 2937 11062 2943
rect 10324 2916 10328 2924
rect 1293 2897 1324 2903
rect 5818 2897 5836 2903
rect 11780 2897 11795 2903
rect 2568 2877 2588 2883
rect 9709 2877 9756 2883
rect 5165 2837 5196 2843
rect 6484 2837 6548 2843
rect 11018 2836 11020 2844
rect 676 2757 707 2763
rect 2644 2756 2648 2764
rect 7828 2757 7848 2763
rect 9140 2757 9155 2763
rect 7876 2736 7880 2744
rect 10986 2736 10988 2744
rect 1818 2716 1820 2724
rect 6493 2717 6548 2723
rect 8444 2717 8499 2723
rect 9085 2717 9100 2723
rect 9828 2723 9830 2724
rect 9828 2717 9843 2723
rect 9828 2716 9830 2717
rect 9100 2697 9116 2703
rect 9100 2686 9108 2697
rect 88 2676 92 2684
rect 5204 2677 5219 2683
rect 12276 2676 12278 2684
rect 12317 2637 12348 2643
rect 618 2576 620 2584
rect 644 2577 707 2583
rect 3213 2577 3260 2583
rect 4596 2576 4598 2584
rect 5892 2577 5907 2583
rect 3338 2536 3340 2544
rect 8452 2537 8467 2543
rect 9748 2537 9763 2543
rect 10388 2537 10451 2543
rect 10488 2536 10492 2544
rect 1869 2497 1884 2503
rect 3821 2497 3836 2503
rect 7946 2496 7948 2504
rect 5288 2476 5292 2484
rect 3940 2437 3955 2443
rect 5892 2437 5907 2443
rect 618 2376 620 2384
rect 4596 2376 4598 2384
rect 9796 2376 9798 2384
rect 10436 2377 10451 2383
rect 644 2357 707 2363
rect 2628 2357 2648 2363
rect 11076 2357 11107 2363
rect 2676 2336 2680 2344
rect 7736 2336 7740 2344
rect 7946 2316 7948 2324
rect 11780 2317 11795 2323
rect 4637 2297 4684 2303
rect 5197 2277 5219 2283
rect 6500 2277 6515 2283
rect 7796 2277 7812 2283
rect 10397 2277 10412 2283
rect 3236 2177 3299 2183
rect 11661 2157 11676 2163
rect 1988 2137 2003 2143
rect 3338 2136 3340 2144
rect 5197 2137 5219 2143
rect 7188 2137 7203 2143
rect 8452 2137 8467 2143
rect 10324 2136 10328 2144
rect 11700 2137 11715 2143
rect 1948 2123 1956 2134
rect 1948 2117 1964 2123
rect 3900 2123 3908 2134
rect 3900 2117 3916 2123
rect 7148 2123 7156 2134
rect 7148 2117 7164 2123
rect 10412 2123 10420 2128
rect 10404 2117 10420 2123
rect 1869 2097 1884 2103
rect 11780 2097 11795 2103
rect 3908 2077 3955 2083
rect 4628 2076 4630 2084
rect 5786 2076 5788 2084
rect 11018 2077 11036 2083
rect 11629 2077 11644 2083
rect 5818 1976 5820 1984
rect 5892 1977 5907 1983
rect 7796 1977 7848 1983
rect 88 1936 92 1944
rect 2676 1936 2680 1944
rect 5786 1936 5788 1944
rect 7117 1937 7148 1943
rect 10356 1936 10360 1944
rect 12276 1936 12278 1944
rect 5165 1917 5196 1923
rect 6493 1917 6531 1923
rect 9021 1917 9036 1923
rect 11844 1916 11848 1924
rect 4548 1877 4563 1883
rect 11700 1877 11715 1883
rect 676 1777 707 1783
rect 1988 1777 2003 1783
rect 2628 1777 2648 1783
rect 3940 1777 3955 1783
rect 5165 1777 5196 1783
rect 8436 1777 8499 1783
rect 9709 1777 9724 1783
rect 7768 1757 7788 1763
rect 1876 1736 1878 1744
rect 5124 1736 5128 1744
rect 5844 1737 5862 1743
rect 6500 1737 6515 1743
rect 8538 1736 8540 1744
rect 9732 1737 9798 1743
rect 10488 1736 10492 1744
rect 3900 1723 3908 1734
rect 3900 1717 3916 1723
rect 7076 1716 7078 1724
rect 10396 1723 10404 1728
rect 11708 1724 11716 1734
rect 10396 1717 10412 1723
rect 1380 1697 1395 1703
rect 3821 1697 3836 1703
rect 9021 1697 9036 1703
rect 9181 1697 9196 1703
rect 10986 1703 10988 1704
rect 10973 1697 10988 1703
rect 10986 1696 10988 1697
rect 11060 1697 11107 1703
rect 7117 1677 7148 1683
rect 9828 1676 9830 1684
rect 12308 1676 12310 1684
rect 8413 1657 8476 1663
rect 3940 1637 3955 1643
rect 1917 1577 1948 1583
rect 3213 1577 3228 1583
rect 7844 1576 7848 1584
rect 10365 1577 10380 1583
rect 11700 1577 11748 1583
rect 9092 1557 9155 1563
rect 10388 1557 10451 1563
rect 724 1537 739 1543
rect 1876 1536 1878 1544
rect 2536 1536 2540 1544
rect 7220 1537 7235 1543
rect 7876 1536 7880 1544
rect 634 1517 707 1523
rect 3981 1517 3996 1523
rect 4509 1517 4556 1523
rect 6420 1517 6435 1523
rect 10986 1523 10988 1524
rect 10973 1517 10988 1523
rect 10986 1516 10988 1517
rect 3252 1477 3267 1483
rect 4548 1477 4563 1483
rect 5204 1477 5219 1483
rect 7149 1477 7164 1483
rect 618 1376 620 1384
rect 1917 1377 1932 1383
rect 3213 1377 3228 1383
rect 3252 1377 3299 1383
rect 4580 1377 4598 1383
rect 8436 1377 8499 1383
rect 1300 1337 1315 1343
rect 1876 1336 1878 1344
rect 3940 1337 3955 1343
rect 7076 1336 7078 1344
rect 9748 1337 9763 1343
rect 3900 1323 3908 1334
rect 3900 1317 3916 1323
rect 10412 1323 10420 1328
rect 10404 1317 10420 1323
rect 11708 1323 11716 1334
rect 11700 1317 11716 1323
rect 7768 1297 7788 1303
rect 8968 1296 8972 1304
rect 10356 1276 10360 1284
rect 11018 1277 11036 1283
rect 12308 1276 12310 1284
rect 5220 1237 5251 1243
rect 618 1177 636 1183
rect 1917 1177 1932 1183
rect 6461 1177 6524 1183
rect 9709 1177 9724 1183
rect 1261 1157 1292 1163
rect 3213 1157 3244 1163
rect 7188 1157 7203 1163
rect 1229 1137 1244 1143
rect 2536 1136 2540 1144
rect 4628 1136 4630 1144
rect 9068 1137 9100 1143
rect 7668 1116 7670 1124
rect 1300 1077 1315 1083
rect 7149 1077 7164 1083
rect 10397 1077 10412 1083
rect 4509 1037 4524 1043
rect 9796 1036 9798 1044
rect 10436 1037 10451 1043
rect 2568 976 2572 984
rect 3213 977 3228 983
rect 3940 977 3955 983
rect 11018 977 11036 983
rect 5165 957 5228 963
rect 3338 936 3340 944
rect 3900 923 3908 934
rect 11708 924 11716 934
rect 3900 917 3916 923
rect 7069 897 7084 903
rect 618 877 684 883
rect 5288 876 5292 884
rect 9068 877 9100 883
rect 9677 877 9692 883
rect 12308 876 12310 884
rect 1917 837 1948 843
rect 618 777 636 783
rect 1261 777 1276 783
rect 7768 776 7772 784
rect 586 736 588 744
rect 2536 736 2540 744
rect 4509 737 4556 743
rect 7736 736 7740 744
rect 9709 737 9772 743
rect 10986 736 10988 744
rect 2568 697 2588 703
rect 4548 677 4563 683
rect 5124 676 5128 684
rect 7796 677 7812 683
rect 10397 677 10419 683
rect 11788 677 11804 683
rect 9732 637 9798 643
rect 11661 637 11676 643
rect 618 576 620 584
rect 2568 576 2572 584
rect 4532 577 4598 583
rect 7140 577 7203 583
rect 9068 577 9084 583
rect 9709 577 9740 583
rect 5197 537 5219 543
rect 10412 523 10420 528
rect 10404 517 10420 523
rect 11588 517 11635 523
rect 5818 497 5852 503
rect 10365 497 10380 503
rect 4468 477 4483 483
rect 7876 476 7880 484
rect 12308 476 12310 484
rect 4509 437 4572 443
rect 7117 437 7132 443
rect 6461 377 6492 383
rect 12317 377 12380 383
rect 618 357 636 363
rect 11076 357 11107 363
rect 586 336 588 344
rect 4532 337 4598 343
rect 4628 336 4630 344
rect 9677 337 9692 343
rect 3981 317 3996 323
rect 7768 317 7788 323
rect 9092 317 9123 323
rect 3338 296 3340 304
rect 8413 297 8444 303
rect 4509 277 4572 283
rect 9837 277 9852 283
rect 1917 237 1980 243
rect 3213 237 3228 243
rect 7117 237 7132 243
rect 618 177 684 183
rect 1332 177 1348 183
rect 3892 177 3955 183
rect 4580 177 4598 183
rect 11684 177 11748 183
rect 6461 157 6524 163
rect 11661 157 11692 163
rect 5197 137 5219 143
rect 10404 137 10419 143
rect 10365 117 10396 123
rect 9709 97 9756 103
rect 2536 76 2540 84
rect 3181 77 3196 83
rect 7768 77 7804 83
rect 11018 77 11052 83
<< m2contact >>
rect 11628 8990 11636 8998
rect 11660 8990 11668 8998
rect 7116 8976 7124 8984
rect 11740 8976 11748 8984
rect 3292 8956 3300 8964
rect 7132 8956 7140 8964
rect 7820 8956 7828 8964
rect 732 8936 740 8944
rect 1980 8936 1988 8944
rect 2684 8936 2692 8944
rect 3340 8936 3348 8944
rect 5196 8936 5204 8944
rect 7068 8936 7076 8944
rect 7884 8936 7892 8944
rect 8540 8936 8548 8944
rect 11788 8936 11796 8944
rect 2620 8916 2628 8924
rect 4476 8916 4484 8924
rect 8492 8916 8500 8924
rect 1884 8896 1892 8904
rect 3996 8896 4004 8904
rect 5276 8896 5284 8904
rect 6572 8896 6580 8904
rect 9036 8896 9044 8904
rect 5788 8876 5796 8884
rect 6444 8876 6452 8884
rect 9692 8876 9700 8884
rect 10396 8876 10404 8884
rect 10988 8876 10996 8884
rect 44 8836 52 8844
rect 588 8836 596 8844
rect 1324 8836 1332 8844
rect 1884 8836 1892 8844
rect 2540 8836 2548 8844
rect 7740 8836 7748 8844
rect 9036 8836 9044 8844
rect 588 8776 596 8784
rect 1884 8776 1892 8784
rect 2540 8776 2548 8784
rect 5932 8776 5940 8784
rect 7228 8776 7236 8784
rect 7740 8776 7748 8784
rect 9036 8776 9044 8784
rect 9148 8776 9156 8784
rect 668 8756 676 8764
rect 732 8756 740 8764
rect 1340 8756 1348 8764
rect 1964 8756 1972 8764
rect 2028 8756 2036 8764
rect 4572 8756 4580 8764
rect 5868 8756 5876 8764
rect 7164 8756 7172 8764
rect 8492 8756 8500 8764
rect 9772 8756 9780 8764
rect 10428 8756 10436 8764
rect 1388 8736 1396 8744
rect 3900 8736 3908 8744
rect 6572 8736 6580 8744
rect 8524 8736 8532 8744
rect 10476 8736 10484 8744
rect 12268 8736 12276 8744
rect 1164 8716 1172 8724
rect 1212 8716 1220 8724
rect 1884 8716 1892 8724
rect 3324 8716 3332 8724
rect 5132 8716 5140 8724
rect 7084 8716 7092 8724
rect 7724 8716 7732 8724
rect 7884 8716 7892 8724
rect 10332 8716 10340 8724
rect 11772 8716 11780 8724
rect 3228 8696 3236 8704
rect 3244 8696 3252 8704
rect 3820 8696 3828 8704
rect 5212 8696 5220 8704
rect 11692 8696 11700 8704
rect 10412 8676 10420 8684
rect 44 8636 52 8644
rect 4572 8636 4580 8644
rect 5244 8636 5252 8644
rect 8380 8636 8388 8644
rect 8412 8636 8420 8644
rect 636 8576 644 8584
rect 1324 8576 1332 8584
rect 2588 8576 2596 8584
rect 4540 8576 4548 8584
rect 5836 8576 5844 8584
rect 6428 8576 6436 8584
rect 6460 8576 6468 8584
rect 8460 8576 8468 8584
rect 10364 8576 10372 8584
rect 11676 8576 11684 8584
rect 12316 8576 12324 8584
rect 6540 8556 6548 8564
rect 7788 8556 7796 8564
rect 1388 8536 1396 8544
rect 2524 8536 2532 8544
rect 2684 8536 2692 8544
rect 8540 8536 8548 8544
rect 9740 8536 9748 8544
rect 10316 8536 10324 8544
rect 11036 8536 11044 8544
rect 12220 8536 12228 8544
rect 4588 8516 4596 8524
rect 9676 8516 9684 8524
rect 10972 8516 10980 8524
rect 76 8496 84 8504
rect 2040 8496 2048 8504
rect 3116 8496 3124 8504
rect 3168 8496 3176 8504
rect 3324 8496 3332 8504
rect 5132 8496 5140 8504
rect 5276 8496 5284 8504
rect 7240 8496 7248 8504
rect 9036 8496 9044 8504
rect 9820 8496 9828 8504
rect 11772 8496 11780 8504
rect 684 8476 692 8484
rect 3836 8476 3844 8484
rect 7740 8476 7748 8484
rect 7868 8476 7876 8484
rect 11036 8476 11044 8484
rect 1884 8436 1892 8444
rect 5276 8436 5284 8444
rect 5918 8436 5926 8444
rect 10476 8436 10484 8444
rect 11772 8436 11780 8444
rect 732 8376 740 8384
rect 1884 8376 1892 8384
rect 1996 8376 2004 8384
rect 3180 8376 3188 8384
rect 3228 8376 3236 8384
rect 3980 8376 3988 8384
rect 5196 8376 5204 8384
rect 5276 8376 5284 8384
rect 5918 8376 5926 8384
rect 7132 8376 7140 8384
rect 7228 8376 7236 8384
rect 9068 8376 9076 8384
rect 9708 8376 9716 8384
rect 9788 8376 9796 8384
rect 10476 8376 10484 8384
rect 11772 8376 11780 8384
rect 668 8356 676 8364
rect 2028 8356 2036 8364
rect 3932 8356 3940 8364
rect 7820 8356 7828 8364
rect 1372 8336 1380 8344
rect 5788 8336 5796 8344
rect 7868 8336 7876 8344
rect 9036 8336 9044 8344
rect 9820 8336 9828 8344
rect 10988 8336 10996 8344
rect 11004 8336 11012 8344
rect 11036 8336 11044 8344
rect 1884 8316 1892 8324
rect 3836 8316 3844 8324
rect 3900 8316 3908 8324
rect 5276 8316 5284 8324
rect 6508 8316 6516 8324
rect 8524 8316 8532 8324
rect 10332 8316 10340 8324
rect 11676 8316 11684 8324
rect 1964 8296 1972 8304
rect 4556 8296 4564 8304
rect 6492 8296 6500 8304
rect 11692 8296 11700 8304
rect 1964 8276 1972 8284
rect 3916 8276 3924 8284
rect 11692 8276 11700 8284
rect 12268 8276 12276 8284
rect 44 8236 52 8244
rect 12332 8236 12340 8244
rect 2572 8176 2580 8184
rect 5180 8176 5188 8184
rect 5244 8176 5252 8184
rect 8428 8176 8436 8184
rect 9068 8176 9076 8184
rect 9724 8176 9732 8184
rect 11628 8176 11636 8184
rect 11676 8176 11684 8184
rect 2524 8136 2532 8144
rect 2684 8136 2692 8144
rect 4540 8136 4548 8144
rect 5116 8136 5124 8144
rect 5292 8136 5300 8144
rect 5932 8136 5940 8144
rect 6588 8136 6596 8144
rect 9020 8136 9028 8144
rect 11788 8136 11796 8144
rect 732 8116 740 8124
rect 1868 8116 1876 8124
rect 3820 8116 3828 8124
rect 4476 8116 4484 8124
rect 6540 8116 6548 8124
rect 7788 8116 7796 8124
rect 9772 8116 9780 8124
rect 76 8096 84 8104
rect 1212 8096 1220 8104
rect 3900 8096 3908 8104
rect 4620 8096 4628 8104
rect 8524 8096 8532 8104
rect 10332 8096 10340 8104
rect 11020 8096 11028 8104
rect 11036 8096 11044 8104
rect 12284 8096 12292 8104
rect 572 8076 580 8084
rect 1948 8076 1956 8084
rect 7740 8076 7748 8084
rect 10988 8076 10996 8084
rect 4620 8036 4628 8044
rect 7868 8036 7876 8044
rect 12284 8036 12292 8044
rect 700 7976 708 7984
rect 732 7976 740 7984
rect 2620 7976 2628 7984
rect 2636 7976 2644 7984
rect 4476 7976 4484 7984
rect 4620 7976 4628 7984
rect 6428 7976 6436 7984
rect 7116 7976 7124 7984
rect 7868 7976 7876 7984
rect 8380 7976 8388 7984
rect 8428 7976 8436 7984
rect 9676 7976 9684 7984
rect 10380 7976 10388 7984
rect 12284 7976 12292 7984
rect 1340 7956 1348 7964
rect 10380 7956 10388 7964
rect 1372 7936 1380 7944
rect 2684 7936 2692 7944
rect 3324 7936 3332 7944
rect 10316 7936 10324 7944
rect 1820 7916 1828 7924
rect 4044 7916 4052 7924
rect 4620 7916 4628 7924
rect 5276 7916 5284 7924
rect 7724 7916 7732 7924
rect 12284 7916 12292 7924
rect 92 7876 100 7884
rect 6492 7876 6500 7884
rect 5820 7836 5828 7844
rect 7180 7836 7188 7844
rect 11628 7836 11636 7844
rect 11660 7836 11668 7844
rect 11740 7836 11748 7844
rect 1260 7776 1268 7784
rect 2636 7776 2644 7784
rect 4476 7776 4484 7784
rect 4508 7776 4516 7784
rect 5228 7776 5236 7784
rect 8428 7776 8436 7784
rect 9068 7776 9076 7784
rect 9676 7776 9684 7784
rect 9740 7776 9748 7784
rect 11020 7776 11028 7784
rect 12 7756 20 7764
rect 2028 7756 2036 7764
rect 5278 7756 5286 7764
rect 92 7736 100 7744
rect 1388 7736 1396 7744
rect 2684 7736 2692 7744
rect 4636 7736 4644 7744
rect 5212 7736 5220 7744
rect 9020 7736 9028 7744
rect 10316 7736 10324 7744
rect 12268 7736 12276 7744
rect 7068 7716 7076 7724
rect 7788 7716 7796 7724
rect 8380 7716 8388 7724
rect 1884 7696 1892 7704
rect 2524 7696 2532 7704
rect 3168 7696 3176 7704
rect 3996 7696 4004 7704
rect 5132 7696 5140 7704
rect 7148 7696 7156 7704
rect 8524 7696 8532 7704
rect 9084 7696 9092 7704
rect 9884 7696 9892 7704
rect 10396 7696 10404 7704
rect 10476 7696 10484 7704
rect 3324 7676 3332 7684
rect 4524 7676 4532 7684
rect 7740 7676 7748 7684
rect 2540 7636 2548 7644
rect 5788 7636 5796 7644
rect 5884 7636 5892 7644
rect 7868 7636 7876 7644
rect 9820 7636 9828 7644
rect 10476 7636 10484 7644
rect 11100 7636 11108 7644
rect 11772 7636 11780 7644
rect 1228 7576 1236 7584
rect 1276 7576 1284 7584
rect 1996 7576 2004 7584
rect 2028 7576 2036 7584
rect 2540 7576 2548 7584
rect 3180 7576 3188 7584
rect 4476 7576 4484 7584
rect 5164 7576 5172 7584
rect 5180 7576 5188 7584
rect 5788 7576 5796 7584
rect 6540 7576 6548 7584
rect 7868 7576 7876 7584
rect 8380 7576 8388 7584
rect 8428 7576 8436 7584
rect 9820 7576 9828 7584
rect 10476 7576 10484 7584
rect 11036 7576 11044 7584
rect 11772 7576 11780 7584
rect 7180 7556 7188 7564
rect 7228 7556 7236 7564
rect 8492 7556 8500 7564
rect 588 7536 596 7544
rect 1980 7536 1988 7544
rect 3836 7536 3844 7544
rect 5276 7536 5284 7544
rect 11644 7536 11652 7544
rect 1372 7516 1380 7524
rect 1932 7516 1940 7524
rect 3324 7516 3332 7524
rect 3996 7516 4004 7524
rect 4620 7516 4628 7524
rect 7084 7516 7092 7524
rect 10476 7516 10484 7524
rect 11772 7516 11780 7524
rect 1292 7496 1300 7504
rect 3244 7496 3252 7504
rect 8540 7496 8548 7504
rect 9676 7496 9684 7504
rect 9740 7496 9748 7504
rect 2028 7476 2036 7484
rect 7164 7476 7172 7484
rect 11692 7476 11700 7484
rect 6428 7436 6436 7444
rect 6460 7436 6468 7444
rect 10364 7436 10372 7444
rect 12316 7436 12324 7444
rect 28 7376 36 7384
rect 700 7376 708 7384
rect 732 7376 740 7384
rect 1996 7376 2004 7384
rect 2028 7376 2036 7384
rect 4524 7376 4532 7384
rect 7228 7376 7236 7384
rect 8380 7376 8388 7384
rect 8412 7376 8420 7384
rect 9084 7376 9092 7384
rect 11100 7376 11108 7384
rect 11132 7376 11140 7384
rect 1340 7356 1348 7364
rect 4540 7356 4548 7364
rect 9772 7356 9780 7364
rect 1388 7336 1396 7344
rect 2684 7336 2692 7344
rect 5340 7336 5348 7344
rect 7068 7336 7076 7344
rect 9020 7336 9028 7344
rect 12268 7336 12276 7344
rect 3820 7316 3828 7324
rect 5212 7316 5220 7324
rect 1884 7296 1892 7304
rect 3116 7296 3124 7304
rect 3168 7296 3176 7304
rect 5132 7296 5140 7304
rect 6572 7296 6580 7304
rect 7660 7296 7668 7304
rect 10332 7296 10340 7304
rect 10476 7296 10484 7304
rect 11772 7296 11780 7304
rect 3884 7276 3892 7284
rect 5276 7276 5284 7284
rect 9804 7276 9812 7284
rect 9676 7256 9684 7264
rect 1884 7236 1892 7244
rect 2540 7236 2548 7244
rect 5132 7236 5140 7244
rect 5868 7236 5876 7244
rect 8524 7236 8532 7244
rect 10476 7236 10484 7244
rect 11020 7236 11028 7244
rect 11772 7236 11780 7244
rect 700 7176 708 7184
rect 1340 7176 1348 7184
rect 1884 7176 1892 7184
rect 2028 7176 2036 7184
rect 2540 7176 2548 7184
rect 3980 7176 3988 7184
rect 4588 7176 4596 7184
rect 5132 7176 5140 7184
rect 5932 7176 5940 7184
rect 7836 7176 7844 7184
rect 8524 7176 8532 7184
rect 9724 7176 9732 7184
rect 10476 7176 10484 7184
rect 11772 7176 11780 7184
rect 1964 7156 1972 7164
rect 5836 7156 5844 7164
rect 572 7136 580 7144
rect 1372 7136 1380 7144
rect 4620 7136 4628 7144
rect 5804 7136 5812 7144
rect 7740 7136 7748 7144
rect 7884 7136 7892 7144
rect 9100 7136 9108 7144
rect 9692 7136 9700 7144
rect 10332 7136 10340 7144
rect 10988 7136 10996 7144
rect 11644 7136 11652 7144
rect 76 7116 84 7124
rect 1884 7116 1892 7124
rect 2460 7116 2468 7124
rect 6508 7116 6516 7124
rect 7084 7116 7092 7124
rect 10476 7116 10484 7124
rect 11772 7116 11780 7124
rect 3340 7096 3348 7104
rect 6588 7096 6596 7104
rect 9020 7096 9028 7104
rect 2684 7076 2692 7084
rect 11692 7076 11700 7084
rect 12268 7076 12276 7084
rect 2620 7036 2628 7044
rect 10380 7036 10388 7044
rect 12332 7036 12340 7044
rect 700 6976 708 6984
rect 3932 6976 3940 6984
rect 5180 6976 5188 6984
rect 6476 6976 6484 6984
rect 7788 6976 7796 6984
rect 10396 6976 10404 6984
rect 11676 6976 11684 6984
rect 11708 6976 11716 6984
rect 7820 6956 7828 6964
rect 1388 6936 1396 6944
rect 2588 6936 2596 6944
rect 3244 6936 3252 6944
rect 5772 6936 5780 6944
rect 6492 6936 6500 6944
rect 10316 6936 10324 6944
rect 10972 6936 10980 6944
rect 2588 6916 2596 6924
rect 3820 6916 3828 6924
rect 7068 6916 7076 6924
rect 9020 6916 9028 6924
rect 1324 6896 1332 6904
rect 1884 6896 1892 6904
rect 3324 6896 3332 6904
rect 4620 6896 4628 6904
rect 5276 6896 5284 6904
rect 9100 6896 9108 6904
rect 9884 6896 9892 6904
rect 11036 6896 11044 6904
rect 92 6876 100 6884
rect 2540 6876 2548 6884
rect 3196 6876 3204 6884
rect 7148 6876 7156 6884
rect 9740 6876 9748 6884
rect 2668 6836 2676 6844
rect 3324 6836 3332 6844
rect 4620 6836 4628 6844
rect 5276 6836 5284 6844
rect 8524 6836 8532 6844
rect 10476 6836 10484 6844
rect 12284 6836 12292 6844
rect 620 6776 628 6784
rect 2572 6776 2580 6784
rect 2668 6776 2676 6784
rect 3324 6776 3332 6784
rect 4476 6776 4484 6784
rect 4508 6776 4516 6784
rect 4620 6776 4628 6784
rect 5276 6776 5284 6784
rect 5900 6776 5908 6784
rect 8380 6776 8388 6784
rect 8524 6776 8532 6784
rect 9708 6776 9716 6784
rect 10476 6776 10484 6784
rect 11036 6776 11044 6784
rect 11740 6776 11748 6784
rect 12284 6776 12292 6784
rect 3180 6756 3188 6764
rect 6540 6756 6548 6764
rect 11628 6756 11636 6764
rect 1948 6736 1956 6744
rect 5948 6736 5956 6744
rect 6572 6736 6580 6744
rect 7724 6736 7732 6744
rect 9100 6736 9108 6744
rect 10988 6736 10996 6744
rect 11788 6736 11796 6744
rect 12924 6736 12932 6744
rect 76 6716 84 6724
rect 3868 6716 3876 6724
rect 5276 6716 5284 6724
rect 8524 6716 8532 6724
rect 10396 6716 10404 6724
rect 10476 6716 10484 6724
rect 11036 6716 11044 6724
rect 11196 6716 11204 6724
rect 1868 6696 1876 6704
rect 3820 6696 3828 6704
rect 5116 6696 5124 6704
rect 9020 6696 9028 6704
rect 10316 6696 10324 6704
rect 8444 6676 8452 6684
rect 10396 6676 10404 6684
rect 732 6636 740 6644
rect 11660 6636 11668 6644
rect 2028 6576 2036 6584
rect 4524 6576 4532 6584
rect 8460 6576 8468 6584
rect 12316 6576 12324 6584
rect 1340 6556 1348 6564
rect 9132 6556 9140 6564
rect 1388 6536 1396 6544
rect 1964 6536 1972 6544
rect 6492 6536 6500 6544
rect 7836 6536 7844 6544
rect 7884 6536 7892 6544
rect 9116 6536 9124 6544
rect 11132 6536 11140 6544
rect 3820 6516 3828 6524
rect 5772 6516 5780 6524
rect 9180 6516 9188 6524
rect 11068 6516 11076 6524
rect 76 6496 84 6504
rect 1884 6496 1892 6504
rect 2524 6496 2532 6504
rect 3324 6496 3332 6504
rect 4572 6496 4580 6504
rect 5132 6496 5140 6504
rect 5340 6496 5348 6504
rect 6572 6496 6580 6504
rect 8316 6496 8324 6504
rect 10332 6496 10340 6504
rect 3244 6476 3252 6484
rect 3900 6476 3908 6484
rect 5852 6476 5860 6484
rect 7084 6476 7092 6484
rect 9820 6476 9828 6484
rect 10460 6476 10468 6484
rect 620 6436 628 6444
rect 684 6436 692 6444
rect 1884 6436 1892 6444
rect 2668 6436 2676 6444
rect 5276 6436 5284 6444
rect 5918 6436 5926 6444
rect 6428 6436 6436 6444
rect 6460 6436 6468 6444
rect 7180 6436 7188 6444
rect 44 6376 52 6384
rect 732 6376 740 6384
rect 1884 6376 1892 6384
rect 2668 6376 2676 6384
rect 3292 6376 3300 6384
rect 5276 6376 5284 6384
rect 5918 6376 5926 6384
rect 6428 6376 6436 6384
rect 6476 6376 6484 6384
rect 7820 6376 7828 6384
rect 11724 6376 11732 6384
rect 668 6356 676 6364
rect 76 6336 84 6344
rect 1372 6336 1380 6344
rect 4524 6336 4532 6344
rect 5788 6336 5796 6344
rect 8524 6336 8532 6344
rect 9692 6336 9700 6344
rect 10332 6336 10340 6344
rect 10988 6336 10996 6344
rect 11788 6336 11796 6344
rect 1820 6316 1828 6324
rect 2092 6316 2100 6324
rect 2748 6316 2756 6324
rect 3996 6316 4004 6324
rect 5132 6316 5140 6324
rect 5276 6316 5284 6324
rect 7084 6316 7092 6324
rect 7820 6316 7828 6324
rect 10476 6316 10484 6324
rect 12284 6316 12292 6324
rect 9740 6296 9748 6304
rect 10396 6296 10404 6304
rect 2508 6276 2516 6284
rect 2588 6276 2596 6284
rect 6588 6276 6596 6284
rect 2572 6236 2580 6244
rect 3180 6236 3188 6244
rect 4524 6236 4532 6244
rect 6476 6236 6484 6244
rect 44 6176 52 6184
rect 2028 6176 2036 6184
rect 3868 6176 3876 6184
rect 5164 6176 5172 6184
rect 5244 6176 5252 6184
rect 7116 6176 7124 6184
rect 7228 6176 7236 6184
rect 9084 6176 9092 6184
rect 9180 6176 9188 6184
rect 12316 6176 12324 6184
rect 1964 6156 1972 6164
rect 2620 6156 2628 6164
rect 5932 6156 5940 6164
rect 92 6136 100 6144
rect 684 6136 692 6144
rect 2684 6136 2692 6144
rect 3820 6136 3828 6144
rect 5292 6136 5300 6144
rect 7068 6136 7076 6144
rect 9020 6136 9028 6144
rect 9836 6136 9844 6144
rect 4540 6116 4548 6124
rect 10972 6116 10980 6124
rect 11692 6116 11700 6124
rect 1324 6096 1332 6104
rect 1884 6096 1892 6104
rect 3168 6096 3176 6104
rect 4044 6096 4052 6104
rect 8524 6096 8532 6104
rect 1340 6076 1348 6084
rect 4556 6076 4564 6084
rect 7868 6076 7876 6084
rect 11036 6076 11044 6084
rect 588 6036 596 6044
rect 1884 6036 1892 6044
rect 6572 6036 6580 6044
rect 7836 6036 7844 6044
rect 10476 6036 10484 6044
rect 11772 6036 11780 6044
rect 44 5976 52 5984
rect 588 5976 596 5984
rect 1884 5976 1892 5984
rect 2588 5976 2596 5984
rect 3260 5976 3268 5984
rect 6572 5976 6580 5984
rect 7148 5976 7156 5984
rect 8412 5976 8420 5984
rect 8476 5976 8484 5984
rect 9676 5976 9684 5984
rect 10476 5976 10484 5984
rect 11772 5976 11780 5984
rect 92 5936 100 5944
rect 1388 5936 1396 5944
rect 3324 5936 3332 5944
rect 4636 5936 4644 5944
rect 5788 5936 5796 5944
rect 6444 5936 6452 5944
rect 7740 5936 7748 5944
rect 10988 5936 10996 5944
rect 11644 5936 11652 5944
rect 2040 5916 2048 5924
rect 4044 5916 4052 5924
rect 5132 5916 5140 5924
rect 5276 5916 5284 5924
rect 6492 5916 6500 5924
rect 10396 5916 10404 5924
rect 11772 5916 11780 5924
rect 1324 5896 1332 5904
rect 6460 5896 6468 5904
rect 7788 5896 7796 5904
rect 9740 5896 9748 5904
rect 2588 5876 2596 5884
rect 5836 5876 5844 5884
rect 7788 5876 7796 5884
rect 8556 5876 8564 5884
rect 10316 5876 10324 5884
rect 12268 5876 12276 5884
rect 4476 5836 4484 5844
rect 5820 5836 5828 5844
rect 8444 5836 8452 5844
rect 12316 5836 12324 5844
rect 700 5776 708 5784
rect 732 5776 740 5784
rect 1324 5776 1332 5784
rect 3276 5776 3284 5784
rect 3948 5776 3956 5784
rect 6476 5776 6484 5784
rect 6492 5776 6500 5784
rect 8380 5776 8388 5784
rect 11692 5776 11700 5784
rect 5278 5756 5286 5764
rect 7180 5756 7188 5764
rect 1388 5736 1396 5744
rect 2684 5736 2692 5744
rect 4636 5736 4644 5744
rect 5228 5736 5236 5744
rect 6588 5736 6596 5744
rect 7164 5736 7172 5744
rect 10316 5736 10324 5744
rect 12364 5736 12372 5744
rect 5212 5716 5220 5724
rect 10972 5716 10980 5724
rect 3836 5696 3844 5704
rect 5132 5696 5140 5704
rect 7084 5696 7092 5704
rect 7724 5696 7732 5704
rect 8524 5696 8532 5704
rect 10540 5696 10548 5704
rect 12284 5696 12292 5704
rect 9020 5676 9028 5684
rect 9740 5676 9748 5684
rect 11052 5676 11060 5684
rect 44 5636 52 5644
rect 1884 5636 1892 5644
rect 1980 5636 1988 5644
rect 2540 5636 2548 5644
rect 3836 5636 3844 5644
rect 5788 5636 5796 5644
rect 7084 5636 7092 5644
rect 7740 5636 7748 5644
rect 8524 5636 8532 5644
rect 9068 5636 9076 5644
rect 10476 5636 10484 5644
rect 11740 5636 11748 5644
rect 732 5576 740 5584
rect 1324 5576 1332 5584
rect 1884 5576 1892 5584
rect 2028 5576 2036 5584
rect 2540 5576 2548 5584
rect 3836 5576 3844 5584
rect 3948 5576 3956 5584
rect 5180 5576 5188 5584
rect 5788 5576 5796 5584
rect 7084 5576 7092 5584
rect 7740 5576 7748 5584
rect 8524 5576 8532 5584
rect 9084 5576 9092 5584
rect 10476 5576 10484 5584
rect 12 5556 20 5564
rect 2636 5556 2644 5564
rect 7228 5556 7236 5564
rect 12972 5556 12980 5564
rect 76 5536 84 5544
rect 1372 5536 1380 5544
rect 2684 5536 2692 5544
rect 5132 5536 5140 5544
rect 5276 5536 5284 5544
rect 5852 5536 5860 5544
rect 10988 5536 10996 5544
rect 12284 5536 12292 5544
rect 1884 5516 1892 5524
rect 3836 5516 3844 5524
rect 4556 5516 4564 5524
rect 7084 5516 7092 5524
rect 7948 5516 7956 5524
rect 8444 5516 8452 5524
rect 8524 5516 8532 5524
rect 10332 5516 10340 5524
rect 7164 5496 7172 5504
rect 11708 5496 11716 5504
rect 3340 5476 3348 5484
rect 8380 5476 8388 5484
rect 8412 5436 8420 5444
rect 9676 5436 9684 5444
rect 9724 5436 9732 5444
rect 11100 5436 11108 5444
rect 11132 5436 11140 5444
rect 620 5376 628 5384
rect 732 5376 740 5384
rect 1964 5376 1972 5384
rect 3980 5376 3988 5384
rect 5820 5376 5828 5384
rect 6460 5376 6468 5384
rect 6476 5376 6484 5384
rect 7804 5376 7812 5384
rect 8476 5376 8484 5384
rect 11036 5376 11044 5384
rect 9788 5356 9796 5364
rect 572 5336 580 5344
rect 1388 5336 1396 5344
rect 3388 5336 3396 5344
rect 5772 5336 5780 5344
rect 6588 5336 6596 5344
rect 9116 5336 9124 5344
rect 9836 5336 9844 5344
rect 3916 5316 3924 5324
rect 5116 5316 5124 5324
rect 12268 5316 12276 5324
rect 76 5296 84 5304
rect 1884 5296 1892 5304
rect 3836 5296 3844 5304
rect 4684 5296 4692 5304
rect 7084 5296 7092 5304
rect 9772 5296 9780 5304
rect 10268 5296 10276 5304
rect 10540 5296 10548 5304
rect 684 5276 692 5284
rect 5836 5276 5844 5284
rect 7740 5276 7748 5284
rect 10988 5276 10996 5284
rect 12348 5276 12356 5284
rect 12924 5276 12932 5284
rect 9116 5256 9124 5264
rect 76 5236 84 5244
rect 1884 5236 1892 5244
rect 2540 5236 2548 5244
rect 3212 5236 3220 5244
rect 4620 5236 4628 5244
rect 5276 5236 5284 5244
rect 9036 5236 9044 5244
rect 9180 5236 9188 5244
rect 10476 5236 10484 5244
rect 12972 5236 12980 5244
rect 76 5176 84 5184
rect 636 5176 644 5184
rect 732 5176 740 5184
rect 1884 5176 1892 5184
rect 2028 5176 2036 5184
rect 2540 5176 2548 5184
rect 3884 5176 3892 5184
rect 4476 5176 4484 5184
rect 4508 5176 4516 5184
rect 4620 5176 4628 5184
rect 5276 5176 5284 5184
rect 5932 5176 5940 5184
rect 9036 5176 9044 5184
rect 10476 5176 10484 5184
rect 11740 5176 11748 5184
rect 636 5156 644 5164
rect 9788 5156 9796 5164
rect 588 5136 596 5144
rect 2012 5136 2020 5144
rect 7148 5136 7156 5144
rect 9820 5136 9828 5144
rect 10988 5136 10996 5144
rect 3228 5116 3236 5124
rect 3324 5116 3332 5124
rect 3996 5116 4004 5124
rect 5276 5116 5284 5124
rect 9772 5116 9780 5124
rect 11724 5116 11732 5124
rect 12284 5116 12292 5124
rect 3180 5096 3188 5104
rect 5868 5096 5876 5104
rect 7068 5096 7076 5104
rect 1388 5076 1396 5084
rect 3244 5076 3252 5084
rect 3820 5076 3828 5084
rect 4540 5076 4548 5084
rect 5116 5076 5124 5084
rect 7724 5076 7732 5084
rect 12364 5076 12372 5084
rect 3868 5036 3876 5044
rect 5836 5036 5844 5044
rect 7772 5036 7780 5044
rect 8380 5036 8388 5044
rect 8492 5036 8500 5044
rect 9116 5036 9124 5044
rect 44 4976 52 4984
rect 3260 4976 3268 4984
rect 3980 4976 3988 4984
rect 4588 4976 4596 4984
rect 7132 4976 7140 4984
rect 9068 4976 9076 4984
rect 12972 4976 12980 4984
rect 6476 4956 6484 4964
rect 732 4936 740 4944
rect 1388 4936 1396 4944
rect 2028 4936 2036 4944
rect 2636 4936 2644 4944
rect 4636 4936 4644 4944
rect 6492 4936 6500 4944
rect 9740 4936 9748 4944
rect 11628 4936 11636 4944
rect 12876 4936 12884 4944
rect 1340 4916 1348 4924
rect 2684 4916 2692 4924
rect 3916 4916 3924 4924
rect 5772 4916 5780 4924
rect 8380 4916 8388 4924
rect 1884 4896 1892 4904
rect 3116 4896 3124 4904
rect 3168 4896 3176 4904
rect 5132 4896 5140 4904
rect 5852 4896 5860 4904
rect 6572 4896 6580 4904
rect 8524 4896 8532 4904
rect 10476 4896 10484 4904
rect 11196 4896 11204 4904
rect 11692 4896 11700 4904
rect 2684 4876 2692 4884
rect 6444 4876 6452 4884
rect 10396 4876 10404 4884
rect 11628 4856 11636 4864
rect 1884 4836 1892 4844
rect 5918 4836 5926 4844
rect 7132 4836 7140 4844
rect 7740 4836 7748 4844
rect 8524 4836 8532 4844
rect 9708 4836 9716 4844
rect 11020 4836 11028 4844
rect 11660 4836 11668 4844
rect 12316 4836 12324 4844
rect 700 4776 708 4784
rect 1884 4776 1892 4784
rect 3948 4776 3956 4784
rect 5164 4776 5172 4784
rect 5918 4776 5926 4784
rect 6540 4776 6548 4784
rect 7180 4776 7188 4784
rect 7740 4776 7748 4784
rect 7836 4776 7844 4784
rect 8524 4776 8532 4784
rect 9788 4776 9796 4784
rect 11628 4776 11636 4784
rect 11676 4776 11684 4784
rect 5196 4756 5204 4764
rect 10428 4756 10436 4764
rect 92 4736 100 4744
rect 1308 4736 1316 4744
rect 2540 4736 2548 4744
rect 2684 4736 2692 4744
rect 3836 4736 3844 4744
rect 7212 4736 7220 4744
rect 9820 4736 9828 4744
rect 10476 4736 10484 4744
rect 1884 4716 1892 4724
rect 3324 4716 3332 4724
rect 4620 4716 4628 4724
rect 7084 4716 7092 4724
rect 8588 4716 8596 4724
rect 10332 4716 10340 4724
rect 12284 4716 12292 4724
rect 1388 4696 1396 4704
rect 10412 4696 10420 4704
rect 11724 4696 11732 4704
rect 12364 4696 12372 4704
rect 5100 4676 5108 4684
rect 7164 4676 7172 4684
rect 9020 4676 9028 4684
rect 6428 4636 6436 4644
rect 6460 4636 6468 4644
rect 9724 4636 9732 4644
rect 2028 4576 2036 4584
rect 5820 4576 5828 4584
rect 5836 4576 5844 4584
rect 7116 4576 7124 4584
rect 7820 4576 7828 4584
rect 9180 4576 9188 4584
rect 9772 4576 9780 4584
rect 11052 4576 11060 4584
rect 11740 4576 11748 4584
rect 12 4556 20 4564
rect 7228 4556 7236 4564
rect 9084 4556 9092 4564
rect 92 4536 100 4544
rect 732 4536 740 4544
rect 4540 4536 4548 4544
rect 7884 4536 7892 4544
rect 9020 4536 9028 4544
rect 9836 4536 9844 4544
rect 12364 4536 12372 4544
rect 3820 4516 3828 4524
rect 5196 4516 5204 4524
rect 1212 4496 1220 4504
rect 1884 4496 1892 4504
rect 3324 4496 3332 4504
rect 5276 4496 5284 4504
rect 6572 4496 6580 4504
rect 9772 4496 9780 4504
rect 10476 4496 10484 4504
rect 12284 4496 12292 4504
rect 4492 4476 4500 4484
rect 588 4436 596 4444
rect 1340 4436 1348 4444
rect 1884 4436 1892 4444
rect 2540 4436 2548 4444
rect 3228 4436 3236 4444
rect 3324 4436 3332 4444
rect 4508 4436 4516 4444
rect 5164 4436 5172 4444
rect 6572 4436 6580 4444
rect 10476 4436 10484 4444
rect 11020 4436 11028 4444
rect 44 4376 52 4384
rect 588 4376 596 4384
rect 732 4376 740 4384
rect 1340 4376 1348 4384
rect 1884 4376 1892 4384
rect 2028 4376 2036 4384
rect 2540 4376 2548 4384
rect 2620 4376 2628 4384
rect 3324 4376 3332 4384
rect 3868 4376 3876 4384
rect 3980 4376 3988 4384
rect 5244 4376 5252 4384
rect 5884 4376 5892 4384
rect 6572 4376 6580 4384
rect 8380 4376 8388 4384
rect 8412 4376 8420 4384
rect 9180 4376 9188 4384
rect 10476 4376 10484 4384
rect 11628 4376 11636 4384
rect 11660 4376 11668 4384
rect 3884 4356 3892 4364
rect 9132 4356 9140 4364
rect 76 4336 84 4344
rect 2684 4336 2692 4344
rect 4604 4336 4612 4344
rect 7724 4336 7732 4344
rect 9820 4336 9828 4344
rect 12348 4336 12356 4344
rect 1884 4316 1892 4324
rect 2460 4316 2468 4324
rect 3116 4316 3124 4324
rect 3324 4316 3332 4324
rect 5132 4316 5140 4324
rect 6364 4316 6372 4324
rect 6412 4316 6420 4324
rect 9036 4316 9044 4324
rect 9100 4316 9108 4324
rect 10332 4316 10340 4324
rect 10476 4316 10484 4324
rect 11708 4316 11716 4324
rect 7788 4296 7796 4304
rect 9116 4296 9124 4304
rect 11692 4296 11700 4304
rect 7068 4276 7076 4284
rect 11036 4276 11044 4284
rect 8492 4256 8500 4264
rect 11020 4236 11028 4244
rect 12972 4236 12980 4244
rect 44 4176 52 4184
rect 1964 4176 1972 4184
rect 2028 4176 2036 4184
rect 3180 4176 3188 4184
rect 4476 4176 4484 4184
rect 4508 4176 4516 4184
rect 4524 4176 4532 4184
rect 5820 4176 5828 4184
rect 7116 4176 7124 4184
rect 9708 4176 9716 4184
rect 10364 4176 10372 4184
rect 10444 4176 10452 4184
rect 12396 4176 12404 4184
rect 12428 4176 12436 4184
rect 1340 4156 1348 4164
rect 5932 4156 5940 4164
rect 11628 4156 11636 4164
rect 1388 4136 1396 4144
rect 3244 4136 3252 4144
rect 5772 4136 5780 4144
rect 7068 4136 7076 4144
rect 8444 4136 8452 4144
rect 9020 4136 9028 4144
rect 9740 4136 9748 4144
rect 10316 4136 10324 4144
rect 10492 4136 10500 4144
rect 11676 4136 11684 4144
rect 11788 4136 11796 4144
rect 12364 4136 12372 4144
rect 3820 4116 3828 4124
rect 7724 4116 7732 4124
rect 2524 4096 2532 4104
rect 3324 4096 3332 4104
rect 5132 4096 5140 4104
rect 6636 4096 6644 4104
rect 12284 4096 12292 4104
rect 7788 4076 7796 4084
rect 11724 4076 11732 4084
rect 684 4056 692 4064
rect 1884 4036 1892 4044
rect 3180 4036 3188 4044
rect 5276 4036 5284 4044
rect 6572 4036 6580 4044
rect 8412 4036 8420 4044
rect 10988 4036 10996 4044
rect 12940 4036 12948 4044
rect 620 3976 628 3984
rect 1228 3976 1236 3984
rect 1884 3976 1892 3984
rect 2636 3976 2644 3984
rect 3292 3976 3300 3984
rect 4508 3976 4516 3984
rect 5276 3976 5284 3984
rect 5868 3976 5876 3984
rect 5900 3976 5908 3984
rect 6572 3976 6580 3984
rect 7116 3976 7124 3984
rect 7788 3976 7796 3984
rect 10988 3976 10996 3984
rect 11084 3976 11092 3984
rect 12396 3976 12404 3984
rect 12940 3976 12948 3984
rect 9132 3956 9140 3964
rect 9788 3956 9796 3964
rect 572 3936 580 3944
rect 1372 3936 1380 3944
rect 3340 3936 3348 3944
rect 5212 3936 5220 3944
rect 7084 3936 7092 3944
rect 7740 3936 7748 3944
rect 8460 3936 8468 3944
rect 12300 3936 12308 3944
rect 76 3916 84 3924
rect 1884 3916 1892 3924
rect 5276 3916 5284 3924
rect 6572 3916 6580 3924
rect 6636 3916 6644 3924
rect 11612 3916 11620 3924
rect 11836 3916 11844 3924
rect 5116 3896 5124 3904
rect 8540 3896 8548 3904
rect 9116 3896 9124 3904
rect 9836 3896 9844 3904
rect 9996 3896 10004 3904
rect 11708 3896 11716 3904
rect 2508 3876 2516 3884
rect 10412 3876 10420 3884
rect 10492 3876 10500 3884
rect 12268 3876 12276 3884
rect 9996 3856 10004 3864
rect 5932 3836 5940 3844
rect 10428 3836 10436 3844
rect 12364 3836 12372 3844
rect 44 3776 52 3784
rect 2620 3776 2628 3784
rect 3868 3776 3876 3784
rect 4540 3776 4548 3784
rect 5164 3776 5172 3784
rect 6428 3776 6436 3784
rect 6460 3776 6468 3784
rect 7772 3776 7780 3784
rect 8380 3776 8388 3784
rect 8412 3776 8420 3784
rect 9180 3776 9188 3784
rect 11628 3776 11636 3784
rect 11660 3776 11668 3784
rect 11740 3776 11748 3784
rect 92 3736 100 3744
rect 3820 3736 3828 3744
rect 6492 3736 6500 3744
rect 8444 3736 8452 3744
rect 8636 3736 8644 3744
rect 1372 3696 1380 3704
rect 3168 3696 3176 3704
rect 3324 3696 3332 3704
rect 3900 3696 3908 3704
rect 4620 3696 4628 3704
rect 7948 3696 7956 3704
rect 8524 3696 8532 3704
rect 10476 3696 10484 3704
rect 12284 3696 12292 3704
rect 1244 3676 1252 3684
rect 1948 3676 1956 3684
rect 7068 3676 7076 3684
rect 7724 3676 7732 3684
rect 9020 3676 9028 3684
rect 10332 3676 10340 3684
rect 10988 3676 10996 3684
rect 2588 3656 2596 3664
rect 5196 3636 5204 3644
rect 5918 3636 5926 3644
rect 7868 3636 7876 3644
rect 8524 3636 8532 3644
rect 9068 3636 9076 3644
rect 10476 3636 10484 3644
rect 12284 3636 12292 3644
rect 12380 3636 12388 3644
rect 12428 3636 12436 3644
rect 636 3576 644 3584
rect 2604 3576 2612 3584
rect 4476 3576 4484 3584
rect 5180 3576 5188 3584
rect 5836 3576 5844 3584
rect 5918 3576 5926 3584
rect 7868 3576 7876 3584
rect 8524 3576 8532 3584
rect 10476 3576 10484 3584
rect 12284 3576 12292 3584
rect 572 3536 580 3544
rect 1372 3536 1380 3544
rect 2668 3536 2676 3544
rect 5116 3536 5124 3544
rect 10988 3536 10996 3544
rect 76 3516 84 3524
rect 3900 3516 3908 3524
rect 4684 3516 4692 3524
rect 5180 3516 5188 3524
rect 6492 3516 6500 3524
rect 6572 3516 6580 3524
rect 7804 3516 7812 3524
rect 8524 3516 8532 3524
rect 10332 3516 10340 3524
rect 10540 3516 10548 3524
rect 12284 3516 12292 3524
rect 6428 3496 6436 3504
rect 8380 3496 8388 3504
rect 8444 3496 8452 3504
rect 2524 3476 2532 3484
rect 4540 3476 4548 3484
rect 6492 3476 6500 3484
rect 7724 3476 7732 3484
rect 9084 3476 9092 3484
rect 11788 3476 11796 3484
rect 12364 3476 12372 3484
rect 9676 3456 9684 3464
rect 3292 3436 3300 3444
rect 7132 3436 7140 3444
rect 9708 3436 9716 3444
rect 9788 3436 9796 3444
rect 11628 3436 11636 3444
rect 11740 3436 11748 3444
rect 44 3376 52 3384
rect 3916 3376 3924 3384
rect 3932 3376 3940 3384
rect 3980 3376 3988 3384
rect 5868 3376 5876 3384
rect 10380 3376 10388 3384
rect 12972 3376 12980 3384
rect 2028 3356 2036 3364
rect 9132 3356 9140 3364
rect 11132 3356 11140 3364
rect 92 3336 100 3344
rect 732 3336 740 3344
rect 1388 3336 1396 3344
rect 1980 3336 1988 3344
rect 5228 3336 5236 3344
rect 6588 3336 6596 3344
rect 9116 3336 9124 3344
rect 10492 3336 10500 3344
rect 1340 3316 1348 3324
rect 3180 3316 3188 3324
rect 6540 3316 6548 3324
rect 7724 3316 7732 3324
rect 9756 3316 9764 3324
rect 12268 3316 12276 3324
rect 1884 3296 1892 3304
rect 7084 3296 7092 3304
rect 7804 3296 7812 3304
rect 10428 3296 10436 3304
rect 8380 3276 8388 3284
rect 8524 3276 8532 3284
rect 12348 3276 12356 3284
rect 588 3236 596 3244
rect 2540 3236 2548 3244
rect 7868 3236 7876 3244
rect 11772 3236 11780 3244
rect 588 3176 596 3184
rect 1964 3176 1972 3184
rect 2540 3176 2548 3184
rect 3292 3176 3300 3184
rect 3932 3176 3940 3184
rect 3980 3176 3988 3184
rect 5228 3176 5236 3184
rect 5932 3176 5940 3184
rect 7868 3176 7876 3184
rect 9708 3176 9716 3184
rect 11036 3176 11044 3184
rect 11772 3176 11780 3184
rect 12972 3176 12980 3184
rect 2028 3156 2036 3164
rect 2620 3156 2628 3164
rect 4588 3156 4596 3164
rect 5868 3156 5876 3164
rect 92 3136 100 3144
rect 1884 3136 1892 3144
rect 3324 3136 3332 3144
rect 4636 3136 4644 3144
rect 7148 3136 7156 3144
rect 9036 3136 9044 3144
rect 10988 3136 10996 3144
rect 11644 3136 11652 3144
rect 12348 3136 12356 3144
rect 12924 3136 12932 3144
rect 2524 3116 2532 3124
rect 6572 3116 6580 3124
rect 8524 3116 8532 3124
rect 10332 3116 10340 3124
rect 10476 3116 10484 3124
rect 11772 3116 11780 3124
rect 1292 3096 1300 3104
rect 4636 3096 4644 3104
rect 7068 3096 7076 3104
rect 8380 3096 8388 3104
rect 3356 3076 3364 3084
rect 5212 3076 5220 3084
rect 8444 3076 8452 3084
rect 9852 3076 9860 3084
rect 11692 3076 11700 3084
rect 1228 3036 1236 3044
rect 7788 3036 7796 3044
rect 9788 3036 9796 3044
rect 44 2976 52 2984
rect 1340 2976 1348 2984
rect 3276 2976 3284 2984
rect 3292 2976 3300 2984
rect 3948 2976 3956 2984
rect 3980 2976 3988 2984
rect 6540 2976 6548 2984
rect 7836 2976 7844 2984
rect 9068 2976 9076 2984
rect 11628 2976 11636 2984
rect 668 2956 676 2964
rect 6428 2956 6436 2964
rect 12316 2956 12324 2964
rect 732 2936 740 2944
rect 1388 2936 1396 2944
rect 2588 2936 2596 2944
rect 5116 2936 5124 2944
rect 6588 2936 6596 2944
rect 7724 2936 7732 2944
rect 11036 2936 11044 2944
rect 2524 2916 2532 2924
rect 10316 2916 10324 2924
rect 1324 2896 1332 2904
rect 1884 2896 1892 2904
rect 2040 2896 2048 2904
rect 5276 2896 5284 2904
rect 5836 2896 5844 2904
rect 5996 2896 6004 2904
rect 7084 2896 7092 2904
rect 8524 2896 8532 2904
rect 10476 2896 10484 2904
rect 11772 2896 11780 2904
rect 2588 2876 2596 2884
rect 9756 2876 9764 2884
rect 1884 2836 1892 2844
rect 4620 2836 4628 2844
rect 5196 2836 5204 2844
rect 5276 2836 5284 2844
rect 6476 2836 6484 2844
rect 7084 2836 7092 2844
rect 9820 2836 9828 2844
rect 10476 2836 10484 2844
rect 11020 2836 11028 2844
rect 11772 2836 11780 2844
rect 1884 2776 1892 2784
rect 2028 2776 2036 2784
rect 3980 2776 3988 2784
rect 4620 2776 4628 2784
rect 5276 2776 5284 2784
rect 5900 2776 5908 2784
rect 5932 2776 5940 2784
rect 7084 2776 7092 2784
rect 7196 2776 7204 2784
rect 9180 2776 9188 2784
rect 9820 2776 9828 2784
rect 10476 2776 10484 2784
rect 11100 2776 11108 2784
rect 11772 2776 11780 2784
rect 668 2756 676 2764
rect 1340 2756 1348 2764
rect 2636 2756 2644 2764
rect 7820 2756 7828 2764
rect 9132 2756 9140 2764
rect 1372 2736 1380 2744
rect 2684 2736 2692 2744
rect 3836 2736 3844 2744
rect 6572 2736 6580 2744
rect 7868 2736 7876 2744
rect 8524 2736 8532 2744
rect 10332 2736 10340 2744
rect 10988 2736 10996 2744
rect 1820 2716 1828 2724
rect 3324 2716 3332 2724
rect 5276 2716 5284 2724
rect 9036 2716 9044 2724
rect 9100 2716 9108 2724
rect 9820 2716 9828 2724
rect 9884 2716 9892 2724
rect 10476 2716 10484 2724
rect 9116 2696 9124 2704
rect 92 2676 100 2684
rect 5196 2676 5204 2684
rect 5772 2676 5780 2684
rect 12268 2676 12276 2684
rect 12348 2636 12356 2644
rect 620 2576 628 2584
rect 636 2576 644 2584
rect 732 2576 740 2584
rect 3260 2576 3268 2584
rect 3980 2576 3988 2584
rect 4588 2576 4596 2584
rect 5884 2576 5892 2584
rect 5932 2576 5940 2584
rect 7228 2576 7236 2584
rect 9068 2576 9076 2584
rect 9676 2576 9684 2584
rect 9708 2576 9716 2584
rect 10364 2576 10372 2584
rect 11628 2576 11636 2584
rect 5278 2556 5286 2564
rect 8380 2556 8388 2564
rect 1388 2536 1396 2544
rect 2028 2536 2036 2544
rect 3340 2536 3348 2544
rect 4636 2536 4644 2544
rect 5244 2536 5252 2544
rect 8444 2536 8452 2544
rect 9740 2536 9748 2544
rect 10380 2536 10388 2544
rect 10492 2536 10500 2544
rect 11788 2536 11796 2544
rect 76 2496 84 2504
rect 1884 2496 1892 2504
rect 2684 2496 2692 2504
rect 3836 2496 3844 2504
rect 5132 2496 5140 2504
rect 7948 2496 7956 2504
rect 8524 2496 8532 2504
rect 5292 2476 5300 2484
rect 12924 2476 12932 2484
rect 76 2436 84 2444
rect 1884 2436 1892 2444
rect 2540 2436 2548 2444
rect 3180 2436 3188 2444
rect 3836 2436 3844 2444
rect 3932 2436 3940 2444
rect 5132 2436 5140 2444
rect 5884 2436 5892 2444
rect 6572 2436 6580 2444
rect 7868 2436 7876 2444
rect 8524 2436 8532 2444
rect 10988 2436 10996 2444
rect 76 2376 84 2384
rect 620 2376 628 2384
rect 1884 2376 1892 2384
rect 2028 2376 2036 2384
rect 2540 2376 2548 2384
rect 3292 2376 3300 2384
rect 3836 2376 3844 2384
rect 3948 2376 3956 2384
rect 4588 2376 4596 2384
rect 5132 2376 5140 2384
rect 6460 2376 6468 2384
rect 6572 2376 6580 2384
rect 7868 2376 7876 2384
rect 8380 2376 8388 2384
rect 8524 2376 8532 2384
rect 9788 2376 9796 2384
rect 10428 2376 10436 2384
rect 10988 2376 10996 2384
rect 12316 2376 12324 2384
rect 636 2356 644 2364
rect 1340 2356 1348 2364
rect 2620 2356 2628 2364
rect 11068 2356 11076 2364
rect 11132 2356 11140 2364
rect 1372 2336 1380 2344
rect 2668 2336 2676 2344
rect 3324 2336 3332 2344
rect 7084 2336 7092 2344
rect 7740 2336 7748 2344
rect 9036 2336 9044 2344
rect 9836 2336 9844 2344
rect 12284 2336 12292 2344
rect 76 2316 84 2324
rect 3116 2316 3124 2324
rect 5132 2316 5140 2324
rect 5276 2316 5284 2324
rect 7948 2316 7956 2324
rect 10332 2316 10340 2324
rect 11772 2316 11780 2324
rect 4684 2296 4692 2304
rect 9676 2296 9684 2304
rect 5772 2276 5780 2284
rect 6492 2276 6500 2284
rect 7788 2276 7796 2284
rect 10412 2276 10420 2284
rect 44 2176 52 2184
rect 3228 2176 3236 2184
rect 8380 2176 8388 2184
rect 9676 2176 9684 2184
rect 10364 2176 10372 2184
rect 2028 2156 2036 2164
rect 3980 2156 3988 2164
rect 6540 2156 6548 2164
rect 7228 2156 7236 2164
rect 11676 2156 11684 2164
rect 732 2136 740 2144
rect 1388 2136 1396 2144
rect 1980 2136 1988 2144
rect 3340 2136 3348 2144
rect 6588 2136 6596 2144
rect 7180 2136 7188 2144
rect 8444 2136 8452 2144
rect 9020 2136 9028 2144
rect 10316 2136 10324 2144
rect 11692 2136 11700 2144
rect 1964 2116 1972 2124
rect 3916 2116 3924 2124
rect 7164 2116 7172 2124
rect 10396 2116 10404 2124
rect 10972 2116 10980 2124
rect 1884 2096 1892 2104
rect 5276 2096 5284 2104
rect 7084 2096 7092 2104
rect 8524 2096 8532 2104
rect 9884 2096 9892 2104
rect 11772 2096 11780 2104
rect 3900 2076 3908 2084
rect 4604 2076 4612 2084
rect 4620 2076 4628 2084
rect 5788 2076 5796 2084
rect 11036 2076 11044 2084
rect 11644 2076 11652 2084
rect 2540 2036 2548 2044
rect 3180 2036 3188 2044
rect 3292 2036 3300 2044
rect 5276 2036 5284 2044
rect 9820 2036 9828 2044
rect 11772 2036 11780 2044
rect 12316 2036 12324 2044
rect 44 1976 52 1984
rect 1916 1976 1924 1984
rect 2028 1976 2036 1984
rect 2540 1976 2548 1984
rect 5276 1976 5284 1984
rect 5820 1976 5828 1984
rect 5884 1976 5892 1984
rect 7788 1976 7796 1984
rect 8492 1976 8500 1984
rect 9820 1976 9828 1984
rect 10444 1976 10452 1984
rect 11628 1976 11636 1984
rect 11772 1976 11780 1984
rect 732 1956 740 1964
rect 92 1936 100 1944
rect 2668 1936 2676 1944
rect 3836 1936 3844 1944
rect 5788 1936 5796 1944
rect 7148 1936 7156 1944
rect 7724 1936 7732 1944
rect 10348 1936 10356 1944
rect 12268 1936 12276 1944
rect 3324 1916 3332 1924
rect 5196 1916 5204 1924
rect 5276 1916 5284 1924
rect 9036 1916 9044 1924
rect 11836 1916 11844 1924
rect 4476 1896 4484 1904
rect 4540 1876 4548 1884
rect 11692 1876 11700 1884
rect 9708 1836 9716 1844
rect 44 1776 52 1784
rect 668 1776 676 1784
rect 1980 1776 1988 1784
rect 2028 1776 2036 1784
rect 2620 1776 2628 1784
rect 3932 1776 3940 1784
rect 3980 1776 3988 1784
rect 5196 1776 5204 1784
rect 6428 1776 6436 1784
rect 6460 1776 6468 1784
rect 8428 1776 8436 1784
rect 9724 1776 9732 1784
rect 732 1756 740 1764
rect 7788 1756 7796 1764
rect 11132 1756 11140 1764
rect 1868 1736 1876 1744
rect 2684 1736 2692 1744
rect 5116 1736 5124 1744
rect 5772 1736 5780 1744
rect 5836 1736 5844 1744
rect 6492 1736 6500 1744
rect 8540 1736 8548 1744
rect 9724 1736 9732 1744
rect 10492 1736 10500 1744
rect 3916 1716 3924 1724
rect 7068 1716 7076 1724
rect 10412 1716 10420 1724
rect 11708 1716 11716 1724
rect 1372 1696 1380 1704
rect 3836 1696 3844 1704
rect 5276 1696 5284 1704
rect 7884 1696 7892 1704
rect 9036 1696 9044 1704
rect 9196 1696 9204 1704
rect 9244 1696 9252 1704
rect 10332 1696 10340 1704
rect 10988 1696 10996 1704
rect 11052 1696 11060 1704
rect 11564 1696 11572 1704
rect 3324 1676 3332 1684
rect 7148 1676 7156 1684
rect 9820 1676 9828 1684
rect 12284 1676 12292 1684
rect 12300 1676 12308 1684
rect 8476 1656 8484 1664
rect 1372 1636 1380 1644
rect 3932 1636 3940 1644
rect 4620 1636 4628 1644
rect 5276 1636 5284 1644
rect 10988 1636 10996 1644
rect 44 1576 52 1584
rect 1372 1576 1380 1584
rect 1948 1576 1956 1584
rect 3228 1576 3236 1584
rect 4620 1576 4628 1584
rect 5276 1576 5284 1584
rect 7836 1576 7844 1584
rect 9180 1576 9188 1584
rect 10380 1576 10388 1584
rect 10988 1576 10996 1584
rect 11692 1576 11700 1584
rect 3180 1556 3188 1564
rect 9084 1556 9092 1564
rect 10380 1556 10388 1564
rect 716 1536 724 1544
rect 1868 1536 1876 1544
rect 2540 1536 2548 1544
rect 6572 1536 6580 1544
rect 7212 1536 7220 1544
rect 7868 1536 7876 1544
rect 9036 1536 9044 1544
rect 10332 1536 10340 1544
rect 10476 1536 10484 1544
rect 3996 1516 4004 1524
rect 4556 1516 4564 1524
rect 5276 1516 5284 1524
rect 6412 1516 6420 1524
rect 9740 1516 9748 1524
rect 9884 1516 9892 1524
rect 10988 1516 10996 1524
rect 12284 1516 12292 1524
rect 3820 1496 3828 1504
rect 11628 1496 11636 1504
rect 3244 1476 3252 1484
rect 4540 1476 4548 1484
rect 5196 1476 5204 1484
rect 5772 1476 5780 1484
rect 7164 1476 7172 1484
rect 700 1436 708 1444
rect 732 1436 740 1444
rect 5164 1436 5172 1444
rect 5900 1436 5908 1444
rect 5932 1436 5940 1444
rect 620 1376 628 1384
rect 1260 1376 1268 1384
rect 1932 1376 1940 1384
rect 1996 1376 2004 1384
rect 3228 1376 3236 1384
rect 3244 1376 3252 1384
rect 4572 1376 4580 1384
rect 8412 1376 8420 1384
rect 8428 1376 8436 1384
rect 1292 1336 1300 1344
rect 1868 1336 1876 1344
rect 3932 1336 3940 1344
rect 4636 1336 4644 1344
rect 7068 1336 7076 1344
rect 9740 1336 9748 1344
rect 3916 1316 3924 1324
rect 6428 1316 6436 1324
rect 7724 1316 7732 1324
rect 10396 1316 10404 1324
rect 10972 1316 10980 1324
rect 11692 1316 11700 1324
rect 1372 1296 1380 1304
rect 5132 1296 5140 1304
rect 6572 1296 6580 1304
rect 7788 1296 7796 1304
rect 8972 1296 8980 1304
rect 8524 1276 8532 1284
rect 10332 1276 10340 1284
rect 10348 1276 10356 1284
rect 11036 1276 11044 1284
rect 12284 1276 12292 1284
rect 12300 1276 12308 1284
rect 76 1236 84 1244
rect 2668 1236 2676 1244
rect 5132 1236 5140 1244
rect 5212 1236 5220 1244
rect 5788 1236 5796 1244
rect 9676 1236 9684 1244
rect 11660 1236 11668 1244
rect 76 1176 84 1184
rect 636 1176 644 1184
rect 1932 1176 1940 1184
rect 2668 1176 2676 1184
rect 5132 1176 5140 1184
rect 5788 1176 5796 1184
rect 6428 1176 6436 1184
rect 6524 1176 6532 1184
rect 6540 1176 6548 1184
rect 7228 1176 7236 1184
rect 9724 1176 9732 1184
rect 11660 1176 11668 1184
rect 11740 1176 11748 1184
rect 1292 1156 1300 1164
rect 3244 1156 3252 1164
rect 7180 1156 7188 1164
rect 11628 1156 11636 1164
rect 1244 1136 1252 1144
rect 2540 1136 2548 1144
rect 2556 1136 2564 1144
rect 3820 1136 3828 1144
rect 4620 1136 4628 1144
rect 5276 1136 5284 1144
rect 6572 1136 6580 1144
rect 7884 1136 7892 1144
rect 9100 1136 9108 1144
rect 76 1116 84 1124
rect 1372 1116 1380 1124
rect 5132 1116 5140 1124
rect 7084 1116 7092 1124
rect 7660 1116 7668 1124
rect 10332 1116 10340 1124
rect 11196 1116 11204 1124
rect 12284 1116 12292 1124
rect 9020 1096 9028 1104
rect 1292 1076 1300 1084
rect 7164 1076 7172 1084
rect 10412 1076 10420 1084
rect 4524 1036 4532 1044
rect 9788 1036 9796 1044
rect 10428 1036 10436 1044
rect 732 976 740 984
rect 1916 976 1924 984
rect 2572 976 2580 984
rect 3228 976 3236 984
rect 3292 976 3300 984
rect 3932 976 3940 984
rect 3980 976 3988 984
rect 6460 976 6468 984
rect 7196 976 7204 984
rect 11036 976 11044 984
rect 11132 976 11140 984
rect 5228 956 5236 964
rect 3340 936 3348 944
rect 7884 936 7892 944
rect 3916 916 3924 924
rect 9020 916 9028 924
rect 11708 916 11716 924
rect 76 896 84 904
rect 1372 896 1380 904
rect 7084 896 7092 904
rect 8524 896 8532 904
rect 10476 896 10484 904
rect 684 876 692 884
rect 5292 876 5300 884
rect 9100 876 9108 884
rect 9692 876 9700 884
rect 10332 876 10340 884
rect 12284 876 12292 884
rect 12300 876 12308 884
rect 76 836 84 844
rect 1372 836 1380 844
rect 1948 836 1956 844
rect 2668 836 2676 844
rect 4620 836 4628 844
rect 5788 836 5796 844
rect 7084 836 7092 844
rect 8524 836 8532 844
rect 10476 836 10484 844
rect 76 776 84 784
rect 636 776 644 784
rect 1276 776 1284 784
rect 1372 776 1380 784
rect 1916 776 1924 784
rect 2668 776 2676 784
rect 3212 776 3220 784
rect 4620 776 4628 784
rect 5788 776 5796 784
rect 6428 776 6436 784
rect 7084 776 7092 784
rect 7772 776 7780 784
rect 8524 776 8532 784
rect 10476 776 10484 784
rect 588 736 596 744
rect 2540 736 2548 744
rect 3836 736 3844 744
rect 4556 736 4564 744
rect 5276 736 5284 744
rect 6588 736 6596 744
rect 7740 736 7748 744
rect 9036 736 9044 744
rect 9772 736 9780 744
rect 10988 736 10996 744
rect 10332 716 10340 724
rect 10476 716 10484 724
rect 11196 716 11204 724
rect 12284 716 12292 724
rect 2588 696 2596 704
rect 4476 696 4484 704
rect 6540 696 6548 704
rect 11628 696 11636 704
rect 4540 676 4548 684
rect 5116 676 5124 684
rect 7788 676 7796 684
rect 11804 676 11812 684
rect 9676 656 9684 664
rect 8380 636 8388 644
rect 9724 636 9732 644
rect 11676 636 11684 644
rect 620 576 628 584
rect 1260 576 1268 584
rect 2572 576 2580 584
rect 3180 576 3188 584
rect 4524 576 4532 584
rect 6428 576 6436 584
rect 7132 576 7140 584
rect 7228 576 7236 584
rect 9084 576 9092 584
rect 9740 576 9748 584
rect 11628 556 11636 564
rect 4636 536 4644 544
rect 3820 516 3828 524
rect 10396 516 10404 524
rect 11580 516 11588 524
rect 76 496 84 504
rect 2684 496 2692 504
rect 5132 496 5140 504
rect 5276 496 5284 504
rect 5852 496 5860 504
rect 8368 496 8376 504
rect 10380 496 10388 504
rect 10476 496 10484 504
rect 1884 476 1892 484
rect 3836 476 3844 484
rect 4460 476 4468 484
rect 7868 476 7876 484
rect 11004 476 11012 484
rect 12300 476 12308 484
rect 76 436 84 444
rect 1372 436 1380 444
rect 2668 436 2676 444
rect 4572 436 4580 444
rect 5132 436 5140 444
rect 5918 436 5926 444
rect 6572 436 6580 444
rect 7132 436 7140 444
rect 8524 436 8532 444
rect 11772 436 11780 444
rect 76 376 84 384
rect 1372 376 1380 384
rect 2028 376 2036 384
rect 2668 376 2676 384
rect 5132 376 5140 384
rect 5918 376 5926 384
rect 6492 376 6500 384
rect 6572 376 6580 384
rect 8524 376 8532 384
rect 9068 376 9076 384
rect 10444 376 10452 384
rect 11132 376 11140 384
rect 11772 376 11780 384
rect 12380 376 12388 384
rect 636 356 644 364
rect 11068 356 11076 364
rect 588 336 596 344
rect 4524 336 4532 344
rect 4620 336 4628 344
rect 9020 336 9028 344
rect 9692 336 9700 344
rect 3836 316 3844 324
rect 3996 316 4004 324
rect 5068 316 5076 324
rect 7788 316 7796 324
rect 8524 316 8532 324
rect 9084 316 9092 324
rect 10268 316 10276 324
rect 11692 316 11700 324
rect 3340 296 3348 304
rect 7724 296 7732 304
rect 8380 296 8388 304
rect 8444 296 8452 304
rect 3292 276 3300 284
rect 4572 276 4580 284
rect 9852 276 9860 284
rect 5278 256 5286 264
rect 1980 236 1988 244
rect 3228 236 3236 244
rect 7132 236 7140 244
rect 684 176 692 184
rect 700 176 708 184
rect 1324 176 1332 184
rect 3868 176 3876 184
rect 3884 176 3892 184
rect 4572 176 4580 184
rect 6540 176 6548 184
rect 9068 176 9076 184
rect 11628 176 11636 184
rect 11676 176 11684 184
rect 6524 156 6532 164
rect 11692 156 11700 164
rect 1388 136 1396 144
rect 4636 136 4644 144
rect 6588 136 6596 144
rect 9020 136 9028 144
rect 10396 136 10404 144
rect 11788 136 11796 144
rect 5772 116 5780 124
rect 7724 116 7732 124
rect 8380 116 8388 124
rect 10396 116 10404 124
rect 10972 116 10980 124
rect 76 96 84 104
rect 1884 96 1892 104
rect 3324 96 3332 104
rect 7084 96 7092 104
rect 8524 96 8532 104
rect 9756 96 9764 104
rect 12284 96 12292 104
rect 2540 76 2548 84
rect 3196 76 3204 84
rect 7804 76 7812 84
rect 11052 76 11060 84
<< metal2 >>
rect 6413 9024 6419 9083
rect 6445 9024 6451 9083
rect 7069 9077 7091 9083
rect 3341 8944 3347 8976
rect 7069 8944 7075 9077
rect 7117 8984 7123 9083
rect 10317 9024 10323 9083
rect 10349 9024 10355 9083
rect 11629 8998 11635 9083
rect 11661 8998 11667 9083
rect 11741 9077 11763 9083
rect 11741 8984 11747 9077
rect 8541 8944 8547 8956
rect 11789 8944 11795 9083
rect 524 8890 532 8896
rect 1213 8884 1219 8904
rect 45 8664 51 8836
rect 589 8784 595 8836
rect 653 8757 668 8763
rect 524 8724 532 8730
rect 557 8716 563 8756
rect 653 8704 659 8757
rect 1213 8744 1219 8856
rect 1213 8724 1219 8736
rect 45 8604 51 8636
rect 637 8584 643 8596
rect 653 8544 659 8683
rect 1277 8537 1283 8683
rect 1293 8677 1299 8943
rect 1885 8884 1891 8896
rect 1325 8684 1331 8836
rect 1341 8764 1347 8816
rect 1389 8744 1395 8836
rect 1885 8784 1891 8836
rect 1901 8824 1907 8923
rect 2541 8784 2547 8836
rect 1949 8757 1964 8763
rect 1885 8724 1891 8756
rect 1949 8703 1955 8757
rect 3245 8704 3251 8943
rect 3885 8937 3923 8943
rect 3772 8890 3780 8896
rect 3316 8717 3324 8723
rect 1933 8697 1955 8703
rect 2605 8683 2612 8684
rect 1325 8584 1331 8656
rect 1389 8544 1395 8616
rect 77 8484 83 8496
rect 524 8324 532 8330
rect 557 8316 563 8376
rect 45 8204 51 8236
rect 77 8104 83 8116
rect 573 7944 579 8076
rect 524 7924 532 7930
rect 93 7804 99 7876
rect 93 7744 99 7776
rect 637 7737 643 7883
rect 653 7744 659 8536
rect 1213 8484 1219 8504
rect 1261 8384 1267 8523
rect 1213 8316 1219 8356
rect 1293 8284 1299 8543
rect 1933 8537 1939 8683
rect 2589 8677 2612 8683
rect 2605 8676 2612 8677
rect 2589 8584 2595 8596
rect 2525 8544 2531 8576
rect 1949 8537 1971 8543
rect 1885 8384 1891 8436
rect 1997 8384 2003 8436
rect 2045 8364 2051 8496
rect 1373 8344 1379 8356
rect 1885 8324 1891 8356
rect 2605 8284 2611 8676
rect 2685 8544 2691 8616
rect 3261 8543 3267 8683
rect 3245 8537 3267 8543
rect 3165 8496 3168 8504
rect 3165 8484 3171 8496
rect 3165 8364 3171 8476
rect 3181 8384 3187 8456
rect 3229 8384 3235 8416
rect 3261 8284 3267 8537
rect 3325 8464 3331 8496
rect 3772 8324 3780 8330
rect 3837 8324 3843 8376
rect 3901 8324 3907 8356
rect 3917 8284 3923 8937
rect 3997 8884 4003 8896
rect 3997 8864 4003 8876
rect 3997 8716 4003 8736
rect 4541 8584 4547 8676
rect 3997 8484 4003 8504
rect 4461 8316 4467 8336
rect 4557 8304 4563 8943
rect 4684 8890 4692 8896
rect 5140 8717 5148 8723
rect 5213 8704 5219 8943
rect 5869 8923 5875 8943
rect 5853 8917 5875 8923
rect 5277 8904 5283 8916
rect 5757 8716 5763 8776
rect 4573 8344 4579 8636
rect 5197 8537 5203 8683
rect 5245 8604 5251 8636
rect 5837 8584 5843 8636
rect 5853 8544 5859 8917
rect 5949 8884 5955 8904
rect 6573 8884 6579 8896
rect 6636 8890 6644 8896
rect 7741 8784 7747 8836
rect 6413 8716 6419 8756
rect 6573 8744 6579 8756
rect 7085 8724 7091 8756
rect 7149 8703 7155 8776
rect 7709 8724 7715 8736
rect 7901 8724 7907 8736
rect 7724 8710 7732 8716
rect 7884 8710 7892 8716
rect 7133 8697 7155 8703
rect 6509 8684 6515 8696
rect 7784 8696 7788 8704
rect 6496 8683 6515 8684
rect 6493 8676 6515 8683
rect 7805 8683 7812 8684
rect 6429 8584 6435 8616
rect 6461 8584 6467 8616
rect 5853 8536 5862 8544
rect 5133 8484 5139 8496
rect 5149 8484 5155 8523
rect 5277 8484 5283 8496
rect 5949 8484 5955 8504
rect 4684 8324 4692 8330
rect 1277 8137 1283 8283
rect 1293 8277 1308 8284
rect 1296 8276 1308 8277
rect 2605 8276 2612 8284
rect 4541 8277 4563 8283
rect 1293 8137 1315 8143
rect 1213 8084 1219 8096
rect 701 7984 707 7996
rect 733 7984 739 8076
rect 1261 8004 1267 8123
rect 1213 7916 1219 7956
rect 1261 7897 1267 7976
rect 1261 7784 1267 7796
rect 653 7736 662 7744
rect 669 7723 675 7743
rect 653 7717 675 7723
rect 524 7690 532 7696
rect 589 7544 595 7676
rect 653 7484 659 7717
rect 1277 7584 1283 7736
rect 1293 7504 1299 8137
rect 1436 8090 1444 8096
rect 1373 7944 1379 7976
rect 1389 7744 1395 7896
rect 1965 7883 1971 8276
rect 2525 8144 2531 8196
rect 2573 8184 2579 8256
rect 2045 8084 2051 8104
rect 2045 7916 2051 7976
rect 1949 7877 1971 7883
rect 1885 7704 1891 7716
rect 1373 7524 1379 7536
rect 1436 7524 1444 7530
rect 1933 7524 1939 7536
rect 1549 7484 1555 7502
rect 660 7476 662 7484
rect 669 7463 675 7483
rect 653 7457 675 7463
rect 29 7384 35 7456
rect 524 7290 532 7296
rect 557 7283 563 7304
rect 557 7277 579 7283
rect 573 7144 579 7277
rect 77 7124 83 7136
rect 524 6890 532 6896
rect 93 6744 99 6876
rect 605 6764 611 6923
rect 621 6784 627 6816
rect 68 6717 76 6723
rect 77 6504 83 6516
rect 45 6384 51 6396
rect 77 6344 83 6496
rect 621 6404 627 6436
rect 524 6324 532 6330
rect 557 6316 563 6376
rect 621 6343 627 6356
rect 605 6337 627 6343
rect 605 6297 611 6337
rect 45 6184 51 6196
rect 93 6144 99 6156
rect 653 6137 659 7457
rect 701 7384 707 7396
rect 733 7384 739 7396
rect 1309 7344 1315 7483
rect 1389 7344 1395 7376
rect 1296 7343 1315 7344
rect 1293 7336 1315 7343
rect 1949 7337 1955 7877
rect 2589 7737 2595 8276
rect 2621 7984 2627 8236
rect 3261 8143 3267 8276
rect 3245 8137 3267 8143
rect 3165 8084 3171 8104
rect 3213 8064 3219 8123
rect 2637 7984 2643 8016
rect 2637 7784 2643 7956
rect 2685 7944 2691 8056
rect 3165 7916 3171 7936
rect 2685 7744 2691 7756
rect 3229 7737 3235 7883
rect 3245 7877 3251 8137
rect 3325 7944 3331 8016
rect 3917 7883 3923 8276
rect 4541 8144 4547 8277
rect 5117 8144 5123 8296
rect 5181 8184 5187 8476
rect 5197 8384 5203 8476
rect 5917 8436 5918 8443
rect 5277 8384 5283 8436
rect 5917 8384 5923 8436
rect 5917 8377 5918 8384
rect 5949 8316 5955 8336
rect 6493 8304 6499 8676
rect 7133 8537 7139 8683
rect 7789 8677 7812 8683
rect 7805 8676 7812 8677
rect 7149 8537 7171 8543
rect 7069 8384 7075 8504
rect 7133 8384 7139 8396
rect 6636 8324 6644 8330
rect 7165 8284 7171 8537
rect 7389 8518 7395 8536
rect 7245 8344 7251 8496
rect 7709 8316 7715 8356
rect 7805 8284 7811 8676
rect 8381 8604 8387 8636
rect 8413 8604 8419 8636
rect 7869 8424 7875 8476
rect 7869 8344 7875 8376
rect 8221 8284 8227 8302
rect 5213 8144 5219 8283
rect 5869 8263 5875 8283
rect 5853 8257 5875 8263
rect 5245 8184 5251 8196
rect 5293 8144 5299 8196
rect 4621 8104 4627 8116
rect 4684 8090 4692 8096
rect 4621 7984 4627 8036
rect 4684 7924 4692 7930
rect 4061 7884 4067 7902
rect 3885 7877 3923 7883
rect 2365 7718 2371 7736
rect 2524 7704 2532 7710
rect 1997 7584 2003 7636
rect 2029 7584 2035 7596
rect 2509 7584 2515 7696
rect 3165 7644 3171 7696
rect 2541 7584 2547 7636
rect 3213 7604 3219 7723
rect 1997 7384 2003 7556
rect 3245 7504 3251 7743
rect 3885 7737 3891 7877
rect 3772 7690 3780 7696
rect 3853 7664 3859 7723
rect 3837 7544 3843 7556
rect 3485 7484 3491 7502
rect 2029 7384 2035 7436
rect 2573 7337 2579 7483
rect 2685 7344 2691 7396
rect 3261 7343 3267 7483
rect 3917 7344 3923 7877
rect 4477 7784 4483 7816
rect 4509 7784 4515 7816
rect 3997 7684 4003 7696
rect 4525 7384 4531 7436
rect 4541 7364 4547 7896
rect 4557 7744 4563 7883
rect 4637 7744 4643 7776
rect 5213 7744 5219 8136
rect 5277 7924 5283 7936
rect 5853 7903 5859 8257
rect 6509 8144 6515 8283
rect 7804 8276 7811 8284
rect 8445 8283 8451 8943
rect 9101 8937 9123 8943
rect 9053 8904 9059 8923
rect 8972 8890 8980 8896
rect 9037 8884 9043 8896
rect 9037 8784 9043 8836
rect 9149 8784 9155 8896
rect 9197 8884 9203 8904
rect 8972 8724 8980 8730
rect 9709 8697 9715 8756
rect 9757 8684 9763 8943
rect 9853 8884 9859 8904
rect 9884 8890 9892 8896
rect 10333 8724 10339 8776
rect 10397 8703 10403 8756
rect 10381 8697 10403 8703
rect 10413 8684 10419 8943
rect 11069 8923 11075 8943
rect 11053 8917 11075 8923
rect 10477 8744 10483 8776
rect 10924 8724 10932 8730
rect 10957 8716 10963 8736
rect 11053 8684 11059 8917
rect 11149 8884 11155 8904
rect 8541 8544 8547 8556
rect 9085 8537 9091 8683
rect 9101 8544 9107 8683
rect 9741 8544 9747 8683
rect 9754 8676 9763 8684
rect 11053 8676 11062 8684
rect 10317 8544 10323 8616
rect 10365 8584 10371 8616
rect 9101 8543 9120 8544
rect 9101 8536 9123 8543
rect 8972 8490 8980 8496
rect 9037 8484 9043 8496
rect 9069 8384 9075 8456
rect 8516 8317 8524 8323
rect 8445 8277 8467 8283
rect 6589 8144 6595 8156
rect 6496 8143 6515 8144
rect 6493 8136 6515 8143
rect 7165 8143 7171 8276
rect 7149 8137 7171 8143
rect 6429 7984 6435 8036
rect 5949 7916 5955 7936
rect 5405 7884 5411 7902
rect 5853 7897 5875 7903
rect 5853 7876 5862 7884
rect 5869 7877 5875 7897
rect 6093 7884 6099 7902
rect 6493 7884 6499 8136
rect 7069 8024 7075 8104
rect 7117 7984 7123 8016
rect 6636 7924 6644 7930
rect 5229 7784 5235 7796
rect 5277 7764 5283 7816
rect 5821 7764 5827 7836
rect 5277 7757 5278 7764
rect 3245 7337 3267 7343
rect 3901 7337 3923 7344
rect 701 7184 707 7276
rect 1213 7116 1219 7156
rect 701 6984 707 7016
rect 1277 6937 1283 7083
rect 1293 7077 1299 7336
rect 1341 7184 1347 7336
rect 1885 7284 1891 7296
rect 1885 7184 1891 7236
rect 2541 7184 2547 7236
rect 1373 7144 1379 7156
rect 1885 7124 1891 7156
rect 1949 7103 1955 7176
rect 3213 7124 3219 7323
rect 1933 7097 1955 7103
rect 1389 6944 1395 7036
rect 1213 6884 1219 6904
rect 1293 6683 1299 6943
rect 1933 6937 1939 7083
rect 2589 6944 2595 7083
rect 2621 7004 2627 7036
rect 2685 7024 2691 7076
rect 3245 6944 3251 7337
rect 3901 7336 3920 7337
rect 3772 7124 3780 7130
rect 1949 6937 1971 6943
rect 1325 6904 1331 6936
rect 1885 6884 1891 6896
rect 1436 6724 1444 6730
rect 733 6604 739 6636
rect 1277 6537 1283 6683
rect 1293 6677 1315 6683
rect 1389 6544 1395 6576
rect 1965 6544 1971 6937
rect 2045 6884 2051 6904
rect 2701 6884 2707 6904
rect 3325 6884 3331 6896
rect 2573 6784 2579 6796
rect 2669 6784 2675 6836
rect 3325 6784 3331 6836
rect 2045 6716 2051 6736
rect 2605 6676 2612 6684
rect 2029 6584 2035 6596
rect 2605 6544 2611 6676
rect 1213 6316 1219 6336
rect 1277 6137 1283 6283
rect 1293 6277 1299 6543
rect 2605 6536 2612 6544
rect 2524 6504 2532 6510
rect 1885 6484 1891 6496
rect 1373 6344 1379 6416
rect 1885 6384 1891 6436
rect 2557 6404 2563 6523
rect 2701 6484 2707 6504
rect 2669 6384 2675 6436
rect 2045 6316 2051 6336
rect 2189 6284 2195 6302
rect 524 6090 532 6096
rect 45 5984 51 6016
rect 93 5944 99 6056
rect 589 5984 595 6036
rect 524 5924 532 5930
rect 557 5916 563 5936
rect 621 5737 627 5883
rect 701 5784 707 5816
rect 733 5784 739 5796
rect 524 5690 532 5696
rect 45 5404 51 5636
rect 557 5604 563 5704
rect 77 5544 83 5576
rect 524 5524 532 5530
rect 573 5344 579 5416
rect 621 5384 627 5456
rect 653 5344 659 5743
rect 733 5584 739 5596
rect 1213 5516 1219 5536
rect 1277 5337 1283 5483
rect 1293 5477 1299 6143
rect 1933 6137 1939 6283
rect 1949 6277 1971 6283
rect 2509 6204 2515 6276
rect 2573 6224 2579 6236
rect 2589 6137 2595 6276
rect 3181 6204 3187 6236
rect 2685 6144 2691 6176
rect 2604 6136 2611 6144
rect 3261 6143 3267 6683
rect 3325 6484 3331 6496
rect 3293 6384 3299 6456
rect 3885 6344 3891 7056
rect 3901 6703 3907 7336
rect 3997 7284 4003 7304
rect 3981 7184 3987 7196
rect 4557 7103 4563 7736
rect 5133 7684 5139 7696
rect 5149 7664 5155 7723
rect 5149 7644 5155 7656
rect 5165 7584 5171 7656
rect 4653 7524 4659 7576
rect 4684 7524 4692 7530
rect 5197 7337 5203 7743
rect 5853 7737 5859 7876
rect 6493 7743 6499 7876
rect 6493 7737 6515 7743
rect 5789 7584 5795 7636
rect 5885 7624 5891 7636
rect 5949 7516 5955 7536
rect 5341 7344 5347 7356
rect 5821 7337 5827 7483
rect 6429 7404 6435 7436
rect 6461 7404 6467 7436
rect 6493 7343 6499 7737
rect 6541 7584 6547 7676
rect 7085 7524 7091 7556
rect 7165 7484 7171 8137
rect 7805 8144 7811 8276
rect 7805 8136 7812 8144
rect 7901 8084 7907 8104
rect 7869 7984 7875 8036
rect 8429 7984 8435 7996
rect 7724 7910 7732 7916
rect 7949 7884 7955 7902
rect 7805 7883 7812 7884
rect 7789 7877 7812 7883
rect 7805 7876 7812 7877
rect 7805 7744 7811 7876
rect 7805 7736 7812 7744
rect 7757 7683 7763 7696
rect 7748 7677 7763 7683
rect 7869 7584 7875 7636
rect 8381 7584 8387 7636
rect 7069 7344 7075 7416
rect 5133 7284 5139 7296
rect 4589 7184 4595 7216
rect 4621 7144 4627 7256
rect 5133 7184 5139 7236
rect 5117 7116 5123 7176
rect 5197 7103 5203 7156
rect 5805 7144 5811 7296
rect 4541 7097 4563 7103
rect 5181 7097 5203 7103
rect 3933 6984 3939 7076
rect 4525 6937 4531 7083
rect 4541 7077 4547 7097
rect 4541 6937 4563 6943
rect 5213 6937 5219 7083
rect 5773 6944 5779 7036
rect 5853 6963 5859 7343
rect 6493 7337 6515 7343
rect 5869 7024 5875 7236
rect 6477 6984 6483 7016
rect 5853 6957 5875 6963
rect 5853 6936 5862 6944
rect 5869 6937 5875 6957
rect 6493 6944 6499 7337
rect 6573 7144 6579 7296
rect 6636 7290 6644 7296
rect 7092 7117 7100 7123
rect 7165 7083 7171 7476
rect 7229 7384 7235 7396
rect 7773 7337 7779 7483
rect 7789 7477 7812 7483
rect 8381 7384 8387 7476
rect 8413 7384 8419 7816
rect 8429 7784 8435 7836
rect 8429 7584 8435 7756
rect 8461 7337 8467 8277
rect 9021 8144 9027 8236
rect 9069 8184 9075 8256
rect 8525 8084 8531 8096
rect 8972 7924 8980 7930
rect 9117 7883 9123 8536
rect 9709 8384 9715 8416
rect 9197 8316 9203 8336
rect 9725 8184 9731 8216
rect 9677 7984 9683 8016
rect 9085 7877 9123 7883
rect 9021 7744 9027 7816
rect 9069 7784 9075 7856
rect 8525 7704 8531 7716
rect 9085 7704 9091 7736
rect 8972 7524 8980 7530
rect 8541 7404 8547 7496
rect 9117 7483 9123 7877
rect 9677 7784 9683 7796
rect 9741 7784 9747 7936
rect 9757 7737 9763 8543
rect 10413 8537 10419 8676
rect 11037 8544 11043 8676
rect 11677 8584 11683 8756
rect 12269 8744 12275 8904
rect 11836 8724 11844 8730
rect 11069 8523 11075 8543
rect 11709 8537 11715 8683
rect 12317 8584 12323 8616
rect 12221 8544 12227 8556
rect 11053 8517 11075 8523
rect 9821 8504 9827 8516
rect 9884 8490 9892 8496
rect 9789 8384 9795 8476
rect 9821 8344 9827 8476
rect 10477 8384 10483 8436
rect 10333 8324 10339 8356
rect 10989 8344 10995 8376
rect 11005 8344 11011 8456
rect 11053 8284 11059 8517
rect 11149 8484 11155 8504
rect 11836 8490 11844 8496
rect 11773 8384 11779 8436
rect 11101 8297 11107 8376
rect 11149 8316 11155 8336
rect 11836 8324 11844 8330
rect 10333 8024 10339 8096
rect 10317 7944 10323 7996
rect 10381 7984 10387 8076
rect 9853 7916 9859 7936
rect 9884 7924 9892 7930
rect 10413 7884 10419 8283
rect 11053 8276 11062 8284
rect 11069 8263 11075 8283
rect 11053 8257 11075 8263
rect 11053 8144 11059 8257
rect 11629 8184 11635 8196
rect 11677 8184 11683 8316
rect 11053 8136 11062 8144
rect 10637 8118 10643 8136
rect 11069 8123 11075 8143
rect 11053 8117 11075 8123
rect 10924 7924 10932 7930
rect 10957 7916 10963 7936
rect 10989 7904 10995 8076
rect 11021 8044 11027 8096
rect 11037 8084 11043 8096
rect 11053 7884 11059 8117
rect 11293 7884 11299 7902
rect 11693 7884 11699 8276
rect 11789 8144 11795 8216
rect 12269 8204 12275 8276
rect 12333 8164 12339 8236
rect 12349 8137 12355 8943
rect 12285 8084 12291 8096
rect 12285 7984 12291 8036
rect 12285 7924 12291 7936
rect 11053 7876 11062 7884
rect 10413 7737 10419 7876
rect 11021 7784 11027 7856
rect 9341 7718 9347 7736
rect 9981 7718 9987 7736
rect 10637 7718 10643 7736
rect 9197 7684 9203 7704
rect 9853 7684 9859 7704
rect 9884 7690 9892 7696
rect 9261 7484 9267 7502
rect 9085 7477 9123 7483
rect 9021 7344 9027 7416
rect 7741 7144 7747 7156
rect 7757 7104 7763 7323
rect 8685 7318 8691 7336
rect 7149 7077 7171 7083
rect 4461 6884 4467 6904
rect 4509 6784 4515 6923
rect 4621 6904 4627 6916
rect 4684 6890 4692 6896
rect 5277 6884 5283 6896
rect 4621 6784 4627 6836
rect 5277 6784 5283 6836
rect 4509 6764 4515 6776
rect 4653 6716 4659 6776
rect 4684 6724 4692 6730
rect 3901 6697 3923 6703
rect 3772 6324 3780 6330
rect 3917 6283 3923 6697
rect 4525 6584 4531 6616
rect 3997 6484 4003 6504
rect 3997 6324 4003 6336
rect 3885 6277 3923 6283
rect 3821 6144 3827 6196
rect 3869 6184 3875 6216
rect 3245 6137 3267 6143
rect 1325 6104 1331 6136
rect 1885 6104 1891 6116
rect 2509 6084 2515 6104
rect 1405 6043 1411 6076
rect 1389 6037 1411 6043
rect 1389 5944 1395 6037
rect 1885 5984 1891 6036
rect 2589 5984 2595 6056
rect 2605 5884 2611 6136
rect 1325 5784 1331 5836
rect 1389 5744 1395 5816
rect 1933 5737 1939 5883
rect 1949 5877 1971 5883
rect 2605 5876 2612 5884
rect 2589 5737 2595 5876
rect 2685 5744 2691 5756
rect 1901 5704 1907 5723
rect 1325 5584 1331 5636
rect 1373 5544 1379 5616
rect 1885 5584 1891 5636
rect 1885 5524 1891 5536
rect 1389 5344 1395 5456
rect 77 5284 83 5296
rect 77 5184 83 5236
rect 589 5144 595 5256
rect 637 5184 643 5216
rect 524 4890 532 4896
rect 93 4744 99 4856
rect 524 4724 532 4730
rect 557 4716 563 4736
rect 93 4544 99 4576
rect 653 4537 659 5336
rect 733 5184 739 5196
rect 1277 4937 1283 5083
rect 1293 5077 1299 5343
rect 1933 5337 1939 5483
rect 1965 5384 1971 5396
rect 1885 5284 1891 5296
rect 1885 5184 1891 5236
rect 1389 4964 1395 5076
rect 1213 4716 1219 4736
rect 1277 4537 1283 4683
rect 1293 4677 1299 4943
rect 1933 4937 1939 5083
rect 1885 4904 1891 4916
rect 1885 4784 1891 4836
rect 1981 4764 1987 5636
rect 2029 5584 2035 5596
rect 2541 5584 2547 5636
rect 2685 5544 2691 5596
rect 3165 5516 3171 5536
rect 2445 5484 2451 5502
rect 2573 5337 2579 5483
rect 2013 5144 2019 5256
rect 2029 5184 2035 5216
rect 2541 5184 2547 5236
rect 2573 4937 2579 5083
rect 3213 5004 3219 5236
rect 3245 5084 3251 6137
rect 3261 5984 3267 6116
rect 3885 6064 3891 6256
rect 3325 5944 3331 5956
rect 3772 5924 3780 5930
rect 3853 5924 3859 6056
rect 3277 5784 3283 5896
rect 3917 5884 3923 6277
rect 4525 6104 4531 6236
rect 4557 6137 4563 6683
rect 5213 6537 5219 6683
rect 5853 6563 5859 6936
rect 5901 6784 5907 6923
rect 5949 6744 5955 6904
rect 6413 6716 6419 6756
rect 6461 6697 6467 6776
rect 6509 6684 6515 6943
rect 6636 6890 6644 6896
rect 6573 6744 6579 6776
rect 6925 6684 6931 6702
rect 6496 6683 6515 6684
rect 6493 6676 6515 6683
rect 7165 6683 7171 7077
rect 7789 6984 7795 6996
rect 7821 6964 7827 7256
rect 7885 7144 7891 7196
rect 7901 7184 7907 7304
rect 8525 7184 8531 7236
rect 8429 6937 8435 7083
rect 8461 6943 8467 7083
rect 8445 6937 8467 6943
rect 8685 6918 8691 6936
rect 7245 6884 7251 6904
rect 8365 6884 8371 6904
rect 9101 6884 9107 6896
rect 7725 6744 7731 6796
rect 8381 6784 8387 6796
rect 8525 6784 8531 6836
rect 8516 6717 8524 6723
rect 7149 6677 7171 6683
rect 5853 6557 5875 6563
rect 5869 6537 5875 6557
rect 6493 6544 6499 6676
rect 7165 6544 7171 6677
rect 7805 6676 7812 6684
rect 7805 6544 7811 6676
rect 7885 6544 7891 6556
rect 7804 6536 7811 6544
rect 5133 6484 5139 6496
rect 5949 6484 5955 6504
rect 5917 6436 5918 6443
rect 5277 6384 5283 6436
rect 5917 6384 5923 6436
rect 6429 6404 6435 6436
rect 6461 6404 6467 6436
rect 6477 6384 6483 6496
rect 5917 6377 5918 6384
rect 6429 6364 6435 6376
rect 5133 6324 5139 6336
rect 5277 6324 5283 6356
rect 5949 6316 5955 6336
rect 5165 6184 5171 6216
rect 3997 5916 4003 5936
rect 3885 5737 3891 5883
rect 3901 5877 3923 5884
rect 3901 5876 3920 5877
rect 3901 5737 3907 5876
rect 4477 5804 4483 5836
rect 3837 5684 3843 5696
rect 4461 5664 4467 5704
rect 3837 5584 3843 5636
rect 3949 5584 3955 5656
rect 3772 5524 3780 5530
rect 4461 5516 4467 5596
rect 4541 5483 4547 6116
rect 4653 6084 4659 6104
rect 4684 6090 4692 6096
rect 4637 5944 4643 6056
rect 4637 5744 4643 5756
rect 5197 5737 5203 5883
rect 5213 5877 5219 6283
rect 5853 6276 5862 6284
rect 5245 6184 5251 6216
rect 5293 6144 5299 6216
rect 5853 5903 5859 6276
rect 6477 6164 6483 6236
rect 6493 6143 6499 6536
rect 6573 6484 6579 6496
rect 6636 6490 6644 6496
rect 7165 6283 7171 6536
rect 7181 6404 7187 6436
rect 7245 6316 7251 6336
rect 7149 6277 7171 6283
rect 6589 6224 6595 6276
rect 7117 6184 7123 6216
rect 7069 6144 7075 6176
rect 6493 6137 6515 6143
rect 6636 6090 6644 6096
rect 5949 5916 5955 5936
rect 5853 5897 5875 5903
rect 5869 5877 5875 5897
rect 5837 5744 5843 5876
rect 6477 5784 6483 6056
rect 6573 5984 6579 6036
rect 7149 5984 7155 6156
rect 6636 5924 6644 5930
rect 6493 5784 6499 5916
rect 5133 5704 5139 5716
rect 4557 5524 4563 5576
rect 4653 5516 4659 5556
rect 5133 5544 5139 5596
rect 3341 5364 3347 5476
rect 3389 5344 3395 5356
rect 3885 5337 3891 5483
rect 3981 5384 3987 5416
rect 4525 5337 4531 5483
rect 4541 5477 4563 5483
rect 4541 5337 4563 5343
rect 5213 5337 5219 5716
rect 5949 5684 5955 5704
rect 5789 5584 5795 5636
rect 6509 5484 6515 5883
rect 6589 5744 6595 5816
rect 7165 5744 7171 6277
rect 7805 6223 7811 6536
rect 8428 6504 8436 6510
rect 7821 6384 7827 6436
rect 8365 6316 8371 6336
rect 7789 6217 7811 6223
rect 7229 6184 7235 6196
rect 7789 6137 7795 6217
rect 7804 6136 7811 6144
rect 8445 6143 8451 6676
rect 8461 6584 8467 6596
rect 9117 6544 9123 7477
rect 9725 7184 9731 7596
rect 9821 7584 9827 7636
rect 9853 7524 9859 7676
rect 10477 7584 10483 7636
rect 11037 7584 11043 7656
rect 10477 7524 10483 7536
rect 11053 7503 11059 7876
rect 11629 7804 11635 7836
rect 11661 7804 11667 7836
rect 11693 7743 11699 7876
rect 11741 7764 11747 7836
rect 12269 7744 12275 7816
rect 11693 7737 11715 7743
rect 11933 7718 11939 7736
rect 11836 7690 11844 7696
rect 11101 7524 11107 7636
rect 11773 7584 11779 7636
rect 11773 7524 11779 7536
rect 11836 7524 11844 7530
rect 11053 7497 11075 7503
rect 9197 7116 9203 7136
rect 9341 6918 9347 6936
rect 9709 6784 9715 6816
rect 9197 6716 9203 6736
rect 8972 6490 8980 6496
rect 8525 6344 8531 6356
rect 8972 6324 8980 6330
rect 9101 6284 9107 6543
rect 9181 6524 9187 6556
rect 9757 6544 9763 7483
rect 10365 7404 10371 7436
rect 10413 7337 10419 7483
rect 11053 7476 11062 7484
rect 11069 7477 11075 7497
rect 10477 7284 10483 7296
rect 9805 7124 9811 7276
rect 10477 7184 10483 7236
rect 10324 7137 10332 7143
rect 9853 7116 9859 7136
rect 9884 7124 9892 7130
rect 10317 6944 10323 7096
rect 10317 6924 10323 6936
rect 9884 6890 9892 6896
rect 10381 6584 10387 7036
rect 10397 6984 10403 7116
rect 11053 7103 11059 7476
rect 11101 7384 11107 7396
rect 11133 7384 11139 7396
rect 11693 7343 11699 7476
rect 12269 7344 12275 7416
rect 11693 7337 11715 7343
rect 11469 7318 11475 7336
rect 11613 7264 11619 7304
rect 11836 7290 11844 7296
rect 11773 7184 11779 7236
rect 11149 7116 11155 7136
rect 11773 7124 11779 7136
rect 11836 7124 11844 7130
rect 11053 7097 11075 7103
rect 10413 6937 10419 7083
rect 10973 6944 10979 7096
rect 11053 7076 11062 7084
rect 11069 7077 11075 7097
rect 11053 6963 11059 7076
rect 11677 6984 11683 7116
rect 11053 6957 11075 6963
rect 11053 6936 11062 6944
rect 11069 6937 11075 6957
rect 10477 6784 10483 6836
rect 10989 6744 10995 6856
rect 11037 6784 11043 6896
rect 11037 6684 11043 6716
rect 11053 6703 11059 6936
rect 11149 6864 11155 6904
rect 11053 6697 11075 6703
rect 11053 6676 11062 6684
rect 11069 6677 11075 6697
rect 9517 6518 9523 6536
rect 9741 6304 9747 6543
rect 9754 6536 9763 6544
rect 10333 6484 10339 6496
rect 9821 6324 9827 6476
rect 9853 6316 9859 6336
rect 9884 6324 9892 6330
rect 10397 6304 10403 6676
rect 10924 6490 10932 6496
rect 10461 6324 10467 6476
rect 10477 6324 10483 6336
rect 11053 6303 11059 6676
rect 11661 6604 11667 6636
rect 11693 6543 11699 7076
rect 11709 6984 11715 6996
rect 11741 6784 11747 7056
rect 12269 7004 12275 7076
rect 12317 7004 12323 7436
rect 12333 6964 12339 7036
rect 11789 6744 11795 6816
rect 12269 6804 12275 6904
rect 12285 6784 12291 6836
rect 12925 6744 12931 6796
rect 12445 6716 12451 6736
rect 12397 6697 12403 6716
rect 12349 6677 12371 6683
rect 12317 6584 12323 6616
rect 11693 6537 11715 6543
rect 11693 6523 11699 6537
rect 11693 6517 11715 6523
rect 11149 6316 11155 6336
rect 11053 6297 11075 6303
rect 9101 6283 9120 6284
rect 9085 6277 9123 6283
rect 9101 6276 9123 6277
rect 9021 6144 9027 6156
rect 8445 6137 8467 6143
rect 7565 6118 7571 6136
rect 7245 5916 7251 5936
rect 7805 5884 7811 6136
rect 7869 6064 7875 6076
rect 7837 5944 7843 6036
rect 8413 5984 8419 6016
rect 7805 5876 7812 5884
rect 7789 5744 7795 5876
rect 8381 5784 8387 5816
rect 7565 5718 7571 5736
rect 7724 5704 7732 5710
rect 7709 5644 7715 5696
rect 7901 5684 7907 5704
rect 8445 5684 8451 5836
rect 8461 5737 8467 6137
rect 8525 6084 8531 6096
rect 8477 5984 8483 6056
rect 8972 5924 8980 5930
rect 9117 5883 9123 6276
rect 9181 6184 9187 6196
rect 9757 6144 9763 6283
rect 9837 6144 9843 6176
rect 9677 5984 9683 6056
rect 9741 5904 9747 6143
rect 9754 6136 9763 6144
rect 10413 6137 10419 6283
rect 11053 6276 11062 6284
rect 11069 6277 11075 6297
rect 11053 6163 11059 6276
rect 11053 6157 11075 6163
rect 11053 6136 11062 6144
rect 11069 6137 11075 6157
rect 11709 6137 11715 6517
rect 11725 6384 11731 6476
rect 11789 6344 11795 6510
rect 11836 6490 11844 6496
rect 12292 6317 12300 6323
rect 12317 6184 12323 6216
rect 10477 5984 10483 6036
rect 9884 5924 9892 5930
rect 9085 5877 9123 5883
rect 8557 5864 8563 5876
rect 8685 5718 8691 5736
rect 8525 5684 8531 5696
rect 7085 5584 7091 5636
rect 7741 5584 7747 5636
rect 8525 5584 8531 5636
rect 9021 5564 9027 5676
rect 9069 5604 9075 5636
rect 7085 5524 7091 5556
rect 7757 5497 7763 5556
rect 7901 5516 7907 5536
rect 8605 5484 8611 5502
rect 6496 5483 6515 5484
rect 6493 5476 6515 5483
rect 5773 5344 5779 5416
rect 5821 5384 5827 5436
rect 5853 5363 5859 5476
rect 6477 5384 6483 5456
rect 5853 5357 5875 5363
rect 5853 5336 5862 5344
rect 5869 5337 5875 5357
rect 3772 5290 3780 5296
rect 3917 5084 3923 5316
rect 4684 5290 4692 5296
rect 4509 5184 4515 5196
rect 4621 5184 4627 5236
rect 5277 5184 5283 5236
rect 3997 5124 4003 5136
rect 4684 5124 4692 5130
rect 3901 5077 3923 5084
rect 3901 5076 3920 5077
rect 2604 4936 2611 4944
rect 1885 4724 1891 4736
rect 2045 4716 2051 4736
rect 2189 4684 2195 4702
rect 524 4490 532 4496
rect 1213 4484 1219 4496
rect 45 4384 51 4416
rect 45 4184 51 4356
rect 77 4344 83 4476
rect 589 4384 595 4436
rect 733 4384 739 4416
rect 524 4324 532 4330
rect 557 4316 563 4336
rect 524 4090 532 4096
rect 557 4084 563 4104
rect 573 3944 579 4036
rect 621 3984 627 4076
rect 653 3884 659 4283
rect 1277 4137 1283 4283
rect 1293 4277 1299 4543
rect 1933 4537 1939 4683
rect 1949 4677 1971 4683
rect 2029 4584 2035 4616
rect 2605 4544 2611 4936
rect 2685 4824 2691 4876
rect 2685 4744 2691 4796
rect 3165 4784 3171 4896
rect 3165 4716 3171 4736
rect 3245 4683 3251 5076
rect 3821 5004 3827 5076
rect 3869 4964 3875 5036
rect 3901 4937 3907 5076
rect 3981 4984 3987 5016
rect 3772 4890 3780 4896
rect 3325 4724 3331 4856
rect 3837 4744 3843 4776
rect 3245 4677 3267 4683
rect 2605 4543 2612 4544
rect 2589 4537 2612 4543
rect 3261 4537 3267 4677
rect 2605 4536 2612 4537
rect 1885 4504 1891 4516
rect 1933 4464 1939 4510
rect 1341 4404 1347 4436
rect 1885 4384 1891 4436
rect 2029 4384 2035 4396
rect 2541 4384 2547 4436
rect 2621 4384 2627 4476
rect 2653 4464 2659 4523
rect 2685 4344 2691 4456
rect 3229 4364 3235 4436
rect 3325 4384 3331 4436
rect 3869 4384 3875 4576
rect 2557 4297 2563 4336
rect 3332 4317 3340 4323
rect 1389 4144 1395 4176
rect 1293 4123 1299 4143
rect 1933 4137 1939 4283
rect 1965 4184 1971 4196
rect 2573 4137 2579 4283
rect 3181 4184 3187 4216
rect 3245 4144 3251 4283
rect 3261 4137 3267 4283
rect 1293 4117 1315 4123
rect 1229 3984 1235 4016
rect 660 3876 662 3884
rect 669 3863 675 3883
rect 653 3857 675 3863
rect 45 3784 51 3796
rect 93 3744 99 3796
rect 653 3744 659 3857
rect 653 3743 662 3744
rect 637 3737 662 3743
rect 653 3736 662 3737
rect 669 3723 675 3743
rect 653 3717 675 3723
rect 524 3690 532 3696
rect 557 3604 563 3704
rect 573 3544 579 3616
rect 637 3584 643 3596
rect 45 3384 51 3396
rect 93 3344 99 3396
rect 653 3337 659 3717
rect 1213 3516 1219 3536
rect 1309 3484 1315 4117
rect 2524 4104 2532 4110
rect 1373 3944 1379 3996
rect 1885 3984 1891 4036
rect 2557 3984 2563 4123
rect 2605 4044 2611 4096
rect 2701 4084 2707 4104
rect 1885 3924 1891 3936
rect 1949 3877 1971 3883
rect 1373 3664 1379 3696
rect 1436 3690 1444 3696
rect 1373 3544 1379 3576
rect 1277 3337 1283 3483
rect 1304 3476 1315 3484
rect 1965 3483 1971 3877
rect 2509 3724 2515 3876
rect 2605 3584 2611 4036
rect 2621 3784 2627 4056
rect 2637 3984 2643 4016
rect 3181 3964 3187 4036
rect 3229 3737 3235 3883
rect 3245 3877 3251 4136
rect 3293 3984 3299 4036
rect 3332 3937 3340 3943
rect 3772 3924 3780 3930
rect 3661 3884 3667 3902
rect 3917 3883 3923 4916
rect 4461 4864 4467 4904
rect 3949 4784 3955 4796
rect 4461 4716 4467 4736
rect 4541 4683 4547 5076
rect 4589 4984 4595 5056
rect 4637 4944 4643 5016
rect 5117 5004 5123 5076
rect 5133 4884 5139 4896
rect 4684 4724 4692 4730
rect 4541 4677 4563 4683
rect 4541 4544 4547 4677
rect 5101 4664 5107 4676
rect 4493 4297 4499 4476
rect 4509 4324 4515 4436
rect 4541 4277 4547 4536
rect 4605 4344 4611 4496
rect 4684 4490 4692 4496
rect 5165 4344 5171 4436
rect 5181 4310 5187 4876
rect 5213 4537 5219 5083
rect 5437 4926 5443 4936
rect 5837 4884 5843 5036
rect 5853 4963 5859 5336
rect 5949 5284 5955 5304
rect 6493 5083 6499 5476
rect 6589 5344 6595 5416
rect 7133 5337 7139 5483
rect 7149 5337 7171 5343
rect 7085 5304 7091 5316
rect 6636 5124 6644 5130
rect 6557 5097 6563 5116
rect 6493 5077 6515 5083
rect 5853 4957 5875 4963
rect 5869 4937 5875 4957
rect 6493 4944 6499 5077
rect 5917 4836 5918 4843
rect 5917 4784 5923 4836
rect 5917 4777 5918 4784
rect 5757 4716 5763 4756
rect 5901 4697 5907 4716
rect 5853 4683 5862 4684
rect 5837 4677 5862 4683
rect 5853 4676 5862 4677
rect 5821 4584 5827 4616
rect 5837 4584 5843 4596
rect 4554 4276 4563 4284
rect 4477 4184 4483 4196
rect 4509 4184 4515 4196
rect 4525 4184 4531 4216
rect 4509 4084 4515 4136
rect 4509 3984 4515 4076
rect 3885 3877 3923 3883
rect 3821 3744 3827 3816
rect 3869 3784 3875 3856
rect 3245 3737 3267 3743
rect 2669 3544 2675 3656
rect 1949 3477 1971 3483
rect 1389 3344 1395 3356
rect 524 3290 532 3296
rect 93 3144 99 3256
rect 589 3184 595 3236
rect 1293 3104 1299 3343
rect 1885 3304 1891 3316
rect 1885 3144 1891 3256
rect 1436 3124 1444 3130
rect 45 2984 51 3016
rect 621 2937 627 3083
rect 1229 3004 1235 3036
rect 1309 2944 1315 3083
rect 1389 2944 1395 3016
rect 524 2890 532 2896
rect 524 2724 532 2730
rect 93 2604 99 2676
rect 621 2584 627 2616
rect 637 2584 643 2596
rect 653 2544 659 2943
rect 1296 2943 1315 2944
rect 1293 2936 1315 2943
rect 1949 2943 1955 3477
rect 2525 3404 2531 3476
rect 3229 3344 3235 3483
rect 3245 3477 3251 3737
rect 3325 3544 3331 3696
rect 3772 3524 3780 3530
rect 3901 3524 3907 3696
rect 3661 3484 3667 3502
rect 3917 3484 3923 3877
rect 4541 3784 4547 3916
rect 4477 3584 4483 3676
rect 4141 3484 4147 3502
rect 3901 3483 3923 3484
rect 3885 3477 3923 3483
rect 3901 3476 3920 3477
rect 4557 3477 4563 4276
rect 5181 4137 5187 4283
rect 5197 4277 5203 4516
rect 5277 4484 5283 4496
rect 5245 4384 5251 4476
rect 5805 4324 5811 4356
rect 5773 4144 5779 4196
rect 5821 4184 5827 4256
rect 4605 3924 4611 4036
rect 4684 3924 4692 3930
rect 4653 3644 4659 3696
rect 4684 3690 4692 3696
rect 5117 3544 5123 3656
rect 5181 3584 5187 4056
rect 5293 4044 5299 4104
rect 5277 3984 5283 4036
rect 5277 3924 5283 3936
rect 4684 3524 4692 3530
rect 3293 3404 3299 3436
rect 1965 3184 1971 3316
rect 2509 3284 2515 3304
rect 2509 3124 2515 3256
rect 2541 3184 2547 3236
rect 2524 3110 2532 3116
rect 3229 3110 3235 3136
rect 2589 2944 2595 3083
rect 1949 2937 1971 2943
rect 2605 2936 2612 2944
rect 1213 2716 1219 2756
rect 1261 2697 1267 2776
rect 1277 2537 1283 2683
rect 1293 2677 1299 2936
rect 1325 2904 1331 2936
rect 1885 2884 1891 2896
rect 2013 2864 2019 2923
rect 2045 2884 2051 2896
rect 1885 2784 1891 2836
rect 2029 2784 2035 2796
rect 1373 2744 1379 2776
rect 2509 2716 2515 2736
rect 2605 2684 2611 2936
rect 2701 2884 2707 2904
rect 2685 2744 2691 2776
rect 1389 2544 1395 2616
rect 77 2504 83 2516
rect 77 2384 83 2436
rect 621 2384 627 2416
rect 77 2324 83 2336
rect 45 2184 51 2216
rect 524 2090 532 2096
rect 45 1984 51 1996
rect 93 1944 99 2036
rect 524 1924 532 1930
rect 557 1916 563 1936
rect 45 1784 51 1796
rect 524 1690 532 1696
rect 557 1684 563 1704
rect 45 1584 51 1596
rect 524 1524 532 1530
rect 557 1516 563 1536
rect 621 1384 627 1456
rect 77 1184 83 1236
rect 637 1184 643 1416
rect 653 1344 659 2536
rect 1213 2484 1219 2504
rect 1213 2316 1219 2356
rect 1261 2297 1267 2376
rect 1277 2137 1283 2283
rect 1293 2277 1299 2543
rect 1933 2537 1939 2683
rect 2573 2537 2579 2683
rect 2604 2676 2611 2684
rect 3245 2683 3251 3336
rect 3293 3184 3299 3276
rect 3277 2984 3283 3156
rect 3325 3144 3331 3296
rect 3772 3124 3780 3130
rect 3357 3064 3363 3076
rect 3293 2984 3299 3016
rect 3885 2937 3891 3083
rect 3901 3077 3907 3476
rect 3917 3384 3923 3456
rect 3933 3384 3939 3436
rect 3933 3184 3939 3296
rect 3949 2984 3955 3416
rect 3981 3384 3987 3396
rect 4541 3343 4547 3476
rect 4541 3337 4563 3343
rect 4509 3284 4515 3323
rect 3981 3184 3987 3276
rect 4461 3116 4467 3156
rect 3981 2984 3987 3016
rect 3325 2724 3331 2756
rect 3837 2744 3843 2876
rect 3853 2864 3859 2923
rect 3245 2677 3267 2683
rect 1885 2484 1891 2496
rect 1885 2384 1891 2436
rect 1901 2404 1907 2523
rect 1924 2516 1926 2524
rect 2509 2484 2515 2504
rect 2557 2464 2563 2523
rect 2684 2504 2692 2510
rect 2029 2384 2035 2416
rect 2541 2384 2547 2436
rect 2701 2404 2707 2496
rect 3181 2424 3187 2436
rect 1373 2344 1379 2376
rect 2605 2357 2620 2363
rect 2509 2316 2515 2356
rect 1932 2310 1940 2316
rect 2605 2304 2611 2357
rect 2669 2344 2675 2356
rect 3165 2316 3171 2336
rect 1725 2284 1731 2302
rect 1389 2144 1395 2176
rect 1213 1916 1219 1936
rect 1261 1897 1267 2096
rect 1293 1883 1299 2143
rect 1933 2137 1939 2283
rect 2573 2137 2579 2283
rect 3229 2184 3235 2256
rect 1892 2097 1900 2103
rect 1917 1984 1923 2076
rect 1357 1897 1363 1936
rect 1436 1924 1444 1930
rect 1549 1884 1555 1902
rect 1293 1877 1315 1883
rect 669 1784 675 1796
rect 1293 1743 1299 1877
rect 1869 1744 1875 1816
rect 1293 1737 1315 1743
rect 1213 1516 1219 1536
rect 1261 1524 1267 1723
rect 1436 1690 1444 1696
rect 1373 1584 1379 1636
rect 1869 1544 1875 1676
rect 1357 1497 1363 1536
rect 1436 1524 1444 1530
rect 1549 1484 1555 1502
rect 1293 1477 1315 1483
rect 701 1404 707 1436
rect 1261 1384 1267 1396
rect 1293 1344 1299 1477
rect 1869 1344 1875 1496
rect 653 1336 662 1344
rect 669 1323 675 1343
rect 653 1317 675 1323
rect 68 1117 76 1123
rect 653 1084 659 1317
rect 701 1097 707 1323
rect 653 1076 662 1084
rect 669 1063 675 1083
rect 1309 1077 1315 1343
rect 1373 1304 1379 1316
rect 1436 1290 1444 1296
rect 1373 1124 1379 1136
rect 1436 1124 1444 1130
rect 653 1057 675 1063
rect 61 937 67 956
rect 237 918 243 936
rect 77 784 83 836
rect 589 744 595 796
rect 61 664 67 683
rect 136 676 140 684
rect 621 584 627 816
rect 653 684 659 1057
rect 733 984 739 1016
rect 1293 943 1299 1076
rect 1917 984 1923 1616
rect 1949 1584 1955 1616
rect 1933 1384 1939 1536
rect 1933 1224 1939 1356
rect 1933 1184 1939 1216
rect 1293 937 1315 943
rect 1373 884 1379 896
rect 1436 890 1444 896
rect 1277 784 1283 876
rect 1373 784 1379 836
rect 1917 784 1923 956
rect 1949 784 1955 836
rect 1436 724 1444 730
rect 653 676 662 684
rect 653 563 659 676
rect 1261 584 1267 616
rect 653 557 675 563
rect 61 537 67 556
rect 653 536 662 544
rect 669 537 675 557
rect 1309 537 1315 683
rect 77 484 83 496
rect 77 384 83 436
rect 589 344 595 456
rect 653 303 659 536
rect 749 464 755 504
rect 1436 490 1444 496
rect 1373 384 1379 436
rect 1885 424 1891 476
rect 1436 324 1444 330
rect 653 297 675 303
rect 61 264 67 283
rect 669 277 675 297
rect 1965 284 1971 2116
rect 1981 1784 1987 2116
rect 2557 2104 2563 2123
rect 2628 2116 2632 2124
rect 2509 2084 2515 2104
rect 2029 1984 2035 2056
rect 2541 1984 2547 2036
rect 2509 1916 2515 1956
rect 2029 1784 2035 1896
rect 2573 1737 2579 1883
rect 2621 1784 2627 2076
rect 3181 1964 3187 2036
rect 2669 1944 2675 1956
rect 3213 1897 3219 2016
rect 3245 1883 3251 2677
rect 3261 2584 3267 2656
rect 3341 2544 3347 2616
rect 3901 2537 3907 2943
rect 4525 2937 4531 3083
rect 4541 3077 4547 3337
rect 4684 3290 4692 3296
rect 5181 3284 5187 3516
rect 4637 3144 4643 3176
rect 5213 3084 5219 3883
rect 5837 3744 5843 4283
rect 5853 4277 5859 4676
rect 6429 4604 6435 4636
rect 6461 4604 6467 4636
rect 6493 4543 6499 4936
rect 6733 4918 6739 4936
rect 6573 4884 6579 4896
rect 6541 4784 6547 4856
rect 7133 4784 7139 4836
rect 7085 4724 7091 4736
rect 7149 4703 7155 4776
rect 7133 4697 7155 4703
rect 7165 4684 7171 5337
rect 7245 5284 7251 5304
rect 7245 5116 7251 5136
rect 7789 5084 7795 5476
rect 7805 5384 7811 5436
rect 8461 5343 8467 5483
rect 8477 5384 8483 5396
rect 9117 5344 9123 5877
rect 9677 5404 9683 5436
rect 9725 5384 9731 5436
rect 9757 5344 9763 5883
rect 10317 5764 10323 5876
rect 10365 5744 10371 5956
rect 11053 5903 11059 6136
rect 11149 6084 11155 6104
rect 11836 6090 11844 6096
rect 11773 5984 11779 6036
rect 11773 5924 11779 5936
rect 11836 5924 11844 5930
rect 10557 5884 10563 5902
rect 11053 5897 11075 5903
rect 9853 5684 9859 5704
rect 9884 5690 9892 5696
rect 10381 5564 10387 5776
rect 10413 5737 10419 5883
rect 11053 5876 11062 5884
rect 11069 5877 11075 5897
rect 11053 5763 11059 5876
rect 11693 5784 11699 5916
rect 11053 5757 11075 5763
rect 11069 5737 11075 5757
rect 11149 5684 11155 5704
rect 10477 5584 10483 5636
rect 10324 5517 10332 5523
rect 10349 5497 10355 5556
rect 10989 5544 10995 5676
rect 11709 5504 11715 5883
rect 12269 5804 12275 5876
rect 12317 5804 12323 5836
rect 12333 5737 12339 6283
rect 12349 6277 12355 6677
rect 12285 5704 12291 5716
rect 11741 5544 11747 5636
rect 11836 5524 11844 5530
rect 8445 5337 8467 5343
rect 8365 5284 8371 5304
rect 7853 5097 7859 5156
rect 7725 5004 7731 5076
rect 7773 4964 7779 5036
rect 7789 4944 7795 5076
rect 8381 4964 8387 5036
rect 7389 4744 7395 4916
rect 7741 4784 7747 4836
rect 7837 4784 7843 4876
rect 7220 4737 7228 4743
rect 8365 4716 8371 4736
rect 8413 4724 8419 4956
rect 8461 4937 8467 5337
rect 8972 5290 8980 5296
rect 9037 5184 9043 5236
rect 8972 5124 8980 5130
rect 9053 5097 9059 5256
rect 9181 5204 9187 5236
rect 9661 5116 9667 5156
rect 8493 5004 8499 5036
rect 9069 4984 9075 5016
rect 9101 4944 9107 5083
rect 9117 4964 9123 5036
rect 9741 4944 9747 5343
rect 9754 5336 9763 5344
rect 9773 5304 9779 5376
rect 9837 5344 9843 5376
rect 10413 5337 10419 5483
rect 11037 5384 11043 5456
rect 10637 5318 10643 5336
rect 10477 5184 10483 5236
rect 9773 5124 9779 5176
rect 9821 5144 9827 5176
rect 11101 5124 11107 5436
rect 11133 5404 11139 5436
rect 11677 5337 11683 5483
rect 11693 5477 11715 5483
rect 11693 5337 11715 5343
rect 11693 5323 11699 5337
rect 11693 5317 11715 5323
rect 11933 5318 11939 5336
rect 12269 5324 12275 5356
rect 11613 5284 11619 5304
rect 9101 4943 9120 4944
rect 9101 4936 9123 4943
rect 8525 4904 8531 4916
rect 8525 4784 8531 4836
rect 8685 4684 8691 4702
rect 7117 4584 7123 4616
rect 6493 4537 6515 4543
rect 5885 4384 5891 4496
rect 6573 4484 6579 4496
rect 6636 4490 6644 4496
rect 6573 4384 6579 4436
rect 6461 4364 6467 4376
rect 6461 4297 6467 4356
rect 6636 4324 6644 4330
rect 6493 4277 6515 4283
rect 5869 3984 5875 4236
rect 6493 4143 6499 4277
rect 7069 4144 7075 4256
rect 7117 4184 7123 4216
rect 6493 4137 6515 4143
rect 6733 4118 6739 4136
rect 5901 3984 5907 3996
rect 6573 3984 6579 4036
rect 7085 3944 7091 4056
rect 7117 3984 7123 4016
rect 6573 3924 6579 3936
rect 6493 3877 6515 3883
rect 5933 3804 5939 3836
rect 6429 3784 6435 3816
rect 6461 3784 6467 3816
rect 6493 3744 6499 3877
rect 5757 3624 5763 3704
rect 5837 3584 5843 3676
rect 5949 3664 5955 3704
rect 5917 3636 5918 3643
rect 5917 3584 5923 3636
rect 5917 3577 5918 3584
rect 5949 3516 5955 3536
rect 5357 3464 5363 3502
rect 5853 3476 5862 3484
rect 6509 3477 6515 3743
rect 6636 3690 6644 3696
rect 6589 3510 6595 3676
rect 7069 3584 7075 3676
rect 6636 3524 6644 3530
rect 5229 3184 5235 3196
rect 5757 3116 5763 3156
rect 5821 3143 5827 3176
rect 5805 3137 5827 3143
rect 5805 3097 5811 3137
rect 4541 2937 4563 2943
rect 5213 2937 5219 3076
rect 5853 2963 5859 3476
rect 6461 3097 6467 3116
rect 6493 3083 6499 3476
rect 6589 3344 6595 3356
rect 7165 3343 7171 4676
rect 7773 4537 7779 4683
rect 7821 4584 7827 4596
rect 7885 4544 7891 4556
rect 7804 4536 7811 4544
rect 8429 4537 8435 4683
rect 8461 4543 8467 4683
rect 9021 4644 9027 4676
rect 9021 4544 9027 4616
rect 8445 4537 8467 4543
rect 7725 4344 7731 4416
rect 7805 4284 7811 4536
rect 8381 4384 8387 4436
rect 8413 4384 8419 4416
rect 7805 4276 7812 4284
rect 7805 4144 7811 4276
rect 8429 4244 8435 4510
rect 8445 4144 8451 4537
rect 8972 4324 8980 4330
rect 9037 4324 9043 4376
rect 9101 4324 9107 4356
rect 9117 4304 9123 4936
rect 9293 4764 9299 4856
rect 9709 4604 9715 4836
rect 9181 4584 9187 4596
rect 9725 4564 9731 4636
rect 9757 4544 9763 4943
rect 9981 4918 9987 4936
rect 9884 4890 9892 4896
rect 9789 4784 9795 4856
rect 9821 4744 9827 4776
rect 10333 4724 10339 4776
rect 10397 4703 10403 4756
rect 10413 4704 10419 5083
rect 11069 5063 11075 5083
rect 11053 5057 11075 5063
rect 11053 4944 11059 5057
rect 11053 4936 11062 4944
rect 11069 4923 11075 4943
rect 11053 4917 11075 4923
rect 10477 4884 10483 4896
rect 10477 4744 10483 4776
rect 10924 4724 10932 4730
rect 10957 4716 10963 4736
rect 10381 4697 10403 4703
rect 11005 4697 11011 4856
rect 11021 4744 11027 4836
rect 11053 4684 11059 4917
rect 11101 4904 11107 4923
rect 11645 4843 11651 4856
rect 11629 4837 11651 4843
rect 11629 4784 11635 4837
rect 11677 4784 11683 4816
rect 11149 4716 11155 4736
rect 9773 4584 9779 4616
rect 9661 4316 9667 4356
rect 9021 4144 9027 4216
rect 9101 4144 9107 4283
rect 9709 4184 9715 4196
rect 9741 4144 9747 4543
rect 9754 4536 9763 4544
rect 9773 4504 9779 4556
rect 9837 4544 9843 4556
rect 10397 4537 10403 4683
rect 11053 4676 11062 4684
rect 10468 4497 10476 4503
rect 10477 4384 10483 4436
rect 9821 4344 9827 4356
rect 10468 4317 10476 4323
rect 10365 4184 10371 4196
rect 10317 4144 10323 4176
rect 7805 4136 7812 4144
rect 9101 4143 9120 4144
rect 9101 4136 9123 4143
rect 7197 4004 7203 4123
rect 7245 4084 7251 4104
rect 7405 3964 7411 4056
rect 7789 3984 7795 4016
rect 7741 3944 7747 3956
rect 7773 3784 7779 3816
rect 7805 3744 7811 4136
rect 7901 4084 7907 4104
rect 8413 4024 8419 4036
rect 8365 3916 8371 3936
rect 8413 3784 8419 3816
rect 8445 3744 8451 4136
rect 8972 3924 8980 3930
rect 9117 3904 9123 4136
rect 9197 4084 9203 4104
rect 9661 3916 9667 3956
rect 8541 3884 8547 3896
rect 9757 3884 9763 4143
rect 9853 4084 9859 4104
rect 9884 4090 9892 4096
rect 9997 3904 10003 3976
rect 10381 3910 10387 4256
rect 10413 3884 10419 4283
rect 11021 4264 11027 4436
rect 11037 4284 11043 4676
rect 11053 4584 11059 4596
rect 11709 4544 11715 5317
rect 11836 5290 11844 5296
rect 11741 5184 11747 5256
rect 12285 5124 12291 5136
rect 12365 5084 12371 5736
rect 12445 5516 12451 5536
rect 12445 5284 12451 5304
rect 11933 4918 11939 4936
rect 11836 4890 11844 4896
rect 12301 4697 12307 4856
rect 12317 4744 12323 4836
rect 12365 4704 12371 5076
rect 12925 4964 12931 5276
rect 12973 5004 12979 5236
rect 12877 4944 12883 4956
rect 11741 4584 11747 4656
rect 11696 4543 11715 4544
rect 11693 4536 11715 4543
rect 12333 4537 12339 4683
rect 11613 4484 11619 4504
rect 11661 4384 11667 4396
rect 11677 4384 11683 4504
rect 11693 4304 11699 4536
rect 12285 4484 12291 4496
rect 11836 4324 11844 4330
rect 11213 4284 11219 4302
rect 11069 4263 11075 4283
rect 11053 4257 11075 4263
rect 10493 4144 10499 4216
rect 11021 4164 11027 4236
rect 11053 4144 11059 4257
rect 11709 4144 11715 4283
rect 11789 4144 11795 4176
rect 12365 4144 12371 4536
rect 12397 4184 12403 4196
rect 12429 4184 12435 4196
rect 12973 4164 12979 4236
rect 11053 4136 11062 4144
rect 10924 4090 10932 4096
rect 11149 4044 11155 4104
rect 10989 3984 10995 4036
rect 11085 3984 11091 4016
rect 10924 3924 10932 3930
rect 11613 3924 11619 3936
rect 11709 3904 11715 4136
rect 12285 4084 12291 4096
rect 11853 3884 11859 3902
rect 7805 3736 7812 3744
rect 8628 3737 8636 3743
rect 8525 3704 8531 3716
rect 7901 3684 7907 3704
rect 7725 3584 7731 3676
rect 7869 3584 7875 3636
rect 8525 3584 8531 3636
rect 9021 3564 9027 3676
rect 9069 3524 9075 3636
rect 7965 3484 7971 3502
rect 9101 3484 9107 3883
rect 9181 3784 9187 3816
rect 9181 3764 9187 3776
rect 9725 3737 9731 3883
rect 9754 3876 9763 3884
rect 9741 3737 9763 3743
rect 10413 3737 10419 3876
rect 10429 3804 10435 3836
rect 10493 3804 10499 3876
rect 11053 3763 11059 3883
rect 11661 3784 11667 3816
rect 11053 3757 11075 3763
rect 9517 3718 9523 3736
rect 7805 3476 7812 3484
rect 7149 3337 7171 3343
rect 7085 3284 7091 3296
rect 6573 3124 6579 3136
rect 6493 3077 6515 3083
rect 5853 2957 5875 2963
rect 5853 2936 5862 2944
rect 5869 2937 5875 2957
rect 5268 2897 5276 2903
rect 4684 2890 4692 2896
rect 5293 2884 5299 2904
rect 4621 2784 4627 2836
rect 5197 2764 5203 2836
rect 5277 2784 5283 2836
rect 5293 2743 5299 2836
rect 5277 2737 5299 2743
rect 4684 2724 4692 2730
rect 5277 2724 5283 2737
rect 5293 2716 5299 2737
rect 4588 2710 4596 2716
rect 4541 2677 4563 2683
rect 3981 2584 3987 2616
rect 3981 2564 3987 2576
rect 3772 2490 3780 2496
rect 3293 2384 3299 2416
rect 3837 2384 3843 2436
rect 3772 2324 3780 2330
rect 3885 2137 3891 2283
rect 3341 2124 3347 2136
rect 3772 2090 3780 2096
rect 3293 1984 3299 2036
rect 3837 1944 3843 2096
rect 3325 1924 3331 1936
rect 3917 1884 3923 2116
rect 3933 1944 3939 2436
rect 3949 2384 3955 2416
rect 4525 2137 4531 2283
rect 4541 2277 4547 2677
rect 4589 2584 4595 2596
rect 4637 2544 4643 2616
rect 5197 2537 5203 2676
rect 5773 2604 5779 2676
rect 5277 2564 5283 2576
rect 5277 2557 5278 2564
rect 4589 2384 4595 2416
rect 5133 2384 5139 2436
rect 4701 2324 4707 2376
rect 5277 2344 5283 2396
rect 5293 2344 5299 2476
rect 5805 2384 5811 2523
rect 5133 2324 5139 2336
rect 5277 2324 5283 2336
rect 5261 2297 5267 2316
rect 5853 2303 5859 2936
rect 5885 2584 5891 2856
rect 5901 2784 5907 2856
rect 5933 2784 5939 2816
rect 6413 2716 6419 2756
rect 5933 2584 5939 2616
rect 6477 2537 6483 2683
rect 6493 2677 6499 3077
rect 6541 2984 6547 3056
rect 6589 2944 6595 3016
rect 7165 2943 7171 3337
rect 7805 3344 7811 3476
rect 7805 3336 7812 3344
rect 7805 3284 7811 3296
rect 7869 3184 7875 3236
rect 7245 3116 7251 3136
rect 7901 3116 7907 3156
rect 7965 3084 7971 3102
rect 7805 3076 7812 3084
rect 7725 2944 7731 2956
rect 7149 2937 7171 2943
rect 7092 2897 7100 2903
rect 6573 2744 6579 2756
rect 7069 2716 7075 2796
rect 7085 2784 7091 2836
rect 7197 2784 7203 2856
rect 7101 2697 7107 2756
rect 7789 2744 7795 3036
rect 7709 2716 7715 2736
rect 7565 2684 7571 2702
rect 7805 2684 7811 3076
rect 7837 2984 7843 3056
rect 8461 2943 8467 3483
rect 9101 3483 9120 3484
rect 9101 3476 9123 3483
rect 9117 3344 9123 3476
rect 8972 3290 8980 3296
rect 8525 3144 8531 3276
rect 9101 3084 9107 3343
rect 9741 3343 9747 3737
rect 11053 3736 11062 3744
rect 11069 3737 11075 3757
rect 9884 3690 9892 3696
rect 10477 3684 10483 3696
rect 9997 3504 10003 3656
rect 10477 3584 10483 3636
rect 10989 3544 10995 3656
rect 11053 3503 11059 3736
rect 11149 3684 11155 3704
rect 10637 3484 10643 3502
rect 11053 3497 11075 3503
rect 9789 3364 9795 3436
rect 10381 3384 10387 3456
rect 9741 3337 9763 3343
rect 9981 3318 9987 3336
rect 9661 3284 9667 3304
rect 9709 3184 9715 3256
rect 9197 3116 9203 3136
rect 9757 3084 9763 3316
rect 9853 3284 9859 3304
rect 9884 3290 9892 3296
rect 10333 3124 10339 3176
rect 9101 3083 9120 3084
rect 9101 3076 9123 3083
rect 10397 3077 10403 3483
rect 11053 3476 11062 3484
rect 11069 3477 11075 3497
rect 10493 3344 10499 3396
rect 11053 3344 11059 3476
rect 11629 3404 11635 3436
rect 11677 3337 11683 3883
rect 11693 3877 11715 3883
rect 11741 3784 11747 3856
rect 12269 3824 12275 3876
rect 12349 3737 12355 4143
rect 12397 3984 12403 4056
rect 12941 3984 12947 4036
rect 12909 3916 12915 3936
rect 12365 3704 12371 3836
rect 12973 3737 12979 3883
rect 12765 3718 12771 3736
rect 12285 3584 12291 3636
rect 12285 3524 12291 3556
rect 12301 3497 12307 3576
rect 12381 3564 12387 3636
rect 12429 3584 12435 3636
rect 11741 3364 11747 3436
rect 11789 3404 11795 3476
rect 11693 3337 11715 3343
rect 10924 3290 10932 3296
rect 11037 3184 11043 3236
rect 10989 3144 10995 3156
rect 10477 3124 10483 3136
rect 11053 3103 11059 3336
rect 11661 3204 11667 3323
rect 11836 3290 11844 3296
rect 11773 3184 11779 3236
rect 11773 3124 11779 3136
rect 11836 3124 11844 3130
rect 11053 3097 11075 3103
rect 9069 2984 9075 3016
rect 8445 2937 8467 2943
rect 7869 2744 7875 2796
rect 8365 2716 8371 2756
rect 6493 2537 6515 2543
rect 6636 2490 6644 2496
rect 5885 2344 5891 2436
rect 6461 2384 6467 2416
rect 6573 2384 6579 2436
rect 6636 2324 6644 2330
rect 5853 2297 5875 2303
rect 4554 2136 4563 2144
rect 5181 2137 5187 2283
rect 5853 2276 5862 2284
rect 5869 2277 5875 2297
rect 7133 2284 7139 2683
rect 7229 2584 7235 2636
rect 7773 2537 7779 2683
rect 7804 2676 7811 2684
rect 8445 2544 8451 2937
rect 8516 2897 8524 2903
rect 8525 2744 8531 2756
rect 8972 2724 8980 2730
rect 9037 2724 9043 2796
rect 9101 2724 9107 2756
rect 9117 2704 9123 3076
rect 9757 2937 9763 3076
rect 9789 2964 9795 3036
rect 9853 3004 9859 3076
rect 10413 2937 10419 3083
rect 11053 3076 11062 3084
rect 11069 3077 11075 3097
rect 11853 3084 11859 3102
rect 11053 2963 11059 3076
rect 11629 2984 11635 3016
rect 11053 2957 11075 2963
rect 11069 2937 11075 2957
rect 11709 2937 11715 3083
rect 10477 2904 10483 2916
rect 9853 2884 9859 2904
rect 9884 2890 9892 2896
rect 9181 2784 9187 2796
rect 9821 2784 9827 2836
rect 10333 2744 10339 2796
rect 10477 2784 10483 2836
rect 10989 2744 10995 2836
rect 9821 2724 9827 2736
rect 9853 2724 9859 2736
rect 9884 2724 9892 2730
rect 10477 2724 10483 2736
rect 9069 2584 9075 2616
rect 9101 2544 9107 2683
rect 9741 2677 9763 2683
rect 9709 2584 9715 2596
rect 9741 2544 9747 2677
rect 10365 2584 10371 2596
rect 9101 2543 9120 2544
rect 9101 2536 9123 2543
rect 7784 2516 7788 2524
rect 8685 2518 8691 2536
rect 7741 2344 7747 2456
rect 7869 2384 7875 2436
rect 7901 2316 7907 2336
rect 8173 2304 8179 2516
rect 8429 2284 8435 2436
rect 8525 2384 8531 2436
rect 9037 2344 9043 2376
rect 5773 2144 5779 2276
rect 4461 2084 4467 2104
rect 2685 1744 2691 1856
rect 2604 1736 2611 1744
rect 3229 1737 3235 1883
rect 3245 1877 3267 1883
rect 3901 1877 3923 1884
rect 3901 1876 3920 1877
rect 2509 1684 2515 1704
rect 2541 1544 2547 1656
rect 2045 1516 2051 1536
rect 2605 1484 2611 1736
rect 3229 1584 3235 1656
rect 2628 1496 2632 1504
rect 2605 1476 2612 1484
rect 1997 1384 2003 1396
rect 2605 1344 2611 1476
rect 2605 1343 2612 1344
rect 2589 1337 2612 1343
rect 2605 1336 2612 1337
rect 2509 1284 2515 1304
rect 2557 1144 2563 1323
rect 2653 1304 2659 1323
rect 2701 1284 2707 1304
rect 2669 1184 2675 1236
rect 2045 1116 2051 1136
rect 1980 1110 1988 1116
rect 2557 1104 2563 1136
rect 2701 1116 2707 1136
rect 2557 924 2563 1096
rect 2605 1076 2612 1084
rect 2573 984 2579 996
rect 2605 944 2611 1076
rect 2605 936 2612 944
rect 2045 884 2051 904
rect 2557 844 2563 916
rect 2701 884 2707 904
rect 2669 784 2675 836
rect 3213 784 3219 1416
rect 3229 1384 3235 1536
rect 3245 1484 3251 1743
rect 3901 1737 3907 1876
rect 4045 1864 4051 1902
rect 4557 1877 4563 2136
rect 5277 2084 5283 2096
rect 4605 1924 4611 2076
rect 4621 1897 4627 2076
rect 5277 1984 5283 2036
rect 5789 2004 5795 2076
rect 5821 1984 5827 2016
rect 5789 1944 5795 1976
rect 4684 1924 4692 1930
rect 5277 1924 5283 1936
rect 3933 1784 3939 1856
rect 3981 1784 3987 1816
rect 4541 1743 4547 1876
rect 5117 1744 5123 1856
rect 5197 1784 5203 1876
rect 4541 1737 4563 1743
rect 5213 1737 5219 1883
rect 5853 1763 5859 2276
rect 5885 1984 5891 2096
rect 6493 1883 6499 2276
rect 6589 2144 6595 2176
rect 7133 2137 7139 2276
rect 7789 2144 7795 2276
rect 8381 2184 8387 2276
rect 7805 2136 7812 2144
rect 8461 2137 8467 2283
rect 9021 2144 9027 2256
rect 7784 2116 7788 2124
rect 7085 2104 7091 2116
rect 6636 1924 6644 1930
rect 6493 1877 6515 1883
rect 6429 1784 6435 1796
rect 6461 1784 6467 1816
rect 5853 1757 5875 1763
rect 5869 1737 5875 1757
rect 6493 1744 6499 1877
rect 4781 1718 4787 1736
rect 5437 1718 5443 1736
rect 3772 1690 3780 1696
rect 3325 1524 3331 1676
rect 3837 1564 3843 1696
rect 3917 1484 3923 1716
rect 5277 1704 5283 1716
rect 4461 1684 4467 1704
rect 4653 1684 4659 1704
rect 4684 1690 4692 1696
rect 5293 1664 5299 1704
rect 3933 1584 3939 1636
rect 4621 1584 4627 1636
rect 5277 1584 5283 1636
rect 4684 1524 4692 1530
rect 5277 1524 5283 1536
rect 3245 1384 3251 1416
rect 3229 984 3235 1096
rect 2541 744 2547 756
rect 2045 716 2051 736
rect 2701 716 2707 736
rect 2605 676 2612 684
rect 2573 584 2579 616
rect 2605 544 2611 676
rect 3181 584 3187 696
rect 2605 536 2612 544
rect 2628 516 2632 524
rect 2684 504 2692 510
rect 2029 384 2035 476
rect 2701 444 2707 496
rect 2669 384 2675 436
rect 2605 276 2612 284
rect 685 184 691 196
rect 701 184 707 216
rect 61 137 67 156
rect 1277 137 1283 276
rect 1325 184 1331 196
rect 1389 144 1395 156
rect 1965 143 1971 276
rect 1981 164 1987 236
rect 1949 137 1971 143
rect 2605 144 2611 276
rect 3229 144 3235 236
rect 2605 136 2612 144
rect 3261 137 3267 1483
rect 3901 1477 3923 1484
rect 3901 1476 3920 1477
rect 3901 1337 3907 1476
rect 3772 1290 3780 1296
rect 3821 1144 3827 1256
rect 3917 1084 3923 1316
rect 3901 1077 3923 1084
rect 3901 1076 3920 1077
rect 3293 984 3299 996
rect 3341 944 3347 996
rect 3901 937 3907 1076
rect 3933 984 3939 1056
rect 3981 984 3987 1016
rect 4525 984 4531 1036
rect 3933 964 3939 976
rect 4541 943 4547 1476
rect 4573 1384 4579 1416
rect 5165 1404 5171 1436
rect 4637 1344 4643 1396
rect 5197 1337 5203 1476
rect 5837 1344 5843 1736
rect 6493 1484 6499 1736
rect 6636 1690 6644 1696
rect 6573 1544 6579 1636
rect 7165 1484 7171 2116
rect 7789 1984 7795 2016
rect 7725 1944 7731 1976
rect 7805 1884 7811 2136
rect 7805 1744 7811 1876
rect 8429 1784 8435 1856
rect 7805 1736 7812 1744
rect 7245 1684 7251 1704
rect 7805 1484 7811 1736
rect 8045 1718 8051 1736
rect 7884 1704 7892 1710
rect 7837 1584 7843 1676
rect 7901 1644 7907 1696
rect 7869 1544 7875 1596
rect 8365 1516 8371 1596
rect 8413 1497 8419 1556
rect 6493 1477 6515 1484
rect 6496 1476 6515 1477
rect 7804 1476 7811 1484
rect 5901 1424 5907 1436
rect 5933 1424 5939 1436
rect 6509 1337 6515 1476
rect 7069 1344 7075 1416
rect 5133 1184 5139 1236
rect 4621 1144 4627 1176
rect 5140 1117 5148 1123
rect 4541 937 4563 943
rect 3772 890 3780 896
rect 3309 697 3315 776
rect 3837 744 3843 836
rect 3772 324 3780 330
rect 3837 324 3843 476
rect 3917 283 3923 916
rect 4461 884 4467 904
rect 4509 883 4515 923
rect 4684 890 4692 896
rect 4509 877 4531 883
rect 4525 584 4531 877
rect 4621 784 4627 836
rect 4653 716 4659 736
rect 4684 724 4692 730
rect 4461 464 4467 476
rect 3997 324 4003 336
rect 3885 277 3923 283
rect 3869 184 3875 256
rect 3885 184 3891 196
rect 4541 137 4547 676
rect 5117 624 5123 676
rect 4637 544 4643 616
rect 5181 537 5187 1083
rect 5213 724 5219 1236
rect 5229 964 5235 1256
rect 5789 1184 5795 1236
rect 5805 1224 5811 1323
rect 6573 1304 6579 1316
rect 6636 1290 6644 1296
rect 5277 1144 5283 1176
rect 5821 1110 5827 1276
rect 6429 1184 6435 1216
rect 6525 1184 6531 1256
rect 6541 1184 6547 1276
rect 6573 1144 6579 1216
rect 5949 1116 5955 1136
rect 7085 1124 7091 1156
rect 7149 1103 7155 1176
rect 7133 1097 7155 1103
rect 7165 1084 7171 1476
rect 7805 1344 7811 1476
rect 8445 1483 8451 2136
rect 8525 2084 8531 2096
rect 8493 1984 8499 2056
rect 8972 1924 8980 1930
rect 8541 1744 8547 1816
rect 9085 1743 9091 1883
rect 9117 1743 9123 2536
rect 9677 2184 9683 2256
rect 9757 2137 9763 2543
rect 9789 2384 9795 2476
rect 9853 2423 9859 2504
rect 9884 2490 9892 2496
rect 9837 2417 9859 2423
rect 9837 2344 9843 2417
rect 10413 2284 10419 2683
rect 11021 2564 11027 2836
rect 10493 2544 10499 2556
rect 11037 2544 11043 2936
rect 11293 2918 11299 2936
rect 11101 2784 11107 2896
rect 11836 2890 11844 2896
rect 11613 2716 11619 2816
rect 11773 2784 11779 2836
rect 11836 2724 11844 2730
rect 11661 2697 11667 2716
rect 11693 2677 11715 2683
rect 11629 2584 11635 2596
rect 10924 2490 10932 2496
rect 10429 2384 10435 2396
rect 10989 2384 10995 2436
rect 11053 2357 11068 2363
rect 10924 2324 10932 2330
rect 10957 2316 10963 2356
rect 11053 2304 11059 2357
rect 11613 2316 11619 2336
rect 11693 2283 11699 2677
rect 11789 2544 11795 2616
rect 12269 2604 12275 2676
rect 12349 2564 12355 2636
rect 12365 2543 12371 3476
rect 12973 3384 12979 3396
rect 12445 3284 12451 3304
rect 12925 3144 12931 3216
rect 12973 3184 12979 3216
rect 12349 2537 12371 2543
rect 12445 2484 12451 2504
rect 12285 2344 12291 2416
rect 12317 2384 12323 2456
rect 11836 2324 11844 2330
rect 10365 2184 10371 2196
rect 10317 2144 10323 2176
rect 10413 2137 10419 2276
rect 11053 2163 11059 2283
rect 11693 2277 11715 2283
rect 11053 2157 11075 2163
rect 11053 2136 11062 2144
rect 11069 2137 11075 2157
rect 11693 2144 11699 2277
rect 10637 2118 10643 2136
rect 9197 2004 9203 2104
rect 9884 2090 9892 2096
rect 9821 1984 9827 2036
rect 10349 1944 10355 1956
rect 9884 1924 9892 1930
rect 9085 1737 9123 1743
rect 8972 1690 8980 1696
rect 9037 1684 9043 1696
rect 9037 1544 9043 1576
rect 8445 1477 8467 1483
rect 8413 1384 8419 1396
rect 8429 1384 8435 1416
rect 7805 1336 7812 1344
rect 7784 1096 7788 1104
rect 7805 1084 7811 1336
rect 7885 1144 7891 1156
rect 5821 937 5827 1083
rect 6461 984 6467 1016
rect 7133 937 7139 1083
rect 7773 937 7779 1083
rect 7804 1076 7811 1084
rect 8445 1083 8451 1477
rect 9117 1343 9123 1737
rect 9341 1718 9347 1736
rect 9197 1684 9203 1696
rect 9197 1644 9203 1676
rect 9181 1584 9187 1596
rect 9661 1516 9667 1596
rect 9709 1524 9715 1836
rect 9741 1524 9747 1556
rect 9757 1503 9763 1883
rect 10397 1737 10403 2116
rect 10445 1984 10451 2036
rect 10924 1924 10932 1930
rect 10957 1916 10963 1936
rect 11053 1903 11059 2136
rect 11933 2118 11939 2136
rect 11149 2084 11155 2104
rect 11773 2084 11779 2096
rect 11836 2090 11844 2096
rect 11053 1897 11075 1903
rect 11101 1897 11107 2056
rect 11629 1984 11635 1996
rect 11773 1984 11779 2036
rect 12269 1944 12275 1956
rect 11149 1916 11155 1936
rect 11037 1737 11043 1883
rect 11053 1876 11062 1884
rect 11069 1877 11075 1897
rect 11053 1737 11059 1876
rect 11693 1743 11699 1876
rect 11693 1737 11715 1743
rect 10333 1704 10339 1716
rect 10333 1544 10339 1636
rect 10381 1584 10387 1596
rect 9884 1524 9892 1530
rect 9741 1497 9763 1503
rect 9741 1483 9747 1497
rect 9741 1477 9763 1483
rect 9741 1344 9747 1477
rect 9085 1337 9123 1343
rect 8525 1264 8531 1276
rect 7885 944 7891 956
rect 7804 936 7811 944
rect 8429 937 8435 1083
rect 8445 1077 8467 1083
rect 8461 937 8467 1077
rect 7085 904 7091 916
rect 5949 884 5955 904
rect 5277 744 5283 856
rect 5293 764 5299 876
rect 5789 784 5795 836
rect 6429 784 6435 816
rect 7085 784 7091 836
rect 7709 804 7715 904
rect 7757 803 7763 923
rect 7741 797 7763 803
rect 7741 744 7747 797
rect 7773 784 7779 796
rect 5869 737 5955 743
rect 5805 697 5811 716
rect 5869 704 5875 737
rect 5949 716 5955 737
rect 7245 716 7251 736
rect 7197 697 7203 716
rect 5853 676 5862 684
rect 5853 563 5859 676
rect 6429 584 6435 696
rect 7805 684 7811 936
rect 8221 918 8227 936
rect 8685 918 8691 936
rect 7901 716 7907 756
rect 7149 677 7171 683
rect 7133 584 7139 596
rect 5853 557 5875 563
rect 5869 537 5875 557
rect 5133 484 5139 496
rect 5277 484 5283 496
rect 5277 444 5283 476
rect 5917 436 5918 443
rect 4573 324 4579 436
rect 4621 344 4627 416
rect 5133 384 5139 436
rect 5917 384 5923 436
rect 6493 384 6499 536
rect 6636 490 6644 496
rect 6573 384 6579 436
rect 5917 377 5918 384
rect 6636 324 6644 330
rect 7133 324 7139 436
rect 5853 283 5862 284
rect 4573 184 4579 196
rect 4637 144 4643 216
rect 5181 137 5187 283
rect 5837 277 5862 283
rect 5853 276 5862 277
rect 5277 256 5278 263
rect 5277 244 5283 256
rect 5853 163 5859 276
rect 5853 157 5875 163
rect 5869 137 5875 157
rect 6589 144 6595 216
rect 7133 164 7139 236
rect 7165 143 7171 677
rect 7805 676 7812 684
rect 7789 537 7795 676
rect 8381 604 8387 636
rect 8429 564 8435 910
rect 8516 897 8524 903
rect 8525 784 8531 836
rect 9028 737 9036 743
rect 7804 536 7811 544
rect 8461 543 8467 683
rect 9085 584 9091 616
rect 9117 544 9123 1337
rect 9677 1204 9683 1236
rect 9725 1184 9731 1196
rect 9197 1116 9203 1136
rect 9197 884 9203 904
rect 9677 644 9683 656
rect 8445 537 8467 543
rect 8586 536 8588 544
rect 7565 518 7571 536
rect 7773 484 7779 510
rect 7149 137 7171 143
rect 7805 284 7811 536
rect 7869 364 7875 476
rect 8365 444 8371 496
rect 8429 484 8435 510
rect 8365 384 8371 436
rect 8525 384 8531 436
rect 9021 344 9027 456
rect 9069 384 9075 416
rect 7805 276 7812 284
rect 7805 144 7811 276
rect 7805 136 7812 144
rect 8461 137 8467 283
rect 9021 144 9027 216
rect 9069 184 9075 356
rect 9085 324 9091 496
rect 9117 137 9123 536
rect 9149 364 9155 523
rect 9693 344 9699 456
rect 9725 384 9731 636
rect 9741 584 9747 776
rect 9757 137 9763 1343
rect 10413 1337 10419 1716
rect 10924 1690 10932 1696
rect 10477 1544 10483 1576
rect 10924 1524 10932 1530
rect 10957 1524 10963 1696
rect 10989 1584 10995 1636
rect 11005 1497 11011 1723
rect 11469 1718 11475 1736
rect 11053 1476 11062 1484
rect 11053 1363 11059 1476
rect 11053 1357 11075 1363
rect 11053 1336 11062 1344
rect 11069 1337 11075 1357
rect 9981 1318 9987 1336
rect 9884 1290 9892 1296
rect 10333 1144 10339 1276
rect 10349 1123 10355 1276
rect 10340 1117 10355 1123
rect 10397 1077 10403 1316
rect 10924 1124 10932 1130
rect 10957 1116 10963 1176
rect 11005 1097 11011 1156
rect 11053 1103 11059 1336
rect 11149 1284 11155 1304
rect 11661 1224 11667 1236
rect 11053 1097 11075 1103
rect 11053 1083 11062 1084
rect 11037 1077 11062 1083
rect 11069 1077 11075 1097
rect 11053 1076 11062 1077
rect 9789 964 9795 1036
rect 10413 937 10419 1076
rect 10429 964 10435 1036
rect 11037 984 11043 1036
rect 9853 884 9859 904
rect 9884 890 9892 896
rect 10477 884 10483 896
rect 10477 784 10483 836
rect 10989 744 10995 856
rect 10333 724 10339 736
rect 10468 717 10476 723
rect 11053 703 11059 1076
rect 11133 984 11139 996
rect 11677 964 11683 1704
rect 11693 1584 11699 1616
rect 11709 1337 11715 1716
rect 11836 1690 11844 1696
rect 12285 1544 12291 1676
rect 12301 1523 12307 1676
rect 12292 1517 12307 1523
rect 11693 943 11699 1316
rect 11836 1290 11844 1296
rect 11741 1184 11747 1276
rect 12285 1144 12291 1276
rect 12301 1123 12307 1276
rect 12292 1117 12307 1123
rect 11693 937 11715 943
rect 11053 697 11075 703
rect 11101 697 11107 736
rect 11693 704 11699 796
rect 10413 537 10419 683
rect 11053 676 11062 684
rect 11069 677 11075 697
rect 11053 563 11059 676
rect 11053 557 11075 563
rect 11053 536 11062 544
rect 11069 537 11075 557
rect 9884 490 9892 496
rect 9853 204 9859 276
rect 10397 144 10403 516
rect 10924 324 10932 330
rect 10957 316 10963 376
rect 11005 324 11011 476
rect 11053 163 11059 536
rect 11677 344 11683 636
rect 11613 316 11619 336
rect 11693 324 11699 696
rect 11709 684 11715 916
rect 11836 890 11844 896
rect 12285 744 12291 876
rect 12301 723 12307 876
rect 12292 717 12307 723
rect 11709 537 11715 676
rect 11805 664 11811 676
rect 11836 490 11844 496
rect 11773 384 11779 436
rect 11836 324 11844 330
rect 11693 277 11715 283
rect 11853 264 11859 302
rect 11629 184 11635 196
rect 11677 184 11683 256
rect 11693 164 11699 256
rect 11053 157 11075 163
rect 11069 137 11075 157
rect 11789 144 11795 216
rect 12349 137 12355 1483
rect 12381 384 12387 576
rect 5437 118 5443 136
rect 6093 118 6099 136
rect 10637 118 10643 136
rect 77 104 83 116
rect 8525 104 8531 116
rect 12925 104 12931 2476
rect 93 24 99 104
rect 2701 84 2707 104
rect 3325 84 3331 96
rect 7085 84 7091 96
rect 7901 84 7907 104
rect 9884 90 9892 96
rect 11149 84 11155 104
rect 141 -43 147 16
rect 205 -43 211 16
rect 781 -43 787 16
rect 1757 -43 1763 16
rect 1805 -43 1811 16
rect 1837 -43 1843 36
rect 2749 -43 2755 16
rect 5965 -43 5971 16
rect 5997 -43 6003 16
rect 7005 -43 7011 16
rect 9213 -43 9219 16
rect 9245 -43 9251 16
<< m3contact >>
rect 6412 9016 6420 9024
rect 6444 9016 6452 9024
rect 3340 8976 3348 8984
rect 3292 8956 3300 8964
rect 10316 9016 10324 9024
rect 10348 9016 10356 9024
rect 7132 8956 7140 8964
rect 7820 8956 7828 8964
rect 8540 8956 8548 8964
rect 732 8936 740 8944
rect 1276 8916 1284 8924
rect 524 8896 532 8904
rect 556 8896 564 8904
rect 1164 8896 1172 8904
rect 1212 8876 1220 8884
rect 1212 8856 1220 8864
rect 556 8756 564 8764
rect 524 8716 532 8724
rect 732 8756 740 8764
rect 1212 8736 1220 8744
rect 1164 8716 1172 8724
rect 1196 8716 1204 8724
rect 620 8696 628 8704
rect 652 8696 660 8704
rect 1276 8696 1284 8704
rect 44 8656 52 8664
rect 44 8596 52 8604
rect 636 8596 644 8604
rect 124 8536 132 8544
rect 652 8536 660 8544
rect 1980 8936 1988 8944
rect 2684 8936 2692 8944
rect 1820 8896 1828 8904
rect 1884 8876 1892 8884
rect 1388 8836 1396 8844
rect 1340 8816 1348 8824
rect 1340 8756 1348 8764
rect 2364 8918 2372 8926
rect 2572 8916 2580 8924
rect 2620 8916 2628 8924
rect 3228 8916 3236 8924
rect 2460 8896 2468 8904
rect 2508 8896 2516 8904
rect 3116 8896 3124 8904
rect 3164 8896 3172 8904
rect 1900 8816 1908 8824
rect 1884 8756 1892 8764
rect 1820 8716 1828 8724
rect 2028 8756 2036 8764
rect 2460 8716 2468 8724
rect 2508 8716 2516 8724
rect 2716 8716 2724 8724
rect 2748 8716 2756 8724
rect 3852 8916 3860 8924
rect 3772 8896 3780 8904
rect 3900 8736 3908 8744
rect 3308 8716 3316 8724
rect 3388 8716 3396 8724
rect 2572 8696 2580 8704
rect 2764 8694 2772 8702
rect 3228 8696 3236 8704
rect 3468 8694 3476 8702
rect 3820 8696 3828 8704
rect 1324 8676 1332 8684
rect 1324 8656 1332 8664
rect 1388 8616 1396 8624
rect 140 8496 148 8504
rect 76 8476 84 8484
rect 556 8376 564 8384
rect 524 8316 532 8324
rect 620 8296 628 8304
rect 44 8196 52 8204
rect 124 8136 132 8144
rect 76 8116 84 8124
rect 140 8096 148 8104
rect 572 7936 580 7944
rect 524 7916 532 7924
rect 620 7896 628 7904
rect 92 7796 100 7804
rect 92 7776 100 7784
rect 12 7756 20 7764
rect 1164 8496 1172 8504
rect 684 8476 692 8484
rect 1212 8476 1220 8484
rect 732 8376 740 8384
rect 1260 8376 1268 8384
rect 668 8356 676 8364
rect 1212 8356 1220 8364
rect 1164 8316 1172 8324
rect 2588 8596 2596 8604
rect 2524 8576 2532 8584
rect 1900 8516 1908 8524
rect 2188 8518 2196 8526
rect 1820 8496 1828 8504
rect 2044 8496 2048 8504
rect 2048 8496 2052 8504
rect 2060 8496 2068 8504
rect 1996 8436 2004 8444
rect 1372 8356 1380 8364
rect 1884 8356 1892 8364
rect 2028 8356 2036 8364
rect 2044 8356 2052 8364
rect 1820 8316 1828 8324
rect 2460 8316 2468 8324
rect 2508 8316 2516 8324
rect 1932 8296 1940 8304
rect 1964 8296 1972 8304
rect 2572 8296 2580 8304
rect 2684 8616 2692 8624
rect 3020 8518 3028 8526
rect 3228 8516 3236 8524
rect 3116 8496 3124 8504
rect 3148 8496 3156 8504
rect 3164 8476 3172 8484
rect 3180 8456 3188 8464
rect 3228 8416 3236 8424
rect 3164 8356 3172 8364
rect 2700 8316 2708 8324
rect 2748 8316 2756 8324
rect 2676 8296 2684 8304
rect 3388 8496 3396 8504
rect 3836 8476 3844 8484
rect 3324 8456 3332 8464
rect 3836 8376 3844 8384
rect 3900 8356 3908 8364
rect 3772 8316 3780 8324
rect 4140 8918 4148 8926
rect 4476 8916 4484 8924
rect 3996 8896 4004 8904
rect 4012 8896 4020 8904
rect 4044 8896 4052 8904
rect 3996 8876 4004 8884
rect 3996 8856 4004 8864
rect 3996 8736 4004 8744
rect 4044 8716 4052 8724
rect 3932 8696 3940 8704
rect 4540 8676 4548 8684
rect 4044 8496 4052 8504
rect 3996 8476 4004 8484
rect 3980 8376 3988 8384
rect 3932 8356 3940 8364
rect 4460 8336 4468 8344
rect 4412 8316 4420 8324
rect 5196 8936 5204 8944
rect 4652 8896 4660 8904
rect 4684 8896 4692 8904
rect 4572 8756 4580 8764
rect 5068 8716 5076 8724
rect 5148 8716 5156 8724
rect 5276 8916 5284 8924
rect 6604 8936 6612 8944
rect 7884 8936 7892 8944
rect 5340 8896 5348 8904
rect 5788 8876 5796 8884
rect 5756 8776 5764 8784
rect 5180 8696 5188 8704
rect 5820 8696 5828 8704
rect 5836 8636 5844 8644
rect 5244 8596 5252 8604
rect 7772 8916 7780 8924
rect 8428 8916 8436 8924
rect 5996 8896 6004 8904
rect 6636 8896 6644 8904
rect 7660 8896 7668 8904
rect 7708 8896 7716 8904
rect 8316 8896 8324 8904
rect 8364 8896 8372 8904
rect 5948 8876 5956 8884
rect 6444 8876 6452 8884
rect 6572 8876 6580 8884
rect 5932 8776 5940 8784
rect 7148 8776 7156 8784
rect 7228 8776 7236 8784
rect 5868 8756 5876 8764
rect 6412 8756 6420 8764
rect 6572 8756 6580 8764
rect 7084 8756 7092 8764
rect 6364 8716 6372 8724
rect 7020 8716 7028 8724
rect 6508 8696 6516 8704
rect 7164 8756 7172 8764
rect 7708 8736 7716 8744
rect 7900 8736 7908 8744
rect 7660 8716 7668 8724
rect 7692 8716 7700 8724
rect 7708 8716 7716 8724
rect 7724 8716 7732 8724
rect 7884 8716 7892 8724
rect 7900 8716 7908 8724
rect 7916 8716 7924 8724
rect 7948 8716 7956 8724
rect 7564 8694 7572 8702
rect 7788 8696 7796 8704
rect 8044 8694 8052 8702
rect 7036 8676 7044 8684
rect 6428 8616 6436 8624
rect 6460 8616 6468 8624
rect 4588 8516 4596 8524
rect 5068 8496 5076 8504
rect 5916 8516 5924 8524
rect 5340 8496 5348 8504
rect 5996 8496 6004 8504
rect 5132 8476 5140 8484
rect 5148 8476 5156 8484
rect 5180 8476 5188 8484
rect 5196 8476 5204 8484
rect 5276 8476 5284 8484
rect 5948 8476 5956 8484
rect 4572 8336 4580 8344
rect 4684 8316 4692 8324
rect 4508 8296 4516 8304
rect 4780 8294 4788 8302
rect 5116 8296 5124 8304
rect 1308 8276 1316 8284
rect 1836 8276 1844 8284
rect 2588 8276 2596 8284
rect 2620 8276 2628 8284
rect 3260 8276 3268 8284
rect 3788 8276 3796 8284
rect 3916 8276 3924 8284
rect 4428 8276 4436 8284
rect 732 8116 740 8124
rect 1164 8096 1172 8104
rect 1196 8096 1204 8104
rect 1212 8096 1220 8104
rect 732 8076 740 8084
rect 1212 8076 1220 8084
rect 700 7996 708 8004
rect 1260 7996 1268 8004
rect 1260 7976 1268 7984
rect 1212 7956 1220 7964
rect 1164 7916 1172 7924
rect 1260 7796 1268 7804
rect 1276 7736 1284 7744
rect 524 7696 532 7704
rect 556 7696 564 7704
rect 588 7676 596 7684
rect 140 7516 148 7524
rect 76 7496 84 7504
rect 684 7716 692 7724
rect 748 7696 756 7704
rect 796 7696 804 7704
rect 1228 7576 1236 7584
rect 748 7516 756 7524
rect 796 7516 804 7524
rect 1532 8118 1540 8126
rect 1868 8116 1876 8124
rect 1436 8096 1444 8104
rect 1948 8076 1956 8084
rect 1372 7976 1380 7984
rect 1340 7956 1348 7964
rect 1820 7916 1828 7924
rect 1388 7896 1396 7904
rect 1932 7896 1940 7904
rect 2572 8256 2580 8264
rect 2524 8196 2532 8204
rect 1980 8116 1988 8124
rect 2092 8096 2100 8104
rect 2044 8076 2052 8084
rect 2044 7976 2052 7984
rect 2092 7916 2100 7924
rect 2188 7894 2196 7902
rect 1884 7716 1892 7724
rect 1820 7696 1828 7704
rect 1372 7536 1380 7544
rect 1932 7536 1940 7544
rect 1436 7516 1444 7524
rect 700 7496 708 7504
rect 124 7476 132 7484
rect 652 7476 660 7484
rect 28 7456 36 7464
rect 524 7296 532 7304
rect 76 7136 84 7144
rect 140 7116 148 7124
rect 204 7094 212 7102
rect 124 7076 132 7084
rect 524 6896 532 6904
rect 620 6816 628 6824
rect 604 6756 612 6764
rect 92 6736 100 6744
rect 60 6716 68 6724
rect 140 6716 148 6724
rect 156 6694 164 6702
rect 124 6676 132 6684
rect 124 6536 132 6544
rect 76 6516 84 6524
rect 236 6518 244 6526
rect 140 6496 148 6504
rect 44 6396 52 6404
rect 620 6396 628 6404
rect 556 6376 564 6384
rect 524 6316 532 6324
rect 620 6356 628 6364
rect 44 6196 52 6204
rect 92 6156 100 6164
rect 700 7396 708 7404
rect 732 7396 740 7404
rect 1548 7476 1556 7484
rect 1388 7376 1396 7384
rect 1340 7356 1348 7364
rect 1340 7336 1348 7344
rect 2028 7756 2036 7764
rect 2364 7736 2372 7744
rect 2620 8236 2628 8244
rect 2684 8136 2692 8144
rect 3020 8118 3028 8126
rect 3116 8096 3124 8104
rect 3164 8076 3172 8084
rect 2684 8056 2692 8064
rect 3212 8056 3220 8064
rect 2636 8016 2644 8024
rect 2636 7956 2644 7964
rect 3164 7936 3172 7944
rect 3116 7916 3124 7924
rect 3228 7896 3236 7904
rect 2684 7756 2692 7764
rect 3484 8118 3492 8126
rect 3820 8116 3828 8124
rect 3388 8096 3396 8104
rect 3900 8096 3908 8104
rect 3324 8016 3332 8024
rect 3836 7896 3844 7904
rect 5788 8336 5796 8344
rect 5948 8336 5956 8344
rect 5276 8316 5284 8324
rect 5340 8316 5348 8324
rect 5996 8316 6004 8324
rect 6540 8556 6548 8564
rect 7788 8556 7796 8564
rect 7020 8496 7028 8504
rect 7132 8396 7140 8404
rect 7068 8376 7076 8384
rect 6508 8316 6516 8324
rect 6604 8316 6612 8324
rect 6636 8316 6644 8324
rect 5260 8296 5268 8304
rect 6636 8294 6644 8302
rect 7388 8536 7396 8544
rect 7180 8516 7188 8524
rect 7244 8496 7248 8504
rect 7248 8496 7252 8504
rect 7260 8496 7268 8504
rect 7292 8496 7300 8504
rect 7228 8376 7236 8384
rect 7740 8476 7748 8484
rect 7708 8356 7716 8364
rect 7244 8336 7252 8344
rect 7660 8316 7668 8324
rect 7772 8296 7780 8304
rect 8380 8596 8388 8604
rect 8412 8596 8420 8604
rect 8428 8516 8436 8524
rect 8316 8496 8324 8504
rect 8364 8496 8372 8504
rect 7868 8416 7876 8424
rect 7868 8376 7876 8384
rect 7820 8356 7828 8364
rect 8316 8316 8324 8324
rect 8348 8316 8356 8324
rect 5244 8196 5252 8204
rect 5292 8196 5300 8204
rect 5212 8136 5220 8144
rect 5724 8136 5732 8144
rect 3932 8116 3940 8124
rect 4476 8116 4484 8124
rect 4620 8116 4628 8124
rect 3996 8096 4004 8104
rect 4044 8096 4052 8104
rect 4684 8096 4692 8104
rect 4476 7976 4484 7984
rect 4044 7916 4052 7924
rect 4620 7916 4628 7924
rect 4652 7916 4660 7924
rect 4668 7916 4676 7924
rect 4684 7916 4692 7924
rect 4540 7896 4548 7904
rect 2460 7696 2468 7704
rect 2492 7696 2500 7704
rect 2508 7696 2516 7704
rect 2524 7696 2532 7704
rect 3116 7696 3124 7704
rect 3148 7696 3156 7704
rect 3164 7696 3168 7704
rect 3168 7696 3172 7704
rect 1996 7636 2004 7644
rect 2028 7596 2036 7604
rect 3164 7636 3172 7644
rect 3212 7596 3220 7604
rect 2508 7576 2516 7584
rect 3180 7576 3188 7584
rect 1996 7556 2004 7564
rect 1980 7536 1988 7544
rect 2460 7516 2468 7524
rect 2748 7516 2756 7524
rect 3772 7696 3780 7704
rect 3804 7696 3812 7704
rect 3324 7676 3332 7684
rect 3852 7656 3860 7664
rect 3836 7556 3844 7564
rect 3324 7516 3332 7524
rect 3388 7516 3396 7524
rect 2364 7494 2372 7502
rect 2572 7496 2580 7504
rect 2828 7494 2836 7502
rect 3276 7496 3284 7504
rect 2028 7476 2036 7484
rect 2028 7436 2036 7444
rect 2588 7476 2596 7484
rect 2620 7476 2628 7484
rect 2684 7396 2692 7404
rect 3484 7476 3492 7484
rect 4060 7876 4068 7884
rect 4476 7816 4484 7824
rect 4508 7816 4516 7824
rect 4140 7718 4148 7726
rect 3996 7696 4004 7704
rect 4012 7696 4020 7704
rect 4044 7696 4052 7704
rect 3996 7676 4004 7684
rect 4524 7676 4532 7684
rect 4476 7576 4484 7584
rect 3996 7516 4004 7524
rect 4012 7516 4020 7524
rect 4044 7516 4052 7524
rect 4060 7494 4068 7502
rect 4524 7436 4532 7444
rect 4796 7894 4804 7902
rect 4636 7776 4644 7784
rect 5756 8096 5764 8104
rect 5276 7936 5284 7944
rect 5228 7896 5236 7904
rect 7164 8276 7172 8284
rect 7676 8276 7684 8284
rect 8220 8276 8228 8284
rect 8492 8916 8500 8924
rect 9340 8918 9348 8926
rect 8972 8896 8980 8904
rect 9052 8896 9060 8904
rect 9132 8896 9140 8904
rect 9148 8896 9156 8904
rect 9036 8876 9044 8884
rect 9244 8896 9252 8904
rect 9196 8876 9204 8884
rect 9692 8876 9700 8884
rect 8492 8756 8500 8764
rect 9708 8756 9716 8764
rect 8524 8736 8532 8744
rect 8972 8716 8980 8724
rect 9612 8716 9620 8724
rect 9068 8696 9076 8704
rect 9516 8694 9524 8702
rect 9884 8896 9892 8904
rect 9852 8876 9860 8884
rect 10396 8876 10404 8884
rect 10332 8776 10340 8784
rect 9772 8756 9780 8764
rect 10396 8756 10404 8764
rect 10268 8716 10276 8724
rect 10636 8918 10644 8926
rect 10540 8896 10548 8904
rect 10988 8876 10996 8884
rect 10476 8776 10484 8784
rect 10428 8756 10436 8764
rect 10956 8736 10964 8744
rect 10924 8716 10932 8724
rect 11004 8696 11012 8704
rect 11196 8896 11204 8904
rect 12220 8896 12228 8904
rect 11148 8876 11156 8884
rect 11676 8756 11684 8764
rect 11196 8716 11204 8724
rect 11292 8694 11300 8702
rect 8460 8576 8468 8584
rect 8540 8556 8548 8564
rect 11036 8676 11044 8684
rect 11068 8676 11076 8684
rect 10316 8616 10324 8624
rect 10364 8616 10372 8624
rect 9052 8516 9060 8524
rect 8972 8496 8980 8504
rect 9036 8476 9044 8484
rect 9068 8456 9076 8464
rect 9036 8336 9044 8344
rect 8508 8316 8516 8324
rect 8588 8316 8596 8324
rect 8476 8296 8484 8304
rect 6588 8156 6596 8164
rect 5932 8136 5940 8144
rect 6476 8116 6484 8124
rect 6364 8096 6372 8104
rect 6412 8096 6420 8104
rect 6428 8036 6436 8044
rect 5948 7936 5956 7944
rect 5996 7916 6004 7924
rect 5404 7876 5412 7884
rect 5884 7896 5892 7904
rect 6540 8116 6548 8124
rect 7020 8096 7028 8104
rect 7068 8016 7076 8024
rect 7116 8016 7124 8024
rect 6604 7916 6612 7924
rect 6636 7916 6644 7924
rect 6540 7896 6548 7904
rect 6732 7894 6740 7902
rect 6092 7876 6100 7884
rect 5276 7816 5284 7824
rect 5228 7796 5236 7804
rect 5820 7756 5828 7764
rect 4556 7736 4564 7744
rect 5084 7736 5092 7744
rect 1276 7316 1284 7324
rect 1164 7296 1172 7304
rect 1212 7296 1220 7304
rect 700 7276 708 7284
rect 1212 7156 1220 7164
rect 1164 7116 1172 7124
rect 700 7016 708 7024
rect 1900 7316 1908 7324
rect 2572 7316 2580 7324
rect 1820 7296 1828 7304
rect 2460 7296 2468 7304
rect 2492 7296 2500 7304
rect 3116 7296 3124 7304
rect 3148 7296 3156 7304
rect 3164 7296 3168 7304
rect 3168 7296 3172 7304
rect 1884 7276 1892 7284
rect 1948 7176 1956 7184
rect 2028 7176 2036 7184
rect 1372 7156 1380 7164
rect 1884 7156 1892 7164
rect 1820 7116 1828 7124
rect 1964 7156 1972 7164
rect 2460 7116 2468 7124
rect 3116 7116 3124 7124
rect 3212 7116 3220 7124
rect 2556 7096 2564 7104
rect 3020 7094 3028 7102
rect 1388 7036 1396 7044
rect 1164 6896 1172 6904
rect 1212 6876 1220 6884
rect 1164 6716 1172 6724
rect 1276 6696 1284 6704
rect 1324 6936 1332 6944
rect 2684 7016 2692 7024
rect 2620 6996 2628 7004
rect 3484 7318 3492 7326
rect 3820 7316 3828 7324
rect 3388 7296 3396 7304
rect 3884 7276 3892 7284
rect 3772 7116 3780 7124
rect 3788 7116 3796 7124
rect 3340 7096 3348 7104
rect 3868 7096 3876 7104
rect 3884 7056 3892 7064
rect 1900 6916 1908 6924
rect 1820 6896 1828 6904
rect 1884 6876 1892 6884
rect 1948 6736 1956 6744
rect 1436 6716 1444 6724
rect 1868 6696 1876 6704
rect 732 6596 740 6604
rect 1388 6576 1396 6584
rect 1340 6556 1348 6564
rect 1980 6916 1988 6924
rect 2188 6918 2196 6926
rect 2588 6916 2596 6924
rect 2636 6916 2644 6924
rect 3820 6916 3828 6924
rect 2092 6896 2100 6904
rect 2748 6896 2756 6904
rect 3388 6896 3396 6904
rect 2044 6876 2052 6884
rect 2540 6876 2548 6884
rect 2700 6876 2708 6884
rect 3196 6876 3204 6884
rect 3324 6876 3332 6884
rect 2572 6796 2580 6804
rect 3180 6756 3188 6764
rect 2044 6736 2052 6744
rect 2092 6716 2100 6724
rect 2716 6716 2724 6724
rect 2748 6716 2756 6724
rect 3388 6716 3396 6724
rect 3868 6716 3876 6724
rect 1980 6696 1988 6704
rect 2636 6696 2644 6704
rect 2812 6694 2820 6702
rect 3276 6696 3284 6704
rect 3820 6696 3828 6704
rect 2028 6596 2036 6604
rect 1276 6516 1284 6524
rect 1164 6496 1172 6504
rect 1212 6496 1220 6504
rect 684 6436 692 6444
rect 732 6376 740 6384
rect 668 6356 676 6364
rect 1212 6336 1220 6344
rect 1164 6316 1172 6324
rect 1276 6296 1284 6304
rect 684 6136 692 6144
rect 1964 6536 1972 6544
rect 2476 6536 2484 6544
rect 2588 6536 2596 6544
rect 2620 6536 2628 6544
rect 1900 6516 1908 6524
rect 1820 6496 1828 6504
rect 2460 6496 2468 6504
rect 2492 6496 2500 6504
rect 2508 6496 2516 6504
rect 2524 6496 2532 6504
rect 1884 6476 1892 6484
rect 1372 6416 1380 6424
rect 2700 6476 2708 6484
rect 3244 6476 3252 6484
rect 2556 6396 2564 6404
rect 2044 6336 2052 6344
rect 1820 6316 1828 6324
rect 2092 6316 2100 6324
rect 2748 6316 2756 6324
rect 524 6096 532 6104
rect 556 6096 564 6104
rect 1164 6096 1172 6104
rect 92 6056 100 6064
rect 44 6016 52 6024
rect 556 5936 564 5944
rect 524 5916 532 5924
rect 748 5916 756 5924
rect 796 5916 804 5924
rect 604 5896 612 5904
rect 726 5896 734 5904
rect 636 5876 644 5884
rect 668 5876 676 5884
rect 700 5816 708 5824
rect 732 5796 740 5804
rect 524 5696 532 5704
rect 12 5556 20 5564
rect 556 5596 564 5604
rect 76 5576 84 5584
rect 524 5516 532 5524
rect 556 5516 564 5524
rect 604 5496 612 5504
rect 620 5456 628 5464
rect 572 5416 580 5424
rect 44 5396 52 5404
rect 1276 5716 1284 5724
rect 1164 5696 1172 5704
rect 732 5596 740 5604
rect 1212 5536 1220 5544
rect 1164 5516 1172 5524
rect 1068 5494 1076 5502
rect 732 5376 740 5384
rect 124 5336 132 5344
rect 652 5336 660 5344
rect 1324 6136 1332 6144
rect 2188 6276 2196 6284
rect 2572 6216 2580 6224
rect 2508 6196 2516 6204
rect 2028 6176 2036 6184
rect 1964 6156 1972 6164
rect 3180 6196 3188 6204
rect 2684 6176 2692 6184
rect 2620 6156 2628 6164
rect 3820 6516 3828 6524
rect 3388 6496 3396 6504
rect 3324 6476 3332 6484
rect 3292 6456 3300 6464
rect 3932 7316 3940 7324
rect 4044 7296 4052 7304
rect 3996 7276 4004 7284
rect 3980 7196 3988 7204
rect 4412 7116 4420 7124
rect 4508 7096 4516 7104
rect 5068 7696 5076 7704
rect 5132 7676 5140 7684
rect 5148 7656 5156 7664
rect 5164 7656 5172 7664
rect 5148 7636 5156 7644
rect 4652 7576 4660 7584
rect 5180 7576 5188 7584
rect 4620 7516 4628 7524
rect 4652 7516 4660 7524
rect 4668 7516 4676 7524
rect 4684 7516 4692 7524
rect 4796 7494 4804 7502
rect 5740 7696 5748 7704
rect 6364 7696 6372 7704
rect 6396 7696 6404 7704
rect 5884 7616 5892 7624
rect 5276 7536 5284 7544
rect 5948 7536 5956 7544
rect 5996 7516 6004 7524
rect 5612 7494 5620 7502
rect 6092 7494 6100 7502
rect 5340 7356 5348 7364
rect 5836 7476 5844 7484
rect 5868 7476 5876 7484
rect 6428 7396 6436 7404
rect 6460 7396 6468 7404
rect 6732 7718 6740 7726
rect 7068 7716 7076 7724
rect 6604 7696 6612 7704
rect 7148 7696 7156 7704
rect 6540 7676 6548 7684
rect 7084 7556 7092 7564
rect 7020 7516 7028 7524
rect 7132 7496 7140 7504
rect 8428 8176 8436 8184
rect 7388 8118 7396 8126
rect 7788 8116 7796 8124
rect 7836 8116 7844 8124
rect 7260 8096 7268 8104
rect 7292 8096 7300 8104
rect 7948 8096 7956 8104
rect 7740 8076 7748 8084
rect 7900 8076 7908 8084
rect 8428 7996 8436 8004
rect 8380 7976 8388 7984
rect 7660 7916 7668 7924
rect 7692 7916 7700 7924
rect 7708 7916 7716 7924
rect 7724 7916 7732 7924
rect 7900 7916 7908 7924
rect 7948 7916 7956 7924
rect 7772 7896 7780 7904
rect 7948 7876 7956 7884
rect 7180 7836 7188 7844
rect 8428 7836 8436 7844
rect 8412 7816 8420 7824
rect 7180 7716 7188 7724
rect 7788 7716 7796 7724
rect 7836 7716 7844 7724
rect 8380 7716 8388 7724
rect 7244 7696 7252 7704
rect 7292 7696 7300 7704
rect 7756 7696 7764 7704
rect 7900 7696 7908 7704
rect 7948 7696 7956 7704
rect 8380 7636 8388 7644
rect 7180 7556 7188 7564
rect 7228 7556 7236 7564
rect 7916 7516 7924 7524
rect 7948 7516 7956 7524
rect 7756 7496 7764 7504
rect 8044 7494 8052 7502
rect 7068 7416 7076 7424
rect 5148 7316 5156 7324
rect 5212 7316 5220 7324
rect 5068 7296 5076 7304
rect 5756 7296 5764 7304
rect 5804 7296 5812 7304
rect 5132 7276 5140 7284
rect 5276 7276 5284 7284
rect 4620 7256 4628 7264
rect 4588 7216 4596 7224
rect 5116 7176 5124 7184
rect 5068 7116 5076 7124
rect 5196 7156 5204 7164
rect 5836 7156 5844 7164
rect 5340 7116 5348 7124
rect 3932 7076 3940 7084
rect 5388 7094 5396 7102
rect 5180 6976 5188 6984
rect 5772 7036 5780 7044
rect 6460 7316 6468 7324
rect 6364 7296 6372 7304
rect 6412 7296 6420 7304
rect 5932 7176 5940 7184
rect 6364 7116 6372 7124
rect 6412 7116 6420 7124
rect 6476 7096 6484 7104
rect 5868 7016 5876 7024
rect 6476 7016 6484 7024
rect 6732 7318 6740 7326
rect 6604 7296 6612 7304
rect 6636 7296 6644 7304
rect 6572 7136 6580 7144
rect 6508 7116 6516 7124
rect 7020 7116 7028 7124
rect 7100 7116 7108 7124
rect 6588 7096 6596 7104
rect 7132 7096 7140 7104
rect 7228 7396 7236 7404
rect 8380 7476 8388 7484
rect 8428 7756 8436 7764
rect 8428 7576 8436 7584
rect 7788 7336 7796 7344
rect 7820 7336 7828 7344
rect 9068 8256 9076 8264
rect 9020 8236 9028 8244
rect 8588 8096 8596 8104
rect 8524 8076 8532 8084
rect 8972 7916 8980 7924
rect 9004 7916 9012 7924
rect 9068 7896 9076 7904
rect 9132 8516 9140 8524
rect 9676 8516 9684 8524
rect 9196 8496 9204 8504
rect 9244 8496 9252 8504
rect 9708 8416 9716 8424
rect 9196 8336 9204 8344
rect 9244 8316 9252 8324
rect 9724 8216 9732 8224
rect 9164 8116 9172 8124
rect 9196 8096 9204 8104
rect 9244 8096 9252 8104
rect 9676 8016 9684 8024
rect 9740 7936 9748 7944
rect 9212 7916 9220 7924
rect 9244 7916 9252 7924
rect 9340 7894 9348 7902
rect 9068 7856 9076 7864
rect 9020 7816 9028 7824
rect 9084 7736 9092 7744
rect 8524 7716 8532 7724
rect 8588 7696 8596 7704
rect 8492 7556 8500 7564
rect 8972 7516 8980 7524
rect 8988 7516 8996 7524
rect 8540 7496 8548 7504
rect 9036 7496 9044 7504
rect 9676 7796 9684 7804
rect 9340 7736 9348 7744
rect 11772 8716 11780 8724
rect 11804 8716 11812 8724
rect 11820 8716 11828 8724
rect 11836 8716 11844 8724
rect 11692 8696 11700 8704
rect 11948 8694 11956 8702
rect 9820 8516 9828 8524
rect 10636 8518 10644 8526
rect 10972 8516 10980 8524
rect 12316 8616 12324 8624
rect 12220 8556 12228 8564
rect 9884 8496 9892 8504
rect 10540 8496 10548 8504
rect 9788 8476 9796 8484
rect 9820 8476 9828 8484
rect 11036 8476 11044 8484
rect 11004 8456 11012 8464
rect 10988 8376 10996 8384
rect 10332 8356 10340 8364
rect 11036 8336 11044 8344
rect 10268 8316 10276 8324
rect 10540 8316 10548 8324
rect 10380 8296 10388 8304
rect 10428 8296 10436 8304
rect 11084 8516 11092 8524
rect 11196 8496 11204 8504
rect 11772 8496 11780 8504
rect 11804 8496 11812 8504
rect 11820 8496 11828 8504
rect 11836 8496 11844 8504
rect 11148 8476 11156 8484
rect 11100 8376 11108 8384
rect 11148 8336 11156 8344
rect 11196 8316 11204 8324
rect 11804 8316 11812 8324
rect 11836 8316 11844 8324
rect 9772 8116 9780 8124
rect 10268 8096 10276 8104
rect 10380 8076 10388 8084
rect 10332 8016 10340 8024
rect 10316 7996 10324 8004
rect 10380 7956 10388 7964
rect 9852 7936 9860 7944
rect 9884 7916 9892 7924
rect 9788 7896 9796 7904
rect 11628 8196 11636 8204
rect 11692 8296 11700 8304
rect 10636 8136 10644 8144
rect 10540 8096 10548 8104
rect 11020 8096 11028 8104
rect 10988 8076 10996 8084
rect 10956 7936 10964 7944
rect 10924 7916 10932 7924
rect 11036 8076 11044 8084
rect 11020 8036 11028 8044
rect 10988 7896 10996 7904
rect 11148 8096 11156 8104
rect 11196 8096 11204 8104
rect 11196 7916 11204 7924
rect 11084 7896 11092 7904
rect 11788 8216 11796 8224
rect 12268 8196 12276 8204
rect 12332 8156 12340 8164
rect 12220 8096 12228 8104
rect 12284 8076 12292 8084
rect 12284 7936 12292 7944
rect 12220 7916 12228 7924
rect 12332 7896 12340 7904
rect 10412 7876 10420 7884
rect 10924 7876 10932 7884
rect 11036 7876 11044 7884
rect 11068 7876 11076 7884
rect 11292 7876 11300 7884
rect 11692 7876 11700 7884
rect 12236 7876 12244 7884
rect 9980 7736 9988 7744
rect 10316 7736 10324 7744
rect 11020 7856 11028 7864
rect 10636 7736 10644 7744
rect 9244 7696 9252 7704
rect 9884 7696 9892 7704
rect 10396 7696 10404 7704
rect 10476 7696 10484 7704
rect 10540 7696 10548 7704
rect 9196 7676 9204 7684
rect 9852 7676 9860 7684
rect 9724 7596 9732 7604
rect 9244 7516 9252 7524
rect 9340 7494 9348 7502
rect 9676 7496 9684 7504
rect 9020 7416 9028 7424
rect 8540 7396 8548 7404
rect 9084 7376 9092 7384
rect 8684 7336 8692 7344
rect 7660 7296 7668 7304
rect 7740 7156 7748 7164
rect 7292 7116 7300 7124
rect 8028 7318 8036 7326
rect 7820 7256 7828 7264
rect 7388 7094 7396 7102
rect 7756 7096 7764 7104
rect 4412 6896 4420 6904
rect 4460 6876 4468 6884
rect 4620 6916 4628 6924
rect 5436 6918 5444 6926
rect 4684 6896 4692 6904
rect 5340 6896 5348 6904
rect 5276 6876 5284 6884
rect 4476 6776 4484 6784
rect 4652 6776 4660 6784
rect 4508 6756 4516 6764
rect 3996 6716 4004 6724
rect 4044 6716 4052 6724
rect 4684 6716 4692 6724
rect 5276 6716 5284 6724
rect 5340 6716 5348 6724
rect 3900 6476 3908 6484
rect 3884 6336 3892 6344
rect 3772 6316 3780 6324
rect 3804 6316 3812 6324
rect 3868 6296 3876 6304
rect 3932 6696 3940 6704
rect 4620 6696 4628 6704
rect 5116 6696 5124 6704
rect 4524 6616 4532 6624
rect 3932 6516 3940 6524
rect 4044 6496 4052 6504
rect 3996 6476 4004 6484
rect 3996 6336 4004 6344
rect 4524 6336 4532 6344
rect 3996 6316 4004 6324
rect 4012 6316 4020 6324
rect 4044 6316 4052 6324
rect 3884 6256 3892 6264
rect 3868 6216 3876 6224
rect 3820 6196 3828 6204
rect 1884 6116 1892 6124
rect 1932 6116 1940 6124
rect 2556 6116 2564 6124
rect 1820 6096 1828 6104
rect 2460 6096 2468 6104
rect 1340 6076 1348 6084
rect 1404 6076 1412 6084
rect 2508 6076 2516 6084
rect 2588 6056 2596 6064
rect 1820 5916 1828 5924
rect 2044 5916 2048 5924
rect 2048 5916 2052 5924
rect 2060 5916 2068 5924
rect 2092 5916 2100 5924
rect 1324 5896 1332 5904
rect 1724 5894 1732 5902
rect 1932 5896 1940 5904
rect 2188 5894 2196 5902
rect 3020 6118 3028 6126
rect 3116 6096 3124 6104
rect 3148 6096 3156 6104
rect 3164 6096 3168 6104
rect 3168 6096 3172 6104
rect 2716 5916 2724 5924
rect 2748 5916 2756 5924
rect 2764 5894 2772 5902
rect 1324 5836 1332 5844
rect 1388 5816 1396 5824
rect 2684 5756 2692 5764
rect 2572 5716 2580 5724
rect 3020 5718 3028 5726
rect 1820 5696 1828 5704
rect 1900 5696 1908 5704
rect 2460 5696 2468 5704
rect 2492 5696 2500 5704
rect 3116 5696 3124 5704
rect 3148 5696 3156 5704
rect 1324 5636 1332 5644
rect 1372 5616 1380 5624
rect 1884 5536 1892 5544
rect 1820 5516 1828 5524
rect 1932 5496 1940 5504
rect 1388 5456 1396 5464
rect 140 5296 148 5304
rect 76 5276 84 5284
rect 588 5256 596 5264
rect 636 5216 644 5224
rect 636 5156 644 5164
rect 140 5116 148 5124
rect 44 4976 52 4984
rect 524 4896 532 4904
rect 556 4896 564 4904
rect 92 4856 100 4864
rect 556 4736 564 4744
rect 524 4716 532 4724
rect 92 4576 100 4584
rect 12 4556 20 4564
rect 1276 5316 1284 5324
rect 1164 5296 1172 5304
rect 684 5276 692 5284
rect 732 5196 740 5204
rect 1164 5116 1172 5124
rect 1212 5116 1220 5124
rect 1276 5096 1284 5104
rect 732 4936 740 4944
rect 1964 5396 1972 5404
rect 1900 5316 1908 5324
rect 1820 5296 1828 5304
rect 1884 5276 1892 5284
rect 1820 5116 1828 5124
rect 1900 5096 1908 5104
rect 1388 4956 1396 4964
rect 1276 4916 1284 4924
rect 1164 4896 1172 4904
rect 1212 4896 1220 4904
rect 700 4776 708 4784
rect 1212 4736 1220 4744
rect 1164 4716 1172 4724
rect 1276 4696 1284 4704
rect 732 4536 740 4544
rect 1388 4936 1396 4944
rect 1340 4916 1348 4924
rect 1884 4916 1892 4924
rect 1820 4896 1828 4904
rect 2028 5596 2036 5604
rect 2684 5596 2692 5604
rect 2636 5556 2644 5564
rect 3164 5536 3172 5544
rect 2460 5516 2468 5524
rect 2508 5516 2516 5524
rect 3116 5516 3124 5524
rect 3212 5496 3220 5504
rect 2444 5476 2452 5484
rect 2588 5336 2596 5344
rect 2620 5336 2628 5344
rect 2364 5318 2372 5326
rect 2828 5318 2836 5326
rect 2460 5296 2468 5304
rect 2492 5296 2500 5304
rect 2716 5296 2724 5304
rect 2748 5296 2756 5304
rect 2012 5256 2020 5264
rect 2028 5216 2036 5224
rect 2460 5116 2468 5124
rect 2748 5116 2756 5124
rect 2572 5096 2580 5104
rect 3180 5096 3188 5104
rect 2028 4936 2036 4944
rect 2588 5076 2596 5084
rect 2620 5076 2628 5084
rect 3228 5116 3236 5124
rect 3260 6116 3268 6124
rect 3484 6118 3492 6126
rect 3388 6096 3396 6104
rect 3852 6056 3860 6064
rect 3884 6056 3892 6064
rect 3324 5956 3332 5964
rect 3772 5916 3780 5924
rect 3852 5916 3860 5924
rect 3276 5896 3284 5904
rect 3852 5896 3860 5904
rect 5884 6916 5892 6924
rect 5996 6896 6004 6904
rect 6460 6776 6468 6784
rect 6412 6756 6420 6764
rect 6364 6716 6372 6724
rect 6732 6918 6740 6926
rect 7068 6916 7076 6924
rect 6636 6896 6644 6904
rect 7148 6876 7156 6884
rect 6572 6776 6580 6784
rect 6540 6756 6548 6764
rect 7020 6716 7028 6724
rect 7132 6696 7140 6704
rect 6924 6676 6932 6684
rect 7788 6996 7796 7004
rect 7884 7196 7892 7204
rect 7836 7176 7844 7184
rect 7948 7296 7956 7304
rect 7900 7176 7908 7184
rect 9100 7136 9108 7144
rect 8316 7116 8324 7124
rect 8588 7116 8596 7124
rect 8220 7094 8228 7102
rect 8428 7096 8436 7104
rect 8668 7094 8676 7102
rect 9020 7096 9028 7104
rect 8684 6936 8692 6944
rect 7180 6916 7188 6924
rect 8428 6916 8436 6924
rect 9020 6916 9028 6924
rect 7292 6896 7300 6904
rect 8316 6896 8324 6904
rect 8588 6896 8596 6904
rect 9100 6896 9108 6904
rect 7244 6876 7252 6884
rect 8364 6876 8372 6884
rect 9100 6876 9108 6884
rect 7724 6796 7732 6804
rect 8380 6796 8388 6804
rect 9100 6736 9108 6744
rect 7292 6716 7300 6724
rect 7948 6716 7956 6724
rect 8508 6716 8516 6724
rect 8588 6716 8596 6724
rect 8476 6696 8484 6704
rect 9020 6696 9028 6704
rect 7884 6556 7892 6564
rect 7164 6536 7172 6544
rect 7676 6536 7684 6544
rect 7836 6536 7844 6544
rect 5148 6516 5156 6524
rect 5436 6518 5444 6526
rect 5772 6516 5780 6524
rect 5884 6516 5892 6524
rect 4572 6496 4580 6504
rect 5068 6496 5076 6504
rect 5340 6496 5348 6504
rect 5996 6496 6004 6504
rect 6476 6496 6484 6504
rect 5132 6476 5140 6484
rect 5852 6476 5860 6484
rect 5948 6476 5956 6484
rect 6428 6396 6436 6404
rect 6460 6396 6468 6404
rect 5276 6356 5284 6364
rect 6428 6356 6436 6364
rect 5132 6336 5140 6344
rect 5788 6336 5796 6344
rect 5948 6336 5956 6344
rect 5068 6316 5076 6324
rect 5276 6316 5284 6324
rect 5340 6316 5348 6324
rect 5996 6316 6004 6324
rect 5180 6296 5188 6304
rect 5260 6296 5268 6304
rect 5164 6216 5172 6224
rect 4012 6096 4020 6104
rect 4044 6096 4052 6104
rect 4524 6096 4532 6104
rect 3996 5936 4004 5944
rect 4044 5916 4052 5924
rect 4476 5796 4484 5804
rect 3948 5776 3956 5784
rect 4524 5716 4532 5724
rect 4412 5696 4420 5704
rect 3836 5676 3844 5684
rect 3948 5656 3956 5664
rect 4460 5656 4468 5664
rect 4460 5596 4468 5604
rect 3772 5516 3780 5524
rect 3788 5516 3796 5524
rect 3804 5516 3812 5524
rect 3836 5516 3844 5524
rect 4412 5516 4420 5524
rect 3660 5494 3668 5502
rect 4684 6096 4692 6104
rect 4556 6076 4564 6084
rect 4652 6076 4660 6084
rect 4636 6056 4644 6064
rect 5068 5916 5076 5924
rect 5132 5916 5140 5924
rect 5180 5896 5188 5904
rect 4636 5756 4644 5764
rect 5244 6216 5252 6224
rect 5292 6216 5300 6224
rect 5756 6096 5764 6104
rect 5788 5936 5796 5944
rect 5276 5916 5284 5924
rect 5340 5916 5348 5924
rect 5932 6156 5940 6164
rect 6476 6156 6484 6164
rect 6732 6518 6740 6526
rect 6636 6496 6644 6504
rect 6572 6476 6580 6484
rect 7084 6476 7092 6484
rect 7020 6316 7028 6324
rect 7084 6316 7092 6324
rect 7100 6296 7108 6304
rect 7772 6516 7780 6524
rect 7660 6496 7668 6504
rect 7708 6496 7716 6504
rect 7180 6396 7188 6404
rect 7244 6336 7252 6344
rect 7292 6316 7300 6324
rect 7388 6294 7396 6302
rect 6588 6216 6596 6224
rect 7116 6216 7124 6224
rect 7068 6176 7076 6184
rect 7148 6156 7156 6164
rect 6460 6116 6468 6124
rect 6732 6118 6740 6126
rect 6364 6096 6372 6104
rect 6412 6096 6420 6104
rect 6636 6096 6644 6104
rect 6476 6056 6484 6064
rect 5948 5936 5956 5944
rect 6444 5936 6452 5944
rect 5996 5916 6004 5924
rect 5436 5894 5444 5902
rect 6092 5894 6100 5902
rect 6460 5896 6468 5904
rect 5820 5836 5828 5844
rect 5276 5756 5278 5764
rect 5278 5756 5284 5764
rect 6492 5916 6500 5924
rect 6604 5916 6612 5924
rect 6636 5916 6644 5924
rect 5228 5736 5236 5744
rect 5836 5736 5844 5744
rect 5868 5736 5876 5744
rect 5132 5716 5140 5724
rect 5148 5716 5156 5724
rect 5804 5716 5812 5724
rect 5068 5696 5076 5704
rect 5132 5596 5140 5604
rect 4556 5576 4564 5584
rect 4652 5556 4660 5564
rect 5180 5576 5188 5584
rect 4588 5496 4596 5504
rect 3340 5356 3348 5364
rect 3388 5356 3396 5364
rect 3980 5416 3988 5424
rect 5740 5696 5748 5704
rect 5996 5696 6004 5704
rect 5948 5676 5956 5684
rect 5276 5536 5284 5544
rect 5852 5536 5860 5544
rect 5740 5516 5748 5524
rect 6364 5516 6372 5524
rect 6412 5516 6420 5524
rect 5820 5496 5828 5504
rect 6476 5496 6484 5504
rect 6588 5816 6596 5824
rect 8220 6518 8228 6526
rect 8316 6496 8324 6504
rect 8428 6496 8436 6504
rect 7820 6436 7828 6444
rect 8364 6336 8372 6344
rect 7820 6316 7828 6324
rect 8316 6316 8324 6324
rect 8428 6296 8436 6304
rect 7228 6196 7236 6204
rect 7564 6136 7572 6144
rect 8460 6596 8468 6604
rect 9260 7476 9268 7484
rect 9164 7316 9172 7324
rect 9212 7296 9220 7304
rect 9244 7296 9252 7304
rect 9676 7256 9684 7264
rect 11036 7656 11044 7664
rect 10476 7536 10484 7544
rect 9852 7516 9860 7524
rect 10540 7516 10548 7524
rect 9740 7496 9748 7504
rect 9980 7494 9988 7502
rect 10428 7496 10436 7504
rect 11628 7836 11636 7844
rect 11628 7796 11636 7804
rect 11660 7796 11668 7804
rect 12268 7816 12276 7824
rect 11740 7756 11748 7764
rect 11932 7736 11940 7744
rect 11644 7716 11652 7724
rect 11564 7696 11572 7704
rect 11612 7696 11620 7704
rect 11836 7696 11844 7704
rect 11644 7536 11652 7544
rect 11772 7536 11780 7544
rect 11100 7516 11108 7524
rect 11148 7516 11156 7524
rect 11196 7516 11204 7524
rect 11836 7516 11844 7524
rect 9196 7136 9204 7144
rect 9692 7136 9700 7144
rect 9244 7116 9252 7124
rect 9132 7096 9140 7104
rect 9340 6936 9348 6944
rect 9132 6916 9140 6924
rect 9196 6896 9204 6904
rect 9244 6896 9252 6904
rect 9740 6876 9748 6884
rect 9708 6816 9716 6824
rect 9196 6736 9204 6744
rect 9244 6716 9252 6724
rect 9132 6696 9140 6704
rect 9132 6556 9140 6564
rect 9180 6556 9188 6564
rect 9052 6516 9060 6524
rect 8972 6496 8980 6504
rect 9004 6496 9012 6504
rect 8524 6356 8532 6364
rect 8972 6316 8980 6324
rect 9052 6296 9060 6304
rect 10364 7396 10372 7404
rect 9772 7356 9780 7364
rect 11100 7496 11108 7504
rect 10268 7296 10276 7304
rect 10332 7296 10340 7304
rect 10540 7296 10548 7304
rect 10476 7276 10484 7284
rect 11020 7236 11028 7244
rect 9852 7136 9860 7144
rect 10316 7136 10324 7144
rect 10988 7136 10996 7144
rect 9804 7116 9812 7124
rect 9884 7116 9892 7124
rect 10396 7116 10404 7124
rect 10476 7116 10484 7124
rect 10540 7116 10548 7124
rect 10316 7096 10324 7104
rect 9980 6918 9988 6926
rect 10316 6916 10324 6924
rect 9852 6896 9860 6904
rect 9884 6896 9892 6904
rect 9820 6696 9828 6704
rect 10316 6696 10324 6704
rect 10428 7096 10436 7104
rect 10972 7096 10980 7104
rect 11100 7396 11108 7404
rect 11132 7396 11140 7404
rect 11468 7336 11476 7344
rect 12268 7416 12276 7424
rect 11932 7318 11940 7326
rect 11564 7296 11572 7304
rect 11772 7296 11780 7304
rect 11804 7296 11812 7304
rect 11820 7296 11828 7304
rect 11836 7296 11844 7304
rect 11612 7256 11620 7264
rect 11148 7136 11156 7144
rect 11644 7136 11652 7144
rect 11772 7136 11780 7144
rect 11196 7116 11204 7124
rect 11676 7116 11684 7124
rect 11836 7116 11844 7124
rect 10636 6918 10644 6926
rect 10540 6896 10548 6904
rect 10988 6856 10996 6864
rect 10396 6716 10404 6724
rect 10476 6716 10484 6724
rect 10540 6716 10548 6724
rect 10428 6696 10436 6704
rect 11196 6896 11204 6904
rect 11148 6856 11156 6864
rect 11628 6756 11636 6764
rect 11196 6716 11204 6724
rect 11036 6676 11044 6684
rect 10380 6576 10388 6584
rect 9516 6536 9524 6544
rect 9180 6516 9188 6524
rect 9724 6516 9732 6524
rect 9612 6496 9620 6504
rect 9692 6336 9700 6344
rect 9244 6316 9252 6324
rect 10348 6516 10356 6524
rect 10268 6496 10276 6504
rect 9820 6476 9828 6484
rect 10332 6476 10340 6484
rect 9852 6336 9860 6344
rect 10332 6336 10340 6344
rect 9820 6316 9828 6324
rect 9884 6316 9892 6324
rect 11020 6516 11028 6524
rect 10924 6496 10932 6504
rect 10956 6496 10964 6504
rect 10476 6336 10484 6344
rect 10988 6336 10996 6344
rect 10460 6316 10468 6324
rect 10540 6316 10548 6324
rect 9340 6294 9348 6302
rect 11660 6596 11668 6604
rect 11132 6536 11140 6544
rect 11740 7056 11748 7064
rect 11708 6996 11716 7004
rect 12268 6996 12276 7004
rect 12316 6996 12324 7004
rect 12332 6956 12340 6964
rect 12220 6896 12228 6904
rect 11788 6816 11796 6824
rect 12268 6796 12276 6804
rect 12924 6796 12932 6804
rect 12444 6736 12452 6744
rect 12220 6716 12228 6724
rect 12396 6716 12404 6724
rect 12492 6716 12500 6724
rect 12124 6694 12132 6702
rect 12332 6696 12340 6704
rect 12316 6616 12324 6624
rect 11068 6516 11076 6524
rect 11660 6516 11668 6524
rect 11564 6496 11572 6504
rect 11612 6496 11620 6504
rect 11148 6336 11156 6344
rect 11196 6316 11204 6324
rect 9084 6176 9092 6184
rect 9020 6156 9028 6164
rect 7772 6116 7780 6124
rect 7660 6096 7668 6104
rect 7692 6096 7700 6104
rect 7244 5936 7252 5944
rect 7740 5936 7748 5944
rect 7292 5916 7300 5924
rect 7180 5896 7188 5904
rect 7788 5896 7796 5904
rect 8428 6116 8436 6124
rect 8316 6096 8324 6104
rect 8364 6096 8372 6104
rect 7868 6056 7876 6064
rect 8412 6016 8420 6024
rect 7836 5936 7844 5944
rect 7900 5916 7908 5924
rect 7948 5916 7956 5924
rect 7836 5896 7844 5904
rect 7180 5756 7188 5764
rect 8380 5816 8388 5824
rect 7564 5736 7572 5744
rect 7788 5736 7796 5744
rect 7820 5736 7828 5744
rect 8028 5718 8036 5726
rect 7020 5696 7028 5704
rect 7084 5696 7092 5704
rect 7660 5696 7668 5704
rect 7692 5696 7700 5704
rect 7708 5696 7716 5704
rect 7724 5696 7732 5704
rect 7948 5696 7956 5704
rect 8588 6096 8596 6104
rect 8524 6076 8532 6084
rect 8476 6056 8484 6064
rect 8972 5916 8980 5924
rect 8860 5894 8868 5902
rect 9180 6196 9188 6204
rect 9836 6176 9844 6184
rect 9724 6116 9732 6124
rect 9612 6096 9620 6104
rect 9676 6056 9684 6064
rect 11724 6476 11732 6484
rect 11836 6496 11844 6504
rect 12220 6316 12228 6324
rect 12300 6316 12308 6324
rect 12300 6296 12308 6304
rect 12316 6216 12324 6224
rect 10348 6116 10356 6124
rect 10636 6118 10644 6126
rect 10972 6116 10980 6124
rect 10268 6096 10276 6104
rect 10540 6096 10548 6104
rect 11036 6076 11044 6084
rect 10364 5956 10372 5964
rect 9852 5916 9860 5924
rect 9884 5916 9892 5924
rect 9340 5894 9348 5902
rect 9788 5896 9796 5904
rect 9980 5894 9988 5902
rect 8556 5856 8564 5864
rect 8684 5736 8692 5744
rect 8588 5696 8596 5704
rect 7900 5676 7908 5684
rect 8444 5676 8452 5684
rect 8524 5676 8532 5684
rect 7708 5636 7716 5644
rect 9068 5596 9076 5604
rect 9084 5576 9092 5584
rect 7084 5556 7092 5564
rect 7228 5556 7236 5564
rect 7756 5556 7764 5564
rect 9020 5556 9028 5564
rect 7020 5516 7028 5524
rect 7660 5516 7668 5524
rect 7708 5516 7716 5524
rect 7132 5496 7140 5504
rect 7164 5496 7172 5504
rect 7900 5536 7908 5544
rect 7948 5516 7956 5524
rect 8444 5516 8452 5524
rect 8524 5516 8532 5524
rect 8588 5516 8596 5524
rect 7836 5496 7844 5504
rect 5852 5476 5860 5484
rect 6380 5476 6388 5484
rect 5820 5436 5828 5444
rect 5772 5416 5780 5424
rect 6476 5456 6484 5464
rect 6460 5376 6468 5384
rect 3852 5316 3860 5324
rect 4508 5316 4516 5324
rect 4780 5318 4788 5326
rect 5116 5316 5124 5324
rect 5436 5318 5444 5326
rect 3772 5296 3780 5304
rect 3788 5296 3796 5304
rect 3804 5296 3812 5304
rect 3836 5296 3844 5304
rect 3884 5176 3892 5184
rect 3324 5116 3332 5124
rect 3388 5116 3396 5124
rect 3276 5096 3284 5104
rect 4412 5296 4420 5304
rect 4668 5296 4676 5304
rect 4684 5296 4692 5304
rect 5340 5296 5348 5304
rect 5836 5276 5844 5284
rect 4508 5196 4516 5204
rect 4476 5176 4484 5184
rect 3996 5136 4004 5144
rect 3996 5116 4004 5124
rect 4012 5116 4020 5124
rect 4044 5116 4052 5124
rect 4684 5116 4692 5124
rect 5276 5116 5284 5124
rect 5340 5116 5348 5124
rect 4140 5094 4148 5102
rect 4796 5094 4804 5102
rect 5436 5094 5444 5102
rect 3212 4996 3220 5004
rect 2636 4936 2644 4944
rect 2572 4916 2580 4924
rect 2460 4896 2468 4904
rect 2508 4896 2516 4904
rect 1980 4756 1988 4764
rect 1308 4736 1316 4744
rect 1884 4736 1892 4744
rect 2044 4736 2052 4744
rect 2540 4736 2548 4744
rect 1820 4716 1828 4724
rect 2060 4716 2068 4724
rect 2092 4716 2100 4724
rect 1388 4696 1396 4704
rect 1932 4696 1940 4704
rect 1980 4696 1988 4704
rect 1244 4516 1252 4524
rect 524 4496 532 4504
rect 556 4496 564 4504
rect 1164 4496 1172 4504
rect 1196 4496 1204 4504
rect 1212 4496 1220 4504
rect 76 4476 84 4484
rect 1212 4476 1220 4484
rect 44 4416 52 4424
rect 44 4356 52 4364
rect 732 4416 740 4424
rect 556 4336 564 4344
rect 524 4316 532 4324
rect 1164 4316 1172 4324
rect 620 4296 628 4304
rect 524 4096 532 4104
rect 556 4076 564 4084
rect 620 4076 628 4084
rect 572 4036 580 4044
rect 76 3916 84 3924
rect 140 3916 148 3924
rect 60 3896 68 3904
rect 2188 4676 2196 4684
rect 2028 4616 2036 4624
rect 2684 4916 2692 4924
rect 3228 4916 3236 4924
rect 3116 4896 3124 4904
rect 3148 4896 3156 4904
rect 3164 4896 3168 4904
rect 3168 4896 3172 4904
rect 2684 4816 2692 4824
rect 2684 4796 2692 4804
rect 3164 4776 3172 4784
rect 3164 4736 3172 4744
rect 3116 4716 3124 4724
rect 3228 4696 3236 4704
rect 3820 4996 3828 5004
rect 3260 4976 3268 4984
rect 3868 4956 3876 4964
rect 3980 5016 3988 5024
rect 3852 4916 3860 4924
rect 4524 4916 4532 4924
rect 3772 4896 3780 4904
rect 3804 4896 3812 4904
rect 3324 4856 3332 4864
rect 3836 4776 3844 4784
rect 3388 4716 3396 4724
rect 3484 4694 3492 4702
rect 3868 4576 3876 4584
rect 1724 4518 1732 4526
rect 1884 4516 1892 4524
rect 1820 4496 1828 4504
rect 2460 4496 2468 4504
rect 2620 4476 2628 4484
rect 1932 4456 1940 4464
rect 1340 4396 1348 4404
rect 2028 4396 2036 4404
rect 3484 4518 3492 4526
rect 3820 4516 3828 4524
rect 2700 4496 2708 4504
rect 2748 4496 2756 4504
rect 3324 4496 3332 4504
rect 3388 4496 3396 4504
rect 2652 4456 2660 4464
rect 2684 4456 2692 4464
rect 1340 4376 1348 4384
rect 3228 4356 3236 4364
rect 3884 4356 3892 4364
rect 2556 4336 2564 4344
rect 1820 4316 1828 4324
rect 1884 4316 1892 4324
rect 2460 4316 2468 4324
rect 1932 4296 1940 4304
rect 2364 4294 2372 4302
rect 3116 4316 3124 4324
rect 3340 4316 3348 4324
rect 3388 4316 3396 4324
rect 3228 4296 3236 4304
rect 3324 4296 3332 4304
rect 1388 4176 1396 4184
rect 1340 4156 1348 4164
rect 1276 4116 1284 4124
rect 1964 4196 1972 4204
rect 2028 4176 2036 4184
rect 3180 4216 3188 4224
rect 2588 4136 2596 4144
rect 2620 4136 2628 4144
rect 1164 4096 1172 4104
rect 1196 4096 1204 4104
rect 684 4056 692 4064
rect 1228 4016 1236 4024
rect 796 3916 804 3924
rect 684 3896 692 3904
rect 892 3894 900 3902
rect 124 3876 132 3884
rect 652 3876 660 3884
rect 44 3796 52 3804
rect 92 3796 100 3804
rect 892 3718 900 3726
rect 524 3696 532 3704
rect 572 3616 580 3624
rect 556 3596 564 3604
rect 636 3596 644 3604
rect 76 3516 84 3524
rect 140 3516 148 3524
rect 60 3496 68 3504
rect 124 3476 132 3484
rect 44 3396 52 3404
rect 92 3396 100 3404
rect 796 3696 804 3704
rect 1244 3676 1252 3684
rect 1212 3536 1220 3544
rect 1164 3516 1172 3524
rect 1260 3496 1268 3504
rect 1820 4096 1828 4104
rect 2460 4096 2468 4104
rect 2492 4096 2500 4104
rect 2508 4096 2516 4104
rect 2524 4096 2532 4104
rect 1372 3996 1380 4004
rect 2828 4118 2836 4126
rect 2604 4096 2612 4104
rect 2748 4096 2756 4104
rect 2700 4076 2708 4084
rect 2620 4056 2628 4064
rect 2604 4036 2612 4044
rect 2556 3976 2564 3984
rect 1884 3936 1892 3944
rect 1820 3916 1828 3924
rect 2092 3916 2100 3924
rect 1932 3896 1940 3904
rect 1436 3696 1444 3704
rect 1948 3676 1956 3684
rect 1372 3656 1380 3664
rect 1372 3576 1380 3584
rect 1820 3516 1828 3524
rect 1932 3496 1940 3504
rect 732 3336 740 3344
rect 2012 3716 2020 3724
rect 2508 3716 2516 3724
rect 2044 3696 2052 3704
rect 2092 3696 2100 3704
rect 2588 3656 2596 3664
rect 2636 4016 2644 4024
rect 3180 3956 3188 3964
rect 3116 3916 3124 3924
rect 3164 3916 3172 3924
rect 3212 3896 3220 3904
rect 3484 4118 3492 4126
rect 3820 4116 3828 4124
rect 3324 4096 3332 4104
rect 3388 4096 3396 4104
rect 3292 4036 3300 4044
rect 3324 3936 3332 3944
rect 3772 3916 3780 3924
rect 3660 3876 3668 3884
rect 4460 4856 4468 4864
rect 3948 4796 3956 4804
rect 4460 4736 4468 4744
rect 4412 4716 4420 4724
rect 4508 4696 4516 4704
rect 4588 5056 4596 5064
rect 4636 5016 4644 5024
rect 5116 4996 5124 5004
rect 5148 4916 5156 4924
rect 5068 4896 5076 4904
rect 5132 4876 5140 4884
rect 5180 4876 5188 4884
rect 5164 4776 5172 4784
rect 4620 4716 4628 4724
rect 4652 4716 4660 4724
rect 4668 4716 4676 4724
rect 4684 4716 4692 4724
rect 4796 4694 4804 4702
rect 5100 4656 5108 4664
rect 3996 4496 4004 4504
rect 4044 4496 4052 4504
rect 3980 4376 3988 4384
rect 4412 4316 4420 4324
rect 4460 4316 4468 4324
rect 4508 4316 4516 4324
rect 4604 4496 4612 4504
rect 4652 4496 4660 4504
rect 4684 4496 4692 4504
rect 5164 4336 5172 4344
rect 5068 4316 5076 4324
rect 5132 4316 5140 4324
rect 5196 4756 5204 4764
rect 5436 4936 5444 4944
rect 5436 4918 5444 4926
rect 5772 4916 5780 4924
rect 5340 4896 5348 4904
rect 6092 5318 6100 5326
rect 5996 5296 6004 5304
rect 5948 5276 5956 5284
rect 5932 5176 5940 5184
rect 6364 5116 6372 5124
rect 5868 5096 5876 5104
rect 6460 5096 6468 5104
rect 6588 5416 6596 5424
rect 7788 5476 7796 5484
rect 7820 5476 7828 5484
rect 8380 5476 8388 5484
rect 7084 5316 7092 5324
rect 7020 5296 7028 5304
rect 7148 5136 7156 5144
rect 6556 5116 6564 5124
rect 6604 5116 6612 5124
rect 6636 5116 6644 5124
rect 6732 5094 6740 5102
rect 7068 5096 7076 5104
rect 6476 4956 6484 4964
rect 7132 4976 7140 4984
rect 6732 4936 6740 4944
rect 5884 4916 5892 4924
rect 5852 4896 5860 4904
rect 5948 4896 5956 4904
rect 5996 4896 6004 4904
rect 5836 4876 5844 4884
rect 6444 4876 6452 4884
rect 5756 4756 5764 4764
rect 5900 4716 5908 4724
rect 5996 4716 6004 4724
rect 5820 4696 5828 4704
rect 6092 4694 6100 4702
rect 5820 4616 5828 4624
rect 5836 4596 5844 4604
rect 5180 4296 5188 4304
rect 4524 4216 4532 4224
rect 4476 4196 4484 4204
rect 4508 4196 4516 4204
rect 4508 4136 4516 4144
rect 3996 4096 4004 4104
rect 4044 4096 4052 4104
rect 4508 4076 4516 4084
rect 4044 3916 4052 3924
rect 4540 3916 4548 3924
rect 3868 3856 3876 3864
rect 3820 3816 3828 3824
rect 3228 3716 3236 3724
rect 3116 3696 3124 3704
rect 3148 3696 3156 3704
rect 3164 3696 3168 3704
rect 3168 3696 3172 3704
rect 2668 3656 2676 3664
rect 2092 3516 2100 3524
rect 3116 3516 3124 3524
rect 3212 3496 3220 3504
rect 1388 3356 1396 3364
rect 1276 3316 1284 3324
rect 524 3296 532 3304
rect 556 3296 564 3304
rect 1164 3296 1172 3304
rect 1212 3296 1220 3304
rect 92 3256 100 3264
rect 1340 3316 1348 3324
rect 1884 3316 1892 3324
rect 1932 3316 1940 3324
rect 1820 3296 1828 3304
rect 1884 3256 1892 3264
rect 1404 3116 1412 3124
rect 1436 3116 1444 3124
rect 1372 3096 1380 3104
rect 44 3016 52 3024
rect 636 3076 644 3084
rect 668 3076 676 3084
rect 1228 2996 1236 3004
rect 668 2956 676 2964
rect 1388 3016 1396 3024
rect 1340 2976 1348 2984
rect 620 2916 628 2924
rect 524 2896 532 2904
rect 556 2896 564 2904
rect 524 2716 532 2724
rect 556 2716 564 2724
rect 620 2696 628 2704
rect 620 2616 628 2624
rect 92 2596 100 2604
rect 636 2596 644 2604
rect 732 2936 740 2944
rect 1324 2936 1332 2944
rect 2524 3396 2532 3404
rect 2028 3356 2036 3364
rect 3388 3696 3396 3704
rect 3324 3536 3332 3544
rect 3772 3516 3780 3524
rect 4140 3718 4148 3726
rect 4044 3696 4052 3704
rect 4476 3676 4484 3684
rect 3932 3516 3940 3524
rect 3996 3516 4004 3524
rect 4044 3516 4052 3524
rect 3660 3476 3668 3484
rect 4140 3476 4148 3484
rect 5340 4496 5348 4504
rect 5244 4476 5252 4484
rect 5276 4476 5284 4484
rect 5804 4356 5812 4364
rect 5740 4316 5748 4324
rect 5804 4316 5812 4324
rect 5804 4296 5812 4304
rect 5820 4256 5828 4264
rect 5772 4196 5780 4204
rect 5148 4116 5156 4124
rect 5068 4096 5076 4104
rect 5132 4096 5140 4104
rect 5180 4056 5188 4064
rect 4604 4036 4612 4044
rect 4604 3916 4612 3924
rect 4684 3916 4692 3924
rect 4780 3894 4788 3902
rect 5116 3896 5124 3904
rect 5164 3776 5172 3784
rect 4620 3696 4628 3704
rect 4652 3696 4660 3704
rect 4668 3696 4676 3704
rect 4684 3696 4692 3704
rect 5116 3656 5124 3664
rect 4652 3636 4660 3644
rect 5340 4096 5348 4104
rect 5292 4036 5300 4044
rect 5212 3936 5220 3944
rect 5276 3936 5284 3944
rect 5340 3916 5348 3924
rect 5228 3896 5236 3904
rect 5196 3636 5204 3644
rect 4652 3516 4660 3524
rect 4684 3516 4692 3524
rect 4796 3494 4804 3502
rect 3292 3396 3300 3404
rect 1980 3336 1988 3344
rect 2588 3336 2596 3344
rect 2620 3336 2628 3344
rect 2732 3336 2740 3344
rect 3228 3336 3236 3344
rect 3244 3336 3252 3344
rect 3260 3336 3268 3344
rect 1964 3316 1972 3324
rect 2572 3316 2580 3324
rect 2668 3316 2676 3324
rect 3180 3316 3188 3324
rect 2460 3296 2468 3304
rect 2716 3296 2724 3304
rect 2748 3296 2756 3304
rect 2508 3276 2516 3284
rect 2508 3256 2516 3264
rect 2028 3156 2036 3164
rect 2620 3156 2628 3164
rect 3228 3136 3236 3144
rect 2460 3116 2468 3124
rect 2492 3116 2500 3124
rect 2508 3116 2516 3124
rect 2524 3116 2532 3124
rect 2572 3096 2580 3104
rect 3084 3094 3092 3102
rect 1068 2918 1076 2926
rect 1164 2896 1172 2904
rect 1260 2776 1268 2784
rect 668 2756 676 2764
rect 1212 2756 1220 2764
rect 1164 2716 1172 2724
rect 732 2576 740 2584
rect 124 2536 132 2544
rect 652 2536 660 2544
rect 1900 2916 1908 2924
rect 1820 2896 1828 2904
rect 1884 2876 1892 2884
rect 2524 2916 2532 2924
rect 2044 2896 2048 2904
rect 2048 2896 2052 2904
rect 2060 2896 2068 2904
rect 2092 2896 2100 2904
rect 2044 2876 2052 2884
rect 2588 2876 2596 2884
rect 2012 2856 2020 2864
rect 2028 2796 2036 2804
rect 1372 2776 1380 2784
rect 1340 2756 1348 2764
rect 2508 2736 2516 2744
rect 1820 2716 1828 2724
rect 1900 2696 1908 2704
rect 2636 2916 2644 2924
rect 2748 2896 2756 2904
rect 2700 2876 2708 2884
rect 2684 2776 2692 2784
rect 2636 2756 2644 2764
rect 3116 2716 3124 2724
rect 3182 2696 3190 2704
rect 1388 2616 1396 2624
rect 76 2516 84 2524
rect 140 2496 148 2504
rect 620 2416 628 2424
rect 636 2356 644 2364
rect 76 2336 84 2344
rect 140 2316 148 2324
rect 140 2294 148 2302
rect 44 2216 52 2224
rect 524 2096 532 2104
rect 556 2096 564 2104
rect 92 2036 100 2044
rect 44 1996 52 2004
rect 556 1936 564 1944
rect 524 1916 532 1924
rect 620 1896 628 1904
rect 44 1796 52 1804
rect 620 1716 628 1724
rect 524 1696 532 1704
rect 556 1676 564 1684
rect 44 1596 52 1604
rect 556 1536 564 1544
rect 524 1516 532 1524
rect 620 1456 628 1464
rect 636 1416 644 1424
rect 236 1318 244 1326
rect 140 1296 148 1304
rect 1276 2516 1284 2524
rect 1164 2496 1172 2504
rect 1212 2476 1220 2484
rect 1260 2376 1268 2384
rect 1212 2356 1220 2364
rect 1164 2316 1172 2324
rect 732 2136 740 2144
rect 2028 2536 2036 2544
rect 3324 3296 3332 3304
rect 3340 3296 3348 3304
rect 3388 3296 3396 3304
rect 3292 3276 3300 3284
rect 3276 3156 3284 3164
rect 3772 3116 3780 3124
rect 3660 3094 3668 3102
rect 3868 3096 3876 3104
rect 3356 3056 3364 3064
rect 3292 3016 3300 3024
rect 3916 3456 3924 3464
rect 3932 3436 3940 3444
rect 3948 3416 3956 3424
rect 3932 3296 3940 3304
rect 3980 3396 3988 3404
rect 4316 3318 4324 3326
rect 3980 3276 3988 3284
rect 4508 3276 4516 3284
rect 4460 3156 4468 3164
rect 4412 3116 4420 3124
rect 4524 3096 4532 3104
rect 3980 3016 3988 3024
rect 3836 2876 3844 2884
rect 3324 2756 3332 2764
rect 3852 2856 3860 2864
rect 3388 2716 3396 2724
rect 3276 2696 3284 2704
rect 3484 2694 3492 2702
rect 2588 2536 2596 2544
rect 2620 2536 2628 2544
rect 1820 2496 1828 2504
rect 1884 2476 1892 2484
rect 1916 2516 1924 2524
rect 2460 2496 2468 2504
rect 2508 2476 2516 2484
rect 2844 2518 2852 2526
rect 2684 2496 2692 2504
rect 2700 2496 2708 2504
rect 2716 2496 2724 2504
rect 2748 2496 2756 2504
rect 2556 2456 2564 2464
rect 2028 2416 2036 2424
rect 1900 2396 1908 2404
rect 3180 2416 3188 2424
rect 2700 2396 2708 2404
rect 1372 2376 1380 2384
rect 1340 2356 1348 2364
rect 2508 2356 2516 2364
rect 1820 2316 1828 2324
rect 1932 2316 1940 2324
rect 2460 2316 2468 2324
rect 2668 2356 2676 2364
rect 3164 2336 3172 2344
rect 3116 2316 3124 2324
rect 2572 2296 2580 2304
rect 2604 2296 2612 2304
rect 3228 2296 3236 2304
rect 1724 2276 1732 2284
rect 1388 2176 1396 2184
rect 1260 2116 1268 2124
rect 1164 2096 1172 2104
rect 1196 2096 1204 2104
rect 1260 2096 1268 2104
rect 732 1956 740 1964
rect 1212 1936 1220 1944
rect 1164 1916 1172 1924
rect 1276 1916 1284 1924
rect 2028 2156 2036 2164
rect 1980 2136 1988 2144
rect 3228 2256 3236 2264
rect 2588 2136 2596 2144
rect 2620 2136 2628 2144
rect 1900 2116 1908 2124
rect 1980 2116 1988 2124
rect 1820 2096 1828 2104
rect 1900 2096 1908 2104
rect 1916 2076 1924 2084
rect 1356 1936 1364 1944
rect 1404 1916 1412 1924
rect 1436 1916 1444 1924
rect 668 1796 676 1804
rect 732 1756 740 1764
rect 1548 1876 1556 1884
rect 1868 1816 1876 1824
rect 716 1536 724 1544
rect 1212 1536 1220 1544
rect 1164 1516 1172 1524
rect 1276 1716 1284 1724
rect 1372 1696 1380 1704
rect 1404 1696 1412 1704
rect 1420 1696 1428 1704
rect 1436 1696 1444 1704
rect 1868 1676 1876 1684
rect 1916 1616 1924 1624
rect 1948 1616 1956 1624
rect 1356 1536 1364 1544
rect 1260 1516 1268 1524
rect 1276 1496 1284 1504
rect 1420 1516 1428 1524
rect 1436 1516 1444 1524
rect 1868 1496 1876 1504
rect 732 1436 740 1444
rect 700 1396 708 1404
rect 1260 1396 1268 1404
rect 1548 1476 1556 1484
rect 60 1116 68 1124
rect 140 1116 148 1124
rect 684 1316 692 1324
rect 796 1296 804 1304
rect 1292 1156 1300 1164
rect 1244 1136 1252 1144
rect 796 1116 804 1124
rect 60 1076 68 1084
rect 1372 1316 1380 1324
rect 1532 1318 1540 1326
rect 1436 1296 1444 1304
rect 1372 1136 1380 1144
rect 1436 1116 1444 1124
rect 1548 1094 1556 1102
rect 60 956 68 964
rect 236 936 244 944
rect 76 896 84 904
rect 140 896 148 904
rect 620 816 628 824
rect 588 796 596 804
rect 140 716 148 724
rect 76 696 84 704
rect 140 676 148 684
rect 60 656 68 664
rect 636 776 644 784
rect 732 1016 740 1024
rect 1932 1536 1940 1544
rect 1932 1356 1940 1364
rect 1932 1216 1940 1224
rect 1916 956 1924 964
rect 1276 916 1284 924
rect 1164 896 1172 904
rect 1196 896 1204 904
rect 1436 896 1444 904
rect 684 876 692 884
rect 1276 876 1284 884
rect 1372 876 1380 884
rect 1948 776 1956 784
rect 764 716 772 724
rect 796 716 804 724
rect 1420 716 1428 724
rect 1436 716 1444 724
rect 892 694 900 702
rect 1548 694 1556 702
rect 668 676 676 684
rect 60 556 68 564
rect 1260 616 1268 624
rect 236 518 244 526
rect 76 496 84 504
rect 140 496 148 504
rect 76 476 84 484
rect 588 456 596 464
rect 636 356 644 364
rect 92 316 100 324
rect 140 316 148 324
rect 892 518 900 526
rect 1532 518 1540 526
rect 796 496 804 504
rect 1404 496 1412 504
rect 1436 496 1444 504
rect 748 456 756 464
rect 1884 416 1892 424
rect 764 316 772 324
rect 796 316 804 324
rect 1404 316 1412 324
rect 1436 316 1444 324
rect 726 296 734 304
rect 892 294 900 302
rect 1340 296 1348 304
rect 1548 294 1556 302
rect 2620 2116 2628 2124
rect 2844 2118 2852 2126
rect 2460 2096 2468 2104
rect 2556 2096 2564 2104
rect 2716 2096 2724 2104
rect 2748 2096 2756 2104
rect 2508 2076 2516 2084
rect 2620 2076 2628 2084
rect 2028 2056 2036 2064
rect 2508 1956 2516 1964
rect 2460 1916 2468 1924
rect 2028 1896 2036 1904
rect 3212 2016 3220 2024
rect 2668 1956 2676 1964
rect 3180 1956 3188 1964
rect 3116 1916 3124 1924
rect 3182 1896 3190 1904
rect 3260 2656 3268 2664
rect 3340 2616 3348 2624
rect 4668 3296 4676 3304
rect 4684 3296 4692 3304
rect 5180 3276 5188 3284
rect 4636 3176 4644 3184
rect 4588 3156 4596 3164
rect 5068 3116 5076 3124
rect 4636 3096 4644 3104
rect 4972 3094 4980 3102
rect 5180 3096 5188 3104
rect 6428 4596 6436 4604
rect 6460 4596 6468 4604
rect 6572 4876 6580 4884
rect 6540 4856 6548 4864
rect 7132 4776 7140 4784
rect 7148 4776 7156 4784
rect 7084 4736 7092 4744
rect 7020 4716 7028 4724
rect 7212 5316 7220 5324
rect 7292 5296 7300 5304
rect 7244 5276 7252 5284
rect 7740 5276 7748 5284
rect 7244 5136 7252 5144
rect 7292 5116 7300 5124
rect 7180 5096 7188 5104
rect 7804 5436 7812 5444
rect 8412 5436 8420 5444
rect 8604 5476 8612 5484
rect 8476 5396 8484 5404
rect 9340 5718 9348 5726
rect 9244 5696 9252 5704
rect 9740 5676 9748 5684
rect 9244 5516 9252 5524
rect 9132 5496 9140 5504
rect 9340 5494 9348 5502
rect 9676 5396 9684 5404
rect 9724 5376 9732 5384
rect 10316 5756 10324 5764
rect 10988 5936 10996 5944
rect 10396 5916 10404 5924
rect 10540 5916 10548 5924
rect 11084 6116 11092 6124
rect 11692 6116 11700 6124
rect 11196 6096 11204 6104
rect 11804 6096 11812 6104
rect 11836 6096 11844 6104
rect 11148 6076 11156 6084
rect 11644 5936 11652 5944
rect 11772 5936 11780 5944
rect 11148 5916 11156 5924
rect 11196 5916 11204 5924
rect 11692 5916 11700 5924
rect 11836 5916 11844 5924
rect 10636 5894 10644 5902
rect 10380 5776 10388 5784
rect 10316 5736 10324 5744
rect 10364 5736 10372 5744
rect 9884 5696 9892 5704
rect 9852 5676 9860 5684
rect 10556 5876 10564 5884
rect 11260 5894 11268 5902
rect 10636 5718 10644 5726
rect 10972 5716 10980 5724
rect 11084 5716 11092 5724
rect 10540 5696 10548 5704
rect 11196 5696 11204 5704
rect 10988 5676 10996 5684
rect 11052 5676 11060 5684
rect 11148 5676 11156 5684
rect 10348 5556 10356 5564
rect 10380 5556 10388 5564
rect 10268 5516 10276 5524
rect 10316 5516 10324 5524
rect 10540 5516 10548 5524
rect 11564 5516 11572 5524
rect 12268 5796 12276 5804
rect 12316 5796 12324 5804
rect 12284 5716 12292 5724
rect 12300 5716 12308 5724
rect 12220 5696 12228 5704
rect 11740 5536 11748 5544
rect 12284 5536 12292 5544
rect 11804 5516 11812 5524
rect 11836 5516 11844 5524
rect 10428 5496 10436 5504
rect 11468 5494 11476 5502
rect 11868 5494 11876 5502
rect 9772 5376 9780 5384
rect 9836 5376 9844 5384
rect 8428 5316 8436 5324
rect 8316 5296 8324 5304
rect 8364 5276 8372 5284
rect 7852 5156 7860 5164
rect 7948 5116 7956 5124
rect 7788 5076 7796 5084
rect 7820 5076 7828 5084
rect 7724 4996 7732 5004
rect 7772 4956 7780 4964
rect 8380 4956 8388 4964
rect 8412 4956 8420 4964
rect 7788 4936 7796 4944
rect 7820 4936 7828 4944
rect 7388 4916 7396 4924
rect 7772 4916 7780 4924
rect 7836 4916 7844 4924
rect 8380 4916 8388 4924
rect 7180 4776 7188 4784
rect 7660 4896 7668 4904
rect 7708 4896 7716 4904
rect 7900 4896 7908 4904
rect 7948 4896 7956 4904
rect 7836 4876 7844 4884
rect 7228 4736 7236 4744
rect 7388 4736 7396 4744
rect 8364 4736 8372 4744
rect 7660 4716 7668 4724
rect 7708 4716 7716 4724
rect 8316 4716 8324 4724
rect 9052 5316 9060 5324
rect 8972 5296 8980 5304
rect 9004 5296 9012 5304
rect 9612 5296 9620 5304
rect 9660 5296 9668 5304
rect 9052 5256 9060 5264
rect 9116 5256 9124 5264
rect 8972 5116 8980 5124
rect 9004 5116 9012 5124
rect 9180 5196 9188 5204
rect 9660 5156 9668 5164
rect 9612 5116 9620 5124
rect 9068 5016 9076 5024
rect 8492 4996 8500 5004
rect 9116 4956 9124 4964
rect 9788 5356 9796 5364
rect 11036 5456 11044 5464
rect 10636 5336 10644 5344
rect 10348 5316 10356 5324
rect 10268 5296 10276 5304
rect 10540 5296 10548 5304
rect 10988 5276 10996 5284
rect 9772 5176 9780 5184
rect 9820 5176 9828 5184
rect 9788 5156 9796 5164
rect 10988 5136 10996 5144
rect 11132 5396 11140 5404
rect 12268 5356 12276 5364
rect 11676 5316 11684 5324
rect 11932 5336 11940 5344
rect 11564 5296 11572 5304
rect 11612 5276 11620 5284
rect 10268 5116 10276 5124
rect 10540 5116 10548 5124
rect 11100 5116 11108 5124
rect 11148 5116 11156 5124
rect 11196 5116 11204 5124
rect 10172 5094 10180 5102
rect 10380 5096 10388 5104
rect 10572 5094 10580 5102
rect 11126 5096 11134 5104
rect 8524 4916 8532 4924
rect 8588 4896 8596 4904
rect 8412 4716 8420 4724
rect 8588 4716 8596 4724
rect 7772 4696 7780 4704
rect 8428 4696 8436 4704
rect 8476 4696 8484 4704
rect 7116 4616 7124 4624
rect 6444 4516 6452 4524
rect 6732 4518 6740 4526
rect 5884 4496 5892 4504
rect 6364 4496 6372 4504
rect 6412 4496 6420 4504
rect 6636 4496 6644 4504
rect 6572 4476 6580 4484
rect 6460 4376 6468 4384
rect 6460 4356 6468 4364
rect 6364 4316 6372 4324
rect 6396 4316 6404 4324
rect 6412 4316 6420 4324
rect 6636 4316 6644 4324
rect 6732 4294 6740 4302
rect 5868 4236 5876 4244
rect 5932 4156 5940 4164
rect 7068 4276 7076 4284
rect 7068 4256 7076 4264
rect 7116 4216 7124 4224
rect 7116 4176 7124 4184
rect 6732 4136 6740 4144
rect 6460 4116 6468 4124
rect 6364 4096 6372 4104
rect 6412 4096 6420 4104
rect 6636 4096 6644 4104
rect 7084 4056 7092 4064
rect 5900 3996 5908 4004
rect 7116 4016 7124 4024
rect 6572 3936 6580 3944
rect 6364 3916 6372 3924
rect 6396 3916 6404 3924
rect 6636 3916 6644 3924
rect 6476 3896 6484 3904
rect 6428 3816 6436 3824
rect 6460 3816 6468 3824
rect 5932 3796 5940 3804
rect 5836 3736 5844 3744
rect 5868 3736 5876 3744
rect 5804 3716 5812 3724
rect 5836 3676 5844 3684
rect 5756 3616 5764 3624
rect 5996 3696 6004 3704
rect 5948 3656 5956 3664
rect 5948 3536 5956 3544
rect 5340 3516 5348 3524
rect 5996 3516 6004 3524
rect 6492 3516 6500 3524
rect 6428 3496 6436 3504
rect 6604 3696 6612 3704
rect 6636 3696 6644 3704
rect 6588 3676 6596 3684
rect 6572 3516 6580 3524
rect 7068 3576 7076 3584
rect 6604 3516 6612 3524
rect 6620 3516 6628 3524
rect 6636 3516 6644 3524
rect 6540 3496 6548 3504
rect 5356 3456 5364 3464
rect 5228 3336 5236 3344
rect 5228 3196 5236 3204
rect 5820 3176 5828 3184
rect 5756 3156 5764 3164
rect 5116 2936 5124 2944
rect 5868 3376 5876 3384
rect 6476 3316 6484 3324
rect 6364 3296 6372 3304
rect 6412 3296 6420 3304
rect 5932 3176 5940 3184
rect 5868 3156 5876 3164
rect 6364 3116 6372 3124
rect 6412 3116 6420 3124
rect 6460 3116 6468 3124
rect 7132 3436 7140 3444
rect 6588 3356 6596 3364
rect 7228 4556 7236 4564
rect 7820 4596 7828 4604
rect 7884 4556 7892 4564
rect 8684 4676 8692 4684
rect 9020 4636 9028 4644
rect 9020 4616 9028 4624
rect 9084 4556 9092 4564
rect 7756 4516 7764 4524
rect 7660 4496 7668 4504
rect 7724 4416 7732 4424
rect 7292 4316 7300 4324
rect 7388 4294 7396 4302
rect 7788 4296 7796 4304
rect 8428 4516 8436 4524
rect 8316 4496 8324 4504
rect 8364 4496 8372 4504
rect 8380 4436 8388 4444
rect 8412 4416 8420 4424
rect 7900 4316 7908 4324
rect 7948 4316 7956 4324
rect 7876 4296 7884 4304
rect 8428 4236 8436 4244
rect 8684 4518 8692 4526
rect 9036 4376 9044 4384
rect 9100 4356 9108 4364
rect 8972 4316 8980 4324
rect 9244 4896 9252 4904
rect 9292 4856 9300 4864
rect 9292 4756 9300 4764
rect 9244 4716 9252 4724
rect 9340 4694 9348 4702
rect 9180 4596 9188 4604
rect 9708 4596 9716 4604
rect 9724 4556 9732 4564
rect 9980 4936 9988 4944
rect 9884 4896 9892 4904
rect 10396 4876 10404 4884
rect 9788 4856 9796 4864
rect 9820 4776 9828 4784
rect 10332 4776 10340 4784
rect 10396 4756 10404 4764
rect 10268 4716 10276 4724
rect 11628 4936 11636 4944
rect 10540 4896 10548 4904
rect 10476 4876 10484 4884
rect 11004 4856 11012 4864
rect 10476 4776 10484 4784
rect 10428 4756 10436 4764
rect 10956 4736 10964 4744
rect 10924 4716 10932 4724
rect 11020 4736 11028 4744
rect 11100 4896 11108 4904
rect 11196 4896 11204 4904
rect 11692 4896 11700 4904
rect 11628 4856 11636 4864
rect 11644 4856 11652 4864
rect 11660 4836 11668 4844
rect 11676 4816 11684 4824
rect 11148 4736 11156 4744
rect 11196 4716 11204 4724
rect 11116 4696 11124 4704
rect 9772 4616 9780 4624
rect 9772 4556 9780 4564
rect 9836 4556 9844 4564
rect 9612 4496 9620 4504
rect 9660 4496 9668 4504
rect 9180 4376 9188 4384
rect 9132 4356 9140 4364
rect 9660 4356 9668 4364
rect 9612 4316 9620 4324
rect 8492 4256 8500 4264
rect 9020 4216 9028 4224
rect 9708 4196 9716 4204
rect 11036 4676 11044 4684
rect 11068 4676 11076 4684
rect 10348 4516 10356 4524
rect 10268 4496 10276 4504
rect 10460 4496 10468 4504
rect 10540 4496 10548 4504
rect 9820 4356 9828 4364
rect 10268 4316 10276 4324
rect 10332 4316 10340 4324
rect 10460 4316 10468 4324
rect 10540 4316 10548 4324
rect 10348 4296 10356 4304
rect 10476 4296 10484 4304
rect 10380 4256 10388 4264
rect 10364 4196 10372 4204
rect 10316 4176 10324 4184
rect 7724 4116 7732 4124
rect 7292 4096 7300 4104
rect 7244 4076 7252 4084
rect 7788 4076 7796 4084
rect 7404 4056 7412 4064
rect 7196 3996 7204 4004
rect 7788 4016 7796 4024
rect 7404 3956 7412 3964
rect 7740 3956 7748 3964
rect 7292 3916 7300 3924
rect 7388 3894 7396 3902
rect 7772 3816 7780 3824
rect 7836 4116 7844 4124
rect 7948 4096 7956 4104
rect 7900 4076 7908 4084
rect 8412 4016 8420 4024
rect 8364 3936 8372 3944
rect 8316 3916 8324 3924
rect 8428 3896 8436 3904
rect 8412 3816 8420 3824
rect 8380 3776 8388 3784
rect 8588 4096 8596 4104
rect 8460 3936 8468 3944
rect 8972 3916 8980 3924
rect 9132 4116 9140 4124
rect 9244 4096 9252 4104
rect 9196 4076 9204 4084
rect 9132 3956 9140 3964
rect 9660 3956 9668 3964
rect 9612 3916 9620 3924
rect 8540 3896 8548 3904
rect 8860 3894 8868 3902
rect 9084 3896 9092 3904
rect 9724 3896 9732 3904
rect 9980 4118 9988 4126
rect 9884 4096 9892 4104
rect 9852 4076 9860 4084
rect 9996 3976 10004 3984
rect 9788 3956 9796 3964
rect 10268 3916 10276 3924
rect 9836 3896 9844 3904
rect 10172 3894 10180 3902
rect 11052 4596 11060 4604
rect 12268 5316 12276 5324
rect 11804 5296 11812 5304
rect 11836 5296 11844 5304
rect 12348 5276 12356 5284
rect 11740 5256 11748 5264
rect 12284 5136 12292 5144
rect 11724 5116 11732 5124
rect 12220 5116 12228 5124
rect 12332 5096 12340 5104
rect 12972 5556 12980 5564
rect 12444 5536 12452 5544
rect 12492 5516 12500 5524
rect 12380 5316 12388 5324
rect 12492 5296 12500 5304
rect 12444 5276 12452 5284
rect 11932 4936 11940 4944
rect 11804 4896 11812 4904
rect 11836 4896 11844 4904
rect 12300 4856 12308 4864
rect 12220 4716 12228 4724
rect 12284 4716 12292 4724
rect 11724 4696 11732 4704
rect 12316 4736 12324 4744
rect 12972 4996 12980 5004
rect 12972 4976 12980 4984
rect 12876 4956 12884 4964
rect 12924 4956 12932 4964
rect 12380 4916 12388 4924
rect 12588 4918 12596 4926
rect 12492 4896 12500 4904
rect 11740 4656 11748 4664
rect 11564 4496 11572 4504
rect 11612 4476 11620 4484
rect 11660 4396 11668 4404
rect 11628 4376 11636 4384
rect 11676 4376 11684 4384
rect 11196 4316 11204 4324
rect 12300 4516 12308 4524
rect 12220 4496 12228 4504
rect 12284 4476 12292 4484
rect 12348 4336 12356 4344
rect 11708 4316 11716 4324
rect 11804 4316 11812 4324
rect 11836 4316 11844 4324
rect 11932 4294 11940 4302
rect 11020 4256 11028 4264
rect 11212 4276 11220 4284
rect 10492 4216 10500 4224
rect 10444 4176 10452 4184
rect 11020 4156 11028 4164
rect 11628 4156 11636 4164
rect 11788 4176 11796 4184
rect 12444 4316 12452 4324
rect 12492 4316 12500 4324
rect 12396 4296 12404 4304
rect 12396 4196 12404 4204
rect 12428 4196 12436 4204
rect 12972 4156 12980 4164
rect 11036 4136 11044 4144
rect 11068 4136 11076 4144
rect 11676 4136 11684 4144
rect 11708 4136 11716 4144
rect 12236 4136 12244 4144
rect 11004 4116 11012 4124
rect 11084 4116 11092 4124
rect 10924 4096 10932 4104
rect 11196 4096 11204 4104
rect 11148 4036 11156 4044
rect 11084 4016 11092 4024
rect 11612 3936 11620 3944
rect 10924 3916 10932 3924
rect 10956 3916 10964 3924
rect 11564 3916 11572 3924
rect 11596 3916 11604 3924
rect 11612 3916 11620 3924
rect 12300 4116 12308 4124
rect 12220 4096 12228 4104
rect 11724 4076 11732 4084
rect 12284 4076 12292 4084
rect 12300 3936 12308 3944
rect 11836 3916 11844 3924
rect 11020 3896 11028 3904
rect 11676 3896 11684 3904
rect 8540 3876 8548 3884
rect 8620 3736 8628 3744
rect 8524 3716 8532 3724
rect 7948 3696 7956 3704
rect 8588 3696 8596 3704
rect 7900 3676 7908 3684
rect 7724 3576 7732 3584
rect 9020 3556 9028 3564
rect 7292 3516 7300 3524
rect 7804 3516 7812 3524
rect 7900 3516 7908 3524
rect 7948 3516 7956 3524
rect 8524 3516 8532 3524
rect 8588 3516 8596 3524
rect 9068 3516 9076 3524
rect 7388 3494 7396 3502
rect 8380 3496 8388 3504
rect 8444 3496 8452 3504
rect 8476 3496 8484 3504
rect 9180 3816 9188 3824
rect 9180 3756 9188 3764
rect 9516 3736 9524 3744
rect 10412 3876 10420 3884
rect 10924 3876 10932 3884
rect 9996 3856 10004 3864
rect 10428 3796 10436 3804
rect 10492 3796 10500 3804
rect 11660 3816 11668 3824
rect 11628 3776 11636 3784
rect 9724 3716 9732 3724
rect 9612 3696 9620 3704
rect 9244 3516 9252 3524
rect 9132 3496 9140 3504
rect 9340 3494 9348 3502
rect 7724 3476 7732 3484
rect 7964 3476 7972 3484
rect 6540 3316 6548 3324
rect 7100 3316 7108 3324
rect 7020 3296 7028 3304
rect 7084 3276 7092 3284
rect 6572 3136 6580 3144
rect 7148 3136 7156 3144
rect 6620 3116 6628 3124
rect 6572 3096 6580 3104
rect 7068 3096 7076 3104
rect 6428 2956 6436 2964
rect 4524 2916 4532 2924
rect 4780 2918 4788 2926
rect 4412 2896 4420 2904
rect 4460 2896 4468 2904
rect 4684 2896 4692 2904
rect 5260 2896 5268 2904
rect 5340 2896 5348 2904
rect 5836 2896 5844 2904
rect 5292 2876 5300 2884
rect 5292 2836 5300 2844
rect 3980 2776 3988 2784
rect 5196 2756 5204 2764
rect 4412 2716 4420 2724
rect 4460 2716 4468 2724
rect 4588 2716 4596 2724
rect 4652 2716 4660 2724
rect 4684 2716 4692 2724
rect 5340 2716 5348 2724
rect 4524 2696 4532 2704
rect 4764 2694 4772 2702
rect 5436 2694 5444 2702
rect 3980 2616 3988 2624
rect 3980 2556 3988 2564
rect 3852 2516 3860 2524
rect 3772 2496 3780 2504
rect 3788 2496 3796 2504
rect 3804 2496 3812 2504
rect 3836 2496 3844 2504
rect 4412 2496 4420 2504
rect 4460 2496 4468 2504
rect 3292 2416 3300 2424
rect 3324 2336 3332 2344
rect 3772 2316 3780 2324
rect 3804 2316 3812 2324
rect 3340 2116 3348 2124
rect 3852 2116 3860 2124
rect 3772 2096 3780 2104
rect 3836 2096 3844 2104
rect 3292 1976 3300 1984
rect 3900 2076 3908 2084
rect 3324 1936 3332 1944
rect 3388 1916 3396 1924
rect 3324 1896 3332 1904
rect 3948 2416 3956 2424
rect 4412 2316 4420 2324
rect 3980 2156 3988 2164
rect 4636 2616 4644 2624
rect 4588 2596 4596 2604
rect 5772 2596 5780 2604
rect 5276 2576 5284 2584
rect 5244 2536 5252 2544
rect 5148 2516 5156 2524
rect 5068 2496 5076 2504
rect 5132 2496 5140 2504
rect 4588 2416 4596 2424
rect 5276 2396 5284 2404
rect 4700 2376 4708 2384
rect 5820 2516 5828 2524
rect 5804 2376 5812 2384
rect 5132 2336 5140 2344
rect 5276 2336 5284 2344
rect 5292 2336 5300 2344
rect 4700 2316 4708 2324
rect 5068 2316 5076 2324
rect 5260 2316 5268 2324
rect 5340 2316 5348 2324
rect 4684 2296 4692 2304
rect 4972 2294 4980 2302
rect 5180 2296 5188 2304
rect 5948 2896 5956 2904
rect 5996 2896 6004 2904
rect 5884 2856 5892 2864
rect 5900 2856 5908 2864
rect 6476 2836 6484 2844
rect 5932 2816 5940 2824
rect 6412 2756 6420 2764
rect 6364 2716 6372 2724
rect 5932 2616 5940 2624
rect 6540 3056 6548 3064
rect 6588 3016 6596 3024
rect 7388 3318 7396 3326
rect 7724 3316 7732 3324
rect 7836 3316 7844 3324
rect 7804 3296 7812 3304
rect 7900 3296 7908 3304
rect 7948 3296 7956 3304
rect 7804 3276 7812 3284
rect 8380 3276 8388 3284
rect 7900 3156 7908 3164
rect 7244 3136 7252 3144
rect 7292 3116 7300 3124
rect 7948 3116 7956 3124
rect 7180 3096 7188 3104
rect 8380 3096 8388 3104
rect 7964 3076 7972 3084
rect 8444 3076 8452 3084
rect 7724 2956 7732 2964
rect 7100 2916 7108 2924
rect 7212 2916 7220 2924
rect 7100 2896 7108 2904
rect 7196 2856 7204 2864
rect 7068 2796 7076 2804
rect 6572 2756 6580 2764
rect 7020 2716 7028 2724
rect 7100 2756 7108 2764
rect 6924 2694 6932 2702
rect 7708 2736 7716 2744
rect 7788 2736 7796 2744
rect 7660 2716 7668 2724
rect 7772 2696 7780 2704
rect 7836 3056 7844 3064
rect 9084 3476 9092 3484
rect 9676 3456 9684 3464
rect 9708 3436 9716 3444
rect 9132 3356 9140 3364
rect 8972 3296 8980 3304
rect 9004 3296 9012 3304
rect 8524 3136 8532 3144
rect 9036 3136 9044 3144
rect 8524 3116 8532 3124
rect 8588 3116 8596 3124
rect 8476 3096 8484 3104
rect 9116 3336 9124 3344
rect 9628 3336 9636 3344
rect 9980 3718 9988 3726
rect 9868 3696 9876 3704
rect 9884 3696 9892 3704
rect 10540 3696 10548 3704
rect 10332 3676 10340 3684
rect 10476 3676 10484 3684
rect 10988 3676 10996 3684
rect 9996 3656 10004 3664
rect 10988 3656 10996 3664
rect 10268 3516 10276 3524
rect 10332 3516 10340 3524
rect 10540 3516 10548 3524
rect 9996 3496 10004 3504
rect 10348 3496 10356 3504
rect 10428 3496 10436 3504
rect 11196 3696 11204 3704
rect 11148 3676 11156 3684
rect 11148 3516 11156 3524
rect 11196 3516 11204 3524
rect 10380 3456 10388 3464
rect 9788 3356 9796 3364
rect 9980 3336 9988 3344
rect 9708 3316 9716 3324
rect 9612 3296 9620 3304
rect 9660 3276 9668 3284
rect 9708 3256 9716 3264
rect 9196 3136 9204 3144
rect 9244 3116 9252 3124
rect 9884 3296 9892 3304
rect 9852 3276 9860 3284
rect 10332 3176 10340 3184
rect 10268 3116 10276 3124
rect 10380 3096 10388 3104
rect 9756 3076 9764 3084
rect 10284 3076 10292 3084
rect 10636 3476 10644 3484
rect 11084 3496 11092 3504
rect 10492 3396 10500 3404
rect 11628 3396 11636 3404
rect 11132 3356 11140 3364
rect 11052 3336 11060 3344
rect 11580 3336 11588 3344
rect 11852 3876 11860 3884
rect 12268 3876 12276 3884
rect 11740 3856 11748 3864
rect 12268 3816 12276 3824
rect 12364 4136 12372 4144
rect 12876 4136 12884 4144
rect 12972 4116 12980 4124
rect 12860 4096 12868 4104
rect 12908 4096 12916 4104
rect 12396 4056 12404 4064
rect 12908 3936 12916 3944
rect 12860 3916 12868 3924
rect 12972 3896 12980 3904
rect 12300 3716 12308 3724
rect 12764 3736 12772 3744
rect 12220 3696 12228 3704
rect 12284 3696 12292 3704
rect 12364 3696 12372 3704
rect 12300 3576 12308 3584
rect 12284 3556 12292 3564
rect 12220 3516 12228 3524
rect 12428 3576 12436 3584
rect 12380 3556 12388 3564
rect 11788 3396 11796 3404
rect 11740 3356 11748 3364
rect 10428 3296 10436 3304
rect 10924 3296 10932 3304
rect 10956 3296 10964 3304
rect 11036 3236 11044 3244
rect 10988 3156 10996 3164
rect 10476 3136 10484 3144
rect 10540 3116 10548 3124
rect 10428 3096 10436 3104
rect 11564 3296 11572 3304
rect 11596 3296 11604 3304
rect 11932 3318 11940 3326
rect 12268 3316 12276 3324
rect 11836 3296 11844 3304
rect 12348 3276 12356 3284
rect 11660 3196 11668 3204
rect 11644 3136 11652 3144
rect 11772 3136 11780 3144
rect 12348 3136 12356 3144
rect 11196 3116 11204 3124
rect 11836 3116 11844 3124
rect 10636 3094 10644 3102
rect 9068 3016 9076 3024
rect 8316 2896 8324 2904
rect 7868 2796 7876 2804
rect 7820 2756 7828 2764
rect 8364 2756 8372 2764
rect 8316 2716 8324 2724
rect 6268 2518 6276 2526
rect 6732 2518 6740 2526
rect 6364 2496 6372 2504
rect 6636 2496 6644 2504
rect 6460 2416 6468 2424
rect 5884 2336 5892 2344
rect 7084 2336 7092 2344
rect 5948 2316 5956 2324
rect 5996 2316 6004 2324
rect 6604 2316 6612 2324
rect 6636 2316 6644 2324
rect 5884 2296 5892 2304
rect 6540 2296 6548 2304
rect 7564 2676 7572 2684
rect 7228 2636 7236 2644
rect 8380 2556 8388 2564
rect 8684 2918 8692 2926
rect 8508 2896 8516 2904
rect 8588 2896 8596 2904
rect 9036 2796 9044 2804
rect 8524 2756 8532 2764
rect 9100 2756 9108 2764
rect 8972 2716 8980 2724
rect 9852 2996 9860 3004
rect 9788 2956 9796 2964
rect 11292 3094 11300 3102
rect 11692 3076 11700 3084
rect 11628 3016 11636 3024
rect 11292 2936 11300 2944
rect 11852 3076 11860 3084
rect 12316 2956 12324 2964
rect 9132 2916 9140 2924
rect 10316 2916 10324 2924
rect 10476 2916 10484 2924
rect 9196 2896 9204 2904
rect 9244 2896 9252 2904
rect 9884 2896 9892 2904
rect 10540 2896 10548 2904
rect 9756 2876 9764 2884
rect 9852 2876 9860 2884
rect 10988 2836 10996 2844
rect 9180 2796 9188 2804
rect 10332 2796 10340 2804
rect 9132 2756 9140 2764
rect 9820 2736 9828 2744
rect 9852 2736 9860 2744
rect 10476 2736 10484 2744
rect 9612 2716 9620 2724
rect 9660 2716 9668 2724
rect 9852 2716 9860 2724
rect 9868 2716 9876 2724
rect 9884 2716 9892 2724
rect 10540 2716 10548 2724
rect 9708 2696 9716 2704
rect 9980 2694 9988 2702
rect 10428 2696 10436 2704
rect 10636 2694 10644 2702
rect 9068 2616 9076 2624
rect 9708 2596 9716 2604
rect 9676 2576 9684 2584
rect 10364 2596 10372 2604
rect 7788 2536 7796 2544
rect 7820 2536 7828 2544
rect 8684 2536 8692 2544
rect 7564 2518 7572 2526
rect 7788 2516 7796 2524
rect 7836 2516 7844 2524
rect 8044 2518 8052 2526
rect 8172 2516 8180 2524
rect 7660 2496 7668 2504
rect 7948 2496 7956 2504
rect 7740 2456 7748 2464
rect 7900 2336 7908 2344
rect 7292 2316 7300 2324
rect 7948 2316 7956 2324
rect 8524 2496 8532 2504
rect 8588 2496 8596 2504
rect 8428 2436 8436 2444
rect 8380 2376 8388 2384
rect 8012 2294 8020 2302
rect 8172 2296 8180 2304
rect 9036 2376 9044 2384
rect 8588 2316 8596 2324
rect 8476 2296 8484 2304
rect 8508 2296 8516 2304
rect 8684 2294 8692 2302
rect 7132 2276 7140 2284
rect 7164 2276 7172 2284
rect 8380 2276 8388 2284
rect 8428 2276 8436 2284
rect 5772 2136 5780 2144
rect 4524 2116 4532 2124
rect 4412 2096 4420 2104
rect 4460 2076 4468 2084
rect 3932 1936 3940 1944
rect 3996 1916 4004 1924
rect 4044 1916 4052 1924
rect 2684 1856 2692 1864
rect 2620 1776 2628 1784
rect 2572 1716 2580 1724
rect 2460 1696 2468 1704
rect 2508 1676 2516 1684
rect 2540 1656 2548 1664
rect 2044 1536 2052 1544
rect 1980 1496 1988 1504
rect 2188 1494 2196 1502
rect 3196 1716 3204 1724
rect 3116 1696 3124 1704
rect 3228 1656 3236 1664
rect 3180 1556 3188 1564
rect 3228 1536 3236 1544
rect 2700 1516 2708 1524
rect 2748 1516 2756 1524
rect 2620 1496 2628 1504
rect 2828 1494 2836 1502
rect 1996 1396 2004 1404
rect 3212 1416 3220 1424
rect 2460 1296 2468 1304
rect 2508 1276 2516 1284
rect 2652 1296 2660 1304
rect 2748 1296 2756 1304
rect 2700 1276 2708 1284
rect 2044 1136 2052 1144
rect 2540 1136 2548 1144
rect 2700 1136 2708 1144
rect 1980 1116 1988 1124
rect 2092 1116 2100 1124
rect 2748 1116 2756 1124
rect 2188 1094 2196 1102
rect 2556 1096 2564 1104
rect 2636 1096 2644 1104
rect 2572 996 2580 1004
rect 2012 916 2020 924
rect 2556 916 2564 924
rect 2636 916 2644 924
rect 2092 896 2100 904
rect 2044 876 2052 884
rect 2748 896 2756 904
rect 2700 876 2708 884
rect 2556 836 2564 844
rect 4476 1896 4484 1904
rect 5148 2116 5156 2124
rect 5068 2096 5076 2104
rect 5340 2096 5348 2104
rect 5276 2076 5284 2084
rect 4604 1916 4612 1924
rect 5820 2016 5828 2024
rect 5788 1996 5796 2004
rect 5788 1976 5796 1984
rect 5276 1936 5284 1944
rect 4652 1916 4660 1924
rect 4684 1916 4692 1924
rect 5196 1916 5204 1924
rect 5228 1896 5236 1904
rect 5196 1876 5204 1884
rect 3932 1856 3940 1864
rect 4044 1856 4052 1864
rect 3980 1816 3988 1824
rect 5116 1856 5124 1864
rect 4780 1736 4788 1744
rect 6476 2116 6484 2124
rect 5884 2096 5892 2104
rect 6364 2096 6372 2104
rect 6412 2096 6420 2104
rect 6364 1916 6372 1924
rect 6412 1916 6420 1924
rect 6588 2176 6596 2184
rect 6540 2156 6548 2164
rect 7228 2156 7236 2164
rect 7180 2136 7188 2144
rect 7788 2136 7796 2144
rect 7820 2136 7828 2144
rect 9020 2256 9028 2264
rect 7084 2116 7092 2124
rect 7132 2116 7140 2124
rect 7564 2118 7572 2126
rect 7788 2116 7796 2124
rect 7020 2096 7028 2104
rect 7148 1936 7156 1944
rect 6604 1916 6612 1924
rect 6636 1916 6644 1924
rect 6572 1896 6580 1904
rect 6460 1816 6468 1824
rect 6428 1796 6436 1804
rect 5436 1736 5444 1744
rect 5772 1736 5780 1744
rect 3852 1716 3860 1724
rect 5276 1716 5284 1724
rect 3772 1696 3780 1704
rect 3788 1696 3796 1704
rect 3804 1696 3812 1704
rect 3836 1696 3844 1704
rect 3836 1556 3844 1564
rect 3324 1516 3332 1524
rect 3388 1516 3396 1524
rect 3484 1494 3492 1502
rect 3820 1496 3828 1504
rect 4412 1696 4420 1704
rect 4684 1696 4692 1704
rect 4460 1676 4468 1684
rect 4652 1676 4660 1684
rect 5340 1696 5348 1704
rect 5292 1656 5300 1664
rect 3932 1576 3940 1584
rect 5276 1536 5284 1544
rect 3996 1516 4004 1524
rect 4012 1516 4020 1524
rect 4044 1516 4052 1524
rect 4556 1516 4564 1524
rect 4684 1516 4692 1524
rect 4140 1494 4148 1502
rect 4780 1494 4788 1502
rect 3244 1416 3252 1424
rect 3244 1156 3252 1164
rect 3228 1096 3236 1104
rect 2540 756 2548 764
rect 2044 736 2052 744
rect 2700 736 2708 744
rect 2092 716 2100 724
rect 2748 716 2756 724
rect 1980 696 1988 704
rect 2188 694 2196 702
rect 2588 696 2596 704
rect 2636 696 2644 704
rect 3180 696 3188 704
rect 2572 616 2580 624
rect 2188 518 2196 526
rect 2620 516 2628 524
rect 2844 518 2852 526
rect 2060 496 2068 504
rect 2092 496 2100 504
rect 2684 496 2692 504
rect 2700 496 2708 504
rect 2716 496 2724 504
rect 2748 496 2756 504
rect 2028 476 2036 484
rect 2700 436 2708 444
rect 2460 316 2468 324
rect 2716 316 2724 324
rect 2748 316 2756 324
rect 2636 296 2644 304
rect 780 276 788 284
rect 1276 276 1284 284
rect 1308 276 1316 284
rect 1964 276 1972 284
rect 2476 276 2484 284
rect 2588 276 2596 284
rect 2620 276 2628 284
rect 60 256 68 264
rect 700 216 708 224
rect 684 196 692 204
rect 60 156 68 164
rect 1324 196 1332 204
rect 1388 156 1396 164
rect 1980 156 1988 164
rect 3228 136 3236 144
rect 5772 1476 5780 1484
rect 3932 1336 3940 1344
rect 4316 1318 4324 1326
rect 3772 1296 3780 1304
rect 3804 1296 3812 1304
rect 3820 1256 3828 1264
rect 3388 1116 3396 1124
rect 3276 1096 3284 1104
rect 3484 1094 3492 1102
rect 4412 1296 4420 1304
rect 4044 1116 4052 1124
rect 4140 1094 4148 1102
rect 3292 996 3300 1004
rect 3340 996 3348 1004
rect 3932 1056 3940 1064
rect 3980 1016 3988 1024
rect 4524 976 4532 984
rect 3932 956 3940 964
rect 4572 1416 4580 1424
rect 4636 1396 4644 1404
rect 5164 1396 5172 1404
rect 5964 1696 5972 1704
rect 5996 1696 6004 1704
rect 6364 1516 6372 1524
rect 6396 1516 6404 1524
rect 6412 1516 6420 1524
rect 6732 1718 6740 1726
rect 7068 1716 7076 1724
rect 6636 1696 6644 1704
rect 7148 1676 7156 1684
rect 6572 1636 6580 1644
rect 7020 1516 7028 1524
rect 7660 2096 7668 2104
rect 7788 2016 7796 2024
rect 7724 1976 7732 1984
rect 7388 1894 7396 1902
rect 7836 2116 7844 2124
rect 7948 2096 7956 2104
rect 8316 1916 8324 1924
rect 8364 1916 8372 1924
rect 8428 1896 8436 1904
rect 7804 1876 7812 1884
rect 8332 1876 8340 1884
rect 7788 1756 7796 1764
rect 8428 1856 8436 1864
rect 8044 1736 8052 1744
rect 7180 1716 7188 1724
rect 7292 1696 7300 1704
rect 7244 1676 7252 1684
rect 7212 1536 7220 1544
rect 7660 1516 7668 1524
rect 7708 1516 7716 1524
rect 7772 1496 7780 1504
rect 7884 1696 7892 1704
rect 7900 1696 7908 1704
rect 7916 1696 7924 1704
rect 7948 1696 7956 1704
rect 7836 1676 7844 1684
rect 7900 1636 7908 1644
rect 7868 1596 7876 1604
rect 8364 1596 8372 1604
rect 8316 1516 8324 1524
rect 8412 1556 8420 1564
rect 5900 1416 5908 1424
rect 5932 1416 5940 1424
rect 5836 1336 5844 1344
rect 5868 1336 5876 1344
rect 7068 1416 7076 1424
rect 5068 1296 5076 1304
rect 5132 1296 5140 1304
rect 5228 1256 5236 1264
rect 4620 1176 4628 1184
rect 5068 1116 5076 1124
rect 5148 1116 5156 1124
rect 4316 918 4324 926
rect 3772 896 3780 904
rect 3804 896 3812 904
rect 3836 836 3844 844
rect 3308 776 3316 784
rect 3388 716 3396 724
rect 3484 694 3492 702
rect 3820 516 3828 524
rect 3772 316 3780 324
rect 3340 296 3348 304
rect 3292 276 3300 284
rect 4412 896 4420 904
rect 4460 876 4468 884
rect 4524 916 4532 924
rect 4652 896 4660 904
rect 4684 896 4692 904
rect 4044 716 4052 724
rect 4140 694 4148 702
rect 4476 696 4484 704
rect 4556 736 4564 744
rect 4652 736 4660 744
rect 4684 716 4692 724
rect 4588 696 4596 704
rect 4524 576 4532 584
rect 3996 496 4004 504
rect 4044 496 4052 504
rect 4460 476 4468 484
rect 4460 456 4468 464
rect 3996 336 4004 344
rect 4524 336 4532 344
rect 3996 316 4004 324
rect 4012 316 4020 324
rect 4044 316 4052 324
rect 4140 294 4148 302
rect 3868 256 3876 264
rect 3884 196 3892 204
rect 4636 616 4644 624
rect 5116 616 5124 624
rect 5820 1316 5828 1324
rect 5916 1316 5924 1324
rect 6428 1316 6436 1324
rect 6572 1316 6580 1324
rect 5948 1296 5956 1304
rect 5996 1296 6004 1304
rect 6636 1296 6644 1304
rect 5820 1276 5828 1284
rect 6540 1276 6548 1284
rect 5804 1216 5812 1224
rect 5276 1176 5284 1184
rect 6524 1256 6532 1264
rect 6428 1216 6436 1224
rect 6572 1216 6580 1224
rect 7148 1176 7156 1184
rect 7084 1156 7092 1164
rect 5948 1136 5956 1144
rect 7020 1116 7028 1124
rect 5612 1094 5620 1102
rect 8524 2076 8532 2084
rect 8492 2056 8500 2064
rect 8972 1916 8980 1924
rect 9004 1916 9012 1924
rect 9036 1916 9044 1924
rect 9052 1896 9060 1904
rect 8540 1816 8548 1824
rect 9132 2516 9140 2524
rect 9196 2496 9204 2504
rect 9244 2496 9252 2504
rect 9244 2316 9252 2324
rect 9132 2296 9140 2304
rect 9340 2294 9348 2302
rect 9676 2296 9684 2304
rect 9676 2256 9684 2264
rect 10380 2536 10388 2544
rect 9980 2518 9988 2526
rect 9788 2476 9796 2484
rect 9884 2496 9892 2504
rect 10268 2316 10276 2324
rect 10332 2316 10340 2324
rect 10380 2296 10388 2304
rect 10492 2556 10500 2564
rect 11020 2556 11028 2564
rect 11084 2916 11092 2924
rect 11948 2918 11956 2926
rect 11100 2896 11108 2904
rect 11196 2896 11204 2904
rect 11772 2896 11780 2904
rect 11804 2896 11812 2904
rect 11820 2896 11828 2904
rect 11836 2896 11844 2904
rect 11612 2816 11620 2824
rect 11564 2716 11572 2724
rect 11660 2716 11668 2724
rect 11836 2716 11844 2724
rect 11948 2694 11956 2702
rect 11628 2596 11636 2604
rect 11036 2536 11044 2544
rect 11068 2536 11076 2544
rect 11004 2516 11012 2524
rect 11084 2516 11092 2524
rect 10924 2496 10932 2504
rect 11196 2496 11204 2504
rect 10428 2396 10436 2404
rect 10956 2356 10964 2364
rect 10924 2316 10932 2324
rect 11132 2356 11140 2364
rect 11612 2336 11620 2344
rect 11564 2316 11572 2324
rect 11020 2296 11028 2304
rect 11052 2296 11060 2304
rect 11676 2296 11684 2304
rect 11788 2616 11796 2624
rect 12268 2596 12276 2604
rect 12348 2556 12356 2564
rect 12972 3396 12980 3404
rect 12380 3316 12388 3324
rect 12492 3296 12500 3304
rect 12444 3276 12452 3284
rect 12924 3216 12932 3224
rect 12972 3216 12980 3224
rect 12444 3116 12452 3124
rect 12492 3116 12500 3124
rect 12426 3096 12434 3104
rect 12300 2516 12308 2524
rect 12380 2516 12388 2524
rect 12220 2496 12228 2504
rect 12492 2496 12500 2504
rect 12444 2476 12452 2484
rect 12316 2456 12324 2464
rect 12284 2416 12292 2424
rect 11772 2316 11780 2324
rect 11804 2316 11812 2324
rect 11820 2316 11828 2324
rect 11836 2316 11844 2324
rect 11948 2294 11956 2302
rect 10364 2196 10372 2204
rect 10316 2176 10324 2184
rect 10636 2136 10644 2144
rect 11676 2156 11684 2164
rect 11932 2136 11940 2144
rect 9164 2116 9172 2124
rect 10972 2116 10980 2124
rect 9244 2096 9252 2104
rect 9884 2096 9892 2104
rect 9196 1996 9204 2004
rect 10348 1956 10356 1964
rect 9196 1916 9204 1924
rect 9244 1916 9252 1924
rect 9852 1916 9860 1924
rect 9884 1916 9892 1924
rect 9132 1896 9140 1904
rect 9788 1896 9796 1904
rect 9052 1716 9060 1724
rect 8972 1696 8980 1704
rect 8988 1696 8996 1704
rect 9004 1696 9012 1704
rect 9036 1676 9044 1684
rect 8476 1656 8484 1664
rect 9036 1576 9044 1584
rect 9084 1556 9092 1564
rect 8668 1494 8676 1502
rect 8428 1416 8436 1424
rect 8412 1396 8420 1404
rect 7180 1316 7188 1324
rect 7388 1318 7396 1326
rect 7724 1316 7732 1324
rect 7292 1296 7300 1304
rect 7788 1296 7796 1304
rect 7228 1176 7236 1184
rect 7180 1156 7188 1164
rect 7660 1116 7668 1124
rect 7564 1094 7572 1102
rect 7788 1096 7796 1104
rect 7836 1316 7844 1324
rect 7900 1296 7908 1304
rect 7948 1296 7956 1304
rect 7884 1156 7892 1164
rect 8316 1116 8324 1124
rect 8428 1096 8436 1104
rect 5836 1076 5844 1084
rect 5868 1076 5876 1084
rect 6460 1016 6468 1024
rect 5836 936 5844 944
rect 5868 936 5876 944
rect 7196 976 7204 984
rect 9340 1736 9348 1744
rect 9212 1696 9220 1704
rect 9244 1696 9252 1704
rect 9196 1676 9204 1684
rect 9196 1636 9204 1644
rect 9180 1596 9188 1604
rect 9660 1596 9668 1604
rect 9612 1516 9620 1524
rect 9724 1776 9732 1784
rect 9724 1736 9732 1744
rect 9740 1556 9748 1564
rect 9708 1516 9716 1524
rect 10540 2096 10548 2104
rect 11036 2076 11044 2084
rect 10444 2036 10452 2044
rect 10956 1936 10964 1944
rect 10924 1916 10932 1924
rect 11004 1896 11012 1904
rect 11084 2116 11092 2124
rect 11196 2096 11204 2104
rect 11836 2096 11844 2104
rect 11148 2076 11156 2084
rect 11644 2076 11652 2084
rect 11772 2076 11780 2084
rect 11100 2056 11108 2064
rect 12316 2036 12324 2044
rect 11628 1996 11636 2004
rect 12268 1956 12276 1964
rect 11148 1936 11156 1944
rect 11196 1916 11204 1924
rect 11836 1916 11844 1924
rect 10492 1736 10500 1744
rect 11932 1894 11940 1902
rect 11132 1756 11140 1764
rect 11468 1736 11476 1744
rect 10332 1716 10340 1724
rect 10268 1696 10276 1704
rect 9820 1676 9828 1684
rect 10332 1636 10340 1644
rect 10380 1596 10388 1604
rect 10380 1556 10388 1564
rect 9884 1516 9892 1524
rect 9996 1494 10004 1502
rect 9052 1316 9060 1324
rect 8972 1296 8980 1304
rect 8524 1276 8532 1284
rect 8524 1256 8532 1264
rect 9100 1136 9108 1144
rect 8588 1116 8596 1124
rect 8476 1096 8484 1104
rect 8684 1094 8692 1102
rect 9020 1096 9028 1104
rect 7884 956 7892 964
rect 8220 936 8228 944
rect 8684 936 8692 944
rect 5804 916 5812 924
rect 6092 918 6100 926
rect 7084 916 7092 924
rect 7100 916 7108 924
rect 5740 896 5748 904
rect 5996 896 6004 904
rect 7020 896 7028 904
rect 7660 896 7668 904
rect 5948 876 5956 884
rect 5276 856 5284 864
rect 6428 816 6436 824
rect 7708 796 7716 804
rect 5292 756 5300 764
rect 7772 796 7780 804
rect 5212 716 5220 724
rect 5740 716 5748 724
rect 5804 716 5812 724
rect 6588 736 6596 744
rect 7244 736 7252 744
rect 5996 716 6004 724
rect 7020 716 7028 724
rect 7196 716 7204 724
rect 7292 716 7300 724
rect 5868 696 5876 704
rect 6044 694 6052 702
rect 6428 696 6436 704
rect 6540 696 6548 704
rect 5836 676 5844 684
rect 5868 676 5876 684
rect 9020 916 9028 924
rect 8316 896 8324 904
rect 7900 756 7908 764
rect 7132 596 7140 604
rect 6492 536 6500 544
rect 5148 516 5156 524
rect 6092 518 6100 526
rect 5068 496 5076 504
rect 5852 496 5860 504
rect 5996 496 6004 504
rect 5132 476 5140 484
rect 5276 476 5284 484
rect 4572 436 4580 444
rect 5276 436 5284 444
rect 4620 416 4628 424
rect 6620 496 6628 504
rect 6636 496 6644 504
rect 4572 316 4580 324
rect 5068 316 5076 324
rect 5964 316 5972 324
rect 5996 316 6004 324
rect 6604 316 6612 324
rect 6636 316 6644 324
rect 7132 316 7140 324
rect 5180 296 5188 304
rect 5820 296 5828 304
rect 5926 296 5934 304
rect 6572 296 6580 304
rect 4572 276 4580 284
rect 4636 216 4644 224
rect 4572 196 4580 204
rect 5980 276 5988 284
rect 6508 276 6516 284
rect 5276 236 5284 244
rect 6588 216 6596 224
rect 6540 176 6548 184
rect 5436 136 5444 144
rect 6524 156 6532 164
rect 7132 156 7140 164
rect 6092 136 6100 144
rect 7228 576 7236 584
rect 7564 536 7572 544
rect 8380 596 8388 604
rect 8508 896 8516 904
rect 8588 896 8596 904
rect 9100 876 9108 884
rect 9020 736 9028 744
rect 8428 556 8436 564
rect 9084 616 9092 624
rect 9164 1316 9172 1324
rect 9212 1296 9220 1304
rect 9244 1296 9252 1304
rect 9676 1196 9684 1204
rect 9724 1196 9732 1204
rect 9196 1136 9204 1144
rect 9244 1116 9252 1124
rect 9132 1096 9140 1104
rect 9132 916 9140 924
rect 9244 896 9252 904
rect 9196 876 9204 884
rect 9692 876 9700 884
rect 9740 776 9748 784
rect 9132 696 9140 704
rect 9676 636 9684 644
rect 8588 536 8596 544
rect 9116 536 9124 544
rect 7660 496 7668 504
rect 7772 476 7780 484
rect 7292 316 7300 324
rect 7788 316 7796 324
rect 7180 296 7188 304
rect 7388 294 7396 302
rect 7724 296 7732 304
rect 8220 518 8228 526
rect 8316 496 8324 504
rect 8348 496 8356 504
rect 8364 496 8368 504
rect 8368 496 8372 504
rect 8588 496 8596 504
rect 9084 496 9092 504
rect 8428 476 8436 484
rect 9020 456 9028 464
rect 8364 436 8372 444
rect 8364 376 8372 384
rect 7868 356 7876 364
rect 9068 416 9076 424
rect 9068 356 9076 364
rect 7900 316 7908 324
rect 7948 316 7956 324
rect 8524 316 8532 324
rect 8588 316 8596 324
rect 7836 296 7844 304
rect 8380 296 8388 304
rect 8444 296 8452 304
rect 8476 296 8484 304
rect 9020 216 9028 224
rect 9196 496 9204 504
rect 9244 496 9252 504
rect 9692 456 9700 464
rect 9148 356 9156 364
rect 9724 376 9732 384
rect 9244 316 9252 324
rect 9980 1336 9988 1344
rect 10924 1696 10932 1704
rect 10940 1696 10948 1704
rect 10956 1696 10964 1704
rect 10988 1696 10996 1704
rect 10476 1576 10484 1584
rect 10924 1516 10932 1524
rect 10940 1516 10948 1524
rect 10956 1516 10964 1524
rect 10988 1516 10996 1524
rect 11020 1716 11028 1724
rect 11932 1718 11940 1726
rect 11052 1696 11060 1704
rect 11564 1696 11572 1704
rect 11196 1516 11204 1524
rect 11084 1496 11092 1504
rect 11628 1496 11636 1504
rect 11036 1476 11044 1484
rect 11068 1476 11076 1484
rect 10636 1318 10644 1326
rect 10972 1316 10980 1324
rect 9852 1296 9860 1304
rect 9884 1296 9892 1304
rect 10332 1136 10340 1144
rect 10268 1116 10276 1124
rect 10332 1096 10340 1104
rect 10540 1296 10548 1304
rect 11036 1276 11044 1284
rect 10956 1176 10964 1184
rect 10924 1116 10932 1124
rect 11004 1156 11012 1164
rect 11084 1316 11092 1324
rect 11196 1296 11204 1304
rect 11148 1276 11156 1284
rect 11660 1216 11668 1224
rect 11660 1176 11668 1184
rect 11628 1156 11636 1164
rect 11164 1116 11172 1124
rect 11196 1116 11204 1124
rect 11084 1096 11092 1104
rect 9788 956 9796 964
rect 11036 1036 11044 1044
rect 10428 956 10436 964
rect 9884 896 9892 904
rect 10540 896 10548 904
rect 9852 876 9860 884
rect 10332 876 10340 884
rect 10476 876 10484 884
rect 10988 856 10996 864
rect 9772 736 9780 744
rect 10332 736 10340 744
rect 10268 716 10276 724
rect 10460 716 10468 724
rect 10540 716 10548 724
rect 10332 696 10340 704
rect 10428 696 10436 704
rect 11132 996 11140 1004
rect 11692 1616 11700 1624
rect 11804 1696 11812 1704
rect 11836 1696 11844 1704
rect 12284 1536 12292 1544
rect 12220 1516 12228 1524
rect 12284 1496 12292 1504
rect 11932 1318 11940 1326
rect 11676 956 11684 964
rect 11820 1296 11828 1304
rect 11836 1296 11844 1304
rect 11740 1276 11748 1284
rect 12284 1136 12292 1144
rect 12220 1116 12228 1124
rect 12284 1096 12292 1104
rect 11468 918 11476 926
rect 11932 918 11940 926
rect 11564 896 11572 904
rect 11692 796 11700 804
rect 11100 736 11108 744
rect 11196 716 11204 724
rect 11628 696 11636 704
rect 11692 696 11700 704
rect 11628 556 11636 564
rect 9980 518 9988 526
rect 9884 496 9892 504
rect 10380 496 10388 504
rect 10268 316 10276 324
rect 10172 294 10180 302
rect 9852 196 9860 204
rect 10476 496 10484 504
rect 10540 496 10548 504
rect 10444 376 10452 384
rect 10956 376 10964 384
rect 10924 316 10932 324
rect 11004 316 11012 324
rect 11020 296 11028 304
rect 11084 516 11092 524
rect 11580 516 11588 524
rect 11196 496 11204 504
rect 11132 376 11140 384
rect 11068 356 11076 364
rect 11612 336 11620 344
rect 11676 336 11684 344
rect 11564 316 11572 324
rect 11820 896 11828 904
rect 11836 896 11844 904
rect 12284 736 12292 744
rect 12220 716 12228 724
rect 12284 696 12292 704
rect 11708 676 11716 684
rect 12236 676 12244 684
rect 11804 656 11812 664
rect 11804 496 11812 504
rect 11836 496 11844 504
rect 12300 476 12308 484
rect 11804 316 11812 324
rect 11836 316 11844 324
rect 11676 256 11684 264
rect 11692 256 11700 264
rect 11852 256 11860 264
rect 11628 196 11636 204
rect 11788 216 11796 224
rect 10636 136 10644 144
rect 12380 576 12388 584
rect 76 116 84 124
rect 1276 116 1284 124
rect 1900 116 1908 124
rect 1980 116 1988 124
rect 2188 118 2196 126
rect 2844 118 2852 126
rect 4524 116 4532 124
rect 5148 116 5156 124
rect 5772 116 5780 124
rect 7212 116 7220 124
rect 7724 116 7732 124
rect 7836 116 7844 124
rect 8380 116 8388 124
rect 8524 116 8532 124
rect 9132 116 9140 124
rect 10396 116 10404 124
rect 10972 116 10980 124
rect 11084 116 11092 124
rect 140 96 148 104
rect 1164 96 1172 104
rect 1212 96 1220 104
rect 1820 96 1828 104
rect 1884 96 1892 104
rect 2092 96 2100 104
rect 2748 96 2756 104
rect 3388 96 3396 104
rect 4412 96 4420 104
rect 4460 96 4468 104
rect 5068 96 5076 104
rect 5340 96 5348 104
rect 5964 96 5972 104
rect 7020 96 7028 104
rect 7292 96 7300 104
rect 7948 96 7956 104
rect 8588 96 8596 104
rect 9196 96 9204 104
rect 9244 96 9252 104
rect 9756 96 9764 104
rect 9852 96 9860 104
rect 9884 96 9892 104
rect 10540 96 10548 104
rect 11196 96 11204 104
rect 12220 96 12228 104
rect 12284 96 12292 104
rect 12924 96 12932 104
rect 2540 76 2548 84
rect 2700 76 2708 84
rect 3196 76 3204 84
rect 3324 76 3332 84
rect 7084 76 7092 84
rect 7804 76 7812 84
rect 7900 76 7908 84
rect 11052 76 11060 84
rect 11148 76 11156 84
rect 1836 36 1844 44
rect 92 16 100 24
rect 140 16 148 24
rect 204 16 212 24
rect 780 16 788 24
rect 1756 16 1764 24
rect 1804 16 1812 24
rect 2748 16 2756 24
rect 5964 16 5972 24
rect 5996 16 6004 24
rect 7004 16 7012 24
rect 9212 16 9220 24
rect 9244 16 9252 24
<< metal3 >>
rect 3252 8977 3340 8983
rect 3188 8957 3292 8963
rect 6148 8957 7132 8963
rect 7780 8957 7820 8963
rect 8388 8957 8540 8963
rect 564 8937 732 8943
rect 1172 8937 1980 8943
rect 2516 8937 2684 8943
rect 5204 8937 6595 8943
rect 1284 8917 1292 8923
rect 1821 8918 2364 8923
rect 1821 8917 2371 8918
rect 1821 8904 1827 8917
rect 2580 8917 2620 8923
rect 3236 8917 3244 8923
rect 4484 8917 5276 8923
rect 6589 8923 6595 8937
rect 7716 8937 7884 8943
rect 6589 8917 6723 8923
rect 516 8897 524 8903
rect 1876 8897 1891 8903
rect 1885 8884 1891 8897
rect 2372 8897 2460 8903
rect 3028 8897 3116 8903
rect 3172 8897 3180 8903
rect 3780 8897 3788 8903
rect 4004 8897 4012 8903
rect 5332 8897 5340 8903
rect 6004 8897 6140 8903
rect 6717 8903 6723 8917
rect 8436 8917 8492 8923
rect 6717 8897 7660 8903
rect 8260 8897 8316 8903
rect 8372 8897 8380 8903
rect 8916 8897 8972 8903
rect 9060 8897 9132 8903
rect 9156 8897 9244 8903
rect 9892 8897 9900 8903
rect 1172 8877 1212 8883
rect 4004 8877 4092 8883
rect 4685 8883 4691 8896
rect 4644 8877 4691 8883
rect 5796 8877 5948 8883
rect 6452 8877 6572 8883
rect 6637 8883 6643 8896
rect 6637 8877 6748 8883
rect 9044 8877 9196 8883
rect 9204 8877 9292 8883
rect 9700 8877 9852 8883
rect 10541 8883 10547 8896
rect 10404 8877 10547 8883
rect 10996 8877 11148 8883
rect 1220 8857 3996 8863
rect 1396 8837 1420 8843
rect 1348 8817 1900 8823
rect 5764 8777 5932 8783
rect 7156 8777 7228 8783
rect 10340 8777 10476 8783
rect 564 8757 732 8763
rect 1188 8757 1340 8763
rect 1892 8757 2028 8763
rect 4580 8757 4956 8763
rect 5828 8757 5868 8763
rect 6420 8757 6572 8763
rect 7092 8757 7164 8763
rect 8052 8757 8492 8763
rect 9716 8757 9772 8763
rect 10404 8757 10428 8763
rect 10644 8757 11292 8763
rect 11300 8757 11676 8763
rect 1197 8737 1212 8743
rect 1197 8724 1203 8737
rect 3908 8737 3996 8743
rect 7284 8737 7708 8743
rect 7908 8737 8524 8743
rect 9300 8737 9820 8743
rect 10884 8737 10956 8743
rect 1172 8717 1180 8723
rect 1812 8717 1820 8723
rect 2724 8717 2732 8723
rect 3316 8717 3324 8723
rect 3453 8717 4044 8723
rect 628 8697 652 8703
rect 2580 8697 2668 8703
rect 2749 8703 2755 8716
rect 2676 8697 2755 8703
rect 3453 8703 3459 8717
rect 5140 8717 5148 8723
rect 5860 8717 6364 8723
rect 6916 8717 7020 8723
rect 7668 8717 7676 8723
rect 7700 8717 7708 8723
rect 7716 8717 7724 8723
rect 7892 8717 7900 8723
rect 7908 8717 7916 8723
rect 8868 8717 8972 8723
rect 10868 8717 10924 8723
rect 11188 8717 11196 8723
rect 11780 8717 11804 8723
rect 11812 8717 11820 8723
rect 3236 8697 3459 8703
rect 3828 8697 3932 8703
rect 6516 8697 6604 8703
rect 7412 8702 7571 8703
rect 7412 8697 7564 8702
rect 9076 8702 9523 8703
rect 9076 8697 9516 8702
rect 11837 8703 11843 8716
rect 11700 8697 11843 8703
rect 1188 8677 1324 8683
rect 4548 8677 4636 8683
rect 6612 8677 7036 8683
rect 11044 8677 11068 8683
rect 52 8657 140 8663
rect 1172 8657 1324 8663
rect 5844 8637 5852 8643
rect 1300 8617 1388 8623
rect 2676 8617 2684 8623
rect 6420 8617 6428 8623
rect 6452 8617 6460 8623
rect 10356 8617 10364 8623
rect 11956 8617 12316 8623
rect 52 8597 60 8603
rect 532 8597 636 8603
rect 2516 8597 2588 8603
rect 5252 8597 5260 8603
rect 8388 8597 8396 8603
rect 2468 8577 2524 8583
rect 8436 8577 8460 8583
rect 4500 8557 6540 8563
rect 7620 8557 7788 8563
rect 8388 8557 8540 8563
rect 11828 8557 12220 8563
rect 132 8537 652 8543
rect 3261 8537 3468 8543
rect 2196 8518 3020 8523
rect 2196 8517 3027 8518
rect 3261 8523 3267 8537
rect 3476 8537 6092 8543
rect 6100 8537 7132 8543
rect 7140 8537 7187 8543
rect 7181 8524 7187 8537
rect 7396 8537 7404 8543
rect 8420 8537 9139 8543
rect 9133 8524 9139 8537
rect 3236 8517 3267 8523
rect 3844 8517 4588 8523
rect 5924 8517 6028 8523
rect 9684 8517 9820 8523
rect 10628 8518 10636 8523
rect 10628 8517 10643 8518
rect 10980 8517 11084 8523
rect 1044 8497 1164 8503
rect 1716 8497 1820 8503
rect 2052 8497 2060 8503
rect 3380 8497 3388 8503
rect 4052 8497 4076 8503
rect 4964 8497 5068 8503
rect 5348 8497 5836 8503
rect 6708 8497 7020 8503
rect 7252 8497 7260 8503
rect 7268 8497 7276 8503
rect 7300 8497 7404 8503
rect 8372 8497 8380 8503
rect 8852 8497 8972 8503
rect 9188 8497 9196 8503
rect 9252 8497 9260 8503
rect 9892 8497 9900 8503
rect 10548 8497 10700 8503
rect 11172 8497 11196 8503
rect 11780 8497 11788 8503
rect 11796 8497 11804 8503
rect 11812 8497 11820 8503
rect 84 8477 636 8483
rect 692 8477 1116 8483
rect 1156 8477 1212 8483
rect 3149 8483 3155 8496
rect 5133 8484 5139 8496
rect 3149 8477 3164 8483
rect 3172 8477 3324 8483
rect 3844 8477 3996 8483
rect 5156 8477 5180 8483
rect 5204 8477 5276 8483
rect 5956 8477 6012 8483
rect 8317 8483 8323 8496
rect 7748 8477 8323 8483
rect 8964 8477 9036 8483
rect 11044 8477 11148 8483
rect 11837 8483 11843 8496
rect 11812 8477 11843 8483
rect 3188 8457 3324 8463
rect 8868 8457 9068 8463
rect 10884 8457 11004 8463
rect 2004 8437 4044 8443
rect 564 8417 3228 8423
rect 7268 8417 7868 8423
rect 8260 8417 9708 8423
rect 7140 8397 11196 8403
rect 564 8377 732 8383
rect 1268 8377 1276 8383
rect 3844 8377 3980 8383
rect 7076 8377 7228 8383
rect 7780 8377 7868 8383
rect 10996 8377 11004 8383
rect 11012 8377 11100 8383
rect 628 8357 668 8363
rect 1220 8357 1372 8363
rect 1892 8357 2028 8363
rect 2052 8357 2524 8363
rect 2532 8357 3164 8363
rect 3908 8357 3932 8363
rect 7716 8357 7820 8363
rect 10260 8357 10332 8363
rect 4420 8337 4460 8343
rect 4580 8337 5347 8343
rect 5341 8324 5347 8337
rect 5796 8337 5948 8343
rect 7092 8337 7244 8343
rect 9044 8337 9196 8343
rect 11044 8337 11148 8343
rect 532 8317 556 8323
rect 1108 8317 1164 8323
rect 1700 8317 1820 8323
rect 2388 8317 2460 8323
rect 2676 8317 2700 8323
rect 2708 8317 2732 8323
rect 2756 8317 2844 8323
rect 3780 8317 3836 8323
rect 4420 8317 4492 8323
rect 4692 8317 4716 8323
rect 5284 8317 5292 8323
rect 5988 8317 5996 8323
rect 6516 8317 6572 8323
rect 6596 8317 6604 8323
rect 6628 8317 6636 8323
rect 7796 8317 8220 8323
rect 8228 8317 8316 8323
rect 8340 8317 8348 8323
rect 8516 8317 8524 8323
rect 8564 8317 8588 8323
rect 9252 8317 9324 8323
rect 10116 8317 10268 8323
rect 10548 8317 10668 8323
rect 11204 8317 11292 8323
rect 11652 8317 11804 8323
rect 1940 8297 1964 8303
rect 2692 8297 2764 8303
rect 5124 8297 5132 8303
rect 6628 8302 6643 8303
rect 6628 8297 6636 8302
rect 8436 8297 8476 8303
rect 10404 8297 10428 8303
rect 11837 8303 11843 8316
rect 11700 8297 11843 8303
rect 1316 8277 1836 8283
rect 2596 8277 2620 8283
rect 3268 8277 3788 8283
rect 3924 8277 4428 8283
rect 7172 8277 7676 8283
rect 7748 8277 8220 8283
rect 8964 8257 9068 8263
rect 2628 8237 7948 8243
rect 9028 8237 9052 8243
rect 9060 8237 9996 8243
rect 8916 8217 9724 8223
rect 52 8197 1116 8203
rect 2516 8197 2524 8203
rect 5252 8197 5260 8203
rect 11636 8197 11644 8203
rect 12276 8197 12284 8203
rect 8436 8177 12220 8183
rect 6436 8157 6588 8163
rect 2180 8137 2684 8143
rect 5220 8137 5724 8143
rect 5764 8137 5932 8143
rect 8084 8137 10636 8143
rect 10644 8137 10652 8143
rect 84 8117 732 8123
rect 1876 8117 1980 8123
rect 2564 8118 3020 8123
rect 2564 8117 3027 8118
rect 3828 8117 3932 8123
rect 4484 8117 4620 8123
rect 6484 8117 6540 8123
rect 7396 8118 7612 8123
rect 7389 8117 7612 8118
rect 7620 8117 7660 8123
rect 7796 8117 7836 8123
rect 9172 8117 9324 8123
rect 9780 8117 12115 8123
rect 8589 8104 8595 8116
rect 1204 8097 1212 8103
rect 1332 8097 1436 8103
rect 2100 8097 2172 8103
rect 3028 8097 3116 8103
rect 3284 8097 3388 8103
rect 3908 8097 3996 8103
rect 4020 8097 4044 8103
rect 4692 8097 4748 8103
rect 6292 8097 6364 8103
rect 6420 8097 6428 8103
rect 6948 8097 7020 8103
rect 7284 8097 7292 8103
rect 7956 8097 7980 8103
rect 8692 8097 9196 8103
rect 10532 8097 10540 8103
rect 11028 8097 11148 8103
rect 11204 8097 11516 8103
rect 12109 8103 12115 8117
rect 12109 8097 12220 8103
rect 141 8083 147 8096
rect 52 8077 147 8083
rect 740 8077 1212 8083
rect 1956 8077 2044 8083
rect 3044 8077 3164 8083
rect 3172 8077 5388 8083
rect 7748 8077 7900 8083
rect 8532 8077 8652 8083
rect 10269 8083 10275 8096
rect 10269 8077 10284 8083
rect 10996 8077 11036 8083
rect 12212 8077 12284 8083
rect 3220 8057 5100 8063
rect 6436 8037 8844 8043
rect 8852 8037 10636 8043
rect 10884 8037 11020 8043
rect 2644 8017 2668 8023
rect 2852 8017 3324 8023
rect 7076 8017 7116 8023
rect 9684 8017 10332 8023
rect 708 7997 1260 8003
rect 1268 7997 1292 8003
rect 6756 7997 8428 8003
rect 10260 7997 10316 8003
rect 1268 7977 1372 7983
rect 2052 7977 2108 7983
rect 4484 7977 4604 7983
rect 8388 7977 10684 7983
rect 10692 7977 11292 7983
rect 1220 7957 1340 7963
rect 1700 7957 2204 7963
rect 2212 7957 2636 7963
rect 2660 7957 10380 7963
rect 3172 7937 3228 7943
rect 3236 7937 4028 7943
rect 5956 7937 6044 7943
rect 6612 7937 8268 7943
rect 8404 7937 9324 7943
rect 9748 7937 9852 7943
rect 10884 7937 10956 7943
rect 532 7917 540 7923
rect 1828 7917 1836 7923
rect 2020 7917 2092 7923
rect 2740 7917 3116 7923
rect 4004 7917 4044 7923
rect 4628 7917 4652 7923
rect 4660 7917 4668 7923
rect 5277 7923 5283 7936
rect 6605 7924 6611 7936
rect 12285 7924 12291 7936
rect 5277 7917 5292 7923
rect 6004 7917 6092 7923
rect 6644 7917 6748 7923
rect 7700 7917 7708 7923
rect 7716 7917 7724 7923
rect 7732 7917 7884 7923
rect 7956 7917 8076 7923
rect 8916 7917 8972 7923
rect 9220 7917 9228 7923
rect 9252 7917 9276 7923
rect 9892 7917 9996 7923
rect 11204 7917 11308 7923
rect 644 7897 1388 7903
rect 2189 7902 2204 7903
rect 2196 7897 2204 7902
rect 3828 7897 3836 7903
rect 4685 7903 4691 7916
rect 4548 7897 4691 7903
rect 5108 7897 5228 7903
rect 5460 7897 5884 7903
rect 6077 7897 6540 7903
rect 3028 7877 4060 7883
rect 4068 7877 4156 7883
rect 6077 7883 6083 7897
rect 6733 7902 7740 7903
rect 6740 7897 7740 7902
rect 7780 7897 7804 7903
rect 9332 7902 9347 7903
rect 9332 7897 9340 7902
rect 9748 7897 9788 7903
rect 11076 7897 11084 7903
rect 5412 7877 6083 7883
rect 6100 7877 7948 7883
rect 7956 7877 8060 7883
rect 10420 7877 10924 7883
rect 11044 7877 11068 7883
rect 11700 7877 12236 7883
rect 10292 7857 11020 7863
rect 7060 7837 7180 7843
rect 7812 7837 8428 7843
rect 10932 7837 11628 7843
rect 4420 7817 4476 7823
rect 4676 7817 5276 7823
rect 8404 7817 8412 7823
rect 9012 7817 9020 7823
rect 10868 7817 12268 7823
rect 84 7797 92 7803
rect 1108 7797 1260 7803
rect 4804 7797 5228 7803
rect 9620 7797 9676 7803
rect 9684 7797 9740 7803
rect 11636 7797 11644 7803
rect -51 7777 92 7783
rect -51 7737 -45 7777
rect 4148 7777 4636 7783
rect -35 7757 12 7763
rect -35 7723 -29 7757
rect 1892 7757 2028 7763
rect 2116 7757 2684 7763
rect 11748 7757 11772 7763
rect 1284 7737 2364 7743
rect 4564 7737 5084 7743
rect 6772 7737 9084 7743
rect 9348 7737 9980 7743
rect 10004 7737 10316 7743
rect 10324 7737 10636 7743
rect 10660 7737 11932 7743
rect 685 7724 691 7736
rect -51 7717 -29 7723
rect 6740 7718 6764 7723
rect 6733 7717 6764 7718
rect 7076 7717 7180 7723
rect 7796 7717 7836 7723
rect 7892 7717 8380 7723
rect 8388 7717 8524 7723
rect 1885 7704 1891 7716
rect 6397 7704 6403 7716
rect 468 7697 524 7703
rect 564 7697 572 7703
rect 740 7697 748 7703
rect 1764 7697 1820 7703
rect 2500 7697 2508 7703
rect 2516 7697 2524 7703
rect 3156 7697 3164 7703
rect 3668 7697 3772 7703
rect 3812 7697 3868 7703
rect 4004 7697 4012 7703
rect 4964 7697 5068 7703
rect 5124 7697 5139 7703
rect 797 7683 803 7696
rect 596 7677 803 7683
rect 3117 7683 3123 7696
rect 5133 7684 5139 7697
rect 5732 7697 5740 7703
rect 7156 7697 7244 7703
rect 7764 7697 7900 7703
rect 7956 7697 8092 7703
rect 8580 7697 8588 7703
rect 9252 7697 9260 7703
rect 9892 7697 10220 7703
rect 10404 7697 10476 7703
rect 10548 7697 10684 7703
rect 11620 7697 11660 7703
rect 11748 7697 11836 7703
rect 3117 7677 3324 7683
rect 4004 7677 4524 7683
rect 6548 7677 6700 7683
rect 7700 7677 9196 7683
rect 9204 7677 9852 7683
rect 2084 7657 3852 7663
rect 3860 7657 5148 7663
rect 5172 7657 7292 7663
rect 11044 7657 11164 7663
rect 2004 7637 3164 7643
rect 5156 7637 7516 7643
rect 8388 7637 8508 7643
rect 2484 7617 5884 7623
rect 2036 7597 3212 7603
rect 6916 7597 9724 7603
rect 1236 7577 2508 7583
rect 3188 7577 4012 7583
rect 4484 7577 4604 7583
rect 4660 7577 5180 7583
rect 6468 7577 8428 7583
rect 2004 7557 2012 7563
rect 3844 7557 4684 7563
rect 7092 7557 7180 7563
rect 7204 7557 7228 7563
rect 7972 7557 8492 7563
rect 1380 7537 1932 7543
rect 1988 7537 2396 7543
rect 3060 7537 4780 7543
rect 4804 7537 5276 7543
rect 5956 7537 6060 7543
rect 9972 7537 10476 7543
rect 11652 7537 11772 7543
rect 804 7517 812 7523
rect 2756 7517 3228 7523
rect 3332 7517 3340 7523
rect 3396 7517 3532 7523
rect 3940 7517 3996 7523
rect 4004 7517 4012 7523
rect 4628 7517 4652 7523
rect 4660 7517 4668 7523
rect 6004 7517 6460 7523
rect 7028 7517 7036 7523
rect 7940 7517 7948 7523
rect 8836 7517 8972 7523
rect 9252 7517 9340 7523
rect 10548 7517 10716 7523
rect 11108 7517 11116 7523
rect 11780 7517 11836 7523
rect 84 7497 92 7503
rect 141 7503 147 7516
rect 7917 7504 7923 7516
rect 116 7497 147 7503
rect 1908 7502 2371 7503
rect 1908 7497 2364 7502
rect 2580 7497 2588 7503
rect 3124 7497 3164 7503
rect 3172 7497 3276 7503
rect 5396 7502 5619 7503
rect 5396 7497 5612 7502
rect 6084 7502 6099 7503
rect 6084 7497 6092 7502
rect 7140 7497 7148 7503
rect 8045 7502 8540 7503
rect 8052 7497 8540 7502
rect 9341 7502 9356 7503
rect 9348 7497 9356 7502
rect 9684 7497 9724 7503
rect 9748 7497 9964 7503
rect 10420 7497 10428 7503
rect 132 7477 652 7483
rect 1556 7477 2028 7483
rect 2596 7477 2620 7483
rect 3492 7477 3820 7483
rect 3828 7477 3996 7483
rect 5844 7477 5868 7483
rect 8388 7477 8684 7483
rect 8708 7477 9260 7483
rect 36 7457 11180 7463
rect 1156 7437 2028 7443
rect 4052 7437 4524 7443
rect 7044 7417 7068 7423
rect 9028 7417 9228 7423
rect 12212 7417 12268 7423
rect 740 7397 748 7403
rect 2468 7397 2684 7403
rect 6420 7397 6428 7403
rect 6948 7397 7228 7403
rect 8548 7397 9356 7403
rect 10356 7397 10364 7403
rect 11140 7397 11148 7403
rect 1300 7377 1388 7383
rect 9092 7377 9212 7383
rect 9220 7377 9244 7383
rect 1236 7357 1340 7363
rect 5348 7357 6060 7363
rect 9780 7357 10492 7363
rect 10500 7357 10531 7363
rect 1348 7337 1436 7343
rect 7796 7337 7820 7343
rect 8452 7337 8684 7343
rect 10525 7343 10531 7357
rect 10525 7337 11468 7343
rect 1284 7317 1292 7323
rect 1908 7317 2556 7323
rect 2580 7317 2604 7323
rect 3492 7318 3500 7323
rect 3485 7317 3500 7318
rect 3828 7317 3932 7323
rect 5156 7317 5212 7323
rect 5220 7317 6076 7323
rect 6740 7318 6764 7323
rect 6733 7317 6764 7318
rect 9172 7317 9228 7323
rect 9236 7317 9324 7323
rect 11924 7318 11932 7323
rect 11924 7317 11939 7318
rect 452 7297 524 7303
rect 1220 7297 1228 7303
rect 1668 7297 1820 7303
rect 2468 7297 2476 7303
rect 3156 7297 3164 7303
rect 3220 7297 3388 7303
rect 4004 7297 4044 7303
rect 4228 7297 5068 7303
rect 5732 7297 5756 7303
rect 5764 7297 5804 7303
rect 6276 7297 6364 7303
rect 6644 7297 6652 7303
rect 7524 7297 7660 7303
rect 7924 7297 7948 7303
rect 9252 7297 9372 7303
rect 10132 7297 10268 7303
rect 10340 7297 10348 7303
rect 10548 7297 10556 7303
rect 11572 7297 11740 7303
rect 11780 7297 11788 7303
rect 11796 7297 11804 7303
rect 11812 7297 11820 7303
rect 11844 7297 11852 7303
rect 708 7277 812 7283
rect 1892 7277 3036 7283
rect 3892 7277 3996 7283
rect 5140 7277 5276 7283
rect 10356 7277 10476 7283
rect 4100 7257 4620 7263
rect 7828 7257 8556 7263
rect 9684 7257 11612 7263
rect 10916 7237 11020 7243
rect 3988 7197 3996 7203
rect 7892 7197 8028 7203
rect 8036 7197 8412 7203
rect 1956 7177 2028 7183
rect 5124 7177 5932 7183
rect 7844 7177 7900 7183
rect 1220 7157 1372 7163
rect 1892 7157 1964 7163
rect 5204 7157 5836 7163
rect 7748 7157 9372 7163
rect 84 7137 172 7143
rect 3652 7137 3779 7143
rect 3773 7124 3779 7137
rect 6580 7137 7692 7143
rect 9108 7137 9196 7143
rect 9700 7137 9852 7143
rect 10324 7137 10332 7143
rect 10996 7137 11148 7143
rect 11652 7137 11772 7143
rect 84 7117 140 7123
rect 1076 7117 1164 7123
rect 1396 7117 1820 7123
rect 1844 7117 2124 7123
rect 2132 7117 2460 7123
rect 3220 7117 3644 7123
rect 3876 7117 3891 7123
rect 3117 7103 3123 7116
rect 3117 7097 3340 7103
rect 3885 7064 3891 7117
rect 5076 7117 5084 7123
rect 5252 7117 5340 7123
rect 5796 7117 6364 7123
rect 6420 7117 6508 7123
rect 6516 7117 6572 7123
rect 6996 7117 7020 7123
rect 7092 7117 7100 7123
rect 8324 7117 8332 7123
rect 8596 7117 8732 7123
rect 9252 7117 9356 7123
rect 9812 7117 9884 7123
rect 10404 7117 10476 7123
rect 10548 7117 10636 7123
rect 11124 7117 11196 7123
rect 11684 7117 11836 7123
rect 6484 7097 6588 7103
rect 6596 7097 6604 7103
rect 7124 7097 7132 7103
rect 7389 7102 7756 7103
rect 7396 7097 7756 7102
rect 7764 7102 8227 7103
rect 7764 7097 8220 7102
rect 8436 7097 8444 7103
rect 9028 7097 9132 7103
rect 10324 7097 10428 7103
rect 10980 7097 11564 7103
rect 3940 7077 4076 7083
rect 11748 7057 11788 7063
rect 5780 7037 5788 7043
rect 708 7017 716 7023
rect 2212 7017 2684 7023
rect 3396 7017 5868 7023
rect 6484 7017 12220 7023
rect 2148 6997 2620 7003
rect 5092 6997 7788 7003
rect 9396 6997 11708 7003
rect 12276 6997 12300 7003
rect 5188 6977 7980 6983
rect 1332 6937 1955 6943
rect 1876 6917 1900 6923
rect 1949 6923 1955 6937
rect 6740 6937 8668 6943
rect 8676 6937 8684 6943
rect 9348 6937 9356 6943
rect 1949 6917 1980 6923
rect 2196 6918 2204 6923
rect 2189 6917 2204 6918
rect 2596 6917 2636 6923
rect 3828 6917 4620 6923
rect 5364 6918 5436 6923
rect 5364 6917 5443 6918
rect 5844 6917 5884 6923
rect 7076 6917 7180 6923
rect 8436 6917 8508 6923
rect 8756 6917 9020 6923
rect 9028 6917 9132 6923
rect 532 6897 540 6903
rect 1156 6897 1164 6903
rect 1716 6897 1820 6903
rect 2100 6897 2204 6903
rect 4340 6897 4412 6903
rect 4692 6897 4828 6903
rect 5348 6897 5452 6903
rect 5844 6897 5996 6903
rect 6644 6897 6668 6903
rect 7300 6897 7388 6903
rect 8596 6897 8604 6903
rect 9108 6897 9196 6903
rect 9252 6897 9372 6903
rect 9892 6897 9939 6903
rect 1220 6877 1612 6883
rect 1748 6877 1884 6883
rect 1924 6877 2044 6883
rect 2052 6877 2140 6883
rect 2548 6877 2700 6883
rect 3204 6877 3324 6883
rect 4372 6877 4460 6883
rect 5284 6877 5404 6883
rect 7156 6877 7244 6883
rect 8372 6877 9100 6883
rect 9748 6877 9836 6883
rect 9933 6883 9939 6897
rect 10148 6897 10540 6903
rect 12164 6897 12220 6903
rect 9933 6877 10748 6883
rect 10996 6857 11148 6863
rect 6612 6837 7372 6843
rect 452 6817 620 6823
rect 9716 6817 10268 6823
rect 11796 6817 11916 6823
rect 2212 6797 2572 6803
rect 7396 6797 7724 6803
rect 8324 6797 8380 6803
rect 12276 6797 12924 6803
rect 4372 6777 4476 6783
rect 4484 6777 4652 6783
rect 6468 6777 6572 6783
rect 612 6757 636 6763
rect 3188 6757 4044 6763
rect 4516 6757 4780 6763
rect 6420 6757 6540 6763
rect 11524 6757 11628 6763
rect 11636 6757 11660 6763
rect 1956 6737 2044 6743
rect 9108 6737 9196 6743
rect 12308 6737 12444 6743
rect 68 6717 76 6723
rect 148 6717 380 6723
rect 1172 6717 1180 6723
rect 2052 6717 2092 6723
rect 2756 6717 2844 6723
rect 3876 6717 3996 6723
rect 4340 6717 4364 6723
rect 4692 6717 4732 6723
rect 5348 6717 5500 6723
rect 6308 6717 6364 6723
rect 7012 6717 7020 6723
rect 7300 6717 7388 6723
rect 7956 6717 8060 6723
rect 8516 6717 8531 6723
rect 8596 6717 8700 6723
rect 9252 6717 9356 6723
rect 10404 6717 10476 6723
rect 10756 6717 11196 6723
rect 12340 6717 12396 6723
rect 12484 6717 12492 6723
rect 1876 6697 1980 6703
rect 2836 6697 3276 6703
rect 3828 6697 3932 6703
rect 4628 6697 4668 6703
rect 5277 6703 5283 6716
rect 5124 6697 5283 6703
rect 8468 6697 8476 6703
rect 9028 6697 9132 6703
rect 9828 6697 9836 6703
rect 10180 6697 10316 6703
rect 10324 6697 10428 6703
rect 10644 6702 12131 6703
rect 10644 6697 12124 6702
rect 2829 6663 2835 6696
rect 2852 6677 3660 6683
rect 3668 6677 5420 6683
rect 5428 6677 6924 6683
rect 9748 6677 10364 6683
rect 10372 6677 11036 6683
rect 2829 6657 2844 6663
rect 1780 6617 4524 6623
rect 10020 6617 12316 6623
rect 740 6597 748 6603
rect 2036 6597 2044 6603
rect 4372 6597 8460 6603
rect 11652 6597 11660 6603
rect 1300 6577 1388 6583
rect 1252 6557 1340 6563
rect 7780 6557 7884 6563
rect 9060 6557 9132 6563
rect 9188 6557 11468 6563
rect 1972 6537 2476 6543
rect 2596 6537 2620 6543
rect 6436 6537 6588 6543
rect 7172 6537 7676 6543
rect 7716 6537 7836 6543
rect 8676 6537 9340 6543
rect 9348 6537 9516 6543
rect 10964 6537 11132 6543
rect 164 6518 236 6523
rect 164 6517 243 6518
rect 1284 6517 1292 6523
rect 1876 6517 1900 6523
rect 3828 6517 3932 6523
rect 5156 6517 5260 6523
rect 5428 6518 5436 6523
rect 5428 6517 5443 6518
rect 5780 6517 5884 6523
rect 6708 6518 6732 6523
rect 6708 6517 6739 6518
rect 9060 6517 9180 6523
rect 9732 6517 9740 6523
rect 10340 6517 10348 6523
rect 11028 6517 11068 6523
rect 11076 6517 11196 6523
rect 100 6497 140 6503
rect 1172 6497 1180 6503
rect 1220 6497 1244 6503
rect 1812 6497 1820 6503
rect 2420 6497 2460 6503
rect 2500 6497 2508 6503
rect 2516 6497 2524 6503
rect 3396 6497 3420 6503
rect 4580 6497 5068 6503
rect 6004 6497 6108 6503
rect 6484 6497 6620 6503
rect 6644 6497 6780 6503
rect 7085 6497 7660 6503
rect 7085 6484 7091 6497
rect 8324 6497 8348 6503
rect 8436 6497 8828 6503
rect 8868 6497 8972 6503
rect 9012 6497 9052 6503
rect 9540 6497 9612 6503
rect 10164 6497 10268 6503
rect 10324 6497 10339 6503
rect 10333 6484 10339 6497
rect 11476 6497 11564 6503
rect 11620 6497 11644 6503
rect 11828 6497 11836 6503
rect 1748 6477 1884 6483
rect 1940 6477 2364 6483
rect 2372 6477 2700 6483
rect 3252 6477 3324 6483
rect 3908 6477 3996 6483
rect 5028 6477 5132 6483
rect 5860 6477 5948 6483
rect 6052 6477 6572 6483
rect 6580 6477 6700 6483
rect 9828 6477 9852 6483
rect 11732 6477 11804 6483
rect 3300 6457 4044 6463
rect 532 6437 684 6443
rect 2388 6437 7820 6443
rect 1188 6417 1372 6423
rect 52 6397 156 6403
rect 612 6397 620 6403
rect 1924 6397 2188 6403
rect 2196 6397 2556 6403
rect 2564 6397 3244 6403
rect 3252 6397 4940 6403
rect 6420 6397 6428 6403
rect 7028 6397 7180 6403
rect 564 6377 732 6383
rect 6429 6364 6435 6376
rect 628 6357 668 6363
rect 5028 6357 5276 6363
rect 6484 6357 7004 6363
rect 7012 6357 8060 6363
rect 8324 6357 8524 6363
rect 1140 6337 1212 6343
rect 2052 6337 3132 6343
rect 4004 6337 4524 6343
rect 5028 6337 5132 6343
rect 5796 6337 5948 6343
rect 7252 6337 7356 6343
rect 8372 6337 8476 6343
rect 8973 6337 9532 6343
rect 756 6317 1164 6323
rect 1828 6317 2012 6323
rect 2020 6317 2076 6323
rect 2100 6317 2124 6323
rect 2756 6317 3164 6323
rect 3684 6317 3772 6323
rect 1284 6297 1292 6303
rect 2196 6277 3004 6283
rect 3869 6243 3875 6296
rect 3885 6264 3891 6336
rect 8973 6324 8979 6337
rect 9700 6337 9852 6343
rect 10340 6337 10476 6343
rect 10996 6337 11148 6343
rect 4004 6317 4012 6323
rect 4788 6317 4956 6323
rect 4964 6317 5068 6323
rect 5284 6317 5292 6323
rect 5348 6317 5468 6323
rect 6004 6317 6012 6323
rect 7076 6317 7084 6323
rect 7300 6317 7580 6323
rect 7828 6317 8300 6323
rect 9252 6317 9820 6323
rect 9876 6317 9884 6323
rect 10468 6317 10540 6323
rect 11204 6317 11212 6323
rect 11924 6317 12220 6323
rect 12292 6317 12300 6323
rect 7380 6302 7395 6303
rect 7380 6297 7388 6302
rect 8436 6297 8556 6303
rect 9341 6302 9356 6303
rect 9348 6297 9356 6302
rect 9364 6297 9724 6303
rect 3869 6237 3891 6243
rect 2068 6217 2572 6223
rect 2580 6217 3148 6223
rect 3812 6217 3868 6223
rect 52 6197 380 6203
rect 3124 6197 3180 6203
rect 3885 6203 3891 6237
rect 5076 6217 5164 6223
rect 5252 6217 5260 6223
rect 5316 6217 6588 6223
rect 7076 6217 7116 6223
rect 11860 6217 12316 6223
rect 3828 6197 3891 6203
rect 6308 6197 7228 6203
rect 8372 6197 9180 6203
rect 1940 6177 2028 6183
rect 2500 6177 2684 6183
rect 7076 6177 7100 6183
rect 8436 6177 9084 6183
rect 9732 6177 9836 6183
rect 100 6157 732 6163
rect 1892 6157 1964 6163
rect 2612 6157 2620 6163
rect 5764 6157 5932 6163
rect 5956 6157 6476 6163
rect 7156 6157 7276 6163
rect 9028 6157 9276 6163
rect 564 6137 684 6143
rect 1332 6137 1900 6143
rect 1908 6137 2556 6143
rect 6772 6137 7564 6143
rect 2564 6117 2636 6123
rect 2980 6118 3020 6123
rect 2980 6117 3027 6118
rect 3268 6117 3372 6123
rect 6580 6118 6732 6123
rect 6580 6117 6739 6118
rect 7652 6117 7667 6123
rect 1885 6104 1891 6116
rect 4013 6104 4019 6116
rect 7661 6104 7667 6117
rect 7780 6117 7788 6123
rect 10356 6117 10380 6123
rect 10980 6117 11084 6123
rect 11700 6117 11843 6123
rect 8589 6104 8595 6116
rect 11837 6104 11843 6117
rect 436 6097 524 6103
rect 1092 6097 1164 6103
rect 2372 6097 2460 6103
rect 3156 6097 3164 6103
rect 4052 6097 4124 6103
rect 4532 6097 4684 6103
rect 6516 6097 6636 6103
rect 6644 6097 6684 6103
rect 8260 6097 8316 6103
rect 9796 6097 10268 6103
rect 10276 6097 10508 6103
rect 10532 6097 10540 6103
rect 11188 6097 11196 6103
rect 980 6077 1340 6083
rect 1821 6083 1827 6096
rect 1412 6077 1827 6083
rect 2516 6077 2572 6083
rect 4564 6077 4652 6083
rect 6068 6077 8524 6083
rect 11044 6077 11148 6083
rect 100 6057 204 6063
rect 2596 6057 3836 6063
rect 3860 6057 3884 6063
rect 4644 6057 4732 6063
rect 7812 6057 7868 6063
rect 9684 6057 11180 6063
rect 2196 6037 2508 6043
rect 2516 6037 2972 6043
rect 52 6017 172 6023
rect 8420 6017 9900 6023
rect 2884 5957 3324 5963
rect 10372 5957 11804 5963
rect 500 5937 556 5943
rect 3892 5937 3996 5943
rect 5796 5937 5948 5943
rect 6452 5937 7244 5943
rect 7748 5937 7827 5943
rect 452 5917 524 5923
rect 804 5917 972 5923
rect 1700 5917 1820 5923
rect 2052 5917 2060 5923
rect 2100 5917 2108 5923
rect 2724 5917 2732 5923
rect 2756 5917 2876 5923
rect 3780 5917 3836 5923
rect 3860 5917 3884 5923
rect 3956 5917 4044 5923
rect 5060 5917 5068 5923
rect 5092 5917 5132 5923
rect 5284 5917 5308 5923
rect 6004 5917 6492 5923
rect 6644 5917 6796 5923
rect 7300 5917 7452 5923
rect 7821 5923 7827 5937
rect 10996 5937 11203 5943
rect 11197 5924 11203 5937
rect 11652 5937 11772 5943
rect 7821 5917 7900 5923
rect 9892 5917 9900 5923
rect 9908 5917 10156 5923
rect 10164 5917 10380 5923
rect 10404 5917 10524 5923
rect 10548 5917 10668 5923
rect 11140 5917 11148 5923
rect 11700 5917 11836 5923
rect 1332 5897 1676 5903
rect 1716 5902 1731 5903
rect 1716 5897 1724 5902
rect 3284 5897 3420 5903
rect 5188 5897 5196 5903
rect 5437 5902 5948 5903
rect 5444 5897 5948 5902
rect 6468 5897 7180 5903
rect 7796 5897 7836 5903
rect 7949 5903 7955 5916
rect 7908 5897 7955 5903
rect 8324 5902 8867 5903
rect 9341 5902 9708 5903
rect 8324 5897 8860 5902
rect 9348 5897 9708 5902
rect 9732 5897 9788 5903
rect 11261 5902 11267 5903
rect 11261 5884 11267 5894
rect 644 5877 668 5883
rect 9364 5877 10556 5883
rect 1140 5837 1324 5843
rect 5828 5837 6092 5843
rect 6100 5837 6908 5843
rect 708 5817 748 5823
rect 1300 5817 1388 5823
rect 6596 5817 6604 5823
rect 8388 5817 12220 5823
rect 4484 5797 4492 5803
rect 12276 5797 12284 5803
rect 12308 5797 12316 5803
rect 3956 5777 5324 5783
rect 10356 5777 10380 5783
rect 2468 5757 2684 5763
rect 4420 5757 4636 5763
rect 5156 5757 5276 5763
rect 7108 5757 7180 5763
rect 10324 5757 10348 5763
rect 5133 5737 5228 5743
rect 1284 5717 1964 5723
rect 2580 5717 2604 5723
rect 3012 5718 3020 5723
rect 5133 5724 5139 5737
rect 5844 5737 5868 5743
rect 7124 5737 7564 5743
rect 7796 5737 7820 5743
rect 8564 5737 8684 5743
rect 10324 5737 10364 5743
rect 3012 5717 3027 5718
rect 8029 5704 8035 5718
rect 9332 5718 9340 5723
rect 10644 5718 10652 5723
rect 9332 5717 9347 5718
rect 10637 5717 10652 5718
rect 10980 5717 11084 5723
rect 12285 5704 12291 5716
rect 68 5697 524 5703
rect 1108 5697 1164 5703
rect 1828 5697 1836 5703
rect 1908 5697 2188 5703
rect 3028 5697 3116 5703
rect 3140 5697 3148 5703
rect 4500 5697 5068 5703
rect 5476 5697 5484 5703
rect 5492 5697 5740 5703
rect 6964 5697 7020 5703
rect 7092 5697 7100 5703
rect 7700 5697 7708 5703
rect 7716 5697 7724 5703
rect 8596 5697 8604 5703
rect 9892 5697 9900 5703
rect 10452 5697 10540 5703
rect 10548 5697 10748 5703
rect 11037 5697 11196 5703
rect 3844 5677 4092 5683
rect 4100 5677 4796 5683
rect 4804 5677 5948 5683
rect 5956 5677 6060 5683
rect 7044 5677 7900 5683
rect 7908 5677 8012 5683
rect 8452 5677 8524 5683
rect 9748 5677 9852 5683
rect 11037 5683 11043 5697
rect 10996 5677 11043 5683
rect 11060 5677 11148 5683
rect 468 5657 3948 5663
rect 4420 5657 4460 5663
rect 500 5637 1324 5643
rect 3956 5637 7084 5643
rect 7092 5637 7708 5643
rect 612 5617 1372 5623
rect 564 5597 732 5603
rect 1092 5597 2028 5603
rect 2692 5597 2764 5603
rect 4468 5597 4652 5603
rect 5140 5597 5164 5603
rect -51 5577 76 5583
rect -51 5537 -45 5577
rect 4564 5577 5180 5583
rect 9092 5577 10924 5583
rect -35 5557 12 5563
rect -35 5523 -29 5557
rect 2644 5557 2732 5563
rect 4436 5557 4652 5563
rect 7092 5557 7228 5563
rect 7764 5557 7836 5563
rect 10356 5557 10380 5563
rect 10404 5557 12972 5563
rect 740 5537 1212 5543
rect 1892 5537 2876 5543
rect 3060 5537 3164 5543
rect 3172 5537 3500 5543
rect 4660 5537 5276 5543
rect 5300 5537 5852 5543
rect 6708 5537 7900 5543
rect 7908 5537 8012 5543
rect 10516 5537 11571 5543
rect 11565 5524 11571 5537
rect 11748 5537 11756 5543
rect 12292 5537 12444 5543
rect -51 5517 -29 5523
rect 1140 5517 1164 5523
rect 1716 5517 1820 5523
rect 2356 5517 2460 5523
rect 2516 5517 2556 5523
rect 3012 5517 3116 5523
rect 3796 5517 3804 5523
rect 3812 5517 3836 5523
rect 3844 5517 3948 5523
rect 4020 5517 4412 5523
rect 5668 5517 5740 5523
rect 6372 5517 6380 5523
rect 6916 5517 7020 5523
rect 7716 5517 7804 5523
rect 7956 5517 8316 5523
rect 8452 5517 8524 5523
rect 8596 5517 8700 5523
rect 8708 5517 8860 5523
rect 9236 5517 9244 5523
rect 10164 5517 10268 5523
rect 10324 5517 10332 5523
rect 10532 5517 10540 5523
rect 11572 5517 11612 5523
rect 11780 5517 11804 5523
rect 12324 5517 12492 5523
rect 11837 5504 11843 5516
rect 708 5502 1075 5503
rect 708 5497 1068 5502
rect 1940 5497 1948 5503
rect 3252 5502 3667 5503
rect 3252 5497 3660 5502
rect 4580 5497 4588 5503
rect 7140 5497 7164 5503
rect 7172 5497 7516 5503
rect 7828 5497 7836 5503
rect 8836 5497 9132 5503
rect 9341 5502 9356 5503
rect 9348 5497 9356 5502
rect 10404 5497 10428 5503
rect 11300 5502 11475 5503
rect 11300 5497 11468 5502
rect 2452 5477 2572 5483
rect 2580 5477 3260 5483
rect 5860 5477 6380 5483
rect 7796 5477 7820 5483
rect 8388 5477 8428 5483
rect 8436 5477 8604 5483
rect 612 5457 620 5463
rect 1108 5457 1388 5463
rect 10116 5457 11036 5463
rect 5668 5437 5820 5443
rect 6292 5437 7804 5443
rect 8276 5437 8412 5443
rect 564 5417 572 5423
rect 3684 5417 3980 5423
rect 5780 5417 5820 5423
rect 5828 5417 6076 5423
rect 6420 5417 6588 5423
rect 52 5397 140 5403
rect 1732 5397 1964 5403
rect 6324 5397 8476 5403
rect 9652 5397 9676 5403
rect 740 5377 1164 5383
rect 4836 5377 6460 5383
rect 8996 5377 9724 5383
rect 9780 5377 9836 5383
rect 3332 5357 3340 5363
rect 9684 5357 9788 5363
rect 11716 5357 12268 5363
rect 132 5337 652 5343
rect 2596 5337 2620 5343
rect 6788 5337 7756 5343
rect 10404 5337 10636 5343
rect 10980 5337 11932 5343
rect 1748 5317 1900 5323
rect 2084 5318 2364 5323
rect 2084 5317 2371 5318
rect 2772 5318 2828 5323
rect 2772 5317 2835 5318
rect 3652 5317 3852 5323
rect 3860 5317 3980 5323
rect 5124 5317 5347 5323
rect 5341 5304 5347 5317
rect 6084 5318 6092 5323
rect 6084 5317 6099 5318
rect 7012 5317 7084 5323
rect 7220 5317 7228 5323
rect 9060 5317 9068 5323
rect 9076 5317 9180 5323
rect 10356 5317 10364 5323
rect 11684 5317 11708 5323
rect 12276 5317 12380 5323
rect 756 5297 1164 5303
rect 1828 5297 1836 5303
rect 2340 5297 2460 5303
rect 2484 5297 2492 5303
rect 2724 5297 2732 5303
rect 2756 5297 2812 5303
rect 3796 5297 3804 5303
rect 3812 5297 3820 5303
rect 3828 5297 3836 5303
rect 3844 5297 3948 5303
rect 4052 5297 4412 5303
rect 6004 5297 6140 5303
rect 7028 5297 7036 5303
rect 7300 5297 7420 5303
rect 8253 5297 8316 5303
rect 77 5284 83 5296
rect 212 5277 684 5283
rect 1876 5277 1884 5283
rect 1892 5277 3212 5283
rect 3773 5283 3779 5296
rect 3556 5277 3779 5283
rect 5844 5277 5948 5283
rect 6420 5277 7244 5283
rect 8253 5283 8259 5297
rect 9012 5297 9020 5303
rect 9620 5297 9644 5303
rect 9668 5297 9676 5303
rect 10228 5297 10268 5303
rect 10532 5297 10540 5303
rect 11844 5297 11852 5303
rect 12500 5297 12604 5303
rect 7748 5277 8259 5283
rect 8276 5277 8364 5283
rect 11565 5283 11571 5296
rect 10996 5277 11571 5283
rect 11620 5277 12348 5283
rect 12356 5277 12444 5283
rect 596 5257 700 5263
rect 2020 5257 2460 5263
rect 8980 5257 9052 5263
rect 9060 5257 9116 5263
rect 11748 5257 12220 5263
rect 4676 5237 5100 5243
rect 5460 5237 5820 5243
rect 5828 5237 9788 5243
rect 644 5217 732 5223
rect 2036 5217 2076 5223
rect 740 5197 748 5203
rect 2340 5197 2860 5203
rect 2868 5197 3324 5203
rect 4420 5197 4508 5203
rect 5812 5197 7068 5203
rect 7076 5197 8076 5203
rect 9012 5197 9180 5203
rect 3892 5177 4220 5183
rect 4484 5177 4524 5183
rect 5812 5177 5836 5183
rect 5844 5177 5932 5183
rect 7124 5177 7676 5183
rect 7684 5177 8860 5183
rect 9780 5177 9820 5183
rect 420 5157 636 5163
rect 644 5157 1708 5163
rect 4132 5157 7852 5163
rect 7860 5157 7948 5163
rect 9668 5157 9788 5163
rect 4004 5137 4684 5143
rect 7156 5137 7244 5143
rect 9613 5137 10172 5143
rect 9613 5124 9619 5137
rect 10996 5137 11203 5143
rect 11197 5124 11203 5137
rect 12285 5124 12291 5136
rect 148 5117 204 5123
rect 1172 5117 1180 5123
rect 1828 5117 1836 5123
rect 2340 5117 2460 5123
rect 2756 5117 3068 5123
rect 3236 5117 3324 5123
rect 4004 5117 4012 5123
rect 4692 5117 5020 5123
rect 5028 5117 5164 5123
rect 5284 5117 5324 5123
rect 5380 5117 6364 5123
rect 6452 5117 6556 5123
rect 6644 5117 6780 5123
rect 7300 5117 7388 5123
rect 7956 5117 7964 5123
rect 8884 5117 8972 5123
rect 10148 5117 10268 5123
rect 10548 5117 10684 5123
rect 11108 5117 11148 5123
rect 11732 5117 12220 5123
rect 1284 5097 1292 5103
rect 3188 5097 3276 5103
rect 4045 5103 4051 5116
rect 4004 5097 4051 5103
rect 4141 5102 4620 5103
rect 4148 5097 4620 5102
rect 5437 5102 5804 5103
rect 5444 5097 5804 5102
rect 5860 5097 5868 5103
rect 6733 5102 6748 5103
rect 6740 5097 6748 5102
rect 7076 5097 7180 5103
rect 9716 5102 10179 5103
rect 9716 5097 10172 5102
rect 10388 5097 10508 5103
rect 10573 5102 10579 5103
rect 12340 5097 12348 5103
rect 10573 5084 10579 5094
rect 2596 5077 2620 5083
rect 7796 5077 7820 5083
rect 4596 5057 4684 5063
rect 3988 5017 4044 5023
rect 4628 5017 4636 5023
rect 7748 5017 9068 5023
rect 1828 4997 3212 5003
rect 5124 4997 7644 5003
rect 8500 4997 8524 5003
rect 52 4977 508 4983
rect 1204 4977 3260 4983
rect 7140 4977 8572 4983
rect 12292 4977 12972 4983
rect 1252 4957 1363 4963
rect 564 4937 732 4943
rect 1357 4943 1363 4957
rect 1380 4957 1388 4963
rect 3860 4957 3868 4963
rect 6484 4957 6636 4963
rect 6644 4957 6675 4963
rect 1357 4937 1388 4943
rect 1885 4937 2028 4943
rect 1885 4924 1891 4937
rect 2516 4937 2636 4943
rect 5444 4937 6460 4943
rect 6669 4943 6675 4957
rect 8388 4957 8396 4963
rect 8420 4957 9116 4963
rect 12356 4957 12876 4963
rect 12916 4957 12924 4963
rect 6669 4937 6732 4943
rect 7796 4937 7820 4943
rect 9588 4937 9980 4943
rect 11636 4937 11932 4943
rect 1284 4917 1340 4923
rect 2580 4917 2684 4923
rect 3236 4917 3244 4923
rect 4532 4917 4540 4923
rect 5092 4917 5148 4923
rect 5332 4917 5347 4923
rect 5341 4904 5347 4917
rect 5428 4918 5436 4923
rect 5428 4917 5443 4918
rect 5492 4917 5772 4923
rect 5780 4917 5884 4923
rect 7780 4917 7836 4923
rect 8388 4917 8524 4923
rect 12340 4917 12380 4923
rect 468 4897 524 4903
rect 1172 4897 1196 4903
rect 1220 4897 1244 4903
rect 2388 4897 2460 4903
rect 3156 4897 3164 4903
rect 3764 4897 3772 4903
rect 3812 4897 3820 4903
rect 5060 4897 5068 4903
rect 5860 4897 5948 4903
rect 7604 4897 7660 4903
rect 7716 4897 7724 4903
rect 7732 4897 7900 4903
rect 7956 4897 7964 4903
rect 8532 4897 8588 4903
rect 8644 4897 9244 4903
rect 9293 4897 9308 4903
rect 5140 4877 5180 4883
rect 5188 4877 5196 4883
rect 5204 4877 5372 4883
rect 5997 4883 6003 4896
rect 5844 4877 6003 4883
rect 6452 4877 6572 4883
rect 7844 4877 8092 4883
rect 9293 4864 9299 4897
rect 10644 4897 11100 4903
rect 11188 4897 11196 4903
rect 11204 4897 11676 4903
rect 11700 4897 11804 4903
rect 11844 4897 11948 4903
rect 10404 4877 10476 4883
rect 100 4857 108 4863
rect 3220 4857 3324 4863
rect 3332 4857 4460 4863
rect 4468 4857 5068 4863
rect 5076 4857 5356 4863
rect 6548 4857 7900 4863
rect 11012 4857 11628 4863
rect 11652 4857 12300 4863
rect 12308 4857 12604 4863
rect 3316 4837 6988 4843
rect 6996 4837 7532 4843
rect 10868 4837 11660 4843
rect 2692 4817 4828 4823
rect 5924 4817 8652 4823
rect 10724 4817 11676 4823
rect 2692 4797 3020 4803
rect 3956 4797 4012 4803
rect 4964 4797 6748 4803
rect 7140 4797 7388 4803
rect 708 4777 1148 4783
rect 1892 4777 2524 4783
rect 2532 4777 3164 4783
rect 3172 4777 3788 4783
rect 3844 4777 4716 4783
rect 4724 4777 4924 4783
rect 5060 4777 5164 4783
rect 6388 4777 7132 4783
rect 7156 4777 7180 4783
rect 8269 4777 9820 4783
rect 3028 4757 5020 4763
rect 5044 4757 5196 4763
rect 8269 4763 8275 4777
rect 10340 4777 10476 4783
rect 5764 4757 8275 4763
rect 10404 4757 10428 4763
rect 484 4737 556 4743
rect 1220 4737 1308 4743
rect 1316 4737 1372 4743
rect 1892 4737 2044 4743
rect 2548 4737 2652 4743
rect 3076 4737 3164 4743
rect 3172 4737 3228 4743
rect 4420 4737 4460 4743
rect 7220 4737 7228 4743
rect 7396 4737 7404 4743
rect 7661 4737 7740 4743
rect 4685 4724 4691 4736
rect 7085 4724 7091 4736
rect 7661 4724 7667 4737
rect 8324 4737 8364 4743
rect 420 4717 524 4723
rect 1684 4717 1820 4723
rect 2100 4717 2188 4723
rect 3124 4717 3260 4723
rect 4420 4717 4428 4723
rect 4628 4717 4652 4723
rect 4660 4717 4668 4723
rect 5284 4717 5388 4723
rect 5396 4717 5900 4723
rect 5988 4717 5996 4723
rect 7028 4717 7036 4723
rect 8324 4717 8412 4723
rect 3389 4704 3395 4716
rect 1284 4697 1388 4703
rect 1396 4697 1580 4703
rect 1940 4697 1980 4703
rect 3236 4697 3244 4703
rect 3485 4702 3500 4703
rect 3492 4697 3500 4702
rect 6093 4702 6572 4703
rect 6100 4697 6572 4702
rect 8452 4697 8476 4703
rect 9293 4703 9299 4756
rect 10868 4737 10956 4743
rect 10980 4737 11020 4743
rect 11156 4737 11244 4743
rect 12228 4737 12316 4743
rect 10852 4717 10924 4723
rect 11204 4717 11292 4723
rect 12116 4717 12220 4723
rect 12269 4717 12284 4723
rect 9293 4697 9315 4703
rect 2196 4677 3292 4683
rect 8429 4683 8435 4696
rect 8429 4677 8444 4683
rect 9309 4683 9315 4697
rect 9332 4702 9347 4703
rect 9332 4697 9340 4702
rect 12269 4703 12275 4717
rect 11732 4697 12275 4703
rect 9309 4677 9324 4683
rect 11044 4677 11068 4683
rect 5108 4657 5324 4663
rect 10164 4657 11740 4663
rect 500 4617 2028 4623
rect 5508 4617 5820 4623
rect 7044 4617 7116 4623
rect 7412 4617 9020 4623
rect 9716 4617 9772 4623
rect 564 4597 5836 4603
rect 7780 4597 7820 4603
rect 8372 4597 9180 4603
rect 9700 4597 9708 4603
rect 10276 4597 11052 4603
rect -67 4577 92 4583
rect -67 4523 -61 4577
rect 3876 4577 11820 4583
rect -35 4557 12 4563
rect -35 4543 -29 4557
rect 1300 4557 4780 4563
rect 5460 4557 7228 4563
rect 7716 4557 7884 4563
rect 8756 4557 9084 4563
rect 9780 4557 9836 4563
rect -51 4537 -29 4543
rect 580 4537 732 4543
rect 1245 4524 1251 4536
rect -67 4517 -45 4523
rect 1124 4517 1171 4523
rect 1165 4504 1171 4517
rect 1588 4518 1724 4523
rect 1588 4517 1731 4518
rect 1812 4517 1884 4523
rect 3485 4504 3491 4518
rect 3828 4517 4003 4523
rect 3997 4504 4003 4517
rect 6436 4517 6444 4523
rect 6740 4518 6764 4523
rect 6733 4517 6764 4518
rect 7652 4517 7667 4523
rect 7661 4504 7667 4517
rect 8436 4517 8556 4523
rect 8676 4518 8684 4523
rect 8676 4517 8691 4518
rect 9748 4517 10348 4523
rect 12116 4517 12300 4523
rect 436 4497 524 4503
rect 564 4497 572 4503
rect 1204 4497 1212 4503
rect 1812 4497 1820 4503
rect 2756 4497 2860 4503
rect 3300 4497 3324 4503
rect 4612 4497 4652 4503
rect 4692 4497 4828 4503
rect 5348 4497 5452 4503
rect 5892 4497 6012 4503
rect 6372 4497 6380 4503
rect 6420 4497 6460 4503
rect 8308 4497 8316 4503
rect 9028 4497 9612 4503
rect 9668 4497 9708 4503
rect 9988 4497 10268 4503
rect 10468 4497 10483 4503
rect 10548 4497 10572 4503
rect 11204 4497 11564 4503
rect 12228 4497 12348 4503
rect 84 4477 1212 4483
rect 2461 4483 2467 4496
rect 2100 4477 2620 4483
rect 3389 4483 3395 4496
rect 3268 4477 3395 4483
rect 5252 4477 5276 4483
rect 6436 4477 6572 4483
rect 11524 4477 11612 4483
rect 1940 4457 2652 4463
rect 2692 4457 2812 4463
rect 8388 4437 8444 4443
rect 8452 4437 10684 4443
rect 52 4417 60 4423
rect 452 4417 732 4423
rect 1828 4417 1980 4423
rect 2484 4417 7724 4423
rect 8324 4417 8412 4423
rect 1812 4397 2028 4403
rect 11524 4397 11660 4403
rect 1348 4377 2444 4383
rect 3476 4377 3980 4383
rect 4180 4377 5436 4383
rect 6468 4377 6764 4383
rect 9044 4377 9180 4383
rect 11636 4377 11676 4383
rect 11684 4377 11932 4383
rect 3444 4357 3884 4363
rect 5812 4357 6460 4363
rect 9108 4357 9132 4363
rect 9668 4357 9820 4363
rect 10628 4357 11276 4363
rect 500 4337 556 4343
rect 2564 4337 3356 4343
rect 3117 4324 3123 4337
rect 5172 4337 5180 4343
rect 12356 4337 12499 4343
rect 12493 4324 12499 4337
rect 532 4317 556 4323
rect 1860 4317 1884 4323
rect 2468 4317 3100 4323
rect 3325 4317 3340 4323
rect 3396 4317 3516 4323
rect 3540 4317 4412 4323
rect 4420 4317 4428 4323
rect 4468 4317 4508 4323
rect 4948 4317 5068 4323
rect 5092 4317 5116 4323
rect 5124 4317 5132 4323
rect 5652 4317 5740 4323
rect 5812 4317 5827 4323
rect 1972 4302 2371 4303
rect 1972 4297 2364 4302
rect 1933 4203 1939 4296
rect 3332 4297 3468 4303
rect 5805 4284 5811 4296
rect 5821 4264 5827 4317
rect 6356 4317 6364 4323
rect 6404 4317 6412 4323
rect 6420 4317 6428 4323
rect 6644 4317 6652 4323
rect 7300 4317 7420 4323
rect 7780 4317 7900 4323
rect 8980 4317 8988 4323
rect 9604 4317 9612 4323
rect 10260 4317 10268 4323
rect 10324 4317 10332 4323
rect 10468 4317 10476 4323
rect 10548 4317 10684 4323
rect 10804 4317 11196 4323
rect 11716 4317 11804 4323
rect 11844 4317 11948 4323
rect 7949 4304 7955 4316
rect 6733 4302 6764 4303
rect 6740 4297 6764 4302
rect 7380 4302 7395 4303
rect 7380 4297 7388 4302
rect 7796 4297 7852 4303
rect 10340 4297 10348 4303
rect 10484 4297 10492 4303
rect 10500 4297 10572 4303
rect 7076 4277 7100 4283
rect 7428 4277 11212 4283
rect 11220 4277 11308 4283
rect 7092 4257 8492 4263
rect 10388 4257 10396 4263
rect 10564 4257 11020 4263
rect 5876 4237 8300 4243
rect 8436 4237 8700 4243
rect 3188 4217 3196 4223
rect 4164 4217 4524 4223
rect 5476 4217 7116 4223
rect 8884 4217 9020 4223
rect 1933 4197 1964 4203
rect 4420 4197 4476 4203
rect 5780 4197 6428 4203
rect 9604 4197 9708 4203
rect 10324 4197 10364 4203
rect 12436 4197 12444 4203
rect 1316 4177 1388 4183
rect 1860 4177 2028 4183
rect 7124 4177 7395 4183
rect 1229 4157 1340 4163
rect 1229 4143 1235 4157
rect 3156 4157 5932 4163
rect 1204 4137 1235 4143
rect 2596 4137 2620 4143
rect 3844 4137 4508 4143
rect 6740 4137 7372 4143
rect 1284 4117 1308 4123
rect 2836 4117 3004 4123
rect 3476 4118 3484 4123
rect 5149 4124 5155 4136
rect 3476 4117 3491 4118
rect 3828 4117 4003 4123
rect 3997 4104 4003 4117
rect 7389 4123 7395 4177
rect 10324 4177 10348 4183
rect 10452 4177 10476 4183
rect 11060 4177 11788 4183
rect 11012 4157 11020 4163
rect 11636 4157 12092 4163
rect 12948 4157 12972 4163
rect 11044 4137 11068 4143
rect 11108 4137 11676 4143
rect 11716 4137 12236 4143
rect 12372 4137 12876 4143
rect 7389 4117 7411 4123
rect 532 4097 588 4103
rect 1828 4097 1868 4103
rect 2500 4097 2508 4103
rect 2516 4097 2524 4103
rect 2532 4097 2604 4103
rect 2756 4097 2876 4103
rect 3188 4097 3324 4103
rect 3380 4097 3388 4103
rect 4964 4097 5068 4103
rect 5140 4097 5148 4103
rect 5204 4097 5340 4103
rect 6244 4097 6364 4103
rect 6372 4097 6380 4103
rect 6628 4097 6636 4103
rect 7293 4084 7299 4096
rect 516 4077 556 4083
rect 2324 4077 2700 4083
rect 2708 4077 3132 4083
rect 4516 4077 6636 4083
rect 6724 4077 7244 4083
rect 7405 4064 7411 4117
rect 7732 4117 7836 4123
rect 8516 4117 9132 4123
rect 9988 4118 10428 4123
rect 9981 4117 10428 4118
rect 10660 4117 11004 4123
rect 11012 4117 11020 4123
rect 12100 4117 12300 4123
rect 8580 4097 8588 4103
rect 9188 4097 9244 4103
rect 9892 4097 9916 4103
rect 10804 4097 10924 4103
rect 11204 4097 11276 4103
rect 7796 4077 7900 4083
rect 8548 4077 9196 4083
rect 9860 4077 9932 4083
rect 11732 4077 12284 4083
rect 180 4057 684 4063
rect 2628 4057 4044 4063
rect 7092 4057 7100 4063
rect 12164 4057 12396 4063
rect 500 4037 572 4043
rect 2612 4037 3180 4043
rect 3204 4037 3292 4043
rect 4612 4037 5292 4043
rect 6964 4037 7139 4043
rect 1172 4017 1228 4023
rect 2468 4017 2636 4023
rect 2644 4017 5452 4023
rect 7133 4023 7139 4037
rect 7316 4037 11148 4043
rect 7133 4017 7788 4023
rect 7812 4017 8412 4023
rect 916 3997 1372 4003
rect 1828 3997 3836 4003
rect 3844 3997 4956 4003
rect 5076 3997 5900 4003
rect 5908 3997 7196 4003
rect 2564 3977 2668 3983
rect 2676 3977 3468 3983
rect 5965 3977 9996 3983
rect 5965 3963 5971 3977
rect 3188 3957 5971 3963
rect 7748 3957 7932 3963
rect 7940 3957 7948 3963
rect 8324 3957 9132 3963
rect 9668 3957 9788 3963
rect 1892 3937 2860 3943
rect 3332 3937 3340 3943
rect 4685 3937 5100 3943
rect 4685 3924 4691 3937
rect 5220 3937 5276 3943
rect 6068 3937 6572 3943
rect 84 3917 92 3923
rect 148 3917 172 3923
rect 804 3917 1100 3923
rect 1108 3917 1324 3923
rect 3124 3917 3148 3923
rect 3172 3917 3196 3923
rect 4052 3917 4316 3923
rect 4548 3917 4604 3923
rect 5348 3917 5452 3923
rect 6132 3917 6364 3923
rect 6628 3917 6636 3923
rect 644 3897 684 3903
rect 893 3902 1676 3903
rect 900 3897 1676 3902
rect 1940 3897 1996 3903
rect 2093 3903 2099 3916
rect 2084 3897 2099 3903
rect 5124 3897 5228 3903
rect 6397 3903 6403 3916
rect 6340 3897 6403 3903
rect 6484 3897 6492 3903
rect 132 3877 652 3883
rect 1684 3877 3484 3883
rect 3492 3877 3660 3883
rect 7405 3863 7411 3956
rect 8372 3937 8460 3943
rect 8468 3937 8524 3943
rect 10925 3937 11004 3943
rect 10925 3924 10931 3937
rect 11620 3937 12300 3943
rect 12852 3937 12908 3943
rect 9204 3917 9612 3923
rect 9636 3917 10268 3923
rect 10276 3917 10284 3923
rect 10964 3917 11052 3923
rect 11460 3917 11564 3923
rect 11604 3917 11612 3923
rect 11684 3917 11820 3923
rect 11828 3917 11836 3923
rect 12868 3917 12940 3923
rect 8436 3897 8540 3903
rect 8692 3902 8867 3903
rect 8692 3897 8860 3902
rect 9732 3897 9836 3903
rect 10004 3902 10179 3903
rect 10004 3897 10172 3902
rect 11028 3897 11100 3903
rect 11684 3897 11987 3903
rect 8548 3877 8684 3883
rect 10420 3877 10924 3883
rect 11316 3877 11852 3883
rect 11860 3877 11964 3883
rect 11981 3883 11987 3897
rect 11981 3877 12268 3883
rect 7396 3857 7411 3863
rect 10852 3857 11740 3863
rect 3828 3817 3836 3823
rect 6420 3817 6428 3823
rect 8420 3817 8540 3823
rect 9188 3817 9196 3823
rect 52 3797 60 3803
rect 5940 3797 5948 3803
rect 5172 3777 6364 3783
rect 8388 3777 8508 3783
rect 6644 3757 9180 3763
rect 5844 3737 5868 3743
rect 8644 3737 9516 3743
rect 900 3718 908 3723
rect 893 3717 908 3718
rect 2020 3717 2060 3723
rect 2516 3717 3123 3723
rect 3117 3704 3123 3717
rect 3236 3717 3324 3723
rect 4132 3718 4140 3723
rect 4132 3717 4147 3718
rect 3156 3697 3164 3703
rect 3396 3697 3628 3703
rect 3860 3697 4044 3703
rect 4628 3697 4652 3703
rect 4660 3697 4668 3703
rect 1437 3683 1443 3696
rect 1252 3677 1443 3683
rect 2093 3683 2099 3696
rect 1956 3677 2099 3683
rect 4685 3683 4691 3696
rect 4484 3677 4691 3683
rect 5645 3683 5651 3736
rect 8621 3724 8627 3736
rect 5956 3717 6515 3723
rect 6004 3697 6124 3703
rect 6509 3703 6515 3717
rect 6621 3717 6716 3723
rect 6509 3697 6604 3703
rect 6621 3703 6627 3717
rect 8532 3717 8572 3723
rect 9732 3717 9740 3723
rect 9860 3718 9980 3723
rect 9860 3717 9987 3718
rect 6612 3697 6627 3703
rect 6644 3697 6748 3703
rect 7405 3697 7948 3703
rect 5645 3677 5788 3683
rect 5844 3677 6508 3683
rect 7405 3683 7411 3697
rect 8596 3697 8732 3703
rect 9620 3697 9628 3703
rect 9869 3684 9875 3696
rect 6596 3677 7411 3683
rect 9997 3664 10003 3856
rect 11668 3817 11804 3823
rect 12276 3817 12316 3823
rect 10420 3797 10428 3803
rect 11636 3777 11756 3783
rect 11972 3737 12300 3743
rect 12308 3737 12588 3743
rect 12596 3737 12764 3743
rect 12308 3717 12316 3723
rect 10548 3697 10972 3703
rect 12292 3697 12364 3703
rect 10340 3677 10476 3683
rect 10996 3677 11148 3683
rect 1380 3657 2588 3663
rect 5860 3657 5948 3663
rect 5956 3657 7900 3663
rect 10996 3657 12220 3663
rect 1716 3637 2332 3643
rect 2340 3637 4588 3643
rect 4660 3637 5196 3643
rect 516 3617 572 3623
rect 3140 3617 5324 3623
rect 5332 3617 5756 3623
rect 5764 3617 6780 3623
rect 6804 3617 8988 3623
rect 8996 3617 11100 3623
rect 564 3597 636 3603
rect 532 3577 1372 3583
rect 7716 3577 7724 3583
rect 12308 3577 12428 3583
rect 12292 3557 12380 3563
rect 1220 3537 1292 3543
rect 3188 3537 3324 3543
rect 5412 3537 5948 3543
rect 5956 3537 6060 3543
rect 7396 3537 9756 3543
rect 84 3517 92 3523
rect 148 3517 156 3523
rect 1140 3517 1164 3523
rect 1700 3517 1820 3523
rect 1828 3517 1852 3523
rect 3780 3517 3932 3523
rect 4052 3517 4172 3523
rect 4628 3517 4652 3523
rect 4692 3517 4844 3523
rect 5348 3517 5692 3523
rect 6004 3517 6092 3523
rect 6500 3517 6572 3523
rect 6580 3517 6604 3523
rect 6612 3517 6620 3523
rect 7300 3517 7436 3523
rect 7812 3517 7900 3523
rect 8429 3517 8524 3523
rect 3117 3503 3123 3516
rect 3117 3497 3132 3503
rect 3220 3497 3532 3503
rect 4797 3502 4803 3503
rect 1933 3483 1939 3496
rect 6436 3497 6540 3503
rect 7396 3497 7756 3503
rect 8429 3503 8435 3517
rect 9181 3523 9187 3537
rect 10004 3537 11203 3543
rect 11197 3524 11203 3537
rect 9181 3517 9244 3523
rect 9284 3517 10268 3523
rect 10324 3517 10332 3523
rect 10356 3517 10444 3523
rect 10452 3517 10540 3523
rect 10612 3517 11148 3523
rect 11156 3517 11180 3523
rect 12228 3517 12236 3523
rect 8388 3497 8435 3503
rect 8452 3497 8476 3503
rect 9076 3497 9132 3503
rect 10356 3497 10371 3503
rect 4797 3484 4803 3494
rect 1933 3477 2364 3483
rect 2372 3477 3228 3483
rect 3364 3477 3532 3483
rect 3540 3477 3660 3483
rect 4125 3477 4140 3483
rect 3924 3457 4028 3463
rect 4125 3443 4131 3477
rect 7732 3477 7756 3483
rect 7764 3477 7964 3483
rect 9092 3477 9276 3483
rect 5364 3457 6124 3463
rect 9684 3457 9708 3463
rect 3940 3437 4131 3443
rect 7140 3437 7148 3443
rect 9572 3437 9708 3443
rect 52 3397 60 3403
rect 3300 3397 3340 3403
rect 3988 3397 3996 3403
rect 532 3377 5868 3383
rect 1268 3357 1388 3363
rect 1956 3357 2028 3363
rect 6436 3357 6588 3363
rect 9028 3357 9132 3363
rect 9796 3357 9820 3363
rect 564 3337 732 3343
rect 1885 3337 1980 3343
rect 1885 3324 1891 3337
rect 2596 3337 2620 3343
rect 2740 3337 3228 3343
rect 3236 3337 3244 3343
rect 3252 3337 3260 3343
rect 4717 3337 5228 3343
rect 1284 3317 1340 3323
rect 1940 3317 1948 3323
rect 1972 3317 2060 3323
rect 2676 3317 2684 3323
rect 2717 3317 2780 3323
rect 2717 3304 2723 3317
rect 3188 3317 3395 3323
rect 3389 3304 3395 3317
rect 4212 3317 4316 3323
rect 4717 3323 4723 3337
rect 9124 3337 9628 3343
rect 9716 3337 9852 3343
rect 9860 3337 9980 3343
rect 4669 3317 4723 3323
rect 4669 3304 4675 3317
rect 6484 3317 6540 3323
rect 7092 3317 7100 3323
rect 7396 3318 7420 3323
rect 7389 3317 7420 3318
rect 7444 3317 7580 3323
rect 7588 3317 7724 3323
rect 7732 3317 7836 3323
rect 9997 3323 10003 3496
rect 10365 3463 10371 3497
rect 10388 3497 10428 3503
rect 11092 3497 11116 3503
rect 10644 3477 10652 3483
rect 10365 3457 10380 3463
rect 10324 3397 10492 3403
rect 11636 3397 11644 3403
rect 11780 3397 11788 3403
rect 12244 3397 12972 3403
rect 10964 3357 11132 3363
rect 11732 3357 11740 3363
rect 11060 3337 11580 3343
rect 9885 3317 10003 3323
rect 9885 3304 9891 3317
rect 11060 3317 11603 3323
rect 11597 3304 11603 3317
rect 11652 3317 11923 3323
rect 1220 3297 1260 3303
rect 1748 3297 1820 3303
rect 2468 3297 2540 3303
rect 2756 3297 2860 3303
rect 2877 3297 3324 3303
rect 2877 3283 2883 3297
rect 3940 3297 4060 3303
rect 4692 3297 4796 3303
rect 6292 3297 6364 3303
rect 6420 3297 6428 3303
rect 7028 3297 7068 3303
rect 7812 3297 7900 3303
rect 7956 3297 7996 3303
rect 8381 3297 8972 3303
rect 8381 3284 8387 3297
rect 9012 3297 9020 3303
rect 9620 3297 9692 3303
rect 10436 3297 10924 3303
rect 11444 3297 11564 3303
rect 11620 3297 11628 3303
rect 11636 3297 11836 3303
rect 11917 3303 11923 3317
rect 12276 3317 12380 3323
rect 11917 3297 12492 3303
rect 2516 3277 2883 3283
rect 3300 3277 3308 3283
rect 3940 3277 3980 3283
rect 4516 3277 5180 3283
rect 7092 3277 7804 3283
rect 9572 3277 9660 3283
rect 9668 3277 9852 3283
rect 9860 3277 9916 3283
rect 12356 3277 12444 3283
rect 100 3257 1740 3263
rect 1892 3257 1980 3263
rect 2020 3257 2508 3263
rect 9716 3257 11196 3263
rect 756 3237 3516 3243
rect 11044 3237 11052 3243
rect 12852 3217 12924 3223
rect 4836 3197 5228 3203
rect 11204 3197 11660 3203
rect 4644 3177 4796 3183
rect 5828 3177 5932 3183
rect 10340 3177 10492 3183
rect 1556 3157 2028 3163
rect 2468 3157 2620 3163
rect 3284 3157 3372 3163
rect 4468 3157 4588 3163
rect 5764 3157 5868 3163
rect 6788 3157 7692 3163
rect 7700 3157 7900 3163
rect 7908 3157 9388 3163
rect 10996 3157 11196 3163
rect 3236 3137 4652 3143
rect 6580 3137 6620 3143
rect 7156 3137 7244 3143
rect 8020 3137 8524 3143
rect 9044 3137 9196 3143
rect 9348 3137 9932 3143
rect 9940 3137 10476 3143
rect 10484 3137 10604 3143
rect 11652 3137 11772 3143
rect 11780 3137 11804 3143
rect 12356 3137 12499 3143
rect 12493 3124 12499 3137
rect 1444 3117 1548 3123
rect 2500 3117 2508 3123
rect 2516 3117 2524 3123
rect 2532 3117 2572 3123
rect 4340 3117 4412 3123
rect 4509 3117 5068 3123
rect 1380 3097 1388 3103
rect 2580 3097 2684 3103
rect 3636 3102 3667 3103
rect 3636 3097 3660 3102
rect 4509 3103 4515 3117
rect 6276 3117 6364 3123
rect 6372 3117 6380 3123
rect 6420 3117 6428 3123
rect 6468 3117 6604 3123
rect 7300 3117 7804 3123
rect 7940 3117 7948 3123
rect 7956 3117 8044 3123
rect 8532 3117 8540 3123
rect 8596 3117 8732 3123
rect 9828 3117 10268 3123
rect 10548 3117 10636 3123
rect 11748 3117 11836 3123
rect 12436 3117 12444 3123
rect 4084 3097 4515 3103
rect 4532 3097 4636 3103
rect 4660 3102 4979 3103
rect 4660 3097 4972 3102
rect 5188 3097 5276 3103
rect 6580 3097 6588 3103
rect 7076 3097 7180 3103
rect 8388 3097 8476 3103
rect 10388 3097 10412 3103
rect 10637 3102 11084 3103
rect 10644 3097 11084 3102
rect 11293 3102 11308 3103
rect 11300 3097 11308 3102
rect 12434 3097 12460 3103
rect 644 3077 668 3083
rect 6388 3077 7964 3083
rect 7972 3077 8028 3083
rect 8452 3077 8540 3083
rect 9764 3077 10284 3083
rect 11700 3077 11852 3083
rect 11860 3077 11964 3083
rect 6548 3057 6620 3063
rect 7844 3057 7996 3063
rect 8548 3037 9347 3043
rect 52 3017 156 3023
rect 3284 3017 3292 3023
rect 9060 3017 9068 3023
rect 1236 2997 2092 3003
rect 1348 2977 1404 2983
rect 612 2957 668 2963
rect 6436 2957 7708 2963
rect 7732 2957 7964 2963
rect 621 2937 732 2943
rect 621 2924 627 2937
rect 740 2937 748 2943
rect 1332 2937 2348 2943
rect 5124 2937 5340 2943
rect 708 2918 1068 2923
rect 708 2917 1075 2918
rect 1908 2917 1948 2923
rect 2532 2917 2636 2923
rect 4532 2917 4540 2923
rect 4788 2918 4812 2923
rect 4781 2917 4812 2918
rect 7108 2917 7116 2923
rect 7220 2917 7228 2923
rect 8580 2918 8684 2923
rect 8692 2918 9132 2923
rect 8580 2917 9132 2918
rect 9341 2923 9347 3037
rect 11620 3017 11628 3023
rect 11652 2957 12316 2963
rect 11284 2937 11292 2943
rect 11300 2937 11932 2943
rect 11085 2924 11091 2936
rect 9245 2917 9347 2923
rect 9245 2904 9251 2917
rect 10324 2917 10476 2923
rect 11956 2918 11964 2923
rect 11949 2917 11964 2918
rect 516 2897 524 2903
rect 564 2897 604 2903
rect 1108 2897 1164 2903
rect 1812 2897 1820 2903
rect 2052 2897 2060 2903
rect 2532 2897 2748 2903
rect 4324 2897 4412 2903
rect 4468 2897 4620 2903
rect 4692 2897 4796 2903
rect 5268 2897 5276 2903
rect 5844 2897 5948 2903
rect 6964 2897 7084 2903
rect 7092 2897 7100 2903
rect 8228 2897 8316 2903
rect 8516 2897 8540 2903
rect 8596 2897 8684 2903
rect 9188 2897 9196 2903
rect 10548 2897 10556 2903
rect 11204 2897 11308 2903
rect 11780 2897 11804 2903
rect 11812 2897 11820 2903
rect 1764 2877 1884 2883
rect 2052 2877 2236 2883
rect 2596 2877 2700 2883
rect 3844 2877 3852 2883
rect 5300 2877 6924 2883
rect 9764 2877 9852 2883
rect 2020 2857 2124 2863
rect 2132 2857 2300 2863
rect 3860 2857 3884 2863
rect 5908 2857 6028 2863
rect 7204 2857 7452 2863
rect 4852 2837 5292 2843
rect 5300 2837 6476 2843
rect 10996 2837 11276 2843
rect 11284 2837 11948 2843
rect 5940 2817 6044 2823
rect 11620 2817 11772 2823
rect 1812 2797 2028 2803
rect 4836 2797 6492 2803
rect 7076 2797 7868 2803
rect 9044 2797 9180 2803
rect 10340 2797 10796 2803
rect 1268 2777 1372 2783
rect 2436 2777 2684 2783
rect 2692 2777 3052 2783
rect 3988 2777 4076 2783
rect 6916 2777 9052 2783
rect 532 2757 668 2763
rect 1220 2757 1340 2763
rect 2644 2757 2668 2763
rect 2676 2757 3324 2763
rect 3332 2757 3420 2763
rect 5204 2757 5340 2763
rect 6420 2757 6572 2763
rect 7108 2757 7820 2763
rect 8372 2757 8524 2763
rect 9108 2757 9132 2763
rect 2196 2737 2508 2743
rect 2516 2737 4780 2743
rect 4685 2724 4691 2737
rect 4797 2737 5916 2743
rect 1828 2717 3004 2723
rect 4420 2717 4428 2723
rect 4468 2717 4588 2723
rect 4644 2717 4652 2723
rect 4797 2723 4803 2737
rect 7588 2737 7708 2743
rect 7780 2737 7788 2743
rect 8132 2737 9820 2743
rect 9828 2737 9852 2743
rect 9860 2737 10348 2743
rect 10484 2737 10588 2743
rect 4708 2717 4803 2723
rect 6276 2717 6364 2723
rect 7668 2717 8012 2723
rect 9524 2717 9612 2723
rect 9860 2717 9868 2723
rect 9892 2717 9916 2723
rect 10548 2717 10636 2723
rect 10644 2717 11004 2723
rect 11572 2717 11644 2723
rect 11668 2717 11724 2723
rect 3117 2683 3123 2716
rect 3485 2702 3548 2703
rect 3492 2697 3548 2702
rect 4532 2697 4636 2703
rect 6356 2702 6931 2703
rect 6356 2697 6924 2702
rect 7780 2697 7788 2703
rect 10404 2697 10428 2703
rect 10637 2702 11548 2703
rect 10644 2697 11548 2702
rect 3117 2677 4204 2683
rect 7028 2677 7564 2683
rect 3268 2657 3388 2663
rect 6116 2637 7228 2643
rect 7236 2637 8732 2643
rect 468 2617 620 2623
rect 1172 2617 1388 2623
rect 3140 2617 3340 2623
rect 3972 2617 3980 2623
rect 5924 2617 5932 2623
rect 8980 2617 9068 2623
rect 10052 2617 11788 2623
rect 84 2597 92 2603
rect 564 2597 636 2603
rect 4596 2597 4764 2603
rect 9668 2597 9708 2603
rect 9748 2597 10364 2603
rect 11636 2597 11836 2603
rect 12276 2597 12284 2603
rect 628 2577 732 2583
rect 3844 2577 5276 2583
rect 9684 2577 9708 2583
rect 3988 2557 5804 2563
rect 8372 2557 8380 2563
rect 8388 2557 8428 2563
rect 9165 2557 10492 2563
rect 132 2537 652 2543
rect 1204 2537 2028 2543
rect 2596 2537 2620 2543
rect 3012 2537 3804 2543
rect 3812 2537 5244 2543
rect 5252 2537 5996 2543
rect 7796 2537 7820 2543
rect 8692 2537 8700 2543
rect 9165 2543 9171 2557
rect 11028 2557 11036 2563
rect 8708 2537 9171 2543
rect 10052 2537 10380 2543
rect 11044 2537 11068 2543
rect 1284 2517 1292 2523
rect 3844 2517 3852 2523
rect 4820 2517 5148 2523
rect 5828 2517 5852 2523
rect 6132 2518 6268 2523
rect 6740 2518 6748 2523
rect 6132 2517 6275 2518
rect 6733 2517 6748 2518
rect 6932 2517 7212 2523
rect 7220 2518 7564 2523
rect 7220 2517 7571 2518
rect 7796 2517 7836 2523
rect 8052 2518 8172 2523
rect 8045 2517 8172 2518
rect 8436 2517 8595 2523
rect 8589 2504 8595 2517
rect 9124 2517 9132 2523
rect 9828 2518 9980 2523
rect 9828 2517 9987 2518
rect 12356 2517 12380 2523
rect 148 2497 252 2503
rect 1156 2497 1164 2503
rect 1716 2497 1820 2503
rect 2356 2497 2460 2503
rect 2468 2497 2476 2503
rect 2692 2497 2700 2503
rect 2708 2497 2716 2503
rect 2756 2497 2796 2503
rect 3796 2497 3804 2503
rect 3812 2497 3836 2503
rect 3988 2497 4316 2503
rect 4324 2497 4412 2503
rect 4628 2497 4940 2503
rect 4964 2497 5068 2503
rect 5092 2497 5132 2503
rect 6356 2497 6364 2503
rect 7540 2497 7660 2503
rect 7700 2497 7948 2503
rect 8532 2497 8572 2503
rect 9252 2497 9372 2503
rect 10932 2497 10940 2503
rect 11188 2497 11196 2503
rect 1885 2484 1891 2496
rect 1220 2477 1756 2483
rect 2516 2477 3468 2483
rect 3476 2477 6428 2483
rect 9796 2477 9820 2483
rect 12292 2477 12444 2483
rect 2564 2457 3292 2463
rect 3300 2457 5244 2463
rect 5252 2457 6604 2463
rect 7748 2457 9884 2463
rect 12324 2457 12444 2463
rect 8436 2437 12492 2443
rect 260 2417 620 2423
rect 1108 2417 2028 2423
rect 3156 2417 3180 2423
rect 3300 2417 3324 2423
rect 3764 2417 3772 2423
rect 3780 2417 3948 2423
rect 3956 2417 3980 2423
rect 6468 2417 7916 2423
rect 12292 2417 12412 2423
rect 2708 2397 4668 2403
rect 4676 2397 5276 2403
rect 8916 2397 10428 2403
rect 1268 2377 1372 2383
rect 4708 2377 5804 2383
rect 8388 2377 8428 2383
rect 9044 2377 11836 2383
rect 260 2357 636 2363
rect 1220 2357 1340 2363
rect 2516 2357 2668 2363
rect 4932 2357 7100 2363
rect 7108 2357 9980 2363
rect 10964 2357 11132 2363
rect 84 2337 156 2343
rect 3076 2337 3164 2343
rect 3181 2337 3324 2343
rect 148 2317 252 2323
rect 1172 2317 1196 2323
rect 1828 2317 1836 2323
rect 1940 2317 2188 2323
rect 3124 2317 3164 2323
rect 3181 2323 3187 2337
rect 4996 2337 5132 2343
rect 5140 2337 5148 2343
rect 7092 2337 7299 2343
rect 5277 2324 5283 2336
rect 3172 2317 3187 2323
rect 3636 2317 3772 2323
rect 3812 2317 3884 2323
rect 3956 2317 4412 2323
rect 4420 2317 4700 2323
rect 4804 2317 5068 2323
rect 5140 2317 5260 2323
rect 5293 2323 5299 2336
rect 7293 2324 7299 2337
rect 7540 2337 7900 2343
rect 7908 2337 7996 2343
rect 11572 2337 11612 2343
rect 5293 2317 5340 2323
rect 5940 2317 5948 2323
rect 6004 2317 6108 2323
rect 7812 2317 7948 2323
rect 8596 2317 8604 2323
rect 9252 2317 9260 2323
rect 10157 2317 10268 2323
rect 2461 2303 2467 2316
rect 2036 2297 2467 2303
rect 2580 2297 2604 2303
rect 3236 2297 3244 2303
rect 4692 2297 4940 2303
rect 4964 2302 4979 2303
rect 4964 2297 4972 2302
rect 5188 2297 5692 2303
rect 5860 2297 5884 2303
rect 6436 2297 6540 2303
rect 8013 2302 8019 2316
rect 8180 2297 8476 2303
rect 8484 2297 8508 2303
rect 8685 2302 9132 2303
rect 8692 2297 9132 2302
rect 9341 2302 9580 2303
rect 9348 2297 9580 2302
rect 10157 2303 10163 2317
rect 10324 2317 10332 2323
rect 11044 2317 11564 2323
rect 11780 2317 11804 2323
rect 11812 2317 11820 2323
rect 9684 2297 10163 2303
rect 11028 2297 11052 2303
rect 1300 2277 1724 2283
rect 7140 2277 7164 2283
rect 8388 2277 8428 2283
rect 3124 2257 3228 2263
rect 9028 2257 9052 2263
rect 9684 2257 12220 2263
rect 52 2217 508 2223
rect 10324 2197 10364 2203
rect 1172 2177 1388 2183
rect 6500 2177 6588 2183
rect 10324 2177 10380 2183
rect 1268 2157 2028 2163
rect 2804 2157 3260 2163
rect 3268 2157 3980 2163
rect 6429 2157 6540 2163
rect 564 2137 732 2143
rect 1204 2137 1980 2143
rect 2596 2137 2620 2143
rect 5780 2137 5788 2143
rect 6429 2143 6435 2157
rect 7156 2157 7228 2163
rect 11684 2157 11875 2163
rect 6420 2137 6435 2143
rect 7085 2137 7180 2143
rect 1908 2117 1980 2123
rect 2564 2117 2620 2123
rect 2717 2117 2796 2123
rect 2717 2104 2723 2117
rect 3341 2124 3347 2136
rect 5149 2124 5155 2136
rect 7085 2124 7091 2137
rect 7796 2137 7820 2143
rect 8644 2137 9980 2143
rect 9988 2137 10636 2143
rect 11869 2143 11875 2157
rect 11869 2137 11932 2143
rect 11940 2137 11948 2143
rect 2852 2118 2956 2123
rect 2845 2117 2956 2118
rect 3860 2117 4204 2123
rect 4532 2117 4540 2123
rect 4548 2117 4988 2123
rect 6484 2117 6492 2123
rect 7140 2117 7148 2123
rect 7204 2118 7564 2123
rect 7204 2117 7571 2118
rect 7796 2117 7804 2123
rect 7828 2117 7836 2123
rect 9172 2117 9340 2123
rect 10980 2117 11084 2123
rect 180 2097 524 2103
rect 1268 2097 1820 2103
rect 1828 2097 1836 2103
rect 1892 2097 1900 2103
rect 2564 2097 2668 2103
rect 2756 2097 2844 2103
rect 3844 2097 3916 2103
rect 5076 2097 5100 2103
rect 5348 2097 5356 2103
rect 5892 2097 6140 2103
rect 6308 2097 6364 2103
rect 6916 2097 7020 2103
rect 7652 2097 7660 2103
rect 7956 2097 8060 2103
rect 9252 2097 9260 2103
rect 10148 2097 10540 2103
rect 10548 2097 10684 2103
rect 11204 2097 11308 2103
rect 11780 2097 11836 2103
rect 4413 2084 4419 2096
rect 1924 2077 2028 2083
rect 2436 2077 2508 2083
rect 2580 2077 2620 2083
rect 2964 2077 3900 2083
rect 4468 2077 4956 2083
rect 5284 2077 5388 2083
rect 5396 2077 6412 2083
rect 8532 2077 8636 2083
rect 11044 2077 11148 2083
rect 11652 2077 11772 2083
rect 11780 2077 11804 2083
rect 2036 2057 2108 2063
rect 6276 2057 8492 2063
rect 10356 2057 11100 2063
rect 100 2037 156 2043
rect 436 2037 5955 2043
rect 3220 2017 3820 2023
rect 3828 2017 3948 2023
rect 5828 2017 5932 2023
rect 5949 2023 5955 2037
rect 6292 2037 10444 2043
rect 12212 2037 12316 2043
rect 5949 2017 7788 2023
rect 52 1997 140 2003
rect 5796 1997 6380 2003
rect 6612 1997 9196 2003
rect 9204 1997 10428 2003
rect 11316 1997 11628 2003
rect 3300 1977 3804 1983
rect 5796 1977 5852 1983
rect 7652 1977 7724 1983
rect 532 1957 732 1963
rect 2516 1957 2668 1963
rect 3188 1957 4028 1963
rect 8324 1957 10348 1963
rect 10948 1957 12268 1963
rect 484 1937 556 1943
rect 1220 1937 1356 1943
rect 3972 1937 5276 1943
rect 5325 1937 6371 1943
rect 1108 1917 1164 1923
rect 1284 1917 1404 1923
rect 1444 1917 1644 1923
rect 2388 1917 2460 1923
rect 3028 1917 3116 1923
rect 3325 1923 3331 1936
rect 3325 1917 3340 1923
rect 3396 1917 3500 1923
rect 3933 1923 3939 1936
rect 3508 1917 3980 1923
rect 4612 1917 4652 1923
rect 5325 1923 5331 1937
rect 6365 1924 6371 1937
rect 7156 1937 7228 1943
rect 9044 1937 9251 1943
rect 9245 1924 9251 1937
rect 10500 1937 10956 1943
rect 11012 1937 11148 1943
rect 11197 1924 11203 1936
rect 5204 1917 5331 1923
rect 6420 1917 6524 1923
rect 6532 1917 6604 1923
rect 8372 1917 8380 1923
rect 8980 1917 8988 1923
rect 9012 1917 9036 1923
rect 9876 1917 9884 1923
rect 10932 1917 10940 1923
rect 11588 1917 11820 1923
rect 11828 1917 11836 1923
rect 1892 1897 2028 1903
rect 3332 1897 3468 1903
rect 4685 1903 4691 1916
rect 4484 1897 4691 1903
rect 9124 1897 9132 1903
rect 1556 1877 1948 1883
rect 1956 1877 3964 1883
rect 5204 1877 5276 1883
rect 7812 1877 8332 1883
rect 8429 1864 8435 1896
rect 3940 1857 4044 1863
rect 5124 1857 5132 1863
rect 7524 1837 7948 1843
rect 1668 1817 1868 1823
rect 3988 1817 3996 1823
rect 6452 1817 6460 1823
rect 8388 1817 8540 1823
rect 52 1797 172 1803
rect 484 1797 668 1803
rect 6404 1797 6428 1803
rect 2628 1777 4556 1783
rect 9732 1777 10924 1783
rect 628 1757 732 1763
rect 3908 1757 5171 1763
rect 4548 1737 4780 1743
rect 4788 1737 4812 1743
rect 5165 1743 5171 1757
rect 7796 1757 9244 1763
rect 11044 1757 11132 1763
rect 5165 1737 5436 1743
rect 5780 1737 6060 1743
rect 8052 1737 9340 1743
rect 9348 1737 9724 1743
rect 10333 1737 10492 1743
rect 10333 1724 10339 1737
rect 11028 1737 11468 1743
rect 1284 1717 1292 1723
rect 3188 1717 3196 1723
rect 3860 1717 3900 1723
rect 4564 1717 5276 1723
rect 5341 1717 5804 1723
rect 5341 1704 5347 1717
rect 7076 1717 7180 1723
rect 11028 1717 11036 1723
rect 11837 1704 11843 1716
rect 468 1697 524 1703
rect 1380 1697 1404 1703
rect 1412 1697 1420 1703
rect 2372 1697 2460 1703
rect 3796 1697 3804 1703
rect 3812 1697 3836 1703
rect 4420 1697 4684 1703
rect 4692 1697 4828 1703
rect 6004 1697 6124 1703
rect 7300 1697 7420 1703
rect 7892 1697 7900 1703
rect 7908 1697 7916 1703
rect 8996 1697 9004 1703
rect 10260 1697 10268 1703
rect 10916 1697 10924 1703
rect 10948 1697 10956 1703
rect 10964 1697 10988 1703
rect 10996 1697 11052 1703
rect 11572 1697 11580 1703
rect 484 1677 556 1683
rect 1437 1683 1443 1696
rect 1437 1677 1868 1683
rect 2516 1677 2636 1683
rect 4372 1677 4460 1683
rect 4628 1677 4652 1683
rect 7156 1677 7244 1683
rect 7844 1677 7852 1683
rect 9012 1677 9036 1683
rect 9213 1683 9219 1696
rect 9204 1677 9820 1683
rect 2548 1657 2604 1663
rect 3236 1657 3468 1663
rect 5300 1657 7692 1663
rect 7700 1657 8460 1663
rect 8484 1657 8972 1663
rect 1764 1637 3324 1643
rect 3332 1637 3772 1643
rect 6308 1637 6572 1643
rect 7908 1637 9196 1643
rect 10340 1637 10924 1643
rect 10932 1637 11004 1643
rect 1428 1617 1916 1623
rect 1956 1617 2812 1623
rect 9652 1617 11692 1623
rect 52 1597 636 1603
rect 3028 1597 3628 1603
rect 7588 1597 7868 1603
rect 8372 1597 9180 1603
rect 9668 1597 9747 1603
rect 1300 1577 2412 1583
rect 2420 1577 3932 1583
rect 9044 1577 9724 1583
rect 9741 1583 9747 1597
rect 10388 1597 10492 1603
rect 9741 1577 10476 1583
rect 3188 1557 3420 1563
rect 3844 1557 7084 1563
rect 7092 1557 8124 1563
rect 8420 1557 9084 1563
rect 9748 1557 10380 1563
rect 564 1537 716 1543
rect 1220 1537 1356 1543
rect 1940 1537 2044 1543
rect 2052 1537 2828 1543
rect 3236 1537 5276 1543
rect 5284 1537 5420 1543
rect 7021 1537 7212 1543
rect 7021 1524 7027 1537
rect 2468 1517 2700 1523
rect 2740 1517 2748 1523
rect 3332 1517 3388 1523
rect 4004 1517 4012 1523
rect 4564 1517 4652 1523
rect 6388 1517 6396 1523
rect 6404 1517 6412 1523
rect 8228 1517 8316 1523
rect 9620 1517 9644 1523
rect 9668 1517 9708 1523
rect 10948 1517 10956 1523
rect 10964 1517 10988 1523
rect 11140 1517 11196 1523
rect 12109 1517 12220 1523
rect 1421 1503 1427 1516
rect 1284 1497 1836 1503
rect 1876 1497 1980 1503
rect 2189 1502 2316 1503
rect 2196 1497 2316 1502
rect 2340 1497 2620 1503
rect 4045 1503 4051 1516
rect 3828 1497 4051 1503
rect 4141 1502 4332 1503
rect 4148 1497 4332 1502
rect 7661 1503 7667 1516
rect 7661 1497 7756 1503
rect 9885 1503 9891 1516
rect 9204 1497 9891 1503
rect 11076 1497 11084 1503
rect 12109 1503 12115 1517
rect 11636 1497 12115 1503
rect 532 1477 604 1483
rect 612 1477 1436 1483
rect 1556 1477 1804 1483
rect 5780 1477 6364 1483
rect 11044 1477 11068 1483
rect 628 1457 1132 1463
rect 740 1437 1500 1443
rect 644 1417 796 1423
rect 3236 1417 3244 1423
rect 4340 1417 4572 1423
rect 5908 1417 5916 1423
rect 7012 1417 7068 1423
rect 7716 1417 8428 1423
rect 708 1397 716 1403
rect 1108 1397 1260 1403
rect 2004 1397 2860 1403
rect 4020 1397 4636 1403
rect 5428 1397 6972 1403
rect 7428 1397 8412 1403
rect 3812 1337 3932 1343
rect 5844 1337 5868 1343
rect 8036 1337 9340 1343
rect 9348 1337 9980 1343
rect 84 1318 236 1323
rect 244 1318 684 1323
rect 84 1317 684 1318
rect 1380 1317 1500 1323
rect 2340 1317 3084 1323
rect 3092 1318 4316 1323
rect 3092 1317 4323 1318
rect 5924 1317 5932 1323
rect 6436 1317 6572 1323
rect 6980 1317 7180 1323
rect 7396 1318 7404 1323
rect 7389 1317 7404 1318
rect 7732 1317 7836 1323
rect 9060 1317 9068 1323
rect 9172 1317 9324 1323
rect 9540 1317 10467 1323
rect 10644 1318 10652 1323
rect 10637 1317 10652 1318
rect 148 1297 172 1303
rect 804 1297 892 1303
rect 1444 1297 1564 1303
rect 2372 1297 2460 1303
rect 2580 1297 2652 1303
rect 2756 1297 2860 1303
rect 4324 1297 4412 1303
rect 5060 1297 5068 1303
rect 5140 1297 5164 1303
rect 5924 1297 5948 1303
rect 7300 1297 7308 1303
rect 7796 1297 7900 1303
rect 7940 1297 7948 1303
rect 8468 1297 8972 1303
rect 8980 1297 9196 1303
rect 9396 1297 9852 1303
rect 9892 1297 10028 1303
rect 10461 1303 10467 1317
rect 10980 1317 11084 1323
rect 11837 1304 11843 1316
rect 10461 1297 10540 1303
rect 11204 1297 11292 1303
rect 2436 1277 2508 1283
rect 2644 1277 2700 1283
rect 5828 1277 5836 1283
rect 6548 1277 6572 1283
rect 7780 1277 8524 1283
rect 11044 1277 11148 1283
rect 3780 1257 3820 1263
rect 5236 1257 5996 1263
rect 6532 1257 6604 1263
rect 8532 1257 9356 1263
rect 2548 1237 8716 1243
rect 1940 1217 5804 1223
rect 6532 1217 6572 1223
rect 148 1197 716 1203
rect 724 1197 908 1203
rect 916 1197 1532 1203
rect 9252 1197 9676 1203
rect 9732 1197 12860 1203
rect 4324 1177 4620 1183
rect 5060 1177 5276 1183
rect 7156 1177 7228 1183
rect 10964 1177 11660 1183
rect 1300 1157 1564 1163
rect 1572 1157 2748 1163
rect 2756 1157 2860 1163
rect 3252 1157 4140 1163
rect 7092 1157 7180 1163
rect 7892 1157 7932 1163
rect 11012 1157 11292 1163
rect 11300 1157 11628 1163
rect 1252 1137 1372 1143
rect 1844 1137 2044 1143
rect 2052 1137 2140 1143
rect 2436 1137 2540 1143
rect 2548 1137 2700 1143
rect 2708 1137 2796 1143
rect 4045 1137 4316 1143
rect 4045 1124 4051 1137
rect 5956 1137 6044 1143
rect 9060 1137 9100 1143
rect 9108 1137 9196 1143
rect 68 1117 76 1123
rect 356 1117 796 1123
rect 1444 1117 1548 1123
rect 1812 1117 1980 1123
rect 2100 1117 2220 1123
rect 3380 1117 3388 1123
rect 4932 1117 5068 1123
rect 5124 1117 5148 1123
rect 6532 1117 7020 1123
rect 7668 1117 7676 1123
rect 8308 1117 8316 1123
rect 8596 1117 8668 1123
rect 9252 1117 9356 1123
rect 9732 1117 10268 1123
rect 11172 1117 11180 1123
rect 11796 1117 12220 1123
rect 1549 1102 1564 1103
rect 1556 1097 1564 1102
rect 2564 1097 2636 1103
rect 3204 1097 3228 1103
rect 3236 1097 3276 1103
rect 3485 1102 4076 1103
rect 3492 1097 4076 1102
rect 5604 1102 5619 1103
rect 5604 1097 5612 1102
rect 7412 1102 7571 1103
rect 7412 1097 7564 1102
rect 8436 1097 8444 1103
rect 8468 1097 8476 1103
rect 9028 1097 9132 1103
rect 10436 1097 11084 1103
rect 5844 1077 5868 1083
rect 11044 1037 11132 1043
rect 468 1017 732 1023
rect 3972 1017 3980 1023
rect 3988 1017 3996 1023
rect 6468 1017 6476 1023
rect 2388 997 2572 1003
rect 3300 997 3308 1003
rect 3332 997 3340 1003
rect 3348 997 4044 1003
rect 10932 997 11132 1003
rect 7204 977 7660 983
rect 3940 957 6812 963
rect 7668 957 7884 963
rect 9796 957 9820 963
rect 10276 957 10428 963
rect 11684 957 11699 963
rect 244 937 252 943
rect 260 937 348 943
rect 5844 937 5868 943
rect 7796 937 8220 943
rect 8388 937 8684 943
rect 8692 937 8700 943
rect 11693 943 11699 957
rect 11693 937 11836 943
rect 1284 917 1292 923
rect 2020 917 2188 923
rect 2564 917 2636 923
rect 3636 918 4316 923
rect 3636 917 4323 918
rect 1197 904 1203 916
rect 3773 904 3779 917
rect 4532 917 4540 923
rect 6100 918 6108 923
rect 6093 917 6108 918
rect 8317 917 8428 923
rect 7085 904 7091 916
rect 8317 904 8323 917
rect 9028 917 9132 923
rect 10660 918 11468 923
rect 10660 917 11475 918
rect 11821 917 11884 923
rect 11821 904 11827 917
rect 84 897 124 903
rect 148 897 172 903
rect 180 897 892 903
rect 1444 897 1548 903
rect 1572 897 2092 903
rect 2100 897 2204 903
rect 2740 897 2748 903
rect 3812 897 3820 903
rect 4420 897 4428 903
rect 4532 897 4652 903
rect 5652 897 5740 903
rect 6004 897 6092 903
rect 6804 897 7020 903
rect 8516 897 8531 903
rect 8596 897 8716 903
rect 9828 897 9884 903
rect 10548 897 10556 903
rect 11556 897 11564 903
rect 1165 883 1171 896
rect 692 877 1171 883
rect 1380 877 1500 883
rect 2052 877 2140 883
rect 2708 877 2796 883
rect 4468 877 4620 883
rect 5956 877 6044 883
rect 9108 877 9196 883
rect 9700 877 9852 883
rect 10340 877 10476 883
rect 3796 857 5276 863
rect 10996 857 11772 863
rect 900 837 2556 843
rect 3844 837 3852 843
rect 628 817 1148 823
rect 6420 817 6428 823
rect 596 797 844 803
rect 852 797 1500 803
rect 7716 797 7772 803
rect 11700 797 11788 803
rect 644 777 876 783
rect 1956 777 3308 783
rect 9748 777 9868 783
rect 2548 757 2636 763
rect 7012 757 7900 763
rect 1908 737 2044 743
rect 2052 737 2140 743
rect 2637 743 2643 756
rect 2637 737 2700 743
rect 4564 737 4652 743
rect 5700 737 6588 743
rect 6596 737 7244 743
rect 9028 737 9036 743
rect 9780 737 10332 743
rect 10516 737 11100 743
rect 11108 737 11196 743
rect 804 717 908 723
rect 1444 717 1532 723
rect 2100 717 2172 723
rect 2756 717 2860 723
rect 4692 717 5212 723
rect 5668 717 5740 723
rect 5812 717 5996 723
rect 6004 717 6092 723
rect 7012 717 7020 723
rect 7117 717 7196 723
rect 765 704 771 716
rect 1421 703 1427 716
rect 884 702 899 703
rect 884 697 892 702
rect 1421 697 1500 703
rect 1844 697 1980 703
rect 2580 697 2588 703
rect 2596 697 2636 703
rect 3389 703 3395 716
rect 3188 697 3395 703
rect 3485 702 3532 703
rect 3492 697 3532 702
rect 4141 702 4364 703
rect 4148 697 4364 702
rect 4484 697 4588 703
rect 5876 697 6028 703
rect 6436 697 6524 703
rect 6548 697 6748 703
rect 7117 703 7123 717
rect 7300 717 7404 723
rect 10468 717 10476 723
rect 10532 717 10540 723
rect 10580 717 11196 723
rect 11204 717 11580 723
rect 12084 717 12220 723
rect 6756 697 7123 703
rect 9092 697 9132 703
rect 11636 697 11692 703
rect 148 677 668 683
rect 5844 677 5868 683
rect 11716 677 12236 683
rect 9677 644 9683 656
rect 2548 617 2572 623
rect 4628 617 4636 623
rect 5124 617 5132 623
rect 9092 617 9532 623
rect 3828 597 7132 603
rect 8324 597 8380 603
rect 4180 577 4524 583
rect 7236 577 9900 583
rect 12388 577 12476 583
rect 11636 557 12076 563
rect 6132 537 6492 543
rect 6500 537 7564 543
rect 8596 537 9116 543
rect 1533 526 1539 536
rect 212 518 236 523
rect 244 518 252 523
rect 212 517 252 518
rect 884 518 892 523
rect 884 517 899 518
rect 1069 517 1276 523
rect -51 497 76 503
rect 148 497 796 503
rect 1069 503 1075 517
rect 1533 517 1539 518
rect 2180 518 2188 523
rect 2180 517 2195 518
rect 2244 517 2620 523
rect 2749 517 2764 523
rect 2749 504 2755 517
rect 2852 518 2860 523
rect 2845 517 2860 518
rect 3828 517 3836 523
rect 3844 517 3923 523
rect 804 497 1075 503
rect 1300 497 1404 503
rect 2068 497 2076 503
rect 2100 497 2204 503
rect 2308 497 2684 503
rect 2692 497 2700 503
rect 2708 497 2716 503
rect 3917 503 3923 517
rect 5156 517 5164 523
rect 6084 518 6092 523
rect 6084 517 6099 518
rect 6621 517 6684 523
rect 6621 504 6627 517
rect 11076 517 11084 523
rect 11476 517 11580 523
rect 11668 517 11843 523
rect 11837 504 11843 517
rect 3917 497 3996 503
rect 4052 497 4172 503
rect 5860 497 5996 503
rect 6644 497 6748 503
rect 7652 497 7660 503
rect 8356 497 8364 503
rect 8413 497 8588 503
rect 84 477 156 483
rect 1437 483 1443 496
rect 1437 477 2028 483
rect 2868 477 4460 483
rect 5140 477 5276 483
rect 8413 483 8419 497
rect 8596 497 9084 503
rect 9156 497 9196 503
rect 9252 497 9660 503
rect 9764 497 9884 503
rect 10388 497 10476 503
rect 11204 497 11628 503
rect 7780 477 8419 483
rect 8436 477 9916 483
rect 9924 477 10476 483
rect 12036 477 12300 483
rect 596 457 748 463
rect 756 457 844 463
rect 4468 457 8220 463
rect 9012 457 9020 463
rect 9700 457 10540 463
rect 2708 437 4572 443
rect 5284 437 5980 443
rect 8372 437 9884 443
rect 9892 437 10428 443
rect 1892 417 2092 423
rect 4148 417 4620 423
rect 9060 417 9068 423
rect 5940 377 8364 383
rect 8596 377 9724 383
rect 10452 377 10556 383
rect 10964 377 11132 383
rect 644 357 764 363
rect 772 357 876 363
rect 7300 357 7868 363
rect 9076 357 9148 363
rect 11028 357 11068 363
rect 1412 337 1500 343
rect 4004 337 4524 343
rect 7396 337 9251 343
rect 1405 324 1411 336
rect 9245 324 9251 337
rect 11620 337 11676 343
rect 84 317 92 323
rect 148 317 156 323
rect 772 317 780 323
rect 804 317 892 323
rect 1444 317 1580 323
rect 2468 317 2476 323
rect 2724 317 2732 323
rect 2756 317 2876 323
rect 3780 317 3820 323
rect 4004 317 4012 323
rect 4580 317 5068 323
rect 5076 317 5932 323
rect 5956 317 5964 323
rect 6004 317 6044 323
rect 6628 317 6636 323
rect 7140 317 7292 323
rect 7796 317 7900 323
rect 8429 317 8524 323
rect 734 297 764 303
rect 893 302 1340 303
rect 900 297 1340 302
rect 2228 297 2636 303
rect 2948 297 3340 303
rect 5828 297 5836 303
rect 5934 297 5980 303
rect 6580 297 6588 303
rect 6756 297 7180 303
rect 7732 297 7836 303
rect 8429 303 8435 317
rect 9252 317 9996 323
rect 10004 317 10179 323
rect 8388 297 8435 303
rect 8452 297 8476 303
rect 10173 302 10179 317
rect 10276 317 10572 323
rect 10932 317 11004 323
rect 11476 317 11564 323
rect 11652 317 11804 323
rect 11844 317 12028 323
rect 788 277 1276 283
rect 1284 277 1308 283
rect 1972 277 2476 283
rect 2596 277 2620 283
rect 2868 277 3292 283
rect 4580 277 5964 283
rect 5988 277 6508 283
rect 3876 257 6636 263
rect 11700 257 11852 263
rect 4420 237 5276 243
rect 4580 217 4636 223
rect 9028 217 9148 223
rect 11572 217 11788 223
rect 612 197 684 203
rect 692 197 1036 203
rect 1284 197 1324 203
rect 3508 197 3884 203
rect 4516 197 4572 203
rect 11636 197 11644 203
rect 6548 177 6604 183
rect 1236 157 1388 163
rect 2852 157 5443 163
rect 5437 144 5443 157
rect 6532 157 6908 163
rect 6916 157 6924 163
rect 7140 157 8588 163
rect 3236 137 4956 143
rect 8436 137 10636 143
rect 10644 137 10652 143
rect 1860 117 1900 123
rect 2196 118 2332 123
rect 2189 117 2332 118
rect 2852 118 2940 123
rect 2845 117 2940 118
rect 4532 117 4572 123
rect 5156 117 5292 123
rect 5300 117 5347 123
rect 77 104 83 116
rect 1821 104 1827 116
rect 5341 104 5347 117
rect 5780 117 5948 123
rect 5965 117 6044 123
rect 5965 104 5971 117
rect 7732 117 7836 123
rect 8388 117 8524 123
rect 8932 117 9132 123
rect 9140 117 9212 123
rect 9860 117 9891 123
rect 9885 104 9891 117
rect 10404 117 10963 123
rect 148 97 204 103
rect 1044 97 1164 103
rect 1220 97 1228 103
rect 1844 97 1884 103
rect 2541 97 2748 103
rect 2541 84 2547 97
rect 3396 97 3500 103
rect 4468 97 4508 103
rect 4964 97 5068 103
rect 6932 97 7020 103
rect 9188 97 9196 103
rect 9252 97 9340 103
rect 9764 97 9852 103
rect 10548 97 10668 103
rect 10957 103 10963 117
rect 10980 117 11084 123
rect 10957 97 11196 103
rect 12212 97 12220 103
rect 12292 97 12924 103
rect 2708 77 2860 83
rect 3204 77 3324 83
rect 7012 77 7084 83
rect 7812 77 7900 83
rect 11060 77 11148 83
rect 1844 37 1852 43
rect 100 17 140 23
rect 772 17 780 23
rect 1812 17 1836 23
rect 2740 17 2748 23
rect 5972 17 5980 23
rect 6004 17 6012 23
<< m4contact >>
rect 6412 9016 6420 9024
rect 6444 9016 6452 9024
rect 10316 9016 10324 9024
rect 10348 9016 10356 9024
rect 3244 8976 3252 8984
rect 3180 8956 3188 8964
rect 6140 8956 6148 8964
rect 7772 8956 7780 8964
rect 8380 8956 8388 8964
rect 556 8936 564 8944
rect 1164 8936 1172 8944
rect 2508 8936 2516 8944
rect 1292 8916 1300 8924
rect 3244 8916 3252 8924
rect 3852 8916 3860 8924
rect 4140 8918 4148 8924
rect 4140 8916 4148 8918
rect 6604 8936 6612 8944
rect 7708 8936 7716 8944
rect 508 8896 516 8904
rect 556 8896 564 8904
rect 1164 8896 1172 8904
rect 1868 8896 1876 8904
rect 2364 8896 2372 8904
rect 2508 8896 2516 8904
rect 3020 8896 3028 8904
rect 3180 8896 3188 8904
rect 3788 8896 3796 8904
rect 4044 8896 4052 8904
rect 4652 8896 4660 8904
rect 5324 8896 5332 8904
rect 6140 8896 6148 8904
rect 7772 8916 7780 8924
rect 9340 8918 9348 8924
rect 9340 8916 9348 8918
rect 10636 8918 10644 8924
rect 10636 8916 10644 8918
rect 7708 8896 7716 8904
rect 8252 8896 8260 8904
rect 8380 8896 8388 8904
rect 8908 8896 8916 8904
rect 9900 8896 9908 8904
rect 11196 8896 11204 8904
rect 12220 8896 12228 8904
rect 1164 8876 1172 8884
rect 4092 8876 4100 8884
rect 4636 8876 4644 8884
rect 6748 8876 6756 8884
rect 9292 8876 9300 8884
rect 1420 8836 1428 8844
rect 1180 8756 1188 8764
rect 4956 8756 4964 8764
rect 5820 8756 5828 8764
rect 8044 8756 8052 8764
rect 10636 8756 10644 8764
rect 11292 8756 11300 8764
rect 7276 8736 7284 8744
rect 9292 8736 9300 8744
rect 9820 8736 9828 8744
rect 10876 8736 10884 8744
rect 524 8716 532 8724
rect 1180 8716 1188 8724
rect 1804 8716 1812 8724
rect 2460 8716 2468 8724
rect 2508 8716 2516 8724
rect 2732 8716 2740 8724
rect 3324 8716 3332 8724
rect 3388 8716 3396 8724
rect 1276 8696 1284 8704
rect 2668 8696 2676 8704
rect 2764 8702 2772 8704
rect 2764 8696 2772 8702
rect 5068 8716 5076 8724
rect 5132 8716 5140 8724
rect 5852 8716 5860 8724
rect 6908 8716 6916 8724
rect 7676 8716 7684 8724
rect 7948 8716 7956 8724
rect 8860 8716 8868 8724
rect 9612 8716 9620 8724
rect 10268 8716 10276 8724
rect 10860 8716 10868 8724
rect 11180 8716 11188 8724
rect 11820 8716 11828 8724
rect 3468 8702 3476 8704
rect 3468 8696 3476 8702
rect 5180 8696 5188 8704
rect 5820 8696 5828 8704
rect 6604 8696 6612 8704
rect 7404 8696 7412 8704
rect 7788 8696 7796 8704
rect 8044 8702 8052 8704
rect 8044 8696 8052 8702
rect 11004 8696 11012 8704
rect 11292 8702 11300 8704
rect 11292 8696 11300 8702
rect 11948 8702 11956 8704
rect 11948 8696 11956 8702
rect 1180 8676 1188 8684
rect 4636 8676 4644 8684
rect 6604 8676 6612 8684
rect 140 8656 148 8664
rect 1164 8656 1172 8664
rect 5852 8636 5860 8644
rect 1292 8616 1300 8624
rect 2668 8616 2676 8624
rect 6412 8616 6420 8624
rect 6444 8616 6452 8624
rect 10316 8616 10324 8624
rect 10348 8616 10356 8624
rect 11948 8616 11956 8624
rect 60 8596 68 8604
rect 524 8596 532 8604
rect 2508 8596 2516 8604
rect 5260 8596 5268 8604
rect 8396 8596 8404 8604
rect 8412 8596 8420 8604
rect 2460 8576 2468 8584
rect 8428 8576 8436 8584
rect 4492 8556 4500 8564
rect 7612 8556 7620 8564
rect 8380 8556 8388 8564
rect 11820 8556 11828 8564
rect 124 8536 132 8544
rect 1900 8516 1908 8524
rect 2188 8518 2196 8524
rect 2188 8516 2196 8518
rect 3468 8536 3476 8544
rect 6092 8536 6100 8544
rect 7132 8536 7140 8544
rect 7404 8536 7412 8544
rect 8412 8536 8420 8544
rect 3836 8516 3844 8524
rect 6028 8516 6036 8524
rect 8428 8516 8436 8524
rect 9052 8516 9060 8524
rect 10620 8516 10628 8524
rect 140 8496 148 8504
rect 1036 8496 1044 8504
rect 1708 8496 1716 8504
rect 3116 8496 3124 8504
rect 3372 8496 3380 8504
rect 4076 8496 4084 8504
rect 4956 8496 4964 8504
rect 5132 8496 5140 8504
rect 5836 8496 5844 8504
rect 5996 8496 6004 8504
rect 6700 8496 6708 8504
rect 7276 8496 7284 8504
rect 7404 8496 7412 8504
rect 8380 8496 8388 8504
rect 8844 8496 8852 8504
rect 9180 8496 9188 8504
rect 9260 8496 9268 8504
rect 9900 8496 9908 8504
rect 10700 8496 10708 8504
rect 11164 8496 11172 8504
rect 11788 8496 11796 8504
rect 636 8476 644 8484
rect 1116 8476 1124 8484
rect 1148 8476 1156 8484
rect 3324 8476 3332 8484
rect 5180 8476 5188 8484
rect 6012 8476 6020 8484
rect 8956 8476 8964 8484
rect 9788 8476 9796 8484
rect 9820 8476 9828 8484
rect 11804 8476 11812 8484
rect 8860 8456 8868 8464
rect 10876 8456 10884 8464
rect 4044 8436 4052 8444
rect 556 8416 564 8424
rect 7260 8416 7268 8424
rect 8252 8416 8260 8424
rect 11196 8396 11204 8404
rect 1276 8376 1284 8384
rect 7772 8376 7780 8384
rect 11004 8376 11012 8384
rect 620 8356 628 8364
rect 2524 8356 2532 8364
rect 10252 8356 10260 8364
rect 4412 8336 4420 8344
rect 7084 8336 7092 8344
rect 556 8316 564 8324
rect 1100 8316 1108 8324
rect 1692 8316 1700 8324
rect 2380 8316 2388 8324
rect 2508 8316 2516 8324
rect 2668 8316 2676 8324
rect 2732 8316 2740 8324
rect 2844 8316 2852 8324
rect 3836 8316 3844 8324
rect 4492 8316 4500 8324
rect 4716 8316 4724 8324
rect 5292 8316 5300 8324
rect 5980 8316 5988 8324
rect 6572 8316 6580 8324
rect 6588 8316 6596 8324
rect 6620 8316 6628 8324
rect 7660 8316 7668 8324
rect 7788 8316 7796 8324
rect 8220 8316 8228 8324
rect 8332 8316 8340 8324
rect 8524 8316 8532 8324
rect 8556 8316 8564 8324
rect 9324 8316 9332 8324
rect 10108 8316 10116 8324
rect 10668 8316 10676 8324
rect 11292 8316 11300 8324
rect 11644 8316 11652 8324
rect 620 8296 628 8304
rect 2572 8296 2580 8304
rect 2684 8296 2692 8304
rect 2764 8296 2772 8304
rect 4508 8296 4516 8304
rect 4780 8302 4788 8304
rect 4780 8296 4788 8302
rect 5132 8296 5140 8304
rect 5260 8296 5268 8304
rect 6620 8296 6628 8304
rect 7772 8296 7780 8304
rect 8428 8296 8436 8304
rect 10380 8296 10388 8304
rect 10396 8296 10404 8304
rect 7740 8276 7748 8284
rect 2572 8256 2580 8264
rect 8956 8256 8964 8264
rect 7948 8236 7956 8244
rect 9052 8236 9060 8244
rect 9996 8236 10004 8244
rect 8908 8216 8916 8224
rect 11788 8216 11796 8224
rect 1116 8196 1124 8204
rect 2508 8196 2516 8204
rect 5260 8196 5268 8204
rect 5292 8196 5300 8204
rect 11644 8196 11652 8204
rect 12284 8196 12292 8204
rect 12220 8176 12228 8184
rect 6428 8156 6436 8164
rect 12332 8156 12340 8164
rect 124 8136 132 8144
rect 2172 8136 2180 8144
rect 5756 8136 5764 8144
rect 8076 8136 8084 8144
rect 10652 8136 10660 8144
rect 1532 8118 1540 8124
rect 1532 8116 1540 8118
rect 2556 8116 2564 8124
rect 3484 8118 3492 8124
rect 3484 8116 3492 8118
rect 7612 8116 7620 8124
rect 7660 8116 7668 8124
rect 8588 8116 8596 8124
rect 9324 8116 9332 8124
rect 1164 8096 1172 8104
rect 1324 8096 1332 8104
rect 2172 8096 2180 8104
rect 3020 8096 3028 8104
rect 3276 8096 3284 8104
rect 4012 8096 4020 8104
rect 4748 8096 4756 8104
rect 5756 8096 5764 8104
rect 6284 8096 6292 8104
rect 6428 8096 6436 8104
rect 6940 8096 6948 8104
rect 7260 8096 7268 8104
rect 7276 8096 7284 8104
rect 7980 8096 7988 8104
rect 8684 8096 8692 8104
rect 9244 8096 9252 8104
rect 10524 8096 10532 8104
rect 11516 8096 11524 8104
rect 44 8076 52 8084
rect 3036 8076 3044 8084
rect 5388 8076 5396 8084
rect 8652 8076 8660 8084
rect 10284 8076 10292 8084
rect 10380 8076 10388 8084
rect 12204 8076 12212 8084
rect 2684 8056 2692 8064
rect 5100 8056 5108 8064
rect 8844 8036 8852 8044
rect 10636 8036 10644 8044
rect 10876 8036 10884 8044
rect 2668 8016 2676 8024
rect 2844 8016 2852 8024
rect 1292 7996 1300 8004
rect 6748 7996 6756 8004
rect 10252 7996 10260 8004
rect 2108 7976 2116 7984
rect 4604 7976 4612 7984
rect 10684 7976 10692 7984
rect 11292 7976 11300 7984
rect 1692 7956 1700 7964
rect 2204 7956 2212 7964
rect 2652 7956 2660 7964
rect 572 7936 580 7944
rect 3228 7936 3236 7944
rect 4028 7936 4036 7944
rect 6044 7936 6052 7944
rect 6604 7936 6612 7944
rect 8268 7936 8276 7944
rect 8396 7936 8404 7944
rect 9324 7936 9332 7944
rect 10876 7936 10884 7944
rect 540 7916 548 7924
rect 1164 7916 1172 7924
rect 1836 7916 1844 7924
rect 2012 7916 2020 7924
rect 2732 7916 2740 7924
rect 3996 7916 4004 7924
rect 4668 7916 4676 7924
rect 5292 7916 5300 7924
rect 6092 7916 6100 7924
rect 6748 7916 6756 7924
rect 7660 7916 7668 7924
rect 7884 7916 7892 7924
rect 7900 7916 7908 7924
rect 7948 7916 7956 7924
rect 8076 7916 8084 7924
rect 8908 7916 8916 7924
rect 9004 7916 9012 7924
rect 9228 7916 9236 7924
rect 9276 7916 9284 7924
rect 9996 7916 10004 7924
rect 10924 7916 10932 7924
rect 11308 7916 11316 7924
rect 12220 7916 12228 7924
rect 12284 7916 12292 7924
rect 620 7896 628 7904
rect 636 7896 644 7904
rect 1932 7896 1940 7904
rect 2204 7896 2212 7904
rect 3228 7896 3236 7904
rect 3820 7896 3828 7904
rect 4796 7902 4804 7904
rect 4796 7896 4804 7902
rect 5100 7896 5108 7904
rect 5452 7896 5460 7904
rect 3020 7876 3028 7884
rect 4156 7876 4164 7884
rect 7740 7896 7748 7904
rect 7804 7896 7812 7904
rect 9068 7896 9076 7904
rect 9324 7896 9332 7904
rect 9740 7896 9748 7904
rect 10988 7896 10996 7904
rect 11068 7896 11076 7904
rect 12332 7896 12340 7904
rect 6092 7876 6100 7884
rect 8060 7876 8068 7884
rect 11292 7876 11300 7884
rect 9068 7856 9076 7864
rect 10284 7856 10292 7864
rect 7052 7836 7060 7844
rect 7804 7836 7812 7844
rect 10924 7836 10932 7844
rect 4412 7816 4420 7824
rect 4508 7816 4516 7824
rect 4668 7816 4676 7824
rect 8396 7816 8404 7824
rect 9004 7816 9012 7824
rect 10860 7816 10868 7824
rect 76 7796 84 7804
rect 1100 7796 1108 7804
rect 4796 7796 4804 7804
rect 9612 7796 9620 7804
rect 9740 7796 9748 7804
rect 11644 7796 11652 7804
rect 11660 7796 11668 7804
rect 4140 7776 4148 7784
rect 1884 7756 1892 7764
rect 2108 7756 2116 7764
rect 5820 7756 5828 7764
rect 8428 7756 8436 7764
rect 11772 7756 11780 7764
rect 684 7736 692 7744
rect 6764 7736 6772 7744
rect 9980 7736 9988 7744
rect 9996 7736 10004 7744
rect 10652 7736 10660 7744
rect 4140 7718 4148 7724
rect 4140 7716 4148 7718
rect 6396 7716 6404 7724
rect 6764 7716 6772 7724
rect 7884 7716 7892 7724
rect 11644 7716 11652 7724
rect 460 7696 468 7704
rect 572 7696 580 7704
rect 732 7696 740 7704
rect 1756 7696 1764 7704
rect 1884 7696 1892 7704
rect 2460 7696 2468 7704
rect 3660 7696 3668 7704
rect 3772 7696 3780 7704
rect 3868 7696 3876 7704
rect 4044 7696 4052 7704
rect 4956 7696 4964 7704
rect 5116 7696 5124 7704
rect 5724 7696 5732 7704
rect 6364 7696 6372 7704
rect 6604 7696 6612 7704
rect 7292 7696 7300 7704
rect 8092 7696 8100 7704
rect 8572 7696 8580 7704
rect 9260 7696 9268 7704
rect 10220 7696 10228 7704
rect 10684 7696 10692 7704
rect 11564 7696 11572 7704
rect 11660 7696 11668 7704
rect 11740 7696 11748 7704
rect 6700 7676 6708 7684
rect 7692 7676 7700 7684
rect 2076 7656 2084 7664
rect 7292 7656 7300 7664
rect 11164 7656 11172 7664
rect 7516 7636 7524 7644
rect 8508 7636 8516 7644
rect 2476 7616 2484 7624
rect 6908 7596 6916 7604
rect 4012 7576 4020 7584
rect 4604 7576 4612 7584
rect 6460 7576 6468 7584
rect 2012 7556 2020 7564
rect 4684 7556 4692 7564
rect 7196 7556 7204 7564
rect 7964 7556 7972 7564
rect 2396 7536 2404 7544
rect 3052 7536 3060 7544
rect 4780 7536 4788 7544
rect 4796 7536 4804 7544
rect 6060 7536 6068 7544
rect 9964 7536 9972 7544
rect 748 7516 756 7524
rect 812 7516 820 7524
rect 1436 7516 1444 7524
rect 2460 7516 2468 7524
rect 3228 7516 3236 7524
rect 3340 7516 3348 7524
rect 3532 7516 3540 7524
rect 3932 7516 3940 7524
rect 4044 7516 4052 7524
rect 4684 7516 4692 7524
rect 6460 7516 6468 7524
rect 7036 7516 7044 7524
rect 7932 7516 7940 7524
rect 8828 7516 8836 7524
rect 8988 7516 8996 7524
rect 9340 7516 9348 7524
rect 9852 7516 9860 7524
rect 10716 7516 10724 7524
rect 11116 7516 11124 7524
rect 11148 7516 11156 7524
rect 11196 7516 11204 7524
rect 11772 7516 11780 7524
rect 92 7496 100 7504
rect 108 7496 116 7504
rect 700 7496 708 7504
rect 1900 7496 1908 7504
rect 2588 7496 2596 7504
rect 2828 7502 2836 7504
rect 2828 7496 2836 7502
rect 3116 7496 3124 7504
rect 3164 7496 3172 7504
rect 4060 7502 4068 7504
rect 4060 7496 4068 7502
rect 4796 7502 4804 7504
rect 4796 7496 4804 7502
rect 5388 7496 5396 7504
rect 6076 7496 6084 7504
rect 7148 7496 7156 7504
rect 7756 7496 7764 7504
rect 7916 7496 7924 7504
rect 9036 7496 9044 7504
rect 9356 7496 9364 7504
rect 9724 7496 9732 7504
rect 9964 7496 9972 7504
rect 9980 7502 9988 7504
rect 9980 7496 9988 7502
rect 10412 7496 10420 7504
rect 11100 7496 11108 7504
rect 124 7476 132 7484
rect 3820 7476 3828 7484
rect 3996 7476 4004 7484
rect 8684 7476 8692 7484
rect 8700 7476 8708 7484
rect 11180 7456 11188 7464
rect 1148 7436 1156 7444
rect 4044 7436 4052 7444
rect 7036 7416 7044 7424
rect 9228 7416 9236 7424
rect 12204 7416 12212 7424
rect 700 7396 708 7404
rect 748 7396 756 7404
rect 2460 7396 2468 7404
rect 6412 7396 6420 7404
rect 6460 7396 6468 7404
rect 6940 7396 6948 7404
rect 9356 7396 9364 7404
rect 10348 7396 10356 7404
rect 11100 7396 11108 7404
rect 11148 7396 11156 7404
rect 1292 7376 1300 7384
rect 9212 7376 9220 7384
rect 9244 7376 9252 7384
rect 1228 7356 1236 7364
rect 6060 7356 6068 7364
rect 10492 7356 10500 7364
rect 1436 7336 1444 7344
rect 8444 7336 8452 7344
rect 1292 7316 1300 7324
rect 2556 7316 2564 7324
rect 2604 7316 2612 7324
rect 3500 7316 3508 7324
rect 6076 7316 6084 7324
rect 6460 7316 6468 7324
rect 6764 7316 6772 7324
rect 8028 7318 8036 7324
rect 8028 7316 8036 7318
rect 9228 7316 9236 7324
rect 9324 7316 9332 7324
rect 11916 7316 11924 7324
rect 444 7296 452 7304
rect 1164 7296 1172 7304
rect 1228 7296 1236 7304
rect 1660 7296 1668 7304
rect 2476 7296 2484 7304
rect 2492 7296 2500 7304
rect 3116 7296 3124 7304
rect 3164 7296 3172 7304
rect 3212 7296 3220 7304
rect 3996 7296 4004 7304
rect 4220 7296 4228 7304
rect 5724 7296 5732 7304
rect 6268 7296 6276 7304
rect 6412 7296 6420 7304
rect 6604 7296 6612 7304
rect 6652 7296 6660 7304
rect 7516 7296 7524 7304
rect 7916 7296 7924 7304
rect 9212 7296 9220 7304
rect 9372 7296 9380 7304
rect 10124 7296 10132 7304
rect 10348 7296 10356 7304
rect 10556 7296 10564 7304
rect 11740 7296 11748 7304
rect 11788 7296 11796 7304
rect 11852 7296 11860 7304
rect 812 7276 820 7284
rect 3036 7276 3044 7284
rect 10348 7276 10356 7284
rect 4092 7256 4100 7264
rect 8556 7256 8564 7264
rect 10908 7236 10916 7244
rect 4588 7216 4596 7224
rect 3996 7196 4004 7204
rect 8028 7196 8036 7204
rect 8412 7196 8420 7204
rect 9372 7156 9380 7164
rect 172 7136 180 7144
rect 3644 7136 3652 7144
rect 7692 7136 7700 7144
rect 10332 7136 10340 7144
rect 76 7116 84 7124
rect 1068 7116 1076 7124
rect 1388 7116 1396 7124
rect 1836 7116 1844 7124
rect 2124 7116 2132 7124
rect 3644 7116 3652 7124
rect 3788 7116 3796 7124
rect 3868 7116 3876 7124
rect 204 7102 212 7104
rect 204 7096 212 7102
rect 2556 7096 2564 7104
rect 3020 7102 3028 7104
rect 3020 7096 3028 7102
rect 3868 7096 3876 7104
rect 124 7076 132 7084
rect 4412 7116 4420 7124
rect 5084 7116 5092 7124
rect 5244 7116 5252 7124
rect 5788 7116 5796 7124
rect 6572 7116 6580 7124
rect 6988 7116 6996 7124
rect 7084 7116 7092 7124
rect 7292 7116 7300 7124
rect 8332 7116 8340 7124
rect 8732 7116 8740 7124
rect 9356 7116 9364 7124
rect 10636 7116 10644 7124
rect 11116 7116 11124 7124
rect 4508 7096 4516 7104
rect 5388 7102 5396 7104
rect 5388 7096 5396 7102
rect 6604 7096 6612 7104
rect 7116 7096 7124 7104
rect 7132 7096 7140 7104
rect 8444 7096 8452 7104
rect 8668 7102 8676 7104
rect 8668 7096 8676 7102
rect 11564 7096 11572 7104
rect 4076 7076 4084 7084
rect 11788 7056 11796 7064
rect 1388 7036 1396 7044
rect 5788 7036 5796 7044
rect 716 7016 724 7024
rect 2204 7016 2212 7024
rect 3388 7016 3396 7024
rect 12220 7016 12228 7024
rect 2140 6996 2148 7004
rect 5084 6996 5092 7004
rect 9388 6996 9396 7004
rect 12300 6996 12308 7004
rect 12316 6996 12324 7004
rect 7980 6976 7988 6984
rect 12332 6956 12340 6964
rect 1868 6916 1876 6924
rect 6732 6936 6740 6944
rect 8668 6936 8676 6944
rect 9356 6936 9364 6944
rect 2204 6916 2212 6924
rect 5356 6916 5364 6924
rect 5836 6916 5844 6924
rect 6732 6918 6740 6924
rect 6732 6916 6740 6918
rect 8508 6916 8516 6924
rect 8748 6916 8756 6924
rect 9980 6918 9988 6924
rect 9980 6916 9988 6918
rect 10316 6916 10324 6924
rect 10636 6918 10644 6924
rect 10636 6916 10644 6918
rect 540 6896 548 6904
rect 1148 6896 1156 6904
rect 1708 6896 1716 6904
rect 2204 6896 2212 6904
rect 2748 6896 2756 6904
rect 3388 6896 3396 6904
rect 4332 6896 4340 6904
rect 4828 6896 4836 6904
rect 5340 6896 5348 6904
rect 5452 6896 5460 6904
rect 5836 6896 5844 6904
rect 6668 6896 6676 6904
rect 7388 6896 7396 6904
rect 8316 6896 8324 6904
rect 8604 6896 8612 6904
rect 9372 6896 9380 6904
rect 9852 6896 9860 6904
rect 1612 6876 1620 6884
rect 1740 6876 1748 6884
rect 1916 6876 1924 6884
rect 2140 6876 2148 6884
rect 4364 6876 4372 6884
rect 5404 6876 5412 6884
rect 9836 6876 9844 6884
rect 10140 6896 10148 6904
rect 11196 6896 11204 6904
rect 12156 6896 12164 6904
rect 10748 6876 10756 6884
rect 6604 6836 6612 6844
rect 7372 6836 7380 6844
rect 444 6816 452 6824
rect 10268 6816 10276 6824
rect 11916 6816 11924 6824
rect 2204 6796 2212 6804
rect 7388 6796 7396 6804
rect 8316 6796 8324 6804
rect 4364 6776 4372 6784
rect 636 6756 644 6764
rect 4044 6756 4052 6764
rect 4780 6756 4788 6764
rect 11516 6756 11524 6764
rect 11660 6756 11668 6764
rect 92 6736 100 6744
rect 12300 6736 12308 6744
rect 76 6716 84 6724
rect 380 6716 388 6724
rect 1180 6716 1188 6724
rect 1436 6716 1444 6724
rect 2044 6716 2052 6724
rect 2716 6716 2724 6724
rect 2844 6716 2852 6724
rect 3388 6716 3396 6724
rect 4044 6716 4052 6724
rect 4332 6716 4340 6724
rect 4364 6716 4372 6724
rect 4732 6716 4740 6724
rect 5500 6716 5508 6724
rect 6300 6716 6308 6724
rect 7004 6716 7012 6724
rect 7292 6716 7300 6724
rect 7388 6716 7396 6724
rect 8060 6716 8068 6724
rect 8508 6716 8516 6724
rect 8700 6716 8708 6724
rect 9356 6716 9364 6724
rect 10540 6716 10548 6724
rect 10748 6716 10756 6724
rect 12220 6716 12228 6724
rect 12332 6716 12340 6724
rect 12476 6716 12484 6724
rect 156 6702 164 6704
rect 156 6696 164 6702
rect 1276 6696 1284 6704
rect 2636 6696 2644 6704
rect 2812 6702 2820 6704
rect 2812 6696 2820 6702
rect 2828 6696 2836 6704
rect 4668 6696 4676 6704
rect 7132 6696 7140 6704
rect 8460 6696 8468 6704
rect 9836 6696 9844 6704
rect 10172 6696 10180 6704
rect 10636 6696 10644 6704
rect 124 6676 132 6684
rect 12332 6696 12340 6704
rect 2844 6676 2852 6684
rect 3660 6676 3668 6684
rect 5420 6676 5428 6684
rect 9740 6676 9748 6684
rect 10364 6676 10372 6684
rect 2844 6656 2852 6664
rect 1772 6616 1780 6624
rect 10012 6616 10020 6624
rect 748 6596 756 6604
rect 2044 6596 2052 6604
rect 4364 6596 4372 6604
rect 11644 6596 11652 6604
rect 1292 6576 1300 6584
rect 10380 6576 10388 6584
rect 1244 6556 1252 6564
rect 7772 6556 7780 6564
rect 9052 6556 9060 6564
rect 11468 6556 11476 6564
rect 124 6536 132 6544
rect 6428 6536 6436 6544
rect 6588 6536 6596 6544
rect 7708 6536 7716 6544
rect 8668 6536 8676 6544
rect 9340 6536 9348 6544
rect 10956 6536 10964 6544
rect 76 6516 84 6524
rect 156 6516 164 6524
rect 1292 6516 1300 6524
rect 1868 6516 1876 6524
rect 5260 6516 5268 6524
rect 5420 6516 5428 6524
rect 6700 6516 6708 6524
rect 7772 6516 7780 6524
rect 8220 6518 8228 6524
rect 8220 6516 8228 6518
rect 9740 6516 9748 6524
rect 10332 6516 10340 6524
rect 11196 6516 11204 6524
rect 11660 6516 11668 6524
rect 92 6496 100 6504
rect 1180 6496 1188 6504
rect 1244 6496 1252 6504
rect 1804 6496 1812 6504
rect 2412 6496 2420 6504
rect 2524 6496 2532 6504
rect 3420 6496 3428 6504
rect 4044 6496 4052 6504
rect 5340 6496 5348 6504
rect 6108 6496 6116 6504
rect 6620 6496 6628 6504
rect 6636 6496 6644 6504
rect 6780 6496 6788 6504
rect 7708 6496 7716 6504
rect 8348 6496 8356 6504
rect 8828 6496 8836 6504
rect 8860 6496 8868 6504
rect 9052 6496 9060 6504
rect 9532 6496 9540 6504
rect 10156 6496 10164 6504
rect 10316 6496 10324 6504
rect 10924 6496 10932 6504
rect 10956 6496 10964 6504
rect 11468 6496 11476 6504
rect 11644 6496 11652 6504
rect 11820 6496 11828 6504
rect 1740 6476 1748 6484
rect 1932 6476 1940 6484
rect 2364 6476 2372 6484
rect 5020 6476 5028 6484
rect 6044 6476 6052 6484
rect 6700 6476 6708 6484
rect 9852 6476 9860 6484
rect 11804 6476 11812 6484
rect 4044 6456 4052 6464
rect 524 6436 532 6444
rect 2380 6436 2388 6444
rect 1180 6416 1188 6424
rect 156 6396 164 6404
rect 604 6396 612 6404
rect 1916 6396 1924 6404
rect 2188 6396 2196 6404
rect 3244 6396 3252 6404
rect 4940 6396 4948 6404
rect 6412 6396 6420 6404
rect 6460 6396 6468 6404
rect 7020 6396 7028 6404
rect 6428 6376 6436 6384
rect 5020 6356 5028 6364
rect 6476 6356 6484 6364
rect 7004 6356 7012 6364
rect 8060 6356 8068 6364
rect 8316 6356 8324 6364
rect 1132 6336 1140 6344
rect 3132 6336 3140 6344
rect 5020 6336 5028 6344
rect 7356 6336 7364 6344
rect 8476 6336 8484 6344
rect 524 6316 532 6324
rect 748 6316 756 6324
rect 2012 6316 2020 6324
rect 2076 6316 2084 6324
rect 2124 6316 2132 6324
rect 3164 6316 3172 6324
rect 3676 6316 3684 6324
rect 3804 6316 3812 6324
rect 1292 6296 1300 6304
rect 3004 6276 3012 6284
rect 9532 6336 9540 6344
rect 4044 6316 4052 6324
rect 4780 6316 4788 6324
rect 4956 6316 4964 6324
rect 5292 6316 5300 6324
rect 5468 6316 5476 6324
rect 6012 6316 6020 6324
rect 7020 6316 7028 6324
rect 7068 6316 7076 6324
rect 7580 6316 7588 6324
rect 8300 6316 8308 6324
rect 8316 6316 8324 6324
rect 9868 6316 9876 6324
rect 11212 6316 11220 6324
rect 11916 6316 11924 6324
rect 12284 6316 12292 6324
rect 5180 6296 5188 6304
rect 5260 6296 5268 6304
rect 7100 6296 7108 6304
rect 7372 6296 7380 6304
rect 8556 6296 8564 6304
rect 9052 6296 9060 6304
rect 9356 6296 9364 6304
rect 9724 6296 9732 6304
rect 12300 6296 12308 6304
rect 2060 6216 2068 6224
rect 3148 6216 3156 6224
rect 3804 6216 3812 6224
rect 380 6196 388 6204
rect 2508 6196 2516 6204
rect 3116 6196 3124 6204
rect 5068 6216 5076 6224
rect 5260 6216 5268 6224
rect 5292 6216 5300 6224
rect 5308 6216 5316 6224
rect 7068 6216 7076 6224
rect 11852 6216 11860 6224
rect 6300 6196 6308 6204
rect 8364 6196 8372 6204
rect 1932 6176 1940 6184
rect 2492 6176 2500 6184
rect 7100 6176 7108 6184
rect 8428 6176 8436 6184
rect 9724 6176 9732 6184
rect 732 6156 740 6164
rect 1884 6156 1892 6164
rect 2604 6156 2612 6164
rect 5756 6156 5764 6164
rect 5948 6156 5956 6164
rect 7276 6156 7284 6164
rect 9276 6156 9284 6164
rect 556 6136 564 6144
rect 1900 6136 1908 6144
rect 2556 6136 2564 6144
rect 6764 6136 6772 6144
rect 1932 6116 1940 6124
rect 2556 6116 2564 6124
rect 2636 6116 2644 6124
rect 2972 6116 2980 6124
rect 3372 6116 3380 6124
rect 3484 6118 3492 6124
rect 3484 6116 3492 6118
rect 4012 6116 4020 6124
rect 6460 6116 6468 6124
rect 6572 6116 6580 6124
rect 7644 6116 7652 6124
rect 7788 6116 7796 6124
rect 8428 6116 8436 6124
rect 8588 6116 8596 6124
rect 9724 6116 9732 6124
rect 10380 6116 10388 6124
rect 10636 6118 10644 6124
rect 10636 6116 10644 6118
rect 428 6096 436 6104
rect 556 6096 564 6104
rect 1084 6096 1092 6104
rect 1884 6096 1892 6104
rect 2364 6096 2372 6104
rect 3116 6096 3124 6104
rect 3148 6096 3156 6104
rect 3388 6096 3396 6104
rect 4124 6096 4132 6104
rect 5756 6096 5764 6104
rect 6364 6096 6372 6104
rect 6412 6096 6420 6104
rect 6508 6096 6516 6104
rect 6684 6096 6692 6104
rect 7692 6096 7700 6104
rect 8252 6096 8260 6104
rect 8364 6096 8372 6104
rect 9612 6096 9620 6104
rect 9788 6096 9796 6104
rect 10508 6096 10516 6104
rect 10524 6096 10532 6104
rect 11180 6096 11188 6104
rect 11804 6096 11812 6104
rect 972 6076 980 6084
rect 2572 6076 2580 6084
rect 6060 6076 6068 6084
rect 204 6056 212 6064
rect 3836 6056 3844 6064
rect 4732 6056 4740 6064
rect 6476 6056 6484 6064
rect 7804 6056 7812 6064
rect 8476 6056 8484 6064
rect 11180 6056 11188 6064
rect 2188 6036 2196 6044
rect 2508 6036 2516 6044
rect 2972 6036 2980 6044
rect 172 6016 180 6024
rect 9900 6016 9908 6024
rect 2876 5956 2884 5964
rect 11804 5956 11812 5964
rect 492 5936 500 5944
rect 3884 5936 3892 5944
rect 444 5916 452 5924
rect 748 5916 756 5924
rect 972 5916 980 5924
rect 1692 5916 1700 5924
rect 2060 5916 2068 5924
rect 2108 5916 2116 5924
rect 2732 5916 2740 5924
rect 2876 5916 2884 5924
rect 3836 5916 3844 5924
rect 3884 5916 3892 5924
rect 3948 5916 3956 5924
rect 5052 5916 5060 5924
rect 5084 5916 5092 5924
rect 5308 5916 5316 5924
rect 5340 5916 5348 5924
rect 6604 5916 6612 5924
rect 6796 5916 6804 5924
rect 7452 5916 7460 5924
rect 7836 5936 7844 5944
rect 8972 5916 8980 5924
rect 9852 5916 9860 5924
rect 9900 5916 9908 5924
rect 10156 5916 10164 5924
rect 10380 5916 10388 5924
rect 10524 5916 10532 5924
rect 10540 5916 10548 5924
rect 10668 5916 10676 5924
rect 11132 5916 11140 5924
rect 604 5896 612 5904
rect 732 5896 734 5904
rect 734 5896 740 5904
rect 1676 5896 1684 5904
rect 1708 5896 1716 5904
rect 1932 5896 1940 5904
rect 2188 5902 2196 5904
rect 2188 5896 2196 5902
rect 2764 5902 2772 5904
rect 2764 5896 2772 5902
rect 3420 5896 3428 5904
rect 3852 5896 3860 5904
rect 5196 5896 5204 5904
rect 5948 5896 5956 5904
rect 6092 5902 6100 5904
rect 6092 5896 6100 5902
rect 7900 5896 7908 5904
rect 8316 5896 8324 5904
rect 9708 5896 9716 5904
rect 9724 5896 9732 5904
rect 9980 5902 9988 5904
rect 9980 5896 9988 5902
rect 10636 5902 10644 5904
rect 10636 5896 10644 5902
rect 9356 5876 9364 5884
rect 11260 5876 11268 5884
rect 8556 5856 8564 5864
rect 1132 5836 1140 5844
rect 6092 5836 6100 5844
rect 6908 5836 6916 5844
rect 748 5816 756 5824
rect 1292 5816 1300 5824
rect 6604 5816 6612 5824
rect 12220 5816 12228 5824
rect 732 5796 740 5804
rect 4492 5796 4500 5804
rect 12284 5796 12292 5804
rect 12300 5796 12308 5804
rect 5324 5776 5332 5784
rect 10348 5776 10356 5784
rect 2460 5756 2468 5764
rect 4412 5756 4420 5764
rect 5148 5756 5156 5764
rect 5276 5756 5284 5764
rect 7100 5756 7108 5764
rect 10348 5756 10356 5764
rect 1964 5716 1972 5724
rect 2604 5716 2612 5724
rect 3004 5716 3012 5724
rect 7116 5736 7124 5744
rect 8556 5736 8564 5744
rect 4524 5716 4532 5724
rect 5148 5716 5156 5724
rect 5804 5716 5812 5724
rect 9324 5716 9332 5724
rect 10652 5716 10660 5724
rect 12300 5716 12308 5724
rect 60 5696 68 5704
rect 1100 5696 1108 5704
rect 1836 5696 1844 5704
rect 1900 5696 1908 5704
rect 2188 5696 2196 5704
rect 2460 5696 2468 5704
rect 2492 5696 2500 5704
rect 3020 5696 3028 5704
rect 3132 5696 3140 5704
rect 4412 5696 4420 5704
rect 4492 5696 4500 5704
rect 5468 5696 5476 5704
rect 5484 5696 5492 5704
rect 5996 5696 6004 5704
rect 6956 5696 6964 5704
rect 7100 5696 7108 5704
rect 7660 5696 7668 5704
rect 7948 5696 7956 5704
rect 8028 5696 8036 5704
rect 8604 5696 8612 5704
rect 9244 5696 9252 5704
rect 9900 5696 9908 5704
rect 10444 5696 10452 5704
rect 10748 5696 10756 5704
rect 4092 5676 4100 5684
rect 4796 5676 4804 5684
rect 6060 5676 6068 5684
rect 7036 5676 7044 5684
rect 8012 5676 8020 5684
rect 12220 5696 12228 5704
rect 12284 5696 12292 5704
rect 460 5656 468 5664
rect 4412 5656 4420 5664
rect 492 5636 500 5644
rect 3948 5636 3956 5644
rect 7084 5636 7092 5644
rect 604 5616 612 5624
rect 1084 5596 1092 5604
rect 2764 5596 2772 5604
rect 4652 5596 4660 5604
rect 5164 5596 5172 5604
rect 9068 5596 9076 5604
rect 10924 5576 10932 5584
rect 2732 5556 2740 5564
rect 4428 5556 4436 5564
rect 7836 5556 7844 5564
rect 9020 5556 9028 5564
rect 10396 5556 10404 5564
rect 732 5536 740 5544
rect 2876 5536 2884 5544
rect 3052 5536 3060 5544
rect 3500 5536 3508 5544
rect 4652 5536 4660 5544
rect 5292 5536 5300 5544
rect 6700 5536 6708 5544
rect 8012 5536 8020 5544
rect 10508 5536 10516 5544
rect 11756 5536 11764 5544
rect 524 5516 532 5524
rect 556 5516 564 5524
rect 1132 5516 1140 5524
rect 1708 5516 1716 5524
rect 2348 5516 2356 5524
rect 2556 5516 2564 5524
rect 3004 5516 3012 5524
rect 3772 5516 3780 5524
rect 3788 5516 3796 5524
rect 3948 5516 3956 5524
rect 4012 5516 4020 5524
rect 5660 5516 5668 5524
rect 6380 5516 6388 5524
rect 6412 5516 6420 5524
rect 6908 5516 6916 5524
rect 7660 5516 7668 5524
rect 7804 5516 7812 5524
rect 7948 5516 7956 5524
rect 8316 5516 8324 5524
rect 8700 5516 8708 5524
rect 8860 5516 8868 5524
rect 9228 5516 9236 5524
rect 10156 5516 10164 5524
rect 10332 5516 10340 5524
rect 10524 5516 10532 5524
rect 11612 5516 11620 5524
rect 11772 5516 11780 5524
rect 12316 5516 12324 5524
rect 604 5496 612 5504
rect 700 5496 708 5504
rect 1948 5496 1956 5504
rect 3212 5496 3220 5504
rect 3244 5496 3252 5504
rect 4572 5496 4580 5504
rect 5820 5496 5828 5504
rect 6476 5496 6484 5504
rect 7516 5496 7524 5504
rect 7820 5496 7828 5504
rect 8828 5496 8836 5504
rect 9356 5496 9364 5504
rect 10396 5496 10404 5504
rect 11292 5496 11300 5504
rect 11836 5496 11844 5504
rect 11868 5502 11876 5504
rect 11868 5496 11876 5502
rect 2572 5476 2580 5484
rect 3260 5476 3268 5484
rect 8428 5476 8436 5484
rect 604 5456 612 5464
rect 1100 5456 1108 5464
rect 6476 5456 6484 5464
rect 10108 5456 10116 5464
rect 5660 5436 5668 5444
rect 6284 5436 6292 5444
rect 8268 5436 8276 5444
rect 556 5416 564 5424
rect 3676 5416 3684 5424
rect 5820 5416 5828 5424
rect 6076 5416 6084 5424
rect 6412 5416 6420 5424
rect 140 5396 148 5404
rect 1724 5396 1732 5404
rect 6316 5396 6324 5404
rect 9644 5396 9652 5404
rect 11132 5396 11140 5404
rect 1164 5376 1172 5384
rect 4828 5376 4836 5384
rect 8988 5376 8996 5384
rect 3324 5356 3332 5364
rect 3388 5356 3396 5364
rect 9676 5356 9684 5364
rect 11708 5356 11716 5364
rect 6780 5336 6788 5344
rect 7756 5336 7764 5344
rect 10396 5336 10404 5344
rect 10972 5336 10980 5344
rect 1276 5316 1284 5324
rect 1740 5316 1748 5324
rect 1900 5316 1908 5324
rect 2076 5316 2084 5324
rect 2764 5316 2772 5324
rect 3644 5316 3652 5324
rect 3980 5316 3988 5324
rect 4508 5316 4516 5324
rect 4780 5318 4788 5324
rect 4780 5316 4788 5318
rect 5436 5318 5444 5324
rect 5436 5316 5444 5318
rect 6076 5316 6084 5324
rect 7004 5316 7012 5324
rect 7228 5316 7236 5324
rect 8428 5316 8436 5324
rect 9068 5316 9076 5324
rect 9180 5316 9188 5324
rect 10364 5316 10372 5324
rect 11708 5316 11716 5324
rect 76 5296 84 5304
rect 140 5296 148 5304
rect 748 5296 756 5304
rect 1836 5296 1844 5304
rect 2332 5296 2340 5304
rect 2476 5296 2484 5304
rect 2732 5296 2740 5304
rect 2812 5296 2820 5304
rect 3820 5296 3828 5304
rect 3948 5296 3956 5304
rect 4044 5296 4052 5304
rect 4668 5296 4676 5304
rect 4684 5296 4692 5304
rect 6140 5296 6148 5304
rect 7036 5296 7044 5304
rect 7420 5296 7428 5304
rect 204 5276 212 5284
rect 1868 5276 1876 5284
rect 3212 5276 3220 5284
rect 3548 5276 3556 5284
rect 6412 5276 6420 5284
rect 8972 5296 8980 5304
rect 9020 5296 9028 5304
rect 9644 5296 9652 5304
rect 9676 5296 9684 5304
rect 10220 5296 10228 5304
rect 10268 5296 10276 5304
rect 10524 5296 10532 5304
rect 11804 5296 11812 5304
rect 11852 5296 11860 5304
rect 12604 5296 12612 5304
rect 8268 5276 8276 5284
rect 700 5256 708 5264
rect 2460 5256 2468 5264
rect 8972 5256 8980 5264
rect 12220 5256 12228 5264
rect 4668 5236 4676 5244
rect 5100 5236 5108 5244
rect 5452 5236 5460 5244
rect 5820 5236 5828 5244
rect 9788 5236 9796 5244
rect 732 5216 740 5224
rect 2076 5216 2084 5224
rect 748 5196 756 5204
rect 2332 5196 2340 5204
rect 2860 5196 2868 5204
rect 3324 5196 3332 5204
rect 4412 5196 4420 5204
rect 5804 5196 5812 5204
rect 7068 5196 7076 5204
rect 8076 5196 8084 5204
rect 9004 5196 9012 5204
rect 4220 5176 4228 5184
rect 4524 5176 4532 5184
rect 5804 5176 5812 5184
rect 5836 5176 5844 5184
rect 7116 5176 7124 5184
rect 7676 5176 7684 5184
rect 8860 5176 8868 5184
rect 412 5156 420 5164
rect 1708 5156 1716 5164
rect 4124 5156 4132 5164
rect 7948 5156 7956 5164
rect 4684 5136 4692 5144
rect 10172 5136 10180 5144
rect 204 5116 212 5124
rect 1180 5116 1188 5124
rect 1212 5116 1220 5124
rect 1836 5116 1844 5124
rect 2332 5116 2340 5124
rect 3068 5116 3076 5124
rect 3388 5116 3396 5124
rect 5020 5116 5028 5124
rect 5164 5116 5172 5124
rect 5324 5116 5332 5124
rect 5340 5116 5348 5124
rect 5372 5116 5380 5124
rect 6444 5116 6452 5124
rect 6604 5116 6612 5124
rect 6780 5116 6788 5124
rect 7388 5116 7396 5124
rect 7964 5116 7972 5124
rect 8876 5116 8884 5124
rect 9004 5116 9012 5124
rect 10140 5116 10148 5124
rect 10540 5116 10548 5124
rect 10684 5116 10692 5124
rect 12284 5116 12292 5124
rect 1292 5096 1300 5104
rect 1900 5096 1908 5104
rect 2572 5096 2580 5104
rect 3996 5096 4004 5104
rect 4620 5096 4628 5104
rect 4796 5102 4804 5104
rect 4796 5096 4804 5102
rect 5804 5096 5812 5104
rect 5852 5096 5860 5104
rect 6460 5096 6468 5104
rect 6748 5096 6756 5104
rect 9708 5096 9716 5104
rect 10508 5096 10516 5104
rect 11132 5096 11134 5104
rect 11134 5096 11140 5104
rect 12348 5096 12356 5104
rect 10572 5076 10580 5084
rect 4684 5056 4692 5064
rect 4044 5016 4052 5024
rect 4620 5016 4628 5024
rect 7740 5016 7748 5024
rect 1820 4996 1828 5004
rect 3820 4996 3828 5004
rect 7644 4996 7652 5004
rect 7724 4996 7732 5004
rect 8524 4996 8532 5004
rect 12972 4996 12980 5004
rect 508 4976 516 4984
rect 1196 4976 1204 4984
rect 8572 4976 8580 4984
rect 12284 4976 12292 4984
rect 1244 4956 1252 4964
rect 556 4936 564 4944
rect 1372 4956 1380 4964
rect 3852 4956 3860 4964
rect 6636 4956 6644 4964
rect 2508 4936 2516 4944
rect 6460 4936 6468 4944
rect 7772 4956 7780 4964
rect 8396 4956 8404 4964
rect 12348 4956 12356 4964
rect 12908 4956 12916 4964
rect 9580 4936 9588 4944
rect 3244 4916 3252 4924
rect 3852 4916 3860 4924
rect 4540 4916 4548 4924
rect 5084 4916 5092 4924
rect 5324 4916 5332 4924
rect 5420 4916 5428 4924
rect 5484 4916 5492 4924
rect 7388 4916 7396 4924
rect 7772 4916 7780 4924
rect 12332 4916 12340 4924
rect 12588 4918 12596 4924
rect 12588 4916 12596 4918
rect 460 4896 468 4904
rect 556 4896 564 4904
rect 1196 4896 1204 4904
rect 1244 4896 1252 4904
rect 1820 4896 1828 4904
rect 2380 4896 2388 4904
rect 2508 4896 2516 4904
rect 3116 4896 3124 4904
rect 3756 4896 3764 4904
rect 3820 4896 3828 4904
rect 5052 4896 5060 4904
rect 7596 4896 7604 4904
rect 7724 4896 7732 4904
rect 7964 4896 7972 4904
rect 8524 4896 8532 4904
rect 8636 4896 8644 4904
rect 5196 4876 5204 4884
rect 5372 4876 5380 4884
rect 8092 4876 8100 4884
rect 9308 4896 9316 4904
rect 9884 4896 9892 4904
rect 10540 4896 10548 4904
rect 10636 4896 10644 4904
rect 11180 4896 11188 4904
rect 11676 4896 11684 4904
rect 11948 4896 11956 4904
rect 12492 4896 12500 4904
rect 108 4856 116 4864
rect 3212 4856 3220 4864
rect 5068 4856 5076 4864
rect 5356 4856 5364 4864
rect 7900 4856 7908 4864
rect 9788 4856 9796 4864
rect 12604 4856 12612 4864
rect 3308 4836 3316 4844
rect 6988 4836 6996 4844
rect 7532 4836 7540 4844
rect 10860 4836 10868 4844
rect 4828 4816 4836 4824
rect 5916 4816 5924 4824
rect 8652 4816 8660 4824
rect 10716 4816 10724 4824
rect 3020 4796 3028 4804
rect 4012 4796 4020 4804
rect 4956 4796 4964 4804
rect 6748 4796 6756 4804
rect 7132 4796 7140 4804
rect 7388 4796 7396 4804
rect 1148 4776 1156 4784
rect 1884 4776 1892 4784
rect 2524 4776 2532 4784
rect 3788 4776 3796 4784
rect 4716 4776 4724 4784
rect 4924 4776 4932 4784
rect 5052 4776 5060 4784
rect 6380 4776 6388 4784
rect 1980 4756 1988 4764
rect 3020 4756 3028 4764
rect 5020 4756 5028 4764
rect 5036 4756 5044 4764
rect 476 4736 484 4744
rect 1372 4736 1380 4744
rect 2652 4736 2660 4744
rect 3068 4736 3076 4744
rect 3228 4736 3236 4744
rect 4412 4736 4420 4744
rect 4684 4736 4692 4744
rect 7212 4736 7220 4744
rect 7404 4736 7412 4744
rect 7740 4736 7748 4744
rect 8316 4736 8324 4744
rect 412 4716 420 4724
rect 1164 4716 1172 4724
rect 1676 4716 1684 4724
rect 2060 4716 2068 4724
rect 2188 4716 2196 4724
rect 3260 4716 3268 4724
rect 4428 4716 4436 4724
rect 4668 4716 4676 4724
rect 5276 4716 5284 4724
rect 5388 4716 5396 4724
rect 5980 4716 5988 4724
rect 7036 4716 7044 4724
rect 7084 4716 7092 4724
rect 7708 4716 7716 4724
rect 8588 4716 8596 4724
rect 9244 4716 9252 4724
rect 1580 4696 1588 4704
rect 3228 4696 3236 4704
rect 3244 4696 3252 4704
rect 3388 4696 3396 4704
rect 3500 4696 3508 4704
rect 4508 4696 4516 4704
rect 4796 4702 4804 4704
rect 4796 4696 4804 4702
rect 5820 4696 5828 4704
rect 6572 4696 6580 4704
rect 7772 4696 7780 4704
rect 8444 4696 8452 4704
rect 10860 4736 10868 4744
rect 10972 4736 10980 4744
rect 11244 4736 11252 4744
rect 12220 4736 12228 4744
rect 10268 4716 10276 4724
rect 10844 4716 10852 4724
rect 11292 4716 11300 4724
rect 12108 4716 12116 4724
rect 3292 4676 3300 4684
rect 8444 4676 8452 4684
rect 8684 4676 8692 4684
rect 9324 4696 9332 4704
rect 11116 4696 11124 4704
rect 9324 4676 9332 4684
rect 5100 4656 5108 4664
rect 5324 4656 5332 4664
rect 10156 4656 10164 4664
rect 9020 4636 9028 4644
rect 492 4616 500 4624
rect 5500 4616 5508 4624
rect 7036 4616 7044 4624
rect 7404 4616 7412 4624
rect 9708 4616 9716 4624
rect 556 4596 564 4604
rect 6428 4596 6436 4604
rect 6460 4596 6468 4604
rect 7772 4596 7780 4604
rect 8364 4596 8372 4604
rect 9692 4596 9700 4604
rect 10268 4596 10276 4604
rect 11820 4576 11828 4584
rect 1292 4556 1300 4564
rect 4780 4556 4788 4564
rect 5452 4556 5460 4564
rect 7708 4556 7716 4564
rect 8748 4556 8756 4564
rect 9724 4556 9732 4564
rect 572 4536 580 4544
rect 1244 4536 1252 4544
rect 1116 4516 1124 4524
rect 1580 4516 1588 4524
rect 1804 4516 1812 4524
rect 6428 4516 6436 4524
rect 6764 4516 6772 4524
rect 7644 4516 7652 4524
rect 7756 4516 7764 4524
rect 8556 4516 8564 4524
rect 8668 4516 8676 4524
rect 9740 4516 9748 4524
rect 10348 4516 10356 4524
rect 12108 4516 12116 4524
rect 12300 4516 12308 4524
rect 428 4496 436 4504
rect 572 4496 580 4504
rect 1804 4496 1812 4504
rect 2700 4496 2708 4504
rect 2860 4496 2868 4504
rect 3292 4496 3300 4504
rect 3484 4496 3492 4504
rect 4044 4496 4052 4504
rect 4828 4496 4836 4504
rect 5452 4496 5460 4504
rect 6012 4496 6020 4504
rect 6380 4496 6388 4504
rect 6460 4496 6468 4504
rect 6636 4496 6644 4504
rect 8300 4496 8308 4504
rect 8364 4496 8372 4504
rect 9020 4496 9028 4504
rect 9708 4496 9716 4504
rect 9980 4496 9988 4504
rect 10460 4496 10468 4504
rect 10572 4496 10580 4504
rect 11196 4496 11204 4504
rect 12348 4496 12356 4504
rect 76 4476 84 4484
rect 2092 4476 2100 4484
rect 3260 4476 3268 4484
rect 6428 4476 6436 4484
rect 11516 4476 11524 4484
rect 12284 4476 12292 4484
rect 2812 4456 2820 4464
rect 8444 4436 8452 4444
rect 10684 4436 10692 4444
rect 60 4416 68 4424
rect 444 4416 452 4424
rect 1820 4416 1828 4424
rect 1980 4416 1988 4424
rect 2476 4416 2484 4424
rect 8316 4416 8324 4424
rect 1340 4396 1348 4404
rect 1804 4396 1812 4404
rect 11516 4396 11524 4404
rect 2444 4376 2452 4384
rect 3468 4376 3476 4384
rect 4172 4376 4180 4384
rect 5436 4376 5444 4384
rect 6764 4376 6772 4384
rect 11932 4376 11940 4384
rect 44 4356 52 4364
rect 3228 4356 3236 4364
rect 3436 4356 3444 4364
rect 10620 4356 10628 4364
rect 11276 4356 11284 4364
rect 492 4336 500 4344
rect 3356 4336 3364 4344
rect 5180 4336 5188 4344
rect 556 4316 564 4324
rect 1164 4316 1172 4324
rect 1820 4316 1828 4324
rect 1852 4316 1860 4324
rect 3100 4316 3108 4324
rect 3340 4316 3348 4324
rect 3516 4316 3524 4324
rect 3532 4316 3540 4324
rect 4428 4316 4436 4324
rect 4940 4316 4948 4324
rect 5084 4316 5092 4324
rect 5116 4316 5124 4324
rect 5644 4316 5652 4324
rect 620 4296 628 4304
rect 1964 4296 1972 4304
rect 3228 4296 3236 4304
rect 3468 4296 3476 4304
rect 5180 4296 5188 4304
rect 5804 4276 5812 4284
rect 6348 4316 6356 4324
rect 6428 4316 6436 4324
rect 6636 4316 6644 4324
rect 6652 4316 6660 4324
rect 7292 4316 7300 4324
rect 7420 4316 7428 4324
rect 7772 4316 7780 4324
rect 8988 4316 8996 4324
rect 9596 4316 9604 4324
rect 10252 4316 10260 4324
rect 10316 4316 10324 4324
rect 10476 4316 10484 4324
rect 10684 4316 10692 4324
rect 10796 4316 10804 4324
rect 11948 4316 11956 4324
rect 12444 4316 12452 4324
rect 6764 4296 6772 4304
rect 7372 4296 7380 4304
rect 7852 4296 7860 4304
rect 7884 4296 7892 4304
rect 7948 4296 7956 4304
rect 10332 4296 10340 4304
rect 10492 4296 10500 4304
rect 10572 4296 10580 4304
rect 11932 4302 11940 4304
rect 11932 4296 11940 4302
rect 12396 4296 12404 4304
rect 7100 4276 7108 4284
rect 7420 4276 7428 4284
rect 11308 4276 11316 4284
rect 7068 4256 7076 4264
rect 7084 4256 7092 4264
rect 10396 4256 10404 4264
rect 10556 4256 10564 4264
rect 8300 4236 8308 4244
rect 8700 4236 8708 4244
rect 3196 4216 3204 4224
rect 4156 4216 4164 4224
rect 5468 4216 5476 4224
rect 8876 4216 8884 4224
rect 10492 4216 10500 4224
rect 4412 4196 4420 4204
rect 4508 4196 4516 4204
rect 6428 4196 6436 4204
rect 9596 4196 9604 4204
rect 10316 4196 10324 4204
rect 12396 4196 12404 4204
rect 12444 4196 12452 4204
rect 1308 4176 1316 4184
rect 1852 4176 1860 4184
rect 1196 4136 1204 4144
rect 3148 4156 3156 4164
rect 3836 4136 3844 4144
rect 5148 4136 5156 4144
rect 7372 4136 7380 4144
rect 1308 4116 1316 4124
rect 2828 4118 2836 4124
rect 2828 4116 2836 4118
rect 3004 4116 3012 4124
rect 3468 4116 3476 4124
rect 6460 4116 6468 4124
rect 10348 4176 10356 4184
rect 10476 4176 10484 4184
rect 11052 4176 11060 4184
rect 11004 4156 11012 4164
rect 12092 4156 12100 4164
rect 12940 4156 12948 4164
rect 11100 4136 11108 4144
rect 588 4096 596 4104
rect 1164 4096 1172 4104
rect 1196 4096 1204 4104
rect 1868 4096 1876 4104
rect 2460 4096 2468 4104
rect 2876 4096 2884 4104
rect 3180 4096 3188 4104
rect 3372 4096 3380 4104
rect 4044 4096 4052 4104
rect 4956 4096 4964 4104
rect 5148 4096 5156 4104
rect 5196 4096 5204 4104
rect 6236 4096 6244 4104
rect 6380 4096 6388 4104
rect 6412 4096 6420 4104
rect 6620 4096 6628 4104
rect 508 4076 516 4084
rect 620 4076 628 4084
rect 2316 4076 2324 4084
rect 3132 4076 3140 4084
rect 6636 4076 6644 4084
rect 6716 4076 6724 4084
rect 7292 4076 7300 4084
rect 8508 4116 8516 4124
rect 10428 4116 10436 4124
rect 10652 4116 10660 4124
rect 11020 4116 11028 4124
rect 11084 4116 11092 4124
rect 12092 4116 12100 4124
rect 12300 4116 12308 4124
rect 12972 4116 12980 4124
rect 7948 4096 7956 4104
rect 8572 4096 8580 4104
rect 9180 4096 9188 4104
rect 9916 4096 9924 4104
rect 10796 4096 10804 4104
rect 11276 4096 11284 4104
rect 12220 4096 12228 4104
rect 12860 4096 12868 4104
rect 12908 4096 12916 4104
rect 8540 4076 8548 4084
rect 9932 4076 9940 4084
rect 12284 4076 12292 4084
rect 172 4056 180 4064
rect 4044 4056 4052 4064
rect 5180 4056 5188 4064
rect 7100 4056 7108 4064
rect 12156 4056 12164 4064
rect 492 4036 500 4044
rect 3180 4036 3188 4044
rect 3196 4036 3204 4044
rect 6956 4036 6964 4044
rect 1164 4016 1172 4024
rect 2460 4016 2468 4024
rect 5452 4016 5460 4024
rect 7116 4016 7124 4024
rect 7308 4036 7316 4044
rect 7804 4016 7812 4024
rect 11084 4016 11092 4024
rect 908 3996 916 4004
rect 1820 3996 1828 4004
rect 3836 3996 3844 4004
rect 4956 3996 4964 4004
rect 5068 3996 5076 4004
rect 2668 3976 2676 3984
rect 3468 3976 3476 3984
rect 7932 3956 7940 3964
rect 7948 3956 7956 3964
rect 8316 3956 8324 3964
rect 2860 3936 2868 3944
rect 3340 3936 3348 3944
rect 5100 3936 5108 3944
rect 6060 3936 6068 3944
rect 92 3916 100 3924
rect 172 3916 180 3924
rect 1100 3916 1108 3924
rect 1324 3916 1332 3924
rect 1820 3916 1828 3924
rect 3148 3916 3156 3924
rect 3196 3916 3204 3924
rect 3772 3916 3780 3924
rect 4316 3916 4324 3924
rect 5452 3916 5460 3924
rect 6124 3916 6132 3924
rect 6620 3916 6628 3924
rect 7292 3916 7300 3924
rect 60 3896 68 3904
rect 636 3896 644 3904
rect 1676 3896 1684 3904
rect 1996 3896 2004 3904
rect 2076 3896 2084 3904
rect 3212 3896 3220 3904
rect 4780 3902 4788 3904
rect 4780 3896 4788 3902
rect 6332 3896 6340 3904
rect 6492 3896 6500 3904
rect 7388 3902 7396 3904
rect 7388 3896 7396 3902
rect 124 3876 132 3884
rect 1676 3876 1684 3884
rect 3484 3876 3492 3884
rect 3868 3856 3876 3864
rect 7388 3856 7396 3864
rect 8524 3936 8532 3944
rect 11004 3936 11012 3944
rect 12844 3936 12852 3944
rect 8316 3916 8324 3924
rect 8972 3916 8980 3924
rect 9196 3916 9204 3924
rect 9628 3916 9636 3924
rect 10284 3916 10292 3924
rect 11052 3916 11060 3924
rect 11452 3916 11460 3924
rect 11676 3916 11684 3924
rect 11820 3916 11828 3924
rect 12940 3916 12948 3924
rect 8684 3896 8692 3904
rect 9084 3896 9092 3904
rect 9836 3896 9844 3904
rect 9996 3896 10004 3904
rect 11100 3896 11108 3904
rect 8684 3876 8692 3884
rect 11308 3876 11316 3884
rect 11964 3876 11972 3884
rect 12972 3896 12980 3904
rect 10844 3856 10852 3864
rect 3836 3816 3844 3824
rect 6412 3816 6420 3824
rect 6460 3816 6468 3824
rect 7772 3816 7780 3824
rect 8540 3816 8548 3824
rect 9196 3816 9204 3824
rect 60 3796 68 3804
rect 92 3796 100 3804
rect 5948 3796 5956 3804
rect 6364 3776 6372 3784
rect 8508 3776 8516 3784
rect 6636 3756 6644 3764
rect 5644 3736 5652 3744
rect 8636 3736 8644 3744
rect 908 3716 916 3724
rect 2060 3716 2068 3724
rect 3324 3716 3332 3724
rect 4124 3716 4132 3724
rect 524 3696 532 3704
rect 796 3696 804 3704
rect 2044 3696 2052 3704
rect 3164 3696 3172 3704
rect 3388 3696 3396 3704
rect 3628 3696 3636 3704
rect 3852 3696 3860 3704
rect 5804 3716 5812 3724
rect 5948 3716 5956 3724
rect 6124 3696 6132 3704
rect 6716 3716 6724 3724
rect 8572 3716 8580 3724
rect 8620 3716 8628 3724
rect 9740 3716 9748 3724
rect 9852 3716 9860 3724
rect 6748 3696 6756 3704
rect 5788 3676 5796 3684
rect 6508 3676 6516 3684
rect 8732 3696 8740 3704
rect 9628 3696 9636 3704
rect 9884 3696 9892 3704
rect 7900 3676 7908 3684
rect 9868 3676 9876 3684
rect 11804 3816 11812 3824
rect 12316 3816 12324 3824
rect 10412 3796 10420 3804
rect 10492 3796 10500 3804
rect 11756 3776 11764 3784
rect 11964 3736 11972 3744
rect 12300 3736 12308 3744
rect 12588 3736 12596 3744
rect 12316 3716 12324 3724
rect 10972 3696 10980 3704
rect 11196 3696 11204 3704
rect 12220 3696 12228 3704
rect 2668 3656 2676 3664
rect 5116 3656 5124 3664
rect 5852 3656 5860 3664
rect 7900 3656 7908 3664
rect 12220 3656 12228 3664
rect 1708 3636 1716 3644
rect 2332 3636 2340 3644
rect 4588 3636 4596 3644
rect 508 3616 516 3624
rect 3132 3616 3140 3624
rect 5324 3616 5332 3624
rect 6780 3616 6788 3624
rect 6796 3616 6804 3624
rect 8988 3616 8996 3624
rect 11100 3616 11108 3624
rect 524 3576 532 3584
rect 7068 3576 7076 3584
rect 7708 3576 7716 3584
rect 9020 3556 9028 3564
rect 1292 3536 1300 3544
rect 3180 3536 3188 3544
rect 5404 3536 5412 3544
rect 6060 3536 6068 3544
rect 7388 3536 7396 3544
rect 92 3516 100 3524
rect 156 3516 164 3524
rect 1132 3516 1140 3524
rect 1692 3516 1700 3524
rect 1852 3516 1860 3524
rect 2092 3516 2100 3524
rect 3996 3516 4004 3524
rect 4172 3516 4180 3524
rect 4620 3516 4628 3524
rect 4844 3516 4852 3524
rect 5692 3516 5700 3524
rect 6092 3516 6100 3524
rect 6636 3516 6644 3524
rect 7436 3516 7444 3524
rect 7948 3516 7956 3524
rect 60 3496 68 3504
rect 1260 3496 1268 3504
rect 3132 3496 3140 3504
rect 3212 3496 3220 3504
rect 3532 3496 3540 3504
rect 124 3476 132 3484
rect 7388 3502 7396 3504
rect 7388 3496 7396 3502
rect 7756 3496 7764 3504
rect 8588 3516 8596 3524
rect 9068 3516 9076 3524
rect 9756 3536 9764 3544
rect 9996 3536 10004 3544
rect 9276 3516 9284 3524
rect 10316 3516 10324 3524
rect 10348 3516 10356 3524
rect 10444 3516 10452 3524
rect 10604 3516 10612 3524
rect 11180 3516 11188 3524
rect 12236 3516 12244 3524
rect 9068 3496 9076 3504
rect 9340 3502 9348 3504
rect 9340 3496 9348 3502
rect 2364 3476 2372 3484
rect 3228 3476 3236 3484
rect 3356 3476 3364 3484
rect 3532 3476 3540 3484
rect 4028 3456 4036 3464
rect 4796 3476 4804 3484
rect 7756 3476 7764 3484
rect 9276 3476 9284 3484
rect 6124 3456 6132 3464
rect 9708 3456 9716 3464
rect 7148 3436 7156 3444
rect 9564 3436 9572 3444
rect 3948 3416 3956 3424
rect 60 3396 68 3404
rect 92 3396 100 3404
rect 2524 3396 2532 3404
rect 3340 3396 3348 3404
rect 3996 3396 4004 3404
rect 524 3376 532 3384
rect 1260 3356 1268 3364
rect 1948 3356 1956 3364
rect 6428 3356 6436 3364
rect 9020 3356 9028 3364
rect 9820 3356 9828 3364
rect 556 3336 564 3344
rect 1948 3316 1956 3324
rect 2060 3316 2068 3324
rect 2572 3316 2580 3324
rect 2684 3316 2692 3324
rect 2780 3316 2788 3324
rect 4204 3316 4212 3324
rect 4316 3318 4324 3324
rect 9708 3336 9716 3344
rect 9852 3336 9860 3344
rect 4316 3316 4324 3318
rect 7084 3316 7092 3324
rect 7420 3316 7428 3324
rect 7436 3316 7444 3324
rect 7580 3316 7588 3324
rect 9708 3316 9716 3324
rect 10380 3496 10388 3504
rect 11084 3496 11092 3504
rect 11116 3496 11124 3504
rect 10652 3476 10660 3484
rect 10316 3396 10324 3404
rect 11644 3396 11652 3404
rect 11772 3396 11780 3404
rect 12236 3396 12244 3404
rect 10956 3356 10964 3364
rect 11724 3356 11732 3364
rect 11052 3316 11060 3324
rect 11644 3316 11652 3324
rect 524 3296 532 3304
rect 556 3296 564 3304
rect 1164 3296 1172 3304
rect 1260 3296 1268 3304
rect 1740 3296 1748 3304
rect 2540 3296 2548 3304
rect 2860 3296 2868 3304
rect 3340 3296 3348 3304
rect 4060 3296 4068 3304
rect 4796 3296 4804 3304
rect 6284 3296 6292 3304
rect 6428 3296 6436 3304
rect 7068 3296 7076 3304
rect 7996 3296 8004 3304
rect 9020 3296 9028 3304
rect 9692 3296 9700 3304
rect 10956 3296 10964 3304
rect 11436 3296 11444 3304
rect 11612 3296 11620 3304
rect 11628 3296 11636 3304
rect 11932 3318 11940 3324
rect 11932 3316 11940 3318
rect 3308 3276 3316 3284
rect 3932 3276 3940 3284
rect 9564 3276 9572 3284
rect 9916 3276 9924 3284
rect 1740 3256 1748 3264
rect 1980 3256 1988 3264
rect 2012 3256 2020 3264
rect 11196 3256 11204 3264
rect 748 3236 756 3244
rect 3516 3236 3524 3244
rect 11052 3236 11060 3244
rect 12844 3216 12852 3224
rect 12972 3216 12980 3224
rect 4828 3196 4836 3204
rect 11196 3196 11204 3204
rect 4796 3176 4804 3184
rect 10492 3176 10500 3184
rect 1548 3156 1556 3164
rect 2460 3156 2468 3164
rect 3372 3156 3380 3164
rect 6780 3156 6788 3164
rect 7692 3156 7700 3164
rect 9388 3156 9396 3164
rect 11196 3156 11204 3164
rect 4652 3136 4660 3144
rect 6620 3136 6628 3144
rect 8012 3136 8020 3144
rect 9340 3136 9348 3144
rect 9932 3136 9940 3144
rect 10604 3136 10612 3144
rect 11804 3136 11812 3144
rect 1404 3116 1412 3124
rect 1548 3116 1556 3124
rect 2460 3116 2468 3124
rect 2572 3116 2580 3124
rect 3772 3116 3780 3124
rect 4332 3116 4340 3124
rect 1388 3096 1396 3104
rect 2684 3096 2692 3104
rect 3084 3102 3092 3104
rect 3084 3096 3092 3102
rect 3628 3096 3636 3104
rect 3868 3096 3876 3104
rect 4076 3096 4084 3104
rect 6268 3116 6276 3124
rect 6380 3116 6388 3124
rect 6428 3116 6436 3124
rect 6604 3116 6612 3124
rect 6620 3116 6628 3124
rect 7804 3116 7812 3124
rect 7932 3116 7940 3124
rect 8044 3116 8052 3124
rect 8540 3116 8548 3124
rect 8732 3116 8740 3124
rect 9244 3116 9252 3124
rect 9820 3116 9828 3124
rect 10636 3116 10644 3124
rect 11196 3116 11204 3124
rect 11740 3116 11748 3124
rect 12428 3116 12436 3124
rect 4652 3096 4660 3104
rect 5276 3096 5284 3104
rect 6588 3096 6596 3104
rect 10412 3096 10420 3104
rect 10428 3096 10436 3104
rect 11084 3096 11092 3104
rect 11308 3096 11316 3104
rect 12460 3096 12468 3104
rect 6380 3076 6388 3084
rect 8028 3076 8036 3084
rect 8540 3076 8548 3084
rect 11964 3076 11972 3084
rect 3356 3056 3364 3064
rect 6620 3056 6628 3064
rect 7996 3056 8004 3064
rect 8540 3036 8548 3044
rect 156 3016 164 3024
rect 1388 3016 1396 3024
rect 3276 3016 3284 3024
rect 3980 3016 3988 3024
rect 6588 3016 6596 3024
rect 9052 3016 9060 3024
rect 2092 2996 2100 3004
rect 1404 2976 1412 2984
rect 604 2956 612 2964
rect 7708 2956 7716 2964
rect 7964 2956 7972 2964
rect 748 2936 756 2944
rect 2348 2936 2356 2944
rect 5340 2936 5348 2944
rect 700 2916 708 2924
rect 1948 2916 1956 2924
rect 4540 2916 4548 2924
rect 4812 2916 4820 2924
rect 7116 2916 7124 2924
rect 7228 2916 7236 2924
rect 8572 2916 8580 2924
rect 11612 3016 11620 3024
rect 9852 2996 9860 3004
rect 9788 2956 9796 2964
rect 11644 2956 11652 2964
rect 11084 2936 11092 2944
rect 11276 2936 11284 2944
rect 11932 2936 11940 2944
rect 11964 2916 11972 2924
rect 508 2896 516 2904
rect 604 2896 612 2904
rect 1100 2896 1108 2904
rect 1804 2896 1812 2904
rect 2092 2896 2100 2904
rect 2524 2896 2532 2904
rect 4316 2896 4324 2904
rect 4620 2896 4628 2904
rect 4796 2896 4804 2904
rect 5276 2896 5284 2904
rect 5340 2896 5348 2904
rect 5996 2896 6004 2904
rect 6956 2896 6964 2904
rect 7084 2896 7092 2904
rect 8220 2896 8228 2904
rect 8540 2896 8548 2904
rect 8588 2896 8596 2904
rect 8684 2896 8692 2904
rect 9180 2896 9188 2904
rect 9884 2896 9892 2904
rect 10556 2896 10564 2904
rect 11100 2896 11108 2904
rect 11308 2896 11316 2904
rect 11804 2896 11812 2904
rect 11836 2896 11844 2904
rect 1756 2876 1764 2884
rect 2236 2876 2244 2884
rect 3852 2876 3860 2884
rect 6924 2876 6932 2884
rect 2124 2856 2132 2864
rect 2300 2856 2308 2864
rect 3884 2856 3892 2864
rect 5884 2856 5892 2864
rect 6028 2856 6036 2864
rect 7452 2856 7460 2864
rect 4844 2836 4852 2844
rect 11276 2836 11284 2844
rect 11948 2836 11956 2844
rect 6044 2816 6052 2824
rect 11772 2816 11780 2824
rect 1804 2796 1812 2804
rect 4828 2796 4836 2804
rect 6492 2796 6500 2804
rect 10796 2796 10804 2804
rect 2428 2776 2436 2784
rect 3052 2776 3060 2784
rect 4076 2776 4084 2784
rect 6908 2776 6916 2784
rect 9052 2776 9060 2784
rect 524 2756 532 2764
rect 2668 2756 2676 2764
rect 3420 2756 3428 2764
rect 5340 2756 5348 2764
rect 2188 2736 2196 2744
rect 4780 2736 4788 2744
rect 524 2716 532 2724
rect 556 2716 564 2724
rect 1164 2716 1172 2724
rect 3004 2716 3012 2724
rect 3388 2716 3396 2724
rect 4428 2716 4436 2724
rect 4636 2716 4644 2724
rect 4700 2716 4708 2724
rect 5916 2736 5924 2744
rect 7580 2736 7588 2744
rect 7772 2736 7780 2744
rect 8124 2736 8132 2744
rect 10348 2736 10356 2744
rect 10588 2736 10596 2744
rect 5340 2716 5348 2724
rect 6268 2716 6276 2724
rect 7020 2716 7028 2724
rect 8012 2716 8020 2724
rect 8316 2716 8324 2724
rect 8972 2716 8980 2724
rect 9516 2716 9524 2724
rect 9660 2716 9668 2724
rect 9916 2716 9924 2724
rect 10540 2716 10548 2724
rect 10636 2716 10644 2724
rect 11004 2716 11012 2724
rect 11644 2716 11652 2724
rect 11724 2716 11732 2724
rect 11836 2716 11844 2724
rect 620 2696 628 2704
rect 1900 2696 1908 2704
rect 3180 2696 3182 2704
rect 3182 2696 3188 2704
rect 3276 2696 3284 2704
rect 3548 2696 3556 2704
rect 4636 2696 4644 2704
rect 4764 2702 4772 2704
rect 4764 2696 4772 2702
rect 5436 2702 5444 2704
rect 5436 2696 5444 2702
rect 6348 2696 6356 2704
rect 7788 2696 7796 2704
rect 9708 2696 9716 2704
rect 9980 2702 9988 2704
rect 9980 2696 9988 2702
rect 10396 2696 10404 2704
rect 11548 2696 11556 2704
rect 11948 2702 11956 2704
rect 11948 2696 11956 2702
rect 4204 2676 4212 2684
rect 7020 2676 7028 2684
rect 3388 2656 3396 2664
rect 6108 2636 6116 2644
rect 8732 2636 8740 2644
rect 460 2616 468 2624
rect 1164 2616 1172 2624
rect 3132 2616 3140 2624
rect 3964 2616 3972 2624
rect 4636 2616 4644 2624
rect 5916 2616 5924 2624
rect 8972 2616 8980 2624
rect 10044 2616 10052 2624
rect 76 2596 84 2604
rect 556 2596 564 2604
rect 4764 2596 4772 2604
rect 5772 2596 5780 2604
rect 9660 2596 9668 2604
rect 9740 2596 9748 2604
rect 11836 2596 11844 2604
rect 12284 2596 12292 2604
rect 620 2576 628 2584
rect 3836 2576 3844 2584
rect 9708 2576 9716 2584
rect 5804 2556 5812 2564
rect 8364 2556 8372 2564
rect 8428 2556 8436 2564
rect 1196 2536 1204 2544
rect 3004 2536 3012 2544
rect 3804 2536 3812 2544
rect 5996 2536 6004 2544
rect 8700 2536 8708 2544
rect 11036 2556 11044 2564
rect 12348 2556 12356 2564
rect 10044 2536 10052 2544
rect 76 2516 84 2524
rect 1292 2516 1300 2524
rect 1916 2516 1924 2524
rect 2844 2518 2852 2524
rect 2844 2516 2852 2518
rect 3836 2516 3844 2524
rect 4812 2516 4820 2524
rect 5852 2516 5860 2524
rect 6124 2516 6132 2524
rect 6748 2516 6756 2524
rect 6924 2516 6932 2524
rect 7212 2516 7220 2524
rect 8428 2516 8436 2524
rect 9116 2516 9124 2524
rect 9820 2516 9828 2524
rect 11004 2516 11012 2524
rect 11084 2516 11092 2524
rect 12300 2516 12308 2524
rect 12348 2516 12356 2524
rect 252 2496 260 2504
rect 1148 2496 1156 2504
rect 1708 2496 1716 2504
rect 1884 2496 1892 2504
rect 2348 2496 2356 2504
rect 2476 2496 2484 2504
rect 2796 2496 2804 2504
rect 3772 2496 3780 2504
rect 3804 2496 3812 2504
rect 3980 2496 3988 2504
rect 4316 2496 4324 2504
rect 4460 2496 4468 2504
rect 4620 2496 4628 2504
rect 4940 2496 4948 2504
rect 4956 2496 4964 2504
rect 5084 2496 5092 2504
rect 6348 2496 6356 2504
rect 6636 2496 6644 2504
rect 7532 2496 7540 2504
rect 7692 2496 7700 2504
rect 8572 2496 8580 2504
rect 9196 2496 9204 2504
rect 9372 2496 9380 2504
rect 9884 2496 9892 2504
rect 10940 2496 10948 2504
rect 11180 2496 11188 2504
rect 12220 2496 12228 2504
rect 12492 2496 12500 2504
rect 1756 2476 1764 2484
rect 3468 2476 3476 2484
rect 6428 2476 6436 2484
rect 9820 2476 9828 2484
rect 12284 2476 12292 2484
rect 3292 2456 3300 2464
rect 5244 2456 5252 2464
rect 6604 2456 6612 2464
rect 9884 2456 9892 2464
rect 12444 2456 12452 2464
rect 12492 2436 12500 2444
rect 252 2416 260 2424
rect 1100 2416 1108 2424
rect 3148 2416 3156 2424
rect 3324 2416 3332 2424
rect 3756 2416 3764 2424
rect 3772 2416 3780 2424
rect 3980 2416 3988 2424
rect 4588 2416 4596 2424
rect 7916 2416 7924 2424
rect 12412 2416 12420 2424
rect 1900 2396 1908 2404
rect 4668 2396 4676 2404
rect 8908 2396 8916 2404
rect 8428 2376 8436 2384
rect 11836 2376 11844 2384
rect 252 2356 260 2364
rect 4924 2356 4932 2364
rect 7100 2356 7108 2364
rect 9980 2356 9988 2364
rect 156 2336 164 2344
rect 3068 2336 3076 2344
rect 252 2316 260 2324
rect 1196 2316 1204 2324
rect 1836 2316 1844 2324
rect 2188 2316 2196 2324
rect 3164 2316 3172 2324
rect 4988 2336 4996 2344
rect 5148 2336 5156 2344
rect 5884 2336 5892 2344
rect 3628 2316 3636 2324
rect 3884 2316 3892 2324
rect 3948 2316 3956 2324
rect 4796 2316 4804 2324
rect 5132 2316 5140 2324
rect 5276 2316 5284 2324
rect 7532 2336 7540 2344
rect 7996 2336 8004 2344
rect 11564 2336 11572 2344
rect 5932 2316 5940 2324
rect 6108 2316 6116 2324
rect 6604 2316 6612 2324
rect 6636 2316 6644 2324
rect 7804 2316 7812 2324
rect 8012 2316 8020 2324
rect 8604 2316 8612 2324
rect 9260 2316 9268 2324
rect 140 2302 148 2304
rect 140 2296 148 2302
rect 2028 2296 2036 2304
rect 3244 2296 3252 2304
rect 4940 2296 4948 2304
rect 4956 2296 4964 2304
rect 5692 2296 5700 2304
rect 5852 2296 5860 2304
rect 6428 2296 6436 2304
rect 9580 2296 9588 2304
rect 10316 2316 10324 2324
rect 10924 2316 10932 2324
rect 11036 2316 11044 2324
rect 11804 2316 11812 2324
rect 11836 2316 11844 2324
rect 10380 2296 10388 2304
rect 11676 2296 11684 2304
rect 11948 2302 11956 2304
rect 11948 2296 11956 2302
rect 1292 2276 1300 2284
rect 3116 2256 3124 2264
rect 9052 2256 9060 2264
rect 12220 2256 12228 2264
rect 508 2216 516 2224
rect 10316 2196 10324 2204
rect 1164 2176 1172 2184
rect 6492 2176 6500 2184
rect 10380 2176 10388 2184
rect 1260 2156 1268 2164
rect 2796 2156 2804 2164
rect 3260 2156 3268 2164
rect 556 2136 564 2144
rect 1196 2136 1204 2144
rect 3340 2136 3348 2144
rect 5148 2136 5156 2144
rect 5788 2136 5796 2144
rect 6412 2136 6420 2144
rect 7148 2156 7156 2164
rect 1260 2116 1268 2124
rect 1900 2116 1908 2124
rect 2556 2116 2564 2124
rect 2796 2116 2804 2124
rect 8636 2136 8644 2144
rect 9980 2136 9988 2144
rect 10636 2136 10644 2144
rect 11948 2136 11956 2144
rect 2956 2116 2964 2124
rect 4204 2116 4212 2124
rect 4540 2116 4548 2124
rect 4988 2116 4996 2124
rect 6492 2116 6500 2124
rect 7148 2116 7156 2124
rect 7196 2116 7204 2124
rect 7804 2116 7812 2124
rect 7820 2116 7828 2124
rect 9340 2116 9348 2124
rect 172 2096 180 2104
rect 556 2096 564 2104
rect 1164 2096 1172 2104
rect 1196 2096 1204 2104
rect 1836 2096 1844 2104
rect 1884 2096 1892 2104
rect 2460 2096 2468 2104
rect 2668 2096 2676 2104
rect 2844 2096 2852 2104
rect 3772 2096 3780 2104
rect 3916 2096 3924 2104
rect 5100 2096 5108 2104
rect 5356 2096 5364 2104
rect 6140 2096 6148 2104
rect 6300 2096 6308 2104
rect 6412 2096 6420 2104
rect 6908 2096 6916 2104
rect 7644 2096 7652 2104
rect 8060 2096 8068 2104
rect 9260 2096 9268 2104
rect 9884 2096 9892 2104
rect 10140 2096 10148 2104
rect 10684 2096 10692 2104
rect 11308 2096 11316 2104
rect 11772 2096 11780 2104
rect 2028 2076 2036 2084
rect 2428 2076 2436 2084
rect 2572 2076 2580 2084
rect 2956 2076 2964 2084
rect 4412 2076 4420 2084
rect 4956 2076 4964 2084
rect 5388 2076 5396 2084
rect 6412 2076 6420 2084
rect 8636 2076 8644 2084
rect 11804 2076 11812 2084
rect 2108 2056 2116 2064
rect 6268 2056 6276 2064
rect 10348 2056 10356 2064
rect 156 2036 164 2044
rect 428 2036 436 2044
rect 3820 2016 3828 2024
rect 3948 2016 3956 2024
rect 5932 2016 5940 2024
rect 6284 2036 6292 2044
rect 12204 2036 12212 2044
rect 140 1996 148 2004
rect 6380 1996 6388 2004
rect 6604 1996 6612 2004
rect 10428 1996 10436 2004
rect 11308 1996 11316 2004
rect 3804 1976 3812 1984
rect 5852 1976 5860 1984
rect 7644 1976 7652 1984
rect 524 1956 532 1964
rect 4028 1956 4036 1964
rect 8316 1956 8324 1964
rect 10940 1956 10948 1964
rect 476 1936 484 1944
rect 3964 1936 3972 1944
rect 524 1916 532 1924
rect 1100 1916 1108 1924
rect 1644 1916 1652 1924
rect 2380 1916 2388 1924
rect 3020 1916 3028 1924
rect 3340 1916 3348 1924
rect 3500 1916 3508 1924
rect 3980 1916 3988 1924
rect 3996 1916 4004 1924
rect 4044 1916 4052 1924
rect 7228 1936 7236 1944
rect 9036 1936 9044 1944
rect 10492 1936 10500 1944
rect 11004 1936 11012 1944
rect 11196 1936 11204 1944
rect 6524 1916 6532 1924
rect 6636 1916 6644 1924
rect 8316 1916 8324 1924
rect 8380 1916 8388 1924
rect 8988 1916 8996 1924
rect 9004 1916 9012 1924
rect 9196 1916 9204 1924
rect 9852 1916 9860 1924
rect 9868 1916 9876 1924
rect 10940 1916 10948 1924
rect 11580 1916 11588 1924
rect 11820 1916 11828 1924
rect 620 1896 628 1904
rect 1884 1896 1892 1904
rect 3180 1896 3182 1904
rect 3182 1896 3188 1904
rect 3468 1896 3476 1904
rect 5228 1896 5236 1904
rect 6572 1896 6580 1904
rect 7388 1902 7396 1904
rect 7388 1896 7396 1902
rect 9052 1896 9060 1904
rect 9116 1896 9124 1904
rect 9788 1896 9796 1904
rect 11004 1896 11012 1904
rect 11932 1902 11940 1904
rect 11932 1896 11940 1902
rect 1948 1876 1956 1884
rect 3964 1876 3972 1884
rect 5276 1876 5284 1884
rect 2684 1856 2692 1864
rect 5132 1856 5140 1864
rect 7516 1836 7524 1844
rect 7948 1836 7956 1844
rect 1660 1816 1668 1824
rect 3996 1816 4004 1824
rect 6444 1816 6452 1824
rect 8380 1816 8388 1824
rect 172 1796 180 1804
rect 476 1796 484 1804
rect 6396 1796 6404 1804
rect 4556 1776 4564 1784
rect 10924 1776 10932 1784
rect 620 1756 628 1764
rect 3900 1756 3908 1764
rect 4540 1736 4548 1744
rect 4812 1736 4820 1744
rect 9244 1756 9252 1764
rect 11036 1756 11044 1764
rect 6060 1736 6068 1744
rect 11020 1736 11028 1744
rect 620 1716 628 1724
rect 1292 1716 1300 1724
rect 2572 1716 2580 1724
rect 3180 1716 3188 1724
rect 3900 1716 3908 1724
rect 4556 1716 4564 1724
rect 5804 1716 5812 1724
rect 6732 1718 6740 1724
rect 6732 1716 6740 1718
rect 9052 1716 9060 1724
rect 11036 1716 11044 1724
rect 11836 1716 11844 1724
rect 11932 1718 11940 1724
rect 11932 1716 11940 1718
rect 460 1696 468 1704
rect 1420 1696 1428 1704
rect 2364 1696 2372 1704
rect 3116 1696 3124 1704
rect 3772 1696 3780 1704
rect 3804 1696 3812 1704
rect 4828 1696 4836 1704
rect 5964 1696 5972 1704
rect 6124 1696 6132 1704
rect 6636 1696 6644 1704
rect 7420 1696 7428 1704
rect 7948 1696 7956 1704
rect 8972 1696 8980 1704
rect 9004 1696 9012 1704
rect 9244 1696 9252 1704
rect 10252 1696 10260 1704
rect 10908 1696 10916 1704
rect 11580 1696 11588 1704
rect 11804 1696 11812 1704
rect 476 1676 484 1684
rect 2636 1676 2644 1684
rect 4364 1676 4372 1684
rect 4620 1676 4628 1684
rect 7852 1676 7860 1684
rect 9004 1676 9012 1684
rect 2604 1656 2612 1664
rect 3468 1656 3476 1664
rect 7692 1656 7700 1664
rect 8460 1656 8468 1664
rect 8972 1656 8980 1664
rect 1756 1636 1764 1644
rect 3324 1636 3332 1644
rect 3772 1636 3780 1644
rect 6300 1636 6308 1644
rect 10924 1636 10932 1644
rect 11004 1636 11012 1644
rect 1420 1616 1428 1624
rect 2812 1616 2820 1624
rect 9644 1616 9652 1624
rect 636 1596 644 1604
rect 3020 1596 3028 1604
rect 3628 1596 3636 1604
rect 7580 1596 7588 1604
rect 1292 1576 1300 1584
rect 2412 1576 2420 1584
rect 9724 1576 9732 1584
rect 10492 1596 10500 1604
rect 3420 1556 3428 1564
rect 7084 1556 7092 1564
rect 8124 1556 8132 1564
rect 2828 1536 2836 1544
rect 3228 1536 3236 1544
rect 5420 1536 5428 1544
rect 12284 1536 12292 1544
rect 524 1516 532 1524
rect 1164 1516 1172 1524
rect 1260 1516 1268 1524
rect 1436 1516 1444 1524
rect 2460 1516 2468 1524
rect 2732 1516 2740 1524
rect 4012 1516 4020 1524
rect 4652 1516 4660 1524
rect 4684 1516 4692 1524
rect 6364 1516 6372 1524
rect 6380 1516 6388 1524
rect 7708 1516 7716 1524
rect 8220 1516 8228 1524
rect 9644 1516 9652 1524
rect 9660 1516 9668 1524
rect 10924 1516 10932 1524
rect 11132 1516 11140 1524
rect 1836 1496 1844 1504
rect 2316 1496 2324 1504
rect 2332 1496 2340 1504
rect 2828 1502 2836 1504
rect 2828 1496 2836 1502
rect 3484 1502 3492 1504
rect 3484 1496 3492 1502
rect 4332 1496 4340 1504
rect 4780 1502 4788 1504
rect 4780 1496 4788 1502
rect 7756 1496 7764 1504
rect 7772 1496 7780 1504
rect 8668 1502 8676 1504
rect 8668 1496 8676 1502
rect 9196 1496 9204 1504
rect 9996 1502 10004 1504
rect 9996 1496 10004 1502
rect 11068 1496 11076 1504
rect 12284 1496 12292 1504
rect 524 1476 532 1484
rect 604 1476 612 1484
rect 1436 1476 1444 1484
rect 1804 1476 1812 1484
rect 6364 1476 6372 1484
rect 1132 1456 1140 1464
rect 1500 1436 1508 1444
rect 796 1416 804 1424
rect 3212 1416 3220 1424
rect 3228 1416 3236 1424
rect 4332 1416 4340 1424
rect 5916 1416 5924 1424
rect 5932 1416 5940 1424
rect 7004 1416 7012 1424
rect 7708 1416 7716 1424
rect 716 1396 724 1404
rect 1100 1396 1108 1404
rect 2860 1396 2868 1404
rect 4012 1396 4020 1404
rect 5164 1396 5172 1404
rect 5420 1396 5428 1404
rect 6972 1396 6980 1404
rect 7420 1396 7428 1404
rect 1932 1356 1940 1364
rect 3804 1336 3812 1344
rect 8028 1336 8036 1344
rect 9340 1336 9348 1344
rect 76 1316 84 1324
rect 1500 1316 1508 1324
rect 1532 1318 1540 1324
rect 1532 1316 1540 1318
rect 2332 1316 2340 1324
rect 3084 1316 3092 1324
rect 5820 1316 5828 1324
rect 5932 1316 5940 1324
rect 6972 1316 6980 1324
rect 7404 1316 7412 1324
rect 9068 1316 9076 1324
rect 9324 1316 9332 1324
rect 9532 1316 9540 1324
rect 172 1296 180 1304
rect 892 1296 900 1304
rect 1564 1296 1572 1304
rect 2364 1296 2372 1304
rect 2572 1296 2580 1304
rect 2860 1296 2868 1304
rect 3772 1296 3780 1304
rect 3804 1296 3812 1304
rect 4316 1296 4324 1304
rect 5052 1296 5060 1304
rect 5164 1296 5172 1304
rect 5916 1296 5924 1304
rect 5996 1296 6004 1304
rect 6636 1296 6644 1304
rect 7308 1296 7316 1304
rect 7932 1296 7940 1304
rect 8460 1296 8468 1304
rect 9196 1296 9204 1304
rect 9212 1296 9220 1304
rect 9244 1296 9252 1304
rect 9388 1296 9396 1304
rect 10028 1296 10036 1304
rect 10652 1316 10660 1324
rect 11836 1316 11844 1324
rect 11932 1318 11940 1324
rect 11932 1316 11940 1318
rect 11292 1296 11300 1304
rect 11820 1296 11828 1304
rect 2428 1276 2436 1284
rect 2636 1276 2644 1284
rect 5836 1276 5844 1284
rect 6572 1276 6580 1284
rect 7772 1276 7780 1284
rect 11740 1276 11748 1284
rect 3772 1256 3780 1264
rect 5996 1256 6004 1264
rect 6604 1256 6612 1264
rect 9356 1256 9364 1264
rect 2540 1236 2548 1244
rect 8716 1236 8724 1244
rect 6428 1216 6436 1224
rect 6524 1216 6532 1224
rect 11660 1216 11668 1224
rect 140 1196 148 1204
rect 716 1196 724 1204
rect 908 1196 916 1204
rect 1532 1196 1540 1204
rect 9244 1196 9252 1204
rect 12860 1196 12868 1204
rect 4316 1176 4324 1184
rect 5052 1176 5060 1184
rect 1564 1156 1572 1164
rect 2748 1156 2756 1164
rect 2860 1156 2868 1164
rect 4140 1156 4148 1164
rect 7932 1156 7940 1164
rect 11292 1156 11300 1164
rect 1836 1136 1844 1144
rect 2140 1136 2148 1144
rect 2428 1136 2436 1144
rect 2796 1136 2804 1144
rect 4316 1136 4324 1144
rect 6044 1136 6052 1144
rect 9052 1136 9060 1144
rect 10332 1136 10340 1144
rect 12284 1136 12292 1144
rect 76 1116 84 1124
rect 140 1116 148 1124
rect 348 1116 356 1124
rect 1548 1116 1556 1124
rect 1804 1116 1812 1124
rect 2220 1116 2228 1124
rect 2748 1116 2756 1124
rect 3372 1116 3380 1124
rect 4924 1116 4932 1124
rect 5116 1116 5124 1124
rect 6524 1116 6532 1124
rect 7676 1116 7684 1124
rect 8300 1116 8308 1124
rect 8588 1116 8596 1124
rect 8668 1116 8676 1124
rect 9356 1116 9364 1124
rect 9724 1116 9732 1124
rect 10924 1116 10932 1124
rect 11180 1116 11188 1124
rect 11196 1116 11204 1124
rect 11788 1116 11796 1124
rect 1564 1096 1572 1104
rect 2188 1102 2196 1104
rect 2188 1096 2196 1102
rect 3196 1096 3204 1104
rect 4076 1096 4084 1104
rect 4140 1102 4148 1104
rect 4140 1096 4148 1102
rect 5596 1096 5604 1104
rect 7404 1096 7412 1104
rect 7788 1096 7796 1104
rect 8444 1096 8452 1104
rect 8460 1096 8468 1104
rect 8684 1102 8692 1104
rect 8684 1096 8692 1102
rect 10332 1096 10340 1104
rect 10428 1096 10436 1104
rect 12284 1096 12292 1104
rect 60 1076 68 1084
rect 3932 1056 3940 1064
rect 11132 1036 11140 1044
rect 460 1016 468 1024
rect 3964 1016 3972 1024
rect 3996 1016 4004 1024
rect 6476 1016 6484 1024
rect 2380 996 2388 1004
rect 3308 996 3316 1004
rect 3324 996 3332 1004
rect 4044 996 4052 1004
rect 10924 996 10932 1004
rect 4524 976 4532 984
rect 7660 976 7668 984
rect 60 956 68 964
rect 1916 956 1924 964
rect 6812 956 6820 964
rect 7660 956 7668 964
rect 9820 956 9828 964
rect 10268 956 10276 964
rect 252 936 260 944
rect 348 936 356 944
rect 7788 936 7796 944
rect 8380 936 8388 944
rect 8700 936 8708 944
rect 11836 936 11844 944
rect 1196 916 1204 924
rect 1292 916 1300 924
rect 2188 916 2196 924
rect 3628 916 3636 924
rect 4540 916 4548 924
rect 5804 916 5812 924
rect 6108 916 6116 924
rect 7100 916 7108 924
rect 8428 916 8436 924
rect 10652 916 10660 924
rect 11884 916 11892 924
rect 11932 918 11940 924
rect 11932 916 11940 918
rect 124 896 132 904
rect 172 896 180 904
rect 892 896 900 904
rect 1548 896 1556 904
rect 1564 896 1572 904
rect 2204 896 2212 904
rect 2732 896 2740 904
rect 3820 896 3828 904
rect 4428 896 4436 904
rect 4524 896 4532 904
rect 4684 896 4692 904
rect 5644 896 5652 904
rect 6092 896 6100 904
rect 6796 896 6804 904
rect 7020 896 7028 904
rect 7084 896 7092 904
rect 7660 896 7668 904
rect 8508 896 8516 904
rect 8716 896 8724 904
rect 9244 896 9252 904
rect 9820 896 9828 904
rect 10556 896 10564 904
rect 11548 896 11556 904
rect 11836 896 11844 904
rect 1276 876 1284 884
rect 1500 876 1508 884
rect 2140 876 2148 884
rect 2796 876 2804 884
rect 4620 876 4628 884
rect 6044 876 6052 884
rect 3788 856 3796 864
rect 11772 856 11780 864
rect 892 836 900 844
rect 3852 836 3860 844
rect 1148 816 1156 824
rect 6412 816 6420 824
rect 844 796 852 804
rect 1500 796 1508 804
rect 11788 796 11796 804
rect 876 776 884 784
rect 9868 776 9876 784
rect 2636 756 2644 764
rect 5292 756 5300 764
rect 7004 756 7012 764
rect 7900 756 7908 764
rect 1900 736 1908 744
rect 2140 736 2148 744
rect 5692 736 5700 744
rect 9036 736 9044 744
rect 10508 736 10516 744
rect 11196 736 11204 744
rect 12284 736 12292 744
rect 140 716 148 724
rect 908 716 916 724
rect 1532 716 1540 724
rect 2172 716 2180 724
rect 2860 716 2868 724
rect 4044 716 4052 724
rect 5660 716 5668 724
rect 6092 716 6100 724
rect 7004 716 7012 724
rect 76 696 84 704
rect 764 696 772 704
rect 876 696 884 704
rect 1500 696 1508 704
rect 1548 702 1556 704
rect 1548 696 1556 702
rect 1836 696 1844 704
rect 2188 702 2196 704
rect 2188 696 2196 702
rect 2572 696 2580 704
rect 3532 696 3540 704
rect 4364 696 4372 704
rect 6028 696 6036 704
rect 6044 702 6052 704
rect 6044 696 6052 702
rect 6524 696 6532 704
rect 6540 696 6548 704
rect 6748 696 6756 704
rect 7404 716 7412 724
rect 10268 716 10276 724
rect 10476 716 10484 724
rect 10524 716 10532 724
rect 10572 716 10580 724
rect 11580 716 11588 724
rect 12076 716 12084 724
rect 9084 696 9092 704
rect 10332 696 10340 704
rect 10428 696 10436 704
rect 12284 696 12292 704
rect 60 656 68 664
rect 9676 656 9684 664
rect 11804 656 11812 664
rect 1260 616 1268 624
rect 2540 616 2548 624
rect 4620 616 4628 624
rect 5132 616 5140 624
rect 9532 616 9540 624
rect 3820 596 3828 604
rect 8316 596 8324 604
rect 4172 576 4180 584
rect 9900 576 9908 584
rect 12476 576 12484 584
rect 60 556 68 564
rect 8428 556 8436 564
rect 12076 556 12084 564
rect 1532 536 1540 544
rect 6124 536 6132 544
rect 204 516 212 524
rect 252 516 260 524
rect 876 516 884 524
rect 1276 516 1284 524
rect 2172 516 2180 524
rect 2236 516 2244 524
rect 2764 516 2772 524
rect 2860 516 2868 524
rect 3836 516 3844 524
rect 1292 496 1300 504
rect 2076 496 2084 504
rect 2204 496 2212 504
rect 2300 496 2308 504
rect 5164 516 5172 524
rect 6076 516 6084 524
rect 6684 516 6692 524
rect 8220 518 8228 524
rect 8220 516 8228 518
rect 9980 518 9988 524
rect 9980 516 9988 518
rect 11068 516 11076 524
rect 11468 516 11476 524
rect 11660 516 11668 524
rect 4172 496 4180 504
rect 5068 496 5076 504
rect 6748 496 6756 504
rect 7644 496 7652 504
rect 8316 496 8324 504
rect 156 476 164 484
rect 2860 476 2868 484
rect 9148 496 9156 504
rect 9660 496 9668 504
rect 9756 496 9764 504
rect 10540 496 10548 504
rect 11628 496 11636 504
rect 11804 496 11812 504
rect 9916 476 9924 484
rect 10476 476 10484 484
rect 12028 476 12036 484
rect 844 456 852 464
rect 8220 456 8228 464
rect 9004 456 9012 464
rect 10540 456 10548 464
rect 5980 436 5988 444
rect 9884 436 9892 444
rect 10428 436 10436 444
rect 2092 416 2100 424
rect 4140 416 4148 424
rect 9052 416 9060 424
rect 5932 376 5940 384
rect 8588 376 8596 384
rect 10556 376 10564 384
rect 764 356 772 364
rect 876 356 884 364
rect 7292 356 7300 364
rect 11020 356 11028 364
rect 1404 336 1412 344
rect 1500 336 1508 344
rect 7388 336 7396 344
rect 76 316 84 324
rect 156 316 164 324
rect 780 316 788 324
rect 892 316 900 324
rect 1580 316 1588 324
rect 2476 316 2484 324
rect 2732 316 2740 324
rect 2876 316 2884 324
rect 3820 316 3828 324
rect 4044 316 4052 324
rect 5932 316 5940 324
rect 5948 316 5956 324
rect 5996 316 6004 324
rect 6044 316 6052 324
rect 6604 316 6612 324
rect 6620 316 6628 324
rect 7948 316 7956 324
rect 764 296 772 304
rect 1548 302 1556 304
rect 1548 296 1556 302
rect 2220 296 2228 304
rect 2940 296 2948 304
rect 4140 302 4148 304
rect 4140 296 4148 302
rect 5180 296 5188 304
rect 5836 296 5844 304
rect 5980 296 5988 304
rect 6588 296 6596 304
rect 6748 296 6756 304
rect 7388 302 7396 304
rect 7388 296 7396 302
rect 8588 316 8596 324
rect 9996 316 10004 324
rect 10572 316 10580 324
rect 11468 316 11476 324
rect 11644 316 11652 324
rect 12028 316 12036 324
rect 11020 296 11028 304
rect 2860 276 2868 284
rect 5964 276 5972 284
rect 60 256 68 264
rect 6636 256 6644 264
rect 11676 256 11684 264
rect 4412 236 4420 244
rect 700 216 708 224
rect 4572 216 4580 224
rect 6588 216 6596 224
rect 9148 216 9156 224
rect 11564 216 11572 224
rect 604 196 612 204
rect 1036 196 1044 204
rect 1276 196 1284 204
rect 3500 196 3508 204
rect 4508 196 4516 204
rect 9852 196 9860 204
rect 11644 196 11652 204
rect 6604 176 6612 184
rect 60 156 68 164
rect 1228 156 1236 164
rect 1980 156 1988 164
rect 2844 156 2852 164
rect 6908 156 6916 164
rect 6924 156 6932 164
rect 8588 156 8596 164
rect 4956 136 4964 144
rect 6092 136 6100 144
rect 8428 136 8436 144
rect 10652 136 10660 144
rect 1276 116 1284 124
rect 1820 116 1828 124
rect 1852 116 1860 124
rect 1900 116 1908 124
rect 1980 116 1988 124
rect 2332 116 2340 124
rect 2940 116 2948 124
rect 4572 116 4580 124
rect 5292 116 5300 124
rect 5948 116 5956 124
rect 6044 116 6052 124
rect 7212 116 7220 124
rect 8924 116 8932 124
rect 9212 116 9220 124
rect 9852 116 9860 124
rect 76 96 84 104
rect 204 96 212 104
rect 1036 96 1044 104
rect 1228 96 1236 104
rect 1836 96 1844 104
rect 2092 96 2100 104
rect 3500 96 3508 104
rect 4412 96 4420 104
rect 4508 96 4516 104
rect 4956 96 4964 104
rect 6924 96 6932 104
rect 7292 96 7300 104
rect 7948 96 7956 104
rect 8588 96 8596 104
rect 9180 96 9188 104
rect 9340 96 9348 104
rect 10668 96 10676 104
rect 12204 96 12212 104
rect 2860 76 2868 84
rect 7004 76 7012 84
rect 1852 36 1860 44
rect 204 16 212 24
rect 764 16 772 24
rect 1756 16 1764 24
rect 1836 16 1844 24
rect 2732 16 2740 24
rect 5980 16 5988 24
rect 6012 16 6020 24
rect 7004 16 7012 24
rect 9212 16 9220 24
rect 9244 16 9252 24
<< metal4 >>
rect 557 8904 563 8936
rect 1165 8904 1171 8936
rect 45 4364 51 8076
rect 61 5704 67 8596
rect 125 8144 131 8536
rect 141 8504 147 8656
rect 77 7124 83 7796
rect 77 6524 83 6716
rect 93 6504 99 6736
rect 61 4424 67 4776
rect 77 4484 83 5296
rect 109 4864 115 7496
rect 125 7084 131 7476
rect 125 6684 131 7076
rect 125 6544 131 6676
rect 157 6524 163 6696
rect 157 6404 163 6516
rect 173 6024 179 7136
rect 205 6064 211 7096
rect 381 6724 387 7716
rect 445 6824 451 7296
rect 381 6204 387 6716
rect 141 5304 147 5396
rect 205 5124 211 5276
rect 413 4724 419 5156
rect 429 4744 435 6096
rect 173 3924 179 4056
rect 61 3804 67 3896
rect 93 3804 99 3916
rect 61 3404 67 3496
rect 93 3404 99 3516
rect 125 3484 131 3876
rect 157 3024 163 3516
rect 77 2524 83 2596
rect 253 2424 259 2496
rect 141 2004 147 2296
rect 157 2044 163 2336
rect 253 2324 259 2356
rect 173 1804 179 2096
rect 429 2044 435 4496
rect 445 4424 451 5916
rect 461 5664 467 7696
rect 493 5644 499 5936
rect 509 4984 515 8896
rect 525 8604 531 8716
rect 1165 8664 1171 8876
rect 1181 8724 1187 8756
rect 557 8324 563 8416
rect 621 8304 627 8356
rect 532 7917 540 7923
rect 573 7704 579 7936
rect 637 7904 643 8476
rect 1037 8084 1043 8496
rect 525 6324 531 6436
rect 541 6404 547 6896
rect 557 6104 563 6136
rect 605 5924 611 6396
rect 605 5624 611 5896
rect 525 5524 531 5556
rect 557 5424 563 5516
rect 605 5464 611 5496
rect 557 4904 563 4936
rect 461 2624 467 4896
rect 621 4764 627 7896
rect 685 7724 691 7736
rect 637 6944 643 7496
rect 701 7404 707 7496
rect 717 7024 723 8076
rect 1101 7804 1107 8316
rect 637 6764 643 6936
rect 477 4124 483 4736
rect 493 4624 499 4736
rect 493 4044 499 4336
rect 557 4324 563 4596
rect 573 4504 579 4536
rect 589 4104 595 4276
rect 621 4084 627 4296
rect 509 3624 515 4076
rect 637 3904 643 6756
rect 733 6164 739 7696
rect 749 7404 755 7516
rect 813 7284 819 7516
rect 1069 6864 1075 7116
rect 749 6324 755 6596
rect 973 5924 979 6076
rect 733 5804 739 5896
rect 749 5824 755 5916
rect 1085 5604 1091 6096
rect 701 5264 707 5496
rect 733 5224 739 5536
rect 1101 5464 1107 5696
rect 749 5204 755 5296
rect 525 3584 531 3696
rect 525 3304 531 3376
rect 557 3304 563 3336
rect 605 2904 611 2956
rect 509 2224 515 2896
rect 525 2724 531 2756
rect 557 2604 563 2716
rect 621 2584 627 2696
rect 557 2104 563 2136
rect 477 1804 483 1936
rect 525 1924 531 1956
rect 77 1124 83 1316
rect 141 1124 147 1196
rect 61 964 67 1076
rect 77 704 83 1116
rect 173 904 179 1296
rect 349 944 355 1116
rect 461 1024 467 1696
rect 477 1684 483 1796
rect 621 1764 627 1896
rect 621 1724 627 1756
rect 637 1604 643 3896
rect 701 2924 707 4756
rect 1117 4524 1123 8196
rect 1149 7444 1155 8476
rect 1181 8103 1187 8676
rect 1277 8404 1283 8696
rect 1293 8624 1299 8916
rect 2509 8904 2515 8936
rect 3181 8904 3187 8956
rect 3245 8924 3251 8976
rect 1876 8897 1884 8903
rect 3780 8897 3788 8903
rect 1421 8844 1427 8896
rect 1812 8717 1820 8723
rect 1172 8097 1187 8103
rect 1277 8004 1283 8376
rect 1293 8004 1299 8036
rect 1165 7924 1171 7956
rect 1229 7304 1235 7356
rect 1293 7324 1299 7376
rect 1133 5844 1139 6336
rect 1133 5524 1139 5536
rect 1149 4784 1155 6896
rect 1165 5384 1171 7296
rect 1181 6704 1187 6716
rect 1277 6704 1283 6716
rect 1245 6504 1251 6556
rect 1181 6424 1187 6496
rect 1277 5324 1283 6696
rect 1293 6524 1299 6576
rect 1293 5824 1299 6296
rect 1213 5104 1219 5116
rect 1197 4904 1203 4976
rect 1245 4904 1251 4956
rect 1165 4724 1171 4836
rect 1245 4524 1251 4536
rect 1165 4324 1171 4336
rect 909 4004 915 4116
rect 1197 4104 1203 4136
rect 1165 4024 1171 4096
rect 909 3724 915 3996
rect 749 2944 755 3236
rect 525 1484 531 1516
rect 157 723 163 896
rect 148 717 163 723
rect 61 564 67 656
rect 77 324 83 696
rect 157 484 163 717
rect 253 524 259 936
rect 157 324 163 476
rect 61 164 67 256
rect 77 104 83 316
rect 205 104 211 516
rect 605 204 611 1476
rect 701 224 707 2916
rect 797 1424 803 3696
rect 1101 3304 1107 3916
rect 1101 2424 1107 2896
rect 1101 1404 1107 1916
rect 1133 1464 1139 3516
rect 1261 3504 1267 5096
rect 1165 3304 1171 3356
rect 1261 3304 1267 3356
rect 1165 2624 1171 2716
rect 717 1204 723 1396
rect 893 1044 899 1296
rect 893 844 899 896
rect 845 724 851 796
rect 877 784 883 836
rect 765 704 771 716
rect 877 704 883 776
rect 765 304 771 356
rect 845 324 851 456
rect 877 364 883 516
rect 893 324 899 836
rect 909 724 915 1196
rect 1149 824 1155 2496
rect 1197 2324 1203 2536
rect 1165 2104 1171 2176
rect 1197 2104 1203 2136
rect 1261 2124 1267 2156
rect 1165 1504 1171 1516
rect 1197 904 1203 916
rect 1261 624 1267 1516
rect 1277 884 1283 5316
rect 1293 4564 1299 5096
rect 1293 3544 1299 4556
rect 1309 4124 1315 4176
rect 1325 3924 1331 8096
rect 1437 7344 1443 7516
rect 1389 7044 1395 7116
rect 1437 6724 1443 6736
rect 1533 6724 1539 8116
rect 1693 7964 1699 8316
rect 1709 7924 1715 8496
rect 1373 4844 1379 4956
rect 1373 4624 1379 4736
rect 1581 4524 1587 4696
rect 1341 3364 1347 4396
rect 1549 3124 1555 3156
rect 1389 3024 1395 3096
rect 1405 2984 1411 3116
rect 1293 2524 1299 2916
rect 1293 1724 1299 2276
rect 1661 1824 1667 7296
rect 1709 7204 1715 7916
rect 1677 5124 1683 5296
rect 1677 3904 1683 4716
rect 1677 3884 1683 3896
rect 1693 3524 1699 5916
rect 1709 5904 1715 6896
rect 1741 6484 1747 6876
rect 1757 6743 1763 7696
rect 1837 7124 1843 7916
rect 1885 7704 1891 7756
rect 1901 7504 1907 8516
rect 2173 8104 2179 8136
rect 2013 7924 2019 7996
rect 1933 7904 1939 7916
rect 1757 6737 1779 6743
rect 1773 6624 1779 6737
rect 1869 6524 1875 6916
rect 1812 6497 1820 6503
rect 1709 5164 1715 5516
rect 1741 5324 1747 6476
rect 1828 5697 1836 5703
rect 1828 5297 1836 5303
rect 1869 5284 1875 6516
rect 1933 6484 1939 7896
rect 2013 7564 2019 7916
rect 2109 7764 2115 7976
rect 2045 6604 2051 6716
rect 1885 6104 1891 6156
rect 1901 5704 1907 6136
rect 1901 5324 1907 5336
rect 1828 5117 1836 5123
rect 1821 4904 1827 4996
rect 1805 4404 1811 4496
rect 1821 4324 1827 4416
rect 1853 4184 1859 4316
rect 1869 4104 1875 5276
rect 1901 4964 1907 5096
rect 1821 3924 1827 3996
rect 1709 2504 1715 3636
rect 1853 3484 1859 3516
rect 1741 3264 1747 3296
rect 1757 2484 1763 2876
rect 1805 2804 1811 2896
rect 1885 2504 1891 4776
rect 1901 2724 1907 3496
rect 1901 2704 1907 2716
rect 1901 2503 1907 2696
rect 1917 2524 1923 6396
rect 2077 6324 2083 7656
rect 2125 6324 2131 7116
rect 2141 6884 2147 6996
rect 2189 6404 2195 8516
rect 2365 8084 2371 8896
rect 3021 8804 3027 8896
rect 3389 8724 3395 8896
rect 2461 8584 2467 8716
rect 2509 8604 2515 8716
rect 2669 8624 2675 8696
rect 2205 7904 2211 7956
rect 2205 6924 2211 7016
rect 2205 6864 2211 6896
rect 2205 6804 2211 6856
rect 1933 6124 1939 6176
rect 1901 2497 1923 2503
rect 1421 1624 1427 1696
rect 1757 1644 1763 2476
rect 1828 2317 1836 2323
rect 1885 2104 1891 2496
rect 1901 2124 1907 2396
rect 1828 2097 1836 2103
rect 1885 1904 1891 2096
rect 1293 924 1299 1576
rect 1437 1484 1443 1516
rect 1501 1324 1507 1436
rect 1533 1204 1539 1316
rect 1277 524 1283 556
rect 205 24 211 96
rect 765 24 771 296
rect 1277 204 1283 516
rect 1293 504 1299 916
rect 1501 804 1507 876
rect 1533 724 1539 1196
rect 1565 1164 1571 1296
rect 1549 904 1555 1116
rect 1565 1104 1571 1156
rect 1805 1124 1811 1476
rect 1837 1144 1843 1496
rect 1549 823 1555 896
rect 1565 844 1571 896
rect 1549 817 1571 823
rect 1501 344 1507 696
rect 1533 524 1539 536
rect 1405 324 1411 336
rect 1549 304 1555 696
rect 1565 564 1571 817
rect 1581 324 1587 1036
rect 1917 964 1923 2497
rect 1933 1364 1939 5896
rect 1949 5484 1955 5496
rect 1965 4304 1971 5716
rect 1981 4424 1987 4756
rect 1997 3884 2003 3896
rect 1949 3324 1955 3356
rect 1981 3264 1987 3356
rect 2013 3264 2019 6316
rect 2061 5924 2067 6216
rect 2077 5224 2083 5316
rect 2061 4704 2067 4716
rect 2045 3364 2051 3696
rect 2061 3324 2067 3716
rect 2093 3524 2099 4476
rect 2093 2904 2099 2996
rect 2029 2084 2035 2296
rect 2109 2064 2115 5916
rect 2125 2864 2131 6316
rect 2365 6104 2371 6476
rect 2381 6444 2387 8316
rect 2509 8204 2515 8316
rect 2445 7697 2460 7703
rect 2413 6504 2419 6696
rect 2189 5904 2195 6036
rect 2189 4724 2195 5696
rect 2349 5304 2355 5516
rect 2333 5204 2339 5296
rect 2189 2744 2195 4716
rect 2317 3904 2323 4076
rect 2189 2324 2195 2736
rect 1949 1884 1955 1936
rect 2141 884 2147 1136
rect 2221 1124 2227 1536
rect 2189 924 2195 1096
rect 2141 744 2147 876
rect 1037 104 1043 196
rect 1229 104 1235 156
rect 1277 124 1283 196
rect 1821 104 1827 116
rect 1837 104 1843 696
rect 1901 124 1907 736
rect 2173 724 2179 796
rect 2173 524 2179 716
rect 2189 704 2195 916
rect 2077 504 2083 516
rect 2205 504 2211 896
rect 2221 524 2227 1116
rect 2237 524 2243 2876
rect 1981 124 1987 156
rect 1757 24 1763 96
rect 1837 24 1843 96
rect 1853 44 1859 116
rect 2093 104 2099 416
rect 2221 304 2227 516
rect 2301 504 2307 2856
rect 2317 1504 2323 3896
rect 2333 3644 2339 5116
rect 2349 3964 2355 5296
rect 2365 3484 2371 6096
rect 2413 6084 2419 6496
rect 2381 4624 2387 4896
rect 2349 2504 2355 2936
rect 2365 1524 2371 1696
rect 2221 104 2227 296
rect 2333 124 2339 1316
rect 2365 1304 2371 1516
rect 2381 1004 2387 1916
rect 2413 1584 2419 6076
rect 2445 4384 2451 7697
rect 2461 7404 2467 7516
rect 2477 7304 2483 7616
rect 2493 6184 2499 7296
rect 2525 6504 2531 8356
rect 2733 8324 2739 8716
rect 2573 8264 2579 8296
rect 2557 7324 2563 8116
rect 2669 8024 2675 8316
rect 2765 8304 2771 8696
rect 2685 8064 2691 8296
rect 2845 8024 2851 8316
rect 3021 7884 3027 8096
rect 2580 7497 2588 7503
rect 2461 5704 2467 5756
rect 2493 5704 2499 6176
rect 2509 6044 2515 6196
rect 2461 5297 2476 5303
rect 2461 5264 2467 5297
rect 2509 4904 2515 4936
rect 2525 4784 2531 6496
rect 2557 6144 2563 7096
rect 2605 6164 2611 7316
rect 2749 6884 2755 6896
rect 2717 6704 2723 6716
rect 2813 6704 2819 7096
rect 2829 6704 2835 7496
rect 3021 7104 3027 7876
rect 3037 7284 3043 8076
rect 3117 7504 3123 8496
rect 3325 8484 3331 8716
rect 3469 8544 3475 8696
rect 3229 7924 3235 7936
rect 3229 7884 3235 7896
rect 3229 7524 3235 7876
rect 3165 7304 3171 7496
rect 3021 6944 3027 7096
rect 2557 5524 2563 6116
rect 2573 6084 2579 6116
rect 2477 4424 2483 4616
rect 2461 4024 2467 4096
rect 2461 3124 2467 3156
rect 2525 2904 2531 3396
rect 2541 3304 2547 3336
rect 2429 2084 2435 2776
rect 2557 2124 2563 5516
rect 2573 5484 2579 6076
rect 2605 5724 2611 6156
rect 2637 6124 2643 6696
rect 2845 6684 2851 6716
rect 2845 6544 2851 6656
rect 3117 6304 3123 7296
rect 2973 6044 2979 6116
rect 2877 5924 2883 5956
rect 2733 5564 2739 5916
rect 2765 5604 2771 5896
rect 3005 5724 3011 6276
rect 3117 6104 3123 6196
rect 2733 5304 2739 5556
rect 2765 5324 2771 5596
rect 2573 5104 2579 5116
rect 2573 3604 2579 5096
rect 2653 4744 2659 5076
rect 2701 4504 2707 4516
rect 2813 4464 2819 5296
rect 2861 4504 2867 5196
rect 2669 3664 2675 3976
rect 2781 3324 2787 3876
rect 2813 3344 2819 4436
rect 2676 3317 2684 3323
rect 2573 3304 2579 3316
rect 2781 3284 2787 3316
rect 2461 2104 2467 2116
rect 2461 1524 2467 1536
rect 2429 1144 2435 1276
rect 2541 1244 2547 2116
rect 2573 2084 2579 3116
rect 2669 2104 2675 2756
rect 2685 1864 2691 3096
rect 2797 2164 2803 2496
rect 2797 2124 2803 2156
rect 2573 1304 2579 1716
rect 2605 1664 2611 1856
rect 2541 624 2547 1236
rect 2573 1044 2579 1296
rect 2637 1284 2643 1676
rect 2740 1517 2748 1523
rect 2573 704 2579 1036
rect 2637 764 2643 1276
rect 2749 1124 2755 1156
rect 2740 897 2748 903
rect 2733 324 2739 796
rect 2765 524 2771 1936
rect 2813 1624 2819 3336
rect 2829 1544 2835 4116
rect 2877 4104 2883 5536
rect 3005 5524 3011 5716
rect 3005 4124 3011 5516
rect 3021 4804 3027 5696
rect 3053 5344 3059 5536
rect 3021 4764 3027 4796
rect 3069 4744 3075 5116
rect 3117 4904 3123 6036
rect 3133 5704 3139 6336
rect 3165 6324 3171 7296
rect 3149 6104 3155 6216
rect 3005 4104 3011 4116
rect 2861 3503 2867 3936
rect 2845 3497 2867 3503
rect 2845 3324 2851 3497
rect 2861 3304 2867 3336
rect 2845 2524 2851 2536
rect 2845 2104 2851 2496
rect 2797 884 2803 1136
rect 2829 804 2835 1496
rect 2468 317 2476 323
rect 2733 24 2739 316
rect 2845 164 2851 2096
rect 2861 1404 2867 3296
rect 2877 2104 2883 4096
rect 3053 2744 3059 2776
rect 3005 2544 3011 2716
rect 3069 2344 3075 4736
rect 3117 4323 3123 4896
rect 3108 4317 3123 4323
rect 2957 2084 2963 2116
rect 3021 1604 3027 1916
rect 2861 1164 2867 1296
rect 2861 724 2867 896
rect 2861 484 2867 516
rect 2877 324 2883 1516
rect 3085 1324 3091 3096
rect 3117 2264 3123 4317
rect 3133 4084 3139 5696
rect 3133 3624 3139 4076
rect 3149 3924 3155 4156
rect 3165 3704 3171 6296
rect 3213 5504 3219 7296
rect 3213 5284 3219 5496
rect 3213 4864 3219 5276
rect 3229 4744 3235 7516
rect 3245 5504 3251 6396
rect 3245 4924 3251 5496
rect 3261 5484 3267 5496
rect 3261 4724 3267 5476
rect 3229 4704 3235 4716
rect 3229 4344 3235 4356
rect 3197 4224 3203 4336
rect 3181 4044 3187 4096
rect 3197 3924 3203 4036
rect 3213 3904 3219 3976
rect 3229 3744 3235 4296
rect 3133 2624 3139 3496
rect 3117 1704 3123 1716
rect 3149 1124 3155 2416
rect 3165 2324 3171 3696
rect 3181 2704 3187 3536
rect 3181 1904 3187 2696
rect 3181 1724 3187 1896
rect 3197 1104 3203 3596
rect 3213 1424 3219 3496
rect 3229 1544 3235 3476
rect 3245 2304 3251 4696
rect 3261 4484 3267 4716
rect 3261 2164 3267 4476
rect 3277 3024 3283 8096
rect 3341 7504 3347 7516
rect 3373 6124 3379 8496
rect 3837 8324 3843 8516
rect 3389 6904 3395 7016
rect 3389 6724 3395 6736
rect 3389 6704 3395 6716
rect 3389 5364 3395 6096
rect 3421 5904 3427 6496
rect 3485 6124 3491 8116
rect 3828 7897 3836 7903
rect 3853 7744 3859 8916
rect 4045 8444 4051 8896
rect 3773 7704 3779 7736
rect 3325 5204 3331 5356
rect 3485 5124 3491 6116
rect 3501 5184 3507 5536
rect 3389 5084 3395 5116
rect 3293 4504 3299 4676
rect 3277 2684 3283 2696
rect 3293 2464 3299 4496
rect 3309 3304 3315 4836
rect 3389 4717 3404 4723
rect 3389 4704 3395 4717
rect 3501 4704 3507 5176
rect 3485 4504 3491 4523
rect 3332 4317 3340 4323
rect 3325 3724 3331 3996
rect 3341 3944 3347 3976
rect 3325 3484 3331 3716
rect 3357 3484 3363 4336
rect 3437 4324 3443 4356
rect 3469 4304 3475 4376
rect 3533 4324 3539 7516
rect 3645 7144 3651 7496
rect 3645 7124 3651 7136
rect 3629 5484 3635 5696
rect 3645 5324 3651 7116
rect 3661 6684 3667 7696
rect 3789 7104 3795 7116
rect 3677 5424 3683 6316
rect 3805 6224 3811 6316
rect 3773 5484 3779 5516
rect 3309 3284 3315 3296
rect 3309 1004 3315 2916
rect 3325 2424 3331 3476
rect 3341 3304 3347 3396
rect 3373 3164 3379 4096
rect 3469 3984 3475 4116
rect 3389 3704 3395 3736
rect 3357 2824 3363 3056
rect 3421 2764 3427 2796
rect 3389 2664 3395 2716
rect 3469 2484 3475 2696
rect 3341 2144 3347 2176
rect 3485 2124 3491 3876
rect 3332 1917 3340 1923
rect 3469 1884 3475 1896
rect 3469 1664 3475 1876
rect 3325 1004 3331 1636
rect 3421 1564 3427 1596
rect 3485 1504 3491 2116
rect 3501 1924 3507 3316
rect 3517 3244 3523 4316
rect 3533 3504 3539 4316
rect 3533 1784 3539 3476
rect 3549 2704 3555 5276
rect 3764 4897 3772 4903
rect 3789 4784 3795 5516
rect 3821 5304 3827 7476
rect 3869 7124 3875 7696
rect 3821 4904 3827 4996
rect 3837 4144 3843 5916
rect 3853 5904 3859 6716
rect 3869 5504 3875 7096
rect 3885 6324 3891 7896
rect 3885 5944 3891 6316
rect 3853 4924 3859 4956
rect 3869 4784 3875 5476
rect 3773 3924 3779 4016
rect 3837 3824 3843 3996
rect 3869 3864 3875 4776
rect 3629 3104 3635 3696
rect 3757 3117 3772 3123
rect 3629 2324 3635 3096
rect 3757 2424 3763 3117
rect 3853 2884 3859 3696
rect 3869 3104 3875 3116
rect 3885 3104 3891 5916
rect 3837 2584 3843 2596
rect 3805 2504 3811 2536
rect 3837 2524 3843 2576
rect 3780 2497 3795 2503
rect 3380 1117 3388 1123
rect 3533 704 3539 1776
rect 3629 1724 3635 2316
rect 3773 2104 3779 2416
rect 3773 1644 3779 1696
rect 3629 924 3635 1596
rect 3773 1264 3779 1296
rect 3629 324 3635 916
rect 3789 864 3795 2497
rect 3885 2324 3891 2856
rect 3805 1704 3811 1976
rect 3805 1304 3811 1336
rect 3821 904 3827 2016
rect 3885 1644 3891 2316
rect 3901 1764 3907 3096
rect 3917 2104 3923 6296
rect 3933 3284 3939 7516
rect 3997 7484 4003 7916
rect 4013 7584 4019 8096
rect 4029 7903 4035 7936
rect 4061 7903 4067 7916
rect 4029 7897 4067 7903
rect 4029 7697 4044 7703
rect 3997 7204 4003 7296
rect 4013 6104 4019 6116
rect 3949 5644 3955 5916
rect 3949 5524 3955 5636
rect 3949 4744 3955 5296
rect 3949 3424 3955 4736
rect 3965 3284 3971 3916
rect 3965 2624 3971 3276
rect 3981 3024 3987 5316
rect 3997 4444 4003 5096
rect 4013 4804 4019 5516
rect 3997 3404 4003 3516
rect 4029 3464 4035 7697
rect 4045 7444 4051 7516
rect 4045 6724 4051 6756
rect 4045 6464 4051 6496
rect 4045 6304 4051 6316
rect 4045 5024 4051 5296
rect 4045 4484 4051 4496
rect 4045 4064 4051 4096
rect 4061 3304 4067 7496
rect 4077 7084 4083 8496
rect 4093 7264 4099 8876
rect 4141 8404 4147 8916
rect 6141 8904 6147 8956
rect 4637 8684 4643 8876
rect 4141 7724 4147 7776
rect 4157 6924 4163 7876
rect 4413 7824 4419 8336
rect 4493 8324 4499 8556
rect 4509 7824 4515 8296
rect 4093 5684 4099 6096
rect 4125 5164 4131 6096
rect 4221 5184 4227 7296
rect 4589 7224 4595 8396
rect 4605 7984 4611 8296
rect 4653 7744 4659 8896
rect 4957 8744 4963 8756
rect 4957 8504 4963 8736
rect 4669 7824 4675 7916
rect 4605 7584 4611 7736
rect 4685 7524 4691 7556
rect 4413 7104 4419 7116
rect 4333 6724 4339 6896
rect 4365 6784 4371 6876
rect 4365 6604 4371 6716
rect 4413 5704 4419 5756
rect 4413 5204 4419 5656
rect 4429 5564 4435 7096
rect 4509 6724 4515 7096
rect 4509 6524 4515 6716
rect 4669 6704 4675 6716
rect 4493 5704 4499 5796
rect 4509 5324 4515 5336
rect 4125 3724 4131 5156
rect 4509 4804 4515 5316
rect 4525 5184 4531 5716
rect 4580 5497 4588 5503
rect 4541 4924 4547 5176
rect 4621 5104 4627 6396
rect 4653 5544 4659 5596
rect 4669 5304 4675 5316
rect 4621 5024 4627 5096
rect 4077 2784 4083 3096
rect 3981 2424 3987 2496
rect 3901 1704 3907 1716
rect 3821 324 3827 596
rect 3837 524 3843 1636
rect 3933 1064 3939 2096
rect 3949 2024 3955 2316
rect 3965 1924 3971 1936
rect 3997 1924 4003 1936
rect 3965 1024 3971 1876
rect 3997 1824 4003 1916
rect 4013 1404 4019 1516
rect 3997 944 4003 1016
rect 3853 844 3859 876
rect 4029 323 4035 1956
rect 4045 1864 4051 1916
rect 4141 1164 4147 4796
rect 4157 4224 4163 4256
rect 4173 3524 4179 4376
rect 4413 4204 4419 4736
rect 4429 4724 4435 4756
rect 4669 4724 4675 5236
rect 4685 5144 4691 5296
rect 4685 5064 4691 5136
rect 4717 4784 4723 8316
rect 4781 8124 4787 8296
rect 4797 7804 4803 7896
rect 4797 7504 4803 7536
rect 4957 7524 4963 7696
rect 4781 6724 4787 6756
rect 4733 6064 4739 6716
rect 4781 5284 4787 5316
rect 4685 4724 4691 4736
rect 4509 4204 4515 4696
rect 4173 3344 4179 3516
rect 4317 3324 4323 3916
rect 4205 2684 4211 3316
rect 4205 2124 4211 2676
rect 4317 2504 4323 2896
rect 4333 1504 4339 3116
rect 4532 2917 4540 2923
rect 4429 2704 4435 2716
rect 4461 2484 4467 2496
rect 4365 1684 4371 2476
rect 4589 2424 4595 3636
rect 4621 2904 4627 3516
rect 4653 3104 4659 3136
rect 4621 2504 4627 2896
rect 4637 2704 4643 2716
rect 4637 2624 4643 2696
rect 4413 2084 4419 2096
rect 4541 1764 4547 2116
rect 4333 1424 4339 1496
rect 4317 1184 4323 1296
rect 4141 1104 4147 1156
rect 4317 1144 4323 1176
rect 4045 724 4051 996
rect 4365 704 4371 1676
rect 4525 904 4531 976
rect 4541 924 4547 1736
rect 4557 1724 4563 1776
rect 4621 1684 4627 2496
rect 4669 2404 4675 4716
rect 4781 4564 4787 5276
rect 4797 5104 4803 5676
rect 4829 5384 4835 6896
rect 4797 4484 4803 4696
rect 4420 897 4428 903
rect 4621 884 4627 1676
rect 4685 1524 4691 3996
rect 4781 3904 4787 3956
rect 4781 2744 4787 3896
rect 4797 3484 4803 3503
rect 4797 3184 4803 3296
rect 4797 2904 4803 3116
rect 4813 2924 4819 5156
rect 4829 4504 4835 4816
rect 4925 4724 4931 4776
rect 4941 4324 4947 6396
rect 5021 6364 5027 6476
rect 4957 4804 4963 6316
rect 5021 5124 5027 6336
rect 5069 6224 5075 8716
rect 5133 8504 5139 8716
rect 5133 8304 5139 8496
rect 5181 8484 5187 8696
rect 5261 8324 5267 8596
rect 5261 8204 5267 8296
rect 5293 8204 5299 8316
rect 5101 7904 5107 8056
rect 5284 7917 5292 7923
rect 5085 7004 5091 7116
rect 5060 5917 5068 5923
rect 5085 4924 5091 5916
rect 5101 5244 5107 7896
rect 5124 7697 5132 7703
rect 5149 5724 5155 5756
rect 5165 5604 5171 6816
rect 5181 6304 5187 6696
rect 5181 5604 5187 6296
rect 5053 4784 5059 4896
rect 5021 4704 5027 4756
rect 4957 4004 4963 4096
rect 5069 4004 5075 4856
rect 5085 4324 5091 4916
rect 5101 3944 5107 4656
rect 4829 3204 4835 3256
rect 4701 2704 4707 2716
rect 4765 2684 4771 2696
rect 4781 1504 4787 2736
rect 4797 2324 4803 2896
rect 4813 2724 4819 2916
rect 4845 2844 4851 3516
rect 4813 2524 4819 2696
rect 4797 2104 4803 2316
rect 4813 1744 4819 2516
rect 4829 1704 4835 2796
rect 4941 2517 4979 2523
rect 4941 2504 4947 2517
rect 4925 2184 4931 2356
rect 4957 2304 4963 2496
rect 4973 2483 4979 2517
rect 5021 2497 5084 2503
rect 4973 2477 4995 2483
rect 4989 2464 4995 2477
rect 5021 2464 5027 2497
rect 4925 1124 4931 2176
rect 4957 2084 4963 2296
rect 4989 2124 4995 2336
rect 5101 2104 5107 3936
rect 5117 3664 5123 4316
rect 5133 2544 5139 4476
rect 5149 4124 5155 4136
rect 5165 4124 5171 5116
rect 5197 4884 5203 5896
rect 5181 4344 5187 4356
rect 5149 4084 5155 4096
rect 5181 4064 5187 4296
rect 5197 4104 5203 4136
rect 5133 2324 5139 2536
rect 5245 2464 5251 7116
rect 5261 6304 5267 6516
rect 5261 6224 5267 6296
rect 5277 5764 5283 7196
rect 5293 6224 5299 6316
rect 5309 5924 5315 6216
rect 5325 5784 5331 8896
rect 5389 7924 5395 8076
rect 5453 7884 5459 7896
rect 5389 7324 5395 7496
rect 5389 7104 5395 7316
rect 5341 6904 5347 6916
rect 5357 6704 5363 6916
rect 5341 6044 5347 6496
rect 5341 5904 5347 5916
rect 5293 5544 5299 5556
rect 5277 3104 5283 4716
rect 5325 4664 5331 4916
rect 5277 2904 5283 3096
rect 5325 2903 5331 3616
rect 5341 2944 5347 5116
rect 5357 4864 5363 6696
rect 5373 4884 5379 5116
rect 5389 4724 5395 7096
rect 5405 6724 5411 6876
rect 5405 5184 5411 6716
rect 5421 6524 5427 6676
rect 5421 5344 5427 6516
rect 5453 5924 5459 6896
rect 5469 5903 5475 6316
rect 5453 5897 5475 5903
rect 5437 5304 5443 5316
rect 5421 5124 5427 5196
rect 5325 2897 5340 2903
rect 5341 2724 5347 2756
rect 5405 2484 5411 3536
rect 5133 1864 5139 2316
rect 5149 2124 5155 2136
rect 5229 1884 5235 1896
rect 5277 1884 5283 2316
rect 5348 2097 5356 2103
rect 5389 2084 5395 2476
rect 5421 1544 5427 4916
rect 5437 4384 5443 5296
rect 5453 5244 5459 5897
rect 5485 5704 5491 8896
rect 5821 8704 5827 8756
rect 5853 8644 5859 8716
rect 6413 8624 6419 9016
rect 6445 8624 6451 9016
rect 6605 8704 6611 8936
rect 7709 8904 7715 8936
rect 7773 8924 7779 8956
rect 8381 8904 8387 8956
rect 6605 8684 6611 8696
rect 5757 8104 5763 8136
rect 5821 7704 5827 7756
rect 5725 7304 5731 7696
rect 5789 7044 5795 7116
rect 5837 6924 5843 8496
rect 5997 8484 6003 8496
rect 5988 8317 5996 8323
rect 5453 4504 5459 4556
rect 5469 4224 5475 5696
rect 5485 4904 5491 4916
rect 5501 4624 5507 6716
rect 5757 6104 5763 6156
rect 5661 5444 5667 5516
rect 5453 3924 5459 4016
rect 5645 3924 5651 4316
rect 5645 3744 5651 3916
rect 5693 3524 5699 5676
rect 5805 5204 5811 5716
rect 5821 5424 5827 5496
rect 5805 5104 5811 5176
rect 5821 4704 5827 5236
rect 5837 5184 5843 6896
rect 6013 6464 6019 8476
rect 5949 5904 5955 6156
rect 5997 5684 6003 5696
rect 5853 5104 5859 5196
rect 5805 4284 5811 4296
rect 5805 3724 5811 4096
rect 5805 3704 5811 3716
rect 5789 3664 5795 3676
rect 5437 2704 5443 2856
rect 5645 1924 5651 2596
rect 5693 2304 5699 3516
rect 5421 1404 5427 1536
rect 5165 1304 5171 1396
rect 5053 1184 5059 1296
rect 5124 1117 5132 1123
rect 5604 1097 5612 1103
rect 4685 884 4691 896
rect 4621 624 4627 876
rect 4173 504 4179 576
rect 5069 504 5075 536
rect 4029 317 4044 323
rect 4141 304 4147 416
rect 5133 344 5139 616
rect 5165 464 5171 516
rect 5181 304 5187 1096
rect 5645 904 5651 1916
rect 2861 84 2867 276
rect 2941 124 2947 296
rect 3501 104 3507 196
rect 4413 104 4419 236
rect 4509 104 4515 196
rect 4573 124 4579 216
rect 4957 104 4963 136
rect 5293 124 5299 756
rect 5693 744 5699 2296
rect 5773 1964 5779 2596
rect 5789 2044 5795 2136
rect 5805 1724 5811 2556
rect 5805 924 5811 1716
rect 5821 1324 5827 4356
rect 5917 4124 5923 4816
rect 5837 1284 5843 3556
rect 5853 2524 5859 3656
rect 5885 2864 5891 4076
rect 5917 2744 5923 4116
rect 5949 3804 5955 5176
rect 5988 4717 5996 4723
rect 6013 4504 6019 6316
rect 5949 3724 5955 3796
rect 5917 2624 5923 2736
rect 5997 2544 6003 2896
rect 6029 2864 6035 8516
rect 6045 6484 6051 7936
rect 6093 7924 6099 8536
rect 6628 8317 6636 8323
rect 6429 8104 6435 8156
rect 6061 7364 6067 7536
rect 6077 7324 6083 7496
rect 6093 6544 6099 7876
rect 6109 6504 6115 7556
rect 6045 2824 6051 6456
rect 6061 5684 6067 6076
rect 6093 5844 6099 5896
rect 6061 3944 6067 5676
rect 6269 5524 6275 7296
rect 6285 5444 6291 8096
rect 6365 7704 6371 7716
rect 6397 7704 6403 7716
rect 6461 7524 6467 7576
rect 6413 7304 6419 7396
rect 6461 7324 6467 7396
rect 6573 6844 6579 7116
rect 6301 6204 6307 6716
rect 6589 6544 6595 8316
rect 6605 7924 6611 7936
rect 6605 7304 6611 7696
rect 6605 6844 6611 7096
rect 6413 6104 6419 6396
rect 6429 6384 6435 6536
rect 6621 6504 6627 8296
rect 6701 7684 6707 8496
rect 6749 8004 6755 8876
rect 6637 6504 6643 6516
rect 6461 6124 6467 6396
rect 6077 5324 6083 5416
rect 6317 5404 6323 5516
rect 6061 3544 6067 3936
rect 6093 3524 6099 3956
rect 6125 3704 6131 3916
rect 6125 3464 6131 3696
rect 5885 2324 5891 2336
rect 5853 1984 5859 2296
rect 5933 2024 5939 2316
rect 5965 1684 5971 1696
rect 5917 1304 5923 1416
rect 5933 1324 5939 1416
rect 5997 1264 6003 1296
rect 6045 1144 6051 1636
rect 5661 544 5667 716
rect 6029 704 6035 736
rect 6045 704 6051 876
rect 5661 364 5667 536
rect 6045 444 6051 696
rect 6077 524 6083 3156
rect 6109 2324 6115 2636
rect 6125 2524 6131 3456
rect 6125 1704 6131 2516
rect 6141 2104 6147 5296
rect 6237 4104 6243 4316
rect 6237 3164 6243 4096
rect 6269 3124 6275 3696
rect 6333 3444 6339 3896
rect 6269 2064 6275 2716
rect 6285 2044 6291 3296
rect 6349 2704 6355 4316
rect 6365 3784 6371 6096
rect 6477 6064 6483 6356
rect 6381 5524 6387 5556
rect 6413 5424 6419 5516
rect 6477 5464 6483 5496
rect 6381 4504 6387 4776
rect 6413 4104 6419 5276
rect 6429 4524 6435 4596
rect 6429 4324 6435 4476
rect 6429 4204 6435 4316
rect 6413 3824 6419 4096
rect 6429 3304 6435 3356
rect 6381 3084 6387 3116
rect 6429 3104 6435 3116
rect 6100 917 6108 923
rect 6093 724 6099 896
rect 6077 504 6083 516
rect 6093 444 6099 716
rect 6125 544 6131 1696
rect 6301 1644 6307 2096
rect 6349 1444 6355 2496
rect 6429 2484 6435 3096
rect 6429 2304 6435 2476
rect 6413 2104 6419 2136
rect 6381 1524 6387 1996
rect 6365 1484 6371 1516
rect 6413 824 6419 2076
rect 6429 1224 6435 2296
rect 6445 1824 6451 5116
rect 6461 5104 6467 5116
rect 6461 4944 6467 5096
rect 6461 4504 6467 4596
rect 6461 3984 6467 4116
rect 6461 3824 6467 3976
rect 6493 2804 6499 3896
rect 6509 3684 6515 6096
rect 6573 4704 6579 6116
rect 6605 5824 6611 5916
rect 6605 5104 6611 5116
rect 6637 4504 6643 4956
rect 6653 4324 6659 7296
rect 6733 6924 6739 6936
rect 6669 5684 6675 6896
rect 6701 6524 6707 6536
rect 6685 6104 6691 6136
rect 6701 5544 6707 6476
rect 6701 5104 6707 5536
rect 6621 3924 6627 4096
rect 6637 4084 6643 4316
rect 6621 3144 6627 3916
rect 6637 3524 6643 3756
rect 6717 3724 6723 4076
rect 6733 3964 6739 6916
rect 6749 6104 6755 7916
rect 6765 7724 6771 7736
rect 6765 7324 6771 7716
rect 6909 7604 6915 8716
rect 6941 7404 6947 8096
rect 7037 7424 7043 7516
rect 6765 6144 6771 7316
rect 6749 5124 6755 6096
rect 6781 5344 6787 6496
rect 6781 5124 6787 5296
rect 6749 5084 6755 5096
rect 6749 3704 6755 4796
rect 6765 4384 6771 4516
rect 6781 4384 6787 5116
rect 6765 4304 6771 4356
rect 6797 3624 6803 5916
rect 6909 5524 6915 5836
rect 6957 4044 6963 5696
rect 6989 4844 6995 7116
rect 7005 6364 7011 6716
rect 7021 6324 7027 6396
rect 7053 5483 7059 7836
rect 7085 7124 7091 8336
rect 7069 6224 7075 6316
rect 7085 5644 7091 7116
rect 7133 7104 7139 8536
rect 7277 8504 7283 8736
rect 7405 8544 7411 8696
rect 7261 8104 7267 8416
rect 7149 7504 7155 7576
rect 7197 7564 7203 7576
rect 7101 6184 7107 6296
rect 7101 5704 7107 5756
rect 7117 5744 7123 7096
rect 7133 6544 7139 6696
rect 7037 5477 7059 5483
rect 6621 3124 6627 3136
rect 6589 3024 6595 3096
rect 6589 2864 6595 3016
rect 6605 2464 6611 3116
rect 6621 3064 6627 3116
rect 6637 2504 6643 3116
rect 6749 2524 6755 3556
rect 6781 3164 6787 3616
rect 6605 2324 6611 2456
rect 6493 2124 6499 2176
rect 6605 2004 6611 2316
rect 6637 2304 6643 2316
rect 6909 2104 6915 2776
rect 6925 2524 6931 2876
rect 6957 2804 6963 2896
rect 6445 1544 6451 1816
rect 6525 1224 6531 1916
rect 6477 1024 6483 1096
rect 6525 704 6531 1116
rect 6541 704 6547 1436
rect 6573 1284 6579 1896
rect 6605 1264 6611 1996
rect 6637 1924 6643 1956
rect 6637 1704 6643 1736
rect 6733 1724 6739 1776
rect 7005 1424 7011 5316
rect 7037 5304 7043 5477
rect 7037 4624 7043 4716
rect 7069 4264 7075 5196
rect 7085 4724 7091 4756
rect 7085 4264 7091 4276
rect 7101 4124 7107 4276
rect 7101 4064 7107 4076
rect 7117 4024 7123 5176
rect 7133 4804 7139 6536
rect 7277 6164 7283 8096
rect 7293 7664 7299 7696
rect 7293 6724 7299 7116
rect 7357 6344 7363 6836
rect 7373 6304 7379 6836
rect 7389 6804 7395 6896
rect 7389 6604 7395 6716
rect 7405 6404 7411 8496
rect 7613 8124 7619 8556
rect 7661 8304 7667 8316
rect 7661 7924 7667 8116
rect 7517 7304 7523 7636
rect 7220 5317 7228 5323
rect 7389 4924 7395 5116
rect 7213 4744 7219 4756
rect 7293 4324 7299 4356
rect 7373 4144 7379 4296
rect 7293 4084 7299 4096
rect 7293 3924 7299 4056
rect 7309 4044 7315 4076
rect 7373 3684 7379 4136
rect 7389 3904 7395 4796
rect 7405 4784 7411 4916
rect 7405 4624 7411 4736
rect 7421 4324 7427 5296
rect 7421 4284 7427 4316
rect 7389 3724 7395 3856
rect 7069 3304 7075 3576
rect 7389 3544 7395 3696
rect 7092 3317 7100 3323
rect 7085 2904 7091 2936
rect 7117 2924 7123 3436
rect 7149 3144 7155 3436
rect 7220 2917 7228 2923
rect 7021 2684 7027 2716
rect 6973 1324 6979 1396
rect 5933 324 5939 376
rect 5956 317 5964 323
rect 5981 304 5987 436
rect 5997 324 6003 356
rect 5828 297 5836 303
rect 5981 24 5987 296
rect 6013 24 6019 316
rect 6045 124 6051 316
rect 6093 144 6099 436
rect 6621 324 6627 336
rect 6589 224 6595 296
rect 6605 184 6611 316
rect 6637 264 6643 1296
rect 6813 944 6819 956
rect 6797 904 6803 936
rect 7085 904 7091 1556
rect 7101 924 7107 2356
rect 7149 2124 7155 2156
rect 7197 2004 7203 2116
rect 7005 724 7011 756
rect 6685 444 6691 516
rect 6749 504 6755 696
rect 6685 144 6691 436
rect 6909 164 6915 396
rect 6045 104 6051 116
rect 6925 104 6931 156
rect 7005 84 7011 716
rect 7213 124 7219 2516
rect 7389 1904 7395 3496
rect 7421 3324 7427 4276
rect 7437 3524 7443 4776
rect 7453 2864 7459 5916
rect 7300 1297 7308 1303
rect 7293 104 7299 356
rect 7389 344 7395 1896
rect 7517 1844 7523 5496
rect 7533 4844 7539 4856
rect 7533 2504 7539 4836
rect 7581 3324 7587 6316
rect 7645 6124 7651 6136
rect 7661 5704 7667 6816
rect 7597 4123 7603 4896
rect 7645 4524 7651 4996
rect 7597 4117 7619 4123
rect 7613 4044 7619 4117
rect 7533 2344 7539 2496
rect 7421 1404 7427 1696
rect 7581 1604 7587 2736
rect 7645 1984 7651 2096
rect 7405 1104 7411 1316
rect 7405 404 7411 716
rect 7565 504 7571 1076
rect 7661 984 7667 5516
rect 7677 5184 7683 8716
rect 7773 8304 7779 8376
rect 7789 8324 7795 8696
rect 7741 7904 7747 8276
rect 7949 8244 7955 8716
rect 8045 8704 8051 8756
rect 8253 8424 8259 8896
rect 8381 8504 8387 8556
rect 8397 8504 8403 8596
rect 8413 8544 8419 8596
rect 8429 8584 8435 8796
rect 8429 8524 8435 8576
rect 8340 8317 8348 8323
rect 7901 7924 7907 7936
rect 7693 7144 7699 7676
rect 7757 7504 7763 7896
rect 7805 7844 7811 7896
rect 7885 7724 7891 7916
rect 7949 7904 7955 7916
rect 7965 7524 7971 7556
rect 7917 7504 7923 7516
rect 7693 6104 7699 7136
rect 7709 6504 7715 6536
rect 7773 6524 7779 6556
rect 7677 1124 7683 4736
rect 7693 3164 7699 6096
rect 7725 4904 7731 4996
rect 7741 4744 7747 5016
rect 7709 4564 7715 4716
rect 7757 4524 7763 5336
rect 7773 4924 7779 4956
rect 7789 4804 7795 6116
rect 7805 5524 7811 6056
rect 7837 5564 7843 5936
rect 7828 5497 7836 5503
rect 7901 4864 7907 5896
rect 7773 4604 7779 4696
rect 7709 3444 7715 3576
rect 7757 3504 7763 4516
rect 7773 3824 7779 4316
rect 7853 4304 7859 4316
rect 7885 4284 7891 4296
rect 7693 1664 7699 2496
rect 7709 1424 7715 1516
rect 7757 1504 7763 3476
rect 7773 2944 7779 3816
rect 7805 3124 7811 4016
rect 7901 3664 7907 3676
rect 7773 2924 7779 2936
rect 7773 1704 7779 2736
rect 7789 2364 7795 2696
rect 7805 2124 7811 2316
rect 7828 2117 7836 2123
rect 7853 1684 7859 2356
rect 7773 1284 7779 1496
rect 7661 904 7667 956
rect 7789 944 7795 1096
rect 7901 764 7907 3656
rect 7917 2424 7923 7296
rect 7933 3964 7939 7516
rect 7981 6984 7987 8096
rect 8013 7504 8019 7936
rect 8077 7924 8083 8136
rect 8221 8104 8227 8316
rect 8269 7944 8275 8316
rect 8061 7524 8067 7876
rect 8397 7824 8403 7936
rect 8429 7764 8435 8296
rect 8525 7743 8531 8316
rect 8509 7737 8531 7743
rect 8029 7204 8035 7316
rect 7949 5704 7955 5736
rect 8013 5684 8019 6516
rect 8061 6364 8067 6716
rect 8029 5704 8035 5723
rect 7949 5164 7955 5516
rect 8013 5244 8019 5536
rect 8077 5204 8083 5736
rect 7956 5117 7964 5123
rect 7949 4304 7955 4316
rect 7949 4104 7955 4116
rect 7949 3524 7955 3956
rect 7965 2964 7971 4896
rect 8093 4884 8099 7696
rect 8509 7644 8515 7737
rect 8317 6804 8323 6896
rect 8221 6524 8227 6536
rect 8317 6324 8323 6356
rect 8253 6064 8259 6096
rect 8333 5904 8339 7116
rect 8317 5524 8323 5896
rect 8349 5504 8355 6496
rect 8365 6104 8371 6196
rect 8269 5284 8275 5436
rect 8397 4944 8403 4956
rect 8413 4904 8419 7196
rect 8445 7104 8451 7336
rect 8557 7264 8563 8316
rect 8589 8104 8595 8116
rect 8429 6124 8435 6176
rect 8429 5324 8435 5476
rect 8445 5164 8451 7096
rect 8516 6717 8524 6723
rect 8468 6697 8476 6703
rect 8477 6064 8483 6336
rect 8557 5864 8563 6296
rect 8557 5744 8563 5856
rect 7997 3064 8003 3296
rect 8013 2724 8019 3136
rect 8029 3084 8035 4796
rect 8301 4244 8307 4496
rect 8317 4424 8323 4736
rect 8445 4704 8451 5156
rect 8525 4904 8531 4996
rect 8573 4984 8579 7696
rect 8596 6897 8604 6903
rect 8589 6104 8595 6116
rect 8653 5944 8659 8076
rect 8685 7484 8691 8096
rect 8845 8044 8851 8496
rect 8861 8464 8867 8716
rect 8909 8224 8915 8896
rect 9293 8744 9299 8876
rect 9341 8724 9347 8916
rect 9892 8897 9900 8903
rect 9613 8724 9619 8736
rect 8957 8264 8963 8476
rect 9053 8244 9059 8516
rect 9188 8497 9196 8503
rect 9252 8497 9260 8503
rect 9789 8484 9795 8716
rect 9821 8484 9827 8736
rect 9325 8124 9331 8316
rect 9245 8044 9251 8096
rect 9325 7944 9331 8116
rect 8669 6944 8675 7096
rect 8669 6544 8675 6936
rect 8701 6724 8707 7476
rect 8701 6104 8707 6716
rect 8596 5697 8604 5703
rect 8653 4824 8659 5936
rect 8589 4724 8595 4736
rect 8365 4504 8371 4596
rect 8445 4444 8451 4676
rect 8557 4524 8563 4536
rect 8669 4524 8675 5076
rect 8701 4964 8707 5516
rect 8045 3984 8051 4116
rect 8317 3924 8323 3956
rect 8509 3784 8515 4116
rect 8580 4097 8588 4103
rect 8525 3864 8531 3936
rect 8541 3824 8547 4076
rect 8621 3724 8627 3736
rect 8637 3564 8643 3736
rect 8589 3464 8595 3516
rect 7997 2344 8003 2496
rect 8013 2304 8019 2316
rect 7949 1704 7955 1836
rect 8029 1344 8035 3076
rect 8045 2944 8051 3116
rect 8541 3084 8547 3116
rect 8541 3044 8547 3076
rect 8589 2904 8595 2936
rect 8532 2897 8540 2903
rect 8061 1484 8067 2096
rect 8125 1564 8131 2736
rect 8221 2684 8227 2896
rect 8317 2604 8323 2716
rect 8365 2564 8371 2676
rect 8429 2524 8435 2556
rect 8429 2384 8435 2476
rect 8221 1504 8227 1516
rect 7933 1164 7939 1296
rect 8301 1124 8307 2036
rect 8317 1924 8323 1956
rect 8381 1824 8387 1916
rect 8429 924 8435 2376
rect 8445 1104 8451 2716
rect 8621 2503 8627 2536
rect 8580 2497 8627 2503
rect 8596 2317 8604 2323
rect 8637 2144 8643 3556
rect 8637 2084 8643 2136
rect 8669 1924 8675 4516
rect 8685 3904 8691 4676
rect 8685 3744 8691 3876
rect 8701 3764 8707 4236
rect 8733 4024 8739 7116
rect 8829 6504 8835 7516
rect 8829 5504 8835 6496
rect 8861 5524 8867 6496
rect 8749 4544 8755 4556
rect 8861 4144 8867 5176
rect 8877 4224 8883 5116
rect 8461 1304 8467 1656
rect 8669 1504 8675 1916
rect 8669 1124 8675 1496
rect 8468 1097 8476 1103
rect 8589 1084 8595 1116
rect 8685 1104 8691 2896
rect 8701 2544 8707 3736
rect 8733 3704 8739 3756
rect 8733 2644 8739 3116
rect 8909 2404 8915 7916
rect 9005 7824 9011 7916
rect 9069 7864 9075 7896
rect 9229 7683 9235 7916
rect 9252 7697 9260 7703
rect 9229 7677 9251 7683
rect 8989 7504 8995 7516
rect 9037 7504 9043 7516
rect 9213 7304 9219 7376
rect 9229 7324 9235 7416
rect 9245 7384 9251 7677
rect 9053 6504 9059 6556
rect 8973 5904 8979 5916
rect 8973 5264 8979 5296
rect 8989 4324 8995 5376
rect 9021 5304 9027 5556
rect 9005 5124 9011 5196
rect 9021 4504 9027 4636
rect 9053 4384 9059 6296
rect 9277 6164 9283 7916
rect 9325 7324 9331 7896
rect 9341 7204 9347 7516
rect 9357 7504 9363 7896
rect 9741 7804 9747 7896
rect 9357 7124 9363 7396
rect 9373 7164 9379 7296
rect 9357 6944 9363 7016
rect 9373 6904 9379 7156
rect 9325 5724 9331 5916
rect 9245 5704 9251 5716
rect 9069 5324 9075 5596
rect 9236 5517 9244 5523
rect 8973 3924 8979 4136
rect 9181 4104 9187 5316
rect 9309 4904 9315 5236
rect 9245 4704 9251 4716
rect 9325 4704 9331 5716
rect 8973 2624 8979 2716
rect 8701 944 8707 2116
rect 8989 1924 8995 3616
rect 9021 3384 9027 3556
rect 9021 3304 9027 3356
rect 9053 3024 9059 4016
rect 9069 3524 9075 3536
rect 9053 2784 9059 2796
rect 9053 2264 9059 2776
rect 9005 1704 9011 1916
rect 9053 1724 9059 1896
rect 8973 1664 8979 1696
rect 9005 1684 9011 1696
rect 8717 904 8723 1236
rect 8516 897 8524 903
rect 7652 497 7660 503
rect 8221 464 8227 516
rect 8317 504 8323 596
rect 7389 304 7395 336
rect 7949 284 7955 316
rect 8429 144 8435 556
rect 9005 464 9011 1676
rect 9053 1504 9059 1716
rect 9053 1144 9059 1476
rect 9069 1324 9075 3496
rect 9037 724 9043 736
rect 9053 424 9059 1116
rect 9069 524 9075 1316
rect 9085 704 9091 3896
rect 9197 3824 9203 3916
rect 9277 3484 9283 3516
rect 9245 3124 9251 3136
rect 9325 3124 9331 4676
rect 9341 3504 9347 6536
rect 9357 6304 9363 6716
rect 9533 6344 9539 6496
rect 9357 5504 9363 5876
rect 9341 3104 9347 3136
rect 9188 2897 9196 2903
rect 9117 2504 9123 2516
rect 9197 2504 9203 2516
rect 9252 2317 9260 2323
rect 9341 2124 9347 3096
rect 9373 2924 9379 4376
rect 9373 2504 9379 2916
rect 9252 2097 9260 2103
rect 9197 1924 9203 1936
rect 9124 1897 9132 1903
rect 9245 1704 9251 1756
rect 9197 1304 9203 1496
rect 9325 1324 9331 1536
rect 9245 1304 9251 1316
rect 9213 1284 9219 1296
rect 9245 904 9251 1196
rect 8589 324 8595 376
rect 9149 224 9155 496
rect 7949 104 7955 116
rect 8589 104 8595 156
rect 8925 124 8931 136
rect 9188 97 9196 103
rect 7005 24 7011 76
rect 9213 24 9219 116
rect 9341 104 9347 1336
rect 9389 1304 9395 3156
rect 9517 2724 9523 3196
rect 9533 1324 9539 6336
rect 9613 6104 9619 7796
rect 9853 6904 9859 7516
rect 9828 6697 9836 6703
rect 9741 6524 9747 6676
rect 9853 6484 9859 6796
rect 9876 6317 9884 6323
rect 9725 6184 9731 6296
rect 9725 6124 9731 6176
rect 9789 6084 9795 6096
rect 9901 6024 9907 8496
rect 9997 7924 10003 8236
rect 9965 7504 9971 7536
rect 9981 7504 9987 7736
rect 9997 7724 10003 7736
rect 9981 6924 9987 7496
rect 10013 6624 10019 6676
rect 9853 5924 9859 5936
rect 9892 5917 9900 5923
rect 9645 5304 9651 5396
rect 9677 5304 9683 5356
rect 9709 5104 9715 5896
rect 9725 5884 9731 5896
rect 9565 3284 9571 3436
rect 9581 2304 9587 4936
rect 9789 4864 9795 5236
rect 9885 4904 9891 4916
rect 9597 4204 9603 4316
rect 9629 3704 9635 3916
rect 9693 3304 9699 4596
rect 9709 4504 9715 4616
rect 9725 4504 9731 4556
rect 9741 3724 9747 4516
rect 9709 3344 9715 3456
rect 9709 3324 9715 3336
rect 9661 2604 9667 2716
rect 9709 2584 9715 2696
rect 9645 1524 9651 1616
rect 9725 1584 9731 3716
rect 9837 3684 9843 3896
rect 9357 1124 9363 1256
rect 9533 624 9539 1316
rect 9661 504 9667 1516
rect 9725 1124 9731 1576
rect 9677 664 9683 676
rect 9757 504 9763 3536
rect 9821 3124 9827 3356
rect 9853 3344 9859 3716
rect 9885 3704 9891 3716
rect 9869 3684 9875 3696
rect 9789 1904 9795 2956
rect 9821 2524 9827 3036
rect 9821 2484 9827 2516
rect 9853 1924 9859 2996
rect 9885 2884 9891 2896
rect 9885 2464 9891 2496
rect 9885 2104 9891 2436
rect 9821 904 9827 956
rect 9869 784 9875 1916
rect 9885 444 9891 2096
rect 9901 584 9907 5696
rect 9981 4884 9987 5896
rect 10109 5464 10115 8316
rect 10253 8004 10259 8356
rect 10125 7024 10131 7296
rect 10141 5124 10147 6896
rect 10157 5924 10163 6496
rect 9981 4504 9987 4876
rect 9917 4084 9923 4096
rect 9917 3284 9923 3296
rect 9933 3144 9939 4076
rect 9997 3544 10003 3896
rect 9917 484 9923 2716
rect 9981 2364 9987 2696
rect 9981 2164 9987 2356
rect 9981 524 9987 2136
rect 9997 1504 10003 3536
rect 9997 1304 10003 1496
rect 10029 1304 10035 4416
rect 10141 2124 10147 5116
rect 10157 4664 10163 5516
rect 10173 5144 10179 6696
rect 10221 5304 10227 7696
rect 10269 6824 10275 8716
rect 10317 8624 10323 9016
rect 10349 8624 10355 9016
rect 10637 8764 10643 8916
rect 10381 8084 10387 8296
rect 10397 8264 10403 8296
rect 10532 8097 10540 8103
rect 10285 7864 10291 8076
rect 10420 7497 10428 7503
rect 10349 7304 10355 7396
rect 10349 7284 10355 7296
rect 10317 6644 10323 6916
rect 10333 6544 10339 7136
rect 10340 6517 10348 6523
rect 10324 6497 10332 6503
rect 10349 5784 10355 6136
rect 10349 5604 10355 5756
rect 10333 5524 10339 5536
rect 10365 5324 10371 6676
rect 10381 6144 10387 6576
rect 10381 5924 10387 6116
rect 10269 4904 10275 5296
rect 10269 4744 10275 4896
rect 10269 4604 10275 4716
rect 10349 4524 10355 4536
rect 10260 4317 10268 4323
rect 10317 4204 10323 4316
rect 10340 4297 10348 4303
rect 10276 3917 10284 3923
rect 10317 3404 10323 3516
rect 10349 2744 10355 3516
rect 10381 3504 10387 5916
rect 10397 5344 10403 5496
rect 10397 4264 10403 5336
rect 10317 2204 10323 2316
rect 10141 2104 10147 2116
rect 10349 2064 10355 2736
rect 10397 2704 10403 3496
rect 10413 3104 10419 3796
rect 10429 3104 10435 4116
rect 10445 3524 10451 5696
rect 10468 4497 10476 4503
rect 10493 4324 10499 7356
rect 10548 7297 10556 7303
rect 10541 6724 10547 6736
rect 10532 6097 10540 6103
rect 10509 5544 10515 6096
rect 10541 5904 10547 5916
rect 10532 5517 10540 5523
rect 10525 5304 10531 5496
rect 10477 4184 10483 4316
rect 10493 4224 10499 4296
rect 10493 3184 10499 3796
rect 10381 2184 10387 2296
rect 10429 2004 10435 3096
rect 10260 1697 10268 1703
rect 9997 324 10003 1296
rect 10333 1104 10339 1136
rect 10429 1104 10435 1996
rect 10493 1604 10499 1936
rect 10269 724 10275 956
rect 10509 744 10515 5096
rect 10525 2444 10531 5296
rect 10541 5084 10547 5116
rect 10573 5084 10579 5096
rect 10541 4904 10547 4936
rect 10573 4304 10579 4496
rect 10621 4364 10627 8516
rect 10637 7124 10643 8036
rect 10653 7744 10659 8136
rect 10637 6704 10643 6916
rect 10637 5904 10643 6116
rect 10637 4904 10643 5896
rect 10653 5724 10659 7736
rect 10669 5924 10675 8316
rect 10685 7724 10691 7976
rect 10685 6804 10691 7696
rect 10701 6824 10707 8496
rect 10861 7824 10867 8716
rect 10877 8464 10883 8736
rect 11005 8384 11011 8696
rect 10877 7944 10883 8036
rect 10925 7844 10931 7916
rect 11076 7897 11084 7903
rect 10989 7564 10995 7896
rect 11165 7664 11171 8496
rect 10557 2904 10563 4256
rect 10589 2744 10595 3636
rect 10605 3144 10611 3516
rect 10637 3124 10643 4896
rect 10653 4124 10659 5716
rect 10685 5124 10691 5296
rect 10717 4824 10723 7516
rect 11101 7404 11107 7496
rect 10749 6724 10755 6876
rect 10749 5704 10755 6716
rect 10861 4744 10867 4836
rect 10685 4324 10691 4436
rect 10797 4104 10803 4316
rect 10637 2724 10643 3116
rect 10653 2544 10659 3476
rect 10637 1504 10643 2136
rect 10653 1324 10659 2536
rect 10685 2523 10691 4016
rect 10797 2804 10803 4096
rect 10845 3864 10851 4716
rect 10669 2517 10691 2523
rect 10532 717 10540 723
rect 10333 684 10339 696
rect 10429 444 10435 696
rect 10477 484 10483 716
rect 10541 464 10547 496
rect 10557 384 10563 896
rect 10573 324 10579 716
rect 9853 124 9859 196
rect 10653 144 10659 916
rect 10669 104 10675 2517
rect 10685 2104 10691 2496
rect 10909 1704 10915 7236
rect 11117 7124 11123 7516
rect 11149 7404 11155 7516
rect 11181 7464 11187 8716
rect 11197 8404 11203 8896
rect 11293 8704 11299 8756
rect 11821 8564 11827 8716
rect 11949 8624 11955 8696
rect 11293 7984 11299 8316
rect 11645 8204 11651 8316
rect 11789 8224 11795 8496
rect 11197 7524 11203 7536
rect 11197 6884 11203 6896
rect 10957 6504 10963 6536
rect 10925 5584 10931 6496
rect 11181 6064 11187 6096
rect 11140 5917 11148 5923
rect 11133 5104 11139 5396
rect 10973 3704 10979 4736
rect 11005 3944 11011 4156
rect 10957 3304 10963 3356
rect 11005 2524 11011 2716
rect 10932 2497 10940 2503
rect 10925 1784 10931 2316
rect 10941 1924 10947 1956
rect 11005 1644 11011 1896
rect 11021 1744 11027 4116
rect 11053 3924 11059 4176
rect 11085 4124 11091 4136
rect 11085 4024 11091 4036
rect 11101 3904 11107 4136
rect 11053 3244 11059 3316
rect 11085 3104 11091 3496
rect 11085 2924 11091 2936
rect 11101 2904 11107 3616
rect 11117 3504 11123 4696
rect 11197 4504 11203 6516
rect 11181 3524 11187 3536
rect 11197 3264 11203 3696
rect 11197 3164 11203 3196
rect 11197 3124 11203 3156
rect 11037 2324 11043 2556
rect 11085 2524 11091 2536
rect 11188 2497 11196 2503
rect 11197 1924 11203 1936
rect 11037 1724 11043 1756
rect 10925 1524 10931 1636
rect 11133 1524 11139 1536
rect 11076 1497 11084 1503
rect 11213 1204 11219 6316
rect 11261 5884 11267 5896
rect 11293 5504 11299 7876
rect 11245 3544 11251 4736
rect 11293 4724 11299 5496
rect 11309 4884 11315 7916
rect 11517 6764 11523 8096
rect 11645 7724 11651 7796
rect 11661 7704 11667 7796
rect 11565 7104 11571 7696
rect 11773 7524 11779 7756
rect 11469 6504 11475 6556
rect 11645 6504 11651 6596
rect 11661 6524 11667 6756
rect 11517 4404 11523 4476
rect 11277 4104 11283 4356
rect 10925 1004 10931 1116
rect 11133 1044 11139 1196
rect 11245 1124 11251 3536
rect 11277 2944 11283 4096
rect 11309 3884 11315 4276
rect 11437 3304 11443 3676
rect 11453 3204 11459 3916
rect 11613 3304 11619 5516
rect 11709 5324 11715 5356
rect 11677 3924 11683 4896
rect 11645 3324 11651 3396
rect 11309 2924 11315 3096
rect 11613 3024 11619 3196
rect 11277 2844 11283 2916
rect 11309 2504 11315 2896
rect 11309 2004 11315 2096
rect 11293 1164 11299 1296
rect 11172 1117 11180 1123
rect 11197 744 11203 1116
rect 11549 904 11555 2696
rect 11076 517 11084 523
rect 11021 304 11027 356
rect 11469 324 11475 516
rect 11565 224 11571 2336
rect 11581 1704 11587 1916
rect 11581 724 11587 1696
rect 11629 504 11635 3296
rect 11645 2724 11651 2956
rect 11725 2724 11731 3356
rect 11741 3124 11747 7296
rect 11789 7064 11795 7296
rect 11805 6484 11811 8476
rect 12221 8184 12227 8896
rect 12205 7424 12211 8076
rect 12285 7924 12291 8196
rect 11805 5964 11811 6096
rect 11757 5524 11763 5536
rect 11773 3943 11779 5516
rect 11805 5304 11811 5316
rect 11757 3937 11779 3943
rect 11757 3784 11763 3937
rect 11805 3824 11811 5276
rect 11821 4584 11827 6496
rect 11853 6224 11859 7296
rect 11917 6824 11923 7316
rect 12221 7024 12227 7916
rect 12333 7904 12339 8156
rect 11917 6324 11923 6816
rect 11837 5504 11843 5516
rect 11844 5297 11852 5303
rect 11869 5284 11875 5496
rect 11949 4904 11955 5596
rect 12109 4524 12115 4716
rect 11933 4304 11939 4376
rect 11661 524 11667 1216
rect 11645 204 11651 316
rect 11677 264 11683 2296
rect 11741 1284 11747 3116
rect 11773 2824 11779 3396
rect 11805 2904 11811 3136
rect 11773 864 11779 2096
rect 11805 2084 11811 2316
rect 11821 1924 11827 3916
rect 11837 2904 11843 2956
rect 11933 2944 11939 3316
rect 11949 3044 11955 4316
rect 12093 4124 12099 4156
rect 12157 4064 12163 6896
rect 12301 6744 12307 6996
rect 12221 5824 12227 6716
rect 12285 5804 12291 6316
rect 12301 5804 12307 6296
rect 12285 5704 12291 5796
rect 12301 5724 12307 5796
rect 12221 5264 12227 5696
rect 12317 5524 12323 6996
rect 12333 6724 12339 6956
rect 12285 4984 12291 5116
rect 12333 4924 12339 6696
rect 12349 4964 12355 5096
rect 12221 4104 12227 4736
rect 12285 4084 12291 4476
rect 12301 4124 12307 4516
rect 11965 3744 11971 3876
rect 12221 3664 12227 3696
rect 12237 3404 12243 3516
rect 11837 2604 11843 2716
rect 11837 2324 11843 2376
rect 11933 1904 11939 2936
rect 11965 2924 11971 3076
rect 11949 2704 11955 2836
rect 11949 2144 11955 2296
rect 12221 2264 12227 2496
rect 12285 2484 12291 2596
rect 12301 2524 12307 3736
rect 12317 3724 12323 3816
rect 12349 2564 12355 4496
rect 12397 4204 12403 4296
rect 12445 4204 12451 4316
rect 12429 2583 12435 3116
rect 12461 2583 12467 3096
rect 12413 2577 12435 2583
rect 12445 2577 12467 2583
rect 12349 2524 12355 2556
rect 12413 2424 12419 2577
rect 12445 2464 12451 2577
rect 11933 1724 11939 1876
rect 11805 1704 11811 1716
rect 11837 1704 11843 1716
rect 11885 1324 11891 1716
rect 11933 1324 11939 1716
rect 11821 1304 11827 1316
rect 11837 1304 11843 1316
rect 11789 804 11795 1116
rect 11837 904 11843 936
rect 11885 924 11891 1316
rect 11933 924 11939 1316
rect 11805 504 11811 656
rect 12077 564 12083 716
rect 12029 324 12035 476
rect 12205 104 12211 2036
rect 12285 1504 12291 1536
rect 12285 1104 12291 1136
rect 12285 704 12291 736
rect 12477 584 12483 6716
rect 12493 4884 12499 4896
rect 12589 3744 12595 4916
rect 12605 4864 12611 5296
rect 12909 4104 12915 4956
rect 12845 3224 12851 3936
rect 12493 2444 12499 2496
rect 12861 1204 12867 4096
rect 12941 3924 12947 4156
rect 12973 4124 12979 4996
rect 12973 3224 12979 3896
rect 9245 24 9251 96
<< m5contact >>
rect 380 7716 388 7724
rect 92 7496 100 7504
rect 60 4776 68 4784
rect 428 4736 436 4744
rect 524 7916 532 7924
rect 1116 8476 1124 8484
rect 716 8076 724 8084
rect 1036 8076 1044 8084
rect 620 7896 628 7904
rect 540 6396 548 6404
rect 604 5916 612 5924
rect 524 5556 532 5564
rect 684 7716 692 7724
rect 636 7496 644 7504
rect 636 6936 644 6944
rect 620 4756 628 4764
rect 492 4736 500 4744
rect 476 4116 484 4124
rect 588 4276 596 4284
rect 1068 6856 1076 6864
rect 700 4756 708 4764
rect 1420 8896 1428 8904
rect 1884 8896 1892 8904
rect 3388 8896 3396 8904
rect 3772 8896 3780 8904
rect 1820 8716 1828 8724
rect 1276 8396 1284 8404
rect 1292 8036 1300 8044
rect 1276 7996 1284 8004
rect 1164 7956 1172 7964
rect 1132 5536 1140 5544
rect 1276 6716 1284 6724
rect 1180 6696 1188 6704
rect 1180 5116 1188 5124
rect 1212 5096 1220 5104
rect 1260 5096 1268 5104
rect 1164 4836 1172 4844
rect 1244 4516 1252 4524
rect 1164 4336 1172 4344
rect 908 4116 916 4124
rect 124 896 132 904
rect 156 896 164 904
rect 1100 3296 1108 3304
rect 1164 3356 1172 3364
rect 892 1036 900 1044
rect 876 836 884 844
rect 764 716 772 724
rect 844 716 852 724
rect 1164 1496 1172 1504
rect 1196 896 1204 904
rect 1436 6736 1444 6744
rect 1708 7916 1716 7924
rect 1612 6876 1620 6884
rect 1532 6716 1540 6724
rect 1372 4836 1380 4844
rect 1372 4616 1380 4624
rect 1340 3356 1348 3364
rect 1292 2916 1300 2924
rect 1644 1916 1652 1924
rect 1708 7196 1716 7204
rect 1676 5896 1684 5904
rect 1676 5296 1684 5304
rect 1676 5116 1684 5124
rect 2012 7996 2020 8004
rect 1932 7916 1940 7924
rect 1916 6876 1924 6884
rect 1820 6496 1828 6504
rect 1724 5396 1732 5404
rect 1820 5696 1828 5704
rect 1820 5296 1828 5304
rect 1900 5336 1908 5344
rect 1820 5116 1828 5124
rect 1804 4516 1812 4524
rect 1900 4956 1908 4964
rect 1852 3476 1860 3484
rect 1900 3496 1908 3504
rect 1900 2716 1908 2724
rect 3020 8796 3028 8804
rect 2364 8076 2372 8084
rect 2204 6856 2212 6864
rect 1820 2316 1828 2324
rect 1820 2096 1828 2104
rect 1436 1516 1444 1524
rect 1276 556 1284 564
rect 780 316 788 324
rect 844 316 852 324
rect 1580 1036 1588 1044
rect 1564 836 1572 844
rect 1532 516 1540 524
rect 1404 316 1412 324
rect 1564 556 1572 564
rect 1948 5476 1956 5484
rect 1996 3876 2004 3884
rect 1980 3356 1988 3364
rect 2060 4696 2068 4704
rect 2076 3896 2084 3904
rect 2044 3356 2052 3364
rect 1948 2916 1956 2924
rect 2396 7536 2404 7544
rect 2412 6696 2420 6704
rect 2348 5296 2356 5304
rect 2332 5116 2340 5124
rect 2316 3896 2324 3904
rect 1948 1936 1956 1944
rect 2220 1536 2228 1544
rect 2172 796 2180 804
rect 2204 896 2212 904
rect 2076 516 2084 524
rect 2220 516 2228 524
rect 1756 96 1764 104
rect 1820 96 1828 104
rect 2348 3956 2356 3964
rect 2412 6076 2420 6084
rect 2380 4616 2388 4624
rect 2364 1516 2372 1524
rect 2332 1496 2340 1504
rect 2652 7956 2660 7964
rect 2732 7916 2740 7924
rect 2572 7496 2580 7504
rect 2812 7096 2820 7104
rect 2748 6876 2756 6884
rect 3052 7536 3060 7544
rect 3228 7916 3236 7924
rect 3228 7876 3236 7884
rect 3020 6936 3028 6944
rect 2716 6696 2724 6704
rect 2572 6116 2580 6124
rect 2476 4616 2484 4624
rect 2540 3336 2548 3344
rect 2476 2496 2484 2504
rect 2844 6536 2852 6544
rect 3116 6296 3124 6304
rect 3116 6036 3124 6044
rect 2572 5116 2580 5124
rect 2652 5076 2660 5084
rect 2700 4516 2708 4524
rect 2812 4436 2820 4444
rect 2780 3876 2788 3884
rect 2572 3596 2580 3604
rect 2812 3336 2820 3344
rect 2668 3316 2676 3324
rect 2572 3296 2580 3304
rect 2780 3276 2788 3284
rect 2460 2116 2468 2124
rect 2540 2116 2548 2124
rect 2460 1536 2468 1544
rect 2684 3096 2692 3104
rect 2764 1936 2772 1944
rect 2604 1856 2612 1864
rect 2748 1516 2756 1524
rect 2572 1036 2580 1044
rect 2748 896 2756 904
rect 2732 796 2740 804
rect 3052 5336 3060 5344
rect 3164 6296 3172 6304
rect 3004 4096 3012 4104
rect 2860 3336 2868 3344
rect 2844 3316 2852 3324
rect 2844 2536 2852 2544
rect 2844 2496 2852 2504
rect 2828 796 2836 804
rect 2460 316 2468 324
rect 2220 96 2228 104
rect 3052 2736 3060 2744
rect 2876 2096 2884 2104
rect 2876 1516 2884 1524
rect 2860 896 2868 904
rect 3260 5496 3268 5504
rect 3228 4716 3236 4724
rect 3196 4336 3204 4344
rect 3228 4336 3236 4344
rect 3212 3976 3220 3984
rect 3228 3736 3236 3744
rect 3116 1716 3124 1724
rect 3196 3596 3204 3604
rect 3148 1116 3156 1124
rect 3340 7496 3348 7504
rect 3484 8116 3492 8124
rect 3388 6736 3396 6744
rect 3388 6696 3396 6704
rect 3836 7896 3844 7904
rect 3884 7896 3892 7904
rect 3772 7736 3780 7744
rect 3852 7736 3860 7744
rect 3868 7696 3876 7704
rect 3532 7516 3540 7524
rect 3500 7316 3508 7324
rect 3500 5176 3508 5184
rect 3484 5116 3492 5124
rect 3388 5076 3396 5084
rect 3276 2676 3284 2684
rect 3404 4716 3412 4724
rect 3484 4496 3492 4504
rect 3324 4316 3332 4324
rect 3324 3996 3332 4004
rect 3340 3976 3348 3984
rect 3436 4316 3444 4324
rect 3644 7496 3652 7504
rect 3628 5696 3636 5704
rect 3628 5476 3636 5484
rect 3788 7096 3796 7104
rect 3772 5476 3780 5484
rect 3324 3476 3332 3484
rect 3308 3296 3316 3304
rect 3308 2916 3316 2924
rect 3228 1416 3236 1424
rect 3388 3736 3396 3744
rect 3356 2816 3364 2824
rect 3420 2796 3428 2804
rect 3468 2696 3476 2704
rect 3340 2176 3348 2184
rect 3500 3316 3508 3324
rect 3484 2116 3492 2124
rect 3324 1916 3332 1924
rect 3468 1876 3476 1884
rect 3420 1596 3428 1604
rect 3772 4896 3780 4904
rect 3852 6716 3860 6724
rect 3836 6056 3844 6064
rect 3884 6316 3892 6324
rect 3916 6296 3924 6304
rect 3868 5496 3876 5504
rect 3868 5476 3876 5484
rect 3868 4776 3876 4784
rect 3772 4016 3780 4024
rect 3868 3116 3876 3124
rect 3884 3096 3892 3104
rect 3900 3096 3908 3104
rect 3836 2596 3844 2604
rect 3532 1776 3540 1784
rect 3388 1116 3396 1124
rect 3628 1716 3636 1724
rect 4060 7916 4068 7924
rect 4012 6096 4020 6104
rect 3948 4736 3956 4744
rect 3964 3916 3972 3924
rect 3964 3276 3972 3284
rect 3996 4436 4004 4444
rect 4044 6296 4052 6304
rect 4044 4476 4052 4484
rect 5484 8896 5492 8904
rect 4140 8396 4148 8404
rect 4588 8396 4596 8404
rect 4156 6916 4164 6924
rect 4092 6096 4100 6104
rect 4604 8296 4612 8304
rect 4956 8736 4964 8744
rect 4604 7736 4612 7744
rect 4652 7736 4660 7744
rect 4412 7096 4420 7104
rect 4428 7096 4436 7104
rect 4508 6716 4516 6724
rect 4668 6716 4676 6724
rect 4508 6516 4516 6524
rect 4620 6396 4628 6404
rect 4508 5336 4516 5344
rect 4588 5496 4596 5504
rect 4540 5176 4548 5184
rect 4668 5316 4676 5324
rect 4140 4796 4148 4804
rect 4508 4796 4516 4804
rect 3932 2096 3940 2104
rect 3900 1696 3908 1704
rect 3836 1636 3844 1644
rect 3884 1636 3892 1644
rect 3996 1936 4004 1944
rect 3964 1916 3972 1924
rect 3980 1916 3988 1924
rect 3996 936 4004 944
rect 3852 876 3860 884
rect 3628 316 3636 324
rect 4044 1856 4052 1864
rect 4428 4756 4436 4764
rect 4156 4256 4164 4264
rect 4780 8116 4788 8124
rect 4748 8096 4756 8104
rect 4780 7536 4788 7544
rect 4956 7516 4964 7524
rect 4780 6716 4788 6724
rect 4780 6316 4788 6324
rect 4780 5276 4788 5284
rect 4684 4716 4692 4724
rect 4428 4316 4436 4324
rect 4172 3336 4180 3344
rect 4524 2916 4532 2924
rect 4428 2696 4436 2704
rect 4364 2476 4372 2484
rect 4460 2476 4468 2484
rect 4412 2096 4420 2104
rect 4540 1756 4548 1764
rect 4076 1096 4084 1104
rect 4812 5156 4820 5164
rect 4796 4476 4804 4484
rect 4684 3996 4692 4004
rect 4412 896 4420 904
rect 4780 3956 4788 3964
rect 4796 3476 4804 3484
rect 4796 3116 4804 3124
rect 4924 4716 4932 4724
rect 5260 8316 5268 8324
rect 5276 7916 5284 7924
rect 5068 5916 5076 5924
rect 5132 7696 5140 7704
rect 5276 7196 5284 7204
rect 5164 6816 5172 6824
rect 5180 6696 5188 6704
rect 5180 5596 5188 5604
rect 5036 4756 5044 4764
rect 5020 4696 5028 4704
rect 5132 4476 5140 4484
rect 4828 3256 4836 3264
rect 4700 2696 4708 2704
rect 4764 2676 4772 2684
rect 4764 2596 4772 2604
rect 4652 1516 4660 1524
rect 4812 2716 4820 2724
rect 4812 2696 4820 2704
rect 4796 2096 4804 2104
rect 4988 2456 4996 2464
rect 5020 2456 5028 2464
rect 4940 2296 4948 2304
rect 4924 2176 4932 2184
rect 5180 4356 5188 4364
rect 5148 4116 5156 4124
rect 5164 4116 5172 4124
rect 5148 4076 5156 4084
rect 5196 4136 5204 4144
rect 5132 2536 5140 2544
rect 5388 7916 5396 7924
rect 5452 7876 5460 7884
rect 5388 7316 5396 7324
rect 5340 6916 5348 6924
rect 5356 6696 5364 6704
rect 5340 6036 5348 6044
rect 5340 5896 5348 5904
rect 5292 5556 5300 5564
rect 5324 5116 5332 5124
rect 5404 6716 5412 6724
rect 5452 5916 5460 5924
rect 5420 5336 5428 5344
rect 5436 5296 5444 5304
rect 5420 5196 5428 5204
rect 5404 5176 5412 5184
rect 5420 5116 5428 5124
rect 5388 2476 5396 2484
rect 5404 2476 5412 2484
rect 5148 2336 5156 2344
rect 5148 2116 5156 2124
rect 5340 2096 5348 2104
rect 5228 1876 5236 1884
rect 5276 1876 5284 1884
rect 5820 7696 5828 7704
rect 5996 8476 6004 8484
rect 5996 8316 6004 8324
rect 5484 4896 5492 4904
rect 5692 5676 5700 5684
rect 5644 3916 5652 3924
rect 6012 6456 6020 6464
rect 5996 5676 6004 5684
rect 5852 5196 5860 5204
rect 5948 5176 5956 5184
rect 5820 4356 5828 4364
rect 5804 4296 5812 4304
rect 5804 4096 5812 4104
rect 5804 3696 5812 3704
rect 5788 3656 5796 3664
rect 5436 2856 5444 2864
rect 5644 2596 5652 2604
rect 5644 1916 5652 1924
rect 5132 1116 5140 1124
rect 5180 1096 5188 1104
rect 5612 1096 5620 1104
rect 4684 876 4692 884
rect 5068 536 5076 544
rect 5164 456 5172 464
rect 5132 336 5140 344
rect 5788 2036 5796 2044
rect 5772 1956 5780 1964
rect 5916 4116 5924 4124
rect 5884 4076 5892 4084
rect 5836 3556 5844 3564
rect 5820 1316 5828 1324
rect 5996 4716 6004 4724
rect 6044 7936 6052 7944
rect 6572 8316 6580 8324
rect 6636 8316 6644 8324
rect 6108 7556 6116 7564
rect 6092 6536 6100 6544
rect 6044 6456 6052 6464
rect 6268 5516 6276 5524
rect 6364 7716 6372 7724
rect 6396 7696 6404 7704
rect 6572 6836 6580 6844
rect 6604 7916 6612 7924
rect 6636 6516 6644 6524
rect 6316 5516 6324 5524
rect 6092 3956 6100 3964
rect 6076 3156 6084 3164
rect 5884 2316 5892 2324
rect 6060 1736 6068 1744
rect 5964 1676 5972 1684
rect 6044 1636 6052 1644
rect 6028 736 6036 744
rect 5660 536 5668 544
rect 6236 4316 6244 4324
rect 6268 3696 6276 3704
rect 6236 3156 6244 3164
rect 6332 3436 6340 3444
rect 6380 5556 6388 5564
rect 6412 5276 6420 5284
rect 6460 5116 6468 5124
rect 6380 4096 6388 4104
rect 6428 3096 6436 3104
rect 6092 916 6100 924
rect 6076 496 6084 504
rect 6380 1996 6388 2004
rect 6396 1796 6404 1804
rect 6348 1436 6356 1444
rect 6460 3976 6468 3984
rect 6604 5096 6612 5104
rect 6700 6536 6708 6544
rect 6700 6516 6708 6524
rect 6684 6136 6692 6144
rect 6668 5676 6676 5684
rect 6700 5096 6708 5104
rect 6748 6096 6756 6104
rect 6780 5296 6788 5304
rect 6748 5116 6756 5124
rect 6748 5076 6756 5084
rect 6732 3956 6740 3964
rect 6780 4376 6788 4384
rect 6764 4356 6772 4364
rect 7036 5676 7044 5684
rect 7148 7576 7156 7584
rect 7196 7576 7204 7584
rect 7132 6536 7140 6544
rect 6748 3556 6756 3564
rect 6636 3116 6644 3124
rect 6588 2856 6596 2864
rect 6492 2796 6500 2804
rect 6636 2296 6644 2304
rect 6956 2796 6964 2804
rect 6444 1536 6452 1544
rect 6540 1436 6548 1444
rect 6476 1096 6484 1104
rect 6636 1956 6644 1964
rect 6732 1776 6740 1784
rect 6636 1736 6644 1744
rect 7084 4756 7092 4764
rect 7084 4276 7092 4284
rect 7100 4116 7108 4124
rect 7100 4076 7108 4084
rect 7356 6836 7364 6844
rect 7388 6596 7396 6604
rect 7660 8296 7668 8304
rect 7660 6816 7668 6824
rect 7404 6396 7412 6404
rect 7212 5316 7220 5324
rect 7404 4916 7412 4924
rect 7212 4756 7220 4764
rect 7292 4356 7300 4364
rect 7292 4096 7300 4104
rect 7308 4076 7316 4084
rect 7292 4056 7300 4064
rect 7404 4776 7412 4784
rect 7436 4776 7444 4784
rect 7388 3716 7396 3724
rect 7388 3696 7396 3704
rect 7372 3676 7380 3684
rect 7116 3436 7124 3444
rect 7100 3316 7108 3324
rect 7084 2936 7092 2944
rect 7148 3136 7156 3144
rect 7212 2916 7220 2924
rect 5980 436 5988 444
rect 6044 436 6052 444
rect 6092 436 6100 444
rect 5660 356 5668 364
rect 5964 316 5972 324
rect 5996 356 6004 364
rect 6012 316 6020 324
rect 5820 296 5828 304
rect 5964 276 5972 284
rect 5948 116 5956 124
rect 6620 336 6628 344
rect 6796 936 6804 944
rect 6812 936 6820 944
rect 7196 1996 7204 2004
rect 7020 896 7028 904
rect 6684 436 6692 444
rect 6908 396 6916 404
rect 6748 296 6756 304
rect 6684 136 6692 144
rect 6044 96 6052 104
rect 7228 1936 7236 1944
rect 7436 3316 7444 3324
rect 7292 1296 7300 1304
rect 7532 4856 7540 4864
rect 7644 6136 7652 6144
rect 7612 4036 7620 4044
rect 7564 1076 7572 1084
rect 8428 8796 8436 8804
rect 8396 8496 8404 8504
rect 8268 8316 8276 8324
rect 8348 8316 8356 8324
rect 7900 7936 7908 7944
rect 7756 7896 7764 7904
rect 7948 7896 7956 7904
rect 7916 7516 7924 7524
rect 7964 7516 7972 7524
rect 7676 4736 7684 4744
rect 7836 5496 7844 5504
rect 7788 4796 7796 4804
rect 7852 4316 7860 4324
rect 7884 4276 7892 4284
rect 7708 3436 7716 3444
rect 7708 2956 7716 2964
rect 7772 2936 7780 2944
rect 7772 2916 7780 2924
rect 7788 2356 7796 2364
rect 7852 2356 7860 2364
rect 7836 2116 7844 2124
rect 7772 1696 7780 1704
rect 8012 7936 8020 7944
rect 8220 8096 8228 8104
rect 8060 7516 8068 7524
rect 8012 7496 8020 7504
rect 8012 6516 8020 6524
rect 7948 5736 7956 5744
rect 8076 5736 8084 5744
rect 8028 5696 8036 5704
rect 8012 5236 8020 5244
rect 7948 5116 7956 5124
rect 7948 4316 7956 4324
rect 7948 4116 7956 4124
rect 7932 3116 7940 3124
rect 8220 6536 8228 6544
rect 8300 6316 8308 6324
rect 8252 6056 8260 6064
rect 8332 5896 8340 5904
rect 8348 5496 8356 5504
rect 8396 4936 8404 4944
rect 8588 8096 8596 8104
rect 8508 6916 8516 6924
rect 8524 6716 8532 6724
rect 8476 6696 8484 6704
rect 8444 5156 8452 5164
rect 8412 4896 8420 4904
rect 8028 4796 8036 4804
rect 8588 6896 8596 6904
rect 8588 6096 8596 6104
rect 9884 8896 9892 8904
rect 9612 8736 9620 8744
rect 9340 8716 9348 8724
rect 9788 8716 9796 8724
rect 9196 8496 9204 8504
rect 9244 8496 9252 8504
rect 9244 8036 9252 8044
rect 8700 6096 8708 6104
rect 8652 5936 8660 5944
rect 8588 5696 8596 5704
rect 8636 4896 8644 4904
rect 8668 5076 8676 5084
rect 8588 4736 8596 4744
rect 8556 4536 8564 4544
rect 8700 4956 8708 4964
rect 8044 4116 8052 4124
rect 8044 3976 8052 3984
rect 8588 4096 8596 4104
rect 8524 3856 8532 3864
rect 8620 3736 8628 3744
rect 8572 3716 8580 3724
rect 8636 3556 8644 3564
rect 8588 3456 8596 3464
rect 7996 2496 8004 2504
rect 8012 2296 8020 2304
rect 8044 2936 8052 2944
rect 8588 2936 8596 2944
rect 8572 2916 8580 2924
rect 8524 2896 8532 2904
rect 8444 2716 8452 2724
rect 8220 2676 8228 2684
rect 8364 2676 8372 2684
rect 8316 2596 8324 2604
rect 8428 2476 8436 2484
rect 8300 2036 8308 2044
rect 8220 1496 8228 1504
rect 8060 1476 8068 1484
rect 8380 936 8388 944
rect 8620 2536 8628 2544
rect 8588 2316 8596 2324
rect 8748 6916 8756 6924
rect 8748 4536 8756 4544
rect 8860 4136 8868 4144
rect 8732 4016 8740 4024
rect 8700 3756 8708 3764
rect 8732 3756 8740 3764
rect 8684 3736 8692 3744
rect 8700 3736 8708 3744
rect 8668 1916 8676 1924
rect 8476 1096 8484 1104
rect 9244 7696 9252 7704
rect 9036 7516 9044 7524
rect 8988 7496 8996 7504
rect 8972 5896 8980 5904
rect 9356 7896 9364 7904
rect 9340 7196 9348 7204
rect 9356 7016 9364 7024
rect 9388 6996 9396 7004
rect 9324 5916 9332 5924
rect 9244 5716 9252 5724
rect 9244 5516 9252 5524
rect 9052 4376 9060 4384
rect 8972 4136 8980 4144
rect 9308 5236 9316 5244
rect 9244 4696 9252 4704
rect 9052 4016 9060 4024
rect 8700 2116 8708 2124
rect 8588 1076 8596 1084
rect 9020 3376 9028 3384
rect 9068 3536 9076 3544
rect 9052 2796 9060 2804
rect 9036 1936 9044 1944
rect 8524 896 8532 904
rect 7564 496 7572 504
rect 7660 496 7668 504
rect 7404 396 7412 404
rect 7948 276 7956 284
rect 9052 1496 9060 1504
rect 9052 1476 9060 1484
rect 9052 1116 9060 1124
rect 9036 716 9044 724
rect 9244 3136 9252 3144
rect 9372 4376 9380 4384
rect 9324 3116 9332 3124
rect 9340 3096 9348 3104
rect 9196 2896 9204 2904
rect 9196 2516 9204 2524
rect 9116 2496 9124 2504
rect 9244 2316 9252 2324
rect 9516 3196 9524 3204
rect 9372 2916 9380 2924
rect 9244 2096 9252 2104
rect 9196 1936 9204 1944
rect 9132 1896 9140 1904
rect 9324 1536 9332 1544
rect 9244 1316 9252 1324
rect 9212 1276 9220 1284
rect 9068 516 9076 524
rect 7948 116 7956 124
rect 8924 136 8932 144
rect 9196 96 9204 104
rect 9724 7496 9732 7504
rect 9836 6876 9844 6884
rect 9852 6796 9860 6804
rect 9820 6696 9828 6704
rect 9884 6316 9892 6324
rect 9788 6076 9796 6084
rect 9996 7716 10004 7724
rect 10012 6676 10020 6684
rect 9852 5936 9860 5944
rect 9884 5916 9892 5924
rect 9724 5876 9732 5884
rect 9884 4916 9892 4924
rect 9724 4496 9732 4504
rect 9724 3716 9732 3724
rect 9884 3716 9892 3724
rect 9836 3676 9844 3684
rect 9740 2596 9748 2604
rect 9676 676 9684 684
rect 9868 3696 9876 3704
rect 9820 3036 9828 3044
rect 9884 2876 9892 2884
rect 9884 2436 9892 2444
rect 10124 7016 10132 7024
rect 10140 6896 10148 6904
rect 9980 4876 9988 4884
rect 10028 4416 10036 4424
rect 9916 4076 9924 4084
rect 9916 3296 9924 3304
rect 9980 2156 9988 2164
rect 10044 2616 10052 2624
rect 10044 2536 10052 2544
rect 10396 8256 10404 8264
rect 10540 8096 10548 8104
rect 10428 7496 10436 7504
rect 10316 6636 10324 6644
rect 10332 6536 10340 6544
rect 10348 6516 10356 6524
rect 10332 6496 10340 6504
rect 10348 6136 10356 6144
rect 10348 5596 10356 5604
rect 10332 5536 10340 5544
rect 10380 6136 10388 6144
rect 10268 4896 10276 4904
rect 10268 4736 10276 4744
rect 10348 4536 10356 4544
rect 10268 4316 10276 4324
rect 10348 4296 10356 4304
rect 10348 4176 10356 4184
rect 10268 3916 10276 3924
rect 10396 5556 10404 5564
rect 10396 3496 10404 3504
rect 10140 2116 10148 2124
rect 10476 4496 10484 4504
rect 10540 7296 10548 7304
rect 10540 6736 10548 6744
rect 10540 6096 10548 6104
rect 10524 5916 10532 5924
rect 10540 5896 10548 5904
rect 10540 5516 10548 5524
rect 10524 5496 10532 5504
rect 10492 4316 10500 4324
rect 10268 1696 10276 1704
rect 9996 1296 10004 1304
rect 10572 5096 10580 5104
rect 10540 5076 10548 5084
rect 10540 4936 10548 4944
rect 10636 6696 10644 6704
rect 10684 7716 10692 7724
rect 11084 7896 11092 7904
rect 10988 7556 10996 7564
rect 10700 6816 10708 6824
rect 10684 6796 10692 6804
rect 10588 3636 10596 3644
rect 10684 5296 10692 5304
rect 10684 4016 10692 4024
rect 10540 2716 10548 2724
rect 10652 2536 10660 2544
rect 10524 2436 10532 2444
rect 10636 1496 10644 1504
rect 10540 716 10548 724
rect 10332 676 10340 684
rect 10684 2496 10692 2504
rect 11196 7536 11204 7544
rect 11196 6876 11204 6884
rect 11148 5916 11156 5924
rect 10972 5336 10980 5344
rect 11180 4896 11188 4904
rect 10924 2496 10932 2504
rect 11004 1936 11012 1944
rect 11084 4136 11092 4144
rect 11084 4036 11092 4044
rect 11084 2916 11092 2924
rect 11180 3536 11188 3544
rect 11084 2536 11092 2544
rect 11196 2496 11204 2504
rect 11196 1916 11204 1924
rect 11132 1536 11140 1544
rect 11084 1496 11092 1504
rect 11260 5896 11268 5904
rect 11740 7696 11748 7704
rect 11308 4876 11316 4884
rect 11244 3536 11252 3544
rect 11132 1196 11140 1204
rect 11212 1196 11220 1204
rect 11436 3676 11444 3684
rect 11452 3196 11460 3204
rect 11612 3196 11620 3204
rect 11276 2916 11284 2924
rect 11308 2916 11316 2924
rect 11308 2496 11316 2504
rect 11164 1116 11172 1124
rect 11244 1116 11252 1124
rect 11084 516 11092 524
rect 11756 5516 11764 5524
rect 11804 5316 11812 5324
rect 11804 5276 11812 5284
rect 11948 5596 11956 5604
rect 11836 5516 11844 5524
rect 11836 5296 11844 5304
rect 11868 5276 11876 5284
rect 11836 2956 11844 2964
rect 11948 3036 11956 3044
rect 11932 1876 11940 1884
rect 11804 1716 11812 1724
rect 11884 1716 11892 1724
rect 11836 1696 11844 1704
rect 11820 1316 11828 1324
rect 11884 1316 11892 1324
rect 11836 1296 11844 1304
rect 12492 4876 12500 4884
rect 9244 96 9252 104
<< metal5 >>
rect 1428 8897 1884 8903
rect 3396 8897 3772 8903
rect 3780 8897 5484 8903
rect 9892 8897 10011 8903
rect 3028 8797 8428 8803
rect 4964 8737 9612 8743
rect 1701 8717 1820 8723
rect 9348 8717 9788 8723
rect 8404 8497 9196 8503
rect 9252 8497 9371 8503
rect 1124 8477 5996 8483
rect 1284 8397 4140 8403
rect 4148 8397 4588 8403
rect 5268 8317 5996 8323
rect 6580 8317 6636 8323
rect 8276 8317 8348 8323
rect 4612 8297 7660 8303
rect 10373 8257 10396 8263
rect 3492 8117 4780 8123
rect 4756 8097 4827 8103
rect 8228 8097 8588 8103
rect 9349 8097 10540 8103
rect 724 8077 1036 8083
rect 1044 8077 2364 8083
rect 1300 8037 9244 8043
rect 1284 7997 2012 8003
rect 1172 7957 2652 7963
rect 4141 7937 6044 7943
rect 532 7917 1708 7923
rect 1940 7917 2732 7923
rect 4141 7923 4147 7937
rect 6052 7937 7900 7943
rect 7908 7937 8012 7943
rect 4068 7917 4147 7923
rect 5284 7917 5388 7923
rect 5396 7917 5403 7923
rect 5413 7917 6604 7923
rect 628 7897 3836 7903
rect 3844 7897 3884 7903
rect 3892 7897 7756 7903
rect 7764 7897 7948 7903
rect 9364 7897 11084 7903
rect 3236 7877 5452 7883
rect 3780 7737 3852 7743
rect 4612 7737 4652 7743
rect 388 7717 684 7723
rect 6372 7717 9996 7723
rect 3876 7697 5132 7703
rect 5828 7697 6396 7703
rect 9252 7697 9339 7703
rect 10661 7697 11740 7703
rect 7156 7577 7196 7583
rect 6116 7557 10988 7563
rect 2404 7537 3052 7543
rect 4788 7537 11196 7543
rect 3540 7517 4956 7523
rect 7924 7517 7964 7523
rect 8068 7517 9036 7523
rect 100 7497 636 7503
rect 2580 7497 2843 7503
rect 3348 7497 3644 7503
rect 8020 7497 8988 7503
rect 9732 7497 10428 7503
rect 3508 7317 5388 7323
rect 10548 7297 10683 7303
rect 1716 7197 5276 7203
rect 5284 7197 9340 7203
rect 2820 7097 3788 7103
rect 3796 7097 4412 7103
rect 4420 7097 4428 7103
rect 9364 7017 10124 7023
rect 9381 6997 9388 7003
rect 644 6937 3020 6943
rect 4164 6917 5340 6923
rect 8516 6917 8748 6923
rect 8596 6897 10140 6903
rect 1620 6877 1916 6883
rect 2756 6877 2875 6883
rect 9844 6877 11196 6883
rect 1076 6857 2204 6863
rect 6580 6837 7356 6843
rect 5172 6817 7660 6823
rect 7668 6817 10700 6823
rect 9860 6797 10683 6803
rect 1444 6737 3388 6743
rect 10548 6737 10683 6743
rect 1284 6717 1532 6723
rect 1540 6717 3852 6723
rect 3860 6717 4508 6723
rect 4676 6717 4780 6723
rect 5412 6717 8524 6723
rect 1188 6697 2412 6703
rect 2724 6697 2779 6703
rect 3396 6697 5180 6703
rect 5364 6697 8476 6703
rect 9828 6697 10636 6703
rect 8741 6637 10316 6643
rect 7396 6597 7419 6603
rect 1925 6537 2844 6543
rect 6100 6537 6700 6543
rect 7140 6537 8220 6543
rect 4516 6517 6636 6523
rect 6708 6517 6747 6523
rect 8020 6517 10348 6523
rect 10356 6517 10395 6523
rect 1828 6497 1915 6503
rect 10221 6497 10332 6503
rect 8037 6477 10203 6483
rect 10221 6483 10227 6497
rect 10213 6477 10227 6483
rect 6020 6457 6044 6463
rect 548 6397 4620 6403
rect 4628 6397 7404 6403
rect 3892 6317 4780 6323
rect 8308 6317 9884 6323
rect 3124 6297 3164 6303
rect 3924 6297 4044 6303
rect 6692 6137 7644 6143
rect 10356 6137 10380 6143
rect 2580 6117 2779 6123
rect 4020 6097 4092 6103
rect 6756 6097 8588 6103
rect 8596 6097 8700 6103
rect 9349 6097 10540 6103
rect 2420 6077 9788 6083
rect 3844 6057 8252 6063
rect 3124 6037 5340 6043
rect 8660 5937 9852 5943
rect 612 5917 635 5923
rect 5076 5917 5452 5923
rect 5460 5917 9324 5923
rect 9332 5917 9884 5923
rect 10532 5917 11148 5923
rect 1684 5897 5340 5903
rect 8340 5897 8859 5903
rect 8869 5897 8972 5903
rect 8980 5897 10540 5903
rect 11268 5897 11291 5903
rect 8709 5877 9724 5883
rect 7956 5737 8076 5743
rect 9252 5717 9371 5723
rect 8029 5704 8035 5715
rect 1828 5697 3628 5703
rect 8596 5697 8731 5703
rect 5700 5677 5996 5683
rect 6676 5677 6779 5683
rect 6789 5677 7036 5683
rect 5029 5597 5180 5603
rect 5188 5597 8699 5603
rect 10356 5597 11291 5603
rect 11301 5597 11948 5603
rect 532 5557 5292 5563
rect 6388 5557 10396 5563
rect 645 5537 1132 5543
rect 6276 5517 6316 5523
rect 8069 5517 9244 5523
rect 9252 5517 9371 5523
rect 9381 5517 10540 5523
rect 11764 5517 11836 5523
rect 3268 5497 3868 5503
rect 3876 5497 4588 5503
rect 6757 5497 7836 5503
rect 8356 5497 10524 5503
rect 1949 5484 1955 5495
rect 3636 5477 3772 5483
rect 3780 5477 3868 5483
rect 1701 5397 1724 5403
rect 1908 5337 3052 5343
rect 4516 5337 5420 5343
rect 10405 5337 10972 5343
rect 4676 5317 4731 5323
rect 4741 5317 7212 5323
rect 7220 5317 7387 5323
rect 10213 5317 10619 5323
rect 10629 5317 11804 5323
rect 1684 5297 1820 5303
rect 1828 5297 2348 5303
rect 5444 5297 6780 5303
rect 10692 5297 11836 5303
rect 4788 5277 6412 5283
rect 11812 5277 11868 5283
rect 8020 5237 9308 5243
rect 5428 5197 5852 5203
rect 3508 5177 4540 5183
rect 4548 5177 5404 5183
rect 5412 5177 5948 5183
rect 4820 5157 8444 5163
rect 1188 5117 1676 5123
rect 1828 5117 2332 5123
rect 2580 5117 3484 5123
rect 5332 5117 5420 5123
rect 6468 5117 6748 5123
rect 7956 5117 8059 5123
rect 1220 5097 1260 5103
rect 1268 5097 4731 5103
rect 6437 5097 6604 5103
rect 6612 5097 6700 5103
rect 10580 5097 10651 5103
rect 6749 5084 6755 5095
rect 2660 5077 3388 5083
rect 8676 5077 10540 5083
rect 1908 4957 1915 4963
rect 8404 4937 10540 4943
rect 7412 4917 9884 4923
rect 3780 4897 5484 4903
rect 8420 4897 8636 4903
rect 10276 4897 11180 4903
rect 9988 4877 11308 4883
rect 11316 4877 12492 4883
rect 7540 4857 9339 4863
rect 1172 4837 1372 4843
rect 4148 4797 4508 4803
rect 7796 4797 8028 4803
rect 68 4777 1275 4783
rect 3876 4777 7404 4783
rect 7412 4777 7436 4783
rect 628 4757 700 4763
rect 4436 4757 5036 4763
rect 7092 4757 7212 4763
rect 436 4737 492 4743
rect 3956 4737 7676 4743
rect 7684 4737 8588 4743
rect 8596 4737 10268 4743
rect 3397 4717 3404 4723
rect 3412 4717 4684 4723
rect 4932 4717 5996 4723
rect 2068 4697 3483 4703
rect 5028 4697 9244 4703
rect 1380 4617 1755 4623
rect 2388 4617 2476 4623
rect 8564 4537 8748 4543
rect 10356 4537 10363 4543
rect 1252 4517 1275 4523
rect 1765 4517 1804 4523
rect 1812 4517 2700 4523
rect 3485 4504 3491 4515
rect 9732 4497 10476 4503
rect 4052 4477 4155 4483
rect 4804 4477 5132 4483
rect 5140 4477 5403 4483
rect 5413 4477 9339 4483
rect 2820 4437 3996 4443
rect 3333 4417 8859 4423
rect 8869 4417 10028 4423
rect 6788 4377 9052 4383
rect 9060 4377 9372 4383
rect 5828 4357 6764 4363
rect 6772 4357 7292 4363
rect 5181 4345 5187 4356
rect 1172 4337 3196 4343
rect 3332 4317 3436 4323
rect 4436 4317 6236 4323
rect 7860 4317 7948 4323
rect 10276 4317 10492 4323
rect 5812 4297 5819 4303
rect 5829 4297 6779 4303
rect 10356 4297 10363 4303
rect 596 4277 7084 4283
rect 7892 4277 8051 4283
rect 5189 4137 5196 4143
rect 8045 4124 8051 4277
rect 10356 4177 10363 4183
rect 8868 4137 8972 4143
rect 8980 4137 11084 4143
rect 484 4117 908 4123
rect 5156 4117 5164 4123
rect 5172 4117 5916 4123
rect 7108 4117 7948 4123
rect 3012 4097 5804 4103
rect 6388 4097 7292 4103
rect 8421 4097 8588 4103
rect 5029 4077 5148 4083
rect 5156 4077 5884 4083
rect 7108 4077 7308 4083
rect 9924 4077 10011 4083
rect 3461 4057 7292 4063
rect 7300 4057 7419 4063
rect 7620 4037 11084 4043
rect 3780 4017 5019 4023
rect 5029 4017 8732 4023
rect 8740 4017 9052 4023
rect 9060 4017 10651 4023
rect 10661 4017 10684 4023
rect 3332 3997 4684 4003
rect 4692 3997 8059 4003
rect 3220 3977 3340 3983
rect 6468 3977 7387 3983
rect 8052 3977 8059 3983
rect 2356 3957 3867 3963
rect 4788 3957 6092 3963
rect 6100 3957 6732 3963
rect 3972 3917 5644 3923
rect 10276 3917 10395 3923
rect 2084 3897 2316 3903
rect 2004 3877 2780 3883
rect 8532 3857 8635 3863
rect 8708 3757 8732 3763
rect 3236 3737 3388 3743
rect 8628 3737 8684 3743
rect 7396 3717 7419 3723
rect 8580 3717 8635 3723
rect 9732 3717 9884 3723
rect 5812 3697 6268 3703
rect 9876 3697 9947 3703
rect 7380 3677 7387 3683
rect 9844 3677 11436 3683
rect 5796 3657 8027 3663
rect 10596 3637 10619 3643
rect 2580 3597 3196 3603
rect 5844 3557 6748 3563
rect 6756 3557 8636 3563
rect 11188 3537 11244 3543
rect 9069 3523 9075 3536
rect 9069 3517 9083 3523
rect 1908 3497 1915 3503
rect 4797 3484 4803 3495
rect 1860 3477 3324 3483
rect 3237 3457 8588 3463
rect 6340 3437 7116 3443
rect 7124 3437 7708 3443
rect 7716 3437 8059 3443
rect 8069 3437 8635 3443
rect 9028 3377 9051 3383
rect 1172 3357 1340 3363
rect 1988 3357 2044 3363
rect 2548 3337 2812 3343
rect 2853 3337 2860 3343
rect 2868 3337 4172 3343
rect 2676 3317 2844 3323
rect 2852 3317 3500 3323
rect 7108 3317 7436 3323
rect 1108 3297 2572 3303
rect 2580 3297 3308 3303
rect 9924 3297 9947 3303
rect 2788 3277 3964 3283
rect 9524 3197 11452 3203
rect 11460 3197 11612 3203
rect 6084 3157 6236 3163
rect 7156 3137 9244 3143
rect 3876 3117 4796 3123
rect 4804 3117 6636 3123
rect 6644 3117 7387 3123
rect 7397 3117 7932 3123
rect 9317 3117 9324 3123
rect 2692 3097 3884 3103
rect 3892 3097 3900 3103
rect 6436 3097 9340 3103
rect 9828 3037 11948 3043
rect 7716 2957 11836 2963
rect 7092 2937 7772 2943
rect 8052 2937 8588 2943
rect 1300 2917 1948 2923
rect 1956 2917 3308 2923
rect 3316 2917 3323 2923
rect 4532 2917 4795 2923
rect 7220 2917 7387 2923
rect 7780 2917 8572 2923
rect 9380 2917 11084 2923
rect 11284 2917 11308 2923
rect 8532 2897 8635 2903
rect 8645 2897 9196 2903
rect 9892 2877 10003 2883
rect 5444 2857 6588 2863
rect 3364 2817 8027 2823
rect 9997 2823 10003 2877
rect 9997 2817 10035 2823
rect 3428 2797 3451 2803
rect 6500 2797 6956 2803
rect 9060 2797 10011 2803
rect 10029 2783 10035 2817
rect 10021 2777 10035 2783
rect 3060 2737 3067 2743
rect 1908 2717 4812 2723
rect 8452 2717 10540 2723
rect 3476 2697 3483 2703
rect 4436 2697 4700 2703
rect 4805 2697 4812 2703
rect 3077 2677 3276 2683
rect 4772 2677 4795 2683
rect 8228 2677 8364 2683
rect 10021 2617 10044 2623
rect 3844 2597 3867 2603
rect 4772 2597 4795 2603
rect 5652 2597 5819 2603
rect 8324 2597 9740 2603
rect 2852 2537 5132 2543
rect 8628 2537 10044 2543
rect 10660 2537 11084 2543
rect 8037 2517 9196 2523
rect 2484 2497 2844 2503
rect 8004 2497 9116 2503
rect 10692 2497 10924 2503
rect 10932 2497 11196 2503
rect 11204 2497 11308 2503
rect 4372 2477 4460 2483
rect 4468 2477 5388 2483
rect 5396 2477 5404 2483
rect 8421 2477 8428 2483
rect 4996 2457 5020 2463
rect 9892 2437 10524 2443
rect 7796 2357 7852 2363
rect 5156 2337 5467 2343
rect 1828 2317 5884 2323
rect 8596 2317 8699 2323
rect 9252 2317 9371 2323
rect 4948 2297 6636 2303
rect 8020 2297 8027 2303
rect 3348 2177 3387 2183
rect 3397 2177 3867 2183
rect 3877 2177 4924 2183
rect 9988 2157 10011 2163
rect 2468 2117 2540 2123
rect 3492 2117 5148 2123
rect 6053 2117 7387 2123
rect 7397 2117 7836 2123
rect 8708 2117 10140 2123
rect 1828 2097 2876 2103
rect 2884 2097 3932 2103
rect 4420 2097 4796 2103
rect 5348 2097 5467 2103
rect 9252 2097 9339 2103
rect 5796 2037 8300 2043
rect 8308 2037 8699 2043
rect 6388 1997 7196 2003
rect 5780 1957 6636 1963
rect 2749 1937 2764 1943
rect 1573 1917 1644 1923
rect 2749 1923 2755 1937
rect 2772 1937 3996 1943
rect 7236 1937 9036 1943
rect 9061 1937 9196 1943
rect 10021 1937 11004 1943
rect 1652 1917 2755 1923
rect 3332 1917 3451 1923
rect 3461 1917 3964 1923
rect 3988 1917 5644 1923
rect 8676 1917 11196 1923
rect 11204 1917 11323 1923
rect 9093 1897 9132 1903
rect 3476 1877 5228 1883
rect 5284 1877 11932 1883
rect 2612 1857 4044 1863
rect 6404 1797 6427 1803
rect 3540 1777 6732 1783
rect 4517 1757 4540 1763
rect 6068 1737 6636 1743
rect 3124 1717 3628 1723
rect 9349 1717 11804 1723
rect 11812 1717 11884 1723
rect 3877 1697 3900 1703
rect 7780 1697 10268 1703
rect 11333 1697 11836 1703
rect 5972 1677 6043 1683
rect 3844 1637 3884 1643
rect 3892 1637 6043 1643
rect 3428 1597 3451 1603
rect 2228 1537 2460 1543
rect 6452 1537 9324 1543
rect 9332 1537 11132 1543
rect 1444 1517 2364 1523
rect 2372 1517 2748 1523
rect 2756 1517 2876 1523
rect 4660 1517 7619 1523
rect 1172 1497 2332 1503
rect 7613 1503 7619 1517
rect 7613 1497 8220 1503
rect 10644 1497 11084 1503
rect 8068 1477 9052 1483
rect 5477 1437 6348 1443
rect 6356 1437 6540 1443
rect 2885 1417 3228 1423
rect 5828 1317 9244 1323
rect 11828 1317 11884 1323
rect 7300 1297 7419 1303
rect 10004 1297 11836 1303
rect 9220 1277 9307 1283
rect 11140 1197 11212 1203
rect 3156 1117 3388 1123
rect 5029 1117 5132 1123
rect 11172 1117 11244 1123
rect 4084 1097 5180 1103
rect 5188 1097 5612 1103
rect 6484 1097 8476 1103
rect 7572 1077 8588 1083
rect 900 1037 1580 1043
rect 1588 1037 2572 1043
rect 4004 937 6796 943
rect 6820 937 8380 943
rect 6053 917 6092 923
rect 132 897 156 903
rect 1204 897 1563 903
rect 2212 897 2748 903
rect 2756 897 2860 903
rect 4420 897 4507 903
rect 7028 897 8524 903
rect 3860 877 4684 883
rect 884 837 1564 843
rect 2180 797 2732 803
rect 2740 797 2828 803
rect 6036 737 6043 743
rect 772 717 844 723
rect 9044 717 10540 723
rect 9684 677 10332 683
rect 1284 557 1564 563
rect 5076 537 5660 543
rect 1540 517 1563 523
rect 2084 517 2220 523
rect 9076 517 11084 523
rect 6084 497 7564 503
rect 7572 497 7660 503
rect 5172 457 6043 463
rect 5988 437 6044 443
rect 6100 437 6684 443
rect 6916 397 7404 403
rect 5668 357 5996 363
rect 5140 337 6620 343
rect 788 317 844 323
rect 852 317 1404 323
rect 2468 317 3628 323
rect 5972 317 6012 323
rect 6020 317 6043 323
rect 5828 297 6748 303
rect 5972 277 7948 283
rect 6692 137 8924 143
rect 5956 117 7948 123
rect 1764 97 1820 103
rect 1828 97 2220 103
rect 6052 97 9196 103
rect 9204 97 9244 103
<< m6contact >>
rect 10011 8895 10021 8905
rect 1691 8715 1701 8725
rect 9371 8495 9381 8505
rect 10363 8255 10373 8265
rect 4827 8095 4837 8105
rect 9339 8095 9349 8105
rect 3227 7924 3237 7925
rect 3227 7916 3228 7924
rect 3228 7916 3236 7924
rect 3236 7916 3237 7924
rect 3227 7915 3237 7916
rect 5403 7915 5413 7925
rect 10683 7724 10693 7725
rect 10683 7716 10684 7724
rect 10684 7716 10692 7724
rect 10692 7716 10693 7724
rect 10683 7715 10693 7716
rect 9339 7695 9349 7705
rect 10651 7695 10661 7705
rect 2843 7495 2853 7505
rect 10683 7295 10693 7305
rect 9371 6995 9381 7005
rect 2875 6875 2885 6885
rect 10683 6804 10693 6805
rect 10683 6796 10684 6804
rect 10684 6796 10692 6804
rect 10692 6796 10693 6804
rect 10683 6795 10693 6796
rect 10683 6735 10693 6745
rect 2779 6695 2789 6705
rect 10011 6684 10021 6685
rect 10011 6676 10012 6684
rect 10012 6676 10020 6684
rect 10020 6676 10021 6684
rect 10011 6675 10021 6676
rect 8731 6635 8741 6645
rect 7419 6595 7429 6605
rect 1915 6535 1925 6545
rect 10331 6544 10341 6545
rect 10331 6536 10332 6544
rect 10332 6536 10340 6544
rect 10340 6536 10341 6544
rect 10331 6535 10341 6536
rect 6747 6515 6757 6525
rect 10395 6515 10405 6525
rect 1915 6495 1925 6505
rect 8027 6475 8037 6485
rect 10203 6475 10213 6485
rect 2779 6115 2789 6125
rect 9339 6095 9349 6105
rect 635 5915 645 5925
rect 8859 5895 8869 5905
rect 11291 5895 11301 5905
rect 8699 5875 8709 5885
rect 8027 5715 8037 5725
rect 9371 5715 9381 5725
rect 8731 5695 8741 5705
rect 6779 5675 6789 5685
rect 5019 5595 5029 5605
rect 8699 5595 8709 5605
rect 11291 5595 11301 5605
rect 635 5535 645 5545
rect 10331 5544 10341 5545
rect 10331 5536 10332 5544
rect 10332 5536 10340 5544
rect 10340 5536 10341 5544
rect 10331 5535 10341 5536
rect 8059 5515 8069 5525
rect 9371 5515 9381 5525
rect 1947 5495 1957 5505
rect 6747 5495 6757 5505
rect 1691 5395 1701 5405
rect 10395 5335 10405 5345
rect 4731 5315 4741 5325
rect 7387 5315 7397 5325
rect 10203 5315 10213 5325
rect 10619 5315 10629 5325
rect 8059 5115 8069 5125
rect 4731 5095 4741 5105
rect 6427 5095 6437 5105
rect 6747 5095 6757 5105
rect 10651 5095 10661 5105
rect 1915 4955 1925 4965
rect 8699 4964 8709 4965
rect 8699 4956 8700 4964
rect 8700 4956 8708 4964
rect 8708 4956 8709 4964
rect 8699 4955 8709 4956
rect 9339 4855 9349 4865
rect 1275 4775 1285 4785
rect 3227 4724 3237 4725
rect 3227 4716 3228 4724
rect 3228 4716 3236 4724
rect 3236 4716 3237 4724
rect 3227 4715 3237 4716
rect 3387 4715 3397 4725
rect 3483 4695 3493 4705
rect 1755 4615 1765 4625
rect 10363 4535 10373 4545
rect 1275 4515 1285 4525
rect 1755 4515 1765 4525
rect 3483 4515 3493 4525
rect 4155 4475 4165 4485
rect 5403 4475 5413 4485
rect 9339 4475 9349 4485
rect 3323 4415 3333 4425
rect 8859 4415 8869 4425
rect 3227 4344 3237 4345
rect 3227 4336 3228 4344
rect 3228 4336 3236 4344
rect 3236 4336 3237 4344
rect 3227 4335 3237 4336
rect 5179 4335 5189 4345
rect 5819 4295 5829 4305
rect 6779 4295 6789 4305
rect 10363 4295 10373 4305
rect 4155 4264 4165 4265
rect 4155 4256 4156 4264
rect 4156 4256 4164 4264
rect 4164 4256 4165 4264
rect 4155 4255 4165 4256
rect 5179 4135 5189 4145
rect 10363 4175 10373 4185
rect 8411 4095 8421 4105
rect 5019 4075 5029 4085
rect 10011 4075 10021 4085
rect 3451 4055 3461 4065
rect 7419 4055 7429 4065
rect 5019 4015 5029 4025
rect 10651 4015 10661 4025
rect 8059 3995 8069 4005
rect 7387 3975 7397 3985
rect 8059 3975 8069 3985
rect 3867 3955 3877 3965
rect 10395 3915 10405 3925
rect 8635 3855 8645 3865
rect 8699 3744 8709 3745
rect 8699 3736 8700 3744
rect 8700 3736 8708 3744
rect 8708 3736 8709 3744
rect 8699 3735 8709 3736
rect 7419 3715 7429 3725
rect 8635 3715 8645 3725
rect 7387 3704 7397 3705
rect 7387 3696 7388 3704
rect 7388 3696 7396 3704
rect 7396 3696 7397 3704
rect 7387 3695 7397 3696
rect 9947 3695 9957 3705
rect 7387 3675 7397 3685
rect 8027 3655 8037 3665
rect 10619 3635 10629 3645
rect 9083 3515 9093 3525
rect 1915 3495 1925 3505
rect 4795 3495 4805 3505
rect 10395 3504 10405 3505
rect 10395 3496 10396 3504
rect 10396 3496 10404 3504
rect 10404 3496 10405 3504
rect 10395 3495 10405 3496
rect 3227 3455 3237 3465
rect 8059 3435 8069 3445
rect 8635 3435 8645 3445
rect 9051 3375 9061 3385
rect 2843 3335 2853 3345
rect 9947 3295 9957 3305
rect 4827 3264 4837 3265
rect 4827 3256 4828 3264
rect 4828 3256 4836 3264
rect 4836 3256 4837 3264
rect 4827 3255 4837 3256
rect 7387 3115 7397 3125
rect 9307 3115 9317 3125
rect 3323 2915 3333 2925
rect 4795 2915 4805 2925
rect 7387 2915 7397 2925
rect 8635 2895 8645 2905
rect 8027 2815 8037 2825
rect 3451 2795 3461 2805
rect 10011 2795 10021 2805
rect 10011 2775 10021 2785
rect 3067 2735 3077 2745
rect 3483 2695 3493 2705
rect 4795 2695 4805 2705
rect 3067 2675 3077 2685
rect 4795 2675 4805 2685
rect 10011 2615 10021 2625
rect 3867 2595 3877 2605
rect 4795 2595 4805 2605
rect 5819 2595 5829 2605
rect 8027 2515 8037 2525
rect 8411 2475 8421 2485
rect 5467 2335 5477 2345
rect 8699 2315 8709 2325
rect 9371 2315 9381 2325
rect 8027 2295 8037 2305
rect 3387 2175 3397 2185
rect 3867 2175 3877 2185
rect 10011 2155 10021 2165
rect 6043 2115 6053 2125
rect 7387 2115 7397 2125
rect 5467 2095 5477 2105
rect 9339 2095 9349 2105
rect 8699 2035 8709 2045
rect 1947 1944 1957 1945
rect 1947 1936 1948 1944
rect 1948 1936 1956 1944
rect 1956 1936 1957 1944
rect 1947 1935 1957 1936
rect 1563 1915 1573 1925
rect 9051 1935 9061 1945
rect 10011 1935 10021 1945
rect 3451 1915 3461 1925
rect 11323 1915 11333 1925
rect 9083 1895 9093 1905
rect 6427 1795 6437 1805
rect 4507 1755 4517 1765
rect 9339 1715 9349 1725
rect 3867 1695 3877 1705
rect 11323 1695 11333 1705
rect 6043 1675 6053 1685
rect 6043 1644 6053 1645
rect 6043 1636 6044 1644
rect 6044 1636 6052 1644
rect 6052 1636 6053 1644
rect 6043 1635 6053 1636
rect 3451 1595 3461 1605
rect 9051 1504 9061 1505
rect 9051 1496 9052 1504
rect 9052 1496 9060 1504
rect 9060 1496 9061 1504
rect 9051 1495 9061 1496
rect 5467 1435 5477 1445
rect 2875 1415 2885 1425
rect 7419 1295 7429 1305
rect 9307 1275 9317 1285
rect 5019 1115 5029 1125
rect 9051 1124 9061 1125
rect 9051 1116 9052 1124
rect 9052 1116 9060 1124
rect 9060 1116 9061 1124
rect 9051 1115 9061 1116
rect 6043 915 6053 925
rect 1563 895 1573 905
rect 4507 895 4517 905
rect 6043 735 6053 745
rect 1563 515 1573 525
rect 6043 455 6053 465
rect 6043 315 6053 325
<< metal6 >>
rect 635 5545 645 5915
rect 1691 5405 1701 8715
rect 1915 6505 1925 6535
rect 1915 4965 1925 6495
rect 2779 6125 2789 6695
rect 1275 4525 1285 4775
rect 1755 4525 1765 4615
rect 1915 3505 1925 4955
rect 1947 1945 1957 5495
rect 2843 3345 2853 7495
rect 1563 905 1573 1915
rect 2875 1425 2885 6875
rect 3227 4725 3237 7915
rect 4731 5105 4741 5315
rect 3227 3465 3237 4335
rect 3323 2925 3333 4415
rect 3067 2685 3077 2735
rect 3387 2185 3397 4715
rect 3483 4525 3493 4695
rect 3451 2805 3461 4055
rect 3483 2705 3493 4515
rect 4155 4265 4165 4475
rect 3867 2605 3877 3955
rect 4795 2925 4805 3495
rect 4827 3265 4837 8095
rect 5019 4085 5029 5595
rect 5403 4485 5413 7915
rect 9339 7705 9349 8095
rect 6747 5505 6757 6515
rect 6747 5105 6757 5495
rect 5179 4145 5189 4335
rect 4795 2705 4805 2915
rect 4795 2605 4805 2675
rect 3451 1605 3461 1915
rect 3867 1705 3877 2175
rect 4507 905 4517 1755
rect 5019 1125 5029 4015
rect 5819 2605 5829 4295
rect 5467 2105 5477 2335
rect 5467 1445 5477 2095
rect 6043 1685 6053 2115
rect 6427 1805 6437 5095
rect 6779 4305 6789 5675
rect 7387 3985 7397 5315
rect 7419 4065 7429 6595
rect 8027 5725 8037 6475
rect 7387 3705 7397 3975
rect 7387 3125 7397 3675
rect 7387 2125 7397 2915
rect 6043 1645 6053 1675
rect 7419 1305 7429 3715
rect 8027 3665 8037 5715
rect 8699 5605 8709 5875
rect 8731 5705 8741 6635
rect 9339 6105 9349 7695
rect 9371 7005 9381 8495
rect 10011 6685 10021 8895
rect 8059 5125 8069 5515
rect 8059 4005 8069 5115
rect 8059 3445 8069 3975
rect 8027 2525 8037 2815
rect 8027 2305 8037 2515
rect 8411 2485 8421 4095
rect 8635 3725 8645 3855
rect 8699 3745 8709 4955
rect 8859 4425 8869 5895
rect 9339 4865 9349 6095
rect 9371 5525 9381 5715
rect 8635 2905 8645 3435
rect 8699 2045 8709 2315
rect 9051 1945 9061 3375
rect 9083 1905 9093 3515
rect 9051 1125 9061 1495
rect 9307 1285 9317 3115
rect 9339 2105 9349 4475
rect 9371 2325 9381 5515
rect 10203 5325 10213 6475
rect 10331 5545 10341 6535
rect 10363 4545 10373 8255
rect 10395 5345 10405 6515
rect 10363 4185 10373 4295
rect 9947 3305 9957 3695
rect 10011 2805 10021 4075
rect 10395 3925 10405 5335
rect 10395 3505 10405 3915
rect 10619 3645 10629 5315
rect 10651 5105 10661 7695
rect 10683 7305 10693 7715
rect 10683 6745 10693 6795
rect 11291 5605 11301 5895
rect 10651 4025 10661 5095
rect 10011 2625 10021 2775
rect 9339 1725 9349 2095
rect 10011 1945 10021 2155
rect 11323 1705 11333 1915
rect 1563 525 1573 895
rect 6043 745 6053 915
rect 6043 465 6053 735
rect 6043 325 6053 455
use SECLIBAND_opt  SECLIBAND_opt_50
timestamp 1602073617
transform 1 0 8 0 -1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_1
timestamp 1602073617
transform 1 0 8 0 1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_51
timestamp 1602073617
transform -1 0 1308 0 -1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_12
timestamp 1602073617
transform 1 0 658 0 1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_30
timestamp 1602073617
transform -1 0 1958 0 -1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_3
timestamp 1602073617
transform 1 0 1308 0 1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_751
timestamp 1602073617
transform 1 0 1958 0 -1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_749
timestamp 1602073617
transform -1 0 2608 0 1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_789
timestamp 1602073617
transform 1 0 2608 0 -1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_752
timestamp 1602073617
transform 1 0 2608 0 1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_793
timestamp 1602073617
transform 1 0 3258 0 -1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_748
timestamp 1602073617
transform -1 0 3908 0 1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_790
timestamp 1602073617
transform -1 0 4558 0 -1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_621
timestamp 1602073617
transform 1 0 3908 0 1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_753
timestamp 1602073617
transform -1 0 5208 0 -1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_616
timestamp 1602073617
transform -1 0 5208 0 1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_816
timestamp 1602073617
transform 1 0 5208 0 -1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_754
timestamp 1602073617
transform -1 0 5858 0 1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_381
timestamp 1602073617
transform 1 0 5858 0 -1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_14
timestamp 1602073617
transform 1 0 5858 0 1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_817
timestamp 1602073617
transform -1 0 7158 0 -1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_847
timestamp 1602073617
transform 1 0 6508 0 1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_815
timestamp 1602073617
transform 1 0 7158 0 -1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_619
timestamp 1602073617
transform 1 0 7158 0 1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_846
timestamp 1602073617
transform 1 0 7808 0 -1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_622
timestamp 1602073617
transform 1 0 7808 0 1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_848
timestamp 1602073617
transform 1 0 8458 0 -1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_624
timestamp 1602073617
transform 1 0 8458 0 1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_529
timestamp 1602073617
transform 1 0 9108 0 -1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_693
timestamp 1602073617
transform 1 0 9108 0 1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_548
timestamp 1602073617
transform 1 0 9758 0 -1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_530
timestamp 1602073617
transform -1 0 10408 0 1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_531
timestamp 1602073617
transform 1 0 10408 0 -1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_713
timestamp 1602073617
transform -1 0 11058 0 1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_549
timestamp 1602073617
transform 1 0 11058 0 -1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_705
timestamp 1602073617
transform -1 0 11708 0 1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_348
timestamp 1602073617
transform -1 0 12358 0 -1 210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_565
timestamp 1602073617
transform 1 0 11708 0 1 210
box -4 -6 618 206
use FILL  FILL_2_1
timestamp 1602073617
transform 1 0 12358 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1
timestamp 1602073617
transform -1 0 12374 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_4
timestamp 1602073617
transform 1 0 12406 0 1 210
box -4 -6 20 206
use FILL  FILL_2_3
timestamp 1602073617
transform 1 0 12390 0 1 210
box -4 -6 20 206
use FILL  FILL_2_2
timestamp 1602073617
transform 1 0 12374 0 1 210
box -4 -6 20 206
use FILL  FILL_1_4
timestamp 1602073617
transform -1 0 12422 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_3
timestamp 1602073617
transform -1 0 12406 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_2
timestamp 1602073617
transform -1 0 12390 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_7
timestamp 1602073617
transform 1 0 12454 0 1 210
box -4 -6 20 206
use FILL  FILL_2_6
timestamp 1602073617
transform 1 0 12438 0 1 210
box -4 -6 20 206
use FILL  FILL_2_5
timestamp 1602073617
transform 1 0 12422 0 1 210
box -4 -6 20 206
use FILL  FILL_1_7
timestamp 1602073617
transform -1 0 12470 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_6
timestamp 1602073617
transform -1 0 12454 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_5
timestamp 1602073617
transform -1 0 12438 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_8
timestamp 1602073617
transform 1 0 12470 0 1 210
box -4 -6 20 206
use FILL  FILL_1_8
timestamp 1602073617
transform -1 0 12486 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_10
timestamp 1602073617
transform 1 0 12502 0 1 210
box -4 -6 20 206
use FILL  FILL_2_9
timestamp 1602073617
transform 1 0 12486 0 1 210
box -4 -6 20 206
use FILL  FILL_1_10
timestamp 1602073617
transform -1 0 12518 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_9
timestamp 1602073617
transform -1 0 12502 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_11
timestamp 1602073617
transform 1 0 12518 0 1 210
box -4 -6 20 206
use FILL  FILL_1_11
timestamp 1602073617
transform -1 0 12534 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_13
timestamp 1602073617
transform 1 0 12550 0 1 210
box -4 -6 20 206
use FILL  FILL_2_12
timestamp 1602073617
transform 1 0 12534 0 1 210
box -4 -6 20 206
use FILL  FILL_1_13
timestamp 1602073617
transform -1 0 12566 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_12
timestamp 1602073617
transform -1 0 12550 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_14
timestamp 1602073617
transform 1 0 12566 0 1 210
box -4 -6 20 206
use FILL  FILL_1_14
timestamp 1602073617
transform -1 0 12582 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_16
timestamp 1602073617
transform 1 0 12598 0 1 210
box -4 -6 20 206
use FILL  FILL_2_15
timestamp 1602073617
transform 1 0 12582 0 1 210
box -4 -6 20 206
use FILL  FILL_1_16
timestamp 1602073617
transform -1 0 12614 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_15
timestamp 1602073617
transform -1 0 12598 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_17
timestamp 1602073617
transform 1 0 12614 0 1 210
box -4 -6 20 206
use FILL  FILL_1_17
timestamp 1602073617
transform -1 0 12630 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_19
timestamp 1602073617
transform 1 0 12646 0 1 210
box -4 -6 20 206
use FILL  FILL_2_18
timestamp 1602073617
transform 1 0 12630 0 1 210
box -4 -6 20 206
use FILL  FILL_1_19
timestamp 1602073617
transform -1 0 12662 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_18
timestamp 1602073617
transform -1 0 12646 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_21
timestamp 1602073617
transform 1 0 12678 0 1 210
box -4 -6 20 206
use FILL  FILL_2_20
timestamp 1602073617
transform 1 0 12662 0 1 210
box -4 -6 20 206
use FILL  FILL_1_21
timestamp 1602073617
transform -1 0 12694 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_20
timestamp 1602073617
transform -1 0 12678 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_22
timestamp 1602073617
transform 1 0 12694 0 1 210
box -4 -6 20 206
use FILL  FILL_1_22
timestamp 1602073617
transform -1 0 12710 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_24
timestamp 1602073617
transform 1 0 12726 0 1 210
box -4 -6 20 206
use FILL  FILL_2_23
timestamp 1602073617
transform 1 0 12710 0 1 210
box -4 -6 20 206
use FILL  FILL_1_24
timestamp 1602073617
transform -1 0 12742 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_23
timestamp 1602073617
transform -1 0 12726 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_25
timestamp 1602073617
transform 1 0 12742 0 1 210
box -4 -6 20 206
use FILL  FILL_1_25
timestamp 1602073617
transform -1 0 12758 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_27
timestamp 1602073617
transform 1 0 12774 0 1 210
box -4 -6 20 206
use FILL  FILL_2_26
timestamp 1602073617
transform 1 0 12758 0 1 210
box -4 -6 20 206
use FILL  FILL_1_27
timestamp 1602073617
transform -1 0 12790 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_26
timestamp 1602073617
transform -1 0 12774 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_28
timestamp 1602073617
transform 1 0 12790 0 1 210
box -4 -6 20 206
use FILL  FILL_1_28
timestamp 1602073617
transform -1 0 12806 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_30
timestamp 1602073617
transform 1 0 12822 0 1 210
box -4 -6 20 206
use FILL  FILL_2_29
timestamp 1602073617
transform 1 0 12806 0 1 210
box -4 -6 20 206
use FILL  FILL_1_30
timestamp 1602073617
transform -1 0 12838 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_29
timestamp 1602073617
transform -1 0 12822 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_31
timestamp 1602073617
transform 1 0 12838 0 1 210
box -4 -6 20 206
use FILL  FILL_1_31
timestamp 1602073617
transform -1 0 12854 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_33
timestamp 1602073617
transform 1 0 12870 0 1 210
box -4 -6 20 206
use FILL  FILL_2_32
timestamp 1602073617
transform 1 0 12854 0 1 210
box -4 -6 20 206
use FILL  FILL_1_33
timestamp 1602073617
transform -1 0 12886 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_32
timestamp 1602073617
transform -1 0 12870 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_34
timestamp 1602073617
transform 1 0 12886 0 1 210
box -4 -6 20 206
use FILL  FILL_1_34
timestamp 1602073617
transform -1 0 12902 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_36
timestamp 1602073617
transform 1 0 12918 0 1 210
box -4 -6 20 206
use FILL  FILL_2_35
timestamp 1602073617
transform 1 0 12902 0 1 210
box -4 -6 20 206
use FILL  FILL_1_36
timestamp 1602073617
transform -1 0 12934 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_35
timestamp 1602073617
transform -1 0 12918 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_37
timestamp 1602073617
transform 1 0 12934 0 1 210
box -4 -6 20 206
use FILL  FILL_1_37
timestamp 1602073617
transform -1 0 12950 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_39
timestamp 1602073617
transform 1 0 12966 0 1 210
box -4 -6 20 206
use FILL  FILL_2_38
timestamp 1602073617
transform 1 0 12950 0 1 210
box -4 -6 20 206
use FILL  FILL_1_39
timestamp 1602073617
transform -1 0 12982 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_38
timestamp 1602073617
transform -1 0 12966 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_40
timestamp 1602073617
transform 1 0 12982 0 1 210
box -4 -6 20 206
use FILL  FILL_1_40
timestamp 1602073617
transform -1 0 12998 0 -1 210
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_587
timestamp 1602073617
transform 1 0 8 0 -1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_31
timestamp 1602073617
transform 1 0 658 0 -1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_750
timestamp 1602073617
transform 1 0 1308 0 -1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_425
timestamp 1602073617
transform 1 0 1958 0 -1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_756
timestamp 1602073617
transform 1 0 2608 0 -1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_4
timestamp 1602073617
transform 1 0 3258 0 -1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_104
timestamp 1602073617
transform 1 0 3908 0 -1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_8
timestamp 1602073617
transform -1 0 5208 0 -1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_671
timestamp 1602073617
transform 1 0 5208 0 -1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_672
timestamp 1602073617
transform 1 0 5858 0 -1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_618
timestamp 1602073617
transform 1 0 6508 0 -1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_699
timestamp 1602073617
transform -1 0 7808 0 -1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_814
timestamp 1602073617
transform -1 0 8458 0 -1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_110
timestamp 1602073617
transform 1 0 8458 0 -1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_859
timestamp 1602073617
transform 1 0 9108 0 -1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_692
timestamp 1602073617
transform 1 0 9758 0 -1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_706
timestamp 1602073617
transform 1 0 10408 0 -1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_526
timestamp 1602073617
transform 1 0 11058 0 -1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_550
timestamp 1602073617
transform 1 0 11708 0 -1 610
box -4 -6 618 206
use FILL  FILL_3_1
timestamp 1602073617
transform -1 0 12374 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_2
timestamp 1602073617
transform -1 0 12390 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_3
timestamp 1602073617
transform -1 0 12406 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_4
timestamp 1602073617
transform -1 0 12422 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_5
timestamp 1602073617
transform -1 0 12438 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_6
timestamp 1602073617
transform -1 0 12454 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_7
timestamp 1602073617
transform -1 0 12470 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_8
timestamp 1602073617
transform -1 0 12486 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_10
timestamp 1602073617
transform -1 0 12518 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_9
timestamp 1602073617
transform -1 0 12502 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_11
timestamp 1602073617
transform -1 0 12534 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_13
timestamp 1602073617
transform -1 0 12566 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_12
timestamp 1602073617
transform -1 0 12550 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_14
timestamp 1602073617
transform -1 0 12582 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_16
timestamp 1602073617
transform -1 0 12614 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_15
timestamp 1602073617
transform -1 0 12598 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_17
timestamp 1602073617
transform -1 0 12630 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_19
timestamp 1602073617
transform -1 0 12662 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_18
timestamp 1602073617
transform -1 0 12646 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_21
timestamp 1602073617
transform -1 0 12694 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_20
timestamp 1602073617
transform -1 0 12678 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_22
timestamp 1602073617
transform -1 0 12710 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_24
timestamp 1602073617
transform -1 0 12742 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_23
timestamp 1602073617
transform -1 0 12726 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_25
timestamp 1602073617
transform -1 0 12758 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_27
timestamp 1602073617
transform -1 0 12790 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_26
timestamp 1602073617
transform -1 0 12774 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_28
timestamp 1602073617
transform -1 0 12806 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_30
timestamp 1602073617
transform -1 0 12838 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_29
timestamp 1602073617
transform -1 0 12822 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_31
timestamp 1602073617
transform -1 0 12854 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_33
timestamp 1602073617
transform -1 0 12886 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_32
timestamp 1602073617
transform -1 0 12870 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_34
timestamp 1602073617
transform -1 0 12902 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_36
timestamp 1602073617
transform -1 0 12934 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_35
timestamp 1602073617
transform -1 0 12918 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_37
timestamp 1602073617
transform -1 0 12950 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_39
timestamp 1602073617
transform -1 0 12982 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_38
timestamp 1602073617
transform -1 0 12966 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_40
timestamp 1602073617
transform -1 0 12998 0 -1 610
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_17
timestamp 1602073617
transform 1 0 8 0 1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_36
timestamp 1602073617
transform 1 0 658 0 1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_22
timestamp 1602073617
transform 1 0 1308 0 1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_2
timestamp 1602073617
transform 1 0 1958 0 1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_157
timestamp 1602073617
transform 1 0 2608 0 1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_757
timestamp 1602073617
transform 1 0 3258 0 1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_818
timestamp 1602073617
transform 1 0 3908 0 1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_820
timestamp 1602073617
transform 1 0 4558 0 1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_414
timestamp 1602073617
transform -1 0 5858 0 1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_5
timestamp 1602073617
transform 1 0 5858 0 1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_28
timestamp 1602073617
transform -1 0 7158 0 1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_382
timestamp 1602073617
transform 1 0 7158 0 1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_225
timestamp 1602073617
transform 1 0 7808 0 1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_260
timestamp 1602073617
transform 1 0 8458 0 1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_615
timestamp 1602073617
transform 1 0 9108 0 1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_623
timestamp 1602073617
transform -1 0 10408 0 1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_261
timestamp 1602073617
transform 1 0 10408 0 1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_485
timestamp 1602073617
transform 1 0 11058 0 1 610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_546
timestamp 1602073617
transform -1 0 12358 0 1 610
box -4 -6 618 206
use FILL  FILL_4_1
timestamp 1602073617
transform 1 0 12358 0 1 610
box -4 -6 20 206
use FILL  FILL_4_2
timestamp 1602073617
transform 1 0 12374 0 1 610
box -4 -6 20 206
use FILL  FILL_4_3
timestamp 1602073617
transform 1 0 12390 0 1 610
box -4 -6 20 206
use FILL  FILL_4_4
timestamp 1602073617
transform 1 0 12406 0 1 610
box -4 -6 20 206
use FILL  FILL_4_5
timestamp 1602073617
transform 1 0 12422 0 1 610
box -4 -6 20 206
use FILL  FILL_4_6
timestamp 1602073617
transform 1 0 12438 0 1 610
box -4 -6 20 206
use FILL  FILL_4_7
timestamp 1602073617
transform 1 0 12454 0 1 610
box -4 -6 20 206
use FILL  FILL_4_8
timestamp 1602073617
transform 1 0 12470 0 1 610
box -4 -6 20 206
use FILL  FILL_4_10
timestamp 1602073617
transform 1 0 12502 0 1 610
box -4 -6 20 206
use FILL  FILL_4_9
timestamp 1602073617
transform 1 0 12486 0 1 610
box -4 -6 20 206
use FILL  FILL_4_11
timestamp 1602073617
transform 1 0 12518 0 1 610
box -4 -6 20 206
use FILL  FILL_4_13
timestamp 1602073617
transform 1 0 12550 0 1 610
box -4 -6 20 206
use FILL  FILL_4_12
timestamp 1602073617
transform 1 0 12534 0 1 610
box -4 -6 20 206
use FILL  FILL_4_14
timestamp 1602073617
transform 1 0 12566 0 1 610
box -4 -6 20 206
use FILL  FILL_4_16
timestamp 1602073617
transform 1 0 12598 0 1 610
box -4 -6 20 206
use FILL  FILL_4_15
timestamp 1602073617
transform 1 0 12582 0 1 610
box -4 -6 20 206
use FILL  FILL_4_17
timestamp 1602073617
transform 1 0 12614 0 1 610
box -4 -6 20 206
use FILL  FILL_4_19
timestamp 1602073617
transform 1 0 12646 0 1 610
box -4 -6 20 206
use FILL  FILL_4_18
timestamp 1602073617
transform 1 0 12630 0 1 610
box -4 -6 20 206
use FILL  FILL_4_21
timestamp 1602073617
transform 1 0 12678 0 1 610
box -4 -6 20 206
use FILL  FILL_4_20
timestamp 1602073617
transform 1 0 12662 0 1 610
box -4 -6 20 206
use FILL  FILL_4_22
timestamp 1602073617
transform 1 0 12694 0 1 610
box -4 -6 20 206
use FILL  FILL_4_24
timestamp 1602073617
transform 1 0 12726 0 1 610
box -4 -6 20 206
use FILL  FILL_4_23
timestamp 1602073617
transform 1 0 12710 0 1 610
box -4 -6 20 206
use FILL  FILL_4_25
timestamp 1602073617
transform 1 0 12742 0 1 610
box -4 -6 20 206
use FILL  FILL_4_27
timestamp 1602073617
transform 1 0 12774 0 1 610
box -4 -6 20 206
use FILL  FILL_4_26
timestamp 1602073617
transform 1 0 12758 0 1 610
box -4 -6 20 206
use FILL  FILL_4_28
timestamp 1602073617
transform 1 0 12790 0 1 610
box -4 -6 20 206
use FILL  FILL_4_30
timestamp 1602073617
transform 1 0 12822 0 1 610
box -4 -6 20 206
use FILL  FILL_4_29
timestamp 1602073617
transform 1 0 12806 0 1 610
box -4 -6 20 206
use FILL  FILL_4_31
timestamp 1602073617
transform 1 0 12838 0 1 610
box -4 -6 20 206
use FILL  FILL_4_33
timestamp 1602073617
transform 1 0 12870 0 1 610
box -4 -6 20 206
use FILL  FILL_4_32
timestamp 1602073617
transform 1 0 12854 0 1 610
box -4 -6 20 206
use FILL  FILL_4_34
timestamp 1602073617
transform 1 0 12886 0 1 610
box -4 -6 20 206
use FILL  FILL_4_36
timestamp 1602073617
transform 1 0 12918 0 1 610
box -4 -6 20 206
use FILL  FILL_4_35
timestamp 1602073617
transform 1 0 12902 0 1 610
box -4 -6 20 206
use FILL  FILL_4_37
timestamp 1602073617
transform 1 0 12934 0 1 610
box -4 -6 20 206
use FILL  FILL_4_39
timestamp 1602073617
transform 1 0 12966 0 1 610
box -4 -6 20 206
use FILL  FILL_4_38
timestamp 1602073617
transform 1 0 12950 0 1 610
box -4 -6 20 206
use FILL  FILL_4_40
timestamp 1602073617
transform 1 0 12982 0 1 610
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_429
timestamp 1602073617
transform 1 0 8 0 -1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_430
timestamp 1602073617
transform -1 0 1308 0 -1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_44
timestamp 1602073617
transform 1 0 1308 0 -1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_386
timestamp 1602073617
transform 1 0 1958 0 -1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_18
timestamp 1602073617
transform 1 0 2608 0 -1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_143
timestamp 1602073617
transform -1 0 3908 0 -1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_133
timestamp 1602073617
transform -1 0 4558 0 -1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_791
timestamp 1602073617
transform 1 0 4558 0 -1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_185
timestamp 1602073617
transform -1 0 5858 0 -1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_37
timestamp 1602073617
transform 1 0 5858 0 -1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_614
timestamp 1602073617
transform -1 0 7158 0 -1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_391
timestamp 1602073617
transform -1 0 7808 0 -1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_384
timestamp 1602073617
transform -1 0 8458 0 -1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_694
timestamp 1602073617
transform 1 0 8458 0 -1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_707
timestamp 1602073617
transform 1 0 9108 0 -1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_712
timestamp 1602073617
transform 1 0 9758 0 -1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_725
timestamp 1602073617
transform 1 0 10408 0 -1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_613
timestamp 1602073617
transform -1 0 11708 0 -1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_525
timestamp 1602073617
transform 1 0 11708 0 -1 1010
box -4 -6 618 206
use FILL  FILL_5_1
timestamp 1602073617
transform -1 0 12374 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_2
timestamp 1602073617
transform -1 0 12390 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_3
timestamp 1602073617
transform -1 0 12406 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_4
timestamp 1602073617
transform -1 0 12422 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_5
timestamp 1602073617
transform -1 0 12438 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_6
timestamp 1602073617
transform -1 0 12454 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_7
timestamp 1602073617
transform -1 0 12470 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_8
timestamp 1602073617
transform -1 0 12486 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_10
timestamp 1602073617
transform -1 0 12518 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_9
timestamp 1602073617
transform -1 0 12502 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_11
timestamp 1602073617
transform -1 0 12534 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_13
timestamp 1602073617
transform -1 0 12566 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_12
timestamp 1602073617
transform -1 0 12550 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_14
timestamp 1602073617
transform -1 0 12582 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_16
timestamp 1602073617
transform -1 0 12614 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_15
timestamp 1602073617
transform -1 0 12598 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_17
timestamp 1602073617
transform -1 0 12630 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_19
timestamp 1602073617
transform -1 0 12662 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_18
timestamp 1602073617
transform -1 0 12646 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_21
timestamp 1602073617
transform -1 0 12694 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_20
timestamp 1602073617
transform -1 0 12678 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_22
timestamp 1602073617
transform -1 0 12710 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_24
timestamp 1602073617
transform -1 0 12742 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_23
timestamp 1602073617
transform -1 0 12726 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_25
timestamp 1602073617
transform -1 0 12758 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_27
timestamp 1602073617
transform -1 0 12790 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_26
timestamp 1602073617
transform -1 0 12774 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_28
timestamp 1602073617
transform -1 0 12806 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_30
timestamp 1602073617
transform -1 0 12838 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_29
timestamp 1602073617
transform -1 0 12822 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_31
timestamp 1602073617
transform -1 0 12854 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_33
timestamp 1602073617
transform -1 0 12886 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_32
timestamp 1602073617
transform -1 0 12870 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_34
timestamp 1602073617
transform -1 0 12902 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_36
timestamp 1602073617
transform -1 0 12934 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_35
timestamp 1602073617
transform -1 0 12918 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_37
timestamp 1602073617
transform -1 0 12950 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_39
timestamp 1602073617
transform -1 0 12982 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_38
timestamp 1602073617
transform -1 0 12966 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_40
timestamp 1602073617
transform -1 0 12998 0 -1 1010
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_408
timestamp 1602073617
transform 1 0 8 0 1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_25
timestamp 1602073617
transform 1 0 658 0 1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_47
timestamp 1602073617
transform 1 0 1308 0 1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_11
timestamp 1602073617
transform 1 0 1958 0 1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_59
timestamp 1602073617
transform 1 0 2608 0 1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_666
timestamp 1602073617
transform 1 0 3258 0 1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_755
timestamp 1602073617
transform 1 0 3908 0 1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_664
timestamp 1602073617
transform -1 0 5208 0 1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_226
timestamp 1602073617
transform -1 0 5858 0 1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_6
timestamp 1602073617
transform 1 0 5858 0 1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_673
timestamp 1602073617
transform -1 0 7158 0 1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_670
timestamp 1602073617
transform -1 0 7808 0 1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_295
timestamp 1602073617
transform -1 0 8458 0 1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_255
timestamp 1602073617
transform 1 0 8458 0 1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_541
timestamp 1602073617
transform 1 0 9108 0 1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_708
timestamp 1602073617
transform -1 0 10408 0 1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_620
timestamp 1602073617
transform -1 0 11058 0 1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_528
timestamp 1602073617
transform 1 0 11058 0 1 1010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_486
timestamp 1602073617
transform -1 0 12358 0 1 1010
box -4 -6 618 206
use FILL  FILL_6_1
timestamp 1602073617
transform 1 0 12358 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_2
timestamp 1602073617
transform 1 0 12374 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_3
timestamp 1602073617
transform 1 0 12390 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_4
timestamp 1602073617
transform 1 0 12406 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_5
timestamp 1602073617
transform 1 0 12422 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_6
timestamp 1602073617
transform 1 0 12438 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_7
timestamp 1602073617
transform 1 0 12454 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_8
timestamp 1602073617
transform 1 0 12470 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_10
timestamp 1602073617
transform 1 0 12502 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_9
timestamp 1602073617
transform 1 0 12486 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_11
timestamp 1602073617
transform 1 0 12518 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_13
timestamp 1602073617
transform 1 0 12550 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_12
timestamp 1602073617
transform 1 0 12534 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_14
timestamp 1602073617
transform 1 0 12566 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_16
timestamp 1602073617
transform 1 0 12598 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_15
timestamp 1602073617
transform 1 0 12582 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_17
timestamp 1602073617
transform 1 0 12614 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_19
timestamp 1602073617
transform 1 0 12646 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_18
timestamp 1602073617
transform 1 0 12630 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_21
timestamp 1602073617
transform 1 0 12678 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_20
timestamp 1602073617
transform 1 0 12662 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_22
timestamp 1602073617
transform 1 0 12694 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_24
timestamp 1602073617
transform 1 0 12726 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_23
timestamp 1602073617
transform 1 0 12710 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_25
timestamp 1602073617
transform 1 0 12742 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_27
timestamp 1602073617
transform 1 0 12774 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_26
timestamp 1602073617
transform 1 0 12758 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_28
timestamp 1602073617
transform 1 0 12790 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_30
timestamp 1602073617
transform 1 0 12822 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_29
timestamp 1602073617
transform 1 0 12806 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_31
timestamp 1602073617
transform 1 0 12838 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_33
timestamp 1602073617
transform 1 0 12870 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_32
timestamp 1602073617
transform 1 0 12854 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_34
timestamp 1602073617
transform 1 0 12886 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_36
timestamp 1602073617
transform 1 0 12918 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_35
timestamp 1602073617
transform 1 0 12902 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_37
timestamp 1602073617
transform 1 0 12934 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_39
timestamp 1602073617
transform 1 0 12966 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_38
timestamp 1602073617
transform 1 0 12950 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_40
timestamp 1602073617
transform 1 0 12982 0 1 1010
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_762
timestamp 1602073617
transform 1 0 8 0 -1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_581
timestamp 1602073617
transform 1 0 658 0 -1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_26
timestamp 1602073617
transform 1 0 1308 0 -1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_95
timestamp 1602073617
transform -1 0 2608 0 -1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_40
timestamp 1602073617
transform 1 0 2608 0 -1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_719
timestamp 1602073617
transform -1 0 3908 0 -1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_665
timestamp 1602073617
transform -1 0 4558 0 -1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_227
timestamp 1602073617
transform -1 0 5208 0 -1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_819
timestamp 1602073617
transform -1 0 5858 0 -1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_792
timestamp 1602073617
transform 1 0 5858 0 -1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_805
timestamp 1602073617
transform 1 0 6508 0 -1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_292
timestamp 1602073617
transform 1 0 7158 0 -1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_346
timestamp 1602073617
transform 1 0 7808 0 -1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_272
timestamp 1602073617
transform -1 0 9108 0 -1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_695
timestamp 1602073617
transform 1 0 9108 0 -1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_696
timestamp 1602073617
transform 1 0 9758 0 -1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_527
timestamp 1602073617
transform 1 0 10408 0 -1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_547
timestamp 1602073617
transform 1 0 11058 0 -1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_484
timestamp 1602073617
transform 1 0 11708 0 -1 1410
box -4 -6 618 206
use FILL  FILL_7_1
timestamp 1602073617
transform -1 0 12374 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_2
timestamp 1602073617
transform -1 0 12390 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_3
timestamp 1602073617
transform -1 0 12406 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_4
timestamp 1602073617
transform -1 0 12422 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_5
timestamp 1602073617
transform -1 0 12438 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_6
timestamp 1602073617
transform -1 0 12454 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_7
timestamp 1602073617
transform -1 0 12470 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_8
timestamp 1602073617
transform -1 0 12486 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_10
timestamp 1602073617
transform -1 0 12518 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_9
timestamp 1602073617
transform -1 0 12502 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_11
timestamp 1602073617
transform -1 0 12534 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_13
timestamp 1602073617
transform -1 0 12566 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_12
timestamp 1602073617
transform -1 0 12550 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_14
timestamp 1602073617
transform -1 0 12582 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_16
timestamp 1602073617
transform -1 0 12614 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_15
timestamp 1602073617
transform -1 0 12598 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_17
timestamp 1602073617
transform -1 0 12630 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_19
timestamp 1602073617
transform -1 0 12662 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_18
timestamp 1602073617
transform -1 0 12646 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_21
timestamp 1602073617
transform -1 0 12694 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_20
timestamp 1602073617
transform -1 0 12678 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_22
timestamp 1602073617
transform -1 0 12710 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_24
timestamp 1602073617
transform -1 0 12742 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_23
timestamp 1602073617
transform -1 0 12726 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_25
timestamp 1602073617
transform -1 0 12758 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_27
timestamp 1602073617
transform -1 0 12790 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_26
timestamp 1602073617
transform -1 0 12774 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_28
timestamp 1602073617
transform -1 0 12806 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_30
timestamp 1602073617
transform -1 0 12838 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_29
timestamp 1602073617
transform -1 0 12822 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_31
timestamp 1602073617
transform -1 0 12854 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_33
timestamp 1602073617
transform -1 0 12886 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_32
timestamp 1602073617
transform -1 0 12870 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_34
timestamp 1602073617
transform -1 0 12902 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_36
timestamp 1602073617
transform -1 0 12934 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_35
timestamp 1602073617
transform -1 0 12918 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_37
timestamp 1602073617
transform -1 0 12950 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_39
timestamp 1602073617
transform -1 0 12982 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_38
timestamp 1602073617
transform -1 0 12966 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_40
timestamp 1602073617
transform -1 0 12998 0 -1 1410
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_64
timestamp 1602073617
transform -1 0 658 0 1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_21
timestamp 1602073617
transform -1 0 1308 0 1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_328
timestamp 1602073617
transform 1 0 1308 0 1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_668
timestamp 1602073617
transform 1 0 1958 0 1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_53
timestamp 1602073617
transform 1 0 2608 0 1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_503
timestamp 1602073617
transform 1 0 3258 0 1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_509
timestamp 1602073617
transform 1 0 3908 0 1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_224
timestamp 1602073617
transform 1 0 4558 0 1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_758
timestamp 1602073617
transform 1 0 5208 0 1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_759
timestamp 1602073617
transform -1 0 6508 0 1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_275
timestamp 1602073617
transform -1 0 7158 0 1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_274
timestamp 1602073617
transform -1 0 7808 0 1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_510
timestamp 1602073617
transform -1 0 8458 0 1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_697
timestamp 1602073617
transform 1 0 8458 0 1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_508
timestamp 1602073617
transform -1 0 9758 0 1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_419
timestamp 1602073617
transform 1 0 9758 0 1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_506
timestamp 1602073617
transform -1 0 11058 0 1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_505
timestamp 1602073617
transform 1 0 11058 0 1 1410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_507
timestamp 1602073617
transform -1 0 12358 0 1 1410
box -4 -6 618 206
use FILL  FILL_8_1
timestamp 1602073617
transform 1 0 12358 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_2
timestamp 1602073617
transform 1 0 12374 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_3
timestamp 1602073617
transform 1 0 12390 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_4
timestamp 1602073617
transform 1 0 12406 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_5
timestamp 1602073617
transform 1 0 12422 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_6
timestamp 1602073617
transform 1 0 12438 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_7
timestamp 1602073617
transform 1 0 12454 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_8
timestamp 1602073617
transform 1 0 12470 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_10
timestamp 1602073617
transform 1 0 12502 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_9
timestamp 1602073617
transform 1 0 12486 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_11
timestamp 1602073617
transform 1 0 12518 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_13
timestamp 1602073617
transform 1 0 12550 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_12
timestamp 1602073617
transform 1 0 12534 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_14
timestamp 1602073617
transform 1 0 12566 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_16
timestamp 1602073617
transform 1 0 12598 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_15
timestamp 1602073617
transform 1 0 12582 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_17
timestamp 1602073617
transform 1 0 12614 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_19
timestamp 1602073617
transform 1 0 12646 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_18
timestamp 1602073617
transform 1 0 12630 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_21
timestamp 1602073617
transform 1 0 12678 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_20
timestamp 1602073617
transform 1 0 12662 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_22
timestamp 1602073617
transform 1 0 12694 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_24
timestamp 1602073617
transform 1 0 12726 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_23
timestamp 1602073617
transform 1 0 12710 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_25
timestamp 1602073617
transform 1 0 12742 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_27
timestamp 1602073617
transform 1 0 12774 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_26
timestamp 1602073617
transform 1 0 12758 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_28
timestamp 1602073617
transform 1 0 12790 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_30
timestamp 1602073617
transform 1 0 12822 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_29
timestamp 1602073617
transform 1 0 12806 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_31
timestamp 1602073617
transform 1 0 12838 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_33
timestamp 1602073617
transform 1 0 12870 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_32
timestamp 1602073617
transform 1 0 12854 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_34
timestamp 1602073617
transform 1 0 12886 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_36
timestamp 1602073617
transform 1 0 12918 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_35
timestamp 1602073617
transform 1 0 12902 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_37
timestamp 1602073617
transform 1 0 12934 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_39
timestamp 1602073617
transform 1 0 12966 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_38
timestamp 1602073617
transform 1 0 12950 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_40
timestamp 1602073617
transform 1 0 12982 0 1 1410
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_451
timestamp 1602073617
transform -1 0 658 0 -1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_428
timestamp 1602073617
transform -1 0 1308 0 -1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_596
timestamp 1602073617
transform 1 0 1308 0 -1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_70
timestamp 1602073617
transform -1 0 2608 0 -1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_42
timestamp 1602073617
transform -1 0 3258 0 -1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_502
timestamp 1602073617
transform -1 0 3908 0 -1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_159
timestamp 1602073617
transform -1 0 4558 0 -1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_10
timestamp 1602073617
transform 1 0 4558 0 -1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_296
timestamp 1602073617
transform 1 0 5208 0 -1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_23
timestamp 1602073617
transform 1 0 5858 0 -1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_297
timestamp 1602073617
transform 1 0 6508 0 -1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_347
timestamp 1602073617
transform 1 0 7158 0 -1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_860
timestamp 1602073617
transform 1 0 7808 0 -1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_861
timestamp 1602073617
transform -1 0 9108 0 -1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_360
timestamp 1602073617
transform 1 0 9108 0 -1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_244
timestamp 1602073617
transform -1 0 10408 0 -1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_242
timestamp 1602073617
transform -1 0 11058 0 -1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_239
timestamp 1602073617
transform -1 0 11708 0 -1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_504
timestamp 1602073617
transform 1 0 11708 0 -1 1810
box -4 -6 618 206
use FILL  FILL_9_1
timestamp 1602073617
transform -1 0 12374 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_2
timestamp 1602073617
transform -1 0 12390 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_3
timestamp 1602073617
transform -1 0 12406 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_4
timestamp 1602073617
transform -1 0 12422 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_5
timestamp 1602073617
transform -1 0 12438 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_6
timestamp 1602073617
transform -1 0 12454 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_7
timestamp 1602073617
transform -1 0 12470 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_8
timestamp 1602073617
transform -1 0 12486 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_10
timestamp 1602073617
transform -1 0 12518 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_9
timestamp 1602073617
transform -1 0 12502 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_11
timestamp 1602073617
transform -1 0 12534 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_13
timestamp 1602073617
transform -1 0 12566 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_12
timestamp 1602073617
transform -1 0 12550 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_14
timestamp 1602073617
transform -1 0 12582 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_16
timestamp 1602073617
transform -1 0 12614 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_15
timestamp 1602073617
transform -1 0 12598 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_17
timestamp 1602073617
transform -1 0 12630 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_19
timestamp 1602073617
transform -1 0 12662 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_18
timestamp 1602073617
transform -1 0 12646 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_21
timestamp 1602073617
transform -1 0 12694 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_20
timestamp 1602073617
transform -1 0 12678 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_22
timestamp 1602073617
transform -1 0 12710 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_24
timestamp 1602073617
transform -1 0 12742 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_23
timestamp 1602073617
transform -1 0 12726 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_25
timestamp 1602073617
transform -1 0 12758 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_27
timestamp 1602073617
transform -1 0 12790 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_26
timestamp 1602073617
transform -1 0 12774 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_28
timestamp 1602073617
transform -1 0 12806 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_30
timestamp 1602073617
transform -1 0 12838 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_29
timestamp 1602073617
transform -1 0 12822 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_31
timestamp 1602073617
transform -1 0 12854 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_33
timestamp 1602073617
transform -1 0 12886 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_32
timestamp 1602073617
transform -1 0 12870 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_34
timestamp 1602073617
transform -1 0 12902 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_36
timestamp 1602073617
transform -1 0 12934 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_35
timestamp 1602073617
transform -1 0 12918 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_37
timestamp 1602073617
transform -1 0 12950 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_39
timestamp 1602073617
transform -1 0 12982 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_38
timestamp 1602073617
transform -1 0 12966 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_40
timestamp 1602073617
transform -1 0 12998 0 -1 1810
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_635
timestamp 1602073617
transform -1 0 658 0 1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_582
timestamp 1602073617
transform -1 0 1308 0 1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_161
timestamp 1602073617
transform 1 0 1308 0 1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_387
timestamp 1602073617
transform -1 0 2608 0 1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_92
timestamp 1602073617
transform -1 0 3258 0 1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_56
timestamp 1602073617
transform 1 0 3258 0 1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_669
timestamp 1602073617
transform 1 0 3908 0 1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_720
timestamp 1602073617
transform 1 0 4558 0 1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_304
timestamp 1602073617
transform 1 0 5208 0 1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_721
timestamp 1602073617
transform -1 0 6508 0 1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_845
timestamp 1602073617
transform 1 0 6508 0 1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_268
timestamp 1602073617
transform 1 0 7158 0 1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_865
timestamp 1602073617
transform -1 0 8458 0 1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_658
timestamp 1602073617
transform -1 0 9108 0 1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_849
timestamp 1602073617
transform 1 0 9108 0 1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_862
timestamp 1602073617
transform 1 0 9758 0 1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_447
timestamp 1602073617
transform -1 0 11058 0 1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_258
timestamp 1602073617
transform 1 0 11058 0 1 1810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_420
timestamp 1602073617
transform 1 0 11708 0 1 1810
box -4 -6 618 206
use FILL  FILL_10_1
timestamp 1602073617
transform 1 0 12358 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_2
timestamp 1602073617
transform 1 0 12374 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_3
timestamp 1602073617
transform 1 0 12390 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_4
timestamp 1602073617
transform 1 0 12406 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_5
timestamp 1602073617
transform 1 0 12422 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_6
timestamp 1602073617
transform 1 0 12438 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_7
timestamp 1602073617
transform 1 0 12454 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_8
timestamp 1602073617
transform 1 0 12470 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_10
timestamp 1602073617
transform 1 0 12502 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_9
timestamp 1602073617
transform 1 0 12486 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_11
timestamp 1602073617
transform 1 0 12518 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_13
timestamp 1602073617
transform 1 0 12550 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_12
timestamp 1602073617
transform 1 0 12534 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_14
timestamp 1602073617
transform 1 0 12566 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_16
timestamp 1602073617
transform 1 0 12598 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_15
timestamp 1602073617
transform 1 0 12582 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_17
timestamp 1602073617
transform 1 0 12614 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_19
timestamp 1602073617
transform 1 0 12646 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_18
timestamp 1602073617
transform 1 0 12630 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_21
timestamp 1602073617
transform 1 0 12678 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_20
timestamp 1602073617
transform 1 0 12662 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_22
timestamp 1602073617
transform 1 0 12694 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_24
timestamp 1602073617
transform 1 0 12726 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_23
timestamp 1602073617
transform 1 0 12710 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_25
timestamp 1602073617
transform 1 0 12742 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_27
timestamp 1602073617
transform 1 0 12774 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_26
timestamp 1602073617
transform 1 0 12758 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_28
timestamp 1602073617
transform 1 0 12790 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_30
timestamp 1602073617
transform 1 0 12822 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_29
timestamp 1602073617
transform 1 0 12806 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_31
timestamp 1602073617
transform 1 0 12838 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_33
timestamp 1602073617
transform 1 0 12870 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_32
timestamp 1602073617
transform 1 0 12854 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_34
timestamp 1602073617
transform 1 0 12886 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_36
timestamp 1602073617
transform 1 0 12918 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_35
timestamp 1602073617
transform 1 0 12902 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_37
timestamp 1602073617
transform 1 0 12934 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_39
timestamp 1602073617
transform 1 0 12966 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_38
timestamp 1602073617
transform 1 0 12950 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_40
timestamp 1602073617
transform 1 0 12982 0 1 1810
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_452
timestamp 1602073617
transform -1 0 658 0 -1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_450
timestamp 1602073617
transform -1 0 1308 0 -1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_427
timestamp 1602073617
transform -1 0 1958 0 -1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_426
timestamp 1602073617
transform -1 0 2608 0 -1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_617
timestamp 1602073617
transform 1 0 2608 0 -1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_77
timestamp 1602073617
transform -1 0 3908 0 -1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_38
timestamp 1602073617
transform -1 0 4558 0 -1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_667
timestamp 1602073617
transform -1 0 5208 0 -1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_236
timestamp 1602073617
transform 1 0 5208 0 -1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_276
timestamp 1602073617
transform -1 0 6508 0 -1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_271
timestamp 1602073617
transform -1 0 7158 0 -1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_269
timestamp 1602073617
transform -1 0 7808 0 -1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_256
timestamp 1602073617
transform 1 0 7808 0 -1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_270
timestamp 1602073617
transform 1 0 8458 0 -1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_247
timestamp 1602073617
transform 1 0 9108 0 -1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_125
timestamp 1602073617
transform 1 0 9758 0 -1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_257
timestamp 1602073617
transform 1 0 10408 0 -1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_259
timestamp 1602073617
transform 1 0 11058 0 -1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_345
timestamp 1602073617
transform 1 0 11708 0 -1 2210
box -4 -6 618 206
use FILL  FILL_11_1
timestamp 1602073617
transform -1 0 12374 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_2
timestamp 1602073617
transform -1 0 12390 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_3
timestamp 1602073617
transform -1 0 12406 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_4
timestamp 1602073617
transform -1 0 12422 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_5
timestamp 1602073617
transform -1 0 12438 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_6
timestamp 1602073617
transform -1 0 12454 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_7
timestamp 1602073617
transform -1 0 12470 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_8
timestamp 1602073617
transform -1 0 12486 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_10
timestamp 1602073617
transform -1 0 12518 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_9
timestamp 1602073617
transform -1 0 12502 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_11
timestamp 1602073617
transform -1 0 12534 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_13
timestamp 1602073617
transform -1 0 12566 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_12
timestamp 1602073617
transform -1 0 12550 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_14
timestamp 1602073617
transform -1 0 12582 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_16
timestamp 1602073617
transform -1 0 12614 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_15
timestamp 1602073617
transform -1 0 12598 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_17
timestamp 1602073617
transform -1 0 12630 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_19
timestamp 1602073617
transform -1 0 12662 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_18
timestamp 1602073617
transform -1 0 12646 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_21
timestamp 1602073617
transform -1 0 12694 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_20
timestamp 1602073617
transform -1 0 12678 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_22
timestamp 1602073617
transform -1 0 12710 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_24
timestamp 1602073617
transform -1 0 12742 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_23
timestamp 1602073617
transform -1 0 12726 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_25
timestamp 1602073617
transform -1 0 12758 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_27
timestamp 1602073617
transform -1 0 12790 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_26
timestamp 1602073617
transform -1 0 12774 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_28
timestamp 1602073617
transform -1 0 12806 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_30
timestamp 1602073617
transform -1 0 12838 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_29
timestamp 1602073617
transform -1 0 12822 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_31
timestamp 1602073617
transform -1 0 12854 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_33
timestamp 1602073617
transform -1 0 12886 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_32
timestamp 1602073617
transform -1 0 12870 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_34
timestamp 1602073617
transform -1 0 12902 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_36
timestamp 1602073617
transform -1 0 12934 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_35
timestamp 1602073617
transform -1 0 12918 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_37
timestamp 1602073617
transform -1 0 12950 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_39
timestamp 1602073617
transform -1 0 12982 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_38
timestamp 1602073617
transform -1 0 12966 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_40
timestamp 1602073617
transform -1 0 12998 0 -1 2210
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_639
timestamp 1602073617
transform 1 0 8 0 1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_636
timestamp 1602073617
transform -1 0 1308 0 1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_583
timestamp 1602073617
transform -1 0 1958 0 1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_162
timestamp 1602073617
transform -1 0 2608 0 1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_160
timestamp 1602073617
transform -1 0 3258 0 1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_126
timestamp 1602073617
transform -1 0 3908 0 1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_54
timestamp 1602073617
transform -1 0 4558 0 1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_129
timestamp 1602073617
transform -1 0 5208 0 1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_294
timestamp 1602073617
transform 1 0 5208 0 1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_307
timestamp 1602073617
transform 1 0 5858 0 1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_130
timestamp 1602073617
transform 1 0 6508 0 1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_131
timestamp 1602073617
transform 1 0 7158 0 1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_383
timestamp 1602073617
transform 1 0 7808 0 1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_481
timestamp 1602073617
transform 1 0 8458 0 1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_127
timestamp 1602073617
transform 1 0 9108 0 1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_128
timestamp 1602073617
transform -1 0 10408 0 1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_363
timestamp 1602073617
transform -1 0 11058 0 1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_359
timestamp 1602073617
transform -1 0 11708 0 1 2210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_555
timestamp 1602073617
transform 1 0 11708 0 1 2210
box -4 -6 618 206
use FILL  FILL_12_1
timestamp 1602073617
transform 1 0 12358 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_2
timestamp 1602073617
transform 1 0 12374 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_3
timestamp 1602073617
transform 1 0 12390 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_4
timestamp 1602073617
transform 1 0 12406 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_5
timestamp 1602073617
transform 1 0 12422 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_6
timestamp 1602073617
transform 1 0 12438 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_7
timestamp 1602073617
transform 1 0 12454 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_8
timestamp 1602073617
transform 1 0 12470 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_10
timestamp 1602073617
transform 1 0 12502 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_9
timestamp 1602073617
transform 1 0 12486 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_11
timestamp 1602073617
transform 1 0 12518 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_13
timestamp 1602073617
transform 1 0 12550 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_12
timestamp 1602073617
transform 1 0 12534 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_14
timestamp 1602073617
transform 1 0 12566 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_16
timestamp 1602073617
transform 1 0 12598 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_15
timestamp 1602073617
transform 1 0 12582 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_17
timestamp 1602073617
transform 1 0 12614 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_19
timestamp 1602073617
transform 1 0 12646 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_18
timestamp 1602073617
transform 1 0 12630 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_21
timestamp 1602073617
transform 1 0 12678 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_20
timestamp 1602073617
transform 1 0 12662 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_22
timestamp 1602073617
transform 1 0 12694 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_24
timestamp 1602073617
transform 1 0 12726 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_23
timestamp 1602073617
transform 1 0 12710 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_25
timestamp 1602073617
transform 1 0 12742 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_27
timestamp 1602073617
transform 1 0 12774 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_26
timestamp 1602073617
transform 1 0 12758 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_28
timestamp 1602073617
transform 1 0 12790 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_30
timestamp 1602073617
transform 1 0 12822 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_29
timestamp 1602073617
transform 1 0 12806 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_31
timestamp 1602073617
transform 1 0 12838 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_33
timestamp 1602073617
transform 1 0 12870 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_32
timestamp 1602073617
transform 1 0 12854 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_34
timestamp 1602073617
transform 1 0 12886 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_36
timestamp 1602073617
transform 1 0 12918 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_35
timestamp 1602073617
transform 1 0 12902 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_37
timestamp 1602073617
transform 1 0 12934 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_39
timestamp 1602073617
transform 1 0 12966 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_38
timestamp 1602073617
transform 1 0 12950 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_40
timestamp 1602073617
transform 1 0 12982 0 1 2210
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_651
timestamp 1602073617
transform 1 0 8 0 -1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_588
timestamp 1602073617
transform -1 0 1308 0 -1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_586
timestamp 1602073617
transform -1 0 1958 0 -1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_584
timestamp 1602073617
transform -1 0 2608 0 -1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_120
timestamp 1602073617
transform 1 0 2608 0 -1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_415
timestamp 1602073617
transform -1 0 3908 0 -1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_55
timestamp 1602073617
transform -1 0 4558 0 -1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_29
timestamp 1602073617
transform -1 0 5208 0 -1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_293
timestamp 1602073617
transform -1 0 5858 0 -1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_49
timestamp 1602073617
transform -1 0 6508 0 -1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_85
timestamp 1602073617
transform 1 0 6508 0 -1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_305
timestamp 1602073617
transform -1 0 7808 0 -1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_136
timestamp 1602073617
transform 1 0 7808 0 -1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_138
timestamp 1602073617
transform 1 0 8458 0 -1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_132
timestamp 1602073617
transform 1 0 9108 0 -1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_140
timestamp 1602073617
transform 1 0 9758 0 -1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_135
timestamp 1602073617
transform -1 0 11058 0 -1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_253
timestamp 1602073617
transform 1 0 11058 0 -1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_248
timestamp 1602073617
transform -1 0 12358 0 -1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_344
timestamp 1602073617
transform 1 0 12358 0 -1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_638
timestamp 1602073617
transform -1 0 658 0 1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_637
timestamp 1602073617
transform -1 0 1308 0 1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_585
timestamp 1602073617
transform -1 0 1958 0 1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_375
timestamp 1602073617
transform -1 0 2608 0 1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_119
timestamp 1602073617
transform -1 0 3258 0 1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_121
timestamp 1602073617
transform 1 0 3258 0 1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_87
timestamp 1602073617
transform -1 0 4558 0 1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_32
timestamp 1602073617
transform 1 0 4558 0 1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_813
timestamp 1602073617
transform 1 0 5208 0 1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_659
timestamp 1602073617
transform -1 0 6508 0 1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_657
timestamp 1602073617
transform -1 0 7158 0 1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_574
timestamp 1602073617
transform -1 0 7808 0 1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_141
timestamp 1602073617
transform -1 0 8458 0 1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_139
timestamp 1602073617
transform -1 0 9108 0 1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_137
timestamp 1602073617
transform -1 0 9758 0 1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_105
timestamp 1602073617
transform 1 0 9758 0 1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_252
timestamp 1602073617
transform 1 0 10408 0 1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_632
timestamp 1602073617
transform -1 0 11708 0 1 2610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_254
timestamp 1602073617
transform 1 0 11708 0 1 2610
box -4 -6 618 206
use FILL  FILL_14_1
timestamp 1602073617
transform 1 0 12358 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_2
timestamp 1602073617
transform 1 0 12374 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_3
timestamp 1602073617
transform 1 0 12390 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_4
timestamp 1602073617
transform 1 0 12406 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_5
timestamp 1602073617
transform 1 0 12422 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_6
timestamp 1602073617
transform 1 0 12438 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_7
timestamp 1602073617
transform 1 0 12454 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_8
timestamp 1602073617
transform 1 0 12470 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_10
timestamp 1602073617
transform 1 0 12502 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_9
timestamp 1602073617
transform 1 0 12486 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_11
timestamp 1602073617
transform 1 0 12518 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_13
timestamp 1602073617
transform 1 0 12550 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_12
timestamp 1602073617
transform 1 0 12534 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_14
timestamp 1602073617
transform 1 0 12566 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_16
timestamp 1602073617
transform 1 0 12598 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_15
timestamp 1602073617
transform 1 0 12582 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_17
timestamp 1602073617
transform 1 0 12614 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_19
timestamp 1602073617
transform 1 0 12646 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_18
timestamp 1602073617
transform 1 0 12630 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_21
timestamp 1602073617
transform 1 0 12678 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_20
timestamp 1602073617
transform 1 0 12662 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_22
timestamp 1602073617
transform 1 0 12694 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_24
timestamp 1602073617
transform 1 0 12726 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_23
timestamp 1602073617
transform 1 0 12710 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_25
timestamp 1602073617
transform 1 0 12742 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_27
timestamp 1602073617
transform 1 0 12774 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_26
timestamp 1602073617
transform 1 0 12758 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_28
timestamp 1602073617
transform 1 0 12790 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_30
timestamp 1602073617
transform 1 0 12822 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_29
timestamp 1602073617
transform 1 0 12806 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_31
timestamp 1602073617
transform 1 0 12838 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_33
timestamp 1602073617
transform 1 0 12870 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_32
timestamp 1602073617
transform 1 0 12854 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_34
timestamp 1602073617
transform 1 0 12886 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_36
timestamp 1602073617
transform 1 0 12918 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_35
timestamp 1602073617
transform 1 0 12902 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_37
timestamp 1602073617
transform 1 0 12934 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_39
timestamp 1602073617
transform 1 0 12966 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_38
timestamp 1602073617
transform 1 0 12950 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_40
timestamp 1602073617
transform 1 0 12982 0 1 2610
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_467
timestamp 1602073617
transform -1 0 658 0 -1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_163
timestamp 1602073617
transform -1 0 1308 0 -1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_376
timestamp 1602073617
transform -1 0 1958 0 -1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_411
timestamp 1602073617
transform 1 0 1958 0 -1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_461
timestamp 1602073617
transform 1 0 2608 0 -1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_19
timestamp 1602073617
transform -1 0 3908 0 -1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_102
timestamp 1602073617
transform -1 0 4558 0 -1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_263
timestamp 1602073617
transform 1 0 4558 0 -1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_66
timestamp 1602073617
transform 1 0 5208 0 -1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_625
timestamp 1602073617
transform 1 0 5858 0 -1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_62
timestamp 1602073617
transform -1 0 7158 0 -1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_490
timestamp 1602073617
transform 1 0 7158 0 -1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_514
timestamp 1602073617
transform -1 0 8458 0 -1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_73
timestamp 1602073617
transform 1 0 8458 0 -1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_246
timestamp 1602073617
transform 1 0 9108 0 -1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_342
timestamp 1602073617
transform 1 0 9758 0 -1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_349
timestamp 1602073617
transform 1 0 10408 0 -1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_134
timestamp 1602073617
transform 1 0 11058 0 -1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_631
timestamp 1602073617
transform 1 0 11708 0 -1 3010
box -4 -6 618 206
use FILL  FILL_15_1
timestamp 1602073617
transform -1 0 12374 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_2
timestamp 1602073617
transform -1 0 12390 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_3
timestamp 1602073617
transform -1 0 12406 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_4
timestamp 1602073617
transform -1 0 12422 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_5
timestamp 1602073617
transform -1 0 12438 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_6
timestamp 1602073617
transform -1 0 12454 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_7
timestamp 1602073617
transform -1 0 12470 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_8
timestamp 1602073617
transform -1 0 12486 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_10
timestamp 1602073617
transform -1 0 12518 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_9
timestamp 1602073617
transform -1 0 12502 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_11
timestamp 1602073617
transform -1 0 12534 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_13
timestamp 1602073617
transform -1 0 12566 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_12
timestamp 1602073617
transform -1 0 12550 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_14
timestamp 1602073617
transform -1 0 12582 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_16
timestamp 1602073617
transform -1 0 12614 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_15
timestamp 1602073617
transform -1 0 12598 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_17
timestamp 1602073617
transform -1 0 12630 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_19
timestamp 1602073617
transform -1 0 12662 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_18
timestamp 1602073617
transform -1 0 12646 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_21
timestamp 1602073617
transform -1 0 12694 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_20
timestamp 1602073617
transform -1 0 12678 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_22
timestamp 1602073617
transform -1 0 12710 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_24
timestamp 1602073617
transform -1 0 12742 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_23
timestamp 1602073617
transform -1 0 12726 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_25
timestamp 1602073617
transform -1 0 12758 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_27
timestamp 1602073617
transform -1 0 12790 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_26
timestamp 1602073617
transform -1 0 12774 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_28
timestamp 1602073617
transform -1 0 12806 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_30
timestamp 1602073617
transform -1 0 12838 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_29
timestamp 1602073617
transform -1 0 12822 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_31
timestamp 1602073617
transform -1 0 12854 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_33
timestamp 1602073617
transform -1 0 12886 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_32
timestamp 1602073617
transform -1 0 12870 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_34
timestamp 1602073617
transform -1 0 12902 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_36
timestamp 1602073617
transform -1 0 12934 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_35
timestamp 1602073617
transform -1 0 12918 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_37
timestamp 1602073617
transform -1 0 12950 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_39
timestamp 1602073617
transform -1 0 12982 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_38
timestamp 1602073617
transform -1 0 12966 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_40
timestamp 1602073617
transform -1 0 12998 0 -1 3010
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_422
timestamp 1602073617
transform -1 0 658 0 1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_410
timestamp 1602073617
transform 1 0 658 0 1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_459
timestamp 1602073617
transform 1 0 1308 0 1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_378
timestamp 1602073617
transform -1 0 2608 0 1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_377
timestamp 1602073617
transform -1 0 3258 0 1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_90
timestamp 1602073617
transform -1 0 3908 0 1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_340
timestamp 1602073617
transform -1 0 4558 0 1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_88
timestamp 1602073617
transform -1 0 5208 0 1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_34
timestamp 1602073617
transform -1 0 5858 0 1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_27
timestamp 1602073617
transform -1 0 6508 0 1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_235
timestamp 1602073617
transform 1 0 6508 0 1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_243
timestamp 1602073617
transform 1 0 7158 0 1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_245
timestamp 1602073617
transform 1 0 7808 0 1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_777
timestamp 1602073617
transform 1 0 8458 0 1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_784
timestamp 1602073617
transform 1 0 9108 0 1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_858
timestamp 1602073617
transform -1 0 10408 0 1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_482
timestamp 1602073617
transform 1 0 10408 0 1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_483
timestamp 1602073617
transform 1 0 11058 0 1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_556
timestamp 1602073617
transform 1 0 11708 0 1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_562
timestamp 1602073617
transform 1 0 12358 0 1 3010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_466
timestamp 1602073617
transform -1 0 658 0 -1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_453
timestamp 1602073617
transform -1 0 1308 0 -1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_448
timestamp 1602073617
transform -1 0 1958 0 -1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_421
timestamp 1602073617
transform -1 0 2608 0 -1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_826
timestamp 1602073617
transform 1 0 2608 0 -1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_837
timestamp 1602073617
transform 1 0 3258 0 -1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_94
timestamp 1602073617
transform -1 0 4558 0 -1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_100
timestamp 1602073617
transform 1 0 4558 0 -1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_86
timestamp 1602073617
transform -1 0 5858 0 -1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_454
timestamp 1602073617
transform -1 0 6508 0 -1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_446
timestamp 1602073617
transform -1 0 7158 0 -1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_417
timestamp 1602073617
transform 1 0 7158 0 -1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_515
timestamp 1602073617
transform 1 0 7808 0 -1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_516
timestamp 1602073617
transform -1 0 9108 0 -1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_513
timestamp 1602073617
transform -1 0 9758 0 -1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_834
timestamp 1602073617
transform 1 0 9758 0 -1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_840
timestamp 1602073617
transform -1 0 11058 0 -1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_833
timestamp 1602073617
transform -1 0 11708 0 -1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_626
timestamp 1602073617
transform 1 0 11708 0 -1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_629
timestamp 1602073617
transform 1 0 12358 0 -1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_470
timestamp 1602073617
transform 1 0 8 0 1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_769
timestamp 1602073617
transform -1 0 658 0 -1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_763
timestamp 1602073617
transform -1 0 1308 0 1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_409
timestamp 1602073617
transform 1 0 658 0 -1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_764
timestamp 1602073617
transform -1 0 1958 0 1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_460
timestamp 1602073617
transform 1 0 1308 0 -1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_413
timestamp 1602073617
transform 1 0 1958 0 1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_463
timestamp 1602073617
transform 1 0 1958 0 -1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_416
timestamp 1602073617
transform -1 0 3258 0 1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_380
timestamp 1602073617
transform -1 0 3258 0 -1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_825
timestamp 1602073617
transform -1 0 3908 0 1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_153
timestamp 1602073617
transform 1 0 3258 0 -1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_96
timestamp 1602073617
transform 1 0 3908 0 1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_122
timestamp 1602073617
transform 1 0 3908 0 -1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_63
timestamp 1602073617
transform 1 0 4558 0 1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_98
timestamp 1602073617
transform 1 0 4558 0 -1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_82
timestamp 1602073617
transform 1 0 5208 0 1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_93
timestamp 1602073617
transform -1 0 5858 0 -1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_371
timestamp 1602073617
transform 1 0 5858 0 1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_46
timestamp 1602073617
transform 1 0 5858 0 -1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_778
timestamp 1602073617
transform 1 0 6508 0 1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_418
timestamp 1602073617
transform 1 0 6508 0 -1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_273
timestamp 1602073617
transform 1 0 7158 0 1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_9
timestamp 1602073617
transform 1 0 7158 0 -1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_831
timestamp 1602073617
transform 1 0 7808 0 1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_372
timestamp 1602073617
transform 1 0 7808 0 -1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_841
timestamp 1602073617
transform 1 0 8458 0 1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_844
timestamp 1602073617
transform 1 0 8458 0 -1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_511
timestamp 1602073617
transform 1 0 9108 0 1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_496
timestamp 1602073617
transform -1 0 9758 0 -1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_851
timestamp 1602073617
transform -1 0 10408 0 1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_779
timestamp 1602073617
transform 1 0 9758 0 -1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_107
timestamp 1602073617
transform 1 0 10408 0 1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_783
timestamp 1602073617
transform 1 0 10408 0 -1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_627
timestamp 1602073617
transform 1 0 11058 0 1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_796
timestamp 1602073617
transform 1 0 11058 0 -1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_630
timestamp 1602073617
transform -1 0 12358 0 1 3410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_113
timestamp 1602073617
transform -1 0 12358 0 -1 3810
box -4 -6 618 206
use FILL  FILL_18_1
timestamp 1602073617
transform 1 0 12358 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_2
timestamp 1602073617
transform 1 0 12374 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_3
timestamp 1602073617
transform 1 0 12390 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_4
timestamp 1602073617
transform 1 0 12406 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_5
timestamp 1602073617
transform 1 0 12422 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_6
timestamp 1602073617
transform 1 0 12438 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_7
timestamp 1602073617
transform 1 0 12454 0 1 3410
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_628
timestamp 1602073617
transform -1 0 13008 0 -1 3810
box -4 -6 618 206
use FILL  FILL_18_8
timestamp 1602073617
transform 1 0 12470 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_10
timestamp 1602073617
transform 1 0 12502 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_9
timestamp 1602073617
transform 1 0 12486 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_11
timestamp 1602073617
transform 1 0 12518 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_13
timestamp 1602073617
transform 1 0 12550 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_12
timestamp 1602073617
transform 1 0 12534 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_14
timestamp 1602073617
transform 1 0 12566 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_16
timestamp 1602073617
transform 1 0 12598 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_15
timestamp 1602073617
transform 1 0 12582 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_17
timestamp 1602073617
transform 1 0 12614 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_19
timestamp 1602073617
transform 1 0 12646 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_18
timestamp 1602073617
transform 1 0 12630 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_21
timestamp 1602073617
transform 1 0 12678 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_20
timestamp 1602073617
transform 1 0 12662 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_22
timestamp 1602073617
transform 1 0 12694 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_24
timestamp 1602073617
transform 1 0 12726 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_23
timestamp 1602073617
transform 1 0 12710 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_25
timestamp 1602073617
transform 1 0 12742 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_27
timestamp 1602073617
transform 1 0 12774 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_26
timestamp 1602073617
transform 1 0 12758 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_28
timestamp 1602073617
transform 1 0 12790 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_30
timestamp 1602073617
transform 1 0 12822 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_29
timestamp 1602073617
transform 1 0 12806 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_31
timestamp 1602073617
transform 1 0 12838 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_33
timestamp 1602073617
transform 1 0 12870 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_32
timestamp 1602073617
transform 1 0 12854 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_34
timestamp 1602073617
transform 1 0 12886 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_36
timestamp 1602073617
transform 1 0 12918 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_35
timestamp 1602073617
transform 1 0 12902 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_37
timestamp 1602073617
transform 1 0 12934 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_39
timestamp 1602073617
transform 1 0 12966 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_38
timestamp 1602073617
transform 1 0 12950 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_40
timestamp 1602073617
transform 1 0 12982 0 1 3410
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_771
timestamp 1602073617
transform 1 0 8 0 1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_766
timestamp 1602073617
transform 1 0 658 0 1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_407
timestamp 1602073617
transform -1 0 1958 0 1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_379
timestamp 1602073617
transform 1 0 1958 0 1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_520
timestamp 1602073617
transform -1 0 3258 0 1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_518
timestamp 1602073617
transform -1 0 3908 0 1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_233
timestamp 1602073617
transform 1 0 3908 0 1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_517
timestamp 1602073617
transform 1 0 4558 0 1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_559
timestamp 1602073617
transform 1 0 5208 0 1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_15
timestamp 1602073617
transform -1 0 6508 0 1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_71
timestamp 1602073617
transform 1 0 6508 0 1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_300
timestamp 1602073617
transform 1 0 7158 0 1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_500
timestamp 1602073617
transform -1 0 8458 0 1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_497
timestamp 1602073617
transform -1 0 9108 0 1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_499
timestamp 1602073617
transform -1 0 9758 0 1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_495
timestamp 1602073617
transform -1 0 10408 0 1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_850
timestamp 1602073617
transform -1 0 11058 0 1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_768
timestamp 1602073617
transform -1 0 11708 0 1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_103
timestamp 1602073617
transform 1 0 11708 0 1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_570
timestamp 1602073617
transform -1 0 13008 0 1 3810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_477
timestamp 1602073617
transform -1 0 658 0 -1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_770
timestamp 1602073617
transform -1 0 1308 0 -1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_765
timestamp 1602073617
transform -1 0 1958 0 -1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_642
timestamp 1602073617
transform -1 0 2608 0 -1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_677
timestamp 1602073617
transform 1 0 2608 0 -1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_462
timestamp 1602073617
transform 1 0 3258 0 -1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_472
timestamp 1602073617
transform 1 0 3908 0 -1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_155
timestamp 1602073617
transform -1 0 5208 0 -1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_124
timestamp 1602073617
transform 1 0 5208 0 -1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_519
timestamp 1602073617
transform -1 0 6508 0 -1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_150
timestamp 1602073617
transform 1 0 6508 0 -1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_232
timestamp 1602073617
transform 1 0 7158 0 -1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_240
timestamp 1602073617
transform 1 0 7808 0 -1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_494
timestamp 1602073617
transform 1 0 8458 0 -1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_458
timestamp 1602073617
transform 1 0 9108 0 -1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_368
timestamp 1602073617
transform 1 0 9758 0 -1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_251
timestamp 1602073617
transform -1 0 11058 0 -1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_184
timestamp 1602073617
transform 1 0 11058 0 -1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_842
timestamp 1602073617
transform -1 0 12358 0 -1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_553
timestamp 1602073617
transform -1 0 13008 0 -1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_774
timestamp 1602073617
transform -1 0 658 0 1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_678
timestamp 1602073617
transform -1 0 1308 0 1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_649
timestamp 1602073617
transform -1 0 1958 0 1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_424
timestamp 1602073617
transform -1 0 2608 0 1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_412
timestamp 1602073617
transform -1 0 3258 0 1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_210
timestamp 1602073617
transform 1 0 3258 0 1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_158
timestamp 1602073617
transform -1 0 4558 0 1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_117
timestamp 1602073617
transform -1 0 5208 0 1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_67
timestamp 1602073617
transform -1 0 5858 0 1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_217
timestamp 1602073617
transform -1 0 6508 0 1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_234
timestamp 1602073617
transform 1 0 6508 0 1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_277
timestamp 1602073617
transform 1 0 7158 0 1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_278
timestamp 1602073617
transform 1 0 7808 0 1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_471
timestamp 1602073617
transform -1 0 9108 0 1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_464
timestamp 1602073617
transform -1 0 9758 0 1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_457
timestamp 1602073617
transform -1 0 10408 0 1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_843
timestamp 1602073617
transform 1 0 10408 0 1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_106
timestamp 1602073617
transform 1 0 11058 0 1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_554
timestamp 1602073617
transform 1 0 11708 0 1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_563
timestamp 1602073617
transform 1 0 12358 0 1 4210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_866
timestamp 1602073617
transform -1 0 658 0 -1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_864
timestamp 1602073617
transform -1 0 1308 0 -1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_449
timestamp 1602073617
transform -1 0 1958 0 -1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_690
timestamp 1602073617
transform -1 0 2608 0 -1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_832
timestamp 1602073617
transform 1 0 2608 0 -1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_154
timestamp 1602073617
transform 1 0 3258 0 -1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_156
timestamp 1602073617
transform 1 0 3908 0 -1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_123
timestamp 1602073617
transform 1 0 4558 0 -1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_202
timestamp 1602073617
transform 1 0 5208 0 -1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_773
timestamp 1602073617
transform -1 0 6508 0 -1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_572
timestamp 1602073617
transform 1 0 6508 0 -1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_69
timestamp 1602073617
transform -1 0 7808 0 -1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_560
timestamp 1602073617
transform -1 0 8458 0 -1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_488
timestamp 1602073617
transform 1 0 8458 0 -1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_523
timestamp 1602073617
transform -1 0 9758 0 -1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_521
timestamp 1602073617
transform -1 0 10408 0 -1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_343
timestamp 1602073617
transform 1 0 10408 0 -1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_115
timestamp 1602073617
transform -1 0 11708 0 -1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_456
timestamp 1602073617
transform -1 0 12358 0 -1 4610
box -4 -6 618 206
use FILL  FILL_23_1
timestamp 1602073617
transform -1 0 12374 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_2
timestamp 1602073617
transform -1 0 12390 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_3
timestamp 1602073617
transform -1 0 12406 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_4
timestamp 1602073617
transform -1 0 12422 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_5
timestamp 1602073617
transform -1 0 12438 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_6
timestamp 1602073617
transform -1 0 12454 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_7
timestamp 1602073617
transform -1 0 12470 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_8
timestamp 1602073617
transform -1 0 12486 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_10
timestamp 1602073617
transform -1 0 12518 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_9
timestamp 1602073617
transform -1 0 12502 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_11
timestamp 1602073617
transform -1 0 12534 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_13
timestamp 1602073617
transform -1 0 12566 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_12
timestamp 1602073617
transform -1 0 12550 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_14
timestamp 1602073617
transform -1 0 12582 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_16
timestamp 1602073617
transform -1 0 12614 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_15
timestamp 1602073617
transform -1 0 12598 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_17
timestamp 1602073617
transform -1 0 12630 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_19
timestamp 1602073617
transform -1 0 12662 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_18
timestamp 1602073617
transform -1 0 12646 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_21
timestamp 1602073617
transform -1 0 12694 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_20
timestamp 1602073617
transform -1 0 12678 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_22
timestamp 1602073617
transform -1 0 12710 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_24
timestamp 1602073617
transform -1 0 12742 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_23
timestamp 1602073617
transform -1 0 12726 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_25
timestamp 1602073617
transform -1 0 12758 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_27
timestamp 1602073617
transform -1 0 12790 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_26
timestamp 1602073617
transform -1 0 12774 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_28
timestamp 1602073617
transform -1 0 12806 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_30
timestamp 1602073617
transform -1 0 12838 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_29
timestamp 1602073617
transform -1 0 12822 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_31
timestamp 1602073617
transform -1 0 12854 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_33
timestamp 1602073617
transform -1 0 12886 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_32
timestamp 1602073617
transform -1 0 12870 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_34
timestamp 1602073617
transform -1 0 12902 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_36
timestamp 1602073617
transform -1 0 12934 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_35
timestamp 1602073617
transform -1 0 12918 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_37
timestamp 1602073617
transform -1 0 12950 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_39
timestamp 1602073617
transform -1 0 12982 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_38
timestamp 1602073617
transform -1 0 12966 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_40
timestamp 1602073617
transform -1 0 12998 0 -1 4610
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_828
timestamp 1602073617
transform -1 0 658 0 1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_592
timestamp 1602073617
transform -1 0 1308 0 1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_423
timestamp 1602073617
transform -1 0 1958 0 1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_230
timestamp 1602073617
transform 1 0 1958 0 1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_249
timestamp 1602073617
transform -1 0 3258 0 1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_78
timestamp 1602073617
transform 1 0 3258 0 1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_476
timestamp 1602073617
transform -1 0 4558 0 1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_264
timestamp 1602073617
transform 1 0 4558 0 1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_473
timestamp 1602073617
transform -1 0 5858 0 1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_767
timestamp 1602073617
transform 1 0 5858 0 1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_576
timestamp 1602073617
transform -1 0 7158 0 1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_571
timestamp 1602073617
transform -1 0 7808 0 1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_287
timestamp 1602073617
transform -1 0 8458 0 1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_522
timestamp 1602073617
transform 1 0 8458 0 1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_250
timestamp 1602073617
transform 1 0 9108 0 1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_116
timestamp 1602073617
transform -1 0 10408 0 1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_114
timestamp 1602073617
transform -1 0 11058 0 1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_183
timestamp 1602073617
transform 1 0 11058 0 1 4610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_190
timestamp 1602073617
transform -1 0 12358 0 1 4610
box -4 -6 618 206
use FILL  FILL_24_1
timestamp 1602073617
transform 1 0 12358 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_2
timestamp 1602073617
transform 1 0 12374 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_3
timestamp 1602073617
transform 1 0 12390 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_4
timestamp 1602073617
transform 1 0 12406 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_5
timestamp 1602073617
transform 1 0 12422 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_6
timestamp 1602073617
transform 1 0 12438 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_7
timestamp 1602073617
transform 1 0 12454 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_8
timestamp 1602073617
transform 1 0 12470 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_10
timestamp 1602073617
transform 1 0 12502 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_9
timestamp 1602073617
transform 1 0 12486 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_11
timestamp 1602073617
transform 1 0 12518 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_13
timestamp 1602073617
transform 1 0 12550 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_12
timestamp 1602073617
transform 1 0 12534 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_14
timestamp 1602073617
transform 1 0 12566 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_16
timestamp 1602073617
transform 1 0 12598 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_15
timestamp 1602073617
transform 1 0 12582 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_17
timestamp 1602073617
transform 1 0 12614 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_19
timestamp 1602073617
transform 1 0 12646 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_18
timestamp 1602073617
transform 1 0 12630 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_21
timestamp 1602073617
transform 1 0 12678 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_20
timestamp 1602073617
transform 1 0 12662 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_22
timestamp 1602073617
transform 1 0 12694 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_24
timestamp 1602073617
transform 1 0 12726 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_23
timestamp 1602073617
transform 1 0 12710 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_25
timestamp 1602073617
transform 1 0 12742 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_27
timestamp 1602073617
transform 1 0 12774 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_26
timestamp 1602073617
transform 1 0 12758 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_28
timestamp 1602073617
transform 1 0 12790 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_30
timestamp 1602073617
transform 1 0 12822 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_29
timestamp 1602073617
transform 1 0 12806 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_31
timestamp 1602073617
transform 1 0 12838 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_33
timestamp 1602073617
transform 1 0 12870 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_32
timestamp 1602073617
transform 1 0 12854 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_34
timestamp 1602073617
transform 1 0 12886 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_36
timestamp 1602073617
transform 1 0 12918 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_35
timestamp 1602073617
transform 1 0 12902 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_37
timestamp 1602073617
transform 1 0 12934 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_39
timestamp 1602073617
transform 1 0 12966 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_38
timestamp 1602073617
transform 1 0 12950 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_40
timestamp 1602073617
transform 1 0 12982 0 1 4610
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_654
timestamp 1602073617
transform -1 0 658 0 -1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_650
timestamp 1602073617
transform -1 0 1308 0 -1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_640
timestamp 1602073617
transform -1 0 1958 0 -1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_633
timestamp 1602073617
transform -1 0 2608 0 -1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_118
timestamp 1602073617
transform -1 0 3258 0 -1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_641
timestamp 1602073617
transform -1 0 3908 0 -1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_608
timestamp 1602073617
transform -1 0 4558 0 -1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_327
timestamp 1602073617
transform -1 0 5208 0 -1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_265
timestamp 1602073617
transform 1 0 5208 0 -1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_267
timestamp 1602073617
transform 1 0 5858 0 -1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_361
timestamp 1602073617
transform 1 0 6508 0 -1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_772
timestamp 1602073617
transform -1 0 7808 0 -1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_557
timestamp 1602073617
transform 1 0 7808 0 -1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_561
timestamp 1602073617
transform 1 0 8458 0 -1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_512
timestamp 1602073617
transform 1 0 9108 0 -1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_743
timestamp 1602073617
transform 1 0 9758 0 -1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_780
timestamp 1602073617
transform 1 0 10408 0 -1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_108
timestamp 1602073617
transform 1 0 11058 0 -1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_830
timestamp 1602073617
transform 1 0 11708 0 -1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_747
timestamp 1602073617
transform 1 0 12358 0 -1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_761
timestamp 1602073617
transform 1 0 8 0 1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_598
timestamp 1602073617
transform -1 0 1308 0 1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_589
timestamp 1602073617
transform -1 0 1958 0 1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_432
timestamp 1602073617
transform -1 0 2608 0 1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_229
timestamp 1602073617
transform 1 0 2608 0 1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_231
timestamp 1602073617
transform 1 0 3258 0 1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_329
timestamp 1602073617
transform 1 0 3908 0 1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_68
timestamp 1602073617
transform 1 0 4558 0 1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_266
timestamp 1602073617
transform 1 0 5208 0 1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_262
timestamp 1602073617
transform -1 0 6508 0 1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_487
timestamp 1602073617
transform 1 0 6508 0 1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_489
timestamp 1602073617
transform 1 0 7158 0 1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_744
timestamp 1602073617
transform 1 0 7808 0 1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_558
timestamp 1602073617
transform -1 0 9108 0 1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_284
timestamp 1602073617
transform -1 0 9758 0 1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_279
timestamp 1602073617
transform -1 0 10408 0 1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_746
timestamp 1602073617
transform 1 0 10408 0 1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_781
timestamp 1602073617
transform 1 0 11058 0 1 5010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_782
timestamp 1602073617
transform -1 0 12358 0 1 5010
box -4 -6 618 206
use FILL  FILL_26_1
timestamp 1602073617
transform 1 0 12358 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_2
timestamp 1602073617
transform 1 0 12374 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_3
timestamp 1602073617
transform 1 0 12390 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_4
timestamp 1602073617
transform 1 0 12406 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_5
timestamp 1602073617
transform 1 0 12422 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_6
timestamp 1602073617
transform 1 0 12438 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_7
timestamp 1602073617
transform 1 0 12454 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_8
timestamp 1602073617
transform 1 0 12470 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_10
timestamp 1602073617
transform 1 0 12502 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_9
timestamp 1602073617
transform 1 0 12486 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_11
timestamp 1602073617
transform 1 0 12518 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_13
timestamp 1602073617
transform 1 0 12550 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_12
timestamp 1602073617
transform 1 0 12534 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_14
timestamp 1602073617
transform 1 0 12566 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_16
timestamp 1602073617
transform 1 0 12598 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_15
timestamp 1602073617
transform 1 0 12582 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_17
timestamp 1602073617
transform 1 0 12614 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_19
timestamp 1602073617
transform 1 0 12646 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_18
timestamp 1602073617
transform 1 0 12630 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_21
timestamp 1602073617
transform 1 0 12678 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_20
timestamp 1602073617
transform 1 0 12662 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_22
timestamp 1602073617
transform 1 0 12694 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_24
timestamp 1602073617
transform 1 0 12726 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_23
timestamp 1602073617
transform 1 0 12710 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_25
timestamp 1602073617
transform 1 0 12742 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_27
timestamp 1602073617
transform 1 0 12774 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_26
timestamp 1602073617
transform 1 0 12758 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_28
timestamp 1602073617
transform 1 0 12790 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_30
timestamp 1602073617
transform 1 0 12822 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_29
timestamp 1602073617
transform 1 0 12806 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_31
timestamp 1602073617
transform 1 0 12838 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_33
timestamp 1602073617
transform 1 0 12870 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_32
timestamp 1602073617
transform 1 0 12854 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_34
timestamp 1602073617
transform 1 0 12886 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_36
timestamp 1602073617
transform 1 0 12918 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_35
timestamp 1602073617
transform 1 0 12902 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_37
timestamp 1602073617
transform 1 0 12934 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_39
timestamp 1602073617
transform 1 0 12966 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_38
timestamp 1602073617
transform 1 0 12950 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_40
timestamp 1602073617
transform 1 0 12982 0 1 5010
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_810
timestamp 1602073617
transform 1 0 8 0 -1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_599
timestamp 1602073617
transform -1 0 1308 0 -1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_398
timestamp 1602073617
transform -1 0 1958 0 -1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_435
timestamp 1602073617
transform -1 0 2608 0 -1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_634
timestamp 1602073617
transform 1 0 2608 0 -1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_606
timestamp 1602073617
transform -1 0 3908 0 -1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_609
timestamp 1602073617
transform -1 0 4558 0 -1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_405
timestamp 1602073617
transform 1 0 4558 0 -1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_406
timestamp 1602073617
transform 1 0 5208 0 -1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_734
timestamp 1602073617
transform 1 0 5858 0 -1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_807
timestamp 1602073617
transform -1 0 7158 0 -1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_48
timestamp 1602073617
transform 1 0 7158 0 -1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_196
timestamp 1602073617
transform -1 0 8458 0 -1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_717
timestamp 1602073617
transform -1 0 9108 0 -1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_493
timestamp 1602073617
transform -1 0 9758 0 -1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_491
timestamp 1602073617
transform -1 0 10408 0 -1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_179
timestamp 1602073617
transform 1 0 10408 0 -1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_181
timestamp 1602073617
transform -1 0 11708 0 -1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_178
timestamp 1602073617
transform 1 0 11708 0 -1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_540
timestamp 1602073617
transform 1 0 12358 0 -1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_812
timestamp 1602073617
transform -1 0 658 0 1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_801
timestamp 1602073617
transform -1 0 1308 0 1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_676
timestamp 1602073617
transform -1 0 1958 0 1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_688
timestamp 1602073617
transform -1 0 2608 0 1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_290
timestamp 1602073617
transform -1 0 3258 0 1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_433
timestamp 1602073617
transform -1 0 3908 0 1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_479
timestamp 1602073617
transform -1 0 4558 0 1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_188
timestamp 1602073617
transform 1 0 4558 0 1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_475
timestamp 1602073617
transform -1 0 5858 0 1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_811
timestamp 1602073617
transform -1 0 6508 0 1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_474
timestamp 1602073617
transform -1 0 7158 0 1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_392
timestamp 1602073617
transform -1 0 7808 0 1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_45
timestamp 1602073617
transform 1 0 7808 0 1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_702
timestamp 1602073617
transform 1 0 8458 0 1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_492
timestamp 1602073617
transform 1 0 9108 0 1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_465
timestamp 1602073617
transform -1 0 10408 0 1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_146
timestamp 1602073617
transform 1 0 10408 0 1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_745
timestamp 1602073617
transform -1 0 11708 0 1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_803
timestamp 1602073617
transform 1 0 11708 0 1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_808
timestamp 1602073617
transform 1 0 12358 0 1 5410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_809
timestamp 1602073617
transform -1 0 658 0 -1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_399
timestamp 1602073617
transform -1 0 1308 0 -1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_681
timestamp 1602073617
transform -1 0 1958 0 -1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_643
timestamp 1602073617
transform -1 0 2608 0 -1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_595
timestamp 1602073617
transform -1 0 3258 0 -1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_611
timestamp 1602073617
transform -1 0 3908 0 -1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_355
timestamp 1602073617
transform -1 0 4558 0 -1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_331
timestamp 1602073617
transform -1 0 5208 0 -1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_186
timestamp 1602073617
transform -1 0 5858 0 -1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_80
timestamp 1602073617
transform 1 0 5858 0 -1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_501
timestamp 1602073617
transform -1 0 7158 0 -1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_498
timestamp 1602073617
transform -1 0 7808 0 -1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_151
timestamp 1602073617
transform 1 0 7808 0 -1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_374
timestamp 1602073617
transform 1 0 8458 0 -1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_698
timestamp 1602073617
transform 1 0 9108 0 -1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_709
timestamp 1602073617
transform 1 0 9758 0 -1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_145
timestamp 1602073617
transform 1 0 10408 0 -1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_148
timestamp 1602073617
transform 1 0 11058 0 -1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_797
timestamp 1602073617
transform -1 0 12358 0 -1 5810
box -4 -6 618 206
use FILL  FILL_29_1
timestamp 1602073617
transform -1 0 12374 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_2
timestamp 1602073617
transform -1 0 12390 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_3
timestamp 1602073617
transform -1 0 12406 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_4
timestamp 1602073617
transform -1 0 12422 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_5
timestamp 1602073617
transform -1 0 12438 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_6
timestamp 1602073617
transform -1 0 12454 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_7
timestamp 1602073617
transform -1 0 12470 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_8
timestamp 1602073617
transform -1 0 12486 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_10
timestamp 1602073617
transform -1 0 12518 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_9
timestamp 1602073617
transform -1 0 12502 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_11
timestamp 1602073617
transform -1 0 12534 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_13
timestamp 1602073617
transform -1 0 12566 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_12
timestamp 1602073617
transform -1 0 12550 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_14
timestamp 1602073617
transform -1 0 12582 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_16
timestamp 1602073617
transform -1 0 12614 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_15
timestamp 1602073617
transform -1 0 12598 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_17
timestamp 1602073617
transform -1 0 12630 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_19
timestamp 1602073617
transform -1 0 12662 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_18
timestamp 1602073617
transform -1 0 12646 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_21
timestamp 1602073617
transform -1 0 12694 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_20
timestamp 1602073617
transform -1 0 12678 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_22
timestamp 1602073617
transform -1 0 12710 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_24
timestamp 1602073617
transform -1 0 12742 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_23
timestamp 1602073617
transform -1 0 12726 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_25
timestamp 1602073617
transform -1 0 12758 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_27
timestamp 1602073617
transform -1 0 12790 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_26
timestamp 1602073617
transform -1 0 12774 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_28
timestamp 1602073617
transform -1 0 12806 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_30
timestamp 1602073617
transform -1 0 12838 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_29
timestamp 1602073617
transform -1 0 12822 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_31
timestamp 1602073617
transform -1 0 12854 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_33
timestamp 1602073617
transform -1 0 12886 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_32
timestamp 1602073617
transform -1 0 12870 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_34
timestamp 1602073617
transform -1 0 12902 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_36
timestamp 1602073617
transform -1 0 12934 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_35
timestamp 1602073617
transform -1 0 12918 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_37
timestamp 1602073617
transform -1 0 12950 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_39
timestamp 1602073617
transform -1 0 12982 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_38
timestamp 1602073617
transform -1 0 12966 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_40
timestamp 1602073617
transform -1 0 12998 0 -1 5810
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_679
timestamp 1602073617
transform -1 0 658 0 1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_403
timestamp 1602073617
transform 1 0 658 0 1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_394
timestamp 1602073617
transform -1 0 1958 0 1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_389
timestamp 1602073617
transform 1 0 1958 0 1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_334
timestamp 1602073617
transform 1 0 2608 0 1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_291
timestamp 1602073617
transform -1 0 3908 0 1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_330
timestamp 1602073617
transform 1 0 3908 0 1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_65
timestamp 1602073617
transform -1 0 5208 0 1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_404
timestamp 1602073617
transform 1 0 5208 0 1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_573
timestamp 1602073617
transform 1 0 5858 0 1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_735
timestamp 1602073617
transform 1 0 6508 0 1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_575
timestamp 1602073617
transform 1 0 7158 0 1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_579
timestamp 1602073617
transform 1 0 7808 0 1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_322
timestamp 1602073617
transform -1 0 9108 0 1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_701
timestamp 1602073617
transform 1 0 9108 0 1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_142
timestamp 1602073617
transform 1 0 9758 0 1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_144
timestamp 1602073617
transform 1 0 10408 0 1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_147
timestamp 1602073617
transform 1 0 11058 0 1 5810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_149
timestamp 1602073617
transform 1 0 11708 0 1 5810
box -4 -6 618 206
use FILL  FILL_30_1
timestamp 1602073617
transform 1 0 12358 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_2
timestamp 1602073617
transform 1 0 12374 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_3
timestamp 1602073617
transform 1 0 12390 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_4
timestamp 1602073617
transform 1 0 12406 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_5
timestamp 1602073617
transform 1 0 12422 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_6
timestamp 1602073617
transform 1 0 12438 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_7
timestamp 1602073617
transform 1 0 12454 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_8
timestamp 1602073617
transform 1 0 12470 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_10
timestamp 1602073617
transform 1 0 12502 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_9
timestamp 1602073617
transform 1 0 12486 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_11
timestamp 1602073617
transform 1 0 12518 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_13
timestamp 1602073617
transform 1 0 12550 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_12
timestamp 1602073617
transform 1 0 12534 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_14
timestamp 1602073617
transform 1 0 12566 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_16
timestamp 1602073617
transform 1 0 12598 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_15
timestamp 1602073617
transform 1 0 12582 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_17
timestamp 1602073617
transform 1 0 12614 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_19
timestamp 1602073617
transform 1 0 12646 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_18
timestamp 1602073617
transform 1 0 12630 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_21
timestamp 1602073617
transform 1 0 12678 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_20
timestamp 1602073617
transform 1 0 12662 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_22
timestamp 1602073617
transform 1 0 12694 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_24
timestamp 1602073617
transform 1 0 12726 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_23
timestamp 1602073617
transform 1 0 12710 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_25
timestamp 1602073617
transform 1 0 12742 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_27
timestamp 1602073617
transform 1 0 12774 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_26
timestamp 1602073617
transform 1 0 12758 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_28
timestamp 1602073617
transform 1 0 12790 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_30
timestamp 1602073617
transform 1 0 12822 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_29
timestamp 1602073617
transform 1 0 12806 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_31
timestamp 1602073617
transform 1 0 12838 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_33
timestamp 1602073617
transform 1 0 12870 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_32
timestamp 1602073617
transform 1 0 12854 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_34
timestamp 1602073617
transform 1 0 12886 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_36
timestamp 1602073617
transform 1 0 12918 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_35
timestamp 1602073617
transform 1 0 12902 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_37
timestamp 1602073617
transform 1 0 12934 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_39
timestamp 1602073617
transform 1 0 12966 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_38
timestamp 1602073617
transform 1 0 12950 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_40
timestamp 1602073617
transform 1 0 12982 0 1 5810
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_691
timestamp 1602073617
transform -1 0 658 0 -1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_689
timestamp 1602073617
transform -1 0 1308 0 -1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_400
timestamp 1602073617
transform -1 0 1958 0 -1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_393
timestamp 1602073617
transform -1 0 2608 0 -1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_537
timestamp 1602073617
transform -1 0 3258 0 -1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_607
timestamp 1602073617
transform 1 0 3258 0 -1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_57
timestamp 1602073617
transform 1 0 3908 0 -1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_198
timestamp 1602073617
transform 1 0 4558 0 -1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_101
timestamp 1602073617
transform -1 0 5858 0 -1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_99
timestamp 1602073617
transform -1 0 6508 0 -1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_397
timestamp 1602073617
transform 1 0 6508 0 -1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_83
timestamp 1602073617
transform -1 0 7808 0 -1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_390
timestamp 1602073617
transform -1 0 8458 0 -1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_310
timestamp 1602073617
transform 1 0 8458 0 -1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_388
timestamp 1602073617
transform -1 0 9758 0 -1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_167
timestamp 1602073617
transform -1 0 10408 0 -1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_700
timestamp 1602073617
transform 1 0 10408 0 -1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_710
timestamp 1602073617
transform 1 0 11058 0 -1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_711
timestamp 1602073617
transform 1 0 11708 0 -1 6210
box -4 -6 618 206
use FILL  FILL_31_1
timestamp 1602073617
transform -1 0 12374 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_2
timestamp 1602073617
transform -1 0 12390 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_3
timestamp 1602073617
transform -1 0 12406 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_4
timestamp 1602073617
transform -1 0 12422 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_5
timestamp 1602073617
transform -1 0 12438 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_6
timestamp 1602073617
transform -1 0 12454 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_7
timestamp 1602073617
transform -1 0 12470 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_8
timestamp 1602073617
transform -1 0 12486 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_10
timestamp 1602073617
transform -1 0 12518 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_9
timestamp 1602073617
transform -1 0 12502 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_11
timestamp 1602073617
transform -1 0 12534 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_13
timestamp 1602073617
transform -1 0 12566 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_12
timestamp 1602073617
transform -1 0 12550 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_14
timestamp 1602073617
transform -1 0 12582 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_16
timestamp 1602073617
transform -1 0 12614 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_15
timestamp 1602073617
transform -1 0 12598 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_17
timestamp 1602073617
transform -1 0 12630 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_19
timestamp 1602073617
transform -1 0 12662 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_18
timestamp 1602073617
transform -1 0 12646 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_21
timestamp 1602073617
transform -1 0 12694 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_20
timestamp 1602073617
transform -1 0 12678 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_22
timestamp 1602073617
transform -1 0 12710 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_24
timestamp 1602073617
transform -1 0 12742 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_23
timestamp 1602073617
transform -1 0 12726 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_25
timestamp 1602073617
transform -1 0 12758 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_27
timestamp 1602073617
transform -1 0 12790 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_26
timestamp 1602073617
transform -1 0 12774 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_28
timestamp 1602073617
transform -1 0 12806 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_30
timestamp 1602073617
transform -1 0 12838 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_29
timestamp 1602073617
transform -1 0 12822 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_31
timestamp 1602073617
transform -1 0 12854 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_33
timestamp 1602073617
transform -1 0 12886 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_32
timestamp 1602073617
transform -1 0 12870 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_34
timestamp 1602073617
transform -1 0 12902 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_36
timestamp 1602073617
transform -1 0 12934 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_35
timestamp 1602073617
transform -1 0 12918 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_37
timestamp 1602073617
transform -1 0 12950 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_39
timestamp 1602073617
transform -1 0 12982 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_38
timestamp 1602073617
transform -1 0 12966 0 -1 6210
box -4 -6 20 206
use FILL  FILL_31_40
timestamp 1602073617
transform -1 0 12998 0 -1 6210
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_687
timestamp 1602073617
transform -1 0 658 0 1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_685
timestamp 1602073617
transform -1 0 1308 0 1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_684
timestamp 1602073617
transform -1 0 1958 0 1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_385
timestamp 1602073617
transform 1 0 1958 0 1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_536
timestamp 1602073617
transform 1 0 2608 0 1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_646
timestamp 1602073617
transform -1 0 3908 0 1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_197
timestamp 1602073617
transform 1 0 3908 0 1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_52
timestamp 1602073617
transform -1 0 5208 0 1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_216
timestamp 1602073617
transform 1 0 5208 0 1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_218
timestamp 1602073617
transform 1 0 5858 0 1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_402
timestamp 1602073617
transform -1 0 7158 0 1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_704
timestamp 1602073617
transform 1 0 7158 0 1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_325
timestamp 1602073617
transform -1 0 8458 0 1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_323
timestamp 1602073617
transform -1 0 9108 0 1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_703
timestamp 1602073617
transform 1 0 9108 0 1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_714
timestamp 1602073617
transform 1 0 9758 0 1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_724
timestamp 1602073617
transform 1 0 10408 0 1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_732
timestamp 1602073617
transform 1 0 11058 0 1 6210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_209
timestamp 1602073617
transform -1 0 12358 0 1 6210
box -4 -6 618 206
use FILL  FILL_32_1
timestamp 1602073617
transform 1 0 12358 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_2
timestamp 1602073617
transform 1 0 12374 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_3
timestamp 1602073617
transform 1 0 12390 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_4
timestamp 1602073617
transform 1 0 12406 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_5
timestamp 1602073617
transform 1 0 12422 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_6
timestamp 1602073617
transform 1 0 12438 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_7
timestamp 1602073617
transform 1 0 12454 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_8
timestamp 1602073617
transform 1 0 12470 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_10
timestamp 1602073617
transform 1 0 12502 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_9
timestamp 1602073617
transform 1 0 12486 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_11
timestamp 1602073617
transform 1 0 12518 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_13
timestamp 1602073617
transform 1 0 12550 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_12
timestamp 1602073617
transform 1 0 12534 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_14
timestamp 1602073617
transform 1 0 12566 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_16
timestamp 1602073617
transform 1 0 12598 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_15
timestamp 1602073617
transform 1 0 12582 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_17
timestamp 1602073617
transform 1 0 12614 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_19
timestamp 1602073617
transform 1 0 12646 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_18
timestamp 1602073617
transform 1 0 12630 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_21
timestamp 1602073617
transform 1 0 12678 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_20
timestamp 1602073617
transform 1 0 12662 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_22
timestamp 1602073617
transform 1 0 12694 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_24
timestamp 1602073617
transform 1 0 12726 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_23
timestamp 1602073617
transform 1 0 12710 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_25
timestamp 1602073617
transform 1 0 12742 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_27
timestamp 1602073617
transform 1 0 12774 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_26
timestamp 1602073617
transform 1 0 12758 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_28
timestamp 1602073617
transform 1 0 12790 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_30
timestamp 1602073617
transform 1 0 12822 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_29
timestamp 1602073617
transform 1 0 12806 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_31
timestamp 1602073617
transform 1 0 12838 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_33
timestamp 1602073617
transform 1 0 12870 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_32
timestamp 1602073617
transform 1 0 12854 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_34
timestamp 1602073617
transform 1 0 12886 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_36
timestamp 1602073617
transform 1 0 12918 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_35
timestamp 1602073617
transform 1 0 12902 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_37
timestamp 1602073617
transform 1 0 12934 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_39
timestamp 1602073617
transform 1 0 12966 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_38
timestamp 1602073617
transform 1 0 12950 0 1 6210
box -4 -6 20 206
use FILL  FILL_32_40
timestamp 1602073617
transform 1 0 12982 0 1 6210
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_800
timestamp 1602073617
transform 1 0 8 0 -1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_686
timestamp 1602073617
transform -1 0 1308 0 -1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_683
timestamp 1602073617
transform -1 0 1958 0 -1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_604
timestamp 1602073617
transform -1 0 2608 0 -1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_610
timestamp 1602073617
transform 1 0 2608 0 -1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_612
timestamp 1602073617
transform 1 0 3258 0 -1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_647
timestamp 1602073617
transform 1 0 3908 0 -1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_656
timestamp 1602073617
transform -1 0 5208 0 -1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_89
timestamp 1602073617
transform 1 0 5208 0 -1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_97
timestamp 1602073617
transform 1 0 5858 0 -1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_396
timestamp 1602073617
transform 1 0 6508 0 -1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_401
timestamp 1602073617
transform -1 0 7808 0 -1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_395
timestamp 1602073617
transform -1 0 8458 0 -1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_332
timestamp 1602073617
transform -1 0 9108 0 -1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_111
timestamp 1602073617
transform -1 0 9758 0 -1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_312
timestamp 1602073617
transform -1 0 10408 0 -1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_715
timestamp 1602073617
transform -1 0 11058 0 -1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_112
timestamp 1602073617
transform -1 0 11708 0 -1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_213
timestamp 1602073617
transform 1 0 11708 0 -1 6610
box -4 -6 618 206
use FILL  FILL_33_1
timestamp 1602073617
transform -1 0 12374 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_2
timestamp 1602073617
transform -1 0 12390 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_3
timestamp 1602073617
transform -1 0 12406 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_4
timestamp 1602073617
transform -1 0 12422 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_5
timestamp 1602073617
transform -1 0 12438 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_6
timestamp 1602073617
transform -1 0 12454 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_7
timestamp 1602073617
transform -1 0 12470 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_8
timestamp 1602073617
transform -1 0 12486 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_10
timestamp 1602073617
transform -1 0 12518 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_9
timestamp 1602073617
transform -1 0 12502 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_11
timestamp 1602073617
transform -1 0 12534 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_13
timestamp 1602073617
transform -1 0 12566 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_12
timestamp 1602073617
transform -1 0 12550 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_14
timestamp 1602073617
transform -1 0 12582 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_16
timestamp 1602073617
transform -1 0 12614 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_15
timestamp 1602073617
transform -1 0 12598 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_17
timestamp 1602073617
transform -1 0 12630 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_19
timestamp 1602073617
transform -1 0 12662 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_18
timestamp 1602073617
transform -1 0 12646 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_21
timestamp 1602073617
transform -1 0 12694 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_20
timestamp 1602073617
transform -1 0 12678 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_22
timestamp 1602073617
transform -1 0 12710 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_24
timestamp 1602073617
transform -1 0 12742 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_23
timestamp 1602073617
transform -1 0 12726 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_25
timestamp 1602073617
transform -1 0 12758 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_27
timestamp 1602073617
transform -1 0 12790 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_26
timestamp 1602073617
transform -1 0 12774 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_28
timestamp 1602073617
transform -1 0 12806 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_30
timestamp 1602073617
transform -1 0 12838 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_29
timestamp 1602073617
transform -1 0 12822 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_31
timestamp 1602073617
transform -1 0 12854 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_33
timestamp 1602073617
transform -1 0 12886 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_32
timestamp 1602073617
transform -1 0 12870 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_34
timestamp 1602073617
transform -1 0 12902 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_36
timestamp 1602073617
transform -1 0 12934 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_35
timestamp 1602073617
transform -1 0 12918 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_37
timestamp 1602073617
transform -1 0 12950 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_39
timestamp 1602073617
transform -1 0 12982 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_38
timestamp 1602073617
transform -1 0 12966 0 -1 6610
box -4 -6 20 206
use FILL  FILL_33_40
timestamp 1602073617
transform -1 0 12998 0 -1 6610
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_729
timestamp 1602073617
transform 1 0 8 0 1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_682
timestamp 1602073617
transform -1 0 1308 0 1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_603
timestamp 1602073617
transform 1 0 1308 0 1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_605
timestamp 1602073617
transform 1 0 1958 0 1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_60
timestamp 1602073617
transform 1 0 2608 0 1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_58
timestamp 1602073617
transform 1 0 3258 0 1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_61
timestamp 1602073617
transform 1 0 3908 0 1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_201
timestamp 1602073617
transform 1 0 4558 0 1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_206
timestamp 1602073617
transform 1 0 5208 0 1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_84
timestamp 1602073617
transform -1 0 6508 0 1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_81
timestamp 1602073617
transform -1 0 7158 0 1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_299
timestamp 1602073617
transform 1 0 7158 0 1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_316
timestamp 1602073617
transform 1 0 7808 0 1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_166
timestamp 1602073617
transform 1 0 8458 0 1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_169
timestamp 1602073617
transform 1 0 9108 0 1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_280
timestamp 1602073617
transform 1 0 9758 0 1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_542
timestamp 1602073617
transform 1 0 10408 0 1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_109
timestamp 1602073617
transform 1 0 11058 0 1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_152
timestamp 1602073617
transform -1 0 12358 0 1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_569
timestamp 1602073617
transform 1 0 12358 0 1 6610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_760
timestamp 1602073617
transform -1 0 658 0 -1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_728
timestamp 1602073617
transform 1 0 8 0 1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_593
timestamp 1602073617
transform -1 0 1308 0 -1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_645
timestamp 1602073617
transform -1 0 1308 0 1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_601
timestamp 1602073617
transform -1 0 1958 0 -1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_602
timestamp 1602073617
transform -1 0 1958 0 1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_718
timestamp 1602073617
transform 1 0 1958 0 -1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_600
timestamp 1602073617
transform -1 0 2608 0 1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_722
timestamp 1602073617
transform 1 0 2608 0 -1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_591
timestamp 1602073617
transform -1 0 3258 0 1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_733
timestamp 1602073617
transform 1 0 3258 0 -1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_590
timestamp 1602073617
transform -1 0 3908 0 1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_339
timestamp 1602073617
transform -1 0 4558 0 -1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_39
timestamp 1602073617
transform -1 0 4558 0 1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_737
timestamp 1602073617
transform 1 0 4558 0 -1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_319
timestamp 1602073617
transform -1 0 5208 0 1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_314
timestamp 1602073617
transform 1 0 5208 0 -1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_7
timestamp 1602073617
transform 1 0 5208 0 1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_786
timestamp 1602073617
transform 1 0 5858 0 -1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_317
timestamp 1602073617
transform -1 0 6508 0 1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_298
timestamp 1602073617
transform 1 0 6508 0 -1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_313
timestamp 1602073617
transform -1 0 7158 0 1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_302
timestamp 1602073617
transform 1 0 7158 0 -1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_369
timestamp 1602073617
transform 1 0 7158 0 1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_318
timestamp 1602073617
transform -1 0 8458 0 -1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_306
timestamp 1602073617
transform -1 0 8458 0 1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_315
timestamp 1602073617
transform 1 0 8458 0 -1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_74
timestamp 1602073617
transform 1 0 8458 0 1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_543
timestamp 1602073617
transform 1 0 9108 0 -1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_76
timestamp 1602073617
transform 1 0 9108 0 1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_373
timestamp 1602073617
transform 1 0 9758 0 -1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_455
timestamp 1602073617
transform 1 0 9758 0 1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_524
timestamp 1602073617
transform 1 0 10408 0 -1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_544
timestamp 1602073617
transform 1 0 10408 0 1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_552
timestamp 1602073617
transform 1 0 11058 0 -1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_551
timestamp 1602073617
transform 1 0 11058 0 1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_577
timestamp 1602073617
transform -1 0 12358 0 -1 7010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_564
timestamp 1602073617
transform 1 0 11708 0 1 7010
box -4 -6 618 206
use FILL  FILL_36_1
timestamp 1602073617
transform 1 0 12358 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_1
timestamp 1602073617
transform -1 0 12374 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_4
timestamp 1602073617
transform 1 0 12406 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_3
timestamp 1602073617
transform 1 0 12390 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_2
timestamp 1602073617
transform 1 0 12374 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_4
timestamp 1602073617
transform -1 0 12422 0 -1 7010
box -4 -6 20 206
use FILL  FILL_35_3
timestamp 1602073617
transform -1 0 12406 0 -1 7010
box -4 -6 20 206
use FILL  FILL_35_2
timestamp 1602073617
transform -1 0 12390 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_7
timestamp 1602073617
transform 1 0 12454 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_6
timestamp 1602073617
transform 1 0 12438 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_5
timestamp 1602073617
transform 1 0 12422 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_7
timestamp 1602073617
transform -1 0 12470 0 -1 7010
box -4 -6 20 206
use FILL  FILL_35_6
timestamp 1602073617
transform -1 0 12454 0 -1 7010
box -4 -6 20 206
use FILL  FILL_35_5
timestamp 1602073617
transform -1 0 12438 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_8
timestamp 1602073617
transform 1 0 12470 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_8
timestamp 1602073617
transform -1 0 12486 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_10
timestamp 1602073617
transform 1 0 12502 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_9
timestamp 1602073617
transform 1 0 12486 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_10
timestamp 1602073617
transform -1 0 12518 0 -1 7010
box -4 -6 20 206
use FILL  FILL_35_9
timestamp 1602073617
transform -1 0 12502 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_11
timestamp 1602073617
transform 1 0 12518 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_11
timestamp 1602073617
transform -1 0 12534 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_13
timestamp 1602073617
transform 1 0 12550 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_12
timestamp 1602073617
transform 1 0 12534 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_13
timestamp 1602073617
transform -1 0 12566 0 -1 7010
box -4 -6 20 206
use FILL  FILL_35_12
timestamp 1602073617
transform -1 0 12550 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_14
timestamp 1602073617
transform 1 0 12566 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_14
timestamp 1602073617
transform -1 0 12582 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_16
timestamp 1602073617
transform 1 0 12598 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_15
timestamp 1602073617
transform 1 0 12582 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_16
timestamp 1602073617
transform -1 0 12614 0 -1 7010
box -4 -6 20 206
use FILL  FILL_35_15
timestamp 1602073617
transform -1 0 12598 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_17
timestamp 1602073617
transform 1 0 12614 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_17
timestamp 1602073617
transform -1 0 12630 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_19
timestamp 1602073617
transform 1 0 12646 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_18
timestamp 1602073617
transform 1 0 12630 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_19
timestamp 1602073617
transform -1 0 12662 0 -1 7010
box -4 -6 20 206
use FILL  FILL_35_18
timestamp 1602073617
transform -1 0 12646 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_21
timestamp 1602073617
transform 1 0 12678 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_20
timestamp 1602073617
transform 1 0 12662 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_21
timestamp 1602073617
transform -1 0 12694 0 -1 7010
box -4 -6 20 206
use FILL  FILL_35_20
timestamp 1602073617
transform -1 0 12678 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_22
timestamp 1602073617
transform 1 0 12694 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_22
timestamp 1602073617
transform -1 0 12710 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_24
timestamp 1602073617
transform 1 0 12726 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_23
timestamp 1602073617
transform 1 0 12710 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_24
timestamp 1602073617
transform -1 0 12742 0 -1 7010
box -4 -6 20 206
use FILL  FILL_35_23
timestamp 1602073617
transform -1 0 12726 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_25
timestamp 1602073617
transform 1 0 12742 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_25
timestamp 1602073617
transform -1 0 12758 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_27
timestamp 1602073617
transform 1 0 12774 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_26
timestamp 1602073617
transform 1 0 12758 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_27
timestamp 1602073617
transform -1 0 12790 0 -1 7010
box -4 -6 20 206
use FILL  FILL_35_26
timestamp 1602073617
transform -1 0 12774 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_28
timestamp 1602073617
transform 1 0 12790 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_28
timestamp 1602073617
transform -1 0 12806 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_30
timestamp 1602073617
transform 1 0 12822 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_29
timestamp 1602073617
transform 1 0 12806 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_30
timestamp 1602073617
transform -1 0 12838 0 -1 7010
box -4 -6 20 206
use FILL  FILL_35_29
timestamp 1602073617
transform -1 0 12822 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_31
timestamp 1602073617
transform 1 0 12838 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_31
timestamp 1602073617
transform -1 0 12854 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_33
timestamp 1602073617
transform 1 0 12870 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_32
timestamp 1602073617
transform 1 0 12854 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_33
timestamp 1602073617
transform -1 0 12886 0 -1 7010
box -4 -6 20 206
use FILL  FILL_35_32
timestamp 1602073617
transform -1 0 12870 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_34
timestamp 1602073617
transform 1 0 12886 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_34
timestamp 1602073617
transform -1 0 12902 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_36
timestamp 1602073617
transform 1 0 12918 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_35
timestamp 1602073617
transform 1 0 12902 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_36
timestamp 1602073617
transform -1 0 12934 0 -1 7010
box -4 -6 20 206
use FILL  FILL_35_35
timestamp 1602073617
transform -1 0 12918 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_37
timestamp 1602073617
transform 1 0 12934 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_37
timestamp 1602073617
transform -1 0 12950 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_39
timestamp 1602073617
transform 1 0 12966 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_38
timestamp 1602073617
transform 1 0 12950 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_39
timestamp 1602073617
transform -1 0 12982 0 -1 7010
box -4 -6 20 206
use FILL  FILL_35_38
timestamp 1602073617
transform -1 0 12966 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_40
timestamp 1602073617
transform 1 0 12982 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_40
timestamp 1602073617
transform -1 0 12998 0 -1 7010
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_730
timestamp 1602073617
transform -1 0 658 0 -1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_644
timestamp 1602073617
transform -1 0 1308 0 -1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_597
timestamp 1602073617
transform -1 0 1958 0 -1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_539
timestamp 1602073617
transform -1 0 2608 0 -1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_532
timestamp 1602073617
transform -1 0 3258 0 -1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_16
timestamp 1602073617
transform 1 0 3258 0 -1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_194
timestamp 1602073617
transform 1 0 3908 0 -1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_341
timestamp 1602073617
transform -1 0 5208 0 -1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_228
timestamp 1602073617
transform -1 0 5858 0 -1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_723
timestamp 1602073617
transform -1 0 6508 0 -1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_824
timestamp 1602073617
transform 1 0 6508 0 -1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_43
timestamp 1602073617
transform -1 0 7808 0 -1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_308
timestamp 1602073617
transform 1 0 7808 0 -1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_309
timestamp 1602073617
transform 1 0 8458 0 -1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_370
timestamp 1602073617
transform 1 0 9108 0 -1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_445
timestamp 1602073617
transform -1 0 10408 0 -1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_241
timestamp 1602073617
transform 1 0 10408 0 -1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_787
timestamp 1602073617
transform -1 0 11708 0 -1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_726
timestamp 1602073617
transform 1 0 11708 0 -1 7410
box -4 -6 618 206
use FILL  FILL_37_1
timestamp 1602073617
transform -1 0 12374 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_2
timestamp 1602073617
transform -1 0 12390 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_3
timestamp 1602073617
transform -1 0 12406 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_4
timestamp 1602073617
transform -1 0 12422 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_5
timestamp 1602073617
transform -1 0 12438 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_6
timestamp 1602073617
transform -1 0 12454 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_7
timestamp 1602073617
transform -1 0 12470 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_8
timestamp 1602073617
transform -1 0 12486 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_10
timestamp 1602073617
transform -1 0 12518 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_9
timestamp 1602073617
transform -1 0 12502 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_11
timestamp 1602073617
transform -1 0 12534 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_13
timestamp 1602073617
transform -1 0 12566 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_12
timestamp 1602073617
transform -1 0 12550 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_14
timestamp 1602073617
transform -1 0 12582 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_16
timestamp 1602073617
transform -1 0 12614 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_15
timestamp 1602073617
transform -1 0 12598 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_17
timestamp 1602073617
transform -1 0 12630 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_19
timestamp 1602073617
transform -1 0 12662 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_18
timestamp 1602073617
transform -1 0 12646 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_21
timestamp 1602073617
transform -1 0 12694 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_20
timestamp 1602073617
transform -1 0 12678 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_22
timestamp 1602073617
transform -1 0 12710 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_24
timestamp 1602073617
transform -1 0 12742 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_23
timestamp 1602073617
transform -1 0 12726 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_25
timestamp 1602073617
transform -1 0 12758 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_27
timestamp 1602073617
transform -1 0 12790 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_26
timestamp 1602073617
transform -1 0 12774 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_28
timestamp 1602073617
transform -1 0 12806 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_30
timestamp 1602073617
transform -1 0 12838 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_29
timestamp 1602073617
transform -1 0 12822 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_31
timestamp 1602073617
transform -1 0 12854 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_33
timestamp 1602073617
transform -1 0 12886 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_32
timestamp 1602073617
transform -1 0 12870 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_34
timestamp 1602073617
transform -1 0 12902 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_36
timestamp 1602073617
transform -1 0 12934 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_35
timestamp 1602073617
transform -1 0 12918 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_37
timestamp 1602073617
transform -1 0 12950 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_39
timestamp 1602073617
transform -1 0 12982 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_38
timestamp 1602073617
transform -1 0 12966 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_40
timestamp 1602073617
transform -1 0 12998 0 -1 7410
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_829
timestamp 1602073617
transform 1 0 8 0 1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_648
timestamp 1602073617
transform 1 0 658 0 1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_788
timestamp 1602073617
transform 1 0 1308 0 1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_533
timestamp 1602073617
transform -1 0 2608 0 1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_24
timestamp 1602073617
transform 1 0 2608 0 1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_282
timestamp 1602073617
transform 1 0 3258 0 1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_350
timestamp 1602073617
transform 1 0 3908 0 1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_285
timestamp 1602073617
transform 1 0 4558 0 1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_281
timestamp 1602073617
transform -1 0 5858 0 1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_716
timestamp 1602073617
transform 1 0 5858 0 1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_836
timestamp 1602073617
transform -1 0 7158 0 1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_823
timestamp 1602073617
transform -1 0 7808 0 1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_301
timestamp 1602073617
transform 1 0 7808 0 1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_75
timestamp 1602073617
transform -1 0 9108 0 1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_187
timestamp 1602073617
transform 1 0 9108 0 1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_237
timestamp 1602073617
transform 1 0 9758 0 1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_191
timestamp 1602073617
transform 1 0 10408 0 1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_794
timestamp 1602073617
transform 1 0 11058 0 1 7410
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_804
timestamp 1602073617
transform 1 0 11708 0 1 7410
box -4 -6 618 206
use FILL  FILL_38_1
timestamp 1602073617
transform 1 0 12358 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_2
timestamp 1602073617
transform 1 0 12374 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_3
timestamp 1602073617
transform 1 0 12390 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_4
timestamp 1602073617
transform 1 0 12406 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_5
timestamp 1602073617
transform 1 0 12422 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_6
timestamp 1602073617
transform 1 0 12438 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_7
timestamp 1602073617
transform 1 0 12454 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_8
timestamp 1602073617
transform 1 0 12470 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_10
timestamp 1602073617
transform 1 0 12502 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_9
timestamp 1602073617
transform 1 0 12486 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_11
timestamp 1602073617
transform 1 0 12518 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_13
timestamp 1602073617
transform 1 0 12550 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_12
timestamp 1602073617
transform 1 0 12534 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_14
timestamp 1602073617
transform 1 0 12566 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_16
timestamp 1602073617
transform 1 0 12598 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_15
timestamp 1602073617
transform 1 0 12582 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_17
timestamp 1602073617
transform 1 0 12614 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_19
timestamp 1602073617
transform 1 0 12646 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_18
timestamp 1602073617
transform 1 0 12630 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_21
timestamp 1602073617
transform 1 0 12678 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_20
timestamp 1602073617
transform 1 0 12662 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_22
timestamp 1602073617
transform 1 0 12694 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_24
timestamp 1602073617
transform 1 0 12726 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_23
timestamp 1602073617
transform 1 0 12710 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_25
timestamp 1602073617
transform 1 0 12742 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_27
timestamp 1602073617
transform 1 0 12774 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_26
timestamp 1602073617
transform 1 0 12758 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_28
timestamp 1602073617
transform 1 0 12790 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_30
timestamp 1602073617
transform 1 0 12822 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_29
timestamp 1602073617
transform 1 0 12806 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_31
timestamp 1602073617
transform 1 0 12838 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_33
timestamp 1602073617
transform 1 0 12870 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_32
timestamp 1602073617
transform 1 0 12854 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_34
timestamp 1602073617
transform 1 0 12886 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_36
timestamp 1602073617
transform 1 0 12918 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_35
timestamp 1602073617
transform 1 0 12902 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_37
timestamp 1602073617
transform 1 0 12934 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_39
timestamp 1602073617
transform 1 0 12966 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_38
timestamp 1602073617
transform 1 0 12950 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_40
timestamp 1602073617
transform 1 0 12982 0 1 7410
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_480
timestamp 1602073617
transform -1 0 658 0 -1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_855
timestamp 1602073617
transform 1 0 658 0 -1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_660
timestamp 1602073617
transform -1 0 1958 0 -1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_655
timestamp 1602073617
transform -1 0 2608 0 -1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_535
timestamp 1602073617
transform -1 0 3258 0 -1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_534
timestamp 1602073617
transform -1 0 3908 0 -1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_838
timestamp 1602073617
transform 1 0 3908 0 -1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_827
timestamp 1602073617
transform -1 0 5208 0 -1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_193
timestamp 1602073617
transform -1 0 5858 0 -1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_538
timestamp 1602073617
transform -1 0 6508 0 -1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_283
timestamp 1602073617
transform 1 0 6508 0 -1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_286
timestamp 1602073617
transform 1 0 7158 0 -1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_288
timestamp 1602073617
transform 1 0 7808 0 -1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_362
timestamp 1602073617
transform 1 0 8458 0 -1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_176
timestamp 1602073617
transform 1 0 9108 0 -1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_311
timestamp 1602073617
transform 1 0 9758 0 -1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_336
timestamp 1602073617
transform 1 0 10408 0 -1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_545
timestamp 1602073617
transform -1 0 11708 0 -1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_165
timestamp 1602073617
transform 1 0 11708 0 -1 7810
box -4 -6 618 206
use FILL  FILL_39_1
timestamp 1602073617
transform -1 0 12374 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_2
timestamp 1602073617
transform -1 0 12390 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_3
timestamp 1602073617
transform -1 0 12406 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_4
timestamp 1602073617
transform -1 0 12422 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_5
timestamp 1602073617
transform -1 0 12438 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_6
timestamp 1602073617
transform -1 0 12454 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_7
timestamp 1602073617
transform -1 0 12470 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_8
timestamp 1602073617
transform -1 0 12486 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_10
timestamp 1602073617
transform -1 0 12518 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_9
timestamp 1602073617
transform -1 0 12502 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_11
timestamp 1602073617
transform -1 0 12534 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_13
timestamp 1602073617
transform -1 0 12566 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_12
timestamp 1602073617
transform -1 0 12550 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_14
timestamp 1602073617
transform -1 0 12582 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_16
timestamp 1602073617
transform -1 0 12614 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_15
timestamp 1602073617
transform -1 0 12598 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_17
timestamp 1602073617
transform -1 0 12630 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_19
timestamp 1602073617
transform -1 0 12662 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_18
timestamp 1602073617
transform -1 0 12646 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_21
timestamp 1602073617
transform -1 0 12694 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_20
timestamp 1602073617
transform -1 0 12678 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_22
timestamp 1602073617
transform -1 0 12710 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_24
timestamp 1602073617
transform -1 0 12742 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_23
timestamp 1602073617
transform -1 0 12726 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_25
timestamp 1602073617
transform -1 0 12758 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_27
timestamp 1602073617
transform -1 0 12790 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_26
timestamp 1602073617
transform -1 0 12774 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_28
timestamp 1602073617
transform -1 0 12806 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_30
timestamp 1602073617
transform -1 0 12838 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_29
timestamp 1602073617
transform -1 0 12822 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_31
timestamp 1602073617
transform -1 0 12854 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_33
timestamp 1602073617
transform -1 0 12886 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_32
timestamp 1602073617
transform -1 0 12870 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_34
timestamp 1602073617
transform -1 0 12902 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_36
timestamp 1602073617
transform -1 0 12934 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_35
timestamp 1602073617
transform -1 0 12918 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_37
timestamp 1602073617
transform -1 0 12950 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_39
timestamp 1602073617
transform -1 0 12982 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_38
timestamp 1602073617
transform -1 0 12966 0 -1 7810
box -4 -6 20 206
use FILL  FILL_39_40
timestamp 1602073617
transform -1 0 12998 0 -1 7810
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_680
timestamp 1602073617
transform -1 0 658 0 1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_444
timestamp 1602073617
transform -1 0 1308 0 1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_442
timestamp 1602073617
transform -1 0 1958 0 1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_567
timestamp 1602073617
transform 1 0 1958 0 1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_171
timestamp 1602073617
transform -1 0 3258 0 1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_289
timestamp 1602073617
transform -1 0 3908 0 1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_822
timestamp 1602073617
transform 1 0 3908 0 1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_200
timestamp 1602073617
transform 1 0 4558 0 1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_13
timestamp 1602073617
transform 1 0 5208 0 1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_438
timestamp 1602073617
transform 1 0 5858 0 1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_41
timestamp 1602073617
transform 1 0 6508 0 1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_806
timestamp 1602073617
transform -1 0 7808 0 1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_238
timestamp 1602073617
transform 1 0 7808 0 1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_366
timestamp 1602073617
transform -1 0 9108 0 1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_335
timestamp 1602073617
transform 1 0 9108 0 1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_180
timestamp 1602073617
transform 1 0 9758 0 1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_443
timestamp 1602073617
transform -1 0 11058 0 1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_441
timestamp 1602073617
transform 1 0 11058 0 1 7810
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_795
timestamp 1602073617
transform -1 0 12358 0 1 7810
box -4 -6 618 206
use FILL  FILL_40_1
timestamp 1602073617
transform 1 0 12358 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_2
timestamp 1602073617
transform 1 0 12374 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_3
timestamp 1602073617
transform 1 0 12390 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_4
timestamp 1602073617
transform 1 0 12406 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_5
timestamp 1602073617
transform 1 0 12422 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_6
timestamp 1602073617
transform 1 0 12438 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_7
timestamp 1602073617
transform 1 0 12454 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_8
timestamp 1602073617
transform 1 0 12470 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_10
timestamp 1602073617
transform 1 0 12502 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_9
timestamp 1602073617
transform 1 0 12486 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_11
timestamp 1602073617
transform 1 0 12518 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_13
timestamp 1602073617
transform 1 0 12550 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_12
timestamp 1602073617
transform 1 0 12534 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_14
timestamp 1602073617
transform 1 0 12566 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_16
timestamp 1602073617
transform 1 0 12598 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_15
timestamp 1602073617
transform 1 0 12582 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_17
timestamp 1602073617
transform 1 0 12614 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_19
timestamp 1602073617
transform 1 0 12646 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_18
timestamp 1602073617
transform 1 0 12630 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_21
timestamp 1602073617
transform 1 0 12678 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_20
timestamp 1602073617
transform 1 0 12662 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_22
timestamp 1602073617
transform 1 0 12694 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_24
timestamp 1602073617
transform 1 0 12726 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_23
timestamp 1602073617
transform 1 0 12710 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_25
timestamp 1602073617
transform 1 0 12742 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_27
timestamp 1602073617
transform 1 0 12774 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_26
timestamp 1602073617
transform 1 0 12758 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_28
timestamp 1602073617
transform 1 0 12790 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_30
timestamp 1602073617
transform 1 0 12822 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_29
timestamp 1602073617
transform 1 0 12806 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_31
timestamp 1602073617
transform 1 0 12838 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_33
timestamp 1602073617
transform 1 0 12870 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_32
timestamp 1602073617
transform 1 0 12854 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_34
timestamp 1602073617
transform 1 0 12886 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_36
timestamp 1602073617
transform 1 0 12918 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_35
timestamp 1602073617
transform 1 0 12902 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_37
timestamp 1602073617
transform 1 0 12934 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_39
timestamp 1602073617
transform 1 0 12966 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_38
timestamp 1602073617
transform 1 0 12950 0 1 7810
box -4 -6 20 206
use FILL  FILL_40_40
timestamp 1602073617
transform 1 0 12982 0 1 7810
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_478
timestamp 1602073617
transform 1 0 8 0 -1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_469
timestamp 1602073617
transform -1 0 1308 0 -1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_320
timestamp 1602073617
transform 1 0 1308 0 -1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_324
timestamp 1602073617
transform 1 0 1958 0 -1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_321
timestamp 1602073617
transform -1 0 3258 0 -1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_20
timestamp 1602073617
transform 1 0 3258 0 -1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_33
timestamp 1602073617
transform 1 0 3908 0 -1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_35
timestamp 1602073617
transform 1 0 4558 0 -1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_207
timestamp 1602073617
transform -1 0 5858 0 -1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_199
timestamp 1602073617
transform -1 0 6508 0 -1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_195
timestamp 1602073617
transform -1 0 7158 0 -1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_736
timestamp 1602073617
transform 1 0 7158 0 -1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_741
timestamp 1602073617
transform 1 0 7808 0 -1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_177
timestamp 1602073617
transform 1 0 8458 0 -1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_727
timestamp 1602073617
transform 1 0 9108 0 -1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_337
timestamp 1602073617
transform -1 0 10408 0 -1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_91
timestamp 1602073617
transform 1 0 10408 0 -1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_775
timestamp 1602073617
transform 1 0 11058 0 -1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_731
timestamp 1602073617
transform -1 0 12358 0 -1 8210
box -4 -6 618 206
use FILL  FILL_41_1
timestamp 1602073617
transform -1 0 12374 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_2
timestamp 1602073617
transform -1 0 12390 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_3
timestamp 1602073617
transform -1 0 12406 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_4
timestamp 1602073617
transform -1 0 12422 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_5
timestamp 1602073617
transform -1 0 12438 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_6
timestamp 1602073617
transform -1 0 12454 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_7
timestamp 1602073617
transform -1 0 12470 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_8
timestamp 1602073617
transform -1 0 12486 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_10
timestamp 1602073617
transform -1 0 12518 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_9
timestamp 1602073617
transform -1 0 12502 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_11
timestamp 1602073617
transform -1 0 12534 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_13
timestamp 1602073617
transform -1 0 12566 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_12
timestamp 1602073617
transform -1 0 12550 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_14
timestamp 1602073617
transform -1 0 12582 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_16
timestamp 1602073617
transform -1 0 12614 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_15
timestamp 1602073617
transform -1 0 12598 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_17
timestamp 1602073617
transform -1 0 12630 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_19
timestamp 1602073617
transform -1 0 12662 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_18
timestamp 1602073617
transform -1 0 12646 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_21
timestamp 1602073617
transform -1 0 12694 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_20
timestamp 1602073617
transform -1 0 12678 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_22
timestamp 1602073617
transform -1 0 12710 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_24
timestamp 1602073617
transform -1 0 12742 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_23
timestamp 1602073617
transform -1 0 12726 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_25
timestamp 1602073617
transform -1 0 12758 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_27
timestamp 1602073617
transform -1 0 12790 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_26
timestamp 1602073617
transform -1 0 12774 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_28
timestamp 1602073617
transform -1 0 12806 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_30
timestamp 1602073617
transform -1 0 12838 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_29
timestamp 1602073617
transform -1 0 12822 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_31
timestamp 1602073617
transform -1 0 12854 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_33
timestamp 1602073617
transform -1 0 12886 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_32
timestamp 1602073617
transform -1 0 12870 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_34
timestamp 1602073617
transform -1 0 12902 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_36
timestamp 1602073617
transform -1 0 12934 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_35
timestamp 1602073617
transform -1 0 12918 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_37
timestamp 1602073617
transform -1 0 12950 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_39
timestamp 1602073617
transform -1 0 12982 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_38
timestamp 1602073617
transform -1 0 12966 0 -1 8210
box -4 -6 20 206
use FILL  FILL_41_40
timestamp 1602073617
transform -1 0 12998 0 -1 8210
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_863
timestamp 1602073617
transform -1 0 658 0 1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_856
timestamp 1602073617
transform -1 0 1308 0 1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_854
timestamp 1602073617
transform -1 0 1958 0 1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_326
timestamp 1602073617
transform -1 0 2608 0 1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_333
timestamp 1602073617
transform 1 0 2608 0 1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_857
timestamp 1602073617
transform -1 0 3908 0 1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_852
timestamp 1602073617
transform -1 0 4558 0 1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_79
timestamp 1602073617
transform 1 0 4558 0 1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_214
timestamp 1602073617
transform 1 0 5208 0 1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_219
timestamp 1602073617
transform 1 0 5858 0 1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_222
timestamp 1602073617
transform 1 0 6508 0 1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_835
timestamp 1602073617
transform -1 0 7808 0 1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_821
timestamp 1602073617
transform -1 0 8458 0 1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_303
timestamp 1602073617
transform 1 0 8458 0 1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_353
timestamp 1602073617
transform 1 0 9108 0 1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_182
timestamp 1602073617
transform -1 0 10408 0 1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_164
timestamp 1602073617
transform 1 0 10408 0 1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_776
timestamp 1602073617
transform 1 0 11058 0 1 8210
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_785
timestamp 1602073617
transform 1 0 11708 0 1 8210
box -4 -6 618 206
use FILL  FILL_42_1
timestamp 1602073617
transform 1 0 12358 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_2
timestamp 1602073617
transform 1 0 12374 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_3
timestamp 1602073617
transform 1 0 12390 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_4
timestamp 1602073617
transform 1 0 12406 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_5
timestamp 1602073617
transform 1 0 12422 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_6
timestamp 1602073617
transform 1 0 12438 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_7
timestamp 1602073617
transform 1 0 12454 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_8
timestamp 1602073617
transform 1 0 12470 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_10
timestamp 1602073617
transform 1 0 12502 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_9
timestamp 1602073617
transform 1 0 12486 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_11
timestamp 1602073617
transform 1 0 12518 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_13
timestamp 1602073617
transform 1 0 12550 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_12
timestamp 1602073617
transform 1 0 12534 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_14
timestamp 1602073617
transform 1 0 12566 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_16
timestamp 1602073617
transform 1 0 12598 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_15
timestamp 1602073617
transform 1 0 12582 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_17
timestamp 1602073617
transform 1 0 12614 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_19
timestamp 1602073617
transform 1 0 12646 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_18
timestamp 1602073617
transform 1 0 12630 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_21
timestamp 1602073617
transform 1 0 12678 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_20
timestamp 1602073617
transform 1 0 12662 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_22
timestamp 1602073617
transform 1 0 12694 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_24
timestamp 1602073617
transform 1 0 12726 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_23
timestamp 1602073617
transform 1 0 12710 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_25
timestamp 1602073617
transform 1 0 12742 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_27
timestamp 1602073617
transform 1 0 12774 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_26
timestamp 1602073617
transform 1 0 12758 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_28
timestamp 1602073617
transform 1 0 12790 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_30
timestamp 1602073617
transform 1 0 12822 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_29
timestamp 1602073617
transform 1 0 12806 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_31
timestamp 1602073617
transform 1 0 12838 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_33
timestamp 1602073617
transform 1 0 12870 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_32
timestamp 1602073617
transform 1 0 12854 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_34
timestamp 1602073617
transform 1 0 12886 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_36
timestamp 1602073617
transform 1 0 12918 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_35
timestamp 1602073617
transform 1 0 12902 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_37
timestamp 1602073617
transform 1 0 12934 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_39
timestamp 1602073617
transform 1 0 12966 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_38
timestamp 1602073617
transform 1 0 12950 0 1 8210
box -4 -6 20 206
use FILL  FILL_42_40
timestamp 1602073617
transform 1 0 12982 0 1 8210
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_662
timestamp 1602073617
transform 1 0 8 0 -1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_799
timestamp 1602073617
transform -1 0 1308 0 -1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_594
timestamp 1602073617
transform -1 0 1958 0 -1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_431
timestamp 1602073617
transform 1 0 1958 0 -1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_172
timestamp 1602073617
transform -1 0 3258 0 -1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_338
timestamp 1602073617
transform 1 0 3258 0 -1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_351
timestamp 1602073617
transform 1 0 3908 0 -1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_853
timestamp 1602073617
transform -1 0 5208 0 -1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_204
timestamp 1602073617
transform 1 0 5208 0 -1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_663
timestamp 1602073617
transform 1 0 5858 0 -1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_839
timestamp 1602073617
transform -1 0 7158 0 -1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_674
timestamp 1602073617
transform 1 0 7158 0 -1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_675
timestamp 1602073617
transform -1 0 8458 0 -1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_439
timestamp 1602073617
transform -1 0 9108 0 -1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_578
timestamp 1602073617
transform 1 0 9108 0 -1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_580
timestamp 1602073617
transform 1 0 9758 0 -1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_189
timestamp 1602073617
transform 1 0 10408 0 -1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_192
timestamp 1602073617
transform 1 0 11058 0 -1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_738
timestamp 1602073617
transform 1 0 11708 0 -1 8610
box -4 -6 618 206
use FILL  FILL_43_1
timestamp 1602073617
transform -1 0 12374 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_2
timestamp 1602073617
transform -1 0 12390 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_3
timestamp 1602073617
transform -1 0 12406 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_4
timestamp 1602073617
transform -1 0 12422 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_5
timestamp 1602073617
transform -1 0 12438 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_6
timestamp 1602073617
transform -1 0 12454 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_7
timestamp 1602073617
transform -1 0 12470 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_8
timestamp 1602073617
transform -1 0 12486 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_10
timestamp 1602073617
transform -1 0 12518 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_9
timestamp 1602073617
transform -1 0 12502 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_11
timestamp 1602073617
transform -1 0 12534 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_13
timestamp 1602073617
transform -1 0 12566 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_12
timestamp 1602073617
transform -1 0 12550 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_14
timestamp 1602073617
transform -1 0 12582 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_16
timestamp 1602073617
transform -1 0 12614 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_15
timestamp 1602073617
transform -1 0 12598 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_17
timestamp 1602073617
transform -1 0 12630 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_19
timestamp 1602073617
transform -1 0 12662 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_18
timestamp 1602073617
transform -1 0 12646 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_21
timestamp 1602073617
transform -1 0 12694 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_20
timestamp 1602073617
transform -1 0 12678 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_22
timestamp 1602073617
transform -1 0 12710 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_24
timestamp 1602073617
transform -1 0 12742 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_23
timestamp 1602073617
transform -1 0 12726 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_25
timestamp 1602073617
transform -1 0 12758 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_27
timestamp 1602073617
transform -1 0 12790 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_26
timestamp 1602073617
transform -1 0 12774 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_28
timestamp 1602073617
transform -1 0 12806 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_30
timestamp 1602073617
transform -1 0 12838 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_29
timestamp 1602073617
transform -1 0 12822 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_31
timestamp 1602073617
transform -1 0 12854 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_33
timestamp 1602073617
transform -1 0 12886 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_32
timestamp 1602073617
transform -1 0 12870 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_34
timestamp 1602073617
transform -1 0 12902 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_36
timestamp 1602073617
transform -1 0 12934 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_35
timestamp 1602073617
transform -1 0 12918 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_37
timestamp 1602073617
transform -1 0 12950 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_39
timestamp 1602073617
transform -1 0 12982 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_38
timestamp 1602073617
transform -1 0 12966 0 -1 8610
box -4 -6 20 206
use FILL  FILL_43_40
timestamp 1602073617
transform -1 0 12998 0 -1 8610
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_802
timestamp 1602073617
transform -1 0 658 0 1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_798
timestamp 1602073617
transform -1 0 1308 0 1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_436
timestamp 1602073617
transform -1 0 1958 0 1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_434
timestamp 1602073617
transform -1 0 2608 0 1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_174
timestamp 1602073617
transform 1 0 2608 0 1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_173
timestamp 1602073617
transform 1 0 3258 0 1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_175
timestamp 1602073617
transform 1 0 3908 0 1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_208
timestamp 1602073617
transform -1 0 5208 0 1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_215
timestamp 1602073617
transform -1 0 5858 0 1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_205
timestamp 1602073617
transform -1 0 6508 0 1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_203
timestamp 1602073617
transform -1 0 7158 0 1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_72
timestamp 1602073617
transform -1 0 7808 0 1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_568
timestamp 1602073617
transform 1 0 7808 0 1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_566
timestamp 1602073617
transform -1 0 9108 0 1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_211
timestamp 1602073617
transform -1 0 9758 0 1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_170
timestamp 1602073617
transform -1 0 10408 0 1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_168
timestamp 1602073617
transform -1 0 11058 0 1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_739
timestamp 1602073617
transform 1 0 11058 0 1 8610
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_740
timestamp 1602073617
transform 1 0 11708 0 1 8610
box -4 -6 618 206
use FILL  FILL_44_1
timestamp 1602073617
transform 1 0 12358 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_2
timestamp 1602073617
transform 1 0 12374 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_3
timestamp 1602073617
transform 1 0 12390 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_4
timestamp 1602073617
transform 1 0 12406 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_5
timestamp 1602073617
transform 1 0 12422 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_6
timestamp 1602073617
transform 1 0 12438 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_7
timestamp 1602073617
transform 1 0 12454 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_8
timestamp 1602073617
transform 1 0 12470 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_10
timestamp 1602073617
transform 1 0 12502 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_9
timestamp 1602073617
transform 1 0 12486 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_11
timestamp 1602073617
transform 1 0 12518 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_13
timestamp 1602073617
transform 1 0 12550 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_12
timestamp 1602073617
transform 1 0 12534 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_14
timestamp 1602073617
transform 1 0 12566 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_16
timestamp 1602073617
transform 1 0 12598 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_15
timestamp 1602073617
transform 1 0 12582 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_17
timestamp 1602073617
transform 1 0 12614 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_19
timestamp 1602073617
transform 1 0 12646 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_18
timestamp 1602073617
transform 1 0 12630 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_21
timestamp 1602073617
transform 1 0 12678 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_20
timestamp 1602073617
transform 1 0 12662 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_22
timestamp 1602073617
transform 1 0 12694 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_24
timestamp 1602073617
transform 1 0 12726 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_23
timestamp 1602073617
transform 1 0 12710 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_25
timestamp 1602073617
transform 1 0 12742 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_27
timestamp 1602073617
transform 1 0 12774 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_26
timestamp 1602073617
transform 1 0 12758 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_28
timestamp 1602073617
transform 1 0 12790 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_30
timestamp 1602073617
transform 1 0 12822 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_29
timestamp 1602073617
transform 1 0 12806 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_31
timestamp 1602073617
transform 1 0 12838 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_33
timestamp 1602073617
transform 1 0 12870 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_32
timestamp 1602073617
transform 1 0 12854 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_34
timestamp 1602073617
transform 1 0 12886 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_36
timestamp 1602073617
transform 1 0 12918 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_35
timestamp 1602073617
transform 1 0 12902 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_37
timestamp 1602073617
transform 1 0 12934 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_39
timestamp 1602073617
transform 1 0 12966 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_38
timestamp 1602073617
transform 1 0 12950 0 1 8610
box -4 -6 20 206
use FILL  FILL_44_40
timestamp 1602073617
transform 1 0 12982 0 1 8610
box -4 -6 20 206
use SECLIBAND_opt  SECLIBAND_opt_661
timestamp 1602073617
transform -1 0 658 0 -1 9010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_653
timestamp 1602073617
transform -1 0 1308 0 -1 9010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_468
timestamp 1602073617
transform -1 0 1958 0 -1 9010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_652
timestamp 1602073617
transform -1 0 2608 0 -1 9010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_440
timestamp 1602073617
transform -1 0 3258 0 -1 9010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_437
timestamp 1602073617
transform -1 0 3908 0 -1 9010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_354
timestamp 1602073617
transform 1 0 3908 0 -1 9010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_358
timestamp 1602073617
transform 1 0 4558 0 -1 9010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_356
timestamp 1602073617
transform 1 0 5208 0 -1 9010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_365
timestamp 1602073617
transform 1 0 5858 0 -1 9010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_367
timestamp 1602073617
transform 1 0 6508 0 -1 9010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_364
timestamp 1602073617
transform -1 0 7808 0 -1 9010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_357
timestamp 1602073617
transform -1 0 8458 0 -1 9010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_352
timestamp 1602073617
transform -1 0 9108 0 -1 9010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_212
timestamp 1602073617
transform 1 0 9108 0 -1 9010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_220
timestamp 1602073617
transform 1 0 9758 0 -1 9010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_221
timestamp 1602073617
transform 1 0 10408 0 -1 9010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_223
timestamp 1602073617
transform 1 0 11058 0 -1 9010
box -4 -6 618 206
use SECLIBAND_opt  SECLIBAND_opt_742
timestamp 1602073617
transform -1 0 12358 0 -1 9010
box -4 -6 618 206
use FILL  FILL_45_1
timestamp 1602073617
transform -1 0 12374 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_2
timestamp 1602073617
transform -1 0 12390 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_3
timestamp 1602073617
transform -1 0 12406 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_4
timestamp 1602073617
transform -1 0 12422 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_5
timestamp 1602073617
transform -1 0 12438 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_6
timestamp 1602073617
transform -1 0 12454 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_7
timestamp 1602073617
transform -1 0 12470 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_8
timestamp 1602073617
transform -1 0 12486 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_10
timestamp 1602073617
transform -1 0 12518 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_9
timestamp 1602073617
transform -1 0 12502 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_11
timestamp 1602073617
transform -1 0 12534 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_13
timestamp 1602073617
transform -1 0 12566 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_12
timestamp 1602073617
transform -1 0 12550 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_14
timestamp 1602073617
transform -1 0 12582 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_16
timestamp 1602073617
transform -1 0 12614 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_15
timestamp 1602073617
transform -1 0 12598 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_17
timestamp 1602073617
transform -1 0 12630 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_19
timestamp 1602073617
transform -1 0 12662 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_18
timestamp 1602073617
transform -1 0 12646 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_21
timestamp 1602073617
transform -1 0 12694 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_20
timestamp 1602073617
transform -1 0 12678 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_22
timestamp 1602073617
transform -1 0 12710 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_24
timestamp 1602073617
transform -1 0 12742 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_23
timestamp 1602073617
transform -1 0 12726 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_25
timestamp 1602073617
transform -1 0 12758 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_27
timestamp 1602073617
transform -1 0 12790 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_26
timestamp 1602073617
transform -1 0 12774 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_28
timestamp 1602073617
transform -1 0 12806 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_30
timestamp 1602073617
transform -1 0 12838 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_29
timestamp 1602073617
transform -1 0 12822 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_31
timestamp 1602073617
transform -1 0 12854 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_33
timestamp 1602073617
transform -1 0 12886 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_32
timestamp 1602073617
transform -1 0 12870 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_34
timestamp 1602073617
transform -1 0 12902 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_36
timestamp 1602073617
transform -1 0 12934 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_35
timestamp 1602073617
transform -1 0 12918 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_37
timestamp 1602073617
transform -1 0 12950 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_39
timestamp 1602073617
transform -1 0 12982 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_38
timestamp 1602073617
transform -1 0 12966 0 -1 9010
box -4 -6 20 206
use FILL  FILL_45_40
timestamp 1602073617
transform -1 0 12998 0 -1 9010
box -4 -6 20 206
<< labels >>
rlabel metal3 s -48 5120 -48 5120 4 INPUT_0
port 0 nsew
rlabel metal3 s -48 5100 -48 5100 4 D_INPUT_0
port 1 nsew
rlabel metal2 s 7008 -40 7008 -40 8 INPUT_1
port 2 nsew
rlabel metal2 s 7040 -40 7040 -40 8 D_INPUT_1
port 3 nsew
rlabel metal2 s 6000 -40 6000 -40 8 INPUT_2
port 4 nsew
rlabel metal2 s 5968 -40 5968 -40 8 D_INPUT_2
port 5 nsew
rlabel metal2 s 9216 -40 9216 -40 8 INPUT_3
port 6 nsew
rlabel metal2 s 9248 -40 9248 -40 8 D_INPUT_3
port 7 nsew
rlabel metal2 s 1840 -40 1840 -40 8 INPUT_4
port 8 nsew
rlabel metal2 s 1808 -40 1808 -40 8 D_INPUT_4
port 9 nsew
rlabel metal2 s 1760 -40 1760 -40 8 INPUT_5
port 10 nsew
rlabel metal2 s 2752 -40 2752 -40 8 D_INPUT_5
port 11 nsew
rlabel metal2 s 144 -40 144 -40 8 INPUT_6
port 12 nsew
rlabel metal2 s 176 -40 176 -40 8 D_INPUT_6
port 13 nsew
rlabel metal3 s -48 500 -48 500 4 INPUT_7
port 14 nsew
rlabel metal2 s 208 -40 208 -40 8 D_INPUT_7
port 15 nsew
rlabel metal2 s 11632 9080 11632 9080 6 D_GATE_222
port 16 nsew
rlabel metal2 s 7088 9080 7088 9080 6 D_GATE_366
port 17 nsew
rlabel metal3 s -48 7740 -48 7740 4 D_GATE_479
port 18 nsew
rlabel metal2 s 10320 9080 10320 9080 6 D_GATE_579
port 19 nsew
rlabel metal2 s 6416 9080 6416 9080 6 D_GATE_662
port 20 nsew
rlabel metal2 s 11792 9080 11792 9080 6 D_GATE_741
port 21 nsew
rlabel metal3 s -48 5540 -48 5540 4 D_GATE_811
port 22 nsew
rlabel metal3 s -48 4520 -48 4520 4 D_GATE_865
port 23 nsew
rlabel metal2 s 11664 9080 11664 9080 6 GATE_222
port 24 nsew
rlabel metal2 s 7120 9080 7120 9080 6 GATE_366
port 25 nsew
rlabel metal3 s -48 7720 -48 7720 4 GATE_479
port 26 nsew
rlabel metal2 s 10352 9080 10352 9080 6 GATE_579
port 27 nsew
rlabel metal2 s 6448 9080 6448 9080 6 GATE_662
port 28 nsew
rlabel metal2 s 11760 9080 11760 9080 6 GATE_741
port 29 nsew
rlabel metal3 s -48 5520 -48 5520 4 GATE_811
port 30 nsew
rlabel metal3 s -48 4540 -48 4540 4 GATE_865
port 31 nsew
rlabel metal3 s 13072 7220 13072 7220 6 gate
port 32 nsew
rlabel metal3 s -48 1540 -48 1540 4 type:
port 33 nsew
rlabel metal3 s -48 3800 -48 3800 4 dual-rail
port 34 nsew
rlabel metal2 s 7968 9080 7968 9080 6 AND;
port 35 nsew
rlabel metal3 s -48 3540 -48 3540 4 name:
port 36 nsew
rlabel metal2 s 784 -40 784 -40 8 GATE_0
port 37 nsew
<< end >>
