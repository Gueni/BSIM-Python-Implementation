* SPICE3 file created from dualRailAS.ext - technology: scmos
*
* drain/source ordering enforced by hand
*

.subckt NAND2X1_LOC a_36_24# Y VSS VDD A B
X0 a_36_24# A VSS VSS NMOS_MAGIC ad=0.6p pd=4.6u as=1p ps=5u w=2u l=0.2u
X1 Y B a_36_24# VSS NMOS_MAGIC ad=1p pd=5u as=0p ps=0u w=2u l=0.2u
X2 Y B VDD VDD PMOS_MAGIC ad=2p pd=10u as=1.2p ps=5.2u w=2u l=0.2u
X3 Y A VDD VDD PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=2u l=0.2u
C0 B Y 0.10fF
C1 Y a_36_24# 0.01fF
C2 VDD A 0.20fF
C3 VDD B 0.27fF
C4 A B 0.22fF
C5 VDD Y 0.57fF
C6 A Y 0.08fF
C7 Y VSS 0.20fF
C8 B VSS 0.19fF
C9 A VSS 0.30fF
C10 VDD VSS 1.73fF
.ends

.subckt INVX1_LOC Y VSS VDD A
X0 Y A VSS VSS NMOS_MAGIC ad=0.5p pd=3u as=0.5p ps=3u w=1u l=0.2u
X1 Y A VDD VDD PMOS_MAGIC ad=1p pd=5u as=1p ps=5u w=2u l=0.2u

C0 VDD A 0.20fF
C1 VDD Y 0.39fF
C2 A Y 0.08fF
C3 Y VSS 0.07fF
C4 A VSS 0.37fF
C5 VDD VSS 1.52fF
.ends 

.subckt NOR2X1_LOC a_36_216# Y VSS VDD A B
X0 Y B a_36_216# VDD PMOS_MAGIC ad=2p pd=9u as=1.2p ps=8.6u w=4u l=0.2u
X1 Y B VSS VSS NMOS_MAGIC ad=1p pd=6u as=0.6p ps=3.2u w=1u l=0.2u
X2 Y A VSS VSS NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=1u l=0.2u
X3 a_36_216# A VDD VDD PMOS_MAGIC ad=0p pd=0u as=2p ps=9u w=4u l=0.2u

C0 VDD A 0.07fF
C1 VDD B 0.12fF
C2 A B 0.18fF
C3 VDD Y 0.17fF
C4 A Y 0.07fF
C5 B Y 0.12fF
C6 a_36_216# Y 0.01fF
C7 Y VSS 0.11fF
C8 B VSS 0.28fF
C9 A VSS 0.37fF
C10 VDD VSS 1.73fF
.ends

.subckt AES_SBOX INPUT_0 INPUT_1 INPUT_2 INPUT_3 INPUT_4 INPUT_5 INPUT_6 INPUT_7 
+ D_INPUT_0 D_INPUT_1 D_INPUT_2 D_INPUT_3 D_INPUT_4 D_INPUT_5 D_INPUT_6 D_INPUT_7 
+ GATE_222 GATE_366 GATE_479 GATE_579 GATE_662 GATE_741 GATE_811 GATE_865 
+ D_GATE_222 D_GATE_366 D_GATE_479 D_GATE_579 D_GATE_662 D_GATE_741 D_GATE_811 D_GATE_865 
+ VDD VSS 

XNAND2X1_LOC_580 NAND2X1_LOC_580/a_36_24# GATE_579 VSS VDD INVX1_LOC_240/Y INVX1_LOC_242/Y
+ NAND2X1_LOC
XNAND2X1_LOC_591 NAND2X1_LOC_591/a_36_24# NOR2X1_LOC_718/B VSS VDD INVX1_LOC_50/Y
+ NOR2X1_LOC_590/Y NAND2X1_LOC
XNOR2X1_LOC_815 NOR2X1_LOC_815/a_36_216# NOR2X1_LOC_815/Y VSS VDD NOR2X1_LOC_815/A
+ INVX1_LOC_2/A NOR2X1_LOC
XNOR2X1_LOC_804 NOR2X1_LOC_804/a_36_216# NOR2X1_LOC_808/A VSS VDD NOR2X1_LOC_795/Y
+ NOR2X1_LOC_804/B NOR2X1_LOC
XNOR2X1_LOC_826 NOR2X1_LOC_826/a_36_216# NOR2X1_LOC_826/Y VSS VDD INVX1_LOC_58/A INVX1_LOC_42/A
+ NOR2X1_LOC
XNOR2X1_LOC_848 NOR2X1_LOC_848/a_36_216# NOR2X1_LOC_848/Y VSS VDD INVX1_LOC_315/Y
+ NOR2X1_LOC_846/Y NOR2X1_LOC
XNOR2X1_LOC_859 NOR2X1_LOC_859/a_36_216# NOR2X1_LOC_859/Y VSS VDD NOR2X1_LOC_859/A
+ NOR2X1_LOC_848/Y NOR2X1_LOC
XNOR2X1_LOC_837 NOR2X1_LOC_837/a_36_216# NOR2X1_LOC_837/Y VSS VDD NOR2X1_LOC_837/A
+ NOR2X1_LOC_837/B NOR2X1_LOC
XINVX1_LOC_210 INVX1_LOC_210/Y VSS VDD INVX1_LOC_210/A INVX1_LOC
XINVX1_LOC_232 INVX1_LOC_232/Y VSS VDD INVX1_LOC_232/A INVX1_LOC
XINVX1_LOC_221 INVX1_LOC_221/Y VSS VDD INVX1_LOC_221/A INVX1_LOC
XINVX1_LOC_243 INVX1_LOC_243/Y VSS VDD INVX1_LOC_243/A INVX1_LOC
XNAND2X1_LOC_10 NAND2X1_LOC_10/a_36_24# INVX1_LOC_9/A VSS VDD INVX1_LOC_7/A NAND2X1_LOC_9/Y
+ NAND2X1_LOC
XNAND2X1_LOC_32 NAND2X1_LOC_32/a_36_24# NOR2X1_LOC_34/A VSS VDD NOR2X1_LOC_87/B INVX1_LOC_21/A
+ NAND2X1_LOC
XNAND2X1_LOC_43 NAND2X1_LOC_43/a_36_24# NOR2X1_LOC_195/A VSS VDD INVX1_LOC_17/A INVX1_LOC_31/A
+ NAND2X1_LOC
XNAND2X1_LOC_21 NAND2X1_LOC_21/a_36_24# NAND2X1_LOC_21/Y VSS VDD INPUT_4 D_INPUT_5
+ NAND2X1_LOC
XINVX1_LOC_254 INVX1_LOC_254/Y VSS VDD INVX1_LOC_254/A INVX1_LOC
XINVX1_LOC_265 INVX1_LOC_265/Y VSS VDD INVX1_LOC_265/A INVX1_LOC
XINVX1_LOC_276 INVX1_LOC_276/Y VSS VDD INVX1_LOC_276/A INVX1_LOC
XINVX1_LOC_298 INVX1_LOC_298/Y VSS VDD INVX1_LOC_298/A INVX1_LOC
XINVX1_LOC_287 INVX1_LOC_287/Y VSS VDD INVX1_LOC_287/A INVX1_LOC
XNOR2X1_LOC_601 NOR2X1_LOC_601/a_36_216# NOR2X1_LOC_601/Y VSS VDD INVX1_LOC_36/A NOR2X1_LOC_15/Y
+ NOR2X1_LOC
XNOR2X1_LOC_678 NOR2X1_LOC_678/a_36_216# INVX1_LOC_272/A VSS VDD NOR2X1_LOC_678/A
+ INVX1_LOC_12/Y NOR2X1_LOC
XNOR2X1_LOC_667 NOR2X1_LOC_667/a_36_216# NOR2X1_LOC_667/Y VSS VDD NOR2X1_LOC_667/A
+ INVX1_LOC_49/Y NOR2X1_LOC
XNOR2X1_LOC_645 NOR2X1_LOC_645/a_36_216# INVX1_LOC_264/A VSS VDD INVX1_LOC_250/A INVX1_LOC_248/A
+ NOR2X1_LOC
XNOR2X1_LOC_634 NOR2X1_LOC_634/a_36_216# NOR2X1_LOC_634/Y VSS VDD NOR2X1_LOC_634/A
+ NOR2X1_LOC_634/B NOR2X1_LOC
XNAND2X1_LOC_54 NAND2X1_LOC_54/a_36_24# INVX1_LOC_39/A VSS VDD INPUT_0 INPUT_1
+ NAND2X1_LOC
XNAND2X1_LOC_65 NAND2X1_LOC_65/a_36_24# NOR2X1_LOC_201/A VSS VDD NAND2X1_LOC_63/Y
+ INVX1_LOC_50/Y NAND2X1_LOC
XNAND2X1_LOC_87 NAND2X1_LOC_87/a_36_24# NOR2X1_LOC_88/A VSS VDD NOR2X1_LOC_32/B NOR2X1_LOC_52/B
+ NAND2X1_LOC
XNAND2X1_LOC_98 NAND2X1_LOC_98/a_36_24# INVX1_LOC_59/A VSS VDD NOR2X1_LOC_93/Y NOR2X1_LOC_96/Y
+ NAND2X1_LOC
XNAND2X1_LOC_76 NAND2X1_LOC_76/a_36_24# INVX1_LOC_55/A VSS VDD NOR2X1_LOC_74/Y NOR2X1_LOC_75/Y
+ NAND2X1_LOC
XNOR2X1_LOC_656 NOR2X1_LOC_656/a_36_216# NOR2X1_LOC_656/Y VSS VDD NOR2X1_LOC_647/Y
+ NOR2X1_LOC_216/B NOR2X1_LOC
XNOR2X1_LOC_623 NOR2X1_LOC_623/a_36_216# NOR2X1_LOC_624/A VSS VDD NOR2X1_LOC_620/Y
+ NOR2X1_LOC_623/B NOR2X1_LOC
XNOR2X1_LOC_612 NOR2X1_LOC_612/a_36_216# NOR2X1_LOC_612/Y VSS VDD INVX1_LOC_251/Y
+ NOR2X1_LOC_612/B NOR2X1_LOC
XNOR2X1_LOC_689 NOR2X1_LOC_689/a_36_216# NOR2X1_LOC_689/Y VSS VDD NOR2X1_LOC_689/A
+ INVX1_LOC_22/A NOR2X1_LOC
XNAND2X1_LOC_409 NAND2X1_LOC_409/a_36_24# NOR2X1_LOC_460/A VSS VDD NOR2X1_LOC_828/B
+ INVX1_LOC_174/Y NAND2X1_LOC
XNOR2X1_LOC_453 NOR2X1_LOC_453/a_36_216# NOR2X1_LOC_453/Y VSS VDD INVX1_LOC_189/Y
+ NOR2X1_LOC_448/Y NOR2X1_LOC
XNOR2X1_LOC_486 NOR2X1_LOC_486/a_36_216# NOR2X1_LOC_486/Y VSS VDD NOR2X1_LOC_705/B
+ NOR2X1_LOC_486/B NOR2X1_LOC
XNOR2X1_LOC_431 NOR2X1_LOC_431/a_36_216# NOR2X1_LOC_431/Y VSS VDD INVX1_LOC_118/A
+ INVX1_LOC_54/A NOR2X1_LOC
XNOR2X1_LOC_464 NOR2X1_LOC_464/a_36_216# NOR2X1_LOC_464/Y VSS VDD NOR2X1_LOC_458/Y
+ NOR2X1_LOC_464/B NOR2X1_LOC
XNOR2X1_LOC_475 NOR2X1_LOC_475/a_36_216# NOR2X1_LOC_479/B VSS VDD NOR2X1_LOC_475/A
+ INVX1_LOC_172/Y NOR2X1_LOC
XNOR2X1_LOC_497 NOR2X1_LOC_497/a_36_216# NOR2X1_LOC_497/Y VSS VDD NOR2X1_LOC_71/Y
+ INVX1_LOC_17/Y NOR2X1_LOC
XNOR2X1_LOC_420 NOR2X1_LOC_420/a_36_216# NOR2X1_LOC_420/Y VSS VDD NOR2X1_LOC_536/A
+ INVX1_LOC_58/A NOR2X1_LOC
XNOR2X1_LOC_442 NOR2X1_LOC_442/a_36_216# INVX1_LOC_184/A VSS VDD INVX1_LOC_64/A INVX1_LOC_30/A
+ NOR2X1_LOC
XNAND2X1_LOC_206 NAND2X1_LOC_206/a_36_24# NAND2X1_LOC_206/Y VSS VDD INVX1_LOC_110/Y
+ NAND2X1_LOC_206/B NAND2X1_LOC
XNAND2X1_LOC_217 NAND2X1_LOC_217/a_36_24# NAND2X1_LOC_218/B VSS VDD INVX1_LOC_74/Y
+ NAND2X1_LOC_141/Y NAND2X1_LOC
XNAND2X1_LOC_239 NAND2X1_LOC_239/a_36_24# INVX1_LOC_119/A VSS VDD INVX1_LOC_37/A NOR2X1_LOC_590/A
+ NAND2X1_LOC
XNAND2X1_LOC_228 NAND2X1_LOC_228/a_36_24# NAND2X1_LOC_341/A VSS VDD NOR2X1_LOC_7/Y
+ NOR2X1_LOC_52/Y NAND2X1_LOC
XNOR2X1_LOC_261 NOR2X1_LOC_261/a_36_216# NOR2X1_LOC_261/Y VSS VDD NOR2X1_LOC_261/A
+ INVX1_LOC_63/Y NOR2X1_LOC
XNOR2X1_LOC_272 NOR2X1_LOC_272/a_36_216# NOR2X1_LOC_272/Y VSS VDD INVX1_LOC_32/A INVX1_LOC_22/A
+ NOR2X1_LOC
XNOR2X1_LOC_250 NOR2X1_LOC_250/a_36_216# NOR2X1_LOC_250/Y VSS VDD NOR2X1_LOC_250/A
+ INVX1_LOC_49/Y NOR2X1_LOC
XNOR2X1_LOC_294 NOR2X1_LOC_294/a_36_216# NOR2X1_LOC_294/Y VSS VDD INVX1_LOC_135/A
+ INVX1_LOC_9/A NOR2X1_LOC
XNOR2X1_LOC_283 NOR2X1_LOC_283/a_36_216# INVX1_LOC_132/A VSS VDD NOR2X1_LOC_226/A
+ INVX1_LOC_20/A NOR2X1_LOC
XNAND2X1_LOC_795 NAND2X1_LOC_795/a_36_24# NAND2X1_LOC_795/Y VSS VDD NAND2X1_LOC_785/Y
+ INVX1_LOC_304/Y NAND2X1_LOC
XNAND2X1_LOC_773 NAND2X1_LOC_773/a_36_24# NAND2X1_LOC_773/Y VSS VDD INVX1_LOC_293/Y
+ NAND2X1_LOC_773/B NAND2X1_LOC
XNAND2X1_LOC_751 NAND2X1_LOC_751/a_36_24# NOR2X1_LOC_789/A VSS VDD INVX1_LOC_2/Y NOR2X1_LOC_750/Y
+ NAND2X1_LOC
XNAND2X1_LOC_784 NAND2X1_LOC_784/a_36_24# NAND2X1_LOC_796/B VSS VDD NAND2X1_LOC_784/A
+ NAND2X1_LOC_778/Y NAND2X1_LOC
XNAND2X1_LOC_740 NAND2X1_LOC_740/a_36_24# NAND2X1_LOC_740/Y VSS VDD NAND2X1_LOC_740/A
+ NAND2X1_LOC_740/B NAND2X1_LOC
XNAND2X1_LOC_762 NAND2X1_LOC_762/a_36_24# NAND2X1_LOC_763/B VSS VDD INPUT_6 NAND2X1_LOC_11/Y
+ NAND2X1_LOC
XINVX1_LOC_6 INVX1_LOC_6/Y VSS VDD INVX1_LOC_6/A INVX1_LOC
XNAND2X1_LOC_570 NAND2X1_LOC_570/a_36_24# NAND2X1_LOC_570/Y VSS VDD NAND2X1_LOC_562/Y
+ NAND2X1_LOC_563/Y NAND2X1_LOC
XNAND2X1_LOC_592 NAND2X1_LOC_592/a_36_24# INVX1_LOC_245/A VSS VDD NOR2X1_LOC_423/Y
+ NOR2X1_LOC_589/Y NAND2X1_LOC
XNAND2X1_LOC_581 NAND2X1_LOC_581/a_36_24# NAND2X1_LOC_581/Y VSS VDD INPUT_6 NAND2X1_LOC_3/B
+ NAND2X1_LOC
XNOR2X1_LOC_816 NOR2X1_LOC_816/a_36_216# NOR2X1_LOC_816/Y VSS VDD NOR2X1_LOC_816/A
+ INVX1_LOC_38/A NOR2X1_LOC
XNOR2X1_LOC_805 NOR2X1_LOC_805/a_36_216# NOR2X1_LOC_807/B VSS VDD NOR2X1_LOC_793/Y
+ INVX1_LOC_307/Y NOR2X1_LOC
XNOR2X1_LOC_849 NOR2X1_LOC_849/a_36_216# NOR2X1_LOC_859/A VSS VDD NOR2X1_LOC_849/A
+ NOR2X1_LOC_844/Y NOR2X1_LOC
XNOR2X1_LOC_838 NOR2X1_LOC_838/a_36_216# NOR2X1_LOC_852/B VSS VDD NOR2X1_LOC_837/Y
+ INVX1_LOC_310/Y NOR2X1_LOC
XNOR2X1_LOC_827 NOR2X1_LOC_827/a_36_216# INVX1_LOC_310/A VSS VDD INVX1_LOC_90/A INVX1_LOC_31/Y
+ NOR2X1_LOC
XINVX1_LOC_255 INVX1_LOC_255/Y VSS VDD INVX1_LOC_255/A INVX1_LOC
XINVX1_LOC_200 INVX1_LOC_200/Y VSS VDD INVX1_LOC_200/A INVX1_LOC
XINVX1_LOC_233 INVX1_LOC_233/Y VSS VDD INVX1_LOC_233/A INVX1_LOC
XINVX1_LOC_222 INVX1_LOC_222/Y VSS VDD INVX1_LOC_222/A INVX1_LOC
XINVX1_LOC_266 INVX1_LOC_266/Y VSS VDD INVX1_LOC_266/A INVX1_LOC
XINVX1_LOC_211 INVX1_LOC_211/Y VSS VDD INVX1_LOC_211/A INVX1_LOC
XINVX1_LOC_277 INVX1_LOC_277/Y VSS VDD INVX1_LOC_277/A INVX1_LOC
XINVX1_LOC_244 INVX1_LOC_244/Y VSS VDD INVX1_LOC_244/A INVX1_LOC
XNAND2X1_LOC_55 NAND2X1_LOC_55/a_36_24# INVX1_LOC_41/A VSS VDD INVX1_LOC_3/A INVX1_LOC_39/A
+ NAND2X1_LOC
XNAND2X1_LOC_66 NAND2X1_LOC_66/a_36_24# NOR2X1_LOC_67/A VSS VDD INVX1_LOC_2/A INVX1_LOC_20/A
+ NAND2X1_LOC
XNAND2X1_LOC_77 NAND2X1_LOC_77/a_36_24# NOR2X1_LOC_78/A VSS VDD INVX1_LOC_13/A INVX1_LOC_39/A
+ NAND2X1_LOC
XNAND2X1_LOC_33 NAND2X1_LOC_33/a_36_24# NAND2X1_LOC_33/Y VSS VDD NOR2X1_LOC_20/Y NOR2X1_LOC_24/Y
+ NAND2X1_LOC
XNAND2X1_LOC_44 NAND2X1_LOC_44/a_36_24# INVX1_LOC_33/A VSS VDD NAND2X1_LOC_36/A NAND2X1_LOC_30/Y
+ NAND2X1_LOC
XNAND2X1_LOC_22 NAND2X1_LOC_22/a_36_24# INVX1_LOC_17/A VSS VDD NAND2X1_LOC_1/Y NAND2X1_LOC_21/Y
+ NAND2X1_LOC
XNAND2X1_LOC_11 NAND2X1_LOC_11/a_36_24# NAND2X1_LOC_11/Y VSS VDD D_INPUT_4 INPUT_5
+ NAND2X1_LOC
XINVX1_LOC_299 INVX1_LOC_299/Y VSS VDD INVX1_LOC_299/A INVX1_LOC
XINVX1_LOC_288 INVX1_LOC_288/Y VSS VDD INVX1_LOC_288/A INVX1_LOC
XNOR2X1_LOC_635 NOR2X1_LOC_635/a_36_216# NOR2X1_LOC_639/B VSS VDD NOR2X1_LOC_635/A
+ NOR2X1_LOC_635/B NOR2X1_LOC
XNOR2X1_LOC_657 NOR2X1_LOC_657/a_36_216# NOR2X1_LOC_657/Y VSS VDD NOR2X1_LOC_510/Y
+ NOR2X1_LOC_657/B NOR2X1_LOC
XNOR2X1_LOC_679 NOR2X1_LOC_679/a_36_216# NOR2X1_LOC_679/Y VSS VDD INVX1_LOC_272/Y
+ NOR2X1_LOC_679/B NOR2X1_LOC
XNOR2X1_LOC_602 NOR2X1_LOC_602/a_36_216# INVX1_LOC_248/A VSS VDD NOR2X1_LOC_602/A
+ NOR2X1_LOC_602/B NOR2X1_LOC
XNAND2X1_LOC_99 NAND2X1_LOC_99/a_36_24# NAND2X1_LOC_99/Y VSS VDD NAND2X1_LOC_99/A
+ INVX1_LOC_60/Y NAND2X1_LOC
XNAND2X1_LOC_88 NAND2X1_LOC_88/a_36_24# NOR2X1_LOC_100/A VSS VDD INVX1_LOC_2/Y NOR2X1_LOC_87/Y
+ NAND2X1_LOC
XNOR2X1_LOC_646 NOR2X1_LOC_646/a_36_216# NOR2X1_LOC_647/A VSS VDD NOR2X1_LOC_646/A
+ NOR2X1_LOC_646/B NOR2X1_LOC
XNOR2X1_LOC_668 NOR2X1_LOC_668/a_36_216# NOR2X1_LOC_668/Y VSS VDD INVX1_LOC_89/A INVX1_LOC_19/A
+ NOR2X1_LOC
XNOR2X1_LOC_613 NOR2X1_LOC_613/a_36_216# NOR2X1_LOC_613/Y VSS VDD INVX1_LOC_42/A INVX1_LOC_30/A
+ NOR2X1_LOC
XNOR2X1_LOC_624 NOR2X1_LOC_624/a_36_216# INVX1_LOC_256/A VSS VDD NOR2X1_LOC_624/A
+ NOR2X1_LOC_624/B NOR2X1_LOC
XNOR2X1_LOC_410 NOR2X1_LOC_410/a_36_216# NOR2X1_LOC_410/Y VSS VDD INVX1_LOC_37/A INVX1_LOC_11/A
+ NOR2X1_LOC
XNOR2X1_LOC_454 NOR2X1_LOC_454/a_36_216# NOR2X1_LOC_454/Y VSS VDD NOR2X1_LOC_447/Y
+ INVX1_LOC_187/Y NOR2X1_LOC
XNOR2X1_LOC_432 NOR2X1_LOC_432/a_36_216# NOR2X1_LOC_432/Y VSS VDD NOR2X1_LOC_589/A
+ INVX1_LOC_16/A NOR2X1_LOC
XNOR2X1_LOC_421 NOR2X1_LOC_421/a_36_216# NOR2X1_LOC_421/Y VSS VDD NOR2X1_LOC_328/Y
+ NOR2X1_LOC_91/A NOR2X1_LOC
XNOR2X1_LOC_465 NOR2X1_LOC_465/a_36_216# NOR2X1_LOC_465/Y VSS VDD NOR2X1_LOC_456/Y
+ NOR2X1_LOC_455/Y NOR2X1_LOC
XNOR2X1_LOC_476 NOR2X1_LOC_476/a_36_216# NOR2X1_LOC_476/Y VSS VDD INVX1_LOC_201/Y
+ NOR2X1_LOC_476/B NOR2X1_LOC
XNOR2X1_LOC_443 NOR2X1_LOC_443/a_36_216# NOR2X1_LOC_443/Y VSS VDD NOR2X1_LOC_545/B
+ NOR2X1_LOC_97/A NOR2X1_LOC
XNOR2X1_LOC_487 NOR2X1_LOC_487/a_36_216# NOR2X1_LOC_487/Y VSS VDD INVX1_LOC_57/Y NOR2X1_LOC_45/B
+ NOR2X1_LOC
XNOR2X1_LOC_498 NOR2X1_LOC_498/a_36_216# NOR2X1_LOC_498/Y VSS VDD NOR2X1_LOC_189/A
+ INVX1_LOC_54/A NOR2X1_LOC
XNAND2X1_LOC_229 NAND2X1_LOC_229/a_36_24# NOR2X1_LOC_231/B VSS VDD INVX1_LOC_11/A
+ NOR2X1_LOC_160/B NAND2X1_LOC
XNAND2X1_LOC_218 NAND2X1_LOC_218/a_36_24# NAND2X1_LOC_222/A VSS VDD NAND2X1_LOC_218/A
+ NAND2X1_LOC_218/B NAND2X1_LOC
XNAND2X1_LOC_207 NAND2X1_LOC_207/a_36_24# NAND2X1_LOC_207/Y VSS VDD INVX1_LOC_108/Y
+ NAND2X1_LOC_207/B NAND2X1_LOC
XNOR2X1_LOC_251 NOR2X1_LOC_251/a_36_216# NOR2X1_LOC_251/Y VSS VDD NOR2X1_LOC_106/A
+ INVX1_LOC_38/A NOR2X1_LOC
XNOR2X1_LOC_240 NOR2X1_LOC_240/a_36_216# NOR2X1_LOC_240/Y VSS VDD NOR2X1_LOC_240/A
+ NOR2X1_LOC_240/B NOR2X1_LOC
XNOR2X1_LOC_273 NOR2X1_LOC_273/a_36_216# NOR2X1_LOC_273/Y VSS VDD NOR2X1_LOC_433/A
+ INVX1_LOC_24/A NOR2X1_LOC
XNOR2X1_LOC_295 NOR2X1_LOC_295/a_36_216# NOR2X1_LOC_295/Y VSS VDD NOR2X1_LOC_481/A
+ INVX1_LOC_45/Y NOR2X1_LOC
XNOR2X1_LOC_284 NOR2X1_LOC_284/a_36_216# NOR2X1_LOC_287/A VSS VDD NOR2X1_LOC_542/B
+ NOR2X1_LOC_284/B NOR2X1_LOC
XNOR2X1_LOC_262 NOR2X1_LOC_262/a_36_216# NOR2X1_LOC_262/Y VSS VDD NOR2X1_LOC_65/B
+ INVX1_LOC_29/Y NOR2X1_LOC
XNAND2X1_LOC_785 NAND2X1_LOC_785/a_36_24# NAND2X1_LOC_785/Y VSS VDD NAND2X1_LOC_785/A
+ NAND2X1_LOC_785/B NAND2X1_LOC
XNAND2X1_LOC_774 NAND2X1_LOC_774/a_36_24# INVX1_LOC_299/A VSS VDD INVX1_LOC_298/Y
+ NAND2X1_LOC_773/Y NAND2X1_LOC
XNAND2X1_LOC_796 NAND2X1_LOC_796/a_36_24# NAND2X1_LOC_796/Y VSS VDD NAND2X1_LOC_783/Y
+ NAND2X1_LOC_796/B NAND2X1_LOC
XNAND2X1_LOC_730 NAND2X1_LOC_730/a_36_24# NAND2X1_LOC_739/B VSS VDD NAND2X1_LOC_728/Y
+ NAND2X1_LOC_729/Y NAND2X1_LOC
XNAND2X1_LOC_741 NAND2X1_LOC_741/a_36_24# NAND2X1_LOC_741/Y VSS VDD NAND2X1_LOC_736/Y
+ NAND2X1_LOC_741/B NAND2X1_LOC
XNAND2X1_LOC_752 NAND2X1_LOC_752/a_36_24# INVX1_LOC_289/A VSS VDD INPUT_5 NAND2X1_LOC_51/B
+ NAND2X1_LOC
XNAND2X1_LOC_763 NAND2X1_LOC_763/a_36_24# NOR2X1_LOC_769/B VSS VDD NOR2X1_LOC_598/B
+ NAND2X1_LOC_763/B NAND2X1_LOC
XINVX1_LOC_7 INVX1_LOC_7/Y VSS VDD INVX1_LOC_7/A INVX1_LOC
XNAND2X1_LOC_560 NAND2X1_LOC_560/a_36_24# INVX1_LOC_229/A VSS VDD NAND2X1_LOC_560/A
+ NAND2X1_LOC_559/Y NAND2X1_LOC
XNAND2X1_LOC_571 NAND2X1_LOC_571/a_36_24# NAND2X1_LOC_571/Y VSS VDD INVX1_LOC_230/Y
+ NAND2X1_LOC_571/B NAND2X1_LOC
XNAND2X1_LOC_593 NAND2X1_LOC_593/a_36_24# NAND2X1_LOC_593/Y VSS VDD NOR2X1_LOC_591/Y
+ INVX1_LOC_246/Y NAND2X1_LOC
XNAND2X1_LOC_582 NAND2X1_LOC_582/a_36_24# NOR2X1_LOC_635/A VSS VDD INVX1_LOC_77/A
+ NAND2X1_LOC_581/Y NAND2X1_LOC
XNAND2X1_LOC_390 NAND2X1_LOC_390/a_36_24# NAND2X1_LOC_392/A VSS VDD NAND2X1_LOC_390/A
+ INVX1_LOC_162/Y NAND2X1_LOC
XNOR2X1_LOC_828 NOR2X1_LOC_828/a_36_216# NOR2X1_LOC_828/Y VSS VDD NOR2X1_LOC_828/A
+ NOR2X1_LOC_828/B NOR2X1_LOC
XNOR2X1_LOC_806 NOR2X1_LOC_806/a_36_216# NOR2X1_LOC_806/Y VSS VDD INVX1_LOC_269/Y
+ INVX1_LOC_134/A NOR2X1_LOC
XNOR2X1_LOC_817 NOR2X1_LOC_817/a_36_216# NOR2X1_LOC_817/Y VSS VDD NOR2X1_LOC_381/Y
+ INPUT_1 NOR2X1_LOC
XNOR2X1_LOC_839 NOR2X1_LOC_839/a_36_216# NOR2X1_LOC_852/A VSS VDD NOR2X1_LOC_836/Y
+ NOR2X1_LOC_839/B NOR2X1_LOC
XINVX1_LOC_212 INVX1_LOC_212/Y VSS VDD INVX1_LOC_212/A INVX1_LOC
XINVX1_LOC_201 INVX1_LOC_201/Y VSS VDD INVX1_LOC_201/A INVX1_LOC
XINVX1_LOC_267 INVX1_LOC_267/Y VSS VDD INVX1_LOC_267/A INVX1_LOC
XINVX1_LOC_234 INVX1_LOC_234/Y VSS VDD INVX1_LOC_234/A INVX1_LOC
XINVX1_LOC_256 INVX1_LOC_256/Y VSS VDD INVX1_LOC_256/A INVX1_LOC
XINVX1_LOC_278 INVX1_LOC_278/Y VSS VDD INVX1_LOC_278/A INVX1_LOC
XINVX1_LOC_223 INVX1_LOC_223/Y VSS VDD INVX1_LOC_223/A INVX1_LOC
XINVX1_LOC_289 INVX1_LOC_289/Y VSS VDD INVX1_LOC_289/A INVX1_LOC
XINVX1_LOC_245 INVX1_LOC_245/Y VSS VDD INVX1_LOC_245/A INVX1_LOC
XNAND2X1_LOC_89 NAND2X1_LOC_89/a_36_24# NOR2X1_LOC_97/B VSS VDD INVX1_LOC_45/A NOR2X1_LOC_78/A
+ NAND2X1_LOC
XNAND2X1_LOC_45 NAND2X1_LOC_45/a_36_24# NAND2X1_LOC_45/Y VSS VDD NOR2X1_LOC_160/B
+ INVX1_LOC_33/A NAND2X1_LOC
XNAND2X1_LOC_34 NAND2X1_LOC_34/a_36_24# NAND2X1_LOC_35/B VSS VDD NOR2X1_LOC_27/Y NOR2X1_LOC_32/Y
+ NAND2X1_LOC
XNAND2X1_LOC_23 NAND2X1_LOC_23/a_36_24# NOR2X1_LOC_160/B VSS VDD NOR2X1_LOC_19/B INVX1_LOC_13/A
+ NAND2X1_LOC
XNAND2X1_LOC_78 NAND2X1_LOC_78/a_36_24# NOR2X1_LOC_79/A VSS VDD NOR2X1_LOC_15/Y NOR2X1_LOC_89/A
+ NAND2X1_LOC
XNAND2X1_LOC_67 NAND2X1_LOC_67/a_36_24# NAND2X1_LOC_67/Y VSS VDD INVX1_LOC_42/Y NOR2X1_LOC_66/Y
+ NAND2X1_LOC
XNAND2X1_LOC_56 NAND2X1_LOC_56/a_36_24# NOR2X1_LOC_197/A VSS VDD NAND2X1_LOC_53/Y
+ INVX1_LOC_41/A NAND2X1_LOC
XNAND2X1_LOC_12 NAND2X1_LOC_12/a_36_24# INVX1_LOC_11/A VSS VDD NAND2X1_LOC_1/Y NAND2X1_LOC_11/Y
+ NAND2X1_LOC
XNOR2X1_LOC_636 NOR2X1_LOC_636/a_36_216# INVX1_LOC_262/A VSS VDD NOR2X1_LOC_636/A
+ NOR2X1_LOC_636/B NOR2X1_LOC
XNOR2X1_LOC_603 NOR2X1_LOC_603/a_36_216# NOR2X1_LOC_603/Y VSS VDD NOR2X1_LOC_52/B
+ INVX1_LOC_12/A NOR2X1_LOC
XNOR2X1_LOC_658 NOR2X1_LOC_658/a_36_216# NOR2X1_LOC_658/Y VSS VDD NOR2X1_LOC_632/Y
+ INVX1_LOC_256/A NOR2X1_LOC
XNOR2X1_LOC_614 NOR2X1_LOC_614/a_36_216# NOR2X1_LOC_614/Y VSS VDD INVX1_LOC_77/A NOR2X1_LOC_78/A
+ NOR2X1_LOC
XNOR2X1_LOC_669 NOR2X1_LOC_669/a_36_216# NOR2X1_LOC_669/Y VSS VDD NOR2X1_LOC_669/A
+ INVX1_LOC_92/A NOR2X1_LOC
XNOR2X1_LOC_647 NOR2X1_LOC_647/a_36_216# NOR2X1_LOC_647/Y VSS VDD NOR2X1_LOC_647/A
+ NOR2X1_LOC_647/B NOR2X1_LOC
XNOR2X1_LOC_625 NOR2X1_LOC_625/a_36_216# NOR2X1_LOC_625/Y VSS VDD INVX1_LOC_136/A
+ NOR2X1_LOC_67/A NOR2X1_LOC
XNOR2X1_LOC_433 NOR2X1_LOC_433/a_36_216# NOR2X1_LOC_433/Y VSS VDD NOR2X1_LOC_433/A
+ INVX1_LOC_54/A NOR2X1_LOC
XNOR2X1_LOC_422 NOR2X1_LOC_422/a_36_216# NOR2X1_LOC_422/Y VSS VDD NOR2X1_LOC_92/Y
+ INVX1_LOC_12/A NOR2X1_LOC
XNOR2X1_LOC_400 NOR2X1_LOC_400/a_36_216# INVX1_LOC_166/A VSS VDD NOR2X1_LOC_400/A
+ NOR2X1_LOC_400/B NOR2X1_LOC
XNOR2X1_LOC_411 NOR2X1_LOC_411/a_36_216# NOR2X1_LOC_411/Y VSS VDD NOR2X1_LOC_411/A
+ INVX1_LOC_64/A NOR2X1_LOC
XNOR2X1_LOC_466 NOR2X1_LOC_466/a_36_216# NOR2X1_LOC_470/B VSS VDD NOR2X1_LOC_454/Y
+ NOR2X1_LOC_453/Y NOR2X1_LOC
XNOR2X1_LOC_477 NOR2X1_LOC_477/a_36_216# NOR2X1_LOC_478/A VSS VDD NOR2X1_LOC_471/Y
+ NOR2X1_LOC_477/B NOR2X1_LOC
XNOR2X1_LOC_499 NOR2X1_LOC_499/a_36_216# NOR2X1_LOC_500/A VSS VDD NOR2X1_LOC_778/A
+ NOR2X1_LOC_499/B NOR2X1_LOC
XNOR2X1_LOC_455 NOR2X1_LOC_455/a_36_216# NOR2X1_LOC_455/Y VSS VDD NOR2X1_LOC_445/Y
+ INVX1_LOC_55/Y NOR2X1_LOC
XNOR2X1_LOC_488 NOR2X1_LOC_488/a_36_216# NOR2X1_LOC_488/Y VSS VDD NOR2X1_LOC_226/A
+ INVX1_LOC_90/A NOR2X1_LOC
XNOR2X1_LOC_444 NOR2X1_LOC_444/a_36_216# INVX1_LOC_186/A VSS VDD NOR2X1_LOC_443/Y
+ INVX1_LOC_184/Y NOR2X1_LOC
XNAND2X1_LOC_208 NAND2X1_LOC_208/a_36_24# NAND2X1_LOC_214/B VSS VDD NAND2X1_LOC_35/Y
+ NAND2X1_LOC_208/B NAND2X1_LOC
XNAND2X1_LOC_219 NAND2X1_LOC_219/a_36_24# NAND2X1_LOC_222/B VSS VDD NAND2X1_LOC_214/Y
+ NAND2X1_LOC_219/B NAND2X1_LOC
XNOR2X1_LOC_230 NOR2X1_LOC_230/a_36_216# NOR2X1_LOC_230/Y VSS VDD INVX1_LOC_22/A INVX1_LOC_6/A
+ NOR2X1_LOC
XNOR2X1_LOC_274 NOR2X1_LOC_274/a_36_216# NOR2X1_LOC_274/Y VSS VDD NOR2X1_LOC_831/B
+ NOR2X1_LOC_274/B NOR2X1_LOC
XNOR2X1_LOC_263 NOR2X1_LOC_263/a_36_216# INVX1_LOC_124/A VSS VDD INVX1_LOC_25/Y INVX1_LOC_18/A
+ NOR2X1_LOC
XNOR2X1_LOC_252 NOR2X1_LOC_252/a_36_216# NOR2X1_LOC_252/Y VSS VDD INVX1_LOC_46/A INVX1_LOC_42/A
+ NOR2X1_LOC
XNOR2X1_LOC_285 NOR2X1_LOC_285/a_36_216# NOR2X1_LOC_285/Y VSS VDD NOR2X1_LOC_285/A
+ NOR2X1_LOC_285/B NOR2X1_LOC
XNOR2X1_LOC_241 NOR2X1_LOC_241/a_36_216# NOR2X1_LOC_242/A VSS VDD NOR2X1_LOC_241/A
+ NOR2X1_LOC_445/B NOR2X1_LOC
XNOR2X1_LOC_296 NOR2X1_LOC_296/a_36_216# NOR2X1_LOC_296/Y VSS VDD INVX1_LOC_41/A INVX1_LOC_31/A
+ NOR2X1_LOC
XNAND2X1_LOC_720 NAND2X1_LOC_720/a_36_24# NAND2X1_LOC_721/B VSS VDD NOR2X1_LOC_667/Y
+ NOR2X1_LOC_669/Y NAND2X1_LOC
XNAND2X1_LOC_786 NAND2X1_LOC_786/a_36_24# INVX1_LOC_303/A VSS VDD NAND2X1_LOC_84/Y
+ NOR2X1_LOC_262/Y NAND2X1_LOC
XNAND2X1_LOC_775 NAND2X1_LOC_775/a_36_24# NAND2X1_LOC_785/A VSS VDD NOR2X1_LOC_91/Y
+ NOR2X1_LOC_109/Y NAND2X1_LOC
XNAND2X1_LOC_731 NAND2X1_LOC_731/a_36_24# NAND2X1_LOC_731/Y VSS VDD NAND2X1_LOC_726/Y
+ NAND2X1_LOC_727/Y NAND2X1_LOC
XNAND2X1_LOC_753 NAND2X1_LOC_753/a_36_24# NOR2X1_LOC_790/B VSS VDD NOR2X1_LOC_188/A
+ INVX1_LOC_290/Y NAND2X1_LOC
XNAND2X1_LOC_742 NAND2X1_LOC_742/a_36_24# GATE_741 VSS VDD NAND2X1_LOC_740/Y NAND2X1_LOC_741/Y
+ NAND2X1_LOC
XNAND2X1_LOC_797 NAND2X1_LOC_797/a_36_24# NAND2X1_LOC_803/B VSS VDD NAND2X1_LOC_149/Y
+ INVX1_LOC_302/Y NAND2X1_LOC
XNAND2X1_LOC_764 NAND2X1_LOC_764/a_36_24# NOR2X1_LOC_769/A VSS VDD INVX1_LOC_29/A
+ INVX1_LOC_75/A NAND2X1_LOC
XINVX1_LOC_8 INVX1_LOC_8/Y VSS VDD INVX1_LOC_8/A INVX1_LOC
XNAND2X1_LOC_572 NAND2X1_LOC_572/a_36_24# INVX1_LOC_233/A VSS VDD INVX1_LOC_73/A NAND2X1_LOC_572/B
+ NAND2X1_LOC
XNAND2X1_LOC_550 NAND2X1_LOC_550/a_36_24# NAND2X1_LOC_565/B VSS VDD NAND2X1_LOC_550/A
+ INVX1_LOC_226/Y NAND2X1_LOC
XNAND2X1_LOC_561 NAND2X1_LOC_561/a_36_24# NAND2X1_LOC_571/B VSS VDD NAND2X1_LOC_557/Y
+ NAND2X1_LOC_561/B NAND2X1_LOC
XNAND2X1_LOC_594 NAND2X1_LOC_594/a_36_24# NOR2X1_LOC_653/B VSS VDD INVX1_LOC_57/A
+ NOR2X1_LOC_186/Y NAND2X1_LOC
XNAND2X1_LOC_583 NAND2X1_LOC_583/a_36_24# NOR2X1_LOC_636/B VSS VDD INVX1_LOC_21/A
+ NOR2X1_LOC_68/A NAND2X1_LOC
XNAND2X1_LOC_391 NAND2X1_LOC_391/a_36_24# NAND2X1_LOC_391/Y VSS VDD NOR2X1_LOC_382/Y
+ NOR2X1_LOC_384/Y NAND2X1_LOC
XNAND2X1_LOC_380 NAND2X1_LOC_380/a_36_24# NOR2X1_LOC_460/B VSS VDD INVX1_LOC_76/Y
+ NOR2X1_LOC_379/Y NAND2X1_LOC
XNOR2X1_LOC_807 NOR2X1_LOC_807/a_36_216# NOR2X1_LOC_811/B VSS VDD NOR2X1_LOC_806/Y
+ NOR2X1_LOC_807/B NOR2X1_LOC
XNOR2X1_LOC_829 NOR2X1_LOC_829/a_36_216# NOR2X1_LOC_829/Y VSS VDD NOR2X1_LOC_829/A
+ INVX1_LOC_50/A NOR2X1_LOC
XNOR2X1_LOC_818 NOR2X1_LOC_818/a_36_216# NOR2X1_LOC_818/Y VSS VDD INVX1_LOC_83/A INVX1_LOC_4/Y
+ NOR2X1_LOC
XINVX1_LOC_235 INVX1_LOC_235/Y VSS VDD INVX1_LOC_235/A INVX1_LOC
XINVX1_LOC_224 INVX1_LOC_224/Y VSS VDD INVX1_LOC_224/A INVX1_LOC
XINVX1_LOC_279 INVX1_LOC_279/Y VSS VDD INVX1_LOC_279/A INVX1_LOC
XINVX1_LOC_246 INVX1_LOC_246/Y VSS VDD INVX1_LOC_246/A INVX1_LOC
XINVX1_LOC_202 INVX1_LOC_202/Y VSS VDD INVX1_LOC_202/A INVX1_LOC
XINVX1_LOC_213 INVX1_LOC_213/Y VSS VDD INVX1_LOC_213/A INVX1_LOC
XINVX1_LOC_257 INVX1_LOC_257/Y VSS VDD INVX1_LOC_257/A INVX1_LOC
XINVX1_LOC_268 INVX1_LOC_268/Y VSS VDD INVX1_LOC_268/A INVX1_LOC
XNOR2X1_LOC_604 NOR2X1_LOC_604/a_36_216# NOR2X1_LOC_604/Y VSS VDD INVX1_LOC_92/A INVX1_LOC_54/A
+ NOR2X1_LOC
XNOR2X1_LOC_626 NOR2X1_LOC_626/a_36_216# NOR2X1_LOC_626/Y VSS VDD INVX1_LOC_92/A INVX1_LOC_58/A
+ NOR2X1_LOC
XNAND2X1_LOC_13 NAND2X1_LOC_13/a_36_24# NOR2X1_LOC_538/B VSS VDD INVX1_LOC_9/A INVX1_LOC_11/A
+ NAND2X1_LOC
XNAND2X1_LOC_57 NAND2X1_LOC_57/a_36_24# INVX1_LOC_43/A VSS VDD INVX1_LOC_4/Y INVX1_LOC_33/A
+ NAND2X1_LOC
XNAND2X1_LOC_79 NAND2X1_LOC_79/a_36_24# NAND2X1_LOC_79/Y VSS VDD INVX1_LOC_16/Y NOR2X1_LOC_78/Y
+ NAND2X1_LOC
XNAND2X1_LOC_35 NAND2X1_LOC_35/a_36_24# NAND2X1_LOC_35/Y VSS VDD NAND2X1_LOC_33/Y
+ NAND2X1_LOC_35/B NAND2X1_LOC
XNAND2X1_LOC_24 NAND2X1_LOC_24/a_36_24# NOR2X1_LOC_33/A VSS VDD INVX1_LOC_17/A NOR2X1_LOC_160/B
+ NAND2X1_LOC
XNAND2X1_LOC_46 NAND2X1_LOC_46/a_36_24# NOR2X1_LOC_598/B VSS VDD D_INPUT_1 INVX1_LOC_13/A
+ NAND2X1_LOC
XNAND2X1_LOC_68 NAND2X1_LOC_68/a_36_24# NOR2X1_LOC_69/A VSS VDD INVX1_LOC_4/A NOR2X1_LOC_52/B
+ NAND2X1_LOC
XNOR2X1_LOC_615 NOR2X1_LOC_615/a_36_216# NOR2X1_LOC_615/Y VSS VDD NOR2X1_LOC_754/A
+ INVX1_LOC_17/Y NOR2X1_LOC
XNOR2X1_LOC_659 NOR2X1_LOC_659/a_36_216# INVX1_LOC_268/A VSS VDD NOR2X1_LOC_658/Y
+ NOR2X1_LOC_657/Y NOR2X1_LOC
XNOR2X1_LOC_637 NOR2X1_LOC_637/a_36_216# NOR2X1_LOC_637/Y VSS VDD NOR2X1_LOC_637/A
+ NOR2X1_LOC_637/B NOR2X1_LOC
XNOR2X1_LOC_648 NOR2X1_LOC_648/a_36_216# NOR2X1_LOC_655/B VSS VDD INVX1_LOC_263/Y
+ NOR2X1_LOC_644/Y NOR2X1_LOC
XNOR2X1_LOC_467 NOR2X1_LOC_467/a_36_216# NOR2X1_LOC_470/A VSS VDD NOR2X1_LOC_467/A
+ NOR2X1_LOC_210/A NOR2X1_LOC
XNOR2X1_LOC_423 NOR2X1_LOC_423/a_36_216# NOR2X1_LOC_423/Y VSS VDD INVX1_LOC_50/A INVX1_LOC_6/A
+ NOR2X1_LOC
XNOR2X1_LOC_456 NOR2X1_LOC_456/a_36_216# NOR2X1_LOC_456/Y VSS VDD NOR2X1_LOC_254/Y
+ INVX1_LOC_99/A NOR2X1_LOC
XNOR2X1_LOC_445 NOR2X1_LOC_445/a_36_216# NOR2X1_LOC_445/Y VSS VDD NOR2X1_LOC_318/B
+ NOR2X1_LOC_445/B NOR2X1_LOC
XNOR2X1_LOC_434 NOR2X1_LOC_434/a_36_216# NOR2X1_LOC_434/Y VSS VDD NOR2X1_LOC_434/A
+ NOR2X1_LOC_174/A NOR2X1_LOC
XNOR2X1_LOC_412 NOR2X1_LOC_412/a_36_216# NOR2X1_LOC_690/A VSS VDD INVX1_LOC_34/A INVX1_LOC_25/Y
+ NOR2X1_LOC
XNOR2X1_LOC_401 NOR2X1_LOC_401/a_36_216# NOR2X1_LOC_401/Y VSS VDD NOR2X1_LOC_401/A
+ NOR2X1_LOC_401/B NOR2X1_LOC
XNOR2X1_LOC_478 NOR2X1_LOC_478/a_36_216# INVX1_LOC_204/A VSS VDD NOR2X1_LOC_478/A
+ INVX1_LOC_199/Y NOR2X1_LOC
XNOR2X1_LOC_489 NOR2X1_LOC_489/a_36_216# NOR2X1_LOC_772/B VSS VDD NOR2X1_LOC_489/A
+ NOR2X1_LOC_489/B NOR2X1_LOC
XNAND2X1_LOC_209 NAND2X1_LOC_209/a_36_24# NAND2X1_LOC_213/A VSS VDD NAND2X1_LOC_149/Y
+ NOR2X1_LOC_152/Y NAND2X1_LOC
XNOR2X1_LOC_275 NOR2X1_LOC_275/a_36_216# INVX1_LOC_130/A VSS VDD NOR2X1_LOC_275/A
+ INPUT_0 NOR2X1_LOC
XNOR2X1_LOC_220 NOR2X1_LOC_220/a_36_216# INVX1_LOC_116/A VSS VDD NOR2X1_LOC_220/A
+ NOR2X1_LOC_220/B NOR2X1_LOC
XNOR2X1_LOC_297 NOR2X1_LOC_297/a_36_216# INVX1_LOC_138/A VSS VDD NOR2X1_LOC_297/A
+ INVX1_LOC_34/A NOR2X1_LOC
XNOR2X1_LOC_242 NOR2X1_LOC_242/a_36_216# NOR2X1_LOC_244/B VSS VDD NOR2X1_LOC_242/A
+ INVX1_LOC_120/Y NOR2X1_LOC
XNOR2X1_LOC_253 NOR2X1_LOC_253/a_36_216# NOR2X1_LOC_253/Y VSS VDD INVX1_LOC_78/A INVX1_LOC_50/A
+ NOR2X1_LOC
XNOR2X1_LOC_286 NOR2X1_LOC_286/a_36_216# NOR2X1_LOC_286/Y VSS VDD NOR2X1_LOC_285/Y
+ INVX1_LOC_132/Y NOR2X1_LOC
XNOR2X1_LOC_264 NOR2X1_LOC_264/a_36_216# NOR2X1_LOC_264/Y VSS VDD NOR2X1_LOC_78/A
+ INVX1_LOC_9/A NOR2X1_LOC
XNOR2X1_LOC_231 NOR2X1_LOC_231/a_36_216# NOR2X1_LOC_641/B VSS VDD NOR2X1_LOC_231/A
+ NOR2X1_LOC_231/B NOR2X1_LOC
XNAND2X1_LOC_710 NAND2X1_LOC_710/a_36_24# NAND2X1_LOC_711/B VSS VDD NOR2X1_LOC_700/Y
+ NOR2X1_LOC_701/Y NAND2X1_LOC
XNAND2X1_LOC_721 NAND2X1_LOC_721/a_36_24# NAND2X1_LOC_734/B VSS VDD NAND2X1_LOC_721/A
+ NAND2X1_LOC_721/B NAND2X1_LOC
XNAND2X1_LOC_754 NAND2X1_LOC_754/a_36_24# NOR2X1_LOC_790/A VSS VDD INVX1_LOC_24/Y
+ NOR2X1_LOC_614/Y NAND2X1_LOC
XNAND2X1_LOC_732 NAND2X1_LOC_732/a_36_24# NAND2X1_LOC_738/B VSS VDD NAND2X1_LOC_724/Y
+ NAND2X1_LOC_725/Y NAND2X1_LOC
XNAND2X1_LOC_743 NAND2X1_LOC_743/a_36_24# NOR2X1_LOC_780/B VSS VDD INVX1_LOC_1/A NOR2X1_LOC_155/A
+ NAND2X1_LOC
XNAND2X1_LOC_787 NAND2X1_LOC_787/a_36_24# NAND2X1_LOC_787/Y VSS VDD NAND2X1_LOC_787/A
+ NAND2X1_LOC_787/B NAND2X1_LOC
XNAND2X1_LOC_776 NAND2X1_LOC_776/a_36_24# NAND2X1_LOC_785/B VSS VDD NOR2X1_LOC_164/Y
+ NOR2X1_LOC_238/Y NAND2X1_LOC
XNAND2X1_LOC_798 NAND2X1_LOC_798/a_36_24# NAND2X1_LOC_802/A VSS VDD NAND2X1_LOC_798/A
+ NAND2X1_LOC_798/B NAND2X1_LOC
XNAND2X1_LOC_765 NAND2X1_LOC_765/a_36_24# NOR2X1_LOC_770/B VSS VDD INVX1_LOC_11/A
+ NOR2X1_LOC_78/B NAND2X1_LOC
XINVX1_LOC_9 INVX1_LOC_9/Y VSS VDD INVX1_LOC_9/A INVX1_LOC
XNAND2X1_LOC_551 NAND2X1_LOC_551/a_36_24# NAND2X1_LOC_564/A VSS VDD NAND2X1_LOC_551/A
+ INVX1_LOC_224/Y NAND2X1_LOC
XNAND2X1_LOC_540 NAND2X1_LOC_540/a_36_24# NAND2X1_LOC_553/A VSS VDD NOR2X1_LOC_178/Y
+ INVX1_LOC_98/A NAND2X1_LOC
XNAND2X1_LOC_595 NAND2X1_LOC_595/a_36_24# NOR2X1_LOC_643/A VSS VDD INVX1_LOC_20/Y
+ NOR2X1_LOC_249/Y NAND2X1_LOC
XNAND2X1_LOC_562 NAND2X1_LOC_562/a_36_24# NAND2X1_LOC_562/Y VSS VDD NAND2X1_LOC_555/Y
+ NAND2X1_LOC_562/B NAND2X1_LOC
XNAND2X1_LOC_573 NAND2X1_LOC_573/a_36_24# NAND2X1_LOC_573/Y VSS VDD NAND2X1_LOC_573/A
+ INVX1_LOC_208/Y NAND2X1_LOC
XNAND2X1_LOC_584 NAND2X1_LOC_584/a_36_24# NOR2X1_LOC_636/A VSS VDD INVX1_LOC_5/A INVX1_LOC_37/A
+ NAND2X1_LOC
XNOR2X1_LOC_808 NOR2X1_LOC_808/a_36_216# NOR2X1_LOC_811/A VSS VDD NOR2X1_LOC_808/A
+ NOR2X1_LOC_808/B NOR2X1_LOC
XNAND2X1_LOC_370 NAND2X1_LOC_370/a_36_24# NAND2X1_LOC_787/A VSS VDD NOR2X1_LOC_309/Y
+ NOR2X1_LOC_369/Y NAND2X1_LOC
XNAND2X1_LOC_392 NAND2X1_LOC_392/a_36_24# NAND2X1_LOC_392/Y VSS VDD NAND2X1_LOC_392/A
+ NAND2X1_LOC_391/Y NAND2X1_LOC
XNAND2X1_LOC_381 NAND2X1_LOC_381/a_36_24# NAND2X1_LOC_381/Y VSS VDD INPUT_3 INVX1_LOC_11/A
+ NAND2X1_LOC
XNOR2X1_LOC_819 NOR2X1_LOC_819/a_36_216# NOR2X1_LOC_820/A VSS VDD INVX1_LOC_40/Y INVX1_LOC_36/A
+ NOR2X1_LOC
XINVX1_LOC_203 INVX1_LOC_203/Y VSS VDD INVX1_LOC_203/A INVX1_LOC
XINVX1_LOC_225 INVX1_LOC_225/Y VSS VDD INVX1_LOC_225/A INVX1_LOC
XINVX1_LOC_214 INVX1_LOC_214/Y VSS VDD INVX1_LOC_214/A INVX1_LOC
XNAND2X1_LOC_14 NAND2X1_LOC_14/a_36_24# INVX1_LOC_13/A VSS VDD D_INPUT_2 D_INPUT_3
+ NAND2X1_LOC
XNAND2X1_LOC_25 NAND2X1_LOC_25/a_36_24# NAND2X1_LOC_59/B VSS VDD INPUT_6 D_INPUT_7
+ NAND2X1_LOC
XINVX1_LOC_258 INVX1_LOC_258/Y VSS VDD INVX1_LOC_258/A INVX1_LOC
XINVX1_LOC_269 INVX1_LOC_269/Y VSS VDD INVX1_LOC_269/A INVX1_LOC
XINVX1_LOC_236 INVX1_LOC_236/Y VSS VDD INVX1_LOC_236/A INVX1_LOC
XINVX1_LOC_247 INVX1_LOC_247/Y VSS VDD INVX1_LOC_247/A INVX1_LOC
XNOR2X1_LOC_638 NOR2X1_LOC_638/a_36_216# NOR2X1_LOC_638/Y VSS VDD NOR2X1_LOC_637/Y
+ INVX1_LOC_244/Y NOR2X1_LOC
XNOR2X1_LOC_627 NOR2X1_LOC_627/a_36_216# NOR2X1_LOC_627/Y VSS VDD INVX1_LOC_24/A INVX1_LOC_6/A
+ NOR2X1_LOC
XNOR2X1_LOC_605 NOR2X1_LOC_605/a_36_216# INVX1_LOC_250/A VSS VDD NOR2X1_LOC_605/A
+ NOR2X1_LOC_605/B NOR2X1_LOC
XNAND2X1_LOC_69 NAND2X1_LOC_69/a_36_24# INVX1_LOC_51/A VSS VDD INVX1_LOC_24/Y NOR2X1_LOC_68/Y
+ NAND2X1_LOC
XNAND2X1_LOC_58 NAND2X1_LOC_58/a_36_24# NOR2X1_LOC_61/B VSS VDD INVX1_LOC_17/A NOR2X1_LOC_68/A
+ NAND2X1_LOC
XNAND2X1_LOC_47 NAND2X1_LOC_47/a_36_24# INVX1_LOC_35/A VSS VDD NAND2X1_LOC_59/B NAND2X1_LOC_30/Y
+ NAND2X1_LOC
XNAND2X1_LOC_36 NAND2X1_LOC_36/a_36_24# INVX1_LOC_23/A VSS VDD NAND2X1_LOC_36/A NAND2X1_LOC_21/Y
+ NAND2X1_LOC
XNOR2X1_LOC_649 NOR2X1_LOC_649/a_36_216# NOR2X1_LOC_649/Y VSS VDD NOR2X1_LOC_643/Y
+ NOR2X1_LOC_649/B NOR2X1_LOC
XNOR2X1_LOC_616 NOR2X1_LOC_616/a_36_216# NOR2X1_LOC_616/Y VSS VDD INVX1_LOC_64/A INVX1_LOC_15/Y
+ NOR2X1_LOC
XNOR2X1_LOC_424 NOR2X1_LOC_424/a_36_216# NOR2X1_LOC_424/Y VSS VDD NOR2X1_LOC_89/A
+ INVX1_LOC_34/A NOR2X1_LOC
XNOR2X1_LOC_435 NOR2X1_LOC_435/a_36_216# INVX1_LOC_180/A VSS VDD NOR2X1_LOC_435/A
+ NOR2X1_LOC_435/B NOR2X1_LOC
XNOR2X1_LOC_457 NOR2X1_LOC_457/a_36_216# NOR2X1_LOC_464/B VSS VDD NOR2X1_LOC_457/A
+ NOR2X1_LOC_457/B NOR2X1_LOC
XNOR2X1_LOC_446 NOR2X1_LOC_446/a_36_216# INVX1_LOC_188/A VSS VDD NOR2X1_LOC_446/A
+ INVX1_LOC_177/A NOR2X1_LOC
XNOR2X1_LOC_479 NOR2X1_LOC_479/a_36_216# NOR2X1_LOC_480/A VSS VDD NOR2X1_LOC_476/Y
+ NOR2X1_LOC_479/B NOR2X1_LOC
XNOR2X1_LOC_413 NOR2X1_LOC_413/a_36_216# NOR2X1_LOC_413/Y VSS VDD NOR2X1_LOC_690/A
+ D_INPUT_0 NOR2X1_LOC
XNOR2X1_LOC_402 NOR2X1_LOC_402/a_36_216# INVX1_LOC_168/A VSS VDD NOR2X1_LOC_401/Y
+ INVX1_LOC_164/Y NOR2X1_LOC
XNOR2X1_LOC_468 NOR2X1_LOC_468/a_36_216# NOR2X1_LOC_468/Y VSS VDD NOR2X1_LOC_440/Y
+ NOR2X1_LOC_798/A NOR2X1_LOC
XNOR2X1_LOC_221 NOR2X1_LOC_221/a_36_216# NOR2X1_LOC_223/B VSS VDD INVX1_LOC_115/Y
+ INVX1_LOC_103/Y NOR2X1_LOC
XNOR2X1_LOC_210 NOR2X1_LOC_210/a_36_216# INVX1_LOC_114/A VSS VDD NOR2X1_LOC_210/A
+ NOR2X1_LOC_210/B NOR2X1_LOC
XNOR2X1_LOC_254 NOR2X1_LOC_254/a_36_216# NOR2X1_LOC_254/Y VSS VDD NOR2X1_LOC_254/A
+ NOR2X1_LOC_483/B NOR2X1_LOC
XNOR2X1_LOC_276 NOR2X1_LOC_276/a_36_216# NOR2X1_LOC_276/Y VSS VDD INVX1_LOC_130/Y
+ NOR2X1_LOC_276/B NOR2X1_LOC
XNOR2X1_LOC_287 NOR2X1_LOC_287/a_36_216# NOR2X1_LOC_288/A VSS VDD NOR2X1_LOC_287/A
+ NOR2X1_LOC_843/A NOR2X1_LOC
XNOR2X1_LOC_265 NOR2X1_LOC_265/a_36_216# INVX1_LOC_126/A VSS VDD NOR2X1_LOC_667/A
+ INVX1_LOC_30/A NOR2X1_LOC
XNOR2X1_LOC_298 NOR2X1_LOC_298/a_36_216# NOR2X1_LOC_298/Y VSS VDD INVX1_LOC_42/A INVX1_LOC_22/A
+ NOR2X1_LOC
XNOR2X1_LOC_243 NOR2X1_LOC_243/a_36_216# NOR2X1_LOC_243/Y VSS VDD NOR2X1_LOC_240/Y
+ NOR2X1_LOC_243/B NOR2X1_LOC
XNOR2X1_LOC_232 NOR2X1_LOC_232/a_36_216# NOR2X1_LOC_232/Y VSS VDD INVX1_LOC_90/A NOR2X1_LOC_15/Y
+ NOR2X1_LOC
XNAND2X1_LOC_722 NAND2X1_LOC_722/a_36_24# NAND2X1_LOC_733/A VSS VDD NAND2X1_LOC_722/A
+ INVX1_LOC_284/Y NAND2X1_LOC
XNAND2X1_LOC_733 NAND2X1_LOC_733/a_36_24# NAND2X1_LOC_733/Y VSS VDD NAND2X1_LOC_733/A
+ NAND2X1_LOC_733/B NAND2X1_LOC
XNAND2X1_LOC_755 NAND2X1_LOC_755/a_36_24# NOR2X1_LOC_791/B VSS VDD INVX1_LOC_46/Y
+ NOR2X1_LOC_664/Y NAND2X1_LOC
XNAND2X1_LOC_711 NAND2X1_LOC_711/a_36_24# NAND2X1_LOC_711/Y VSS VDD INVX1_LOC_278/Y
+ NAND2X1_LOC_711/B NAND2X1_LOC
XNAND2X1_LOC_777 NAND2X1_LOC_777/a_36_24# NAND2X1_LOC_784/A VSS VDD NOR2X1_LOC_246/A
+ NOR2X1_LOC_305/Y NAND2X1_LOC
XNAND2X1_LOC_788 NAND2X1_LOC_788/a_36_24# NAND2X1_LOC_794/B VSS VDD NOR2X1_LOC_533/Y
+ INVX1_LOC_248/Y NAND2X1_LOC
XNAND2X1_LOC_700 NAND2X1_LOC_700/a_36_24# NOR2X1_LOC_710/B VSS VDD INVX1_LOC_45/A
+ NOR2X1_LOC_383/B NAND2X1_LOC
XNAND2X1_LOC_744 NAND2X1_LOC_744/a_36_24# NOR2X1_LOC_780/A VSS VDD INVX1_LOC_33/A
+ INVX1_LOC_75/A NAND2X1_LOC
XNAND2X1_LOC_766 NAND2X1_LOC_766/a_36_24# NOR2X1_LOC_770/A VSS VDD INVX1_LOC_49/A
+ NOR2X1_LOC_383/B NAND2X1_LOC
XNAND2X1_LOC_799 NAND2X1_LOC_799/a_36_24# NAND2X1_LOC_799/Y VSS VDD NAND2X1_LOC_799/A
+ NAND2X1_LOC_593/Y NAND2X1_LOC
XNAND2X1_LOC_552 NAND2X1_LOC_552/a_36_24# NAND2X1_LOC_564/B VSS VDD NAND2X1_LOC_552/A
+ NAND2X1_LOC_543/Y NAND2X1_LOC
XNAND2X1_LOC_541 NAND2X1_LOC_541/a_36_24# NAND2X1_LOC_541/Y VSS VDD NOR2X1_LOC_255/Y
+ NOR2X1_LOC_272/Y NAND2X1_LOC
XNAND2X1_LOC_574 NAND2X1_LOC_574/a_36_24# INVX1_LOC_235/A VSS VDD NAND2X1_LOC_574/A
+ NOR2X1_LOC_516/Y NAND2X1_LOC
XNAND2X1_LOC_563 NAND2X1_LOC_563/a_36_24# NAND2X1_LOC_563/Y VSS VDD NAND2X1_LOC_563/A
+ INVX1_LOC_228/Y NAND2X1_LOC
XNAND2X1_LOC_530 NAND2X1_LOC_530/a_36_24# NOR2X1_LOC_548/A VSS VDD INVX1_LOC_23/A
+ NOR2X1_LOC_590/A NAND2X1_LOC
XNAND2X1_LOC_585 NAND2X1_LOC_585/a_36_24# NOR2X1_LOC_637/B VSS VDD INVX1_LOC_17/A
+ INVX1_LOC_135/A NAND2X1_LOC
XNAND2X1_LOC_596 NAND2X1_LOC_596/a_36_24# NOR2X1_LOC_597/A VSS VDD INVX1_LOC_34/A
+ NOR2X1_LOC_328/Y NAND2X1_LOC
XNOR2X1_LOC_809 NOR2X1_LOC_809/a_36_216# NOR2X1_LOC_810/A VSS VDD NOR2X1_LOC_809/A
+ NOR2X1_LOC_809/B NOR2X1_LOC
XNAND2X1_LOC_360 NAND2X1_LOC_360/a_36_24# NAND2X1_LOC_363/B VSS VDD NAND2X1_LOC_860/A
+ NAND2X1_LOC_360/B NAND2X1_LOC
XNAND2X1_LOC_393 NAND2X1_LOC_393/a_36_24# NOR2X1_LOC_400/B VSS VDD INVX1_LOC_27/A
+ INVX1_LOC_29/A NAND2X1_LOC
XNAND2X1_LOC_382 NAND2X1_LOC_382/a_36_24# NOR2X1_LOC_391/B VSS VDD NOR2X1_LOC_82/A
+ NAND2X1_LOC_381/Y NAND2X1_LOC
XNAND2X1_LOC_371 NAND2X1_LOC_371/a_36_24# NOR2X1_LOC_778/B VSS VDD INVX1_LOC_4/Y INVX1_LOC_21/A
+ NAND2X1_LOC
XINVX1_LOC_237 INVX1_LOC_237/Y VSS VDD INVX1_LOC_237/A INVX1_LOC
XINVX1_LOC_226 INVX1_LOC_226/Y VSS VDD INVX1_LOC_226/A INVX1_LOC
XINVX1_LOC_248 INVX1_LOC_248/Y VSS VDD INVX1_LOC_248/A INVX1_LOC
XINVX1_LOC_215 INVX1_LOC_215/Y VSS VDD INVX1_LOC_215/A INVX1_LOC
XINVX1_LOC_259 INVX1_LOC_259/Y VSS VDD INVX1_LOC_259/A INVX1_LOC
XINVX1_LOC_204 INVX1_LOC_204/Y VSS VDD INVX1_LOC_204/A INVX1_LOC
XNAND2X1_LOC_15 NAND2X1_LOC_15/a_36_24# NOR2X1_LOC_78/B VSS VDD NAND2X1_LOC_9/Y INVX1_LOC_13/A
+ NAND2X1_LOC
XNAND2X1_LOC_37 NAND2X1_LOC_37/a_36_24# INVX1_LOC_25/A VSS VDD INPUT_2 INPUT_3
+ NAND2X1_LOC
XNAND2X1_LOC_48 NAND2X1_LOC_48/a_36_24# NOR2X1_LOC_196/A VSS VDD NOR2X1_LOC_598/B
+ INVX1_LOC_35/A NAND2X1_LOC
XNAND2X1_LOC_26 NAND2X1_LOC_26/a_36_24# INVX1_LOC_19/A VSS VDD NAND2X1_LOC_21/Y NAND2X1_LOC_59/B
+ NAND2X1_LOC
XNAND2X1_LOC_59 NAND2X1_LOC_59/a_36_24# INVX1_LOC_45/A VSS VDD NAND2X1_LOC_11/Y NAND2X1_LOC_59/B
+ NAND2X1_LOC
XNOR2X1_LOC_639 NOR2X1_LOC_639/a_36_216# NOR2X1_LOC_639/Y VSS VDD INVX1_LOC_261/Y
+ NOR2X1_LOC_639/B NOR2X1_LOC
XNAND2X1_LOC_190 NAND2X1_LOC_190/a_36_24# NAND2X1_LOC_190/Y VSS VDD INVX1_LOC_97/Y
+ INVX1_LOC_99/Y NAND2X1_LOC
XNOR2X1_LOC_628 NOR2X1_LOC_628/a_36_216# INVX1_LOC_258/A VSS VDD NOR2X1_LOC_92/Y INVX1_LOC_36/A
+ NOR2X1_LOC
XNOR2X1_LOC_606 NOR2X1_LOC_606/a_36_216# NOR2X1_LOC_606/Y VSS VDD INVX1_LOC_71/A NOR2X1_LOC_590/A
+ NOR2X1_LOC
XNOR2X1_LOC_617 NOR2X1_LOC_617/a_36_216# NOR2X1_LOC_617/Y VSS VDD INVX1_LOC_37/Y INVX1_LOC_28/A
+ NOR2X1_LOC
XNOR2X1_LOC_425 NOR2X1_LOC_425/a_36_216# NOR2X1_LOC_425/Y VSS VDD NOR2X1_LOC_36/B
+ INPUT_5 NOR2X1_LOC
XNOR2X1_LOC_447 NOR2X1_LOC_447/a_36_216# NOR2X1_LOC_447/Y VSS VDD NOR2X1_LOC_447/A
+ NOR2X1_LOC_447/B NOR2X1_LOC
XNOR2X1_LOC_458 NOR2X1_LOC_458/a_36_216# NOR2X1_LOC_458/Y VSS VDD NOR2X1_LOC_717/B
+ NOR2X1_LOC_458/B NOR2X1_LOC
XNOR2X1_LOC_436 NOR2X1_LOC_436/a_36_216# NOR2X1_LOC_798/A VSS VDD INVX1_LOC_179/Y
+ NOR2X1_LOC_434/Y NOR2X1_LOC
XNOR2X1_LOC_469 NOR2X1_LOC_469/a_36_216# INVX1_LOC_200/A VSS VDD NOR2X1_LOC_468/Y
+ INVX1_LOC_185/Y NOR2X1_LOC
XNOR2X1_LOC_414 NOR2X1_LOC_414/a_36_216# NOR2X1_LOC_414/Y VSS VDD NOR2X1_LOC_6/B D_INPUT_3
+ NOR2X1_LOC
XNOR2X1_LOC_403 NOR2X1_LOC_403/a_36_216# INVX1_LOC_170/A VSS VDD INVX1_LOC_165/Y NOR2X1_LOC_403/B
+ NOR2X1_LOC
XNOR2X1_LOC_200 NOR2X1_LOC_200/a_36_216# NOR2X1_LOC_207/A VSS VDD NOR2X1_LOC_194/Y
+ INVX1_LOC_105/Y NOR2X1_LOC
XNOR2X1_LOC_222 NOR2X1_LOC_222/a_36_216# NOR2X1_LOC_222/Y VSS VDD NOR2X1_LOC_219/Y
+ NOR2X1_LOC_218/Y NOR2X1_LOC
XNOR2X1_LOC_211 NOR2X1_LOC_211/a_36_216# NOR2X1_LOC_211/Y VSS VDD NOR2X1_LOC_211/A
+ INVX1_LOC_93/Y NOR2X1_LOC
XNOR2X1_LOC_233 NOR2X1_LOC_233/a_36_216# NOR2X1_LOC_824/A VSS VDD INVX1_LOC_13/Y D_INPUT_0
+ NOR2X1_LOC
XNOR2X1_LOC_288 NOR2X1_LOC_288/a_36_216# INVX1_LOC_134/A VSS VDD NOR2X1_LOC_288/A
+ NOR2X1_LOC_286/Y NOR2X1_LOC
XNOR2X1_LOC_266 NOR2X1_LOC_266/a_36_216# NOR2X1_LOC_267/A VSS VDD INVX1_LOC_124/Y
+ NOR2X1_LOC_266/B NOR2X1_LOC
XNOR2X1_LOC_299 NOR2X1_LOC_299/a_36_216# NOR2X1_LOC_299/Y VSS VDD INVX1_LOC_72/A INVX1_LOC_11/Y
+ NOR2X1_LOC
XNOR2X1_LOC_244 NOR2X1_LOC_244/a_36_216# NOR2X1_LOC_860/B VSS VDD NOR2X1_LOC_243/Y
+ NOR2X1_LOC_244/B NOR2X1_LOC
XNOR2X1_LOC_255 NOR2X1_LOC_255/a_36_216# NOR2X1_LOC_255/Y VSS VDD INVX1_LOC_89/Y INVX1_LOC_25/Y
+ NOR2X1_LOC
XNOR2X1_LOC_277 NOR2X1_LOC_277/a_36_216# NOR2X1_LOC_278/A VSS VDD INVX1_LOC_36/A INVX1_LOC_25/Y
+ NOR2X1_LOC
XNAND2X1_LOC_778 NAND2X1_LOC_778/a_36_24# NAND2X1_LOC_778/Y VSS VDD NOR2X1_LOC_372/A
+ NOR2X1_LOC_496/Y NAND2X1_LOC
XNAND2X1_LOC_767 NAND2X1_LOC_767/a_36_24# INVX1_LOC_293/A VSS VDD INVX1_LOC_2/Y NOR2X1_LOC_78/Y
+ NAND2X1_LOC
XNAND2X1_LOC_789 NAND2X1_LOC_789/a_36_24# INVX1_LOC_305/A VSS VDD NOR2X1_LOC_748/Y
+ NOR2X1_LOC_751/Y NAND2X1_LOC
XNAND2X1_LOC_734 NAND2X1_LOC_734/a_36_24# INVX1_LOC_285/A VSS VDD INVX1_LOC_172/A
+ NAND2X1_LOC_734/B NAND2X1_LOC
XNAND2X1_LOC_723 NAND2X1_LOC_723/a_36_24# NAND2X1_LOC_733/B VSS VDD INVX1_LOC_282/Y
+ NAND2X1_LOC_717/Y NAND2X1_LOC
XNAND2X1_LOC_756 NAND2X1_LOC_756/a_36_24# NOR2X1_LOC_757/A VSS VDD INVX1_LOC_64/A
+ INVX1_LOC_92/A NAND2X1_LOC
XNAND2X1_LOC_712 NAND2X1_LOC_712/a_36_24# NAND2X1_LOC_725/A VSS VDD NAND2X1_LOC_712/A
+ NAND2X1_LOC_708/Y NAND2X1_LOC
XNAND2X1_LOC_745 NAND2X1_LOC_745/a_36_24# NOR2X1_LOC_781/B VSS VDD INVX1_LOC_29/A
+ INVX1_LOC_91/A NAND2X1_LOC
XNAND2X1_LOC_701 NAND2X1_LOC_701/a_36_24# NOR2X1_LOC_710/A VSS VDD INVX1_LOC_33/A
+ INVX1_LOC_117/A NAND2X1_LOC
XNAND2X1_LOC_520 NAND2X1_LOC_520/a_36_24# INVX1_LOC_217/A VSS VDD NOR2X1_LOC_518/Y
+ NOR2X1_LOC_519/Y NAND2X1_LOC
XNAND2X1_LOC_564 NAND2X1_LOC_564/a_36_24# NAND2X1_LOC_569/A VSS VDD NAND2X1_LOC_564/A
+ NAND2X1_LOC_564/B NAND2X1_LOC
XNAND2X1_LOC_553 NAND2X1_LOC_553/a_36_24# NAND2X1_LOC_563/A VSS VDD NAND2X1_LOC_553/A
+ NAND2X1_LOC_541/Y NAND2X1_LOC
XNAND2X1_LOC_531 NAND2X1_LOC_531/a_36_24# INVX1_LOC_219/A VSS VDD INVX1_LOC_29/A NAND2X1_LOC_74/B
+ NAND2X1_LOC
XNAND2X1_LOC_542 NAND2X1_LOC_542/a_36_24# NAND2X1_LOC_552/A VSS VDD NOR2X1_LOC_280/Y
+ NOR2X1_LOC_312/Y NAND2X1_LOC
XNAND2X1_LOC_575 NAND2X1_LOC_575/a_36_24# NAND2X1_LOC_579/A VSS VDD NAND2X1_LOC_573/Y
+ INVX1_LOC_236/Y NAND2X1_LOC
XNAND2X1_LOC_597 NAND2X1_LOC_597/a_36_24# NOR2X1_LOC_644/B VSS VDD INVX1_LOC_10/Y
+ NOR2X1_LOC_596/Y NAND2X1_LOC
XNAND2X1_LOC_586 NAND2X1_LOC_586/a_36_24# NOR2X1_LOC_637/A VSS VDD INVX1_LOC_53/A
+ NOR2X1_LOC_130/A NAND2X1_LOC
XNAND2X1_LOC_361 NAND2X1_LOC_361/a_36_24# NAND2X1_LOC_361/Y VSS VDD NAND2X1_LOC_572/B
+ NAND2X1_LOC_276/Y NAND2X1_LOC
XNAND2X1_LOC_372 NAND2X1_LOC_372/a_36_24# NOR2X1_LOC_458/B VSS VDD D_INPUT_1 NOR2X1_LOC_778/B
+ NAND2X1_LOC
XNAND2X1_LOC_350 NAND2X1_LOC_350/a_36_24# INVX1_LOC_157/A VSS VDD NAND2X1_LOC_350/A
+ NAND2X1_LOC_350/B NAND2X1_LOC
XNAND2X1_LOC_383 NAND2X1_LOC_383/a_36_24# NOR2X1_LOC_384/A VSS VDD NOR2X1_LOC_91/A
+ INVX1_LOC_118/A NAND2X1_LOC
XNAND2X1_LOC_394 NAND2X1_LOC_394/a_36_24# NOR2X1_LOC_400/A VSS VDD INVX1_LOC_35/A
+ INVX1_LOC_75/A NAND2X1_LOC
XINVX1_LOC_205 INVX1_LOC_205/Y VSS VDD INVX1_LOC_205/A INVX1_LOC
XINVX1_LOC_216 INVX1_LOC_216/Y VSS VDD INVX1_LOC_216/A INVX1_LOC
XINVX1_LOC_238 INVX1_LOC_238/Y VSS VDD INVX1_LOC_238/A INVX1_LOC
XINVX1_LOC_227 INVX1_LOC_227/Y VSS VDD INVX1_LOC_227/A INVX1_LOC
XINVX1_LOC_249 INVX1_LOC_249/Y VSS VDD INVX1_LOC_249/A INVX1_LOC
XNAND2X1_LOC_180 NAND2X1_LOC_180/a_36_24# NAND2X1_LOC_182/A VSS VDD NOR2X1_LOC_176/Y
+ NOR2X1_LOC_177/Y NAND2X1_LOC
XNAND2X1_LOC_49 NAND2X1_LOC_49/a_36_24# NOR2X1_LOC_68/A VSS VDD INVX1_LOC_13/A NOR2X1_LOC_82/A
+ NAND2X1_LOC
XNAND2X1_LOC_38 NAND2X1_LOC_38/a_36_24# INVX1_LOC_27/A VSS VDD NOR2X1_LOC_82/A INVX1_LOC_25/A
+ NAND2X1_LOC
XNAND2X1_LOC_27 NAND2X1_LOC_27/a_36_24# NOR2X1_LOC_34/B VSS VDD INVX1_LOC_5/A INVX1_LOC_19/A
+ NAND2X1_LOC
XNAND2X1_LOC_191 NAND2X1_LOC_191/a_36_24# NAND2X1_LOC_192/B VSS VDD NOR2X1_LOC_187/Y
+ NAND2X1_LOC_190/Y NAND2X1_LOC
XNAND2X1_LOC_16 NAND2X1_LOC_16/a_36_24# NAND2X1_LOC_16/Y VSS VDD INVX1_LOC_1/A NOR2X1_LOC_78/B
+ NAND2X1_LOC
XNOR2X1_LOC_607 NOR2X1_LOC_607/a_36_216# NOR2X1_LOC_607/Y VSS VDD NOR2X1_LOC_607/A
+ INVX1_LOC_16/A NOR2X1_LOC
XNOR2X1_LOC_629 NOR2X1_LOC_629/a_36_216# NOR2X1_LOC_629/Y VSS VDD NOR2X1_LOC_629/A
+ NOR2X1_LOC_629/B NOR2X1_LOC
XNOR2X1_LOC_618 NOR2X1_LOC_618/a_36_216# NOR2X1_LOC_619/A VSS VDD NOR2X1_LOC_38/B
+ INPUT_3 NOR2X1_LOC
XNOR2X1_LOC_415 NOR2X1_LOC_415/a_36_216# NOR2X1_LOC_415/Y VSS VDD NOR2X1_LOC_415/A
+ INVX1_LOC_135/A NOR2X1_LOC
XNOR2X1_LOC_404 NOR2X1_LOC_404/a_36_216# NOR2X1_LOC_474/A VSS VDD INVX1_LOC_169/Y
+ INVX1_LOC_167/Y NOR2X1_LOC
XNOR2X1_LOC_448 NOR2X1_LOC_448/a_36_216# NOR2X1_LOC_448/Y VSS VDD NOR2X1_LOC_448/A
+ NOR2X1_LOC_448/B NOR2X1_LOC
XNOR2X1_LOC_426 NOR2X1_LOC_426/a_36_216# NOR2X1_LOC_426/Y VSS VDD NOR2X1_LOC_425/Y
+ INVX1_LOC_72/A NOR2X1_LOC
XNOR2X1_LOC_437 NOR2X1_LOC_437/a_36_216# NOR2X1_LOC_437/Y VSS VDD INVX1_LOC_88/A INVX1_LOC_45/Y
+ NOR2X1_LOC
XNOR2X1_LOC_459 NOR2X1_LOC_459/a_36_216# INVX1_LOC_194/A VSS VDD NOR2X1_LOC_459/A
+ NOR2X1_LOC_459/B NOR2X1_LOC
XNOR2X1_LOC_223 NOR2X1_LOC_223/a_36_216# D_GATE_222 VSS VDD NOR2X1_LOC_222/Y NOR2X1_LOC_223/B
+ NOR2X1_LOC
XNOR2X1_LOC_245 NOR2X1_LOC_245/a_36_216# NOR2X1_LOC_246/A VSS VDD INVX1_LOC_25/Y INVX1_LOC_20/A
+ NOR2X1_LOC
XNOR2X1_LOC_212 NOR2X1_LOC_212/a_36_216# NOR2X1_LOC_220/B VSS VDD NOR2X1_LOC_211/Y
+ INVX1_LOC_95/Y NOR2X1_LOC
XNOR2X1_LOC_267 NOR2X1_LOC_267/a_36_216# NOR2X1_LOC_361/B VSS VDD NOR2X1_LOC_267/A
+ INVX1_LOC_126/Y NOR2X1_LOC
XNOR2X1_LOC_201 NOR2X1_LOC_201/a_36_216# INVX1_LOC_110/A VSS VDD NOR2X1_LOC_201/A
+ NOR2X1_LOC_61/Y NOR2X1_LOC
XNOR2X1_LOC_256 NOR2X1_LOC_256/a_36_216# NOR2X1_LOC_256/Y VSS VDD NOR2X1_LOC_255/Y
+ NOR2X1_LOC_19/B NOR2X1_LOC
XNOR2X1_LOC_234 NOR2X1_LOC_234/a_36_216# NOR2X1_LOC_234/Y VSS VDD NOR2X1_LOC_824/A
+ INVX1_LOC_35/Y NOR2X1_LOC
XNOR2X1_LOC_289 NOR2X1_LOC_289/a_36_216# NOR2X1_LOC_289/Y VSS VDD NOR2X1_LOC_226/A
+ INVX1_LOC_38/A NOR2X1_LOC
XNOR2X1_LOC_278 NOR2X1_LOC_278/a_36_216# NOR2X1_LOC_278/Y VSS VDD NOR2X1_LOC_278/A
+ NAND2X1_LOC_9/Y NOR2X1_LOC
XNAND2X1_LOC_702 NAND2X1_LOC_702/a_36_24# NAND2X1_LOC_715/B VSS VDD NOR2X1_LOC_45/Y
+ NOR2X1_LOC_135/Y NAND2X1_LOC
XNAND2X1_LOC_713 NAND2X1_LOC_713/a_36_24# NAND2X1_LOC_725/B VSS VDD NAND2X1_LOC_705/Y
+ NAND2X1_LOC_706/Y NAND2X1_LOC
XNAND2X1_LOC_768 NAND2X1_LOC_768/a_36_24# NAND2X1_LOC_768/Y VSS VDD NOR2X1_LOC_103/Y
+ NOR2X1_LOC_134/Y NAND2X1_LOC
XNAND2X1_LOC_757 NAND2X1_LOC_757/a_36_24# NOR2X1_LOC_791/A VSS VDD INVX1_LOC_34/Y
+ NOR2X1_LOC_756/Y NAND2X1_LOC
XNAND2X1_LOC_735 NAND2X1_LOC_735/a_36_24# NAND2X1_LOC_736/B VSS VDD INVX1_LOC_207/A
+ NAND2X1_LOC_735/B NAND2X1_LOC
XNAND2X1_LOC_724 NAND2X1_LOC_724/a_36_24# NAND2X1_LOC_724/Y VSS VDD NAND2X1_LOC_724/A
+ INVX1_LOC_280/Y NAND2X1_LOC
XNAND2X1_LOC_779 NAND2X1_LOC_779/a_36_24# NAND2X1_LOC_783/A VSS VDD INVX1_LOC_214/A
+ NOR2X1_LOC_697/Y NAND2X1_LOC
XNAND2X1_LOC_746 NAND2X1_LOC_746/a_36_24# NOR2X1_LOC_781/A VSS VDD NAND2X1_LOC_74/B
+ INVX1_LOC_89/A NAND2X1_LOC
XNOR2X1_LOC_790 NOR2X1_LOC_790/a_36_216# NOR2X1_LOC_793/A VSS VDD NOR2X1_LOC_790/A
+ NOR2X1_LOC_790/B NOR2X1_LOC
XNAND2X1_LOC_543 NAND2X1_LOC_543/a_36_24# NAND2X1_LOC_543/Y VSS VDD NOR2X1_LOC_315/Y
+ NOR2X1_LOC_369/Y NAND2X1_LOC
XNAND2X1_LOC_521 NAND2X1_LOC_521/a_36_24# NOR2X1_LOC_523/B VSS VDD INVX1_LOC_15/A
+ NOR2X1_LOC_68/A NAND2X1_LOC
XNAND2X1_LOC_510 NAND2X1_LOC_510/a_36_24# NAND2X1_LOC_574/A VSS VDD NAND2X1_LOC_510/A
+ INVX1_LOC_212/Y NAND2X1_LOC
XNAND2X1_LOC_532 NAND2X1_LOC_532/a_36_24# NOR2X1_LOC_533/A VSS VDD NOR2X1_LOC_536/A
+ INVX1_LOC_76/A NAND2X1_LOC
XNAND2X1_LOC_554 NAND2X1_LOC_554/a_36_24# INVX1_LOC_227/A VSS VDD NOR2X1_LOC_106/Y
+ NAND2X1_LOC_140/A NAND2X1_LOC
XNAND2X1_LOC_565 NAND2X1_LOC_565/a_36_24# NAND2X1_LOC_569/B VSS VDD NAND2X1_LOC_549/Y
+ NAND2X1_LOC_565/B NAND2X1_LOC
XNAND2X1_LOC_576 NAND2X1_LOC_576/a_36_24# INVX1_LOC_237/A VSS VDD NAND2X1_LOC_571/Y
+ INVX1_LOC_234/Y NAND2X1_LOC
XNAND2X1_LOC_598 NAND2X1_LOC_598/a_36_24# NOR2X1_LOC_599/A VSS VDD NOR2X1_LOC_48/B
+ INVX1_LOC_136/A NAND2X1_LOC
XNAND2X1_LOC_587 NAND2X1_LOC_587/a_36_24# NAND2X1_LOC_588/B VSS VDD D_INPUT_7
+ NAND2X1_LOC_30/Y NAND2X1_LOC
XNAND2X1_LOC_362 NAND2X1_LOC_362/a_36_24# NAND2X1_LOC_366/A VSS VDD INVX1_LOC_134/Y
+ NAND2X1_LOC_361/Y NAND2X1_LOC
XNAND2X1_LOC_395 NAND2X1_LOC_395/a_36_24# NOR2X1_LOC_401/B VSS VDD INVX1_LOC_45/A
+ INVX1_LOC_63/A NAND2X1_LOC
XNAND2X1_LOC_384 NAND2X1_LOC_384/a_36_24# NOR2X1_LOC_391/A VSS VDD INVX1_LOC_30/Y
+ NOR2X1_LOC_383/Y NAND2X1_LOC
XNAND2X1_LOC_351 NAND2X1_LOC_351/a_36_24# NAND2X1_LOC_358/B VSS VDD NAND2X1_LOC_351/A
+ INVX1_LOC_152/Y NAND2X1_LOC
XNAND2X1_LOC_373 NAND2X1_LOC_373/a_36_24# NOR2X1_LOC_374/A VSS VDD INVX1_LOC_19/A
+ NOR2X1_LOC_78/A NAND2X1_LOC
XNAND2X1_LOC_340 NAND2X1_LOC_340/a_36_24# NAND2X1_LOC_350/A VSS VDD NOR2X1_LOC_88/Y
+ NAND2X1_LOC_227/Y NAND2X1_LOC
XINVX1_LOC_239 INVX1_LOC_239/Y VSS VDD INVX1_LOC_239/A INVX1_LOC
XINVX1_LOC_228 INVX1_LOC_228/Y VSS VDD INVX1_LOC_228/A INVX1_LOC
XINVX1_LOC_217 INVX1_LOC_217/Y VSS VDD INVX1_LOC_217/A INVX1_LOC
XINVX1_LOC_206 INVX1_LOC_206/Y VSS VDD INVX1_LOC_206/A INVX1_LOC
XNAND2X1_LOC_181 NAND2X1_LOC_181/a_36_24# NAND2X1_LOC_181/Y VSS VDD NOR2X1_LOC_178/Y
+ NOR2X1_LOC_179/Y NAND2X1_LOC
XNAND2X1_LOC_28 NAND2X1_LOC_28/a_36_24# NOR2X1_LOC_82/A VSS VDD D_INPUT_0 INPUT_1
+ NAND2X1_LOC
XNAND2X1_LOC_170 NAND2X1_LOC_170/a_36_24# INVX1_LOC_93/A VSS VDD NAND2X1_LOC_170/A
+ NAND2X1_LOC_169/Y NAND2X1_LOC
XNAND2X1_LOC_192 NAND2X1_LOC_192/a_36_24# INVX1_LOC_103/A VSS VDD INVX1_LOC_101/Y
+ NAND2X1_LOC_192/B NAND2X1_LOC
XNAND2X1_LOC_39 NAND2X1_LOC_39/a_36_24# NAND2X1_LOC_39/Y VSS VDD INVX1_LOC_23/A INVX1_LOC_27/A
+ NAND2X1_LOC
XNAND2X1_LOC_17 NAND2X1_LOC_17/a_36_24# NAND2X1_LOC_36/A VSS VDD INPUT_6 INPUT_7
+ NAND2X1_LOC
XNOR2X1_LOC_608 NOR2X1_LOC_608/a_36_216# NOR2X1_LOC_608/Y VSS VDD NAND2X1_LOC_74/B
+ NOR2X1_LOC_78/B NOR2X1_LOC
XNOR2X1_LOC_619 NOR2X1_LOC_619/a_36_216# INVX1_LOC_254/A VSS VDD NOR2X1_LOC_619/A
+ INVX1_LOC_24/A NOR2X1_LOC
XNOR2X1_LOC_427 NOR2X1_LOC_427/a_36_216# NOR2X1_LOC_427/Y VSS VDD INVX1_LOC_78/A INVX1_LOC_54/A
+ NOR2X1_LOC
XNOR2X1_LOC_449 NOR2X1_LOC_449/a_36_216# INVX1_LOC_190/A VSS VDD NOR2X1_LOC_449/A
+ NOR2X1_LOC_592/B NOR2X1_LOC
XNOR2X1_LOC_405 NOR2X1_LOC_405/a_36_216# NOR2X1_LOC_405/Y VSS VDD NOR2X1_LOC_405/A
+ NOR2X1_LOC_598/B NOR2X1_LOC
XNOR2X1_LOC_416 NOR2X1_LOC_416/a_36_216# INVX1_LOC_176/A VSS VDD NOR2X1_LOC_416/A
+ INVX1_LOC_90/A NOR2X1_LOC
XNOR2X1_LOC_438 NOR2X1_LOC_438/a_36_216# NOR2X1_LOC_438/Y VSS VDD INVX1_LOC_54/A NOR2X1_LOC_45/B
+ NOR2X1_LOC
XNOR2X1_LOC_257 NOR2X1_LOC_257/a_36_216# NOR2X1_LOC_257/Y VSS VDD INVX1_LOC_78/A INVX1_LOC_16/A
+ NOR2X1_LOC
XNOR2X1_LOC_213 NOR2X1_LOC_213/a_36_216# NOR2X1_LOC_220/A VSS VDD INVX1_LOC_113/Y
+ NOR2X1_LOC_209/Y NOR2X1_LOC
XNOR2X1_LOC_224 NOR2X1_LOC_224/a_36_216# NOR2X1_LOC_224/Y VSS VDD INVX1_LOC_76/A INVX1_LOC_22/A
+ NOR2X1_LOC
XNOR2X1_LOC_202 NOR2X1_LOC_202/a_36_216# NOR2X1_LOC_202/Y VSS VDD INVX1_LOC_52/Y NAND2X1_LOC_67/Y
+ NOR2X1_LOC
XNOR2X1_LOC_268 NOR2X1_LOC_268/a_36_216# INVX1_LOC_128/A VSS VDD NOR2X1_LOC_92/Y INVX1_LOC_24/A
+ NOR2X1_LOC
XNOR2X1_LOC_279 NOR2X1_LOC_279/a_36_216# NOR2X1_LOC_279/Y VSS VDD INVX1_LOC_78/A INVX1_LOC_33/Y
+ NOR2X1_LOC
XNOR2X1_LOC_246 NOR2X1_LOC_246/a_36_216# NOR2X1_LOC_246/Y VSS VDD NOR2X1_LOC_246/A
+ NOR2X1_LOC_9/Y NOR2X1_LOC
XNOR2X1_LOC_235 NOR2X1_LOC_235/a_36_216# NOR2X1_LOC_235/Y VSS VDD NOR2X1_LOC_86/A
+ INVX1_LOC_48/Y NOR2X1_LOC
XNAND2X1_LOC_736 NAND2X1_LOC_736/a_36_24# NAND2X1_LOC_736/Y VSS VDD INVX1_LOC_269/A
+ NAND2X1_LOC_736/B NAND2X1_LOC
XNAND2X1_LOC_725 NAND2X1_LOC_725/a_36_24# NAND2X1_LOC_725/Y VSS VDD NAND2X1_LOC_725/A
+ NAND2X1_LOC_725/B NAND2X1_LOC
XNAND2X1_LOC_703 NAND2X1_LOC_703/a_36_24# NAND2X1_LOC_703/Y VSS VDD NOR2X1_LOC_167/Y
+ NOR2X1_LOC_312/Y NAND2X1_LOC
XNAND2X1_LOC_714 NAND2X1_LOC_714/a_36_24# NAND2X1_LOC_724/A VSS VDD NAND2X1_LOC_703/Y
+ NAND2X1_LOC_714/B NAND2X1_LOC
XNAND2X1_LOC_758 NAND2X1_LOC_758/a_36_24# NOR2X1_LOC_759/A VSS VDD INVX1_LOC_30/A
+ INVX1_LOC_58/A NAND2X1_LOC
XNAND2X1_LOC_747 NAND2X1_LOC_747/a_36_24# INVX1_LOC_287/A VSS VDD INVX1_LOC_35/A NOR2X1_LOC_68/A
+ NAND2X1_LOC
XNAND2X1_LOC_769 NAND2X1_LOC_769/a_36_24# INVX1_LOC_295/A VSS VDD NOR2X1_LOC_763/Y
+ NOR2X1_LOC_764/Y NAND2X1_LOC
XNOR2X1_LOC_780 NOR2X1_LOC_780/a_36_216# NOR2X1_LOC_783/A VSS VDD NOR2X1_LOC_780/A
+ NOR2X1_LOC_780/B NOR2X1_LOC
XNOR2X1_LOC_791 NOR2X1_LOC_791/a_36_216# NOR2X1_LOC_791/Y VSS VDD NOR2X1_LOC_791/A
+ NOR2X1_LOC_791/B NOR2X1_LOC
XNAND2X1_LOC_500 NAND2X1_LOC_500/a_36_24# NAND2X1_LOC_500/Y VSS VDD NOR2X1_LOC_497/Y
+ NAND2X1_LOC_500/B NAND2X1_LOC
XNAND2X1_LOC_544 NAND2X1_LOC_544/a_36_24# NAND2X1_LOC_551/A VSS VDD NOR2X1_LOC_373/Y
+ NOR2X1_LOC_438/Y NAND2X1_LOC
XNAND2X1_LOC_522 NAND2X1_LOC_522/a_36_24# NOR2X1_LOC_523/A VSS VDD INVX1_LOC_17/A
+ NOR2X1_LOC_590/A NAND2X1_LOC
XNAND2X1_LOC_555 NAND2X1_LOC_555/a_36_24# NAND2X1_LOC_555/Y VSS VDD INVX1_LOC_122/Y
+ INVX1_LOC_205/Y NAND2X1_LOC
XNAND2X1_LOC_577 NAND2X1_LOC_577/a_36_24# NAND2X1_LOC_578/B VSS VDD NAND2X1_LOC_577/A
+ NAND2X1_LOC_570/Y NAND2X1_LOC
XNAND2X1_LOC_533 NAND2X1_LOC_533/a_36_24# NOR2X1_LOC_788/B VSS VDD INVX1_LOC_58/Y
+ NOR2X1_LOC_532/Y NAND2X1_LOC
XNAND2X1_LOC_566 NAND2X1_LOC_566/a_36_24# NAND2X1_LOC_568/A VSS VDD INVX1_LOC_94/Y
+ NAND2X1_LOC_303/Y NAND2X1_LOC
XNAND2X1_LOC_511 NAND2X1_LOC_511/a_36_24# INVX1_LOC_213/A VSS VDD INVX1_LOC_21/A NOR2X1_LOC_598/B
+ NAND2X1_LOC
XNAND2X1_LOC_588 NAND2X1_LOC_588/a_36_24# INVX1_LOC_243/A VSS VDD INVX1_LOC_83/A NAND2X1_LOC_588/B
+ NAND2X1_LOC
XNAND2X1_LOC_599 NAND2X1_LOC_599/a_36_24# NOR2X1_LOC_644/A VSS VDD INVX1_LOC_24/Y
+ NOR2X1_LOC_828/A NAND2X1_LOC
XNAND2X1_LOC_396 NAND2X1_LOC_396/a_36_24# NOR2X1_LOC_401/A VSS VDD NOR2X1_LOC_160/B
+ INVX1_LOC_23/A NAND2X1_LOC
XNAND2X1_LOC_374 NAND2X1_LOC_374/a_36_24# NAND2X1_LOC_374/Y VSS VDD NOR2X1_LOC_322/Y
+ NOR2X1_LOC_373/Y NAND2X1_LOC
XNAND2X1_LOC_363 NAND2X1_LOC_363/a_36_24# NAND2X1_LOC_363/Y VSS VDD NAND2X1_LOC_359/Y
+ NAND2X1_LOC_363/B NAND2X1_LOC
XNAND2X1_LOC_385 NAND2X1_LOC_385/a_36_24# NOR2X1_LOC_389/B VSS VDD INVX1_LOC_19/A
+ INVX1_LOC_63/A NAND2X1_LOC
XNAND2X1_LOC_352 NAND2X1_LOC_352/a_36_24# NAND2X1_LOC_357/A VSS VDD INVX1_LOC_95/A
+ NAND2X1_LOC_352/B NAND2X1_LOC
XNAND2X1_LOC_330 NAND2X1_LOC_330/a_36_24# INVX1_LOC_145/A VSS VDD INVX1_LOC_38/A INVX1_LOC_53/Y
+ NAND2X1_LOC
XNAND2X1_LOC_341 NAND2X1_LOC_341/a_36_24# NAND2X1_LOC_350/B VSS VDD NAND2X1_LOC_341/A
+ NAND2X1_LOC_231/Y NAND2X1_LOC
XINVX1_LOC_207 INVX1_LOC_207/Y VSS VDD INVX1_LOC_207/A INVX1_LOC
XINVX1_LOC_229 INVX1_LOC_229/Y VSS VDD INVX1_LOC_229/A INVX1_LOC
XINVX1_LOC_218 INVX1_LOC_218/Y VSS VDD INVX1_LOC_218/A INVX1_LOC
XNOR2X1_LOC_609 NOR2X1_LOC_609/a_36_216# NOR2X1_LOC_609/Y VSS VDD NOR2X1_LOC_609/A
+ INVX1_LOC_45/Y NOR2X1_LOC
XNAND2X1_LOC_182 NAND2X1_LOC_182/a_36_24# INVX1_LOC_95/A VSS VDD NAND2X1_LOC_182/A
+ NAND2X1_LOC_181/Y NAND2X1_LOC
XNAND2X1_LOC_29 NAND2X1_LOC_29/a_36_24# NOR2X1_LOC_87/B VSS VDD INVX1_LOC_7/A NOR2X1_LOC_38/B
+ NAND2X1_LOC
XNAND2X1_LOC_171 NAND2X1_LOC_171/a_36_24# NOR2X1_LOC_174/B VSS VDD NOR2X1_LOC_160/B
+ INVX1_LOC_29/A NAND2X1_LOC
XNAND2X1_LOC_193 NAND2X1_LOC_193/a_36_24# INVX1_LOC_105/A VSS VDD NOR2X1_LOC_7/Y NOR2X1_LOC_13/Y
+ NAND2X1_LOC
XNAND2X1_LOC_160 NAND2X1_LOC_160/a_36_24# NAND2X1_LOC_162/A VSS VDD NOR2X1_LOC_45/B
+ INVX1_LOC_76/A NAND2X1_LOC
XNAND2X1_LOC_18 NAND2X1_LOC_18/a_36_24# INVX1_LOC_15/A VSS VDD NAND2X1_LOC_11/Y NAND2X1_LOC_36/A
+ NAND2X1_LOC
XNOR2X1_LOC_428 NOR2X1_LOC_428/a_36_216# NOR2X1_LOC_428/Y VSS VDD INVX1_LOC_118/A
+ INVX1_LOC_22/A NOR2X1_LOC
XNOR2X1_LOC_417 NOR2X1_LOC_417/a_36_216# INVX1_LOC_178/A VSS VDD NOR2X1_LOC_226/A
+ INVX1_LOC_36/A NOR2X1_LOC
XNOR2X1_LOC_439 NOR2X1_LOC_439/a_36_216# INVX1_LOC_182/A VSS VDD NOR2X1_LOC_544/A
+ NOR2X1_LOC_439/B NOR2X1_LOC
XNOR2X1_LOC_406 NOR2X1_LOC_406/a_36_216# INVX1_LOC_172/A VSS VDD NOR2X1_LOC_406/A
+ INVX1_LOC_58/A NOR2X1_LOC
XNOR2X1_LOC_258 NOR2X1_LOC_258/a_36_216# NOR2X1_LOC_258/Y VSS VDD INVX1_LOC_90/A NOR2X1_LOC_89/A
+ NOR2X1_LOC
XNOR2X1_LOC_214 NOR2X1_LOC_214/a_36_216# NOR2X1_LOC_219/B VSS VDD NOR2X1_LOC_208/Y
+ NOR2X1_LOC_214/B NOR2X1_LOC
XNOR2X1_LOC_269 NOR2X1_LOC_269/a_36_216# NOR2X1_LOC_269/Y VSS VDD INVX1_LOC_128/Y
+ INVX1_LOC_118/Y NOR2X1_LOC
XNOR2X1_LOC_203 NOR2X1_LOC_203/a_36_216# NOR2X1_LOC_203/Y VSS VDD INVX1_LOC_55/Y NAND2X1_LOC_72/Y
+ NOR2X1_LOC
XNOR2X1_LOC_225 NOR2X1_LOC_225/a_36_216# NOR2X1_LOC_226/A VSS VDD INVX1_LOC_4/A INPUT_1
+ NOR2X1_LOC
XNOR2X1_LOC_247 NOR2X1_LOC_247/a_36_216# NOR2X1_LOC_247/Y VSS VDD INVX1_LOC_9/A INVX1_LOC_5/A
+ NOR2X1_LOC
XNOR2X1_LOC_236 NOR2X1_LOC_236/a_36_216# INVX1_LOC_118/A VSS VDD NOR2X1_LOC_38/B INVX1_LOC_3/Y
+ NOR2X1_LOC
XNAND2X1_LOC_748 NAND2X1_LOC_748/a_36_24# NOR2X1_LOC_789/B VSS VDD NOR2X1_LOC_19/B
+ NOR2X1_LOC_709/A NAND2X1_LOC
XNAND2X1_LOC_726 NAND2X1_LOC_726/a_36_24# NAND2X1_LOC_726/Y VSS VDD NOR2X1_LOC_152/Y
+ NAND2X1_LOC_711/Y NAND2X1_LOC
XNAND2X1_LOC_759 NAND2X1_LOC_759/a_36_24# NOR2X1_LOC_792/B VSS VDD INVX1_LOC_118/Y
+ NOR2X1_LOC_758/Y NAND2X1_LOC
XNAND2X1_LOC_715 NAND2X1_LOC_715/a_36_24# INVX1_LOC_279/A VSS VDD NAND2X1_LOC_112/Y
+ NAND2X1_LOC_715/B NAND2X1_LOC
XNAND2X1_LOC_704 NAND2X1_LOC_704/a_36_24# NAND2X1_LOC_714/B VSS VDD NOR2X1_LOC_313/Y
+ INVX1_LOC_178/A NAND2X1_LOC
XNAND2X1_LOC_737 NAND2X1_LOC_737/a_36_24# NAND2X1_LOC_741/B VSS VDD NAND2X1_LOC_733/Y
+ INVX1_LOC_286/Y NAND2X1_LOC
XNOR2X1_LOC_770 NOR2X1_LOC_770/a_36_216# NOR2X1_LOC_770/Y VSS VDD NOR2X1_LOC_770/A
+ NOR2X1_LOC_770/B NOR2X1_LOC
XNOR2X1_LOC_781 NOR2X1_LOC_781/a_36_216# NOR2X1_LOC_781/Y VSS VDD NOR2X1_LOC_781/A
+ NOR2X1_LOC_781/B NOR2X1_LOC
XNOR2X1_LOC_792 NOR2X1_LOC_792/a_36_216# INVX1_LOC_308/A VSS VDD NOR2X1_LOC_791/Y
+ NOR2X1_LOC_792/B NOR2X1_LOC
XNAND2X1_LOC_501 NAND2X1_LOC_501/a_36_24# INVX1_LOC_207/A VSS VDD NOR2X1_LOC_498/Y
+ NAND2X1_LOC_500/Y NAND2X1_LOC
XNAND2X1_LOC_556 NAND2X1_LOC_556/a_36_24# NAND2X1_LOC_562/B VSS VDD NAND2X1_LOC_483/Y
+ NAND2X1_LOC_787/B NAND2X1_LOC
XNAND2X1_LOC_523 NAND2X1_LOC_523/a_36_24# NAND2X1_LOC_560/A VSS VDD NOR2X1_LOC_521/Y
+ NOR2X1_LOC_522/Y NAND2X1_LOC
XNAND2X1_LOC_578 NAND2X1_LOC_578/a_36_24# INVX1_LOC_239/A VSS VDD INVX1_LOC_232/Y
+ NAND2X1_LOC_578/B NAND2X1_LOC
XNAND2X1_LOC_545 NAND2X1_LOC_545/a_36_24# INVX1_LOC_223/A VSS VDD NOR2X1_LOC_441/Y
+ NOR2X1_LOC_524/Y NAND2X1_LOC
XNAND2X1_LOC_534 NAND2X1_LOC_534/a_36_24# INVX1_LOC_221/A VSS VDD INVX1_LOC_31/A INVX1_LOC_45/A
+ NAND2X1_LOC
XNAND2X1_LOC_567 NAND2X1_LOC_567/a_36_24# NAND2X1_LOC_567/Y VSS VDD NAND2X1_LOC_854/B
+ NAND2X1_LOC_799/A NAND2X1_LOC
XNAND2X1_LOC_512 NAND2X1_LOC_512/a_36_24# NAND2X1_LOC_513/B VSS VDD INPUT_0 INVX1_LOC_142/A
+ NAND2X1_LOC
XNAND2X1_LOC_589 NAND2X1_LOC_589/a_36_24# NOR2X1_LOC_592/A VSS VDD INVX1_LOC_17/A
+ NOR2X1_LOC_130/A NAND2X1_LOC
XNAND2X1_LOC_320 NAND2X1_LOC_320/a_36_24# NOR2X1_LOC_324/B VSS VDD INVX1_LOC_23/A
+ NOR2X1_LOC_383/B NAND2X1_LOC
XNAND2X1_LOC_364 NAND2X1_LOC_364/a_36_24# NAND2X1_LOC_364/Y VSS VDD NAND2X1_LOC_364/A
+ NAND2X1_LOC_358/Y NAND2X1_LOC
XNAND2X1_LOC_397 NAND2X1_LOC_397/a_36_24# INVX1_LOC_163/A VSS VDD INVX1_LOC_1/A NAND2X1_LOC_82/Y
+ NAND2X1_LOC
XNAND2X1_LOC_342 NAND2X1_LOC_342/a_36_24# NAND2X1_LOC_342/Y VSS VDD NOR2X1_LOC_246/Y
+ NOR2X1_LOC_248/Y NAND2X1_LOC
XNAND2X1_LOC_353 NAND2X1_LOC_353/a_36_24# NAND2X1_LOC_357/B VSS VDD NAND2X1_LOC_303/Y
+ NAND2X1_LOC_308/Y NAND2X1_LOC
XNAND2X1_LOC_331 NAND2X1_LOC_331/a_36_24# NOR2X1_LOC_355/A VSS VDD NOR2X1_LOC_186/Y
+ INVX1_LOC_145/Y NAND2X1_LOC
XNAND2X1_LOC_375 NAND2X1_LOC_375/a_36_24# NOR2X1_LOC_376/A VSS VDD INVX1_LOC_22/A
+ INVX1_LOC_90/A NAND2X1_LOC
XNAND2X1_LOC_386 NAND2X1_LOC_386/a_36_24# NAND2X1_LOC_387/B VSS VDD D_INPUT_4
+ NAND2X1_LOC_36/A NAND2X1_LOC
XINVX1_LOC_219 INVX1_LOC_219/Y VSS VDD INVX1_LOC_219/A INVX1_LOC
XINVX1_LOC_208 INVX1_LOC_208/Y VSS VDD INVX1_LOC_208/A INVX1_LOC
XNAND2X1_LOC_150 NAND2X1_LOC_150/a_36_24# INVX1_LOC_87/A VSS VDD INVX1_LOC_26/Y INVX1_LOC_47/A
+ NAND2X1_LOC
XNAND2X1_LOC_19 NAND2X1_LOC_19/a_36_24# NAND2X1_LOC_20/B VSS VDD NOR2X1_LOC_6/B INVX1_LOC_3/A
+ NAND2X1_LOC
XNAND2X1_LOC_161 NAND2X1_LOC_161/a_36_24# NAND2X1_LOC_162/B VSS VDD INVX1_LOC_78/A
+ INVX1_LOC_92/A NAND2X1_LOC
XNAND2X1_LOC_194 NAND2X1_LOC_194/a_36_24# NAND2X1_LOC_200/B VSS VDD NOR2X1_LOC_16/Y
+ NOR2X1_LOC_39/Y NAND2X1_LOC
XNAND2X1_LOC_172 NAND2X1_LOC_172/a_36_24# NOR2X1_LOC_174/A VSS VDD INVX1_LOC_53/A
+ NOR2X1_LOC_590/A NAND2X1_LOC
XNAND2X1_LOC_183 NAND2X1_LOC_183/a_36_24# INVX1_LOC_97/A VSS VDD INVX1_LOC_5/A INVX1_LOC_29/A
+ NAND2X1_LOC
XNOR2X1_LOC_429 NOR2X1_LOC_429/a_36_216# NOR2X1_LOC_430/A VSS VDD NOR2X1_LOC_11/Y
+ INPUT_7 NOR2X1_LOC
XNOR2X1_LOC_418 NOR2X1_LOC_418/a_36_216# NOR2X1_LOC_418/Y VSS VDD INVX1_LOC_38/A NOR2X1_LOC_15/Y
+ NOR2X1_LOC
XNOR2X1_LOC_407 NOR2X1_LOC_407/a_36_216# NOR2X1_LOC_828/B VSS VDD NOR2X1_LOC_155/A
+ INVX1_LOC_41/A NOR2X1_LOC
XNOR2X1_LOC_215 NOR2X1_LOC_215/a_36_216# NOR2X1_LOC_215/Y VSS VDD NOR2X1_LOC_215/A
+ NOR2X1_LOC_205/Y NOR2X1_LOC
XNOR2X1_LOC_204 NOR2X1_LOC_204/a_36_216# INVX1_LOC_112/A VSS VDD NOR2X1_LOC_84/Y NAND2X1_LOC_79/Y
+ NOR2X1_LOC
XNOR2X1_LOC_226 NOR2X1_LOC_226/a_36_216# NOR2X1_LOC_226/Y VSS VDD NOR2X1_LOC_226/A
+ INVX1_LOC_16/A NOR2X1_LOC
XNOR2X1_LOC_248 NOR2X1_LOC_248/a_36_216# NOR2X1_LOC_248/Y VSS VDD NOR2X1_LOC_248/A
+ INVX1_LOC_36/A NOR2X1_LOC
XNOR2X1_LOC_259 NOR2X1_LOC_259/a_36_216# INVX1_LOC_122/A VSS VDD NOR2X1_LOC_259/A
+ NOR2X1_LOC_259/B NOR2X1_LOC
XNOR2X1_LOC_237 NOR2X1_LOC_237/a_36_216# NOR2X1_LOC_237/Y VSS VDD INVX1_LOC_118/A
+ INVX1_LOC_20/A NOR2X1_LOC
XNAND2X1_LOC_705 NAND2X1_LOC_705/a_36_24# NAND2X1_LOC_705/Y VSS VDD NOR2X1_LOC_485/Y
+ NOR2X1_LOC_526/Y NAND2X1_LOC
XNAND2X1_LOC_749 NAND2X1_LOC_749/a_36_24# NOR2X1_LOC_750/A VSS VDD D_INPUT_0 INVX1_LOC_7/A
+ NAND2X1_LOC
XNAND2X1_LOC_727 NAND2X1_LOC_727/a_36_24# NAND2X1_LOC_727/Y VSS VDD NAND2X1_LOC_308/Y
+ INVX1_LOC_185/A NAND2X1_LOC
XNAND2X1_LOC_738 NAND2X1_LOC_738/a_36_24# NAND2X1_LOC_740/A VSS VDD NAND2X1_LOC_731/Y
+ NAND2X1_LOC_738/B NAND2X1_LOC
XNAND2X1_LOC_716 NAND2X1_LOC_716/a_36_24# INVX1_LOC_281/A VSS VDD NAND2X1_LOC_341/A
+ INVX1_LOC_139/A NAND2X1_LOC
XNOR2X1_LOC_771 NOR2X1_LOC_771/a_36_216# INVX1_LOC_298/A VSS VDD NOR2X1_LOC_770/Y
+ INVX1_LOC_295/Y NOR2X1_LOC
XNOR2X1_LOC_760 NOR2X1_LOC_760/a_36_216# INVX1_LOC_292/A VSS VDD NOR2X1_LOC_329/B
+ INVX1_LOC_50/A NOR2X1_LOC
XNOR2X1_LOC_782 NOR2X1_LOC_782/a_36_216# INVX1_LOC_302/A VSS VDD NOR2X1_LOC_781/Y
+ INVX1_LOC_288/Y NOR2X1_LOC
XNOR2X1_LOC_793 NOR2X1_LOC_793/a_36_216# NOR2X1_LOC_793/Y VSS VDD NOR2X1_LOC_793/A
+ INVX1_LOC_305/Y NOR2X1_LOC
XNAND2X1_LOC_502 NAND2X1_LOC_502/a_36_24# NOR2X1_LOC_503/A VSS VDD NOR2X1_LOC_89/A
+ INVX1_LOC_84/A NAND2X1_LOC
XNAND2X1_LOC_546 NAND2X1_LOC_546/a_36_24# NAND2X1_LOC_550/A VSS VDD NOR2X1_LOC_525/Y
+ NOR2X1_LOC_526/Y NAND2X1_LOC
XNAND2X1_LOC_524 NAND2X1_LOC_524/a_36_24# NOR2X1_LOC_545/A VSS VDD INVX1_LOC_35/A
+ INVX1_LOC_77/A NAND2X1_LOC
XNAND2X1_LOC_579 NAND2X1_LOC_579/a_36_24# INVX1_LOC_241/A VSS VDD NAND2X1_LOC_579/A
+ INVX1_LOC_238/Y NAND2X1_LOC
XNAND2X1_LOC_557 NAND2X1_LOC_557/a_36_24# NAND2X1_LOC_557/Y VSS VDD NAND2X1_LOC_489/Y
+ NOR2X1_LOC_490/Y NAND2X1_LOC
XNAND2X1_LOC_535 NAND2X1_LOC_535/a_36_24# NAND2X1_LOC_854/B VSS VDD NOR2X1_LOC_533/Y
+ INVX1_LOC_221/Y NAND2X1_LOC
XNAND2X1_LOC_568 NAND2X1_LOC_568/a_36_24# INVX1_LOC_231/A VSS VDD NAND2X1_LOC_568/A
+ NAND2X1_LOC_567/Y NAND2X1_LOC
XNAND2X1_LOC_513 NAND2X1_LOC_513/a_36_24# NOR2X1_LOC_516/B VSS VDD INVX1_LOC_213/Y
+ NAND2X1_LOC_513/B NAND2X1_LOC
XNOR2X1_LOC_590 NOR2X1_LOC_590/a_36_216# NOR2X1_LOC_590/Y VSS VDD NOR2X1_LOC_590/A
+ INVX1_LOC_27/A NOR2X1_LOC
XNAND2X1_LOC_321 NAND2X1_LOC_321/a_36_24# NOR2X1_LOC_324/A VSS VDD INVX1_LOC_9/A INVX1_LOC_49/A
+ NAND2X1_LOC
XNAND2X1_LOC_310 NAND2X1_LOC_310/a_36_24# NOR2X1_LOC_335/A VSS VDD INVX1_LOC_4/Y INVX1_LOC_29/A
+ NAND2X1_LOC
XNAND2X1_LOC_343 NAND2X1_LOC_343/a_36_24# NAND2X1_LOC_349/B VSS VDD NOR2X1_LOC_250/Y
+ NOR2X1_LOC_251/Y NAND2X1_LOC
XNAND2X1_LOC_332 NAND2X1_LOC_332/a_36_24# NAND2X1_LOC_332/Y VSS VDD NOR2X1_LOC_111/Y
+ NOR2X1_LOC_135/Y NAND2X1_LOC
XNAND2X1_LOC_354 NAND2X1_LOC_354/a_36_24# NAND2X1_LOC_354/Y VSS VDD NAND2X1_LOC_798/A
+ NAND2X1_LOC_354/B NAND2X1_LOC
XNAND2X1_LOC_365 NAND2X1_LOC_365/a_36_24# NAND2X1_LOC_367/A VSS VDD INVX1_LOC_160/Y
+ NAND2X1_LOC_364/Y NAND2X1_LOC
XNAND2X1_LOC_376 NAND2X1_LOC_376/a_36_24# NOR2X1_LOC_459/B VSS VDD INVX1_LOC_84/Y
+ NOR2X1_LOC_375/Y NAND2X1_LOC
XNAND2X1_LOC_398 NAND2X1_LOC_398/a_36_24# NOR2X1_LOC_399/A VSS VDD NOR2X1_LOC_15/Y
+ INVX1_LOC_135/Y NAND2X1_LOC
XNAND2X1_LOC_387 NAND2X1_LOC_387/a_36_24# NOR2X1_LOC_389/A VSS VDD NAND2X1_LOC_93/B
+ NAND2X1_LOC_387/B NAND2X1_LOC
XINVX1_LOC_209 INVX1_LOC_209/Y VSS VDD INVX1_LOC_209/A INVX1_LOC
XNAND2X1_LOC_173 NAND2X1_LOC_173/a_36_24# NOR2X1_LOC_175/B VSS VDD INVX1_LOC_54/Y
+ INVX1_LOC_87/A NAND2X1_LOC
XNAND2X1_LOC_184 NAND2X1_LOC_184/a_36_24# INVX1_LOC_99/A VSS VDD NAND2X1_LOC_72/B
+ INVX1_LOC_58/Y NAND2X1_LOC
XNAND2X1_LOC_151 NAND2X1_LOC_151/a_36_24# NOR2X1_LOC_152/A VSS VDD INVX1_LOC_42/A
+ INVX1_LOC_88/A NAND2X1_LOC
XNAND2X1_LOC_140 NAND2X1_LOC_140/a_36_24# INVX1_LOC_81/A VSS VDD NAND2X1_LOC_140/A
+ NOR2X1_LOC_131/Y NAND2X1_LOC
XNAND2X1_LOC_195 NAND2X1_LOC_195/a_36_24# NAND2X1_LOC_195/Y VSS VDD NOR2X1_LOC_41/Y
+ NOR2X1_LOC_43/Y NAND2X1_LOC
XNAND2X1_LOC_162 NAND2X1_LOC_162/a_36_24# NOR2X1_LOC_163/A VSS VDD NAND2X1_LOC_162/A
+ NAND2X1_LOC_162/B NAND2X1_LOC
XNOR2X1_LOC_408 NOR2X1_LOC_408/a_36_216# INVX1_LOC_174/A VSS VDD NOR2X1_LOC_36/A INPUT_6
+ NOR2X1_LOC
XNOR2X1_LOC_419 NOR2X1_LOC_419/a_36_216# NOR2X1_LOC_419/Y VSS VDD INVX1_LOC_32/A INVX1_LOC_24/A
+ NOR2X1_LOC
XNOR2X1_LOC_205 NOR2X1_LOC_205/a_36_216# NOR2X1_LOC_205/Y VSS VDD INVX1_LOC_111/Y
+ NOR2X1_LOC_203/Y NOR2X1_LOC
XNOR2X1_LOC_216 NOR2X1_LOC_216/a_36_216# NOR2X1_LOC_216/Y VSS VDD NOR2X1_LOC_473/B
+ NOR2X1_LOC_216/B NOR2X1_LOC
XNOR2X1_LOC_227 NOR2X1_LOC_227/a_36_216# NOR2X1_LOC_340/A VSS VDD NOR2X1_LOC_227/A
+ NOR2X1_LOC_227/B NOR2X1_LOC
XNOR2X1_LOC_249 NOR2X1_LOC_249/a_36_216# NOR2X1_LOC_249/Y VSS VDD INVX1_LOC_27/A NOR2X1_LOC_160/B
+ NOR2X1_LOC
XNOR2X1_LOC_238 NOR2X1_LOC_238/a_36_216# NOR2X1_LOC_238/Y VSS VDD INVX1_LOC_37/Y NOR2X1_LOC_45/B
+ NOR2X1_LOC
XNAND2X1_LOC_706 NAND2X1_LOC_706/a_36_24# NAND2X1_LOC_706/Y VSS VDD NOR2X1_LOC_692/Y
+ NOR2X1_LOC_693/Y NAND2X1_LOC
XNAND2X1_LOC_717 NAND2X1_LOC_717/a_36_24# NAND2X1_LOC_717/Y VSS VDD NAND2X1_LOC_374/Y
+ NAND2X1_LOC_493/Y NAND2X1_LOC
XNAND2X1_LOC_728 NAND2X1_LOC_728/a_36_24# NAND2X1_LOC_728/Y VSS VDD NOR2X1_LOC_679/Y
+ INVX1_LOC_273/Y NAND2X1_LOC
XNAND2X1_LOC_739 NAND2X1_LOC_739/a_36_24# NAND2X1_LOC_740/B VSS VDD INVX1_LOC_103/A
+ NAND2X1_LOC_739/B NAND2X1_LOC
XNOR2X1_LOC_783 NOR2X1_LOC_783/a_36_216# NOR2X1_LOC_796/B VSS VDD NOR2X1_LOC_783/A
+ NOR2X1_LOC_779/Y NOR2X1_LOC
XNOR2X1_LOC_761 NOR2X1_LOC_761/a_36_216# NOR2X1_LOC_761/Y VSS VDD NOR2X1_LOC_599/Y
+ INPUT_0 NOR2X1_LOC
XNOR2X1_LOC_794 NOR2X1_LOC_794/a_36_216# NOR2X1_LOC_804/B VSS VDD NOR2X1_LOC_794/A
+ NOR2X1_LOC_794/B NOR2X1_LOC
XNOR2X1_LOC_772 NOR2X1_LOC_772/a_36_216# NOR2X1_LOC_772/Y VSS VDD NOR2X1_LOC_772/A
+ NOR2X1_LOC_772/B NOR2X1_LOC
XNOR2X1_LOC_750 NOR2X1_LOC_750/a_36_216# NOR2X1_LOC_750/Y VSS VDD NOR2X1_LOC_750/A
+ INVX1_LOC_91/A NOR2X1_LOC
XNAND2X1_LOC_503 NAND2X1_LOC_503/a_36_24# NOR2X1_LOC_509/A VSS VDD INVX1_LOC_50/Y
+ NOR2X1_LOC_502/Y NAND2X1_LOC
XNAND2X1_LOC_536 NAND2X1_LOC_536/a_36_24# NOR2X1_LOC_537/A VSS VDD INVX1_LOC_11/A
+ NOR2X1_LOC_590/A NAND2X1_LOC
XNAND2X1_LOC_514 NAND2X1_LOC_514/a_36_24# NAND2X1_LOC_514/Y VSS VDD D_INPUT_0
+ NOR2X1_LOC_136/Y NAND2X1_LOC
XNAND2X1_LOC_525 NAND2X1_LOC_525/a_36_24# NOR2X1_LOC_546/B VSS VDD INVX1_LOC_9/A INVX1_LOC_37/A
+ NAND2X1_LOC
XNAND2X1_LOC_558 NAND2X1_LOC_558/a_36_24# NAND2X1_LOC_561/B VSS VDD NAND2X1_LOC_493/Y
+ NOR2X1_LOC_494/Y NAND2X1_LOC
XNAND2X1_LOC_569 NAND2X1_LOC_569/a_36_24# NAND2X1_LOC_577/A VSS VDD NAND2X1_LOC_569/A
+ NAND2X1_LOC_569/B NAND2X1_LOC
XNAND2X1_LOC_547 NAND2X1_LOC_547/a_36_24# INVX1_LOC_225/A VSS VDD NOR2X1_LOC_527/Y
+ NOR2X1_LOC_528/Y NAND2X1_LOC
XNOR2X1_LOC_591 NOR2X1_LOC_591/a_36_216# NOR2X1_LOC_591/Y VSS VDD NOR2X1_LOC_591/A
+ INVX1_LOC_49/Y NOR2X1_LOC
XNOR2X1_LOC_580 NOR2X1_LOC_580/a_36_216# D_GATE_579 VSS VDD INVX1_LOC_241/Y INVX1_LOC_239/Y
+ NOR2X1_LOC
XNAND2X1_LOC_366 NAND2X1_LOC_366/a_36_24# NAND2X1_LOC_367/B VSS VDD NAND2X1_LOC_366/A
+ NAND2X1_LOC_363/Y NAND2X1_LOC
XNAND2X1_LOC_344 NAND2X1_LOC_344/a_36_24# NAND2X1_LOC_348/A VSS VDD NAND2X1_LOC_254/Y
+ NOR2X1_LOC_256/Y NAND2X1_LOC
XNAND2X1_LOC_377 NAND2X1_LOC_377/a_36_24# NAND2X1_LOC_377/Y VSS VDD INVX1_LOC_1/A
+ INVX1_LOC_14/A NAND2X1_LOC
XNAND2X1_LOC_311 NAND2X1_LOC_311/a_36_24# NOR2X1_LOC_336/B VSS VDD INVX1_LOC_19/A
+ NOR2X1_LOC_590/A NAND2X1_LOC
XNAND2X1_LOC_300 NAND2X1_LOC_300/a_36_24# NOR2X1_LOC_301/A VSS VDD INVX1_LOC_45/A
+ INVX1_LOC_71/A NAND2X1_LOC
XNAND2X1_LOC_322 NAND2X1_LOC_322/a_36_24# NOR2X1_LOC_374/B VSS VDD INVX1_LOC_33/A
+ INVX1_LOC_83/A NAND2X1_LOC
XNAND2X1_LOC_333 NAND2X1_LOC_333/a_36_24# INVX1_LOC_147/A VSS VDD NOR2X1_LOC_171/Y
+ NOR2X1_LOC_289/Y NAND2X1_LOC
XNAND2X1_LOC_355 NAND2X1_LOC_355/a_36_24# NAND2X1_LOC_355/Y VSS VDD NOR2X1_LOC_329/Y
+ NOR2X1_LOC_331/Y NAND2X1_LOC
XNAND2X1_LOC_399 NAND2X1_LOC_399/a_36_24# NOR2X1_LOC_403/B VSS VDD INVX1_LOC_34/Y
+ NOR2X1_LOC_398/Y NAND2X1_LOC
XNAND2X1_LOC_388 NAND2X1_LOC_388/a_36_24# NAND2X1_LOC_390/A VSS VDD NOR2X1_LOC_167/Y
+ NOR2X1_LOC_176/Y NAND2X1_LOC
XNAND2X1_LOC_141 NAND2X1_LOC_141/a_36_24# NAND2X1_LOC_141/Y VSS VDD NAND2X1_LOC_141/A
+ INVX1_LOC_82/Y NAND2X1_LOC
XNAND2X1_LOC_185 NAND2X1_LOC_185/a_36_24# NOR2X1_LOC_816/A VSS VDD INVX1_LOC_41/Y
+ NOR2X1_LOC_74/A NAND2X1_LOC
XNAND2X1_LOC_174 NAND2X1_LOC_174/a_36_24# NAND2X1_LOC_175/B VSS VDD NOR2X1_LOC_171/Y
+ NOR2X1_LOC_172/Y NAND2X1_LOC
XNAND2X1_LOC_130 NAND2X1_LOC_130/a_36_24# NOR2X1_LOC_131/A VSS VDD INVX1_LOC_6/A NOR2X1_LOC_589/A
+ NAND2X1_LOC
XNAND2X1_LOC_152 NAND2X1_LOC_152/a_36_24# NOR2X1_LOC_209/A VSS VDD INVX1_LOC_35/A
+ NOR2X1_LOC_151/Y NAND2X1_LOC
XNAND2X1_LOC_196 NAND2X1_LOC_196/a_36_24# NAND2X1_LOC_199/B VSS VDD NOR2X1_LOC_45/Y
+ NOR2X1_LOC_48/Y NAND2X1_LOC
XNAND2X1_LOC_163 NAND2X1_LOC_163/a_36_24# NOR2X1_LOC_210/A VSS VDD INVX1_LOC_37/A
+ NOR2X1_LOC_162/Y NAND2X1_LOC
XNOR2X1_LOC_409 NOR2X1_LOC_409/a_36_216# NOR2X1_LOC_409/Y VSS VDD INVX1_LOC_173/Y
+ NOR2X1_LOC_409/B NOR2X1_LOC
XNOR2X1_LOC_206 NOR2X1_LOC_206/a_36_216# NOR2X1_LOC_215/A VSS VDD NOR2X1_LOC_202/Y
+ INVX1_LOC_109/Y NOR2X1_LOC
XNOR2X1_LOC_217 NOR2X1_LOC_217/a_36_216# NOR2X1_LOC_218/A VSS VDD NOR2X1_LOC_657/B
+ INVX1_LOC_73/Y NOR2X1_LOC
XNOR2X1_LOC_239 NOR2X1_LOC_239/a_36_216# INVX1_LOC_120/A VSS VDD NOR2X1_LOC_536/A
+ INVX1_LOC_38/A NOR2X1_LOC
XNOR2X1_LOC_228 NOR2X1_LOC_228/a_36_216# NOR2X1_LOC_716/B VSS VDD NOR2X1_LOC_197/B
+ NAND2X1_LOC_7/Y NOR2X1_LOC
XNAND2X1_LOC_718 NAND2X1_LOC_718/a_36_24# NAND2X1_LOC_722/A VSS VDD NOR2X1_LOC_591/Y
+ INVX1_LOC_250/Y NAND2X1_LOC
XNAND2X1_LOC_707 NAND2X1_LOC_707/a_36_24# NAND2X1_LOC_712/A VSS VDD NOR2X1_LOC_694/Y
+ NOR2X1_LOC_695/Y NAND2X1_LOC
XNAND2X1_LOC_729 NAND2X1_LOC_729/a_36_24# NAND2X1_LOC_729/Y VSS VDD NAND2X1_LOC_800/A
+ NAND2X1_LOC_729/B NAND2X1_LOC
XNOR2X1_LOC_762 NOR2X1_LOC_762/a_36_216# NOR2X1_LOC_763/A VSS VDD NOR2X1_LOC_11/Y
+ D_INPUT_6 NOR2X1_LOC
XNOR2X1_LOC_740 NOR2X1_LOC_740/a_36_216# NOR2X1_LOC_740/Y VSS VDD NOR2X1_LOC_739/Y
+ NOR2X1_LOC_738/Y NOR2X1_LOC
XNOR2X1_LOC_784 NOR2X1_LOC_784/a_36_216# NOR2X1_LOC_784/Y VSS VDD NOR2X1_LOC_778/Y
+ NOR2X1_LOC_784/B NOR2X1_LOC
XNOR2X1_LOC_773 NOR2X1_LOC_773/a_36_216# NOR2X1_LOC_773/Y VSS VDD NOR2X1_LOC_772/Y
+ INVX1_LOC_294/Y NOR2X1_LOC
XNOR2X1_LOC_795 NOR2X1_LOC_795/a_36_216# NOR2X1_LOC_795/Y VSS VDD INVX1_LOC_303/Y
+ NOR2X1_LOC_785/Y NOR2X1_LOC
XNOR2X1_LOC_751 NOR2X1_LOC_751/a_36_216# NOR2X1_LOC_751/Y VSS VDD NOR2X1_LOC_751/A
+ INVX1_LOC_1/Y NOR2X1_LOC
XNAND2X1_LOC_559 NAND2X1_LOC_559/a_36_24# NAND2X1_LOC_559/Y VSS VDD NOR2X1_LOC_517/Y
+ INVX1_LOC_217/A NAND2X1_LOC
XNAND2X1_LOC_548 NAND2X1_LOC_548/a_36_24# NAND2X1_LOC_549/B VSS VDD NOR2X1_LOC_529/Y
+ NOR2X1_LOC_530/Y NAND2X1_LOC
XNAND2X1_LOC_504 NAND2X1_LOC_504/a_36_24# NOR2X1_LOC_507/B VSS VDD INVX1_LOC_9/A INVX1_LOC_89/A
+ NAND2X1_LOC
XNAND2X1_LOC_537 NAND2X1_LOC_537/a_36_24# NAND2X1_LOC_537/Y VSS VDD NOR2X1_LOC_385/Y
+ NOR2X1_LOC_536/Y NAND2X1_LOC
XNAND2X1_LOC_515 NAND2X1_LOC_515/a_36_24# INVX1_LOC_215/A VSS VDD INVX1_LOC_177/Y
+ NAND2X1_LOC_514/Y NAND2X1_LOC
XNAND2X1_LOC_526 NAND2X1_LOC_526/a_36_24# NOR2X1_LOC_546/A VSS VDD INVX1_LOC_21/A
+ INVX1_LOC_91/A NAND2X1_LOC
XINVX1_LOC_190 INVX1_LOC_190/Y VSS VDD INVX1_LOC_190/A INVX1_LOC
XNOR2X1_LOC_581 NOR2X1_LOC_581/a_36_216# NOR2X1_LOC_582/A VSS VDD NOR2X1_LOC_2/Y D_INPUT_6
+ NOR2X1_LOC
XNOR2X1_LOC_592 NOR2X1_LOC_592/a_36_216# INVX1_LOC_246/A VSS VDD NOR2X1_LOC_592/A
+ NOR2X1_LOC_592/B NOR2X1_LOC
XNOR2X1_LOC_570 NOR2X1_LOC_570/a_36_216# NOR2X1_LOC_570/Y VSS VDD NOR2X1_LOC_570/A
+ NOR2X1_LOC_570/B NOR2X1_LOC
XNAND2X1_LOC_367 NAND2X1_LOC_367/a_36_24# GATE_366 VSS VDD NAND2X1_LOC_367/A NAND2X1_LOC_367/B
+ NAND2X1_LOC
XNAND2X1_LOC_334 NAND2X1_LOC_334/a_36_24# NAND2X1_LOC_338/B VSS VDD NOR2X1_LOC_290/Y
+ NOR2X1_LOC_291/Y NAND2X1_LOC
XNAND2X1_LOC_378 NAND2X1_LOC_378/a_36_24# NOR2X1_LOC_459/A VSS VDD INVX1_LOC_32/A
+ NAND2X1_LOC_377/Y NAND2X1_LOC
XNAND2X1_LOC_323 NAND2X1_LOC_323/a_36_24# NOR2X1_LOC_325/A VSS VDD INVX1_LOC_57/A
+ NAND2X1_LOC_323/B NAND2X1_LOC
XNAND2X1_LOC_312 NAND2X1_LOC_312/a_36_24# NOR2X1_LOC_703/A VSS VDD INVX1_LOC_41/A
+ INVX1_LOC_49/A NAND2X1_LOC
XNAND2X1_LOC_389 NAND2X1_LOC_389/a_36_24# INVX1_LOC_161/A VSS VDD NOR2X1_LOC_385/Y
+ NOR2X1_LOC_387/Y NAND2X1_LOC
XNAND2X1_LOC_356 NAND2X1_LOC_356/a_36_24# INVX1_LOC_159/A VSS VDD NAND2X1_LOC_354/Y
+ NAND2X1_LOC_355/Y NAND2X1_LOC
XNAND2X1_LOC_301 NAND2X1_LOC_301/a_36_24# INVX1_LOC_139/A VSS VDD NOR2X1_LOC_75/Y
+ NOR2X1_LOC_300/Y NAND2X1_LOC
XNAND2X1_LOC_345 NAND2X1_LOC_345/a_36_24# INVX1_LOC_153/A VSS VDD INVX1_LOC_121/A
+ NOR2X1_LOC_261/Y NAND2X1_LOC
XNAND2X1_LOC_131 NAND2X1_LOC_131/a_36_24# NOR2X1_LOC_140/A VSS VDD INVX1_LOC_12/Y
+ NOR2X1_LOC_130/Y NAND2X1_LOC
XNAND2X1_LOC_153 NAND2X1_LOC_153/a_36_24# NOR2X1_LOC_155/A VSS VDD D_INPUT_1 INVX1_LOC_25/A
+ NAND2X1_LOC
XNAND2X1_LOC_164 NAND2X1_LOC_164/a_36_24# NOR2X1_LOC_168/B VSS VDD INVX1_LOC_15/A
+ INVX1_LOC_83/A NAND2X1_LOC
XNAND2X1_LOC_186 NAND2X1_LOC_186/a_36_24# NOR2X1_LOC_331/B VSS VDD INVX1_LOC_88/A
+ NOR2X1_LOC_816/A NAND2X1_LOC
XNAND2X1_LOC_175 NAND2X1_LOC_175/a_36_24# NAND2X1_LOC_175/Y VSS VDD NOR2X1_LOC_173/Y
+ NAND2X1_LOC_175/B NAND2X1_LOC
XNAND2X1_LOC_120 NAND2X1_LOC_120/a_36_24# NOR2X1_LOC_666/A VSS VDD INVX1_LOC_10/A
+ INVX1_LOC_28/A NAND2X1_LOC
XNAND2X1_LOC_197 NAND2X1_LOC_197/a_36_24# NAND2X1_LOC_198/B VSS VDD NOR2X1_LOC_52/Y
+ NOR2X1_LOC_56/Y NAND2X1_LOC
XNAND2X1_LOC_142 NAND2X1_LOC_142/a_36_24# NOR2X1_LOC_147/B VSS VDD NOR2X1_LOC_68/A
+ INVX1_LOC_49/A NAND2X1_LOC
XNOR2X1_LOC_229 NOR2X1_LOC_229/a_36_216# NOR2X1_LOC_229/Y VSS VDD NOR2X1_LOC_45/B
+ INVX1_LOC_12/A NOR2X1_LOC
XNOR2X1_LOC_207 NOR2X1_LOC_207/a_36_216# NOR2X1_LOC_214/B VSS VDD NOR2X1_LOC_207/A
+ INVX1_LOC_107/Y NOR2X1_LOC
XNOR2X1_LOC_218 NOR2X1_LOC_218/a_36_216# NOR2X1_LOC_218/Y VSS VDD NOR2X1_LOC_218/A
+ NOR2X1_LOC_216/Y NOR2X1_LOC
XNAND2X1_LOC_719 NAND2X1_LOC_719/a_36_24# INVX1_LOC_283/A VSS VDD NOR2X1_LOC_665/Y
+ NOR2X1_LOC_666/Y NAND2X1_LOC
XNAND2X1_LOC_708 NAND2X1_LOC_708/a_36_24# NAND2X1_LOC_708/Y VSS VDD NOR2X1_LOC_696/Y
+ NOR2X1_LOC_697/Y NAND2X1_LOC
XNOR2X1_LOC_763 NOR2X1_LOC_763/a_36_216# NOR2X1_LOC_763/Y VSS VDD NOR2X1_LOC_763/A
+ NOR2X1_LOC_48/B NOR2X1_LOC
XNOR2X1_LOC_752 NOR2X1_LOC_752/a_36_216# INVX1_LOC_290/A VSS VDD NOR2X1_LOC_51/A D_INPUT_5
+ NOR2X1_LOC
XNOR2X1_LOC_741 NOR2X1_LOC_741/a_36_216# NOR2X1_LOC_742/A VSS VDD NOR2X1_LOC_741/A
+ NOR2X1_LOC_736/Y NOR2X1_LOC
XNOR2X1_LOC_796 NOR2X1_LOC_796/a_36_216# NOR2X1_LOC_803/B VSS VDD NOR2X1_LOC_784/Y
+ NOR2X1_LOC_796/B NOR2X1_LOC
XNOR2X1_LOC_730 NOR2X1_LOC_730/a_36_216# NOR2X1_LOC_730/Y VSS VDD NOR2X1_LOC_730/A
+ NOR2X1_LOC_730/B NOR2X1_LOC
XNOR2X1_LOC_774 NOR2X1_LOC_774/a_36_216# INVX1_LOC_300/A VSS VDD NOR2X1_LOC_773/Y
+ INVX1_LOC_297/Y NOR2X1_LOC
XNOR2X1_LOC_785 NOR2X1_LOC_785/a_36_216# NOR2X1_LOC_785/Y VSS VDD NOR2X1_LOC_785/A
+ NOR2X1_LOC_775/Y NOR2X1_LOC
XNAND2X1_LOC_527 NAND2X1_LOC_527/a_36_24# NOR2X1_LOC_547/B VSS VDD INVX1_LOC_49/A
+ NAND2X1_LOC_323/B NAND2X1_LOC
XNAND2X1_LOC_549 NAND2X1_LOC_549/a_36_24# NAND2X1_LOC_549/Y VSS VDD INVX1_LOC_219/Y
+ NAND2X1_LOC_549/B NAND2X1_LOC
XNAND2X1_LOC_505 NAND2X1_LOC_505/a_36_24# NOR2X1_LOC_507/A VSS VDD INVX1_LOC_15/A
+ NOR2X1_LOC_160/B NAND2X1_LOC
XNAND2X1_LOC_538 NAND2X1_LOC_538/a_36_24# NAND2X1_LOC_538/Y VSS VDD NOR2X1_LOC_13/Y
+ NOR2X1_LOC_311/Y NAND2X1_LOC
XNAND2X1_LOC_516 NAND2X1_LOC_516/a_36_24# NOR2X1_LOC_574/A VSS VDD NOR2X1_LOC_513/Y
+ INVX1_LOC_215/Y NAND2X1_LOC
XINVX1_LOC_180 INVX1_LOC_180/Y VSS VDD INVX1_LOC_180/A INVX1_LOC
XINVX1_LOC_191 INVX1_LOC_191/Y VSS VDD INVX1_LOC_191/A INVX1_LOC
XNOR2X1_LOC_571 NOR2X1_LOC_571/a_36_216# NOR2X1_LOC_576/B VSS VDD NOR2X1_LOC_561/Y
+ INVX1_LOC_229/Y NOR2X1_LOC
XNOR2X1_LOC_560 NOR2X1_LOC_560/a_36_216# INVX1_LOC_230/A VSS VDD NOR2X1_LOC_560/A
+ NOR2X1_LOC_844/A NOR2X1_LOC
XNOR2X1_LOC_582 NOR2X1_LOC_582/a_36_216# NOR2X1_LOC_582/Y VSS VDD NOR2X1_LOC_582/A
+ INVX1_LOC_78/A NOR2X1_LOC
XNOR2X1_LOC_593 NOR2X1_LOC_593/a_36_216# NOR2X1_LOC_593/Y VSS VDD INVX1_LOC_245/Y
+ NOR2X1_LOC_718/B NOR2X1_LOC
XNAND2X1_LOC_302 NAND2X1_LOC_302/a_36_24# NAND2X1_LOC_303/B VSS VDD NOR2X1_LOC_298/Y
+ NOR2X1_LOC_299/Y NAND2X1_LOC
XNAND2X1_LOC_346 NAND2X1_LOC_346/a_36_24# NAND2X1_LOC_347/B VSS VDD NOR2X1_LOC_292/Y
+ NOR2X1_LOC_295/Y NAND2X1_LOC
XNAND2X1_LOC_357 NAND2X1_LOC_357/a_36_24# NAND2X1_LOC_364/A VSS VDD NAND2X1_LOC_357/A
+ NAND2X1_LOC_357/B NAND2X1_LOC
XNAND2X1_LOC_335 NAND2X1_LOC_335/a_36_24# INVX1_LOC_149/A VSS VDD NOR2X1_LOC_309/Y
+ NOR2X1_LOC_310/Y NAND2X1_LOC
XNAND2X1_LOC_379 NAND2X1_LOC_379/a_36_24# NOR2X1_LOC_380/A VSS VDD INVX1_LOC_11/Y
+ INVX1_LOC_20/A NAND2X1_LOC
XNAND2X1_LOC_324 NAND2X1_LOC_324/a_36_24# NAND2X1_LOC_326/A VSS VDD NOR2X1_LOC_320/Y
+ NOR2X1_LOC_321/Y NAND2X1_LOC
XNAND2X1_LOC_313 NAND2X1_LOC_313/a_36_24# NOR2X1_LOC_317/B VSS VDD INVX1_LOC_53/A
+ NOR2X1_LOC_383/B NAND2X1_LOC
XNAND2X1_LOC_368 NAND2X1_LOC_368/a_36_24# NOR2X1_LOC_457/B VSS VDD INVX1_LOC_6/Y NOR2X1_LOC_270/Y
+ NAND2X1_LOC
XNOR2X1_LOC_390 NOR2X1_LOC_390/a_36_216# NOR2X1_LOC_392/B VSS VDD INVX1_LOC_161/Y
+ NOR2X1_LOC_388/Y NOR2X1_LOC
XNAND2X1_LOC_110 NAND2X1_LOC_110/a_36_24# NAND2X1_LOC_323/B VSS VDD D_INPUT_0
+ INVX1_LOC_13/A NAND2X1_LOC
XNAND2X1_LOC_143 NAND2X1_LOC_143/a_36_24# INVX1_LOC_83/A VSS VDD D_INPUT_1 INVX1_LOC_7/A
+ NAND2X1_LOC
XNAND2X1_LOC_132 NAND2X1_LOC_132/a_36_24# NOR2X1_LOC_137/B VSS VDD NOR2X1_LOC_383/B
+ INVX1_LOC_57/A NAND2X1_LOC
XNAND2X1_LOC_121 NAND2X1_LOC_121/a_36_24# NOR2X1_LOC_122/A VSS VDD INVX1_LOC_72/A
+ NOR2X1_LOC_666/A NAND2X1_LOC
XNAND2X1_LOC_198 NAND2X1_LOC_198/a_36_24# NAND2X1_LOC_208/B VSS VDD INVX1_LOC_43/Y
+ NAND2X1_LOC_198/B NAND2X1_LOC
XNAND2X1_LOC_187 NAND2X1_LOC_187/a_36_24# NOR2X1_LOC_191/B VSS VDD INVX1_LOC_29/A
+ NOR2X1_LOC_186/Y NAND2X1_LOC
XNAND2X1_LOC_165 NAND2X1_LOC_165/a_36_24# NOR2X1_LOC_168/A VSS VDD INVX1_LOC_37/A
+ NAND2X1_LOC_74/B NAND2X1_LOC
XNAND2X1_LOC_176 NAND2X1_LOC_176/a_36_24# NOR2X1_LOC_180/B VSS VDD INVX1_LOC_19/A
+ NOR2X1_LOC_383/B NAND2X1_LOC
XNAND2X1_LOC_154 NAND2X1_LOC_154/a_36_24# NAND2X1_LOC_154/Y VSS VDD INVX1_LOC_6/A
+ INVX1_LOC_28/A NAND2X1_LOC
XNOR2X1_LOC_219 NOR2X1_LOC_219/a_36_216# NOR2X1_LOC_219/Y VSS VDD NOR2X1_LOC_215/Y
+ NOR2X1_LOC_219/B NOR2X1_LOC
XNOR2X1_LOC_208 NOR2X1_LOC_208/a_36_216# NOR2X1_LOC_208/Y VSS VDD NOR2X1_LOC_208/A
+ NOR2X1_LOC_35/Y NOR2X1_LOC
XNAND2X1_LOC_709 NAND2X1_LOC_709/a_36_24# INVX1_LOC_277/A VSS VDD NOR2X1_LOC_698/Y
+ NOR2X1_LOC_748/A NAND2X1_LOC
XNOR2X1_LOC_742 NOR2X1_LOC_742/a_36_216# D_GATE_741 VSS VDD NOR2X1_LOC_742/A NOR2X1_LOC_740/Y
+ NOR2X1_LOC
XNOR2X1_LOC_731 NOR2X1_LOC_731/a_36_216# NOR2X1_LOC_731/Y VSS VDD NOR2X1_LOC_731/A
+ NOR2X1_LOC_726/Y NOR2X1_LOC
XNOR2X1_LOC_753 NOR2X1_LOC_753/a_36_216# NOR2X1_LOC_753/Y VSS VDD INVX1_LOC_289/Y
+ NOR2X1_LOC_816/A NOR2X1_LOC
XNOR2X1_LOC_720 NOR2X1_LOC_720/a_36_216# NOR2X1_LOC_721/A VSS VDD NOR2X1_LOC_720/A
+ NOR2X1_LOC_720/B NOR2X1_LOC
XNOR2X1_LOC_764 NOR2X1_LOC_764/a_36_216# NOR2X1_LOC_764/Y VSS VDD INVX1_LOC_76/A INVX1_LOC_30/A
+ NOR2X1_LOC
XNOR2X1_LOC_797 NOR2X1_LOC_797/a_36_216# NOR2X1_LOC_803/A VSS VDD INVX1_LOC_301/Y
+ NOR2X1_LOC_209/B NOR2X1_LOC
XNOR2X1_LOC_775 NOR2X1_LOC_775/a_36_216# NOR2X1_LOC_775/Y VSS VDD NOR2X1_LOC_112/B
+ NOR2X1_LOC_97/A NOR2X1_LOC
XNOR2X1_LOC_786 NOR2X1_LOC_786/a_36_216# INVX1_LOC_304/A VSS VDD NOR2X1_LOC_266/B
+ NOR2X1_LOC_84/Y NOR2X1_LOC
XINVX1_LOC_170 INVX1_LOC_170/Y VSS VDD INVX1_LOC_170/A INVX1_LOC
XNAND2X1_LOC_517 NAND2X1_LOC_517/a_36_24# NOR2X1_LOC_559/B VSS VDD INVX1_LOC_22/Y
+ NOR2X1_LOC_264/Y NAND2X1_LOC
XNAND2X1_LOC_528 NAND2X1_LOC_528/a_36_24# NOR2X1_LOC_620/B VSS VDD INVX1_LOC_5/A INVX1_LOC_33/A
+ NAND2X1_LOC
XNAND2X1_LOC_506 NAND2X1_LOC_506/a_36_24# NAND2X1_LOC_508/A VSS VDD INVX1_LOC_120/A
+ NOR2X1_LOC_419/Y NAND2X1_LOC
XNAND2X1_LOC_539 NAND2X1_LOC_539/a_36_24# NAND2X1_LOC_799/A VSS VDD NAND2X1_LOC_537/Y
+ NAND2X1_LOC_538/Y NAND2X1_LOC
XINVX1_LOC_181 INVX1_LOC_181/Y VSS VDD INVX1_LOC_181/A INVX1_LOC
XINVX1_LOC_192 INVX1_LOC_192/Y VSS VDD INVX1_LOC_192/A INVX1_LOC
XNOR2X1_LOC_583 NOR2X1_LOC_583/a_36_216# NOR2X1_LOC_583/Y VSS VDD NOR2X1_LOC_52/B
+ INVX1_LOC_22/A NOR2X1_LOC
XNOR2X1_LOC_594 NOR2X1_LOC_594/a_36_216# NOR2X1_LOC_594/Y VSS VDD NOR2X1_LOC_331/B
+ INVX1_LOC_58/A NOR2X1_LOC
XNOR2X1_LOC_550 NOR2X1_LOC_550/a_36_216# NOR2X1_LOC_565/A VSS VDD INVX1_LOC_225/Y
+ NOR2X1_LOC_550/B NOR2X1_LOC
XNOR2X1_LOC_561 NOR2X1_LOC_561/a_36_216# NOR2X1_LOC_561/Y VSS VDD NOR2X1_LOC_561/A
+ NOR2X1_LOC_557/Y NOR2X1_LOC
XNOR2X1_LOC_572 NOR2X1_LOC_572/a_36_216# INVX1_LOC_234/A VSS VDD NOR2X1_LOC_361/B
+ INVX1_LOC_74/A NOR2X1_LOC
XNAND2X1_LOC_325 NAND2X1_LOC_325/a_36_24# NAND2X1_LOC_325/Y VSS VDD NOR2X1_LOC_322/Y
+ NOR2X1_LOC_323/Y NAND2X1_LOC
XNAND2X1_LOC_336 NAND2X1_LOC_336/a_36_24# NAND2X1_LOC_337/B VSS VDD NOR2X1_LOC_311/Y
+ NOR2X1_LOC_312/Y NAND2X1_LOC
XNAND2X1_LOC_314 NAND2X1_LOC_314/a_36_24# NOR2X1_LOC_317/A VSS VDD NOR2X1_LOC_78/B
+ INVX1_LOC_49/A NAND2X1_LOC
XNAND2X1_LOC_303 NAND2X1_LOC_303/a_36_24# NAND2X1_LOC_303/Y VSS VDD INVX1_LOC_140/Y
+ NAND2X1_LOC_303/B NAND2X1_LOC
XNAND2X1_LOC_347 NAND2X1_LOC_347/a_36_24# NAND2X1_LOC_360/B VSS VDD INVX1_LOC_137/Y
+ NAND2X1_LOC_347/B NAND2X1_LOC
XNAND2X1_LOC_358 NAND2X1_LOC_358/a_36_24# NAND2X1_LOC_358/Y VSS VDD INVX1_LOC_158/Y
+ NAND2X1_LOC_358/B NAND2X1_LOC
XNAND2X1_LOC_369 NAND2X1_LOC_369/a_36_24# NOR2X1_LOC_543/A VSS VDD INVX1_LOC_17/A
+ INVX1_LOC_71/A NAND2X1_LOC
XNOR2X1_LOC_391 NOR2X1_LOC_391/a_36_216# NOR2X1_LOC_391/Y VSS VDD NOR2X1_LOC_391/A
+ NOR2X1_LOC_391/B NOR2X1_LOC
XNOR2X1_LOC_380 NOR2X1_LOC_380/a_36_216# NOR2X1_LOC_380/Y VSS VDD NOR2X1_LOC_380/A
+ INVX1_LOC_76/A NOR2X1_LOC
XNAND2X1_LOC_100 NAND2X1_LOC_100/a_36_24# INVX1_LOC_61/A VSS VDD NOR2X1_LOC_86/Y NOR2X1_LOC_88/Y
+ NAND2X1_LOC
XNAND2X1_LOC_122 NAND2X1_LOC_122/a_36_24# NOR2X1_LOC_124/B VSS VDD INVX1_LOC_33/A
+ NOR2X1_LOC_121/Y NAND2X1_LOC
XNAND2X1_LOC_133 NAND2X1_LOC_133/a_36_24# INVX1_LOC_77/A VSS VDD INVX1_LOC_7/A NOR2X1_LOC_82/A
+ NAND2X1_LOC
XNAND2X1_LOC_111 NAND2X1_LOC_111/a_36_24# NOR2X1_LOC_332/B VSS VDD INVX1_LOC_21/A
+ NAND2X1_LOC_323/B NAND2X1_LOC
XNAND2X1_LOC_166 NAND2X1_LOC_166/a_36_24# NOR2X1_LOC_169/B VSS VDD NOR2X1_LOC_78/B
+ INVX1_LOC_29/A NAND2X1_LOC
XNAND2X1_LOC_177 NAND2X1_LOC_177/a_36_24# NOR2X1_LOC_439/B VSS VDD NOR2X1_LOC_68/A
+ INVX1_LOC_53/A NAND2X1_LOC
XNAND2X1_LOC_155 NAND2X1_LOC_155/a_36_24# NAND2X1_LOC_156/B VSS VDD NOR2X1_LOC_52/B
+ NOR2X1_LOC_433/A NAND2X1_LOC
XNAND2X1_LOC_144 NAND2X1_LOC_144/a_36_24# NOR2X1_LOC_147/A VSS VDD INVX1_LOC_45/A
+ INVX1_LOC_83/A NAND2X1_LOC
XNAND2X1_LOC_188 NAND2X1_LOC_188/a_36_24# NOR2X1_LOC_189/A VSS VDD INVX1_LOC_28/A
+ NOR2X1_LOC_816/A NAND2X1_LOC
XNAND2X1_LOC_199 NAND2X1_LOC_199/a_36_24# INVX1_LOC_107/A VSS VDD NAND2X1_LOC_195/Y
+ NAND2X1_LOC_199/B NAND2X1_LOC
XINVX1_LOC_90 INVX1_LOC_90/Y VSS VDD INVX1_LOC_90/A INVX1_LOC
XNOR2X1_LOC_1 NOR2X1_LOC_1/a_36_216# NOR2X1_LOC_1/Y VSS VDD D_INPUT_7 INPUT_6
+ NOR2X1_LOC
XNOR2X1_LOC_209 NOR2X1_LOC_209/a_36_216# NOR2X1_LOC_209/Y VSS VDD NOR2X1_LOC_209/A
+ NOR2X1_LOC_209/B NOR2X1_LOC
XNOR2X1_LOC_732 NOR2X1_LOC_732/a_36_216# NOR2X1_LOC_738/A VSS VDD NOR2X1_LOC_732/A
+ NOR2X1_LOC_724/Y NOR2X1_LOC
XNOR2X1_LOC_710 NOR2X1_LOC_710/a_36_216# NOR2X1_LOC_711/A VSS VDD NOR2X1_LOC_710/A
+ NOR2X1_LOC_710/B NOR2X1_LOC
XNOR2X1_LOC_787 NOR2X1_LOC_787/a_36_216# NOR2X1_LOC_794/B VSS VDD NOR2X1_LOC_486/Y
+ NOR2X1_LOC_457/A NOR2X1_LOC
XNOR2X1_LOC_765 NOR2X1_LOC_765/a_36_216# NOR2X1_LOC_765/Y VSS VDD NOR2X1_LOC_15/Y
+ INVX1_LOC_11/Y NOR2X1_LOC
XNOR2X1_LOC_743 NOR2X1_LOC_743/a_36_216# NOR2X1_LOC_743/Y VSS VDD NOR2X1_LOC_433/A
+ INVX1_LOC_1/Y NOR2X1_LOC
XNOR2X1_LOC_721 NOR2X1_LOC_721/a_36_216# NOR2X1_LOC_721/Y VSS VDD NOR2X1_LOC_721/A
+ NOR2X1_LOC_721/B NOR2X1_LOC
XNOR2X1_LOC_754 NOR2X1_LOC_754/a_36_216# NOR2X1_LOC_754/Y VSS VDD NOR2X1_LOC_754/A
+ INVX1_LOC_24/A NOR2X1_LOC
XNOR2X1_LOC_776 NOR2X1_LOC_776/a_36_216# NOR2X1_LOC_785/A VSS VDD NOR2X1_LOC_241/A
+ NOR2X1_LOC_168/B NOR2X1_LOC
XNOR2X1_LOC_798 NOR2X1_LOC_798/a_36_216# NOR2X1_LOC_798/Y VSS VDD NOR2X1_LOC_798/A
+ NOR2X1_LOC_354/B NOR2X1_LOC
XNAND2X1_LOC_518 NAND2X1_LOC_518/a_36_24# NOR2X1_LOC_520/B VSS VDD INVX1_LOC_49/A
+ NAND2X1_LOC_74/B NAND2X1_LOC
XNAND2X1_LOC_507 NAND2X1_LOC_507/a_36_24# INVX1_LOC_209/A VSS VDD NOR2X1_LOC_504/Y
+ NOR2X1_LOC_505/Y NAND2X1_LOC
XINVX1_LOC_160 INVX1_LOC_160/Y VSS VDD INVX1_LOC_160/A INVX1_LOC
XINVX1_LOC_171 INVX1_LOC_171/Y VSS VDD INVX1_LOC_171/A INVX1_LOC
XINVX1_LOC_182 INVX1_LOC_182/Y VSS VDD INVX1_LOC_182/A INVX1_LOC
XINVX1_LOC_193 INVX1_LOC_193/Y VSS VDD INVX1_LOC_193/A INVX1_LOC
XNAND2X1_LOC_529 NAND2X1_LOC_529/a_36_24# NOR2X1_LOC_548/B VSS VDD INPUT_3 INVX1_LOC_19/A
+ NAND2X1_LOC
XNOR2X1_LOC_584 NOR2X1_LOC_584/a_36_216# NOR2X1_LOC_584/Y VSS VDD INVX1_LOC_38/A INVX1_LOC_6/A
+ NOR2X1_LOC
XNOR2X1_LOC_562 NOR2X1_LOC_562/a_36_216# NOR2X1_LOC_570/B VSS VDD NOR2X1_LOC_562/A
+ NOR2X1_LOC_562/B NOR2X1_LOC
XNOR2X1_LOC_540 NOR2X1_LOC_540/a_36_216# NOR2X1_LOC_553/B VSS VDD INVX1_LOC_97/A NOR2X1_LOC_540/B
+ NOR2X1_LOC
XNOR2X1_LOC_551 NOR2X1_LOC_551/a_36_216# NOR2X1_LOC_551/Y VSS VDD INVX1_LOC_223/Y
+ NOR2X1_LOC_551/B NOR2X1_LOC
XNOR2X1_LOC_595 NOR2X1_LOC_595/a_36_216# NOR2X1_LOC_595/Y VSS VDD NOR2X1_LOC_250/A
+ INVX1_LOC_20/A NOR2X1_LOC
XNOR2X1_LOC_573 NOR2X1_LOC_573/a_36_216# NOR2X1_LOC_573/Y VSS VDD INVX1_LOC_207/Y
+ NOR2X1_LOC_474/A NOR2X1_LOC
XNAND2X1_LOC_359 NAND2X1_LOC_359/a_36_24# NAND2X1_LOC_359/Y VSS VDD NAND2X1_LOC_359/A
+ INVX1_LOC_156/Y NAND2X1_LOC
XNAND2X1_LOC_348 NAND2X1_LOC_348/a_36_24# NAND2X1_LOC_359/A VSS VDD NAND2X1_LOC_348/A
+ INVX1_LOC_154/Y NAND2X1_LOC
XNAND2X1_LOC_337 NAND2X1_LOC_337/a_36_24# NAND2X1_LOC_352/B VSS VDD INVX1_LOC_150/Y
+ NAND2X1_LOC_337/B NAND2X1_LOC
XNAND2X1_LOC_315 NAND2X1_LOC_315/a_36_24# NOR2X1_LOC_318/B VSS VDD INVX1_LOC_21/A
+ INVX1_LOC_77/A NAND2X1_LOC
XNAND2X1_LOC_326 NAND2X1_LOC_326/a_36_24# NAND2X1_LOC_354/B VSS VDD NAND2X1_LOC_326/A
+ NAND2X1_LOC_325/Y NAND2X1_LOC
XNAND2X1_LOC_304 NAND2X1_LOC_304/a_36_24# NOR2X1_LOC_307/B VSS VDD NAND2X1_LOC_53/Y
+ INVX1_LOC_117/A NAND2X1_LOC
XNOR2X1_LOC_370 NOR2X1_LOC_370/a_36_216# NOR2X1_LOC_457/A VSS VDD NOR2X1_LOC_543/A
+ NOR2X1_LOC_335/B NOR2X1_LOC
XNOR2X1_LOC_381 NOR2X1_LOC_381/a_36_216# NOR2X1_LOC_381/Y VSS VDD INVX1_LOC_12/A D_INPUT_3
+ NOR2X1_LOC
XNOR2X1_LOC_392 NOR2X1_LOC_392/a_36_216# NOR2X1_LOC_392/Y VSS VDD NOR2X1_LOC_391/Y
+ NOR2X1_LOC_392/B NOR2X1_LOC
XNAND2X1_LOC_860 NAND2X1_LOC_860/a_36_24# NAND2X1_LOC_860/Y VSS VDD NAND2X1_LOC_860/A
+ NAND2X1_LOC_392/Y NAND2X1_LOC
XNAND2X1_LOC_101 NAND2X1_LOC_101/a_36_24# NAND2X1_LOC_656/A VSS VDD NAND2X1_LOC_99/Y
+ INVX1_LOC_62/Y NAND2X1_LOC
XNAND2X1_LOC_134 NAND2X1_LOC_134/a_36_24# NOR2X1_LOC_137/A VSS VDD INVX1_LOC_57/A
+ INVX1_LOC_77/A NAND2X1_LOC
XNAND2X1_LOC_189 NAND2X1_LOC_189/a_36_24# INVX1_LOC_101/A VSS VDD INVX1_LOC_57/A NOR2X1_LOC_188/Y
+ NAND2X1_LOC
XNAND2X1_LOC_123 NAND2X1_LOC_123/a_36_24# NAND2X1_LOC_123/Y VSS VDD NOR2X1_LOC_117/Y
+ INVX1_LOC_69/Y NAND2X1_LOC
XNAND2X1_LOC_167 NAND2X1_LOC_167/a_36_24# NOR2X1_LOC_703/B VSS VDD INVX1_LOC_49/A
+ INVX1_LOC_91/A NAND2X1_LOC
XNAND2X1_LOC_112 NAND2X1_LOC_112/a_36_24# NAND2X1_LOC_112/Y VSS VDD NOR2X1_LOC_109/Y
+ NOR2X1_LOC_111/Y NAND2X1_LOC
XNAND2X1_LOC_145 NAND2X1_LOC_145/a_36_24# NOR2X1_LOC_148/B VSS VDD INVX1_LOC_37/A
+ NOR2X1_LOC_78/A NAND2X1_LOC
XNAND2X1_LOC_178 NAND2X1_LOC_178/a_36_24# NOR2X1_LOC_540/B VSS VDD INVX1_LOC_41/A
+ INVX1_LOC_89/A NAND2X1_LOC
XNAND2X1_LOC_156 NAND2X1_LOC_156/a_36_24# NOR2X1_LOC_158/B VSS VDD NAND2X1_LOC_154/Y
+ NAND2X1_LOC_156/B NAND2X1_LOC
XNAND2X1_LOC_690 NAND2X1_LOC_690/a_36_24# NOR2X1_LOC_691/A VSS VDD D_INPUT_0 NOR2X1_LOC_634/A
+ NAND2X1_LOC
XINVX1_LOC_80 INVX1_LOC_80/Y VSS VDD INVX1_LOC_80/A INVX1_LOC
XINVX1_LOC_91 INVX1_LOC_91/Y VSS VDD INVX1_LOC_91/A INVX1_LOC
XNOR2X1_LOC_2 NOR2X1_LOC_2/a_36_216# NOR2X1_LOC_2/Y VSS VDD INPUT_5 INPUT_4 NOR2X1_LOC
XNOR2X1_LOC_733 NOR2X1_LOC_733/a_36_216# NOR2X1_LOC_733/Y VSS VDD NOR2X1_LOC_723/Y
+ NOR2X1_LOC_722/Y NOR2X1_LOC
XNOR2X1_LOC_722 NOR2X1_LOC_722/a_36_216# NOR2X1_LOC_722/Y VSS VDD INVX1_LOC_283/Y
+ NOR2X1_LOC_718/Y NOR2X1_LOC
XNOR2X1_LOC_711 NOR2X1_LOC_711/a_36_216# NOR2X1_LOC_711/Y VSS VDD NOR2X1_LOC_711/A
+ INVX1_LOC_277/Y NOR2X1_LOC
XNOR2X1_LOC_777 NOR2X1_LOC_777/a_36_216# NOR2X1_LOC_784/B VSS VDD NOR2X1_LOC_307/A
+ NOR2X1_LOC_777/B NOR2X1_LOC
XNOR2X1_LOC_755 NOR2X1_LOC_755/a_36_216# NOR2X1_LOC_755/Y VSS VDD NOR2X1_LOC_665/A
+ INVX1_LOC_45/Y NOR2X1_LOC
XNOR2X1_LOC_788 NOR2X1_LOC_788/a_36_216# NOR2X1_LOC_794/A VSS VDD INVX1_LOC_247/Y
+ NOR2X1_LOC_788/B NOR2X1_LOC
XNOR2X1_LOC_766 NOR2X1_LOC_766/a_36_216# NOR2X1_LOC_766/Y VSS VDD NOR2X1_LOC_91/A
+ INVX1_LOC_50/A NOR2X1_LOC
XNOR2X1_LOC_744 NOR2X1_LOC_744/a_36_216# NOR2X1_LOC_744/Y VSS VDD INVX1_LOC_76/A INVX1_LOC_33/Y
+ NOR2X1_LOC
XNOR2X1_LOC_799 NOR2X1_LOC_799/a_36_216# NOR2X1_LOC_802/A VSS VDD NOR2X1_LOC_593/Y
+ NOR2X1_LOC_799/B NOR2X1_LOC
XNOR2X1_LOC_700 NOR2X1_LOC_700/a_36_216# NOR2X1_LOC_700/Y VSS VDD NOR2X1_LOC_91/A
+ INVX1_LOC_46/A NOR2X1_LOC
XNAND2X1_LOC_519 NAND2X1_LOC_519/a_36_24# NOR2X1_LOC_520/A VSS VDD NOR2X1_LOC_598/B
+ INVX1_LOC_89/A NAND2X1_LOC
XNAND2X1_LOC_508 NAND2X1_LOC_508/a_36_24# NAND2X1_LOC_510/A VSS VDD NAND2X1_LOC_508/A
+ INVX1_LOC_210/Y NAND2X1_LOC
XINVX1_LOC_194 INVX1_LOC_194/Y VSS VDD INVX1_LOC_194/A INVX1_LOC
XINVX1_LOC_172 INVX1_LOC_172/Y VSS VDD INVX1_LOC_172/A INVX1_LOC
XINVX1_LOC_183 INVX1_LOC_183/Y VSS VDD INVX1_LOC_183/A INVX1_LOC
XINVX1_LOC_150 INVX1_LOC_150/Y VSS VDD INVX1_LOC_150/A INVX1_LOC
XINVX1_LOC_161 INVX1_LOC_161/Y VSS VDD INVX1_LOC_161/A INVX1_LOC
XNOR2X1_LOC_585 NOR2X1_LOC_585/a_36_216# NOR2X1_LOC_585/Y VSS VDD INVX1_LOC_136/A
+ INVX1_LOC_18/A NOR2X1_LOC
XNOR2X1_LOC_596 NOR2X1_LOC_596/a_36_216# NOR2X1_LOC_596/Y VSS VDD NOR2X1_LOC_596/A
+ INVX1_LOC_33/A NOR2X1_LOC
XNOR2X1_LOC_574 NOR2X1_LOC_574/a_36_216# INVX1_LOC_236/A VSS VDD NOR2X1_LOC_574/A
+ NOR2X1_LOC_510/Y NOR2X1_LOC
XNOR2X1_LOC_563 NOR2X1_LOC_563/a_36_216# NOR2X1_LOC_570/A VSS VDD INVX1_LOC_227/Y
+ NOR2X1_LOC_553/Y NOR2X1_LOC
XNOR2X1_LOC_552 NOR2X1_LOC_552/a_36_216# NOR2X1_LOC_552/Y VSS VDD NOR2X1_LOC_552/A
+ NOR2X1_LOC_542/Y NOR2X1_LOC
XNOR2X1_LOC_541 NOR2X1_LOC_541/a_36_216# NOR2X1_LOC_541/Y VSS VDD NOR2X1_LOC_274/B
+ NOR2X1_LOC_541/B NOR2X1_LOC
XNOR2X1_LOC_530 NOR2X1_LOC_530/a_36_216# NOR2X1_LOC_530/Y VSS VDD NOR2X1_LOC_536/A
+ INVX1_LOC_23/Y NOR2X1_LOC
XNAND2X1_LOC_338 NAND2X1_LOC_338/a_36_24# NAND2X1_LOC_351/A VSS VDD INVX1_LOC_148/Y
+ NAND2X1_LOC_338/B NAND2X1_LOC
XNAND2X1_LOC_316 NAND2X1_LOC_316/a_36_24# NOR2X1_LOC_318/A VSS VDD INVX1_LOC_11/A
+ NAND2X1_LOC_81/B NAND2X1_LOC
XNAND2X1_LOC_349 NAND2X1_LOC_349/a_36_24# INVX1_LOC_155/A VSS VDD NAND2X1_LOC_342/Y
+ NAND2X1_LOC_349/B NAND2X1_LOC
XNAND2X1_LOC_327 NAND2X1_LOC_327/a_36_24# NOR2X1_LOC_329/B VSS VDD NOR2X1_LOC_65/B
+ NOR2X1_LOC_667/A NAND2X1_LOC
XNAND2X1_LOC_305 NAND2X1_LOC_305/a_36_24# NOR2X1_LOC_307/A VSS VDD INVX1_LOC_1/A NOR2X1_LOC_383/B
+ NAND2X1_LOC
XNOR2X1_LOC_360 NOR2X1_LOC_360/a_36_216# NOR2X1_LOC_360/Y VSS VDD NOR2X1_LOC_360/A
+ NOR2X1_LOC_860/B NOR2X1_LOC
XNOR2X1_LOC_382 NOR2X1_LOC_382/a_36_216# NOR2X1_LOC_382/Y VSS VDD NOR2X1_LOC_381/Y
+ NOR2X1_LOC_38/B NOR2X1_LOC
XNOR2X1_LOC_393 NOR2X1_LOC_393/a_36_216# NOR2X1_LOC_393/Y VSS VDD INVX1_LOC_30/A INVX1_LOC_28/A
+ NOR2X1_LOC
XNOR2X1_LOC_371 NOR2X1_LOC_371/a_36_216# NOR2X1_LOC_372/A VSS VDD INVX1_LOC_22/A INVX1_LOC_3/Y
+ NOR2X1_LOC
XNAND2X1_LOC_850 NAND2X1_LOC_850/a_36_24# NAND2X1_LOC_850/Y VSS VDD NAND2X1_LOC_850/A
+ INVX1_LOC_314/Y NAND2X1_LOC
XNAND2X1_LOC_861 NAND2X1_LOC_861/a_36_24# NAND2X1_LOC_861/Y VSS VDD INVX1_LOC_256/Y
+ NAND2X1_LOC_860/Y NAND2X1_LOC
XNAND2X1_LOC_102 NAND2X1_LOC_102/a_36_24# NOR2X1_LOC_590/A VSS VDD INVX1_LOC_7/A INVX1_LOC_39/A
+ NAND2X1_LOC
XNAND2X1_LOC_113 NAND2X1_LOC_113/a_36_24# NAND2X1_LOC_114/B VSS VDD NOR2X1_LOC_103/Y
+ NOR2X1_LOC_107/Y NAND2X1_LOC
XNAND2X1_LOC_135 NAND2X1_LOC_135/a_36_24# NOR2X1_LOC_332/A VSS VDD INVX1_LOC_45/A
+ INVX1_LOC_77/A NAND2X1_LOC
XNAND2X1_LOC_168 NAND2X1_LOC_168/a_36_24# NAND2X1_LOC_170/A VSS VDD NOR2X1_LOC_164/Y
+ NOR2X1_LOC_165/Y NAND2X1_LOC
XNAND2X1_LOC_124 NAND2X1_LOC_124/a_36_24# INVX1_LOC_73/A VSS VDD NOR2X1_LOC_122/Y
+ NAND2X1_LOC_123/Y NAND2X1_LOC
XNAND2X1_LOC_179 NAND2X1_LOC_179/a_36_24# NOR2X1_LOC_181/A VSS VDD INVX1_LOC_23/A
+ INVX1_LOC_63/A NAND2X1_LOC
XNAND2X1_LOC_146 NAND2X1_LOC_146/a_36_24# NOR2X1_LOC_148/A VSS VDD INVX1_LOC_23/A
+ INVX1_LOC_75/A NAND2X1_LOC
XNAND2X1_LOC_157 NAND2X1_LOC_157/a_36_24# INVX1_LOC_89/A VSS VDD NAND2X1_LOC_3/B NAND2X1_LOC_36/A
+ NAND2X1_LOC
XNOR2X1_LOC_190 NOR2X1_LOC_190/a_36_216# NOR2X1_LOC_191/A VSS VDD INVX1_LOC_100/Y
+ INVX1_LOC_98/Y NOR2X1_LOC
XNAND2X1_LOC_691 NAND2X1_LOC_691/a_36_24# NAND2X1_LOC_729/B VSS VDD NOR2X1_LOC_689/Y
+ NOR2X1_LOC_690/Y NAND2X1_LOC
XNAND2X1_LOC_680 NAND2X1_LOC_680/a_36_24# INVX1_LOC_273/A VSS VDD INVX1_LOC_37/A NOR2X1_LOC_186/Y
+ NAND2X1_LOC
XINVX1_LOC_92 INVX1_LOC_92/Y VSS VDD INVX1_LOC_92/A INVX1_LOC
XINVX1_LOC_70 INVX1_LOC_70/Y VSS VDD INVX1_LOC_70/A INVX1_LOC
XINVX1_LOC_81 INVX1_LOC_81/Y VSS VDD INVX1_LOC_81/A INVX1_LOC
XNOR2X1_LOC_3 NOR2X1_LOC_3/a_36_216# INVX1_LOC_2/A VSS VDD NOR2X1_LOC_2/Y NOR2X1_LOC_1/Y
+ NOR2X1_LOC
XINVX1_LOC_310 INVX1_LOC_310/Y VSS VDD INVX1_LOC_310/A INVX1_LOC
XNOR2X1_LOC_701 NOR2X1_LOC_701/a_36_216# NOR2X1_LOC_701/Y VSS VDD INVX1_LOC_118/A
+ INVX1_LOC_34/A NOR2X1_LOC
XNOR2X1_LOC_712 NOR2X1_LOC_712/a_36_216# NOR2X1_LOC_712/Y VSS VDD NOR2X1_LOC_708/Y
+ NOR2X1_LOC_712/B NOR2X1_LOC
XNOR2X1_LOC_745 NOR2X1_LOC_745/a_36_216# NOR2X1_LOC_745/Y VSS VDD INVX1_LOC_92/A INVX1_LOC_30/A
+ NOR2X1_LOC
XNOR2X1_LOC_723 NOR2X1_LOC_723/a_36_216# NOR2X1_LOC_723/Y VSS VDD NOR2X1_LOC_717/Y
+ INVX1_LOC_281/Y NOR2X1_LOC
XNOR2X1_LOC_778 NOR2X1_LOC_778/a_36_216# NOR2X1_LOC_778/Y VSS VDD NOR2X1_LOC_778/A
+ NOR2X1_LOC_778/B NOR2X1_LOC
XNOR2X1_LOC_767 NOR2X1_LOC_767/a_36_216# INVX1_LOC_294/A VSS VDD NOR2X1_LOC_79/A INVX1_LOC_1/Y
+ NOR2X1_LOC
XNOR2X1_LOC_789 NOR2X1_LOC_789/a_36_216# INVX1_LOC_306/A VSS VDD NOR2X1_LOC_789/A
+ NOR2X1_LOC_789/B NOR2X1_LOC
XNOR2X1_LOC_756 NOR2X1_LOC_756/a_36_216# NOR2X1_LOC_756/Y VSS VDD INVX1_LOC_91/A INVX1_LOC_63/A
+ NOR2X1_LOC
XNOR2X1_LOC_734 NOR2X1_LOC_734/a_36_216# INVX1_LOC_286/A VSS VDD NOR2X1_LOC_721/Y
+ INVX1_LOC_171/A NOR2X1_LOC
XNAND2X1_LOC_509 NAND2X1_LOC_509/a_36_24# INVX1_LOC_211/A VSS VDD NAND2X1_LOC_227/Y
+ NOR2X1_LOC_503/Y NAND2X1_LOC
XINVX1_LOC_195 INVX1_LOC_195/Y VSS VDD INVX1_LOC_195/A INVX1_LOC
XINVX1_LOC_184 INVX1_LOC_184/Y VSS VDD INVX1_LOC_184/A INVX1_LOC
XINVX1_LOC_162 INVX1_LOC_162/Y VSS VDD INVX1_LOC_162/A INVX1_LOC
XINVX1_LOC_151 INVX1_LOC_151/Y VSS VDD INVX1_LOC_151/A INVX1_LOC
XINVX1_LOC_173 INVX1_LOC_173/Y VSS VDD INVX1_LOC_173/A INVX1_LOC
XINVX1_LOC_140 INVX1_LOC_140/Y VSS VDD INVX1_LOC_140/A INVX1_LOC
XNOR2X1_LOC_553 NOR2X1_LOC_553/a_36_216# NOR2X1_LOC_553/Y VSS VDD NOR2X1_LOC_541/Y
+ NOR2X1_LOC_553/B NOR2X1_LOC
XNOR2X1_LOC_531 NOR2X1_LOC_531/a_36_216# INVX1_LOC_220/A VSS VDD NOR2X1_LOC_74/A INVX1_LOC_30/A
+ NOR2X1_LOC
XNOR2X1_LOC_542 NOR2X1_LOC_542/a_36_216# NOR2X1_LOC_542/Y VSS VDD NOR2X1_LOC_703/A
+ NOR2X1_LOC_542/B NOR2X1_LOC
XNOR2X1_LOC_520 NOR2X1_LOC_520/a_36_216# INVX1_LOC_218/A VSS VDD NOR2X1_LOC_520/A
+ NOR2X1_LOC_520/B NOR2X1_LOC
XNOR2X1_LOC_586 NOR2X1_LOC_586/a_36_216# NOR2X1_LOC_586/Y VSS VDD NOR2X1_LOC_589/A
+ INVX1_LOC_54/A NOR2X1_LOC
XNOR2X1_LOC_597 NOR2X1_LOC_597/a_36_216# NOR2X1_LOC_597/Y VSS VDD NOR2X1_LOC_597/A
+ INVX1_LOC_10/A NOR2X1_LOC
XNOR2X1_LOC_564 NOR2X1_LOC_564/a_36_216# NOR2X1_LOC_564/Y VSS VDD NOR2X1_LOC_552/Y
+ NOR2X1_LOC_551/Y NOR2X1_LOC
XNOR2X1_LOC_575 NOR2X1_LOC_575/a_36_216# NOR2X1_LOC_575/Y VSS VDD INVX1_LOC_235/Y
+ NOR2X1_LOC_573/Y NOR2X1_LOC
XNAND2X1_LOC_306 NAND2X1_LOC_306/a_36_24# INVX1_LOC_141/A VSS VDD INVX1_LOC_17/A INVX1_LOC_83/A
+ NAND2X1_LOC
XNAND2X1_LOC_339 NAND2X1_LOC_339/a_36_24# INVX1_LOC_151/A VSS VDD NAND2X1_LOC_61/Y
+ NAND2X1_LOC_332/Y NAND2X1_LOC
XNAND2X1_LOC_317 NAND2X1_LOC_317/a_36_24# NAND2X1_LOC_319/A VSS VDD NOR2X1_LOC_313/Y
+ NOR2X1_LOC_314/Y NAND2X1_LOC
XNAND2X1_LOC_328 NAND2X1_LOC_328/a_36_24# NOR2X1_LOC_596/A VSS VDD D_INPUT_4 NAND2X1_LOC_51/B
+ NAND2X1_LOC
XNOR2X1_LOC_361 NOR2X1_LOC_361/a_36_216# NOR2X1_LOC_361/Y VSS VDD NOR2X1_LOC_276/Y
+ NOR2X1_LOC_361/B NOR2X1_LOC
XNOR2X1_LOC_350 NOR2X1_LOC_350/a_36_216# INVX1_LOC_158/A VSS VDD NOR2X1_LOC_350/A
+ NOR2X1_LOC_340/Y NOR2X1_LOC
XNOR2X1_LOC_383 NOR2X1_LOC_383/a_36_216# NOR2X1_LOC_383/Y VSS VDD INVX1_LOC_117/A
+ NOR2X1_LOC_383/B NOR2X1_LOC
XNOR2X1_LOC_394 NOR2X1_LOC_394/a_36_216# NOR2X1_LOC_394/Y VSS VDD INVX1_LOC_76/A INVX1_LOC_36/A
+ NOR2X1_LOC
XNOR2X1_LOC_372 NOR2X1_LOC_372/a_36_216# NOR2X1_LOC_372/Y VSS VDD NOR2X1_LOC_372/A
+ INPUT_1 NOR2X1_LOC
XNAND2X1_LOC_840 NAND2X1_LOC_840/a_36_24# NAND2X1_LOC_840/Y VSS VDD NAND2X1_LOC_833/Y
+ NAND2X1_LOC_840/B NAND2X1_LOC
XNAND2X1_LOC_862 NAND2X1_LOC_862/a_36_24# NAND2X1_LOC_862/Y VSS VDD NAND2X1_LOC_862/A
+ NAND2X1_LOC_859/Y NAND2X1_LOC
XNAND2X1_LOC_851 NAND2X1_LOC_851/a_36_24# NAND2X1_LOC_858/B VSS VDD NAND2X1_LOC_840/Y
+ INVX1_LOC_312/Y NAND2X1_LOC
XNOR2X1_LOC_90 NOR2X1_LOC_90/a_36_216# NOR2X1_LOC_91/A VSS VDD INVX1_LOC_39/Y INVX1_LOC_26/A
+ NOR2X1_LOC
XNAND2X1_LOC_114 NAND2X1_LOC_114/a_36_24# NAND2X1_LOC_116/A VSS VDD INVX1_LOC_65/Y
+ NAND2X1_LOC_114/B NAND2X1_LOC
XNAND2X1_LOC_125 NAND2X1_LOC_125/a_36_24# NOR2X1_LOC_128/B VSS VDD INVX1_LOC_57/A
+ INVX1_LOC_63/A NAND2X1_LOC
XNAND2X1_LOC_103 NAND2X1_LOC_103/a_36_24# NOR2X1_LOC_113/B VSS VDD INVX1_LOC_35/A
+ NOR2X1_LOC_590/A NAND2X1_LOC
XNAND2X1_LOC_136 NAND2X1_LOC_136/a_36_24# NOR2X1_LOC_514/A VSS VDD INVX1_LOC_1/A INVX1_LOC_31/A
+ NAND2X1_LOC
XNAND2X1_LOC_169 NAND2X1_LOC_169/a_36_24# NAND2X1_LOC_169/Y VSS VDD NOR2X1_LOC_166/Y
+ NOR2X1_LOC_167/Y NAND2X1_LOC
XNAND2X1_LOC_147 NAND2X1_LOC_147/a_36_24# INVX1_LOC_85/A VSS VDD NOR2X1_LOC_142/Y
+ NOR2X1_LOC_144/Y NAND2X1_LOC
XNAND2X1_LOC_158 NAND2X1_LOC_158/a_36_24# NOR2X1_LOC_210/B VSS VDD NOR2X1_LOC_156/Y
+ INVX1_LOC_89/A NAND2X1_LOC
XNAND2X1_LOC_1 NAND2X1_LOC_1/a_36_24# NAND2X1_LOC_1/Y VSS VDD D_INPUT_6 INPUT_7
+ NAND2X1_LOC
XNOR2X1_LOC_180 NOR2X1_LOC_180/a_36_216# NOR2X1_LOC_180/Y VSS VDD NOR2X1_LOC_439/B
+ NOR2X1_LOC_180/B NOR2X1_LOC
XNOR2X1_LOC_191 NOR2X1_LOC_191/a_36_216# NOR2X1_LOC_192/A VSS VDD NOR2X1_LOC_191/A
+ NOR2X1_LOC_191/B NOR2X1_LOC
XNAND2X1_LOC_670 NAND2X1_LOC_670/a_36_24# NOR2X1_LOC_673/B VSS VDD INVX1_LOC_29/A
+ NOR2X1_LOC_590/A NAND2X1_LOC
XNAND2X1_LOC_681 NAND2X1_LOC_681/a_36_24# NOR2X1_LOC_685/B VSS VDD INVX1_LOC_21/A
+ NOR2X1_LOC_155/A NAND2X1_LOC
XINVX1_LOC_60 INVX1_LOC_60/Y VSS VDD INVX1_LOC_60/A INVX1_LOC
XNAND2X1_LOC_692 NAND2X1_LOC_692/a_36_24# NOR2X1_LOC_706/B VSS VDD INVX1_LOC_15/A
+ NOR2X1_LOC_598/B NAND2X1_LOC
XINVX1_LOC_82 INVX1_LOC_82/Y VSS VDD INVX1_LOC_82/A INVX1_LOC
XINVX1_LOC_71 INVX1_LOC_71/Y VSS VDD INVX1_LOC_71/A INVX1_LOC
XINVX1_LOC_93 INVX1_LOC_93/Y VSS VDD INVX1_LOC_93/A INVX1_LOC
XNOR2X1_LOC_4 NOR2X1_LOC_4/a_36_216# NOR2X1_LOC_6/B VSS VDD INPUT_1 D_INPUT_0
+ NOR2X1_LOC
XINVX1_LOC_300 INVX1_LOC_300/Y VSS VDD INVX1_LOC_300/A INVX1_LOC
XINVX1_LOC_311 INVX1_LOC_311/Y VSS VDD INVX1_LOC_311/A INVX1_LOC
XNOR2X1_LOC_713 NOR2X1_LOC_713/a_36_216# NOR2X1_LOC_725/A VSS VDD NOR2X1_LOC_706/Y
+ NOR2X1_LOC_713/B NOR2X1_LOC
XNOR2X1_LOC_735 NOR2X1_LOC_735/a_36_216# NOR2X1_LOC_735/Y VSS VDD NOR2X1_LOC_632/Y
+ INVX1_LOC_208/A NOR2X1_LOC
XNOR2X1_LOC_724 NOR2X1_LOC_724/a_36_216# NOR2X1_LOC_724/Y VSS VDD INVX1_LOC_279/Y
+ NOR2X1_LOC_714/Y NOR2X1_LOC
XNOR2X1_LOC_702 NOR2X1_LOC_702/a_36_216# NOR2X1_LOC_702/Y VSS VDD NOR2X1_LOC_332/A
+ NAND2X1_LOC_45/Y NOR2X1_LOC
XNOR2X1_LOC_746 NOR2X1_LOC_746/a_36_216# NOR2X1_LOC_746/Y VSS VDD INVX1_LOC_90/A NOR2X1_LOC_74/A
+ NOR2X1_LOC
XNOR2X1_LOC_779 NOR2X1_LOC_779/a_36_216# NOR2X1_LOC_779/Y VSS VDD NOR2X1_LOC_708/A
+ INVX1_LOC_213/A NOR2X1_LOC
XNOR2X1_LOC_757 NOR2X1_LOC_757/a_36_216# NOR2X1_LOC_757/Y VSS VDD NOR2X1_LOC_757/A
+ INVX1_LOC_34/A NOR2X1_LOC
XNOR2X1_LOC_768 NOR2X1_LOC_768/a_36_216# NOR2X1_LOC_772/A VSS VDD NOR2X1_LOC_137/A
+ NOR2X1_LOC_113/B NOR2X1_LOC
XINVX1_LOC_152 INVX1_LOC_152/Y VSS VDD INVX1_LOC_152/A INVX1_LOC
XINVX1_LOC_141 INVX1_LOC_141/Y VSS VDD INVX1_LOC_141/A INVX1_LOC
XINVX1_LOC_130 INVX1_LOC_130/Y VSS VDD INVX1_LOC_130/A INVX1_LOC
XINVX1_LOC_163 INVX1_LOC_163/Y VSS VDD INVX1_LOC_163/A INVX1_LOC
XINVX1_LOC_185 INVX1_LOC_185/Y VSS VDD INVX1_LOC_185/A INVX1_LOC
XINVX1_LOC_196 INVX1_LOC_196/Y VSS VDD INVX1_LOC_196/A INVX1_LOC
XINVX1_LOC_174 INVX1_LOC_174/Y VSS VDD INVX1_LOC_174/A INVX1_LOC
XNOR2X1_LOC_510 NOR2X1_LOC_510/a_36_216# NOR2X1_LOC_510/Y VSS VDD INVX1_LOC_211/Y
+ NOR2X1_LOC_510/B NOR2X1_LOC
XNOR2X1_LOC_565 NOR2X1_LOC_565/a_36_216# NOR2X1_LOC_569/A VSS VDD NOR2X1_LOC_565/A
+ NOR2X1_LOC_565/B NOR2X1_LOC
XNOR2X1_LOC_543 NOR2X1_LOC_543/a_36_216# NOR2X1_LOC_552/A VSS VDD NOR2X1_LOC_543/A
+ NOR2X1_LOC_318/B NOR2X1_LOC
XNOR2X1_LOC_532 NOR2X1_LOC_532/a_36_216# NOR2X1_LOC_532/Y VSS VDD INVX1_LOC_75/A NOR2X1_LOC_590/A
+ NOR2X1_LOC
XNOR2X1_LOC_554 NOR2X1_LOC_554/a_36_216# INVX1_LOC_228/A VSS VDD NOR2X1_LOC_554/A
+ NOR2X1_LOC_554/B NOR2X1_LOC
XNOR2X1_LOC_521 NOR2X1_LOC_521/a_36_216# NOR2X1_LOC_521/Y VSS VDD NOR2X1_LOC_52/B
+ INVX1_LOC_15/Y NOR2X1_LOC
XNOR2X1_LOC_576 NOR2X1_LOC_576/a_36_216# INVX1_LOC_238/A VSS VDD INVX1_LOC_233/Y NOR2X1_LOC_576/B
+ NOR2X1_LOC
XNOR2X1_LOC_587 NOR2X1_LOC_587/a_36_216# NOR2X1_LOC_588/A VSS VDD NOR2X1_LOC_30/Y
+ INPUT_7 NOR2X1_LOC
XNOR2X1_LOC_598 NOR2X1_LOC_598/a_36_216# NOR2X1_LOC_828/A VSS VDD INVX1_LOC_135/A
+ NOR2X1_LOC_598/B NOR2X1_LOC
XNAND2X1_LOC_318 NAND2X1_LOC_318/a_36_24# INVX1_LOC_143/A VSS VDD NOR2X1_LOC_315/Y
+ NOR2X1_LOC_316/Y NAND2X1_LOC
XNAND2X1_LOC_307 NAND2X1_LOC_307/a_36_24# NAND2X1_LOC_308/B VSS VDD NOR2X1_LOC_304/Y
+ NOR2X1_LOC_305/Y NAND2X1_LOC
XNAND2X1_LOC_329 NAND2X1_LOC_329/a_36_24# NOR2X1_LOC_355/B VSS VDD NOR2X1_LOC_405/A
+ NOR2X1_LOC_596/A NAND2X1_LOC
XNOR2X1_LOC_351 NOR2X1_LOC_351/a_36_216# NOR2X1_LOC_351/Y VSS VDD INVX1_LOC_151/Y
+ NOR2X1_LOC_338/Y NOR2X1_LOC
XNOR2X1_LOC_362 NOR2X1_LOC_362/a_36_216# NOR2X1_LOC_366/B VSS VDD NOR2X1_LOC_361/Y
+ INVX1_LOC_133/Y NOR2X1_LOC
XNOR2X1_LOC_395 NOR2X1_LOC_395/a_36_216# NOR2X1_LOC_395/Y VSS VDD INVX1_LOC_64/A INVX1_LOC_46/A
+ NOR2X1_LOC
XNOR2X1_LOC_340 NOR2X1_LOC_340/a_36_216# NOR2X1_LOC_340/Y VSS VDD NOR2X1_LOC_340/A
+ NOR2X1_LOC_100/A NOR2X1_LOC
XNOR2X1_LOC_384 NOR2X1_LOC_384/a_36_216# NOR2X1_LOC_384/Y VSS VDD NOR2X1_LOC_384/A
+ INVX1_LOC_30/A NOR2X1_LOC
XNOR2X1_LOC_373 NOR2X1_LOC_373/a_36_216# NOR2X1_LOC_373/Y VSS VDD NOR2X1_LOC_89/A
+ INVX1_LOC_19/Y NOR2X1_LOC
XNAND2X1_LOC_852 NAND2X1_LOC_852/a_36_24# NAND2X1_LOC_852/Y VSS VDD NAND2X1_LOC_838/Y
+ NAND2X1_LOC_839/Y NAND2X1_LOC
XNAND2X1_LOC_863 NAND2X1_LOC_863/a_36_24# NAND2X1_LOC_863/Y VSS VDD NAND2X1_LOC_863/A
+ NAND2X1_LOC_863/B NAND2X1_LOC
XNAND2X1_LOC_830 NAND2X1_LOC_830/a_36_24# NAND2X1_LOC_842/B VSS VDD INVX1_LOC_66/A
+ NOR2X1_LOC_142/Y NAND2X1_LOC
XNAND2X1_LOC_841 NAND2X1_LOC_841/a_36_24# INVX1_LOC_311/A VSS VDD NAND2X1_LOC_841/A
+ NAND2X1_LOC_832/Y NAND2X1_LOC
XNOR2X1_LOC_80 NOR2X1_LOC_80/a_36_216# NOR2X1_LOC_80/Y VSS VDD NOR2X1_LOC_82/A INVX1_LOC_4/A
+ NOR2X1_LOC
XNOR2X1_LOC_91 NOR2X1_LOC_91/a_36_216# NOR2X1_LOC_91/Y VSS VDD NOR2X1_LOC_91/A INVX1_LOC_38/A
+ NOR2X1_LOC
XNAND2X1_LOC_137 NAND2X1_LOC_137/a_36_24# NAND2X1_LOC_139/A VSS VDD NOR2X1_LOC_132/Y
+ NOR2X1_LOC_134/Y NAND2X1_LOC
XNAND2X1_LOC_159 NAND2X1_LOC_159/a_36_24# INVX1_LOC_91/A VSS VDD INVX1_LOC_3/A NAND2X1_LOC_9/Y
+ NAND2X1_LOC
XNAND2X1_LOC_126 NAND2X1_LOC_126/a_36_24# INVX1_LOC_75/A VSS VDD NOR2X1_LOC_19/B INVX1_LOC_25/A
+ NAND2X1_LOC
XNAND2X1_LOC_104 NAND2X1_LOC_104/a_36_24# INVX1_LOC_63/A VSS VDD NOR2X1_LOC_19/B INVX1_LOC_7/A
+ NAND2X1_LOC
XNAND2X1_LOC_115 NAND2X1_LOC_115/a_36_24# INVX1_LOC_67/A VSS VDD NOR2X1_LOC_106/Y
+ NAND2X1_LOC_112/Y NAND2X1_LOC
XNAND2X1_LOC_148 NAND2X1_LOC_148/a_36_24# NAND2X1_LOC_149/B VSS VDD NOR2X1_LOC_145/Y
+ NOR2X1_LOC_146/Y NAND2X1_LOC
XNAND2X1_LOC_2 NAND2X1_LOC_2/a_36_24# NAND2X1_LOC_3/B VSS VDD D_INPUT_4 D_INPUT_5
+ NAND2X1_LOC
XNOR2X1_LOC_181 NOR2X1_LOC_181/a_36_216# NOR2X1_LOC_181/Y VSS VDD NOR2X1_LOC_181/A
+ NOR2X1_LOC_540/B NOR2X1_LOC
XNOR2X1_LOC_170 NOR2X1_LOC_170/a_36_216# INVX1_LOC_94/A VSS VDD NOR2X1_LOC_170/A NOR2X1_LOC_168/Y
+ NOR2X1_LOC
XNOR2X1_LOC_192 NOR2X1_LOC_192/a_36_216# INVX1_LOC_104/A VSS VDD NOR2X1_LOC_192/A
+ INVX1_LOC_102/Y NOR2X1_LOC
XNAND2X1_LOC_671 NAND2X1_LOC_671/a_36_24# NAND2X1_LOC_672/B VSS VDD INPUT_2 NOR2X1_LOC_19/B
+ NAND2X1_LOC
XNAND2X1_LOC_660 NAND2X1_LOC_660/a_36_24# NAND2X1_LOC_660/Y VSS VDD NAND2X1_LOC_660/A
+ NAND2X1_LOC_656/Y NAND2X1_LOC
XNAND2X1_LOC_693 NAND2X1_LOC_693/a_36_24# NOR2X1_LOC_706/A VSS VDD INVX1_LOC_14/Y
+ INVX1_LOC_23/A NAND2X1_LOC
XNAND2X1_LOC_682 NAND2X1_LOC_682/a_36_24# NOR2X1_LOC_685/A VSS VDD INVX1_LOC_23/A
+ INVX1_LOC_91/A NAND2X1_LOC
XINVX1_LOC_61 INVX1_LOC_61/Y VSS VDD INVX1_LOC_61/A INVX1_LOC
XINVX1_LOC_72 INVX1_LOC_72/Y VSS VDD INVX1_LOC_72/A INVX1_LOC
XINVX1_LOC_94 INVX1_LOC_94/Y VSS VDD INVX1_LOC_94/A INVX1_LOC
XINVX1_LOC_50 INVX1_LOC_50/Y VSS VDD INVX1_LOC_50/A INVX1_LOC
XINVX1_LOC_83 INVX1_LOC_83/Y VSS VDD INVX1_LOC_83/A INVX1_LOC
XNOR2X1_LOC_5 NOR2X1_LOC_5/a_36_216# INVX1_LOC_4/A VSS VDD D_INPUT_3 INPUT_2 NOR2X1_LOC
XNAND2X1_LOC_490 NAND2X1_LOC_490/a_36_24# NOR2X1_LOC_557/A VSS VDD NOR2X1_LOC_6/B
+ NAND2X1_LOC_85/Y NAND2X1_LOC
XINVX1_LOC_312 INVX1_LOC_312/Y VSS VDD INVX1_LOC_312/A INVX1_LOC
XINVX1_LOC_301 INVX1_LOC_301/Y VSS VDD INVX1_LOC_301/A INVX1_LOC
XNOR2X1_LOC_725 NOR2X1_LOC_725/a_36_216# NOR2X1_LOC_732/A VSS VDD NOR2X1_LOC_725/A
+ NOR2X1_LOC_712/Y NOR2X1_LOC
XNOR2X1_LOC_769 NOR2X1_LOC_769/a_36_216# INVX1_LOC_296/A VSS VDD NOR2X1_LOC_769/A
+ NOR2X1_LOC_769/B NOR2X1_LOC
XNOR2X1_LOC_747 NOR2X1_LOC_747/a_36_216# INVX1_LOC_288/A VSS VDD NOR2X1_LOC_52/B INVX1_LOC_36/A
+ NOR2X1_LOC
XNOR2X1_LOC_736 NOR2X1_LOC_736/a_36_216# NOR2X1_LOC_736/Y VSS VDD NOR2X1_LOC_735/Y
+ INVX1_LOC_270/A NOR2X1_LOC
XNOR2X1_LOC_714 NOR2X1_LOC_714/a_36_216# NOR2X1_LOC_714/Y VSS VDD NOR2X1_LOC_704/Y
+ NOR2X1_LOC_703/Y NOR2X1_LOC
XNOR2X1_LOC_703 NOR2X1_LOC_703/a_36_216# NOR2X1_LOC_703/Y VSS VDD NOR2X1_LOC_703/A
+ NOR2X1_LOC_703/B NOR2X1_LOC
XNOR2X1_LOC_758 NOR2X1_LOC_758/a_36_216# NOR2X1_LOC_758/Y VSS VDD INVX1_LOC_57/A INVX1_LOC_29/A
+ NOR2X1_LOC
XINVX1_LOC_175 INVX1_LOC_175/Y VSS VDD INVX1_LOC_175/A INVX1_LOC
XINVX1_LOC_120 INVX1_LOC_120/Y VSS VDD INVX1_LOC_120/A INVX1_LOC
XINVX1_LOC_164 INVX1_LOC_164/Y VSS VDD INVX1_LOC_164/A INVX1_LOC
XINVX1_LOC_131 INVX1_LOC_131/Y VSS VDD INVX1_LOC_131/A INVX1_LOC
XINVX1_LOC_186 INVX1_LOC_186/Y VSS VDD INVX1_LOC_186/A INVX1_LOC
XINVX1_LOC_142 INVX1_LOC_142/Y VSS VDD INVX1_LOC_142/A INVX1_LOC
XINVX1_LOC_153 INVX1_LOC_153/Y VSS VDD INVX1_LOC_153/A INVX1_LOC
XINVX1_LOC_197 INVX1_LOC_197/Y VSS VDD INVX1_LOC_197/A INVX1_LOC
XNOR2X1_LOC_588 NOR2X1_LOC_588/a_36_216# INVX1_LOC_244/A VSS VDD NOR2X1_LOC_588/A
+ INVX1_LOC_84/A NOR2X1_LOC
XNOR2X1_LOC_555 NOR2X1_LOC_555/a_36_216# NOR2X1_LOC_562/B VSS VDD INVX1_LOC_206/Y
+ INVX1_LOC_121/Y NOR2X1_LOC
XNOR2X1_LOC_599 NOR2X1_LOC_599/a_36_216# NOR2X1_LOC_599/Y VSS VDD NOR2X1_LOC_599/A
+ INVX1_LOC_24/A NOR2X1_LOC
XNOR2X1_LOC_544 NOR2X1_LOC_544/a_36_216# NOR2X1_LOC_551/B VSS VDD NOR2X1_LOC_544/A
+ NOR2X1_LOC_374/A NOR2X1_LOC
XNOR2X1_LOC_511 NOR2X1_LOC_511/a_36_216# INVX1_LOC_214/A VSS VDD NOR2X1_LOC_48/B INVX1_LOC_21/Y
+ NOR2X1_LOC
XNOR2X1_LOC_577 NOR2X1_LOC_577/a_36_216# NOR2X1_LOC_577/Y VSS VDD NOR2X1_LOC_570/Y
+ NOR2X1_LOC_569/Y NOR2X1_LOC
XNOR2X1_LOC_533 NOR2X1_LOC_533/a_36_216# NOR2X1_LOC_533/Y VSS VDD NOR2X1_LOC_533/A
+ INVX1_LOC_58/A NOR2X1_LOC
XNOR2X1_LOC_500 NOR2X1_LOC_500/a_36_216# NOR2X1_LOC_500/Y VSS VDD NOR2X1_LOC_500/A
+ NOR2X1_LOC_500/B NOR2X1_LOC
XNOR2X1_LOC_566 NOR2X1_LOC_566/a_36_216# NOR2X1_LOC_566/Y VSS VDD NOR2X1_LOC_303/Y
+ INVX1_LOC_93/Y NOR2X1_LOC
XNOR2X1_LOC_522 NOR2X1_LOC_522/a_36_216# NOR2X1_LOC_522/Y VSS VDD NOR2X1_LOC_536/A
+ INVX1_LOC_18/A NOR2X1_LOC
XNAND2X1_LOC_308 NAND2X1_LOC_308/a_36_24# NAND2X1_LOC_308/Y VSS VDD INVX1_LOC_141/Y
+ NAND2X1_LOC_308/B NAND2X1_LOC
XNAND2X1_LOC_319 NAND2X1_LOC_319/a_36_24# NAND2X1_LOC_798/A VSS VDD NAND2X1_LOC_319/A
+ INVX1_LOC_144/Y NAND2X1_LOC
XNOR2X1_LOC_330 NOR2X1_LOC_330/a_36_216# INVX1_LOC_146/A VSS VDD INVX1_LOC_53/A INVX1_LOC_37/A
+ NOR2X1_LOC
XNOR2X1_LOC_352 NOR2X1_LOC_352/a_36_216# NOR2X1_LOC_352/Y VSS VDD NOR2X1_LOC_337/Y
+ INVX1_LOC_96/A NOR2X1_LOC
XNOR2X1_LOC_363 NOR2X1_LOC_363/a_36_216# NOR2X1_LOC_363/Y VSS VDD NOR2X1_LOC_360/Y
+ NOR2X1_LOC_359/Y NOR2X1_LOC
XNOR2X1_LOC_374 NOR2X1_LOC_374/a_36_216# NOR2X1_LOC_717/B VSS VDD NOR2X1_LOC_374/A
+ NOR2X1_LOC_374/B NOR2X1_LOC
XNOR2X1_LOC_385 NOR2X1_LOC_385/a_36_216# NOR2X1_LOC_385/Y VSS VDD INVX1_LOC_64/A INVX1_LOC_20/A
+ NOR2X1_LOC
XNOR2X1_LOC_396 NOR2X1_LOC_396/a_36_216# NOR2X1_LOC_396/Y VSS VDD INVX1_LOC_24/A NOR2X1_LOC_45/B
+ NOR2X1_LOC
XNOR2X1_LOC_341 NOR2X1_LOC_341/a_36_216# NOR2X1_LOC_350/A VSS VDD NOR2X1_LOC_641/B
+ NOR2X1_LOC_716/B NOR2X1_LOC
XNAND2X1_LOC_820 NAND2X1_LOC_820/a_36_24# NOR2X1_LOC_847/A VSS VDD NOR2X1_LOC_818/Y
+ NAND2X1_LOC_819/Y NAND2X1_LOC
XNAND2X1_LOC_842 NAND2X1_LOC_842/a_36_24# NAND2X1_LOC_850/A VSS VDD INVX1_LOC_100/A
+ NAND2X1_LOC_842/B NAND2X1_LOC
XNAND2X1_LOC_853 NAND2X1_LOC_853/a_36_24# NAND2X1_LOC_853/Y VSS VDD NAND2X1_LOC_35/Y
+ NAND2X1_LOC_175/Y NAND2X1_LOC
XNAND2X1_LOC_864 NAND2X1_LOC_864/a_36_24# NAND2X1_LOC_866/A VSS VDD INVX1_LOC_300/Y
+ NAND2X1_LOC_863/Y NAND2X1_LOC
XNAND2X1_LOC_831 NAND2X1_LOC_831/a_36_24# NAND2X1_LOC_841/A VSS VDD NOR2X1_LOC_273/Y
+ NOR2X1_LOC_300/Y NAND2X1_LOC
XNOR2X1_LOC_70 NOR2X1_LOC_70/a_36_216# INVX1_LOC_54/A VSS VDD NOR2X1_LOC_51/A NOR2X1_LOC_2/Y
+ NOR2X1_LOC
XNOR2X1_LOC_92 NOR2X1_LOC_92/a_36_216# NOR2X1_LOC_92/Y VSS VDD INVX1_LOC_8/A D_INPUT_1
+ NOR2X1_LOC
XNOR2X1_LOC_81 NOR2X1_LOC_81/a_36_216# NOR2X1_LOC_81/Y VSS VDD NOR2X1_LOC_80/Y INVX1_LOC_46/A
+ NOR2X1_LOC
XNAND2X1_LOC_127 NAND2X1_LOC_127/a_36_24# NOR2X1_LOC_128/A VSS VDD INVX1_LOC_1/A INVX1_LOC_75/A
+ NAND2X1_LOC
XNAND2X1_LOC_116 NAND2X1_LOC_116/a_36_24# NAND2X1_LOC_473/A VSS VDD NAND2X1_LOC_116/A
+ INVX1_LOC_68/Y NAND2X1_LOC
XNAND2X1_LOC_105 NAND2X1_LOC_105/a_36_24# NOR2X1_LOC_106/A VSS VDD NOR2X1_LOC_89/A
+ INVX1_LOC_64/A NAND2X1_LOC
XNAND2X1_LOC_138 NAND2X1_LOC_138/a_36_24# INVX1_LOC_79/A VSS VDD NOR2X1_LOC_135/Y
+ NOR2X1_LOC_136/Y NAND2X1_LOC
XNAND2X1_LOC_149 NAND2X1_LOC_149/a_36_24# NAND2X1_LOC_149/Y VSS VDD INVX1_LOC_86/Y
+ NAND2X1_LOC_149/B NAND2X1_LOC
XNAND2X1_LOC_3 NAND2X1_LOC_3/a_36_24# INVX1_LOC_1/A VSS VDD NAND2X1_LOC_1/Y NAND2X1_LOC_3/B
+ NAND2X1_LOC
XNOR2X1_LOC_160 NOR2X1_LOC_160/a_36_216# NOR2X1_LOC_160/Y VSS VDD INVX1_LOC_75/A NOR2X1_LOC_160/B
+ NOR2X1_LOC
XNOR2X1_LOC_182 NOR2X1_LOC_182/a_36_216# INVX1_LOC_96/A VSS VDD NOR2X1_LOC_181/Y NOR2X1_LOC_180/Y
+ NOR2X1_LOC
XNOR2X1_LOC_171 NOR2X1_LOC_171/a_36_216# NOR2X1_LOC_171/Y VSS VDD INVX1_LOC_30/A NOR2X1_LOC_45/B
+ NOR2X1_LOC
XNOR2X1_LOC_193 NOR2X1_LOC_193/a_36_216# INVX1_LOC_106/A VSS VDD NOR2X1_LOC_538/B
+ NAND2X1_LOC_7/Y NOR2X1_LOC
XNAND2X1_LOC_672 NAND2X1_LOC_672/a_36_24# NOR2X1_LOC_673/A VSS VDD INVX1_LOC_89/A
+ NAND2X1_LOC_672/B NAND2X1_LOC
XNAND2X1_LOC_650 NAND2X1_LOC_650/a_36_24# INVX1_LOC_265/A VSS VDD NAND2X1_LOC_640/Y
+ NAND2X1_LOC_650/B NAND2X1_LOC
XNAND2X1_LOC_683 NAND2X1_LOC_683/a_36_24# NOR2X1_LOC_686/B VSS VDD NOR2X1_LOC_78/B
+ INVX1_LOC_17/A NAND2X1_LOC
XNAND2X1_LOC_661 NAND2X1_LOC_661/a_36_24# NAND2X1_LOC_662/B VSS VDD NAND2X1_LOC_661/A
+ NAND2X1_LOC_661/B NAND2X1_LOC
XNAND2X1_LOC_694 NAND2X1_LOC_694/a_36_24# NOR2X1_LOC_707/B VSS VDD INVX1_LOC_77/A
+ NAND2X1_LOC_425/Y NAND2X1_LOC
XINVX1_LOC_84 INVX1_LOC_84/Y VSS VDD INVX1_LOC_84/A INVX1_LOC
XINVX1_LOC_40 INVX1_LOC_40/Y VSS VDD INVX1_LOC_40/A INVX1_LOC
XINVX1_LOC_62 INVX1_LOC_62/Y VSS VDD INVX1_LOC_62/A INVX1_LOC
XINVX1_LOC_51 INVX1_LOC_51/Y VSS VDD INVX1_LOC_51/A INVX1_LOC
XINVX1_LOC_95 INVX1_LOC_95/Y VSS VDD INVX1_LOC_95/A INVX1_LOC
XINVX1_LOC_73 INVX1_LOC_73/Y VSS VDD INVX1_LOC_73/A INVX1_LOC
XNOR2X1_LOC_6 NOR2X1_LOC_6/a_36_216# INVX1_LOC_6/A VSS VDD INVX1_LOC_4/A NOR2X1_LOC_6/B
+ NOR2X1_LOC
XNAND2X1_LOC_491 NAND2X1_LOC_491/a_36_24# NOR2X1_LOC_493/B VSS VDD INVX1_LOC_21/A
+ NOR2X1_LOC_590/A NAND2X1_LOC
XNAND2X1_LOC_480 NAND2X1_LOC_480/a_36_24# GATE_479 VSS VDD INVX1_LOC_204/Y NAND2X1_LOC_479/Y
+ NAND2X1_LOC
XINVX1_LOC_313 INVX1_LOC_313/Y VSS VDD INVX1_LOC_313/A INVX1_LOC
XINVX1_LOC_302 INVX1_LOC_302/Y VSS VDD INVX1_LOC_302/A INVX1_LOC
XNOR2X1_LOC_737 NOR2X1_LOC_737/a_36_216# NOR2X1_LOC_741/A VSS VDD INVX1_LOC_285/Y
+ NOR2X1_LOC_733/Y NOR2X1_LOC
XNOR2X1_LOC_726 NOR2X1_LOC_726/a_36_216# NOR2X1_LOC_726/Y VSS VDD NOR2X1_LOC_711/Y
+ NOR2X1_LOC_209/A NOR2X1_LOC
XNOR2X1_LOC_759 NOR2X1_LOC_759/a_36_216# NOR2X1_LOC_759/Y VSS VDD NOR2X1_LOC_759/A
+ INVX1_LOC_117/Y NOR2X1_LOC
XNOR2X1_LOC_704 NOR2X1_LOC_704/a_36_216# NOR2X1_LOC_704/Y VSS VDD INVX1_LOC_177/A
+ NOR2X1_LOC_317/B NOR2X1_LOC
XNOR2X1_LOC_748 NOR2X1_LOC_748/a_36_216# NOR2X1_LOC_748/Y VSS VDD NOR2X1_LOC_748/A
+ NOR2X1_LOC_6/B NOR2X1_LOC
XNOR2X1_LOC_715 NOR2X1_LOC_715/a_36_216# INVX1_LOC_280/A VSS VDD NOR2X1_LOC_702/Y
+ NOR2X1_LOC_112/Y NOR2X1_LOC
XINVX1_LOC_154 INVX1_LOC_154/Y VSS VDD INVX1_LOC_154/A INVX1_LOC
XINVX1_LOC_110 INVX1_LOC_110/Y VSS VDD INVX1_LOC_110/A INVX1_LOC
XINVX1_LOC_176 INVX1_LOC_176/Y VSS VDD INVX1_LOC_176/A INVX1_LOC
XINVX1_LOC_165 INVX1_LOC_165/Y VSS VDD INVX1_LOC_165/A INVX1_LOC
XINVX1_LOC_132 INVX1_LOC_132/Y VSS VDD INVX1_LOC_132/A INVX1_LOC
XINVX1_LOC_143 INVX1_LOC_143/Y VSS VDD INVX1_LOC_143/A INVX1_LOC
XINVX1_LOC_187 INVX1_LOC_187/Y VSS VDD INVX1_LOC_187/A INVX1_LOC
XINVX1_LOC_198 INVX1_LOC_198/Y VSS VDD INVX1_LOC_198/A INVX1_LOC
XINVX1_LOC_121 INVX1_LOC_121/Y VSS VDD INVX1_LOC_121/A INVX1_LOC
XNOR2X1_LOC_501 NOR2X1_LOC_501/a_36_216# INVX1_LOC_208/A VSS VDD NOR2X1_LOC_500/Y
+ NOR2X1_LOC_501/B NOR2X1_LOC
XNOR2X1_LOC_589 NOR2X1_LOC_589/a_36_216# NOR2X1_LOC_589/Y VSS VDD NOR2X1_LOC_589/A
+ INVX1_LOC_18/A NOR2X1_LOC
XNOR2X1_LOC_556 NOR2X1_LOC_556/a_36_216# NOR2X1_LOC_562/A VSS VDD NOR2X1_LOC_486/Y
+ NOR2X1_LOC_631/B NOR2X1_LOC
XNOR2X1_LOC_578 NOR2X1_LOC_578/a_36_216# INVX1_LOC_240/A VSS VDD NOR2X1_LOC_577/Y
+ INVX1_LOC_231/Y NOR2X1_LOC
XNOR2X1_LOC_512 NOR2X1_LOC_512/a_36_216# NOR2X1_LOC_512/Y VSS VDD INVX1_LOC_141/A
+ D_INPUT_0 NOR2X1_LOC
XNOR2X1_LOC_534 NOR2X1_LOC_534/a_36_216# INVX1_LOC_222/A VSS VDD INVX1_LOC_46/A INVX1_LOC_32/A
+ NOR2X1_LOC
XNOR2X1_LOC_567 NOR2X1_LOC_567/a_36_216# NOR2X1_LOC_568/A VSS VDD NOR2X1_LOC_799/B
+ NOR2X1_LOC_567/B NOR2X1_LOC
XNOR2X1_LOC_523 NOR2X1_LOC_523/a_36_216# NOR2X1_LOC_844/A VSS VDD NOR2X1_LOC_523/A
+ NOR2X1_LOC_523/B NOR2X1_LOC
XNOR2X1_LOC_545 NOR2X1_LOC_545/a_36_216# INVX1_LOC_224/A VSS VDD NOR2X1_LOC_545/A
+ NOR2X1_LOC_545/B NOR2X1_LOC
XNAND2X1_LOC_309 NAND2X1_LOC_309/a_36_24# NOR2X1_LOC_335/B VSS VDD INVX1_LOC_17/A
+ NOR2X1_LOC_814/A NAND2X1_LOC
XNOR2X1_LOC_331 NOR2X1_LOC_331/a_36_216# NOR2X1_LOC_331/Y VSS VDD INVX1_LOC_146/Y
+ NOR2X1_LOC_331/B NOR2X1_LOC
XNOR2X1_LOC_320 NOR2X1_LOC_320/a_36_216# NOR2X1_LOC_320/Y VSS VDD NOR2X1_LOC_91/A
+ INVX1_LOC_24/A NOR2X1_LOC
XNOR2X1_LOC_342 NOR2X1_LOC_342/a_36_216# NOR2X1_LOC_349/B VSS VDD NOR2X1_LOC_342/A
+ NOR2X1_LOC_342/B NOR2X1_LOC
XNOR2X1_LOC_386 NOR2X1_LOC_386/a_36_216# NOR2X1_LOC_387/A VSS VDD NOR2X1_LOC_36/B
+ INPUT_4 NOR2X1_LOC
XNOR2X1_LOC_364 NOR2X1_LOC_364/a_36_216# NOR2X1_LOC_364/Y VSS VDD NOR2X1_LOC_364/A
+ NOR2X1_LOC_357/Y NOR2X1_LOC
XNOR2X1_LOC_353 NOR2X1_LOC_353/a_36_216# NOR2X1_LOC_353/Y VSS VDD NOR2X1_LOC_727/B
+ NOR2X1_LOC_303/Y NOR2X1_LOC
XNOR2X1_LOC_375 NOR2X1_LOC_375/a_36_216# NOR2X1_LOC_375/Y VSS VDD INVX1_LOC_89/A INVX1_LOC_21/A
+ NOR2X1_LOC
XNOR2X1_LOC_397 NOR2X1_LOC_397/a_36_216# INVX1_LOC_164/A VSS VDD NOR2X1_LOC_82/Y INVX1_LOC_1/Y
+ NOR2X1_LOC
XNAND2X1_LOC_865 NAND2X1_LOC_865/a_36_24# NAND2X1_LOC_866/B VSS VDD NAND2X1_LOC_861/Y
+ NAND2X1_LOC_862/Y NAND2X1_LOC
XNAND2X1_LOC_821 NAND2X1_LOC_821/a_36_24# NOR2X1_LOC_835/B VSS VDD INVX1_LOC_9/A INVX1_LOC_53/A
+ NAND2X1_LOC
XNAND2X1_LOC_843 NAND2X1_LOC_843/a_36_24# INVX1_LOC_313/A VSS VDD NOR2X1_LOC_251/Y
+ NOR2X1_LOC_278/Y NAND2X1_LOC
XNAND2X1_LOC_854 NAND2X1_LOC_854/a_36_24# NAND2X1_LOC_856/A VSS VDD NAND2X1_LOC_354/B
+ NAND2X1_LOC_854/B NAND2X1_LOC
XNAND2X1_LOC_810 NAND2X1_LOC_810/a_36_24# NAND2X1_LOC_812/A VSS VDD INVX1_LOC_300/Y
+ NAND2X1_LOC_810/B NAND2X1_LOC
XNAND2X1_LOC_832 NAND2X1_LOC_832/a_36_24# NAND2X1_LOC_832/Y VSS VDD NOR2X1_LOC_423/Y
+ NOR2X1_LOC_433/Y NAND2X1_LOC
XNOR2X1_LOC_60 NOR2X1_LOC_60/a_36_216# NOR2X1_LOC_60/Y VSS VDD INVX1_LOC_46/A INVX1_LOC_28/A
+ NOR2X1_LOC
XNOR2X1_LOC_71 NOR2X1_LOC_71/a_36_216# NOR2X1_LOC_71/Y VSS VDD INVX1_LOC_47/Y INVX1_LOC_4/A
+ NOR2X1_LOC
XNOR2X1_LOC_82 NOR2X1_LOC_82/a_36_216# NOR2X1_LOC_82/Y VSS VDD NOR2X1_LOC_82/A INVX1_LOC_14/A
+ NOR2X1_LOC
XNOR2X1_LOC_93 NOR2X1_LOC_93/a_36_216# NOR2X1_LOC_93/Y VSS VDD NOR2X1_LOC_92/Y INVX1_LOC_20/A
+ NOR2X1_LOC
XNAND2X1_LOC_117 NAND2X1_LOC_117/a_36_24# NOR2X1_LOC_123/B VSS VDD NAND2X1_LOC_63/Y
+ INVX1_LOC_54/Y NAND2X1_LOC
XNAND2X1_LOC_4 NAND2X1_LOC_4/a_36_24# NOR2X1_LOC_19/B VSS VDD INPUT_0 D_INPUT_1
+ NAND2X1_LOC
XNAND2X1_LOC_106 NAND2X1_LOC_106/a_36_24# NOR2X1_LOC_554/B VSS VDD INVX1_LOC_36/Y
+ NOR2X1_LOC_105/Y NAND2X1_LOC
XNAND2X1_LOC_139 NAND2X1_LOC_139/a_36_24# NAND2X1_LOC_141/A VSS VDD NAND2X1_LOC_139/A
+ INVX1_LOC_80/Y NAND2X1_LOC
XNAND2X1_LOC_128 NAND2X1_LOC_128/a_36_24# NAND2X1_LOC_140/A VSS VDD NOR2X1_LOC_125/Y
+ NOR2X1_LOC_127/Y NAND2X1_LOC
XNOR2X1_LOC_161 NOR2X1_LOC_161/a_36_216# NOR2X1_LOC_161/Y VSS VDD INVX1_LOC_91/A INVX1_LOC_77/A
+ NOR2X1_LOC
XNOR2X1_LOC_194 NOR2X1_LOC_194/a_36_216# NOR2X1_LOC_194/Y VSS VDD NAND2X1_LOC_39/Y
+ NAND2X1_LOC_16/Y NOR2X1_LOC
XNOR2X1_LOC_172 NOR2X1_LOC_172/a_36_216# NOR2X1_LOC_172/Y VSS VDD NOR2X1_LOC_536/A
+ INVX1_LOC_53/Y NOR2X1_LOC
XNOR2X1_LOC_150 NOR2X1_LOC_150/a_36_216# INVX1_LOC_88/A VSS VDD INVX1_LOC_47/Y INVX1_LOC_25/Y
+ NOR2X1_LOC
XNOR2X1_LOC_183 NOR2X1_LOC_183/a_36_216# INVX1_LOC_98/A VSS VDD INVX1_LOC_29/Y INVX1_LOC_6/A
+ NOR2X1_LOC
XNAND2X1_LOC_640 NAND2X1_LOC_640/a_36_24# NAND2X1_LOC_640/Y VSS VDD NAND2X1_LOC_633/Y
+ NAND2X1_LOC_634/Y NAND2X1_LOC
XNAND2X1_LOC_673 NAND2X1_LOC_673/a_36_24# NAND2X1_LOC_721/A VSS VDD NOR2X1_LOC_670/Y
+ NOR2X1_LOC_672/Y NAND2X1_LOC
XNAND2X1_LOC_684 NAND2X1_LOC_684/a_36_24# NOR2X1_LOC_686/A VSS VDD INVX1_LOC_11/A
+ INVX1_LOC_31/A NAND2X1_LOC
XNAND2X1_LOC_662 NAND2X1_LOC_662/a_36_24# NAND2X1_LOC_662/Y VSS VDD NAND2X1_LOC_660/Y
+ NAND2X1_LOC_662/B NAND2X1_LOC
XNAND2X1_LOC_651 NAND2X1_LOC_651/a_36_24# NAND2X1_LOC_654/B VSS VDD NAND2X1_LOC_638/Y
+ NAND2X1_LOC_651/B NAND2X1_LOC
XNAND2X1_LOC_695 NAND2X1_LOC_695/a_36_24# NOR2X1_LOC_707/A VSS VDD NOR2X1_LOC_160/B
+ INVX1_LOC_35/A NAND2X1_LOC
XINVX1_LOC_74 INVX1_LOC_74/Y VSS VDD INVX1_LOC_74/A INVX1_LOC
XINVX1_LOC_30 INVX1_LOC_30/Y VSS VDD INVX1_LOC_30/A INVX1_LOC
XINVX1_LOC_41 INVX1_LOC_41/Y VSS VDD INVX1_LOC_41/A INVX1_LOC
XINVX1_LOC_63 INVX1_LOC_63/Y VSS VDD INVX1_LOC_63/A INVX1_LOC
XINVX1_LOC_96 INVX1_LOC_96/Y VSS VDD INVX1_LOC_96/A INVX1_LOC
XINVX1_LOC_52 INVX1_LOC_52/Y VSS VDD INVX1_LOC_52/A INVX1_LOC
XINVX1_LOC_85 INVX1_LOC_85/Y VSS VDD INVX1_LOC_85/A INVX1_LOC
XNOR2X1_LOC_7 NOR2X1_LOC_7/a_36_216# NOR2X1_LOC_7/Y VSS VDD INVX1_LOC_6/A INVX1_LOC_2/A
+ NOR2X1_LOC
XNAND2X1_LOC_481 NAND2X1_LOC_481/a_36_24# INVX1_LOC_205/A VSS VDD INVX1_LOC_2/Y NOR2X1_LOC_294/Y
+ NAND2X1_LOC
XNAND2X1_LOC_470 NAND2X1_LOC_470/a_36_24# NAND2X1_LOC_477/A VSS VDD NAND2X1_LOC_466/Y
+ NAND2X1_LOC_470/B NAND2X1_LOC
XNAND2X1_LOC_492 NAND2X1_LOC_492/a_36_24# NOR2X1_LOC_493/A VSS VDD INVX1_LOC_45/A
+ INVX1_LOC_75/A NAND2X1_LOC
XINVX1_LOC_303 INVX1_LOC_303/Y VSS VDD INVX1_LOC_303/A INVX1_LOC
XINVX1_LOC_314 INVX1_LOC_314/Y VSS VDD INVX1_LOC_314/A INVX1_LOC
XNOR2X1_LOC_705 NOR2X1_LOC_705/a_36_216# NOR2X1_LOC_713/B VSS VDD NOR2X1_LOC_546/A
+ NOR2X1_LOC_705/B NOR2X1_LOC
XNOR2X1_LOC_727 NOR2X1_LOC_727/a_36_216# NOR2X1_LOC_731/A VSS VDD INVX1_LOC_186/A
+ NOR2X1_LOC_727/B NOR2X1_LOC
XNOR2X1_LOC_738 NOR2X1_LOC_738/a_36_216# NOR2X1_LOC_738/Y VSS VDD NOR2X1_LOC_738/A
+ NOR2X1_LOC_731/Y NOR2X1_LOC
XNOR2X1_LOC_749 NOR2X1_LOC_749/a_36_216# NOR2X1_LOC_749/Y VSS VDD INVX1_LOC_8/A INPUT_0
+ NOR2X1_LOC
XNOR2X1_LOC_716 NOR2X1_LOC_716/a_36_216# INVX1_LOC_282/A VSS VDD INVX1_LOC_140/A NOR2X1_LOC_716/B
+ NOR2X1_LOC
XINVX1_LOC_100 INVX1_LOC_100/Y VSS VDD INVX1_LOC_100/A INVX1_LOC
XINVX1_LOC_122 INVX1_LOC_122/Y VSS VDD INVX1_LOC_122/A INVX1_LOC
XINVX1_LOC_166 INVX1_LOC_166/Y VSS VDD INVX1_LOC_166/A INVX1_LOC
XINVX1_LOC_111 INVX1_LOC_111/Y VSS VDD INVX1_LOC_111/A INVX1_LOC
XINVX1_LOC_155 INVX1_LOC_155/Y VSS VDD INVX1_LOC_155/A INVX1_LOC
XINVX1_LOC_177 INVX1_LOC_177/Y VSS VDD INVX1_LOC_177/A INVX1_LOC
XINVX1_LOC_133 INVX1_LOC_133/Y VSS VDD INVX1_LOC_133/A INVX1_LOC
XINVX1_LOC_188 INVX1_LOC_188/Y VSS VDD INVX1_LOC_188/A INVX1_LOC
XINVX1_LOC_144 INVX1_LOC_144/Y VSS VDD INVX1_LOC_144/A INVX1_LOC
XINVX1_LOC_199 INVX1_LOC_199/Y VSS VDD INVX1_LOC_199/A INVX1_LOC
XNOR2X1_LOC_513 NOR2X1_LOC_513/a_36_216# NOR2X1_LOC_513/Y VSS VDD NOR2X1_LOC_512/Y
+ INVX1_LOC_214/Y NOR2X1_LOC
XNOR2X1_LOC_524 NOR2X1_LOC_524/a_36_216# NOR2X1_LOC_524/Y VSS VDD INVX1_LOC_78/A INVX1_LOC_36/A
+ NOR2X1_LOC
XNOR2X1_LOC_535 NOR2X1_LOC_535/a_36_216# NOR2X1_LOC_567/B VSS VDD INVX1_LOC_222/Y
+ NOR2X1_LOC_788/B NOR2X1_LOC
XNOR2X1_LOC_502 NOR2X1_LOC_502/a_36_216# NOR2X1_LOC_502/Y VSS VDD INVX1_LOC_83/A NOR2X1_LOC_78/A
+ NOR2X1_LOC
XNOR2X1_LOC_546 NOR2X1_LOC_546/a_36_216# NOR2X1_LOC_550/B VSS VDD NOR2X1_LOC_546/A
+ NOR2X1_LOC_546/B NOR2X1_LOC
XNOR2X1_LOC_568 NOR2X1_LOC_568/a_36_216# INVX1_LOC_232/A VSS VDD NOR2X1_LOC_568/A
+ NOR2X1_LOC_566/Y NOR2X1_LOC
XNOR2X1_LOC_579 NOR2X1_LOC_579/a_36_216# INVX1_LOC_242/A VSS VDD INVX1_LOC_237/Y NOR2X1_LOC_575/Y
+ NOR2X1_LOC
XNOR2X1_LOC_557 NOR2X1_LOC_557/a_36_216# NOR2X1_LOC_557/Y VSS VDD NOR2X1_LOC_557/A
+ NOR2X1_LOC_772/B NOR2X1_LOC
XNOR2X1_LOC_376 NOR2X1_LOC_376/a_36_216# NOR2X1_LOC_376/Y VSS VDD NOR2X1_LOC_376/A
+ INVX1_LOC_84/A NOR2X1_LOC
XNOR2X1_LOC_365 NOR2X1_LOC_365/a_36_216# NOR2X1_LOC_367/B VSS VDD NOR2X1_LOC_364/Y
+ INVX1_LOC_159/Y NOR2X1_LOC
XNOR2X1_LOC_321 NOR2X1_LOC_321/a_36_216# NOR2X1_LOC_321/Y VSS VDD INVX1_LOC_50/A INVX1_LOC_9/Y
+ NOR2X1_LOC
XNOR2X1_LOC_354 NOR2X1_LOC_354/a_36_216# NOR2X1_LOC_354/Y VSS VDD NOR2X1_LOC_326/Y
+ NOR2X1_LOC_354/B NOR2X1_LOC
XNOR2X1_LOC_310 NOR2X1_LOC_310/a_36_216# NOR2X1_LOC_310/Y VSS VDD INVX1_LOC_30/A INVX1_LOC_4/A
+ NOR2X1_LOC
XNOR2X1_LOC_343 NOR2X1_LOC_343/a_36_216# NOR2X1_LOC_349/A VSS VDD NOR2X1_LOC_843/B
+ NOR2X1_LOC_343/B NOR2X1_LOC
XNOR2X1_LOC_332 NOR2X1_LOC_332/a_36_216# NOR2X1_LOC_332/Y VSS VDD NOR2X1_LOC_332/A
+ NOR2X1_LOC_332/B NOR2X1_LOC
XNOR2X1_LOC_387 NOR2X1_LOC_387/a_36_216# NOR2X1_LOC_387/Y VSS VDD NOR2X1_LOC_387/A
+ NOR2X1_LOC_92/Y NOR2X1_LOC
XNOR2X1_LOC_398 NOR2X1_LOC_398/a_36_216# NOR2X1_LOC_398/Y VSS VDD INVX1_LOC_135/A
+ NOR2X1_LOC_78/B NOR2X1_LOC
XNAND2X1_LOC_822 NAND2X1_LOC_822/a_36_24# NOR2X1_LOC_835/A VSS VDD INVX1_LOC_49/A
+ NOR2X1_LOC_590/A NAND2X1_LOC
XNAND2X1_LOC_811 NAND2X1_LOC_811/a_36_24# NAND2X1_LOC_811/Y VSS VDD NAND2X1_LOC_807/Y
+ NAND2X1_LOC_811/B NAND2X1_LOC
XNAND2X1_LOC_800 NAND2X1_LOC_800/a_36_24# NAND2X1_LOC_800/Y VSS VDD NAND2X1_LOC_800/A
+ INVX1_LOC_291/Y NAND2X1_LOC
XNAND2X1_LOC_833 NAND2X1_LOC_833/a_36_24# NAND2X1_LOC_833/Y VSS VDD NOR2X1_LOC_482/Y
+ NOR2X1_LOC_495/Y NAND2X1_LOC
XNAND2X1_LOC_866 NAND2X1_LOC_866/a_36_24# GATE_865 VSS VDD NAND2X1_LOC_866/A NAND2X1_LOC_866/B
+ NAND2X1_LOC
XNAND2X1_LOC_844 NAND2X1_LOC_844/a_36_24# NAND2X1_LOC_849/A VSS VDD NOR2X1_LOC_497/Y
+ NAND2X1_LOC_560/A NAND2X1_LOC
XNAND2X1_LOC_855 NAND2X1_LOC_855/a_36_24# NAND2X1_LOC_855/Y VSS VDD NAND2X1_LOC_729/B
+ NOR2X1_LOC_829/Y NAND2X1_LOC
XNOR2X1_LOC_50 NOR2X1_LOC_50/a_36_216# NOR2X1_LOC_51/A VSS VDD INPUT_7 INPUT_6
+ NOR2X1_LOC
XNOR2X1_LOC_61 NOR2X1_LOC_61/a_36_216# NOR2X1_LOC_61/Y VSS VDD NOR2X1_LOC_61/A NOR2X1_LOC_61/B
+ NOR2X1_LOC
XNOR2X1_LOC_94 NOR2X1_LOC_94/a_36_216# NOR2X1_LOC_94/Y VSS VDD INVX1_LOC_39/A INVX1_LOC_14/A
+ NOR2X1_LOC
XNOR2X1_LOC_72 NOR2X1_LOC_72/a_36_216# NOR2X1_LOC_72/Y VSS VDD NOR2X1_LOC_71/Y INVX1_LOC_53/Y
+ NOR2X1_LOC
XNOR2X1_LOC_83 NOR2X1_LOC_83/a_36_216# NOR2X1_LOC_83/Y VSS VDD NOR2X1_LOC_82/Y INVX1_LOC_20/A
+ NOR2X1_LOC
XNAND2X1_LOC_107 NAND2X1_LOC_107/a_36_24# NOR2X1_LOC_113/A VSS VDD INVX1_LOC_49/A
+ NOR2X1_LOC_78/A NAND2X1_LOC
XNAND2X1_LOC_129 NAND2X1_LOC_129/a_36_24# NOR2X1_LOC_130/A VSS VDD NOR2X1_LOC_38/B
+ INVX1_LOC_25/A NAND2X1_LOC
XNAND2X1_LOC_5 NAND2X1_LOC_5/a_36_24# INVX1_LOC_3/A VSS VDD D_INPUT_2 INPUT_3
+ NAND2X1_LOC
XNAND2X1_LOC_118 NAND2X1_LOC_118/a_36_24# INVX1_LOC_69/A VSS VDD INVX1_LOC_53/A NOR2X1_LOC_78/A
+ NAND2X1_LOC
XNOR2X1_LOC_162 NOR2X1_LOC_162/a_36_216# NOR2X1_LOC_162/Y VSS VDD NOR2X1_LOC_161/Y
+ NOR2X1_LOC_160/Y NOR2X1_LOC
XNOR2X1_LOC_151 NOR2X1_LOC_151/a_36_216# NOR2X1_LOC_151/Y VSS VDD INVX1_LOC_88/Y INVX1_LOC_42/Y
+ NOR2X1_LOC
XNOR2X1_LOC_173 NOR2X1_LOC_173/a_36_216# NOR2X1_LOC_173/Y VSS VDD INVX1_LOC_88/A INVX1_LOC_54/A
+ NOR2X1_LOC
XNOR2X1_LOC_140 NOR2X1_LOC_140/a_36_216# INVX1_LOC_82/A VSS VDD NOR2X1_LOC_140/A NOR2X1_LOC_554/A
+ NOR2X1_LOC
XNOR2X1_LOC_195 NOR2X1_LOC_195/a_36_216# NOR2X1_LOC_199/B VSS VDD NOR2X1_LOC_195/A
+ NAND2X1_LOC_41/Y NOR2X1_LOC
XNOR2X1_LOC_184 NOR2X1_LOC_184/a_36_216# INVX1_LOC_100/A VSS VDD INVX1_LOC_58/A NOR2X1_LOC_71/Y
+ NOR2X1_LOC
XNAND2X1_LOC_641 NAND2X1_LOC_641/a_36_24# NAND2X1_LOC_650/B VSS VDD NAND2X1_LOC_231/Y
+ INVX1_LOC_126/A NAND2X1_LOC
XNAND2X1_LOC_652 NAND2X1_LOC_652/a_36_24# NAND2X1_LOC_652/Y VSS VDD NAND2X1_LOC_468/B
+ NAND2X1_LOC_593/Y NAND2X1_LOC
XNAND2X1_LOC_630 NAND2X1_LOC_630/a_36_24# INVX1_LOC_259/A VSS VDD INVX1_LOC_257/Y
+ NAND2X1_LOC_629/Y NAND2X1_LOC
XNAND2X1_LOC_663 NAND2X1_LOC_663/a_36_24# GATE_662 VSS VDD INVX1_LOC_268/Y NAND2X1_LOC_662/Y
+ NAND2X1_LOC
XINVX1_LOC_20 INVX1_LOC_20/Y VSS VDD INVX1_LOC_20/A INVX1_LOC
XINVX1_LOC_31 INVX1_LOC_31/Y VSS VDD INVX1_LOC_31/A INVX1_LOC
XINVX1_LOC_42 INVX1_LOC_42/Y VSS VDD INVX1_LOC_42/A INVX1_LOC
XNAND2X1_LOC_674 NAND2X1_LOC_674/a_36_24# NOR2X1_LOC_675/A VSS VDD INVX1_LOC_53/A
+ NOR2X1_LOC_405/A NAND2X1_LOC
XNAND2X1_LOC_685 NAND2X1_LOC_685/a_36_24# NAND2X1_LOC_687/A VSS VDD NOR2X1_LOC_681/Y
+ NOR2X1_LOC_682/Y NAND2X1_LOC
XNAND2X1_LOC_696 NAND2X1_LOC_696/a_36_24# NOR2X1_LOC_708/B VSS VDD INVX1_LOC_19/A
+ INVX1_LOC_83/A NAND2X1_LOC
XINVX1_LOC_64 INVX1_LOC_64/Y VSS VDD INVX1_LOC_64/A INVX1_LOC
XINVX1_LOC_53 INVX1_LOC_53/Y VSS VDD INVX1_LOC_53/A INVX1_LOC
XINVX1_LOC_97 INVX1_LOC_97/Y VSS VDD INVX1_LOC_97/A INVX1_LOC
XINVX1_LOC_86 INVX1_LOC_86/Y VSS VDD INVX1_LOC_86/A INVX1_LOC
XINVX1_LOC_75 INVX1_LOC_75/Y VSS VDD INVX1_LOC_75/A INVX1_LOC
XNOR2X1_LOC_8 NOR2X1_LOC_8/a_36_216# INVX1_LOC_8/A VSS VDD INPUT_3 D_INPUT_2 NOR2X1_LOC
XNAND2X1_LOC_471 NAND2X1_LOC_471/a_36_24# NAND2X1_LOC_471/Y VSS VDD NAND2X1_LOC_464/Y
+ NAND2X1_LOC_465/Y NAND2X1_LOC
XNAND2X1_LOC_493 NAND2X1_LOC_493/a_36_24# NAND2X1_LOC_493/Y VSS VDD NOR2X1_LOC_491/Y
+ NOR2X1_LOC_492/Y NAND2X1_LOC
XNAND2X1_LOC_482 NAND2X1_LOC_482/a_36_24# NOR2X1_LOC_833/B VSS VDD INVX1_LOC_5/A INVX1_LOC_45/A
+ NAND2X1_LOC
XNAND2X1_LOC_460 NAND2X1_LOC_460/a_36_24# NAND2X1_LOC_463/B VSS VDD NOR2X1_LOC_380/Y
+ NOR2X1_LOC_409/Y NAND2X1_LOC
XINVX1_LOC_315 INVX1_LOC_315/Y VSS VDD INVX1_LOC_315/A INVX1_LOC
XINVX1_LOC_304 INVX1_LOC_304/Y VSS VDD INVX1_LOC_304/A INVX1_LOC
XNOR2X1_LOC_706 NOR2X1_LOC_706/a_36_216# NOR2X1_LOC_706/Y VSS VDD NOR2X1_LOC_706/A
+ NOR2X1_LOC_706/B NOR2X1_LOC
XNOR2X1_LOC_717 NOR2X1_LOC_717/a_36_216# NOR2X1_LOC_717/Y VSS VDD NOR2X1_LOC_717/A
+ NOR2X1_LOC_717/B NOR2X1_LOC
XNAND2X1_LOC_290 NAND2X1_LOC_290/a_36_24# NOR2X1_LOC_634/B VSS VDD NOR2X1_LOC_78/B
+ INVX1_LOC_19/A NAND2X1_LOC
XNOR2X1_LOC_739 NOR2X1_LOC_739/a_36_216# NOR2X1_LOC_739/Y VSS VDD NOR2X1_LOC_730/Y
+ INVX1_LOC_104/A NOR2X1_LOC
XNOR2X1_LOC_728 NOR2X1_LOC_728/a_36_216# NOR2X1_LOC_730/B VSS VDD INVX1_LOC_274/Y
+ NOR2X1_LOC_728/B NOR2X1_LOC
XINVX1_LOC_112 INVX1_LOC_112/Y VSS VDD INVX1_LOC_112/A INVX1_LOC
XINVX1_LOC_123 INVX1_LOC_123/Y VSS VDD INVX1_LOC_123/A INVX1_LOC
XINVX1_LOC_134 INVX1_LOC_134/Y VSS VDD INVX1_LOC_134/A INVX1_LOC
XINVX1_LOC_101 INVX1_LOC_101/Y VSS VDD INVX1_LOC_101/A INVX1_LOC
XINVX1_LOC_156 INVX1_LOC_156/Y VSS VDD INVX1_LOC_156/A INVX1_LOC
XINVX1_LOC_167 INVX1_LOC_167/Y VSS VDD INVX1_LOC_167/A INVX1_LOC
XINVX1_LOC_178 INVX1_LOC_178/Y VSS VDD INVX1_LOC_178/A INVX1_LOC
XINVX1_LOC_145 INVX1_LOC_145/Y VSS VDD INVX1_LOC_145/A INVX1_LOC
XINVX1_LOC_189 INVX1_LOC_189/Y VSS VDD INVX1_LOC_189/A INVX1_LOC
XNOR2X1_LOC_503 NOR2X1_LOC_503/a_36_216# NOR2X1_LOC_503/Y VSS VDD NOR2X1_LOC_503/A
+ INVX1_LOC_49/Y NOR2X1_LOC
XNOR2X1_LOC_536 NOR2X1_LOC_536/a_36_216# NOR2X1_LOC_536/Y VSS VDD NOR2X1_LOC_536/A
+ INVX1_LOC_12/A NOR2X1_LOC
XNOR2X1_LOC_558 NOR2X1_LOC_558/a_36_216# NOR2X1_LOC_561/A VSS VDD NOR2X1_LOC_558/A
+ NOR2X1_LOC_717/A NOR2X1_LOC
XNOR2X1_LOC_514 NOR2X1_LOC_514/a_36_216# NOR2X1_LOC_514/Y VSS VDD NOR2X1_LOC_514/A
+ INPUT_0 NOR2X1_LOC
XNOR2X1_LOC_547 NOR2X1_LOC_547/a_36_216# INVX1_LOC_226/A VSS VDD NOR2X1_LOC_620/B
+ NOR2X1_LOC_547/B NOR2X1_LOC
XNOR2X1_LOC_525 NOR2X1_LOC_525/a_36_216# NOR2X1_LOC_525/Y VSS VDD INVX1_LOC_38/A INVX1_LOC_10/A
+ NOR2X1_LOC
XNOR2X1_LOC_569 NOR2X1_LOC_569/a_36_216# NOR2X1_LOC_569/Y VSS VDD NOR2X1_LOC_569/A
+ NOR2X1_LOC_564/Y NOR2X1_LOC
XNOR2X1_LOC_377 NOR2X1_LOC_377/a_36_216# NOR2X1_LOC_377/Y VSS VDD INVX1_LOC_14/Y INVX1_LOC_2/A
+ NOR2X1_LOC
XNOR2X1_LOC_300 NOR2X1_LOC_300/a_36_216# NOR2X1_LOC_300/Y VSS VDD INVX1_LOC_72/A INVX1_LOC_46/A
+ NOR2X1_LOC
XNOR2X1_LOC_366 NOR2X1_LOC_366/a_36_216# NOR2X1_LOC_366/Y VSS VDD NOR2X1_LOC_363/Y
+ NOR2X1_LOC_366/B NOR2X1_LOC
XNOR2X1_LOC_344 NOR2X1_LOC_344/a_36_216# NOR2X1_LOC_348/B VSS VDD NOR2X1_LOC_344/A
+ NOR2X1_LOC_254/Y NOR2X1_LOC
XNOR2X1_LOC_388 NOR2X1_LOC_388/a_36_216# NOR2X1_LOC_388/Y VSS VDD NOR2X1_LOC_180/B
+ NOR2X1_LOC_703/B NOR2X1_LOC
XNOR2X1_LOC_355 NOR2X1_LOC_355/a_36_216# NOR2X1_LOC_356/A VSS VDD NOR2X1_LOC_355/A
+ NOR2X1_LOC_355/B NOR2X1_LOC
XNOR2X1_LOC_311 NOR2X1_LOC_311/a_36_216# NOR2X1_LOC_311/Y VSS VDD NOR2X1_LOC_536/A
+ INVX1_LOC_20/A NOR2X1_LOC
XNOR2X1_LOC_322 NOR2X1_LOC_322/a_36_216# NOR2X1_LOC_322/Y VSS VDD INVX1_LOC_84/A INVX1_LOC_33/Y
+ NOR2X1_LOC
XNOR2X1_LOC_399 NOR2X1_LOC_399/a_36_216# NOR2X1_LOC_399/Y VSS VDD NOR2X1_LOC_399/A
+ INVX1_LOC_34/A NOR2X1_LOC
XNOR2X1_LOC_333 NOR2X1_LOC_333/a_36_216# INVX1_LOC_148/A VSS VDD NOR2X1_LOC_333/A
+ NOR2X1_LOC_174/B NOR2X1_LOC
XNAND2X1_LOC_823 NAND2X1_LOC_823/a_36_24# NOR2X1_LOC_836/B VSS VDD INVX1_LOC_37/A
+ INVX1_LOC_117/A NAND2X1_LOC
XNAND2X1_LOC_845 NAND2X1_LOC_845/a_36_24# NAND2X1_LOC_849/B VSS VDD NAND2X1_LOC_721/A
+ NOR2X1_LOC_813/Y NAND2X1_LOC
XNAND2X1_LOC_812 NAND2X1_LOC_812/a_36_24# GATE_811 VSS VDD NAND2X1_LOC_812/A NAND2X1_LOC_811/Y
+ NAND2X1_LOC
XNAND2X1_LOC_834 NAND2X1_LOC_834/a_36_24# NAND2X1_LOC_840/B VSS VDD INVX1_LOC_214/A
+ NOR2X1_LOC_677/Y NAND2X1_LOC
XNAND2X1_LOC_801 NAND2X1_LOC_801/a_36_24# NAND2X1_LOC_809/A VSS VDD NOR2X1_LOC_761/Y
+ NAND2X1_LOC_800/Y NAND2X1_LOC
XNAND2X1_LOC_856 NAND2X1_LOC_856/a_36_24# NAND2X1_LOC_863/A VSS VDD NAND2X1_LOC_856/A
+ NAND2X1_LOC_855/Y NAND2X1_LOC
XNOR2X1_LOC_51 NOR2X1_LOC_51/a_36_216# INVX1_LOC_38/A VSS VDD NOR2X1_LOC_51/A NOR2X1_LOC_30/Y
+ NOR2X1_LOC
XNOR2X1_LOC_40 NOR2X1_LOC_40/a_36_216# INVX1_LOC_30/A VSS VDD NOR2X1_LOC_25/Y NOR2X1_LOC_2/Y
+ NOR2X1_LOC
XNOR2X1_LOC_95 NOR2X1_LOC_95/a_36_216# INVX1_LOC_58/A VSS VDD NOR2X1_LOC_51/A NOR2X1_LOC_11/Y
+ NOR2X1_LOC
XNOR2X1_LOC_84 NOR2X1_LOC_84/a_36_216# NOR2X1_LOC_84/Y VSS VDD NOR2X1_LOC_84/A NOR2X1_LOC_84/B
+ NOR2X1_LOC
XNOR2X1_LOC_62 NOR2X1_LOC_62/a_36_216# INVX1_LOC_48/A VSS VDD INVX1_LOC_39/A NAND2X1_LOC_9/Y
+ NOR2X1_LOC
XNOR2X1_LOC_73 NOR2X1_LOC_73/a_36_216# NOR2X1_LOC_74/A VSS VDD INVX1_LOC_26/A NOR2X1_LOC_9/Y
+ NOR2X1_LOC
XNAND2X1_LOC_108 NAND2X1_LOC_108/a_36_24# INVX1_LOC_65/A VSS VDD INVX1_LOC_45/A NOR2X1_LOC_590/A
+ NAND2X1_LOC
XNAND2X1_LOC_119 NAND2X1_LOC_119/a_36_24# INVX1_LOC_71/A VSS VDD INPUT_1 INVX1_LOC_13/A
+ NAND2X1_LOC
XNAND2X1_LOC_6 NAND2X1_LOC_6/a_36_24# INVX1_LOC_5/A VSS VDD NOR2X1_LOC_19/B INVX1_LOC_3/A
+ NAND2X1_LOC
XNOR2X1_LOC_163 NOR2X1_LOC_163/a_36_216# NOR2X1_LOC_163/Y VSS VDD NOR2X1_LOC_163/A
+ INVX1_LOC_38/A NOR2X1_LOC
XNOR2X1_LOC_141 NOR2X1_LOC_141/a_36_216# NOR2X1_LOC_657/B VSS VDD INVX1_LOC_81/Y NOR2X1_LOC_139/Y
+ NOR2X1_LOC
XNOR2X1_LOC_152 NOR2X1_LOC_152/a_36_216# NOR2X1_LOC_152/Y VSS VDD NOR2X1_LOC_152/A
+ INVX1_LOC_36/A NOR2X1_LOC
XNOR2X1_LOC_174 NOR2X1_LOC_174/a_36_216# NOR2X1_LOC_175/A VSS VDD NOR2X1_LOC_174/A
+ NOR2X1_LOC_174/B NOR2X1_LOC
XNOR2X1_LOC_196 NOR2X1_LOC_196/a_36_216# NOR2X1_LOC_196/Y VSS VDD NOR2X1_LOC_196/A
+ NAND2X1_LOC_45/Y NOR2X1_LOC
XNOR2X1_LOC_130 NOR2X1_LOC_130/a_36_216# NOR2X1_LOC_130/Y VSS VDD NOR2X1_LOC_130/A
+ INVX1_LOC_5/A NOR2X1_LOC
XNOR2X1_LOC_185 NOR2X1_LOC_185/a_36_216# NOR2X1_LOC_188/A VSS VDD NAND2X1_LOC_74/B
+ INVX1_LOC_41/A NOR2X1_LOC
XNAND2X1_LOC_620 NAND2X1_LOC_620/a_36_24# NAND2X1_LOC_623/B VSS VDD NOR2X1_LOC_528/Y
+ NOR2X1_LOC_613/Y NAND2X1_LOC
XNAND2X1_LOC_642 NAND2X1_LOC_642/a_36_24# NAND2X1_LOC_642/Y VSS VDD INVX1_LOC_176/A
+ INVX1_LOC_218/Y NAND2X1_LOC
XNAND2X1_LOC_631 NAND2X1_LOC_631/a_36_24# NAND2X1_LOC_632/B VSS VDD NAND2X1_LOC_483/Y
+ NOR2X1_LOC_625/Y NAND2X1_LOC
XNAND2X1_LOC_675 NAND2X1_LOC_675/a_36_24# INVX1_LOC_269/A VSS VDD INVX1_LOC_182/Y
+ NOR2X1_LOC_674/Y NAND2X1_LOC
XNAND2X1_LOC_664 NAND2X1_LOC_664/a_36_24# NOR2X1_LOC_665/A VSS VDD NOR2X1_LOC_74/A
+ NOR2X1_LOC_89/A NAND2X1_LOC
XNAND2X1_LOC_653 NAND2X1_LOC_653/a_36_24# NAND2X1_LOC_661/A VSS VDD NOR2X1_LOC_594/Y
+ NAND2X1_LOC_652/Y NAND2X1_LOC
XNAND2X1_LOC_697 NAND2X1_LOC_697/a_36_24# NOR2X1_LOC_708/A VSS VDD INVX1_LOC_89/A
+ INVX1_LOC_117/A NAND2X1_LOC
XNAND2X1_LOC_686 NAND2X1_LOC_686/a_36_24# INVX1_LOC_275/A VSS VDD NOR2X1_LOC_683/Y
+ NOR2X1_LOC_684/Y NAND2X1_LOC
XINVX1_LOC_43 INVX1_LOC_43/Y VSS VDD INVX1_LOC_43/A INVX1_LOC
XINVX1_LOC_65 INVX1_LOC_65/Y VSS VDD INVX1_LOC_65/A INVX1_LOC
XINVX1_LOC_54 INVX1_LOC_54/Y VSS VDD INVX1_LOC_54/A INVX1_LOC
XINVX1_LOC_21 INVX1_LOC_21/Y VSS VDD INVX1_LOC_21/A INVX1_LOC
XINVX1_LOC_10 INVX1_LOC_10/Y VSS VDD INVX1_LOC_10/A INVX1_LOC
XINVX1_LOC_76 INVX1_LOC_76/Y VSS VDD INVX1_LOC_76/A INVX1_LOC
XINVX1_LOC_32 INVX1_LOC_32/Y VSS VDD INVX1_LOC_32/A INVX1_LOC
XINVX1_LOC_87 INVX1_LOC_87/Y VSS VDD INVX1_LOC_87/A INVX1_LOC
XINVX1_LOC_98 INVX1_LOC_98/Y VSS VDD INVX1_LOC_98/A INVX1_LOC
XNOR2X1_LOC_9 NOR2X1_LOC_9/a_36_216# NOR2X1_LOC_9/Y VSS VDD INPUT_1 INPUT_0 NOR2X1_LOC
XNAND2X1_LOC_494 NAND2X1_LOC_494/a_36_24# NOR2X1_LOC_558/A VSS VDD INVX1_LOC_12/Y
+ NOR2X1_LOC_383/Y NAND2X1_LOC
XNAND2X1_LOC_483 NAND2X1_LOC_483/a_36_24# NAND2X1_LOC_483/Y VSS VDD NOR2X1_LOC_252/Y
+ NOR2X1_LOC_482/Y NAND2X1_LOC
XNAND2X1_LOC_461 NAND2X1_LOC_461/a_36_24# NAND2X1_LOC_462/B VSS VDD NOR2X1_LOC_411/Y
+ NOR2X1_LOC_413/Y NAND2X1_LOC
XNAND2X1_LOC_472 NAND2X1_LOC_472/a_36_24# NAND2X1_LOC_472/Y VSS VDD INVX1_LOC_196/Y
+ INVX1_LOC_198/Y NAND2X1_LOC
XNAND2X1_LOC_450 NAND2X1_LOC_450/a_36_24# INVX1_LOC_191/A VSS VDD NOR2X1_LOC_426/Y
+ NOR2X1_LOC_427/Y NAND2X1_LOC
XINVX1_LOC_316 INVX1_LOC_316/Y VSS VDD INVX1_LOC_316/A INVX1_LOC
XINVX1_LOC_305 INVX1_LOC_305/Y VSS VDD INVX1_LOC_305/A INVX1_LOC
XNOR2X1_LOC_707 NOR2X1_LOC_707/a_36_216# NOR2X1_LOC_712/B VSS VDD NOR2X1_LOC_707/A
+ NOR2X1_LOC_707/B NOR2X1_LOC
XNOR2X1_LOC_718 NOR2X1_LOC_718/a_36_216# NOR2X1_LOC_718/Y VSS VDD INVX1_LOC_249/Y
+ NOR2X1_LOC_718/B NOR2X1_LOC
XNOR2X1_LOC_729 NOR2X1_LOC_729/a_36_216# NOR2X1_LOC_730/A VSS VDD NOR2X1_LOC_729/A
+ NOR2X1_LOC_687/Y NOR2X1_LOC
XNAND2X1_LOC_291 NAND2X1_LOC_291/a_36_24# NOR2X1_LOC_334/A VSS VDD INVX1_LOC_23/A
+ NAND2X1_LOC_291/B NAND2X1_LOC
XNAND2X1_LOC_280 NAND2X1_LOC_280/a_36_24# NOR2X1_LOC_542/B VSS VDD INVX1_LOC_35/A
+ INVX1_LOC_117/A NAND2X1_LOC
XINVX1_LOC_135 INVX1_LOC_135/Y VSS VDD INVX1_LOC_135/A INVX1_LOC
XINVX1_LOC_168 INVX1_LOC_168/Y VSS VDD INVX1_LOC_168/A INVX1_LOC
XINVX1_LOC_124 INVX1_LOC_124/Y VSS VDD INVX1_LOC_124/A INVX1_LOC
XINVX1_LOC_102 INVX1_LOC_102/Y VSS VDD INVX1_LOC_102/A INVX1_LOC
XINVX1_LOC_157 INVX1_LOC_157/Y VSS VDD INVX1_LOC_157/A INVX1_LOC
XINVX1_LOC_146 INVX1_LOC_146/Y VSS VDD INVX1_LOC_146/A INVX1_LOC
XINVX1_LOC_113 INVX1_LOC_113/Y VSS VDD INVX1_LOC_113/A INVX1_LOC
XINVX1_LOC_179 INVX1_LOC_179/Y VSS VDD INVX1_LOC_179/A INVX1_LOC
XNOR2X1_LOC_504 NOR2X1_LOC_504/a_36_216# NOR2X1_LOC_504/Y VSS VDD INVX1_LOC_90/A INVX1_LOC_10/A
+ NOR2X1_LOC
XNOR2X1_LOC_548 NOR2X1_LOC_548/a_36_216# NOR2X1_LOC_548/Y VSS VDD NOR2X1_LOC_548/A
+ NOR2X1_LOC_548/B NOR2X1_LOC
XNOR2X1_LOC_537 NOR2X1_LOC_537/a_36_216# NOR2X1_LOC_537/Y VSS VDD NOR2X1_LOC_537/A
+ NOR2X1_LOC_389/B NOR2X1_LOC
XNOR2X1_LOC_515 NOR2X1_LOC_515/a_36_216# INVX1_LOC_216/A VSS VDD NOR2X1_LOC_514/Y
+ INVX1_LOC_178/Y NOR2X1_LOC
XNOR2X1_LOC_559 NOR2X1_LOC_559/a_36_216# NOR2X1_LOC_560/A VSS VDD INVX1_LOC_218/A
+ NOR2X1_LOC_559/B NOR2X1_LOC
XNOR2X1_LOC_526 NOR2X1_LOC_526/a_36_216# NOR2X1_LOC_526/Y VSS VDD INVX1_LOC_91/Y INVX1_LOC_22/A
+ NOR2X1_LOC
XNOR2X1_LOC_301 NOR2X1_LOC_301/a_36_216# INVX1_LOC_140/A VSS VDD NOR2X1_LOC_301/A
+ NOR2X1_LOC_76/A NOR2X1_LOC
XNOR2X1_LOC_378 NOR2X1_LOC_378/a_36_216# NOR2X1_LOC_378/Y VSS VDD NOR2X1_LOC_377/Y
+ INVX1_LOC_32/Y NOR2X1_LOC
XNOR2X1_LOC_367 NOR2X1_LOC_367/a_36_216# D_GATE_366 VSS VDD NOR2X1_LOC_366/Y NOR2X1_LOC_367/B
+ NOR2X1_LOC
XNOR2X1_LOC_356 NOR2X1_LOC_356/a_36_216# INVX1_LOC_160/A VSS VDD NOR2X1_LOC_356/A
+ NOR2X1_LOC_354/Y NOR2X1_LOC
XNOR2X1_LOC_323 NOR2X1_LOC_323/a_36_216# NOR2X1_LOC_323/Y VSS VDD NOR2X1_LOC_111/A
+ INVX1_LOC_57/Y NOR2X1_LOC
XNOR2X1_LOC_312 NOR2X1_LOC_312/a_36_216# NOR2X1_LOC_312/Y VSS VDD INVX1_LOC_50/A INVX1_LOC_42/A
+ NOR2X1_LOC
XNOR2X1_LOC_389 NOR2X1_LOC_389/a_36_216# INVX1_LOC_162/A VSS VDD NOR2X1_LOC_389/A
+ NOR2X1_LOC_389/B NOR2X1_LOC
XNOR2X1_LOC_334 NOR2X1_LOC_334/a_36_216# NOR2X1_LOC_334/Y VSS VDD NOR2X1_LOC_334/A
+ NOR2X1_LOC_634/B NOR2X1_LOC
XNOR2X1_LOC_345 NOR2X1_LOC_345/a_36_216# INVX1_LOC_154/A VSS VDD NOR2X1_LOC_345/A
+ INVX1_LOC_122/A NOR2X1_LOC
XNAND2X1_LOC_835 NAND2X1_LOC_835/a_36_24# NAND2X1_LOC_839/A VSS VDD NOR2X1_LOC_821/Y
+ NOR2X1_LOC_822/Y NAND2X1_LOC
XNAND2X1_LOC_824 NAND2X1_LOC_824/a_36_24# NOR2X1_LOC_836/A VSS VDD INVX1_LOC_19/A
+ NAND2X1_LOC_291/B NAND2X1_LOC
XNAND2X1_LOC_813 NAND2X1_LOC_813/a_36_24# NOR2X1_LOC_845/A VSS VDD INVX1_LOC_48/A
+ INVX1_LOC_123/A NAND2X1_LOC
XNAND2X1_LOC_846 NAND2X1_LOC_846/a_36_24# NAND2X1_LOC_848/A VSS VDD NOR2X1_LOC_815/Y
+ NOR2X1_LOC_816/Y NAND2X1_LOC
XNAND2X1_LOC_802 NAND2X1_LOC_802/a_36_24# NAND2X1_LOC_802/Y VSS VDD NAND2X1_LOC_802/A
+ NAND2X1_LOC_799/Y NAND2X1_LOC
XNAND2X1_LOC_857 NAND2X1_LOC_857/a_36_24# NAND2X1_LOC_863/B VSS VDD NAND2X1_LOC_852/Y
+ NAND2X1_LOC_853/Y NAND2X1_LOC
XNOR2X1_LOC_30 NOR2X1_LOC_30/a_36_216# NOR2X1_LOC_30/Y VSS VDD D_INPUT_5 D_INPUT_4
+ NOR2X1_LOC
XNOR2X1_LOC_74 NOR2X1_LOC_74/a_36_216# NOR2X1_LOC_74/Y VSS VDD NOR2X1_LOC_74/A INVX1_LOC_22/A
+ NOR2X1_LOC
XNOR2X1_LOC_41 NOR2X1_LOC_41/a_36_216# NOR2X1_LOC_41/Y VSS VDD INVX1_LOC_30/A INVX1_LOC_10/A
+ NOR2X1_LOC
XNOR2X1_LOC_52 NOR2X1_LOC_52/a_36_216# NOR2X1_LOC_52/Y VSS VDD INVX1_LOC_38/A NOR2X1_LOC_52/B
+ NOR2X1_LOC
XNOR2X1_LOC_96 NOR2X1_LOC_96/a_36_216# NOR2X1_LOC_96/Y VSS VDD INVX1_LOC_58/A NOR2X1_LOC_94/Y
+ NOR2X1_LOC
XNOR2X1_LOC_63 NOR2X1_LOC_63/a_36_216# NOR2X1_LOC_65/B VSS VDD INVX1_LOC_48/A INVX1_LOC_7/Y
+ NOR2X1_LOC
XNOR2X1_LOC_85 NOR2X1_LOC_85/a_36_216# NOR2X1_LOC_86/A VSS VDD INVX1_LOC_25/Y INVX1_LOC_16/A
+ NOR2X1_LOC
XNAND2X1_LOC_7 NAND2X1_LOC_7/a_36_24# NAND2X1_LOC_7/Y VSS VDD INVX1_LOC_1/A INVX1_LOC_5/A
+ NAND2X1_LOC
XNAND2X1_LOC_109 NAND2X1_LOC_109/a_36_24# NOR2X1_LOC_112/B VSS VDD INVX1_LOC_21/A
+ NOR2X1_LOC_78/A NAND2X1_LOC
XNOR2X1_LOC_142 NOR2X1_LOC_142/a_36_216# NOR2X1_LOC_142/Y VSS VDD INVX1_LOC_50/A NOR2X1_LOC_52/B
+ NOR2X1_LOC
XNOR2X1_LOC_131 NOR2X1_LOC_131/a_36_216# NOR2X1_LOC_131/Y VSS VDD NOR2X1_LOC_131/A
+ INVX1_LOC_12/A NOR2X1_LOC
XNOR2X1_LOC_120 NOR2X1_LOC_120/a_36_216# NOR2X1_LOC_121/A VSS VDD INVX1_LOC_27/A INVX1_LOC_9/A
+ NOR2X1_LOC
XNOR2X1_LOC_197 NOR2X1_LOC_197/a_36_216# NOR2X1_LOC_197/Y VSS VDD NOR2X1_LOC_197/A
+ NOR2X1_LOC_197/B NOR2X1_LOC
XNOR2X1_LOC_186 NOR2X1_LOC_186/a_36_216# NOR2X1_LOC_186/Y VSS VDD NOR2X1_LOC_188/A
+ INVX1_LOC_87/A NOR2X1_LOC
XNOR2X1_LOC_175 NOR2X1_LOC_175/a_36_216# NOR2X1_LOC_211/A VSS VDD NOR2X1_LOC_175/A
+ NOR2X1_LOC_175/B NOR2X1_LOC
XNOR2X1_LOC_153 NOR2X1_LOC_153/a_36_216# NOR2X1_LOC_433/A VSS VDD INVX1_LOC_26/A INPUT_1
+ NOR2X1_LOC
XNOR2X1_LOC_164 NOR2X1_LOC_164/a_36_216# NOR2X1_LOC_164/Y VSS VDD INVX1_LOC_84/A INVX1_LOC_16/A
+ NOR2X1_LOC
XNAND2X1_LOC_698 NAND2X1_LOC_698/a_36_24# NOR2X1_LOC_709/B VSS VDD INVX1_LOC_49/A
+ INVX1_LOC_75/A NAND2X1_LOC
XNAND2X1_LOC_610 NAND2X1_LOC_610/a_36_24# NOR2X1_LOC_612/B VSS VDD INVX1_LOC_30/A
+ INVX1_LOC_36/A NAND2X1_LOC
XNAND2X1_LOC_632 NAND2X1_LOC_632/a_36_24# NAND2X1_LOC_735/B VSS VDD INVX1_LOC_260/Y
+ NAND2X1_LOC_632/B NAND2X1_LOC
XNAND2X1_LOC_665 NAND2X1_LOC_665/a_36_24# NOR2X1_LOC_719/B VSS VDD INVX1_LOC_2/Y NOR2X1_LOC_664/Y
+ NAND2X1_LOC
XNAND2X1_LOC_621 NAND2X1_LOC_621/a_36_24# NAND2X1_LOC_622/B VSS VDD NOR2X1_LOC_616/Y
+ NOR2X1_LOC_617/Y NAND2X1_LOC
XNAND2X1_LOC_643 NAND2X1_LOC_643/a_36_24# NAND2X1_LOC_649/B VSS VDD NAND2X1_LOC_537/Y
+ NOR2X1_LOC_595/Y NAND2X1_LOC
XNAND2X1_LOC_687 NAND2X1_LOC_687/a_36_24# NAND2X1_LOC_800/A VSS VDD NAND2X1_LOC_687/A
+ INVX1_LOC_276/Y NAND2X1_LOC
XNAND2X1_LOC_676 NAND2X1_LOC_676/a_36_24# NOR2X1_LOC_679/B VSS VDD INVX1_LOC_78/A
+ NOR2X1_LOC_599/A NAND2X1_LOC
XNAND2X1_LOC_654 NAND2X1_LOC_654/a_36_24# NAND2X1_LOC_661/B VSS VDD INVX1_LOC_266/Y
+ NAND2X1_LOC_654/B NAND2X1_LOC
XINVX1_LOC_22 INVX1_LOC_22/Y VSS VDD INVX1_LOC_22/A INVX1_LOC
XINVX1_LOC_66 INVX1_LOC_66/Y VSS VDD INVX1_LOC_66/A INVX1_LOC
XINVX1_LOC_33 INVX1_LOC_33/Y VSS VDD INVX1_LOC_33/A INVX1_LOC
XINVX1_LOC_11 INVX1_LOC_11/Y VSS VDD INVX1_LOC_11/A INVX1_LOC
XINVX1_LOC_99 INVX1_LOC_99/Y VSS VDD INVX1_LOC_99/A INVX1_LOC
XINVX1_LOC_88 INVX1_LOC_88/Y VSS VDD INVX1_LOC_88/A INVX1_LOC
XINVX1_LOC_44 INVX1_LOC_44/Y VSS VDD INVX1_LOC_44/A INVX1_LOC
XINVX1_LOC_77 INVX1_LOC_77/Y VSS VDD INVX1_LOC_77/A INVX1_LOC
XINVX1_LOC_55 INVX1_LOC_55/Y VSS VDD INVX1_LOC_55/A INVX1_LOC
XNAND2X1_LOC_462 NAND2X1_LOC_462/a_36_24# INVX1_LOC_195/A VSS VDD INVX1_LOC_175/Y
+ NAND2X1_LOC_462/B NAND2X1_LOC
XNAND2X1_LOC_473 NAND2X1_LOC_473/a_36_24# INVX1_LOC_201/A VSS VDD NAND2X1_LOC_473/A
+ NAND2X1_LOC_276/Y NAND2X1_LOC
XNAND2X1_LOC_440 NAND2X1_LOC_440/a_36_24# NAND2X1_LOC_468/B VSS VDD NOR2X1_LOC_437/Y
+ INVX1_LOC_182/Y NAND2X1_LOC
XNAND2X1_LOC_495 NAND2X1_LOC_495/a_36_24# NOR2X1_LOC_499/B VSS VDD INVX1_LOC_23/A
+ INVX1_LOC_41/A NAND2X1_LOC
XNAND2X1_LOC_484 NAND2X1_LOC_484/a_36_24# NOR2X1_LOC_486/B VSS VDD INVX1_LOC_9/A INVX1_LOC_23/A
+ NAND2X1_LOC
XNAND2X1_LOC_451 NAND2X1_LOC_451/a_36_24# NAND2X1_LOC_451/Y VSS VDD NOR2X1_LOC_428/Y
+ NOR2X1_LOC_430/Y NAND2X1_LOC
XINVX1_LOC_306 INVX1_LOC_306/Y VSS VDD INVX1_LOC_306/A INVX1_LOC
XNAND2X1_LOC_270 NAND2X1_LOC_270/a_36_24# NOR2X1_LOC_368/A VSS VDD INVX1_LOC_16/A
+ INVX1_LOC_24/A NAND2X1_LOC
XNOR2X1_LOC_708 NOR2X1_LOC_708/a_36_216# NOR2X1_LOC_708/Y VSS VDD NOR2X1_LOC_708/A
+ NOR2X1_LOC_708/B NOR2X1_LOC
XNAND2X1_LOC_281 NAND2X1_LOC_281/a_36_24# NOR2X1_LOC_285/B VSS VDD INVX1_LOC_1/A INVX1_LOC_117/A
+ NAND2X1_LOC
XNAND2X1_LOC_292 NAND2X1_LOC_292/a_36_24# NOR2X1_LOC_346/B VSS VDD INVX1_LOC_30/Y
+ INVX1_LOC_87/A NAND2X1_LOC
XNOR2X1_LOC_719 NOR2X1_LOC_719/a_36_216# INVX1_LOC_284/A VSS VDD NOR2X1_LOC_719/A
+ NOR2X1_LOC_719/B NOR2X1_LOC
XINVX1_LOC_169 INVX1_LOC_169/Y VSS VDD INVX1_LOC_169/A INVX1_LOC
XINVX1_LOC_158 INVX1_LOC_158/Y VSS VDD INVX1_LOC_158/A INVX1_LOC
XINVX1_LOC_125 INVX1_LOC_125/Y VSS VDD INVX1_LOC_125/A INVX1_LOC
XINVX1_LOC_147 INVX1_LOC_147/Y VSS VDD INVX1_LOC_147/A INVX1_LOC
XINVX1_LOC_136 INVX1_LOC_136/Y VSS VDD INVX1_LOC_136/A INVX1_LOC
XINVX1_LOC_114 INVX1_LOC_114/Y VSS VDD INVX1_LOC_114/A INVX1_LOC
XINVX1_LOC_103 INVX1_LOC_103/Y VSS VDD INVX1_LOC_103/A INVX1_LOC
XNOR2X1_LOC_505 NOR2X1_LOC_505/a_36_216# NOR2X1_LOC_505/Y VSS VDD NOR2X1_LOC_45/B
+ INVX1_LOC_16/A NOR2X1_LOC
XNOR2X1_LOC_549 NOR2X1_LOC_549/a_36_216# NOR2X1_LOC_565/B VSS VDD NOR2X1_LOC_548/Y
+ INVX1_LOC_220/Y NOR2X1_LOC
XNOR2X1_LOC_527 NOR2X1_LOC_527/a_36_216# NOR2X1_LOC_527/Y VSS VDD NOR2X1_LOC_111/A
+ INVX1_LOC_50/A NOR2X1_LOC
XNOR2X1_LOC_538 NOR2X1_LOC_538/a_36_216# NOR2X1_LOC_538/Y VSS VDD NOR2X1_LOC_336/B
+ NOR2X1_LOC_538/B NOR2X1_LOC
XNOR2X1_LOC_516 NOR2X1_LOC_516/a_36_216# NOR2X1_LOC_516/Y VSS VDD INVX1_LOC_216/Y
+ NOR2X1_LOC_516/B NOR2X1_LOC
XNOR2X1_LOC_302 NOR2X1_LOC_302/a_36_216# NOR2X1_LOC_302/Y VSS VDD NOR2X1_LOC_302/A
+ NOR2X1_LOC_302/B NOR2X1_LOC
XNOR2X1_LOC_313 NOR2X1_LOC_313/a_36_216# NOR2X1_LOC_313/Y VSS VDD NOR2X1_LOC_91/A
+ INVX1_LOC_54/A NOR2X1_LOC
XNOR2X1_LOC_324 NOR2X1_LOC_324/a_36_216# NOR2X1_LOC_324/Y VSS VDD NOR2X1_LOC_324/A
+ NOR2X1_LOC_324/B NOR2X1_LOC
XNOR2X1_LOC_379 NOR2X1_LOC_379/a_36_216# NOR2X1_LOC_379/Y VSS VDD INVX1_LOC_19/A INVX1_LOC_11/A
+ NOR2X1_LOC
XNOR2X1_LOC_357 NOR2X1_LOC_357/a_36_216# NOR2X1_LOC_357/Y VSS VDD NOR2X1_LOC_353/Y
+ NOR2X1_LOC_352/Y NOR2X1_LOC
XNOR2X1_LOC_335 NOR2X1_LOC_335/a_36_216# INVX1_LOC_150/A VSS VDD NOR2X1_LOC_335/A
+ NOR2X1_LOC_335/B NOR2X1_LOC
XNOR2X1_LOC_346 NOR2X1_LOC_346/a_36_216# NOR2X1_LOC_346/Y VSS VDD NOR2X1_LOC_346/A
+ NOR2X1_LOC_346/B NOR2X1_LOC
XNOR2X1_LOC_368 NOR2X1_LOC_368/a_36_216# NOR2X1_LOC_368/Y VSS VDD NOR2X1_LOC_368/A
+ INVX1_LOC_6/A NOR2X1_LOC
XNAND2X1_LOC_836 NAND2X1_LOC_836/a_36_24# NAND2X1_LOC_836/Y VSS VDD NOR2X1_LOC_823/Y
+ NOR2X1_LOC_824/Y NAND2X1_LOC
XNAND2X1_LOC_825 NAND2X1_LOC_825/a_36_24# NOR2X1_LOC_837/B VSS VDD INVX1_LOC_33/A
+ NAND2X1_LOC_96/A NAND2X1_LOC
XNAND2X1_LOC_847 NAND2X1_LOC_847/a_36_24# INVX1_LOC_315/A VSS VDD NOR2X1_LOC_817/Y
+ NOR2X1_LOC_820/Y NAND2X1_LOC
XNAND2X1_LOC_858 NAND2X1_LOC_858/a_36_24# NAND2X1_LOC_862/A VSS VDD NAND2X1_LOC_850/Y
+ NAND2X1_LOC_858/B NAND2X1_LOC
XNAND2X1_LOC_803 NAND2X1_LOC_803/a_36_24# NAND2X1_LOC_808/A VSS VDD NAND2X1_LOC_796/Y
+ NAND2X1_LOC_803/B NAND2X1_LOC
XNAND2X1_LOC_814 NAND2X1_LOC_814/a_36_24# NOR2X1_LOC_815/A VSS VDD INVX1_LOC_63/Y
+ NOR2X1_LOC_226/A NAND2X1_LOC
XNOR2X1_LOC_31 NOR2X1_LOC_31/a_36_216# INVX1_LOC_22/A VSS VDD NOR2X1_LOC_30/Y NOR2X1_LOC_1/Y
+ NOR2X1_LOC
XNOR2X1_LOC_64 NOR2X1_LOC_64/a_36_216# INVX1_LOC_50/A VSS VDD NOR2X1_LOC_51/A NOR2X1_LOC_36/A
+ NOR2X1_LOC
XNOR2X1_LOC_53 NOR2X1_LOC_53/a_36_216# NOR2X1_LOC_53/Y VSS VDD NOR2X1_LOC_51/A INPUT_5
+ NOR2X1_LOC
XNOR2X1_LOC_20 NOR2X1_LOC_20/a_36_216# NOR2X1_LOC_20/Y VSS VDD NOR2X1_LOC_19/Y INVX1_LOC_15/Y
+ NOR2X1_LOC
XNOR2X1_LOC_42 NOR2X1_LOC_42/a_36_216# INVX1_LOC_32/A VSS VDD INVX1_LOC_26/A D_INPUT_1
+ NOR2X1_LOC
XNOR2X1_LOC_75 NOR2X1_LOC_75/a_36_216# NOR2X1_LOC_75/Y VSS VDD INVX1_LOC_46/A NOR2X1_LOC_45/B
+ NOR2X1_LOC
XNOR2X1_LOC_97 NOR2X1_LOC_97/a_36_216# NOR2X1_LOC_99/B VSS VDD NOR2X1_LOC_97/A NOR2X1_LOC_97/B
+ NOR2X1_LOC
XNOR2X1_LOC_86 NOR2X1_LOC_86/a_36_216# NOR2X1_LOC_86/Y VSS VDD NOR2X1_LOC_86/A D_INPUT_0
+ NOR2X1_LOC
XNAND2X1_LOC_8 NAND2X1_LOC_8/a_36_24# INVX1_LOC_7/A VSS VDD INPUT_2 D_INPUT_3
+ NAND2X1_LOC
XNOR2X1_LOC_154 NOR2X1_LOC_154/a_36_216# NOR2X1_LOC_156/B VSS VDD INVX1_LOC_27/A INVX1_LOC_5/A
+ NOR2X1_LOC
XNOR2X1_LOC_110 NOR2X1_LOC_110/a_36_216# NOR2X1_LOC_111/A VSS VDD INVX1_LOC_14/A INPUT_0
+ NOR2X1_LOC
XNOR2X1_LOC_165 NOR2X1_LOC_165/a_36_216# NOR2X1_LOC_165/Y VSS VDD NOR2X1_LOC_74/A
+ INVX1_LOC_38/A NOR2X1_LOC
XNOR2X1_LOC_176 NOR2X1_LOC_176/a_36_216# NOR2X1_LOC_176/Y VSS VDD NOR2X1_LOC_91/A
+ INVX1_LOC_20/A NOR2X1_LOC
XNOR2X1_LOC_143 NOR2X1_LOC_143/a_36_216# INVX1_LOC_84/A VSS VDD INVX1_LOC_8/A INPUT_1
+ NOR2X1_LOC
XNOR2X1_LOC_121 NOR2X1_LOC_121/a_36_216# NOR2X1_LOC_121/Y VSS VDD NOR2X1_LOC_121/A
+ INVX1_LOC_72/Y NOR2X1_LOC
XNOR2X1_LOC_132 NOR2X1_LOC_132/a_36_216# NOR2X1_LOC_132/Y VSS VDD INVX1_LOC_58/A NOR2X1_LOC_91/A
+ NOR2X1_LOC
XNOR2X1_LOC_198 NOR2X1_LOC_198/a_36_216# NOR2X1_LOC_208/A VSS VDD NOR2X1_LOC_197/Y
+ INVX1_LOC_44/Y NOR2X1_LOC
XNOR2X1_LOC_187 NOR2X1_LOC_187/a_36_216# NOR2X1_LOC_187/Y VSS VDD NOR2X1_LOC_331/B
+ INVX1_LOC_29/Y NOR2X1_LOC
XNAND2X1_LOC_611 NAND2X1_LOC_611/a_36_24# INVX1_LOC_251/A VSS VDD INVX1_LOC_3/A INVX1_LOC_40/A
+ NAND2X1_LOC
XNAND2X1_LOC_600 NAND2X1_LOC_600/a_36_24# NOR2X1_LOC_602/B VSS VDD INVX1_LOC_21/A
+ INVX1_LOC_63/A NAND2X1_LOC
XNAND2X1_LOC_633 NAND2X1_LOC_633/a_36_24# NAND2X1_LOC_633/Y VSS VDD INVX1_LOC_70/A
+ NOR2X1_LOC_278/A NAND2X1_LOC
XNAND2X1_LOC_666 NAND2X1_LOC_666/a_36_24# NOR2X1_LOC_719/A VSS VDD INVX1_LOC_16/Y
+ NOR2X1_LOC_121/A NAND2X1_LOC
XNAND2X1_LOC_622 NAND2X1_LOC_622/a_36_24# NAND2X1_LOC_624/A VSS VDD INVX1_LOC_253/Y
+ NAND2X1_LOC_622/B NAND2X1_LOC
XNAND2X1_LOC_688 NAND2X1_LOC_688/a_36_24# NOR2X1_LOC_689/A VSS VDD INVX1_LOC_28/A
+ INVX1_LOC_136/A NAND2X1_LOC
XNAND2X1_LOC_699 NAND2X1_LOC_699/a_36_24# NOR2X1_LOC_709/A VSS VDD INVX1_LOC_14/Y
+ INVX1_LOC_89/A NAND2X1_LOC
XNAND2X1_LOC_655 NAND2X1_LOC_655/a_36_24# NAND2X1_LOC_660/A VSS VDD NAND2X1_LOC_655/A
+ NAND2X1_LOC_655/B NAND2X1_LOC
XNAND2X1_LOC_644 NAND2X1_LOC_644/a_36_24# NAND2X1_LOC_648/A VSS VDD NOR2X1_LOC_597/Y
+ NOR2X1_LOC_599/Y NAND2X1_LOC
XNAND2X1_LOC_677 NAND2X1_LOC_677/a_36_24# NOR2X1_LOC_678/A VSS VDD INVX1_LOC_19/A
+ INVX1_LOC_77/A NAND2X1_LOC
XINVX1_LOC_12 INVX1_LOC_12/Y VSS VDD INVX1_LOC_12/A INVX1_LOC
XINVX1_LOC_89 INVX1_LOC_89/Y VSS VDD INVX1_LOC_89/A INVX1_LOC
XINVX1_LOC_34 INVX1_LOC_34/Y VSS VDD INVX1_LOC_34/A INVX1_LOC
XINVX1_LOC_56 INVX1_LOC_56/Y VSS VDD INVX1_LOC_56/A INVX1_LOC
XINVX1_LOC_23 INVX1_LOC_23/Y VSS VDD INVX1_LOC_23/A INVX1_LOC
XINVX1_LOC_45 INVX1_LOC_45/Y VSS VDD INVX1_LOC_45/A INVX1_LOC
XINVX1_LOC_67 INVX1_LOC_67/Y VSS VDD INVX1_LOC_67/A INVX1_LOC
XINVX1_LOC_78 INVX1_LOC_78/Y VSS VDD INVX1_LOC_78/A INVX1_LOC
XNAND2X1_LOC_441 NAND2X1_LOC_441/a_36_24# NOR2X1_LOC_545/B VSS VDD INVX1_LOC_29/A
+ NOR2X1_LOC_68/A NAND2X1_LOC
XNAND2X1_LOC_463 NAND2X1_LOC_463/a_36_24# INVX1_LOC_197/A VSS VDD INVX1_LOC_194/Y
+ NAND2X1_LOC_463/B NAND2X1_LOC
XNAND2X1_LOC_430 NAND2X1_LOC_430/a_36_24# NOR2X1_LOC_451/A VSS VDD INVX1_LOC_91/A
+ NAND2X1_LOC_430/B NAND2X1_LOC
XNAND2X1_LOC_452 NAND2X1_LOC_452/a_36_24# NAND2X1_LOC_452/Y VSS VDD INVX1_LOC_192/Y
+ NAND2X1_LOC_451/Y NAND2X1_LOC
XNAND2X1_LOC_474 NAND2X1_LOC_474/a_36_24# NAND2X1_LOC_474/Y VSS VDD NAND2X1_LOC_392/Y
+ NAND2X1_LOC_573/A NAND2X1_LOC
XNAND2X1_LOC_496 NAND2X1_LOC_496/a_36_24# NOR2X1_LOC_778/A VSS VDD INVX1_LOC_15/A
+ INVX1_LOC_41/A NAND2X1_LOC
XNAND2X1_LOC_485 NAND2X1_LOC_485/a_36_24# NOR2X1_LOC_705/B VSS VDD INVX1_LOC_33/A
+ NOR2X1_LOC_590/A NAND2X1_LOC
XINVX1_LOC_307 INVX1_LOC_307/Y VSS VDD INVX1_LOC_307/A INVX1_LOC
XNAND2X1_LOC_282 NAND2X1_LOC_282/a_36_24# NOR2X1_LOC_285/A VSS VDD NOR2X1_LOC_590/A
+ INVX1_LOC_89/A NAND2X1_LOC
XNAND2X1_LOC_293 NAND2X1_LOC_293/a_36_24# INVX1_LOC_135/A VSS VDD INPUT_1 INVX1_LOC_3/A
+ NAND2X1_LOC
XNAND2X1_LOC_271 NAND2X1_LOC_271/a_36_24# NOR2X1_LOC_276/B VSS VDD NOR2X1_LOC_269/Y
+ NOR2X1_LOC_270/Y NAND2X1_LOC
XNAND2X1_LOC_260 NAND2X1_LOC_260/a_36_24# NOR2X1_LOC_261/A VSS VDD INVX1_LOC_12/A
+ INVX1_LOC_90/A NAND2X1_LOC
XNOR2X1_LOC_709 NOR2X1_LOC_709/a_36_216# INVX1_LOC_278/A VSS VDD NOR2X1_LOC_709/A
+ NOR2X1_LOC_709/B NOR2X1_LOC
XINVX1_LOC_137 INVX1_LOC_137/Y VSS VDD INVX1_LOC_137/A INVX1_LOC
XINVX1_LOC_148 INVX1_LOC_148/Y VSS VDD INVX1_LOC_148/A INVX1_LOC
XINVX1_LOC_104 INVX1_LOC_104/Y VSS VDD INVX1_LOC_104/A INVX1_LOC
XINVX1_LOC_126 INVX1_LOC_126/Y VSS VDD INVX1_LOC_126/A INVX1_LOC
XINVX1_LOC_159 INVX1_LOC_159/Y VSS VDD INVX1_LOC_159/A INVX1_LOC
XINVX1_LOC_115 INVX1_LOC_115/Y VSS VDD INVX1_LOC_115/A INVX1_LOC
XNOR2X1_LOC_506 NOR2X1_LOC_506/a_36_216# NOR2X1_LOC_506/Y VSS VDD NOR2X1_LOC_447/B
+ INVX1_LOC_119/A NOR2X1_LOC
XNOR2X1_LOC_517 NOR2X1_LOC_517/a_36_216# NOR2X1_LOC_517/Y VSS VDD NOR2X1_LOC_667/A
+ INVX1_LOC_22/A NOR2X1_LOC
XNOR2X1_LOC_539 NOR2X1_LOC_539/a_36_216# NOR2X1_LOC_799/B VSS VDD NOR2X1_LOC_538/Y
+ NOR2X1_LOC_537/Y NOR2X1_LOC
XNOR2X1_LOC_528 NOR2X1_LOC_528/a_36_216# NOR2X1_LOC_528/Y VSS VDD INVX1_LOC_34/A INVX1_LOC_6/A
+ NOR2X1_LOC
XNOR2X1_LOC_303 NOR2X1_LOC_303/a_36_216# NOR2X1_LOC_303/Y VSS VDD NOR2X1_LOC_302/Y
+ INVX1_LOC_139/Y NOR2X1_LOC
XNOR2X1_LOC_314 NOR2X1_LOC_314/a_36_216# NOR2X1_LOC_314/Y VSS VDD INVX1_LOC_50/A NOR2X1_LOC_15/Y
+ NOR2X1_LOC
XNOR2X1_LOC_358 NOR2X1_LOC_358/a_36_216# NOR2X1_LOC_364/A VSS VDD NOR2X1_LOC_351/Y
+ INVX1_LOC_157/Y NOR2X1_LOC
XNOR2X1_LOC_325 NOR2X1_LOC_325/a_36_216# NOR2X1_LOC_325/Y VSS VDD NOR2X1_LOC_325/A
+ NOR2X1_LOC_374/B NOR2X1_LOC
XNOR2X1_LOC_336 NOR2X1_LOC_336/a_36_216# NOR2X1_LOC_337/A VSS VDD NOR2X1_LOC_703/A
+ NOR2X1_LOC_336/B NOR2X1_LOC
XNOR2X1_LOC_347 NOR2X1_LOC_347/a_36_216# NOR2X1_LOC_360/A VSS VDD NOR2X1_LOC_346/Y
+ INVX1_LOC_138/Y NOR2X1_LOC
XNOR2X1_LOC_369 NOR2X1_LOC_369/a_36_216# NOR2X1_LOC_369/Y VSS VDD INVX1_LOC_71/Y INVX1_LOC_18/A
+ NOR2X1_LOC
XNAND2X1_LOC_804 NAND2X1_LOC_804/a_36_24# NAND2X1_LOC_804/Y VSS VDD NAND2X1_LOC_804/A
+ NAND2X1_LOC_795/Y NAND2X1_LOC
XNAND2X1_LOC_826 NAND2X1_LOC_826/a_36_24# NOR2X1_LOC_837/A VSS VDD INVX1_LOC_41/A
+ INVX1_LOC_57/A NAND2X1_LOC
XNAND2X1_LOC_837 NAND2X1_LOC_837/a_36_24# NAND2X1_LOC_837/Y VSS VDD NOR2X1_LOC_825/Y
+ NOR2X1_LOC_826/Y NAND2X1_LOC
XNAND2X1_LOC_859 NAND2X1_LOC_859/a_36_24# NAND2X1_LOC_859/Y VSS VDD NAND2X1_LOC_848/Y
+ NAND2X1_LOC_859/B NAND2X1_LOC
XNAND2X1_LOC_848 NAND2X1_LOC_848/a_36_24# NAND2X1_LOC_848/Y VSS VDD NAND2X1_LOC_848/A
+ INVX1_LOC_316/Y NAND2X1_LOC
XNAND2X1_LOC_815 NAND2X1_LOC_815/a_36_24# NOR2X1_LOC_846/B VSS VDD INVX1_LOC_2/Y NOR2X1_LOC_814/Y
+ NAND2X1_LOC
XNOR2X1_LOC_21 NOR2X1_LOC_21/a_36_216# NOR2X1_LOC_36/A VSS VDD INPUT_5 D_INPUT_4
+ NOR2X1_LOC
XNOR2X1_LOC_43 NOR2X1_LOC_43/a_36_216# NOR2X1_LOC_43/Y VSS VDD INVX1_LOC_32/A INVX1_LOC_18/A
+ NOR2X1_LOC
XNOR2X1_LOC_65 NOR2X1_LOC_65/a_36_216# NOR2X1_LOC_65/Y VSS VDD INVX1_LOC_49/Y NOR2X1_LOC_65/B
+ NOR2X1_LOC
XNOR2X1_LOC_54 NOR2X1_LOC_54/a_36_216# INVX1_LOC_40/A VSS VDD D_INPUT_1 D_INPUT_0
+ NOR2X1_LOC
XNOR2X1_LOC_87 NOR2X1_LOC_87/a_36_216# NOR2X1_LOC_87/Y VSS VDD NOR2X1_LOC_68/A NOR2X1_LOC_87/B
+ NOR2X1_LOC
XNOR2X1_LOC_32 NOR2X1_LOC_32/a_36_216# NOR2X1_LOC_32/Y VSS VDD INVX1_LOC_22/A NOR2X1_LOC_32/B
+ NOR2X1_LOC
XNOR2X1_LOC_76 NOR2X1_LOC_76/a_36_216# INVX1_LOC_56/A VSS VDD NOR2X1_LOC_76/A NOR2X1_LOC_76/B
+ NOR2X1_LOC
XNOR2X1_LOC_10 NOR2X1_LOC_10/a_36_216# INVX1_LOC_10/A VSS VDD NOR2X1_LOC_9/Y INVX1_LOC_8/A
+ NOR2X1_LOC
XNOR2X1_LOC_98 NOR2X1_LOC_98/a_36_216# INVX1_LOC_60/A VSS VDD NOR2X1_LOC_98/A NOR2X1_LOC_98/B
+ NOR2X1_LOC
XNAND2X1_LOC_9 NAND2X1_LOC_9/a_36_24# NAND2X1_LOC_9/Y VSS VDD D_INPUT_0 D_INPUT_1
+ NAND2X1_LOC
XNOR2X1_LOC_155 NOR2X1_LOC_155/a_36_216# NOR2X1_LOC_156/A VSS VDD NOR2X1_LOC_155/A
+ NOR2X1_LOC_68/A NOR2X1_LOC
XNOR2X1_LOC_144 NOR2X1_LOC_144/a_36_216# NOR2X1_LOC_144/Y VSS VDD INVX1_LOC_84/A INVX1_LOC_46/A
+ NOR2X1_LOC
XNOR2X1_LOC_122 NOR2X1_LOC_122/a_36_216# NOR2X1_LOC_122/Y VSS VDD NOR2X1_LOC_122/A
+ INVX1_LOC_34/A NOR2X1_LOC
XNOR2X1_LOC_111 NOR2X1_LOC_111/a_36_216# NOR2X1_LOC_111/Y VSS VDD NOR2X1_LOC_111/A
+ INVX1_LOC_22/A NOR2X1_LOC
XNOR2X1_LOC_188 NOR2X1_LOC_188/a_36_216# NOR2X1_LOC_188/Y VSS VDD NOR2X1_LOC_188/A
+ INVX1_LOC_28/Y NOR2X1_LOC
XNOR2X1_LOC_166 NOR2X1_LOC_166/a_36_216# NOR2X1_LOC_166/Y VSS VDD INVX1_LOC_30/A NOR2X1_LOC_15/Y
+ NOR2X1_LOC
XNOR2X1_LOC_199 NOR2X1_LOC_199/a_36_216# INVX1_LOC_108/A VSS VDD NOR2X1_LOC_196/Y
+ NOR2X1_LOC_199/B NOR2X1_LOC
XNOR2X1_LOC_100 NOR2X1_LOC_100/a_36_216# INVX1_LOC_62/A VSS VDD NOR2X1_LOC_100/A NAND2X1_LOC_86/Y
+ NOR2X1_LOC
XNOR2X1_LOC_133 NOR2X1_LOC_133/a_36_216# INVX1_LOC_78/A VSS VDD NOR2X1_LOC_38/B INVX1_LOC_8/A
+ NOR2X1_LOC
XNOR2X1_LOC_177 NOR2X1_LOC_177/a_36_216# NOR2X1_LOC_177/Y VSS VDD INVX1_LOC_54/A NOR2X1_LOC_52/B
+ NOR2X1_LOC
XNAND2X1_LOC_623 NAND2X1_LOC_623/a_36_24# NAND2X1_LOC_624/B VSS VDD NOR2X1_LOC_615/Y
+ NAND2X1_LOC_623/B NAND2X1_LOC
XNAND2X1_LOC_634 NAND2X1_LOC_634/a_36_24# NAND2X1_LOC_634/Y VSS VDD NOR2X1_LOC_290/Y
+ NOR2X1_LOC_690/A NAND2X1_LOC
XNAND2X1_LOC_612 NAND2X1_LOC_612/a_36_24# NOR2X1_LOC_647/B VSS VDD NOR2X1_LOC_610/Y
+ INVX1_LOC_252/Y NAND2X1_LOC
XNAND2X1_LOC_601 NAND2X1_LOC_601/a_36_24# NOR2X1_LOC_602/A VSS VDD NOR2X1_LOC_78/B
+ INVX1_LOC_35/A NAND2X1_LOC
XNAND2X1_LOC_645 NAND2X1_LOC_645/a_36_24# INVX1_LOC_263/A VSS VDD INVX1_LOC_247/A
+ INVX1_LOC_249/A NAND2X1_LOC
XINVX1_LOC_13 INVX1_LOC_13/Y VSS VDD INVX1_LOC_13/A INVX1_LOC
XINVX1_LOC_24 INVX1_LOC_24/Y VSS VDD INVX1_LOC_24/A INVX1_LOC
XNAND2X1_LOC_689 NAND2X1_LOC_689/a_36_24# NOR2X1_LOC_691/B VSS VDD INVX1_LOC_22/Y
+ NOR2X1_LOC_688/Y NAND2X1_LOC
XNAND2X1_LOC_667 NAND2X1_LOC_667/a_36_24# NOR2X1_LOC_720/B VSS VDD INVX1_LOC_50/Y
+ NOR2X1_LOC_264/Y NAND2X1_LOC
XNAND2X1_LOC_656 NAND2X1_LOC_656/a_36_24# NAND2X1_LOC_656/Y VSS VDD NAND2X1_LOC_656/A
+ NAND2X1_LOC_656/B NAND2X1_LOC
XNAND2X1_LOC_678 NAND2X1_LOC_678/a_36_24# INVX1_LOC_271/A VSS VDD INVX1_LOC_12/A NOR2X1_LOC_677/Y
+ NAND2X1_LOC
XINVX1_LOC_68 INVX1_LOC_68/Y VSS VDD INVX1_LOC_68/A INVX1_LOC
XINVX1_LOC_46 INVX1_LOC_46/Y VSS VDD INVX1_LOC_46/A INVX1_LOC
XINVX1_LOC_35 INVX1_LOC_35/Y VSS VDD INVX1_LOC_35/A INVX1_LOC
XINVX1_LOC_57 INVX1_LOC_57/Y VSS VDD INVX1_LOC_57/A INVX1_LOC
XINVX1_LOC_79 INVX1_LOC_79/Y VSS VDD INVX1_LOC_79/A INVX1_LOC
XNAND2X1_LOC_486 NAND2X1_LOC_486/a_36_24# NAND2X1_LOC_787/B VSS VDD NOR2X1_LOC_484/Y
+ NOR2X1_LOC_485/Y NAND2X1_LOC
XNAND2X1_LOC_464 NAND2X1_LOC_464/a_36_24# NAND2X1_LOC_464/Y VSS VDD NAND2X1_LOC_464/A
+ NAND2X1_LOC_464/B NAND2X1_LOC
XNAND2X1_LOC_442 NAND2X1_LOC_442/a_36_24# INVX1_LOC_183/A VSS VDD INVX1_LOC_29/A INVX1_LOC_63/A
+ NAND2X1_LOC
XNAND2X1_LOC_431 NAND2X1_LOC_431/a_36_24# NOR2X1_LOC_434/A VSS VDD INVX1_LOC_53/A
+ INVX1_LOC_117/A NAND2X1_LOC
XNAND2X1_LOC_475 NAND2X1_LOC_475/a_36_24# NAND2X1_LOC_475/Y VSS VDD INVX1_LOC_171/Y
+ NAND2X1_LOC_474/Y NAND2X1_LOC
XNAND2X1_LOC_497 NAND2X1_LOC_497/a_36_24# NOR2X1_LOC_500/B VSS VDD INVX1_LOC_18/Y
+ NAND2X1_LOC_72/B NAND2X1_LOC
XNAND2X1_LOC_453 NAND2X1_LOC_453/a_36_24# NAND2X1_LOC_466/A VSS VDD NAND2X1_LOC_453/A
+ INVX1_LOC_190/Y NAND2X1_LOC
XNAND2X1_LOC_420 NAND2X1_LOC_420/a_36_24# NOR2X1_LOC_447/A VSS VDD INVX1_LOC_57/A
+ NOR2X1_LOC_590/A NAND2X1_LOC
XINVX1_LOC_308 INVX1_LOC_308/Y VSS VDD INVX1_LOC_308/A INVX1_LOC
XNAND2X1_LOC_250 NAND2X1_LOC_250/a_36_24# NOR2X1_LOC_343/B VSS VDD INVX1_LOC_50/Y
+ NOR2X1_LOC_249/Y NAND2X1_LOC
XNAND2X1_LOC_261 NAND2X1_LOC_261/a_36_24# NOR2X1_LOC_345/A VSS VDD INVX1_LOC_64/Y
+ NOR2X1_LOC_260/Y NAND2X1_LOC
XNAND2X1_LOC_272 NAND2X1_LOC_272/a_36_24# NOR2X1_LOC_274/B VSS VDD INVX1_LOC_21/A
+ INVX1_LOC_31/A NAND2X1_LOC
XNAND2X1_LOC_283 NAND2X1_LOC_283/a_36_24# INVX1_LOC_131/A VSS VDD INVX1_LOC_19/A NOR2X1_LOC_814/A
+ NAND2X1_LOC
XNAND2X1_LOC_294 NAND2X1_LOC_294/a_36_24# NOR2X1_LOC_481/A VSS VDD INVX1_LOC_10/A
+ INVX1_LOC_136/A NAND2X1_LOC
XINVX1_LOC_116 INVX1_LOC_116/Y VSS VDD INVX1_LOC_116/A INVX1_LOC
XINVX1_LOC_105 INVX1_LOC_105/Y VSS VDD INVX1_LOC_105/A INVX1_LOC
XINVX1_LOC_138 INVX1_LOC_138/Y VSS VDD INVX1_LOC_138/A INVX1_LOC
XINVX1_LOC_127 INVX1_LOC_127/Y VSS VDD INVX1_LOC_127/A INVX1_LOC
XINVX1_LOC_149 INVX1_LOC_149/Y VSS VDD INVX1_LOC_149/A INVX1_LOC
XNOR2X1_LOC_518 NOR2X1_LOC_518/a_36_216# NOR2X1_LOC_518/Y VSS VDD NOR2X1_LOC_74/A
+ INVX1_LOC_50/A NOR2X1_LOC
XNOR2X1_LOC_507 NOR2X1_LOC_507/a_36_216# INVX1_LOC_210/A VSS VDD NOR2X1_LOC_507/A
+ NOR2X1_LOC_507/B NOR2X1_LOC
XNOR2X1_LOC_529 NOR2X1_LOC_529/a_36_216# NOR2X1_LOC_529/Y VSS VDD INVX1_LOC_20/A D_INPUT_3
+ NOR2X1_LOC
XNOR2X1_LOC_304 NOR2X1_LOC_304/a_36_216# NOR2X1_LOC_304/Y VSS VDD INVX1_LOC_118/A
+ NOR2X1_LOC_53/Y NOR2X1_LOC
XNOR2X1_LOC_359 NOR2X1_LOC_359/a_36_216# NOR2X1_LOC_359/Y VSS VDD INVX1_LOC_155/Y
+ NOR2X1_LOC_348/Y NOR2X1_LOC
XNOR2X1_LOC_348 NOR2X1_LOC_348/a_36_216# NOR2X1_LOC_348/Y VSS VDD INVX1_LOC_153/Y
+ NOR2X1_LOC_348/B NOR2X1_LOC
XNOR2X1_LOC_326 NOR2X1_LOC_326/a_36_216# NOR2X1_LOC_326/Y VSS VDD NOR2X1_LOC_325/Y
+ NOR2X1_LOC_324/Y NOR2X1_LOC
XNOR2X1_LOC_337 NOR2X1_LOC_337/a_36_216# NOR2X1_LOC_337/Y VSS VDD NOR2X1_LOC_337/A
+ INVX1_LOC_149/Y NOR2X1_LOC
XNOR2X1_LOC_315 NOR2X1_LOC_315/a_36_216# NOR2X1_LOC_315/Y VSS VDD INVX1_LOC_78/A INVX1_LOC_22/A
+ NOR2X1_LOC
XNAND2X1_LOC_827 NAND2X1_LOC_827/a_36_24# INVX1_LOC_309/A VSS VDD INVX1_LOC_31/A INVX1_LOC_89/A
+ NAND2X1_LOC
XNAND2X1_LOC_816 NAND2X1_LOC_816/a_36_24# NOR2X1_LOC_846/A VSS VDD INVX1_LOC_38/Y
+ NOR2X1_LOC_188/A NAND2X1_LOC
XNAND2X1_LOC_805 NAND2X1_LOC_805/a_36_24# NAND2X1_LOC_807/A VSS VDD INVX1_LOC_308/Y
+ NAND2X1_LOC_793/Y NAND2X1_LOC
XNAND2X1_LOC_838 NAND2X1_LOC_838/a_36_24# NAND2X1_LOC_838/Y VSS VDD INVX1_LOC_309/Y
+ NAND2X1_LOC_837/Y NAND2X1_LOC
XNAND2X1_LOC_849 NAND2X1_LOC_849/a_36_24# NAND2X1_LOC_859/B VSS VDD NAND2X1_LOC_849/A
+ NAND2X1_LOC_849/B NAND2X1_LOC
XNOR2X1_LOC_860 NOR2X1_LOC_860/a_36_216# NOR2X1_LOC_860/Y VSS VDD NOR2X1_LOC_392/Y
+ NOR2X1_LOC_860/B NOR2X1_LOC
XNOR2X1_LOC_22 NOR2X1_LOC_22/a_36_216# INVX1_LOC_18/A VSS VDD NOR2X1_LOC_36/A NOR2X1_LOC_1/Y
+ NOR2X1_LOC
XNOR2X1_LOC_11 NOR2X1_LOC_11/a_36_216# NOR2X1_LOC_11/Y VSS VDD D_INPUT_5 INPUT_4
+ NOR2X1_LOC
XNOR2X1_LOC_44 NOR2X1_LOC_44/a_36_216# INVX1_LOC_34/A VSS VDD NOR2X1_LOC_30/Y NOR2X1_LOC_36/B
+ NOR2X1_LOC
XNOR2X1_LOC_66 NOR2X1_LOC_66/a_36_216# NOR2X1_LOC_66/Y VSS VDD INVX1_LOC_19/A INVX1_LOC_1/A
+ NOR2X1_LOC
XNOR2X1_LOC_33 NOR2X1_LOC_33/a_36_216# NOR2X1_LOC_33/Y VSS VDD NOR2X1_LOC_33/A NOR2X1_LOC_33/B
+ NOR2X1_LOC
XNOR2X1_LOC_99 NOR2X1_LOC_99/a_36_216# NOR2X1_LOC_99/Y VSS VDD INVX1_LOC_59/Y NOR2X1_LOC_99/B
+ NOR2X1_LOC
XNOR2X1_LOC_88 NOR2X1_LOC_88/a_36_216# NOR2X1_LOC_88/Y VSS VDD NOR2X1_LOC_88/A INVX1_LOC_2/A
+ NOR2X1_LOC
XNOR2X1_LOC_77 NOR2X1_LOC_77/a_36_216# NOR2X1_LOC_89/A VSS VDD INVX1_LOC_40/A INVX1_LOC_14/A
+ NOR2X1_LOC
XNOR2X1_LOC_55 NOR2X1_LOC_55/a_36_216# INVX1_LOC_42/A VSS VDD INVX1_LOC_40/A INVX1_LOC_3/Y
+ NOR2X1_LOC
XNOR2X1_LOC_145 NOR2X1_LOC_145/a_36_216# NOR2X1_LOC_145/Y VSS VDD NOR2X1_LOC_89/A
+ INVX1_LOC_38/A NOR2X1_LOC
XNOR2X1_LOC_156 NOR2X1_LOC_156/a_36_216# NOR2X1_LOC_156/Y VSS VDD NOR2X1_LOC_156/A
+ NOR2X1_LOC_156/B NOR2X1_LOC
XNOR2X1_LOC_189 NOR2X1_LOC_189/a_36_216# INVX1_LOC_102/A VSS VDD NOR2X1_LOC_189/A
+ INVX1_LOC_58/A NOR2X1_LOC
XNOR2X1_LOC_167 NOR2X1_LOC_167/a_36_216# NOR2X1_LOC_167/Y VSS VDD INVX1_LOC_92/A INVX1_LOC_50/A
+ NOR2X1_LOC
XNOR2X1_LOC_112 NOR2X1_LOC_112/a_36_216# NOR2X1_LOC_112/Y VSS VDD NOR2X1_LOC_332/B
+ NOR2X1_LOC_112/B NOR2X1_LOC
XNOR2X1_LOC_101 NOR2X1_LOC_101/a_36_216# NOR2X1_LOC_216/B VSS VDD INVX1_LOC_61/Y NOR2X1_LOC_99/Y
+ NOR2X1_LOC
XNOR2X1_LOC_178 NOR2X1_LOC_178/a_36_216# NOR2X1_LOC_178/Y VSS VDD INVX1_LOC_90/A INVX1_LOC_42/A
+ NOR2X1_LOC
XNOR2X1_LOC_134 NOR2X1_LOC_134/a_36_216# NOR2X1_LOC_134/Y VSS VDD INVX1_LOC_78/A INVX1_LOC_57/Y
+ NOR2X1_LOC
XNOR2X1_LOC_123 NOR2X1_LOC_123/a_36_216# NOR2X1_LOC_124/A VSS VDD INVX1_LOC_70/Y NOR2X1_LOC_123/B
+ NOR2X1_LOC
XNAND2X1_LOC_613 NAND2X1_LOC_613/a_36_24# NOR2X1_LOC_620/A VSS VDD INVX1_LOC_29/A
+ INVX1_LOC_41/A NAND2X1_LOC
XNAND2X1_LOC_624 NAND2X1_LOC_624/a_36_24# INVX1_LOC_255/A VSS VDD NAND2X1_LOC_624/A
+ NAND2X1_LOC_624/B NAND2X1_LOC
XNAND2X1_LOC_657 NAND2X1_LOC_657/a_36_24# NAND2X1_LOC_659/A VSS VDD NAND2X1_LOC_141/Y
+ NAND2X1_LOC_574/A NAND2X1_LOC
XNAND2X1_LOC_668 NAND2X1_LOC_668/a_36_24# NOR2X1_LOC_669/A VSS VDD INVX1_LOC_20/A
+ INVX1_LOC_90/A NAND2X1_LOC
XNAND2X1_LOC_646 NAND2X1_LOC_646/a_36_24# NAND2X1_LOC_647/B VSS VDD NOR2X1_LOC_607/Y
+ NOR2X1_LOC_609/Y NAND2X1_LOC
XNAND2X1_LOC_679 NAND2X1_LOC_679/a_36_24# NOR2X1_LOC_728/B VSS VDD NOR2X1_LOC_676/Y
+ INVX1_LOC_271/Y NAND2X1_LOC
XNAND2X1_LOC_602 NAND2X1_LOC_602/a_36_24# INVX1_LOC_247/A VSS VDD NOR2X1_LOC_600/Y
+ NOR2X1_LOC_601/Y NAND2X1_LOC
XNAND2X1_LOC_635 NAND2X1_LOC_635/a_36_24# NAND2X1_LOC_639/A VSS VDD NOR2X1_LOC_428/Y
+ NOR2X1_LOC_582/Y NAND2X1_LOC
XINVX1_LOC_36 INVX1_LOC_36/Y VSS VDD INVX1_LOC_36/A INVX1_LOC
XINVX1_LOC_25 INVX1_LOC_25/Y VSS VDD INVX1_LOC_25/A INVX1_LOC
XINVX1_LOC_47 INVX1_LOC_47/Y VSS VDD INVX1_LOC_47/A INVX1_LOC
XINVX1_LOC_58 INVX1_LOC_58/Y VSS VDD INVX1_LOC_58/A INVX1_LOC
XINVX1_LOC_14 INVX1_LOC_14/Y VSS VDD INVX1_LOC_14/A INVX1_LOC
XINVX1_LOC_69 INVX1_LOC_69/Y VSS VDD INVX1_LOC_69/A INVX1_LOC
XNOR2X1_LOC_690 NOR2X1_LOC_690/a_36_216# NOR2X1_LOC_690/Y VSS VDD NOR2X1_LOC_690/A
+ INPUT_0 NOR2X1_LOC
XNAND2X1_LOC_487 NAND2X1_LOC_487/a_36_24# NOR2X1_LOC_489/B VSS VDD NOR2X1_LOC_160/B
+ INVX1_LOC_57/A NAND2X1_LOC
XNAND2X1_LOC_465 NAND2X1_LOC_465/a_36_24# NAND2X1_LOC_465/Y VSS VDD NAND2X1_LOC_465/A
+ NAND2X1_LOC_456/Y NAND2X1_LOC
XNAND2X1_LOC_410 NAND2X1_LOC_410/a_36_24# NOR2X1_LOC_411/A VSS VDD INVX1_LOC_12/A
+ INVX1_LOC_38/A NAND2X1_LOC
XNAND2X1_LOC_443 NAND2X1_LOC_443/a_36_24# NAND2X1_LOC_444/B VSS VDD NOR2X1_LOC_91/Y
+ NOR2X1_LOC_441/Y NAND2X1_LOC
XNAND2X1_LOC_498 NAND2X1_LOC_498/a_36_24# NOR2X1_LOC_501/B VSS VDD INVX1_LOC_53/A
+ NOR2X1_LOC_188/Y NAND2X1_LOC
XNAND2X1_LOC_454 NAND2X1_LOC_454/a_36_24# NAND2X1_LOC_454/Y VSS VDD INVX1_LOC_188/Y
+ NAND2X1_LOC_447/Y NAND2X1_LOC
XNAND2X1_LOC_476 NAND2X1_LOC_476/a_36_24# NAND2X1_LOC_476/Y VSS VDD NAND2X1_LOC_472/Y
+ INVX1_LOC_202/Y NAND2X1_LOC
XNAND2X1_LOC_432 NAND2X1_LOC_432/a_36_24# NOR2X1_LOC_435/B VSS VDD INVX1_LOC_15/A
+ NOR2X1_LOC_130/A NAND2X1_LOC
XNAND2X1_LOC_421 NAND2X1_LOC_421/a_36_24# NOR2X1_LOC_448/B VSS VDD NOR2X1_LOC_383/B
+ NOR2X1_LOC_596/A NAND2X1_LOC
XINVX1_LOC_309 INVX1_LOC_309/Y VSS VDD INVX1_LOC_309/A INVX1_LOC
XNAND2X1_LOC_262 NAND2X1_LOC_262/a_36_24# NOR2X1_LOC_266/B VSS VDD INVX1_LOC_30/Y
+ NAND2X1_LOC_63/Y NAND2X1_LOC
XNAND2X1_LOC_240 NAND2X1_LOC_240/a_36_24# NAND2X1_LOC_243/B VSS VDD NOR2X1_LOC_232/Y
+ NOR2X1_LOC_234/Y NAND2X1_LOC
XNAND2X1_LOC_295 NAND2X1_LOC_295/a_36_24# NOR2X1_LOC_346/A VSS VDD INVX1_LOC_46/Y
+ NOR2X1_LOC_294/Y NAND2X1_LOC
XNAND2X1_LOC_251 NAND2X1_LOC_251/a_36_24# NOR2X1_LOC_843/B VSS VDD INVX1_LOC_38/Y
+ NOR2X1_LOC_105/Y NAND2X1_LOC
XNAND2X1_LOC_284 NAND2X1_LOC_284/a_36_24# NAND2X1_LOC_287/B VSS VDD NOR2X1_LOC_279/Y
+ NOR2X1_LOC_280/Y NAND2X1_LOC
XNAND2X1_LOC_273 NAND2X1_LOC_273/a_36_24# NOR2X1_LOC_831/B VSS VDD INVX1_LOC_23/A
+ NOR2X1_LOC_155/A NAND2X1_LOC
XINVX1_LOC_106 INVX1_LOC_106/Y VSS VDD INVX1_LOC_106/A INVX1_LOC
XINVX1_LOC_128 INVX1_LOC_128/Y VSS VDD INVX1_LOC_128/A INVX1_LOC
XINVX1_LOC_117 INVX1_LOC_117/Y VSS VDD INVX1_LOC_117/A INVX1_LOC
XINVX1_LOC_139 INVX1_LOC_139/Y VSS VDD INVX1_LOC_139/A INVX1_LOC
XNOR2X1_LOC_508 NOR2X1_LOC_508/a_36_216# NOR2X1_LOC_510/B VSS VDD INVX1_LOC_209/Y
+ NOR2X1_LOC_506/Y NOR2X1_LOC
XNOR2X1_LOC_519 NOR2X1_LOC_519/a_36_216# NOR2X1_LOC_519/Y VSS VDD INVX1_LOC_90/A NOR2X1_LOC_48/B
+ NOR2X1_LOC
XNOR2X1_LOC_338 NOR2X1_LOC_338/a_36_216# NOR2X1_LOC_338/Y VSS VDD NOR2X1_LOC_334/Y
+ INVX1_LOC_147/Y NOR2X1_LOC
XNOR2X1_LOC_305 NOR2X1_LOC_305/a_36_216# NOR2X1_LOC_305/Y VSS VDD NOR2X1_LOC_91/A
+ INVX1_LOC_2/A NOR2X1_LOC
XNOR2X1_LOC_349 NOR2X1_LOC_349/a_36_216# INVX1_LOC_156/A VSS VDD NOR2X1_LOC_349/A
+ NOR2X1_LOC_349/B NOR2X1_LOC
XNOR2X1_LOC_327 NOR2X1_LOC_327/a_36_216# NOR2X1_LOC_405/A VSS VDD NOR2X1_LOC_264/Y
+ NAND2X1_LOC_63/Y NOR2X1_LOC
XNOR2X1_LOC_316 NOR2X1_LOC_316/a_36_216# NOR2X1_LOC_316/Y VSS VDD NOR2X1_LOC_80/Y
+ INVX1_LOC_12/A NOR2X1_LOC
XNAND2X1_LOC_839 NAND2X1_LOC_839/a_36_24# NAND2X1_LOC_839/Y VSS VDD NAND2X1_LOC_839/A
+ NAND2X1_LOC_836/Y NAND2X1_LOC
XNAND2X1_LOC_817 NAND2X1_LOC_817/a_36_24# NOR2X1_LOC_847/B VSS VDD D_INPUT_1 NAND2X1_LOC_381/Y
+ NAND2X1_LOC
XNAND2X1_LOC_806 NAND2X1_LOC_806/a_36_24# NAND2X1_LOC_807/B VSS VDD INVX1_LOC_133/A
+ INVX1_LOC_270/Y NAND2X1_LOC
XNAND2X1_LOC_828 NAND2X1_LOC_828/a_36_24# NOR2X1_LOC_829/A VSS VDD NOR2X1_LOC_409/B
+ NOR2X1_LOC_599/A NAND2X1_LOC
XNOR2X1_LOC_850 NOR2X1_LOC_850/a_36_216# NOR2X1_LOC_858/B VSS VDD INVX1_LOC_313/Y
+ NOR2X1_LOC_850/B NOR2X1_LOC
XNOR2X1_LOC_861 NOR2X1_LOC_861/a_36_216# NOR2X1_LOC_861/Y VSS VDD NOR2X1_LOC_860/Y
+ INVX1_LOC_255/Y NOR2X1_LOC
XNOR2X1_LOC_12 NOR2X1_LOC_12/a_36_216# INVX1_LOC_12/A VSS VDD NOR2X1_LOC_11/Y NOR2X1_LOC_1/Y
+ NOR2X1_LOC
XNOR2X1_LOC_45 NOR2X1_LOC_45/a_36_216# NOR2X1_LOC_45/Y VSS VDD INVX1_LOC_34/A NOR2X1_LOC_45/B
+ NOR2X1_LOC
XNOR2X1_LOC_56 NOR2X1_LOC_56/a_36_216# NOR2X1_LOC_56/Y VSS VDD INVX1_LOC_42/A NOR2X1_LOC_53/Y
+ NOR2X1_LOC
XNOR2X1_LOC_34 NOR2X1_LOC_34/a_36_216# NOR2X1_LOC_34/Y VSS VDD NOR2X1_LOC_34/A NOR2X1_LOC_34/B
+ NOR2X1_LOC
XNOR2X1_LOC_78 NOR2X1_LOC_78/a_36_216# NOR2X1_LOC_78/Y VSS VDD NOR2X1_LOC_78/A NOR2X1_LOC_78/B
+ NOR2X1_LOC
XNOR2X1_LOC_23 NOR2X1_LOC_23/a_36_216# NOR2X1_LOC_45/B VSS VDD INVX1_LOC_14/A NOR2X1_LOC_6/B
+ NOR2X1_LOC
XNOR2X1_LOC_67 NOR2X1_LOC_67/a_36_216# NOR2X1_LOC_67/Y VSS VDD NOR2X1_LOC_67/A INVX1_LOC_42/A
+ NOR2X1_LOC
XNOR2X1_LOC_89 NOR2X1_LOC_89/a_36_216# NOR2X1_LOC_89/Y VSS VDD NOR2X1_LOC_89/A INVX1_LOC_46/A
+ NOR2X1_LOC
XNOR2X1_LOC_113 NOR2X1_LOC_113/a_36_216# NOR2X1_LOC_114/A VSS VDD NOR2X1_LOC_113/A
+ NOR2X1_LOC_113/B NOR2X1_LOC
XNOR2X1_LOC_124 NOR2X1_LOC_124/a_36_216# INVX1_LOC_74/A VSS VDD NOR2X1_LOC_124/A NOR2X1_LOC_124/B
+ NOR2X1_LOC
XNOR2X1_LOC_102 NOR2X1_LOC_102/a_36_216# NOR2X1_LOC_536/A VSS VDD INVX1_LOC_39/Y INVX1_LOC_8/A
+ NOR2X1_LOC
XNOR2X1_LOC_146 NOR2X1_LOC_146/a_36_216# NOR2X1_LOC_146/Y VSS VDD INVX1_LOC_75/Y INVX1_LOC_24/A
+ NOR2X1_LOC
XNOR2X1_LOC_157 NOR2X1_LOC_157/a_36_216# INVX1_LOC_90/A VSS VDD NOR2X1_LOC_36/B NOR2X1_LOC_2/Y
+ NOR2X1_LOC
XNOR2X1_LOC_135 NOR2X1_LOC_135/a_36_216# NOR2X1_LOC_135/Y VSS VDD INVX1_LOC_78/A INVX1_LOC_46/A
+ NOR2X1_LOC
XNOR2X1_LOC_168 NOR2X1_LOC_168/a_36_216# NOR2X1_LOC_168/Y VSS VDD NOR2X1_LOC_168/A
+ NOR2X1_LOC_168/B NOR2X1_LOC
XNOR2X1_LOC_179 NOR2X1_LOC_179/a_36_216# NOR2X1_LOC_179/Y VSS VDD INVX1_LOC_64/A INVX1_LOC_24/A
+ NOR2X1_LOC
XNAND2X1_LOC_614 NAND2X1_LOC_614/a_36_24# NOR2X1_LOC_754/A VSS VDD NOR2X1_LOC_89/A
+ INVX1_LOC_78/A NAND2X1_LOC
XNAND2X1_LOC_669 NAND2X1_LOC_669/a_36_24# NOR2X1_LOC_720/A VSS VDD INVX1_LOC_92/Y
+ NOR2X1_LOC_668/Y NAND2X1_LOC
XNAND2X1_LOC_658 NAND2X1_LOC_658/a_36_24# NAND2X1_LOC_659/B VSS VDD INVX1_LOC_255/A
+ NAND2X1_LOC_735/B NAND2X1_LOC
XNAND2X1_LOC_603 NAND2X1_LOC_603/a_36_24# NOR2X1_LOC_605/B VSS VDD INVX1_LOC_11/A
+ NOR2X1_LOC_68/A NAND2X1_LOC
XNAND2X1_LOC_647 NAND2X1_LOC_647/a_36_24# NAND2X1_LOC_656/B VSS VDD NOR2X1_LOC_612/Y
+ NAND2X1_LOC_647/B NAND2X1_LOC
XNAND2X1_LOC_625 NAND2X1_LOC_625/a_36_24# NOR2X1_LOC_631/A VSS VDD NOR2X1_LOC_66/Y
+ INVX1_LOC_136/Y NAND2X1_LOC
XNAND2X1_LOC_636 NAND2X1_LOC_636/a_36_24# INVX1_LOC_261/A VSS VDD NOR2X1_LOC_583/Y
+ NOR2X1_LOC_584/Y NAND2X1_LOC
XINVX1_LOC_15 INVX1_LOC_15/Y VSS VDD INVX1_LOC_15/A INVX1_LOC
XINVX1_LOC_26 INVX1_LOC_26/Y VSS VDD INVX1_LOC_26/A INVX1_LOC
XINVX1_LOC_48 INVX1_LOC_48/Y VSS VDD INVX1_LOC_48/A INVX1_LOC
XINVX1_LOC_59 INVX1_LOC_59/Y VSS VDD INVX1_LOC_59/A INVX1_LOC
XINVX1_LOC_37 INVX1_LOC_37/Y VSS VDD INVX1_LOC_37/A INVX1_LOC
XNOR2X1_LOC_680 NOR2X1_LOC_680/a_36_216# INVX1_LOC_274/A VSS VDD NOR2X1_LOC_331/B
+ INVX1_LOC_38/A NOR2X1_LOC
XNOR2X1_LOC_691 NOR2X1_LOC_691/a_36_216# NOR2X1_LOC_729/A VSS VDD NOR2X1_LOC_691/A
+ NOR2X1_LOC_691/B NOR2X1_LOC
XNAND2X1_LOC_400 NAND2X1_LOC_400/a_36_24# INVX1_LOC_165/A VSS VDD NOR2X1_LOC_393/Y
+ NOR2X1_LOC_394/Y NAND2X1_LOC
XNAND2X1_LOC_411 NAND2X1_LOC_411/a_36_24# NOR2X1_LOC_461/B VSS VDD INVX1_LOC_64/Y
+ NOR2X1_LOC_410/Y NAND2X1_LOC
XNAND2X1_LOC_488 NAND2X1_LOC_488/a_36_24# NOR2X1_LOC_489/A VSS VDD INVX1_LOC_89/A
+ NOR2X1_LOC_814/A NAND2X1_LOC
XNAND2X1_LOC_499 NAND2X1_LOC_499/a_36_24# NAND2X1_LOC_500/B VSS VDD NOR2X1_LOC_495/Y
+ NOR2X1_LOC_496/Y NAND2X1_LOC
XNAND2X1_LOC_477 NAND2X1_LOC_477/a_36_24# NAND2X1_LOC_477/Y VSS VDD NAND2X1_LOC_477/A
+ NAND2X1_LOC_471/Y NAND2X1_LOC
XNAND2X1_LOC_455 NAND2X1_LOC_455/a_36_24# NAND2X1_LOC_465/A VSS VDD INVX1_LOC_56/Y
+ NAND2X1_LOC_455/B NAND2X1_LOC
XNAND2X1_LOC_444 NAND2X1_LOC_444/a_36_24# INVX1_LOC_185/A VSS VDD INVX1_LOC_183/Y
+ NAND2X1_LOC_444/B NAND2X1_LOC
XNAND2X1_LOC_433 NAND2X1_LOC_433/a_36_24# NOR2X1_LOC_435/A VSS VDD INVX1_LOC_53/A
+ NOR2X1_LOC_155/A NAND2X1_LOC
XNAND2X1_LOC_466 NAND2X1_LOC_466/a_36_24# NAND2X1_LOC_466/Y VSS VDD NAND2X1_LOC_466/A
+ NAND2X1_LOC_454/Y NAND2X1_LOC
XNAND2X1_LOC_422 NAND2X1_LOC_422/a_36_24# NOR2X1_LOC_448/A VSS VDD INVX1_LOC_11/A
+ NAND2X1_LOC_93/B NAND2X1_LOC
XNAND2X1_LOC_230 NAND2X1_LOC_230/a_36_24# NOR2X1_LOC_231/A VSS VDD INVX1_LOC_5/A INVX1_LOC_21/A
+ NAND2X1_LOC
XNAND2X1_LOC_241 NAND2X1_LOC_241/a_36_24# NAND2X1_LOC_241/Y VSS VDD NOR2X1_LOC_237/Y
+ NOR2X1_LOC_238/Y NAND2X1_LOC
XNAND2X1_LOC_252 NAND2X1_LOC_252/a_36_24# NOR2X1_LOC_483/B VSS VDD INVX1_LOC_41/A
+ INVX1_LOC_45/A NAND2X1_LOC
XNAND2X1_LOC_263 NAND2X1_LOC_263/a_36_24# INVX1_LOC_123/A VSS VDD INVX1_LOC_17/A INVX1_LOC_26/Y
+ NAND2X1_LOC
XNAND2X1_LOC_296 NAND2X1_LOC_296/a_36_24# NOR2X1_LOC_297/A VSS VDD INVX1_LOC_32/A
+ INVX1_LOC_42/A NAND2X1_LOC
XNAND2X1_LOC_285 NAND2X1_LOC_285/a_36_24# NAND2X1_LOC_286/B VSS VDD NOR2X1_LOC_281/Y
+ NOR2X1_LOC_282/Y NAND2X1_LOC
XNAND2X1_LOC_274 NAND2X1_LOC_274/a_36_24# NOR2X1_LOC_275/A VSS VDD NOR2X1_LOC_272/Y
+ NOR2X1_LOC_273/Y NAND2X1_LOC
XINVX1_LOC_129 INVX1_LOC_129/Y VSS VDD INVX1_LOC_129/A INVX1_LOC
XINVX1_LOC_118 INVX1_LOC_118/Y VSS VDD INVX1_LOC_118/A INVX1_LOC
XINVX1_LOC_107 INVX1_LOC_107/Y VSS VDD INVX1_LOC_107/A INVX1_LOC
XNOR2X1_LOC_509 NOR2X1_LOC_509/a_36_216# INVX1_LOC_212/A VSS VDD NOR2X1_LOC_509/A
+ NOR2X1_LOC_340/A NOR2X1_LOC
XNOR2X1_LOC_306 NOR2X1_LOC_306/a_36_216# INVX1_LOC_142/A VSS VDD INVX1_LOC_83/Y INVX1_LOC_18/A
+ NOR2X1_LOC
XNOR2X1_LOC_328 NOR2X1_LOC_328/a_36_216# NOR2X1_LOC_328/Y VSS VDD NOR2X1_LOC_51/A
+ INPUT_4 NOR2X1_LOC
XNOR2X1_LOC_317 NOR2X1_LOC_317/a_36_216# NOR2X1_LOC_319/B VSS VDD NOR2X1_LOC_317/A
+ NOR2X1_LOC_317/B NOR2X1_LOC
XNOR2X1_LOC_339 NOR2X1_LOC_339/a_36_216# INVX1_LOC_152/A VSS VDD NOR2X1_LOC_332/Y
+ NOR2X1_LOC_61/Y NOR2X1_LOC
XNAND2X1_LOC_818 NAND2X1_LOC_818/a_36_24# NOR2X1_LOC_820/B VSS VDD INVX1_LOC_4/A INVX1_LOC_84/A
+ NAND2X1_LOC
XNAND2X1_LOC_807 NAND2X1_LOC_807/a_36_24# NAND2X1_LOC_807/Y VSS VDD NAND2X1_LOC_807/A
+ NAND2X1_LOC_807/B NAND2X1_LOC
XNAND2X1_LOC_829 NAND2X1_LOC_829/a_36_24# NOR2X1_LOC_855/A VSS VDD INVX1_LOC_49/A
+ NOR2X1_LOC_828/Y NAND2X1_LOC
XNOR2X1_LOC_851 NOR2X1_LOC_851/a_36_216# NOR2X1_LOC_858/A VSS VDD INVX1_LOC_311/Y
+ NOR2X1_LOC_840/Y NOR2X1_LOC
XNOR2X1_LOC_840 NOR2X1_LOC_840/a_36_216# NOR2X1_LOC_840/Y VSS VDD NOR2X1_LOC_840/A
+ NOR2X1_LOC_833/Y NOR2X1_LOC
XNOR2X1_LOC_862 NOR2X1_LOC_862/a_36_216# NOR2X1_LOC_865/A VSS VDD NOR2X1_LOC_859/Y
+ NOR2X1_LOC_862/B NOR2X1_LOC
XNOR2X1_LOC_13 NOR2X1_LOC_13/a_36_216# NOR2X1_LOC_13/Y VSS VDD INVX1_LOC_12/A INVX1_LOC_10/A
+ NOR2X1_LOC
XNOR2X1_LOC_46 NOR2X1_LOC_46/a_36_216# NOR2X1_LOC_48/B VSS VDD INVX1_LOC_14/A INPUT_1
+ NOR2X1_LOC
XNOR2X1_LOC_35 NOR2X1_LOC_35/a_36_216# NOR2X1_LOC_35/Y VSS VDD NOR2X1_LOC_34/Y NOR2X1_LOC_33/Y
+ NOR2X1_LOC
XNOR2X1_LOC_24 NOR2X1_LOC_24/a_36_216# NOR2X1_LOC_24/Y VSS VDD NOR2X1_LOC_45/B INVX1_LOC_18/A
+ NOR2X1_LOC
XNOR2X1_LOC_57 NOR2X1_LOC_57/a_36_216# INVX1_LOC_44/A VSS VDD INVX1_LOC_34/A INVX1_LOC_4/A
+ NOR2X1_LOC
XNOR2X1_LOC_79 NOR2X1_LOC_79/a_36_216# NOR2X1_LOC_79/Y VSS VDD NOR2X1_LOC_79/A INVX1_LOC_16/A
+ NOR2X1_LOC
XNOR2X1_LOC_68 NOR2X1_LOC_68/a_36_216# NOR2X1_LOC_68/Y VSS VDD NOR2X1_LOC_68/A INVX1_LOC_4/Y
+ NOR2X1_LOC
XNOR2X1_LOC_147 NOR2X1_LOC_147/a_36_216# INVX1_LOC_86/A VSS VDD NOR2X1_LOC_147/A NOR2X1_LOC_147/B
+ NOR2X1_LOC
XNOR2X1_LOC_158 NOR2X1_LOC_158/a_36_216# NOR2X1_LOC_158/Y VSS VDD INVX1_LOC_90/A NOR2X1_LOC_158/B
+ NOR2X1_LOC
XNOR2X1_LOC_125 NOR2X1_LOC_125/a_36_216# NOR2X1_LOC_125/Y VSS VDD INVX1_LOC_64/A INVX1_LOC_58/A
+ NOR2X1_LOC
XNOR2X1_LOC_136 NOR2X1_LOC_136/a_36_216# NOR2X1_LOC_136/Y VSS VDD INVX1_LOC_32/A INVX1_LOC_2/A
+ NOR2X1_LOC
XNOR2X1_LOC_114 NOR2X1_LOC_114/a_36_216# NOR2X1_LOC_114/Y VSS VDD NOR2X1_LOC_114/A
+ INVX1_LOC_66/Y NOR2X1_LOC
XNOR2X1_LOC_103 NOR2X1_LOC_103/a_36_216# NOR2X1_LOC_103/Y VSS VDD NOR2X1_LOC_536/A
+ INVX1_LOC_35/Y NOR2X1_LOC
XNOR2X1_LOC_169 NOR2X1_LOC_169/a_36_216# NOR2X1_LOC_170/A VSS VDD NOR2X1_LOC_703/B
+ NOR2X1_LOC_169/B NOR2X1_LOC
XNAND2X1_LOC_626 NAND2X1_LOC_626/a_36_24# NOR2X1_LOC_629/B VSS VDD INVX1_LOC_57/A
+ INVX1_LOC_91/A NAND2X1_LOC
XNAND2X1_LOC_659 NAND2X1_LOC_659/a_36_24# INVX1_LOC_267/A VSS VDD NAND2X1_LOC_659/A
+ NAND2X1_LOC_659/B NAND2X1_LOC
XNAND2X1_LOC_604 NAND2X1_LOC_604/a_36_24# NOR2X1_LOC_605/A VSS VDD INVX1_LOC_53/A
+ INVX1_LOC_91/A NAND2X1_LOC
XNAND2X1_LOC_615 NAND2X1_LOC_615/a_36_24# NOR2X1_LOC_623/B VSS VDD INVX1_LOC_18/Y
+ NOR2X1_LOC_614/Y NAND2X1_LOC
XNAND2X1_LOC_648 NAND2X1_LOC_648/a_36_24# NAND2X1_LOC_655/A VSS VDD NAND2X1_LOC_648/A
+ INVX1_LOC_264/Y NAND2X1_LOC
XNAND2X1_LOC_637 NAND2X1_LOC_637/a_36_24# NAND2X1_LOC_637/Y VSS VDD NOR2X1_LOC_585/Y
+ NOR2X1_LOC_586/Y NAND2X1_LOC
XINVX1_LOC_38 INVX1_LOC_38/Y VSS VDD INVX1_LOC_38/A INVX1_LOC
XINVX1_LOC_16 INVX1_LOC_16/Y VSS VDD INVX1_LOC_16/A INVX1_LOC
XINVX1_LOC_27 INVX1_LOC_27/Y VSS VDD INVX1_LOC_27/A INVX1_LOC
XINVX1_LOC_49 INVX1_LOC_49/Y VSS VDD INVX1_LOC_49/A INVX1_LOC
XINVX1_LOC_290 INVX1_LOC_290/Y VSS VDD INVX1_LOC_290/A INVX1_LOC
XNOR2X1_LOC_681 NOR2X1_LOC_681/a_36_216# NOR2X1_LOC_681/Y VSS VDD NOR2X1_LOC_433/A
+ INVX1_LOC_21/Y NOR2X1_LOC
XNAND2X1_LOC_90 NAND2X1_LOC_90/a_36_24# NOR2X1_LOC_383/B VSS VDD INVX1_LOC_25/A INVX1_LOC_39/A
+ NAND2X1_LOC
XNOR2X1_LOC_670 NOR2X1_LOC_670/a_36_216# NOR2X1_LOC_670/Y VSS VDD NOR2X1_LOC_536/A
+ INVX1_LOC_30/A NOR2X1_LOC
XNOR2X1_LOC_692 NOR2X1_LOC_692/a_36_216# NOR2X1_LOC_692/Y VSS VDD NOR2X1_LOC_48/B
+ INVX1_LOC_16/A NOR2X1_LOC
XNAND2X1_LOC_412 NAND2X1_LOC_412/a_36_24# NOR2X1_LOC_634/A VSS VDD INVX1_LOC_26/Y
+ INVX1_LOC_33/A NAND2X1_LOC
XNAND2X1_LOC_445 NAND2X1_LOC_445/a_36_24# NAND2X1_LOC_455/B VSS VDD NOR2X1_LOC_237/Y
+ NOR2X1_LOC_315/Y NAND2X1_LOC
XNAND2X1_LOC_401 NAND2X1_LOC_401/a_36_24# NAND2X1_LOC_402/B VSS VDD NOR2X1_LOC_395/Y
+ NOR2X1_LOC_396/Y NAND2X1_LOC
XNAND2X1_LOC_434 NAND2X1_LOC_434/a_36_24# NAND2X1_LOC_434/Y VSS VDD NOR2X1_LOC_172/Y
+ NOR2X1_LOC_431/Y NAND2X1_LOC
XNAND2X1_LOC_423 NAND2X1_LOC_423/a_36_24# NOR2X1_LOC_592/B VSS VDD INVX1_LOC_5/A INVX1_LOC_49/A
+ NAND2X1_LOC
XNAND2X1_LOC_489 NAND2X1_LOC_489/a_36_24# NAND2X1_LOC_489/Y VSS VDD NOR2X1_LOC_487/Y
+ NOR2X1_LOC_488/Y NAND2X1_LOC
XNAND2X1_LOC_478 NAND2X1_LOC_478/a_36_24# INVX1_LOC_203/A VSS VDD INVX1_LOC_200/Y
+ NAND2X1_LOC_477/Y NAND2X1_LOC
XNAND2X1_LOC_456 NAND2X1_LOC_456/a_36_24# NAND2X1_LOC_456/Y VSS VDD INVX1_LOC_100/A
+ NAND2X1_LOC_254/Y NAND2X1_LOC
XNAND2X1_LOC_467 NAND2X1_LOC_467/a_36_24# NAND2X1_LOC_470/B VSS VDD NOR2X1_LOC_163/Y
+ NAND2X1_LOC_452/Y NAND2X1_LOC
XNAND2X1_LOC_275 NAND2X1_LOC_275/a_36_24# INVX1_LOC_129/A VSS VDD D_INPUT_0 NOR2X1_LOC_274/Y
+ NAND2X1_LOC
XNAND2X1_LOC_242 NAND2X1_LOC_242/a_36_24# NAND2X1_LOC_244/A VSS VDD INVX1_LOC_119/Y
+ NAND2X1_LOC_241/Y NAND2X1_LOC
XNAND2X1_LOC_264 NAND2X1_LOC_264/a_36_24# NOR2X1_LOC_667/A VSS VDD INVX1_LOC_10/A
+ NOR2X1_LOC_89/A NAND2X1_LOC
XNAND2X1_LOC_286 NAND2X1_LOC_286/a_36_24# NAND2X1_LOC_288/A VSS VDD INVX1_LOC_131/Y
+ NAND2X1_LOC_286/B NAND2X1_LOC
XNAND2X1_LOC_253 NAND2X1_LOC_253/a_36_24# NOR2X1_LOC_254/A VSS VDD INVX1_LOC_49/A
+ INVX1_LOC_77/A NAND2X1_LOC
XNAND2X1_LOC_231 NAND2X1_LOC_231/a_36_24# NAND2X1_LOC_231/Y VSS VDD NOR2X1_LOC_229/Y
+ NOR2X1_LOC_230/Y NAND2X1_LOC
XNAND2X1_LOC_220 NAND2X1_LOC_220/a_36_24# INVX1_LOC_115/A VSS VDD NAND2X1_LOC_212/Y
+ NAND2X1_LOC_220/B NAND2X1_LOC
XNAND2X1_LOC_297 NAND2X1_LOC_297/a_36_24# INVX1_LOC_137/A VSS VDD INVX1_LOC_34/Y NOR2X1_LOC_296/Y
+ NAND2X1_LOC
XINVX1_LOC_108 INVX1_LOC_108/Y VSS VDD INVX1_LOC_108/A INVX1_LOC
XINVX1_LOC_119 INVX1_LOC_119/Y VSS VDD INVX1_LOC_119/A INVX1_LOC
XNOR2X1_LOC_307 NOR2X1_LOC_307/a_36_216# NOR2X1_LOC_307/Y VSS VDD NOR2X1_LOC_307/A
+ NOR2X1_LOC_307/B NOR2X1_LOC
XNOR2X1_LOC_329 NOR2X1_LOC_329/a_36_216# NOR2X1_LOC_329/Y VSS VDD NOR2X1_LOC_328/Y
+ NOR2X1_LOC_329/B NOR2X1_LOC
XNOR2X1_LOC_318 NOR2X1_LOC_318/a_36_216# INVX1_LOC_144/A VSS VDD NOR2X1_LOC_318/A
+ NOR2X1_LOC_318/B NOR2X1_LOC
XNAND2X1_LOC_819 NAND2X1_LOC_819/a_36_24# NAND2X1_LOC_819/Y VSS VDD INVX1_LOC_35/A
+ INVX1_LOC_40/A NAND2X1_LOC
XNAND2X1_LOC_808 NAND2X1_LOC_808/a_36_24# NAND2X1_LOC_811/B VSS VDD NAND2X1_LOC_808/A
+ NAND2X1_LOC_804/Y NAND2X1_LOC
XNOR2X1_LOC_830 NOR2X1_LOC_830/a_36_216# NOR2X1_LOC_830/Y VSS VDD NOR2X1_LOC_147/B
+ INVX1_LOC_65/A NOR2X1_LOC
XNOR2X1_LOC_841 NOR2X1_LOC_841/a_36_216# INVX1_LOC_312/A VSS VDD NOR2X1_LOC_841/A
+ NOR2X1_LOC_831/Y NOR2X1_LOC
XNOR2X1_LOC_863 NOR2X1_LOC_863/a_36_216# NOR2X1_LOC_863/Y VSS VDD NOR2X1_LOC_863/A
+ NOR2X1_LOC_863/B NOR2X1_LOC
XNOR2X1_LOC_852 NOR2X1_LOC_852/a_36_216# NOR2X1_LOC_852/Y VSS VDD NOR2X1_LOC_852/A
+ NOR2X1_LOC_852/B NOR2X1_LOC
XNOR2X1_LOC_36 NOR2X1_LOC_36/a_36_216# INVX1_LOC_24/A VSS VDD NOR2X1_LOC_36/A NOR2X1_LOC_36/B
+ NOR2X1_LOC
XNOR2X1_LOC_25 NOR2X1_LOC_25/a_36_216# NOR2X1_LOC_25/Y VSS VDD INPUT_7 D_INPUT_6
+ NOR2X1_LOC
XNOR2X1_LOC_47 NOR2X1_LOC_47/a_36_216# INVX1_LOC_36/A VSS VDD NOR2X1_LOC_30/Y NOR2X1_LOC_25/Y
+ NOR2X1_LOC
XNOR2X1_LOC_69 NOR2X1_LOC_69/a_36_216# INVX1_LOC_52/A VSS VDD NOR2X1_LOC_69/A INVX1_LOC_24/A
+ NOR2X1_LOC
XNOR2X1_LOC_58 NOR2X1_LOC_58/a_36_216# NOR2X1_LOC_58/Y VSS VDD NOR2X1_LOC_52/B INVX1_LOC_18/A
+ NOR2X1_LOC
XNOR2X1_LOC_14 NOR2X1_LOC_14/a_36_216# INVX1_LOC_14/A VSS VDD INPUT_3 INPUT_2
+ NOR2X1_LOC
XNOR2X1_LOC_148 NOR2X1_LOC_148/a_36_216# NOR2X1_LOC_148/Y VSS VDD NOR2X1_LOC_148/A
+ NOR2X1_LOC_148/B NOR2X1_LOC
XNOR2X1_LOC_137 NOR2X1_LOC_137/a_36_216# NOR2X1_LOC_137/Y VSS VDD NOR2X1_LOC_137/A
+ NOR2X1_LOC_137/B NOR2X1_LOC
XNOR2X1_LOC_115 NOR2X1_LOC_115/a_36_216# INVX1_LOC_68/A VSS VDD NOR2X1_LOC_112/Y NOR2X1_LOC_554/B
+ NOR2X1_LOC
XNOR2X1_LOC_104 NOR2X1_LOC_104/a_36_216# INVX1_LOC_64/A VSS VDD INVX1_LOC_8/A NOR2X1_LOC_6/B
+ NOR2X1_LOC
XNOR2X1_LOC_126 NOR2X1_LOC_126/a_36_216# INVX1_LOC_76/A VSS VDD INVX1_LOC_26/A NOR2X1_LOC_6/B
+ NOR2X1_LOC
XNOR2X1_LOC_159 NOR2X1_LOC_159/a_36_216# INVX1_LOC_92/A VSS VDD NOR2X1_LOC_9/Y INVX1_LOC_4/A
+ NOR2X1_LOC
XNAND2X1_LOC_616 NAND2X1_LOC_616/a_36_24# NOR2X1_LOC_621/B VSS VDD INVX1_LOC_15/A
+ INVX1_LOC_63/A NAND2X1_LOC
XNAND2X1_LOC_627 NAND2X1_LOC_627/a_36_24# NOR2X1_LOC_629/A VSS VDD INVX1_LOC_5/A INVX1_LOC_23/A
+ NAND2X1_LOC
XNAND2X1_LOC_605 NAND2X1_LOC_605/a_36_24# INVX1_LOC_249/A VSS VDD NOR2X1_LOC_603/Y
+ NOR2X1_LOC_604/Y NAND2X1_LOC
XINVX1_LOC_280 INVX1_LOC_280/Y VSS VDD INVX1_LOC_280/A INVX1_LOC
XINVX1_LOC_291 INVX1_LOC_291/Y VSS VDD INVX1_LOC_291/A INVX1_LOC
XNAND2X1_LOC_80 NAND2X1_LOC_80/a_36_24# NAND2X1_LOC_81/B VSS VDD INVX1_LOC_3/A NOR2X1_LOC_38/B
+ NAND2X1_LOC
XNAND2X1_LOC_91 NAND2X1_LOC_91/a_36_24# NOR2X1_LOC_97/A VSS VDD INVX1_LOC_37/A NOR2X1_LOC_383/B
+ NAND2X1_LOC
XNAND2X1_LOC_649 NAND2X1_LOC_649/a_36_24# NAND2X1_LOC_655/B VSS VDD NAND2X1_LOC_642/Y
+ NAND2X1_LOC_649/B NAND2X1_LOC
XNAND2X1_LOC_638 NAND2X1_LOC_638/a_36_24# NAND2X1_LOC_638/Y VSS VDD INVX1_LOC_243/Y
+ NAND2X1_LOC_637/Y NAND2X1_LOC
XINVX1_LOC_39 INVX1_LOC_39/Y VSS VDD INVX1_LOC_39/A INVX1_LOC
XINVX1_LOC_17 INVX1_LOC_17/Y VSS VDD INVX1_LOC_17/A INVX1_LOC
XINVX1_LOC_28 INVX1_LOC_28/Y VSS VDD INVX1_LOC_28/A INVX1_LOC
XNOR2X1_LOC_682 NOR2X1_LOC_682/a_36_216# NOR2X1_LOC_682/Y VSS VDD INVX1_LOC_92/A INVX1_LOC_24/A
+ NOR2X1_LOC
XNOR2X1_LOC_660 NOR2X1_LOC_660/a_36_216# NOR2X1_LOC_660/Y VSS VDD NOR2X1_LOC_656/Y
+ NOR2X1_LOC_655/Y NOR2X1_LOC
XNOR2X1_LOC_671 NOR2X1_LOC_671/a_36_216# NOR2X1_LOC_671/Y VSS VDD NOR2X1_LOC_6/B D_INPUT_2
+ NOR2X1_LOC
XNOR2X1_LOC_693 NOR2X1_LOC_693/a_36_216# NOR2X1_LOC_693/Y VSS VDD INVX1_LOC_23/Y INVX1_LOC_13/Y
+ NOR2X1_LOC
XNAND2X1_LOC_457 NAND2X1_LOC_457/a_36_24# NAND2X1_LOC_464/A VSS VDD NOR2X1_LOC_368/Y
+ NAND2X1_LOC_787/A NAND2X1_LOC
XNAND2X1_LOC_413 NAND2X1_LOC_413/a_36_24# NOR2X1_LOC_461/A VSS VDD INPUT_0 NOR2X1_LOC_634/A
+ NAND2X1_LOC
XNAND2X1_LOC_402 NAND2X1_LOC_402/a_36_24# INVX1_LOC_167/A VSS VDD INVX1_LOC_163/Y
+ NAND2X1_LOC_402/B NAND2X1_LOC
XNAND2X1_LOC_424 NAND2X1_LOC_424/a_36_24# NOR2X1_LOC_449/A VSS VDD INVX1_LOC_33/A
+ NOR2X1_LOC_78/A NAND2X1_LOC
XNAND2X1_LOC_468 NAND2X1_LOC_468/a_36_24# NAND2X1_LOC_469/B VSS VDD NAND2X1_LOC_798/B
+ NAND2X1_LOC_468/B NAND2X1_LOC
XNAND2X1_LOC_446 NAND2X1_LOC_446/a_36_24# INVX1_LOC_187/A VSS VDD INVX1_LOC_178/A
+ NOR2X1_LOC_418/Y NAND2X1_LOC
XNAND2X1_LOC_435 NAND2X1_LOC_435/a_36_24# INVX1_LOC_179/A VSS VDD NOR2X1_LOC_432/Y
+ NOR2X1_LOC_433/Y NAND2X1_LOC
XNAND2X1_LOC_479 NAND2X1_LOC_479/a_36_24# NAND2X1_LOC_479/Y VSS VDD NAND2X1_LOC_475/Y
+ NAND2X1_LOC_476/Y NAND2X1_LOC
XNOR2X1_LOC_490 NOR2X1_LOC_490/a_36_216# NOR2X1_LOC_490/Y VSS VDD NOR2X1_LOC_86/A
+ NOR2X1_LOC_19/B NOR2X1_LOC
XNAND2X1_LOC_221 NAND2X1_LOC_221/a_36_24# NAND2X1_LOC_223/A VSS VDD INVX1_LOC_104/Y
+ INVX1_LOC_116/Y NAND2X1_LOC
XNAND2X1_LOC_265 NAND2X1_LOC_265/a_36_24# INVX1_LOC_125/A VSS VDD INVX1_LOC_30/Y NOR2X1_LOC_264/Y
+ NAND2X1_LOC
XNAND2X1_LOC_254 NAND2X1_LOC_254/a_36_24# NAND2X1_LOC_254/Y VSS VDD NOR2X1_LOC_252/Y
+ NOR2X1_LOC_253/Y NAND2X1_LOC
XNAND2X1_LOC_276 NAND2X1_LOC_276/a_36_24# NAND2X1_LOC_276/Y VSS VDD NOR2X1_LOC_271/Y
+ INVX1_LOC_129/Y NAND2X1_LOC
XNAND2X1_LOC_243 NAND2X1_LOC_243/a_36_24# NAND2X1_LOC_243/Y VSS VDD NOR2X1_LOC_235/Y
+ NAND2X1_LOC_243/B NAND2X1_LOC
XNAND2X1_LOC_232 NAND2X1_LOC_232/a_36_24# NOR2X1_LOC_240/B VSS VDD NOR2X1_LOC_78/B
+ INVX1_LOC_89/A NAND2X1_LOC
XNAND2X1_LOC_287 NAND2X1_LOC_287/a_36_24# NAND2X1_LOC_288/B VSS VDD NOR2X1_LOC_278/Y
+ NAND2X1_LOC_287/B NAND2X1_LOC
XNAND2X1_LOC_298 NAND2X1_LOC_298/a_36_24# NOR2X1_LOC_302/B VSS VDD INVX1_LOC_21/A
+ INVX1_LOC_41/A NAND2X1_LOC
XNAND2X1_LOC_210 NAND2X1_LOC_210/a_36_24# INVX1_LOC_113/A VSS VDD NOR2X1_LOC_158/Y
+ NOR2X1_LOC_163/Y NAND2X1_LOC
XINVX1_LOC_109 INVX1_LOC_109/Y VSS VDD INVX1_LOC_109/A INVX1_LOC
XNOR2X1_LOC_308 NOR2X1_LOC_308/a_36_216# NOR2X1_LOC_727/B VSS VDD NOR2X1_LOC_307/Y
+ INVX1_LOC_142/Y NOR2X1_LOC
XNOR2X1_LOC_319 NOR2X1_LOC_319/a_36_216# NOR2X1_LOC_354/B VSS VDD INVX1_LOC_143/Y
+ NOR2X1_LOC_319/B NOR2X1_LOC
XNAND2X1_LOC_809 NAND2X1_LOC_809/a_36_24# NAND2X1_LOC_810/B VSS VDD NAND2X1_LOC_809/A
+ NAND2X1_LOC_802/Y NAND2X1_LOC
XNOR2X1_LOC_842 NOR2X1_LOC_842/a_36_216# NOR2X1_LOC_850/B VSS VDD NOR2X1_LOC_830/Y
+ INVX1_LOC_99/A NOR2X1_LOC
XNOR2X1_LOC_831 NOR2X1_LOC_831/a_36_216# NOR2X1_LOC_831/Y VSS VDD NOR2X1_LOC_301/A
+ NOR2X1_LOC_831/B NOR2X1_LOC
XNOR2X1_LOC_853 NOR2X1_LOC_853/a_36_216# NOR2X1_LOC_857/A VSS VDD NOR2X1_LOC_211/A
+ NOR2X1_LOC_35/Y NOR2X1_LOC
XNOR2X1_LOC_864 NOR2X1_LOC_864/a_36_216# NOR2X1_LOC_866/B VSS VDD NOR2X1_LOC_863/Y
+ INVX1_LOC_299/Y NOR2X1_LOC
XNOR2X1_LOC_820 NOR2X1_LOC_820/a_36_216# NOR2X1_LOC_820/Y VSS VDD NOR2X1_LOC_820/A
+ NOR2X1_LOC_820/B NOR2X1_LOC
XNOR2X1_LOC_48 NOR2X1_LOC_48/a_36_216# NOR2X1_LOC_48/Y VSS VDD INVX1_LOC_36/A NOR2X1_LOC_48/B
+ NOR2X1_LOC
XNOR2X1_LOC_59 NOR2X1_LOC_59/a_36_216# INVX1_LOC_46/A VSS VDD NOR2X1_LOC_25/Y NOR2X1_LOC_11/Y
+ NOR2X1_LOC
XNOR2X1_LOC_26 NOR2X1_LOC_26/a_36_216# INVX1_LOC_20/A VSS VDD NOR2X1_LOC_25/Y NOR2X1_LOC_36/A
+ NOR2X1_LOC
XNOR2X1_LOC_15 NOR2X1_LOC_15/a_36_216# NOR2X1_LOC_15/Y VSS VDD INVX1_LOC_14/A NOR2X1_LOC_9/Y
+ NOR2X1_LOC
XNOR2X1_LOC_37 NOR2X1_LOC_37/a_36_216# INVX1_LOC_26/A VSS VDD D_INPUT_3 D_INPUT_2
+ NOR2X1_LOC
XNOR2X1_LOC_149 NOR2X1_LOC_149/a_36_216# NOR2X1_LOC_209/B VSS VDD NOR2X1_LOC_148/Y
+ INVX1_LOC_85/Y NOR2X1_LOC
XNOR2X1_LOC_127 NOR2X1_LOC_127/a_36_216# NOR2X1_LOC_127/Y VSS VDD INVX1_LOC_76/A INVX1_LOC_2/A
+ NOR2X1_LOC
XNOR2X1_LOC_116 NOR2X1_LOC_116/a_36_216# NOR2X1_LOC_473/B VSS VDD INVX1_LOC_67/Y NOR2X1_LOC_114/Y
+ NOR2X1_LOC
XNOR2X1_LOC_105 NOR2X1_LOC_105/a_36_216# NOR2X1_LOC_105/Y VSS VDD INVX1_LOC_63/A NOR2X1_LOC_78/A
+ NOR2X1_LOC
XNOR2X1_LOC_138 NOR2X1_LOC_138/a_36_216# INVX1_LOC_80/A VSS VDD NOR2X1_LOC_514/A NOR2X1_LOC_332/A
+ NOR2X1_LOC
XNAND2X1_LOC_617 NAND2X1_LOC_617/a_36_24# NOR2X1_LOC_621/A VSS VDD INVX1_LOC_27/A
+ INVX1_LOC_37/A NAND2X1_LOC
XNAND2X1_LOC_606 NAND2X1_LOC_606/a_36_24# NOR2X1_LOC_607/A VSS VDD NOR2X1_LOC_536/A
+ INVX1_LOC_72/A NAND2X1_LOC
XNAND2X1_LOC_639 NAND2X1_LOC_639/a_36_24# NAND2X1_LOC_651/B VSS VDD NAND2X1_LOC_639/A
+ INVX1_LOC_262/Y NAND2X1_LOC
XNAND2X1_LOC_628 NAND2X1_LOC_628/a_36_24# INVX1_LOC_257/A VSS VDD INVX1_LOC_35/A NAND2X1_LOC_93/B
+ NAND2X1_LOC
XINVX1_LOC_18 INVX1_LOC_18/Y VSS VDD INVX1_LOC_18/A INVX1_LOC
XINVX1_LOC_270 INVX1_LOC_270/Y VSS VDD INVX1_LOC_270/A INVX1_LOC
XINVX1_LOC_292 INVX1_LOC_292/Y VSS VDD INVX1_LOC_292/A INVX1_LOC
XINVX1_LOC_29 INVX1_LOC_29/Y VSS VDD INVX1_LOC_29/A INVX1_LOC
XINVX1_LOC_281 INVX1_LOC_281/Y VSS VDD INVX1_LOC_281/A INVX1_LOC
XNAND2X1_LOC_92 NAND2X1_LOC_92/a_36_24# NAND2X1_LOC_93/B VSS VDD INPUT_1 INVX1_LOC_7/A
+ NAND2X1_LOC
XNAND2X1_LOC_81 NAND2X1_LOC_81/a_36_24# NOR2X1_LOC_84/B VSS VDD INVX1_LOC_45/A NAND2X1_LOC_81/B
+ NAND2X1_LOC
XNAND2X1_LOC_70 NAND2X1_LOC_70/a_36_24# INVX1_LOC_53/A VSS VDD NAND2X1_LOC_3/B NAND2X1_LOC_51/B
+ NAND2X1_LOC
XNOR2X1_LOC_683 NOR2X1_LOC_683/a_36_216# NOR2X1_LOC_683/Y VSS VDD INVX1_LOC_18/A NOR2X1_LOC_15/Y
+ NOR2X1_LOC
XNOR2X1_LOC_694 NOR2X1_LOC_694/a_36_216# NOR2X1_LOC_694/Y VSS VDD NOR2X1_LOC_425/Y
+ INVX1_LOC_77/Y NOR2X1_LOC
XNOR2X1_LOC_650 NOR2X1_LOC_650/a_36_216# INVX1_LOC_266/A VSS VDD NOR2X1_LOC_641/Y
+ NOR2X1_LOC_640/Y NOR2X1_LOC
XNOR2X1_LOC_661 NOR2X1_LOC_661/a_36_216# NOR2X1_LOC_662/A VSS VDD NOR2X1_LOC_661/A
+ NOR2X1_LOC_653/Y NOR2X1_LOC
XNOR2X1_LOC_672 NOR2X1_LOC_672/a_36_216# NOR2X1_LOC_672/Y VSS VDD NOR2X1_LOC_671/Y
+ INVX1_LOC_90/A NOR2X1_LOC
XNAND2X1_LOC_447 NAND2X1_LOC_447/a_36_24# NAND2X1_LOC_447/Y VSS VDD NOR2X1_LOC_419/Y
+ NOR2X1_LOC_420/Y NAND2X1_LOC
XNAND2X1_LOC_458 NAND2X1_LOC_458/a_36_24# NAND2X1_LOC_464/B VSS VDD NOR2X1_LOC_372/Y
+ NAND2X1_LOC_374/Y NAND2X1_LOC
XNAND2X1_LOC_414 NAND2X1_LOC_414/a_36_24# NOR2X1_LOC_415/A VSS VDD INPUT_3 NOR2X1_LOC_19/B
+ NAND2X1_LOC
XNAND2X1_LOC_403 NAND2X1_LOC_403/a_36_24# INVX1_LOC_169/A VSS VDD NOR2X1_LOC_399/Y
+ INVX1_LOC_166/Y NAND2X1_LOC
XNAND2X1_LOC_436 NAND2X1_LOC_436/a_36_24# NAND2X1_LOC_798/B VSS VDD NAND2X1_LOC_434/Y
+ INVX1_LOC_180/Y NAND2X1_LOC
XNAND2X1_LOC_469 NAND2X1_LOC_469/a_36_24# INVX1_LOC_199/A VSS VDD INVX1_LOC_186/Y
+ NAND2X1_LOC_469/B NAND2X1_LOC
XNAND2X1_LOC_425 NAND2X1_LOC_425/a_36_24# NAND2X1_LOC_425/Y VSS VDD D_INPUT_5
+ NAND2X1_LOC_36/A NAND2X1_LOC
XNOR2X1_LOC_480 NOR2X1_LOC_480/a_36_216# D_GATE_479 VSS VDD NOR2X1_LOC_480/A INVX1_LOC_203/Y
+ NOR2X1_LOC
XNOR2X1_LOC_491 NOR2X1_LOC_491/a_36_216# NOR2X1_LOC_491/Y VSS VDD NOR2X1_LOC_536/A
+ INVX1_LOC_22/A NOR2X1_LOC
XNAND2X1_LOC_200 NAND2X1_LOC_200/a_36_24# NAND2X1_LOC_207/B VSS VDD INVX1_LOC_106/Y
+ NAND2X1_LOC_200/B NAND2X1_LOC
XNAND2X1_LOC_211 NAND2X1_LOC_211/a_36_24# NAND2X1_LOC_211/Y VSS VDD INVX1_LOC_94/Y
+ NAND2X1_LOC_175/Y NAND2X1_LOC
XNAND2X1_LOC_266 NAND2X1_LOC_266/a_36_24# NAND2X1_LOC_267/B VSS VDD NOR2X1_LOC_262/Y
+ INVX1_LOC_124/A NAND2X1_LOC
XNAND2X1_LOC_244 NAND2X1_LOC_244/a_36_24# NAND2X1_LOC_860/A VSS VDD NAND2X1_LOC_244/A
+ NAND2X1_LOC_243/Y NAND2X1_LOC
XNAND2X1_LOC_233 NAND2X1_LOC_233/a_36_24# NAND2X1_LOC_291/B VSS VDD INPUT_0 INVX1_LOC_13/A
+ NAND2X1_LOC
XNAND2X1_LOC_222 NAND2X1_LOC_222/a_36_24# NAND2X1_LOC_223/B VSS VDD NAND2X1_LOC_222/A
+ NAND2X1_LOC_222/B NAND2X1_LOC
XNAND2X1_LOC_277 NAND2X1_LOC_277/a_36_24# NOR2X1_LOC_633/A VSS VDD INVX1_LOC_26/Y
+ INVX1_LOC_35/A NAND2X1_LOC
XNAND2X1_LOC_255 NAND2X1_LOC_255/a_36_24# NOR2X1_LOC_541/B VSS VDD INVX1_LOC_26/Y
+ INVX1_LOC_89/A NAND2X1_LOC
XNAND2X1_LOC_288 NAND2X1_LOC_288/a_36_24# INVX1_LOC_133/A VSS VDD NAND2X1_LOC_288/A
+ NAND2X1_LOC_288/B NAND2X1_LOC
XNAND2X1_LOC_299 NAND2X1_LOC_299/a_36_24# NOR2X1_LOC_302/A VSS VDD INVX1_LOC_11/A
+ INVX1_LOC_71/A NAND2X1_LOC
XNOR2X1_LOC_309 NOR2X1_LOC_309/a_36_216# NOR2X1_LOC_309/Y VSS VDD NOR2X1_LOC_226/A
+ INVX1_LOC_18/A NOR2X1_LOC
XNOR2X1_LOC_810 NOR2X1_LOC_810/a_36_216# NOR2X1_LOC_810/Y VSS VDD NOR2X1_LOC_810/A
+ INVX1_LOC_299/Y NOR2X1_LOC
XNOR2X1_LOC_832 NOR2X1_LOC_832/a_36_216# NOR2X1_LOC_841/A VSS VDD NOR2X1_LOC_435/A
+ NOR2X1_LOC_592/B NOR2X1_LOC
XNOR2X1_LOC_854 NOR2X1_LOC_854/a_36_216# NOR2X1_LOC_856/B VSS VDD NOR2X1_LOC_567/B
+ NOR2X1_LOC_326/Y NOR2X1_LOC
XNOR2X1_LOC_865 NOR2X1_LOC_865/a_36_216# NOR2X1_LOC_865/Y VSS VDD NOR2X1_LOC_865/A
+ NOR2X1_LOC_861/Y NOR2X1_LOC
XNOR2X1_LOC_821 NOR2X1_LOC_821/a_36_216# NOR2X1_LOC_821/Y VSS VDD INVX1_LOC_54/A INVX1_LOC_10/A
+ NOR2X1_LOC
XNOR2X1_LOC_843 NOR2X1_LOC_843/a_36_216# INVX1_LOC_314/A VSS VDD NOR2X1_LOC_843/A
+ NOR2X1_LOC_843/B NOR2X1_LOC
XNOR2X1_LOC_27 NOR2X1_LOC_27/a_36_216# NOR2X1_LOC_27/Y VSS VDD INVX1_LOC_20/A INVX1_LOC_5/Y
+ NOR2X1_LOC
XNOR2X1_LOC_16 NOR2X1_LOC_16/a_36_216# NOR2X1_LOC_16/Y VSS VDD NOR2X1_LOC_15/Y INVX1_LOC_1/Y
+ NOR2X1_LOC
XNOR2X1_LOC_49 NOR2X1_LOC_49/a_36_216# NOR2X1_LOC_52/B VSS VDD NOR2X1_LOC_38/B INVX1_LOC_14/A
+ NOR2X1_LOC
XNOR2X1_LOC_38 NOR2X1_LOC_38/a_36_216# INVX1_LOC_28/A VSS VDD INVX1_LOC_26/A NOR2X1_LOC_38/B
+ NOR2X1_LOC
XNOR2X1_LOC_106 NOR2X1_LOC_106/a_36_216# NOR2X1_LOC_106/Y VSS VDD NOR2X1_LOC_106/A
+ INVX1_LOC_36/A NOR2X1_LOC
XNOR2X1_LOC_139 NOR2X1_LOC_139/a_36_216# NOR2X1_LOC_139/Y VSS VDD INVX1_LOC_79/Y NOR2X1_LOC_137/Y
+ NOR2X1_LOC
XNOR2X1_LOC_117 NOR2X1_LOC_117/a_36_216# NOR2X1_LOC_117/Y VSS VDD INVX1_LOC_54/A NOR2X1_LOC_65/B
+ NOR2X1_LOC
XNOR2X1_LOC_128 NOR2X1_LOC_128/a_36_216# NOR2X1_LOC_554/A VSS VDD NOR2X1_LOC_128/A
+ NOR2X1_LOC_128/B NOR2X1_LOC
XNAND2X1_LOC_607 NAND2X1_LOC_607/a_36_24# NOR2X1_LOC_646/B VSS VDD INVX1_LOC_16/Y
+ NOR2X1_LOC_606/Y NAND2X1_LOC
XNAND2X1_LOC_618 NAND2X1_LOC_618/a_36_24# NAND2X1_LOC_618/Y VSS VDD D_INPUT_3
+ NOR2X1_LOC_82/A NAND2X1_LOC
XNAND2X1_LOC_629 NAND2X1_LOC_629/a_36_24# NAND2X1_LOC_629/Y VSS VDD NOR2X1_LOC_626/Y
+ NOR2X1_LOC_627/Y NAND2X1_LOC
XINVX1_LOC_260 INVX1_LOC_260/Y VSS VDD INVX1_LOC_260/A INVX1_LOC
XINVX1_LOC_293 INVX1_LOC_293/Y VSS VDD INVX1_LOC_293/A INVX1_LOC
XINVX1_LOC_282 INVX1_LOC_282/Y VSS VDD INVX1_LOC_282/A INVX1_LOC
XINVX1_LOC_19 INVX1_LOC_19/Y VSS VDD INVX1_LOC_19/A INVX1_LOC
XINVX1_LOC_271 INVX1_LOC_271/Y VSS VDD INVX1_LOC_271/A INVX1_LOC
XNOR2X1_LOC_651 NOR2X1_LOC_651/a_36_216# NOR2X1_LOC_654/A VSS VDD NOR2X1_LOC_639/Y
+ NOR2X1_LOC_638/Y NOR2X1_LOC
XNOR2X1_LOC_640 NOR2X1_LOC_640/a_36_216# NOR2X1_LOC_640/Y VSS VDD NOR2X1_LOC_634/Y
+ NOR2X1_LOC_640/B NOR2X1_LOC
XNAND2X1_LOC_93 NAND2X1_LOC_93/a_36_24# NOR2X1_LOC_98/B VSS VDD INVX1_LOC_19/A NAND2X1_LOC_93/B
+ NAND2X1_LOC
XNAND2X1_LOC_60 NAND2X1_LOC_60/a_36_24# NOR2X1_LOC_61/A VSS VDD INVX1_LOC_27/A INVX1_LOC_45/A
+ NAND2X1_LOC
XNAND2X1_LOC_82 NAND2X1_LOC_82/a_36_24# NAND2X1_LOC_82/Y VSS VDD INVX1_LOC_13/A NOR2X1_LOC_38/B
+ NAND2X1_LOC
XNAND2X1_LOC_71 NAND2X1_LOC_71/a_36_24# NAND2X1_LOC_72/B VSS VDD INVX1_LOC_4/Y INVX1_LOC_47/A
+ NAND2X1_LOC
XNOR2X1_LOC_662 NOR2X1_LOC_662/a_36_216# NOR2X1_LOC_663/A VSS VDD NOR2X1_LOC_662/A
+ NOR2X1_LOC_660/Y NOR2X1_LOC
XNOR2X1_LOC_684 NOR2X1_LOC_684/a_36_216# NOR2X1_LOC_684/Y VSS VDD INVX1_LOC_32/A INVX1_LOC_12/A
+ NOR2X1_LOC
XNOR2X1_LOC_695 NOR2X1_LOC_695/a_36_216# NOR2X1_LOC_695/Y VSS VDD INVX1_LOC_36/A NOR2X1_LOC_45/B
+ NOR2X1_LOC
XNOR2X1_LOC_673 NOR2X1_LOC_673/a_36_216# NOR2X1_LOC_721/B VSS VDD NOR2X1_LOC_673/A
+ NOR2X1_LOC_673/B NOR2X1_LOC
XNAND2X1_LOC_404 NAND2X1_LOC_404/a_36_24# NAND2X1_LOC_573/A VSS VDD INVX1_LOC_168/Y
+ INVX1_LOC_170/Y NAND2X1_LOC
XNAND2X1_LOC_437 NAND2X1_LOC_437/a_36_24# NOR2X1_LOC_440/B VSS VDD INVX1_LOC_46/Y
+ INVX1_LOC_87/A NAND2X1_LOC
XNAND2X1_LOC_415 NAND2X1_LOC_415/a_36_24# NOR2X1_LOC_416/A VSS VDD INVX1_LOC_136/A
+ NOR2X1_LOC_414/Y NAND2X1_LOC
XNAND2X1_LOC_448 NAND2X1_LOC_448/a_36_24# NAND2X1_LOC_453/A VSS VDD NOR2X1_LOC_421/Y
+ NOR2X1_LOC_422/Y NAND2X1_LOC
XNAND2X1_LOC_459 NAND2X1_LOC_459/a_36_24# INVX1_LOC_193/A VSS VDD NOR2X1_LOC_376/Y
+ NOR2X1_LOC_378/Y NAND2X1_LOC
XNAND2X1_LOC_426 NAND2X1_LOC_426/a_36_24# NOR2X1_LOC_450/B VSS VDD INVX1_LOC_71/A
+ NAND2X1_LOC_425/Y NAND2X1_LOC
XNOR2X1_LOC_470 NOR2X1_LOC_470/a_36_216# NOR2X1_LOC_477/B VSS VDD NOR2X1_LOC_470/A
+ NOR2X1_LOC_470/B NOR2X1_LOC
XNOR2X1_LOC_481 NOR2X1_LOC_481/a_36_216# INVX1_LOC_206/A VSS VDD NOR2X1_LOC_481/A
+ INVX1_LOC_1/Y NOR2X1_LOC
XNOR2X1_LOC_492 NOR2X1_LOC_492/a_36_216# NOR2X1_LOC_492/Y VSS VDD INVX1_LOC_76/A INVX1_LOC_46/A
+ NOR2X1_LOC
XNAND2X1_LOC_234 NAND2X1_LOC_234/a_36_24# NOR2X1_LOC_240/A VSS VDD INVX1_LOC_35/A
+ NAND2X1_LOC_291/B NAND2X1_LOC
XNAND2X1_LOC_223 NAND2X1_LOC_223/a_36_24# GATE_222 VSS VDD NAND2X1_LOC_223/A NAND2X1_LOC_223/B
+ NAND2X1_LOC
XNAND2X1_LOC_201 NAND2X1_LOC_201/a_36_24# INVX1_LOC_109/A VSS VDD NAND2X1_LOC_61/Y
+ NOR2X1_LOC_65/Y NAND2X1_LOC
XNAND2X1_LOC_212 NAND2X1_LOC_212/a_36_24# NAND2X1_LOC_212/Y VSS VDD INVX1_LOC_96/Y
+ NAND2X1_LOC_211/Y NAND2X1_LOC
XNAND2X1_LOC_289 NAND2X1_LOC_289/a_36_24# NOR2X1_LOC_333/A VSS VDD INVX1_LOC_37/A
+ NOR2X1_LOC_814/A NAND2X1_LOC
XNAND2X1_LOC_267 NAND2X1_LOC_267/a_36_24# NAND2X1_LOC_572/B VSS VDD INVX1_LOC_125/Y
+ NAND2X1_LOC_267/B NAND2X1_LOC
XNAND2X1_LOC_245 NAND2X1_LOC_245/a_36_24# NOR2X1_LOC_777/B VSS VDD INVX1_LOC_19/A
+ INVX1_LOC_26/Y NAND2X1_LOC
XNAND2X1_LOC_278 NAND2X1_LOC_278/a_36_24# NOR2X1_LOC_843/A VSS VDD NOR2X1_LOC_9/Y
+ NOR2X1_LOC_633/A NAND2X1_LOC
XNAND2X1_LOC_256 NAND2X1_LOC_256/a_36_24# NOR2X1_LOC_344/A VSS VDD NOR2X1_LOC_6/B
+ NOR2X1_LOC_541/B NAND2X1_LOC
XNAND2X1_LOC_790 NAND2X1_LOC_790/a_36_24# NAND2X1_LOC_793/B VSS VDD NOR2X1_LOC_753/Y
+ NOR2X1_LOC_754/Y NAND2X1_LOC
XINVX1_LOC_1 INVX1_LOC_1/Y VSS VDD INVX1_LOC_1/A INVX1_LOC
XNOR2X1_LOC_833 NOR2X1_LOC_833/a_36_216# NOR2X1_LOC_833/Y VSS VDD NOR2X1_LOC_499/B
+ NOR2X1_LOC_833/B NOR2X1_LOC
XNOR2X1_LOC_800 NOR2X1_LOC_800/a_36_216# NOR2X1_LOC_801/A VSS VDD INVX1_LOC_292/Y
+ NOR2X1_LOC_687/Y NOR2X1_LOC
XNOR2X1_LOC_811 NOR2X1_LOC_811/a_36_216# NOR2X1_LOC_812/A VSS VDD NOR2X1_LOC_811/A
+ NOR2X1_LOC_811/B NOR2X1_LOC
XNOR2X1_LOC_844 NOR2X1_LOC_844/a_36_216# NOR2X1_LOC_844/Y VSS VDD NOR2X1_LOC_844/A
+ NOR2X1_LOC_500/B NOR2X1_LOC
XNOR2X1_LOC_822 NOR2X1_LOC_822/a_36_216# NOR2X1_LOC_822/Y VSS VDD NOR2X1_LOC_536/A
+ INVX1_LOC_50/A NOR2X1_LOC
XNOR2X1_LOC_855 NOR2X1_LOC_855/a_36_216# NOR2X1_LOC_856/A VSS VDD NOR2X1_LOC_855/A
+ NOR2X1_LOC_729/A NOR2X1_LOC
XNOR2X1_LOC_866 NOR2X1_LOC_866/a_36_216# D_GATE_865 VSS VDD NOR2X1_LOC_865/Y NOR2X1_LOC_866/B
+ NOR2X1_LOC
XNOR2X1_LOC_17 NOR2X1_LOC_17/a_36_216# NOR2X1_LOC_36/B VSS VDD D_INPUT_7 D_INPUT_6
+ NOR2X1_LOC
XNOR2X1_LOC_28 NOR2X1_LOC_28/a_36_216# NOR2X1_LOC_38/B VSS VDD D_INPUT_1 INPUT_0
+ NOR2X1_LOC
XNOR2X1_LOC_39 NOR2X1_LOC_39/a_36_216# NOR2X1_LOC_39/Y VSS VDD INVX1_LOC_27/Y INVX1_LOC_23/Y
+ NOR2X1_LOC
XNOR2X1_LOC_129 NOR2X1_LOC_129/a_36_216# NOR2X1_LOC_589/A VSS VDD INVX1_LOC_26/A NOR2X1_LOC_82/A
+ NOR2X1_LOC
XNOR2X1_LOC_107 NOR2X1_LOC_107/a_36_216# NOR2X1_LOC_107/Y VSS VDD NOR2X1_LOC_89/A
+ INVX1_LOC_50/A NOR2X1_LOC
XNOR2X1_LOC_118 NOR2X1_LOC_118/a_36_216# INVX1_LOC_70/A VSS VDD NOR2X1_LOC_89/A INVX1_LOC_54/A
+ NOR2X1_LOC
XINVX1_LOC_250 INVX1_LOC_250/Y VSS VDD INVX1_LOC_250/A INVX1_LOC
XINVX1_LOC_261 INVX1_LOC_261/Y VSS VDD INVX1_LOC_261/A INVX1_LOC
XNAND2X1_LOC_619 NAND2X1_LOC_619/a_36_24# INVX1_LOC_253/A VSS VDD INVX1_LOC_23/A NAND2X1_LOC_618/Y
+ NAND2X1_LOC
XNAND2X1_LOC_608 NAND2X1_LOC_608/a_36_24# NOR2X1_LOC_609/A VSS VDD NOR2X1_LOC_15/Y
+ NOR2X1_LOC_74/A NAND2X1_LOC
XNAND2X1_LOC_61 NAND2X1_LOC_61/a_36_24# NAND2X1_LOC_61/Y VSS VDD NOR2X1_LOC_58/Y NOR2X1_LOC_60/Y
+ NAND2X1_LOC
XNAND2X1_LOC_50 NAND2X1_LOC_50/a_36_24# NAND2X1_LOC_51/B VSS VDD D_INPUT_6 D_INPUT_7
+ NAND2X1_LOC
XINVX1_LOC_294 INVX1_LOC_294/Y VSS VDD INVX1_LOC_294/A INVX1_LOC
XINVX1_LOC_272 INVX1_LOC_272/Y VSS VDD INVX1_LOC_272/A INVX1_LOC
XINVX1_LOC_283 INVX1_LOC_283/Y VSS VDD INVX1_LOC_283/A INVX1_LOC
XNOR2X1_LOC_685 NOR2X1_LOC_685/a_36_216# NOR2X1_LOC_685/Y VSS VDD NOR2X1_LOC_685/A
+ NOR2X1_LOC_685/B NOR2X1_LOC
XNOR2X1_LOC_696 NOR2X1_LOC_696/a_36_216# NOR2X1_LOC_696/Y VSS VDD INVX1_LOC_84/A INVX1_LOC_20/A
+ NOR2X1_LOC
XNOR2X1_LOC_674 NOR2X1_LOC_674/a_36_216# NOR2X1_LOC_674/Y VSS VDD NOR2X1_LOC_329/B
+ INVX1_LOC_54/A NOR2X1_LOC
XNOR2X1_LOC_652 NOR2X1_LOC_652/a_36_216# NOR2X1_LOC_652/Y VSS VDD NOR2X1_LOC_593/Y
+ NOR2X1_LOC_440/Y NOR2X1_LOC
XNAND2X1_LOC_94 NAND2X1_LOC_94/a_36_24# NAND2X1_LOC_96/A VSS VDD INVX1_LOC_13/A INVX1_LOC_40/A
+ NAND2X1_LOC
XNAND2X1_LOC_83 NAND2X1_LOC_83/a_36_24# NOR2X1_LOC_84/A VSS VDD INVX1_LOC_19/A NAND2X1_LOC_82/Y
+ NAND2X1_LOC
XNAND2X1_LOC_72 NAND2X1_LOC_72/a_36_24# NAND2X1_LOC_72/Y VSS VDD INVX1_LOC_54/Y NAND2X1_LOC_72/B
+ NAND2X1_LOC
XNOR2X1_LOC_663 NOR2X1_LOC_663/a_36_216# D_GATE_662 VSS VDD NOR2X1_LOC_663/A INVX1_LOC_267/Y
+ NOR2X1_LOC
XNOR2X1_LOC_630 NOR2X1_LOC_630/a_36_216# INVX1_LOC_260/A VSS VDD NOR2X1_LOC_629/Y
+ INVX1_LOC_258/Y NOR2X1_LOC
XNOR2X1_LOC_641 NOR2X1_LOC_641/a_36_216# NOR2X1_LOC_641/Y VSS VDD INVX1_LOC_125/A
+ NOR2X1_LOC_641/B NOR2X1_LOC
XNAND2X1_LOC_416 NAND2X1_LOC_416/a_36_24# INVX1_LOC_175/A VSS VDD INVX1_LOC_90/Y NOR2X1_LOC_415/Y
+ NAND2X1_LOC
XNAND2X1_LOC_405 NAND2X1_LOC_405/a_36_24# NOR2X1_LOC_406/A VSS VDD NOR2X1_LOC_48/B
+ NOR2X1_LOC_329/B NAND2X1_LOC
XNAND2X1_LOC_427 NAND2X1_LOC_427/a_36_24# NOR2X1_LOC_450/A VSS VDD INVX1_LOC_53/A
+ INVX1_LOC_77/A NAND2X1_LOC
XNAND2X1_LOC_438 NAND2X1_LOC_438/a_36_24# NOR2X1_LOC_544/A VSS VDD NOR2X1_LOC_160/B
+ INVX1_LOC_53/A NAND2X1_LOC
XNAND2X1_LOC_449 NAND2X1_LOC_449/a_36_24# INVX1_LOC_189/A VSS VDD NOR2X1_LOC_423/Y
+ NOR2X1_LOC_424/Y NAND2X1_LOC
XNOR2X1_LOC_460 NOR2X1_LOC_460/a_36_216# NOR2X1_LOC_460/Y VSS VDD NOR2X1_LOC_460/A
+ NOR2X1_LOC_460/B NOR2X1_LOC
XNOR2X1_LOC_471 NOR2X1_LOC_471/a_36_216# NOR2X1_LOC_471/Y VSS VDD NOR2X1_LOC_465/Y
+ NOR2X1_LOC_464/Y NOR2X1_LOC
XNOR2X1_LOC_493 NOR2X1_LOC_493/a_36_216# NOR2X1_LOC_717/A VSS VDD NOR2X1_LOC_493/A
+ NOR2X1_LOC_493/B NOR2X1_LOC
XNOR2X1_LOC_482 NOR2X1_LOC_482/a_36_216# NOR2X1_LOC_482/Y VSS VDD INVX1_LOC_46/A INVX1_LOC_6/A
+ NOR2X1_LOC
XNAND2X1_LOC_268 NAND2X1_LOC_268/a_36_24# INVX1_LOC_127/A VSS VDD INVX1_LOC_23/A NAND2X1_LOC_93/B
+ NAND2X1_LOC
XNAND2X1_LOC_235 NAND2X1_LOC_235/a_36_24# NOR2X1_LOC_243/B VSS VDD INVX1_LOC_48/A
+ NAND2X1_LOC_85/Y NAND2X1_LOC
XNAND2X1_LOC_202 NAND2X1_LOC_202/a_36_24# NAND2X1_LOC_206/B VSS VDD NOR2X1_LOC_67/Y
+ INVX1_LOC_51/Y NAND2X1_LOC
XNAND2X1_LOC_246 NAND2X1_LOC_246/a_36_24# NOR2X1_LOC_342/B VSS VDD NAND2X1_LOC_9/Y
+ NOR2X1_LOC_777/B NAND2X1_LOC
XNAND2X1_LOC_224 NAND2X1_LOC_224/a_36_24# NOR2X1_LOC_227/B VSS VDD INVX1_LOC_21/A
+ INVX1_LOC_75/A NAND2X1_LOC
XNAND2X1_LOC_257 NAND2X1_LOC_257/a_36_24# NOR2X1_LOC_259/B VSS VDD INVX1_LOC_15/A
+ INVX1_LOC_77/A NAND2X1_LOC
XNAND2X1_LOC_213 NAND2X1_LOC_213/a_36_24# NAND2X1_LOC_220/B VSS VDD NAND2X1_LOC_213/A
+ INVX1_LOC_114/Y NAND2X1_LOC
XNAND2X1_LOC_279 NAND2X1_LOC_279/a_36_24# NOR2X1_LOC_284/B VSS VDD INVX1_LOC_33/A
+ INVX1_LOC_77/A NAND2X1_LOC
XNOR2X1_LOC_290 NOR2X1_LOC_290/a_36_216# NOR2X1_LOC_290/Y VSS VDD INVX1_LOC_20/A NOR2X1_LOC_15/Y
+ NOR2X1_LOC
XNAND2X1_LOC_780 NAND2X1_LOC_780/a_36_24# NAND2X1_LOC_780/Y VSS VDD NOR2X1_LOC_743/Y
+ NOR2X1_LOC_744/Y NAND2X1_LOC
XNAND2X1_LOC_791 NAND2X1_LOC_791/a_36_24# NAND2X1_LOC_792/B VSS VDD NOR2X1_LOC_755/Y
+ NOR2X1_LOC_757/Y NAND2X1_LOC
XINVX1_LOC_2 INVX1_LOC_2/Y VSS VDD INVX1_LOC_2/A INVX1_LOC
XNOR2X1_LOC_834 NOR2X1_LOC_834/a_36_216# NOR2X1_LOC_840/A VSS VDD NOR2X1_LOC_678/A
+ INVX1_LOC_213/A NOR2X1_LOC
XNOR2X1_LOC_801 NOR2X1_LOC_801/a_36_216# NOR2X1_LOC_809/B VSS VDD NOR2X1_LOC_801/A
+ NOR2X1_LOC_801/B NOR2X1_LOC
XNOR2X1_LOC_812 NOR2X1_LOC_812/a_36_216# D_GATE_811 VSS VDD NOR2X1_LOC_812/A NOR2X1_LOC_810/Y
+ NOR2X1_LOC
XNOR2X1_LOC_856 NOR2X1_LOC_856/a_36_216# NOR2X1_LOC_863/B VSS VDD NOR2X1_LOC_856/A
+ NOR2X1_LOC_856/B NOR2X1_LOC
XNOR2X1_LOC_845 NOR2X1_LOC_845/a_36_216# NOR2X1_LOC_849/A VSS VDD NOR2X1_LOC_845/A
+ NOR2X1_LOC_721/B NOR2X1_LOC
XNOR2X1_LOC_823 NOR2X1_LOC_823/a_36_216# NOR2X1_LOC_823/Y VSS VDD INVX1_LOC_118/A
+ INVX1_LOC_38/A NOR2X1_LOC
XNOR2X1_LOC_18 NOR2X1_LOC_18/a_36_216# INVX1_LOC_16/A VSS VDD NOR2X1_LOC_36/B NOR2X1_LOC_11/Y
+ NOR2X1_LOC
XNOR2X1_LOC_29 NOR2X1_LOC_29/a_36_216# NOR2X1_LOC_32/B VSS VDD NOR2X1_LOC_82/A INVX1_LOC_8/A
+ NOR2X1_LOC
XNOR2X1_LOC_108 NOR2X1_LOC_108/a_36_216# INVX1_LOC_66/A VSS VDD NOR2X1_LOC_536/A INVX1_LOC_46/A
+ NOR2X1_LOC
XNOR2X1_LOC_119 NOR2X1_LOC_119/a_36_216# INVX1_LOC_72/A VSS VDD INVX1_LOC_14/A D_INPUT_1
+ NOR2X1_LOC
XNAND2X1_LOC_609 NAND2X1_LOC_609/a_36_24# NOR2X1_LOC_646/A VSS VDD INVX1_LOC_46/Y
+ NOR2X1_LOC_608/Y NAND2X1_LOC
XINVX1_LOC_240 INVX1_LOC_240/Y VSS VDD INVX1_LOC_240/A INVX1_LOC
XINVX1_LOC_284 INVX1_LOC_284/Y VSS VDD INVX1_LOC_284/A INVX1_LOC
XINVX1_LOC_251 INVX1_LOC_251/Y VSS VDD INVX1_LOC_251/A INVX1_LOC
XINVX1_LOC_273 INVX1_LOC_273/Y VSS VDD INVX1_LOC_273/A INVX1_LOC
XINVX1_LOC_262 INVX1_LOC_262/Y VSS VDD INVX1_LOC_262/A INVX1_LOC
XINVX1_LOC_295 INVX1_LOC_295/Y VSS VDD INVX1_LOC_295/A INVX1_LOC
XNAND2X1_LOC_84 NAND2X1_LOC_84/a_36_24# NAND2X1_LOC_84/Y VSS VDD NOR2X1_LOC_81/Y NOR2X1_LOC_83/Y
+ NAND2X1_LOC
XNAND2X1_LOC_62 NAND2X1_LOC_62/a_36_24# INVX1_LOC_47/A VSS VDD NOR2X1_LOC_9/Y INVX1_LOC_40/A
+ NAND2X1_LOC
XNAND2X1_LOC_73 NAND2X1_LOC_73/a_36_24# NAND2X1_LOC_74/B VSS VDD NAND2X1_LOC_9/Y INVX1_LOC_25/A
+ NAND2X1_LOC
XNAND2X1_LOC_95 NAND2X1_LOC_95/a_36_24# INVX1_LOC_57/A VSS VDD NAND2X1_LOC_11/Y NAND2X1_LOC_51/B
+ NAND2X1_LOC
XNAND2X1_LOC_40 NAND2X1_LOC_40/a_36_24# INVX1_LOC_29/A VSS VDD NAND2X1_LOC_3/B NAND2X1_LOC_59/B
+ NAND2X1_LOC
XNAND2X1_LOC_51 NAND2X1_LOC_51/a_36_24# INVX1_LOC_37/A VSS VDD NAND2X1_LOC_30/Y NAND2X1_LOC_51/B
+ NAND2X1_LOC
XNOR2X1_LOC_697 NOR2X1_LOC_697/a_36_216# NOR2X1_LOC_697/Y VSS VDD INVX1_LOC_117/Y
+ INVX1_LOC_90/A NOR2X1_LOC
XNOR2X1_LOC_631 NOR2X1_LOC_631/a_36_216# NOR2X1_LOC_631/Y VSS VDD NOR2X1_LOC_631/A
+ NOR2X1_LOC_631/B NOR2X1_LOC
XNOR2X1_LOC_686 NOR2X1_LOC_686/a_36_216# INVX1_LOC_276/A VSS VDD NOR2X1_LOC_686/A
+ NOR2X1_LOC_686/B NOR2X1_LOC
XNOR2X1_LOC_653 NOR2X1_LOC_653/a_36_216# NOR2X1_LOC_653/Y VSS VDD NOR2X1_LOC_652/Y
+ NOR2X1_LOC_653/B NOR2X1_LOC
XNOR2X1_LOC_675 NOR2X1_LOC_675/a_36_216# INVX1_LOC_270/A VSS VDD NOR2X1_LOC_675/A
+ INVX1_LOC_181/Y NOR2X1_LOC
XNOR2X1_LOC_642 NOR2X1_LOC_642/a_36_216# NOR2X1_LOC_649/B VSS VDD INVX1_LOC_217/Y
+ INVX1_LOC_175/A NOR2X1_LOC
XNOR2X1_LOC_664 NOR2X1_LOC_664/a_36_216# NOR2X1_LOC_664/Y VSS VDD NOR2X1_LOC_78/A
+ NAND2X1_LOC_74/B NOR2X1_LOC
XNOR2X1_LOC_620 NOR2X1_LOC_620/a_36_216# NOR2X1_LOC_620/Y VSS VDD NOR2X1_LOC_620/A
+ NOR2X1_LOC_620/B NOR2X1_LOC
XNAND2X1_LOC_439 NAND2X1_LOC_439/a_36_24# INVX1_LOC_181/A VSS VDD NOR2X1_LOC_177/Y
+ NOR2X1_LOC_438/Y NAND2X1_LOC
XNAND2X1_LOC_406 NAND2X1_LOC_406/a_36_24# INVX1_LOC_171/A VSS VDD INVX1_LOC_58/Y NOR2X1_LOC_405/Y
+ NAND2X1_LOC
XNAND2X1_LOC_417 NAND2X1_LOC_417/a_36_24# INVX1_LOC_177/A VSS VDD INVX1_LOC_35/A NOR2X1_LOC_814/A
+ NAND2X1_LOC
XNAND2X1_LOC_428 NAND2X1_LOC_428/a_36_24# NOR2X1_LOC_635/B VSS VDD INVX1_LOC_21/A
+ INVX1_LOC_117/A NAND2X1_LOC
XNOR2X1_LOC_450 NOR2X1_LOC_450/a_36_216# INVX1_LOC_192/A VSS VDD NOR2X1_LOC_450/A
+ NOR2X1_LOC_450/B NOR2X1_LOC
XNOR2X1_LOC_483 NOR2X1_LOC_483/a_36_216# NOR2X1_LOC_631/B VSS VDD NOR2X1_LOC_833/B
+ NOR2X1_LOC_483/B NOR2X1_LOC
XNOR2X1_LOC_472 NOR2X1_LOC_472/a_36_216# NOR2X1_LOC_476/B VSS VDD INVX1_LOC_197/Y
+ INVX1_LOC_195/Y NOR2X1_LOC
XNOR2X1_LOC_494 NOR2X1_LOC_494/a_36_216# NOR2X1_LOC_494/Y VSS VDD NOR2X1_LOC_384/A
+ INVX1_LOC_12/A NOR2X1_LOC
XNOR2X1_LOC_461 NOR2X1_LOC_461/a_36_216# NOR2X1_LOC_461/Y VSS VDD NOR2X1_LOC_461/A
+ NOR2X1_LOC_461/B NOR2X1_LOC
XNAND2X1_LOC_269 NAND2X1_LOC_269/a_36_24# NOR2X1_LOC_271/B VSS VDD INVX1_LOC_118/A
+ INVX1_LOC_127/Y NAND2X1_LOC
XNAND2X1_LOC_203 NAND2X1_LOC_203/a_36_24# NAND2X1_LOC_205/A VSS VDD NOR2X1_LOC_72/Y
+ INVX1_LOC_56/Y NAND2X1_LOC
XNAND2X1_LOC_236 NAND2X1_LOC_236/a_36_24# INVX1_LOC_117/A VSS VDD INVX1_LOC_3/A NOR2X1_LOC_82/A
+ NAND2X1_LOC
XNAND2X1_LOC_258 NAND2X1_LOC_258/a_36_24# NOR2X1_LOC_259/A VSS VDD NOR2X1_LOC_78/A
+ INVX1_LOC_89/A NAND2X1_LOC
XNAND2X1_LOC_225 NAND2X1_LOC_225/a_36_24# NOR2X1_LOC_814/A VSS VDD D_INPUT_1 INVX1_LOC_3/A
+ NAND2X1_LOC
XNAND2X1_LOC_214 NAND2X1_LOC_214/a_36_24# NAND2X1_LOC_214/Y VSS VDD NAND2X1_LOC_207/Y
+ NAND2X1_LOC_214/B NAND2X1_LOC
XNAND2X1_LOC_247 NAND2X1_LOC_247/a_36_24# NOR2X1_LOC_248/A VSS VDD INVX1_LOC_6/A INVX1_LOC_10/A
+ NAND2X1_LOC
XNOR2X1_LOC_280 NOR2X1_LOC_280/a_36_216# NOR2X1_LOC_280/Y VSS VDD INVX1_LOC_118/A
+ INVX1_LOC_36/A NOR2X1_LOC
XNOR2X1_LOC_291 NOR2X1_LOC_291/a_36_216# NOR2X1_LOC_291/Y VSS VDD NOR2X1_LOC_824/A
+ INVX1_LOC_24/A NOR2X1_LOC
XNAND2X1_LOC_770 NAND2X1_LOC_770/a_36_24# NAND2X1_LOC_770/Y VSS VDD NOR2X1_LOC_765/Y
+ NOR2X1_LOC_766/Y NAND2X1_LOC
XNAND2X1_LOC_792 NAND2X1_LOC_792/a_36_24# INVX1_LOC_307/A VSS VDD NOR2X1_LOC_759/Y
+ NAND2X1_LOC_792/B NAND2X1_LOC
XNAND2X1_LOC_781 NAND2X1_LOC_781/a_36_24# NAND2X1_LOC_782/B VSS VDD NOR2X1_LOC_745/Y
+ NOR2X1_LOC_746/Y NAND2X1_LOC
XINVX1_LOC_3 INVX1_LOC_3/Y VSS VDD INVX1_LOC_3/A INVX1_LOC
XNOR2X1_LOC_802 NOR2X1_LOC_802/a_36_216# NOR2X1_LOC_809/A VSS VDD NOR2X1_LOC_802/A
+ NOR2X1_LOC_798/Y NOR2X1_LOC
XNOR2X1_LOC_857 NOR2X1_LOC_857/a_36_216# NOR2X1_LOC_863/A VSS VDD NOR2X1_LOC_857/A
+ NOR2X1_LOC_852/Y NOR2X1_LOC
XNOR2X1_LOC_846 NOR2X1_LOC_846/a_36_216# NOR2X1_LOC_846/Y VSS VDD NOR2X1_LOC_846/A
+ NOR2X1_LOC_846/B NOR2X1_LOC
XNOR2X1_LOC_813 NOR2X1_LOC_813/a_36_216# NOR2X1_LOC_813/Y VSS VDD INVX1_LOC_123/Y
+ INVX1_LOC_48/Y NOR2X1_LOC
XNOR2X1_LOC_824 NOR2X1_LOC_824/a_36_216# NOR2X1_LOC_824/Y VSS VDD NOR2X1_LOC_824/A
+ INVX1_LOC_20/A NOR2X1_LOC
XNOR2X1_LOC_835 NOR2X1_LOC_835/a_36_216# NOR2X1_LOC_839/B VSS VDD NOR2X1_LOC_835/A
+ NOR2X1_LOC_835/B NOR2X1_LOC
XNOR2X1_LOC_19 NOR2X1_LOC_19/a_36_216# NOR2X1_LOC_19/Y VSS VDD INVX1_LOC_3/Y NOR2X1_LOC_19/B
+ NOR2X1_LOC
XNOR2X1_LOC_109 NOR2X1_LOC_109/a_36_216# NOR2X1_LOC_109/Y VSS VDD NOR2X1_LOC_89/A
+ INVX1_LOC_22/A NOR2X1_LOC
XINVX1_LOC_252 INVX1_LOC_252/Y VSS VDD INVX1_LOC_252/A INVX1_LOC
XINVX1_LOC_230 INVX1_LOC_230/Y VSS VDD INVX1_LOC_230/A INVX1_LOC
XINVX1_LOC_241 INVX1_LOC_241/Y VSS VDD INVX1_LOC_241/A INVX1_LOC
XINVX1_LOC_285 INVX1_LOC_285/Y VSS VDD INVX1_LOC_285/A INVX1_LOC
XINVX1_LOC_263 INVX1_LOC_263/Y VSS VDD INVX1_LOC_263/A INVX1_LOC
XINVX1_LOC_274 INVX1_LOC_274/Y VSS VDD INVX1_LOC_274/A INVX1_LOC
XINVX1_LOC_296 INVX1_LOC_296/Y VSS VDD INVX1_LOC_296/A INVX1_LOC
XNAND2X1_LOC_63 NAND2X1_LOC_63/a_36_24# NAND2X1_LOC_63/Y VSS VDD INVX1_LOC_8/Y INVX1_LOC_47/A
+ NAND2X1_LOC
XNAND2X1_LOC_52 NAND2X1_LOC_52/a_36_24# NOR2X1_LOC_197/B VSS VDD NOR2X1_LOC_68/A INVX1_LOC_37/A
+ NAND2X1_LOC
XNAND2X1_LOC_74 NAND2X1_LOC_74/a_36_24# NOR2X1_LOC_76/B VSS VDD INVX1_LOC_21/A NAND2X1_LOC_74/B
+ NAND2X1_LOC
XNAND2X1_LOC_96 NAND2X1_LOC_96/a_36_24# NOR2X1_LOC_98/A VSS VDD NAND2X1_LOC_96/A INVX1_LOC_57/A
+ NAND2X1_LOC
XNAND2X1_LOC_85 NAND2X1_LOC_85/a_36_24# NAND2X1_LOC_85/Y VSS VDD INVX1_LOC_15/A INVX1_LOC_26/Y
+ NAND2X1_LOC
XNAND2X1_LOC_41 NAND2X1_LOC_41/a_36_24# NAND2X1_LOC_41/Y VSS VDD INVX1_LOC_9/A INVX1_LOC_29/A
+ NAND2X1_LOC
XNAND2X1_LOC_30 NAND2X1_LOC_30/a_36_24# NAND2X1_LOC_30/Y VSS VDD INPUT_4 INPUT_5
+ NAND2X1_LOC
XNOR2X1_LOC_610 NOR2X1_LOC_610/a_36_216# NOR2X1_LOC_610/Y VSS VDD INVX1_LOC_35/A INVX1_LOC_29/A
+ NOR2X1_LOC
XNOR2X1_LOC_687 NOR2X1_LOC_687/a_36_216# NOR2X1_LOC_687/Y VSS VDD INVX1_LOC_275/Y
+ NOR2X1_LOC_685/Y NOR2X1_LOC
XNOR2X1_LOC_632 NOR2X1_LOC_632/a_36_216# NOR2X1_LOC_632/Y VSS VDD NOR2X1_LOC_631/Y
+ INVX1_LOC_259/Y NOR2X1_LOC
XNOR2X1_LOC_665 NOR2X1_LOC_665/a_36_216# NOR2X1_LOC_665/Y VSS VDD NOR2X1_LOC_665/A
+ INVX1_LOC_2/A NOR2X1_LOC
XNOR2X1_LOC_698 NOR2X1_LOC_698/a_36_216# NOR2X1_LOC_698/Y VSS VDD INVX1_LOC_76/A INVX1_LOC_50/A
+ NOR2X1_LOC
XNOR2X1_LOC_676 NOR2X1_LOC_676/a_36_216# NOR2X1_LOC_676/Y VSS VDD NOR2X1_LOC_828/A
+ INVX1_LOC_78/Y NOR2X1_LOC
XNOR2X1_LOC_654 NOR2X1_LOC_654/a_36_216# NOR2X1_LOC_661/A VSS VDD NOR2X1_LOC_654/A
+ INVX1_LOC_265/Y NOR2X1_LOC
XNOR2X1_LOC_643 NOR2X1_LOC_643/a_36_216# NOR2X1_LOC_643/Y VSS VDD NOR2X1_LOC_643/A
+ NOR2X1_LOC_537/Y NOR2X1_LOC
XNOR2X1_LOC_621 NOR2X1_LOC_621/a_36_216# NOR2X1_LOC_622/A VSS VDD NOR2X1_LOC_621/A
+ NOR2X1_LOC_621/B NOR2X1_LOC
XNAND2X1_LOC_418 NAND2X1_LOC_418/a_36_24# NOR2X1_LOC_446/A VSS VDD NOR2X1_LOC_78/B
+ INVX1_LOC_37/A NAND2X1_LOC
XNAND2X1_LOC_407 NAND2X1_LOC_407/a_36_24# NOR2X1_LOC_409/B VSS VDD INVX1_LOC_42/A
+ NOR2X1_LOC_433/A NAND2X1_LOC
XNAND2X1_LOC_429 NAND2X1_LOC_429/a_36_24# NAND2X1_LOC_430/B VSS VDD D_INPUT_7
+ NAND2X1_LOC_11/Y NAND2X1_LOC
XNOR2X1_LOC_451 NOR2X1_LOC_451/a_36_216# NOR2X1_LOC_452/A VSS VDD NOR2X1_LOC_451/A
+ NOR2X1_LOC_635/B NOR2X1_LOC
XNOR2X1_LOC_440 NOR2X1_LOC_440/a_36_216# NOR2X1_LOC_440/Y VSS VDD INVX1_LOC_181/Y
+ NOR2X1_LOC_440/B NOR2X1_LOC
XNOR2X1_LOC_473 NOR2X1_LOC_473/a_36_216# INVX1_LOC_202/A VSS VDD NOR2X1_LOC_276/Y
+ NOR2X1_LOC_473/B NOR2X1_LOC
XNOR2X1_LOC_462 NOR2X1_LOC_462/a_36_216# INVX1_LOC_196/A VSS VDD NOR2X1_LOC_461/Y
+ INVX1_LOC_176/Y NOR2X1_LOC
XNOR2X1_LOC_484 NOR2X1_LOC_484/a_36_216# NOR2X1_LOC_484/Y VSS VDD INVX1_LOC_24/A INVX1_LOC_10/A
+ NOR2X1_LOC
XNOR2X1_LOC_495 NOR2X1_LOC_495/a_36_216# NOR2X1_LOC_495/Y VSS VDD INVX1_LOC_41/Y INVX1_LOC_24/A
+ NOR2X1_LOC
XNAND2X1_LOC_215 NAND2X1_LOC_215/a_36_24# NAND2X1_LOC_219/B VSS VDD NAND2X1_LOC_215/A
+ NAND2X1_LOC_206/Y NAND2X1_LOC
XNAND2X1_LOC_226 NAND2X1_LOC_226/a_36_24# NOR2X1_LOC_227/A VSS VDD INVX1_LOC_15/A
+ NOR2X1_LOC_814/A NAND2X1_LOC
XNAND2X1_LOC_248 NAND2X1_LOC_248/a_36_24# NOR2X1_LOC_342/A VSS VDD INVX1_LOC_36/Y
+ NOR2X1_LOC_247/Y NAND2X1_LOC
XNAND2X1_LOC_204 NAND2X1_LOC_204/a_36_24# INVX1_LOC_111/A VSS VDD NOR2X1_LOC_79/Y
+ NAND2X1_LOC_84/Y NAND2X1_LOC
XNAND2X1_LOC_237 NAND2X1_LOC_237/a_36_24# NOR2X1_LOC_445/B VSS VDD INVX1_LOC_19/A
+ INVX1_LOC_117/A NAND2X1_LOC
XNAND2X1_LOC_259 NAND2X1_LOC_259/a_36_24# INVX1_LOC_121/A VSS VDD NOR2X1_LOC_257/Y
+ NOR2X1_LOC_258/Y NAND2X1_LOC
XNOR2X1_LOC_270 NOR2X1_LOC_270/a_36_216# NOR2X1_LOC_270/Y VSS VDD INVX1_LOC_23/A INVX1_LOC_15/A
+ NOR2X1_LOC
XNOR2X1_LOC_281 NOR2X1_LOC_281/a_36_216# NOR2X1_LOC_281/Y VSS VDD INVX1_LOC_118/A
+ INVX1_LOC_2/A NOR2X1_LOC
XNOR2X1_LOC_292 NOR2X1_LOC_292/a_36_216# NOR2X1_LOC_292/Y VSS VDD INVX1_LOC_87/Y INVX1_LOC_29/Y
+ NOR2X1_LOC
XNAND2X1_LOC_793 NAND2X1_LOC_793/a_36_24# NAND2X1_LOC_793/Y VSS VDD INVX1_LOC_306/Y
+ NAND2X1_LOC_793/B NAND2X1_LOC
XNAND2X1_LOC_760 NAND2X1_LOC_760/a_36_24# INVX1_LOC_291/A VSS VDD INVX1_LOC_49/A NOR2X1_LOC_405/A
+ NAND2X1_LOC
XNAND2X1_LOC_771 NAND2X1_LOC_771/a_36_24# INVX1_LOC_297/A VSS VDD INVX1_LOC_296/Y
+ NAND2X1_LOC_770/Y NAND2X1_LOC
XNAND2X1_LOC_782 NAND2X1_LOC_782/a_36_24# INVX1_LOC_301/A VSS VDD INVX1_LOC_287/Y
+ NAND2X1_LOC_782/B NAND2X1_LOC
XINVX1_LOC_4 INVX1_LOC_4/Y VSS VDD INVX1_LOC_4/A INVX1_LOC
XNAND2X1_LOC_590 NAND2X1_LOC_590/a_36_24# NOR2X1_LOC_591/A VSS VDD INVX1_LOC_28/A
+ NOR2X1_LOC_536/A NAND2X1_LOC
XNOR2X1_LOC_803 NOR2X1_LOC_803/a_36_216# NOR2X1_LOC_808/B VSS VDD NOR2X1_LOC_803/A
+ NOR2X1_LOC_803/B NOR2X1_LOC
XNOR2X1_LOC_858 NOR2X1_LOC_858/a_36_216# NOR2X1_LOC_862/B VSS VDD NOR2X1_LOC_858/A
+ NOR2X1_LOC_858/B NOR2X1_LOC
XNOR2X1_LOC_814 NOR2X1_LOC_814/a_36_216# NOR2X1_LOC_814/Y VSS VDD NOR2X1_LOC_814/A
+ INVX1_LOC_63/A NOR2X1_LOC
XNOR2X1_LOC_847 NOR2X1_LOC_847/a_36_216# INVX1_LOC_316/A VSS VDD NOR2X1_LOC_847/A
+ NOR2X1_LOC_847/B NOR2X1_LOC
XNOR2X1_LOC_825 NOR2X1_LOC_825/a_36_216# NOR2X1_LOC_825/Y VSS VDD NOR2X1_LOC_94/Y
+ INVX1_LOC_34/A NOR2X1_LOC
XNOR2X1_LOC_836 NOR2X1_LOC_836/a_36_216# NOR2X1_LOC_836/Y VSS VDD NOR2X1_LOC_836/A
+ NOR2X1_LOC_836/B NOR2X1_LOC
XINVX1_LOC_253 INVX1_LOC_253/Y VSS VDD INVX1_LOC_253/A INVX1_LOC
XINVX1_LOC_242 INVX1_LOC_242/Y VSS VDD INVX1_LOC_242/A INVX1_LOC
XINVX1_LOC_286 INVX1_LOC_286/Y VSS VDD INVX1_LOC_286/A INVX1_LOC
XINVX1_LOC_297 INVX1_LOC_297/Y VSS VDD INVX1_LOC_297/A INVX1_LOC
XINVX1_LOC_220 INVX1_LOC_220/Y VSS VDD INVX1_LOC_220/A INVX1_LOC
XINVX1_LOC_264 INVX1_LOC_264/Y VSS VDD INVX1_LOC_264/A INVX1_LOC
XINVX1_LOC_231 INVX1_LOC_231/Y VSS VDD INVX1_LOC_231/A INVX1_LOC
XINVX1_LOC_275 INVX1_LOC_275/Y VSS VDD INVX1_LOC_275/A INVX1_LOC
XNOR2X1_LOC_644 NOR2X1_LOC_644/a_36_216# NOR2X1_LOC_644/Y VSS VDD NOR2X1_LOC_644/A
+ NOR2X1_LOC_644/B NOR2X1_LOC
XNOR2X1_LOC_600 NOR2X1_LOC_600/a_36_216# NOR2X1_LOC_600/Y VSS VDD INVX1_LOC_64/A INVX1_LOC_22/A
+ NOR2X1_LOC
XNOR2X1_LOC_633 NOR2X1_LOC_633/a_36_216# NOR2X1_LOC_640/B VSS VDD NOR2X1_LOC_633/A
+ INVX1_LOC_69/A NOR2X1_LOC
XNAND2X1_LOC_97 NAND2X1_LOC_97/a_36_24# NAND2X1_LOC_99/A VSS VDD NOR2X1_LOC_89/Y NOR2X1_LOC_91/Y
+ NAND2X1_LOC
XNAND2X1_LOC_75 NAND2X1_LOC_75/a_36_24# NOR2X1_LOC_76/A VSS VDD NOR2X1_LOC_160/B INVX1_LOC_45/A
+ NAND2X1_LOC
XNAND2X1_LOC_86 NAND2X1_LOC_86/a_36_24# NAND2X1_LOC_86/Y VSS VDD INPUT_0 NAND2X1_LOC_85/Y
+ NAND2X1_LOC
XNAND2X1_LOC_42 NAND2X1_LOC_42/a_36_24# INVX1_LOC_31/A VSS VDD INPUT_1 INVX1_LOC_25/A
+ NAND2X1_LOC
XNAND2X1_LOC_20 NAND2X1_LOC_20/a_36_24# NOR2X1_LOC_33/B VSS VDD INVX1_LOC_15/A NAND2X1_LOC_20/B
+ NAND2X1_LOC
XNAND2X1_LOC_53 NAND2X1_LOC_53/a_36_24# NAND2X1_LOC_53/Y VSS VDD D_INPUT_5 NAND2X1_LOC_51/B
+ NAND2X1_LOC
XNAND2X1_LOC_64 NAND2X1_LOC_64/a_36_24# INVX1_LOC_49/A VSS VDD NAND2X1_LOC_21/Y NAND2X1_LOC_51/B
+ NAND2X1_LOC
XNAND2X1_LOC_31 NAND2X1_LOC_31/a_36_24# INVX1_LOC_21/A VSS VDD NAND2X1_LOC_1/Y NAND2X1_LOC_30/Y
+ NAND2X1_LOC
XNOR2X1_LOC_611 NOR2X1_LOC_611/a_36_216# INVX1_LOC_252/A VSS VDD INVX1_LOC_40/Y INVX1_LOC_3/Y
+ NOR2X1_LOC
XNOR2X1_LOC_622 NOR2X1_LOC_622/a_36_216# NOR2X1_LOC_624/B VSS VDD NOR2X1_LOC_622/A
+ INVX1_LOC_254/Y NOR2X1_LOC
XNOR2X1_LOC_666 NOR2X1_LOC_666/a_36_216# NOR2X1_LOC_666/Y VSS VDD NOR2X1_LOC_666/A
+ INVX1_LOC_16/A NOR2X1_LOC
XNOR2X1_LOC_677 NOR2X1_LOC_677/a_36_216# NOR2X1_LOC_677/Y VSS VDD INVX1_LOC_78/A INVX1_LOC_20/A
+ NOR2X1_LOC
XNOR2X1_LOC_699 NOR2X1_LOC_699/a_36_216# NOR2X1_LOC_748/A VSS VDD INVX1_LOC_90/A INVX1_LOC_13/Y
+ NOR2X1_LOC
XNOR2X1_LOC_655 NOR2X1_LOC_655/a_36_216# NOR2X1_LOC_655/Y VSS VDD NOR2X1_LOC_649/Y
+ NOR2X1_LOC_655/B NOR2X1_LOC
XNOR2X1_LOC_688 NOR2X1_LOC_688/a_36_216# NOR2X1_LOC_688/Y VSS VDD INVX1_LOC_135/A
+ INVX1_LOC_27/A NOR2X1_LOC
XNAND2X1_LOC_419 NAND2X1_LOC_419/a_36_24# NOR2X1_LOC_447/B VSS VDD INVX1_LOC_23/A
+ INVX1_LOC_31/A NAND2X1_LOC
XNAND2X1_LOC_408 NAND2X1_LOC_408/a_36_24# INVX1_LOC_173/A VSS VDD D_INPUT_6 NAND2X1_LOC_21/Y
+ NAND2X1_LOC
XNOR2X1_LOC_463 NOR2X1_LOC_463/a_36_216# INVX1_LOC_198/A VSS VDD NOR2X1_LOC_460/Y
+ INVX1_LOC_193/Y NOR2X1_LOC
XNOR2X1_LOC_430 NOR2X1_LOC_430/a_36_216# NOR2X1_LOC_430/Y VSS VDD NOR2X1_LOC_430/A
+ INVX1_LOC_92/A NOR2X1_LOC
XNOR2X1_LOC_452 NOR2X1_LOC_452/a_36_216# NOR2X1_LOC_467/A VSS VDD NOR2X1_LOC_452/A
+ INVX1_LOC_191/Y NOR2X1_LOC
XNOR2X1_LOC_441 NOR2X1_LOC_441/a_36_216# NOR2X1_LOC_441/Y VSS VDD NOR2X1_LOC_52/B
+ INVX1_LOC_30/A NOR2X1_LOC
XNOR2X1_LOC_474 NOR2X1_LOC_474/a_36_216# NOR2X1_LOC_475/A VSS VDD NOR2X1_LOC_474/A
+ NOR2X1_LOC_392/Y NOR2X1_LOC
XNOR2X1_LOC_485 NOR2X1_LOC_485/a_36_216# NOR2X1_LOC_485/Y VSS VDD NOR2X1_LOC_536/A
+ INVX1_LOC_34/A NOR2X1_LOC
XNOR2X1_LOC_496 NOR2X1_LOC_496/a_36_216# NOR2X1_LOC_496/Y VSS VDD INVX1_LOC_42/A INVX1_LOC_16/A
+ NOR2X1_LOC
XNAND2X1_LOC_205 NAND2X1_LOC_205/a_36_24# NAND2X1_LOC_215/A VSS VDD NAND2X1_LOC_205/A
+ INVX1_LOC_112/Y NAND2X1_LOC
XNAND2X1_LOC_216 NAND2X1_LOC_216/a_36_24# NAND2X1_LOC_218/A VSS VDD NAND2X1_LOC_656/A
+ NAND2X1_LOC_473/A NAND2X1_LOC
XNAND2X1_LOC_238 NAND2X1_LOC_238/a_36_24# NOR2X1_LOC_241/A VSS VDD NOR2X1_LOC_160/B
+ INVX1_LOC_37/A NAND2X1_LOC
XNAND2X1_LOC_249 NAND2X1_LOC_249/a_36_24# NOR2X1_LOC_250/A VSS VDD NOR2X1_LOC_45/B
+ INVX1_LOC_28/A NAND2X1_LOC
XNAND2X1_LOC_227 NAND2X1_LOC_227/a_36_24# NAND2X1_LOC_227/Y VSS VDD NOR2X1_LOC_224/Y
+ NOR2X1_LOC_226/Y NAND2X1_LOC
XNOR2X1_LOC_282 NOR2X1_LOC_282/a_36_216# NOR2X1_LOC_282/Y VSS VDD INVX1_LOC_90/A NOR2X1_LOC_536/A
+ NOR2X1_LOC
XNOR2X1_LOC_260 NOR2X1_LOC_260/a_36_216# NOR2X1_LOC_260/Y VSS VDD INVX1_LOC_89/A INVX1_LOC_11/A
+ NOR2X1_LOC
XNOR2X1_LOC_293 NOR2X1_LOC_293/a_36_216# INVX1_LOC_136/A VSS VDD INVX1_LOC_3/Y D_INPUT_1
+ NOR2X1_LOC
XNOR2X1_LOC_271 NOR2X1_LOC_271/a_36_216# NOR2X1_LOC_271/Y VSS VDD NOR2X1_LOC_368/A
+ NOR2X1_LOC_271/B NOR2X1_LOC
XNAND2X1_LOC_750 NAND2X1_LOC_750/a_36_24# NOR2X1_LOC_751/A VSS VDD INVX1_LOC_92/A
+ NOR2X1_LOC_749/Y NAND2X1_LOC
XNAND2X1_LOC_772 NAND2X1_LOC_772/a_36_24# NAND2X1_LOC_773/B VSS VDD NAND2X1_LOC_489/Y
+ NAND2X1_LOC_768/Y NAND2X1_LOC
XNAND2X1_LOC_761 NAND2X1_LOC_761/a_36_24# NOR2X1_LOC_801/B VSS VDD D_INPUT_0 NOR2X1_LOC_644/A
+ NAND2X1_LOC
XNAND2X1_LOC_794 NAND2X1_LOC_794/a_36_24# NAND2X1_LOC_804/A VSS VDD NAND2X1_LOC_787/Y
+ NAND2X1_LOC_794/B NAND2X1_LOC
XNAND2X1_LOC_783 NAND2X1_LOC_783/a_36_24# NAND2X1_LOC_783/Y VSS VDD NAND2X1_LOC_783/A
+ NAND2X1_LOC_780/Y NAND2X1_LOC
XINVX1_LOC_5 INVX1_LOC_5/Y VSS VDD INVX1_LOC_5/A INVX1_LOC
C0 NOR2X1_LOC_843/A INVX1_LOC_37/A 0.05fF
C1 INVX1_LOC_30/A NAND2X1_LOC_798/B 0.15fF
C2 NAND2X1_LOC_154/Y INVX1_LOC_117/Y 0.01fF
C3 NAND2X1_LOC_705/Y INVX1_LOC_12/A 0.06fF
C4 INVX1_LOC_13/A INVX1_LOC_123/A 0.00fF
C5 NAND2X1_LOC_350/A NAND2X1_LOC_432/a_36_24# 0.00fF
C6 NAND2X1_LOC_337/B INVX1_LOC_63/A 2.22fF
C7 INPUT_3 INVX1_LOC_84/A 0.09fF
C8 INVX1_LOC_60/A NOR2X1_LOC_98/A 0.00fF
C9 INVX1_LOC_312/A NOR2X1_LOC_841/A 0.15fF
C10 NAND2X1_LOC_303/Y INVX1_LOC_12/A 0.24fF
C11 NOR2X1_LOC_65/B INVX1_LOC_270/A 0.43fF
C12 NAND2X1_LOC_361/Y NOR2X1_LOC_536/A 0.04fF
C13 NAND2X1_LOC_569/A NOR2X1_LOC_813/Y 0.04fF
C14 INVX1_LOC_58/A INVX1_LOC_23/Y 0.00fF
C15 NOR2X1_LOC_318/B NOR2X1_LOC_188/a_36_216# 0.00fF
C16 INVX1_LOC_276/A INVX1_LOC_76/A 0.10fF
C17 NOR2X1_LOC_197/A INVX1_LOC_186/Y 0.01fF
C18 INVX1_LOC_75/A NOR2X1_LOC_156/A 0.02fF
C19 INVX1_LOC_303/A NAND2X1_LOC_617/a_36_24# 0.00fF
C20 NAND2X1_LOC_16/Y INVX1_LOC_113/A -0.03fF
C21 INVX1_LOC_313/Y NOR2X1_LOC_74/A 0.47fF
C22 INVX1_LOC_25/Y NOR2X1_LOC_124/A 0.03fF
C23 NAND2X1_LOC_579/A NAND2X1_LOC_254/Y 0.03fF
C24 INVX1_LOC_35/A NOR2X1_LOC_415/Y 0.01fF
C25 NOR2X1_LOC_67/A INVX1_LOC_76/A 2.80fF
C26 INVX1_LOC_2/A INVX1_LOC_46/A 11.62fF
C27 NAND2X1_LOC_116/A INVX1_LOC_117/A 0.02fF
C28 INVX1_LOC_95/Y INVX1_LOC_56/Y 0.10fF
C29 INVX1_LOC_78/A NOR2X1_LOC_109/Y 0.07fF
C30 INVX1_LOC_26/A NOR2X1_LOC_717/A 0.01fF
C31 NAND2X1_LOC_717/Y VDD 0.17fF
C32 NAND2X1_LOC_852/Y NAND2X1_LOC_836/Y 0.05fF
C33 INVX1_LOC_101/Y INVX1_LOC_290/Y 0.04fF
C34 NAND2X1_LOC_569/A INVX1_LOC_280/A 0.00fF
C35 INVX1_LOC_16/A NOR2X1_LOC_56/Y 0.08fF
C36 NOR2X1_LOC_759/Y NOR2X1_LOC_364/A 0.02fF
C37 NOR2X1_LOC_226/A INVX1_LOC_46/A 0.17fF
C38 NOR2X1_LOC_687/Y NOR2X1_LOC_833/Y 0.07fF
C39 NAND2X1_LOC_811/Y NAND2X1_LOC_264/a_36_24# 0.01fF
C40 NOR2X1_LOC_370/a_36_216# NOR2X1_LOC_318/B 0.00fF
C41 NOR2X1_LOC_218/A NOR2X1_LOC_89/A 0.00fF
C42 INVX1_LOC_50/A NOR2X1_LOC_754/Y 0.04fF
C43 INVX1_LOC_64/Y NAND2X1_LOC_96/A 0.02fF
C44 NOR2X1_LOC_86/A NOR2X1_LOC_670/Y 0.23fF
C45 INVX1_LOC_266/Y INVX1_LOC_38/A 0.07fF
C46 INVX1_LOC_90/A INVX1_LOC_125/Y 0.04fF
C47 NOR2X1_LOC_65/B NOR2X1_LOC_109/Y 0.07fF
C48 NAND2X1_LOC_120/a_36_24# INVX1_LOC_12/A 0.01fF
C49 VDD INVX1_LOC_16/A 1.27fF
C50 NAND2X1_LOC_661/A INVX1_LOC_6/A 0.02fF
C51 INVX1_LOC_135/A NOR2X1_LOC_346/Y 0.01fF
C52 NOR2X1_LOC_667/a_36_216# INVX1_LOC_42/A 0.00fF
C53 INVX1_LOC_16/A NAND2X1_LOC_800/A 0.03fF
C54 INVX1_LOC_63/Y INVX1_LOC_117/Y 0.01fF
C55 NOR2X1_LOC_590/A NAND2X1_LOC_206/B 0.01fF
C56 INVX1_LOC_64/A INVX1_LOC_29/Y 0.02fF
C57 INVX1_LOC_208/A INVX1_LOC_281/A 0.00fF
C58 INVX1_LOC_232/A INVX1_LOC_117/A 0.01fF
C59 INVX1_LOC_224/Y INVX1_LOC_306/Y 0.42fF
C60 NAND2X1_LOC_214/B NAND2X1_LOC_215/A 0.13fF
C61 NOR2X1_LOC_78/B INVX1_LOC_118/A 0.07fF
C62 INVX1_LOC_174/A NAND2X1_LOC_628/a_36_24# 0.00fF
C63 INVX1_LOC_83/A NOR2X1_LOC_586/Y 0.06fF
C64 INVX1_LOC_75/A INVX1_LOC_96/A 0.03fF
C65 INVX1_LOC_316/Y INVX1_LOC_280/A 0.03fF
C66 NOR2X1_LOC_94/Y INVX1_LOC_316/Y 0.01fF
C67 INVX1_LOC_1/A NAND2X1_LOC_70/a_36_24# 0.01fF
C68 INVX1_LOC_36/A INVX1_LOC_42/A 0.11fF
C69 NAND2X1_LOC_198/B NAND2X1_LOC_81/B 0.11fF
C70 NOR2X1_LOC_383/Y INVX1_LOC_117/A 0.01fF
C71 INVX1_LOC_73/A NOR2X1_LOC_78/A 0.00fF
C72 NOR2X1_LOC_76/A NAND2X1_LOC_464/A 0.02fF
C73 NOR2X1_LOC_92/Y NAND2X1_LOC_99/A 0.02fF
C74 INVX1_LOC_28/A NOR2X1_LOC_56/Y 0.07fF
C75 NOR2X1_LOC_429/a_36_216# NOR2X1_LOC_11/Y 0.00fF
C76 NOR2X1_LOC_103/Y NAND2X1_LOC_477/a_36_24# 0.00fF
C77 INPUT_1 INVX1_LOC_46/A 0.03fF
C78 NAND2X1_LOC_464/Y NAND2X1_LOC_489/Y 0.01fF
C79 INVX1_LOC_75/A NOR2X1_LOC_124/A 0.03fF
C80 INVX1_LOC_30/A INVX1_LOC_47/Y 0.18fF
C81 NOR2X1_LOC_709/A NAND2X1_LOC_572/B 0.32fF
C82 NOR2X1_LOC_172/Y INVX1_LOC_19/A 0.03fF
C83 INVX1_LOC_85/A NOR2X1_LOC_66/Y 0.00fF
C84 NAND2X1_LOC_842/B NOR2X1_LOC_266/B 0.15fF
C85 NOR2X1_LOC_716/B INVX1_LOC_125/A 0.04fF
C86 NOR2X1_LOC_704/Y NOR2X1_LOC_78/A 0.01fF
C87 INVX1_LOC_28/A VDD 1.03fF
C88 NAND2X1_LOC_147/a_36_24# INVX1_LOC_84/A 0.01fF
C89 INVX1_LOC_132/A INVX1_LOC_106/A -0.01fF
C90 NAND2X1_LOC_538/Y NOR2X1_LOC_654/A 0.10fF
C91 NOR2X1_LOC_147/B INVX1_LOC_19/A 2.35fF
C92 NOR2X1_LOC_325/A NOR2X1_LOC_809/B 0.32fF
C93 NAND2X1_LOC_323/B NOR2X1_LOC_865/Y 0.01fF
C94 INVX1_LOC_92/Y NAND2X1_LOC_642/Y 0.02fF
C95 NOR2X1_LOC_392/B INVX1_LOC_19/A 0.02fF
C96 INVX1_LOC_182/Y NOR2X1_LOC_137/Y 0.02fF
C97 NOR2X1_LOC_516/B NOR2X1_LOC_862/B 0.07fF
C98 NAND2X1_LOC_323/B NOR2X1_LOC_243/B 0.02fF
C99 INVX1_LOC_77/A NOR2X1_LOC_114/Y 0.00fF
C100 INVX1_LOC_83/A INVX1_LOC_118/A 0.10fF
C101 INVX1_LOC_215/Y NOR2X1_LOC_686/a_36_216# 0.01fF
C102 NOR2X1_LOC_690/A INVX1_LOC_12/A 0.07fF
C103 NOR2X1_LOC_15/Y NOR2X1_LOC_392/Y 1.49fF
C104 INVX1_LOC_36/A INVX1_LOC_78/A 1.57fF
C105 NOR2X1_LOC_332/A NOR2X1_LOC_656/Y 0.03fF
C106 INVX1_LOC_155/Y NOR2X1_LOC_89/A 0.02fF
C107 NOR2X1_LOC_591/Y INVX1_LOC_264/A 0.15fF
C108 INVX1_LOC_119/A INVX1_LOC_49/Y 0.19fF
C109 NAND2X1_LOC_564/B NOR2X1_LOC_88/Y 0.06fF
C110 NAND2X1_LOC_466/Y INVX1_LOC_12/A 0.01fF
C111 NOR2X1_LOC_413/Y INVX1_LOC_12/A 0.21fF
C112 NOR2X1_LOC_773/Y NOR2X1_LOC_654/a_36_216# 0.00fF
C113 INVX1_LOC_17/A NOR2X1_LOC_598/B 0.15fF
C114 NOR2X1_LOC_844/A NOR2X1_LOC_340/A 0.00fF
C115 NOR2X1_LOC_718/Y INVX1_LOC_283/A 0.06fF
C116 INVX1_LOC_51/Y INVX1_LOC_176/A 0.03fF
C117 NOR2X1_LOC_194/Y INVX1_LOC_12/A 0.03fF
C118 NOR2X1_LOC_773/Y INVX1_LOC_63/A 0.14fF
C119 INVX1_LOC_58/A NOR2X1_LOC_596/Y 0.07fF
C120 INVX1_LOC_288/A INVX1_LOC_36/A 0.02fF
C121 NOR2X1_LOC_337/Y NOR2X1_LOC_35/Y 0.27fF
C122 INVX1_LOC_94/A INVX1_LOC_94/Y 0.04fF
C123 NOR2X1_LOC_309/Y INVX1_LOC_42/A 0.14fF
C124 NOR2X1_LOC_471/Y NOR2X1_LOC_598/B 0.08fF
C125 NOR2X1_LOC_65/B INVX1_LOC_36/A 0.22fF
C126 NOR2X1_LOC_441/Y INVX1_LOC_271/A 0.05fF
C127 NAND2X1_LOC_564/B INVX1_LOC_84/A 0.03fF
C128 D_INPUT_0 NAND2X1_LOC_243/B 0.08fF
C129 INVX1_LOC_25/A NAND2X1_LOC_37/a_36_24# 0.02fF
C130 NOR2X1_LOC_772/A INVX1_LOC_54/A 0.00fF
C131 NOR2X1_LOC_208/Y INVX1_LOC_78/A 0.03fF
C132 NOR2X1_LOC_456/Y NOR2X1_LOC_590/A 0.07fF
C133 INVX1_LOC_122/Y NOR2X1_LOC_843/B 0.00fF
C134 NOR2X1_LOC_71/Y INVX1_LOC_35/Y 0.00fF
C135 INVX1_LOC_124/A NOR2X1_LOC_114/Y 0.27fF
C136 NOR2X1_LOC_598/B NAND2X1_LOC_555/Y 0.03fF
C137 INVX1_LOC_85/Y INVX1_LOC_179/A 0.29fF
C138 NOR2X1_LOC_818/a_36_216# INPUT_3 0.01fF
C139 NOR2X1_LOC_643/Y NAND2X1_LOC_223/A 0.03fF
C140 NOR2X1_LOC_237/Y INVX1_LOC_78/A 0.43fF
C141 NOR2X1_LOC_657/B NAND2X1_LOC_274/a_36_24# 0.00fF
C142 NOR2X1_LOC_103/Y INVX1_LOC_306/Y 0.17fF
C143 INVX1_LOC_14/A NAND2X1_LOC_474/Y 0.03fF
C144 NOR2X1_LOC_68/A NOR2X1_LOC_383/B 0.19fF
C145 NOR2X1_LOC_242/a_36_216# NAND2X1_LOC_291/B 0.00fF
C146 INVX1_LOC_11/Y NOR2X1_LOC_305/a_36_216# 0.00fF
C147 NOR2X1_LOC_567/B NOR2X1_LOC_640/Y 0.62fF
C148 NAND2X1_LOC_26/a_36_24# NAND2X1_LOC_3/B 0.00fF
C149 NOR2X1_LOC_778/B NOR2X1_LOC_850/B 0.01fF
C150 NOR2X1_LOC_311/a_36_216# NOR2X1_LOC_111/A 0.01fF
C151 NOR2X1_LOC_65/B INVX1_LOC_145/A 0.05fF
C152 NOR2X1_LOC_373/Y NAND2X1_LOC_477/Y 0.20fF
C153 INVX1_LOC_191/A INVX1_LOC_38/A 0.39fF
C154 NOR2X1_LOC_637/Y NOR2X1_LOC_638/Y 0.01fF
C155 INVX1_LOC_161/A NOR2X1_LOC_304/Y 0.10fF
C156 NOR2X1_LOC_16/Y INVX1_LOC_32/A 0.01fF
C157 NOR2X1_LOC_332/A INVX1_LOC_63/A 0.20fF
C158 INVX1_LOC_186/A INVX1_LOC_117/A 0.11fF
C159 INPUT_6 D_INPUT_7 2.95fF
C160 NOR2X1_LOC_613/Y NAND2X1_LOC_550/A 0.03fF
C161 INVX1_LOC_25/A INVX1_LOC_24/A 0.07fF
C162 INVX1_LOC_90/A NOR2X1_LOC_653/Y 0.06fF
C163 NOR2X1_LOC_309/Y INVX1_LOC_78/A 0.11fF
C164 VDD NOR2X1_LOC_253/Y 0.35fF
C165 INVX1_LOC_41/A NAND2X1_LOC_99/A 0.01fF
C166 VDD NOR2X1_LOC_35/Y 4.78fF
C167 INVX1_LOC_191/A NOR2X1_LOC_51/A 0.04fF
C168 INVX1_LOC_45/A INVX1_LOC_306/Y 0.08fF
C169 INVX1_LOC_27/A NOR2X1_LOC_441/Y 0.03fF
C170 NAND2X1_LOC_213/A INVX1_LOC_174/A 0.49fF
C171 NAND2X1_LOC_725/Y INVX1_LOC_209/Y 0.03fF
C172 NOR2X1_LOC_496/Y NAND2X1_LOC_500/Y 0.18fF
C173 INVX1_LOC_232/A INVX1_LOC_3/Y 0.10fF
C174 NOR2X1_LOC_111/A INVX1_LOC_20/A 0.10fF
C175 INVX1_LOC_90/A INVX1_LOC_19/A 6.33fF
C176 NOR2X1_LOC_528/Y INVX1_LOC_54/A 0.10fF
C177 INVX1_LOC_91/A NOR2X1_LOC_629/Y 0.04fF
C178 NAND2X1_LOC_564/B INVX1_LOC_15/A 0.07fF
C179 INVX1_LOC_90/A NOR2X1_LOC_11/Y 0.03fF
C180 NOR2X1_LOC_65/B NOR2X1_LOC_309/Y 0.03fF
C181 NOR2X1_LOC_388/Y INVX1_LOC_57/A 0.03fF
C182 NOR2X1_LOC_389/B INVX1_LOC_19/A 0.11fF
C183 D_INPUT_0 INVX1_LOC_284/A 0.28fF
C184 NOR2X1_LOC_346/Y INVX1_LOC_280/A 0.05fF
C185 INVX1_LOC_25/A NOR2X1_LOC_557/Y 0.38fF
C186 NOR2X1_LOC_142/Y INVX1_LOC_271/A 0.10fF
C187 INVX1_LOC_58/A NOR2X1_LOC_722/a_36_216# 0.00fF
C188 NAND2X1_LOC_9/Y INVX1_LOC_49/A 0.01fF
C189 INVX1_LOC_286/A NOR2X1_LOC_216/B 0.10fF
C190 NOR2X1_LOC_694/Y INVX1_LOC_20/A 0.00fF
C191 NAND2X1_LOC_303/Y NAND2X1_LOC_733/Y 0.20fF
C192 INVX1_LOC_28/A INVX1_LOC_133/A 0.07fF
C193 NOR2X1_LOC_664/Y NAND2X1_LOC_215/A 0.01fF
C194 INVX1_LOC_103/A NOR2X1_LOC_389/A 0.10fF
C195 INVX1_LOC_281/A NAND2X1_LOC_211/Y 0.00fF
C196 INVX1_LOC_143/A INVX1_LOC_116/Y 0.00fF
C197 NOR2X1_LOC_152/Y NOR2X1_LOC_109/Y 0.01fF
C198 INVX1_LOC_256/Y INVX1_LOC_26/A 0.07fF
C199 INVX1_LOC_17/A NOR2X1_LOC_372/A 0.20fF
C200 NOR2X1_LOC_368/Y INVX1_LOC_118/A 0.02fF
C201 NOR2X1_LOC_420/a_36_216# INVX1_LOC_314/Y 0.01fF
C202 INVX1_LOC_7/Y NAND2X1_LOC_656/A 0.06fF
C203 NOR2X1_LOC_188/A NAND2X1_LOC_206/Y 0.07fF
C204 INVX1_LOC_71/A INVX1_LOC_306/Y 0.10fF
C205 INVX1_LOC_83/A INVX1_LOC_257/A 0.03fF
C206 INVX1_LOC_266/A NOR2X1_LOC_274/B 0.01fF
C207 INVX1_LOC_306/A INVX1_LOC_251/A 0.03fF
C208 NAND2X1_LOC_348/A INVX1_LOC_19/A 0.03fF
C209 NOR2X1_LOC_289/Y INVX1_LOC_272/A 0.03fF
C210 INVX1_LOC_223/A INVX1_LOC_88/A 0.10fF
C211 NAND2X1_LOC_9/Y INVX1_LOC_60/A 0.01fF
C212 NOR2X1_LOC_863/Y NOR2X1_LOC_863/A 0.00fF
C213 NAND2X1_LOC_53/Y NOR2X1_LOC_717/Y 0.10fF
C214 INVX1_LOC_269/A NOR2X1_LOC_703/B 0.01fF
C215 NOR2X1_LOC_32/B NOR2X1_LOC_52/B 0.24fF
C216 INVX1_LOC_35/A INVX1_LOC_104/A 0.04fF
C217 NOR2X1_LOC_798/A INVX1_LOC_49/A 0.03fF
C218 NAND2X1_LOC_212/Y INVX1_LOC_92/A 0.03fF
C219 INVX1_LOC_46/A INVX1_LOC_118/A 0.43fF
C220 NOR2X1_LOC_716/B NOR2X1_LOC_81/Y 0.02fF
C221 NOR2X1_LOC_815/a_36_216# NOR2X1_LOC_510/Y 0.00fF
C222 NOR2X1_LOC_639/B NOR2X1_LOC_52/B 0.04fF
C223 NOR2X1_LOC_193/a_36_216# NAND2X1_LOC_63/Y 0.00fF
C224 NAND2X1_LOC_9/Y INVX1_LOC_2/A 0.01fF
C225 INVX1_LOC_24/A INVX1_LOC_1/A 0.22fF
C226 INVX1_LOC_36/A NOR2X1_LOC_503/Y 0.00fF
C227 INVX1_LOC_64/A NOR2X1_LOC_361/Y 0.06fF
C228 INVX1_LOC_95/Y NOR2X1_LOC_179/a_36_216# 0.01fF
C229 INVX1_LOC_233/A INVX1_LOC_2/A 0.07fF
C230 INPUT_0 INVX1_LOC_106/Y 0.02fF
C231 INVX1_LOC_21/A NOR2X1_LOC_445/Y 0.00fF
C232 NAND2X1_LOC_9/Y NOR2X1_LOC_226/A 0.01fF
C233 INVX1_LOC_27/A NOR2X1_LOC_340/Y 0.02fF
C234 NOR2X1_LOC_570/Y NOR2X1_LOC_383/B 0.01fF
C235 NAND2X1_LOC_705/Y NAND2X1_LOC_787/B 0.42fF
C236 INVX1_LOC_103/A NOR2X1_LOC_596/A 0.01fF
C237 NOR2X1_LOC_197/A INVX1_LOC_18/A 0.01fF
C238 NOR2X1_LOC_231/B INVX1_LOC_30/A 0.01fF
C239 INVX1_LOC_14/Y INVX1_LOC_92/A 0.11fF
C240 INVX1_LOC_233/A NOR2X1_LOC_226/A 0.19fF
C241 NOR2X1_LOC_736/Y INVX1_LOC_4/A 0.04fF
C242 INVX1_LOC_266/A NOR2X1_LOC_577/Y 0.28fF
C243 NAND2X1_LOC_573/Y NAND2X1_LOC_833/Y 0.03fF
C244 INVX1_LOC_58/A INVX1_LOC_232/A 0.19fF
C245 NOR2X1_LOC_836/Y NOR2X1_LOC_852/A 0.00fF
C246 NOR2X1_LOC_156/Y INVX1_LOC_37/A 0.01fF
C247 NAND2X1_LOC_714/B NAND2X1_LOC_354/B 0.03fF
C248 NAND2X1_LOC_149/Y INVX1_LOC_153/Y 0.12fF
C249 INVX1_LOC_17/A NOR2X1_LOC_513/a_36_216# 0.00fF
C250 INVX1_LOC_13/A D_INPUT_1 1.50fF
C251 INVX1_LOC_24/A NOR2X1_LOC_794/B 0.03fF
C252 INVX1_LOC_1/A NOR2X1_LOC_557/Y 0.31fF
C253 NAND2X1_LOC_214/B NOR2X1_LOC_655/B 0.01fF
C254 NAND2X1_LOC_149/Y INVX1_LOC_121/Y 0.03fF
C255 INVX1_LOC_2/A NOR2X1_LOC_798/A 0.03fF
C256 NOR2X1_LOC_331/B INVX1_LOC_274/A 0.04fF
C257 INVX1_LOC_292/A NOR2X1_LOC_596/A 0.12fF
C258 INVX1_LOC_278/A NAND2X1_LOC_564/B 0.01fF
C259 NOR2X1_LOC_218/A NOR2X1_LOC_433/A 0.01fF
C260 NOR2X1_LOC_626/Y NOR2X1_LOC_627/Y 0.02fF
C261 INVX1_LOC_90/A INVX1_LOC_26/Y 0.13fF
C262 INVX1_LOC_36/A NOR2X1_LOC_554/B 0.21fF
C263 NOR2X1_LOC_226/A NOR2X1_LOC_798/A 0.03fF
C264 INVX1_LOC_135/A INVX1_LOC_57/A 0.16fF
C265 NOR2X1_LOC_454/Y NOR2X1_LOC_200/a_36_216# 0.01fF
C266 NOR2X1_LOC_274/a_36_216# NOR2X1_LOC_590/A 0.00fF
C267 NOR2X1_LOC_667/Y NOR2X1_LOC_152/a_36_216# 0.01fF
C268 NOR2X1_LOC_655/B INVX1_LOC_27/A 0.01fF
C269 NAND2X1_LOC_214/B NAND2X1_LOC_553/a_36_24# 0.01fF
C270 INVX1_LOC_57/Y NOR2X1_LOC_68/A 0.06fF
C271 INVX1_LOC_256/A NAND2X1_LOC_361/Y 0.01fF
C272 INVX1_LOC_39/A NOR2X1_LOC_78/B 0.06fF
C273 NOR2X1_LOC_172/Y INVX1_LOC_161/Y 0.02fF
C274 NOR2X1_LOC_27/Y NAND2X1_LOC_725/B 0.02fF
C275 INVX1_LOC_2/A NAND2X1_LOC_703/Y 0.30fF
C276 NOR2X1_LOC_528/Y NOR2X1_LOC_48/B 0.02fF
C277 NOR2X1_LOC_598/B NOR2X1_LOC_199/B 0.03fF
C278 INVX1_LOC_25/A NOR2X1_LOC_130/A 0.00fF
C279 D_INPUT_0 NAND2X1_LOC_275/a_36_24# 0.01fF
C280 INVX1_LOC_224/A NOR2X1_LOC_720/B 0.40fF
C281 INVX1_LOC_225/Y INVX1_LOC_33/A 0.03fF
C282 NOR2X1_LOC_381/Y NOR2X1_LOC_84/a_36_216# 0.00fF
C283 INVX1_LOC_5/A INVX1_LOC_1/Y 0.00fF
C284 INVX1_LOC_166/A INVX1_LOC_90/A 0.05fF
C285 INVX1_LOC_84/A NAND2X1_LOC_804/Y 0.11fF
C286 INVX1_LOC_123/A INVX1_LOC_32/A 0.07fF
C287 NOR2X1_LOC_590/A NOR2X1_LOC_550/B 3.74fF
C288 INVX1_LOC_144/A INVX1_LOC_94/Y 0.03fF
C289 NOR2X1_LOC_226/A NAND2X1_LOC_703/Y 0.12fF
C290 INVX1_LOC_22/A INVX1_LOC_50/Y 0.05fF
C291 NOR2X1_LOC_272/Y NOR2X1_LOC_131/Y 0.03fF
C292 NAND2X1_LOC_860/A NOR2X1_LOC_71/Y 1.11fF
C293 NOR2X1_LOC_389/A INVX1_LOC_67/A 0.03fF
C294 INVX1_LOC_64/A NAND2X1_LOC_461/a_36_24# 0.00fF
C295 NOR2X1_LOC_392/B INVX1_LOC_161/Y 0.19fF
C296 INVX1_LOC_6/A NOR2X1_LOC_89/a_36_216# 0.00fF
C297 NOR2X1_LOC_788/B INVX1_LOC_23/A 0.01fF
C298 NOR2X1_LOC_68/A NOR2X1_LOC_512/Y 0.03fF
C299 INVX1_LOC_1/A INVX1_LOC_143/A 0.08fF
C300 NOR2X1_LOC_248/a_36_216# INVX1_LOC_57/A 0.00fF
C301 INVX1_LOC_286/Y INVX1_LOC_231/Y 0.03fF
C302 INVX1_LOC_36/A NOR2X1_LOC_152/Y 0.08fF
C303 NAND2X1_LOC_455/B NOR2X1_LOC_368/Y 0.13fF
C304 D_INPUT_1 INVX1_LOC_55/Y 0.03fF
C305 INVX1_LOC_269/A NAND2X1_LOC_578/B 0.02fF
C306 NOR2X1_LOC_658/Y NOR2X1_LOC_214/a_36_216# 0.01fF
C307 NAND2X1_LOC_149/Y NAND2X1_LOC_162/A 0.06fF
C308 NAND2X1_LOC_63/Y INVX1_LOC_46/A 0.09fF
C309 NOR2X1_LOC_813/Y NOR2X1_LOC_662/A 0.18fF
C310 D_INPUT_7 NOR2X1_LOC_50/a_36_216# 0.00fF
C311 NAND2X1_LOC_468/B INVX1_LOC_290/Y 0.01fF
C312 INVX1_LOC_17/A NAND2X1_LOC_660/A 0.16fF
C313 NOR2X1_LOC_690/A NAND2X1_LOC_733/Y 0.10fF
C314 NOR2X1_LOC_401/Y NOR2X1_LOC_401/A 0.00fF
C315 NOR2X1_LOC_19/B NAND2X1_LOC_215/A 0.02fF
C316 NAND2X1_LOC_9/Y INPUT_1 0.06fF
C317 NOR2X1_LOC_272/Y NOR2X1_LOC_589/A 0.07fF
C318 INVX1_LOC_35/Y NAND2X1_LOC_243/Y 0.00fF
C319 VDD INVX1_LOC_109/A 0.00fF
C320 INVX1_LOC_233/A INPUT_1 0.36fF
C321 NOR2X1_LOC_489/A NAND2X1_LOC_572/B 0.00fF
C322 INVX1_LOC_235/Y NAND2X1_LOC_376/a_36_24# 0.00fF
C323 INVX1_LOC_255/Y NAND2X1_LOC_473/A 0.03fF
C324 NOR2X1_LOC_135/Y INVX1_LOC_23/A 0.00fF
C325 NOR2X1_LOC_474/A INVX1_LOC_195/Y 0.02fF
C326 NAND2X1_LOC_214/B NOR2X1_LOC_99/B 0.14fF
C327 NOR2X1_LOC_15/Y INVX1_LOC_25/Y 1.23fF
C328 INVX1_LOC_280/A NOR2X1_LOC_662/A 0.07fF
C329 NOR2X1_LOC_99/Y INVX1_LOC_123/Y 0.00fF
C330 NAND2X1_LOC_802/Y NAND2X1_LOC_810/B 0.02fF
C331 INVX1_LOC_266/A INVX1_LOC_22/A 0.07fF
C332 INVX1_LOC_226/Y INVX1_LOC_14/A 0.12fF
C333 NOR2X1_LOC_123/B INVX1_LOC_306/Y 0.00fF
C334 NOR2X1_LOC_246/A NOR2X1_LOC_652/Y 1.11fF
C335 NOR2X1_LOC_401/Y NOR2X1_LOC_160/B 0.01fF
C336 INVX1_LOC_38/A INVX1_LOC_19/A 0.16fF
C337 NOR2X1_LOC_361/B INVX1_LOC_16/A 0.03fF
C338 INVX1_LOC_33/A INVX1_LOC_72/Y 0.11fF
C339 NOR2X1_LOC_690/A INVX1_LOC_217/A 1.71fF
C340 NAND2X1_LOC_11/Y INVX1_LOC_174/A 0.29fF
C341 NAND2X1_LOC_553/A INPUT_1 0.03fF
C342 INVX1_LOC_27/A NOR2X1_LOC_99/B 0.17fF
C343 INVX1_LOC_38/A NOR2X1_LOC_11/Y 0.03fF
C344 GATE_741 NOR2X1_LOC_380/A 0.51fF
C345 NAND2X1_LOC_733/A NAND2X1_LOC_722/A 0.03fF
C346 NOR2X1_LOC_220/A INVX1_LOC_292/A 0.10fF
C347 NOR2X1_LOC_205/Y NOR2X1_LOC_665/A 0.03fF
C348 INVX1_LOC_41/A NAND2X1_LOC_656/A 0.02fF
C349 INVX1_LOC_27/A NOR2X1_LOC_846/B 0.01fF
C350 NAND2X1_LOC_848/A INVX1_LOC_284/A 0.03fF
C351 INVX1_LOC_37/A D_INPUT_5 0.04fF
C352 NAND2X1_LOC_337/B INVX1_LOC_1/Y 0.01fF
C353 NOR2X1_LOC_147/A INVX1_LOC_23/A 0.01fF
C354 NAND2X1_LOC_656/Y NOR2X1_LOC_359/a_36_216# 0.01fF
C355 NOR2X1_LOC_168/Y NOR2X1_LOC_337/a_36_216# 0.00fF
C356 NOR2X1_LOC_510/Y INVX1_LOC_28/A 0.42fF
C357 NOR2X1_LOC_570/B NOR2X1_LOC_303/Y 0.10fF
C358 NOR2X1_LOC_498/Y NOR2X1_LOC_484/Y 0.05fF
C359 INVX1_LOC_249/A NOR2X1_LOC_142/Y 0.52fF
C360 NOR2X1_LOC_51/A NOR2X1_LOC_11/Y 0.91fF
C361 INVX1_LOC_221/A INVX1_LOC_24/A 0.16fF
C362 INVX1_LOC_223/A NOR2X1_LOC_203/Y 0.00fF
C363 INVX1_LOC_136/A NAND2X1_LOC_342/Y 0.01fF
C364 NAND2X1_LOC_218/B NOR2X1_LOC_6/B 0.06fF
C365 INVX1_LOC_230/Y NOR2X1_LOC_789/A 0.02fF
C366 NOR2X1_LOC_791/A NAND2X1_LOC_338/B 0.01fF
C367 NOR2X1_LOC_140/A NOR2X1_LOC_130/Y 0.09fF
C368 NAND2X1_LOC_131/a_36_24# NOR2X1_LOC_130/A 0.00fF
C369 INVX1_LOC_292/A NOR2X1_LOC_548/Y 0.03fF
C370 NOR2X1_LOC_186/Y INVX1_LOC_73/A 0.03fF
C371 NAND2X1_LOC_833/Y NAND2X1_LOC_640/Y 0.38fF
C372 NOR2X1_LOC_656/Y NOR2X1_LOC_847/A 0.03fF
C373 NOR2X1_LOC_690/A NAND2X1_LOC_787/B 0.10fF
C374 NAND2X1_LOC_350/B NOR2X1_LOC_52/Y 0.07fF
C375 NOR2X1_LOC_7/Y INVX1_LOC_53/A 0.11fF
C376 NOR2X1_LOC_92/Y NOR2X1_LOC_329/B 0.14fF
C377 INVX1_LOC_35/A INVX1_LOC_86/Y 0.07fF
C378 NOR2X1_LOC_640/Y NOR2X1_LOC_633/a_36_216# 0.00fF
C379 INVX1_LOC_225/A NAND2X1_LOC_833/Y 0.12fF
C380 INVX1_LOC_227/Y NOR2X1_LOC_500/Y 0.02fF
C381 NAND2X1_LOC_565/B NOR2X1_LOC_384/Y 0.01fF
C382 NOR2X1_LOC_361/B INVX1_LOC_28/A 0.19fF
C383 INVX1_LOC_21/A NOR2X1_LOC_335/B 0.04fF
C384 NAND2X1_LOC_727/Y INVX1_LOC_72/A 0.01fF
C385 INVX1_LOC_90/A INVX1_LOC_161/Y 0.07fF
C386 INVX1_LOC_58/A NAND2X1_LOC_447/Y 0.19fF
C387 NOR2X1_LOC_716/B NOR2X1_LOC_709/A 0.28fF
C388 NOR2X1_LOC_246/A NAND2X1_LOC_805/a_36_24# 0.01fF
C389 INVX1_LOC_33/A INVX1_LOC_266/Y 2.49fF
C390 NOR2X1_LOC_52/B NOR2X1_LOC_364/Y 0.01fF
C391 NOR2X1_LOC_2/Y NOR2X1_LOC_582/A 0.00fF
C392 NOR2X1_LOC_15/Y INVX1_LOC_75/A 0.21fF
C393 INVX1_LOC_93/A INVX1_LOC_286/A 0.10fF
C394 NAND2X1_LOC_74/B INVX1_LOC_285/A 0.07fF
C395 INVX1_LOC_76/A NAND2X1_LOC_787/Y 0.13fF
C396 NOR2X1_LOC_541/Y NOR2X1_LOC_356/A 0.06fF
C397 INVX1_LOC_314/Y INVX1_LOC_43/A 0.02fF
C398 NOR2X1_LOC_589/A NAND2X1_LOC_364/A 0.03fF
C399 NAND2X1_LOC_1/Y INVX1_LOC_23/A 0.30fF
C400 NAND2X1_LOC_802/A NAND2X1_LOC_798/A 0.25fF
C401 NOR2X1_LOC_544/A INVX1_LOC_77/A 0.07fF
C402 NAND2X1_LOC_74/B NOR2X1_LOC_814/A 0.10fF
C403 NOR2X1_LOC_643/Y INVX1_LOC_40/A 0.05fF
C404 NOR2X1_LOC_778/B NOR2X1_LOC_551/B 0.03fF
C405 INVX1_LOC_170/A NOR2X1_LOC_76/A 0.01fF
C406 NAND2X1_LOC_731/Y NOR2X1_LOC_690/Y 0.02fF
C407 NOR2X1_LOC_384/Y NOR2X1_LOC_130/A 0.07fF
C408 NOR2X1_LOC_4/a_36_216# INVX1_LOC_216/A 0.00fF
C409 INVX1_LOC_13/A D_INPUT_2 0.01fF
C410 NOR2X1_LOC_561/Y INVX1_LOC_181/Y 0.02fF
C411 INVX1_LOC_26/Y INVX1_LOC_38/A 0.10fF
C412 INVX1_LOC_63/A NOR2X1_LOC_847/A 0.03fF
C413 INVX1_LOC_14/Y INVX1_LOC_53/A 0.10fF
C414 NAND2X1_LOC_739/B INVX1_LOC_10/A 0.09fF
C415 NAND2X1_LOC_44/a_36_24# INVX1_LOC_295/A 0.01fF
C416 INVX1_LOC_63/A INVX1_LOC_42/A 0.17fF
C417 INVX1_LOC_45/A NOR2X1_LOC_356/A 0.36fF
C418 INVX1_LOC_93/A INVX1_LOC_95/A 0.12fF
C419 NAND2X1_LOC_364/A INVX1_LOC_171/A 0.10fF
C420 NOR2X1_LOC_6/B NOR2X1_LOC_346/B 0.03fF
C421 NOR2X1_LOC_718/Y INVX1_LOC_22/A 0.05fF
C422 NOR2X1_LOC_541/Y NOR2X1_LOC_74/A 0.03fF
C423 INVX1_LOC_50/A NOR2X1_LOC_536/A 0.63fF
C424 NOR2X1_LOC_132/Y INVX1_LOC_16/A 0.03fF
C425 INVX1_LOC_136/A NOR2X1_LOC_246/Y 0.01fF
C426 NOR2X1_LOC_360/A INVX1_LOC_138/Y 0.06fF
C427 NAND2X1_LOC_726/Y NAND2X1_LOC_811/Y 0.01fF
C428 INVX1_LOC_153/Y INVX1_LOC_16/A 0.01fF
C429 NOR2X1_LOC_155/A INVX1_LOC_94/Y 0.03fF
C430 NOR2X1_LOC_655/B INVX1_LOC_206/A 0.10fF
C431 NAND2X1_LOC_740/B INVX1_LOC_141/Y 0.10fF
C432 INVX1_LOC_120/A INVX1_LOC_62/Y 0.24fF
C433 INVX1_LOC_57/A INVX1_LOC_280/A 0.07fF
C434 NAND2X1_LOC_21/Y GATE_662 0.02fF
C435 INVX1_LOC_5/A INVX1_LOC_139/A 0.02fF
C436 NOR2X1_LOC_315/Y INVX1_LOC_56/A 0.03fF
C437 INVX1_LOC_269/A INVX1_LOC_91/A 0.17fF
C438 NOR2X1_LOC_78/Y INVX1_LOC_16/Y 0.00fF
C439 INVX1_LOC_255/Y NOR2X1_LOC_516/Y 0.02fF
C440 NOR2X1_LOC_487/Y NOR2X1_LOC_693/Y 0.03fF
C441 NOR2X1_LOC_6/B INVX1_LOC_22/A 0.03fF
C442 NAND2X1_LOC_717/Y INVX1_LOC_280/Y 0.03fF
C443 NAND2X1_LOC_711/Y INPUT_0 0.02fF
C444 NOR2X1_LOC_272/Y INVX1_LOC_20/A 0.03fF
C445 NAND2X1_LOC_552/A NAND2X1_LOC_721/A 0.05fF
C446 NAND2X1_LOC_724/A NAND2X1_LOC_729/B 0.01fF
C447 INVX1_LOC_21/A NOR2X1_LOC_825/Y 0.68fF
C448 INVX1_LOC_5/A NAND2X1_LOC_721/A 0.00fF
C449 NOR2X1_LOC_261/Y NOR2X1_LOC_261/A 0.03fF
C450 INVX1_LOC_111/Y NOR2X1_LOC_500/Y 0.01fF
C451 INVX1_LOC_45/A NOR2X1_LOC_74/A 0.17fF
C452 NAND2X1_LOC_794/B VDD 0.63fF
C453 INVX1_LOC_177/A INVX1_LOC_16/A 0.03fF
C454 NOR2X1_LOC_590/A NOR2X1_LOC_334/A 0.02fF
C455 NOR2X1_LOC_68/A NOR2X1_LOC_163/Y 0.03fF
C456 INVX1_LOC_269/A INVX1_LOC_11/Y 0.03fF
C457 INPUT_3 INVX1_LOC_123/A 0.07fF
C458 NAND2X1_LOC_555/Y INVX1_LOC_201/A 0.11fF
C459 NOR2X1_LOC_67/Y NAND2X1_LOC_206/B -0.00fF
C460 INVX1_LOC_1/A NOR2X1_LOC_209/A 0.00fF
C461 NOR2X1_LOC_781/Y NAND2X1_LOC_654/B 0.01fF
C462 NOR2X1_LOC_568/A NOR2X1_LOC_74/A 0.07fF
C463 INVX1_LOC_50/A NAND2X1_LOC_93/B 0.03fF
C464 NOR2X1_LOC_356/A INVX1_LOC_71/A 0.15fF
C465 NOR2X1_LOC_552/a_36_216# INVX1_LOC_77/A 0.02fF
C466 NOR2X1_LOC_770/A NOR2X1_LOC_770/Y 0.17fF
C467 NOR2X1_LOC_322/Y NOR2X1_LOC_91/Y 0.01fF
C468 NAND2X1_LOC_9/Y INVX1_LOC_118/A 0.08fF
C469 INVX1_LOC_45/A NOR2X1_LOC_9/Y 0.41fF
C470 INVX1_LOC_240/A NAND2X1_LOC_795/Y 0.01fF
C471 INVX1_LOC_233/A INVX1_LOC_118/A 0.07fF
C472 NAND2X1_LOC_736/Y NOR2X1_LOC_576/B 0.06fF
C473 INVX1_LOC_280/Y INVX1_LOC_16/A 0.03fF
C474 INVX1_LOC_78/A INVX1_LOC_63/A 0.13fF
C475 NOR2X1_LOC_68/A NOR2X1_LOC_74/Y 0.03fF
C476 INVX1_LOC_178/A NAND2X1_LOC_721/A 0.14fF
C477 INVX1_LOC_49/A NAND2X1_LOC_842/B 0.21fF
C478 INVX1_LOC_34/A INVX1_LOC_89/A 1.81fF
C479 NAND2X1_LOC_860/A NAND2X1_LOC_243/Y 0.01fF
C480 INVX1_LOC_48/Y VDD 1.04fF
C481 NOR2X1_LOC_216/B NAND2X1_LOC_215/A 0.12fF
C482 INVX1_LOC_103/A NAND2X1_LOC_469/B 0.08fF
C483 NOR2X1_LOC_544/A NOR2X1_LOC_687/Y 0.03fF
C484 NOR2X1_LOC_773/Y INVX1_LOC_1/Y 0.07fF
C485 INVX1_LOC_13/A NOR2X1_LOC_620/B 0.05fF
C486 NOR2X1_LOC_15/Y NAND2X1_LOC_453/A 0.03fF
C487 NOR2X1_LOC_309/Y NAND2X1_LOC_861/Y 0.01fF
C488 NAND2X1_LOC_223/A INVX1_LOC_19/A 0.03fF
C489 INVX1_LOC_174/A NAND2X1_LOC_422/a_36_24# 0.00fF
C490 NAND2X1_LOC_477/Y NOR2X1_LOC_438/Y 0.04fF
C491 INVX1_LOC_120/A NOR2X1_LOC_844/A 0.02fF
C492 NAND2X1_LOC_371/a_36_24# NOR2X1_LOC_337/A 0.00fF
C493 NOR2X1_LOC_309/Y NOR2X1_LOC_150/a_36_216# 0.00fF
C494 INVX1_LOC_14/A INVX1_LOC_178/Y 0.35fF
C495 NAND2X1_LOC_23/a_36_24# INVX1_LOC_3/A 0.00fF
C496 NOR2X1_LOC_210/B NAND2X1_LOC_158/a_36_24# 0.01fF
C497 INVX1_LOC_255/Y INVX1_LOC_172/Y 0.21fF
C498 INVX1_LOC_246/A NOR2X1_LOC_56/Y 0.00fF
C499 INVX1_LOC_18/Y INVX1_LOC_19/A 0.32fF
C500 NAND2X1_LOC_553/A INVX1_LOC_118/A 0.02fF
C501 INVX1_LOC_24/A NOR2X1_LOC_188/A 0.03fF
C502 NAND2X1_LOC_352/B INVX1_LOC_95/Y 0.00fF
C503 NOR2X1_LOC_142/Y NOR2X1_LOC_772/A 0.02fF
C504 INVX1_LOC_256/Y INVX1_LOC_164/A 0.16fF
C505 INVX1_LOC_71/A NOR2X1_LOC_74/A 0.25fF
C506 NOR2X1_LOC_639/a_36_216# INVX1_LOC_191/Y 0.00fF
C507 NOR2X1_LOC_65/B INVX1_LOC_63/A 0.17fF
C508 D_INPUT_0 NOR2X1_LOC_537/Y 0.03fF
C509 INVX1_LOC_103/A NOR2X1_LOC_447/B 0.03fF
C510 D_INPUT_0 NAND2X1_LOC_338/B 0.23fF
C511 INVX1_LOC_93/A INVX1_LOC_54/A 0.07fF
C512 INVX1_LOC_193/Y NOR2X1_LOC_713/B 0.16fF
C513 INVX1_LOC_50/A NOR2X1_LOC_661/A 0.18fF
C514 NOR2X1_LOC_856/B NOR2X1_LOC_863/B 0.09fF
C515 NOR2X1_LOC_301/A INVX1_LOC_29/A 0.03fF
C516 INVX1_LOC_71/A NOR2X1_LOC_9/Y 0.10fF
C517 NAND2X1_LOC_231/Y INVX1_LOC_89/A 0.61fF
C518 INVX1_LOC_33/A INVX1_LOC_42/Y 0.05fF
C519 D_INPUT_0 NAND2X1_LOC_323/B 0.13fF
C520 INVX1_LOC_5/A INVX1_LOC_117/Y 0.26fF
C521 NOR2X1_LOC_666/Y INVX1_LOC_10/Y 0.05fF
C522 NOR2X1_LOC_329/B NAND2X1_LOC_477/A 0.09fF
C523 INVX1_LOC_246/A VDD 0.12fF
C524 INVX1_LOC_286/A NOR2X1_LOC_303/Y 0.01fF
C525 INVX1_LOC_225/A INVX1_LOC_73/A 0.07fF
C526 NOR2X1_LOC_120/a_36_216# NOR2X1_LOC_709/A 0.01fF
C527 INVX1_LOC_28/A INVX1_LOC_177/A 0.03fF
C528 NOR2X1_LOC_704/Y NOR2X1_LOC_374/A 0.02fF
C529 NOR2X1_LOC_209/Y NOR2X1_LOC_738/A 0.02fF
C530 INVX1_LOC_271/Y NOR2X1_LOC_270/a_36_216# 0.01fF
C531 INVX1_LOC_101/Y INVX1_LOC_9/A 0.00fF
C532 NOR2X1_LOC_784/Y NOR2X1_LOC_148/Y 0.04fF
C533 INVX1_LOC_280/Y INVX1_LOC_28/A 0.03fF
C534 INVX1_LOC_75/A NAND2X1_LOC_141/A 0.01fF
C535 NOR2X1_LOC_226/A INVX1_LOC_146/A 0.03fF
C536 INVX1_LOC_75/A INVX1_LOC_96/Y 0.05fF
C537 INVX1_LOC_161/Y INVX1_LOC_38/A 0.14fF
C538 NOR2X1_LOC_315/Y NOR2X1_LOC_83/Y 0.04fF
C539 INVX1_LOC_200/Y NOR2X1_LOC_89/A 0.03fF
C540 NOR2X1_LOC_620/Y NOR2X1_LOC_78/A 0.07fF
C541 NAND2X1_LOC_9/Y NAND2X1_LOC_63/Y 0.19fF
C542 INVX1_LOC_201/Y NAND2X1_LOC_4/a_36_24# 0.03fF
C543 INVX1_LOC_208/A NOR2X1_LOC_755/a_36_216# -0.01fF
C544 NOR2X1_LOC_137/A INVX1_LOC_10/A 0.03fF
C545 NOR2X1_LOC_513/Y INVX1_LOC_54/A 0.05fF
C546 INVX1_LOC_61/Y NOR2X1_LOC_536/A 0.03fF
C547 INVX1_LOC_181/Y INVX1_LOC_76/A 0.10fF
C548 INVX1_LOC_30/A INVX1_LOC_33/Y 0.01fF
C549 NAND2X1_LOC_773/Y NOR2X1_LOC_831/B 0.01fF
C550 NAND2X1_LOC_569/A NOR2X1_LOC_45/B -0.02fF
C551 INVX1_LOC_1/A NOR2X1_LOC_197/B 0.03fF
C552 INVX1_LOC_21/A INVX1_LOC_84/A 0.10fF
C553 INVX1_LOC_143/A NOR2X1_LOC_188/A 0.10fF
C554 INVX1_LOC_17/A INVX1_LOC_152/A 0.26fF
C555 INVX1_LOC_49/A NOR2X1_LOC_545/B 0.05fF
C556 INVX1_LOC_43/Y INVX1_LOC_127/A 0.01fF
C557 INVX1_LOC_207/A NOR2X1_LOC_396/Y -0.01fF
C558 INVX1_LOC_143/A NOR2X1_LOC_548/B 0.10fF
C559 NOR2X1_LOC_844/Y NOR2X1_LOC_865/A 0.06fF
C560 INVX1_LOC_50/Y INVX1_LOC_186/Y 0.15fF
C561 NAND2X1_LOC_9/Y NAND2X1_LOC_455/B 0.70fF
C562 INVX1_LOC_54/Y INVX1_LOC_286/A 0.01fF
C563 NOR2X1_LOC_392/Y NOR2X1_LOC_672/a_36_216# 0.01fF
C564 INVX1_LOC_63/A NOR2X1_LOC_655/a_36_216# 0.00fF
C565 INVX1_LOC_90/A INVX1_LOC_62/A 0.18fF
C566 D_INPUT_1 INVX1_LOC_32/A 9.91fF
C567 NOR2X1_LOC_350/A VDD 0.43fF
C568 NOR2X1_LOC_189/A VDD -0.00fF
C569 INVX1_LOC_34/A NOR2X1_LOC_24/Y 0.04fF
C570 INVX1_LOC_21/A NAND2X1_LOC_651/B 0.61fF
C571 INVX1_LOC_78/A NOR2X1_LOC_65/Y 0.03fF
C572 INVX1_LOC_17/A NAND2X1_LOC_606/a_36_24# 0.00fF
C573 NOR2X1_LOC_281/Y NOR2X1_LOC_301/A 0.01fF
C574 NOR2X1_LOC_794/B NOR2X1_LOC_197/B 0.07fF
C575 NOR2X1_LOC_19/B NOR2X1_LOC_99/B 0.01fF
C576 NOR2X1_LOC_510/Y INVX1_LOC_109/A 0.01fF
C577 NOR2X1_LOC_348/B INVX1_LOC_188/Y 0.01fF
C578 INVX1_LOC_285/Y INVX1_LOC_16/A 0.03fF
C579 INVX1_LOC_231/Y VDD 0.44fF
C580 NOR2X1_LOC_460/B VDD -0.00fF
C581 NOR2X1_LOC_89/A NOR2X1_LOC_406/A 0.00fF
C582 NAND2X1_LOC_181/Y INVX1_LOC_98/A 0.30fF
C583 NAND2X1_LOC_842/B INPUT_1 0.01fF
C584 INVX1_LOC_269/A INVX1_LOC_203/A 0.03fF
C585 INVX1_LOC_39/A NOR2X1_LOC_671/Y 0.00fF
C586 INVX1_LOC_223/Y INVX1_LOC_99/A 0.01fF
C587 NOR2X1_LOC_232/Y INVX1_LOC_203/A 0.02fF
C588 INVX1_LOC_207/Y NOR2X1_LOC_575/Y 0.15fF
C589 NOR2X1_LOC_554/B NOR2X1_LOC_656/Y 0.02fF
C590 NAND2X1_LOC_845/a_36_24# NOR2X1_LOC_536/A 0.00fF
C591 INVX1_LOC_36/A INVX1_LOC_291/A 0.07fF
C592 INVX1_LOC_45/A NOR2X1_LOC_650/a_36_216# 0.00fF
C593 INVX1_LOC_18/A NAND2X1_LOC_260/a_36_24# 0.00fF
C594 NOR2X1_LOC_828/B INVX1_LOC_85/Y 0.03fF
C595 NAND2X1_LOC_348/A INVX1_LOC_62/A 0.32fF
C596 NOR2X1_LOC_568/A NOR2X1_LOC_650/a_36_216# 0.00fF
C597 INVX1_LOC_36/A NAND2X1_LOC_802/Y 0.04fF
C598 INVX1_LOC_93/A NOR2X1_LOC_48/B 0.01fF
C599 NOR2X1_LOC_45/B INVX1_LOC_316/Y 0.01fF
C600 INVX1_LOC_34/A NOR2X1_LOC_425/Y 0.04fF
C601 INVX1_LOC_177/A NOR2X1_LOC_35/Y 0.01fF
C602 NOR2X1_LOC_229/Y NOR2X1_LOC_45/B 0.29fF
C603 NOR2X1_LOC_773/Y INVX1_LOC_93/Y 1.13fF
C604 INVX1_LOC_80/Y D_INPUT_3 0.01fF
C605 NOR2X1_LOC_163/A NOR2X1_LOC_163/Y 0.01fF
C606 NOR2X1_LOC_123/B NOR2X1_LOC_74/A 0.00fF
C607 NOR2X1_LOC_78/B NAND2X1_LOC_212/Y 0.02fF
C608 INVX1_LOC_45/A NOR2X1_LOC_865/Y 0.24fF
C609 NOR2X1_LOC_371/a_36_216# NAND2X1_LOC_489/Y 0.00fF
C610 INVX1_LOC_32/A NOR2X1_LOC_652/Y 0.10fF
C611 NOR2X1_LOC_61/B NOR2X1_LOC_861/Y 0.15fF
C612 INVX1_LOC_23/A NAND2X1_LOC_61/Y 0.42fF
C613 INVX1_LOC_61/Y INVX1_LOC_3/A 0.07fF
C614 NAND2X1_LOC_562/B NAND2X1_LOC_721/A 0.02fF
C615 NOR2X1_LOC_543/A NOR2X1_LOC_355/B 0.04fF
C616 INVX1_LOC_89/A INPUT_0 0.20fF
C617 NOR2X1_LOC_84/Y VDD 2.14fF
C618 INVX1_LOC_45/A NOR2X1_LOC_243/B 0.02fF
C619 NOR2X1_LOC_68/A INVX1_LOC_179/A 0.06fF
C620 INVX1_LOC_14/A INVX1_LOC_12/A 0.09fF
C621 INVX1_LOC_31/A NAND2X1_LOC_42/a_36_24# 0.03fF
C622 NAND2X1_LOC_354/Y NOR2X1_LOC_88/Y 0.03fF
C623 INVX1_LOC_17/A INVX1_LOC_29/A 0.23fF
C624 INVX1_LOC_126/A NAND2X1_LOC_850/Y 0.05fF
C625 NOR2X1_LOC_123/B NOR2X1_LOC_9/Y 0.11fF
C626 NAND2X1_LOC_359/Y VDD 0.24fF
C627 NOR2X1_LOC_482/Y VDD 0.42fF
C628 INVX1_LOC_21/A INVX1_LOC_15/A 0.86fF
C629 NOR2X1_LOC_590/A INVX1_LOC_293/Y 0.05fF
C630 INVX1_LOC_216/A VDD 0.25fF
C631 INVX1_LOC_30/A INVX1_LOC_220/A 0.36fF
C632 NOR2X1_LOC_589/A NOR2X1_LOC_405/A 0.07fF
C633 INVX1_LOC_22/A INVX1_LOC_188/Y 0.01fF
C634 NOR2X1_LOC_483/B INVX1_LOC_19/A 0.02fF
C635 NOR2X1_LOC_769/B INVX1_LOC_296/A 0.02fF
C636 NOR2X1_LOC_773/a_36_216# NOR2X1_LOC_536/A 0.01fF
C637 NAND2X1_LOC_508/A INPUT_0 0.03fF
C638 NAND2X1_LOC_451/Y INVX1_LOC_37/A 0.01fF
C639 INVX1_LOC_16/A NOR2X1_LOC_137/B 0.12fF
C640 INVX1_LOC_136/A INVX1_LOC_285/A 0.31fF
C641 NOR2X1_LOC_78/B INVX1_LOC_14/Y 0.03fF
C642 INVX1_LOC_88/A INVX1_LOC_290/Y 0.79fF
C643 NOR2X1_LOC_598/B INVX1_LOC_296/A 0.03fF
C644 INVX1_LOC_136/A NOR2X1_LOC_814/A 0.20fF
C645 NOR2X1_LOC_816/A NOR2X1_LOC_669/A 0.03fF
C646 INVX1_LOC_102/Y NOR2X1_LOC_74/A 0.07fF
C647 INVX1_LOC_28/A INVX1_LOC_285/Y 0.01fF
C648 NAND2X1_LOC_555/Y INVX1_LOC_29/A 0.09fF
C649 INVX1_LOC_196/Y INVX1_LOC_78/Y 0.06fF
C650 NOR2X1_LOC_590/A NAND2X1_LOC_74/B 1.63fF
C651 NOR2X1_LOC_232/a_36_216# INVX1_LOC_3/Y 0.02fF
C652 INVX1_LOC_239/Y VDD -0.00fF
C653 NOR2X1_LOC_773/Y NAND2X1_LOC_721/A 0.08fF
C654 NOR2X1_LOC_299/Y INPUT_4 0.03fF
C655 NOR2X1_LOC_582/Y INVX1_LOC_84/A 0.00fF
C656 INVX1_LOC_83/A NOR2X1_LOC_448/A 0.01fF
C657 NOR2X1_LOC_554/B INVX1_LOC_63/A 0.49fF
C658 NOR2X1_LOC_86/A INVX1_LOC_20/A 0.05fF
C659 NOR2X1_LOC_134/Y INVX1_LOC_284/A 0.01fF
C660 VDD NOR2X1_LOC_374/B 0.22fF
C661 INVX1_LOC_171/A NOR2X1_LOC_405/A 0.08fF
C662 NAND2X1_LOC_113/a_36_24# NOR2X1_LOC_89/A 0.00fF
C663 INVX1_LOC_178/A NAND2X1_LOC_619/a_36_24# 0.00fF
C664 NOR2X1_LOC_709/B NOR2X1_LOC_709/A 0.00fF
C665 NOR2X1_LOC_791/Y INVX1_LOC_23/Y 0.02fF
C666 NAND2X1_LOC_735/B INVX1_LOC_46/A 0.03fF
C667 INVX1_LOC_290/A VDD 2.27fF
C668 NOR2X1_LOC_773/Y NOR2X1_LOC_323/a_36_216# 0.01fF
C669 INVX1_LOC_178/A INVX1_LOC_175/A 0.02fF
C670 INVX1_LOC_50/Y NOR2X1_LOC_843/B 0.06fF
C671 NOR2X1_LOC_717/Y INVX1_LOC_12/A 0.34fF
C672 NOR2X1_LOC_792/B NOR2X1_LOC_743/Y 0.03fF
C673 NAND2X1_LOC_390/A NOR2X1_LOC_176/a_36_216# 0.00fF
C674 NOR2X1_LOC_172/Y NOR2X1_LOC_841/A 0.01fF
C675 NOR2X1_LOC_68/A NAND2X1_LOC_215/a_36_24# 0.00fF
C676 NOR2X1_LOC_459/A D_GATE_479 0.01fF
C677 NOR2X1_LOC_152/Y INVX1_LOC_63/A 0.07fF
C678 INVX1_LOC_250/A NOR2X1_LOC_89/A 0.04fF
C679 INVX1_LOC_83/A D_INPUT_3 0.07fF
C680 INVX1_LOC_28/A NOR2X1_LOC_137/B 0.03fF
C681 INVX1_LOC_58/A NAND2X1_LOC_796/B -0.01fF
C682 INVX1_LOC_73/A NAND2X1_LOC_642/Y 0.68fF
C683 INVX1_LOC_17/A INVX1_LOC_298/Y 0.02fF
C684 NOR2X1_LOC_537/Y INVX1_LOC_46/Y 0.07fF
C685 NAND2X1_LOC_739/B INVX1_LOC_12/A 0.05fF
C686 NAND2X1_LOC_338/B INVX1_LOC_46/Y 0.01fF
C687 NOR2X1_LOC_718/Y INVX1_LOC_186/Y 0.03fF
C688 NOR2X1_LOC_440/B INVX1_LOC_29/Y 0.10fF
C689 INVX1_LOC_41/A NOR2X1_LOC_691/B 0.03fF
C690 NAND2X1_LOC_9/Y INVX1_LOC_39/A 0.07fF
C691 INVX1_LOC_21/A INVX1_LOC_108/Y 0.03fF
C692 INVX1_LOC_214/A NOR2X1_LOC_88/Y 0.03fF
C693 INVX1_LOC_75/A NOR2X1_LOC_708/A 0.09fF
C694 NAND2X1_LOC_785/Y INVX1_LOC_84/A 0.01fF
C695 NOR2X1_LOC_860/B NAND2X1_LOC_291/B 0.02fF
C696 INVX1_LOC_33/A INVX1_LOC_19/A 0.31fF
C697 NOR2X1_LOC_667/A NOR2X1_LOC_88/Y 0.07fF
C698 INVX1_LOC_21/A INVX1_LOC_278/A 0.10fF
C699 INVX1_LOC_248/A NOR2X1_LOC_88/Y 0.07fF
C700 INVX1_LOC_298/Y NOR2X1_LOC_471/Y 0.12fF
C701 INVX1_LOC_222/A NOR2X1_LOC_405/A 0.06fF
C702 NOR2X1_LOC_272/Y INVX1_LOC_64/A 0.22fF
C703 NOR2X1_LOC_87/B NAND2X1_LOC_206/Y 0.00fF
C704 INVX1_LOC_2/A INVX1_LOC_119/Y 0.02fF
C705 INVX1_LOC_62/A INVX1_LOC_38/A 0.12fF
C706 INVX1_LOC_100/A NOR2X1_LOC_124/A 0.24fF
C707 NAND2X1_LOC_53/Y NOR2X1_LOC_383/B 0.07fF
C708 NOR2X1_LOC_793/Y INVX1_LOC_23/A 0.21fF
C709 NAND2X1_LOC_364/A INVX1_LOC_4/A 0.14fF
C710 NAND2X1_LOC_518/a_36_24# NAND2X1_LOC_74/B 0.01fF
C711 NAND2X1_LOC_361/Y NOR2X1_LOC_89/A 0.01fF
C712 NOR2X1_LOC_700/Y INVX1_LOC_118/A 0.11fF
C713 INVX1_LOC_35/A NOR2X1_LOC_92/Y 0.06fF
C714 NOR2X1_LOC_226/A INVX1_LOC_119/Y 0.07fF
C715 NAND2X1_LOC_555/Y NOR2X1_LOC_33/Y -0.00fF
C716 INVX1_LOC_256/A INVX1_LOC_50/A 0.20fF
C717 INVX1_LOC_299/A NOR2X1_LOC_598/B 0.27fF
C718 INVX1_LOC_39/A NAND2X1_LOC_553/A 0.02fF
C719 INVX1_LOC_140/A NAND2X1_LOC_721/A 0.07fF
C720 NAND2X1_LOC_538/Y NOR2X1_LOC_591/A 0.06fF
C721 NOR2X1_LOC_667/A INVX1_LOC_84/A 0.10fF
C722 NOR2X1_LOC_296/Y D_INPUT_1 0.65fF
C723 NOR2X1_LOC_403/B INVX1_LOC_32/A 0.02fF
C724 INVX1_LOC_35/A INVX1_LOC_24/Y 0.01fF
C725 NOR2X1_LOC_471/Y INVX1_LOC_204/A 0.04fF
C726 INVX1_LOC_248/A INVX1_LOC_84/A 0.03fF
C727 D_INPUT_2 INVX1_LOC_32/A 0.02fF
C728 NOR2X1_LOC_714/Y INVX1_LOC_19/A 0.06fF
C729 NOR2X1_LOC_453/Y NOR2X1_LOC_223/B 0.01fF
C730 INVX1_LOC_30/A INVX1_LOC_23/Y 0.01fF
C731 NOR2X1_LOC_609/A NOR2X1_LOC_334/Y 0.02fF
C732 NOR2X1_LOC_285/A NOR2X1_LOC_590/A 0.00fF
C733 NOR2X1_LOC_802/A INVX1_LOC_69/A 0.19fF
C734 D_INPUT_1 INPUT_3 0.87fF
C735 INVX1_LOC_17/A NAND2X1_LOC_385/a_36_24# 0.01fF
C736 NOR2X1_LOC_612/B INVX1_LOC_12/A 0.07fF
C737 NOR2X1_LOC_93/a_36_216# NOR2X1_LOC_671/Y 0.00fF
C738 NOR2X1_LOC_237/Y NOR2X1_LOC_89/a_36_216# 0.00fF
C739 NAND2X1_LOC_139/A INVX1_LOC_3/Y 0.02fF
C740 INVX1_LOC_40/A INVX1_LOC_19/A 0.07fF
C741 INVX1_LOC_2/A INVX1_LOC_284/A -0.00fF
C742 INVX1_LOC_105/A NAND2X1_LOC_470/B 0.07fF
C743 NOR2X1_LOC_357/Y NOR2X1_LOC_144/a_36_216# 0.01fF
C744 INVX1_LOC_41/A NOR2X1_LOC_620/a_36_216# 0.00fF
C745 NOR2X1_LOC_7/Y INVX1_LOC_46/A 0.01fF
C746 NOR2X1_LOC_824/A NAND2X1_LOC_579/A 0.10fF
C747 NOR2X1_LOC_82/A INVX1_LOC_5/A 0.13fF
C748 INVX1_LOC_289/Y INVX1_LOC_178/A 0.55fF
C749 NOR2X1_LOC_172/Y INVX1_LOC_128/A 0.01fF
C750 NOR2X1_LOC_141/a_36_216# NAND2X1_LOC_469/B 0.00fF
C751 INVX1_LOC_224/Y NOR2X1_LOC_791/A 0.00fF
C752 INVX1_LOC_89/A NAND2X1_LOC_240/a_36_24# 0.01fF
C753 INVX1_LOC_309/A NOR2X1_LOC_492/Y 0.01fF
C754 NOR2X1_LOC_74/A NOR2X1_LOC_331/B 1.55fF
C755 INVX1_LOC_96/Y INVX1_LOC_283/A 0.15fF
C756 NOR2X1_LOC_577/Y INVX1_LOC_273/A -0.01fF
C757 INVX1_LOC_160/A VDD 0.09fF
C758 INVX1_LOC_12/Y NOR2X1_LOC_114/A 0.20fF
C759 NOR2X1_LOC_360/Y NAND2X1_LOC_96/a_36_24# 0.01fF
C760 INVX1_LOC_11/A NOR2X1_LOC_406/A 0.01fF
C761 INVX1_LOC_16/A NAND2X1_LOC_81/B 0.01fF
C762 INVX1_LOC_90/A NOR2X1_LOC_841/A 0.08fF
C763 INVX1_LOC_12/Y INVX1_LOC_91/A 0.10fF
C764 INVX1_LOC_78/Y INVX1_LOC_44/A 0.00fF
C765 NOR2X1_LOC_361/B INVX1_LOC_48/Y 0.01fF
C766 NOR2X1_LOC_590/A NOR2X1_LOC_845/a_36_216# 0.00fF
C767 NOR2X1_LOC_510/Y INVX1_LOC_246/A 0.03fF
C768 INVX1_LOC_103/A INVX1_LOC_52/Y 0.04fF
C769 NOR2X1_LOC_590/a_36_216# INVX1_LOC_179/A 0.00fF
C770 NOR2X1_LOC_78/A INVX1_LOC_117/A 0.10fF
C771 NOR2X1_LOC_152/Y NOR2X1_LOC_65/Y 0.03fF
C772 NOR2X1_LOC_99/B NOR2X1_LOC_126/a_36_216# 0.01fF
C773 NOR2X1_LOC_91/A NOR2X1_LOC_753/Y 2.27fF
C774 NOR2X1_LOC_825/Y NOR2X1_LOC_670/Y 0.00fF
C775 NOR2X1_LOC_272/Y INVX1_LOC_43/Y 0.01fF
C776 NAND2X1_LOC_212/Y INVX1_LOC_46/A 0.10fF
C777 NOR2X1_LOC_667/A INVX1_LOC_15/A 0.07fF
C778 INVX1_LOC_25/A NOR2X1_LOC_191/B 0.14fF
C779 INVX1_LOC_33/A INVX1_LOC_26/Y 0.03fF
C780 INVX1_LOC_1/Y INVX1_LOC_42/A 0.03fF
C781 INVX1_LOC_93/A NOR2X1_LOC_441/Y 0.00fF
C782 INVX1_LOC_248/A INVX1_LOC_15/A 0.94fF
C783 NOR2X1_LOC_589/A INVX1_LOC_109/Y 0.20fF
C784 NOR2X1_LOC_199/B INVX1_LOC_29/A 0.03fF
C785 INVX1_LOC_64/A NAND2X1_LOC_364/A 0.09fF
C786 INVX1_LOC_11/Y NOR2X1_LOC_492/Y 0.03fF
C787 NOR2X1_LOC_97/B NAND2X1_LOC_291/B 0.04fF
C788 NOR2X1_LOC_591/Y NAND2X1_LOC_175/Y 0.09fF
C789 INVX1_LOC_200/A INVX1_LOC_14/A 0.01fF
C790 NAND2X1_LOC_660/A INVX1_LOC_94/Y 0.29fF
C791 NAND2X1_LOC_21/Y INVX1_LOC_173/A 0.16fF
C792 NOR2X1_LOC_106/Y INVX1_LOC_53/A 0.04fF
C793 INVX1_LOC_289/Y NOR2X1_LOC_816/A 0.00fF
C794 NOR2X1_LOC_139/Y INVX1_LOC_9/A 0.01fF
C795 NAND2X1_LOC_465/Y NAND2X1_LOC_99/A 0.01fF
C796 NOR2X1_LOC_497/Y NAND2X1_LOC_489/Y 0.01fF
C797 INVX1_LOC_14/Y INVX1_LOC_46/A 0.03fF
C798 NOR2X1_LOC_687/Y NOR2X1_LOC_685/Y 0.14fF
C799 INVX1_LOC_224/Y NOR2X1_LOC_121/Y 0.01fF
C800 NOR2X1_LOC_208/Y NOR2X1_LOC_665/a_36_216# 0.01fF
C801 INVX1_LOC_18/A INVX1_LOC_50/Y 0.12fF
C802 NOR2X1_LOC_828/B NAND2X1_LOC_782/B 0.07fF
C803 NAND2X1_LOC_363/B NAND2X1_LOC_517/a_36_24# 0.00fF
C804 NOR2X1_LOC_313/Y NOR2X1_LOC_697/Y 0.01fF
C805 INVX1_LOC_58/A NAND2X1_LOC_139/A 0.03fF
C806 NAND2X1_LOC_51/B INVX1_LOC_84/A 0.08fF
C807 NOR2X1_LOC_446/A NOR2X1_LOC_457/A 0.03fF
C808 NOR2X1_LOC_52/B NOR2X1_LOC_113/a_36_216# 0.01fF
C809 NOR2X1_LOC_307/B NOR2X1_LOC_307/Y 0.01fF
C810 INVX1_LOC_224/A NAND2X1_LOC_113/a_36_24# 0.00fF
C811 INVX1_LOC_28/A NAND2X1_LOC_81/B 0.00fF
C812 INPUT_1 INVX1_LOC_284/A 0.11fF
C813 INVX1_LOC_200/Y NOR2X1_LOC_52/B 0.03fF
C814 INVX1_LOC_21/A NOR2X1_LOC_168/Y 0.73fF
C815 NOR2X1_LOC_772/B INVX1_LOC_77/A 0.07fF
C816 INVX1_LOC_311/A INVX1_LOC_84/A 0.07fF
C817 NAND2X1_LOC_466/Y INVX1_LOC_53/A 0.07fF
C818 INVX1_LOC_34/A NOR2X1_LOC_392/Y 0.04fF
C819 NOR2X1_LOC_91/A NOR2X1_LOC_67/A 0.04fF
C820 INVX1_LOC_35/A INVX1_LOC_41/A 0.13fF
C821 INVX1_LOC_1/Y INVX1_LOC_78/A 5.95fF
C822 INVX1_LOC_35/A INVX1_LOC_201/Y 0.32fF
C823 INVX1_LOC_251/Y INVX1_LOC_57/A 0.00fF
C824 INVX1_LOC_13/Y INVX1_LOC_77/A 0.03fF
C825 INVX1_LOC_266/A INVX1_LOC_18/A 0.00fF
C826 NOR2X1_LOC_636/B INVX1_LOC_30/A 0.05fF
C827 INVX1_LOC_133/Y INVX1_LOC_23/A 0.00fF
C828 NOR2X1_LOC_439/B INVX1_LOC_99/A 0.03fF
C829 NOR2X1_LOC_250/Y INVX1_LOC_45/A 0.09fF
C830 INVX1_LOC_56/A NAND2X1_LOC_99/A 0.11fF
C831 NAND2X1_LOC_363/B NAND2X1_LOC_116/A 0.03fF
C832 INVX1_LOC_17/A NAND2X1_LOC_634/Y 0.39fF
C833 INVX1_LOC_24/A NAND2X1_LOC_326/A 0.12fF
C834 INVX1_LOC_75/A INVX1_LOC_99/A 0.03fF
C835 NOR2X1_LOC_67/A INVX1_LOC_23/A 0.07fF
C836 INVX1_LOC_250/A INVX1_LOC_11/A 0.02fF
C837 NOR2X1_LOC_500/Y NOR2X1_LOC_383/B 0.08fF
C838 INVX1_LOC_226/Y NOR2X1_LOC_383/B 0.01fF
C839 NOR2X1_LOC_65/B INVX1_LOC_1/Y 0.17fF
C840 INVX1_LOC_1/A NOR2X1_LOC_191/B 0.26fF
C841 INVX1_LOC_21/A NAND2X1_LOC_21/Y 0.08fF
C842 NOR2X1_LOC_411/Y NAND2X1_LOC_33/Y 0.07fF
C843 NOR2X1_LOC_88/Y NOR2X1_LOC_670/Y 0.01fF
C844 INVX1_LOC_35/A INVX1_LOC_64/Y 0.03fF
C845 INVX1_LOC_124/A NOR2X1_LOC_772/B -0.04fF
C846 NOR2X1_LOC_45/B NOR2X1_LOC_662/A 0.10fF
C847 NOR2X1_LOC_632/Y INVX1_LOC_270/A 0.00fF
C848 NOR2X1_LOC_828/A NOR2X1_LOC_334/Y 0.03fF
C849 NOR2X1_LOC_19/B NOR2X1_LOC_28/a_36_216# 0.02fF
C850 INVX1_LOC_48/Y NOR2X1_LOC_132/Y 0.01fF
C851 NOR2X1_LOC_15/Y NOR2X1_LOC_577/Y 0.13fF
C852 INVX1_LOC_304/A INVX1_LOC_84/A 0.02fF
C853 INVX1_LOC_45/A INVX1_LOC_124/Y 0.07fF
C854 INVX1_LOC_136/A NOR2X1_LOC_590/A 0.13fF
C855 INVX1_LOC_88/A INVX1_LOC_77/A 0.13fF
C856 INVX1_LOC_1/A INVX1_LOC_283/Y 0.04fF
C857 INVX1_LOC_124/A INVX1_LOC_13/Y 0.06fF
C858 INVX1_LOC_28/A INVX1_LOC_4/Y 0.02fF
C859 NOR2X1_LOC_250/Y INVX1_LOC_71/A 0.02fF
C860 NOR2X1_LOC_644/A NAND2X1_LOC_454/Y 0.05fF
C861 INVX1_LOC_10/A NOR2X1_LOC_383/B 0.10fF
C862 NOR2X1_LOC_122/A INVX1_LOC_33/A 0.00fF
C863 NOR2X1_LOC_246/A NOR2X1_LOC_318/A 0.04fF
C864 INVX1_LOC_84/A NOR2X1_LOC_670/Y 0.07fF
C865 NOR2X1_LOC_598/B INVX1_LOC_268/Y 0.03fF
C866 NAND2X1_LOC_51/B INVX1_LOC_15/A 0.01fF
C867 INVX1_LOC_235/Y INVX1_LOC_194/A 0.37fF
C868 NAND2X1_LOC_363/B INVX1_LOC_232/A 0.01fF
C869 INVX1_LOC_35/A NOR2X1_LOC_211/A 0.49fF
C870 NAND2X1_LOC_570/a_36_24# INVX1_LOC_178/A 0.00fF
C871 INVX1_LOC_235/Y NOR2X1_LOC_399/A 0.02fF
C872 NAND2X1_LOC_563/Y INVX1_LOC_163/A 0.02fF
C873 NOR2X1_LOC_641/B NOR2X1_LOC_68/A 0.02fF
C874 INPUT_3 D_INPUT_2 0.11fF
C875 NOR2X1_LOC_486/Y INVX1_LOC_19/A 0.03fF
C876 INVX1_LOC_233/Y INVX1_LOC_16/A 0.40fF
C877 INVX1_LOC_224/Y D_INPUT_0 0.05fF
C878 NAND2X1_LOC_739/B NAND2X1_LOC_733/Y 0.05fF
C879 INVX1_LOC_11/A NAND2X1_LOC_361/Y 0.07fF
C880 INVX1_LOC_17/A NAND2X1_LOC_310/a_36_24# 0.00fF
C881 INVX1_LOC_103/A INVX1_LOC_63/Y 0.21fF
C882 NOR2X1_LOC_567/B NAND2X1_LOC_72/B 0.01fF
C883 NAND2X1_LOC_794/B INVX1_LOC_280/Y 0.27fF
C884 NOR2X1_LOC_742/A INVX1_LOC_78/A 0.07fF
C885 INVX1_LOC_33/A INVX1_LOC_161/Y 0.07fF
C886 NOR2X1_LOC_318/B INVX1_LOC_42/A 0.07fF
C887 INVX1_LOC_17/A INVX1_LOC_8/A 0.00fF
C888 NOR2X1_LOC_751/Y NOR2X1_LOC_68/A 0.05fF
C889 NOR2X1_LOC_315/Y NOR2X1_LOC_271/a_36_216# 0.01fF
C890 INVX1_LOC_58/A NOR2X1_LOC_207/a_36_216# 0.00fF
C891 NAND2X1_LOC_331/a_36_24# INVX1_LOC_23/A 0.00fF
C892 NOR2X1_LOC_468/a_36_216# NOR2X1_LOC_717/A 0.01fF
C893 INVX1_LOC_27/A INVX1_LOC_43/A 0.04fF
C894 INVX1_LOC_59/A NAND2X1_LOC_549/B 0.01fF
C895 INVX1_LOC_124/A INVX1_LOC_88/A 0.01fF
C896 INVX1_LOC_38/A NOR2X1_LOC_841/A 0.03fF
C897 D_INPUT_0 NAND2X1_LOC_415/a_36_24# 0.01fF
C898 INVX1_LOC_93/Y INVX1_LOC_42/A 0.19fF
C899 NOR2X1_LOC_361/B NOR2X1_LOC_84/Y 0.10fF
C900 D_INPUT_0 NAND2X1_LOC_793/B 0.05fF
C901 NAND2X1_LOC_778/Y INVX1_LOC_22/A 0.00fF
C902 INVX1_LOC_27/A INVX1_LOC_208/Y 0.06fF
C903 NOR2X1_LOC_78/A INVX1_LOC_3/Y 0.01fF
C904 INVX1_LOC_34/A NOR2X1_LOC_599/Y 0.03fF
C905 INVX1_LOC_77/A NOR2X1_LOC_500/B 3.69fF
C906 NAND2X1_LOC_325/Y INVX1_LOC_31/A 0.01fF
C907 NAND2X1_LOC_187/a_36_24# INVX1_LOC_18/A 0.01fF
C908 NAND2X1_LOC_711/Y NAND2X1_LOC_811/Y 0.00fF
C909 INVX1_LOC_49/A INVX1_LOC_72/A 0.07fF
C910 INVX1_LOC_180/Y NAND2X1_LOC_798/B 0.21fF
C911 INVX1_LOC_1/A NOR2X1_LOC_568/a_36_216# 0.00fF
C912 D_INPUT_3 NOR2X1_LOC_671/Y 0.05fF
C913 VDD INVX1_LOC_261/Y 0.33fF
C914 NOR2X1_LOC_215/Y NOR2X1_LOC_759/Y 0.01fF
C915 INVX1_LOC_55/Y NOR2X1_LOC_678/A 0.03fF
C916 NOR2X1_LOC_240/Y INVX1_LOC_89/A 0.04fF
C917 INVX1_LOC_304/A INVX1_LOC_15/A 0.07fF
C918 INVX1_LOC_255/A INVX1_LOC_15/A 0.11fF
C919 VDD INVX1_LOC_114/Y 0.26fF
C920 NOR2X1_LOC_405/A INVX1_LOC_4/A 0.07fF
C921 NOR2X1_LOC_468/Y INVX1_LOC_56/Y -0.03fF
C922 INVX1_LOC_258/Y NOR2X1_LOC_32/Y 0.00fF
C923 NOR2X1_LOC_15/Y INVX1_LOC_22/A 13.29fF
C924 NAND2X1_LOC_714/B NAND2X1_LOC_854/B 0.30fF
C925 INVX1_LOC_286/Y INVX1_LOC_221/A -0.02fF
C926 NAND2X1_LOC_363/B NOR2X1_LOC_775/Y 0.03fF
C927 NOR2X1_LOC_82/A NOR2X1_LOC_773/Y 0.00fF
C928 NOR2X1_LOC_318/B INVX1_LOC_78/A 0.08fF
C929 INVX1_LOC_34/A NOR2X1_LOC_86/Y 0.01fF
C930 NOR2X1_LOC_205/Y INVX1_LOC_16/A 0.06fF
C931 NAND2X1_LOC_833/Y NOR2X1_LOC_91/Y 0.73fF
C932 NOR2X1_LOC_134/Y NAND2X1_LOC_338/B 0.19fF
C933 INVX1_LOC_217/Y INVX1_LOC_217/A -0.03fF
C934 NAND2X1_LOC_721/A INVX1_LOC_42/A 0.05fF
C935 NOR2X1_LOC_74/A NOR2X1_LOC_493/A 0.03fF
C936 INVX1_LOC_276/A INVX1_LOC_31/A 0.08fF
C937 INVX1_LOC_50/A INVX1_LOC_69/Y 0.07fF
C938 INVX1_LOC_93/Y INVX1_LOC_78/A 0.07fF
C939 INVX1_LOC_278/Y NOR2X1_LOC_816/A 0.03fF
C940 NAND2X1_LOC_392/A NAND2X1_LOC_793/Y 0.02fF
C941 NAND2X1_LOC_783/A NAND2X1_LOC_326/A 0.10fF
C942 INVX1_LOC_303/A INVX1_LOC_77/A 0.14fF
C943 INVX1_LOC_116/A NOR2X1_LOC_593/Y 0.08fF
C944 NOR2X1_LOC_67/A INVX1_LOC_31/A 0.56fF
C945 INVX1_LOC_291/A INVX1_LOC_63/A 0.07fF
C946 INVX1_LOC_38/A INPUT_7 0.12fF
C947 NOR2X1_LOC_6/B INVX1_LOC_18/A -0.01fF
C948 INVX1_LOC_99/Y INVX1_LOC_182/A 0.01fF
C949 VDD NOR2X1_LOC_467/A 0.22fF
C950 NOR2X1_LOC_35/Y INVX1_LOC_4/Y 0.11fF
C951 NAND2X1_LOC_462/a_36_24# INVX1_LOC_253/Y 0.00fF
C952 INPUT_0 NOR2X1_LOC_392/Y 0.14fF
C953 NOR2X1_LOC_65/B NOR2X1_LOC_318/B 0.72fF
C954 NOR2X1_LOC_792/B NAND2X1_LOC_198/B 0.02fF
C955 NOR2X1_LOC_292/Y NOR2X1_LOC_717/A 0.03fF
C956 NOR2X1_LOC_620/Y INVX1_LOC_132/A 0.06fF
C957 INVX1_LOC_2/A INVX1_LOC_72/A 0.14fF
C958 INVX1_LOC_58/A NOR2X1_LOC_737/a_36_216# 0.00fF
C959 INVX1_LOC_77/Y D_INPUT_5 0.09fF
C960 NAND2X1_LOC_59/B INVX1_LOC_77/A 0.22fF
C961 NAND2X1_LOC_321/a_36_24# NOR2X1_LOC_325/A 0.00fF
C962 NOR2X1_LOC_456/Y INVX1_LOC_206/Y 0.07fF
C963 NAND2X1_LOC_860/A INVX1_LOC_286/A 1.66fF
C964 NAND2X1_LOC_208/B INVX1_LOC_25/Y 0.42fF
C965 INVX1_LOC_262/Y INVX1_LOC_92/A 0.03fF
C966 NOR2X1_LOC_160/B INVX1_LOC_137/Y 0.01fF
C967 INVX1_LOC_118/A INVX1_LOC_284/A 0.00fF
C968 NOR2X1_LOC_226/A INVX1_LOC_72/A 0.10fF
C969 NOR2X1_LOC_65/B INVX1_LOC_93/Y 0.09fF
C970 NOR2X1_LOC_211/a_36_216# INVX1_LOC_286/A 0.02fF
C971 NOR2X1_LOC_45/B INVX1_LOC_57/A 0.51fF
C972 INVX1_LOC_95/A NAND2X1_LOC_286/B 0.03fF
C973 NOR2X1_LOC_51/A INPUT_7 0.04fF
C974 NAND2X1_LOC_66/a_36_24# INVX1_LOC_136/A 0.01fF
C975 D_INPUT_0 NOR2X1_LOC_103/Y 0.07fF
C976 NOR2X1_LOC_82/A NOR2X1_LOC_332/A 0.48fF
C977 INVX1_LOC_58/A NOR2X1_LOC_78/A 0.03fF
C978 NAND2X1_LOC_341/A NOR2X1_LOC_658/Y 0.04fF
C979 NOR2X1_LOC_433/A NAND2X1_LOC_799/Y 0.01fF
C980 NOR2X1_LOC_711/Y NOR2X1_LOC_383/B 0.15fF
C981 NAND2X1_LOC_72/Y INVX1_LOC_69/Y 0.02fF
C982 INVX1_LOC_30/A INVX1_LOC_232/A 0.17fF
C983 INVX1_LOC_104/A NOR2X1_LOC_550/B 0.18fF
C984 NAND2X1_LOC_721/A INVX1_LOC_78/A 0.03fF
C985 NOR2X1_LOC_218/Y INVX1_LOC_72/A 0.05fF
C986 INVX1_LOC_223/Y INPUT_0 0.03fF
C987 NAND2X1_LOC_579/A NOR2X1_LOC_19/B 0.16fF
C988 NOR2X1_LOC_516/B NOR2X1_LOC_703/B 0.03fF
C989 INVX1_LOC_279/A INVX1_LOC_81/Y 0.01fF
C990 NOR2X1_LOC_456/Y NOR2X1_LOC_600/Y 0.01fF
C991 VDD INVX1_LOC_116/Y 0.71fF
C992 NOR2X1_LOC_615/a_36_216# NAND2X1_LOC_866/B 0.00fF
C993 NOR2X1_LOC_78/B NOR2X1_LOC_106/Y 0.24fF
C994 NAND2X1_LOC_733/B NAND2X1_LOC_866/A 0.02fF
C995 NAND2X1_LOC_860/A INVX1_LOC_95/A 0.03fF
C996 NAND2X1_LOC_206/Y NAND2X1_LOC_219/B 0.04fF
C997 NOR2X1_LOC_860/B NOR2X1_LOC_346/B 0.09fF
C998 INVX1_LOC_49/A INVX1_LOC_192/Y 0.02fF
C999 INVX1_LOC_255/Y NOR2X1_LOC_68/A 0.00fF
C1000 NOR2X1_LOC_705/B INVX1_LOC_90/A 0.03fF
C1001 INVX1_LOC_11/A NAND2X1_LOC_654/B 0.03fF
C1002 NAND2X1_LOC_338/B INVX1_LOC_49/A 0.09fF
C1003 NOR2X1_LOC_189/A INVX1_LOC_280/Y 0.01fF
C1004 INVX1_LOC_30/A NOR2X1_LOC_366/Y 0.02fF
C1005 INVX1_LOC_124/Y NOR2X1_LOC_123/B 0.63fF
C1006 NOR2X1_LOC_419/Y INVX1_LOC_218/A 0.01fF
C1007 INVX1_LOC_136/A INVX1_LOC_227/A 0.10fF
C1008 NOR2X1_LOC_360/Y NOR2X1_LOC_665/A 0.20fF
C1009 INVX1_LOC_45/A D_INPUT_0 0.25fF
C1010 NOR2X1_LOC_781/a_36_216# INVX1_LOC_72/A 0.00fF
C1011 INVX1_LOC_287/Y VDD 0.27fF
C1012 NAND2X1_LOC_323/B INVX1_LOC_49/A 0.18fF
C1013 NOR2X1_LOC_447/B NOR2X1_LOC_677/Y 0.05fF
C1014 NAND2X1_LOC_53/Y NOR2X1_LOC_163/Y 0.00fF
C1015 NOR2X1_LOC_577/Y NAND2X1_LOC_840/B 0.02fF
C1016 NOR2X1_LOC_15/Y INVX1_LOC_100/A 0.01fF
C1017 INVX1_LOC_25/A VDD 1.90fF
C1018 NAND2X1_LOC_86/Y INVX1_LOC_50/Y 0.01fF
C1019 INVX1_LOC_233/Y NOR2X1_LOC_253/Y 0.01fF
C1020 NOR2X1_LOC_632/Y NOR2X1_LOC_208/Y 0.02fF
C1021 INVX1_LOC_44/A NOR2X1_LOC_727/B 0.01fF
C1022 NOR2X1_LOC_209/Y NOR2X1_LOC_731/A 0.48fF
C1023 NAND2X1_LOC_338/B INVX1_LOC_60/A 0.04fF
C1024 INVX1_LOC_5/A NOR2X1_LOC_124/a_36_216# 0.00fF
C1025 INVX1_LOC_64/A NOR2X1_LOC_682/a_36_216# 0.00fF
C1026 INVX1_LOC_72/A NAND2X1_LOC_648/A 0.05fF
C1027 INVX1_LOC_5/A INVX1_LOC_112/A 0.02fF
C1028 INVX1_LOC_5/A INVX1_LOC_59/Y 0.11fF
C1029 INVX1_LOC_305/A NOR2X1_LOC_174/B 0.03fF
C1030 INVX1_LOC_72/A INPUT_1 0.07fF
C1031 INVX1_LOC_64/A NOR2X1_LOC_857/A 0.07fF
C1032 INVX1_LOC_106/Y INVX1_LOC_19/A 0.03fF
C1033 INVX1_LOC_89/A INVX1_LOC_72/Y 0.00fF
C1034 INVX1_LOC_34/A INVX1_LOC_25/Y 0.21fF
C1035 INVX1_LOC_45/A NOR2X1_LOC_216/a_36_216# 0.00fF
C1036 NOR2X1_LOC_91/Y NOR2X1_LOC_76/A 0.06fF
C1037 INVX1_LOC_78/A INVX1_LOC_117/Y 0.03fF
C1038 NAND2X1_LOC_579/A NOR2X1_LOC_528/Y 0.02fF
C1039 INVX1_LOC_34/A NAND2X1_LOC_716/a_36_24# 0.00fF
C1040 INVX1_LOC_124/Y INVX1_LOC_102/Y 0.15fF
C1041 NAND2X1_LOC_785/A NAND2X1_LOC_850/Y 0.28fF
C1042 INVX1_LOC_5/A INVX1_LOC_176/A 0.03fF
C1043 INVX1_LOC_2/A NAND2X1_LOC_338/B 0.22fF
C1044 NOR2X1_LOC_655/B INVX1_LOC_54/Y 0.01fF
C1045 D_INPUT_0 INVX1_LOC_71/A 0.07fF
C1046 NOR2X1_LOC_12/a_36_216# NOR2X1_LOC_11/Y 0.00fF
C1047 NOR2X1_LOC_226/A NAND2X1_LOC_633/a_36_24# 0.01fF
C1048 NOR2X1_LOC_598/B NAND2X1_LOC_96/A 0.75fF
C1049 NOR2X1_LOC_68/A NOR2X1_LOC_644/A 0.01fF
C1050 NAND2X1_LOC_740/Y INVX1_LOC_20/A 0.03fF
C1051 NOR2X1_LOC_599/Y INPUT_0 0.29fF
C1052 NAND2X1_LOC_114/B INVX1_LOC_92/Y 0.05fF
C1053 INVX1_LOC_51/A NAND2X1_LOC_96/A 0.03fF
C1054 NAND2X1_LOC_717/Y NOR2X1_LOC_526/Y 0.10fF
C1055 INVX1_LOC_290/Y INVX1_LOC_272/A 0.02fF
C1056 INVX1_LOC_279/A NOR2X1_LOC_344/A 0.02fF
C1057 NOR2X1_LOC_798/A NOR2X1_LOC_853/a_36_216# 0.00fF
C1058 INVX1_LOC_45/A NAND2X1_LOC_538/a_36_24# 0.01fF
C1059 INVX1_LOC_291/A NOR2X1_LOC_65/Y 0.02fF
C1060 NAND2X1_LOC_647/B NOR2X1_LOC_814/A 0.20fF
C1061 NAND2X1_LOC_848/A NAND2X1_LOC_793/B 0.01fF
C1062 NAND2X1_LOC_347/B INVX1_LOC_95/Y 0.01fF
C1063 NOR2X1_LOC_68/A NOR2X1_LOC_828/B 0.07fF
C1064 NOR2X1_LOC_254/A INVX1_LOC_78/Y 0.01fF
C1065 NOR2X1_LOC_383/B NOR2X1_LOC_801/a_36_216# 0.00fF
C1066 INVX1_LOC_23/A NOR2X1_LOC_729/A 0.23fF
C1067 NOR2X1_LOC_160/B NOR2X1_LOC_114/A 0.02fF
C1068 NOR2X1_LOC_794/B NOR2X1_LOC_337/Y 0.03fF
C1069 INVX1_LOC_96/Y INVX1_LOC_22/A 0.07fF
C1070 NOR2X1_LOC_215/A INVX1_LOC_139/A 0.01fF
C1071 NOR2X1_LOC_383/B INVX1_LOC_307/A 0.10fF
C1072 NAND2X1_LOC_550/A INVX1_LOC_91/A 0.07fF
C1073 INVX1_LOC_1/A NAND2X1_LOC_659/B 0.00fF
C1074 NOR2X1_LOC_858/A NOR2X1_LOC_676/a_36_216# 0.03fF
C1075 NOR2X1_LOC_78/Y NAND2X1_LOC_215/A 0.04fF
C1076 NAND2X1_LOC_860/A INVX1_LOC_54/A 0.15fF
C1077 INVX1_LOC_49/A INVX1_LOC_313/Y 0.03fF
C1078 NOR2X1_LOC_216/a_36_216# INVX1_LOC_71/A 0.00fF
C1079 INVX1_LOC_93/A NOR2X1_LOC_176/Y 0.01fF
C1080 NOR2X1_LOC_160/B INVX1_LOC_91/A 5.76fF
C1081 INVX1_LOC_224/Y INVX1_LOC_46/Y 0.11fF
C1082 INVX1_LOC_121/A INVX1_LOC_257/Y 0.03fF
C1083 NAND2X1_LOC_740/Y NOR2X1_LOC_765/Y 0.00fF
C1084 NOR2X1_LOC_383/B NOR2X1_LOC_445/B 0.03fF
C1085 INVX1_LOC_57/A NOR2X1_LOC_862/B 0.10fF
C1086 INVX1_LOC_90/A NOR2X1_LOC_172/Y 0.03fF
C1087 NOR2X1_LOC_788/B NOR2X1_LOC_804/B 0.03fF
C1088 NOR2X1_LOC_394/Y NAND2X1_LOC_773/B 0.06fF
C1089 INVX1_LOC_182/A NOR2X1_LOC_303/Y 0.10fF
C1090 INVX1_LOC_90/A NOR2X1_LOC_772/Y 0.07fF
C1091 NOR2X1_LOC_753/Y NAND2X1_LOC_807/Y 0.07fF
C1092 NOR2X1_LOC_218/A NOR2X1_LOC_657/B 0.23fF
C1093 NAND2X1_LOC_167/a_36_24# INPUT_0 0.01fF
C1094 NOR2X1_LOC_457/A NAND2X1_LOC_447/Y 0.19fF
C1095 INVX1_LOC_90/A NOR2X1_LOC_147/B 0.01fF
C1096 NOR2X1_LOC_389/B NOR2X1_LOC_772/Y 0.02fF
C1097 NAND2X1_LOC_623/a_36_24# INVX1_LOC_118/A 0.00fF
C1098 INVX1_LOC_43/A INVX1_LOC_137/A 0.15fF
C1099 NOR2X1_LOC_67/A NAND2X1_LOC_859/Y 0.30fF
C1100 INVX1_LOC_1/A VDD 3.00fF
C1101 NOR2X1_LOC_52/B NAND2X1_LOC_660/a_36_24# 0.00fF
C1102 INVX1_LOC_90/A NOR2X1_LOC_392/B 0.01fF
C1103 NAND2X1_LOC_725/a_36_24# NOR2X1_LOC_298/Y 0.09fF
C1104 NOR2X1_LOC_246/a_36_216# NOR2X1_LOC_309/Y 0.00fF
C1105 NAND2X1_LOC_325/Y NAND2X1_LOC_807/Y 0.02fF
C1106 INVX1_LOC_45/A NOR2X1_LOC_191/a_36_216# 0.01fF
C1107 NOR2X1_LOC_742/A INVX1_LOC_113/Y 0.04fF
C1108 INVX1_LOC_94/Y INVX1_LOC_29/A 0.21fF
C1109 NOR2X1_LOC_389/B NOR2X1_LOC_392/B 0.10fF
C1110 INVX1_LOC_89/A INVX1_LOC_266/Y 0.03fF
C1111 NOR2X1_LOC_784/Y VDD 0.24fF
C1112 INVX1_LOC_182/A NOR2X1_LOC_254/Y 0.01fF
C1113 INVX1_LOC_19/Y INVX1_LOC_15/A 0.06fF
C1114 NAND2X1_LOC_21/Y NAND2X1_LOC_51/B 0.48fF
C1115 INVX1_LOC_118/A NOR2X1_LOC_384/A 0.00fF
C1116 INVX1_LOC_19/A NOR2X1_LOC_635/B 0.09fF
C1117 INVX1_LOC_2/A INVX1_LOC_313/Y 0.07fF
C1118 INVX1_LOC_34/A INVX1_LOC_75/A 0.15fF
C1119 INVX1_LOC_277/A NOR2X1_LOC_209/A 0.02fF
C1120 INVX1_LOC_277/Y NOR2X1_LOC_711/Y 0.33fF
C1121 NOR2X1_LOC_794/B VDD 0.42fF
C1122 INVX1_LOC_279/A NOR2X1_LOC_540/a_36_216# 0.00fF
C1123 NOR2X1_LOC_246/Y NAND2X1_LOC_342/Y 0.19fF
C1124 INVX1_LOC_87/A INVX1_LOC_42/A 0.03fF
C1125 NAND2X1_LOC_338/B INPUT_1 0.46fF
C1126 INVX1_LOC_35/A NAND2X1_LOC_574/A 0.02fF
C1127 INVX1_LOC_30/A NAND2X1_LOC_447/Y 2.28fF
C1128 INVX1_LOC_19/A INVX1_LOC_275/Y 0.06fF
C1129 NOR2X1_LOC_90/a_36_216# INVX1_LOC_59/Y 0.01fF
C1130 NOR2X1_LOC_735/Y INVX1_LOC_96/Y 0.12fF
C1131 NAND2X1_LOC_198/B NOR2X1_LOC_269/Y 0.38fF
C1132 NOR2X1_LOC_388/Y NOR2X1_LOC_74/A 0.13fF
C1133 INVX1_LOC_19/A NOR2X1_LOC_748/A 0.56fF
C1134 INVX1_LOC_159/A NOR2X1_LOC_43/Y 0.01fF
C1135 INVX1_LOC_181/A INVX1_LOC_29/A 0.07fF
C1136 INVX1_LOC_106/Y INVX1_LOC_26/Y 0.03fF
C1137 INVX1_LOC_161/Y NOR2X1_LOC_816/Y 0.06fF
C1138 INVX1_LOC_296/A INVX1_LOC_29/A 0.08fF
C1139 NOR2X1_LOC_488/Y NAND2X1_LOC_862/Y 0.26fF
C1140 NOR2X1_LOC_576/B INVX1_LOC_22/A 0.06fF
C1141 NOR2X1_LOC_341/a_36_216# NOR2X1_LOC_78/A 0.00fF
C1142 NAND2X1_LOC_807/B NAND2X1_LOC_286/B 0.00fF
C1143 INVX1_LOC_88/A INVX1_LOC_9/A 0.10fF
C1144 INVX1_LOC_86/Y NOR2X1_LOC_550/B 0.02fF
C1145 INVX1_LOC_12/A NOR2X1_LOC_383/B 0.13fF
C1146 NAND2X1_LOC_74/B NOR2X1_LOC_441/a_36_216# 0.02fF
C1147 INVX1_LOC_17/A INVX1_LOC_118/Y 0.08fF
C1148 INVX1_LOC_45/A NOR2X1_LOC_266/B 0.03fF
C1149 NAND2X1_LOC_785/A INVX1_LOC_282/A 0.03fF
C1150 NAND2X1_LOC_537/Y INVX1_LOC_54/A 0.68fF
C1151 INVX1_LOC_50/A NOR2X1_LOC_89/A 1.27fF
C1152 NAND2X1_LOC_149/Y NOR2X1_LOC_156/Y 0.06fF
C1153 NAND2X1_LOC_357/B NAND2X1_LOC_858/B 0.07fF
C1154 INVX1_LOC_28/A NAND2X1_LOC_862/A 0.04fF
C1155 INVX1_LOC_72/A NOR2X1_LOC_586/Y 0.20fF
C1156 NOR2X1_LOC_136/Y NOR2X1_LOC_329/B 0.06fF
C1157 NOR2X1_LOC_392/Y NOR2X1_LOC_84/B 0.00fF
C1158 NOR2X1_LOC_384/Y VDD 0.91fF
C1159 INVX1_LOC_17/Y NAND2X1_LOC_254/Y 0.01fF
C1160 INVX1_LOC_278/Y INVX1_LOC_140/A 0.10fF
C1161 NOR2X1_LOC_584/Y INVX1_LOC_23/A 0.03fF
C1162 NOR2X1_LOC_464/B NOR2X1_LOC_155/A 0.01fF
C1163 NOR2X1_LOC_454/Y INVX1_LOC_107/Y 0.07fF
C1164 NAND2X1_LOC_312/a_36_24# NOR2X1_LOC_862/B 0.06fF
C1165 INVX1_LOC_133/Y INVX1_LOC_6/A 0.06fF
C1166 INVX1_LOC_78/A INVX1_LOC_87/A 0.03fF
C1167 NAND2X1_LOC_729/Y VDD 0.01fF
C1168 NOR2X1_LOC_720/B NOR2X1_LOC_557/A 0.21fF
C1169 NOR2X1_LOC_468/Y NOR2X1_LOC_179/a_36_216# 0.00fF
C1170 INVX1_LOC_45/A NAND2X1_LOC_848/A 0.03fF
C1171 NOR2X1_LOC_473/B NAND2X1_LOC_656/Y 0.42fF
C1172 INVX1_LOC_208/A INVX1_LOC_79/A 0.10fF
C1173 INVX1_LOC_206/A NOR2X1_LOC_501/B 0.01fF
C1174 NAND2X1_LOC_785/B INVX1_LOC_38/A 0.66fF
C1175 INVX1_LOC_17/A NAND2X1_LOC_244/a_36_24# 0.00fF
C1176 NAND2X1_LOC_544/a_36_24# NOR2X1_LOC_89/A 0.00fF
C1177 NOR2X1_LOC_103/Y INVX1_LOC_46/Y 0.02fF
C1178 NOR2X1_LOC_577/Y NOR2X1_LOC_137/a_36_216# 0.01fF
C1179 NOR2X1_LOC_52/B INVX1_LOC_159/Y 0.01fF
C1180 NAND2X1_LOC_53/Y INVX1_LOC_179/A 0.48fF
C1181 NAND2X1_LOC_9/Y NOR2X1_LOC_38/a_36_216# 0.00fF
C1182 INVX1_LOC_64/A INVX1_LOC_109/Y 0.31fF
C1183 INVX1_LOC_36/A NAND2X1_LOC_297/a_36_24# 0.01fF
C1184 INPUT_0 INVX1_LOC_25/Y 0.21fF
C1185 INVX1_LOC_5/A NOR2X1_LOC_340/A 0.03fF
C1186 INVX1_LOC_135/A NOR2X1_LOC_356/A 0.07fF
C1187 NAND2X1_LOC_67/Y NOR2X1_LOC_66/Y 0.16fF
C1188 INVX1_LOC_18/A NOR2X1_LOC_684/Y 0.31fF
C1189 INVX1_LOC_189/A INVX1_LOC_91/A 0.00fF
C1190 NOR2X1_LOC_65/B INVX1_LOC_87/A 0.02fF
C1191 INVX1_LOC_278/A INVX1_LOC_19/Y 0.03fF
C1192 INVX1_LOC_72/A INVX1_LOC_118/A 0.21fF
C1193 NOR2X1_LOC_360/Y NOR2X1_LOC_652/a_36_216# 0.01fF
C1194 INVX1_LOC_32/A NOR2X1_LOC_678/A 0.03fF
C1195 INVX1_LOC_90/A NOR2X1_LOC_389/B 0.07fF
C1196 NAND2X1_LOC_500/a_36_24# INVX1_LOC_91/A 0.00fF
C1197 NOR2X1_LOC_389/A NOR2X1_LOC_831/B 0.10fF
C1198 NOR2X1_LOC_409/B INVX1_LOC_296/Y 0.03fF
C1199 NOR2X1_LOC_15/Y INVX1_LOC_186/Y 0.07fF
C1200 INVX1_LOC_34/A NAND2X1_LOC_453/A 0.03fF
C1201 NOR2X1_LOC_690/A INVX1_LOC_46/A 0.07fF
C1202 INVX1_LOC_39/A INVX1_LOC_284/A 0.44fF
C1203 NOR2X1_LOC_717/Y INVX1_LOC_92/A 0.06fF
C1204 INVX1_LOC_71/A NAND2X1_LOC_848/A 0.10fF
C1205 INVX1_LOC_132/A INVX1_LOC_117/A 0.47fF
C1206 INVX1_LOC_48/Y NAND2X1_LOC_81/B 0.02fF
C1207 NOR2X1_LOC_140/a_36_216# D_INPUT_3 0.00fF
C1208 NOR2X1_LOC_657/B NOR2X1_LOC_131/A 0.01fF
C1209 INVX1_LOC_208/A INVX1_LOC_91/A 0.03fF
C1210 NOR2X1_LOC_160/B NOR2X1_LOC_179/Y 0.01fF
C1211 INVX1_LOC_135/A NOR2X1_LOC_74/A 0.10fF
C1212 NAND2X1_LOC_184/a_36_24# NOR2X1_LOC_356/A 0.00fF
C1213 NOR2X1_LOC_194/Y INVX1_LOC_46/A 0.01fF
C1214 INVX1_LOC_174/A INVX1_LOC_84/A 0.09fF
C1215 INVX1_LOC_299/A INVX1_LOC_29/A 0.68fF
C1216 NOR2X1_LOC_639/Y NOR2X1_LOC_654/A 0.08fF
C1217 INVX1_LOC_26/Y NOR2X1_LOC_748/A 0.46fF
C1218 NAND2X1_LOC_550/A INVX1_LOC_203/A 0.09fF
C1219 INVX1_LOC_90/A NAND2X1_LOC_348/A 0.08fF
C1220 NOR2X1_LOC_130/A NOR2X1_LOC_815/A 0.01fF
C1221 NOR2X1_LOC_91/A NAND2X1_LOC_787/Y 0.00fF
C1222 NAND2X1_LOC_853/Y INVX1_LOC_11/Y 0.03fF
C1223 INVX1_LOC_303/A INVX1_LOC_9/A 0.41fF
C1224 NOR2X1_LOC_663/A NAND2X1_LOC_618/Y 0.01fF
C1225 NOR2X1_LOC_172/Y INVX1_LOC_38/A 0.03fF
C1226 NOR2X1_LOC_288/A INVX1_LOC_117/A 0.15fF
C1227 INVX1_LOC_61/A NAND2X1_LOC_243/B 0.11fF
C1228 INVX1_LOC_289/Y INVX1_LOC_42/A 0.03fF
C1229 NOR2X1_LOC_561/Y NOR2X1_LOC_139/Y 0.00fF
C1230 NAND2X1_LOC_390/A NAND2X1_LOC_642/Y 0.78fF
C1231 NAND2X1_LOC_149/Y D_INPUT_5 0.07fF
C1232 NAND2X1_LOC_84/Y INVX1_LOC_92/A 3.06fF
C1233 INVX1_LOC_75/A INVX1_LOC_131/A 0.63fF
C1234 NAND2X1_LOC_537/Y NOR2X1_LOC_48/B 0.07fF
C1235 NOR2X1_LOC_329/B INVX1_LOC_144/A 0.14fF
C1236 NOR2X1_LOC_82/A NOR2X1_LOC_847/A 0.32fF
C1237 INVX1_LOC_50/A NAND2X1_LOC_804/A 0.01fF
C1238 NOR2X1_LOC_152/Y INVX1_LOC_117/Y 0.03fF
C1239 NAND2X1_LOC_133/a_36_24# INVX1_LOC_91/A 0.00fF
C1240 NOR2X1_LOC_209/Y INVX1_LOC_117/A 1.27fF
C1241 NOR2X1_LOC_638/a_36_216# INVX1_LOC_92/A 0.02fF
C1242 INVX1_LOC_89/A INVX1_LOC_125/Y 0.08fF
C1243 NAND2X1_LOC_193/a_36_24# INVX1_LOC_117/Y 0.00fF
C1244 NOR2X1_LOC_309/Y NOR2X1_LOC_186/a_36_216# 0.00fF
C1245 NOR2X1_LOC_82/A INVX1_LOC_42/A 0.14fF
C1246 NOR2X1_LOC_791/B INVX1_LOC_3/A 0.00fF
C1247 NOR2X1_LOC_561/Y NAND2X1_LOC_468/B 0.01fF
C1248 INVX1_LOC_75/A INPUT_0 0.89fF
C1249 INVX1_LOC_192/A NAND2X1_LOC_93/B 0.05fF
C1250 NAND2X1_LOC_721/A NAND2X1_LOC_859/B 0.27fF
C1251 NAND2X1_LOC_528/a_36_24# NAND2X1_LOC_96/A 0.00fF
C1252 NOR2X1_LOC_721/Y NOR2X1_LOC_188/A 0.02fF
C1253 INVX1_LOC_72/A NAND2X1_LOC_63/Y 0.06fF
C1254 NOR2X1_LOC_298/Y INVX1_LOC_76/A 0.20fF
C1255 NAND2X1_LOC_181/Y NOR2X1_LOC_271/Y 0.01fF
C1256 INVX1_LOC_289/Y INVX1_LOC_78/A 0.03fF
C1257 NOR2X1_LOC_552/A NOR2X1_LOC_356/A -0.02fF
C1258 NOR2X1_LOC_721/Y NOR2X1_LOC_548/B 0.03fF
C1259 NAND2X1_LOC_500/Y INVX1_LOC_42/A 0.01fF
C1260 INVX1_LOC_192/A NAND2X1_LOC_425/Y 0.23fF
C1261 NOR2X1_LOC_203/Y INVX1_LOC_9/A 0.03fF
C1262 NAND2X1_LOC_338/B INVX1_LOC_118/A 0.01fF
C1263 NOR2X1_LOC_295/Y NOR2X1_LOC_831/B 0.02fF
C1264 INVX1_LOC_174/A INVX1_LOC_15/A 0.08fF
C1265 NOR2X1_LOC_715/a_36_216# NOR2X1_LOC_78/A 0.02fF
C1266 NOR2X1_LOC_191/a_36_216# INVX1_LOC_102/Y 0.00fF
C1267 NOR2X1_LOC_794/A NOR2X1_LOC_74/A 0.02fF
C1268 NOR2X1_LOC_226/A NOR2X1_LOC_506/Y 0.72fF
C1269 INVX1_LOC_254/Y NOR2X1_LOC_68/a_36_216# 0.00fF
C1270 INVX1_LOC_153/A INVX1_LOC_84/A 0.01fF
C1271 NOR2X1_LOC_706/A INVX1_LOC_91/A 0.44fF
C1272 INVX1_LOC_298/Y INVX1_LOC_299/A 0.07fF
C1273 NOR2X1_LOC_767/a_36_216# NAND2X1_LOC_93/B 0.01fF
C1274 NOR2X1_LOC_123/B NOR2X1_LOC_266/B 0.19fF
C1275 NAND2X1_LOC_228/a_36_24# INVX1_LOC_38/A 0.01fF
C1276 INVX1_LOC_35/A NAND2X1_LOC_35/Y 0.08fF
C1277 NAND2X1_LOC_799/A INVX1_LOC_273/A 0.03fF
C1278 INVX1_LOC_111/Y INVX1_LOC_92/A 0.10fF
C1279 NOR2X1_LOC_82/A INVX1_LOC_78/A 0.15fF
C1280 INVX1_LOC_61/A INVX1_LOC_284/A 0.05fF
C1281 INVX1_LOC_21/A D_INPUT_1 0.03fF
C1282 NAND2X1_LOC_751/a_36_24# NAND2X1_LOC_214/B 0.00fF
C1283 NAND2X1_LOC_124/a_36_24# NOR2X1_LOC_269/Y 0.00fF
C1284 NOR2X1_LOC_590/A NAND2X1_LOC_647/B 0.02fF
C1285 NAND2X1_LOC_672/B NOR2X1_LOC_655/Y 0.25fF
C1286 NOR2X1_LOC_717/B NAND2X1_LOC_472/Y 0.40fF
C1287 NAND2X1_LOC_660/Y NOR2X1_LOC_331/B 0.07fF
C1288 NAND2X1_LOC_861/Y NAND2X1_LOC_721/A 0.07fF
C1289 INVX1_LOC_222/Y NOR2X1_LOC_598/B 0.01fF
C1290 NOR2X1_LOC_577/Y INVX1_LOC_49/Y 0.10fF
C1291 NOR2X1_LOC_512/a_36_216# INVX1_LOC_38/A 0.00fF
C1292 NOR2X1_LOC_168/A NOR2X1_LOC_445/B 0.01fF
C1293 NOR2X1_LOC_552/A NOR2X1_LOC_74/A 0.07fF
C1294 INVX1_LOC_143/A NAND2X1_LOC_572/B 0.00fF
C1295 NAND2X1_LOC_632/B INVX1_LOC_12/A 0.04fF
C1296 INVX1_LOC_58/A NAND2X1_LOC_724/A 0.06fF
C1297 INVX1_LOC_224/A INVX1_LOC_50/A 0.00fF
C1298 NOR2X1_LOC_65/B NOR2X1_LOC_82/A 0.12fF
C1299 NAND2X1_LOC_342/Y INVX1_LOC_285/A 0.01fF
C1300 INVX1_LOC_305/A NOR2X1_LOC_623/B 0.07fF
C1301 NOR2X1_LOC_32/B INVX1_LOC_237/A 0.11fF
C1302 INVX1_LOC_59/A NAND2X1_LOC_549/Y 0.02fF
C1303 INVX1_LOC_102/Y NOR2X1_LOC_266/B 0.20fF
C1304 NOR2X1_LOC_495/Y NAND2X1_LOC_254/Y 0.23fF
C1305 INVX1_LOC_50/A INVX1_LOC_11/A 0.13fF
C1306 INVX1_LOC_90/A NAND2X1_LOC_849/B 0.05fF
C1307 INVX1_LOC_162/A INVX1_LOC_29/A 0.25fF
C1308 NOR2X1_LOC_254/A NOR2X1_LOC_727/B 0.09fF
C1309 INVX1_LOC_14/A INVX1_LOC_53/A 0.00fF
C1310 INVX1_LOC_79/A NAND2X1_LOC_211/Y 0.46fF
C1311 NOR2X1_LOC_411/A NAND2X1_LOC_725/B 0.00fF
C1312 INVX1_LOC_90/A INVX1_LOC_38/A 1.36fF
C1313 NOR2X1_LOC_218/A INVX1_LOC_271/A 0.05fF
C1314 INVX1_LOC_64/A NAND2X1_LOC_706/Y 0.04fF
C1315 INVX1_LOC_96/Y INVX1_LOC_186/Y 0.06fF
C1316 INVX1_LOC_21/A NOR2X1_LOC_652/Y 0.07fF
C1317 NAND2X1_LOC_68/a_36_24# INVX1_LOC_5/A 0.00fF
C1318 NAND2X1_LOC_660/Y NOR2X1_LOC_592/B 0.06fF
C1319 NOR2X1_LOC_441/Y NAND2X1_LOC_286/B 0.31fF
C1320 INVX1_LOC_299/A NAND2X1_LOC_385/a_36_24# 0.00fF
C1321 INVX1_LOC_18/A INVX1_LOC_273/A 0.03fF
C1322 NOR2X1_LOC_315/Y INVX1_LOC_29/A 0.03fF
C1323 NAND2X1_LOC_672/B INVX1_LOC_3/A 0.02fF
C1324 INVX1_LOC_90/A NOR2X1_LOC_96/Y 0.14fF
C1325 NOR2X1_LOC_84/Y NAND2X1_LOC_81/B 0.03fF
C1326 NOR2X1_LOC_74/A INVX1_LOC_139/Y 0.03fF
C1327 NOR2X1_LOC_418/Y INVX1_LOC_84/A 0.02fF
C1328 NOR2X1_LOC_151/Y NAND2X1_LOC_472/Y 0.04fF
C1329 NAND2X1_LOC_514/Y INVX1_LOC_78/A 0.01fF
C1330 NOR2X1_LOC_188/A VDD 1.59fF
C1331 INVX1_LOC_58/A NOR2X1_LOC_45/Y 0.03fF
C1332 NOR2X1_LOC_435/a_36_216# INVX1_LOC_103/A 0.00fF
C1333 NOR2X1_LOC_837/Y NOR2X1_LOC_839/B 0.14fF
C1334 INVX1_LOC_34/A INVX1_LOC_283/A 0.03fF
C1335 INVX1_LOC_24/A NOR2X1_LOC_394/Y 0.26fF
C1336 NOR2X1_LOC_548/B VDD 1.82fF
C1337 NOR2X1_LOC_537/Y NAND2X1_LOC_63/Y 0.03fF
C1338 NAND2X1_LOC_338/B NAND2X1_LOC_63/Y 0.10fF
C1339 NAND2X1_LOC_738/B NAND2X1_LOC_733/Y 0.05fF
C1340 NAND2X1_LOC_579/A INVX1_LOC_93/A 0.10fF
C1341 NOR2X1_LOC_68/A INVX1_LOC_16/Y 0.01fF
C1342 NOR2X1_LOC_350/A INVX1_LOC_4/Y 0.00fF
C1343 INVX1_LOC_5/A INVX1_LOC_103/A 0.10fF
C1344 NOR2X1_LOC_427/Y INVX1_LOC_77/Y 0.07fF
C1345 INVX1_LOC_10/Y NOR2X1_LOC_74/A 0.03fF
C1346 NAND2X1_LOC_198/B INVX1_LOC_26/A 0.03fF
C1347 NAND2X1_LOC_348/A INVX1_LOC_38/A 0.01fF
C1348 INVX1_LOC_264/Y INVX1_LOC_20/A 0.01fF
C1349 NOR2X1_LOC_92/Y NAND2X1_LOC_714/B 0.07fF
C1350 INVX1_LOC_2/A NOR2X1_LOC_226/Y 0.01fF
C1351 INVX1_LOC_191/Y NOR2X1_LOC_584/Y 0.01fF
C1352 INVX1_LOC_58/A INVX1_LOC_170/A 0.11fF
C1353 INVX1_LOC_25/Y NOR2X1_LOC_84/B 0.00fF
C1354 NAND2X1_LOC_655/A INVX1_LOC_76/A 0.10fF
C1355 INVX1_LOC_135/A NOR2X1_LOC_243/B 0.07fF
C1356 INVX1_LOC_91/A NAND2X1_LOC_211/Y 0.01fF
C1357 NOR2X1_LOC_84/A NOR2X1_LOC_28/a_36_216# 0.00fF
C1358 INVX1_LOC_161/Y NOR2X1_LOC_304/Y 0.04fF
C1359 NOR2X1_LOC_91/A INVX1_LOC_181/Y 0.17fF
C1360 NOR2X1_LOC_223/B INVX1_LOC_174/A 0.01fF
C1361 NOR2X1_LOC_590/A NOR2X1_LOC_109/a_36_216# 0.00fF
C1362 INVX1_LOC_103/A INVX1_LOC_178/A 0.09fF
C1363 INVX1_LOC_5/A INVX1_LOC_292/A 0.07fF
C1364 NOR2X1_LOC_68/A NAND2X1_LOC_205/A 0.38fF
C1365 VDD NOR2X1_LOC_43/Y 0.13fF
C1366 NOR2X1_LOC_302/Y INVX1_LOC_179/A 0.01fF
C1367 INVX1_LOC_268/Y INVX1_LOC_29/A 0.09fF
C1368 NOR2X1_LOC_329/B NOR2X1_LOC_155/A 0.07fF
C1369 NOR2X1_LOC_860/B NOR2X1_LOC_843/B 0.07fF
C1370 NOR2X1_LOC_560/A NOR2X1_LOC_243/B 0.16fF
C1371 NAND2X1_LOC_661/A INVX1_LOC_117/Y 0.01fF
C1372 NAND2X1_LOC_468/B INVX1_LOC_76/A 0.05fF
C1373 INVX1_LOC_269/A NOR2X1_LOC_140/A 0.07fF
C1374 INVX1_LOC_24/A NOR2X1_LOC_654/A 0.01fF
C1375 INVX1_LOC_171/A INVX1_LOC_84/A 0.03fF
C1376 NAND2X1_LOC_332/Y INVX1_LOC_78/A 0.05fF
C1377 INVX1_LOC_177/A NOR2X1_LOC_801/B 0.27fF
C1378 NOR2X1_LOC_246/Y INVX1_LOC_285/A 0.02fF
C1379 INVX1_LOC_227/Y INVX1_LOC_53/A 0.01fF
C1380 NOR2X1_LOC_99/B NOR2X1_LOC_721/B 0.04fF
C1381 INVX1_LOC_181/Y INVX1_LOC_23/A 0.07fF
C1382 NOR2X1_LOC_431/Y INVX1_LOC_271/A 0.01fF
C1383 NOR2X1_LOC_85/a_36_216# INVX1_LOC_284/A 0.00fF
C1384 INVX1_LOC_150/A INVX1_LOC_19/A 0.02fF
C1385 NOR2X1_LOC_191/A INVX1_LOC_32/A 0.01fF
C1386 NAND2X1_LOC_642/Y INVX1_LOC_117/A 0.04fF
C1387 INVX1_LOC_50/A NOR2X1_LOC_433/A 0.13fF
C1388 NOR2X1_LOC_599/A NOR2X1_LOC_304/Y 0.20fF
C1389 NOR2X1_LOC_598/B NAND2X1_LOC_656/A 0.17fF
C1390 NOR2X1_LOC_181/A NAND2X1_LOC_472/Y 0.01fF
C1391 INVX1_LOC_24/A INVX1_LOC_58/Y 0.07fF
C1392 NAND2X1_LOC_375/a_36_24# INVX1_LOC_174/A 0.00fF
C1393 INVX1_LOC_89/A INVX1_LOC_19/A 15.63fF
C1394 INVX1_LOC_149/A NAND2X1_LOC_72/B 0.06fF
C1395 NOR2X1_LOC_131/Y INVX1_LOC_15/A 0.04fF
C1396 INVX1_LOC_50/A NOR2X1_LOC_593/Y 0.09fF
C1397 INVX1_LOC_289/Y NOR2X1_LOC_503/Y 0.10fF
C1398 NOR2X1_LOC_332/A NOR2X1_LOC_340/A 0.07fF
C1399 NAND2X1_LOC_162/A NOR2X1_LOC_467/A 0.08fF
C1400 INVX1_LOC_58/A INVX1_LOC_132/A 0.08fF
C1401 NAND2X1_LOC_9/Y INVX1_LOC_254/A 0.03fF
C1402 INVX1_LOC_82/Y INVX1_LOC_3/A 0.22fF
C1403 INVX1_LOC_278/A NAND2X1_LOC_169/a_36_24# 0.00fF
C1404 NAND2X1_LOC_214/Y INVX1_LOC_31/A 0.05fF
C1405 NOR2X1_LOC_261/Y INVX1_LOC_153/A 0.12fF
C1406 INVX1_LOC_86/Y INVX1_LOC_75/Y 0.08fF
C1407 INVX1_LOC_306/A INVX1_LOC_42/A 0.01fF
C1408 NOR2X1_LOC_589/A INVX1_LOC_15/A 0.06fF
C1409 NAND2X1_LOC_684/a_36_24# INVX1_LOC_78/A 0.01fF
C1410 INVX1_LOC_286/Y NAND2X1_LOC_326/A 0.00fF
C1411 INVX1_LOC_224/Y INVX1_LOC_60/A 0.20fF
C1412 INVX1_LOC_41/A NOR2X1_LOC_456/Y 0.01fF
C1413 INVX1_LOC_50/A NOR2X1_LOC_52/B 1.24fF
C1414 INVX1_LOC_58/A INVX1_LOC_225/A 0.11fF
C1415 INVX1_LOC_226/Y INVX1_LOC_165/A 0.01fF
C1416 NOR2X1_LOC_134/Y NOR2X1_LOC_103/Y 0.01fF
C1417 NAND2X1_LOC_563/Y INVX1_LOC_23/A 0.04fF
C1418 INVX1_LOC_11/A INVX1_LOC_61/Y 0.07fF
C1419 GATE_741 INVX1_LOC_300/Y 0.01fF
C1420 INVX1_LOC_267/A INVX1_LOC_166/A 0.03fF
C1421 INVX1_LOC_268/A NOR2X1_LOC_158/Y 0.05fF
C1422 INVX1_LOC_247/A INVX1_LOC_274/A 0.06fF
C1423 NAND2X1_LOC_72/Y NOR2X1_LOC_593/Y 1.10fF
C1424 INVX1_LOC_2/A INVX1_LOC_224/Y 0.03fF
C1425 INVX1_LOC_256/A INVX1_LOC_130/A 0.01fF
C1426 INVX1_LOC_227/A NAND2X1_LOC_647/B 0.04fF
C1427 NAND2X1_LOC_354/Y NAND2X1_LOC_175/a_36_24# 0.00fF
C1428 NOR2X1_LOC_15/Y INVX1_LOC_18/A 0.38fF
C1429 INVX1_LOC_53/Y INVX1_LOC_26/A 0.07fF
C1430 NOR2X1_LOC_163/Y INVX1_LOC_12/A 0.02fF
C1431 NOR2X1_LOC_389/A NAND2X1_LOC_352/B 0.28fF
C1432 INVX1_LOC_35/A NAND2X1_LOC_465/Y 0.09fF
C1433 NAND2X1_LOC_728/Y NOR2X1_LOC_15/Y 0.07fF
C1434 INVX1_LOC_45/A NAND2X1_LOC_30/Y 0.03fF
C1435 INVX1_LOC_21/A NOR2X1_LOC_607/Y 0.01fF
C1436 NOR2X1_LOC_619/A INVX1_LOC_26/A 0.01fF
C1437 NOR2X1_LOC_598/B NOR2X1_LOC_423/Y 0.23fF
C1438 NOR2X1_LOC_778/B NOR2X1_LOC_858/A 0.00fF
C1439 INVX1_LOC_57/Y INVX1_LOC_200/A 0.10fF
C1440 NOR2X1_LOC_733/Y INVX1_LOC_186/Y 0.02fF
C1441 INVX1_LOC_117/A NOR2X1_LOC_271/Y 0.02fF
C1442 INVX1_LOC_111/Y INVX1_LOC_53/A 0.01fF
C1443 INVX1_LOC_2/A NAND2X1_LOC_793/B 0.07fF
C1444 NOR2X1_LOC_82/A NOR2X1_LOC_554/B 0.09fF
C1445 NOR2X1_LOC_703/Y INVX1_LOC_19/A 0.09fF
C1446 NAND2X1_LOC_112/Y NOR2X1_LOC_135/a_36_216# 0.00fF
C1447 INVX1_LOC_5/A INVX1_LOC_240/A 0.10fF
C1448 INPUT_6 NAND2X1_LOC_11/Y 0.03fF
C1449 INVX1_LOC_284/Y NAND2X1_LOC_733/A 0.48fF
C1450 NAND2X1_LOC_561/B NAND2X1_LOC_837/Y 0.03fF
C1451 INVX1_LOC_233/Y NOR2X1_LOC_482/Y 0.01fF
C1452 INVX1_LOC_91/A NOR2X1_LOC_605/A 0.01fF
C1453 NOR2X1_LOC_111/A INVX1_LOC_185/A 0.01fF
C1454 INVX1_LOC_1/A INVX1_LOC_184/Y 0.04fF
C1455 NOR2X1_LOC_598/B NOR2X1_LOC_222/Y 0.07fF
C1456 NOR2X1_LOC_226/A NAND2X1_LOC_793/B 0.14fF
C1457 NAND2X1_LOC_391/Y NAND2X1_LOC_569/A 0.07fF
C1458 NOR2X1_LOC_88/Y INVX1_LOC_20/A 0.39fF
C1459 INVX1_LOC_289/Y NOR2X1_LOC_152/Y 0.07fF
C1460 NOR2X1_LOC_15/Y INVX1_LOC_172/A 0.03fF
C1461 NOR2X1_LOC_87/B INVX1_LOC_38/Y 0.12fF
C1462 INVX1_LOC_90/A NAND2X1_LOC_223/A 0.03fF
C1463 INVX1_LOC_6/A NOR2X1_LOC_584/Y 0.11fF
C1464 NAND2X1_LOC_773/a_36_24# INVX1_LOC_306/A 0.00fF
C1465 INVX1_LOC_237/Y NAND2X1_LOC_725/B 0.11fF
C1466 NOR2X1_LOC_75/Y INVX1_LOC_24/A 0.00fF
C1467 NAND2X1_LOC_182/A NAND2X1_LOC_793/a_36_24# 0.00fF
C1468 NOR2X1_LOC_740/Y INVX1_LOC_77/A 0.07fF
C1469 NOR2X1_LOC_45/Y NOR2X1_LOC_338/Y 0.01fF
C1470 NOR2X1_LOC_363/Y NAND2X1_LOC_93/B 0.79fF
C1471 INVX1_LOC_251/Y INVX1_LOC_306/Y 0.01fF
C1472 INVX1_LOC_256/A INVX1_LOC_81/A 0.03fF
C1473 INVX1_LOC_1/A INVX1_LOC_153/Y 0.29fF
C1474 NOR2X1_LOC_66/Y INVX1_LOC_76/A 0.02fF
C1475 INVX1_LOC_295/A NAND2X1_LOC_425/a_36_24# 0.01fF
C1476 INVX1_LOC_89/A INVX1_LOC_26/Y 0.17fF
C1477 INVX1_LOC_84/A INVX1_LOC_20/A 0.19fF
C1478 NOR2X1_LOC_51/A INVX1_LOC_38/A 5.07fF
C1479 NAND2X1_LOC_190/Y NOR2X1_LOC_344/A 0.15fF
C1480 NOR2X1_LOC_790/B NOR2X1_LOC_548/Y 0.00fF
C1481 INVX1_LOC_150/Y INVX1_LOC_77/A 0.20fF
C1482 NAND2X1_LOC_36/a_36_24# NAND2X1_LOC_36/A 0.00fF
C1483 NAND2X1_LOC_581/Y INVX1_LOC_1/A 0.02fF
C1484 NOR2X1_LOC_506/Y INVX1_LOC_118/A 0.01fF
C1485 INVX1_LOC_2/Y INVX1_LOC_3/A 0.05fF
C1486 NAND2X1_LOC_11/a_36_24# D_INPUT_6 0.00fF
C1487 NOR2X1_LOC_355/A INVX1_LOC_270/Y 0.07fF
C1488 INVX1_LOC_1/A INVX1_LOC_121/Y 0.01fF
C1489 INVX1_LOC_166/A INVX1_LOC_89/A 0.98fF
C1490 NAND2X1_LOC_715/B NOR2X1_LOC_269/a_36_216# 0.00fF
C1491 NAND2X1_LOC_348/A NAND2X1_LOC_223/A 0.03fF
C1492 INVX1_LOC_25/A NAND2X1_LOC_143/a_36_24# 0.00fF
C1493 NOR2X1_LOC_32/B INVX1_LOC_234/A 0.28fF
C1494 INVX1_LOC_64/A NOR2X1_LOC_32/Y 0.00fF
C1495 NAND2X1_LOC_149/Y NAND2X1_LOC_451/Y 0.13fF
C1496 INVX1_LOC_161/A NOR2X1_LOC_577/Y 0.18fF
C1497 NOR2X1_LOC_705/B INVX1_LOC_33/A 0.01fF
C1498 NAND2X1_LOC_21/Y INVX1_LOC_174/A 0.05fF
C1499 INVX1_LOC_224/Y INPUT_1 0.14fF
C1500 INVX1_LOC_89/A NAND2X1_LOC_265/a_36_24# 0.00fF
C1501 INVX1_LOC_269/A NOR2X1_LOC_709/A 0.10fF
C1502 NAND2X1_LOC_276/Y NOR2X1_LOC_160/B 0.08fF
C1503 INVX1_LOC_274/A NOR2X1_LOC_676/Y 0.01fF
C1504 NOR2X1_LOC_137/A INVX1_LOC_53/A 0.01fF
C1505 NOR2X1_LOC_305/Y INVX1_LOC_264/A 0.01fF
C1506 NOR2X1_LOC_15/Y NOR2X1_LOC_709/a_36_216# 0.00fF
C1507 VDD NOR2X1_LOC_810/Y 0.09fF
C1508 NOR2X1_LOC_658/Y NOR2X1_LOC_219/a_36_216# 0.01fF
C1509 INVX1_LOC_59/Y NOR2X1_LOC_847/A 0.01fF
C1510 INVX1_LOC_119/A INVX1_LOC_161/Y 0.03fF
C1511 INVX1_LOC_45/A INVX1_LOC_49/A 0.26fF
C1512 NOR2X1_LOC_536/A NOR2X1_LOC_485/Y 0.02fF
C1513 NOR2X1_LOC_816/A INVX1_LOC_240/A 0.14fF
C1514 NAND2X1_LOC_833/Y INVX1_LOC_141/Y 0.02fF
C1515 NAND2X1_LOC_563/A NOR2X1_LOC_140/A 0.07fF
C1516 INVX1_LOC_256/A NOR2X1_LOC_802/A 0.03fF
C1517 NOR2X1_LOC_78/B INVX1_LOC_14/A 0.08fF
C1518 INVX1_LOC_59/Y INVX1_LOC_42/A 3.04fF
C1519 INVX1_LOC_124/A INVX1_LOC_150/Y 0.23fF
C1520 INVX1_LOC_2/A NOR2X1_LOC_103/Y 0.10fF
C1521 INPUT_1 NAND2X1_LOC_793/B 0.07fF
C1522 NOR2X1_LOC_209/Y NOR2X1_LOC_738/Y 0.02fF
C1523 INVX1_LOC_13/Y INVX1_LOC_7/A 0.01fF
C1524 NOR2X1_LOC_425/Y NOR2X1_LOC_11/Y 0.01fF
C1525 INVX1_LOC_179/A INVX1_LOC_307/A 0.04fF
C1526 INVX1_LOC_110/Y NAND2X1_LOC_116/A 0.74fF
C1527 NOR2X1_LOC_48/Y INVX1_LOC_117/A 0.02fF
C1528 INVX1_LOC_232/Y INVX1_LOC_216/Y 0.01fF
C1529 NOR2X1_LOC_794/B INVX1_LOC_177/A 0.55fF
C1530 NAND2X1_LOC_563/Y INVX1_LOC_31/A 0.70fF
C1531 INVX1_LOC_5/A INVX1_LOC_120/A 0.03fF
C1532 NOR2X1_LOC_32/B NOR2X1_LOC_19/B 0.07fF
C1533 NAND2X1_LOC_550/A NAND2X1_LOC_374/Y 1.30fF
C1534 NAND2X1_LOC_96/A INVX1_LOC_29/A 0.07fF
C1535 INVX1_LOC_21/A NOR2X1_LOC_747/a_36_216# 0.02fF
C1536 INVX1_LOC_24/A NOR2X1_LOC_419/Y 0.69fF
C1537 NOR2X1_LOC_666/A NOR2X1_LOC_665/A 0.01fF
C1538 NOR2X1_LOC_590/A NAND2X1_LOC_342/Y 0.02fF
C1539 INVX1_LOC_20/A INVX1_LOC_15/A 14.58fF
C1540 INVX1_LOC_24/A NOR2X1_LOC_716/B 0.07fF
C1541 NOR2X1_LOC_588/A NOR2X1_LOC_25/Y 0.01fF
C1542 INVX1_LOC_304/Y INVX1_LOC_57/Y 0.03fF
C1543 INVX1_LOC_49/A INVX1_LOC_71/A 0.23fF
C1544 INVX1_LOC_136/A INVX1_LOC_104/A 0.18fF
C1545 NOR2X1_LOC_659/a_36_216# NOR2X1_LOC_52/B 0.00fF
C1546 NOR2X1_LOC_376/A INVX1_LOC_83/A 0.03fF
C1547 INVX1_LOC_14/A NAND2X1_LOC_392/Y 0.03fF
C1548 NOR2X1_LOC_735/a_36_216# INVX1_LOC_63/Y 0.01fF
C1549 NOR2X1_LOC_635/A INVX1_LOC_18/A 0.01fF
C1550 NAND2X1_LOC_330/a_36_24# INVX1_LOC_49/A 0.00fF
C1551 INVX1_LOC_1/A NOR2X1_LOC_785/Y 0.04fF
C1552 INVX1_LOC_2/A INVX1_LOC_45/A 0.13fF
C1553 NOR2X1_LOC_315/Y NAND2X1_LOC_634/Y 0.06fF
C1554 NOR2X1_LOC_457/B INVX1_LOC_88/Y 0.01fF
C1555 NOR2X1_LOC_336/B NOR2X1_LOC_538/Y 0.00fF
C1556 NOR2X1_LOC_119/a_36_216# NAND2X1_LOC_74/B 0.00fF
C1557 INVX1_LOC_14/A NOR2X1_LOC_459/A 0.07fF
C1558 INVX1_LOC_88/A NOR2X1_LOC_561/Y 0.48fF
C1559 NAND2X1_LOC_361/Y INVX1_LOC_314/Y 0.08fF
C1560 INVX1_LOC_2/A NOR2X1_LOC_568/A 0.10fF
C1561 INVX1_LOC_276/A INVX1_LOC_36/A 0.07fF
C1562 INVX1_LOC_35/A INVX1_LOC_144/A 2.75fF
C1563 NOR2X1_LOC_78/B NOR2X1_LOC_717/Y 0.11fF
C1564 NOR2X1_LOC_846/B NAND2X1_LOC_473/A 0.03fF
C1565 NOR2X1_LOC_433/A NOR2X1_LOC_679/B 0.01fF
C1566 INVX1_LOC_45/A NOR2X1_LOC_226/A 0.11fF
C1567 INVX1_LOC_14/A INVX1_LOC_83/A 0.18fF
C1568 NAND2X1_LOC_765/a_36_24# INVX1_LOC_18/A 0.00fF
C1569 NOR2X1_LOC_67/A INVX1_LOC_36/A 0.07fF
C1570 NAND2X1_LOC_454/a_36_24# NAND2X1_LOC_454/Y 0.02fF
C1571 INVX1_LOC_179/Y NOR2X1_LOC_500/B 0.05fF
C1572 NAND2X1_LOC_332/Y NOR2X1_LOC_152/Y 0.03fF
C1573 INVX1_LOC_41/A NOR2X1_LOC_550/B 0.01fF
C1574 NAND2X1_LOC_567/Y NAND2X1_LOC_354/B 0.03fF
C1575 INVX1_LOC_285/A INVX1_LOC_265/Y 0.00fF
C1576 INVX1_LOC_34/A NOR2X1_LOC_577/Y 0.14fF
C1577 NOR2X1_LOC_172/Y INVX1_LOC_33/A 0.01fF
C1578 INVX1_LOC_26/A NAND2X1_LOC_465/A 0.00fF
C1579 INVX1_LOC_285/A NOR2X1_LOC_814/A 0.00fF
C1580 NAND2X1_LOC_785/A INVX1_LOC_41/Y 0.03fF
C1581 NOR2X1_LOC_147/B INVX1_LOC_33/A 0.01fF
C1582 NOR2X1_LOC_355/B NOR2X1_LOC_717/A 0.23fF
C1583 INVX1_LOC_3/Y NOR2X1_LOC_271/Y 0.00fF
C1584 INVX1_LOC_50/A NOR2X1_LOC_601/Y 0.05fF
C1585 NAND2X1_LOC_783/Y NAND2X1_LOC_783/A 0.02fF
C1586 INVX1_LOC_2/A INVX1_LOC_71/A 0.12fF
C1587 NOR2X1_LOC_392/B INVX1_LOC_33/A 0.01fF
C1588 INVX1_LOC_12/A INVX1_LOC_179/A 0.05fF
C1589 INVX1_LOC_26/Y NOR2X1_LOC_852/a_36_216# 0.00fF
C1590 NOR2X1_LOC_103/Y INPUT_1 0.07fF
C1591 NAND2X1_LOC_363/B NOR2X1_LOC_78/A 0.07fF
C1592 NOR2X1_LOC_203/a_36_216# INVX1_LOC_206/Y 0.00fF
C1593 INVX1_LOC_72/Y INVX1_LOC_25/Y 0.00fF
C1594 NOR2X1_LOC_226/A INVX1_LOC_71/A 1.33fF
C1595 INVX1_LOC_72/A NAND2X1_LOC_735/B 0.03fF
C1596 NOR2X1_LOC_833/Y INVX1_LOC_23/A 0.01fF
C1597 INVX1_LOC_64/A INVX1_LOC_264/Y 0.01fF
C1598 INVX1_LOC_278/Y NAND2X1_LOC_520/a_36_24# 0.00fF
C1599 NOR2X1_LOC_360/Y INVX1_LOC_16/A 0.01fF
C1600 NAND2X1_LOC_231/Y NOR2X1_LOC_577/Y 0.10fF
C1601 NOR2X1_LOC_315/Y INVX1_LOC_8/A 0.07fF
C1602 INVX1_LOC_103/A INVX1_LOC_140/A 0.10fF
C1603 INVX1_LOC_72/A INPUT_5 1.36fF
C1604 NOR2X1_LOC_716/B INVX1_LOC_143/A 0.33fF
C1605 NAND2X1_LOC_717/Y INVX1_LOC_207/A 0.01fF
C1606 INVX1_LOC_118/Y INVX1_LOC_94/Y 0.08fF
C1607 NOR2X1_LOC_791/Y INVX1_LOC_98/A 0.13fF
C1608 NAND2X1_LOC_725/Y VDD 4.53fF
C1609 NOR2X1_LOC_218/Y INVX1_LOC_71/A 0.04fF
C1610 INVX1_LOC_57/Y NAND2X1_LOC_808/A 0.00fF
C1611 NAND2X1_LOC_59/B INVX1_LOC_243/A 0.02fF
C1612 NOR2X1_LOC_78/a_36_216# NOR2X1_LOC_38/B 0.00fF
C1613 INVX1_LOC_94/A NOR2X1_LOC_188/Y 0.00fF
C1614 NAND2X1_LOC_454/Y INVX1_LOC_54/A 0.07fF
C1615 INVX1_LOC_1/A INVX1_LOC_285/Y 0.08fF
C1616 INVX1_LOC_278/A INVX1_LOC_20/A 0.08fF
C1617 NOR2X1_LOC_617/Y NOR2X1_LOC_86/A 0.02fF
C1618 INVX1_LOC_45/A INPUT_1 0.10fF
C1619 INVX1_LOC_152/Y INVX1_LOC_176/A 0.02fF
C1620 INVX1_LOC_225/Y INVX1_LOC_75/A 0.01fF
C1621 INVX1_LOC_45/Y INVX1_LOC_10/A 0.01fF
C1622 INVX1_LOC_38/A NAND2X1_LOC_256/a_36_24# 0.01fF
C1623 INVX1_LOC_64/A NOR2X1_LOC_825/Y 0.01fF
C1624 NOR2X1_LOC_717/a_36_216# INVX1_LOC_16/A 0.00fF
C1625 NOR2X1_LOC_717/B INVX1_LOC_24/A 0.03fF
C1626 NAND2X1_LOC_276/Y NOR2X1_LOC_516/B 0.18fF
C1627 NOR2X1_LOC_392/B INVX1_LOC_40/A 0.08fF
C1628 INVX1_LOC_248/A NOR2X1_LOC_591/Y 0.03fF
C1629 NAND2X1_LOC_740/A INVX1_LOC_10/A 0.01fF
C1630 INVX1_LOC_34/A INVX1_LOC_22/A 0.89fF
C1631 NOR2X1_LOC_536/A INVX1_LOC_29/Y 0.03fF
C1632 NOR2X1_LOC_570/B NOR2X1_LOC_570/Y 0.05fF
C1633 INVX1_LOC_145/A NAND2X1_LOC_331/a_36_24# 0.00fF
C1634 INVX1_LOC_13/Y INVX1_LOC_76/A 0.15fF
C1635 INVX1_LOC_84/A INVX1_LOC_4/A 1.48fF
C1636 INVX1_LOC_224/Y INVX1_LOC_118/A 0.08fF
C1637 NAND2X1_LOC_500/a_36_24# NAND2X1_LOC_374/Y 0.01fF
C1638 INVX1_LOC_1/A INVX1_LOC_65/A 0.02fF
C1639 INVX1_LOC_71/A INPUT_1 0.35fF
C1640 NOR2X1_LOC_716/B NOR2X1_LOC_130/A 0.07fF
C1641 INVX1_LOC_1/A INVX1_LOC_316/A 0.19fF
C1642 NOR2X1_LOC_690/A NOR2X1_LOC_700/Y 0.06fF
C1643 NOR2X1_LOC_383/B INVX1_LOC_92/A 0.10fF
C1644 INVX1_LOC_204/Y INVX1_LOC_117/A 0.03fF
C1645 INVX1_LOC_14/A NOR2X1_LOC_368/Y 0.01fF
C1646 NOR2X1_LOC_503/A INVX1_LOC_24/A 0.01fF
C1647 INVX1_LOC_202/A NOR2X1_LOC_122/Y 0.04fF
C1648 INVX1_LOC_256/A NOR2X1_LOC_192/A 0.01fF
C1649 NAND2X1_LOC_231/Y INVX1_LOC_22/A 0.01fF
C1650 NAND2X1_LOC_793/B INVX1_LOC_118/A 0.01fF
C1651 NOR2X1_LOC_810/A NOR2X1_LOC_802/A 0.10fF
C1652 NAND2X1_LOC_93/B INVX1_LOC_29/Y 0.05fF
C1653 INVX1_LOC_90/A INVX1_LOC_33/A 0.14fF
C1654 INVX1_LOC_24/A NOR2X1_LOC_151/Y 0.03fF
C1655 NOR2X1_LOC_440/Y NOR2X1_LOC_767/a_36_216# 0.00fF
C1656 NAND2X1_LOC_326/A VDD 0.08fF
C1657 NOR2X1_LOC_389/B INVX1_LOC_33/A 0.07fF
C1658 NOR2X1_LOC_433/A NAND2X1_LOC_652/Y 0.02fF
C1659 INVX1_LOC_88/A INVX1_LOC_76/A 0.07fF
C1660 NAND2X1_LOC_198/B NOR2X1_LOC_368/A 0.16fF
C1661 INVX1_LOC_136/A INVX1_LOC_206/Y 0.03fF
C1662 NOR2X1_LOC_705/B NOR2X1_LOC_486/Y 0.00fF
C1663 INVX1_LOC_14/A INVX1_LOC_46/A 0.30fF
C1664 NOR2X1_LOC_103/Y NAND2X1_LOC_455/a_36_24# 0.00fF
C1665 INVX1_LOC_49/A INVX1_LOC_102/Y 0.15fF
C1666 INVX1_LOC_17/A INVX1_LOC_36/Y 0.18fF
C1667 NAND2X1_LOC_392/A NAND2X1_LOC_390/a_36_24# 0.02fF
C1668 NAND2X1_LOC_218/B INPUT_0 0.07fF
C1669 INVX1_LOC_34/A NOR2X1_LOC_735/Y 0.00fF
C1670 INVX1_LOC_30/A NOR2X1_LOC_78/A 0.19fF
C1671 INVX1_LOC_58/Y NOR2X1_LOC_197/B 0.10fF
C1672 INVX1_LOC_181/Y INVX1_LOC_6/A 0.21fF
C1673 INVX1_LOC_35/A NOR2X1_LOC_155/A 1.08fF
C1674 NAND2X1_LOC_656/A INVX1_LOC_201/A 0.04fF
C1675 NOR2X1_LOC_795/Y NOR2X1_LOC_356/A 0.10fF
C1676 NAND2X1_LOC_785/A NAND2X1_LOC_865/a_36_24# 0.00fF
C1677 NOR2X1_LOC_226/A NOR2X1_LOC_123/B 1.48fF
C1678 INVX1_LOC_64/A NOR2X1_LOC_88/Y 0.07fF
C1679 NOR2X1_LOC_577/Y INPUT_0 0.07fF
C1680 VDD NAND2X1_LOC_807/A -0.00fF
C1681 NAND2X1_LOC_698/a_36_24# NAND2X1_LOC_474/Y 0.01fF
C1682 INVX1_LOC_81/Y NAND2X1_LOC_469/B 0.01fF
C1683 INVX1_LOC_53/A NOR2X1_LOC_127/Y 0.07fF
C1684 INVX1_LOC_21/A NOR2X1_LOC_61/Y 0.21fF
C1685 INVX1_LOC_245/Y INVX1_LOC_139/Y 0.02fF
C1686 INVX1_LOC_15/A INVX1_LOC_4/A 0.07fF
C1687 NOR2X1_LOC_808/A INVX1_LOC_196/Y 0.01fF
C1688 INVX1_LOC_29/A NAND2X1_LOC_99/A 0.07fF
C1689 INVX1_LOC_102/A NOR2X1_LOC_301/A 0.07fF
C1690 INVX1_LOC_90/A NAND2X1_LOC_798/A 0.02fF
C1691 NOR2X1_LOC_329/B NAND2X1_LOC_660/A 0.09fF
C1692 INVX1_LOC_72/A NAND2X1_LOC_212/Y 0.57fF
C1693 INVX1_LOC_30/A NAND2X1_LOC_464/A 0.03fF
C1694 NOR2X1_LOC_804/B NOR2X1_LOC_551/Y 0.03fF
C1695 INVX1_LOC_90/A INVX1_LOC_40/A 0.00fF
C1696 INVX1_LOC_64/A INVX1_LOC_84/A 1.89fF
C1697 INVX1_LOC_75/A INVX1_LOC_266/Y 0.10fF
C1698 INVX1_LOC_41/A NOR2X1_LOC_334/A 0.03fF
C1699 INVX1_LOC_277/A VDD 0.00fF
C1700 NOR2X1_LOC_763/A INVX1_LOC_92/A 0.02fF
C1701 NOR2X1_LOC_644/B NAND2X1_LOC_472/Y 0.05fF
C1702 NOR2X1_LOC_614/Y NOR2X1_LOC_356/A 0.02fF
C1703 INVX1_LOC_36/A NOR2X1_LOC_558/A 0.00fF
C1704 INVX1_LOC_236/Y INVX1_LOC_33/Y 0.00fF
C1705 NOR2X1_LOC_852/A VDD 0.24fF
C1706 NOR2X1_LOC_192/a_36_216# INVX1_LOC_6/A 0.00fF
C1707 NOR2X1_LOC_392/Y INVX1_LOC_19/A 0.07fF
C1708 NAND2X1_LOC_361/Y NOR2X1_LOC_557/A 0.16fF
C1709 NOR2X1_LOC_103/Y INVX1_LOC_118/A 0.14fF
C1710 INVX1_LOC_224/Y NAND2X1_LOC_455/B 0.06fF
C1711 INVX1_LOC_50/A NAND2X1_LOC_254/Y 0.01fF
C1712 INVX1_LOC_251/Y NOR2X1_LOC_74/A 0.01fF
C1713 INVX1_LOC_177/A NOR2X1_LOC_188/A 0.00fF
C1714 INVX1_LOC_155/A INVX1_LOC_91/A 0.21fF
C1715 NOR2X1_LOC_590/A NOR2X1_LOC_862/a_36_216# 0.00fF
C1716 INVX1_LOC_289/Y NAND2X1_LOC_802/Y 0.39fF
C1717 INVX1_LOC_5/A NOR2X1_LOC_631/A 0.03fF
C1718 NOR2X1_LOC_577/Y NAND2X1_LOC_649/B 0.01fF
C1719 NOR2X1_LOC_186/Y NAND2X1_LOC_475/Y 0.02fF
C1720 INVX1_LOC_69/Y NOR2X1_LOC_802/A 0.02fF
C1721 INVX1_LOC_135/A D_INPUT_0 0.17fF
C1722 NOR2X1_LOC_453/a_36_216# NAND2X1_LOC_425/Y 0.01fF
C1723 NOR2X1_LOC_681/a_36_216# NAND2X1_LOC_175/Y 0.00fF
C1724 NOR2X1_LOC_807/B INVX1_LOC_307/Y 0.04fF
C1725 INVX1_LOC_229/A NOR2X1_LOC_491/Y 0.02fF
C1726 INVX1_LOC_30/A NOR2X1_LOC_60/Y 0.00fF
C1727 INVX1_LOC_23/A NOR2X1_LOC_114/Y 0.02fF
C1728 INVX1_LOC_251/Y NOR2X1_LOC_9/Y 0.15fF
C1729 NAND2X1_LOC_348/A INVX1_LOC_40/A 0.03fF
C1730 INVX1_LOC_120/A NOR2X1_LOC_332/A 0.03fF
C1731 NOR2X1_LOC_826/Y INVX1_LOC_284/A 0.04fF
C1732 INPUT_0 NOR2X1_LOC_346/B 0.00fF
C1733 INVX1_LOC_116/Y INVX1_LOC_4/Y 0.09fF
C1734 NOR2X1_LOC_758/Y NOR2X1_LOC_405/A 0.03fF
C1735 NOR2X1_LOC_130/A NOR2X1_LOC_130/Y 0.02fF
C1736 INVX1_LOC_35/A NOR2X1_LOC_833/B 0.23fF
C1737 NAND2X1_LOC_84/Y INVX1_LOC_46/A 0.01fF
C1738 D_INPUT_0 NOR2X1_LOC_560/A -0.00fF
C1739 INVX1_LOC_223/Y INVX1_LOC_19/A 0.03fF
C1740 NOR2X1_LOC_632/Y NOR2X1_LOC_742/A 0.02fF
C1741 NOR2X1_LOC_598/B NOR2X1_LOC_477/B 0.04fF
C1742 NOR2X1_LOC_123/B INPUT_1 0.12fF
C1743 NAND2X1_LOC_802/A NAND2X1_LOC_453/A 0.06fF
C1744 INVX1_LOC_45/A INVX1_LOC_118/A 0.11fF
C1745 INPUT_0 INVX1_LOC_22/A 0.16fF
C1746 NOR2X1_LOC_625/Y VDD 0.23fF
C1747 INVX1_LOC_5/A NAND2X1_LOC_469/a_36_24# 0.00fF
C1748 NAND2X1_LOC_661/B INVX1_LOC_91/A 0.01fF
C1749 NOR2X1_LOC_151/Y NOR2X1_LOC_739/a_36_216# 0.00fF
C1750 INVX1_LOC_73/A NAND2X1_LOC_656/Y 0.03fF
C1751 INVX1_LOC_25/A INVX1_LOC_4/Y 0.03fF
C1752 INVX1_LOC_239/A INVX1_LOC_163/Y 0.13fF
C1753 INVX1_LOC_227/A INVX1_LOC_67/Y 0.13fF
C1754 D_INPUT_1 NOR2X1_LOC_248/A 0.04fF
C1755 NOR2X1_LOC_380/A NAND2X1_LOC_560/A 4.66fF
C1756 NAND2X1_LOC_61/Y NOR2X1_LOC_65/Y 0.00fF
C1757 INVX1_LOC_64/A INVX1_LOC_15/A 0.54fF
C1758 NOR2X1_LOC_68/A INVX1_LOC_54/A 0.14fF
C1759 NOR2X1_LOC_301/A NOR2X1_LOC_280/a_36_216# 0.01fF
C1760 NOR2X1_LOC_92/Y NAND2X1_LOC_74/B 0.57fF
C1761 INVX1_LOC_102/Y INPUT_1 0.00fF
C1762 INVX1_LOC_168/A INVX1_LOC_76/A 0.19fF
C1763 NOR2X1_LOC_590/A INVX1_LOC_285/A 0.00fF
C1764 INVX1_LOC_33/A NOR2X1_LOC_561/A 0.01fF
C1765 NOR2X1_LOC_300/Y VDD 0.22fF
C1766 INVX1_LOC_71/A INVX1_LOC_118/A 0.33fF
C1767 INVX1_LOC_49/A NOR2X1_LOC_331/B 0.07fF
C1768 VDD NOR2X1_LOC_87/B 0.38fF
C1769 D_INPUT_0 NOR2X1_LOC_391/B 0.00fF
C1770 NAND2X1_LOC_96/A INVX1_LOC_8/A 0.13fF
C1771 INVX1_LOC_14/A NOR2X1_LOC_671/Y 0.02fF
C1772 NAND2X1_LOC_799/A INVX1_LOC_49/Y 0.07fF
C1773 NOR2X1_LOC_590/A NOR2X1_LOC_814/A 0.32fF
C1774 NOR2X1_LOC_538/Y NOR2X1_LOC_857/A 0.01fF
C1775 NOR2X1_LOC_860/B NOR2X1_LOC_860/Y 0.00fF
C1776 INVX1_LOC_33/A INVX1_LOC_38/A 0.22fF
C1777 NOR2X1_LOC_324/A NOR2X1_LOC_325/A 0.47fF
C1778 INVX1_LOC_111/Y INVX1_LOC_46/A 0.01fF
C1779 INVX1_LOC_77/A NOR2X1_LOC_612/Y 0.00fF
C1780 NAND2X1_LOC_360/B VDD 0.15fF
C1781 INVX1_LOC_12/Y NOR2X1_LOC_709/A 0.10fF
C1782 NOR2X1_LOC_532/Y INVX1_LOC_69/Y 0.03fF
C1783 INVX1_LOC_308/A NAND2X1_LOC_286/B 0.01fF
C1784 NOR2X1_LOC_140/A NOR2X1_LOC_554/A 0.06fF
C1785 NOR2X1_LOC_652/Y NOR2X1_LOC_248/A 0.03fF
C1786 NOR2X1_LOC_160/B INVX1_LOC_125/A 0.01fF
C1787 INVX1_LOC_17/A INVX1_LOC_102/A 0.07fF
C1788 INVX1_LOC_60/Y NOR2X1_LOC_536/A 0.07fF
C1789 INVX1_LOC_103/A INVX1_LOC_42/A 0.03fF
C1790 INVX1_LOC_13/A INVX1_LOC_95/Y 0.06fF
C1791 INVX1_LOC_53/A NOR2X1_LOC_383/B 0.77fF
C1792 NOR2X1_LOC_103/Y NAND2X1_LOC_455/B 0.09fF
C1793 NAND2X1_LOC_397/a_36_24# INVX1_LOC_15/A 0.00fF
C1794 NOR2X1_LOC_165/Y VDD 0.35fF
C1795 NOR2X1_LOC_510/Y NOR2X1_LOC_338/a_36_216# 0.01fF
C1796 INVX1_LOC_49/A NOR2X1_LOC_592/B 0.03fF
C1797 NAND2X1_LOC_577/A INVX1_LOC_29/A 0.06fF
C1798 NOR2X1_LOC_722/Y INVX1_LOC_186/Y 0.03fF
C1799 INVX1_LOC_2/A NOR2X1_LOC_331/B 0.17fF
C1800 INVX1_LOC_34/A NOR2X1_LOC_88/A 0.00fF
C1801 INVX1_LOC_292/A INVX1_LOC_42/A 1.20fF
C1802 INVX1_LOC_255/Y INVX1_LOC_178/Y 0.04fF
C1803 NOR2X1_LOC_716/B NOR2X1_LOC_197/B 0.00fF
C1804 NOR2X1_LOC_537/Y INVX1_LOC_230/A 0.05fF
C1805 INVX1_LOC_174/Y VDD 0.40fF
C1806 NOR2X1_LOC_180/Y INVX1_LOC_274/A 0.33fF
C1807 INVX1_LOC_1/A INVX1_LOC_4/Y 0.03fF
C1808 NOR2X1_LOC_87/B NOR2X1_LOC_846/a_36_216# 0.00fF
C1809 NOR2X1_LOC_246/A INVX1_LOC_95/Y 0.08fF
C1810 GATE_479 INVX1_LOC_37/A 0.01fF
C1811 INVX1_LOC_61/Y NAND2X1_LOC_254/Y 0.07fF
C1812 INVX1_LOC_21/A NOR2X1_LOC_318/A 0.04fF
C1813 NOR2X1_LOC_226/A NOR2X1_LOC_331/B 0.18fF
C1814 INVX1_LOC_124/A NOR2X1_LOC_612/Y 0.02fF
C1815 INVX1_LOC_18/A INVX1_LOC_49/Y 0.03fF
C1816 INVX1_LOC_36/Y NOR2X1_LOC_199/B 0.01fF
C1817 INVX1_LOC_35/A NOR2X1_LOC_598/B 0.22fF
C1818 INPUT_0 INVX1_LOC_100/A 0.04fF
C1819 INVX1_LOC_269/A NOR2X1_LOC_334/Y 0.08fF
C1820 NAND2X1_LOC_728/Y INVX1_LOC_49/Y 0.07fF
C1821 NAND2X1_LOC_594/a_36_24# NAND2X1_LOC_286/B 0.00fF
C1822 INVX1_LOC_90/A NOR2X1_LOC_486/Y 5.33fF
C1823 NOR2X1_LOC_554/B NOR2X1_LOC_340/A 0.03fF
C1824 INVX1_LOC_180/A INVX1_LOC_63/A 0.11fF
C1825 INVX1_LOC_103/A INVX1_LOC_78/A 0.22fF
C1826 INVX1_LOC_188/A INVX1_LOC_32/A 0.01fF
C1827 INVX1_LOC_39/A INVX1_LOC_224/Y 0.89fF
C1828 NAND2X1_LOC_633/Y NOR2X1_LOC_130/A 0.07fF
C1829 INVX1_LOC_18/A INVX1_LOC_99/A 0.03fF
C1830 NOR2X1_LOC_272/Y INVX1_LOC_270/Y 0.10fF
C1831 NOR2X1_LOC_218/Y NOR2X1_LOC_331/B 0.01fF
C1832 NOR2X1_LOC_481/A NAND2X1_LOC_475/Y 0.07fF
C1833 NOR2X1_LOC_137/A INVX1_LOC_46/A 0.05fF
C1834 NOR2X1_LOC_357/Y NOR2X1_LOC_367/a_36_216# 0.01fF
C1835 INVX1_LOC_17/Y NOR2X1_LOC_824/A 0.03fF
C1836 NAND2X1_LOC_833/a_36_24# INVX1_LOC_84/A 0.00fF
C1837 NOR2X1_LOC_91/A NAND2X1_LOC_725/B 2.27fF
C1838 NOR2X1_LOC_520/B INVX1_LOC_63/A 0.07fF
C1839 INVX1_LOC_71/A NAND2X1_LOC_63/Y 0.01fF
C1840 NOR2X1_LOC_146/Y INVX1_LOC_193/A 0.01fF
C1841 INVX1_LOC_45/Y INVX1_LOC_12/A 0.03fF
C1842 NOR2X1_LOC_45/B NOR2X1_LOC_74/A 0.07fF
C1843 NAND2X1_LOC_684/a_36_24# INVX1_LOC_291/A 0.01fF
C1844 INVX1_LOC_135/A NOR2X1_LOC_859/Y 0.01fF
C1845 NAND2X1_LOC_350/A NAND2X1_LOC_454/Y 0.03fF
C1846 NOR2X1_LOC_644/A NOR2X1_LOC_850/a_36_216# 0.00fF
C1847 INVX1_LOC_86/A INVX1_LOC_91/A 0.00fF
C1848 NAND2X1_LOC_656/Y NOR2X1_LOC_122/a_36_216# 0.01fF
C1849 NOR2X1_LOC_68/A NOR2X1_LOC_48/B 0.32fF
C1850 INVX1_LOC_225/A NAND2X1_LOC_475/Y 0.00fF
C1851 D_INPUT_0 NOR2X1_LOC_813/Y 0.26fF
C1852 INVX1_LOC_292/A INVX1_LOC_78/A 0.07fF
C1853 INVX1_LOC_313/Y INVX1_LOC_14/Y 0.10fF
C1854 NOR2X1_LOC_226/A NOR2X1_LOC_592/B 0.03fF
C1855 NOR2X1_LOC_151/Y NOR2X1_LOC_209/A 0.06fF
C1856 NOR2X1_LOC_312/Y INVX1_LOC_33/Y 0.01fF
C1857 INVX1_LOC_196/Y INVX1_LOC_37/A 0.00fF
C1858 INVX1_LOC_60/Y INVX1_LOC_3/A 0.06fF
C1859 INVX1_LOC_21/A NOR2X1_LOC_678/A 0.03fF
C1860 INVX1_LOC_34/A INVX1_LOC_186/Y 0.13fF
C1861 NOR2X1_LOC_348/Y INVX1_LOC_29/Y 0.01fF
C1862 NAND2X1_LOC_740/A INVX1_LOC_12/A 0.01fF
C1863 NOR2X1_LOC_719/A NOR2X1_LOC_99/Y 0.00fF
C1864 D_INPUT_0 INVX1_LOC_280/A 0.21fF
C1865 INVX1_LOC_144/Y NOR2X1_LOC_697/Y 0.59fF
C1866 NOR2X1_LOC_160/Y NAND2X1_LOC_93/B 0.04fF
C1867 INVX1_LOC_130/Y INVX1_LOC_15/A 0.06fF
C1868 INVX1_LOC_10/A NAND2X1_LOC_698/a_36_24# 0.00fF
C1869 INVX1_LOC_41/A NAND2X1_LOC_74/B 0.14fF
C1870 NOR2X1_LOC_815/A NOR2X1_LOC_56/Y 0.00fF
C1871 INVX1_LOC_16/A NOR2X1_LOC_79/Y 0.09fF
C1872 NOR2X1_LOC_368/A NAND2X1_LOC_465/A 0.11fF
C1873 NOR2X1_LOC_78/B NOR2X1_LOC_127/Y 0.07fF
C1874 NAND2X1_LOC_9/Y INVX1_LOC_14/A 0.05fF
C1875 NOR2X1_LOC_160/Y NAND2X1_LOC_425/Y 0.04fF
C1876 INVX1_LOC_126/A INVX1_LOC_126/Y 0.10fF
C1877 NOR2X1_LOC_690/A INVX1_LOC_284/A 0.03fF
C1878 INVX1_LOC_176/A INVX1_LOC_158/Y 0.01fF
C1879 INVX1_LOC_5/A INVX1_LOC_234/Y 0.01fF
C1880 INVX1_LOC_233/A INVX1_LOC_14/A 0.11fF
C1881 NOR2X1_LOC_67/A INVX1_LOC_63/A 0.07fF
C1882 NAND2X1_LOC_578/B NOR2X1_LOC_662/A 0.15fF
C1883 INVX1_LOC_256/A INVX1_LOC_29/Y 0.05fF
C1884 NAND2X1_LOC_665/a_36_24# INVX1_LOC_280/A 0.01fF
C1885 NOR2X1_LOC_413/Y INVX1_LOC_284/A 0.01fF
C1886 NOR2X1_LOC_8/a_36_216# NOR2X1_LOC_38/B 0.00fF
C1887 NAND2X1_LOC_477/A NAND2X1_LOC_74/B 0.03fF
C1888 VDD NOR2X1_LOC_527/Y 0.24fF
C1889 NAND2X1_LOC_35/Y NAND2X1_LOC_561/B 0.03fF
C1890 NOR2X1_LOC_355/A NAND2X1_LOC_93/B 0.07fF
C1891 NOR2X1_LOC_262/Y INVX1_LOC_4/A 0.01fF
C1892 INVX1_LOC_25/Y NOR2X1_LOC_653/Y 0.11fF
C1893 INVX1_LOC_123/A INVX1_LOC_20/A 0.07fF
C1894 INVX1_LOC_286/Y NOR2X1_LOC_654/A 0.10fF
C1895 INVX1_LOC_135/A INVX1_LOC_46/Y 0.03fF
C1896 NOR2X1_LOC_717/B NOR2X1_LOC_197/B 0.03fF
C1897 NAND2X1_LOC_553/A INVX1_LOC_14/A 0.01fF
C1898 INVX1_LOC_217/A NOR2X1_LOC_693/Y 0.89fF
C1899 NOR2X1_LOC_74/A INVX1_LOC_281/A 0.07fF
C1900 NOR2X1_LOC_798/A INVX1_LOC_14/A 0.03fF
C1901 INVX1_LOC_298/Y NAND2X1_LOC_656/A 0.03fF
C1902 NAND2X1_LOC_361/Y NOR2X1_LOC_839/B 0.02fF
C1903 INVX1_LOC_25/Y INVX1_LOC_19/A 0.16fF
C1904 INVX1_LOC_266/Y INVX1_LOC_283/A 0.00fF
C1905 NOR2X1_LOC_644/A INVX1_LOC_307/A 0.02fF
C1906 INVX1_LOC_16/A NOR2X1_LOC_36/B 0.02fF
C1907 INVX1_LOC_49/A NAND2X1_LOC_467/a_36_24# 0.01fF
C1908 NOR2X1_LOC_356/A NOR2X1_LOC_862/B 0.10fF
C1909 NAND2X1_LOC_364/A INVX1_LOC_270/Y 0.11fF
C1910 NAND2X1_LOC_338/B NOR2X1_LOC_38/a_36_216# 0.00fF
C1911 NOR2X1_LOC_87/Y NOR2X1_LOC_861/Y 0.09fF
C1912 NOR2X1_LOC_468/Y NAND2X1_LOC_347/B 0.45fF
C1913 NOR2X1_LOC_68/A NAND2X1_LOC_215/A 1.06fF
C1914 INVX1_LOC_67/A INVX1_LOC_78/A 0.04fF
C1915 NOR2X1_LOC_391/A NAND2X1_LOC_773/B 0.07fF
C1916 INVX1_LOC_49/A NOR2X1_LOC_449/A 0.03fF
C1917 INVX1_LOC_104/A NAND2X1_LOC_647/B 0.01fF
C1918 INVX1_LOC_181/Y INVX1_LOC_270/A 0.00fF
C1919 INVX1_LOC_58/A NOR2X1_LOC_91/Y 0.03fF
C1920 NOR2X1_LOC_142/Y NAND2X1_LOC_454/Y 0.19fF
C1921 NOR2X1_LOC_2/Y INVX1_LOC_54/A 0.09fF
C1922 NOR2X1_LOC_589/A NAND2X1_LOC_449/a_36_24# 0.00fF
C1923 NOR2X1_LOC_163/Y INVX1_LOC_92/A 0.06fF
C1924 INVX1_LOC_255/Y INVX1_LOC_12/A 0.09fF
C1925 INVX1_LOC_220/Y INVX1_LOC_29/A 0.03fF
C1926 INVX1_LOC_50/A INVX1_LOC_314/Y 0.07fF
C1927 NOR2X1_LOC_231/B INVX1_LOC_50/Y 0.05fF
C1928 INVX1_LOC_233/Y NOR2X1_LOC_384/Y 0.03fF
C1929 NAND2X1_LOC_850/Y INVX1_LOC_15/A 0.07fF
C1930 NOR2X1_LOC_151/Y NOR2X1_LOC_197/B 0.10fF
C1931 NOR2X1_LOC_457/B NOR2X1_LOC_717/A 0.01fF
C1932 INVX1_LOC_162/Y NOR2X1_LOC_301/A 0.12fF
C1933 NOR2X1_LOC_15/Y NAND2X1_LOC_793/Y 0.12fF
C1934 NOR2X1_LOC_434/Y NOR2X1_LOC_500/B 0.03fF
C1935 INVX1_LOC_8/A NAND2X1_LOC_99/A 0.64fF
C1936 NOR2X1_LOC_186/Y INVX1_LOC_30/A 0.55fF
C1937 NOR2X1_LOC_123/B NAND2X1_LOC_63/Y 0.02fF
C1938 NOR2X1_LOC_607/a_36_216# INVX1_LOC_53/A 0.01fF
C1939 NOR2X1_LOC_703/A NOR2X1_LOC_814/A 0.00fF
C1940 INVX1_LOC_39/A INVX1_LOC_45/A 0.03fF
C1941 INVX1_LOC_311/A NAND2X1_LOC_435/a_36_24# 0.00fF
C1942 NOR2X1_LOC_749/Y NAND2X1_LOC_63/Y 0.01fF
C1943 NAND2X1_LOC_866/B NAND2X1_LOC_500/B 0.02fF
C1944 NOR2X1_LOC_631/B INVX1_LOC_44/A 0.28fF
C1945 INVX1_LOC_85/A NOR2X1_LOC_302/A 0.00fF
C1946 NOR2X1_LOC_147/B INVX1_LOC_275/Y 0.01fF
C1947 NOR2X1_LOC_71/Y INVX1_LOC_12/A 0.08fF
C1948 INVX1_LOC_7/Y INVX1_LOC_136/A 0.01fF
C1949 NOR2X1_LOC_486/Y INVX1_LOC_38/A 0.03fF
C1950 NOR2X1_LOC_147/B NOR2X1_LOC_748/A 0.12fF
C1951 INVX1_LOC_103/A NOR2X1_LOC_503/Y 0.14fF
C1952 INVX1_LOC_290/A D_INPUT_5 0.22fF
C1953 INVX1_LOC_2/A NOR2X1_LOC_449/A 0.03fF
C1954 INVX1_LOC_122/Y NOR2X1_LOC_249/Y 0.13fF
C1955 NOR2X1_LOC_596/a_36_216# NOR2X1_LOC_678/A 0.00fF
C1956 NOR2X1_LOC_533/Y NOR2X1_LOC_816/A 0.08fF
C1957 NAND2X1_LOC_573/Y INVX1_LOC_30/A 0.10fF
C1958 INVX1_LOC_126/A NOR2X1_LOC_536/A 0.03fF
C1959 INVX1_LOC_282/A INVX1_LOC_84/A 0.01fF
C1960 INVX1_LOC_33/Y NAND2X1_LOC_287/B 0.01fF
C1961 NAND2X1_LOC_787/A NAND2X1_LOC_640/Y 0.01fF
C1962 NOR2X1_LOC_274/Y NOR2X1_LOC_772/B 0.00fF
C1963 INVX1_LOC_90/A INVX1_LOC_106/Y 0.01fF
C1964 NAND2X1_LOC_214/Y INVX1_LOC_36/A 0.02fF
C1965 NOR2X1_LOC_209/A NOR2X1_LOC_209/B 0.27fF
C1966 NOR2X1_LOC_329/B INVX1_LOC_29/A 0.07fF
C1967 INVX1_LOC_136/A NOR2X1_LOC_92/Y 0.22fF
C1968 INVX1_LOC_37/A INVX1_LOC_44/A 0.46fF
C1969 INVX1_LOC_1/A NOR2X1_LOC_723/Y 0.02fF
C1970 INVX1_LOC_75/A INVX1_LOC_19/A 0.08fF
C1971 NOR2X1_LOC_703/Y NOR2X1_LOC_801/A 0.02fF
C1972 NOR2X1_LOC_274/Y INVX1_LOC_13/Y 0.02fF
C1973 NAND2X1_LOC_803/B NOR2X1_LOC_590/A 0.02fF
C1974 NAND2X1_LOC_84/Y NOR2X1_LOC_798/A 0.03fF
C1975 NAND2X1_LOC_303/Y INVX1_LOC_72/A 0.10fF
C1976 NOR2X1_LOC_634/B NOR2X1_LOC_383/B 0.03fF
C1977 D_INPUT_4 INVX1_LOC_29/A 0.00fF
C1978 NOR2X1_LOC_111/A NOR2X1_LOC_536/A 0.05fF
C1979 INVX1_LOC_39/A INVX1_LOC_71/A 0.02fF
C1980 NAND2X1_LOC_555/Y INPUT_2 0.03fF
C1981 NOR2X1_LOC_78/B NOR2X1_LOC_383/B 0.13fF
C1982 NOR2X1_LOC_279/a_36_216# INVX1_LOC_57/A 0.00fF
C1983 NOR2X1_LOC_598/B INVX1_LOC_257/Y -0.00fF
C1984 INVX1_LOC_50/A NOR2X1_LOC_778/B 0.03fF
C1985 INVX1_LOC_17/A INVX1_LOC_223/A 0.01fF
C1986 INVX1_LOC_16/A INVX1_LOC_26/A 0.11fF
C1987 NAND2X1_LOC_555/Y NAND2X1_LOC_612/a_36_24# 0.00fF
C1988 NAND2X1_LOC_785/A NOR2X1_LOC_754/Y 0.01fF
C1989 NOR2X1_LOC_813/Y NAND2X1_LOC_848/A 0.07fF
C1990 NOR2X1_LOC_540/B INVX1_LOC_307/A 0.01fF
C1991 INVX1_LOC_47/A INVX1_LOC_32/A 0.03fF
C1992 NOR2X1_LOC_859/Y INVX1_LOC_280/A 0.02fF
C1993 INVX1_LOC_226/Y NOR2X1_LOC_39/Y 0.21fF
C1994 NOR2X1_LOC_824/A NOR2X1_LOC_495/Y 0.01fF
C1995 INVX1_LOC_11/A D_INPUT_7 0.01fF
C1996 NOR2X1_LOC_99/Y INVX1_LOC_76/A 0.09fF
C1997 NOR2X1_LOC_816/Y INVX1_LOC_38/A 0.01fF
C1998 NOR2X1_LOC_590/A INVX1_LOC_22/Y 0.03fF
C1999 INVX1_LOC_37/A NOR2X1_LOC_641/Y 0.11fF
C2000 INVX1_LOC_11/A NOR2X1_LOC_791/B 0.03fF
C2001 INVX1_LOC_27/A NAND2X1_LOC_361/Y 0.02fF
C2002 NOR2X1_LOC_45/Y INVX1_LOC_30/A 0.03fF
C2003 INVX1_LOC_225/Y NOR2X1_LOC_274/B 0.34fF
C2004 NAND2X1_LOC_848/A INVX1_LOC_280/A 0.01fF
C2005 NOR2X1_LOC_599/Y NOR2X1_LOC_599/A 0.03fF
C2006 INVX1_LOC_226/Y NAND2X1_LOC_205/A 0.03fF
C2007 INVX1_LOC_225/A NOR2X1_LOC_791/Y 0.02fF
C2008 NOR2X1_LOC_242/A NAND2X1_LOC_281/a_36_24# 0.00fF
C2009 NOR2X1_LOC_68/A NAND2X1_LOC_350/A 0.03fF
C2010 INVX1_LOC_107/Y INVX1_LOC_76/A 0.52fF
C2011 NOR2X1_LOC_598/B INVX1_LOC_305/Y 0.13fF
C2012 NOR2X1_LOC_91/A NOR2X1_LOC_298/Y 0.03fF
C2013 NOR2X1_LOC_255/Y INVX1_LOC_16/A 0.02fF
C2014 NOR2X1_LOC_589/A NAND2X1_LOC_231/a_36_24# 0.00fF
C2015 NOR2X1_LOC_351/Y INVX1_LOC_38/A 0.05fF
C2016 INVX1_LOC_103/A NOR2X1_LOC_152/Y 0.17fF
C2017 INVX1_LOC_55/Y INVX1_LOC_271/Y 0.07fF
C2018 NAND2X1_LOC_728/Y INVX1_LOC_161/A 0.37fF
C2019 NOR2X1_LOC_810/A NOR2X1_LOC_809/A 0.10fF
C2020 NOR2X1_LOC_331/B INVX1_LOC_118/A 0.16fF
C2021 NOR2X1_LOC_148/Y NOR2X1_LOC_209/B 0.01fF
C2022 NOR2X1_LOC_798/A NOR2X1_LOC_612/B 0.01fF
C2023 INVX1_LOC_103/A INVX1_LOC_113/Y 0.03fF
C2024 INVX1_LOC_6/A NOR2X1_LOC_114/Y 0.07fF
C2025 NOR2X1_LOC_440/Y INVX1_LOC_29/Y 0.21fF
C2026 INVX1_LOC_58/A NOR2X1_LOC_543/A 0.06fF
C2027 NOR2X1_LOC_68/A NOR2X1_LOC_441/Y 0.10fF
C2028 NOR2X1_LOC_295/Y NAND2X1_LOC_347/B 0.06fF
C2029 NOR2X1_LOC_401/Y INVX1_LOC_306/Y 0.01fF
C2030 INVX1_LOC_37/A NOR2X1_LOC_461/B 0.42fF
C2031 VDD NAND2X1_LOC_572/B 0.55fF
C2032 INVX1_LOC_34/A NOR2X1_LOC_536/Y 0.05fF
C2033 INVX1_LOC_83/A NOR2X1_LOC_383/B 0.42fF
C2034 NOR2X1_LOC_843/A INVX1_LOC_1/A 0.09fF
C2035 NOR2X1_LOC_269/Y INVX1_LOC_109/A 0.03fF
C2036 NOR2X1_LOC_310/a_36_216# INVX1_LOC_4/A 0.00fF
C2037 NAND2X1_LOC_650/B INVX1_LOC_265/Y 0.08fF
C2038 INVX1_LOC_14/A NOR2X1_LOC_140/a_36_216# 0.01fF
C2039 NAND2X1_LOC_724/Y NOR2X1_LOC_576/B 4.65fF
C2040 NAND2X1_LOC_571/B INVX1_LOC_234/A 0.17fF
C2041 INVX1_LOC_259/Y INVX1_LOC_121/A 0.08fF
C2042 INVX1_LOC_28/A INVX1_LOC_26/A 0.12fF
C2043 INVX1_LOC_97/A NOR2X1_LOC_748/A 0.01fF
C2044 INVX1_LOC_280/A INVX1_LOC_46/Y 0.38fF
C2045 NOR2X1_LOC_92/Y NAND2X1_LOC_859/a_36_24# 0.01fF
C2046 INVX1_LOC_21/A NOR2X1_LOC_191/A 0.05fF
C2047 INVX1_LOC_11/A INVX1_LOC_192/A 0.09fF
C2048 INVX1_LOC_90/A INVX1_LOC_275/Y 0.84fF
C2049 INVX1_LOC_36/A INVX1_LOC_181/Y 0.06fF
C2050 NOR2X1_LOC_369/Y NOR2X1_LOC_716/B 0.12fF
C2051 NAND2X1_LOC_93/B INVX1_LOC_127/A 0.01fF
C2052 NOR2X1_LOC_188/A INVX1_LOC_4/Y 0.32fF
C2053 NOR2X1_LOC_336/a_36_216# NAND2X1_LOC_72/B 0.00fF
C2054 INVX1_LOC_212/A NAND2X1_LOC_510/A 0.03fF
C2055 INVX1_LOC_11/A NOR2X1_LOC_124/B 0.01fF
C2056 INVX1_LOC_90/A NOR2X1_LOC_748/A 0.24fF
C2057 NOR2X1_LOC_220/B INVX1_LOC_22/A 0.01fF
C2058 NAND2X1_LOC_724/A NAND2X1_LOC_722/A 0.02fF
C2059 VDD NAND2X1_LOC_219/B 0.26fF
C2060 NOR2X1_LOC_548/B INVX1_LOC_4/Y 0.14fF
C2061 NOR2X1_LOC_267/A INVX1_LOC_181/Y 0.18fF
C2062 NAND2X1_LOC_453/A INVX1_LOC_19/A 0.07fF
C2063 INVX1_LOC_123/A INVX1_LOC_4/A 0.07fF
C2064 NOR2X1_LOC_592/B INVX1_LOC_118/A 0.01fF
C2065 INVX1_LOC_161/Y NOR2X1_LOC_320/a_36_216# 0.01fF
C2066 INVX1_LOC_76/A INVX1_LOC_272/A 1.07fF
C2067 NOR2X1_LOC_118/a_36_216# INVX1_LOC_70/A 0.02fF
C2068 INVX1_LOC_136/A NAND2X1_LOC_837/Y 0.19fF
C2069 NOR2X1_LOC_589/A NOR2X1_LOC_652/Y 0.07fF
C2070 INVX1_LOC_132/A INVX1_LOC_30/A 0.02fF
C2071 INVX1_LOC_152/Y INVX1_LOC_120/A 0.02fF
C2072 INVX1_LOC_50/A NAND2X1_LOC_123/Y 0.09fF
C2073 NOR2X1_LOC_471/Y INVX1_LOC_85/A 0.02fF
C2074 NOR2X1_LOC_481/A INVX1_LOC_30/A 0.43fF
C2075 NAND2X1_LOC_29/a_36_24# INVX1_LOC_83/A 0.01fF
C2076 INVX1_LOC_50/A NOR2X1_LOC_597/Y 0.01fF
C2077 INVX1_LOC_179/A INVX1_LOC_92/A 0.06fF
C2078 INVX1_LOC_30/A NAND2X1_LOC_640/Y 0.16fF
C2079 NOR2X1_LOC_516/B NAND2X1_LOC_218/A 0.00fF
C2080 NOR2X1_LOC_673/A INVX1_LOC_9/A 0.02fF
C2081 NOR2X1_LOC_516/B NOR2X1_LOC_140/A 0.12fF
C2082 INPUT_0 NOR2X1_LOC_843/B 0.03fF
C2083 INVX1_LOC_166/A INVX1_LOC_75/A 0.03fF
C2084 NOR2X1_LOC_160/B NOR2X1_LOC_709/A 0.24fF
C2085 NOR2X1_LOC_712/Y NOR2X1_LOC_707/B 0.16fF
C2086 NOR2X1_LOC_666/A INVX1_LOC_16/A 0.35fF
C2087 NOR2X1_LOC_624/A INVX1_LOC_45/A 0.00fF
C2088 NOR2X1_LOC_382/Y NAND2X1_LOC_139/A 0.35fF
C2089 INVX1_LOC_41/A INVX1_LOC_136/A 0.08fF
C2090 NOR2X1_LOC_690/A INVX1_LOC_72/A 0.07fF
C2091 INVX1_LOC_225/A INVX1_LOC_30/A 1.47fF
C2092 INVX1_LOC_232/Y NAND2X1_LOC_563/a_36_24# -0.03fF
C2093 NOR2X1_LOC_89/A INVX1_LOC_37/Y 0.02fF
C2094 NAND2X1_LOC_773/Y INVX1_LOC_13/A 0.17fF
C2095 NOR2X1_LOC_163/Y INVX1_LOC_53/A 0.00fF
C2096 INVX1_LOC_171/A NOR2X1_LOC_652/Y 0.00fF
C2097 INVX1_LOC_36/A NOR2X1_LOC_192/a_36_216# 0.00fF
C2098 INVX1_LOC_90/A NOR2X1_LOC_304/Y 0.03fF
C2099 NOR2X1_LOC_68/A NOR2X1_LOC_340/Y 0.01fF
C2100 INVX1_LOC_34/A INVX1_LOC_18/A 0.33fF
C2101 NOR2X1_LOC_363/Y NOR2X1_LOC_89/A 0.19fF
C2102 INVX1_LOC_255/Y NOR2X1_LOC_643/A 0.01fF
C2103 NOR2X1_LOC_243/B NOR2X1_LOC_862/B 0.00fF
C2104 INVX1_LOC_73/A NOR2X1_LOC_717/A 0.44fF
C2105 NAND2X1_LOC_728/Y INVX1_LOC_34/A 0.07fF
C2106 INVX1_LOC_110/A NOR2X1_LOC_844/A 0.00fF
C2107 NOR2X1_LOC_274/Y INVX1_LOC_303/A -0.03fF
C2108 NOR2X1_LOC_194/Y INVX1_LOC_72/A 0.02fF
C2109 NOR2X1_LOC_538/B NOR2X1_LOC_748/Y 0.16fF
C2110 INVX1_LOC_255/Y INVX1_LOC_228/Y 0.05fF
C2111 INVX1_LOC_309/A INVX1_LOC_57/A 0.06fF
C2112 INVX1_LOC_136/A NAND2X1_LOC_477/A 0.10fF
C2113 INVX1_LOC_69/Y INVX1_LOC_29/Y 0.07fF
C2114 NOR2X1_LOC_209/Y INVX1_LOC_30/A 0.07fF
C2115 INVX1_LOC_106/Y INVX1_LOC_38/A 0.12fF
C2116 NOR2X1_LOC_791/B NOR2X1_LOC_52/B 0.00fF
C2117 INVX1_LOC_34/A NAND2X1_LOC_711/B 0.03fF
C2118 INVX1_LOC_225/Y INVX1_LOC_22/A 0.03fF
C2119 NAND2X1_LOC_656/A INVX1_LOC_8/A 0.01fF
C2120 INVX1_LOC_58/A NAND2X1_LOC_450/a_36_24# 0.00fF
C2121 NOR2X1_LOC_309/Y INVX1_LOC_181/Y 0.02fF
C2122 INVX1_LOC_13/A INVX1_LOC_252/Y 0.02fF
C2123 NOR2X1_LOC_448/Y INVX1_LOC_295/A 0.01fF
C2124 NOR2X1_LOC_637/B NAND2X1_LOC_585/a_36_24# 0.02fF
C2125 INVX1_LOC_72/A NAND2X1_LOC_675/a_36_24# 0.01fF
C2126 INVX1_LOC_50/A NOR2X1_LOC_557/A 0.07fF
C2127 INVX1_LOC_200/Y NOR2X1_LOC_528/Y 0.69fF
C2128 INVX1_LOC_34/A INVX1_LOC_172/A 0.10fF
C2129 NOR2X1_LOC_561/Y INVX1_LOC_150/Y 0.10fF
C2130 NAND2X1_LOC_9/Y INVX1_LOC_48/A 0.10fF
C2131 NAND2X1_LOC_231/Y INVX1_LOC_18/A 0.02fF
C2132 INVX1_LOC_57/A INVX1_LOC_91/A 0.31fF
C2133 VDD NOR2X1_LOC_394/Y 0.27fF
C2134 NOR2X1_LOC_669/Y INVX1_LOC_90/A 0.57fF
C2135 NAND2X1_LOC_725/B NAND2X1_LOC_866/B 0.07fF
C2136 NOR2X1_LOC_419/a_36_216# NOR2X1_LOC_6/B 0.00fF
C2137 NOR2X1_LOC_655/B NOR2X1_LOC_68/A 0.03fF
C2138 NOR2X1_LOC_647/A NAND2X1_LOC_819/a_36_24# 0.00fF
C2139 NOR2X1_LOC_113/A INVX1_LOC_270/Y 0.16fF
C2140 NOR2X1_LOC_305/Y NAND2X1_LOC_175/Y 0.07fF
C2141 INVX1_LOC_89/Y INVX1_LOC_12/A 0.01fF
C2142 NOR2X1_LOC_139/Y INVX1_LOC_23/A 0.05fF
C2143 NOR2X1_LOC_405/A INVX1_LOC_270/Y 0.33fF
C2144 NOR2X1_LOC_675/A INVX1_LOC_270/A 0.07fF
C2145 NOR2X1_LOC_496/Y NAND2X1_LOC_849/A 0.06fF
C2146 INVX1_LOC_256/A NOR2X1_LOC_355/A 0.15fF
C2147 NAND2X1_LOC_363/B NAND2X1_LOC_669/a_36_24# 0.00fF
C2148 INVX1_LOC_12/Y NOR2X1_LOC_334/Y 0.10fF
C2149 NOR2X1_LOC_666/A INVX1_LOC_28/A 0.12fF
C2150 INVX1_LOC_14/A NAND2X1_LOC_842/B 0.16fF
C2151 NOR2X1_LOC_56/Y NOR2X1_LOC_654/A 0.02fF
C2152 NAND2X1_LOC_30/Y INVX1_LOC_295/A 0.08fF
C2153 NOR2X1_LOC_590/A INVX1_LOC_227/A 0.08fF
C2154 INVX1_LOC_136/A NOR2X1_LOC_211/A 0.04fF
C2155 NOR2X1_LOC_510/Y NOR2X1_LOC_815/A 0.00fF
C2156 NOR2X1_LOC_577/Y INVX1_LOC_266/Y 0.18fF
C2157 NOR2X1_LOC_705/B INVX1_LOC_89/A 0.01fF
C2158 INVX1_LOC_254/A NAND2X1_LOC_338/B 0.01fF
C2159 NOR2X1_LOC_689/A INVX1_LOC_46/A 0.03fF
C2160 NAND2X1_LOC_468/B INVX1_LOC_23/A 0.06fF
C2161 NOR2X1_LOC_593/Y NOR2X1_LOC_802/A 0.10fF
C2162 NOR2X1_LOC_133/a_36_216# INVX1_LOC_26/A 0.00fF
C2163 NAND2X1_LOC_363/B NAND2X1_LOC_642/Y 0.02fF
C2164 NOR2X1_LOC_533/A NOR2X1_LOC_152/Y 0.09fF
C2165 NOR2X1_LOC_383/B INVX1_LOC_46/A 0.13fF
C2166 INVX1_LOC_146/Y NOR2X1_LOC_654/A 0.04fF
C2167 INVX1_LOC_247/Y INVX1_LOC_220/Y 0.02fF
C2168 NOR2X1_LOC_533/Y INVX1_LOC_140/A 0.35fF
C2169 D_INPUT_1 INVX1_LOC_20/A 0.13fF
C2170 VDD NOR2X1_LOC_654/A 1.22fF
C2171 INVX1_LOC_286/A NAND2X1_LOC_474/Y 0.19fF
C2172 INVX1_LOC_2/A NOR2X1_LOC_388/Y 0.07fF
C2173 INVX1_LOC_277/Y INVX1_LOC_83/A 0.01fF
C2174 NAND2X1_LOC_182/a_36_24# INVX1_LOC_71/A 0.00fF
C2175 INVX1_LOC_34/A INVX1_LOC_34/Y 0.15fF
C2176 NOR2X1_LOC_844/Y INVX1_LOC_120/A 0.01fF
C2177 NOR2X1_LOC_122/Y NOR2X1_LOC_276/Y 0.00fF
C2178 NAND2X1_LOC_738/B INVX1_LOC_46/A 0.03fF
C2179 NOR2X1_LOC_156/Y NOR2X1_LOC_467/A 0.02fF
C2180 NOR2X1_LOC_348/B INVX1_LOC_266/Y 0.10fF
C2181 INVX1_LOC_276/Y NAND2X1_LOC_354/B 0.00fF
C2182 INVX1_LOC_276/A NAND2X1_LOC_326/a_36_24# 0.00fF
C2183 INVX1_LOC_57/A NOR2X1_LOC_653/a_36_216# 0.00fF
C2184 NOR2X1_LOC_327/a_36_216# INVX1_LOC_63/A 0.01fF
C2185 INVX1_LOC_28/A INVX1_LOC_141/A 0.05fF
C2186 NOR2X1_LOC_480/A NOR2X1_LOC_459/A 0.01fF
C2187 NOR2X1_LOC_13/Y NOR2X1_LOC_781/A 0.28fF
C2188 INVX1_LOC_161/Y INVX1_LOC_75/A 0.10fF
C2189 NOR2X1_LOC_391/A INVX1_LOC_24/A 0.03fF
C2190 NOR2X1_LOC_68/A NOR2X1_LOC_99/B 0.14fF
C2191 INVX1_LOC_217/A NOR2X1_LOC_71/Y 0.01fF
C2192 NAND2X1_LOC_766/a_36_24# INVX1_LOC_22/A 0.00fF
C2193 NAND2X1_LOC_342/Y INVX1_LOC_104/A 0.05fF
C2194 NOR2X1_LOC_791/Y NAND2X1_LOC_642/Y 0.02fF
C2195 NAND2X1_LOC_708/Y INVX1_LOC_76/A 0.06fF
C2196 VDD INVX1_LOC_58/Y 0.68fF
C2197 INVX1_LOC_315/Y NAND2X1_LOC_218/A 0.02fF
C2198 NOR2X1_LOC_570/B NOR2X1_LOC_500/Y 0.07fF
C2199 INVX1_LOC_83/A NOR2X1_LOC_512/Y 0.02fF
C2200 INVX1_LOC_256/A NOR2X1_LOC_541/a_36_216# 0.00fF
C2201 NAND2X1_LOC_738/B NOR2X1_LOC_766/Y 0.41fF
C2202 NAND2X1_LOC_854/B NAND2X1_LOC_567/Y 0.01fF
C2203 INVX1_LOC_38/A NOR2X1_LOC_748/A 0.03fF
C2204 INVX1_LOC_95/A NAND2X1_LOC_474/Y 0.00fF
C2205 NAND2X1_LOC_811/Y INVX1_LOC_22/A 0.03fF
C2206 INVX1_LOC_311/Y INVX1_LOC_142/A 0.34fF
C2207 NAND2X1_LOC_787/A NOR2X1_LOC_495/a_36_216# 0.00fF
C2208 NAND2X1_LOC_722/A NAND2X1_LOC_852/Y 0.10fF
C2209 INVX1_LOC_34/A NOR2X1_LOC_690/Y 0.03fF
C2210 INVX1_LOC_135/A INVX1_LOC_49/A 0.10fF
C2211 INVX1_LOC_164/Y INVX1_LOC_256/Y 0.04fF
C2212 NOR2X1_LOC_821/Y INVX1_LOC_22/A 0.20fF
C2213 NOR2X1_LOC_68/A INVX1_LOC_182/A 0.10fF
C2214 INVX1_LOC_131/A INVX1_LOC_18/A 0.01fF
C2215 INVX1_LOC_70/A INVX1_LOC_181/A 0.05fF
C2216 INVX1_LOC_266/Y INVX1_LOC_22/A 0.18fF
C2217 INVX1_LOC_295/A INVX1_LOC_49/A 0.19fF
C2218 NAND2X1_LOC_363/B NOR2X1_LOC_271/Y 0.33fF
C2219 INVX1_LOC_2/A NAND2X1_LOC_479/Y 0.03fF
C2220 NAND2X1_LOC_367/B GATE_366 0.01fF
C2221 INVX1_LOC_219/Y INVX1_LOC_234/A 0.02fF
C2222 INVX1_LOC_177/Y INVX1_LOC_67/Y 0.06fF
C2223 INVX1_LOC_49/A NOR2X1_LOC_560/A 0.00fF
C2224 NOR2X1_LOC_392/B INVX1_LOC_150/A 0.26fF
C2225 INVX1_LOC_76/A INVX1_LOC_198/A 0.14fF
C2226 INVX1_LOC_78/A NOR2X1_LOC_631/A 0.07fF
C2227 INVX1_LOC_136/A NAND2X1_LOC_662/B 0.05fF
C2228 INVX1_LOC_18/A INPUT_0 0.15fF
C2229 INVX1_LOC_89/A NOR2X1_LOC_147/B 0.08fF
C2230 NOR2X1_LOC_248/a_36_216# INVX1_LOC_49/A 0.01fF
C2231 NOR2X1_LOC_296/Y INVX1_LOC_95/Y 0.11fF
C2232 NAND2X1_LOC_728/Y INPUT_0 0.07fF
C2233 INVX1_LOC_89/A NOR2X1_LOC_392/B 0.00fF
C2234 NAND2X1_LOC_341/A NOR2X1_LOC_219/Y 0.13fF
C2235 NOR2X1_LOC_437/Y INVX1_LOC_75/A 0.10fF
C2236 INVX1_LOC_31/A NAND2X1_LOC_655/A 0.07fF
C2237 NOR2X1_LOC_740/Y INVX1_LOC_76/A 0.17fF
C2238 NOR2X1_LOC_272/Y NOR2X1_LOC_536/A 0.01fF
C2239 INVX1_LOC_53/A INVX1_LOC_179/A 0.12fF
C2240 NOR2X1_LOC_791/Y NOR2X1_LOC_271/Y 0.03fF
C2241 NOR2X1_LOC_254/A NOR2X1_LOC_631/B 0.12fF
C2242 NAND2X1_LOC_711/B INPUT_0 0.06fF
C2243 NAND2X1_LOC_338/B NAND2X1_LOC_358/a_36_24# 0.00fF
C2244 INVX1_LOC_2/A INVX1_LOC_135/A 0.13fF
C2245 NOR2X1_LOC_179/Y INVX1_LOC_57/A 0.04fF
C2246 NOR2X1_LOC_246/Y INVX1_LOC_104/A 0.03fF
C2247 INVX1_LOC_119/A INVX1_LOC_90/A 0.04fF
C2248 NOR2X1_LOC_178/Y NOR2X1_LOC_99/Y 0.01fF
C2249 NOR2X1_LOC_135/Y NAND2X1_LOC_332/Y 0.09fF
C2250 NAND2X1_LOC_63/Y NOR2X1_LOC_621/B 0.04fF
C2251 NOR2X1_LOC_419/Y NOR2X1_LOC_721/Y 0.00fF
C2252 NOR2X1_LOC_371/a_36_216# INVX1_LOC_20/A 0.00fF
C2253 NOR2X1_LOC_226/A INVX1_LOC_135/A 0.10fF
C2254 INVX1_LOC_172/A INPUT_0 0.07fF
C2255 NOR2X1_LOC_299/Y NAND2X1_LOC_507/a_36_24# 0.01fF
C2256 INVX1_LOC_30/A NAND2X1_LOC_642/Y 0.99fF
C2257 NOR2X1_LOC_75/Y VDD 0.91fF
C2258 NOR2X1_LOC_334/Y NOR2X1_LOC_842/a_36_216# 0.01fF
C2259 INVX1_LOC_36/A NAND2X1_LOC_107/a_36_24# 0.01fF
C2260 D_INPUT_5 NOR2X1_LOC_467/A 0.72fF
C2261 INVX1_LOC_161/Y NOR2X1_LOC_65/a_36_216# 0.01fF
C2262 INVX1_LOC_50/A NAND2X1_LOC_625/a_36_24# 0.00fF
C2263 NOR2X1_LOC_716/B NOR2X1_LOC_721/Y 0.02fF
C2264 NAND2X1_LOC_783/Y VDD 0.00fF
C2265 NAND2X1_LOC_36/A NAND2X1_LOC_1/Y 0.89fF
C2266 NAND2X1_LOC_402/B INVX1_LOC_167/A 0.01fF
C2267 INVX1_LOC_265/A NOR2X1_LOC_74/A 0.04fF
C2268 INVX1_LOC_21/A NAND2X1_LOC_60/a_36_24# 0.01fF
C2269 INVX1_LOC_104/A INVX1_LOC_67/Y 0.00fF
C2270 NAND2X1_LOC_114/B INVX1_LOC_117/A 0.15fF
C2271 INVX1_LOC_32/A INVX1_LOC_271/Y 0.07fF
C2272 INVX1_LOC_295/A NOR2X1_LOC_161/Y 0.04fF
C2273 INVX1_LOC_2/A NOR2X1_LOC_202/Y 0.02fF
C2274 NOR2X1_LOC_134/Y NOR2X1_LOC_813/Y 0.04fF
C2275 INVX1_LOC_45/A INVX1_LOC_14/Y 0.05fF
C2276 NOR2X1_LOC_805/a_36_216# NOR2X1_LOC_729/A 0.02fF
C2277 INVX1_LOC_57/Y INVX1_LOC_46/A 0.02fF
C2278 INVX1_LOC_135/A NAND2X1_LOC_462/B 0.05fF
C2279 NOR2X1_LOC_523/A NOR2X1_LOC_61/Y 0.01fF
C2280 NOR2X1_LOC_114/Y INVX1_LOC_270/A 0.10fF
C2281 NOR2X1_LOC_89/A INVX1_LOC_29/Y 1.61fF
C2282 INPUT_0 INVX1_LOC_34/Y 0.07fF
C2283 NAND2X1_LOC_53/Y INVX1_LOC_54/A 0.48fF
C2284 INVX1_LOC_1/A NOR2X1_LOC_156/Y 0.01fF
C2285 NAND2X1_LOC_361/a_36_24# INVX1_LOC_125/Y 0.00fF
C2286 NAND2X1_LOC_863/A NAND2X1_LOC_853/Y 0.30fF
C2287 INVX1_LOC_35/A INVX1_LOC_29/A 0.92fF
C2288 NOR2X1_LOC_716/B NOR2X1_LOC_123/a_36_216# 0.01fF
C2289 NOR2X1_LOC_298/Y NAND2X1_LOC_866/B 0.10fF
C2290 INVX1_LOC_103/A NAND2X1_LOC_802/Y 0.07fF
C2291 INVX1_LOC_55/Y INVX1_LOC_279/A 0.07fF
C2292 INVX1_LOC_84/A NOR2X1_LOC_440/B 0.07fF
C2293 NAND2X1_LOC_35/Y NAND2X1_LOC_74/B 0.07fF
C2294 INVX1_LOC_89/A INVX1_LOC_97/A 0.03fF
C2295 INVX1_LOC_135/A INPUT_1 0.41fF
C2296 NAND2X1_LOC_162/B VDD 0.01fF
C2297 NAND2X1_LOC_703/a_36_24# NAND2X1_LOC_808/A 0.01fF
C2298 INVX1_LOC_42/Y INVX1_LOC_22/A 0.06fF
C2299 INVX1_LOC_71/A INVX1_LOC_14/Y 0.50fF
C2300 NOR2X1_LOC_646/B NOR2X1_LOC_38/B 0.00fF
C2301 NOR2X1_LOC_258/a_36_216# NAND2X1_LOC_93/B 0.00fF
C2302 INVX1_LOC_23/A NOR2X1_LOC_685/Y 0.01fF
C2303 INVX1_LOC_90/A INVX1_LOC_89/A 3.17fF
C2304 NAND2X1_LOC_364/A NOR2X1_LOC_536/A 0.05fF
C2305 NOR2X1_LOC_238/Y NAND2X1_LOC_804/Y 0.01fF
C2306 INVX1_LOC_16/A NOR2X1_LOC_368/A 0.02fF
C2307 NOR2X1_LOC_310/Y NOR2X1_LOC_405/A 0.01fF
C2308 NOR2X1_LOC_309/Y NOR2X1_LOC_675/A 0.01fF
C2309 NOR2X1_LOC_419/Y VDD 1.84fF
C2310 NAND2X1_LOC_769/a_36_24# INVX1_LOC_89/A 0.00fF
C2311 NAND2X1_LOC_214/Y INVX1_LOC_63/A 0.01fF
C2312 NAND2X1_LOC_337/B NOR2X1_LOC_831/B 0.01fF
C2313 NOR2X1_LOC_546/B INVX1_LOC_117/A 0.00fF
C2314 NOR2X1_LOC_389/B INVX1_LOC_89/A 0.07fF
C2315 D_INPUT_1 INVX1_LOC_4/A 0.07fF
C2316 INVX1_LOC_49/A INVX1_LOC_139/Y 0.03fF
C2317 NOR2X1_LOC_124/B INVX1_LOC_74/A 0.03fF
C2318 NOR2X1_LOC_391/Y INVX1_LOC_232/A 0.01fF
C2319 INVX1_LOC_159/A NAND2X1_LOC_423/a_36_24# 0.00fF
C2320 INPUT_6 INVX1_LOC_15/A 0.02fF
C2321 NOR2X1_LOC_258/a_36_216# NAND2X1_LOC_425/Y 0.01fF
C2322 NOR2X1_LOC_329/B NAND2X1_LOC_140/A 0.02fF
C2323 NOR2X1_LOC_716/B VDD 2.91fF
C2324 NAND2X1_LOC_100/a_36_24# NOR2X1_LOC_536/A 0.00fF
C2325 INVX1_LOC_83/A NOR2X1_LOC_163/Y 0.02fF
C2326 NOR2X1_LOC_677/Y INVX1_LOC_78/A 0.10fF
C2327 NOR2X1_LOC_690/Y INPUT_0 0.47fF
C2328 NAND2X1_LOC_20/B NOR2X1_LOC_673/A 0.13fF
C2329 NOR2X1_LOC_321/Y INVX1_LOC_49/Y 0.01fF
C2330 NAND2X1_LOC_348/A NOR2X1_LOC_719/a_36_216# 0.00fF
C2331 NOR2X1_LOC_144/Y NOR2X1_LOC_357/Y 0.05fF
C2332 NOR2X1_LOC_433/A NOR2X1_LOC_363/Y 0.04fF
C2333 NOR2X1_LOC_383/a_36_216# INPUT_0 0.00fF
C2334 INVX1_LOC_269/A NAND2X1_LOC_773/B 0.10fF
C2335 INVX1_LOC_253/A NOR2X1_LOC_476/B 0.00fF
C2336 NAND2X1_LOC_624/B INVX1_LOC_15/A 0.01fF
C2337 INVX1_LOC_69/Y INVX1_LOC_101/A 0.03fF
C2338 NOR2X1_LOC_591/Y INVX1_LOC_20/A 0.05fF
C2339 NAND2X1_LOC_325/Y NAND2X1_LOC_721/A 0.01fF
C2340 INVX1_LOC_275/A INVX1_LOC_117/A 0.03fF
C2341 NOR2X1_LOC_233/a_36_216# INVX1_LOC_42/A 0.00fF
C2342 NOR2X1_LOC_191/B NOR2X1_LOC_709/B 0.01fF
C2343 NAND2X1_LOC_348/A INVX1_LOC_89/A 0.17fF
C2344 NOR2X1_LOC_529/Y INVX1_LOC_20/A 0.07fF
C2345 INVX1_LOC_55/Y INVX1_LOC_182/Y 0.03fF
C2346 NAND2X1_LOC_364/A NAND2X1_LOC_93/B 0.03fF
C2347 INVX1_LOC_234/Y INVX1_LOC_42/A 0.10fF
C2348 INVX1_LOC_286/A INVX1_LOC_10/A 0.07fF
C2349 NOR2X1_LOC_849/A INVX1_LOC_15/A 0.03fF
C2350 INVX1_LOC_290/A NOR2X1_LOC_269/Y 0.00fF
C2351 NOR2X1_LOC_355/A INVX1_LOC_69/Y 0.01fF
C2352 NOR2X1_LOC_815/Y NOR2X1_LOC_331/B 0.02fF
C2353 NAND2X1_LOC_348/A NAND2X1_LOC_508/A 0.12fF
C2354 INVX1_LOC_14/A INVX1_LOC_284/A 0.57fF
C2355 INVX1_LOC_31/A NOR2X1_LOC_820/B 0.04fF
C2356 INVX1_LOC_296/A INVX1_LOC_296/Y 0.02fF
C2357 NOR2X1_LOC_652/Y INVX1_LOC_4/A -0.04fF
C2358 NOR2X1_LOC_52/B INVX1_LOC_37/Y 0.14fF
C2359 INVX1_LOC_45/Y INVX1_LOC_92/A 0.14fF
C2360 INVX1_LOC_2/A INVX1_LOC_139/Y 0.03fF
C2361 INVX1_LOC_50/A INVX1_LOC_271/A 0.07fF
C2362 INVX1_LOC_35/A INVX1_LOC_298/Y 0.00fF
C2363 INVX1_LOC_98/Y VDD 0.02fF
C2364 NOR2X1_LOC_717/B NOR2X1_LOC_337/Y 0.02fF
C2365 NOR2X1_LOC_273/Y NOR2X1_LOC_155/A 0.02fF
C2366 INVX1_LOC_53/A NAND2X1_LOC_288/B 0.05fF
C2367 INVX1_LOC_33/A NOR2X1_LOC_351/Y 0.03fF
C2368 NOR2X1_LOC_775/Y NOR2X1_LOC_97/A 0.42fF
C2369 NOR2X1_LOC_759/Y NOR2X1_LOC_155/A 0.05fF
C2370 INVX1_LOC_127/Y NOR2X1_LOC_271/B 0.17fF
C2371 INVX1_LOC_41/Y NOR2X1_LOC_88/Y 0.03fF
C2372 NOR2X1_LOC_168/B INVX1_LOC_117/A 0.06fF
C2373 INVX1_LOC_202/A NOR2X1_LOC_155/A 0.01fF
C2374 NOR2X1_LOC_757/Y VDD 0.39fF
C2375 NAND2X1_LOC_9/Y NOR2X1_LOC_383/B 0.01fF
C2376 INVX1_LOC_2/A NOR2X1_LOC_813/Y 0.10fF
C2377 D_INPUT_0 NOR2X1_LOC_45/B 0.07fF
C2378 NAND2X1_LOC_311/a_36_24# INVX1_LOC_63/A 0.01fF
C2379 NOR2X1_LOC_67/A NAND2X1_LOC_721/A 0.03fF
C2380 INVX1_LOC_136/A INVX1_LOC_136/Y 0.04fF
C2381 INVX1_LOC_119/A INVX1_LOC_38/A 0.09fF
C2382 INVX1_LOC_272/Y NOR2X1_LOC_48/B 0.62fF
C2383 NAND2X1_LOC_331/a_36_24# NOR2X1_LOC_318/B 0.00fF
C2384 INVX1_LOC_1/A D_INPUT_5 0.06fF
C2385 NOR2X1_LOC_520/A NAND2X1_LOC_96/A -0.02fF
C2386 NOR2X1_LOC_15/Y INVX1_LOC_47/Y 0.09fF
C2387 NOR2X1_LOC_668/a_36_216# INVX1_LOC_57/A 0.00fF
C2388 NAND2X1_LOC_11/Y NAND2X1_LOC_639/A 0.25fF
C2389 NAND2X1_LOC_593/Y NOR2X1_LOC_88/Y 0.03fF
C2390 NOR2X1_LOC_550/B NOR2X1_LOC_155/A 0.03fF
C2391 INVX1_LOC_313/A NOR2X1_LOC_139/Y 0.00fF
C2392 INVX1_LOC_30/A NOR2X1_LOC_48/Y 0.05fF
C2393 INVX1_LOC_72/A NAND2X1_LOC_479/a_36_24# 0.00fF
C2394 INVX1_LOC_2/A INVX1_LOC_280/A 0.01fF
C2395 INVX1_LOC_233/Y NAND2X1_LOC_725/Y 0.39fF
C2396 NOR2X1_LOC_590/A NOR2X1_LOC_67/Y 0.36fF
C2397 INVX1_LOC_45/A NOR2X1_LOC_831/Y 0.01fF
C2398 NOR2X1_LOC_274/B INVX1_LOC_19/A 0.42fF
C2399 NOR2X1_LOC_575/Y INVX1_LOC_167/Y 0.01fF
C2400 INVX1_LOC_41/Y INVX1_LOC_84/A 2.61fF
C2401 INPUT_0 NOR2X1_LOC_185/a_36_216# 0.00fF
C2402 NOR2X1_LOC_91/A INVX1_LOC_13/Y 0.07fF
C2403 NAND2X1_LOC_763/B NOR2X1_LOC_48/Y 0.00fF
C2404 NOR2X1_LOC_262/a_36_216# NOR2X1_LOC_772/B 0.00fF
C2405 INVX1_LOC_181/Y INVX1_LOC_63/A 0.07fF
C2406 INVX1_LOC_232/A INVX1_LOC_129/Y 0.03fF
C2407 NAND2X1_LOC_213/A NAND2X1_LOC_470/B 0.36fF
C2408 INVX1_LOC_64/A D_INPUT_1 0.32fF
C2409 NOR2X1_LOC_470/A VDD 0.15fF
C2410 INVX1_LOC_77/A NOR2X1_LOC_450/B 0.00fF
C2411 NOR2X1_LOC_798/A NOR2X1_LOC_383/B 0.03fF
C2412 NOR2X1_LOC_424/Y VDD 0.32fF
C2413 NOR2X1_LOC_151/Y NOR2X1_LOC_337/Y 0.00fF
C2414 NOR2X1_LOC_510/Y NOR2X1_LOC_654/A 0.03fF
C2415 NOR2X1_LOC_567/B INVX1_LOC_160/A 0.02fF
C2416 INVX1_LOC_48/Y INVX1_LOC_26/A 0.02fF
C2417 NOR2X1_LOC_360/a_36_216# NAND2X1_LOC_206/Y 0.01fF
C2418 NOR2X1_LOC_326/Y VDD 0.45fF
C2419 NOR2X1_LOC_717/B VDD 0.12fF
C2420 INVX1_LOC_50/A INVX1_LOC_27/A 0.03fF
C2421 INVX1_LOC_292/A NOR2X1_LOC_609/Y 0.02fF
C2422 INVX1_LOC_13/Y INVX1_LOC_23/A 0.08fF
C2423 INVX1_LOC_13/A NOR2X1_LOC_98/B 0.02fF
C2424 NOR2X1_LOC_106/A NAND2X1_LOC_211/Y 0.08fF
C2425 NOR2X1_LOC_790/B INVX1_LOC_5/A 0.68fF
C2426 NOR2X1_LOC_86/A NOR2X1_LOC_536/A 0.84fF
C2427 INVX1_LOC_251/Y INVX1_LOC_46/Y 0.15fF
C2428 INVX1_LOC_90/A NAND2X1_LOC_244/A 0.07fF
C2429 INVX1_LOC_71/A NOR2X1_LOC_831/Y 0.12fF
C2430 NOR2X1_LOC_160/B NOR2X1_LOC_334/Y 0.15fF
C2431 INVX1_LOC_104/A INVX1_LOC_285/A 0.07fF
C2432 NOR2X1_LOC_577/Y INVX1_LOC_19/A 0.07fF
C2433 NOR2X1_LOC_130/Y VDD 0.23fF
C2434 NOR2X1_LOC_78/B INVX1_LOC_179/A 2.16fF
C2435 NOR2X1_LOC_379/Y INVX1_LOC_19/A 0.27fF
C2436 NOR2X1_LOC_828/A VDD 0.25fF
C2437 NOR2X1_LOC_497/Y INVX1_LOC_20/A 0.02fF
C2438 INVX1_LOC_142/A INVX1_LOC_15/A 0.05fF
C2439 INVX1_LOC_104/A NOR2X1_LOC_814/A 0.09fF
C2440 NOR2X1_LOC_859/A INVX1_LOC_15/A 0.10fF
C2441 NOR2X1_LOC_255/Y INVX1_LOC_48/Y 0.19fF
C2442 NOR2X1_LOC_139/Y INVX1_LOC_6/A 4.14fF
C2443 NAND2X1_LOC_214/B NAND2X1_LOC_749/a_36_24# 0.00fF
C2444 NOR2X1_LOC_753/a_36_216# NOR2X1_LOC_89/A 0.02fF
C2445 INVX1_LOC_16/A NOR2X1_LOC_235/Y 0.02fF
C2446 NOR2X1_LOC_813/Y INPUT_1 0.15fF
C2447 INVX1_LOC_135/Y VDD 0.26fF
C2448 NAND2X1_LOC_199/B NOR2X1_LOC_158/Y 0.05fF
C2449 INVX1_LOC_89/A NAND2X1_LOC_849/B 0.17fF
C2450 NAND2X1_LOC_638/Y INVX1_LOC_117/A 0.02fF
C2451 INVX1_LOC_88/A INVX1_LOC_23/A 0.19fF
C2452 NOR2X1_LOC_264/Y INVX1_LOC_125/A 0.13fF
C2453 NOR2X1_LOC_163/Y INVX1_LOC_46/A 0.00fF
C2454 INVX1_LOC_10/A INVX1_LOC_54/A 0.61fF
C2455 INVX1_LOC_89/A INVX1_LOC_38/A 0.13fF
C2456 INVX1_LOC_223/A INVX1_LOC_94/Y 0.00fF
C2457 INVX1_LOC_135/A INVX1_LOC_118/A 0.10fF
C2458 INVX1_LOC_41/Y INVX1_LOC_15/A 0.03fF
C2459 INVX1_LOC_266/Y INVX1_LOC_186/Y 0.10fF
C2460 NOR2X1_LOC_151/Y VDD 1.35fF
C2461 NOR2X1_LOC_322/Y INVX1_LOC_37/A 0.07fF
C2462 NAND2X1_LOC_468/B INVX1_LOC_6/A 0.03fF
C2463 NAND2X1_LOC_391/Y INVX1_LOC_306/Y 0.02fF
C2464 NAND2X1_LOC_550/A NAND2X1_LOC_464/B 0.65fF
C2465 INPUT_1 INVX1_LOC_280/A 0.09fF
C2466 NAND2X1_LOC_169/Y INVX1_LOC_178/A 0.06fF
C2467 INVX1_LOC_217/Y INVX1_LOC_284/A -0.02fF
C2468 INVX1_LOC_89/A NOR2X1_LOC_96/Y 0.03fF
C2469 NOR2X1_LOC_617/Y INVX1_LOC_15/A 0.00fF
C2470 NOR2X1_LOC_515/a_36_216# NAND2X1_LOC_82/Y 0.00fF
C2471 NOR2X1_LOC_483/B NOR2X1_LOC_748/A 0.01fF
C2472 NOR2X1_LOC_178/Y NOR2X1_LOC_271/B 0.11fF
C2473 INVX1_LOC_107/A NOR2X1_LOC_158/Y 0.04fF
C2474 NAND2X1_LOC_725/A NAND2X1_LOC_561/B 0.13fF
C2475 D_INPUT_1 INVX1_LOC_43/Y -0.00fF
C2476 NOR2X1_LOC_212/a_36_216# INVX1_LOC_1/A 0.00fF
C2477 NOR2X1_LOC_346/B INVX1_LOC_19/A 5.55fF
C2478 NOR2X1_LOC_329/B INVX1_LOC_118/Y 0.07fF
C2479 D_INPUT_0 NOR2X1_LOC_862/B 0.01fF
C2480 NOR2X1_LOC_361/Y NOR2X1_LOC_89/A 0.01fF
C2481 NOR2X1_LOC_562/B NOR2X1_LOC_631/B 0.27fF
C2482 INVX1_LOC_147/A NAND2X1_LOC_61/a_36_24# 0.01fF
C2483 INVX1_LOC_174/A INVX1_LOC_295/Y 0.01fF
C2484 INVX1_LOC_286/Y NOR2X1_LOC_591/A 0.02fF
C2485 INVX1_LOC_7/A NOR2X1_LOC_673/A 0.03fF
C2486 NOR2X1_LOC_500/B INVX1_LOC_23/A 0.00fF
C2487 INVX1_LOC_22/A INVX1_LOC_19/A 0.25fF
C2488 INVX1_LOC_186/A NOR2X1_LOC_858/B 0.07fF
C2489 NOR2X1_LOC_544/a_36_216# NOR2X1_LOC_334/Y 0.01fF
C2490 INVX1_LOC_56/A NAND2X1_LOC_74/B 0.05fF
C2491 INVX1_LOC_22/A NOR2X1_LOC_11/Y 2.75fF
C2492 INVX1_LOC_78/Y INVX1_LOC_117/A 0.03fF
C2493 INVX1_LOC_93/Y NOR2X1_LOC_558/A 0.01fF
C2494 NOR2X1_LOC_689/A NAND2X1_LOC_866/A 0.16fF
C2495 NOR2X1_LOC_272/Y INVX1_LOC_256/A 0.37fF
C2496 INVX1_LOC_17/A NOR2X1_LOC_454/Y 0.07fF
C2497 INVX1_LOC_244/Y INVX1_LOC_57/A 0.02fF
C2498 INVX1_LOC_233/A INVX1_LOC_57/Y 0.10fF
C2499 NAND2X1_LOC_214/B INVX1_LOC_61/Y 0.01fF
C2500 NOR2X1_LOC_188/Y INVX1_LOC_29/A 0.36fF
C2501 NOR2X1_LOC_121/a_36_216# INVX1_LOC_42/A 0.00fF
C2502 INVX1_LOC_152/Y NAND2X1_LOC_351/A 0.00fF
C2503 INVX1_LOC_249/A INVX1_LOC_50/A 0.05fF
C2504 NAND2X1_LOC_451/Y NOR2X1_LOC_467/A 0.92fF
C2505 INVX1_LOC_299/A NAND2X1_LOC_774/a_36_24# 0.01fF
C2506 INVX1_LOC_248/Y INVX1_LOC_141/Y 0.02fF
C2507 INVX1_LOC_13/Y INVX1_LOC_31/A 0.13fF
C2508 NAND2X1_LOC_787/A NOR2X1_LOC_91/Y 0.83fF
C2509 NOR2X1_LOC_152/Y NOR2X1_LOC_677/Y 0.04fF
C2510 NOR2X1_LOC_45/B NAND2X1_LOC_848/A 0.10fF
C2511 NAND2X1_LOC_865/a_36_24# INVX1_LOC_84/A 0.00fF
C2512 NOR2X1_LOC_751/A INVX1_LOC_92/A 0.19fF
C2513 INVX1_LOC_202/A NOR2X1_LOC_125/Y 0.19fF
C2514 NOR2X1_LOC_728/B INVX1_LOC_274/A -0.06fF
C2515 INVX1_LOC_136/A NAND2X1_LOC_35/Y 0.59fF
C2516 NOR2X1_LOC_647/A INVX1_LOC_34/A 0.01fF
C2517 NOR2X1_LOC_454/Y NOR2X1_LOC_471/Y 0.18fF
C2518 INVX1_LOC_45/Y INVX1_LOC_53/A 0.08fF
C2519 NOR2X1_LOC_113/A NOR2X1_LOC_536/A 0.09fF
C2520 INVX1_LOC_105/A INVX1_LOC_105/Y 0.10fF
C2521 NOR2X1_LOC_405/A NOR2X1_LOC_536/A 0.16fF
C2522 NAND2X1_LOC_360/B INVX1_LOC_4/Y 0.49fF
C2523 INVX1_LOC_214/Y INVX1_LOC_21/Y 0.96fF
C2524 INVX1_LOC_278/A INVX1_LOC_41/Y 0.45fF
C2525 INVX1_LOC_33/A INVX1_LOC_275/Y 0.04fF
C2526 INVX1_LOC_33/A NOR2X1_LOC_748/A 0.03fF
C2527 NAND2X1_LOC_633/Y VDD 0.43fF
C2528 NAND2X1_LOC_738/B NAND2X1_LOC_812/A 0.00fF
C2529 NOR2X1_LOC_355/A NOR2X1_LOC_89/A 0.03fF
C2530 NOR2X1_LOC_84/Y INVX1_LOC_26/A 0.06fF
C2531 INVX1_LOC_64/A NOR2X1_LOC_403/B 0.16fF
C2532 INVX1_LOC_274/A INVX1_LOC_91/A 0.07fF
C2533 INVX1_LOC_10/A NOR2X1_LOC_48/B 0.21fF
C2534 NOR2X1_LOC_598/B NOR2X1_LOC_550/B 0.12fF
C2535 INVX1_LOC_64/A D_INPUT_2 0.05fF
C2536 NOR2X1_LOC_731/A NOR2X1_LOC_727/B 0.00fF
C2537 INVX1_LOC_208/A NOR2X1_LOC_334/Y 1.77fF
C2538 NAND2X1_LOC_231/Y NAND2X1_LOC_466/a_36_24# 0.06fF
C2539 NOR2X1_LOC_434/a_36_216# NOR2X1_LOC_798/A 0.00fF
C2540 INVX1_LOC_233/Y NOR2X1_LOC_625/Y 0.01fF
C2541 INPUT_6 NAND2X1_LOC_21/Y 0.29fF
C2542 NOR2X1_LOC_226/A NAND2X1_LOC_437/a_36_24# 0.00fF
C2543 INVX1_LOC_88/A INVX1_LOC_31/A 0.02fF
C2544 NOR2X1_LOC_516/B NOR2X1_LOC_334/Y 0.07fF
C2545 INVX1_LOC_279/A INVX1_LOC_32/A 0.14fF
C2546 INVX1_LOC_13/A NOR2X1_LOC_38/B 0.13fF
C2547 INVX1_LOC_13/Y INVX1_LOC_111/A 0.01fF
C2548 NOR2X1_LOC_52/B INVX1_LOC_29/Y 0.03fF
C2549 NOR2X1_LOC_405/A NAND2X1_LOC_93/B 0.03fF
C2550 NAND2X1_LOC_337/B NAND2X1_LOC_352/B 0.04fF
C2551 NOR2X1_LOC_346/B INVX1_LOC_26/Y 1.79fF
C2552 NAND2X1_LOC_303/Y NAND2X1_LOC_856/A 0.01fF
C2553 NOR2X1_LOC_707/A VDD -0.00fF
C2554 INVX1_LOC_168/A INVX1_LOC_23/A 0.19fF
C2555 NOR2X1_LOC_166/Y INVX1_LOC_102/A 0.04fF
C2556 NOR2X1_LOC_392/B NOR2X1_LOC_392/Y 0.06fF
C2557 NOR2X1_LOC_255/Y NOR2X1_LOC_84/Y 0.10fF
C2558 INVX1_LOC_14/Y NOR2X1_LOC_331/B 0.10fF
C2559 INVX1_LOC_73/Y INVX1_LOC_30/A 0.02fF
C2560 INVX1_LOC_14/A INVX1_LOC_72/A 0.06fF
C2561 NAND2X1_LOC_579/A NOR2X1_LOC_68/A 0.03fF
C2562 NOR2X1_LOC_780/A NOR2X1_LOC_783/A 0.08fF
C2563 VDD NOR2X1_LOC_709/B -0.00fF
C2564 NAND2X1_LOC_374/Y INVX1_LOC_57/A 0.07fF
C2565 INVX1_LOC_1/A NOR2X1_LOC_360/Y 0.17fF
C2566 INVX1_LOC_256/A NOR2X1_LOC_336/B 0.01fF
C2567 INVX1_LOC_50/A NAND2X1_LOC_200/B 0.00fF
C2568 VDD NOR2X1_LOC_209/B 0.14fF
C2569 INVX1_LOC_22/A INVX1_LOC_26/Y 0.04fF
C2570 INVX1_LOC_144/A NAND2X1_LOC_74/B 0.02fF
C2571 INVX1_LOC_298/Y NOR2X1_LOC_188/Y 0.18fF
C2572 INVX1_LOC_64/A NOR2X1_LOC_591/Y 0.02fF
C2573 INVX1_LOC_50/A NOR2X1_LOC_251/Y 0.01fF
C2574 NAND2X1_LOC_738/B NOR2X1_LOC_505/Y 0.02fF
C2575 NAND2X1_LOC_454/a_36_24# INVX1_LOC_307/A 0.00fF
C2576 INVX1_LOC_269/A INVX1_LOC_24/A 0.08fF
C2577 INVX1_LOC_64/A NOR2X1_LOC_529/Y 0.01fF
C2578 NAND2X1_LOC_552/A NAND2X1_LOC_357/B 0.00fF
C2579 INVX1_LOC_256/A NAND2X1_LOC_364/A 0.08fF
C2580 NOR2X1_LOC_58/a_36_216# INVX1_LOC_76/A 0.01fF
C2581 VDD INVX1_LOC_71/Y 0.21fF
C2582 NOR2X1_LOC_299/Y NOR2X1_LOC_395/Y 0.04fF
C2583 NAND2X1_LOC_662/Y INVX1_LOC_296/A 0.05fF
C2584 NOR2X1_LOC_51/A NOR2X1_LOC_425/Y 0.43fF
C2585 INVX1_LOC_225/Y INVX1_LOC_18/A 0.02fF
C2586 NAND2X1_LOC_116/A INVX1_LOC_50/Y 0.03fF
C2587 INVX1_LOC_89/A NAND2X1_LOC_223/A 0.02fF
C2588 NOR2X1_LOC_383/Y NOR2X1_LOC_72/Y -0.02fF
C2589 INVX1_LOC_182/Y INVX1_LOC_32/A 0.03fF
C2590 NOR2X1_LOC_643/Y NAND2X1_LOC_216/a_36_24# 0.00fF
C2591 INVX1_LOC_289/Y NOR2X1_LOC_753/Y 0.06fF
C2592 INVX1_LOC_16/A NOR2X1_LOC_696/Y 0.26fF
C2593 INVX1_LOC_286/A INVX1_LOC_12/A 0.07fF
C2594 NOR2X1_LOC_32/B INVX1_LOC_172/Y 0.03fF
C2595 INVX1_LOC_21/A NOR2X1_LOC_574/A 0.03fF
C2596 NOR2X1_LOC_533/Y NOR2X1_LOC_152/Y 0.03fF
C2597 INVX1_LOC_178/A NAND2X1_LOC_357/B 0.10fF
C2598 NOR2X1_LOC_841/A NAND2X1_LOC_453/A 0.11fF
C2599 NAND2X1_LOC_568/A NAND2X1_LOC_567/Y 0.03fF
C2600 NOR2X1_LOC_441/Y NAND2X1_LOC_545/a_36_24# 0.01fF
C2601 INVX1_LOC_17/A INVX1_LOC_77/A 0.14fF
C2602 NOR2X1_LOC_524/Y INVX1_LOC_223/A 0.09fF
C2603 NAND2X1_LOC_267/B NAND2X1_LOC_572/B 0.02fF
C2604 INVX1_LOC_13/Y NOR2X1_LOC_290/Y 0.04fF
C2605 INVX1_LOC_28/A NAND2X1_LOC_471/Y 0.02fF
C2606 NOR2X1_LOC_361/B NOR2X1_LOC_716/B 0.10fF
C2607 INVX1_LOC_5/A NAND2X1_LOC_549/B 0.01fF
C2608 NAND2X1_LOC_802/A NAND2X1_LOC_799/A 0.38fF
C2609 INVX1_LOC_35/A INVX1_LOC_151/Y 0.01fF
C2610 NOR2X1_LOC_849/a_36_216# NOR2X1_LOC_500/B 0.00fF
C2611 NOR2X1_LOC_859/Y NOR2X1_LOC_862/B 0.01fF
C2612 INVX1_LOC_269/A NOR2X1_LOC_557/Y 0.10fF
C2613 INVX1_LOC_233/A NAND2X1_LOC_170/A 0.00fF
C2614 NOR2X1_LOC_536/Y NAND2X1_LOC_811/Y 0.01fF
C2615 INVX1_LOC_80/A INVX1_LOC_23/A 0.05fF
C2616 NOR2X1_LOC_710/B INVX1_LOC_33/A 0.40fF
C2617 INVX1_LOC_161/Y NOR2X1_LOC_577/Y 0.31fF
C2618 INVX1_LOC_299/A INVX1_LOC_149/Y 0.00fF
C2619 NOR2X1_LOC_471/Y INVX1_LOC_77/A 2.07fF
C2620 INVX1_LOC_58/A NAND2X1_LOC_656/Y 0.01fF
C2621 INVX1_LOC_30/A NOR2X1_LOC_91/Y 0.80fF
C2622 INVX1_LOC_12/Y NOR2X1_LOC_813/a_36_216# 0.01fF
C2623 NAND2X1_LOC_231/Y NOR2X1_LOC_321/Y 0.10fF
C2624 INVX1_LOC_303/A INVX1_LOC_31/A 0.07fF
C2625 NOR2X1_LOC_45/B NOR2X1_LOC_754/A 0.03fF
C2626 NAND2X1_LOC_8/a_36_24# NOR2X1_LOC_814/A 0.01fF
C2627 NAND2X1_LOC_739/B INVX1_LOC_72/A 0.01fF
C2628 NOR2X1_LOC_160/B NOR2X1_LOC_162/Y 0.00fF
C2629 INVX1_LOC_136/A INVX1_LOC_94/A 0.10fF
C2630 NAND2X1_LOC_218/B NAND2X1_LOC_672/a_36_24# 0.00fF
C2631 NOR2X1_LOC_238/a_36_216# INVX1_LOC_217/A 0.06fF
C2632 INVX1_LOC_1/A NAND2X1_LOC_451/Y 0.02fF
C2633 INVX1_LOC_137/Y INVX1_LOC_306/Y 0.01fF
C2634 INVX1_LOC_135/A INVX1_LOC_138/A 0.01fF
C2635 INVX1_LOC_216/Y NAND2X1_LOC_141/A 0.01fF
C2636 NAND2X1_LOC_858/B NAND2X1_LOC_175/Y 0.04fF
C2637 NOR2X1_LOC_361/B INVX1_LOC_98/Y 0.04fF
C2638 INVX1_LOC_14/A NAND2X1_LOC_338/B 1.33fF
C2639 INVX1_LOC_12/Y NAND2X1_LOC_773/B 0.10fF
C2640 NOR2X1_LOC_144/a_36_216# INVX1_LOC_4/A 0.00fF
C2641 NAND2X1_LOC_357/B NOR2X1_LOC_816/A 0.07fF
C2642 NOR2X1_LOC_88/Y INVX1_LOC_185/A 0.03fF
C2643 NOR2X1_LOC_638/a_36_216# INVX1_LOC_72/A -0.02fF
C2644 NAND2X1_LOC_387/B INVX1_LOC_49/A 0.02fF
C2645 NAND2X1_LOC_652/Y INVX1_LOC_271/A 0.02fF
C2646 INVX1_LOC_90/A NOR2X1_LOC_392/Y 0.07fF
C2647 NOR2X1_LOC_644/A INVX1_LOC_53/A 0.07fF
C2648 NOR2X1_LOC_479/B NOR2X1_LOC_15/Y 0.02fF
C2649 NOR2X1_LOC_590/A INVX1_LOC_104/A 0.19fF
C2650 INVX1_LOC_106/A INVX1_LOC_37/A 0.05fF
C2651 NAND2X1_LOC_149/Y GATE_479 0.01fF
C2652 NOR2X1_LOC_328/Y NOR2X1_LOC_15/Y 0.03fF
C2653 INVX1_LOC_201/Y INVX1_LOC_40/Y 0.02fF
C2654 NOR2X1_LOC_67/A NOR2X1_LOC_82/A 0.15fF
C2655 NOR2X1_LOC_828/B INVX1_LOC_53/A 0.00fF
C2656 INVX1_LOC_116/A NOR2X1_LOC_303/Y 0.03fF
C2657 INVX1_LOC_39/A INVX1_LOC_135/A 0.03fF
C2658 INVX1_LOC_185/A INVX1_LOC_84/A 0.03fF
C2659 NAND2X1_LOC_796/B NOR2X1_LOC_312/Y 0.03fF
C2660 NAND2X1_LOC_843/a_36_24# INVX1_LOC_94/Y 0.01fF
C2661 NOR2X1_LOC_559/B NAND2X1_LOC_517/a_36_24# 0.02fF
C2662 INVX1_LOC_37/Y NAND2X1_LOC_254/Y 0.01fF
C2663 NAND2X1_LOC_348/A NOR2X1_LOC_392/Y 0.42fF
C2664 INVX1_LOC_11/A NOR2X1_LOC_160/Y 0.03fF
C2665 NOR2X1_LOC_530/Y INVX1_LOC_316/Y 0.15fF
C2666 INVX1_LOC_161/Y INVX1_LOC_22/A 0.20fF
C2667 INVX1_LOC_34/A NOR2X1_LOC_607/A 0.09fF
C2668 INVX1_LOC_72/A NOR2X1_LOC_612/B 0.10fF
C2669 INVX1_LOC_18/A INVX1_LOC_266/Y 0.11fF
C2670 INVX1_LOC_226/Y INVX1_LOC_218/Y 0.01fF
C2671 NOR2X1_LOC_457/A NOR2X1_LOC_543/A 0.24fF
C2672 INVX1_LOC_50/A NOR2X1_LOC_528/Y 0.53fF
C2673 NAND2X1_LOC_726/Y NAND2X1_LOC_711/Y 0.04fF
C2674 NOR2X1_LOC_124/A INVX1_LOC_23/Y 0.02fF
C2675 NAND2X1_LOC_785/Y NOR2X1_LOC_238/Y 0.02fF
C2676 NOR2X1_LOC_334/Y NAND2X1_LOC_211/Y 0.03fF
C2677 INVX1_LOC_12/A INVX1_LOC_54/A 7.36fF
C2678 INVX1_LOC_72/Y INVX1_LOC_34/Y 0.11fF
C2679 NOR2X1_LOC_609/A INVX1_LOC_177/A 0.01fF
C2680 NOR2X1_LOC_468/Y NAND2X1_LOC_551/A 0.02fF
C2681 INVX1_LOC_278/A NOR2X1_LOC_368/a_36_216# 0.00fF
C2682 NAND2X1_LOC_350/A INVX1_LOC_10/A 0.23fF
C2683 INVX1_LOC_178/A NAND2X1_LOC_849/A 0.01fF
C2684 NOR2X1_LOC_599/A INVX1_LOC_22/A 0.05fF
C2685 INVX1_LOC_116/A INVX1_LOC_54/Y 0.01fF
C2686 NAND2X1_LOC_190/Y INVX1_LOC_55/Y 0.07fF
C2687 NOR2X1_LOC_795/Y INVX1_LOC_49/A 0.03fF
C2688 INVX1_LOC_90/A NAND2X1_LOC_357/A 0.01fF
C2689 NAND2X1_LOC_20/B INVX1_LOC_20/Y 0.02fF
C2690 INVX1_LOC_80/A INVX1_LOC_31/A 0.03fF
C2691 NOR2X1_LOC_433/A NOR2X1_LOC_361/Y 0.03fF
C2692 INVX1_LOC_139/Y NOR2X1_LOC_631/Y 0.00fF
C2693 INVX1_LOC_1/A NOR2X1_LOC_567/B 0.07fF
C2694 NOR2X1_LOC_693/Y INVX1_LOC_46/A 0.05fF
C2695 INVX1_LOC_13/Y INVX1_LOC_6/A 0.03fF
C2696 NAND2X1_LOC_563/A INVX1_LOC_24/A 0.01fF
C2697 NAND2X1_LOC_288/B INVX1_LOC_46/A 0.11fF
C2698 NOR2X1_LOC_101/a_36_216# INVX1_LOC_42/A 0.00fF
C2699 NOR2X1_LOC_246/A NOR2X1_LOC_389/A 0.02fF
C2700 NOR2X1_LOC_831/B INVX1_LOC_42/A 0.70fF
C2701 NAND2X1_LOC_465/a_36_24# NAND2X1_LOC_773/B 0.00fF
C2702 NOR2X1_LOC_788/B INVX1_LOC_292/A 0.02fF
C2703 INVX1_LOC_181/Y INVX1_LOC_1/Y 0.03fF
C2704 NOR2X1_LOC_301/a_36_216# NOR2X1_LOC_438/Y 0.00fF
C2705 INVX1_LOC_91/A INVX1_LOC_306/Y 0.10fF
C2706 INVX1_LOC_186/Y INVX1_LOC_19/A 0.07fF
C2707 NOR2X1_LOC_863/Y NOR2X1_LOC_863/B 0.02fF
C2708 INVX1_LOC_13/A INVX1_LOC_62/Y 0.01fF
C2709 INVX1_LOC_278/Y NOR2X1_LOC_753/Y 0.07fF
C2710 INVX1_LOC_227/A INVX1_LOC_177/Y 0.17fF
C2711 INVX1_LOC_48/A NAND2X1_LOC_85/a_36_24# 0.00fF
C2712 NOR2X1_LOC_219/Y NOR2X1_LOC_219/a_36_216# 0.01fF
C2713 NOR2X1_LOC_727/B INVX1_LOC_117/A 0.05fF
C2714 INVX1_LOC_209/Y NAND2X1_LOC_853/Y 0.00fF
C2715 INVX1_LOC_33/A NOR2X1_LOC_524/a_36_216# 0.00fF
C2716 NOR2X1_LOC_315/Y NOR2X1_LOC_316/Y 0.00fF
C2717 INVX1_LOC_232/Y NAND2X1_LOC_139/A 0.02fF
C2718 NOR2X1_LOC_777/B INVX1_LOC_19/A 0.07fF
C2719 NOR2X1_LOC_19/B INVX1_LOC_61/Y 0.00fF
C2720 NOR2X1_LOC_705/B INVX1_LOC_75/A 0.03fF
C2721 INVX1_LOC_214/A NOR2X1_LOC_574/A 0.16fF
C2722 INVX1_LOC_88/A INVX1_LOC_6/A 0.03fF
C2723 INPUT_0 NAND2X1_LOC_793/Y 0.01fF
C2724 NAND2X1_LOC_386/a_36_24# INVX1_LOC_89/A 0.00fF
C2725 INVX1_LOC_90/A NOR2X1_LOC_86/Y 0.00fF
C2726 INVX1_LOC_54/A NOR2X1_LOC_686/A 0.01fF
C2727 NAND2X1_LOC_357/B NOR2X1_LOC_773/Y 0.15fF
C2728 NOR2X1_LOC_92/Y INVX1_LOC_70/Y 0.03fF
C2729 NOR2X1_LOC_703/B NOR2X1_LOC_356/A 0.01fF
C2730 NOR2X1_LOC_75/Y INVX1_LOC_285/Y 0.00fF
C2731 INVX1_LOC_200/A INVX1_LOC_286/A 0.00fF
C2732 INVX1_LOC_251/Y NOR2X1_LOC_226/A 0.15fF
C2733 INVX1_LOC_78/A NOR2X1_LOC_831/B 0.42fF
C2734 NAND2X1_LOC_326/A NOR2X1_LOC_595/Y 0.01fF
C2735 INVX1_LOC_90/A NOR2X1_LOC_744/a_36_216# 0.00fF
C2736 NOR2X1_LOC_716/B NAND2X1_LOC_573/A 0.02fF
C2737 NAND2X1_LOC_206/B INVX1_LOC_29/A 0.01fF
C2738 NOR2X1_LOC_355/A NOR2X1_LOC_433/A 0.01fF
C2739 INVX1_LOC_255/Y INVX1_LOC_80/Y 0.03fF
C2740 NOR2X1_LOC_222/a_36_216# NOR2X1_LOC_52/B 0.00fF
C2741 NAND2X1_LOC_21/a_36_24# INVX1_LOC_140/A 0.01fF
C2742 NAND2X1_LOC_854/B NAND2X1_LOC_354/B 0.00fF
C2743 INVX1_LOC_55/Y NOR2X1_LOC_596/A 0.07fF
C2744 NAND2X1_LOC_181/Y INVX1_LOC_256/Y 0.01fF
C2745 NOR2X1_LOC_142/Y INVX1_LOC_10/A 0.01fF
C2746 INVX1_LOC_21/A NOR2X1_LOC_305/Y 0.02fF
C2747 NOR2X1_LOC_458/Y NOR2X1_LOC_717/B -0.01fF
C2748 INVX1_LOC_12/A NOR2X1_LOC_48/B 0.15fF
C2749 NOR2X1_LOC_677/Y INVX1_LOC_291/A 0.01fF
C2750 VDD NOR2X1_LOC_343/B -0.00fF
C2751 INVX1_LOC_226/Y NOR2X1_LOC_655/B 0.10fF
C2752 INVX1_LOC_138/A INVX1_LOC_280/A 0.03fF
C2753 NOR2X1_LOC_519/Y NOR2X1_LOC_48/B 0.06fF
C2754 INVX1_LOC_285/A NOR2X1_LOC_281/a_36_216# 0.00fF
C2755 INVX1_LOC_136/A INVX1_LOC_144/A 0.10fF
C2756 NOR2X1_LOC_65/B NOR2X1_LOC_831/B 0.01fF
C2757 NOR2X1_LOC_750/a_36_216# NAND2X1_LOC_656/A 0.11fF
C2758 INVX1_LOC_89/A INVX1_LOC_33/A 1.23fF
C2759 INVX1_LOC_227/A INVX1_LOC_104/A 1.07fF
C2760 INVX1_LOC_35/A INVX1_LOC_118/Y 0.02fF
C2761 NOR2X1_LOC_96/Y NOR2X1_LOC_392/Y 0.02fF
C2762 NOR2X1_LOC_703/B NOR2X1_LOC_74/A 2.11fF
C2763 INVX1_LOC_256/A NOR2X1_LOC_405/A 0.38fF
C2764 NOR2X1_LOC_336/B INVX1_LOC_69/Y 0.01fF
C2765 INVX1_LOC_217/A NOR2X1_LOC_754/a_36_216# 0.01fF
C2766 NOR2X1_LOC_134/Y NOR2X1_LOC_45/B 0.05fF
C2767 INVX1_LOC_164/A NOR2X1_LOC_84/Y 0.03fF
C2768 NOR2X1_LOC_622/A NOR2X1_LOC_624/B 0.06fF
C2769 INVX1_LOC_39/A NOR2X1_LOC_813/Y 0.07fF
C2770 D_INPUT_1 NAND2X1_LOC_817/a_36_24# 0.00fF
C2771 NOR2X1_LOC_20/Y NOR2X1_LOC_24/Y 0.00fF
C2772 NOR2X1_LOC_355/A NOR2X1_LOC_52/B 0.10fF
C2773 NOR2X1_LOC_360/Y NOR2X1_LOC_188/A 0.26fF
C2774 INVX1_LOC_201/Y NAND2X1_LOC_28/a_36_24# 0.00fF
C2775 NOR2X1_LOC_589/A NOR2X1_LOC_191/A 0.06fF
C2776 INVX1_LOC_41/A INVX1_LOC_87/Y 0.01fF
C2777 INVX1_LOC_64/A NOR2X1_LOC_61/Y 0.01fF
C2778 NOR2X1_LOC_394/Y NAND2X1_LOC_81/B 0.06fF
C2779 NOR2X1_LOC_717/B INVX1_LOC_177/A 0.00fF
C2780 INVX1_LOC_39/A INVX1_LOC_280/A 0.03fF
C2781 NOR2X1_LOC_609/A INVX1_LOC_285/Y 0.01fF
C2782 NAND2X1_LOC_848/Y NOR2X1_LOC_392/Y -0.03fF
C2783 NAND2X1_LOC_734/a_36_24# NAND2X1_LOC_807/Y 0.01fF
C2784 INVX1_LOC_39/A NOR2X1_LOC_94/Y 0.00fF
C2785 NAND2X1_LOC_734/B INVX1_LOC_90/A 0.01fF
C2786 INVX1_LOC_130/A NOR2X1_LOC_657/B 0.04fF
C2787 INVX1_LOC_30/Y INVX1_LOC_232/A 0.05fF
C2788 NOR2X1_LOC_67/A INVX1_LOC_306/A 0.03fF
C2789 INVX1_LOC_36/A NOR2X1_LOC_139/Y 0.02fF
C2790 INVX1_LOC_256/A NOR2X1_LOC_857/A 0.07fF
C2791 INVX1_LOC_36/A NAND2X1_LOC_655/A 0.07fF
C2792 INVX1_LOC_5/A NOR2X1_LOC_78/a_36_216# 0.00fF
C2793 INVX1_LOC_282/A NAND2X1_LOC_631/a_36_24# 0.00fF
C2794 NOR2X1_LOC_78/B NOR2X1_LOC_71/Y 0.07fF
C2795 INVX1_LOC_122/Y NOR2X1_LOC_78/A 0.28fF
C2796 INVX1_LOC_35/A NOR2X1_LOC_240/A 0.01fF
C2797 NOR2X1_LOC_458/Y NOR2X1_LOC_151/Y 0.01fF
C2798 INVX1_LOC_13/Y NOR2X1_LOC_79/A 0.15fF
C2799 NOR2X1_LOC_151/Y INVX1_LOC_153/Y 0.03fF
C2800 INVX1_LOC_11/A NOR2X1_LOC_111/A 0.10fF
C2801 NOR2X1_LOC_705/B NAND2X1_LOC_485/a_36_24# 0.02fF
C2802 INVX1_LOC_104/A NOR2X1_LOC_703/A 0.01fF
C2803 INVX1_LOC_24/A NOR2X1_LOC_741/A 0.01fF
C2804 NOR2X1_LOC_582/Y NOR2X1_LOC_588/A 0.14fF
C2805 INVX1_LOC_26/Y NOR2X1_LOC_777/B 0.08fF
C2806 INVX1_LOC_30/Y NOR2X1_LOC_383/Y 0.02fF
C2807 NAND2X1_LOC_357/B INVX1_LOC_140/A 0.10fF
C2808 NOR2X1_LOC_389/A NOR2X1_LOC_357/Y 0.10fF
C2809 INVX1_LOC_211/Y NOR2X1_LOC_447/B 0.86fF
C2810 NOR2X1_LOC_448/B INVX1_LOC_38/A 0.02fF
C2811 NOR2X1_LOC_392/B INVX1_LOC_75/A 0.10fF
C2812 INVX1_LOC_36/A NAND2X1_LOC_468/B 0.03fF
C2813 NAND2X1_LOC_536/a_36_24# INVX1_LOC_222/A 0.01fF
C2814 INVX1_LOC_84/A NOR2X1_LOC_754/Y 0.00fF
C2815 INVX1_LOC_32/A NOR2X1_LOC_38/B 1.21fF
C2816 INVX1_LOC_89/A INVX1_LOC_40/A 0.15fF
C2817 NOR2X1_LOC_78/B NOR2X1_LOC_644/A 0.08fF
C2818 INVX1_LOC_255/Y INVX1_LOC_83/A 0.01fF
C2819 INVX1_LOC_135/A NAND2X1_LOC_735/B 0.03fF
C2820 INVX1_LOC_181/Y INVX1_LOC_93/Y 0.91fF
C2821 INVX1_LOC_90/A INVX1_LOC_25/Y 0.00fF
C2822 INVX1_LOC_17/A INVX1_LOC_9/A 0.21fF
C2823 INVX1_LOC_23/A INVX1_LOC_272/A 0.39fF
C2824 NAND2X1_LOC_7/Y NOR2X1_LOC_78/A 0.01fF
C2825 NOR2X1_LOC_609/A NOR2X1_LOC_137/B 0.05fF
C2826 INVX1_LOC_48/Y NOR2X1_LOC_235/Y 0.04fF
C2827 INVX1_LOC_49/A NOR2X1_LOC_45/B 0.14fF
C2828 NOR2X1_LOC_389/B INVX1_LOC_25/Y 0.12fF
C2829 NOR2X1_LOC_84/Y NOR2X1_LOC_368/A 0.12fF
C2830 NOR2X1_LOC_456/Y INVX1_LOC_29/A 0.21fF
C2831 INVX1_LOC_14/A NAND2X1_LOC_444/a_36_24# 0.00fF
C2832 NOR2X1_LOC_128/B NOR2X1_LOC_332/A 0.01fF
C2833 INVX1_LOC_81/A NOR2X1_LOC_657/B 0.06fF
C2834 NOR2X1_LOC_598/B NAND2X1_LOC_74/B 0.12fF
C2835 NOR2X1_LOC_739/Y INVX1_LOC_274/A 0.00fF
C2836 INVX1_LOC_134/A NOR2X1_LOC_729/A 0.21fF
C2837 INVX1_LOC_200/A INVX1_LOC_54/A 0.18fF
C2838 NOR2X1_LOC_598/B NAND2X1_LOC_207/Y 0.02fF
C2839 INVX1_LOC_27/A NAND2X1_LOC_235/a_36_24# 0.00fF
C2840 INVX1_LOC_1/A NOR2X1_LOC_79/Y 0.08fF
C2841 NOR2X1_LOC_564/a_36_216# INVX1_LOC_104/A 0.00fF
C2842 INVX1_LOC_269/A NOR2X1_LOC_197/B 0.10fF
C2843 NOR2X1_LOC_596/A NOR2X1_LOC_357/Y 0.05fF
C2844 NOR2X1_LOC_714/Y NOR2X1_LOC_703/Y 0.13fF
C2845 NAND2X1_LOC_740/B INVX1_LOC_16/A 0.06fF
C2846 NAND2X1_LOC_348/A INVX1_LOC_25/Y 0.01fF
C2847 NOR2X1_LOC_256/Y INVX1_LOC_16/A 0.06fF
C2848 NOR2X1_LOC_92/Y INVX1_LOC_285/A 0.57fF
C2849 INVX1_LOC_269/A NAND2X1_LOC_237/a_36_24# 0.00fF
C2850 INVX1_LOC_48/A NOR2X1_LOC_537/Y 0.07fF
C2851 INVX1_LOC_11/A NOR2X1_LOC_600/a_36_216# 0.01fF
C2852 NAND2X1_LOC_363/B NOR2X1_LOC_461/Y 0.03fF
C2853 INVX1_LOC_268/A NAND2X1_LOC_51/B 0.02fF
C2854 NOR2X1_LOC_317/A NOR2X1_LOC_319/B 0.00fF
C2855 NAND2X1_LOC_733/Y INVX1_LOC_54/A 0.20fF
C2856 NOR2X1_LOC_332/A NOR2X1_LOC_702/Y 0.16fF
C2857 NOR2X1_LOC_137/A INVX1_LOC_313/Y 0.00fF
C2858 NOR2X1_LOC_192/a_36_216# INVX1_LOC_93/Y 0.01fF
C2859 INVX1_LOC_61/A NOR2X1_LOC_813/Y 0.03fF
C2860 NOR2X1_LOC_307/A NOR2X1_LOC_155/A 0.03fF
C2861 INVX1_LOC_24/A INVX1_LOC_12/Y 0.98fF
C2862 INVX1_LOC_88/A NOR2X1_LOC_117/Y 0.29fF
C2863 NOR2X1_LOC_357/a_36_216# INVX1_LOC_78/Y 0.00fF
C2864 INVX1_LOC_286/A NOR2X1_LOC_566/Y 0.03fF
C2865 INVX1_LOC_24/Y NOR2X1_LOC_814/A 0.10fF
C2866 INVX1_LOC_2/A NOR2X1_LOC_45/B 6.19fF
C2867 NOR2X1_LOC_716/B NAND2X1_LOC_267/B 0.03fF
C2868 NOR2X1_LOC_6/B INVX1_LOC_74/Y 0.06fF
C2869 NOR2X1_LOC_520/B INVX1_LOC_176/A 0.02fF
C2870 NOR2X1_LOC_828/B INVX1_LOC_83/A 0.03fF
C2871 NAND2X1_LOC_564/B NAND2X1_LOC_858/B 0.00fF
C2872 NOR2X1_LOC_276/Y NOR2X1_LOC_155/A 0.05fF
C2873 INVX1_LOC_61/A INVX1_LOC_280/A 0.60fF
C2874 NOR2X1_LOC_172/Y NAND2X1_LOC_453/A 0.01fF
C2875 INVX1_LOC_314/Y NAND2X1_LOC_230/a_36_24# 0.00fF
C2876 NOR2X1_LOC_226/A NOR2X1_LOC_45/B 0.14fF
C2877 NOR2X1_LOC_667/Y NOR2X1_LOC_88/Y 0.01fF
C2878 NAND2X1_LOC_833/Y INVX1_LOC_37/A 0.06fF
C2879 INVX1_LOC_13/A INVX1_LOC_51/Y 0.02fF
C2880 NOR2X1_LOC_272/Y NOR2X1_LOC_89/A 0.03fF
C2881 NOR2X1_LOC_388/Y INVX1_LOC_14/Y 0.10fF
C2882 NOR2X1_LOC_678/A INVX1_LOC_4/A 0.03fF
C2883 INVX1_LOC_217/A INVX1_LOC_54/A 0.14fF
C2884 NOR2X1_LOC_843/B INVX1_LOC_26/Y 0.03fF
C2885 NAND2X1_LOC_364/Y INVX1_LOC_117/A 2.10fF
C2886 NOR2X1_LOC_789/B INVX1_LOC_42/A 0.01fF
C2887 NAND2X1_LOC_9/Y INVX1_LOC_165/A 0.01fF
C2888 D_INPUT_4 D_GATE_366 0.06fF
C2889 INVX1_LOC_90/A INVX1_LOC_75/A 0.18fF
C2890 NOR2X1_LOC_78/B NOR2X1_LOC_540/B 0.02fF
C2891 NAND2X1_LOC_74/B NOR2X1_LOC_271/a_36_216# 0.00fF
C2892 INVX1_LOC_25/A INVX1_LOC_26/A 0.07fF
C2893 NOR2X1_LOC_392/Y NAND2X1_LOC_223/A 0.07fF
C2894 NOR2X1_LOC_67/A INVX1_LOC_59/Y 0.10fF
C2895 INVX1_LOC_136/A NOR2X1_LOC_155/A 0.04fF
C2896 NOR2X1_LOC_796/B INVX1_LOC_301/A 0.14fF
C2897 NOR2X1_LOC_504/Y NOR2X1_LOC_422/Y -0.00fF
C2898 NAND2X1_LOC_149/B INVX1_LOC_91/A 0.01fF
C2899 INVX1_LOC_227/A INVX1_LOC_206/Y 0.01fF
C2900 INVX1_LOC_183/Y NOR2X1_LOC_74/A 0.01fF
C2901 NOR2X1_LOC_389/B INVX1_LOC_75/A 0.07fF
C2902 NOR2X1_LOC_52/B NOR2X1_LOC_111/A 0.10fF
C2903 INVX1_LOC_40/Y NAND2X1_LOC_574/A 0.01fF
C2904 NOR2X1_LOC_160/B NAND2X1_LOC_773/B 0.07fF
C2905 NOR2X1_LOC_679/Y INVX1_LOC_49/Y 0.22fF
C2906 NOR2X1_LOC_627/a_36_216# INVX1_LOC_139/Y 0.00fF
C2907 NOR2X1_LOC_401/Y NOR2X1_LOC_266/B 0.00fF
C2908 INVX1_LOC_282/A NOR2X1_LOC_497/Y 0.07fF
C2909 NOR2X1_LOC_667/A NOR2X1_LOC_305/Y 0.07fF
C2910 NAND2X1_LOC_30/Y NOR2X1_LOC_1/Y 0.04fF
C2911 INVX1_LOC_248/A NOR2X1_LOC_305/Y 0.74fF
C2912 NOR2X1_LOC_220/A NOR2X1_LOC_357/Y 0.03fF
C2913 NAND2X1_LOC_787/B INVX1_LOC_54/A 0.01fF
C2914 INVX1_LOC_36/A NOR2X1_LOC_820/B 0.02fF
C2915 NAND2X1_LOC_348/A INVX1_LOC_75/A 0.03fF
C2916 NAND2X1_LOC_350/A INVX1_LOC_12/A 0.12fF
C2917 INVX1_LOC_30/Y NAND2X1_LOC_447/Y 0.00fF
C2918 NOR2X1_LOC_468/Y INVX1_LOC_32/A 0.10fF
C2919 INVX1_LOC_17/A NOR2X1_LOC_861/Y 0.25fF
C2920 INVX1_LOC_2/A INVX1_LOC_281/A 0.02fF
C2921 INVX1_LOC_21/A INVX1_LOC_271/Y 0.07fF
C2922 NOR2X1_LOC_258/a_36_216# NOR2X1_LOC_89/A 0.00fF
C2923 NOR2X1_LOC_93/a_36_216# INVX1_LOC_280/A 0.00fF
C2924 INVX1_LOC_49/A NOR2X1_LOC_862/B 0.32fF
C2925 NAND2X1_LOC_190/Y INVX1_LOC_32/A 0.03fF
C2926 NOR2X1_LOC_186/Y NOR2X1_LOC_278/Y 0.21fF
C2927 INVX1_LOC_45/A INVX1_LOC_262/Y 0.01fF
C2928 NOR2X1_LOC_82/A NAND2X1_LOC_445/a_36_24# 0.01fF
C2929 INVX1_LOC_34/A NOR2X1_LOC_433/Y 0.05fF
C2930 NOR2X1_LOC_45/B INPUT_1 0.06fF
C2931 NOR2X1_LOC_52/B INVX1_LOC_127/A 0.00fF
C2932 NOR2X1_LOC_441/Y INVX1_LOC_12/A 0.00fF
C2933 INVX1_LOC_208/A NAND2X1_LOC_472/Y 0.10fF
C2934 NOR2X1_LOC_598/B INVX1_LOC_259/Y 0.02fF
C2935 INVX1_LOC_33/Y NAND2X1_LOC_840/B 0.00fF
C2936 INVX1_LOC_304/Y INVX1_LOC_54/A 0.03fF
C2937 NOR2X1_LOC_577/Y NOR2X1_LOC_841/A 0.10fF
C2938 NOR2X1_LOC_356/A INVX1_LOC_91/A 0.09fF
C2939 NOR2X1_LOC_500/B NOR2X1_LOC_633/A 0.01fF
C2940 NOR2X1_LOC_208/Y NOR2X1_LOC_66/Y 0.03fF
C2941 NAND2X1_LOC_396/a_36_24# INVX1_LOC_32/A 0.06fF
C2942 NAND2X1_LOC_361/Y NAND2X1_LOC_412/a_36_24# 0.00fF
C2943 INVX1_LOC_18/A INVX1_LOC_19/A 0.71fF
C2944 NOR2X1_LOC_71/Y NOR2X1_LOC_368/Y 0.06fF
C2945 NOR2X1_LOC_516/B NAND2X1_LOC_472/Y 0.13fF
C2946 INVX1_LOC_89/A NOR2X1_LOC_486/Y 0.05fF
C2947 NAND2X1_LOC_573/Y NOR2X1_LOC_278/Y 0.07fF
C2948 NOR2X1_LOC_840/Y NOR2X1_LOC_840/A 0.10fF
C2949 NOR2X1_LOC_222/Y NOR2X1_LOC_142/a_36_216# 0.00fF
C2950 NOR2X1_LOC_391/A VDD 0.01fF
C2951 NAND2X1_LOC_466/Y NOR2X1_LOC_592/B 0.09fF
C2952 NOR2X1_LOC_561/A INVX1_LOC_25/Y 0.18fF
C2953 NAND2X1_LOC_35/B NOR2X1_LOC_629/Y 0.00fF
C2954 NOR2X1_LOC_218/Y INVX1_LOC_281/A 0.05fF
C2955 NOR2X1_LOC_598/B NAND2X1_LOC_358/B 0.01fF
C2956 INVX1_LOC_50/A INVX1_LOC_93/A 0.02fF
C2957 NOR2X1_LOC_813/Y NOR2X1_LOC_85/a_36_216# 0.01fF
C2958 INVX1_LOC_248/A NAND2X1_LOC_600/a_36_24# 0.00fF
C2959 NOR2X1_LOC_372/a_36_216# INVX1_LOC_42/A 0.01fF
C2960 NOR2X1_LOC_242/A NAND2X1_LOC_246/a_36_24# 0.00fF
C2961 INVX1_LOC_64/A NOR2X1_LOC_678/A 0.68fF
C2962 INVX1_LOC_135/A D_GATE_479 0.02fF
C2963 INVX1_LOC_214/Y INVX1_LOC_54/A 0.03fF
C2964 INVX1_LOC_135/A D_INPUT_3 0.24fF
C2965 INVX1_LOC_1/A INVX1_LOC_26/A 0.03fF
C2966 NAND2X1_LOC_364/A NOR2X1_LOC_89/A 2.23fF
C2967 NOR2X1_LOC_15/Y INVX1_LOC_23/Y 0.07fF
C2968 NOR2X1_LOC_718/a_36_216# INVX1_LOC_179/A 0.00fF
C2969 NOR2X1_LOC_71/Y INVX1_LOC_46/A 0.01fF
C2970 INPUT_3 NOR2X1_LOC_38/B 0.57fF
C2971 NAND2X1_LOC_349/B INVX1_LOC_38/A 0.08fF
C2972 INVX1_LOC_5/A NAND2X1_LOC_549/Y 0.00fF
C2973 NOR2X1_LOC_218/A NAND2X1_LOC_454/Y 0.02fF
C2974 INVX1_LOC_41/A NOR2X1_LOC_814/A 0.11fF
C2975 NAND2X1_LOC_735/B INVX1_LOC_280/A 0.81fF
C2976 NOR2X1_LOC_74/A INVX1_LOC_91/A 0.81fF
C2977 NAND2X1_LOC_231/Y NAND2X1_LOC_798/B 0.19fF
C2978 NOR2X1_LOC_68/A NOR2X1_LOC_470/a_36_216# 0.00fF
C2979 NOR2X1_LOC_655/B INVX1_LOC_307/A 0.01fF
C2980 INVX1_LOC_90/A NAND2X1_LOC_485/a_36_24# 0.00fF
C2981 NOR2X1_LOC_130/A INVX1_LOC_12/Y 0.02fF
C2982 INVX1_LOC_90/A NAND2X1_LOC_453/A 0.07fF
C2983 INVX1_LOC_217/A NOR2X1_LOC_48/B 0.03fF
C2984 NOR2X1_LOC_400/B INVX1_LOC_14/A 0.04fF
C2985 NAND2X1_LOC_477/A INVX1_LOC_285/A 0.10fF
C2986 NOR2X1_LOC_644/A INVX1_LOC_46/A 0.03fF
C2987 INVX1_LOC_5/A INVX1_LOC_213/A 0.27fF
C2988 NOR2X1_LOC_180/B INVX1_LOC_37/A 0.12fF
C2989 NAND2X1_LOC_795/Y NOR2X1_LOC_692/Y 0.06fF
C2990 NOR2X1_LOC_9/Y INVX1_LOC_91/A 0.23fF
C2991 NOR2X1_LOC_550/B INVX1_LOC_29/A 0.01fF
C2992 NOR2X1_LOC_716/B NAND2X1_LOC_81/B 0.07fF
C2993 INVX1_LOC_88/A INVX1_LOC_270/A 0.12fF
C2994 INVX1_LOC_23/A INVX1_LOC_198/A 0.00fF
C2995 INVX1_LOC_224/Y INVX1_LOC_14/A 1.48fF
C2996 NAND2X1_LOC_51/B INVX1_LOC_187/Y 0.07fF
C2997 INVX1_LOC_23/A NOR2X1_LOC_271/B 0.01fF
C2998 NOR2X1_LOC_199/B INVX1_LOC_9/A 0.06fF
C2999 INVX1_LOC_316/Y NOR2X1_LOC_104/a_36_216# 0.00fF
C3000 NAND2X1_LOC_538/Y INVX1_LOC_57/A 0.07fF
C3001 INVX1_LOC_135/A INVX1_LOC_230/A 0.01fF
C3002 NAND2X1_LOC_632/B INVX1_LOC_284/A 0.01fF
C3003 INVX1_LOC_62/Y INVX1_LOC_32/A 0.07fF
C3004 NAND2X1_LOC_38/a_36_24# INVX1_LOC_14/A 0.01fF
C3005 NOR2X1_LOC_740/Y INVX1_LOC_23/A 0.98fF
C3006 NAND2X1_LOC_364/A INVX1_LOC_104/Y 0.01fF
C3007 NAND2X1_LOC_593/Y NOR2X1_LOC_677/a_36_216# 0.00fF
C3008 NOR2X1_LOC_142/Y INVX1_LOC_12/A 0.07fF
C3009 NAND2X1_LOC_123/Y NOR2X1_LOC_363/Y 0.03fF
C3010 NOR2X1_LOC_560/A INVX1_LOC_230/A 0.01fF
C3011 NAND2X1_LOC_787/B NOR2X1_LOC_48/B 0.02fF
C3012 NOR2X1_LOC_216/Y INVX1_LOC_12/Y 0.25fF
C3013 INVX1_LOC_94/A NAND2X1_LOC_647/B 0.03fF
C3014 NOR2X1_LOC_338/Y INVX1_LOC_128/Y 0.05fF
C3015 NOR2X1_LOC_598/a_36_216# NOR2X1_LOC_334/Y 0.01fF
C3016 NAND2X1_LOC_680/a_36_24# NOR2X1_LOC_152/A 0.00fF
C3017 NOR2X1_LOC_276/Y NOR2X1_LOC_125/Y 0.15fF
C3018 INVX1_LOC_251/Y NAND2X1_LOC_63/Y 0.28fF
C3019 NOR2X1_LOC_186/Y NAND2X1_LOC_475/a_36_24# 0.00fF
C3020 INVX1_LOC_57/Y NOR2X1_LOC_134/a_36_216# 0.02fF
C3021 NOR2X1_LOC_598/B NOR2X1_LOC_307/A 0.03fF
C3022 NOR2X1_LOC_76/A NOR2X1_LOC_177/Y 0.17fF
C3023 NAND2X1_LOC_785/A NOR2X1_LOC_89/A 0.07fF
C3024 INVX1_LOC_2/A NOR2X1_LOC_1/Y -0.00fF
C3025 NAND2X1_LOC_357/B INVX1_LOC_42/A 0.07fF
C3026 NOR2X1_LOC_74/A NOR2X1_LOC_698/Y 0.03fF
C3027 NOR2X1_LOC_826/a_36_216# INVX1_LOC_230/Y 0.00fF
C3028 NOR2X1_LOC_419/Y INVX1_LOC_4/Y 0.10fF
C3029 INVX1_LOC_75/A INVX1_LOC_38/A 0.13fF
C3030 NAND2X1_LOC_363/B NAND2X1_LOC_114/B 0.32fF
C3031 INVX1_LOC_34/A INVX1_LOC_47/Y 0.19fF
C3032 INVX1_LOC_304/Y NOR2X1_LOC_48/B 0.00fF
C3033 INVX1_LOC_77/A INVX1_LOC_94/Y 0.03fF
C3034 INVX1_LOC_72/A NOR2X1_LOC_383/B 0.10fF
C3035 NOR2X1_LOC_632/Y NOR2X1_LOC_631/A 0.00fF
C3036 NOR2X1_LOC_716/B INVX1_LOC_4/Y 0.10fF
C3037 NOR2X1_LOC_474/A INVX1_LOC_253/A 0.28fF
C3038 NOR2X1_LOC_596/a_36_216# INVX1_LOC_271/Y 0.01fF
C3039 NOR2X1_LOC_689/Y INVX1_LOC_136/A 0.06fF
C3040 INVX1_LOC_155/A NOR2X1_LOC_334/Y 0.02fF
C3041 NAND2X1_LOC_656/Y NAND2X1_LOC_475/Y 0.10fF
C3042 NOR2X1_LOC_78/A NOR2X1_LOC_858/B 0.03fF
C3043 NAND2X1_LOC_557/Y INVX1_LOC_18/A 0.04fF
C3044 INVX1_LOC_91/Y INVX1_LOC_118/A 0.02fF
C3045 NOR2X1_LOC_272/Y INVX1_LOC_11/A 0.10fF
C3046 NOR2X1_LOC_860/B NOR2X1_LOC_342/B 0.17fF
C3047 INVX1_LOC_182/A INVX1_LOC_307/A 0.03fF
C3048 INVX1_LOC_25/A NOR2X1_LOC_820/A 0.06fF
C3049 INVX1_LOC_22/A INPUT_7 0.18fF
C3050 NOR2X1_LOC_78/A INVX1_LOC_129/Y 0.01fF
C3051 INVX1_LOC_187/A VDD -0.00fF
C3052 NOR2X1_LOC_456/Y INVX1_LOC_247/Y 0.06fF
C3053 NAND2X1_LOC_342/a_36_24# INVX1_LOC_53/A 0.00fF
C3054 INVX1_LOC_50/A NOR2X1_LOC_303/Y 0.15fF
C3055 NOR2X1_LOC_357/Y NAND2X1_LOC_469/B 0.04fF
C3056 INVX1_LOC_77/A INVX1_LOC_296/A 0.04fF
C3057 NAND2X1_LOC_751/a_36_24# NOR2X1_LOC_68/A 0.00fF
C3058 INVX1_LOC_58/A NOR2X1_LOC_13/Y 0.57fF
C3059 NAND2X1_LOC_357/B INVX1_LOC_78/A 0.08fF
C3060 NOR2X1_LOC_335/B NAND2X1_LOC_93/B 0.23fF
C3061 INVX1_LOC_130/Y NOR2X1_LOC_678/A 0.13fF
C3062 NAND2X1_LOC_466/Y NOR2X1_LOC_449/A 0.04fF
C3063 INVX1_LOC_1/Y NOR2X1_LOC_114/Y 0.00fF
C3064 INVX1_LOC_136/A NAND2X1_LOC_725/A 0.01fF
C3065 NAND2X1_LOC_803/B NOR2X1_LOC_92/Y 0.02fF
C3066 NOR2X1_LOC_220/A INVX1_LOC_32/A 0.05fF
C3067 INVX1_LOC_64/A INVX1_LOC_305/A 0.07fF
C3068 NOR2X1_LOC_639/B NOR2X1_LOC_68/A 0.08fF
C3069 INVX1_LOC_124/A INVX1_LOC_94/Y 0.01fF
C3070 INVX1_LOC_225/A NOR2X1_LOC_278/Y 0.04fF
C3071 INVX1_LOC_14/A NOR2X1_LOC_103/Y 0.18fF
C3072 INVX1_LOC_36/A INVX1_LOC_13/Y 0.15fF
C3073 NOR2X1_LOC_128/B NOR2X1_LOC_847/A 0.08fF
C3074 NOR2X1_LOC_131/A NAND2X1_LOC_454/Y 0.03fF
C3075 NOR2X1_LOC_511/a_36_216# INVX1_LOC_273/A 0.00fF
C3076 NOR2X1_LOC_45/B INVX1_LOC_118/A 0.99fF
C3077 NAND2X1_LOC_725/Y INVX1_LOC_207/A 0.06fF
C3078 NOR2X1_LOC_92/Y NOR2X1_LOC_590/A 0.10fF
C3079 NAND2X1_LOC_214/B NOR2X1_LOC_791/B 0.07fF
C3080 NOR2X1_LOC_15/Y NOR2X1_LOC_596/Y 0.03fF
C3081 INVX1_LOC_286/A INVX1_LOC_92/A 0.07fF
C3082 INVX1_LOC_50/A NOR2X1_LOC_254/Y 0.14fF
C3083 NOR2X1_LOC_756/a_36_216# NAND2X1_LOC_773/B 0.01fF
C3084 NOR2X1_LOC_286/Y INVX1_LOC_134/A 0.04fF
C3085 NOR2X1_LOC_798/A NOR2X1_LOC_751/Y 0.02fF
C3086 INVX1_LOC_14/Y INVX1_LOC_139/Y 0.03fF
C3087 NOR2X1_LOC_577/Y NOR2X1_LOC_493/a_36_216# 0.01fF
C3088 NOR2X1_LOC_196/A INVX1_LOC_5/A 0.01fF
C3089 NOR2X1_LOC_590/A INVX1_LOC_24/Y 0.08fF
C3090 INVX1_LOC_149/A INVX1_LOC_116/Y 0.00fF
C3091 NAND2X1_LOC_799/A INVX1_LOC_161/Y 0.03fF
C3092 INVX1_LOC_89/A INVX1_LOC_106/Y 0.01fF
C3093 INVX1_LOC_44/A NOR2X1_LOC_35/Y 0.06fF
C3094 NOR2X1_LOC_313/a_36_216# INVX1_LOC_84/A 0.02fF
C3095 INVX1_LOC_6/A INVX1_LOC_107/Y 0.06fF
C3096 VDD INVX1_LOC_122/A 0.14fF
C3097 INVX1_LOC_24/Y INVX1_LOC_22/Y 0.31fF
C3098 NAND2X1_LOC_808/A NOR2X1_LOC_48/B 0.14fF
C3099 INVX1_LOC_22/A INVX1_LOC_128/A 0.00fF
C3100 NOR2X1_LOC_78/B INVX1_LOC_16/Y 0.10fF
C3101 NOR2X1_LOC_570/B INVX1_LOC_53/A 0.07fF
C3102 NOR2X1_LOC_476/Y INVX1_LOC_239/A 0.03fF
C3103 NAND2X1_LOC_555/Y NAND2X1_LOC_20/B 0.03fF
C3104 INVX1_LOC_10/Y INVX1_LOC_14/Y 0.23fF
C3105 INVX1_LOC_45/A INVX1_LOC_14/A 0.00fF
C3106 NOR2X1_LOC_709/A INVX1_LOC_57/A 0.03fF
C3107 INVX1_LOC_200/A NOR2X1_LOC_441/Y 0.00fF
C3108 INVX1_LOC_38/A NAND2X1_LOC_453/A 0.07fF
C3109 NOR2X1_LOC_773/Y NOR2X1_LOC_282/Y 0.03fF
C3110 NAND2X1_LOC_863/B NAND2X1_LOC_175/Y 0.03fF
C3111 D_INPUT_3 INVX1_LOC_280/A 0.02fF
C3112 INVX1_LOC_50/A NOR2X1_LOC_353/Y 0.02fF
C3113 INVX1_LOC_36/A INVX1_LOC_88/A 0.13fF
C3114 NAND2X1_LOC_338/B NOR2X1_LOC_383/B 0.02fF
C3115 INVX1_LOC_13/Y NOR2X1_LOC_237/Y 0.01fF
C3116 INVX1_LOC_27/A INVX1_LOC_81/A 0.06fF
C3117 NAND2X1_LOC_468/B NOR2X1_LOC_435/A 0.50fF
C3118 NAND2X1_LOC_323/B NOR2X1_LOC_383/B 0.03fF
C3119 NOR2X1_LOC_78/B NAND2X1_LOC_205/A 0.03fF
C3120 NOR2X1_LOC_272/Y NOR2X1_LOC_433/A 0.12fF
C3121 INVX1_LOC_36/A NAND2X1_LOC_537/a_36_24# 0.01fF
C3122 NOR2X1_LOC_602/A NAND2X1_LOC_337/B 0.01fF
C3123 VDD NOR2X1_LOC_629/Y 0.57fF
C3124 NAND2X1_LOC_348/A NAND2X1_LOC_291/B 0.03fF
C3125 NOR2X1_LOC_75/Y NOR2X1_LOC_723/Y 0.00fF
C3126 INVX1_LOC_223/Y INVX1_LOC_33/A 0.01fF
C3127 NAND2X1_LOC_724/A NAND2X1_LOC_731/Y 0.00fF
C3128 NOR2X1_LOC_772/B NOR2X1_LOC_309/Y 0.03fF
C3129 NAND2X1_LOC_849/A INVX1_LOC_42/A 0.05fF
C3130 NAND2X1_LOC_214/B NOR2X1_LOC_124/B 0.04fF
C3131 INVX1_LOC_11/A NAND2X1_LOC_364/A 0.21fF
C3132 INVX1_LOC_161/Y INVX1_LOC_18/A 0.34fF
C3133 INVX1_LOC_6/A INVX1_LOC_272/A 0.07fF
C3134 INVX1_LOC_35/A NOR2X1_LOC_520/A 0.02fF
C3135 INVX1_LOC_14/A INVX1_LOC_71/A 0.29fF
C3136 INVX1_LOC_13/Y NOR2X1_LOC_309/Y 0.05fF
C3137 NAND2X1_LOC_728/Y INVX1_LOC_161/Y 0.03fF
C3138 NAND2X1_LOC_72/Y INVX1_LOC_54/Y 0.04fF
C3139 INVX1_LOC_280/A INVX1_LOC_230/A 0.18fF
C3140 NOR2X1_LOC_295/Y INVX1_LOC_171/Y 0.08fF
C3141 INVX1_LOC_299/A INVX1_LOC_77/A 0.20fF
C3142 INVX1_LOC_103/A INVX1_LOC_180/A 0.04fF
C3143 INVX1_LOC_40/A NOR2X1_LOC_392/Y 0.07fF
C3144 NOR2X1_LOC_272/Y NOR2X1_LOC_52/B 0.30fF
C3145 NAND2X1_LOC_550/A INVX1_LOC_24/A 0.75fF
C3146 INVX1_LOC_30/A INVX1_LOC_312/Y 0.05fF
C3147 NOR2X1_LOC_92/Y NAND2X1_LOC_354/B 0.01fF
C3148 INPUT_3 INVX1_LOC_62/Y 0.09fF
C3149 NAND2X1_LOC_468/B INVX1_LOC_63/A 0.03fF
C3150 NOR2X1_LOC_314/Y NOR2X1_LOC_697/Y 0.00fF
C3151 INVX1_LOC_62/A NOR2X1_LOC_843/B 0.48fF
C3152 NOR2X1_LOC_406/a_36_216# NOR2X1_LOC_773/Y 0.01fF
C3153 INVX1_LOC_24/A NOR2X1_LOC_160/B 0.16fF
C3154 INVX1_LOC_215/A INVX1_LOC_53/A 0.08fF
C3155 NAND2X1_LOC_756/a_36_24# INVX1_LOC_271/A 0.00fF
C3156 INVX1_LOC_35/A NOR2X1_LOC_748/Y 0.07fF
C3157 INVX1_LOC_269/A NOR2X1_LOC_4/a_36_216# 0.01fF
C3158 INVX1_LOC_89/A INVX1_LOC_275/Y 0.01fF
C3159 NAND2X1_LOC_568/A NAND2X1_LOC_354/B 0.02fF
C3160 INVX1_LOC_75/A NAND2X1_LOC_223/A 0.02fF
C3161 INVX1_LOC_302/Y NOR2X1_LOC_158/Y 0.23fF
C3162 NOR2X1_LOC_405/A NOR2X1_LOC_89/A 0.17fF
C3163 INVX1_LOC_89/A NOR2X1_LOC_748/A 0.08fF
C3164 INVX1_LOC_88/A NOR2X1_LOC_309/Y 0.01fF
C3165 INVX1_LOC_70/Y INVX1_LOC_168/Y 0.00fF
C3166 NOR2X1_LOC_88/Y NOR2X1_LOC_536/A 0.04fF
C3167 NOR2X1_LOC_646/A NAND2X1_LOC_214/B -0.00fF
C3168 INVX1_LOC_313/Y NOR2X1_LOC_383/B 0.39fF
C3169 NOR2X1_LOC_635/A NOR2X1_LOC_636/B 0.06fF
C3170 INVX1_LOC_54/A INVX1_LOC_92/A 0.03fF
C3171 INVX1_LOC_27/A NAND2X1_LOC_672/B 0.04fF
C3172 NOR2X1_LOC_160/B NOR2X1_LOC_557/Y 1.09fF
C3173 NOR2X1_LOC_826/Y INVX1_LOC_135/A 0.03fF
C3174 NAND2X1_LOC_9/Y NOR2X1_LOC_71/Y 0.07fF
C3175 NAND2X1_LOC_563/Y NOR2X1_LOC_82/A 0.68fF
C3176 NOR2X1_LOC_524/Y INVX1_LOC_77/A 0.08fF
C3177 INVX1_LOC_31/Y INVX1_LOC_26/Y 0.21fF
C3178 INVX1_LOC_230/Y NOR2X1_LOC_413/a_36_216# 0.00fF
C3179 NAND2X1_LOC_35/B INVX1_LOC_269/A 0.01fF
C3180 INVX1_LOC_41/A NOR2X1_LOC_590/A 0.13fF
C3181 INVX1_LOC_233/A NOR2X1_LOC_71/Y 0.02fF
C3182 NOR2X1_LOC_536/A INVX1_LOC_84/A 0.10fF
C3183 NOR2X1_LOC_431/Y NOR2X1_LOC_68/A 0.01fF
C3184 INVX1_LOC_41/A INVX1_LOC_22/Y 0.01fF
C3185 NAND2X1_LOC_603/a_36_24# NOR2X1_LOC_605/A 0.00fF
C3186 INVX1_LOC_35/A INVX1_LOC_65/Y 0.25fF
C3187 INVX1_LOC_230/Y NOR2X1_LOC_629/a_36_216# 0.00fF
C3188 INVX1_LOC_11/A NOR2X1_LOC_627/Y 0.02fF
C3189 NOR2X1_LOC_167/Y NOR2X1_LOC_301/A 0.03fF
C3190 NAND2X1_LOC_563/a_36_24# NAND2X1_LOC_141/A -0.01fF
C3191 NOR2X1_LOC_471/Y NAND2X1_LOC_629/Y 0.70fF
C3192 NAND2X1_LOC_364/A NOR2X1_LOC_433/A 1.62fF
C3193 NOR2X1_LOC_548/B INVX1_LOC_26/A 0.01fF
C3194 NAND2X1_LOC_483/Y INVX1_LOC_30/A 0.07fF
C3195 INVX1_LOC_21/A INVX1_LOC_279/A 0.07fF
C3196 INVX1_LOC_11/A NAND2X1_LOC_11/Y 0.09fF
C3197 NOR2X1_LOC_590/A NAND2X1_LOC_477/A 0.03fF
C3198 NOR2X1_LOC_15/Y INVX1_LOC_232/A 0.03fF
C3199 INVX1_LOC_230/Y NOR2X1_LOC_84/Y 0.73fF
C3200 NAND2X1_LOC_553/A NOR2X1_LOC_71/Y 0.03fF
C3201 NOR2X1_LOC_197/A NOR2X1_LOC_209/Y 0.02fF
C3202 NAND2X1_LOC_564/B NOR2X1_LOC_468/Y 0.25fF
C3203 NAND2X1_LOC_364/A NOR2X1_LOC_593/Y 0.05fF
C3204 NOR2X1_LOC_186/Y NOR2X1_LOC_312/Y 0.10fF
C3205 NOR2X1_LOC_814/Y INVX1_LOC_38/Y 0.03fF
C3206 NOR2X1_LOC_653/B NOR2X1_LOC_130/A 0.06fF
C3207 NOR2X1_LOC_160/B INVX1_LOC_143/A 0.13fF
C3208 NAND2X1_LOC_391/Y D_INPUT_0 0.02fF
C3209 NAND2X1_LOC_624/B NOR2X1_LOC_497/Y 0.00fF
C3210 NOR2X1_LOC_239/a_36_216# NOR2X1_LOC_6/B 0.00fF
C3211 NOR2X1_LOC_759/A INVX1_LOC_63/Y 0.01fF
C3212 NAND2X1_LOC_722/A INVX1_LOC_141/Y 0.01fF
C3213 INVX1_LOC_32/A NAND2X1_LOC_414/a_36_24# 0.00fF
C3214 INVX1_LOC_84/A NAND2X1_LOC_93/B 0.22fF
C3215 INVX1_LOC_136/A NAND2X1_LOC_308/Y 0.07fF
C3216 NOR2X1_LOC_664/Y NOR2X1_LOC_791/B 0.01fF
C3217 NOR2X1_LOC_590/A NOR2X1_LOC_405/a_36_216# 0.00fF
C3218 INVX1_LOC_1/A INVX1_LOC_164/A 0.05fF
C3219 INVX1_LOC_12/A NAND2X1_LOC_61/a_36_24# 0.00fF
C3220 INVX1_LOC_36/A INVX1_LOC_168/A 0.44fF
C3221 NOR2X1_LOC_720/B NOR2X1_LOC_68/A 0.05fF
C3222 NOR2X1_LOC_168/B INVX1_LOC_30/A 0.05fF
C3223 INVX1_LOC_177/Y INVX1_LOC_104/A 0.06fF
C3224 INVX1_LOC_224/Y INVX1_LOC_48/A 0.01fF
C3225 INVX1_LOC_45/A INVX1_LOC_111/Y 0.01fF
C3226 NAND2X1_LOC_573/Y NOR2X1_LOC_312/Y 0.10fF
C3227 INVX1_LOC_132/A NAND2X1_LOC_7/Y 0.12fF
C3228 NAND2X1_LOC_364/A NOR2X1_LOC_52/B 0.03fF
C3229 NAND2X1_LOC_642/Y NOR2X1_LOC_278/Y 0.03fF
C3230 NAND2X1_LOC_16/Y INVX1_LOC_266/Y 0.01fF
C3231 INVX1_LOC_84/A NAND2X1_LOC_425/Y 0.01fF
C3232 INVX1_LOC_284/Y NAND2X1_LOC_852/Y 0.05fF
C3233 INVX1_LOC_17/A NOR2X1_LOC_561/Y 0.09fF
C3234 INVX1_LOC_136/A NAND2X1_LOC_660/A 0.10fF
C3235 NAND2X1_LOC_555/Y NOR2X1_LOC_375/Y 0.01fF
C3236 INVX1_LOC_2/A NOR2X1_LOC_52/Y 0.09fF
C3237 NAND2X1_LOC_649/a_36_24# INVX1_LOC_94/Y 0.00fF
C3238 NOR2X1_LOC_172/Y NOR2X1_LOC_577/Y 0.03fF
C3239 NAND2X1_LOC_703/a_36_24# NAND2X1_LOC_703/Y 0.02fF
C3240 INVX1_LOC_14/A NOR2X1_LOC_123/B 0.10fF
C3241 NAND2X1_LOC_574/A NOR2X1_LOC_814/A 0.23fF
C3242 NOR2X1_LOC_860/B NAND2X1_LOC_116/A 0.07fF
C3243 INVX1_LOC_21/A INVX1_LOC_182/Y -0.00fF
C3244 INVX1_LOC_84/A NOR2X1_LOC_649/B 0.09fF
C3245 INVX1_LOC_27/A INVX1_LOC_82/Y 0.03fF
C3246 NAND2X1_LOC_63/Y NOR2X1_LOC_862/B 0.04fF
C3247 INVX1_LOC_84/A INVX1_LOC_3/A 0.10fF
C3248 NOR2X1_LOC_536/A INVX1_LOC_15/A 0.12fF
C3249 NAND2X1_LOC_468/B NOR2X1_LOC_65/Y 0.00fF
C3250 NOR2X1_LOC_392/B NOR2X1_LOC_577/Y 0.02fF
C3251 NAND2X1_LOC_357/B NOR2X1_LOC_152/Y 0.01fF
C3252 INVX1_LOC_71/A NOR2X1_LOC_612/B 0.10fF
C3253 NOR2X1_LOC_710/B INVX1_LOC_89/A 0.04fF
C3254 INPUT_4 INVX1_LOC_296/Y 0.12fF
C3255 NOR2X1_LOC_591/Y NAND2X1_LOC_593/Y 0.07fF
C3256 NAND2X1_LOC_555/Y INVX1_LOC_7/A 0.03fF
C3257 INVX1_LOC_111/Y INVX1_LOC_71/A 0.50fF
C3258 INVX1_LOC_24/Y NOR2X1_LOC_703/A 0.08fF
C3259 NOR2X1_LOC_820/B INVX1_LOC_63/A 0.00fF
C3260 INVX1_LOC_48/Y NOR2X1_LOC_256/Y 0.02fF
C3261 NOR2X1_LOC_806/Y INVX1_LOC_49/A 0.00fF
C3262 NOR2X1_LOC_6/B NAND2X1_LOC_139/A 1.31fF
C3263 NOR2X1_LOC_48/B INVX1_LOC_92/A 5.50fF
C3264 NOR2X1_LOC_850/B INVX1_LOC_307/A 0.07fF
C3265 INVX1_LOC_95/A INVX1_LOC_53/A 0.00fF
C3266 INVX1_LOC_14/A INVX1_LOC_102/Y 0.05fF
C3267 INVX1_LOC_133/Y INVX1_LOC_67/A 0.01fF
C3268 NOR2X1_LOC_98/A NOR2X1_LOC_39/Y 0.01fF
C3269 INVX1_LOC_30/A NAND2X1_LOC_656/Y 0.30fF
C3270 NOR2X1_LOC_244/B NOR2X1_LOC_860/B 0.00fF
C3271 NOR2X1_LOC_457/B NOR2X1_LOC_665/A 0.07fF
C3272 NAND2X1_LOC_93/B INVX1_LOC_15/A 0.03fF
C3273 INVX1_LOC_45/A NOR2X1_LOC_137/A 0.03fF
C3274 NAND2X1_LOC_741/B NOR2X1_LOC_576/B 0.02fF
C3275 NOR2X1_LOC_78/A INVX1_LOC_50/Y 0.43fF
C3276 NOR2X1_LOC_128/B NOR2X1_LOC_554/B 0.03fF
C3277 NOR2X1_LOC_78/B NOR2X1_LOC_570/B 0.16fF
C3278 INVX1_LOC_54/Y NOR2X1_LOC_773/a_36_216# 0.12fF
C3279 NOR2X1_LOC_716/B NAND2X1_LOC_862/A 0.01fF
C3280 INVX1_LOC_39/A NOR2X1_LOC_45/B 0.03fF
C3281 NOR2X1_LOC_593/a_36_216# INVX1_LOC_266/Y 0.01fF
C3282 INVX1_LOC_6/A NOR2X1_LOC_271/B 0.08fF
C3283 NOR2X1_LOC_160/B NOR2X1_LOC_216/Y 0.10fF
C3284 INVX1_LOC_216/Y INPUT_0 0.01fF
C3285 INVX1_LOC_35/A INVX1_LOC_36/Y 0.05fF
C3286 NOR2X1_LOC_363/Y INVX1_LOC_271/A 0.31fF
C3287 INVX1_LOC_30/A NAND2X1_LOC_638/Y 0.06fF
C3288 INVX1_LOC_33/A INVX1_LOC_25/Y 0.26fF
C3289 NOR2X1_LOC_196/A NOR2X1_LOC_332/A 0.02fF
C3290 INVX1_LOC_90/A NOR2X1_LOC_274/B 0.10fF
C3291 NOR2X1_LOC_673/a_36_216# INVX1_LOC_42/A 0.00fF
C3292 INVX1_LOC_17/A NOR2X1_LOC_167/Y 0.03fF
C3293 INVX1_LOC_256/A NOR2X1_LOC_335/B 0.10fF
C3294 INVX1_LOC_41/A NOR2X1_LOC_82/Y 0.03fF
C3295 NAND2X1_LOC_349/B INVX1_LOC_33/A 0.20fF
C3296 NAND2X1_LOC_74/B INVX1_LOC_29/A 0.06fF
C3297 NOR2X1_LOC_328/Y INVX1_LOC_34/A 0.03fF
C3298 NAND2X1_LOC_116/A INVX1_LOC_226/A 0.27fF
C3299 INVX1_LOC_17/A NAND2X1_LOC_251/a_36_24# 0.00fF
C3300 INVX1_LOC_269/A NOR2X1_LOC_337/Y 0.02fF
C3301 NOR2X1_LOC_649/B INVX1_LOC_15/A 0.08fF
C3302 NOR2X1_LOC_107/Y NOR2X1_LOC_548/B 0.05fF
C3303 NAND2X1_LOC_198/B NOR2X1_LOC_76/A 0.05fF
C3304 INVX1_LOC_223/A NOR2X1_LOC_329/B 0.00fF
C3305 NOR2X1_LOC_646/A NOR2X1_LOC_664/Y 0.09fF
C3306 NOR2X1_LOC_759/Y NAND2X1_LOC_140/A 0.00fF
C3307 INVX1_LOC_238/Y NAND2X1_LOC_463/B 3.76fF
C3308 INVX1_LOC_35/A NOR2X1_LOC_706/a_36_216# 0.00fF
C3309 NOR2X1_LOC_392/B INVX1_LOC_22/A 0.01fF
C3310 NOR2X1_LOC_137/A INVX1_LOC_71/A 0.27fF
C3311 INVX1_LOC_150/Y INVX1_LOC_6/A 0.07fF
C3312 NAND2X1_LOC_214/B INVX1_LOC_2/Y 0.04fF
C3313 INVX1_LOC_202/A NAND2X1_LOC_140/A 0.02fF
C3314 NOR2X1_LOC_226/A NOR2X1_LOC_401/Y 0.02fF
C3315 NOR2X1_LOC_209/Y INVX1_LOC_83/Y 0.04fF
C3316 INVX1_LOC_136/A NAND2X1_LOC_560/A 0.06fF
C3317 INVX1_LOC_278/A NOR2X1_LOC_536/A 0.07fF
C3318 INVX1_LOC_72/A NOR2X1_LOC_163/Y 0.00fF
C3319 NOR2X1_LOC_186/Y NAND2X1_LOC_287/B 0.07fF
C3320 NOR2X1_LOC_489/A INVX1_LOC_57/A 0.01fF
C3321 INVX1_LOC_292/A NOR2X1_LOC_551/Y 0.02fF
C3322 NOR2X1_LOC_548/Y NOR2X1_LOC_337/a_36_216# 0.00fF
C3323 NOR2X1_LOC_191/A NAND2X1_LOC_850/Y 0.11fF
C3324 NOR2X1_LOC_826/Y INVX1_LOC_280/A 0.01fF
C3325 NOR2X1_LOC_607/a_36_216# INVX1_LOC_313/Y 0.00fF
C3326 NOR2X1_LOC_250/Y INVX1_LOC_91/A 0.04fF
C3327 NOR2X1_LOC_295/a_36_216# INVX1_LOC_10/A 0.00fF
C3328 NOR2X1_LOC_267/a_36_216# INVX1_LOC_95/A 0.00fF
C3329 NOR2X1_LOC_52/B NOR2X1_LOC_86/A 0.72fF
C3330 INVX1_LOC_27/A INVX1_LOC_2/Y 0.03fF
C3331 INVX1_LOC_34/A INVX1_LOC_219/A 0.03fF
C3332 INVX1_LOC_200/Y NOR2X1_LOC_487/Y 0.01fF
C3333 NOR2X1_LOC_93/Y VDD 0.00fF
C3334 NOR2X1_LOC_690/A INVX1_LOC_135/A 0.02fF
C3335 NAND2X1_LOC_444/B NOR2X1_LOC_662/A 0.10fF
C3336 INVX1_LOC_90/A NOR2X1_LOC_577/Y 0.07fF
C3337 NOR2X1_LOC_516/B INVX1_LOC_143/A 0.10fF
C3338 INVX1_LOC_269/A NAND2X1_LOC_659/B 0.01fF
C3339 INVX1_LOC_21/A NAND2X1_LOC_298/a_36_24# 0.01fF
C3340 INVX1_LOC_53/A INVX1_LOC_54/A 1.40fF
C3341 INVX1_LOC_52/Y NOR2X1_LOC_357/Y -0.00fF
C3342 NOR2X1_LOC_413/Y INVX1_LOC_135/A 0.09fF
C3343 NOR2X1_LOC_346/A NOR2X1_LOC_861/Y 0.05fF
C3344 INVX1_LOC_11/A NAND2X1_LOC_422/a_36_24# 0.01fF
C3345 NAND2X1_LOC_37/a_36_24# INVX1_LOC_315/Y 0.00fF
C3346 INVX1_LOC_24/A NOR2X1_LOC_706/A 0.07fF
C3347 INVX1_LOC_225/A NOR2X1_LOC_312/Y 0.01fF
C3348 NOR2X1_LOC_824/A INVX1_LOC_37/Y 0.02fF
C3349 INVX1_LOC_30/A INVX1_LOC_78/Y 0.03fF
C3350 INVX1_LOC_215/A NOR2X1_LOC_78/B 1.74fF
C3351 INVX1_LOC_119/Y NOR2X1_LOC_693/Y 0.01fF
C3352 NAND2X1_LOC_456/Y INVX1_LOC_23/Y 0.01fF
C3353 INVX1_LOC_55/Y INVX1_LOC_63/Y 0.00fF
C3354 INVX1_LOC_265/A INPUT_1 0.03fF
C3355 NOR2X1_LOC_487/a_36_216# INVX1_LOC_6/A 0.00fF
C3356 NOR2X1_LOC_604/Y INVX1_LOC_179/A 0.01fF
C3357 INVX1_LOC_17/A INVX1_LOC_76/A 0.30fF
C3358 INVX1_LOC_124/Y INVX1_LOC_91/A 0.51fF
C3359 INVX1_LOC_269/A VDD 3.85fF
C3360 NOR2X1_LOC_123/B NOR2X1_LOC_612/B 0.03fF
C3361 NOR2X1_LOC_160/B NOR2X1_LOC_209/A 0.06fF
C3362 NOR2X1_LOC_589/A NAND2X1_LOC_841/A 0.04fF
C3363 NOR2X1_LOC_232/Y VDD 0.02fF
C3364 INVX1_LOC_90/A NOR2X1_LOC_348/B 0.46fF
C3365 INVX1_LOC_41/A NOR2X1_LOC_703/A 0.12fF
C3366 NAND2X1_LOC_341/A INVX1_LOC_290/A 0.01fF
C3367 INVX1_LOC_11/A NOR2X1_LOC_857/A 0.07fF
C3368 INVX1_LOC_58/A NOR2X1_LOC_697/Y 0.01fF
C3369 INVX1_LOC_267/A INVX1_LOC_89/A 0.02fF
C3370 NOR2X1_LOC_174/B NOR2X1_LOC_175/A 0.02fF
C3371 NOR2X1_LOC_471/Y INVX1_LOC_76/A 0.02fF
C3372 INVX1_LOC_268/A NOR2X1_LOC_589/A 0.03fF
C3373 NOR2X1_LOC_223/B NAND2X1_LOC_93/B 0.05fF
C3374 INVX1_LOC_57/A INVX1_LOC_294/A 0.03fF
C3375 INVX1_LOC_33/A INVX1_LOC_75/A 0.27fF
C3376 NOR2X1_LOC_284/a_36_216# INVX1_LOC_83/A 0.00fF
C3377 NOR2X1_LOC_662/A NAND2X1_LOC_464/B 0.10fF
C3378 NAND2X1_LOC_149/Y INVX1_LOC_193/A 0.01fF
C3379 NAND2X1_LOC_223/A GATE_222 0.02fF
C3380 INVX1_LOC_84/A NOR2X1_LOC_476/B 0.00fF
C3381 INVX1_LOC_61/A NOR2X1_LOC_45/B 0.07fF
C3382 NOR2X1_LOC_382/a_36_216# NOR2X1_LOC_332/A 0.00fF
C3383 NOR2X1_LOC_401/Y INPUT_1 0.05fF
C3384 NOR2X1_LOC_223/B NAND2X1_LOC_425/Y 0.03fF
C3385 NAND2X1_LOC_214/B NOR2X1_LOC_608/Y 0.01fF
C3386 INVX1_LOC_135/Y NOR2X1_LOC_399/A 0.05fF
C3387 NOR2X1_LOC_781/A NOR2X1_LOC_781/B 0.03fF
C3388 INVX1_LOC_90/A NOR2X1_LOC_175/B 0.08fF
C3389 NOR2X1_LOC_190/a_36_216# NAND2X1_LOC_842/B 0.00fF
C3390 INVX1_LOC_299/A INVX1_LOC_9/A 0.10fF
C3391 NOR2X1_LOC_445/Y INVX1_LOC_69/Y 0.02fF
C3392 NAND2X1_LOC_470/B INVX1_LOC_15/A 0.00fF
C3393 NOR2X1_LOC_538/B INVX1_LOC_9/A 0.34fF
C3394 NAND2X1_LOC_740/Y INVX1_LOC_297/A 0.02fF
C3395 INVX1_LOC_90/A INVX1_LOC_22/A 0.26fF
C3396 NOR2X1_LOC_772/B INVX1_LOC_63/A 0.02fF
C3397 NOR2X1_LOC_19/B NAND2X1_LOC_672/B 0.17fF
C3398 NOR2X1_LOC_389/B INVX1_LOC_22/A 0.39fF
C3399 NOR2X1_LOC_815/Y NOR2X1_LOC_45/B 0.08fF
C3400 INVX1_LOC_226/Y NOR2X1_LOC_756/Y 0.01fF
C3401 INVX1_LOC_149/A NOR2X1_LOC_188/A 0.10fF
C3402 NOR2X1_LOC_433/A NOR2X1_LOC_405/A 0.06fF
C3403 NOR2X1_LOC_187/Y INVX1_LOC_307/A 0.01fF
C3404 NAND2X1_LOC_348/A NOR2X1_LOC_346/B 0.00fF
C3405 INVX1_LOC_104/A INVX1_LOC_206/Y 0.02fF
C3406 NOR2X1_LOC_646/A NOR2X1_LOC_19/B 0.39fF
C3407 NOR2X1_LOC_432/Y NAND2X1_LOC_832/Y 0.05fF
C3408 INVX1_LOC_149/A NOR2X1_LOC_548/B 0.34fF
C3409 NOR2X1_LOC_660/Y INVX1_LOC_29/A 0.07fF
C3410 NOR2X1_LOC_464/a_36_216# INVX1_LOC_96/A 0.01fF
C3411 INVX1_LOC_208/A NOR2X1_LOC_216/Y 0.08fF
C3412 INVX1_LOC_13/Y INVX1_LOC_63/A 0.08fF
C3413 NOR2X1_LOC_593/Y NOR2X1_LOC_405/A 0.98fF
C3414 INVX1_LOC_53/A NAND2X1_LOC_807/B 0.04fF
C3415 NOR2X1_LOC_667/A NAND2X1_LOC_858/B 0.03fF
C3416 NOR2X1_LOC_793/A NAND2X1_LOC_237/a_36_24# 0.00fF
C3417 NOR2X1_LOC_824/A NOR2X1_LOC_485/Y 0.04fF
C3418 INVX1_LOC_73/A INVX1_LOC_53/Y 0.03fF
C3419 INVX1_LOC_248/A NAND2X1_LOC_858/B 0.01fF
C3420 NOR2X1_LOC_6/B NOR2X1_LOC_78/A 0.01fF
C3421 NAND2X1_LOC_354/B NAND2X1_LOC_648/a_36_24# 0.00fF
C3422 NOR2X1_LOC_496/Y NAND2X1_LOC_489/Y 0.00fF
C3423 NOR2X1_LOC_717/Y NOR2X1_LOC_331/B 0.00fF
C3424 INVX1_LOC_150/Y INVX1_LOC_131/Y 0.03fF
C3425 INVX1_LOC_53/A NOR2X1_LOC_48/B 0.10fF
C3426 INVX1_LOC_35/A INVX1_LOC_102/A 1.81fF
C3427 NOR2X1_LOC_500/B NOR2X1_LOC_865/A 0.15fF
C3428 NOR2X1_LOC_78/B INVX1_LOC_286/A 0.07fF
C3429 INVX1_LOC_47/A INVX1_LOC_171/A 0.16fF
C3430 NAND2X1_LOC_350/A INVX1_LOC_92/A 0.17fF
C3431 INVX1_LOC_72/A NAND2X1_LOC_476/a_36_24# 0.00fF
C3432 NOR2X1_LOC_52/B NOR2X1_LOC_405/A 0.10fF
C3433 NOR2X1_LOC_76/A NOR2X1_LOC_76/a_36_216# 0.01fF
C3434 INVX1_LOC_240/Y INVX1_LOC_242/A 0.10fF
C3435 NOR2X1_LOC_355/A NAND2X1_LOC_123/Y 0.04fF
C3436 D_INPUT_6 NOR2X1_LOC_11/Y 0.19fF
C3437 NOR2X1_LOC_553/B NOR2X1_LOC_74/A 0.00fF
C3438 NOR2X1_LOC_160/B NOR2X1_LOC_197/B 0.02fF
C3439 NOR2X1_LOC_334/Y INVX1_LOC_57/A 0.00fF
C3440 INVX1_LOC_41/A NAND2X1_LOC_650/B 0.03fF
C3441 NOR2X1_LOC_620/Y INVX1_LOC_37/A 0.03fF
C3442 NOR2X1_LOC_321/Y INVX1_LOC_19/A 0.06fF
C3443 NOR2X1_LOC_357/Y INVX1_LOC_63/Y 0.13fF
C3444 INVX1_LOC_88/A INVX1_LOC_63/A 0.03fF
C3445 NOR2X1_LOC_291/Y INVX1_LOC_42/A 0.03fF
C3446 INVX1_LOC_53/A NAND2X1_LOC_3/B 0.41fF
C3447 NOR2X1_LOC_473/B INVX1_LOC_28/A -0.09fF
C3448 INVX1_LOC_132/A INVX1_LOC_129/Y 0.00fF
C3449 INVX1_LOC_77/A NAND2X1_LOC_96/A 0.07fF
C3450 INVX1_LOC_36/A NOR2X1_LOC_99/Y 0.06fF
C3451 NOR2X1_LOC_859/A NOR2X1_LOC_61/Y 0.01fF
C3452 INVX1_LOC_256/A INVX1_LOC_84/A 0.01fF
C3453 NOR2X1_LOC_664/Y INVX1_LOC_2/Y 0.59fF
C3454 D_INPUT_0 INVX1_LOC_79/A 0.02fF
C3455 INVX1_LOC_50/A NOR2X1_LOC_829/A 0.00fF
C3456 INVX1_LOC_225/A NAND2X1_LOC_287/B 0.09fF
C3457 INVX1_LOC_219/A INPUT_0 0.02fF
C3458 NAND2X1_LOC_466/A NAND2X1_LOC_453/A -0.01fF
C3459 NAND2X1_LOC_400/a_36_24# INVX1_LOC_23/A 0.00fF
C3460 NOR2X1_LOC_384/Y NOR2X1_LOC_235/Y 0.03fF
C3461 NAND2X1_LOC_477/A NAND2X1_LOC_650/B 0.80fF
C3462 INVX1_LOC_286/A NAND2X1_LOC_392/Y 0.03fF
C3463 NAND2X1_LOC_541/Y NOR2X1_LOC_124/A 0.22fF
C3464 NAND2X1_LOC_579/A INVX1_LOC_12/A 0.26fF
C3465 NOR2X1_LOC_577/Y INVX1_LOC_38/A 0.17fF
C3466 NOR2X1_LOC_690/A NOR2X1_LOC_813/Y 0.02fF
C3467 NAND2X1_LOC_717/Y NAND2X1_LOC_836/Y 0.01fF
C3468 INVX1_LOC_31/A NOR2X1_LOC_673/A 0.07fF
C3469 NOR2X1_LOC_45/B NAND2X1_LOC_735/B 0.01fF
C3470 INVX1_LOC_136/A NOR2X1_LOC_58/Y 0.03fF
C3471 NAND2X1_LOC_793/Y INVX1_LOC_19/A 0.03fF
C3472 NAND2X1_LOC_392/A NAND2X1_LOC_642/Y 0.01fF
C3473 NAND2X1_LOC_660/Y INVX1_LOC_91/A 0.92fF
C3474 INVX1_LOC_30/Y NOR2X1_LOC_78/A 0.12fF
C3475 NOR2X1_LOC_791/B NOR2X1_LOC_216/B 0.03fF
C3476 NOR2X1_LOC_78/B NAND2X1_LOC_454/a_36_24# 0.00fF
C3477 NOR2X1_LOC_15/Y NOR2X1_LOC_46/a_36_216# 0.00fF
C3478 INVX1_LOC_224/Y NOR2X1_LOC_383/B 0.02fF
C3479 INVX1_LOC_82/Y NOR2X1_LOC_19/B 0.10fF
C3480 NOR2X1_LOC_322/Y INVX1_LOC_28/A 0.89fF
C3481 NOR2X1_LOC_606/Y INVX1_LOC_84/A 0.01fF
C3482 NOR2X1_LOC_816/A INVX1_LOC_264/A 0.04fF
C3483 NOR2X1_LOC_690/A INVX1_LOC_280/A 0.00fF
C3484 NOR2X1_LOC_45/B INPUT_5 0.03fF
C3485 INVX1_LOC_18/A NOR2X1_LOC_841/A 0.12fF
C3486 NAND2X1_LOC_727/Y INVX1_LOC_11/Y 0.01fF
C3487 NOR2X1_LOC_616/Y VDD 0.12fF
C3488 INVX1_LOC_5/A NOR2X1_LOC_158/Y 0.07fF
C3489 NAND2X1_LOC_725/A NOR2X1_LOC_395/Y 0.12fF
C3490 NOR2X1_LOC_413/Y INVX1_LOC_280/A 0.01fF
C3491 NAND2X1_LOC_9/Y NOR2X1_LOC_39/Y 0.01fF
C3492 NAND2X1_LOC_798/A NAND2X1_LOC_453/A 0.04fF
C3493 NOR2X1_LOC_589/A INVX1_LOC_95/Y 0.03fF
C3494 NAND2X1_LOC_192/B INVX1_LOC_290/Y 0.03fF
C3495 INVX1_LOC_95/A NAND2X1_LOC_392/Y 0.01fF
C3496 D_INPUT_0 INVX1_LOC_91/A 0.23fF
C3497 NAND2X1_LOC_563/A VDD 0.38fF
C3498 NAND2X1_LOC_802/A NAND2X1_LOC_798/B 0.03fF
C3499 INVX1_LOC_73/A NAND2X1_LOC_124/a_36_24# 0.02fF
C3500 NAND2X1_LOC_500/Y NAND2X1_LOC_500/B 0.15fF
C3501 NAND2X1_LOC_9/Y NAND2X1_LOC_205/A 0.03fF
C3502 INVX1_LOC_62/A NAND2X1_LOC_86/Y 0.00fF
C3503 INVX1_LOC_73/A NOR2X1_LOC_113/B 0.03fF
C3504 NOR2X1_LOC_382/Y NAND2X1_LOC_82/Y 0.01fF
C3505 NOR2X1_LOC_781/A NOR2X1_LOC_585/Y 0.03fF
C3506 NOR2X1_LOC_312/Y NAND2X1_LOC_642/Y 0.00fF
C3507 NOR2X1_LOC_551/B INVX1_LOC_307/A 0.01fF
C3508 NOR2X1_LOC_142/Y INVX1_LOC_92/A 1.50fF
C3509 INVX1_LOC_36/A INVX1_LOC_272/A 0.49fF
C3510 INVX1_LOC_215/A INVX1_LOC_46/A 0.16fF
C3511 INVX1_LOC_94/A NOR2X1_LOC_814/A 0.07fF
C3512 INVX1_LOC_171/A INVX1_LOC_95/Y 0.05fF
C3513 INVX1_LOC_256/A INVX1_LOC_15/A 0.24fF
C3514 NOR2X1_LOC_216/a_36_216# INVX1_LOC_91/A 0.01fF
C3515 INVX1_LOC_136/A INVX1_LOC_29/A 0.20fF
C3516 NOR2X1_LOC_124/B NOR2X1_LOC_216/B 0.04fF
C3517 INVX1_LOC_69/Y NOR2X1_LOC_335/B 0.13fF
C3518 INVX1_LOC_266/Y NOR2X1_LOC_433/Y 0.02fF
C3519 NOR2X1_LOC_76/A NAND2X1_LOC_465/A 0.02fF
C3520 NOR2X1_LOC_561/A INVX1_LOC_22/A 0.03fF
C3521 INVX1_LOC_18/A INPUT_7 0.02fF
C3522 INVX1_LOC_223/Y NOR2X1_LOC_748/A 0.03fF
C3523 INVX1_LOC_280/Y NOR2X1_LOC_629/Y 0.02fF
C3524 NOR2X1_LOC_78/B INVX1_LOC_54/A 2.10fF
C3525 INVX1_LOC_303/A INVX1_LOC_63/A 0.15fF
C3526 NOR2X1_LOC_373/Y INVX1_LOC_46/A 0.11fF
C3527 INVX1_LOC_76/Y NAND2X1_LOC_425/Y 0.04fF
C3528 INVX1_LOC_22/A INVX1_LOC_38/A 0.99fF
C3529 NAND2X1_LOC_451/Y NAND2X1_LOC_638/a_36_24# 0.00fF
C3530 NAND2X1_LOC_795/Y NAND2X1_LOC_804/Y 0.02fF
C3531 INVX1_LOC_188/A INVX1_LOC_4/A 0.01fF
C3532 NOR2X1_LOC_95/a_36_216# NOR2X1_LOC_11/Y 0.02fF
C3533 INVX1_LOC_24/A NAND2X1_LOC_207/B 0.03fF
C3534 VDD NOR2X1_LOC_814/Y 0.15fF
C3535 NOR2X1_LOC_655/B INVX1_LOC_92/A 0.38fF
C3536 NOR2X1_LOC_214/B VDD 0.19fF
C3537 NAND2X1_LOC_342/Y NOR2X1_LOC_155/A 0.03fF
C3538 NOR2X1_LOC_105/Y NAND2X1_LOC_473/A 0.02fF
C3539 INVX1_LOC_88/A NOR2X1_LOC_65/Y 0.02fF
C3540 NOR2X1_LOC_778/B NOR2X1_LOC_600/a_36_216# 0.00fF
C3541 INVX1_LOC_75/A NOR2X1_LOC_486/Y 0.03fF
C3542 INVX1_LOC_8/A INVX1_LOC_293/Y 0.14fF
C3543 NOR2X1_LOC_112/B NAND2X1_LOC_109/a_36_24# 0.00fF
C3544 NOR2X1_LOC_147/B INVX1_LOC_186/Y 0.08fF
C3545 INVX1_LOC_228/A NOR2X1_LOC_847/B 0.01fF
C3546 NOR2X1_LOC_51/A INVX1_LOC_22/A 4.91fF
C3547 INVX1_LOC_50/A NAND2X1_LOC_537/Y 0.00fF
C3548 NAND2X1_LOC_569/A NAND2X1_LOC_773/B 0.10fF
C3549 NOR2X1_LOC_19/B INVX1_LOC_2/Y 0.03fF
C3550 NOR2X1_LOC_312/a_36_216# INVX1_LOC_285/A 0.00fF
C3551 NAND2X1_LOC_392/Y INVX1_LOC_54/A 0.01fF
C3552 NOR2X1_LOC_433/A INVX1_LOC_109/Y 0.98fF
C3553 INVX1_LOC_30/A INVX1_LOC_128/Y 0.01fF
C3554 NAND2X1_LOC_198/B NAND2X1_LOC_404/a_36_24# 0.00fF
C3555 NOR2X1_LOC_103/Y NOR2X1_LOC_383/B 0.01fF
C3556 INVX1_LOC_308/Y INVX1_LOC_57/A 0.01fF
C3557 INVX1_LOC_168/A INVX1_LOC_63/A 0.04fF
C3558 NOR2X1_LOC_216/Y NAND2X1_LOC_211/Y 1.68fF
C3559 NOR2X1_LOC_541/Y NOR2X1_LOC_383/B 0.00fF
C3560 INVX1_LOC_33/A NAND2X1_LOC_291/B 0.07fF
C3561 INVX1_LOC_8/A NAND2X1_LOC_74/B 1.16fF
C3562 NOR2X1_LOC_781/Y INVX1_LOC_15/A 0.03fF
C3563 INVX1_LOC_150/Y INVX1_LOC_270/A 0.15fF
C3564 NAND2X1_LOC_208/B INVX1_LOC_23/Y 0.11fF
C3565 INVX1_LOC_83/A INVX1_LOC_54/A 0.55fF
C3566 NOR2X1_LOC_121/A INVX1_LOC_123/Y 0.34fF
C3567 NAND2X1_LOC_778/Y NAND2X1_LOC_796/B 0.03fF
C3568 INVX1_LOC_35/A NAND2X1_LOC_774/a_36_24# 0.00fF
C3569 NOR2X1_LOC_589/Y INVX1_LOC_37/A 0.02fF
C3570 INVX1_LOC_25/A INVX1_LOC_230/Y 1.15fF
C3571 INVX1_LOC_136/A NOR2X1_LOC_281/Y 0.02fF
C3572 NOR2X1_LOC_52/B INVX1_LOC_109/Y 0.53fF
C3573 NAND2X1_LOC_350/A INVX1_LOC_53/A 0.64fF
C3574 NAND2X1_LOC_842/B NAND2X1_LOC_698/a_36_24# 0.01fF
C3575 INVX1_LOC_256/A INVX1_LOC_278/A 0.02fF
C3576 INVX1_LOC_30/A NOR2X1_LOC_727/B 0.03fF
C3577 NOR2X1_LOC_5/a_36_216# NOR2X1_LOC_655/Y 0.00fF
C3578 INVX1_LOC_311/A NAND2X1_LOC_298/a_36_24# 0.00fF
C3579 INVX1_LOC_45/A NOR2X1_LOC_383/B 0.07fF
C3580 INVX1_LOC_13/A INVX1_LOC_27/Y 0.01fF
C3581 INVX1_LOC_286/A INVX1_LOC_46/A 0.14fF
C3582 NOR2X1_LOC_298/Y NAND2X1_LOC_770/Y 0.04fF
C3583 NAND2X1_LOC_724/Y NOR2X1_LOC_599/A 0.05fF
C3584 INVX1_LOC_63/Y INVX1_LOC_32/A 0.02fF
C3585 NOR2X1_LOC_741/A VDD 0.24fF
C3586 NOR2X1_LOC_440/Y INVX1_LOC_84/A 0.98fF
C3587 INVX1_LOC_58/A NOR2X1_LOC_426/Y 0.20fF
C3588 NOR2X1_LOC_145/a_36_216# INVX1_LOC_91/A 0.00fF
C3589 INVX1_LOC_21/A NOR2X1_LOC_468/Y 0.07fF
C3590 NOR2X1_LOC_441/Y INVX1_LOC_53/A 0.05fF
C3591 NAND2X1_LOC_35/Y NOR2X1_LOC_615/Y 0.03fF
C3592 INVX1_LOC_313/Y INVX1_LOC_179/A 0.00fF
C3593 INVX1_LOC_120/Y NAND2X1_LOC_291/B 0.01fF
C3594 NOR2X1_LOC_195/A INVX1_LOC_5/A 0.01fF
C3595 INVX1_LOC_21/A NAND2X1_LOC_190/Y 0.05fF
C3596 NOR2X1_LOC_266/B INVX1_LOC_91/A 0.01fF
C3597 NOR2X1_LOC_45/B D_INPUT_3 0.03fF
C3598 INVX1_LOC_64/A INVX1_LOC_188/A 0.09fF
C3599 NAND2X1_LOC_738/B NAND2X1_LOC_856/A 0.00fF
C3600 INVX1_LOC_95/Y INVX1_LOC_20/A 0.10fF
C3601 INVX1_LOC_30/A NOR2X1_LOC_717/A 0.12fF
C3602 NOR2X1_LOC_528/Y INVX1_LOC_37/Y 0.06fF
C3603 NAND2X1_LOC_287/B NAND2X1_LOC_642/Y 0.07fF
C3604 INVX1_LOC_57/Y NAND2X1_LOC_793/B 0.10fF
C3605 NOR2X1_LOC_19/B NOR2X1_LOC_608/Y 0.01fF
C3606 INVX1_LOC_123/A NOR2X1_LOC_536/A 0.01fF
C3607 NOR2X1_LOC_103/Y NAND2X1_LOC_75/a_36_24# 0.01fF
C3608 D_INPUT_0 INVX1_LOC_203/A 0.03fF
C3609 NOR2X1_LOC_175/A NOR2X1_LOC_623/B 0.10fF
C3610 INVX1_LOC_142/A NOR2X1_LOC_678/A 0.02fF
C3611 INVX1_LOC_71/A NOR2X1_LOC_383/B 0.11fF
C3612 INVX1_LOC_36/A NAND2X1_LOC_708/Y 0.01fF
C3613 INVX1_LOC_211/Y INVX1_LOC_178/A 0.41fF
C3614 NAND2X1_LOC_555/Y NOR2X1_LOC_34/B 0.05fF
C3615 INVX1_LOC_201/Y NOR2X1_LOC_415/Y 0.04fF
C3616 INVX1_LOC_217/A NAND2X1_LOC_827/a_36_24# 0.05fF
C3617 INVX1_LOC_129/Y NAND2X1_LOC_642/Y 0.03fF
C3618 NAND2X1_LOC_391/Y NOR2X1_LOC_134/Y 0.03fF
C3619 NAND2X1_LOC_848/A INVX1_LOC_91/A 0.10fF
C3620 INPUT_5 NOR2X1_LOC_1/Y 0.43fF
C3621 NOR2X1_LOC_321/Y INVX1_LOC_161/Y 0.03fF
C3622 NOR2X1_LOC_768/a_36_216# NOR2X1_LOC_814/A 0.00fF
C3623 NOR2X1_LOC_326/Y NOR2X1_LOC_856/B 0.17fF
C3624 INVX1_LOC_21/A NOR2X1_LOC_389/A 0.03fF
C3625 INVX1_LOC_200/A NAND2X1_LOC_579/A 0.10fF
C3626 NOR2X1_LOC_305/Y INVX1_LOC_20/A 0.21fF
C3627 INVX1_LOC_34/A INVX1_LOC_23/Y 0.08fF
C3628 NOR2X1_LOC_589/A NAND2X1_LOC_806/a_36_24# 0.01fF
C3629 INVX1_LOC_255/Y NOR2X1_LOC_643/a_36_216# 0.01fF
C3630 INVX1_LOC_90/A INVX1_LOC_186/Y 0.07fF
C3631 INVX1_LOC_136/A NAND2X1_LOC_557/a_36_24# 0.01fF
C3632 NAND2X1_LOC_555/Y INVX1_LOC_163/A 0.07fF
C3633 INVX1_LOC_228/A NOR2X1_LOC_660/Y 0.10fF
C3634 NAND2X1_LOC_338/B INVX1_LOC_165/A 0.03fF
C3635 NAND2X1_LOC_212/Y INVX1_LOC_281/A 0.19fF
C3636 NAND2X1_LOC_326/A INVX1_LOC_141/A 0.02fF
C3637 INVX1_LOC_230/Y INVX1_LOC_1/A 0.10fF
C3638 INVX1_LOC_5/A NOR2X1_LOC_759/A 0.07fF
C3639 NOR2X1_LOC_68/A NOR2X1_LOC_406/A 0.00fF
C3640 VDD INVX1_LOC_12/Y 2.86fF
C3641 INVX1_LOC_230/Y NAND2X1_LOC_131/a_36_24# 0.01fF
C3642 NOR2X1_LOC_835/A NOR2X1_LOC_839/B 0.03fF
C3643 INVX1_LOC_83/A NOR2X1_LOC_48/B 0.10fF
C3644 NAND2X1_LOC_725/B NAND2X1_LOC_500/Y 0.01fF
C3645 VDD NOR2X1_LOC_492/Y 0.21fF
C3646 INVX1_LOC_37/A INVX1_LOC_117/A 1.33fF
C3647 INVX1_LOC_140/A INVX1_LOC_264/A 0.37fF
C3648 NOR2X1_LOC_142/Y INVX1_LOC_53/A 0.10fF
C3649 INVX1_LOC_91/A INVX1_LOC_46/Y 0.08fF
C3650 INVX1_LOC_21/A INVX1_LOC_62/Y 0.19fF
C3651 INVX1_LOC_157/A INVX1_LOC_15/A 0.02fF
C3652 NOR2X1_LOC_164/Y INVX1_LOC_54/A 0.04fF
C3653 NOR2X1_LOC_361/Y INVX1_LOC_271/A 0.01fF
C3654 INVX1_LOC_69/Y INVX1_LOC_84/A 0.45fF
C3655 INVX1_LOC_37/A NOR2X1_LOC_808/B 0.13fF
C3656 INVX1_LOC_276/A NOR2X1_LOC_677/Y 0.00fF
C3657 NAND2X1_LOC_579/A INVX1_LOC_217/A 0.10fF
C3658 INVX1_LOC_206/A INVX1_LOC_29/Y 0.07fF
C3659 INVX1_LOC_243/A INVX1_LOC_296/A 0.03fF
C3660 NOR2X1_LOC_602/B INVX1_LOC_46/A 0.00fF
C3661 INVX1_LOC_35/A INVX1_LOC_149/Y 0.01fF
C3662 INVX1_LOC_35/A INVX1_LOC_162/Y 0.05fF
C3663 NOR2X1_LOC_272/Y INVX1_LOC_314/Y 0.03fF
C3664 INVX1_LOC_132/A INVX1_LOC_50/Y 0.10fF
C3665 INVX1_LOC_123/A INVX1_LOC_3/A 0.14fF
C3666 INVX1_LOC_222/Y INVX1_LOC_77/A 0.95fF
C3667 NOR2X1_LOC_561/Y INVX1_LOC_94/Y 0.01fF
C3668 INVX1_LOC_83/A NAND2X1_LOC_3/B 0.89fF
C3669 INVX1_LOC_111/Y NOR2X1_LOC_493/A 0.04fF
C3670 NOR2X1_LOC_78/B NAND2X1_LOC_215/A 0.13fF
C3671 NOR2X1_LOC_393/a_36_216# NAND2X1_LOC_254/Y 0.01fF
C3672 INVX1_LOC_46/A INVX1_LOC_54/A 1.75fF
C3673 INVX1_LOC_36/A INVX1_LOC_150/Y 0.59fF
C3674 INVX1_LOC_196/Y NOR2X1_LOC_801/B 0.09fF
C3675 NOR2X1_LOC_9/Y INVX1_LOC_125/A -0.00fF
C3676 NAND2X1_LOC_96/A INVX1_LOC_9/A 0.07fF
C3677 NOR2X1_LOC_335/B NOR2X1_LOC_89/A 0.07fF
C3678 NAND2X1_LOC_741/B INVX1_LOC_161/A 0.01fF
C3679 NAND2X1_LOC_787/A INVX1_LOC_256/Y 0.00fF
C3680 INVX1_LOC_58/A INVX1_LOC_289/A 0.06fF
C3681 NAND2X1_LOC_848/A NAND2X1_LOC_783/a_36_24# 0.06fF
C3682 INVX1_LOC_11/Y INVX1_LOC_5/Y 0.03fF
C3683 NAND2X1_LOC_579/A NAND2X1_LOC_787/B 0.01fF
C3684 NOR2X1_LOC_607/A INVX1_LOC_161/Y 0.04fF
C3685 NOR2X1_LOC_709/A INVX1_LOC_306/Y 0.06fF
C3686 NOR2X1_LOC_346/Y NAND2X1_LOC_206/Y 0.04fF
C3687 INVX1_LOC_17/A NOR2X1_LOC_274/Y 0.02fF
C3688 NOR2X1_LOC_658/Y INVX1_LOC_30/A 0.21fF
C3689 NAND2X1_LOC_67/a_36_24# INVX1_LOC_153/Y 0.06fF
C3690 INVX1_LOC_58/A NOR2X1_LOC_605/a_36_216# 0.00fF
C3691 INVX1_LOC_254/Y INVX1_LOC_224/A 0.00fF
C3692 NAND2X1_LOC_725/Y NAND2X1_LOC_863/a_36_24# 0.07fF
C3693 NOR2X1_LOC_533/Y NOR2X1_LOC_753/Y 0.23fF
C3694 NOR2X1_LOC_209/Y INVX1_LOC_50/Y 0.01fF
C3695 NOR2X1_LOC_21/a_36_216# D_INPUT_5 0.00fF
C3696 INVX1_LOC_85/Y NOR2X1_LOC_306/a_36_216# 0.00fF
C3697 NOR2X1_LOC_705/B NOR2X1_LOC_713/B 0.14fF
C3698 NAND2X1_LOC_849/B NOR2X1_LOC_88/A 0.02fF
C3699 NOR2X1_LOC_464/a_36_216# NOR2X1_LOC_15/Y 0.00fF
C3700 NOR2X1_LOC_590/A INVX1_LOC_94/A 0.07fF
C3701 INVX1_LOC_64/A INVX1_LOC_268/A 0.02fF
C3702 NOR2X1_LOC_791/Y INVX1_LOC_256/Y 0.02fF
C3703 INVX1_LOC_35/A NAND2X1_LOC_662/Y 3.82fF
C3704 INVX1_LOC_90/A NOR2X1_LOC_843/B 0.03fF
C3705 INVX1_LOC_24/Y INVX1_LOC_104/A 0.07fF
C3706 INVX1_LOC_35/A NOR2X1_LOC_730/Y 0.77fF
C3707 INVX1_LOC_304/Y NAND2X1_LOC_579/A 0.07fF
C3708 NOR2X1_LOC_226/A NAND2X1_LOC_391/Y 0.00fF
C3709 INVX1_LOC_45/A NOR2X1_LOC_512/Y 0.01fF
C3710 NOR2X1_LOC_772/B INVX1_LOC_1/Y 0.11fF
C3711 INVX1_LOC_148/A INVX1_LOC_26/Y 0.00fF
C3712 INVX1_LOC_255/Y NOR2X1_LOC_663/A 0.02fF
C3713 INVX1_LOC_21/A NOR2X1_LOC_220/A 0.53fF
C3714 INVX1_LOC_159/A NAND2X1_LOC_195/Y 0.01fF
C3715 NOR2X1_LOC_612/Y NOR2X1_LOC_79/A 0.04fF
C3716 NOR2X1_LOC_754/A INVX1_LOC_91/A 0.06fF
C3717 NOR2X1_LOC_516/B INVX1_LOC_38/Y 0.04fF
C3718 NOR2X1_LOC_719/a_36_216# NOR2X1_LOC_392/Y 0.00fF
C3719 NOR2X1_LOC_13/Y INVX1_LOC_30/A 1.33fF
C3720 INVX1_LOC_13/A INVX1_LOC_5/A 0.26fF
C3721 INVX1_LOC_199/A INVX1_LOC_109/Y 0.01fF
C3722 INPUT_5 NOR2X1_LOC_53/Y 0.03fF
C3723 INVX1_LOC_269/A INVX1_LOC_177/A 0.02fF
C3724 INVX1_LOC_45/Y INVX1_LOC_72/A 0.03fF
C3725 INVX1_LOC_13/Y INVX1_LOC_1/Y 0.04fF
C3726 INVX1_LOC_303/A NOR2X1_LOC_688/Y 0.03fF
C3727 NOR2X1_LOC_453/Y INVX1_LOC_189/Y 0.01fF
C3728 NOR2X1_LOC_609/A NOR2X1_LOC_360/Y 0.01fF
C3729 NOR2X1_LOC_430/A INVX1_LOC_30/A 0.05fF
C3730 NOR2X1_LOC_667/A NOR2X1_LOC_468/Y 0.70fF
C3731 INVX1_LOC_239/A INVX1_LOC_197/Y 0.04fF
C3732 INVX1_LOC_89/A NOR2X1_LOC_392/Y 0.24fF
C3733 NAND2X1_LOC_243/B NAND2X1_LOC_243/Y 0.01fF
C3734 INVX1_LOC_299/A INVX1_LOC_179/Y 0.02fF
C3735 INVX1_LOC_88/A NOR2X1_LOC_362/a_36_216# 0.00fF
C3736 NAND2X1_LOC_348/A NOR2X1_LOC_843/B 0.07fF
C3737 NOR2X1_LOC_790/B NOR2X1_LOC_788/B 0.02fF
C3738 INPUT_0 INVX1_LOC_23/Y 0.07fF
C3739 NOR2X1_LOC_331/B NOR2X1_LOC_127/Y 0.02fF
C3740 INVX1_LOC_21/A NOR2X1_LOC_548/Y 0.11fF
C3741 NAND2X1_LOC_364/A INVX1_LOC_314/Y 0.02fF
C3742 NOR2X1_LOC_164/Y NOR2X1_LOC_48/B 0.14fF
C3743 NAND2X1_LOC_67/Y INVX1_LOC_52/A 0.03fF
C3744 NOR2X1_LOC_487/a_36_216# NOR2X1_LOC_237/Y 0.03fF
C3745 NOR2X1_LOC_364/A NOR2X1_LOC_155/A 0.15fF
C3746 INVX1_LOC_49/A NOR2X1_LOC_703/B 0.82fF
C3747 INVX1_LOC_134/A INVX1_LOC_134/Y 0.00fF
C3748 NAND2X1_LOC_552/A NOR2X1_LOC_246/A 0.01fF
C3749 NAND2X1_LOC_807/B INVX1_LOC_46/A 0.03fF
C3750 INVX1_LOC_75/A NOR2X1_LOC_748/A 0.05fF
C3751 NOR2X1_LOC_419/Y NOR2X1_LOC_360/Y 0.08fF
C3752 NAND2X1_LOC_347/a_36_24# NOR2X1_LOC_103/Y 0.00fF
C3753 NAND2X1_LOC_656/A NAND2X1_LOC_101/a_36_24# 0.02fF
C3754 NAND2X1_LOC_1/Y NAND2X1_LOC_430/B 0.04fF
C3755 INVX1_LOC_182/A INVX1_LOC_53/A 0.23fF
C3756 INVX1_LOC_38/A INVX1_LOC_186/Y 0.07fF
C3757 NOR2X1_LOC_172/Y INVX1_LOC_18/A 0.03fF
C3758 NOR2X1_LOC_68/A NAND2X1_LOC_361/Y 0.07fF
C3759 NOR2X1_LOC_716/B NOR2X1_LOC_360/Y 0.07fF
C3760 NAND2X1_LOC_656/A INVX1_LOC_77/A 0.00fF
C3761 INVX1_LOC_95/Y INVX1_LOC_4/A 1.76fF
C3762 INVX1_LOC_88/A INVX1_LOC_1/Y 0.10fF
C3763 INVX1_LOC_136/A INVX1_LOC_8/A 0.22fF
C3764 NOR2X1_LOC_567/B INVX1_LOC_58/Y 0.01fF
C3765 NOR2X1_LOC_48/B INVX1_LOC_46/A 0.06fF
C3766 INVX1_LOC_27/A NOR2X1_LOC_355/A 0.03fF
C3767 INVX1_LOC_227/Y NOR2X1_LOC_388/Y 0.01fF
C3768 NOR2X1_LOC_590/Y INVX1_LOC_85/Y 0.13fF
C3769 INVX1_LOC_5/A INVX1_LOC_55/Y 0.07fF
C3770 INVX1_LOC_223/Y INVX1_LOC_89/A 0.03fF
C3771 VDD NOR2X1_LOC_554/A 0.00fF
C3772 INVX1_LOC_258/A NAND2X1_LOC_735/B 0.02fF
C3773 INVX1_LOC_38/A INVX1_LOC_261/A 0.18fF
C3774 NOR2X1_LOC_155/A INVX1_LOC_285/A 0.01fF
C3775 NOR2X1_LOC_392/B INVX1_LOC_18/A 0.10fF
C3776 INVX1_LOC_235/A INVX1_LOC_89/A 0.02fF
C3777 NOR2X1_LOC_78/B NOR2X1_LOC_441/Y 0.03fF
C3778 INVX1_LOC_37/A INVX1_LOC_3/Y 0.00fF
C3779 NAND2X1_LOC_391/Y INPUT_1 0.01fF
C3780 NAND2X1_LOC_569/A INVX1_LOC_24/A 0.03fF
C3781 INVX1_LOC_25/A NOR2X1_LOC_391/a_36_216# 0.00fF
C3782 NAND2X1_LOC_579/A NAND2X1_LOC_808/A 0.02fF
C3783 NOR2X1_LOC_264/Y INVX1_LOC_24/A 0.03fF
C3784 NAND2X1_LOC_568/A NAND2X1_LOC_854/B 0.01fF
C3785 NAND2X1_LOC_393/a_36_24# INVX1_LOC_89/A 0.00fF
C3786 INVX1_LOC_64/A NOR2X1_LOC_594/a_36_216# 0.00fF
C3787 NAND2X1_LOC_773/Y INVX1_LOC_171/A 0.01fF
C3788 INVX1_LOC_135/A INVX1_LOC_14/A 0.37fF
C3789 INVX1_LOC_33/A NOR2X1_LOC_577/Y 0.10fF
C3790 INVX1_LOC_94/Y INVX1_LOC_76/A 0.03fF
C3791 INVX1_LOC_27/A NOR2X1_LOC_736/Y 0.08fF
C3792 NAND2X1_LOC_798/B INVX1_LOC_19/A 0.07fF
C3793 NAND2X1_LOC_9/Y INVX1_LOC_286/A 0.07fF
C3794 INVX1_LOC_124/A NAND2X1_LOC_656/A 0.10fF
C3795 NAND2X1_LOC_842/a_36_24# NAND2X1_LOC_474/Y 0.01fF
C3796 INVX1_LOC_161/Y NOR2X1_LOC_686/B 0.06fF
C3797 NOR2X1_LOC_445/Y NOR2X1_LOC_593/Y 0.23fF
C3798 NAND2X1_LOC_794/B NOR2X1_LOC_322/Y 0.08fF
C3799 INVX1_LOC_233/A INVX1_LOC_286/A 0.19fF
C3800 NOR2X1_LOC_195/A NOR2X1_LOC_332/A 0.02fF
C3801 NAND2X1_LOC_243/Y INVX1_LOC_284/A 0.21fF
C3802 INVX1_LOC_132/A NOR2X1_LOC_6/B 0.10fF
C3803 INVX1_LOC_89/Y INVX1_LOC_284/A 0.13fF
C3804 VDD NOR2X1_LOC_89/Y 0.12fF
C3805 NAND2X1_LOC_350/A INVX1_LOC_83/A 0.10fF
C3806 NAND2X1_LOC_350/B INVX1_LOC_159/A 0.01fF
C3807 NAND2X1_LOC_99/Y INVX1_LOC_60/Y 0.08fF
C3808 NAND2X1_LOC_181/Y NAND2X1_LOC_198/B 0.03fF
C3809 NAND2X1_LOC_162/B NAND2X1_LOC_451/Y 0.02fF
C3810 INVX1_LOC_46/A NOR2X1_LOC_438/Y 0.00fF
C3811 INVX1_LOC_33/A NOR2X1_LOC_348/B 0.42fF
C3812 NOR2X1_LOC_9/Y NOR2X1_LOC_81/Y 0.04fF
C3813 INVX1_LOC_41/A INVX1_LOC_104/A 0.17fF
C3814 NOR2X1_LOC_276/Y NAND2X1_LOC_140/A 0.03fF
C3815 INVX1_LOC_223/A NOR2X1_LOC_188/Y 0.01fF
C3816 NOR2X1_LOC_88/Y NOR2X1_LOC_89/A 0.07fF
C3817 INVX1_LOC_90/A NOR2X1_LOC_787/a_36_216# 0.01fF
C3818 INVX1_LOC_8/Y INVX1_LOC_143/A 0.01fF
C3819 NOR2X1_LOC_457/B INVX1_LOC_16/A 0.02fF
C3820 NOR2X1_LOC_798/A INVX1_LOC_286/A 0.36fF
C3821 NOR2X1_LOC_222/Y INVX1_LOC_77/A 0.03fF
C3822 NOR2X1_LOC_273/Y NAND2X1_LOC_831/a_36_24# 0.01fF
C3823 INVX1_LOC_233/A INVX1_LOC_95/A 0.00fF
C3824 NAND2X1_LOC_139/A NAND2X1_LOC_141/A 0.02fF
C3825 NAND2X1_LOC_792/B NAND2X1_LOC_792/a_36_24# 0.00fF
C3826 INVX1_LOC_272/A INVX1_LOC_63/A 0.07fF
C3827 INVX1_LOC_111/Y NOR2X1_LOC_388/Y 0.02fF
C3828 NOR2X1_LOC_590/A NOR2X1_LOC_768/a_36_216# 0.00fF
C3829 NAND2X1_LOC_182/A NAND2X1_LOC_477/A 0.17fF
C3830 INVX1_LOC_31/A INVX1_LOC_20/Y 0.03fF
C3831 NOR2X1_LOC_772/B INVX1_LOC_93/Y 0.96fF
C3832 INVX1_LOC_64/A INVX1_LOC_95/Y 0.01fF
C3833 NOR2X1_LOC_89/A INVX1_LOC_84/A 0.41fF
C3834 INVX1_LOC_58/A INVX1_LOC_37/A 0.10fF
C3835 NOR2X1_LOC_263/a_36_216# INVX1_LOC_124/A 0.03fF
C3836 NOR2X1_LOC_78/B NOR2X1_LOC_142/Y 0.76fF
C3837 INVX1_LOC_72/A NOR2X1_LOC_71/Y 0.08fF
C3838 INVX1_LOC_14/A NOR2X1_LOC_391/B 0.03fF
C3839 INVX1_LOC_303/A INVX1_LOC_1/Y 0.21fF
C3840 INVX1_LOC_50/Y NAND2X1_LOC_642/Y 0.02fF
C3841 INVX1_LOC_269/A INVX1_LOC_285/Y 0.10fF
C3842 INVX1_LOC_256/A NOR2X1_LOC_310/a_36_216# 0.01fF
C3843 INVX1_LOC_13/Y INVX1_LOC_93/Y 0.23fF
C3844 INVX1_LOC_227/A INVX1_LOC_94/A 0.07fF
C3845 INVX1_LOC_89/A NOR2X1_LOC_86/Y 0.01fF
C3846 INVX1_LOC_33/A NOR2X1_LOC_325/A 0.00fF
C3847 NAND2X1_LOC_803/B INVX1_LOC_144/A 0.02fF
C3848 NOR2X1_LOC_431/Y INVX1_LOC_10/A 0.02fF
C3849 NAND2X1_LOC_656/a_36_24# NOR2X1_LOC_360/Y 0.06fF
C3850 INVX1_LOC_33/A INVX1_LOC_22/A 0.25fF
C3851 INVX1_LOC_64/A NOR2X1_LOC_305/Y 0.05fF
C3852 NAND2X1_LOC_833/Y INVX1_LOC_16/A 0.03fF
C3853 INVX1_LOC_132/A INVX1_LOC_30/Y 0.03fF
C3854 NOR2X1_LOC_509/A NOR2X1_LOC_340/A 0.03fF
C3855 NOR2X1_LOC_331/B NOR2X1_LOC_383/B 0.07fF
C3856 NOR2X1_LOC_448/Y INVX1_LOC_91/A 0.01fF
C3857 INVX1_LOC_34/A INVX1_LOC_232/A 0.08fF
C3858 INVX1_LOC_90/A INVX1_LOC_18/A 3.68fF
C3859 NOR2X1_LOC_431/a_36_216# NOR2X1_LOC_130/A 0.00fF
C3860 NOR2X1_LOC_272/Y NOR2X1_LOC_657/B 0.30fF
C3861 NOR2X1_LOC_15/Y INVX1_LOC_98/A 0.01fF
C3862 NOR2X1_LOC_160/B NOR2X1_LOC_721/Y 0.01fF
C3863 INVX1_LOC_226/Y NOR2X1_LOC_720/B 0.04fF
C3864 D_INPUT_1 NOR2X1_LOC_536/A 3.70fF
C3865 NOR2X1_LOC_15/Y NOR2X1_LOC_78/A 3.34fF
C3866 NOR2X1_LOC_389/B INVX1_LOC_18/A 0.07fF
C3867 NAND2X1_LOC_303/Y NOR2X1_LOC_45/B 0.10fF
C3868 INVX1_LOC_5/A NOR2X1_LOC_357/Y 0.12fF
C3869 NOR2X1_LOC_409/B NAND2X1_LOC_810/B 0.01fF
C3870 INVX1_LOC_243/Y NAND2X1_LOC_637/Y 0.00fF
C3871 NOR2X1_LOC_590/A INVX1_LOC_144/A 0.08fF
C3872 INVX1_LOC_104/A NOR2X1_LOC_211/A 0.03fF
C3873 INVX1_LOC_88/A NOR2X1_LOC_318/B 0.10fF
C3874 NOR2X1_LOC_304/Y NAND2X1_LOC_453/A 0.02fF
C3875 INVX1_LOC_22/A NAND2X1_LOC_466/A 0.08fF
C3876 INVX1_LOC_289/Y NAND2X1_LOC_655/A 0.07fF
C3877 INVX1_LOC_34/A NOR2X1_LOC_383/Y 0.07fF
C3878 NOR2X1_LOC_68/A NAND2X1_LOC_654/B 0.01fF
C3879 INVX1_LOC_45/Y INVX1_LOC_313/Y 0.05fF
C3880 NOR2X1_LOC_637/B NOR2X1_LOC_130/A 0.46fF
C3881 INVX1_LOC_155/Y INVX1_LOC_10/A 0.03fF
C3882 NOR2X1_LOC_637/Y INVX1_LOC_90/A 0.01fF
C3883 INVX1_LOC_269/A INVX1_LOC_65/A 0.10fF
C3884 NOR2X1_LOC_468/Y INVX1_LOC_304/A 0.02fF
C3885 NOR2X1_LOC_490/Y NOR2X1_LOC_522/Y 0.08fF
C3886 NOR2X1_LOC_401/a_36_216# NAND2X1_LOC_181/Y 0.00fF
C3887 INVX1_LOC_58/A INVX1_LOC_157/Y 0.06fF
C3888 NOR2X1_LOC_653/B VDD -0.00fF
C3889 NAND2X1_LOC_741/B INPUT_0 0.03fF
C3890 NAND2X1_LOC_574/A NOR2X1_LOC_415/Y 0.16fF
C3891 INVX1_LOC_269/A INVX1_LOC_316/A -0.02fF
C3892 INVX1_LOC_34/A NOR2X1_LOC_366/Y 0.00fF
C3893 NOR2X1_LOC_316/a_36_216# NAND2X1_LOC_572/B 0.01fF
C3894 INVX1_LOC_59/A INVX1_LOC_20/A 0.05fF
C3895 NAND2X1_LOC_276/Y D_INPUT_0 0.06fF
C3896 D_INPUT_1 NOR2X1_LOC_655/Y 0.17fF
C3897 INVX1_LOC_172/A INVX1_LOC_90/A 0.09fF
C3898 NOR2X1_LOC_67/A NOR2X1_LOC_121/a_36_216# 0.00fF
C3899 INVX1_LOC_135/A INVX1_LOC_217/Y -0.01fF
C3900 INVX1_LOC_206/A INVX1_LOC_101/A 0.01fF
C3901 INVX1_LOC_249/A NOR2X1_LOC_736/Y 0.01fF
C3902 NAND2X1_LOC_773/Y INVX1_LOC_20/A 0.49fF
C3903 NAND2X1_LOC_785/Y NAND2X1_LOC_795/Y 0.04fF
C3904 INVX1_LOC_255/Y NOR2X1_LOC_537/Y 0.08fF
C3905 D_INPUT_1 NAND2X1_LOC_93/B 0.04fF
C3906 NOR2X1_LOC_590/A NOR2X1_LOC_845/A 0.01fF
C3907 NOR2X1_LOC_606/Y INVX1_LOC_123/A 0.01fF
C3908 NAND2X1_LOC_840/B NAND2X1_LOC_834/a_36_24# 0.02fF
C3909 INVX1_LOC_233/A INVX1_LOC_54/A 0.12fF
C3910 NAND2X1_LOC_647/B INVX1_LOC_29/A 0.03fF
C3911 NOR2X1_LOC_536/A NOR2X1_LOC_652/Y 0.07fF
C3912 NOR2X1_LOC_89/A INVX1_LOC_15/A 0.06fF
C3913 NOR2X1_LOC_114/Y NOR2X1_LOC_116/a_36_216# -0.00fF
C3914 INVX1_LOC_233/Y NOR2X1_LOC_629/Y 0.02fF
C3915 NAND2X1_LOC_198/B NAND2X1_LOC_138/a_36_24# 0.06fF
C3916 NOR2X1_LOC_286/Y INVX1_LOC_143/Y 0.03fF
C3917 NOR2X1_LOC_238/Y INVX1_LOC_282/A 0.02fF
C3918 NOR2X1_LOC_216/B INVX1_LOC_29/Y 0.01fF
C3919 NOR2X1_LOC_596/A NAND2X1_LOC_51/B 0.03fF
C3920 NOR2X1_LOC_793/A VDD 0.24fF
C3921 INVX1_LOC_10/A NOR2X1_LOC_822/Y 0.29fF
C3922 INVX1_LOC_28/A NAND2X1_LOC_833/Y 0.05fF
C3923 INVX1_LOC_77/A D_INPUT_4 0.07fF
C3924 NAND2X1_LOC_726/Y INVX1_LOC_22/A 0.08fF
C3925 NOR2X1_LOC_15/Y NOR2X1_LOC_176/a_36_216# 0.00fF
C3926 INVX1_LOC_10/A NOR2X1_LOC_131/A 0.01fF
C3927 INVX1_LOC_206/A NOR2X1_LOC_355/A 0.00fF
C3928 NOR2X1_LOC_459/B INVX1_LOC_175/Y 0.26fF
C3929 INVX1_LOC_43/Y INVX1_LOC_95/Y 0.05fF
C3930 NOR2X1_LOC_763/A NAND2X1_LOC_635/a_36_24# 0.00fF
C3931 NOR2X1_LOC_55/a_36_216# NAND2X1_LOC_773/B 0.01fF
C3932 INVX1_LOC_209/Y NOR2X1_LOC_380/Y 0.22fF
C3933 INVX1_LOC_69/Y NOR2X1_LOC_168/Y 0.01fF
C3934 NOR2X1_LOC_596/A INVX1_LOC_311/A 0.29fF
C3935 NOR2X1_LOC_667/A NAND2X1_LOC_795/Y 0.01fF
C3936 NOR2X1_LOC_655/B INVX1_LOC_83/A 0.10fF
C3937 INVX1_LOC_222/Y INVX1_LOC_9/A 0.03fF
C3938 NAND2X1_LOC_90/a_36_24# INVX1_LOC_3/A 0.00fF
C3939 NOR2X1_LOC_216/Y INVX1_LOC_155/A 0.10fF
C3940 INVX1_LOC_293/A INVX1_LOC_76/A 0.01fF
C3941 NOR2X1_LOC_666/Y NAND2X1_LOC_472/Y 0.01fF
C3942 INVX1_LOC_279/A NOR2X1_LOC_131/Y 0.01fF
C3943 NOR2X1_LOC_151/Y NOR2X1_LOC_717/a_36_216# 0.00fF
C3944 NAND2X1_LOC_338/B NOR2X1_LOC_71/Y 0.85fF
C3945 NOR2X1_LOC_254/Y NOR2X1_LOC_197/Y 0.03fF
C3946 NAND2X1_LOC_391/Y INVX1_LOC_118/A 0.07fF
C3947 INVX1_LOC_14/A NOR2X1_LOC_813/Y 0.07fF
C3948 D_INPUT_1 NOR2X1_LOC_649/B 0.15fF
C3949 NAND2X1_LOC_364/A NOR2X1_LOC_557/A 0.00fF
C3950 INVX1_LOC_170/A NOR2X1_LOC_124/A 0.03fF
C3951 NOR2X1_LOC_673/A NOR2X1_LOC_416/A 0.07fF
C3952 D_INPUT_1 INVX1_LOC_3/A 1.03fF
C3953 INVX1_LOC_27/A INVX1_LOC_127/A 0.03fF
C3954 NAND2X1_LOC_550/A VDD -0.00fF
C3955 NOR2X1_LOC_497/a_36_216# NAND2X1_LOC_489/Y 0.00fF
C3956 NOR2X1_LOC_246/A NOR2X1_LOC_773/Y 0.03fF
C3957 NAND2X1_LOC_93/B NOR2X1_LOC_652/Y 0.03fF
C3958 INVX1_LOC_5/A INVX1_LOC_260/A 0.01fF
C3959 NOR2X1_LOC_160/B VDD 2.98fF
C3960 NOR2X1_LOC_690/A INVX1_LOC_91/Y 0.01fF
C3961 INVX1_LOC_57/A NAND2X1_LOC_773/B 0.07fF
C3962 NOR2X1_LOC_65/Y INVX1_LOC_272/A 0.01fF
C3963 INVX1_LOC_279/A NOR2X1_LOC_589/A 0.07fF
C3964 INVX1_LOC_14/A INVX1_LOC_280/A 0.22fF
C3965 NOR2X1_LOC_598/B NOR2X1_LOC_814/A 0.26fF
C3966 NOR2X1_LOC_134/Y NOR2X1_LOC_290/a_36_216# 0.00fF
C3967 INVX1_LOC_14/A NOR2X1_LOC_94/Y 0.13fF
C3968 NOR2X1_LOC_548/Y NOR2X1_LOC_565/B 0.02fF
C3969 NOR2X1_LOC_441/Y INVX1_LOC_46/A 0.08fF
C3970 INVX1_LOC_89/A INVX1_LOC_25/Y 0.23fF
C3971 INVX1_LOC_13/A NOR2X1_LOC_332/A 0.18fF
C3972 NOR2X1_LOC_860/B NOR2X1_LOC_78/A 0.07fF
C3973 INVX1_LOC_16/A NOR2X1_LOC_76/A 0.02fF
C3974 INVX1_LOC_1/A NOR2X1_LOC_641/Y 0.01fF
C3975 NAND2X1_LOC_116/A INPUT_0 3.80fF
C3976 NOR2X1_LOC_78/B INVX1_LOC_182/A 0.13fF
C3977 NOR2X1_LOC_717/Y INVX1_LOC_139/Y 0.00fF
C3978 INVX1_LOC_49/A INVX1_LOC_91/A 0.87fF
C3979 INVX1_LOC_271/Y INVX1_LOC_4/A 0.07fF
C3980 NOR2X1_LOC_561/Y INVX1_LOC_66/A -0.02fF
C3981 INVX1_LOC_314/Y NOR2X1_LOC_405/A 0.02fF
C3982 INVX1_LOC_2/A INVX1_LOC_79/A 0.07fF
C3983 NOR2X1_LOC_74/A NOR2X1_LOC_709/A 0.10fF
C3984 NOR2X1_LOC_646/B INVX1_LOC_42/A 0.00fF
C3985 INVX1_LOC_284/A NAND2X1_LOC_205/A 0.04fF
C3986 NOR2X1_LOC_455/a_36_216# INVX1_LOC_206/Y 0.00fF
C3987 INVX1_LOC_303/A INVX1_LOC_93/Y 0.04fF
C3988 INVX1_LOC_174/A NOR2X1_LOC_450/A 0.01fF
C3989 NOR2X1_LOC_187/Y INVX1_LOC_92/A 0.01fF
C3990 NOR2X1_LOC_261/Y NOR2X1_LOC_89/A 0.12fF
C3991 INVX1_LOC_83/A NOR2X1_LOC_99/B 0.07fF
C3992 NOR2X1_LOC_11/a_36_216# INPUT_4 0.01fF
C3993 NAND2X1_LOC_354/Y NOR2X1_LOC_447/B 0.03fF
C3994 NOR2X1_LOC_709/A NOR2X1_LOC_9/Y 0.35fF
C3995 NOR2X1_LOC_690/A NOR2X1_LOC_45/B 0.07fF
C3996 NOR2X1_LOC_321/Y NOR2X1_LOC_841/A 0.03fF
C3997 NOR2X1_LOC_32/B INVX1_LOC_12/A 0.07fF
C3998 INVX1_LOC_78/A NOR2X1_LOC_158/Y 0.30fF
C3999 NOR2X1_LOC_717/Y INVX1_LOC_10/Y 0.03fF
C4000 NOR2X1_LOC_556/a_36_216# NOR2X1_LOC_303/Y 0.00fF
C4001 NOR2X1_LOC_109/a_36_216# INVX1_LOC_29/A 0.02fF
C4002 INVX1_LOC_278/A NOR2X1_LOC_89/A 1.06fF
C4003 INVX1_LOC_83/A NOR2X1_LOC_846/B 0.03fF
C4004 INVX1_LOC_26/A NOR2X1_LOC_394/Y 0.01fF
C4005 INVX1_LOC_178/A NAND2X1_LOC_489/Y 0.03fF
C4006 NOR2X1_LOC_725/A INVX1_LOC_76/Y 0.04fF
C4007 NOR2X1_LOC_220/A INVX1_LOC_311/A 0.04fF
C4008 INVX1_LOC_53/A NOR2X1_LOC_850/B 0.16fF
C4009 INVX1_LOC_11/A NOR2X1_LOC_88/Y 0.03fF
C4010 NOR2X1_LOC_329/B NAND2X1_LOC_796/Y 0.01fF
C4011 NOR2X1_LOC_6/B NAND2X1_LOC_642/Y 0.03fF
C4012 INPUT_0 INVX1_LOC_232/A 0.12fF
C4013 NAND2X1_LOC_332/Y NAND2X1_LOC_468/B 0.00fF
C4014 INVX1_LOC_18/A NAND2X1_LOC_849/B 0.10fF
C4015 INVX1_LOC_233/A NOR2X1_LOC_48/B 0.01fF
C4016 INVX1_LOC_2/A INVX1_LOC_91/A 0.48fF
C4017 NAND2X1_LOC_391/a_36_24# NOR2X1_LOC_536/A 0.00fF
C4018 INVX1_LOC_18/A INVX1_LOC_38/A 0.27fF
C4019 NOR2X1_LOC_82/A NAND2X1_LOC_141/Y 0.02fF
C4020 INVX1_LOC_63/A NOR2X1_LOC_271/B 0.03fF
C4021 NOR2X1_LOC_486/Y NOR2X1_LOC_348/B 0.09fF
C4022 NOR2X1_LOC_567/B NOR2X1_LOC_326/Y 0.00fF
C4023 NOR2X1_LOC_91/A NOR2X1_LOC_301/A 0.06fF
C4024 NOR2X1_LOC_226/A INVX1_LOC_91/A 0.19fF
C4025 INVX1_LOC_50/A NAND2X1_LOC_454/Y 0.07fF
C4026 NOR2X1_LOC_590/A NOR2X1_LOC_155/A 0.07fF
C4027 NOR2X1_LOC_644/A INVX1_LOC_313/Y 0.67fF
C4028 NOR2X1_LOC_383/Y INPUT_0 0.23fF
C4029 INVX1_LOC_162/A INVX1_LOC_76/A 0.04fF
C4030 NAND2X1_LOC_33/Y NOR2X1_LOC_24/Y 0.10fF
C4031 INVX1_LOC_30/A NOR2X1_LOC_640/Y 0.10fF
C4032 D_INPUT_6 INPUT_7 0.68fF
C4033 INVX1_LOC_11/A INVX1_LOC_84/A 0.13fF
C4034 INVX1_LOC_75/A INVX1_LOC_150/A 0.01fF
C4035 NOR2X1_LOC_672/Y NAND2X1_LOC_721/A 0.00fF
C4036 INVX1_LOC_2/A INVX1_LOC_11/Y 0.04fF
C4037 NOR2X1_LOC_142/Y INVX1_LOC_46/A 0.01fF
C4038 INVX1_LOC_49/A NOR2X1_LOC_698/Y 0.19fF
C4039 NOR2X1_LOC_759/Y NOR2X1_LOC_142/a_36_216# 0.00fF
C4040 NOR2X1_LOC_637/Y INVX1_LOC_38/A 0.03fF
C4041 INVX1_LOC_45/A INVX1_LOC_179/A 0.02fF
C4042 NAND2X1_LOC_656/A INVX1_LOC_9/A 0.06fF
C4043 NOR2X1_LOC_315/Y INVX1_LOC_76/A 0.07fF
C4044 INVX1_LOC_18/A NOR2X1_LOC_51/A 0.01fF
C4045 NOR2X1_LOC_351/a_36_216# NOR2X1_LOC_351/Y 0.00fF
C4046 INVX1_LOC_89/A INVX1_LOC_75/A 0.42fF
C4047 NAND2X1_LOC_734/a_36_24# NAND2X1_LOC_721/A 0.00fF
C4048 INVX1_LOC_5/A INVX1_LOC_32/A 0.57fF
C4049 NOR2X1_LOC_161/Y INVX1_LOC_91/A 0.00fF
C4050 NOR2X1_LOC_344/a_36_216# INVX1_LOC_37/A 0.00fF
C4051 INVX1_LOC_90/A INVX1_LOC_31/Y 0.09fF
C4052 INVX1_LOC_119/A NAND2X1_LOC_453/A 0.64fF
C4053 INVX1_LOC_172/A INVX1_LOC_38/A 0.02fF
C4054 NAND2X1_LOC_631/a_36_24# NOR2X1_LOC_536/A 0.00fF
C4055 NAND2X1_LOC_350/B NOR2X1_LOC_56/Y 0.29fF
C4056 NAND2X1_LOC_563/A INVX1_LOC_316/A 0.12fF
C4057 INVX1_LOC_207/Y NAND2X1_LOC_463/B 0.00fF
C4058 INVX1_LOC_28/A INVX1_LOC_73/A 0.07fF
C4059 INVX1_LOC_11/A NAND2X1_LOC_651/B 0.03fF
C4060 NAND2X1_LOC_508/A INVX1_LOC_75/A 0.02fF
C4061 NAND2X1_LOC_703/Y NOR2X1_LOC_48/B 0.27fF
C4062 INVX1_LOC_189/A VDD 0.00fF
C4063 NOR2X1_LOC_483/B INVX1_LOC_186/Y 0.01fF
C4064 INVX1_LOC_90/A NOR2X1_LOC_548/A 0.05fF
C4065 NOR2X1_LOC_486/Y INVX1_LOC_22/A 0.00fF
C4066 NOR2X1_LOC_78/A NOR2X1_LOC_97/B 0.10fF
C4067 NOR2X1_LOC_655/B INVX1_LOC_46/A 0.30fF
C4068 INVX1_LOC_217/Y INVX1_LOC_280/A 0.64fF
C4069 NOR2X1_LOC_383/B NOR2X1_LOC_493/A 0.01fF
C4070 NOR2X1_LOC_772/B INVX1_LOC_87/A 0.10fF
C4071 INVX1_LOC_30/Y NAND2X1_LOC_642/Y 0.14fF
C4072 INVX1_LOC_36/A NOR2X1_LOC_673/A 0.03fF
C4073 NOR2X1_LOC_781/a_36_216# INVX1_LOC_91/A 0.00fF
C4074 INVX1_LOC_52/A INVX1_LOC_76/A 0.02fF
C4075 NAND2X1_LOC_350/B VDD 0.22fF
C4076 INVX1_LOC_298/Y NOR2X1_LOC_665/Y 0.05fF
C4077 NOR2X1_LOC_775/Y INPUT_0 0.64fF
C4078 INVX1_LOC_71/A INVX1_LOC_179/A 0.00fF
C4079 NOR2X1_LOC_591/Y NOR2X1_LOC_536/A 0.29fF
C4080 NOR2X1_LOC_186/Y INVX1_LOC_273/A 0.10fF
C4081 INVX1_LOC_13/Y INVX1_LOC_87/A 0.03fF
C4082 VDD NAND2X1_LOC_853/Y 1.95fF
C4083 INVX1_LOC_286/A NAND2X1_LOC_842/B 0.39fF
C4084 INVX1_LOC_208/A VDD 2.50fF
C4085 NOR2X1_LOC_240/Y NOR2X1_LOC_342/B 0.02fF
C4086 NAND2X1_LOC_773/Y INVX1_LOC_4/A 0.17fF
C4087 NOR2X1_LOC_516/B VDD 3.93fF
C4088 NOR2X1_LOC_433/A NOR2X1_LOC_88/Y 0.03fF
C4089 NOR2X1_LOC_238/a_36_216# INVX1_LOC_119/Y -0.00fF
C4090 INPUT_1 INVX1_LOC_91/A 0.01fF
C4091 INVX1_LOC_224/A INVX1_LOC_15/A 0.03fF
C4092 NOR2X1_LOC_309/Y NOR2X1_LOC_612/Y 0.02fF
C4093 INVX1_LOC_178/A NAND2X1_LOC_175/Y 0.10fF
C4094 INVX1_LOC_155/Y INVX1_LOC_307/A 0.00fF
C4095 NAND2X1_LOC_276/Y INVX1_LOC_46/Y 0.07fF
C4096 D_INPUT_2 NOR2X1_LOC_649/B 0.07fF
C4097 NOR2X1_LOC_399/A NOR2X1_LOC_629/Y 0.00fF
C4098 INVX1_LOC_11/A INVX1_LOC_15/A 1.48fF
C4099 NAND2X1_LOC_30/Y NAND2X1_LOC_429/a_36_24# 0.00fF
C4100 NOR2X1_LOC_403/B INVX1_LOC_3/A 0.19fF
C4101 D_INPUT_2 INVX1_LOC_3/A 0.00fF
C4102 INVX1_LOC_269/A INVX1_LOC_4/Y 1.45fF
C4103 NAND2X1_LOC_337/B INVX1_LOC_32/A 0.08fF
C4104 INVX1_LOC_24/A NOR2X1_LOC_662/A 0.01fF
C4105 NOR2X1_LOC_537/a_36_216# INVX1_LOC_22/A 0.00fF
C4106 NOR2X1_LOC_264/Y NOR2X1_LOC_197/B 0.02fF
C4107 NOR2X1_LOC_433/A INVX1_LOC_84/A 0.40fF
C4108 INVX1_LOC_28/A NAND2X1_LOC_729/B 0.01fF
C4109 NAND2X1_LOC_842/B INVX1_LOC_95/A 0.00fF
C4110 NOR2X1_LOC_540/B INVX1_LOC_313/Y 0.00fF
C4111 NOR2X1_LOC_52/B NOR2X1_LOC_88/Y 0.03fF
C4112 NOR2X1_LOC_272/Y INVX1_LOC_271/A 0.04fF
C4113 NOR2X1_LOC_180/B NOR2X1_LOC_35/Y 0.10fF
C4114 NOR2X1_LOC_740/Y NOR2X1_LOC_307/Y 0.02fF
C4115 INVX1_LOC_33/A NAND2X1_LOC_476/Y 0.06fF
C4116 INVX1_LOC_143/A NAND2X1_LOC_487/a_36_24# 0.00fF
C4117 INVX1_LOC_69/Y NOR2X1_LOC_548/a_36_216# 0.01fF
C4118 NOR2X1_LOC_152/Y INVX1_LOC_264/A 0.01fF
C4119 INVX1_LOC_285/Y NOR2X1_LOC_741/A 0.00fF
C4120 NOR2X1_LOC_351/Y INVX1_LOC_22/A 0.77fF
C4121 NOR2X1_LOC_67/A NOR2X1_LOC_101/a_36_216# 0.00fF
C4122 NOR2X1_LOC_516/B NOR2X1_LOC_846/a_36_216# 0.00fF
C4123 NAND2X1_LOC_337/B NAND2X1_LOC_175/Y 0.14fF
C4124 NOR2X1_LOC_816/A NAND2X1_LOC_175/Y 1.09fF
C4125 NOR2X1_LOC_91/A INVX1_LOC_17/A 0.10fF
C4126 INVX1_LOC_17/A NOR2X1_LOC_668/Y 0.01fF
C4127 NOR2X1_LOC_52/B INVX1_LOC_84/A 0.07fF
C4128 NOR2X1_LOC_706/Y INVX1_LOC_91/A 0.01fF
C4129 D_INPUT_1 NOR2X1_LOC_348/Y 0.13fF
C4130 NOR2X1_LOC_262/Y NOR2X1_LOC_89/A 0.13fF
C4131 INVX1_LOC_33/A NOR2X1_LOC_777/B 11.16fF
C4132 INPUT_0 INVX1_LOC_74/Y 0.01fF
C4133 INVX1_LOC_35/A NOR2X1_LOC_454/Y 0.07fF
C4134 INVX1_LOC_22/A INVX1_LOC_241/Y 0.03fF
C4135 INVX1_LOC_59/A INVX1_LOC_64/A 0.00fF
C4136 INVX1_LOC_155/Y INVX1_LOC_12/A 0.03fF
C4137 INVX1_LOC_36/A NOR2X1_LOC_409/B 0.03fF
C4138 NOR2X1_LOC_272/Y NAND2X1_LOC_214/B 0.00fF
C4139 INVX1_LOC_17/A INVX1_LOC_23/A 2.59fF
C4140 NOR2X1_LOC_366/B NOR2X1_LOC_127/Y 0.02fF
C4141 NAND2X1_LOC_858/B INVX1_LOC_20/A 0.00fF
C4142 INVX1_LOC_256/A D_INPUT_1 0.01fF
C4143 NOR2X1_LOC_261/Y INVX1_LOC_11/A 0.04fF
C4144 NOR2X1_LOC_557/A NOR2X1_LOC_405/A 0.00fF
C4145 INVX1_LOC_39/A NAND2X1_LOC_391/Y 0.11fF
C4146 NOR2X1_LOC_272/Y INVX1_LOC_27/A 0.03fF
C4147 NOR2X1_LOC_647/B D_INPUT_1 0.01fF
C4148 NOR2X1_LOC_433/A INVX1_LOC_15/A 0.14fF
C4149 INVX1_LOC_120/A NAND2X1_LOC_86/a_36_24# 0.00fF
C4150 NOR2X1_LOC_474/A INVX1_LOC_15/A 0.03fF
C4151 NOR2X1_LOC_411/a_36_216# INVX1_LOC_269/A 0.00fF
C4152 NAND2X1_LOC_555/Y INVX1_LOC_23/A 0.03fF
C4153 INVX1_LOC_232/Y NAND2X1_LOC_82/Y 0.29fF
C4154 NOR2X1_LOC_593/Y INVX1_LOC_15/A 0.03fF
C4155 NOR2X1_LOC_329/B INVX1_LOC_9/A 0.04fF
C4156 NAND2X1_LOC_842/B INVX1_LOC_54/A 0.00fF
C4157 NAND2X1_LOC_342/Y INVX1_LOC_29/A 0.00fF
C4158 NOR2X1_LOC_186/Y NOR2X1_LOC_15/Y 0.05fF
C4159 NOR2X1_LOC_16/Y NOR2X1_LOC_89/A 0.01fF
C4160 INVX1_LOC_72/Y INVX1_LOC_23/Y 0.02fF
C4161 NOR2X1_LOC_598/B NOR2X1_LOC_590/A 0.12fF
C4162 NAND2X1_LOC_213/A INVX1_LOC_27/A 0.04fF
C4163 INVX1_LOC_11/A NOR2X1_LOC_223/B 0.01fF
C4164 D_INPUT_1 NOR2X1_LOC_606/Y 0.01fF
C4165 NAND2X1_LOC_9/Y INVX1_LOC_218/Y 0.03fF
C4166 INVX1_LOC_208/A INVX1_LOC_133/A 0.23fF
C4167 NOR2X1_LOC_152/Y NOR2X1_LOC_158/Y 0.07fF
C4168 INVX1_LOC_315/Y VDD 0.35fF
C4169 INVX1_LOC_236/A INVX1_LOC_42/A 0.00fF
C4170 NOR2X1_LOC_315/Y INVX1_LOC_127/Y 0.02fF
C4171 NOR2X1_LOC_757/A NAND2X1_LOC_475/Y 0.04fF
C4172 INVX1_LOC_91/A NOR2X1_LOC_586/Y 0.42fF
C4173 NAND2X1_LOC_84/Y NAND2X1_LOC_437/a_36_24# 0.00fF
C4174 INVX1_LOC_303/A INVX1_LOC_87/A -0.04fF
C4175 INVX1_LOC_90/A NAND2X1_LOC_489/a_36_24# 0.01fF
C4176 NOR2X1_LOC_144/Y INVX1_LOC_4/A 0.04fF
C4177 INVX1_LOC_72/A NAND2X1_LOC_205/A 0.02fF
C4178 NOR2X1_LOC_328/Y NOR2X1_LOC_11/Y 0.01fF
C4179 INVX1_LOC_50/A NOR2X1_LOC_68/A 4.89fF
C4180 INVX1_LOC_233/A NOR2X1_LOC_441/Y 0.00fF
C4181 NOR2X1_LOC_82/A INVX1_LOC_13/Y 2.82fF
C4182 INVX1_LOC_51/A INVX1_LOC_22/Y 0.15fF
C4183 NOR2X1_LOC_52/B INVX1_LOC_15/A 0.17fF
C4184 INVX1_LOC_256/A NOR2X1_LOC_652/Y 0.07fF
C4185 INVX1_LOC_269/A NOR2X1_LOC_790/A 0.03fF
C4186 NOR2X1_LOC_528/Y NOR2X1_LOC_111/A 0.01fF
C4187 INPUT_3 INVX1_LOC_5/A 0.07fF
C4188 NOR2X1_LOC_419/Y INVX1_LOC_26/A 0.16fF
C4189 NAND2X1_LOC_348/A NOR2X1_LOC_860/Y 0.01fF
C4190 NOR2X1_LOC_78/B NOR2X1_LOC_850/B 0.01fF
C4191 NAND2X1_LOC_374/Y NOR2X1_LOC_754/A 0.01fF
C4192 INVX1_LOC_45/A NOR2X1_LOC_405/Y 0.01fF
C4193 NOR2X1_LOC_748/Y NAND2X1_LOC_74/B 0.05fF
C4194 NOR2X1_LOC_74/A NOR2X1_LOC_489/A 0.03fF
C4195 NOR2X1_LOC_15/Y NAND2X1_LOC_724/A 0.07fF
C4196 NAND2X1_LOC_796/a_36_24# NOR2X1_LOC_109/Y 0.01fF
C4197 NOR2X1_LOC_716/B INVX1_LOC_26/A 0.14fF
C4198 INVX1_LOC_24/A INVX1_LOC_57/A 5.48fF
C4199 NAND2X1_LOC_88/a_36_24# INVX1_LOC_15/A 0.00fF
C4200 NOR2X1_LOC_228/a_36_216# INVX1_LOC_26/Y 0.00fF
C4201 NAND2X1_LOC_808/A NAND2X1_LOC_604/a_36_24# 0.00fF
C4202 NOR2X1_LOC_32/B INVX1_LOC_217/A 0.08fF
C4203 NAND2X1_LOC_693/a_36_24# INVX1_LOC_92/A 0.01fF
C4204 INVX1_LOC_309/A INVX1_LOC_118/A 0.00fF
C4205 INVX1_LOC_13/A NOR2X1_LOC_847/A 0.30fF
C4206 NOR2X1_LOC_773/Y INVX1_LOC_32/A 0.10fF
C4207 INPUT_1 INVX1_LOC_203/A 0.03fF
C4208 INVX1_LOC_13/A INVX1_LOC_42/A 0.12fF
C4209 NAND2X1_LOC_578/B NAND2X1_LOC_618/Y 0.58fF
C4210 INVX1_LOC_21/A NOR2X1_LOC_550/a_36_216# 0.01fF
C4211 INVX1_LOC_287/A INVX1_LOC_33/A 0.04fF
C4212 INVX1_LOC_236/A INVX1_LOC_78/A 0.17fF
C4213 VDD NAND2X1_LOC_211/Y 0.22fF
C4214 INVX1_LOC_34/A INVX1_LOC_112/Y 0.03fF
C4215 NOR2X1_LOC_388/Y NOR2X1_LOC_383/B 0.06fF
C4216 INVX1_LOC_91/A INVX1_LOC_118/A 1.00fF
C4217 NOR2X1_LOC_68/A NAND2X1_LOC_749/a_36_24# 0.00fF
C4218 NOR2X1_LOC_557/Y INVX1_LOC_57/A 0.29fF
C4219 NOR2X1_LOC_250/Y NOR2X1_LOC_250/A 0.05fF
C4220 INVX1_LOC_101/Y INVX1_LOC_292/A 0.01fF
C4221 NOR2X1_LOC_361/B NOR2X1_LOC_160/B 0.03fF
C4222 INVX1_LOC_35/A INVX1_LOC_77/A 13.26fF
C4223 NOR2X1_LOC_246/Y INVX1_LOC_29/A 0.07fF
C4224 INVX1_LOC_89/A NAND2X1_LOC_291/B 0.04fF
C4225 NOR2X1_LOC_619/a_36_216# NOR2X1_LOC_419/Y 0.00fF
C4226 NAND2X1_LOC_103/a_36_24# NOR2X1_LOC_831/B 0.00fF
C4227 INVX1_LOC_98/Y INVX1_LOC_26/A 0.01fF
C4228 INVX1_LOC_11/Y INVX1_LOC_118/A 0.03fF
C4229 INVX1_LOC_27/A NAND2X1_LOC_364/A 0.03fF
C4230 NOR2X1_LOC_551/B INVX1_LOC_53/A 0.03fF
C4231 NOR2X1_LOC_679/Y INVX1_LOC_161/Y 0.02fF
C4232 NOR2X1_LOC_773/Y NAND2X1_LOC_175/Y 0.01fF
C4233 NOR2X1_LOC_246/A INVX1_LOC_42/A 0.03fF
C4234 NOR2X1_LOC_503/a_36_216# INVX1_LOC_42/A -0.00fF
C4235 NOR2X1_LOC_750/A NAND2X1_LOC_74/B 0.04fF
C4236 NAND2X1_LOC_391/Y INVX1_LOC_61/A 0.02fF
C4237 NAND2X1_LOC_9/Y NOR2X1_LOC_340/Y 0.02fF
C4238 INVX1_LOC_17/A INVX1_LOC_31/A 0.36fF
C4239 INVX1_LOC_279/A INVX1_LOC_4/A 0.07fF
C4240 NAND2X1_LOC_338/B NOR2X1_LOC_39/Y 0.42fF
C4241 NOR2X1_LOC_332/A INVX1_LOC_32/A 0.07fF
C4242 INVX1_LOC_207/Y INVX1_LOC_42/A 0.18fF
C4243 INVX1_LOC_55/Y INVX1_LOC_42/A 4.02fF
C4244 INVX1_LOC_13/A INVX1_LOC_78/A 0.03fF
C4245 INVX1_LOC_35/A NOR2X1_LOC_732/A 0.01fF
C4246 NOR2X1_LOC_389/A INVX1_LOC_174/A 0.42fF
C4247 INVX1_LOC_201/A NOR2X1_LOC_814/A 0.19fF
C4248 INVX1_LOC_54/Y INVX1_LOC_29/Y 0.05fF
C4249 INVX1_LOC_143/A INVX1_LOC_57/A 0.07fF
C4250 NAND2X1_LOC_338/B NAND2X1_LOC_205/A 0.03fF
C4251 INVX1_LOC_278/A NOR2X1_LOC_52/B 0.07fF
C4252 NOR2X1_LOC_175/B NOR2X1_LOC_748/A 0.09fF
C4253 INVX1_LOC_146/A NOR2X1_LOC_48/B 0.15fF
C4254 INVX1_LOC_149/A INVX1_LOC_58/Y 0.02fF
C4255 NOR2X1_LOC_802/A NOR2X1_LOC_634/Y 0.07fF
C4256 INVX1_LOC_35/A INVX1_LOC_124/A 0.33fF
C4257 NOR2X1_LOC_92/Y NAND2X1_LOC_837/Y 0.20fF
C4258 NOR2X1_LOC_479/B INVX1_LOC_166/A 0.05fF
C4259 NOR2X1_LOC_289/a_36_216# INVX1_LOC_271/A 0.01fF
C4260 NOR2X1_LOC_178/Y NOR2X1_LOC_315/Y 0.02fF
C4261 NAND2X1_LOC_9/Y NOR2X1_LOC_655/B 0.05fF
C4262 NOR2X1_LOC_827/a_36_216# INVX1_LOC_64/A 0.01fF
C4263 NOR2X1_LOC_195/A NOR2X1_LOC_554/B 0.01fF
C4264 INVX1_LOC_17/A NAND2X1_LOC_106/a_36_24# 0.00fF
C4265 INVX1_LOC_2/Y NOR2X1_LOC_78/Y 0.51fF
C4266 NOR2X1_LOC_65/B INVX1_LOC_13/A 0.03fF
C4267 NOR2X1_LOC_454/a_36_216# NOR2X1_LOC_454/Y 0.02fF
C4268 NAND2X1_LOC_656/Y NOR2X1_LOC_278/Y 0.02fF
C4269 INVX1_LOC_11/A NOR2X1_LOC_168/Y 0.03fF
C4270 INVX1_LOC_299/A NOR2X1_LOC_274/Y 0.02fF
C4271 NOR2X1_LOC_246/A INVX1_LOC_78/A 0.07fF
C4272 INVX1_LOC_22/A NOR2X1_LOC_748/A 0.06fF
C4273 INVX1_LOC_5/A NAND2X1_LOC_147/a_36_24# 0.00fF
C4274 INVX1_LOC_50/A NOR2X1_LOC_570/Y 0.03fF
C4275 NAND2X1_LOC_472/Y INVX1_LOC_274/A 0.14fF
C4276 NOR2X1_LOC_172/Y NOR2X1_LOC_321/Y 0.03fF
C4277 INVX1_LOC_7/A NAND2X1_LOC_99/A 0.00fF
C4278 NOR2X1_LOC_483/B INVX1_LOC_18/A 0.01fF
C4279 NOR2X1_LOC_356/A NOR2X1_LOC_334/Y 0.07fF
C4280 INVX1_LOC_41/A NOR2X1_LOC_92/Y 0.03fF
C4281 INVX1_LOC_208/Y INVX1_LOC_53/A 0.03fF
C4282 NOR2X1_LOC_15/Y NAND2X1_LOC_640/Y -0.00fF
C4283 INVX1_LOC_55/Y INVX1_LOC_78/A 0.64fF
C4284 NAND2X1_LOC_63/Y INVX1_LOC_91/A 0.03fF
C4285 INVX1_LOC_74/A INVX1_LOC_84/A 0.02fF
C4286 INVX1_LOC_41/A INVX1_LOC_24/Y 3.38fF
C4287 NOR2X1_LOC_19/B INVX1_LOC_253/A 0.01fF
C4288 INVX1_LOC_174/A NOR2X1_LOC_596/A 0.13fF
C4289 NOR2X1_LOC_486/Y INVX1_LOC_186/Y 0.07fF
C4290 INVX1_LOC_21/A NOR2X1_LOC_175/A 0.07fF
C4291 INVX1_LOC_135/A NOR2X1_LOC_383/B 0.03fF
C4292 NOR2X1_LOC_244/B NOR2X1_LOC_240/Y 0.02fF
C4293 INVX1_LOC_35/A NOR2X1_LOC_687/Y 0.03fF
C4294 NOR2X1_LOC_655/B NOR2X1_LOC_798/A 0.01fF
C4295 INVX1_LOC_225/A NOR2X1_LOC_15/Y 0.73fF
C4296 NOR2X1_LOC_845/A NOR2X1_LOC_67/Y 0.02fF
C4297 INVX1_LOC_88/A NAND2X1_LOC_332/Y 0.39fF
C4298 NOR2X1_LOC_160/B INVX1_LOC_184/Y 0.03fF
C4299 NOR2X1_LOC_627/Y INVX1_LOC_27/A 0.02fF
C4300 INVX1_LOC_11/A NAND2X1_LOC_21/Y 0.33fF
C4301 INVX1_LOC_13/A INVX1_LOC_152/Y 0.01fF
C4302 NOR2X1_LOC_130/A INVX1_LOC_57/A 0.06fF
C4303 NAND2X1_LOC_725/B INVX1_LOC_240/A 0.03fF
C4304 NAND2X1_LOC_807/Y NOR2X1_LOC_301/A 0.01fF
C4305 INVX1_LOC_224/Y NOR2X1_LOC_71/Y 0.08fF
C4306 NOR2X1_LOC_92/Y NAND2X1_LOC_477/A 0.13fF
C4307 NOR2X1_LOC_769/B NOR2X1_LOC_763/Y 0.04fF
C4308 NAND2X1_LOC_9/Y NAND2X1_LOC_358/Y 0.01fF
C4309 INVX1_LOC_140/A NAND2X1_LOC_175/Y 0.10fF
C4310 NOR2X1_LOC_67/A NOR2X1_LOC_789/B 0.02fF
C4311 NOR2X1_LOC_280/Y NOR2X1_LOC_662/A 0.01fF
C4312 NOR2X1_LOC_74/A NAND2X1_LOC_444/B 0.02fF
C4313 INVX1_LOC_45/A INVX1_LOC_45/Y 1.01fF
C4314 NAND2X1_LOC_564/B NAND2X1_LOC_552/A -0.00fF
C4315 NOR2X1_LOC_523/A NOR2X1_LOC_844/A 0.37fF
C4316 INVX1_LOC_22/A NOR2X1_LOC_304/Y 0.20fF
C4317 INVX1_LOC_272/Y NAND2X1_LOC_799/Y 0.10fF
C4318 NOR2X1_LOC_74/A NOR2X1_LOC_334/Y 0.18fF
C4319 NOR2X1_LOC_598/B NOR2X1_LOC_763/Y 0.89fF
C4320 INVX1_LOC_269/A NOR2X1_LOC_399/A 0.00fF
C4321 NOR2X1_LOC_477/a_36_216# INVX1_LOC_113/Y 0.00fF
C4322 NOR2X1_LOC_793/A INVX1_LOC_177/A 0.01fF
C4323 INVX1_LOC_64/A INVX1_LOC_279/A 0.37fF
C4324 NAND2X1_LOC_9/Y NOR2X1_LOC_99/B 0.03fF
C4325 INVX1_LOC_11/A INVX1_LOC_76/Y 0.09fF
C4326 INVX1_LOC_33/Y NOR2X1_LOC_653/Y 0.07fF
C4327 NOR2X1_LOC_320/Y INVX1_LOC_78/A 0.01fF
C4328 INVX1_LOC_251/Y INVX1_LOC_14/A 1.45fF
C4329 INVX1_LOC_133/A NAND2X1_LOC_211/Y 0.03fF
C4330 INVX1_LOC_6/A NOR2X1_LOC_158/B 0.00fF
C4331 INVX1_LOC_91/A INVX1_LOC_257/A 0.01fF
C4332 INVX1_LOC_224/A NOR2X1_LOC_16/Y 0.01fF
C4333 NAND2X1_LOC_198/B NOR2X1_LOC_338/Y 0.05fF
C4334 NAND2X1_LOC_573/Y NAND2X1_LOC_840/B 0.00fF
C4335 NOR2X1_LOC_647/A NAND2X1_LOC_348/A 0.02fF
C4336 NAND2X1_LOC_740/A NAND2X1_LOC_856/A 0.07fF
C4337 NAND2X1_LOC_569/B D_INPUT_0 0.07fF
C4338 NOR2X1_LOC_440/Y NOR2X1_LOC_652/Y 0.34fF
C4339 INVX1_LOC_223/A NOR2X1_LOC_550/B 0.00fF
C4340 INVX1_LOC_17/A INVX1_LOC_191/Y 0.03fF
C4341 VDD NAND2X1_LOC_207/B 0.36fF
C4342 NAND2X1_LOC_59/B NAND2X1_LOC_36/A 0.18fF
C4343 INVX1_LOC_33/A NOR2X1_LOC_532/a_36_216# 0.00fF
C4344 NOR2X1_LOC_179/Y INVX1_LOC_118/A 0.07fF
C4345 INVX1_LOC_33/Y INVX1_LOC_19/A 0.04fF
C4346 NOR2X1_LOC_171/Y INVX1_LOC_23/A 0.03fF
C4347 NAND2X1_LOC_583/a_36_24# NAND2X1_LOC_451/Y 0.00fF
C4348 NOR2X1_LOC_238/Y INVX1_LOC_41/Y 0.00fF
C4349 NOR2X1_LOC_601/Y INVX1_LOC_15/A 0.03fF
C4350 NOR2X1_LOC_160/B INVX1_LOC_177/A 2.04fF
C4351 INVX1_LOC_45/Y INVX1_LOC_71/A 0.01fF
C4352 INVX1_LOC_125/Y NAND2X1_LOC_447/a_36_24# 0.00fF
C4353 INVX1_LOC_119/Y INVX1_LOC_54/A 0.07fF
C4354 INVX1_LOC_33/A INVX1_LOC_18/A 0.16fF
C4355 INVX1_LOC_280/Y NAND2X1_LOC_550/A 0.03fF
C4356 GATE_741 NOR2X1_LOC_299/Y 0.14fF
C4357 INVX1_LOC_203/A INVX1_LOC_118/A 0.07fF
C4358 NAND2X1_LOC_798/B NOR2X1_LOC_841/A 0.10fF
C4359 INVX1_LOC_174/A INVX1_LOC_189/Y 0.02fF
C4360 NOR2X1_LOC_711/A NOR2X1_LOC_383/B 0.16fF
C4361 NOR2X1_LOC_465/a_36_216# INVX1_LOC_182/Y 0.00fF
C4362 NAND2X1_LOC_733/Y NOR2X1_LOC_822/Y 0.02fF
C4363 INVX1_LOC_75/A NOR2X1_LOC_392/Y 0.07fF
C4364 INVX1_LOC_64/A INVX1_LOC_182/Y 0.00fF
C4365 INVX1_LOC_37/A NOR2X1_LOC_452/a_36_216# 0.00fF
C4366 INVX1_LOC_20/A NOR2X1_LOC_38/B 0.03fF
C4367 NOR2X1_LOC_794/A NOR2X1_LOC_383/B 0.01fF
C4368 NOR2X1_LOC_791/a_36_216# INVX1_LOC_8/A 0.01fF
C4369 INVX1_LOC_150/Y INVX1_LOC_1/Y 0.13fF
C4370 D_INPUT_1 INVX1_LOC_69/Y 0.03fF
C4371 D_INPUT_0 NOR2X1_LOC_140/A 0.01fF
C4372 NOR2X1_LOC_250/A NAND2X1_LOC_660/Y 0.36fF
C4373 INVX1_LOC_291/A INVX1_LOC_264/A 0.06fF
C4374 INVX1_LOC_163/A NAND2X1_LOC_624/A 0.03fF
C4375 INVX1_LOC_94/A INVX1_LOC_104/A 0.07fF
C4376 NOR2X1_LOC_82/A INVX1_LOC_80/A 0.01fF
C4377 NOR2X1_LOC_790/B NOR2X1_LOC_551/Y 0.06fF
C4378 D_INPUT_0 NAND2X1_LOC_538/Y 0.17fF
C4379 NAND2X1_LOC_35/Y NOR2X1_LOC_394/a_36_216# 0.00fF
C4380 NAND2X1_LOC_711/Y INVX1_LOC_22/A 0.00fF
C4381 NOR2X1_LOC_357/Y INVX1_LOC_78/A 0.03fF
C4382 NOR2X1_LOC_389/A NOR2X1_LOC_589/A 0.08fF
C4383 INVX1_LOC_159/A NAND2X1_LOC_661/B 0.02fF
C4384 NOR2X1_LOC_243/Y NOR2X1_LOC_860/B 0.28fF
C4385 INVX1_LOC_223/Y INVX1_LOC_75/A 0.91fF
C4386 D_INPUT_0 NOR2X1_LOC_250/A 0.03fF
C4387 NOR2X1_LOC_103/Y NOR2X1_LOC_71/Y 1.19fF
C4388 INVX1_LOC_17/A INVX1_LOC_313/A 0.09fF
C4389 NOR2X1_LOC_160/B NOR2X1_LOC_785/Y 0.05fF
C4390 NAND2X1_LOC_357/B NOR2X1_LOC_753/Y 0.07fF
C4391 INVX1_LOC_235/A INVX1_LOC_75/A 0.03fF
C4392 NOR2X1_LOC_589/A NAND2X1_LOC_199/B 0.04fF
C4393 INVX1_LOC_251/Y NAND2X1_LOC_84/Y 0.10fF
C4394 NOR2X1_LOC_673/A INVX1_LOC_63/A 0.03fF
C4395 INVX1_LOC_85/A NOR2X1_LOC_550/B 0.07fF
C4396 NOR2X1_LOC_607/A NAND2X1_LOC_294/a_36_24# 0.00fF
C4397 INVX1_LOC_34/A NAND2X1_LOC_139/A 0.01fF
C4398 INVX1_LOC_76/A NAND2X1_LOC_99/A 0.07fF
C4399 INVX1_LOC_119/A NOR2X1_LOC_577/Y 0.10fF
C4400 D_INPUT_0 NOR2X1_LOC_530/Y 0.01fF
C4401 INPUT_3 NOR2X1_LOC_332/A 0.41fF
C4402 INVX1_LOC_236/A NOR2X1_LOC_152/Y 0.40fF
C4403 NOR2X1_LOC_716/B NOR2X1_LOC_369/a_36_216# 0.01fF
C4404 NOR2X1_LOC_537/A INVX1_LOC_149/A 0.08fF
C4405 INVX1_LOC_90/A NAND2X1_LOC_793/Y 0.00fF
C4406 NAND2X1_LOC_357/B NAND2X1_LOC_325/Y 0.02fF
C4407 INVX1_LOC_255/Y NOR2X1_LOC_819/a_36_216# 0.00fF
C4408 INVX1_LOC_72/Y INVX1_LOC_232/A 0.02fF
C4409 NOR2X1_LOC_493/B NOR2X1_LOC_577/Y 0.02fF
C4410 INVX1_LOC_41/A NAND2X1_LOC_477/A 0.03fF
C4411 INVX1_LOC_17/A NAND2X1_LOC_807/Y 0.07fF
C4412 NOR2X1_LOC_757/A INVX1_LOC_30/A 0.08fF
C4413 NOR2X1_LOC_437/a_36_216# NOR2X1_LOC_757/Y 0.00fF
C4414 INVX1_LOC_58/A NAND2X1_LOC_465/A 0.53fF
C4415 INVX1_LOC_285/A INVX1_LOC_29/A 0.32fF
C4416 INVX1_LOC_49/A NOR2X1_LOC_352/Y 0.04fF
C4417 NOR2X1_LOC_722/a_36_216# INVX1_LOC_266/Y 0.01fF
C4418 NOR2X1_LOC_88/Y NAND2X1_LOC_254/Y 0.03fF
C4419 NAND2X1_LOC_149/Y NOR2X1_LOC_589/Y 0.14fF
C4420 INVX1_LOC_33/A INVX1_LOC_34/Y 0.07fF
C4421 NAND2X1_LOC_833/Y NOR2X1_LOC_482/Y 0.00fF
C4422 NOR2X1_LOC_280/Y INVX1_LOC_57/A 0.02fF
C4423 NOR2X1_LOC_691/B NOR2X1_LOC_691/a_36_216# 0.02fF
C4424 NOR2X1_LOC_589/A INVX1_LOC_107/A 0.06fF
C4425 NOR2X1_LOC_446/a_36_216# INVX1_LOC_313/Y 0.00fF
C4426 INVX1_LOC_139/Y NOR2X1_LOC_383/B 0.03fF
C4427 INVX1_LOC_85/A INVX1_LOC_249/Y 0.01fF
C4428 INVX1_LOC_29/A NOR2X1_LOC_814/A 0.32fF
C4429 NAND2X1_LOC_736/Y INVX1_LOC_282/Y 0.13fF
C4430 INVX1_LOC_45/A NOR2X1_LOC_71/Y 0.08fF
C4431 INVX1_LOC_57/Y INVX1_LOC_135/A 0.10fF
C4432 INVX1_LOC_279/A INVX1_LOC_130/Y 0.00fF
C4433 NOR2X1_LOC_78/B NOR2X1_LOC_551/B 0.01fF
C4434 NOR2X1_LOC_599/A NAND2X1_LOC_801/a_36_24# 0.00fF
C4435 NOR2X1_LOC_589/A NOR2X1_LOC_596/A 0.64fF
C4436 NOR2X1_LOC_536/A NOR2X1_LOC_318/A 1.22fF
C4437 INVX1_LOC_30/Y NOR2X1_LOC_81/a_36_216# 0.00fF
C4438 NOR2X1_LOC_615/Y NAND2X1_LOC_560/A 0.01fF
C4439 NAND2X1_LOC_562/Y NAND2X1_LOC_578/B 0.21fF
C4440 INVX1_LOC_1/A INVX1_LOC_92/Y 0.12fF
C4441 NOR2X1_LOC_65/B INVX1_LOC_66/Y 0.01fF
C4442 INVX1_LOC_84/A NAND2X1_LOC_254/Y 0.03fF
C4443 NOR2X1_LOC_726/Y NOR2X1_LOC_724/Y 0.01fF
C4444 NOR2X1_LOC_706/B INVX1_LOC_23/A 0.01fF
C4445 NOR2X1_LOC_48/B INVX1_LOC_119/Y 0.15fF
C4446 INVX1_LOC_7/A NAND2X1_LOC_656/A 0.03fF
C4447 INVX1_LOC_36/A INVX1_LOC_20/Y 0.01fF
C4448 NOR2X1_LOC_709/B INVX1_LOC_26/A 0.01fF
C4449 NAND2X1_LOC_787/A INVX1_LOC_37/A 0.03fF
C4450 INVX1_LOC_45/A NOR2X1_LOC_644/A 0.03fF
C4451 INVX1_LOC_58/A INVX1_LOC_77/Y 0.04fF
C4452 INVX1_LOC_251/Y NOR2X1_LOC_612/B 0.05fF
C4453 NOR2X1_LOC_480/A INVX1_LOC_135/A 0.03fF
C4454 NOR2X1_LOC_372/Y INPUT_1 0.30fF
C4455 INVX1_LOC_42/A NAND2X1_LOC_489/Y 0.04fF
C4456 INVX1_LOC_27/A NOR2X1_LOC_405/A 0.07fF
C4457 NOR2X1_LOC_220/B NAND2X1_LOC_447/Y 0.02fF
C4458 NAND2X1_LOC_363/B INVX1_LOC_37/A 0.60fF
C4459 INVX1_LOC_17/A INVX1_LOC_6/A 0.10fF
C4460 NOR2X1_LOC_299/Y NAND2X1_LOC_837/Y 0.01fF
C4461 INVX1_LOC_45/A NOR2X1_LOC_828/B 0.03fF
C4462 INVX1_LOC_136/A NOR2X1_LOC_750/A 0.05fF
C4463 INVX1_LOC_2/A NAND2X1_LOC_374/Y 0.07fF
C4464 INVX1_LOC_1/A NOR2X1_LOC_562/B 0.10fF
C4465 INVX1_LOC_11/A NOR2X1_LOC_548/a_36_216# 0.00fF
C4466 INVX1_LOC_93/A INVX1_LOC_126/A 0.05fF
C4467 INVX1_LOC_233/A NOR2X1_LOC_176/Y 0.01fF
C4468 NOR2X1_LOC_637/A INVX1_LOC_90/A 0.02fF
C4469 INVX1_LOC_14/A NOR2X1_LOC_45/B 6.76fF
C4470 NAND2X1_LOC_364/A NOR2X1_LOC_772/A 0.01fF
C4471 NOR2X1_LOC_716/B INVX1_LOC_164/A 0.21fF
C4472 INVX1_LOC_102/A NAND2X1_LOC_74/B 0.07fF
C4473 NAND2X1_LOC_218/B INVX1_LOC_89/A 0.14fF
C4474 INVX1_LOC_57/A NOR2X1_LOC_16/a_36_216# 0.00fF
C4475 INVX1_LOC_33/A NOR2X1_LOC_383/a_36_216# 0.00fF
C4476 INVX1_LOC_208/A INVX1_LOC_177/A 0.03fF
C4477 NOR2X1_LOC_15/Y NAND2X1_LOC_642/Y 0.11fF
C4478 INVX1_LOC_40/A INVX1_LOC_34/Y 0.29fF
C4479 NOR2X1_LOC_197/A INVX1_LOC_78/Y 0.00fF
C4480 INVX1_LOC_103/A NOR2X1_LOC_139/Y 0.00fF
C4481 NOR2X1_LOC_516/B INVX1_LOC_177/A 0.03fF
C4482 NAND2X1_LOC_578/a_36_24# NAND2X1_LOC_659/B 0.00fF
C4483 NOR2X1_LOC_644/A INVX1_LOC_71/A 0.03fF
C4484 NOR2X1_LOC_215/A NOR2X1_LOC_357/Y 0.05fF
C4485 INVX1_LOC_203/A NAND2X1_LOC_618/Y 0.10fF
C4486 INVX1_LOC_28/A NAND2X1_LOC_306/a_36_24# 0.00fF
C4487 NAND2X1_LOC_67/Y NOR2X1_LOC_69/A 0.03fF
C4488 NOR2X1_LOC_78/B INVX1_LOC_208/Y 0.03fF
C4489 INVX1_LOC_35/A INVX1_LOC_9/A 0.06fF
C4490 NOR2X1_LOC_604/Y INVX1_LOC_54/A 0.01fF
C4491 INVX1_LOC_2/Y NAND2X1_LOC_473/A 0.04fF
C4492 NOR2X1_LOC_41/Y NAND2X1_LOC_662/Y 0.04fF
C4493 INVX1_LOC_13/A NOR2X1_LOC_721/A 0.01fF
C4494 INVX1_LOC_55/Y INVX1_LOC_113/Y 0.03fF
C4495 INVX1_LOC_103/A NAND2X1_LOC_468/B 0.00fF
C4496 NOR2X1_LOC_858/A INVX1_LOC_307/A 0.03fF
C4497 NOR2X1_LOC_281/Y INVX1_LOC_285/A 0.04fF
C4498 NOR2X1_LOC_468/Y INVX1_LOC_20/A 0.10fF
C4499 INVX1_LOC_78/A NAND2X1_LOC_489/Y 0.01fF
C4500 NAND2X1_LOC_656/B INVX1_LOC_29/Y 0.03fF
C4501 NAND2X1_LOC_787/A NOR2X1_LOC_177/Y 0.01fF
C4502 NAND2X1_LOC_223/B NOR2X1_LOC_673/A 0.14fF
C4503 INVX1_LOC_298/A INVX1_LOC_38/A 0.01fF
C4504 NOR2X1_LOC_794/a_36_216# NOR2X1_LOC_564/Y 0.00fF
C4505 INVX1_LOC_298/Y NOR2X1_LOC_814/A 0.02fF
C4506 NAND2X1_LOC_361/a_36_24# INVX1_LOC_89/A 0.00fF
C4507 NAND2X1_LOC_579/A INVX1_LOC_46/A 0.11fF
C4508 NOR2X1_LOC_570/B INVX1_LOC_313/Y 0.07fF
C4509 NOR2X1_LOC_160/B INVX1_LOC_65/A 0.01fF
C4510 INVX1_LOC_286/A INVX1_LOC_72/A 0.10fF
C4511 NOR2X1_LOC_33/Y NOR2X1_LOC_814/A -0.03fF
C4512 INVX1_LOC_179/Y INVX1_LOC_220/Y 0.08fF
C4513 NAND2X1_LOC_93/B NOR2X1_LOC_678/A 0.03fF
C4514 NAND2X1_LOC_254/Y INVX1_LOC_15/A 0.03fF
C4515 NOR2X1_LOC_361/B NAND2X1_LOC_211/Y 0.11fF
C4516 INVX1_LOC_32/A INVX1_LOC_42/A 0.49fF
C4517 NAND2X1_LOC_149/Y INVX1_LOC_117/A 4.43fF
C4518 NOR2X1_LOC_142/Y NAND2X1_LOC_842/B 0.03fF
C4519 NAND2X1_LOC_93/B INVX1_LOC_295/Y 0.11fF
C4520 NOR2X1_LOC_639/B INVX1_LOC_92/A 0.02fF
C4521 NOR2X1_LOC_757/a_36_216# NAND2X1_LOC_656/Y 0.01fF
C4522 D_INPUT_6 INVX1_LOC_38/A 0.03fF
C4523 NOR2X1_LOC_84/Y NOR2X1_LOC_76/A 0.48fF
C4524 INVX1_LOC_193/Y NOR2X1_LOC_546/B 0.00fF
C4525 INVX1_LOC_77/A NOR2X1_LOC_534/a_36_216# 0.00fF
C4526 NAND2X1_LOC_726/Y NOR2X1_LOC_690/Y 0.01fF
C4527 NOR2X1_LOC_173/Y INVX1_LOC_38/A 0.04fF
C4528 INVX1_LOC_23/Y INVX1_LOC_19/A 0.07fF
C4529 INVX1_LOC_54/A NOR2X1_LOC_674/Y 0.61fF
C4530 NOR2X1_LOC_500/A NOR2X1_LOC_552/Y 0.03fF
C4531 INVX1_LOC_23/A NOR2X1_LOC_430/Y 0.05fF
C4532 NAND2X1_LOC_425/Y INVX1_LOC_295/Y 0.04fF
C4533 NOR2X1_LOC_320/Y NOR2X1_LOC_152/Y 0.05fF
C4534 NOR2X1_LOC_760/a_36_216# NOR2X1_LOC_137/Y 0.00fF
C4535 NOR2X1_LOC_457/A INVX1_LOC_37/A 0.01fF
C4536 NOR2X1_LOC_321/Y INVX1_LOC_38/A 0.09fF
C4537 INVX1_LOC_94/A INVX1_LOC_206/Y 0.00fF
C4538 NOR2X1_LOC_781/A INVX1_LOC_290/A 0.02fF
C4539 INVX1_LOC_1/A INVX1_LOC_281/Y 0.01fF
C4540 INVX1_LOC_229/Y NAND2X1_LOC_863/B 0.07fF
C4541 NOR2X1_LOC_220/A INVX1_LOC_171/A 0.43fF
C4542 INVX1_LOC_186/Y NOR2X1_LOC_748/A 0.08fF
C4543 NOR2X1_LOC_791/Y NOR2X1_LOC_743/Y 0.00fF
C4544 NOR2X1_LOC_843/a_36_216# NOR2X1_LOC_814/A 0.01fF
C4545 NAND2X1_LOC_374/Y INPUT_1 0.19fF
C4546 NOR2X1_LOC_15/Y NOR2X1_LOC_271/Y 0.02fF
C4547 NAND2X1_LOC_175/Y INVX1_LOC_42/A 0.03fF
C4548 D_INPUT_6 NOR2X1_LOC_51/A 0.03fF
C4549 NAND2X1_LOC_538/Y NAND2X1_LOC_848/A 0.10fF
C4550 NAND2X1_LOC_537/Y NAND2X1_LOC_846/a_36_24# 0.00fF
C4551 INVX1_LOC_33/A NOR2X1_LOC_548/A 0.01fF
C4552 INVX1_LOC_53/A NOR2X1_LOC_691/A 0.07fF
C4553 NOR2X1_LOC_816/A NAND2X1_LOC_804/Y 0.02fF
C4554 NAND2X1_LOC_579/a_36_24# NOR2X1_LOC_299/Y 0.00fF
C4555 NAND2X1_LOC_139/A INPUT_0 0.02fF
C4556 NOR2X1_LOC_264/Y NOR2X1_LOC_721/Y 0.01fF
C4557 NOR2X1_LOC_38/B INVX1_LOC_4/A 0.03fF
C4558 INVX1_LOC_195/A NAND2X1_LOC_659/B 0.00fF
C4559 INVX1_LOC_18/A NOR2X1_LOC_486/Y 0.03fF
C4560 INVX1_LOC_311/A INVX1_LOC_63/Y 0.22fF
C4561 INVX1_LOC_176/A NOR2X1_LOC_500/B 0.02fF
C4562 NOR2X1_LOC_78/B NOR2X1_LOC_756/Y 0.05fF
C4563 NAND2X1_LOC_319/A INVX1_LOC_10/A 0.01fF
C4564 INVX1_LOC_89/A INVX1_LOC_22/A 0.22fF
C4565 NAND2X1_LOC_40/a_36_24# INVX1_LOC_29/A 0.02fF
C4566 INVX1_LOC_78/A INVX1_LOC_32/A 0.16fF
C4567 NOR2X1_LOC_354/B INVX1_LOC_143/Y 0.01fF
C4568 INVX1_LOC_210/Y VDD 0.27fF
C4569 NOR2X1_LOC_283/a_36_216# NOR2X1_LOC_78/A 0.00fF
C4570 NOR2X1_LOC_190/a_36_216# INVX1_LOC_102/Y 0.00fF
C4571 INVX1_LOC_30/A INVX1_LOC_37/A 0.22fF
C4572 INVX1_LOC_243/A D_INPUT_4 0.01fF
C4573 NOR2X1_LOC_592/A INVX1_LOC_118/A 0.00fF
C4574 INVX1_LOC_30/A NOR2X1_LOC_231/A 0.01fF
C4575 NOR2X1_LOC_67/A NAND2X1_LOC_849/A 0.09fF
C4576 INVX1_LOC_195/A VDD 0.00fF
C4577 INVX1_LOC_284/A NAND2X1_LOC_215/A 0.18fF
C4578 D_INPUT_1 NOR2X1_LOC_89/A 1.59fF
C4579 NAND2X1_LOC_763/B INVX1_LOC_37/A 0.00fF
C4580 INVX1_LOC_67/A NOR2X1_LOC_139/Y 0.01fF
C4581 INVX1_LOC_312/A INVX1_LOC_33/Y 0.24fF
C4582 NAND2X1_LOC_656/A INVX1_LOC_76/A 0.10fF
C4583 INVX1_LOC_34/A NOR2X1_LOC_78/A 0.04fF
C4584 NOR2X1_LOC_65/B INVX1_LOC_32/A 0.03fF
C4585 D_INPUT_0 NOR2X1_LOC_106/A 0.27fF
C4586 NOR2X1_LOC_123/B NOR2X1_LOC_71/Y 0.01fF
C4587 NOR2X1_LOC_637/B NOR2X1_LOC_56/Y 0.01fF
C4588 NOR2X1_LOC_82/A NOR2X1_LOC_99/Y 0.01fF
C4589 INVX1_LOC_306/Y NAND2X1_LOC_773/B 0.17fF
C4590 NAND2X1_LOC_564/B INVX1_LOC_140/A -0.01fF
C4591 INVX1_LOC_75/A INVX1_LOC_25/Y 0.03fF
C4592 INVX1_LOC_78/A NAND2X1_LOC_175/Y 0.09fF
C4593 NOR2X1_LOC_456/Y INVX1_LOC_290/Y 0.02fF
C4594 NAND2X1_LOC_858/B NAND2X1_LOC_850/Y 0.18fF
C4595 NOR2X1_LOC_484/Y INVX1_LOC_76/A 0.04fF
C4596 NOR2X1_LOC_19/B NOR2X1_LOC_86/A 0.03fF
C4597 NOR2X1_LOC_220/A INVX1_LOC_222/A 0.03fF
C4598 NAND2X1_LOC_727/Y NAND2X1_LOC_863/A 0.04fF
C4599 INVX1_LOC_18/A NOR2X1_LOC_816/Y 0.01fF
C4600 NOR2X1_LOC_561/Y NOR2X1_LOC_329/B 0.07fF
C4601 NAND2X1_LOC_785/A NOR2X1_LOC_528/Y 0.10fF
C4602 INVX1_LOC_197/Y NAND2X1_LOC_622/B 0.21fF
C4603 INVX1_LOC_75/A NOR2X1_LOC_302/B 0.02fF
C4604 NOR2X1_LOC_186/Y INVX1_LOC_49/Y 0.00fF
C4605 NOR2X1_LOC_91/A INVX1_LOC_94/Y 0.06fF
C4606 INVX1_LOC_35/A NOR2X1_LOC_861/Y 1.44fF
C4607 INVX1_LOC_208/A INVX1_LOC_285/Y 0.10fF
C4608 INVX1_LOC_8/Y VDD 0.21fF
C4609 INVX1_LOC_17/A NOR2X1_LOC_117/Y 0.00fF
C4610 NOR2X1_LOC_637/B VDD 0.14fF
C4611 NOR2X1_LOC_569/Y NOR2X1_LOC_74/A 0.01fF
C4612 NOR2X1_LOC_372/Y INVX1_LOC_118/A 0.01fF
C4613 INVX1_LOC_13/A INVX1_LOC_158/Y 0.06fF
C4614 NOR2X1_LOC_89/A NOR2X1_LOC_652/Y 0.35fF
C4615 NOR2X1_LOC_590/A NOR2X1_LOC_634/A 0.02fF
C4616 NAND2X1_LOC_837/Y NOR2X1_LOC_494/a_36_216# 0.01fF
C4617 INVX1_LOC_155/A VDD 0.15fF
C4618 INVX1_LOC_72/A INVX1_LOC_54/A 0.46fF
C4619 NOR2X1_LOC_218/a_36_216# NAND2X1_LOC_656/Y 0.01fF
C4620 NOR2X1_LOC_168/A NOR2X1_LOC_552/A 0.02fF
C4621 INVX1_LOC_50/A NOR2X1_LOC_36/A -0.01fF
C4622 NOR2X1_LOC_134/Y NOR2X1_LOC_103/a_36_216# 0.00fF
C4623 INVX1_LOC_30/A NOR2X1_LOC_743/Y 0.03fF
C4624 INVX1_LOC_45/Y NOR2X1_LOC_331/B 0.02fF
C4625 INVX1_LOC_23/A INVX1_LOC_94/Y 0.80fF
C4626 NOR2X1_LOC_186/Y NAND2X1_LOC_288/a_36_24# 0.00fF
C4627 NOR2X1_LOC_788/B NOR2X1_LOC_564/Y 0.00fF
C4628 NAND2X1_LOC_569/A VDD 0.27fF
C4629 INVX1_LOC_27/A INVX1_LOC_109/Y 0.07fF
C4630 INVX1_LOC_295/A NOR2X1_LOC_163/Y 0.03fF
C4631 NOR2X1_LOC_264/Y VDD 0.87fF
C4632 INVX1_LOC_232/A INVX1_LOC_125/Y 0.10fF
C4633 NOR2X1_LOC_836/Y NOR2X1_LOC_865/Y 0.03fF
C4634 NOR2X1_LOC_91/A INVX1_LOC_181/A 0.00fF
C4635 NOR2X1_LOC_381/Y NAND2X1_LOC_82/Y 0.26fF
C4636 INVX1_LOC_64/A NOR2X1_LOC_38/B 0.11fF
C4637 INVX1_LOC_224/Y INVX1_LOC_16/Y 0.01fF
C4638 NOR2X1_LOC_423/Y INVX1_LOC_76/A 0.01fF
C4639 NAND2X1_LOC_493/Y INVX1_LOC_12/A 0.03fF
C4640 INVX1_LOC_35/A INVX1_LOC_274/Y 0.12fF
C4641 NOR2X1_LOC_589/A INVX1_LOC_100/Y 0.02fF
C4642 NOR2X1_LOC_707/A NOR2X1_LOC_712/B 0.14fF
C4643 NOR2X1_LOC_751/A NOR2X1_LOC_749/Y 0.12fF
C4644 INVX1_LOC_224/Y NOR2X1_LOC_39/Y 0.04fF
C4645 NAND2X1_LOC_623/B INVX1_LOC_16/A 0.08fF
C4646 NOR2X1_LOC_709/A NOR2X1_LOC_266/B 0.21fF
C4647 NAND2X1_LOC_735/B INVX1_LOC_91/A 0.00fF
C4648 INVX1_LOC_177/Y NOR2X1_LOC_155/A 0.03fF
C4649 NOR2X1_LOC_590/A NOR2X1_LOC_673/B 0.05fF
C4650 NOR2X1_LOC_92/Y INVX1_LOC_168/Y 0.07fF
C4651 INVX1_LOC_24/A NAND2X1_LOC_241/a_36_24# 0.00fF
C4652 NOR2X1_LOC_516/B INVX1_LOC_65/A 0.07fF
C4653 NOR2X1_LOC_420/Y INVX1_LOC_4/A 0.03fF
C4654 NAND2X1_LOC_364/A NOR2X1_LOC_216/B 0.03fF
C4655 NOR2X1_LOC_516/B INVX1_LOC_316/A 0.00fF
C4656 NOR2X1_LOC_773/Y NOR2X1_LOC_279/Y 0.03fF
C4657 NAND2X1_LOC_13/a_36_24# NAND2X1_LOC_74/B 0.06fF
C4658 INVX1_LOC_230/Y NAND2X1_LOC_219/B 0.02fF
C4659 VDD NAND2X1_LOC_661/B 0.01fF
C4660 NOR2X1_LOC_222/Y INVX1_LOC_76/A 0.09fF
C4661 NAND2X1_LOC_721/B INVX1_LOC_285/A 0.01fF
C4662 NOR2X1_LOC_131/Y NAND2X1_LOC_469/B 0.04fF
C4663 INVX1_LOC_224/Y NAND2X1_LOC_205/A 0.10fF
C4664 INVX1_LOC_23/A INVX1_LOC_296/A 0.07fF
C4665 INVX1_LOC_147/A NAND2X1_LOC_652/Y 0.07fF
C4666 NOR2X1_LOC_791/B NOR2X1_LOC_49/a_36_216# 0.00fF
C4667 NAND2X1_LOC_735/B INVX1_LOC_11/Y 0.03fF
C4668 INVX1_LOC_286/Y NOR2X1_LOC_662/A 0.28fF
C4669 NOR2X1_LOC_301/A NOR2X1_LOC_109/Y 0.18fF
C4670 NOR2X1_LOC_68/A NAND2X1_LOC_235/a_36_24# 0.01fF
C4671 NOR2X1_LOC_561/Y INPUT_4 0.00fF
C4672 NOR2X1_LOC_816/A NOR2X1_LOC_519/a_36_216# 0.00fF
C4673 NAND2X1_LOC_863/B INVX1_LOC_20/A 0.02fF
C4674 NOR2X1_LOC_269/a_36_216# INVX1_LOC_76/A 0.00fF
C4675 INVX1_LOC_225/A NAND2X1_LOC_204/a_36_24# 0.00fF
C4676 NOR2X1_LOC_296/Y INVX1_LOC_42/A 0.01fF
C4677 NOR2X1_LOC_148/B NOR2X1_LOC_78/A 0.01fF
C4678 NOR2X1_LOC_457/a_36_216# INVX1_LOC_4/A 0.02fF
C4679 NOR2X1_LOC_589/A NAND2X1_LOC_469/B 0.05fF
C4680 NOR2X1_LOC_590/A INVX1_LOC_29/A 8.49fF
C4681 NOR2X1_LOC_178/Y NAND2X1_LOC_99/A 0.28fF
C4682 NOR2X1_LOC_529/a_36_216# NOR2X1_LOC_392/Y 0.00fF
C4683 VDD INVX1_LOC_316/Y 0.84fF
C4684 INVX1_LOC_208/Y INVX1_LOC_46/A 0.00fF
C4685 NOR2X1_LOC_773/Y NAND2X1_LOC_804/Y 0.01fF
C4686 NOR2X1_LOC_229/Y VDD 0.24fF
C4687 NOR2X1_LOC_52/a_36_216# INVX1_LOC_22/A 0.01fF
C4688 INVX1_LOC_22/Y INVX1_LOC_29/A 0.09fF
C4689 NOR2X1_LOC_468/Y INVX1_LOC_4/A 0.07fF
C4690 INPUT_3 NOR2X1_LOC_847/A 0.04fF
C4691 NOR2X1_LOC_172/Y NAND2X1_LOC_798/B 0.05fF
C4692 NAND2X1_LOC_789/a_36_24# INVX1_LOC_63/A 0.01fF
C4693 INVX1_LOC_155/Y INVX1_LOC_92/A 0.02fF
C4694 NAND2X1_LOC_190/Y INVX1_LOC_4/A 0.04fF
C4695 NAND2X1_LOC_741/B NOR2X1_LOC_11/Y 0.03fF
C4696 INPUT_3 INVX1_LOC_42/A 0.00fF
C4697 NAND2X1_LOC_737/a_36_24# NOR2X1_LOC_36/B 0.00fF
C4698 NOR2X1_LOC_332/A NOR2X1_LOC_332/B 0.02fF
C4699 NOR2X1_LOC_752/a_36_216# INVX1_LOC_77/Y 0.01fF
C4700 INVX1_LOC_314/Y INVX1_LOC_84/A 0.07fF
C4701 INVX1_LOC_160/Y VDD 0.56fF
C4702 INVX1_LOC_16/A INVX1_LOC_117/A 0.02fF
C4703 NAND2X1_LOC_863/B NOR2X1_LOC_765/Y 0.05fF
C4704 NOR2X1_LOC_278/A INVX1_LOC_70/A 0.18fF
C4705 INVX1_LOC_33/A NAND2X1_LOC_210/a_36_24# 0.01fF
C4706 NOR2X1_LOC_65/B INVX1_LOC_171/Y 0.26fF
C4707 NOR2X1_LOC_594/Y INVX1_LOC_6/A 0.28fF
C4708 NOR2X1_LOC_772/A NOR2X1_LOC_405/A 0.01fF
C4709 NAND2X1_LOC_374/Y INVX1_LOC_118/A 0.27fF
C4710 INVX1_LOC_92/Y NOR2X1_LOC_188/A 0.02fF
C4711 INVX1_LOC_104/A NOR2X1_LOC_155/A 0.09fF
C4712 INVX1_LOC_131/A NOR2X1_LOC_78/A 0.08fF
C4713 INVX1_LOC_236/A INVX1_LOC_291/A 0.12fF
C4714 NOR2X1_LOC_160/B NAND2X1_LOC_269/a_36_24# 0.00fF
C4715 INVX1_LOC_136/A INVX1_LOC_102/A 0.07fF
C4716 INVX1_LOC_201/Y NAND2X1_LOC_574/A 0.05fF
C4717 NOR2X1_LOC_709/A INVX1_LOC_46/Y 0.30fF
C4718 NOR2X1_LOC_168/B NOR2X1_LOC_809/B 0.16fF
C4719 NOR2X1_LOC_355/B NOR2X1_LOC_188/A 0.08fF
C4720 NOR2X1_LOC_457/A NAND2X1_LOC_72/B 0.03fF
C4721 INPUT_0 INVX1_LOC_98/A 0.12fF
C4722 NOR2X1_LOC_121/A INVX1_LOC_9/A 0.11fF
C4723 INVX1_LOC_72/A NOR2X1_LOC_48/B 2.59fF
C4724 NOR2X1_LOC_160/B INVX1_LOC_4/Y 0.26fF
C4725 INPUT_0 NOR2X1_LOC_78/A 0.39fF
C4726 INVX1_LOC_8/A NOR2X1_LOC_814/A 0.01fF
C4727 INVX1_LOC_1/A NOR2X1_LOC_699/a_36_216# 0.00fF
C4728 NAND2X1_LOC_562/Y INVX1_LOC_203/A 0.14fF
C4729 NOR2X1_LOC_329/B INVX1_LOC_76/A 0.27fF
C4730 INVX1_LOC_1/Y NOR2X1_LOC_612/Y 0.01fF
C4731 INVX1_LOC_17/A INVX1_LOC_28/Y 0.01fF
C4732 NOR2X1_LOC_686/B INVX1_LOC_38/A 0.01fF
C4733 INVX1_LOC_31/A INVX1_LOC_94/Y 0.28fF
C4734 INVX1_LOC_130/A NAND2X1_LOC_454/Y 0.03fF
C4735 NOR2X1_LOC_759/Y INVX1_LOC_290/Y 0.02fF
C4736 NAND2X1_LOC_850/A VDD -0.00fF
C4737 NOR2X1_LOC_103/Y NOR2X1_LOC_39/Y 0.07fF
C4738 D_INPUT_4 INVX1_LOC_76/A 0.00fF
C4739 INVX1_LOC_17/A INVX1_LOC_270/A 0.03fF
C4740 INVX1_LOC_299/A INVX1_LOC_23/A 0.03fF
C4741 INVX1_LOC_263/A NOR2X1_LOC_155/A 0.01fF
C4742 INVX1_LOC_287/A NOR2X1_LOC_710/B 0.32fF
C4743 INVX1_LOC_202/A INVX1_LOC_290/Y 0.02fF
C4744 NAND2X1_LOC_276/Y NAND2X1_LOC_63/Y 0.02fF
C4745 INVX1_LOC_36/A NOR2X1_LOC_158/B 0.03fF
C4746 INVX1_LOC_298/Y NOR2X1_LOC_590/A 0.18fF
C4747 INVX1_LOC_161/Y NOR2X1_LOC_686/a_36_216# 0.01fF
C4748 NAND2X1_LOC_332/Y INVX1_LOC_272/A 0.01fF
C4749 INVX1_LOC_75/A NOR2X1_LOC_309/a_36_216# 0.00fF
C4750 INVX1_LOC_64/A NOR2X1_LOC_456/a_36_216# 0.01fF
C4751 NAND2X1_LOC_479/Y INVX1_LOC_179/A 0.03fF
C4752 INVX1_LOC_30/A NAND2X1_LOC_72/B 0.03fF
C4753 INVX1_LOC_21/A INVX1_LOC_5/A 0.34fF
C4754 INVX1_LOC_200/Y INVX1_LOC_200/A 0.03fF
C4755 NOR2X1_LOC_197/A NOR2X1_LOC_727/B 0.02fF
C4756 NOR2X1_LOC_6/B NAND2X1_LOC_82/Y 0.10fF
C4757 NAND2X1_LOC_462/B NAND2X1_LOC_624/a_36_24# 0.00fF
C4758 NOR2X1_LOC_103/Y NAND2X1_LOC_205/A 0.03fF
C4759 INVX1_LOC_233/A NAND2X1_LOC_579/A 0.10fF
C4760 INVX1_LOC_36/A NOR2X1_LOC_30/Y 0.01fF
C4761 NOR2X1_LOC_641/B NOR2X1_LOC_621/B 0.04fF
C4762 INVX1_LOC_142/A INVX1_LOC_271/Y 0.02fF
C4763 NOR2X1_LOC_433/A NOR2X1_LOC_677/a_36_216# 0.00fF
C4764 NOR2X1_LOC_142/Y NOR2X1_LOC_755/Y 0.09fF
C4765 INVX1_LOC_162/Y NAND2X1_LOC_74/B 0.01fF
C4766 D_INPUT_0 NOR2X1_LOC_489/A 0.03fF
C4767 D_INPUT_1 INVX1_LOC_11/A 0.30fF
C4768 NAND2X1_LOC_35/Y NOR2X1_LOC_92/Y 0.14fF
C4769 NOR2X1_LOC_67/A NOR2X1_LOC_673/a_36_216# 0.01fF
C4770 NOR2X1_LOC_465/a_36_216# NAND2X1_LOC_190/Y 0.00fF
C4771 INVX1_LOC_64/A NOR2X1_LOC_468/Y 0.00fF
C4772 NOR2X1_LOC_596/A INVX1_LOC_4/A 0.07fF
C4773 INVX1_LOC_314/Y INVX1_LOC_15/A 0.07fF
C4774 D_INPUT_1 NAND2X1_LOC_381/Y 0.02fF
C4775 INVX1_LOC_36/A NOR2X1_LOC_301/A 0.04fF
C4776 NOR2X1_LOC_448/A INVX1_LOC_91/A 0.01fF
C4777 NOR2X1_LOC_152/Y INVX1_LOC_32/A 0.01fF
C4778 NAND2X1_LOC_464/Y NAND2X1_LOC_254/Y 0.01fF
C4779 INVX1_LOC_64/A NAND2X1_LOC_190/Y 0.10fF
C4780 INVX1_LOC_86/A VDD 0.12fF
C4781 INVX1_LOC_113/Y INVX1_LOC_32/A 0.03fF
C4782 INVX1_LOC_125/Y NAND2X1_LOC_447/Y 0.17fF
C4783 NOR2X1_LOC_284/B INVX1_LOC_19/A 0.02fF
C4784 NOR2X1_LOC_387/A INVX1_LOC_46/A 0.03fF
C4785 INVX1_LOC_313/Y INVX1_LOC_54/A 0.03fF
C4786 INVX1_LOC_256/A NOR2X1_LOC_678/A 1.31fF
C4787 NOR2X1_LOC_74/A NAND2X1_LOC_472/Y 0.17fF
C4788 INVX1_LOC_17/A NOR2X1_LOC_109/Y 0.14fF
C4789 INVX1_LOC_286/Y INVX1_LOC_57/A 0.08fF
C4790 INVX1_LOC_89/A NOR2X1_LOC_88/A 0.00fF
C4791 NOR2X1_LOC_503/a_36_216# NAND2X1_LOC_802/Y -0.02fF
C4792 INVX1_LOC_233/Y NAND2X1_LOC_550/A 0.10fF
C4793 INVX1_LOC_81/A NAND2X1_LOC_454/Y 0.03fF
C4794 INVX1_LOC_82/A NOR2X1_LOC_554/A 0.24fF
C4795 NOR2X1_LOC_92/Y NAND2X1_LOC_571/Y 0.34fF
C4796 INVX1_LOC_18/A NOR2X1_LOC_635/B 0.03fF
C4797 INVX1_LOC_90/A NAND2X1_LOC_798/B 0.25fF
C4798 NOR2X1_LOC_524/Y INVX1_LOC_23/A 0.00fF
C4799 INVX1_LOC_232/A INVX1_LOC_19/A 0.14fF
C4800 NAND2X1_LOC_53/Y NOR2X1_LOC_590/Y 0.01fF
C4801 NOR2X1_LOC_392/B INVX1_LOC_47/Y 0.10fF
C4802 NOR2X1_LOC_152/Y NAND2X1_LOC_175/Y 0.60fF
C4803 NOR2X1_LOC_181/Y INVX1_LOC_15/A 0.11fF
C4804 INVX1_LOC_17/Y INVX1_LOC_217/A 0.02fF
C4805 INVX1_LOC_64/A NOR2X1_LOC_389/A 0.22fF
C4806 NAND2X1_LOC_725/B INVX1_LOC_234/Y 0.06fF
C4807 NOR2X1_LOC_790/A NOR2X1_LOC_793/A 0.02fF
C4808 NAND2X1_LOC_579/A NAND2X1_LOC_703/Y 0.03fF
C4809 INVX1_LOC_11/A NOR2X1_LOC_652/Y -0.03fF
C4810 INVX1_LOC_18/A NOR2X1_LOC_748/A 0.17fF
C4811 NOR2X1_LOC_139/Y NOR2X1_LOC_137/Y 0.10fF
C4812 NOR2X1_LOC_15/Y INVX1_LOC_239/A 0.07fF
C4813 NAND2X1_LOC_844/a_36_24# INVX1_LOC_118/A 0.00fF
C4814 NOR2X1_LOC_516/B NOR2X1_LOC_830/Y 0.01fF
C4815 NAND2X1_LOC_553/a_36_24# INVX1_LOC_284/A 0.00fF
C4816 NAND2X1_LOC_468/B NAND2X1_LOC_440/a_36_24# 0.02fF
C4817 NAND2X1_LOC_655/B INVX1_LOC_20/A 0.00fF
C4818 NAND2X1_LOC_540/a_36_24# NOR2X1_LOC_160/B 0.00fF
C4819 NAND2X1_LOC_114/B INVX1_LOC_50/Y 0.32fF
C4820 NAND2X1_LOC_662/Y NAND2X1_LOC_74/B 0.02fF
C4821 INVX1_LOC_21/A NAND2X1_LOC_337/B 0.34fF
C4822 NOR2X1_LOC_69/A INVX1_LOC_76/A 0.03fF
C4823 VDD NOR2X1_LOC_346/Y 0.24fF
C4824 INVX1_LOC_21/A NOR2X1_LOC_816/A 0.12fF
C4825 NOR2X1_LOC_191/B INVX1_LOC_57/A 0.20fF
C4826 NOR2X1_LOC_196/Y INVX1_LOC_108/A 0.14fF
C4827 NOR2X1_LOC_778/B INVX1_LOC_15/A 0.28fF
C4828 INPUT_3 NOR2X1_LOC_655/a_36_216# 0.00fF
C4829 NOR2X1_LOC_320/Y INVX1_LOC_291/A 0.02fF
C4830 INVX1_LOC_227/A INVX1_LOC_29/A 0.06fF
C4831 NAND2X1_LOC_564/B INVX1_LOC_42/A 0.07fF
C4832 INVX1_LOC_20/Y INVX1_LOC_63/A 0.01fF
C4833 INVX1_LOC_89/A INVX1_LOC_186/Y 0.07fF
C4834 NAND2X1_LOC_319/A INVX1_LOC_12/A 0.01fF
C4835 INVX1_LOC_103/A INVX1_LOC_88/A 0.12fF
C4836 NOR2X1_LOC_82/A NOR2X1_LOC_271/B 0.07fF
C4837 NOR2X1_LOC_309/Y NOR2X1_LOC_301/A 0.07fF
C4838 NOR2X1_LOC_763/Y INVX1_LOC_29/A 0.02fF
C4839 NOR2X1_LOC_238/Y NOR2X1_LOC_754/Y 0.17fF
C4840 NOR2X1_LOC_431/Y INVX1_LOC_53/A 0.01fF
C4841 INVX1_LOC_16/A INVX1_LOC_3/Y 4.58fF
C4842 NOR2X1_LOC_468/Y INVX1_LOC_43/Y 0.33fF
C4843 INVX1_LOC_278/A INVX1_LOC_314/Y 0.01fF
C4844 INVX1_LOC_64/A NOR2X1_LOC_596/A 0.07fF
C4845 INVX1_LOC_286/A NOR2X1_LOC_79/a_36_216# 0.01fF
C4846 NOR2X1_LOC_35/Y INVX1_LOC_117/A 0.10fF
C4847 NAND2X1_LOC_728/Y NOR2X1_LOC_304/Y 0.02fF
C4848 D_INPUT_1 NOR2X1_LOC_593/Y 0.03fF
C4849 NOR2X1_LOC_91/A NOR2X1_LOC_315/Y 0.03fF
C4850 INVX1_LOC_206/Y NOR2X1_LOC_155/A 0.03fF
C4851 INVX1_LOC_163/A NAND2X1_LOC_577/A 0.07fF
C4852 INVX1_LOC_208/A INVX1_LOC_4/Y 0.01fF
C4853 NAND2X1_LOC_35/Y NAND2X1_LOC_837/Y 0.07fF
C4854 NOR2X1_LOC_458/a_36_216# NOR2X1_LOC_570/B 0.02fF
C4855 INVX1_LOC_299/A INVX1_LOC_31/A 0.10fF
C4856 INVX1_LOC_162/A INVX1_LOC_23/A 0.02fF
C4857 NAND2X1_LOC_778/Y NOR2X1_LOC_91/Y 0.01fF
C4858 NOR2X1_LOC_516/B INVX1_LOC_4/Y 0.15fF
C4859 INVX1_LOC_178/A NAND2X1_LOC_354/Y 0.53fF
C4860 INVX1_LOC_256/Y NOR2X1_LOC_278/Y 0.04fF
C4861 NOR2X1_LOC_795/Y NOR2X1_LOC_383/B 0.00fF
C4862 NOR2X1_LOC_791/Y NAND2X1_LOC_198/B 0.01fF
C4863 INVX1_LOC_155/Y INVX1_LOC_53/A 0.02fF
C4864 INVX1_LOC_93/Y NOR2X1_LOC_612/Y 0.02fF
C4865 NAND2X1_LOC_338/B NOR2X1_LOC_438/Y 0.02fF
C4866 INVX1_LOC_9/Y INVX1_LOC_78/A 0.43fF
C4867 INVX1_LOC_304/Y INVX1_LOC_200/Y 0.00fF
C4868 NOR2X1_LOC_113/B NAND2X1_LOC_475/Y 0.40fF
C4869 NAND2X1_LOC_370/a_36_24# NAND2X1_LOC_833/Y 0.00fF
C4870 NOR2X1_LOC_703/A INVX1_LOC_29/A 0.03fF
C4871 D_INPUT_1 NOR2X1_LOC_52/B 0.07fF
C4872 NOR2X1_LOC_315/Y INVX1_LOC_23/A 0.08fF
C4873 NAND2X1_LOC_564/B INVX1_LOC_78/A 0.07fF
C4874 INVX1_LOC_191/Y INVX1_LOC_296/A 0.01fF
C4875 NOR2X1_LOC_647/A INVX1_LOC_40/A 0.14fF
C4876 NOR2X1_LOC_600/Y NOR2X1_LOC_155/A 0.00fF
C4877 INVX1_LOC_259/Y INVX1_LOC_85/A 0.00fF
C4878 NOR2X1_LOC_598/B INVX1_LOC_104/A 1.46fF
C4879 NOR2X1_LOC_113/A NOR2X1_LOC_216/B 0.04fF
C4880 NOR2X1_LOC_433/A NOR2X1_LOC_652/Y 0.07fF
C4881 NOR2X1_LOC_405/A NOR2X1_LOC_216/B 0.10fF
C4882 INVX1_LOC_293/A INVX1_LOC_31/A 0.03fF
C4883 NOR2X1_LOC_273/Y NOR2X1_LOC_454/Y 0.37fF
C4884 INVX1_LOC_17/A INVX1_LOC_36/A 2.12fF
C4885 NOR2X1_LOC_498/Y NAND2X1_LOC_35/Y 0.01fF
C4886 NOR2X1_LOC_99/Y INVX1_LOC_59/Y 0.01fF
C4887 NOR2X1_LOC_15/Y NOR2X1_LOC_91/Y 0.04fF
C4888 INVX1_LOC_83/Y NOR2X1_LOC_727/B 0.01fF
C4889 INVX1_LOC_303/Y NOR2X1_LOC_691/B 0.10fF
C4890 INVX1_LOC_117/A NAND2X1_LOC_236/a_36_24# 0.00fF
C4891 NOR2X1_LOC_510/B NOR2X1_LOC_56/Y 0.13fF
C4892 NOR2X1_LOC_510/Y NOR2X1_LOC_637/B 0.01fF
C4893 NOR2X1_LOC_84/a_36_216# NOR2X1_LOC_392/Y 0.00fF
C4894 INVX1_LOC_161/A NAND2X1_LOC_389/a_36_24# 0.00fF
C4895 INVX1_LOC_269/A NOR2X1_LOC_360/Y 0.10fF
C4896 INVX1_LOC_64/A NOR2X1_LOC_844/A 0.53fF
C4897 INVX1_LOC_90/A INVX1_LOC_47/Y 0.21fF
C4898 NOR2X1_LOC_15/Y NOR2X1_LOC_359/Y 0.03fF
C4899 NOR2X1_LOC_724/Y INVX1_LOC_15/A 0.74fF
C4900 D_INPUT_0 NOR2X1_LOC_334/Y 0.00fF
C4901 INVX1_LOC_50/A NOR2X1_LOC_500/Y 0.07fF
C4902 INVX1_LOC_299/A INVX1_LOC_111/A 0.11fF
C4903 NOR2X1_LOC_186/Y INVX1_LOC_34/A 0.03fF
C4904 NOR2X1_LOC_471/Y INVX1_LOC_36/A 0.01fF
C4905 NOR2X1_LOC_389/B INVX1_LOC_47/Y 0.02fF
C4906 NAND2X1_LOC_55/a_36_24# INVX1_LOC_13/Y 0.00fF
C4907 INVX1_LOC_75/A GATE_222 0.03fF
C4908 INVX1_LOC_28/A INVX1_LOC_3/Y 0.23fF
C4909 INVX1_LOC_256/A INVX1_LOC_305/A 0.03fF
C4910 INVX1_LOC_298/Y INVX1_LOC_227/A 0.02fF
C4911 NOR2X1_LOC_441/Y NOR2X1_LOC_361/a_36_216# 0.01fF
C4912 NAND2X1_LOC_503/a_36_24# NAND2X1_LOC_510/A 0.00fF
C4913 INVX1_LOC_313/A INVX1_LOC_94/Y 0.04fF
C4914 NAND2X1_LOC_208/B NAND2X1_LOC_198/a_36_24# 0.02fF
C4915 NOR2X1_LOC_67/A NAND2X1_LOC_549/Y 0.01fF
C4916 VDD NOR2X1_LOC_510/B 0.18fF
C4917 NOR2X1_LOC_685/A INVX1_LOC_19/A 0.01fF
C4918 NAND2X1_LOC_493/Y NAND2X1_LOC_787/B 0.03fF
C4919 INVX1_LOC_17/A INVX1_LOC_145/A 0.02fF
C4920 NOR2X1_LOC_321/Y INVX1_LOC_33/A 0.15fF
C4921 NOR2X1_LOC_52/B NOR2X1_LOC_652/Y 0.07fF
C4922 INPUT_3 NOR2X1_LOC_554/B 0.08fF
C4923 INVX1_LOC_25/A NOR2X1_LOC_62/a_36_216# 0.00fF
C4924 INVX1_LOC_186/A INVX1_LOC_19/A 0.10fF
C4925 NAND2X1_LOC_153/a_36_24# INVX1_LOC_150/Y 0.00fF
C4926 INVX1_LOC_35/A INVX1_LOC_179/Y 0.00fF
C4927 INVX1_LOC_58/A INVX1_LOC_16/A 0.19fF
C4928 INVX1_LOC_139/Y INVX1_LOC_179/A 2.28fF
C4929 NOR2X1_LOC_773/a_36_216# NAND2X1_LOC_474/Y 0.00fF
C4930 INVX1_LOC_64/A NOR2X1_LOC_399/Y 0.03fF
C4931 NOR2X1_LOC_165/a_36_216# INVX1_LOC_102/A 0.01fF
C4932 INVX1_LOC_135/A NOR2X1_LOC_693/Y 0.10fF
C4933 INVX1_LOC_64/A NOR2X1_LOC_220/A 0.03fF
C4934 NAND2X1_LOC_785/A INVX1_LOC_93/A 0.09fF
C4935 NAND2X1_LOC_741/B NOR2X1_LOC_599/A 0.03fF
C4936 NOR2X1_LOC_168/B INVX1_LOC_50/Y 3.03fF
C4937 INVX1_LOC_17/A NOR2X1_LOC_237/Y 0.07fF
C4938 NOR2X1_LOC_332/Y INVX1_LOC_280/A 0.00fF
C4939 NOR2X1_LOC_667/A NAND2X1_LOC_552/A 0.03fF
C4940 INVX1_LOC_50/A INVX1_LOC_10/A 0.69fF
C4941 INVX1_LOC_269/A INVX1_LOC_207/A 0.03fF
C4942 NAND2X1_LOC_53/Y INVX1_LOC_105/A 0.06fF
C4943 NOR2X1_LOC_471/Y NOR2X1_LOC_208/Y 0.02fF
C4944 INVX1_LOC_34/A NAND2X1_LOC_724/A 0.07fF
C4945 NOR2X1_LOC_186/Y NAND2X1_LOC_231/Y 0.10fF
C4946 NAND2X1_LOC_659/B NOR2X1_LOC_662/A 0.10fF
C4947 INVX1_LOC_49/Y NAND2X1_LOC_642/Y 0.00fF
C4948 INVX1_LOC_20/Y NAND2X1_LOC_223/B 0.23fF
C4949 NOR2X1_LOC_202/a_36_216# INVX1_LOC_63/Y 0.01fF
C4950 INVX1_LOC_159/Y INVX1_LOC_12/A 0.03fF
C4951 NAND2X1_LOC_72/Y NOR2X1_LOC_500/Y 0.01fF
C4952 INVX1_LOC_49/A NOR2X1_LOC_250/A 0.06fF
C4953 INVX1_LOC_89/A NOR2X1_LOC_843/B 0.06fF
C4954 INVX1_LOC_136/A INVX1_LOC_223/A 0.03fF
C4955 NOR2X1_LOC_226/A NOR2X1_LOC_81/Y 0.03fF
C4956 INVX1_LOC_25/A NOR2X1_LOC_719/B 0.02fF
C4957 NAND2X1_LOC_643/a_36_24# INVX1_LOC_49/Y 0.00fF
C4958 NOR2X1_LOC_559/B NAND2X1_LOC_114/B 0.08fF
C4959 INVX1_LOC_265/A INVX1_LOC_14/A 0.22fF
C4960 D_INPUT_0 NAND2X1_LOC_464/B 0.07fF
C4961 NAND2X1_LOC_447/Y INVX1_LOC_19/A 0.03fF
C4962 NOR2X1_LOC_506/Y INVX1_LOC_54/A 0.29fF
C4963 NAND2X1_LOC_711/B NAND2X1_LOC_711/Y 0.04fF
C4964 INVX1_LOC_33/Y NOR2X1_LOC_841/A 0.09fF
C4965 INVX1_LOC_287/A INVX1_LOC_89/A 0.01fF
C4966 INVX1_LOC_38/A NAND2X1_LOC_798/B 0.07fF
C4967 NOR2X1_LOC_667/A INVX1_LOC_178/A 0.10fF
C4968 INVX1_LOC_5/A NAND2X1_LOC_6/a_36_24# 0.02fF
C4969 NOR2X1_LOC_91/A NOR2X1_LOC_166/Y 0.03fF
C4970 INVX1_LOC_248/A INVX1_LOC_178/A 0.10fF
C4971 INVX1_LOC_21/A NOR2X1_LOC_773/Y 0.14fF
C4972 INVX1_LOC_35/A NOR2X1_LOC_561/Y 0.08fF
C4973 NAND2X1_LOC_573/Y NAND2X1_LOC_231/Y 0.10fF
C4974 NOR2X1_LOC_775/Y INVX1_LOC_26/Y 0.02fF
C4975 VDD NOR2X1_LOC_662/A 1.24fF
C4976 NOR2X1_LOC_68/A NOR2X1_LOC_791/B 0.03fF
C4977 INVX1_LOC_17/A NOR2X1_LOC_309/Y 0.20fF
C4978 NAND2X1_LOC_559/Y NAND2X1_LOC_722/A 0.07fF
C4979 NOR2X1_LOC_329/B NOR2X1_LOC_447/A 0.00fF
C4980 INVX1_LOC_5/A NOR2X1_LOC_521/Y 0.01fF
C4981 INVX1_LOC_34/A NOR2X1_LOC_45/Y 0.12fF
C4982 INVX1_LOC_11/A NOR2X1_LOC_591/Y 0.34fF
C4983 NOR2X1_LOC_843/A NOR2X1_LOC_160/B 0.22fF
C4984 INVX1_LOC_2/A NAND2X1_LOC_538/Y 0.07fF
C4985 INVX1_LOC_245/Y NOR2X1_LOC_718/B 0.03fF
C4986 NOR2X1_LOC_468/Y NAND2X1_LOC_850/Y 0.04fF
C4987 INVX1_LOC_6/A INVX1_LOC_94/Y 0.03fF
C4988 NAND2X1_LOC_650/B INVX1_LOC_29/A 0.02fF
C4989 INVX1_LOC_274/A NOR2X1_LOC_197/B 0.06fF
C4990 NAND2X1_LOC_114/B NOR2X1_LOC_6/B 0.07fF
C4991 INVX1_LOC_140/A INVX1_LOC_173/A 0.08fF
C4992 INVX1_LOC_5/A NOR2X1_LOC_565/B 0.03fF
C4993 NOR2X1_LOC_590/A INVX1_LOC_8/A 0.12fF
C4994 INVX1_LOC_58/A INVX1_LOC_28/A 0.40fF
C4995 NOR2X1_LOC_226/A NAND2X1_LOC_538/Y 0.10fF
C4996 INVX1_LOC_217/A NOR2X1_LOC_495/Y 0.15fF
C4997 INVX1_LOC_135/A INVX1_LOC_253/Y 0.30fF
C4998 INVX1_LOC_178/A NOR2X1_LOC_521/Y 0.26fF
C4999 NOR2X1_LOC_657/B INVX1_LOC_15/A 0.07fF
C5000 INVX1_LOC_161/Y NOR2X1_LOC_511/a_36_216# 0.00fF
C5001 NAND2X1_LOC_9/Y NOR2X1_LOC_756/Y 0.01fF
C5002 INVX1_LOC_11/A NOR2X1_LOC_620/B 0.01fF
C5003 NOR2X1_LOC_130/A INVX1_LOC_306/Y 0.03fF
C5004 NAND2X1_LOC_808/A NOR2X1_LOC_406/A 0.02fF
C5005 NAND2X1_LOC_569/B INPUT_1 0.04fF
C5006 INVX1_LOC_25/A INVX1_LOC_73/A 0.07fF
C5007 INVX1_LOC_208/A NOR2X1_LOC_205/Y 0.01fF
C5008 NAND2X1_LOC_720/a_36_24# NAND2X1_LOC_325/Y 0.01fF
C5009 INVX1_LOC_18/A NAND2X1_LOC_283/a_36_24# 0.01fF
C5010 NOR2X1_LOC_274/Y NAND2X1_LOC_656/A 0.00fF
C5011 NOR2X1_LOC_448/B INVX1_LOC_22/A 0.01fF
C5012 NOR2X1_LOC_273/Y INVX1_LOC_77/A 0.03fF
C5013 INVX1_LOC_214/A NOR2X1_LOC_816/A 0.03fF
C5014 INVX1_LOC_256/A NOR2X1_LOC_191/A 0.00fF
C5015 NOR2X1_LOC_142/Y INVX1_LOC_72/A 0.26fF
C5016 INVX1_LOC_237/A NOR2X1_LOC_32/Y 0.09fF
C5017 NAND2X1_LOC_231/Y NOR2X1_LOC_45/Y 0.07fF
C5018 NOR2X1_LOC_667/A NOR2X1_LOC_816/A 0.10fF
C5019 NOR2X1_LOC_721/Y INVX1_LOC_57/A 0.03fF
C5020 INVX1_LOC_21/A NOR2X1_LOC_332/A 0.14fF
C5021 INVX1_LOC_248/A NAND2X1_LOC_337/B 0.03fF
C5022 INVX1_LOC_77/A NOR2X1_LOC_759/Y 0.03fF
C5023 INVX1_LOC_248/A NOR2X1_LOC_816/A 0.03fF
C5024 NOR2X1_LOC_274/a_36_216# INVX1_LOC_77/A 0.00fF
C5025 INVX1_LOC_202/A INVX1_LOC_77/A 0.07fF
C5026 INVX1_LOC_292/A NOR2X1_LOC_203/Y 0.02fF
C5027 INVX1_LOC_136/A INVX1_LOC_162/Y 0.00fF
C5028 INVX1_LOC_218/Y NAND2X1_LOC_338/B 0.04fF
C5029 INVX1_LOC_11/A NOR2X1_LOC_553/Y 0.03fF
C5030 NOR2X1_LOC_68/A NOR2X1_LOC_124/B 0.02fF
C5031 NOR2X1_LOC_791/Y NOR2X1_LOC_76/a_36_216# 0.00fF
C5032 NAND2X1_LOC_553/A NOR2X1_LOC_756/Y 0.31fF
C5033 INVX1_LOC_45/Y NOR2X1_LOC_388/Y 0.18fF
C5034 NOR2X1_LOC_68/A NOR2X1_LOC_802/A 0.01fF
C5035 INVX1_LOC_78/A NOR2X1_LOC_279/Y 0.07fF
C5036 INVX1_LOC_226/Y INVX1_LOC_61/Y 0.40fF
C5037 INVX1_LOC_255/Y NOR2X1_LOC_647/a_36_216# 0.00fF
C5038 INVX1_LOC_54/Y NAND2X1_LOC_364/A 0.04fF
C5039 NOR2X1_LOC_186/Y INVX1_LOC_131/A 0.02fF
C5040 NAND2X1_LOC_384/a_36_24# NOR2X1_LOC_103/Y 0.00fF
C5041 INVX1_LOC_30/Y NAND2X1_LOC_114/B 0.02fF
C5042 INVX1_LOC_41/A NAND2X1_LOC_786/a_36_24# 0.00fF
C5043 NAND2X1_LOC_227/Y INVX1_LOC_10/A 0.01fF
C5044 INVX1_LOC_21/A INVX1_LOC_140/A 0.07fF
C5045 NOR2X1_LOC_677/Y NAND2X1_LOC_655/A 0.01fF
C5046 INVX1_LOC_286/A NAND2X1_LOC_793/B 0.05fF
C5047 INVX1_LOC_119/A NOR2X1_LOC_637/Y 0.00fF
C5048 NOR2X1_LOC_219/Y INVX1_LOC_30/A 0.00fF
C5049 NOR2X1_LOC_561/A INVX1_LOC_47/Y 0.02fF
C5050 NOR2X1_LOC_778/B NOR2X1_LOC_168/Y 0.04fF
C5051 INVX1_LOC_304/Y NOR2X1_LOC_495/Y 0.04fF
C5052 NOR2X1_LOC_506/Y NOR2X1_LOC_48/B 0.08fF
C5053 NOR2X1_LOC_66/Y NOR2X1_LOC_631/A 0.13fF
C5054 INVX1_LOC_1/A NOR2X1_LOC_738/A 0.03fF
C5055 NOR2X1_LOC_591/Y NOR2X1_LOC_433/A 0.02fF
C5056 NOR2X1_LOC_186/Y INPUT_0 0.04fF
C5057 NOR2X1_LOC_846/Y NOR2X1_LOC_188/A 0.08fF
C5058 NOR2X1_LOC_56/Y INVX1_LOC_57/A 0.03fF
C5059 INVX1_LOC_34/A INVX1_LOC_225/A 0.07fF
C5060 NOR2X1_LOC_361/B NAND2X1_LOC_850/A 0.16fF
C5061 NOR2X1_LOC_646/A NOR2X1_LOC_68/A -0.01fF
C5062 INVX1_LOC_136/A NAND2X1_LOC_662/Y 0.06fF
C5063 INVX1_LOC_1/A INVX1_LOC_73/A 0.07fF
C5064 NOR2X1_LOC_769/A GATE_662 0.07fF
C5065 INVX1_LOC_155/A INVX1_LOC_177/A 0.00fF
C5066 NOR2X1_LOC_287/a_36_216# NOR2X1_LOC_288/A 0.00fF
C5067 NOR2X1_LOC_530/Y INPUT_1 0.01fF
C5068 D_INPUT_1 INVX1_LOC_74/A 0.02fF
C5069 INVX1_LOC_243/Y VDD 0.21fF
C5070 NOR2X1_LOC_180/B NOR2X1_LOC_794/B 0.03fF
C5071 NAND2X1_LOC_573/Y INPUT_0 0.01fF
C5072 INVX1_LOC_78/Y INVX1_LOC_50/Y 0.02fF
C5073 NOR2X1_LOC_831/B NOR2X1_LOC_114/Y 0.02fF
C5074 NAND2X1_LOC_563/Y NOR2X1_LOC_514/Y 0.03fF
C5075 INVX1_LOC_230/Y NOR2X1_LOC_130/Y 0.02fF
C5076 INVX1_LOC_146/Y INVX1_LOC_57/A 0.01fF
C5077 NOR2X1_LOC_15/Y NOR2X1_LOC_151/a_36_216# 0.00fF
C5078 INVX1_LOC_83/A NAND2X1_LOC_510/A 0.15fF
C5079 VDD INVX1_LOC_57/A 3.74fF
C5080 NOR2X1_LOC_261/A INVX1_LOC_78/A 0.01fF
C5081 INVX1_LOC_215/Y INVX1_LOC_28/A 0.78fF
C5082 NAND2X1_LOC_863/Y NAND2X1_LOC_863/B 0.03fF
C5083 NAND2X1_LOC_724/A INPUT_0 0.07fF
C5084 NAND2X1_LOC_338/B NOR2X1_LOC_340/Y 0.02fF
C5085 INVX1_LOC_9/Y NOR2X1_LOC_152/Y 0.08fF
C5086 NOR2X1_LOC_524/Y INVX1_LOC_313/A 0.10fF
C5087 INVX1_LOC_250/A NAND2X1_LOC_808/A 0.04fF
C5088 NOR2X1_LOC_721/a_36_216# INVX1_LOC_62/Y 0.01fF
C5089 INVX1_LOC_120/A NOR2X1_LOC_500/B 0.00fF
C5090 NAND2X1_LOC_552/A INVX1_LOC_304/A 0.04fF
C5091 INVX1_LOC_225/A NAND2X1_LOC_231/Y 0.01fF
C5092 INVX1_LOC_18/A INVX1_LOC_150/A 0.02fF
C5093 INVX1_LOC_64/A NAND2X1_LOC_469/B 0.04fF
C5094 NOR2X1_LOC_383/B INVX1_LOC_281/A 1.48fF
C5095 INVX1_LOC_35/A INVX1_LOC_76/A 0.09fF
C5096 NOR2X1_LOC_612/Y INVX1_LOC_87/A 0.00fF
C5097 INVX1_LOC_34/A NAND2X1_LOC_852/Y 0.10fF
C5098 NOR2X1_LOC_358/a_36_216# NAND2X1_LOC_454/Y 0.01fF
C5099 NAND2X1_LOC_63/Y INVX1_LOC_125/A 0.03fF
C5100 NOR2X1_LOC_357/Y NOR2X1_LOC_665/a_36_216# 0.00fF
C5101 INVX1_LOC_89/A INVX1_LOC_18/A 0.36fF
C5102 INVX1_LOC_5/A NOR2X1_LOC_670/Y 0.00fF
C5103 NAND2X1_LOC_848/A NAND2X1_LOC_464/B 0.07fF
C5104 NAND2X1_LOC_345/a_36_24# INVX1_LOC_18/A 0.00fF
C5105 NAND2X1_LOC_96/A INVX1_LOC_23/A 0.14fF
C5106 INVX1_LOC_291/A NAND2X1_LOC_175/Y 0.07fF
C5107 NAND2X1_LOC_263/a_36_24# INVX1_LOC_19/A 0.01fF
C5108 NOR2X1_LOC_100/A NOR2X1_LOC_87/Y 0.03fF
C5109 NOR2X1_LOC_843/A NOR2X1_LOC_516/B 0.03fF
C5110 INVX1_LOC_178/A INVX1_LOC_255/A 0.07fF
C5111 NOR2X1_LOC_383/B NOR2X1_LOC_499/B 0.02fF
C5112 INVX1_LOC_64/A NOR2X1_LOC_447/B 0.11fF
C5113 NOR2X1_LOC_226/A NOR2X1_LOC_709/A 0.33fF
C5114 NAND2X1_LOC_181/Y NOR2X1_LOC_84/Y 0.23fF
C5115 NAND2X1_LOC_432/a_36_24# INVX1_LOC_15/A 0.01fF
C5116 NOR2X1_LOC_589/A INVX1_LOC_63/Y 0.19fF
C5117 NOR2X1_LOC_655/B NAND2X1_LOC_338/B 0.10fF
C5118 NOR2X1_LOC_67/Y INVX1_LOC_29/A 0.36fF
C5119 NOR2X1_LOC_78/B NOR2X1_LOC_131/A 0.01fF
C5120 NAND2X1_LOC_389/a_36_24# INPUT_0 0.01fF
C5121 INVX1_LOC_247/Y NOR2X1_LOC_703/A 0.00fF
C5122 NOR2X1_LOC_496/Y INVX1_LOC_20/A 0.16fF
C5123 INVX1_LOC_94/Y NOR2X1_LOC_117/Y 0.07fF
C5124 INVX1_LOC_24/A NOR2X1_LOC_356/A 0.07fF
C5125 INVX1_LOC_49/A NOR2X1_LOC_106/A 0.03fF
C5126 NOR2X1_LOC_570/A INVX1_LOC_104/A 0.08fF
C5127 NAND2X1_LOC_303/Y INVX1_LOC_11/Y 0.05fF
C5128 NAND2X1_LOC_351/a_36_24# NAND2X1_LOC_96/A 0.00fF
C5129 NOR2X1_LOC_456/Y INVX1_LOC_9/A 0.07fF
C5130 NAND2X1_LOC_562/B NOR2X1_LOC_521/Y 0.00fF
C5131 NOR2X1_LOC_667/A NOR2X1_LOC_773/Y 0.15fF
C5132 INVX1_LOC_170/A INPUT_0 0.00fF
C5133 NAND2X1_LOC_659/B NOR2X1_LOC_475/A 0.03fF
C5134 VDD INVX1_LOC_252/A 0.12fF
C5135 NOR2X1_LOC_113/B INVX1_LOC_30/A 0.04fF
C5136 NOR2X1_LOC_383/B NOR2X1_LOC_862/B 0.02fF
C5137 INVX1_LOC_50/A INVX1_LOC_307/A 0.08fF
C5138 NAND2X1_LOC_392/A INVX1_LOC_256/Y 0.02fF
C5139 NOR2X1_LOC_861/Y NAND2X1_LOC_206/B 0.17fF
C5140 NAND2X1_LOC_303/Y NOR2X1_LOC_421/Y 0.07fF
C5141 NAND2X1_LOC_736/B NOR2X1_LOC_576/B 0.03fF
C5142 NOR2X1_LOC_641/Y INVX1_LOC_58/Y 0.01fF
C5143 NAND2X1_LOC_793/B INVX1_LOC_54/A 0.12fF
C5144 INVX1_LOC_45/A INVX1_LOC_286/A 1.07fF
C5145 NOR2X1_LOC_576/B GATE_811 0.02fF
C5146 INVX1_LOC_50/A NOR2X1_LOC_445/B 0.07fF
C5147 NOR2X1_LOC_474/A NOR2X1_LOC_575/Y 0.15fF
C5148 NAND2X1_LOC_607/a_36_24# INVX1_LOC_46/Y 0.01fF
C5149 INVX1_LOC_84/Y NOR2X1_LOC_375/Y 0.01fF
C5150 INVX1_LOC_286/A NOR2X1_LOC_568/A 0.01fF
C5151 NAND2X1_LOC_218/B INVX1_LOC_75/A 0.34fF
C5152 INVX1_LOC_271/A NOR2X1_LOC_88/Y 0.12fF
C5153 NOR2X1_LOC_142/Y INVX1_LOC_313/Y 0.02fF
C5154 NOR2X1_LOC_301/A INVX1_LOC_63/A 0.09fF
C5155 NAND2X1_LOC_358/Y NAND2X1_LOC_338/B 0.08fF
C5156 INVX1_LOC_24/A NOR2X1_LOC_74/A 0.13fF
C5157 NOR2X1_LOC_666/Y VDD 0.15fF
C5158 INVX1_LOC_88/A NOR2X1_LOC_137/Y 0.01fF
C5159 NOR2X1_LOC_273/Y NAND2X1_LOC_832/Y 0.03fF
C5160 INVX1_LOC_278/Y NAND2X1_LOC_168/a_36_24# 0.00fF
C5161 NAND2X1_LOC_564/B NAND2X1_LOC_860/Y 0.01fF
C5162 INVX1_LOC_25/Y INVX1_LOC_22/A 0.06fF
C5163 NOR2X1_LOC_106/Y INVX1_LOC_79/A 0.30fF
C5164 NAND2X1_LOC_207/B INVX1_LOC_4/Y 0.00fF
C5165 NOR2X1_LOC_207/a_36_216# INVX1_LOC_266/Y 0.01fF
C5166 NOR2X1_LOC_121/A NOR2X1_LOC_719/A 0.03fF
C5167 NAND2X1_LOC_358/Y NAND2X1_LOC_323/B 0.01fF
C5168 INVX1_LOC_75/A NOR2X1_LOC_577/Y 0.10fF
C5169 NOR2X1_LOC_99/B NOR2X1_LOC_537/Y 0.07fF
C5170 NOR2X1_LOC_379/Y INVX1_LOC_75/A 0.22fF
C5171 INVX1_LOC_57/Y NOR2X1_LOC_45/B 0.19fF
C5172 INVX1_LOC_24/A NOR2X1_LOC_9/Y 0.03fF
C5173 INVX1_LOC_94/A NAND2X1_LOC_309/a_36_24# 0.07fF
C5174 NOR2X1_LOC_415/Y INVX1_LOC_29/A 0.02fF
C5175 INPUT_1 NOR2X1_LOC_709/A 0.12fF
C5176 NAND2X1_LOC_257/a_36_24# NOR2X1_LOC_342/A 0.00fF
C5177 INVX1_LOC_132/A INPUT_0 0.08fF
C5178 NAND2X1_LOC_323/B NOR2X1_LOC_99/B 0.50fF
C5179 NAND2X1_LOC_72/Y NOR2X1_LOC_445/B 0.04fF
C5180 INVX1_LOC_225/A INVX1_LOC_131/A 0.03fF
C5181 D_INPUT_0 INVX1_LOC_218/A 0.51fF
C5182 INVX1_LOC_286/A INVX1_LOC_71/A 0.19fF
C5183 INVX1_LOC_7/A NOR2X1_LOC_121/A 0.03fF
C5184 NOR2X1_LOC_667/Y NOR2X1_LOC_305/Y 0.02fF
C5185 NAND2X1_LOC_640/Y INPUT_0 0.01fF
C5186 NOR2X1_LOC_557/Y NOR2X1_LOC_74/A 1.36fF
C5187 NOR2X1_LOC_406/A INVX1_LOC_92/A 0.03fF
C5188 NOR2X1_LOC_655/B INVX1_LOC_313/Y 0.01fF
C5189 NOR2X1_LOC_45/B NOR2X1_LOC_512/Y 0.01fF
C5190 NOR2X1_LOC_335/A INVX1_LOC_69/Y 0.01fF
C5191 NAND2X1_LOC_353/a_36_24# INVX1_LOC_28/A 0.00fF
C5192 INVX1_LOC_30/A NAND2X1_LOC_465/A 0.01fF
C5193 NOR2X1_LOC_89/A NOR2X1_LOC_318/A 0.12fF
C5194 INVX1_LOC_212/A NOR2X1_LOC_349/A 0.01fF
C5195 INVX1_LOC_255/Y INVX1_LOC_135/A 0.13fF
C5196 NOR2X1_LOC_740/a_36_216# INVX1_LOC_117/A 0.00fF
C5197 INVX1_LOC_72/A NAND2X1_LOC_274/a_36_24# 0.00fF
C5198 INVX1_LOC_17/A NOR2X1_LOC_865/A 0.04fF
C5199 INVX1_LOC_225/A INPUT_0 0.10fF
C5200 INVX1_LOC_41/A NOR2X1_LOC_730/B 0.01fF
C5201 NAND2X1_LOC_564/B NAND2X1_LOC_861/Y -0.02fF
C5202 INVX1_LOC_50/A INVX1_LOC_12/A 0.29fF
C5203 NOR2X1_LOC_690/A INVX1_LOC_309/A 0.10fF
C5204 NAND2X1_LOC_538/Y INVX1_LOC_118/A 0.10fF
C5205 INVX1_LOC_18/A NOR2X1_LOC_24/Y 0.04fF
C5206 NOR2X1_LOC_328/Y INVX1_LOC_90/A 2.81fF
C5207 NAND2X1_LOC_477/A INVX1_LOC_144/A 0.01fF
C5208 INVX1_LOC_50/A NOR2X1_LOC_519/Y 0.02fF
C5209 INVX1_LOC_158/A INVX1_LOC_158/Y 0.27fF
C5210 NOR2X1_LOC_667/A INVX1_LOC_140/A 0.10fF
C5211 NOR2X1_LOC_303/Y NOR2X1_LOC_405/A 0.07fF
C5212 NOR2X1_LOC_45/B NAND2X1_LOC_632/B 0.18fF
C5213 NOR2X1_LOC_824/A NOR2X1_LOC_88/Y 0.07fF
C5214 INVX1_LOC_58/A INVX1_LOC_109/A 0.03fF
C5215 INVX1_LOC_248/A INVX1_LOC_140/A 0.20fF
C5216 INVX1_LOC_31/A NAND2X1_LOC_96/A 0.07fF
C5217 INVX1_LOC_95/A INVX1_LOC_71/A 0.03fF
C5218 NAND2X1_LOC_214/B INVX1_LOC_84/A 0.42fF
C5219 INVX1_LOC_206/A NOR2X1_LOC_335/B 0.34fF
C5220 NAND2X1_LOC_338/B NAND2X1_LOC_102/a_36_24# 0.00fF
C5221 NOR2X1_LOC_315/Y INVX1_LOC_6/A 0.28fF
C5222 NOR2X1_LOC_68/A INVX1_LOC_2/Y 1.81fF
C5223 NOR2X1_LOC_632/Y INVX1_LOC_55/Y 0.03fF
C5224 INVX1_LOC_143/A NOR2X1_LOC_74/A 0.01fF
C5225 NOR2X1_LOC_690/A INVX1_LOC_91/A 0.08fF
C5226 INVX1_LOC_135/A NOR2X1_LOC_71/Y 0.01fF
C5227 D_INPUT_1 NAND2X1_LOC_254/Y 0.12fF
C5228 NOR2X1_LOC_346/A NOR2X1_LOC_416/A 0.05fF
C5229 NOR2X1_LOC_32/B NOR2X1_LOC_671/Y 0.13fF
C5230 NOR2X1_LOC_298/Y INVX1_LOC_173/Y 1.91fF
C5231 NOR2X1_LOC_798/A NOR2X1_LOC_691/A 0.00fF
C5232 NOR2X1_LOC_224/Y INVX1_LOC_12/A 0.01fF
C5233 INVX1_LOC_27/A INVX1_LOC_84/A 0.14fF
C5234 NAND2X1_LOC_350/A NOR2X1_LOC_506/Y 0.02fF
C5235 NAND2X1_LOC_597/a_36_24# NOR2X1_LOC_331/B 0.00fF
C5236 NOR2X1_LOC_590/A INVX1_LOC_118/Y 0.02fF
C5237 NOR2X1_LOC_68/A NAND2X1_LOC_129/a_36_24# 0.00fF
C5238 NOR2X1_LOC_737/a_36_216# INVX1_LOC_266/Y 0.01fF
C5239 NOR2X1_LOC_824/A INVX1_LOC_84/A 0.42fF
C5240 NOR2X1_LOC_89/A NOR2X1_LOC_678/A 0.03fF
C5241 INVX1_LOC_219/A INVX1_LOC_90/A 0.01fF
C5242 INVX1_LOC_143/A NOR2X1_LOC_9/Y -0.02fF
C5243 INVX1_LOC_34/A NAND2X1_LOC_642/Y 0.03fF
C5244 NOR2X1_LOC_89/A INVX1_LOC_295/Y 0.01fF
C5245 INVX1_LOC_75/A INVX1_LOC_22/A 0.08fF
C5246 NOR2X1_LOC_690/A INVX1_LOC_11/Y 0.07fF
C5247 NOR2X1_LOC_717/B INVX1_LOC_196/Y 0.03fF
C5248 NOR2X1_LOC_387/A NOR2X1_LOC_505/Y 0.00fF
C5249 NAND2X1_LOC_850/A NAND2X1_LOC_573/A 0.02fF
C5250 INVX1_LOC_271/A INVX1_LOC_15/A 1.98fF
C5251 INVX1_LOC_45/A NOR2X1_LOC_602/B 0.01fF
C5252 INVX1_LOC_135/A NOR2X1_LOC_644/A 0.09fF
C5253 NAND2X1_LOC_63/Y NOR2X1_LOC_81/Y 0.01fF
C5254 INVX1_LOC_10/A NAND2X1_LOC_652/Y 0.02fF
C5255 INVX1_LOC_278/A INVX1_LOC_170/Y 0.00fF
C5256 INVX1_LOC_45/A INVX1_LOC_54/A 0.16fF
C5257 INVX1_LOC_100/Y NAND2X1_LOC_850/Y 0.02fF
C5258 NOR2X1_LOC_68/A NAND2X1_LOC_846/a_36_24# 0.01fF
C5259 INVX1_LOC_270/A INVX1_LOC_94/Y 0.03fF
C5260 NOR2X1_LOC_828/A INVX1_LOC_196/Y 0.06fF
C5261 INVX1_LOC_255/Y NOR2X1_LOC_391/B 0.04fF
C5262 NAND2X1_LOC_333/a_36_24# INVX1_LOC_12/A 0.00fF
C5263 INVX1_LOC_54/Y NOR2X1_LOC_405/A 0.08fF
C5264 NAND2X1_LOC_562/B NOR2X1_LOC_670/Y 0.01fF
C5265 NOR2X1_LOC_350/A INVX1_LOC_117/A 0.02fF
C5266 NAND2X1_LOC_231/Y NAND2X1_LOC_642/Y 0.03fF
C5267 NOR2X1_LOC_91/A NAND2X1_LOC_99/A 0.19fF
C5268 INVX1_LOC_17/A INVX1_LOC_63/A 0.46fF
C5269 INVX1_LOC_182/A INVX1_LOC_313/Y 0.02fF
C5270 INVX1_LOC_89/A INVX1_LOC_31/Y 0.03fF
C5271 INVX1_LOC_21/A INVX1_LOC_42/A 0.17fF
C5272 NOR2X1_LOC_130/A NOR2X1_LOC_74/A 0.07fF
C5273 INVX1_LOC_27/A NAND2X1_LOC_220/B 0.13fF
C5274 INVX1_LOC_207/A NOR2X1_LOC_492/Y 0.06fF
C5275 NAND2X1_LOC_348/A NOR2X1_LOC_130/a_36_216# 0.00fF
C5276 INVX1_LOC_299/A NOR2X1_LOC_633/A 0.02fF
C5277 NOR2X1_LOC_151/Y INVX1_LOC_196/Y 0.02fF
C5278 NAND2X1_LOC_364/A NAND2X1_LOC_656/B 0.01fF
C5279 INVX1_LOC_275/A NOR2X1_LOC_684/Y 0.22fF
C5280 NAND2X1_LOC_579/A INVX1_LOC_284/A 0.02fF
C5281 INVX1_LOC_71/A INVX1_LOC_54/A 0.38fF
C5282 NOR2X1_LOC_434/a_36_216# NOR2X1_LOC_862/B 0.15fF
C5283 INVX1_LOC_23/A NAND2X1_LOC_99/A 0.20fF
C5284 INVX1_LOC_316/A INVX1_LOC_316/Y 0.00fF
C5285 INVX1_LOC_94/Y NOR2X1_LOC_109/Y 0.03fF
C5286 NOR2X1_LOC_68/A NOR2X1_LOC_608/Y 0.05fF
C5287 INVX1_LOC_27/A INVX1_LOC_15/A 7.03fF
C5288 NOR2X1_LOC_781/A NOR2X1_LOC_43/Y 0.02fF
C5289 NOR2X1_LOC_180/B NOR2X1_LOC_188/A 0.18fF
C5290 INVX1_LOC_286/A NOR2X1_LOC_123/B 0.10fF
C5291 NAND2X1_LOC_793/B NOR2X1_LOC_438/Y 0.05fF
C5292 INVX1_LOC_34/A NOR2X1_LOC_271/Y 0.05fF
C5293 GATE_811 NAND2X1_LOC_770/a_36_24# 0.00fF
C5294 INVX1_LOC_48/Y INVX1_LOC_3/Y 0.13fF
C5295 NAND2X1_LOC_227/Y INVX1_LOC_12/A 0.04fF
C5296 NOR2X1_LOC_121/A INVX1_LOC_76/A 0.20fF
C5297 INVX1_LOC_53/A NOR2X1_LOC_858/A 0.00fF
C5298 NAND2X1_LOC_415/a_36_24# NAND2X1_LOC_215/A 0.00fF
C5299 INVX1_LOC_55/A NOR2X1_LOC_89/A 0.01fF
C5300 INVX1_LOC_21/A INVX1_LOC_78/A 0.18fF
C5301 NAND2X1_LOC_361/Y INVX1_LOC_92/A 0.38fF
C5302 INVX1_LOC_22/A NAND2X1_LOC_453/A 0.03fF
C5303 NOR2X1_LOC_551/Y NOR2X1_LOC_564/Y 0.02fF
C5304 NOR2X1_LOC_371/a_36_216# NAND2X1_LOC_254/Y 0.00fF
C5305 INVX1_LOC_61/Y INVX1_LOC_12/A 1.23fF
C5306 NOR2X1_LOC_632/Y NOR2X1_LOC_357/Y 0.01fF
C5307 NOR2X1_LOC_791/A NAND2X1_LOC_773/B -0.01fF
C5308 NOR2X1_LOC_276/Y INVX1_LOC_290/Y 0.00fF
C5309 INVX1_LOC_41/A NOR2X1_LOC_155/A 1.51fF
C5310 INVX1_LOC_286/A INVX1_LOC_102/Y 0.10fF
C5311 NAND2X1_LOC_54/a_36_24# NOR2X1_LOC_536/A 0.00fF
C5312 NAND2X1_LOC_116/A INVX1_LOC_108/A 0.06fF
C5313 INVX1_LOC_249/A INVX1_LOC_84/A 0.29fF
C5314 INVX1_LOC_50/Y NOR2X1_LOC_727/B 0.16fF
C5315 INVX1_LOC_234/A NOR2X1_LOC_825/Y 0.10fF
C5316 INVX1_LOC_21/A INVX1_LOC_288/A 0.06fF
C5317 INVX1_LOC_45/A NAND2X1_LOC_807/B 0.01fF
C5318 NOR2X1_LOC_454/Y NOR2X1_LOC_45/a_36_216# 0.01fF
C5319 NAND2X1_LOC_466/A NAND2X1_LOC_798/B 0.05fF
C5320 INVX1_LOC_21/A NOR2X1_LOC_65/B 0.08fF
C5321 INVX1_LOC_290/A INVX1_LOC_117/A 0.07fF
C5322 NOR2X1_LOC_45/B NOR2X1_LOC_163/Y 1.20fF
C5323 NOR2X1_LOC_510/Y INVX1_LOC_57/A 0.03fF
C5324 INVX1_LOC_45/A NOR2X1_LOC_48/B 0.07fF
C5325 NOR2X1_LOC_338/Y INVX1_LOC_109/A 0.03fF
C5326 INVX1_LOC_288/Y NOR2X1_LOC_454/Y 0.05fF
C5327 INVX1_LOC_58/A NAND2X1_LOC_794/B 0.03fF
C5328 INVX1_LOC_136/A INVX1_LOC_290/Y 0.09fF
C5329 INVX1_LOC_269/A INVX1_LOC_26/A 0.10fF
C5330 INVX1_LOC_255/Y INVX1_LOC_280/A 0.07fF
C5331 NOR2X1_LOC_207/A NOR2X1_LOC_155/A 0.04fF
C5332 NAND2X1_LOC_122/a_36_24# INVX1_LOC_123/Y 0.00fF
C5333 INVX1_LOC_95/A INVX1_LOC_102/Y 0.24fF
C5334 INVX1_LOC_140/A INVX1_LOC_304/A 0.11fF
C5335 INVX1_LOC_53/A NOR2X1_LOC_406/A 0.03fF
C5336 INVX1_LOC_18/A NOR2X1_LOC_490/a_36_216# 0.00fF
C5337 INVX1_LOC_35/A NOR2X1_LOC_434/Y 0.54fF
C5338 NOR2X1_LOC_272/Y NAND2X1_LOC_860/A 0.19fF
C5339 NOR2X1_LOC_690/A INVX1_LOC_203/A 0.03fF
C5340 NOR2X1_LOC_664/Y INVX1_LOC_84/A 0.04fF
C5341 INVX1_LOC_77/A NAND2X1_LOC_74/B 0.10fF
C5342 INVX1_LOC_108/Y INVX1_LOC_27/A 0.03fF
C5343 INVX1_LOC_11/A NOR2X1_LOC_318/A 0.01fF
C5344 INVX1_LOC_58/A INVX1_LOC_48/Y 0.02fF
C5345 NOR2X1_LOC_328/Y NOR2X1_LOC_51/A 0.01fF
C5346 INVX1_LOC_71/A NAND2X1_LOC_807/B 0.03fF
C5347 INPUT_0 NAND2X1_LOC_642/Y 2.63fF
C5348 INVX1_LOC_21/A INVX1_LOC_152/Y 0.08fF
C5349 INVX1_LOC_278/A INVX1_LOC_27/A 0.10fF
C5350 INVX1_LOC_105/A INVX1_LOC_12/A 0.09fF
C5351 INVX1_LOC_45/A NAND2X1_LOC_3/B 0.02fF
C5352 INVX1_LOC_96/A INVX1_LOC_78/Y 0.17fF
C5353 INVX1_LOC_223/A NAND2X1_LOC_647/B 0.03fF
C5354 NOR2X1_LOC_403/B NAND2X1_LOC_254/Y 0.00fF
C5355 INVX1_LOC_39/A NAND2X1_LOC_569/B 0.04fF
C5356 NOR2X1_LOC_361/B INVX1_LOC_57/A 0.05fF
C5357 INVX1_LOC_206/A INVX1_LOC_84/A 0.38fF
C5358 INVX1_LOC_90/A INVX1_LOC_33/Y 0.07fF
C5359 NAND2X1_LOC_570/Y INVX1_LOC_84/A 0.02fF
C5360 NOR2X1_LOC_380/Y VDD 0.61fF
C5361 NOR2X1_LOC_78/A INVX1_LOC_125/Y 0.01fF
C5362 NAND2X1_LOC_555/Y NAND2X1_LOC_223/B 0.03fF
C5363 NOR2X1_LOC_598/B INVX1_LOC_24/Y 0.48fF
C5364 INVX1_LOC_36/A INVX1_LOC_94/Y 0.67fF
C5365 INVX1_LOC_248/Y NAND2X1_LOC_794/B 0.20fF
C5366 INVX1_LOC_258/Y INVX1_LOC_5/A 0.03fF
C5367 INVX1_LOC_31/A NAND2X1_LOC_99/A 0.00fF
C5368 NAND2X1_LOC_182/A INVX1_LOC_29/A 0.03fF
C5369 NOR2X1_LOC_92/Y NAND2X1_LOC_725/A 0.19fF
C5370 NAND2X1_LOC_174/a_36_24# INVX1_LOC_12/A 0.00fF
C5371 INVX1_LOC_104/A INVX1_LOC_29/A 0.17fF
C5372 NAND2X1_LOC_787/A NOR2X1_LOC_438/a_36_216# 0.00fF
C5373 D_INPUT_7 NOR2X1_LOC_36/A 0.17fF
C5374 NAND2X1_LOC_354/Y INVX1_LOC_78/A 0.04fF
C5375 INVX1_LOC_249/A INVX1_LOC_15/A 0.00fF
C5376 NAND2X1_LOC_141/A NAND2X1_LOC_82/Y 0.04fF
C5377 NOR2X1_LOC_428/a_36_216# INVX1_LOC_23/A 0.02fF
C5378 INVX1_LOC_135/A NAND2X1_LOC_243/Y 0.03fF
C5379 NOR2X1_LOC_134/Y NAND2X1_LOC_464/B 0.03fF
C5380 NOR2X1_LOC_709/A NAND2X1_LOC_63/Y 0.08fF
C5381 NOR2X1_LOC_582/Y INVX1_LOC_78/A 0.00fF
C5382 INVX1_LOC_6/Y INVX1_LOC_15/A 0.02fF
C5383 INVX1_LOC_50/A NAND2X1_LOC_733/Y 0.11fF
C5384 INVX1_LOC_11/A NOR2X1_LOC_678/A 0.03fF
C5385 NOR2X1_LOC_239/a_36_216# INVX1_LOC_26/Y 0.00fF
C5386 INVX1_LOC_11/A INVX1_LOC_295/Y 0.09fF
C5387 INVX1_LOC_16/A NAND2X1_LOC_475/Y 0.39fF
C5388 NAND2X1_LOC_649/B NAND2X1_LOC_642/Y 0.03fF
C5389 INVX1_LOC_145/A INVX1_LOC_94/Y 0.04fF
C5390 INVX1_LOC_36/A INVX1_LOC_181/A 0.62fF
C5391 INVX1_LOC_137/A INVX1_LOC_84/A 0.01fF
C5392 NOR2X1_LOC_778/Y NOR2X1_LOC_383/B 0.20fF
C5393 INVX1_LOC_36/A INVX1_LOC_296/A 0.09fF
C5394 NOR2X1_LOC_303/a_36_216# INVX1_LOC_38/A 0.02fF
C5395 NAND2X1_LOC_573/A NAND2X1_LOC_286/a_36_24# 0.00fF
C5396 NAND2X1_LOC_577/A INVX1_LOC_23/A 0.09fF
C5397 INVX1_LOC_49/A NOR2X1_LOC_334/Y 5.96fF
C5398 NAND2X1_LOC_579/A NOR2X1_LOC_384/A 0.02fF
C5399 INVX1_LOC_201/A NAND2X1_LOC_8/a_36_24# 0.00fF
C5400 INVX1_LOC_63/Y INVX1_LOC_4/A 0.10fF
C5401 D_GATE_366 NOR2X1_LOC_364/A 0.00fF
C5402 NOR2X1_LOC_302/B INVX1_LOC_186/Y 0.03fF
C5403 INVX1_LOC_234/A INVX1_LOC_84/A 0.27fF
C5404 INVX1_LOC_50/A INVX1_LOC_217/A 0.10fF
C5405 NOR2X1_LOC_468/Y NOR2X1_LOC_440/B 0.19fF
C5406 INPUT_0 NOR2X1_LOC_271/Y 0.04fF
C5407 NOR2X1_LOC_245/a_36_216# INVX1_LOC_285/A 0.00fF
C5408 INVX1_LOC_62/Y NOR2X1_LOC_720/A 0.02fF
C5409 NAND2X1_LOC_654/B INVX1_LOC_92/A 0.02fF
C5410 INVX1_LOC_71/A NOR2X1_LOC_438/Y 0.01fF
C5411 NOR2X1_LOC_667/A INVX1_LOC_42/A 0.10fF
C5412 NOR2X1_LOC_356/A NOR2X1_LOC_197/B 0.10fF
C5413 NOR2X1_LOC_84/Y INVX1_LOC_3/Y 0.12fF
C5414 INVX1_LOC_248/A INVX1_LOC_42/A 0.07fF
C5415 NOR2X1_LOC_264/Y INVX1_LOC_4/Y 0.02fF
C5416 NOR2X1_LOC_356/A NAND2X1_LOC_237/a_36_24# 0.01fF
C5417 INVX1_LOC_12/Y NOR2X1_LOC_269/Y 0.02fF
C5418 NOR2X1_LOC_333/A NOR2X1_LOC_814/A 0.02fF
C5419 NAND2X1_LOC_570/Y INVX1_LOC_15/A 0.01fF
C5420 NOR2X1_LOC_780/B NOR2X1_LOC_796/B 0.01fF
C5421 INVX1_LOC_39/A NOR2X1_LOC_530/Y 0.01fF
C5422 NOR2X1_LOC_20/a_36_216# NOR2X1_LOC_629/Y 0.00fF
C5423 INVX1_LOC_64/A NAND2X1_LOC_154/Y 0.02fF
C5424 INVX1_LOC_288/Y INVX1_LOC_77/A 0.01fF
C5425 NOR2X1_LOC_334/A INVX1_LOC_9/A 0.02fF
C5426 NAND2X1_LOC_858/B INVX1_LOC_185/A 0.03fF
C5427 NAND2X1_LOC_640/Y INVX1_LOC_183/A 0.00fF
C5428 D_INPUT_1 INVX1_LOC_314/Y 0.04fF
C5429 INVX1_LOC_2/A NOR2X1_LOC_334/Y 0.36fF
C5430 INVX1_LOC_50/A NAND2X1_LOC_787/B 0.03fF
C5431 INVX1_LOC_298/Y INVX1_LOC_104/A 0.15fF
C5432 NOR2X1_LOC_392/B INVX1_LOC_23/Y 0.10fF
C5433 INVX1_LOC_28/A NAND2X1_LOC_475/Y 0.10fF
C5434 NOR2X1_LOC_74/A NOR2X1_LOC_197/B 0.01fF
C5435 NOR2X1_LOC_19/B INVX1_LOC_84/A 0.26fF
C5436 INVX1_LOC_190/A NAND2X1_LOC_74/B 0.00fF
C5437 NAND2X1_LOC_569/B INVX1_LOC_61/A 0.21fF
C5438 NOR2X1_LOC_337/Y INVX1_LOC_274/A 0.08fF
C5439 INVX1_LOC_95/Y NOR2X1_LOC_536/A 0.07fF
C5440 NOR2X1_LOC_112/B NOR2X1_LOC_243/B 0.01fF
C5441 NOR2X1_LOC_52/B NOR2X1_LOC_318/A 0.00fF
C5442 INVX1_LOC_214/A INVX1_LOC_78/A 0.01fF
C5443 NOR2X1_LOC_667/A INVX1_LOC_78/A 0.21fF
C5444 INVX1_LOC_35/A NOR2X1_LOC_274/Y 0.01fF
C5445 NOR2X1_LOC_9/Y NOR2X1_LOC_197/B 0.04fF
C5446 NAND2X1_LOC_725/A NAND2X1_LOC_837/Y 0.10fF
C5447 INVX1_LOC_248/A INVX1_LOC_78/A 0.03fF
C5448 NOR2X1_LOC_632/Y INVX1_LOC_32/A 0.03fF
C5449 NAND2X1_LOC_149/Y INVX1_LOC_30/A 1.21fF
C5450 INVX1_LOC_223/Y INVX1_LOC_18/A 0.03fF
C5451 INVX1_LOC_144/A NOR2X1_LOC_435/B 0.02fF
C5452 NOR2X1_LOC_433/A NOR2X1_LOC_678/A 0.04fF
C5453 INVX1_LOC_21/A NOR2X1_LOC_554/B 0.10fF
C5454 INVX1_LOC_172/Y INVX1_LOC_253/A 0.00fF
C5455 NOR2X1_LOC_796/B NOR2X1_LOC_803/B 0.02fF
C5456 NOR2X1_LOC_180/Y NOR2X1_LOC_383/B 0.09fF
C5457 INVX1_LOC_41/A NOR2X1_LOC_598/B 0.23fF
C5458 NOR2X1_LOC_750/Y INVX1_LOC_34/A 0.03fF
C5459 NAND2X1_LOC_763/B NAND2X1_LOC_149/Y 0.02fF
C5460 INVX1_LOC_55/A INVX1_LOC_11/A 0.02fF
C5461 NAND2X1_LOC_850/A NAND2X1_LOC_81/B 0.03fF
C5462 NOR2X1_LOC_593/Y NOR2X1_LOC_678/A 0.06fF
C5463 NOR2X1_LOC_555/a_36_216# INVX1_LOC_179/A 0.00fF
C5464 INVX1_LOC_136/A NOR2X1_LOC_454/Y 0.01fF
C5465 INVX1_LOC_234/A INVX1_LOC_15/A 0.07fF
C5466 INVX1_LOC_75/A INVX1_LOC_186/Y 0.48fF
C5467 INVX1_LOC_268/A NAND2X1_LOC_470/B 0.02fF
C5468 INVX1_LOC_41/A INVX1_LOC_51/A 0.01fF
C5469 NOR2X1_LOC_528/Y NOR2X1_LOC_88/Y 0.07fF
C5470 NAND2X1_LOC_579/A INVX1_LOC_72/A 0.07fF
C5471 INVX1_LOC_177/A INVX1_LOC_57/A 0.00fF
C5472 NOR2X1_LOC_405/A NAND2X1_LOC_656/B 0.01fF
C5473 NAND2X1_LOC_9/Y NOR2X1_LOC_720/B 0.01fF
C5474 INVX1_LOC_64/A INVX1_LOC_63/Y 0.43fF
C5475 NAND2X1_LOC_652/Y INVX1_LOC_12/A 0.03fF
C5476 INVX1_LOC_313/Y NOR2X1_LOC_850/B 0.07fF
C5477 INVX1_LOC_95/Y NAND2X1_LOC_93/B 0.17fF
C5478 NOR2X1_LOC_655/B INVX1_LOC_224/Y 0.05fF
C5479 NOR2X1_LOC_498/Y NAND2X1_LOC_725/A 0.10fF
C5480 NOR2X1_LOC_67/A NOR2X1_LOC_646/B 0.00fF
C5481 INVX1_LOC_144/Y NOR2X1_LOC_654/A 0.22fF
C5482 NOR2X1_LOC_497/Y NAND2X1_LOC_254/Y 0.01fF
C5483 INVX1_LOC_233/Y NAND2X1_LOC_735/a_36_24# 0.01fF
C5484 INVX1_LOC_21/A NOR2X1_LOC_152/Y 0.06fF
C5485 NAND2X1_LOC_347/B INVX1_LOC_181/Y 0.00fF
C5486 INVX1_LOC_135/A INVX1_LOC_21/Y 0.01fF
C5487 NOR2X1_LOC_78/B NOR2X1_LOC_858/A 0.04fF
C5488 INVX1_LOC_34/A INVX1_LOC_204/Y 0.07fF
C5489 NOR2X1_LOC_528/Y INVX1_LOC_84/A 0.01fF
C5490 INVX1_LOC_33/Y INVX1_LOC_38/A 0.03fF
C5491 NOR2X1_LOC_388/a_36_216# NOR2X1_LOC_383/B 0.00fF
C5492 NAND2X1_LOC_35/Y NAND2X1_LOC_465/Y 0.03fF
C5493 INVX1_LOC_45/A NAND2X1_LOC_350/A 0.07fF
C5494 INVX1_LOC_269/A NAND2X1_LOC_371/a_36_24# 0.00fF
C5495 NAND2X1_LOC_35/Y NOR2X1_LOC_234/Y 0.02fF
C5496 VDD INVX1_LOC_274/A 0.24fF
C5497 NOR2X1_LOC_468/Y INVX1_LOC_41/Y 0.00fF
C5498 NOR2X1_LOC_242/A NAND2X1_LOC_361/Y 0.07fF
C5499 INVX1_LOC_36/A INVX1_LOC_293/A 0.04fF
C5500 NOR2X1_LOC_222/Y INVX1_LOC_23/A 0.08fF
C5501 NAND2X1_LOC_67/Y NOR2X1_LOC_759/Y 0.09fF
C5502 NOR2X1_LOC_240/Y NOR2X1_LOC_243/Y 0.19fF
C5503 INVX1_LOC_64/A NOR2X1_LOC_175/A 0.03fF
C5504 NAND2X1_LOC_577/A INVX1_LOC_31/A 0.09fF
C5505 INVX1_LOC_225/A NOR2X1_LOC_220/B 0.01fF
C5506 NAND2X1_LOC_489/a_36_24# NAND2X1_LOC_244/A 0.00fF
C5507 NOR2X1_LOC_19/B INVX1_LOC_15/A 0.07fF
C5508 NOR2X1_LOC_135/Y INVX1_LOC_32/A 0.00fF
C5509 INVX1_LOC_45/A NOR2X1_LOC_441/Y 0.02fF
C5510 NOR2X1_LOC_844/A NOR2X1_LOC_849/A 0.53fF
C5511 INVX1_LOC_206/Y INVX1_LOC_29/A 0.06fF
C5512 NAND2X1_LOC_600/a_36_24# NOR2X1_LOC_536/A 0.00fF
C5513 NOR2X1_LOC_186/Y NAND2X1_LOC_759/a_36_24# 0.00fF
C5514 INVX1_LOC_95/Y INVX1_LOC_3/A 0.03fF
C5515 INVX1_LOC_61/A NOR2X1_LOC_530/Y 0.01fF
C5516 INVX1_LOC_135/A INVX1_LOC_16/Y 0.01fF
C5517 NOR2X1_LOC_620/Y INVX1_LOC_1/A 0.01fF
C5518 NOR2X1_LOC_160/B NOR2X1_LOC_360/Y 0.07fF
C5519 NOR2X1_LOC_846/Y NOR2X1_LOC_87/B 0.00fF
C5520 NOR2X1_LOC_78/A INVX1_LOC_19/A 0.25fF
C5521 NOR2X1_LOC_813/Y NAND2X1_LOC_243/Y 0.02fF
C5522 INVX1_LOC_58/A INVX1_LOC_290/A 0.12fF
C5523 NOR2X1_LOC_798/A NOR2X1_LOC_174/a_36_216# 0.00fF
C5524 INVX1_LOC_245/Y INVX1_LOC_24/A 0.00fF
C5525 INVX1_LOC_36/A NOR2X1_LOC_524/Y 0.04fF
C5526 NOR2X1_LOC_813/Y INVX1_LOC_89/Y 0.03fF
C5527 VDD NOR2X1_LOC_820/Y 0.19fF
C5528 NAND2X1_LOC_787/A INVX1_LOC_16/A 0.04fF
C5529 NOR2X1_LOC_331/B INVX1_LOC_54/A 0.26fF
C5530 INVX1_LOC_220/Y INVX1_LOC_23/A 0.03fF
C5531 NAND2X1_LOC_573/A INVX1_LOC_57/A 0.02fF
C5532 INVX1_LOC_39/A NOR2X1_LOC_709/A 0.03fF
C5533 NOR2X1_LOC_91/A NOR2X1_LOC_380/A 0.08fF
C5534 NOR2X1_LOC_785/Y INVX1_LOC_57/A 0.11fF
C5535 NAND2X1_LOC_573/Y NAND2X1_LOC_759/a_36_24# 0.01fF
C5536 INVX1_LOC_179/A INVX1_LOC_281/A 0.00fF
C5537 NOR2X1_LOC_15/Y INVX1_LOC_88/Y 0.01fF
C5538 INVX1_LOC_50/A NAND2X1_LOC_808/A 0.00fF
C5539 NAND2X1_LOC_724/A NAND2X1_LOC_811/Y 0.02fF
C5540 INVX1_LOC_66/A INVX1_LOC_270/A 0.03fF
C5541 NOR2X1_LOC_600/Y INVX1_LOC_29/A 0.01fF
C5542 INVX1_LOC_36/Y NOR2X1_LOC_814/A 0.03fF
C5543 NAND2X1_LOC_656/A INVX1_LOC_31/A 0.25fF
C5544 NOR2X1_LOC_443/Y INVX1_LOC_148/Y 0.27fF
C5545 INVX1_LOC_224/Y NOR2X1_LOC_99/B 0.04fF
C5546 INVX1_LOC_280/A NOR2X1_LOC_61/A 0.00fF
C5547 INVX1_LOC_135/A NAND2X1_LOC_205/A 0.01fF
C5548 INVX1_LOC_1/A NOR2X1_LOC_731/A 0.03fF
C5549 INVX1_LOC_77/A NOR2X1_LOC_276/Y 0.11fF
C5550 NOR2X1_LOC_657/Y INVX1_LOC_159/A 0.02fF
C5551 NOR2X1_LOC_598/B INVX1_LOC_121/A 0.02fF
C5552 NOR2X1_LOC_441/Y INVX1_LOC_71/A 0.00fF
C5553 INVX1_LOC_207/A NAND2X1_LOC_550/A 0.01fF
C5554 NAND2X1_LOC_51/B INVX1_LOC_78/A 0.92fF
C5555 NAND2X1_LOC_464/A INVX1_LOC_19/A 0.02fF
C5556 INPUT_1 NAND2X1_LOC_464/B 0.08fF
C5557 NOR2X1_LOC_91/A NOR2X1_LOC_329/B 0.10fF
C5558 NAND2X1_LOC_705/Y NAND2X1_LOC_374/Y 0.10fF
C5559 INVX1_LOC_5/A NOR2X1_LOC_589/A 0.14fF
C5560 NOR2X1_LOC_791/Y INVX1_LOC_16/A 0.00fF
C5561 NOR2X1_LOC_294/Y NOR2X1_LOC_860/B 0.01fF
C5562 INVX1_LOC_178/A NOR2X1_LOC_418/Y 0.40fF
C5563 INVX1_LOC_304/A INVX1_LOC_42/A 0.03fF
C5564 INVX1_LOC_311/A INVX1_LOC_78/A 0.03fF
C5565 NOR2X1_LOC_592/B INVX1_LOC_54/A 0.07fF
C5566 NOR2X1_LOC_742/A NOR2X1_LOC_302/A 0.04fF
C5567 NAND2X1_LOC_725/A NOR2X1_LOC_299/Y 0.07fF
C5568 INVX1_LOC_175/Y NOR2X1_LOC_476/B 0.71fF
C5569 INVX1_LOC_174/A NOR2X1_LOC_377/Y 0.02fF
C5570 NOR2X1_LOC_565/A NOR2X1_LOC_550/B 0.03fF
C5571 INVX1_LOC_75/A NOR2X1_LOC_843/B 0.01fF
C5572 NAND2X1_LOC_348/A NOR2X1_LOC_342/B 0.28fF
C5573 INVX1_LOC_163/A INVX1_LOC_84/Y 0.04fF
C5574 INVX1_LOC_35/A NAND2X1_LOC_45/Y 0.01fF
C5575 NAND2X1_LOC_181/Y INVX1_LOC_1/A 0.64fF
C5576 NOR2X1_LOC_670/Y INVX1_LOC_42/A 0.02fF
C5577 INVX1_LOC_136/A INVX1_LOC_77/A 0.11fF
C5578 NOR2X1_LOC_329/B INVX1_LOC_23/A 4.64fF
C5579 NAND2X1_LOC_656/A INVX1_LOC_111/A 0.04fF
C5580 VDD NOR2X1_LOC_33/B -0.00fF
C5581 NOR2X1_LOC_655/B NOR2X1_LOC_103/Y 0.10fF
C5582 NOR2X1_LOC_391/B INVX1_LOC_16/Y 0.06fF
C5583 INVX1_LOC_287/A INVX1_LOC_75/A 0.00fF
C5584 NOR2X1_LOC_60/Y INVX1_LOC_19/A 0.06fF
C5585 NOR2X1_LOC_623/a_36_216# INVX1_LOC_30/A 0.00fF
C5586 NOR2X1_LOC_545/B NOR2X1_LOC_620/A 0.05fF
C5587 INVX1_LOC_45/A NOR2X1_LOC_142/Y 0.01fF
C5588 NAND2X1_LOC_787/A INVX1_LOC_28/A 0.03fF
C5589 NOR2X1_LOC_45/Y INVX1_LOC_266/Y 0.01fF
C5590 INVX1_LOC_104/A NOR2X1_LOC_703/a_36_216# 0.00fF
C5591 D_INPUT_4 INVX1_LOC_23/A 0.01fF
C5592 NOR2X1_LOC_565/a_36_216# NOR2X1_LOC_383/B 0.00fF
C5593 NAND2X1_LOC_714/B NOR2X1_LOC_561/Y 0.01fF
C5594 INVX1_LOC_298/A INVX1_LOC_89/A 0.00fF
C5595 NOR2X1_LOC_690/A NOR2X1_LOC_372/Y 0.01fF
C5596 INVX1_LOC_265/A INVX1_LOC_57/Y 0.41fF
C5597 INVX1_LOC_6/A NAND2X1_LOC_99/A 0.09fF
C5598 NOR2X1_LOC_341/a_36_216# NOR2X1_LOC_350/A 0.02fF
C5599 NOR2X1_LOC_590/A NOR2X1_LOC_520/A 0.01fF
C5600 INVX1_LOC_114/Y INVX1_LOC_117/A 0.03fF
C5601 INVX1_LOC_14/A INVX1_LOC_137/Y 0.00fF
C5602 INVX1_LOC_21/A NAND2X1_LOC_861/Y 0.07fF
C5603 INVX1_LOC_36/A NOR2X1_LOC_315/Y 0.07fF
C5604 NOR2X1_LOC_817/Y NAND2X1_LOC_820/a_36_24# 0.00fF
C5605 INVX1_LOC_17/A INVX1_LOC_1/Y 0.03fF
C5606 INVX1_LOC_194/A INVX1_LOC_195/A 0.01fF
C5607 NOR2X1_LOC_859/A NOR2X1_LOC_844/A 0.02fF
C5608 INVX1_LOC_285/Y INVX1_LOC_57/A 0.74fF
C5609 INVX1_LOC_247/Y INVX1_LOC_104/A 0.01fF
C5610 INVX1_LOC_304/A INVX1_LOC_78/A 0.07fF
C5611 NOR2X1_LOC_15/Y NAND2X1_LOC_656/Y 0.20fF
C5612 NOR2X1_LOC_78/A INVX1_LOC_26/Y 0.09fF
C5613 NOR2X1_LOC_45/B NOR2X1_LOC_693/Y 0.09fF
C5614 NOR2X1_LOC_307/A NOR2X1_LOC_687/Y 0.03fF
C5615 INVX1_LOC_46/Y NAND2X1_LOC_206/Y 0.01fF
C5616 NAND2X1_LOC_74/B INVX1_LOC_9/A 0.28fF
C5617 INVX1_LOC_136/A INVX1_LOC_124/A 0.04fF
C5618 NOR2X1_LOC_216/B INVX1_LOC_84/A 0.07fF
C5619 INVX1_LOC_24/A NOR2X1_LOC_121/Y 0.01fF
C5620 NAND2X1_LOC_112/Y INVX1_LOC_161/Y 0.01fF
C5621 NAND2X1_LOC_806/a_36_24# NOR2X1_LOC_536/A 0.00fF
C5622 NAND2X1_LOC_207/Y INVX1_LOC_9/A 0.02fF
C5623 INVX1_LOC_45/A NOR2X1_LOC_655/B 0.69fF
C5624 INVX1_LOC_213/Y INVX1_LOC_198/Y 0.01fF
C5625 NOR2X1_LOC_142/Y INVX1_LOC_71/A 0.10fF
C5626 NOR2X1_LOC_589/A NAND2X1_LOC_337/B 0.07fF
C5627 NOR2X1_LOC_655/B NOR2X1_LOC_568/A 0.64fF
C5628 INVX1_LOC_119/A NOR2X1_LOC_637/A 0.03fF
C5629 INVX1_LOC_141/Y NAND2X1_LOC_840/B 0.00fF
C5630 NOR2X1_LOC_405/A NAND2X1_LOC_286/B 0.01fF
C5631 INVX1_LOC_46/Y NAND2X1_LOC_773/B 0.02fF
C5632 NOR2X1_LOC_162/Y INVX1_LOC_49/A 0.02fF
C5633 INVX1_LOC_117/A NOR2X1_LOC_467/A 0.03fF
C5634 NAND2X1_LOC_536/a_36_24# NOR2X1_LOC_593/Y 0.00fF
C5635 INVX1_LOC_14/A INVX1_LOC_183/Y 0.01fF
C5636 NOR2X1_LOC_817/Y INVX1_LOC_135/A 0.47fF
C5637 NOR2X1_LOC_778/A NOR2X1_LOC_778/B 0.21fF
C5638 INVX1_LOC_72/A INVX1_LOC_43/A 0.01fF
C5639 INVX1_LOC_58/A NOR2X1_LOC_41/a_36_216# 0.00fF
C5640 INVX1_LOC_230/Y NOR2X1_LOC_391/A 0.70fF
C5641 NAND2X1_LOC_734/B INVX1_LOC_172/A 0.27fF
C5642 INVX1_LOC_30/A INVX1_LOC_16/A 1.31fF
C5643 NOR2X1_LOC_388/Y NOR2X1_LOC_570/B 0.36fF
C5644 NOR2X1_LOC_237/Y NOR2X1_LOC_315/Y 0.41fF
C5645 NOR2X1_LOC_337/A INVX1_LOC_50/Y 0.03fF
C5646 NOR2X1_LOC_496/Y INVX1_LOC_282/A 0.01fF
C5647 INVX1_LOC_278/A NOR2X1_LOC_528/Y 0.12fF
C5648 INVX1_LOC_22/A NOR2X1_LOC_274/B 0.07fF
C5649 NOR2X1_LOC_82/A NOR2X1_LOC_72/a_36_216# 0.00fF
C5650 INVX1_LOC_18/A INVX1_LOC_25/Y 0.03fF
C5651 NAND2X1_LOC_866/A NOR2X1_LOC_822/Y 0.06fF
C5652 INVX1_LOC_226/Y NOR2X1_LOC_791/B 0.03fF
C5653 NOR2X1_LOC_655/B INVX1_LOC_71/A 0.01fF
C5654 INVX1_LOC_208/A NOR2X1_LOC_360/Y 0.10fF
C5655 INVX1_LOC_57/A NOR2X1_LOC_137/B 0.11fF
C5656 INVX1_LOC_51/Y NOR2X1_LOC_849/A 0.02fF
C5657 NAND2X1_LOC_214/B INVX1_LOC_123/A 0.39fF
C5658 INVX1_LOC_214/A NOR2X1_LOC_152/Y 0.10fF
C5659 NOR2X1_LOC_309/Y INVX1_LOC_162/A 0.02fF
C5660 NAND2X1_LOC_388/a_36_24# INVX1_LOC_30/A 0.00fF
C5661 INVX1_LOC_2/A INVX1_LOC_209/Y 0.03fF
C5662 NOR2X1_LOC_759/Y NOR2X1_LOC_131/a_36_216# 0.00fF
C5663 INVX1_LOC_18/A NOR2X1_LOC_302/B 0.01fF
C5664 NOR2X1_LOC_221/a_36_216# INVX1_LOC_91/A 0.00fF
C5665 INVX1_LOC_12/Y INVX1_LOC_26/A 0.10fF
C5666 NOR2X1_LOC_667/A NOR2X1_LOC_152/Y 0.18fF
C5667 NOR2X1_LOC_590/A NOR2X1_LOC_333/A 0.01fF
C5668 NOR2X1_LOC_497/a_36_216# INVX1_LOC_20/A 0.00fF
C5669 NOR2X1_LOC_219/B INVX1_LOC_96/Y 0.03fF
C5670 NOR2X1_LOC_601/Y NOR2X1_LOC_678/A 0.01fF
C5671 INVX1_LOC_57/A NAND2X1_LOC_267/B 0.01fF
C5672 NOR2X1_LOC_433/A NOR2X1_LOC_191/A 0.02fF
C5673 INVX1_LOC_45/A NOR2X1_LOC_99/B 0.11fF
C5674 NAND2X1_LOC_361/Y NOR2X1_LOC_78/B 2.25fF
C5675 INVX1_LOC_27/A INVX1_LOC_123/A 0.02fF
C5676 NAND2X1_LOC_537/a_36_24# NOR2X1_LOC_385/Y 0.00fF
C5677 INVX1_LOC_22/Y INVX1_LOC_65/Y 0.02fF
C5678 INVX1_LOC_200/Y INVX1_LOC_46/A 0.80fF
C5679 INVX1_LOC_49/A INVX1_LOC_218/A 0.01fF
C5680 NOR2X1_LOC_15/Y NAND2X1_LOC_622/B 0.38fF
C5681 NOR2X1_LOC_690/A NAND2X1_LOC_374/Y 0.06fF
C5682 NOR2X1_LOC_48/a_36_216# NOR2X1_LOC_48/Y 0.00fF
C5683 INVX1_LOC_24/A NAND2X1_LOC_660/Y 0.10fF
C5684 INVX1_LOC_102/A INVX1_LOC_265/Y 0.01fF
C5685 INVX1_LOC_2/A NOR2X1_LOC_718/B 0.01fF
C5686 NAND2X1_LOC_363/B NOR2X1_LOC_35/Y 0.10fF
C5687 INVX1_LOC_280/A INVX1_LOC_16/Y 0.01fF
C5688 INVX1_LOC_269/A NOR2X1_LOC_20/a_36_216# 0.00fF
C5689 INVX1_LOC_174/A INVX1_LOC_140/A 0.31fF
C5690 NOR2X1_LOC_273/Y NOR2X1_LOC_561/Y 0.01fF
C5691 NOR2X1_LOC_160/B NOR2X1_LOC_567/B 0.07fF
C5692 NOR2X1_LOC_833/Y INVX1_LOC_213/A 0.01fF
C5693 NOR2X1_LOC_123/a_36_216# INVX1_LOC_306/Y 0.00fF
C5694 NAND2X1_LOC_477/A NAND2X1_LOC_660/A 0.12fF
C5695 NOR2X1_LOC_471/Y NOR2X1_LOC_742/A 0.02fF
C5696 INVX1_LOC_90/A NAND2X1_LOC_741/B 0.06fF
C5697 NOR2X1_LOC_577/Y INVX1_LOC_22/A 2.63fF
C5698 NOR2X1_LOC_329/B INVX1_LOC_31/A 0.07fF
C5699 INVX1_LOC_177/Y NAND2X1_LOC_140/A 0.01fF
C5700 NOR2X1_LOC_468/Y NOR2X1_LOC_368/a_36_216# 0.00fF
C5701 NOR2X1_LOC_158/B INVX1_LOC_117/Y 0.12fF
C5702 NAND2X1_LOC_811/Y NAND2X1_LOC_852/Y 0.06fF
C5703 NOR2X1_LOC_857/A NOR2X1_LOC_634/Y 0.00fF
C5704 NOR2X1_LOC_192/A NAND2X1_LOC_474/Y 0.02fF
C5705 NOR2X1_LOC_255/Y INVX1_LOC_12/Y 0.02fF
C5706 INVX1_LOC_202/A NOR2X1_LOC_561/Y 0.10fF
C5707 NAND2X1_LOC_93/B INVX1_LOC_271/Y 0.23fF
C5708 NOR2X1_LOC_376/A INVX1_LOC_91/A 0.01fF
C5709 INVX1_LOC_25/A INVX1_LOC_117/A 0.05fF
C5710 NOR2X1_LOC_817/Y NOR2X1_LOC_391/B 0.50fF
C5711 NOR2X1_LOC_515/a_36_216# INVX1_LOC_216/A 0.02fF
C5712 INVX1_LOC_14/A NOR2X1_LOC_114/A 0.00fF
C5713 INVX1_LOC_28/A INVX1_LOC_30/A 1.17fF
C5714 INVX1_LOC_81/A INVX1_LOC_10/A 0.03fF
C5715 NAND2X1_LOC_717/Y NAND2X1_LOC_722/A 0.07fF
C5716 INVX1_LOC_276/A INVX1_LOC_236/A 0.19fF
C5717 D_INPUT_0 INVX1_LOC_24/A 0.15fF
C5718 INVX1_LOC_5/A INVX1_LOC_20/A 1.70fF
C5719 INVX1_LOC_45/A INVX1_LOC_182/A 0.07fF
C5720 NOR2X1_LOC_821/Y NAND2X1_LOC_852/Y 0.36fF
C5721 INVX1_LOC_13/A NOR2X1_LOC_520/B 0.46fF
C5722 NOR2X1_LOC_278/Y NOR2X1_LOC_743/Y 0.70fF
C5723 NAND2X1_LOC_291/B NOR2X1_LOC_777/B 0.06fF
C5724 NOR2X1_LOC_176/Y NAND2X1_LOC_793/B 0.04fF
C5725 INVX1_LOC_280/A NAND2X1_LOC_205/A 0.02fF
C5726 INVX1_LOC_5/A NOR2X1_LOC_360/A 0.06fF
C5727 INVX1_LOC_186/Y INVX1_LOC_283/A 0.05fF
C5728 NOR2X1_LOC_16/Y NAND2X1_LOC_200/B 0.02fF
C5729 NAND2X1_LOC_477/Y INVX1_LOC_15/A 0.07fF
C5730 NAND2X1_LOC_464/B INVX1_LOC_118/A 0.10fF
C5731 NOR2X1_LOC_348/B INVX1_LOC_22/A 0.10fF
C5732 NOR2X1_LOC_500/A NOR2X1_LOC_542/Y -0.09fF
C5733 NOR2X1_LOC_445/a_36_216# INVX1_LOC_69/Y 0.01fF
C5734 INVX1_LOC_286/Y NOR2X1_LOC_74/A -0.02fF
C5735 VDD INVX1_LOC_306/Y 2.22fF
C5736 INVX1_LOC_178/A INVX1_LOC_20/A 0.07fF
C5737 INVX1_LOC_17/A NOR2X1_LOC_318/B 0.20fF
C5738 NAND2X1_LOC_360/a_36_24# INVX1_LOC_117/A 0.00fF
C5739 NOR2X1_LOC_439/B INVX1_LOC_18/A 0.03fF
C5740 NAND2X1_LOC_338/B INVX1_LOC_43/A 0.06fF
C5741 NAND2X1_LOC_361/Y INVX1_LOC_83/A 0.07fF
C5742 INVX1_LOC_223/A INVX1_LOC_67/Y 0.07fF
C5743 INVX1_LOC_25/Y INVX1_LOC_34/Y 0.02fF
C5744 NAND2X1_LOC_714/B INVX1_LOC_76/A 0.19fF
C5745 NAND2X1_LOC_722/A INVX1_LOC_16/A 0.10fF
C5746 NOR2X1_LOC_632/Y NAND2X1_LOC_147/a_36_24# 0.00fF
C5747 D_INPUT_0 NOR2X1_LOC_557/Y 0.14fF
C5748 INVX1_LOC_161/Y NOR2X1_LOC_78/A 0.07fF
C5749 INVX1_LOC_75/A INVX1_LOC_18/A 0.25fF
C5750 INVX1_LOC_17/A INVX1_LOC_93/Y 0.03fF
C5751 NAND2X1_LOC_206/B NAND2X1_LOC_202/a_36_24# 0.02fF
C5752 INVX1_LOC_50/A INVX1_LOC_92/A 0.53fF
C5753 INVX1_LOC_94/Y INVX1_LOC_63/A 0.03fF
C5754 NOR2X1_LOC_451/A NOR2X1_LOC_452/A 0.06fF
C5755 NOR2X1_LOC_778/B NOR2X1_LOC_553/Y 0.03fF
C5756 INVX1_LOC_182/A INVX1_LOC_71/A 0.07fF
C5757 NOR2X1_LOC_160/B NOR2X1_LOC_269/Y 0.07fF
C5758 D_INPUT_3 NOR2X1_LOC_611/a_36_216# 0.00fF
C5759 NOR2X1_LOC_595/a_36_216# INVX1_LOC_91/A 0.01fF
C5760 NAND2X1_LOC_560/A NAND2X1_LOC_837/Y 0.01fF
C5761 D_INPUT_3 NAND2X1_LOC_218/A 0.07fF
C5762 NOR2X1_LOC_392/Y NOR2X1_LOC_860/Y 0.20fF
C5763 NOR2X1_LOC_175/B INVX1_LOC_22/A 0.68fF
C5764 NAND2X1_LOC_493/Y INVX1_LOC_46/A 0.01fF
C5765 NOR2X1_LOC_140/A D_INPUT_3 0.00fF
C5766 NOR2X1_LOC_67/A INVX1_LOC_13/A 0.08fF
C5767 NOR2X1_LOC_91/Y INPUT_0 0.31fF
C5768 INVX1_LOC_256/A INVX1_LOC_95/Y 0.40fF
C5769 INVX1_LOC_104/A NAND2X1_LOC_140/A 0.01fF
C5770 NOR2X1_LOC_810/A INVX1_LOC_196/A 0.39fF
C5771 INVX1_LOC_75/A NOR2X1_LOC_713/B 0.03fF
C5772 NOR2X1_LOC_589/A NOR2X1_LOC_773/Y 0.09fF
C5773 NOR2X1_LOC_191/B NOR2X1_LOC_74/A 0.16fF
C5774 NOR2X1_LOC_197/A NOR2X1_LOC_631/B 0.01fF
C5775 NAND2X1_LOC_719/a_36_24# INVX1_LOC_76/A 0.01fF
C5776 NOR2X1_LOC_280/a_36_216# INVX1_LOC_285/A 0.00fF
C5777 NOR2X1_LOC_522/Y INVX1_LOC_309/A 0.01fF
C5778 INVX1_LOC_59/A NOR2X1_LOC_536/A 0.03fF
C5779 NOR2X1_LOC_716/B NOR2X1_LOC_322/Y 0.10fF
C5780 INVX1_LOC_1/A INVX1_LOC_117/A 0.36fF
C5781 NOR2X1_LOC_816/A INVX1_LOC_20/A 0.09fF
C5782 D_INPUT_0 INVX1_LOC_143/A 0.11fF
C5783 NAND2X1_LOC_656/A INVX1_LOC_6/A 0.02fF
C5784 NOR2X1_LOC_191/B NOR2X1_LOC_9/Y 0.19fF
C5785 NOR2X1_LOC_498/Y NAND2X1_LOC_560/A 0.00fF
C5786 INVX1_LOC_17/A NAND2X1_LOC_721/A 0.03fF
C5787 NOR2X1_LOC_78/B NAND2X1_LOC_660/a_36_24# 0.01fF
C5788 NOR2X1_LOC_621/a_36_216# INVX1_LOC_63/A 0.01fF
C5789 INVX1_LOC_81/Y NAND2X1_LOC_468/B 0.01fF
C5790 NAND2X1_LOC_773/Y NOR2X1_LOC_536/A 0.05fF
C5791 NOR2X1_LOC_598/B NAND2X1_LOC_574/A 0.02fF
C5792 INVX1_LOC_50/Y NOR2X1_LOC_640/Y 0.09fF
C5793 INVX1_LOC_311/A INVX1_LOC_113/Y 0.02fF
C5794 NOR2X1_LOC_522/Y INVX1_LOC_91/A 0.05fF
C5795 NAND2X1_LOC_833/Y NOR2X1_LOC_527/Y 0.09fF
C5796 NAND2X1_LOC_722/A INVX1_LOC_28/A 0.02fF
C5797 INVX1_LOC_21/A INVX1_LOC_291/A 0.03fF
C5798 NOR2X1_LOC_716/B INVX1_LOC_92/Y 0.01fF
C5799 NAND2X1_LOC_565/B D_INPUT_0 0.03fF
C5800 NAND2X1_LOC_348/A NAND2X1_LOC_116/A 0.07fF
C5801 INVX1_LOC_30/A NOR2X1_LOC_35/Y 0.03fF
C5802 INVX1_LOC_278/A NAND2X1_LOC_477/Y 0.02fF
C5803 INVX1_LOC_78/A INVX1_LOC_19/Y 0.08fF
C5804 NAND2X1_LOC_338/B NOR2X1_LOC_756/Y 0.01fF
C5805 INVX1_LOC_185/Y NOR2X1_LOC_74/A 0.02fF
C5806 INVX1_LOC_93/A NOR2X1_LOC_88/Y 0.07fF
C5807 INVX1_LOC_57/A NAND2X1_LOC_81/B 0.99fF
C5808 INVX1_LOC_50/Y NAND2X1_LOC_85/Y 0.08fF
C5809 NOR2X1_LOC_186/Y NAND2X1_LOC_288/A 0.98fF
C5810 NOR2X1_LOC_296/Y NAND2X1_LOC_297/a_36_24# 0.00fF
C5811 INVX1_LOC_132/A INVX1_LOC_125/Y 0.02fF
C5812 NAND2X1_LOC_660/Y NOR2X1_LOC_130/A 0.03fF
C5813 INVX1_LOC_90/A INVX1_LOC_232/A 0.03fF
C5814 INVX1_LOC_75/A INVX1_LOC_34/Y 0.07fF
C5815 INVX1_LOC_201/Y INVX1_LOC_201/A 0.26fF
C5816 NOR2X1_LOC_657/Y VDD 0.35fF
C5817 INVX1_LOC_266/A NOR2X1_LOC_640/Y 0.03fF
C5818 INVX1_LOC_308/Y INVX1_LOC_118/A 0.12fF
C5819 NAND2X1_LOC_773/Y NAND2X1_LOC_93/B 0.03fF
C5820 INVX1_LOC_58/A INVX1_LOC_261/Y 0.03fF
C5821 NOR2X1_LOC_389/B INVX1_LOC_232/A 0.15fF
C5822 NAND2X1_LOC_350/A NOR2X1_LOC_331/B 0.17fF
C5823 INVX1_LOC_269/A NOR2X1_LOC_660/a_36_216# 0.01fF
C5824 INVX1_LOC_32/A NAND2X1_LOC_61/Y 0.01fF
C5825 INVX1_LOC_18/A NAND2X1_LOC_453/A 0.12fF
C5826 NOR2X1_LOC_92/Y NOR2X1_LOC_58/Y 0.02fF
C5827 NAND2X1_LOC_573/Y NAND2X1_LOC_288/A 0.65fF
C5828 NOR2X1_LOC_186/Y NOR2X1_LOC_653/Y 0.08fF
C5829 NOR2X1_LOC_383/Y INVX1_LOC_90/A 0.02fF
C5830 INVX1_LOC_15/Y NAND2X1_LOC_622/B 0.01fF
C5831 NOR2X1_LOC_418/Y INVX1_LOC_140/A 0.15fF
C5832 NOR2X1_LOC_423/Y INVX1_LOC_6/A 0.09fF
C5833 INVX1_LOC_9/Y NOR2X1_LOC_135/Y 0.18fF
C5834 NOR2X1_LOC_273/Y INVX1_LOC_76/A 0.07fF
C5835 D_INPUT_0 NOR2X1_LOC_130/A 0.99fF
C5836 NOR2X1_LOC_495/Y NOR2X1_LOC_164/Y 0.11fF
C5837 NOR2X1_LOC_516/B NOR2X1_LOC_567/B 0.10fF
C5838 NOR2X1_LOC_244/B NAND2X1_LOC_348/A 0.01fF
C5839 NOR2X1_LOC_759/Y INVX1_LOC_76/A 0.01fF
C5840 NOR2X1_LOC_441/Y NOR2X1_LOC_331/B 0.07fF
C5841 INVX1_LOC_252/Y NOR2X1_LOC_655/Y 0.01fF
C5842 NOR2X1_LOC_68/A NOR2X1_LOC_111/A 0.10fF
C5843 NOR2X1_LOC_32/B INVX1_LOC_284/A 1.02fF
C5844 INVX1_LOC_88/A NOR2X1_LOC_831/B 0.24fF
C5845 INVX1_LOC_230/Y NOR2X1_LOC_629/Y 0.00fF
C5846 NAND2X1_LOC_348/A INVX1_LOC_232/A 0.00fF
C5847 NOR2X1_LOC_637/Y NAND2X1_LOC_453/A 0.02fF
C5848 NOR2X1_LOC_186/Y INVX1_LOC_19/A 0.11fF
C5849 INVX1_LOC_24/A NOR2X1_LOC_682/Y 0.08fF
C5850 INVX1_LOC_25/A INVX1_LOC_3/Y 3.72fF
C5851 NOR2X1_LOC_222/Y INVX1_LOC_6/A 0.07fF
C5852 NAND2X1_LOC_194/a_36_24# NOR2X1_LOC_188/A 0.00fF
C5853 NOR2X1_LOC_380/A NAND2X1_LOC_866/B 0.02fF
C5854 NOR2X1_LOC_550/B INVX1_LOC_76/A 0.03fF
C5855 INVX1_LOC_14/A NOR2X1_LOC_179/Y 0.00fF
C5856 NOR2X1_LOC_495/Y INVX1_LOC_46/A 0.05fF
C5857 INVX1_LOC_83/A NAND2X1_LOC_654/B 0.03fF
C5858 NAND2X1_LOC_593/Y NOR2X1_LOC_447/B 0.01fF
C5859 NAND2X1_LOC_350/A NOR2X1_LOC_592/B 0.03fF
C5860 NOR2X1_LOC_526/Y NOR2X1_LOC_526/a_36_216# 0.00fF
C5861 INVX1_LOC_136/A INVX1_LOC_9/A 0.11fF
C5862 INVX1_LOC_57/A INVX1_LOC_4/Y 1.28fF
C5863 INVX1_LOC_71/A NOR2X1_LOC_176/Y 0.01fF
C5864 NOR2X1_LOC_299/Y NAND2X1_LOC_560/A 6.13fF
C5865 NAND2X1_LOC_573/Y INVX1_LOC_19/A 0.16fF
C5866 INVX1_LOC_299/A INVX1_LOC_63/A 0.07fF
C5867 INVX1_LOC_89/A INVX1_LOC_148/A 0.00fF
C5868 NOR2X1_LOC_557/Y NOR2X1_LOC_266/B 0.00fF
C5869 NAND2X1_LOC_741/B NOR2X1_LOC_51/A 0.06fF
C5870 INVX1_LOC_24/A NAND2X1_LOC_848/A 0.04fF
C5871 NOR2X1_LOC_329/B INVX1_LOC_313/A 0.00fF
C5872 NAND2X1_LOC_320/a_36_24# NOR2X1_LOC_324/A 0.00fF
C5873 NOR2X1_LOC_802/A NOR2X1_LOC_799/B 0.25fF
C5874 INVX1_LOC_49/A NAND2X1_LOC_472/Y 0.07fF
C5875 NOR2X1_LOC_538/B INVX1_LOC_63/A 0.01fF
C5876 NOR2X1_LOC_19/B NOR2X1_LOC_5/a_36_216# 0.00fF
C5877 INVX1_LOC_294/Y VDD 0.19fF
C5878 NOR2X1_LOC_92/Y INVX1_LOC_29/A 0.10fF
C5879 INVX1_LOC_252/Y INVX1_LOC_3/A 0.01fF
C5880 INVX1_LOC_256/Y NOR2X1_LOC_124/A 0.11fF
C5881 INPUT_2 NOR2X1_LOC_814/A 0.05fF
C5882 INVX1_LOC_24/Y INVX1_LOC_29/A 1.34fF
C5883 INVX1_LOC_5/A INVX1_LOC_4/A 0.31fF
C5884 INVX1_LOC_93/A INVX1_LOC_15/A 0.07fF
C5885 NAND2X1_LOC_860/Y INVX1_LOC_304/A 0.03fF
C5886 INVX1_LOC_14/Y NOR2X1_LOC_709/A 0.07fF
C5887 INVX1_LOC_209/Y INVX1_LOC_118/A 0.09fF
C5888 INVX1_LOC_49/A NAND2X1_LOC_637/Y 0.05fF
C5889 NOR2X1_LOC_773/Y INVX1_LOC_20/A 0.08fF
C5890 NOR2X1_LOC_134/Y NAND2X1_LOC_773/B 0.01fF
C5891 INVX1_LOC_21/A NOR2X1_LOC_609/Y 0.01fF
C5892 NOR2X1_LOC_142/Y NOR2X1_LOC_331/B 0.10fF
C5893 INVX1_LOC_33/A NOR2X1_LOC_149/a_36_216# 0.02fF
C5894 INVX1_LOC_24/A INVX1_LOC_46/Y 0.14fF
C5895 NOR2X1_LOC_647/A NOR2X1_LOC_392/Y 0.03fF
C5896 NAND2X1_LOC_513/B INVX1_LOC_15/A 0.04fF
C5897 NAND2X1_LOC_859/B NOR2X1_LOC_670/Y 0.25fF
C5898 INVX1_LOC_223/A NOR2X1_LOC_814/A 0.00fF
C5899 NOR2X1_LOC_91/A INVX1_LOC_35/A 0.03fF
C5900 INVX1_LOC_2/A NAND2X1_LOC_472/Y 0.07fF
C5901 INVX1_LOC_35/A NOR2X1_LOC_201/A 0.04fF
C5902 INVX1_LOC_50/A INVX1_LOC_53/A 0.27fF
C5903 INVX1_LOC_1/A INVX1_LOC_3/Y 0.10fF
C5904 NOR2X1_LOC_137/A INVX1_LOC_91/A 0.07fF
C5905 NOR2X1_LOC_45/B NOR2X1_LOC_71/Y 0.07fF
C5906 NOR2X1_LOC_249/Y NAND2X1_LOC_223/A 0.02fF
C5907 INVX1_LOC_141/Y INVX1_LOC_49/Y 0.01fF
C5908 NOR2X1_LOC_272/Y NAND2X1_LOC_454/Y 0.01fF
C5909 NOR2X1_LOC_626/Y INVX1_LOC_78/A 0.06fF
C5910 NOR2X1_LOC_329/B INVX1_LOC_6/A 0.03fF
C5911 NOR2X1_LOC_337/Y NOR2X1_LOC_356/A 0.01fF
C5912 NAND2X1_LOC_740/Y NOR2X1_LOC_829/A 0.37fF
C5913 NOR2X1_LOC_773/Y NOR2X1_LOC_765/Y 0.00fF
C5914 INVX1_LOC_75/A NOR2X1_LOC_548/A 0.15fF
C5915 INVX1_LOC_77/A NOR2X1_LOC_117/a_36_216# 0.01fF
C5916 NOR2X1_LOC_342/A NOR2X1_LOC_260/Y 0.01fF
C5917 NOR2X1_LOC_19/B INVX1_LOC_123/A 0.05fF
C5918 NAND2X1_LOC_149/B VDD 0.01fF
C5919 NOR2X1_LOC_456/Y NOR2X1_LOC_455/Y 0.02fF
C5920 INVX1_LOC_35/A INVX1_LOC_23/A 0.78fF
C5921 INVX1_LOC_41/A NOR2X1_LOC_634/A 0.02fF
C5922 NOR2X1_LOC_210/A INVX1_LOC_37/A 0.04fF
C5923 NAND2X1_LOC_861/Y INVX1_LOC_304/A 0.47fF
C5924 INVX1_LOC_30/A INVX1_LOC_109/A 0.12fF
C5925 NOR2X1_LOC_332/A INVX1_LOC_20/A 0.08fF
C5926 NOR2X1_LOC_721/Y NOR2X1_LOC_9/Y 0.00fF
C5927 NOR2X1_LOC_613/Y NOR2X1_LOC_693/Y 0.04fF
C5928 NAND2X1_LOC_135/a_36_24# NOR2X1_LOC_243/B 0.01fF
C5929 NAND2X1_LOC_72/Y INVX1_LOC_53/A 0.01fF
C5930 NOR2X1_LOC_180/Y INVX1_LOC_179/A 0.02fF
C5931 D_INPUT_0 NOR2X1_LOC_280/Y 0.03fF
C5932 NAND2X1_LOC_214/B D_INPUT_1 0.03fF
C5933 INVX1_LOC_119/A NAND2X1_LOC_798/B 0.28fF
C5934 INVX1_LOC_90/A NAND2X1_LOC_447/Y 0.01fF
C5935 NOR2X1_LOC_791/B INVX1_LOC_12/A 0.03fF
C5936 NOR2X1_LOC_644/A INVX1_LOC_247/A 0.00fF
C5937 NOR2X1_LOC_337/Y NOR2X1_LOC_74/A 0.02fF
C5938 NAND2X1_LOC_463/B INVX1_LOC_167/Y 0.01fF
C5939 NOR2X1_LOC_389/B NAND2X1_LOC_447/Y 0.01fF
C5940 INVX1_LOC_17/A INVX1_LOC_87/A 0.02fF
C5941 NOR2X1_LOC_6/B NAND2X1_LOC_85/Y 0.16fF
C5942 INVX1_LOC_214/A INVX1_LOC_291/A 0.05fF
C5943 NOR2X1_LOC_802/A NOR2X1_LOC_445/B 0.04fF
C5944 INVX1_LOC_10/A NOR2X1_LOC_363/Y 0.08fF
C5945 NOR2X1_LOC_226/A NAND2X1_LOC_434/Y 0.01fF
C5946 INVX1_LOC_256/A INVX1_LOC_271/Y 0.09fF
C5947 NOR2X1_LOC_808/A NOR2X1_LOC_809/B 0.01fF
C5948 INVX1_LOC_162/Y INVX1_LOC_285/A 0.15fF
C5949 NAND2X1_LOC_35/Y NAND2X1_LOC_725/A 0.10fF
C5950 NAND2X1_LOC_474/Y INVX1_LOC_29/Y 0.04fF
C5951 D_INPUT_1 INVX1_LOC_27/A 2.38fF
C5952 NOR2X1_LOC_84/A INVX1_LOC_84/A 0.16fF
C5953 INVX1_LOC_132/A INVX1_LOC_19/A 0.07fF
C5954 INVX1_LOC_64/A INVX1_LOC_5/A 0.54fF
C5955 INVX1_LOC_124/A NOR2X1_LOC_117/a_36_216# 0.00fF
C5956 NOR2X1_LOC_374/A INVX1_LOC_19/A 0.03fF
C5957 INVX1_LOC_225/A NOR2X1_LOC_653/Y 0.01fF
C5958 INVX1_LOC_278/A INVX1_LOC_93/A 0.09fF
C5959 NOR2X1_LOC_238/Y NOR2X1_LOC_89/A 0.14fF
C5960 NAND2X1_LOC_783/A NAND2X1_LOC_848/A 0.03fF
C5961 NAND2X1_LOC_479/Y INVX1_LOC_54/A 0.03fF
C5962 NOR2X1_LOC_384/Y INVX1_LOC_3/Y 0.01fF
C5963 NOR2X1_LOC_121/a_36_216# NOR2X1_LOC_99/Y 0.01fF
C5964 NOR2X1_LOC_356/A VDD 0.12fF
C5965 NAND2X1_LOC_175/a_36_24# INVX1_LOC_271/A 0.01fF
C5966 INVX1_LOC_223/Y NAND2X1_LOC_533/a_36_24# 0.00fF
C5967 INVX1_LOC_140/A INVX1_LOC_20/A 0.03fF
C5968 NAND2X1_LOC_350/A NOR2X1_LOC_449/A 0.08fF
C5969 INVX1_LOC_48/A INVX1_LOC_91/A 0.35fF
C5970 INVX1_LOC_58/A INVX1_LOC_1/A 0.21fF
C5971 INVX1_LOC_24/A NOR2X1_LOC_754/A 0.47fF
C5972 NOR2X1_LOC_315/Y INVX1_LOC_63/A 0.07fF
C5973 INVX1_LOC_64/A INVX1_LOC_178/A 0.07fF
C5974 NOR2X1_LOC_160/B INVX1_LOC_26/A 0.13fF
C5975 NOR2X1_LOC_716/B INVX1_LOC_106/A 0.01fF
C5976 NOR2X1_LOC_496/Y NAND2X1_LOC_624/B 0.06fF
C5977 INVX1_LOC_54/Y INVX1_LOC_84/A 0.46fF
C5978 NAND2X1_LOC_555/Y INVX1_LOC_175/A 0.20fF
C5979 INVX1_LOC_225/A INVX1_LOC_19/A 0.12fF
C5980 INVX1_LOC_41/A INVX1_LOC_29/A 0.08fF
C5981 NOR2X1_LOC_288/A INVX1_LOC_19/A 1.02fF
C5982 NAND2X1_LOC_581/a_36_24# INVX1_LOC_1/A 0.01fF
C5983 NAND2X1_LOC_579/A NAND2X1_LOC_793/B 0.10fF
C5984 INVX1_LOC_201/Y INVX1_LOC_29/A 0.17fF
C5985 NOR2X1_LOC_15/Y NOR2X1_LOC_717/A 0.08fF
C5986 INVX1_LOC_279/A NAND2X1_LOC_93/B 0.07fF
C5987 INVX1_LOC_135/A INVX1_LOC_54/A 0.10fF
C5988 NOR2X1_LOC_500/A INVX1_LOC_15/A 0.09fF
C5989 NAND2X1_LOC_739/B INVX1_LOC_231/A 0.32fF
C5990 NAND2X1_LOC_548/a_36_24# INVX1_LOC_84/A 0.00fF
C5991 INVX1_LOC_286/A NOR2X1_LOC_566/a_36_216# 0.01fF
C5992 INVX1_LOC_27/A NOR2X1_LOC_652/Y 0.12fF
C5993 INVX1_LOC_64/A NOR2X1_LOC_494/Y 0.05fF
C5994 NOR2X1_LOC_67/A NAND2X1_LOC_489/Y 0.02fF
C5995 NOR2X1_LOC_303/Y INVX1_LOC_15/A 0.07fF
C5996 INVX1_LOC_266/Y NOR2X1_LOC_48/Y 0.72fF
C5997 INVX1_LOC_219/Y NOR2X1_LOC_671/Y 0.01fF
C5998 VDD NOR2X1_LOC_74/A 2.19fF
C5999 NAND2X1_LOC_477/A INVX1_LOC_29/A 0.03fF
C6000 NOR2X1_LOC_209/Y INVX1_LOC_19/A 0.46fF
C6001 NOR2X1_LOC_97/A INVX1_LOC_37/A 0.08fF
C6002 NOR2X1_LOC_389/A INVX1_LOC_270/Y 1.16fF
C6003 NAND2X1_LOC_703/Y NOR2X1_LOC_406/A 0.02fF
C6004 INVX1_LOC_36/A NAND2X1_LOC_99/A 0.48fF
C6005 NOR2X1_LOC_312/Y NOR2X1_LOC_743/Y 0.01fF
C6006 NOR2X1_LOC_322/Y NOR2X1_LOC_322/a_36_216# 0.01fF
C6007 VDD NOR2X1_LOC_9/Y 1.14fF
C6008 INVX1_LOC_77/A NAND2X1_LOC_647/B 0.18fF
C6009 NOR2X1_LOC_828/B NOR2X1_LOC_499/B 0.96fF
C6010 NAND2X1_LOC_198/B NOR2X1_LOC_278/Y 0.40fF
C6011 NOR2X1_LOC_188/A INVX1_LOC_117/A 0.89fF
C6012 NOR2X1_LOC_361/B INVX1_LOC_306/Y 0.19fF
C6013 NOR2X1_LOC_128/B NAND2X1_LOC_141/Y 0.01fF
C6014 NAND2X1_LOC_740/Y NAND2X1_LOC_537/Y 0.16fF
C6015 NOR2X1_LOC_91/Y INVX1_LOC_183/A 0.02fF
C6016 NOR2X1_LOC_254/Y INVX1_LOC_15/A 0.07fF
C6017 INVX1_LOC_64/A NOR2X1_LOC_816/A 0.03fF
C6018 NOR2X1_LOC_548/B INVX1_LOC_117/A 0.07fF
C6019 INVX1_LOC_22/A INVX1_LOC_186/Y 0.07fF
C6020 NOR2X1_LOC_703/B NOR2X1_LOC_383/B 0.01fF
C6021 NOR2X1_LOC_532/Y NOR2X1_LOC_445/B 0.01fF
C6022 NOR2X1_LOC_269/Y NAND2X1_LOC_211/Y 0.07fF
C6023 NOR2X1_LOC_540/B INVX1_LOC_247/A 0.03fF
C6024 NOR2X1_LOC_644/A NOR2X1_LOC_862/B 0.03fF
C6025 INVX1_LOC_35/A INVX1_LOC_31/A 12.01fF
C6026 NOR2X1_LOC_753/Y NAND2X1_LOC_175/Y 0.07fF
C6027 INVX1_LOC_58/A NOR2X1_LOC_384/Y 0.06fF
C6028 INVX1_LOC_153/A INVX1_LOC_78/A 0.01fF
C6029 INVX1_LOC_7/A INVX1_LOC_293/Y 0.07fF
C6030 NAND2X1_LOC_35/Y NOR2X1_LOC_372/A 0.03fF
C6031 INVX1_LOC_182/Y NAND2X1_LOC_93/B 0.03fF
C6032 NAND2X1_LOC_325/Y NAND2X1_LOC_175/Y 0.07fF
C6033 NOR2X1_LOC_237/Y NAND2X1_LOC_99/A 0.01fF
C6034 INVX1_LOC_124/A NAND2X1_LOC_647/B 0.00fF
C6035 INVX1_LOC_132/A INVX1_LOC_26/Y 0.07fF
C6036 NAND2X1_LOC_392/a_36_24# NAND2X1_LOC_793/Y 0.00fF
C6037 INVX1_LOC_56/Y NOR2X1_LOC_76/B 0.01fF
C6038 INPUT_1 NOR2X1_LOC_813/a_36_216# 0.00fF
C6039 NOR2X1_LOC_639/B INVX1_LOC_72/A 0.63fF
C6040 INVX1_LOC_33/A INVX1_LOC_23/Y 0.07fF
C6041 NOR2X1_LOC_67/A INVX1_LOC_32/A 0.47fF
C6042 NOR2X1_LOC_43/Y INVX1_LOC_117/A 0.00fF
C6043 NOR2X1_LOC_561/Y NAND2X1_LOC_74/B 0.03fF
C6044 NOR2X1_LOC_731/a_36_216# INVX1_LOC_213/A 0.01fF
C6045 NAND2X1_LOC_656/Y INVX1_LOC_49/Y 0.03fF
C6046 NOR2X1_LOC_93/Y INVX1_LOC_230/Y 0.06fF
C6047 INVX1_LOC_7/A NAND2X1_LOC_74/B 0.07fF
C6048 INVX1_LOC_5/A NOR2X1_LOC_585/a_36_216# 0.02fF
C6049 INVX1_LOC_7/A NAND2X1_LOC_207/Y 0.01fF
C6050 NOR2X1_LOC_784/B NOR2X1_LOC_777/B 0.02fF
C6051 INVX1_LOC_1/A NOR2X1_LOC_738/Y 0.01fF
C6052 NOR2X1_LOC_594/Y INVX1_LOC_117/Y 0.02fF
C6053 NOR2X1_LOC_186/Y INVX1_LOC_312/A -0.03fF
C6054 NOR2X1_LOC_718/B NOR2X1_LOC_631/Y 0.06fF
C6055 NOR2X1_LOC_68/A INVX1_LOC_138/Y 0.69fF
C6056 INVX1_LOC_259/A INVX1_LOC_78/A 0.06fF
C6057 NOR2X1_LOC_773/Y INVX1_LOC_4/A 0.00fF
C6058 INVX1_LOC_73/A NAND2X1_LOC_572/B 0.02fF
C6059 INPUT_1 NAND2X1_LOC_773/B 0.10fF
C6060 NAND2X1_LOC_833/Y NOR2X1_LOC_654/A 0.06fF
C6061 INVX1_LOC_35/A INVX1_LOC_111/A 0.05fF
C6062 NAND2X1_LOC_794/B INVX1_LOC_30/A 0.01fF
C6063 NOR2X1_LOC_510/Y NOR2X1_LOC_657/Y 0.01fF
C6064 NAND2X1_LOC_99/Y D_INPUT_1 0.01fF
C6065 INVX1_LOC_64/A NOR2X1_LOC_759/a_36_216# 0.01fF
C6066 INVX1_LOC_105/A INVX1_LOC_53/A 0.07fF
C6067 NOR2X1_LOC_730/B NOR2X1_LOC_155/A 0.01fF
C6068 NOR2X1_LOC_189/A NAND2X1_LOC_787/A 0.00fF
C6069 INVX1_LOC_276/A NAND2X1_LOC_175/Y 0.98fF
C6070 NOR2X1_LOC_764/a_36_216# D_INPUT_5 0.00fF
C6071 INVX1_LOC_230/Y INVX1_LOC_269/A 0.10fF
C6072 NAND2X1_LOC_573/Y INVX1_LOC_312/A -0.01fF
C6073 NAND2X1_LOC_559/Y INVX1_LOC_284/Y 0.03fF
C6074 INVX1_LOC_235/Y NOR2X1_LOC_476/Y 0.04fF
C6075 NOR2X1_LOC_246/A NAND2X1_LOC_807/a_36_24# 0.01fF
C6076 INVX1_LOC_171/A INVX1_LOC_42/A 0.03fF
C6077 NOR2X1_LOC_418/Y INVX1_LOC_78/A 0.01fF
C6078 NAND2X1_LOC_848/A NOR2X1_LOC_280/Y 0.05fF
C6079 NOR2X1_LOC_647/B INVX1_LOC_252/Y 0.20fF
C6080 INVX1_LOC_36/A NOR2X1_LOC_464/B 0.01fF
C6081 INVX1_LOC_201/A NAND2X1_LOC_574/A 0.01fF
C6082 NAND2X1_LOC_555/Y NOR2X1_LOC_82/A 0.03fF
C6083 INVX1_LOC_116/A NOR2X1_LOC_798/A 0.01fF
C6084 NAND2X1_LOC_858/B NOR2X1_LOC_661/A 0.03fF
C6085 INVX1_LOC_40/A INVX1_LOC_23/Y 0.02fF
C6086 INVX1_LOC_17/A NAND2X1_LOC_36/A 0.71fF
C6087 INVX1_LOC_53/Y NOR2X1_LOC_278/Y 0.03fF
C6088 INVX1_LOC_165/Y INVX1_LOC_23/Y 0.01fF
C6089 NAND2X1_LOC_213/A NOR2X1_LOC_68/A 0.04fF
C6090 NOR2X1_LOC_589/A INVX1_LOC_78/A 0.91fF
C6091 NOR2X1_LOC_15/Y NOR2X1_LOC_518/Y 0.01fF
C6092 INVX1_LOC_27/A D_INPUT_2 0.08fF
C6093 NOR2X1_LOC_332/A INVX1_LOC_4/A 0.09fF
C6094 NOR2X1_LOC_181/Y NOR2X1_LOC_678/A 0.01fF
C6095 INVX1_LOC_50/A NOR2X1_LOC_78/B 5.51fF
C6096 NOR2X1_LOC_586/Y NAND2X1_LOC_637/Y 0.07fF
C6097 INVX1_LOC_89/A INVX1_LOC_47/Y 0.08fF
C6098 INPUT_0 NAND2X1_LOC_82/Y 0.66fF
C6099 INVX1_LOC_64/A NAND2X1_LOC_562/B 0.03fF
C6100 NOR2X1_LOC_655/B NOR2X1_LOC_493/A 0.31fF
C6101 NOR2X1_LOC_626/Y INVX1_LOC_113/Y 0.01fF
C6102 NAND2X1_LOC_787/A NOR2X1_LOC_482/Y 0.02fF
C6103 INVX1_LOC_22/A NOR2X1_LOC_843/B 0.17fF
C6104 NAND2X1_LOC_862/A INVX1_LOC_57/A 0.01fF
C6105 NOR2X1_LOC_218/A INVX1_LOC_72/A 0.00fF
C6106 NOR2X1_LOC_603/Y INVX1_LOC_179/A 0.01fF
C6107 INVX1_LOC_305/Y INVX1_LOC_23/A 0.00fF
C6108 NAND2X1_LOC_287/B NOR2X1_LOC_743/Y 0.00fF
C6109 INVX1_LOC_47/A INVX1_LOC_104/Y 0.01fF
C6110 NOR2X1_LOC_112/Y INVX1_LOC_15/A 0.12fF
C6111 NOR2X1_LOC_65/B NOR2X1_LOC_589/A 0.07fF
C6112 NOR2X1_LOC_331/B NAND2X1_LOC_61/a_36_24# 0.01fF
C6113 NOR2X1_LOC_590/A INVX1_LOC_223/A 0.07fF
C6114 NAND2X1_LOC_642/Y NOR2X1_LOC_653/Y 0.01fF
C6115 NOR2X1_LOC_319/B NOR2X1_LOC_729/A 0.05fF
C6116 D_INPUT_3 NOR2X1_LOC_104/a_36_216# 0.00fF
C6117 INVX1_LOC_137/A NAND2X1_LOC_90/a_36_24# 0.00fF
C6118 NAND2X1_LOC_30/Y INVX1_LOC_24/A 0.04fF
C6119 NAND2X1_LOC_36/a_36_24# INVX1_LOC_174/A 0.00fF
C6120 NAND2X1_LOC_363/B NAND2X1_LOC_292/a_36_24# 0.01fF
C6121 D_INPUT_1 INVX1_LOC_137/A 0.01fF
C6122 INVX1_LOC_314/A NOR2X1_LOC_814/A 0.03fF
C6123 INVX1_LOC_64/A NOR2X1_LOC_773/Y 0.07fF
C6124 NOR2X1_LOC_644/A NOR2X1_LOC_465/Y 0.18fF
C6125 INVX1_LOC_5/A INVX1_LOC_44/Y 0.01fF
C6126 NOR2X1_LOC_791/Y NOR2X1_LOC_84/Y 0.04fF
C6127 VDD NOR2X1_LOC_865/Y 0.66fF
C6128 NOR2X1_LOC_363/Y INVX1_LOC_307/A 0.12fF
C6129 NOR2X1_LOC_188/Y INVX1_LOC_23/A 0.01fF
C6130 NOR2X1_LOC_92/Y INVX1_LOC_8/A 0.26fF
C6131 NAND2X1_LOC_794/B NAND2X1_LOC_722/A 0.02fF
C6132 NAND2X1_LOC_642/Y INVX1_LOC_19/A 0.07fF
C6133 NAND2X1_LOC_93/B NOR2X1_LOC_98/B 0.03fF
C6134 NAND2X1_LOC_276/Y INVX1_LOC_14/A 0.04fF
C6135 NOR2X1_LOC_134/Y INVX1_LOC_24/A 1.38fF
C6136 NAND2X1_LOC_799/A NOR2X1_LOC_577/Y 0.07fF
C6137 NOR2X1_LOC_65/B INVX1_LOC_171/A 0.03fF
C6138 D_INPUT_1 INVX1_LOC_234/A 0.17fF
C6139 NOR2X1_LOC_609/a_36_216# INVX1_LOC_292/A 0.00fF
C6140 INVX1_LOC_83/A NOR2X1_LOC_105/Y 0.01fF
C6141 INVX1_LOC_135/A NAND2X1_LOC_215/A -0.02fF
C6142 INVX1_LOC_293/Y INVX1_LOC_76/A -0.02fF
C6143 NAND2X1_LOC_93/B NOR2X1_LOC_450/A 0.02fF
C6144 INVX1_LOC_167/Y INVX1_LOC_42/A 0.75fF
C6145 NOR2X1_LOC_481/A INVX1_LOC_161/Y 0.09fF
C6146 INVX1_LOC_18/A NOR2X1_LOC_274/B 0.59fF
C6147 NOR2X1_LOC_160/B NOR2X1_LOC_712/B 0.06fF
C6148 NOR2X1_LOC_841/A NOR2X1_LOC_60/Y 0.04fF
C6149 NAND2X1_LOC_434/Y INVX1_LOC_118/A 0.04fF
C6150 INVX1_LOC_124/Y NOR2X1_LOC_191/B 0.04fF
C6151 INVX1_LOC_27/A NOR2X1_LOC_620/B 0.04fF
C6152 NOR2X1_LOC_151/Y NOR2X1_LOC_464/Y 0.29fF
C6153 INVX1_LOC_36/A NAND2X1_LOC_656/A 0.13fF
C6154 NOR2X1_LOC_445/a_36_216# NOR2X1_LOC_593/Y 0.03fF
C6155 NOR2X1_LOC_68/A NAND2X1_LOC_364/A 0.64fF
C6156 NAND2X1_LOC_425/Y NOR2X1_LOC_450/A 0.01fF
C6157 NOR2X1_LOC_596/Y INVX1_LOC_33/A 0.02fF
C6158 INVX1_LOC_95/Y NOR2X1_LOC_89/A 0.03fF
C6159 INVX1_LOC_222/A INVX1_LOC_78/A 0.07fF
C6160 INVX1_LOC_76/A NAND2X1_LOC_74/B 0.18fF
C6161 INVX1_LOC_64/A NOR2X1_LOC_332/A 0.56fF
C6162 INVX1_LOC_41/A NOR2X1_LOC_181/a_36_216# 0.00fF
C6163 INVX1_LOC_224/Y NOR2X1_LOC_756/Y 0.06fF
C6164 NAND2X1_LOC_96/A INVX1_LOC_63/A 0.07fF
C6165 NOR2X1_LOC_447/Y INVX1_LOC_72/A 0.02fF
C6166 D_GATE_579 INVX1_LOC_242/A 0.01fF
C6167 NOR2X1_LOC_590/A INVX1_LOC_149/Y 0.54fF
C6168 NAND2X1_LOC_573/A INVX1_LOC_306/Y 0.01fF
C6169 INVX1_LOC_208/A NOR2X1_LOC_666/A 0.01fF
C6170 NOR2X1_LOC_89/A NOR2X1_LOC_305/Y 0.07fF
C6171 NAND2X1_LOC_348/A INVX1_LOC_112/Y 0.01fF
C6172 D_INPUT_1 NOR2X1_LOC_19/B 1.96fF
C6173 NOR2X1_LOC_510/Y NOR2X1_LOC_171/a_36_216# 0.00fF
C6174 NOR2X1_LOC_34/A NAND2X1_LOC_24/a_36_24# 0.01fF
C6175 INVX1_LOC_20/A INVX1_LOC_42/A 0.32fF
C6176 NOR2X1_LOC_590/A INVX1_LOC_85/A 0.29fF
C6177 NAND2X1_LOC_588/B INVX1_LOC_77/A 0.03fF
C6178 NAND2X1_LOC_349/B NOR2X1_LOC_321/Y 0.01fF
C6179 NAND2X1_LOC_650/B INVX1_LOC_102/A 0.09fF
C6180 INVX1_LOC_18/A NOR2X1_LOC_577/Y 0.07fF
C6181 INVX1_LOC_56/Y NOR2X1_LOC_271/B 0.46fF
C6182 NAND2X1_LOC_652/Y INVX1_LOC_53/A 0.02fF
C6183 NAND2X1_LOC_728/Y NOR2X1_LOC_577/Y 0.08fF
C6184 NOR2X1_LOC_318/B INVX1_LOC_94/Y 0.05fF
C6185 NOR2X1_LOC_103/Y INVX1_LOC_43/A 0.10fF
C6186 INVX1_LOC_35/A NAND2X1_LOC_807/Y 0.98fF
C6187 INVX1_LOC_45/A INVX1_LOC_213/Y 0.01fF
C6188 NOR2X1_LOC_363/Y INVX1_LOC_12/A 0.07fF
C6189 INVX1_LOC_24/A INVX1_LOC_49/A 2.32fF
C6190 INVX1_LOC_279/A NOR2X1_LOC_348/Y 0.45fF
C6191 INVX1_LOC_118/A NAND2X1_LOC_773/B 0.01fF
C6192 NOR2X1_LOC_263/a_36_216# INVX1_LOC_36/A 0.00fF
C6193 INVX1_LOC_58/A NOR2X1_LOC_188/A 0.19fF
C6194 INVX1_LOC_64/A INVX1_LOC_140/A 0.01fF
C6195 NOR2X1_LOC_391/B NAND2X1_LOC_215/A 0.00fF
C6196 NOR2X1_LOC_78/Y INVX1_LOC_84/A 0.02fF
C6197 NOR2X1_LOC_329/B NOR2X1_LOC_109/Y 0.02fF
C6198 INVX1_LOC_25/Y NAND2X1_LOC_793/Y 0.00fF
C6199 INVX1_LOC_310/A NOR2X1_LOC_688/Y 0.01fF
C6200 NOR2X1_LOC_658/Y INVX1_LOC_96/Y 0.08fF
C6201 NAND2X1_LOC_561/a_36_24# INVX1_LOC_282/A 0.00fF
C6202 INVX1_LOC_230/Y NAND2X1_LOC_563/A 0.03fF
C6203 NAND2X1_LOC_802/A NAND2X1_LOC_798/a_36_24# 0.02fF
C6204 NAND2X1_LOC_814/a_36_24# INVX1_LOC_271/A 0.00fF
C6205 NAND2X1_LOC_533/a_36_24# INVX1_LOC_75/A 0.00fF
C6206 NAND2X1_LOC_35/Y NAND2X1_LOC_560/A 0.26fF
C6207 NAND2X1_LOC_796/B INVX1_LOC_90/A 0.00fF
C6208 NOR2X1_LOC_441/Y NOR2X1_LOC_366/B 0.10fF
C6209 NOR2X1_LOC_295/a_36_216# INVX1_LOC_71/A 0.00fF
C6210 INVX1_LOC_26/Y NAND2X1_LOC_642/Y 0.03fF
C6211 INVX1_LOC_91/A NOR2X1_LOC_383/B 0.20fF
C6212 NAND2X1_LOC_565/B NOR2X1_LOC_134/Y 0.01fF
C6213 NOR2X1_LOC_598/B NOR2X1_LOC_730/B 0.00fF
C6214 NOR2X1_LOC_309/Y NAND2X1_LOC_656/A 0.03fF
C6215 NAND2X1_LOC_47/a_36_24# GATE_662 0.00fF
C6216 INVX1_LOC_78/A INVX1_LOC_20/A 0.14fF
C6217 VDD NOR2X1_LOC_855/A 0.13fF
C6218 NAND2X1_LOC_740/Y NAND2X1_LOC_855/Y 0.00fF
C6219 NOR2X1_LOC_405/A NOR2X1_LOC_831/a_36_216# 0.01fF
C6220 NOR2X1_LOC_599/A NAND2X1_LOC_852/Y 0.05fF
C6221 INVX1_LOC_31/A NOR2X1_LOC_121/A 0.03fF
C6222 INVX1_LOC_256/A INVX1_LOC_279/A 0.12fF
C6223 INVX1_LOC_238/Y INVX1_LOC_241/A 0.09fF
C6224 NOR2X1_LOC_238/Y NOR2X1_LOC_52/B 0.03fF
C6225 INVX1_LOC_50/A NOR2X1_LOC_311/Y 0.22fF
C6226 INVX1_LOC_93/Y INVX1_LOC_181/A 0.00fF
C6227 NOR2X1_LOC_716/B NAND2X1_LOC_833/Y 0.00fF
C6228 NOR2X1_LOC_824/A NOR2X1_LOC_497/Y 0.04fF
C6229 INVX1_LOC_21/A NOR2X1_LOC_135/Y 0.01fF
C6230 INVX1_LOC_35/A INVX1_LOC_6/A 0.10fF
C6231 INVX1_LOC_14/Y NOR2X1_LOC_334/Y 0.10fF
C6232 NAND2X1_LOC_213/A NOR2X1_LOC_163/A 0.06fF
C6233 INVX1_LOC_174/A NAND2X1_LOC_148/a_36_24# 0.01fF
C6234 NAND2X1_LOC_11/Y NOR2X1_LOC_68/A 0.00fF
C6235 INVX1_LOC_45/A INVX1_LOC_208/Y 0.04fF
C6236 INVX1_LOC_172/A NOR2X1_LOC_629/B 0.00fF
C6237 NOR2X1_LOC_561/Y NOR2X1_LOC_276/Y -0.02fF
C6238 INVX1_LOC_2/A INVX1_LOC_24/A 0.29fF
C6239 INVX1_LOC_34/A NOR2X1_LOC_219/B 0.07fF
C6240 NOR2X1_LOC_848/Y NOR2X1_LOC_846/B 0.01fF
C6241 NOR2X1_LOC_382/Y INVX1_LOC_16/A 0.02fF
C6242 INVX1_LOC_58/A NOR2X1_LOC_43/Y 0.01fF
C6243 NOR2X1_LOC_168/a_36_216# NAND2X1_LOC_72/B 0.00fF
C6244 INVX1_LOC_34/A NAND2X1_LOC_483/Y 0.00fF
C6245 NAND2X1_LOC_773/a_36_24# INVX1_LOC_20/A 0.01fF
C6246 NOR2X1_LOC_388/Y NOR2X1_LOC_142/Y 0.10fF
C6247 INVX1_LOC_41/A INVX1_LOC_8/A 0.18fF
C6248 INVX1_LOC_290/A INVX1_LOC_30/A 0.25fF
C6249 NOR2X1_LOC_536/A NOR2X1_LOC_38/B 0.03fF
C6250 INVX1_LOC_50/A NOR2X1_LOC_164/Y 0.00fF
C6251 NOR2X1_LOC_226/A INVX1_LOC_24/A 0.10fF
C6252 INVX1_LOC_182/Y NOR2X1_LOC_348/Y 0.01fF
C6253 NAND2X1_LOC_738/B INVX1_LOC_11/Y 0.93fF
C6254 NOR2X1_LOC_189/A NAND2X1_LOC_722/A 0.09fF
C6255 INVX1_LOC_238/Y NOR2X1_LOC_298/Y 0.04fF
C6256 NOR2X1_LOC_134/Y NOR2X1_LOC_130/A 0.03fF
C6257 INVX1_LOC_64/A NOR2X1_LOC_187/a_36_216# 0.01fF
C6258 NOR2X1_LOC_820/A NOR2X1_LOC_516/B 0.04fF
C6259 INVX1_LOC_18/A INVX1_LOC_22/A 0.28fF
C6260 NAND2X1_LOC_811/Y GATE_811 0.03fF
C6261 NOR2X1_LOC_155/A NOR2X1_LOC_833/B 0.08fF
C6262 NAND2X1_LOC_342/Y INVX1_LOC_77/A 0.02fF
C6263 NAND2X1_LOC_574/A INVX1_LOC_29/A 0.07fF
C6264 NOR2X1_LOC_222/Y NOR2X1_LOC_208/Y 0.02fF
C6265 NAND2X1_LOC_647/B INVX1_LOC_9/A 0.04fF
C6266 NAND2X1_LOC_728/Y INVX1_LOC_22/A 0.07fF
C6267 NAND2X1_LOC_303/Y NAND2X1_LOC_863/A 0.14fF
C6268 INVX1_LOC_314/Y NOR2X1_LOC_191/A 0.39fF
C6269 NOR2X1_LOC_454/a_36_216# INVX1_LOC_191/Y 0.00fF
C6270 INVX1_LOC_49/A INVX1_LOC_143/A 0.03fF
C6271 NAND2X1_LOC_53/Y NOR2X1_LOC_736/Y 0.03fF
C6272 INVX1_LOC_21/A NOR2X1_LOC_147/A 0.03fF
C6273 NOR2X1_LOC_437/a_36_216# INVX1_LOC_208/A 0.00fF
C6274 INVX1_LOC_227/A INVX1_LOC_223/A 0.00fF
C6275 NOR2X1_LOC_657/B NOR2X1_LOC_678/A 0.15fF
C6276 NOR2X1_LOC_494/Y INVX1_LOC_282/A 0.01fF
C6277 INVX1_LOC_2/A NOR2X1_LOC_557/Y 0.08fF
C6278 INVX1_LOC_136/A NOR2X1_LOC_561/Y 0.11fF
C6279 INVX1_LOC_166/A D_GATE_662 0.02fF
C6280 INVX1_LOC_50/A INVX1_LOC_46/A 1.08fF
C6281 INVX1_LOC_136/A INVX1_LOC_7/A 0.36fF
C6282 INVX1_LOC_164/Y NOR2X1_LOC_716/B 0.04fF
C6283 NOR2X1_LOC_398/Y INVX1_LOC_8/A 0.02fF
C6284 NOR2X1_LOC_574/A NOR2X1_LOC_52/B 0.17fF
C6285 INVX1_LOC_159/A NAND2X1_LOC_660/Y -0.02fF
C6286 INVX1_LOC_208/Y INVX1_LOC_71/A 0.15fF
C6287 NOR2X1_LOC_637/Y INVX1_LOC_22/A 0.00fF
C6288 INVX1_LOC_77/Y NOR2X1_LOC_638/Y 0.03fF
C6289 NOR2X1_LOC_226/A NOR2X1_LOC_557/Y 0.07fF
C6290 INVX1_LOC_256/A INVX1_LOC_182/Y 0.03fF
C6291 NOR2X1_LOC_655/B NOR2X1_LOC_388/Y 0.03fF
C6292 NAND2X1_LOC_748/a_36_24# INVX1_LOC_48/A 0.00fF
C6293 NOR2X1_LOC_570/A INVX1_LOC_94/A 0.01fF
C6294 NOR2X1_LOC_361/B NOR2X1_LOC_74/A 0.18fF
C6295 NAND2X1_LOC_391/a_36_24# INVX1_LOC_234/A 0.00fF
C6296 NAND2X1_LOC_545/a_36_24# NOR2X1_LOC_355/A 0.00fF
C6297 INVX1_LOC_35/Y INVX1_LOC_15/A 0.07fF
C6298 INVX1_LOC_172/A INVX1_LOC_22/A 0.03fF
C6299 NOR2X1_LOC_726/Y INVX1_LOC_85/Y 0.01fF
C6300 NOR2X1_LOC_720/B NAND2X1_LOC_338/B 0.04fF
C6301 NOR2X1_LOC_717/B NOR2X1_LOC_457/B 0.02fF
C6302 INVX1_LOC_50/A NOR2X1_LOC_766/Y 0.01fF
C6303 NOR2X1_LOC_589/A NOR2X1_LOC_152/Y 0.07fF
C6304 INVX1_LOC_91/A NOR2X1_LOC_463/a_36_216# 0.00fF
C6305 INVX1_LOC_33/A INVX1_LOC_232/A 0.16fF
C6306 NOR2X1_LOC_175/A NOR2X1_LOC_538/Y 0.03fF
C6307 INVX1_LOC_234/A D_INPUT_2 0.00fF
C6308 NOR2X1_LOC_589/A INVX1_LOC_113/Y 0.04fF
C6309 NAND2X1_LOC_722/A NOR2X1_LOC_482/Y 0.01fF
C6310 NOR2X1_LOC_631/B INVX1_LOC_50/Y 0.00fF
C6311 NAND2X1_LOC_112/Y NOR2X1_LOC_172/Y 0.30fF
C6312 NOR2X1_LOC_639/Y INVX1_LOC_118/A 0.06fF
C6313 NAND2X1_LOC_72/Y INVX1_LOC_46/A 0.91fF
C6314 NOR2X1_LOC_516/B INVX1_LOC_315/A 0.03fF
C6315 NAND2X1_LOC_114/B INPUT_0 0.04fF
C6316 NOR2X1_LOC_160/B NOR2X1_LOC_368/A 0.45fF
C6317 INVX1_LOC_2/A INVX1_LOC_143/A 0.10fF
C6318 INVX1_LOC_36/A NOR2X1_LOC_329/B 0.16fF
C6319 NOR2X1_LOC_142/Y NAND2X1_LOC_479/Y 0.07fF
C6320 NOR2X1_LOC_820/Y INVX1_LOC_4/Y 0.14fF
C6321 INVX1_LOC_280/A NAND2X1_LOC_215/A -0.03fF
C6322 NAND2X1_LOC_324/a_36_24# INVX1_LOC_91/A 0.01fF
C6323 NOR2X1_LOC_804/B INVX1_LOC_220/Y 0.18fF
C6324 INVX1_LOC_34/A NOR2X1_LOC_789/A 0.01fF
C6325 NOR2X1_LOC_383/Y INVX1_LOC_33/A 0.19fF
C6326 INVX1_LOC_226/Y INVX1_LOC_60/Y 0.34fF
C6327 NOR2X1_LOC_38/B NOR2X1_LOC_649/B 0.03fF
C6328 INVX1_LOC_24/A NAND2X1_LOC_648/A 0.01fF
C6329 NOR2X1_LOC_106/Y NOR2X1_LOC_106/A 0.02fF
C6330 INVX1_LOC_21/A NAND2X1_LOC_1/Y 0.14fF
C6331 NOR2X1_LOC_226/A INVX1_LOC_143/A 0.09fF
C6332 NOR2X1_LOC_38/B INVX1_LOC_3/A 0.10fF
C6333 NOR2X1_LOC_229/a_36_216# INVX1_LOC_266/Y 0.00fF
C6334 INVX1_LOC_24/A INPUT_1 1.23fF
C6335 INVX1_LOC_268/A NOR2X1_LOC_52/B 0.01fF
C6336 NOR2X1_LOC_418/a_36_216# INVX1_LOC_191/Y 0.00fF
C6337 INVX1_LOC_72/A INVX1_LOC_302/A 0.08fF
C6338 INVX1_LOC_299/A INVX1_LOC_93/Y 0.00fF
C6339 INVX1_LOC_33/A NOR2X1_LOC_366/Y 0.02fF
C6340 NAND2X1_LOC_563/Y INVX1_LOC_13/A 0.20fF
C6341 INVX1_LOC_50/Y INVX1_LOC_37/A 0.15fF
C6342 NOR2X1_LOC_773/Y NAND2X1_LOC_850/Y 0.02fF
C6343 INVX1_LOC_34/A NAND2X1_LOC_656/Y 0.09fF
C6344 INVX1_LOC_75/A INVX1_LOC_205/A 0.01fF
C6345 NAND2X1_LOC_74/B INVX1_LOC_127/Y 0.03fF
C6346 INVX1_LOC_135/A NOR2X1_LOC_340/Y 0.01fF
C6347 NOR2X1_LOC_244/B INVX1_LOC_120/Y 0.24fF
C6348 NOR2X1_LOC_716/B NOR2X1_LOC_76/A 0.00fF
C6349 NOR2X1_LOC_151/Y NOR2X1_LOC_457/B 0.02fF
C6350 NAND2X1_LOC_574/A NOR2X1_LOC_33/Y 0.06fF
C6351 NOR2X1_LOC_19/B D_INPUT_2 0.15fF
C6352 NOR2X1_LOC_474/A INVX1_LOC_175/Y 0.24fF
C6353 D_INPUT_0 NOR2X1_LOC_4/a_36_216# 0.00fF
C6354 INVX1_LOC_11/A INVX1_LOC_95/Y 1.12fF
C6355 INVX1_LOC_307/A INVX1_LOC_29/Y 0.00fF
C6356 NOR2X1_LOC_321/Y NOR2X1_LOC_65/a_36_216# 0.00fF
C6357 NOR2X1_LOC_155/A NOR2X1_LOC_125/Y 0.07fF
C6358 NOR2X1_LOC_420/Y NOR2X1_LOC_536/A 0.04fF
C6359 INVX1_LOC_40/A INVX1_LOC_232/A 0.10fF
C6360 INVX1_LOC_313/Y INVX1_LOC_155/Y 0.21fF
C6361 INVX1_LOC_45/A NOR2X1_LOC_501/B 0.01fF
C6362 INVX1_LOC_90/A NAND2X1_LOC_139/A 0.02fF
C6363 NOR2X1_LOC_226/A NAND2X1_LOC_552/a_36_24# 0.01fF
C6364 NOR2X1_LOC_488/Y NAND2X1_LOC_543/Y 0.01fF
C6365 D_INPUT_1 NOR2X1_LOC_216/B 0.10fF
C6366 INVX1_LOC_266/A INVX1_LOC_37/A 0.49fF
C6367 NAND2X1_LOC_670/a_36_24# INVX1_LOC_123/A 0.01fF
C6368 INVX1_LOC_2/A NAND2X1_LOC_783/A 0.45fF
C6369 NOR2X1_LOC_775/Y INVX1_LOC_33/A 0.01fF
C6370 NOR2X1_LOC_52/B NOR2X1_LOC_367/a_36_216# 0.00fF
C6371 NAND2X1_LOC_231/Y NAND2X1_LOC_656/Y 0.10fF
C6372 NOR2X1_LOC_598/B NOR2X1_LOC_155/A 0.27fF
C6373 NOR2X1_LOC_524/Y NOR2X1_LOC_318/B 0.03fF
C6374 INVX1_LOC_35/A INVX1_LOC_131/Y 0.27fF
C6375 INVX1_LOC_63/A NAND2X1_LOC_99/A 0.07fF
C6376 INVX1_LOC_2/A NOR2X1_LOC_130/A 0.07fF
C6377 INVX1_LOC_4/A INVX1_LOC_42/A 0.10fF
C6378 NOR2X1_LOC_576/B NOR2X1_LOC_504/Y 0.01fF
C6379 INPUT_5 NOR2X1_LOC_44/a_36_216# 0.02fF
C6380 INVX1_LOC_77/A INVX1_LOC_67/Y 0.01fF
C6381 INVX1_LOC_11/A NOR2X1_LOC_305/Y 0.01fF
C6382 NOR2X1_LOC_669/Y INVX1_LOC_33/Y 0.01fF
C6383 NOR2X1_LOC_716/B INVX1_LOC_73/A 0.01fF
C6384 NOR2X1_LOC_655/B INVX1_LOC_135/A 0.03fF
C6385 INVX1_LOC_200/Y INVX1_LOC_119/Y 0.17fF
C6386 NOR2X1_LOC_250/Y VDD 0.18fF
C6387 NOR2X1_LOC_89/A INVX1_LOC_271/Y 0.07fF
C6388 NOR2X1_LOC_226/A NOR2X1_LOC_130/A 1.17fF
C6389 INVX1_LOC_312/Y NAND2X1_LOC_649/B 0.02fF
C6390 NOR2X1_LOC_690/Y INVX1_LOC_22/A 0.00fF
C6391 NOR2X1_LOC_202/Y NOR2X1_LOC_142/Y 0.09fF
C6392 NAND2X1_LOC_454/Y INVX1_LOC_109/Y 0.02fF
C6393 NOR2X1_LOC_468/Y NOR2X1_LOC_536/A 0.21fF
C6394 NOR2X1_LOC_717/B NAND2X1_LOC_372/a_36_24# 0.00fF
C6395 INVX1_LOC_25/A NAND2X1_LOC_475/Y 0.00fF
C6396 INVX1_LOC_245/Y VDD 0.79fF
C6397 INVX1_LOC_177/A NOR2X1_LOC_356/A 0.04fF
C6398 NOR2X1_LOC_232/a_36_216# NAND2X1_LOC_849/B 0.00fF
C6399 NAND2X1_LOC_860/A INVX1_LOC_84/A 0.12fF
C6400 NOR2X1_LOC_355/A NOR2X1_LOC_500/Y 0.12fF
C6401 NOR2X1_LOC_512/Y INVX1_LOC_91/A 0.02fF
C6402 INVX1_LOC_71/A NOR2X1_LOC_501/B 0.00fF
C6403 NOR2X1_LOC_208/Y NOR2X1_LOC_66/a_36_216# 0.00fF
C6404 NOR2X1_LOC_187/Y NOR2X1_LOC_331/B 0.02fF
C6405 INVX1_LOC_72/A NAND2X1_LOC_271/a_36_24# 0.00fF
C6406 NAND2X1_LOC_632/B INVX1_LOC_309/A 0.02fF
C6407 NOR2X1_LOC_216/B NOR2X1_LOC_652/Y 0.18fF
C6408 INVX1_LOC_1/Y INVX1_LOC_66/A 0.01fF
C6409 INVX1_LOC_249/A NOR2X1_LOC_144/a_36_216# 0.00fF
C6410 NOR2X1_LOC_763/Y NAND2X1_LOC_662/Y 0.05fF
C6411 NAND2X1_LOC_562/B INVX1_LOC_282/A 0.04fF
C6412 NOR2X1_LOC_458/B NOR2X1_LOC_644/A 0.01fF
C6413 INVX1_LOC_230/Y INVX1_LOC_12/Y 0.00fF
C6414 NOR2X1_LOC_151/Y NOR2X1_LOC_182/a_36_216# 0.00fF
C6415 INVX1_LOC_138/A NAND2X1_LOC_206/Y 0.06fF
C6416 INVX1_LOC_124/Y VDD 0.49fF
C6417 INVX1_LOC_157/A INVX1_LOC_279/A 0.10fF
C6418 NAND2X1_LOC_276/Y INVX1_LOC_48/A 0.08fF
C6419 NOR2X1_LOC_186/Y NOR2X1_LOC_841/A 0.00fF
C6420 INVX1_LOC_136/A INVX1_LOC_76/A 0.33fF
C6421 INVX1_LOC_299/A NOR2X1_LOC_856/A 0.15fF
C6422 NOR2X1_LOC_554/B INVX1_LOC_20/A 0.08fF
C6423 NAND2X1_LOC_565/B INPUT_1 0.12fF
C6424 D_INPUT_1 NAND2X1_LOC_82/a_36_24# 0.00fF
C6425 INVX1_LOC_78/A INVX1_LOC_4/A 3.07fF
C6426 INVX1_LOC_33/A NOR2X1_LOC_685/A 0.01fF
C6427 INVX1_LOC_177/A NOR2X1_LOC_74/A 0.08fF
C6428 INVX1_LOC_12/A INVX1_LOC_29/Y 0.03fF
C6429 NOR2X1_LOC_468/Y NAND2X1_LOC_93/B 0.67fF
C6430 NOR2X1_LOC_355/A INVX1_LOC_10/A 0.10fF
C6431 INVX1_LOC_33/A INVX1_LOC_186/A 0.03fF
C6432 INVX1_LOC_119/Y NOR2X1_LOC_406/A 0.02fF
C6433 NOR2X1_LOC_389/A NOR2X1_LOC_536/A 0.03fF
C6434 NOR2X1_LOC_168/B INPUT_0 0.03fF
C6435 NOR2X1_LOC_791/A VDD 0.00fF
C6436 NOR2X1_LOC_409/Y NOR2X1_LOC_505/Y 0.06fF
C6437 NOR2X1_LOC_68/A NOR2X1_LOC_857/A 0.10fF
C6438 INVX1_LOC_277/A INVX1_LOC_117/A 0.08fF
C6439 NAND2X1_LOC_579/A NOR2X1_LOC_491/Y 0.14fF
C6440 INVX1_LOC_315/Y INVX1_LOC_315/A 0.03fF
C6441 NAND2X1_LOC_573/Y NOR2X1_LOC_841/A 0.34fF
C6442 INVX1_LOC_39/A NOR2X1_LOC_813/a_36_216# 0.00fF
C6443 INVX1_LOC_135/A NOR2X1_LOC_99/B 0.07fF
C6444 INVX1_LOC_286/Y NAND2X1_LOC_848/A 0.23fF
C6445 NAND2X1_LOC_571/B INVX1_LOC_284/A 0.07fF
C6446 NOR2X1_LOC_778/B NAND2X1_LOC_496/a_36_24# 0.00fF
C6447 NOR2X1_LOC_147/B NOR2X1_LOC_78/A 0.00fF
C6448 INVX1_LOC_14/A NAND2X1_LOC_647/a_36_24# 0.01fF
C6449 INVX1_LOC_35/A NOR2X1_LOC_633/A 0.01fF
C6450 NAND2X1_LOC_363/B NAND2X1_LOC_245/a_36_24# 0.00fF
C6451 NAND2X1_LOC_198/B NAND2X1_LOC_287/B 0.10fF
C6452 NOR2X1_LOC_637/A NAND2X1_LOC_453/A 0.04fF
C6453 NAND2X1_LOC_537/Y NOR2X1_LOC_88/Y 0.07fF
C6454 INVX1_LOC_222/Y INVX1_LOC_63/A 0.03fF
C6455 NOR2X1_LOC_598/B NOR2X1_LOC_833/B 0.16fF
C6456 NOR2X1_LOC_218/Y NOR2X1_LOC_216/Y 0.03fF
C6457 INVX1_LOC_64/A INVX1_LOC_263/Y 0.01fF
C6458 NOR2X1_LOC_392/B NOR2X1_LOC_78/A 0.01fF
C6459 NOR2X1_LOC_562/a_36_216# NOR2X1_LOC_486/Y 0.02fF
C6460 NAND2X1_LOC_800/Y NAND2X1_LOC_648/A 0.31fF
C6461 NOR2X1_LOC_65/B INVX1_LOC_4/A 0.03fF
C6462 NAND2X1_LOC_35/Y INVX1_LOC_29/A 0.07fF
C6463 NOR2X1_LOC_591/a_36_216# INVX1_LOC_91/A 0.01fF
C6464 NOR2X1_LOC_178/Y NAND2X1_LOC_74/B 0.01fF
C6465 NOR2X1_LOC_152/Y INVX1_LOC_20/A 0.10fF
C6466 NOR2X1_LOC_593/Y INVX1_LOC_95/Y 0.00fF
C6467 NOR2X1_LOC_15/Y NOR2X1_LOC_697/Y 0.03fF
C6468 NAND2X1_LOC_743/a_36_24# NAND2X1_LOC_782/B 0.01fF
C6469 NOR2X1_LOC_717/B NOR2X1_LOC_180/B 0.03fF
C6470 NOR2X1_LOC_560/A NOR2X1_LOC_99/B 0.02fF
C6471 NOR2X1_LOC_130/A INPUT_1 0.12fF
C6472 INVX1_LOC_24/A NAND2X1_LOC_605/a_36_24# 0.00fF
C6473 INVX1_LOC_39/A NAND2X1_LOC_773/B 0.05fF
C6474 NOR2X1_LOC_239/a_36_216# INVX1_LOC_38/A 0.02fF
C6475 NOR2X1_LOC_570/B INVX1_LOC_247/A 0.02fF
C6476 NAND2X1_LOC_81/B INVX1_LOC_306/Y 0.03fF
C6477 NOR2X1_LOC_160/B NOR2X1_LOC_660/a_36_216# 0.02fF
C6478 INVX1_LOC_64/A INVX1_LOC_42/A 0.35fF
C6479 INVX1_LOC_105/A INVX1_LOC_46/A 0.10fF
C6480 NOR2X1_LOC_389/A NAND2X1_LOC_93/B 0.00fF
C6481 NAND2X1_LOC_364/A NOR2X1_LOC_114/a_36_216# 0.00fF
C6482 INVX1_LOC_150/Y NOR2X1_LOC_831/B 0.31fF
C6483 INVX1_LOC_1/A NAND2X1_LOC_475/Y 0.01fF
C6484 NAND2X1_LOC_860/A INVX1_LOC_15/A 0.03fF
C6485 NOR2X1_LOC_34/B NAND2X1_LOC_207/Y 0.06fF
C6486 NOR2X1_LOC_548/A INVX1_LOC_22/A 0.09fF
C6487 NAND2X1_LOC_537/Y INVX1_LOC_84/A 1.30fF
C6488 NOR2X1_LOC_168/A INVX1_LOC_91/A 0.05fF
C6489 INVX1_LOC_62/Y NOR2X1_LOC_536/A 0.07fF
C6490 NOR2X1_LOC_52/B INVX1_LOC_95/Y 0.01fF
C6491 NOR2X1_LOC_540/B NOR2X1_LOC_180/Y 0.02fF
C6492 NOR2X1_LOC_632/Y INVX1_LOC_311/A 0.01fF
C6493 NOR2X1_LOC_389/A NAND2X1_LOC_425/Y 0.02fF
C6494 NOR2X1_LOC_355/A NAND2X1_LOC_132/a_36_24# 0.00fF
C6495 NOR2X1_LOC_74/A NAND2X1_LOC_573/A 0.02fF
C6496 INVX1_LOC_311/Y INVX1_LOC_85/Y 0.94fF
C6497 NOR2X1_LOC_121/Y VDD 0.25fF
C6498 NAND2X1_LOC_656/Y INPUT_0 0.08fF
C6499 INVX1_LOC_138/A NOR2X1_LOC_297/A 0.00fF
C6500 INVX1_LOC_77/A NOR2X1_LOC_862/a_36_216# 0.01fF
C6501 NOR2X1_LOC_828/B NOR2X1_LOC_732/a_36_216# 0.02fF
C6502 D_INPUT_0 NOR2X1_LOC_721/Y 0.37fF
C6503 NAND2X1_LOC_170/A INVX1_LOC_91/A 0.03fF
C6504 NOR2X1_LOC_172/Y NOR2X1_LOC_60/Y 0.01fF
C6505 INVX1_LOC_24/A INVX1_LOC_118/A 1.53fF
C6506 NOR2X1_LOC_718/B INVX1_LOC_14/Y 0.06fF
C6507 NOR2X1_LOC_6/B INVX1_LOC_37/A 3.90fF
C6508 INVX1_LOC_18/A NOR2X1_LOC_88/A 0.02fF
C6509 NAND2X1_LOC_325/a_36_24# NAND2X1_LOC_808/A 0.00fF
C6510 NOR2X1_LOC_285/B INVX1_LOC_117/A 0.01fF
C6511 NAND2X1_LOC_119/a_36_24# NOR2X1_LOC_271/Y 0.00fF
C6512 NOR2X1_LOC_151/Y NOR2X1_LOC_180/B 0.02fF
C6513 INVX1_LOC_90/A NAND2X1_LOC_840/Y 0.01fF
C6514 NAND2X1_LOC_773/Y NOR2X1_LOC_89/A 0.03fF
C6515 NAND2X1_LOC_269/a_36_24# INVX1_LOC_306/Y 0.06fF
C6516 NAND2X1_LOC_841/A INVX1_LOC_199/A 0.12fF
C6517 INVX1_LOC_215/A NOR2X1_LOC_45/B 0.18fF
C6518 NOR2X1_LOC_315/Y NAND2X1_LOC_721/A 0.03fF
C6519 INVX1_LOC_64/A INVX1_LOC_78/A 0.24fF
C6520 INVX1_LOC_17/A NOR2X1_LOC_340/A 0.07fF
C6521 NOR2X1_LOC_340/Y INVX1_LOC_280/A 0.02fF
C6522 NOR2X1_LOC_596/A NAND2X1_LOC_93/B 0.20fF
C6523 INVX1_LOC_306/Y INVX1_LOC_4/Y 0.01fF
C6524 INVX1_LOC_15/A NAND2X1_LOC_473/A 0.23fF
C6525 INVX1_LOC_140/A INVX1_LOC_282/A 0.03fF
C6526 NAND2X1_LOC_860/Y INVX1_LOC_20/A 0.02fF
C6527 INVX1_LOC_52/A INVX1_LOC_139/A 0.01fF
C6528 NOR2X1_LOC_596/A NAND2X1_LOC_425/Y 0.01fF
C6529 NOR2X1_LOC_373/Y NOR2X1_LOC_45/B 0.07fF
C6530 INVX1_LOC_50/Y NAND2X1_LOC_72/B 0.03fF
C6531 NAND2X1_LOC_660/Y NOR2X1_LOC_56/Y 0.07fF
C6532 INVX1_LOC_58/A NAND2X1_LOC_784/A 0.00fF
C6533 NOR2X1_LOC_285/Y INVX1_LOC_26/Y 0.01fF
C6534 INVX1_LOC_57/Y INVX1_LOC_203/A 0.00fF
C6535 NAND2X1_LOC_360/B INVX1_LOC_117/A 0.05fF
C6536 NOR2X1_LOC_65/B INVX1_LOC_64/A 0.02fF
C6537 INVX1_LOC_233/A INVX1_LOC_50/A 0.02fF
C6538 NOR2X1_LOC_456/Y INVX1_LOC_23/A 1.95fF
C6539 INVX1_LOC_35/A INVX1_LOC_270/A 0.07fF
C6540 INVX1_LOC_271/A NOR2X1_LOC_678/A 0.03fF
C6541 NOR2X1_LOC_769/B NOR2X1_LOC_598/B 0.03fF
C6542 INVX1_LOC_280/Y NOR2X1_LOC_690/a_36_216# 0.00fF
C6543 INVX1_LOC_49/A NOR2X1_LOC_197/B 0.12fF
C6544 NAND2X1_LOC_727/Y VDD 0.01fF
C6545 INVX1_LOC_90/A NOR2X1_LOC_78/A 0.17fF
C6546 INVX1_LOC_43/Y INVX1_LOC_42/A 0.02fF
C6547 NOR2X1_LOC_689/Y NAND2X1_LOC_725/A 0.05fF
C6548 INVX1_LOC_27/A NOR2X1_LOC_34/Y 0.03fF
C6549 INVX1_LOC_5/A NOR2X1_LOC_720/A 0.02fF
C6550 INVX1_LOC_18/A INVX1_LOC_186/Y 0.03fF
C6551 NOR2X1_LOC_655/B INVX1_LOC_280/A 0.10fF
C6552 NOR2X1_LOC_480/A INVX1_LOC_203/A 0.00fF
C6553 NOR2X1_LOC_389/B NOR2X1_LOC_78/A 0.07fF
C6554 NAND2X1_LOC_660/Y VDD 0.10fF
C6555 INVX1_LOC_278/A NAND2X1_LOC_860/A 0.22fF
C6556 NAND2X1_LOC_656/A INVX1_LOC_63/A 0.56fF
C6557 INVX1_LOC_77/A INVX1_LOC_285/A 0.00fF
C6558 INVX1_LOC_266/A NAND2X1_LOC_72/B 0.08fF
C6559 INVX1_LOC_289/Y INVX1_LOC_94/Y 0.03fF
C6560 NOR2X1_LOC_91/Y INVX1_LOC_19/A 0.00fF
C6561 NAND2X1_LOC_464/Y INVX1_LOC_35/Y 0.06fF
C6562 NOR2X1_LOC_356/A INVX1_LOC_65/A 0.10fF
C6563 INVX1_LOC_16/A INVX1_LOC_202/Y 0.10fF
C6564 INVX1_LOC_77/A NOR2X1_LOC_814/A 0.72fF
C6565 INVX1_LOC_50/A NOR2X1_LOC_798/A 0.03fF
C6566 NAND2X1_LOC_861/Y INVX1_LOC_20/A 0.08fF
C6567 INVX1_LOC_5/A NOR2X1_LOC_629/A 0.01fF
C6568 INVX1_LOC_64/A INVX1_LOC_152/Y 0.17fF
C6569 NAND2X1_LOC_787/B NOR2X1_LOC_485/Y 0.19fF
C6570 D_INPUT_0 VDD 1.55fF
C6571 INVX1_LOC_24/A NAND2X1_LOC_63/Y 0.07fF
C6572 INVX1_LOC_11/A INVX1_LOC_271/Y 0.07fF
C6573 NAND2X1_LOC_348/A NOR2X1_LOC_78/A 0.08fF
C6574 NOR2X1_LOC_13/Y INVX1_LOC_49/Y 0.17fF
C6575 INVX1_LOC_35/A NOR2X1_LOC_109/Y 0.11fF
C6576 NAND2X1_LOC_112/Y INVX1_LOC_38/A 0.03fF
C6577 INVX1_LOC_191/A NAND2X1_LOC_450/a_36_24# 0.01fF
C6578 INVX1_LOC_94/A INVX1_LOC_29/A 0.16fF
C6579 INVX1_LOC_50/A NAND2X1_LOC_703/Y 0.01fF
C6580 NAND2X1_LOC_11/Y NAND2X1_LOC_430/a_36_24# 0.00fF
C6581 INVX1_LOC_21/A NOR2X1_LOC_452/A 0.02fF
C6582 INVX1_LOC_189/Y NAND2X1_LOC_93/B 0.03fF
C6583 INVX1_LOC_166/A INVX1_LOC_239/A 2.28fF
C6584 NOR2X1_LOC_91/A NAND2X1_LOC_561/B 0.03fF
C6585 NAND2X1_LOC_624/B INVX1_LOC_5/A 0.03fF
C6586 INVX1_LOC_30/A NOR2X1_LOC_467/A 0.40fF
C6587 NAND2X1_LOC_35/Y NOR2X1_LOC_291/a_36_216# 0.01fF
C6588 INVX1_LOC_124/A INVX1_LOC_285/A 0.20fF
C6589 INVX1_LOC_189/Y NAND2X1_LOC_425/Y 0.03fF
C6590 NAND2X1_LOC_763/B NOR2X1_LOC_467/A 0.69fF
C6591 NOR2X1_LOC_238/Y NAND2X1_LOC_254/Y 0.00fF
C6592 NOR2X1_LOC_156/A INVX1_LOC_37/A 0.01fF
C6593 NOR2X1_LOC_516/B NOR2X1_LOC_660/a_36_216# 0.00fF
C6594 NOR2X1_LOC_636/B NOR2X1_LOC_635/B 0.08fF
C6595 NOR2X1_LOC_82/A INVX1_LOC_181/A 0.04fF
C6596 INVX1_LOC_108/Y NAND2X1_LOC_473/A 0.09fF
C6597 NAND2X1_LOC_22/a_36_24# INPUT_7 0.00fF
C6598 INVX1_LOC_124/A NOR2X1_LOC_814/A 0.04fF
C6599 NOR2X1_LOC_557/Y NAND2X1_LOC_63/Y 0.08fF
C6600 NOR2X1_LOC_99/B INVX1_LOC_280/A 0.11fF
C6601 NOR2X1_LOC_514/a_36_216# NAND2X1_LOC_82/Y 0.00fF
C6602 INVX1_LOC_5/A NOR2X1_LOC_849/A 0.03fF
C6603 NAND2X1_LOC_624/B INVX1_LOC_178/A 0.02fF
C6604 NOR2X1_LOC_554/B INVX1_LOC_4/A 0.09fF
C6605 NAND2X1_LOC_51/B NAND2X1_LOC_1/Y 0.01fF
C6606 NAND2X1_LOC_783/A INVX1_LOC_118/A 0.19fF
C6607 NOR2X1_LOC_433/A NAND2X1_LOC_806/a_36_24# 0.01fF
C6608 INVX1_LOC_13/Y NOR2X1_LOC_291/Y 0.14fF
C6609 INVX1_LOC_181/Y INVX1_LOC_32/A 0.10fF
C6610 INVX1_LOC_163/A NOR2X1_LOC_660/Y 0.33fF
C6611 NOR2X1_LOC_130/A INVX1_LOC_118/A 0.18fF
C6612 NOR2X1_LOC_74/A NAND2X1_LOC_267/B 0.00fF
C6613 INVX1_LOC_290/A INVX1_LOC_113/A 0.04fF
C6614 NOR2X1_LOC_665/A NAND2X1_LOC_792/a_36_24# 0.00fF
C6615 NAND2X1_LOC_67/Y NOR2X1_LOC_665/Y 0.33fF
C6616 INVX1_LOC_30/A INVX1_LOC_116/Y 0.00fF
C6617 NOR2X1_LOC_272/Y NAND2X1_LOC_474/Y 0.10fF
C6618 NOR2X1_LOC_9/Y NAND2X1_LOC_267/B 0.01fF
C6619 NOR2X1_LOC_74/a_36_216# INVX1_LOC_117/A 0.00fF
C6620 NOR2X1_LOC_456/Y NAND2X1_LOC_179/a_36_24# 0.02fF
C6621 INVX1_LOC_143/A NAND2X1_LOC_63/Y 0.02fF
C6622 NOR2X1_LOC_106/Y NOR2X1_LOC_334/Y 0.03fF
C6623 INVX1_LOC_14/A NOR2X1_LOC_81/Y 0.02fF
C6624 NOR2X1_LOC_791/Y INVX1_LOC_1/A 0.41fF
C6625 INVX1_LOC_298/Y INVX1_LOC_94/A 0.02fF
C6626 INVX1_LOC_24/A NOR2X1_LOC_631/Y 0.12fF
C6627 INPUT_5 NAND2X1_LOC_30/a_36_24# 0.01fF
C6628 INVX1_LOC_25/A INVX1_LOC_30/A 0.07fF
C6629 INVX1_LOC_1/A NAND2X1_LOC_63/a_36_24# 0.01fF
C6630 INVX1_LOC_220/Y INVX1_LOC_63/A 0.03fF
C6631 INVX1_LOC_96/A INVX1_LOC_37/A 0.08fF
C6632 NOR2X1_LOC_91/A INVX1_LOC_300/Y 2.46fF
C6633 INVX1_LOC_67/Y INVX1_LOC_9/A 0.01fF
C6634 INVX1_LOC_28/A INVX1_LOC_180/Y 0.01fF
C6635 NOR2X1_LOC_593/Y INVX1_LOC_271/Y 0.07fF
C6636 NAND2X1_LOC_850/Y INVX1_LOC_42/A 0.07fF
C6637 INVX1_LOC_14/A NOR2X1_LOC_611/a_36_216# 0.01fF
C6638 INVX1_LOC_58/A NOR2X1_LOC_194/a_36_216# 0.00fF
C6639 NOR2X1_LOC_360/Y INVX1_LOC_57/A 0.10fF
C6640 INVX1_LOC_121/A NOR2X1_LOC_258/Y 0.09fF
C6641 NAND2X1_LOC_190/Y NOR2X1_LOC_348/Y 0.17fF
C6642 INVX1_LOC_14/A NOR2X1_LOC_140/A 0.02fF
C6643 INVX1_LOC_35/A INVX1_LOC_36/A 0.06fF
C6644 NAND2X1_LOC_553/A INVX1_LOC_61/Y 0.00fF
C6645 NOR2X1_LOC_443/Y INVX1_LOC_303/A 0.03fF
C6646 NOR2X1_LOC_454/Y NAND2X1_LOC_803/B 0.04fF
C6647 NOR2X1_LOC_759/Y INVX1_LOC_23/A 0.03fF
C6648 D_GATE_741 INVX1_LOC_198/A 0.59fF
C6649 INVX1_LOC_157/A NAND2X1_LOC_433/a_36_24# 0.00fF
C6650 INVX1_LOC_202/A INVX1_LOC_23/A 0.52fF
C6651 NOR2X1_LOC_78/A INVX1_LOC_38/A 0.07fF
C6652 D_INPUT_1 NOR2X1_LOC_303/Y 0.07fF
C6653 NAND2X1_LOC_35/Y NAND2X1_LOC_634/Y 0.02fF
C6654 INVX1_LOC_279/A NOR2X1_LOC_89/A 0.24fF
C6655 INVX1_LOC_5/A INVX1_LOC_142/A 0.02fF
C6656 INVX1_LOC_215/Y NAND2X1_LOC_326/A 0.29fF
C6657 INVX1_LOC_299/A INVX1_LOC_134/A 0.94fF
C6658 INVX1_LOC_17/A INVX1_LOC_103/A 0.09fF
C6659 NAND2X1_LOC_231/Y INVX1_LOC_128/Y 0.14fF
C6660 INVX1_LOC_172/Y INVX1_LOC_15/A 0.00fF
C6661 INVX1_LOC_174/Y NOR2X1_LOC_460/A 0.09fF
C6662 NOR2X1_LOC_405/A NOR2X1_LOC_114/a_36_216# 0.01fF
C6663 INVX1_LOC_256/A NAND2X1_LOC_190/Y 0.10fF
C6664 NAND2X1_LOC_214/Y INPUT_3 0.01fF
C6665 NOR2X1_LOC_550/B INVX1_LOC_23/A 0.01fF
C6666 NOR2X1_LOC_355/A INVX1_LOC_12/A 0.07fF
C6667 INVX1_LOC_14/A NOR2X1_LOC_530/Y 0.03fF
C6668 NOR2X1_LOC_740/Y D_GATE_741 0.03fF
C6669 NOR2X1_LOC_329/B INVX1_LOC_63/A 0.08fF
C6670 INVX1_LOC_249/A NOR2X1_LOC_678/A 0.02fF
C6671 NOR2X1_LOC_690/A NAND2X1_LOC_464/B 0.01fF
C6672 NOR2X1_LOC_45/B INVX1_LOC_54/A 0.69fF
C6673 INVX1_LOC_32/Y INVX1_LOC_32/A 0.01fF
C6674 NOR2X1_LOC_682/Y VDD 0.19fF
C6675 NAND2X1_LOC_850/Y INVX1_LOC_78/A 0.07fF
C6676 NOR2X1_LOC_536/A NAND2X1_LOC_655/B 0.01fF
C6677 NOR2X1_LOC_552/Y NOR2X1_LOC_445/B 0.00fF
C6678 NOR2X1_LOC_471/Y INVX1_LOC_103/A 0.10fF
C6679 NAND2X1_LOC_564/A NAND2X1_LOC_569/A 0.12fF
C6680 INVX1_LOC_6/Y NOR2X1_LOC_678/A 0.01fF
C6681 NAND2X1_LOC_180/a_36_24# INVX1_LOC_181/A 0.00fF
C6682 NAND2X1_LOC_552/A INVX1_LOC_41/Y 0.21fF
C6683 INVX1_LOC_35/A NOR2X1_LOC_237/Y 0.07fF
C6684 NOR2X1_LOC_689/Y NAND2X1_LOC_308/Y 0.50fF
C6685 INVX1_LOC_64/A NOR2X1_LOC_152/Y 0.30fF
C6686 VDD NOR2X1_LOC_859/Y 0.12fF
C6687 NOR2X1_LOC_382/Y INVX1_LOC_48/Y 0.00fF
C6688 NOR2X1_LOC_792/B INVX1_LOC_57/A 0.00fF
C6689 INVX1_LOC_14/Y NAND2X1_LOC_472/Y 0.10fF
C6690 D_INPUT_1 NOR2X1_LOC_84/A 0.01fF
C6691 NAND2X1_LOC_644/a_36_24# INVX1_LOC_12/A 0.01fF
C6692 NOR2X1_LOC_457/A NOR2X1_LOC_794/B 0.05fF
C6693 NOR2X1_LOC_617/Y INVX1_LOC_5/A 0.02fF
C6694 INVX1_LOC_35/A NOR2X1_LOC_804/B 0.07fF
C6695 INVX1_LOC_91/A INVX1_LOC_179/A 0.03fF
C6696 INVX1_LOC_1/A INVX1_LOC_30/A 0.31fF
C6697 INVX1_LOC_192/A INVX1_LOC_53/A 0.11fF
C6698 INVX1_LOC_124/Y NOR2X1_LOC_361/B 1.17fF
C6699 NAND2X1_LOC_84/Y NOR2X1_LOC_81/Y 0.10fF
C6700 INVX1_LOC_150/Y NAND2X1_LOC_352/B 0.04fF
C6701 NAND2X1_LOC_493/Y INVX1_LOC_72/A 1.73fF
C6702 INVX1_LOC_256/A NOR2X1_LOC_389/A 0.25fF
C6703 NAND2X1_LOC_562/B NOR2X1_LOC_629/A 0.03fF
C6704 INVX1_LOC_39/A INVX1_LOC_24/A 0.05fF
C6705 NOR2X1_LOC_736/Y INVX1_LOC_12/A 0.05fF
C6706 INVX1_LOC_58/A NOR2X1_LOC_300/Y 0.05fF
C6707 VDD NAND2X1_LOC_848/A 0.98fF
C6708 INVX1_LOC_243/Y NAND2X1_LOC_451/Y 0.06fF
C6709 NAND2X1_LOC_763/B INVX1_LOC_1/A 0.22fF
C6710 NOR2X1_LOC_613/a_36_216# NOR2X1_LOC_238/Y 0.00fF
C6711 INVX1_LOC_37/A NOR2X1_LOC_684/Y 0.60fF
C6712 INVX1_LOC_178/A INVX1_LOC_41/Y 0.03fF
C6713 INVX1_LOC_230/Y NOR2X1_LOC_160/B 0.07fF
C6714 INVX1_LOC_316/Y INVX1_LOC_26/A 0.09fF
C6715 INVX1_LOC_244/Y NOR2X1_LOC_763/A 0.02fF
C6716 NOR2X1_LOC_91/A INVX1_LOC_297/Y 0.01fF
C6717 NOR2X1_LOC_280/Y INVX1_LOC_118/A 0.05fF
C6718 D_INPUT_1 INVX1_LOC_54/Y 0.17fF
C6719 NOR2X1_LOC_617/Y INVX1_LOC_178/A 0.05fF
C6720 INVX1_LOC_182/Y NOR2X1_LOC_89/A 0.03fF
C6721 INVX1_LOC_35/A NOR2X1_LOC_309/Y 0.10fF
C6722 NOR2X1_LOC_802/A INVX1_LOC_53/A 0.05fF
C6723 NAND2X1_LOC_35/Y INVX1_LOC_8/A 0.07fF
C6724 INVX1_LOC_178/A NAND2X1_LOC_593/Y 0.05fF
C6725 NOR2X1_LOC_598/B NOR2X1_LOC_156/B 0.03fF
C6726 NOR2X1_LOC_74/A NAND2X1_LOC_81/B 0.07fF
C6727 NOR2X1_LOC_596/A NOR2X1_LOC_348/Y 0.72fF
C6728 NAND2X1_LOC_725/A NAND2X1_LOC_308/Y 0.03fF
C6729 NAND2X1_LOC_624/B NAND2X1_LOC_562/B 0.07fF
C6730 INVX1_LOC_291/A INVX1_LOC_20/A 0.07fF
C6731 NAND2X1_LOC_9/Y NOR2X1_LOC_720/a_36_216# 0.01fF
C6732 INVX1_LOC_85/Y INVX1_LOC_15/A 0.03fF
C6733 NOR2X1_LOC_460/B NOR2X1_LOC_460/Y 0.01fF
C6734 NOR2X1_LOC_186/Y NOR2X1_LOC_772/Y 0.01fF
C6735 NAND2X1_LOC_468/a_36_24# NOR2X1_LOC_435/A 0.00fF
C6736 INVX1_LOC_53/Y NOR2X1_LOC_72/Y 0.05fF
C6737 INVX1_LOC_123/A NOR2X1_LOC_721/B 0.03fF
C6738 INVX1_LOC_21/A NOR2X1_LOC_520/B 0.03fF
C6739 NAND2X1_LOC_366/A NOR2X1_LOC_852/Y 0.61fF
C6740 INVX1_LOC_282/A INVX1_LOC_42/A 0.13fF
C6741 NOR2X1_LOC_321/Y NOR2X1_LOC_577/Y 0.08fF
C6742 NOR2X1_LOC_337/A INVX1_LOC_99/A 0.02fF
C6743 NOR2X1_LOC_188/Y INVX1_LOC_28/Y 0.05fF
C6744 NAND2X1_LOC_724/Y INVX1_LOC_22/A 0.05fF
C6745 NOR2X1_LOC_186/Y NOR2X1_LOC_392/B 0.03fF
C6746 INVX1_LOC_11/Y INVX1_LOC_250/Y 0.23fF
C6747 INVX1_LOC_89/A NAND2X1_LOC_447/a_36_24# 0.00fF
C6748 NAND2X1_LOC_798/B NAND2X1_LOC_453/A 0.17fF
C6749 VDD INVX1_LOC_46/Y 1.61fF
C6750 INVX1_LOC_281/A INVX1_LOC_54/A 0.07fF
C6751 INVX1_LOC_173/Y NOR2X1_LOC_409/B 0.03fF
C6752 NOR2X1_LOC_553/B NOR2X1_LOC_383/B 0.02fF
C6753 NOR2X1_LOC_356/A INVX1_LOC_4/Y 0.01fF
C6754 NAND2X1_LOC_303/Y INVX1_LOC_209/Y 0.03fF
C6755 NOR2X1_LOC_470/B INVX1_LOC_49/A 0.01fF
C6756 INVX1_LOC_122/A NOR2X1_LOC_259/A 0.12fF
C6757 NAND2X1_LOC_687/A INVX1_LOC_92/A 0.03fF
C6758 INVX1_LOC_5/A NOR2X1_LOC_538/Y 0.04fF
C6759 NAND2X1_LOC_773/Y NOR2X1_LOC_593/Y 0.03fF
C6760 INVX1_LOC_256/A NOR2X1_LOC_596/A 1.35fF
C6761 NOR2X1_LOC_218/A INVX1_LOC_71/A 0.01fF
C6762 NOR2X1_LOC_845/A INVX1_LOC_29/A 0.01fF
C6763 NOR2X1_LOC_363/Y INVX1_LOC_92/A 0.08fF
C6764 NAND2X1_LOC_655/A INVX1_LOC_264/A 0.00fF
C6765 INVX1_LOC_89/A INVX1_LOC_23/Y 0.07fF
C6766 NOR2X1_LOC_644/B NOR2X1_LOC_457/B 0.02fF
C6767 INVX1_LOC_54/Y NOR2X1_LOC_652/Y 0.10fF
C6768 INVX1_LOC_30/A NOR2X1_LOC_384/Y 0.05fF
C6769 INVX1_LOC_89/A NOR2X1_LOC_342/B 0.02fF
C6770 INVX1_LOC_7/A NOR2X1_LOC_414/Y 0.11fF
C6771 INVX1_LOC_21/A INVX1_LOC_133/Y 0.00fF
C6772 INVX1_LOC_64/A NAND2X1_LOC_859/B 0.00fF
C6773 D_INPUT_4 NAND2X1_LOC_452/Y 0.03fF
C6774 NOR2X1_LOC_816/A NAND2X1_LOC_593/Y 0.09fF
C6775 INVX1_LOC_21/A INVX1_LOC_276/A 0.38fF
C6776 INVX1_LOC_28/A NOR2X1_LOC_278/Y 0.01fF
C6777 INVX1_LOC_223/A INVX1_LOC_177/Y 0.01fF
C6778 VDD INVX1_LOC_5/Y 0.41fF
C6779 INVX1_LOC_30/A NOR2X1_LOC_522/a_36_216# 0.00fF
C6780 INVX1_LOC_21/A NOR2X1_LOC_67/A 0.30fF
C6781 D_INPUT_3 NAND2X1_LOC_206/Y 0.31fF
C6782 D_INPUT_1 NAND2X1_LOC_125/a_36_24# 0.00fF
C6783 NAND2X1_LOC_850/A INVX1_LOC_26/A 0.77fF
C6784 NOR2X1_LOC_74/A INVX1_LOC_4/Y 0.20fF
C6785 NOR2X1_LOC_590/A INVX1_LOC_77/A 0.23fF
C6786 INVX1_LOC_298/A INVX1_LOC_22/A 0.02fF
C6787 INVX1_LOC_282/A INVX1_LOC_78/A 0.06fF
C6788 NOR2X1_LOC_45/B NOR2X1_LOC_48/B 0.05fF
C6789 NAND2X1_LOC_564/a_36_24# NOR2X1_LOC_103/Y -0.00fF
C6790 NAND2X1_LOC_346/a_36_24# NOR2X1_LOC_612/B 0.00fF
C6791 INVX1_LOC_41/A NOR2X1_LOC_443/a_36_216# 0.00fF
C6792 INVX1_LOC_22/Y INVX1_LOC_77/A 0.03fF
C6793 INVX1_LOC_245/Y INVX1_LOC_153/Y 0.04fF
C6794 NOR2X1_LOC_758/Y NAND2X1_LOC_337/B 0.04fF
C6795 INVX1_LOC_219/A NOR2X1_LOC_392/Y 0.02fF
C6796 INVX1_LOC_14/A NOR2X1_LOC_709/A 0.28fF
C6797 NOR2X1_LOC_329/B NOR2X1_LOC_65/Y 0.04fF
C6798 NOR2X1_LOC_272/Y INVX1_LOC_226/Y 0.03fF
C6799 NOR2X1_LOC_9/Y INVX1_LOC_4/Y 0.10fF
C6800 INVX1_LOC_235/Y INVX1_LOC_197/Y 0.06fF
C6801 INVX1_LOC_39/A NAND2X1_LOC_565/B 0.17fF
C6802 NOR2X1_LOC_82/A NOR2X1_LOC_315/Y 1.16fF
C6803 NOR2X1_LOC_220/a_36_216# NOR2X1_LOC_360/Y 0.01fF
C6804 D_INPUT_6 INVX1_LOC_22/A 0.03fF
C6805 NOR2X1_LOC_778/A NOR2X1_LOC_500/A 0.01fF
C6806 NOR2X1_LOC_130/a_36_216# NOR2X1_LOC_392/Y 0.01fF
C6807 NOR2X1_LOC_831/B NOR2X1_LOC_612/Y 0.01fF
C6808 NAND2X1_LOC_563/Y INPUT_3 0.00fF
C6809 NOR2X1_LOC_567/B INVX1_LOC_57/A 0.07fF
C6810 INVX1_LOC_230/A NAND2X1_LOC_206/Y 0.06fF
C6811 NAND2X1_LOC_53/Y NOR2X1_LOC_627/Y 0.03fF
C6812 NOR2X1_LOC_321/Y INVX1_LOC_22/A 0.07fF
C6813 NOR2X1_LOC_174/A INVX1_LOC_53/A 0.20fF
C6814 NAND2X1_LOC_736/Y NAND2X1_LOC_733/A 0.17fF
C6815 INVX1_LOC_172/A INVX1_LOC_18/A 0.07fF
C6816 NOR2X1_LOC_658/Y INVX1_LOC_34/A 0.08fF
C6817 NOR2X1_LOC_210/A NAND2X1_LOC_149/Y 0.04fF
C6818 INVX1_LOC_208/A NOR2X1_LOC_359/a_36_216# 0.00fF
C6819 INVX1_LOC_254/Y NOR2X1_LOC_68/A 0.09fF
C6820 NOR2X1_LOC_364/a_36_216# INVX1_LOC_109/Y 0.00fF
C6821 INVX1_LOC_9/A NOR2X1_LOC_814/A 0.12fF
C6822 NOR2X1_LOC_272/Y INVX1_LOC_10/A 0.05fF
C6823 INVX1_LOC_124/A NOR2X1_LOC_590/A 0.10fF
C6824 INVX1_LOC_2/A NOR2X1_LOC_369/Y 0.06fF
C6825 INVX1_LOC_159/A INVX1_LOC_49/A 0.07fF
C6826 NAND2X1_LOC_338/B NAND2X1_LOC_529/a_36_24# 0.00fF
C6827 NOR2X1_LOC_78/A NAND2X1_LOC_223/A 0.02fF
C6828 INPUT_6 INVX1_LOC_140/A 0.02fF
C6829 INVX1_LOC_256/A NOR2X1_LOC_220/A 0.10fF
C6830 INVX1_LOC_39/A NOR2X1_LOC_130/A 0.03fF
C6831 NOR2X1_LOC_607/A NOR2X1_LOC_577/Y 0.01fF
C6832 NOR2X1_LOC_226/A NOR2X1_LOC_369/Y 0.02fF
C6833 INVX1_LOC_223/A INVX1_LOC_104/A 0.03fF
C6834 NAND2X1_LOC_391/Y NOR2X1_LOC_71/Y 0.07fF
C6835 NOR2X1_LOC_191/B INVX1_LOC_49/A 0.13fF
C6836 NOR2X1_LOC_440/Y NOR2X1_LOC_468/Y 0.18fF
C6837 INVX1_LOC_58/A NOR2X1_LOC_527/Y 0.01fF
C6838 INVX1_LOC_2/A INVX1_LOC_286/Y 0.17fF
C6839 NOR2X1_LOC_815/Y INVX1_LOC_24/A 0.22fF
C6840 NOR2X1_LOC_186/Y INVX1_LOC_90/A 1.08fF
C6841 INVX1_LOC_284/Y NAND2X1_LOC_717/Y 2.33fF
C6842 NOR2X1_LOC_89/A NOR2X1_LOC_98/B 0.01fF
C6843 INVX1_LOC_64/A NAND2X1_LOC_661/A 0.03fF
C6844 NOR2X1_LOC_234/Y NAND2X1_LOC_634/Y 0.05fF
C6845 NAND2X1_LOC_725/A NAND2X1_LOC_560/A 0.01fF
C6846 NOR2X1_LOC_601/Y INVX1_LOC_271/Y 0.03fF
C6847 NOR2X1_LOC_45/B NOR2X1_LOC_438/Y 0.01fF
C6848 INVX1_LOC_91/A NOR2X1_LOC_693/Y 0.07fF
C6849 NOR2X1_LOC_186/Y NOR2X1_LOC_389/B 0.01fF
C6850 NOR2X1_LOC_226/A INVX1_LOC_286/Y 0.10fF
C6851 NAND2X1_LOC_470/B NAND2X1_LOC_469/B 0.04fF
C6852 INVX1_LOC_66/Y NOR2X1_LOC_114/Y 0.18fF
C6853 INVX1_LOC_49/A INVX1_LOC_283/Y 0.02fF
C6854 NOR2X1_LOC_334/A INVX1_LOC_23/A 6.27fF
C6855 NAND2X1_LOC_363/B NOR2X1_LOC_188/A 0.91fF
C6856 NAND2X1_LOC_86/Y NOR2X1_LOC_843/B 0.01fF
C6857 INVX1_LOC_11/A INVX1_LOC_279/A 0.07fF
C6858 D_INPUT_2 NOR2X1_LOC_84/A 0.07fF
C6859 NAND2X1_LOC_573/Y INVX1_LOC_90/A 0.07fF
C6860 INVX1_LOC_57/Y NAND2X1_LOC_374/Y 0.08fF
C6861 INVX1_LOC_186/A NOR2X1_LOC_748/A 0.01fF
C6862 NOR2X1_LOC_361/B D_INPUT_0 0.00fF
C6863 NOR2X1_LOC_667/A NAND2X1_LOC_726/a_36_24# 0.00fF
C6864 NAND2X1_LOC_363/B NOR2X1_LOC_548/B 0.03fF
C6865 NOR2X1_LOC_790/A NOR2X1_LOC_356/A 0.03fF
C6866 NAND2X1_LOC_803/B NAND2X1_LOC_796/Y 0.03fF
C6867 NOR2X1_LOC_617/Y NAND2X1_LOC_562/B 0.02fF
C6868 INVX1_LOC_2/A INVX1_LOC_159/A 0.01fF
C6869 NOR2X1_LOC_423/a_36_216# INVX1_LOC_6/A 0.01fF
C6870 NAND2X1_LOC_725/B INVX1_LOC_207/Y 0.01fF
C6871 NAND2X1_LOC_588/B INVX1_LOC_243/A 0.30fF
C6872 NOR2X1_LOC_78/B NOR2X1_LOC_791/B 0.10fF
C6873 NOR2X1_LOC_681/Y INVX1_LOC_273/A 0.53fF
C6874 INVX1_LOC_17/A INVX1_LOC_120/A 0.02fF
C6875 INVX1_LOC_37/A INVX1_LOC_273/A 0.03fF
C6876 NAND2X1_LOC_84/Y NOR2X1_LOC_709/A 0.16fF
C6877 NOR2X1_LOC_248/Y INVX1_LOC_53/Y 0.01fF
C6878 NOR2X1_LOC_226/A INVX1_LOC_159/A 0.02fF
C6879 NOR2X1_LOC_155/A INVX1_LOC_29/A 0.01fF
C6880 NAND2X1_LOC_785/Y NOR2X1_LOC_753/Y 0.00fF
C6881 NAND2X1_LOC_63/Y NOR2X1_LOC_197/B 0.00fF
C6882 INVX1_LOC_36/A NOR2X1_LOC_121/A 0.03fF
C6883 NOR2X1_LOC_481/A NOR2X1_LOC_392/B 0.23fF
C6884 NAND2X1_LOC_796/B NOR2X1_LOC_323/Y 0.00fF
C6885 NAND2X1_LOC_579/A NOR2X1_LOC_490/Y 0.03fF
C6886 NOR2X1_LOC_590/A NAND2X1_LOC_796/Y 0.01fF
C6887 NAND2X1_LOC_231/Y NOR2X1_LOC_13/Y 0.12fF
C6888 INVX1_LOC_225/A NOR2X1_LOC_772/Y 0.01fF
C6889 NAND2X1_LOC_16/Y INVX1_LOC_22/A 0.20fF
C6890 NOR2X1_LOC_92/Y NOR2X1_LOC_289/Y 0.01fF
C6891 INVX1_LOC_225/A NOR2X1_LOC_392/B 0.10fF
C6892 NAND2X1_LOC_565/B INVX1_LOC_61/A 0.01fF
C6893 NOR2X1_LOC_667/A NOR2X1_LOC_753/Y 0.07fF
C6894 INVX1_LOC_254/A INVX1_LOC_218/A 0.03fF
C6895 NAND2X1_LOC_361/Y NOR2X1_LOC_537/Y 0.07fF
C6896 NOR2X1_LOC_160/B INVX1_LOC_196/Y 0.03fF
C6897 NAND2X1_LOC_347/B NOR2X1_LOC_83/a_36_216# 0.03fF
C6898 NAND2X1_LOC_93/B INVX1_LOC_251/A 0.01fF
C6899 NAND2X1_LOC_656/A INVX1_LOC_1/Y 0.01fF
C6900 NOR2X1_LOC_209/Y NOR2X1_LOC_147/B 0.02fF
C6901 NAND2X1_LOC_181/Y NOR2X1_LOC_716/B 0.20fF
C6902 NAND2X1_LOC_364/A INVX1_LOC_10/A 0.03fF
C6903 INVX1_LOC_24/A NAND2X1_LOC_735/B 0.00fF
C6904 INVX1_LOC_286/Y NAND2X1_LOC_648/A 0.05fF
C6905 NAND2X1_LOC_361/Y NAND2X1_LOC_323/B 0.07fF
C6906 NOR2X1_LOC_667/A NAND2X1_LOC_325/Y 0.01fF
C6907 NOR2X1_LOC_624/A INVX1_LOC_143/A 0.03fF
C6908 NOR2X1_LOC_205/Y NOR2X1_LOC_74/A 0.04fF
C6909 INVX1_LOC_248/A NAND2X1_LOC_325/Y 0.07fF
C6910 INVX1_LOC_19/A NAND2X1_LOC_82/Y 0.78fF
C6911 INVX1_LOC_24/A NOR2X1_LOC_302/a_36_216# 0.02fF
C6912 NOR2X1_LOC_458/B NOR2X1_LOC_570/B 0.65fF
C6913 INVX1_LOC_236/Y INVX1_LOC_28/A 0.01fF
C6914 NAND2X1_LOC_711/B NOR2X1_LOC_690/Y 0.22fF
C6915 INVX1_LOC_24/A INPUT_5 0.05fF
C6916 NOR2X1_LOC_612/B NOR2X1_LOC_709/A 0.13fF
C6917 INVX1_LOC_271/Y NOR2X1_LOC_676/a_36_216# 0.00fF
C6918 INVX1_LOC_119/A NOR2X1_LOC_511/a_36_216# 0.12fF
C6919 INVX1_LOC_61/A NOR2X1_LOC_130/A 0.07fF
C6920 INVX1_LOC_11/A NAND2X1_LOC_858/B 0.01fF
C6921 NOR2X1_LOC_861/Y NOR2X1_LOC_814/A 0.07fF
C6922 INVX1_LOC_76/A NOR2X1_LOC_665/Y 0.03fF
C6923 NOR2X1_LOC_457/A NOR2X1_LOC_188/A 0.22fF
C6924 INVX1_LOC_8/A INVX1_LOC_56/A 0.02fF
C6925 NAND2X1_LOC_112/Y INVX1_LOC_33/A 0.04fF
C6926 INVX1_LOC_227/A INVX1_LOC_77/A 0.07fF
C6927 INVX1_LOC_279/A NOR2X1_LOC_433/A 0.04fF
C6928 INVX1_LOC_269/A NOR2X1_LOC_355/B 0.08fF
C6929 INVX1_LOC_19/A NOR2X1_LOC_461/Y 0.04fF
C6930 INVX1_LOC_251/A INVX1_LOC_3/A 0.04fF
C6931 INVX1_LOC_72/A NAND2X1_LOC_654/B 0.07fF
C6932 INVX1_LOC_276/A INVX1_LOC_214/A 0.06fF
C6933 NOR2X1_LOC_763/Y INVX1_LOC_77/A 0.13fF
C6934 NAND2X1_LOC_487/a_36_24# INVX1_LOC_26/A 0.00fF
C6935 INVX1_LOC_279/A NOR2X1_LOC_593/Y 0.07fF
C6936 NOR2X1_LOC_619/A NOR2X1_LOC_6/B 0.44fF
C6937 INVX1_LOC_298/Y NOR2X1_LOC_155/A 0.03fF
C6938 NOR2X1_LOC_68/A INVX1_LOC_311/Y 0.03fF
C6939 NOR2X1_LOC_815/Y NAND2X1_LOC_783/A 0.09fF
C6940 INVX1_LOC_209/A NOR2X1_LOC_505/Y 0.07fF
C6941 NAND2X1_LOC_122/a_36_24# NOR2X1_LOC_719/A 0.00fF
C6942 INVX1_LOC_47/A INVX1_LOC_314/Y 0.02fF
C6943 INVX1_LOC_104/A NOR2X1_LOC_730/Y 0.05fF
C6944 NAND2X1_LOC_731/Y INVX1_LOC_28/A 0.07fF
C6945 INVX1_LOC_35/A NOR2X1_LOC_865/A 0.37fF
C6946 INVX1_LOC_135/A NOR2X1_LOC_551/B 0.03fF
C6947 NOR2X1_LOC_15/Y NOR2X1_LOC_631/B 0.06fF
C6948 INVX1_LOC_30/A NOR2X1_LOC_188/A 0.89fF
C6949 NAND2X1_LOC_775/a_36_24# NAND2X1_LOC_564/B 0.00fF
C6950 INVX1_LOC_190/Y INVX1_LOC_49/A 0.05fF
C6951 NAND2X1_LOC_454/Y INVX1_LOC_84/A 0.07fF
C6952 INVX1_LOC_132/A INVX1_LOC_90/A 0.42fF
C6953 NAND2X1_LOC_350/A NOR2X1_LOC_45/B 0.14fF
C6954 INVX1_LOC_83/A INVX1_LOC_192/A 0.06fF
C6955 INVX1_LOC_279/A NOR2X1_LOC_52/B 0.03fF
C6956 INVX1_LOC_30/A NOR2X1_LOC_548/B 0.03fF
C6957 NOR2X1_LOC_646/A NOR2X1_LOC_78/B 0.03fF
C6958 INVX1_LOC_41/Y INVX1_LOC_140/A 0.04fF
C6959 INVX1_LOC_255/Y NAND2X1_LOC_578/B 0.03fF
C6960 NOR2X1_LOC_518/Y INPUT_0 0.14fF
C6961 INVX1_LOC_41/A INVX1_LOC_65/Y 0.02fF
C6962 INVX1_LOC_29/Y INVX1_LOC_92/A 0.02fF
C6963 NOR2X1_LOC_448/Y VDD 0.14fF
C6964 INVX1_LOC_77/A NOR2X1_LOC_703/A 0.03fF
C6965 NOR2X1_LOC_2/Y NOR2X1_LOC_3/a_36_216# 0.00fF
C6966 INVX1_LOC_223/A INVX1_LOC_206/Y 0.00fF
C6967 NOR2X1_LOC_598/B INVX1_LOC_152/A 0.12fF
C6968 INVX1_LOC_140/A NAND2X1_LOC_593/Y 0.04fF
C6969 INVX1_LOC_278/A NOR2X1_LOC_487/Y 0.03fF
C6970 NOR2X1_LOC_67/A NOR2X1_LOC_521/Y 0.01fF
C6971 NOR2X1_LOC_441/Y NOR2X1_LOC_45/B 0.03fF
C6972 INVX1_LOC_83/A NOR2X1_LOC_802/A 0.07fF
C6973 NOR2X1_LOC_15/Y INVX1_LOC_37/A 0.08fF
C6974 NOR2X1_LOC_186/Y INVX1_LOC_38/A 0.05fF
C6975 INVX1_LOC_89/A NAND2X1_LOC_116/A 0.03fF
C6976 NOR2X1_LOC_433/A INVX1_LOC_182/Y 0.04fF
C6977 INVX1_LOC_229/A VDD 0.26fF
C6978 INVX1_LOC_225/A INVX1_LOC_90/A 0.10fF
C6979 INVX1_LOC_256/A NAND2X1_LOC_469/B 0.21fF
C6980 NOR2X1_LOC_598/B NOR2X1_LOC_634/A 0.12fF
C6981 NOR2X1_LOC_361/B NOR2X1_LOC_266/B 0.05fF
C6982 NAND2X1_LOC_15/a_36_24# INVX1_LOC_37/A 0.00fF
C6983 D_INPUT_0 INVX1_LOC_177/A 0.24fF
C6984 INVX1_LOC_35/A NOR2X1_LOC_435/A 0.03fF
C6985 INVX1_LOC_64/A INVX1_LOC_291/A 0.00fF
C6986 INVX1_LOC_203/A NOR2X1_LOC_693/Y 0.00fF
C6987 INVX1_LOC_225/A NOR2X1_LOC_389/B 1.21fF
C6988 INVX1_LOC_182/Y NOR2X1_LOC_593/Y 0.03fF
C6989 INVX1_LOC_50/A INVX1_LOC_119/Y 0.20fF
C6990 NAND2X1_LOC_552/A INVX1_LOC_185/A 0.02fF
C6991 NAND2X1_LOC_717/Y NOR2X1_LOC_525/Y 0.33fF
C6992 NOR2X1_LOC_273/Y INVX1_LOC_6/A 0.03fF
C6993 INVX1_LOC_174/A NAND2X1_LOC_1/Y 0.69fF
C6994 INVX1_LOC_30/A NOR2X1_LOC_43/Y 0.23fF
C6995 NAND2X1_LOC_508/A NAND2X1_LOC_116/A 0.03fF
C6996 NAND2X1_LOC_30/Y VDD 0.59fF
C6997 NOR2X1_LOC_759/Y INVX1_LOC_6/A 0.14fF
C6998 NOR2X1_LOC_207/A D_GATE_366 0.06fF
C6999 INVX1_LOC_202/A INVX1_LOC_6/A 0.10fF
C7000 INVX1_LOC_90/A NOR2X1_LOC_209/Y 0.41fF
C7001 INVX1_LOC_174/A NOR2X1_LOC_145/Y 0.02fF
C7002 NOR2X1_LOC_297/a_36_216# NAND2X1_LOC_348/A 0.00fF
C7003 NOR2X1_LOC_91/A NAND2X1_LOC_74/B 0.06fF
C7004 NAND2X1_LOC_724/A INVX1_LOC_38/A 0.07fF
C7005 INVX1_LOC_178/A INVX1_LOC_185/A 0.05fF
C7006 NOR2X1_LOC_134/Y VDD 0.63fF
C7007 NOR2X1_LOC_668/Y NAND2X1_LOC_74/B 0.03fF
C7008 NAND2X1_LOC_46/a_36_24# NOR2X1_LOC_673/A 0.00fF
C7009 INVX1_LOC_45/Y INVX1_LOC_91/A 0.01fF
C7010 NOR2X1_LOC_244/B INVX1_LOC_89/A 0.02fF
C7011 NOR2X1_LOC_75/Y INVX1_LOC_117/A 0.07fF
C7012 INVX1_LOC_24/Y NAND2X1_LOC_617/a_36_24# 0.06fF
C7013 NOR2X1_LOC_243/Y NAND2X1_LOC_348/A 0.04fF
C7014 INVX1_LOC_89/A INVX1_LOC_232/A 0.16fF
C7015 NOR2X1_LOC_391/A NOR2X1_LOC_719/B 0.21fF
C7016 NOR2X1_LOC_78/B NOR2X1_LOC_111/Y 0.02fF
C7017 NAND2X1_LOC_454/Y INVX1_LOC_15/A 0.18fF
C7018 NOR2X1_LOC_68/A NOR2X1_LOC_683/a_36_216# 0.00fF
C7019 INVX1_LOC_35/A INVX1_LOC_63/A 0.13fF
C7020 NAND2X1_LOC_198/B NOR2X1_LOC_124/A 0.00fF
C7021 NAND2X1_LOC_656/A INVX1_LOC_93/Y 0.10fF
C7022 NOR2X1_LOC_843/A NOR2X1_LOC_9/Y 0.04fF
C7023 INVX1_LOC_11/A NOR2X1_LOC_450/A 0.08fF
C7024 NAND2X1_LOC_120/a_36_24# NAND2X1_LOC_472/Y 0.00fF
C7025 NOR2X1_LOC_13/Y NAND2X1_LOC_649/B 0.19fF
C7026 INVX1_LOC_278/Y NOR2X1_LOC_166/Y 0.13fF
C7027 NOR2X1_LOC_295/Y INVX1_LOC_69/Y 0.03fF
C7028 NOR2X1_LOC_769/B INVX1_LOC_29/A 0.02fF
C7029 NOR2X1_LOC_218/A NOR2X1_LOC_331/B 0.03fF
C7030 INVX1_LOC_23/A NAND2X1_LOC_74/B 0.07fF
C7031 INVX1_LOC_249/Y INVX1_LOC_6/A 0.01fF
C7032 D_INPUT_1 NOR2X1_LOC_610/Y 0.01fF
C7033 INVX1_LOC_286/Y NOR2X1_LOC_694/a_36_216# 0.01fF
C7034 NOR2X1_LOC_598/B INVX1_LOC_29/A 0.25fF
C7035 INVX1_LOC_314/Y INVX1_LOC_95/Y 0.57fF
C7036 INVX1_LOC_33/A NOR2X1_LOC_78/A 1.90fF
C7037 NAND2X1_LOC_740/A INVX1_LOC_11/Y 0.01fF
C7038 INVX1_LOC_85/A INVX1_LOC_206/Y 0.03fF
C7039 INVX1_LOC_226/Y NOR2X1_LOC_393/a_36_216# 0.00fF
C7040 INVX1_LOC_129/A INVX1_LOC_42/A 0.01fF
C7041 INVX1_LOC_256/Y INPUT_0 0.07fF
C7042 INVX1_LOC_48/A NOR2X1_LOC_709/A 0.03fF
C7043 INVX1_LOC_49/A NOR2X1_LOC_56/Y 0.07fF
C7044 NOR2X1_LOC_590/A INVX1_LOC_9/A 0.17fF
C7045 INVX1_LOC_1/A INVX1_LOC_113/A 0.18fF
C7046 INVX1_LOC_97/Y INVX1_LOC_29/A 0.01fF
C7047 NOR2X1_LOC_816/A INVX1_LOC_185/A 0.03fF
C7048 INVX1_LOC_11/A NOR2X1_LOC_624/B 0.00fF
C7049 NOR2X1_LOC_160/B NOR2X1_LOC_641/Y 0.00fF
C7050 NAND2X1_LOC_862/A NOR2X1_LOC_74/A 0.02fF
C7051 NAND2X1_LOC_7/Y NOR2X1_LOC_35/Y 0.08fF
C7052 INVX1_LOC_24/A INVX1_LOC_14/Y 0.03fF
C7053 NOR2X1_LOC_401/Y INVX1_LOC_286/A 0.01fF
C7054 NAND2X1_LOC_567/Y INVX1_LOC_76/A 0.01fF
C7055 NOR2X1_LOC_354/B NOR2X1_LOC_319/B -0.01fF
C7056 INVX1_LOC_151/Y INVX1_LOC_144/A 0.04fF
C7057 NOR2X1_LOC_392/B NAND2X1_LOC_642/Y 0.10fF
C7058 NOR2X1_LOC_220/A INVX1_LOC_69/Y 0.10fF
C7059 NOR2X1_LOC_174/A INVX1_LOC_83/A 0.00fF
C7060 NOR2X1_LOC_660/Y NOR2X1_LOC_847/a_36_216# 0.00fF
C7061 NAND2X1_LOC_624/B INVX1_LOC_42/A 0.04fF
C7062 NOR2X1_LOC_714/Y NOR2X1_LOC_78/A 0.01fF
C7063 NOR2X1_LOC_263/a_36_216# INVX1_LOC_93/Y 0.01fF
C7064 INVX1_LOC_49/A VDD 1.51fF
C7065 NAND2X1_LOC_162/B INVX1_LOC_117/A 0.03fF
C7066 INVX1_LOC_236/A NAND2X1_LOC_655/A 0.10fF
C7067 NOR2X1_LOC_420/Y NOR2X1_LOC_89/A 0.06fF
C7068 NOR2X1_LOC_391/Y INVX1_LOC_16/A 0.02fF
C7069 INVX1_LOC_89/A NOR2X1_LOC_775/Y 0.02fF
C7070 NOR2X1_LOC_181/a_36_216# NOR2X1_LOC_155/A 0.00fF
C7071 NOR2X1_LOC_272/Y INVX1_LOC_12/A 0.00fF
C7072 NOR2X1_LOC_419/Y INVX1_LOC_117/A 0.10fF
C7073 NOR2X1_LOC_78/B NOR2X1_LOC_192/A 0.01fF
C7074 NOR2X1_LOC_350/a_36_216# INVX1_LOC_176/A 0.00fF
C7075 NAND2X1_LOC_20/B NOR2X1_LOC_814/A 0.04fF
C7076 INVX1_LOC_69/Y NOR2X1_LOC_548/Y 0.43fF
C7077 INVX1_LOC_2/A NOR2X1_LOC_56/Y 0.03fF
C7078 INVX1_LOC_40/A NOR2X1_LOC_78/A 0.11fF
C7079 NOR2X1_LOC_665/a_36_216# INVX1_LOC_4/A 0.00fF
C7080 INVX1_LOC_26/A INVX1_LOC_57/A 0.17fF
C7081 INVX1_LOC_60/A VDD 0.12fF
C7082 NOR2X1_LOC_336/B NOR2X1_LOC_445/B 0.01fF
C7083 NAND2X1_LOC_555/Y NAND2X1_LOC_659/A -0.02fF
C7084 NOR2X1_LOC_635/A INVX1_LOC_37/A 0.00fF
C7085 NOR2X1_LOC_226/A NOR2X1_LOC_56/Y 0.11fF
C7086 NOR2X1_LOC_423/Y INVX1_LOC_139/A 0.02fF
C7087 NOR2X1_LOC_471/Y NOR2X1_LOC_631/A 0.02fF
C7088 INVX1_LOC_132/A INVX1_LOC_38/A 0.07fF
C7089 NOR2X1_LOC_500/Y NOR2X1_LOC_405/A 0.26fF
C7090 NOR2X1_LOC_554/B NAND2X1_LOC_817/a_36_24# -0.01fF
C7091 NOR2X1_LOC_468/Y NOR2X1_LOC_89/A 0.07fF
C7092 NAND2X1_LOC_84/Y NOR2X1_LOC_489/A 0.01fF
C7093 NOR2X1_LOC_67/A NOR2X1_LOC_670/Y 0.03fF
C7094 NOR2X1_LOC_142/Y INVX1_LOC_281/A 0.01fF
C7095 INVX1_LOC_298/Y NOR2X1_LOC_598/B 0.02fF
C7096 NOR2X1_LOC_717/B NAND2X1_LOC_679/a_36_24# 0.00fF
C7097 INVX1_LOC_2/A NOR2X1_LOC_69/a_36_216# 0.00fF
C7098 NAND2X1_LOC_190/Y NOR2X1_LOC_89/A 0.27fF
C7099 NOR2X1_LOC_65/B INVX1_LOC_129/A 0.19fF
C7100 INVX1_LOC_2/A VDD 4.96fF
C7101 NOR2X1_LOC_818/Y VDD 0.12fF
C7102 NOR2X1_LOC_68/A NOR2X1_LOC_88/Y 0.07fF
C7103 INVX1_LOC_155/Y NOR2X1_LOC_331/B 0.02fF
C7104 NAND2X1_LOC_114/B INVX1_LOC_19/A 0.08fF
C7105 INVX1_LOC_2/A NAND2X1_LOC_800/A 0.03fF
C7106 NOR2X1_LOC_78/B INVX1_LOC_2/Y 0.18fF
C7107 NOR2X1_LOC_226/A INVX1_LOC_146/Y 0.01fF
C7108 NOR2X1_LOC_222/Y INVX1_LOC_139/A 0.03fF
C7109 NOR2X1_LOC_226/A VDD 1.40fF
C7110 INVX1_LOC_58/A NOR2X1_LOC_654/A 0.04fF
C7111 INVX1_LOC_300/Y NAND2X1_LOC_810/B 0.00fF
C7112 NOR2X1_LOC_285/A INVX1_LOC_23/A 0.01fF
C7113 NOR2X1_LOC_392/B NOR2X1_LOC_271/Y 0.01fF
C7114 NAND2X1_LOC_181/Y NAND2X1_LOC_633/Y 0.22fF
C7115 NOR2X1_LOC_113/A INVX1_LOC_10/A 0.01fF
C7116 NOR2X1_LOC_255/Y INVX1_LOC_57/A 0.01fF
C7117 NOR2X1_LOC_431/Y NOR2X1_LOC_592/B 0.01fF
C7118 NOR2X1_LOC_688/Y NOR2X1_LOC_691/B 0.10fF
C7119 NOR2X1_LOC_405/A INVX1_LOC_10/A 0.07fF
C7120 NOR2X1_LOC_598/B INVX1_LOC_204/A 0.02fF
C7121 NOR2X1_LOC_71/Y INVX1_LOC_91/A 0.10fF
C7122 INVX1_LOC_89/A NOR2X1_LOC_685/A 0.00fF
C7123 NOR2X1_LOC_681/Y NAND2X1_LOC_840/B 0.00fF
C7124 NOR2X1_LOC_748/Y NOR2X1_LOC_538/a_36_216# 0.00fF
C7125 NOR2X1_LOC_68/A INVX1_LOC_84/A 0.51fF
C7126 INVX1_LOC_185/Y INVX1_LOC_118/A 0.01fF
C7127 INVX1_LOC_31/A NAND2X1_LOC_74/B 0.35fF
C7128 D_INPUT_1 NAND2X1_LOC_860/A 0.03fF
C7129 NOR2X1_LOC_328/Y NAND2X1_LOC_453/A 0.04fF
C7130 INVX1_LOC_53/A INVX1_LOC_29/Y 2.03fF
C7131 INVX1_LOC_200/Y NAND2X1_LOC_793/B 0.01fF
C7132 INVX1_LOC_31/A NAND2X1_LOC_207/Y 0.04fF
C7133 NAND2X1_LOC_462/B NAND2X1_LOC_659/B 0.21fF
C7134 NOR2X1_LOC_218/Y VDD 0.17fF
C7135 INVX1_LOC_312/Y INVX1_LOC_19/A 0.08fF
C7136 INVX1_LOC_47/A NOR2X1_LOC_557/A 0.00fF
C7137 NOR2X1_LOC_161/Y VDD 0.24fF
C7138 NOR2X1_LOC_389/A NOR2X1_LOC_89/A 0.01fF
C7139 INVX1_LOC_63/Y NAND2X1_LOC_93/B 0.07fF
C7140 INVX1_LOC_61/Y INVX1_LOC_284/A 0.03fF
C7141 NOR2X1_LOC_644/A INVX1_LOC_91/A 0.03fF
C7142 INVX1_LOC_23/A NOR2X1_LOC_660/Y 0.02fF
C7143 INVX1_LOC_157/A NAND2X1_LOC_469/B 0.01fF
C7144 NOR2X1_LOC_589/A NAND2X1_LOC_39/Y 0.14fF
C7145 NAND2X1_LOC_286/B NOR2X1_LOC_652/Y 0.11fF
C7146 INVX1_LOC_31/A NOR2X1_LOC_847/B 0.01fF
C7147 INVX1_LOC_90/A NAND2X1_LOC_642/Y 0.15fF
C7148 INVX1_LOC_14/A NAND2X1_LOC_444/B 0.02fF
C7149 INVX1_LOC_11/A NOR2X1_LOC_38/B 0.06fF
C7150 NAND2X1_LOC_462/B VDD 0.01fF
C7151 NOR2X1_LOC_68/A NAND2X1_LOC_651/B 0.04fF
C7152 NOR2X1_LOC_828/B INVX1_LOC_91/A 0.00fF
C7153 INVX1_LOC_50/A NOR2X1_LOC_674/Y 0.18fF
C7154 INVX1_LOC_89/A NAND2X1_LOC_447/Y 0.01fF
C7155 NOR2X1_LOC_367/B NOR2X1_LOC_364/A 0.01fF
C7156 INVX1_LOC_83/A INVX1_LOC_2/Y 0.02fF
C7157 NAND2X1_LOC_364/A INVX1_LOC_12/A 0.03fF
C7158 NOR2X1_LOC_795/a_36_216# INVX1_LOC_37/A 0.00fF
C7159 NOR2X1_LOC_130/A D_INPUT_3 0.03fF
C7160 NOR2X1_LOC_470/A INVX1_LOC_117/A 0.18fF
C7161 NOR2X1_LOC_78/B INVX1_LOC_307/Y 0.01fF
C7162 NOR2X1_LOC_111/A NAND2X1_LOC_808/A 0.10fF
C7163 NOR2X1_LOC_424/Y INVX1_LOC_117/A 0.18fF
C7164 NOR2X1_LOC_773/Y INVX1_LOC_185/A 0.01fF
C7165 INVX1_LOC_182/A INVX1_LOC_247/A 0.01fF
C7166 VDD NAND2X1_LOC_648/A 0.32fF
C7167 NOR2X1_LOC_717/B INVX1_LOC_117/A 0.03fF
C7168 NAND2X1_LOC_562/a_36_24# INVX1_LOC_15/A 0.00fF
C7169 NOR2X1_LOC_68/A NAND2X1_LOC_220/B 0.18fF
C7170 INVX1_LOC_49/A INVX1_LOC_133/A 0.03fF
C7171 NOR2X1_LOC_596/A NOR2X1_LOC_89/A 0.07fF
C7172 NOR2X1_LOC_92/Y INVX1_LOC_296/Y 0.05fF
C7173 VDD INPUT_1 0.99fF
C7174 D_INPUT_1 NAND2X1_LOC_473/A 0.04fF
C7175 NOR2X1_LOC_78/B NOR2X1_LOC_608/Y -0.01fF
C7176 NAND2X1_LOC_800/A NAND2X1_LOC_648/A 0.00fF
C7177 INVX1_LOC_77/A NOR2X1_LOC_77/a_36_216# 0.01fF
C7178 NAND2X1_LOC_845/a_36_24# INVX1_LOC_284/A 0.01fF
C7179 INVX1_LOC_215/A NAND2X1_LOC_760/a_36_24# -0.02fF
C7180 INVX1_LOC_41/Y INVX1_LOC_42/A 0.03fF
C7181 NOR2X1_LOC_82/A NAND2X1_LOC_99/A 0.18fF
C7182 NOR2X1_LOC_473/B INVX1_LOC_12/Y 0.36fF
C7183 INVX1_LOC_22/A NOR2X1_LOC_433/Y 0.01fF
C7184 NOR2X1_LOC_111/Y INVX1_LOC_46/A 0.02fF
C7185 INVX1_LOC_227/A INVX1_LOC_9/A 1.08fF
C7186 NAND2X1_LOC_513/B NOR2X1_LOC_678/A 0.01fF
C7187 NOR2X1_LOC_208/Y NOR2X1_LOC_631/a_36_216# 0.00fF
C7188 NOR2X1_LOC_68/A INVX1_LOC_15/A 6.96fF
C7189 INVX1_LOC_21/A INVX1_LOC_68/A 0.05fF
C7190 NAND2X1_LOC_114/B INVX1_LOC_26/Y 0.07fF
C7191 NAND2X1_LOC_319/A NOR2X1_LOC_506/Y 0.16fF
C7192 INVX1_LOC_22/A NAND2X1_LOC_798/B 0.07fF
C7193 NAND2X1_LOC_593/Y INVX1_LOC_42/A 0.01fF
C7194 NAND2X1_LOC_805/a_36_24# NAND2X1_LOC_286/B 0.00fF
C7195 NOR2X1_LOC_107/Y INVX1_LOC_57/A 0.07fF
C7196 INVX1_LOC_171/A NOR2X1_LOC_186/a_36_216# 0.00fF
C7197 NAND2X1_LOC_337/B INVX1_LOC_270/Y 0.27fF
C7198 INVX1_LOC_227/Y NOR2X1_LOC_334/Y 0.02fF
C7199 INVX1_LOC_41/A INVX1_LOC_102/A 0.16fF
C7200 NOR2X1_LOC_561/Y NOR2X1_LOC_364/A 0.10fF
C7201 INVX1_LOC_279/A NOR2X1_LOC_858/a_36_216# 0.00fF
C7202 INVX1_LOC_28/A NAND2X1_LOC_808/a_36_24# 0.00fF
C7203 NAND2X1_LOC_863/B INVX1_LOC_297/A 0.39fF
C7204 INVX1_LOC_58/A NOR2X1_LOC_75/Y 0.01fF
C7205 NOR2X1_LOC_307/A INVX1_LOC_23/A 0.03fF
C7206 NOR2X1_LOC_168/B INVX1_LOC_19/A 0.23fF
C7207 INVX1_LOC_13/A NAND2X1_LOC_141/Y 0.08fF
C7208 NOR2X1_LOC_151/Y INVX1_LOC_117/A 0.07fF
C7209 NOR2X1_LOC_355/A INVX1_LOC_92/A 0.03fF
C7210 NOR2X1_LOC_276/Y INVX1_LOC_23/A 0.04fF
C7211 INVX1_LOC_265/A NOR2X1_LOC_48/B 0.09fF
C7212 NAND2X1_LOC_43/a_36_24# INVX1_LOC_108/Y 0.01fF
C7213 NOR2X1_LOC_647/Y NOR2X1_LOC_647/A 0.11fF
C7214 NAND2X1_LOC_33/Y NAND2X1_LOC_410/a_36_24# 0.00fF
C7215 NOR2X1_LOC_706/Y VDD 0.24fF
C7216 NOR2X1_LOC_99/B NOR2X1_LOC_862/B 0.10fF
C7217 NAND2X1_LOC_656/A INVX1_LOC_87/A 0.02fF
C7218 INVX1_LOC_41/Y INVX1_LOC_78/A 0.03fF
C7219 NAND2X1_LOC_477/A INVX1_LOC_102/A 0.10fF
C7220 INVX1_LOC_104/A INVX1_LOC_290/Y 0.01fF
C7221 NOR2X1_LOC_91/A INVX1_LOC_136/A 0.16fF
C7222 NAND2X1_LOC_140/A NOR2X1_LOC_155/A 0.00fF
C7223 INVX1_LOC_255/Y INVX1_LOC_203/A 0.10fF
C7224 INVX1_LOC_45/A NOR2X1_LOC_858/A 0.01fF
C7225 INVX1_LOC_50/A INVX1_LOC_72/A 0.18fF
C7226 NAND2X1_LOC_593/Y INVX1_LOC_78/A 0.02fF
C7227 NOR2X1_LOC_561/Y NOR2X1_LOC_814/A 0.01fF
C7228 NOR2X1_LOC_387/Y NOR2X1_LOC_409/B 0.01fF
C7229 NAND2X1_LOC_336/a_36_24# NOR2X1_LOC_109/Y 0.01fF
C7230 INVX1_LOC_89/A NAND2X1_LOC_750/a_36_24# 0.00fF
C7231 INVX1_LOC_140/A INVX1_LOC_185/A 0.05fF
C7232 INVX1_LOC_7/A NOR2X1_LOC_814/A 0.04fF
C7233 INVX1_LOC_31/A NOR2X1_LOC_660/Y 0.18fF
C7234 NOR2X1_LOC_736/Y INVX1_LOC_92/A 0.03fF
C7235 NOR2X1_LOC_71/Y NOR2X1_LOC_179/Y 0.01fF
C7236 INVX1_LOC_154/A VDD 0.12fF
C7237 NOR2X1_LOC_456/Y INVX1_LOC_36/A 0.01fF
C7238 INVX1_LOC_136/A INVX1_LOC_23/A 0.15fF
C7239 INVX1_LOC_63/Y NAND2X1_LOC_470/B 0.03fF
C7240 NOR2X1_LOC_666/Y NOR2X1_LOC_666/A 0.03fF
C7241 NOR2X1_LOC_799/B NOR2X1_LOC_857/A 0.01fF
C7242 NOR2X1_LOC_261/Y NOR2X1_LOC_68/A 0.20fF
C7243 NOR2X1_LOC_71/Y INVX1_LOC_203/A 0.03fF
C7244 NAND2X1_LOC_108/a_36_24# INVX1_LOC_37/A 0.00fF
C7245 NAND2X1_LOC_9/Y NOR2X1_LOC_791/B 1.40fF
C7246 INVX1_LOC_139/A NOR2X1_LOC_69/A 0.04fF
C7247 INVX1_LOC_263/A INVX1_LOC_290/Y 0.02fF
C7248 NOR2X1_LOC_181/Y INVX1_LOC_271/Y 0.05fF
C7249 NOR2X1_LOC_577/Y NAND2X1_LOC_211/a_36_24# 0.00fF
C7250 NAND2X1_LOC_656/Y INVX1_LOC_19/A 0.01fF
C7251 INPUT_0 NOR2X1_LOC_640/Y 0.07fF
C7252 NAND2X1_LOC_632/a_36_24# INVX1_LOC_12/A 0.01fF
C7253 INVX1_LOC_55/Y NOR2X1_LOC_66/Y 0.04fF
C7254 INVX1_LOC_11/A NOR2X1_LOC_468/Y 0.07fF
C7255 NOR2X1_LOC_562/A INVX1_LOC_76/A 0.03fF
C7256 NAND2X1_LOC_324/a_36_24# NOR2X1_LOC_250/A 0.00fF
C7257 INVX1_LOC_277/A NOR2X1_LOC_840/A 0.03fF
C7258 NOR2X1_LOC_561/A NAND2X1_LOC_642/Y 0.03fF
C7259 INVX1_LOC_11/A NAND2X1_LOC_190/Y 0.05fF
C7260 INVX1_LOC_111/Y NOR2X1_LOC_334/Y 0.02fF
C7261 VDD NOR2X1_LOC_586/Y 0.38fF
C7262 INVX1_LOC_10/A INVX1_LOC_109/Y 0.02fF
C7263 INVX1_LOC_38/A NAND2X1_LOC_642/Y 0.21fF
C7264 INVX1_LOC_298/A INVX1_LOC_18/A 0.01fF
C7265 NAND2X1_LOC_553/A NOR2X1_LOC_791/B 0.02fF
C7266 NOR2X1_LOC_78/A NOR2X1_LOC_351/Y 0.01fF
C7267 INVX1_LOC_58/A NOR2X1_LOC_716/B 0.07fF
C7268 INVX1_LOC_22/A INVX1_LOC_47/Y 0.10fF
C7269 NOR2X1_LOC_303/Y NOR2X1_LOC_678/A 0.03fF
C7270 NAND2X1_LOC_638/Y INVX1_LOC_19/A 0.11fF
C7271 NOR2X1_LOC_762/a_36_216# INVX1_LOC_30/A 0.01fF
C7272 NOR2X1_LOC_581/a_36_216# INVX1_LOC_30/A 0.01fF
C7273 INVX1_LOC_45/A NOR2X1_LOC_698/a_36_216# 0.00fF
C7274 INVX1_LOC_176/A NAND2X1_LOC_96/A 0.02fF
C7275 INVX1_LOC_37/Y INVX1_LOC_46/A 0.00fF
C7276 NOR2X1_LOC_632/Y INVX1_LOC_4/A 0.01fF
C7277 D_INPUT_6 INVX1_LOC_18/A 0.00fF
C7278 NOR2X1_LOC_56/Y INVX1_LOC_118/A 0.08fF
C7279 NAND2X1_LOC_584/a_36_24# INVX1_LOC_296/A 0.01fF
C7280 NOR2X1_LOC_167/Y INVX1_LOC_285/A 0.02fF
C7281 NAND2X1_LOC_807/Y NAND2X1_LOC_74/B 0.07fF
C7282 NOR2X1_LOC_709/A NOR2X1_LOC_383/B 0.12fF
C7283 NOR2X1_LOC_382/Y INVX1_LOC_1/A 0.01fF
C7284 INVX1_LOC_11/A NOR2X1_LOC_389/A 0.28fF
C7285 NAND2X1_LOC_374/Y NOR2X1_LOC_693/Y 0.13fF
C7286 NOR2X1_LOC_721/A NOR2X1_LOC_720/A 0.14fF
C7287 NOR2X1_LOC_167/Y INVX1_LOC_265/Y 0.01fF
C7288 INVX1_LOC_21/A INVX1_LOC_181/Y 0.07fF
C7289 INVX1_LOC_288/Y INVX1_LOC_191/Y 0.01fF
C7290 NAND2X1_LOC_47/a_36_24# INVX1_LOC_174/A 0.00fF
C7291 NOR2X1_LOC_254/Y NOR2X1_LOC_678/A 0.03fF
C7292 NOR2X1_LOC_667/Y NOR2X1_LOC_816/A 0.03fF
C7293 NAND2X1_LOC_725/Y NAND2X1_LOC_722/A 0.47fF
C7294 INVX1_LOC_50/A NOR2X1_LOC_537/Y 0.03fF
C7295 NOR2X1_LOC_82/A NAND2X1_LOC_577/A 0.04fF
C7296 INVX1_LOC_25/Y INVX1_LOC_23/Y 0.13fF
C7297 INVX1_LOC_146/Y INVX1_LOC_118/A 0.03fF
C7298 NOR2X1_LOC_277/a_36_216# NOR2X1_LOC_278/A 0.02fF
C7299 NOR2X1_LOC_510/Y INVX1_LOC_49/A 0.07fF
C7300 NAND2X1_LOC_705/Y INVX1_LOC_24/A 0.02fF
C7301 NOR2X1_LOC_667/A NAND2X1_LOC_787/Y 0.03fF
C7302 VDD INVX1_LOC_118/A 2.61fF
C7303 NOR2X1_LOC_721/Y NAND2X1_LOC_63/Y 0.02fF
C7304 NOR2X1_LOC_15/Y NAND2X1_LOC_198/B 0.03fF
C7305 D_INPUT_0 INVX1_LOC_4/Y 0.10fF
C7306 NOR2X1_LOC_186/Y INVX1_LOC_33/A 0.08fF
C7307 NOR2X1_LOC_91/A NOR2X1_LOC_701/Y 0.01fF
C7308 NAND2X1_LOC_303/Y INVX1_LOC_24/A 3.13fF
C7309 NOR2X1_LOC_15/Y NAND2X1_LOC_368/a_36_24# 0.01fF
C7310 NOR2X1_LOC_137/A NOR2X1_LOC_334/Y 0.00fF
C7311 NOR2X1_LOC_298/Y NAND2X1_LOC_175/Y 0.09fF
C7312 NOR2X1_LOC_364/A INVX1_LOC_76/A 0.01fF
C7313 NAND2X1_LOC_538/Y NOR2X1_LOC_512/Y 0.03fF
C7314 NAND2X1_LOC_773/Y INVX1_LOC_314/Y 0.10fF
C7315 INVX1_LOC_290/A NOR2X1_LOC_638/Y 0.01fF
C7316 NOR2X1_LOC_251/a_36_216# INVX1_LOC_77/A -0.01fF
C7317 INVX1_LOC_78/Y INVX1_LOC_19/A 0.03fF
C7318 NAND2X1_LOC_741/B NOR2X1_LOC_599/Y 0.03fF
C7319 NAND2X1_LOC_733/Y NOR2X1_LOC_761/Y 0.12fF
C7320 NAND2X1_LOC_363/B NAND2X1_LOC_360/B 0.00fF
C7321 NAND2X1_LOC_267/B INVX1_LOC_46/Y 0.26fF
C7322 INVX1_LOC_6/A NAND2X1_LOC_74/B 0.16fF
C7323 NOR2X1_LOC_209/B INVX1_LOC_117/A 0.20fF
C7324 NAND2X1_LOC_544/a_36_24# NAND2X1_LOC_338/B 0.01fF
C7325 NAND2X1_LOC_573/Y INVX1_LOC_33/A 0.01fF
C7326 INVX1_LOC_268/A INVX1_LOC_105/Y 0.16fF
C7327 NOR2X1_LOC_82/A NAND2X1_LOC_656/A 0.02fF
C7328 INVX1_LOC_11/A NOR2X1_LOC_596/A 0.06fF
C7329 NOR2X1_LOC_857/A NOR2X1_LOC_445/B 0.06fF
C7330 NOR2X1_LOC_790/a_36_216# INVX1_LOC_33/A 0.00fF
C7331 INVX1_LOC_136/A INVX1_LOC_31/A 1.29fF
C7332 INVX1_LOC_21/A NAND2X1_LOC_563/Y 0.07fF
C7333 INVX1_LOC_312/A INVX1_LOC_312/Y 0.09fF
C7334 INVX1_LOC_306/A NAND2X1_LOC_99/A 0.03fF
C7335 NOR2X1_LOC_361/B INVX1_LOC_49/A 0.05fF
C7336 INVX1_LOC_224/Y NOR2X1_LOC_789/a_36_216# 0.00fF
C7337 INVX1_LOC_147/A INVX1_LOC_15/A 0.07fF
C7338 INVX1_LOC_76/A INVX1_LOC_285/A 0.10fF
C7339 INVX1_LOC_235/Y NOR2X1_LOC_6/B 0.07fF
C7340 NOR2X1_LOC_844/Y NOR2X1_LOC_859/A 0.09fF
C7341 INVX1_LOC_164/A INVX1_LOC_57/A 0.03fF
C7342 NAND2X1_LOC_190/Y NOR2X1_LOC_593/Y 0.15fF
C7343 INVX1_LOC_232/A NOR2X1_LOC_392/Y 0.14fF
C7344 INVX1_LOC_2/A NOR2X1_LOC_510/Y 0.11fF
C7345 NOR2X1_LOC_92/Y INVX1_LOC_162/Y 0.02fF
C7346 NOR2X1_LOC_798/A NOR2X1_LOC_767/a_36_216# 0.00fF
C7347 INVX1_LOC_206/Y INVX1_LOC_290/Y 0.07fF
C7348 INVX1_LOC_132/Y INVX1_LOC_26/Y 0.01fF
C7349 NOR2X1_LOC_357/Y NOR2X1_LOC_66/Y 0.06fF
C7350 INVX1_LOC_101/A INVX1_LOC_53/A 0.29fF
C7351 INVX1_LOC_83/A NOR2X1_LOC_809/A 0.01fF
C7352 INVX1_LOC_35/A INVX1_LOC_1/Y 0.04fF
C7353 NOR2X1_LOC_78/A INVX1_LOC_106/Y 0.01fF
C7354 NOR2X1_LOC_510/Y NOR2X1_LOC_226/A 0.00fF
C7355 NOR2X1_LOC_679/Y NOR2X1_LOC_577/Y 0.02fF
C7356 INVX1_LOC_58/A NOR2X1_LOC_717/B 0.01fF
C7357 NOR2X1_LOC_468/Y NOR2X1_LOC_52/B 0.12fF
C7358 NOR2X1_LOC_405/A INVX1_LOC_12/A 0.03fF
C7359 INVX1_LOC_18/A NAND2X1_LOC_16/Y 0.03fF
C7360 NAND2X1_LOC_140/A NOR2X1_LOC_125/Y 0.02fF
C7361 INVX1_LOC_256/A INVX1_LOC_63/Y 0.07fF
C7362 NOR2X1_LOC_591/Y NAND2X1_LOC_537/Y 0.08fF
C7363 NOR2X1_LOC_591/a_36_216# NAND2X1_LOC_538/Y 0.01fF
C7364 NOR2X1_LOC_389/A NOR2X1_LOC_433/A 0.22fF
C7365 INVX1_LOC_50/A INVX1_LOC_313/Y 0.12fF
C7366 NOR2X1_LOC_355/A INVX1_LOC_53/A 0.25fF
C7367 NAND2X1_LOC_581/Y NAND2X1_LOC_30/Y 0.03fF
C7368 NOR2X1_LOC_600/Y INVX1_LOC_290/Y 0.00fF
C7369 NOR2X1_LOC_852/B NOR2X1_LOC_590/A 0.04fF
C7370 INVX1_LOC_36/A NOR2X1_LOC_759/Y 0.02fF
C7371 INVX1_LOC_27/A NAND2X1_LOC_841/A 0.03fF
C7372 NOR2X1_LOC_32/B INVX1_LOC_135/A 0.10fF
C7373 INVX1_LOC_136/A INVX1_LOC_111/A 0.01fF
C7374 INVX1_LOC_202/A INVX1_LOC_36/A 0.10fF
C7375 INVX1_LOC_75/A INVX1_LOC_23/Y 0.07fF
C7376 INVX1_LOC_204/Y NAND2X1_LOC_480/a_36_24# 0.00fF
C7377 INVX1_LOC_299/A NAND2X1_LOC_118/a_36_24# 0.00fF
C7378 INVX1_LOC_13/A INVX1_LOC_13/Y 0.16fF
C7379 INVX1_LOC_30/A NOR2X1_LOC_625/Y 0.02fF
C7380 NOR2X1_LOC_536/A INVX1_LOC_27/Y 0.01fF
C7381 INVX1_LOC_75/A NAND2X1_LOC_72/a_36_24# 0.00fF
C7382 NOR2X1_LOC_689/A NAND2X1_LOC_863/A 0.01fF
C7383 NOR2X1_LOC_242/A NOR2X1_LOC_835/A 0.00fF
C7384 INVX1_LOC_201/Y NAND2X1_LOC_612/a_36_24# 0.00fF
C7385 NAND2X1_LOC_785/A INVX1_LOC_200/A 0.18fF
C7386 INVX1_LOC_37/A INVX1_LOC_49/Y 0.12fF
C7387 VDD NAND2X1_LOC_63/Y 2.50fF
C7388 INVX1_LOC_105/A INVX1_LOC_72/A 0.08fF
C7389 NOR2X1_LOC_226/A NOR2X1_LOC_361/B 0.10fF
C7390 INVX1_LOC_45/A NAND2X1_LOC_361/Y 0.07fF
C7391 INVX1_LOC_256/A NOR2X1_LOC_175/A 0.03fF
C7392 NOR2X1_LOC_112/a_36_216# NAND2X1_LOC_291/B 0.00fF
C7393 NAND2X1_LOC_740/Y INVX1_LOC_10/A 0.03fF
C7394 NOR2X1_LOC_637/Y NOR2X1_LOC_637/A 0.16fF
C7395 NOR2X1_LOC_389/A NOR2X1_LOC_52/B 0.11fF
C7396 NAND2X1_LOC_190/a_36_24# NOR2X1_LOC_717/B 0.00fF
C7397 NAND2X1_LOC_726/Y NAND2X1_LOC_724/A 0.03fF
C7398 INVX1_LOC_11/A INVX1_LOC_189/Y 0.02fF
C7399 NOR2X1_LOC_15/Y INVX1_LOC_53/Y 0.02fF
C7400 NAND2X1_LOC_736/Y NAND2X1_LOC_741/B 0.00fF
C7401 NAND2X1_LOC_468/B INVX1_LOC_32/A 1.00fF
C7402 NOR2X1_LOC_208/Y NOR2X1_LOC_759/Y 0.02fF
C7403 NAND2X1_LOC_350/A NAND2X1_LOC_470/a_36_24# 0.00fF
C7404 VDD NAND2X1_LOC_455/B 0.10fF
C7405 INVX1_LOC_58/A NOR2X1_LOC_151/Y 0.03fF
C7406 INVX1_LOC_11/A NOR2X1_LOC_220/A 0.08fF
C7407 INVX1_LOC_254/A INVX1_LOC_24/A 0.06fF
C7408 NOR2X1_LOC_91/A NOR2X1_LOC_165/a_36_216# 0.00fF
C7409 NOR2X1_LOC_483/B NOR2X1_LOC_209/Y 0.02fF
C7410 INVX1_LOC_202/A NOR2X1_LOC_208/Y 0.02fF
C7411 NOR2X1_LOC_605/B NAND2X1_LOC_724/A 0.05fF
C7412 NOR2X1_LOC_570/B NOR2X1_LOC_703/B 0.16fF
C7413 NOR2X1_LOC_15/Y NOR2X1_LOC_665/A 0.14fF
C7414 NOR2X1_LOC_846/Y NOR2X1_LOC_814/Y 0.04fF
C7415 INVX1_LOC_166/A NAND2X1_LOC_622/B 0.02fF
C7416 NOR2X1_LOC_433/A NOR2X1_LOC_596/A 0.06fF
C7417 NOR2X1_LOC_750/Y NAND2X1_LOC_348/A 0.01fF
C7418 NOR2X1_LOC_270/Y NOR2X1_LOC_142/Y 0.03fF
C7419 NAND2X1_LOC_655/A NAND2X1_LOC_175/Y 0.07fF
C7420 NAND2X1_LOC_642/Y NAND2X1_LOC_223/A 0.16fF
C7421 INVX1_LOC_74/A NOR2X1_LOC_38/B 0.17fF
C7422 INVX1_LOC_203/A NAND2X1_LOC_243/Y 0.03fF
C7423 NAND2X1_LOC_659/B NAND2X1_LOC_618/Y 0.02fF
C7424 INVX1_LOC_42/Y NOR2X1_LOC_717/A 0.08fF
C7425 NOR2X1_LOC_590/A INVX1_LOC_179/Y 0.08fF
C7426 NOR2X1_LOC_690/A INVX1_LOC_24/A 0.03fF
C7427 INVX1_LOC_269/A NOR2X1_LOC_719/B 0.01fF
C7428 NOR2X1_LOC_122/A NAND2X1_LOC_656/Y 0.01fF
C7429 INVX1_LOC_11/A NOR2X1_LOC_548/Y 0.08fF
C7430 INVX1_LOC_91/A NOR2X1_LOC_39/Y 0.46fF
C7431 NOR2X1_LOC_433/Y INVX1_LOC_186/Y 0.01fF
C7432 NOR2X1_LOC_798/A NOR2X1_LOC_174/A 0.01fF
C7433 INVX1_LOC_230/Y INVX1_LOC_316/Y 0.72fF
C7434 NAND2X1_LOC_559/Y NOR2X1_LOC_576/B 0.25fF
C7435 VDD NAND2X1_LOC_618/Y 0.53fF
C7436 NOR2X1_LOC_575/Y INVX1_LOC_242/A 0.18fF
C7437 NOR2X1_LOC_67/Y INVX1_LOC_9/A 0.09fF
C7438 INVX1_LOC_33/A NOR2X1_LOC_374/A 0.03fF
C7439 NAND2X1_LOC_803/B NOR2X1_LOC_561/Y 0.03fF
C7440 NOR2X1_LOC_274/a_36_216# NOR2X1_LOC_309/Y 0.00fF
C7441 INVX1_LOC_49/A INVX1_LOC_153/Y 0.01fF
C7442 NOR2X1_LOC_596/A NOR2X1_LOC_52/B 0.05fF
C7443 NAND2X1_LOC_149/Y NOR2X1_LOC_156/A 0.06fF
C7444 D_INPUT_2 NOR2X1_LOC_143/a_36_216# 0.00fF
C7445 NOR2X1_LOC_307/B INVX1_LOC_142/A 0.12fF
C7446 INVX1_LOC_147/Y NAND2X1_LOC_61/Y 0.36fF
C7447 INVX1_LOC_161/Y NAND2X1_LOC_656/Y 0.07fF
C7448 INVX1_LOC_27/Y INVX1_LOC_3/A 0.14fF
C7449 NAND2X1_LOC_363/B NOR2X1_LOC_837/A 0.02fF
C7450 INVX1_LOC_75/A NOR2X1_LOC_249/Y 0.29fF
C7451 INVX1_LOC_77/A INVX1_LOC_104/A 0.67fF
C7452 NOR2X1_LOC_361/B INPUT_1 0.04fF
C7453 NOR2X1_LOC_388/Y INVX1_LOC_155/Y 0.00fF
C7454 NAND2X1_LOC_364/A NOR2X1_LOC_566/Y 0.00fF
C7455 INVX1_LOC_185/A INVX1_LOC_42/A 0.03fF
C7456 NOR2X1_LOC_590/A NOR2X1_LOC_561/Y 0.09fF
C7457 INVX1_LOC_225/A INVX1_LOC_33/A 0.07fF
C7458 NOR2X1_LOC_590/A INVX1_LOC_7/A 0.09fF
C7459 VDD NOR2X1_LOC_631/Y 0.26fF
C7460 NOR2X1_LOC_288/A INVX1_LOC_33/A 0.12fF
C7461 INVX1_LOC_41/A INVX1_LOC_162/Y 0.00fF
C7462 NAND2X1_LOC_288/a_36_24# NOR2X1_LOC_743/Y 0.00fF
C7463 INVX1_LOC_87/A NOR2X1_LOC_107/a_36_216# 0.00fF
C7464 INVX1_LOC_13/A NOR2X1_LOC_500/B 0.02fF
C7465 INVX1_LOC_286/Y INPUT_5 0.27fF
C7466 INVX1_LOC_49/A INVX1_LOC_177/A 0.10fF
C7467 INVX1_LOC_41/A INVX1_LOC_85/A 0.00fF
C7468 NOR2X1_LOC_714/Y NOR2X1_LOC_374/A 0.01fF
C7469 NOR2X1_LOC_795/Y NOR2X1_LOC_551/B 0.00fF
C7470 INVX1_LOC_136/A NAND2X1_LOC_859/Y 0.10fF
C7471 INVX1_LOC_217/A NOR2X1_LOC_86/A 0.04fF
C7472 NAND2X1_LOC_53/Y INVX1_LOC_311/Y 0.01fF
C7473 INVX1_LOC_227/Y NOR2X1_LOC_569/Y 0.20fF
C7474 INVX1_LOC_54/Y NAND2X1_LOC_536/a_36_24# 0.01fF
C7475 NAND2X1_LOC_391/Y INVX1_LOC_286/A 0.00fF
C7476 INVX1_LOC_2/A INVX1_LOC_153/Y 0.01fF
C7477 NAND2X1_LOC_83/a_36_24# NOR2X1_LOC_649/B 0.01fF
C7478 NOR2X1_LOC_474/A NOR2X1_LOC_399/Y 0.00fF
C7479 NOR2X1_LOC_617/Y NAND2X1_LOC_859/B 0.02fF
C7480 NOR2X1_LOC_573/Y NOR2X1_LOC_575/Y 0.11fF
C7481 INVX1_LOC_132/A INVX1_LOC_40/A 0.01fF
C7482 INVX1_LOC_48/Y NOR2X1_LOC_391/Y -0.01fF
C7483 INVX1_LOC_46/A INVX1_LOC_29/Y 0.10fF
C7484 INVX1_LOC_18/A NOR2X1_LOC_686/B 0.01fF
C7485 NOR2X1_LOC_220/A NOR2X1_LOC_593/Y 0.49fF
C7486 INVX1_LOC_174/Y NOR2X1_LOC_705/a_36_216# 0.00fF
C7487 INVX1_LOC_304/Y NAND2X1_LOC_785/A 0.01fF
C7488 NOR2X1_LOC_372/Y NOR2X1_LOC_71/Y 0.01fF
C7489 INVX1_LOC_135/A INVX1_LOC_195/Y 0.01fF
C7490 NOR2X1_LOC_174/B NOR2X1_LOC_500/B 0.09fF
C7491 NAND2X1_LOC_550/A NOR2X1_LOC_322/Y 0.02fF
C7492 NAND2X1_LOC_141/Y INVX1_LOC_32/A 0.04fF
C7493 NOR2X1_LOC_445/Y NOR2X1_LOC_500/Y 0.01fF
C7494 INVX1_LOC_46/Y INVX1_LOC_4/Y 0.10fF
C7495 INVX1_LOC_2/A INVX1_LOC_177/A 0.03fF
C7496 INVX1_LOC_136/A NAND2X1_LOC_866/B 0.07fF
C7497 VDD INVX1_LOC_138/A 0.12fF
C7498 INVX1_LOC_58/A NOR2X1_LOC_322/a_36_216# 0.00fF
C7499 INVX1_LOC_11/A INVX1_LOC_51/Y 0.03fF
C7500 INVX1_LOC_232/Y NOR2X1_LOC_84/Y 0.01fF
C7501 NOR2X1_LOC_437/Y NAND2X1_LOC_656/Y 0.04fF
C7502 INVX1_LOC_255/Y NAND2X1_LOC_276/Y 0.21fF
C7503 NAND2X1_LOC_579/A NOR2X1_LOC_45/B 0.08fF
C7504 INVX1_LOC_27/A INVX1_LOC_95/Y 1.01fF
C7505 INVX1_LOC_90/A NOR2X1_LOC_91/Y 0.05fF
C7506 NAND2X1_LOC_861/Y INVX1_LOC_41/Y 0.00fF
C7507 NAND2X1_LOC_36/A D_INPUT_4 0.07fF
C7508 INVX1_LOC_41/A NOR2X1_LOC_730/Y 0.02fF
C7509 INVX1_LOC_136/A NAND2X1_LOC_807/Y 0.02fF
C7510 NOR2X1_LOC_785/Y INVX1_LOC_49/A 0.02fF
C7511 INVX1_LOC_232/Y INVX1_LOC_216/A 1.00fF
C7512 INVX1_LOC_107/Y NOR2X1_LOC_158/Y 0.03fF
C7513 NOR2X1_LOC_590/A NOR2X1_LOC_835/B 0.00fF
C7514 INVX1_LOC_12/A INVX1_LOC_109/Y 0.07fF
C7515 NAND2X1_LOC_561/a_36_24# NOR2X1_LOC_536/A 0.00fF
C7516 NOR2X1_LOC_276/Y INVX1_LOC_6/A 0.03fF
C7517 INVX1_LOC_34/A NOR2X1_LOC_757/A 0.03fF
C7518 NAND2X1_LOC_852/a_36_24# NAND2X1_LOC_852/Y 0.03fF
C7519 NOR2X1_LOC_219/Y INVX1_LOC_96/Y 0.77fF
C7520 NOR2X1_LOC_471/Y NOR2X1_LOC_377/a_36_216# 0.00fF
C7521 NAND2X1_LOC_514/Y NOR2X1_LOC_329/B 0.04fF
C7522 NOR2X1_LOC_831/B NOR2X1_LOC_301/A 0.01fF
C7523 NAND2X1_LOC_722/A NOR2X1_LOC_165/Y 0.25fF
C7524 NOR2X1_LOC_590/A INVX1_LOC_303/Y 0.01fF
C7525 NOR2X1_LOC_32/B INVX1_LOC_280/A 0.05fF
C7526 NOR2X1_LOC_32/B NOR2X1_LOC_94/Y 0.13fF
C7527 INVX1_LOC_299/A NOR2X1_LOC_542/B 0.01fF
C7528 NOR2X1_LOC_690/A NOR2X1_LOC_525/a_36_216# 0.16fF
C7529 INVX1_LOC_39/A VDD 1.45fF
C7530 INVX1_LOC_282/Y GATE_865 0.52fF
C7531 NOR2X1_LOC_453/Y INVX1_LOC_115/A 0.00fF
C7532 NAND2X1_LOC_798/a_36_24# INVX1_LOC_90/A 0.00fF
C7533 INVX1_LOC_104/A NOR2X1_LOC_549/a_36_216# 0.00fF
C7534 NAND2X1_LOC_361/Y NOR2X1_LOC_749/Y 0.00fF
C7535 INVX1_LOC_266/A NOR2X1_LOC_35/Y 0.10fF
C7536 NOR2X1_LOC_589/A INVX1_LOC_133/Y 0.07fF
C7537 INVX1_LOC_96/Y NOR2X1_LOC_665/A 0.50fF
C7538 NAND2X1_LOC_466/Y NOR2X1_LOC_130/A 0.01fF
C7539 INVX1_LOC_5/A NOR2X1_LOC_536/A 0.03fF
C7540 INVX1_LOC_299/A INVX1_LOC_143/Y 0.02fF
C7541 INVX1_LOC_223/A NAND2X1_LOC_309/a_36_24# 0.01fF
C7542 NOR2X1_LOC_132/Y INPUT_1 0.01fF
C7543 NOR2X1_LOC_781/Y INVX1_LOC_302/Y 0.01fF
C7544 NOR2X1_LOC_360/Y NOR2X1_LOC_74/A 0.07fF
C7545 NAND2X1_LOC_715/B INVX1_LOC_118/Y 0.02fF
C7546 INVX1_LOC_136/A INVX1_LOC_6/A 0.11fF
C7547 INVX1_LOC_38/Y INVX1_LOC_230/A 0.01fF
C7548 NAND2X1_LOC_222/A NOR2X1_LOC_673/A 0.01fF
C7549 NOR2X1_LOC_360/Y NOR2X1_LOC_9/Y 0.03fF
C7550 NOR2X1_LOC_778/B INVX1_LOC_279/A 0.01fF
C7551 INVX1_LOC_178/A NOR2X1_LOC_536/A 0.06fF
C7552 NOR2X1_LOC_328/Y INVX1_LOC_22/A 0.03fF
C7553 NOR2X1_LOC_226/A NAND2X1_LOC_573/A 0.07fF
C7554 INVX1_LOC_35/A INVX1_LOC_117/Y 0.03fF
C7555 NOR2X1_LOC_615/a_36_216# INVX1_LOC_20/A 0.00fF
C7556 NAND2X1_LOC_803/B INVX1_LOC_76/A 0.02fF
C7557 INVX1_LOC_5/A NOR2X1_LOC_655/Y 0.02fF
C7558 NOR2X1_LOC_15/Y INVX1_LOC_77/Y 0.02fF
C7559 NOR2X1_LOC_763/Y INVX1_LOC_243/A 0.02fF
C7560 NOR2X1_LOC_329/B NAND2X1_LOC_332/Y 0.03fF
C7561 NAND2X1_LOC_254/Y NOR2X1_LOC_38/B 0.01fF
C7562 NAND2X1_LOC_149/Y NOR2X1_LOC_684/Y 0.08fF
C7563 NOR2X1_LOC_510/Y INVX1_LOC_118/A 0.05fF
C7564 INVX1_LOC_30/Y INVX1_LOC_16/A 0.07fF
C7565 NOR2X1_LOC_82/A NOR2X1_LOC_42/a_36_216# 0.00fF
C7566 NOR2X1_LOC_383/Y INVX1_LOC_25/Y 0.07fF
C7567 NOR2X1_LOC_550/B NOR2X1_LOC_208/A 0.03fF
C7568 NOR2X1_LOC_78/B NOR2X1_LOC_355/A 0.03fF
C7569 INVX1_LOC_99/A NAND2X1_LOC_72/B 0.01fF
C7570 NAND2X1_LOC_374/Y NOR2X1_LOC_71/Y 0.14fF
C7571 INVX1_LOC_5/A NAND2X1_LOC_93/B 0.07fF
C7572 INVX1_LOC_298/Y INVX1_LOC_29/A 0.02fF
C7573 INVX1_LOC_159/A NOR2X1_LOC_7/Y 0.01fF
C7574 NOR2X1_LOC_439/a_36_216# INVX1_LOC_279/A 0.00fF
C7575 NAND2X1_LOC_391/Y INVX1_LOC_54/A 0.00fF
C7576 NOR2X1_LOC_494/Y NOR2X1_LOC_536/A 0.07fF
C7577 NOR2X1_LOC_727/B INVX1_LOC_19/A 0.03fF
C7578 NOR2X1_LOC_590/A INVX1_LOC_76/A 0.30fF
C7579 NAND2X1_LOC_541/Y INVX1_LOC_89/A 0.01fF
C7580 INVX1_LOC_88/A INVX1_LOC_66/Y 0.32fF
C7581 NOR2X1_LOC_238/Y NOR2X1_LOC_528/Y 0.16fF
C7582 NOR2X1_LOC_456/Y INVX1_LOC_63/A 0.12fF
C7583 NOR2X1_LOC_638/Y INVX1_LOC_261/Y 0.01fF
C7584 INVX1_LOC_55/Y NOR2X1_LOC_203/Y 0.30fF
C7585 NAND2X1_LOC_291/B NOR2X1_LOC_342/B 0.01fF
C7586 INVX1_LOC_83/A NOR2X1_LOC_160/Y 0.03fF
C7587 INVX1_LOC_208/A NOR2X1_LOC_473/B 0.10fF
C7588 INVX1_LOC_227/A NOR2X1_LOC_561/Y 0.10fF
C7589 NOR2X1_LOC_78/B NOR2X1_LOC_736/Y 0.05fF
C7590 NOR2X1_LOC_551/a_36_216# INVX1_LOC_177/A 0.00fF
C7591 NAND2X1_LOC_337/B NOR2X1_LOC_536/A 0.08fF
C7592 NOR2X1_LOC_361/B INVX1_LOC_118/A 0.80fF
C7593 INVX1_LOC_179/Y NOR2X1_LOC_703/A 0.02fF
C7594 NAND2X1_LOC_741/B NAND2X1_LOC_453/A 0.05fF
C7595 INVX1_LOC_5/A NOR2X1_LOC_649/B 0.07fF
C7596 NOR2X1_LOC_816/A NOR2X1_LOC_536/A 0.12fF
C7597 INVX1_LOC_5/A INVX1_LOC_3/A 0.25fF
C7598 NOR2X1_LOC_458/B INVX1_LOC_182/A 0.01fF
C7599 INVX1_LOC_19/A NOR2X1_LOC_717/A 0.03fF
C7600 NOR2X1_LOC_596/A INVX1_LOC_199/A 0.11fF
C7601 NAND2X1_LOC_213/A INVX1_LOC_92/A 0.04fF
C7602 NAND2X1_LOC_552/A NOR2X1_LOC_661/A 0.03fF
C7603 NAND2X1_LOC_859/Y NAND2X1_LOC_862/Y 0.17fF
C7604 INVX1_LOC_6/A NOR2X1_LOC_278/A 0.07fF
C7605 NOR2X1_LOC_717/Y NAND2X1_LOC_472/Y 0.01fF
C7606 INVX1_LOC_49/A INVX1_LOC_65/A 0.08fF
C7607 NOR2X1_LOC_34/B NOR2X1_LOC_814/A 0.07fF
C7608 NOR2X1_LOC_644/A NOR2X1_LOC_553/B 0.03fF
C7609 INVX1_LOC_178/A NOR2X1_LOC_649/B 0.02fF
C7610 INVX1_LOC_61/A VDD 0.00fF
C7611 INVX1_LOC_13/Y NAND2X1_LOC_489/Y 0.02fF
C7612 INVX1_LOC_2/A INVX1_LOC_285/Y 0.03fF
C7613 INVX1_LOC_33/A NAND2X1_LOC_642/Y 0.06fF
C7614 NOR2X1_LOC_45/Y NOR2X1_LOC_351/Y 0.01fF
C7615 INVX1_LOC_75/A INVX1_LOC_232/A 0.07fF
C7616 NAND2X1_LOC_74/B NOR2X1_LOC_109/Y 0.07fF
C7617 NOR2X1_LOC_597/A INVX1_LOC_10/A 0.04fF
C7618 NAND2X1_LOC_515/a_36_24# NAND2X1_LOC_211/Y 0.01fF
C7619 NOR2X1_LOC_754/Y INVX1_LOC_42/A 0.01fF
C7620 INVX1_LOC_272/Y NOR2X1_LOC_88/Y 0.07fF
C7621 INVX1_LOC_17/A NOR2X1_LOC_831/B 0.72fF
C7622 NOR2X1_LOC_773/Y INVX1_LOC_126/Y 0.52fF
C7623 NOR2X1_LOC_500/Y NOR2X1_LOC_335/B 0.06fF
C7624 INVX1_LOC_279/A NAND2X1_LOC_123/Y 0.01fF
C7625 NAND2X1_LOC_18/a_36_24# INPUT_7 0.00fF
C7626 NAND2X1_LOC_862/Y NAND2X1_LOC_866/B 0.01fF
C7627 INVX1_LOC_215/A INVX1_LOC_79/A 0.06fF
C7628 INVX1_LOC_21/A NOR2X1_LOC_509/A 0.01fF
C7629 NAND2X1_LOC_562/Y NAND2X1_LOC_659/B 0.04fF
C7630 NOR2X1_LOC_334/Y NOR2X1_LOC_383/B 0.21fF
C7631 NAND2X1_LOC_325/Y INVX1_LOC_20/A 0.03fF
C7632 NOR2X1_LOC_401/B INVX1_LOC_98/A 0.06fF
C7633 NOR2X1_LOC_433/A NOR2X1_LOC_447/B 0.01fF
C7634 NAND2X1_LOC_647/B INVX1_LOC_23/A 0.02fF
C7635 NAND2X1_LOC_740/Y INVX1_LOC_12/A 0.03fF
C7636 NAND2X1_LOC_662/B NAND2X1_LOC_662/Y 0.00fF
C7637 NOR2X1_LOC_91/Y INVX1_LOC_38/A 0.10fF
C7638 NOR2X1_LOC_815/Y VDD 0.31fF
C7639 INVX1_LOC_177/Y INVX1_LOC_9/A 0.22fF
C7640 NAND2X1_LOC_354/B INVX1_LOC_76/A 0.01fF
C7641 INVX1_LOC_272/Y INVX1_LOC_84/A 0.03fF
C7642 NOR2X1_LOC_52/B NAND2X1_LOC_655/B 0.01fF
C7643 INVX1_LOC_78/A INVX1_LOC_270/Y 0.08fF
C7644 INVX1_LOC_271/A INVX1_LOC_271/Y 0.00fF
C7645 NOR2X1_LOC_6/B NOR2X1_LOC_35/Y 0.01fF
C7646 NOR2X1_LOC_52/B NAND2X1_LOC_469/B 0.06fF
C7647 INVX1_LOC_208/A NOR2X1_LOC_355/B 0.00fF
C7648 NAND2X1_LOC_53/Y INVX1_LOC_84/A 0.07fF
C7649 INPUT_2 NAND2X1_LOC_574/A 0.10fF
C7650 INPUT_3 NAND2X1_LOC_141/Y 0.27fF
C7651 INVX1_LOC_69/Y NOR2X1_LOC_188/a_36_216# 0.01fF
C7652 NAND2X1_LOC_286/B NOR2X1_LOC_318/A 0.17fF
C7653 NOR2X1_LOC_624/A VDD 0.24fF
C7654 NOR2X1_LOC_372/Y NAND2X1_LOC_243/Y 0.01fF
C7655 INVX1_LOC_14/A NAND2X1_LOC_773/B 0.20fF
C7656 NOR2X1_LOC_335/B INVX1_LOC_10/A 0.06fF
C7657 NOR2X1_LOC_209/Y NOR2X1_LOC_486/Y 0.07fF
C7658 NAND2X1_LOC_562/Y VDD 0.01fF
C7659 INVX1_LOC_34/A INVX1_LOC_37/A 0.38fF
C7660 D_INPUT_1 NAND2X1_LOC_454/Y 0.01fF
C7661 NOR2X1_LOC_808/A NOR2X1_LOC_324/A 0.00fF
C7662 INVX1_LOC_136/A NOR2X1_LOC_79/A 0.04fF
C7663 INVX1_LOC_18/A NOR2X1_LOC_433/Y 0.03fF
C7664 NOR2X1_LOC_483/B NAND2X1_LOC_252/a_36_24# 0.02fF
C7665 INVX1_LOC_40/A NAND2X1_LOC_642/Y 0.03fF
C7666 NOR2X1_LOC_220/A NOR2X1_LOC_601/Y 0.01fF
C7667 NAND2X1_LOC_364/A INVX1_LOC_92/A 0.07fF
C7668 INVX1_LOC_13/Y INVX1_LOC_32/A 0.13fF
C7669 INPUT_3 NOR2X1_LOC_820/B 0.01fF
C7670 INVX1_LOC_276/A INVX1_LOC_20/A 0.03fF
C7671 INVX1_LOC_18/A NAND2X1_LOC_798/B 0.07fF
C7672 NOR2X1_LOC_370/a_36_216# INVX1_LOC_69/Y 0.01fF
C7673 INVX1_LOC_312/Y NOR2X1_LOC_841/A 0.10fF
C7674 NOR2X1_LOC_65/B INVX1_LOC_270/Y 0.17fF
C7675 NOR2X1_LOC_598/B NAND2X1_LOC_91/a_36_24# 0.08fF
C7676 NOR2X1_LOC_318/B NOR2X1_LOC_188/Y 0.04fF
C7677 INVX1_LOC_230/Y NOR2X1_LOC_662/A 0.03fF
C7678 INVX1_LOC_182/Y NAND2X1_LOC_123/Y 0.08fF
C7679 NOR2X1_LOC_67/A INVX1_LOC_20/A 0.40fF
C7680 INVX1_LOC_33/A NOR2X1_LOC_271/Y 0.01fF
C7681 NAND2X1_LOC_56/a_36_24# INVX1_LOC_186/Y 0.01fF
C7682 INVX1_LOC_16/A NOR2X1_LOC_124/A 0.05fF
C7683 NOR2X1_LOC_226/A NAND2X1_LOC_267/B 0.00fF
C7684 NOR2X1_LOC_152/Y INVX1_LOC_185/A 0.00fF
C7685 INVX1_LOC_5/A NAND2X1_LOC_470/B 0.03fF
C7686 NOR2X1_LOC_820/A NOR2X1_LOC_820/Y 0.01fF
C7687 INVX1_LOC_224/A NAND2X1_LOC_200/a_36_24# 0.00fF
C7688 NAND2X1_LOC_733/B VDD 0.33fF
C7689 INVX1_LOC_95/Y INVX1_LOC_137/A 0.01fF
C7690 NAND2X1_LOC_562/B NOR2X1_LOC_536/A 0.03fF
C7691 NOR2X1_LOC_637/Y NAND2X1_LOC_798/B 0.00fF
C7692 NAND2X1_LOC_735/B NAND2X1_LOC_659/B 0.03fF
C7693 NOR2X1_LOC_78/B NOR2X1_LOC_111/A 0.09fF
C7694 NOR2X1_LOC_392/Y INVX1_LOC_112/Y 0.02fF
C7695 INVX1_LOC_279/A NOR2X1_LOC_657/B 0.36fF
C7696 NOR2X1_LOC_553/B NOR2X1_LOC_540/B 0.03fF
C7697 NAND2X1_LOC_227/Y NOR2X1_LOC_226/Y 0.10fF
C7698 INVX1_LOC_104/A INVX1_LOC_9/A 0.15fF
C7699 D_INPUT_0 NOR2X1_LOC_595/Y 0.02fF
C7700 INVX1_LOC_89/A NOR2X1_LOC_78/A 2.79fF
C7701 NOR2X1_LOC_546/a_36_216# NAND2X1_LOC_425/Y 0.01fF
C7702 INVX1_LOC_26/A INVX1_LOC_306/Y 0.03fF
C7703 INVX1_LOC_88/A INVX1_LOC_32/A 0.22fF
C7704 NOR2X1_LOC_551/B NOR2X1_LOC_862/B 0.02fF
C7705 VDD NAND2X1_LOC_735/B 0.47fF
C7706 NAND2X1_LOC_802/A NOR2X1_LOC_697/Y 0.01fF
C7707 NOR2X1_LOC_667/Y INVX1_LOC_42/A 0.17fF
C7708 INVX1_LOC_36/A NAND2X1_LOC_74/B 0.10fF
C7709 NAND2X1_LOC_53/Y INVX1_LOC_15/A 0.07fF
C7710 NAND2X1_LOC_508/A NOR2X1_LOC_78/A 0.03fF
C7711 NOR2X1_LOC_773/Y NOR2X1_LOC_536/A 0.18fF
C7712 NOR2X1_LOC_192/A NAND2X1_LOC_842/B 0.01fF
C7713 NOR2X1_LOC_751/Y INVX1_LOC_125/A 0.01fF
C7714 NOR2X1_LOC_377/Y NAND2X1_LOC_93/B 0.02fF
C7715 INVX1_LOC_36/A NAND2X1_LOC_207/Y 0.39fF
C7716 INVX1_LOC_213/Y NOR2X1_LOC_676/Y 0.02fF
C7717 NOR2X1_LOC_445/Y NOR2X1_LOC_445/B 0.08fF
C7718 VDD INPUT_5 0.52fF
C7719 NOR2X1_LOC_274/Y NOR2X1_LOC_814/A 0.06fF
C7720 INVX1_LOC_316/A INPUT_1 0.03fF
C7721 INVX1_LOC_247/Y INVX1_LOC_29/A 0.09fF
C7722 INVX1_LOC_40/A NOR2X1_LOC_271/Y 1.29fF
C7723 INVX1_LOC_280/Y INVX1_LOC_118/A 0.03fF
C7724 INVX1_LOC_75/A NOR2X1_LOC_685/A 0.01fF
C7725 INVX1_LOC_315/A NOR2X1_LOC_820/Y 0.11fF
C7726 NOR2X1_LOC_377/Y NAND2X1_LOC_425/Y 0.01fF
C7727 NOR2X1_LOC_533/Y INVX1_LOC_94/Y 0.01fF
C7728 INVX1_LOC_16/A NOR2X1_LOC_684/Y 0.08fF
C7729 NOR2X1_LOC_13/Y INVX1_LOC_19/A 0.07fF
C7730 INVX1_LOC_28/A NOR2X1_LOC_124/A 0.02fF
C7731 NOR2X1_LOC_96/a_36_216# INVX1_LOC_316/Y 0.00fF
C7732 NAND2X1_LOC_231/Y NOR2X1_LOC_743/Y 0.01fF
C7733 NOR2X1_LOC_798/A INVX1_LOC_29/Y 0.76fF
C7734 NAND2X1_LOC_374/Y NAND2X1_LOC_243/Y 0.00fF
C7735 NOR2X1_LOC_148/B INVX1_LOC_37/A 0.01fF
C7736 NOR2X1_LOC_516/B NOR2X1_LOC_54/a_36_216# 0.00fF
C7737 NAND2X1_LOC_11/Y INVX1_LOC_92/A 0.00fF
C7738 NAND2X1_LOC_364/Y INVX1_LOC_19/A 0.03fF
C7739 NAND2X1_LOC_562/B NOR2X1_LOC_649/B 0.09fF
C7740 NOR2X1_LOC_430/A NOR2X1_LOC_11/Y 0.11fF
C7741 NOR2X1_LOC_272/Y INVX1_LOC_53/A 0.14fF
C7742 INVX1_LOC_75/A INVX1_LOC_74/Y 0.06fF
C7743 NOR2X1_LOC_237/Y NAND2X1_LOC_74/B 0.26fF
C7744 NOR2X1_LOC_234/a_36_216# NAND2X1_LOC_489/Y 0.01fF
C7745 NOR2X1_LOC_709/A NAND2X1_LOC_267/a_36_24# 0.07fF
C7746 NOR2X1_LOC_500/B NOR2X1_LOC_623/B 0.40fF
C7747 INVX1_LOC_75/A NAND2X1_LOC_447/Y 0.03fF
C7748 INVX1_LOC_278/A NAND2X1_LOC_474/Y 0.01fF
C7749 INVX1_LOC_286/A INVX1_LOC_91/A 0.17fF
C7750 NOR2X1_LOC_703/Y NOR2X1_LOC_78/A 0.03fF
C7751 NOR2X1_LOC_795/Y NOR2X1_LOC_691/A 0.40fF
C7752 INVX1_LOC_132/A INVX1_LOC_106/Y 0.00fF
C7753 INVX1_LOC_13/A NOR2X1_LOC_99/Y 0.14fF
C7754 NOR2X1_LOC_772/B INVX1_LOC_171/Y 0.13fF
C7755 INVX1_LOC_63/Y NOR2X1_LOC_89/A 1.90fF
C7756 NOR2X1_LOC_590/A NOR2X1_LOC_447/A 0.01fF
C7757 NOR2X1_LOC_272/a_36_216# NOR2X1_LOC_510/Y 0.00fF
C7758 NOR2X1_LOC_309/Y NAND2X1_LOC_74/B 0.07fF
C7759 NOR2X1_LOC_332/A NOR2X1_LOC_655/Y 0.02fF
C7760 NOR2X1_LOC_757/Y NAND2X1_LOC_475/Y 0.11fF
C7761 INVX1_LOC_233/Y INVX1_LOC_229/A 0.05fF
C7762 NOR2X1_LOC_124/B INVX1_LOC_284/A 0.06fF
C7763 NAND2X1_LOC_709/a_36_24# INVX1_LOC_117/A 0.01fF
C7764 NOR2X1_LOC_773/Y NOR2X1_LOC_661/A 0.18fF
C7765 INVX1_LOC_303/A INVX1_LOC_32/A 0.07fF
C7766 INVX1_LOC_230/Y INVX1_LOC_57/A 0.07fF
C7767 NOR2X1_LOC_636/a_36_216# NOR2X1_LOC_48/B 0.00fF
C7768 INPUT_0 INVX1_LOC_37/A 0.14fF
C7769 NOR2X1_LOC_500/Y INVX1_LOC_84/A 0.07fF
C7770 NAND2X1_LOC_650/B NOR2X1_LOC_167/Y 0.27fF
C7771 INVX1_LOC_226/Y INVX1_LOC_84/A 0.98fF
C7772 INVX1_LOC_140/A NOR2X1_LOC_536/A 0.03fF
C7773 INVX1_LOC_21/A NOR2X1_LOC_61/B 0.03fF
C7774 INVX1_LOC_10/A NOR2X1_LOC_88/Y 0.59fF
C7775 INVX1_LOC_256/Y INVX1_LOC_19/A 0.05fF
C7776 INVX1_LOC_35/A NOR2X1_LOC_82/A 0.07fF
C7777 INVX1_LOC_58/A NOR2X1_LOC_644/B 0.03fF
C7778 INVX1_LOC_288/Y INVX1_LOC_36/A 0.02fF
C7779 NOR2X1_LOC_607/a_36_216# NOR2X1_LOC_334/Y 0.00fF
C7780 INVX1_LOC_96/A NOR2X1_LOC_35/Y 0.45fF
C7781 NOR2X1_LOC_226/A NAND2X1_LOC_81/B 0.07fF
C7782 INVX1_LOC_45/A INVX1_LOC_50/A 0.28fF
C7783 INVX1_LOC_249/A INVX1_LOC_271/Y 0.03fF
C7784 INVX1_LOC_50/A NOR2X1_LOC_568/A 0.07fF
C7785 NAND2X1_LOC_773/Y INVX1_LOC_27/A 0.39fF
C7786 NOR2X1_LOC_706/A INVX1_LOC_193/A -0.00fF
C7787 NAND2X1_LOC_46/a_36_24# NAND2X1_LOC_555/Y 0.00fF
C7788 INVX1_LOC_6/Y INVX1_LOC_271/Y 0.04fF
C7789 NOR2X1_LOC_7/Y VDD 0.14fF
C7790 NOR2X1_LOC_272/a_36_216# NOR2X1_LOC_361/B 0.00fF
C7791 INVX1_LOC_21/A INVX1_LOC_101/Y 0.01fF
C7792 INVX1_LOC_136/A INVX1_LOC_270/A 0.08fF
C7793 INVX1_LOC_39/A NOR2X1_LOC_361/B 0.03fF
C7794 INVX1_LOC_235/Y NOR2X1_LOC_15/Y 0.23fF
C7795 INVX1_LOC_256/A INVX1_LOC_5/A 0.08fF
C7796 D_GATE_366 NOR2X1_LOC_155/A 4.84fF
C7797 INVX1_LOC_10/A INVX1_LOC_84/A 0.07fF
C7798 NOR2X1_LOC_542/Y NOR2X1_LOC_445/B -0.00fF
C7799 NAND2X1_LOC_149/Y NOR2X1_LOC_15/Y 0.08fF
C7800 NOR2X1_LOC_78/A NOR2X1_LOC_52/a_36_216# 0.00fF
C7801 NOR2X1_LOC_296/Y INVX1_LOC_13/Y 0.28fF
C7802 NOR2X1_LOC_332/A NOR2X1_LOC_649/B 0.04fF
C7803 INVX1_LOC_199/A NAND2X1_LOC_469/B 0.02fF
C7804 NOR2X1_LOC_332/A INVX1_LOC_3/A 0.14fF
C7805 NOR2X1_LOC_244/B NAND2X1_LOC_291/B 0.01fF
C7806 INVX1_LOC_168/A INVX1_LOC_32/A 0.10fF
C7807 INVX1_LOC_35/A NAND2X1_LOC_36/A 0.01fF
C7808 NAND2X1_LOC_21/Y NOR2X1_LOC_36/A 0.33fF
C7809 VDD NOR2X1_LOC_448/A -0.00fF
C7810 D_INPUT_1 NOR2X1_LOC_68/A 0.03fF
C7811 NOR2X1_LOC_311/Y NOR2X1_LOC_111/A 0.03fF
C7812 NAND2X1_LOC_361/Y NOR2X1_LOC_621/B 0.06fF
C7813 NOR2X1_LOC_373/Y INVX1_LOC_203/A 0.04fF
C7814 NAND2X1_LOC_450/a_36_24# INVX1_LOC_38/A 0.00fF
C7815 NOR2X1_LOC_91/A NAND2X1_LOC_567/Y 0.08fF
C7816 NOR2X1_LOC_590/A NOR2X1_LOC_434/Y 0.41fF
C7817 NOR2X1_LOC_332/A NOR2X1_LOC_814/a_36_216# 0.01fF
C7818 INVX1_LOC_27/A INVX1_LOC_252/Y 0.05fF
C7819 NAND2X1_LOC_364/A INVX1_LOC_53/A 0.14fF
C7820 NAND2X1_LOC_364/Y INVX1_LOC_26/Y 0.01fF
C7821 INVX1_LOC_50/A INVX1_LOC_71/A 0.10fF
C7822 NAND2X1_LOC_642/a_36_24# NAND2X1_LOC_642/Y 0.02fF
C7823 NAND2X1_LOC_72/Y NOR2X1_LOC_568/A 0.01fF
C7824 NOR2X1_LOC_42/a_36_216# INVX1_LOC_59/Y 0.00fF
C7825 VDD NAND2X1_LOC_212/Y 0.16fF
C7826 INVX1_LOC_206/Y INVX1_LOC_9/A 0.02fF
C7827 NAND2X1_LOC_740/Y NAND2X1_LOC_733/Y 0.05fF
C7828 INVX1_LOC_305/A NOR2X1_LOC_634/Y 0.04fF
C7829 INPUT_0 NOR2X1_LOC_743/Y 0.03fF
C7830 INVX1_LOC_126/A INVX1_LOC_46/A 0.03fF
C7831 NOR2X1_LOC_558/A INVX1_LOC_20/A 0.00fF
C7832 NOR2X1_LOC_67/A INVX1_LOC_4/A 0.07fF
C7833 INVX1_LOC_2/A INVX1_LOC_4/Y 0.18fF
C7834 INVX1_LOC_136/A NOR2X1_LOC_109/Y 0.10fF
C7835 NOR2X1_LOC_636/A INVX1_LOC_296/A 0.03fF
C7836 NOR2X1_LOC_818/Y INVX1_LOC_4/Y 0.01fF
C7837 NAND2X1_LOC_192/B INVX1_LOC_103/A 0.12fF
C7838 NAND2X1_LOC_55/a_36_24# NAND2X1_LOC_99/A 0.00fF
C7839 NAND2X1_LOC_357/B NOR2X1_LOC_301/A 0.07fF
C7840 INVX1_LOC_303/A NOR2X1_LOC_622/A 0.03fF
C7841 INVX1_LOC_226/Y INVX1_LOC_15/A 0.03fF
C7842 NOR2X1_LOC_197/A INVX1_LOC_1/A 0.05fF
C7843 VDD D_GATE_479 0.09fF
C7844 NAND2X1_LOC_738/B INVX1_LOC_209/Y 0.02fF
C7845 VDD D_INPUT_3 1.46fF
C7846 VDD INVX1_LOC_14/Y 2.09fF
C7847 INVX1_LOC_90/A NAND2X1_LOC_82/Y 0.07fF
C7848 INVX1_LOC_91/A INVX1_LOC_54/A 0.29fF
C7849 NOR2X1_LOC_111/A INVX1_LOC_46/A 0.07fF
C7850 INPUT_1 NAND2X1_LOC_81/B 0.03fF
C7851 NAND2X1_LOC_363/B NOR2X1_LOC_419/Y 0.10fF
C7852 NOR2X1_LOC_210/A NOR2X1_LOC_467/A 0.18fF
C7853 NAND2X1_LOC_72/Y INVX1_LOC_71/A 0.00fF
C7854 NAND2X1_LOC_724/A NAND2X1_LOC_711/Y 0.01fF
C7855 NAND2X1_LOC_787/A NOR2X1_LOC_716/B 0.12fF
C7856 INVX1_LOC_256/A NAND2X1_LOC_337/B 0.10fF
C7857 NOR2X1_LOC_391/A INVX1_LOC_3/Y 0.07fF
C7858 NAND2X1_LOC_303/Y INVX1_LOC_286/Y 0.09fF
C7859 INVX1_LOC_11/Y INVX1_LOC_54/A 0.07fF
C7860 NOR2X1_LOC_597/A INVX1_LOC_12/A 0.02fF
C7861 INVX1_LOC_10/A INVX1_LOC_15/A 1.39fF
C7862 NAND2X1_LOC_139/A NOR2X1_LOC_392/Y 0.02fF
C7863 INVX1_LOC_84/Y INVX1_LOC_175/A 0.01fF
C7864 NOR2X1_LOC_489/B NOR2X1_LOC_557/Y 0.10fF
C7865 NOR2X1_LOC_420/Y INVX1_LOC_314/Y 0.05fF
C7866 NOR2X1_LOC_405/A INVX1_LOC_92/A 0.16fF
C7867 INVX1_LOC_35/A NAND2X1_LOC_332/Y 0.03fF
C7868 VDD INVX1_LOC_230/A 0.17fF
C7869 NOR2X1_LOC_350/A INVX1_LOC_50/Y 0.05fF
C7870 INVX1_LOC_299/A NAND2X1_LOC_497/a_36_24# 0.00fF
C7871 NOR2X1_LOC_122/Y INVX1_LOC_290/Y 0.04fF
C7872 NAND2X1_LOC_9/Y INVX1_LOC_60/Y 0.10fF
C7873 NOR2X1_LOC_459/A INVX1_LOC_253/A 0.15fF
C7874 NOR2X1_LOC_751/A INVX1_LOC_125/A 0.03fF
C7875 NAND2X1_LOC_342/Y INVX1_LOC_23/A 0.01fF
C7876 NOR2X1_LOC_186/Y NAND2X1_LOC_283/a_36_24# 0.00fF
C7877 INVX1_LOC_95/Y NOR2X1_LOC_216/B 0.07fF
C7878 NOR2X1_LOC_815/Y NOR2X1_LOC_510/Y 0.03fF
C7879 INVX1_LOC_39/A NOR2X1_LOC_132/Y 0.01fF
C7880 INVX1_LOC_24/A INVX1_LOC_14/A 0.07fF
C7881 INVX1_LOC_36/A INVX1_LOC_211/A 0.08fF
C7882 INPUT_0 NOR2X1_LOC_178/a_36_216# 0.00fF
C7883 NOR2X1_LOC_468/Y INVX1_LOC_314/Y 0.15fF
C7884 INVX1_LOC_36/A NOR2X1_LOC_276/Y 0.04fF
C7885 INVX1_LOC_64/A INVX1_LOC_133/Y 0.15fF
C7886 INVX1_LOC_51/A NOR2X1_LOC_520/A 0.07fF
C7887 INVX1_LOC_40/Y INVX1_LOC_31/A 0.03fF
C7888 INVX1_LOC_45/A INVX1_LOC_61/Y 0.07fF
C7889 INVX1_LOC_276/A INVX1_LOC_64/A 0.00fF
C7890 NOR2X1_LOC_569/Y NOR2X1_LOC_383/B 0.01fF
C7891 INVX1_LOC_24/Y INVX1_LOC_77/A 0.20fF
C7892 NOR2X1_LOC_489/B INVX1_LOC_143/A 0.01fF
C7893 NOR2X1_LOC_679/Y NAND2X1_LOC_728/Y 0.11fF
C7894 NOR2X1_LOC_67/A INVX1_LOC_64/A 0.02fF
C7895 INVX1_LOC_130/A INVX1_LOC_72/A 0.04fF
C7896 NOR2X1_LOC_76/A NOR2X1_LOC_89/Y 0.02fF
C7897 NOR2X1_LOC_13/Y INVX1_LOC_161/Y 0.10fF
C7898 NAND2X1_LOC_308/B NAND2X1_LOC_175/Y 0.05fF
C7899 NOR2X1_LOC_298/Y INVX1_LOC_173/A 0.17fF
C7900 NAND2X1_LOC_456/Y NAND2X1_LOC_465/A 0.18fF
C7901 INVX1_LOC_279/A INVX1_LOC_271/A 0.12fF
C7902 INVX1_LOC_28/A INVX1_LOC_273/A -0.06fF
C7903 NAND2X1_LOC_703/Y NAND2X1_LOC_840/a_36_24# 0.00fF
C7904 INVX1_LOC_14/A NOR2X1_LOC_557/Y 0.17fF
C7905 NOR2X1_LOC_468/a_36_216# INVX1_LOC_57/A 0.00fF
C7906 NOR2X1_LOC_432/a_36_216# INVX1_LOC_27/A 0.01fF
C7907 INVX1_LOC_136/A INVX1_LOC_36/A 0.22fF
C7908 INVX1_LOC_235/Y NAND2X1_LOC_141/A 0.47fF
C7909 INVX1_LOC_52/Y NOR2X1_LOC_52/B 0.00fF
C7910 NOR2X1_LOC_208/Y NOR2X1_LOC_276/Y -0.00fF
C7911 INVX1_LOC_73/Y INVX1_LOC_33/A 0.01fF
C7912 NAND2X1_LOC_198/B NAND2X1_LOC_208/B 0.27fF
C7913 INVX1_LOC_65/A NAND2X1_LOC_63/Y 0.02fF
C7914 INVX1_LOC_200/Y INVX1_LOC_135/A 0.03fF
C7915 NOR2X1_LOC_272/Y NOR2X1_LOC_78/B 0.08fF
C7916 INVX1_LOC_136/A NOR2X1_LOC_267/A 0.94fF
C7917 NOR2X1_LOC_454/Y NOR2X1_LOC_207/A 0.03fF
C7918 NOR2X1_LOC_274/Y NOR2X1_LOC_590/A 0.00fF
C7919 INVX1_LOC_11/A INVX1_LOC_63/Y 0.12fF
C7920 NOR2X1_LOC_667/Y NOR2X1_LOC_152/Y 0.03fF
C7921 INVX1_LOC_50/A NOR2X1_LOC_749/Y 0.01fF
C7922 NOR2X1_LOC_791/B INVX1_LOC_72/A 0.00fF
C7923 NOR2X1_LOC_455/Y INVX1_LOC_227/A 0.01fF
C7924 INVX1_LOC_24/A NOR2X1_LOC_717/Y 0.03fF
C7925 NOR2X1_LOC_705/B INVX1_LOC_275/A 0.04fF
C7926 INVX1_LOC_106/Y NAND2X1_LOC_642/Y 0.02fF
C7927 NOR2X1_LOC_48/B INVX1_LOC_91/A 0.20fF
C7928 INVX1_LOC_37/Y INVX1_LOC_119/Y 0.07fF
C7929 INVX1_LOC_278/A INVX1_LOC_10/A 0.00fF
C7930 NOR2X1_LOC_456/a_36_216# NOR2X1_LOC_778/B 0.00fF
C7931 INVX1_LOC_223/A INVX1_LOC_94/A 0.75fF
C7932 NOR2X1_LOC_381/Y NOR2X1_LOC_84/Y 0.00fF
C7933 INVX1_LOC_17/A NAND2X1_LOC_357/B 0.07fF
C7934 NOR2X1_LOC_846/Y NOR2X1_LOC_516/B 0.01fF
C7935 INVX1_LOC_103/A NOR2X1_LOC_423/Y 0.03fF
C7936 NAND2X1_LOC_778/Y INVX1_LOC_16/A 0.02fF
C7937 INVX1_LOC_37/A NOR2X1_LOC_48/a_36_216# 0.00fF
C7938 NAND2X1_LOC_63/Y NAND2X1_LOC_267/B 0.00fF
C7939 INVX1_LOC_135/A INVX1_LOC_292/Y 0.19fF
C7940 INVX1_LOC_232/Y INVX1_LOC_1/A 0.91fF
C7941 INVX1_LOC_136/A NOR2X1_LOC_208/Y 0.03fF
C7942 INVX1_LOC_2/A NOR2X1_LOC_205/Y 0.16fF
C7943 INVX1_LOC_14/A INVX1_LOC_143/A 0.07fF
C7944 INVX1_LOC_199/Y NOR2X1_LOC_470/a_36_216# 0.00fF
C7945 INVX1_LOC_81/A INVX1_LOC_72/A 0.05fF
C7946 NOR2X1_LOC_446/A NOR2X1_LOC_348/B 0.02fF
C7947 NAND2X1_LOC_842/B INVX1_LOC_29/Y 0.07fF
C7948 INVX1_LOC_11/A NOR2X1_LOC_175/A 0.07fF
C7949 NAND2X1_LOC_741/B NOR2X1_LOC_577/Y 0.39fF
C7950 INVX1_LOC_174/Y NOR2X1_LOC_460/Y 0.01fF
C7951 VDD NOR2X1_LOC_831/Y 0.19fF
C7952 NAND2X1_LOC_364/A INVX1_LOC_184/A 0.04fF
C7953 NOR2X1_LOC_74/A INVX1_LOC_26/A 0.06fF
C7954 NOR2X1_LOC_778/B NAND2X1_LOC_190/Y 0.09fF
C7955 NOR2X1_LOC_598/B D_GATE_366 0.07fF
C7956 NOR2X1_LOC_716/B INVX1_LOC_30/A 0.20fF
C7957 INVX1_LOC_1/A INVX1_LOC_83/Y 0.02fF
C7958 NAND2X1_LOC_742/a_36_24# NAND2X1_LOC_863/B 0.01fF
C7959 INVX1_LOC_164/A INVX1_LOC_306/Y 0.02fF
C7960 VDD INVX1_LOC_167/A -0.00fF
C7961 INVX1_LOC_100/A INVX1_LOC_23/Y -0.04fF
C7962 NOR2X1_LOC_222/Y INVX1_LOC_103/A 1.42fF
C7963 NOR2X1_LOC_9/Y INVX1_LOC_26/A 0.55fF
C7964 INVX1_LOC_27/A INVX1_LOC_279/A 0.07fF
C7965 INVX1_LOC_255/Y NAND2X1_LOC_218/A 0.04fF
C7966 NOR2X1_LOC_15/Y INVX1_LOC_16/A 1.31fF
C7967 INVX1_LOC_255/Y NOR2X1_LOC_140/A 0.19fF
C7968 NOR2X1_LOC_508/a_36_216# NOR2X1_LOC_697/Y 0.00fF
C7969 INVX1_LOC_256/A NOR2X1_LOC_773/Y 0.01fF
C7970 INVX1_LOC_61/A NOR2X1_LOC_132/Y 0.02fF
C7971 NOR2X1_LOC_363/Y NOR2X1_LOC_755/Y -0.04fF
C7972 INVX1_LOC_67/Y INVX1_LOC_23/A 0.04fF
C7973 NOR2X1_LOC_565/A INVX1_LOC_104/A 0.04fF
C7974 NOR2X1_LOC_292/Y INVX1_LOC_57/A 0.01fF
C7975 INVX1_LOC_164/Y NOR2X1_LOC_160/B 0.00fF
C7976 INVX1_LOC_59/A INVX1_LOC_234/A 0.64fF
C7977 INVX1_LOC_36/A NOR2X1_LOC_278/A 0.03fF
C7978 INVX1_LOC_158/A NOR2X1_LOC_500/B 0.22fF
C7979 NOR2X1_LOC_559/B NOR2X1_LOC_350/A 0.01fF
C7980 INVX1_LOC_136/A NOR2X1_LOC_309/Y 4.22fF
C7981 NAND2X1_LOC_722/a_36_24# NAND2X1_LOC_722/A 0.00fF
C7982 INVX1_LOC_84/A INVX1_LOC_307/A 0.07fF
C7983 NAND2X1_LOC_574/a_36_24# INVX1_LOC_89/A 0.00fF
C7984 INVX1_LOC_118/Y INVX1_LOC_29/A 0.02fF
C7985 INVX1_LOC_178/Y INVX1_LOC_15/A 0.04fF
C7986 NOR2X1_LOC_446/A INVX1_LOC_22/A 0.01fF
C7987 INVX1_LOC_25/A NOR2X1_LOC_391/Y 0.03fF
C7988 NAND2X1_LOC_84/Y NOR2X1_LOC_557/Y 0.17fF
C7989 NOR2X1_LOC_68/A NOR2X1_LOC_154/a_36_216# 0.00fF
C7990 NAND2X1_LOC_81/B INVX1_LOC_118/A 0.08fF
C7991 NOR2X1_LOC_91/A INVX1_LOC_70/Y 0.06fF
C7992 NOR2X1_LOC_536/A INVX1_LOC_42/A 0.42fF
C7993 NAND2X1_LOC_778/Y INVX1_LOC_28/A 0.10fF
C7994 NOR2X1_LOC_640/Y INVX1_LOC_19/A 0.35fF
C7995 INVX1_LOC_114/A NAND2X1_LOC_220/B 0.10fF
C7996 INVX1_LOC_174/A INVX1_LOC_32/Y -0.03fF
C7997 INVX1_LOC_41/A INVX1_LOC_77/A 0.22fF
C7998 INVX1_LOC_14/A NOR2X1_LOC_130/A 0.15fF
C7999 INVX1_LOC_249/A NOR2X1_LOC_144/Y 0.04fF
C8000 NOR2X1_LOC_757/Y INVX1_LOC_30/A 0.19fF
C8001 NOR2X1_LOC_433/A INVX1_LOC_63/Y 1.51fF
C8002 INVX1_LOC_90/A NAND2X1_LOC_780/Y 0.01fF
C8003 INVX1_LOC_91/A NAND2X1_LOC_215/A 0.00fF
C8004 NOR2X1_LOC_791/B NAND2X1_LOC_338/B 0.03fF
C8005 INVX1_LOC_292/A INVX1_LOC_220/Y 0.01fF
C8006 NOR2X1_LOC_78/B NAND2X1_LOC_364/A 0.03fF
C8007 NOR2X1_LOC_717/B NOR2X1_LOC_457/A 0.06fF
C8008 NOR2X1_LOC_435/A NAND2X1_LOC_74/B 0.03fF
C8009 NOR2X1_LOC_655/Y NOR2X1_LOC_847/A 0.09fF
C8010 NOR2X1_LOC_160/B NOR2X1_LOC_719/B 0.01fF
C8011 INVX1_LOC_19/A NAND2X1_LOC_85/Y 0.00fF
C8012 INVX1_LOC_225/A NAND2X1_LOC_283/a_36_24# 0.01fF
C8013 NOR2X1_LOC_647/B NOR2X1_LOC_332/A 0.00fF
C8014 NOR2X1_LOC_15/Y INVX1_LOC_28/A 0.96fF
C8015 NOR2X1_LOC_500/A INVX1_LOC_196/A 0.10fF
C8016 INVX1_LOC_5/A INVX1_LOC_69/Y 0.07fF
C8017 INVX1_LOC_58/A INVX1_LOC_187/A 0.05fF
C8018 NOR2X1_LOC_32/B NOR2X1_LOC_45/B 0.11fF
C8019 NAND2X1_LOC_555/Y NOR2X1_LOC_128/B 0.14fF
C8020 NOR2X1_LOC_78/A NOR2X1_LOC_392/Y 0.01fF
C8021 NAND2X1_LOC_84/Y INVX1_LOC_143/A 0.02fF
C8022 NAND2X1_LOC_93/B INVX1_LOC_42/A 0.03fF
C8023 INVX1_LOC_208/A NOR2X1_LOC_457/B 0.10fF
C8024 NOR2X1_LOC_88/Y INVX1_LOC_12/A 1.69fF
C8025 NOR2X1_LOC_405/A INVX1_LOC_53/A 0.08fF
C8026 NOR2X1_LOC_52/B INVX1_LOC_63/Y 0.04fF
C8027 INVX1_LOC_312/Y NOR2X1_LOC_512/a_36_216# 0.00fF
C8028 INVX1_LOC_103/A NOR2X1_LOC_329/B 0.07fF
C8029 INVX1_LOC_78/A NOR2X1_LOC_536/A 0.10fF
C8030 NOR2X1_LOC_511/a_36_216# NOR2X1_LOC_577/Y 0.01fF
C8031 INVX1_LOC_41/A INVX1_LOC_124/A 0.04fF
C8032 NOR2X1_LOC_557/Y NOR2X1_LOC_612/B 0.04fF
C8033 INVX1_LOC_90/A NAND2X1_LOC_114/B 0.07fF
C8034 NOR2X1_LOC_405/a_36_216# INVX1_LOC_77/A 0.00fF
C8035 NOR2X1_LOC_717/B INVX1_LOC_30/A 0.03fF
C8036 NOR2X1_LOC_328/Y NOR2X1_LOC_637/Y 0.10fF
C8037 INVX1_LOC_12/A INVX1_LOC_84/A 0.21fF
C8038 INVX1_LOC_252/Y NOR2X1_LOC_19/B 0.03fF
C8039 INPUT_6 NAND2X1_LOC_1/Y 0.03fF
C8040 NAND2X1_LOC_756/a_36_24# INVX1_LOC_72/A 0.01fF
C8041 NOR2X1_LOC_589/A INVX1_LOC_181/Y 0.08fF
C8042 INVX1_LOC_307/A INVX1_LOC_15/A 0.46fF
C8043 NAND2X1_LOC_74/B INVX1_LOC_63/A 0.20fF
C8044 NOR2X1_LOC_649/B NOR2X1_LOC_847/A 0.04fF
C8045 NOR2X1_LOC_620/A NOR2X1_LOC_862/B 0.05fF
C8046 INVX1_LOC_35/A INVX1_LOC_59/Y 0.00fF
C8047 NOR2X1_LOC_570/B NOR2X1_LOC_352/Y 0.03fF
C8048 INVX1_LOC_192/A INVX1_LOC_192/Y 0.01fF
C8049 INVX1_LOC_90/A INVX1_LOC_141/Y 0.07fF
C8050 NAND2X1_LOC_207/Y INVX1_LOC_63/A 0.27fF
C8051 NOR2X1_LOC_809/B NOR2X1_LOC_801/B 0.16fF
C8052 INVX1_LOC_223/Y NOR2X1_LOC_78/A 0.03fF
C8053 NOR2X1_LOC_598/B INVX1_LOC_36/Y 0.04fF
C8054 NOR2X1_LOC_151/Y NOR2X1_LOC_457/A 0.00fF
C8055 NAND2X1_LOC_472/Y NOR2X1_LOC_383/B 0.14fF
C8056 INVX1_LOC_53/A NOR2X1_LOC_857/A 0.03fF
C8057 NAND2X1_LOC_364/A INVX1_LOC_83/A 0.07fF
C8058 INVX1_LOC_15/A NOR2X1_LOC_445/B 0.14fF
C8059 INVX1_LOC_3/A INVX1_LOC_42/A 0.45fF
C8060 NOR2X1_LOC_6/B INVX1_LOC_216/A 0.28fF
C8061 NOR2X1_LOC_65/B NOR2X1_LOC_536/A 0.68fF
C8062 INVX1_LOC_35/A INVX1_LOC_176/A 0.03fF
C8063 INVX1_LOC_21/A NOR2X1_LOC_139/Y 0.01fF
C8064 INVX1_LOC_90/A INVX1_LOC_312/Y 0.10fF
C8065 NAND2X1_LOC_787/A NAND2X1_LOC_633/Y 0.00fF
C8066 INVX1_LOC_21/A NAND2X1_LOC_655/A 0.06fF
C8067 NOR2X1_LOC_160/B INVX1_LOC_73/A 0.39fF
C8068 D_INPUT_0 NOR2X1_LOC_360/Y 0.03fF
C8069 INVX1_LOC_63/A NOR2X1_LOC_847/B -0.01fF
C8070 NOR2X1_LOC_826/Y VDD 0.23fF
C8071 NOR2X1_LOC_661/A INVX1_LOC_42/A 0.03fF
C8072 INVX1_LOC_34/A NOR2X1_LOC_219/Y 1.10fF
C8073 INVX1_LOC_78/A NAND2X1_LOC_93/B 0.03fF
C8074 NOR2X1_LOC_334/Y INVX1_LOC_179/A 0.01fF
C8075 NAND2X1_LOC_739/B NAND2X1_LOC_800/Y 0.01fF
C8076 INVX1_LOC_226/Y NAND2X1_LOC_464/Y 0.01fF
C8077 NAND2X1_LOC_139/A INVX1_LOC_25/Y 0.03fF
C8078 INVX1_LOC_143/A NOR2X1_LOC_612/B 0.20fF
C8079 INVX1_LOC_34/A INVX1_LOC_53/Y 0.03fF
C8080 INVX1_LOC_41/A NOR2X1_LOC_687/Y 0.05fF
C8081 INVX1_LOC_50/A NOR2X1_LOC_331/B 0.14fF
C8082 INVX1_LOC_45/A NAND2X1_LOC_652/Y 0.02fF
C8083 NAND2X1_LOC_323/B NOR2X1_LOC_802/A 0.07fF
C8084 NAND2X1_LOC_59/B GATE_662 0.10fF
C8085 INVX1_LOC_34/A NOR2X1_LOC_665/A 0.01fF
C8086 NAND2X1_LOC_466/a_36_24# NAND2X1_LOC_798/B 0.01fF
C8087 NOR2X1_LOC_577/Y NOR2X1_LOC_366/Y 0.00fF
C8088 NOR2X1_LOC_315/Y INVX1_LOC_56/Y 0.33fF
C8089 INVX1_LOC_48/Y NOR2X1_LOC_124/A 1.12fF
C8090 NOR2X1_LOC_151/Y INVX1_LOC_30/A 0.07fF
C8091 INVX1_LOC_90/A NOR2X1_LOC_546/B 0.03fF
C8092 NOR2X1_LOC_828/B NAND2X1_LOC_694/a_36_24# 0.00fF
C8093 NAND2X1_LOC_371/a_36_24# NOR2X1_LOC_356/A 0.00fF
C8094 NOR2X1_LOC_172/Y NAND2X1_LOC_656/Y 0.02fF
C8095 NOR2X1_LOC_65/B NAND2X1_LOC_93/B 0.04fF
C8096 NOR2X1_LOC_294/Y NAND2X1_LOC_348/A 0.02fF
C8097 NOR2X1_LOC_481/A INVX1_LOC_150/A 0.00fF
C8098 INVX1_LOC_47/A NOR2X1_LOC_303/Y 0.00fF
C8099 NOR2X1_LOC_778/B NOR2X1_LOC_220/A 0.03fF
C8100 INVX1_LOC_135/A NAND2X1_LOC_361/Y 0.24fF
C8101 INVX1_LOC_256/A NOR2X1_LOC_187/a_36_216# 0.12fF
C8102 INVX1_LOC_96/Y INVX1_LOC_16/A 0.14fF
C8103 INVX1_LOC_132/A INVX1_LOC_89/A 0.29fF
C8104 NOR2X1_LOC_272/Y INVX1_LOC_46/A 0.01fF
C8105 NOR2X1_LOC_226/A NAND2X1_LOC_862/A 0.01fF
C8106 NOR2X1_LOC_561/Y INVX1_LOC_104/A 0.10fF
C8107 NAND2X1_LOC_350/A INVX1_LOC_91/A 0.07fF
C8108 NAND2X1_LOC_214/Y INVX1_LOC_20/A 0.02fF
C8109 INVX1_LOC_32/A INVX1_LOC_272/A 0.01fF
C8110 INVX1_LOC_26/Y NAND2X1_LOC_85/Y 0.06fF
C8111 INVX1_LOC_194/A NAND2X1_LOC_462/B 0.09fF
C8112 NAND2X1_LOC_766/a_36_24# NOR2X1_LOC_770/Y 0.00fF
C8113 INVX1_LOC_77/A NOR2X1_LOC_122/Y 0.03fF
C8114 INVX1_LOC_90/A INVX1_LOC_275/A 0.41fF
C8115 NOR2X1_LOC_399/A NAND2X1_LOC_462/B 0.02fF
C8116 NOR2X1_LOC_783/A NOR2X1_LOC_708/A 0.10fF
C8117 INVX1_LOC_286/Y NOR2X1_LOC_536/a_36_216# 0.02fF
C8118 NOR2X1_LOC_473/B INVX1_LOC_155/A 0.01fF
C8119 INVX1_LOC_233/Y INVX1_LOC_118/A 0.03fF
C8120 NOR2X1_LOC_656/Y NOR2X1_LOC_660/Y 0.17fF
C8121 INVX1_LOC_12/A INVX1_LOC_15/A 0.28fF
C8122 NAND2X1_LOC_703/Y NOR2X1_LOC_111/A 0.07fF
C8123 NOR2X1_LOC_91/A INVX1_LOC_285/A 0.07fF
C8124 NAND2X1_LOC_503/a_36_24# NOR2X1_LOC_349/A 0.00fF
C8125 INVX1_LOC_280/Y NAND2X1_LOC_735/B 0.54fF
C8126 INVX1_LOC_88/A NOR2X1_LOC_173/a_36_216# 0.00fF
C8127 NOR2X1_LOC_778/B NOR2X1_LOC_548/Y 0.08fF
C8128 NOR2X1_LOC_266/a_36_216# INVX1_LOC_6/A -0.00fF
C8129 INVX1_LOC_225/A INVX1_LOC_89/A 0.07fF
C8130 NAND2X1_LOC_63/Y INVX1_LOC_4/Y 0.03fF
C8131 NOR2X1_LOC_441/Y INVX1_LOC_91/A 0.03fF
C8132 NOR2X1_LOC_91/A INVX1_LOC_265/Y 0.03fF
C8133 NAND2X1_LOC_303/Y VDD 1.52fF
C8134 INVX1_LOC_190/Y NAND2X1_LOC_466/Y 0.12fF
C8135 NAND2X1_LOC_787/A INVX1_LOC_71/Y 0.01fF
C8136 NAND2X1_LOC_198/B INPUT_0 0.01fF
C8137 INVX1_LOC_32/A NOR2X1_LOC_76/B 0.10fF
C8138 INVX1_LOC_57/A NOR2X1_LOC_461/B 0.00fF
C8139 INVX1_LOC_55/Y NOR2X1_LOC_770/B 0.11fF
C8140 NOR2X1_LOC_65/B INVX1_LOC_3/A 1.91fF
C8141 NOR2X1_LOC_329/B INVX1_LOC_67/A 0.01fF
C8142 NAND2X1_LOC_303/Y NAND2X1_LOC_800/A 0.02fF
C8143 INVX1_LOC_82/A INPUT_1 0.26fF
C8144 NOR2X1_LOC_243/Y INVX1_LOC_89/A 0.02fF
C8145 NAND2X1_LOC_333/a_36_24# NOR2X1_LOC_331/B 0.01fF
C8146 INVX1_LOC_232/A INVX1_LOC_22/A 0.12fF
C8147 NOR2X1_LOC_389/A NOR2X1_LOC_657/B 0.03fF
C8148 NOR2X1_LOC_742/A NOR2X1_LOC_550/B 0.10fF
C8149 INVX1_LOC_7/Y INVX1_LOC_9/A 0.00fF
C8150 NOR2X1_LOC_553/Y NOR2X1_LOC_570/Y 0.07fF
C8151 NAND2X1_LOC_550/A NAND2X1_LOC_241/Y 0.01fF
C8152 NAND2X1_LOC_175/Y INVX1_LOC_272/A 0.01fF
C8153 NOR2X1_LOC_373/Y NAND2X1_LOC_374/Y 0.09fF
C8154 NOR2X1_LOC_753/Y INVX1_LOC_282/A 0.04fF
C8155 NAND2X1_LOC_717/Y NOR2X1_LOC_576/B 2.22fF
C8156 INVX1_LOC_23/A INVX1_LOC_285/A 0.07fF
C8157 INVX1_LOC_174/A INVX1_LOC_115/A 0.67fF
C8158 NOR2X1_LOC_209/Y INVX1_LOC_89/A 0.07fF
C8159 INVX1_LOC_269/A INVX1_LOC_117/A 0.07fF
C8160 INVX1_LOC_24/A INVX1_LOC_48/A 0.02fF
C8161 NAND2X1_LOC_342/Y INVX1_LOC_313/A 0.22fF
C8162 D_GATE_366 NOR2X1_LOC_156/B 0.04fF
C8163 NOR2X1_LOC_15/Y NAND2X1_LOC_236/a_36_24# 0.00fF
C8164 INVX1_LOC_23/A NOR2X1_LOC_814/A 0.01fF
C8165 NOR2X1_LOC_383/B NAND2X1_LOC_773/B 0.03fF
C8166 NOR2X1_LOC_237/a_36_216# INVX1_LOC_6/A 0.00fF
C8167 INVX1_LOC_62/Y NOR2X1_LOC_557/A 0.09fF
C8168 NOR2X1_LOC_742/A INVX1_LOC_249/Y 0.01fF
C8169 NOR2X1_LOC_65/Y NAND2X1_LOC_74/B 0.04fF
C8170 NOR2X1_LOC_703/Y NOR2X1_LOC_374/A 0.12fF
C8171 NOR2X1_LOC_274/B NAND2X1_LOC_447/Y 0.19fF
C8172 INVX1_LOC_34/A NOR2X1_LOC_113/B 0.03fF
C8173 NOR2X1_LOC_576/B INVX1_LOC_16/A 0.05fF
C8174 NOR2X1_LOC_447/Y NOR2X1_LOC_45/B 0.03fF
C8175 NOR2X1_LOC_660/Y INVX1_LOC_63/A 0.11fF
C8176 INVX1_LOC_150/Y INVX1_LOC_66/Y 0.02fF
C8177 NOR2X1_LOC_264/Y INVX1_LOC_92/Y 0.06fF
C8178 INVX1_LOC_30/A NAND2X1_LOC_633/Y 0.10fF
C8179 INVX1_LOC_28/A NAND2X1_LOC_840/B 0.13fF
C8180 INVX1_LOC_128/A INVX1_LOC_128/Y 0.09fF
C8181 NOR2X1_LOC_147/B INVX1_LOC_78/Y 0.03fF
C8182 INVX1_LOC_149/A NOR2X1_LOC_74/A 0.46fF
C8183 NAND2X1_LOC_114/B INVX1_LOC_38/A 0.07fF
C8184 NAND2X1_LOC_218/B INVX1_LOC_74/Y 0.00fF
C8185 NOR2X1_LOC_316/Y NOR2X1_LOC_83/Y 0.05fF
C8186 NOR2X1_LOC_592/A INVX1_LOC_54/A 0.01fF
C8187 NOR2X1_LOC_261/Y INVX1_LOC_12/A 0.20fF
C8188 INVX1_LOC_95/Y NOR2X1_LOC_303/Y 0.02fF
C8189 NAND2X1_LOC_837/Y NOR2X1_LOC_670/a_36_216# 0.01fF
C8190 NAND2X1_LOC_364/A INVX1_LOC_46/A 0.09fF
C8191 INVX1_LOC_217/A NOR2X1_LOC_482/a_36_216# 0.01fF
C8192 NOR2X1_LOC_67/A INVX1_LOC_282/A 0.09fF
C8193 NOR2X1_LOC_142/Y INVX1_LOC_91/A 0.10fF
C8194 NOR2X1_LOC_215/Y INVX1_LOC_76/A 0.03fF
C8195 INVX1_LOC_296/A NAND2X1_LOC_430/B 0.05fF
C8196 INVX1_LOC_208/A INVX1_LOC_73/A 0.02fF
C8197 NOR2X1_LOC_273/Y INVX1_LOC_139/A 0.04fF
C8198 INVX1_LOC_299/A NOR2X1_LOC_831/B 0.02fF
C8199 NOR2X1_LOC_296/Y NOR2X1_LOC_99/Y 0.06fF
C8200 INVX1_LOC_53/A INVX1_LOC_109/Y 0.04fF
C8201 NOR2X1_LOC_860/B NOR2X1_LOC_35/Y 0.10fF
C8202 INVX1_LOC_72/A NOR2X1_LOC_363/Y 0.05fF
C8203 INVX1_LOC_141/Y INVX1_LOC_38/A 0.04fF
C8204 INVX1_LOC_176/Y NOR2X1_LOC_78/A 0.11fF
C8205 NOR2X1_LOC_577/Y NAND2X1_LOC_447/Y 0.10fF
C8206 INVX1_LOC_43/Y NAND2X1_LOC_268/a_36_24# 0.00fF
C8207 INVX1_LOC_49/A INVX1_LOC_115/Y 0.01fF
C8208 NAND2X1_LOC_351/A NAND2X1_LOC_96/A 0.07fF
C8209 NOR2X1_LOC_624/A INVX1_LOC_65/A 0.03fF
C8210 INVX1_LOC_18/A INVX1_LOC_33/Y 0.03fF
C8211 NOR2X1_LOC_294/Y INVX1_LOC_38/A 0.00fF
C8212 INVX1_LOC_63/Y INVX1_LOC_199/A 0.01fF
C8213 NOR2X1_LOC_106/Y VDD 0.14fF
C8214 INVX1_LOC_200/A NOR2X1_LOC_88/Y 0.12fF
C8215 NAND2X1_LOC_348/A NOR2X1_LOC_789/A 0.00fF
C8216 NAND2X1_LOC_755/a_36_24# NOR2X1_LOC_78/A 0.00fF
C8217 INVX1_LOC_254/A VDD 0.12fF
C8218 NOR2X1_LOC_349/B INVX1_LOC_156/A 0.03fF
C8219 INPUT_0 INVX1_LOC_53/Y 0.07fF
C8220 NAND2X1_LOC_725/A INVX1_LOC_102/A 0.19fF
C8221 NAND2X1_LOC_466/Y NOR2X1_LOC_56/Y 0.05fF
C8222 INVX1_LOC_5/A NOR2X1_LOC_89/A 0.07fF
C8223 NOR2X1_LOC_75/Y INVX1_LOC_113/A 0.01fF
C8224 INVX1_LOC_39/A NAND2X1_LOC_81/B 0.02fF
C8225 NOR2X1_LOC_655/B INVX1_LOC_91/A 0.10fF
C8226 NOR2X1_LOC_282/Y NOR2X1_LOC_301/A 0.01fF
C8227 D_INPUT_0 NOR2X1_LOC_567/B 0.07fF
C8228 NOR2X1_LOC_84/Y NOR2X1_LOC_124/A 0.07fF
C8229 INVX1_LOC_161/Y NOR2X1_LOC_697/Y 0.02fF
C8230 NOR2X1_LOC_348/B NAND2X1_LOC_447/Y 0.17fF
C8231 INVX1_LOC_214/A NAND2X1_LOC_655/A 0.17fF
C8232 NOR2X1_LOC_689/a_36_216# NAND2X1_LOC_175/Y 0.01fF
C8233 INVX1_LOC_200/A INVX1_LOC_84/A 1.51fF
C8234 NOR2X1_LOC_690/A VDD 2.04fF
C8235 NOR2X1_LOC_730/Y NOR2X1_LOC_730/B 0.04fF
C8236 INVX1_LOC_178/A NOR2X1_LOC_89/A 0.10fF
C8237 NOR2X1_LOC_554/B NOR2X1_LOC_655/Y 0.11fF
C8238 NOR2X1_LOC_78/B NOR2X1_LOC_405/A 0.10fF
C8239 INVX1_LOC_54/Y INVX1_LOC_95/Y 0.00fF
C8240 NAND2X1_LOC_466/Y VDD 0.00fF
C8241 NOR2X1_LOC_413/Y VDD 0.92fF
C8242 NOR2X1_LOC_152/Y NOR2X1_LOC_536/A 0.02fF
C8243 NOR2X1_LOC_91/Y NOR2X1_LOC_177/a_36_216# 0.00fF
C8244 NOR2X1_LOC_68/A NOR2X1_LOC_61/Y 0.17fF
C8245 NOR2X1_LOC_496/Y NAND2X1_LOC_254/Y 0.04fF
C8246 NOR2X1_LOC_78/A INVX1_LOC_25/Y 0.17fF
C8247 INVX1_LOC_136/A NOR2X1_LOC_435/A 0.01fF
C8248 INVX1_LOC_164/A NOR2X1_LOC_9/Y 0.19fF
C8249 NOR2X1_LOC_194/Y VDD 0.24fF
C8250 INVX1_LOC_121/Y INVX1_LOC_14/Y 0.01fF
C8251 INVX1_LOC_313/A INVX1_LOC_67/Y 0.30fF
C8252 NOR2X1_LOC_693/Y NAND2X1_LOC_464/B 0.00fF
C8253 INVX1_LOC_31/A INVX1_LOC_285/A 0.07fF
C8254 NAND2X1_LOC_454/Y NOR2X1_LOC_678/A 0.07fF
C8255 INVX1_LOC_50/A NOR2X1_LOC_106/a_36_216# 0.00fF
C8256 NAND2X1_LOC_214/B NOR2X1_LOC_38/B 0.10fF
C8257 NAND2X1_LOC_58/a_36_24# NOR2X1_LOC_861/Y 0.07fF
C8258 NOR2X1_LOC_360/Y INVX1_LOC_46/Y 0.07fF
C8259 INVX1_LOC_31/A NOR2X1_LOC_814/A 0.10fF
C8260 INVX1_LOC_177/A INVX1_LOC_14/Y 0.01fF
C8261 NOR2X1_LOC_93/Y INVX1_LOC_3/Y 0.03fF
C8262 INVX1_LOC_2/Y NOR2X1_LOC_537/Y 0.03fF
C8263 NAND2X1_LOC_463/B INVX1_LOC_169/A 0.01fF
C8264 NOR2X1_LOC_634/B NOR2X1_LOC_857/A 0.03fF
C8265 INPUT_0 NOR2X1_LOC_76/a_36_216# 0.00fF
C8266 INVX1_LOC_21/A NOR2X1_LOC_685/Y 0.05fF
C8267 NOR2X1_LOC_637/A NAND2X1_LOC_798/B 0.04fF
C8268 NOR2X1_LOC_34/A INVX1_LOC_15/A 0.01fF
C8269 NOR2X1_LOC_78/B NOR2X1_LOC_857/A 0.03fF
C8270 NOR2X1_LOC_168/Y NOR2X1_LOC_445/B 0.02fF
C8271 INVX1_LOC_41/A INVX1_LOC_9/A 0.11fF
C8272 NOR2X1_LOC_468/Y INVX1_LOC_170/Y 0.00fF
C8273 NOR2X1_LOC_121/A INVX1_LOC_59/Y 0.00fF
C8274 INVX1_LOC_22/A NAND2X1_LOC_447/Y 0.10fF
C8275 INVX1_LOC_27/A NOR2X1_LOC_38/B 0.07fF
C8276 NOR2X1_LOC_502/Y NOR2X1_LOC_340/A 0.03fF
C8277 NAND2X1_LOC_174/a_36_24# NOR2X1_LOC_331/B 0.01fF
C8278 NAND2X1_LOC_535/a_36_24# INVX1_LOC_49/Y 0.00fF
C8279 INVX1_LOC_39/A INVX1_LOC_4/Y 0.03fF
C8280 INVX1_LOC_219/Y INVX1_LOC_280/A 0.03fF
C8281 INVX1_LOC_300/Y NAND2X1_LOC_770/Y 0.65fF
C8282 NOR2X1_LOC_554/B NOR2X1_LOC_649/B 1.06fF
C8283 INVX1_LOC_18/A INVX1_LOC_220/A 0.09fF
C8284 INVX1_LOC_25/Y NAND2X1_LOC_464/A 0.02fF
C8285 INVX1_LOC_72/A NOR2X1_LOC_485/Y 0.01fF
C8286 NOR2X1_LOC_99/B INVX1_LOC_91/A 0.09fF
C8287 NOR2X1_LOC_414/Y NOR2X1_LOC_416/A 0.33fF
C8288 NAND2X1_LOC_337/B NOR2X1_LOC_89/A 0.01fF
C8289 NOR2X1_LOC_554/B INVX1_LOC_3/A 0.07fF
C8290 INVX1_LOC_113/Y NAND2X1_LOC_93/B 0.03fF
C8291 INVX1_LOC_83/A NOR2X1_LOC_349/A 0.30fF
C8292 INVX1_LOC_272/Y NOR2X1_LOC_677/a_36_216# 0.00fF
C8293 NOR2X1_LOC_816/A NOR2X1_LOC_89/A 0.06fF
C8294 INVX1_LOC_217/A INVX1_LOC_84/A 0.05fF
C8295 NOR2X1_LOC_13/Y NOR2X1_LOC_841/A 0.10fF
C8296 INVX1_LOC_256/A INVX1_LOC_42/A 0.07fF
C8297 NOR2X1_LOC_647/B NOR2X1_LOC_847/A 0.04fF
C8298 INVX1_LOC_269/A INVX1_LOC_3/Y 0.13fF
C8299 INVX1_LOC_136/A INVX1_LOC_63/A 0.23fF
C8300 NOR2X1_LOC_232/Y INVX1_LOC_3/Y 0.08fF
C8301 NOR2X1_LOC_426/Y NOR2X1_LOC_11/Y 0.26fF
C8302 NOR2X1_LOC_554/B NOR2X1_LOC_814/a_36_216# 0.00fF
C8303 NAND2X1_LOC_513/B INVX1_LOC_271/Y 0.01fF
C8304 NAND2X1_LOC_854/B INVX1_LOC_76/A 1.02fF
C8305 INVX1_LOC_89/A NAND2X1_LOC_642/Y 0.76fF
C8306 INVX1_LOC_111/A NOR2X1_LOC_814/A 0.10fF
C8307 NAND2X1_LOC_30/Y D_INPUT_5 0.37fF
C8308 INVX1_LOC_208/A NOR2X1_LOC_122/a_36_216# 0.01fF
C8309 NOR2X1_LOC_53/a_36_216# INVX1_LOC_20/A 0.00fF
C8310 NAND2X1_LOC_759/a_36_24# NOR2X1_LOC_743/Y 0.01fF
C8311 INVX1_LOC_182/A INVX1_LOC_91/A 0.07fF
C8312 NOR2X1_LOC_606/Y INVX1_LOC_42/A 0.00fF
C8313 NOR2X1_LOC_718/B INVX1_LOC_179/A 0.02fF
C8314 NAND2X1_LOC_508/a_36_24# NOR2X1_LOC_340/A 0.00fF
C8315 NAND2X1_LOC_859/B NOR2X1_LOC_536/A 0.01fF
C8316 INVX1_LOC_83/A NOR2X1_LOC_857/A 0.07fF
C8317 NOR2X1_LOC_526/Y INVX1_LOC_118/A 0.04fF
C8318 INVX1_LOC_75/A INVX1_LOC_98/A 0.07fF
C8319 INVX1_LOC_304/Y NOR2X1_LOC_88/Y 0.07fF
C8320 INVX1_LOC_75/A NOR2X1_LOC_78/A 0.16fF
C8321 NOR2X1_LOC_41/Y INVX1_LOC_117/Y 0.01fF
C8322 NOR2X1_LOC_211/A INVX1_LOC_9/A 0.01fF
C8323 INVX1_LOC_89/A D_GATE_662 0.01fF
C8324 NOR2X1_LOC_106/Y INVX1_LOC_133/A 0.01fF
C8325 NOR2X1_LOC_315/Y NOR2X1_LOC_179/a_36_216# 0.01fF
C8326 INVX1_LOC_256/A INVX1_LOC_78/A 0.08fF
C8327 D_INPUT_1 NAND2X1_LOC_474/Y 0.07fF
C8328 NAND2X1_LOC_858/B NOR2X1_LOC_528/Y 0.15fF
C8329 INVX1_LOC_225/Y NAND2X1_LOC_72/B 0.10fF
C8330 INVX1_LOC_144/Y NOR2X1_LOC_510/B 0.00fF
C8331 NOR2X1_LOC_307/A NOR2X1_LOC_307/Y 0.05fF
C8332 NAND2X1_LOC_9/Y NOR2X1_LOC_272/Y 0.05fF
C8333 NOR2X1_LOC_272/Y INVX1_LOC_233/A 0.10fF
C8334 INVX1_LOC_304/Y INVX1_LOC_84/A 0.02fF
C8335 NAND2X1_LOC_656/Y INVX1_LOC_38/A 0.17fF
C8336 INVX1_LOC_244/Y NOR2X1_LOC_48/B 0.03fF
C8337 NOR2X1_LOC_329/B NOR2X1_LOC_137/Y 0.61fF
C8338 INVX1_LOC_256/A NOR2X1_LOC_65/B 0.01fF
C8339 INVX1_LOC_58/A INVX1_LOC_269/A 0.10fF
C8340 NOR2X1_LOC_848/Y NOR2X1_LOC_105/Y 0.21fF
C8341 INVX1_LOC_58/A NOR2X1_LOC_232/Y 0.00fF
C8342 NOR2X1_LOC_773/Y INVX1_LOC_297/A 0.03fF
C8343 INPUT_0 NAND2X1_LOC_465/A 0.00fF
C8344 NOR2X1_LOC_91/A NOR2X1_LOC_590/A 0.03fF
C8345 NOR2X1_LOC_264/Y INVX1_LOC_106/A -0.00fF
C8346 NOR2X1_LOC_730/Y NOR2X1_LOC_155/A 0.01fF
C8347 NAND2X1_LOC_537/Y NAND2X1_LOC_590/a_36_24# 0.00fF
C8348 INVX1_LOC_181/Y INVX1_LOC_4/A -0.00fF
C8349 INVX1_LOC_21/A INVX1_LOC_13/Y 0.03fF
C8350 NAND2X1_LOC_222/A NAND2X1_LOC_555/Y 0.02fF
C8351 NOR2X1_LOC_201/A NOR2X1_LOC_590/A 0.01fF
C8352 INVX1_LOC_124/Y INVX1_LOC_26/A 0.35fF
C8353 NAND2X1_LOC_87/a_36_24# NOR2X1_LOC_92/Y 0.01fF
C8354 NAND2X1_LOC_474/Y NOR2X1_LOC_652/Y 0.07fF
C8355 NAND2X1_LOC_803/B INVX1_LOC_23/A 0.02fF
C8356 NOR2X1_LOC_377/Y NOR2X1_LOC_89/A 0.00fF
C8357 NOR2X1_LOC_6/B NOR2X1_LOC_641/a_36_216# 0.02fF
C8358 INVX1_LOC_35/A INVX1_LOC_103/A 0.07fF
C8359 INVX1_LOC_49/A D_INPUT_5 0.07fF
C8360 NOR2X1_LOC_389/A INVX1_LOC_271/A 0.01fF
C8361 INVX1_LOC_45/Y NOR2X1_LOC_334/Y 0.07fF
C8362 INVX1_LOC_206/Y INVX1_LOC_76/A 0.07fF
C8363 NAND2X1_LOC_652/Y NOR2X1_LOC_331/B 0.03fF
C8364 INVX1_LOC_11/A NOR2X1_LOC_435/a_36_216# 0.02fF
C8365 NOR2X1_LOC_590/A INVX1_LOC_23/A 0.43fF
C8366 INVX1_LOC_196/Y INVX1_LOC_274/A 0.20fF
C8367 INVX1_LOC_13/A NOR2X1_LOC_673/A 0.01fF
C8368 NAND2X1_LOC_222/B INVX1_LOC_5/A 0.00fF
C8369 INVX1_LOC_1/A INVX1_LOC_50/Y 0.13fF
C8370 NAND2X1_LOC_808/A NOR2X1_LOC_88/Y 0.07fF
C8371 INVX1_LOC_66/A NOR2X1_LOC_831/B 0.01fF
C8372 INVX1_LOC_224/A INVX1_LOC_5/A 0.03fF
C8373 NOR2X1_LOC_15/Y NAND2X1_LOC_794/B 0.14fF
C8374 NOR2X1_LOC_303/Y INVX1_LOC_271/Y 0.07fF
C8375 NOR2X1_LOC_100/A NAND2X1_LOC_206/B 0.36fF
C8376 NOR2X1_LOC_152/Y NAND2X1_LOC_470/B 2.68fF
C8377 INVX1_LOC_27/A NOR2X1_LOC_468/Y 0.46fF
C8378 INVX1_LOC_17/A NOR2X1_LOC_291/Y 0.13fF
C8379 INVX1_LOC_11/A INVX1_LOC_5/A 0.20fF
C8380 INVX1_LOC_18/A NOR2X1_LOC_686/a_36_216# 0.00fF
C8381 INVX1_LOC_62/A NAND2X1_LOC_85/Y 0.05fF
C8382 NOR2X1_LOC_644/A NOR2X1_LOC_830/a_36_216# 0.00fF
C8383 INVX1_LOC_25/A NOR2X1_LOC_248/Y 0.05fF
C8384 INVX1_LOC_289/Y NAND2X1_LOC_714/B 0.41fF
C8385 INVX1_LOC_21/A INVX1_LOC_88/A 0.16fF
C8386 NOR2X1_LOC_78/B INVX1_LOC_109/Y 0.07fF
C8387 NOR2X1_LOC_172/Y INVX1_LOC_128/Y 0.09fF
C8388 NOR2X1_LOC_657/B NAND2X1_LOC_469/B 0.02fF
C8389 INVX1_LOC_41/A INVX1_LOC_274/Y 0.10fF
C8390 NOR2X1_LOC_773/Y NOR2X1_LOC_89/A 0.15fF
C8391 INVX1_LOC_224/Y NOR2X1_LOC_791/B 0.23fF
C8392 INVX1_LOC_72/A INVX1_LOC_29/Y 0.03fF
C8393 NOR2X1_LOC_664/Y NOR2X1_LOC_38/B 0.23fF
C8394 NOR2X1_LOC_61/B NOR2X1_LOC_523/A 0.04fF
C8395 NAND2X1_LOC_808/A INVX1_LOC_84/A 0.09fF
C8396 NOR2X1_LOC_113/A INVX1_LOC_46/A 0.01fF
C8397 NOR2X1_LOC_405/A INVX1_LOC_46/A 0.25fF
C8398 INVX1_LOC_11/A INVX1_LOC_178/A 0.01fF
C8399 NOR2X1_LOC_794/B INVX1_LOC_50/Y 0.03fF
C8400 INVX1_LOC_24/A NOR2X1_LOC_383/B 0.06fF
C8401 NOR2X1_LOC_254/Y INVX1_LOC_271/Y 0.07fF
C8402 NAND2X1_LOC_652/Y NOR2X1_LOC_592/B 0.02fF
C8403 INVX1_LOC_316/A D_INPUT_3 0.01fF
C8404 NOR2X1_LOC_381/Y INVX1_LOC_1/A 0.06fF
C8405 INVX1_LOC_78/Y INVX1_LOC_38/A 0.01fF
C8406 NOR2X1_LOC_616/Y INVX1_LOC_3/Y 0.10fF
C8407 INVX1_LOC_278/A INVX1_LOC_217/A 0.17fF
C8408 NOR2X1_LOC_596/A INVX1_LOC_105/Y 0.05fF
C8409 NOR2X1_LOC_817/Y NOR2X1_LOC_140/A 0.07fF
C8410 NOR2X1_LOC_68/A NOR2X1_LOC_678/A 0.03fF
C8411 INVX1_LOC_91/A NAND2X1_LOC_61/a_36_24# 0.01fF
C8412 NAND2X1_LOC_807/Y INVX1_LOC_285/A 0.03fF
C8413 INVX1_LOC_27/A NOR2X1_LOC_389/A 4.21fF
C8414 NOR2X1_LOC_824/A NAND2X1_LOC_546/a_36_24# 0.01fF
C8415 NOR2X1_LOC_335/B INVX1_LOC_92/A 0.20fF
C8416 NAND2X1_LOC_807/Y INVX1_LOC_265/Y 0.01fF
C8417 NOR2X1_LOC_91/A NAND2X1_LOC_354/B 0.03fF
C8418 INVX1_LOC_28/A NAND2X1_LOC_456/Y 0.08fF
C8419 NOR2X1_LOC_557/Y NOR2X1_LOC_383/B 0.07fF
C8420 INVX1_LOC_89/A NOR2X1_LOC_48/Y 0.03fF
C8421 NOR2X1_LOC_798/A NOR2X1_LOC_336/B 0.00fF
C8422 NAND2X1_LOC_655/a_36_24# INVX1_LOC_94/Y 0.00fF
C8423 NOR2X1_LOC_147/B NOR2X1_LOC_727/B 0.03fF
C8424 INVX1_LOC_6/A NOR2X1_LOC_364/A 0.02fF
C8425 INVX1_LOC_50/A NOR2X1_LOC_388/Y 0.03fF
C8426 NOR2X1_LOC_168/B INVX1_LOC_18/Y 0.01fF
C8427 NAND2X1_LOC_276/Y NAND2X1_LOC_215/A 0.07fF
C8428 INVX1_LOC_236/Y NAND2X1_LOC_326/A 0.12fF
C8429 INVX1_LOC_65/Y INVX1_LOC_29/A 0.03fF
C8430 NOR2X1_LOC_709/A INVX1_LOC_16/Y 0.02fF
C8431 NOR2X1_LOC_798/A NAND2X1_LOC_364/A 0.09fF
C8432 NOR2X1_LOC_208/Y NOR2X1_LOC_665/Y 0.03fF
C8433 INVX1_LOC_11/A NAND2X1_LOC_337/B 0.96fF
C8434 INVX1_LOC_224/Y NOR2X1_LOC_124/B 0.02fF
C8435 NOR2X1_LOC_730/A INVX1_LOC_15/A 0.03fF
C8436 INVX1_LOC_34/Y INVX1_LOC_23/Y 0.04fF
C8437 INVX1_LOC_11/A NOR2X1_LOC_816/A 0.04fF
C8438 NAND2X1_LOC_350/A NOR2X1_LOC_592/A -0.02fF
C8439 INVX1_LOC_28/A INVX1_LOC_49/Y 0.47fF
C8440 INVX1_LOC_58/A NAND2X1_LOC_137/a_36_24# 0.00fF
C8441 NOR2X1_LOC_445/Y INVX1_LOC_53/A 0.01fF
C8442 INVX1_LOC_286/Y INVX1_LOC_14/A -0.01fF
C8443 INVX1_LOC_25/A NOR2X1_LOC_6/B 0.06fF
C8444 INVX1_LOC_6/A INVX1_LOC_285/A 0.00fF
C8445 INVX1_LOC_27/A INVX1_LOC_62/Y 0.00fF
C8446 NOR2X1_LOC_168/B NAND2X1_LOC_279/a_36_24# 0.00fF
C8447 NOR2X1_LOC_442/a_36_216# INVX1_LOC_30/A 0.00fF
C8448 NOR2X1_LOC_598/B INVX1_LOC_149/Y 0.00fF
C8449 INVX1_LOC_5/A NOR2X1_LOC_433/A 0.07fF
C8450 INVX1_LOC_21/A NOR2X1_LOC_758/a_36_216# 0.00fF
C8451 NOR2X1_LOC_297/a_36_216# NOR2X1_LOC_392/Y 0.01fF
C8452 NOR2X1_LOC_392/B NOR2X1_LOC_717/A 0.10fF
C8453 INVX1_LOC_234/A NOR2X1_LOC_38/B 0.01fF
C8454 INVX1_LOC_27/A NOR2X1_LOC_596/A 0.11fF
C8455 INVX1_LOC_143/A NOR2X1_LOC_383/B 0.07fF
C8456 NAND2X1_LOC_72/Y NOR2X1_LOC_388/Y 0.00fF
C8457 NOR2X1_LOC_455/Y INVX1_LOC_104/A 0.03fF
C8458 NAND2X1_LOC_573/Y NOR2X1_LOC_744/a_36_216# 0.00fF
C8459 INVX1_LOC_140/A NOR2X1_LOC_89/A 0.12fF
C8460 INVX1_LOC_5/A NOR2X1_LOC_593/Y 0.02fF
C8461 INVX1_LOC_17/A INVX1_LOC_110/A 0.00fF
C8462 INVX1_LOC_144/Y INVX1_LOC_57/A 0.03fF
C8463 INVX1_LOC_304/Y INVX1_LOC_278/A 0.07fF
C8464 INVX1_LOC_21/A INVX1_LOC_303/A 0.07fF
C8465 INVX1_LOC_56/Y NAND2X1_LOC_99/A 0.01fF
C8466 NAND2X1_LOC_363/B NAND2X1_LOC_114/a_36_24# 0.00fF
C8467 INVX1_LOC_178/A NOR2X1_LOC_433/A 0.05fF
C8468 NOR2X1_LOC_590/A INVX1_LOC_31/A 6.27fF
C8469 INVX1_LOC_233/A NAND2X1_LOC_785/A 0.08fF
C8470 INVX1_LOC_157/A INVX1_LOC_78/A 0.03fF
C8471 NOR2X1_LOC_795/Y INVX1_LOC_292/Y 0.31fF
C8472 INVX1_LOC_178/A NOR2X1_LOC_474/A 0.03fF
C8473 INVX1_LOC_22/Y INVX1_LOC_31/A 0.13fF
C8474 NOR2X1_LOC_156/A NOR2X1_LOC_467/A 0.04fF
C8475 INVX1_LOC_5/A NOR2X1_LOC_52/B 0.20fF
C8476 INVX1_LOC_64/A NAND2X1_LOC_35/a_36_24# 0.00fF
C8477 INVX1_LOC_50/A NAND2X1_LOC_479/Y 0.03fF
C8478 NOR2X1_LOC_647/B NOR2X1_LOC_554/B -0.02fF
C8479 NOR2X1_LOC_849/a_36_216# NOR2X1_LOC_590/A 0.00fF
C8480 NOR2X1_LOC_65/B NOR2X1_LOC_440/Y -0.00fF
C8481 INVX1_LOC_226/Y D_INPUT_1 0.33fF
C8482 NOR2X1_LOC_67/A NAND2X1_LOC_624/B 0.02fF
C8483 INVX1_LOC_55/A NOR2X1_LOC_68/A 0.01fF
C8484 NAND2X1_LOC_149/Y INVX1_LOC_34/A 0.08fF
C8485 NOR2X1_LOC_644/A NOR2X1_LOC_334/Y 0.05fF
C8486 D_INPUT_0 INVX1_LOC_26/A 0.56fF
C8487 NOR2X1_LOC_19/B NOR2X1_LOC_38/B 0.19fF
C8488 INVX1_LOC_27/A NOR2X1_LOC_844/A 0.03fF
C8489 INVX1_LOC_1/A NOR2X1_LOC_718/Y 0.01fF
C8490 INVX1_LOC_25/A INVX1_LOC_30/Y 0.07fF
C8491 NOR2X1_LOC_287/A NOR2X1_LOC_634/Y 0.04fF
C8492 INVX1_LOC_69/Y INVX1_LOC_42/A 0.07fF
C8493 INVX1_LOC_229/A INVX1_LOC_207/A 0.02fF
C8494 INVX1_LOC_21/A INVX1_LOC_168/A 0.03fF
C8495 INVX1_LOC_299/A NOR2X1_LOC_344/A 0.01fF
C8496 INVX1_LOC_45/A D_INPUT_7 0.00fF
C8497 NOR2X1_LOC_598/B NAND2X1_LOC_662/Y 0.01fF
C8498 NOR2X1_LOC_598/B NOR2X1_LOC_730/Y 0.07fF
C8499 NOR2X1_LOC_590/A INVX1_LOC_111/A 0.00fF
C8500 INVX1_LOC_50/A INVX1_LOC_135/A 0.01fF
C8501 INVX1_LOC_227/A INVX1_LOC_23/A 0.08fF
C8502 NAND2X1_LOC_337/B NOR2X1_LOC_433/A 0.06fF
C8503 D_INPUT_1 INVX1_LOC_10/A 4.04fF
C8504 NOR2X1_LOC_78/A NAND2X1_LOC_291/B 0.05fF
C8505 NOR2X1_LOC_246/A NAND2X1_LOC_287/a_36_24# 0.01fF
C8506 INVX1_LOC_1/A NOR2X1_LOC_6/B 0.16fF
C8507 NOR2X1_LOC_631/B INVX1_LOC_19/A 0.32fF
C8508 NOR2X1_LOC_816/A NOR2X1_LOC_433/A 0.01fF
C8509 NOR2X1_LOC_71/Y NAND2X1_LOC_464/B 0.34fF
C8510 NAND2X1_LOC_739/B INVX1_LOC_286/Y 0.03fF
C8511 NOR2X1_LOC_223/B D_GATE_222 0.03fF
C8512 NAND2X1_LOC_728/Y NAND2X1_LOC_741/B 0.00fF
C8513 NOR2X1_LOC_266/a_36_216# NOR2X1_LOC_267/A 0.01fF
C8514 INVX1_LOC_14/A INVX1_LOC_185/Y 0.04fF
C8515 INVX1_LOC_233/Y NAND2X1_LOC_735/B 0.03fF
C8516 NAND2X1_LOC_734/B NAND2X1_LOC_724/A 0.02fF
C8517 NOR2X1_LOC_620/Y NOR2X1_LOC_160/B 0.01fF
C8518 INVX1_LOC_305/A NOR2X1_LOC_68/A 0.05fF
C8519 INVX1_LOC_27/A NOR2X1_LOC_220/A 0.10fF
C8520 INVX1_LOC_225/A NAND2X1_LOC_357/A 0.18fF
C8521 NOR2X1_LOC_186/Y INVX1_LOC_25/Y 0.05fF
C8522 NAND2X1_LOC_500/B INVX1_LOC_20/A 0.01fF
C8523 NAND2X1_LOC_773/Y INVX1_LOC_54/Y 0.01fF
C8524 INVX1_LOC_58/A NOR2X1_LOC_214/B 0.09fF
C8525 INVX1_LOC_57/Y INVX1_LOC_24/A -0.00fF
C8526 INVX1_LOC_269/A NOR2X1_LOC_515/a_36_216# 0.00fF
C8527 INVX1_LOC_272/Y NOR2X1_LOC_591/Y 0.04fF
C8528 INVX1_LOC_59/A NAND2X1_LOC_548/a_36_24# 0.01fF
C8529 NOR2X1_LOC_173/a_36_216# INVX1_LOC_272/A 0.01fF
C8530 NOR2X1_LOC_186/Y NAND2X1_LOC_349/B 0.43fF
C8531 INVX1_LOC_313/Y INVX1_LOC_29/Y 0.01fF
C8532 VDD INVX1_LOC_262/Y 0.26fF
C8533 INVX1_LOC_37/A INVX1_LOC_19/A 0.27fF
C8534 INVX1_LOC_99/Y INVX1_LOC_279/A 0.07fF
C8535 INVX1_LOC_36/Y INVX1_LOC_29/A 0.03fF
C8536 NAND2X1_LOC_352/B INVX1_LOC_162/A 0.18fF
C8537 NOR2X1_LOC_542/Y INVX1_LOC_53/A 0.03fF
C8538 INVX1_LOC_24/Y INVX1_LOC_179/Y 0.19fF
C8539 INVX1_LOC_283/Y NOR2X1_LOC_717/Y 0.18fF
C8540 NOR2X1_LOC_657/a_36_216# INVX1_LOC_22/A 0.00fF
C8541 INVX1_LOC_69/Y INVX1_LOC_78/A 0.07fF
C8542 INVX1_LOC_214/A INVX1_LOC_88/A 0.02fF
C8543 INVX1_LOC_35/A INVX1_LOC_120/A 0.03fF
C8544 NOR2X1_LOC_816/A NOR2X1_LOC_52/B 4.06fF
C8545 NAND2X1_LOC_354/B INVX1_LOC_31/A 0.00fF
C8546 NOR2X1_LOC_791/B INVX1_LOC_71/A 0.00fF
C8547 INVX1_LOC_90/A NOR2X1_LOC_717/A 0.07fF
C8548 INVX1_LOC_24/A NOR2X1_LOC_512/Y 0.00fF
C8549 INVX1_LOC_50/A NOR2X1_LOC_202/Y 0.10fF
C8550 NOR2X1_LOC_703/A INVX1_LOC_23/A 0.07fF
C8551 INVX1_LOC_10/A NOR2X1_LOC_652/Y 0.01fF
C8552 NOR2X1_LOC_389/B NOR2X1_LOC_717/A 0.10fF
C8553 INVX1_LOC_7/Y INVX1_LOC_7/A 0.10fF
C8554 NOR2X1_LOC_401/A NAND2X1_LOC_181/Y 0.01fF
C8555 NOR2X1_LOC_285/Y INVX1_LOC_89/A 0.02fF
C8556 NAND2X1_LOC_30/Y NAND2X1_LOC_451/Y 0.17fF
C8557 NAND2X1_LOC_741/Y INVX1_LOC_229/Y 0.00fF
C8558 NOR2X1_LOC_88/Y INVX1_LOC_92/A 5.65fF
C8559 NAND2X1_LOC_288/A NOR2X1_LOC_743/Y 0.03fF
C8560 NOR2X1_LOC_322/Y INVX1_LOC_57/A 0.13fF
C8561 INVX1_LOC_291/Y INVX1_LOC_231/A 0.01fF
C8562 NOR2X1_LOC_355/A NOR2X1_LOC_674/Y 0.01fF
C8563 INVX1_LOC_249/A NOR2X1_LOC_596/A 0.07fF
C8564 INVX1_LOC_204/Y INVX1_LOC_89/A 0.01fF
C8565 INVX1_LOC_11/A NOR2X1_LOC_773/Y 0.08fF
C8566 NOR2X1_LOC_703/B NOR2X1_LOC_551/B 0.50fF
C8567 NOR2X1_LOC_15/Y INVX1_LOC_290/A 0.00fF
C8568 NAND2X1_LOC_9/Y NOR2X1_LOC_393/a_36_216# 0.00fF
C8569 INVX1_LOC_259/Y NOR2X1_LOC_742/A 0.02fF
C8570 NOR2X1_LOC_753/Y INVX1_LOC_41/Y 0.03fF
C8571 NOR2X1_LOC_92/Y NOR2X1_LOC_561/Y 0.02fF
C8572 INVX1_LOC_45/A NOR2X1_LOC_802/A 0.16fF
C8573 NAND2X1_LOC_181/Y NOR2X1_LOC_160/B 0.03fF
C8574 NOR2X1_LOC_757/A NOR2X1_LOC_122/A 0.12fF
C8575 NOR2X1_LOC_237/a_36_216# NOR2X1_LOC_237/Y 0.03fF
C8576 INVX1_LOC_92/Y INVX1_LOC_57/A 0.05fF
C8577 INVX1_LOC_84/A INVX1_LOC_92/A 0.06fF
C8578 NOR2X1_LOC_802/A NOR2X1_LOC_568/A 0.11fF
C8579 NOR2X1_LOC_13/Y NOR2X1_LOC_172/Y 0.01fF
C8580 NOR2X1_LOC_37/a_36_216# INVX1_LOC_3/Y 0.01fF
C8581 NOR2X1_LOC_540/B NOR2X1_LOC_334/Y 0.01fF
C8582 NOR2X1_LOC_599/Y NAND2X1_LOC_852/Y 0.43fF
C8583 NOR2X1_LOC_770/A INVX1_LOC_49/A 0.02fF
C8584 NOR2X1_LOC_335/B INVX1_LOC_53/A 0.01fF
C8585 NAND2X1_LOC_66/a_36_24# INVX1_LOC_31/A 0.00fF
C8586 INVX1_LOC_31/A NAND2X1_LOC_819/Y 0.04fF
C8587 INVX1_LOC_215/A NOR2X1_LOC_250/A 0.07fF
C8588 NOR2X1_LOC_272/Y NAND2X1_LOC_842/B 0.10fF
C8589 INVX1_LOC_36/A NAND2X1_LOC_342/Y 0.02fF
C8590 INVX1_LOC_12/Y INVX1_LOC_3/Y 0.10fF
C8591 NOR2X1_LOC_488/Y INVX1_LOC_31/A 0.94fF
C8592 INVX1_LOC_24/A NAND2X1_LOC_706/a_36_24# 0.00fF
C8593 INVX1_LOC_19/A NOR2X1_LOC_743/Y 0.71fF
C8594 INVX1_LOC_161/A INVX1_LOC_16/A 0.42fF
C8595 NAND2X1_LOC_222/B NOR2X1_LOC_332/A 0.02fF
C8596 INVX1_LOC_58/A NOR2X1_LOC_741/A 0.03fF
C8597 INVX1_LOC_14/Y INVX1_LOC_4/Y 0.02fF
C8598 INVX1_LOC_33/A INVX1_LOC_275/A 0.15fF
C8599 INVX1_LOC_2/A NOR2X1_LOC_360/Y 0.10fF
C8600 NAND2X1_LOC_651/B INVX1_LOC_92/A 0.03fF
C8601 NOR2X1_LOC_455/Y INVX1_LOC_206/Y 0.02fF
C8602 NAND2X1_LOC_367/A GATE_366 0.00fF
C8603 INVX1_LOC_200/Y NOR2X1_LOC_45/B 0.07fF
C8604 NAND2X1_LOC_208/B INVX1_LOC_16/A 0.00fF
C8605 INVX1_LOC_50/A NOR2X1_LOC_552/A 0.07fF
C8606 NOR2X1_LOC_186/Y INVX1_LOC_75/A 0.15fF
C8607 INVX1_LOC_11/A NOR2X1_LOC_332/A 0.08fF
C8608 NOR2X1_LOC_172/Y NAND2X1_LOC_175/B 0.10fF
C8609 INVX1_LOC_124/A INVX1_LOC_94/A 0.01fF
C8610 INVX1_LOC_117/Y NAND2X1_LOC_74/B 0.00fF
C8611 NOR2X1_LOC_226/A NOR2X1_LOC_360/Y 0.07fF
C8612 NAND2X1_LOC_381/Y NOR2X1_LOC_332/A 0.03fF
C8613 NAND2X1_LOC_722/A NAND2X1_LOC_559/a_36_24# 0.00fF
C8614 NAND2X1_LOC_341/A NOR2X1_LOC_657/Y 0.00fF
C8615 INVX1_LOC_33/A INVX1_LOC_88/Y 0.03fF
C8616 NOR2X1_LOC_188/A INVX1_LOC_50/Y 0.18fF
C8617 INVX1_LOC_181/Y NAND2X1_LOC_850/Y 0.03fF
C8618 NOR2X1_LOC_767/a_36_216# INVX1_LOC_71/A 0.12fF
C8619 INVX1_LOC_93/A NAND2X1_LOC_858/B 0.00fF
C8620 NOR2X1_LOC_266/B INVX1_LOC_26/A 0.02fF
C8621 INVX1_LOC_25/A NOR2X1_LOC_124/A 0.00fF
C8622 INVX1_LOC_223/A NOR2X1_LOC_570/A 0.00fF
C8623 NOR2X1_LOC_91/A NAND2X1_LOC_650/B 0.12fF
C8624 INVX1_LOC_136/A INVX1_LOC_1/Y 0.21fF
C8625 INVX1_LOC_124/Y INVX1_LOC_164/A 0.23fF
C8626 NOR2X1_LOC_67/A NOR2X1_LOC_617/Y 0.02fF
C8627 NAND2X1_LOC_220/B INVX1_LOC_92/A 0.30fF
C8628 INVX1_LOC_26/Y INVX1_LOC_37/A 0.07fF
C8629 INVX1_LOC_135/A INVX1_LOC_61/Y 0.10fF
C8630 NOR2X1_LOC_615/Y NAND2X1_LOC_866/B 0.02fF
C8631 INVX1_LOC_27/A INVX1_LOC_51/Y 0.00fF
C8632 NAND2X1_LOC_717/Y NAND2X1_LOC_864/a_36_24# 0.01fF
C8633 NAND2X1_LOC_357/B INVX1_LOC_162/A 0.34fF
C8634 NAND2X1_LOC_860/A INVX1_LOC_95/Y 0.21fF
C8635 INVX1_LOC_49/A NAND2X1_LOC_451/Y 0.10fF
C8636 NOR2X1_LOC_590/A INVX1_LOC_313/A 0.36fF
C8637 NOR2X1_LOC_168/B INVX1_LOC_33/A 0.13fF
C8638 INVX1_LOC_83/A NOR2X1_LOC_726/Y 0.01fF
C8639 NAND2X1_LOC_72/Y NOR2X1_LOC_552/A 0.05fF
C8640 NOR2X1_LOC_350/A INVX1_LOC_226/A 0.17fF
C8641 INVX1_LOC_226/Y NOR2X1_LOC_403/B 0.01fF
C8642 INVX1_LOC_11/A INVX1_LOC_140/A 0.05fF
C8643 NAND2X1_LOC_562/B NOR2X1_LOC_52/B 0.09fF
C8644 INVX1_LOC_35/A NOR2X1_LOC_542/B 0.01fF
C8645 NOR2X1_LOC_773/Y NOR2X1_LOC_433/A 0.02fF
C8646 INVX1_LOC_15/A INVX1_LOC_92/A 0.11fF
C8647 INVX1_LOC_266/A NOR2X1_LOC_188/A 0.08fF
C8648 NOR2X1_LOC_655/B NAND2X1_LOC_276/Y 0.02fF
C8649 NOR2X1_LOC_355/A INVX1_LOC_72/A 0.07fF
C8650 INVX1_LOC_266/A NOR2X1_LOC_548/B 0.10fF
C8651 NOR2X1_LOC_328/Y NOR2X1_LOC_417/a_36_216# 0.00fF
C8652 INVX1_LOC_45/A NOR2X1_LOC_532/Y 0.02fF
C8653 NOR2X1_LOC_667/A NAND2X1_LOC_734/a_36_24# 0.00fF
C8654 NOR2X1_LOC_690/A INVX1_LOC_280/Y 0.07fF
C8655 NOR2X1_LOC_644/Y NOR2X1_LOC_348/B 0.38fF
C8656 INVX1_LOC_5/A INVX1_LOC_199/A 0.02fF
C8657 NOR2X1_LOC_309/Y NAND2X1_LOC_342/Y 0.01fF
C8658 NAND2X1_LOC_579/A INVX1_LOC_309/A -0.01fF
C8659 NOR2X1_LOC_100/a_36_216# INVX1_LOC_50/Y 0.00fF
C8660 NOR2X1_LOC_620/Y NOR2X1_LOC_516/B 0.03fF
C8661 NOR2X1_LOC_798/A NOR2X1_LOC_405/A 0.03fF
C8662 NAND2X1_LOC_112/Y NOR2X1_LOC_577/Y 1.59fF
C8663 NAND2X1_LOC_338/B INVX1_LOC_60/Y 0.16fF
C8664 NOR2X1_LOC_216/B NOR2X1_LOC_38/B 6.20fF
C8665 NOR2X1_LOC_757/A NOR2X1_LOC_437/Y 0.01fF
C8666 INVX1_LOC_5/A INVX1_LOC_74/A 0.67fF
C8667 INVX1_LOC_279/A NOR2X1_LOC_303/Y 0.10fF
C8668 NAND2X1_LOC_141/A INVX1_LOC_216/A 0.01fF
C8669 NOR2X1_LOC_489/B VDD -0.00fF
C8670 INVX1_LOC_201/Y NOR2X1_LOC_375/Y 0.06fF
C8671 NOR2X1_LOC_518/Y INVX1_LOC_90/A 0.21fF
C8672 NOR2X1_LOC_773/Y NOR2X1_LOC_52/B 0.14fF
C8673 INVX1_LOC_34/A INVX1_LOC_16/A 0.25fF
C8674 NAND2X1_LOC_579/A INVX1_LOC_91/A 0.07fF
C8675 INVX1_LOC_32/A NOR2X1_LOC_673/A 1.38fF
C8676 INVX1_LOC_157/A NOR2X1_LOC_152/Y 0.05fF
C8677 INVX1_LOC_225/A INVX1_LOC_25/Y 0.04fF
C8678 NAND2X1_LOC_803/B INVX1_LOC_6/A 0.02fF
C8679 NAND2X1_LOC_364/A NAND2X1_LOC_842/B 0.01fF
C8680 INVX1_LOC_134/A NOR2X1_LOC_334/A 0.00fF
C8681 INVX1_LOC_27/A NAND2X1_LOC_469/B 0.07fF
C8682 INVX1_LOC_7/Y INVX1_LOC_76/A 0.02fF
C8683 NOR2X1_LOC_582/Y INVX1_LOC_244/A 0.03fF
C8684 INVX1_LOC_102/A INVX1_LOC_29/A 0.04fF
C8685 NOR2X1_LOC_561/A NOR2X1_LOC_717/A 0.01fF
C8686 INVX1_LOC_41/A NOR2X1_LOC_561/Y 0.00fF
C8687 INVX1_LOC_26/A INVX1_LOC_46/Y 0.01fF
C8688 INPUT_2 INVX1_LOC_201/A 0.02fF
C8689 NAND2X1_LOC_740/Y INVX1_LOC_46/A 0.03fF
C8690 NOR2X1_LOC_798/A NOR2X1_LOC_857/A 0.08fF
C8691 INVX1_LOC_33/A NAND2X1_LOC_656/Y 1.12fF
C8692 NAND2X1_LOC_579/A INVX1_LOC_11/Y 0.07fF
C8693 INVX1_LOC_279/A NOR2X1_LOC_254/Y 0.01fF
C8694 INVX1_LOC_1/A NOR2X1_LOC_124/A 0.08fF
C8695 NOR2X1_LOC_590/A INVX1_LOC_6/A 0.03fF
C8696 NOR2X1_LOC_89/A INVX1_LOC_42/A 0.35fF
C8697 NAND2X1_LOC_464/B NAND2X1_LOC_243/Y 0.00fF
C8698 NOR2X1_LOC_483/B INVX1_LOC_78/Y 0.01fF
C8699 NOR2X1_LOC_644/Y INVX1_LOC_22/A 0.01fF
C8700 NAND2X1_LOC_276/Y NOR2X1_LOC_99/B 0.07fF
C8701 INVX1_LOC_14/A NAND2X1_LOC_659/B 0.02fF
C8702 NOR2X1_LOC_561/Y NAND2X1_LOC_477/A 0.01fF
C8703 NOR2X1_LOC_209/Y NOR2X1_LOC_302/B 0.00fF
C8704 NOR2X1_LOC_858/A NOR2X1_LOC_676/Y 0.20fF
C8705 NOR2X1_LOC_92/Y INVX1_LOC_76/A 0.17fF
C8706 INVX1_LOC_33/A INVX1_LOC_132/Y 0.03fF
C8707 NAND2X1_LOC_550/A NAND2X1_LOC_623/B 0.05fF
C8708 NOR2X1_LOC_383/B NOR2X1_LOC_197/B 0.01fF
C8709 NAND2X1_LOC_725/B INVX1_LOC_20/A 0.07fF
C8710 NOR2X1_LOC_376/A VDD -0.00fF
C8711 NAND2X1_LOC_740/Y NOR2X1_LOC_766/Y 0.02fF
C8712 NOR2X1_LOC_781/A NAND2X1_LOC_661/B 0.09fF
C8713 NOR2X1_LOC_781/B INVX1_LOC_266/Y 0.00fF
C8714 NAND2X1_LOC_569/A NOR2X1_LOC_76/A -0.02fF
C8715 INVX1_LOC_90/A NAND2X1_LOC_175/B 0.12fF
C8716 NAND2X1_LOC_706/Y INVX1_LOC_46/A 0.10fF
C8717 D_INPUT_1 INVX1_LOC_307/A 0.01fF
C8718 INVX1_LOC_165/A NAND2X1_LOC_773/B 0.01fF
C8719 NOR2X1_LOC_433/A INVX1_LOC_140/A 0.03fF
C8720 NOR2X1_LOC_779/Y VDD 0.14fF
C8721 NOR2X1_LOC_553/Y NOR2X1_LOC_500/Y 0.03fF
C8722 NAND2X1_LOC_72/B INVX1_LOC_19/A 0.03fF
C8723 INVX1_LOC_90/A NAND2X1_LOC_142/a_36_24# 0.00fF
C8724 NAND2X1_LOC_568/A INVX1_LOC_76/A 0.01fF
C8725 INVX1_LOC_49/A NOR2X1_LOC_567/B 0.07fF
C8726 INVX1_LOC_14/A VDD 5.40fF
C8727 NOR2X1_LOC_772/a_36_216# INVX1_LOC_16/A 0.00fF
C8728 INVX1_LOC_270/A INVX1_LOC_285/A 0.02fF
C8729 NOR2X1_LOC_763/Y INVX1_LOC_191/Y 0.01fF
C8730 INVX1_LOC_34/A INVX1_LOC_28/A 0.14fF
C8731 NOR2X1_LOC_246/Y NOR2X1_LOC_309/Y 0.01fF
C8732 INVX1_LOC_53/A NOR2X1_LOC_88/Y 0.15fF
C8733 NOR2X1_LOC_205/Y INVX1_LOC_14/Y 0.06fF
C8734 NOR2X1_LOC_295/Y NOR2X1_LOC_772/A 0.53fF
C8735 INVX1_LOC_45/A NOR2X1_LOC_192/A 0.05fF
C8736 NOR2X1_LOC_488/Y NAND2X1_LOC_859/Y 0.02fF
C8737 NAND2X1_LOC_112/Y INVX1_LOC_22/A 0.05fF
C8738 INVX1_LOC_36/A INVX1_LOC_70/Y 0.17fF
C8739 INVX1_LOC_73/A INVX1_LOC_155/A 2.49fF
C8740 NOR2X1_LOC_474/A NAND2X1_LOC_463/B 0.01fF
C8741 NOR2X1_LOC_793/A INVX1_LOC_117/A 0.03fF
C8742 INVX1_LOC_270/A NOR2X1_LOC_814/A 0.07fF
C8743 INVX1_LOC_136/A NOR2X1_LOC_318/B 0.05fF
C8744 INVX1_LOC_90/A NOR2X1_LOC_504/Y 0.07fF
C8745 NOR2X1_LOC_89/A INVX1_LOC_78/A 0.26fF
C8746 INVX1_LOC_161/Y NOR2X1_LOC_681/Y 0.01fF
C8747 NAND2X1_LOC_807/A NAND2X1_LOC_287/B 0.04fF
C8748 INVX1_LOC_161/Y INVX1_LOC_37/A 0.03fF
C8749 NAND2X1_LOC_59/B NAND2X1_LOC_51/B 0.30fF
C8750 INVX1_LOC_241/A INVX1_LOC_229/Y 0.14fF
C8751 INVX1_LOC_136/A INVX1_LOC_93/Y 0.29fF
C8752 INVX1_LOC_53/A INVX1_LOC_84/A 0.13fF
C8753 NOR2X1_LOC_52/B INVX1_LOC_140/A 0.80fF
C8754 INVX1_LOC_225/A INVX1_LOC_75/A 0.07fF
C8755 INVX1_LOC_35/A NAND2X1_LOC_659/A 0.21fF
C8756 NAND2X1_LOC_231/Y INVX1_LOC_28/A 0.10fF
C8757 INVX1_LOC_174/A NAND2X1_LOC_51/a_36_24# 0.01fF
C8758 NOR2X1_LOC_383/Y NOR2X1_LOC_383/a_36_216# 0.02fF
C8759 INVX1_LOC_294/Y NOR2X1_LOC_292/Y 0.00fF
C8760 NOR2X1_LOC_109/Y INVX1_LOC_285/A 0.07fF
C8761 NOR2X1_LOC_65/B NOR2X1_LOC_89/A 0.17fF
C8762 INVX1_LOC_78/A NOR2X1_LOC_170/A 0.04fF
C8763 INVX1_LOC_18/A NAND2X1_LOC_447/Y 0.10fF
C8764 NOR2X1_LOC_160/B INVX1_LOC_117/A 9.06fF
C8765 NOR2X1_LOC_6/B NOR2X1_LOC_188/A 0.86fF
C8766 NOR2X1_LOC_717/Y VDD 0.25fF
C8767 INVX1_LOC_229/Y NOR2X1_LOC_298/Y 0.93fF
C8768 INVX1_LOC_215/A NOR2X1_LOC_106/A 0.01fF
C8769 NOR2X1_LOC_393/Y INVX1_LOC_165/A 0.00fF
C8770 NOR2X1_LOC_103/Y NAND2X1_LOC_276/a_36_24# 0.00fF
C8771 NAND2X1_LOC_538/Y INVX1_LOC_54/A 0.07fF
C8772 NOR2X1_LOC_209/Y INVX1_LOC_75/A 0.07fF
C8773 NOR2X1_LOC_577/Y NOR2X1_LOC_78/A 0.07fF
C8774 NOR2X1_LOC_486/Y NOR2X1_LOC_546/B 0.03fF
C8775 INVX1_LOC_61/Y NOR2X1_LOC_813/Y 0.49fF
C8776 NOR2X1_LOC_454/Y NOR2X1_LOC_155/A 0.07fF
C8777 INVX1_LOC_213/Y NOR2X1_LOC_728/B 0.05fF
C8778 D_INPUT_1 INVX1_LOC_12/A 0.12fF
C8779 INVX1_LOC_78/A INVX1_LOC_104/Y 0.01fF
C8780 INVX1_LOC_313/Y INVX1_LOC_101/A 0.01fF
C8781 NOR2X1_LOC_158/B NOR2X1_LOC_158/Y 0.01fF
C8782 NOR2X1_LOC_497/a_36_216# NAND2X1_LOC_254/Y 0.00fF
C8783 INVX1_LOC_227/Y VDD 0.41fF
C8784 INVX1_LOC_227/A INVX1_LOC_313/A 0.10fF
C8785 NOR2X1_LOC_468/Y NOR2X1_LOC_216/B 0.01fF
C8786 NOR2X1_LOC_295/a_36_216# INVX1_LOC_91/A 0.01fF
C8787 INVX1_LOC_136/A NAND2X1_LOC_721/A 0.02fF
C8788 INVX1_LOC_61/Y INVX1_LOC_280/A 0.02fF
C8789 INVX1_LOC_286/A NOR2X1_LOC_709/A 0.10fF
C8790 NAND2X1_LOC_837/Y INVX1_LOC_76/A 0.08fF
C8791 NOR2X1_LOC_522/Y VDD 0.13fF
C8792 NOR2X1_LOC_486/Y INVX1_LOC_275/A 0.14fF
C8793 NOR2X1_LOC_561/Y NOR2X1_LOC_122/Y 0.03fF
C8794 NAND2X1_LOC_739/B VDD 0.01fF
C8795 NOR2X1_LOC_208/Y NOR2X1_LOC_562/A 0.01fF
C8796 INVX1_LOC_182/A NOR2X1_LOC_553/B 0.02fF
C8797 NOR2X1_LOC_30/Y NOR2X1_LOC_25/Y 0.17fF
C8798 NAND2X1_LOC_739/B NAND2X1_LOC_800/A 0.47fF
C8799 NOR2X1_LOC_355/A INVX1_LOC_313/Y 0.00fF
C8800 NAND2X1_LOC_84/Y VDD 0.08fF
C8801 NAND2X1_LOC_116/A NAND2X1_LOC_86/Y 0.08fF
C8802 NAND2X1_LOC_53/Y NAND2X1_LOC_435/a_36_24# 0.01fF
C8803 NOR2X1_LOC_241/A NOR2X1_LOC_445/B 0.00fF
C8804 INPUT_0 INVX1_LOC_16/A 0.47fF
C8805 INVX1_LOC_217/Y NAND2X1_LOC_659/B -0.02fF
C8806 INVX1_LOC_83/A INVX1_LOC_311/Y 0.03fF
C8807 NOR2X1_LOC_590/A INVX1_LOC_131/Y 0.01fF
C8808 INVX1_LOC_34/A NOR2X1_LOC_253/Y 0.04fF
C8809 INVX1_LOC_2/A NOR2X1_LOC_269/Y 0.15fF
C8810 NOR2X1_LOC_488/Y INVX1_LOC_6/A 0.01fF
C8811 INVX1_LOC_12/A NOR2X1_LOC_652/Y 0.03fF
C8812 INVX1_LOC_41/A INVX1_LOC_76/A 0.04fF
C8813 INVX1_LOC_21/A INVX1_LOC_272/A 0.07fF
C8814 INVX1_LOC_269/A NAND2X1_LOC_475/Y 0.10fF
C8815 NAND2X1_LOC_20/B NAND2X1_LOC_574/A 0.06fF
C8816 NAND2X1_LOC_149/Y NOR2X1_LOC_48/a_36_216# 0.01fF
C8817 INVX1_LOC_53/A INVX1_LOC_15/A 2.79fF
C8818 NOR2X1_LOC_363/Y INVX1_LOC_71/A 0.02fF
C8819 NOR2X1_LOC_82/Y INVX1_LOC_6/A 0.06fF
C8820 NOR2X1_LOC_498/Y INVX1_LOC_76/A 0.07fF
C8821 INVX1_LOC_72/A INVX1_LOC_127/A 0.01fF
C8822 INVX1_LOC_30/Y NOR2X1_LOC_188/A 0.07fF
C8823 NOR2X1_LOC_730/B NOR2X1_LOC_687/Y 0.04fF
C8824 INVX1_LOC_304/A INVX1_LOC_168/A 0.11fF
C8825 INVX1_LOC_312/A NOR2X1_LOC_743/Y 0.00fF
C8826 INVX1_LOC_30/Y NOR2X1_LOC_548/B 0.03fF
C8827 NOR2X1_LOC_445/Y INVX1_LOC_46/A 0.01fF
C8828 INVX1_LOC_193/Y INVX1_LOC_174/Y 0.89fF
C8829 INVX1_LOC_217/Y VDD 0.87fF
C8830 NOR2X1_LOC_13/Y INVX1_LOC_38/A 0.06fF
C8831 INVX1_LOC_94/A INVX1_LOC_9/A 0.90fF
C8832 NAND2X1_LOC_477/A INVX1_LOC_76/A 0.07fF
C8833 NOR2X1_LOC_82/A INVX1_LOC_293/Y 0.15fF
C8834 INVX1_LOC_178/A NAND2X1_LOC_254/Y 0.01fF
C8835 INVX1_LOC_82/A D_INPUT_3 0.01fF
C8836 NOR2X1_LOC_139/Y NOR2X1_LOC_131/Y 0.02fF
C8837 INVX1_LOC_208/Y INVX1_LOC_91/A 0.01fF
C8838 INVX1_LOC_98/A INVX1_LOC_22/A 0.10fF
C8839 INVX1_LOC_190/A INVX1_LOC_144/A 0.03fF
C8840 INVX1_LOC_136/A INVX1_LOC_117/Y 0.05fF
C8841 INPUT_3 NOR2X1_LOC_673/A 0.07fF
C8842 INVX1_LOC_13/Y INVX1_LOC_19/Y 0.00fF
C8843 INVX1_LOC_266/Y NOR2X1_LOC_585/Y 0.01fF
C8844 NOR2X1_LOC_218/Y NOR2X1_LOC_269/Y 0.01fF
C8845 INVX1_LOC_227/A INVX1_LOC_6/A 0.01fF
C8846 NAND2X1_LOC_175/a_36_24# INVX1_LOC_12/A 0.00fF
C8847 NOR2X1_LOC_78/A INVX1_LOC_22/A 0.71fF
C8848 NOR2X1_LOC_638/Y NOR2X1_LOC_654/A 0.02fF
C8849 INVX1_LOC_25/Y NAND2X1_LOC_642/Y 0.02fF
C8850 NAND2X1_LOC_30/Y NOR2X1_LOC_36/B 0.01fF
C8851 VDD NOR2X1_LOC_612/B 0.00fF
C8852 NOR2X1_LOC_589/A NOR2X1_LOC_139/Y 0.01fF
C8853 NAND2X1_LOC_175/B INVX1_LOC_38/A 0.46fF
C8854 NOR2X1_LOC_131/Y NAND2X1_LOC_468/B 0.01fF
C8855 INVX1_LOC_223/A NAND2X1_LOC_606/a_36_24# 0.00fF
C8856 NOR2X1_LOC_242/A INVX1_LOC_15/A 0.04fF
C8857 INVX1_LOC_27/A INVX1_LOC_251/A 0.01fF
C8858 NAND2X1_LOC_51/B INVX1_LOC_244/A 0.23fF
C8859 INVX1_LOC_111/Y VDD 0.07fF
C8860 INVX1_LOC_36/A INVX1_LOC_285/A 0.14fF
C8861 NOR2X1_LOC_82/A NAND2X1_LOC_74/B 0.33fF
C8862 NAND2X1_LOC_721/A NAND2X1_LOC_859/a_36_24# 0.00fF
C8863 NOR2X1_LOC_660/Y INVX1_LOC_175/A 0.70fF
C8864 INVX1_LOC_24/A INVX1_LOC_179/A 0.04fF
C8865 NAND2X1_LOC_483/a_36_24# INVX1_LOC_46/A 0.00fF
C8866 NOR2X1_LOC_753/Y INVX1_LOC_185/A 0.03fF
C8867 INVX1_LOC_207/A INVX1_LOC_118/A 0.69fF
C8868 INVX1_LOC_28/A INPUT_0 0.49fF
C8869 INVX1_LOC_36/A NOR2X1_LOC_814/A 0.03fF
C8870 INVX1_LOC_40/Y INVX1_LOC_63/A 0.04fF
C8871 INVX1_LOC_11/A NOR2X1_LOC_847/A 0.00fF
C8872 NAND2X1_LOC_656/A NOR2X1_LOC_831/B 0.01fF
C8873 NAND2X1_LOC_538/Y NOR2X1_LOC_48/B 0.07fF
C8874 INVX1_LOC_189/A INVX1_LOC_117/A -0.02fF
C8875 NOR2X1_LOC_589/A NAND2X1_LOC_468/B 0.03fF
C8876 INVX1_LOC_11/A INVX1_LOC_42/A 2.01fF
C8877 NAND2X1_LOC_381/Y NOR2X1_LOC_847/A 0.03fF
C8878 NOR2X1_LOC_82/A NOR2X1_LOC_847/B -0.00fF
C8879 NOR2X1_LOC_503/Y NOR2X1_LOC_89/A 0.19fF
C8880 NOR2X1_LOC_590/A NOR2X1_LOC_633/A 0.03fF
C8881 INVX1_LOC_77/A NOR2X1_LOC_155/A 0.13fF
C8882 NAND2X1_LOC_325/Y INVX1_LOC_185/A 0.00fF
C8883 NAND2X1_LOC_114/B INVX1_LOC_106/Y 0.01fF
C8884 INVX1_LOC_140/Y INVX1_LOC_140/A 0.10fF
C8885 NAND2X1_LOC_361/Y NOR2X1_LOC_862/B 0.10fF
C8886 NAND2X1_LOC_514/a_36_24# NAND2X1_LOC_211/Y 0.01fF
C8887 NOR2X1_LOC_750/Y NOR2X1_LOC_392/Y 0.02fF
C8888 NOR2X1_LOC_292/Y NOR2X1_LOC_74/A 0.01fF
C8889 INVX1_LOC_173/Y INPUT_4 0.03fF
C8890 NOR2X1_LOC_332/A INVX1_LOC_74/A 0.02fF
C8891 INVX1_LOC_223/A INVX1_LOC_29/A 0.81fF
C8892 NOR2X1_LOC_298/Y INVX1_LOC_20/A 0.03fF
C8893 NOR2X1_LOC_516/B INVX1_LOC_117/A 4.19fF
C8894 NOR2X1_LOC_756/Y INVX1_LOC_91/A 0.26fF
C8895 NOR2X1_LOC_732/A NOR2X1_LOC_155/A 0.02fF
C8896 NAND2X1_LOC_354/Y INVX1_LOC_272/A 0.00fF
C8897 INVX1_LOC_164/A NOR2X1_LOC_266/B 0.16fF
C8898 NOR2X1_LOC_299/Y INVX1_LOC_76/A 0.03fF
C8899 NAND2X1_LOC_842/B NOR2X1_LOC_405/A 0.08fF
C8900 NAND2X1_LOC_198/B INVX1_LOC_19/A 0.03fF
C8901 NOR2X1_LOC_160/B INVX1_LOC_3/Y 0.07fF
C8902 INVX1_LOC_72/A NOR2X1_LOC_583/Y 0.03fF
C8903 NOR2X1_LOC_360/Y NAND2X1_LOC_63/Y 0.05fF
C8904 INVX1_LOC_28/A NAND2X1_LOC_649/B 0.04fF
C8905 NOR2X1_LOC_136/Y INVX1_LOC_9/A 0.01fF
C8906 NOR2X1_LOC_192/A INVX1_LOC_102/Y 0.05fF
C8907 INVX1_LOC_25/Y NOR2X1_LOC_271/Y 0.10fF
C8908 INVX1_LOC_224/A INVX1_LOC_78/A 0.06fF
C8909 INVX1_LOC_254/Y NOR2X1_LOC_68/Y 0.03fF
C8910 NOR2X1_LOC_137/A VDD 0.15fF
C8911 INVX1_LOC_11/A INVX1_LOC_78/A 9.55fF
C8912 NAND2X1_LOC_117/a_36_24# NOR2X1_LOC_266/B 0.00fF
C8913 INVX1_LOC_196/A NOR2X1_LOC_461/A 0.01fF
C8914 NOR2X1_LOC_309/Y INVX1_LOC_285/A 0.12fF
C8915 INVX1_LOC_75/A NAND2X1_LOC_642/Y 0.03fF
C8916 NAND2X1_LOC_671/a_36_24# NOR2X1_LOC_655/Y 0.01fF
C8917 NOR2X1_LOC_309/Y INVX1_LOC_265/Y 0.04fF
C8918 NOR2X1_LOC_226/A NOR2X1_LOC_79/Y 0.03fF
C8919 NOR2X1_LOC_309/Y NOR2X1_LOC_814/A 0.03fF
C8920 INVX1_LOC_310/Y INVX1_LOC_19/A 0.06fF
C8921 NOR2X1_LOC_19/B NAND2X1_LOC_414/a_36_24# 0.01fF
C8922 NAND2X1_LOC_785/A INVX1_LOC_119/Y 0.07fF
C8923 NOR2X1_LOC_152/Y NOR2X1_LOC_89/A 0.07fF
C8924 NOR2X1_LOC_454/Y NOR2X1_LOC_598/B 0.10fF
C8925 INVX1_LOC_245/A NAND2X1_LOC_93/B 0.01fF
C8926 NAND2X1_LOC_756/a_36_24# NOR2X1_LOC_331/B 0.01fF
C8927 INVX1_LOC_25/A NOR2X1_LOC_15/Y 0.01fF
C8928 NOR2X1_LOC_808/A NOR2X1_LOC_801/A 0.07fF
C8929 NOR2X1_LOC_501/B INVX1_LOC_91/A 0.03fF
C8930 INVX1_LOC_77/A NOR2X1_LOC_833/B 0.04fF
C8931 INVX1_LOC_113/Y NOR2X1_LOC_89/A 0.03fF
C8932 INVX1_LOC_64/A NOR2X1_LOC_61/B 0.27fF
C8933 NOR2X1_LOC_687/Y NOR2X1_LOC_155/A 7.28fF
C8934 NOR2X1_LOC_433/A INVX1_LOC_42/A 0.24fF
C8935 INPUT_0 NOR2X1_LOC_35/Y 0.03fF
C8936 NOR2X1_LOC_474/A INVX1_LOC_42/A 0.00fF
C8937 D_INPUT_1 INVX1_LOC_228/Y 0.04fF
C8938 NOR2X1_LOC_78/B INVX1_LOC_84/A 5.89fF
C8939 INVX1_LOC_53/Y NAND2X1_LOC_288/A 0.07fF
C8940 INVX1_LOC_162/Y INVX1_LOC_29/A 0.26fF
C8941 NOR2X1_LOC_86/A NAND2X1_LOC_243/B 0.15fF
C8942 NOR2X1_LOC_483/B NOR2X1_LOC_727/B 0.02fF
C8943 NOR2X1_LOC_593/Y INVX1_LOC_42/A 0.03fF
C8944 NAND2X1_LOC_138/a_36_24# NAND2X1_LOC_211/Y 0.01fF
C8945 INVX1_LOC_184/A INVX1_LOC_15/A 0.05fF
C8946 INVX1_LOC_64/A NAND2X1_LOC_725/B 0.18fF
C8947 INVX1_LOC_136/A INVX1_LOC_87/A 0.10fF
C8948 INVX1_LOC_58/A NAND2X1_LOC_550/A 0.07fF
C8949 INVX1_LOC_64/A INVX1_LOC_101/Y 0.01fF
C8950 NOR2X1_LOC_15/Y NAND2X1_LOC_360/a_36_24# 0.00fF
C8951 NOR2X1_LOC_335/B INVX1_LOC_46/A 0.05fF
C8952 NOR2X1_LOC_387/A NOR2X1_LOC_421/Y 0.00fF
C8953 NAND2X1_LOC_660/Y NOR2X1_LOC_832/a_36_216# 0.02fF
C8954 NOR2X1_LOC_590/A INVX1_LOC_270/A 0.04fF
C8955 NOR2X1_LOC_441/Y NAND2X1_LOC_285/a_36_24# 0.00fF
C8956 NOR2X1_LOC_706/A INVX1_LOC_117/A 0.02fF
C8957 INVX1_LOC_58/A NOR2X1_LOC_160/B 0.07fF
C8958 INVX1_LOC_236/Y NOR2X1_LOC_654/A 0.00fF
C8959 NOR2X1_LOC_824/A NOR2X1_LOC_496/Y 0.04fF
C8960 INVX1_LOC_11/A INVX1_LOC_152/Y 0.01fF
C8961 D_INPUT_0 NOR2X1_LOC_235/Y 0.02fF
C8962 NOR2X1_LOC_82/A NOR2X1_LOC_660/Y 0.30fF
C8963 INVX1_LOC_24/A INVX1_LOC_165/A 0.01fF
C8964 INVX1_LOC_254/A INVX1_LOC_4/Y 0.02fF
C8965 NOR2X1_LOC_52/B INVX1_LOC_42/A 8.06fF
C8966 NAND2X1_LOC_231/Y INVX1_LOC_109/A 0.06fF
C8967 INVX1_LOC_255/Y NAND2X1_LOC_206/Y 0.08fF
C8968 NOR2X1_LOC_468/Y INVX1_LOC_93/A 0.04fF
C8969 VDD INVX1_LOC_48/A 0.12fF
C8970 NAND2X1_LOC_724/Y NAND2X1_LOC_741/B 0.03fF
C8971 INVX1_LOC_7/A NAND2X1_LOC_574/A 0.02fF
C8972 NOR2X1_LOC_561/Y NOR2X1_LOC_435/B 0.05fF
C8973 INVX1_LOC_21/A INVX1_LOC_198/A 0.03fF
C8974 INVX1_LOC_75/A NOR2X1_LOC_271/Y 0.06fF
C8975 NAND2X1_LOC_763/B NAND2X1_LOC_64/a_36_24# -0.02fF
C8976 NAND2X1_LOC_803/B NOR2X1_LOC_109/Y 0.00fF
C8977 INVX1_LOC_191/A INVX1_LOC_77/Y 0.04fF
C8978 INVX1_LOC_45/A INVX1_LOC_29/Y 0.03fF
C8979 NAND2X1_LOC_655/A INVX1_LOC_20/A 0.28fF
C8980 INVX1_LOC_53/Y INVX1_LOC_19/A 0.03fF
C8981 NOR2X1_LOC_459/A INVX1_LOC_84/A 0.47fF
C8982 NOR2X1_LOC_433/A INVX1_LOC_78/A 0.14fF
C8983 NOR2X1_LOC_619/A INVX1_LOC_19/A 0.06fF
C8984 D_INPUT_2 NOR2X1_LOC_29/a_36_216# 0.00fF
C8985 INVX1_LOC_16/A NOR2X1_LOC_84/B -0.01fF
C8986 INVX1_LOC_313/Y NOR2X1_LOC_600/a_36_216# 0.00fF
C8987 NOR2X1_LOC_635/A NOR2X1_LOC_467/A 0.01fF
C8988 INVX1_LOC_24/A NOR2X1_LOC_693/Y 0.11fF
C8989 NOR2X1_LOC_337/A INVX1_LOC_38/A 0.03fF
C8990 NOR2X1_LOC_84/A NOR2X1_LOC_38/B 0.06fF
C8991 NAND2X1_LOC_468/B INVX1_LOC_147/Y 0.48fF
C8992 INVX1_LOC_58/A NAND2X1_LOC_195/Y 0.01fF
C8993 NOR2X1_LOC_771/a_36_216# NAND2X1_LOC_93/B 0.00fF
C8994 NOR2X1_LOC_593/Y INVX1_LOC_78/A 0.07fF
C8995 INVX1_LOC_90/A NAND2X1_LOC_85/Y 0.03fF
C8996 INVX1_LOC_83/A INVX1_LOC_84/A 0.03fF
C8997 NOR2X1_LOC_570/B NOR2X1_LOC_334/Y 0.08fF
C8998 NOR2X1_LOC_590/A NOR2X1_LOC_109/Y 0.04fF
C8999 INVX1_LOC_103/A NAND2X1_LOC_714/B 0.01fF
C9000 INVX1_LOC_90/A NOR2X1_LOC_697/Y 0.12fF
C9001 INVX1_LOC_58/A NOR2X1_LOC_733/a_36_216# 0.00fF
C9002 NOR2X1_LOC_15/Y INVX1_LOC_1/A 0.14fF
C9003 INVX1_LOC_49/A INVX1_LOC_26/A 0.00fF
C9004 NOR2X1_LOC_716/B NOR2X1_LOC_278/Y 0.02fF
C9005 NAND2X1_LOC_662/Y INVX1_LOC_29/A 0.00fF
C9006 INVX1_LOC_306/A INVX1_LOC_293/Y 0.09fF
C9007 NOR2X1_LOC_771/a_36_216# NAND2X1_LOC_425/Y 0.01fF
C9008 NOR2X1_LOC_634/B INVX1_LOC_15/A 0.03fF
C9009 INVX1_LOC_177/A NAND2X1_LOC_761/a_36_24# 0.02fF
C9010 NOR2X1_LOC_65/B NOR2X1_LOC_433/A 0.10fF
C9011 NOR2X1_LOC_687/Y NOR2X1_LOC_833/B 0.05fF
C9012 NOR2X1_LOC_78/B INVX1_LOC_15/A 0.36fF
C9013 NOR2X1_LOC_9/Y NOR2X1_LOC_641/Y 0.03fF
C9014 NOR2X1_LOC_86/A INVX1_LOC_284/A 0.19fF
C9015 NOR2X1_LOC_52/B INVX1_LOC_78/A 2.97fF
C9016 INVX1_LOC_310/Y INVX1_LOC_26/Y 0.25fF
C9017 INVX1_LOC_71/A INVX1_LOC_29/Y 1.00fF
C9018 NOR2X1_LOC_65/B NOR2X1_LOC_593/Y 0.22fF
C9019 INVX1_LOC_83/A NAND2X1_LOC_651/B 0.03fF
C9020 INVX1_LOC_178/A NAND2X1_LOC_354/a_36_24# 0.06fF
C9021 INVX1_LOC_306/A NAND2X1_LOC_74/B 0.02fF
C9022 NAND2X1_LOC_51/B INVX1_LOC_107/Y 0.02fF
C9023 NOR2X1_LOC_540/B NAND2X1_LOC_472/Y 0.04fF
C9024 INVX1_LOC_269/A NOR2X1_LOC_457/A 0.28fF
C9025 INVX1_LOC_60/A INVX1_LOC_26/A 0.03fF
C9026 NOR2X1_LOC_516/B INVX1_LOC_3/Y 0.07fF
C9027 INVX1_LOC_149/A NAND2X1_LOC_71/a_36_24# 0.00fF
C9028 NAND2X1_LOC_833/Y INVX1_LOC_57/A 0.05fF
C9029 NAND2X1_LOC_160/a_36_24# NOR2X1_LOC_467/A 0.00fF
C9030 NOR2X1_LOC_598/B INVX1_LOC_77/A 0.98fF
C9031 INVX1_LOC_48/Y NAND2X1_LOC_208/B 0.02fF
C9032 INVX1_LOC_288/A NOR2X1_LOC_52/B 0.00fF
C9033 INVX1_LOC_63/Y INVX1_LOC_271/A 0.00fF
C9034 NOR2X1_LOC_753/Y NOR2X1_LOC_754/Y 0.01fF
C9035 NOR2X1_LOC_272/Y INVX1_LOC_72/A 0.04fF
C9036 NOR2X1_LOC_65/B NOR2X1_LOC_52/B 0.12fF
C9037 INVX1_LOC_205/A NOR2X1_LOC_249/Y 0.20fF
C9038 INVX1_LOC_2/A INVX1_LOC_26/A 0.01fF
C9039 INVX1_LOC_1/Y NAND2X1_LOC_647/B 0.01fF
C9040 NOR2X1_LOC_669/Y INVX1_LOC_141/Y 0.01fF
C9041 NAND2X1_LOC_21/Y INVX1_LOC_53/A 0.07fF
C9042 NAND2X1_LOC_794/B NOR2X1_LOC_518/a_36_216# 0.01fF
C9043 NAND2X1_LOC_796/B INVX1_LOC_18/A 0.68fF
C9044 INVX1_LOC_120/A NAND2X1_LOC_206/B 0.12fF
C9045 INPUT_5 D_INPUT_5 2.31fF
C9046 INVX1_LOC_33/A NOR2X1_LOC_717/A 0.00fF
C9047 INVX1_LOC_89/A NOR2X1_LOC_461/Y 0.07fF
C9048 NOR2X1_LOC_226/A INVX1_LOC_26/A 0.12fF
C9049 INVX1_LOC_5/A INVX1_LOC_314/Y 0.34fF
C9050 INVX1_LOC_104/A INVX1_LOC_23/A 0.27fF
C9051 INVX1_LOC_269/A INVX1_LOC_30/A 0.19fF
C9052 INVX1_LOC_215/A NOR2X1_LOC_334/Y 0.01fF
C9053 NOR2X1_LOC_455/Y NOR2X1_LOC_455/a_36_216# 0.02fF
C9054 NOR2X1_LOC_441/Y NOR2X1_LOC_250/A 0.03fF
C9055 INVX1_LOC_133/Y INVX1_LOC_270/Y 0.00fF
C9056 NOR2X1_LOC_168/B NOR2X1_LOC_748/A 0.14fF
C9057 INVX1_LOC_83/A INVX1_LOC_15/A 0.79fF
C9058 NOR2X1_LOC_15/Y NOR2X1_LOC_384/Y 0.15fF
C9059 INVX1_LOC_233/Y NOR2X1_LOC_690/A 0.10fF
C9060 INVX1_LOC_267/Y INVX1_LOC_166/A 0.06fF
C9061 NAND2X1_LOC_262/a_36_24# NOR2X1_LOC_536/A 0.01fF
C9062 INVX1_LOC_41/A NOR2X1_LOC_178/Y 0.07fF
C9063 NOR2X1_LOC_471/Y NOR2X1_LOC_477/a_36_216# 0.02fF
C9064 INVX1_LOC_227/A NAND2X1_LOC_646/a_36_24# 0.00fF
C9065 NOR2X1_LOC_318/B NOR2X1_LOC_117/a_36_216# 0.00fF
C9066 INVX1_LOC_286/A INVX1_LOC_294/A 0.02fF
C9067 NOR2X1_LOC_667/a_36_216# NOR2X1_LOC_590/A 0.02fF
C9068 NOR2X1_LOC_186/Y NOR2X1_LOC_577/Y 0.01fF
C9069 NOR2X1_LOC_232/a_36_216# INVX1_LOC_18/A 0.00fF
C9070 NAND2X1_LOC_222/B NOR2X1_LOC_554/B 0.00fF
C9071 NAND2X1_LOC_740/Y NAND2X1_LOC_812/A 0.02fF
C9072 NOR2X1_LOC_113/B INVX1_LOC_19/A 0.76fF
C9073 NOR2X1_LOC_619/A INVX1_LOC_26/Y 0.03fF
C9074 NOR2X1_LOC_666/Y NOR2X1_LOC_457/B 0.20fF
C9075 NAND2X1_LOC_803/B INVX1_LOC_36/A 0.03fF
C9076 NOR2X1_LOC_363/Y NOR2X1_LOC_331/B 0.81fF
C9077 INVX1_LOC_136/A NOR2X1_LOC_82/A 0.04fF
C9078 NAND2X1_LOC_563/Y NOR2X1_LOC_662/a_36_216# 0.01fF
C9079 INVX1_LOC_58/A NAND2X1_LOC_350/B 0.01fF
C9080 INVX1_LOC_11/A NOR2X1_LOC_554/B 0.00fF
C9081 INVX1_LOC_64/A NOR2X1_LOC_398/a_36_216# 0.00fF
C9082 NOR2X1_LOC_756/a_36_216# INVX1_LOC_3/Y 0.00fF
C9083 NOR2X1_LOC_27/Y NAND2X1_LOC_725/A 0.02fF
C9084 NOR2X1_LOC_261/Y NOR2X1_LOC_78/B 0.01fF
C9085 NOR2X1_LOC_828/Y NOR2X1_LOC_778/B 0.13fF
C9086 INVX1_LOC_222/Y NOR2X1_LOC_344/A 0.14fF
C9087 INVX1_LOC_95/Y NOR2X1_LOC_49/a_36_216# 0.00fF
C9088 INVX1_LOC_34/A NAND2X1_LOC_794/B 0.07fF
C9089 NAND2X1_LOC_381/Y NOR2X1_LOC_554/B 0.04fF
C9090 NOR2X1_LOC_273/Y INVX1_LOC_103/A 0.00fF
C9091 NOR2X1_LOC_145/Y NAND2X1_LOC_93/B 0.06fF
C9092 INVX1_LOC_27/A INVX1_LOC_63/Y 0.17fF
C9093 D_INPUT_4 NAND2X1_LOC_430/B 0.01fF
C9094 NOR2X1_LOC_91/A NAND2X1_LOC_854/B 0.68fF
C9095 INVX1_LOC_278/A NOR2X1_LOC_78/B 0.63fF
C9096 INVX1_LOC_36/A NOR2X1_LOC_590/A 0.10fF
C9097 INVX1_LOC_103/A NOR2X1_LOC_759/Y 0.21fF
C9098 NAND2X1_LOC_190/Y NOR2X1_LOC_303/Y 0.01fF
C9099 NAND2X1_LOC_391/Y NAND2X1_LOC_564/a_36_24# 0.00fF
C9100 NAND2X1_LOC_198/B INVX1_LOC_161/Y 0.10fF
C9101 NOR2X1_LOC_537/Y INVX1_LOC_138/Y 0.03fF
C9102 INVX1_LOC_202/A INVX1_LOC_103/A 0.00fF
C9103 INVX1_LOC_237/Y NOR2X1_LOC_92/Y 0.01fF
C9104 NOR2X1_LOC_246/A NOR2X1_LOC_301/A 0.07fF
C9105 NOR2X1_LOC_88/Y INVX1_LOC_46/A 0.03fF
C9106 NOR2X1_LOC_145/Y NAND2X1_LOC_425/Y 0.03fF
C9107 NOR2X1_LOC_164/Y INVX1_LOC_84/A 0.31fF
C9108 INVX1_LOC_34/A INVX1_LOC_48/Y 0.07fF
C9109 INVX1_LOC_227/A INVX1_LOC_270/A 0.10fF
C9110 INVX1_LOC_201/Y INVX1_LOC_163/A 0.11fF
C9111 INVX1_LOC_136/A NAND2X1_LOC_500/Y 0.02fF
C9112 NOR2X1_LOC_215/A NOR2X1_LOC_52/B 0.01fF
C9113 INVX1_LOC_11/A NOR2X1_LOC_152/Y 0.08fF
C9114 NOR2X1_LOC_598/B NOR2X1_LOC_687/Y 0.24fF
C9115 NOR2X1_LOC_78/A NOR2X1_LOC_777/B 0.06fF
C9116 NOR2X1_LOC_778/B INVX1_LOC_5/A 0.03fF
C9117 INVX1_LOC_11/A INVX1_LOC_113/Y 0.04fF
C9118 INPUT_1 INVX1_LOC_26/A 0.05fF
C9119 NOR2X1_LOC_614/a_36_216# NOR2X1_LOC_516/B 0.14fF
C9120 INVX1_LOC_136/Y INVX1_LOC_76/A 0.01fF
C9121 NAND2X1_LOC_190/Y NOR2X1_LOC_254/Y 0.13fF
C9122 INVX1_LOC_36/A NAND2X1_LOC_589/a_36_24# 0.01fF
C9123 NAND2X1_LOC_149/Y INVX1_LOC_266/Y 0.34fF
C9124 NOR2X1_LOC_433/A NOR2X1_LOC_503/Y 0.01fF
C9125 VDD NOR2X1_LOC_127/Y 0.39fF
C9126 NOR2X1_LOC_790/B INVX1_LOC_220/Y 0.04fF
C9127 NAND2X1_LOC_347/B NOR2X1_LOC_315/Y 0.17fF
C9128 NOR2X1_LOC_272/Y NAND2X1_LOC_338/B 0.01fF
C9129 NOR2X1_LOC_635/A INVX1_LOC_1/A 0.04fF
C9130 INVX1_LOC_84/A INVX1_LOC_46/A 0.17fF
C9131 INVX1_LOC_129/Y NAND2X1_LOC_572/B 0.21fF
C9132 NAND2X1_LOC_465/A INVX1_LOC_19/A 0.01fF
C9133 NAND2X1_LOC_364/A INVX1_LOC_72/A 0.03fF
C9134 INVX1_LOC_40/A NOR2X1_LOC_649/Y 0.22fF
C9135 NOR2X1_LOC_296/a_36_216# INVX1_LOC_8/A 0.01fF
C9136 NOR2X1_LOC_641/B INVX1_LOC_24/A 0.03fF
C9137 NAND2X1_LOC_638/Y NOR2X1_LOC_635/B 0.14fF
C9138 INVX1_LOC_292/A NOR2X1_LOC_550/B 0.01fF
C9139 NOR2X1_LOC_123/B INVX1_LOC_29/Y 0.01fF
C9140 NOR2X1_LOC_191/A NAND2X1_LOC_474/Y 0.02fF
C9141 INVX1_LOC_1/A NAND2X1_LOC_141/A 0.39fF
C9142 INVX1_LOC_10/A NOR2X1_LOC_678/A 0.01fF
C9143 NOR2X1_LOC_155/A INVX1_LOC_9/A 0.06fF
C9144 INVX1_LOC_213/Y NOR2X1_LOC_739/Y 0.01fF
C9145 INVX1_LOC_1/A INVX1_LOC_96/Y 0.14fF
C9146 INVX1_LOC_161/A INVX1_LOC_231/Y 0.01fF
C9147 INVX1_LOC_108/Y INVX1_LOC_83/A 0.56fF
C9148 NAND2X1_LOC_59/B INVX1_LOC_174/A 0.27fF
C9149 NOR2X1_LOC_186/Y INVX1_LOC_22/A 0.00fF
C9150 NOR2X1_LOC_751/Y INVX1_LOC_24/A 0.03fF
C9151 NAND2X1_LOC_17/a_36_24# NAND2X1_LOC_36/A 0.02fF
C9152 NAND2X1_LOC_705/Y NOR2X1_LOC_526/Y 0.06fF
C9153 NOR2X1_LOC_82/A NOR2X1_LOC_278/A 0.03fF
C9154 NOR2X1_LOC_103/Y INVX1_LOC_60/Y 0.16fF
C9155 NOR2X1_LOC_730/B INVX1_LOC_274/Y 0.29fF
C9156 NAND2X1_LOC_579/A NAND2X1_LOC_374/Y 0.10fF
C9157 INVX1_LOC_38/A NOR2X1_LOC_697/Y 0.03fF
C9158 NOR2X1_LOC_255/Y INPUT_1 0.01fF
C9159 INVX1_LOC_74/A NOR2X1_LOC_847/A 0.02fF
C9160 NOR2X1_LOC_311/Y INVX1_LOC_15/A 0.03fF
C9161 NOR2X1_LOC_825/Y NOR2X1_LOC_671/Y 0.03fF
C9162 NAND2X1_LOC_297/a_36_24# INVX1_LOC_3/A 0.00fF
C9163 NOR2X1_LOC_318/B NAND2X1_LOC_647/B 0.01fF
C9164 NOR2X1_LOC_865/A NOR2X1_LOC_814/A 0.03fF
C9165 NOR2X1_LOC_223/B INVX1_LOC_83/A 0.06fF
C9166 NAND2X1_LOC_573/Y INVX1_LOC_22/A 0.02fF
C9167 NOR2X1_LOC_590/A NOR2X1_LOC_309/Y 0.01fF
C9168 NOR2X1_LOC_717/Y INVX1_LOC_153/Y 0.01fF
C9169 INVX1_LOC_37/A INPUT_7 0.51fF
C9170 INVX1_LOC_73/A INVX1_LOC_57/A 0.03fF
C9171 INVX1_LOC_77/Y NOR2X1_LOC_11/Y 0.08fF
C9172 NAND2X1_LOC_577/A NOR2X1_LOC_514/Y 0.06fF
C9173 NOR2X1_LOC_841/A NOR2X1_LOC_743/Y 0.01fF
C9174 NAND2X1_LOC_563/Y NOR2X1_LOC_514/A 0.06fF
C9175 INVX1_LOC_286/Y NOR2X1_LOC_591/a_36_216# 0.01fF
C9176 NAND2X1_LOC_724/A INVX1_LOC_22/A 0.28fF
C9177 NAND2X1_LOC_207/B INVX1_LOC_117/A 0.02fF
C9178 INVX1_LOC_13/Y INVX1_LOC_171/A 0.06fF
C9179 INVX1_LOC_2/A INVX1_LOC_141/A 0.02fF
C9180 NAND2X1_LOC_208/B NOR2X1_LOC_84/Y 0.03fF
C9181 NOR2X1_LOC_122/A NOR2X1_LOC_665/A 0.08fF
C9182 NOR2X1_LOC_307/A NOR2X1_LOC_731/Y 0.01fF
C9183 INVX1_LOC_225/A NOR2X1_LOC_274/B 0.02fF
C9184 INVX1_LOC_88/A NOR2X1_LOC_589/A 0.03fF
C9185 INVX1_LOC_17/A INVX1_LOC_13/A 0.02fF
C9186 NOR2X1_LOC_433/A NOR2X1_LOC_152/Y 0.67fF
C9187 INVX1_LOC_78/A NOR2X1_LOC_601/Y 0.01fF
C9188 INVX1_LOC_46/A INVX1_LOC_15/A 0.52fF
C9189 INVX1_LOC_199/A INVX1_LOC_78/A 0.00fF
C9190 NOR2X1_LOC_337/Y NOR2X1_LOC_383/B 0.02fF
C9191 NOR2X1_LOC_641/B INVX1_LOC_143/A 0.13fF
C9192 NAND2X1_LOC_577/A NAND2X1_LOC_549/B 0.08fF
C9193 INVX1_LOC_78/Y NOR2X1_LOC_748/A 0.05fF
C9194 NOR2X1_LOC_78/A NOR2X1_LOC_843/B 0.03fF
C9195 NAND2X1_LOC_7/Y NOR2X1_LOC_716/B 0.09fF
C9196 INVX1_LOC_41/A NOR2X1_LOC_274/Y -0.00fF
C9197 INVX1_LOC_249/A INVX1_LOC_63/Y 0.18fF
C9198 NOR2X1_LOC_251/a_36_216# INVX1_LOC_313/A -0.00fF
C9199 NOR2X1_LOC_45/Y INVX1_LOC_22/A 0.00fF
C9200 INVX1_LOC_227/Y INVX1_LOC_177/A 0.01fF
C9201 NOR2X1_LOC_593/Y INVX1_LOC_113/Y 0.00fF
C9202 INVX1_LOC_50/A NOR2X1_LOC_45/B 0.13fF
C9203 NOR2X1_LOC_751/Y INVX1_LOC_143/A 0.01fF
C9204 NAND2X1_LOC_364/Y INVX1_LOC_33/A 0.03fF
C9205 NOR2X1_LOC_820/A NOR2X1_LOC_818/Y 0.03fF
C9206 NAND2X1_LOC_364/A NOR2X1_LOC_537/Y 0.07fF
C9207 INVX1_LOC_49/A INVX1_LOC_103/Y 0.00fF
C9208 INVX1_LOC_285/A NOR2X1_LOC_654/a_36_216# 0.01fF
C9209 INVX1_LOC_13/A NAND2X1_LOC_555/Y 0.08fF
C9210 INVX1_LOC_201/Y INVX1_LOC_203/Y 0.01fF
C9211 INVX1_LOC_34/A INVX1_LOC_231/Y 0.03fF
C9212 INVX1_LOC_17/A NOR2X1_LOC_246/A 0.07fF
C9213 NOR2X1_LOC_52/B NOR2X1_LOC_152/Y 0.14fF
C9214 INVX1_LOC_285/A INVX1_LOC_63/A 0.14fF
C9215 INVX1_LOC_136/A INVX1_LOC_278/Y 0.07fF
C9216 NOR2X1_LOC_68/A NOR2X1_LOC_769/a_36_216# 0.00fF
C9217 NOR2X1_LOC_78/B NOR2X1_LOC_168/Y 0.00fF
C9218 NAND2X1_LOC_555/Y NAND2X1_LOC_14/a_36_24# 0.00fF
C9219 NOR2X1_LOC_32/B INVX1_LOC_91/A 0.16fF
C9220 INVX1_LOC_50/A INVX1_LOC_247/A 0.06fF
C9221 NOR2X1_LOC_89/A NAND2X1_LOC_802/Y 0.59fF
C9222 NOR2X1_LOC_814/A INVX1_LOC_63/A 0.29fF
C9223 NAND2X1_LOC_794/B INPUT_0 0.00fF
C9224 NAND2X1_LOC_736/Y NAND2X1_LOC_736/B 0.01fF
C9225 NOR2X1_LOC_224/Y NOR2X1_LOC_45/B 0.01fF
C9226 INVX1_LOC_45/A INVX1_LOC_101/A 0.03fF
C9227 INVX1_LOC_230/Y D_INPUT_0 0.42fF
C9228 INVX1_LOC_256/A NOR2X1_LOC_246/a_36_216# 0.01fF
C9229 NAND2X1_LOC_736/Y GATE_811 0.03fF
C9230 NOR2X1_LOC_639/B INVX1_LOC_91/A 0.03fF
C9231 NOR2X1_LOC_91/Y INVX1_LOC_25/Y 0.08fF
C9232 INVX1_LOC_174/A NAND2X1_LOC_1/a_36_24# 0.01fF
C9233 INVX1_LOC_89/A NAND2X1_LOC_114/B 0.08fF
C9234 INVX1_LOC_72/Y INVX1_LOC_16/A 0.00fF
C9235 INVX1_LOC_2/A NOR2X1_LOC_214/a_36_216# 0.00fF
C9236 INVX1_LOC_268/A NOR2X1_LOC_68/A 0.02fF
C9237 INVX1_LOC_64/A NOR2X1_LOC_139/Y 0.07fF
C9238 NAND2X1_LOC_141/Y NOR2X1_LOC_128/A 0.03fF
C9239 INVX1_LOC_64/A NAND2X1_LOC_655/A 0.01fF
C9240 NOR2X1_LOC_205/Y NOR2X1_LOC_736/a_36_216# 0.00fF
C9241 NOR2X1_LOC_220/A NOR2X1_LOC_303/Y 0.12fF
C9242 NOR2X1_LOC_773/Y INVX1_LOC_314/Y 0.01fF
C9243 NAND2X1_LOC_725/B INVX1_LOC_282/A 0.07fF
C9244 INPUT_3 INVX1_LOC_20/Y 0.02fF
C9245 INVX1_LOC_34/A NOR2X1_LOC_84/Y 0.01fF
C9246 VDD NOR2X1_LOC_383/B 2.10fF
C9247 INVX1_LOC_5/A NOR2X1_LOC_557/A 4.37fF
C9248 INVX1_LOC_48/Y INPUT_0 0.07fF
C9249 NOR2X1_LOC_471/Y INVX1_LOC_55/Y 0.04fF
C9250 NOR2X1_LOC_413/Y NOR2X1_LOC_399/A 0.02fF
C9251 INVX1_LOC_36/A NOR2X1_LOC_763/Y 0.02fF
C9252 INVX1_LOC_45/A NOR2X1_LOC_355/A 0.64fF
C9253 INVX1_LOC_278/A NOR2X1_LOC_368/Y 0.02fF
C9254 INVX1_LOC_230/Y NAND2X1_LOC_665/a_36_24# 0.00fF
C9255 NOR2X1_LOC_351/Y INVX1_LOC_128/Y 0.12fF
C9256 NOR2X1_LOC_716/B NAND2X1_LOC_318/a_36_24# 0.07fF
C9257 INVX1_LOC_34/A NOR2X1_LOC_482/Y 0.15fF
C9258 NOR2X1_LOC_15/Y NOR2X1_LOC_188/A 3.30fF
C9259 NAND2X1_LOC_444/B INVX1_LOC_54/A 0.01fF
C9260 INVX1_LOC_84/A NOR2X1_LOC_671/Y 0.03fF
C9261 NOR2X1_LOC_295/Y INVX1_LOC_54/Y 0.02fF
C9262 NOR2X1_LOC_818/Y INVX1_LOC_315/A 0.53fF
C9263 INVX1_LOC_59/Y NOR2X1_LOC_660/Y 0.01fF
C9264 NOR2X1_LOC_334/Y INVX1_LOC_54/A 0.07fF
C9265 NOR2X1_LOC_488/Y NOR2X1_LOC_237/Y 0.20fF
C9266 NAND2X1_LOC_738/B VDD 0.51fF
C9267 INVX1_LOC_64/A NAND2X1_LOC_468/B 0.09fF
C9268 INVX1_LOC_223/A NAND2X1_LOC_140/A 0.00fF
C9269 NOR2X1_LOC_78/Y NOR2X1_LOC_38/B 0.48fF
C9270 NOR2X1_LOC_690/A NOR2X1_LOC_526/Y 0.12fF
C9271 NAND2X1_LOC_738/B NAND2X1_LOC_800/A 0.00fF
C9272 NAND2X1_LOC_35/Y NOR2X1_LOC_824/Y 0.03fF
C9273 INVX1_LOC_135/A NOR2X1_LOC_791/B 0.03fF
C9274 INVX1_LOC_101/A INVX1_LOC_71/A 0.00fF
C9275 INVX1_LOC_132/A INVX1_LOC_22/A 0.02fF
C9276 INVX1_LOC_1/A NOR2X1_LOC_733/Y 0.02fF
C9277 NAND2X1_LOC_392/A NOR2X1_LOC_716/B 0.01fF
C9278 INVX1_LOC_50/A INVX1_LOC_281/A 0.01fF
C9279 INVX1_LOC_11/A INVX1_LOC_158/Y 0.01fF
C9280 NAND2X1_LOC_358/B INVX1_LOC_176/A 0.01fF
C9281 INVX1_LOC_278/A INVX1_LOC_46/A 0.08fF
C9282 INVX1_LOC_26/A INVX1_LOC_118/A 0.08fF
C9283 INVX1_LOC_177/Y INVX1_LOC_313/A 1.04fF
C9284 INVX1_LOC_124/Y NOR2X1_LOC_153/a_36_216# 0.00fF
C9285 INVX1_LOC_2/A INVX1_LOC_149/A 0.12fF
C9286 NOR2X1_LOC_155/A INVX1_LOC_274/Y 0.21fF
C9287 NAND2X1_LOC_639/A NOR2X1_LOC_452/A 0.04fF
C9288 INVX1_LOC_111/Y INVX1_LOC_177/A 0.00fF
C9289 NOR2X1_LOC_541/a_36_216# NOR2X1_LOC_541/Y 0.02fF
C9290 NOR2X1_LOC_298/Y NAND2X1_LOC_863/Y 0.04fF
C9291 NAND2X1_LOC_35/Y INVX1_LOC_76/A 0.14fF
C9292 INVX1_LOC_18/Y NOR2X1_LOC_640/Y 0.06fF
C9293 NOR2X1_LOC_254/A NOR2X1_LOC_74/A 0.10fF
C9294 INVX1_LOC_207/A NAND2X1_LOC_735/B 0.05fF
C9295 NOR2X1_LOC_351/Y NAND2X1_LOC_424/a_36_24# 0.00fF
C9296 INVX1_LOC_221/A NAND2X1_LOC_840/B 0.20fF
C9297 INVX1_LOC_24/A NOR2X1_LOC_71/Y 0.17fF
C9298 NAND2X1_LOC_811/Y INVX1_LOC_16/A 3.27fF
C9299 NOR2X1_LOC_590/A NOR2X1_LOC_208/A 0.03fF
C9300 NOR2X1_LOC_355/A INVX1_LOC_71/A 0.07fF
C9301 INVX1_LOC_34/A INVX1_LOC_290/A 0.03fF
C9302 INVX1_LOC_13/Y INVX1_LOC_20/A 0.06fF
C9303 INVX1_LOC_89/A NOR2X1_LOC_546/B 0.01fF
C9304 NOR2X1_LOC_570/B NOR2X1_LOC_569/Y 0.01fF
C9305 NOR2X1_LOC_335/A INVX1_LOC_10/A 0.01fF
C9306 NOR2X1_LOC_66/Y INVX1_LOC_4/A 0.07fF
C9307 NOR2X1_LOC_331/B INVX1_LOC_29/Y 0.01fF
C9308 INVX1_LOC_32/A NOR2X1_LOC_257/Y 0.04fF
C9309 NOR2X1_LOC_220/A INVX1_LOC_54/Y 0.34fF
C9310 NOR2X1_LOC_52/B NAND2X1_LOC_859/B 0.23fF
C9311 INVX1_LOC_290/Y INVX1_LOC_29/A 0.07fF
C9312 NAND2X1_LOC_564/A INVX1_LOC_118/A 0.02fF
C9313 NOR2X1_LOC_644/A INVX1_LOC_24/A 0.03fF
C9314 INVX1_LOC_303/A INVX1_LOC_171/A 0.02fF
C9315 NOR2X1_LOC_757/a_36_216# NOR2X1_LOC_757/Y 0.01fF
C9316 INVX1_LOC_16/A INVX1_LOC_266/Y 0.03fF
C9317 NAND2X1_LOC_21/Y INVX1_LOC_83/A 0.56fF
C9318 NAND2X1_LOC_156/B INVX1_LOC_63/Y 0.00fF
C9319 INVX1_LOC_45/A NOR2X1_LOC_541/a_36_216# 0.00fF
C9320 NOR2X1_LOC_721/B NOR2X1_LOC_38/B 0.03fF
C9321 NOR2X1_LOC_598/B INVX1_LOC_9/A 0.19fF
C9322 NAND2X1_LOC_227/Y NOR2X1_LOC_45/B 0.18fF
C9323 INVX1_LOC_89/A INVX1_LOC_275/A 0.01fF
C9324 INVX1_LOC_206/A NOR2X1_LOC_188/a_36_216# 0.00fF
C9325 NAND2X1_LOC_840/Y INVX1_LOC_18/A 0.01fF
C9326 NOR2X1_LOC_541/a_36_216# NOR2X1_LOC_568/A 0.00fF
C9327 INVX1_LOC_170/A INVX1_LOC_100/A 0.16fF
C9328 NAND2X1_LOC_254/Y INVX1_LOC_42/A 0.05fF
C9329 NAND2X1_LOC_178/a_36_24# INVX1_LOC_247/A 0.00fF
C9330 INVX1_LOC_88/A INVX1_LOC_147/Y 0.01fF
C9331 NAND2X1_LOC_231/Y INVX1_LOC_290/A 0.04fF
C9332 INVX1_LOC_45/Y NOR2X1_LOC_216/Y 0.02fF
C9333 NOR2X1_LOC_582/A VDD 0.24fF
C9334 NOR2X1_LOC_671/Y INVX1_LOC_15/A 0.03fF
C9335 D_INPUT_1 INVX1_LOC_92/A 0.06fF
C9336 INVX1_LOC_295/A INVX1_LOC_192/A 0.10fF
C9337 NAND2X1_LOC_852/Y INVX1_LOC_22/A 1.97fF
C9338 INVX1_LOC_94/Y INVX1_LOC_264/A 0.02fF
C9339 NAND2X1_LOC_223/B NOR2X1_LOC_814/A 0.15fF
C9340 INVX1_LOC_282/A INVX1_LOC_309/Y 0.01fF
C9341 INVX1_LOC_135/A NOR2X1_LOC_802/A 0.07fF
C9342 INVX1_LOC_206/A NOR2X1_LOC_370/a_36_216# 0.02fF
C9343 INVX1_LOC_177/Y INVX1_LOC_6/A 0.07fF
C9344 INVX1_LOC_104/A INVX1_LOC_313/A 0.02fF
C9345 NOR2X1_LOC_52/B NAND2X1_LOC_861/Y 0.08fF
C9346 NOR2X1_LOC_99/B NOR2X1_LOC_709/A 0.91fF
C9347 NOR2X1_LOC_804/B NOR2X1_LOC_703/A 0.01fF
C9348 NOR2X1_LOC_848/Y INVX1_LOC_2/Y 0.02fF
C9349 NOR2X1_LOC_226/A INVX1_LOC_164/A 0.06fF
C9350 NOR2X1_LOC_137/A INVX1_LOC_177/A 0.00fF
C9351 INVX1_LOC_28/A NAND2X1_LOC_811/Y 0.32fF
C9352 INVX1_LOC_225/Y NOR2X1_LOC_35/Y 0.03fF
C9353 NOR2X1_LOC_860/B NOR2X1_LOC_188/A 0.07fF
C9354 NOR2X1_LOC_215/Y INVX1_LOC_6/A 0.01fF
C9355 NAND2X1_LOC_63/Y NOR2X1_LOC_316/a_36_216# 0.00fF
C9356 NOR2X1_LOC_350/A INPUT_0 0.05fF
C9357 NAND2X1_LOC_45/Y INVX1_LOC_64/Y 0.27fF
C9358 INVX1_LOC_233/A NOR2X1_LOC_88/Y 0.07fF
C9359 INVX1_LOC_35/A NOR2X1_LOC_831/B 0.07fF
C9360 NOR2X1_LOC_189/A INPUT_0 0.02fF
C9361 NAND2X1_LOC_63/Y INVX1_LOC_26/A 0.05fF
C9362 NOR2X1_LOC_471/Y NOR2X1_LOC_357/Y 0.02fF
C9363 NOR2X1_LOC_68/A NOR2X1_LOC_746/a_36_216# 0.00fF
C9364 NAND2X1_LOC_656/A NAND2X1_LOC_473/a_36_24# 0.00fF
C9365 NOR2X1_LOC_6/a_36_216# INPUT_0 0.00fF
C9366 INVX1_LOC_72/A NOR2X1_LOC_405/A 0.03fF
C9367 INVX1_LOC_30/A NOR2X1_LOC_275/A 0.01fF
C9368 NOR2X1_LOC_266/a_36_216# INVX1_LOC_93/Y -0.01fF
C9369 NOR2X1_LOC_210/A NOR2X1_LOC_470/A 0.12fF
C9370 INVX1_LOC_58/A NOR2X1_LOC_605/A 0.01fF
C9371 INVX1_LOC_33/A NOR2X1_LOC_337/A 0.01fF
C9372 INVX1_LOC_234/A NAND2X1_LOC_848/a_36_24# 0.01fF
C9373 NAND2X1_LOC_9/Y INVX1_LOC_84/A 0.03fF
C9374 NAND2X1_LOC_205/A NAND2X1_LOC_773/B 0.10fF
C9375 NOR2X1_LOC_646/A INVX1_LOC_135/A 0.46fF
C9376 INVX1_LOC_26/A NAND2X1_LOC_455/B 0.72fF
C9377 INVX1_LOC_298/Y INVX1_LOC_290/Y 0.07fF
C9378 INVX1_LOC_233/A INVX1_LOC_84/A 0.19fF
C9379 NOR2X1_LOC_32/B INVX1_LOC_203/A 0.10fF
C9380 INVX1_LOC_136/A INVX1_LOC_59/Y 0.04fF
C9381 NOR2X1_LOC_250/a_36_216# INVX1_LOC_38/A 0.00fF
C9382 NOR2X1_LOC_554/B INVX1_LOC_74/A 0.02fF
C9383 INVX1_LOC_130/Y NAND2X1_LOC_468/B 0.00fF
C9384 NOR2X1_LOC_759/Y NOR2X1_LOC_141/a_36_216# 0.00fF
C9385 INVX1_LOC_89/A NOR2X1_LOC_789/A 0.04fF
C9386 INVX1_LOC_277/Y VDD -0.00fF
C9387 NOR2X1_LOC_34/B NAND2X1_LOC_574/A 0.02fF
C9388 NAND2X1_LOC_597/a_36_24# NAND2X1_LOC_472/Y 0.00fF
C9389 INVX1_LOC_57/Y VDD 1.94fF
C9390 INPUT_0 NOR2X1_LOC_84/Y 0.11fF
C9391 INVX1_LOC_230/Y NAND2X1_LOC_848/A 0.00fF
C9392 INVX1_LOC_45/A NOR2X1_LOC_111/A 0.22fF
C9393 NOR2X1_LOC_103/Y INVX1_LOC_127/A 0.02fF
C9394 INVX1_LOC_1/Y INVX1_LOC_87/Y 0.00fF
C9395 INVX1_LOC_104/A INVX1_LOC_6/A 0.08fF
C9396 NAND2X1_LOC_703/Y NOR2X1_LOC_88/Y 0.07fF
C9397 NOR2X1_LOC_510/Y NOR2X1_LOC_127/Y 0.08fF
C9398 INVX1_LOC_2/A NOR2X1_LOC_313/Y 0.00fF
C9399 NOR2X1_LOC_577/Y NAND2X1_LOC_642/Y 0.00fF
C9400 NOR2X1_LOC_751/A INVX1_LOC_143/A 0.10fF
C9401 NOR2X1_LOC_798/A INVX1_LOC_84/A 0.07fF
C9402 INPUT_0 INVX1_LOC_216/A 0.07fF
C9403 NOR2X1_LOC_590/A NOR2X1_LOC_865/A 0.01fF
C9404 INVX1_LOC_5/A NAND2X1_LOC_625/a_36_24# 0.00fF
C9405 NOR2X1_LOC_577/Y NAND2X1_LOC_643/a_36_24# 0.00fF
C9406 INVX1_LOC_27/A INVX1_LOC_27/Y 0.10fF
C9407 NAND2X1_LOC_454/Y INVX1_LOC_271/Y 0.87fF
C9408 NOR2X1_LOC_71/Y NOR2X1_LOC_130/A 0.07fF
C9409 INVX1_LOC_12/A NOR2X1_LOC_678/A 0.03fF
C9410 INVX1_LOC_199/A INVX1_LOC_113/Y 0.05fF
C9411 INVX1_LOC_11/A INVX1_LOC_291/A 0.09fF
C9412 INVX1_LOC_26/Y NAND2X1_LOC_278/a_36_24# 0.00fF
C9413 INVX1_LOC_164/A INPUT_1 0.06fF
C9414 NOR2X1_LOC_480/A VDD 0.12fF
C9415 NOR2X1_LOC_512/Y VDD 0.12fF
C9416 NAND2X1_LOC_223/A NAND2X1_LOC_221/a_36_24# 0.02fF
C9417 INVX1_LOC_141/A INVX1_LOC_118/A 0.04fF
C9418 NAND2X1_LOC_84/Y NAND2X1_LOC_267/B 0.03fF
C9419 INVX1_LOC_241/A INVX1_LOC_282/A 0.06fF
C9420 INVX1_LOC_18/A NOR2X1_LOC_60/Y 0.02fF
C9421 INVX1_LOC_42/Y INVX1_LOC_16/A 0.03fF
C9422 INVX1_LOC_89/A INVX1_LOC_132/Y 0.01fF
C9423 INVX1_LOC_68/Y NOR2X1_LOC_199/a_36_216# 0.00fF
C9424 NOR2X1_LOC_78/B INVX1_LOC_123/A 0.06fF
C9425 INVX1_LOC_71/A NOR2X1_LOC_111/A 0.18fF
C9426 NAND2X1_LOC_798/a_36_24# NAND2X1_LOC_453/A 0.00fF
C9427 NOR2X1_LOC_543/A INVX1_LOC_75/A 0.16fF
C9428 NAND2X1_LOC_632/B VDD 0.07fF
C9429 NOR2X1_LOC_791/B INVX1_LOC_280/A 0.58fF
C9430 INVX1_LOC_230/Y INVX1_LOC_46/Y 0.51fF
C9431 NOR2X1_LOC_361/B NOR2X1_LOC_127/Y 0.26fF
C9432 NAND2X1_LOC_342/Y NOR2X1_LOC_318/B 0.03fF
C9433 NAND2X1_LOC_9/Y INVX1_LOC_15/A 0.07fF
C9434 NAND2X1_LOC_149/Y INVX1_LOC_19/A 0.07fF
C9435 INVX1_LOC_90/A NOR2X1_LOC_770/Y 0.02fF
C9436 NOR2X1_LOC_78/A NOR2X1_LOC_709/a_36_216# 0.01fF
C9437 NOR2X1_LOC_360/Y INVX1_LOC_230/A 0.02fF
C9438 NOR2X1_LOC_426/Y NOR2X1_LOC_51/A 0.81fF
C9439 INVX1_LOC_233/A INVX1_LOC_15/A 0.49fF
C9440 INVX1_LOC_135/A INVX1_LOC_82/Y 0.04fF
C9441 INVX1_LOC_48/Y NOR2X1_LOC_84/B 0.00fF
C9442 NOR2X1_LOC_792/a_36_216# NAND2X1_LOC_81/B 0.00fF
C9443 NOR2X1_LOC_298/Y INVX1_LOC_282/A 0.05fF
C9444 NOR2X1_LOC_561/Y INVX1_LOC_144/A 1.64fF
C9445 NAND2X1_LOC_303/B INVX1_LOC_140/A 0.07fF
C9446 NOR2X1_LOC_454/Y INVX1_LOC_29/A 0.11fF
C9447 NOR2X1_LOC_25/Y INVX1_LOC_296/A 0.08fF
C9448 D_INPUT_1 NAND2X1_LOC_247/a_36_24# 0.00fF
C9449 NOR2X1_LOC_716/B INVX1_LOC_129/Y 0.01fF
C9450 INVX1_LOC_17/A NAND2X1_LOC_489/Y 0.02fF
C9451 NOR2X1_LOC_147/B INVX1_LOC_37/A 0.01fF
C9452 NOR2X1_LOC_598/B INVX1_LOC_274/Y 0.51fF
C9453 NOR2X1_LOC_346/B NAND2X1_LOC_642/Y 0.01fF
C9454 INVX1_LOC_168/A INVX1_LOC_20/A 0.08fF
C9455 NOR2X1_LOC_753/Y NOR2X1_LOC_536/A 0.01fF
C9456 NOR2X1_LOC_772/B INVX1_LOC_4/A 0.10fF
C9457 NOR2X1_LOC_570/B NAND2X1_LOC_472/Y 0.02fF
C9458 NOR2X1_LOC_489/B INVX1_LOC_4/Y 0.04fF
C9459 NOR2X1_LOC_751/Y NOR2X1_LOC_197/B 0.30fF
C9460 NOR2X1_LOC_264/Y INVX1_LOC_117/A 0.02fF
C9461 NOR2X1_LOC_798/A INVX1_LOC_15/A 0.03fF
C9462 INVX1_LOC_103/A NAND2X1_LOC_74/B 0.03fF
C9463 NAND2X1_LOC_325/Y NOR2X1_LOC_536/A 0.00fF
C9464 INVX1_LOC_24/A NAND2X1_LOC_243/Y 0.00fF
C9465 NOR2X1_LOC_235/a_36_216# INVX1_LOC_284/A 0.00fF
C9466 INVX1_LOC_22/A NAND2X1_LOC_642/Y 0.15fF
C9467 INVX1_LOC_13/Y INVX1_LOC_4/A 5.52fF
C9468 NAND2X1_LOC_539/a_36_24# INVX1_LOC_49/Y 0.00fF
C9469 NOR2X1_LOC_590/A INVX1_LOC_63/A 0.11fF
C9470 INVX1_LOC_305/A NOR2X1_LOC_445/B 0.09fF
C9471 NOR2X1_LOC_537/Y NOR2X1_LOC_857/A 0.12fF
C9472 INVX1_LOC_308/Y NAND2X1_LOC_807/B 0.14fF
C9473 INVX1_LOC_209/Y INVX1_LOC_54/A 0.07fF
C9474 NOR2X1_LOC_788/B INVX1_LOC_69/Y 0.02fF
C9475 NAND2X1_LOC_323/B NOR2X1_LOC_857/A 0.07fF
C9476 NOR2X1_LOC_124/B INVX1_LOC_280/A 0.01fF
C9477 INVX1_LOC_89/A INVX1_LOC_78/Y 0.03fF
C9478 NOR2X1_LOC_433/A INVX1_LOC_291/A 0.01fF
C9479 NOR2X1_LOC_652/Y NAND2X1_LOC_247/a_36_24# 0.01fF
C9480 NOR2X1_LOC_38/B NAND2X1_LOC_473/A 0.02fF
C9481 NAND2X1_LOC_303/Y D_INPUT_5 0.01fF
C9482 NOR2X1_LOC_433/A NAND2X1_LOC_802/Y 0.02fF
C9483 NOR2X1_LOC_794/B INVX1_LOC_99/A 0.04fF
C9484 NOR2X1_LOC_816/a_36_216# INVX1_LOC_78/A 0.00fF
C9485 NOR2X1_LOC_322/Y NOR2X1_LOC_74/A 0.10fF
C9486 NOR2X1_LOC_613/a_36_216# INVX1_LOC_78/A 0.00fF
C9487 INVX1_LOC_283/Y INVX1_LOC_179/A -0.00fF
C9488 NOR2X1_LOC_361/Y NOR2X1_LOC_331/B 0.04fF
C9489 NAND2X1_LOC_392/A NAND2X1_LOC_633/Y 0.01fF
C9490 D_INPUT_1 INVX1_LOC_53/A 0.08fF
C9491 NAND2X1_LOC_170/A VDD 0.25fF
C9492 NOR2X1_LOC_355/B NOR2X1_LOC_356/A 0.02fF
C9493 INVX1_LOC_17/A INVX1_LOC_32/A 0.10fF
C9494 INVX1_LOC_50/A NOR2X1_LOC_53/Y 0.20fF
C9495 NOR2X1_LOC_67/A NOR2X1_LOC_536/A 0.23fF
C9496 NOR2X1_LOC_532/Y NOR2X1_LOC_552/A 0.03fF
C9497 NOR2X1_LOC_34/A NOR2X1_LOC_34/Y 0.00fF
C9498 INVX1_LOC_39/A INVX1_LOC_26/A 0.02fF
C9499 NOR2X1_LOC_137/A NOR2X1_LOC_137/B 0.00fF
C9500 NAND2X1_LOC_326/A INVX1_LOC_273/A 0.04fF
C9501 INVX1_LOC_14/A INVX1_LOC_4/Y 2.10fF
C9502 INVX1_LOC_62/Y NOR2X1_LOC_721/B 0.09fF
C9503 NAND2X1_LOC_9/Y INVX1_LOC_278/A 0.07fF
C9504 INVX1_LOC_313/Y NOR2X1_LOC_405/A 0.00fF
C9505 NOR2X1_LOC_52/B INVX1_LOC_291/A 0.14fF
C9506 INVX1_LOC_104/A INVX1_LOC_131/Y 0.10fF
C9507 INVX1_LOC_17/A NOR2X1_LOC_329/Y 0.07fF
C9508 NOR2X1_LOC_471/Y INVX1_LOC_32/A 0.03fF
C9509 INVX1_LOC_93/Y INVX1_LOC_87/Y 0.02fF
C9510 INVX1_LOC_233/A INVX1_LOC_278/A 0.44fF
C9511 NAND2X1_LOC_99/Y INVX1_LOC_27/Y 0.01fF
C9512 INVX1_LOC_90/A NOR2X1_LOC_631/B 0.72fF
C9513 INVX1_LOC_289/A INVX1_LOC_38/A 0.01fF
C9514 NOR2X1_LOC_478/a_36_216# INVX1_LOC_37/A 0.00fF
C9515 INVX1_LOC_302/A INVX1_LOC_91/A 0.01fF
C9516 INVX1_LOC_72/A INVX1_LOC_109/Y 0.07fF
C9517 INVX1_LOC_135/A INVX1_LOC_2/Y 1.59fF
C9518 NOR2X1_LOC_272/Y INVX1_LOC_224/Y 0.10fF
C9519 NOR2X1_LOC_78/A INVX1_LOC_31/Y 0.23fF
C9520 NAND2X1_LOC_555/Y INVX1_LOC_32/A 0.07fF
C9521 NOR2X1_LOC_646/A INVX1_LOC_280/A 0.24fF
C9522 INVX1_LOC_160/Y INVX1_LOC_117/A 0.05fF
C9523 NOR2X1_LOC_91/A NOR2X1_LOC_92/Y 0.10fF
C9524 NOR2X1_LOC_411/A NAND2X1_LOC_35/Y 0.02fF
C9525 NOR2X1_LOC_355/B NOR2X1_LOC_74/A 0.00fF
C9526 INVX1_LOC_166/A INVX1_LOC_235/Y 0.65fF
C9527 INVX1_LOC_17/A NAND2X1_LOC_175/Y 0.08fF
C9528 NOR2X1_LOC_318/B INVX1_LOC_67/Y 0.01fF
C9529 INVX1_LOC_53/A NOR2X1_LOC_652/Y 0.17fF
C9530 INVX1_LOC_39/A NOR2X1_LOC_255/Y 0.01fF
C9531 NOR2X1_LOC_828/B NOR2X1_LOC_209/A 0.01fF
C9532 NOR2X1_LOC_2/Y NOR2X1_LOC_588/A 0.02fF
C9533 INVX1_LOC_50/Y INVX1_LOC_58/Y 0.08fF
C9534 NAND2X1_LOC_149/B INVX1_LOC_193/A 0.01fF
C9535 NOR2X1_LOC_134/Y NAND2X1_LOC_471/Y 0.01fF
C9536 NOR2X1_LOC_570/A INVX1_LOC_9/A 0.02fF
C9537 INVX1_LOC_90/A INVX1_LOC_37/A 4.82fF
C9538 INVX1_LOC_77/A INVX1_LOC_29/A 0.91fF
C9539 NOR2X1_LOC_440/Y NOR2X1_LOC_186/a_36_216# 0.00fF
C9540 NOR2X1_LOC_441/Y NAND2X1_LOC_444/B 0.17fF
C9541 NOR2X1_LOC_374/A NOR2X1_LOC_777/B 0.06fF
C9542 INVX1_LOC_126/A INVX1_LOC_102/Y 0.12fF
C9543 NOR2X1_LOC_92/Y INVX1_LOC_23/A 0.37fF
C9544 NOR2X1_LOC_441/Y NOR2X1_LOC_334/Y 0.03fF
C9545 NOR2X1_LOC_131/a_36_216# NOR2X1_LOC_155/A 0.00fF
C9546 NAND2X1_LOC_214/B INVX1_LOC_5/A 0.00fF
C9547 NAND2X1_LOC_354/a_36_24# INVX1_LOC_78/A 0.00fF
C9548 INVX1_LOC_2/Y NOR2X1_LOC_346/a_36_216# 0.00fF
C9549 INVX1_LOC_100/A NAND2X1_LOC_642/Y 0.03fF
C9550 NOR2X1_LOC_335/A INVX1_LOC_12/A 0.01fF
C9551 INVX1_LOC_24/Y INVX1_LOC_23/A 0.53fF
C9552 INVX1_LOC_314/Y INVX1_LOC_42/A 0.07fF
C9553 NOR2X1_LOC_6/B NAND2X1_LOC_219/B 0.21fF
C9554 NAND2X1_LOC_860/A NOR2X1_LOC_468/Y 0.09fF
C9555 NAND2X1_LOC_798/A NOR2X1_LOC_697/Y 0.01fF
C9556 NOR2X1_LOC_163/Y VDD 0.30fF
C9557 INVX1_LOC_266/A INVX1_LOC_58/Y 0.02fF
C9558 NOR2X1_LOC_368/A NAND2X1_LOC_455/a_36_24# 0.00fF
C9559 INVX1_LOC_27/A INVX1_LOC_5/A 0.24fF
C9560 NOR2X1_LOC_67/A INVX1_LOC_3/A 0.22fF
C9561 INVX1_LOC_221/A INVX1_LOC_49/Y 0.63fF
C9562 INVX1_LOC_144/A INVX1_LOC_76/A 0.18fF
C9563 NOR2X1_LOC_770/Y INVX1_LOC_38/A 0.00fF
C9564 NOR2X1_LOC_15/Y NOR2X1_LOC_129/a_36_216# 0.00fF
C9565 NOR2X1_LOC_84/Y NOR2X1_LOC_84/B 0.24fF
C9566 VDD NOR2X1_LOC_74/Y 0.12fF
C9567 NOR2X1_LOC_162/a_36_216# NAND2X1_LOC_425/Y 0.01fF
C9568 NOR2X1_LOC_209/Y INVX1_LOC_186/Y 0.00fF
C9569 NOR2X1_LOC_816/A INVX1_LOC_271/A 0.01fF
C9570 INVX1_LOC_5/A INVX1_LOC_237/A 0.21fF
C9571 NOR2X1_LOC_68/A INVX1_LOC_271/Y 0.19fF
C9572 NOR2X1_LOC_561/Y NOR2X1_LOC_155/A 0.09fF
C9573 NOR2X1_LOC_589/A INVX1_LOC_107/Y 0.04fF
C9574 INVX1_LOC_24/A INVX1_LOC_21/Y 0.05fF
C9575 NOR2X1_LOC_334/A INVX1_LOC_143/Y 0.02fF
C9576 NAND2X1_LOC_819/Y INVX1_LOC_63/A 0.08fF
C9577 NAND2X1_LOC_662/a_36_24# INVX1_LOC_117/Y 0.00fF
C9578 INVX1_LOC_208/A NAND2X1_LOC_475/Y 0.10fF
C9579 INVX1_LOC_64/A INVX1_LOC_88/A 0.19fF
C9580 INVX1_LOC_124/A INVX1_LOC_29/A 0.10fF
C9581 INVX1_LOC_1/Y INVX1_LOC_285/A 0.09fF
C9582 INVX1_LOC_160/A NOR2X1_LOC_324/A 0.01fF
C9583 INVX1_LOC_30/Y NAND2X1_LOC_572/B 0.04fF
C9584 NOR2X1_LOC_836/Y NOR2X1_LOC_836/A 0.02fF
C9585 NOR2X1_LOC_824/A INVX1_LOC_178/A 0.10fF
C9586 INVX1_LOC_303/A INVX1_LOC_4/A 0.07fF
C9587 INVX1_LOC_35/A D_GATE_741 0.02fF
C9588 NOR2X1_LOC_180/B INVX1_LOC_274/A 0.02fF
C9589 INVX1_LOC_1/Y NOR2X1_LOC_814/A 0.45fF
C9590 INVX1_LOC_135/A NOR2X1_LOC_608/Y 0.02fF
C9591 INVX1_LOC_90/A NOR2X1_LOC_743/Y 0.09fF
C9592 INVX1_LOC_86/A INVX1_LOC_117/A 0.02fF
C9593 INVX1_LOC_314/Y INVX1_LOC_78/A 0.07fF
C9594 NAND2X1_LOC_363/B NOR2X1_LOC_160/B 0.19fF
C9595 INPUT_1 NOR2X1_LOC_235/Y 0.07fF
C9596 NOR2X1_LOC_389/B NOR2X1_LOC_743/Y 0.00fF
C9597 INVX1_LOC_35/A NAND2X1_LOC_352/B 0.03fF
C9598 INVX1_LOC_24/A INVX1_LOC_16/Y 0.48fF
C9599 INVX1_LOC_16/A INVX1_LOC_19/A 0.13fF
C9600 NOR2X1_LOC_214/B INVX1_LOC_113/A 0.01fF
C9601 INVX1_LOC_16/A NOR2X1_LOC_11/Y 0.16fF
C9602 NOR2X1_LOC_644/A NOR2X1_LOC_197/B 0.03fF
C9603 NOR2X1_LOC_65/B NAND2X1_LOC_315/a_36_24# 0.00fF
C9604 INVX1_LOC_298/Y INVX1_LOC_77/A 0.02fF
C9605 NOR2X1_LOC_91/A NAND2X1_LOC_837/Y 0.05fF
C9606 NOR2X1_LOC_142/Y NOR2X1_LOC_334/Y 0.10fF
C9607 NOR2X1_LOC_272/Y NOR2X1_LOC_103/Y 0.10fF
C9608 NOR2X1_LOC_242/A NOR2X1_LOC_241/A 0.06fF
C9609 NOR2X1_LOC_368/A INVX1_LOC_118/A 0.51fF
C9610 NAND2X1_LOC_714/B NOR2X1_LOC_533/Y 0.06fF
C9611 NOR2X1_LOC_313/Y INVX1_LOC_118/A 0.02fF
C9612 NOR2X1_LOC_65/B INVX1_LOC_314/Y 0.10fF
C9613 NOR2X1_LOC_589/A INVX1_LOC_272/A 0.07fF
C9614 INVX1_LOC_245/A NOR2X1_LOC_89/A 0.01fF
C9615 INPUT_5 NOR2X1_LOC_36/B 0.34fF
C9616 INVX1_LOC_27/A NAND2X1_LOC_337/B 0.43fF
C9617 NOR2X1_LOC_791/Y NOR2X1_LOC_160/B 0.04fF
C9618 NOR2X1_LOC_778/A INVX1_LOC_53/A 0.24fF
C9619 INVX1_LOC_64/A NOR2X1_LOC_500/B 3.79fF
C9620 INVX1_LOC_24/A NAND2X1_LOC_205/A 0.03fF
C9621 INVX1_LOC_132/A NOR2X1_LOC_843/B 0.07fF
C9622 NOR2X1_LOC_632/Y NOR2X1_LOC_89/A 0.03fF
C9623 NOR2X1_LOC_703/B INVX1_LOC_292/Y -0.00fF
C9624 NOR2X1_LOC_231/a_36_216# INVX1_LOC_50/Y 0.12fF
C9625 NOR2X1_LOC_91/A INVX1_LOC_41/A 0.06fF
C9626 INVX1_LOC_41/A NOR2X1_LOC_668/Y 0.17fF
C9627 INVX1_LOC_111/Y INVX1_LOC_4/Y 0.02fF
C9628 NOR2X1_LOC_455/Y INVX1_LOC_94/A 0.01fF
C9629 INVX1_LOC_236/A INVX1_LOC_94/Y 0.03fF
C9630 INVX1_LOC_316/Y INVX1_LOC_3/Y 0.72fF
C9631 NOR2X1_LOC_793/Y NOR2X1_LOC_807/B 0.00fF
C9632 NOR2X1_LOC_620/Y INVX1_LOC_57/A 0.04fF
C9633 NOR2X1_LOC_655/B NOR2X1_LOC_334/Y 0.02fF
C9634 NAND2X1_LOC_117/a_36_24# NAND2X1_LOC_63/Y 0.00fF
C9635 NOR2X1_LOC_272/Y INVX1_LOC_45/A 0.01fF
C9636 NOR2X1_LOC_607/Y INVX1_LOC_53/A 0.03fF
C9637 INVX1_LOC_232/A INVX1_LOC_47/Y 0.10fF
C9638 NAND2X1_LOC_740/Y INVX1_LOC_72/A 0.45fF
C9639 NOR2X1_LOC_92/Y INVX1_LOC_31/A 0.09fF
C9640 NOR2X1_LOC_91/A NAND2X1_LOC_477/A 0.01fF
C9641 NAND2X1_LOC_142/a_36_24# INVX1_LOC_275/Y 0.00fF
C9642 NOR2X1_LOC_186/Y INVX1_LOC_18/A 0.04fF
C9643 INVX1_LOC_41/A INVX1_LOC_23/A 0.17fF
C9644 INVX1_LOC_28/A INVX1_LOC_19/A 0.49fF
C9645 NOR2X1_LOC_388/Y INVX1_LOC_29/Y 0.09fF
C9646 INVX1_LOC_24/Y INVX1_LOC_31/A 0.01fF
C9647 INVX1_LOC_122/Y NOR2X1_LOC_343/B 0.03fF
C9648 INVX1_LOC_25/A INVX1_LOC_34/A 0.66fF
C9649 INVX1_LOC_58/A NAND2X1_LOC_569/A 0.00fF
C9650 INVX1_LOC_103/A NOR2X1_LOC_276/Y -0.03fF
C9651 INVX1_LOC_104/A INVX1_LOC_270/A 0.10fF
C9652 INVX1_LOC_64/A INVX1_LOC_303/A 0.07fF
C9653 INVX1_LOC_249/A INVX1_LOC_5/A 0.09fF
C9654 INVX1_LOC_64/A NOR2X1_LOC_672/Y 0.01fF
C9655 INVX1_LOC_177/A NOR2X1_LOC_383/B 5.98fF
C9656 NOR2X1_LOC_273/a_36_216# INVX1_LOC_27/A 0.01fF
C9657 NAND2X1_LOC_573/Y INVX1_LOC_18/A 0.03fF
C9658 NOR2X1_LOC_382/Y INVX1_LOC_269/A 0.04fF
C9659 NOR2X1_LOC_689/A INVX1_LOC_280/Y 0.00fF
C9660 NAND2X1_LOC_477/A INVX1_LOC_23/A 0.03fF
C9661 INVX1_LOC_2/Y INVX1_LOC_280/A 0.52fF
C9662 INVX1_LOC_50/A NOR2X1_LOC_172/a_36_216# 0.00fF
C9663 INVX1_LOC_1/A NOR2X1_LOC_722/Y 0.02fF
C9664 INVX1_LOC_48/Y INVX1_LOC_72/Y 0.00fF
C9665 NOR2X1_LOC_419/Y INVX1_LOC_50/Y 0.05fF
C9666 NOR2X1_LOC_771/a_36_216# NOR2X1_LOC_89/A 0.01fF
C9667 NOR2X1_LOC_272/Y INVX1_LOC_71/A 0.10fF
C9668 INVX1_LOC_37/A INVX1_LOC_38/A 0.28fF
C9669 NOR2X1_LOC_6/B INVX1_LOC_58/Y -0.04fF
C9670 NAND2X1_LOC_863/B NOR2X1_LOC_829/A 0.18fF
C9671 NOR2X1_LOC_816/a_36_216# NOR2X1_LOC_152/Y 0.01fF
C9672 NAND2X1_LOC_555/Y INPUT_3 0.13fF
C9673 INVX1_LOC_269/A NAND2X1_LOC_530/a_36_24# 0.00fF
C9674 NAND2X1_LOC_564/B NOR2X1_LOC_301/A 0.07fF
C9675 INVX1_LOC_58/A NAND2X1_LOC_661/B 0.00fF
C9676 NOR2X1_LOC_598/B NAND2X1_LOC_629/Y 0.01fF
C9677 INVX1_LOC_136/A INVX1_LOC_103/A 0.10fF
C9678 INVX1_LOC_35/A NAND2X1_LOC_357/B 0.07fF
C9679 INVX1_LOC_279/A NAND2X1_LOC_454/Y 0.02fF
C9680 NAND2X1_LOC_181/Y INVX1_LOC_57/A 0.03fF
C9681 NAND2X1_LOC_785/A NAND2X1_LOC_793/B 0.05fF
C9682 VDD NOR2X1_LOC_332/Y 0.12fF
C9683 NAND2X1_LOC_550/A INVX1_LOC_30/A 0.09fF
C9684 D_INPUT_1 NOR2X1_LOC_78/B 1.10fF
C9685 NOR2X1_LOC_493/B NOR2X1_LOC_717/A 0.09fF
C9686 NOR2X1_LOC_664/Y INVX1_LOC_5/A 0.07fF
C9687 NOR2X1_LOC_318/B NOR2X1_LOC_814/A 0.01fF
C9688 NOR2X1_LOC_160/B INVX1_LOC_30/A 0.63fF
C9689 NOR2X1_LOC_155/A INVX1_LOC_76/A 0.09fF
C9690 NOR2X1_LOC_598/B INVX1_LOC_179/Y 0.14fF
C9691 NOR2X1_LOC_368/A NAND2X1_LOC_455/B 0.01fF
C9692 INVX1_LOC_58/A INVX1_LOC_316/Y 0.00fF
C9693 INVX1_LOC_136/A INVX1_LOC_292/A 0.10fF
C9694 NOR2X1_LOC_240/Y NAND2X1_LOC_359/Y 0.00fF
C9695 INVX1_LOC_266/A NOR2X1_LOC_537/A 0.01fF
C9696 VDD INVX1_LOC_179/A 0.51fF
C9697 INVX1_LOC_93/Y NOR2X1_LOC_814/A 0.09fF
C9698 INVX1_LOC_172/A NAND2X1_LOC_724/A 0.02fF
C9699 NAND2X1_LOC_705/Y INVX1_LOC_207/A 0.01fF
C9700 NOR2X1_LOC_45/Y INVX1_LOC_18/A 0.02fF
C9701 NOR2X1_LOC_598/B NOR2X1_LOC_793/a_36_216# 0.16fF
C9702 INVX1_LOC_90/A NAND2X1_LOC_72/B 0.03fF
C9703 NOR2X1_LOC_91/A NOR2X1_LOC_299/Y 0.03fF
C9704 INVX1_LOC_45/A NOR2X1_LOC_336/B 0.03fF
C9705 NOR2X1_LOC_785/Y NOR2X1_LOC_383/B 0.03fF
C9706 NOR2X1_LOC_553/Y INVX1_LOC_53/A 0.03fF
C9707 NOR2X1_LOC_389/B NAND2X1_LOC_72/B 0.01fF
C9708 NOR2X1_LOC_723/Y NOR2X1_LOC_717/Y 0.00fF
C9709 NOR2X1_LOC_336/B NOR2X1_LOC_568/A 0.04fF
C9710 INVX1_LOC_157/Y INVX1_LOC_38/A 0.01fF
C9711 INVX1_LOC_1/Y NOR2X1_LOC_292/a_36_216# 0.00fF
C9712 INVX1_LOC_87/Y INVX1_LOC_87/A 0.10fF
C9713 INVX1_LOC_246/Y INVX1_LOC_246/A 0.09fF
C9714 NAND2X1_LOC_729/Y INVX1_LOC_161/A 0.00fF
C9715 NAND2X1_LOC_363/B NOR2X1_LOC_516/B 0.10fF
C9716 INVX1_LOC_34/A INVX1_LOC_1/A 0.47fF
C9717 INVX1_LOC_182/A NOR2X1_LOC_334/Y 0.88fF
C9718 INVX1_LOC_223/Y NOR2X1_LOC_168/B 0.00fF
C9719 NAND2X1_LOC_195/Y INVX1_LOC_30/A 0.04fF
C9720 INVX1_LOC_5/A NAND2X1_LOC_200/B 0.03fF
C9721 INVX1_LOC_164/Y INVX1_LOC_306/Y 0.04fF
C9722 NOR2X1_LOC_78/B NOR2X1_LOC_652/Y 0.07fF
C9723 NOR2X1_LOC_789/A NOR2X1_LOC_392/Y 0.01fF
C9724 NAND2X1_LOC_588/B NAND2X1_LOC_36/A 0.02fF
C9725 INVX1_LOC_45/A NAND2X1_LOC_364/A 0.19fF
C9726 VDD INVX1_LOC_250/Y 0.17fF
C9727 NAND2X1_LOC_807/Y NOR2X1_LOC_281/a_36_216# 0.00fF
C9728 INVX1_LOC_89/A NOR2X1_LOC_727/B 0.03fF
C9729 NAND2X1_LOC_570/Y INVX1_LOC_178/A 0.03fF
C9730 NAND2X1_LOC_802/A INVX1_LOC_246/A 0.06fF
C9731 INVX1_LOC_182/Y NAND2X1_LOC_454/Y 0.00fF
C9732 INVX1_LOC_36/A INVX1_LOC_177/Y 0.98fF
C9733 NAND2X1_LOC_637/Y INVX1_LOC_54/A 0.07fF
C9734 NAND2X1_LOC_364/A NOR2X1_LOC_568/A 0.00fF
C9735 INVX1_LOC_31/A NAND2X1_LOC_837/Y 0.19fF
C9736 INVX1_LOC_14/A INVX1_LOC_82/A 0.04fF
C9737 NOR2X1_LOC_99/B NAND2X1_LOC_607/a_36_24# 0.01fF
C9738 NAND2X1_LOC_721/A INVX1_LOC_285/A 0.08fF
C9739 NAND2X1_LOC_650/B INVX1_LOC_63/A 0.08fF
C9740 NAND2X1_LOC_725/Y NOR2X1_LOC_576/B 0.16fF
C9741 NOR2X1_LOC_598/B INVX1_LOC_7/A 0.02fF
C9742 D_INPUT_1 INVX1_LOC_83/A 0.24fF
C9743 NAND2X1_LOC_350/A INVX1_LOC_209/Y 0.72fF
C9744 NAND2X1_LOC_721/A INVX1_LOC_265/Y 0.14fF
C9745 NOR2X1_LOC_92/Y NOR2X1_LOC_290/Y 0.03fF
C9746 INVX1_LOC_280/A NOR2X1_LOC_608/Y 0.39fF
C9747 NOR2X1_LOC_35/Y INVX1_LOC_19/A 0.05fF
C9748 INVX1_LOC_204/Y INVX1_LOC_22/A 0.09fF
C9749 INVX1_LOC_147/Y INVX1_LOC_272/A 0.07fF
C9750 INVX1_LOC_27/A NOR2X1_LOC_773/Y 0.10fF
C9751 NAND2X1_LOC_178/a_36_24# NOR2X1_LOC_180/Y 0.00fF
C9752 NOR2X1_LOC_323/a_36_216# INVX1_LOC_285/A 0.00fF
C9753 NAND2X1_LOC_725/A NOR2X1_LOC_561/Y 0.05fF
C9754 INVX1_LOC_35/A NOR2X1_LOC_128/B 0.18fF
C9755 NOR2X1_LOC_770/B INVX1_LOC_174/A 0.02fF
C9756 NOR2X1_LOC_15/Y NAND2X1_LOC_360/B 0.09fF
C9757 INVX1_LOC_48/A INVX1_LOC_4/Y 0.10fF
C9758 NOR2X1_LOC_205/Y INVX1_LOC_111/Y 0.01fF
C9759 INVX1_LOC_41/A INVX1_LOC_31/A 0.15fF
C9760 INVX1_LOC_5/A INVX1_LOC_234/A 0.10fF
C9761 NAND2X1_LOC_364/A INVX1_LOC_71/A 0.03fF
C9762 NAND2X1_LOC_326/A NAND2X1_LOC_840/B 0.03fF
C9763 NOR2X1_LOC_825/Y INVX1_LOC_284/A 0.15fF
C9764 INVX1_LOC_76/A NOR2X1_LOC_833/B 0.48fF
C9765 INVX1_LOC_232/Y NOR2X1_LOC_817/a_36_216# 0.00fF
C9766 NAND2X1_LOC_214/B NOR2X1_LOC_332/A 0.01fF
C9767 NOR2X1_LOC_15/Y NOR2X1_LOC_165/Y 0.01fF
C9768 NOR2X1_LOC_89/A NOR2X1_LOC_145/Y 0.17fF
C9769 NAND2X1_LOC_112/Y NOR2X1_LOC_321/Y 0.02fF
C9770 INVX1_LOC_64/A NAND2X1_LOC_308/B 0.02fF
C9771 INVX1_LOC_278/A NAND2X1_LOC_842/B 0.01fF
C9772 NOR2X1_LOC_772/a_36_216# INVX1_LOC_1/A 0.00fF
C9773 NOR2X1_LOC_673/B INVX1_LOC_9/A 0.01fF
C9774 NOR2X1_LOC_717/B INVX1_LOC_50/Y 0.03fF
C9775 NOR2X1_LOC_122/A INVX1_LOC_16/A 0.04fF
C9776 INVX1_LOC_178/A INVX1_LOC_234/A 0.10fF
C9777 NOR2X1_LOC_557/A INVX1_LOC_78/A 0.07fF
C9778 INVX1_LOC_2/A INVX1_LOC_230/Y 0.01fF
C9779 NAND2X1_LOC_438/a_36_24# INVX1_LOC_307/A 0.00fF
C9780 INVX1_LOC_256/A NAND2X1_LOC_229/a_36_24# 0.00fF
C9781 INVX1_LOC_47/Y NAND2X1_LOC_447/Y 0.03fF
C9782 NOR2X1_LOC_92/Y NAND2X1_LOC_859/Y 0.38fF
C9783 INVX1_LOC_34/A NOR2X1_LOC_384/Y 0.10fF
C9784 INVX1_LOC_89/A NOR2X1_LOC_649/Y 0.72fF
C9785 INVX1_LOC_27/A NOR2X1_LOC_332/A 0.07fF
C9786 NAND2X1_LOC_53/Y NAND2X1_LOC_841/A 0.24fF
C9787 NOR2X1_LOC_337/A NOR2X1_LOC_748/A 0.03fF
C9788 NOR2X1_LOC_272/Y NOR2X1_LOC_123/B 0.10fF
C9789 INVX1_LOC_36/A INVX1_LOC_104/A 0.09fF
C9790 INVX1_LOC_285/Y NOR2X1_LOC_383/B 0.03fF
C9791 NOR2X1_LOC_124/A NOR2X1_LOC_394/Y 0.09fF
C9792 INVX1_LOC_25/A INPUT_0 0.13fF
C9793 NAND2X1_LOC_724/A NOR2X1_LOC_690/Y 0.01fF
C9794 NOR2X1_LOC_419/Y NOR2X1_LOC_559/B -0.00fF
C9795 INVX1_LOC_17/A NAND2X1_LOC_564/B 0.07fF
C9796 INVX1_LOC_136/A INVX1_LOC_240/A 0.02fF
C9797 INVX1_LOC_225/A INVX1_LOC_18/A 0.13fF
C9798 NAND2X1_LOC_53/Y INVX1_LOC_268/A 0.02fF
C9799 INVX1_LOC_161/Y INVX1_LOC_16/A 2.25fF
C9800 INVX1_LOC_5/A NOR2X1_LOC_19/B 0.15fF
C9801 NOR2X1_LOC_647/A NOR2X1_LOC_78/A 0.01fF
C9802 INVX1_LOC_218/Y INVX1_LOC_218/A 0.32fF
C9803 NOR2X1_LOC_67/A NOR2X1_LOC_606/Y 0.03fF
C9804 NOR2X1_LOC_632/Y INVX1_LOC_11/A 0.01fF
C9805 INVX1_LOC_9/A INVX1_LOC_29/A 0.28fF
C9806 NOR2X1_LOC_88/Y INVX1_LOC_119/Y 0.01fF
C9807 INVX1_LOC_45/A NAND2X1_LOC_11/Y 0.28fF
C9808 NOR2X1_LOC_264/Y NOR2X1_LOC_341/a_36_216# 0.00fF
C9809 INVX1_LOC_39/Y INVX1_LOC_25/Y 0.06fF
C9810 NAND2X1_LOC_571/B INVX1_LOC_309/A 0.05fF
C9811 NAND2X1_LOC_350/B INVX1_LOC_30/A 0.02fF
C9812 INVX1_LOC_31/A NOR2X1_LOC_211/A 0.22fF
C9813 NOR2X1_LOC_209/Y INVX1_LOC_18/A 0.27fF
C9814 NOR2X1_LOC_590/A INVX1_LOC_1/Y 0.04fF
C9815 INVX1_LOC_17/Y INVX1_LOC_91/A 0.03fF
C9816 INVX1_LOC_77/A INVX1_LOC_8/A 0.07fF
C9817 INVX1_LOC_178/A NOR2X1_LOC_19/B 0.19fF
C9818 INVX1_LOC_208/A INVX1_LOC_30/A 0.10fF
C9819 INVX1_LOC_65/A NOR2X1_LOC_383/B 0.03fF
C9820 NAND2X1_LOC_9/Y INVX1_LOC_123/A 0.07fF
C9821 NOR2X1_LOC_784/Y NOR2X1_LOC_148/B 0.00fF
C9822 NOR2X1_LOC_279/Y NOR2X1_LOC_301/A 0.01fF
C9823 NOR2X1_LOC_272/Y INVX1_LOC_102/Y 0.23fF
C9824 VDD INVX1_LOC_165/A -0.00fF
C9825 INVX1_LOC_84/A INVX1_LOC_119/Y 0.03fF
C9826 NOR2X1_LOC_419/Y NOR2X1_LOC_6/B 1.24fF
C9827 NOR2X1_LOC_860/B NOR2X1_LOC_87/B 0.02fF
C9828 INVX1_LOC_36/A INVX1_LOC_263/A -0.00fF
C9829 NOR2X1_LOC_690/A INVX1_LOC_207/A 0.08fF
C9830 NOR2X1_LOC_92/Y NAND2X1_LOC_807/Y 0.95fF
C9831 NOR2X1_LOC_516/B INVX1_LOC_30/A 0.15fF
C9832 NOR2X1_LOC_599/A INVX1_LOC_16/A 0.05fF
C9833 NOR2X1_LOC_328/Y NAND2X1_LOC_741/B 0.36fF
C9834 NOR2X1_LOC_48/B NAND2X1_LOC_637/Y 0.00fF
C9835 NOR2X1_LOC_607/a_36_216# INVX1_LOC_177/A 0.00fF
C9836 INVX1_LOC_26/Y NOR2X1_LOC_35/Y 0.29fF
C9837 NOR2X1_LOC_383/B NOR2X1_LOC_137/B 0.08fF
C9838 NOR2X1_LOC_716/B NOR2X1_LOC_6/B 0.03fF
C9839 D_INPUT_3 INVX1_LOC_26/A 0.18fF
C9840 NOR2X1_LOC_804/B INVX1_LOC_104/A 0.41fF
C9841 NOR2X1_LOC_82/A NAND2X1_LOC_28/a_36_24# 0.02fF
C9842 NOR2X1_LOC_403/B NOR2X1_LOC_78/B 0.30fF
C9843 INVX1_LOC_93/Y NOR2X1_LOC_292/a_36_216# 0.01fF
C9844 VDD NOR2X1_LOC_693/Y 1.07fF
C9845 NOR2X1_LOC_88/Y INVX1_LOC_284/A 0.19fF
C9846 VDD NAND2X1_LOC_288/B 0.01fF
C9847 NOR2X1_LOC_689/Y INVX1_LOC_76/A 0.03fF
C9848 NAND2X1_LOC_552/A NOR2X1_LOC_528/Y 0.01fF
C9849 INVX1_LOC_122/Y NAND2X1_LOC_41/Y 0.02fF
C9850 INVX1_LOC_72/A NOR2X1_LOC_32/Y 0.01fF
C9851 INVX1_LOC_38/A NAND2X1_LOC_72/B 0.03fF
C9852 NOR2X1_LOC_309/Y INVX1_LOC_104/A 0.03fF
C9853 INVX1_LOC_280/Y NAND2X1_LOC_632/B 0.20fF
C9854 INVX1_LOC_230/Y INPUT_1 1.61fF
C9855 INVX1_LOC_161/Y INVX1_LOC_28/A 0.10fF
C9856 NOR2X1_LOC_808/A INVX1_LOC_33/A 0.03fF
C9857 NAND2X1_LOC_471/Y INVX1_LOC_118/A 0.01fF
C9858 INVX1_LOC_1/A INPUT_0 0.21fF
C9859 NOR2X1_LOC_68/A INVX1_LOC_279/A 0.10fF
C9860 NOR2X1_LOC_514/a_36_216# INVX1_LOC_216/A 0.00fF
C9861 INVX1_LOC_50/A NOR2X1_LOC_139/a_36_216# 0.00fF
C9862 NOR2X1_LOC_437/Y INVX1_LOC_16/A 0.98fF
C9863 INVX1_LOC_215/A INVX1_LOC_24/A 0.00fF
C9864 INVX1_LOC_84/A INVX1_LOC_284/A 1.35fF
C9865 NOR2X1_LOC_598/B INVX1_LOC_76/A 0.13fF
C9866 INVX1_LOC_243/Y INVX1_LOC_117/A 0.02fF
C9867 NOR2X1_LOC_92/Y INVX1_LOC_6/A 0.12fF
C9868 D_INPUT_1 INVX1_LOC_46/A 0.18fF
C9869 NAND2X1_LOC_243/B INVX1_LOC_15/A 0.02fF
C9870 NOR2X1_LOC_795/Y NOR2X1_LOC_802/A 0.10fF
C9871 NAND2X1_LOC_493/Y INVX1_LOC_309/A 0.01fF
C9872 NOR2X1_LOC_778/A INVX1_LOC_83/A 0.16fF
C9873 NAND2X1_LOC_859/Y NAND2X1_LOC_837/Y 0.13fF
C9874 INVX1_LOC_298/Y INVX1_LOC_9/A 0.03fF
C9875 NOR2X1_LOC_67/Y INVX1_LOC_63/A 0.01fF
C9876 INVX1_LOC_57/A INVX1_LOC_117/A 1.17fF
C9877 NAND2X1_LOC_708/Y INVX1_LOC_20/A 0.28fF
C9878 INVX1_LOC_30/Y NOR2X1_LOC_419/Y 0.02fF
C9879 NOR2X1_LOC_172/Y INVX1_LOC_53/Y 0.06fF
C9880 NOR2X1_LOC_558/a_36_216# INVX1_LOC_29/Y 0.02fF
C9881 NAND2X1_LOC_725/A INVX1_LOC_76/A 0.10fF
C9882 NOR2X1_LOC_181/A INVX1_LOC_50/Y 0.00fF
C9883 INVX1_LOC_49/A GATE_479 0.03fF
C9884 VDD NOR2X1_LOC_405/Y 0.23fF
C9885 NOR2X1_LOC_590/A NOR2X1_LOC_742/A 0.09fF
C9886 NOR2X1_LOC_373/Y INVX1_LOC_24/A 0.00fF
C9887 INVX1_LOC_30/Y NOR2X1_LOC_716/B 0.03fF
C9888 NAND2X1_LOC_715/B INVX1_LOC_76/A 0.89fF
C9889 NOR2X1_LOC_632/Y NOR2X1_LOC_593/Y 0.02fF
C9890 INVX1_LOC_95/Y NAND2X1_LOC_474/Y 0.07fF
C9891 NOR2X1_LOC_361/Y NOR2X1_LOC_366/B 0.27fF
C9892 INVX1_LOC_90/A NAND2X1_LOC_198/B 0.01fF
C9893 INVX1_LOC_43/A NOR2X1_LOC_709/A 0.05fF
C9894 VDD INVX1_LOC_253/Y 0.21fF
C9895 INVX1_LOC_311/Y INVX1_LOC_142/Y 0.28fF
C9896 NOR2X1_LOC_388/Y INVX1_LOC_101/A 0.02fF
C9897 INVX1_LOC_255/Y NOR2X1_LOC_4/a_36_216# 0.00fF
C9898 NOR2X1_LOC_13/Y INVX1_LOC_89/A 0.13fF
C9899 NOR2X1_LOC_662/A INVX1_LOC_3/Y 0.07fF
C9900 NOR2X1_LOC_401/B INVX1_LOC_256/Y 0.12fF
C9901 INVX1_LOC_46/A NOR2X1_LOC_652/Y 0.07fF
C9902 NAND2X1_LOC_320/a_36_24# NOR2X1_LOC_325/A 0.00fF
C9903 NAND2X1_LOC_364/Y NAND2X1_LOC_363/Y 0.01fF
C9904 INVX1_LOC_311/Y INVX1_LOC_198/Y 0.05fF
C9905 NOR2X1_LOC_861/Y INVX1_LOC_29/A 0.07fF
C9906 INVX1_LOC_1/A NOR2X1_LOC_324/A 0.06fF
C9907 NOR2X1_LOC_451/A INVX1_LOC_296/A 0.21fF
C9908 NAND2X1_LOC_341/A INVX1_LOC_2/A 0.12fF
C9909 NAND2X1_LOC_364/Y INVX1_LOC_89/A 0.01fF
C9910 NOR2X1_LOC_640/Y NOR2X1_LOC_748/A 0.27fF
C9911 INVX1_LOC_290/A INVX1_LOC_266/Y 0.90fF
C9912 NOR2X1_LOC_355/A NOR2X1_LOC_388/Y 0.00fF
C9913 NAND2X1_LOC_562/B INVX1_LOC_234/A 1.17fF
C9914 INVX1_LOC_49/A INVX1_LOC_196/Y 0.05fF
C9915 INVX1_LOC_87/A NOR2X1_LOC_814/A 0.04fF
C9916 NOR2X1_LOC_384/Y INPUT_0 0.01fF
C9917 NOR2X1_LOC_78/B NOR2X1_LOC_553/Y 0.03fF
C9918 NOR2X1_LOC_246/A INVX1_LOC_162/A 0.04fF
C9919 NOR2X1_LOC_590/A NOR2X1_LOC_318/B 0.07fF
C9920 NOR2X1_LOC_457/B NOR2X1_LOC_74/A 0.07fF
C9921 INVX1_LOC_75/A NOR2X1_LOC_546/B 0.55fF
C9922 INVX1_LOC_284/A INVX1_LOC_15/A 0.03fF
C9923 INVX1_LOC_36/A INVX1_LOC_206/Y 0.03fF
C9924 NOR2X1_LOC_68/A NAND2X1_LOC_858/B 0.07fF
C9925 NOR2X1_LOC_498/Y NAND2X1_LOC_866/B 0.01fF
C9926 NAND2X1_LOC_729/Y INPUT_0 0.03fF
C9927 NOR2X1_LOC_135/Y NOR2X1_LOC_433/A 0.04fF
C9928 INVX1_LOC_11/A NAND2X1_LOC_1/Y 0.13fF
C9929 NAND2X1_LOC_341/A NOR2X1_LOC_218/Y 0.07fF
C9930 NOR2X1_LOC_678/A INVX1_LOC_92/A 0.03fF
C9931 NOR2X1_LOC_698/a_36_216# NOR2X1_LOC_698/Y 0.00fF
C9932 INVX1_LOC_181/Y INVX1_LOC_126/Y 0.45fF
C9933 NOR2X1_LOC_82/Y INVX1_LOC_1/Y 0.13fF
C9934 INVX1_LOC_132/A INVX1_LOC_31/Y 0.01fF
C9935 NOR2X1_LOC_272/Y NOR2X1_LOC_331/B 0.44fF
C9936 NOR2X1_LOC_483/B NOR2X1_LOC_631/B 0.24fF
C9937 NAND2X1_LOC_551/A NOR2X1_LOC_315/Y 0.01fF
C9938 INVX1_LOC_75/A INVX1_LOC_275/A 0.07fF
C9939 NAND2X1_LOC_239/a_36_24# INVX1_LOC_90/A 0.00fF
C9940 INVX1_LOC_242/Y VDD 0.26fF
C9941 INVX1_LOC_45/A NOR2X1_LOC_405/A 1.16fF
C9942 NOR2X1_LOC_276/Y NAND2X1_LOC_440/a_36_24# 0.00fF
C9943 INVX1_LOC_36/A NOR2X1_LOC_600/Y 0.06fF
C9944 NOR2X1_LOC_219/B INVX1_LOC_75/A 0.11fF
C9945 NOR2X1_LOC_568/A NOR2X1_LOC_405/A 0.03fF
C9946 NAND2X1_LOC_206/Y NAND2X1_LOC_215/A 0.02fF
C9947 NAND2X1_LOC_562/B NOR2X1_LOC_19/B 0.09fF
C9948 INVX1_LOC_299/A NOR2X1_LOC_319/B 0.00fF
C9949 NOR2X1_LOC_443/Y NOR2X1_LOC_691/B 0.21fF
C9950 NOR2X1_LOC_560/a_36_216# INVX1_LOC_230/A 0.02fF
C9951 NAND2X1_LOC_477/A NAND2X1_LOC_807/Y 0.19fF
C9952 NOR2X1_LOC_334/Y NOR2X1_LOC_850/B 0.02fF
C9953 INVX1_LOC_133/A NAND2X1_LOC_288/B 0.06fF
C9954 INVX1_LOC_200/Y INVX1_LOC_203/A 0.09fF
C9955 NOR2X1_LOC_208/Y INVX1_LOC_206/Y 0.03fF
C9956 INVX1_LOC_5/A NOR2X1_LOC_216/B 0.03fF
C9957 INVX1_LOC_40/Y INVX1_LOC_59/Y 0.00fF
C9958 INVX1_LOC_58/A NOR2X1_LOC_662/A 0.10fF
C9959 INVX1_LOC_250/A INVX1_LOC_11/Y 0.09fF
C9960 INVX1_LOC_18/A NAND2X1_LOC_642/Y 0.09fF
C9961 INVX1_LOC_278/A INVX1_LOC_119/Y 2.79fF
C9962 NAND2X1_LOC_349/B NAND2X1_LOC_656/Y 0.11fF
C9963 INVX1_LOC_39/A NOR2X1_LOC_235/Y 0.04fF
C9964 INVX1_LOC_208/Y NOR2X1_LOC_106/A 0.01fF
C9965 INVX1_LOC_32/A INVX1_LOC_94/Y 0.07fF
C9966 INVX1_LOC_41/A INVX1_LOC_6/A 0.10fF
C9967 INVX1_LOC_26/A NOR2X1_LOC_38/a_36_216# 0.00fF
C9968 INVX1_LOC_45/A NOR2X1_LOC_857/A 0.07fF
C9969 INVX1_LOC_30/A NAND2X1_LOC_211/Y 0.03fF
C9970 INVX1_LOC_215/A NOR2X1_LOC_130/A 0.07fF
C9971 NOR2X1_LOC_641/B VDD 0.12fF
C9972 NOR2X1_LOC_557/Y INVX1_LOC_286/A 0.24fF
C9973 NOR2X1_LOC_495/Y INVX1_LOC_91/A 0.02fF
C9974 INVX1_LOC_295/A NOR2X1_LOC_160/Y 0.03fF
C9975 NOR2X1_LOC_168/B INVX1_LOC_75/A 0.00fF
C9976 INVX1_LOC_90/A INVX1_LOC_53/Y 0.01fF
C9977 NOR2X1_LOC_619/A INVX1_LOC_90/A 0.01fF
C9978 NOR2X1_LOC_405/A INVX1_LOC_71/A 0.20fF
C9979 NOR2X1_LOC_389/B INVX1_LOC_53/Y 0.00fF
C9980 NOR2X1_LOC_55/a_36_216# INVX1_LOC_3/Y 0.01fF
C9981 NAND2X1_LOC_361/Y INVX1_LOC_91/A 0.03fF
C9982 NOR2X1_LOC_807/B NOR2X1_LOC_729/A 0.06fF
C9983 NOR2X1_LOC_751/Y VDD 0.60fF
C9984 NOR2X1_LOC_471/Y NOR2X1_LOC_261/A 0.01fF
C9985 NAND2X1_LOC_477/A INVX1_LOC_6/A 0.05fF
C9986 NOR2X1_LOC_114/Y INVX1_LOC_270/Y 0.10fF
C9987 NOR2X1_LOC_607/a_36_216# NOR2X1_LOC_137/B 0.00fF
C9988 NAND2X1_LOC_3/B NAND2X1_LOC_70/a_36_24# 0.00fF
C9989 NAND2X1_LOC_162/A NOR2X1_LOC_163/Y 0.00fF
C9990 INVX1_LOC_64/A INVX1_LOC_272/A 0.11fF
C9991 NAND2X1_LOC_363/B NAND2X1_LOC_207/B 0.05fF
C9992 INVX1_LOC_94/Y NAND2X1_LOC_175/Y 0.07fF
C9993 NOR2X1_LOC_716/B NOR2X1_LOC_124/A 0.02fF
C9994 INVX1_LOC_122/Y INVX1_LOC_122/A 0.10fF
C9995 INVX1_LOC_34/A NOR2X1_LOC_43/Y 0.02fF
C9996 NOR2X1_LOC_299/Y NAND2X1_LOC_866/B 0.07fF
C9997 INVX1_LOC_45/Y VDD 0.04fF
C9998 INVX1_LOC_18/Y NAND2X1_LOC_72/B 0.14fF
C9999 NOR2X1_LOC_564/Y INVX1_LOC_220/Y 0.04fF
C10000 NOR2X1_LOC_15/Y NAND2X1_LOC_572/B 0.07fF
C10001 INVX1_LOC_57/A INVX1_LOC_3/Y 0.07fF
C10002 NAND2X1_LOC_803/B INVX1_LOC_117/Y 0.02fF
C10003 NAND2X1_LOC_350/A NAND2X1_LOC_434/Y 0.02fF
C10004 INVX1_LOC_286/A INVX1_LOC_143/A 0.01fF
C10005 INVX1_LOC_43/Y NOR2X1_LOC_99/Y 0.61fF
C10006 INVX1_LOC_23/A NOR2X1_LOC_687/a_36_216# 0.00fF
C10007 NOR2X1_LOC_332/A NOR2X1_LOC_19/B 0.17fF
C10008 INVX1_LOC_275/A NAND2X1_LOC_485/a_36_24# 0.00fF
C10009 INVX1_LOC_188/A INVX1_LOC_307/A -0.03fF
C10010 INVX1_LOC_181/Y NOR2X1_LOC_536/A 0.03fF
C10011 NAND2X1_LOC_198/B INVX1_LOC_38/A 0.03fF
C10012 NOR2X1_LOC_654/A INVX1_LOC_273/A 0.03fF
C10013 INVX1_LOC_48/Y INVX1_LOC_19/A 0.03fF
C10014 NAND2X1_LOC_214/B INVX1_LOC_42/A 0.45fF
C10015 NAND2X1_LOC_231/Y NOR2X1_LOC_43/Y 0.36fF
C10016 INVX1_LOC_75/A NAND2X1_LOC_656/Y 0.11fF
C10017 NOR2X1_LOC_773/Y NOR2X1_LOC_528/Y 0.08fF
C10018 INVX1_LOC_81/A INVX1_LOC_281/A 0.02fF
C10019 INVX1_LOC_290/A INVX1_LOC_191/A 0.07fF
C10020 INVX1_LOC_33/A INVX1_LOC_37/A 7.32fF
C10021 INVX1_LOC_271/A INVX1_LOC_78/A 0.03fF
C10022 NAND2X1_LOC_19/a_36_24# NOR2X1_LOC_673/A 0.00fF
C10023 NAND2X1_LOC_326/A INVX1_LOC_49/Y 0.16fF
C10024 NAND2X1_LOC_308/Y INVX1_LOC_76/A 0.27fF
C10025 NAND2X1_LOC_303/Y NOR2X1_LOC_36/B 0.04fF
C10026 NOR2X1_LOC_391/A NOR2X1_LOC_391/Y 0.00fF
C10027 INVX1_LOC_49/A INVX1_LOC_44/A 0.25fF
C10028 INVX1_LOC_27/A INVX1_LOC_42/A 0.12fF
C10029 NOR2X1_LOC_663/A INVX1_LOC_15/A 0.01fF
C10030 INVX1_LOC_24/Y NOR2X1_LOC_633/A 0.01fF
C10031 NOR2X1_LOC_824/A INVX1_LOC_42/A 0.30fF
C10032 NOR2X1_LOC_256/Y INPUT_1 0.01fF
C10033 INVX1_LOC_24/A INVX1_LOC_54/A 0.27fF
C10034 NOR2X1_LOC_142/Y NAND2X1_LOC_472/Y 0.19fF
C10035 INVX1_LOC_7/A INVX1_LOC_201/A 0.03fF
C10036 INVX1_LOC_77/A INVX1_LOC_118/Y 0.04fF
C10037 INVX1_LOC_262/A INVX1_LOC_296/A 0.08fF
C10038 INVX1_LOC_61/A NOR2X1_LOC_235/Y 0.03fF
C10039 INVX1_LOC_89/A NOR2X1_LOC_337/A 0.03fF
C10040 NOR2X1_LOC_180/B NOR2X1_LOC_74/A 0.89fF
C10041 INVX1_LOC_149/A INVX1_LOC_14/Y 0.01fF
C10042 INVX1_LOC_226/Y INVX1_LOC_95/Y 0.04fF
C10043 INVX1_LOC_3/Y INVX1_LOC_252/A 0.04fF
C10044 INVX1_LOC_286/A NOR2X1_LOC_130/A 0.07fF
C10045 NOR2X1_LOC_741/a_36_216# NOR2X1_LOC_742/A 0.01fF
C10046 INVX1_LOC_278/A NOR2X1_LOC_134/a_36_216# 0.01fF
C10047 NOR2X1_LOC_717/B INVX1_LOC_96/A 0.00fF
C10048 INVX1_LOC_58/A INVX1_LOC_57/A 0.55fF
C10049 NOR2X1_LOC_357/Y INVX1_LOC_52/A 0.03fF
C10050 INVX1_LOC_33/A INVX1_LOC_157/Y 0.02fF
C10051 INVX1_LOC_255/Y NAND2X1_LOC_659/B 0.02fF
C10052 INVX1_LOC_8/A INVX1_LOC_9/A 0.12fF
C10053 INVX1_LOC_72/A INVX1_LOC_84/A 0.07fF
C10054 INVX1_LOC_3/Y NOR2X1_LOC_475/A 0.02fF
C10055 INVX1_LOC_299/A INVX1_LOC_32/A 0.07fF
C10056 INVX1_LOC_73/A NOR2X1_LOC_74/A 0.07fF
C10057 INVX1_LOC_136/A NOR2X1_LOC_631/A 0.07fF
C10058 NOR2X1_LOC_91/A NAND2X1_LOC_35/Y 0.22fF
C10059 INVX1_LOC_33/A NOR2X1_LOC_743/Y 0.02fF
C10060 NOR2X1_LOC_644/A NOR2X1_LOC_337/Y 0.02fF
C10061 INVX1_LOC_27/A INVX1_LOC_78/A 3.04fF
C10062 NAND2X1_LOC_11/Y NAND2X1_LOC_635/a_36_24# 0.00fF
C10063 INVX1_LOC_299/A NOR2X1_LOC_623/B 0.05fF
C10064 NAND2X1_LOC_9/Y D_INPUT_1 0.93fF
C10065 NOR2X1_LOC_488/Y NAND2X1_LOC_721/A 0.01fF
C10066 INVX1_LOC_95/A NOR2X1_LOC_130/A 0.03fF
C10067 NOR2X1_LOC_454/Y NOR2X1_LOC_158/a_36_216# 0.00fF
C10068 NOR2X1_LOC_717/B INVX1_LOC_188/Y 0.01fF
C10069 INVX1_LOC_64/A NOR2X1_LOC_125/a_36_216# 0.00fF
C10070 INVX1_LOC_34/Y NOR2X1_LOC_271/Y 0.00fF
C10071 INVX1_LOC_255/Y VDD 3.83fF
C10072 INVX1_LOC_73/A NOR2X1_LOC_9/Y 0.14fF
C10073 INVX1_LOC_233/A D_INPUT_1 0.07fF
C10074 INVX1_LOC_21/A NOR2X1_LOC_301/A 0.01fF
C10075 INVX1_LOC_153/Y INVX1_LOC_179/A 0.01fF
C10076 NOR2X1_LOC_569/A NOR2X1_LOC_74/A 0.05fF
C10077 INVX1_LOC_45/A NOR2X1_LOC_841/a_36_216# 0.00fF
C10078 NOR2X1_LOC_169/B INVX1_LOC_29/A 0.04fF
C10079 INPUT_0 NOR2X1_LOC_188/A 0.03fF
C10080 INVX1_LOC_53/A NOR2X1_LOC_678/A 0.00fF
C10081 INVX1_LOC_18/A NOR2X1_LOC_48/Y 0.01fF
C10082 NAND2X1_LOC_654/B INVX1_LOC_91/A 0.61fF
C10083 NOR2X1_LOC_772/B INVX1_LOC_129/A -0.03fF
C10084 NOR2X1_LOC_78/A INVX1_LOC_148/A 0.00fF
C10085 NAND2X1_LOC_35/Y INVX1_LOC_23/A 0.09fF
C10086 INPUT_0 NOR2X1_LOC_548/B 0.08fF
C10087 INVX1_LOC_75/A INVX1_LOC_78/Y 0.03fF
C10088 INVX1_LOC_140/A NOR2X1_LOC_528/Y 0.10fF
C10089 INVX1_LOC_293/A INVX1_LOC_32/A 0.02fF
C10090 D_INPUT_7 NOR2X1_LOC_1/Y 0.29fF
C10091 INVX1_LOC_121/Y INVX1_LOC_179/A 0.08fF
C10092 INVX1_LOC_77/A NOR2X1_LOC_450/a_36_216# 0.00fF
C10093 NOR2X1_LOC_65/B INVX1_LOC_27/A 0.06fF
C10094 NAND2X1_LOC_190/Y NAND2X1_LOC_454/Y 0.04fF
C10095 NAND2X1_LOC_662/B INVX1_LOC_6/A 0.15fF
C10096 NOR2X1_LOC_225/a_36_216# INVX1_LOC_47/Y 0.01fF
C10097 NOR2X1_LOC_151/Y INVX1_LOC_96/A 0.07fF
C10098 INVX1_LOC_13/A NAND2X1_LOC_96/A 0.11fF
C10099 INVX1_LOC_298/Y NAND2X1_LOC_67/Y 0.03fF
C10100 NOR2X1_LOC_802/A NOR2X1_LOC_862/B 0.10fF
C10101 INVX1_LOC_53/Y INVX1_LOC_38/A 0.06fF
C10102 NOR2X1_LOC_619/A INVX1_LOC_38/A 0.03fF
C10103 NOR2X1_LOC_71/Y VDD 0.51fF
C10104 INVX1_LOC_35/A INVX1_LOC_213/A 0.10fF
C10105 INVX1_LOC_292/A NAND2X1_LOC_647/B 0.01fF
C10106 INVX1_LOC_135/A NOR2X1_LOC_111/A 0.10fF
C10107 NOR2X1_LOC_350/A INVX1_LOC_19/A 0.12fF
C10108 NOR2X1_LOC_598/B NOR2X1_LOC_34/B 0.02fF
C10109 NOR2X1_LOC_469/a_36_216# NOR2X1_LOC_301/A 0.02fF
C10110 INVX1_LOC_119/A NOR2X1_LOC_697/Y 0.01fF
C10111 NAND2X1_LOC_563/Y NOR2X1_LOC_649/B 1.07fF
C10112 NOR2X1_LOC_361/B NAND2X1_LOC_288/B 0.87fF
C10113 NAND2X1_LOC_560/A NOR2X1_LOC_824/Y 0.01fF
C10114 D_INPUT_2 NOR2X1_LOC_671/Y 0.02fF
C10115 NAND2X1_LOC_20/B NOR2X1_LOC_33/Y 0.04fF
C10116 NOR2X1_LOC_460/B INVX1_LOC_19/A 0.02fF
C10117 NOR2X1_LOC_644/A VDD 0.63fF
C10118 NOR2X1_LOC_185/a_36_216# NAND2X1_LOC_642/Y 0.00fF
C10119 NOR2X1_LOC_389/A NAND2X1_LOC_454/Y 0.10fF
C10120 INVX1_LOC_99/Y INVX1_LOC_5/A 0.11fF
C10121 NAND2X1_LOC_724/Y NAND2X1_LOC_724/A 0.00fF
C10122 INVX1_LOC_71/A INVX1_LOC_109/Y 0.07fF
C10123 INVX1_LOC_72/A INVX1_LOC_15/A 0.81fF
C10124 INVX1_LOC_66/A INVX1_LOC_66/Y 0.12fF
C10125 NOR2X1_LOC_773/Y NOR2X1_LOC_216/B 0.10fF
C10126 INVX1_LOC_27/A INVX1_LOC_152/Y 0.14fF
C10127 NOR2X1_LOC_205/Y NOR2X1_LOC_383/B 0.06fF
C10128 INVX1_LOC_13/Y NOR2X1_LOC_211/Y 0.01fF
C10129 INVX1_LOC_104/A INVX1_LOC_63/A 0.07fF
C10130 NAND2X1_LOC_560/A INVX1_LOC_76/A 0.03fF
C10131 NOR2X1_LOC_810/A NOR2X1_LOC_729/A 0.03fF
C10132 INVX1_LOC_24/A NOR2X1_LOC_48/B 3.35fF
C10133 NOR2X1_LOC_315/Y NAND2X1_LOC_489/Y 0.01fF
C10134 NOR2X1_LOC_736/Y INVX1_LOC_139/Y 0.05fF
C10135 NOR2X1_LOC_828/B VDD 0.27fF
C10136 NOR2X1_LOC_753/Y NOR2X1_LOC_89/A 0.11fF
C10137 INVX1_LOC_32/Y NAND2X1_LOC_93/B 0.03fF
C10138 INVX1_LOC_33/A NOR2X1_LOC_178/a_36_216# 0.00fF
C10139 INVX1_LOC_198/Y INVX1_LOC_15/A 0.01fF
C10140 NAND2X1_LOC_722/A NOR2X1_LOC_605/A 0.02fF
C10141 NAND2X1_LOC_338/B INVX1_LOC_84/A 0.07fF
C10142 NAND2X1_LOC_783/A INVX1_LOC_54/A 0.30fF
C10143 NOR2X1_LOC_68/A NOR2X1_LOC_38/B 0.07fF
C10144 NAND2X1_LOC_140/A INVX1_LOC_9/A 0.00fF
C10145 NOR2X1_LOC_772/B NOR2X1_LOC_440/B 0.01fF
C10146 NOR2X1_LOC_798/A NOR2X1_LOC_652/Y 0.04fF
C10147 INVX1_LOC_32/Y NAND2X1_LOC_425/Y 0.03fF
C10148 INVX1_LOC_50/Y NOR2X1_LOC_343/B 0.09fF
C10149 NOR2X1_LOC_130/A INVX1_LOC_54/A 0.07fF
C10150 INVX1_LOC_83/A NOR2X1_LOC_61/Y 0.07fF
C10151 NOR2X1_LOC_92/Y NOR2X1_LOC_109/Y 0.07fF
C10152 NAND2X1_LOC_25/a_36_24# INVX1_LOC_1/A 0.01fF
C10153 NAND2X1_LOC_735/B INVX1_LOC_260/Y 0.02fF
C10154 INVX1_LOC_171/A NOR2X1_LOC_612/Y 0.02fF
C10155 NOR2X1_LOC_664/Y NOR2X1_LOC_847/A 0.01fF
C10156 NOR2X1_LOC_254/a_36_216# NOR2X1_LOC_748/A 0.00fF
C10157 INVX1_LOC_162/Y INVX1_LOC_102/A 0.04fF
C10158 NAND2X1_LOC_451/Y INVX1_LOC_262/Y 0.02fF
C10159 NOR2X1_LOC_204/a_36_216# NOR2X1_LOC_38/B 0.00fF
C10160 INVX1_LOC_89/A NOR2X1_LOC_640/Y 0.03fF
C10161 NOR2X1_LOC_529/Y NOR2X1_LOC_671/Y 0.01fF
C10162 INVX1_LOC_286/A NOR2X1_LOC_280/Y 0.01fF
C10163 INVX1_LOC_30/A NAND2X1_LOC_442/a_36_24# 0.00fF
C10164 NOR2X1_LOC_32/B NOR2X1_LOC_530/Y 0.01fF
C10165 NOR2X1_LOC_220/B INVX1_LOC_1/A 0.01fF
C10166 NOR2X1_LOC_332/A NOR2X1_LOC_216/B 0.07fF
C10167 NOR2X1_LOC_596/A NAND2X1_LOC_454/Y 0.08fF
C10168 INVX1_LOC_133/Y NOR2X1_LOC_89/A 0.03fF
C10169 NOR2X1_LOC_561/Y NAND2X1_LOC_606/a_36_24# 0.06fF
C10170 NOR2X1_LOC_723/Y NOR2X1_LOC_383/B 0.01fF
C10171 INVX1_LOC_179/Y INVX1_LOC_29/A 0.02fF
C10172 INVX1_LOC_206/A INVX1_LOC_42/A 0.07fF
C10173 INVX1_LOC_162/A INVX1_LOC_32/A 0.01fF
C10174 INVX1_LOC_230/Y INVX1_LOC_138/A 0.03fF
C10175 INVX1_LOC_50/A NOR2X1_LOC_703/B 0.03fF
C10176 NOR2X1_LOC_486/Y NOR2X1_LOC_631/B 0.13fF
C10177 NOR2X1_LOC_374/B INVX1_LOC_19/A 0.01fF
C10178 NOR2X1_LOC_531/a_36_216# NOR2X1_LOC_383/B 0.01fF
C10179 NOR2X1_LOC_216/Y INVX1_LOC_54/A 0.60fF
C10180 NOR2X1_LOC_315/Y INVX1_LOC_32/A 0.10fF
C10181 INVX1_LOC_290/A INVX1_LOC_19/A 0.07fF
C10182 INVX1_LOC_75/A NOR2X1_LOC_680/a_36_216# 0.02fF
C10183 NAND2X1_LOC_841/A INVX1_LOC_12/A 0.05fF
C10184 NOR2X1_LOC_551/B NOR2X1_LOC_334/Y 0.02fF
C10185 NOR2X1_LOC_174/A NOR2X1_LOC_862/B 0.11fF
C10186 INVX1_LOC_21/A INVX1_LOC_17/A 0.38fF
C10187 INVX1_LOC_56/Y NAND2X1_LOC_74/B 1.34fF
C10188 INVX1_LOC_33/A NAND2X1_LOC_72/B 2.35fF
C10189 NAND2X1_LOC_35/Y INVX1_LOC_31/A 0.07fF
C10190 NOR2X1_LOC_635/a_36_216# INVX1_LOC_30/A 0.00fF
C10191 INVX1_LOC_35/A NOR2X1_LOC_602/A 0.02fF
C10192 NOR2X1_LOC_433/A NAND2X1_LOC_61/Y 0.15fF
C10193 NOR2X1_LOC_350/A INVX1_LOC_26/Y 0.03fF
C10194 NOR2X1_LOC_45/B INVX1_LOC_37/Y 0.00fF
C10195 INVX1_LOC_268/A INVX1_LOC_12/A 0.02fF
C10196 INVX1_LOC_35/A NOR2X1_LOC_707/B 0.01fF
C10197 NOR2X1_LOC_597/Y NAND2X1_LOC_802/Y 0.02fF
C10198 NAND2X1_LOC_78/a_36_24# INVX1_LOC_30/A 0.00fF
C10199 INVX1_LOC_305/A INVX1_LOC_53/A 0.11fF
C10200 INVX1_LOC_28/A NOR2X1_LOC_841/A 0.03fF
C10201 INVX1_LOC_35/A INVX1_LOC_110/A 0.04fF
C10202 NAND2X1_LOC_338/B INVX1_LOC_15/A 0.08fF
C10203 NOR2X1_LOC_486/Y INVX1_LOC_37/A 0.07fF
C10204 INVX1_LOC_39/A INVX1_LOC_230/Y 0.02fF
C10205 NOR2X1_LOC_540/B VDD -0.00fF
C10206 NAND2X1_LOC_99/Y NOR2X1_LOC_65/B 0.01fF
C10207 NAND2X1_LOC_358/B NAND2X1_LOC_351/A 0.07fF
C10208 INVX1_LOC_313/Y INVX1_LOC_84/A 0.07fF
C10209 NOR2X1_LOC_561/Y INVX1_LOC_29/A 0.10fF
C10210 INVX1_LOC_94/A INVX1_LOC_23/A 0.80fF
C10211 INVX1_LOC_21/A NAND2X1_LOC_555/Y 0.16fF
C10212 NOR2X1_LOC_152/Y INVX1_LOC_271/A 0.03fF
C10213 INVX1_LOC_35/A NOR2X1_LOC_546/A 0.01fF
C10214 NAND2X1_LOC_323/B INVX1_LOC_15/A 6.75fF
C10215 NOR2X1_LOC_309/Y NOR2X1_LOC_281/a_36_216# 0.01fF
C10216 NAND2X1_LOC_679/a_36_24# INVX1_LOC_274/A 0.00fF
C10217 NOR2X1_LOC_828/Y NOR2X1_LOC_500/A 0.01fF
C10218 INVX1_LOC_240/A NOR2X1_LOC_395/Y 0.09fF
C10219 INVX1_LOC_35/A NOR2X1_LOC_196/A 0.00fF
C10220 INVX1_LOC_303/A INVX1_LOC_129/A -0.07fF
C10221 NAND2X1_LOC_107/a_36_24# NOR2X1_LOC_536/A 0.00fF
C10222 NAND2X1_LOC_740/a_36_24# NOR2X1_LOC_15/Y 0.00fF
C10223 NAND2X1_LOC_9/Y NOR2X1_LOC_403/B 0.01fF
C10224 NOR2X1_LOC_500/B NOR2X1_LOC_849/A 0.01fF
C10225 NOR2X1_LOC_844/Y INVX1_LOC_27/A 0.03fF
C10226 NAND2X1_LOC_214/B NOR2X1_LOC_554/B 0.01fF
C10227 INVX1_LOC_285/Y INVX1_LOC_179/A 0.00fF
C10228 NAND2X1_LOC_740/Y NAND2X1_LOC_856/A 0.01fF
C10229 INVX1_LOC_43/Y NOR2X1_LOC_271/B 0.02fF
C10230 INVX1_LOC_234/A INVX1_LOC_42/A 0.36fF
C10231 NOR2X1_LOC_790/B NOR2X1_LOC_550/B 0.00fF
C10232 NAND2X1_LOC_200/B INVX1_LOC_78/A 0.03fF
C10233 NAND2X1_LOC_35/Y NOR2X1_LOC_617/a_36_216# -0.01fF
C10234 INVX1_LOC_11/A NAND2X1_LOC_47/a_36_24# 0.00fF
C10235 INVX1_LOC_27/A NOR2X1_LOC_554/B 0.07fF
C10236 NAND2X1_LOC_800/Y NOR2X1_LOC_48/B 0.00fF
C10237 NOR2X1_LOC_513/Y NOR2X1_LOC_816/A 0.01fF
C10238 INVX1_LOC_17/A NOR2X1_LOC_428/Y 0.05fF
C10239 NOR2X1_LOC_510/Y NOR2X1_LOC_268/a_36_216# -0.02fF
C10240 NOR2X1_LOC_667/A NOR2X1_LOC_301/A 0.06fF
C10241 INVX1_LOC_233/Y NAND2X1_LOC_632/B 0.01fF
C10242 INVX1_LOC_36/A NOR2X1_LOC_92/Y 1.44fF
C10243 INPUT_6 NAND2X1_LOC_59/B 0.13fF
C10244 INVX1_LOC_5/A NOR2X1_LOC_303/Y 0.08fF
C10245 NAND2X1_LOC_465/Y INVX1_LOC_23/A 0.27fF
C10246 INVX1_LOC_225/Y NOR2X1_LOC_794/B -0.00fF
C10247 NOR2X1_LOC_82/A NOR2X1_LOC_590/A 0.03fF
C10248 INVX1_LOC_237/Y NAND2X1_LOC_725/A 0.07fF
C10249 NOR2X1_LOC_92/Y NOR2X1_LOC_267/A 0.04fF
C10250 NAND2X1_LOC_292/a_36_24# INVX1_LOC_26/Y 0.01fF
C10251 NAND2X1_LOC_363/B NOR2X1_LOC_264/Y 0.01fF
C10252 NOR2X1_LOC_396/Y INVX1_LOC_241/Y 0.06fF
C10253 NOR2X1_LOC_244/B NOR2X1_LOC_342/B 0.04fF
C10254 INVX1_LOC_251/Y INVX1_LOC_29/Y 0.09fF
C10255 INVX1_LOC_17/Y NAND2X1_LOC_374/Y 0.04fF
C10256 INVX1_LOC_232/A INVX1_LOC_23/Y 0.10fF
C10257 NOR2X1_LOC_280/Y INVX1_LOC_54/A 0.03fF
C10258 NAND2X1_LOC_177/a_36_24# INVX1_LOC_53/A 0.01fF
C10259 NOR2X1_LOC_65/B NOR2X1_LOC_251/Y 0.24fF
C10260 INVX1_LOC_200/Y NAND2X1_LOC_374/Y 0.22fF
C10261 NOR2X1_LOC_19/B INVX1_LOC_42/A 0.50fF
C10262 NOR2X1_LOC_15/Y NOR2X1_LOC_609/A 0.03fF
C10263 INVX1_LOC_14/A NOR2X1_LOC_360/Y 0.01fF
C10264 INVX1_LOC_38/A INVX1_LOC_77/Y 0.11fF
C10265 INVX1_LOC_5/A NOR2X1_LOC_254/Y 0.54fF
C10266 NAND2X1_LOC_724/Y NAND2X1_LOC_852/Y 0.47fF
C10267 INVX1_LOC_10/A INVX1_LOC_271/Y 0.04fF
C10268 INVX1_LOC_229/Y NOR2X1_LOC_409/B 0.03fF
C10269 NAND2X1_LOC_778/Y NOR2X1_LOC_716/B 0.10fF
C10270 INVX1_LOC_17/A NAND2X1_LOC_354/Y 0.34fF
C10271 INVX1_LOC_115/A NAND2X1_LOC_93/B 0.01fF
C10272 INVX1_LOC_5/A NOR2X1_LOC_84/A 0.08fF
C10273 INVX1_LOC_27/A INVX1_LOC_113/Y 0.14fF
C10274 NAND2X1_LOC_840/B NOR2X1_LOC_654/A 0.01fF
C10275 INVX1_LOC_135/A INVX1_LOC_253/A 0.05fF
C10276 NAND2X1_LOC_690/a_36_24# INVX1_LOC_53/A 0.00fF
C10277 NAND2X1_LOC_22/a_36_24# D_INPUT_6 0.00fF
C10278 INVX1_LOC_135/A INVX1_LOC_90/Y 0.03fF
C10279 NAND2X1_LOC_564/B INVX1_LOC_181/A 0.08fF
C10280 INVX1_LOC_13/A NAND2X1_LOC_99/A 0.12fF
C10281 NAND2X1_LOC_477/A NOR2X1_LOC_109/Y 0.10fF
C10282 VDD NAND2X1_LOC_243/Y 0.48fF
C10283 NOR2X1_LOC_136/Y INVX1_LOC_23/A 0.00fF
C10284 NOR2X1_LOC_302/B NOR2X1_LOC_727/B 0.00fF
C10285 NOR2X1_LOC_167/Y INVX1_LOC_29/A 0.02fF
C10286 VDD INVX1_LOC_89/Y -0.00fF
C10287 NOR2X1_LOC_92/Y NOR2X1_LOC_237/Y 0.07fF
C10288 NAND2X1_LOC_9/Y NOR2X1_LOC_620/B 0.01fF
C10289 INVX1_LOC_115/A NAND2X1_LOC_425/Y 0.01fF
C10290 NOR2X1_LOC_15/Y NOR2X1_LOC_419/Y 0.01fF
C10291 NOR2X1_LOC_78/B NOR2X1_LOC_678/A 0.03fF
C10292 NOR2X1_LOC_58/Y INVX1_LOC_76/A 0.03fF
C10293 NAND2X1_LOC_35/Y NOR2X1_LOC_290/Y 0.04fF
C10294 INVX1_LOC_274/A INVX1_LOC_117/A 0.72fF
C10295 NOR2X1_LOC_51/A INVX1_LOC_77/Y 0.17fF
C10296 NOR2X1_LOC_528/a_36_216# NOR2X1_LOC_693/Y 0.01fF
C10297 INVX1_LOC_256/A INVX1_LOC_181/Y 0.18fF
C10298 INVX1_LOC_88/A NAND2X1_LOC_593/Y 0.24fF
C10299 NOR2X1_LOC_15/Y NOR2X1_LOC_716/B 0.14fF
C10300 INVX1_LOC_45/A NOR2X1_LOC_726/Y 0.05fF
C10301 INVX1_LOC_5/A NOR2X1_LOC_353/Y 0.03fF
C10302 NOR2X1_LOC_68/A NOR2X1_LOC_389/A 0.10fF
C10303 INVX1_LOC_24/Y NOR2X1_LOC_804/B 0.07fF
C10304 INVX1_LOC_103/A NAND2X1_LOC_567/Y 0.73fF
C10305 INVX1_LOC_118/Y INVX1_LOC_9/A 0.03fF
C10306 INVX1_LOC_11/A INVX1_LOC_180/A 0.06fF
C10307 NAND2X1_LOC_566/a_36_24# NAND2X1_LOC_567/Y 0.00fF
C10308 INVX1_LOC_20/A NOR2X1_LOC_673/A 0.03fF
C10309 INVX1_LOC_289/Y NAND2X1_LOC_354/B 0.03fF
C10310 NOR2X1_LOC_859/A NOR2X1_LOC_500/B 0.04fF
C10311 NOR2X1_LOC_92/Y NOR2X1_LOC_309/Y 0.57fF
C10312 NOR2X1_LOC_588/A INVX1_LOC_12/A 0.01fF
C10313 INVX1_LOC_218/Y INVX1_LOC_24/A 0.23fF
C10314 INVX1_LOC_176/A NOR2X1_LOC_814/A 0.03fF
C10315 NAND2X1_LOC_181/Y INVX1_LOC_306/Y 1.93fF
C10316 NAND2X1_LOC_551/A NAND2X1_LOC_99/A 0.33fF
C10317 INVX1_LOC_11/A NOR2X1_LOC_520/B 0.71fF
C10318 NOR2X1_LOC_441/Y INVX1_LOC_24/A 0.05fF
C10319 NOR2X1_LOC_528/Y INVX1_LOC_42/A 0.01fF
C10320 INVX1_LOC_11/A NAND2X1_LOC_325/Y 0.03fF
C10321 NOR2X1_LOC_254/A INVX1_LOC_49/A 0.17fF
C10322 INVX1_LOC_93/A NOR2X1_LOC_773/Y 0.01fF
C10323 INVX1_LOC_81/Y NOR2X1_LOC_759/Y 0.00fF
C10324 NOR2X1_LOC_272/Y NOR2X1_LOC_366/B 0.03fF
C10325 INVX1_LOC_1/A INVX1_LOC_266/Y 0.17fF
C10326 INVX1_LOC_95/Y INVX1_LOC_12/A 0.07fF
C10327 NAND2X1_LOC_35/Y NAND2X1_LOC_859/Y 0.10fF
C10328 NOR2X1_LOC_65/B NOR2X1_LOC_772/A 0.02fF
C10329 NAND2X1_LOC_392/a_36_24# INVX1_LOC_256/Y 0.00fF
C10330 NOR2X1_LOC_91/Y INVX1_LOC_18/A 0.68fF
C10331 INVX1_LOC_36/A NAND2X1_LOC_837/Y 0.07fF
C10332 INVX1_LOC_225/A NAND2X1_LOC_793/Y 0.03fF
C10333 NOR2X1_LOC_15/Y INVX1_LOC_98/Y 0.01fF
C10334 INVX1_LOC_256/A NOR2X1_LOC_192/a_36_216# 0.02fF
C10335 INVX1_LOC_141/Y NOR2X1_LOC_577/Y 0.00fF
C10336 INVX1_LOC_83/A INVX1_LOC_295/Y 0.01fF
C10337 INVX1_LOC_76/A INVX1_LOC_29/A 0.10fF
C10338 INVX1_LOC_8/Y INVX1_LOC_30/A 0.02fF
C10339 NOR2X1_LOC_238/Y INVX1_LOC_217/A 0.44fF
C10340 NOR2X1_LOC_88/Y NOR2X1_LOC_506/Y 0.28fF
C10341 D_INPUT_1 NAND2X1_LOC_842/B 0.10fF
C10342 NOR2X1_LOC_742/A NOR2X1_LOC_632/a_36_216# 0.01fF
C10343 NOR2X1_LOC_68/A NOR2X1_LOC_596/A 0.56fF
C10344 NOR2X1_LOC_78/A INVX1_LOC_47/Y 0.00fF
C10345 INVX1_LOC_135/A INVX1_LOC_138/Y 0.01fF
C10346 INVX1_LOC_232/Y INVX1_LOC_269/A 0.08fF
C10347 NOR2X1_LOC_766/a_36_216# NAND2X1_LOC_811/Y 0.00fF
C10348 NOR2X1_LOC_717/Y NOR2X1_LOC_717/a_36_216# 0.02fF
C10349 INVX1_LOC_135/A NOR2X1_LOC_860/a_36_216# 0.00fF
C10350 INVX1_LOC_75/A NOR2X1_LOC_727/B 0.03fF
C10351 NAND2X1_LOC_84/Y NOR2X1_LOC_360/Y 0.08fF
C10352 INVX1_LOC_171/A NAND2X1_LOC_406/a_36_24# 0.02fF
C10353 NOR2X1_LOC_475/a_36_216# INVX1_LOC_269/A 0.00fF
C10354 INVX1_LOC_17/A NOR2X1_LOC_667/A 0.08fF
C10355 NAND2X1_LOC_773/Y INVX1_LOC_226/Y 0.03fF
C10356 NOR2X1_LOC_67/A INVX1_LOC_11/A 0.07fF
C10357 INVX1_LOC_17/A INVX1_LOC_248/A 0.07fF
C10358 INVX1_LOC_41/A INVX1_LOC_36/A 0.10fF
C10359 INVX1_LOC_172/A NOR2X1_LOC_91/Y 0.03fF
C10360 INVX1_LOC_230/Y NOR2X1_LOC_93/a_36_216# 0.01fF
C10361 INVX1_LOC_311/A NOR2X1_LOC_302/A 0.03fF
C10362 INVX1_LOC_50/A INVX1_LOC_79/A 0.02fF
C10363 NOR2X1_LOC_445/Y NOR2X1_LOC_568/A 0.01fF
C10364 NOR2X1_LOC_498/Y INVX1_LOC_36/A 0.07fF
C10365 NAND2X1_LOC_35/Y NAND2X1_LOC_866/B 0.07fF
C10366 NOR2X1_LOC_528/Y INVX1_LOC_78/A 0.30fF
C10367 NOR2X1_LOC_100/A NOR2X1_LOC_590/A 0.00fF
C10368 INVX1_LOC_300/Y NOR2X1_LOC_387/Y 0.00fF
C10369 INVX1_LOC_41/A NOR2X1_LOC_267/A 0.41fF
C10370 NOR2X1_LOC_478/a_36_216# NAND2X1_LOC_149/Y 0.01fF
C10371 NAND2X1_LOC_114/B NOR2X1_LOC_346/B 0.00fF
C10372 NAND2X1_LOC_198/B INVX1_LOC_33/A 0.03fF
C10373 INVX1_LOC_144/A INVX1_LOC_23/A 0.08fF
C10374 NOR2X1_LOC_481/A NOR2X1_LOC_607/A 0.07fF
C10375 NOR2X1_LOC_434/a_36_216# NOR2X1_LOC_843/A 0.00fF
C10376 INVX1_LOC_36/A NAND2X1_LOC_477/A 0.03fF
C10377 INVX1_LOC_75/A NOR2X1_LOC_717/A 1.03fF
C10378 NOR2X1_LOC_82/A NOR2X1_LOC_82/Y 0.00fF
C10379 INVX1_LOC_5/A NOR2X1_LOC_112/Y 0.03fF
C10380 INVX1_LOC_249/A INVX1_LOC_113/Y 0.00fF
C10381 INVX1_LOC_279/Y NOR2X1_LOC_778/B 0.01fF
C10382 NAND2X1_LOC_729/Y NAND2X1_LOC_811/Y 0.00fF
C10383 NAND2X1_LOC_842/B NOR2X1_LOC_652/Y 0.08fF
C10384 NOR2X1_LOC_68/A NOR2X1_LOC_844/A 0.06fF
C10385 INVX1_LOC_24/A NOR2X1_LOC_142/Y 0.07fF
C10386 NOR2X1_LOC_758/Y NOR2X1_LOC_758/a_36_216# 0.00fF
C10387 NOR2X1_LOC_15/Y NOR2X1_LOC_717/B 0.02fF
C10388 INPUT_4 NOR2X1_LOC_25/Y 0.07fF
C10389 NOR2X1_LOC_445/Y INVX1_LOC_71/A 0.00fF
C10390 NAND2X1_LOC_447/Y NAND2X1_LOC_447/a_36_24# 0.02fF
C10391 INVX1_LOC_235/Y INVX1_LOC_90/A 0.51fF
C10392 NAND2X1_LOC_114/B INVX1_LOC_22/A 0.02fF
C10393 NAND2X1_LOC_454/Y NAND2X1_LOC_469/B 0.22fF
C10394 NOR2X1_LOC_536/A NOR2X1_LOC_114/Y 0.01fF
C10395 NOR2X1_LOC_791/Y NAND2X1_LOC_850/A 0.42fF
C10396 INVX1_LOC_304/A NOR2X1_LOC_301/A 0.02fF
C10397 NAND2X1_LOC_149/Y INVX1_LOC_90/A 0.15fF
C10398 NOR2X1_LOC_15/Y NAND2X1_LOC_656/a_36_24# 0.01fF
C10399 VDD INVX1_LOC_21/Y 0.05fF
C10400 NOR2X1_LOC_409/B INVX1_LOC_20/A 0.03fF
C10401 INVX1_LOC_50/A INVX1_LOC_91/A 0.52fF
C10402 NOR2X1_LOC_454/Y D_GATE_366 0.07fF
C10403 NAND2X1_LOC_555/Y NAND2X1_LOC_6/a_36_24# 0.00fF
C10404 INVX1_LOC_34/A NOR2X1_LOC_625/Y 0.02fF
C10405 NOR2X1_LOC_361/B NOR2X1_LOC_71/Y 0.10fF
C10406 INVX1_LOC_230/Y NAND2X1_LOC_735/B 0.00fF
C10407 NAND2X1_LOC_96/A INVX1_LOC_32/A 0.01fF
C10408 INVX1_LOC_304/Y NOR2X1_LOC_238/Y 0.02fF
C10409 NOR2X1_LOC_139/Y INVX1_LOC_270/Y 0.01fF
C10410 INVX1_LOC_222/A NAND2X1_LOC_406/a_36_24# 0.01fF
C10411 INVX1_LOC_41/A NOR2X1_LOC_804/B 0.08fF
C10412 NAND2X1_LOC_276/Y NAND2X1_LOC_361/Y 0.00fF
C10413 INVX1_LOC_33/A INVX1_LOC_310/Y 0.07fF
C10414 INVX1_LOC_45/Y INVX1_LOC_177/A 0.03fF
C10415 INVX1_LOC_57/Y NAND2X1_LOC_862/A 0.17fF
C10416 INVX1_LOC_39/A NOR2X1_LOC_256/Y 0.01fF
C10417 INVX1_LOC_298/Y INVX1_LOC_76/A 0.15fF
C10418 NAND2X1_LOC_785/B INVX1_LOC_16/A 0.23fF
C10419 NOR2X1_LOC_382/Y NOR2X1_LOC_516/B 0.03fF
C10420 INVX1_LOC_50/A INVX1_LOC_11/Y 0.10fF
C10421 NOR2X1_LOC_557/Y NOR2X1_LOC_142/Y 0.00fF
C10422 NOR2X1_LOC_220/B NOR2X1_LOC_188/A 0.06fF
C10423 NOR2X1_LOC_237/Y NAND2X1_LOC_477/A 0.10fF
C10424 NOR2X1_LOC_655/B INVX1_LOC_24/A 0.01fF
C10425 INVX1_LOC_136/A INVX1_LOC_56/Y 0.03fF
C10426 NAND2X1_LOC_350/A NOR2X1_LOC_130/A 0.10fF
C10427 NOR2X1_LOC_631/B NOR2X1_LOC_748/A 0.03fF
C10428 INVX1_LOC_223/Y NOR2X1_LOC_337/A 0.01fF
C10429 VDD INVX1_LOC_16/Y 0.45fF
C10430 NOR2X1_LOC_15/Y INVX1_LOC_135/Y 0.09fF
C10431 NOR2X1_LOC_252/a_36_216# INVX1_LOC_217/A 0.15fF
C10432 NOR2X1_LOC_590/A INVX1_LOC_306/A 0.02fF
C10433 INVX1_LOC_27/A INVX1_LOC_158/Y 0.03fF
C10434 INVX1_LOC_80/A NOR2X1_LOC_514/A 0.20fF
C10435 NOR2X1_LOC_433/A INVX1_LOC_133/Y 0.09fF
C10436 NOR2X1_LOC_179/a_36_216# NAND2X1_LOC_74/B 0.00fF
C10437 NOR2X1_LOC_216/B NOR2X1_LOC_847/A 0.02fF
C10438 INVX1_LOC_2/A NOR2X1_LOC_219/a_36_216# 0.00fF
C10439 NOR2X1_LOC_829/Y INVX1_LOC_76/A 0.09fF
C10440 INVX1_LOC_77/A NOR2X1_LOC_520/A 0.08fF
C10441 INVX1_LOC_50/A NOR2X1_LOC_421/Y 0.16fF
C10442 INVX1_LOC_276/A NOR2X1_LOC_433/A 0.16fF
C10443 NAND2X1_LOC_72/Y INVX1_LOC_91/A 0.02fF
C10444 NOR2X1_LOC_667/A NAND2X1_LOC_547/a_36_24# 0.00fF
C10445 NAND2X1_LOC_374/Y NOR2X1_LOC_495/Y 0.00fF
C10446 VDD NOR2X1_LOC_39/Y 0.18fF
C10447 NOR2X1_LOC_15/Y NOR2X1_LOC_151/Y 0.14fF
C10448 NOR2X1_LOC_216/B INVX1_LOC_42/A 0.04fF
C10449 NOR2X1_LOC_441/Y NOR2X1_LOC_130/A 0.14fF
C10450 INVX1_LOC_37/A NOR2X1_LOC_635/B 0.02fF
C10451 NOR2X1_LOC_763/Y NAND2X1_LOC_36/A 0.00fF
C10452 NOR2X1_LOC_350/a_36_216# INVX1_LOC_158/A 0.02fF
C10453 NOR2X1_LOC_419/Y INVX1_LOC_226/A 0.00fF
C10454 INVX1_LOC_44/A NOR2X1_LOC_631/Y 0.25fF
C10455 NOR2X1_LOC_309/Y NAND2X1_LOC_477/A 0.10fF
C10456 NOR2X1_LOC_655/B NOR2X1_LOC_557/Y 0.10fF
C10457 INVX1_LOC_37/A NOR2X1_LOC_748/A 0.06fF
C10458 NOR2X1_LOC_340/A NOR2X1_LOC_814/A 0.05fF
C10459 NAND2X1_LOC_691/a_36_24# INVX1_LOC_72/A 0.00fF
C10460 VDD NAND2X1_LOC_205/A 0.67fF
C10461 INVX1_LOC_13/A NAND2X1_LOC_656/A 0.01fF
C10462 NAND2X1_LOC_338/B NAND2X1_LOC_464/Y 0.06fF
C10463 INVX1_LOC_17/A NAND2X1_LOC_51/B 0.03fF
C10464 NOR2X1_LOC_440/Y INVX1_LOC_181/Y 0.00fF
C10465 NOR2X1_LOC_234/Y NOR2X1_LOC_290/Y 0.06fF
C10466 INVX1_LOC_305/A INVX1_LOC_83/A 0.07fF
C10467 INVX1_LOC_84/A NOR2X1_LOC_226/Y 0.07fF
C10468 INVX1_LOC_135/A NAND2X1_LOC_364/A 2.53fF
C10469 INVX1_LOC_50/A NOR2X1_LOC_698/Y 0.11fF
C10470 INVX1_LOC_276/A NOR2X1_LOC_52/B 0.10fF
C10471 INVX1_LOC_46/A NOR2X1_LOC_678/A 0.03fF
C10472 INVX1_LOC_33/A INVX1_LOC_53/Y 0.37fF
C10473 NOR2X1_LOC_67/A NOR2X1_LOC_52/B 0.07fF
C10474 INVX1_LOC_214/Y NOR2X1_LOC_574/A 0.00fF
C10475 NOR2X1_LOC_772/Y INVX1_LOC_16/A 0.09fF
C10476 NOR2X1_LOC_126/a_36_216# INVX1_LOC_42/A 0.00fF
C10477 INVX1_LOC_45/A INVX1_LOC_311/Y 0.04fF
C10478 INVX1_LOC_24/A NOR2X1_LOC_99/B 0.17fF
C10479 NAND2X1_LOC_483/Y INVX1_LOC_22/A 0.12fF
C10480 INVX1_LOC_225/Y NOR2X1_LOC_188/A 0.13fF
C10481 NOR2X1_LOC_216/B INVX1_LOC_78/A 1.27fF
C10482 INVX1_LOC_33/A NOR2X1_LOC_665/A 0.03fF
C10483 NOR2X1_LOC_471/Y INVX1_LOC_311/A 0.02fF
C10484 NOR2X1_LOC_392/B INVX1_LOC_16/A 0.12fF
C10485 INVX1_LOC_225/Y NOR2X1_LOC_548/B 0.02fF
C10486 NOR2X1_LOC_655/B INVX1_LOC_143/A 0.10fF
C10487 NOR2X1_LOC_75/Y NOR2X1_LOC_733/Y 0.00fF
C10488 NAND2X1_LOC_157/a_36_24# GATE_662 0.00fF
C10489 NAND2X1_LOC_739/a_36_24# INVX1_LOC_76/A 0.01fF
C10490 NAND2X1_LOC_326/A NAND2X1_LOC_649/B 0.03fF
C10491 NAND2X1_LOC_656/Y NOR2X1_LOC_577/Y 0.10fF
C10492 NOR2X1_LOC_658/Y INVX1_LOC_75/A 0.10fF
C10493 INVX1_LOC_90/A NOR2X1_LOC_744/Y 0.01fF
C10494 INVX1_LOC_54/Y NOR2X1_LOC_773/Y 0.40fF
C10495 NOR2X1_LOC_19/B NOR2X1_LOC_554/B 0.08fF
C10496 INVX1_LOC_104/A INVX1_LOC_1/Y 0.09fF
C10497 NOR2X1_LOC_226/A INVX1_LOC_144/Y 0.06fF
C10498 INVX1_LOC_145/Y INVX1_LOC_33/A 0.01fF
C10499 NAND2X1_LOC_173/a_36_24# INVX1_LOC_149/A 0.01fF
C10500 NAND2X1_LOC_564/B NOR2X1_LOC_315/Y 0.22fF
C10501 INVX1_LOC_232/Y NAND2X1_LOC_563/A 0.07fF
C10502 INVX1_LOC_7/A INVX1_LOC_8/A 0.09fF
C10503 NOR2X1_LOC_616/Y INVX1_LOC_197/Y -0.04fF
C10504 INVX1_LOC_45/A NOR2X1_LOC_335/B 0.04fF
C10505 INVX1_LOC_19/A NOR2X1_LOC_467/A 0.02fF
C10506 INVX1_LOC_77/A D_GATE_366 0.08fF
C10507 INVX1_LOC_24/A INVX1_LOC_182/A 0.07fF
C10508 NOR2X1_LOC_65/B NOR2X1_LOC_216/B 0.42fF
C10509 INVX1_LOC_58/A NAND2X1_LOC_241/a_36_24# 0.01fF
C10510 NOR2X1_LOC_332/A NOR2X1_LOC_84/A 0.24fF
C10511 INVX1_LOC_256/Y INVX1_LOC_25/Y 0.00fF
C10512 INVX1_LOC_117/A INVX1_LOC_306/Y 0.35fF
C10513 INVX1_LOC_138/Y INVX1_LOC_280/A 0.03fF
C10514 INVX1_LOC_78/A NAND2X1_LOC_477/Y 0.25fF
C10515 INVX1_LOC_17/A INVX1_LOC_304/A 0.03fF
C10516 INVX1_LOC_286/Y INVX1_LOC_286/A 0.29fF
C10517 INVX1_LOC_21/A NOR2X1_LOC_706/B 0.01fF
C10518 NAND2X1_LOC_793/Y NAND2X1_LOC_642/Y 0.02fF
C10519 NOR2X1_LOC_860/a_36_216# INVX1_LOC_280/A 0.01fF
C10520 NOR2X1_LOC_272/Y NOR2X1_LOC_813/Y 0.03fF
C10521 NAND2X1_LOC_796/B INVX1_LOC_33/Y 0.50fF
C10522 INVX1_LOC_300/A NAND2X1_LOC_852/Y 0.01fF
C10523 NOR2X1_LOC_281/a_36_216# INVX1_LOC_63/A 0.01fF
C10524 NOR2X1_LOC_15/Y NAND2X1_LOC_633/Y 0.07fF
C10525 NOR2X1_LOC_155/A INVX1_LOC_23/A 4.96fF
C10526 NOR2X1_LOC_172/Y INVX1_LOC_28/A 0.09fF
C10527 NAND2X1_LOC_331/a_36_24# NOR2X1_LOC_52/B 0.00fF
C10528 NAND2X1_LOC_358/Y INVX1_LOC_143/A 0.00fF
C10529 INVX1_LOC_58/A NAND2X1_LOC_243/a_36_24# 0.00fF
C10530 INVX1_LOC_128/A INVX1_LOC_109/A 0.03fF
C10531 NAND2X1_LOC_99/A NAND2X1_LOC_489/Y 0.00fF
C10532 NOR2X1_LOC_360/Y INVX1_LOC_48/A 0.07fF
C10533 NOR2X1_LOC_335/B INVX1_LOC_71/A 0.03fF
C10534 NOR2X1_LOC_88/Y NAND2X1_LOC_793/B 0.07fF
C10535 INVX1_LOC_224/Y INVX1_LOC_84/A 0.03fF
C10536 NOR2X1_LOC_392/B INVX1_LOC_28/A 0.07fF
C10537 NOR2X1_LOC_817/Y VDD 0.32fF
C10538 NOR2X1_LOC_336/B NOR2X1_LOC_552/A 0.01fF
C10539 NOR2X1_LOC_589/a_36_216# INVX1_LOC_113/Y 0.00fF
C10540 NAND2X1_LOC_149/Y INVX1_LOC_38/A 0.68fF
C10541 INVX1_LOC_57/A NAND2X1_LOC_475/Y 0.00fF
C10542 INVX1_LOC_5/A NOR2X1_LOC_78/Y 0.05fF
C10543 INVX1_LOC_268/Y GATE_662 0.00fF
C10544 NOR2X1_LOC_191/B INVX1_LOC_286/A 0.01fF
C10545 NAND2X1_LOC_725/B NOR2X1_LOC_536/A 0.03fF
C10546 NOR2X1_LOC_644/A INVX1_LOC_177/A 0.06fF
C10547 INVX1_LOC_234/A NAND2X1_LOC_859/B 0.06fF
C10548 NOR2X1_LOC_590/A INVX1_LOC_176/A 0.09fF
C10549 INVX1_LOC_230/Y D_INPUT_3 0.45fF
C10550 NAND2X1_LOC_656/Y INVX1_LOC_22/A 0.07fF
C10551 INVX1_LOC_33/A NOR2X1_LOC_113/B 0.03fF
C10552 NAND2X1_LOC_507/a_36_24# INVX1_LOC_173/Y 0.01fF
C10553 INVX1_LOC_209/Y NOR2X1_LOC_387/A 0.00fF
C10554 INVX1_LOC_49/Y NOR2X1_LOC_654/A 0.03fF
C10555 NOR2X1_LOC_441/Y NOR2X1_LOC_280/Y 0.04fF
C10556 NAND2X1_LOC_807/Y NOR2X1_LOC_312/a_36_216# 0.01fF
C10557 INVX1_LOC_84/A NAND2X1_LOC_793/B 0.08fF
C10558 INVX1_LOC_236/A NOR2X1_LOC_329/B 0.15fF
C10559 NOR2X1_LOC_15/Y NOR2X1_LOC_709/B 0.01fF
C10560 NAND2X1_LOC_787/A NOR2X1_LOC_662/A 0.02fF
C10561 INVX1_LOC_28/A NAND2X1_LOC_294/a_36_24# 0.01fF
C10562 NOR2X1_LOC_152/a_36_216# INVX1_LOC_91/A 0.00fF
C10563 INVX1_LOC_279/A INVX1_LOC_10/A 0.14fF
C10564 INVX1_LOC_135/A NOR2X1_LOC_86/A 0.10fF
C10565 NOR2X1_LOC_413/Y NOR2X1_LOC_20/a_36_216# 0.01fF
C10566 INPUT_3 NAND2X1_LOC_96/A 0.02fF
C10567 INVX1_LOC_2/A NOR2X1_LOC_322/Y 0.07fF
C10568 NOR2X1_LOC_486/a_36_216# INVX1_LOC_117/A 0.01fF
C10569 INVX1_LOC_90/A INVX1_LOC_16/A 0.17fF
C10570 INVX1_LOC_49/A NOR2X1_LOC_562/B 0.12fF
C10571 INVX1_LOC_77/A NOR2X1_LOC_746/Y 0.04fF
C10572 NOR2X1_LOC_228/a_36_216# NOR2X1_LOC_78/A 0.00fF
C10573 NOR2X1_LOC_426/Y NOR2X1_LOC_425/Y 0.00fF
C10574 NOR2X1_LOC_426/a_36_216# INVX1_LOC_77/Y 0.02fF
C10575 INVX1_LOC_45/Y NOR2X1_LOC_137/B 0.03fF
C10576 INVX1_LOC_284/Y NOR2X1_LOC_492/Y 0.01fF
C10577 D_INPUT_0 NOR2X1_LOC_719/B 0.27fF
C10578 NOR2X1_LOC_561/Y NAND2X1_LOC_140/A 0.02fF
C10579 NOR2X1_LOC_389/B INVX1_LOC_16/A 0.08fF
C10580 NOR2X1_LOC_226/A NOR2X1_LOC_322/Y 0.20fF
C10581 NOR2X1_LOC_188/A INVX1_LOC_266/Y 0.01fF
C10582 NOR2X1_LOC_272/Y NOR2X1_LOC_473/a_36_216# 0.12fF
C10583 D_INPUT_1 NOR2X1_LOC_755/Y 0.02fF
C10584 INVX1_LOC_230/Y INVX1_LOC_230/A 0.07fF
C10585 D_INPUT_1 INVX1_LOC_284/A 0.08fF
C10586 NAND2X1_LOC_140/a_36_24# NOR2X1_LOC_657/B 0.00fF
C10587 INVX1_LOC_5/A NOR2X1_LOC_721/B 0.03fF
C10588 INVX1_LOC_269/A NOR2X1_LOC_809/B 0.03fF
C10589 INVX1_LOC_32/A NAND2X1_LOC_99/A 0.10fF
C10590 INVX1_LOC_23/A NOR2X1_LOC_833/B 0.07fF
C10591 NAND2X1_LOC_360/B INPUT_0 0.01fF
C10592 INVX1_LOC_50/A NOR2X1_LOC_483/a_36_216# 0.00fF
C10593 NOR2X1_LOC_215/Y INVX1_LOC_139/A 0.01fF
C10594 INVX1_LOC_99/A INVX1_LOC_58/Y 0.03fF
C10595 INVX1_LOC_103/A NOR2X1_LOC_364/A 0.14fF
C10596 NOR2X1_LOC_490/Y NOR2X1_LOC_86/A 0.01fF
C10597 NOR2X1_LOC_388/Y NOR2X1_LOC_405/A 0.02fF
C10598 NOR2X1_LOC_369/Y INVX1_LOC_54/A 0.05fF
C10599 NOR2X1_LOC_318/B INVX1_LOC_104/A 0.01fF
C10600 NOR2X1_LOC_808/A NOR2X1_LOC_703/Y 0.12fF
C10601 NOR2X1_LOC_13/Y NAND2X1_LOC_453/A 0.29fF
C10602 NAND2X1_LOC_348/A INVX1_LOC_16/A 0.01fF
C10603 NOR2X1_LOC_789/B INVX1_LOC_293/Y 0.03fF
C10604 NOR2X1_LOC_165/Y INPUT_0 0.01fF
C10605 NAND2X1_LOC_181/Y NOR2X1_LOC_9/Y 0.02fF
C10606 INVX1_LOC_123/A NOR2X1_LOC_537/Y 0.07fF
C10607 NOR2X1_LOC_415/Y INVX1_LOC_175/A 0.10fF
C10608 INVX1_LOC_286/Y INVX1_LOC_54/A 0.10fF
C10609 NOR2X1_LOC_332/A NOR2X1_LOC_112/Y 2.23fF
C10610 INVX1_LOC_104/A INVX1_LOC_93/Y 0.02fF
C10611 NOR2X1_LOC_92/Y INVX1_LOC_63/A 0.14fF
C10612 NOR2X1_LOC_15/Y NOR2X1_LOC_666/a_36_216# 0.00fF
C10613 NOR2X1_LOC_614/Y NOR2X1_LOC_552/Y 0.02fF
C10614 INVX1_LOC_182/Y INVX1_LOC_10/A 0.03fF
C10615 NAND2X1_LOC_329/a_36_24# NOR2X1_LOC_493/B 0.01fF
C10616 INVX1_LOC_286/A NOR2X1_LOC_568/a_36_216# 0.01fF
C10617 NAND2X1_LOC_390/A NOR2X1_LOC_74/A 0.31fF
C10618 NOR2X1_LOC_246/A NOR2X1_LOC_329/B 0.01fF
C10619 NAND2X1_LOC_793/B INVX1_LOC_15/A 0.01fF
C10620 NOR2X1_LOC_789/B NAND2X1_LOC_74/B 0.05fF
C10621 INVX1_LOC_8/A INVX1_LOC_76/A 0.07fF
C10622 INVX1_LOC_309/Y NOR2X1_LOC_536/A -0.00fF
C10623 NAND2X1_LOC_175/B NAND2X1_LOC_453/A 0.05fF
C10624 NAND2X1_LOC_72/B NOR2X1_LOC_748/A 0.03fF
C10625 INVX1_LOC_90/A INVX1_LOC_28/A 0.32fF
C10626 NOR2X1_LOC_103/Y INVX1_LOC_84/A 0.07fF
C10627 NOR2X1_LOC_570/B VDD 0.40fF
C10628 INVX1_LOC_93/A INVX1_LOC_42/A 0.07fF
C10629 INVX1_LOC_1/A INVX1_LOC_19/A 3.29fF
C10630 NOR2X1_LOC_802/A NAND2X1_LOC_280/a_36_24# 0.00fF
C10631 NAND2X1_LOC_341/A NOR2X1_LOC_7/Y 0.20fF
C10632 NAND2X1_LOC_198/B NOR2X1_LOC_351/Y 0.07fF
C10633 INVX1_LOC_21/A NOR2X1_LOC_346/A 0.02fF
C10634 NOR2X1_LOC_52/Y NOR2X1_LOC_358/a_36_216# 0.00fF
C10635 NOR2X1_LOC_97/A NOR2X1_LOC_97/a_36_216# 0.00fF
C10636 INVX1_LOC_159/A INVX1_LOC_54/A 0.07fF
C10637 INVX1_LOC_174/A NOR2X1_LOC_450/B 0.01fF
C10638 INVX1_LOC_83/A NAND2X1_LOC_496/a_36_24# 0.01fF
C10639 NAND2X1_LOC_367/A INVX1_LOC_117/A 0.02fF
C10640 INVX1_LOC_13/A NAND2X1_LOC_4/a_36_24# 0.00fF
C10641 NOR2X1_LOC_723/Y INVX1_LOC_179/A 0.01fF
C10642 NOR2X1_LOC_428/Y NOR2X1_LOC_430/Y 0.23fF
C10643 INVX1_LOC_45/A NOR2X1_LOC_88/Y 0.03fF
C10644 NOR2X1_LOC_620/B NOR2X1_LOC_545/B 0.18fF
C10645 NOR2X1_LOC_322/Y INPUT_1 0.07fF
C10646 INVX1_LOC_3/Y INVX1_LOC_306/Y 0.19fF
C10647 NOR2X1_LOC_357/Y NOR2X1_LOC_423/Y 0.02fF
C10648 NOR2X1_LOC_91/A NOR2X1_LOC_689/Y 0.03fF
C10649 INVX1_LOC_119/A NOR2X1_LOC_681/Y 0.10fF
C10650 INVX1_LOC_119/A INVX1_LOC_37/A 0.31fF
C10651 INVX1_LOC_174/A NOR2X1_LOC_257/Y 0.02fF
C10652 INVX1_LOC_136/A NOR2X1_LOC_831/B 0.03fF
C10653 INVX1_LOC_35/A NOR2X1_LOC_158/Y 0.07fF
C10654 NOR2X1_LOC_186/Y INVX1_LOC_47/Y 0.00fF
C10655 NOR2X1_LOC_554/B NOR2X1_LOC_216/B 0.01fF
C10656 NAND2X1_LOC_819/Y INVX1_LOC_59/Y 0.02fF
C10657 NOR2X1_LOC_504/Y NAND2X1_LOC_453/A 0.01fF
C10658 INVX1_LOC_296/A INVX1_LOC_173/A 0.16fF
C10659 INVX1_LOC_213/Y NAND2X1_LOC_472/Y 0.06fF
C10660 INVX1_LOC_45/A INVX1_LOC_84/A 0.03fF
C10661 NOR2X1_LOC_627/Y INVX1_LOC_139/Y 0.01fF
C10662 NOR2X1_LOC_510/Y INVX1_LOC_21/Y 0.02fF
C10663 INVX1_LOC_164/Y NOR2X1_LOC_266/B 0.00fF
C10664 INVX1_LOC_158/A NAND2X1_LOC_96/A 0.01fF
C10665 INVX1_LOC_255/Y INVX1_LOC_316/A -0.01fF
C10666 NOR2X1_LOC_222/Y NOR2X1_LOC_357/Y 0.10fF
C10667 NOR2X1_LOC_489/B INVX1_LOC_26/A 0.02fF
C10668 INVX1_LOC_151/Y INVX1_LOC_76/A 0.03fF
C10669 INVX1_LOC_233/Y NOR2X1_LOC_693/Y 0.10fF
C10670 NOR2X1_LOC_125/Y INVX1_LOC_23/A 0.43fF
C10671 NOR2X1_LOC_320/Y NOR2X1_LOC_329/B 0.01fF
C10672 NAND2X1_LOC_861/Y NOR2X1_LOC_528/Y 0.10fF
C10673 NAND2X1_LOC_787/Y NAND2X1_LOC_804/A 0.33fF
C10674 INVX1_LOC_30/A NOR2X1_LOC_662/A 0.02fF
C10675 INVX1_LOC_93/A INVX1_LOC_78/A 0.07fF
C10676 INVX1_LOC_36/A NAND2X1_LOC_818/a_36_24# 0.00fF
C10677 NOR2X1_LOC_582/Y NOR2X1_LOC_430/Y 0.18fF
C10678 NAND2X1_LOC_787/A INVX1_LOC_57/A 0.03fF
C10679 NOR2X1_LOC_91/A NAND2X1_LOC_725/A 0.14fF
C10680 INVX1_LOC_21/A INVX1_LOC_94/Y 0.88fF
C10681 NOR2X1_LOC_615/a_36_216# NAND2X1_LOC_254/Y 0.00fF
C10682 INVX1_LOC_278/A INVX1_LOC_224/Y 0.23fF
C10683 NOR2X1_LOC_598/B INVX1_LOC_23/A 0.20fF
C10684 INVX1_LOC_291/Y NAND2X1_LOC_800/Y 0.06fF
C10685 NAND2X1_LOC_363/B INVX1_LOC_57/A 0.04fF
C10686 INVX1_LOC_75/A NOR2X1_LOC_337/A 1.00fF
C10687 INVX1_LOC_45/A NAND2X1_LOC_651/B 0.07fF
C10688 NAND2X1_LOC_717/Y INVX1_LOC_38/A 0.02fF
C10689 NAND2X1_LOC_123/a_36_24# INVX1_LOC_28/A 0.00fF
C10690 INVX1_LOC_215/A VDD 0.00fF
C10691 NOR2X1_LOC_283/a_36_216# NAND2X1_LOC_572/B 0.01fF
C10692 INVX1_LOC_279/A NOR2X1_LOC_850/a_36_216# 0.00fF
C10693 NOR2X1_LOC_742/A INVX1_LOC_206/Y 0.02fF
C10694 INVX1_LOC_71/A INVX1_LOC_84/A 1.47fF
C10695 NOR2X1_LOC_208/Y INVX1_LOC_136/Y 0.01fF
C10696 NOR2X1_LOC_500/B INVX1_LOC_69/A 0.02fF
C10697 INVX1_LOC_278/A NAND2X1_LOC_793/B 0.07fF
C10698 NAND2X1_LOC_513/a_36_24# NAND2X1_LOC_472/Y 0.00fF
C10699 INVX1_LOC_226/Y NOR2X1_LOC_98/B 0.01fF
C10700 INVX1_LOC_89/A NOR2X1_LOC_631/B 0.07fF
C10701 NOR2X1_LOC_644/A INVX1_LOC_65/A 0.03fF
C10702 NAND2X1_LOC_715/B INVX1_LOC_23/A 0.01fF
C10703 INVX1_LOC_144/Y INVX1_LOC_118/A -0.01fF
C10704 NAND2X1_LOC_477/A NOR2X1_LOC_435/A 0.12fF
C10705 INVX1_LOC_286/Y NOR2X1_LOC_48/B 0.07fF
C10706 INVX1_LOC_135/A NOR2X1_LOC_857/A 0.07fF
C10707 INVX1_LOC_21/A INVX1_LOC_296/A 0.58fF
C10708 NOR2X1_LOC_791/Y INVX1_LOC_57/A 0.05fF
C10709 INVX1_LOC_36/A INVX1_LOC_168/Y 0.01fF
C10710 NOR2X1_LOC_813/Y NOR2X1_LOC_86/A 0.04fF
C10711 NOR2X1_LOC_373/Y VDD 0.41fF
C10712 INVX1_LOC_223/A INVX1_LOC_290/Y 0.00fF
C10713 INVX1_LOC_16/A INVX1_LOC_38/A 0.53fF
C10714 INVX1_LOC_90/A NOR2X1_LOC_35/Y 0.05fF
C10715 INVX1_LOC_20/Y INVX1_LOC_20/A 0.01fF
C10716 INVX1_LOC_14/A INVX1_LOC_26/A 0.05fF
C10717 NOR2X1_LOC_513/Y INVX1_LOC_78/A 0.01fF
C10718 NOR2X1_LOC_92/Y NOR2X1_LOC_65/Y 0.01fF
C10719 INVX1_LOC_1/A INVX1_LOC_26/Y 0.09fF
C10720 NOR2X1_LOC_68/A NAND2X1_LOC_200/a_36_24# 0.01fF
C10721 NAND2X1_LOC_363/Y INVX1_LOC_37/A 0.05fF
C10722 INVX1_LOC_181/Y NOR2X1_LOC_89/A 0.07fF
C10723 INVX1_LOC_89/A INVX1_LOC_37/A 6.15fF
C10724 INVX1_LOC_41/A INVX1_LOC_63/A 0.26fF
C10725 INVX1_LOC_136/A NAND2X1_LOC_74/a_36_24# 0.01fF
C10726 INVX1_LOC_45/A INVX1_LOC_15/A 6.61fF
C10727 NAND2X1_LOC_593/Y INVX1_LOC_272/A 0.74fF
C10728 NOR2X1_LOC_219/B INVX1_LOC_186/Y 0.04fF
C10729 INVX1_LOC_269/A NOR2X1_LOC_72/Y 0.06fF
C10730 NOR2X1_LOC_400/a_36_216# INVX1_LOC_14/A 0.01fF
C10731 INVX1_LOC_166/A INVX1_LOC_1/A 0.04fF
C10732 INVX1_LOC_16/A NOR2X1_LOC_51/A 0.00fF
C10733 INVX1_LOC_34/A NAND2X1_LOC_219/B 0.01fF
C10734 NAND2X1_LOC_361/Y INVX1_LOC_125/A 0.05fF
C10735 NOR2X1_LOC_296/Y NAND2X1_LOC_99/A 0.01fF
C10736 NOR2X1_LOC_78/B NAND2X1_LOC_438/a_36_24# 0.00fF
C10737 NAND2X1_LOC_564/A INVX1_LOC_14/A 0.07fF
C10738 NAND2X1_LOC_477/A INVX1_LOC_63/A 0.10fF
C10739 NAND2X1_LOC_348/A NOR2X1_LOC_35/Y 0.05fF
C10740 INVX1_LOC_268/A INVX1_LOC_92/A 0.02fF
C10741 NOR2X1_LOC_172/Y INVX1_LOC_109/A 0.00fF
C10742 NAND2X1_LOC_337/B NAND2X1_LOC_286/B 0.04fF
C10743 NOR2X1_LOC_62/a_36_216# INVX1_LOC_46/Y 0.00fF
C10744 NOR2X1_LOC_356/A INVX1_LOC_117/A 0.09fF
C10745 NAND2X1_LOC_631/a_36_24# INVX1_LOC_284/A 0.00fF
C10746 INVX1_LOC_73/A NOR2X1_LOC_266/B 0.03fF
C10747 NAND2X1_LOC_114/B NOR2X1_LOC_843/B 0.46fF
C10748 INVX1_LOC_286/A NOR2X1_LOC_123/a_36_216# 0.00fF
C10749 NAND2X1_LOC_656/A INVX1_LOC_32/A 0.10fF
C10750 INVX1_LOC_67/Y NOR2X1_LOC_137/Y 0.01fF
C10751 NOR2X1_LOC_736/Y INVX1_LOC_281/A 0.08fF
C10752 INVX1_LOC_71/A INVX1_LOC_15/A 0.21fF
C10753 NAND2X1_LOC_357/B NAND2X1_LOC_74/B 0.07fF
C10754 INVX1_LOC_5/A NAND2X1_LOC_473/A 0.13fF
C10755 NOR2X1_LOC_428/Y INVX1_LOC_296/A 0.17fF
C10756 INVX1_LOC_279/A INVX1_LOC_307/A 0.01fF
C10757 NOR2X1_LOC_803/A NOR2X1_LOC_148/Y 0.03fF
C10758 INVX1_LOC_154/Y VDD 0.26fF
C10759 NAND2X1_LOC_860/A NOR2X1_LOC_786/a_36_216# 0.01fF
C10760 INVX1_LOC_28/A INVX1_LOC_38/A 1.95fF
C10761 NOR2X1_LOC_91/Y NAND2X1_LOC_443/a_36_24# 0.00fF
C10762 NOR2X1_LOC_84/A INVX1_LOC_42/A 0.00fF
C10763 INVX1_LOC_28/A NAND2X1_LOC_264/a_36_24# 0.00fF
C10764 NAND2X1_LOC_840/Y INVX1_LOC_33/Y 0.01fF
C10765 NOR2X1_LOC_52/B NOR2X1_LOC_584/Y 0.04fF
C10766 INVX1_LOC_243/Y INVX1_LOC_30/A 0.06fF
C10767 INVX1_LOC_205/Y INVX1_LOC_21/A 0.01fF
C10768 INVX1_LOC_35/A NOR2X1_LOC_195/A 0.01fF
C10769 NOR2X1_LOC_74/A INVX1_LOC_117/A 0.26fF
C10770 INVX1_LOC_286/A VDD 3.00fF
C10771 NOR2X1_LOC_357/Y NOR2X1_LOC_66/a_36_216# 0.00fF
C10772 INVX1_LOC_269/A INVX1_LOC_50/Y 0.07fF
C10773 INVX1_LOC_243/Y NAND2X1_LOC_763/B 0.25fF
C10774 NOR2X1_LOC_826/Y INVX1_LOC_230/Y 0.01fF
C10775 NOR2X1_LOC_303/Y INVX1_LOC_78/A 0.10fF
C10776 INVX1_LOC_313/A NOR2X1_LOC_155/A 0.03fF
C10777 INVX1_LOC_30/A INVX1_LOC_57/A 0.43fF
C10778 INVX1_LOC_47/A INVX1_LOC_92/A 0.05fF
C10779 NOR2X1_LOC_598/B INVX1_LOC_31/A 0.04fF
C10780 INVX1_LOC_21/A INVX1_LOC_299/A 0.08fF
C10781 INVX1_LOC_54/Y INVX1_LOC_42/A 0.03fF
C10782 NOR2X1_LOC_632/Y NAND2X1_LOC_625/a_36_24# 0.00fF
C10783 INVX1_LOC_225/A INVX1_LOC_47/Y 0.02fF
C10784 INVX1_LOC_178/A NAND2X1_LOC_537/Y 0.10fF
C10785 INVX1_LOC_51/A INVX1_LOC_31/A 0.03fF
C10786 NAND2X1_LOC_557/Y NOR2X1_LOC_384/Y 0.01fF
C10787 NOR2X1_LOC_78/A NOR2X1_LOC_112/a_36_216# 0.00fF
C10788 NAND2X1_LOC_84/Y INVX1_LOC_26/A 0.33fF
C10789 NOR2X1_LOC_360/Y NOR2X1_LOC_383/B 0.01fF
C10790 NOR2X1_LOC_582/Y INVX1_LOC_296/A 0.19fF
C10791 NOR2X1_LOC_67/A NAND2X1_LOC_254/Y 0.08fF
C10792 INVX1_LOC_21/A NOR2X1_LOC_538/B 0.03fF
C10793 INVX1_LOC_155/Y NOR2X1_LOC_334/Y 0.21fF
C10794 INVX1_LOC_94/A INVX1_LOC_28/Y 0.01fF
C10795 D_INPUT_1 INVX1_LOC_72/A 0.57fF
C10796 NOR2X1_LOC_400/A NAND2X1_LOC_555/Y 0.02fF
C10797 NOR2X1_LOC_45/B NOR2X1_LOC_111/A 0.07fF
C10798 INVX1_LOC_101/Y NOR2X1_LOC_348/Y 0.17fF
C10799 INVX1_LOC_278/A INVX1_LOC_45/A 0.15fF
C10800 INVX1_LOC_182/Y INVX1_LOC_307/A 0.02fF
C10801 INVX1_LOC_95/A VDD 0.60fF
C10802 INVX1_LOC_266/A INVX1_LOC_269/A 0.10fF
C10803 INVX1_LOC_120/A NOR2X1_LOC_814/A 0.03fF
C10804 INVX1_LOC_182/A NOR2X1_LOC_197/B 0.10fF
C10805 NOR2X1_LOC_471/Y NOR2X1_LOC_626/Y 0.25fF
C10806 NOR2X1_LOC_357/Y NOR2X1_LOC_69/A 0.02fF
C10807 INVX1_LOC_32/Y NOR2X1_LOC_89/A 0.01fF
C10808 NOR2X1_LOC_381/Y INVX1_LOC_269/A 0.05fF
C10809 NOR2X1_LOC_45/B NOR2X1_LOC_694/Y 0.02fF
C10810 NOR2X1_LOC_770/A NOR2X1_LOC_383/B 0.02fF
C10811 NAND2X1_LOC_35/Y INVX1_LOC_36/A 0.07fF
C10812 INVX1_LOC_104/A INVX1_LOC_87/A 0.08fF
C10813 INVX1_LOC_279/A INVX1_LOC_12/A 0.07fF
C10814 NOR2X1_LOC_536/A NAND2X1_LOC_655/A 0.03fF
C10815 INVX1_LOC_17/A NOR2X1_LOC_523/A 0.00fF
C10816 NOR2X1_LOC_425/a_36_216# NOR2X1_LOC_25/Y 0.00fF
C10817 INVX1_LOC_37/A NAND2X1_LOC_244/A 0.02fF
C10818 NOR2X1_LOC_71/Y NAND2X1_LOC_81/B 0.40fF
C10819 INVX1_LOC_25/A NAND2X1_LOC_119/a_36_24# 0.00fF
C10820 INVX1_LOC_54/Y INVX1_LOC_78/A 0.03fF
C10821 NOR2X1_LOC_717/B INVX1_LOC_99/A 0.01fF
C10822 INVX1_LOC_72/A NOR2X1_LOC_652/Y 0.01fF
C10823 NAND2X1_LOC_537/Y NOR2X1_LOC_816/A 0.57fF
C10824 NAND2X1_LOC_552/A NAND2X1_LOC_640/a_36_24# 0.01fF
C10825 NAND2X1_LOC_803/B INVX1_LOC_103/A 0.03fF
C10826 NOR2X1_LOC_667/A INVX1_LOC_94/Y 0.04fF
C10827 NOR2X1_LOC_128/B NOR2X1_LOC_847/B 0.01fF
C10828 NAND2X1_LOC_125/a_36_24# NOR2X1_LOC_847/A 0.00fF
C10829 INVX1_LOC_6/A NOR2X1_LOC_155/A 0.15fF
C10830 NOR2X1_LOC_612/B INVX1_LOC_26/A 0.35fF
C10831 NOR2X1_LOC_15/Y NOR2X1_LOC_644/B 0.02fF
C10832 INVX1_LOC_226/Y NOR2X1_LOC_38/B 0.13fF
C10833 NOR2X1_LOC_756/Y NAND2X1_LOC_773/B 0.03fF
C10834 INVX1_LOC_249/A NOR2X1_LOC_665/a_36_216# 0.00fF
C10835 NOR2X1_LOC_798/A INVX1_LOC_305/A 0.01fF
C10836 NAND2X1_LOC_724/Y GATE_811 0.03fF
C10837 NOR2X1_LOC_577/Y NOR2X1_LOC_717/A 0.09fF
C10838 INVX1_LOC_17/A INVX1_LOC_174/A 0.08fF
C10839 NOR2X1_LOC_91/A NAND2X1_LOC_660/A 0.07fF
C10840 NOR2X1_LOC_590/A INVX1_LOC_103/A 0.09fF
C10841 NOR2X1_LOC_644/A NOR2X1_LOC_830/Y 0.01fF
C10842 INVX1_LOC_22/A INVX1_LOC_128/Y 0.22fF
C10843 INVX1_LOC_38/A NOR2X1_LOC_35/Y 0.05fF
C10844 NOR2X1_LOC_65/B INVX1_LOC_54/Y 0.67fF
C10845 INVX1_LOC_255/Y INVX1_LOC_4/Y 0.34fF
C10846 NAND2X1_LOC_53/Y NOR2X1_LOC_389/A 0.01fF
C10847 NOR2X1_LOC_56/Y INVX1_LOC_54/A 0.22fF
C10848 INVX1_LOC_224/Y NOR2X1_LOC_63/a_36_216# 0.00fF
C10849 NAND2X1_LOC_555/Y NAND2X1_LOC_19/a_36_24# 0.00fF
C10850 INVX1_LOC_118/Y INVX1_LOC_76/A 0.13fF
C10851 NOR2X1_LOC_794/B NOR2X1_LOC_553/a_36_216# 0.00fF
C10852 INVX1_LOC_304/A NOR2X1_LOC_118/a_36_216# 0.01fF
C10853 INVX1_LOC_36/Y INVX1_LOC_9/A 0.07fF
C10854 NOR2X1_LOC_773/Y NAND2X1_LOC_286/B 0.01fF
C10855 INVX1_LOC_50/A NOR2X1_LOC_352/Y 0.00fF
C10856 VDD NOR2X1_LOC_602/B -0.00fF
C10857 INVX1_LOC_182/Y INVX1_LOC_12/A 0.03fF
C10858 INVX1_LOC_95/Y INVX1_LOC_92/A 0.10fF
C10859 NOR2X1_LOC_348/B NOR2X1_LOC_717/A 0.03fF
C10860 NOR2X1_LOC_514/Y NOR2X1_LOC_660/Y 0.01fF
C10861 NOR2X1_LOC_71/Y NAND2X1_LOC_269/a_36_24# 0.01fF
C10862 NOR2X1_LOC_590/A INVX1_LOC_292/A 0.16fF
C10863 NOR2X1_LOC_740/Y INVX1_LOC_142/A 0.07fF
C10864 NOR2X1_LOC_188/A INVX1_LOC_19/A 0.20fF
C10865 NAND2X1_LOC_96/A NAND2X1_LOC_825/a_36_24# 0.01fF
C10866 D_INPUT_1 NAND2X1_LOC_338/B 0.15fF
C10867 NOR2X1_LOC_372/A INVX1_LOC_31/A 0.09fF
C10868 VDD INVX1_LOC_54/A 1.49fF
C10869 NOR2X1_LOC_548/B INVX1_LOC_19/A 0.07fF
C10870 NAND2X1_LOC_579/A INVX1_LOC_24/A 0.10fF
C10871 NOR2X1_LOC_269/Y NOR2X1_LOC_127/Y 0.06fF
C10872 INVX1_LOC_196/A INVX1_LOC_53/A 0.03fF
C10873 INVX1_LOC_78/Y INVX1_LOC_186/Y 0.00fF
C10874 NOR2X1_LOC_75/Y NOR2X1_LOC_722/Y 0.00fF
C10875 INVX1_LOC_92/Y NAND2X1_LOC_63/Y 0.04fF
C10876 NOR2X1_LOC_121/A NOR2X1_LOC_646/B 0.01fF
C10877 NOR2X1_LOC_305/Y INVX1_LOC_92/A 0.07fF
C10878 INVX1_LOC_194/A INVX1_LOC_253/Y 0.20fF
C10879 INVX1_LOC_286/Y NOR2X1_LOC_441/Y 0.07fF
C10880 NOR2X1_LOC_329/B INVX1_LOC_32/A 0.01fF
C10881 NOR2X1_LOC_91/Y NAND2X1_LOC_793/Y 0.01fF
C10882 INVX1_LOC_21/A INVX1_LOC_162/A 0.03fF
C10883 NAND2X1_LOC_149/Y INVX1_LOC_33/A 0.07fF
C10884 INVX1_LOC_11/A INVX1_LOC_181/Y 0.03fF
C10885 INVX1_LOC_122/Y NOR2X1_LOC_160/B 0.63fF
C10886 INVX1_LOC_136/A NAND2X1_LOC_352/B 0.11fF
C10887 INVX1_LOC_89/A NAND2X1_LOC_72/B 0.03fF
C10888 NOR2X1_LOC_541/Y NOR2X1_LOC_168/Y 0.02fF
C10889 NOR2X1_LOC_163/Y D_INPUT_5 0.01fF
C10890 NOR2X1_LOC_287/A INVX1_LOC_53/A 0.04fF
C10891 NAND2X1_LOC_53/Y NOR2X1_LOC_596/A 0.46fF
C10892 NOR2X1_LOC_542/B NOR2X1_LOC_814/A 0.25fF
C10893 NOR2X1_LOC_329/B NOR2X1_LOC_329/Y 0.15fF
C10894 NOR2X1_LOC_533/Y NAND2X1_LOC_567/Y 0.01fF
C10895 INVX1_LOC_21/A NOR2X1_LOC_315/Y 0.17fF
C10896 NOR2X1_LOC_43/Y INVX1_LOC_19/A 0.42fF
C10897 INVX1_LOC_268/A INVX1_LOC_53/A 0.03fF
C10898 INVX1_LOC_141/Y INVX1_LOC_18/A 0.03fF
C10899 INVX1_LOC_22/A NOR2X1_LOC_717/A 0.43fF
C10900 NOR2X1_LOC_513/Y NOR2X1_LOC_152/Y 0.03fF
C10901 INPUT_3 NAND2X1_LOC_656/A 0.10fF
C10902 INVX1_LOC_48/Y NOR2X1_LOC_392/B 0.10fF
C10903 NAND2X1_LOC_453/A NOR2X1_LOC_697/Y 0.02fF
C10904 INVX1_LOC_14/A INVX1_LOC_315/A 0.07fF
C10905 NOR2X1_LOC_329/B NAND2X1_LOC_175/Y 0.16fF
C10906 NOR2X1_LOC_242/A INVX1_LOC_196/A 0.09fF
C10907 INVX1_LOC_35/A INVX1_LOC_13/A 0.13fF
C10908 NOR2X1_LOC_865/Y INVX1_LOC_117/A 0.66fF
C10909 INVX1_LOC_103/A NAND2X1_LOC_354/B 0.12fF
C10910 INVX1_LOC_5/A INVX1_LOC_172/Y 0.01fF
C10911 INVX1_LOC_269/A NOR2X1_LOC_6/B 0.11fF
C10912 INVX1_LOC_31/A NOR2X1_LOC_513/a_36_216# 0.00fF
C10913 NOR2X1_LOC_168/Y NOR2X1_LOC_568/A -0.03fF
C10914 NOR2X1_LOC_471/Y INVX1_LOC_153/A 0.01fF
C10915 INVX1_LOC_2/A NOR2X1_LOC_669/a_36_216# 0.00fF
C10916 NOR2X1_LOC_768/a_36_216# INVX1_LOC_270/A 0.01fF
C10917 NOR2X1_LOC_75/Y INVX1_LOC_34/A 0.03fF
C10918 NOR2X1_LOC_128/B NOR2X1_LOC_660/Y 0.29fF
C10919 NOR2X1_LOC_83/Y NOR2X1_LOC_80/Y 0.40fF
C10920 NOR2X1_LOC_635/A NAND2X1_LOC_583/a_36_24# 0.00fF
C10921 NOR2X1_LOC_669/a_36_216# NOR2X1_LOC_226/A 0.13fF
C10922 NOR2X1_LOC_91/A NAND2X1_LOC_560/A 0.06fF
C10923 INVX1_LOC_178/A INVX1_LOC_172/Y 0.01fF
C10924 NOR2X1_LOC_160/B NOR2X1_LOC_561/a_36_216# 0.01fF
C10925 INVX1_LOC_230/Y NOR2X1_LOC_690/A 0.00fF
C10926 INVX1_LOC_278/A NOR2X1_LOC_123/B 0.02fF
C10927 D_INPUT_1 INVX1_LOC_313/Y 0.02fF
C10928 INVX1_LOC_223/A INVX1_LOC_77/A 0.03fF
C10929 INVX1_LOC_58/A NOR2X1_LOC_356/A 0.03fF
C10930 INVX1_LOC_35/A NOR2X1_LOC_246/A 0.07fF
C10931 INVX1_LOC_230/Y NOR2X1_LOC_413/Y 0.01fF
C10932 NOR2X1_LOC_567/B NOR2X1_LOC_383/B 0.07fF
C10933 NOR2X1_LOC_16/Y NOR2X1_LOC_103/Y 0.10fF
C10934 NOR2X1_LOC_56/Y NOR2X1_LOC_48/B 0.05fF
C10935 INVX1_LOC_35/A NOR2X1_LOC_174/B 0.32fF
C10936 NOR2X1_LOC_632/Y INVX1_LOC_27/A 0.01fF
C10937 INVX1_LOC_45/A NAND2X1_LOC_21/Y 0.02fF
C10938 NOR2X1_LOC_135/Y INVX1_LOC_271/A 0.00fF
C10939 NOR2X1_LOC_331/B INVX1_LOC_84/A 0.07fF
C10940 NOR2X1_LOC_155/A INVX1_LOC_131/Y 0.81fF
C10941 INVX1_LOC_176/A NOR2X1_LOC_67/Y 0.13fF
C10942 INVX1_LOC_47/Y NAND2X1_LOC_642/Y 0.10fF
C10943 INVX1_LOC_35/A NAND2X1_LOC_551/A 0.07fF
C10944 NOR2X1_LOC_381/Y NAND2X1_LOC_563/A 0.17fF
C10945 NOR2X1_LOC_168/Y INVX1_LOC_71/A 0.01fF
C10946 NOR2X1_LOC_188/A INVX1_LOC_26/Y 0.10fF
C10947 NOR2X1_LOC_454/Y NAND2X1_LOC_662/Y 0.07fF
C10948 NAND2X1_LOC_51/B INVX1_LOC_296/A 0.02fF
C10949 VDD NAND2X1_LOC_807/B 0.36fF
C10950 NAND2X1_LOC_725/A NAND2X1_LOC_866/B 0.10fF
C10951 NOR2X1_LOC_548/B INVX1_LOC_26/Y 0.92fF
C10952 INVX1_LOC_18/A INVX1_LOC_275/A 0.05fF
C10953 NOR2X1_LOC_546/A NOR2X1_LOC_550/B 0.05fF
C10954 INVX1_LOC_48/A INVX1_LOC_26/A 0.02fF
C10955 NAND2X1_LOC_323/B NOR2X1_LOC_241/A 0.01fF
C10956 NAND2X1_LOC_540/a_36_24# NOR2X1_LOC_71/Y 0.00fF
C10957 NAND2X1_LOC_53/Y NOR2X1_LOC_220/A 0.10fF
C10958 INVX1_LOC_181/Y NOR2X1_LOC_433/A 0.15fF
C10959 NOR2X1_LOC_814/Y INVX1_LOC_50/Y 0.08fF
C10960 VDD NOR2X1_LOC_48/B 3.18fF
C10961 NOR2X1_LOC_264/a_36_216# INVX1_LOC_30/Y 0.00fF
C10962 INVX1_LOC_58/A NOR2X1_LOC_74/A 0.29fF
C10963 NOR2X1_LOC_68/A INVX1_LOC_63/Y 0.13fF
C10964 NAND2X1_LOC_594/a_36_24# NOR2X1_LOC_130/A 0.01fF
C10965 NOR2X1_LOC_846/B INVX1_LOC_38/Y 0.10fF
C10966 NOR2X1_LOC_13/Y NOR2X1_LOC_577/Y 0.10fF
C10967 INVX1_LOC_188/A NOR2X1_LOC_78/B 0.04fF
C10968 INVX1_LOC_215/A NOR2X1_LOC_361/B 0.78fF
C10969 INVX1_LOC_289/Y NAND2X1_LOC_854/B 0.08fF
C10970 NOR2X1_LOC_332/A NAND2X1_LOC_473/A 0.05fF
C10971 NOR2X1_LOC_303/Y INVX1_LOC_113/Y 0.00fF
C10972 INVX1_LOC_136/A NAND2X1_LOC_357/B 1.18fF
C10973 NAND2X1_LOC_794/B INVX1_LOC_90/A 0.01fF
C10974 INVX1_LOC_38/A INVX1_LOC_109/A 0.08fF
C10975 NOR2X1_LOC_78/A INVX1_LOC_23/Y 0.07fF
C10976 NOR2X1_LOC_42/a_36_216# INVX1_LOC_32/A 0.01fF
C10977 NAND2X1_LOC_785/B NOR2X1_LOC_482/Y 0.09fF
C10978 INVX1_LOC_17/A NOR2X1_LOC_589/A 0.07fF
C10979 INVX1_LOC_6/A NOR2X1_LOC_125/Y 0.07fF
C10980 NAND2X1_LOC_468/B NAND2X1_LOC_470/B 0.07fF
C10981 INVX1_LOC_58/A NOR2X1_LOC_9/Y 0.08fF
C10982 INVX1_LOC_224/Y INVX1_LOC_123/A 0.02fF
C10983 NOR2X1_LOC_283/a_36_216# NOR2X1_LOC_716/B 0.00fF
C10984 NOR2X1_LOC_194/a_36_216# INVX1_LOC_266/Y 0.01fF
C10985 VDD NAND2X1_LOC_3/B 0.30fF
C10986 NAND2X1_LOC_141/Y INVX1_LOC_3/A 0.05fF
C10987 INVX1_LOC_181/Y NOR2X1_LOC_52/B 0.03fF
C10988 NOR2X1_LOC_68/A NOR2X1_LOC_175/A 0.05fF
C10989 NOR2X1_LOC_168/B INVX1_LOC_18/A 0.07fF
C10990 NOR2X1_LOC_471/Y NOR2X1_LOC_589/A 0.14fF
C10991 INVX1_LOC_2/A NOR2X1_LOC_457/B 0.07fF
C10992 INVX1_LOC_77/A INVX1_LOC_149/Y 0.37fF
C10993 INVX1_LOC_304/A INVX1_LOC_181/A 0.02fF
C10994 INVX1_LOC_34/A NOR2X1_LOC_716/B 0.07fF
C10995 NOR2X1_LOC_372/A NAND2X1_LOC_859/Y 0.11fF
C10996 NOR2X1_LOC_382/Y INVX1_LOC_316/Y 0.80fF
C10997 NOR2X1_LOC_301/A INVX1_LOC_20/A 0.03fF
C10998 INVX1_LOC_36/A INVX1_LOC_56/A 0.01fF
C10999 NOR2X1_LOC_820/B NOR2X1_LOC_649/B 0.04fF
C11000 NOR2X1_LOC_155/A INVX1_LOC_301/A 0.18fF
C11001 NOR2X1_LOC_435/B INVX1_LOC_63/A 0.15fF
C11002 INVX1_LOC_17/A INVX1_LOC_171/A 0.07fF
C11003 NOR2X1_LOC_658/Y INVX1_LOC_22/A 0.02fF
C11004 NAND2X1_LOC_555/Y NAND2X1_LOC_377/Y 0.02fF
C11005 NOR2X1_LOC_458/Y NOR2X1_LOC_570/B 0.14fF
C11006 INVX1_LOC_227/A INVX1_LOC_292/A 0.71fF
C11007 NOR2X1_LOC_445/Y NOR2X1_LOC_388/Y 0.00fF
C11008 NAND2X1_LOC_550/A NOR2X1_LOC_525/Y 0.00fF
C11009 NAND2X1_LOC_464/A INVX1_LOC_23/Y 0.00fF
C11010 INVX1_LOC_257/A INVX1_LOC_193/A 0.01fF
C11011 NOR2X1_LOC_331/B INVX1_LOC_15/A 0.60fF
C11012 NOR2X1_LOC_389/A INVX1_LOC_10/A 0.10fF
C11013 NAND2X1_LOC_463/B INVX1_LOC_242/A 0.01fF
C11014 NAND2X1_LOC_16/a_36_24# NOR2X1_LOC_589/A 0.00fF
C11015 NOR2X1_LOC_403/B NAND2X1_LOC_338/B 0.05fF
C11016 VDD NOR2X1_LOC_438/Y 0.66fF
C11017 NAND2X1_LOC_303/Y NAND2X1_LOC_740/B 0.17fF
C11018 INVX1_LOC_48/Y NAND2X1_LOC_348/A 0.01fF
C11019 NAND2X1_LOC_537/Y INVX1_LOC_140/A 0.10fF
C11020 NOR2X1_LOC_414/a_36_216# INVX1_LOC_7/A 0.00fF
C11021 NAND2X1_LOC_350/A INVX1_LOC_190/Y 0.01fF
C11022 NAND2X1_LOC_229/a_36_24# INVX1_LOC_314/Y 0.00fF
C11023 INVX1_LOC_226/Y INVX1_LOC_62/Y 0.01fF
C11024 NOR2X1_LOC_590/A INVX1_LOC_120/A 0.01fF
C11025 INVX1_LOC_90/A INVX1_LOC_246/A 0.03fF
C11026 INVX1_LOC_95/Y INVX1_LOC_53/A 0.01fF
C11027 INVX1_LOC_35/Y INVX1_LOC_42/A -0.01fF
C11028 INVX1_LOC_2/A NAND2X1_LOC_833/Y 0.07fF
C11029 NOR2X1_LOC_570/B INVX1_LOC_177/A 0.03fF
C11030 NOR2X1_LOC_810/A NOR2X1_LOC_354/B 0.01fF
C11031 NAND2X1_LOC_182/A NAND2X1_LOC_180/a_36_24# 0.02fF
C11032 NOR2X1_LOC_13/Y INVX1_LOC_22/A 0.07fF
C11033 NAND2X1_LOC_79/Y NOR2X1_LOC_719/A 0.03fF
C11034 NOR2X1_LOC_226/A NAND2X1_LOC_833/Y 0.00fF
C11035 INVX1_LOC_72/A NOR2X1_LOC_747/a_36_216# 0.00fF
C11036 INVX1_LOC_100/Y NAND2X1_LOC_474/Y 0.03fF
C11037 INVX1_LOC_119/A NAND2X1_LOC_239/a_36_24# 0.03fF
C11038 NAND2X1_LOC_656/Y INVX1_LOC_18/A 0.01fF
C11039 NOR2X1_LOC_592/B INVX1_LOC_15/A 0.28fF
C11040 NAND2X1_LOC_125/a_36_24# NOR2X1_LOC_554/B 0.00fF
C11041 NOR2X1_LOC_300/Y INVX1_LOC_266/Y 0.02fF
C11042 INVX1_LOC_292/A NOR2X1_LOC_703/A 0.19fF
C11043 NOR2X1_LOC_309/Y NOR2X1_LOC_312/a_36_216# 0.01fF
C11044 INVX1_LOC_53/A NOR2X1_LOC_305/Y 0.07fF
C11045 INVX1_LOC_249/A NOR2X1_LOC_632/Y 0.02fF
C11046 INVX1_LOC_34/A NOR2X1_LOC_757/Y 0.09fF
C11047 NOR2X1_LOC_596/A INVX1_LOC_10/A 0.09fF
C11048 NAND2X1_LOC_647/B NOR2X1_LOC_831/B 0.02fF
C11049 INVX1_LOC_200/A NAND2X1_LOC_858/B 0.03fF
C11050 INVX1_LOC_33/A INVX1_LOC_16/A 2.40fF
C11051 NOR2X1_LOC_361/B INVX1_LOC_286/A 0.10fF
C11052 NOR2X1_LOC_721/B INVX1_LOC_42/A 0.28fF
C11053 NOR2X1_LOC_573/Y NAND2X1_LOC_463/B 0.01fF
C11054 INVX1_LOC_90/A NAND2X1_LOC_272/a_36_24# 0.01fF
C11055 INVX1_LOC_41/A INVX1_LOC_1/Y 0.07fF
C11056 INVX1_LOC_106/A NAND2X1_LOC_63/Y 0.01fF
C11057 NOR2X1_LOC_493/B NAND2X1_LOC_491/a_36_24# 0.02fF
C11058 NAND2X1_LOC_114/B NOR2X1_LOC_185/a_36_216# 0.00fF
C11059 INVX1_LOC_133/A NAND2X1_LOC_807/B 0.18fF
C11060 NAND2X1_LOC_213/A NOR2X1_LOC_45/B 0.02fF
C11061 NOR2X1_LOC_801/A NOR2X1_LOC_801/B 0.01fF
C11062 NAND2X1_LOC_562/B INVX1_LOC_172/Y 0.02fF
C11063 NAND2X1_LOC_717/Y NAND2X1_LOC_852/a_36_24# 0.00fF
C11064 INVX1_LOC_196/A NOR2X1_LOC_634/B 0.16fF
C11065 NOR2X1_LOC_92/Y INVX1_LOC_93/Y 0.07fF
C11066 INVX1_LOC_227/A INVX1_LOC_67/A 0.14fF
C11067 NAND2X1_LOC_338/B NOR2X1_LOC_620/B 0.05fF
C11068 NOR2X1_LOC_226/A INVX1_LOC_164/Y 0.03fF
C11069 INVX1_LOC_45/A NOR2X1_LOC_310/a_36_216# 0.00fF
C11070 INVX1_LOC_35/A INVX1_LOC_66/Y 0.06fF
C11071 INVX1_LOC_136/A NAND2X1_LOC_849/A 0.08fF
C11072 NOR2X1_LOC_227/A NOR2X1_LOC_814/A 0.10fF
C11073 NOR2X1_LOC_568/A NOR2X1_LOC_310/a_36_216# 0.01fF
C11074 NOR2X1_LOC_653/B NAND2X1_LOC_287/B 0.03fF
C11075 NOR2X1_LOC_89/a_36_216# NAND2X1_LOC_477/Y 0.00fF
C11076 INVX1_LOC_223/Y INVX1_LOC_37/A 0.31fF
C11077 INVX1_LOC_36/A INVX1_LOC_144/A 0.07fF
C11078 INVX1_LOC_27/A NAND2X1_LOC_39/Y 0.04fF
C11079 NOR2X1_LOC_78/B NAND2X1_LOC_841/A 0.01fF
C11080 NOR2X1_LOC_607/Y INVX1_LOC_313/Y 0.03fF
C11081 INVX1_LOC_208/A NOR2X1_LOC_757/a_36_216# 0.01fF
C11082 NOR2X1_LOC_295/Y INVX1_LOC_10/A 0.03fF
C11083 NOR2X1_LOC_361/B INVX1_LOC_95/A 0.06fF
C11084 INVX1_LOC_90/A NOR2X1_LOC_350/A 0.04fF
C11085 INVX1_LOC_31/A INVX1_LOC_201/A 0.03fF
C11086 NOR2X1_LOC_68/A INVX1_LOC_302/Y 0.03fF
C11087 INVX1_LOC_256/A NOR2X1_LOC_139/Y 0.14fF
C11088 INVX1_LOC_36/A NOR2X1_LOC_83/Y 0.01fF
C11089 NOR2X1_LOC_180/B INVX1_LOC_49/A 0.47fF
C11090 INVX1_LOC_232/Y NOR2X1_LOC_516/B 0.22fF
C11091 NOR2X1_LOC_220/A NOR2X1_LOC_500/Y 0.10fF
C11092 NOR2X1_LOC_155/A INVX1_LOC_270/A 0.03fF
C11093 NAND2X1_LOC_574/A NAND2X1_LOC_223/B 0.06fF
C11094 NOR2X1_LOC_186/Y INVX1_LOC_33/Y 0.26fF
C11095 INVX1_LOC_89/A INVX1_LOC_310/Y 0.04fF
C11096 NOR2X1_LOC_817/Y INVX1_LOC_316/A 0.03fF
C11097 NAND2X1_LOC_541/Y INVX1_LOC_232/A 0.01fF
C11098 NAND2X1_LOC_833/Y INPUT_1 0.02fF
C11099 INVX1_LOC_13/Y NOR2X1_LOC_536/A 0.17fF
C11100 INVX1_LOC_34/A NOR2X1_LOC_130/Y 0.03fF
C11101 INVX1_LOC_21/A NAND2X1_LOC_96/A 0.08fF
C11102 INVX1_LOC_40/A INVX1_LOC_16/A 2.20fF
C11103 NAND2X1_LOC_584/a_36_24# NOR2X1_LOC_763/Y 0.00fF
C11104 NOR2X1_LOC_568/A NOR2X1_LOC_548/a_36_216# 0.01fF
C11105 INVX1_LOC_256/A NAND2X1_LOC_468/B 0.03fF
C11106 NAND2X1_LOC_726/Y INVX1_LOC_16/A 0.01fF
C11107 INVX1_LOC_12/A NOR2X1_LOC_38/B 0.06fF
C11108 INVX1_LOC_33/A INVX1_LOC_28/A 0.10fF
C11109 NOR2X1_LOC_58/Y INVX1_LOC_23/A 0.04fF
C11110 INVX1_LOC_17/A INVX1_LOC_20/A 0.02fF
C11111 NOR2X1_LOC_92/Y NAND2X1_LOC_721/A 0.12fF
C11112 NOR2X1_LOC_381/Y NOR2X1_LOC_37/a_36_216# 0.00fF
C11113 INVX1_LOC_11/A INVX1_LOC_115/A 0.12fF
C11114 NAND2X1_LOC_350/A NOR2X1_LOC_56/Y 0.17fF
C11115 NAND2X1_LOC_794/B INVX1_LOC_38/A 3.82fF
C11116 NAND2X1_LOC_573/Y INVX1_LOC_33/Y 0.02fF
C11117 INVX1_LOC_17/A NOR2X1_LOC_360/A 0.03fF
C11118 INVX1_LOC_18/A INVX1_LOC_78/Y 0.03fF
C11119 NOR2X1_LOC_500/Y NOR2X1_LOC_548/Y 0.00fF
C11120 INVX1_LOC_83/A INVX1_LOC_196/A 0.03fF
C11121 NOR2X1_LOC_367/B D_GATE_366 0.01fF
C11122 INVX1_LOC_13/A NOR2X1_LOC_121/A 0.21fF
C11123 INVX1_LOC_24/A NOR2X1_LOC_387/A 0.00fF
C11124 INVX1_LOC_272/Y NOR2X1_LOC_447/B 0.00fF
C11125 INVX1_LOC_23/A NAND2X1_LOC_606/a_36_24# 0.00fF
C11126 NOR2X1_LOC_772/B NAND2X1_LOC_93/B 0.07fF
C11127 NOR2X1_LOC_419/Y INPUT_0 0.05fF
C11128 NAND2X1_LOC_724/A INVX1_LOC_33/Y 0.07fF
C11129 NOR2X1_LOC_235/a_36_216# NOR2X1_LOC_813/Y 0.01fF
C11130 INVX1_LOC_267/Y INVX1_LOC_89/A 0.01fF
C11131 NOR2X1_LOC_730/Y NOR2X1_LOC_687/Y 0.11fF
C11132 INVX1_LOC_41/A NOR2X1_LOC_742/A 0.76fF
C11133 NOR2X1_LOC_510/Y INVX1_LOC_54/A 0.64fF
C11134 NOR2X1_LOC_278/a_36_216# NAND2X1_LOC_181/Y 0.00fF
C11135 NOR2X1_LOC_727/B INVX1_LOC_186/Y 0.13fF
C11136 NOR2X1_LOC_590/A INVX1_LOC_143/Y 0.01fF
C11137 INVX1_LOC_90/A INVX1_LOC_216/A 0.03fF
C11138 NAND2X1_LOC_350/A VDD -0.00fF
C11139 NOR2X1_LOC_226/A NOR2X1_LOC_76/A 0.01fF
C11140 NOR2X1_LOC_716/B INPUT_0 0.14fF
C11141 INVX1_LOC_71/A NOR2X1_LOC_548/a_36_216# 0.00fF
C11142 NOR2X1_LOC_287/A INVX1_LOC_83/A 0.00fF
C11143 INVX1_LOC_13/Y NAND2X1_LOC_93/B 0.05fF
C11144 INVX1_LOC_88/A NOR2X1_LOC_536/A 0.05fF
C11145 NOR2X1_LOC_91/A INVX1_LOC_29/A 0.06fF
C11146 INVX1_LOC_164/Y INPUT_1 0.01fF
C11147 NOR2X1_LOC_201/A INVX1_LOC_29/A 0.01fF
C11148 NOR2X1_LOC_612/Y NOR2X1_LOC_440/B 0.03fF
C11149 INVX1_LOC_218/Y VDD 0.22fF
C11150 INVX1_LOC_50/A INVX1_LOC_125/A 0.07fF
C11151 INVX1_LOC_245/Y INVX1_LOC_117/A 0.03fF
C11152 NOR2X1_LOC_441/Y VDD 0.92fF
C11153 NOR2X1_LOC_191/A NAND2X1_LOC_842/B 0.09fF
C11154 INVX1_LOC_35/A NAND2X1_LOC_489/Y 0.03fF
C11155 NAND2X1_LOC_348/A NOR2X1_LOC_84/Y 0.00fF
C11156 INVX1_LOC_49/Y NOR2X1_LOC_591/A 0.22fF
C11157 NAND2X1_LOC_359/Y NAND2X1_LOC_348/A 0.04fF
C11158 NOR2X1_LOC_163/Y NAND2X1_LOC_451/Y 0.07fF
C11159 INVX1_LOC_23/A INVX1_LOC_29/A 4.83fF
C11160 NAND2X1_LOC_13/a_36_24# INVX1_LOC_9/A 0.00fF
C11161 NOR2X1_LOC_82/A NOR2X1_LOC_119/a_36_216# 0.00fF
C11162 NOR2X1_LOC_220/A NOR2X1_LOC_302/Y 0.03fF
C11163 NOR2X1_LOC_621/B INVX1_LOC_15/A 0.04fF
C11164 INVX1_LOC_28/A INVX1_LOC_165/Y 0.02fF
C11165 INVX1_LOC_90/A INVX1_LOC_290/A 0.01fF
C11166 NAND2X1_LOC_726/Y INVX1_LOC_28/A 0.02fF
C11167 NOR2X1_LOC_226/A INVX1_LOC_73/A 0.08fF
C11168 INVX1_LOC_246/A INVX1_LOC_38/A 0.07fF
C11169 NOR2X1_LOC_449/A INVX1_LOC_15/A 0.04fF
C11170 NOR2X1_LOC_238/Y NOR2X1_LOC_164/Y 0.00fF
C11171 NOR2X1_LOC_520/B NOR2X1_LOC_557/A 0.18fF
C11172 NOR2X1_LOC_598/B NOR2X1_LOC_633/A 0.01fF
C11173 INVX1_LOC_13/Y INVX1_LOC_3/A 0.14fF
C11174 INVX1_LOC_9/Y NOR2X1_LOC_329/B 0.09fF
C11175 INVX1_LOC_88/A NAND2X1_LOC_93/B 0.03fF
C11176 NAND2X1_LOC_190/Y INVX1_LOC_307/A 0.02fF
C11177 NOR2X1_LOC_605/B INVX1_LOC_28/A 0.01fF
C11178 NOR2X1_LOC_432/Y INVX1_LOC_311/A 0.06fF
C11179 NAND2X1_LOC_357/A NOR2X1_LOC_743/Y 0.01fF
C11180 INVX1_LOC_208/A NOR2X1_LOC_218/a_36_216# 0.00fF
C11181 NOR2X1_LOC_445/Y NOR2X1_LOC_552/A 0.09fF
C11182 NOR2X1_LOC_513/Y INVX1_LOC_291/A 0.02fF
C11183 NOR2X1_LOC_459/A INVX1_LOC_175/Y 0.02fF
C11184 INVX1_LOC_41/A INVX1_LOC_93/Y 0.01fF
C11185 NAND2X1_LOC_363/Y NAND2X1_LOC_367/B 0.00fF
C11186 NAND2X1_LOC_860/A INVX1_LOC_42/A 0.01fF
C11187 INVX1_LOC_256/Y INVX1_LOC_100/A 0.07fF
C11188 INVX1_LOC_135/A NOR2X1_LOC_542/Y 0.07fF
C11189 NOR2X1_LOC_238/Y INVX1_LOC_46/A 0.01fF
C11190 NOR2X1_LOC_750/A INVX1_LOC_7/A 0.01fF
C11191 INVX1_LOC_314/Y NOR2X1_LOC_558/A 0.01fF
C11192 D_INPUT_4 GATE_662 0.03fF
C11193 NOR2X1_LOC_39/Y INVX1_LOC_4/Y 0.08fF
C11194 INVX1_LOC_89/A NOR2X1_LOC_507/B 0.03fF
C11195 NOR2X1_LOC_750/a_36_216# INVX1_LOC_7/A 0.00fF
C11196 NAND2X1_LOC_721/A NAND2X1_LOC_837/Y 0.10fF
C11197 INVX1_LOC_33/A NOR2X1_LOC_35/Y 0.01fF
C11198 INVX1_LOC_223/A INVX1_LOC_9/A 0.59fF
C11199 INVX1_LOC_226/Y INVX1_LOC_51/Y 0.03fF
C11200 NAND2X1_LOC_714/B INVX1_LOC_264/A 0.18fF
C11201 INVX1_LOC_30/A INVX1_LOC_274/A 0.07fF
C11202 NOR2X1_LOC_762/a_36_216# NOR2X1_LOC_11/Y 0.00fF
C11203 NOR2X1_LOC_334/Y NOR2X1_LOC_858/A 0.01fF
C11204 NOR2X1_LOC_581/a_36_216# NOR2X1_LOC_11/Y 0.00fF
C11205 INVX1_LOC_35/A INVX1_LOC_32/A 0.16fF
C11206 NOR2X1_LOC_91/A NOR2X1_LOC_281/Y 0.03fF
C11207 INVX1_LOC_41/A NAND2X1_LOC_641/a_36_24# 0.00fF
C11208 NOR2X1_LOC_364/a_36_216# INVX1_LOC_63/Y 0.01fF
C11209 NOR2X1_LOC_592/a_36_216# NOR2X1_LOC_697/Y 0.00fF
C11210 NAND2X1_LOC_326/A INVX1_LOC_19/A 0.02fF
C11211 NOR2X1_LOC_340/Y VDD 0.37fF
C11212 NOR2X1_LOC_142/Y VDD 2.04fF
C11213 INVX1_LOC_35/A NOR2X1_LOC_623/B 0.06fF
C11214 INVX1_LOC_26/A NOR2X1_LOC_383/B 0.07fF
C11215 NAND2X1_LOC_347/B NAND2X1_LOC_74/B 0.02fF
C11216 NOR2X1_LOC_510/Y NOR2X1_LOC_48/B 0.08fF
C11217 NAND2X1_LOC_866/B NAND2X1_LOC_560/A 0.08fF
C11218 NAND2X1_LOC_508/A NAND2X1_LOC_506/a_36_24# 0.02fF
C11219 NOR2X1_LOC_717/B INPUT_0 0.03fF
C11220 NOR2X1_LOC_78/B INVX1_LOC_95/Y 6.21fF
C11221 INVX1_LOC_53/A INVX1_LOC_271/Y 0.02fF
C11222 INVX1_LOC_36/A NOR2X1_LOC_155/A 0.03fF
C11223 NAND2X1_LOC_860/A INVX1_LOC_78/A 0.00fF
C11224 NAND2X1_LOC_858/B NAND2X1_LOC_808/A 0.03fF
C11225 INVX1_LOC_242/A INVX1_LOC_42/A 0.20fF
C11226 NOR2X1_LOC_78/A INVX1_LOC_232/A 0.16fF
C11227 INVX1_LOC_73/A INPUT_1 1.09fF
C11228 NOR2X1_LOC_189/A INVX1_LOC_38/A 0.45fF
C11229 NOR2X1_LOC_795/Y NOR2X1_LOC_857/A 0.10fF
C11230 INVX1_LOC_298/Y INVX1_LOC_23/A 0.02fF
C11231 INVX1_LOC_271/A NAND2X1_LOC_61/Y 0.26fF
C11232 NAND2X1_LOC_563/A NOR2X1_LOC_124/A 0.04fF
C11233 INVX1_LOC_62/A NOR2X1_LOC_188/A 0.02fF
C11234 INVX1_LOC_64/A NOR2X1_LOC_158/B 0.01fF
C11235 NAND2X1_LOC_477/A NAND2X1_LOC_641/a_36_24# 0.06fF
C11236 NOR2X1_LOC_468/Y INVX1_LOC_12/A 0.19fF
C11237 INVX1_LOC_286/A NAND2X1_LOC_573/A 0.02fF
C11238 NAND2X1_LOC_364/A NOR2X1_LOC_862/B 0.10fF
C11239 INVX1_LOC_101/Y NOR2X1_LOC_89/A 0.02fF
C11240 INVX1_LOC_225/A INVX1_LOC_33/Y 0.00fF
C11241 NOR2X1_LOC_45/B NAND2X1_LOC_632/a_36_24# 0.00fF
C11242 INVX1_LOC_35/A NAND2X1_LOC_175/Y 0.02fF
C11243 NOR2X1_LOC_383/Y NOR2X1_LOC_78/A 0.02fF
C11244 NOR2X1_LOC_361/B NAND2X1_LOC_807/B 0.15fF
C11245 NOR2X1_LOC_431/Y NAND2X1_LOC_434/Y 0.09fF
C11246 NOR2X1_LOC_655/B VDD 2.72fF
C11247 NOR2X1_LOC_596/A INVX1_LOC_307/A 0.03fF
C11248 NAND2X1_LOC_537/Y INVX1_LOC_42/A 0.08fF
C11249 NAND2X1_LOC_361/Y NOR2X1_LOC_489/A 0.01fF
C11250 D_INPUT_1 INVX1_LOC_224/Y 0.75fF
C11251 NAND2X1_LOC_181/Y NOR2X1_LOC_266/B 0.00fF
C11252 NOR2X1_LOC_78/A NOR2X1_LOC_366/Y 0.02fF
C11253 NOR2X1_LOC_208/Y NOR2X1_LOC_155/A 0.28fF
C11254 INVX1_LOC_95/A NAND2X1_LOC_573/A 0.01fF
C11255 NOR2X1_LOC_658/Y INVX1_LOC_186/Y 0.01fF
C11256 INVX1_LOC_223/Y NAND2X1_LOC_72/B 0.01fF
C11257 INVX1_LOC_277/A INVX1_LOC_19/A 0.11fF
C11258 INVX1_LOC_31/A INVX1_LOC_29/A 0.31fF
C11259 INVX1_LOC_85/A INVX1_LOC_9/A 0.03fF
C11260 NOR2X1_LOC_389/A INVX1_LOC_12/A 0.10fF
C11261 NOR2X1_LOC_151/Y INPUT_0 -0.00fF
C11262 NOR2X1_LOC_532/Y INVX1_LOC_91/A 0.05fF
C11263 NOR2X1_LOC_326/Y NOR2X1_LOC_324/A 0.37fF
C11264 INVX1_LOC_268/A INVX1_LOC_46/A 0.02fF
C11265 NAND2X1_LOC_555/Y NOR2X1_LOC_128/A 0.04fF
C11266 NOR2X1_LOC_516/B NOR2X1_LOC_858/B 0.04fF
C11267 INVX1_LOC_157/A NAND2X1_LOC_468/B 0.31fF
C11268 NOR2X1_LOC_482/Y INVX1_LOC_38/A 0.03fF
C11269 NOR2X1_LOC_848/Y INVX1_LOC_15/A 0.03fF
C11270 INVX1_LOC_193/Y NOR2X1_LOC_706/A 0.01fF
C11271 NOR2X1_LOC_573/Y INVX1_LOC_42/A 0.01fF
C11272 INVX1_LOC_10/A NAND2X1_LOC_469/B 0.27fF
C11273 NAND2X1_LOC_199/B INVX1_LOC_12/A 0.03fF
C11274 NOR2X1_LOC_781/A NOR2X1_LOC_586/Y 0.03fF
C11275 INVX1_LOC_17/A INVX1_LOC_4/A 0.10fF
C11276 NAND2X1_LOC_624/A INVX1_LOC_255/A 0.25fF
C11277 INVX1_LOC_177/A INVX1_LOC_54/A 0.03fF
C11278 INVX1_LOC_15/Y NOR2X1_LOC_629/Y 0.01fF
C11279 NAND2X1_LOC_358/Y VDD 0.10fF
C11280 NOR2X1_LOC_775/Y NOR2X1_LOC_78/A 0.02fF
C11281 INVX1_LOC_180/A NAND2X1_LOC_432/a_36_24# 0.01fF
C11282 INVX1_LOC_227/A NOR2X1_LOC_137/Y 0.02fF
C11283 NOR2X1_LOC_778/B NOR2X1_LOC_729/A 0.18fF
C11284 NOR2X1_LOC_309/Y NOR2X1_LOC_155/A 0.01fF
C11285 INVX1_LOC_135/A NOR2X1_LOC_825/Y 0.16fF
C11286 INVX1_LOC_10/A NOR2X1_LOC_447/B 0.01fF
C11287 NOR2X1_LOC_471/Y INVX1_LOC_4/A 0.16fF
C11288 INVX1_LOC_280/Y INVX1_LOC_54/A 0.07fF
C11289 INVX1_LOC_107/A INVX1_LOC_12/A 0.01fF
C11290 NAND2X1_LOC_149/Y NOR2X1_LOC_635/B 0.04fF
C11291 VDD NOR2X1_LOC_99/B 2.17fF
C11292 NOR2X1_LOC_388/Y INVX1_LOC_84/A 0.07fF
C11293 NAND2X1_LOC_555/Y INVX1_LOC_4/A 0.03fF
C11294 INVX1_LOC_290/A INVX1_LOC_38/A 0.08fF
C11295 NAND2X1_LOC_787/A INVX1_LOC_306/Y 0.40fF
C11296 D_GATE_366 INVX1_LOC_76/A 0.03fF
C11297 VDD NOR2X1_LOC_846/B -0.00fF
C11298 NOR2X1_LOC_666/A NOR2X1_LOC_383/B 0.01fF
C11299 NOR2X1_LOC_596/A INVX1_LOC_12/A 0.17fF
C11300 NAND2X1_LOC_363/B INVX1_LOC_306/Y 0.01fF
C11301 D_INPUT_0 INVX1_LOC_117/A 0.52fF
C11302 INVX1_LOC_25/Y NOR2X1_LOC_177/Y 0.09fF
C11303 NOR2X1_LOC_220/A INVX1_LOC_307/A 0.10fF
C11304 NOR2X1_LOC_552/A NOR2X1_LOC_335/B 0.03fF
C11305 INVX1_LOC_314/Y NOR2X1_LOC_327/a_36_216# 0.01fF
C11306 NAND2X1_LOC_364/Y NOR2X1_LOC_777/B 0.46fF
C11307 NOR2X1_LOC_791/A INVX1_LOC_3/Y -0.01fF
C11308 INVX1_LOC_75/A NOR2X1_LOC_631/B 0.07fF
C11309 NOR2X1_LOC_803/A VDD 0.24fF
C11310 NOR2X1_LOC_220/A NOR2X1_LOC_445/B 0.10fF
C11311 NOR2X1_LOC_289/Y INVX1_LOC_76/A 0.03fF
C11312 INVX1_LOC_50/A NAND2X1_LOC_538/Y 0.28fF
C11313 INVX1_LOC_182/A VDD 0.64fF
C11314 INVX1_LOC_33/A INVX1_LOC_109/A 0.05fF
C11315 NAND2X1_LOC_337/B NOR2X1_LOC_831/a_36_216# 0.00fF
C11316 INVX1_LOC_77/A INVX1_LOC_290/Y 0.07fF
C11317 NOR2X1_LOC_439/B INVX1_LOC_37/A 0.01fF
C11318 INVX1_LOC_50/A NOR2X1_LOC_250/A 0.01fF
C11319 NOR2X1_LOC_791/Y INVX1_LOC_306/Y 0.02fF
C11320 INVX1_LOC_186/A NOR2X1_LOC_78/A 0.08fF
C11321 NOR2X1_LOC_160/B NOR2X1_LOC_72/Y 0.03fF
C11322 NOR2X1_LOC_87/B INVX1_LOC_19/A 0.03fF
C11323 INVX1_LOC_28/A NOR2X1_LOC_816/Y 0.07fF
C11324 NAND2X1_LOC_18/a_36_24# D_INPUT_6 0.00fF
C11325 D_INPUT_1 NOR2X1_LOC_103/Y 0.53fF
C11326 INVX1_LOC_75/A INVX1_LOC_37/A 14.95fF
C11327 INVX1_LOC_150/Y INVX1_LOC_270/Y 0.00fF
C11328 NOR2X1_LOC_745/a_36_216# INVX1_LOC_23/A 0.00fF
C11329 INVX1_LOC_279/A INVX1_LOC_92/A 0.08fF
C11330 NOR2X1_LOC_848/Y INVX1_LOC_108/Y 0.00fF
C11331 NOR2X1_LOC_719/A INVX1_LOC_123/Y 0.11fF
C11332 NOR2X1_LOC_548/Y NOR2X1_LOC_445/B 0.15fF
C11333 NOR2X1_LOC_76/A INVX1_LOC_118/A 0.14fF
C11334 INVX1_LOC_170/A INVX1_LOC_23/Y 0.02fF
C11335 NOR2X1_LOC_45/B NOR2X1_LOC_405/A 0.02fF
C11336 INPUT_0 NAND2X1_LOC_633/Y 0.11fF
C11337 INVX1_LOC_21/A INVX1_LOC_222/Y 0.03fF
C11338 INVX1_LOC_22/A NOR2X1_LOC_697/Y 0.00fF
C11339 NOR2X1_LOC_852/A INVX1_LOC_26/Y 0.04fF
C11340 INVX1_LOC_17/A INVX1_LOC_64/A 0.10fF
C11341 INVX1_LOC_43/Y NAND2X1_LOC_203/a_36_24# 0.00fF
C11342 INVX1_LOC_136/A NOR2X1_LOC_282/Y 0.03fF
C11343 INVX1_LOC_225/Y INVX1_LOC_58/Y 0.29fF
C11344 NOR2X1_LOC_78/A NAND2X1_LOC_447/Y 0.01fF
C11345 NOR2X1_LOC_52/B NOR2X1_LOC_114/Y 0.04fF
C11346 INVX1_LOC_135/A NOR2X1_LOC_88/Y 0.10fF
C11347 NOR2X1_LOC_689/Y INVX1_LOC_36/A 0.03fF
C11348 NOR2X1_LOC_415/A NAND2X1_LOC_141/Y 0.03fF
C11349 NOR2X1_LOC_6/B NOR2X1_LOC_554/A 0.06fF
C11350 INVX1_LOC_35/A INPUT_3 0.06fF
C11351 INVX1_LOC_80/A NOR2X1_LOC_649/B 0.08fF
C11352 NAND2X1_LOC_482/a_36_24# NOR2X1_LOC_155/A 0.01fF
C11353 INVX1_LOC_18/A NOR2X1_LOC_727/B 0.03fF
C11354 NOR2X1_LOC_307/A INVX1_LOC_213/A 0.05fF
C11355 INVX1_LOC_45/A D_INPUT_1 0.30fF
C11356 INVX1_LOC_36/A NOR2X1_LOC_125/Y 0.15fF
C11357 INVX1_LOC_2/Y INVX1_LOC_91/A 0.00fF
C11358 NOR2X1_LOC_315/Y INVX1_LOC_19/Y 0.29fF
C11359 INVX1_LOC_35/A NOR2X1_LOC_201/a_36_216# 0.02fF
C11360 NAND2X1_LOC_581/Y NAND2X1_LOC_3/B 0.20fF
C11361 INVX1_LOC_7/Y NOR2X1_LOC_82/A 0.01fF
C11362 INVX1_LOC_174/Y INVX1_LOC_19/A 0.00fF
C11363 INVX1_LOC_199/A INVX1_LOC_115/A 0.01fF
C11364 INVX1_LOC_289/Y NOR2X1_LOC_92/Y 0.10fF
C11365 NOR2X1_LOC_598/B INVX1_LOC_36/A 0.04fF
C11366 INVX1_LOC_135/A INVX1_LOC_84/A 0.31fF
C11367 INVX1_LOC_247/Y INVX1_LOC_23/A 0.04fF
C11368 INVX1_LOC_280/Y NOR2X1_LOC_48/B 0.10fF
C11369 INVX1_LOC_41/A INVX1_LOC_87/A 2.61fF
C11370 INVX1_LOC_182/Y INVX1_LOC_92/A 0.03fF
C11371 NOR2X1_LOC_160/B INVX1_LOC_50/Y 0.10fF
C11372 NOR2X1_LOC_510/Y NAND2X1_LOC_350/A 0.03fF
C11373 INVX1_LOC_291/Y VDD 0.33fF
C11374 INVX1_LOC_88/A NOR2X1_LOC_348/Y 0.07fF
C11375 INVX1_LOC_269/A NOR2X1_LOC_15/Y 0.13fF
C11376 INVX1_LOC_95/Y INVX1_LOC_46/A 0.07fF
C11377 INVX1_LOC_72/A NOR2X1_LOC_678/A 0.07fF
C11378 INVX1_LOC_291/Y NAND2X1_LOC_800/A 0.01fF
C11379 NOR2X1_LOC_226/A NAND2X1_LOC_404/a_36_24# 0.00fF
C11380 INVX1_LOC_224/Y NOR2X1_LOC_403/B 0.00fF
C11381 NOR2X1_LOC_15/Y NOR2X1_LOC_232/Y 0.03fF
C11382 INVX1_LOC_136/A NAND2X1_LOC_549/Y 0.04fF
C11383 INVX1_LOC_18/A NOR2X1_LOC_717/A 0.10fF
C11384 INVX1_LOC_36/A NAND2X1_LOC_725/A 0.01fF
C11385 INVX1_LOC_285/Y INVX1_LOC_54/A 0.09fF
C11386 NOR2X1_LOC_82/A NOR2X1_LOC_92/Y 0.03fF
C11387 INVX1_LOC_201/Y INVX1_LOC_175/A 0.03fF
C11388 INVX1_LOC_33/Y NAND2X1_LOC_642/Y 0.03fF
C11389 INVX1_LOC_12/Y NOR2X1_LOC_124/A 0.08fF
C11390 INVX1_LOC_144/A NOR2X1_LOC_435/A 0.01fF
C11391 NOR2X1_LOC_510/Y NOR2X1_LOC_441/Y 0.13fF
C11392 INVX1_LOC_180/A INVX1_LOC_271/A 0.20fF
C11393 NOR2X1_LOC_606/Y INVX1_LOC_13/Y 0.01fF
C11394 NAND2X1_LOC_326/A INVX1_LOC_161/Y 0.01fF
C11395 NOR2X1_LOC_285/B INVX1_LOC_26/Y 0.00fF
C11396 D_INPUT_1 INVX1_LOC_71/A 0.23fF
C11397 INVX1_LOC_30/A INVX1_LOC_306/Y 0.03fF
C11398 INVX1_LOC_198/Y NOR2X1_LOC_678/A 0.05fF
C11399 NAND2X1_LOC_662/B INVX1_LOC_117/Y 0.01fF
C11400 INVX1_LOC_45/A NOR2X1_LOC_652/Y 0.07fF
C11401 NAND2X1_LOC_573/A NAND2X1_LOC_807/B 0.03fF
C11402 NOR2X1_LOC_91/A INVX1_LOC_8/A 0.19fF
C11403 INVX1_LOC_21/A NAND2X1_LOC_577/A 0.07fF
C11404 INVX1_LOC_256/A INVX1_LOC_88/A 0.06fF
C11405 NAND2X1_LOC_552/A NOR2X1_LOC_68/A 0.00fF
C11406 NAND2X1_LOC_579/A NOR2X1_LOC_369/Y 0.11fF
C11407 INVX1_LOC_5/A NOR2X1_LOC_68/A 0.45fF
C11408 INVX1_LOC_37/A NAND2X1_LOC_453/A 0.00fF
C11409 NOR2X1_LOC_78/B INVX1_LOC_271/Y 0.07fF
C11410 NAND2X1_LOC_479/Y INVX1_LOC_15/A 0.01fF
C11411 INVX1_LOC_230/Y INVX1_LOC_14/A 0.22fF
C11412 NOR2X1_LOC_243/Y NOR2X1_LOC_342/B 0.26fF
C11413 NAND2X1_LOC_310/a_36_24# INVX1_LOC_23/A 0.00fF
C11414 INVX1_LOC_25/A NOR2X1_LOC_772/Y 0.08fF
C11415 NOR2X1_LOC_516/a_36_216# INVX1_LOC_23/A 0.02fF
C11416 VDD NOR2X1_LOC_176/Y 0.01fF
C11417 INVX1_LOC_120/A NOR2X1_LOC_67/Y 0.00fF
C11418 INVX1_LOC_269/A NAND2X1_LOC_321/a_36_24# 0.00fF
C11419 INVX1_LOC_8/A INVX1_LOC_23/A 0.13fF
C11420 NAND2X1_LOC_850/Y NOR2X1_LOC_301/A 0.07fF
C11421 NOR2X1_LOC_76/A NAND2X1_LOC_455/B 0.03fF
C11422 INVX1_LOC_25/A NOR2X1_LOC_392/B 0.03fF
C11423 NOR2X1_LOC_68/A INVX1_LOC_178/A 0.10fF
C11424 NOR2X1_LOC_361/B NOR2X1_LOC_441/Y 0.45fF
C11425 INVX1_LOC_5/A NOR2X1_LOC_204/a_36_216# 0.00fF
C11426 NOR2X1_LOC_554/B NAND2X1_LOC_473/A 0.19fF
C11427 NOR2X1_LOC_825/Y INVX1_LOC_280/A 0.35fF
C11428 INVX1_LOC_144/A INVX1_LOC_63/A 0.01fF
C11429 NOR2X1_LOC_425/Y INVX1_LOC_77/Y 0.01fF
C11430 NOR2X1_LOC_211/A INVX1_LOC_87/A 0.00fF
C11431 NOR2X1_LOC_94/Y NOR2X1_LOC_825/Y 0.19fF
C11432 NOR2X1_LOC_391/B INVX1_LOC_84/A 0.01fF
C11433 INVX1_LOC_71/A NOR2X1_LOC_652/Y 0.11fF
C11434 NOR2X1_LOC_730/Y INVX1_LOC_274/Y 0.88fF
C11435 D_INPUT_0 INVX1_LOC_3/Y 0.20fF
C11436 NOR2X1_LOC_589/A INVX1_LOC_94/Y 0.39fF
C11437 INVX1_LOC_135/A INVX1_LOC_15/A 0.14fF
C11438 INVX1_LOC_133/Y INVX1_LOC_271/A 0.00fF
C11439 INVX1_LOC_125/Y NAND2X1_LOC_572/B 0.03fF
C11440 INVX1_LOC_35/A INVX1_LOC_158/A 0.03fF
C11441 NOR2X1_LOC_560/A INVX1_LOC_15/A 0.28fF
C11442 NOR2X1_LOC_454/Y INVX1_LOC_77/A 1.48fF
C11443 NOR2X1_LOC_845/A INVX1_LOC_63/A 0.12fF
C11444 NOR2X1_LOC_837/A INVX1_LOC_19/A 0.01fF
C11445 NOR2X1_LOC_589/A INVX1_LOC_181/A 0.01fF
C11446 INVX1_LOC_6/A INVX1_LOC_29/A 1.02fF
C11447 NOR2X1_LOC_857/A NOR2X1_LOC_862/B 0.10fF
C11448 INVX1_LOC_286/A NAND2X1_LOC_81/B 0.07fF
C11449 INVX1_LOC_151/Y INVX1_LOC_23/A 0.01fF
C11450 INVX1_LOC_58/A NAND2X1_LOC_752/a_36_24# 0.00fF
C11451 NOR2X1_LOC_68/A NOR2X1_LOC_816/A 0.06fF
C11452 NAND2X1_LOC_537/Y NOR2X1_LOC_152/Y 0.17fF
C11453 NAND2X1_LOC_538/Y NOR2X1_LOC_152/a_36_216# 0.00fF
C11454 INVX1_LOC_76/A INVX1_LOC_123/Y 0.07fF
C11455 NAND2X1_LOC_860/A NAND2X1_LOC_860/Y 0.03fF
C11456 INVX1_LOC_48/Y INVX1_LOC_33/A 0.08fF
C11457 INVX1_LOC_102/A NOR2X1_LOC_167/Y 0.05fF
C11458 NOR2X1_LOC_561/Y INVX1_LOC_296/Y 3.83fF
C11459 NOR2X1_LOC_657/Y INVX1_LOC_30/A 0.02fF
C11460 INVX1_LOC_58/A NAND2X1_LOC_660/Y 0.03fF
C11461 INVX1_LOC_223/A NOR2X1_LOC_565/A 0.00fF
C11462 INVX1_LOC_1/A NOR2X1_LOC_772/Y 0.11fF
C11463 NAND2X1_LOC_736/Y NAND2X1_LOC_559/Y 0.06fF
C11464 NOR2X1_LOC_67/A NAND2X1_LOC_214/B 0.00fF
C11465 INVX1_LOC_141/A NOR2X1_LOC_512/Y 0.12fF
C11466 INVX1_LOC_46/Y INVX1_LOC_117/A 0.32fF
C11467 INVX1_LOC_1/A NOR2X1_LOC_147/B 0.07fF
C11468 INVX1_LOC_122/Y INVX1_LOC_210/Y 0.03fF
C11469 INVX1_LOC_256/A INVX1_LOC_303/A 0.04fF
C11470 NOR2X1_LOC_798/A INVX1_LOC_196/A 0.03fF
C11471 INVX1_LOC_35/A NAND2X1_LOC_564/B 0.06fF
C11472 INVX1_LOC_1/A NOR2X1_LOC_392/B 0.10fF
C11473 NOR2X1_LOC_294/Y INVX1_LOC_205/A 0.00fF
C11474 NOR2X1_LOC_813/Y NOR2X1_LOC_88/Y 0.03fF
C11475 INVX1_LOC_267/A INVX1_LOC_235/Y 0.03fF
C11476 NOR2X1_LOC_389/B INVX1_LOC_116/Y 0.00fF
C11477 NOR2X1_LOC_139/Y NOR2X1_LOC_89/A 0.03fF
C11478 INVX1_LOC_228/A INVX1_LOC_31/A 0.04fF
C11479 INVX1_LOC_50/A NOR2X1_LOC_106/A 0.36fF
C11480 INVX1_LOC_95/A NAND2X1_LOC_81/B 0.05fF
C11481 NAND2X1_LOC_850/A NOR2X1_LOC_278/Y 0.06fF
C11482 INVX1_LOC_279/A INVX1_LOC_53/A 0.54fF
C11483 INVX1_LOC_35/A GATE_662 0.22fF
C11484 NOR2X1_LOC_533/Y NAND2X1_LOC_354/B 0.00fF
C11485 NAND2X1_LOC_807/Y NOR2X1_LOC_281/Y 0.01fF
C11486 INVX1_LOC_139/Y INVX1_LOC_84/A 0.03fF
C11487 INVX1_LOC_58/A D_INPUT_0 0.93fF
C11488 NOR2X1_LOC_67/A INVX1_LOC_27/A 0.12fF
C11489 INVX1_LOC_41/A NOR2X1_LOC_82/A 0.14fF
C11490 NAND2X1_LOC_53/Y INVX1_LOC_63/Y 0.10fF
C11491 INVX1_LOC_75/A NAND2X1_LOC_72/B 0.01fF
C11492 NAND2X1_LOC_140/A INVX1_LOC_23/A 0.03fF
C11493 D_INPUT_1 NOR2X1_LOC_123/B 0.07fF
C11494 INVX1_LOC_201/Y NOR2X1_LOC_82/A 0.09fF
C11495 NOR2X1_LOC_287/A NOR2X1_LOC_798/A 0.00fF
C11496 NOR2X1_LOC_516/B INVX1_LOC_50/Y 0.03fF
C11497 INVX1_LOC_45/A NOR2X1_LOC_403/B 0.05fF
C11498 NAND2X1_LOC_559/Y INVX1_LOC_282/Y 0.13fF
C11499 INVX1_LOC_269/A NAND2X1_LOC_141/A 0.01fF
C11500 NOR2X1_LOC_798/A NOR2X1_LOC_748/a_36_216# 0.00fF
C11501 NOR2X1_LOC_772/B NOR2X1_LOC_440/Y 0.13fF
C11502 INVX1_LOC_174/A NAND2X1_LOC_157/a_36_24# 0.01fF
C11503 NAND2X1_LOC_740/a_36_24# NAND2X1_LOC_811/Y 0.01fF
C11504 NAND2X1_LOC_860/A NAND2X1_LOC_861/Y 0.13fF
C11505 NOR2X1_LOC_32/B NOR2X1_LOC_130/A 0.02fF
C11506 NAND2X1_LOC_468/B NOR2X1_LOC_89/A 0.00fF
C11507 NOR2X1_LOC_813/Y INVX1_LOC_84/A 0.05fF
C11508 INVX1_LOC_278/A INVX1_LOC_135/A 0.10fF
C11509 INVX1_LOC_269/A INVX1_LOC_15/Y 0.58fF
C11510 INVX1_LOC_12/A NAND2X1_LOC_469/B 0.03fF
C11511 INVX1_LOC_25/A INVX1_LOC_90/A 0.10fF
C11512 INVX1_LOC_230/Y INVX1_LOC_217/Y 0.00fF
C11513 NOR2X1_LOC_453/Y NOR2X1_LOC_222/Y 0.38fF
C11514 INVX1_LOC_286/A INVX1_LOC_4/Y 0.07fF
C11515 INVX1_LOC_10/Y INVX1_LOC_84/A 0.07fF
C11516 INVX1_LOC_31/A NOR2X1_LOC_516/a_36_216# 0.01fF
C11517 INVX1_LOC_25/A NOR2X1_LOC_389/B 0.89fF
C11518 INVX1_LOC_48/Y INVX1_LOC_40/A 0.07fF
C11519 NOR2X1_LOC_479/B INVX1_LOC_239/A 0.09fF
C11520 NOR2X1_LOC_440/Y INVX1_LOC_13/Y 0.46fF
C11521 NOR2X1_LOC_759/A NOR2X1_LOC_759/Y 0.02fF
C11522 NOR2X1_LOC_160/B NOR2X1_LOC_6/B 0.19fF
C11523 INVX1_LOC_31/A INVX1_LOC_8/A 0.07fF
C11524 INVX1_LOC_84/A INVX1_LOC_280/A 0.33fF
C11525 NOR2X1_LOC_75/Y INVX1_LOC_266/Y 0.36fF
C11526 INVX1_LOC_292/A INVX1_LOC_104/A 0.65fF
C11527 NOR2X1_LOC_94/Y INVX1_LOC_84/A 0.03fF
C11528 NOR2X1_LOC_155/A NOR2X1_LOC_435/A 0.02fF
C11529 INVX1_LOC_50/A NAND2X1_LOC_863/A 0.07fF
C11530 INVX1_LOC_298/Y INVX1_LOC_6/A 0.03fF
C11531 INVX1_LOC_17/A NAND2X1_LOC_850/Y 0.07fF
C11532 NOR2X1_LOC_447/B INVX1_LOC_12/A 0.02fF
C11533 INVX1_LOC_37/A NAND2X1_LOC_291/B 0.00fF
C11534 INVX1_LOC_181/Y INVX1_LOC_314/Y 0.01fF
C11535 NOR2X1_LOC_223/B INVX1_LOC_295/A 0.02fF
C11536 NAND2X1_LOC_542/a_36_24# NOR2X1_LOC_246/A 0.00fF
C11537 NOR2X1_LOC_357/Y NOR2X1_LOC_631/a_36_216# 0.00fF
C11538 NAND2X1_LOC_806/a_36_24# INVX1_LOC_46/A 0.00fF
C11539 INVX1_LOC_294/Y INVX1_LOC_30/A 0.04fF
C11540 NOR2X1_LOC_527/a_36_216# INVX1_LOC_57/A 0.00fF
C11541 NOR2X1_LOC_716/B NOR2X1_LOC_91/a_36_216# 0.01fF
C11542 NAND2X1_LOC_254/Y NAND2X1_LOC_254/a_36_24# 0.02fF
C11543 NOR2X1_LOC_381/Y NOR2X1_LOC_516/B 0.09fF
C11544 INVX1_LOC_177/Y INVX1_LOC_67/A 0.11fF
C11545 NOR2X1_LOC_123/B NOR2X1_LOC_652/Y 0.00fF
C11546 INVX1_LOC_25/A NAND2X1_LOC_348/A 0.10fF
C11547 INVX1_LOC_182/Y INVX1_LOC_53/A -0.04fF
C11548 VDD NOR2X1_LOC_850/B 0.28fF
C11549 NAND2X1_LOC_352/B NAND2X1_LOC_342/Y 0.38fF
C11550 INVX1_LOC_36/A NAND2X1_LOC_308/Y 0.01fF
C11551 NOR2X1_LOC_99/Y INVX1_LOC_3/A 0.05fF
C11552 NOR2X1_LOC_294/a_36_216# NOR2X1_LOC_87/B 0.00fF
C11553 INVX1_LOC_246/A NAND2X1_LOC_798/A 0.22fF
C11554 NOR2X1_LOC_321/Y NAND2X1_LOC_656/Y 0.11fF
C11555 INVX1_LOC_109/Y INVX1_LOC_281/A 0.01fF
C11556 NOR2X1_LOC_798/A INVX1_LOC_47/A 0.03fF
C11557 INVX1_LOC_38/A INVX1_LOC_261/Y 0.04fF
C11558 NOR2X1_LOC_68/A NOR2X1_LOC_377/Y 0.03fF
C11559 NOR2X1_LOC_553/Y NOR2X1_LOC_541/Y 0.00fF
C11560 NOR2X1_LOC_831/B INVX1_LOC_285/A 0.01fF
C11561 INVX1_LOC_235/Y INVX1_LOC_89/A 0.06fF
C11562 NAND2X1_LOC_149/Y INVX1_LOC_89/A 0.12fF
C11563 NAND2X1_LOC_776/a_36_24# NAND2X1_LOC_722/A 0.00fF
C11564 NOR2X1_LOC_155/A INVX1_LOC_63/A 0.01fF
C11565 NOR2X1_LOC_831/B NOR2X1_LOC_814/A 0.31fF
C11566 NOR2X1_LOC_351/Y INVX1_LOC_109/A 0.04fF
C11567 NOR2X1_LOC_290/Y NAND2X1_LOC_634/Y 0.15fF
C11568 INVX1_LOC_94/Y INVX1_LOC_20/A 0.07fF
C11569 NOR2X1_LOC_720/B INVX1_LOC_24/A 0.00fF
C11570 INVX1_LOC_64/A NOR2X1_LOC_594/Y 0.03fF
C11571 NOR2X1_LOC_550/a_36_216# NOR2X1_LOC_500/Y 0.01fF
C11572 INVX1_LOC_215/Y NAND2X1_LOC_660/Y 0.07fF
C11573 NOR2X1_LOC_415/a_36_216# INVX1_LOC_14/A 0.01fF
C11574 INVX1_LOC_21/A NOR2X1_LOC_329/B 0.33fF
C11575 INVX1_LOC_299/A INVX1_LOC_171/A 0.01fF
C11576 INVX1_LOC_30/Y NOR2X1_LOC_160/B 0.05fF
C11577 NOR2X1_LOC_813/Y INVX1_LOC_15/A 0.07fF
C11578 NAND2X1_LOC_711/Y INVX1_LOC_16/A 0.03fF
C11579 NAND2X1_LOC_741/B NAND2X1_LOC_852/Y 0.05fF
C11580 NOR2X1_LOC_264/Y NAND2X1_LOC_7/Y 0.03fF
C11581 INVX1_LOC_290/Y INVX1_LOC_9/A 0.00fF
C11582 INVX1_LOC_271/Y INVX1_LOC_46/A 0.07fF
C11583 INVX1_LOC_91/A INVX1_LOC_29/Y 0.07fF
C11584 INVX1_LOC_90/A INVX1_LOC_1/A 4.91fF
C11585 NAND2X1_LOC_848/A INVX1_LOC_3/Y 0.01fF
C11586 INVX1_LOC_10/Y INVX1_LOC_15/A 0.04fF
C11587 INPUT_2 INVX1_LOC_7/A 0.08fF
C11588 INVX1_LOC_21/A D_INPUT_4 0.01fF
C11589 NOR2X1_LOC_426/Y INVX1_LOC_22/A 0.03fF
C11590 INPUT_4 INVX1_LOC_173/A 0.03fF
C11591 NOR2X1_LOC_389/B INVX1_LOC_1/A 1.55fF
C11592 INVX1_LOC_24/A NOR2X1_LOC_822/Y 0.02fF
C11593 INVX1_LOC_38/A NOR2X1_LOC_467/A 0.07fF
C11594 INVX1_LOC_280/A INVX1_LOC_15/A 0.22fF
C11595 NOR2X1_LOC_68/A NOR2X1_LOC_773/Y 0.01fF
C11596 NOR2X1_LOC_94/Y INVX1_LOC_15/A 0.03fF
C11597 NOR2X1_LOC_142/Y INVX1_LOC_153/Y 0.10fF
C11598 INVX1_LOC_124/A INVX1_LOC_77/A 0.17fF
C11599 NOR2X1_LOC_596/A NAND2X1_LOC_832/a_36_24# 0.00fF
C11600 INVX1_LOC_20/A INVX1_LOC_181/A 0.03fF
C11601 NAND2X1_LOC_341/a_36_24# INVX1_LOC_159/A 0.00fF
C11602 INVX1_LOC_67/A INVX1_LOC_104/A 0.23fF
C11603 NAND2X1_LOC_161/a_36_24# NAND2X1_LOC_451/Y 0.01fF
C11604 NOR2X1_LOC_794/B INVX1_LOC_97/A 0.01fF
C11605 NAND2X1_LOC_733/Y NAND2X1_LOC_795/Y 0.03fF
C11606 NOR2X1_LOC_368/A NAND2X1_LOC_75/a_36_24# 0.00fF
C11607 NOR2X1_LOC_457/A NOR2X1_LOC_356/A 0.07fF
C11608 NOR2X1_LOC_35/Y NOR2X1_LOC_748/A 0.05fF
C11609 INVX1_LOC_223/A NOR2X1_LOC_561/Y 0.10fF
C11610 INVX1_LOC_90/A NOR2X1_LOC_794/B 0.10fF
C11611 NAND2X1_LOC_9/Y INVX1_LOC_95/Y 0.04fF
C11612 NAND2X1_LOC_348/A INVX1_LOC_1/A 0.03fF
C11613 NOR2X1_LOC_454/Y NAND2X1_LOC_832/Y 0.02fF
C11614 NAND2X1_LOC_349/B NAND2X1_LOC_198/B 0.20fF
C11615 NOR2X1_LOC_246/Y NAND2X1_LOC_352/B 0.00fF
C11616 NOR2X1_LOC_142/Y INVX1_LOC_177/A 0.05fF
C11617 INVX1_LOC_233/A INVX1_LOC_95/Y 0.07fF
C11618 INVX1_LOC_238/A NAND2X1_LOC_866/B 0.13fF
C11619 INVX1_LOC_94/A INVX1_LOC_1/Y 0.18fF
C11620 NOR2X1_LOC_553/Y INVX1_LOC_71/A 0.03fF
C11621 INVX1_LOC_35/A NOR2X1_LOC_332/B 0.01fF
C11622 NOR2X1_LOC_655/B INVX1_LOC_153/Y 0.10fF
C11623 INVX1_LOC_85/A NAND2X1_LOC_629/Y 0.00fF
C11624 INVX1_LOC_217/A NAND2X1_LOC_795/Y 0.12fF
C11625 INVX1_LOC_40/A NOR2X1_LOC_6/a_36_216# 0.00fF
C11626 NOR2X1_LOC_218/A NOR2X1_LOC_216/Y 0.01fF
C11627 INVX1_LOC_299/A INVX1_LOC_222/A 0.85fF
C11628 INVX1_LOC_14/A NOR2X1_LOC_292/Y 0.03fF
C11629 INVX1_LOC_132/A INVX1_LOC_232/A 0.10fF
C11630 NAND2X1_LOC_711/Y INVX1_LOC_28/A 0.00fF
C11631 NOR2X1_LOC_657/a_36_216# NOR2X1_LOC_78/A 0.00fF
C11632 VDD INVX1_LOC_308/A 0.12fF
C11633 NAND2X1_LOC_553/A INVX1_LOC_95/Y 0.20fF
C11634 NOR2X1_LOC_457/A NOR2X1_LOC_74/A 0.10fF
C11635 INVX1_LOC_78/A NOR2X1_LOC_487/Y 0.01fF
C11636 NOR2X1_LOC_423/a_36_216# NOR2X1_LOC_357/Y 0.00fF
C11637 INVX1_LOC_30/A NOR2X1_LOC_356/A 0.10fF
C11638 INVX1_LOC_90/A NOR2X1_LOC_384/Y 0.12fF
C11639 INVX1_LOC_33/A NOR2X1_LOC_374/B 0.07fF
C11640 NOR2X1_LOC_790/a_36_216# INVX1_LOC_186/A 0.02fF
C11641 NOR2X1_LOC_798/A INVX1_LOC_95/Y 0.06fF
C11642 INVX1_LOC_29/A NOR2X1_LOC_633/A 0.02fF
C11643 INVX1_LOC_224/Y NOR2X1_LOC_99/a_36_216# 0.01fF
C11644 INVX1_LOC_290/A INVX1_LOC_33/A 0.18fF
C11645 NOR2X1_LOC_655/B INVX1_LOC_177/A 0.02fF
C11646 NOR2X1_LOC_453/a_36_216# INVX1_LOC_91/A 0.00fF
C11647 NOR2X1_LOC_431/Y NOR2X1_LOC_130/A 0.01fF
C11648 INVX1_LOC_58/A NAND2X1_LOC_848/A 0.33fF
C11649 INVX1_LOC_15/Y NOR2X1_LOC_616/Y 0.09fF
C11650 NOR2X1_LOC_432/a_36_216# NOR2X1_LOC_78/B 0.00fF
C11651 NAND2X1_LOC_807/B NAND2X1_LOC_81/B 0.19fF
C11652 NAND2X1_LOC_500/B NAND2X1_LOC_254/Y 0.01fF
C11653 INVX1_LOC_209/Y NAND2X1_LOC_319/A 0.43fF
C11654 INVX1_LOC_225/A INVX1_LOC_232/A 0.15fF
C11655 NOR2X1_LOC_516/B NOR2X1_LOC_6/B 0.02fF
C11656 INVX1_LOC_36/A NAND2X1_LOC_560/A 0.03fF
C11657 INVX1_LOC_107/Y NAND2X1_LOC_470/B 0.02fF
C11658 NAND2X1_LOC_563/A NAND2X1_LOC_141/A 0.01fF
C11659 NOR2X1_LOC_409/B NAND2X1_LOC_809/a_36_24# 0.00fF
C11660 D_INPUT_1 NOR2X1_LOC_331/B 0.09fF
C11661 NAND2X1_LOC_354/Y NOR2X1_LOC_329/B 0.03fF
C11662 NAND2X1_LOC_795/Y NAND2X1_LOC_787/B 0.31fF
C11663 NOR2X1_LOC_596/A NOR2X1_LOC_155/a_36_216# 0.02fF
C11664 NOR2X1_LOC_636/A NOR2X1_LOC_763/Y 0.02fF
C11665 INVX1_LOC_118/Y INVX1_LOC_23/A 0.00fF
C11666 INVX1_LOC_289/Y NAND2X1_LOC_648/a_36_24# 0.01fF
C11667 INVX1_LOC_165/Y NOR2X1_LOC_84/Y 0.06fF
C11668 INVX1_LOC_22/A NAND2X1_LOC_453/a_36_24# 0.01fF
C11669 INVX1_LOC_34/A NOR2X1_LOC_391/A 0.00fF
C11670 INVX1_LOC_63/Y INVX1_LOC_10/A 0.17fF
C11671 NOR2X1_LOC_226/A NAND2X1_LOC_181/Y 0.00fF
C11672 NOR2X1_LOC_68/A INVX1_LOC_140/A 0.03fF
C11673 NOR2X1_LOC_742/A NOR2X1_LOC_723/a_36_216# 0.01fF
C11674 NOR2X1_LOC_637/a_36_216# NOR2X1_LOC_130/A 0.00fF
C11675 NOR2X1_LOC_473/B NOR2X1_LOC_106/Y 0.02fF
C11676 INVX1_LOC_292/A INVX1_LOC_206/Y 0.02fF
C11677 INVX1_LOC_30/A NOR2X1_LOC_74/A 0.43fF
C11678 NOR2X1_LOC_808/A NOR2X1_LOC_325/A 0.00fF
C11679 NAND2X1_LOC_659/A NOR2X1_LOC_415/Y 0.02fF
C11680 INVX1_LOC_232/Y INVX1_LOC_316/Y 0.00fF
C11681 NOR2X1_LOC_222/Y NOR2X1_LOC_223/a_36_216# 0.00fF
C11682 NAND2X1_LOC_703/Y NOR2X1_LOC_305/Y 0.01fF
C11683 NOR2X1_LOC_843/B NAND2X1_LOC_85/Y 0.03fF
C11684 NAND2X1_LOC_739/B NAND2X1_LOC_740/B 0.04fF
C11685 NAND2X1_LOC_601/a_36_24# INVX1_LOC_90/A 0.01fF
C11686 INVX1_LOC_30/A NOR2X1_LOC_9/Y 0.73fF
C11687 INVX1_LOC_69/Y NOR2X1_LOC_500/B 0.35fF
C11688 NOR2X1_LOC_612/a_36_216# INVX1_LOC_22/A 0.00fF
C11689 INVX1_LOC_304/Y NAND2X1_LOC_795/Y 0.17fF
C11690 INVX1_LOC_11/A NAND2X1_LOC_468/B 0.03fF
C11691 INVX1_LOC_36/A INVX1_LOC_201/A 0.01fF
C11692 NOR2X1_LOC_703/B NOR2X1_LOC_552/Y 0.00fF
C11693 NAND2X1_LOC_579/A VDD 1.52fF
C11694 NAND2X1_LOC_773/Y INVX1_LOC_46/A 0.13fF
C11695 INVX1_LOC_233/Y INVX1_LOC_54/A 0.02fF
C11696 NAND2X1_LOC_634/Y INVX1_LOC_6/A 0.03fF
C11697 NOR2X1_LOC_383/B NOR2X1_LOC_800/a_36_216# 0.00fF
C11698 NOR2X1_LOC_717/B INVX1_LOC_266/Y 0.01fF
C11699 INVX1_LOC_289/A INVX1_LOC_22/A 0.00fF
C11700 NOR2X1_LOC_187/Y VDD 0.12fF
C11701 NAND2X1_LOC_516/a_36_24# NOR2X1_LOC_45/B 0.01fF
C11702 INVX1_LOC_62/A NOR2X1_LOC_87/B 0.02fF
C11703 INVX1_LOC_53/Y INVX1_LOC_25/Y 0.02fF
C11704 NOR2X1_LOC_78/B INVX1_LOC_279/A 0.18fF
C11705 INVX1_LOC_269/A NOR2X1_LOC_27/a_36_216# 0.00fF
C11706 NOR2X1_LOC_411/Y NOR2X1_LOC_629/Y 0.00fF
C11707 NOR2X1_LOC_422/a_36_216# NOR2X1_LOC_561/Y 0.01fF
C11708 NAND2X1_LOC_349/B INVX1_LOC_53/Y 0.00fF
C11709 NOR2X1_LOC_15/Y INVX1_LOC_12/Y 0.62fF
C11710 INVX1_LOC_209/Y NOR2X1_LOC_409/Y 0.29fF
C11711 INVX1_LOC_55/Y INVX1_LOC_249/Y 0.02fF
C11712 INVX1_LOC_69/Y NOR2X1_LOC_170/a_36_216# 0.01fF
C11713 NAND2X1_LOC_35/Y NOR2X1_LOC_823/a_36_216# 0.01fF
C11714 NOR2X1_LOC_214/B INVX1_LOC_96/Y 0.11fF
C11715 NOR2X1_LOC_596/A NAND2X1_LOC_841/a_36_24# 0.00fF
C11716 INVX1_LOC_77/A NAND2X1_LOC_832/Y 0.01fF
C11717 NAND2X1_LOC_363/B NOR2X1_LOC_865/Y 0.03fF
C11718 INVX1_LOC_119/A INVX1_LOC_28/A 0.34fF
C11719 NAND2X1_LOC_454/Y INVX1_LOC_42/A 0.01fF
C11720 NOR2X1_LOC_307/Y NOR2X1_LOC_833/B 0.31fF
C11721 INVX1_LOC_1/A INVX1_LOC_38/A 1.25fF
C11722 NOR2X1_LOC_420/Y INVX1_LOC_92/A 0.01fF
C11723 INVX1_LOC_145/Y NAND2X1_LOC_349/B 0.23fF
C11724 INVX1_LOC_28/Y INVX1_LOC_29/A 0.02fF
C11725 NOR2X1_LOC_307/B INVX1_LOC_85/Y 0.01fF
C11726 NOR2X1_LOC_318/B INVX1_LOC_94/A 0.08fF
C11727 NOR2X1_LOC_552/A NOR2X1_LOC_168/Y 0.01fF
C11728 NAND2X1_LOC_181/Y INPUT_1 0.00fF
C11729 NOR2X1_LOC_598/B INVX1_LOC_63/A 0.23fF
C11730 NAND2X1_LOC_46/a_36_24# NOR2X1_LOC_814/A 0.00fF
C11731 NOR2X1_LOC_614/Y NOR2X1_LOC_542/Y 0.17fF
C11732 INVX1_LOC_270/A INVX1_LOC_29/A 0.64fF
C11733 NOR2X1_LOC_419/Y INVX1_LOC_125/Y 0.10fF
C11734 INVX1_LOC_214/A NOR2X1_LOC_329/B 0.03fF
C11735 NOR2X1_LOC_142/Y INVX1_LOC_285/Y 0.07fF
C11736 NOR2X1_LOC_151/Y INVX1_LOC_266/Y 0.05fF
C11737 INVX1_LOC_89/A INVX1_LOC_16/A 2.14fF
C11738 NOR2X1_LOC_667/A NOR2X1_LOC_329/B 0.22fF
C11739 NOR2X1_LOC_67/A NOR2X1_LOC_19/B 0.01fF
C11740 INVX1_LOC_150/Y NOR2X1_LOC_536/A 0.12fF
C11741 INVX1_LOC_248/A NOR2X1_LOC_329/B 0.03fF
C11742 INVX1_LOC_215/Y NAND2X1_LOC_848/A 0.01fF
C11743 NOR2X1_LOC_716/B INVX1_LOC_125/Y 0.04fF
C11744 NOR2X1_LOC_78/B INVX1_LOC_182/Y 0.01fF
C11745 NOR2X1_LOC_433/A NOR2X1_LOC_139/Y 0.16fF
C11746 NOR2X1_LOC_770/Y INVX1_LOC_22/A 0.05fF
C11747 INVX1_LOC_19/A INVX1_LOC_58/Y 0.11fF
C11748 NOR2X1_LOC_794/B INVX1_LOC_38/A 0.03fF
C11749 NOR2X1_LOC_433/A NAND2X1_LOC_655/A 0.08fF
C11750 NAND2X1_LOC_722/A NOR2X1_LOC_74/A 0.02fF
C11751 NOR2X1_LOC_292/Y NOR2X1_LOC_612/B 0.04fF
C11752 NAND2X1_LOC_537/Y INVX1_LOC_291/A 0.43fF
C11753 INVX1_LOC_311/A NOR2X1_LOC_423/Y 0.02fF
C11754 INVX1_LOC_33/A INVX1_LOC_160/A 0.01fF
C11755 INVX1_LOC_177/Y NOR2X1_LOC_137/Y 0.02fF
C11756 INVX1_LOC_174/A NAND2X1_LOC_427/a_36_24# 0.00fF
C11757 NAND2X1_LOC_190/Y INVX1_LOC_92/A 0.09fF
C11758 NAND2X1_LOC_425/Y INVX1_LOC_198/A 0.02fF
C11759 INVX1_LOC_78/A NAND2X1_LOC_454/Y 0.07fF
C11760 NOR2X1_LOC_273/Y NOR2X1_LOC_357/Y 0.14fF
C11761 NAND2X1_LOC_326/A NOR2X1_LOC_841/A 0.38fF
C11762 NOR2X1_LOC_457/B INVX1_LOC_14/Y 0.10fF
C11763 NOR2X1_LOC_6/B INVX1_LOC_315/Y 0.02fF
C11764 NOR2X1_LOC_433/A NAND2X1_LOC_468/B 0.02fF
C11765 NOR2X1_LOC_219/Y INVX1_LOC_75/A 0.10fF
C11766 NOR2X1_LOC_759/Y NOR2X1_LOC_357/Y 0.05fF
C11767 INVX1_LOC_132/A NAND2X1_LOC_447/Y 0.00fF
C11768 NOR2X1_LOC_109/Y INVX1_LOC_29/A 0.02fF
C11769 INVX1_LOC_75/A INVX1_LOC_53/Y 0.03fF
C11770 NOR2X1_LOC_222/Y INVX1_LOC_311/A 0.03fF
C11771 INVX1_LOC_60/Y INVX1_LOC_91/A 0.46fF
C11772 INVX1_LOC_83/A NAND2X1_LOC_815/a_36_24# 0.01fF
C11773 INVX1_LOC_26/A INVX1_LOC_165/A 0.01fF
C11774 NOR2X1_LOC_45/a_36_216# NOR2X1_LOC_158/Y 0.01fF
C11775 INVX1_LOC_116/Y NAND2X1_LOC_223/A 0.09fF
C11776 NOR2X1_LOC_384/Y NAND2X1_LOC_849/B 0.08fF
C11777 NOR2X1_LOC_52/B NAND2X1_LOC_655/A 0.77fF
C11778 NOR2X1_LOC_772/B NOR2X1_LOC_89/A 0.08fF
C11779 NOR2X1_LOC_142/Y NOR2X1_LOC_137/B 0.01fF
C11780 INVX1_LOC_28/A INVX1_LOC_150/A 0.04fF
C11781 NOR2X1_LOC_384/Y INVX1_LOC_38/A 0.08fF
C11782 NOR2X1_LOC_209/Y INVX1_LOC_186/A 0.00fF
C11783 NOR2X1_LOC_456/Y INVX1_LOC_32/A 1.27fF
C11784 INVX1_LOC_151/A NAND2X1_LOC_468/B 0.00fF
C11785 NOR2X1_LOC_389/A INVX1_LOC_92/A 0.01fF
C11786 NOR2X1_LOC_577/Y NOR2X1_LOC_681/Y 0.05fF
C11787 INVX1_LOC_50/A NOR2X1_LOC_334/Y 0.15fF
C11788 INVX1_LOC_225/A NAND2X1_LOC_447/Y 0.23fF
C11789 INVX1_LOC_4/Y NAND2X1_LOC_215/A 0.10fF
C11790 NOR2X1_LOC_577/Y INVX1_LOC_37/A 0.07fF
C11791 INVX1_LOC_41/A INVX1_LOC_176/A 0.00fF
C11792 NOR2X1_LOC_82/A NAND2X1_LOC_574/A 0.04fF
C11793 INVX1_LOC_13/Y NOR2X1_LOC_89/A 0.72fF
C11794 NOR2X1_LOC_52/B NAND2X1_LOC_468/B 0.04fF
C11795 INVX1_LOC_132/Y INVX1_LOC_148/A 0.27fF
C11796 NAND2X1_LOC_276/Y INVX1_LOC_2/Y 0.06fF
C11797 NOR2X1_LOC_551/B VDD 0.70fF
C11798 NOR2X1_LOC_590/A NOR2X1_LOC_831/B 0.01fF
C11799 NOR2X1_LOC_391/A INPUT_0 0.00fF
C11800 NOR2X1_LOC_837/B NAND2X1_LOC_825/a_36_24# 0.02fF
C11801 NOR2X1_LOC_799/B NOR2X1_LOC_175/A 0.03fF
C11802 INVX1_LOC_49/A INVX1_LOC_117/A 0.24fF
C11803 NOR2X1_LOC_144/Y INVX1_LOC_46/A 0.05fF
C11804 INVX1_LOC_85/A INVX1_LOC_76/A 0.16fF
C11805 NOR2X1_LOC_315/Y INVX1_LOC_20/A 0.07fF
C11806 INVX1_LOC_59/A NOR2X1_LOC_671/Y 0.04fF
C11807 INVX1_LOC_57/A NOR2X1_LOC_278/Y 1.48fF
C11808 NAND2X1_LOC_352/B INVX1_LOC_285/A 0.00fF
C11809 INVX1_LOC_213/Y VDD 0.24fF
C11810 INVX1_LOC_104/A NOR2X1_LOC_137/Y 0.03fF
C11811 INVX1_LOC_18/A NOR2X1_LOC_640/Y 0.06fF
C11812 NOR2X1_LOC_348/B INVX1_LOC_37/A 0.05fF
C11813 NAND2X1_LOC_239/a_36_24# NAND2X1_LOC_453/A 0.00fF
C11814 INVX1_LOC_77/A INVX1_LOC_9/A 0.18fF
C11815 INVX1_LOC_216/Y NAND2X1_LOC_82/Y 0.01fF
C11816 INVX1_LOC_57/A NOR2X1_LOC_638/Y 0.03fF
C11817 NAND2X1_LOC_72/Y NOR2X1_LOC_334/Y 0.00fF
C11818 INVX1_LOC_64/A INVX1_LOC_94/Y 0.03fF
C11819 INVX1_LOC_232/A NAND2X1_LOC_642/Y 0.10fF
C11820 INVX1_LOC_101/A INVX1_LOC_91/A 0.01fF
C11821 INVX1_LOC_269/A INVX1_LOC_99/A 0.01fF
C11822 NOR2X1_LOC_329/B NAND2X1_LOC_327/a_36_24# 0.01fF
C11823 NAND2X1_LOC_140/A INVX1_LOC_6/A 0.02fF
C11824 INVX1_LOC_88/A NOR2X1_LOC_89/A 0.09fF
C11825 NOR2X1_LOC_396/Y INVX1_LOC_22/A -0.01fF
C11826 NOR2X1_LOC_45/B NOR2X1_LOC_32/Y 0.00fF
C11827 INVX1_LOC_90/A NOR2X1_LOC_188/A 6.93fF
C11828 INVX1_LOC_256/A INVX1_LOC_272/A 0.10fF
C11829 NAND2X1_LOC_369/a_36_24# INVX1_LOC_75/A 0.00fF
C11830 NOR2X1_LOC_596/A INVX1_LOC_92/A 2.38fF
C11831 NOR2X1_LOC_254/a_36_216# INVX1_LOC_186/Y 0.00fF
C11832 NAND2X1_LOC_276/Y NAND2X1_LOC_276/a_36_24# 0.01fF
C11833 INVX1_LOC_90/A NOR2X1_LOC_548/B 0.01fF
C11834 NOR2X1_LOC_389/B NOR2X1_LOC_188/A 0.02fF
C11835 NOR2X1_LOC_383/Y NAND2X1_LOC_642/Y 0.22fF
C11836 INVX1_LOC_18/A NOR2X1_LOC_697/Y 0.02fF
C11837 INVX1_LOC_2/A INVX1_LOC_117/A 0.24fF
C11838 INVX1_LOC_221/A INVX1_LOC_38/A 0.01fF
C11839 NOR2X1_LOC_355/A INVX1_LOC_91/A 0.02fF
C11840 INVX1_LOC_43/A VDD 0.00fF
C11841 D_INPUT_4 NAND2X1_LOC_51/B 5.27fF
C11842 NAND2X1_LOC_735/B NOR2X1_LOC_24/a_36_216# 0.00fF
C11843 INVX1_LOC_34/A NOR2X1_LOC_629/Y 0.03fF
C11844 NAND2X1_LOC_374/Y INVX1_LOC_37/Y 0.01fF
C11845 NOR2X1_LOC_151/Y INVX1_LOC_42/Y 0.03fF
C11846 INVX1_LOC_16/A NAND2X1_LOC_244/A 0.01fF
C11847 INVX1_LOC_208/Y VDD 0.68fF
C11848 NAND2X1_LOC_348/A NOR2X1_LOC_188/A 2.27fF
C11849 NOR2X1_LOC_637/Y NOR2X1_LOC_697/Y 0.03fF
C11850 NOR2X1_LOC_113/B INVX1_LOC_75/A 0.06fF
C11851 INVX1_LOC_299/A INVX1_LOC_4/A 0.31fF
C11852 INVX1_LOC_22/A INVX1_LOC_37/A 0.87fF
C11853 NOR2X1_LOC_458/a_36_216# NOR2X1_LOC_678/A -0.00fF
C11854 NOR2X1_LOC_770/B NAND2X1_LOC_93/B -0.03fF
C11855 NOR2X1_LOC_238/Y INVX1_LOC_119/Y 0.26fF
C11856 NAND2X1_LOC_632/B INVX1_LOC_260/Y 0.00fF
C11857 NAND2X1_LOC_714/B NAND2X1_LOC_175/Y 0.09fF
C11858 INVX1_LOC_36/A INVX1_LOC_29/A 0.30fF
C11859 INVX1_LOC_279/A INVX1_LOC_46/A 0.07fF
C11860 NOR2X1_LOC_770/B NAND2X1_LOC_425/Y -0.01fF
C11861 NOR2X1_LOC_267/A INVX1_LOC_29/A 0.00fF
C11862 INVX1_LOC_193/Y INVX1_LOC_86/A 0.00fF
C11863 NOR2X1_LOC_724/Y NOR2X1_LOC_833/Y 0.16fF
C11864 INVX1_LOC_89/A NOR2X1_LOC_35/Y 0.21fF
C11865 NAND2X1_LOC_181/Y INVX1_LOC_118/A 0.02fF
C11866 NAND2X1_LOC_842/B INVX1_LOC_95/Y 0.07fF
C11867 NOR2X1_LOC_52/Y INVX1_LOC_109/Y 0.29fF
C11868 NAND2X1_LOC_712/A NOR2X1_LOC_694/Y 0.16fF
C11869 NOR2X1_LOC_593/Y NOR2X1_LOC_66/Y 0.24fF
C11870 NAND2X1_LOC_45/Y INVX1_LOC_36/Y 0.06fF
C11871 INVX1_LOC_212/Y NOR2X1_LOC_814/A 0.05fF
C11872 NAND2X1_LOC_862/A INVX1_LOC_54/A 0.01fF
C11873 NOR2X1_LOC_318/B INVX1_LOC_144/A 0.00fF
C11874 NOR2X1_LOC_419/Y INVX1_LOC_19/A 0.03fF
C11875 NOR2X1_LOC_537/A INVX1_LOC_19/A 0.01fF
C11876 NOR2X1_LOC_68/A INVX1_LOC_42/A 0.12fF
C11877 NAND2X1_LOC_377/a_36_24# INVX1_LOC_175/A 0.00fF
C11878 NOR2X1_LOC_733/Y NOR2X1_LOC_741/A 0.02fF
C11879 NOR2X1_LOC_758/a_36_216# NOR2X1_LOC_89/A 0.00fF
C11880 NAND2X1_LOC_357/B INVX1_LOC_285/A 0.02fF
C11881 NOR2X1_LOC_716/B INVX1_LOC_19/A 0.09fF
C11882 INVX1_LOC_28/A NAND2X1_LOC_244/A 0.02fF
C11883 NOR2X1_LOC_67/A NOR2X1_LOC_216/B 0.09fF
C11884 NOR2X1_LOC_237/Y INVX1_LOC_29/A 0.07fF
C11885 NOR2X1_LOC_620/Y NAND2X1_LOC_63/Y 0.20fF
C11886 INVX1_LOC_35/A INVX1_LOC_21/A 1.97fF
C11887 INVX1_LOC_17/A NOR2X1_LOC_720/A 0.15fF
C11888 INVX1_LOC_22/A NOR2X1_LOC_743/Y 0.01fF
C11889 NOR2X1_LOC_756/Y VDD 0.08fF
C11890 NOR2X1_LOC_478/A INVX1_LOC_78/A 0.01fF
C11891 NOR2X1_LOC_804/B INVX1_LOC_29/A 0.07fF
C11892 INVX1_LOC_83/A NOR2X1_LOC_450/A 0.01fF
C11893 INVX1_LOC_182/Y INVX1_LOC_46/A 0.03fF
C11894 NOR2X1_LOC_552/A NOR2X1_LOC_548/a_36_216# 0.01fF
C11895 NAND2X1_LOC_9/Y NAND2X1_LOC_773/Y 0.01fF
C11896 INVX1_LOC_1/Y NOR2X1_LOC_155/A 0.27fF
C11897 NAND2X1_LOC_660/A INVX1_LOC_63/A 0.07fF
C11898 INVX1_LOC_98/A NOR2X1_LOC_78/A 0.08fF
C11899 INVX1_LOC_17/A INVX1_LOC_129/A -0.00fF
C11900 INVX1_LOC_161/Y NOR2X1_LOC_654/A 0.03fF
C11901 INVX1_LOC_77/A NOR2X1_LOC_861/Y 0.05fF
C11902 INVX1_LOC_63/Y INVX1_LOC_12/A 0.34fF
C11903 NOR2X1_LOC_274/B NAND2X1_LOC_72/B 0.07fF
C11904 NOR2X1_LOC_309/Y INVX1_LOC_29/A 0.07fF
C11905 NAND2X1_LOC_77/a_36_24# NAND2X1_LOC_214/B 0.00fF
C11906 INVX1_LOC_136/A NOR2X1_LOC_158/Y 0.01fF
C11907 NAND2X1_LOC_796/B NOR2X1_LOC_186/Y 0.07fF
C11908 NOR2X1_LOC_6/B NAND2X1_LOC_207/B 0.03fF
C11909 INVX1_LOC_298/Y INVX1_LOC_36/A 0.03fF
C11910 INVX1_LOC_299/A INVX1_LOC_64/A 0.03fF
C11911 INVX1_LOC_232/Y NOR2X1_LOC_662/A 0.06fF
C11912 NOR2X1_LOC_67/A NOR2X1_LOC_126/a_36_216# 0.00fF
C11913 INVX1_LOC_17/A INPUT_6 0.04fF
C11914 NOR2X1_LOC_68/A INVX1_LOC_78/A 0.14fF
C11915 INVX1_LOC_45/A NOR2X1_LOC_318/A 0.06fF
C11916 INVX1_LOC_36/A NOR2X1_LOC_281/Y 0.01fF
C11917 INVX1_LOC_226/Y INVX1_LOC_27/Y 0.03fF
C11918 NAND2X1_LOC_214/B NAND2X1_LOC_214/Y 0.02fF
C11919 NAND2X1_LOC_581/a_36_24# NAND2X1_LOC_30/Y 0.00fF
C11920 NOR2X1_LOC_645/a_36_216# NAND2X1_LOC_175/Y 0.01fF
C11921 NOR2X1_LOC_387/A VDD 0.15fF
C11922 NOR2X1_LOC_808/A NOR2X1_LOC_777/B 0.03fF
C11923 NOR2X1_LOC_411/Y INVX1_LOC_269/A 0.00fF
C11924 NAND2X1_LOC_796/B NAND2X1_LOC_573/Y 0.01fF
C11925 INVX1_LOC_303/A INVX1_LOC_104/Y 0.04fF
C11926 INVX1_LOC_33/A NOR2X1_LOC_467/A 0.07fF
C11927 NOR2X1_LOC_706/A NOR2X1_LOC_684/Y 0.04fF
C11928 INVX1_LOC_300/Y NAND2X1_LOC_175/Y 0.15fF
C11929 NAND2X1_LOC_773/Y NOR2X1_LOC_798/A 0.01fF
C11930 NOR2X1_LOC_829/Y INVX1_LOC_36/A 0.04fF
C11931 NAND2X1_LOC_654/B NAND2X1_LOC_637/Y 0.01fF
C11932 NAND2X1_LOC_35/Y NOR2X1_LOC_82/A 0.07fF
C11933 NOR2X1_LOC_389/A INVX1_LOC_53/A 0.14fF
C11934 VDD NOR2X1_LOC_501/B -0.00fF
C11935 NOR2X1_LOC_790/B NOR2X1_LOC_590/A 0.03fF
C11936 INVX1_LOC_235/Y NAND2X1_LOC_393/a_36_24# 0.00fF
C11937 NOR2X1_LOC_542/Y NOR2X1_LOC_862/B 0.05fF
C11938 NOR2X1_LOC_152/Y NAND2X1_LOC_454/Y 0.10fF
C11939 INVX1_LOC_41/Y NOR2X1_LOC_301/A 0.03fF
C11940 NAND2X1_LOC_53/Y INVX1_LOC_5/A 0.03fF
C11941 INVX1_LOC_13/A INVX1_LOC_293/Y 0.04fF
C11942 NOR2X1_LOC_360/Y NOR2X1_LOC_39/Y 0.01fF
C11943 INVX1_LOC_298/Y NOR2X1_LOC_208/Y 0.07fF
C11944 INVX1_LOC_208/Y INVX1_LOC_133/A 0.07fF
C11945 INVX1_LOC_11/A INVX1_LOC_13/Y 0.07fF
C11946 NAND2X1_LOC_786/a_36_24# INVX1_LOC_87/A 0.00fF
C11947 NOR2X1_LOC_188/A INVX1_LOC_38/A 0.13fF
C11948 INVX1_LOC_71/A NOR2X1_LOC_318/A 0.09fF
C11949 NOR2X1_LOC_142/Y INVX1_LOC_4/Y 0.06fF
C11950 INVX1_LOC_272/Y INVX1_LOC_178/A 0.10fF
C11951 NOR2X1_LOC_795/Y INVX1_LOC_15/A 0.04fF
C11952 NOR2X1_LOC_111/A INVX1_LOC_91/A 0.07fF
C11953 INVX1_LOC_45/A NOR2X1_LOC_678/A 0.04fF
C11954 NOR2X1_LOC_455/Y INVX1_LOC_223/A 0.00fF
C11955 NOR2X1_LOC_315/Y INVX1_LOC_4/A 0.08fF
C11956 NAND2X1_LOC_778/Y NAND2X1_LOC_550/A 0.09fF
C11957 NOR2X1_LOC_419/Y INVX1_LOC_26/Y 0.03fF
C11958 NOR2X1_LOC_678/a_36_216# INVX1_LOC_88/A 0.00fF
C11959 INVX1_LOC_2/A INVX1_LOC_3/Y 0.10fF
C11960 NOR2X1_LOC_818/Y INVX1_LOC_3/Y 0.19fF
C11961 INVX1_LOC_21/A NOR2X1_LOC_502/Y 0.01fF
C11962 NAND2X1_LOC_35/Y NAND2X1_LOC_500/Y 0.03fF
C11963 INVX1_LOC_13/A NAND2X1_LOC_74/B 0.62fF
C11964 NOR2X1_LOC_92/Y INVX1_LOC_103/A 0.07fF
C11965 INVX1_LOC_200/Y INVX1_LOC_24/A 0.75fF
C11966 INVX1_LOC_123/A INVX1_LOC_280/A 0.16fF
C11967 INVX1_LOC_107/A INVX1_LOC_53/A 0.01fF
C11968 NOR2X1_LOC_312/Y NOR2X1_LOC_662/A 0.01fF
C11969 NOR2X1_LOC_716/B INVX1_LOC_26/Y 0.08fF
C11970 NOR2X1_LOC_717/B INVX1_LOC_19/A 0.04fF
C11971 NAND2X1_LOC_794/B NAND2X1_LOC_711/Y 0.00fF
C11972 INVX1_LOC_50/A INVX1_LOC_209/Y 0.02fF
C11973 NOR2X1_LOC_596/A INVX1_LOC_53/A 0.09fF
C11974 NOR2X1_LOC_78/B NOR2X1_LOC_38/B 0.07fF
C11975 NOR2X1_LOC_15/Y NAND2X1_LOC_550/A 0.60fF
C11976 NOR2X1_LOC_655/B INVX1_LOC_4/Y 0.19fF
C11977 INVX1_LOC_11/A INVX1_LOC_88/A 0.03fF
C11978 NOR2X1_LOC_309/Y NOR2X1_LOC_281/Y 0.03fF
C11979 INVX1_LOC_58/A INVX1_LOC_49/A 0.22fF
C11980 NOR2X1_LOC_15/Y NOR2X1_LOC_160/B 0.10fF
C11981 NAND2X1_LOC_568/A NAND2X1_LOC_566/a_36_24# 0.02fF
C11982 NOR2X1_LOC_561/Y INVX1_LOC_290/Y 0.10fF
C11983 NOR2X1_LOC_246/A NAND2X1_LOC_74/B 0.07fF
C11984 NOR2X1_LOC_828/A INVX1_LOC_19/A 0.01fF
C11985 INVX1_LOC_71/A NOR2X1_LOC_678/A 0.03fF
C11986 NOR2X1_LOC_483/B INVX1_LOC_1/A 0.01fF
C11987 NOR2X1_LOC_390/a_36_216# NOR2X1_LOC_383/B 0.00fF
C11988 INVX1_LOC_24/Y INVX1_LOC_292/A 0.00fF
C11989 NAND2X1_LOC_15/a_36_24# NOR2X1_LOC_160/B 0.01fF
C11990 NAND2X1_LOC_623/B INVX1_LOC_118/A 0.03fF
C11991 INVX1_LOC_25/A INVX1_LOC_33/A 0.10fF
C11992 NOR2X1_LOC_791/A NOR2X1_LOC_791/Y 0.00fF
C11993 NAND2X1_LOC_551/A NAND2X1_LOC_74/B 0.03fF
C11994 NOR2X1_LOC_405/A NAND2X1_LOC_760/a_36_24# 0.01fF
C11995 NOR2X1_LOC_586/Y INVX1_LOC_117/A 0.03fF
C11996 INVX1_LOC_256/A INVX1_LOC_150/Y 0.91fF
C11997 NAND2X1_LOC_462/B INVX1_LOC_3/Y 0.00fF
C11998 NOR2X1_LOC_763/Y NAND2X1_LOC_430/B 0.02fF
C11999 NOR2X1_LOC_687/Y INVX1_LOC_274/Y 0.53fF
C12000 INVX1_LOC_24/A NOR2X1_LOC_406/A 0.03fF
C12001 INVX1_LOC_297/Y NAND2X1_LOC_175/Y 0.04fF
C12002 NOR2X1_LOC_318/B NOR2X1_LOC_155/A 1.24fF
C12003 NOR2X1_LOC_492/a_36_216# NOR2X1_LOC_492/Y 0.00fF
C12004 INVX1_LOC_22/A NAND2X1_LOC_72/B 0.05fF
C12005 NAND2X1_LOC_724/Y NOR2X1_LOC_504/Y 0.23fF
C12006 INVX1_LOC_27/A INVX1_LOC_181/Y 0.01fF
C12007 NOR2X1_LOC_151/Y INVX1_LOC_19/A 0.09fF
C12008 NOR2X1_LOC_570/Y INVX1_LOC_78/A 0.03fF
C12009 NOR2X1_LOC_45/B NOR2X1_LOC_88/Y 0.03fF
C12010 NAND2X1_LOC_850/Y INVX1_LOC_181/A 0.04fF
C12011 INVX1_LOC_224/A NOR2X1_LOC_500/B 0.03fF
C12012 NOR2X1_LOC_590/A NOR2X1_LOC_785/A 0.01fF
C12013 NOR2X1_LOC_314/Y INVX1_LOC_118/A 0.01fF
C12014 INVX1_LOC_58/A INVX1_LOC_2/A 16.60fF
C12015 NOR2X1_LOC_30/a_36_216# D_INPUT_5 0.00fF
C12016 INVX1_LOC_83/A NOR2X1_LOC_38/B 0.02fF
C12017 NOR2X1_LOC_590/A NAND2X1_LOC_352/B 0.00fF
C12018 INVX1_LOC_11/A NOR2X1_LOC_500/B 0.02fF
C12019 INVX1_LOC_201/A INVX1_LOC_63/A 0.01fF
C12020 NAND2X1_LOC_86/Y NAND2X1_LOC_85/Y 0.07fF
C12021 INVX1_LOC_17/A NOR2X1_LOC_859/A 0.00fF
C12022 INPUT_1 INVX1_LOC_3/Y 0.13fF
C12023 NOR2X1_LOC_13/Y NOR2X1_LOC_321/Y 0.10fF
C12024 INVX1_LOC_13/Y NOR2X1_LOC_593/Y 0.00fF
C12025 INVX1_LOC_58/A NOR2X1_LOC_226/A 0.21fF
C12026 NOR2X1_LOC_99/B INVX1_LOC_4/Y 0.10fF
C12027 INVX1_LOC_64/A NOR2X1_LOC_315/Y 0.01fF
C12028 NOR2X1_LOC_45/B INVX1_LOC_84/A 0.07fF
C12029 NOR2X1_LOC_264/Y INVX1_LOC_50/Y 0.05fF
C12030 NOR2X1_LOC_590/Y NOR2X1_LOC_718/B 0.04fF
C12031 NOR2X1_LOC_275/a_36_216# INVX1_LOC_30/A 0.01fF
C12032 INVX1_LOC_25/A INVX1_LOC_40/A 0.29fF
C12033 NOR2X1_LOC_793/Y NOR2X1_LOC_500/A 0.11fF
C12034 INVX1_LOC_310/A INVX1_LOC_64/A 0.06fF
C12035 NAND2X1_LOC_43/a_36_24# NOR2X1_LOC_554/B 0.00fF
C12036 NOR2X1_LOC_220/A INVX1_LOC_53/A 0.10fF
C12037 NOR2X1_LOC_93/Y INVX1_LOC_34/A 0.12fF
C12038 INVX1_LOC_17/A INVX1_LOC_41/Y 0.03fF
C12039 NAND2X1_LOC_141/Y INVX1_LOC_74/A 0.01fF
C12040 NAND2X1_LOC_175/B NOR2X1_LOC_173/Y 0.14fF
C12041 INVX1_LOC_11/A NOR2X1_LOC_170/a_36_216# 0.00fF
C12042 INVX1_LOC_50/A NOR2X1_LOC_569/Y 0.07fF
C12043 NOR2X1_LOC_558/A NOR2X1_LOC_216/B 0.21fF
C12044 INVX1_LOC_13/Y NOR2X1_LOC_52/B 0.06fF
C12045 NAND2X1_LOC_796/B INVX1_LOC_225/A 0.04fF
C12046 NOR2X1_LOC_71/Y INVX1_LOC_26/A 0.07fF
C12047 NOR2X1_LOC_163/A INVX1_LOC_78/A 0.03fF
C12048 INVX1_LOC_88/A NOR2X1_LOC_433/A 0.39fF
C12049 NAND2X1_LOC_67/a_36_24# INVX1_LOC_34/A 0.00fF
C12050 INVX1_LOC_2/A INVX1_LOC_248/Y 0.02fF
C12051 INVX1_LOC_1/A INVX1_LOC_33/A 0.21fF
C12052 INVX1_LOC_17/A NAND2X1_LOC_593/Y 0.09fF
C12053 INVX1_LOC_303/A INVX1_LOC_11/A 0.07fF
C12054 INVX1_LOC_16/A NOR2X1_LOC_392/Y 0.03fF
C12055 NOR2X1_LOC_548/Y INVX1_LOC_53/A 0.01fF
C12056 INVX1_LOC_45/A INVX1_LOC_305/A 0.07fF
C12057 INVX1_LOC_34/A INVX1_LOC_269/A 0.23fF
C12058 NOR2X1_LOC_92/Y INVX1_LOC_240/A 0.10fF
C12059 NOR2X1_LOC_160/B NOR2X1_LOC_860/B 0.10fF
C12060 NOR2X1_LOC_784/Y INVX1_LOC_33/A 0.03fF
C12061 NOR2X1_LOC_631/B INVX1_LOC_186/Y 0.08fF
C12062 INVX1_LOC_34/A NOR2X1_LOC_232/Y 0.30fF
C12063 NOR2X1_LOC_205/Y NOR2X1_LOC_142/Y 0.05fF
C12064 INVX1_LOC_209/Y NAND2X1_LOC_227/Y 0.04fF
C12065 INVX1_LOC_13/A NOR2X1_LOC_660/Y 0.74fF
C12066 INVX1_LOC_5/A NOR2X1_LOC_500/Y 0.03fF
C12067 INVX1_LOC_140/A NOR2X1_LOC_36/A 1.68fF
C12068 INVX1_LOC_88/A INVX1_LOC_151/A 0.01fF
C12069 INVX1_LOC_226/Y INVX1_LOC_5/A 0.07fF
C12070 INVX1_LOC_11/A NAND2X1_LOC_59/B 0.21fF
C12071 NOR2X1_LOC_312/Y INVX1_LOC_57/A 0.27fF
C12072 INVX1_LOC_13/A NAND2X1_LOC_358/B 0.05fF
C12073 NAND2X1_LOC_564/A NOR2X1_LOC_71/Y 0.05fF
C12074 D_INPUT_1 INVX1_LOC_135/A 0.05fF
C12075 NOR2X1_LOC_769/A NOR2X1_LOC_68/A 0.01fF
C12076 INVX1_LOC_88/A NOR2X1_LOC_52/B 0.18fF
C12077 INVX1_LOC_196/Y NOR2X1_LOC_383/B 0.37fF
C12078 NOR2X1_LOC_773/Y NAND2X1_LOC_474/Y 0.10fF
C12079 NAND2X1_LOC_787/A D_INPUT_0 0.03fF
C12080 NOR2X1_LOC_612/Y NAND2X1_LOC_93/B 0.03fF
C12081 NOR2X1_LOC_82/A NAND2X1_LOC_465/Y 0.03fF
C12082 INVX1_LOC_58/A NAND2X1_LOC_648/A 0.03fF
C12083 INVX1_LOC_103/A NAND2X1_LOC_477/A 0.01fF
C12084 NOR2X1_LOC_478/A INVX1_LOC_113/Y 0.01fF
C12085 INVX1_LOC_41/A INVX1_LOC_292/A 0.12fF
C12086 NAND2X1_LOC_35/Y NOR2X1_LOC_236/a_36_216# 0.00fF
C12087 NOR2X1_LOC_188/A NAND2X1_LOC_223/A 0.07fF
C12088 INVX1_LOC_37/A INVX1_LOC_186/Y 0.07fF
C12089 NAND2X1_LOC_633/Y INVX1_LOC_19/A 0.07fF
C12090 INVX1_LOC_65/A NOR2X1_LOC_850/B 0.09fF
C12091 INVX1_LOC_58/A INPUT_1 0.08fF
C12092 NAND2X1_LOC_363/B D_INPUT_0 0.10fF
C12093 NAND2X1_LOC_784/A INVX1_LOC_90/A 0.01fF
C12094 NOR2X1_LOC_590/A NOR2X1_LOC_344/A 0.04fF
C12095 NAND2X1_LOC_579/A INVX1_LOC_280/Y 0.07fF
C12096 NOR2X1_LOC_468/Y NOR2X1_LOC_78/B 0.07fF
C12097 NOR2X1_LOC_476/a_36_216# NOR2X1_LOC_375/Y 0.00fF
C12098 NOR2X1_LOC_536/A NOR2X1_LOC_673/A 0.03fF
C12099 NOR2X1_LOC_45/B INVX1_LOC_15/A 0.17fF
C12100 INVX1_LOC_45/A NOR2X1_LOC_335/A 0.08fF
C12101 INVX1_LOC_5/A INVX1_LOC_10/A 0.03fF
C12102 INVX1_LOC_166/A INVX1_LOC_135/Y 0.05fF
C12103 NOR2X1_LOC_655/B NOR2X1_LOC_205/Y 0.01fF
C12104 NAND2X1_LOC_190/Y NOR2X1_LOC_78/B 0.05fF
C12105 INVX1_LOC_37/A NOR2X1_LOC_777/B 0.08fF
C12106 NOR2X1_LOC_122/A NOR2X1_LOC_757/Y 0.00fF
C12107 INVX1_LOC_119/A INVX1_LOC_246/A 0.10fF
C12108 NOR2X1_LOC_237/Y NAND2X1_LOC_634/Y 0.10fF
C12109 INVX1_LOC_43/Y NOR2X1_LOC_315/Y -0.01fF
C12110 NOR2X1_LOC_15/Y INVX1_LOC_208/A 0.17fF
C12111 INVX1_LOC_276/A NOR2X1_LOC_513/Y 0.03fF
C12112 D_INPUT_3 NOR2X1_LOC_14/a_36_216# 0.00fF
C12113 NOR2X1_LOC_68/A NOR2X1_LOC_152/Y 0.08fF
C12114 NOR2X1_LOC_437/a_36_216# INVX1_LOC_45/Y 0.02fF
C12115 INVX1_LOC_2/A INVX1_LOC_215/Y 0.03fF
C12116 NAND2X1_LOC_63/Y INVX1_LOC_117/A 0.10fF
C12117 NOR2X1_LOC_289/Y INVX1_LOC_23/A 0.32fF
C12118 NOR2X1_LOC_381/Y INVX1_LOC_316/Y 0.12fF
C12119 NOR2X1_LOC_160/B INVX1_LOC_96/Y 0.19fF
C12120 NOR2X1_LOC_449/a_36_216# NOR2X1_LOC_13/Y 0.12fF
C12121 INVX1_LOC_247/A INVX1_LOC_15/A 0.05fF
C12122 INVX1_LOC_247/Y NOR2X1_LOC_804/B 0.01fF
C12123 INVX1_LOC_256/Y NAND2X1_LOC_793/Y 0.36fF
C12124 NOR2X1_LOC_790/B NOR2X1_LOC_703/A 0.03fF
C12125 INVX1_LOC_36/A INVX1_LOC_8/A 0.14fF
C12126 INVX1_LOC_178/A INVX1_LOC_10/A 0.10fF
C12127 NOR2X1_LOC_292/Y NOR2X1_LOC_383/B 0.03fF
C12128 NAND2X1_LOC_758/a_36_24# INVX1_LOC_105/A 0.00fF
C12129 NOR2X1_LOC_361/B INVX1_LOC_208/Y 0.12fF
C12130 NAND2X1_LOC_198/B NOR2X1_LOC_577/Y 0.03fF
C12131 NOR2X1_LOC_574/a_36_216# INVX1_LOC_31/A 0.00fF
C12132 INVX1_LOC_24/A NOR2X1_LOC_495/Y 0.30fF
C12133 NOR2X1_LOC_349/A NAND2X1_LOC_226/a_36_24# 0.00fF
C12134 NOR2X1_LOC_707/A INVX1_LOC_19/A 0.18fF
C12135 NOR2X1_LOC_97/A INVX1_LOC_57/A 0.02fF
C12136 NOR2X1_LOC_598/B NOR2X1_LOC_742/A 0.03fF
C12137 NAND2X1_LOC_742/a_36_24# NOR2X1_LOC_298/Y 0.08fF
C12138 INVX1_LOC_186/Y NAND2X1_LOC_629/a_36_24# 0.00fF
C12139 NOR2X1_LOC_222/Y INVX1_LOC_174/A 0.07fF
C12140 NOR2X1_LOC_520/A INVX1_LOC_31/A 0.01fF
C12141 NOR2X1_LOC_468/Y NAND2X1_LOC_392/Y 0.06fF
C12142 NOR2X1_LOC_78/B NOR2X1_LOC_389/A 0.08fF
C12143 NAND2X1_LOC_361/Y INVX1_LOC_24/A 0.07fF
C12144 NOR2X1_LOC_865/A INVX1_LOC_29/A 0.05fF
C12145 NOR2X1_LOC_335/A INVX1_LOC_71/A 0.02fF
C12146 NAND2X1_LOC_733/Y NAND2X1_LOC_839/A 0.00fF
C12147 VDD NOR2X1_LOC_620/A 0.00fF
C12148 D_INPUT_1 NOR2X1_LOC_391/B 0.10fF
C12149 INVX1_LOC_160/A NOR2X1_LOC_798/Y 0.11fF
C12150 INVX1_LOC_35/A NAND2X1_LOC_51/B 0.00fF
C12151 NAND2X1_LOC_854/B NOR2X1_LOC_533/Y 0.09fF
C12152 INVX1_LOC_48/Y INVX1_LOC_89/A 0.01fF
C12153 INVX1_LOC_24/A NAND2X1_LOC_799/Y 0.01fF
C12154 NOR2X1_LOC_607/Y NOR2X1_LOC_388/Y 0.20fF
C12155 INVX1_LOC_233/A NAND2X1_LOC_858/B 0.01fF
C12156 NOR2X1_LOC_58/Y INVX1_LOC_63/A 0.03fF
C12157 INVX1_LOC_257/A INVX1_LOC_117/A 0.02fF
C12158 NOR2X1_LOC_67/A NAND2X1_LOC_670/a_36_24# 0.00fF
C12159 NOR2X1_LOC_705/B INVX1_LOC_174/Y 0.09fF
C12160 NOR2X1_LOC_264/Y NOR2X1_LOC_559/B 0.03fF
C12161 INVX1_LOC_163/A NAND2X1_LOC_622/a_36_24# 0.00fF
C12162 INVX1_LOC_90/A NAND2X1_LOC_326/A 0.98fF
C12163 INVX1_LOC_240/A NAND2X1_LOC_837/Y 0.10fF
C12164 NOR2X1_LOC_828/B NAND2X1_LOC_152/a_36_24# 0.00fF
C12165 INVX1_LOC_2/A NOR2X1_LOC_338/Y 0.04fF
C12166 NOR2X1_LOC_620/Y NOR2X1_LOC_624/A 0.16fF
C12167 NOR2X1_LOC_78/B NOR2X1_LOC_317/A 0.01fF
C12168 NOR2X1_LOC_861/Y INVX1_LOC_9/A 0.19fF
C12169 NOR2X1_LOC_435/A INVX1_LOC_29/A 0.03fF
C12170 NOR2X1_LOC_673/A INVX1_LOC_3/A 0.05fF
C12171 NOR2X1_LOC_160/B NOR2X1_LOC_97/B 0.10fF
C12172 NOR2X1_LOC_746/Y INVX1_LOC_23/A 0.01fF
C12173 INVX1_LOC_41/A NAND2X1_LOC_55/a_36_24# 0.02fF
C12174 NOR2X1_LOC_272/Y INVX1_LOC_79/A 0.05fF
C12175 INVX1_LOC_20/A NAND2X1_LOC_99/A 0.07fF
C12176 INVX1_LOC_235/Y INVX1_LOC_75/A 0.01fF
C12177 NOR2X1_LOC_499/B INVX1_LOC_15/A 0.01fF
C12178 INVX1_LOC_268/A INVX1_LOC_72/A 0.02fF
C12179 NOR2X1_LOC_78/B NOR2X1_LOC_596/A 0.25fF
C12180 NAND2X1_LOC_149/Y INVX1_LOC_75/A 0.22fF
C12181 INVX1_LOC_278/A NOR2X1_LOC_45/B 0.08fF
C12182 INVX1_LOC_118/A INVX1_LOC_3/Y 0.09fF
C12183 INVX1_LOC_30/A NAND2X1_LOC_660/Y 0.04fF
C12184 NOR2X1_LOC_389/A INVX1_LOC_83/A 0.01fF
C12185 NAND2X1_LOC_573/Y NAND2X1_LOC_840/Y 0.02fF
C12186 NOR2X1_LOC_212/a_36_216# INVX1_LOC_286/A 0.01fF
C12187 NOR2X1_LOC_498/Y INVX1_LOC_240/A 0.10fF
C12188 NAND2X1_LOC_276/Y INVX1_LOC_60/Y 0.01fF
C12189 INVX1_LOC_13/A INVX1_LOC_136/A 0.01fF
C12190 INVX1_LOC_54/A D_INPUT_5 0.02fF
C12191 INVX1_LOC_90/A NAND2X1_LOC_807/A 0.02fF
C12192 NOR2X1_LOC_264/Y NOR2X1_LOC_6/B 1.52fF
C12193 INVX1_LOC_243/A INVX1_LOC_77/A 0.01fF
C12194 NOR2X1_LOC_843/B INVX1_LOC_37/A 0.03fF
C12195 INVX1_LOC_255/Y NOR2X1_LOC_820/A 0.01fF
C12196 NOR2X1_LOC_437/Y NOR2X1_LOC_757/Y 0.03fF
C12197 INVX1_LOC_77/A INVX1_LOC_179/Y 0.02fF
C12198 NOR2X1_LOC_551/B INVX1_LOC_177/A 0.05fF
C12199 NAND2X1_LOC_198/B INVX1_LOC_22/A 0.06fF
C12200 INVX1_LOC_272/Y INVX1_LOC_140/A 0.10fF
C12201 INVX1_LOC_209/Y INVX1_LOC_209/A 0.02fF
C12202 NAND2X1_LOC_703/Y NAND2X1_LOC_858/B -0.07fF
C12203 INVX1_LOC_58/A NAND2X1_LOC_455/a_36_24# 0.01fF
C12204 INVX1_LOC_35/A INVX1_LOC_304/A 0.07fF
C12205 INVX1_LOC_31/A INVX1_LOC_65/Y 0.50fF
C12206 INVX1_LOC_53/A NAND2X1_LOC_469/B 0.03fF
C12207 NOR2X1_LOC_589/A NAND2X1_LOC_199/a_36_24# 0.00fF
C12208 INVX1_LOC_188/A INVX1_LOC_313/Y -0.02fF
C12209 D_INPUT_0 INVX1_LOC_30/A 0.19fF
C12210 NAND2X1_LOC_287/B INVX1_LOC_57/A 0.09fF
C12211 NOR2X1_LOC_676/Y INVX1_LOC_15/A 0.03fF
C12212 NAND2X1_LOC_74/B NAND2X1_LOC_489/Y 0.03fF
C12213 NOR2X1_LOC_516/B NOR2X1_LOC_860/B 0.10fF
C12214 NOR2X1_LOC_203/Y NOR2X1_LOC_593/Y 0.04fF
C12215 INVX1_LOC_29/A INVX1_LOC_63/A 1.64fF
C12216 NAND2X1_LOC_736/Y NAND2X1_LOC_717/Y 0.06fF
C12217 NAND2X1_LOC_734/B NAND2X1_LOC_721/a_36_24# 0.02fF
C12218 INVX1_LOC_269/A INPUT_0 0.27fF
C12219 INVX1_LOC_36/A NAND2X1_LOC_140/A 0.07fF
C12220 NOR2X1_LOC_186/Y NOR2X1_LOC_78/A 0.03fF
C12221 INVX1_LOC_15/A NOR2X1_LOC_862/B 0.10fF
C12222 INVX1_LOC_50/A NAND2X1_LOC_472/Y 0.07fF
C12223 NOR2X1_LOC_272/Y INVX1_LOC_91/A 0.10fF
C12224 NAND2X1_LOC_563/Y NAND2X1_LOC_570/Y 0.06fF
C12225 NOR2X1_LOC_577/Y INVX1_LOC_53/Y 0.00fF
C12226 INVX1_LOC_136/A NOR2X1_LOC_246/A 0.10fF
C12227 INVX1_LOC_174/A D_INPUT_4 0.05fF
C12228 INVX1_LOC_5/A NOR2X1_LOC_799/B 0.05fF
C12229 INVX1_LOC_34/A NAND2X1_LOC_563/A 0.02fF
C12230 NOR2X1_LOC_447/B INVX1_LOC_53/A 0.08fF
C12231 NAND2X1_LOC_698/a_36_24# INVX1_LOC_26/A 0.00fF
C12232 NOR2X1_LOC_639/B VDD 0.25fF
C12233 NOR2X1_LOC_82/A NOR2X1_LOC_83/Y 0.35fF
C12234 INVX1_LOC_42/A NAND2X1_LOC_768/Y 0.02fF
C12235 D_INPUT_1 NOR2X1_LOC_813/Y 0.08fF
C12236 NOR2X1_LOC_561/Y INVX1_LOC_77/A 0.26fF
C12237 INVX1_LOC_83/A NOR2X1_LOC_596/A 0.09fF
C12238 NOR2X1_LOC_388/Y NOR2X1_LOC_553/Y 0.31fF
C12239 NOR2X1_LOC_401/B NOR2X1_LOC_84/Y 0.00fF
C12240 NOR2X1_LOC_725/A INVX1_LOC_198/A 0.08fF
C12241 NOR2X1_LOC_89/A INVX1_LOC_272/A 0.01fF
C12242 NOR2X1_LOC_403/B INVX1_LOC_135/A 0.14fF
C12243 INVX1_LOC_171/A NAND2X1_LOC_656/A 0.03fF
C12244 INVX1_LOC_135/A D_INPUT_2 0.03fF
C12245 NAND2X1_LOC_530/a_36_24# NOR2X1_LOC_356/A 0.02fF
C12246 NOR2X1_LOC_402/a_36_216# NOR2X1_LOC_84/Y 0.00fF
C12247 NOR2X1_LOC_6/B INVX1_LOC_316/Y 0.02fF
C12248 INVX1_LOC_255/Y INVX1_LOC_315/A 0.01fF
C12249 D_INPUT_1 INVX1_LOC_280/A 0.16fF
C12250 NAND2X1_LOC_9/Y NOR2X1_LOC_98/B 0.00fF
C12251 NAND2X1_LOC_586/a_36_24# INVX1_LOC_90/A 0.00fF
C12252 NOR2X1_LOC_264/Y INVX1_LOC_30/Y 0.37fF
C12253 NAND2X1_LOC_787/A NAND2X1_LOC_848/A 0.03fF
C12254 NAND2X1_LOC_303/Y NAND2X1_LOC_729/B 0.02fF
C12255 INVX1_LOC_64/A NAND2X1_LOC_96/A 0.07fF
C12256 INVX1_LOC_208/A INVX1_LOC_96/Y 0.01fF
C12257 INVX1_LOC_58/A INVX1_LOC_118/A 0.16fF
C12258 NOR2X1_LOC_516/B NAND2X1_LOC_141/A 0.00fF
C12259 INVX1_LOC_89/A NOR2X1_LOC_350/A 0.04fF
C12260 NOR2X1_LOC_78/B NOR2X1_LOC_220/A 0.01fF
C12261 NOR2X1_LOC_778/B NOR2X1_LOC_544/A 0.02fF
C12262 NOR2X1_LOC_830/Y NOR2X1_LOC_850/B 0.26fF
C12263 INVX1_LOC_1/A NOR2X1_LOC_486/Y 0.07fF
C12264 NOR2X1_LOC_331/B NOR2X1_LOC_678/A 0.14fF
C12265 NOR2X1_LOC_468/Y NOR2X1_LOC_368/Y 0.01fF
C12266 INVX1_LOC_269/A NOR2X1_LOC_324/A 0.01fF
C12267 NOR2X1_LOC_454/Y INVX1_LOC_76/A 0.10fF
C12268 NAND2X1_LOC_11/Y NAND2X1_LOC_451/a_36_24# 0.00fF
C12269 NOR2X1_LOC_589/A NOR2X1_LOC_423/Y 0.01fF
C12270 NAND2X1_LOC_724/a_36_24# NAND2X1_LOC_852/Y 0.06fF
C12271 INVX1_LOC_57/A NOR2X1_LOC_809/B 0.14fF
C12272 INVX1_LOC_32/A NAND2X1_LOC_74/B 0.17fF
C12273 NOR2X1_LOC_258/a_36_216# INVX1_LOC_91/A 0.00fF
C12274 INVX1_LOC_124/A NOR2X1_LOC_561/Y 0.10fF
C12275 INVX1_LOC_136/A NOR2X1_LOC_320/Y 0.06fF
C12276 NOR2X1_LOC_619/A NOR2X1_LOC_346/B 0.10fF
C12277 NOR2X1_LOC_299/Y INVX1_LOC_240/A 0.07fF
C12278 NOR2X1_LOC_255/Y INVX1_LOC_89/Y 0.34fF
C12279 INVX1_LOC_34/A NOR2X1_LOC_214/B 0.12fF
C12280 INVX1_LOC_83/A NOR2X1_LOC_844/A 0.03fF
C12281 NOR2X1_LOC_68/A INVX1_LOC_158/Y 0.03fF
C12282 NOR2X1_LOC_516/B INVX1_LOC_226/A 0.03fF
C12283 NOR2X1_LOC_282/Y INVX1_LOC_285/A 0.04fF
C12284 NOR2X1_LOC_78/B NOR2X1_LOC_548/Y 0.05fF
C12285 NOR2X1_LOC_171/Y NAND2X1_LOC_593/Y 0.03fF
C12286 NOR2X1_LOC_468/Y INVX1_LOC_46/A 0.06fF
C12287 NOR2X1_LOC_222/Y NOR2X1_LOC_589/A 0.03fF
C12288 NOR2X1_LOC_281/Y INVX1_LOC_63/A 0.05fF
C12289 NOR2X1_LOC_160/B NAND2X1_LOC_108/a_36_24# 0.00fF
C12290 NAND2X1_LOC_190/Y INVX1_LOC_46/A 0.19fF
C12291 NOR2X1_LOC_78/B NAND2X1_LOC_322/a_36_24# 0.00fF
C12292 INVX1_LOC_25/Y INVX1_LOC_16/A 0.18fF
C12293 NAND2X1_LOC_198/B INVX1_LOC_100/A 0.07fF
C12294 INVX1_LOC_53/Y INVX1_LOC_22/A 0.10fF
C12295 NAND2X1_LOC_222/A NOR2X1_LOC_814/A 0.03fF
C12296 INVX1_LOC_135/A NOR2X1_LOC_87/a_36_216# 0.00fF
C12297 NOR2X1_LOC_336/B INVX1_LOC_91/A 0.04fF
C12298 NAND2X1_LOC_364/A NOR2X1_LOC_114/A 0.01fF
C12299 INVX1_LOC_286/A NOR2X1_LOC_360/Y 0.80fF
C12300 INVX1_LOC_89/A NOR2X1_LOC_84/Y 0.07fF
C12301 INVX1_LOC_33/Y NAND2X1_LOC_780/Y 0.07fF
C12302 INVX1_LOC_239/A INVX1_LOC_166/Y 0.01fF
C12303 NOR2X1_LOC_210/a_36_216# INVX1_LOC_117/A -0.01fF
C12304 NOR2X1_LOC_443/Y NOR2X1_LOC_814/A 0.05fF
C12305 NOR2X1_LOC_773/Y INVX1_LOC_10/A 0.15fF
C12306 INVX1_LOC_1/A NOR2X1_LOC_537/a_36_216# 0.00fF
C12307 NOR2X1_LOC_454/a_36_216# NAND2X1_LOC_51/B 0.00fF
C12308 NAND2X1_LOC_175/Y NAND2X1_LOC_74/B 0.07fF
C12309 INVX1_LOC_120/A INVX1_LOC_64/Y 0.17fF
C12310 INVX1_LOC_83/A INVX1_LOC_189/Y 0.03fF
C12311 INVX1_LOC_28/A NOR2X1_LOC_320/a_36_216# 0.00fF
C12312 NAND2X1_LOC_734/B INVX1_LOC_28/A 0.10fF
C12313 NAND2X1_LOC_364/A INVX1_LOC_91/A 0.08fF
C12314 NAND2X1_LOC_178/a_36_24# NAND2X1_LOC_472/Y 0.01fF
C12315 INVX1_LOC_208/Y NAND2X1_LOC_573/A 0.01fF
C12316 NAND2X1_LOC_563/Y NOR2X1_LOC_19/B 2.03fF
C12317 INVX1_LOC_5/A INVX1_LOC_307/A 0.09fF
C12318 NOR2X1_LOC_787/a_36_216# INVX1_LOC_37/A 0.00fF
C12319 NAND2X1_LOC_326/A INVX1_LOC_38/A 0.82fF
C12320 NOR2X1_LOC_781/B INVX1_LOC_22/A 0.21fF
C12321 INVX1_LOC_47/A NOR2X1_LOC_537/Y 0.08fF
C12322 INVX1_LOC_27/A NAND2X1_LOC_86/a_36_24# 0.00fF
C12323 NAND2X1_LOC_3/B D_INPUT_5 0.11fF
C12324 INVX1_LOC_33/A NOR2X1_LOC_188/A 0.08fF
C12325 INVX1_LOC_31/A INVX1_LOC_36/Y 0.43fF
C12326 NOR2X1_LOC_576/B NAND2X1_LOC_853/Y 0.48fF
C12327 NAND2X1_LOC_577/A INVX1_LOC_20/A 0.03fF
C12328 INVX1_LOC_5/A NOR2X1_LOC_445/B 0.07fF
C12329 NOR2X1_LOC_389/A INVX1_LOC_46/A 0.02fF
C12330 NAND2X1_LOC_618/Y INVX1_LOC_3/Y 0.10fF
C12331 NAND2X1_LOC_332/Y INVX1_LOC_144/A 0.15fF
C12332 INVX1_LOC_72/A INVX1_LOC_95/Y 0.19fF
C12333 INVX1_LOC_72/A INVX1_LOC_187/Y 0.01fF
C12334 INVX1_LOC_33/A NOR2X1_LOC_548/B 0.12fF
C12335 INVX1_LOC_195/Y NAND2X1_LOC_659/B 0.01fF
C12336 NAND2X1_LOC_348/A NOR2X1_LOC_87/B 0.93fF
C12337 NOR2X1_LOC_372/A NAND2X1_LOC_721/A 0.23fF
C12338 NOR2X1_LOC_91/A INVX1_LOC_102/A 1.14fF
C12339 NOR2X1_LOC_465/Y INVX1_LOC_15/A 0.00fF
C12340 INVX1_LOC_90/A NOR2X1_LOC_165/Y 0.00fF
C12341 INVX1_LOC_58/A NAND2X1_LOC_63/Y 0.00fF
C12342 INVX1_LOC_89/A INVX1_LOC_290/A 0.07fF
C12343 INVX1_LOC_52/Y INVX1_LOC_92/A 0.01fF
C12344 INVX1_LOC_136/A NOR2X1_LOC_357/Y 0.06fF
C12345 INVX1_LOC_190/A NOR2X1_LOC_561/Y 0.05fF
C12346 INVX1_LOC_132/A NOR2X1_LOC_78/A 0.11fF
C12347 NOR2X1_LOC_374/A NOR2X1_LOC_78/A 0.71fF
C12348 NOR2X1_LOC_191/A INVX1_LOC_102/Y 0.01fF
C12349 INVX1_LOC_141/Y INVX1_LOC_33/Y 1.69fF
C12350 INVX1_LOC_28/A INVX1_LOC_25/Y 0.07fF
C12351 NOR2X1_LOC_848/Y NOR2X1_LOC_61/Y 0.03fF
C12352 NOR2X1_LOC_431/Y NOR2X1_LOC_56/Y 0.02fF
C12353 INVX1_LOC_308/A NAND2X1_LOC_81/B 0.01fF
C12354 INVX1_LOC_17/A INVX1_LOC_185/A 0.03fF
C12355 INVX1_LOC_195/Y VDD -0.00fF
C12356 NOR2X1_LOC_272/Y NOR2X1_LOC_179/Y 0.27fF
C12357 NOR2X1_LOC_298/Y NAND2X1_LOC_303/B 0.83fF
C12358 INVX1_LOC_229/Y NOR2X1_LOC_380/A 0.25fF
C12359 INVX1_LOC_197/A NAND2X1_LOC_463/B 0.01fF
C12360 INVX1_LOC_58/A NAND2X1_LOC_455/B 0.01fF
C12361 INVX1_LOC_215/Y INVX1_LOC_118/A 0.01fF
C12362 NOR2X1_LOC_173/Y NOR2X1_LOC_697/Y 0.06fF
C12363 NAND2X1_LOC_656/A INVX1_LOC_20/A 0.09fF
C12364 INVX1_LOC_18/A INVX1_LOC_37/A 18.97fF
C12365 NAND2X1_LOC_349/B INVX1_LOC_28/A 0.14fF
C12366 INVX1_LOC_312/Y INVX1_LOC_33/Y 0.01fF
C12367 INVX1_LOC_4/A NAND2X1_LOC_99/A 0.07fF
C12368 NOR2X1_LOC_635/B NOR2X1_LOC_467/A 0.93fF
C12369 NOR2X1_LOC_735/Y NOR2X1_LOC_665/A 0.02fF
C12370 NOR2X1_LOC_589/A NOR2X1_LOC_329/B 0.07fF
C12371 INVX1_LOC_225/A NOR2X1_LOC_78/A 0.07fF
C12372 INVX1_LOC_30/A NAND2X1_LOC_848/A 0.01fF
C12373 INVX1_LOC_62/Y NOR2X1_LOC_98/A -0.00fF
C12374 NAND2X1_LOC_563/A INPUT_0 0.11fF
C12375 INVX1_LOC_54/Y NAND2X1_LOC_103/a_36_24# 0.00fF
C12376 NAND2X1_LOC_338/B NAND2X1_LOC_519/a_36_24# 0.01fF
C12377 INVX1_LOC_75/A INVX1_LOC_16/A 0.10fF
C12378 NOR2X1_LOC_596/A INVX1_LOC_46/A 0.09fF
C12379 NOR2X1_LOC_431/Y VDD 0.23fF
C12380 INVX1_LOC_77/A INVX1_LOC_76/A 0.18fF
C12381 NOR2X1_LOC_837/Y VDD 0.42fF
C12382 NAND2X1_LOC_785/A INVX1_LOC_91/A 0.68fF
C12383 NOR2X1_LOC_637/Y INVX1_LOC_37/A 0.03fF
C12384 INVX1_LOC_111/Y NOR2X1_LOC_355/B 0.33fF
C12385 INVX1_LOC_197/Y NAND2X1_LOC_621/a_36_24# 0.00fF
C12386 INVX1_LOC_5/A INVX1_LOC_12/A 2.03fF
C12387 INVX1_LOC_140/A INVX1_LOC_10/A 0.10fF
C12388 NOR2X1_LOC_245/a_36_216# NAND2X1_LOC_807/Y 0.01fF
C12389 INVX1_LOC_103/A NOR2X1_LOC_435/B 0.03fF
C12390 NOR2X1_LOC_824/A NAND2X1_LOC_500/B 0.03fF
C12391 NAND2X1_LOC_391/a_36_24# INVX1_LOC_280/A 0.01fF
C12392 NAND2X1_LOC_11/Y INVX1_LOC_91/A 0.00fF
C12393 INVX1_LOC_47/Y NOR2X1_LOC_717/A 1.04fF
C12394 INVX1_LOC_32/A NOR2X1_LOC_660/Y 0.04fF
C12395 INVX1_LOC_155/Y VDD 0.33fF
C12396 INVX1_LOC_26/A NOR2X1_LOC_39/Y 2.27fF
C12397 INVX1_LOC_178/A INVX1_LOC_12/A 0.04fF
C12398 INVX1_LOC_13/Y NAND2X1_LOC_254/Y 0.00fF
C12399 NAND2X1_LOC_9/Y NOR2X1_LOC_38/B 0.10fF
C12400 NOR2X1_LOC_86/A INVX1_LOC_309/A 0.40fF
C12401 NOR2X1_LOC_295/Y INVX1_LOC_46/A 0.03fF
C12402 INVX1_LOC_5/A NAND2X1_LOC_253/a_36_24# 0.00fF
C12403 NAND2X1_LOC_338/B INVX1_LOC_95/Y 0.11fF
C12404 INVX1_LOC_59/A INVX1_LOC_284/A 0.01fF
C12405 INVX1_LOC_34/A INVX1_LOC_12/Y 0.03fF
C12406 NAND2X1_LOC_562/B INVX1_LOC_178/Y 0.09fF
C12407 NOR2X1_LOC_71/Y NOR2X1_LOC_368/A 0.31fF
C12408 NOR2X1_LOC_68/A INVX1_LOC_291/A 0.07fF
C12409 NOR2X1_LOC_500/A NOR2X1_LOC_729/A 0.07fF
C12410 NOR2X1_LOC_494/Y INVX1_LOC_12/A 0.05fF
C12411 INVX1_LOC_61/Y NOR2X1_LOC_813/a_36_216# 0.00fF
C12412 NOR2X1_LOC_78/B NAND2X1_LOC_469/B 0.03fF
C12413 NAND2X1_LOC_553/A NOR2X1_LOC_38/B 0.02fF
C12414 INVX1_LOC_39/A INVX1_LOC_3/Y 0.22fF
C12415 INVX1_LOC_8/A NOR2X1_LOC_102/a_36_216# 0.01fF
C12416 INVX1_LOC_11/A INVX1_LOC_272/A 0.07fF
C12417 INVX1_LOC_28/A INVX1_LOC_75/A 0.10fF
C12418 VDD NOR2X1_LOC_822/Y 0.32fF
C12419 NOR2X1_LOC_420/a_36_216# INVX1_LOC_4/Y 0.12fF
C12420 INVX1_LOC_90/A NOR2X1_LOC_815/A 0.01fF
C12421 VDD NOR2X1_LOC_131/A 0.00fF
C12422 INVX1_LOC_181/Y NOR2X1_LOC_216/B 0.01fF
C12423 NOR2X1_LOC_13/Y NAND2X1_LOC_798/B 0.10fF
C12424 D_GATE_366 INVX1_LOC_6/A 0.05fF
C12425 INVX1_LOC_272/Y INVX1_LOC_42/A 0.00fF
C12426 NOR2X1_LOC_816/A INVX1_LOC_12/A 0.03fF
C12427 INVX1_LOC_64/A NAND2X1_LOC_99/A 0.01fF
C12428 INPUT_3 NAND2X1_LOC_74/B 0.05fF
C12429 INVX1_LOC_75/A NAND2X1_LOC_126/a_36_24# -0.00fF
C12430 INPUT_3 NAND2X1_LOC_207/Y 0.02fF
C12431 NOR2X1_LOC_637/A NOR2X1_LOC_697/Y 0.01fF
C12432 INVX1_LOC_229/Y INPUT_4 0.00fF
C12433 NOR2X1_LOC_816/A NOR2X1_LOC_519/Y 0.01fF
C12434 INVX1_LOC_22/A NOR2X1_LOC_585/Y 0.29fF
C12435 NOR2X1_LOC_572/a_36_216# INVX1_LOC_59/Y 0.00fF
C12436 NOR2X1_LOC_278/Y INVX1_LOC_306/Y 0.01fF
C12437 INVX1_LOC_136/A NAND2X1_LOC_489/Y 0.02fF
C12438 NOR2X1_LOC_464/B INVX1_LOC_4/A 0.06fF
C12439 INVX1_LOC_16/A NAND2X1_LOC_453/A 0.03fF
C12440 NAND2X1_LOC_474/Y INVX1_LOC_78/A 0.07fF
C12441 NAND2X1_LOC_863/B INVX1_LOC_46/A 0.06fF
C12442 NOR2X1_LOC_87/a_36_216# INVX1_LOC_280/A 0.01fF
C12443 INPUT_3 NOR2X1_LOC_847/B -0.00fF
C12444 INVX1_LOC_63/Y INVX1_LOC_92/A 0.08fF
C12445 NAND2X1_LOC_361/Y NOR2X1_LOC_197/B 0.03fF
C12446 INVX1_LOC_31/A INVX1_LOC_102/A 0.07fF
C12447 INVX1_LOC_83/A NAND2X1_LOC_655/B 0.06fF
C12448 INVX1_LOC_22/A INVX1_LOC_77/Y 0.10fF
C12449 NOR2X1_LOC_329/B NOR2X1_LOC_311/a_36_216# 0.01fF
C12450 NAND2X1_LOC_863/B NOR2X1_LOC_766/Y 0.02fF
C12451 NOR2X1_LOC_65/B NAND2X1_LOC_474/Y 0.00fF
C12452 INVX1_LOC_50/Y INVX1_LOC_57/A 0.12fF
C12453 NOR2X1_LOC_380/A INVX1_LOC_20/A 0.00fF
C12454 NOR2X1_LOC_165/Y INVX1_LOC_38/A 0.10fF
C12455 INVX1_LOC_104/A NOR2X1_LOC_831/B 0.10fF
C12456 INVX1_LOC_272/Y INVX1_LOC_78/A 0.56fF
C12457 NOR2X1_LOC_487/a_36_216# NOR2X1_LOC_89/A 0.01fF
C12458 INVX1_LOC_35/A NOR2X1_LOC_400/A 0.02fF
C12459 INVX1_LOC_58/A NOR2X1_LOC_272/a_36_216# 0.03fF
C12460 NOR2X1_LOC_392/B NAND2X1_LOC_572/B 0.10fF
C12461 NAND2X1_LOC_53/Y INVX1_LOC_78/A 0.10fF
C12462 INVX1_LOC_201/Y NAND2X1_LOC_659/A 2.41fF
C12463 INVX1_LOC_58/A INVX1_LOC_39/A 0.05fF
C12464 INVX1_LOC_1/A NOR2X1_LOC_798/Y 0.02fF
C12465 NOR2X1_LOC_341/a_36_216# NAND2X1_LOC_63/Y 0.01fF
C12466 INVX1_LOC_244/Y NOR2X1_LOC_583/Y 0.03fF
C12467 INVX1_LOC_21/A NOR2X1_LOC_456/Y 0.07fF
C12468 NOR2X1_LOC_92/Y NOR2X1_LOC_677/Y 0.01fF
C12469 INVX1_LOC_8/A INVX1_LOC_63/A 0.17fF
C12470 NOR2X1_LOC_433/A INVX1_LOC_272/A 2.52fF
C12471 NOR2X1_LOC_329/B INVX1_LOC_20/A 0.07fF
C12472 INVX1_LOC_1/A NOR2X1_LOC_748/A 0.01fF
C12473 INVX1_LOC_136/A INVX1_LOC_32/A 6.63fF
C12474 NOR2X1_LOC_561/Y INVX1_LOC_9/A 0.10fF
C12475 INVX1_LOC_28/A NAND2X1_LOC_453/A 0.07fF
C12476 NOR2X1_LOC_52/Y INVX1_LOC_15/A 0.04fF
C12477 INVX1_LOC_7/A INVX1_LOC_9/A 0.07fF
C12478 INVX1_LOC_28/A NOR2X1_LOC_65/a_36_216# 0.00fF
C12479 INVX1_LOC_75/A NOR2X1_LOC_35/Y 0.08fF
C12480 NOR2X1_LOC_270/Y INVX1_LOC_15/A 0.01fF
C12481 INVX1_LOC_255/Y NOR2X1_LOC_660/a_36_216# 0.00fF
C12482 NAND2X1_LOC_21/Y NOR2X1_LOC_1/Y 0.06fF
C12483 INVX1_LOC_17/A INVX1_LOC_270/Y 0.17fF
C12484 INVX1_LOC_287/A NAND2X1_LOC_700/a_36_24# 0.00fF
C12485 INVX1_LOC_48/Y NOR2X1_LOC_392/Y 0.02fF
C12486 INVX1_LOC_43/Y NAND2X1_LOC_99/A 0.02fF
C12487 NAND2X1_LOC_9/Y NOR2X1_LOC_468/Y 0.07fF
C12488 INVX1_LOC_302/A VDD 0.00fF
C12489 INVX1_LOC_151/A INVX1_LOC_272/A 0.07fF
C12490 NOR2X1_LOC_405/A NOR2X1_LOC_114/A 0.03fF
C12491 NOR2X1_LOC_532/a_36_216# NAND2X1_LOC_72/B 0.00fF
C12492 NAND2X1_LOC_56/a_36_24# NOR2X1_LOC_727/B 0.00fF
C12493 INVX1_LOC_233/A NOR2X1_LOC_468/Y 0.03fF
C12494 INVX1_LOC_233/Y NAND2X1_LOC_579/A 0.10fF
C12495 NOR2X1_LOC_770/B NOR2X1_LOC_89/A 0.00fF
C12496 NAND2X1_LOC_656/A INVX1_LOC_4/A 0.30fF
C12497 NOR2X1_LOC_794/B NOR2X1_LOC_748/A 0.03fF
C12498 NOR2X1_LOC_52/B INVX1_LOC_272/A 0.22fF
C12499 INVX1_LOC_98/A NAND2X1_LOC_642/Y 0.01fF
C12500 INVX1_LOC_135/A NOR2X1_LOC_61/Y 0.07fF
C12501 NAND2X1_LOC_545/a_36_24# INVX1_LOC_78/A 0.00fF
C12502 INVX1_LOC_140/A NOR2X1_LOC_301/a_36_216# 0.04fF
C12503 INVX1_LOC_18/A NAND2X1_LOC_72/B 0.09fF
C12504 NOR2X1_LOC_405/A INVX1_LOC_91/A 0.21fF
C12505 NOR2X1_LOC_377/Y INVX1_LOC_12/A 0.01fF
C12506 INVX1_LOC_35/A NOR2X1_LOC_523/A 0.00fF
C12507 NOR2X1_LOC_443/Y NOR2X1_LOC_590/A 0.00fF
C12508 INVX1_LOC_136/A NAND2X1_LOC_175/Y 0.19fF
C12509 NOR2X1_LOC_67/A NOR2X1_LOC_721/B 0.13fF
C12510 NAND2X1_LOC_562/B INVX1_LOC_12/A 0.49fF
C12511 NOR2X1_LOC_78/A NAND2X1_LOC_642/Y 0.11fF
C12512 NOR2X1_LOC_792/B NAND2X1_LOC_807/B 0.00fF
C12513 INVX1_LOC_64/A NAND2X1_LOC_192/B 0.04fF
C12514 NOR2X1_LOC_186/Y NAND2X1_LOC_573/Y 0.72fF
C12515 NOR2X1_LOC_234/a_36_216# NAND2X1_LOC_254/Y 0.00fF
C12516 INVX1_LOC_198/Y INVX1_LOC_271/Y 0.05fF
C12517 NOR2X1_LOC_139/Y NOR2X1_LOC_657/B 0.08fF
C12518 NAND2X1_LOC_553/A NOR2X1_LOC_468/Y 0.00fF
C12519 INPUT_0 INVX1_LOC_12/Y 1.05fF
C12520 NOR2X1_LOC_643/A INVX1_LOC_5/A 0.00fF
C12521 NOR2X1_LOC_811/B NOR2X1_LOC_777/B 0.04fF
C12522 NOR2X1_LOC_311/Y NAND2X1_LOC_655/B 0.01fF
C12523 NOR2X1_LOC_72/a_36_216# NAND2X1_LOC_93/B 0.00fF
C12524 NOR2X1_LOC_219/Y INVX1_LOC_186/Y 0.01fF
C12525 NOR2X1_LOC_798/A NOR2X1_LOC_468/Y 0.00fF
C12526 INVX1_LOC_30/A NOR2X1_LOC_451/a_36_216# 0.01fF
C12527 INVX1_LOC_176/A NOR2X1_LOC_845/A 0.26fF
C12528 INVX1_LOC_35/A INVX1_LOC_174/A 0.05fF
C12529 INVX1_LOC_200/A NAND2X1_LOC_552/A 0.30fF
C12530 NOR2X1_LOC_248/Y INVX1_LOC_57/A 0.10fF
C12531 INPUT_3 NOR2X1_LOC_660/Y 0.60fF
C12532 NOR2X1_LOC_86/A INVX1_LOC_203/A 0.10fF
C12533 NOR2X1_LOC_824/A NAND2X1_LOC_725/B 0.12fF
C12534 NOR2X1_LOC_657/B NAND2X1_LOC_468/B 0.15fF
C12535 NOR2X1_LOC_550/a_36_216# INVX1_LOC_53/A 0.01fF
C12536 NOR2X1_LOC_92/Y INVX1_LOC_234/Y 0.04fF
C12537 NOR2X1_LOC_773/Y INVX1_LOC_12/A 0.07fF
C12538 INVX1_LOC_223/A INVX1_LOC_23/A 0.09fF
C12539 NOR2X1_LOC_180/Y INVX1_LOC_15/A 0.05fF
C12540 NAND2X1_LOC_575/a_36_24# NAND2X1_LOC_703/Y 0.00fF
C12541 NAND2X1_LOC_725/B INVX1_LOC_237/A 0.06fF
C12542 NOR2X1_LOC_93/a_36_216# INVX1_LOC_3/Y 0.01fF
C12543 NAND2X1_LOC_451/Y NOR2X1_LOC_48/B 0.04fF
C12544 INVX1_LOC_41/Y INVX1_LOC_181/A 0.25fF
C12545 INVX1_LOC_1/Y INVX1_LOC_29/A 0.15fF
C12546 NAND2X1_LOC_560/A NOR2X1_LOC_823/a_36_216# 0.00fF
C12547 INVX1_LOC_64/A NAND2X1_LOC_577/A 0.03fF
C12548 NAND2X1_LOC_564/B NAND2X1_LOC_74/B 2.77fF
C12549 INVX1_LOC_90/A NAND2X1_LOC_572/B 0.06fF
C12550 INVX1_LOC_58/A INVX1_LOC_61/A 0.13fF
C12551 INVX1_LOC_50/A INVX1_LOC_24/A 2.16fF
C12552 NOR2X1_LOC_500/Y INVX1_LOC_42/A 0.07fF
C12553 NOR2X1_LOC_473/B NOR2X1_LOC_127/Y 0.32fF
C12554 INVX1_LOC_226/Y INVX1_LOC_42/A 0.25fF
C12555 NOR2X1_LOC_427/Y INVX1_LOC_54/A 0.00fF
C12556 NOR2X1_LOC_187/Y NOR2X1_LOC_205/Y 0.01fF
C12557 NAND2X1_LOC_300/a_36_24# NOR2X1_LOC_301/A 0.02fF
C12558 NOR2X1_LOC_354/Y NOR2X1_LOC_729/A 0.02fF
C12559 NOR2X1_LOC_802/A NOR2X1_LOC_334/Y 0.07fF
C12560 NAND2X1_LOC_469/B INVX1_LOC_46/A 0.03fF
C12561 NOR2X1_LOC_710/B INVX1_LOC_1/A 0.15fF
C12562 INVX1_LOC_11/A INVX1_LOC_198/A 0.02fF
C12563 NOR2X1_LOC_559/B INVX1_LOC_57/A 0.03fF
C12564 INVX1_LOC_134/Y NOR2X1_LOC_839/B 0.04fF
C12565 INVX1_LOC_11/A NOR2X1_LOC_271/B 0.03fF
C12566 NOR2X1_LOC_458/B INVX1_LOC_15/A 0.01fF
C12567 NAND2X1_LOC_9/Y INVX1_LOC_62/Y 0.71fF
C12568 NOR2X1_LOC_433/A NOR2X1_LOC_125/a_36_216# 0.01fF
C12569 INVX1_LOC_279/A NOR2X1_LOC_755/Y -0.00fF
C12570 NOR2X1_LOC_78/A NOR2X1_LOC_271/Y 0.03fF
C12571 NAND2X1_LOC_568/A NOR2X1_LOC_533/Y 0.01fF
C12572 NAND2X1_LOC_212/Y INVX1_LOC_117/A 0.02fF
C12573 INVX1_LOC_6/A INVX1_LOC_70/A 0.03fF
C12574 NOR2X1_LOC_332/A INVX1_LOC_12/A 0.08fF
C12575 INVX1_LOC_5/A INVX1_LOC_217/A 0.00fF
C12576 NOR2X1_LOC_91/A INVX1_LOC_162/Y 0.03fF
C12577 INVX1_LOC_269/A INVX1_LOC_225/Y 0.10fF
C12578 INVX1_LOC_10/A INVX1_LOC_42/A 0.01fF
C12579 NAND2X1_LOC_746/a_36_24# INVX1_LOC_159/A 0.00fF
C12580 NOR2X1_LOC_269/Y INVX1_LOC_54/A 0.07fF
C12581 NAND2X1_LOC_735/B INVX1_LOC_3/Y 0.00fF
C12582 INVX1_LOC_272/Y NOR2X1_LOC_503/Y 0.12fF
C12583 INVX1_LOC_286/A NOR2X1_LOC_79/Y 0.03fF
C12584 INVX1_LOC_136/A INVX1_LOC_171/Y 0.02fF
C12585 NAND2X1_LOC_363/B INVX1_LOC_49/A 0.07fF
C12586 NAND2X1_LOC_397/a_36_24# NAND2X1_LOC_577/A 0.01fF
C12587 INVX1_LOC_89/A INVX1_LOC_114/Y 0.01fF
C12588 INVX1_LOC_178/A INVX1_LOC_217/A 0.10fF
C12589 NOR2X1_LOC_6/B INVX1_LOC_57/A 0.10fF
C12590 INVX1_LOC_14/Y INVX1_LOC_117/A 0.11fF
C12591 INVX1_LOC_149/Y INVX1_LOC_23/A 0.00fF
C12592 NOR2X1_LOC_500/Y INVX1_LOC_78/A 0.07fF
C12593 INVX1_LOC_63/Y INVX1_LOC_53/A 0.09fF
C12594 INVX1_LOC_226/Y INVX1_LOC_78/A 0.03fF
C12595 NAND2X1_LOC_348/A NAND2X1_LOC_219/B 0.05fF
C12596 INVX1_LOC_13/Y INVX1_LOC_314/Y 0.07fF
C12597 NOR2X1_LOC_434/Y INVX1_LOC_77/A 0.03fF
C12598 NOR2X1_LOC_15/Y INVX1_LOC_195/A 0.01fF
C12599 INVX1_LOC_76/A INVX1_LOC_9/A 0.14fF
C12600 NOR2X1_LOC_709/A INVX1_LOC_29/Y 0.07fF
C12601 INVX1_LOC_140/A INVX1_LOC_12/A 0.05fF
C12602 INVX1_LOC_50/A INVX1_LOC_143/A 0.07fF
C12603 NOR2X1_LOC_790/B INVX1_LOC_104/A 0.00fF
C12604 INVX1_LOC_182/Y NOR2X1_LOC_755/Y 0.01fF
C12605 NAND2X1_LOC_767/a_36_24# INVX1_LOC_31/A 0.00fF
C12606 NAND2X1_LOC_30/Y INVX1_LOC_30/A 0.03fF
C12607 INVX1_LOC_89/A NOR2X1_LOC_467/A 0.24fF
C12608 NOR2X1_LOC_160/B NAND2X1_LOC_208/B 0.01fF
C12609 NOR2X1_LOC_65/B INVX1_LOC_226/Y 0.14fF
C12610 INVX1_LOC_21/A NOR2X1_LOC_550/B 0.02fF
C12611 INVX1_LOC_10/A INVX1_LOC_78/A 0.21fF
C12612 NOR2X1_LOC_84/Y NOR2X1_LOC_392/Y 0.02fF
C12613 NAND2X1_LOC_763/B NAND2X1_LOC_30/Y 0.03fF
C12614 INVX1_LOC_2/A NAND2X1_LOC_787/A 0.04fF
C12615 NAND2X1_LOC_35/Y INVX1_LOC_240/A 0.10fF
C12616 NOR2X1_LOC_634/a_36_216# NOR2X1_LOC_798/A 0.00fF
C12617 NOR2X1_LOC_71/Y NAND2X1_LOC_471/Y 0.02fF
C12618 INVX1_LOC_2/A NAND2X1_LOC_363/B 0.01fF
C12619 NOR2X1_LOC_817/Y NOR2X1_LOC_820/A 0.01fF
C12620 NOR2X1_LOC_445/a_36_216# NOR2X1_LOC_568/A 0.00fF
C12621 NAND2X1_LOC_774/a_36_24# INVX1_LOC_111/A 0.01fF
C12622 NOR2X1_LOC_134/Y INVX1_LOC_30/A 0.14fF
C12623 NOR2X1_LOC_602/A NOR2X1_LOC_590/A 0.01fF
C12624 NOR2X1_LOC_226/A NAND2X1_LOC_787/A 0.02fF
C12625 INVX1_LOC_304/Y NAND2X1_LOC_552/A 0.02fF
C12626 INVX1_LOC_278/A NOR2X1_LOC_401/Y 0.01fF
C12627 NOR2X1_LOC_188/A INVX1_LOC_106/Y 0.13fF
C12628 NOR2X1_LOC_32/B INVX1_LOC_280/Y 0.18fF
C12629 NOR2X1_LOC_186/Y INVX1_LOC_225/A 0.44fF
C12630 INVX1_LOC_217/A NOR2X1_LOC_816/A 0.01fF
C12631 NOR2X1_LOC_598/B NOR2X1_LOC_731/Y 0.00fF
C12632 INPUT_0 NOR2X1_LOC_842/a_36_216# 0.02fF
C12633 NAND2X1_LOC_682/a_36_24# INVX1_LOC_19/A 0.00fF
C12634 INVX1_LOC_30/Y INVX1_LOC_57/A 0.12fF
C12635 NOR2X1_LOC_494/Y NAND2X1_LOC_787/B 0.17fF
C12636 NOR2X1_LOC_753/Y NAND2X1_LOC_537/Y 0.00fF
C12637 NOR2X1_LOC_65/B INVX1_LOC_10/A 0.09fF
C12638 INVX1_LOC_64/A NOR2X1_LOC_222/Y 0.04fF
C12639 NOR2X1_LOC_6/B INVX1_LOC_252/A 0.03fF
C12640 NOR2X1_LOC_92/Y NAND2X1_LOC_673/a_36_24# 0.01fF
C12641 INPUT_0 NOR2X1_LOC_554/A 0.00fF
C12642 INVX1_LOC_304/Y INVX1_LOC_178/A 0.10fF
C12643 NOR2X1_LOC_471/Y NOR2X1_LOC_257/a_36_216# 0.00fF
C12644 INVX1_LOC_251/Y NOR2X1_LOC_652/Y 0.00fF
C12645 NAND2X1_LOC_775/a_36_24# INVX1_LOC_93/A 0.01fF
C12646 NOR2X1_LOC_318/B INVX1_LOC_29/A 0.43fF
C12647 INVX1_LOC_50/A NAND2X1_LOC_783/A 0.15fF
C12648 NOR2X1_LOC_667/A NAND2X1_LOC_542/a_36_24# 0.00fF
C12649 NOR2X1_LOC_61/Y INVX1_LOC_280/A 0.01fF
C12650 INVX1_LOC_58/A INPUT_5 0.02fF
C12651 NAND2X1_LOC_537/Y NAND2X1_LOC_325/Y 0.00fF
C12652 INVX1_LOC_269/A NOR2X1_LOC_514/a_36_216# 0.01fF
C12653 NAND2X1_LOC_479/Y NOR2X1_LOC_678/A 0.11fF
C12654 NAND2X1_LOC_53/Y INVX1_LOC_113/Y 0.03fF
C12655 NOR2X1_LOC_445/a_36_216# INVX1_LOC_71/A 0.00fF
C12656 INVX1_LOC_50/A NOR2X1_LOC_130/A 0.03fF
C12657 INVX1_LOC_24/A INVX1_LOC_61/Y 0.09fF
C12658 INVX1_LOC_25/A NOR2X1_LOC_719/a_36_216# 0.00fF
C12659 NOR2X1_LOC_457/B NOR2X1_LOC_717/Y 0.00fF
C12660 INVX1_LOC_93/Y INVX1_LOC_29/A 0.08fF
C12661 NAND2X1_LOC_517/a_36_24# NAND2X1_LOC_114/B 0.00fF
C12662 INVX1_LOC_35/A NOR2X1_LOC_589/A 0.10fF
C12663 NOR2X1_LOC_798/A NOR2X1_LOC_220/A 0.00fF
C12664 INVX1_LOC_186/A NOR2X1_LOC_640/B 0.05fF
C12665 INVX1_LOC_21/A NAND2X1_LOC_526/a_36_24# 0.00fF
C12666 NOR2X1_LOC_815/Y INVX1_LOC_215/Y 0.02fF
C12667 NOR2X1_LOC_817/Y INVX1_LOC_315/A 0.10fF
C12668 INVX1_LOC_90/A NOR2X1_LOC_654/A 0.05fF
C12669 INVX1_LOC_66/Y NOR2X1_LOC_117/a_36_216# 0.01fF
C12670 NAND2X1_LOC_392/A INVX1_LOC_306/Y 0.00fF
C12671 NOR2X1_LOC_426/Y NOR2X1_LOC_95/a_36_216# 0.00fF
C12672 NOR2X1_LOC_703/Y NOR2X1_LOC_801/B 0.00fF
C12673 INVX1_LOC_298/Y NOR2X1_LOC_742/A 0.07fF
C12674 INVX1_LOC_25/A INVX1_LOC_89/A 0.06fF
C12675 INVX1_LOC_248/A NAND2X1_LOC_714/B 0.02fF
C12676 INVX1_LOC_34/A NAND2X1_LOC_550/A 0.09fF
C12677 INVX1_LOC_34/A NOR2X1_LOC_160/B 11.29fF
C12678 NAND2X1_LOC_773/Y NAND2X1_LOC_338/B 0.28fF
C12679 NOR2X1_LOC_548/A NAND2X1_LOC_72/B 0.01fF
C12680 NAND2X1_LOC_807/Y NOR2X1_LOC_280/a_36_216# 0.01fF
C12681 INVX1_LOC_276/A NAND2X1_LOC_537/Y 0.27fF
C12682 NOR2X1_LOC_74/A NOR2X1_LOC_278/Y 0.07fF
C12683 NOR2X1_LOC_66/a_36_216# INVX1_LOC_4/A 0.00fF
C12684 INVX1_LOC_150/Y NOR2X1_LOC_52/B 0.07fF
C12685 INVX1_LOC_49/A INVX1_LOC_30/A 0.19fF
C12686 NOR2X1_LOC_538/B NOR2X1_LOC_538/Y 0.01fF
C12687 INVX1_LOC_35/A INVX1_LOC_171/A 0.01fF
C12688 NAND2X1_LOC_787/a_36_24# NAND2X1_LOC_722/A 0.00fF
C12689 NAND2X1_LOC_564/B NAND2X1_LOC_793/a_36_24# 0.00fF
C12690 NAND2X1_LOC_787/A INPUT_1 0.03fF
C12691 NOR2X1_LOC_501/B INVX1_LOC_4/Y 0.05fF
C12692 NAND2X1_LOC_114/B NAND2X1_LOC_116/A 0.04fF
C12693 INVX1_LOC_90/A INVX1_LOC_58/Y 0.07fF
C12694 NAND2X1_LOC_352/B INVX1_LOC_104/A 0.32fF
C12695 INVX1_LOC_48/Y INVX1_LOC_25/Y 1.71fF
C12696 NAND2X1_LOC_149/Y INVX1_LOC_22/A 0.17fF
C12697 NAND2X1_LOC_552/A NAND2X1_LOC_808/A 0.06fF
C12698 NOR2X1_LOC_606/a_36_216# INVX1_LOC_8/A 0.01fF
C12699 INVX1_LOC_50/A NOR2X1_LOC_216/Y 0.03fF
C12700 NAND2X1_LOC_763/B INVX1_LOC_49/A 0.05fF
C12701 INVX1_LOC_2/A NOR2X1_LOC_457/A 0.06fF
C12702 INVX1_LOC_31/A INVX1_LOC_149/Y 0.09fF
C12703 NOR2X1_LOC_92/Y INVX1_LOC_56/Y 0.07fF
C12704 NAND2X1_LOC_624/B NAND2X1_LOC_624/A 0.01fF
C12705 INVX1_LOC_77/Y INVX1_LOC_261/A 0.04fF
C12706 INVX1_LOC_118/Y INVX1_LOC_63/A 0.02fF
C12707 NAND2X1_LOC_53/Y NOR2X1_LOC_307/B 0.06fF
C12708 INVX1_LOC_41/A NAND2X1_LOC_351/A 0.01fF
C12709 INVX1_LOC_286/A INVX1_LOC_26/A 0.82fF
C12710 INVX1_LOC_34/A NAND2X1_LOC_195/Y 0.03fF
C12711 INVX1_LOC_214/Y NOR2X1_LOC_816/A 0.05fF
C12712 NAND2X1_LOC_784/A NOR2X1_LOC_323/Y 0.01fF
C12713 INVX1_LOC_178/A NAND2X1_LOC_808/A 0.10fF
C12714 NOR2X1_LOC_112/Y INVX1_LOC_68/A 0.00fF
C12715 INVX1_LOC_64/A NOR2X1_LOC_329/B 0.10fF
C12716 NAND2X1_LOC_798/B NOR2X1_LOC_697/Y 0.00fF
C12717 NAND2X1_LOC_93/B NOR2X1_LOC_450/B 0.04fF
C12718 INVX1_LOC_248/A NAND2X1_LOC_336/a_36_24# 0.00fF
C12719 INVX1_LOC_303/A INVX1_LOC_314/Y 0.07fF
C12720 INVX1_LOC_298/Y NOR2X1_LOC_318/B 0.02fF
C12721 NOR2X1_LOC_274/Y INVX1_LOC_77/A 0.01fF
C12722 INVX1_LOC_24/A NOR2X1_LOC_679/B 0.01fF
C12723 D_INPUT_3 INVX1_LOC_3/Y 1.34fF
C12724 NAND2X1_LOC_562/B INVX1_LOC_217/A 0.01fF
C12725 INVX1_LOC_2/A INVX1_LOC_30/A 0.37fF
C12726 INVX1_LOC_54/A NOR2X1_LOC_36/B 0.01fF
C12727 NAND2X1_LOC_425/Y NOR2X1_LOC_450/B 0.10fF
C12728 NAND2X1_LOC_93/B NOR2X1_LOC_257/Y 0.02fF
C12729 NAND2X1_LOC_733/Y NOR2X1_LOC_773/Y 0.10fF
C12730 NOR2X1_LOC_355/B NOR2X1_LOC_383/B 0.01fF
C12731 NOR2X1_LOC_226/A INVX1_LOC_30/A 0.42fF
C12732 INVX1_LOC_95/A INVX1_LOC_26/A 0.01fF
C12733 NAND2X1_LOC_9/Y INVX1_LOC_51/Y 0.05fF
C12734 NAND2X1_LOC_574/A NAND2X1_LOC_659/A 0.12fF
C12735 NOR2X1_LOC_643/A NOR2X1_LOC_332/A 0.01fF
C12736 NAND2X1_LOC_231/Y NAND2X1_LOC_195/Y 0.02fF
C12737 INVX1_LOC_182/Y NOR2X1_LOC_674/Y 0.05fF
C12738 INVX1_LOC_35/A INVX1_LOC_222/A 0.16fF
C12739 INVX1_LOC_255/Y INVX1_LOC_230/Y 0.05fF
C12740 NAND2X1_LOC_425/Y NOR2X1_LOC_257/Y 0.01fF
C12741 NAND2X1_LOC_543/Y INVX1_LOC_31/A 0.03fF
C12742 INVX1_LOC_58/A NOR2X1_LOC_7/Y 0.01fF
C12743 INVX1_LOC_1/A INVX1_LOC_89/A 0.47fF
C12744 NOR2X1_LOC_315/Y INVX1_LOC_41/Y 0.00fF
C12745 INVX1_LOC_228/Y NOR2X1_LOC_332/A 0.03fF
C12746 NOR2X1_LOC_45/B NAND2X1_LOC_231/a_36_24# 0.00fF
C12747 INVX1_LOC_14/A NOR2X1_LOC_76/A 0.07fF
C12748 NOR2X1_LOC_89/A NOR2X1_LOC_612/Y 0.46fF
C12749 NOR2X1_LOC_139/Y INVX1_LOC_271/A 0.03fF
C12750 NOR2X1_LOC_503/Y INVX1_LOC_10/A 0.07fF
C12751 NOR2X1_LOC_655/B NOR2X1_LOC_360/Y 0.10fF
C12752 INVX1_LOC_54/Y INVX1_LOC_181/Y 0.01fF
C12753 INVX1_LOC_24/A NOR2X1_LOC_720/a_36_216# 0.00fF
C12754 INVX1_LOC_117/Y INVX1_LOC_29/A 0.03fF
C12755 NOR2X1_LOC_218/Y INVX1_LOC_30/A 0.09fF
C12756 INVX1_LOC_307/A INVX1_LOC_263/Y 0.03fF
C12757 INVX1_LOC_314/Y INVX1_LOC_168/A 0.11fF
C12758 NOR2X1_LOC_716/B NOR2X1_LOC_392/B 0.10fF
C12759 NOR2X1_LOC_816/A NAND2X1_LOC_808/A 0.07fF
C12760 NAND2X1_LOC_562/B NAND2X1_LOC_787/B 0.04fF
C12761 INVX1_LOC_224/Y INVX1_LOC_95/Y 0.97fF
C12762 NOR2X1_LOC_124/A INVX1_LOC_57/A 0.03fF
C12763 NOR2X1_LOC_15/Y NAND2X1_LOC_850/A 0.01fF
C12764 INVX1_LOC_13/A INVX1_LOC_40/Y 0.00fF
C12765 INVX1_LOC_244/Y NAND2X1_LOC_11/Y 0.01fF
C12766 INVX1_LOC_136/Y NOR2X1_LOC_631/A 0.07fF
C12767 INVX1_LOC_208/A INVX1_LOC_79/Y 0.00fF
C12768 NAND2X1_LOC_468/B INVX1_LOC_271/A 2.27fF
C12769 NOR2X1_LOC_391/Y INVX1_LOC_306/Y -0.01fF
C12770 INVX1_LOC_18/A INVX1_LOC_53/Y 0.03fF
C12771 INVX1_LOC_48/Y INVX1_LOC_75/A 0.07fF
C12772 INVX1_LOC_89/A NOR2X1_LOC_794/B 0.03fF
C12773 INVX1_LOC_307/A INVX1_LOC_42/A 0.19fF
C12774 INVX1_LOC_58/A NAND2X1_LOC_212/Y 0.02fF
C12775 INVX1_LOC_245/A NOR2X1_LOC_68/A 0.03fF
C12776 INVX1_LOC_88/A NAND2X1_LOC_123/Y 0.18fF
C12777 NOR2X1_LOC_361/B NAND2X1_LOC_842/a_36_24# 0.00fF
C12778 NAND2X1_LOC_563/Y NOR2X1_LOC_84/A 0.01fF
C12779 NOR2X1_LOC_285/Y NOR2X1_LOC_78/A 0.00fF
C12780 NOR2X1_LOC_216/B NOR2X1_LOC_114/Y 0.02fF
C12781 INVX1_LOC_50/A NOR2X1_LOC_280/Y 0.14fF
C12782 NOR2X1_LOC_769/A NAND2X1_LOC_663/a_36_24# 0.00fF
C12783 INVX1_LOC_114/A INVX1_LOC_78/A -0.01fF
C12784 NAND2X1_LOC_841/A INVX1_LOC_71/A 0.03fF
C12785 NAND2X1_LOC_541/a_36_24# NOR2X1_LOC_124/A 0.01fF
C12786 INVX1_LOC_155/Y INVX1_LOC_177/A 1.05fF
C12787 NAND2X1_LOC_783/Y INVX1_LOC_90/A 0.00fF
C12788 INVX1_LOC_279/A INVX1_LOC_72/A 0.07fF
C12789 INVX1_LOC_200/A INVX1_LOC_140/A 0.19fF
C12790 NAND2X1_LOC_360/B INVX1_LOC_33/A 0.01fF
C12791 INVX1_LOC_17/Y VDD 0.50fF
C12792 NOR2X1_LOC_382/Y D_INPUT_0 0.01fF
C12793 INVX1_LOC_119/A INVX1_LOC_221/A 0.03fF
C12794 NOR2X1_LOC_536/A NOR2X1_LOC_301/A 0.38fF
C12795 VDD NOR2X1_LOC_858/A 0.08fF
C12796 NOR2X1_LOC_781/B INVX1_LOC_18/A 0.14fF
C12797 INVX1_LOC_200/Y VDD 0.36fF
C12798 INVX1_LOC_35/A INVX1_LOC_147/Y 0.05fF
C12799 NAND2X1_LOC_866/A NAND2X1_LOC_863/B 0.02fF
C12800 NOR2X1_LOC_78/B INVX1_LOC_63/Y 0.20fF
C12801 INVX1_LOC_58/A INVX1_LOC_14/Y 0.27fF
C12802 NAND2X1_LOC_96/A NOR2X1_LOC_720/A 0.01fF
C12803 NOR2X1_LOC_598/B INVX1_LOC_176/A 0.03fF
C12804 INVX1_LOC_103/A INVX1_LOC_144/A 0.02fF
C12805 INVX1_LOC_307/Y NOR2X1_LOC_334/Y 0.11fF
C12806 INVX1_LOC_223/A INVX1_LOC_313/A 0.03fF
C12807 NAND2X1_LOC_860/A NOR2X1_LOC_558/A 0.03fF
C12808 INVX1_LOC_305/A INVX1_LOC_135/A 0.07fF
C12809 INVX1_LOC_34/A NAND2X1_LOC_350/B 0.01fF
C12810 INVX1_LOC_257/Y INVX1_LOC_259/A 0.21fF
C12811 INVX1_LOC_35/A INVX1_LOC_20/A 0.09fF
C12812 NAND2X1_LOC_571/B VDD 0.02fF
C12813 INVX1_LOC_51/A INVX1_LOC_176/A 0.00fF
C12814 NOR2X1_LOC_186/Y NAND2X1_LOC_642/Y 0.07fF
C12815 NOR2X1_LOC_577/Y INVX1_LOC_16/A 0.14fF
C12816 INVX1_LOC_30/A INPUT_1 0.03fF
C12817 INVX1_LOC_27/A NOR2X1_LOC_139/Y 0.06fF
C12818 INVX1_LOC_89/A NOR2X1_LOC_384/Y 0.13fF
C12819 NOR2X1_LOC_67/a_36_216# NOR2X1_LOC_721/B 0.00fF
C12820 NOR2X1_LOC_360/Y NOR2X1_LOC_99/B 0.07fF
C12821 NAND2X1_LOC_812/A NAND2X1_LOC_863/B 0.05fF
C12822 NAND2X1_LOC_740/Y INVX1_LOC_11/Y 0.37fF
C12823 INVX1_LOC_163/Y INVX1_LOC_167/A 0.02fF
C12824 INVX1_LOC_34/A INVX1_LOC_208/A 0.08fF
C12825 INVX1_LOC_182/Y NOR2X1_LOC_348/a_36_216# 0.00fF
C12826 INVX1_LOC_2/A NAND2X1_LOC_722/A 0.01fF
C12827 NAND2X1_LOC_529/a_36_24# NOR2X1_LOC_721/Y 0.00fF
C12828 NOR2X1_LOC_357/Y NOR2X1_LOC_665/Y 0.27fF
C12829 VDD INVX1_LOC_292/Y 0.59fF
C12830 INVX1_LOC_78/A INVX1_LOC_307/A 0.07fF
C12831 INVX1_LOC_38/A NOR2X1_LOC_654/A 0.05fF
C12832 NAND2X1_LOC_500/Y NAND2X1_LOC_560/A 0.01fF
C12833 INVX1_LOC_10/A NOR2X1_LOC_152/Y 0.10fF
C12834 NOR2X1_LOC_68/A NOR2X1_LOC_788/B 0.11fF
C12835 NOR2X1_LOC_160/B INPUT_0 0.19fF
C12836 NOR2X1_LOC_284/B NOR2X1_LOC_168/B 0.01fF
C12837 INVX1_LOC_1/Y INVX1_LOC_8/A 0.00fF
C12838 NAND2X1_LOC_573/Y NAND2X1_LOC_642/Y 0.07fF
C12839 INVX1_LOC_27/A NAND2X1_LOC_468/B 0.03fF
C12840 NOR2X1_LOC_550/B NOR2X1_LOC_565/B 0.02fF
C12841 INVX1_LOC_78/A NOR2X1_LOC_445/B 0.07fF
C12842 NOR2X1_LOC_380/A NAND2X1_LOC_863/Y 0.02fF
C12843 INVX1_LOC_298/A INVX1_LOC_37/A 0.00fF
C12844 INVX1_LOC_182/Y INVX1_LOC_72/A 0.03fF
C12845 INVX1_LOC_10/Y NOR2X1_LOC_678/A 0.54fF
C12846 NOR2X1_LOC_84/Y INVX1_LOC_25/Y 0.06fF
C12847 NAND2X1_LOC_141/A INVX1_LOC_316/Y 0.02fF
C12848 INVX1_LOC_57/Y NOR2X1_LOC_322/Y 0.18fF
C12849 INVX1_LOC_77/A NAND2X1_LOC_45/Y 0.15fF
C12850 NOR2X1_LOC_617/Y NAND2X1_LOC_624/A 0.00fF
C12851 INVX1_LOC_38/A INVX1_LOC_58/Y 0.07fF
C12852 INVX1_LOC_12/A INVX1_LOC_42/A 0.17fF
C12853 NOR2X1_LOC_328/Y NOR2X1_LOC_504/Y 0.08fF
C12854 INVX1_LOC_226/Y NOR2X1_LOC_721/A 0.05fF
C12855 INVX1_LOC_90/A NOR2X1_LOC_419/Y 0.06fF
C12856 NOR2X1_LOC_455/Y INVX1_LOC_9/A 0.01fF
C12857 INVX1_LOC_83/A INVX1_LOC_63/Y 0.03fF
C12858 NOR2X1_LOC_717/B NOR2X1_LOC_147/B 0.01fF
C12859 NAND2X1_LOC_787/A INVX1_LOC_118/A 0.04fF
C12860 NAND2X1_LOC_717/Y INVX1_LOC_22/A 0.07fF
C12861 D_INPUT_6 INVX1_LOC_37/A 0.49fF
C12862 NOR2X1_LOC_173/Y INVX1_LOC_37/A 0.03fF
C12863 NOR2X1_LOC_634/Y NOR2X1_LOC_729/A 0.00fF
C12864 INVX1_LOC_90/A NOR2X1_LOC_716/B 0.20fF
C12865 NAND2X1_LOC_863/B NOR2X1_LOC_505/Y 0.01fF
C12866 INVX1_LOC_223/A INVX1_LOC_6/A 0.03fF
C12867 NOR2X1_LOC_103/Y INVX1_LOC_95/Y 0.19fF
C12868 NOR2X1_LOC_227/B VDD -0.00fF
C12869 INVX1_LOC_50/A NOR2X1_LOC_197/B 0.00fF
C12870 NAND2X1_LOC_67/Y INVX1_LOC_76/A 0.03fF
C12871 NAND2X1_LOC_810/B INVX1_LOC_296/Y 0.05fF
C12872 NOR2X1_LOC_245/a_36_216# NOR2X1_LOC_309/Y 0.01fF
C12873 INVX1_LOC_28/A NOR2X1_LOC_577/Y 0.47fF
C12874 NOR2X1_LOC_113/B INVX1_LOC_18/A 0.03fF
C12875 NAND2X1_LOC_493/Y VDD 0.09fF
C12876 NOR2X1_LOC_443/Y NOR2X1_LOC_688/a_36_216# 0.00fF
C12877 INVX1_LOC_113/Y NOR2X1_LOC_302/Y 0.04fF
C12878 INVX1_LOC_163/A INVX1_LOC_194/Y 0.03fF
C12879 NAND2X1_LOC_678/a_36_24# NOR2X1_LOC_88/Y 0.01fF
C12880 NOR2X1_LOC_441/Y NOR2X1_LOC_269/Y 0.08fF
C12881 NAND2X1_LOC_218/B NAND2X1_LOC_126/a_36_24# -0.02fF
C12882 NAND2X1_LOC_217/a_36_24# INVX1_LOC_75/A 0.00fF
C12883 NOR2X1_LOC_38/a_36_216# INVX1_LOC_3/Y 0.00fF
C12884 NOR2X1_LOC_68/A NOR2X1_LOC_147/A 0.05fF
C12885 NOR2X1_LOC_38/B INVX1_LOC_284/A 0.62fF
C12886 NOR2X1_LOC_34/B INVX1_LOC_9/A 0.01fF
C12887 NOR2X1_LOC_273/Y INVX1_LOC_311/A 0.02fF
C12888 INVX1_LOC_16/A INVX1_LOC_22/A 0.93fF
C12889 NOR2X1_LOC_789/A INVX1_LOC_232/A 0.03fF
C12890 NOR2X1_LOC_561/Y NOR2X1_LOC_131/a_36_216# 0.01fF
C12891 NOR2X1_LOC_214/B INVX1_LOC_266/Y 0.01fF
C12892 NOR2X1_LOC_791/Y INVX1_LOC_118/A 0.02fF
C12893 INVX1_LOC_78/A INVX1_LOC_12/A 4.39fF
C12894 NOR2X1_LOC_246/A NAND2X1_LOC_342/Y 0.04fF
C12895 NOR2X1_LOC_460/B INVX1_LOC_75/A 0.02fF
C12896 NOR2X1_LOC_773/Y NAND2X1_LOC_808/A 0.01fF
C12897 INVX1_LOC_5/A INVX1_LOC_92/A 0.17fF
C12898 INVX1_LOC_294/A INVX1_LOC_29/Y 0.00fF
C12899 INVX1_LOC_45/A INVX1_LOC_95/Y 0.03fF
C12900 NOR2X1_LOC_151/Y NOR2X1_LOC_147/B 0.10fF
C12901 INVX1_LOC_311/A NOR2X1_LOC_550/B 0.10fF
C12902 INVX1_LOC_246/A NAND2X1_LOC_453/A 0.04fF
C12903 INVX1_LOC_17/A NAND2X1_LOC_639/A 0.07fF
C12904 INVX1_LOC_304/Y INVX1_LOC_140/A 0.85fF
C12905 INVX1_LOC_21/A INVX1_LOC_75/Y 0.13fF
C12906 INVX1_LOC_17/A NOR2X1_LOC_536/A 0.33fF
C12907 NOR2X1_LOC_81/a_36_216# NOR2X1_LOC_78/A 0.00fF
C12908 NOR2X1_LOC_65/B INVX1_LOC_12/A 0.03fF
C12909 INVX1_LOC_178/A INVX1_LOC_92/A 1.37fF
C12910 INVX1_LOC_285/Y INVX1_LOC_155/Y 0.03fF
C12911 INVX1_LOC_75/A NOR2X1_LOC_84/Y 0.07fF
C12912 NOR2X1_LOC_60/a_36_216# NAND2X1_LOC_660/Y 0.03fF
C12913 INVX1_LOC_303/A NOR2X1_LOC_557/A 0.03fF
C12914 NAND2X1_LOC_286/B NAND2X1_LOC_807/a_36_24# 0.00fF
C12915 INVX1_LOC_311/A INVX1_LOC_249/Y 0.01fF
C12916 INVX1_LOC_162/Y INVX1_LOC_6/A 0.13fF
C12917 NAND2X1_LOC_856/A NOR2X1_LOC_305/Y 0.02fF
C12918 INVX1_LOC_18/A NOR2X1_LOC_585/Y 0.11fF
C12919 INVX1_LOC_27/A NAND2X1_LOC_141/Y 1.37fF
C12920 NAND2X1_LOC_656/Y NOR2X1_LOC_366/Y 0.03fF
C12921 NOR2X1_LOC_45/B NAND2X1_LOC_631/a_36_24# 0.01fF
C12922 INVX1_LOC_250/A VDD 0.12fF
C12923 NOR2X1_LOC_860/B NOR2X1_LOC_346/Y 0.01fF
C12924 INVX1_LOC_85/A INVX1_LOC_6/A 0.00fF
C12925 INVX1_LOC_95/Y INVX1_LOC_71/A 0.20fF
C12926 NOR2X1_LOC_392/B NOR2X1_LOC_392/a_36_216# 0.00fF
C12927 NAND2X1_LOC_721/B NAND2X1_LOC_721/A 0.02fF
C12928 NAND2X1_LOC_363/B NAND2X1_LOC_63/Y 0.10fF
C12929 NOR2X1_LOC_598/B NOR2X1_LOC_340/A 0.07fF
C12930 NOR2X1_LOC_445/Y INVX1_LOC_91/A 0.04fF
C12931 INVX1_LOC_28/A INVX1_LOC_22/A 0.36fF
C12932 NOR2X1_LOC_602/a_36_216# NOR2X1_LOC_111/A 0.01fF
C12933 NOR2X1_LOC_315/Y NOR2X1_LOC_368/a_36_216# 0.00fF
C12934 NOR2X1_LOC_142/Y NOR2X1_LOC_269/Y 0.26fF
C12935 INVX1_LOC_290/Y INVX1_LOC_23/A 0.07fF
C12936 INVX1_LOC_17/A NAND2X1_LOC_93/B 0.03fF
C12937 INVX1_LOC_136/A NAND2X1_LOC_804/Y 0.03fF
C12938 NOR2X1_LOC_717/B INVX1_LOC_97/A 0.47fF
C12939 INVX1_LOC_279/A INVX1_LOC_313/Y 0.01fF
C12940 NOR2X1_LOC_355/A NOR2X1_LOC_106/A 0.10fF
C12941 NOR2X1_LOC_690/A NAND2X1_LOC_623/B 0.08fF
C12942 NAND2X1_LOC_555/Y NAND2X1_LOC_659/a_36_24# 0.00fF
C12943 INVX1_LOC_272/Y NAND2X1_LOC_802/Y 0.54fF
C12944 NOR2X1_LOC_299/Y INVX1_LOC_173/Y 4.95fF
C12945 NAND2X1_LOC_510/a_36_24# NOR2X1_LOC_349/A 0.00fF
C12946 NAND2X1_LOC_295/a_36_24# NOR2X1_LOC_416/A 0.00fF
C12947 INVX1_LOC_35/A NOR2X1_LOC_128/A 0.01fF
C12948 INVX1_LOC_64/A NOR2X1_LOC_671/a_36_216# 0.00fF
C12949 INVX1_LOC_103/A NOR2X1_LOC_155/A 0.11fF
C12950 NOR2X1_LOC_717/B INVX1_LOC_90/A 0.03fF
C12951 NOR2X1_LOC_741/A INVX1_LOC_266/Y 0.02fF
C12952 INVX1_LOC_141/A INVX1_LOC_54/A 0.02fF
C12953 INVX1_LOC_116/A VDD 0.12fF
C12954 NOR2X1_LOC_410/Y NAND2X1_LOC_96/A 0.03fF
C12955 NOR2X1_LOC_67/A NOR2X1_LOC_86/a_36_216# 0.00fF
C12956 INVX1_LOC_208/A INPUT_0 0.07fF
C12957 INVX1_LOC_225/A NAND2X1_LOC_642/Y 0.03fF
C12958 NAND2X1_LOC_555/Y NOR2X1_LOC_655/Y 0.09fF
C12959 NOR2X1_LOC_471/Y NAND2X1_LOC_93/B 0.07fF
C12960 INVX1_LOC_32/A NOR2X1_LOC_414/Y 0.28fF
C12961 INVX1_LOC_78/A NOR2X1_LOC_686/A 0.10fF
C12962 INVX1_LOC_155/Y NOR2X1_LOC_137/B 0.09fF
C12963 NOR2X1_LOC_816/A INVX1_LOC_92/A 0.08fF
C12964 NAND2X1_LOC_392/A NOR2X1_LOC_74/A 0.00fF
C12965 NOR2X1_LOC_168/B INVX1_LOC_186/A 0.03fF
C12966 NOR2X1_LOC_516/B INPUT_0 0.11fF
C12967 NOR2X1_LOC_495/Y VDD 0.41fF
C12968 INVX1_LOC_102/A NOR2X1_LOC_109/Y 0.08fF
C12969 INVX1_LOC_30/A INVX1_LOC_118/A 0.35fF
C12970 NAND2X1_LOC_222/B NOR2X1_LOC_673/A 0.04fF
C12971 NOR2X1_LOC_826/Y INVX1_LOC_3/Y 0.08fF
C12972 NOR2X1_LOC_637/Y INVX1_LOC_77/Y 0.01fF
C12973 NOR2X1_LOC_334/Y NOR2X1_LOC_809/A 0.00fF
C12974 NOR2X1_LOC_15/Y NOR2X1_LOC_662/A 0.11fF
C12975 NOR2X1_LOC_130/A NAND2X1_LOC_652/Y 0.02fF
C12976 INVX1_LOC_140/A NAND2X1_LOC_808/A 0.10fF
C12977 NAND2X1_LOC_63/Y NAND2X1_LOC_63/a_36_24# 0.02fF
C12978 INVX1_LOC_21/A NAND2X1_LOC_74/B 0.18fF
C12979 NAND2X1_LOC_361/Y VDD 0.01fF
C12980 INVX1_LOC_270/Y INVX1_LOC_94/Y 0.04fF
C12981 NOR2X1_LOC_775/Y INVX1_LOC_132/Y 0.15fF
C12982 INVX1_LOC_254/A INVX1_LOC_117/A 0.02fF
C12983 INVX1_LOC_57/A INVX1_LOC_273/A 0.03fF
C12984 INVX1_LOC_34/A NAND2X1_LOC_211/Y 0.00fF
C12985 NOR2X1_LOC_334/Y INVX1_LOC_29/Y 0.08fF
C12986 NOR2X1_LOC_751/Y NOR2X1_LOC_641/Y 0.02fF
C12987 INVX1_LOC_63/Y INVX1_LOC_46/A 0.03fF
C12988 INVX1_LOC_17/A NOR2X1_LOC_661/A 0.03fF
C12989 NAND2X1_LOC_662/Y INVX1_LOC_6/A 0.11fF
C12990 INVX1_LOC_26/Y NOR2X1_LOC_621/A 0.01fF
C12991 NOR2X1_LOC_348/B NOR2X1_LOC_35/Y 0.02fF
C12992 NOR2X1_LOC_458/a_36_216# INVX1_LOC_271/Y -0.01fF
C12993 D_INPUT_1 NOR2X1_LOC_465/Y 0.04fF
C12994 INVX1_LOC_35/A INVX1_LOC_4/A 0.07fF
C12995 INVX1_LOC_36/A INVX1_LOC_70/A 0.04fF
C12996 NOR2X1_LOC_367/B INVX1_LOC_76/A 0.02fF
C12997 INVX1_LOC_269/A INVX1_LOC_19/A 0.16fF
C12998 VDD NAND2X1_LOC_799/Y 0.07fF
C12999 INVX1_LOC_219/Y VDD 0.21fF
C13000 INVX1_LOC_182/Y INVX1_LOC_313/Y 0.98fF
C13001 NOR2X1_LOC_419/Y INVX1_LOC_38/A 0.03fF
C13002 INVX1_LOC_90/A NOR2X1_LOC_151/Y 0.03fF
C13003 INVX1_LOC_113/Y INVX1_LOC_114/A 0.01fF
C13004 INVX1_LOC_286/A INVX1_LOC_164/A 0.18fF
C13005 NAND2X1_LOC_348/A NOR2X1_LOC_130/Y -0.00fF
C13006 NAND2X1_LOC_555/Y NOR2X1_LOC_649/B 2.76fF
C13007 INVX1_LOC_27/A NAND2X1_LOC_213/a_36_24# 0.00fF
C13008 NOR2X1_LOC_564/Y NOR2X1_LOC_703/A 0.00fF
C13009 NAND2X1_LOC_555/Y INVX1_LOC_3/A 1.13fF
C13010 INVX1_LOC_299/A INVX1_LOC_69/A 0.01fF
C13011 NOR2X1_LOC_716/B INVX1_LOC_38/A 0.08fF
C13012 INVX1_LOC_89/A NOR2X1_LOC_188/A 0.05fF
C13013 INVX1_LOC_14/A NOR2X1_LOC_14/a_36_216# 0.03fF
C13014 NOR2X1_LOC_346/B NOR2X1_LOC_35/Y 0.01fF
C13015 NAND2X1_LOC_231/Y NAND2X1_LOC_211/Y 0.44fF
C13016 INVX1_LOC_223/A NOR2X1_LOC_117/Y 0.01fF
C13017 INVX1_LOC_89/A NOR2X1_LOC_548/B 0.01fF
C13018 NOR2X1_LOC_710/A NAND2X1_LOC_782/B 0.03fF
C13019 NOR2X1_LOC_82/A INVX1_LOC_29/A 0.07fF
C13020 NOR2X1_LOC_45/Y NOR2X1_LOC_48/Y 0.00fF
C13021 NOR2X1_LOC_503/Y INVX1_LOC_12/A 0.03fF
C13022 INVX1_LOC_28/A INVX1_LOC_100/A 0.09fF
C13023 INVX1_LOC_22/A NOR2X1_LOC_35/Y 0.05fF
C13024 INVX1_LOC_200/A INVX1_LOC_42/A 0.17fF
C13025 INVX1_LOC_120/A NOR2X1_LOC_845/A 0.14fF
C13026 NOR2X1_LOC_719/A INVX1_LOC_76/A 0.00fF
C13027 NOR2X1_LOC_68/A NAND2X1_LOC_42/a_36_24# 0.00fF
C13028 NAND2X1_LOC_319/A NOR2X1_LOC_56/Y 0.01fF
C13029 NAND2X1_LOC_338/B NOR2X1_LOC_98/B 0.04fF
C13030 NAND2X1_LOC_842/B INVX1_LOC_100/Y 0.01fF
C13031 INVX1_LOC_58/A NOR2X1_LOC_826/Y 0.04fF
C13032 INVX1_LOC_89/A NOR2X1_LOC_43/Y 0.13fF
C13033 NOR2X1_LOC_564/a_36_216# NOR2X1_LOC_564/Y 0.02fF
C13034 INVX1_LOC_25/A NOR2X1_LOC_392/Y 0.29fF
C13035 NOR2X1_LOC_828/Y INVX1_LOC_53/A 0.13fF
C13036 INVX1_LOC_67/A NOR2X1_LOC_155/A 0.03fF
C13037 NAND2X1_LOC_36/A INVX1_LOC_29/A 0.00fF
C13038 INVX1_LOC_30/A NAND2X1_LOC_63/Y 0.49fF
C13039 NOR2X1_LOC_561/Y INVX1_LOC_76/A 0.17fF
C13040 NOR2X1_LOC_791/B NAND2X1_LOC_773/B 0.08fF
C13041 INVX1_LOC_95/Y NOR2X1_LOC_123/B 0.07fF
C13042 NAND2X1_LOC_722/A INVX1_LOC_118/A 0.07fF
C13043 INVX1_LOC_7/A INVX1_LOC_76/A 0.09fF
C13044 INVX1_LOC_249/A NOR2X1_LOC_66/Y 0.03fF
C13045 NOR2X1_LOC_377/Y INVX1_LOC_92/A 0.06fF
C13046 NAND2X1_LOC_319/A VDD -0.00fF
C13047 NAND2X1_LOC_364/A INVX1_LOC_125/A 0.02fF
C13048 NOR2X1_LOC_32/B INVX1_LOC_233/Y 0.00fF
C13049 NAND2X1_LOC_453/a_36_24# NAND2X1_LOC_798/B 0.00fF
C13050 INVX1_LOC_35/A INVX1_LOC_64/A 0.20fF
C13051 NAND2X1_LOC_778/Y INVX1_LOC_57/A 0.27fF
C13052 INVX1_LOC_212/A NOR2X1_LOC_509/A 0.00fF
C13053 INVX1_LOC_5/A INVX1_LOC_53/A 2.62fF
C13054 NOR2X1_LOC_384/Y NOR2X1_LOC_490/a_36_216# 0.00fF
C13055 INVX1_LOC_217/A INVX1_LOC_42/A 0.13fF
C13056 NAND2X1_LOC_803/B NOR2X1_LOC_158/Y 0.02fF
C13057 NOR2X1_LOC_335/B INVX1_LOC_91/A 0.52fF
C13058 INVX1_LOC_95/Y INVX1_LOC_102/Y 0.13fF
C13059 NOR2X1_LOC_773/Y INVX1_LOC_92/A 0.07fF
C13060 NOR2X1_LOC_620/B NOR2X1_LOC_862/B 0.04fF
C13061 INVX1_LOC_178/A INVX1_LOC_53/A 0.05fF
C13062 NOR2X1_LOC_454/Y INVX1_LOC_23/A 0.08fF
C13063 NOR2X1_LOC_667/Y INVX1_LOC_94/Y 0.00fF
C13064 NAND2X1_LOC_861/Y NOR2X1_LOC_301/a_36_216# 0.00fF
C13065 NAND2X1_LOC_598/a_36_24# NOR2X1_LOC_409/B 0.00fF
C13066 NOR2X1_LOC_15/Y INVX1_LOC_57/A 0.24fF
C13067 NOR2X1_LOC_152/Y INVX1_LOC_12/A 0.07fF
C13068 NOR2X1_LOC_45/B NAND2X1_LOC_814/a_36_24# 0.01fF
C13069 INVX1_LOC_186/A INVX1_LOC_78/Y 0.03fF
C13070 NAND2X1_LOC_654/B VDD 0.22fF
C13071 NOR2X1_LOC_717/B INVX1_LOC_38/A 0.03fF
C13072 INVX1_LOC_58/A NAND2X1_LOC_303/Y 0.11fF
C13073 INVX1_LOC_113/Y INVX1_LOC_12/A 0.06fF
C13074 NAND2X1_LOC_354/B INVX1_LOC_264/A 0.03fF
C13075 INVX1_LOC_148/A INVX1_LOC_37/A 0.03fF
C13076 INVX1_LOC_88/A INVX1_LOC_271/A 1.81fF
C13077 INVX1_LOC_223/A NAND2X1_LOC_646/a_36_24# 0.00fF
C13078 NOR2X1_LOC_403/a_36_216# NAND2X1_LOC_254/Y 0.01fF
C13079 NAND2X1_LOC_139/A NAND2X1_LOC_82/Y 0.02fF
C13080 INVX1_LOC_72/A NOR2X1_LOC_38/B 0.17fF
C13081 INVX1_LOC_230/Y INVX1_LOC_16/Y 0.01fF
C13082 INVX1_LOC_146/A NOR2X1_LOC_447/B 0.01fF
C13083 NAND2X1_LOC_35/Y NOR2X1_LOC_233/a_36_216# 0.01fF
C13084 NAND2X1_LOC_41/Y INVX1_LOC_108/A 0.13fF
C13085 INVX1_LOC_45/A INVX1_LOC_271/Y 0.07fF
C13086 NOR2X1_LOC_790/B INVX1_LOC_24/Y 0.05fF
C13087 NOR2X1_LOC_409/Y VDD 0.31fF
C13088 INVX1_LOC_1/A NOR2X1_LOC_392/Y 0.07fF
C13089 NAND2X1_LOC_787/B INVX1_LOC_42/A 0.07fF
C13090 NAND2X1_LOC_45/Y INVX1_LOC_9/A 0.09fF
C13091 NOR2X1_LOC_598/B INVX1_LOC_103/A 0.10fF
C13092 INVX1_LOC_27/A INVX1_LOC_13/Y 0.14fF
C13093 NOR2X1_LOC_328/Y NOR2X1_LOC_697/Y 0.02fF
C13094 INVX1_LOC_217/A INVX1_LOC_78/A 0.01fF
C13095 INVX1_LOC_13/Y NOR2X1_LOC_824/A 0.00fF
C13096 INVX1_LOC_10/A NAND2X1_LOC_802/Y 0.07fF
C13097 INVX1_LOC_230/Y NAND2X1_LOC_205/A 0.05fF
C13098 NOR2X1_LOC_781/Y NOR2X1_LOC_158/B 0.02fF
C13099 NAND2X1_LOC_337/B INVX1_LOC_53/A 0.07fF
C13100 NOR2X1_LOC_309/Y INVX1_LOC_102/A 0.10fF
C13101 NOR2X1_LOC_100/A INVX1_LOC_29/A 0.00fF
C13102 INVX1_LOC_50/A INVX1_LOC_286/Y 0.04fF
C13103 NOR2X1_LOC_816/A INVX1_LOC_53/A 0.07fF
C13104 INVX1_LOC_223/A INVX1_LOC_28/Y 0.02fF
C13105 INVX1_LOC_16/A NAND2X1_LOC_476/Y 0.01fF
C13106 INVX1_LOC_277/A NOR2X1_LOC_748/A 0.11fF
C13107 INVX1_LOC_304/Y INVX1_LOC_42/A 0.01fF
C13108 NOR2X1_LOC_690/A INVX1_LOC_3/Y 0.02fF
C13109 NAND2X1_LOC_571/Y INVX1_LOC_234/Y 0.09fF
C13110 INVX1_LOC_71/A INVX1_LOC_271/Y 0.07fF
C13111 INVX1_LOC_223/A INVX1_LOC_270/A 0.01fF
C13112 INVX1_LOC_13/A NOR2X1_LOC_814/A 0.08fF
C13113 NOR2X1_LOC_151/Y INVX1_LOC_38/A 0.12fF
C13114 NOR2X1_LOC_524/Y INVX1_LOC_270/Y 0.12fF
C13115 NOR2X1_LOC_748/Y INVX1_LOC_63/A 0.03fF
C13116 NOR2X1_LOC_9/Y INVX1_LOC_129/Y 0.00fF
C13117 NOR2X1_LOC_413/Y INVX1_LOC_3/Y 0.01fF
C13118 INVX1_LOC_16/A INVX1_LOC_186/Y 0.15fF
C13119 NOR2X1_LOC_419/Y NAND2X1_LOC_223/A 0.07fF
C13120 NAND2X1_LOC_214/Y NAND2X1_LOC_473/A 0.03fF
C13121 NOR2X1_LOC_433/A NOR2X1_LOC_409/B 0.02fF
C13122 NOR2X1_LOC_356/A NOR2X1_LOC_809/B 0.03fF
C13123 INVX1_LOC_27/A INVX1_LOC_88/A 0.03fF
C13124 VDD INVX1_LOC_159/Y 0.00fF
C13125 NOR2X1_LOC_324/A NOR2X1_LOC_324/B 0.03fF
C13126 NOR2X1_LOC_457/B NOR2X1_LOC_383/B 0.07fF
C13127 NOR2X1_LOC_253/a_36_216# INVX1_LOC_217/A 0.01fF
C13128 INVX1_LOC_269/A NOR2X1_LOC_474/a_36_216# 0.00fF
C13129 NOR2X1_LOC_246/A INVX1_LOC_285/A 0.01fF
C13130 NOR2X1_LOC_444/a_36_216# NAND2X1_LOC_364/A 0.01fF
C13131 NOR2X1_LOC_152/Y NOR2X1_LOC_686/A 0.02fF
C13132 NOR2X1_LOC_15/Y NOR2X1_LOC_475/A 0.01fF
C13133 INVX1_LOC_22/A INVX1_LOC_109/A 0.01fF
C13134 NOR2X1_LOC_720/B INVX1_LOC_4/Y 0.01fF
C13135 NOR2X1_LOC_824/Y INVX1_LOC_76/A 0.03fF
C13136 NOR2X1_LOC_15/Y NOR2X1_LOC_666/Y 0.35fF
C13137 INVX1_LOC_316/Y NOR2X1_LOC_672/a_36_216# 0.00fF
C13138 NOR2X1_LOC_313/Y INVX1_LOC_54/A 0.05fF
C13139 INVX1_LOC_8/A INVX1_LOC_87/A 2.43fF
C13140 NOR2X1_LOC_201/A INVX1_LOC_77/A 0.06fF
C13141 NOR2X1_LOC_174/B NOR2X1_LOC_814/A 0.01fF
C13142 NAND2X1_LOC_578/B INVX1_LOC_15/A 0.12fF
C13143 NOR2X1_LOC_802/A NAND2X1_LOC_615/a_36_24# 0.00fF
C13144 NAND2X1_LOC_656/A INVX1_LOC_129/A 0.54fF
C13145 NOR2X1_LOC_19/B NAND2X1_LOC_141/Y 0.32fF
C13146 NAND2X1_LOC_773/Y NOR2X1_LOC_103/Y 0.10fF
C13147 NOR2X1_LOC_316/Y NOR2X1_LOC_80/Y 0.02fF
C13148 NOR2X1_LOC_612/a_36_216# INVX1_LOC_47/Y 0.01fF
C13149 NOR2X1_LOC_537/Y NOR2X1_LOC_38/B 4.58fF
C13150 NAND2X1_LOC_338/B NOR2X1_LOC_38/B 0.19fF
C13151 NOR2X1_LOC_604/Y NOR2X1_LOC_596/A 0.01fF
C13152 NAND2X1_LOC_357/B NOR2X1_LOC_281/a_36_216# 0.00fF
C13153 NOR2X1_LOC_562/A NOR2X1_LOC_357/Y 0.01fF
C13154 NAND2X1_LOC_796/B INVX1_LOC_141/Y 0.57fF
C13155 INVX1_LOC_77/A INVX1_LOC_23/A 0.41fF
C13156 NOR2X1_LOC_318/B INVX1_LOC_118/Y 0.04fF
C13157 INVX1_LOC_269/A INVX1_LOC_161/Y 0.01fF
C13158 NOR2X1_LOC_97/A NOR2X1_LOC_865/Y 0.02fF
C13159 NAND2X1_LOC_565/a_36_24# INVX1_LOC_61/A 0.01fF
C13160 NAND2X1_LOC_642/Y NOR2X1_LOC_271/Y 0.01fF
C13161 INVX1_LOC_96/A INVX1_LOC_274/A 0.20fF
C13162 INVX1_LOC_17/A INVX1_LOC_256/A 0.19fF
C13163 INVX1_LOC_27/A NOR2X1_LOC_500/B 0.03fF
C13164 NOR2X1_LOC_97/A NOR2X1_LOC_243/B 0.02fF
C13165 NOR2X1_LOC_121/A INVX1_LOC_4/A 0.03fF
C13166 INVX1_LOC_214/Y INVX1_LOC_78/A 0.52fF
C13167 NAND2X1_LOC_808/A INVX1_LOC_42/A 0.11fF
C13168 INVX1_LOC_21/A INVX1_LOC_136/A 6.93fF
C13169 INVX1_LOC_58/A NOR2X1_LOC_690/A 0.04fF
C13170 NOR2X1_LOC_309/Y NOR2X1_LOC_280/a_36_216# 0.01fF
C13171 INVX1_LOC_165/Y NOR2X1_LOC_394/Y 0.05fF
C13172 NOR2X1_LOC_689/Y INVX1_LOC_240/A 0.02fF
C13173 NOR2X1_LOC_655/B INVX1_LOC_26/A 0.03fF
C13174 NOR2X1_LOC_187/a_36_216# INVX1_LOC_92/A 0.00fF
C13175 NAND2X1_LOC_190/Y NOR2X1_LOC_348/a_36_216# 0.00fF
C13176 INVX1_LOC_33/A INVX1_LOC_58/Y 0.04fF
C13177 INVX1_LOC_58/A NOR2X1_LOC_194/Y 0.02fF
C13178 NAND2X1_LOC_76/a_36_24# INVX1_LOC_11/A 0.00fF
C13179 NOR2X1_LOC_562/B INVX1_LOC_179/A 0.18fF
C13180 NAND2X1_LOC_149/Y INVX1_LOC_18/A 0.25fF
C13181 NOR2X1_LOC_88/Y INVX1_LOC_91/A 0.07fF
C13182 NOR2X1_LOC_363/Y NAND2X1_LOC_472/Y 0.29fF
C13183 NOR2X1_LOC_468/Y INVX1_LOC_72/A 0.15fF
C13184 INVX1_LOC_101/A NOR2X1_LOC_334/Y 0.02fF
C13185 NOR2X1_LOC_593/Y NAND2X1_LOC_406/a_36_24# 0.00fF
C13186 NOR2X1_LOC_792/B INVX1_LOC_308/A 0.03fF
C13187 INVX1_LOC_15/Y INVX1_LOC_57/A 0.03fF
C13188 NOR2X1_LOC_647/B NAND2X1_LOC_555/Y 0.06fF
C13189 NAND2X1_LOC_198/B NOR2X1_LOC_321/Y 0.10fF
C13190 NOR2X1_LOC_604/a_36_216# NOR2X1_LOC_423/Y 0.01fF
C13191 NOR2X1_LOC_141/a_36_216# NOR2X1_LOC_155/A 0.00fF
C13192 NOR2X1_LOC_643/A NOR2X1_LOC_554/B 0.01fF
C13193 NAND2X1_LOC_28/a_36_24# INVX1_LOC_32/A 0.00fF
C13194 INVX1_LOC_303/A INVX1_LOC_27/A 0.04fF
C13195 NAND2X1_LOC_725/A INVX1_LOC_240/A 0.53fF
C13196 INVX1_LOC_75/A INVX1_LOC_114/Y 0.03fF
C13197 INVX1_LOC_84/A INVX1_LOC_91/A 0.14fF
C13198 NAND2X1_LOC_840/B INVX1_LOC_57/A 0.13fF
C13199 INPUT_0 NAND2X1_LOC_207/B 0.00fF
C13200 INVX1_LOC_40/Y INPUT_3 0.01fF
C13201 INVX1_LOC_177/A INVX1_LOC_292/Y 0.08fF
C13202 NAND2X1_LOC_571/B INVX1_LOC_280/Y 0.08fF
C13203 NOR2X1_LOC_202/a_36_216# NOR2X1_LOC_759/Y 0.00fF
C13204 NAND2X1_LOC_577/A NOR2X1_LOC_514/A 0.09fF
C13205 NOR2X1_LOC_92/Y NOR2X1_LOC_387/Y 0.01fF
C13206 NOR2X1_LOC_773/Y INVX1_LOC_53/A 0.01fF
C13207 INVX1_LOC_25/A INVX1_LOC_25/Y 0.11fF
C13208 D_INPUT_0 NOR2X1_LOC_278/Y 0.01fF
C13209 INVX1_LOC_35/A NAND2X1_LOC_850/Y 0.07fF
C13210 NOR2X1_LOC_389/A INVX1_LOC_72/A 0.10fF
C13211 NOR2X1_LOC_687/Y INVX1_LOC_23/A 0.06fF
C13212 INVX1_LOC_37/A NAND2X1_LOC_798/B 0.02fF
C13213 INVX1_LOC_13/Y NAND2X1_LOC_471/a_36_24# 0.01fF
C13214 INVX1_LOC_269/A NAND2X1_LOC_119/a_36_24# 0.07fF
C13215 NOR2X1_LOC_160/B INVX1_LOC_72/Y 0.02fF
C13216 NOR2X1_LOC_99/B INVX1_LOC_26/A 0.04fF
C13217 NOR2X1_LOC_82/A INVX1_LOC_228/A 0.02fF
C13218 NAND2X1_LOC_579/A INVX1_LOC_207/A 0.07fF
C13219 NOR2X1_LOC_848/a_36_216# NOR2X1_LOC_87/B 0.00fF
C13220 NAND2X1_LOC_199/B INVX1_LOC_72/A 0.03fF
C13221 INVX1_LOC_75/A NOR2X1_LOC_467/A 0.22fF
C13222 NOR2X1_LOC_798/A NOR2X1_LOC_175/A 0.04fF
C13223 NOR2X1_LOC_706/B NAND2X1_LOC_425/Y 0.01fF
C13224 INVX1_LOC_5/A NOR2X1_LOC_78/B 0.71fF
C13225 NOR2X1_LOC_454/Y NOR2X1_LOC_75/a_36_216# 0.01fF
C13226 NOR2X1_LOC_405/A INVX1_LOC_125/A 0.08fF
C13227 NOR2X1_LOC_534/a_36_216# INVX1_LOC_4/A 0.00fF
C13228 NOR2X1_LOC_92/Y NAND2X1_LOC_357/B 0.07fF
C13229 INVX1_LOC_179/A INVX1_LOC_281/Y 0.01fF
C13230 NOR2X1_LOC_778/A NOR2X1_LOC_778/Y 0.04fF
C13231 INVX1_LOC_119/A NAND2X1_LOC_326/A 0.01fF
C13232 NOR2X1_LOC_825/Y INVX1_LOC_203/A 0.10fF
C13233 INVX1_LOC_2/Y NAND2X1_LOC_206/Y 0.39fF
C13234 NOR2X1_LOC_274/B NAND2X1_LOC_272/a_36_24# 0.00fF
C13235 NOR2X1_LOC_86/Y NOR2X1_LOC_384/Y 0.03fF
C13236 NOR2X1_LOC_728/B INVX1_LOC_15/A -0.01fF
C13237 INVX1_LOC_304/A NAND2X1_LOC_74/B 0.07fF
C13238 NOR2X1_LOC_82/A NOR2X1_LOC_516/a_36_216# 0.00fF
C13239 INVX1_LOC_174/A NOR2X1_LOC_550/B 0.06fF
C13240 NOR2X1_LOC_75/Y INVX1_LOC_33/A 0.03fF
C13241 INVX1_LOC_299/A NOR2X1_LOC_310/Y 0.16fF
C13242 INVX1_LOC_107/A INVX1_LOC_72/A 0.01fF
C13243 NOR2X1_LOC_828/Y INVX1_LOC_83/A 0.07fF
C13244 NOR2X1_LOC_454/Y INVX1_LOC_191/Y 0.00fF
C13245 NOR2X1_LOC_180/B NOR2X1_LOC_383/B 0.20fF
C13246 NOR2X1_LOC_82/A INVX1_LOC_8/A 0.56fF
C13247 INVX1_LOC_286/Y NOR2X1_LOC_152/a_36_216# 0.00fF
C13248 INVX1_LOC_77/A INVX1_LOC_31/A 0.02fF
C13249 NOR2X1_LOC_78/A NOR2X1_LOC_640/B 0.06fF
C13250 NAND2X1_LOC_639/A NOR2X1_LOC_430/Y 0.03fF
C13251 NAND2X1_LOC_457/a_36_24# INVX1_LOC_19/A 0.00fF
C13252 NOR2X1_LOC_666/Y INVX1_LOC_96/Y 0.01fF
C13253 VDD INVX1_LOC_240/Y 0.21fF
C13254 NOR2X1_LOC_596/A INVX1_LOC_72/A 0.12fF
C13255 INVX1_LOC_13/Y INVX1_LOC_137/A 0.04fF
C13256 INVX1_LOC_280/Y NAND2X1_LOC_493/Y 0.03fF
C13257 NOR2X1_LOC_598/B INVX1_LOC_120/A 0.03fF
C13258 NAND2X1_LOC_520/a_36_24# INVX1_LOC_217/A 0.02fF
C13259 INVX1_LOC_176/A INVX1_LOC_29/A 0.08fF
C13260 NOR2X1_LOC_791/B INVX1_LOC_24/A 0.03fF
C13261 INVX1_LOC_91/A INVX1_LOC_15/A 0.21fF
C13262 INVX1_LOC_147/A NAND2X1_LOC_61/Y 0.08fF
C13263 NOR2X1_LOC_322/Y NOR2X1_LOC_693/Y 0.10fF
C13264 NOR2X1_LOC_849/a_36_216# INVX1_LOC_77/A 0.01fF
C13265 INVX1_LOC_66/Y NOR2X1_LOC_814/A 0.03fF
C13266 INVX1_LOC_12/Y INVX1_LOC_19/A 0.11fF
C13267 INVX1_LOC_163/A NOR2X1_LOC_375/Y 0.00fF
C13268 NOR2X1_LOC_267/a_36_216# NOR2X1_LOC_773/Y 0.00fF
C13269 NAND2X1_LOC_181/Y INVX1_LOC_14/A 0.11fF
C13270 INVX1_LOC_5/A INVX1_LOC_83/A 8.22fF
C13271 INVX1_LOC_57/Y NAND2X1_LOC_833/Y 0.37fF
C13272 NOR2X1_LOC_160/B INVX1_LOC_266/Y 0.07fF
C13273 INVX1_LOC_1/A INVX1_LOC_25/Y 0.01fF
C13274 INVX1_LOC_105/A INVX1_LOC_159/A 0.15fF
C13275 INVX1_LOC_287/Y INVX1_LOC_75/A 0.01fF
C13276 NOR2X1_LOC_624/A INVX1_LOC_30/A 0.00fF
C13277 INVX1_LOC_126/Y INVX1_LOC_181/A 0.01fF
C13278 INVX1_LOC_140/A INVX1_LOC_53/A 0.05fF
C13279 INVX1_LOC_25/A INVX1_LOC_75/A 0.15fF
C13280 NOR2X1_LOC_569/A NOR2X1_LOC_383/B 0.01fF
C13281 NOR2X1_LOC_78/B NAND2X1_LOC_337/B 0.15fF
C13282 INVX1_LOC_1/A NOR2X1_LOC_302/B 0.02fF
C13283 INVX1_LOC_77/A INVX1_LOC_111/A 0.00fF
C13284 NOR2X1_LOC_68/A NOR2X1_LOC_520/B 0.07fF
C13285 INVX1_LOC_36/A INVX1_LOC_162/Y 0.15fF
C13286 NOR2X1_LOC_389/A INVX1_LOC_192/Y 0.03fF
C13287 NOR2X1_LOC_91/Y NAND2X1_LOC_640/Y 0.02fF
C13288 NOR2X1_LOC_295/Y INVX1_LOC_72/A 0.02fF
C13289 INPUT_6 D_INPUT_4 0.12fF
C13290 NOR2X1_LOC_68/A NAND2X1_LOC_325/Y 0.02fF
C13291 INVX1_LOC_14/A NAND2X1_LOC_390/A 0.11fF
C13292 NOR2X1_LOC_704/Y NOR2X1_LOC_383/B 0.01fF
C13293 INVX1_LOC_36/A NOR2X1_LOC_316/Y 0.00fF
C13294 NAND2X1_LOC_141/a_36_24# INVX1_LOC_89/A 0.00fF
C13295 INVX1_LOC_41/A NOR2X1_LOC_499/a_36_216# 0.00fF
C13296 NOR2X1_LOC_356/A INVX1_LOC_50/Y 0.07fF
C13297 INVX1_LOC_194/A INVX1_LOC_195/Y 0.02fF
C13298 NAND2X1_LOC_741/B NOR2X1_LOC_504/Y 0.29fF
C13299 NAND2X1_LOC_162/B INVX1_LOC_33/A 0.01fF
C13300 NOR2X1_LOC_795/Y INVX1_LOC_305/A 0.10fF
C13301 NAND2X1_LOC_53/Y NOR2X1_LOC_632/Y 0.02fF
C13302 NAND2X1_LOC_195/Y INVX1_LOC_266/Y -0.00fF
C13303 INVX1_LOC_2/Y NOR2X1_LOC_297/A 0.07fF
C13304 INVX1_LOC_186/A NOR2X1_LOC_727/B 0.15fF
C13305 INVX1_LOC_259/Y INVX1_LOC_311/A 0.00fF
C13306 INVX1_LOC_24/A NOR2X1_LOC_124/B 0.01fF
C13307 NOR2X1_LOC_577/Y INVX1_LOC_231/Y 0.04fF
C13308 NAND2X1_LOC_364/A NOR2X1_LOC_709/A 0.01fF
C13309 NOR2X1_LOC_456/a_36_216# INVX1_LOC_313/Y 0.00fF
C13310 NOR2X1_LOC_88/Y INVX1_LOC_203/A 0.26fF
C13311 NOR2X1_LOC_733/a_36_216# INVX1_LOC_266/Y 0.00fF
C13312 NOR2X1_LOC_379/Y NOR2X1_LOC_460/B 0.07fF
C13313 INVX1_LOC_119/A NAND2X1_LOC_586/a_36_24# 0.02fF
C13314 NOR2X1_LOC_716/B INVX1_LOC_33/A 0.08fF
C13315 INVX1_LOC_292/A NOR2X1_LOC_570/A 0.03fF
C13316 INVX1_LOC_276/A NOR2X1_LOC_68/A 0.72fF
C13317 INVX1_LOC_123/Y INVX1_LOC_63/A 0.03fF
C13318 NOR2X1_LOC_698/Y INVX1_LOC_15/A 0.09fF
C13319 INVX1_LOC_136/A NOR2X1_LOC_667/A 0.56fF
C13320 NOR2X1_LOC_208/Y INVX1_LOC_85/A 0.03fF
C13321 INVX1_LOC_24/A NOR2X1_LOC_802/A 0.33fF
C13322 INVX1_LOC_136/A INVX1_LOC_248/A 0.01fF
C13323 INVX1_LOC_13/A NOR2X1_LOC_590/A 0.17fF
C13324 INVX1_LOC_266/A NOR2X1_LOC_356/A 0.10fF
C13325 INVX1_LOC_34/A INVX1_LOC_155/A 0.03fF
C13326 INVX1_LOC_62/Y NOR2X1_LOC_537/Y 0.07fF
C13327 NOR2X1_LOC_74/A INVX1_LOC_50/Y 0.03fF
C13328 NAND2X1_LOC_190/Y INVX1_LOC_313/Y 0.01fF
C13329 NAND2X1_LOC_851/a_36_24# NOR2X1_LOC_109/Y 0.01fF
C13330 INVX1_LOC_200/A NAND2X1_LOC_861/Y 0.62fF
C13331 NOR2X1_LOC_273/a_36_216# NOR2X1_LOC_78/B 0.00fF
C13332 NOR2X1_LOC_596/A INVX1_LOC_192/Y 0.11fF
C13333 INVX1_LOC_12/A NAND2X1_LOC_802/Y 0.07fF
C13334 NAND2X1_LOC_738/B NAND2X1_LOC_729/B 0.03fF
C13335 INVX1_LOC_84/A INVX1_LOC_203/A 0.10fF
C13336 INVX1_LOC_50/A NOR2X1_LOC_56/Y 0.01fF
C13337 NOR2X1_LOC_384/Y INVX1_LOC_25/Y 0.57fF
C13338 NOR2X1_LOC_726/Y NOR2X1_LOC_209/a_36_216# 0.00fF
C13339 INVX1_LOC_278/A INVX1_LOC_91/A 0.10fF
C13340 NAND2X1_LOC_555/Y NOR2X1_LOC_415/A 0.04fF
C13341 INVX1_LOC_217/A NAND2X1_LOC_859/B 0.27fF
C13342 NOR2X1_LOC_9/Y INVX1_LOC_50/Y 0.03fF
C13343 INVX1_LOC_42/A INVX1_LOC_92/A 0.10fF
C13344 INVX1_LOC_18/A INVX1_LOC_16/A 0.33fF
C13345 NAND2X1_LOC_866/A NAND2X1_LOC_839/A 0.77fF
C13346 INVX1_LOC_191/Y INVX1_LOC_77/A 0.00fF
C13347 INVX1_LOC_30/A INPUT_5 0.07fF
C13348 INVX1_LOC_45/A INVX1_LOC_279/A 0.07fF
C13349 NOR2X1_LOC_536/A INVX1_LOC_94/Y 3.50fF
C13350 NAND2X1_LOC_728/Y INVX1_LOC_16/A 0.07fF
C13351 NOR2X1_LOC_590/A NOR2X1_LOC_246/A 0.00fF
C13352 INVX1_LOC_136/A NOR2X1_LOC_521/Y 0.05fF
C13353 INVX1_LOC_1/A INVX1_LOC_75/A 0.32fF
C13354 NAND2X1_LOC_563/Y NOR2X1_LOC_516/Y 0.01fF
C13355 INVX1_LOC_214/Y NOR2X1_LOC_152/Y 0.04fF
C13356 NOR2X1_LOC_598/B NOR2X1_LOC_542/B 0.01fF
C13357 NOR2X1_LOC_309/Y INVX1_LOC_162/Y 0.01fF
C13358 NOR2X1_LOC_759/Y NOR2X1_LOC_131/Y 0.01fF
C13359 NAND2X1_LOC_308/Y INVX1_LOC_240/A 0.02fF
C13360 NOR2X1_LOC_658/Y NOR2X1_LOC_366/Y 0.02fF
C13361 NOR2X1_LOC_223/B INVX1_LOC_91/A 0.01fF
C13362 NOR2X1_LOC_590/A NOR2X1_LOC_174/B 0.10fF
C13363 NOR2X1_LOC_843/A NOR2X1_LOC_174/a_36_216# 0.00fF
C13364 NOR2X1_LOC_331/B INVX1_LOC_271/Y 0.02fF
C13365 INVX1_LOC_50/A VDD 1.93fF
C13366 INVX1_LOC_266/A NOR2X1_LOC_74/A 0.04fF
C13367 NAND2X1_LOC_727/Y NAND2X1_LOC_731/Y 0.09fF
C13368 INVX1_LOC_247/A NOR2X1_LOC_678/A 0.01fF
C13369 NOR2X1_LOC_419/Y INVX1_LOC_40/A 0.12fF
C13370 INVX1_LOC_72/A NAND2X1_LOC_795/Y 0.03fF
C13371 NOR2X1_LOC_598/B INVX1_LOC_143/Y 0.42fF
C13372 NAND2X1_LOC_357/B NAND2X1_LOC_477/A 0.10fF
C13373 NOR2X1_LOC_784/Y INVX1_LOC_75/A 0.03fF
C13374 VDD NOR2X1_LOC_105/Y 0.33fF
C13375 NOR2X1_LOC_454/Y INVX1_LOC_6/A 0.04fF
C13376 NOR2X1_LOC_273/Y NOR2X1_LOC_589/A 0.79fF
C13377 NAND2X1_LOC_366/A NOR2X1_LOC_78/B 0.10fF
C13378 NOR2X1_LOC_794/a_36_216# NOR2X1_LOC_500/Y -0.00fF
C13379 NOR2X1_LOC_589/A NOR2X1_LOC_759/Y 0.19fF
C13380 NOR2X1_LOC_716/B INVX1_LOC_40/A 0.05fF
C13381 INVX1_LOC_203/Y NOR2X1_LOC_375/Y 0.01fF
C13382 NOR2X1_LOC_643/Y NOR2X1_LOC_516/B 0.01fF
C13383 NAND2X1_LOC_639/A INVX1_LOC_296/A 0.12fF
C13384 NOR2X1_LOC_350/A INVX1_LOC_22/A 0.02fF
C13385 INVX1_LOC_172/A INVX1_LOC_16/A 0.07fF
C13386 INVX1_LOC_57/Y NOR2X1_LOC_76/A 0.05fF
C13387 NOR2X1_LOC_536/A INVX1_LOC_181/A 0.07fF
C13388 NOR2X1_LOC_382/Y INPUT_1 0.07fF
C13389 NOR2X1_LOC_89/A NOR2X1_LOC_257/Y 0.00fF
C13390 NOR2X1_LOC_84/B NAND2X1_LOC_81/a_36_24# 0.02fF
C13391 NOR2X1_LOC_833/Y NOR2X1_LOC_834/a_36_216# 0.00fF
C13392 INVX1_LOC_102/A INVX1_LOC_63/A 0.08fF
C13393 NOR2X1_LOC_124/A INVX1_LOC_306/Y 0.01fF
C13394 NOR2X1_LOC_794/B INVX1_LOC_75/A 0.03fF
C13395 NOR2X1_LOC_795/Y NAND2X1_LOC_690/a_36_24# 0.06fF
C13396 INVX1_LOC_279/A INVX1_LOC_71/A 0.14fF
C13397 NAND2X1_LOC_555/Y NAND2X1_LOC_293/a_36_24# 0.01fF
C13398 NOR2X1_LOC_224/Y VDD 0.26fF
C13399 INVX1_LOC_224/Y NOR2X1_LOC_98/B 0.36fF
C13400 GATE_811 NAND2X1_LOC_852/Y 0.52fF
C13401 NOR2X1_LOC_261/a_36_216# INVX1_LOC_117/A 0.01fF
C13402 INVX1_LOC_34/A INVX1_LOC_316/Y 0.00fF
C13403 INVX1_LOC_151/Y NAND2X1_LOC_332/Y 0.01fF
C13404 NOR2X1_LOC_459/B INVX1_LOC_84/Y 0.00fF
C13405 INVX1_LOC_17/A INVX1_LOC_69/Y 0.09fF
C13406 INVX1_LOC_32/A INVX1_LOC_285/A 0.10fF
C13407 INVX1_LOC_78/A INVX1_LOC_92/A 0.34fF
C13408 NOR2X1_LOC_334/Y NOR2X1_LOC_600/a_36_216# 0.08fF
C13409 NOR2X1_LOC_340/A INVX1_LOC_29/A 0.03fF
C13410 NOR2X1_LOC_162/Y NOR2X1_LOC_160/Y 0.12fF
C13411 INVX1_LOC_206/A NOR2X1_LOC_203/Y 0.00fF
C13412 INVX1_LOC_32/A NOR2X1_LOC_814/A 0.07fF
C13413 INVX1_LOC_291/A NOR2X1_LOC_686/A 0.05fF
C13414 NAND2X1_LOC_840/Y INVX1_LOC_141/Y 0.01fF
C13415 INVX1_LOC_5/A INVX1_LOC_46/A 0.07fF
C13416 INVX1_LOC_28/A INVX1_LOC_18/A 0.42fF
C13417 INVX1_LOC_234/A NOR2X1_LOC_672/Y 0.03fF
C13418 NAND2X1_LOC_361/Y NOR2X1_LOC_785/Y 0.00fF
C13419 INVX1_LOC_203/A INVX1_LOC_15/A 0.28fF
C13420 NOR2X1_LOC_590/Y VDD 0.15fF
C13421 INVX1_LOC_38/A NOR2X1_LOC_591/A 0.01fF
C13422 NOR2X1_LOC_623/B NOR2X1_LOC_814/A 0.07fF
C13423 INVX1_LOC_23/A INVX1_LOC_9/A 0.41fF
C13424 NAND2X1_LOC_458/a_36_24# INVX1_LOC_118/A 0.00fF
C13425 NOR2X1_LOC_596/A INVX1_LOC_313/Y 0.03fF
C13426 INVX1_LOC_77/A INVX1_LOC_313/A 0.25fF
C13427 INVX1_LOC_33/A NOR2X1_LOC_326/Y 0.02fF
C13428 NOR2X1_LOC_78/B NOR2X1_LOC_773/Y 0.36fF
C13429 NOR2X1_LOC_717/B INVX1_LOC_33/A 0.06fF
C13430 NOR2X1_LOC_65/B INVX1_LOC_92/A 0.17fF
C13431 NAND2X1_LOC_714/B INVX1_LOC_20/A 0.03fF
C13432 INVX1_LOC_159/A NAND2X1_LOC_652/Y 0.00fF
C13433 NOR2X1_LOC_391/A NOR2X1_LOC_392/B 0.07fF
C13434 INVX1_LOC_16/A INVX1_LOC_34/Y 0.07fF
C13435 INVX1_LOC_201/Y NOR2X1_LOC_128/B 0.09fF
C13436 NAND2X1_LOC_711/B INVX1_LOC_28/A 0.00fF
C13437 NOR2X1_LOC_160/B INVX1_LOC_125/Y 0.12fF
C13438 INVX1_LOC_178/A INVX1_LOC_46/A 0.01fF
C13439 NOR2X1_LOC_513/Y NAND2X1_LOC_655/A 0.03fF
C13440 INVX1_LOC_306/A INVX1_LOC_8/A 0.02fF
C13441 NOR2X1_LOC_250/A NOR2X1_LOC_405/A 0.06fF
C13442 NOR2X1_LOC_248/Y NOR2X1_LOC_9/Y 0.02fF
C13443 INVX1_LOC_83/A NOR2X1_LOC_377/Y 0.01fF
C13444 INVX1_LOC_89/A NOR2X1_LOC_285/B 0.23fF
C13445 INVX1_LOC_172/A INVX1_LOC_28/A 3.28fF
C13446 NOR2X1_LOC_329/B NAND2X1_LOC_593/Y 0.19fF
C13447 INVX1_LOC_135/A NOR2X1_LOC_574/A 0.03fF
C13448 NOR2X1_LOC_445/a_36_216# NOR2X1_LOC_552/A 0.01fF
C13449 NAND2X1_LOC_849/A NAND2X1_LOC_837/Y 0.20fF
C13450 NOR2X1_LOC_609/Y INVX1_LOC_12/A 0.04fF
C13451 INVX1_LOC_58/A NOR2X1_LOC_88/a_36_216# 0.01fF
C13452 NAND2X1_LOC_227/Y NOR2X1_LOC_56/Y 0.02fF
C13453 NAND2X1_LOC_364/Y NOR2X1_LOC_775/Y 0.00fF
C13454 INVX1_LOC_56/A INVX1_LOC_56/Y 0.10fF
C13455 NOR2X1_LOC_494/Y INVX1_LOC_46/A 0.17fF
C13456 NOR2X1_LOC_328/Y INVX1_LOC_289/A 0.00fF
C13457 D_INPUT_4 NOR2X1_LOC_50/a_36_216# 0.00fF
C13458 NOR2X1_LOC_553/Y NOR2X1_LOC_388/a_36_216# 0.00fF
C13459 INVX1_LOC_30/A NOR2X1_LOC_7/Y 0.20fF
C13460 NOR2X1_LOC_354/B NOR2X1_LOC_354/Y 0.25fF
C13461 INVX1_LOC_105/Y INVX1_LOC_107/Y 0.25fF
C13462 INVX1_LOC_304/Y NAND2X1_LOC_861/Y 0.14fF
C13463 NOR2X1_LOC_816/A NOR2X1_LOC_164/Y 0.00fF
C13464 INVX1_LOC_2/A NOR2X1_LOC_60/a_36_216# 0.00fF
C13465 NOR2X1_LOC_773/Y NAND2X1_LOC_392/Y 0.01fF
C13466 INVX1_LOC_19/A NOR2X1_LOC_89/Y 0.00fF
C13467 INVX1_LOC_24/A NAND2X1_LOC_325/a_36_24# 0.01fF
C13468 NOR2X1_LOC_776/a_36_216# INVX1_LOC_143/Y 0.00fF
C13469 INVX1_LOC_290/A INVX1_LOC_22/A 0.17fF
C13470 NAND2X1_LOC_53/Y NAND2X1_LOC_39/Y 0.08fF
C13471 INVX1_LOC_232/Y D_INPUT_0 0.15fF
C13472 NOR2X1_LOC_779/Y INVX1_LOC_117/A 0.04fF
C13473 INVX1_LOC_86/Y NOR2X1_LOC_546/A -0.01fF
C13474 NOR2X1_LOC_507/A NAND2X1_LOC_505/a_36_24# 0.02fF
C13475 NOR2X1_LOC_151/Y INVX1_LOC_33/A 0.01fF
C13476 INVX1_LOC_14/A INVX1_LOC_117/A 0.07fF
C13477 NAND2X1_LOC_214/B NOR2X1_LOC_99/Y 0.04fF
C13478 NAND2X1_LOC_227/Y VDD 0.41fF
C13479 NAND2X1_LOC_89/a_36_24# NOR2X1_LOC_78/A 0.01fF
C13480 NOR2X1_LOC_828/A NOR2X1_LOC_714/Y -0.00fF
C13481 NAND2X1_LOC_429/a_36_24# INVX1_LOC_15/A 0.00fF
C13482 INVX1_LOC_104/A NOR2X1_LOC_564/Y 0.05fF
C13483 NAND2X1_LOC_337/B INVX1_LOC_46/A 0.14fF
C13484 NOR2X1_LOC_816/A INVX1_LOC_46/A 0.00fF
C13485 NOR2X1_LOC_168/Y INVX1_LOC_91/A 0.03fF
C13486 INVX1_LOC_77/A INVX1_LOC_6/A 0.13fF
C13487 INPUT_0 INVX1_LOC_155/A 0.03fF
C13488 INVX1_LOC_240/A NAND2X1_LOC_560/A 0.01fF
C13489 NAND2X1_LOC_9/Y INVX1_LOC_27/Y 0.07fF
C13490 INVX1_LOC_161/Y INVX1_LOC_12/Y 0.10fF
C13491 INVX1_LOC_136/A INVX1_LOC_304/A 0.04fF
C13492 NAND2X1_LOC_112/Y NAND2X1_LOC_656/Y 0.03fF
C13493 INVX1_LOC_50/A INVX1_LOC_133/A 0.00fF
C13494 INVX1_LOC_31/A NOR2X1_LOC_138/a_36_216# 0.01fF
C13495 NOR2X1_LOC_103/Y NOR2X1_LOC_98/B 0.03fF
C13496 INVX1_LOC_61/Y VDD 0.86fF
C13497 INVX1_LOC_57/A INVX1_LOC_49/Y 0.03fF
C13498 INVX1_LOC_13/Y NOR2X1_LOC_216/B 0.10fF
C13499 NOR2X1_LOC_220/A INVX1_LOC_313/Y 0.10fF
C13500 NOR2X1_LOC_264/Y INPUT_0 0.69fF
C13501 INVX1_LOC_284/Y NAND2X1_LOC_839/a_36_24# 0.00fF
C13502 INVX1_LOC_72/A NAND2X1_LOC_469/B 0.07fF
C13503 INVX1_LOC_85/A NOR2X1_LOC_208/A 0.20fF
C13504 NOR2X1_LOC_643/Y INVX1_LOC_315/Y 0.23fF
C13505 INVX1_LOC_271/A INVX1_LOC_272/A 0.13fF
C13506 NOR2X1_LOC_788/B NOR2X1_LOC_500/Y 0.00fF
C13507 INVX1_LOC_278/A INVX1_LOC_203/A 0.01fF
C13508 INVX1_LOC_136/A NOR2X1_LOC_670/Y 0.28fF
C13509 INVX1_LOC_50/Y NOR2X1_LOC_243/B 0.46fF
C13510 INVX1_LOC_18/A NOR2X1_LOC_35/Y 0.10fF
C13511 NOR2X1_LOC_6/B NOR2X1_LOC_9/Y 0.03fF
C13512 NOR2X1_LOC_201/A NOR2X1_LOC_861/Y 0.09fF
C13513 INVX1_LOC_266/A NOR2X1_LOC_650/a_36_216# 0.02fF
C13514 INVX1_LOC_290/Y INVX1_LOC_270/A 0.10fF
C13515 NOR2X1_LOC_780/B NOR2X1_LOC_155/A 0.00fF
C13516 NOR2X1_LOC_590/A INVX1_LOC_66/Y 0.04fF
C13517 INVX1_LOC_171/Y INVX1_LOC_285/A 0.08fF
C13518 INVX1_LOC_172/A NAND2X1_LOC_626/a_36_24# 0.01fF
C13519 INVX1_LOC_83/A NOR2X1_LOC_332/A 0.07fF
C13520 INVX1_LOC_300/Y INVX1_LOC_20/A 0.10fF
C13521 INVX1_LOC_124/A INVX1_LOC_6/A 0.44fF
C13522 INVX1_LOC_13/Y NAND2X1_LOC_477/Y 0.01fF
C13523 NOR2X1_LOC_653/B NOR2X1_LOC_653/Y 0.19fF
C13524 NAND2X1_LOC_361/Y INVX1_LOC_65/A 0.01fF
C13525 D_INPUT_0 NOR2X1_LOC_312/Y 0.07fF
C13526 INVX1_LOC_88/A NOR2X1_LOC_216/B 0.09fF
C13527 INVX1_LOC_31/A INVX1_LOC_9/A 0.12fF
C13528 INVX1_LOC_28/A NOR2X1_LOC_690/Y 0.00fF
C13529 NAND2X1_LOC_338/B INVX1_LOC_51/Y 0.03fF
C13530 INVX1_LOC_227/A INVX1_LOC_55/Y -0.00fF
C13531 INVX1_LOC_53/A INVX1_LOC_42/A 0.10fF
C13532 INVX1_LOC_76/Y INVX1_LOC_91/A 0.28fF
C13533 INVX1_LOC_135/A INVX1_LOC_175/Y 0.01fF
C13534 INPUT_0 INVX1_LOC_316/Y 0.04fF
C13535 INVX1_LOC_80/A NOR2X1_LOC_19/B 0.01fF
C13536 INVX1_LOC_174/A INVX1_LOC_75/Y 0.13fF
C13537 INVX1_LOC_5/A NOR2X1_LOC_671/Y 0.06fF
C13538 INVX1_LOC_24/A INVX1_LOC_37/Y 0.22fF
C13539 INVX1_LOC_224/Y NOR2X1_LOC_38/B 0.10fF
C13540 INVX1_LOC_105/A VDD 0.00fF
C13541 INVX1_LOC_300/Y NOR2X1_LOC_765/Y 0.28fF
C13542 NOR2X1_LOC_168/B NOR2X1_LOC_78/A 0.03fF
C13543 INVX1_LOC_304/A NOR2X1_LOC_278/A 0.04fF
C13544 INVX1_LOC_8/A INVX1_LOC_59/Y 0.12fF
C13545 NOR2X1_LOC_95/a_36_216# INVX1_LOC_77/Y 0.01fF
C13546 INVX1_LOC_27/A INVX1_LOC_272/A 0.07fF
C13547 NOR2X1_LOC_391/A NAND2X1_LOC_348/A 0.00fF
C13548 NOR2X1_LOC_405/A NOR2X1_LOC_709/A 0.01fF
C13549 VDD NOR2X1_LOC_679/B -0.00fF
C13550 NOR2X1_LOC_456/Y INVX1_LOC_4/A 0.07fF
C13551 NAND2X1_LOC_733/Y NAND2X1_LOC_802/Y 0.03fF
C13552 INVX1_LOC_279/Y INVX1_LOC_307/A 0.02fF
C13553 INVX1_LOC_11/A NOR2X1_LOC_450/B -0.02fF
C13554 NOR2X1_LOC_178/Y INVX1_LOC_127/Y 0.08fF
C13555 INVX1_LOC_28/A NAND2X1_LOC_105/a_36_24# 0.00fF
C13556 INVX1_LOC_30/Y NOR2X1_LOC_9/Y 0.04fF
C13557 NOR2X1_LOC_793/A INVX1_LOC_19/A 0.12fF
C13558 INVX1_LOC_89/A NAND2X1_LOC_291/a_36_24# 0.01fF
C13559 NAND2X1_LOC_859/a_36_24# NOR2X1_LOC_670/Y 0.00fF
C13560 NAND2X1_LOC_402/a_36_24# INVX1_LOC_242/A 0.01fF
C13561 NOR2X1_LOC_769/A INVX1_LOC_92/A 0.01fF
C13562 INVX1_LOC_160/A NOR2X1_LOC_325/A 0.04fF
C13563 D_INPUT_0 NOR2X1_LOC_97/A 0.02fF
C13564 INVX1_LOC_53/A INVX1_LOC_78/A 0.35fF
C13565 NOR2X1_LOC_615/Y NAND2X1_LOC_489/Y 0.06fF
C13566 INPUT_3 NOR2X1_LOC_814/A 0.27fF
C13567 NOR2X1_LOC_465/Y NOR2X1_LOC_678/A 0.00fF
C13568 INVX1_LOC_305/A NOR2X1_LOC_862/B 0.10fF
C13569 INVX1_LOC_103/A INVX1_LOC_29/A 0.07fF
C13570 D_INPUT_0 NOR2X1_LOC_391/Y 0.00fF
C13571 NOR2X1_LOC_570/B INVX1_LOC_44/A 0.01fF
C13572 NOR2X1_LOC_160/B INVX1_LOC_19/A 1.06fF
C13573 INVX1_LOC_209/A VDD 0.00fF
C13574 INVX1_LOC_17/A NOR2X1_LOC_89/A 0.13fF
C13575 INVX1_LOC_1/A INVX1_LOC_283/A 0.01fF
C13576 INVX1_LOC_21/A NAND2X1_LOC_647/B 0.04fF
C13577 NOR2X1_LOC_65/B INVX1_LOC_53/A 0.12fF
C13578 INVX1_LOC_33/A NOR2X1_LOC_209/B 0.22fF
C13579 NAND2X1_LOC_656/Y NOR2X1_LOC_78/A 0.07fF
C13580 NOR2X1_LOC_716/B NOR2X1_LOC_177/a_36_216# 0.01fF
C13581 NOR2X1_LOC_773/Y INVX1_LOC_46/A 0.10fF
C13582 NOR2X1_LOC_315/Y NOR2X1_LOC_536/A 0.12fF
C13583 NOR2X1_LOC_372/Y INVX1_LOC_84/A 0.07fF
C13584 NOR2X1_LOC_152/Y INVX1_LOC_92/A 0.08fF
C13585 INVX1_LOC_292/A INVX1_LOC_29/A 0.14fF
C13586 NOR2X1_LOC_272/Y NOR2X1_LOC_334/Y 0.10fF
C13587 INVX1_LOC_143/A NAND2X1_LOC_230/a_36_24# 0.01fF
C13588 NAND2X1_LOC_859/Y NOR2X1_LOC_670/a_36_216# 0.01fF
C13589 INVX1_LOC_113/Y INVX1_LOC_92/A 0.05fF
C13590 NOR2X1_LOC_471/Y NOR2X1_LOC_89/A 0.20fF
C13591 INVX1_LOC_58/Y NOR2X1_LOC_748/A 0.10fF
C13592 INVX1_LOC_14/A INVX1_LOC_3/Y 0.17fF
C13593 INVX1_LOC_132/Y NOR2X1_LOC_78/A 0.01fF
C13594 INVX1_LOC_75/A NOR2X1_LOC_188/A 0.26fF
C13595 NOR2X1_LOC_328/Y INVX1_LOC_37/A 0.02fF
C13596 NOR2X1_LOC_717/B NOR2X1_LOC_486/Y 0.05fF
C13597 NAND2X1_LOC_741/Y NOR2X1_LOC_829/A 0.02fF
C13598 NOR2X1_LOC_739/Y INVX1_LOC_15/A 0.01fF
C13599 INVX1_LOC_75/A NOR2X1_LOC_548/B 0.00fF
C13600 INVX1_LOC_297/Y NOR2X1_LOC_765/Y 0.01fF
C13601 INVX1_LOC_24/A NOR2X1_LOC_485/Y 0.03fF
C13602 INVX1_LOC_58/A NOR2X1_LOC_489/B 0.02fF
C13603 INVX1_LOC_77/A NOR2X1_LOC_117/Y 0.03fF
C13604 NOR2X1_LOC_456/Y NOR2X1_LOC_465/a_36_216# 0.00fF
C13605 NOR2X1_LOC_467/a_36_216# INVX1_LOC_37/A 0.00fF
C13606 NAND2X1_LOC_5/a_36_24# NAND2X1_LOC_141/Y 0.00fF
C13607 INVX1_LOC_124/A NOR2X1_LOC_79/A 0.16fF
C13608 NOR2X1_LOC_456/Y INVX1_LOC_64/A 0.05fF
C13609 INVX1_LOC_17/A INVX1_LOC_104/Y 0.01fF
C13610 INVX1_LOC_31/A NOR2X1_LOC_861/Y 0.07fF
C13611 NOR2X1_LOC_315/Y NAND2X1_LOC_93/B 0.46fF
C13612 NOR2X1_LOC_424/a_36_216# INVX1_LOC_37/A 0.00fF
C13613 NAND2X1_LOC_832/Y INVX1_LOC_6/A 0.02fF
C13614 INVX1_LOC_212/Y NAND2X1_LOC_574/A 0.11fF
C13615 INVX1_LOC_135/A NOR2X1_LOC_305/Y 0.10fF
C13616 NOR2X1_LOC_292/Y INVX1_LOC_286/A 0.13fF
C13617 INVX1_LOC_95/A NOR2X1_LOC_153/a_36_216# 0.00fF
C13618 NAND2X1_LOC_239/a_36_24# NAND2X1_LOC_798/B 0.00fF
C13619 NOR2X1_LOC_590/A INVX1_LOC_32/A 0.26fF
C13620 NAND2X1_LOC_9/Y INVX1_LOC_5/A 0.11fF
C13621 NAND2X1_LOC_116/A NAND2X1_LOC_85/Y 0.01fF
C13622 NOR2X1_LOC_310/a_36_216# INVX1_LOC_91/A 0.01fF
C13623 INVX1_LOC_256/A INVX1_LOC_94/Y 0.29fF
C13624 INVX1_LOC_233/A NAND2X1_LOC_552/A 0.02fF
C13625 NOR2X1_LOC_590/A NOR2X1_LOC_623/B 0.20fF
C13626 NAND2X1_LOC_129/a_36_24# NOR2X1_LOC_130/A 0.00fF
C13627 INVX1_LOC_214/Y INVX1_LOC_291/A 0.03fF
C13628 NAND2X1_LOC_652/Y NOR2X1_LOC_56/Y 0.02fF
C13629 NOR2X1_LOC_590/A NOR2X1_LOC_329/Y 0.18fF
C13630 NOR2X1_LOC_226/A INVX1_LOC_180/Y 0.02fF
C13631 INVX1_LOC_11/A NOR2X1_LOC_301/A 0.03fF
C13632 NAND2X1_LOC_803/B NAND2X1_LOC_175/Y 0.05fF
C13633 INVX1_LOC_255/Y NOR2X1_LOC_54/a_36_216# 0.03fF
C13634 INVX1_LOC_35/A NOR2X1_LOC_849/A 0.03fF
C13635 INVX1_LOC_124/A NOR2X1_LOC_117/Y 0.02fF
C13636 NOR2X1_LOC_669/Y NOR2X1_LOC_654/A 0.03fF
C13637 INVX1_LOC_34/A NOR2X1_LOC_662/A 0.08fF
C13638 NOR2X1_LOC_151/Y NOR2X1_LOC_486/Y 0.03fF
C13639 INVX1_LOC_77/A NOR2X1_LOC_633/A 0.03fF
C13640 NAND2X1_LOC_374/Y NOR2X1_LOC_88/Y 0.07fF
C13641 INVX1_LOC_279/A NOR2X1_LOC_331/B 0.14fF
C13642 INVX1_LOC_225/A NOR2X1_LOC_661/a_36_216# 0.00fF
C13643 INVX1_LOC_278/A NAND2X1_LOC_170/a_36_24# 0.00fF
C13644 INVX1_LOC_224/Y NOR2X1_LOC_468/Y 0.02fF
C13645 INVX1_LOC_45/A NOR2X1_LOC_38/B 0.03fF
C13646 INVX1_LOC_11/A NOR2X1_LOC_302/A 0.08fF
C13647 NOR2X1_LOC_359/Y NAND2X1_LOC_792/B 0.15fF
C13648 INVX1_LOC_66/A NOR2X1_LOC_536/A 0.07fF
C13649 INVX1_LOC_50/A NOR2X1_LOC_361/B 0.03fF
C13650 INVX1_LOC_233/A INVX1_LOC_178/A 0.10fF
C13651 NOR2X1_LOC_317/B INVX1_LOC_19/A 0.07fF
C13652 NOR2X1_LOC_548/a_36_216# INVX1_LOC_91/A 0.01fF
C13653 INVX1_LOC_298/Y INVX1_LOC_292/A 0.03fF
C13654 NOR2X1_LOC_590/A NAND2X1_LOC_175/Y 0.33fF
C13655 INVX1_LOC_21/A NOR2X1_LOC_109/a_36_216# 0.00fF
C13656 NOR2X1_LOC_312/Y NAND2X1_LOC_848/A 0.10fF
C13657 INVX1_LOC_123/A INVX1_LOC_91/A 0.02fF
C13658 INVX1_LOC_137/A NOR2X1_LOC_99/Y 0.32fF
C13659 INVX1_LOC_58/A INVX1_LOC_14/A 0.03fF
C13660 NAND2X1_LOC_652/Y VDD 0.26fF
C13661 INVX1_LOC_24/A NAND2X1_LOC_614/a_36_24# 0.00fF
C13662 NOR2X1_LOC_242/a_36_216# NOR2X1_LOC_865/Y 0.03fF
C13663 NOR2X1_LOC_798/A INVX1_LOC_5/A 0.03fF
C13664 INVX1_LOC_64/A NAND2X1_LOC_714/B 0.03fF
C13665 NOR2X1_LOC_160/B INVX1_LOC_26/Y 0.06fF
C13666 NOR2X1_LOC_716/B INVX1_LOC_106/Y 0.26fF
C13667 INVX1_LOC_136/A NOR2X1_LOC_248/A 0.01fF
C13668 NAND2X1_LOC_374/Y INVX1_LOC_84/A 0.94fF
C13669 INVX1_LOC_313/A INVX1_LOC_9/A 0.14fF
C13670 NAND2X1_LOC_149/Y INVX1_LOC_298/A 0.01fF
C13671 NOR2X1_LOC_763/Y NOR2X1_LOC_451/A 0.03fF
C13672 INVX1_LOC_64/A NAND2X1_LOC_561/B 0.03fF
C13673 NOR2X1_LOC_216/Y NOR2X1_LOC_363/Y 0.23fF
C13674 INVX1_LOC_230/Y NAND2X1_LOC_215/A 0.87fF
C13675 INPUT_6 NOR2X1_LOC_408/a_36_216# 0.00fF
C13676 INVX1_LOC_116/A INVX1_LOC_4/Y 0.01fF
C13677 NOR2X1_LOC_92/Y NOR2X1_LOC_291/Y 0.01fF
C13678 NOR2X1_LOC_488/Y NAND2X1_LOC_489/Y 0.06fF
C13679 NAND2X1_LOC_21/Y NAND2X1_LOC_429/a_36_24# 0.00fF
C13680 NOR2X1_LOC_186/Y NAND2X1_LOC_780/Y 0.01fF
C13681 NOR2X1_LOC_15/Y INVX1_LOC_306/Y 0.04fF
C13682 INVX1_LOC_182/Y NOR2X1_LOC_331/B 0.00fF
C13683 NAND2X1_LOC_703/Y INVX1_LOC_178/A 0.37fF
C13684 INVX1_LOC_217/Y INVX1_LOC_3/Y 0.03fF
C13685 INVX1_LOC_233/A NOR2X1_LOC_816/A 0.02fF
C13686 NOR2X1_LOC_225/a_36_216# NOR2X1_LOC_717/A 0.01fF
C13687 NOR2X1_LOC_78/B INVX1_LOC_263/Y 0.03fF
C13688 NOR2X1_LOC_128/B NAND2X1_LOC_574/A 0.01fF
C13689 INVX1_LOC_58/A NOR2X1_LOC_717/Y 0.01fF
C13690 INVX1_LOC_27/A NOR2X1_LOC_271/B 0.02fF
C13691 INVX1_LOC_316/Y NOR2X1_LOC_84/B 0.00fF
C13692 NAND2X1_LOC_361/Y INVX1_LOC_4/Y 0.08fF
C13693 NOR2X1_LOC_516/B INVX1_LOC_19/A 0.14fF
C13694 NOR2X1_LOC_180/B INVX1_LOC_179/A 0.01fF
C13695 NOR2X1_LOC_169/B INVX1_LOC_23/A 0.01fF
C13696 NAND2X1_LOC_573/Y NAND2X1_LOC_780/Y 0.14fF
C13697 NOR2X1_LOC_151/Y NOR2X1_LOC_833/a_36_216# 0.01fF
C13698 NOR2X1_LOC_788/B NOR2X1_LOC_445/B 0.02fF
C13699 INVX1_LOC_35/A NOR2X1_LOC_514/A 0.03fF
C13700 NOR2X1_LOC_78/B INVX1_LOC_42/A 0.03fF
C13701 INVX1_LOC_89/A NAND2X1_LOC_572/B 0.00fF
C13702 INVX1_LOC_49/A NOR2X1_LOC_278/Y 0.00fF
C13703 INVX1_LOC_22/A INVX1_LOC_261/Y 0.37fF
C13704 NOR2X1_LOC_769/A INVX1_LOC_53/A 0.11fF
C13705 INVX1_LOC_290/A INVX1_LOC_261/A 0.01fF
C13706 NAND2X1_LOC_854/B INVX1_LOC_264/A 0.10fF
C13707 NOR2X1_LOC_598/B NAND2X1_LOC_351/A 0.16fF
C13708 NOR2X1_LOC_350/A NOR2X1_LOC_843/B 0.03fF
C13709 INVX1_LOC_27/A INVX1_LOC_150/Y 0.12fF
C13710 INVX1_LOC_6/A INVX1_LOC_9/A 0.15fF
C13711 NAND2X1_LOC_35/Y NOR2X1_LOC_372/a_36_216# 0.01fF
C13712 INVX1_LOC_58/A NAND2X1_LOC_739/B 0.03fF
C13713 INVX1_LOC_35/A NOR2X1_LOC_859/A 0.00fF
C13714 NOR2X1_LOC_197/Y NOR2X1_LOC_197/B 0.03fF
C13715 NOR2X1_LOC_352/Y INVX1_LOC_15/A 0.00fF
C13716 INVX1_LOC_77/A INVX1_LOC_270/A 0.19fF
C13717 NOR2X1_LOC_270/Y NOR2X1_LOC_678/A 0.01fF
C13718 NAND2X1_LOC_218/B INVX1_LOC_25/A 0.11fF
C13719 NOR2X1_LOC_186/Y INVX1_LOC_141/Y 0.03fF
C13720 NAND2X1_LOC_703/Y NOR2X1_LOC_816/A 0.02fF
C13721 INVX1_LOC_17/A INVX1_LOC_224/A 0.03fF
C13722 INVX1_LOC_256/A INVX1_LOC_299/A 0.72fF
C13723 NOR2X1_LOC_186/Y INVX1_LOC_312/Y 0.07fF
C13724 INVX1_LOC_41/A NOR2X1_LOC_443/Y 0.04fF
C13725 NOR2X1_LOC_273/Y INVX1_LOC_64/A 0.07fF
C13726 INVX1_LOC_17/A INVX1_LOC_11/A 0.10fF
C13727 INVX1_LOC_39/A NOR2X1_LOC_382/Y 0.00fF
C13728 NOR2X1_LOC_152/Y INVX1_LOC_53/A 0.08fF
C13729 INVX1_LOC_50/A INVX1_LOC_153/Y 0.01fF
C13730 INVX1_LOC_120/A INVX1_LOC_29/A 0.49fF
C13731 INVX1_LOC_187/A INVX1_LOC_38/A 0.18fF
C13732 INVX1_LOC_53/Y INVX1_LOC_47/Y 0.09fF
C13733 INVX1_LOC_64/A NOR2X1_LOC_759/Y 1.02fF
C13734 NAND2X1_LOC_573/Y INVX1_LOC_141/Y 0.55fF
C13735 NAND2X1_LOC_477/A NOR2X1_LOC_282/Y 0.12fF
C13736 INVX1_LOC_34/A INVX1_LOC_57/A 0.22fF
C13737 NOR2X1_LOC_454/Y NOR2X1_LOC_230/a_36_216# 0.01fF
C13738 NOR2X1_LOC_78/B INVX1_LOC_78/A 0.18fF
C13739 INVX1_LOC_254/A NAND2X1_LOC_363/B 0.00fF
C13740 NOR2X1_LOC_773/Y NOR2X1_LOC_282/a_36_216# 0.01fF
C13741 NOR2X1_LOC_557/Y INVX1_LOC_29/Y 0.23fF
C13742 INVX1_LOC_64/A INVX1_LOC_202/A 0.03fF
C13743 NAND2X1_LOC_736/Y NAND2X1_LOC_725/Y 6.71fF
C13744 INVX1_LOC_186/A NOR2X1_LOC_640/Y 0.19fF
C13745 NOR2X1_LOC_817/Y NAND2X1_LOC_381/a_36_24# 0.01fF
C13746 INVX1_LOC_58/A INVX1_LOC_217/Y 0.00fF
C13747 NAND2X1_LOC_573/Y INVX1_LOC_312/Y 0.00fF
C13748 NAND2X1_LOC_222/B NAND2X1_LOC_555/Y 0.02fF
C13749 NOR2X1_LOC_471/Y INVX1_LOC_11/A 0.04fF
C13750 NOR2X1_LOC_454/Y INVX1_LOC_36/A 0.08fF
C13751 NOR2X1_LOC_226/A NOR2X1_LOC_278/Y 0.09fF
C13752 NAND2X1_LOC_559/Y NAND2X1_LOC_733/A 0.05fF
C13753 NOR2X1_LOC_361/B INVX1_LOC_61/Y 0.10fF
C13754 NAND2X1_LOC_724/A INVX1_LOC_141/Y 0.04fF
C13755 NOR2X1_LOC_817/Y NAND2X1_LOC_382/a_36_24# 0.00fF
C13756 INVX1_LOC_119/A NOR2X1_LOC_654/A 0.75fF
C13757 INVX1_LOC_33/Y INVX1_LOC_37/A 0.03fF
C13758 INVX1_LOC_64/A NOR2X1_LOC_550/B 0.10fF
C13759 INVX1_LOC_227/A INVX1_LOC_32/A 0.07fF
C13760 NOR2X1_LOC_411/A INVX1_LOC_237/Y 0.00fF
C13761 INVX1_LOC_124/A INVX1_LOC_270/A 0.10fF
C13762 NOR2X1_LOC_690/A NAND2X1_LOC_787/A 0.25fF
C13763 INVX1_LOC_45/A NOR2X1_LOC_468/Y 0.07fF
C13764 NOR2X1_LOC_160/B INVX1_LOC_161/Y 0.07fF
C13765 INVX1_LOC_50/A INVX1_LOC_177/A 0.09fF
C13766 NAND2X1_LOC_711/B NAND2X1_LOC_794/B 0.01fF
C13767 INPUT_0 NOR2X1_LOC_662/A 0.03fF
C13768 INVX1_LOC_13/Y NOR2X1_LOC_303/Y 0.00fF
C13769 NOR2X1_LOC_65/B NOR2X1_LOC_78/B 0.11fF
C13770 INVX1_LOC_35/A NOR2X1_LOC_758/Y 0.35fF
C13771 NAND2X1_LOC_725/Y INVX1_LOC_282/Y 0.12fF
C13772 NAND2X1_LOC_231/Y INVX1_LOC_57/A 0.01fF
C13773 INVX1_LOC_50/A INVX1_LOC_280/Y 0.10fF
C13774 INPUT_3 NOR2X1_LOC_590/A 0.03fF
C13775 NOR2X1_LOC_180/Y NOR2X1_LOC_678/A 0.01fF
C13776 INVX1_LOC_22/A INVX1_LOC_116/Y 0.00fF
C13777 NOR2X1_LOC_516/B INVX1_LOC_26/Y 0.03fF
C13778 INVX1_LOC_259/Y INVX1_LOC_259/A 0.06fF
C13779 INVX1_LOC_143/A INVX1_LOC_29/Y 0.01fF
C13780 NOR2X1_LOC_644/Y NOR2X1_LOC_717/A 0.12fF
C13781 INVX1_LOC_179/Y INVX1_LOC_23/A 0.02fF
C13782 NOR2X1_LOC_387/A NOR2X1_LOC_36/B 0.00fF
C13783 NOR2X1_LOC_447/B NOR2X1_LOC_506/Y 0.10fF
C13784 NOR2X1_LOC_634/A INVX1_LOC_143/Y 0.04fF
C13785 INVX1_LOC_83/A INVX1_LOC_78/A 1.11fF
C13786 NOR2X1_LOC_468/Y INVX1_LOC_71/A 0.03fF
C13787 INVX1_LOC_35/A NOR2X1_LOC_538/Y 0.01fF
C13788 INVX1_LOC_45/A NOR2X1_LOC_389/A 0.08fF
C13789 NOR2X1_LOC_772/a_36_216# INVX1_LOC_57/A 0.00fF
C13790 NAND2X1_LOC_724/Y INVX1_LOC_16/A 0.10fF
C13791 NAND2X1_LOC_72/Y INVX1_LOC_177/A 0.00fF
C13792 INVX1_LOC_203/Y INVX1_LOC_163/A 0.03fF
C13793 NOR2X1_LOC_298/Y NOR2X1_LOC_829/A 1.05fF
C13794 INVX1_LOC_64/A NOR2X1_LOC_41/Y 0.03fF
C13795 INVX1_LOC_278/A NAND2X1_LOC_374/Y 0.01fF
C13796 NAND2X1_LOC_190/Y INVX1_LOC_71/A 0.03fF
C13797 NOR2X1_LOC_639/B NAND2X1_LOC_451/Y 0.03fF
C13798 NOR2X1_LOC_91/A NOR2X1_LOC_561/Y 0.03fF
C13799 INVX1_LOC_315/Y INVX1_LOC_19/A 0.06fF
C13800 INVX1_LOC_237/Y INVX1_LOC_163/A -0.01fF
C13801 NOR2X1_LOC_458/B NOR2X1_LOC_678/A 0.00fF
C13802 INVX1_LOC_247/Y INVX1_LOC_292/A 0.01fF
C13803 INVX1_LOC_25/A INVX1_LOC_22/A 0.03fF
C13804 INVX1_LOC_41/A NAND2X1_LOC_347/B 0.03fF
C13805 INVX1_LOC_33/Y NOR2X1_LOC_743/Y 0.01fF
C13806 NOR2X1_LOC_279/Y INVX1_LOC_285/A 0.03fF
C13807 INVX1_LOC_38/A NOR2X1_LOC_629/Y 0.02fF
C13808 INVX1_LOC_17/A NOR2X1_LOC_433/A 0.17fF
C13809 INVX1_LOC_13/Y INVX1_LOC_54/Y 0.00fF
C13810 NOR2X1_LOC_763/Y INVX1_LOC_262/A 0.02fF
C13811 NOR2X1_LOC_561/Y INVX1_LOC_23/A 0.24fF
C13812 INVX1_LOC_34/A NOR2X1_LOC_666/Y 0.00fF
C13813 NOR2X1_LOC_15/Y INVX1_LOC_294/Y 0.04fF
C13814 NOR2X1_LOC_717/B NOR2X1_LOC_748/A 0.03fF
C13815 INVX1_LOC_17/A NOR2X1_LOC_593/Y 0.03fF
C13816 NOR2X1_LOC_437/Y NOR2X1_LOC_160/B 0.24fF
C13817 NAND2X1_LOC_17/a_36_24# INVX1_LOC_174/A 0.01fF
C13818 INVX1_LOC_90/A NOR2X1_LOC_621/A 0.38fF
C13819 NOR2X1_LOC_389/A INVX1_LOC_71/A 0.35fF
C13820 INVX1_LOC_27/A NOR2X1_LOC_87/Y 0.04fF
C13821 NOR2X1_LOC_597/Y NOR2X1_LOC_409/B 0.02fF
C13822 NOR2X1_LOC_197/A INVX1_LOC_49/A 0.00fF
C13823 INVX1_LOC_269/A NOR2X1_LOC_392/B 0.22fF
C13824 NOR2X1_LOC_382/Y INVX1_LOC_61/A 0.01fF
C13825 INVX1_LOC_147/Y NAND2X1_LOC_74/B 0.03fF
C13826 NOR2X1_LOC_151/Y NOR2X1_LOC_471/a_36_216# 0.00fF
C13827 NOR2X1_LOC_500/A NOR2X1_LOC_500/B 0.00fF
C13828 INVX1_LOC_17/A NOR2X1_LOC_52/B 0.46fF
C13829 NAND2X1_LOC_425/Y NAND2X1_LOC_427/a_36_24# 0.00fF
C13830 INVX1_LOC_20/A NAND2X1_LOC_74/B 0.56fF
C13831 NOR2X1_LOC_644/B INVX1_LOC_33/A 0.01fF
C13832 NAND2X1_LOC_703/Y NOR2X1_LOC_773/Y 0.03fF
C13833 NAND2X1_LOC_796/Y NOR2X1_LOC_109/Y 0.03fF
C13834 NOR2X1_LOC_526/Y NAND2X1_LOC_493/Y 0.38fF
C13835 INVX1_LOC_20/A NAND2X1_LOC_207/Y 0.16fF
C13836 INVX1_LOC_36/A INVX1_LOC_77/A 0.17fF
C13837 INVX1_LOC_221/Y NOR2X1_LOC_591/Y 0.02fF
C13838 INVX1_LOC_89/A INVX1_LOC_58/Y 0.07fF
C13839 INVX1_LOC_291/A INVX1_LOC_92/A 0.07fF
C13840 INVX1_LOC_69/Y INVX1_LOC_94/Y 0.00fF
C13841 NOR2X1_LOC_175/B INVX1_LOC_1/A 0.05fF
C13842 NOR2X1_LOC_794/B NOR2X1_LOC_348/B 0.00fF
C13843 NAND2X1_LOC_794/B NOR2X1_LOC_690/Y 0.02fF
C13844 NOR2X1_LOC_99/Y NOR2X1_LOC_216/B 0.94fF
C13845 NAND2X1_LOC_39/Y INVX1_LOC_12/A 0.03fF
C13846 INVX1_LOC_208/A NOR2X1_LOC_122/A 0.00fF
C13847 NOR2X1_LOC_690/A INVX1_LOC_30/A 0.10fF
C13848 NOR2X1_LOC_151/Y NOR2X1_LOC_748/A 0.10fF
C13849 NOR2X1_LOC_557/a_36_216# INVX1_LOC_47/Y 0.00fF
C13850 NOR2X1_LOC_590/A INVX1_LOC_158/A 0.09fF
C13851 INVX1_LOC_1/A NOR2X1_LOC_325/A 0.46fF
C13852 NOR2X1_LOC_596/A INVX1_LOC_71/A 0.03fF
C13853 D_INPUT_0 INVX1_LOC_50/Y 0.03fF
C13854 INVX1_LOC_1/A INVX1_LOC_22/A 0.55fF
C13855 INVX1_LOC_30/A NAND2X1_LOC_466/Y 0.02fF
C13856 NOR2X1_LOC_295/Y INVX1_LOC_45/A 0.01fF
C13857 INVX1_LOC_56/Y NOR2X1_LOC_271/a_36_216# 0.00fF
C13858 NOR2X1_LOC_155/A NOR2X1_LOC_831/B 0.16fF
C13859 NOR2X1_LOC_91/A NOR2X1_LOC_167/Y 0.03fF
C13860 INVX1_LOC_46/A INVX1_LOC_42/A 5.49fF
C13861 INVX1_LOC_72/A INVX1_LOC_63/Y 0.07fF
C13862 NAND2X1_LOC_729/Y NOR2X1_LOC_577/Y 0.32fF
C13863 NAND2X1_LOC_728/Y INVX1_LOC_231/Y 0.03fF
C13864 NAND2X1_LOC_721/A INVX1_LOC_102/A 0.02fF
C13865 NOR2X1_LOC_405/A NOR2X1_LOC_334/Y 0.00fF
C13866 INVX1_LOC_145/A INVX1_LOC_77/A 0.01fF
C13867 INPUT_0 INVX1_LOC_57/A 0.53fF
C13868 INVX1_LOC_230/Y NOR2X1_LOC_655/B 0.10fF
C13869 INVX1_LOC_2/A INVX1_LOC_236/Y 0.01fF
C13870 NOR2X1_LOC_189/A NAND2X1_LOC_711/B 0.03fF
C13871 NOR2X1_LOC_602/A NAND2X1_LOC_477/A 0.03fF
C13872 NOR2X1_LOC_208/Y INVX1_LOC_77/A 0.07fF
C13873 INVX1_LOC_233/A INVX1_LOC_140/A 0.10fF
C13874 NOR2X1_LOC_360/Y INVX1_LOC_155/Y 0.34fF
C13875 INVX1_LOC_50/A INVX1_LOC_285/Y 0.03fF
C13876 INPUT_3 NAND2X1_LOC_819/Y 0.01fF
C13877 INVX1_LOC_299/A NOR2X1_LOC_810/A 0.01fF
C13878 INVX1_LOC_124/A INVX1_LOC_36/A 0.21fF
C13879 NAND2X1_LOC_725/A NOR2X1_LOC_385/Y 0.34fF
C13880 NOR2X1_LOC_93/Y INVX1_LOC_90/A 0.02fF
C13881 INVX1_LOC_1/A NOR2X1_LOC_784/B 0.04fF
C13882 INVX1_LOC_278/A NOR2X1_LOC_184/a_36_216# 0.00fF
C13883 NAND2X1_LOC_35/Y NAND2X1_LOC_849/A 0.03fF
C13884 NOR2X1_LOC_794/B INVX1_LOC_22/A 0.07fF
C13885 NOR2X1_LOC_804/B INVX1_LOC_77/A 0.07fF
C13886 NOR2X1_LOC_468/Y NOR2X1_LOC_123/B 0.13fF
C13887 NOR2X1_LOC_381/Y D_INPUT_0 0.05fF
C13888 NOR2X1_LOC_712/Y NOR2X1_LOC_707/a_36_216# 0.00fF
C13889 NOR2X1_LOC_510/Y NAND2X1_LOC_652/Y 0.01fF
C13890 NOR2X1_LOC_295/Y INVX1_LOC_71/A 0.05fF
C13891 INVX1_LOC_45/A NOR2X1_LOC_220/A 0.01fF
C13892 NOR2X1_LOC_334/Y NOR2X1_LOC_857/A 0.01fF
C13893 NOR2X1_LOC_784/Y NOR2X1_LOC_784/B -0.00fF
C13894 NOR2X1_LOC_220/A NOR2X1_LOC_568/A 0.53fF
C13895 NOR2X1_LOC_589/A NOR2X1_LOC_276/Y 0.06fF
C13896 NAND2X1_LOC_740/Y NAND2X1_LOC_863/A 0.01fF
C13897 NOR2X1_LOC_599/A NAND2X1_LOC_853/Y 0.08fF
C13898 INVX1_LOC_103/A NAND2X1_LOC_140/A 0.00fF
C13899 D_INPUT_1 INVX1_LOC_91/A 0.20fF
C13900 INVX1_LOC_78/A INVX1_LOC_46/A 0.56fF
C13901 NOR2X1_LOC_321/Y INVX1_LOC_28/A 0.35fF
C13902 NOR2X1_LOC_309/Y INVX1_LOC_77/A 0.34fF
C13903 INVX1_LOC_269/A INVX1_LOC_90/A 0.17fF
C13904 NOR2X1_LOC_294/a_36_216# NOR2X1_LOC_516/B 0.00fF
C13905 NAND2X1_LOC_396/a_36_24# NOR2X1_LOC_123/B 0.00fF
C13906 NOR2X1_LOC_89/A NOR2X1_LOC_118/a_36_216# 0.01fF
C13907 NOR2X1_LOC_232/Y INVX1_LOC_90/A 0.10fF
C13908 NAND2X1_LOC_241/Y NOR2X1_LOC_693/Y 0.01fF
C13909 INVX1_LOC_269/A NOR2X1_LOC_389/B 0.10fF
C13910 NAND2X1_LOC_778/Y NOR2X1_LOC_74/A 0.10fF
C13911 INVX1_LOC_21/A INVX1_LOC_67/Y 0.02fF
C13912 NOR2X1_LOC_91/A INVX1_LOC_76/A 0.13fF
C13913 INVX1_LOC_7/A INVX1_LOC_31/A 0.19fF
C13914 NOR2X1_LOC_390/a_36_216# NOR2X1_LOC_142/Y 0.12fF
C13915 NOR2X1_LOC_75/Y INVX1_LOC_89/A 0.00fF
C13916 NOR2X1_LOC_679/a_36_216# NAND2X1_LOC_648/A 0.00fF
C13917 NOR2X1_LOC_703/B NOR2X1_LOC_553/Y 0.04fF
C13918 NOR2X1_LOC_568/A NOR2X1_LOC_548/Y 0.01fF
C13919 NAND2X1_LOC_475/Y NAND2X1_LOC_479/a_36_24# 0.07fF
C13920 INVX1_LOC_238/Y NOR2X1_LOC_299/Y 0.07fF
C13921 INVX1_LOC_10/Y INVX1_LOC_271/Y 0.13fF
C13922 INVX1_LOC_136/A NOR2X1_LOC_589/A 0.10fF
C13923 NOR2X1_LOC_65/B INVX1_LOC_46/A 0.11fF
C13924 NOR2X1_LOC_220/A INVX1_LOC_71/A 0.01fF
C13925 INVX1_LOC_290/A INVX1_LOC_18/A 0.17fF
C13926 NOR2X1_LOC_78/B NOR2X1_LOC_152/Y 0.01fF
C13927 NOR2X1_LOC_550/B INVX1_LOC_44/Y 0.39fF
C13928 NAND2X1_LOC_574/A NOR2X1_LOC_610/a_36_216# 0.01fF
C13929 NAND2X1_LOC_659/A INVX1_LOC_29/A 0.09fF
C13930 NAND2X1_LOC_646/a_36_24# INVX1_LOC_9/A 0.01fF
C13931 NOR2X1_LOC_774/a_36_216# INVX1_LOC_300/Y 0.01fF
C13932 NOR2X1_LOC_567/a_36_216# NOR2X1_LOC_748/A 0.12fF
C13933 NAND2X1_LOC_624/a_36_24# INVX1_LOC_15/A 0.00fF
C13934 NOR2X1_LOC_78/B INVX1_LOC_113/Y 0.04fF
C13935 INVX1_LOC_150/Y NOR2X1_LOC_772/A 0.02fF
C13936 NOR2X1_LOC_690/A NAND2X1_LOC_722/A 0.10fF
C13937 INVX1_LOC_269/A NAND2X1_LOC_348/A 0.01fF
C13938 NOR2X1_LOC_437/Y INVX1_LOC_208/A 0.03fF
C13939 NAND2X1_LOC_554/a_36_24# INVX1_LOC_223/A 0.00fF
C13940 NOR2X1_LOC_401/B NOR2X1_LOC_716/B 0.02fF
C13941 INVX1_LOC_23/A INVX1_LOC_76/A 4.40fF
C13942 NOR2X1_LOC_15/Y NOR2X1_LOC_74/A 0.22fF
C13943 NAND2X1_LOC_561/B INVX1_LOC_282/A 0.36fF
C13944 NOR2X1_LOC_155/A NOR2X1_LOC_270/a_36_216# 0.00fF
C13945 INVX1_LOC_49/A INVX1_LOC_83/Y 0.10fF
C13946 INVX1_LOC_124/A NOR2X1_LOC_309/Y 0.04fF
C13947 NOR2X1_LOC_402/a_36_216# NOR2X1_LOC_716/B 0.01fF
C13948 INVX1_LOC_91/A NOR2X1_LOC_652/Y 0.10fF
C13949 INVX1_LOC_77/Y NOR2X1_LOC_651/a_36_216# 0.01fF
C13950 NOR2X1_LOC_618/a_36_216# NOR2X1_LOC_419/Y 0.01fF
C13951 NAND2X1_LOC_177/a_36_24# NOR2X1_LOC_180/Y 0.00fF
C13952 NAND2X1_LOC_321/a_36_24# NOR2X1_LOC_356/A 0.00fF
C13953 NOR2X1_LOC_288/A NOR2X1_LOC_168/B 0.16fF
C13954 NOR2X1_LOC_637/Y INVX1_LOC_290/A 0.00fF
C13955 INVX1_LOC_83/A NOR2X1_LOC_554/B 0.20fF
C13956 NAND2X1_LOC_748/a_36_24# INVX1_LOC_123/A 0.01fF
C13957 NOR2X1_LOC_15/Y NOR2X1_LOC_9/Y 0.24fF
C13958 NOR2X1_LOC_536/A NAND2X1_LOC_99/A 0.06fF
C13959 NOR2X1_LOC_383/B INVX1_LOC_117/A 0.37fF
C13960 NOR2X1_LOC_667/Y NOR2X1_LOC_329/B 0.26fF
C13961 NOR2X1_LOC_627/Y NOR2X1_LOC_718/B 0.01fF
C13962 INVX1_LOC_71/A NOR2X1_LOC_548/Y 0.10fF
C13963 NAND2X1_LOC_36/A D_GATE_366 0.07fF
C13964 NAND2X1_LOC_357/B NOR2X1_LOC_312/a_36_216# 0.00fF
C13965 INVX1_LOC_299/A INVX1_LOC_69/Y 0.00fF
C13966 INVX1_LOC_136/A INVX1_LOC_171/A 0.04fF
C13967 NOR2X1_LOC_731/a_36_216# INVX1_LOC_85/Y 0.00fF
C13968 INVX1_LOC_226/Y NOR2X1_LOC_520/B 0.21fF
C13969 NOR2X1_LOC_68/A INVX1_LOC_148/Y 0.10fF
C13970 NAND2X1_LOC_207/B INVX1_LOC_19/A 0.22fF
C13971 NOR2X1_LOC_210/A INVX1_LOC_49/A 0.03fF
C13972 NOR2X1_LOC_804/B NOR2X1_LOC_687/Y 0.18fF
C13973 INVX1_LOC_266/Y NAND2X1_LOC_661/B 0.00fF
C13974 NOR2X1_LOC_189/A NOR2X1_LOC_690/Y 0.03fF
C13975 NOR2X1_LOC_246/A NAND2X1_LOC_357/a_36_24# 0.01fF
C13976 NOR2X1_LOC_175/A NOR2X1_LOC_537/Y 0.02fF
C13977 INVX1_LOC_180/A INVX1_LOC_10/A 0.02fF
C13978 INVX1_LOC_261/A INVX1_LOC_261/Y 0.15fF
C13979 NAND2X1_LOC_364/A NOR2X1_LOC_333/a_36_216# 0.01fF
C13980 INVX1_LOC_270/A INVX1_LOC_9/A 0.10fF
C13981 D_INPUT_0 NOR2X1_LOC_559/B 0.02fF
C13982 INVX1_LOC_83/A NOR2X1_LOC_152/Y 0.10fF
C13983 NOR2X1_LOC_391/A INVX1_LOC_33/A 0.01fF
C13984 INVX1_LOC_2/Y INVX1_LOC_38/Y 0.05fF
C13985 NAND2X1_LOC_93/B NAND2X1_LOC_99/A 0.01fF
C13986 NOR2X1_LOC_331/Y INVX1_LOC_6/A 0.01fF
C13987 NOR2X1_LOC_226/A NAND2X1_LOC_318/a_36_24# 0.01fF
C13988 NOR2X1_LOC_416/A INVX1_LOC_9/A 0.07fF
C13989 NOR2X1_LOC_229/Y INVX1_LOC_266/Y 0.01fF
C13990 INVX1_LOC_293/Y INVX1_LOC_4/A 0.07fF
C13991 INVX1_LOC_31/A NOR2X1_LOC_167/Y 0.03fF
C13992 NOR2X1_LOC_419/Y INVX1_LOC_89/A 0.00fF
C13993 INVX1_LOC_72/A INVX1_LOC_302/Y 0.07fF
C13994 NOR2X1_LOC_607/A INVX1_LOC_28/A 0.03fF
C13995 INVX1_LOC_24/A NOR2X1_LOC_736/Y 0.03fF
C13996 NOR2X1_LOC_558/A NAND2X1_LOC_474/Y 0.04fF
C13997 NOR2X1_LOC_218/A NOR2X1_LOC_269/Y 0.02fF
C13998 INVX1_LOC_67/A NAND2X1_LOC_140/A 0.00fF
C13999 INVX1_LOC_280/Y NOR2X1_LOC_701/a_36_216# 0.00fF
C14000 NOR2X1_LOC_716/B INVX1_LOC_89/A 0.08fF
C14001 NAND2X1_LOC_392/A NOR2X1_LOC_226/A 0.01fF
C14002 NOR2X1_LOC_188/A NOR2X1_LOC_274/B 0.10fF
C14003 NOR2X1_LOC_419/Y NAND2X1_LOC_508/A 0.03fF
C14004 NAND2X1_LOC_588/B NAND2X1_LOC_51/B 0.01fF
C14005 INVX1_LOC_45/Y INVX1_LOC_73/A 0.03fF
C14006 INVX1_LOC_136/A INVX1_LOC_222/A 0.01fF
C14007 INVX1_LOC_271/A NOR2X1_LOC_58/a_36_216# 0.00fF
C14008 D_INPUT_0 NOR2X1_LOC_6/B 0.39fF
C14009 NOR2X1_LOC_548/B NOR2X1_LOC_274/B 0.34fF
C14010 NAND2X1_LOC_74/B INVX1_LOC_4/A 0.03fF
C14011 INVX1_LOC_53/A INVX1_LOC_291/A 0.07fF
C14012 NAND2X1_LOC_222/A NAND2X1_LOC_574/A 0.04fF
C14013 NOR2X1_LOC_1/a_36_216# INPUT_5 0.00fF
C14014 NAND2X1_LOC_114/B NAND2X1_LOC_642/Y 0.04fF
C14015 NOR2X1_LOC_67/Y INVX1_LOC_32/A 0.04fF
C14016 NOR2X1_LOC_171/Y NOR2X1_LOC_433/A 0.05fF
C14017 INVX1_LOC_296/Y NAND2X1_LOC_770/Y 0.45fF
C14018 INVX1_LOC_3/A NAND2X1_LOC_99/A 0.01fF
C14019 INVX1_LOC_45/A NAND2X1_LOC_498/a_36_24# 0.00fF
C14020 NOR2X1_LOC_294/a_36_216# INVX1_LOC_315/Y 0.00fF
C14021 NOR2X1_LOC_488/Y NAND2X1_LOC_564/B 0.00fF
C14022 INVX1_LOC_59/A NOR2X1_LOC_813/Y 0.02fF
C14023 NAND2X1_LOC_672/a_36_24# INVX1_LOC_315/Y 0.00fF
C14024 NAND2X1_LOC_348/A NOR2X1_LOC_360/a_36_216# 0.00fF
C14025 INVX1_LOC_223/A NOR2X1_LOC_318/B 0.00fF
C14026 INVX1_LOC_2/A NOR2X1_LOC_312/Y 0.15fF
C14027 INVX1_LOC_55/Y INVX1_LOC_104/A 0.07fF
C14028 INVX1_LOC_197/Y NAND2X1_LOC_462/B 0.35fF
C14029 NOR2X1_LOC_636/B INVX1_LOC_37/A 0.01fF
C14030 NOR2X1_LOC_89/A INVX1_LOC_94/Y 0.08fF
C14031 NAND2X1_LOC_860/Y NAND2X1_LOC_392/Y 0.15fF
C14032 D_INPUT_1 NOR2X1_LOC_179/Y 0.03fF
C14033 NAND2X1_LOC_555/Y INVX1_LOC_74/A 0.05fF
C14034 INVX1_LOC_59/A INVX1_LOC_280/A 0.13fF
C14035 INVX1_LOC_64/A NOR2X1_LOC_13/a_36_216# 0.01fF
C14036 INVX1_LOC_83/A NOR2X1_LOC_307/B 0.51fF
C14037 INVX1_LOC_58/A NOR2X1_LOC_127/Y 0.08fF
C14038 NOR2X1_LOC_93/Y NOR2X1_LOC_96/Y 0.01fF
C14039 INVX1_LOC_59/A NOR2X1_LOC_94/Y 0.01fF
C14040 INVX1_LOC_312/Y NAND2X1_LOC_642/Y 0.39fF
C14041 INVX1_LOC_11/A NOR2X1_LOC_706/B 0.02fF
C14042 NAND2X1_LOC_395/a_36_24# NOR2X1_LOC_123/B 0.00fF
C14043 NOR2X1_LOC_446/A INVX1_LOC_37/A 0.02fF
C14044 NOR2X1_LOC_577/Y NOR2X1_LOC_188/A 0.01fF
C14045 NOR2X1_LOC_478/A INVX1_LOC_115/A 0.03fF
C14046 INVX1_LOC_31/A INVX1_LOC_76/A 0.45fF
C14047 INVX1_LOC_26/Y NAND2X1_LOC_207/B 0.03fF
C14048 INVX1_LOC_12/A NAND2X1_LOC_61/Y 0.02fF
C14049 INVX1_LOC_232/Y INPUT_1 0.08fF
C14050 NOR2X1_LOC_232/Y NAND2X1_LOC_849/B 0.06fF
C14051 INVX1_LOC_269/A INVX1_LOC_38/A 0.09fF
C14052 NOR2X1_LOC_742/A INVX1_LOC_85/A 0.02fF
C14053 NAND2X1_LOC_190/Y NOR2X1_LOC_331/B 0.03fF
C14054 INVX1_LOC_130/A VDD 0.12fF
C14055 NOR2X1_LOC_238/Y NOR2X1_LOC_45/B 0.00fF
C14056 NAND2X1_LOC_631/a_36_24# INVX1_LOC_309/A 0.00fF
C14057 NOR2X1_LOC_191/B NOR2X1_LOC_192/A 0.02fF
C14058 INVX1_LOC_13/Y INVX1_LOC_35/Y 0.05fF
C14059 NOR2X1_LOC_403/B INVX1_LOC_91/A 0.04fF
C14060 NOR2X1_LOC_89/A INVX1_LOC_181/A 0.11fF
C14061 INVX1_LOC_75/A NOR2X1_LOC_87/B 0.01fF
C14062 NOR2X1_LOC_763/Y GATE_662 0.33fF
C14063 NOR2X1_LOC_773/Y NAND2X1_LOC_842/B 0.21fF
C14064 INVX1_LOC_30/Y D_INPUT_0 0.03fF
C14065 INVX1_LOC_138/Y NAND2X1_LOC_206/Y 0.04fF
C14066 INVX1_LOC_136/A INVX1_LOC_20/A 0.17fF
C14067 NOR2X1_LOC_382/Y D_INPUT_3 0.07fF
C14068 INVX1_LOC_32/A NOR2X1_LOC_415/Y 0.00fF
C14069 NOR2X1_LOC_860/a_36_216# NAND2X1_LOC_206/Y 0.01fF
C14070 NOR2X1_LOC_392/Y NAND2X1_LOC_219/B 0.02fF
C14071 INVX1_LOC_245/Y NOR2X1_LOC_684/Y 0.02fF
C14072 NAND2X1_LOC_276/Y INVX1_LOC_123/A 0.07fF
C14073 INVX1_LOC_135/A INVX1_LOC_279/A 0.02fF
C14074 NAND2X1_LOC_214/B NOR2X1_LOC_673/A 0.06fF
C14075 NOR2X1_LOC_20/Y NOR2X1_LOC_629/Y 0.01fF
C14076 NOR2X1_LOC_68/A INVX1_LOC_115/A 0.01fF
C14077 NAND2X1_LOC_740/A NAND2X1_LOC_729/B 0.01fF
C14078 NAND2X1_LOC_364/Y NOR2X1_LOC_78/A 0.01fF
C14079 INVX1_LOC_96/Y NOR2X1_LOC_74/A 0.18fF
C14080 NAND2X1_LOC_861/Y NAND2X1_LOC_392/Y 0.01fF
C14081 D_INPUT_7 VDD 1.05fF
C14082 NOR2X1_LOC_367/B INVX1_LOC_6/A 0.13fF
C14083 NOR2X1_LOC_470/A INVX1_LOC_89/A 0.04fF
C14084 NAND2X1_LOC_79/Y INVX1_LOC_112/A 0.00fF
C14085 NAND2X1_LOC_79/Y INVX1_LOC_59/Y 0.00fF
C14086 INVX1_LOC_21/A INVX1_LOC_285/A 0.14fF
C14087 NOR2X1_LOC_791/B VDD 0.24fF
C14088 NOR2X1_LOC_389/A NOR2X1_LOC_331/B 0.10fF
C14089 NOR2X1_LOC_272/Y NOR2X1_LOC_813/a_36_216# 0.01fF
C14090 INVX1_LOC_277/Y INVX1_LOC_117/A 0.04fF
C14091 NOR2X1_LOC_424/Y INVX1_LOC_89/A 0.04fF
C14092 INVX1_LOC_305/A NAND2X1_LOC_277/a_36_24# 0.01fF
C14093 NAND2X1_LOC_563/A NAND2X1_LOC_348/A 0.03fF
C14094 INVX1_LOC_71/A NAND2X1_LOC_469/B 2.00fF
C14095 NOR2X1_LOC_547/B INVX1_LOC_158/Y 0.01fF
C14096 INVX1_LOC_27/A NOR2X1_LOC_673/A 0.21fF
C14097 NAND2X1_LOC_577/A NOR2X1_LOC_536/A 0.06fF
C14098 NOR2X1_LOC_215/Y NOR2X1_LOC_357/Y 0.05fF
C14099 NOR2X1_LOC_717/B INVX1_LOC_89/A 0.03fF
C14100 INVX1_LOC_64/A NAND2X1_LOC_74/B 0.03fF
C14101 INVX1_LOC_21/A NOR2X1_LOC_814/A 0.52fF
C14102 NOR2X1_LOC_188/A NOR2X1_LOC_346/B 0.04fF
C14103 NOR2X1_LOC_861/Y NOR2X1_LOC_416/A 0.02fF
C14104 NAND2X1_LOC_586/a_36_24# NAND2X1_LOC_453/A 0.00fF
C14105 NOR2X1_LOC_82/A INVX1_LOC_70/A 0.03fF
C14106 NAND2X1_LOC_538/Y NOR2X1_LOC_88/Y 0.07fF
C14107 NOR2X1_LOC_71/Y NOR2X1_LOC_76/A 0.04fF
C14108 INVX1_LOC_23/A INVX1_LOC_127/Y 0.01fF
C14109 NAND2X1_LOC_9/Y INVX1_LOC_42/A 0.46fF
C14110 NOR2X1_LOC_574/A NOR2X1_LOC_45/B 0.04fF
C14111 NOR2X1_LOC_591/Y INVX1_LOC_91/A 0.03fF
C14112 NOR2X1_LOC_175/B NOR2X1_LOC_548/B 0.16fF
C14113 INVX1_LOC_284/Y INVX1_LOC_118/A 0.16fF
C14114 NOR2X1_LOC_717/B NAND2X1_LOC_176/a_36_24# 0.00fF
C14115 INVX1_LOC_233/A INVX1_LOC_42/A 0.07fF
C14116 NOR2X1_LOC_272/Y NAND2X1_LOC_773/B 0.10fF
C14117 NOR2X1_LOC_444/a_36_216# INVX1_LOC_15/A 0.01fF
C14118 INVX1_LOC_81/A VDD 0.37fF
C14119 INVX1_LOC_162/Y INVX1_LOC_93/Y 0.06fF
C14120 NOR2X1_LOC_140/A INVX1_LOC_84/A 0.03fF
C14121 NOR2X1_LOC_172/Y NAND2X1_LOC_434/a_36_24# 0.00fF
C14122 INVX1_LOC_174/Y INVX1_LOC_75/A 0.01fF
C14123 NOR2X1_LOC_152/Y INVX1_LOC_46/A 0.08fF
C14124 INVX1_LOC_150/Y NOR2X1_LOC_216/B 0.10fF
C14125 INVX1_LOC_36/A INVX1_LOC_9/A 1.82fF
C14126 NOR2X1_LOC_82/A INVX1_LOC_123/Y 0.03fF
C14127 NOR2X1_LOC_188/A INVX1_LOC_22/A 0.10fF
C14128 INVX1_LOC_50/A INVX1_LOC_4/Y 0.10fF
C14129 INVX1_LOC_5/A INVX1_LOC_284/A 0.31fF
C14130 INVX1_LOC_113/Y INVX1_LOC_46/A 0.01fF
C14131 NAND2X1_LOC_352/B NOR2X1_LOC_155/A 0.02fF
C14132 INVX1_LOC_256/Y INVX1_LOC_98/A 0.21fF
C14133 NAND2X1_LOC_538/Y INVX1_LOC_84/A 0.72fF
C14134 NOR2X1_LOC_548/B INVX1_LOC_22/A 0.10fF
C14135 NAND2X1_LOC_27/a_36_24# NAND2X1_LOC_207/Y 0.01fF
C14136 INVX1_LOC_53/A NOR2X1_LOC_609/Y 0.03fF
C14137 NOR2X1_LOC_644/A NOR2X1_LOC_180/B 0.03fF
C14138 NAND2X1_LOC_656/A NOR2X1_LOC_536/A 0.02fF
C14139 NAND2X1_LOC_553/A INVX1_LOC_42/A 0.02fF
C14140 NOR2X1_LOC_355/A NOR2X1_LOC_216/Y 0.03fF
C14141 NOR2X1_LOC_373/Y NOR2X1_LOC_322/Y 0.01fF
C14142 INVX1_LOC_1/A INVX1_LOC_186/Y 0.07fF
C14143 NAND2X1_LOC_206/B NOR2X1_LOC_849/A 0.01fF
C14144 INVX1_LOC_81/Y NOR2X1_LOC_155/A 0.01fF
C14145 NOR2X1_LOC_278/A INVX1_LOC_20/A 0.05fF
C14146 INVX1_LOC_251/Y INVX1_LOC_95/Y 0.01fF
C14147 NOR2X1_LOC_484/Y NOR2X1_LOC_536/A 0.02fF
C14148 INVX1_LOC_178/A INVX1_LOC_284/A 0.10fF
C14149 NOR2X1_LOC_798/A INVX1_LOC_42/A 0.03fF
C14150 NOR2X1_LOC_596/A NOR2X1_LOC_331/B 1.86fF
C14151 INVX1_LOC_192/A VDD 0.12fF
C14152 NOR2X1_LOC_816/A INVX1_LOC_119/Y 0.02fF
C14153 NOR2X1_LOC_124/B VDD 0.00fF
C14154 NOR2X1_LOC_151/Y INVX1_LOC_89/A 0.22fF
C14155 NOR2X1_LOC_530/Y INVX1_LOC_84/A 0.07fF
C14156 INVX1_LOC_1/A NOR2X1_LOC_777/B 0.05fF
C14157 NOR2X1_LOC_561/Y INVX1_LOC_6/A 0.08fF
C14158 INVX1_LOC_83/A INVX1_LOC_158/Y 0.13fF
C14159 NOR2X1_LOC_384/Y NOR2X1_LOC_88/A 0.15fF
C14160 NOR2X1_LOC_208/Y INVX1_LOC_9/A 0.03fF
C14161 INVX1_LOC_77/A NOR2X1_LOC_865/A 0.04fF
C14162 NAND2X1_LOC_9/Y INVX1_LOC_78/A 0.01fF
C14163 INVX1_LOC_135/A NAND2X1_LOC_858/B 0.10fF
C14164 INVX1_LOC_268/A NOR2X1_LOC_45/B 0.20fF
C14165 NOR2X1_LOC_828/B NOR2X1_LOC_738/A 0.07fF
C14166 NAND2X1_LOC_72/Y INVX1_LOC_4/Y 0.02fF
C14167 NOR2X1_LOC_802/A VDD 0.24fF
C14168 INVX1_LOC_233/A INVX1_LOC_78/A 0.08fF
C14169 NOR2X1_LOC_43/Y INVX1_LOC_22/A 0.07fF
C14170 NOR2X1_LOC_784/Y NOR2X1_LOC_777/B 0.01fF
C14171 NOR2X1_LOC_494/Y INVX1_LOC_284/A 0.01fF
C14172 NOR2X1_LOC_520/A INVX1_LOC_176/A 0.01fF
C14173 NAND2X1_LOC_577/A NOR2X1_LOC_649/B 0.08fF
C14174 NOR2X1_LOC_447/A INVX1_LOC_23/A 0.08fF
C14175 INVX1_LOC_2/A NAND2X1_LOC_287/B 0.08fF
C14176 NAND2X1_LOC_656/A NAND2X1_LOC_93/B 0.02fF
C14177 NOR2X1_LOC_763/A NAND2X1_LOC_95/a_36_24# 0.01fF
C14178 INVX1_LOC_58/A NOR2X1_LOC_383/B 0.08fF
C14179 NAND2X1_LOC_9/Y NOR2X1_LOC_65/B 0.09fF
C14180 NOR2X1_LOC_251/a_36_216# INVX1_LOC_32/A 0.01fF
C14181 INVX1_LOC_17/A NAND2X1_LOC_254/Y 0.00fF
C14182 INVX1_LOC_43/Y NAND2X1_LOC_74/B 0.01fF
C14183 NAND2X1_LOC_802/A NOR2X1_LOC_510/B 0.10fF
C14184 NAND2X1_LOC_672/B VDD 0.01fF
C14185 NAND2X1_LOC_807/Y NOR2X1_LOC_167/Y 0.02fF
C14186 NOR2X1_LOC_798/A INVX1_LOC_78/A 0.03fF
C14187 INVX1_LOC_55/Y INVX1_LOC_206/Y 0.09fF
C14188 INVX1_LOC_49/A NOR2X1_LOC_809/B 0.07fF
C14189 NAND2X1_LOC_860/Y INVX1_LOC_46/A 0.02fF
C14190 INVX1_LOC_61/Y NAND2X1_LOC_81/B 0.02fF
C14191 NAND2X1_LOC_347/a_36_24# INVX1_LOC_117/A 0.00fF
C14192 NOR2X1_LOC_646/A VDD 0.21fF
C14193 INVX1_LOC_30/A INVX1_LOC_262/Y 0.06fF
C14194 INVX1_LOC_233/Y INVX1_LOC_50/A 0.01fF
C14195 INPUT_3 NOR2X1_LOC_67/Y 0.01fF
C14196 INVX1_LOC_35/A INVX1_LOC_270/Y 0.05fF
C14197 NAND2X1_LOC_656/A NOR2X1_LOC_649/B 0.01fF
C14198 NOR2X1_LOC_860/B NOR2X1_LOC_243/B 0.21fF
C14199 D_INPUT_0 NOR2X1_LOC_124/A 0.00fF
C14200 NAND2X1_LOC_656/A INVX1_LOC_3/A 1.10fF
C14201 NOR2X1_LOC_103/Y INVX1_LOC_251/A 0.01fF
C14202 NOR2X1_LOC_598/B NAND2X1_LOC_46/a_36_24# 0.02fF
C14203 NOR2X1_LOC_497/Y INVX1_LOC_91/A 0.04fF
C14204 NOR2X1_LOC_65/B NOR2X1_LOC_798/A 0.03fF
C14205 INVX1_LOC_100/Y INVX1_LOC_102/Y 0.01fF
C14206 NOR2X1_LOC_178/Y INVX1_LOC_23/A 0.21fF
C14207 NAND2X1_LOC_9/Y INVX1_LOC_152/Y 0.02fF
C14208 INVX1_LOC_126/A NOR2X1_LOC_130/A 0.03fF
C14209 NOR2X1_LOC_90/a_36_216# INVX1_LOC_284/A 0.01fF
C14210 NOR2X1_LOC_220/A NOR2X1_LOC_331/B 0.10fF
C14211 NOR2X1_LOC_264/a_36_216# NAND2X1_LOC_223/A 0.03fF
C14212 NOR2X1_LOC_6/B INVX1_LOC_46/Y 0.23fF
C14213 NOR2X1_LOC_733/Y NOR2X1_LOC_74/A 0.05fF
C14214 NOR2X1_LOC_234/a_36_216# INVX1_LOC_35/Y 0.01fF
C14215 NAND2X1_LOC_866/B NOR2X1_LOC_824/Y 0.10fF
C14216 NOR2X1_LOC_180/B NOR2X1_LOC_540/B 0.01fF
C14217 INVX1_LOC_77/A INVX1_LOC_63/A 0.10fF
C14218 INVX1_LOC_144/Y INVX1_LOC_54/A 0.00fF
C14219 NOR2X1_LOC_601/a_36_216# NOR2X1_LOC_678/A 0.00fF
C14220 INVX1_LOC_313/A INVX1_LOC_76/A 0.01fF
C14221 INVX1_LOC_193/Y NOR2X1_LOC_706/Y 0.01fF
C14222 INVX1_LOC_11/A INVX1_LOC_94/Y 0.03fF
C14223 NOR2X1_LOC_194/Y INVX1_LOC_113/A 0.01fF
C14224 NAND2X1_LOC_783/A NOR2X1_LOC_111/A 0.12fF
C14225 NAND2X1_LOC_140/A NOR2X1_LOC_137/Y 0.26fF
C14226 NAND2X1_LOC_861/Y INVX1_LOC_46/A 0.03fF
C14227 NAND2X1_LOC_866/B INVX1_LOC_76/A 0.07fF
C14228 NOR2X1_LOC_78/B INVX1_LOC_291/A 0.08fF
C14229 NAND2X1_LOC_860/A INVX1_LOC_13/Y 0.68fF
C14230 NAND2X1_LOC_740/B INVX1_LOC_291/Y 0.01fF
C14231 NOR2X1_LOC_130/A NOR2X1_LOC_111/A 0.07fF
C14232 INVX1_LOC_1/A NOR2X1_LOC_843/B 0.17fF
C14233 NOR2X1_LOC_532/Y VDD 0.34fF
C14234 NOR2X1_LOC_222/Y NAND2X1_LOC_93/B 0.10fF
C14235 NOR2X1_LOC_45/Y INVX1_LOC_128/Y 0.21fF
C14236 NOR2X1_LOC_637/Y INVX1_LOC_261/Y 0.00fF
C14237 INVX1_LOC_223/Y INVX1_LOC_58/Y 0.03fF
C14238 NAND2X1_LOC_7/Y NAND2X1_LOC_63/Y 0.02fF
C14239 NAND2X1_LOC_67/Y INVX1_LOC_270/A 0.08fF
C14240 INVX1_LOC_163/A INVX1_LOC_23/A 0.00fF
C14241 INVX1_LOC_188/A NOR2X1_LOC_465/Y 0.13fF
C14242 NOR2X1_LOC_174/A VDD 0.02fF
C14243 NAND2X1_LOC_35/Y NOR2X1_LOC_291/Y 0.03fF
C14244 NOR2X1_LOC_222/Y NAND2X1_LOC_425/Y 0.01fF
C14245 INVX1_LOC_90/A INVX1_LOC_12/Y 0.01fF
C14246 INVX1_LOC_16/A NOR2X1_LOC_433/Y 0.17fF
C14247 INVX1_LOC_50/A NOR2X1_LOC_205/Y 0.01fF
C14248 NAND2X1_LOC_569/A INVX1_LOC_19/A -0.00fF
C14249 NOR2X1_LOC_111/Y VDD 0.23fF
C14250 INVX1_LOC_18/A NOR2X1_LOC_467/A 0.42fF
C14251 NOR2X1_LOC_709/A INVX1_LOC_84/A 0.07fF
C14252 INVX1_LOC_136/A INVX1_LOC_4/A 0.20fF
C14253 NOR2X1_LOC_264/Y INVX1_LOC_19/A 0.22fF
C14254 NOR2X1_LOC_775/Y INVX1_LOC_37/A 0.03fF
C14255 NOR2X1_LOC_389/B INVX1_LOC_12/Y 0.10fF
C14256 INVX1_LOC_11/A INVX1_LOC_296/A 0.07fF
C14257 VDD NOR2X1_LOC_197/Y 0.24fF
C14258 INVX1_LOC_82/Y VDD 0.33fF
C14259 NOR2X1_LOC_667/A INVX1_LOC_285/A 0.13fF
C14260 NAND2X1_LOC_357/a_36_24# INVX1_LOC_32/A 0.06fF
C14261 NAND2X1_LOC_338/B INVX1_LOC_27/Y 0.03fF
C14262 NAND2X1_LOC_662/Y INVX1_LOC_117/Y 0.21fF
C14263 NOR2X1_LOC_667/A INVX1_LOC_265/Y 0.02fF
C14264 NOR2X1_LOC_525/Y INVX1_LOC_118/A 0.02fF
C14265 NAND2X1_LOC_397/a_36_24# NOR2X1_LOC_660/Y 0.01fF
C14266 INVX1_LOC_295/A NOR2X1_LOC_450/A 0.10fF
C14267 INVX1_LOC_30/Y INVX1_LOC_46/Y -0.01fF
C14268 NOR2X1_LOC_312/Y INVX1_LOC_118/A 0.38fF
C14269 NOR2X1_LOC_237/a_36_216# INVX1_LOC_19/Y 0.02fF
C14270 INVX1_LOC_162/A NOR2X1_LOC_89/A 0.07fF
C14271 NAND2X1_LOC_363/B INVX1_LOC_14/A 0.01fF
C14272 NOR2X1_LOC_606/Y NAND2X1_LOC_99/A 0.01fF
C14273 NOR2X1_LOC_163/Y INVX1_LOC_117/A 0.07fF
C14274 INVX1_LOC_83/A INVX1_LOC_291/A 0.10fF
C14275 NAND2X1_LOC_747/a_36_24# NAND2X1_LOC_782/B 0.01fF
C14276 NOR2X1_LOC_329/B NOR2X1_LOC_536/A 0.08fF
C14277 NAND2X1_LOC_348/A INVX1_LOC_12/Y 0.00fF
C14278 INVX1_LOC_6/A INVX1_LOC_76/A 1.00fF
C14279 NOR2X1_LOC_815/A NAND2X1_LOC_453/A 0.01fF
C14280 NOR2X1_LOC_318/B NAND2X1_LOC_843/a_36_24# 0.00fF
C14281 NOR2X1_LOC_791/Y NOR2X1_LOC_792/a_36_216# 0.03fF
C14282 NAND2X1_LOC_562/B INVX1_LOC_284/A 0.10fF
C14283 INVX1_LOC_190/A NOR2X1_LOC_435/A 0.01fF
C14284 NOR2X1_LOC_315/Y NOR2X1_LOC_89/A 0.15fF
C14285 NOR2X1_LOC_97/B NOR2X1_LOC_865/Y 0.00fF
C14286 INVX1_LOC_70/Y INVX1_LOC_304/A 0.02fF
C14287 INVX1_LOC_206/Y NOR2X1_LOC_357/Y 0.03fF
C14288 NOR2X1_LOC_74/Y INVX1_LOC_117/A 0.06fF
C14289 NOR2X1_LOC_97/B NOR2X1_LOC_243/B 0.04fF
C14290 INVX1_LOC_77/A NAND2X1_LOC_452/Y 0.03fF
C14291 NAND2X1_LOC_850/Y NAND2X1_LOC_74/B 0.07fF
C14292 INVX1_LOC_179/Y NOR2X1_LOC_633/A 0.04fF
C14293 NOR2X1_LOC_791/Y INVX1_LOC_14/A 0.09fF
C14294 INVX1_LOC_316/Y INVX1_LOC_19/A 0.03fF
C14295 NOR2X1_LOC_67/A INVX1_LOC_12/A 0.09fF
C14296 INVX1_LOC_166/A INVX1_LOC_195/A 0.03fF
C14297 NOR2X1_LOC_433/A INVX1_LOC_94/Y 0.01fF
C14298 INVX1_LOC_64/A NOR2X1_LOC_276/Y 0.14fF
C14299 INVX1_LOC_58/A INVX1_LOC_57/Y 0.09fF
C14300 INVX1_LOC_104/A INVX1_LOC_32/A 0.07fF
C14301 INVX1_LOC_77/A NOR2X1_LOC_307/Y 0.06fF
C14302 INVX1_LOC_186/A INVX1_LOC_37/A 0.04fF
C14303 NAND2X1_LOC_730/a_36_24# NOR2X1_LOC_829/A 0.00fF
C14304 INVX1_LOC_17/A NOR2X1_LOC_816/a_36_216# 0.00fF
C14305 NOR2X1_LOC_322/Y INVX1_LOC_54/A 0.10fF
C14306 NOR2X1_LOC_647/Y INVX1_LOC_25/A 0.44fF
C14307 NOR2X1_LOC_445/Y NOR2X1_LOC_334/Y 0.00fF
C14308 NOR2X1_LOC_192/A VDD 0.24fF
C14309 INVX1_LOC_28/A NAND2X1_LOC_798/B 0.13fF
C14310 INVX1_LOC_144/Y NOR2X1_LOC_48/B 0.05fF
C14311 INVX1_LOC_25/A INVX1_LOC_18/A 0.07fF
C14312 INVX1_LOC_222/Y INVX1_LOC_256/A 0.08fF
C14313 INVX1_LOC_278/Y INVX1_LOC_102/A 0.03fF
C14314 INVX1_LOC_21/A NAND2X1_LOC_803/B 0.05fF
C14315 INVX1_LOC_8/Y INVX1_LOC_26/Y 0.01fF
C14316 NAND2X1_LOC_192/B NOR2X1_LOC_348/Y 0.03fF
C14317 INPUT_0 INVX1_LOC_274/A -0.01fF
C14318 NOR2X1_LOC_721/a_36_216# NAND2X1_LOC_74/B 0.00fF
C14319 NOR2X1_LOC_34/B INVX1_LOC_31/A 0.03fF
C14320 INVX1_LOC_88/A NAND2X1_LOC_537/Y 0.00fF
C14321 NOR2X1_LOC_52/B INVX1_LOC_94/Y 0.55fF
C14322 INVX1_LOC_136/A INVX1_LOC_64/A 0.23fF
C14323 NOR2X1_LOC_252/Y NAND2X1_LOC_254/Y -0.00fF
C14324 NOR2X1_LOC_383/Y NOR2X1_LOC_178/a_36_216# 0.01fF
C14325 NOR2X1_LOC_45/B NAND2X1_LOC_446/a_36_24# 0.00fF
C14326 INVX1_LOC_246/A NOR2X1_LOC_173/Y 0.01fF
C14327 NOR2X1_LOC_20/Y INVX1_LOC_269/A 0.01fF
C14328 INVX1_LOC_21/A NOR2X1_LOC_590/A 0.19fF
C14329 INVX1_LOC_299/A INVX1_LOC_11/A 0.11fF
C14330 NOR2X1_LOC_264/Y INVX1_LOC_26/Y 0.66fF
C14331 INVX1_LOC_5/A INVX1_LOC_72/A 0.29fF
C14332 INVX1_LOC_232/Y NAND2X1_LOC_618/Y 0.03fF
C14333 INVX1_LOC_140/A INVX1_LOC_119/Y 0.07fF
C14334 INVX1_LOC_2/Y VDD 1.06fF
C14335 NOR2X1_LOC_538/B INVX1_LOC_11/A 0.01fF
C14336 NOR2X1_LOC_147/A INVX1_LOC_92/A 0.03fF
C14337 INVX1_LOC_16/A INVX1_LOC_47/Y 0.07fF
C14338 NOR2X1_LOC_475/a_36_216# NAND2X1_LOC_618/Y 0.00fF
C14339 NOR2X1_LOC_794/a_36_216# INVX1_LOC_53/A -0.01fF
C14340 NOR2X1_LOC_742/a_36_216# D_GATE_741 0.02fF
C14341 NAND2X1_LOC_638/Y NOR2X1_LOC_48/Y 0.01fF
C14342 INVX1_LOC_5/A INVX1_LOC_198/Y 0.05fF
C14343 NOR2X1_LOC_708/Y INVX1_LOC_301/A 0.03fF
C14344 NAND2X1_LOC_656/Y NAND2X1_LOC_792/B 0.01fF
C14345 NAND2X1_LOC_799/A NAND2X1_LOC_539/a_36_24# 0.02fF
C14346 NAND2X1_LOC_687/A VDD 0.00fF
C14347 D_INPUT_1 NAND2X1_LOC_276/Y 0.03fF
C14348 VDD INVX1_LOC_37/Y 0.21fF
C14349 NOR2X1_LOC_332/A NOR2X1_LOC_643/a_36_216# 0.01fF
C14350 NOR2X1_LOC_363/Y VDD 0.12fF
C14351 NOR2X1_LOC_78/A NOR2X1_LOC_640/Y 0.21fF
C14352 NOR2X1_LOC_689/Y NAND2X1_LOC_357/B 0.02fF
C14353 NOR2X1_LOC_15/Y INVX1_LOC_124/Y 0.01fF
C14354 NOR2X1_LOC_598/B NOR2X1_LOC_344/A 0.00fF
C14355 NOR2X1_LOC_787/a_36_216# NOR2X1_LOC_794/B 0.02fF
C14356 NOR2X1_LOC_61/B NOR2X1_LOC_68/A 0.02fF
C14357 NOR2X1_LOC_356/A INVX1_LOC_99/A 0.01fF
C14358 NOR2X1_LOC_209/Y NOR2X1_LOC_727/B 0.02fF
C14359 NOR2X1_LOC_166/Y NOR2X1_LOC_89/A 0.01fF
C14360 INVX1_LOC_14/A INVX1_LOC_30/A 0.39fF
C14361 INVX1_LOC_181/Y NAND2X1_LOC_474/Y 0.32fF
C14362 NOR2X1_LOC_272/Y INVX1_LOC_24/A 0.16fF
C14363 INVX1_LOC_150/Y NAND2X1_LOC_337/a_36_24# 0.00fF
C14364 INVX1_LOC_225/A NOR2X1_LOC_717/A 0.10fF
C14365 NAND2X1_LOC_762/a_36_24# INVX1_LOC_1/A 0.01fF
C14366 NOR2X1_LOC_613/Y NOR2X1_LOC_238/Y 0.01fF
C14367 INVX1_LOC_1/A INVX1_LOC_18/A 0.31fF
C14368 INVX1_LOC_49/A INVX1_LOC_50/Y 0.04fF
C14369 NOR2X1_LOC_658/Y NOR2X1_LOC_215/a_36_216# 0.01fF
C14370 NAND2X1_LOC_4/a_36_24# INVX1_LOC_3/A 0.01fF
C14371 VDD NOR2X1_LOC_866/B 0.09fF
C14372 NAND2X1_LOC_860/A INVX1_LOC_168/A 0.04fF
C14373 INVX1_LOC_25/A INVX1_LOC_34/Y 0.41fF
C14374 INVX1_LOC_135/A NOR2X1_LOC_38/B 0.68fF
C14375 NAND2X1_LOC_287/B INVX1_LOC_118/A 0.18fF
C14376 INVX1_LOC_35/A NOR2X1_LOC_310/Y 0.01fF
C14377 NAND2X1_LOC_729/Y NOR2X1_LOC_536/Y 0.05fF
C14378 NAND2X1_LOC_714/B NAND2X1_LOC_593/Y 0.01fF
C14379 INVX1_LOC_50/A NAND2X1_LOC_862/A 0.01fF
C14380 INVX1_LOC_278/A NOR2X1_LOC_709/A 0.19fF
C14381 NAND2X1_LOC_725/A NAND2X1_LOC_357/B 0.31fF
C14382 INVX1_LOC_34/A INVX1_LOC_306/Y 0.07fF
C14383 NAND2X1_LOC_9/Y NOR2X1_LOC_721/A 0.05fF
C14384 INVX1_LOC_131/Y INVX1_LOC_76/A 0.10fF
C14385 VDD INVX1_LOC_307/Y 0.18fF
C14386 NAND2X1_LOC_380/a_36_24# NOR2X1_LOC_460/Y 0.00fF
C14387 NOR2X1_LOC_74/A INVX1_LOC_99/A 0.22fF
C14388 NAND2X1_LOC_67/Y NOR2X1_LOC_208/Y 0.01fF
C14389 INVX1_LOC_36/A NOR2X1_LOC_331/Y 0.00fF
C14390 INVX1_LOC_291/A INVX1_LOC_46/A 0.07fF
C14391 NOR2X1_LOC_816/A INVX1_LOC_72/A 0.01fF
C14392 NOR2X1_LOC_322/Y NOR2X1_LOC_48/B 0.12fF
C14393 NOR2X1_LOC_234/Y NOR2X1_LOC_291/Y -0.03fF
C14394 NOR2X1_LOC_719/B INVX1_LOC_16/Y 0.16fF
C14395 NAND2X1_LOC_362/a_36_24# NOR2X1_LOC_852/Y 0.01fF
C14396 NAND2X1_LOC_326/A NOR2X1_LOC_577/Y 0.35fF
C14397 NAND2X1_LOC_588/B INVX1_LOC_174/A 0.01fF
C14398 VDD NOR2X1_LOC_608/Y 0.37fF
C14399 NAND2X1_LOC_436/a_36_24# NAND2X1_LOC_453/A 0.01fF
C14400 INVX1_LOC_17/A INVX1_LOC_314/Y 0.07fF
C14401 NOR2X1_LOC_590/A NAND2X1_LOC_354/Y 0.06fF
C14402 INVX1_LOC_207/A NAND2X1_LOC_493/Y 0.06fF
C14403 INVX1_LOC_215/Y NOR2X1_LOC_512/Y 0.00fF
C14404 NOR2X1_LOC_561/Y INVX1_LOC_270/A 0.17fF
C14405 INVX1_LOC_5/A NOR2X1_LOC_537/Y 0.09fF
C14406 NAND2X1_LOC_685/a_36_24# INVX1_LOC_92/A 0.00fF
C14407 NAND2X1_LOC_842/B INVX1_LOC_78/A 0.05fF
C14408 INVX1_LOC_45/A NAND2X1_LOC_154/Y 0.08fF
C14409 INVX1_LOC_299/A NOR2X1_LOC_593/Y 0.56fF
C14410 INVX1_LOC_233/A NAND2X1_LOC_860/Y 0.03fF
C14411 INVX1_LOC_5/A NAND2X1_LOC_338/B 0.08fF
C14412 NOR2X1_LOC_750/Y NOR2X1_LOC_789/A 0.09fF
C14413 INVX1_LOC_269/A INVX1_LOC_33/A 0.47fF
C14414 NOR2X1_LOC_588/A NOR2X1_LOC_1/Y 0.02fF
C14415 NOR2X1_LOC_719/B NAND2X1_LOC_205/A 0.05fF
C14416 NOR2X1_LOC_13/Y NOR2X1_LOC_45/Y 0.01fF
C14417 INVX1_LOC_6/A INVX1_LOC_127/Y 0.00fF
C14418 INVX1_LOC_7/A NOR2X1_LOC_416/A 0.08fF
C14419 D_INPUT_4 NAND2X1_LOC_470/B 0.00fF
C14420 VDD NOR2X1_LOC_485/Y 0.23fF
C14421 INVX1_LOC_161/Y INVX1_LOC_155/A 0.01fF
C14422 INPUT_1 NOR2X1_LOC_72/Y 0.01fF
C14423 NOR2X1_LOC_384/Y INVX1_LOC_18/A 0.07fF
C14424 INVX1_LOC_30/A NOR2X1_LOC_522/Y 0.18fF
C14425 INVX1_LOC_11/A NAND2X1_LOC_157/a_36_24# 0.00fF
C14426 INVX1_LOC_24/A NOR2X1_LOC_761/Y 0.26fF
C14427 NOR2X1_LOC_65/B NAND2X1_LOC_842/B 0.02fF
C14428 INVX1_LOC_206/Y INVX1_LOC_32/A 0.03fF
C14429 NOR2X1_LOC_391/B NOR2X1_LOC_38/B 0.02fF
C14430 INVX1_LOC_24/A NOR2X1_LOC_336/B 0.04fF
C14431 INVX1_LOC_11/A INVX1_LOC_162/A 0.43fF
C14432 NAND2X1_LOC_842/a_36_24# INVX1_LOC_26/A 0.00fF
C14433 NOR2X1_LOC_848/Y NOR2X1_LOC_844/A 0.00fF
C14434 INVX1_LOC_28/A NAND2X1_LOC_211/a_36_24# 0.01fF
C14435 INVX1_LOC_11/A NOR2X1_LOC_350/a_36_216# 0.00fF
C14436 INVX1_LOC_286/Y NOR2X1_LOC_753/a_36_216# 0.00fF
C14437 NAND2X1_LOC_84/Y INVX1_LOC_30/A 0.00fF
C14438 INVX1_LOC_1/A INVX1_LOC_34/Y 0.10fF
C14439 NAND2X1_LOC_534/a_36_24# NAND2X1_LOC_537/Y 0.00fF
C14440 INVX1_LOC_11/A NOR2X1_LOC_315/Y 0.07fF
C14441 INVX1_LOC_27/A NOR2X1_LOC_210/B 0.16fF
C14442 NOR2X1_LOC_479/B INVX1_LOC_235/Y 0.97fF
C14443 NAND2X1_LOC_728/Y NAND2X1_LOC_729/Y 0.05fF
C14444 INVX1_LOC_24/A NAND2X1_LOC_364/A 0.07fF
C14445 NOR2X1_LOC_160/B NOR2X1_LOC_392/B 0.10fF
C14446 NOR2X1_LOC_508/a_36_216# NOR2X1_LOC_510/B 0.01fF
C14447 NOR2X1_LOC_248/Y INVX1_LOC_49/A 0.05fF
C14448 INVX1_LOC_233/A NAND2X1_LOC_861/Y 0.02fF
C14449 NOR2X1_LOC_788/B INVX1_LOC_53/A 0.00fF
C14450 INVX1_LOC_116/A NOR2X1_LOC_360/Y 0.05fF
C14451 INVX1_LOC_172/A NOR2X1_LOC_384/Y 0.03fF
C14452 NOR2X1_LOC_130/Y NOR2X1_LOC_392/Y -0.03fF
C14453 NOR2X1_LOC_558/A INVX1_LOC_12/A 0.01fF
C14454 NAND2X1_LOC_11/a_36_24# NAND2X1_LOC_30/Y 0.00fF
C14455 NOR2X1_LOC_541/Y NOR2X1_LOC_175/A 0.01fF
C14456 NAND2X1_LOC_63/Y INVX1_LOC_129/Y 0.03fF
C14457 INVX1_LOC_45/A INVX1_LOC_63/Y 0.03fF
C14458 INVX1_LOC_54/Y INVX1_LOC_150/Y 0.01fF
C14459 NAND2X1_LOC_736/Y NAND2X1_LOC_722/a_36_24# 0.01fF
C14460 INVX1_LOC_58/A NOR2X1_LOC_163/Y -0.00fF
C14461 NOR2X1_LOC_657/Y INVX1_LOC_34/A 0.00fF
C14462 NOR2X1_LOC_467/a_36_216# NAND2X1_LOC_149/Y 0.01fF
C14463 INVX1_LOC_21/A INVX1_LOC_227/A 0.18fF
C14464 INVX1_LOC_9/A INVX1_LOC_63/A 0.13fF
C14465 NAND2X1_LOC_711/B NAND2X1_LOC_710/a_36_24# 0.02fF
C14466 NAND2X1_LOC_149/Y NOR2X1_LOC_424/a_36_216# 0.00fF
C14467 INVX1_LOC_21/A NOR2X1_LOC_763/Y 0.04fF
C14468 NAND2X1_LOC_754/a_36_24# INVX1_LOC_269/A 0.00fF
C14469 NAND2X1_LOC_803/B INVX1_LOC_248/A 0.01fF
C14470 NAND2X1_LOC_361/Y NOR2X1_LOC_360/Y 0.03fF
C14471 NOR2X1_LOC_139/Y NAND2X1_LOC_454/Y 0.00fF
C14472 NAND2X1_LOC_350/A INVX1_LOC_144/Y -0.08fF
C14473 NAND2X1_LOC_364/A NOR2X1_LOC_557/Y 0.01fF
C14474 NAND2X1_LOC_354/Y NAND2X1_LOC_354/B 0.03fF
C14475 INVX1_LOC_5/A INVX1_LOC_313/Y 0.07fF
C14476 NOR2X1_LOC_524/Y NOR2X1_LOC_52/B 0.01fF
C14477 NAND2X1_LOC_581/Y D_INPUT_7 0.01fF
C14478 INVX1_LOC_214/A NOR2X1_LOC_590/A 0.03fF
C14479 INVX1_LOC_75/A INVX1_LOC_58/Y 0.00fF
C14480 NOR2X1_LOC_667/A NOR2X1_LOC_590/A 0.21fF
C14481 INVX1_LOC_30/A NOR2X1_LOC_612/B 0.20fF
C14482 INVX1_LOC_45/A NOR2X1_LOC_175/A 0.03fF
C14483 NOR2X1_LOC_559/B INVX1_LOC_49/A 0.03fF
C14484 INVX1_LOC_279/Y NOR2X1_LOC_78/B 0.04fF
C14485 INVX1_LOC_248/A NOR2X1_LOC_590/A 0.00fF
C14486 NOR2X1_LOC_653/B INVX1_LOC_90/A 0.05fF
C14487 NAND2X1_LOC_733/A NAND2X1_LOC_717/Y 0.02fF
C14488 INVX1_LOC_91/A NOR2X1_LOC_318/A 0.08fF
C14489 NOR2X1_LOC_89/A NAND2X1_LOC_93/a_36_24# 0.00fF
C14490 NOR2X1_LOC_389/A NOR2X1_LOC_366/B 0.04fF
C14491 INVX1_LOC_27/A NOR2X1_LOC_72/a_36_216# 0.01fF
C14492 NAND2X1_LOC_860/A NOR2X1_LOC_83/a_36_216# 0.01fF
C14493 INVX1_LOC_27/A INVX1_LOC_20/Y 0.03fF
C14494 INVX1_LOC_247/A INVX1_LOC_271/Y 0.05fF
C14495 NAND2X1_LOC_468/B NAND2X1_LOC_454/Y 0.02fF
C14496 NOR2X1_LOC_388/Y NOR2X1_LOC_596/A 0.14fF
C14497 NAND2X1_LOC_288/A NAND2X1_LOC_286/a_36_24# 0.04fF
C14498 NAND2X1_LOC_9/Y INVX1_LOC_158/Y 0.01fF
C14499 NAND2X1_LOC_623/B NOR2X1_LOC_693/Y 0.00fF
C14500 NOR2X1_LOC_92/Y NOR2X1_LOC_246/A 0.07fF
C14501 INVX1_LOC_63/Y INVX1_LOC_71/A 0.07fF
C14502 NOR2X1_LOC_15/Y D_INPUT_0 0.22fF
C14503 INVX1_LOC_125/Y INVX1_LOC_57/A 0.07fF
C14504 NOR2X1_LOC_114/a_36_216# NOR2X1_LOC_114/Y 0.03fF
C14505 NOR2X1_LOC_100/a_36_216# NOR2X1_LOC_843/B 0.01fF
C14506 NOR2X1_LOC_92/Y NAND2X1_LOC_551/A 0.04fF
C14507 NOR2X1_LOC_865/A NOR2X1_LOC_861/Y 0.03fF
C14508 INVX1_LOC_24/Y NOR2X1_LOC_174/B 0.47fF
C14509 NOR2X1_LOC_449/A NAND2X1_LOC_469/B 0.73fF
C14510 INVX1_LOC_136/A NAND2X1_LOC_850/Y 0.07fF
C14511 NOR2X1_LOC_433/A INVX1_LOC_162/A 0.01fF
C14512 INVX1_LOC_50/A NOR2X1_LOC_595/Y 0.02fF
C14513 NAND2X1_LOC_364/A INVX1_LOC_143/A 0.02fF
C14514 NOR2X1_LOC_67/A INVX1_LOC_217/A 0.10fF
C14515 NAND2X1_LOC_785/A INVX1_LOC_24/A 0.07fF
C14516 NAND2X1_LOC_465/A INVX1_LOC_23/Y 0.00fF
C14517 NOR2X1_LOC_773/Y INVX1_LOC_72/A 0.08fF
C14518 NOR2X1_LOC_381/Y INPUT_1 0.03fF
C14519 NOR2X1_LOC_167/Y NOR2X1_LOC_109/Y 0.12fF
C14520 INVX1_LOC_84/A INVX1_LOC_294/A 0.05fF
C14521 NOR2X1_LOC_817/a_36_216# INVX1_LOC_89/A 0.02fF
C14522 NOR2X1_LOC_682/Y INVX1_LOC_273/A 0.30fF
C14523 INPUT_0 INVX1_LOC_306/Y 0.07fF
C14524 NOR2X1_LOC_178/Y INVX1_LOC_6/A 0.16fF
C14525 INVX1_LOC_49/A NOR2X1_LOC_6/B 0.03fF
C14526 NOR2X1_LOC_627/Y INVX1_LOC_24/A 0.02fF
C14527 NOR2X1_LOC_262/Y NOR2X1_LOC_709/A 0.06fF
C14528 NOR2X1_LOC_226/A NAND2X1_LOC_356/a_36_24# 0.00fF
C14529 NOR2X1_LOC_831/B INVX1_LOC_29/A 0.11fF
C14530 INVX1_LOC_304/Y NOR2X1_LOC_753/Y 0.01fF
C14531 NOR2X1_LOC_78/A NOR2X1_LOC_247/Y 0.05fF
C14532 NOR2X1_LOC_590/A NOR2X1_LOC_565/B 0.01fF
C14533 NOR2X1_LOC_763/Y NOR2X1_LOC_428/Y 0.14fF
C14534 INVX1_LOC_91/A NOR2X1_LOC_678/A 0.03fF
C14535 NOR2X1_LOC_653/Y NOR2X1_LOC_662/A 0.03fF
C14536 INVX1_LOC_280/A NOR2X1_LOC_38/B 0.40fF
C14537 INVX1_LOC_91/A INVX1_LOC_295/Y 0.56fF
C14538 NOR2X1_LOC_718/a_36_216# INVX1_LOC_113/Y 0.00fF
C14539 NOR2X1_LOC_194/a_36_216# INVX1_LOC_22/A 0.02fF
C14540 INVX1_LOC_290/A NAND2X1_LOC_16/Y 0.02fF
C14541 INVX1_LOC_90/A NAND2X1_LOC_550/A 0.07fF
C14542 INVX1_LOC_270/A INVX1_LOC_76/A 0.01fF
C14543 NAND2X1_LOC_642/Y NOR2X1_LOC_717/A 0.00fF
C14544 INVX1_LOC_36/A NOR2X1_LOC_561/Y 0.16fF
C14545 INVX1_LOC_39/A NOR2X1_LOC_391/Y 0.00fF
C14546 INVX1_LOC_36/A INVX1_LOC_7/A 0.02fF
C14547 INVX1_LOC_295/A NOR2X1_LOC_389/A 0.03fF
C14548 INVX1_LOC_17/A NAND2X1_LOC_123/Y 0.01fF
C14549 INVX1_LOC_90/A NOR2X1_LOC_160/B 0.21fF
C14550 NAND2X1_LOC_308/Y NAND2X1_LOC_357/B 0.01fF
C14551 INVX1_LOC_239/A NAND2X1_LOC_622/B 0.12fF
C14552 NOR2X1_LOC_666/Y INVX1_LOC_42/Y 0.02fF
C14553 VDD NOR2X1_LOC_809/A 0.24fF
C14554 INVX1_LOC_256/A NOR2X1_LOC_329/B 0.10fF
C14555 NOR2X1_LOC_389/B NOR2X1_LOC_160/B 0.30fF
C14556 NAND2X1_LOC_347/B NOR2X1_LOC_83/Y 0.20fF
C14557 NOR2X1_LOC_137/A INVX1_LOC_30/A 0.10fF
C14558 NOR2X1_LOC_804/B INVX1_LOC_179/Y 0.02fF
C14559 NOR2X1_LOC_596/A NAND2X1_LOC_479/Y 0.03fF
C14560 NOR2X1_LOC_52/B NOR2X1_LOC_315/Y 0.11fF
C14561 VDD INVX1_LOC_29/Y 0.87fF
C14562 INVX1_LOC_214/A NAND2X1_LOC_354/B 0.01fF
C14563 INVX1_LOC_119/Y INVX1_LOC_42/A 0.14fF
C14564 INVX1_LOC_71/A NOR2X1_LOC_188/a_36_216# 0.00fF
C14565 INVX1_LOC_77/A INVX1_LOC_1/Y 0.07fF
C14566 NOR2X1_LOC_75/Y INVX1_LOC_75/A 0.03fF
C14567 INVX1_LOC_181/Y INVX1_LOC_10/A 0.16fF
C14568 INVX1_LOC_30/A NOR2X1_LOC_588/a_36_216# 0.01fF
C14569 NOR2X1_LOC_716/B INVX1_LOC_25/Y 0.22fF
C14570 NOR2X1_LOC_705/B NOR2X1_LOC_706/A 0.03fF
C14571 NOR2X1_LOC_208/Y NOR2X1_LOC_561/Y 0.10fF
C14572 NAND2X1_LOC_656/Y NOR2X1_LOC_359/Y -0.02fF
C14573 NOR2X1_LOC_160/B NAND2X1_LOC_348/A 0.13fF
C14574 INVX1_LOC_59/A NOR2X1_LOC_45/B 0.12fF
C14575 INVX1_LOC_271/Y NOR2X1_LOC_676/Y 0.01fF
C14576 INVX1_LOC_76/A NOR2X1_LOC_109/Y 0.14fF
C14577 NOR2X1_LOC_861/Y INVX1_LOC_63/A 0.07fF
C14578 NOR2X1_LOC_379/Y INVX1_LOC_174/Y 0.01fF
C14579 NOR2X1_LOC_516/B NOR2X1_LOC_147/B 0.18fF
C14580 NAND2X1_LOC_660/A NAND2X1_LOC_655/a_36_24# 0.01fF
C14581 INVX1_LOC_8/A INVX1_LOC_56/Y 0.04fF
C14582 NOR2X1_LOC_370/a_36_216# INVX1_LOC_71/A 0.00fF
C14583 NAND2X1_LOC_405/a_36_24# NOR2X1_LOC_109/Y 0.01fF
C14584 NOR2X1_LOC_15/Y NOR2X1_LOC_191/a_36_216# 0.00fF
C14585 NOR2X1_LOC_52/B INVX1_LOC_52/A 0.07fF
C14586 INVX1_LOC_304/Y NOR2X1_LOC_488/a_36_216# 0.00fF
C14587 INVX1_LOC_41/A INVX1_LOC_13/A 0.01fF
C14588 INVX1_LOC_295/A NOR2X1_LOC_596/A 0.04fF
C14589 INVX1_LOC_201/Y INVX1_LOC_13/A 0.58fF
C14590 NOR2X1_LOC_504/Y NAND2X1_LOC_852/Y 0.08fF
C14591 INVX1_LOC_276/A INVX1_LOC_214/Y 0.02fF
C14592 NOR2X1_LOC_753/Y NAND2X1_LOC_808/A 0.07fF
C14593 INVX1_LOC_72/A INVX1_LOC_140/A 0.10fF
C14594 NAND2X1_LOC_182/A NAND2X1_LOC_564/B 0.01fF
C14595 NOR2X1_LOC_590/A INVX1_LOC_311/A 0.79fF
C14596 INVX1_LOC_17/A NOR2X1_LOC_557/A 0.07fF
C14597 NOR2X1_LOC_248/A INVX1_LOC_285/A 0.01fF
C14598 NOR2X1_LOC_300/Y INVX1_LOC_22/A 0.01fF
C14599 INVX1_LOC_298/Y NOR2X1_LOC_831/B 0.01fF
C14600 NAND2X1_LOC_338/B NAND2X1_LOC_9/a_36_24# 0.00fF
C14601 NAND2X1_LOC_782/B NOR2X1_LOC_685/Y 0.02fF
C14602 INVX1_LOC_35/A NOR2X1_LOC_536/A 2.94fF
C14603 INVX1_LOC_21/A NAND2X1_LOC_650/B 0.07fF
C14604 INVX1_LOC_124/A INVX1_LOC_1/Y 0.18fF
C14605 INVX1_LOC_201/Y NAND2X1_LOC_14/a_36_24# 0.01fF
C14606 NOR2X1_LOC_334/Y INVX1_LOC_84/A 0.07fF
C14607 INVX1_LOC_284/A INVX1_LOC_42/A 0.24fF
C14608 INVX1_LOC_72/A NAND2X1_LOC_463/B 0.00fF
C14609 INVX1_LOC_80/A NOR2X1_LOC_516/Y 0.06fF
C14610 NAND2X1_LOC_325/Y NAND2X1_LOC_808/A 0.14fF
C14611 INVX1_LOC_78/A INVX1_LOC_119/Y 0.04fF
C14612 NOR2X1_LOC_561/Y NOR2X1_LOC_309/Y 0.02fF
C14613 INVX1_LOC_136/A INVX1_LOC_282/A 0.36fF
C14614 NOR2X1_LOC_474/A NAND2X1_LOC_624/A 0.01fF
C14615 NAND2X1_LOC_796/B INVX1_LOC_37/A 0.03fF
C14616 NOR2X1_LOC_454/Y INVX1_LOC_139/A 0.01fF
C14617 NAND2X1_LOC_785/A NAND2X1_LOC_552/a_36_24# 0.00fF
C14618 INVX1_LOC_2/A INVX1_LOC_30/Y 0.03fF
C14619 INVX1_LOC_41/A NOR2X1_LOC_174/B 0.01fF
C14620 INVX1_LOC_209/Y NOR2X1_LOC_597/A 0.01fF
C14621 NOR2X1_LOC_452/A INVX1_LOC_92/A 0.03fF
C14622 INVX1_LOC_18/A NOR2X1_LOC_188/A 0.17fF
C14623 INVX1_LOC_36/A NAND2X1_LOC_251/a_36_24# 0.00fF
C14624 INVX1_LOC_58/A INVX1_LOC_179/A 0.02fF
C14625 INVX1_LOC_135/A NOR2X1_LOC_844/A 0.01fF
C14626 NOR2X1_LOC_632/Y NOR2X1_LOC_78/B 0.03fF
C14627 NOR2X1_LOC_551/B INVX1_LOC_196/Y 0.06fF
C14628 NOR2X1_LOC_226/A INVX1_LOC_30/Y 0.01fF
C14629 INVX1_LOC_35/A NOR2X1_LOC_655/Y 0.03fF
C14630 NOR2X1_LOC_15/Y NOR2X1_LOC_266/B 0.00fF
C14631 NAND2X1_LOC_162/B INVX1_LOC_75/A 0.04fF
C14632 INVX1_LOC_18/A NOR2X1_LOC_548/B 0.10fF
C14633 NOR2X1_LOC_246/A NAND2X1_LOC_477/A 0.10fF
C14634 D_INPUT_0 NAND2X1_LOC_141/A 0.02fF
C14635 INVX1_LOC_35/A NAND2X1_LOC_93/B 0.03fF
C14636 NAND2X1_LOC_252/a_36_24# NOR2X1_LOC_727/B 0.00fF
C14637 NOR2X1_LOC_328/Y INVX1_LOC_16/A 0.07fF
C14638 NOR2X1_LOC_469/a_36_216# NAND2X1_LOC_650/B 0.01fF
C14639 NOR2X1_LOC_775/Y INVX1_LOC_310/Y 0.02fF
C14640 NOR2X1_LOC_6/B INPUT_1 0.19fF
C14641 INVX1_LOC_213/Y INVX1_LOC_196/Y 0.29fF
C14642 NAND2X1_LOC_817/a_36_24# NOR2X1_LOC_660/Y -0.00fF
C14643 NOR2X1_LOC_332/A NOR2X1_LOC_537/Y 0.08fF
C14644 NOR2X1_LOC_844/A NOR2X1_LOC_560/A 0.36fF
C14645 NAND2X1_LOC_551/A NAND2X1_LOC_477/A 0.00fF
C14646 NOR2X1_LOC_716/B INVX1_LOC_75/A 0.07fF
C14647 NOR2X1_LOC_32/B INVX1_LOC_260/Y 0.05fF
C14648 INVX1_LOC_35/A NAND2X1_LOC_425/Y 0.12fF
C14649 INVX1_LOC_57/A NOR2X1_LOC_653/Y 0.49fF
C14650 NOR2X1_LOC_383/Y INVX1_LOC_53/Y 0.07fF
C14651 NOR2X1_LOC_667/a_36_216# INVX1_LOC_76/A 0.00fF
C14652 NAND2X1_LOC_352/a_36_24# NAND2X1_LOC_287/B 0.00fF
C14653 NOR2X1_LOC_15/Y NAND2X1_LOC_848/A 0.12fF
C14654 NOR2X1_LOC_155/A INVX1_LOC_213/A 0.06fF
C14655 NAND2X1_LOC_181/Y NOR2X1_LOC_71/Y 0.02fF
C14656 D_INPUT_0 INVX1_LOC_226/A 0.03fF
C14657 INVX1_LOC_178/A NOR2X1_LOC_506/Y 0.29fF
C14658 INVX1_LOC_243/Y INVX1_LOC_19/A 0.02fF
C14659 NOR2X1_LOC_219/Y NOR2X1_LOC_366/Y 0.15fF
C14660 INVX1_LOC_49/A NAND2X1_LOC_328/a_36_24# 0.00fF
C14661 INVX1_LOC_295/A INVX1_LOC_189/Y 0.04fF
C14662 INVX1_LOC_18/A NOR2X1_LOC_43/Y 0.05fF
C14663 INVX1_LOC_90/A NOR2X1_LOC_213/a_36_216# 0.02fF
C14664 NOR2X1_LOC_68/A NAND2X1_LOC_655/A 0.07fF
C14665 INVX1_LOC_36/A NOR2X1_LOC_824/Y 0.03fF
C14666 INVX1_LOC_34/A NOR2X1_LOC_74/A 0.11fF
C14667 INVX1_LOC_11/A NAND2X1_LOC_96/A 0.09fF
C14668 INVX1_LOC_35/A NOR2X1_LOC_649/B 0.12fF
C14669 INVX1_LOC_57/A INVX1_LOC_19/A 0.37fF
C14670 NOR2X1_LOC_720/A NAND2X1_LOC_74/B 0.01fF
C14671 INVX1_LOC_35/A INVX1_LOC_3/A 0.15fF
C14672 NOR2X1_LOC_89/A NAND2X1_LOC_99/A 0.03fF
C14673 NOR2X1_LOC_334/Y INVX1_LOC_15/A 0.07fF
C14674 NAND2X1_LOC_654/B NAND2X1_LOC_451/Y 0.05fF
C14675 NAND2X1_LOC_374/Y NOR2X1_LOC_497/Y 0.06fF
C14676 INVX1_LOC_34/A NOR2X1_LOC_9/Y 0.07fF
C14677 INVX1_LOC_36/A INVX1_LOC_76/A 0.64fF
C14678 INVX1_LOC_24/A NOR2X1_LOC_405/A 0.04fF
C14679 INVX1_LOC_77/A NOR2X1_LOC_318/B 1.11fF
C14680 INVX1_LOC_49/A INVX1_LOC_96/A 0.02fF
C14681 NOR2X1_LOC_78/B NOR2X1_LOC_135/Y 0.04fF
C14682 INVX1_LOC_286/Y NOR2X1_LOC_111/A 0.10fF
C14683 NOR2X1_LOC_160/B NOR2X1_LOC_561/A 0.01fF
C14684 NOR2X1_LOC_68/A NOR2X1_LOC_683/Y 0.02fF
C14685 NOR2X1_LOC_13/Y NAND2X1_LOC_642/Y 0.01fF
C14686 NAND2X1_LOC_550/A INVX1_LOC_38/A 0.15fF
C14687 INVX1_LOC_11/A NAND2X1_LOC_427/a_36_24# 0.00fF
C14688 NOR2X1_LOC_335/A INVX1_LOC_91/A 0.03fF
C14689 NOR2X1_LOC_309/Y NOR2X1_LOC_167/Y 0.05fF
C14690 NOR2X1_LOC_160/B INVX1_LOC_38/A 0.10fF
C14691 NOR2X1_LOC_92/Y INVX1_LOC_260/A 0.03fF
C14692 INVX1_LOC_77/A INVX1_LOC_93/Y 0.15fF
C14693 NOR2X1_LOC_391/A INVX1_LOC_89/A 0.03fF
C14694 NOR2X1_LOC_790/B INVX1_LOC_29/A 0.07fF
C14695 NOR2X1_LOC_15/Y INVX1_LOC_46/Y 0.02fF
C14696 NAND2X1_LOC_231/Y NOR2X1_LOC_74/A 0.97fF
C14697 INVX1_LOC_27/A NAND2X1_LOC_73/a_36_24# 0.00fF
C14698 INVX1_LOC_286/Y NOR2X1_LOC_694/Y 0.11fF
C14699 INVX1_LOC_269/A INVX1_LOC_241/Y 0.02fF
C14700 INVX1_LOC_271/Y NOR2X1_LOC_465/Y 0.02fF
C14701 INVX1_LOC_24/A NOR2X1_LOC_682/a_36_216# 0.01fF
C14702 INVX1_LOC_145/A INVX1_LOC_76/A 0.05fF
C14703 NOR2X1_LOC_557/Y NOR2X1_LOC_405/A 0.20fF
C14704 NOR2X1_LOC_373/Y NOR2X1_LOC_76/A 0.00fF
C14705 INVX1_LOC_24/A NOR2X1_LOC_857/A 0.07fF
C14706 NOR2X1_LOC_208/Y INVX1_LOC_76/A 0.02fF
C14707 INVX1_LOC_123/A NOR2X1_LOC_709/A 0.02fF
C14708 NOR2X1_LOC_516/B NAND2X1_LOC_348/A 0.51fF
C14709 NAND2X1_LOC_464/B INVX1_LOC_15/A 0.07fF
C14710 INVX1_LOC_33/A NOR2X1_LOC_275/A 0.01fF
C14711 NAND2X1_LOC_567/Y INVX1_LOC_20/A 0.12fF
C14712 NOR2X1_LOC_596/A INVX1_LOC_139/Y 0.04fF
C14713 NOR2X1_LOC_286/Y NOR2X1_LOC_445/B 0.03fF
C14714 INVX1_LOC_124/A NOR2X1_LOC_318/B 0.13fF
C14715 INVX1_LOC_164/Y INVX1_LOC_286/A 0.03fF
C14716 INVX1_LOC_77/A INVX1_LOC_139/A 0.03fF
C14717 NOR2X1_LOC_434/Y NOR2X1_LOC_633/A 0.00fF
C14718 INVX1_LOC_50/Y NAND2X1_LOC_63/Y 0.10fF
C14719 INVX1_LOC_78/A NOR2X1_LOC_134/a_36_216# 0.00fF
C14720 NOR2X1_LOC_655/B NOR2X1_LOC_355/B 0.05fF
C14721 NOR2X1_LOC_92/Y NAND2X1_LOC_489/Y 0.03fF
C14722 INVX1_LOC_213/A NOR2X1_LOC_833/B 0.17fF
C14723 INVX1_LOC_246/A NAND2X1_LOC_798/B 0.02fF
C14724 NOR2X1_LOC_744/Y INVX1_LOC_33/Y 0.01fF
C14725 NOR2X1_LOC_785/A NOR2X1_LOC_634/A 0.04fF
C14726 NOR2X1_LOC_470/A INVX1_LOC_75/A 0.52fF
C14727 NOR2X1_LOC_802/A INVX1_LOC_65/A 0.10fF
C14728 NOR2X1_LOC_724/a_36_216# NOR2X1_LOC_78/A 0.00fF
C14729 NOR2X1_LOC_172/Y NAND2X1_LOC_211/Y 0.02fF
C14730 NOR2X1_LOC_860/B NOR2X1_LOC_859/Y 0.00fF
C14731 NOR2X1_LOC_717/B NOR2X1_LOC_439/B 0.03fF
C14732 INVX1_LOC_124/A INVX1_LOC_93/Y 0.04fF
C14733 NOR2X1_LOC_523/A NOR2X1_LOC_814/A 0.04fF
C14734 NOR2X1_LOC_596/A INVX1_LOC_10/Y 0.02fF
C14735 NOR2X1_LOC_717/B INVX1_LOC_75/A 0.03fF
C14736 INVX1_LOC_143/A NOR2X1_LOC_405/A 0.07fF
C14737 NOR2X1_LOC_309/Y INVX1_LOC_76/A 0.01fF
C14738 NOR2X1_LOC_763/Y NAND2X1_LOC_51/B 0.00fF
C14739 NOR2X1_LOC_764/Y D_INPUT_4 0.02fF
C14740 INVX1_LOC_21/A NOR2X1_LOC_67/Y 0.07fF
C14741 INVX1_LOC_33/A INVX1_LOC_12/Y 1.19fF
C14742 NAND2X1_LOC_19/a_36_24# NOR2X1_LOC_814/A 0.01fF
C14743 NOR2X1_LOC_220/A NOR2X1_LOC_552/A 0.10fF
C14744 NOR2X1_LOC_226/A NOR2X1_LOC_124/A 0.01fF
C14745 NOR2X1_LOC_665/Y INVX1_LOC_4/A 0.07fF
C14746 NAND2X1_LOC_563/Y INVX1_LOC_178/Y 0.03fF
C14747 INVX1_LOC_90/A NOR2X1_LOC_706/A 0.35fF
C14748 INVX1_LOC_60/Y VDD 0.49fF
C14749 INVX1_LOC_26/Y INVX1_LOC_57/A 0.10fF
C14750 INVX1_LOC_35/A NAND2X1_LOC_470/B 0.07fF
C14751 NAND2X1_LOC_555/Y NAND2X1_LOC_657/a_36_24# 0.01fF
C14752 INVX1_LOC_58/A NOR2X1_LOC_693/Y 0.07fF
C14753 INVX1_LOC_25/A NOR2X1_LOC_647/A 0.05fF
C14754 NOR2X1_LOC_250/Y INVX1_LOC_49/Y 0.23fF
C14755 INVX1_LOC_83/A NOR2X1_LOC_147/A 0.02fF
C14756 NAND2X1_LOC_738/B NAND2X1_LOC_828/a_36_24# 0.00fF
C14757 NOR2X1_LOC_91/A INVX1_LOC_23/A 0.09fF
C14758 NAND2X1_LOC_364/A NOR2X1_LOC_197/B 0.08fF
C14759 NOR2X1_LOC_498/Y NOR2X1_LOC_692/Y 0.02fF
C14760 NAND2X1_LOC_192/B NOR2X1_LOC_89/A 0.02fF
C14761 NOR2X1_LOC_552/A NOR2X1_LOC_548/Y 0.02fF
C14762 NOR2X1_LOC_65/B NAND2X1_LOC_275/a_36_24# 0.02fF
C14763 NOR2X1_LOC_667/A NAND2X1_LOC_650/B 0.05fF
C14764 INPUT_0 NOR2X1_LOC_356/A 0.07fF
C14765 NAND2X1_LOC_560/A NAND2X1_LOC_849/A 0.10fF
C14766 INVX1_LOC_232/Y D_INPUT_3 0.23fF
C14767 NOR2X1_LOC_78/B NAND2X1_LOC_39/Y 0.03fF
C14768 NOR2X1_LOC_151/Y NOR2X1_LOC_439/B 0.03fF
C14769 NOR2X1_LOC_608/a_36_216# INVX1_LOC_2/Y 0.00fF
C14770 NOR2X1_LOC_860/B INVX1_LOC_46/Y 0.01fF
C14771 NAND2X1_LOC_833/Y INVX1_LOC_54/A 0.16fF
C14772 NOR2X1_LOC_92/Y INVX1_LOC_32/A 0.00fF
C14773 NOR2X1_LOC_151/Y INVX1_LOC_75/A 0.07fF
C14774 NOR2X1_LOC_844/A INVX1_LOC_280/A 0.02fF
C14775 NAND2X1_LOC_352/B INVX1_LOC_29/A 0.08fF
C14776 NAND2X1_LOC_363/B NOR2X1_LOC_383/B 0.01fF
C14777 INVX1_LOC_279/A INVX1_LOC_247/A 0.01fF
C14778 NAND2X1_LOC_633/Y INVX1_LOC_25/Y 0.37fF
C14779 INVX1_LOC_24/Y NOR2X1_LOC_623/B 0.02fF
C14780 GATE_741 NAND2X1_LOC_175/Y 0.09fF
C14781 NAND2X1_LOC_462/B NAND2X1_LOC_658/a_36_24# 0.00fF
C14782 INVX1_LOC_189/A INVX1_LOC_38/A 0.00fF
C14783 INVX1_LOC_209/Y NOR2X1_LOC_88/Y 0.08fF
C14784 NOR2X1_LOC_160/Y VDD 0.00fF
C14785 INPUT_0 NOR2X1_LOC_74/A 2.14fF
C14786 NOR2X1_LOC_632/Y INVX1_LOC_46/A 0.00fF
C14787 NOR2X1_LOC_852/A NOR2X1_LOC_777/B 0.04fF
C14788 INVX1_LOC_101/A VDD 0.00fF
C14789 INVX1_LOC_73/A INVX1_LOC_286/A 0.07fF
C14790 INVX1_LOC_63/Y NOR2X1_LOC_592/B 0.07fF
C14791 INVX1_LOC_31/A NOR2X1_LOC_847/a_36_216# 0.01fF
C14792 NAND2X1_LOC_45/a_36_24# NOR2X1_LOC_243/B 0.01fF
C14793 INVX1_LOC_27/A NOR2X1_LOC_302/A 0.03fF
C14794 NOR2X1_LOC_92/Y NAND2X1_LOC_175/Y 0.05fF
C14795 NAND2X1_LOC_837/Y NAND2X1_LOC_489/Y 0.02fF
C14796 INPUT_1 NOR2X1_LOC_124/A 0.02fF
C14797 INVX1_LOC_177/A INVX1_LOC_307/Y 0.02fF
C14798 INPUT_0 NOR2X1_LOC_9/Y 0.14fF
C14799 INVX1_LOC_54/Y NOR2X1_LOC_612/Y 0.34fF
C14800 INVX1_LOC_88/A NAND2X1_LOC_454/Y 0.01fF
C14801 INVX1_LOC_8/A NOR2X1_LOC_179/a_36_216# 0.01fF
C14802 INVX1_LOC_209/Y INVX1_LOC_84/A 0.03fF
C14803 NOR2X1_LOC_598/B INVX1_LOC_213/A 3.39fF
C14804 NOR2X1_LOC_356/A NOR2X1_LOC_324/A 0.13fF
C14805 INVX1_LOC_83/A NOR2X1_LOC_145/Y 0.02fF
C14806 NAND2X1_LOC_552/A NAND2X1_LOC_793/B 0.01fF
C14807 INVX1_LOC_72/A INVX1_LOC_42/A 0.06fF
C14808 INVX1_LOC_276/A INVX1_LOC_92/A 0.03fF
C14809 NOR2X1_LOC_576/B NAND2X1_LOC_839/a_36_24# 0.01fF
C14810 INVX1_LOC_1/Y INVX1_LOC_9/A 1.74fF
C14811 NOR2X1_LOC_554/B NOR2X1_LOC_643/a_36_216# 0.00fF
C14812 NAND2X1_LOC_656/A NOR2X1_LOC_89/A 0.09fF
C14813 NOR2X1_LOC_718/B INVX1_LOC_84/A 0.01fF
C14814 NAND2X1_LOC_20/B NAND2X1_LOC_223/B 0.23fF
C14815 NOR2X1_LOC_160/B NAND2X1_LOC_223/A 0.00fF
C14816 INVX1_LOC_89/A INVX1_LOC_122/A 0.16fF
C14817 NOR2X1_LOC_730/A NOR2X1_LOC_729/A 0.00fF
C14818 INVX1_LOC_11/A NAND2X1_LOC_99/A 0.07fF
C14819 INVX1_LOC_178/A NAND2X1_LOC_793/B 0.10fF
C14820 D_INPUT_1 NAND2X1_LOC_218/A 0.34fF
C14821 INVX1_LOC_147/A NAND2X1_LOC_468/B 0.18fF
C14822 D_INPUT_1 NOR2X1_LOC_140/A 0.03fF
C14823 NOR2X1_LOC_131/Y NOR2X1_LOC_364/A 0.02fF
C14824 INVX1_LOC_269/A NOR2X1_LOC_748/A 0.10fF
C14825 NOR2X1_LOC_781/A INVX1_LOC_54/A 0.78fF
C14826 NOR2X1_LOC_736/Y VDD 0.42fF
C14827 NOR2X1_LOC_68/A NOR2X1_LOC_685/Y 0.06fF
C14828 NOR2X1_LOC_135/Y INVX1_LOC_46/A 0.41fF
C14829 NAND2X1_LOC_554/a_36_24# INVX1_LOC_9/A 0.00fF
C14830 NOR2X1_LOC_845/a_36_216# NOR2X1_LOC_849/A 0.03fF
C14831 NOR2X1_LOC_344/A INVX1_LOC_29/A 0.02fF
C14832 NOR2X1_LOC_457/A NOR2X1_LOC_383/B 0.03fF
C14833 NOR2X1_LOC_644/A INVX1_LOC_117/A 0.03fF
C14834 INVX1_LOC_17/A INVX1_LOC_271/A 0.02fF
C14835 NOR2X1_LOC_208/A INVX1_LOC_76/A 0.23fF
C14836 NOR2X1_LOC_589/A NOR2X1_LOC_364/A 0.55fF
C14837 INVX1_LOC_28/A INVX1_LOC_33/Y 0.05fF
C14838 NOR2X1_LOC_6/B NAND2X1_LOC_63/Y 0.01fF
C14839 INVX1_LOC_161/Y INVX1_LOC_57/A 0.03fF
C14840 INVX1_LOC_280/Y NOR2X1_LOC_485/Y 0.07fF
C14841 NOR2X1_LOC_91/A INVX1_LOC_31/A 0.03fF
C14842 NAND2X1_LOC_840/Y INVX1_LOC_37/A 0.00fF
C14843 NOR2X1_LOC_828/B INVX1_LOC_117/A 0.03fF
C14844 NOR2X1_LOC_561/Y NOR2X1_LOC_435/A 0.05fF
C14845 INVX1_LOC_72/A INVX1_LOC_78/A 0.12fF
C14846 INVX1_LOC_31/A NOR2X1_LOC_668/Y 0.03fF
C14847 NOR2X1_LOC_201/A INVX1_LOC_31/A 0.05fF
C14848 INVX1_LOC_174/A NAND2X1_LOC_40/a_36_24# 0.00fF
C14849 NAND2X1_LOC_357/B INVX1_LOC_29/A 0.10fF
C14850 NOR2X1_LOC_270/Y INVX1_LOC_271/Y 0.07fF
C14851 INVX1_LOC_279/A NOR2X1_LOC_862/B 0.03fF
C14852 NOR2X1_LOC_76/A INVX1_LOC_54/A 0.00fF
C14853 NOR2X1_LOC_739/Y NOR2X1_LOC_678/A 0.03fF
C14854 INVX1_LOC_13/A NAND2X1_LOC_574/A -0.07fF
C14855 NAND2X1_LOC_315/a_36_24# INVX1_LOC_94/Y 0.00fF
C14856 INVX1_LOC_36/A NOR2X1_LOC_447/A 0.03fF
C14857 NAND2X1_LOC_47/a_36_24# INVX1_LOC_53/A 0.00fF
C14858 INVX1_LOC_8/A NAND2X1_LOC_74/a_36_24# 0.00fF
C14859 NOR2X1_LOC_589/A INVX1_LOC_285/A 0.07fF
C14860 NOR2X1_LOC_423/Y NOR2X1_LOC_89/A 0.26fF
C14861 INVX1_LOC_35/A INVX1_LOC_256/A 0.04fF
C14862 INVX1_LOC_288/A INVX1_LOC_72/A 0.06fF
C14863 INVX1_LOC_31/A INVX1_LOC_23/A 0.08fF
C14864 INVX1_LOC_30/A NOR2X1_LOC_383/B 2.59fF
C14865 INVX1_LOC_41/A INVX1_LOC_32/A 0.05fF
C14866 NOR2X1_LOC_65/B INVX1_LOC_72/A 0.12fF
C14867 NAND2X1_LOC_549/B INVX1_LOC_29/A 0.01fF
C14868 INVX1_LOC_35/A NOR2X1_LOC_647/B 0.53fF
C14869 NOR2X1_LOC_32/B INVX1_LOC_230/Y 0.17fF
C14870 INVX1_LOC_75/A NOR2X1_LOC_707/A 0.14fF
C14871 INVX1_LOC_201/Y INVX1_LOC_32/A 0.72fF
C14872 NOR2X1_LOC_742/A INVX1_LOC_9/A 0.07fF
C14873 INVX1_LOC_70/Y INVX1_LOC_20/A 0.10fF
C14874 INVX1_LOC_285/Y NOR2X1_LOC_363/Y 0.10fF
C14875 INVX1_LOC_77/A INVX1_LOC_87/A 0.03fF
C14876 NOR2X1_LOC_557/a_36_216# NAND2X1_LOC_447/Y 0.03fF
C14877 INVX1_LOC_75/A NOR2X1_LOC_709/B 0.01fF
C14878 NOR2X1_LOC_168/B NOR2X1_LOC_640/B 0.01fF
C14879 NOR2X1_LOC_537/Y INVX1_LOC_42/A 0.06fF
C14880 NOR2X1_LOC_222/Y NOR2X1_LOC_89/A 0.03fF
C14881 INVX1_LOC_73/A INVX1_LOC_54/A 0.07fF
C14882 NOR2X1_LOC_561/Y INVX1_LOC_63/A 0.02fF
C14883 INVX1_LOC_75/A NOR2X1_LOC_209/B 0.03fF
C14884 INVX1_LOC_217/A NAND2X1_LOC_787/Y 0.02fF
C14885 NAND2X1_LOC_338/B INVX1_LOC_42/A 0.09fF
C14886 NAND2X1_LOC_477/A INVX1_LOC_32/A 0.03fF
C14887 INVX1_LOC_7/A INVX1_LOC_63/A 0.39fF
C14888 NOR2X1_LOC_514/A NOR2X1_LOC_660/Y 0.03fF
C14889 NOR2X1_LOC_78/A INVX1_LOC_37/A 0.22fF
C14890 INVX1_LOC_222/Y INVX1_LOC_11/A 0.03fF
C14891 INVX1_LOC_17/A INVX1_LOC_27/A 0.20fF
C14892 INVX1_LOC_171/A INVX1_LOC_285/A 0.01fF
C14893 INVX1_LOC_57/Y NAND2X1_LOC_787/A 0.03fF
C14894 INVX1_LOC_17/A NOR2X1_LOC_824/A 0.34fF
C14895 NAND2X1_LOC_784/A INVX1_LOC_18/A 0.07fF
C14896 NAND2X1_LOC_861/Y INVX1_LOC_119/Y 0.07fF
C14897 NOR2X1_LOC_540/a_36_216# INVX1_LOC_29/A 0.00fF
C14898 NAND2X1_LOC_660/Y INVX1_LOC_49/Y 0.03fF
C14899 INVX1_LOC_30/Y NAND2X1_LOC_63/Y 1.44fF
C14900 NOR2X1_LOC_636/B NAND2X1_LOC_149/Y 0.02fF
C14901 NOR2X1_LOC_274/B INVX1_LOC_58/Y 0.15fF
C14902 NAND2X1_LOC_859/B INVX1_LOC_284/A 0.37fF
C14903 INVX1_LOC_171/A NOR2X1_LOC_814/A 0.11fF
C14904 NAND2X1_LOC_361/Y INVX1_LOC_26/A 0.03fF
C14905 NOR2X1_LOC_790/B INVX1_LOC_247/Y 0.01fF
C14906 NOR2X1_LOC_471/Y INVX1_LOC_27/A 0.02fF
C14907 NOR2X1_LOC_180/Y INVX1_LOC_271/Y 0.04fF
C14908 INVX1_LOC_136/A NAND2X1_LOC_624/B 0.03fF
C14909 NOR2X1_LOC_598/B NOR2X1_LOC_196/A 0.05fF
C14910 INVX1_LOC_45/A INVX1_LOC_5/A 0.07fF
C14911 NAND2X1_LOC_725/Y NAND2X1_LOC_733/a_36_24# 0.09fF
C14912 NOR2X1_LOC_355/A INVX1_LOC_133/A 0.12fF
C14913 NAND2X1_LOC_555/Y INVX1_LOC_27/A 0.16fF
C14914 D_INPUT_0 INVX1_LOC_49/Y 0.03fF
C14915 INVX1_LOC_126/A VDD 0.28fF
C14916 INVX1_LOC_136/A NOR2X1_LOC_211/Y 0.05fF
C14917 NOR2X1_LOC_577/Y NOR2X1_LOC_654/A 0.10fF
C14918 INVX1_LOC_5/A NOR2X1_LOC_568/A 0.03fF
C14919 INVX1_LOC_218/A INVX1_LOC_15/A 0.03fF
C14920 NOR2X1_LOC_128/B INVX1_LOC_29/A 0.14fF
C14921 INVX1_LOC_124/A INVX1_LOC_87/A 0.00fF
C14922 NAND2X1_LOC_477/A NAND2X1_LOC_175/Y 0.10fF
C14923 INVX1_LOC_36/A NOR2X1_LOC_34/B 0.01fF
C14924 NAND2X1_LOC_357/B NOR2X1_LOC_281/Y 0.02fF
C14925 NOR2X1_LOC_211/A INVX1_LOC_32/A 0.03fF
C14926 NAND2X1_LOC_39/Y INVX1_LOC_46/A 0.01fF
C14927 INVX1_LOC_180/A INVX1_LOC_53/A 0.05fF
C14928 NOR2X1_LOC_537/Y INVX1_LOC_78/A 9.50fF
C14929 INVX1_LOC_255/Y INVX1_LOC_3/Y 0.16fF
C14930 NAND2X1_LOC_338/B INVX1_LOC_78/A 0.23fF
C14931 NOR2X1_LOC_15/Y NOR2X1_LOC_134/Y 0.11fF
C14932 NOR2X1_LOC_78/A INVX1_LOC_157/Y 0.00fF
C14933 INVX1_LOC_10/A NOR2X1_LOC_114/Y 0.02fF
C14934 NAND2X1_LOC_464/Y NAND2X1_LOC_464/B 0.02fF
C14935 NOR2X1_LOC_52/B NAND2X1_LOC_99/A 0.00fF
C14936 NOR2X1_LOC_226/A INVX1_LOC_273/A 0.03fF
C14937 INPUT_0 NOR2X1_LOC_243/B 0.05fF
C14938 INVX1_LOC_72/Y INVX1_LOC_306/Y 0.35fF
C14939 NOR2X1_LOC_458/B INVX1_LOC_271/Y 0.00fF
C14940 NOR2X1_LOC_111/A VDD 0.92fF
C14941 NOR2X1_LOC_763/A INVX1_LOC_30/A 0.06fF
C14942 NOR2X1_LOC_582/A INVX1_LOC_30/A 0.04fF
C14943 INVX1_LOC_313/Y INVX1_LOC_263/Y 0.01fF
C14944 NOR2X1_LOC_646/A INVX1_LOC_4/Y 0.07fF
C14945 INVX1_LOC_64/A NAND2X1_LOC_567/Y 0.00fF
C14946 INVX1_LOC_21/A INVX1_LOC_177/Y 0.08fF
C14947 INVX1_LOC_114/A INVX1_LOC_115/A 0.11fF
C14948 NAND2X1_LOC_552/A INVX1_LOC_71/A 0.18fF
C14949 NAND2X1_LOC_325/Y INVX1_LOC_53/A 0.07fF
C14950 INVX1_LOC_5/A INVX1_LOC_71/A 0.14fF
C14951 INVX1_LOC_121/A INVX1_LOC_32/A 0.02fF
C14952 NAND2X1_LOC_773/a_36_24# NAND2X1_LOC_338/B 0.00fF
C14953 VDD NOR2X1_LOC_694/Y 0.24fF
C14954 NOR2X1_LOC_516/B NAND2X1_LOC_223/A 0.03fF
C14955 NOR2X1_LOC_285/Y NAND2X1_LOC_364/Y 0.02fF
C14956 NOR2X1_LOC_307/A NAND2X1_LOC_305/a_36_24# 0.02fF
C14957 NOR2X1_LOC_382/Y INVX1_LOC_14/A 0.06fF
C14958 NOR2X1_LOC_65/B NAND2X1_LOC_338/B 0.10fF
C14959 INVX1_LOC_38/A NAND2X1_LOC_211/Y 0.08fF
C14960 INVX1_LOC_313/Y INVX1_LOC_42/A 0.07fF
C14961 NOR2X1_LOC_272/Y NOR2X1_LOC_191/B 0.31fF
C14962 NAND2X1_LOC_326/A INVX1_LOC_18/A 0.07fF
C14963 NOR2X1_LOC_24/Y NOR2X1_LOC_629/Y 0.02fF
C14964 INVX1_LOC_1/A NAND2X1_LOC_16/Y 0.12fF
C14965 INVX1_LOC_41/Y NAND2X1_LOC_793/a_36_24# 0.00fF
C14966 NOR2X1_LOC_71/Y INVX1_LOC_3/Y 0.00fF
C14967 NOR2X1_LOC_329/B NOR2X1_LOC_89/A 0.07fF
C14968 NAND2X1_LOC_538/a_36_24# INVX1_LOC_49/Y 0.00fF
C14969 NOR2X1_LOC_167/Y INVX1_LOC_63/A 0.94fF
C14970 D_INPUT_1 NOR2X1_LOC_709/A 0.03fF
C14971 INVX1_LOC_177/A INVX1_LOC_29/Y 0.04fF
C14972 NAND2X1_LOC_251/a_36_24# INVX1_LOC_63/A 0.00fF
C14973 INVX1_LOC_16/A INVX1_LOC_23/Y 0.25fF
C14974 INVX1_LOC_191/Y INVX1_LOC_23/A 0.03fF
C14975 NAND2X1_LOC_348/A NAND2X1_LOC_207/B 0.02fF
C14976 NAND2X1_LOC_156/B NOR2X1_LOC_158/B 0.04fF
C14977 INVX1_LOC_279/A NOR2X1_LOC_465/Y 0.10fF
C14978 VDD INVX1_LOC_127/A 0.00fF
C14979 NOR2X1_LOC_68/A INVX1_LOC_88/A 0.03fF
C14980 INVX1_LOC_133/Y INVX1_LOC_53/A 0.02fF
C14981 INVX1_LOC_45/A NAND2X1_LOC_337/B 0.27fF
C14982 NAND2X1_LOC_706/Y INVX1_LOC_24/A 0.05fF
C14983 INVX1_LOC_45/A NOR2X1_LOC_816/A 0.03fF
C14984 INVX1_LOC_276/A INVX1_LOC_53/A 0.03fF
C14985 NOR2X1_LOC_333/a_36_216# INVX1_LOC_15/A 0.01fF
C14986 INVX1_LOC_222/Y NOR2X1_LOC_593/Y 0.04fF
C14987 NOR2X1_LOC_435/A INVX1_LOC_76/A 0.34fF
C14988 NOR2X1_LOC_352/Y NOR2X1_LOC_678/A 0.03fF
C14989 INVX1_LOC_22/A NOR2X1_LOC_654/A 0.32fF
C14990 NOR2X1_LOC_807/B NOR2X1_LOC_325/Y 0.05fF
C14991 INVX1_LOC_290/A NOR2X1_LOC_651/a_36_216# 0.00fF
C14992 INVX1_LOC_84/Y NOR2X1_LOC_476/B 0.01fF
C14993 NAND2X1_LOC_387/B NOR2X1_LOC_389/A 0.11fF
C14994 INVX1_LOC_54/Y NAND2X1_LOC_406/a_36_24# 0.00fF
C14995 NOR2X1_LOC_368/a_36_216# NAND2X1_LOC_74/B 0.00fF
C14996 NOR2X1_LOC_15/Y INVX1_LOC_49/A 0.07fF
C14997 NAND2X1_LOC_648/A INVX1_LOC_273/A 0.26fF
C14998 INVX1_LOC_141/Y INVX1_LOC_312/Y 0.12fF
C14999 NOR2X1_LOC_538/B INVX1_LOC_314/Y 0.05fF
C15000 INVX1_LOC_152/Y NAND2X1_LOC_323/B 0.00fF
C15001 INVX1_LOC_313/Y INVX1_LOC_78/A 0.07fF
C15002 INVX1_LOC_21/A INVX1_LOC_104/A 0.14fF
C15003 NOR2X1_LOC_709/A NOR2X1_LOC_652/Y 0.02fF
C15004 NOR2X1_LOC_510/Y NOR2X1_LOC_361/Y 0.04fF
C15005 NOR2X1_LOC_793/A INVX1_LOC_33/A 0.01fF
C15006 INVX1_LOC_20/A INVX1_LOC_285/A 0.07fF
C15007 INVX1_LOC_57/Y INVX1_LOC_30/A 0.04fF
C15008 INVX1_LOC_22/A INVX1_LOC_58/Y 0.07fF
C15009 NAND2X1_LOC_337/B INVX1_LOC_71/A 0.21fF
C15010 NOR2X1_LOC_76/A NOR2X1_LOC_438/Y 0.04fF
C15011 NOR2X1_LOC_82/A INVX1_LOC_77/A 0.07fF
C15012 NOR2X1_LOC_719/B NAND2X1_LOC_215/A 0.21fF
C15013 INVX1_LOC_13/Y NAND2X1_LOC_464/a_36_24# 0.01fF
C15014 NAND2X1_LOC_123/Y INVX1_LOC_94/Y 0.01fF
C15015 INVX1_LOC_89/A NOR2X1_LOC_621/A 0.01fF
C15016 INVX1_LOC_76/A INVX1_LOC_63/A 0.24fF
C15017 NOR2X1_LOC_357/Y INVX1_LOC_136/Y 0.01fF
C15018 INVX1_LOC_182/Y NOR2X1_LOC_465/Y 0.00fF
C15019 NOR2X1_LOC_91/A NAND2X1_LOC_866/B 0.11fF
C15020 NAND2X1_LOC_778/Y NOR2X1_LOC_226/A 0.10fF
C15021 INVX1_LOC_41/A NOR2X1_LOC_296/Y 0.01fF
C15022 NAND2X1_LOC_574/A NOR2X1_LOC_34/a_36_216# 0.01fF
C15023 INVX1_LOC_28/A INVX1_LOC_23/Y 0.10fF
C15024 NOR2X1_LOC_391/A NOR2X1_LOC_392/Y 0.00fF
C15025 INVX1_LOC_58/A NOR2X1_LOC_71/Y 0.18fF
C15026 NOR2X1_LOC_91/A NAND2X1_LOC_807/Y 0.79fF
C15027 NOR2X1_LOC_160/B INVX1_LOC_33/A 9.43fF
C15028 INVX1_LOC_313/A INVX1_LOC_23/A 1.01fF
C15029 NOR2X1_LOC_591/Y NAND2X1_LOC_538/Y 0.10fF
C15030 NAND2X1_LOC_563/Y INVX1_LOC_228/Y 0.00fF
C15031 INVX1_LOC_2/A NOR2X1_LOC_15/Y 3.79fF
C15032 NAND2X1_LOC_472/Y INVX1_LOC_84/A 0.07fF
C15033 NOR2X1_LOC_361/B NOR2X1_LOC_361/Y 0.07fF
C15034 NOR2X1_LOC_831/B INVX1_LOC_118/Y 0.03fF
C15035 INVX1_LOC_100/A NOR2X1_LOC_394/Y 0.01fF
C15036 INVX1_LOC_35/A NOR2X1_LOC_415/A 0.01fF
C15037 NOR2X1_LOC_635/A NAND2X1_LOC_30/Y 0.02fF
C15038 INVX1_LOC_136/A INVX1_LOC_41/Y 0.03fF
C15039 NAND2X1_LOC_36/A INVX1_LOC_77/A 0.56fF
C15040 INVX1_LOC_201/Y INPUT_3 0.08fF
C15041 NOR2X1_LOC_226/A NOR2X1_LOC_15/Y 0.88fF
C15042 INVX1_LOC_58/A NOR2X1_LOC_644/A 0.27fF
C15043 INVX1_LOC_17/A INVX1_LOC_206/A 0.09fF
C15044 NOR2X1_LOC_806/Y INVX1_LOC_269/Y 0.00fF
C15045 NOR2X1_LOC_545/A NOR2X1_LOC_500/B 0.03fF
C15046 INVX1_LOC_30/A NAND2X1_LOC_632/B 0.01fF
C15047 NOR2X1_LOC_690/A INVX1_LOC_284/Y 0.17fF
C15048 INVX1_LOC_72/A NOR2X1_LOC_152/Y 0.07fF
C15049 NAND2X1_LOC_463/B NAND2X1_LOC_402/B 0.00fF
C15050 NOR2X1_LOC_74/A INVX1_LOC_183/A 0.03fF
C15051 NOR2X1_LOC_537/A NOR2X1_LOC_274/B 0.01fF
C15052 INVX1_LOC_216/Y INVX1_LOC_216/A 0.18fF
C15053 NOR2X1_LOC_250/Y NAND2X1_LOC_231/Y 0.03fF
C15054 INVX1_LOC_72/A INVX1_LOC_113/Y 0.02fF
C15055 VDD NOR2X1_LOC_583/Y 0.12fF
C15056 INVX1_LOC_223/A INVX1_LOC_67/A 0.00fF
C15057 INVX1_LOC_303/A NOR2X1_LOC_68/A 0.08fF
C15058 INVX1_LOC_17/A NAND2X1_LOC_200/B 0.03fF
C15059 NAND2X1_LOC_79/a_36_24# NOR2X1_LOC_68/A 0.01fF
C15060 NAND2X1_LOC_564/B NOR2X1_LOC_92/Y 0.00fF
C15061 INVX1_LOC_315/Y NAND2X1_LOC_223/A 0.03fF
C15062 NOR2X1_LOC_160/B NOR2X1_LOC_714/Y 0.03fF
C15063 INVX1_LOC_11/A NOR2X1_LOC_222/Y 0.06fF
C15064 INVX1_LOC_17/A NOR2X1_LOC_251/Y 0.04fF
C15065 NAND2X1_LOC_848/A INVX1_LOC_49/Y 0.01fF
C15066 NOR2X1_LOC_91/A INVX1_LOC_6/A 0.03fF
C15067 NOR2X1_LOC_609/A NOR2X1_LOC_577/Y 0.03fF
C15068 INVX1_LOC_140/A NAND2X1_LOC_793/B 0.18fF
C15069 INVX1_LOC_96/A NOR2X1_LOC_631/Y 0.25fF
C15070 NAND2X1_LOC_721/B NAND2X1_LOC_357/B 0.08fF
C15071 NOR2X1_LOC_846/Y NOR2X1_LOC_846/B 0.00fF
C15072 NOR2X1_LOC_546/B INVX1_LOC_275/A 0.03fF
C15073 NAND2X1_LOC_656/A NOR2X1_LOC_593/Y 0.01fF
C15074 NOR2X1_LOC_15/Y NAND2X1_LOC_462/B 0.02fF
C15075 NOR2X1_LOC_160/B INVX1_LOC_40/A 0.12fF
C15076 NAND2X1_LOC_659/B INVX1_LOC_253/A 0.05fF
C15077 NOR2X1_LOC_75/Y INVX1_LOC_22/A 2.02fF
C15078 INVX1_LOC_274/A INVX1_LOC_19/A 0.08fF
C15079 NOR2X1_LOC_300/Y INVX1_LOC_18/A 0.02fF
C15080 INVX1_LOC_6/A INVX1_LOC_23/A 0.64fF
C15081 NOR2X1_LOC_226/A NAND2X1_LOC_355/a_36_24# 0.00fF
C15082 INVX1_LOC_123/A NAND2X1_LOC_607/a_36_24# 0.00fF
C15083 NOR2X1_LOC_596/Y INVX1_LOC_16/A 0.02fF
C15084 INVX1_LOC_269/A INVX1_LOC_150/A 0.01fF
C15085 INVX1_LOC_2/Y INVX1_LOC_4/Y 0.03fF
C15086 INVX1_LOC_45/A NOR2X1_LOC_773/Y 0.07fF
C15087 INVX1_LOC_229/A NOR2X1_LOC_576/B 0.03fF
C15088 INVX1_LOC_50/A NOR2X1_LOC_269/Y 0.07fF
C15089 NAND2X1_LOC_472/Y INVX1_LOC_15/A 0.04fF
C15090 NOR2X1_LOC_554/B NOR2X1_LOC_537/Y 0.07fF
C15091 NOR2X1_LOC_15/Y NAND2X1_LOC_648/A 0.03fF
C15092 VDD INVX1_LOC_253/A -0.00fF
C15093 INVX1_LOC_269/A INVX1_LOC_89/A 0.24fF
C15094 NOR2X1_LOC_626/a_36_216# NOR2X1_LOC_742/A 0.01fF
C15095 NOR2X1_LOC_274/Y NOR2X1_LOC_309/Y 0.08fF
C15096 VDD INVX1_LOC_90/Y 0.21fF
C15097 NOR2X1_LOC_606/Y NOR2X1_LOC_121/A 0.01fF
C15098 NOR2X1_LOC_15/Y INPUT_1 0.14fF
C15099 NOR2X1_LOC_590/A NOR2X1_LOC_589/A 0.03fF
C15100 INVX1_LOC_257/A NOR2X1_LOC_684/Y 0.01fF
C15101 NOR2X1_LOC_232/Y INVX1_LOC_89/A 0.11fF
C15102 NAND2X1_LOC_304/a_36_24# INVX1_LOC_142/A 0.00fF
C15103 NOR2X1_LOC_307/B INVX1_LOC_142/Y 0.01fF
C15104 INVX1_LOC_314/Y NOR2X1_LOC_315/Y 0.07fF
C15105 INVX1_LOC_116/A INVX1_LOC_149/A 0.01fF
C15106 NOR2X1_LOC_220/B NOR2X1_LOC_74/A 0.01fF
C15107 NAND2X1_LOC_859/Y INVX1_LOC_31/A 3.12fF
C15108 INVX1_LOC_33/A NOR2X1_LOC_317/B 0.03fF
C15109 NAND2X1_LOC_170/A INVX1_LOC_30/A 0.01fF
C15110 NAND2X1_LOC_363/B NAND2X1_LOC_826/a_36_24# 0.01fF
C15111 INVX1_LOC_75/A NOR2X1_LOC_343/B 0.02fF
C15112 NAND2X1_LOC_741/B INVX1_LOC_16/A 0.02fF
C15113 NOR2X1_LOC_763/Y INVX1_LOC_174/A 0.57fF
C15114 NOR2X1_LOC_740/Y INVX1_LOC_85/Y 0.13fF
C15115 NOR2X1_LOC_390/a_36_216# INVX1_LOC_155/Y 0.00fF
C15116 NAND2X1_LOC_364/A NOR2X1_LOC_568/a_36_216# 0.01fF
C15117 INVX1_LOC_1/A INVX1_LOC_148/A 0.01fF
C15118 INVX1_LOC_34/A NOR2X1_LOC_121/Y 0.04fF
C15119 NOR2X1_LOC_584/Y INVX1_LOC_92/A 0.03fF
C15120 INVX1_LOC_24/A NAND2X1_LOC_483/a_36_24# 0.00fF
C15121 INVX1_LOC_52/Y NOR2X1_LOC_202/Y 0.33fF
C15122 INVX1_LOC_76/A NOR2X1_LOC_65/Y 0.01fF
C15123 NOR2X1_LOC_606/a_36_216# INVX1_LOC_7/A 0.00fF
C15124 INVX1_LOC_35/A NOR2X1_LOC_725/A 0.02fF
C15125 INVX1_LOC_84/A NAND2X1_LOC_773/B 0.07fF
C15126 INVX1_LOC_49/A INVX1_LOC_96/Y 0.21fF
C15127 NAND2X1_LOC_783/A NAND2X1_LOC_516/a_36_24# 0.00fF
C15128 NOR2X1_LOC_812/A NOR2X1_LOC_856/A 0.01fF
C15129 NAND2X1_LOC_579/A NOR2X1_LOC_322/Y 0.10fF
C15130 NOR2X1_LOC_773/Y INVX1_LOC_71/A 0.10fF
C15131 NOR2X1_LOC_724/a_36_216# NOR2X1_LOC_374/A 0.00fF
C15132 NOR2X1_LOC_590/A INVX1_LOC_171/A 0.00fF
C15133 NOR2X1_LOC_419/Y NOR2X1_LOC_346/B 0.03fF
C15134 INVX1_LOC_11/A NOR2X1_LOC_329/B 0.07fF
C15135 INVX1_LOC_225/Y NOR2X1_LOC_356/A 0.36fF
C15136 INVX1_LOC_81/Y NAND2X1_LOC_140/A 0.00fF
C15137 NAND2X1_LOC_656/Y INVX1_LOC_312/Y 0.21fF
C15138 NAND2X1_LOC_112/Y NAND2X1_LOC_198/B 0.03fF
C15139 NOR2X1_LOC_222/Y NOR2X1_LOC_433/A 0.03fF
C15140 INVX1_LOC_45/A NOR2X1_LOC_332/A 0.01fF
C15141 INVX1_LOC_279/A NOR2X1_LOC_52/Y 0.00fF
C15142 INVX1_LOC_88/A INVX1_LOC_147/A 0.01fF
C15143 NAND2X1_LOC_267/B INVX1_LOC_29/Y 0.05fF
C15144 INVX1_LOC_49/A INVX1_LOC_226/A 0.01fF
C15145 INVX1_LOC_11/A D_INPUT_4 0.03fF
C15146 INVX1_LOC_21/A INVX1_LOC_86/Y 0.22fF
C15147 INVX1_LOC_87/A INVX1_LOC_9/A 0.03fF
C15148 NOR2X1_LOC_39/Y INVX1_LOC_117/A 0.09fF
C15149 NOR2X1_LOC_52/B NOR2X1_LOC_423/Y 0.00fF
C15150 NOR2X1_LOC_819/a_36_216# NOR2X1_LOC_332/A 0.01fF
C15151 NOR2X1_LOC_269/a_36_216# NOR2X1_LOC_433/A 0.01fF
C15152 INVX1_LOC_31/A NAND2X1_LOC_807/Y 0.07fF
C15153 INVX1_LOC_174/Y NOR2X1_LOC_713/B 0.25fF
C15154 NOR2X1_LOC_537/A INVX1_LOC_22/A 0.01fF
C15155 NAND2X1_LOC_555/Y NOR2X1_LOC_19/B 0.24fF
C15156 INVX1_LOC_208/A INVX1_LOC_33/A 0.03fF
C15157 INVX1_LOC_256/A NOR2X1_LOC_534/a_36_216# 0.01fF
C15158 NOR2X1_LOC_716/B INVX1_LOC_22/A 0.05fF
C15159 NOR2X1_LOC_516/B INVX1_LOC_33/A 0.05fF
C15160 NAND2X1_LOC_574/A INVX1_LOC_32/A 0.01fF
C15161 INVX1_LOC_2/A INVX1_LOC_96/Y 0.94fF
C15162 NOR2X1_LOC_471/Y NOR2X1_LOC_589/a_36_216# 0.01fF
C15163 INVX1_LOC_225/Y NOR2X1_LOC_74/A 0.15fF
C15164 INVX1_LOC_39/A NOR2X1_LOC_124/A 1.52fF
C15165 NOR2X1_LOC_222/Y NOR2X1_LOC_52/B 0.05fF
C15166 NAND2X1_LOC_341/A NOR2X1_LOC_364/Y 0.02fF
C15167 VDD INVX1_LOC_138/Y 0.02fF
C15168 NAND2X1_LOC_479/Y INVX1_LOC_63/Y 0.07fF
C15169 NAND2X1_LOC_727/Y INVX1_LOC_34/A 0.01fF
C15170 NOR2X1_LOC_78/B INVX1_LOC_133/Y 0.98fF
C15171 NAND2X1_LOC_338/B NOR2X1_LOC_721/A 0.04fF
C15172 INVX1_LOC_136/Y INVX1_LOC_32/A 0.02fF
C15173 NAND2X1_LOC_206/Y INVX1_LOC_15/A 0.08fF
C15174 INVX1_LOC_180/A INVX1_LOC_83/A 0.13fF
C15175 INVX1_LOC_276/A NOR2X1_LOC_78/B 0.05fF
C15176 NAND2X1_LOC_862/Y INVX1_LOC_41/Y 0.01fF
C15177 NOR2X1_LOC_249/Y NOR2X1_LOC_35/Y 0.01fF
C15178 INVX1_LOC_4/A NOR2X1_LOC_814/A 0.26fF
C15179 NOR2X1_LOC_590/A INVX1_LOC_222/A 0.02fF
C15180 INVX1_LOC_226/Y NOR2X1_LOC_398/a_36_216# 0.00fF
C15181 NOR2X1_LOC_67/A NOR2X1_LOC_78/B 0.07fF
C15182 INVX1_LOC_2/A NAND2X1_LOC_840/B 0.01fF
C15183 INVX1_LOC_55/Y INVX1_LOC_94/A -0.03fF
C15184 NAND2X1_LOC_564/B NAND2X1_LOC_477/A 0.10fF
C15185 NOR2X1_LOC_65/B NOR2X1_LOC_79/a_36_216# 0.01fF
C15186 NAND2X1_LOC_722/A NAND2X1_LOC_170/A 0.02fF
C15187 NOR2X1_LOC_454/Y NOR2X1_LOC_300/a_36_216# 0.01fF
C15188 INVX1_LOC_31/A INVX1_LOC_6/A 0.03fF
C15189 INVX1_LOC_255/Y NOR2X1_LOC_515/a_36_216# 0.01fF
C15190 NOR2X1_LOC_272/Y VDD 2.99fF
C15191 INVX1_LOC_53/A NOR2X1_LOC_729/A 0.37fF
C15192 INVX1_LOC_8/Y INVX1_LOC_90/A 0.01fF
C15193 NOR2X1_LOC_690/A NOR2X1_LOC_525/Y 0.42fF
C15194 NOR2X1_LOC_637/B INVX1_LOC_90/A 0.02fF
C15195 INVX1_LOC_34/A D_INPUT_0 3.01fF
C15196 INVX1_LOC_58/A NAND2X1_LOC_243/Y 0.01fF
C15197 INVX1_LOC_177/A INVX1_LOC_101/A 0.00fF
C15198 INVX1_LOC_104/A NOR2X1_LOC_565/B 0.01fF
C15199 NOR2X1_LOC_507/A INVX1_LOC_210/A 0.10fF
C15200 NOR2X1_LOC_445/a_36_216# INVX1_LOC_91/A 0.01fF
C15201 NOR2X1_LOC_791/A INPUT_0 0.01fF
C15202 INVX1_LOC_269/A NOR2X1_LOC_24/Y 0.16fF
C15203 INVX1_LOC_131/Y INVX1_LOC_23/A 0.08fF
C15204 NAND2X1_LOC_794/B INVX1_LOC_33/Y 0.20fF
C15205 NAND2X1_LOC_364/A NOR2X1_LOC_721/Y 0.00fF
C15206 INVX1_LOC_96/Y NAND2X1_LOC_664/a_36_24# 0.00fF
C15207 INVX1_LOC_18/A NOR2X1_LOC_527/Y 0.01fF
C15208 INVX1_LOC_140/A INVX1_LOC_71/A 0.03fF
C15209 NAND2X1_LOC_573/Y INVX1_LOC_37/A 0.03fF
C15210 NOR2X1_LOC_717/B NOR2X1_LOC_348/B 0.05fF
C15211 NOR2X1_LOC_590/A NOR2X1_LOC_311/a_36_216# 0.00fF
C15212 NAND2X1_LOC_67/Y INVX1_LOC_139/A 0.00fF
C15213 INVX1_LOC_303/A NAND2X1_LOC_150/a_36_24# -0.02fF
C15214 INVX1_LOC_15/Y NAND2X1_LOC_462/B 0.01fF
C15215 NOR2X1_LOC_516/B INVX1_LOC_40/A 0.20fF
C15216 NAND2X1_LOC_11/a_36_24# INPUT_5 0.01fF
C15217 NOR2X1_LOC_433/A NOR2X1_LOC_329/B 1.67fF
C15218 NOR2X1_LOC_731/Y NOR2X1_LOC_687/Y 0.03fF
C15219 NOR2X1_LOC_264/Y INVX1_LOC_90/A 1.54fF
C15220 INVX1_LOC_50/Y INVX1_LOC_230/A 0.07fF
C15221 NOR2X1_LOC_381/Y D_INPUT_3 0.03fF
C15222 NAND2X1_LOC_199/B NOR2X1_LOC_45/B 0.03fF
C15223 NAND2X1_LOC_652/a_36_24# NAND2X1_LOC_652/Y 0.02fF
C15224 NOR2X1_LOC_355/A INVX1_LOC_177/A 0.00fF
C15225 INVX1_LOC_84/A NOR2X1_LOC_481/a_36_216# 0.00fF
C15226 INVX1_LOC_232/A INVX1_LOC_16/A 0.17fF
C15227 NOR2X1_LOC_843/A NOR2X1_LOC_174/A 0.02fF
C15228 INVX1_LOC_235/Y INVX1_LOC_166/Y 0.03fF
C15229 NAND2X1_LOC_218/a_36_24# NOR2X1_LOC_673/A 0.00fF
C15230 NAND2X1_LOC_477/a_36_24# INVX1_LOC_19/A 0.00fF
C15231 NAND2X1_LOC_714/B NOR2X1_LOC_536/A 0.04fF
C15232 NOR2X1_LOC_458/B INVX1_LOC_279/A 0.01fF
C15233 NAND2X1_LOC_803/B INVX1_LOC_20/A 0.00fF
C15234 NAND2X1_LOC_708/a_36_24# NOR2X1_LOC_45/B 0.00fF
C15235 NOR2X1_LOC_644/A NOR2X1_LOC_344/a_36_216# 0.00fF
C15236 NOR2X1_LOC_798/A NOR2X1_LOC_186/a_36_216# 0.00fF
C15237 D_INPUT_0 NAND2X1_LOC_231/Y 0.10fF
C15238 INVX1_LOC_64/A NOR2X1_LOC_364/A 0.08fF
C15239 INVX1_LOC_23/A NOR2X1_LOC_117/Y 0.01fF
C15240 NOR2X1_LOC_615/Y INVX1_LOC_20/A 0.01fF
C15241 NOR2X1_LOC_82/A NOR2X1_LOC_138/a_36_216# 0.00fF
C15242 NAND2X1_LOC_778/Y INVX1_LOC_118/A 0.01fF
C15243 INVX1_LOC_33/A NOR2X1_LOC_706/A 0.49fF
C15244 NAND2X1_LOC_141/A INPUT_1 0.08fF
C15245 NOR2X1_LOC_383/Y INVX1_LOC_16/A 0.07fF
C15246 NOR2X1_LOC_202/Y INVX1_LOC_63/Y 0.04fF
C15247 NOR2X1_LOC_435/a_36_216# NOR2X1_LOC_592/B 0.00fF
C15248 INVX1_LOC_49/A NAND2X1_LOC_2/a_36_24# 0.00fF
C15249 NAND2X1_LOC_35/Y INVX1_LOC_260/A 0.02fF
C15250 INVX1_LOC_73/A NOR2X1_LOC_142/Y 0.75fF
C15251 NOR2X1_LOC_590/A INVX1_LOC_20/A 0.06fF
C15252 NOR2X1_LOC_561/Y INVX1_LOC_1/Y 0.10fF
C15253 NOR2X1_LOC_726/Y NOR2X1_LOC_209/A 0.18fF
C15254 INVX1_LOC_107/A NOR2X1_LOC_45/B 0.01fF
C15255 NOR2X1_LOC_329/B NOR2X1_LOC_52/B 0.18fF
C15256 NOR2X1_LOC_773/Y NOR2X1_LOC_123/B 0.01fF
C15257 NOR2X1_LOC_186/Y NOR2X1_LOC_743/Y 0.20fF
C15258 NAND2X1_LOC_561/B NOR2X1_LOC_536/A 0.08fF
C15259 NOR2X1_LOC_424/Y INVX1_LOC_22/A 0.03fF
C15260 NOR2X1_LOC_326/Y NOR2X1_LOC_325/A 0.03fF
C15261 INVX1_LOC_5/A NOR2X1_LOC_592/B 0.01fF
C15262 NOR2X1_LOC_716/B INVX1_LOC_100/A 0.07fF
C15263 NAND2X1_LOC_563/A INVX1_LOC_89/A 0.08fF
C15264 NOR2X1_LOC_717/B INVX1_LOC_22/A 0.00fF
C15265 NOR2X1_LOC_238/Y INVX1_LOC_91/A 0.03fF
C15266 NOR2X1_LOC_62/a_36_216# NOR2X1_LOC_99/B 0.01fF
C15267 NOR2X1_LOC_15/Y INVX1_LOC_118/A 0.16fF
C15268 NOR2X1_LOC_147/B INVX1_LOC_86/A 0.00fF
C15269 NOR2X1_LOC_742/A NAND2X1_LOC_629/Y 0.01fF
C15270 INVX1_LOC_55/Y NOR2X1_LOC_205/a_36_216# 0.00fF
C15271 INVX1_LOC_265/A NAND2X1_LOC_858/B 0.02fF
C15272 NOR2X1_LOC_651/a_36_216# INVX1_LOC_261/Y 0.00fF
C15273 NAND2X1_LOC_573/Y NOR2X1_LOC_743/Y 0.58fF
C15274 INVX1_LOC_64/A NOR2X1_LOC_814/A 0.11fF
C15275 INVX1_LOC_90/A INVX1_LOC_316/Y 0.03fF
C15276 NOR2X1_LOC_761/Y VDD 0.12fF
C15277 NAND2X1_LOC_254/Y NAND2X1_LOC_99/A 0.00fF
C15278 NAND2X1_LOC_402/B INVX1_LOC_42/A 0.02fF
C15279 NOR2X1_LOC_336/B VDD 0.15fF
C15280 NOR2X1_LOC_593/Y NOR2X1_LOC_66/a_36_216# 0.03fF
C15281 INVX1_LOC_223/A NOR2X1_LOC_137/Y 0.02fF
C15282 NAND2X1_LOC_336/a_36_24# NOR2X1_LOC_536/A 0.00fF
C15283 INVX1_LOC_266/Y NOR2X1_LOC_74/A 0.08fF
C15284 NOR2X1_LOC_82/A INVX1_LOC_9/A 0.03fF
C15285 INVX1_LOC_1/A NOR2X1_LOC_433/Y 0.08fF
C15286 NAND2X1_LOC_35/Y NAND2X1_LOC_489/Y 0.34fF
C15287 NOR2X1_LOC_816/A NOR2X1_LOC_331/B 0.09fF
C15288 INVX1_LOC_134/A INVX1_LOC_9/A 0.03fF
C15289 INVX1_LOC_16/Y INVX1_LOC_3/Y 0.45fF
C15290 NOR2X1_LOC_773/Y INVX1_LOC_102/Y 0.16fF
C15291 INVX1_LOC_224/Y INVX1_LOC_42/A 0.32fF
C15292 INVX1_LOC_101/Y INVX1_LOC_307/A 0.00fF
C15293 INVX1_LOC_294/A NOR2X1_LOC_652/Y 0.00fF
C15294 NAND2X1_LOC_364/A VDD 2.68fF
C15295 INVX1_LOC_310/Y NOR2X1_LOC_78/A 0.01fF
C15296 NAND2X1_LOC_549/Y INVX1_LOC_29/A 0.01fF
C15297 NOR2X1_LOC_552/Y INVX1_LOC_177/A 0.00fF
C15298 NAND2X1_LOC_338/B INVX1_LOC_158/Y 0.14fF
C15299 NOR2X1_LOC_34/B INVX1_LOC_63/A 0.03fF
C15300 NOR2X1_LOC_503/Y NOR2X1_LOC_506/Y 0.02fF
C15301 INVX1_LOC_13/Y NAND2X1_LOC_768/Y 0.02fF
C15302 INVX1_LOC_191/Y INVX1_LOC_6/A 0.00fF
C15303 NAND2X1_LOC_323/B INVX1_LOC_158/Y 0.19fF
C15304 INVX1_LOC_35/A NOR2X1_LOC_89/A 0.09fF
C15305 INVX1_LOC_19/A INVX1_LOC_306/Y 0.03fF
C15306 NOR2X1_LOC_673/A NAND2X1_LOC_473/A 0.07fF
C15307 NOR2X1_LOC_151/Y INVX1_LOC_22/A 0.03fF
C15308 INVX1_LOC_17/A NOR2X1_LOC_216/B 0.09fF
C15309 NAND2X1_LOC_183/a_36_24# INVX1_LOC_307/A 0.01fF
C15310 NAND2X1_LOC_205/A INVX1_LOC_3/Y 0.10fF
C15311 INVX1_LOC_77/A INVX1_LOC_176/A 0.03fF
C15312 NAND2X1_LOC_793/B INVX1_LOC_42/A 0.07fF
C15313 NOR2X1_LOC_409/B NOR2X1_LOC_829/A 0.01fF
C15314 INVX1_LOC_33/A NOR2X1_LOC_324/B 0.01fF
C15315 INVX1_LOC_75/A NAND2X1_LOC_41/Y 0.02fF
C15316 INVX1_LOC_25/A INVX1_LOC_47/Y 0.10fF
C15317 NAND2X1_LOC_181/Y INVX1_LOC_286/A 0.02fF
C15318 NOR2X1_LOC_272/Y INVX1_LOC_133/A 0.23fF
C15319 NAND2X1_LOC_182/A INVX1_LOC_304/A 0.03fF
C15320 INVX1_LOC_132/A INVX1_LOC_37/A 0.15fF
C15321 NAND2X1_LOC_354/B INVX1_LOC_20/A 0.10fF
C15322 NOR2X1_LOC_596/A INVX1_LOC_281/A 0.03fF
C15323 INVX1_LOC_33/A NAND2X1_LOC_211/Y 0.11fF
C15324 NAND2X1_LOC_22/a_36_24# INVX1_LOC_37/A 0.00fF
C15325 INVX1_LOC_29/Y INVX1_LOC_4/Y 0.07fF
C15326 NOR2X1_LOC_52/B NOR2X1_LOC_69/A 0.00fF
C15327 NAND2X1_LOC_514/Y INVX1_LOC_9/A 0.01fF
C15328 D_INPUT_1 NOR2X1_LOC_334/Y 0.07fF
C15329 INVX1_LOC_34/A NOR2X1_LOC_266/B 0.03fF
C15330 INVX1_LOC_40/A INVX1_LOC_315/Y 0.01fF
C15331 NAND2X1_LOC_319/A NOR2X1_LOC_313/Y 0.02fF
C15332 INVX1_LOC_136/A INVX1_LOC_185/A 0.06fF
C15333 INVX1_LOC_63/Y INVX1_LOC_139/Y 0.03fF
C15334 INVX1_LOC_69/Y NOR2X1_LOC_188/Y 0.04fF
C15335 NAND2X1_LOC_859/Y INVX1_LOC_6/A 0.03fF
C15336 NAND2X1_LOC_35/Y INVX1_LOC_32/A 0.03fF
C15337 INPUT_3 NAND2X1_LOC_574/A 0.06fF
C15338 NAND2X1_LOC_390/A INVX1_LOC_286/A 0.10fF
C15339 NOR2X1_LOC_594/Y NAND2X1_LOC_156/B 0.06fF
C15340 INVX1_LOC_30/A INVX1_LOC_179/A 0.02fF
C15341 NOR2X1_LOC_180/B INVX1_LOC_182/A 0.07fF
C15342 NOR2X1_LOC_15/Y NAND2X1_LOC_63/Y 0.03fF
C15343 NOR2X1_LOC_6/B D_INPUT_3 0.25fF
C15344 INVX1_LOC_72/A NAND2X1_LOC_802/Y 0.10fF
C15345 D_INPUT_0 INPUT_0 1.57fF
C15346 NOR2X1_LOC_78/A INVX1_LOC_53/Y 0.06fF
C15347 NOR2X1_LOC_222/Y INVX1_LOC_199/A 0.01fF
C15348 NOR2X1_LOC_557/Y NOR2X1_LOC_440/a_36_216# 0.00fF
C15349 INVX1_LOC_78/A NAND2X1_LOC_793/B 0.01fF
C15350 NAND2X1_LOC_725/B INVX1_LOC_12/A 0.03fF
C15351 NOR2X1_LOC_637/B INVX1_LOC_38/A 0.07fF
C15352 NOR2X1_LOC_220/A INVX1_LOC_247/A 0.01fF
C15353 NOR2X1_LOC_65/B INVX1_LOC_224/Y 0.01fF
C15354 NOR2X1_LOC_355/A INVX1_LOC_285/Y 0.10fF
C15355 INVX1_LOC_182/Y NOR2X1_LOC_755/a_36_216# -0.00fF
C15356 INVX1_LOC_276/Y INVX1_LOC_20/A 0.01fF
C15357 NOR2X1_LOC_601/a_36_216# INVX1_LOC_271/Y 0.01fF
C15358 INVX1_LOC_23/A INVX1_LOC_28/Y 0.01fF
C15359 INVX1_LOC_34/A NAND2X1_LOC_848/A 0.03fF
C15360 NOR2X1_LOC_561/Y NOR2X1_LOC_318/B 0.10fF
C15361 NOR2X1_LOC_627/Y VDD 0.34fF
C15362 INVX1_LOC_90/A INVX1_LOC_86/A 0.03fF
C15363 INVX1_LOC_313/A INVX1_LOC_6/A 0.46fF
C15364 NOR2X1_LOC_209/Y INVX1_LOC_37/A 0.07fF
C15365 NOR2X1_LOC_264/Y INVX1_LOC_38/A 0.07fF
C15366 INVX1_LOC_23/A INVX1_LOC_270/A 0.10fF
C15367 NOR2X1_LOC_400/A NOR2X1_LOC_415/Y 0.01fF
C15368 NAND2X1_LOC_11/Y VDD 0.06fF
C15369 NAND2X1_LOC_390/A INVX1_LOC_95/A 0.14fF
C15370 NAND2X1_LOC_866/B INVX1_LOC_6/A 0.03fF
C15371 INVX1_LOC_10/A NOR2X1_LOC_139/Y 0.10fF
C15372 NAND2X1_LOC_502/a_36_24# INVX1_LOC_78/A 0.00fF
C15373 NOR2X1_LOC_216/a_36_216# INPUT_0 0.01fF
C15374 D_INPUT_2 NOR2X1_LOC_104/a_36_216# 0.00fF
C15375 INVX1_LOC_24/A NOR2X1_LOC_88/Y 0.06fF
C15376 INVX1_LOC_103/A INVX1_LOC_290/Y 0.02fF
C15377 INVX1_LOC_95/Y INVX1_LOC_137/Y 0.03fF
C15378 NOR2X1_LOC_561/Y INVX1_LOC_93/Y 0.02fF
C15379 NOR2X1_LOC_82/Y INVX1_LOC_20/A 0.21fF
C15380 NOR2X1_LOC_103/Y INVX1_LOC_42/A 0.09fF
C15381 INVX1_LOC_27/A INVX1_LOC_94/Y 0.03fF
C15382 NOR2X1_LOC_91/A NOR2X1_LOC_109/Y 0.13fF
C15383 INVX1_LOC_1/A INVX1_LOC_47/Y 0.01fF
C15384 INVX1_LOC_273/Y INVX1_LOC_291/Y 0.02fF
C15385 D_INPUT_0 NAND2X1_LOC_649/B 0.08fF
C15386 INVX1_LOC_93/A NOR2X1_LOC_301/A 0.07fF
C15387 NAND2X1_LOC_33/Y NOR2X1_LOC_629/Y 0.00fF
C15388 INVX1_LOC_10/A NAND2X1_LOC_468/B 0.06fF
C15389 NOR2X1_LOC_507/B NOR2X1_LOC_78/A 0.01fF
C15390 NOR2X1_LOC_550/B NAND2X1_LOC_425/Y 0.02fF
C15391 NOR2X1_LOC_817/Y INVX1_LOC_3/Y 0.03fF
C15392 INVX1_LOC_45/Y NAND2X1_LOC_475/Y 0.01fF
C15393 NOR2X1_LOC_15/Y NAND2X1_LOC_618/Y 0.07fF
C15394 INVX1_LOC_24/A INVX1_LOC_84/A 0.17fF
C15395 NAND2X1_LOC_377/a_36_24# INVX1_LOC_32/A 0.00fF
C15396 INVX1_LOC_34/A INVX1_LOC_46/Y 0.00fF
C15397 NOR2X1_LOC_355/A NOR2X1_LOC_137/B 0.03fF
C15398 INVX1_LOC_225/A NOR2X1_LOC_743/Y 0.02fF
C15399 VDD NOR2X1_LOC_86/A 0.12fF
C15400 NAND2X1_LOC_364/A INVX1_LOC_133/A 0.38fF
C15401 NOR2X1_LOC_634/B NOR2X1_LOC_729/A 0.02fF
C15402 NOR2X1_LOC_68/A INVX1_LOC_272/A 0.07fF
C15403 NOR2X1_LOC_78/B NOR2X1_LOC_729/A 0.06fF
C15404 NAND2X1_LOC_190/Y NOR2X1_LOC_465/Y 0.04fF
C15405 INVX1_LOC_45/A INVX1_LOC_42/A 2.82fF
C15406 INVX1_LOC_48/Y INVX1_LOC_23/Y 0.02fF
C15407 NOR2X1_LOC_568/A INVX1_LOC_42/A 1.75fF
C15408 NAND2X1_LOC_181/Y INVX1_LOC_54/A 0.01fF
C15409 INVX1_LOC_311/A INVX1_LOC_206/Y 0.05fF
C15410 NOR2X1_LOC_557/Y INVX1_LOC_84/A 0.07fF
C15411 NOR2X1_LOC_103/Y INVX1_LOC_78/A 0.05fF
C15412 INVX1_LOC_83/A NAND2X1_LOC_637/a_36_24# 0.07fF
C15413 NAND2X1_LOC_151/a_36_24# INVX1_LOC_94/Y 0.00fF
C15414 NOR2X1_LOC_96/Y INVX1_LOC_316/Y 0.10fF
C15415 NOR2X1_LOC_590/A INVX1_LOC_4/A 0.03fF
C15416 INVX1_LOC_159/A INVX1_LOC_109/Y 0.02fF
C15417 NOR2X1_LOC_92/Y NAND2X1_LOC_97/a_36_24# 0.00fF
C15418 NAND2X1_LOC_538/a_36_24# NAND2X1_LOC_649/B 0.01fF
C15419 INVX1_LOC_125/Y NOR2X1_LOC_9/Y 0.05fF
C15420 INVX1_LOC_49/A INVX1_LOC_49/Y 0.10fF
C15421 NOR2X1_LOC_706/A NOR2X1_LOC_486/Y 0.18fF
C15422 NOR2X1_LOC_544/A INVX1_LOC_307/A 0.20fF
C15423 NAND2X1_LOC_348/A NOR2X1_LOC_346/Y 0.01fF
C15424 INVX1_LOC_89/A INVX1_LOC_12/Y 0.03fF
C15425 D_INPUT_7 D_INPUT_5 0.11fF
C15426 NOR2X1_LOC_93/Y NOR2X1_LOC_392/Y 0.02fF
C15427 NAND2X1_LOC_465/Y NAND2X1_LOC_489/Y 0.03fF
C15428 NOR2X1_LOC_234/Y NAND2X1_LOC_489/Y 0.02fF
C15429 NOR2X1_LOC_65/B NOR2X1_LOC_103/Y 0.10fF
C15430 NAND2X1_LOC_722/A INVX1_LOC_250/Y 0.06fF
C15431 NAND2X1_LOC_848/Y INVX1_LOC_316/Y 0.11fF
C15432 INVX1_LOC_71/A INVX1_LOC_42/A 0.07fF
C15433 INVX1_LOC_49/A INVX1_LOC_99/A 0.03fF
C15434 NOR2X1_LOC_714/a_36_216# NOR2X1_LOC_78/A 0.00fF
C15435 INVX1_LOC_306/A INVX1_LOC_9/A 0.01fF
C15436 NOR2X1_LOC_205/Y INVX1_LOC_29/Y 0.00fF
C15437 INVX1_LOC_45/A INVX1_LOC_78/A 0.13fF
C15438 INVX1_LOC_83/A NOR2X1_LOC_729/A 0.06fF
C15439 INVX1_LOC_143/A INVX1_LOC_84/A 0.19fF
C15440 INVX1_LOC_50/A NOR2X1_LOC_107/Y 0.05fF
C15441 INVX1_LOC_61/Y INVX1_LOC_26/A 0.09fF
C15442 NAND2X1_LOC_850/Y INVX1_LOC_265/Y 0.01fF
C15443 INVX1_LOC_24/A INVX1_LOC_15/A 8.83fF
C15444 NOR2X1_LOC_568/A INVX1_LOC_78/A 0.07fF
C15445 INVX1_LOC_94/A INVX1_LOC_32/A 0.07fF
C15446 INVX1_LOC_77/A NOR2X1_LOC_116/a_36_216# -0.01fF
C15447 NOR2X1_LOC_526/Y NOR2X1_LOC_485/Y 0.01fF
C15448 INVX1_LOC_269/A NOR2X1_LOC_392/Y 0.41fF
C15449 NOR2X1_LOC_272/Y NOR2X1_LOC_510/Y 0.08fF
C15450 NOR2X1_LOC_286/Y INVX1_LOC_53/A 0.00fF
C15451 INPUT_0 NOR2X1_LOC_266/B 0.03fF
C15452 INVX1_LOC_2/A INVX1_LOC_49/Y 4.62fF
C15453 INVX1_LOC_35/A INVX1_LOC_224/A 0.03fF
C15454 INVX1_LOC_30/A NOR2X1_LOC_693/Y 0.07fF
C15455 NOR2X1_LOC_195/A NOR2X1_LOC_598/B 0.03fF
C15456 INVX1_LOC_34/A NOR2X1_LOC_754/A 0.04fF
C15457 INVX1_LOC_95/Y INVX1_LOC_91/A 3.02fF
C15458 NOR2X1_LOC_91/A INVX1_LOC_36/A 0.27fF
C15459 INVX1_LOC_35/A INVX1_LOC_11/A 0.16fF
C15460 NOR2X1_LOC_65/B INVX1_LOC_45/A 0.06fF
C15461 NOR2X1_LOC_226/A INVX1_LOC_49/Y 0.03fF
C15462 INPUT_0 NOR2X1_LOC_859/Y 0.01fF
C15463 INVX1_LOC_205/Y INVX1_LOC_27/A 0.03fF
C15464 INVX1_LOC_230/Y NAND2X1_LOC_571/B 0.11fF
C15465 NAND2X1_LOC_793/Y NOR2X1_LOC_129/a_36_216# 0.02fF
C15466 NAND2X1_LOC_721/A NOR2X1_LOC_167/Y 0.02fF
C15467 NAND2X1_LOC_103/a_36_24# INVX1_LOC_46/A 0.01fF
C15468 NOR2X1_LOC_255/Y INVX1_LOC_61/Y 0.02fF
C15469 INVX1_LOC_21/A NOR2X1_LOC_92/Y 0.17fF
C15470 INVX1_LOC_64/A NAND2X1_LOC_803/B 0.02fF
C15471 NOR2X1_LOC_848/Y INVX1_LOC_5/A 0.26fF
C15472 NOR2X1_LOC_607/Y NOR2X1_LOC_334/Y 0.01fF
C15473 NOR2X1_LOC_91/A NOR2X1_LOC_267/A 0.56fF
C15474 INVX1_LOC_71/A INVX1_LOC_78/A 0.32fF
C15475 NOR2X1_LOC_605/B NOR2X1_LOC_605/A 0.04fF
C15476 NAND2X1_LOC_552/a_36_24# INVX1_LOC_84/A 0.00fF
C15477 NOR2X1_LOC_318/B INVX1_LOC_76/A 0.01fF
C15478 INVX1_LOC_226/A NAND2X1_LOC_63/Y 0.03fF
C15479 NOR2X1_LOC_315/Y INVX1_LOC_170/Y 0.01fF
C15480 INVX1_LOC_90/A NOR2X1_LOC_510/B 0.25fF
C15481 INVX1_LOC_223/Y INVX1_LOC_269/A 0.09fF
C15482 INPUT_0 NAND2X1_LOC_848/A 0.10fF
C15483 NOR2X1_LOC_305/Y INVX1_LOC_91/A 0.07fF
C15484 INVX1_LOC_308/Y NOR2X1_LOC_652/Y 0.03fF
C15485 INVX1_LOC_17/A INVX1_LOC_93/A 0.07fF
C15486 NOR2X1_LOC_100/A NOR2X1_LOC_861/Y 0.08fF
C15487 NOR2X1_LOC_272/Y NOR2X1_LOC_361/B 0.03fF
C15488 INVX1_LOC_36/A INVX1_LOC_23/A 8.05fF
C15489 INVX1_LOC_18/A NOR2X1_LOC_654/A 0.49fF
C15490 NOR2X1_LOC_321/Y NAND2X1_LOC_326/A 0.06fF
C15491 INVX1_LOC_64/A NOR2X1_LOC_590/A 2.53fF
C15492 INVX1_LOC_55/Y NOR2X1_LOC_155/A 0.03fF
C15493 INVX1_LOC_93/Y INVX1_LOC_76/A 0.10fF
C15494 NAND2X1_LOC_502/a_36_24# NOR2X1_LOC_503/Y 0.01fF
C15495 NOR2X1_LOC_242/A NOR2X1_LOC_286/Y 0.15fF
C15496 NOR2X1_LOC_349/A VDD 0.12fF
C15497 NAND2X1_LOC_214/B INVX1_LOC_293/A 0.01fF
C15498 NOR2X1_LOC_45/B NOR2X1_LOC_447/B 0.00fF
C15499 NOR2X1_LOC_163/A INVX1_LOC_107/Y 0.00fF
C15500 INVX1_LOC_64/A INVX1_LOC_22/Y 0.03fF
C15501 NOR2X1_LOC_130/A INVX1_LOC_84/A 1.33fF
C15502 NOR2X1_LOC_405/A VDD 1.83fF
C15503 INVX1_LOC_45/A INVX1_LOC_152/Y 0.24fF
C15504 INVX1_LOC_11/Y NOR2X1_LOC_305/Y 0.02fF
C15505 NOR2X1_LOC_65/B INVX1_LOC_71/A 0.20fF
C15506 INVX1_LOC_136/A NOR2X1_LOC_754/Y 0.08fF
C15507 NOR2X1_LOC_557/A NAND2X1_LOC_96/A 0.02fF
C15508 NOR2X1_LOC_419/Y NOR2X1_LOC_843/B 0.03fF
C15509 NAND2X1_LOC_361/Y NAND2X1_LOC_616/a_36_24# 0.00fF
C15510 NOR2X1_LOC_264/Y NAND2X1_LOC_223/A 0.12fF
C15511 NOR2X1_LOC_637/Y NOR2X1_LOC_654/A 0.00fF
C15512 NOR2X1_LOC_590/A NOR2X1_LOC_436/a_36_216# 0.00fF
C15513 INVX1_LOC_18/A INVX1_LOC_58/Y 0.02fF
C15514 INVX1_LOC_143/A INVX1_LOC_15/A 0.09fF
C15515 INVX1_LOC_145/A INVX1_LOC_23/A 0.02fF
C15516 NOR2X1_LOC_163/Y INVX1_LOC_113/A 0.08fF
C15517 NOR2X1_LOC_188/Y NOR2X1_LOC_89/A 0.15fF
C15518 NAND2X1_LOC_650/B INVX1_LOC_20/A 0.09fF
C15519 INVX1_LOC_216/Y INVX1_LOC_1/A 0.03fF
C15520 D_INPUT_0 NOR2X1_LOC_84/B 0.02fF
C15521 INVX1_LOC_139/A INVX1_LOC_76/A 0.16fF
C15522 NOR2X1_LOC_326/Y NOR2X1_LOC_777/B 0.05fF
C15523 INVX1_LOC_90/A NOR2X1_LOC_662/A 0.03fF
C15524 NOR2X1_LOC_136/Y INVX1_LOC_32/A 0.06fF
C15525 INPUT_0 INVX1_LOC_46/Y 0.02fF
C15526 INVX1_LOC_68/Y INVX1_LOC_15/A 0.01fF
C15527 INVX1_LOC_56/A INVX1_LOC_32/A 0.29fF
C15528 INVX1_LOC_278/A INVX1_LOC_24/A 0.07fF
C15529 VDD NOR2X1_LOC_857/A 0.12fF
C15530 NAND2X1_LOC_648/A INVX1_LOC_49/Y 0.03fF
C15531 NAND2X1_LOC_634/Y NOR2X1_LOC_291/Y 0.67fF
C15532 NOR2X1_LOC_91/A NOR2X1_LOC_309/Y 0.10fF
C15533 NAND2X1_LOC_56/a_36_24# INVX1_LOC_1/A 0.00fF
C15534 INVX1_LOC_17/A NOR2X1_LOC_513/Y 0.01fF
C15535 NOR2X1_LOC_772/Y INVX1_LOC_57/A 0.54fF
C15536 NOR2X1_LOC_804/B INVX1_LOC_23/A 0.46fF
C15537 NOR2X1_LOC_84/Y INVX1_LOC_23/Y 0.19fF
C15538 INVX1_LOC_96/Y NOR2X1_LOC_631/Y 0.08fF
C15539 NAND2X1_LOC_469/B INVX1_LOC_281/A 0.00fF
C15540 NOR2X1_LOC_356/A INVX1_LOC_19/A 0.09fF
C15541 NOR2X1_LOC_175/A NOR2X1_LOC_541/B 0.22fF
C15542 NOR2X1_LOC_82/Y INVX1_LOC_4/A 0.32fF
C15543 NOR2X1_LOC_231/B INVX1_LOC_1/A 0.02fF
C15544 NOR2X1_LOC_349/A NAND2X1_LOC_41/a_36_24# 0.01fF
C15545 NOR2X1_LOC_392/B INVX1_LOC_57/A 0.09fF
C15546 NOR2X1_LOC_251/Y INVX1_LOC_94/Y 0.00fF
C15547 INVX1_LOC_35/A NOR2X1_LOC_433/A 0.10fF
C15548 INVX1_LOC_233/A NOR2X1_LOC_753/Y 0.08fF
C15549 NAND2X1_LOC_793/Y NAND2X1_LOC_807/A 0.01fF
C15550 NOR2X1_LOC_186/Y NAND2X1_LOC_198/B 0.10fF
C15551 NAND2X1_LOC_9/Y NOR2X1_LOC_520/B 0.04fF
C15552 NOR2X1_LOC_553/Y NOR2X1_LOC_334/Y 0.02fF
C15553 INVX1_LOC_35/A NOR2X1_LOC_593/Y 0.09fF
C15554 NOR2X1_LOC_309/Y INVX1_LOC_23/A 0.03fF
C15555 NOR2X1_LOC_564/Y INVX1_LOC_29/A 0.03fF
C15556 NAND2X1_LOC_642/Y NOR2X1_LOC_743/Y 0.03fF
C15557 INVX1_LOC_50/A INVX1_LOC_149/A 0.39fF
C15558 INVX1_LOC_101/A INVX1_LOC_4/Y 0.02fF
C15559 INVX1_LOC_227/A INVX1_LOC_4/A 0.42fF
C15560 NOR2X1_LOC_92/Y NAND2X1_LOC_354/Y 0.02fF
C15561 INVX1_LOC_14/Y NOR2X1_LOC_684/Y 0.26fF
C15562 INVX1_LOC_254/A INVX1_LOC_50/Y 0.06fF
C15563 NOR2X1_LOC_375/Y INVX1_LOC_175/A 0.01fF
C15564 NOR2X1_LOC_130/A INVX1_LOC_15/A 0.06fF
C15565 INVX1_LOC_64/A NAND2X1_LOC_354/B 0.03fF
C15566 NAND2X1_LOC_573/Y NAND2X1_LOC_198/B 0.10fF
C15567 NOR2X1_LOC_68/A INVX1_LOC_198/A -0.01fF
C15568 NOR2X1_LOC_74/A INVX1_LOC_19/A 0.13fF
C15569 INVX1_LOC_147/A INVX1_LOC_272/A 0.02fF
C15570 NOR2X1_LOC_824/Y NOR2X1_LOC_823/a_36_216# 0.00fF
C15571 NOR2X1_LOC_232/Y NOR2X1_LOC_86/Y 0.10fF
C15572 NOR2X1_LOC_314/Y INVX1_LOC_54/A 0.02fF
C15573 INVX1_LOC_35/A NOR2X1_LOC_52/B 0.06fF
C15574 NOR2X1_LOC_361/B NAND2X1_LOC_364/A 1.25fF
C15575 NOR2X1_LOC_355/A INVX1_LOC_4/Y 0.01fF
C15576 NOR2X1_LOC_9/Y INVX1_LOC_19/A 0.03fF
C15577 INVX1_LOC_238/A INVX1_LOC_238/Y 0.20fF
C15578 NOR2X1_LOC_267/a_36_216# INVX1_LOC_181/Y 0.01fF
C15579 INVX1_LOC_115/A INVX1_LOC_92/A 0.01fF
C15580 INVX1_LOC_76/A INVX1_LOC_117/Y 0.02fF
C15581 INVX1_LOC_313/Y NOR2X1_LOC_609/Y 0.03fF
C15582 INVX1_LOC_110/Y NAND2X1_LOC_206/a_36_24# 0.01fF
C15583 NAND2X1_LOC_9/Y NOR2X1_LOC_67/A 0.09fF
C15584 INVX1_LOC_21/A INVX1_LOC_41/A 4.44fF
C15585 NOR2X1_LOC_75/Y INVX1_LOC_18/A 0.04fF
C15586 INVX1_LOC_36/A NAND2X1_LOC_509/a_36_24# 0.00fF
C15587 NOR2X1_LOC_123/B INVX1_LOC_78/A 0.00fF
C15588 INVX1_LOC_95/Y NOR2X1_LOC_179/Y 0.03fF
C15589 INVX1_LOC_54/A INVX1_LOC_117/A 1.16fF
C15590 INVX1_LOC_21/A INVX1_LOC_201/Y 0.21fF
C15591 INVX1_LOC_36/A INVX1_LOC_31/A 0.22fF
C15592 INVX1_LOC_276/Y INVX1_LOC_64/A 0.01fF
C15593 NAND2X1_LOC_703/Y NAND2X1_LOC_325/Y 0.07fF
C15594 NOR2X1_LOC_577/a_36_216# NOR2X1_LOC_383/B 0.00fF
C15595 NAND2X1_LOC_563/A NOR2X1_LOC_392/Y 0.12fF
C15596 NAND2X1_LOC_725/B NAND2X1_LOC_787/B 0.07fF
C15597 INVX1_LOC_256/A NOR2X1_LOC_273/Y 0.02fF
C15598 INVX1_LOC_269/A NOR2X1_LOC_554/a_36_216# 0.01fF
C15599 NOR2X1_LOC_641/B INVX1_LOC_30/A 0.03fF
C15600 NAND2X1_LOC_579/A NAND2X1_LOC_833/Y 0.06fF
C15601 INVX1_LOC_103/A INVX1_LOC_77/A 0.07fF
C15602 INVX1_LOC_256/A NOR2X1_LOC_759/Y 0.53fF
C15603 INVX1_LOC_256/A NOR2X1_LOC_274/a_36_216# 0.00fF
C15604 INVX1_LOC_21/A NAND2X1_LOC_477/A 0.01fF
C15605 INVX1_LOC_27/A NOR2X1_LOC_315/Y 0.90fF
C15606 NOR2X1_LOC_45/Y NAND2X1_LOC_198/B 0.10fF
C15607 INVX1_LOC_256/A INVX1_LOC_202/A 0.00fF
C15608 NOR2X1_LOC_67/A NAND2X1_LOC_553/A 0.04fF
C15609 INVX1_LOC_144/A INVX1_LOC_32/A 0.08fF
C15610 NOR2X1_LOC_299/Y INVX1_LOC_173/A 0.05fF
C15611 NOR2X1_LOC_405/A INVX1_LOC_133/A 0.02fF
C15612 NOR2X1_LOC_751/Y INVX1_LOC_30/A 0.00fF
C15613 INVX1_LOC_13/A NOR2X1_LOC_598/B 0.91fF
C15614 INVX1_LOC_14/A NOR2X1_LOC_561/a_36_216# 0.00fF
C15615 INVX1_LOC_310/A INVX1_LOC_27/A 0.49fF
C15616 NOR2X1_LOC_188/A INVX1_LOC_47/Y 0.40fF
C15617 NOR2X1_LOC_432/Y INVX1_LOC_27/A 0.03fF
C15618 INVX1_LOC_13/A INVX1_LOC_51/A 0.01fF
C15619 INVX1_LOC_292/A INVX1_LOC_77/A 0.10fF
C15620 NAND2X1_LOC_33/Y INVX1_LOC_269/A -0.00fF
C15621 NOR2X1_LOC_510/Y NOR2X1_LOC_289/a_36_216# 0.01fF
C15622 INVX1_LOC_45/Y INVX1_LOC_30/A 0.07fF
C15623 INVX1_LOC_226/Y INVX1_LOC_13/Y 0.01fF
C15624 NAND2X1_LOC_656/Y NOR2X1_LOC_717/A 0.10fF
C15625 INVX1_LOC_5/A NAND2X1_LOC_479/Y 0.07fF
C15626 NOR2X1_LOC_476/Y NOR2X1_LOC_480/A 0.14fF
C15627 INVX1_LOC_90/A INVX1_LOC_57/A 0.29fF
C15628 NAND2X1_LOC_468/B INVX1_LOC_12/A 0.06fF
C15629 NOR2X1_LOC_13/Y INVX1_LOC_312/Y 0.00fF
C15630 NOR2X1_LOC_186/Y INVX1_LOC_53/Y 0.07fF
C15631 INVX1_LOC_224/A NAND2X1_LOC_667/a_36_24# 0.00fF
C15632 INVX1_LOC_196/Y NOR2X1_LOC_858/A 0.16fF
C15633 NAND2X1_LOC_555/Y NAND2X1_LOC_5/a_36_24# 0.00fF
C15634 NAND2X1_LOC_787/A NOR2X1_LOC_71/Y 0.02fF
C15635 NOR2X1_LOC_389/B INVX1_LOC_57/A 0.32fF
C15636 NOR2X1_LOC_848/a_36_216# NOR2X1_LOC_516/B 0.00fF
C15637 INVX1_LOC_278/A NOR2X1_LOC_130/A 0.07fF
C15638 INVX1_LOC_45/A NOR2X1_LOC_152/Y 0.07fF
C15639 INVX1_LOC_21/A NOR2X1_LOC_211/A 0.02fF
C15640 NAND2X1_LOC_861/Y NAND2X1_LOC_793/B 1.06fF
C15641 NOR2X1_LOC_728/B INVX1_LOC_271/Y 0.09fF
C15642 INVX1_LOC_37/A NOR2X1_LOC_48/Y 0.01fF
C15643 INVX1_LOC_17/A INVX1_LOC_54/Y 0.03fF
C15644 NAND2X1_LOC_856/A NOR2X1_LOC_152/Y 0.03fF
C15645 INVX1_LOC_232/Y INVX1_LOC_14/A 0.02fF
C15646 INVX1_LOC_24/A NOR2X1_LOC_168/Y 0.03fF
C15647 INVX1_LOC_230/Y INVX1_LOC_219/Y 0.05fF
C15648 NAND2X1_LOC_364/A INVX1_LOC_184/Y 0.04fF
C15649 NOR2X1_LOC_286/Y NOR2X1_LOC_634/B 0.36fF
C15650 NAND2X1_LOC_552/A INVX1_LOC_135/A 0.08fF
C15651 NOR2X1_LOC_658/Y NOR2X1_LOC_219/B 0.02fF
C15652 NOR2X1_LOC_598/B INVX1_LOC_55/Y 0.08fF
C15653 NAND2X1_LOC_213/A NAND2X1_LOC_162/A 0.04fF
C15654 NOR2X1_LOC_458/B NAND2X1_LOC_190/Y 0.06fF
C15655 INVX1_LOC_49/A NOR2X1_LOC_722/Y 0.01fF
C15656 INVX1_LOC_48/Y INVX1_LOC_232/A 0.00fF
C15657 INVX1_LOC_245/Y INVX1_LOC_266/Y 0.35fF
C15658 NOR2X1_LOC_706/A INVX1_LOC_275/Y 0.04fF
C15659 INVX1_LOC_5/A INVX1_LOC_135/A 0.41fF
C15660 INVX1_LOC_75/Y NAND2X1_LOC_425/Y 0.03fF
C15661 NOR2X1_LOC_644/B NOR2X1_LOC_348/B 0.00fF
C15662 NOR2X1_LOC_537/A INVX1_LOC_18/A 0.00fF
C15663 NAND2X1_LOC_708/Y NOR2X1_LOC_224/a_36_216# 0.00fF
C15664 NAND2X1_LOC_689/a_36_24# NAND2X1_LOC_361/Y 0.00fF
C15665 VDD INVX1_LOC_109/Y 0.87fF
C15666 INVX1_LOC_196/Y INVX1_LOC_292/Y 0.00fF
C15667 NAND2X1_LOC_348/A INVX1_LOC_57/A 0.03fF
C15668 INVX1_LOC_176/A NOR2X1_LOC_861/Y 0.03fF
C15669 NOR2X1_LOC_9/Y INVX1_LOC_26/Y 0.02fF
C15670 NOR2X1_LOC_716/B INVX1_LOC_18/A 0.08fF
C15671 INVX1_LOC_91/A INVX1_LOC_271/Y 0.07fF
C15672 NAND2X1_LOC_392/A INVX1_LOC_14/A 0.01fF
C15673 NOR2X1_LOC_232/Y INVX1_LOC_25/Y 0.14fF
C15674 NOR2X1_LOC_498/a_36_216# INVX1_LOC_217/A -0.02fF
C15675 NOR2X1_LOC_92/Y NOR2X1_LOC_521/Y 0.04fF
C15676 NOR2X1_LOC_401/B NOR2X1_LOC_160/B 0.06fF
C15677 INVX1_LOC_135/A INVX1_LOC_178/A 0.10fF
C15678 NAND2X1_LOC_807/Y NOR2X1_LOC_109/Y 0.04fF
C15679 NOR2X1_LOC_536/A NAND2X1_LOC_74/B 0.20fF
C15680 INVX1_LOC_64/A NOR2X1_LOC_703/A 0.03fF
C15681 NOR2X1_LOC_590/A INVX1_LOC_44/Y 0.10fF
C15682 NOR2X1_LOC_68/A NOR2X1_LOC_770/B 0.00fF
C15683 NOR2X1_LOC_402/a_36_216# NOR2X1_LOC_160/B 0.00fF
C15684 NAND2X1_LOC_98/a_36_24# INVX1_LOC_234/A 0.01fF
C15685 NOR2X1_LOC_121/Y INVX1_LOC_72/Y 0.19fF
C15686 INVX1_LOC_6/A INVX1_LOC_270/A 0.07fF
C15687 INVX1_LOC_289/Y NOR2X1_LOC_561/Y 0.04fF
C15688 INVX1_LOC_71/A INVX1_LOC_113/Y 0.03fF
C15689 NAND2X1_LOC_21/Y INVX1_LOC_24/A 0.02fF
C15690 INVX1_LOC_78/Y NOR2X1_LOC_727/B 0.00fF
C15691 NOR2X1_LOC_280/Y INVX1_LOC_15/A 0.01fF
C15692 INVX1_LOC_49/Y INVX1_LOC_118/A 0.03fF
C15693 NAND2X1_LOC_214/Y INVX1_LOC_83/A 0.03fF
C15694 NOR2X1_LOC_48/B INVX1_LOC_117/A 0.14fF
C15695 NAND2X1_LOC_655/A NOR2X1_LOC_686/A 0.05fF
C15696 NAND2X1_LOC_93/B INVX1_LOC_293/Y 0.03fF
C15697 INVX1_LOC_24/A NAND2X1_LOC_464/Y 0.02fF
C15698 INVX1_LOC_225/A NAND2X1_LOC_198/B 0.01fF
C15699 INVX1_LOC_205/A NOR2X1_LOC_87/B 0.45fF
C15700 INVX1_LOC_243/A NAND2X1_LOC_36/A 0.00fF
C15701 NOR2X1_LOC_340/A INVX1_LOC_9/A 0.05fF
C15702 INVX1_LOC_88/A INVX1_LOC_10/A 0.13fF
C15703 INVX1_LOC_58/A INVX1_LOC_286/A 0.07fF
C15704 INVX1_LOC_172/A NOR2X1_LOC_716/B 0.07fF
C15705 INVX1_LOC_36/A INVX1_LOC_191/Y 0.00fF
C15706 NOR2X1_LOC_262/Y NOR2X1_LOC_557/Y 0.04fF
C15707 INVX1_LOC_5/A NOR2X1_LOC_202/Y 0.05fF
C15708 INVX1_LOC_20/Y NAND2X1_LOC_473/A 0.02fF
C15709 NOR2X1_LOC_309/Y INVX1_LOC_111/A 0.01fF
C15710 NOR2X1_LOC_331/B INVX1_LOC_42/A 0.03fF
C15711 NOR2X1_LOC_644/B INVX1_LOC_22/A 0.03fF
C15712 INVX1_LOC_87/Y NOR2X1_LOC_440/B 0.03fF
C15713 INVX1_LOC_178/A NOR2X1_LOC_490/Y 0.01fF
C15714 NOR2X1_LOC_848/Y NOR2X1_LOC_332/A 0.22fF
C15715 NOR2X1_LOC_82/A INVX1_LOC_7/A 0.01fF
C15716 INVX1_LOC_34/A INVX1_LOC_49/A 0.03fF
C15717 INVX1_LOC_103/A INVX1_LOC_190/A 0.04fF
C15718 NOR2X1_LOC_68/A NOR2X1_LOC_87/Y 0.25fF
C15719 INVX1_LOC_33/A INVX1_LOC_155/A 0.97fF
C15720 NAND2X1_LOC_93/B NAND2X1_LOC_74/B 0.10fF
C15721 NOR2X1_LOC_500/Y NOR2X1_LOC_500/B 0.01fF
C15722 NAND2X1_LOC_116/A NOR2X1_LOC_350/A 0.58fF
C15723 INVX1_LOC_5/A NOR2X1_LOC_391/B 0.02fF
C15724 NOR2X1_LOC_78/B INVX1_LOC_181/Y 0.07fF
C15725 INVX1_LOC_135/A NOR2X1_LOC_816/A 0.36fF
C15726 INVX1_LOC_293/Y INVX1_LOC_3/A 0.07fF
C15727 NOR2X1_LOC_647/a_36_216# NOR2X1_LOC_332/A 0.01fF
C15728 NAND2X1_LOC_733/Y NOR2X1_LOC_298/Y 0.03fF
C15729 NOR2X1_LOC_751/A NAND2X1_LOC_63/a_36_24# 0.00fF
C15730 NOR2X1_LOC_640/Y NOR2X1_LOC_640/B 0.06fF
C15731 NOR2X1_LOC_205/Y NOR2X1_LOC_736/Y 0.00fF
C15732 NOR2X1_LOC_262/Y INVX1_LOC_143/A 0.02fF
C15733 NOR2X1_LOC_644/A NOR2X1_LOC_457/A 0.03fF
C15734 NOR2X1_LOC_160/B INVX1_LOC_89/A 0.80fF
C15735 NAND2X1_LOC_231/Y INVX1_LOC_49/A 0.01fF
C15736 NAND2X1_LOC_731/a_36_24# INVX1_LOC_72/A 0.01fF
C15737 NOR2X1_LOC_589/A INVX1_LOC_177/Y 0.03fF
C15738 NOR2X1_LOC_863/B NOR2X1_LOC_863/A 0.02fF
C15739 INVX1_LOC_249/A INVX1_LOC_52/A 0.02fF
C15740 INVX1_LOC_269/A INVX1_LOC_75/A 0.29fF
C15741 NAND2X1_LOC_74/B INVX1_LOC_3/A 0.15fF
C15742 NOR2X1_LOC_52/B NOR2X1_LOC_365/a_36_216# 0.00fF
C15743 INVX1_LOC_78/A NOR2X1_LOC_331/B 0.20fF
C15744 NAND2X1_LOC_860/Y INVX1_LOC_71/A 0.05fF
C15745 NAND2X1_LOC_563/Y INVX1_LOC_80/Y 0.06fF
C15746 INVX1_LOC_2/A INVX1_LOC_34/A 0.14fF
C15747 NOR2X1_LOC_751/a_36_216# NOR2X1_LOC_9/Y 0.00fF
C15748 INVX1_LOC_46/A NAND2X1_LOC_787/Y 0.00fF
C15749 NOR2X1_LOC_160/B NAND2X1_LOC_508/A 0.01fF
C15750 NOR2X1_LOC_27/Y INVX1_LOC_240/A 0.03fF
C15751 INVX1_LOC_30/A NOR2X1_LOC_71/Y 0.10fF
C15752 INVX1_LOC_5/A NOR2X1_LOC_552/A 0.07fF
C15753 NOR2X1_LOC_639/a_36_216# INVX1_LOC_72/A 0.00fF
C15754 INVX1_LOC_35/A INVX1_LOC_74/A 0.00fF
C15755 INVX1_LOC_41/A NOR2X1_LOC_667/A 0.03fF
C15756 NAND2X1_LOC_208/B INPUT_1 0.16fF
C15757 NOR2X1_LOC_155/A INVX1_LOC_32/A 0.03fF
C15758 NOR2X1_LOC_274/Y INVX1_LOC_1/Y 0.02fF
C15759 NOR2X1_LOC_226/A INVX1_LOC_34/A 0.07fF
C15760 NOR2X1_LOC_649/B NOR2X1_LOC_847/B -0.03fF
C15761 INVX1_LOC_181/Y NAND2X1_LOC_392/Y 0.01fF
C15762 NOR2X1_LOC_498/Y NOR2X1_LOC_667/A -0.01fF
C15763 NOR2X1_LOC_717/B INVX1_LOC_18/A 0.03fF
C15764 NOR2X1_LOC_197/B INVX1_LOC_15/A 0.10fF
C15765 INVX1_LOC_36/A INVX1_LOC_313/A 0.11fF
C15766 NOR2X1_LOC_521/Y NAND2X1_LOC_837/Y 0.01fF
C15767 INVX1_LOC_286/Y NOR2X1_LOC_597/A 0.02fF
C15768 NOR2X1_LOC_496/Y NOR2X1_LOC_45/B 0.01fF
C15769 INVX1_LOC_36/A NAND2X1_LOC_866/B 0.07fF
C15770 NAND2X1_LOC_656/a_36_24# INVX1_LOC_18/A 0.00fF
C15771 NOR2X1_LOC_644/A INVX1_LOC_30/A 0.03fF
C15772 INVX1_LOC_233/A NOR2X1_LOC_558/A 0.03fF
C15773 NOR2X1_LOC_392/Y NOR2X1_LOC_37/a_36_216# 0.01fF
C15774 NAND2X1_LOC_849/B INVX1_LOC_57/A 0.98fF
C15775 INVX1_LOC_134/A NOR2X1_LOC_835/B 0.00fF
C15776 INVX1_LOC_34/A NOR2X1_LOC_218/Y 0.00fF
C15777 INVX1_LOC_36/A NAND2X1_LOC_807/Y 0.76fF
C15778 INVX1_LOC_2/A NAND2X1_LOC_231/Y 0.10fF
C15779 NAND2X1_LOC_139/A INVX1_LOC_16/A 0.02fF
C15780 INVX1_LOC_57/A INVX1_LOC_38/A 0.13fF
C15781 NOR2X1_LOC_216/B INVX1_LOC_94/Y 0.20fF
C15782 INVX1_LOC_201/Y NAND2X1_LOC_6/a_36_24# 0.00fF
C15783 INVX1_LOC_12/Y NOR2X1_LOC_392/Y 0.00fF
C15784 INVX1_LOC_41/A NOR2X1_LOC_729/a_36_216# 0.00fF
C15785 INVX1_LOC_225/A INVX1_LOC_53/Y 0.01fF
C15786 INVX1_LOC_174/Y NOR2X1_LOC_379/a_36_216# 0.00fF
C15787 INVX1_LOC_145/A INVX1_LOC_313/A 0.03fF
C15788 NAND2X1_LOC_861/Y INVX1_LOC_71/A 0.06fF
C15789 INVX1_LOC_247/Y NOR2X1_LOC_564/Y 0.02fF
C15790 NOR2X1_LOC_643/Y D_INPUT_0 0.00fF
C15791 NOR2X1_LOC_92/Y INVX1_LOC_304/A 0.46fF
C15792 INVX1_LOC_34/A NAND2X1_LOC_664/a_36_24# 0.00fF
C15793 INVX1_LOC_204/Y INVX1_LOC_37/A 0.01fF
C15794 NOR2X1_LOC_220/a_36_216# NOR2X1_LOC_389/B 0.00fF
C15795 NOR2X1_LOC_160/B NOR2X1_LOC_703/Y 0.21fF
C15796 INVX1_LOC_208/A NOR2X1_LOC_493/B 0.16fF
C15797 INVX1_LOC_34/A NAND2X1_LOC_462/B 0.00fF
C15798 INVX1_LOC_120/A INVX1_LOC_77/A 0.03fF
C15799 INVX1_LOC_49/A NOR2X1_LOC_148/B 0.10fF
C15800 NAND2X1_LOC_740/Y VDD 0.11fF
C15801 INVX1_LOC_35/A NAND2X1_LOC_699/a_36_24# 0.00fF
C15802 INVX1_LOC_232/A NOR2X1_LOC_84/Y 0.02fF
C15803 NOR2X1_LOC_361/B NOR2X1_LOC_405/A 0.10fF
C15804 NOR2X1_LOC_751/A INVX1_LOC_30/A 0.00fF
C15805 NOR2X1_LOC_340/A NOR2X1_LOC_861/Y 0.13fF
C15806 INVX1_LOC_58/A INVX1_LOC_54/A 0.64fF
C15807 INVX1_LOC_174/A INVX1_LOC_86/Y 0.03fF
C15808 NOR2X1_LOC_92/Y NOR2X1_LOC_670/Y 0.01fF
C15809 NOR2X1_LOC_151/Y INVX1_LOC_18/A 0.07fF
C15810 NAND2X1_LOC_364/Y INVX1_LOC_132/Y 0.03fF
C15811 NAND2X1_LOC_725/A NOR2X1_LOC_692/Y 0.05fF
C15812 NOR2X1_LOC_203/Y NOR2X1_LOC_500/Y 0.03fF
C15813 NAND2X1_LOC_579/A NAND2X1_LOC_241/Y 0.07fF
C15814 INVX1_LOC_15/Y NAND2X1_LOC_735/B 0.03fF
C15815 INVX1_LOC_289/Y INVX1_LOC_76/A 0.00fF
C15816 NAND2X1_LOC_541/Y INVX1_LOC_16/A 0.01fF
C15817 INVX1_LOC_90/A NAND2X1_LOC_686/a_36_24# 0.00fF
C15818 INVX1_LOC_36/A INVX1_LOC_6/A 2.59fF
C15819 INVX1_LOC_135/A NAND2X1_LOC_562/B 0.10fF
C15820 INVX1_LOC_5/A INVX1_LOC_280/A 1.18fF
C15821 INVX1_LOC_9/Y NOR2X1_LOC_136/Y 0.05fF
C15822 NAND2X1_LOC_35/B NOR2X1_LOC_32/Y 0.06fF
C15823 INVX1_LOC_5/A NOR2X1_LOC_94/Y 0.15fF
C15824 NOR2X1_LOC_542/Y NOR2X1_LOC_542/a_36_216# -0.00fF
C15825 NAND2X1_LOC_706/Y VDD 0.08fF
C15826 NOR2X1_LOC_245/a_36_216# NAND2X1_LOC_357/B 0.00fF
C15827 INVX1_LOC_27/A NAND2X1_LOC_96/A 0.07fF
C15828 INVX1_LOC_34/A INPUT_1 0.15fF
C15829 NOR2X1_LOC_15/Y INVX1_LOC_14/Y 0.10fF
C15830 NAND2X1_LOC_364/A INVX1_LOC_285/Y 0.03fF
C15831 NOR2X1_LOC_267/A INVX1_LOC_6/A 0.08fF
C15832 INVX1_LOC_14/A NAND2X1_LOC_287/B 0.07fF
C15833 INVX1_LOC_49/A INVX1_LOC_131/A 0.08fF
C15834 NAND2X1_LOC_470/B NAND2X1_LOC_74/B 0.12fF
C15835 NOR2X1_LOC_82/A INVX1_LOC_76/A 0.08fF
C15836 NOR2X1_LOC_91/A INVX1_LOC_63/A 4.75fF
C15837 INVX1_LOC_178/A INVX1_LOC_280/A 0.05fF
C15838 INVX1_LOC_52/Y INVX1_LOC_281/A 0.01fF
C15839 NOR2X1_LOC_158/Y INVX1_LOC_29/A 0.08fF
C15840 NOR2X1_LOC_798/A NOR2X1_LOC_729/A 0.00fF
C15841 NAND2X1_LOC_550/A NAND2X1_LOC_244/A 0.07fF
C15842 INVX1_LOC_14/A INVX1_LOC_129/Y 0.00fF
C15843 NOR2X1_LOC_553/Y NOR2X1_LOC_569/Y 0.01fF
C15844 INVX1_LOC_89/A INVX1_LOC_189/A 0.00fF
C15845 NOR2X1_LOC_309/Y NAND2X1_LOC_807/Y 0.87fF
C15846 INVX1_LOC_49/A INPUT_0 0.10fF
C15847 NOR2X1_LOC_208/Y INVX1_LOC_6/A 0.10fF
C15848 INVX1_LOC_135/A NOR2X1_LOC_773/Y 0.10fF
C15849 INVX1_LOC_24/A INVX1_LOC_123/A 0.01fF
C15850 NOR2X1_LOC_593/Y NOR2X1_LOC_534/a_36_216# 0.03fF
C15851 INVX1_LOC_129/A NOR2X1_LOC_814/A 0.07fF
C15852 INVX1_LOC_23/A INVX1_LOC_63/A 0.22fF
C15853 NOR2X1_LOC_237/Y INVX1_LOC_6/A 0.09fF
C15854 INVX1_LOC_33/A INVX1_LOC_86/A 0.02fF
C15855 NAND2X1_LOC_364/A INVX1_LOC_65/A 0.03fF
C15856 NOR2X1_LOC_660/Y NOR2X1_LOC_649/B 1.84fF
C15857 NOR2X1_LOC_802/A NOR2X1_LOC_567/B 0.08fF
C15858 INVX1_LOC_41/A INVX1_LOC_311/A 0.21fF
C15859 NOR2X1_LOC_660/Y INVX1_LOC_3/A 0.03fF
C15860 NAND2X1_LOC_36/A INVX1_LOC_76/A 0.00fF
C15861 INVX1_LOC_83/A INVX1_LOC_32/Y 0.02fF
C15862 D_INPUT_1 NAND2X1_LOC_773/B 0.55fF
C15863 NAND2X1_LOC_198/B NAND2X1_LOC_642/Y 0.01fF
C15864 NOR2X1_LOC_714/a_36_216# NOR2X1_LOC_374/A 0.00fF
C15865 NOR2X1_LOC_516/B INVX1_LOC_89/A 0.09fF
C15866 NOR2X1_LOC_816/A NOR2X1_LOC_152/A 0.01fF
C15867 NOR2X1_LOC_52/Y NAND2X1_LOC_469/B 0.03fF
C15868 NOR2X1_LOC_576/B NAND2X1_LOC_735/B 0.10fF
C15869 NOR2X1_LOC_726/Y VDD 0.04fF
C15870 INVX1_LOC_150/Y NOR2X1_LOC_114/a_36_216# 0.00fF
C15871 INVX1_LOC_104/A INVX1_LOC_222/A 0.72fF
C15872 NOR2X1_LOC_274/Y INVX1_LOC_93/Y 0.09fF
C15873 INVX1_LOC_72/A NAND2X1_LOC_39/Y 0.03fF
C15874 NOR2X1_LOC_309/Y INVX1_LOC_6/A 0.02fF
C15875 NOR2X1_LOC_516/B NAND2X1_LOC_508/A 0.07fF
C15876 NAND2X1_LOC_514/Y INVX1_LOC_76/A 0.01fF
C15877 INVX1_LOC_21/A NAND2X1_LOC_574/A -0.02fF
C15878 INVX1_LOC_2/A INPUT_0 0.10fF
C15879 INVX1_LOC_101/Y INVX1_LOC_92/A 0.02fF
C15880 NOR2X1_LOC_168/B NOR2X1_LOC_337/A 0.00fF
C15881 INVX1_LOC_135/A NOR2X1_LOC_332/A 0.12fF
C15882 NOR2X1_LOC_45/B INVX1_LOC_63/Y 0.03fF
C15883 NOR2X1_LOC_360/Y INVX1_LOC_2/Y 0.03fF
C15884 INVX1_LOC_77/A NOR2X1_LOC_542/B 0.01fF
C15885 NOR2X1_LOC_90/a_36_216# NOR2X1_LOC_813/Y 0.01fF
C15886 NAND2X1_LOC_837/Y NOR2X1_LOC_670/Y 0.17fF
C15887 NAND2X1_LOC_563/A INVX1_LOC_75/A 0.07fF
C15888 NOR2X1_LOC_493/A INVX1_LOC_42/A 0.01fF
C15889 NOR2X1_LOC_596/A NOR2X1_LOC_603/Y 0.01fF
C15890 INVX1_LOC_88/A INVX1_LOC_307/A 0.07fF
C15891 INVX1_LOC_292/A INVX1_LOC_9/A 1.08fF
C15892 INVX1_LOC_49/A NOR2X1_LOC_324/A 0.04fF
C15893 NOR2X1_LOC_91/Y INVX1_LOC_37/A 0.03fF
C15894 NOR2X1_LOC_584/a_36_216# INVX1_LOC_77/Y 0.01fF
C15895 INVX1_LOC_215/Y INVX1_LOC_54/A 0.04fF
C15896 NOR2X1_LOC_226/A INPUT_0 0.22fF
C15897 INVX1_LOC_58/A NOR2X1_LOC_48/B 0.23fF
C15898 INVX1_LOC_181/Y INVX1_LOC_46/A 0.07fF
C15899 INVX1_LOC_3/Y NAND2X1_LOC_215/A 0.23fF
C15900 INVX1_LOC_31/A NOR2X1_LOC_656/Y 0.05fF
C15901 NAND2X1_LOC_276/Y INVX1_LOC_95/Y 0.15fF
C15902 NAND2X1_LOC_208/B INVX1_LOC_118/A 0.02fF
C15903 NOR2X1_LOC_772/B INVX1_LOC_12/A 0.07fF
C15904 NOR2X1_LOC_360/Y NOR2X1_LOC_363/Y 0.23fF
C15905 INVX1_LOC_136/A NOR2X1_LOC_536/A 1.94fF
C15906 INVX1_LOC_35/A NAND2X1_LOC_254/Y 0.03fF
C15907 INVX1_LOC_77/A NOR2X1_LOC_137/Y 0.06fF
C15908 NAND2X1_LOC_53/Y INVX1_LOC_107/Y 0.00fF
C15909 INVX1_LOC_254/Y VDD 0.62fF
C15910 INVX1_LOC_13/Y INVX1_LOC_12/A 0.07fF
C15911 NOR2X1_LOC_598/B INVX1_LOC_32/A 0.08fF
C15912 INVX1_LOC_78/A NOR2X1_LOC_106/a_36_216# 0.00fF
C15913 NAND2X1_LOC_477/A INVX1_LOC_304/A 0.10fF
C15914 INVX1_LOC_177/A NOR2X1_LOC_405/A 0.00fF
C15915 INVX1_LOC_135/A INVX1_LOC_140/A 0.10fF
C15916 NAND2X1_LOC_332/Y INVX1_LOC_76/A 0.01fF
C15917 NOR2X1_LOC_598/B NOR2X1_LOC_623/B 0.00fF
C15918 NAND2X1_LOC_169/Y INVX1_LOC_102/A 0.02fF
C15919 NAND2X1_LOC_286/B NOR2X1_LOC_301/A 0.04fF
C15920 INVX1_LOC_45/A INVX1_LOC_291/A 0.07fF
C15921 INVX1_LOC_57/A NAND2X1_LOC_223/A 0.07fF
C15922 NOR2X1_LOC_445/Y VDD 0.12fF
C15923 NOR2X1_LOC_19/B NAND2X1_LOC_624/A 0.00fF
C15924 INVX1_LOC_214/Y NAND2X1_LOC_655/A 0.01fF
C15925 NOR2X1_LOC_689/Y NAND2X1_LOC_175/Y 0.08fF
C15926 NAND2X1_LOC_182/A INVX1_LOC_20/A 0.12fF
C15927 INVX1_LOC_13/A INVX1_LOC_201/A 0.00fF
C15928 INVX1_LOC_135/A NAND2X1_LOC_463/B 0.00fF
C15929 INVX1_LOC_96/Y NAND2X1_LOC_212/Y 0.00fF
C15930 INVX1_LOC_286/Y NOR2X1_LOC_88/Y 0.07fF
C15931 INVX1_LOC_89/A NOR2X1_LOC_706/A 0.01fF
C15932 NAND2X1_LOC_601/a_36_24# INVX1_LOC_33/Y 0.00fF
C15933 INVX1_LOC_17/A NOR2X1_LOC_721/B 0.02fF
C15934 NOR2X1_LOC_860/B INVX1_LOC_230/A 0.59fF
C15935 INVX1_LOC_136/A NAND2X1_LOC_93/B 0.08fF
C15936 NAND2X1_LOC_715/B INVX1_LOC_32/A 0.24fF
C15937 NOR2X1_LOC_214/B INVX1_LOC_75/A 0.06fF
C15938 NAND2X1_LOC_341/A INVX1_LOC_159/Y 0.01fF
C15939 NOR2X1_LOC_91/Y NOR2X1_LOC_177/Y 0.35fF
C15940 NOR2X1_LOC_523/B NOR2X1_LOC_61/Y 0.03fF
C15941 NOR2X1_LOC_369/Y INVX1_LOC_84/A 0.01fF
C15942 NOR2X1_LOC_152/Y NOR2X1_LOC_331/B 0.10fF
C15943 NOR2X1_LOC_78/A INVX1_LOC_16/A 0.03fF
C15944 NOR2X1_LOC_500/B NOR2X1_LOC_445/B 0.01fF
C15945 NOR2X1_LOC_391/B NOR2X1_LOC_332/A 0.08fF
C15946 INVX1_LOC_25/A INVX1_LOC_23/Y 0.03fF
C15947 INVX1_LOC_38/Y INVX1_LOC_15/A 0.04fF
C15948 NOR2X1_LOC_797/a_36_216# INVX1_LOC_75/A 0.02fF
C15949 NAND2X1_LOC_141/A D_INPUT_3 0.08fF
C15950 INVX1_LOC_63/Y INVX1_LOC_281/A 0.03fF
C15951 INVX1_LOC_272/Y INVX1_LOC_272/A 0.12fF
C15952 INVX1_LOC_53/Y NAND2X1_LOC_642/Y 0.07fF
C15953 INVX1_LOC_88/A INVX1_LOC_12/A 0.01fF
C15954 NOR2X1_LOC_372/A NAND2X1_LOC_489/Y 0.14fF
C15955 INVX1_LOC_96/Y INVX1_LOC_14/Y 0.10fF
C15956 INVX1_LOC_187/A INVX1_LOC_22/A 0.01fF
C15957 INPUT_0 INPUT_1 0.41fF
C15958 INVX1_LOC_286/Y INVX1_LOC_84/A 0.07fF
C15959 INVX1_LOC_267/Y D_GATE_662 0.24fF
C15960 INVX1_LOC_23/A NOR2X1_LOC_65/Y 0.00fF
C15961 INVX1_LOC_31/A INVX1_LOC_63/A 1.17fF
C15962 INVX1_LOC_279/A INVX1_LOC_91/A 0.07fF
C15963 NOR2X1_LOC_168/Y NOR2X1_LOC_197/B 0.01fF
C15964 INVX1_LOC_67/A INVX1_LOC_9/A 0.02fF
C15965 NAND2X1_LOC_725/A NAND2X1_LOC_175/Y 0.10fF
C15966 INVX1_LOC_256/A NAND2X1_LOC_74/B 0.07fF
C15967 NAND2X1_LOC_463/B INVX1_LOC_169/Y 0.01fF
C15968 NAND2X1_LOC_586/a_36_24# NAND2X1_LOC_798/B 0.00fF
C15969 NAND2X1_LOC_650/B NAND2X1_LOC_850/Y 0.83fF
C15970 NOR2X1_LOC_606/Y INVX1_LOC_293/Y 0.14fF
C15971 D_INPUT_0 INVX1_LOC_125/Y 0.07fF
C15972 NOR2X1_LOC_719/A INVX1_LOC_59/Y 0.00fF
C15973 NOR2X1_LOC_405/A NAND2X1_LOC_573/A 0.01fF
C15974 INVX1_LOC_136/A INVX1_LOC_3/A 0.10fF
C15975 NAND2X1_LOC_562/B INVX1_LOC_280/A 0.10fF
C15976 INVX1_LOC_34/A INVX1_LOC_118/A 0.03fF
C15977 NAND2X1_LOC_363/B NOR2X1_LOC_39/Y 0.07fF
C15978 INVX1_LOC_300/Y INVX1_LOC_297/A 1.97fF
C15979 INVX1_LOC_89/A INVX1_LOC_315/Y 0.03fF
C15980 NOR2X1_LOC_68/A NOR2X1_LOC_673/A 0.12fF
C15981 NOR2X1_LOC_655/B INVX1_LOC_117/A 0.03fF
C15982 NOR2X1_LOC_147/B INVX1_LOC_274/A 0.10fF
C15983 NOR2X1_LOC_629/B NOR2X1_LOC_629/Y 0.03fF
C15984 NOR2X1_LOC_773/Y NOR2X1_LOC_558/a_36_216# 0.01fF
C15985 NAND2X1_LOC_555/Y NOR2X1_LOC_610/Y 0.03fF
C15986 NOR2X1_LOC_82/A INVX1_LOC_127/Y 0.03fF
C15987 D_GATE_579 VDD 0.06fF
C15988 NOR2X1_LOC_224/Y NOR2X1_LOC_696/Y 0.25fF
C15989 INVX1_LOC_25/Y INVX1_LOC_12/Y 1.15fF
C15990 NOR2X1_LOC_636/B NOR2X1_LOC_467/A 0.07fF
C15991 NOR2X1_LOC_309/Y NOR2X1_LOC_79/A 0.02fF
C15992 VDD NOR2X1_LOC_32/Y 0.23fF
C15993 INVX1_LOC_28/A NOR2X1_LOC_78/A 0.07fF
C15994 INVX1_LOC_27/A NAND2X1_LOC_99/A 1.37fF
C15995 NAND2X1_LOC_231/Y INVX1_LOC_118/A 0.10fF
C15996 INVX1_LOC_83/A INVX1_LOC_115/A 0.01fF
C15997 INVX1_LOC_306/A INVX1_LOC_76/A 0.01fF
C15998 INVX1_LOC_163/A INVX1_LOC_175/A 0.13fF
C15999 NAND2X1_LOC_390/A NOR2X1_LOC_176/Y 0.08fF
C16000 NOR2X1_LOC_168/B NOR2X1_LOC_640/Y 0.47fF
C16001 NOR2X1_LOC_403/B NAND2X1_LOC_773/B 0.40fF
C16002 NAND2X1_LOC_849/a_36_24# NOR2X1_LOC_536/A 0.00fF
C16003 NOR2X1_LOC_315/Y NOR2X1_LOC_216/B 0.11fF
C16004 NOR2X1_LOC_739/Y INVX1_LOC_271/Y 0.12fF
C16005 INVX1_LOC_1/A INVX1_LOC_23/Y 0.10fF
C16006 INVX1_LOC_207/A NOR2X1_LOC_485/Y 0.03fF
C16007 INVX1_LOC_108/Y INVX1_LOC_38/Y 0.02fF
C16008 NOR2X1_LOC_542/Y VDD 0.16fF
C16009 INVX1_LOC_308/Y NOR2X1_LOC_318/A 0.01fF
C16010 NOR2X1_LOC_283/a_36_216# NAND2X1_LOC_63/Y 0.00fF
C16011 NOR2X1_LOC_67/A NAND2X1_LOC_243/B 0.01fF
C16012 NAND2X1_LOC_798/A NOR2X1_LOC_510/B 0.05fF
C16013 NOR2X1_LOC_759/Y NOR2X1_LOC_89/A 0.00fF
C16014 INVX1_LOC_28/A NAND2X1_LOC_464/A 0.01fF
C16015 NAND2X1_LOC_842/B NOR2X1_LOC_558/A 0.00fF
C16016 NOR2X1_LOC_597/A VDD 0.00fF
C16017 INVX1_LOC_226/Y NOR2X1_LOC_99/Y 0.05fF
C16018 INVX1_LOC_202/A NOR2X1_LOC_89/A 0.25fF
C16019 INVX1_LOC_311/Y VDD 0.31fF
C16020 NOR2X1_LOC_315/Y NAND2X1_LOC_477/Y 0.01fF
C16021 NOR2X1_LOC_332/A INVX1_LOC_280/A 0.04fF
C16022 INVX1_LOC_285/Y NOR2X1_LOC_405/A 0.01fF
C16023 INVX1_LOC_21/A NAND2X1_LOC_35/Y 0.07fF
C16024 INVX1_LOC_159/A INVX1_LOC_15/A 0.03fF
C16025 NOR2X1_LOC_87/a_36_216# NAND2X1_LOC_206/Y 0.01fF
C16026 D_INPUT_4 NOR2X1_LOC_31/a_36_216# 0.00fF
C16027 INVX1_LOC_36/A NOR2X1_LOC_80/Y 0.06fF
C16028 NOR2X1_LOC_826/Y NOR2X1_LOC_15/Y 0.01fF
C16029 INVX1_LOC_101/Y INVX1_LOC_53/A 0.01fF
C16030 INVX1_LOC_297/Y INVX1_LOC_297/A 0.01fF
C16031 NOR2X1_LOC_443/a_36_216# NOR2X1_LOC_443/Y 0.02fF
C16032 NAND2X1_LOC_364/A INVX1_LOC_4/Y 0.17fF
C16033 INVX1_LOC_120/A INVX1_LOC_9/A 0.03fF
C16034 INVX1_LOC_28/A NOR2X1_LOC_60/Y 0.11fF
C16035 NOR2X1_LOC_264/Y INVX1_LOC_106/Y 0.03fF
C16036 INVX1_LOC_17/A NAND2X1_LOC_860/A 0.11fF
C16037 NOR2X1_LOC_456/Y INVX1_LOC_11/A 0.07fF
C16038 NAND2X1_LOC_218/a_36_24# NAND2X1_LOC_555/Y 0.00fF
C16039 NOR2X1_LOC_388/Y INVX1_LOC_42/A 0.07fF
C16040 INVX1_LOC_75/A INVX1_LOC_12/Y 0.27fF
C16041 NOR2X1_LOC_335/B VDD 0.40fF
C16042 NOR2X1_LOC_760/a_36_216# INVX1_LOC_53/A 0.01fF
C16043 INVX1_LOC_30/A NOR2X1_LOC_39/Y 0.07fF
C16044 NOR2X1_LOC_384/Y INVX1_LOC_23/Y 0.09fF
C16045 INVX1_LOC_58/A NOR2X1_LOC_441/Y 0.40fF
C16046 NAND2X1_LOC_25/a_36_24# NAND2X1_LOC_30/Y 0.00fF
C16047 INVX1_LOC_36/A INVX1_LOC_270/A 0.03fF
C16048 NOR2X1_LOC_160/B NOR2X1_LOC_392/Y 0.07fF
C16049 NOR2X1_LOC_178/Y NOR2X1_LOC_82/A 0.08fF
C16050 NOR2X1_LOC_78/A NOR2X1_LOC_35/Y 0.01fF
C16051 NAND2X1_LOC_391/Y NOR2X1_LOC_468/Y 0.02fF
C16052 NOR2X1_LOC_615/Y NAND2X1_LOC_624/B 0.07fF
C16053 INVX1_LOC_258/Y NOR2X1_LOC_92/Y -0.01fF
C16054 NOR2X1_LOC_274/Y INVX1_LOC_87/A -0.00fF
C16055 NOR2X1_LOC_67/A INVX1_LOC_284/A 0.51fF
C16056 INVX1_LOC_62/A NOR2X1_LOC_243/B 0.37fF
C16057 NOR2X1_LOC_798/A NOR2X1_LOC_286/Y 0.03fF
C16058 VDD INVX1_LOC_264/Y 0.26fF
C16059 NOR2X1_LOC_152/Y NOR2X1_LOC_449/A 0.06fF
C16060 INVX1_LOC_65/A NOR2X1_LOC_857/A 0.07fF
C16061 INVX1_LOC_104/A INVX1_LOC_4/A 0.07fF
C16062 NAND2X1_LOC_660/Y INVX1_LOC_19/A 0.03fF
C16063 NAND2X1_LOC_800/A INVX1_LOC_264/Y 0.01fF
C16064 D_INPUT_0 NOR2X1_LOC_653/Y 0.05fF
C16065 INVX1_LOC_203/Y INVX1_LOC_175/A 0.01fF
C16066 NOR2X1_LOC_790/B INVX1_LOC_223/A 0.00fF
C16067 NAND2X1_LOC_107/a_36_24# INVX1_LOC_46/A 0.00fF
C16068 INPUT_0 INVX1_LOC_118/A 0.22fF
C16069 NOR2X1_LOC_15/Y NAND2X1_LOC_303/Y 0.07fF
C16070 NOR2X1_LOC_388/Y INVX1_LOC_78/A 0.03fF
C16071 NOR2X1_LOC_360/Y INVX1_LOC_29/Y 0.46fF
C16072 INVX1_LOC_13/A INVX1_LOC_29/A 0.34fF
C16073 INVX1_LOC_17/A NAND2X1_LOC_473/A 1.04fF
C16074 NAND2X1_LOC_112/Y INVX1_LOC_109/A 0.00fF
C16075 INVX1_LOC_11/A NAND2X1_LOC_714/B 0.00fF
C16076 INVX1_LOC_59/Y INVX1_LOC_76/A 0.01fF
C16077 NOR2X1_LOC_208/Y INVX1_LOC_270/A 0.07fF
C16078 NOR2X1_LOC_363/Y NOR2X1_LOC_269/Y 0.00fF
C16079 INVX1_LOC_194/A INVX1_LOC_253/A 0.05fF
C16080 NOR2X1_LOC_590/A NOR2X1_LOC_849/A 0.69fF
C16081 NAND2X1_LOC_738/B NAND2X1_LOC_731/Y 0.00fF
C16082 INVX1_LOC_36/A NOR2X1_LOC_109/Y 0.07fF
C16083 D_INPUT_1 INVX1_LOC_24/A 0.22fF
C16084 INVX1_LOC_10/A INVX1_LOC_272/A 0.03fF
C16085 NAND2X1_LOC_434/a_36_24# NAND2X1_LOC_453/A 0.00fF
C16086 NAND2X1_LOC_308/Y NAND2X1_LOC_175/Y 0.03fF
C16087 D_INPUT_0 INVX1_LOC_19/A 0.25fF
C16088 NOR2X1_LOC_583/a_36_216# NOR2X1_LOC_584/Y 0.00fF
C16089 INVX1_LOC_17/A NAND2X1_LOC_537/Y 0.11fF
C16090 NOR2X1_LOC_387/Y INVX1_LOC_296/Y 0.10fF
C16091 INVX1_LOC_39/A NAND2X1_LOC_208/B 0.02fF
C16092 VDD NOR2X1_LOC_825/Y 0.28fF
C16093 NAND2X1_LOC_807/Y NOR2X1_LOC_654/a_36_216# 0.01fF
C16094 NOR2X1_LOC_815/A NAND2X1_LOC_798/B 0.02fF
C16095 NOR2X1_LOC_665/A NAND2X1_LOC_792/B 0.09fF
C16096 NAND2X1_LOC_563/a_36_24# INVX1_LOC_1/A -0.02fF
C16097 INVX1_LOC_278/A NOR2X1_LOC_191/B 0.02fF
C16098 NAND2X1_LOC_254/a_36_24# INVX1_LOC_46/A 0.00fF
C16099 NAND2X1_LOC_807/Y INVX1_LOC_63/A 0.03fF
C16100 NAND2X1_LOC_53/Y NOR2X1_LOC_740/Y 0.25fF
C16101 INVX1_LOC_33/A INVX1_LOC_57/A 0.14fF
C16102 NOR2X1_LOC_246/A INVX1_LOC_29/A 0.07fF
C16103 NOR2X1_LOC_352/Y INVX1_LOC_271/Y 0.05fF
C16104 INPUT_1 NOR2X1_LOC_84/B -0.00fF
C16105 INVX1_LOC_47/A INVX1_LOC_125/A 0.14fF
C16106 NOR2X1_LOC_174/B INVX1_LOC_29/A 0.05fF
C16107 NAND2X1_LOC_560/A NAND2X1_LOC_489/Y 0.22fF
C16108 NAND2X1_LOC_471/a_36_24# NAND2X1_LOC_99/A 0.00fF
C16109 D_INPUT_1 NOR2X1_LOC_557/Y 0.19fF
C16110 NAND2X1_LOC_551/A INVX1_LOC_29/A 0.03fF
C16111 INVX1_LOC_135/A INVX1_LOC_42/A 0.22fF
C16112 NOR2X1_LOC_309/Y INVX1_LOC_270/A 0.01fF
C16113 NAND2X1_LOC_214/B NAND2X1_LOC_656/A 0.03fF
C16114 NAND2X1_LOC_357/B NOR2X1_LOC_280/a_36_216# 0.00fF
C16115 NOR2X1_LOC_84/Y INVX1_LOC_112/Y 0.03fF
C16116 NOR2X1_LOC_446/a_36_216# NOR2X1_LOC_457/A 0.02fF
C16117 NAND2X1_LOC_680/a_36_24# INVX1_LOC_49/Y 0.00fF
C16118 NOR2X1_LOC_186/Y NOR2X1_LOC_744/Y 0.01fF
C16119 INVX1_LOC_120/A NOR2X1_LOC_861/Y 0.03fF
C16120 INVX1_LOC_256/A NOR2X1_LOC_276/Y 0.00fF
C16121 INVX1_LOC_143/Y INVX1_LOC_9/A 0.03fF
C16122 NAND2X1_LOC_655/A INVX1_LOC_92/A 0.08fF
C16123 NOR2X1_LOC_385/a_36_216# INVX1_LOC_12/A 0.02fF
C16124 INVX1_LOC_25/Y NOR2X1_LOC_89/Y -0.00fF
C16125 INVX1_LOC_27/A NAND2X1_LOC_656/A 0.23fF
C16126 NAND2X1_LOC_479/Y INVX1_LOC_78/A 0.00fF
C16127 INVX1_LOC_21/A INVX1_LOC_94/A 0.27fF
C16128 INVX1_LOC_34/A INVX1_LOC_138/A 0.02fF
C16129 NOR2X1_LOC_285/Y INVX1_LOC_310/Y 0.01fF
C16130 NOR2X1_LOC_137/Y INVX1_LOC_9/A 0.01fF
C16131 NAND2X1_LOC_342/Y INVX1_LOC_270/Y 0.14fF
C16132 NOR2X1_LOC_598/B INVX1_LOC_158/A 0.12fF
C16133 INVX1_LOC_6/A INVX1_LOC_63/A 0.03fF
C16134 NAND2X1_LOC_573/Y NOR2X1_LOC_744/Y 0.05fF
C16135 NOR2X1_LOC_400/A INVX1_LOC_201/Y 0.03fF
C16136 INVX1_LOC_64/A INVX1_LOC_104/A 0.07fF
C16137 NOR2X1_LOC_848/Y NOR2X1_LOC_554/B 0.31fF
C16138 INVX1_LOC_190/Y INVX1_LOC_15/A 0.15fF
C16139 INPUT_0 NAND2X1_LOC_63/Y 0.12fF
C16140 INVX1_LOC_22/A NOR2X1_LOC_621/A 0.02fF
C16141 NOR2X1_LOC_683/Y INVX1_LOC_92/A 0.03fF
C16142 NOR2X1_LOC_557/Y NOR2X1_LOC_652/Y 0.54fF
C16143 NOR2X1_LOC_88/Y NOR2X1_LOC_56/Y 0.00fF
C16144 INVX1_LOC_137/A NAND2X1_LOC_99/A 0.03fF
C16145 NAND2X1_LOC_714/B NOR2X1_LOC_433/A 0.03fF
C16146 INVX1_LOC_40/A INVX1_LOC_57/A 0.20fF
C16147 INVX1_LOC_256/A INVX1_LOC_136/A 0.13fF
C16148 INVX1_LOC_233/A NAND2X1_LOC_775/a_36_24# 0.00fF
C16149 INVX1_LOC_233/Y NAND2X1_LOC_785/A 0.09fF
C16150 NOR2X1_LOC_10/a_36_216# INVX1_LOC_63/A 0.00fF
C16151 NOR2X1_LOC_75/Y NAND2X1_LOC_16/Y 0.01fF
C16152 INVX1_LOC_292/A NOR2X1_LOC_565/A 0.01fF
C16153 NOR2X1_LOC_83/a_36_216# INVX1_LOC_12/A 0.00fF
C16154 INVX1_LOC_135/A INVX1_LOC_78/A 0.13fF
C16155 NOR2X1_LOC_667/a_36_216# INVX1_LOC_36/A 0.00fF
C16156 NAND2X1_LOC_778/Y NOR2X1_LOC_690/A 0.02fF
C16157 NOR2X1_LOC_392/B INVX1_LOC_306/Y 0.39fF
C16158 INVX1_LOC_39/A INVX1_LOC_34/A 0.04fF
C16159 INVX1_LOC_69/Y NAND2X1_LOC_74/B 0.08fF
C16160 INVX1_LOC_299/A NOR2X1_LOC_303/Y 0.10fF
C16161 NOR2X1_LOC_262/a_36_216# INVX1_LOC_1/Y 0.00fF
C16162 NOR2X1_LOC_544/A INVX1_LOC_53/A 0.05fF
C16163 INPUT_0 NAND2X1_LOC_455/B 0.01fF
C16164 INVX1_LOC_35/A NOR2X1_LOC_778/B 0.03fF
C16165 INVX1_LOC_25/A INVX1_LOC_232/A 0.14fF
C16166 INVX1_LOC_75/A NOR2X1_LOC_554/A 0.07fF
C16167 NOR2X1_LOC_391/B NOR2X1_LOC_847/A 0.10fF
C16168 NOR2X1_LOC_859/A NOR2X1_LOC_590/A 0.01fF
C16169 INVX1_LOC_1/Y INVX1_LOC_23/A 0.01fF
C16170 NOR2X1_LOC_56/Y INVX1_LOC_84/A 0.03fF
C16171 INVX1_LOC_21/A NOR2X1_LOC_234/Y 0.05fF
C16172 VDD NOR2X1_LOC_88/Y 0.80fF
C16173 INVX1_LOC_269/A NOR2X1_LOC_577/Y 0.00fF
C16174 D_INPUT_0 INVX1_LOC_26/Y 0.06fF
C16175 NOR2X1_LOC_246/A NOR2X1_LOC_281/Y 0.01fF
C16176 NAND2X1_LOC_659/B INVX1_LOC_84/A 0.07fF
C16177 INVX1_LOC_48/Y NAND2X1_LOC_139/A 0.01fF
C16178 NOR2X1_LOC_666/Y INVX1_LOC_33/A 0.12fF
C16179 INVX1_LOC_25/A NOR2X1_LOC_383/Y 0.72fF
C16180 NOR2X1_LOC_690/A NOR2X1_LOC_15/Y 0.06fF
C16181 INVX1_LOC_27/A NOR2X1_LOC_423/Y 0.02fF
C16182 INVX1_LOC_274/A INVX1_LOC_38/A 0.00fF
C16183 INVX1_LOC_64/A INVX1_LOC_263/A 0.16fF
C16184 NAND2X1_LOC_803/B NAND2X1_LOC_593/Y 0.04fF
C16185 INVX1_LOC_11/A NOR2X1_LOC_550/B 0.01fF
C16186 NOR2X1_LOC_78/A INVX1_LOC_109/A 0.00fF
C16187 NOR2X1_LOC_441/Y NOR2X1_LOC_338/Y -0.00fF
C16188 INVX1_LOC_298/Y INVX1_LOC_55/Y 0.91fF
C16189 NOR2X1_LOC_598/B GATE_662 0.02fF
C16190 INPUT_1 INVX1_LOC_183/A 0.02fF
C16191 NOR2X1_LOC_716/B NAND2X1_LOC_793/Y 0.02fF
C16192 VDD INVX1_LOC_84/A 1.43fF
C16193 INVX1_LOC_13/Y NOR2X1_LOC_566/Y 0.04fF
C16194 INVX1_LOC_14/A NOR2X1_LOC_6/B 2.70fF
C16195 NOR2X1_LOC_71/Y NAND2X1_LOC_458/a_36_24# 0.00fF
C16196 NAND2X1_LOC_729/Y NAND2X1_LOC_741/B 0.03fF
C16197 NAND2X1_LOC_800/A INVX1_LOC_84/A 0.03fF
C16198 NOR2X1_LOC_590/A NAND2X1_LOC_593/Y 0.07fF
C16199 NOR2X1_LOC_457/A NOR2X1_LOC_570/B 0.12fF
C16200 D_INPUT_1 NOR2X1_LOC_130/A 0.09fF
C16201 INVX1_LOC_233/Y NAND2X1_LOC_632/a_36_24# 0.01fF
C16202 INVX1_LOC_27/A NOR2X1_LOC_222/Y 0.07fF
C16203 INVX1_LOC_21/A NOR2X1_LOC_136/Y 0.01fF
C16204 INVX1_LOC_206/Y INVX1_LOC_4/A 0.03fF
C16205 INVX1_LOC_11/A INVX1_LOC_249/Y 0.01fF
C16206 NOR2X1_LOC_337/Y INVX1_LOC_15/A 0.01fF
C16207 NOR2X1_LOC_186/Y INVX1_LOC_16/A 0.05fF
C16208 INVX1_LOC_299/A INVX1_LOC_54/Y 0.19fF
C16209 INVX1_LOC_223/Y NOR2X1_LOC_516/B 0.06fF
C16210 INVX1_LOC_304/A INVX1_LOC_168/Y 0.01fF
C16211 NAND2X1_LOC_541/Y INVX1_LOC_48/Y 0.02fF
C16212 NOR2X1_LOC_763/a_36_216# INVX1_LOC_30/A 0.01fF
C16213 VDD NAND2X1_LOC_651/B 0.01fF
C16214 NOR2X1_LOC_160/B INVX1_LOC_176/Y 0.03fF
C16215 NOR2X1_LOC_590/A NOR2X1_LOC_758/Y 0.01fF
C16216 NAND2X1_LOC_848/A NOR2X1_LOC_653/Y 0.07fF
C16217 NOR2X1_LOC_329/B INVX1_LOC_271/A 0.19fF
C16218 NAND2X1_LOC_555/Y NOR2X1_LOC_516/Y 0.14fF
C16219 NOR2X1_LOC_718/Y NOR2X1_LOC_717/Y 0.03fF
C16220 NOR2X1_LOC_567/B NOR2X1_LOC_809/A 0.05fF
C16221 INVX1_LOC_214/Y INVX1_LOC_88/A 0.24fF
C16222 INVX1_LOC_91/A NOR2X1_LOC_38/B 0.16fF
C16223 NAND2X1_LOC_53/Y NAND2X1_LOC_301/a_36_24# 0.00fF
C16224 NOR2X1_LOC_793/Y NAND2X1_LOC_323/B -0.01fF
C16225 INVX1_LOC_35/A NOR2X1_LOC_724/Y 5.12fF
C16226 INVX1_LOC_223/A NOR2X1_LOC_344/A 0.02fF
C16227 NAND2X1_LOC_798/B NAND2X1_LOC_436/a_36_24# 0.00fF
C16228 INVX1_LOC_200/Y NOR2X1_LOC_322/Y 0.38fF
C16229 NOR2X1_LOC_403/B INVX1_LOC_24/A 0.25fF
C16230 INVX1_LOC_103/A NOR2X1_LOC_131/a_36_216# 0.00fF
C16231 INVX1_LOC_1/A INVX1_LOC_232/A 0.12fF
C16232 NOR2X1_LOC_742/A INVX1_LOC_23/A 1.49fF
C16233 NAND2X1_LOC_44/a_36_24# INVX1_LOC_33/A 0.02fF
C16234 NOR2X1_LOC_78/B NAND2X1_LOC_183/a_36_24# 0.00fF
C16235 GATE_741 INVX1_LOC_229/Y 1.78fF
C16236 NOR2X1_LOC_323/Y INVX1_LOC_57/A 0.26fF
C16237 NAND2X1_LOC_182/A NAND2X1_LOC_860/a_36_24# 0.00fF
C16238 NOR2X1_LOC_97/A NOR2X1_LOC_383/B 0.00fF
C16239 NAND2X1_LOC_724/A INVX1_LOC_16/A 0.07fF
C16240 NOR2X1_LOC_56/Y INVX1_LOC_15/A 0.17fF
C16241 INVX1_LOC_269/A NOR2X1_LOC_325/A 0.21fF
C16242 INVX1_LOC_185/A INVX1_LOC_285/A 0.39fF
C16243 NOR2X1_LOC_92/Y NOR2X1_LOC_589/A 0.07fF
C16244 NOR2X1_LOC_243/a_36_216# INVX1_LOC_89/A 0.00fF
C16245 NAND2X1_LOC_475/Y INVX1_LOC_54/A 0.10fF
C16246 NAND2X1_LOC_659/B INVX1_LOC_15/A 0.01fF
C16247 NOR2X1_LOC_114/Y INVX1_LOC_46/A 0.01fF
C16248 INVX1_LOC_185/A INVX1_LOC_265/Y 0.02fF
C16249 INVX1_LOC_269/A INVX1_LOC_22/A 0.13fF
C16250 NOR2X1_LOC_405/A INVX1_LOC_4/Y 0.08fF
C16251 D_INPUT_3 NOR2X1_LOC_128/a_36_216# 0.00fF
C16252 NOR2X1_LOC_52/Y INVX1_LOC_63/Y 0.02fF
C16253 VDD NAND2X1_LOC_220/B 0.01fF
C16254 NOR2X1_LOC_273/Y NOR2X1_LOC_433/A 0.01fF
C16255 NAND2X1_LOC_131/a_36_24# INVX1_LOC_232/A 0.00fF
C16256 INVX1_LOC_86/A INVX1_LOC_275/Y 0.02fF
C16257 INVX1_LOC_36/A NOR2X1_LOC_309/Y 0.11fF
C16258 NAND2X1_LOC_99/Y NAND2X1_LOC_656/A 0.01fF
C16259 NOR2X1_LOC_433/A NOR2X1_LOC_759/Y 0.03fF
C16260 NOR2X1_LOC_199/B NAND2X1_LOC_473/A 0.11fF
C16261 INVX1_LOC_30/Y INVX1_LOC_14/A 0.19fF
C16262 NOR2X1_LOC_552/A INVX1_LOC_78/A 0.07fF
C16263 NOR2X1_LOC_843/A NAND2X1_LOC_364/A 0.09fF
C16264 INVX1_LOC_292/A INVX1_LOC_179/Y 0.01fF
C16265 NOR2X1_LOC_361/a_36_216# INVX1_LOC_133/Y 0.00fF
C16266 NOR2X1_LOC_177/a_36_216# NOR2X1_LOC_662/A 0.00fF
C16267 INVX1_LOC_202/A NOR2X1_LOC_433/A 0.09fF
C16268 INVX1_LOC_34/A INVX1_LOC_61/A 0.07fF
C16269 NOR2X1_LOC_240/A NAND2X1_LOC_234/a_36_24# 0.02fF
C16270 NAND2X1_LOC_768/a_36_24# NAND2X1_LOC_338/B 0.00fF
C16271 NAND2X1_LOC_550/A INVX1_LOC_25/Y 0.07fF
C16272 NOR2X1_LOC_813/Y INVX1_LOC_42/A 0.08fF
C16273 NOR2X1_LOC_192/A INVX1_LOC_26/A 0.01fF
C16274 VDD INVX1_LOC_15/A 2.04fF
C16275 NOR2X1_LOC_152/A INVX1_LOC_42/A 0.01fF
C16276 INVX1_LOC_131/Y INVX1_LOC_63/A 0.28fF
C16277 INVX1_LOC_10/Y INVX1_LOC_42/A 0.00fF
C16278 NOR2X1_LOC_160/B INVX1_LOC_25/Y 0.12fF
C16279 INVX1_LOC_103/A NOR2X1_LOC_561/Y 4.37fF
C16280 NAND2X1_LOC_766/a_36_24# INVX1_LOC_49/A 0.01fF
C16281 NOR2X1_LOC_186/Y INVX1_LOC_28/A 0.01fF
C16282 INVX1_LOC_280/A INVX1_LOC_42/A 0.32fF
C16283 NOR2X1_LOC_273/Y NOR2X1_LOC_52/B 0.12fF
C16284 NOR2X1_LOC_250/a_36_216# NAND2X1_LOC_656/Y 0.01fF
C16285 NOR2X1_LOC_91/A INVX1_LOC_93/Y 0.52fF
C16286 NAND2X1_LOC_354/B NAND2X1_LOC_593/Y 0.02fF
C16287 INVX1_LOC_27/A NOR2X1_LOC_329/B 0.07fF
C16288 INVX1_LOC_19/A INVX1_LOC_46/Y 0.07fF
C16289 NAND2X1_LOC_787/A INVX1_LOC_286/A 0.03fF
C16290 INVX1_LOC_24/A NOR2X1_LOC_591/Y 0.03fF
C16291 INVX1_LOC_31/A INVX1_LOC_1/Y 0.05fF
C16292 NOR2X1_LOC_52/B NOR2X1_LOC_759/Y 0.04fF
C16293 NOR2X1_LOC_322/Y NOR2X1_LOC_406/A 0.02fF
C16294 INVX1_LOC_150/Y INVX1_LOC_10/A 0.07fF
C16295 NOR2X1_LOC_318/B INVX1_LOC_23/A 0.24fF
C16296 NOR2X1_LOC_220/A NOR2X1_LOC_703/B 0.03fF
C16297 INVX1_LOC_292/A NOR2X1_LOC_561/Y 0.01fF
C16298 INVX1_LOC_174/A INVX1_LOC_121/A 0.16fF
C16299 NOR2X1_LOC_262/a_36_216# INVX1_LOC_93/Y 0.01fF
C16300 INVX1_LOC_78/A INVX1_LOC_139/Y 0.03fF
C16301 INVX1_LOC_298/Y NOR2X1_LOC_357/Y 0.03fF
C16302 INVX1_LOC_64/A INVX1_LOC_206/Y 0.10fF
C16303 NOR2X1_LOC_202/Y NOR2X1_LOC_215/A 0.17fF
C16304 D_INPUT_0 INVX1_LOC_161/Y 0.01fF
C16305 NOR2X1_LOC_772/Y INVX1_LOC_294/Y 0.25fF
C16306 INVX1_LOC_255/Y NOR2X1_LOC_382/Y 0.05fF
C16307 INVX1_LOC_119/A NOR2X1_LOC_637/B 0.25fF
C16308 INVX1_LOC_58/A INVX1_LOC_291/Y 0.03fF
C16309 INVX1_LOC_93/Y INVX1_LOC_23/A 0.07fF
C16310 NOR2X1_LOC_139/Y INVX1_LOC_53/A 0.03fF
C16311 NAND2X1_LOC_724/A INVX1_LOC_28/A 1.09fF
C16312 NOR2X1_LOC_344/A INVX1_LOC_149/Y 0.03fF
C16313 INVX1_LOC_53/A NAND2X1_LOC_655/A 0.07fF
C16314 INVX1_LOC_21/A INVX1_LOC_144/A 0.07fF
C16315 INVX1_LOC_215/A INVX1_LOC_30/A 0.46fF
C16316 INVX1_LOC_39/A INPUT_0 0.03fF
C16317 INVX1_LOC_49/A INVX1_LOC_266/Y 0.12fF
C16318 NAND2X1_LOC_820/a_36_24# NOR2X1_LOC_554/B 0.01fF
C16319 NOR2X1_LOC_188/A NOR2X1_LOC_846/A 0.00fF
C16320 NOR2X1_LOC_68/A NOR2X1_LOC_210/B 0.08fF
C16321 INVX1_LOC_12/A INVX1_LOC_107/Y 0.01fF
C16322 INVX1_LOC_294/Y NOR2X1_LOC_392/B 0.48fF
C16323 NAND2X1_LOC_577/A INVX1_LOC_234/A 0.02fF
C16324 NOR2X1_LOC_456/Y NOR2X1_LOC_601/Y 0.03fF
C16325 NOR2X1_LOC_226/A NAND2X1_LOC_802/A 0.03fF
C16326 NOR2X1_LOC_703/B NOR2X1_LOC_548/Y 0.16fF
C16327 NOR2X1_LOC_791/Y INVX1_LOC_286/A 0.07fF
C16328 NOR2X1_LOC_488/Y INVX1_LOC_41/Y 0.00fF
C16329 INVX1_LOC_64/A NOR2X1_LOC_600/Y 0.04fF
C16330 INVX1_LOC_136/A NOR2X1_LOC_440/Y 0.12fF
C16331 NOR2X1_LOC_91/A NAND2X1_LOC_721/A 0.11fF
C16332 NAND2X1_LOC_468/B INVX1_LOC_53/A 0.06fF
C16333 NOR2X1_LOC_445/Y INVX1_LOC_177/A 0.00fF
C16334 NAND2X1_LOC_552/A NOR2X1_LOC_45/B 0.16fF
C16335 NAND2X1_LOC_357/B INVX1_LOC_162/Y 0.01fF
C16336 INVX1_LOC_5/A NOR2X1_LOC_45/B 0.04fF
C16337 INVX1_LOC_24/A NOR2X1_LOC_553/Y 0.08fF
C16338 NAND2X1_LOC_338/B NOR2X1_LOC_520/B 0.18fF
C16339 INVX1_LOC_226/Y NOR2X1_LOC_403/a_36_216# 0.00fF
C16340 INVX1_LOC_29/A NAND2X1_LOC_489/Y 0.03fF
C16341 INVX1_LOC_15/Y NOR2X1_LOC_413/Y 0.22fF
C16342 NAND2X1_LOC_139/A INVX1_LOC_216/A 0.14fF
C16343 NAND2X1_LOC_647/B NAND2X1_LOC_93/B 0.04fF
C16344 INVX1_LOC_13/A INVX1_LOC_228/A 0.03fF
C16345 NAND2X1_LOC_341/A INVX1_LOC_105/A 0.02fF
C16346 NOR2X1_LOC_359/Y NOR2X1_LOC_665/A 0.01fF
C16347 INVX1_LOC_155/A NOR2X1_LOC_524/a_36_216# 0.00fF
C16348 INVX1_LOC_21/A NOR2X1_LOC_845/A 0.19fF
C16349 INVX1_LOC_83/A NOR2X1_LOC_354/B 0.02fF
C16350 INVX1_LOC_45/A NOR2X1_LOC_246/a_36_216# 0.01fF
C16351 NAND2X1_LOC_84/Y INVX1_LOC_30/Y 0.01fF
C16352 INVX1_LOC_135/A NOR2X1_LOC_554/B 0.02fF
C16353 NOR2X1_LOC_516/B NOR2X1_LOC_554/a_36_216# 0.00fF
C16354 NOR2X1_LOC_261/Y VDD 0.28fF
C16355 INVX1_LOC_32/A NOR2X1_LOC_58/Y 0.08fF
C16356 NOR2X1_LOC_590/A NOR2X1_LOC_535/a_36_216# 0.00fF
C16357 INVX1_LOC_45/A NOR2X1_LOC_788/B 0.04fF
C16358 INVX1_LOC_178/A NOR2X1_LOC_45/B 0.10fF
C16359 NOR2X1_LOC_648/a_36_216# NOR2X1_LOC_348/B 0.00fF
C16360 INVX1_LOC_5/A INVX1_LOC_247/A 0.00fF
C16361 NOR2X1_LOC_355/A NOR2X1_LOC_360/Y 0.10fF
C16362 INVX1_LOC_108/Y VDD 0.01fF
C16363 NAND2X1_LOC_479/Y INVX1_LOC_113/Y 0.12fF
C16364 INVX1_LOC_50/A INVX1_LOC_44/A 0.11fF
C16365 NOR2X1_LOC_481/A INVX1_LOC_16/A 1.24fF
C16366 INVX1_LOC_2/A INVX1_LOC_266/Y 0.07fF
C16367 NOR2X1_LOC_160/B INVX1_LOC_75/A 0.95fF
C16368 NOR2X1_LOC_791/Y INVX1_LOC_95/A 0.14fF
C16369 INVX1_LOC_278/A VDD 2.00fF
C16370 INVX1_LOC_47/Y NAND2X1_LOC_572/B 0.01fF
C16371 NAND2X1_LOC_577/A NOR2X1_LOC_19/B 0.15fF
C16372 NAND2X1_LOC_784/A INVX1_LOC_33/Y 0.02fF
C16373 INVX1_LOC_170/A INVX1_LOC_28/A 0.00fF
C16374 NOR2X1_LOC_256/Y INVX1_LOC_61/Y 0.01fF
C16375 INVX1_LOC_12/A INVX1_LOC_272/A 0.06fF
C16376 INVX1_LOC_1/A INVX1_LOC_186/A 0.04fF
C16377 NOR2X1_LOC_389/A INVX1_LOC_79/A 0.07fF
C16378 INVX1_LOC_72/Y INPUT_1 0.02fF
C16379 NOR2X1_LOC_468/Y INVX1_LOC_91/A 0.10fF
C16380 INVX1_LOC_11/A NOR2X1_LOC_334/A 0.01fF
C16381 D_INPUT_2 NOR2X1_LOC_130/A 0.04fF
C16382 INVX1_LOC_41/A NOR2X1_LOC_589/A 0.00fF
C16383 INVX1_LOC_32/A NOR2X1_LOC_673/B 0.04fF
C16384 NAND2X1_LOC_472/Y NOR2X1_LOC_678/A 0.02fF
C16385 NOR2X1_LOC_89/A NAND2X1_LOC_74/B 0.07fF
C16386 INVX1_LOC_34/A NAND2X1_LOC_735/B 0.03fF
C16387 INVX1_LOC_225/A INVX1_LOC_16/A 0.09fF
C16388 NOR2X1_LOC_78/B INVX1_LOC_134/Y 0.01fF
C16389 INVX1_LOC_135/A NOR2X1_LOC_152/Y 0.10fF
C16390 NOR2X1_LOC_67/A NOR2X1_LOC_537/Y 0.01fF
C16391 INVX1_LOC_121/A INVX1_LOC_153/A 0.00fF
C16392 NOR2X1_LOC_172/Y NOR2X1_LOC_171/a_36_216# 0.03fF
C16393 NAND2X1_LOC_785/A NAND2X1_LOC_862/A 0.04fF
C16394 NAND2X1_LOC_347/B NOR2X1_LOC_80/a_36_216# 0.00fF
C16395 INVX1_LOC_13/A INVX1_LOC_8/A 0.46fF
C16396 NAND2X1_LOC_725/A NAND2X1_LOC_804/Y 0.27fF
C16397 GATE_741 INVX1_LOC_20/A 0.02fF
C16398 INVX1_LOC_34/A INPUT_5 1.80fF
C16399 INVX1_LOC_181/Y NAND2X1_LOC_842/B 0.86fF
C16400 NAND2X1_LOC_717/Y NAND2X1_LOC_852/Y 0.18fF
C16401 INVX1_LOC_201/Y NAND2X1_LOC_377/Y 0.01fF
C16402 INPUT_3 INVX1_LOC_201/A 0.18fF
C16403 NOR2X1_LOC_828/Y NOR2X1_LOC_499/B 0.03fF
C16404 INVX1_LOC_26/Y INVX1_LOC_46/Y 0.11fF
C16405 NOR2X1_LOC_78/B NOR2X1_LOC_544/A 0.62fF
C16406 NOR2X1_LOC_598/B NOR2X1_LOC_261/A 0.03fF
C16407 NOR2X1_LOC_92/Y INVX1_LOC_147/Y 0.01fF
C16408 NOR2X1_LOC_216/B NAND2X1_LOC_99/A 0.10fF
C16409 INVX1_LOC_152/Y INVX1_LOC_280/A 0.01fF
C16410 NAND2X1_LOC_68/a_36_24# INVX1_LOC_76/A 0.01fF
C16411 INVX1_LOC_1/A NAND2X1_LOC_447/Y 0.01fF
C16412 NOR2X1_LOC_383/B NOR2X1_LOC_809/B 0.02fF
C16413 NOR2X1_LOC_254/a_36_216# INVX1_LOC_78/Y 0.00fF
C16414 NAND2X1_LOC_734/a_36_24# NAND2X1_LOC_808/A 0.00fF
C16415 INVX1_LOC_235/Y D_GATE_662 0.07fF
C16416 NOR2X1_LOC_92/Y INVX1_LOC_20/A 2.24fF
C16417 INVX1_LOC_5/A INVX1_LOC_281/A 0.09fF
C16418 NOR2X1_LOC_816/A NOR2X1_LOC_45/B 0.04fF
C16419 NOR2X1_LOC_207/A NOR2X1_LOC_589/A 0.04fF
C16420 INVX1_LOC_41/A INVX1_LOC_171/A 0.00fF
C16421 INVX1_LOC_32/A INVX1_LOC_29/A 0.30fF
C16422 NOR2X1_LOC_745/Y NOR2X1_LOC_746/Y 0.10fF
C16423 NAND2X1_LOC_787/A INVX1_LOC_54/A 0.04fF
C16424 INVX1_LOC_45/A NOR2X1_LOC_147/A 0.06fF
C16425 NAND2X1_LOC_550/A NAND2X1_LOC_620/a_36_24# 0.01fF
C16426 NOR2X1_LOC_389/A INVX1_LOC_91/A 0.18fF
C16427 INVX1_LOC_286/A INVX1_LOC_30/A 0.61fF
C16428 NAND2X1_LOC_860/A NOR2X1_LOC_118/a_36_216# 0.00fF
C16429 NOR2X1_LOC_264/Y INVX1_LOC_89/A 0.07fF
C16430 NOR2X1_LOC_391/A INVX1_LOC_34/Y 0.07fF
C16431 NOR2X1_LOC_391/B NOR2X1_LOC_554/B 0.02fF
C16432 NOR2X1_LOC_781/a_36_216# INVX1_LOC_266/Y 0.00fF
C16433 INVX1_LOC_61/A INPUT_0 0.05fF
C16434 INVX1_LOC_136/A INVX1_LOC_69/Y 0.15fF
C16435 NAND2X1_LOC_725/B INVX1_LOC_46/A 0.19fF
C16436 NOR2X1_LOC_481/A INVX1_LOC_28/A 0.30fF
C16437 INVX1_LOC_90/A INVX1_LOC_294/Y 0.08fF
C16438 INVX1_LOC_103/A INVX1_LOC_76/A 7.06fF
C16439 NOR2X1_LOC_48/B NOR2X1_LOC_452/a_36_216# 0.00fF
C16440 NAND2X1_LOC_568/A INVX1_LOC_20/A 0.00fF
C16441 INVX1_LOC_280/Y NOR2X1_LOC_32/Y 0.03fF
C16442 NOR2X1_LOC_208/Y NOR2X1_LOC_208/A 0.09fF
C16443 NOR2X1_LOC_563/a_36_216# NOR2X1_LOC_500/Y 0.01fF
C16444 NAND2X1_LOC_477/Y NAND2X1_LOC_99/A 0.01fF
C16445 NOR2X1_LOC_529/Y NOR2X1_LOC_130/A -0.09fF
C16446 NOR2X1_LOC_389/B INVX1_LOC_294/Y 0.02fF
C16447 INVX1_LOC_49/A INVX1_LOC_42/Y 0.02fF
C16448 NOR2X1_LOC_226/A NAND2X1_LOC_862/a_36_24# 0.01fF
C16449 NOR2X1_LOC_772/B INVX1_LOC_92/A 0.07fF
C16450 NAND2X1_LOC_633/Y NAND2X1_LOC_793/Y 0.04fF
C16451 NOR2X1_LOC_414/Y INVX1_LOC_3/A 0.07fF
C16452 NOR2X1_LOC_573/a_36_216# NAND2X1_LOC_463/B 0.00fF
C16453 NOR2X1_LOC_168/Y NOR2X1_LOC_337/Y 0.01fF
C16454 INVX1_LOC_30/A INVX1_LOC_95/A 0.17fF
C16455 INVX1_LOC_182/A NOR2X1_LOC_344/a_36_216# 0.01fF
C16456 INVX1_LOC_161/Y NOR2X1_LOC_682/Y 0.27fF
C16457 INVX1_LOC_5/A NOR2X1_LOC_862/B 0.01fF
C16458 INVX1_LOC_13/Y INVX1_LOC_92/A 0.03fF
C16459 INVX1_LOC_62/Y INVX1_LOC_91/A 0.07fF
C16460 NOR2X1_LOC_416/A INVX1_LOC_63/A 0.05fF
C16461 INVX1_LOC_135/A NAND2X1_LOC_859/B 0.11fF
C16462 NOR2X1_LOC_147/B NOR2X1_LOC_74/A 0.69fF
C16463 INVX1_LOC_89/A NAND2X1_LOC_452/a_36_24# 0.00fF
C16464 INVX1_LOC_249/A NOR2X1_LOC_66/a_36_216# 0.00fF
C16465 NOR2X1_LOC_624/A INPUT_0 0.03fF
C16466 NOR2X1_LOC_596/A INVX1_LOC_91/A 0.09fF
C16467 INVX1_LOC_279/A NOR2X1_LOC_553/B 0.03fF
C16468 NAND2X1_LOC_361/Y INVX1_LOC_92/Y 0.00fF
C16469 NOR2X1_LOC_392/B NOR2X1_LOC_74/A 0.10fF
C16470 INVX1_LOC_89/A INVX1_LOC_316/Y 0.03fF
C16471 INVX1_LOC_171/A NOR2X1_LOC_211/A 0.11fF
C16472 INVX1_LOC_21/A NOR2X1_LOC_155/A 0.08fF
C16473 NOR2X1_LOC_510/Y NOR2X1_LOC_88/Y 0.05fF
C16474 INVX1_LOC_141/Y INVX1_LOC_37/A 0.03fF
C16475 NOR2X1_LOC_214/B INVX1_LOC_22/A 0.99fF
C16476 INVX1_LOC_161/Y NAND2X1_LOC_848/A 0.02fF
C16477 INVX1_LOC_31/A NAND2X1_LOC_721/A 0.46fF
C16478 NOR2X1_LOC_207/a_36_216# INVX1_LOC_290/A 0.01fF
C16479 NOR2X1_LOC_757/A NAND2X1_LOC_656/Y 0.03fF
C16480 NOR2X1_LOC_350/A NOR2X1_LOC_78/A 0.01fF
C16481 NOR2X1_LOC_273/Y INVX1_LOC_199/A 0.03fF
C16482 NOR2X1_LOC_392/B NOR2X1_LOC_9/Y 0.10fF
C16483 INVX1_LOC_229/Y NOR2X1_LOC_299/Y 7.78fF
C16484 INVX1_LOC_2/A INVX1_LOC_42/Y 0.03fF
C16485 INVX1_LOC_106/Y INVX1_LOC_57/A 0.04fF
C16486 NOR2X1_LOC_759/Y INVX1_LOC_199/A 0.03fF
C16487 NOR2X1_LOC_109/Y INVX1_LOC_63/A 0.15fF
C16488 NAND2X1_LOC_213/A NOR2X1_LOC_156/Y 0.04fF
C16489 INVX1_LOC_34/A NOR2X1_LOC_7/Y 0.01fF
C16490 NOR2X1_LOC_291/a_36_216# NAND2X1_LOC_489/Y 0.02fF
C16491 NOR2X1_LOC_6/B INVX1_LOC_48/A 0.01fF
C16492 NOR2X1_LOC_196/A INVX1_LOC_36/Y 0.01fF
C16493 INVX1_LOC_88/A INVX1_LOC_92/A 1.59fF
C16494 INVX1_LOC_249/A NOR2X1_LOC_69/A 0.01fF
C16495 NOR2X1_LOC_158/a_36_216# NOR2X1_LOC_158/Y 0.01fF
C16496 NAND2X1_LOC_554/a_36_24# INVX1_LOC_313/A 0.00fF
C16497 NOR2X1_LOC_168/Y VDD 0.19fF
C16498 NAND2X1_LOC_837/Y INVX1_LOC_20/A 0.07fF
C16499 NOR2X1_LOC_295/Y INVX1_LOC_91/A 0.06fF
C16500 INVX1_LOC_135/A NAND2X1_LOC_861/Y 0.10fF
C16501 INVX1_LOC_208/A INVX1_LOC_75/A 0.10fF
C16502 INVX1_LOC_2/A INVX1_LOC_191/A 0.19fF
C16503 INVX1_LOC_11/A INVX1_LOC_75/Y 0.01fF
C16504 INVX1_LOC_41/Y NAND2X1_LOC_650/B 0.03fF
C16505 NOR2X1_LOC_516/B INVX1_LOC_75/A 0.03fF
C16506 NAND2X1_LOC_562/B NOR2X1_LOC_45/B 0.11fF
C16507 NAND2X1_LOC_708/Y INVX1_LOC_12/A 0.02fF
C16508 NOR2X1_LOC_75/Y NOR2X1_LOC_433/Y 0.01fF
C16509 INVX1_LOC_309/Y INVX1_LOC_46/A 0.04fF
C16510 NOR2X1_LOC_790/B INVX1_LOC_290/Y 0.08fF
C16511 NOR2X1_LOC_546/B INVX1_LOC_37/A 0.06fF
C16512 INVX1_LOC_132/A NOR2X1_LOC_35/Y 0.10fF
C16513 INVX1_LOC_293/A NOR2X1_LOC_78/Y 0.01fF
C16514 NAND2X1_LOC_787/A NOR2X1_LOC_48/B 0.00fF
C16515 NOR2X1_LOC_468/Y NOR2X1_LOC_179/Y 0.02fF
C16516 INVX1_LOC_27/A NOR2X1_LOC_691/B 0.07fF
C16517 INVX1_LOC_2/A INVX1_LOC_125/Y 0.10fF
C16518 NOR2X1_LOC_561/Y NOR2X1_LOC_597/a_36_216# 0.01fF
C16519 NOR2X1_LOC_262/Y VDD 0.23fF
C16520 NOR2X1_LOC_361/Y NOR2X1_LOC_269/Y 0.01fF
C16521 NAND2X1_LOC_231/Y NOR2X1_LOC_7/Y 0.15fF
C16522 NOR2X1_LOC_197/A INVX1_LOC_179/A 0.04fF
C16523 INVX1_LOC_34/A NAND2X1_LOC_212/Y 0.17fF
C16524 INVX1_LOC_39/A NOR2X1_LOC_84/B 0.00fF
C16525 INVX1_LOC_41/A INVX1_LOC_20/A 0.29fF
C16526 NOR2X1_LOC_226/A INVX1_LOC_125/Y 0.06fF
C16527 INVX1_LOC_30/A INVX1_LOC_54/A 2.56fF
C16528 INVX1_LOC_40/Y NOR2X1_LOC_655/Y 0.00fF
C16529 NOR2X1_LOC_361/B INVX1_LOC_84/A 0.01fF
C16530 INVX1_LOC_171/Y INVX1_LOC_29/A 0.13fF
C16531 NOR2X1_LOC_498/Y INVX1_LOC_20/A 0.00fF
C16532 INVX1_LOC_113/Y INVX1_LOC_139/Y 1.75fF
C16533 NAND2X1_LOC_149/Y NOR2X1_LOC_48/Y 0.02fF
C16534 INVX1_LOC_90/A NOR2X1_LOC_356/A 0.07fF
C16535 INVX1_LOC_275/A INVX1_LOC_37/A 0.01fF
C16536 NAND2X1_LOC_21/Y VDD 0.06fF
C16537 INVX1_LOC_189/Y INVX1_LOC_91/A 0.01fF
C16538 INVX1_LOC_1/Y INVX1_LOC_6/A 3.51fF
C16539 NOR2X1_LOC_829/Y NAND2X1_LOC_175/Y 0.04fF
C16540 NOR2X1_LOC_791/Y NAND2X1_LOC_807/B 0.02fF
C16541 NOR2X1_LOC_67/Y NOR2X1_LOC_849/A 0.01fF
C16542 NOR2X1_LOC_220/A INVX1_LOC_91/A 0.10fF
C16543 NOR2X1_LOC_577/Y INVX1_LOC_12/Y 0.10fF
C16544 INVX1_LOC_95/Y NOR2X1_LOC_709/A 0.17fF
C16545 NOR2X1_LOC_78/B NAND2X1_LOC_655/A 0.25fF
C16546 NOR2X1_LOC_843/A NOR2X1_LOC_857/A 0.04fF
C16547 NOR2X1_LOC_773/Y NOR2X1_LOC_45/B 0.07fF
C16548 INVX1_LOC_34/A D_INPUT_3 0.19fF
C16549 INVX1_LOC_312/Y NOR2X1_LOC_743/Y 0.01fF
C16550 NOR2X1_LOC_152/A NOR2X1_LOC_152/Y 0.00fF
C16551 NAND2X1_LOC_464/Y VDD -0.00fF
C16552 INVX1_LOC_34/A INVX1_LOC_14/Y 0.03fF
C16553 INVX1_LOC_240/A INVX1_LOC_76/A 0.02fF
C16554 NOR2X1_LOC_843/B NOR2X1_LOC_621/A 0.03fF
C16555 NAND2X1_LOC_477/A INVX1_LOC_20/A 0.03fF
C16556 NAND2X1_LOC_567/Y NOR2X1_LOC_536/A 0.01fF
C16557 INVX1_LOC_135/A INVX1_LOC_158/Y 0.03fF
C16558 NOR2X1_LOC_551/B INVX1_LOC_117/A 0.03fF
C16559 INVX1_LOC_23/A INVX1_LOC_175/A 0.02fF
C16560 INVX1_LOC_76/Y VDD 0.09fF
C16561 INVX1_LOC_243/Y NOR2X1_LOC_635/B 0.32fF
C16562 NOR2X1_LOC_78/B NAND2X1_LOC_468/B 0.03fF
C16563 NOR2X1_LOC_78/A NOR2X1_LOC_374/B 0.08fF
C16564 INVX1_LOC_26/A INVX1_LOC_29/Y 0.03fF
C16565 INVX1_LOC_266/Y NOR2X1_LOC_586/Y 0.01fF
C16566 NAND2X1_LOC_30/Y INVX1_LOC_19/A 0.02fF
C16567 INVX1_LOC_290/A NOR2X1_LOC_78/A 0.18fF
C16568 INVX1_LOC_30/A NOR2X1_LOC_430/a_36_216# 0.01fF
C16569 NOR2X1_LOC_548/Y INVX1_LOC_91/A 0.02fF
C16570 NAND2X1_LOC_802/A INVX1_LOC_118/A 0.03fF
C16571 NOR2X1_LOC_510/Y INVX1_LOC_15/A 0.09fF
C16572 NAND2X1_LOC_550/A NAND2X1_LOC_478/a_36_24# 0.00fF
C16573 INVX1_LOC_224/A NAND2X1_LOC_74/B 0.07fF
C16574 INVX1_LOC_89/A INVX1_LOC_86/A 0.01fF
C16575 INVX1_LOC_90/A NOR2X1_LOC_74/A 1.10fF
C16576 NOR2X1_LOC_16/Y VDD -0.00fF
C16577 NOR2X1_LOC_756/a_36_216# INVX1_LOC_75/A 0.02fF
C16578 INVX1_LOC_16/A NAND2X1_LOC_642/Y 1.17fF
C16579 NOR2X1_LOC_175/A NAND2X1_LOC_277/a_36_24# 0.00fF
C16580 NAND2X1_LOC_863/B INVX1_LOC_11/Y 0.31fF
C16581 INVX1_LOC_40/Y NOR2X1_LOC_649/B 0.06fF
C16582 NOR2X1_LOC_533/A INVX1_LOC_76/A 0.04fF
C16583 INVX1_LOC_11/A NAND2X1_LOC_74/B 0.14fF
C16584 NOR2X1_LOC_168/B INVX1_LOC_37/A 0.02fF
C16585 NAND2X1_LOC_787/A NOR2X1_LOC_438/Y 0.04fF
C16586 NOR2X1_LOC_389/B NOR2X1_LOC_74/A 0.03fF
C16587 INVX1_LOC_40/Y INVX1_LOC_3/A 0.02fF
C16588 INVX1_LOC_25/A INVX1_LOC_112/Y 0.03fF
C16589 NAND2X1_LOC_177/a_36_24# NAND2X1_LOC_472/Y 0.00fF
C16590 NAND2X1_LOC_860/A INVX1_LOC_181/A 0.53fF
C16591 INVX1_LOC_27/A NOR2X1_LOC_620/a_36_216# 0.02fF
C16592 INVX1_LOC_61/A NAND2X1_LOC_240/a_36_24# 0.01fF
C16593 NOR2X1_LOC_299/Y INVX1_LOC_167/Y 0.25fF
C16594 INVX1_LOC_90/A NOR2X1_LOC_9/Y 0.39fF
C16595 NOR2X1_LOC_192/A INVX1_LOC_164/A 0.02fF
C16596 INVX1_LOC_24/A NAND2X1_LOC_435/a_36_24# 0.00fF
C16597 NOR2X1_LOC_561/Y NOR2X1_LOC_141/a_36_216# 0.01fF
C16598 NOR2X1_LOC_377/Y NOR2X1_LOC_378/Y 0.01fF
C16599 INVX1_LOC_75/A NOR2X1_LOC_706/A 0.11fF
C16600 NOR2X1_LOC_389/B NOR2X1_LOC_9/Y 0.10fF
C16601 INVX1_LOC_303/A INVX1_LOC_92/A 0.07fF
C16602 INPUT_3 INVX1_LOC_29/A 0.06fF
C16603 INVX1_LOC_36/A INVX1_LOC_63/A 2.19fF
C16604 INVX1_LOC_11/A NOR2X1_LOC_847/B 0.00fF
C16605 NAND2X1_LOC_213/A D_INPUT_5 0.13fF
C16606 NOR2X1_LOC_45/Y INVX1_LOC_109/A 0.11fF
C16607 INVX1_LOC_83/A NAND2X1_LOC_655/A 0.01fF
C16608 NAND2X1_LOC_363/B NOR2X1_LOC_836/A 0.46fF
C16609 NAND2X1_LOC_381/Y NOR2X1_LOC_847/B 0.21fF
C16610 NOR2X1_LOC_596/a_36_216# NOR2X1_LOC_155/A 0.00fF
C16611 NOR2X1_LOC_160/B NAND2X1_LOC_291/B 0.03fF
C16612 NOR2X1_LOC_318/B INVX1_LOC_313/A 0.08fF
C16613 NAND2X1_LOC_634/Y NAND2X1_LOC_489/Y 0.02fF
C16614 INVX1_LOC_11/Y NAND2X1_LOC_795/Y 0.01fF
C16615 NOR2X1_LOC_276/Y NOR2X1_LOC_89/A 0.01fF
C16616 INVX1_LOC_77/A NOR2X1_LOC_831/B 0.17fF
C16617 NAND2X1_LOC_342/Y NOR2X1_LOC_536/A 0.02fF
C16618 NAND2X1_LOC_349/B NAND2X1_LOC_211/Y 0.53fF
C16619 INVX1_LOC_35/A INVX1_LOC_271/A 0.03fF
C16620 INVX1_LOC_43/A INVX1_LOC_117/A 0.04fF
C16621 NOR2X1_LOC_68/A NOR2X1_LOC_257/Y 0.03fF
C16622 INVX1_LOC_83/A NAND2X1_LOC_468/B 0.01fF
C16623 NOR2X1_LOC_742/A INVX1_LOC_6/A 0.07fF
C16624 NOR2X1_LOC_545/B INVX1_LOC_148/Y 0.00fF
C16625 INVX1_LOC_12/Y INVX1_LOC_22/A 0.27fF
C16626 NOR2X1_LOC_299/Y INVX1_LOC_20/A 0.03fF
C16627 NOR2X1_LOC_561/Y NOR2X1_LOC_137/Y 0.01fF
C16628 NAND2X1_LOC_722/A INVX1_LOC_54/A 0.94fF
C16629 INVX1_LOC_50/Y NOR2X1_LOC_383/B 0.03fF
C16630 INVX1_LOC_285/Y NOR2X1_LOC_335/B 0.11fF
C16631 D_INPUT_4 NOR2X1_LOC_51/a_36_216# 0.00fF
C16632 NAND2X1_LOC_513/a_36_24# INVX1_LOC_117/A 0.01fF
C16633 NAND2X1_LOC_537/Y INVX1_LOC_94/Y 0.09fF
C16634 NAND2X1_LOC_859/Y NAND2X1_LOC_721/A 0.10fF
C16635 NOR2X1_LOC_298/Y INVX1_LOC_46/A 0.03fF
C16636 NAND2X1_LOC_842/B NOR2X1_LOC_675/A 0.28fF
C16637 NOR2X1_LOC_45/B INVX1_LOC_140/A 0.20fF
C16638 NAND2X1_LOC_175/B NOR2X1_LOC_697/Y 0.02fF
C16639 INVX1_LOC_136/A NOR2X1_LOC_89/A 1.06fF
C16640 NAND2X1_LOC_323/B NOR2X1_LOC_729/A 0.07fF
C16641 INVX1_LOC_72/A NOR2X1_LOC_584/Y 0.18fF
C16642 NAND2X1_LOC_859/B INVX1_LOC_280/A 0.01fF
C16643 INVX1_LOC_28/A NAND2X1_LOC_643/a_36_24# 0.00fF
C16644 INVX1_LOC_30/A NOR2X1_LOC_48/B 0.15fF
C16645 INVX1_LOC_16/A NOR2X1_LOC_271/Y 0.03fF
C16646 INVX1_LOC_124/A NOR2X1_LOC_831/B 0.07fF
C16647 INVX1_LOC_153/Y INVX1_LOC_84/A 0.39fF
C16648 NOR2X1_LOC_804/B INVX1_LOC_63/A 0.02fF
C16649 NOR2X1_LOC_142/Y NAND2X1_LOC_475/Y 0.10fF
C16650 NOR2X1_LOC_123/B NAND2X1_LOC_262/a_36_24# 0.00fF
C16651 INVX1_LOC_41/A NOR2X1_LOC_68/a_36_216# 0.00fF
C16652 INVX1_LOC_132/Y INVX1_LOC_37/A 0.03fF
C16653 INVX1_LOC_49/A INVX1_LOC_19/A 3.33fF
C16654 NOR2X1_LOC_298/Y NOR2X1_LOC_766/Y 0.10fF
C16655 INVX1_LOC_266/A NOR2X1_LOC_383/B 0.00fF
C16656 INVX1_LOC_21/A NOR2X1_LOC_598/B 0.32fF
C16657 NOR2X1_LOC_309/Y NOR2X1_LOC_654/a_36_216# 0.01fF
C16658 NOR2X1_LOC_669/Y INVX1_LOC_57/A 0.06fF
C16659 NOR2X1_LOC_433/A NAND2X1_LOC_74/B 0.07fF
C16660 NAND2X1_LOC_638/Y INVX1_LOC_37/A 0.01fF
C16661 NOR2X1_LOC_318/B INVX1_LOC_6/A 0.07fF
C16662 NOR2X1_LOC_309/Y INVX1_LOC_63/A 0.12fF
C16663 INVX1_LOC_58/A NAND2X1_LOC_579/A 0.02fF
C16664 INVX1_LOC_35/A INVX1_LOC_27/A 0.97fF
C16665 NOR2X1_LOC_91/A NOR2X1_LOC_82/A 0.03fF
C16666 INVX1_LOC_31/A INVX1_LOC_87/A 0.01fF
C16667 INVX1_LOC_21/A INVX1_LOC_97/Y 0.03fF
C16668 INVX1_LOC_177/A INVX1_LOC_84/A 0.03fF
C16669 INVX1_LOC_1/Y INVX1_LOC_131/Y 0.22fF
C16670 NOR2X1_LOC_593/Y NAND2X1_LOC_74/B 0.45fF
C16671 NAND2X1_LOC_763/B NAND2X1_LOC_3/B 0.40fF
C16672 NAND2X1_LOC_361/Y INVX1_LOC_106/A -0.01fF
C16673 NAND2X1_LOC_807/Y NAND2X1_LOC_721/A 0.40fF
C16674 INVX1_LOC_2/A NOR2X1_LOC_653/Y 0.04fF
C16675 INVX1_LOC_93/Y INVX1_LOC_6/A 0.01fF
C16676 NOR2X1_LOC_188/A NAND2X1_LOC_447/Y 0.10fF
C16677 INVX1_LOC_40/A NOR2X1_LOC_820/Y 0.25fF
C16678 NOR2X1_LOC_706/A NAND2X1_LOC_485/a_36_24# 0.00fF
C16679 INVX1_LOC_64/A NAND2X1_LOC_58/a_36_24# 0.00fF
C16680 INVX1_LOC_59/A NAND2X1_LOC_569/B 0.19fF
C16681 NOR2X1_LOC_78/B NOR2X1_LOC_66/Y 0.03fF
C16682 NOR2X1_LOC_729/a_36_216# NOR2X1_LOC_155/A 0.00fF
C16683 NOR2X1_LOC_835/B INVX1_LOC_143/Y 0.24fF
C16684 INVX1_LOC_64/A NOR2X1_LOC_92/Y 0.14fF
C16685 NOR2X1_LOC_770/B INVX1_LOC_12/A 0.01fF
C16686 INVX1_LOC_88/A INVX1_LOC_53/A 0.15fF
C16687 INVX1_LOC_201/Y NOR2X1_LOC_128/A 0.07fF
C16688 INVX1_LOC_50/A NOR2X1_LOC_254/A 0.01fF
C16689 NOR2X1_LOC_68/A NOR2X1_LOC_158/B 0.02fF
C16690 NAND2X1_LOC_721/B NAND2X1_LOC_175/Y -0.02fF
C16691 INVX1_LOC_299/A NOR2X1_LOC_634/Y 0.02fF
C16692 NOR2X1_LOC_82/A INVX1_LOC_23/A 5.58fF
C16693 INVX1_LOC_278/A NOR2X1_LOC_361/B 0.03fF
C16694 INVX1_LOC_64/A INVX1_LOC_24/Y 0.08fF
C16695 INVX1_LOC_134/A INVX1_LOC_23/A 0.03fF
C16696 NAND2X1_LOC_149/Y INVX1_LOC_204/Y 0.05fF
C16697 NOR2X1_LOC_356/A INVX1_LOC_38/A 0.07fF
C16698 NOR2X1_LOC_344/A INVX1_LOC_290/Y 0.42fF
C16699 NOR2X1_LOC_52/B NAND2X1_LOC_74/B 0.08fF
C16700 INPUT_0 D_INPUT_3 0.76fF
C16701 NOR2X1_LOC_631/B INVX1_LOC_78/Y 0.00fF
C16702 INVX1_LOC_184/Y INVX1_LOC_15/A 0.05fF
C16703 INVX1_LOC_2/A INVX1_LOC_19/A 0.08fF
C16704 INVX1_LOC_11/A INVX1_LOC_259/Y 0.03fF
C16705 NOR2X1_LOC_91/A NAND2X1_LOC_500/Y 0.01fF
C16706 INVX1_LOC_135/A INVX1_LOC_291/A 0.10fF
C16707 NOR2X1_LOC_387/A NOR2X1_LOC_422/Y 0.00fF
C16708 NAND2X1_LOC_660/Y NOR2X1_LOC_841/A 0.29fF
C16709 NOR2X1_LOC_278/A NOR2X1_LOC_89/A 0.14fF
C16710 INVX1_LOC_2/A NOR2X1_LOC_11/Y 0.01fF
C16711 NOR2X1_LOC_590/A INVX1_LOC_270/Y 0.28fF
C16712 INVX1_LOC_6/A INVX1_LOC_139/A 0.06fF
C16713 INVX1_LOC_11/A NOR2X1_LOC_660/Y 0.00fF
C16714 INVX1_LOC_64/A NAND2X1_LOC_568/A 0.00fF
C16715 NOR2X1_LOC_226/A INVX1_LOC_19/A 0.09fF
C16716 NOR2X1_LOC_613/Y INVX1_LOC_178/A 0.06fF
C16717 INVX1_LOC_11/A NAND2X1_LOC_358/B 0.02fF
C16718 NAND2X1_LOC_231/Y NOR2X1_LOC_831/Y 0.10fF
C16719 NOR2X1_LOC_135/Y NOR2X1_LOC_331/B 0.00fF
C16720 INVX1_LOC_91/A NAND2X1_LOC_655/B 0.02fF
C16721 NOR2X1_LOC_716/B INVX1_LOC_47/Y 0.01fF
C16722 INVX1_LOC_62/A INVX1_LOC_46/Y 0.04fF
C16723 NAND2X1_LOC_381/Y NOR2X1_LOC_660/Y 0.01fF
C16724 INVX1_LOC_258/A INVX1_LOC_5/A 0.00fF
C16725 NOR2X1_LOC_458/Y INVX1_LOC_15/A -0.01fF
C16726 NOR2X1_LOC_455/Y INVX1_LOC_292/A 0.01fF
C16727 INVX1_LOC_254/Y INVX1_LOC_4/Y 0.02fF
C16728 INVX1_LOC_153/Y INVX1_LOC_15/A 0.01fF
C16729 NAND2X1_LOC_721/A INVX1_LOC_6/A 0.03fF
C16730 VDD INVX1_LOC_123/A 0.03fF
C16731 NOR2X1_LOC_561/A NOR2X1_LOC_74/A 0.01fF
C16732 NAND2X1_LOC_866/B NOR2X1_LOC_823/a_36_216# 0.00fF
C16733 NAND2X1_LOC_794/B NAND2X1_LOC_724/A 0.07fF
C16734 INVX1_LOC_235/Y INVX1_LOC_239/A 1.41fF
C16735 INVX1_LOC_8/A INVX1_LOC_32/A 0.17fF
C16736 INVX1_LOC_78/Y INVX1_LOC_37/A 0.06fF
C16737 NAND2X1_LOC_725/Y NAND2X1_LOC_741/B 0.03fF
C16738 D_INPUT_0 NOR2X1_LOC_841/A 0.10fF
C16739 NAND2X1_LOC_36/A INVX1_LOC_23/A 0.12fF
C16740 NOR2X1_LOC_388/Y NOR2X1_LOC_609/Y 0.03fF
C16741 INVX1_LOC_41/A INVX1_LOC_4/A 0.16fF
C16742 NAND2X1_LOC_276/Y NOR2X1_LOC_38/B 0.03fF
C16743 NAND2X1_LOC_581/Y INVX1_LOC_15/A 0.01fF
C16744 NOR2X1_LOC_74/A INVX1_LOC_38/A 0.62fF
C16745 NAND2X1_LOC_722/A NOR2X1_LOC_48/B 0.21fF
C16746 NAND2X1_LOC_642/Y NOR2X1_LOC_35/Y 0.01fF
C16747 INVX1_LOC_2/A NAND2X1_LOC_227/a_36_24# 0.01fF
C16748 NOR2X1_LOC_445/Y INVX1_LOC_4/Y 0.00fF
C16749 NOR2X1_LOC_828/Y NOR2X1_LOC_778/Y 0.02fF
C16750 NOR2X1_LOC_9/Y INVX1_LOC_38/A 0.03fF
C16751 NAND2X1_LOC_564/B INVX1_LOC_29/A 0.07fF
C16752 INVX1_LOC_177/A INVX1_LOC_15/A 0.03fF
C16753 NAND2X1_LOC_514/Y INVX1_LOC_23/A 0.06fF
C16754 INVX1_LOC_49/A INVX1_LOC_26/Y 0.03fF
C16755 NOR2X1_LOC_15/Y INVX1_LOC_14/A 1.98fF
C16756 GATE_662 INVX1_LOC_29/A 0.01fF
C16757 NAND2X1_LOC_653/a_36_24# INVX1_LOC_117/Y 0.00fF
C16758 NAND2X1_LOC_468/B INVX1_LOC_46/A 0.03fF
C16759 NAND2X1_LOC_11/Y D_INPUT_5 0.02fF
C16760 INVX1_LOC_89/A NOR2X1_LOC_662/A 0.06fF
C16761 D_INPUT_1 NOR2X1_LOC_191/B 0.09fF
C16762 INVX1_LOC_59/A NOR2X1_LOC_530/Y 0.12fF
C16763 NOR2X1_LOC_214/B INVX1_LOC_186/Y 0.31fF
C16764 INVX1_LOC_24/A NOR2X1_LOC_678/A 0.03fF
C16765 NOR2X1_LOC_360/Y INVX1_LOC_138/Y 0.53fF
C16766 INVX1_LOC_5/A NOR2X1_LOC_52/Y 0.00fF
C16767 INVX1_LOC_151/Y INVX1_LOC_32/A 0.01fF
C16768 INVX1_LOC_196/A NOR2X1_LOC_334/Y 1.88fF
C16769 NOR2X1_LOC_168/B NAND2X1_LOC_72/B 0.12fF
C16770 INVX1_LOC_162/A NAND2X1_LOC_286/B 0.00fF
C16771 NAND2X1_LOC_348/A NOR2X1_LOC_243/B 0.09fF
C16772 INPUT_1 INVX1_LOC_19/A 7.08fF
C16773 INVX1_LOC_6/A INVX1_LOC_117/Y 0.11fF
C16774 INVX1_LOC_200/Y NAND2X1_LOC_833/Y 0.02fF
C16775 NOR2X1_LOC_790/B INVX1_LOC_77/A 0.31fF
C16776 NAND2X1_LOC_303/Y INVX1_LOC_161/A 0.51fF
C16777 INVX1_LOC_64/A NAND2X1_LOC_837/Y 0.08fF
C16778 NOR2X1_LOC_753/Y NAND2X1_LOC_793/B 0.03fF
C16779 NAND2X1_LOC_332/Y INVX1_LOC_23/A 0.00fF
C16780 NOR2X1_LOC_261/Y INVX1_LOC_153/Y 0.11fF
C16781 INVX1_LOC_39/A INVX1_LOC_72/Y 0.02fF
C16782 NAND2X1_LOC_59/B INVX1_LOC_53/A 0.10fF
C16783 INVX1_LOC_120/A NAND2X1_LOC_202/a_36_24# 0.00fF
C16784 NOR2X1_LOC_15/Y NOR2X1_LOC_717/Y 0.01fF
C16785 INVX1_LOC_119/A INVX1_LOC_57/A 0.14fF
C16786 NOR2X1_LOC_191/B NOR2X1_LOC_652/Y 0.37fF
C16787 NOR2X1_LOC_785/Y INVX1_LOC_15/A 0.02fF
C16788 NOR2X1_LOC_82/A INVX1_LOC_31/A 0.40fF
C16789 NOR2X1_LOC_456/Y NOR2X1_LOC_181/Y 0.02fF
C16790 INVX1_LOC_285/Y INVX1_LOC_84/A 0.62fF
C16791 INVX1_LOC_41/A INVX1_LOC_64/A 0.03fF
C16792 INVX1_LOC_140/A NOR2X1_LOC_1/Y 0.02fF
C16793 NOR2X1_LOC_498/Y INVX1_LOC_64/A 1.10fF
C16794 GATE_741 NAND2X1_LOC_863/Y 0.03fF
C16795 NAND2X1_LOC_860/A NOR2X1_LOC_315/Y 0.25fF
C16796 NOR2X1_LOC_647/Y INVX1_LOC_269/A 0.05fF
C16797 NOR2X1_LOC_91/A INVX1_LOC_278/Y 0.19fF
C16798 NOR2X1_LOC_471/Y NOR2X1_LOC_478/A 0.14fF
C16799 INVX1_LOC_269/A INVX1_LOC_18/A 0.17fF
C16800 INVX1_LOC_28/A NAND2X1_LOC_792/B 0.07fF
C16801 NOR2X1_LOC_318/B NOR2X1_LOC_117/Y 0.02fF
C16802 NAND2X1_LOC_9/Y NOR2X1_LOC_398/a_36_216# 0.00fF
C16803 NOR2X1_LOC_667/Y NOR2X1_LOC_590/A 0.04fF
C16804 INVX1_LOC_33/A INVX1_LOC_306/Y 0.11fF
C16805 NOR2X1_LOC_232/Y INVX1_LOC_18/A 0.02fF
C16806 NAND2X1_LOC_534/a_36_24# INVX1_LOC_53/A 0.01fF
C16807 INVX1_LOC_10/A NOR2X1_LOC_409/B 0.03fF
C16808 NAND2X1_LOC_67/Y NOR2X1_LOC_735/a_36_216# 0.00fF
C16809 INPUT_0 NOR2X1_LOC_831/Y 0.01fF
C16810 NAND2X1_LOC_650/B INVX1_LOC_185/A 0.01fF
C16811 NAND2X1_LOC_739/B NOR2X1_LOC_15/Y 0.07fF
C16812 INVX1_LOC_136/A INVX1_LOC_11/A 0.05fF
C16813 NOR2X1_LOC_420/Y NAND2X1_LOC_276/Y 0.04fF
C16814 NAND2X1_LOC_350/A INVX1_LOC_30/A 0.07fF
C16815 INVX1_LOC_1/Y INVX1_LOC_28/Y 0.04fF
C16816 INVX1_LOC_17/A NOR2X1_LOC_68/A 0.90fF
C16817 NAND2X1_LOC_84/Y NOR2X1_LOC_15/Y 0.03fF
C16818 NAND2X1_LOC_563/Y NOR2X1_LOC_663/A 0.04fF
C16819 NOR2X1_LOC_456/Y NOR2X1_LOC_778/B 0.01fF
C16820 NOR2X1_LOC_741/A INVX1_LOC_186/Y 0.02fF
C16821 INVX1_LOC_64/A NOR2X1_LOC_398/Y 0.20fF
C16822 NOR2X1_LOC_756/Y INVX1_LOC_3/Y 0.03fF
C16823 NOR2X1_LOC_328/Y NOR2X1_LOC_654/A 0.02fF
C16824 NOR2X1_LOC_203/Y INVX1_LOC_53/A 0.03fF
C16825 INVX1_LOC_5/A NOR2X1_LOC_180/Y 0.03fF
C16826 INVX1_LOC_104/A NOR2X1_LOC_674/a_36_216# 0.00fF
C16827 INVX1_LOC_1/Y INVX1_LOC_270/A 0.17fF
C16828 NOR2X1_LOC_655/B NAND2X1_LOC_363/B 0.01fF
C16829 INVX1_LOC_64/A INVX1_LOC_64/Y 0.05fF
C16830 INVX1_LOC_30/Y NOR2X1_LOC_383/B 0.07fF
C16831 NOR2X1_LOC_612/a_36_216# NOR2X1_LOC_717/A 0.01fF
C16832 NOR2X1_LOC_441/Y INVX1_LOC_30/A 0.12fF
C16833 NOR2X1_LOC_471/Y NOR2X1_LOC_68/A 0.08fF
C16834 INVX1_LOC_230/Y NOR2X1_LOC_791/B 0.17fF
C16835 NOR2X1_LOC_488/a_36_216# NAND2X1_LOC_793/B 0.01fF
C16836 INVX1_LOC_125/Y NAND2X1_LOC_63/Y 0.01fF
C16837 NOR2X1_LOC_667/A NAND2X1_LOC_725/A 0.01fF
C16838 INVX1_LOC_34/A NAND2X1_LOC_705/Y 0.01fF
C16839 NOR2X1_LOC_87/B NOR2X1_LOC_249/Y 0.18fF
C16840 INVX1_LOC_166/A NAND2X1_LOC_462/B 0.01fF
C16841 NOR2X1_LOC_87/B NOR2X1_LOC_846/A 0.01fF
C16842 INVX1_LOC_316/Y NOR2X1_LOC_392/Y 0.07fF
C16843 NOR2X1_LOC_15/Y INVX1_LOC_217/Y 0.03fF
C16844 INVX1_LOC_227/A INVX1_LOC_270/Y 0.06fF
C16845 INVX1_LOC_34/A NAND2X1_LOC_303/Y 0.07fF
C16846 INVX1_LOC_1/A NAND2X1_LOC_139/A 0.01fF
C16847 NOR2X1_LOC_91/A NOR2X1_LOC_132/a_36_216# 0.00fF
C16848 NAND2X1_LOC_218/B NOR2X1_LOC_160/B 0.03fF
C16849 INPUT_3 INVX1_LOC_228/A 0.05fF
C16850 INVX1_LOC_13/Y NOR2X1_LOC_78/B 0.08fF
C16851 INVX1_LOC_197/Y INVX1_LOC_253/Y 0.23fF
C16852 INVX1_LOC_49/A INVX1_LOC_161/Y 0.08fF
C16853 INVX1_LOC_150/A INVX1_LOC_57/A 0.96fF
C16854 NOR2X1_LOC_250/Y NOR2X1_LOC_172/Y 0.02fF
C16855 NOR2X1_LOC_66/Y INVX1_LOC_46/A 0.06fF
C16856 NOR2X1_LOC_631/A INVX1_LOC_76/A 0.03fF
C16857 INVX1_LOC_285/Y INVX1_LOC_15/A 0.03fF
C16858 NAND2X1_LOC_347/B NOR2X1_LOC_316/Y 0.01fF
C16859 INVX1_LOC_40/A INVX1_LOC_306/Y 0.11fF
C16860 NAND2X1_LOC_582/a_36_24# INVX1_LOC_1/A 0.01fF
C16861 NOR2X1_LOC_160/B NOR2X1_LOC_577/Y 0.07fF
C16862 NOR2X1_LOC_433/A NOR2X1_LOC_276/Y 0.05fF
C16863 NOR2X1_LOC_45/B INVX1_LOC_42/A 9.66fF
C16864 NAND2X1_LOC_363/B NAND2X1_LOC_358/Y 0.03fF
C16865 INVX1_LOC_89/A INVX1_LOC_57/A 0.71fF
C16866 NOR2X1_LOC_15/Y NOR2X1_LOC_612/B 0.12fF
C16867 NAND2X1_LOC_214/B NOR2X1_LOC_121/A 0.01fF
C16868 NAND2X1_LOC_455/a_36_24# INVX1_LOC_19/A 0.01fF
C16869 NOR2X1_LOC_296/Y INVX1_LOC_8/A 0.03fF
C16870 INVX1_LOC_233/Y NOR2X1_LOC_32/Y 0.01fF
C16871 NOR2X1_LOC_335/B INVX1_LOC_4/Y 0.08fF
C16872 INVX1_LOC_50/A NOR2X1_LOC_473/B 0.01fF
C16873 NOR2X1_LOC_798/A NOR2X1_LOC_175/a_36_216# 0.00fF
C16874 INVX1_LOC_278/A NOR2X1_LOC_528/a_36_216# 0.01fF
C16875 NOR2X1_LOC_132/a_36_216# INVX1_LOC_23/A 0.02fF
C16876 INVX1_LOC_35/A INVX1_LOC_234/A 0.03fF
C16877 INVX1_LOC_69/Y NAND2X1_LOC_647/B 0.02fF
C16878 NAND2X1_LOC_364/A NOR2X1_LOC_360/Y 0.17fF
C16879 INVX1_LOC_14/A NAND2X1_LOC_141/A 0.02fF
C16880 INVX1_LOC_1/A NAND2X1_LOC_139/a_36_24# 0.00fF
C16881 INVX1_LOC_181/Y INVX1_LOC_72/A 0.00fF
C16882 INVX1_LOC_41/A INVX1_LOC_43/Y 0.24fF
C16883 NAND2X1_LOC_746/a_36_24# NOR2X1_LOC_781/A 0.02fF
C16884 NOR2X1_LOC_586/Y INVX1_LOC_19/A 0.15fF
C16885 NOR2X1_LOC_2/Y NOR2X1_LOC_30/Y 0.01fF
C16886 NAND2X1_LOC_213/A NAND2X1_LOC_451/Y 0.21fF
C16887 INVX1_LOC_45/A INVX1_LOC_180/A 0.05fF
C16888 NOR2X1_LOC_92/Y NAND2X1_LOC_850/Y 0.07fF
C16889 INVX1_LOC_269/A INVX1_LOC_34/Y 0.10fF
C16890 NOR2X1_LOC_536/A INVX1_LOC_285/A 0.15fF
C16891 NAND2X1_LOC_35/Y INVX1_LOC_229/Y 2.73fF
C16892 INVX1_LOC_27/A NOR2X1_LOC_121/A 0.04fF
C16893 INPUT_3 INVX1_LOC_8/A 0.11fF
C16894 NOR2X1_LOC_9/Y NAND2X1_LOC_223/A 0.01fF
C16895 NAND2X1_LOC_541/Y INVX1_LOC_1/A 0.07fF
C16896 INVX1_LOC_230/Y NOR2X1_LOC_124/B 0.04fF
C16897 NAND2X1_LOC_541/a_36_24# INVX1_LOC_89/A 0.00fF
C16898 INVX1_LOC_74/A NOR2X1_LOC_847/B 0.02fF
C16899 INVX1_LOC_113/A INVX1_LOC_54/A 0.01fF
C16900 NOR2X1_LOC_536/A NOR2X1_LOC_814/A 0.02fF
C16901 NAND2X1_LOC_96/A NOR2X1_LOC_721/B 0.01fF
C16902 NOR2X1_LOC_78/B INVX1_LOC_88/A 0.03fF
C16903 NAND2X1_LOC_469/a_36_24# INVX1_LOC_76/A 0.00fF
C16904 NOR2X1_LOC_106/Y INVX1_LOC_79/Y 0.01fF
C16905 INVX1_LOC_136/A NOR2X1_LOC_433/A 0.13fF
C16906 INVX1_LOC_65/A INVX1_LOC_15/A 0.02fF
C16907 NAND2X1_LOC_188/a_36_24# INVX1_LOC_240/A 0.00fF
C16908 INVX1_LOC_20/A INVX1_LOC_168/Y 0.01fF
C16909 INVX1_LOC_50/A NOR2X1_LOC_322/Y 0.05fF
C16910 NOR2X1_LOC_657/Y INVX1_LOC_33/A 0.03fF
C16911 INVX1_LOC_2/A INVX1_LOC_161/Y 0.18fF
C16912 INVX1_LOC_45/A NAND2X1_LOC_325/Y 0.26fF
C16913 NOR2X1_LOC_590/A NOR2X1_LOC_310/Y 0.01fF
C16914 INVX1_LOC_256/A NAND2X1_LOC_342/Y 0.15fF
C16915 NOR2X1_LOC_142/Y INVX1_LOC_30/A 0.19fF
C16916 INVX1_LOC_136/A NOR2X1_LOC_593/Y 0.10fF
C16917 INVX1_LOC_107/Y INVX1_LOC_92/A 0.00fF
C16918 NOR2X1_LOC_653/Y INVX1_LOC_118/A 0.13fF
C16919 NOR2X1_LOC_226/A INVX1_LOC_161/Y 0.03fF
C16920 NAND2X1_LOC_731/Y NAND2X1_LOC_740/A 0.14fF
C16921 INVX1_LOC_35/A NOR2X1_LOC_772/A 0.01fF
C16922 NOR2X1_LOC_45/B INVX1_LOC_78/A 0.34fF
C16923 INVX1_LOC_64/A NOR2X1_LOC_122/Y 0.23fF
C16924 INVX1_LOC_286/Y NOR2X1_LOC_591/Y 0.08fF
C16925 NOR2X1_LOC_655/Y NOR2X1_LOC_814/A 0.03fF
C16926 INVX1_LOC_35/A NOR2X1_LOC_19/B 0.13fF
C16927 NOR2X1_LOC_656/Y INVX1_LOC_63/A 0.05fF
C16928 NOR2X1_LOC_454/Y NOR2X1_LOC_586/a_36_216# 0.01fF
C16929 NAND2X1_LOC_810/B NAND2X1_LOC_770/Y 0.15fF
C16930 NOR2X1_LOC_419/a_36_216# NOR2X1_LOC_419/Y 0.01fF
C16931 INVX1_LOC_170/A NOR2X1_LOC_84/Y 0.03fF
C16932 NOR2X1_LOC_598/B NAND2X1_LOC_51/B 0.07fF
C16933 NOR2X1_LOC_717/Y INVX1_LOC_96/Y 0.68fF
C16934 NAND2X1_LOC_93/B NOR2X1_LOC_814/A 0.03fF
C16935 NOR2X1_LOC_470/a_36_216# INVX1_LOC_117/A 0.01fF
C16936 INVX1_LOC_19/A INVX1_LOC_118/A 0.19fF
C16937 INVX1_LOC_136/A NOR2X1_LOC_52/B 0.11fF
C16938 NAND2X1_LOC_348/A NOR2X1_LOC_342/A 0.00fF
C16939 NOR2X1_LOC_435/A INVX1_LOC_63/A 0.10fF
C16940 INVX1_LOC_132/A NOR2X1_LOC_350/A 0.02fF
C16941 INVX1_LOC_276/A INVX1_LOC_45/A 0.07fF
C16942 NAND2X1_LOC_550/A INVX1_LOC_22/A 0.01fF
C16943 INVX1_LOC_199/Y INVX1_LOC_78/A 0.01fF
C16944 INVX1_LOC_78/A INVX1_LOC_247/A 0.04fF
C16945 NOR2X1_LOC_318/B INVX1_LOC_28/Y 0.00fF
C16946 NOR2X1_LOC_655/B INVX1_LOC_30/A 0.11fF
C16947 NOR2X1_LOC_65/B NOR2X1_LOC_45/B 0.01fF
C16948 NOR2X1_LOC_790/A NOR2X1_LOC_542/Y 0.01fF
C16949 NAND2X1_LOC_577/A NAND2X1_LOC_548/a_36_24# 0.02fF
C16950 NOR2X1_LOC_160/B INVX1_LOC_22/A 0.12fF
C16951 NOR2X1_LOC_646/A INVX1_LOC_230/Y 0.27fF
C16952 NOR2X1_LOC_67/A INVX1_LOC_45/A 0.15fF
C16953 NAND2X1_LOC_833/Y NOR2X1_LOC_495/Y 0.00fF
C16954 NOR2X1_LOC_228/a_36_216# NOR2X1_LOC_716/B 0.00fF
C16955 INVX1_LOC_77/A NOR2X1_LOC_344/A 0.01fF
C16956 INVX1_LOC_88/A INVX1_LOC_83/A 0.03fF
C16957 NAND2X1_LOC_182/A INVX1_LOC_41/Y 0.20fF
C16958 NOR2X1_LOC_318/B INVX1_LOC_270/A 0.10fF
C16959 NOR2X1_LOC_620/A INVX1_LOC_117/A 0.01fF
C16960 INVX1_LOC_64/A NAND2X1_LOC_662/B 0.03fF
C16961 INVX1_LOC_50/A NOR2X1_LOC_562/B 0.73fF
C16962 NOR2X1_LOC_45/Y INVX1_LOC_290/A 0.06fF
C16963 INVX1_LOC_25/A NOR2X1_LOC_78/A 0.18fF
C16964 INVX1_LOC_285/A NOR2X1_LOC_661/A 0.03fF
C16965 NOR2X1_LOC_91/A INVX1_LOC_59/Y 0.03fF
C16966 INVX1_LOC_54/Y NAND2X1_LOC_656/A 0.04fF
C16967 INVX1_LOC_3/A NOR2X1_LOC_814/A 0.09fF
C16968 INVX1_LOC_265/Y NOR2X1_LOC_661/A 0.19fF
C16969 NOR2X1_LOC_631/B NOR2X1_LOC_727/B 0.01fF
C16970 NAND2X1_LOC_581/Y NAND2X1_LOC_21/Y 0.03fF
C16971 NOR2X1_LOC_690/A INVX1_LOC_34/A 0.11fF
C16972 INVX1_LOC_36/A INVX1_LOC_1/Y 0.10fF
C16973 INVX1_LOC_32/A INVX1_LOC_118/Y 0.00fF
C16974 NAND2X1_LOC_329/a_36_24# NOR2X1_LOC_717/A 0.01fF
C16975 INVX1_LOC_237/Y INVX1_LOC_240/A 0.74fF
C16976 INVX1_LOC_34/A NOR2X1_LOC_413/Y 0.09fF
C16977 INVX1_LOC_161/Y NAND2X1_LOC_648/A 0.02fF
C16978 INVX1_LOC_290/A NOR2X1_LOC_584/a_36_216# 0.00fF
C16979 NAND2X1_LOC_564/B NAND2X1_LOC_634/Y 0.00fF
C16980 INVX1_LOC_256/A NOR2X1_LOC_246/Y 0.03fF
C16981 NAND2X1_LOC_287/B NAND2X1_LOC_288/B 0.19fF
C16982 INVX1_LOC_245/Y INVX1_LOC_90/A 0.00fF
C16983 INVX1_LOC_200/Y NAND2X1_LOC_241/Y 0.01fF
C16984 INVX1_LOC_37/A NOR2X1_LOC_727/B 0.03fF
C16985 NOR2X1_LOC_778/B NOR2X1_LOC_550/B 0.01fF
C16986 NAND2X1_LOC_574/A NOR2X1_LOC_128/A 0.03fF
C16987 NOR2X1_LOC_457/A INVX1_LOC_182/A 0.07fF
C16988 NOR2X1_LOC_468/Y NOR2X1_LOC_184/a_36_216# 0.00fF
C16989 INVX1_LOC_83/A NOR2X1_LOC_500/B 0.01fF
C16990 NAND2X1_LOC_303/Y INPUT_0 1.59fF
C16991 NAND2X1_LOC_341/A INVX1_LOC_81/A 0.00fF
C16992 INVX1_LOC_74/A NOR2X1_LOC_660/Y 0.02fF
C16993 INVX1_LOC_208/A NOR2X1_LOC_577/Y 0.37fF
C16994 NAND2X1_LOC_231/Y NAND2X1_LOC_466/Y 0.39fF
C16995 D_INPUT_1 VDD 0.98fF
C16996 INVX1_LOC_41/A NAND2X1_LOC_850/Y 0.02fF
C16997 NAND2X1_LOC_500/Y NAND2X1_LOC_866/B 0.04fF
C16998 INVX1_LOC_269/A NOR2X1_LOC_548/A 0.11fF
C16999 NAND2X1_LOC_63/Y INVX1_LOC_19/A 0.07fF
C17000 NOR2X1_LOC_599/A NAND2X1_LOC_648/A 0.04fF
C17001 NOR2X1_LOC_331/B NAND2X1_LOC_61/Y 0.04fF
C17002 NOR2X1_LOC_496/Y INVX1_LOC_91/A 0.02fF
C17003 INVX1_LOC_33/Y NOR2X1_LOC_654/A 0.25fF
C17004 NOR2X1_LOC_272/Y NOR2X1_LOC_269/Y 0.08fF
C17005 NAND2X1_LOC_198/B NAND2X1_LOC_656/Y 0.10fF
C17006 NOR2X1_LOC_219/Y NOR2X1_LOC_219/B 0.12fF
C17007 NAND2X1_LOC_44/a_36_24# INVX1_LOC_89/A 0.00fF
C17008 NOR2X1_LOC_374/A NOR2X1_LOC_374/B 0.01fF
C17009 NOR2X1_LOC_667/A NAND2X1_LOC_308/Y 0.00fF
C17010 NOR2X1_LOC_574/a_36_216# INVX1_LOC_236/A 0.14fF
C17011 NOR2X1_LOC_214/B INVX1_LOC_18/A 0.07fF
C17012 NAND2X1_LOC_35/Y INVX1_LOC_20/A 0.17fF
C17013 NAND2X1_LOC_569/A INVX1_LOC_25/Y -0.01fF
C17014 NAND2X1_LOC_477/A NAND2X1_LOC_850/Y 0.10fF
C17015 INVX1_LOC_1/A INVX1_LOC_98/A 0.20fF
C17016 NOR2X1_LOC_298/Y NAND2X1_LOC_866/A 1.16fF
C17017 NOR2X1_LOC_299/Y NAND2X1_LOC_863/Y 0.03fF
C17018 NAND2X1_LOC_787/A NOR2X1_LOC_176/Y 0.00fF
C17019 NOR2X1_LOC_172/Y NAND2X1_LOC_660/Y 0.02fF
C17020 NAND2X1_LOC_574/A INVX1_LOC_4/A 0.02fF
C17021 INVX1_LOC_182/A INVX1_LOC_30/A 0.41fF
C17022 NAND2X1_LOC_455/B INVX1_LOC_19/A 0.14fF
C17023 NOR2X1_LOC_82/A INVX1_LOC_6/A 0.10fF
C17024 NOR2X1_LOC_667/A NAND2X1_LOC_660/A 0.00fF
C17025 NOR2X1_LOC_336/B NOR2X1_LOC_567/B 0.06fF
C17026 INVX1_LOC_1/A NOR2X1_LOC_78/A 0.18fF
C17027 INVX1_LOC_303/A INVX1_LOC_83/A 0.07fF
C17028 NAND2X1_LOC_721/A NOR2X1_LOC_109/Y 0.07fF
C17029 INVX1_LOC_210/Y INVX1_LOC_75/A 0.19fF
C17030 NAND2X1_LOC_11/Y NAND2X1_LOC_451/Y 0.09fF
C17031 NOR2X1_LOC_309/Y INVX1_LOC_1/Y 0.09fF
C17032 NAND2X1_LOC_254/Y NAND2X1_LOC_74/B 0.03fF
C17033 INVX1_LOC_28/A NOR2X1_LOC_91/Y 0.03fF
C17034 INVX1_LOC_136/Y INVX1_LOC_4/A 0.10fF
C17035 NOR2X1_LOC_665/A INVX1_LOC_88/Y 0.01fF
C17036 NAND2X1_LOC_182/A NAND2X1_LOC_861/a_36_24# 0.00fF
C17037 INVX1_LOC_13/Y INVX1_LOC_46/A 2.52fF
C17038 INVX1_LOC_64/A NOR2X1_LOC_494/a_36_216# 0.02fF
C17039 VDD NOR2X1_LOC_652/Y 0.94fF
C17040 NOR2X1_LOC_68/A NOR2X1_LOC_171/Y 0.03fF
C17041 INVX1_LOC_84/A INVX1_LOC_4/Y 1.27fF
C17042 INVX1_LOC_274/A NOR2X1_LOC_748/A 0.10fF
C17043 D_INPUT_0 NOR2X1_LOC_172/Y 0.01fF
C17044 NOR2X1_LOC_779/Y NOR2X1_LOC_708/A 0.02fF
C17045 NAND2X1_LOC_59/B INVX1_LOC_83/A 0.54fF
C17046 NOR2X1_LOC_790/B INVX1_LOC_9/A 0.05fF
C17047 INVX1_LOC_35/Y NAND2X1_LOC_99/A 0.01fF
C17048 INVX1_LOC_189/A INVX1_LOC_22/A 0.02fF
C17049 NOR2X1_LOC_503/Y NOR2X1_LOC_45/B 0.00fF
C17050 INVX1_LOC_80/A INVX1_LOC_80/Y -0.00fF
C17051 INVX1_LOC_77/A NOR2X1_LOC_702/Y 0.01fF
C17052 INVX1_LOC_206/A NOR2X1_LOC_188/Y 0.02fF
C17053 INVX1_LOC_310/Y INVX1_LOC_132/Y 0.08fF
C17054 INVX1_LOC_202/A NAND2X1_LOC_123/Y 0.15fF
C17055 INVX1_LOC_13/A NOR2X1_LOC_520/A 0.03fF
C17056 INVX1_LOC_232/Y INVX1_LOC_255/Y 0.14fF
C17057 NOR2X1_LOC_68/A NOR2X1_LOC_594/Y 0.07fF
C17058 INVX1_LOC_33/A NOR2X1_LOC_356/A 0.01fF
C17059 NAND2X1_LOC_93/B NOR2X1_LOC_292/a_36_216# 0.02fF
C17060 NAND2X1_LOC_853/Y INVX1_LOC_22/A 0.04fF
C17061 NOR2X1_LOC_475/a_36_216# INVX1_LOC_255/Y 0.01fF
C17062 INVX1_LOC_277/A INVX1_LOC_186/A 0.04fF
C17063 INVX1_LOC_282/A NAND2X1_LOC_837/Y 0.07fF
C17064 NOR2X1_LOC_215/A INVX1_LOC_281/A 0.02fF
C17065 NOR2X1_LOC_533/Y INVX1_LOC_76/A 0.10fF
C17066 INVX1_LOC_88/A INVX1_LOC_46/A 0.24fF
C17067 INVX1_LOC_36/A NOR2X1_LOC_318/B 0.13fF
C17068 NAND2X1_LOC_359/Y NAND2X1_LOC_359/a_36_24# 0.02fF
C17069 INVX1_LOC_19/A NOR2X1_LOC_631/Y 0.05fF
C17070 NOR2X1_LOC_298/Y NOR2X1_LOC_505/Y 0.01fF
C17071 NOR2X1_LOC_678/A NOR2X1_LOC_197/B 0.03fF
C17072 NOR2X1_LOC_195/A INVX1_LOC_36/Y 0.01fF
C17073 INVX1_LOC_254/A INPUT_0 0.00fF
C17074 NOR2X1_LOC_241/A VDD 0.00fF
C17075 INVX1_LOC_12/A NOR2X1_LOC_409/B 0.03fF
C17076 INVX1_LOC_35/A NOR2X1_LOC_216/B 0.03fF
C17077 INVX1_LOC_75/A INVX1_LOC_155/A 0.01fF
C17078 NOR2X1_LOC_789/B INVX1_LOC_9/A 0.01fF
C17079 NAND2X1_LOC_338/B INVX1_LOC_148/Y 0.05fF
C17080 INVX1_LOC_31/A INVX1_LOC_59/Y 0.07fF
C17081 INVX1_LOC_36/A INVX1_LOC_93/Y 0.08fF
C17082 NAND2X1_LOC_63/Y INVX1_LOC_26/Y 0.92fF
C17083 INVX1_LOC_33/A NOR2X1_LOC_74/A 3.18fF
C17084 INVX1_LOC_230/Y INVX1_LOC_2/Y 0.03fF
C17085 INVX1_LOC_31/A INVX1_LOC_176/A 0.03fF
C17086 NAND2X1_LOC_656/Y INVX1_LOC_53/Y 0.10fF
C17087 NOR2X1_LOC_267/A INVX1_LOC_93/Y 0.10fF
C17088 INVX1_LOC_50/Y INVX1_LOC_179/A 0.05fF
C17089 NOR2X1_LOC_467/a_36_216# NOR2X1_LOC_470/A 0.01fF
C17090 NAND2X1_LOC_218/B INVX1_LOC_315/Y 0.00fF
C17091 NOR2X1_LOC_360/Y NOR2X1_LOC_405/A 4.19fF
C17092 INVX1_LOC_21/A INVX1_LOC_152/A 0.07fF
C17093 NOR2X1_LOC_201/A NOR2X1_LOC_340/A 0.15fF
C17094 INVX1_LOC_230/Y NAND2X1_LOC_129/a_36_24# 0.00fF
C17095 INVX1_LOC_145/A NOR2X1_LOC_318/B 0.01fF
C17096 INVX1_LOC_33/A NOR2X1_LOC_9/Y 0.07fF
C17097 INVX1_LOC_15/A INVX1_LOC_4/Y 0.07fF
C17098 INVX1_LOC_29/A NAND2X1_LOC_97/a_36_24# 0.01fF
C17099 INVX1_LOC_64/A NOR2X1_LOC_23/a_36_216# 0.00fF
C17100 INVX1_LOC_172/Y NAND2X1_LOC_624/A 0.00fF
C17101 NAND2X1_LOC_656/Y NOR2X1_LOC_665/A 0.01fF
C17102 INVX1_LOC_233/Y INVX1_LOC_84/A 0.01fF
C17103 INVX1_LOC_90/A NAND2X1_LOC_319/a_36_24# 0.00fF
C17104 NAND2X1_LOC_327/a_36_24# NAND2X1_LOC_660/A 0.01fF
C17105 NOR2X1_LOC_392/Y NOR2X1_LOC_662/A 0.07fF
C17106 NAND2X1_LOC_803/B NOR2X1_LOC_536/A 0.02fF
C17107 NOR2X1_LOC_250/Y INVX1_LOC_38/A 0.43fF
C17108 NAND2X1_LOC_783/Y INVX1_LOC_33/Y 0.01fF
C17109 NOR2X1_LOC_45/B NOR2X1_LOC_152/Y 0.18fF
C17110 NOR2X1_LOC_273/Y NOR2X1_LOC_657/B 0.01fF
C17111 NOR2X1_LOC_555/a_36_216# INVX1_LOC_113/Y 0.00fF
C17112 NOR2X1_LOC_759/Y NOR2X1_LOC_657/B 0.01fF
C17113 NOR2X1_LOC_298/Y NOR2X1_LOC_700/Y 0.03fF
C17114 INVX1_LOC_208/A NOR2X1_LOC_735/Y 0.07fF
C17115 INVX1_LOC_198/A INVX1_LOC_92/A -0.04fF
C17116 INVX1_LOC_53/A INVX1_LOC_272/A 0.07fF
C17117 NAND2X1_LOC_754/a_36_24# NOR2X1_LOC_356/A 0.00fF
C17118 NOR2X1_LOC_350/A NAND2X1_LOC_642/Y 0.25fF
C17119 NOR2X1_LOC_590/A NOR2X1_LOC_536/A 0.12fF
C17120 INVX1_LOC_161/Y INVX1_LOC_118/A 0.10fF
C17121 NOR2X1_LOC_103/Y NAND2X1_LOC_268/a_36_24# 0.00fF
C17122 INVX1_LOC_278/A NAND2X1_LOC_81/B 0.07fF
C17123 INVX1_LOC_30/A NOR2X1_LOC_176/Y 0.30fF
C17124 NOR2X1_LOC_778/A VDD 0.00fF
C17125 INVX1_LOC_63/Y INVX1_LOC_91/A 0.03fF
C17126 NOR2X1_LOC_6/a_36_216# NAND2X1_LOC_642/Y 0.00fF
C17127 NOR2X1_LOC_68/A NOR2X1_LOC_706/B 0.01fF
C17128 NOR2X1_LOC_781/A NAND2X1_LOC_654/B 0.00fF
C17129 INVX1_LOC_18/A INVX1_LOC_12/Y 0.18fF
C17130 INVX1_LOC_199/Y INVX1_LOC_113/Y 0.01fF
C17131 NOR2X1_LOC_30/Y NOR2X1_LOC_36/A 0.11fF
C17132 INVX1_LOC_30/A NAND2X1_LOC_61/a_36_24# 0.00fF
C17133 NOR2X1_LOC_208/Y INVX1_LOC_139/A 0.00fF
C17134 INVX1_LOC_120/A NAND2X1_LOC_45/Y 0.03fF
C17135 NOR2X1_LOC_394/Y INVX1_LOC_23/Y 0.03fF
C17136 D_INPUT_0 INVX1_LOC_90/A 0.26fF
C17137 INVX1_LOC_256/A NOR2X1_LOC_364/A 0.22fF
C17138 NOR2X1_LOC_403/B VDD 0.03fF
C17139 NOR2X1_LOC_521/Y NAND2X1_LOC_560/A 0.01fF
C17140 D_INPUT_2 VDD 0.79fF
C17141 NOR2X1_LOC_89/A NOR2X1_LOC_665/Y 0.12fF
C17142 NOR2X1_LOC_792/B NOR2X1_LOC_405/A 0.03fF
C17143 NAND2X1_LOC_579/a_36_24# INVX1_LOC_282/A 0.00fF
C17144 NOR2X1_LOC_151/a_36_216# INVX1_LOC_16/A 0.00fF
C17145 INVX1_LOC_39/A INVX1_LOC_19/A 0.03fF
C17146 NOR2X1_LOC_607/Y VDD 0.24fF
C17147 NOR2X1_LOC_309/Y INVX1_LOC_93/Y 0.10fF
C17148 NOR2X1_LOC_643/Y D_INPUT_3 0.05fF
C17149 NOR2X1_LOC_577/Y NAND2X1_LOC_211/Y 0.08fF
C17150 NOR2X1_LOC_590/A NAND2X1_LOC_93/B 0.03fF
C17151 NOR2X1_LOC_53/Y INVX1_LOC_42/A 0.00fF
C17152 NOR2X1_LOC_430/A INVX1_LOC_37/A 0.03fF
C17153 NOR2X1_LOC_637/B NAND2X1_LOC_453/A 0.03fF
C17154 NOR2X1_LOC_32/B INVX1_LOC_3/Y 0.12fF
C17155 NAND2X1_LOC_364/Y INVX1_LOC_37/A 0.03fF
C17156 INVX1_LOC_230/Y NOR2X1_LOC_608/Y 0.05fF
C17157 INVX1_LOC_21/A INVX1_LOC_29/A 12.34fF
C17158 NOR2X1_LOC_205/Y INVX1_LOC_84/A 0.03fF
C17159 NOR2X1_LOC_237/Y NAND2X1_LOC_721/A 0.06fF
C17160 INVX1_LOC_256/A INVX1_LOC_285/A 0.27fF
C17161 INVX1_LOC_136/A NOR2X1_LOC_675/a_36_216# 0.00fF
C17162 NOR2X1_LOC_299/Y INVX1_LOC_282/A 0.11fF
C17163 NAND2X1_LOC_175/B INVX1_LOC_37/A 0.07fF
C17164 NAND2X1_LOC_302/a_36_24# INVX1_LOC_140/A 0.00fF
C17165 NOR2X1_LOC_234/Y INVX1_LOC_20/A 0.05fF
C17166 INVX1_LOC_266/Y NAND2X1_LOC_212/Y 0.02fF
C17167 D_INPUT_0 NAND2X1_LOC_348/A 0.04fF
C17168 NOR2X1_LOC_844/Y NOR2X1_LOC_862/B 0.13fF
C17169 INVX1_LOC_256/A NOR2X1_LOC_814/A 0.50fF
C17170 INVX1_LOC_27/A NAND2X1_LOC_206/B 0.01fF
C17171 NOR2X1_LOC_25/Y INVX1_LOC_296/Y 0.09fF
C17172 INVX1_LOC_113/Y INVX1_LOC_281/A 0.00fF
C17173 NOR2X1_LOC_510/Y NOR2X1_LOC_677/a_36_216# 0.03fF
C17174 NOR2X1_LOC_591/Y VDD 0.43fF
C17175 NOR2X1_LOC_590/A INVX1_LOC_3/A 0.09fF
C17176 NOR2X1_LOC_309/Y NAND2X1_LOC_721/A 0.99fF
C17177 NOR2X1_LOC_188/a_36_216# INVX1_LOC_91/A 0.00fF
C17178 INVX1_LOC_306/A INVX1_LOC_6/A 0.00fF
C17179 NOR2X1_LOC_591/Y NAND2X1_LOC_800/A 0.03fF
C17180 NAND2X1_LOC_725/B INVX1_LOC_284/A 0.07fF
C17181 NOR2X1_LOC_529/Y VDD 0.24fF
C17182 NAND2X1_LOC_364/A NOR2X1_LOC_79/Y 0.08fF
C17183 INVX1_LOC_266/Y INVX1_LOC_14/Y 0.07fF
C17184 NOR2X1_LOC_720/B INVX1_LOC_117/A 0.02fF
C17185 NOR2X1_LOC_160/B INVX1_LOC_186/Y 0.07fF
C17186 NAND2X1_LOC_354/B NOR2X1_LOC_536/A 0.04fF
C17187 NAND2X1_LOC_860/A NAND2X1_LOC_99/A 0.01fF
C17188 INVX1_LOC_28/A NAND2X1_LOC_811/a_36_24# 0.00fF
C17189 NAND2X1_LOC_30/Y INPUT_7 0.09fF
C17190 NOR2X1_LOC_171/Y INVX1_LOC_147/A 0.00fF
C17191 NOR2X1_LOC_324/B NOR2X1_LOC_325/A 0.01fF
C17192 NOR2X1_LOC_344/A INVX1_LOC_9/A 0.02fF
C17193 NOR2X1_LOC_203/Y INVX1_LOC_46/A 0.03fF
C17194 INVX1_LOC_14/A NOR2X1_LOC_128/a_36_216# 0.01fF
C17195 INVX1_LOC_12/Y INVX1_LOC_34/Y 0.10fF
C17196 NOR2X1_LOC_370/a_36_216# INVX1_LOC_91/A 0.00fF
C17197 INVX1_LOC_56/Y INVX1_LOC_76/A 0.03fF
C17198 INVX1_LOC_180/A NOR2X1_LOC_592/B 0.01fF
C17199 NOR2X1_LOC_45/B NAND2X1_LOC_861/Y 0.08fF
C17200 NAND2X1_LOC_618/Y NOR2X1_LOC_474/a_36_216# 0.00fF
C17201 NOR2X1_LOC_103/Y NAND2X1_LOC_445/a_36_24# 0.00fF
C17202 NOR2X1_LOC_392/Y INVX1_LOC_57/A 0.07fF
C17203 INVX1_LOC_22/A NAND2X1_LOC_211/Y 0.09fF
C17204 INVX1_LOC_31/A NOR2X1_LOC_340/A 0.03fF
C17205 NOR2X1_LOC_140/A NOR2X1_LOC_38/B 0.03fF
C17206 INVX1_LOC_58/A NOR2X1_LOC_32/B 0.03fF
C17207 NOR2X1_LOC_553/Y VDD 0.27fF
C17208 NOR2X1_LOC_613/Y INVX1_LOC_78/A 0.02fF
C17209 NOR2X1_LOC_205/Y INVX1_LOC_15/A 0.03fF
C17210 NOR2X1_LOC_718/Y INVX1_LOC_179/A 0.01fF
C17211 INVX1_LOC_133/Y NOR2X1_LOC_331/B 0.02fF
C17212 INVX1_LOC_75/A INVX1_LOC_86/A 0.00fF
C17213 INVX1_LOC_58/A NOR2X1_LOC_639/B 0.02fF
C17214 INVX1_LOC_21/A INVX1_LOC_298/Y 0.02fF
C17215 NOR2X1_LOC_272/Y INVX1_LOC_26/A 0.03fF
C17216 NAND2X1_LOC_66/a_36_24# NOR2X1_LOC_536/A 0.00fF
C17217 NOR2X1_LOC_788/B NOR2X1_LOC_552/A 0.02fF
C17218 NOR2X1_LOC_632/Y INVX1_LOC_139/Y 0.01fF
C17219 INVX1_LOC_33/A NOR2X1_LOC_865/Y 0.15fF
C17220 INVX1_LOC_49/A NAND2X1_LOC_426/a_36_24# -0.01fF
C17221 NOR2X1_LOC_315/Y NOR2X1_LOC_487/Y 0.01fF
C17222 INVX1_LOC_49/A NOR2X1_LOC_801/A 0.01fF
C17223 INVX1_LOC_33/A NOR2X1_LOC_243/B 0.01fF
C17224 NOR2X1_LOC_82/Y NOR2X1_LOC_536/A 0.00fF
C17225 NOR2X1_LOC_210/B INVX1_LOC_114/A 0.25fF
C17226 NAND2X1_LOC_99/a_36_24# INVX1_LOC_27/Y 0.01fF
C17227 NAND2X1_LOC_752/a_36_24# INVX1_LOC_38/A 0.00fF
C17228 NOR2X1_LOC_140/a_36_216# NAND2X1_LOC_141/Y 0.01fF
C17229 INVX1_LOC_302/Y INVX1_LOC_91/A 0.04fF
C17230 NOR2X1_LOC_123/B NOR2X1_LOC_558/A 0.01fF
C17231 INVX1_LOC_25/A NOR2X1_LOC_186/Y 0.06fF
C17232 NOR2X1_LOC_82/A NOR2X1_LOC_80/Y 0.27fF
C17233 INVX1_LOC_136/A NAND2X1_LOC_254/Y 0.10fF
C17234 INVX1_LOC_9/Y INVX1_LOC_118/Y 0.13fF
C17235 NOR2X1_LOC_78/B NOR2X1_LOC_99/Y 0.03fF
C17236 INVX1_LOC_64/A NAND2X1_LOC_35/Y 6.36fF
C17237 NOR2X1_LOC_647/A INVX1_LOC_269/A 0.01fF
C17238 NOR2X1_LOC_68/A NOR2X1_LOC_346/A 0.01fF
C17239 NOR2X1_LOC_272/Y NOR2X1_LOC_255/Y 0.02fF
C17240 NAND2X1_LOC_796/B NAND2X1_LOC_784/A 0.29fF
C17241 NAND2X1_LOC_9/Y INVX1_LOC_13/Y 0.08fF
C17242 NAND2X1_LOC_660/Y INVX1_LOC_38/A 0.01fF
C17243 NOR2X1_LOC_357/Y D_GATE_366 0.03fF
C17244 NOR2X1_LOC_763/Y NAND2X1_LOC_639/A 0.55fF
C17245 NOR2X1_LOC_791/Y INVX1_LOC_308/A 0.19fF
C17246 INVX1_LOC_314/Y NAND2X1_LOC_74/B 0.05fF
C17247 NOR2X1_LOC_78/A NOR2X1_LOC_188/A 0.03fF
C17248 NOR2X1_LOC_15/Y NOR2X1_LOC_383/B 0.13fF
C17249 INVX1_LOC_2/A NOR2X1_LOC_841/A 0.10fF
C17250 INVX1_LOC_35/A INVX1_LOC_93/A 0.07fF
C17251 NOR2X1_LOC_91/A INVX1_LOC_103/A 0.07fF
C17252 NOR2X1_LOC_78/A NOR2X1_LOC_548/B 0.01fF
C17253 NOR2X1_LOC_644/A NOR2X1_LOC_858/B 0.01fF
C17254 NAND2X1_LOC_53/Y NOR2X1_LOC_302/A 0.02fF
C17255 NOR2X1_LOC_385/Y INVX1_LOC_76/A 0.02fF
C17256 INVX1_LOC_120/Y NOR2X1_LOC_865/Y 0.05fF
C17257 NOR2X1_LOC_497/Y VDD 0.12fF
C17258 NAND2X1_LOC_733/Y NOR2X1_LOC_409/B 0.03fF
C17259 NAND2X1_LOC_738/B NOR2X1_LOC_15/Y 0.00fF
C17260 NOR2X1_LOC_92/Y NOR2X1_LOC_629/A 0.06fF
C17261 NOR2X1_LOC_131/Y NOR2X1_LOC_155/A 0.02fF
C17262 D_INPUT_0 INVX1_LOC_38/A 0.97fF
C17263 NOR2X1_LOC_772/B NOR2X1_LOC_798/A 0.02fF
C17264 NAND2X1_LOC_862/A NOR2X1_LOC_88/Y 0.07fF
C17265 INVX1_LOC_144/A INVX1_LOC_147/Y 0.01fF
C17266 NOR2X1_LOC_317/B NOR2X1_LOC_777/B 0.05fF
C17267 INVX1_LOC_258/Y NAND2X1_LOC_725/A 0.03fF
C17268 NAND2X1_LOC_787/A NAND2X1_LOC_579/A 0.01fF
C17269 D_INPUT_1 NOR2X1_LOC_361/B 0.10fF
C17270 NAND2X1_LOC_357/A INVX1_LOC_57/A 0.03fF
C17271 INVX1_LOC_103/A INVX1_LOC_23/A 0.15fF
C17272 NOR2X1_LOC_160/B NOR2X1_LOC_843/B 0.17fF
C17273 NOR2X1_LOC_392/Y NOR2X1_LOC_475/A 0.06fF
C17274 INVX1_LOC_90/A NAND2X1_LOC_848/A 0.27fF
C17275 NAND2X1_LOC_79/Y INVX1_LOC_32/A 0.07fF
C17276 INVX1_LOC_266/A NOR2X1_LOC_405/Y 0.02fF
C17277 NOR2X1_LOC_798/A INVX1_LOC_13/Y 0.03fF
C17278 NAND2X1_LOC_819/Y NOR2X1_LOC_649/B 0.04fF
C17279 NOR2X1_LOC_92/Y NAND2X1_LOC_624/B 0.07fF
C17280 NOR2X1_LOC_589/A NOR2X1_LOC_155/A 0.15fF
C17281 NOR2X1_LOC_83/Y INVX1_LOC_20/A 0.14fF
C17282 INVX1_LOC_227/A NAND2X1_LOC_93/B 0.07fF
C17283 NOR2X1_LOC_52/Y INVX1_LOC_78/A 0.09fF
C17284 INVX1_LOC_287/A NOR2X1_LOC_160/B 0.06fF
C17285 INVX1_LOC_279/A NOR2X1_LOC_830/a_36_216# 0.00fF
C17286 INVX1_LOC_232/A NAND2X1_LOC_572/B 0.03fF
C17287 INVX1_LOC_94/A INVX1_LOC_4/A 0.07fF
C17288 NOR2X1_LOC_168/Y INVX1_LOC_4/Y 0.03fF
C17289 NOR2X1_LOC_68/A INVX1_LOC_94/Y 0.03fF
C17290 INVX1_LOC_269/A NAND2X1_LOC_533/a_36_24# 0.00fF
C17291 NAND2X1_LOC_862/A INVX1_LOC_84/A 0.04fF
C17292 NOR2X1_LOC_83/a_36_216# INVX1_LOC_46/A 0.00fF
C17293 INVX1_LOC_13/A INVX1_LOC_123/Y 0.01fF
C17294 INVX1_LOC_157/A NOR2X1_LOC_364/A 0.02fF
C17295 NAND2X1_LOC_198/B INVX1_LOC_128/Y 0.04fF
C17296 NOR2X1_LOC_561/Y NOR2X1_LOC_831/B 0.04fF
C17297 NAND2X1_LOC_348/A NOR2X1_LOC_859/Y 0.01fF
C17298 INVX1_LOC_89/A INVX1_LOC_274/A 0.08fF
C17299 NOR2X1_LOC_337/A INVX1_LOC_37/A 0.03fF
C17300 INVX1_LOC_150/Y INVX1_LOC_53/A 0.14fF
C17301 INVX1_LOC_292/A INVX1_LOC_23/A 0.10fF
C17302 NOR2X1_LOC_383/Y NAND2X1_LOC_572/B 0.15fF
C17303 D_INPUT_0 NAND2X1_LOC_848/Y 0.03fF
C17304 NAND2X1_LOC_364/A INVX1_LOC_26/A 0.00fF
C17305 INVX1_LOC_25/Y NOR2X1_LOC_662/A 0.01fF
C17306 INVX1_LOC_196/Y INVX1_LOC_307/Y 0.04fF
C17307 NOR2X1_LOC_78/B INVX1_LOC_272/A 0.07fF
C17308 NOR2X1_LOC_186/Y INVX1_LOC_1/A 0.02fF
C17309 NAND2X1_LOC_276/Y INVX1_LOC_251/A 0.08fF
C17310 INVX1_LOC_1/Y INVX1_LOC_63/A 0.19fF
C17311 INVX1_LOC_49/A INVX1_LOC_128/A 0.01fF
C17312 NOR2X1_LOC_667/A INVX1_LOC_29/A 0.02fF
C17313 NOR2X1_LOC_361/B NOR2X1_LOC_652/Y 0.22fF
C17314 NOR2X1_LOC_843/A INVX1_LOC_15/A 0.09fF
C17315 NOR2X1_LOC_346/B NAND2X1_LOC_207/B 0.09fF
C17316 INVX1_LOC_90/A INVX1_LOC_46/Y 0.03fF
C17317 NAND2X1_LOC_725/B NOR2X1_LOC_384/A 0.12fF
C17318 NOR2X1_LOC_68/A INVX1_LOC_296/A 0.15fF
C17319 INVX1_LOC_177/Y INVX1_LOC_270/Y 0.11fF
C17320 NOR2X1_LOC_790/B NOR2X1_LOC_565/A 0.01fF
C17321 INVX1_LOC_290/A NOR2X1_LOC_48/Y 0.04fF
C17322 NAND2X1_LOC_9/Y NOR2X1_LOC_500/B 0.02fF
C17323 NOR2X1_LOC_68/A NAND2X1_LOC_205/a_36_24# 0.00fF
C17324 NOR2X1_LOC_468/Y NAND2X1_LOC_346/a_36_24# 0.01fF
C17325 INPUT_5 NOR2X1_LOC_11/Y 0.07fF
C17326 NOR2X1_LOC_759/Y INVX1_LOC_271/A 0.07fF
C17327 NAND2X1_LOC_348/A INVX1_LOC_46/Y 0.04fF
C17328 NOR2X1_LOC_309/Y INVX1_LOC_87/A 0.03fF
C17329 INVX1_LOC_202/A INVX1_LOC_271/A 0.07fF
C17330 NOR2X1_LOC_97/A NOR2X1_LOC_61/A 0.04fF
C17331 NOR2X1_LOC_16/Y INVX1_LOC_4/Y 0.05fF
C17332 INVX1_LOC_2/A INVX1_LOC_128/A -0.02fF
C17333 INVX1_LOC_58/A NOR2X1_LOC_447/Y 0.13fF
C17334 NOR2X1_LOC_641/B INVX1_LOC_50/Y 0.44fF
C17335 NOR2X1_LOC_624/A INVX1_LOC_26/Y 0.00fF
C17336 INVX1_LOC_56/Y INVX1_LOC_127/Y 0.03fF
C17337 INVX1_LOC_83/A INVX1_LOC_272/A 0.10fF
C17338 INVX1_LOC_158/Y NOR2X1_LOC_862/B 0.01fF
C17339 INVX1_LOC_5/A NOR2X1_LOC_703/B 0.03fF
C17340 INVX1_LOC_50/A NAND2X1_LOC_833/Y 0.02fF
C17341 NOR2X1_LOC_798/A NOR2X1_LOC_500/B 0.03fF
C17342 INVX1_LOC_35/A NOR2X1_LOC_500/A 0.05fF
C17343 NOR2X1_LOC_751/Y INVX1_LOC_50/Y 0.45fF
C17344 NOR2X1_LOC_91/A INVX1_LOC_240/A 0.03fF
C17345 INVX1_LOC_35/A NOR2X1_LOC_303/Y 0.03fF
C17346 NAND2X1_LOC_624/B NAND2X1_LOC_837/Y 0.02fF
C17347 INVX1_LOC_41/A INVX1_LOC_129/A 0.03fF
C17348 NOR2X1_LOC_458/B INVX1_LOC_78/A 0.02fF
C17349 NOR2X1_LOC_556/a_36_216# INVX1_LOC_44/A 0.00fF
C17350 INVX1_LOC_85/A NAND2X1_LOC_299/a_36_24# 0.00fF
C17351 NOR2X1_LOC_598/B INVX1_LOC_153/A 0.01fF
C17352 D_INPUT_1 INVX1_LOC_153/Y 0.09fF
C17353 INVX1_LOC_176/Y INVX1_LOC_57/A 0.02fF
C17354 NOR2X1_LOC_45/B INVX1_LOC_291/A 0.08fF
C17355 NAND2X1_LOC_53/Y NOR2X1_LOC_471/Y 0.02fF
C17356 INVX1_LOC_104/A INVX1_LOC_270/Y 0.10fF
C17357 NOR2X1_LOC_667/A NOR2X1_LOC_281/Y 0.02fF
C17358 NAND2X1_LOC_650/B NOR2X1_LOC_536/A 0.91fF
C17359 NOR2X1_LOC_713/a_36_216# NAND2X1_LOC_425/Y 0.01fF
C17360 NOR2X1_LOC_561/A NOR2X1_LOC_266/B 0.00fF
C17361 NAND2X1_LOC_579/A INVX1_LOC_30/A 0.08fF
C17362 INVX1_LOC_96/Y NOR2X1_LOC_383/B 0.01fF
C17363 INVX1_LOC_289/Y INVX1_LOC_36/A 0.01fF
C17364 INVX1_LOC_57/Y NOR2X1_LOC_15/Y 0.04fF
C17365 NOR2X1_LOC_357/Y NOR2X1_LOC_142/a_36_216# 0.01fF
C17366 NOR2X1_LOC_273/Y INVX1_LOC_27/A 0.03fF
C17367 INVX1_LOC_256/A NOR2X1_LOC_590/A 0.07fF
C17368 NAND2X1_LOC_725/B INVX1_LOC_72/A 0.03fF
C17369 NAND2X1_LOC_662/Y NOR2X1_LOC_158/Y 0.07fF
C17370 INVX1_LOC_27/A NOR2X1_LOC_759/Y 0.03fF
C17371 INVX1_LOC_69/Y NOR2X1_LOC_814/A 0.08fF
C17372 D_INPUT_1 INVX1_LOC_177/A 0.09fF
C17373 INVX1_LOC_202/A INVX1_LOC_27/A 0.96fF
C17374 INVX1_LOC_279/A NOR2X1_LOC_334/Y 0.01fF
C17375 NAND2X1_LOC_656/A NAND2X1_LOC_473/A 0.24fF
C17376 INVX1_LOC_299/A NOR2X1_LOC_68/A 0.35fF
C17377 NAND2X1_LOC_53/Y NAND2X1_LOC_16/a_36_24# 0.00fF
C17378 NAND2X1_LOC_51/B INVX1_LOC_29/A 0.00fF
C17379 INVX1_LOC_36/A NOR2X1_LOC_82/A 0.06fF
C17380 NOR2X1_LOC_186/Y NAND2X1_LOC_601/a_36_24# 0.00fF
C17381 NAND2X1_LOC_241/a_36_24# NAND2X1_LOC_244/A 0.00fF
C17382 NOR2X1_LOC_598/B INVX1_LOC_259/A 0.03fF
C17383 NOR2X1_LOC_732/A INVX1_LOC_213/A 0.04fF
C17384 NOR2X1_LOC_744/Y NAND2X1_LOC_780/Y 0.20fF
C17385 NOR2X1_LOC_516/B NOR2X1_LOC_843/B 0.69fF
C17386 INVX1_LOC_233/A INVX1_LOC_168/A 0.04fF
C17387 INVX1_LOC_91/A INVX1_LOC_27/Y 0.02fF
C17388 NOR2X1_LOC_538/B NOR2X1_LOC_68/A 0.03fF
C17389 NOR2X1_LOC_692/a_36_216# NOR2X1_LOC_692/Y 0.00fF
C17390 VDD NOR2X1_LOC_61/Y 0.02fF
C17391 NOR2X1_LOC_92/Y NOR2X1_LOC_617/Y 0.02fF
C17392 INVX1_LOC_269/A NOR2X1_LOC_607/A 0.00fF
C17393 NOR2X1_LOC_590/A NOR2X1_LOC_606/Y 0.00fF
C17394 INVX1_LOC_316/Y NOR2X1_LOC_529/a_36_216# 0.00fF
C17395 NAND2X1_LOC_491/a_36_24# NOR2X1_LOC_717/A 0.00fF
C17396 INVX1_LOC_11/A NAND2X1_LOC_588/B 0.05fF
C17397 INVX1_LOC_35/A INVX1_LOC_54/Y 0.52fF
C17398 D_INPUT_0 NAND2X1_LOC_223/A 0.03fF
C17399 NOR2X1_LOC_750/A INVX1_LOC_32/A 0.03fF
C17400 NAND2X1_LOC_848/A INVX1_LOC_38/A 0.01fF
C17401 NOR2X1_LOC_92/Y NAND2X1_LOC_593/Y 0.03fF
C17402 INVX1_LOC_25/Y INVX1_LOC_57/A 0.28fF
C17403 NAND2X1_LOC_550/A INVX1_LOC_18/A 0.07fF
C17404 NAND2X1_LOC_149/Y INVX1_LOC_275/A 0.31fF
C17405 INVX1_LOC_37/A NOR2X1_LOC_640/Y 0.02fF
C17406 NOR2X1_LOC_403/B NOR2X1_LOC_361/B 0.01fF
C17407 NOR2X1_LOC_647/Y NOR2X1_LOC_160/B 0.46fF
C17408 NAND2X1_LOC_573/Y NAND2X1_LOC_601/a_36_24# 0.00fF
C17409 NOR2X1_LOC_831/B INVX1_LOC_76/A 0.10fF
C17410 NOR2X1_LOC_510/B NAND2X1_LOC_453/A 0.02fF
C17411 INVX1_LOC_21/A INVX1_LOC_8/A 0.01fF
C17412 INVX1_LOC_293/A NOR2X1_LOC_68/A 0.02fF
C17413 INVX1_LOC_41/A NOR2X1_LOC_440/B 0.03fF
C17414 NOR2X1_LOC_160/B INVX1_LOC_18/A 0.14fF
C17415 NOR2X1_LOC_599/Y NOR2X1_LOC_599/a_36_216# 0.01fF
C17416 NOR2X1_LOC_2/Y NOR2X1_LOC_157/a_36_216# 0.00fF
C17417 INVX1_LOC_132/A INVX1_LOC_1/A 0.17fF
C17418 NAND2X1_LOC_848/A NOR2X1_LOC_96/Y 0.02fF
C17419 INVX1_LOC_1/A NOR2X1_LOC_374/A 0.10fF
C17420 INVX1_LOC_93/Y INVX1_LOC_63/A 0.19fF
C17421 NAND2X1_LOC_803/B NOR2X1_LOC_781/Y 0.01fF
C17422 INVX1_LOC_27/A INVX1_LOC_249/Y 0.01fF
C17423 INVX1_LOC_107/Y INVX1_LOC_46/A 0.03fF
C17424 INVX1_LOC_64/A NOR2X1_LOC_136/Y 0.16fF
C17425 INVX1_LOC_53/Y NOR2X1_LOC_717/A 0.07fF
C17426 NOR2X1_LOC_557/A NAND2X1_LOC_74/B 0.03fF
C17427 NOR2X1_LOC_689/A NOR2X1_LOC_576/B 0.05fF
C17428 NOR2X1_LOC_689/Y INVX1_LOC_229/Y 0.10fF
C17429 NOR2X1_LOC_563/a_36_216# INVX1_LOC_53/A 0.01fF
C17430 NOR2X1_LOC_722/Y NOR2X1_LOC_717/Y 0.11fF
C17431 NAND2X1_LOC_729/Y NAND2X1_LOC_389/a_36_24# 0.00fF
C17432 NAND2X1_LOC_739/B INVX1_LOC_161/A 0.49fF
C17433 NOR2X1_LOC_401/B INVX1_LOC_306/Y 0.03fF
C17434 INVX1_LOC_95/Y NAND2X1_LOC_773/B 0.93fF
C17435 NAND2X1_LOC_303/Y NAND2X1_LOC_811/Y 0.03fF
C17436 NOR2X1_LOC_71/Y NOR2X1_LOC_72/Y 0.06fF
C17437 INVX1_LOC_34/A INVX1_LOC_14/A 0.28fF
C17438 NOR2X1_LOC_201/A INVX1_LOC_120/A 0.02fF
C17439 INVX1_LOC_37/A NOR2X1_LOC_697/Y 0.02fF
C17440 NOR2X1_LOC_598/B NOR2X1_LOC_589/A 0.08fF
C17441 INVX1_LOC_182/Y NOR2X1_LOC_334/Y -0.04fF
C17442 INVX1_LOC_172/A NAND2X1_LOC_550/A 0.07fF
C17443 INVX1_LOC_225/A INVX1_LOC_1/A 0.01fF
C17444 NOR2X1_LOC_402/a_36_216# INVX1_LOC_306/Y 0.02fF
C17445 NOR2X1_LOC_211/Y NOR2X1_LOC_211/A 0.00fF
C17446 NOR2X1_LOC_178/Y INVX1_LOC_56/Y 0.03fF
C17447 NOR2X1_LOC_250/Y INVX1_LOC_33/A 0.00fF
C17448 NAND2X1_LOC_578/B INVX1_LOC_178/A 0.38fF
C17449 NOR2X1_LOC_815/Y INVX1_LOC_161/Y 0.04fF
C17450 NOR2X1_LOC_496/Y NAND2X1_LOC_374/Y 0.03fF
C17451 INVX1_LOC_304/A INVX1_LOC_29/A 0.07fF
C17452 NOR2X1_LOC_687/Y INVX1_LOC_213/A 3.29fF
C17453 NAND2X1_LOC_195/Y INVX1_LOC_18/A -0.01fF
C17454 NOR2X1_LOC_83/Y INVX1_LOC_4/A 0.46fF
C17455 INVX1_LOC_38/A INVX1_LOC_46/Y 0.41fF
C17456 INVX1_LOC_45/A INVX1_LOC_181/Y 0.07fF
C17457 NAND2X1_LOC_738/B NOR2X1_LOC_576/B 0.35fF
C17458 NOR2X1_LOC_468/Y NOR2X1_LOC_709/A 0.02fF
C17459 NOR2X1_LOC_393/a_36_216# INVX1_LOC_26/A 0.00fF
C17460 NOR2X1_LOC_302/Y NOR2X1_LOC_302/A 0.10fF
C17461 NOR2X1_LOC_209/Y INVX1_LOC_1/A 0.01fF
C17462 NOR2X1_LOC_356/A NOR2X1_LOC_748/A 0.10fF
C17463 D_INPUT_3 INVX1_LOC_19/A 0.07fF
C17464 NOR2X1_LOC_337/A NAND2X1_LOC_72/B 0.01fF
C17465 INVX1_LOC_14/Y INVX1_LOC_19/A 0.07fF
C17466 INVX1_LOC_110/Y NOR2X1_LOC_340/Y 0.01fF
C17467 NAND2X1_LOC_231/Y INVX1_LOC_14/A 0.01fF
C17468 INVX1_LOC_136/A INVX1_LOC_314/Y 0.10fF
C17469 INVX1_LOC_46/A INVX1_LOC_272/A 0.15fF
C17470 INVX1_LOC_123/A INVX1_LOC_4/Y 0.10fF
C17471 INVX1_LOC_239/A INVX1_LOC_239/Y 0.04fF
C17472 NOR2X1_LOC_52/Y NOR2X1_LOC_152/Y 0.01fF
C17473 NOR2X1_LOC_595/Y INVX1_LOC_15/A 0.03fF
C17474 INVX1_LOC_298/Y INVX1_LOC_311/A 0.07fF
C17475 NAND2X1_LOC_573/A NOR2X1_LOC_652/Y 0.10fF
C17476 INVX1_LOC_50/A INVX1_LOC_73/A 0.06fF
C17477 INVX1_LOC_11/A NAND2X1_LOC_342/Y 0.00fF
C17478 INVX1_LOC_34/A NOR2X1_LOC_717/Y 0.03fF
C17479 INVX1_LOC_24/A NOR2X1_LOC_238/Y 0.03fF
C17480 INVX1_LOC_232/Y NOR2X1_LOC_817/Y 0.00fF
C17481 NOR2X1_LOC_272/Y INVX1_LOC_164/A 0.10fF
C17482 NOR2X1_LOC_391/Y INVX1_LOC_16/Y 0.37fF
C17483 NOR2X1_LOC_295/a_36_216# INVX1_LOC_30/A 0.12fF
C17484 INVX1_LOC_75/A INVX1_LOC_57/A 18.40fF
C17485 NOR2X1_LOC_15/Y NAND2X1_LOC_170/A 0.03fF
C17486 INVX1_LOC_286/A NOR2X1_LOC_278/Y 0.01fF
C17487 NOR2X1_LOC_2/Y INVX1_LOC_296/A 0.14fF
C17488 INVX1_LOC_41/A INVX1_LOC_142/A 0.03fF
C17489 NAND2X1_LOC_552/A INVX1_LOC_183/Y 0.34fF
C17490 NOR2X1_LOC_160/B INVX1_LOC_34/Y 0.23fF
C17491 NOR2X1_LOC_74/A INVX1_LOC_275/Y 0.00fF
C17492 INVX1_LOC_249/A NOR2X1_LOC_759/Y 0.25fF
C17493 INVX1_LOC_35/A NOR2X1_LOC_112/Y 0.02fF
C17494 NOR2X1_LOC_641/B NOR2X1_LOC_6/B 0.14fF
C17495 NOR2X1_LOC_74/A NOR2X1_LOC_748/A 0.11fF
C17496 NOR2X1_LOC_617/Y NAND2X1_LOC_837/Y 0.02fF
C17497 NOR2X1_LOC_732/A NOR2X1_LOC_707/B 0.01fF
C17498 INVX1_LOC_19/A INVX1_LOC_230/A 0.07fF
C17499 INVX1_LOC_17/A NOR2X1_LOC_500/Y 0.03fF
C17500 INVX1_LOC_17/A INVX1_LOC_226/Y 0.12fF
C17501 INVX1_LOC_255/Y NOR2X1_LOC_381/Y 0.11fF
C17502 NOR2X1_LOC_647/B NAND2X1_LOC_819/Y 0.04fF
C17503 INVX1_LOC_21/A NAND2X1_LOC_140/A 0.00fF
C17504 NOR2X1_LOC_751/Y NOR2X1_LOC_6/B 0.01fF
C17505 NOR2X1_LOC_292/Y INVX1_LOC_29/Y 0.21fF
C17506 NOR2X1_LOC_124/A INVX1_LOC_165/A 0.04fF
C17507 INVX1_LOC_34/A NOR2X1_LOC_522/Y 0.19fF
C17508 NOR2X1_LOC_644/A INVX1_LOC_50/Y 0.03fF
C17509 INVX1_LOC_13/A NOR2X1_LOC_296/a_36_216# 0.00fF
C17510 INVX1_LOC_41/A INVX1_LOC_41/Y 0.01fF
C17511 NAND2X1_LOC_739/B INVX1_LOC_34/A 0.03fF
C17512 D_INPUT_1 INVX1_LOC_285/Y 0.03fF
C17513 NOR2X1_LOC_67/Y NOR2X1_LOC_536/A 0.04fF
C17514 INVX1_LOC_95/A NOR2X1_LOC_278/Y 0.03fF
C17515 NOR2X1_LOC_598/B INVX1_LOC_222/A 0.02fF
C17516 NOR2X1_LOC_791/Y NOR2X1_LOC_756/Y 0.03fF
C17517 NAND2X1_LOC_35/Y INVX1_LOC_282/A 0.14fF
C17518 INVX1_LOC_17/A INVX1_LOC_10/A 0.18fF
C17519 NOR2X1_LOC_172/Y INVX1_LOC_49/A 0.06fF
C17520 INVX1_LOC_13/A INPUT_2 0.06fF
C17521 NOR2X1_LOC_577/Y INVX1_LOC_155/A 0.01fF
C17522 NAND2X1_LOC_149/Y NAND2X1_LOC_638/Y 0.06fF
C17523 INVX1_LOC_24/A NOR2X1_LOC_574/A 0.01fF
C17524 INVX1_LOC_39/Y INVX1_LOC_16/A 0.02fF
C17525 NAND2X1_LOC_721/B INVX1_LOC_248/A -0.02fF
C17526 NAND2X1_LOC_561/a_36_24# INVX1_LOC_309/A 0.00fF
C17527 INVX1_LOC_83/A NOR2X1_LOC_740/Y 0.01fF
C17528 NAND2X1_LOC_364/Y INVX1_LOC_310/Y 0.57fF
C17529 INVX1_LOC_256/A INVX1_LOC_227/A 0.10fF
C17530 NOR2X1_LOC_213/a_36_216# INVX1_LOC_18/A 0.00fF
C17531 NOR2X1_LOC_147/B INVX1_LOC_49/A 0.04fF
C17532 INVX1_LOC_17/Y NAND2X1_LOC_623/B 0.04fF
C17533 NOR2X1_LOC_658/Y NOR2X1_LOC_219/Y 0.03fF
C17534 NOR2X1_LOC_77/a_36_216# NAND2X1_LOC_93/B 0.00fF
C17535 INPUT_5 NOR2X1_LOC_22/a_36_216# -0.00fF
C17536 NOR2X1_LOC_419/Y NAND2X1_LOC_116/A 0.03fF
C17537 NAND2X1_LOC_10/a_36_24# INVX1_LOC_48/A 0.01fF
C17538 INVX1_LOC_101/Y INVX1_LOC_313/Y 0.32fF
C17539 NOR2X1_LOC_446/A NOR2X1_LOC_717/B 0.01fF
C17540 INVX1_LOC_33/A NOR2X1_LOC_121/Y 0.05fF
C17541 NOR2X1_LOC_337/Y NOR2X1_LOC_678/A 0.00fF
C17542 NAND2X1_LOC_198/B INVX1_LOC_256/Y 0.24fF
C17543 VDD NOR2X1_LOC_34/Y 0.24fF
C17544 INVX1_LOC_75/A INVX1_LOC_252/A 0.02fF
C17545 INVX1_LOC_25/A NAND2X1_LOC_642/Y 0.07fF
C17546 NOR2X1_LOC_141/a_36_216# INVX1_LOC_23/A 0.02fF
C17547 NOR2X1_LOC_607/Y INVX1_LOC_177/A 0.01fF
C17548 NOR2X1_LOC_186/Y NOR2X1_LOC_188/A 0.00fF
C17549 NOR2X1_LOC_647/Y NOR2X1_LOC_516/B 0.02fF
C17550 NAND2X1_LOC_472/Y INVX1_LOC_271/Y 0.03fF
C17551 NAND2X1_LOC_169/Y NOR2X1_LOC_167/Y 0.11fF
C17552 NOR2X1_LOC_272/Y NOR2X1_LOC_368/A 0.01fF
C17553 NOR2X1_LOC_561/Y INVX1_LOC_81/Y 0.02fF
C17554 INVX1_LOC_11/A NOR2X1_LOC_246/Y 0.04fF
C17555 NAND2X1_LOC_537/Y NOR2X1_LOC_329/B 0.07fF
C17556 D_INPUT_1 INVX1_LOC_316/A 0.49fF
C17557 VDD NOR2X1_LOC_318/A 0.11fF
C17558 NOR2X1_LOC_542/B INVX1_LOC_23/A 0.00fF
C17559 NAND2X1_LOC_796/B NOR2X1_LOC_527/Y 0.01fF
C17560 D_INPUT_1 NOR2X1_LOC_137/B 0.06fF
C17561 NOR2X1_LOC_724/Y NOR2X1_LOC_307/A 0.03fF
C17562 NOR2X1_LOC_433/A NAND2X1_LOC_342/Y 0.29fF
C17563 NOR2X1_LOC_68/A INVX1_LOC_268/Y 0.01fF
C17564 NOR2X1_LOC_760/a_36_216# INVX1_LOC_313/Y 0.00fF
C17565 NOR2X1_LOC_500/A INVX1_LOC_305/Y 0.02fF
C17566 INVX1_LOC_235/Y NAND2X1_LOC_622/B 0.02fF
C17567 NOR2X1_LOC_183/a_36_216# NOR2X1_LOC_652/Y 0.08fF
C17568 NOR2X1_LOC_486/a_36_216# INVX1_LOC_89/A 0.02fF
C17569 INVX1_LOC_2/A NOR2X1_LOC_172/Y 0.14fF
C17570 INVX1_LOC_23/A INVX1_LOC_143/Y 0.03fF
C17571 INVX1_LOC_120/A INVX1_LOC_31/A 0.06fF
C17572 INVX1_LOC_178/A INVX1_LOC_309/A 0.05fF
C17573 INVX1_LOC_166/A D_GATE_479 0.02fF
C17574 INVX1_LOC_5/A INVX1_LOC_91/A 0.34fF
C17575 NOR2X1_LOC_89/A INVX1_LOC_285/A 0.07fF
C17576 INVX1_LOC_57/A NAND2X1_LOC_453/A 0.07fF
C17577 NOR2X1_LOC_295/Y NOR2X1_LOC_709/A 0.01fF
C17578 INVX1_LOC_176/A NOR2X1_LOC_416/A 0.01fF
C17579 NOR2X1_LOC_226/A NOR2X1_LOC_172/Y 0.01fF
C17580 NOR2X1_LOC_598/B INVX1_LOC_20/A 0.04fF
C17581 NOR2X1_LOC_194/Y INVX1_LOC_266/Y 0.02fF
C17582 INVX1_LOC_14/A INPUT_0 10.23fF
C17583 NOR2X1_LOC_89/A NOR2X1_LOC_814/A 0.03fF
C17584 NOR2X1_LOC_78/B NOR2X1_LOC_770/B 0.03fF
C17585 INVX1_LOC_5/A INVX1_LOC_11/Y 0.03fF
C17586 NAND2X1_LOC_123/Y NOR2X1_LOC_276/Y 0.00fF
C17587 NOR2X1_LOC_155/A INVX1_LOC_4/A 0.03fF
C17588 INVX1_LOC_178/A INVX1_LOC_91/A 0.10fF
C17589 NOR2X1_LOC_831/Y INVX1_LOC_19/A 0.06fF
C17590 NOR2X1_LOC_494/Y INVX1_LOC_309/A 0.01fF
C17591 NOR2X1_LOC_226/A NOR2X1_LOC_392/B 0.10fF
C17592 NAND2X1_LOC_578/B NAND2X1_LOC_562/B 0.06fF
C17593 NOR2X1_LOC_716/B INVX1_LOC_232/A 0.10fF
C17594 NOR2X1_LOC_214/B NAND2X1_LOC_16/Y 0.01fF
C17595 INVX1_LOC_28/A INVX1_LOC_141/Y 1.47fF
C17596 NAND2X1_LOC_342/Y NOR2X1_LOC_52/B 0.00fF
C17597 NOR2X1_LOC_520/A INVX1_LOC_158/A 0.11fF
C17598 NAND2X1_LOC_725/A INVX1_LOC_20/A 0.19fF
C17599 NOR2X1_LOC_640/Y NAND2X1_LOC_72/B 0.06fF
C17600 VDD NOR2X1_LOC_678/A 0.80fF
C17601 NOR2X1_LOC_596/Y NOR2X1_LOC_151/Y 0.01fF
C17602 INVX1_LOC_55/Y INVX1_LOC_223/A -0.00fF
C17603 INVX1_LOC_103/A INVX1_LOC_6/A 0.16fF
C17604 VDD INVX1_LOC_295/Y 0.32fF
C17605 NAND2X1_LOC_338/B NOR2X1_LOC_398/a_36_216# 0.00fF
C17606 INVX1_LOC_181/Y NOR2X1_LOC_123/B 0.02fF
C17607 NAND2X1_LOC_223/A INVX1_LOC_46/Y 0.07fF
C17608 NAND2X1_LOC_702/a_36_24# INVX1_LOC_76/A 0.01fF
C17609 NOR2X1_LOC_383/Y NOR2X1_LOC_716/B 0.01fF
C17610 INVX1_LOC_16/A INVX1_LOC_88/Y 0.11fF
C17611 NAND2X1_LOC_738/B NAND2X1_LOC_770/a_36_24# 0.01fF
C17612 INVX1_LOC_207/A NOR2X1_LOC_32/Y 0.00fF
C17613 INVX1_LOC_25/A NOR2X1_LOC_271/Y 0.82fF
C17614 INVX1_LOC_133/Y NOR2X1_LOC_366/B 0.19fF
C17615 NOR2X1_LOC_84/a_36_216# INVX1_LOC_316/Y 0.01fF
C17616 INVX1_LOC_292/Y INVX1_LOC_117/A 0.00fF
C17617 INVX1_LOC_1/A NAND2X1_LOC_642/Y 0.03fF
C17618 INVX1_LOC_255/Y NOR2X1_LOC_6/B 0.19fF
C17619 NOR2X1_LOC_279/a_36_216# NOR2X1_LOC_773/Y 0.01fF
C17620 NOR2X1_LOC_710/A NOR2X1_LOC_711/A 0.00fF
C17621 NOR2X1_LOC_789/B INVX1_LOC_76/A 0.03fF
C17622 INVX1_LOC_104/Y NOR2X1_LOC_814/A 0.04fF
C17623 NOR2X1_LOC_590/A INVX1_LOC_69/Y 0.30fF
C17624 NOR2X1_LOC_652/a_36_216# NOR2X1_LOC_717/A 0.12fF
C17625 INVX1_LOC_170/Y NAND2X1_LOC_74/B 0.01fF
C17626 NOR2X1_LOC_553/Y INVX1_LOC_177/A 0.01fF
C17627 NOR2X1_LOC_175/a_36_216# NOR2X1_LOC_537/Y 0.00fF
C17628 NAND2X1_LOC_364/Y NAND2X1_LOC_367/B 0.01fF
C17629 NAND2X1_LOC_367/A NAND2X1_LOC_363/Y 0.00fF
C17630 D_INPUT_0 INVX1_LOC_33/A 0.11fF
C17631 NAND2X1_LOC_337/B INVX1_LOC_91/A 0.45fF
C17632 INVX1_LOC_5/A NOR2X1_LOC_698/Y 0.01fF
C17633 NOR2X1_LOC_48/Y NOR2X1_LOC_467/A 0.02fF
C17634 NAND2X1_LOC_661/B INVX1_LOC_22/A 0.01fF
C17635 NOR2X1_LOC_770/B INVX1_LOC_83/A 0.05fF
C17636 INVX1_LOC_90/A INVX1_LOC_49/A 0.10fF
C17637 NOR2X1_LOC_816/A INVX1_LOC_91/A 2.44fF
C17638 INVX1_LOC_67/A INVX1_LOC_313/A 0.21fF
C17639 INVX1_LOC_181/Y INVX1_LOC_102/Y 0.94fF
C17640 NAND2X1_LOC_769/a_36_24# INVX1_LOC_49/A 0.00fF
C17641 NOR2X1_LOC_389/B INVX1_LOC_49/A 0.07fF
C17642 INVX1_LOC_87/A INVX1_LOC_63/A 0.10fF
C17643 NAND2X1_LOC_783/A NOR2X1_LOC_574/A 0.02fF
C17644 INVX1_LOC_77/A NOR2X1_LOC_564/Y 0.03fF
C17645 NOR2X1_LOC_520/B NOR2X1_LOC_560/A -0.02fF
C17646 NOR2X1_LOC_246/A INVX1_LOC_162/Y 0.02fF
C17647 NOR2X1_LOC_360/Y NOR2X1_LOC_335/B 0.10fF
C17648 NAND2X1_LOC_9/Y NOR2X1_LOC_99/Y 0.05fF
C17649 NOR2X1_LOC_706/A NOR2X1_LOC_713/B 0.17fF
C17650 NAND2X1_LOC_739/B INPUT_0 0.03fF
C17651 NOR2X1_LOC_216/a_36_216# INVX1_LOC_33/A 0.00fF
C17652 NOR2X1_LOC_248/A INVX1_LOC_29/A 0.01fF
C17653 NOR2X1_LOC_392/B INPUT_1 0.01fF
C17654 NOR2X1_LOC_229/Y INVX1_LOC_22/A 0.22fF
C17655 NOR2X1_LOC_229/a_36_216# INVX1_LOC_290/A 0.01fF
C17656 INVX1_LOC_240/A NAND2X1_LOC_866/B 0.10fF
C17657 INVX1_LOC_35/A NAND2X1_LOC_656/B 0.01fF
C17658 D_GATE_741 INVX1_LOC_76/A 1.51fF
C17659 INVX1_LOC_276/A INVX1_LOC_135/A 0.10fF
C17660 INVX1_LOC_21/A INVX1_LOC_118/Y 0.05fF
C17661 NAND2X1_LOC_114/B NOR2X1_LOC_35/Y 0.10fF
C17662 INVX1_LOC_64/A NOR2X1_LOC_155/A 2.35fF
C17663 NOR2X1_LOC_67/A INVX1_LOC_135/A 0.19fF
C17664 NAND2X1_LOC_736/Y NOR2X1_LOC_380/Y 0.02fF
C17665 GATE_579 VDD 0.14fF
C17666 NAND2X1_LOC_352/B INVX1_LOC_76/A 0.10fF
C17667 INVX1_LOC_15/A D_INPUT_5 0.01fF
C17668 INVX1_LOC_150/Y INVX1_LOC_46/A 0.09fF
C17669 NOR2X1_LOC_448/Y INVX1_LOC_38/A 0.10fF
C17670 INVX1_LOC_2/A INVX1_LOC_90/A 1.07fF
C17671 INVX1_LOC_132/A NOR2X1_LOC_188/A 0.10fF
C17672 NOR2X1_LOC_372/A INVX1_LOC_20/A 0.04fF
C17673 INVX1_LOC_47/A INVX1_LOC_143/A 0.01fF
C17674 D_INPUT_0 INVX1_LOC_40/A 0.15fF
C17675 INVX1_LOC_2/A NOR2X1_LOC_389/B 0.01fF
C17676 INVX1_LOC_45/A NOR2X1_LOC_833/Y 0.26fF
C17677 NAND2X1_LOC_807/B NOR2X1_LOC_278/Y 0.17fF
C17678 INVX1_LOC_1/A NOR2X1_LOC_271/Y 0.01fF
C17679 INVX1_LOC_132/A NOR2X1_LOC_548/B 0.10fF
C17680 INVX1_LOC_55/A VDD -0.00fF
C17681 NAND2X1_LOC_656/Y INVX1_LOC_16/A 0.07fF
C17682 NOR2X1_LOC_226/A INVX1_LOC_90/A 6.92fF
C17683 NAND2X1_LOC_634/Y INVX1_LOC_304/A 0.03fF
C17684 NAND2X1_LOC_555/Y INVX1_LOC_178/Y 0.00fF
C17685 NOR2X1_LOC_157/a_36_216# NOR2X1_LOC_36/A 0.00fF
C17686 NOR2X1_LOC_226/A NOR2X1_LOC_389/B 0.07fF
C17687 NOR2X1_LOC_544/A INVX1_LOC_313/Y 0.02fF
C17688 INVX1_LOC_67/A INVX1_LOC_6/A 0.03fF
C17689 NOR2X1_LOC_294/Y NOR2X1_LOC_35/Y 0.34fF
C17690 NOR2X1_LOC_329/a_36_216# NOR2X1_LOC_329/Y 0.00fF
C17691 NOR2X1_LOC_52/B INVX1_LOC_67/Y 0.02fF
C17692 NOR2X1_LOC_67/A NOR2X1_LOC_490/Y 0.15fF
C17693 INVX1_LOC_282/Y NOR2X1_LOC_380/Y 4.24fF
C17694 INVX1_LOC_225/A NOR2X1_LOC_188/A 0.01fF
C17695 NAND2X1_LOC_30/Y INVX1_LOC_38/A 0.01fF
C17696 INVX1_LOC_271/A NAND2X1_LOC_74/B 0.03fF
C17697 NOR2X1_LOC_383/B INVX1_LOC_99/A 0.06fF
C17698 INVX1_LOC_232/A NOR2X1_LOC_130/Y 0.01fF
C17699 NOR2X1_LOC_546/a_36_216# INVX1_LOC_91/A 0.00fF
C17700 D_INPUT_1 NAND2X1_LOC_81/B 0.10fF
C17701 INVX1_LOC_2/A NAND2X1_LOC_348/A 0.00fF
C17702 INVX1_LOC_24/A INVX1_LOC_95/Y 0.00fF
C17703 NAND2X1_LOC_357/B NOR2X1_LOC_167/Y 0.05fF
C17704 NOR2X1_LOC_493/B NOR2X1_LOC_74/A 0.06fF
C17705 NOR2X1_LOC_536/a_36_216# NAND2X1_LOC_811/Y 0.00fF
C17706 NAND2X1_LOC_562/B INVX1_LOC_309/A 0.02fF
C17707 INVX1_LOC_5/A INVX1_LOC_203/A 0.03fF
C17708 NOR2X1_LOC_15/Y INVX1_LOC_179/A 0.03fF
C17709 NAND2X1_LOC_349/a_36_24# INVX1_LOC_28/A 0.01fF
C17710 INVX1_LOC_305/A VDD 0.00fF
C17711 NAND2X1_LOC_214/B INVX1_LOC_293/Y -0.09fF
C17712 NOR2X1_LOC_607/Y NOR2X1_LOC_137/B 0.21fF
C17713 NAND2X1_LOC_30/Y NOR2X1_LOC_51/A 0.37fF
C17714 NOR2X1_LOC_419/Y NAND2X1_LOC_447/Y 0.01fF
C17715 INVX1_LOC_71/A INVX1_LOC_115/A 0.03fF
C17716 INVX1_LOC_24/A NOR2X1_LOC_305/Y 0.07fF
C17717 NOR2X1_LOC_516/B INVX1_LOC_31/Y 0.19fF
C17718 NOR2X1_LOC_377/Y INVX1_LOC_91/A 0.00fF
C17719 NAND2X1_LOC_863/A NAND2X1_LOC_863/B 0.24fF
C17720 INVX1_LOC_35/A NOR2X1_LOC_610/Y 0.06fF
C17721 NAND2X1_LOC_562/B INVX1_LOC_91/A 0.02fF
C17722 INVX1_LOC_178/A INVX1_LOC_203/A 0.15fF
C17723 NOR2X1_LOC_716/B NAND2X1_LOC_447/Y 0.02fF
C17724 INVX1_LOC_27/A INVX1_LOC_293/Y 0.08fF
C17725 NOR2X1_LOC_557/Y INVX1_LOC_95/Y 0.06fF
C17726 NOR2X1_LOC_68/A NAND2X1_LOC_96/A 0.14fF
C17727 NAND2X1_LOC_207/a_36_24# NAND2X1_LOC_207/Y 0.01fF
C17728 NAND2X1_LOC_214/B NAND2X1_LOC_74/B 0.11fF
C17729 NAND2X1_LOC_350/A INVX1_LOC_180/Y 0.03fF
C17730 INVX1_LOC_28/A NAND2X1_LOC_656/Y 0.17fF
C17731 INVX1_LOC_1/A NAND2X1_LOC_252/a_36_24# 0.00fF
C17732 NAND2X1_LOC_550/A NAND2X1_LOC_489/a_36_24# 0.00fF
C17733 NAND2X1_LOC_81/B NOR2X1_LOC_652/Y 0.01fF
C17734 INVX1_LOC_229/Y NAND2X1_LOC_560/A 0.01fF
C17735 INVX1_LOC_30/Y NOR2X1_LOC_751/A 0.00fF
C17736 INVX1_LOC_89/A NOR2X1_LOC_356/A 0.07fF
C17737 NAND2X1_LOC_360/B NOR2X1_LOC_78/A 0.07fF
C17738 INVX1_LOC_149/A NOR2X1_LOC_405/A 0.08fF
C17739 INVX1_LOC_33/A NOR2X1_LOC_266/B 0.03fF
C17740 NAND2X1_LOC_222/B NOR2X1_LOC_814/A 0.02fF
C17741 INVX1_LOC_27/A NAND2X1_LOC_74/B 0.47fF
C17742 INVX1_LOC_11/A INVX1_LOC_285/A 0.05fF
C17743 NAND2X1_LOC_363/B NOR2X1_LOC_620/A 0.04fF
C17744 NAND2X1_LOC_392/A INVX1_LOC_286/A 0.00fF
C17745 D_INPUT_1 INVX1_LOC_4/Y 0.03fF
C17746 NOR2X1_LOC_36/A INVX1_LOC_296/A 0.07fF
C17747 NAND2X1_LOC_773/Y NAND2X1_LOC_773/B 0.01fF
C17748 INVX1_LOC_23/Y NOR2X1_LOC_39/a_36_216# 0.02fF
C17749 NAND2X1_LOC_208/a_36_24# INVX1_LOC_42/A 0.00fF
C17750 NOR2X1_LOC_773/Y INVX1_LOC_91/A 0.17fF
C17751 NAND2X1_LOC_35/Y NOR2X1_LOC_496/a_36_216# 0.01fF
C17752 NOR2X1_LOC_196/A INVX1_LOC_9/A 0.11fF
C17753 INVX1_LOC_11/A NOR2X1_LOC_814/A 0.13fF
C17754 NAND2X1_LOC_357/B INVX1_LOC_76/A 0.01fF
C17755 NAND2X1_LOC_391/Y INVX1_LOC_42/A 0.07fF
C17756 NOR2X1_LOC_82/A INVX1_LOC_63/A 0.33fF
C17757 NAND2X1_LOC_303/Y NOR2X1_LOC_11/Y 0.05fF
C17758 NAND2X1_LOC_361/Y INVX1_LOC_117/A 0.16fF
C17759 INVX1_LOC_143/A INVX1_LOC_95/Y 0.10fF
C17760 INVX1_LOC_85/A NOR2X1_LOC_357/Y 0.04fF
C17761 NOR2X1_LOC_433/A NOR2X1_LOC_366/a_36_216# 0.01fF
C17762 NOR2X1_LOC_346/B NOR2X1_LOC_346/Y 0.02fF
C17763 NOR2X1_LOC_318/B INVX1_LOC_1/Y 0.01fF
C17764 NAND2X1_LOC_660/A INVX1_LOC_20/A 0.00fF
C17765 NOR2X1_LOC_773/Y INVX1_LOC_11/Y 0.07fF
C17766 NOR2X1_LOC_718/B NAND2X1_LOC_298/a_36_24# 0.01fF
C17767 INVX1_LOC_89/A NOR2X1_LOC_74/A 0.38fF
C17768 INVX1_LOC_49/A INVX1_LOC_38/A 2.68fF
C17769 INVX1_LOC_24/Y INVX1_LOC_69/A 0.02fF
C17770 NAND2X1_LOC_348/A INPUT_1 0.01fF
C17771 NOR2X1_LOC_860/B NOR2X1_LOC_332/Y 0.03fF
C17772 NOR2X1_LOC_328/Y INVX1_LOC_187/A 0.01fF
C17773 NAND2X1_LOC_392/A INVX1_LOC_95/A 0.34fF
C17774 INVX1_LOC_130/Y NOR2X1_LOC_155/A 0.01fF
C17775 INVX1_LOC_88/A NOR2X1_LOC_755/Y 0.01fF
C17776 INVX1_LOC_93/Y INVX1_LOC_1/Y 0.16fF
C17777 INVX1_LOC_17/A INVX1_LOC_12/A 0.19fF
C17778 NAND2X1_LOC_176/a_36_24# NOR2X1_LOC_74/A 0.08fF
C17779 INVX1_LOC_89/A NOR2X1_LOC_9/Y 0.38fF
C17780 NOR2X1_LOC_172/Y INVX1_LOC_118/A 0.01fF
C17781 NOR2X1_LOC_677/Y INVX1_LOC_23/A 0.09fF
C17782 NOR2X1_LOC_717/B INVX1_LOC_186/A 0.03fF
C17783 INVX1_LOC_104/A NOR2X1_LOC_536/A 0.01fF
C17784 NOR2X1_LOC_666/Y INVX1_LOC_283/A 0.10fF
C17785 NOR2X1_LOC_191/A VDD 0.16fF
C17786 INVX1_LOC_58/A INVX1_LOC_200/Y 0.03fF
C17787 INVX1_LOC_174/A INVX1_LOC_29/A 0.04fF
C17788 INVX1_LOC_35/A NAND2X1_LOC_286/B 0.03fF
C17789 NAND2X1_LOC_850/A INVX1_LOC_100/A 0.20fF
C17790 NOR2X1_LOC_471/Y INVX1_LOC_12/A 0.04fF
C17791 D_INPUT_0 NAND2X1_LOC_490/a_36_24# 0.00fF
C17792 NOR2X1_LOC_750/Y INVX1_LOC_25/A 0.02fF
C17793 INVX1_LOC_2/A NAND2X1_LOC_849/B 0.09fF
C17794 NOR2X1_LOC_67/A NOR2X1_LOC_813/Y 0.39fF
C17795 NOR2X1_LOC_360/Y INVX1_LOC_84/A 0.01fF
C17796 INVX1_LOC_69/Y NOR2X1_LOC_703/A 0.01fF
C17797 INVX1_LOC_269/A INVX1_LOC_47/Y 0.10fF
C17798 NOR2X1_LOC_456/a_36_216# NOR2X1_LOC_334/Y 0.01fF
C17799 INVX1_LOC_2/A INVX1_LOC_38/A 0.18fF
C17800 NOR2X1_LOC_590/A NOR2X1_LOC_89/A 4.34fF
C17801 NOR2X1_LOC_71/Y NOR2X1_LOC_124/A 0.13fF
C17802 NOR2X1_LOC_454/Y NOR2X1_LOC_158/Y 1.69fF
C17803 INVX1_LOC_64/A NOR2X1_LOC_125/Y 0.06fF
C17804 NOR2X1_LOC_717/B NAND2X1_LOC_447/Y 0.00fF
C17805 NOR2X1_LOC_226/A INVX1_LOC_38/A 0.10fF
C17806 NAND2X1_LOC_778/Y NOR2X1_LOC_693/Y 0.10fF
C17807 NAND2X1_LOC_319/A NOR2X1_LOC_314/Y 0.09fF
C17808 INVX1_LOC_311/Y NAND2X1_LOC_677/a_36_24# 0.01fF
C17809 INVX1_LOC_35/A NAND2X1_LOC_860/A 0.07fF
C17810 INVX1_LOC_36/A NOR2X1_LOC_340/A 0.05fF
C17811 INVX1_LOC_104/A NAND2X1_LOC_93/B 0.07fF
C17812 NOR2X1_LOC_433/A INVX1_LOC_285/A 0.07fF
C17813 NAND2X1_LOC_190/Y NOR2X1_LOC_334/Y 0.01fF
C17814 INVX1_LOC_236/Y NOR2X1_LOC_48/B 0.00fF
C17815 INVX1_LOC_64/A NOR2X1_LOC_598/B 0.56fF
C17816 INVX1_LOC_140/A INVX1_LOC_91/A 0.03fF
C17817 NOR2X1_LOC_52/B NOR2X1_LOC_364/A 0.10fF
C17818 INVX1_LOC_35/A NOR2X1_LOC_634/Y 0.41fF
C17819 INVX1_LOC_2/A NOR2X1_LOC_51/A 0.44fF
C17820 NOR2X1_LOC_512/Y INVX1_LOC_49/Y 0.03fF
C17821 NOR2X1_LOC_151/Y INVX1_LOC_186/A 0.07fF
C17822 NOR2X1_LOC_644/A INVX1_LOC_188/Y 0.01fF
C17823 INVX1_LOC_45/A NOR2X1_LOC_114/Y 0.02fF
C17824 NOR2X1_LOC_632/Y INVX1_LOC_281/A 0.16fF
C17825 NAND2X1_LOC_796/B NOR2X1_LOC_654/A 0.30fF
C17826 INVX1_LOC_58/A NOR2X1_LOC_406/A 0.00fF
C17827 NOR2X1_LOC_161/Y INVX1_LOC_38/A 0.01fF
C17828 INVX1_LOC_64/A INVX1_LOC_97/Y 0.01fF
C17829 NOR2X1_LOC_186/Y NAND2X1_LOC_784/A 0.01fF
C17830 NAND2X1_LOC_276/Y INVX1_LOC_27/Y 0.05fF
C17831 NOR2X1_LOC_593/Y NOR2X1_LOC_814/A 0.03fF
C17832 NOR2X1_LOC_188/A NAND2X1_LOC_669/a_36_24# 0.00fF
C17833 INVX1_LOC_64/A NAND2X1_LOC_725/A 0.02fF
C17834 INVX1_LOC_155/Y NAND2X1_LOC_475/Y 0.03fF
C17835 NAND2X1_LOC_348/A INVX1_LOC_154/A 0.00fF
C17836 INVX1_LOC_110/A NOR2X1_LOC_861/Y 0.17fF
C17837 INVX1_LOC_313/A NOR2X1_LOC_137/Y 0.01fF
C17838 NAND2X1_LOC_725/B NAND2X1_LOC_402/B 0.00fF
C17839 INVX1_LOC_14/A INVX1_LOC_183/A 0.03fF
C17840 NAND2X1_LOC_35/Y NAND2X1_LOC_624/B 0.03fF
C17841 NOR2X1_LOC_403/B NAND2X1_LOC_81/B 0.08fF
C17842 D_INPUT_0 NAND2X1_LOC_642/a_36_24# 0.00fF
C17843 NAND2X1_LOC_854/B NOR2X1_LOC_536/A 0.22fF
C17844 NOR2X1_LOC_392/Y INVX1_LOC_306/Y 0.02fF
C17845 INVX1_LOC_200/A NOR2X1_LOC_301/A 0.10fF
C17846 NAND2X1_LOC_392/A INVX1_LOC_54/A 0.03fF
C17847 NOR2X1_LOC_52/B INVX1_LOC_285/A 0.14fF
C17848 INVX1_LOC_223/A INVX1_LOC_32/A 0.03fF
C17849 NOR2X1_LOC_389/A NOR2X1_LOC_334/Y 0.10fF
C17850 INVX1_LOC_27/A INVX1_LOC_259/Y 0.03fF
C17851 NAND2X1_LOC_462/B INVX1_LOC_38/A 0.00fF
C17852 NOR2X1_LOC_91/A NOR2X1_LOC_533/Y 0.03fF
C17853 NAND2X1_LOC_463/B INVX1_LOC_11/Y 0.00fF
C17854 NAND2X1_LOC_784/A NAND2X1_LOC_573/Y 0.05fF
C17855 INVX1_LOC_133/Y NOR2X1_LOC_473/a_36_216# 0.00fF
C17856 NAND2X1_LOC_380/a_36_24# INVX1_LOC_19/A 0.00fF
C17857 NAND2X1_LOC_99/Y NAND2X1_LOC_74/B 0.01fF
C17858 NOR2X1_LOC_52/B NOR2X1_LOC_814/A 0.03fF
C17859 NOR2X1_LOC_188/A NAND2X1_LOC_642/Y 0.05fF
C17860 INVX1_LOC_40/A INVX1_LOC_46/Y 0.03fF
C17861 NAND2X1_LOC_560/A INVX1_LOC_20/A 0.06fF
C17862 NAND2X1_LOC_562/B INVX1_LOC_203/A 0.10fF
C17863 INVX1_LOC_27/A NOR2X1_LOC_660/Y 0.09fF
C17864 NOR2X1_LOC_210/B INVX1_LOC_92/A 0.18fF
C17865 INVX1_LOC_103/A INVX1_LOC_270/A 0.07fF
C17866 NAND2X1_LOC_36/A NAND2X1_LOC_452/Y 0.05fF
C17867 NOR2X1_LOC_473/B NOR2X1_LOC_363/Y 0.02fF
C17868 NOR2X1_LOC_548/B NAND2X1_LOC_642/Y 0.03fF
C17869 INVX1_LOC_71/A NOR2X1_LOC_114/Y 0.12fF
C17870 INVX1_LOC_62/A INVX1_LOC_230/A 0.02fF
C17871 NOR2X1_LOC_303/Y NOR2X1_LOC_631/a_36_216# 0.02fF
C17872 INVX1_LOC_35/A NAND2X1_LOC_473/A 0.13fF
C17873 NOR2X1_LOC_214/a_36_216# INVX1_LOC_109/Y 0.01fF
C17874 D_INPUT_1 NOR2X1_LOC_205/Y 0.02fF
C17875 INVX1_LOC_11/A NAND2X1_LOC_40/a_36_24# 0.00fF
C17876 NOR2X1_LOC_86/A NOR2X1_LOC_235/Y 0.06fF
C17877 NOR2X1_LOC_392/B NAND2X1_LOC_63/Y 0.01fF
C17878 NOR2X1_LOC_664/Y NAND2X1_LOC_74/B 0.04fF
C17879 NAND2X1_LOC_354/B NOR2X1_LOC_89/A 0.03fF
C17880 NOR2X1_LOC_619/A NAND2X1_LOC_85/Y 0.02fF
C17881 INVX1_LOC_292/A INVX1_LOC_270/A 0.01fF
C17882 NOR2X1_LOC_312/Y INVX1_LOC_54/A 0.24fF
C17883 NOR2X1_LOC_249/Y NOR2X1_LOC_343/B 0.09fF
C17884 NOR2X1_LOC_322/Y INVX1_LOC_37/Y 0.01fF
C17885 INVX1_LOC_90/A INVX1_LOC_118/A 5.50fF
C17886 NOR2X1_LOC_276/Y INVX1_LOC_271/A 1.01fF
C17887 INVX1_LOC_201/A INVX1_LOC_20/A 0.01fF
C17888 NAND2X1_LOC_632/a_36_24# INVX1_LOC_260/Y 0.00fF
C17889 NOR2X1_LOC_846/A NAND2X1_LOC_816/a_36_24# 0.00fF
C17890 NOR2X1_LOC_15/Y INVX1_LOC_253/Y 0.42fF
C17891 INVX1_LOC_31/A NOR2X1_LOC_677/Y 0.28fF
C17892 INVX1_LOC_216/A NAND2X1_LOC_82/Y 0.03fF
C17893 INVX1_LOC_78/Y NOR2X1_LOC_35/Y 0.40fF
C17894 NOR2X1_LOC_596/A NOR2X1_LOC_334/Y 0.07fF
C17895 NAND2X1_LOC_553/A NOR2X1_LOC_271/B 0.06fF
C17896 INVX1_LOC_6/A NOR2X1_LOC_137/Y 0.23fF
C17897 NAND2X1_LOC_451/Y NAND2X1_LOC_651/B 0.13fF
C17898 INVX1_LOC_24/A INVX1_LOC_271/Y 0.07fF
C17899 NAND2X1_LOC_21/Y D_INPUT_5 0.30fF
C17900 INVX1_LOC_83/A NOR2X1_LOC_58/a_36_216# 0.14fF
C17901 NOR2X1_LOC_186/Y NAND2X1_LOC_326/A -0.01fF
C17902 INVX1_LOC_286/A NAND2X1_LOC_287/B 0.00fF
C17903 INVX1_LOC_5/A NOR2X1_LOC_739/Y 0.12fF
C17904 INVX1_LOC_88/A NOR2X1_LOC_674/Y 0.15fF
C17905 NOR2X1_LOC_722/Y NOR2X1_LOC_383/B 0.01fF
C17906 NAND2X1_LOC_363/Y NOR2X1_LOC_865/Y 4.02fF
C17907 INVX1_LOC_219/Y INVX1_LOC_3/Y 0.03fF
C17908 INVX1_LOC_89/A NOR2X1_LOC_865/Y 0.07fF
C17909 NOR2X1_LOC_439/B INVX1_LOC_274/A 0.01fF
C17910 INVX1_LOC_136/A INVX1_LOC_271/A 0.01fF
C17911 INVX1_LOC_230/Y INVX1_LOC_138/Y 0.93fF
C17912 INVX1_LOC_85/A INVX1_LOC_32/A 0.03fF
C17913 INVX1_LOC_58/A INVX1_LOC_250/A 0.01fF
C17914 INVX1_LOC_83/A NOR2X1_LOC_673/A 0.07fF
C17915 INVX1_LOC_89/A NOR2X1_LOC_243/B 0.16fF
C17916 INVX1_LOC_75/A INVX1_LOC_274/A 0.06fF
C17917 NOR2X1_LOC_34/A INVX1_LOC_17/A 0.10fF
C17918 NOR2X1_LOC_488/Y NOR2X1_LOC_89/A 0.03fF
C17919 INVX1_LOC_137/A NAND2X1_LOC_74/B 0.00fF
C17920 NOR2X1_LOC_639/B INVX1_LOC_30/A 0.08fF
C17921 INVX1_LOC_95/A NAND2X1_LOC_287/B 0.01fF
C17922 INVX1_LOC_89/A NOR2X1_LOC_461/a_36_216# 0.02fF
C17923 NOR2X1_LOC_589/A INVX1_LOC_29/A 0.22fF
C17924 INVX1_LOC_160/Y NOR2X1_LOC_777/B 0.03fF
C17925 NAND2X1_LOC_508/A NOR2X1_LOC_243/B 0.03fF
C17926 NAND2X1_LOC_451/Y INVX1_LOC_15/A 0.07fF
C17927 NOR2X1_LOC_631/B INVX1_LOC_37/A 0.07fF
C17928 INVX1_LOC_27/A NOR2X1_LOC_276/Y 0.03fF
C17929 INPUT_5 INPUT_7 0.09fF
C17930 NAND2X1_LOC_351/a_36_24# NAND2X1_LOC_351/A 0.00fF
C17931 INVX1_LOC_234/A NAND2X1_LOC_74/B 0.07fF
C17932 NAND2X1_LOC_794/B INVX1_LOC_141/Y 0.01fF
C17933 NOR2X1_LOC_772/B INVX1_LOC_72/A 0.10fF
C17934 NOR2X1_LOC_34/A NAND2X1_LOC_555/Y -0.01fF
C17935 NOR2X1_LOC_381/Y NOR2X1_LOC_817/Y 0.08fF
C17936 INVX1_LOC_216/Y INVX1_LOC_269/A 0.03fF
C17937 NOR2X1_LOC_689/A INVX1_LOC_34/A 0.01fF
C17938 NOR2X1_LOC_577/Y INVX1_LOC_57/A 0.08fF
C17939 INVX1_LOC_227/A NOR2X1_LOC_89/A 0.07fF
C17940 NOR2X1_LOC_456/Y NOR2X1_LOC_303/Y 0.07fF
C17941 INVX1_LOC_136/A NAND2X1_LOC_214/B 0.01fF
C17942 NOR2X1_LOC_609/a_36_216# INVX1_LOC_53/A 0.01fF
C17943 INVX1_LOC_303/A NAND2X1_LOC_275/a_36_24# 0.00fF
C17944 INVX1_LOC_34/A NOR2X1_LOC_383/B 0.03fF
C17945 INVX1_LOC_17/A INVX1_LOC_200/A 0.03fF
C17946 NAND2X1_LOC_9/Y NOR2X1_LOC_403/a_36_216# 0.00fF
C17947 INVX1_LOC_48/Y INVX1_LOC_39/Y 0.01fF
C17948 INVX1_LOC_13/Y INVX1_LOC_72/A 0.01fF
C17949 INVX1_LOC_58/A NAND2X1_LOC_361/Y 0.14fF
C17950 NOR2X1_LOC_837/Y NAND2X1_LOC_363/B 0.01fF
C17951 NOR2X1_LOC_102/a_36_216# INVX1_LOC_59/Y 0.00fF
C17952 NOR2X1_LOC_6/B NOR2X1_LOC_39/Y 0.17fF
C17953 NOR2X1_LOC_733/Y INVX1_LOC_179/A 0.01fF
C17954 NOR2X1_LOC_19/B INVX1_LOC_293/Y 0.01fF
C17955 NOR2X1_LOC_220/A NOR2X1_LOC_334/Y 0.10fF
C17956 INVX1_LOC_90/A NAND2X1_LOC_63/Y 0.27fF
C17957 NAND2X1_LOC_662/Y INVX1_LOC_32/A 0.01fF
C17958 NAND2X1_LOC_803/B INVX1_LOC_11/A 0.00fF
C17959 INVX1_LOC_34/A NAND2X1_LOC_738/B 0.03fF
C17960 INVX1_LOC_136/A INVX1_LOC_27/A 0.12fF
C17961 INVX1_LOC_136/A NOR2X1_LOC_824/A 0.07fF
C17962 NOR2X1_LOC_643/A NAND2X1_LOC_555/Y 0.05fF
C17963 NAND2X1_LOC_35/Y NOR2X1_LOC_617/Y 0.05fF
C17964 INVX1_LOC_224/A NOR2X1_LOC_590/A 0.03fF
C17965 INVX1_LOC_86/Y NAND2X1_LOC_425/Y 0.08fF
C17966 NOR2X1_LOC_456/Y NOR2X1_LOC_254/Y 0.07fF
C17967 INVX1_LOC_225/A NAND2X1_LOC_784/A -0.02fF
C17968 NAND2X1_LOC_464/a_36_24# NAND2X1_LOC_99/A 0.00fF
C17969 NAND2X1_LOC_303/Y NOR2X1_LOC_599/A 0.03fF
C17970 INVX1_LOC_88/A NOR2X1_LOC_361/a_36_216# 0.00fF
C17971 INVX1_LOC_11/A NOR2X1_LOC_590/A 0.81fF
C17972 INVX1_LOC_224/A INVX1_LOC_22/Y 0.01fF
C17973 NOR2X1_LOC_458/Y NOR2X1_LOC_678/A 0.01fF
C17974 INVX1_LOC_153/Y NOR2X1_LOC_678/A 0.03fF
C17975 NOR2X1_LOC_19/B NAND2X1_LOC_74/B 0.02fF
C17976 NAND2X1_LOC_715/a_36_24# INVX1_LOC_32/A 0.00fF
C17977 INVX1_LOC_99/Y NOR2X1_LOC_550/B 0.01fF
C17978 INVX1_LOC_59/Y NOR2X1_LOC_656/Y 0.00fF
C17979 INVX1_LOC_1/Y INVX1_LOC_87/A 2.81fF
C17980 NAND2X1_LOC_634/a_36_24# NAND2X1_LOC_634/Y 0.02fF
C17981 INPUT_2 INPUT_3 0.33fF
C17982 INVX1_LOC_11/A INVX1_LOC_22/Y 0.01fF
C17983 INVX1_LOC_89/Y NOR2X1_LOC_124/A 0.01fF
C17984 INVX1_LOC_55/Y INVX1_LOC_290/Y 0.07fF
C17985 NOR2X1_LOC_171/Y INVX1_LOC_12/A 0.04fF
C17986 INVX1_LOC_35/A NOR2X1_LOC_516/Y 0.03fF
C17987 INVX1_LOC_36/A INVX1_LOC_103/A 0.10fF
C17988 NAND2X1_LOC_218/B INVX1_LOC_252/A 0.04fF
C17989 NAND2X1_LOC_363/B NOR2X1_LOC_720/B 0.04fF
C17990 INVX1_LOC_88/A INVX1_LOC_72/A 0.03fF
C17991 NOR2X1_LOC_596/Y NOR2X1_LOC_644/B 0.12fF
C17992 NOR2X1_LOC_78/A NAND2X1_LOC_572/B 0.79fF
C17993 INVX1_LOC_64/A NAND2X1_LOC_308/Y 0.03fF
C17994 NAND2X1_LOC_276/Y INVX1_LOC_5/A 0.00fF
C17995 NOR2X1_LOC_647/A NOR2X1_LOC_516/B 0.04fF
C17996 INVX1_LOC_90/A INVX1_LOC_257/A 0.02fF
C17997 NOR2X1_LOC_91/A INVX1_LOC_56/Y 0.03fF
C17998 INVX1_LOC_75/A NOR2X1_LOC_33/B 0.02fF
C17999 NOR2X1_LOC_218/A INVX1_LOC_30/A 0.00fF
C18000 INVX1_LOC_10/A INVX1_LOC_94/Y 0.06fF
C18001 INVX1_LOC_14/A INVX1_LOC_72/Y 0.04fF
C18002 NOR2X1_LOC_346/B INVX1_LOC_57/A 0.02fF
C18003 NOR2X1_LOC_816/Y NAND2X1_LOC_848/A 0.13fF
C18004 NAND2X1_LOC_724/Y NAND2X1_LOC_853/Y 3.89fF
C18005 NOR2X1_LOC_612/Y INVX1_LOC_46/A 0.04fF
C18006 NAND2X1_LOC_434/a_36_24# NAND2X1_LOC_798/B 0.00fF
C18007 NOR2X1_LOC_391/A INVX1_LOC_23/Y 0.07fF
C18008 NOR2X1_LOC_415/A NOR2X1_LOC_415/Y 0.00fF
C18009 NAND2X1_LOC_564/B NAND2X1_LOC_439/a_36_24# 0.00fF
C18010 NOR2X1_LOC_15/Y NAND2X1_LOC_740/A 0.02fF
C18011 INVX1_LOC_22/A INVX1_LOC_57/A 1.44fF
C18012 NOR2X1_LOC_160/B INVX1_LOC_205/A 0.00fF
C18013 INVX1_LOC_56/Y INVX1_LOC_23/A 0.20fF
C18014 INVX1_LOC_103/A NOR2X1_LOC_208/Y 0.27fF
C18015 NAND2X1_LOC_562/a_36_24# NAND2X1_LOC_577/A 0.01fF
C18016 INVX1_LOC_204/A NOR2X1_LOC_589/A 0.05fF
C18017 INVX1_LOC_39/A NOR2X1_LOC_392/B 0.01fF
C18018 NOR2X1_LOC_567/B INVX1_LOC_15/A 0.12fF
C18019 NAND2X1_LOC_599/a_36_24# NOR2X1_LOC_544/A 0.00fF
C18020 INVX1_LOC_305/Y NOR2X1_LOC_634/Y 0.16fF
C18021 INVX1_LOC_38/A INVX1_LOC_118/A 0.30fF
C18022 NAND2X1_LOC_848/A NOR2X1_LOC_177/a_36_216# 0.13fF
C18023 NAND2X1_LOC_773/Y NOR2X1_LOC_557/Y 0.10fF
C18024 INVX1_LOC_5/A NOR2X1_LOC_352/Y 0.01fF
C18025 INVX1_LOC_309/A INVX1_LOC_42/A 0.03fF
C18026 INVX1_LOC_161/Y NOR2X1_LOC_106/Y 0.05fF
C18027 INVX1_LOC_16/A NOR2X1_LOC_717/A 0.10fF
C18028 INVX1_LOC_59/Y INVX1_LOC_63/A 0.03fF
C18029 INVX1_LOC_89/A NAND2X1_LOC_425/a_36_24# 0.00fF
C18030 INVX1_LOC_13/Y NOR2X1_LOC_537/Y 0.32fF
C18031 INVX1_LOC_69/Y NOR2X1_LOC_169/a_36_216# 0.01fF
C18032 NAND2X1_LOC_374/a_36_24# NAND2X1_LOC_550/A 0.00fF
C18033 INVX1_LOC_13/Y NAND2X1_LOC_338/B 2.20fF
C18034 NOR2X1_LOC_99/B NOR2X1_LOC_844/a_36_216# 0.01fF
C18035 NAND2X1_LOC_803/B NOR2X1_LOC_433/A 0.03fF
C18036 INVX1_LOC_176/A INVX1_LOC_63/A 1.97fF
C18037 NAND2X1_LOC_114/B NOR2X1_LOC_350/A 0.35fF
C18038 NAND2X1_LOC_30/Y INVX1_LOC_33/A 0.05fF
C18039 NAND2X1_LOC_93/B NOR2X1_LOC_119/a_36_216# 0.00fF
C18040 INVX1_LOC_178/A NAND2X1_LOC_374/Y 0.10fF
C18041 INVX1_LOC_91/A INVX1_LOC_42/A 1.25fF
C18042 NOR2X1_LOC_483/B INVX1_LOC_49/A 0.09fF
C18043 INVX1_LOC_291/A NAND2X1_LOC_760/a_36_24# 0.01fF
C18044 INVX1_LOC_25/Y INVX1_LOC_306/Y 0.06fF
C18045 INVX1_LOC_79/A INVX1_LOC_78/A 0.01fF
C18046 NOR2X1_LOC_590/A NOR2X1_LOC_433/A 0.10fF
C18047 INVX1_LOC_292/A NOR2X1_LOC_804/B -0.00fF
C18048 INVX1_LOC_201/A INVX1_LOC_4/A 0.04fF
C18049 NAND2X1_LOC_773/Y INVX1_LOC_143/A 0.10fF
C18050 NOR2X1_LOC_590/A NOR2X1_LOC_593/Y 0.03fF
C18051 INVX1_LOC_20/A INVX1_LOC_29/A 1.19fF
C18052 INVX1_LOC_11/Y INVX1_LOC_42/A 0.03fF
C18053 INVX1_LOC_225/A NAND2X1_LOC_807/A 0.01fF
C18054 NOR2X1_LOC_15/Y NOR2X1_LOC_190/a_36_216# 0.00fF
C18055 INVX1_LOC_256/A INVX1_LOC_104/A 1.02fF
C18056 NOR2X1_LOC_68/A NAND2X1_LOC_656/A 0.05fF
C18057 NAND2X1_LOC_803/B NOR2X1_LOC_52/B 0.05fF
C18058 NOR2X1_LOC_269/Y INVX1_LOC_15/A 0.05fF
C18059 INVX1_LOC_89/A NOR2X1_LOC_342/A 0.34fF
C18060 NAND2X1_LOC_149/Y NOR2X1_LOC_146/Y 0.05fF
C18061 NOR2X1_LOC_361/B NOR2X1_LOC_191/A 0.03fF
C18062 NOR2X1_LOC_432/Y NAND2X1_LOC_53/Y 0.02fF
C18063 INVX1_LOC_35/A INVX1_LOC_85/Y 0.03fF
C18064 INVX1_LOC_36/A INVX1_LOC_67/A 0.18fF
C18065 INVX1_LOC_30/A INVX1_LOC_155/Y 0.03fF
C18066 INVX1_LOC_17/A INVX1_LOC_214/Y 0.05fF
C18067 NAND2X1_LOC_287/B NAND2X1_LOC_807/B 0.02fF
C18068 NOR2X1_LOC_590/A NOR2X1_LOC_52/B 0.06fF
C18069 NAND2X1_LOC_386/a_36_24# INVX1_LOC_49/A 0.01fF
C18070 NAND2X1_LOC_840/Y NOR2X1_LOC_654/A 0.01fF
C18071 NOR2X1_LOC_675/a_36_216# INVX1_LOC_285/A 0.00fF
C18072 NOR2X1_LOC_479/B INVX1_LOC_269/A 0.01fF
C18073 INVX1_LOC_30/A NOR2X1_LOC_364/Y 0.00fF
C18074 INPUT_0 NOR2X1_LOC_383/B 0.51fF
C18075 INVX1_LOC_255/Y NOR2X1_LOC_15/Y 0.07fF
C18076 INVX1_LOC_78/A INVX1_LOC_91/A 0.25fF
C18077 NOR2X1_LOC_290/a_36_216# INVX1_LOC_42/A 0.01fF
C18078 NOR2X1_LOC_19/B NOR2X1_LOC_660/Y 0.08fF
C18079 INVX1_LOC_102/A NAND2X1_LOC_804/Y 0.03fF
C18080 NAND2X1_LOC_738/B INPUT_0 0.03fF
C18081 INVX1_LOC_11/A NOR2X1_LOC_82/Y 0.01fF
C18082 NAND2X1_LOC_63/Y INVX1_LOC_38/A 0.03fF
C18083 NOR2X1_LOC_637/B NOR2X1_LOC_637/Y 0.07fF
C18084 NOR2X1_LOC_717/Y INVX1_LOC_266/Y 0.00fF
C18085 NOR2X1_LOC_65/B NOR2X1_LOC_114/A 0.16fF
C18086 INVX1_LOC_64/A NAND2X1_LOC_560/A 0.03fF
C18087 INVX1_LOC_93/Y INVX1_LOC_87/A 0.08fF
C18088 INVX1_LOC_59/A NOR2X1_LOC_130/A 1.41fF
C18089 NOR2X1_LOC_391/Y NAND2X1_LOC_215/A 0.03fF
C18090 INVX1_LOC_39/A INVX1_LOC_90/A 0.00fF
C18091 NAND2X1_LOC_348/A INVX1_LOC_138/A 0.01fF
C18092 INVX1_LOC_288/A INVX1_LOC_91/A 0.00fF
C18093 INVX1_LOC_223/Y NOR2X1_LOC_356/A 0.09fF
C18094 NOR2X1_LOC_257/Y INVX1_LOC_92/A 0.03fF
C18095 NOR2X1_LOC_65/B INVX1_LOC_91/A 0.16fF
C18096 NOR2X1_LOC_20/Y NAND2X1_LOC_462/B 0.01fF
C18097 NOR2X1_LOC_523/B NOR2X1_LOC_844/A 0.01fF
C18098 NAND2X1_LOC_338/B NOR2X1_LOC_500/B 0.12fF
C18099 NAND2X1_LOC_725/A INVX1_LOC_282/A 0.10fF
C18100 NOR2X1_LOC_68/A NOR2X1_LOC_423/Y 0.09fF
C18101 NOR2X1_LOC_15/Y NOR2X1_LOC_71/Y 0.68fF
C18102 INVX1_LOC_33/A INVX1_LOC_49/A 0.26fF
C18103 NOR2X1_LOC_791/Y NAND2X1_LOC_842/a_36_24# 0.01fF
C18104 INVX1_LOC_285/Y NOR2X1_LOC_678/A 0.03fF
C18105 NOR2X1_LOC_815/Y NOR2X1_LOC_172/Y 0.08fF
C18106 NOR2X1_LOC_815/a_36_216# NAND2X1_LOC_175/B 0.01fF
C18107 INVX1_LOC_75/A INVX1_LOC_306/Y 0.07fF
C18108 INVX1_LOC_17/A NAND2X1_LOC_808/A 0.68fF
C18109 NOR2X1_LOC_433/A NAND2X1_LOC_354/B 0.02fF
C18110 INVX1_LOC_34/A NAND2X1_LOC_632/B 0.02fF
C18111 NOR2X1_LOC_550/B NOR2X1_LOC_254/Y 0.01fF
C18112 INVX1_LOC_11/A NOR2X1_LOC_763/Y 0.08fF
C18113 NOR2X1_LOC_409/B INVX1_LOC_46/A 0.03fF
C18114 NOR2X1_LOC_658/Y INVX1_LOC_16/A 0.07fF
C18115 INVX1_LOC_37/A NAND2X1_LOC_72/B 0.03fF
C18116 NOR2X1_LOC_324/A NOR2X1_LOC_383/B 0.04fF
C18117 NOR2X1_LOC_222/Y NOR2X1_LOC_68/A 0.07fF
C18118 NOR2X1_LOC_99/Y INVX1_LOC_284/A 0.01fF
C18119 INVX1_LOC_39/A NAND2X1_LOC_348/A 0.01fF
C18120 INVX1_LOC_88/A INVX1_LOC_313/Y 0.01fF
C18121 NOR2X1_LOC_216/B NAND2X1_LOC_74/B 0.01fF
C18122 NOR2X1_LOC_75/Y NOR2X1_LOC_207/a_36_216# 0.00fF
C18123 INVX1_LOC_179/A INVX1_LOC_99/A 0.00fF
C18124 NOR2X1_LOC_516/B INVX1_LOC_205/A 0.01fF
C18125 NOR2X1_LOC_727/B NOR2X1_LOC_35/Y 0.00fF
C18126 NOR2X1_LOC_229/Y INVX1_LOC_18/A 0.02fF
C18127 NOR2X1_LOC_831/Y NOR2X1_LOC_841/A 0.05fF
C18128 INVX1_LOC_245/Y INVX1_LOC_89/A 0.01fF
C18129 INVX1_LOC_90/A NAND2X1_LOC_352/a_36_24# 0.00fF
C18130 NAND2X1_LOC_170/A NOR2X1_LOC_518/a_36_216# 0.00fF
C18131 NOR2X1_LOC_252/Y INVX1_LOC_217/A 0.16fF
C18132 INVX1_LOC_303/A NOR2X1_LOC_537/Y 0.07fF
C18133 NOR2X1_LOC_524/Y INVX1_LOC_10/A 0.09fF
C18134 INVX1_LOC_268/A INVX1_LOC_159/A 0.04fF
C18135 INVX1_LOC_50/A NOR2X1_LOC_314/Y 0.02fF
C18136 INVX1_LOC_150/Y NAND2X1_LOC_842/B 0.01fF
C18137 INVX1_LOC_2/A INVX1_LOC_33/A 0.10fF
C18138 NOR2X1_LOC_312/Y NOR2X1_LOC_441/Y 0.08fF
C18139 NOR2X1_LOC_220/a_36_216# INVX1_LOC_22/A 0.00fF
C18140 NOR2X1_LOC_68/A INVX1_LOC_220/Y 0.01fF
C18141 NAND2X1_LOC_483/Y NOR2X1_LOC_482/Y 0.06fF
C18142 INVX1_LOC_136/A INVX1_LOC_234/A 0.01fF
C18143 NAND2X1_LOC_477/Y NAND2X1_LOC_74/B 0.43fF
C18144 NOR2X1_LOC_845/A NOR2X1_LOC_849/A 0.01fF
C18145 NOR2X1_LOC_226/A INVX1_LOC_33/A 0.07fF
C18146 INVX1_LOC_85/A NAND2X1_LOC_147/a_36_24# 0.02fF
C18147 NOR2X1_LOC_160/B INVX1_LOC_148/A 0.00fF
C18148 INVX1_LOC_38/A NOR2X1_LOC_631/Y 0.15fF
C18149 NOR2X1_LOC_509/a_36_216# NOR2X1_LOC_814/A 0.01fF
C18150 INVX1_LOC_45/A NAND2X1_LOC_189/a_36_24# 0.00fF
C18151 INVX1_LOC_50/A INVX1_LOC_117/A 0.01fF
C18152 INVX1_LOC_279/A INVX1_LOC_24/A 0.07fF
C18153 INVX1_LOC_209/Y NAND2X1_LOC_863/B 0.00fF
C18154 INVX1_LOC_13/A INVX1_LOC_77/A 0.17fF
C18155 INVX1_LOC_21/A NOR2X1_LOC_746/Y 0.26fF
C18156 NOR2X1_LOC_218/Y INVX1_LOC_33/A 0.02fF
C18157 INVX1_LOC_203/A INVX1_LOC_42/A 0.10fF
C18158 NOR2X1_LOC_220/A NOR2X1_LOC_718/B 0.24fF
C18159 INVX1_LOC_60/A INVX1_LOC_40/A 0.01fF
C18160 INVX1_LOC_271/Y NOR2X1_LOC_197/B 0.10fF
C18161 NOR2X1_LOC_128/A INVX1_LOC_29/A 0.01fF
C18162 INVX1_LOC_136/A NOR2X1_LOC_772/A 0.01fF
C18163 INVX1_LOC_90/A INVX1_LOC_61/A 0.15fF
C18164 NAND2X1_LOC_547/a_36_24# NAND2X1_LOC_808/A 0.00fF
C18165 NOR2X1_LOC_488/Y NOR2X1_LOC_52/B 0.94fF
C18166 NOR2X1_LOC_77/a_36_216# NOR2X1_LOC_89/A 0.03fF
C18167 NOR2X1_LOC_808/A NOR2X1_LOC_811/B 0.02fF
C18168 INVX1_LOC_136/A NOR2X1_LOC_19/B 0.08fF
C18169 NAND2X1_LOC_326/A NAND2X1_LOC_642/Y 0.06fF
C18170 NOR2X1_LOC_52/B NOR2X1_LOC_82/Y 0.03fF
C18171 INVX1_LOC_227/A NOR2X1_LOC_593/Y 0.07fF
C18172 NOR2X1_LOC_75/Y NOR2X1_LOC_737/a_36_216# 0.00fF
C18173 NOR2X1_LOC_717/Y INVX1_LOC_42/Y 0.29fF
C18174 NAND2X1_LOC_326/A NAND2X1_LOC_643/a_36_24# 0.01fF
C18175 INVX1_LOC_2/A INVX1_LOC_40/A 0.12fF
C18176 NOR2X1_LOC_68/A NOR2X1_LOC_329/B 0.07fF
C18177 INVX1_LOC_102/A NOR2X1_LOC_519/a_36_216# 0.01fF
C18178 NOR2X1_LOC_38/B NAND2X1_LOC_206/Y 0.13fF
C18179 NOR2X1_LOC_818/Y INVX1_LOC_40/A 0.92fF
C18180 INVX1_LOC_21/A INVX1_LOC_36/Y 0.03fF
C18181 NOR2X1_LOC_226/A NAND2X1_LOC_798/A 0.10fF
C18182 INVX1_LOC_77/A NOR2X1_LOC_174/B 0.09fF
C18183 NAND2X1_LOC_276/Y NOR2X1_LOC_332/A 0.08fF
C18184 INVX1_LOC_255/Y NAND2X1_LOC_141/A 0.01fF
C18185 NAND2X1_LOC_428/a_36_24# INVX1_LOC_296/A 0.02fF
C18186 INVX1_LOC_299/A NOR2X1_LOC_799/B 0.02fF
C18187 NOR2X1_LOC_13/Y INVX1_LOC_28/A 0.01fF
C18188 INVX1_LOC_57/Y INPUT_0 0.10fF
C18189 NOR2X1_LOC_38/B NAND2X1_LOC_773/B 0.26fF
C18190 NOR2X1_LOC_321/Y NAND2X1_LOC_211/Y 0.01fF
C18191 NOR2X1_LOC_82/A INVX1_LOC_93/Y 0.09fF
C18192 NOR2X1_LOC_538/B NOR2X1_LOC_799/B 0.11fF
C18193 NOR2X1_LOC_815/Y INVX1_LOC_90/A 0.05fF
C18194 INVX1_LOC_78/A INVX1_LOC_203/A 0.01fF
C18195 INVX1_LOC_33/A INPUT_1 0.10fF
C18196 INVX1_LOC_89/A NOR2X1_LOC_121/Y 0.00fF
C18197 INVX1_LOC_29/A INVX1_LOC_4/A 5.18fF
C18198 INVX1_LOC_234/A NAND2X1_LOC_859/a_36_24# 0.00fF
C18199 INVX1_LOC_26/A INVX1_LOC_84/A 0.23fF
C18200 NOR2X1_LOC_624/A INVX1_LOC_90/A 0.47fF
C18201 NOR2X1_LOC_831/B INVX1_LOC_23/A 0.61fF
C18202 NOR2X1_LOC_220/A NOR2X1_LOC_569/Y 0.10fF
C18203 NOR2X1_LOC_644/Y NOR2X1_LOC_717/B 0.00fF
C18204 INVX1_LOC_32/A INVX1_LOC_290/Y 0.07fF
C18205 NAND2X1_LOC_63/Y NAND2X1_LOC_223/A 0.02fF
C18206 INVX1_LOC_128/Y INVX1_LOC_109/A 0.35fF
C18207 NAND2X1_LOC_543/Y NAND2X1_LOC_564/B 0.00fF
C18208 INVX1_LOC_64/A INVX1_LOC_152/A 0.22fF
C18209 NAND2X1_LOC_99/A NAND2X1_LOC_768/Y 0.01fF
C18210 INVX1_LOC_45/A NAND2X1_LOC_655/A 0.07fF
C18211 NOR2X1_LOC_360/Y INVX1_LOC_123/A 0.21fF
C18212 INVX1_LOC_205/A INVX1_LOC_315/Y 0.22fF
C18213 NOR2X1_LOC_713/B INVX1_LOC_86/A 0.04fF
C18214 NOR2X1_LOC_216/B NOR2X1_LOC_660/Y 0.00fF
C18215 INVX1_LOC_90/A NOR2X1_LOC_93/a_36_216# 0.00fF
C18216 NOR2X1_LOC_92/Y NOR2X1_LOC_536/A 0.13fF
C18217 NOR2X1_LOC_798/A NOR2X1_LOC_612/Y 0.02fF
C18218 NOR2X1_LOC_391/A INVX1_LOC_232/A 0.09fF
C18219 NAND2X1_LOC_662/Y GATE_662 0.03fF
C18220 NOR2X1_LOC_569/Y NOR2X1_LOC_548/Y 0.00fF
C18221 NOR2X1_LOC_318/A NAND2X1_LOC_81/B 0.01fF
C18222 NOR2X1_LOC_464/a_36_216# NOR2X1_LOC_151/Y 0.00fF
C18223 INVX1_LOC_305/A INVX1_LOC_65/A 0.18fF
C18224 INVX1_LOC_178/A NAND2X1_LOC_624/a_36_24# 0.00fF
C18225 INVX1_LOC_101/Y NOR2X1_LOC_331/B 0.01fF
C18226 INVX1_LOC_188/A VDD 0.12fF
C18227 NAND2X1_LOC_84/Y INVX1_LOC_125/Y 0.27fF
C18228 NAND2X1_LOC_568/A NOR2X1_LOC_536/A 0.01fF
C18229 NOR2X1_LOC_383/Y NOR2X1_LOC_391/A 0.03fF
C18230 INVX1_LOC_290/A NAND2X1_LOC_656/Y 0.01fF
C18231 INVX1_LOC_41/A INVX1_LOC_126/Y 0.01fF
C18232 NOR2X1_LOC_297/A NOR2X1_LOC_38/B 0.01fF
C18233 NOR2X1_LOC_441/Y NAND2X1_LOC_287/B 0.00fF
C18234 NAND2X1_LOC_721/B INVX1_LOC_20/A 0.00fF
C18235 INVX1_LOC_40/A INPUT_1 0.02fF
C18236 INVX1_LOC_225/A NOR2X1_LOC_527/Y 0.00fF
C18237 INVX1_LOC_12/A INVX1_LOC_296/A 0.03fF
C18238 NOR2X1_LOC_152/Y INVX1_LOC_91/A 0.09fF
C18239 NOR2X1_LOC_564/Y INVX1_LOC_179/Y 0.02fF
C18240 NAND2X1_LOC_288/B NAND2X1_LOC_288/a_36_24# 0.00fF
C18241 NOR2X1_LOC_419/Y NOR2X1_LOC_78/A 0.02fF
C18242 INVX1_LOC_232/Y NOR2X1_LOC_381/a_36_216# 0.00fF
C18243 NOR2X1_LOC_716/B INVX1_LOC_98/A 0.10fF
C18244 INVX1_LOC_35/A NAND2X1_LOC_782/B 0.09fF
C18245 INVX1_LOC_36/A NOR2X1_LOC_137/Y 0.06fF
C18246 NOR2X1_LOC_15/Y NAND2X1_LOC_243/Y 0.06fF
C18247 NOR2X1_LOC_191/B INVX1_LOC_95/Y 0.68fF
C18248 NOR2X1_LOC_195/A INVX1_LOC_9/A 0.01fF
C18249 INVX1_LOC_69/Y INVX1_LOC_104/A 0.07fF
C18250 INVX1_LOC_21/Y INVX1_LOC_273/A 0.07fF
C18251 NOR2X1_LOC_716/B NOR2X1_LOC_78/A 0.99fF
C18252 NOR2X1_LOC_426/Y INVX1_LOC_77/Y 0.05fF
C18253 NOR2X1_LOC_570/B INVX1_LOC_96/A 0.02fF
C18254 NOR2X1_LOC_788/a_36_216# INVX1_LOC_104/A 0.00fF
C18255 NOR2X1_LOC_152/Y INVX1_LOC_11/Y 0.03fF
C18256 INVX1_LOC_71/A NAND2X1_LOC_468/B 0.03fF
C18257 INVX1_LOC_7/Y INVX1_LOC_3/A 0.01fF
C18258 INVX1_LOC_298/Y INVX1_LOC_4/A 0.10fF
C18259 INVX1_LOC_90/A INPUT_5 0.01fF
C18260 INVX1_LOC_134/A NOR2X1_LOC_856/A 0.23fF
C18261 NAND2X1_LOC_82/a_36_24# NOR2X1_LOC_660/Y 0.01fF
C18262 INVX1_LOC_103/A NOR2X1_LOC_435/A 0.01fF
C18263 INVX1_LOC_49/A NOR2X1_LOC_486/Y 0.03fF
C18264 INVX1_LOC_135/A INVX1_LOC_148/Y 0.08fF
C18265 INVX1_LOC_299/A NOR2X1_LOC_445/B 0.02fF
C18266 INVX1_LOC_17/A INVX1_LOC_92/A 0.10fF
C18267 INVX1_LOC_64/A INVX1_LOC_29/A 0.38fF
C18268 D_INPUT_0 INVX1_LOC_89/A 4.24fF
C18269 INVX1_LOC_5/A INVX1_LOC_125/A 0.22fF
C18270 INVX1_LOC_83/A INVX1_LOC_20/Y 0.02fF
C18271 NOR2X1_LOC_238/Y VDD 0.56fF
C18272 NOR2X1_LOC_355/A NOR2X1_LOC_473/B 0.13fF
C18273 INVX1_LOC_25/Y NOR2X1_LOC_74/A 0.11fF
C18274 INVX1_LOC_77/A NOR2X1_LOC_357/Y 0.07fF
C18275 INVX1_LOC_218/A INVX1_LOC_51/Y 0.03fF
C18276 NOR2X1_LOC_471/Y INVX1_LOC_92/A 0.19fF
C18277 INVX1_LOC_181/Y NOR2X1_LOC_558/a_36_216# 0.00fF
C18278 NAND2X1_LOC_170/A INPUT_0 0.04fF
C18279 INVX1_LOC_93/A NAND2X1_LOC_74/B 0.07fF
C18280 NAND2X1_LOC_45/Y NOR2X1_LOC_702/Y 0.04fF
C18281 NOR2X1_LOC_596/A NAND2X1_LOC_472/Y 0.38fF
C18282 INVX1_LOC_276/A NOR2X1_LOC_45/B 0.08fF
C18283 INVX1_LOC_25/Y NOR2X1_LOC_9/Y 0.08fF
C18284 INVX1_LOC_6/A INVX1_LOC_56/Y 0.12fF
C18285 NOR2X1_LOC_67/A NOR2X1_LOC_45/B 0.07fF
C18286 INVX1_LOC_8/A INVX1_LOC_20/A 0.11fF
C18287 NAND2X1_LOC_859/B INVX1_LOC_309/A 0.33fF
C18288 NAND2X1_LOC_501/a_36_24# INVX1_LOC_118/A 0.00fF
C18289 NAND2X1_LOC_358/Y NOR2X1_LOC_97/A 0.15fF
C18290 NOR2X1_LOC_543/A NOR2X1_LOC_188/A 0.04fF
C18291 NOR2X1_LOC_419/Y NOR2X1_LOC_98/a_36_216# 0.00fF
C18292 NAND2X1_LOC_837/Y NOR2X1_LOC_536/A 0.13fF
C18293 INVX1_LOC_310/Y INVX1_LOC_37/A 0.07fF
C18294 INVX1_LOC_103/A INVX1_LOC_63/A 0.02fF
C18295 NAND2X1_LOC_360/B NAND2X1_LOC_642/Y 0.44fF
C18296 NOR2X1_LOC_780/B INVX1_LOC_301/A 0.32fF
C18297 NAND2X1_LOC_364/A NOR2X1_LOC_641/Y 0.04fF
C18298 INVX1_LOC_21/A INVX1_LOC_102/A 0.07fF
C18299 INVX1_LOC_1/A NAND2X1_LOC_82/Y 0.06fF
C18300 INVX1_LOC_14/A INVX1_LOC_19/A 0.11fF
C18301 NOR2X1_LOC_52/B NAND2X1_LOC_650/B 0.07fF
C18302 NOR2X1_LOC_97/A NOR2X1_LOC_99/B 0.10fF
C18303 D_INPUT_4 NOR2X1_LOC_163/A 0.00fF
C18304 INVX1_LOC_142/A NOR2X1_LOC_155/A 0.02fF
C18305 NOR2X1_LOC_722/Y INVX1_LOC_179/A 0.01fF
C18306 INVX1_LOC_136/A NOR2X1_LOC_216/B 0.01fF
C18307 INVX1_LOC_35/A NAND2X1_LOC_454/Y 0.07fF
C18308 NOR2X1_LOC_843/B INVX1_LOC_57/A 0.07fF
C18309 INVX1_LOC_292/A INVX1_LOC_63/A 0.07fF
C18310 NAND2X1_LOC_198/B NOR2X1_LOC_743/Y 0.10fF
C18311 INVX1_LOC_75/A NOR2X1_LOC_356/A 0.84fF
C18312 INVX1_LOC_41/A NOR2X1_LOC_536/A 0.06fF
C18313 INVX1_LOC_138/A NAND2X1_LOC_223/A 0.01fF
C18314 INVX1_LOC_72/A INVX1_LOC_107/Y 0.03fF
C18315 INVX1_LOC_174/A NOR2X1_LOC_258/Y 0.02fF
C18316 INVX1_LOC_47/A NOR2X1_LOC_721/Y 0.00fF
C18317 NOR2X1_LOC_498/Y NOR2X1_LOC_536/A 0.19fF
C18318 D_INPUT_0 NOR2X1_LOC_703/Y 0.00fF
C18319 INVX1_LOC_296/Y INVX1_LOC_173/A 0.01fF
C18320 INVX1_LOC_151/Y INVX1_LOC_147/Y 0.03fF
C18321 INVX1_LOC_196/A VDD 1.05fF
C18322 NOR2X1_LOC_401/B NOR2X1_LOC_266/B 0.01fF
C18323 INVX1_LOC_278/A INVX1_LOC_26/A 0.10fF
C18324 INVX1_LOC_298/Y INVX1_LOC_64/A 0.07fF
C18325 INVX1_LOC_58/A INVX1_LOC_50/A 0.11fF
C18326 NOR2X1_LOC_355/A NOR2X1_LOC_355/B 0.05fF
C18327 INVX1_LOC_309/Y NOR2X1_LOC_491/Y 0.01fF
C18328 NOR2X1_LOC_860/B NOR2X1_LOC_61/A 0.01fF
C18329 INVX1_LOC_33/A INVX1_LOC_118/A 0.11fF
C18330 NOR2X1_LOC_469/a_36_216# INVX1_LOC_102/A 0.01fF
C18331 INVX1_LOC_111/A NOR2X1_LOC_831/B 0.01fF
C18332 INVX1_LOC_282/A NAND2X1_LOC_560/A 0.06fF
C18333 NOR2X1_LOC_255/a_36_216# NOR2X1_LOC_124/A 0.00fF
C18334 NOR2X1_LOC_717/B NOR2X1_LOC_78/A 0.01fF
C18335 NAND2X1_LOC_477/A NOR2X1_LOC_536/A 0.45fF
C18336 INVX1_LOC_124/A INVX1_LOC_66/Y 0.06fF
C18337 INVX1_LOC_35/A NOR2X1_LOC_831/a_36_216# 0.00fF
C18338 NOR2X1_LOC_666/A INVX1_LOC_15/A 0.24fF
C18339 NAND2X1_LOC_841/A VDD -0.00fF
C18340 NOR2X1_LOC_287/A VDD 0.12fF
C18341 INVX1_LOC_200/Y NAND2X1_LOC_787/A 0.01fF
C18342 INVX1_LOC_77/A NOR2X1_LOC_259/B 0.03fF
C18343 INVX1_LOC_201/Y NOR2X1_LOC_655/Y 0.05fF
C18344 INVX1_LOC_75/A NOR2X1_LOC_74/A 0.21fF
C18345 NOR2X1_LOC_615/Y NAND2X1_LOC_254/Y 0.01fF
C18346 NOR2X1_LOC_361/a_36_216# INVX1_LOC_272/A 0.08fF
C18347 INVX1_LOC_278/A NAND2X1_LOC_564/A 0.02fF
C18348 INVX1_LOC_41/A NAND2X1_LOC_93/B 0.10fF
C18349 NOR2X1_LOC_220/A NAND2X1_LOC_472/Y 0.10fF
C18350 INVX1_LOC_268/A VDD 0.47fF
C18351 NOR2X1_LOC_790/B INVX1_LOC_23/A 0.09fF
C18352 NOR2X1_LOC_795/Y NOR2X1_LOC_729/A 0.10fF
C18353 NOR2X1_LOC_828/A NOR2X1_LOC_78/A 0.01fF
C18354 INVX1_LOC_289/A INVX1_LOC_77/Y 0.03fF
C18355 INVX1_LOC_45/A NAND2X1_LOC_639/a_36_24# 0.01fF
C18356 NOR2X1_LOC_91/A NAND2X1_LOC_169/Y 0.01fF
C18357 NAND2X1_LOC_360/B NOR2X1_LOC_271/Y 0.31fF
C18358 INVX1_LOC_75/A NOR2X1_LOC_9/Y 0.10fF
C18359 INVX1_LOC_210/A INVX1_LOC_9/A 0.02fF
C18360 INVX1_LOC_132/A NAND2X1_LOC_572/B 0.17fF
C18361 INVX1_LOC_2/A NOR2X1_LOC_351/Y 2.01fF
C18362 INVX1_LOC_226/Y NAND2X1_LOC_96/A 0.62fF
C18363 INVX1_LOC_314/Y NOR2X1_LOC_814/A 0.01fF
C18364 NOR2X1_LOC_208/Y NOR2X1_LOC_631/A 0.01fF
C18365 INVX1_LOC_224/Y INVX1_LOC_13/Y 0.27fF
C18366 NOR2X1_LOC_186/Y NOR2X1_LOC_654/A 0.16fF
C18367 NAND2X1_LOC_214/B NOR2X1_LOC_414/Y 0.28fF
C18368 NAND2X1_LOC_709/a_36_24# INVX1_LOC_186/A 0.00fF
C18369 NOR2X1_LOC_478/A NOR2X1_LOC_477/B 0.09fF
C18370 NOR2X1_LOC_160/B INVX1_LOC_47/Y 0.00fF
C18371 NAND2X1_LOC_798/A INVX1_LOC_118/A 0.03fF
C18372 INVX1_LOC_295/A INVX1_LOC_115/A 0.03fF
C18373 INVX1_LOC_142/A NOR2X1_LOC_833/B 0.02fF
C18374 INVX1_LOC_61/Y INVX1_LOC_3/Y 0.08fF
C18375 INVX1_LOC_176/A NOR2X1_LOC_559/a_36_216# 0.00fF
C18376 NOR2X1_LOC_372/Y INVX1_LOC_42/A 0.01fF
C18377 NAND2X1_LOC_338/B NOR2X1_LOC_99/Y 1.35fF
C18378 INVX1_LOC_41/A INVX1_LOC_3/A 0.02fF
C18379 INVX1_LOC_269/A INVX1_LOC_23/Y 0.10fF
C18380 NAND2X1_LOC_735/B INVX1_LOC_38/A 0.02fF
C18381 INVX1_LOC_201/Y INVX1_LOC_3/A 2.50fF
C18382 INVX1_LOC_269/A NAND2X1_LOC_72/a_36_24# 0.00fF
C18383 NAND2X1_LOC_573/Y NOR2X1_LOC_654/A 0.00fF
C18384 NOR2X1_LOC_15/Y NOR2X1_LOC_39/Y 0.03fF
C18385 INVX1_LOC_90/A D_INPUT_3 0.07fF
C18386 INVX1_LOC_47/A VDD 0.41fF
C18387 INVX1_LOC_13/A INVX1_LOC_9/A 5.72fF
C18388 INPUT_5 INVX1_LOC_38/A 0.02fF
C18389 INVX1_LOC_90/A INVX1_LOC_14/Y 0.03fF
C18390 VDD INVX1_LOC_175/Y 0.01fF
C18391 NOR2X1_LOC_68/A NOR2X1_LOC_477/B 0.03fF
C18392 NOR2X1_LOC_2/Y INPUT_4 0.06fF
C18393 NAND2X1_LOC_21/Y NOR2X1_LOC_36/B 0.04fF
C18394 NOR2X1_LOC_299/Y NOR2X1_LOC_536/A 0.10fF
C18395 NOR2X1_LOC_844/A NAND2X1_LOC_206/Y 0.02fF
C18396 INVX1_LOC_166/A INVX1_LOC_14/A 0.41fF
C18397 INVX1_LOC_64/A NAND2X1_LOC_344/a_36_24# 0.00fF
C18398 INVX1_LOC_53/Y NOR2X1_LOC_743/Y 0.23fF
C18399 INVX1_LOC_170/A NOR2X1_LOC_394/Y 0.05fF
C18400 NOR2X1_LOC_276/B INVX1_LOC_15/A 0.02fF
C18401 NAND2X1_LOC_551/a_36_24# INVX1_LOC_14/A 0.01fF
C18402 INVX1_LOC_89/A NAND2X1_LOC_848/A 0.03fF
C18403 NOR2X1_LOC_685/A NAND2X1_LOC_682/a_36_24# 0.02fF
C18404 INVX1_LOC_120/A NOR2X1_LOC_865/A 0.01fF
C18405 NOR2X1_LOC_51/A INPUT_5 0.05fF
C18406 NAND2X1_LOC_348/A D_INPUT_3 0.03fF
C18407 INVX1_LOC_225/Y NOR2X1_LOC_383/B 0.25fF
C18408 INVX1_LOC_286/A NOR2X1_LOC_124/A 0.03fF
C18409 INVX1_LOC_90/A INVX1_LOC_230/A 0.12fF
C18410 D_GATE_741 INVX1_LOC_23/A 0.02fF
C18411 INVX1_LOC_121/A NAND2X1_LOC_93/B 0.03fF
C18412 INVX1_LOC_17/A INVX1_LOC_53/A 0.15fF
C18413 NOR2X1_LOC_205/Y NOR2X1_LOC_678/A 1.06fF
C18414 NAND2X1_LOC_276/Y INVX1_LOC_42/A 0.07fF
C18415 INVX1_LOC_24/A NOR2X1_LOC_38/B 0.46fF
C18416 INVX1_LOC_16/A NOR2X1_LOC_697/Y 0.00fF
C18417 INVX1_LOC_5/A NAND2X1_LOC_218/A 0.01fF
C18418 INVX1_LOC_111/Y INVX1_LOC_19/A 0.01fF
C18419 INVX1_LOC_77/A INVX1_LOC_32/A 0.10fF
C18420 INVX1_LOC_73/A NOR2X1_LOC_363/Y 0.12fF
C18421 INVX1_LOC_104/A NOR2X1_LOC_89/A 0.07fF
C18422 INVX1_LOC_279/A NOR2X1_LOC_197/B 0.10fF
C18423 INVX1_LOC_5/A NOR2X1_LOC_140/A 0.01fF
C18424 NAND2X1_LOC_733/Y INVX1_LOC_296/A 0.01fF
C18425 INVX1_LOC_55/Y INVX1_LOC_9/A -0.02fF
C18426 NOR2X1_LOC_315/Y INVX1_LOC_12/A 0.17fF
C18427 NOR2X1_LOC_152/Y INVX1_LOC_231/A 0.04fF
C18428 NAND2X1_LOC_352/B INVX1_LOC_23/A 0.07fF
C18429 INVX1_LOC_121/A NAND2X1_LOC_425/Y 0.02fF
C18430 INVX1_LOC_77/A NOR2X1_LOC_623/B 0.06fF
C18431 NOR2X1_LOC_432/Y INVX1_LOC_12/A 0.04fF
C18432 INVX1_LOC_17/Y INVX1_LOC_30/A 0.01fF
C18433 INVX1_LOC_89/A INVX1_LOC_46/Y 0.13fF
C18434 NAND2X1_LOC_850/Y INVX1_LOC_29/A 0.10fF
C18435 NAND2X1_LOC_348/A INVX1_LOC_230/A 0.34fF
C18436 INVX1_LOC_300/Y NOR2X1_LOC_829/A 0.16fF
C18437 NOR2X1_LOC_335/A INVX1_LOC_4/Y 0.01fF
C18438 INVX1_LOC_40/A NAND2X1_LOC_63/Y 0.02fF
C18439 INVX1_LOC_104/A NOR2X1_LOC_170/A 0.00fF
C18440 NAND2X1_LOC_363/B NAND2X1_LOC_113/a_36_24# 0.01fF
C18441 INVX1_LOC_8/A INVX1_LOC_4/A 0.07fF
C18442 NAND2X1_LOC_795/a_36_24# NOR2X1_LOC_48/B 0.00fF
C18443 NOR2X1_LOC_588/A VDD 0.24fF
C18444 INVX1_LOC_13/Y NOR2X1_LOC_103/Y 0.15fF
C18445 NOR2X1_LOC_667/A INVX1_LOC_102/A 0.08fF
C18446 INVX1_LOC_178/A NAND2X1_LOC_538/Y 0.10fF
C18447 NAND2X1_LOC_714/B NAND2X1_LOC_537/Y 0.07fF
C18448 INVX1_LOC_5/A NOR2X1_LOC_530/Y 0.08fF
C18449 INVX1_LOC_83/A NOR2X1_LOC_450/B 0.03fF
C18450 INVX1_LOC_18/A INVX1_LOC_57/A 0.14fF
C18451 NAND2X1_LOC_374/Y INVX1_LOC_42/A 0.18fF
C18452 NAND2X1_LOC_571/B INVX1_LOC_30/A 0.01fF
C18453 NOR2X1_LOC_262/Y INVX1_LOC_26/A 0.01fF
C18454 NOR2X1_LOC_32/B NOR2X1_LOC_382/Y 0.69fF
C18455 NAND2X1_LOC_394/a_36_24# NAND2X1_LOC_555/Y 0.00fF
C18456 NOR2X1_LOC_598/B INVX1_LOC_142/A 0.07fF
C18457 NAND2X1_LOC_557/Y NOR2X1_LOC_522/Y 0.33fF
C18458 INPUT_0 NOR2X1_LOC_332/Y 0.02fF
C18459 INVX1_LOC_83/A NOR2X1_LOC_257/Y 0.01fF
C18460 D_INPUT_1 NOR2X1_LOC_360/Y 0.12fF
C18461 NAND2X1_LOC_341/A INVX1_LOC_109/Y 0.00fF
C18462 NAND2X1_LOC_783/Y NOR2X1_LOC_186/Y 0.01fF
C18463 INVX1_LOC_95/Y VDD 3.03fF
C18464 INVX1_LOC_120/A INVX1_LOC_63/A 0.46fF
C18465 INVX1_LOC_187/Y VDD 0.21fF
C18466 NOR2X1_LOC_637/Y INVX1_LOC_57/A 0.03fF
C18467 NAND2X1_LOC_708/Y INVX1_LOC_72/A 0.05fF
C18468 NAND2X1_LOC_477/A NAND2X1_LOC_470/B 0.04fF
C18469 INVX1_LOC_35/A NOR2X1_LOC_68/A 0.33fF
C18470 INVX1_LOC_64/A INVX1_LOC_247/Y 0.03fF
C18471 INVX1_LOC_49/A INVX1_LOC_275/Y 0.00fF
C18472 NOR2X1_LOC_137/A INVX1_LOC_19/A 0.22fF
C18473 NAND2X1_LOC_854/B NOR2X1_LOC_89/A 0.19fF
C18474 INVX1_LOC_34/A NOR2X1_LOC_693/Y 0.02fF
C18475 INVX1_LOC_172/A INVX1_LOC_57/A 0.17fF
C18476 INVX1_LOC_49/A NOR2X1_LOC_748/A 0.08fF
C18477 INVX1_LOC_45/A INVX1_LOC_13/Y 0.07fF
C18478 NOR2X1_LOC_65/B NAND2X1_LOC_276/Y 0.01fF
C18479 INVX1_LOC_58/A INVX1_LOC_105/A 1.51fF
C18480 NAND2X1_LOC_783/Y NAND2X1_LOC_573/Y 0.01fF
C18481 NOR2X1_LOC_139/Y NOR2X1_LOC_331/B 0.07fF
C18482 VDD NOR2X1_LOC_305/Y 0.65fF
C18483 INVX1_LOC_13/Y NOR2X1_LOC_568/A 0.00fF
C18484 NOR2X1_LOC_78/A NOR2X1_LOC_709/B 0.02fF
C18485 NOR2X1_LOC_448/A INVX1_LOC_38/A 0.00fF
C18486 INVX1_LOC_37/Y NAND2X1_LOC_241/Y 0.00fF
C18487 INVX1_LOC_40/Y INVX1_LOC_27/A 0.02fF
C18488 NAND2X1_LOC_787/A NOR2X1_LOC_495/Y 0.03fF
C18489 NOR2X1_LOC_91/A NAND2X1_LOC_357/B 0.14fF
C18490 INVX1_LOC_21/A INVX1_LOC_223/A 1.38fF
C18491 NAND2X1_LOC_374/Y INVX1_LOC_78/A 0.01fF
C18492 NAND2X1_LOC_538/Y NOR2X1_LOC_816/A 0.77fF
C18493 INVX1_LOC_236/Y NAND2X1_LOC_579/A 0.09fF
C18494 INVX1_LOC_6/A NOR2X1_LOC_831/B 0.07fF
C18495 NOR2X1_LOC_344/A INVX1_LOC_23/A 0.04fF
C18496 NAND2X1_LOC_125/a_36_24# NOR2X1_LOC_847/B 0.00fF
C18497 NAND2X1_LOC_725/Y NAND2X1_LOC_736/B 0.34fF
C18498 INVX1_LOC_225/A NOR2X1_LOC_654/A 0.00fF
C18499 NAND2X1_LOC_794/B NOR2X1_LOC_518/Y 0.03fF
C18500 INVX1_LOC_284/Y NAND2X1_LOC_579/A 0.02fF
C18501 NAND2X1_LOC_468/B NOR2X1_LOC_331/B 0.10fF
C18502 NOR2X1_LOC_360/Y NOR2X1_LOC_652/Y -0.02fF
C18503 INVX1_LOC_91/A INVX1_LOC_291/A 0.07fF
C18504 INVX1_LOC_249/A NOR2X1_LOC_665/Y 0.01fF
C18505 NAND2X1_LOC_725/Y GATE_811 0.03fF
C18506 NOR2X1_LOC_772/B INVX1_LOC_71/A 0.10fF
C18507 NAND2X1_LOC_738/B NAND2X1_LOC_811/Y 0.04fF
C18508 INVX1_LOC_37/A INVX1_LOC_77/Y 0.07fF
C18509 NOR2X1_LOC_514/Y INVX1_LOC_23/A 0.01fF
C18510 NOR2X1_LOC_313/Y INVX1_LOC_84/A 0.05fF
C18511 INVX1_LOC_266/Y NOR2X1_LOC_383/B 0.25fF
C18512 NOR2X1_LOC_644/A INVX1_LOC_99/A 0.04fF
C18513 INVX1_LOC_38/A NOR2X1_LOC_853/a_36_216# 0.02fF
C18514 INVX1_LOC_13/Y INVX1_LOC_71/A 0.08fF
C18515 INVX1_LOC_45/A INVX1_LOC_88/A 0.06fF
C18516 INVX1_LOC_72/A NOR2X1_LOC_271/B 0.03fF
C18517 INVX1_LOC_34/Y INVX1_LOC_57/A 0.07fF
C18518 INVX1_LOC_14/Y INVX1_LOC_38/A 0.03fF
C18519 NOR2X1_LOC_84/A NOR2X1_LOC_660/Y 0.08fF
C18520 INVX1_LOC_304/A INVX1_LOC_70/A 0.01fF
C18521 NOR2X1_LOC_657/B NOR2X1_LOC_364/A 0.13fF
C18522 NOR2X1_LOC_285/Y NOR2X1_LOC_285/B 0.02fF
C18523 INVX1_LOC_64/A INVX1_LOC_8/A 0.90fF
C18524 NOR2X1_LOC_231/B NOR2X1_LOC_160/B 0.09fF
C18525 INVX1_LOC_226/Y NAND2X1_LOC_99/A 0.01fF
C18526 NOR2X1_LOC_223/B INVX1_LOC_103/Y 0.38fF
C18527 NOR2X1_LOC_130/A NOR2X1_LOC_38/B 0.01fF
C18528 NOR2X1_LOC_740/Y INVX1_LOC_142/Y 0.03fF
C18529 NAND2X1_LOC_642/Y NAND2X1_LOC_572/B 0.10fF
C18530 NOR2X1_LOC_340/Y INVX1_LOC_50/Y 0.10fF
C18531 NOR2X1_LOC_468/Y INVX1_LOC_24/A 0.01fF
C18532 NAND2X1_LOC_638/Y NOR2X1_LOC_467/A 0.03fF
C18533 NAND2X1_LOC_796/Y NAND2X1_LOC_175/Y 0.05fF
C18534 NOR2X1_LOC_557/A NOR2X1_LOC_814/A 0.02fF
C18535 NOR2X1_LOC_561/Y NOR2X1_LOC_25/Y 0.18fF
C18536 NOR2X1_LOC_637/B NOR2X1_LOC_173/Y 0.01fF
C18537 NOR2X1_LOC_602/a_36_216# NAND2X1_LOC_337/B 0.00fF
C18538 INVX1_LOC_35/A NAND2X1_LOC_134/a_36_24# 0.00fF
C18539 INVX1_LOC_39/A INVX1_LOC_33/A 0.03fF
C18540 INVX1_LOC_150/Y INVX1_LOC_72/A 0.07fF
C18541 INVX1_LOC_48/A INVX1_LOC_19/A 0.03fF
C18542 NAND2X1_LOC_190/Y INVX1_LOC_24/A 0.05fF
C18543 NAND2X1_LOC_348/A NAND2X1_LOC_233/a_36_24# 0.00fF
C18544 NOR2X1_LOC_740/Y INVX1_LOC_198/Y 0.19fF
C18545 NAND2X1_LOC_844/a_36_24# INVX1_LOC_42/A 0.00fF
C18546 NAND2X1_LOC_560/A NOR2X1_LOC_496/a_36_216# 0.00fF
C18547 NAND2X1_LOC_276/Y NOR2X1_LOC_655/a_36_216# 0.02fF
C18548 NAND2X1_LOC_214/B NAND2X1_LOC_122/a_36_24# 0.00fF
C18549 NOR2X1_LOC_792/B NOR2X1_LOC_652/Y 0.05fF
C18550 INVX1_LOC_88/A INVX1_LOC_71/A 0.13fF
C18551 INVX1_LOC_38/A INVX1_LOC_230/A 0.00fF
C18552 NOR2X1_LOC_348/B NOR2X1_LOC_644/a_36_216# 0.00fF
C18553 INVX1_LOC_21/A INVX1_LOC_149/Y 0.05fF
C18554 NOR2X1_LOC_706/B INVX1_LOC_92/A 0.04fF
C18555 NAND2X1_LOC_739/B INVX1_LOC_161/Y 0.09fF
C18556 INVX1_LOC_21/A INVX1_LOC_85/A 0.03fF
C18557 INVX1_LOC_25/A NOR2X1_LOC_789/A 0.04fF
C18558 INVX1_LOC_45/A NOR2X1_LOC_500/B 0.28fF
C18559 NOR2X1_LOC_468/Y NOR2X1_LOC_557/Y 0.08fF
C18560 NOR2X1_LOC_15/Y NOR2X1_LOC_570/B 0.05fF
C18561 INVX1_LOC_101/Y NOR2X1_LOC_388/Y 0.02fF
C18562 NOR2X1_LOC_617/Y NOR2X1_LOC_372/A -0.01fF
C18563 D_INPUT_4 NOR2X1_LOC_36/A 0.14fF
C18564 INVX1_LOC_41/A INVX1_LOC_256/A 0.02fF
C18565 INVX1_LOC_278/A INVX1_LOC_164/A 0.23fF
C18566 NOR2X1_LOC_170/a_36_216# NOR2X1_LOC_568/A 0.01fF
C18567 INVX1_LOC_39/A INVX1_LOC_40/A 0.12fF
C18568 INVX1_LOC_76/A INVX1_LOC_264/A 0.02fF
C18569 INVX1_LOC_2/A NOR2X1_LOC_669/Y 0.02fF
C18570 NAND2X1_LOC_175/B INVX1_LOC_246/A 0.01fF
C18571 NOR2X1_LOC_318/B NOR2X1_LOC_116/a_36_216# -0.02fF
C18572 INVX1_LOC_70/Y INVX1_LOC_170/Y 0.15fF
C18573 INVX1_LOC_1/A NOR2X1_LOC_168/B 0.01fF
C18574 INVX1_LOC_11/A INVX1_LOC_104/A 0.25fF
C18575 INVX1_LOC_201/Y NOR2X1_LOC_647/B 0.04fF
C18576 D_INPUT_0 NOR2X1_LOC_392/Y 0.18fF
C18577 NOR2X1_LOC_468/Y INVX1_LOC_143/A 0.00fF
C18578 INVX1_LOC_200/A NOR2X1_LOC_315/Y 0.00fF
C18579 NOR2X1_LOC_669/Y NOR2X1_LOC_226/A 0.38fF
C18580 INVX1_LOC_45/A INVX1_LOC_303/A 0.01fF
C18581 INVX1_LOC_43/Y INVX1_LOC_8/A -0.00fF
C18582 NAND2X1_LOC_53/Y NOR2X1_LOC_423/Y 0.01fF
C18583 INVX1_LOC_136/A NOR2X1_LOC_303/Y 0.12fF
C18584 NAND2X1_LOC_361/Y INVX1_LOC_30/A 0.02fF
C18585 INVX1_LOC_24/A INVX1_LOC_62/Y 0.07fF
C18586 INVX1_LOC_299/A NOR2X1_LOC_566/Y 0.01fF
C18587 INVX1_LOC_58/A NAND2X1_LOC_652/Y 0.02fF
C18588 INVX1_LOC_218/Y NOR2X1_LOC_6/B 0.22fF
C18589 INVX1_LOC_17/A NOR2X1_LOC_78/B 0.14fF
C18590 INVX1_LOC_45/A NAND2X1_LOC_59/B 0.03fF
C18591 INVX1_LOC_177/Y NOR2X1_LOC_433/A 0.01fF
C18592 NOR2X1_LOC_337/Y INVX1_LOC_271/Y 0.02fF
C18593 NOR2X1_LOC_208/Y NOR2X1_LOC_735/a_36_216# 0.00fF
C18594 INVX1_LOC_24/A NOR2X1_LOC_596/A 1.97fF
C18595 NOR2X1_LOC_831/B INVX1_LOC_131/Y 0.19fF
C18596 NOR2X1_LOC_170/a_36_216# INVX1_LOC_71/A 0.00fF
C18597 NAND2X1_LOC_357/B INVX1_LOC_31/A 0.07fF
C18598 NAND2X1_LOC_574/A NOR2X1_LOC_655/Y 0.09fF
C18599 NOR2X1_LOC_598/B NOR2X1_LOC_535/a_36_216# 0.01fF
C18600 INVX1_LOC_73/A INVX1_LOC_29/Y 0.04fF
C18601 NOR2X1_LOC_99/B INVX1_LOC_50/Y 0.07fF
C18602 NAND2X1_LOC_53/Y NOR2X1_LOC_222/Y 0.07fF
C18603 INVX1_LOC_40/Y NOR2X1_LOC_664/Y 0.01fF
C18604 INVX1_LOC_256/A NOR2X1_LOC_405/a_36_216# 0.01fF
C18605 INVX1_LOC_269/A INVX1_LOC_232/A 0.10fF
C18606 INVX1_LOC_188/A INVX1_LOC_177/A 0.00fF
C18607 NAND2X1_LOC_483/Y NOR2X1_LOC_384/Y 0.04fF
C18608 NOR2X1_LOC_637/B NOR2X1_LOC_637/A 0.07fF
C18609 NOR2X1_LOC_644/Y NOR2X1_LOC_644/B 0.01fF
C18610 NAND2X1_LOC_648/A NOR2X1_LOC_304/Y 0.02fF
C18611 NAND2X1_LOC_276/Y NOR2X1_LOC_554/B 0.03fF
C18612 INVX1_LOC_48/A INVX1_LOC_26/Y 0.03fF
C18613 INVX1_LOC_123/A INVX1_LOC_26/A 0.04fF
C18614 NOR2X1_LOC_185/a_36_216# INVX1_LOC_57/A 0.00fF
C18615 NOR2X1_LOC_471/Y NOR2X1_LOC_78/B 0.03fF
C18616 NOR2X1_LOC_858/B NOR2X1_LOC_850/B 0.11fF
C18617 NOR2X1_LOC_843/A INVX1_LOC_305/A 0.03fF
C18618 NOR2X1_LOC_430/Y INVX1_LOC_92/A 0.26fF
C18619 NOR2X1_LOC_61/B INVX1_LOC_135/A 0.12fF
C18620 NOR2X1_LOC_590/A NOR2X1_LOC_778/B 0.23fF
C18621 INVX1_LOC_269/A NOR2X1_LOC_383/Y 0.10fF
C18622 NAND2X1_LOC_549/B INVX1_LOC_31/A 0.01fF
C18623 NAND2X1_LOC_624/B NAND2X1_LOC_560/A 0.83fF
C18624 INPUT_4 NOR2X1_LOC_36/A 0.12fF
C18625 NOR2X1_LOC_332/A NAND2X1_LOC_218/A 0.04fF
C18626 INVX1_LOC_34/A INVX1_LOC_45/Y 0.03fF
C18627 NOR2X1_LOC_272/Y NOR2X1_LOC_473/B 0.31fF
C18628 INVX1_LOC_132/A NOR2X1_LOC_419/Y 0.01fF
C18629 NOR2X1_LOC_140/A NOR2X1_LOC_332/A 0.07fF
C18630 NOR2X1_LOC_68/A INVX1_LOC_257/Y -0.00fF
C18631 INVX1_LOC_278/A NOR2X1_LOC_368/A 0.02fF
C18632 INVX1_LOC_250/A NAND2X1_LOC_722/A 0.03fF
C18633 NAND2X1_LOC_667/a_36_24# NOR2X1_LOC_68/A 0.00fF
C18634 NOR2X1_LOC_468/Y NOR2X1_LOC_130/A 0.03fF
C18635 INVX1_LOC_136/A INVX1_LOC_54/Y 0.78fF
C18636 INVX1_LOC_132/A NOR2X1_LOC_716/B 0.04fF
C18637 INVX1_LOC_182/A INVX1_LOC_50/Y 0.07fF
C18638 NOR2X1_LOC_215/Y NOR2X1_LOC_52/B 0.00fF
C18639 NAND2X1_LOC_468/B NOR2X1_LOC_449/A 0.31fF
C18640 NOR2X1_LOC_158/Y INVX1_LOC_76/A 0.10fF
C18641 NAND2X1_LOC_574/A INVX1_LOC_3/A 0.07fF
C18642 NOR2X1_LOC_319/B NOR2X1_LOC_812/A 0.13fF
C18643 NOR2X1_LOC_716/B NAND2X1_LOC_640/Y 0.00fF
C18644 INVX1_LOC_17/A INVX1_LOC_83/A 1.10fF
C18645 INVX1_LOC_211/Y NOR2X1_LOC_561/Y 0.08fF
C18646 NOR2X1_LOC_550/B NOR2X1_LOC_486/B 0.21fF
C18647 INVX1_LOC_90/A NAND2X1_LOC_303/Y 0.05fF
C18648 VDD INVX1_LOC_271/Y 1.66fF
C18649 NOR2X1_LOC_82/A INVX1_LOC_306/A 0.03fF
C18650 NAND2X1_LOC_67/Y INVX1_LOC_55/Y 0.11fF
C18651 INVX1_LOC_77/A INVX1_LOC_158/A 0.03fF
C18652 INVX1_LOC_36/A INVX1_LOC_56/Y 0.03fF
C18653 NAND2X1_LOC_818/a_36_24# NOR2X1_LOC_649/B 0.01fF
C18654 NOR2X1_LOC_657/Y INVX1_LOC_22/A 0.03fF
C18655 INVX1_LOC_161/Y NOR2X1_LOC_137/A 0.19fF
C18656 NOR2X1_LOC_82/A NOR2X1_LOC_132/a_36_216# 0.01fF
C18657 INVX1_LOC_35/Y NAND2X1_LOC_74/B 0.94fF
C18658 NOR2X1_LOC_658/Y INVX1_LOC_290/A 0.10fF
C18659 NOR2X1_LOC_301/A INVX1_LOC_46/A 0.03fF
C18660 NAND2X1_LOC_555/Y NOR2X1_LOC_459/A -0.03fF
C18661 NAND2X1_LOC_30/Y INVX1_LOC_89/A 0.06fF
C18662 NOR2X1_LOC_295/Y NOR2X1_LOC_557/Y 0.04fF
C18663 INVX1_LOC_100/A INVX1_LOC_306/Y 0.03fF
C18664 NOR2X1_LOC_791/A INVX1_LOC_25/Y 0.01fF
C18665 NOR2X1_LOC_593/Y INVX1_LOC_104/A 0.14fF
C18666 NOR2X1_LOC_426/a_36_216# INPUT_5 0.00fF
C18667 NAND2X1_LOC_628/a_36_24# INVX1_LOC_193/A 0.00fF
C18668 INVX1_LOC_32/A INVX1_LOC_9/A 0.28fF
C18669 NAND2X1_LOC_722/A NOR2X1_LOC_495/Y 0.01fF
C18670 NOR2X1_LOC_128/B INVX1_LOC_31/A 0.01fF
C18671 NOR2X1_LOC_220/A INVX1_LOC_24/A 0.02fF
C18672 NOR2X1_LOC_646/B INVX1_LOC_76/A 0.00fF
C18673 NAND2X1_LOC_291/B NOR2X1_LOC_865/Y 0.12fF
C18674 INVX1_LOC_272/Y NOR2X1_LOC_329/B 0.43fF
C18675 INVX1_LOC_12/Y INVX1_LOC_23/Y 0.10fF
C18676 NAND2X1_LOC_198/B INVX1_LOC_53/Y 0.10fF
C18677 NAND2X1_LOC_538/Y INVX1_LOC_140/A 0.10fF
C18678 INVX1_LOC_226/Y NAND2X1_LOC_656/A 0.00fF
C18679 NAND2X1_LOC_291/B NOR2X1_LOC_243/B 0.12fF
C18680 INVX1_LOC_174/A D_GATE_366 0.07fF
C18681 NAND2X1_LOC_208/B NOR2X1_LOC_71/Y 0.04fF
C18682 NOR2X1_LOC_103/a_36_216# INVX1_LOC_42/A 0.01fF
C18683 NOR2X1_LOC_52/B INVX1_LOC_104/A 0.10fF
C18684 INVX1_LOC_314/Y NOR2X1_LOC_82/Y 0.01fF
C18685 INVX1_LOC_304/Y NOR2X1_LOC_315/Y 0.02fF
C18686 INVX1_LOC_24/A NOR2X1_LOC_548/Y 0.07fF
C18687 D_INPUT_0 NOR2X1_LOC_86/Y 0.07fF
C18688 INVX1_LOC_24/Y INVX1_LOC_69/Y 0.02fF
C18689 INVX1_LOC_308/A NAND2X1_LOC_287/B 0.03fF
C18690 NAND2X1_LOC_364/Y NAND2X1_LOC_282/a_36_24# 0.00fF
C18691 INVX1_LOC_263/A NOR2X1_LOC_593/Y 0.07fF
C18692 NOR2X1_LOC_15/Y INVX1_LOC_286/A 0.15fF
C18693 NOR2X1_LOC_782/a_36_216# INVX1_LOC_290/A 0.00fF
C18694 INVX1_LOC_77/A GATE_662 0.07fF
C18695 NAND2X1_LOC_308/B NAND2X1_LOC_856/A 0.01fF
C18696 NOR2X1_LOC_238/Y NOR2X1_LOC_528/a_36_216# 0.00fF
C18697 INVX1_LOC_94/Y INVX1_LOC_92/A 0.07fF
C18698 D_INPUT_0 NOR2X1_LOC_744/a_36_216# 0.02fF
C18699 NOR2X1_LOC_788/B NOR2X1_LOC_703/B 0.02fF
C18700 INVX1_LOC_10/A NOR2X1_LOC_484/Y 0.03fF
C18701 INVX1_LOC_30/A NAND2X1_LOC_654/B 0.06fF
C18702 INVX1_LOC_196/A INVX1_LOC_177/A 0.00fF
C18703 INVX1_LOC_40/Y NOR2X1_LOC_19/B 0.01fF
C18704 INVX1_LOC_222/Y NOR2X1_LOC_799/B 0.01fF
C18705 NOR2X1_LOC_575/a_36_216# NAND2X1_LOC_463/B 0.00fF
C18706 INVX1_LOC_256/Y NOR2X1_LOC_84/Y 0.01fF
C18707 INVX1_LOC_106/Y NAND2X1_LOC_63/Y 0.01fF
C18708 NAND2X1_LOC_114/B NOR2X1_LOC_188/A 0.05fF
C18709 INVX1_LOC_269/A INVX1_LOC_186/A 0.07fF
C18710 INVX1_LOC_11/A INVX1_LOC_206/Y 0.08fF
C18711 NOR2X1_LOC_773/Y NOR2X1_LOC_709/A 0.00fF
C18712 INVX1_LOC_36/A NOR2X1_LOC_385/Y 0.04fF
C18713 INVX1_LOC_124/Y INVX1_LOC_75/A 0.23fF
C18714 NAND2X1_LOC_114/B NOR2X1_LOC_548/B 0.07fF
C18715 INVX1_LOC_41/A NOR2X1_LOC_440/Y 0.01fF
C18716 INVX1_LOC_11/A INVX1_LOC_86/Y 0.23fF
C18717 NOR2X1_LOC_646/a_36_216# NOR2X1_LOC_664/Y 0.00fF
C18718 NOR2X1_LOC_226/A NOR2X1_LOC_401/B 0.03fF
C18719 NOR2X1_LOC_717/B NOR2X1_LOC_374/A 0.07fF
C18720 NOR2X1_LOC_15/Y INVX1_LOC_95/A 0.03fF
C18721 NAND2X1_LOC_848/A NOR2X1_LOC_392/Y 0.00fF
C18722 INVX1_LOC_202/A NAND2X1_LOC_128/a_36_24# 0.00fF
C18723 NOR2X1_LOC_320/a_36_216# NAND2X1_LOC_660/Y 0.03fF
C18724 INVX1_LOC_17/A NOR2X1_LOC_311/Y 0.01fF
C18725 NOR2X1_LOC_689/Y INVX1_LOC_185/A 0.01fF
C18726 INVX1_LOC_35/A NOR2X1_LOC_114/a_36_216# 0.00fF
C18727 INVX1_LOC_89/A INVX1_LOC_49/A 1.58fF
C18728 NAND2X1_LOC_594/a_36_24# NAND2X1_LOC_287/B 0.01fF
C18729 INVX1_LOC_224/Y NOR2X1_LOC_99/Y 0.15fF
C18730 INVX1_LOC_296/A INVX1_LOC_92/A 2.70fF
C18731 INVX1_LOC_201/Y NOR2X1_LOC_415/A 0.06fF
C18732 NAND2X1_LOC_68/a_36_24# INVX1_LOC_139/A 0.01fF
C18733 INVX1_LOC_11/A NOR2X1_LOC_600/Y 0.98fF
C18734 NAND2X1_LOC_35/Y NOR2X1_LOC_536/A 0.13fF
C18735 NOR2X1_LOC_74/A NOR2X1_LOC_274/B 0.07fF
C18736 INVX1_LOC_269/A NAND2X1_LOC_447/Y 0.10fF
C18737 INVX1_LOC_34/A NOR2X1_LOC_71/Y 0.07fF
C18738 NOR2X1_LOC_828/A NOR2X1_LOC_374/A 0.00fF
C18739 NOR2X1_LOC_521/a_36_216# NAND2X1_LOC_735/B 0.00fF
C18740 INVX1_LOC_59/A VDD -0.00fF
C18741 NAND2X1_LOC_149/Y INVX1_LOC_37/A 0.07fF
C18742 NOR2X1_LOC_155/A INVX1_LOC_270/Y 0.08fF
C18743 NOR2X1_LOC_831/B INVX1_LOC_270/A 0.04fF
C18744 NAND2X1_LOC_443/a_36_24# NOR2X1_LOC_662/A 0.01fF
C18745 NOR2X1_LOC_655/B INVX1_LOC_30/Y 0.05fF
C18746 NOR2X1_LOC_6/B NOR2X1_LOC_99/B 0.08fF
C18747 NAND2X1_LOC_563/A INVX1_LOC_232/A 0.00fF
C18748 NAND2X1_LOC_67/Y NOR2X1_LOC_357/Y 0.58fF
C18749 NOR2X1_LOC_690/A INVX1_LOC_90/A 0.12fF
C18750 NOR2X1_LOC_817/Y NAND2X1_LOC_819/a_36_24# 0.00fF
C18751 NAND2X1_LOC_773/Y VDD 1.39fF
C18752 NOR2X1_LOC_82/A INVX1_LOC_59/Y 0.52fF
C18753 NOR2X1_LOC_82/A INVX1_LOC_112/A 0.01fF
C18754 NAND2X1_LOC_725/A INVX1_LOC_185/A 0.05fF
C18755 INVX1_LOC_103/A INVX1_LOC_139/A 0.01fF
C18756 INVX1_LOC_263/A NAND2X1_LOC_645/a_36_24# 0.02fF
C18757 NOR2X1_LOC_123/B INVX1_LOC_168/A 0.64fF
C18758 INVX1_LOC_78/A INVX1_LOC_125/A 0.07fF
C18759 NOR2X1_LOC_304/Y INVX1_LOC_118/A 0.00fF
C18760 INVX1_LOC_30/A INVX1_LOC_159/Y 0.01fF
C18761 NOR2X1_LOC_392/Y INVX1_LOC_46/Y 0.01fF
C18762 INVX1_LOC_17/A INVX1_LOC_46/A 0.24fF
C18763 INVX1_LOC_269/Y VDD 0.41fF
C18764 NOR2X1_LOC_500/Y INVX1_LOC_220/Y 0.01fF
C18765 NOR2X1_LOC_123/B NAND2X1_LOC_610/a_36_24# 0.01fF
C18766 NOR2X1_LOC_61/B INVX1_LOC_280/A 0.01fF
C18767 INVX1_LOC_2/A INVX1_LOC_89/A 0.48fF
C18768 INVX1_LOC_13/A NOR2X1_LOC_719/A 0.07fF
C18769 NOR2X1_LOC_577/Y NOR2X1_LOC_74/A 0.09fF
C18770 NAND2X1_LOC_778/Y INVX1_LOC_54/A 0.10fF
C18771 INVX1_LOC_201/Y NAND2X1_LOC_293/a_36_24# 0.00fF
C18772 NAND2X1_LOC_714/a_36_24# INVX1_LOC_33/Y 0.00fF
C18773 NAND2X1_LOC_357/B NAND2X1_LOC_807/Y 1.18fF
C18774 INVX1_LOC_135/A NOR2X1_LOC_544/A 0.03fF
C18775 INVX1_LOC_84/A NOR2X1_LOC_696/Y 0.07fF
C18776 INVX1_LOC_252/Y VDD 0.26fF
C18777 INVX1_LOC_230/Y NOR2X1_LOC_825/Y 0.32fF
C18778 NOR2X1_LOC_226/A INVX1_LOC_89/A 0.03fF
C18779 NOR2X1_LOC_831/B NOR2X1_LOC_109/Y 0.02fF
C18780 NOR2X1_LOC_174/B INVX1_LOC_179/Y 0.20fF
C18781 NOR2X1_LOC_383/B INVX1_LOC_19/A 0.13fF
C18782 NOR2X1_LOC_401/B INPUT_1 0.01fF
C18783 NAND2X1_LOC_286/B NAND2X1_LOC_74/B 0.03fF
C18784 NOR2X1_LOC_48/B INVX1_LOC_273/A 0.03fF
C18785 INVX1_LOC_13/Y NAND2X1_LOC_92/a_36_24# 0.01fF
C18786 D_INPUT_0 INVX1_LOC_25/Y 13.91fF
C18787 INVX1_LOC_13/A INVX1_LOC_7/A 0.48fF
C18788 INVX1_LOC_12/A NAND2X1_LOC_99/A 1.24fF
C18789 INVX1_LOC_49/A NOR2X1_LOC_703/Y 0.00fF
C18790 INVX1_LOC_88/A NOR2X1_LOC_331/B 0.10fF
C18791 NOR2X1_LOC_163/Y INVX1_LOC_266/Y 0.02fF
C18792 D_INPUT_0 NAND2X1_LOC_349/B 0.04fF
C18793 NOR2X1_LOC_13/Y NOR2X1_LOC_41/a_36_216# 0.01fF
C18794 NAND2X1_LOC_785/A NOR2X1_LOC_322/Y 0.10fF
C18795 NOR2X1_LOC_15/Y INVX1_LOC_54/A 0.13fF
C18796 NOR2X1_LOC_593/Y INVX1_LOC_206/Y 0.03fF
C18797 NAND2X1_LOC_577/A INVX1_LOC_178/Y 0.05fF
C18798 NOR2X1_LOC_348/B NOR2X1_LOC_74/A 0.05fF
C18799 NAND2X1_LOC_35/Y INVX1_LOC_3/A 0.03fF
C18800 NOR2X1_LOC_794/a_36_216# INVX1_LOC_91/A 0.01fF
C18801 NAND2X1_LOC_303/Y NOR2X1_LOC_51/A 0.03fF
C18802 NAND2X1_LOC_361/a_36_24# NOR2X1_LOC_9/Y 0.00fF
C18803 INVX1_LOC_85/A INVX1_LOC_311/A 0.01fF
C18804 NOR2X1_LOC_356/A NOR2X1_LOC_325/A 0.00fF
C18805 NOR2X1_LOC_356/A INVX1_LOC_22/A 0.08fF
C18806 NOR2X1_LOC_759/A INVX1_LOC_76/A 0.10fF
C18807 INVX1_LOC_224/Y NOR2X1_LOC_76/B 0.02fF
C18808 NAND2X1_LOC_860/A NAND2X1_LOC_74/B 0.09fF
C18809 NOR2X1_LOC_419/Y NAND2X1_LOC_642/Y 0.11fF
C18810 INVX1_LOC_299/A INVX1_LOC_92/A 0.07fF
C18811 NOR2X1_LOC_773/Y NAND2X1_LOC_863/A 0.03fF
C18812 NOR2X1_LOC_589/A D_GATE_366 0.10fF
C18813 NAND2X1_LOC_518/a_36_24# NOR2X1_LOC_557/A 0.00fF
C18814 INVX1_LOC_27/A INVX1_LOC_285/A 0.10fF
C18815 NOR2X1_LOC_598/B INVX1_LOC_69/A 0.03fF
C18816 INPUT_3 INVX1_LOC_9/A 0.03fF
C18817 NOR2X1_LOC_716/B NAND2X1_LOC_642/Y 0.10fF
C18818 NOR2X1_LOC_103/Y NOR2X1_LOC_99/Y 0.07fF
C18819 INVX1_LOC_77/A NOR2X1_LOC_332/B 0.02fF
C18820 NAND2X1_LOC_192/B INVX1_LOC_307/A 0.01fF
C18821 INVX1_LOC_27/A NOR2X1_LOC_814/A 0.68fF
C18822 NAND2X1_LOC_190/Y NOR2X1_LOC_197/B 0.37fF
C18823 NOR2X1_LOC_301/A NOR2X1_LOC_282/a_36_216# 0.00fF
C18824 NOR2X1_LOC_33/A INVX1_LOC_75/A 0.03fF
C18825 NOR2X1_LOC_329/B INVX1_LOC_10/A 0.10fF
C18826 INVX1_LOC_227/A NAND2X1_LOC_123/Y 0.02fF
C18827 NOR2X1_LOC_74/A INVX1_LOC_22/A 0.74fF
C18828 NAND2X1_LOC_352/B INVX1_LOC_131/Y 0.15fF
C18829 INVX1_LOC_89/A INPUT_1 0.13fF
C18830 NOR2X1_LOC_849/A INVX1_LOC_29/A 0.04fF
C18831 INVX1_LOC_255/Y INPUT_0 0.13fF
C18832 NAND2X1_LOC_208/B INVX1_LOC_89/Y 0.04fF
C18833 INVX1_LOC_22/A NOR2X1_LOC_9/Y 0.23fF
C18834 NAND2X1_LOC_640/Y NAND2X1_LOC_633/Y 0.00fF
C18835 NOR2X1_LOC_763/A NOR2X1_LOC_11/Y 0.02fF
C18836 INVX1_LOC_33/A INVX1_LOC_14/Y 0.03fF
C18837 NOR2X1_LOC_355/A INVX1_LOC_73/A 0.15fF
C18838 NOR2X1_LOC_582/A NOR2X1_LOC_11/Y 0.31fF
C18839 INVX1_LOC_98/Y NAND2X1_LOC_642/Y 0.32fF
C18840 NOR2X1_LOC_647/B NAND2X1_LOC_574/A 0.02fF
C18841 D_INPUT_0 INVX1_LOC_75/A 0.15fF
C18842 INVX1_LOC_246/A NOR2X1_LOC_697/Y 0.01fF
C18843 NOR2X1_LOC_366/B NOR2X1_LOC_139/Y 0.03fF
C18844 NAND2X1_LOC_833/Y NOR2X1_LOC_111/A 0.02fF
C18845 INVX1_LOC_18/A INVX1_LOC_274/A 0.07fF
C18846 NAND2X1_LOC_207/Y NAND2X1_LOC_473/A 0.37fF
C18847 NOR2X1_LOC_144/Y VDD 0.11fF
C18848 INVX1_LOC_50/A NOR2X1_LOC_167/a_36_216# 0.00fF
C18849 NOR2X1_LOC_357/Y NOR2X1_LOC_367/B 0.88fF
C18850 NAND2X1_LOC_656/Y NOR2X1_LOC_188/A 0.09fF
C18851 INVX1_LOC_53/A INVX1_LOC_94/Y 0.79fF
C18852 INVX1_LOC_26/Y NOR2X1_LOC_383/B 0.02fF
C18853 NAND2X1_LOC_866/B NAND2X1_LOC_849/A 0.02fF
C18854 INVX1_LOC_278/A NAND2X1_LOC_471/Y 0.01fF
C18855 INVX1_LOC_36/A NOR2X1_LOC_831/B 0.07fF
C18856 NOR2X1_LOC_92/Y NOR2X1_LOC_89/A 1.07fF
C18857 NOR2X1_LOC_373/a_36_216# NAND2X1_LOC_848/A 0.12fF
C18858 INPUT_0 NOR2X1_LOC_71/Y 0.09fF
C18859 INVX1_LOC_230/Y INVX1_LOC_84/A 1.36fF
C18860 INVX1_LOC_236/A INVX1_LOC_76/A 0.01fF
C18861 INVX1_LOC_2/A NAND2X1_LOC_244/A 0.03fF
C18862 D_INPUT_1 INVX1_LOC_26/A 0.81fF
C18863 NOR2X1_LOC_140/A NOR2X1_LOC_847/A 0.03fF
C18864 NOR2X1_LOC_78/A NAND2X1_LOC_41/Y 0.01fF
C18865 NOR2X1_LOC_690/A NAND2X1_LOC_849/B 0.07fF
C18866 INVX1_LOC_94/A NAND2X1_LOC_93/B 0.03fF
C18867 INVX1_LOC_233/A NOR2X1_LOC_301/A 0.07fF
C18868 NOR2X1_LOC_396/a_36_216# NAND2X1_LOC_735/B 0.00fF
C18869 INVX1_LOC_62/A INVX1_LOC_48/A 0.02fF
C18870 INVX1_LOC_5/A NOR2X1_LOC_334/Y 0.08fF
C18871 NOR2X1_LOC_690/A INVX1_LOC_38/A 0.10fF
C18872 NOR2X1_LOC_644/A INPUT_0 0.03fF
C18873 INVX1_LOC_71/A NOR2X1_LOC_99/Y 0.07fF
C18874 NOR2X1_LOC_427/a_36_216# INVX1_LOC_12/A 0.02fF
C18875 NOR2X1_LOC_15/Y NOR2X1_LOC_48/B 0.13fF
C18876 NOR2X1_LOC_802/A INVX1_LOC_117/A 0.07fF
C18877 NAND2X1_LOC_465/Y NOR2X1_LOC_536/A 0.54fF
C18878 NOR2X1_LOC_413/Y INVX1_LOC_38/A 0.17fF
C18879 NOR2X1_LOC_735/Y NOR2X1_LOC_74/A -0.01fF
C18880 NOR2X1_LOC_234/Y NOR2X1_LOC_536/A 0.00fF
C18881 NAND2X1_LOC_538/Y INVX1_LOC_42/A 0.11fF
C18882 NOR2X1_LOC_103/Y NOR2X1_LOC_76/B 0.03fF
C18883 INVX1_LOC_50/A NAND2X1_LOC_787/A 0.03fF
C18884 NAND2X1_LOC_319/a_36_24# NAND2X1_LOC_453/A 0.01fF
C18885 INVX1_LOC_135/A NAND2X1_LOC_655/A 0.10fF
C18886 INVX1_LOC_25/Y NOR2X1_LOC_266/B 0.21fF
C18887 NOR2X1_LOC_637/B NAND2X1_LOC_798/B 0.01fF
C18888 INVX1_LOC_50/A NAND2X1_LOC_363/B 0.02fF
C18889 NAND2X1_LOC_640/Y INVX1_LOC_71/Y 0.01fF
C18890 NOR2X1_LOC_81/a_36_216# NAND2X1_LOC_572/B 0.01fF
C18891 INVX1_LOC_13/A INVX1_LOC_76/A 0.08fF
C18892 NOR2X1_LOC_514/A INVX1_LOC_29/A 0.07fF
C18893 NOR2X1_LOC_387/Y NAND2X1_LOC_810/B 0.57fF
C18894 INVX1_LOC_25/A NOR2X1_LOC_717/A 0.07fF
C18895 INVX1_LOC_119/A INVX1_LOC_118/A 0.61fF
C18896 NOR2X1_LOC_788/B INVX1_LOC_91/A 0.06fF
C18897 NOR2X1_LOC_252/Y INVX1_LOC_46/A 0.16fF
C18898 NAND2X1_LOC_462/B NOR2X1_LOC_24/Y 0.00fF
C18899 INVX1_LOC_16/A INVX1_LOC_37/A 0.03fF
C18900 INVX1_LOC_45/A INVX1_LOC_272/A 0.07fF
C18901 NAND2X1_LOC_350/a_36_24# NAND2X1_LOC_468/B 0.00fF
C18902 NAND2X1_LOC_308/Y INVX1_LOC_185/A 0.00fF
C18903 NOR2X1_LOC_806/Y NOR2X1_LOC_729/A 0.01fF
C18904 NAND2X1_LOC_660/Y NAND2X1_LOC_453/A 0.07fF
C18905 INVX1_LOC_232/A INVX1_LOC_12/Y 1.06fF
C18906 INPUT_3 NOR2X1_LOC_861/Y 0.01fF
C18907 NOR2X1_LOC_781/B NOR2X1_LOC_585/Y 0.03fF
C18908 INVX1_LOC_100/A NOR2X1_LOC_74/A 0.02fF
C18909 INVX1_LOC_96/Y INVX1_LOC_54/A 0.07fF
C18910 NOR2X1_LOC_771/a_36_216# INVX1_LOC_91/A 0.00fF
C18911 NOR2X1_LOC_859/A INVX1_LOC_29/A 0.04fF
C18912 INVX1_LOC_23/A INVX1_LOC_213/A 0.12fF
C18913 INVX1_LOC_279/A VDD 0.76fF
C18914 NOR2X1_LOC_616/a_36_216# NOR2X1_LOC_629/Y 0.00fF
C18915 NOR2X1_LOC_245/a_36_216# INVX1_LOC_20/A 0.00fF
C18916 NOR2X1_LOC_237/a_36_216# NAND2X1_LOC_477/Y 0.01fF
C18917 NAND2X1_LOC_848/A INVX1_LOC_25/Y 0.02fF
C18918 INVX1_LOC_230/Y INVX1_LOC_15/A 0.07fF
C18919 NOR2X1_LOC_246/A INVX1_LOC_76/A 0.10fF
C18920 NOR2X1_LOC_309/Y NOR2X1_LOC_831/B 0.14fF
C18921 INVX1_LOC_266/Y INVX1_LOC_179/A 0.04fF
C18922 NOR2X1_LOC_15/Y NOR2X1_LOC_438/Y 0.07fF
C18923 NOR2X1_LOC_250/A INVX1_LOC_78/A 0.01fF
C18924 INVX1_LOC_9/Y INVX1_LOC_9/A 0.01fF
C18925 INVX1_LOC_41/Y INVX1_LOC_29/A 0.01fF
C18926 NOR2X1_LOC_68/A NAND2X1_LOC_206/B 0.23fF
C18927 INVX1_LOC_71/A INVX1_LOC_272/A 0.03fF
C18928 INVX1_LOC_55/Y INVX1_LOC_76/A 0.07fF
C18929 NOR2X1_LOC_561/Y INVX1_LOC_66/Y 0.01fF
C18930 NOR2X1_LOC_750/A INVX1_LOC_20/A 0.02fF
C18931 INVX1_LOC_1/A NOR2X1_LOC_727/B 0.02fF
C18932 NOR2X1_LOC_160/B NAND2X1_LOC_447/a_36_24# 0.01fF
C18933 NOR2X1_LOC_147/A INVX1_LOC_91/A 0.01fF
C18934 NOR2X1_LOC_791/B INVX1_LOC_3/Y 0.24fF
C18935 NAND2X1_LOC_550/A INVX1_LOC_23/Y 0.08fF
C18936 INVX1_LOC_28/A INVX1_LOC_37/A 0.15fF
C18937 NOR2X1_LOC_65/B NOR2X1_LOC_250/A 0.06fF
C18938 INVX1_LOC_33/A NOR2X1_LOC_831/Y 0.04fF
C18939 NOR2X1_LOC_160/B INVX1_LOC_23/Y 0.07fF
C18940 INVX1_LOC_206/A NOR2X1_LOC_814/A 0.07fF
C18941 INVX1_LOC_268/Y INVX1_LOC_92/A 0.02fF
C18942 INVX1_LOC_182/Y VDD 1.15fF
C18943 INVX1_LOC_50/A NOR2X1_LOC_457/A 0.19fF
C18944 INVX1_LOC_161/Y NOR2X1_LOC_383/B 0.06fF
C18945 NOR2X1_LOC_758/Y INVX1_LOC_29/A 0.01fF
C18946 INVX1_LOC_299/A INVX1_LOC_53/A 0.02fF
C18947 NOR2X1_LOC_312/a_36_216# NOR2X1_LOC_661/A 0.00fF
C18948 INVX1_LOC_1/A NOR2X1_LOC_717/A 0.01fF
C18949 INVX1_LOC_75/A NOR2X1_LOC_266/B 0.03fF
C18950 INVX1_LOC_41/A NOR2X1_LOC_89/A 0.05fF
C18951 NAND2X1_LOC_735/B INVX1_LOC_241/Y 0.01fF
C18952 NAND2X1_LOC_793/Y INVX1_LOC_57/A 0.12fF
C18953 NAND2X1_LOC_803/B INVX1_LOC_271/A 0.02fF
C18954 INVX1_LOC_72/A NOR2X1_LOC_409/B 0.05fF
C18955 NOR2X1_LOC_553/a_36_216# NOR2X1_LOC_383/B 0.00fF
C18956 NOR2X1_LOC_548/Y NOR2X1_LOC_197/B 0.10fF
C18957 NAND2X1_LOC_9/Y INVX1_LOC_17/A 0.02fF
C18958 NOR2X1_LOC_745/Y INVX1_LOC_23/A 0.01fF
C18959 INVX1_LOC_30/A NOR2X1_LOC_306/a_36_216# 0.02fF
C18960 INVX1_LOC_17/A INVX1_LOC_233/A 0.07fF
C18961 NAND2X1_LOC_858/B VDD 0.33fF
C18962 NOR2X1_LOC_590/A INVX1_LOC_271/A 0.07fF
C18963 NAND2X1_LOC_796/B NAND2X1_LOC_784/a_36_24# 0.02fF
C18964 NOR2X1_LOC_423/Y INVX1_LOC_12/A 0.01fF
C18965 NAND2X1_LOC_477/A NOR2X1_LOC_89/A 0.10fF
C18966 NOR2X1_LOC_100/A NOR2X1_LOC_340/A 0.03fF
C18967 INVX1_LOC_277/A NOR2X1_LOC_840/Y 0.01fF
C18968 NOR2X1_LOC_273/Y NAND2X1_LOC_454/Y 0.01fF
C18969 INVX1_LOC_21/A NOR2X1_LOC_454/Y 0.07fF
C18970 INVX1_LOC_56/Y INVX1_LOC_63/A 0.03fF
C18971 NOR2X1_LOC_600/Y NOR2X1_LOC_601/Y 0.06fF
C18972 NOR2X1_LOC_201/A INVX1_LOC_110/A 0.00fF
C18973 NOR2X1_LOC_635/A NOR2X1_LOC_48/B 0.01fF
C18974 INVX1_LOC_136/A NAND2X1_LOC_286/B 0.00fF
C18975 INVX1_LOC_50/A INVX1_LOC_30/A 0.19fF
C18976 NAND2X1_LOC_72/Y NOR2X1_LOC_457/A 0.02fF
C18977 INVX1_LOC_225/Y NOR2X1_LOC_405/Y 0.01fF
C18978 INVX1_LOC_202/A NAND2X1_LOC_454/Y 0.01fF
C18979 NAND2X1_LOC_784/A INVX1_LOC_141/Y 0.03fF
C18980 NOR2X1_LOC_709/A INVX1_LOC_42/A 0.00fF
C18981 NOR2X1_LOC_415/A NAND2X1_LOC_574/A 0.06fF
C18982 INVX1_LOC_135/A NAND2X1_LOC_141/Y 0.90fF
C18983 INVX1_LOC_280/Y NOR2X1_LOC_189/a_36_216# 0.02fF
C18984 NAND2X1_LOC_738/B NOR2X1_LOC_599/A 0.07fF
C18985 NOR2X1_LOC_222/Y INVX1_LOC_12/A 0.72fF
C18986 INVX1_LOC_41/A INVX1_LOC_104/Y 0.01fF
C18987 NAND2X1_LOC_784/A INVX1_LOC_312/Y 0.01fF
C18988 NOR2X1_LOC_83/Y NOR2X1_LOC_536/A 0.16fF
C18989 NOR2X1_LOC_45/B NAND2X1_LOC_254/a_36_24# 0.01fF
C18990 NAND2X1_LOC_549/Y INVX1_LOC_31/A 0.04fF
C18991 INVX1_LOC_17/A NOR2X1_LOC_798/A 1.89fF
C18992 NOR2X1_LOC_403/B INVX1_LOC_26/A 0.04fF
C18993 D_INPUT_2 INVX1_LOC_26/A 0.26fF
C18994 NOR2X1_LOC_145/Y INVX1_LOC_91/A 0.01fF
C18995 NOR2X1_LOC_124/a_36_216# INVX1_LOC_59/Y 0.00fF
C18996 INVX1_LOC_303/A NOR2X1_LOC_621/B 0.04fF
C18997 INVX1_LOC_112/A INVX1_LOC_59/Y 0.01fF
C18998 NAND2X1_LOC_464/Y NAND2X1_LOC_471/Y 0.09fF
C18999 INVX1_LOC_166/A NOR2X1_LOC_480/A 0.50fF
C19000 NOR2X1_LOC_458/Y INVX1_LOC_271/Y 0.03fF
C19001 NOR2X1_LOC_635/A NAND2X1_LOC_3/B 0.02fF
C19002 INVX1_LOC_215/A INVX1_LOC_49/Y 0.06fF
C19003 INVX1_LOC_136/A NOR2X1_LOC_15/a_36_216# 0.00fF
C19004 INVX1_LOC_153/Y INVX1_LOC_271/Y 0.10fF
C19005 NOR2X1_LOC_631/B NOR2X1_LOC_35/Y 0.01fF
C19006 INVX1_LOC_199/Y INVX1_LOC_115/A 0.01fF
C19007 INVX1_LOC_136/A NAND2X1_LOC_860/A 0.07fF
C19008 NOR2X1_LOC_757/Y NAND2X1_LOC_792/B 0.02fF
C19009 NOR2X1_LOC_78/A INVX1_LOC_122/A 0.83fF
C19010 INVX1_LOC_17/A NAND2X1_LOC_703/Y 0.01fF
C19011 INVX1_LOC_136/A NOR2X1_LOC_211/a_36_216# 0.00fF
C19012 NOR2X1_LOC_456/Y NOR2X1_LOC_68/A 0.10fF
C19013 NOR2X1_LOC_160/B NOR2X1_LOC_249/Y 0.33fF
C19014 NAND2X1_LOC_840/B NOR2X1_LOC_48/B 0.08fF
C19015 NOR2X1_LOC_615/Y NOR2X1_LOC_824/A 0.04fF
C19016 NOR2X1_LOC_845/A NOR2X1_LOC_536/A 0.02fF
C19017 INVX1_LOC_289/Y INVX1_LOC_103/A 0.02fF
C19018 INVX1_LOC_11/A NOR2X1_LOC_92/Y 0.09fF
C19019 INVX1_LOC_224/A INVX1_LOC_24/Y 0.00fF
C19020 INVX1_LOC_54/Y NAND2X1_LOC_647/B 0.06fF
C19021 NOR2X1_LOC_772/A INVX1_LOC_285/A 0.02fF
C19022 INVX1_LOC_34/A INVX1_LOC_16/Y 0.00fF
C19023 INVX1_LOC_36/A NAND2X1_LOC_712/a_36_24# 0.00fF
C19024 INPUT_0 NOR2X1_LOC_61/A 0.00fF
C19025 NOR2X1_LOC_357/Y INVX1_LOC_76/A -0.03fF
C19026 NOR2X1_LOC_103/Y NOR2X1_LOC_271/B 0.01fF
C19027 INVX1_LOC_27/A NOR2X1_LOC_590/A 0.12fF
C19028 NOR2X1_LOC_83/Y NAND2X1_LOC_93/B 1.47fF
C19029 INVX1_LOC_67/Y NOR2X1_LOC_216/B 0.01fF
C19030 INVX1_LOC_37/A NOR2X1_LOC_35/Y 0.03fF
C19031 NOR2X1_LOC_709/A INVX1_LOC_78/A 0.12fF
C19032 NOR2X1_LOC_772/A NOR2X1_LOC_814/A 0.01fF
C19033 INVX1_LOC_121/A NOR2X1_LOC_89/A 0.01fF
C19034 INVX1_LOC_27/A INVX1_LOC_22/Y 0.02fF
C19035 NOR2X1_LOC_19/B NOR2X1_LOC_814/A 0.08fF
C19036 NAND2X1_LOC_333/a_36_24# INVX1_LOC_30/A 0.00fF
C19037 INVX1_LOC_89/A NAND2X1_LOC_63/Y 0.12fF
C19038 INVX1_LOC_22/A NAND2X1_LOC_421/a_36_24# 0.00fF
C19039 INVX1_LOC_233/Y NOR2X1_LOC_238/Y 0.06fF
C19040 NOR2X1_LOC_78/B INVX1_LOC_94/Y 0.08fF
C19041 NOR2X1_LOC_334/A NOR2X1_LOC_461/A 0.03fF
C19042 NOR2X1_LOC_719/A INVX1_LOC_32/A 0.02fF
C19043 INVX1_LOC_269/A NOR2X1_LOC_225/a_36_216# 0.12fF
C19044 NOR2X1_LOC_709/B NAND2X1_LOC_642/Y 0.03fF
C19045 INVX1_LOC_34/A NAND2X1_LOC_205/A 0.25fF
C19046 NAND2X1_LOC_338/B NAND2X1_LOC_400/a_36_24# 0.00fF
C19047 NAND2X1_LOC_326/A INVX1_LOC_141/Y 0.02fF
C19048 INVX1_LOC_5/A NAND2X1_LOC_758/a_36_24# 0.00fF
C19049 NOR2X1_LOC_15/Y NOR2X1_LOC_441/Y 0.03fF
C19050 NOR2X1_LOC_790/B NOR2X1_LOC_804/B -0.10fF
C19051 NOR2X1_LOC_65/B NOR2X1_LOC_709/A 0.03fF
C19052 NOR2X1_LOC_833/Y NOR2X1_LOC_499/B 0.01fF
C19053 NOR2X1_LOC_561/Y INVX1_LOC_32/A 0.07fF
C19054 NOR2X1_LOC_332/B INVX1_LOC_9/A 0.05fF
C19055 NOR2X1_LOC_349/A NOR2X1_LOC_259/A 0.09fF
C19056 NOR2X1_LOC_717/a_36_216# NOR2X1_LOC_678/A 0.00fF
C19057 NOR2X1_LOC_292/Y INVX1_LOC_84/A 0.03fF
C19058 INVX1_LOC_7/A INVX1_LOC_32/A 0.22fF
C19059 NAND2X1_LOC_157/a_36_24# INVX1_LOC_53/A 0.00fF
C19060 INVX1_LOC_162/A INVX1_LOC_53/A 0.08fF
C19061 INVX1_LOC_50/A NAND2X1_LOC_722/A 0.09fF
C19062 NOR2X1_LOC_122/Y NOR2X1_LOC_89/A 0.32fF
C19063 NOR2X1_LOC_554/B NAND2X1_LOC_218/A 0.00fF
C19064 NOR2X1_LOC_329/B INVX1_LOC_12/A 0.19fF
C19065 NOR2X1_LOC_96/a_36_216# NOR2X1_LOC_825/Y 0.00fF
C19066 NOR2X1_LOC_140/A NOR2X1_LOC_554/B 0.00fF
C19067 NAND2X1_LOC_860/A NOR2X1_LOC_278/A 0.14fF
C19068 NOR2X1_LOC_74/A INVX1_LOC_186/Y 0.10fF
C19069 NAND2X1_LOC_244/A INVX1_LOC_118/A 0.01fF
C19070 NOR2X1_LOC_516/Y NOR2X1_LOC_660/Y 0.06fF
C19071 VDD NOR2X1_LOC_450/A -0.00fF
C19072 INVX1_LOC_136/A NAND2X1_LOC_537/Y 0.10fF
C19073 INVX1_LOC_89/A INVX1_LOC_257/A 0.00fF
C19074 NOR2X1_LOC_528/Y INVX1_LOC_285/A 0.06fF
C19075 INVX1_LOC_223/Y INVX1_LOC_49/A 0.00fF
C19076 INVX1_LOC_21/A INVX1_LOC_77/A 0.20fF
C19077 NOR2X1_LOC_139/Y NOR2X1_LOC_473/a_36_216# 0.00fF
C19078 NOR2X1_LOC_528/Y INVX1_LOC_265/Y 0.02fF
C19079 INVX1_LOC_20/A INVX1_LOC_70/A 0.03fF
C19080 INVX1_LOC_196/Y INVX1_LOC_15/A 0.08fF
C19081 INVX1_LOC_83/A INVX1_LOC_94/Y 0.01fF
C19082 NAND2X1_LOC_357/B NOR2X1_LOC_109/Y 0.07fF
C19083 INVX1_LOC_178/A INVX1_LOC_209/Y 0.02fF
C19084 NAND2X1_LOC_276/a_36_24# INVX1_LOC_117/A 0.00fF
C19085 INVX1_LOC_2/A NOR2X1_LOC_392/Y 0.00fF
C19086 INVX1_LOC_89/A NAND2X1_LOC_618/Y 0.03fF
C19087 NOR2X1_LOC_92/Y NOR2X1_LOC_433/A 1.56fF
C19088 NOR2X1_LOC_106/A INVX1_LOC_78/A 0.00fF
C19089 VDD NOR2X1_LOC_624/B 0.26fF
C19090 NAND2X1_LOC_392/Y INVX1_LOC_181/A 0.23fF
C19091 INVX1_LOC_161/Y NOR2X1_LOC_512/Y 0.02fF
C19092 NOR2X1_LOC_448/B INVX1_LOC_49/A 0.01fF
C19093 INVX1_LOC_36/A INVX1_LOC_81/Y 0.00fF
C19094 NAND2X1_LOC_538/Y NOR2X1_LOC_152/Y 0.02fF
C19095 INVX1_LOC_256/A INVX1_LOC_94/A 0.10fF
C19096 NOR2X1_LOC_626/Y INVX1_LOC_85/A 0.01fF
C19097 NOR2X1_LOC_45/B NAND2X1_LOC_500/B 0.07fF
C19098 NOR2X1_LOC_290/Y NOR2X1_LOC_291/Y 0.26fF
C19099 INVX1_LOC_34/Y INVX1_LOC_306/Y 0.71fF
C19100 INVX1_LOC_150/Y INVX1_LOC_71/A 0.68fF
C19101 NOR2X1_LOC_250/A NOR2X1_LOC_152/Y 0.03fF
C19102 INVX1_LOC_35/A INVX1_LOC_226/Y 0.03fF
C19103 NOR2X1_LOC_659/a_36_216# INVX1_LOC_30/A 0.00fF
C19104 INVX1_LOC_83/A INVX1_LOC_296/A 0.10fF
C19105 NOR2X1_LOC_250/Y NOR2X1_LOC_577/Y -0.04fF
C19106 NOR2X1_LOC_65/B NOR2X1_LOC_106/A 0.01fF
C19107 NAND2X1_LOC_736/Y INVX1_LOC_229/A 0.03fF
C19108 D_INPUT_1 INVX1_LOC_164/A 0.68fF
C19109 INVX1_LOC_122/Y NAND2X1_LOC_510/A 0.12fF
C19110 INVX1_LOC_269/A NAND2X1_LOC_139/A 0.01fF
C19111 D_INPUT_0 NOR2X1_LOC_529/a_36_216# 0.02fF
C19112 INVX1_LOC_41/A INVX1_LOC_224/A 0.01fF
C19113 NOR2X1_LOC_92/Y NOR2X1_LOC_52/B 0.32fF
C19114 NAND2X1_LOC_2/a_36_24# NAND2X1_LOC_3/B 0.02fF
C19115 NOR2X1_LOC_155/A NOR2X1_LOC_536/A 0.03fF
C19116 NAND2X1_LOC_849/B NOR2X1_LOC_88/a_36_216# 0.00fF
C19117 NOR2X1_LOC_756/a_36_216# INVX1_LOC_23/Y 0.01fF
C19118 INVX1_LOC_41/A INVX1_LOC_11/A 0.06fF
C19119 INVX1_LOC_267/Y INVX1_LOC_235/Y 0.07fF
C19120 NOR2X1_LOC_67/A NAND2X1_LOC_391/Y 0.00fF
C19121 NOR2X1_LOC_20/Y NOR2X1_LOC_413/Y 0.04fF
C19122 NAND2X1_LOC_733/Y NOR2X1_LOC_484/Y 0.01fF
C19123 NAND2X1_LOC_807/Y NOR2X1_LOC_282/Y 0.03fF
C19124 NOR2X1_LOC_226/A NAND2X1_LOC_392/a_36_24# 0.01fF
C19125 NAND2X1_LOC_99/Y NOR2X1_LOC_590/A 0.01fF
C19126 INVX1_LOC_35/A INVX1_LOC_10/A 0.10fF
C19127 INVX1_LOC_144/A NAND2X1_LOC_470/B 0.17fF
C19128 INVX1_LOC_5/A NOR2X1_LOC_569/Y 0.03fF
C19129 NAND2X1_LOC_559/Y NAND2X1_LOC_717/Y 0.05fF
C19130 INVX1_LOC_12/A NOR2X1_LOC_69/A 0.01fF
C19131 INVX1_LOC_229/A INVX1_LOC_282/Y 0.05fF
C19132 NOR2X1_LOC_420/a_36_216# INVX1_LOC_30/Y 0.00fF
C19133 NOR2X1_LOC_655/B NOR2X1_LOC_15/Y 0.01fF
C19134 NOR2X1_LOC_516/B NOR2X1_LOC_846/A 0.01fF
C19135 NAND2X1_LOC_634/Y INVX1_LOC_41/Y 0.00fF
C19136 INVX1_LOC_11/A NAND2X1_LOC_477/A 0.05fF
C19137 INVX1_LOC_105/A INVX1_LOC_30/A 0.99fF
C19138 INVX1_LOC_269/A NOR2X1_LOC_616/a_36_216# 0.00fF
C19139 INVX1_LOC_285/Y INVX1_LOC_271/Y 0.53fF
C19140 NOR2X1_LOC_53/a_36_216# NOR2X1_LOC_53/Y 0.02fF
C19141 INVX1_LOC_21/A NOR2X1_LOC_687/Y 0.43fF
C19142 INVX1_LOC_299/A NOR2X1_LOC_78/B 0.03fF
C19143 NOR2X1_LOC_836/Y NAND2X1_LOC_366/A 0.21fF
C19144 INVX1_LOC_159/A NOR2X1_LOC_596/A 0.18fF
C19145 NOR2X1_LOC_309/Y NAND2X1_LOC_352/B 0.01fF
C19146 INVX1_LOC_102/A INVX1_LOC_20/A 0.07fF
C19147 NOR2X1_LOC_155/A NAND2X1_LOC_93/B 0.03fF
C19148 NOR2X1_LOC_265/a_36_216# NOR2X1_LOC_468/Y 0.03fF
C19149 NOR2X1_LOC_564/Y INVX1_LOC_23/A 0.03fF
C19150 INPUT_1 NOR2X1_LOC_392/Y 0.08fF
C19151 NOR2X1_LOC_510/Y INVX1_LOC_279/A 0.47fF
C19152 NOR2X1_LOC_455/Y INVX1_LOC_55/Y 0.03fF
C19153 INVX1_LOC_139/A NAND2X1_LOC_469/a_36_24# 0.00fF
C19154 NOR2X1_LOC_510/B NAND2X1_LOC_798/B 0.29fF
C19155 INVX1_LOC_88/A NOR2X1_LOC_366/B 0.43fF
C19156 INPUT_0 NOR2X1_LOC_39/Y 0.00fF
C19157 NOR2X1_LOC_68/A NOR2X1_LOC_550/B 0.10fF
C19158 INVX1_LOC_64/A D_GATE_366 0.01fF
C19159 INVX1_LOC_21/A NAND2X1_LOC_796/Y 0.01fF
C19160 INVX1_LOC_13/Y INVX1_LOC_135/A 0.01fF
C19161 NOR2X1_LOC_590/A INVX1_LOC_206/A 0.07fF
C19162 NOR2X1_LOC_311/Y INVX1_LOC_94/Y 0.04fF
C19163 NOR2X1_LOC_434/Y NOR2X1_LOC_174/B 0.20fF
C19164 NOR2X1_LOC_716/B NOR2X1_LOC_91/Y -0.01fF
C19165 INVX1_LOC_293/A NOR2X1_LOC_78/B 0.02fF
C19166 NAND2X1_LOC_1/Y NAND2X1_LOC_429/a_36_24# 0.01fF
C19167 INVX1_LOC_256/A NOR2X1_LOC_136/Y 0.10fF
C19168 INPUT_0 NAND2X1_LOC_205/A 0.06fF
C19169 INVX1_LOC_36/A NAND2X1_LOC_357/B 0.18fF
C19170 INVX1_LOC_32/A INVX1_LOC_76/A 0.60fF
C19171 INVX1_LOC_95/Y INVX1_LOC_4/Y 0.11fF
C19172 INVX1_LOC_284/Y NOR2X1_LOC_822/Y 0.16fF
C19173 D_INPUT_1 NOR2X1_LOC_368/A 0.10fF
C19174 NOR2X1_LOC_331/B INVX1_LOC_272/A 0.04fF
C19175 INVX1_LOC_39/A INVX1_LOC_89/A 0.03fF
C19176 NOR2X1_LOC_250/Y INVX1_LOC_22/A 0.04fF
C19177 INVX1_LOC_2/Y INVX1_LOC_3/Y 0.11fF
C19178 NOR2X1_LOC_294/Y NOR2X1_LOC_87/B 0.07fF
C19179 INVX1_LOC_291/Y INVX1_LOC_273/A 0.37fF
C19180 NOR2X1_LOC_716/B NOR2X1_LOC_81/a_36_216# 0.00fF
C19181 NOR2X1_LOC_216/B INVX1_LOC_285/A 0.10fF
C19182 INVX1_LOC_91/A NAND2X1_LOC_61/Y 0.07fF
C19183 INVX1_LOC_24/A INVX1_LOC_63/Y 0.02fF
C19184 INVX1_LOC_49/Y INVX1_LOC_54/A 0.03fF
C19185 NOR2X1_LOC_361/B INVX1_LOC_279/A -0.02fF
C19186 INVX1_LOC_245/Y INVX1_LOC_22/A 0.03fF
C19187 NOR2X1_LOC_78/A NOR2X1_LOC_621/A 0.01fF
C19188 NOR2X1_LOC_160/B INVX1_LOC_232/A 0.53fF
C19189 NOR2X1_LOC_860/B NOR2X1_LOC_340/Y 0.02fF
C19190 NOR2X1_LOC_216/B NOR2X1_LOC_814/A 0.09fF
C19191 NOR2X1_LOC_134/Y INVX1_LOC_25/Y 0.06fF
C19192 NOR2X1_LOC_188/A NOR2X1_LOC_717/A 0.10fF
C19193 INVX1_LOC_299/A INVX1_LOC_83/A 0.03fF
C19194 NOR2X1_LOC_382/a_36_216# INVX1_LOC_31/A 0.01fF
C19195 VDD NOR2X1_LOC_38/B 1.42fF
C19196 INVX1_LOC_90/A NOR2X1_LOC_376/A 0.01fF
C19197 NOR2X1_LOC_35/Y NAND2X1_LOC_72/B 0.01fF
C19198 INVX1_LOC_157/Y INVX1_LOC_109/A 0.11fF
C19199 NOR2X1_LOC_831/B INVX1_LOC_63/A 1.03fF
C19200 INVX1_LOC_185/A INVX1_LOC_29/A 0.03fF
C19201 INVX1_LOC_41/A NOR2X1_LOC_433/A 0.01fF
C19202 INVX1_LOC_207/Y INVX1_LOC_163/A 0.35fF
C19203 INVX1_LOC_179/A INVX1_LOC_19/A 0.03fF
C19204 NOR2X1_LOC_383/Y NOR2X1_LOC_160/B 0.43fF
C19205 NOR2X1_LOC_52/B NAND2X1_LOC_837/Y 0.07fF
C19206 INVX1_LOC_94/Y INVX1_LOC_46/A 0.16fF
C19207 NAND2X1_LOC_175/Y INVX1_LOC_76/A 0.28fF
C19208 NAND2X1_LOC_741/B NAND2X1_LOC_853/Y 0.03fF
C19209 INVX1_LOC_27/A NOR2X1_LOC_741/a_36_216# 0.01fF
C19210 NAND2X1_LOC_803/B NAND2X1_LOC_156/B 0.35fF
C19211 INVX1_LOC_91/A NOR2X1_LOC_452/A 0.04fF
C19212 NOR2X1_LOC_264/Y NOR2X1_LOC_228/a_36_216# 0.00fF
C19213 NAND2X1_LOC_838/Y NAND2X1_LOC_837/Y 0.06fF
C19214 INVX1_LOC_24/A NOR2X1_LOC_175/A 0.19fF
C19215 INVX1_LOC_90/A INVX1_LOC_14/A 0.75fF
C19216 NOR2X1_LOC_489/A INVX1_LOC_42/A 0.03fF
C19217 INPUT_3 INVX1_LOC_7/A 0.11fF
C19218 INVX1_LOC_239/A INVX1_LOC_135/Y 0.05fF
C19219 NOR2X1_LOC_389/B INVX1_LOC_14/A 0.10fF
C19220 NOR2X1_LOC_433/A NAND2X1_LOC_477/A 0.07fF
C19221 NOR2X1_LOC_777/B NOR2X1_LOC_865/Y 0.15fF
C19222 NOR2X1_LOC_269/Y NOR2X1_LOC_678/A 0.08fF
C19223 NAND2X1_LOC_139/A NAND2X1_LOC_137/a_36_24# 0.02fF
C19224 NOR2X1_LOC_441/Y NAND2X1_LOC_130/a_36_24# 0.00fF
C19225 INVX1_LOC_41/A NOR2X1_LOC_52/B 0.03fF
C19226 NOR2X1_LOC_454/Y NAND2X1_LOC_51/B 0.30fF
C19227 INVX1_LOC_20/A NOR2X1_LOC_280/a_36_216# 0.00fF
C19228 NOR2X1_LOC_307/A INVX1_LOC_85/Y 0.03fF
C19229 NAND2X1_LOC_466/Y NAND2X1_LOC_466/A 0.15fF
C19230 NAND2X1_LOC_785/A NAND2X1_LOC_833/Y 0.07fF
C19231 INVX1_LOC_46/A INVX1_LOC_181/A 0.07fF
C19232 NOR2X1_LOC_276/Y NAND2X1_LOC_128/a_36_24# 0.00fF
C19233 NAND2X1_LOC_198/B INVX1_LOC_16/A 0.01fF
C19234 NAND2X1_LOC_733/Y NOR2X1_LOC_380/A 0.01fF
C19235 NOR2X1_LOC_599/Y NAND2X1_LOC_648/A 0.07fF
C19236 NAND2X1_LOC_348/A INVX1_LOC_14/A 0.06fF
C19237 NOR2X1_LOC_454/Y INVX1_LOC_311/A 0.12fF
C19238 NAND2X1_LOC_357/B NOR2X1_LOC_309/Y 0.00fF
C19239 NOR2X1_LOC_142/Y INVX1_LOC_96/Y 1.05fF
C19240 INVX1_LOC_35/A NOR2X1_LOC_799/B 0.03fF
C19241 NOR2X1_LOC_392/B NOR2X1_LOC_612/B 0.10fF
C19242 INVX1_LOC_238/Y NAND2X1_LOC_866/B 0.17fF
C19243 NOR2X1_LOC_52/B NAND2X1_LOC_477/A 0.01fF
C19244 NAND2X1_LOC_347/B INVX1_LOC_6/A 0.00fF
C19245 NOR2X1_LOC_203/Y NOR2X1_LOC_388/Y 0.13fF
C19246 NOR2X1_LOC_590/A NOR2X1_LOC_772/A 0.05fF
C19247 NAND2X1_LOC_647/B NAND2X1_LOC_656/B 0.15fF
C19248 NOR2X1_LOC_340/Y INVX1_LOC_226/A 0.00fF
C19249 INVX1_LOC_255/Y NOR2X1_LOC_643/Y 0.04fF
C19250 NOR2X1_LOC_817/Y INPUT_0 0.12fF
C19251 NAND2X1_LOC_349/B INVX1_LOC_49/A 0.03fF
C19252 NOR2X1_LOC_593/Y NOR2X1_LOC_211/A 0.33fF
C19253 INVX1_LOC_11/A NAND2X1_LOC_662/B 0.07fF
C19254 NOR2X1_LOC_778/B INVX1_LOC_104/A 0.10fF
C19255 NOR2X1_LOC_664/Y NAND2X1_LOC_819/Y 0.00fF
C19256 NOR2X1_LOC_226/A NAND2X1_LOC_734/B 0.03fF
C19257 NOR2X1_LOC_78/B NOR2X1_LOC_315/Y 0.07fF
C19258 NOR2X1_LOC_644/Y NOR2X1_LOC_648/a_36_216# 0.00fF
C19259 NOR2X1_LOC_577/Y NAND2X1_LOC_660/Y 0.01fF
C19260 INVX1_LOC_89/A INVX1_LOC_61/A 0.04fF
C19261 NOR2X1_LOC_155/A NAND2X1_LOC_470/B 0.04fF
C19262 NAND2X1_LOC_190/Y NOR2X1_LOC_337/Y 0.32fF
C19263 NOR2X1_LOC_793/A INVX1_LOC_186/A 1.00fF
C19264 INVX1_LOC_30/A NAND2X1_LOC_652/Y 0.01fF
C19265 NAND2X1_LOC_725/B NOR2X1_LOC_45/B 0.03fF
C19266 INVX1_LOC_255/Y NOR2X1_LOC_514/a_36_216# 0.01fF
C19267 INVX1_LOC_18/A NOR2X1_LOC_356/A 0.07fF
C19268 NOR2X1_LOC_65/B NOR2X1_LOC_489/A 0.05fF
C19269 NOR2X1_LOC_264/a_36_216# NOR2X1_LOC_78/A 0.00fF
C19270 NOR2X1_LOC_432/Y NOR2X1_LOC_78/B 0.01fF
C19271 NOR2X1_LOC_516/B NAND2X1_LOC_116/A 0.01fF
C19272 INVX1_LOC_269/A NOR2X1_LOC_78/A 0.11fF
C19273 NOR2X1_LOC_48/B INVX1_LOC_49/Y 0.19fF
C19274 INVX1_LOC_303/A INVX1_LOC_135/A 0.09fF
C19275 NOR2X1_LOC_15/Y INVX1_LOC_291/Y 0.03fF
C19276 D_INPUT_0 NOR2X1_LOC_577/Y 0.01fF
C19277 INVX1_LOC_279/A INVX1_LOC_153/Y 0.02fF
C19278 NOR2X1_LOC_589/A INVX1_LOC_162/Y 0.15fF
C19279 NOR2X1_LOC_420/Y VDD 0.23fF
C19280 NAND2X1_LOC_84/Y INVX1_LOC_90/A 0.48fF
C19281 NAND2X1_LOC_198/B INVX1_LOC_28/A 0.10fF
C19282 INVX1_LOC_305/A NOR2X1_LOC_567/B 0.01fF
C19283 NOR2X1_LOC_609/a_36_216# INVX1_LOC_313/Y 0.00fF
C19284 NAND2X1_LOC_84/Y NOR2X1_LOC_389/B 0.01fF
C19285 INVX1_LOC_5/A NAND2X1_LOC_472/Y 0.07fF
C19286 NOR2X1_LOC_615/a_36_216# INVX1_LOC_91/A 0.02fF
C19287 NAND2X1_LOC_364/A INVX1_LOC_73/A 0.03fF
C19288 INVX1_LOC_230/Y INVX1_LOC_123/A 0.14fF
C19289 NAND2X1_LOC_541/Y NAND2X1_LOC_563/A 0.11fF
C19290 NAND2X1_LOC_725/A NOR2X1_LOC_536/A 1.69fF
C19291 NAND2X1_LOC_33/Y NAND2X1_LOC_462/B 0.02fF
C19292 INVX1_LOC_63/Y NOR2X1_LOC_130/A 0.13fF
C19293 INVX1_LOC_2/A NAND2X1_LOC_349/B 0.00fF
C19294 NOR2X1_LOC_123/B NAND2X1_LOC_494/a_36_24# 0.00fF
C19295 NOR2X1_LOC_647/A NOR2X1_LOC_820/Y 0.11fF
C19296 NOR2X1_LOC_808/A NOR2X1_LOC_374/B 0.03fF
C19297 NOR2X1_LOC_226/A INVX1_LOC_25/Y 0.08fF
C19298 NOR2X1_LOC_160/B INVX1_LOC_186/A 0.01fF
C19299 NAND2X1_LOC_659/A INVX1_LOC_175/A 0.02fF
C19300 NAND2X1_LOC_288/A NAND2X1_LOC_288/B 0.02fF
C19301 NOR2X1_LOC_222/Y D_GATE_222 0.01fF
C19302 INVX1_LOC_18/A NOR2X1_LOC_74/A 0.34fF
C19303 INVX1_LOC_57/A NAND2X1_LOC_798/B 0.07fF
C19304 NOR2X1_LOC_433/A NOR2X1_LOC_122/Y 0.05fF
C19305 INVX1_LOC_215/A NAND2X1_LOC_231/Y 0.10fF
C19306 INVX1_LOC_237/Y INVX1_LOC_207/Y 0.50fF
C19307 NOR2X1_LOC_624/A INVX1_LOC_89/A 0.00fF
C19308 NOR2X1_LOC_843/B NOR2X1_LOC_243/B 0.07fF
C19309 INVX1_LOC_277/A INVX1_LOC_78/Y 0.00fF
C19310 INVX1_LOC_279/A INVX1_LOC_177/A 0.02fF
C19311 NOR2X1_LOC_392/B NOR2X1_LOC_137/A 0.73fF
C19312 INVX1_LOC_227/A INVX1_LOC_206/A 0.01fF
C19313 NOR2X1_LOC_242/A NAND2X1_LOC_96/A 0.07fF
C19314 NOR2X1_LOC_299/Y NAND2X1_LOC_838/Y 0.02fF
C19315 NOR2X1_LOC_598/B NAND2X1_LOC_93/B 0.07fF
C19316 INVX1_LOC_36/A NAND2X1_LOC_473/a_36_24# 0.00fF
C19317 NOR2X1_LOC_468/Y VDD 1.81fF
C19318 INVX1_LOC_62/Y NOR2X1_LOC_721/Y 0.03fF
C19319 INVX1_LOC_299/A INVX1_LOC_46/A 0.23fF
C19320 INVX1_LOC_18/A NOR2X1_LOC_9/Y 0.28fF
C19321 NOR2X1_LOC_703/B NOR2X1_LOC_551/Y 0.02fF
C19322 INVX1_LOC_209/Y INVX1_LOC_140/A 0.03fF
C19323 NAND2X1_LOC_190/Y VDD 0.39fF
C19324 NOR2X1_LOC_383/B NOR2X1_LOC_801/A 0.01fF
C19325 INVX1_LOC_5/A NAND2X1_LOC_637/Y 0.03fF
C19326 INVX1_LOC_134/A INVX1_LOC_143/Y 0.05fF
C19327 INVX1_LOC_289/A INVX1_LOC_290/A 0.01fF
C19328 NOR2X1_LOC_65/B INVX1_LOC_294/A 0.01fF
C19329 INVX1_LOC_310/A INVX1_LOC_83/A 0.07fF
C19330 INVX1_LOC_35/A INVX1_LOC_307/A 0.07fF
C19331 INVX1_LOC_77/A NAND2X1_LOC_51/B 0.11fF
C19332 INVX1_LOC_49/A INVX1_LOC_75/A 5.82fF
C19333 INVX1_LOC_248/A NAND2X1_LOC_796/Y 0.01fF
C19334 NAND2X1_LOC_727/Y INVX1_LOC_22/A 0.01fF
C19335 NOR2X1_LOC_15/Y NOR2X1_LOC_176/Y 0.10fF
C19336 NOR2X1_LOC_160/B NAND2X1_LOC_447/Y 0.67fF
C19337 NOR2X1_LOC_100/A INVX1_LOC_120/A 0.02fF
C19338 INVX1_LOC_194/A INVX1_LOC_175/Y 0.27fF
C19339 NAND2X1_LOC_538/a_36_24# NOR2X1_LOC_577/Y 0.00fF
C19340 INVX1_LOC_21/A INVX1_LOC_9/A 2.13fF
C19341 INVX1_LOC_209/Y NAND2X1_LOC_463/B 0.06fF
C19342 INVX1_LOC_172/A NOR2X1_LOC_74/A 0.03fF
C19343 INVX1_LOC_182/Y INVX1_LOC_153/Y 0.00fF
C19344 INVX1_LOC_69/Y INVX1_LOC_94/A 0.17fF
C19345 INVX1_LOC_90/A NOR2X1_LOC_612/B 0.02fF
C19346 NOR2X1_LOC_665/A INVX1_LOC_16/A 0.03fF
C19347 NOR2X1_LOC_552/A NOR2X1_LOC_500/B 0.00fF
C19348 NOR2X1_LOC_376/A INVX1_LOC_38/A 0.01fF
C19349 INVX1_LOC_35/A NOR2X1_LOC_445/B 0.03fF
C19350 D_INPUT_0 NOR2X1_LOC_346/B 0.03fF
C19351 NOR2X1_LOC_334/Y INVX1_LOC_42/A 0.07fF
C19352 NAND2X1_LOC_288/B INVX1_LOC_19/A 0.02fF
C19353 NOR2X1_LOC_644/A INVX1_LOC_266/Y 0.08fF
C19354 INVX1_LOC_77/A INVX1_LOC_311/A 0.01fF
C19355 NOR2X1_LOC_589/A NAND2X1_LOC_662/Y 0.07fF
C19356 INVX1_LOC_111/Y NOR2X1_LOC_355/a_36_216# 0.00fF
C19357 NAND2X1_LOC_123/Y INVX1_LOC_104/A 0.08fF
C19358 INVX1_LOC_208/A NOR2X1_LOC_366/Y 0.00fF
C19359 INVX1_LOC_88/A NOR2X1_LOC_152/A 0.31fF
C19360 INVX1_LOC_14/A NOR2X1_LOC_561/A 0.16fF
C19361 NAND2X1_LOC_334/a_36_24# NOR2X1_LOC_71/Y 0.00fF
C19362 INVX1_LOC_219/A INVX1_LOC_316/Y 0.01fF
C19363 INVX1_LOC_246/A INVX1_LOC_37/A 0.85fF
C19364 NOR2X1_LOC_598/B INVX1_LOC_3/A 0.09fF
C19365 NOR2X1_LOC_389/A VDD 2.65fF
C19366 D_INPUT_0 INVX1_LOC_22/A 0.07fF
C19367 NOR2X1_LOC_790/B INVX1_LOC_63/A 0.07fF
C19368 INVX1_LOC_182/Y INVX1_LOC_177/A 0.02fF
C19369 NOR2X1_LOC_552/A NOR2X1_LOC_170/a_36_216# 0.01fF
C19370 NAND2X1_LOC_199/B VDD 0.01fF
C19371 INVX1_LOC_222/A INVX1_LOC_149/Y 0.06fF
C19372 NOR2X1_LOC_13/Y NOR2X1_LOC_43/Y 0.34fF
C19373 INVX1_LOC_25/Y INPUT_1 0.24fF
C19374 INVX1_LOC_2/A INVX1_LOC_75/A 0.13fF
C19375 INVX1_LOC_34/A INVX1_LOC_286/A 0.07fF
C19376 NOR2X1_LOC_753/Y INVX1_LOC_91/A 0.07fF
C19377 INVX1_LOC_133/Y INVX1_LOC_79/A 0.10fF
C19378 NOR2X1_LOC_97/B NOR2X1_LOC_99/B 0.03fF
C19379 INVX1_LOC_5/A NAND2X1_LOC_206/Y 0.07fF
C19380 INVX1_LOC_19/A NOR2X1_LOC_405/Y 0.01fF
C19381 NOR2X1_LOC_226/A INVX1_LOC_75/A 0.08fF
C19382 INVX1_LOC_28/A INVX1_LOC_53/Y 0.01fF
C19383 INVX1_LOC_93/A INVX1_LOC_265/Y 0.01fF
C19384 NAND2X1_LOC_464/B INVX1_LOC_42/A 0.02fF
C19385 NAND2X1_LOC_325/Y INVX1_LOC_91/A 0.09fF
C19386 NOR2X1_LOC_595/a_36_216# INVX1_LOC_38/A 0.00fF
C19387 INVX1_LOC_78/A NOR2X1_LOC_334/Y 0.14fF
C19388 NOR2X1_LOC_91/Y NAND2X1_LOC_633/Y 0.16fF
C19389 NOR2X1_LOC_753/Y INVX1_LOC_11/Y 0.14fF
C19390 NAND2X1_LOC_192/B INVX1_LOC_92/A 0.01fF
C19391 NOR2X1_LOC_250/A INVX1_LOC_291/A 0.18fF
C19392 INVX1_LOC_28/A NOR2X1_LOC_665/A 0.19fF
C19393 INVX1_LOC_62/Y VDD 0.70fF
C19394 INVX1_LOC_35/A INVX1_LOC_12/A 0.10fF
C19395 INVX1_LOC_213/A INVX1_LOC_301/A 0.03fF
C19396 NAND2X1_LOC_324/a_36_24# NOR2X1_LOC_841/A 0.07fF
C19397 INVX1_LOC_2/A NOR2X1_LOC_7/a_36_216# 0.03fF
C19398 NOR2X1_LOC_596/A VDD 0.22fF
C19399 NOR2X1_LOC_447/A NOR2X1_LOC_329/Y 0.01fF
C19400 NOR2X1_LOC_207/a_36_216# NOR2X1_LOC_214/B 0.03fF
C19401 NOR2X1_LOC_562/A NOR2X1_LOC_303/Y 0.02fF
C19402 INVX1_LOC_47/Y INVX1_LOC_57/A 0.10fF
C19403 NOR2X1_LOC_67/A INVX1_LOC_309/A -0.01fF
C19404 INVX1_LOC_145/Y INVX1_LOC_28/A 0.01fF
C19405 INVX1_LOC_64/A INVX1_LOC_102/A 0.07fF
C19406 INVX1_LOC_256/A NOR2X1_LOC_155/A 2.09fF
C19407 NOR2X1_LOC_778/B INVX1_LOC_206/Y 0.01fF
C19408 INVX1_LOC_88/A NOR2X1_LOC_473/a_36_216# 0.00fF
C19409 NAND2X1_LOC_222/B NAND2X1_LOC_574/A 0.02fF
C19410 NOR2X1_LOC_148/A NOR2X1_LOC_148/Y 0.01fF
C19411 INVX1_LOC_49/A NAND2X1_LOC_453/A 0.05fF
C19412 NOR2X1_LOC_350/A INVX1_LOC_37/A 0.01fF
C19413 NOR2X1_LOC_113/B INVX1_LOC_16/A 0.02fF
C19414 NOR2X1_LOC_329/B NAND2X1_LOC_808/A 0.00fF
C19415 INVX1_LOC_201/Y INVX1_LOC_74/A 0.07fF
C19416 NAND2X1_LOC_339/a_36_24# NAND2X1_LOC_468/B 0.00fF
C19417 NOR2X1_LOC_455/Y INVX1_LOC_32/A 0.02fF
C19418 NOR2X1_LOC_577/Y NOR2X1_LOC_682/Y 0.14fF
C19419 NOR2X1_LOC_67/A INVX1_LOC_91/A 0.15fF
C19420 INVX1_LOC_11/A NOR2X1_LOC_435/B 0.03fF
C19421 NOR2X1_LOC_315/Y NOR2X1_LOC_368/Y 0.06fF
C19422 NOR2X1_LOC_590/A NOR2X1_LOC_216/B 0.03fF
C19423 NAND2X1_LOC_721/B INVX1_LOC_185/A 0.00fF
C19424 NOR2X1_LOC_712/Y VDD 0.18fF
C19425 NOR2X1_LOC_778/B NOR2X1_LOC_600/Y 0.01fF
C19426 NAND2X1_LOC_231/Y INVX1_LOC_95/A 0.18fF
C19427 NOR2X1_LOC_488/Y NOR2X1_LOC_528/Y 0.01fF
C19428 NOR2X1_LOC_763/A INPUT_7 0.04fF
C19429 NOR2X1_LOC_550/a_36_216# NOR2X1_LOC_197/B 0.13fF
C19430 INVX1_LOC_27/A NOR2X1_LOC_67/Y 0.02fF
C19431 NOR2X1_LOC_582/A INPUT_7 0.02fF
C19432 NOR2X1_LOC_295/Y VDD 0.49fF
C19433 NAND2X1_LOC_673/a_36_24# NAND2X1_LOC_721/A 0.00fF
C19434 INVX1_LOC_279/A INVX1_LOC_285/Y 0.10fF
C19435 NOR2X1_LOC_392/Y NAND2X1_LOC_618/Y 0.12fF
C19436 INVX1_LOC_64/A NOR2X1_LOC_329/a_36_216# 0.01fF
C19437 NAND2X1_LOC_147/a_36_24# INVX1_LOC_76/A 0.00fF
C19438 NOR2X1_LOC_316/Y INVX1_LOC_20/A 0.01fF
C19439 NOR2X1_LOC_598/B NAND2X1_LOC_470/B 0.02fF
C19440 NOR2X1_LOC_299/Y INVX1_LOC_140/Y 0.08fF
C19441 INVX1_LOC_314/Y NOR2X1_LOC_119/a_36_216# 0.01fF
C19442 NOR2X1_LOC_577/Y NAND2X1_LOC_848/A 0.15fF
C19443 NOR2X1_LOC_844/A VDD 0.12fF
C19444 NOR2X1_LOC_337/Y NOR2X1_LOC_548/Y 0.01fF
C19445 INVX1_LOC_21/A NOR2X1_LOC_861/Y 0.07fF
C19446 INVX1_LOC_75/A INPUT_1 0.33fF
C19447 NOR2X1_LOC_315/Y INVX1_LOC_46/A 0.07fF
C19448 NOR2X1_LOC_434/Y NOR2X1_LOC_623/B 0.03fF
C19449 NAND2X1_LOC_352/B INVX1_LOC_63/A 0.98fF
C19450 NOR2X1_LOC_672/Y INVX1_LOC_280/A 0.05fF
C19451 NOR2X1_LOC_92/Y NAND2X1_LOC_254/Y 0.03fF
C19452 INVX1_LOC_245/Y INVX1_LOC_186/Y 0.00fF
C19453 INVX1_LOC_71/A NOR2X1_LOC_612/Y 0.19fF
C19454 INVX1_LOC_2/A NAND2X1_LOC_453/A 0.03fF
C19455 NAND2X1_LOC_656/A INVX1_LOC_92/A 0.04fF
C19456 NOR2X1_LOC_226/A NAND2X1_LOC_453/A 0.14fF
C19457 INVX1_LOC_189/Y VDD 0.41fF
C19458 NOR2X1_LOC_356/A NOR2X1_LOC_548/A 0.02fF
C19459 NOR2X1_LOC_758/Y INVX1_LOC_118/Y 0.02fF
C19460 NOR2X1_LOC_399/Y VDD 0.12fF
C19461 NOR2X1_LOC_389/A INVX1_LOC_133/A 0.08fF
C19462 INVX1_LOC_279/A INVX1_LOC_65/A 0.30fF
C19463 INVX1_LOC_90/A INVX1_LOC_48/A 0.03fF
C19464 NOR2X1_LOC_220/A VDD 2.41fF
C19465 NOR2X1_LOC_383/B NOR2X1_LOC_493/a_36_216# 0.00fF
C19466 INVX1_LOC_233/A INVX1_LOC_181/A 0.58fF
C19467 NOR2X1_LOC_619/A NOR2X1_LOC_35/Y 0.07fF
C19468 INVX1_LOC_34/A INVX1_LOC_54/A 0.24fF
C19469 NOR2X1_LOC_441/Y INVX1_LOC_49/Y 0.25fF
C19470 NAND2X1_LOC_735/B NOR2X1_LOC_24/Y 0.03fF
C19471 NOR2X1_LOC_641/B INVX1_LOC_19/A 0.03fF
C19472 NAND2X1_LOC_390/A INVX1_LOC_126/A 0.04fF
C19473 NAND2X1_LOC_541/Y INVX1_LOC_12/Y 0.02fF
C19474 NAND2X1_LOC_660/A NOR2X1_LOC_536/A 0.10fF
C19475 INVX1_LOC_41/A NOR2X1_LOC_676/a_36_216# 0.01fF
C19476 NOR2X1_LOC_547/B NAND2X1_LOC_96/A 0.04fF
C19477 INVX1_LOC_22/A NOR2X1_LOC_266/B 0.01fF
C19478 NOR2X1_LOC_78/B NAND2X1_LOC_96/A 1.44fF
C19479 INVX1_LOC_105/A INVX1_LOC_113/A 0.08fF
C19480 VDD NAND2X1_LOC_863/B 0.25fF
C19481 INVX1_LOC_182/Y INVX1_LOC_285/Y 0.03fF
C19482 INVX1_LOC_27/A NOR2X1_LOC_415/Y 0.01fF
C19483 NAND2X1_LOC_773/Y INVX1_LOC_4/Y 0.10fF
C19484 NOR2X1_LOC_751/Y INVX1_LOC_19/A 0.03fF
C19485 NAND2X1_LOC_708/Y NOR2X1_LOC_696/a_36_216# 0.00fF
C19486 NAND2X1_LOC_347/B NOR2X1_LOC_80/Y 0.01fF
C19487 VDD NOR2X1_LOC_548/Y 0.22fF
C19488 INVX1_LOC_290/A INVX1_LOC_37/A 0.03fF
C19489 INVX1_LOC_212/A NOR2X1_LOC_814/A 0.06fF
C19490 NOR2X1_LOC_361/B NOR2X1_LOC_38/B 0.01fF
C19491 INVX1_LOC_217/Y NAND2X1_LOC_848/Y 0.00fF
C19492 NOR2X1_LOC_706/Y INVX1_LOC_75/A 0.01fF
C19493 INVX1_LOC_166/A INVX1_LOC_253/Y 0.17fF
C19494 NAND2X1_LOC_832/Y INVX1_LOC_311/A 0.01fF
C19495 NOR2X1_LOC_655/B NAND2X1_LOC_204/a_36_24# 0.06fF
C19496 NOR2X1_LOC_835/A INVX1_LOC_117/A 0.01fF
C19497 INVX1_LOC_89/A NAND2X1_LOC_212/Y 0.02fF
C19498 NOR2X1_LOC_254/A INVX1_LOC_15/A 0.07fF
C19499 NAND2X1_LOC_231/Y INVX1_LOC_54/A 0.01fF
C19500 INVX1_LOC_138/A NOR2X1_LOC_392/Y 0.02fF
C19501 VDD NAND2X1_LOC_795/Y 0.03fF
C19502 NOR2X1_LOC_205/Y INVX1_LOC_271/Y 0.07fF
C19503 NOR2X1_LOC_68/A NAND2X1_LOC_74/B 1.92fF
C19504 INPUT_5 NOR2X1_LOC_425/Y 0.05fF
C19505 NOR2X1_LOC_423/Y INVX1_LOC_92/A 0.58fF
C19506 INVX1_LOC_286/A INPUT_0 0.27fF
C19507 INPUT_2 INVX1_LOC_4/A 0.09fF
C19508 INVX1_LOC_120/A INVX1_LOC_176/A 0.04fF
C19509 INVX1_LOC_66/A INVX1_LOC_46/A 0.13fF
C19510 INVX1_LOC_16/A NOR2X1_LOC_652/a_36_216# 0.00fF
C19511 NAND2X1_LOC_198/B INVX1_LOC_109/A 0.03fF
C19512 NOR2X1_LOC_355/B NOR2X1_LOC_335/B 0.25fF
C19513 INVX1_LOC_89/A D_INPUT_3 0.03fF
C19514 INVX1_LOC_73/A NOR2X1_LOC_405/A 3.85fF
C19515 NOR2X1_LOC_175/A NOR2X1_LOC_197/B 0.64fF
C19516 INVX1_LOC_25/Y INVX1_LOC_118/A 11.18fF
C19517 INVX1_LOC_28/A NAND2X1_LOC_465/A 0.01fF
C19518 INVX1_LOC_89/A INVX1_LOC_14/Y 1.13fF
C19519 NAND2X1_LOC_345/a_36_24# INVX1_LOC_14/Y 0.00fF
C19520 INVX1_LOC_94/A NOR2X1_LOC_89/A 0.07fF
C19521 NOR2X1_LOC_222/Y INVX1_LOC_92/A 1.04fF
C19522 NOR2X1_LOC_346/B INVX1_LOC_46/Y 0.07fF
C19523 INVX1_LOC_83/A NAND2X1_LOC_96/A 0.07fF
C19524 NOR2X1_LOC_518/a_36_216# NOR2X1_LOC_48/B 0.00fF
C19525 NOR2X1_LOC_391/A NOR2X1_LOC_271/Y 0.03fF
C19526 NOR2X1_LOC_276/Y NAND2X1_LOC_454/Y -0.02fF
C19527 INVX1_LOC_39/A NOR2X1_LOC_392/Y 0.01fF
C19528 INVX1_LOC_144/Y NOR2X1_LOC_88/Y 0.00fF
C19529 NOR2X1_LOC_544/A NOR2X1_LOC_862/B 0.01fF
C19530 NAND2X1_LOC_357/B NOR2X1_LOC_654/a_36_216# 0.00fF
C19531 INVX1_LOC_223/A INVX1_LOC_4/A 0.03fF
C19532 INVX1_LOC_95/A INPUT_0 0.10fF
C19533 NAND2X1_LOC_357/B INVX1_LOC_63/A 0.07fF
C19534 INVX1_LOC_54/Y INVX1_LOC_285/A 0.23fF
C19535 INVX1_LOC_305/Y NOR2X1_LOC_445/B 0.00fF
C19536 NOR2X1_LOC_82/Y NOR2X1_LOC_216/B 0.01fF
C19537 INVX1_LOC_54/Y NOR2X1_LOC_814/A 0.05fF
C19538 NOR2X1_LOC_666/A NOR2X1_LOC_678/A 0.01fF
C19539 INVX1_LOC_72/A NOR2X1_LOC_158/B 0.00fF
C19540 INVX1_LOC_94/A NOR2X1_LOC_170/A 0.11fF
C19541 INVX1_LOC_209/Y INVX1_LOC_42/A 0.00fF
C19542 INVX1_LOC_1/Y NOR2X1_LOC_831/B 1.09fF
C19543 INVX1_LOC_77/A NOR2X1_LOC_865/a_36_216# 0.00fF
C19544 INVX1_LOC_49/A INVX1_LOC_283/A 0.00fF
C19545 NOR2X1_LOC_45/B NAND2X1_LOC_655/A 0.45fF
C19546 NOR2X1_LOC_67/A INVX1_LOC_203/A 0.10fF
C19547 NOR2X1_LOC_365/a_36_216# INVX1_LOC_12/A 0.02fF
C19548 NOR2X1_LOC_641/B INVX1_LOC_26/Y 0.00fF
C19549 INVX1_LOC_31/A NOR2X1_LOC_646/B 0.01fF
C19550 INVX1_LOC_34/A NOR2X1_LOC_48/B 0.10fF
C19551 D_INPUT_0 NOR2X1_LOC_88/A 0.01fF
C19552 INVX1_LOC_157/A NOR2X1_LOC_155/A 0.00fF
C19553 INVX1_LOC_256/A NOR2X1_LOC_598/B 0.07fF
C19554 INVX1_LOC_36/A NOR2X1_LOC_282/Y 0.01fF
C19555 NAND2X1_LOC_560/A NOR2X1_LOC_536/A 0.04fF
C19556 NAND2X1_LOC_303/Y NOR2X1_LOC_304/Y 0.02fF
C19557 INVX1_LOC_230/Y D_INPUT_1 0.15fF
C19558 INVX1_LOC_51/Y VDD 0.85fF
C19559 NOR2X1_LOC_45/B NAND2X1_LOC_468/B 0.03fF
C19560 INVX1_LOC_141/Y NOR2X1_LOC_654/A 0.03fF
C19561 INVX1_LOC_135/A NOR2X1_LOC_861/a_36_216# 0.00fF
C19562 NOR2X1_LOC_751/Y INVX1_LOC_26/Y 0.06fF
C19563 NOR2X1_LOC_152/Y NOR2X1_LOC_334/Y 0.15fF
C19564 INVX1_LOC_312/Y NOR2X1_LOC_654/A 0.00fF
C19565 NOR2X1_LOC_186/Y INVX1_LOC_269/A 0.03fF
C19566 INVX1_LOC_299/A NOR2X1_LOC_798/A 0.06fF
C19567 NAND2X1_LOC_45/Y NOR2X1_LOC_259/B 0.07fF
C19568 NOR2X1_LOC_366/B INVX1_LOC_272/A 0.15fF
C19569 INVX1_LOC_100/Y VDD 0.41fF
C19570 NAND2X1_LOC_231/Y NAND2X1_LOC_807/B 0.04fF
C19571 NOR2X1_LOC_538/B NOR2X1_LOC_798/A 0.02fF
C19572 INVX1_LOC_75/A INVX1_LOC_118/A 0.07fF
C19573 INVX1_LOC_209/Y INVX1_LOC_78/A 0.03fF
C19574 INVX1_LOC_255/Y INVX1_LOC_19/A 0.03fF
C19575 INVX1_LOC_2/A INVX1_LOC_283/A 0.03fF
C19576 NAND2X1_LOC_793/Y INVX1_LOC_306/Y 0.01fF
C19577 NAND2X1_LOC_850/Y INVX1_LOC_102/A 0.03fF
C19578 NOR2X1_LOC_136/Y NOR2X1_LOC_89/A 0.07fF
C19579 NOR2X1_LOC_56/Y NAND2X1_LOC_469/B 0.02fF
C19580 NOR2X1_LOC_128/B INVX1_LOC_63/A 0.03fF
C19581 INVX1_LOC_85/A INVX1_LOC_4/A 0.01fF
C19582 INVX1_LOC_272/Y NAND2X1_LOC_714/B 0.10fF
C19583 NOR2X1_LOC_15/Y NAND2X1_LOC_579/A 0.03fF
C19584 INVX1_LOC_99/Y NOR2X1_LOC_590/A 0.03fF
C19585 NAND2X1_LOC_555/Y NOR2X1_LOC_663/A 0.02fF
C19586 INVX1_LOC_311/A INVX1_LOC_9/A 0.03fF
C19587 NOR2X1_LOC_78/A INVX1_LOC_12/Y 0.05fF
C19588 INPUT_0 INVX1_LOC_54/A 0.10fF
C19589 INVX1_LOC_48/A INVX1_LOC_38/A 0.02fF
C19590 NOR2X1_LOC_316/Y INVX1_LOC_4/A 0.01fF
C19591 NOR2X1_LOC_468/Y NOR2X1_LOC_361/B 0.10fF
C19592 INVX1_LOC_259/Y NOR2X1_LOC_68/A 0.02fF
C19593 NOR2X1_LOC_602/A NOR2X1_LOC_109/Y 0.11fF
C19594 INVX1_LOC_132/A NOR2X1_LOC_621/A 0.02fF
C19595 NOR2X1_LOC_718/B INVX1_LOC_78/A 0.03fF
C19596 INVX1_LOC_21/A NOR2X1_LOC_331/Y 0.05fF
C19597 NOR2X1_LOC_808/A NOR2X1_LOC_801/B 0.03fF
C19598 NOR2X1_LOC_447/B NOR2X1_LOC_56/Y 0.02fF
C19599 VDD NAND2X1_LOC_655/B 0.07fF
C19600 INVX1_LOC_289/Y NOR2X1_LOC_533/Y 0.00fF
C19601 INVX1_LOC_124/A NOR2X1_LOC_248/A 0.04fF
C19602 VDD NAND2X1_LOC_469/B 0.40fF
C19603 NOR2X1_LOC_75/a_36_216# NOR2X1_LOC_158/Y 0.00fF
C19604 NOR2X1_LOC_322/Y NOR2X1_LOC_88/Y 0.07fF
C19605 NAND2X1_LOC_569/A INVX1_LOC_23/Y 0.02fF
C19606 NOR2X1_LOC_276/B NOR2X1_LOC_678/A 0.01fF
C19607 INVX1_LOC_279/A NOR2X1_LOC_830/Y 0.03fF
C19608 NOR2X1_LOC_71/Y INVX1_LOC_19/A 0.08fF
C19609 INVX1_LOC_22/A NOR2X1_LOC_754/A 0.00fF
C19610 NOR2X1_LOC_454/Y INVX1_LOC_174/A 0.12fF
C19611 INVX1_LOC_201/A NOR2X1_LOC_655/Y 0.02fF
C19612 INVX1_LOC_135/A INVX1_LOC_272/A 0.04fF
C19613 NOR2X1_LOC_110/a_36_216# NOR2X1_LOC_831/Y 0.01fF
C19614 NAND2X1_LOC_510/A INVX1_LOC_50/Y 0.18fF
C19615 NOR2X1_LOC_608/a_36_216# NOR2X1_LOC_38/B 0.00fF
C19616 NOR2X1_LOC_772/Y NOR2X1_LOC_383/B 0.03fF
C19617 NOR2X1_LOC_710/a_36_216# NOR2X1_LOC_155/A 0.00fF
C19618 NAND2X1_LOC_783/Y NAND2X1_LOC_780/Y 0.04fF
C19619 NOR2X1_LOC_309/Y NOR2X1_LOC_282/Y 0.03fF
C19620 INVX1_LOC_140/A NAND2X1_LOC_30/a_36_24# 0.01fF
C19621 INVX1_LOC_268/A D_INPUT_5 0.03fF
C19622 INVX1_LOC_21/A NOR2X1_LOC_565/A 0.03fF
C19623 VDD NOR2X1_LOC_447/B 0.27fF
C19624 NOR2X1_LOC_644/A INVX1_LOC_19/A 0.04fF
C19625 INVX1_LOC_21/A NOR2X1_LOC_169/B 0.02fF
C19626 NOR2X1_LOC_188/A NAND2X1_LOC_85/Y 0.03fF
C19627 NOR2X1_LOC_322/Y INVX1_LOC_84/A 0.08fF
C19628 INVX1_LOC_34/A NAND2X1_LOC_215/A 0.23fF
C19629 NOR2X1_LOC_392/B NOR2X1_LOC_383/B 0.02fF
C19630 INVX1_LOC_284/Y NAND2X1_LOC_493/Y 0.24fF
C19631 NOR2X1_LOC_791/B NOR2X1_LOC_791/Y 0.08fF
C19632 NOR2X1_LOC_361/B NOR2X1_LOC_389/A 0.10fF
C19633 INVX1_LOC_5/A INVX1_LOC_24/A 5.47fF
C19634 INVX1_LOC_27/A INVX1_LOC_177/Y 0.03fF
C19635 NOR2X1_LOC_828/B INVX1_LOC_19/A 0.23fF
C19636 INVX1_LOC_36/A NAND2X1_LOC_347/B 0.04fF
C19637 NAND2X1_LOC_96/A NOR2X1_LOC_98/A 0.00fF
C19638 NOR2X1_LOC_191/A INVX1_LOC_26/A 0.02fF
C19639 NOR2X1_LOC_78/B NAND2X1_LOC_99/A 0.07fF
C19640 INVX1_LOC_122/Y NOR2X1_LOC_227/B 0.03fF
C19641 NAND2X1_LOC_9/Y NOR2X1_LOC_350/a_36_216# 0.01fF
C19642 INVX1_LOC_201/A NOR2X1_LOC_649/B 0.10fF
C19643 INVX1_LOC_178/A INVX1_LOC_24/A 0.06fF
C19644 NOR2X1_LOC_195/A INVX1_LOC_31/A 0.01fF
C19645 INVX1_LOC_58/A NOR2X1_LOC_361/Y 0.01fF
C19646 INVX1_LOC_201/A INVX1_LOC_3/A 0.01fF
C19647 NOR2X1_LOC_32/B NOR2X1_LOC_6/B 0.33fF
C19648 NOR2X1_LOC_569/Y INVX1_LOC_78/A 0.43fF
C19649 INVX1_LOC_182/A INVX1_LOC_99/A 0.09fF
C19650 NAND2X1_LOC_9/Y NOR2X1_LOC_315/Y 0.03fF
C19651 NAND2X1_LOC_453/A INVX1_LOC_118/A 0.96fF
C19652 NAND2X1_LOC_387/a_36_24# INVX1_LOC_174/A 0.01fF
C19653 INVX1_LOC_17/A INVX1_LOC_72/A 0.10fF
C19654 NOR2X1_LOC_355/B INVX1_LOC_84/A 0.20fF
C19655 INVX1_LOC_233/A NOR2X1_LOC_315/Y 0.00fF
C19656 NAND2X1_LOC_86/Y NOR2X1_LOC_243/B 0.04fF
C19657 NOR2X1_LOC_93/a_36_216# NOR2X1_LOC_392/Y 0.01fF
C19658 NOR2X1_LOC_366/B NOR2X1_LOC_125/a_36_216# 0.00fF
C19659 NOR2X1_LOC_168/B INVX1_LOC_58/Y 0.07fF
C19660 INVX1_LOC_45/Y NOR2X1_LOC_122/A 0.01fF
C19661 NOR2X1_LOC_599/Y NOR2X1_LOC_761/a_36_216# 0.01fF
C19662 NOR2X1_LOC_13/Y NAND2X1_LOC_326/A 0.23fF
C19663 NAND2X1_LOC_35/Y NOR2X1_LOC_52/B 0.07fF
C19664 INVX1_LOC_126/Y INVX1_LOC_29/A 0.04fF
C19665 NAND2X1_LOC_35/Y NAND2X1_LOC_838/Y 0.02fF
C19666 INPUT_0 NAND2X1_LOC_807/B 0.05fF
C19667 NOR2X1_LOC_328/Y INVX1_LOC_57/A 0.05fF
C19668 NOR2X1_LOC_720/B INVX1_LOC_50/Y 0.04fF
C19669 INVX1_LOC_245/Y INVX1_LOC_18/A 0.03fF
C19670 INVX1_LOC_130/A INVX1_LOC_30/A 0.04fF
C19671 NAND2X1_LOC_553/A NOR2X1_LOC_315/Y 0.01fF
C19672 NOR2X1_LOC_273/Y NAND2X1_LOC_53/Y 0.15fF
C19673 INVX1_LOC_251/Y NOR2X1_LOC_772/B 0.00fF
C19674 NAND2X1_LOC_574/A INVX1_LOC_74/A 0.01fF
C19675 NAND2X1_LOC_567/Y NAND2X1_LOC_537/Y 0.00fF
C19676 INVX1_LOC_11/A INVX1_LOC_94/A 0.01fF
C19677 NOR2X1_LOC_523/A INVX1_LOC_77/A -0.01fF
C19678 INVX1_LOC_45/Y INVX1_LOC_161/Y 0.18fF
C19679 INPUT_0 NOR2X1_LOC_48/B 0.19fF
C19680 INVX1_LOC_27/A INVX1_LOC_104/A 0.07fF
C19681 INVX1_LOC_21/A NOR2X1_LOC_61/a_36_216# 0.02fF
C19682 INVX1_LOC_24/A NOR2X1_LOC_816/A 0.10fF
C19683 INVX1_LOC_5/A INVX1_LOC_143/A 0.07fF
C19684 D_INPUT_0 NOR2X1_LOC_843/B 0.03fF
C19685 INVX1_LOC_251/Y INVX1_LOC_13/Y 1.73fF
C19686 NOR2X1_LOC_441/Y INVX1_LOC_79/Y 0.13fF
C19687 NOR2X1_LOC_481/A INVX1_LOC_269/A 0.09fF
C19688 INVX1_LOC_14/A INVX1_LOC_33/A 0.53fF
C19689 NOR2X1_LOC_91/A NOR2X1_LOC_246/A 0.10fF
C19690 NAND2X1_LOC_16/a_36_24# INVX1_LOC_72/A 0.01fF
C19691 NOR2X1_LOC_829/a_36_216# NAND2X1_LOC_738/B 0.00fF
C19692 NAND2X1_LOC_53/Y NOR2X1_LOC_550/B 0.10fF
C19693 INVX1_LOC_291/Y INVX1_LOC_49/Y 0.03fF
C19694 NAND2X1_LOC_190/Y INVX1_LOC_153/Y 0.02fF
C19695 INVX1_LOC_230/Y D_INPUT_2 0.27fF
C19696 INVX1_LOC_220/Y INVX1_LOC_53/A 0.00fF
C19697 NAND2X1_LOC_763/B D_INPUT_7 0.01fF
C19698 INVX1_LOC_5/A INVX1_LOC_68/Y 0.01fF
C19699 INVX1_LOC_64/A NOR2X1_LOC_94/a_36_216# 0.00fF
C19700 INVX1_LOC_174/A INVX1_LOC_77/A 0.78fF
C19701 INVX1_LOC_225/A INVX1_LOC_269/A 0.10fF
C19702 INVX1_LOC_21/A INVX1_LOC_243/A 0.00fF
C19703 NOR2X1_LOC_590/A NOR2X1_LOC_303/Y 0.03fF
C19704 INVX1_LOC_209/Y NOR2X1_LOC_503/Y 2.52fF
C19705 INVX1_LOC_64/A NAND2X1_LOC_662/Y 0.01fF
C19706 NAND2X1_LOC_140/A INVX1_LOC_270/Y 0.02fF
C19707 NOR2X1_LOC_861/a_36_216# INVX1_LOC_280/A 0.01fF
C19708 INVX1_LOC_159/A NAND2X1_LOC_154/Y 0.01fF
C19709 NOR2X1_LOC_272/Y NAND2X1_LOC_181/Y 0.03fF
C19710 INVX1_LOC_90/A NOR2X1_LOC_383/B 0.06fF
C19711 INVX1_LOC_136/A NOR2X1_LOC_68/A 0.17fF
C19712 NAND2X1_LOC_551/a_36_24# NOR2X1_LOC_71/Y 0.01fF
C19713 NOR2X1_LOC_246/A INVX1_LOC_23/A 0.07fF
C19714 NOR2X1_LOC_86/Y INVX1_LOC_61/A 0.02fF
C19715 NOR2X1_LOC_389/B NOR2X1_LOC_383/B 0.07fF
C19716 INVX1_LOC_225/Y NOR2X1_LOC_570/B 0.05fF
C19717 NAND2X1_LOC_552/a_36_24# NAND2X1_LOC_552/A 0.00fF
C19718 NOR2X1_LOC_363/Y NAND2X1_LOC_475/Y 0.10fF
C19719 NAND2X1_LOC_53/Y INVX1_LOC_249/Y 0.01fF
C19720 INVX1_LOC_272/Y NAND2X1_LOC_802/a_36_24# 0.01fF
C19721 INVX1_LOC_81/A INVX1_LOC_30/A 0.46fF
C19722 NAND2X1_LOC_190/Y INVX1_LOC_177/A 0.15fF
C19723 INVX1_LOC_39/A INVX1_LOC_25/Y 0.09fF
C19724 NOR2X1_LOC_808/A INVX1_LOC_1/A 0.03fF
C19725 NOR2X1_LOC_588/A D_INPUT_5 0.03fF
C19726 NOR2X1_LOC_778/B INVX1_LOC_24/Y 0.02fF
C19727 NOR2X1_LOC_590/A NOR2X1_LOC_254/Y 0.03fF
C19728 NOR2X1_LOC_435/a_36_216# NOR2X1_LOC_130/A 0.00fF
C19729 INVX1_LOC_38/A NOR2X1_LOC_127/Y 0.07fF
C19730 NOR2X1_LOC_536/A NOR2X1_LOC_673/B 0.01fF
C19731 INVX1_LOC_6/A NOR2X1_LOC_158/Y 0.02fF
C19732 INVX1_LOC_58/A NOR2X1_LOC_736/Y 0.07fF
C19733 NOR2X1_LOC_751/A INVX1_LOC_26/Y 0.03fF
C19734 NOR2X1_LOC_852/A NAND2X1_LOC_364/Y 0.04fF
C19735 INVX1_LOC_48/A NAND2X1_LOC_223/A 0.07fF
C19736 INVX1_LOC_17/A NOR2X1_LOC_537/Y 0.03fF
C19737 NAND2X1_LOC_149/Y INVX1_LOC_16/A 0.14fF
C19738 INVX1_LOC_33/A NOR2X1_LOC_717/Y 0.01fF
C19739 NAND2X1_LOC_579/A NAND2X1_LOC_840/B 0.01fF
C19740 INVX1_LOC_17/A NAND2X1_LOC_338/B 0.07fF
C19741 NOR2X1_LOC_479/B NOR2X1_LOC_475/A 0.09fF
C19742 INVX1_LOC_37/A NAND2X1_LOC_245/a_36_24# 0.00fF
C19743 INVX1_LOC_37/A INVX1_LOC_261/Y 0.03fF
C19744 INVX1_LOC_255/Y NOR2X1_LOC_474/a_36_216# 0.01fF
C19745 NOR2X1_LOC_468/a_36_216# NOR2X1_LOC_652/Y 0.00fF
C19746 INVX1_LOC_5/A NOR2X1_LOC_130/A 0.01fF
C19747 NOR2X1_LOC_448/Y INVX1_LOC_22/A 0.02fF
C19748 INVX1_LOC_14/A INVX1_LOC_40/A 0.67fF
C19749 INVX1_LOC_21/A NOR2X1_LOC_561/Y 0.08fF
C19750 INVX1_LOC_37/A NOR2X1_LOC_641/a_36_216# 0.00fF
C19751 INVX1_LOC_230/Y NOR2X1_LOC_529/Y 0.05fF
C19752 INVX1_LOC_37/A INVX1_LOC_114/Y 0.02fF
C19753 NOR2X1_LOC_454/Y NOR2X1_LOC_589/A 0.06fF
C19754 NOR2X1_LOC_329/B INVX1_LOC_53/A 0.64fF
C19755 NOR2X1_LOC_437/Y INVX1_LOC_45/Y 0.03fF
C19756 NOR2X1_LOC_620/Y NAND2X1_LOC_364/A 0.02fF
C19757 NAND2X1_LOC_482/a_36_24# INVX1_LOC_213/A 0.00fF
C19758 NAND2X1_LOC_533/a_36_24# NOR2X1_LOC_356/A 0.00fF
C19759 INVX1_LOC_233/A NOR2X1_LOC_166/Y 0.03fF
C19760 NAND2X1_LOC_350/A NAND2X1_LOC_231/Y 0.10fF
C19761 INVX1_LOC_229/A INVX1_LOC_22/A 0.23fF
C19762 NAND2X1_LOC_577/A INVX1_LOC_80/Y 0.01fF
C19763 NAND2X1_LOC_714/B INVX1_LOC_10/A 0.02fF
C19764 D_INPUT_4 INVX1_LOC_53/A 0.02fF
C19765 NOR2X1_LOC_590/A INVX1_LOC_54/Y 0.05fF
C19766 INPUT_0 NAND2X1_LOC_215/A 0.12fF
C19767 INVX1_LOC_236/A INVX1_LOC_31/A 0.13fF
C19768 NOR2X1_LOC_536/A INVX1_LOC_29/A 1.00fF
C19769 NOR2X1_LOC_802/A INVX1_LOC_30/A 0.02fF
C19770 INVX1_LOC_159/A INVX1_LOC_63/Y 0.00fF
C19771 NOR2X1_LOC_82/A INVX1_LOC_56/Y 0.06fF
C19772 NAND2X1_LOC_231/Y NOR2X1_LOC_441/Y 0.03fF
C19773 INVX1_LOC_278/A NOR2X1_LOC_322/Y 0.10fF
C19774 NOR2X1_LOC_593/Y INVX1_LOC_94/A 0.07fF
C19775 NAND2X1_LOC_30/Y INVX1_LOC_22/A 0.24fF
C19776 NAND2X1_LOC_472/Y INVX1_LOC_42/A 0.09fF
C19777 NAND2X1_LOC_656/B NOR2X1_LOC_814/A 0.02fF
C19778 NOR2X1_LOC_596/A INVX1_LOC_153/Y 0.10fF
C19779 INVX1_LOC_279/A NOR2X1_LOC_205/Y 0.02fF
C19780 INVX1_LOC_37/A NOR2X1_LOC_467/A 0.33fF
C19781 INVX1_LOC_49/A NOR2X1_LOC_577/Y 0.07fF
C19782 INVX1_LOC_41/A INVX1_LOC_314/Y 0.74fF
C19783 NAND2X1_LOC_361/Y NAND2X1_LOC_7/Y 0.03fF
C19784 INVX1_LOC_2/A NOR2X1_LOC_274/B 0.01fF
C19785 NAND2X1_LOC_579/A NOR2X1_LOC_576/B 0.63fF
C19786 NAND2X1_LOC_352/B INVX1_LOC_1/Y 0.08fF
C19787 NOR2X1_LOC_791/A INVX1_LOC_34/Y -0.01fF
C19788 NOR2X1_LOC_655/Y INVX1_LOC_29/A 0.03fF
C19789 NOR2X1_LOC_598/B INVX1_LOC_69/Y 0.00fF
C19790 NAND2X1_LOC_198/B NOR2X1_LOC_84/Y 0.28fF
C19791 NAND2X1_LOC_364/Y NOR2X1_LOC_285/B 0.02fF
C19792 NAND2X1_LOC_93/B INVX1_LOC_29/A 0.04fF
C19793 NOR2X1_LOC_614/Y NOR2X1_LOC_500/B 0.03fF
C19794 INVX1_LOC_2/A NOR2X1_LOC_351/a_36_216# 0.00fF
C19795 INVX1_LOC_13/A INVX1_LOC_31/A 0.30fF
C19796 NOR2X1_LOC_596/A INVX1_LOC_177/A 0.03fF
C19797 INVX1_LOC_39/A INVX1_LOC_75/A 0.03fF
C19798 NAND2X1_LOC_783/A NOR2X1_LOC_816/A 0.34fF
C19799 NOR2X1_LOC_718/B INVX1_LOC_113/Y 0.03fF
C19800 NAND2X1_LOC_337/B NOR2X1_LOC_130/A 0.07fF
C19801 INVX1_LOC_34/A NOR2X1_LOC_142/Y 0.15fF
C19802 NOR2X1_LOC_292/Y NOR2X1_LOC_652/Y 0.01fF
C19803 NAND2X1_LOC_860/A INVX1_LOC_70/Y 0.04fF
C19804 NOR2X1_LOC_518/Y NOR2X1_LOC_165/Y 0.11fF
C19805 NOR2X1_LOC_98/B INVX1_LOC_4/Y 0.03fF
C19806 NOR2X1_LOC_89/A NOR2X1_LOC_155/A 0.06fF
C19807 INVX1_LOC_78/A NAND2X1_LOC_472/Y 0.09fF
C19808 NOR2X1_LOC_589/A NAND2X1_LOC_196/a_36_24# 0.00fF
C19809 INVX1_LOC_41/A NOR2X1_LOC_181/Y 0.13fF
C19810 NOR2X1_LOC_92/Y NOR2X1_LOC_597/Y 0.01fF
C19811 INVX1_LOC_24/A NOR2X1_LOC_773/Y 0.07fF
C19812 INVX1_LOC_272/A NOR2X1_LOC_473/a_36_216# 0.01fF
C19813 INVX1_LOC_46/A NAND2X1_LOC_99/A 0.08fF
C19814 INVX1_LOC_61/A INVX1_LOC_25/Y 0.08fF
C19815 INVX1_LOC_2/A NOR2X1_LOC_577/Y 0.25fF
C19816 NOR2X1_LOC_220/B INVX1_LOC_286/A 0.02fF
C19817 INVX1_LOC_21/A NOR2X1_LOC_167/Y 0.03fF
C19818 NOR2X1_LOC_477/B INVX1_LOC_92/A 0.02fF
C19819 NOR2X1_LOC_205/Y INVX1_LOC_182/Y 0.02fF
C19820 NOR2X1_LOC_720/B NOR2X1_LOC_6/B 0.35fF
C19821 NOR2X1_LOC_649/B INVX1_LOC_29/A 0.07fF
C19822 INVX1_LOC_18/A NAND2X1_LOC_660/Y 0.06fF
C19823 NOR2X1_LOC_226/A NOR2X1_LOC_577/Y 0.10fF
C19824 INVX1_LOC_3/A INVX1_LOC_29/A 0.13fF
C19825 INVX1_LOC_27/A INVX1_LOC_206/Y 0.08fF
C19826 INVX1_LOC_249/A INVX1_LOC_263/A 0.03fF
C19827 NOR2X1_LOC_357/Y INVX1_LOC_23/A 0.07fF
C19828 INVX1_LOC_13/Y NOR2X1_LOC_45/B 0.10fF
C19829 NOR2X1_LOC_655/B INVX1_LOC_34/A 0.01fF
C19830 NOR2X1_LOC_67/A NAND2X1_LOC_276/Y 0.07fF
C19831 INVX1_LOC_41/A NOR2X1_LOC_778/B 0.03fF
C19832 INVX1_LOC_206/A INVX1_LOC_104/A 0.02fF
C19833 NOR2X1_LOC_500/Y NOR2X1_LOC_550/B 0.03fF
C19834 NAND2X1_LOC_736/Y NAND2X1_LOC_733/B 0.85fF
C19835 NOR2X1_LOC_532/Y INVX1_LOC_30/A 0.04fF
C19836 NOR2X1_LOC_773/Y NOR2X1_LOC_557/Y 0.12fF
C19837 INVX1_LOC_49/A NOR2X1_LOC_325/A 0.12fF
C19838 INVX1_LOC_2/A NOR2X1_LOC_348/B 0.03fF
C19839 NAND2X1_LOC_740/Y NAND2X1_LOC_729/B 0.03fF
C19840 INVX1_LOC_58/A NOR2X1_LOC_111/A 0.00fF
C19841 INVX1_LOC_49/A INVX1_LOC_22/A 7.38fF
C19842 INVX1_LOC_11/A INVX1_LOC_144/A 0.07fF
C19843 NAND2X1_LOC_206/Y INVX1_LOC_42/A 0.02fF
C19844 NOR2X1_LOC_609/A NAND2X1_LOC_656/Y 0.02fF
C19845 INVX1_LOC_33/Y INVX1_LOC_57/A 0.03fF
C19846 NAND2X1_LOC_563/Y NAND2X1_LOC_578/B 0.03fF
C19847 INVX1_LOC_85/A INVX1_LOC_44/Y 0.05fF
C19848 INVX1_LOC_162/Y NAND2X1_LOC_850/Y 0.01fF
C19849 NOR2X1_LOC_589/A INVX1_LOC_77/A 3.86fF
C19850 NOR2X1_LOC_74/A NAND2X1_LOC_793/Y 0.01fF
C19851 D_INPUT_3 NOR2X1_LOC_392/Y 0.19fF
C19852 NOR2X1_LOC_759/Y INVX1_LOC_10/A 0.35fF
C19853 NOR2X1_LOC_469/a_36_216# NOR2X1_LOC_167/Y 0.00fF
C19854 NOR2X1_LOC_726/Y NOR2X1_LOC_738/A 0.17fF
C19855 INVX1_LOC_38/A NOR2X1_LOC_383/B 0.24fF
C19856 INVX1_LOC_310/Y NAND2X1_LOC_282/a_36_24# 0.00fF
C19857 INVX1_LOC_202/A INVX1_LOC_10/A 0.07fF
C19858 INVX1_LOC_83/A NAND2X1_LOC_656/A 0.33fF
C19859 NOR2X1_LOC_78/B NOR2X1_LOC_423/Y 0.02fF
C19860 INVX1_LOC_42/A NAND2X1_LOC_773/B 0.05fF
C19861 NOR2X1_LOC_136/Y NOR2X1_LOC_52/B 0.06fF
C19862 NOR2X1_LOC_388/Y NOR2X1_LOC_563/a_36_216# 0.00fF
C19863 NOR2X1_LOC_361/B INVX1_LOC_100/Y 0.03fF
C19864 INVX1_LOC_47/A NOR2X1_LOC_360/Y 0.11fF
C19865 NOR2X1_LOC_401/a_36_216# NOR2X1_LOC_84/Y 0.00fF
C19866 INVX1_LOC_282/Y NAND2X1_LOC_733/B 2.20fF
C19867 NOR2X1_LOC_510/Y NAND2X1_LOC_469/B 0.00fF
C19868 NAND2X1_LOC_9/Y NAND2X1_LOC_96/A 0.03fF
C19869 NOR2X1_LOC_220/A INVX1_LOC_177/A 0.01fF
C19870 INVX1_LOC_90/A NOR2X1_LOC_512/Y 0.04fF
C19871 INVX1_LOC_88/A NOR2X1_LOC_45/B 0.06fF
C19872 NAND2X1_LOC_206/a_36_24# NAND2X1_LOC_348/A 0.01fF
C19873 INVX1_LOC_93/A NAND2X1_LOC_650/B 0.02fF
C19874 NOR2X1_LOC_441/Y INPUT_0 0.17fF
C19875 INVX1_LOC_21/A INVX1_LOC_76/A 0.23fF
C19876 INVX1_LOC_254/A INVX1_LOC_89/A 0.22fF
C19877 INVX1_LOC_171/A INVX1_LOC_77/A 0.04fF
C19878 NOR2X1_LOC_222/Y NOR2X1_LOC_78/B 0.03fF
C19879 INVX1_LOC_269/A NAND2X1_LOC_642/Y 0.10fF
C19880 NOR2X1_LOC_392/Y INVX1_LOC_230/A 0.01fF
C19881 INVX1_LOC_119/Y INVX1_LOC_94/Y 0.00fF
C19882 NOR2X1_LOC_510/Y NOR2X1_LOC_447/B 0.00fF
C19883 INVX1_LOC_136/A INVX1_LOC_147/A 0.01fF
C19884 INVX1_LOC_103/A NOR2X1_LOC_141/a_36_216# 0.00fF
C19885 INVX1_LOC_2/A INVX1_LOC_22/A 0.87fF
C19886 NOR2X1_LOC_496/Y VDD 0.33fF
C19887 NOR2X1_LOC_577/Y NAND2X1_LOC_648/A 0.02fF
C19888 NAND2X1_LOC_363/B NAND2X1_LOC_276/a_36_24# 0.00fF
C19889 NOR2X1_LOC_186/Y INVX1_LOC_12/Y 0.01fF
C19890 NOR2X1_LOC_160/B INVX1_LOC_98/A 0.00fF
C19891 INVX1_LOC_177/A NOR2X1_LOC_548/Y 0.00fF
C19892 NOR2X1_LOC_748/Y NOR2X1_LOC_538/Y 0.02fF
C19893 INVX1_LOC_24/A INVX1_LOC_140/A 0.22fF
C19894 INVX1_LOC_268/A NAND2X1_LOC_451/Y 0.05fF
C19895 NOR2X1_LOC_500/A NOR2X1_LOC_703/A 0.05fF
C19896 NOR2X1_LOC_226/A INVX1_LOC_22/A 2.71fF
C19897 NOR2X1_LOC_160/B NOR2X1_LOC_78/A 2.77fF
C19898 NOR2X1_LOC_690/A INVX1_LOC_89/A 0.04fF
C19899 NAND2X1_LOC_557/a_36_24# NOR2X1_LOC_536/A 0.00fF
C19900 INVX1_LOC_52/Y VDD -0.00fF
C19901 NOR2X1_LOC_550/a_36_216# NOR2X1_LOC_337/Y 0.03fF
C19902 NAND2X1_LOC_81/B NOR2X1_LOC_38/B 0.01fF
C19903 INVX1_LOC_41/A NOR2X1_LOC_724/Y 0.03fF
C19904 NAND2X1_LOC_286/B INVX1_LOC_285/A 0.01fF
C19905 NOR2X1_LOC_861/Y NOR2X1_LOC_865/a_36_216# 0.00fF
C19906 NOR2X1_LOC_41/Y INVX1_LOC_10/A 0.06fF
C19907 NOR2X1_LOC_456/Y INVX1_LOC_307/A 0.18fF
C19908 NOR2X1_LOC_289/Y NAND2X1_LOC_593/Y 0.16fF
C19909 NOR2X1_LOC_340/A NOR2X1_LOC_227/A 0.24fF
C19910 NAND2X1_LOC_222/a_36_24# NOR2X1_LOC_673/A 0.02fF
C19911 INVX1_LOC_1/A INVX1_LOC_37/A 0.31fF
C19912 INVX1_LOC_161/A INVX1_LOC_291/Y 0.01fF
C19913 NOR2X1_LOC_804/B NOR2X1_LOC_564/Y 0.01fF
C19914 INVX1_LOC_1/A NOR2X1_LOC_231/A 0.01fF
C19915 NOR2X1_LOC_662/A INVX1_LOC_23/Y 0.01fF
C19916 NOR2X1_LOC_759/A INVX1_LOC_6/A 0.13fF
C19917 INVX1_LOC_124/A INVX1_LOC_171/A 0.02fF
C19918 NOR2X1_LOC_219/Y INVX1_LOC_290/A 0.10fF
C19919 INVX1_LOC_25/Y NOR2X1_LOC_85/a_36_216# 0.00fF
C19920 INVX1_LOC_35/A INVX1_LOC_92/A 0.06fF
C19921 NAND2X1_LOC_470/B INVX1_LOC_29/A 0.08fF
C19922 NOR2X1_LOC_191/A INVX1_LOC_164/A 0.00fF
C19923 NOR2X1_LOC_393/Y INVX1_LOC_42/A 0.02fF
C19924 INVX1_LOC_290/Y INVX1_LOC_4/A 0.07fF
C19925 NAND2X1_LOC_218/a_36_24# NOR2X1_LOC_814/A 0.01fF
C19926 NOR2X1_LOC_297/A INVX1_LOC_42/A 0.02fF
C19927 NAND2X1_LOC_213/A INVX1_LOC_117/A 0.01fF
C19928 INVX1_LOC_135/A NOR2X1_LOC_87/Y 0.01fF
C19929 INVX1_LOC_280/Y NAND2X1_LOC_795/Y 0.05fF
C19930 NOR2X1_LOC_596/A INVX1_LOC_285/Y 0.03fF
C19931 INVX1_LOC_27/A NOR2X1_LOC_119/a_36_216# 0.01fF
C19932 NOR2X1_LOC_433/A INVX1_LOC_144/A 0.22fF
C19933 NOR2X1_LOC_757/Y NAND2X1_LOC_656/Y 0.23fF
C19934 NOR2X1_LOC_222/Y INVX1_LOC_83/A 0.10fF
C19935 INVX1_LOC_77/A INVX1_LOC_222/A 0.01fF
C19936 NOR2X1_LOC_15/a_36_216# INVX1_LOC_285/A 0.00fF
C19937 NOR2X1_LOC_39/Y INVX1_LOC_19/A 0.12fF
C19938 NOR2X1_LOC_773/Y NOR2X1_LOC_130/A 0.38fF
C19939 INVX1_LOC_314/Y NOR2X1_LOC_71/a_36_216# 0.00fF
C19940 NAND2X1_LOC_721/a_36_24# INVX1_LOC_28/A 0.01fF
C19941 NOR2X1_LOC_332/A INVX1_LOC_68/Y 0.03fF
C19942 INVX1_LOC_262/Y NOR2X1_LOC_635/B 0.01fF
C19943 NOR2X1_LOC_560/A NOR2X1_LOC_87/Y 0.01fF
C19944 INVX1_LOC_292/A NOR2X1_LOC_137/Y 0.38fF
C19945 NOR2X1_LOC_794/B INVX1_LOC_37/A 0.04fF
C19946 INVX1_LOC_181/Y INVX1_LOC_91/A 0.01fF
C19947 INVX1_LOC_5/A NOR2X1_LOC_197/B 0.04fF
C19948 NOR2X1_LOC_781/B INVX1_LOC_290/A 0.05fF
C19949 NOR2X1_LOC_340/Y INPUT_0 0.05fF
C19950 INVX1_LOC_2/A NOR2X1_LOC_735/Y 0.01fF
C19951 INVX1_LOC_269/A NOR2X1_LOC_271/Y 0.03fF
C19952 NAND2X1_LOC_175/B NOR2X1_LOC_815/A 0.02fF
C19953 INVX1_LOC_253/A INVX1_LOC_3/Y 0.02fF
C19954 NOR2X1_LOC_433/a_36_216# NAND2X1_LOC_832/Y 0.00fF
C19955 INVX1_LOC_151/A INVX1_LOC_144/A 0.04fF
C19956 NOR2X1_LOC_52/Y NAND2X1_LOC_468/B 0.00fF
C19957 INVX1_LOC_1/A NAND2X1_LOC_629/a_36_24# 0.00fF
C19958 NOR2X1_LOC_634/Y NOR2X1_LOC_814/A 0.06fF
C19959 INVX1_LOC_53/A NOR2X1_LOC_691/B 0.00fF
C19960 NOR2X1_LOC_609/Y NOR2X1_LOC_334/Y 0.01fF
C19961 NOR2X1_LOC_360/Y INVX1_LOC_95/Y 0.02fF
C19962 NOR2X1_LOC_78/B NOR2X1_LOC_329/B 0.14fF
C19963 NOR2X1_LOC_38/B INVX1_LOC_4/Y 0.03fF
C19964 INVX1_LOC_196/A NOR2X1_LOC_567/B 0.10fF
C19965 NOR2X1_LOC_52/B INVX1_LOC_144/A 0.09fF
C19966 NAND2X1_LOC_648/A INVX1_LOC_22/A 0.03fF
C19967 INVX1_LOC_90/A NAND2X1_LOC_170/A 0.02fF
C19968 NOR2X1_LOC_464/Y INVX1_LOC_15/A 0.02fF
C19969 NAND2X1_LOC_351/A INVX1_LOC_176/A 0.00fF
C19970 INPUT_1 INVX1_LOC_22/A 0.04fF
C19971 NAND2X1_LOC_154/Y VDD -0.00fF
C19972 INVX1_LOC_58/A NOR2X1_LOC_583/Y 0.04fF
C19973 NOR2X1_LOC_89/A NOR2X1_LOC_125/Y 0.15fF
C19974 INVX1_LOC_311/A NAND2X1_LOC_629/Y 0.02fF
C19975 NOR2X1_LOC_544/a_36_216# NOR2X1_LOC_78/A 0.00fF
C19976 INVX1_LOC_243/A NAND2X1_LOC_51/B 0.01fF
C19977 INVX1_LOC_41/A NOR2X1_LOC_557/A 0.02fF
C19978 INVX1_LOC_28/A INVX1_LOC_16/A 1.42fF
C19979 NOR2X1_LOC_287/A NOR2X1_LOC_567/B 0.01fF
C19980 INVX1_LOC_30/A NOR2X1_LOC_363/Y 0.10fF
C19981 NOR2X1_LOC_655/B INPUT_0 0.05fF
C19982 NOR2X1_LOC_299/Y NAND2X1_LOC_303/B 0.08fF
C19983 INVX1_LOC_229/Y NAND2X1_LOC_379/a_36_24# 0.01fF
C19984 NOR2X1_LOC_317/B NOR2X1_LOC_78/A 0.01fF
C19985 NOR2X1_LOC_598/B NOR2X1_LOC_89/A 0.08fF
C19986 NAND2X1_LOC_343/a_36_24# INVX1_LOC_28/A 0.01fF
C19987 NOR2X1_LOC_226/A INVX1_LOC_100/A 0.16fF
C19988 NAND2X1_LOC_656/A INVX1_LOC_46/A 0.17fF
C19989 NOR2X1_LOC_667/A NOR2X1_LOC_167/Y 0.02fF
C19990 NAND2X1_LOC_364/A INVX1_LOC_117/A 0.10fF
C19991 INVX1_LOC_11/A NOR2X1_LOC_155/A 0.04fF
C19992 NOR2X1_LOC_82/A NOR2X1_LOC_101/a_36_216# 0.01fF
C19993 NOR2X1_LOC_814/A NAND2X1_LOC_473/A 0.92fF
C19994 NAND2X1_LOC_858/B NAND2X1_LOC_862/A 0.00fF
C19995 NOR2X1_LOC_465/a_36_216# INVX1_LOC_290/Y 0.00fF
C19996 INVX1_LOC_116/Y NAND2X1_LOC_72/B 0.04fF
C19997 INVX1_LOC_63/Y NOR2X1_LOC_56/Y 0.03fF
C19998 INVX1_LOC_32/A INVX1_LOC_23/A 0.13fF
C19999 NAND2X1_LOC_731/a_36_24# NAND2X1_LOC_863/A 0.06fF
C20000 INVX1_LOC_18/A NAND2X1_LOC_848/A 0.01fF
C20001 NOR2X1_LOC_803/A NOR2X1_LOC_148/B 0.03fF
C20002 INVX1_LOC_64/A INVX1_LOC_290/Y 0.77fF
C20003 NAND2X1_LOC_785/Y NOR2X1_LOC_164/a_36_216# 0.00fF
C20004 NAND2X1_LOC_35/Y NAND2X1_LOC_254/Y 0.04fF
C20005 NOR2X1_LOC_91/A NAND2X1_LOC_175/Y 0.29fF
C20006 NOR2X1_LOC_590/A NAND2X1_LOC_656/B 0.01fF
C20007 NOR2X1_LOC_246/A NAND2X1_LOC_807/Y 0.04fF
C20008 NOR2X1_LOC_55/a_36_216# INVX1_LOC_23/Y 0.01fF
C20009 NOR2X1_LOC_329/Y INVX1_LOC_23/A 0.07fF
C20010 NOR2X1_LOC_413/Y NOR2X1_LOC_24/Y 0.12fF
C20011 NOR2X1_LOC_589/A NAND2X1_LOC_832/Y 0.12fF
C20012 NOR2X1_LOC_690/A NAND2X1_LOC_244/A 0.00fF
C20013 INVX1_LOC_67/A NOR2X1_LOC_137/Y 0.03fF
C20014 INVX1_LOC_83/A D_INPUT_4 0.04fF
C20015 NOR2X1_LOC_512/Y INVX1_LOC_38/A 0.01fF
C20016 NAND2X1_LOC_358/Y INPUT_0 0.03fF
C20017 INVX1_LOC_63/Y NOR2X1_LOC_69/a_36_216# 0.01fF
C20018 NAND2X1_LOC_222/A NAND2X1_LOC_223/B 0.00fF
C20019 INVX1_LOC_63/Y VDD 2.25fF
C20020 NAND2X1_LOC_714/B INVX1_LOC_12/A 0.01fF
C20021 INVX1_LOC_50/A NOR2X1_LOC_278/Y 0.02fF
C20022 NOR2X1_LOC_27/Y INVX1_LOC_20/A 0.05fF
C20023 INVX1_LOC_208/A NOR2X1_LOC_78/A 0.07fF
C20024 NOR2X1_LOC_468/Y NAND2X1_LOC_81/B 0.07fF
C20025 NOR2X1_LOC_500/B NOR2X1_LOC_862/B 0.37fF
C20026 INVX1_LOC_23/A NAND2X1_LOC_175/Y 0.01fF
C20027 INPUT_0 NOR2X1_LOC_99/B 0.09fF
C20028 NOR2X1_LOC_122/Y NAND2X1_LOC_123/Y 0.00fF
C20029 NOR2X1_LOC_516/B NOR2X1_LOC_78/A 4.22fF
C20030 INVX1_LOC_57/A INVX1_LOC_23/Y 0.11fF
C20031 NAND2X1_LOC_632/B INVX1_LOC_38/A 0.14fF
C20032 INVX1_LOC_32/Y INVX1_LOC_91/A 0.01fF
C20033 NOR2X1_LOC_71/Y NAND2X1_LOC_270/a_36_24# 0.01fF
C20034 INVX1_LOC_225/A INVX1_LOC_12/Y 0.10fF
C20035 NAND2X1_LOC_561/B INVX1_LOC_12/A 0.78fF
C20036 NAND2X1_LOC_357/B NAND2X1_LOC_721/A 0.08fF
C20037 NOR2X1_LOC_272/Y INVX1_LOC_3/Y 0.10fF
C20038 NOR2X1_LOC_576/B NOR2X1_LOC_387/A 0.02fF
C20039 NAND2X1_LOC_802/A INVX1_LOC_54/A 0.01fF
C20040 NOR2X1_LOC_667/A INVX1_LOC_76/A 0.04fF
C20041 NOR2X1_LOC_301/A NAND2X1_LOC_793/B 0.10fF
C20042 NOR2X1_LOC_577/Y INVX1_LOC_118/A 0.10fF
C20043 INVX1_LOC_31/A NAND2X1_LOC_489/Y 0.03fF
C20044 INVX1_LOC_8/A NOR2X1_LOC_536/A 0.13fF
C20045 NOR2X1_LOC_717/B INVX1_LOC_78/Y 0.00fF
C20046 INVX1_LOC_248/A INVX1_LOC_76/A 0.10fF
C20047 NOR2X1_LOC_92/Y INVX1_LOC_170/Y 0.05fF
C20048 NOR2X1_LOC_590/A NOR2X1_LOC_721/B 0.12fF
C20049 VDD NAND2X1_LOC_839/A 0.00fF
C20050 INVX1_LOC_256/A INVX1_LOC_29/A 0.06fF
C20051 NAND2X1_LOC_357/B NOR2X1_LOC_323/a_36_216# 0.00fF
C20052 NOR2X1_LOC_420/Y INVX1_LOC_4/Y 0.27fF
C20053 NAND2X1_LOC_9/Y NAND2X1_LOC_99/A 0.03fF
C20054 NAND2X1_LOC_716/a_36_24# NAND2X1_LOC_212/Y 0.01fF
C20055 NOR2X1_LOC_773/Y NOR2X1_LOC_280/Y 0.04fF
C20056 NAND2X1_LOC_551/A INVX1_LOC_6/A 0.01fF
C20057 NOR2X1_LOC_602/A INVX1_LOC_63/A 0.03fF
C20058 INVX1_LOC_16/A NOR2X1_LOC_253/Y 0.01fF
C20059 NOR2X1_LOC_523/A NOR2X1_LOC_861/Y 0.06fF
C20060 NOR2X1_LOC_591/a_36_216# INVX1_LOC_38/A 0.00fF
C20061 INVX1_LOC_55/Y INVX1_LOC_6/A 0.03fF
C20062 INVX1_LOC_182/A INPUT_0 0.12fF
C20063 INVX1_LOC_303/A NOR2X1_LOC_862/B 0.10fF
C20064 NOR2X1_LOC_550/B INVX1_LOC_307/A 0.10fF
C20065 NOR2X1_LOC_572/a_36_216# INVX1_LOC_74/A 0.01fF
C20066 NOR2X1_LOC_433/A NOR2X1_LOC_155/A 0.16fF
C20067 INVX1_LOC_22/A NOR2X1_LOC_586/Y 0.01fF
C20068 NOR2X1_LOC_457/B INVX1_LOC_84/A 0.07fF
C20069 INVX1_LOC_290/A NOR2X1_LOC_585/Y 0.05fF
C20070 NOR2X1_LOC_269/a_36_216# INVX1_LOC_46/A 0.02fF
C20071 NAND2X1_LOC_112/Y NAND2X1_LOC_211/Y 0.02fF
C20072 NAND2X1_LOC_553/A NAND2X1_LOC_99/A 0.00fF
C20073 NOR2X1_LOC_593/Y NOR2X1_LOC_155/A 0.03fF
C20074 INVX1_LOC_228/A NOR2X1_LOC_649/B 0.31fF
C20075 NOR2X1_LOC_773/Y NAND2X1_LOC_811/B 0.03fF
C20076 NOR2X1_LOC_87/Y INVX1_LOC_280/A 0.05fF
C20077 INVX1_LOC_8/A NAND2X1_LOC_93/B 0.00fF
C20078 INVX1_LOC_228/A INVX1_LOC_3/A 0.01fF
C20079 NAND2X1_LOC_577/A NOR2X1_LOC_671/Y 0.03fF
C20080 INPUT_3 NOR2X1_LOC_847/a_36_216# 0.00fF
C20081 NAND2X1_LOC_796/Y INVX1_LOC_20/A 0.01fF
C20082 NAND2X1_LOC_833/Y NOR2X1_LOC_88/Y 0.01fF
C20083 INVX1_LOC_266/Y INVX1_LOC_54/A 0.01fF
C20084 NOR2X1_LOC_826/Y NOR2X1_LOC_392/Y 0.00fF
C20085 INVX1_LOC_35/A INVX1_LOC_53/A 0.97fF
C20086 INVX1_LOC_1/A NAND2X1_LOC_72/B 0.01fF
C20087 NOR2X1_LOC_617/a_36_216# NAND2X1_LOC_489/Y 0.00fF
C20088 NOR2X1_LOC_151/Y INVX1_LOC_78/Y 0.07fF
C20089 INVX1_LOC_290/A INVX1_LOC_77/Y 0.04fF
C20090 NOR2X1_LOC_329/B NOR2X1_LOC_311/Y 0.03fF
C20091 INVX1_LOC_298/Y NOR2X1_LOC_348/Y 0.07fF
C20092 INVX1_LOC_257/Y INVX1_LOC_92/A -0.07fF
C20093 NOR2X1_LOC_52/B NOR2X1_LOC_155/A 0.14fF
C20094 INVX1_LOC_161/Y INVX1_LOC_21/Y 0.54fF
C20095 INVX1_LOC_33/A NOR2X1_LOC_127/Y 0.72fF
C20096 NAND2X1_LOC_170/A INVX1_LOC_38/A 0.03fF
C20097 INVX1_LOC_75/A NOR2X1_LOC_343/a_36_216# 0.00fF
C20098 NOR2X1_LOC_516/a_36_216# NOR2X1_LOC_649/B 0.01fF
C20099 INVX1_LOC_31/A INVX1_LOC_32/A 0.15fF
C20100 NAND2X1_LOC_36/A NAND2X1_LOC_430/B 0.02fF
C20101 NAND2X1_LOC_833/Y INVX1_LOC_84/A 0.30fF
C20102 NOR2X1_LOC_561/Y NOR2X1_LOC_506/a_36_216# 0.01fF
C20103 INVX1_LOC_35/A NAND2X1_LOC_394/a_36_24# 0.01fF
C20104 INVX1_LOC_58/A NOR2X1_LOC_272/Y 0.05fF
C20105 INVX1_LOC_49/A INVX1_LOC_186/Y 0.14fF
C20106 INVX1_LOC_201/Y NAND2X1_LOC_657/a_36_24# 0.03fF
C20107 NOR2X1_LOC_273/Y INVX1_LOC_12/A 0.05fF
C20108 INVX1_LOC_8/A INVX1_LOC_3/A 0.15fF
C20109 NOR2X1_LOC_846/Y INVX1_LOC_108/Y 0.01fF
C20110 INVX1_LOC_22/A INVX1_LOC_118/A 0.24fF
C20111 NOR2X1_LOC_759/Y INVX1_LOC_12/A 0.12fF
C20112 INVX1_LOC_244/Y NOR2X1_LOC_584/Y 0.02fF
C20113 NOR2X1_LOC_589/A INVX1_LOC_9/A 0.03fF
C20114 INVX1_LOC_298/Y INVX1_LOC_256/A 0.07fF
C20115 NOR2X1_LOC_92/Y INVX1_LOC_271/A 0.13fF
C20116 INVX1_LOC_49/A NOR2X1_LOC_777/B 0.03fF
C20117 NOR2X1_LOC_332/A NOR2X1_LOC_115/a_36_216# 0.01fF
C20118 INVX1_LOC_41/Y INVX1_LOC_102/A 0.04fF
C20119 INVX1_LOC_279/Y NOR2X1_LOC_334/Y 0.03fF
C20120 INVX1_LOC_75/A NAND2X1_LOC_212/Y 0.02fF
C20121 INVX1_LOC_24/A INVX1_LOC_42/A 2.44fF
C20122 INVX1_LOC_35/A NOR2X1_LOC_242/A 0.03fF
C20123 NOR2X1_LOC_570/B INVX1_LOC_19/A 0.00fF
C20124 NAND2X1_LOC_563/Y INVX1_LOC_203/A 0.10fF
C20125 INVX1_LOC_246/Y NOR2X1_LOC_48/B 0.01fF
C20126 NOR2X1_LOC_329/B INVX1_LOC_46/A 4.50fF
C20127 INVX1_LOC_5/A INVX1_LOC_38/Y 0.35fF
C20128 INVX1_LOC_31/A NAND2X1_LOC_175/Y 0.19fF
C20129 NOR2X1_LOC_230/a_36_216# NOR2X1_LOC_158/Y 0.01fF
C20130 NOR2X1_LOC_457/B INVX1_LOC_15/A 0.49fF
C20131 NAND2X1_LOC_51/B INVX1_LOC_76/A 0.02fF
C20132 NOR2X1_LOC_303/Y NOR2X1_LOC_169/a_36_216# 0.13fF
C20133 NOR2X1_LOC_290/Y NAND2X1_LOC_489/Y 0.03fF
C20134 NOR2X1_LOC_32/B NOR2X1_LOC_15/Y 0.07fF
C20135 NAND2X1_LOC_802/A NOR2X1_LOC_48/B 0.12fF
C20136 INVX1_LOC_75/A D_INPUT_3 0.17fF
C20137 INVX1_LOC_36/A NOR2X1_LOC_158/Y 0.08fF
C20138 INVX1_LOC_302/Y VDD 0.55fF
C20139 INVX1_LOC_72/A INVX1_LOC_94/Y 0.06fF
C20140 NAND2X1_LOC_222/B NOR2X1_LOC_598/B 0.01fF
C20141 NOR2X1_LOC_197/A INVX1_LOC_50/A 0.03fF
C20142 INVX1_LOC_75/A INVX1_LOC_14/Y 0.25fF
C20143 NOR2X1_LOC_590/A NAND2X1_LOC_286/B 0.00fF
C20144 NOR2X1_LOC_400/B NAND2X1_LOC_555/Y 0.01fF
C20145 INVX1_LOC_2/A INVX1_LOC_186/Y 0.08fF
C20146 NOR2X1_LOC_626/a_36_216# NOR2X1_LOC_626/Y 0.00fF
C20147 INVX1_LOC_45/A NOR2X1_LOC_301/A 0.01fF
C20148 NOR2X1_LOC_557/Y INVX1_LOC_42/A 0.19fF
C20149 NOR2X1_LOC_103/Y NAND2X1_LOC_203/a_36_24# 0.00fF
C20150 INVX1_LOC_7/Y INVX1_LOC_27/A 0.01fF
C20151 INVX1_LOC_36/A NOR2X1_LOC_25/Y 0.01fF
C20152 INVX1_LOC_17/A NAND2X1_LOC_793/B 0.07fF
C20153 D_INPUT_1 NAND2X1_LOC_381/a_36_24# 0.00fF
C20154 NAND2X1_LOC_53/Y INVX1_LOC_259/Y 0.01fF
C20155 NOR2X1_LOC_598/B INVX1_LOC_11/A 0.38fF
C20156 NAND2X1_LOC_308/Y NOR2X1_LOC_89/A 0.00fF
C20157 INVX1_LOC_224/A INVX1_LOC_51/A 0.02fF
C20158 NOR2X1_LOC_357/Y INVX1_LOC_6/A 0.84fF
C20159 INVX1_LOC_10/A NOR2X1_LOC_13/a_36_216# 0.00fF
C20160 NOR2X1_LOC_345/A NOR2X1_LOC_342/A 0.12fF
C20161 D_INPUT_1 NAND2X1_LOC_382/a_36_24# 0.00fF
C20162 INVX1_LOC_11/A INVX1_LOC_51/A 0.00fF
C20163 INVX1_LOC_77/A INVX1_LOC_4/A 0.80fF
C20164 NAND2X1_LOC_465/Y NAND2X1_LOC_254/Y 0.02fF
C20165 NOR2X1_LOC_443/Y NOR2X1_LOC_688/Y 0.06fF
C20166 NOR2X1_LOC_234/Y NAND2X1_LOC_254/Y 0.01fF
C20167 INPUT_0 NOR2X1_LOC_176/Y 0.01fF
C20168 INVX1_LOC_24/A INVX1_LOC_78/A 1.69fF
C20169 INVX1_LOC_226/Y INVX1_LOC_293/Y 0.02fF
C20170 NOR2X1_LOC_163/Y INVX1_LOC_38/A 0.07fF
C20171 INVX1_LOC_21/A INVX1_LOC_163/A 0.08fF
C20172 NAND2X1_LOC_555/Y NAND2X1_LOC_38/a_36_24# 0.00fF
C20173 INVX1_LOC_91/A INVX1_LOC_115/A 0.00fF
C20174 INVX1_LOC_90/A INVX1_LOC_179/A 0.03fF
C20175 NAND2X1_LOC_859/Y NAND2X1_LOC_489/Y 0.03fF
C20176 INVX1_LOC_30/A INVX1_LOC_29/Y 0.09fF
C20177 NOR2X1_LOC_78/A NAND2X1_LOC_211/Y 0.03fF
C20178 NOR2X1_LOC_719/B INVX1_LOC_84/A 0.17fF
C20179 INVX1_LOC_71/A NOR2X1_LOC_301/A 0.17fF
C20180 NOR2X1_LOC_92/Y INVX1_LOC_237/A 0.13fF
C20181 INVX1_LOC_143/A INVX1_LOC_42/A 0.07fF
C20182 INVX1_LOC_245/Y INVX1_LOC_298/A 0.00fF
C20183 NAND2X1_LOC_552/A NOR2X1_LOC_369/Y 0.02fF
C20184 NOR2X1_LOC_151/Y NOR2X1_LOC_680/a_36_216# 0.00fF
C20185 INVX1_LOC_226/Y NAND2X1_LOC_74/B 0.27fF
C20186 NOR2X1_LOC_717/a_36_216# INVX1_LOC_271/Y 0.00fF
C20187 INVX1_LOC_22/A NAND2X1_LOC_63/Y 0.02fF
C20188 INVX1_LOC_135/A NOR2X1_LOC_673/A 0.03fF
C20189 NAND2X1_LOC_348/A NOR2X1_LOC_332/Y 0.03fF
C20190 NOR2X1_LOC_65/B INVX1_LOC_24/A 0.03fF
C20191 INVX1_LOC_71/A NOR2X1_LOC_302/A 0.02fF
C20192 INVX1_LOC_58/A NAND2X1_LOC_364/A 0.08fF
C20193 NOR2X1_LOC_355/A NAND2X1_LOC_475/Y 0.10fF
C20194 INVX1_LOC_269/A INVX1_LOC_239/A 0.01fF
C20195 NOR2X1_LOC_68/A NOR2X1_LOC_414/Y 0.04fF
C20196 NOR2X1_LOC_139/Y NOR2X1_LOC_139/a_36_216# 0.02fF
C20197 INVX1_LOC_41/Y NAND2X1_LOC_439/a_36_24# 0.00fF
C20198 INPUT_4 INVX1_LOC_46/A 0.01fF
C20199 NOR2X1_LOC_82/A NOR2X1_LOC_789/B 0.01fF
C20200 NOR2X1_LOC_186/Y NOR2X1_LOC_160/B 0.03fF
C20201 NAND2X1_LOC_11/Y NAND2X1_LOC_95/a_36_24# 0.00fF
C20202 VDD NOR2X1_LOC_823/Y 0.24fF
C20203 INVX1_LOC_100/A INVX1_LOC_118/A 0.07fF
C20204 NAND2X1_LOC_552/A INVX1_LOC_286/Y 0.02fF
C20205 INVX1_LOC_49/A NOR2X1_LOC_843/B 0.03fF
C20206 INVX1_LOC_12/Y NAND2X1_LOC_642/Y 0.01fF
C20207 NAND2X1_LOC_565/B INVX1_LOC_42/A 0.03fF
C20208 INVX1_LOC_191/A INVX1_LOC_54/A 0.21fF
C20209 NAND2X1_LOC_190/Y NOR2X1_LOC_205/Y 0.00fF
C20210 INVX1_LOC_10/A NAND2X1_LOC_74/B 0.21fF
C20211 INVX1_LOC_157/A INVX1_LOC_29/A 0.03fF
C20212 NOR2X1_LOC_609/A NOR2X1_LOC_717/A 0.21fF
C20213 NOR2X1_LOC_480/a_36_216# D_GATE_479 0.02fF
C20214 NOR2X1_LOC_415/A INVX1_LOC_29/A 0.01fF
C20215 NOR2X1_LOC_65/B NOR2X1_LOC_557/Y 0.28fF
C20216 NAND2X1_LOC_9/Y NAND2X1_LOC_656/A 0.55fF
C20217 INVX1_LOC_33/A NOR2X1_LOC_383/B 7.09fF
C20218 NOR2X1_LOC_433/A NOR2X1_LOC_125/Y 0.07fF
C20219 INVX1_LOC_14/Y NOR2X1_LOC_309/a_36_216# 0.00fF
C20220 INVX1_LOC_178/A INVX1_LOC_286/Y 0.10fF
C20221 NAND2X1_LOC_803/B NAND2X1_LOC_537/Y 0.48fF
C20222 NOR2X1_LOC_564/Y INVX1_LOC_63/A 0.03fF
C20223 INVX1_LOC_143/A INVX1_LOC_78/A 0.07fF
C20224 NOR2X1_LOC_220/A INVX1_LOC_4/Y 0.16fF
C20225 NOR2X1_LOC_315/Y NOR2X1_LOC_134/a_36_216# 0.00fF
C20226 NOR2X1_LOC_174/B NOR2X1_LOC_633/A 0.26fF
C20227 NAND2X1_LOC_303/Y NOR2X1_LOC_599/Y 0.03fF
C20228 INVX1_LOC_5/A INVX1_LOC_159/A 0.10fF
C20229 NOR2X1_LOC_86/A INVX1_LOC_3/Y 0.10fF
C20230 NAND2X1_LOC_800/Y INVX1_LOC_42/A 0.10fF
C20231 NOR2X1_LOC_590/A NAND2X1_LOC_537/Y 0.07fF
C20232 NOR2X1_LOC_454/Y NOR2X1_LOC_585/a_36_216# 0.01fF
C20233 NOR2X1_LOC_857/A INVX1_LOC_117/A 0.08fF
C20234 NOR2X1_LOC_130/A INVX1_LOC_42/A 0.07fF
C20235 NAND2X1_LOC_739/B NOR2X1_LOC_304/Y 0.02fF
C20236 NOR2X1_LOC_815/A NOR2X1_LOC_697/Y 0.01fF
C20237 INVX1_LOC_136/A NAND2X1_LOC_474/Y 0.13fF
C20238 INVX1_LOC_64/A INVX1_LOC_77/A 0.27fF
C20239 NOR2X1_LOC_598/B NOR2X1_LOC_593/Y 0.02fF
C20240 NAND2X1_LOC_116/A INVX1_LOC_57/A 0.02fF
C20241 NAND2X1_LOC_633/a_36_24# INVX1_LOC_181/A 0.00fF
C20242 INVX1_LOC_278/A NAND2X1_LOC_833/Y 0.03fF
C20243 NOR2X1_LOC_798/A NAND2X1_LOC_656/A 0.03fF
C20244 NAND2X1_LOC_477/A INVX1_LOC_271/A 0.03fF
C20245 NOR2X1_LOC_804/a_36_216# NOR2X1_LOC_383/B 0.00fF
C20246 NOR2X1_LOC_548/Y INVX1_LOC_4/Y 0.25fF
C20247 INVX1_LOC_20/A INVX1_LOC_9/A 0.03fF
C20248 NAND2X1_LOC_715/B NOR2X1_LOC_433/A 0.37fF
C20249 NOR2X1_LOC_65/B INVX1_LOC_143/A 0.39fF
C20250 NOR2X1_LOC_296/Y INVX1_LOC_31/A 0.28fF
C20251 NOR2X1_LOC_15/Y INVX1_LOC_195/Y 0.01fF
C20252 NOR2X1_LOC_45/B INVX1_LOC_107/Y 0.04fF
C20253 NOR2X1_LOC_207/A INVX1_LOC_105/Y 0.02fF
C20254 INVX1_LOC_17/A INVX1_LOC_45/A 2.86fF
C20255 INVX1_LOC_6/A NAND2X1_LOC_489/Y 0.01fF
C20256 NAND2X1_LOC_773/Y NOR2X1_LOC_360/Y 0.10fF
C20257 INVX1_LOC_313/A INVX1_LOC_32/A 0.03fF
C20258 NOR2X1_LOC_76/A INVX1_LOC_15/A 0.03fF
C20259 NOR2X1_LOC_601/Y NOR2X1_LOC_155/A 0.01fF
C20260 INPUT_3 INVX1_LOC_31/A 0.21fF
C20261 INVX1_LOC_35/A INVX1_LOC_80/Y 0.09fF
C20262 INVX1_LOC_286/Y NOR2X1_LOC_816/A 1.09fF
C20263 NAND2X1_LOC_361/Y INVX1_LOC_50/Y 0.10fF
C20264 INVX1_LOC_12/Y NOR2X1_LOC_271/Y 0.03fF
C20265 INVX1_LOC_40/A NOR2X1_LOC_383/B 0.03fF
C20266 NOR2X1_LOC_180/B INVX1_LOC_15/A 0.03fF
C20267 NOR2X1_LOC_160/B NAND2X1_LOC_198/a_36_24# 0.00fF
C20268 NOR2X1_LOC_27/Y INVX1_LOC_64/A 0.01fF
C20269 NOR2X1_LOC_32/B INVX1_LOC_15/Y 0.14fF
C20270 NAND2X1_LOC_783/A INVX1_LOC_78/A 0.00fF
C20271 INVX1_LOC_211/Y INVX1_LOC_36/A 0.01fF
C20272 NAND2X1_LOC_762/a_36_24# NAND2X1_LOC_30/Y 0.00fF
C20273 NAND2X1_LOC_30/Y INVX1_LOC_18/A 0.18fF
C20274 INVX1_LOC_286/A INVX1_LOC_19/A 0.08fF
C20275 NOR2X1_LOC_130/A INVX1_LOC_78/A 0.03fF
C20276 NOR2X1_LOC_73/a_36_216# INVX1_LOC_47/Y 0.01fF
C20277 INVX1_LOC_41/A INVX1_LOC_27/A 0.27fF
C20278 NOR2X1_LOC_205/Y NOR2X1_LOC_596/A 0.03fF
C20279 INVX1_LOC_232/A INVX1_LOC_57/A 1.26fF
C20280 INVX1_LOC_69/Y INVX1_LOC_29/A 0.11fF
C20281 NAND2X1_LOC_12/a_36_24# NAND2X1_LOC_30/Y 0.00fF
C20282 NOR2X1_LOC_536/A INVX1_LOC_118/Y 0.00fF
C20283 INVX1_LOC_278/A INVX1_LOC_164/Y 0.02fF
C20284 NOR2X1_LOC_45/Y NAND2X1_LOC_195/Y 0.26fF
C20285 NOR2X1_LOC_788/a_36_216# INVX1_LOC_29/A 0.01fF
C20286 INVX1_LOC_35/A NOR2X1_LOC_78/B 0.17fF
C20287 INVX1_LOC_201/Y INVX1_LOC_27/A 0.64fF
C20288 NOR2X1_LOC_653/B INVX1_LOC_225/A 0.01fF
C20289 NOR2X1_LOC_498/Y NOR2X1_LOC_824/A 0.01fF
C20290 INVX1_LOC_25/A INVX1_LOC_53/Y 0.00fF
C20291 INPUT_0 NOR2X1_LOC_850/B 0.06fF
C20292 INVX1_LOC_17/A INVX1_LOC_71/A 0.54fF
C20293 INVX1_LOC_100/Y NAND2X1_LOC_81/B 0.07fF
C20294 NOR2X1_LOC_67/A NAND2X1_LOC_569/B 0.10fF
C20295 INVX1_LOC_73/A INVX1_LOC_15/A 0.02fF
C20296 NAND2X1_LOC_860/A NOR2X1_LOC_82/Y 0.02fF
C20297 NAND2X1_LOC_500/B INVX1_LOC_91/A 0.01fF
C20298 NOR2X1_LOC_647/A D_INPUT_0 0.01fF
C20299 NAND2X1_LOC_561/B NAND2X1_LOC_787/B 0.02fF
C20300 INVX1_LOC_24/A NOR2X1_LOC_503/Y 0.23fF
C20301 NOR2X1_LOC_753/Y NAND2X1_LOC_538/Y 0.04fF
C20302 INVX1_LOC_58/A NOR2X1_LOC_86/A 0.13fF
C20303 NOR2X1_LOC_626/Y NAND2X1_LOC_629/Y 0.05fF
C20304 NOR2X1_LOC_15/Y INVX1_LOC_155/Y 0.70fF
C20305 NOR2X1_LOC_45/B INVX1_LOC_272/A 1.05fF
C20306 INVX1_LOC_34/A NAND2X1_LOC_579/A 0.07fF
C20307 NOR2X1_LOC_65/B NOR2X1_LOC_130/A 0.03fF
C20308 NOR2X1_LOC_135/Y NOR2X1_LOC_334/Y 0.19fF
C20309 INVX1_LOC_47/A INVX1_LOC_26/A 0.13fF
C20310 NOR2X1_LOC_543/a_36_216# INVX1_LOC_29/A 0.00fF
C20311 NOR2X1_LOC_74/A INVX1_LOC_47/Y 0.33fF
C20312 NOR2X1_LOC_339/a_36_216# INVX1_LOC_280/A 0.00fF
C20313 NAND2X1_LOC_537/Y NAND2X1_LOC_354/B 0.06fF
C20314 NAND2X1_LOC_538/Y NAND2X1_LOC_325/Y 0.09fF
C20315 NOR2X1_LOC_114/A NOR2X1_LOC_114/Y 0.01fF
C20316 NOR2X1_LOC_188/Y INVX1_LOC_53/A 0.00fF
C20317 INVX1_LOC_50/A NOR2X1_LOC_525/Y 0.05fF
C20318 INVX1_LOC_90/A NOR2X1_LOC_693/Y 0.07fF
C20319 INVX1_LOC_269/A NAND2X1_LOC_736/B 0.24fF
C20320 NAND2X1_LOC_802/A NAND2X1_LOC_350/A 0.04fF
C20321 VDD INVX1_LOC_27/Y 0.21fF
C20322 INVX1_LOC_90/A NAND2X1_LOC_288/B 0.22fF
C20323 INVX1_LOC_50/A NOR2X1_LOC_312/Y 0.74fF
C20324 NOR2X1_LOC_203/a_36_216# NOR2X1_LOC_500/Y 0.01fF
C20325 INVX1_LOC_38/A INVX1_LOC_179/A 0.03fF
C20326 INVX1_LOC_6/A INVX1_LOC_32/A 0.03fF
C20327 NOR2X1_LOC_9/Y INVX1_LOC_47/Y 0.38fF
C20328 INVX1_LOC_132/A NOR2X1_LOC_160/B 0.07fF
C20329 INVX1_LOC_91/A NOR2X1_LOC_114/Y 0.00fF
C20330 NOR2X1_LOC_389/B NAND2X1_LOC_288/B 0.01fF
C20331 NOR2X1_LOC_160/B NOR2X1_LOC_374/A 0.34fF
C20332 NOR2X1_LOC_799/B NAND2X1_LOC_74/B 0.16fF
C20333 INVX1_LOC_35/A NAND2X1_LOC_392/Y 0.06fF
C20334 INVX1_LOC_102/Y NOR2X1_LOC_301/A 0.03fF
C20335 INVX1_LOC_269/A NAND2X1_LOC_320/a_36_24# 0.00fF
C20336 NOR2X1_LOC_82/A NOR2X1_LOC_514/Y 0.01fF
C20337 INVX1_LOC_6/A NOR2X1_LOC_329/Y 0.20fF
C20338 NOR2X1_LOC_723/Y NOR2X1_LOC_596/A 0.02fF
C20339 INVX1_LOC_66/Y NOR2X1_LOC_117/Y 0.01fF
C20340 INVX1_LOC_267/A INVX1_LOC_14/A 0.10fF
C20341 NAND2X1_LOC_373/a_36_24# NOR2X1_LOC_78/B 0.00fF
C20342 NAND2X1_LOC_794/B INVX1_LOC_16/A 0.07fF
C20343 INVX1_LOC_35/A INVX1_LOC_83/A 0.22fF
C20344 NAND2X1_LOC_605/a_36_24# INVX1_LOC_186/Y 0.00fF
C20345 NOR2X1_LOC_122/Y INVX1_LOC_271/A 0.01fF
C20346 NOR2X1_LOC_548/B NAND2X1_LOC_72/B 0.03fF
C20347 INVX1_LOC_225/A NOR2X1_LOC_160/B 0.07fF
C20348 NOR2X1_LOC_65/B NOR2X1_LOC_216/Y 0.01fF
C20349 NOR2X1_LOC_775/Y INVX1_LOC_57/A 0.04fF
C20350 INVX1_LOC_278/A NOR2X1_LOC_76/A 0.73fF
C20351 NOR2X1_LOC_590/A NOR2X1_LOC_486/B 0.00fF
C20352 NOR2X1_LOC_288/A NOR2X1_LOC_160/B 0.03fF
C20353 INVX1_LOC_280/A NOR2X1_LOC_673/A 0.07fF
C20354 INVX1_LOC_11/A NAND2X1_LOC_660/A 0.07fF
C20355 NOR2X1_LOC_155/A NOR2X1_LOC_676/a_36_216# 0.00fF
C20356 INVX1_LOC_299/A NAND2X1_LOC_323/B 0.03fF
C20357 INVX1_LOC_2/A NAND2X1_LOC_799/A 0.51fF
C20358 NOR2X1_LOC_246/A NOR2X1_LOC_109/Y 0.01fF
C20359 INVX1_LOC_140/A NAND2X1_LOC_408/a_36_24# 0.00fF
C20360 INVX1_LOC_48/Y INVX1_LOC_16/A 0.12fF
C20361 NOR2X1_LOC_606/Y INVX1_LOC_8/A 0.02fF
C20362 INVX1_LOC_298/Y INVX1_LOC_69/Y 0.02fF
C20363 NAND2X1_LOC_149/Y INVX1_LOC_290/A 0.09fF
C20364 NOR2X1_LOC_533/A NOR2X1_LOC_533/Y 0.01fF
C20365 NOR2X1_LOC_372/A NOR2X1_LOC_52/B 0.03fF
C20366 INVX1_LOC_49/A INVX1_LOC_18/A 0.17fF
C20367 NOR2X1_LOC_332/A INVX1_LOC_38/Y 0.25fF
C20368 INVX1_LOC_1/A INVX1_LOC_53/Y 0.01fF
C20369 NOR2X1_LOC_280/Y INVX1_LOC_42/A 0.17fF
C20370 INVX1_LOC_158/A INVX1_LOC_31/A 0.06fF
C20371 NOR2X1_LOC_321/Y NAND2X1_LOC_660/Y 0.00fF
C20372 INVX1_LOC_77/Y INVX1_LOC_261/Y 0.14fF
C20373 NOR2X1_LOC_360/A NOR2X1_LOC_861/Y 0.02fF
C20374 INVX1_LOC_24/A NOR2X1_LOC_152/Y 0.18fF
C20375 INVX1_LOC_243/A INVX1_LOC_174/A 0.03fF
C20376 NOR2X1_LOC_690/A NOR2X1_LOC_86/Y 0.01fF
C20377 NOR2X1_LOC_67/A NOR2X1_LOC_530/Y 0.01fF
C20378 NOR2X1_LOC_789/B INVX1_LOC_306/A 0.00fF
C20379 NOR2X1_LOC_268/a_36_216# NOR2X1_LOC_172/Y -0.00fF
C20380 INVX1_LOC_24/A INVX1_LOC_113/Y 0.00fF
C20381 NOR2X1_LOC_550/a_36_216# INVX1_LOC_177/A 0.00fF
C20382 NAND2X1_LOC_350/B NOR2X1_LOC_45/Y 0.51fF
C20383 NOR2X1_LOC_92/Y INVX1_LOC_234/A 0.93fF
C20384 NOR2X1_LOC_151/Y NOR2X1_LOC_717/A 0.00fF
C20385 INVX1_LOC_269/A NOR2X1_LOC_543/A 0.02fF
C20386 INVX1_LOC_54/A INVX1_LOC_19/A 0.31fF
C20387 INVX1_LOC_36/A INVX1_LOC_236/A 0.01fF
C20388 INVX1_LOC_54/A NOR2X1_LOC_11/Y 0.88fF
C20389 NAND2X1_LOC_93/B NOR2X1_LOC_258/Y 0.10fF
C20390 NOR2X1_LOC_337/A INVX1_LOC_58/Y 0.08fF
C20391 INVX1_LOC_286/Y NOR2X1_LOC_773/Y 0.10fF
C20392 D_INPUT_7 NOR2X1_LOC_1/a_36_216# 0.00fF
C20393 INVX1_LOC_215/A INVX1_LOC_161/Y 0.02fF
C20394 INVX1_LOC_45/Y NOR2X1_LOC_392/B 0.01fF
C20395 NOR2X1_LOC_609/a_36_216# NOR2X1_LOC_388/Y 0.00fF
C20396 NAND2X1_LOC_794/B INVX1_LOC_28/A 0.21fF
C20397 INVX1_LOC_2/A INVX1_LOC_18/A 0.62fF
C20398 INVX1_LOC_95/Y INVX1_LOC_26/A 0.04fF
C20399 INVX1_LOC_2/A NAND2X1_LOC_728/Y 0.07fF
C20400 NAND2X1_LOC_425/Y NOR2X1_LOC_258/Y 0.03fF
C20401 NAND2X1_LOC_564/B INVX1_LOC_31/A 0.03fF
C20402 NOR2X1_LOC_82/A NOR2X1_LOC_128/B 0.00fF
C20403 INVX1_LOC_14/A INVX1_LOC_89/A 0.16fF
C20404 INVX1_LOC_78/A NOR2X1_LOC_280/Y 0.03fF
C20405 INVX1_LOC_104/A NOR2X1_LOC_303/Y 0.10fF
C20406 NOR2X1_LOC_374/A NOR2X1_LOC_317/B 0.70fF
C20407 NOR2X1_LOC_226/A INVX1_LOC_18/A 0.09fF
C20408 NAND2X1_LOC_703/Y NOR2X1_LOC_329/B 0.00fF
C20409 INVX1_LOC_102/A INVX1_LOC_185/A 0.02fF
C20410 INVX1_LOC_24/A NOR2X1_LOC_721/A 0.02fF
C20411 NOR2X1_LOC_276/Y INVX1_LOC_10/A 0.03fF
C20412 NOR2X1_LOC_92/Y NOR2X1_LOC_19/B 0.07fF
C20413 INVX1_LOC_136/A NOR2X1_LOC_500/Y 0.10fF
C20414 NOR2X1_LOC_222/a_36_216# INVX1_LOC_30/A 0.00fF
C20415 INVX1_LOC_256/A NAND2X1_LOC_140/A 0.01fF
C20416 INVX1_LOC_58/A NOR2X1_LOC_405/A 0.56fF
C20417 INVX1_LOC_136/A INVX1_LOC_226/Y 0.39fF
C20418 INVX1_LOC_68/Y NOR2X1_LOC_554/B 0.01fF
C20419 INVX1_LOC_45/Y NAND2X1_LOC_294/a_36_24# 0.00fF
C20420 NAND2X1_LOC_361/Y NOR2X1_LOC_6/B 0.10fF
C20421 NAND2X1_LOC_50/a_36_24# INPUT_7 0.00fF
C20422 NAND2X1_LOC_74/B NOR2X1_LOC_445/B 0.01fF
C20423 INVX1_LOC_12/A NOR2X1_LOC_13/a_36_216# 0.00fF
C20424 NAND2X1_LOC_799/A NAND2X1_LOC_648/A 0.00fF
C20425 INVX1_LOC_13/A INVX1_LOC_36/A 0.03fF
C20426 NOR2X1_LOC_837/B NOR2X1_LOC_78/B 0.03fF
C20427 NOR2X1_LOC_226/A NOR2X1_LOC_637/Y 0.07fF
C20428 NAND2X1_LOC_49/a_36_24# NOR2X1_LOC_68/A 0.02fF
C20429 INVX1_LOC_9/A INVX1_LOC_4/A 0.07fF
C20430 NAND2X1_LOC_708/Y NOR2X1_LOC_45/B 0.01fF
C20431 INVX1_LOC_88/A NOR2X1_LOC_755/a_36_216# 0.00fF
C20432 NOR2X1_LOC_773/Y NOR2X1_LOC_191/B 0.10fF
C20433 NAND2X1_LOC_33/Y NOR2X1_LOC_413/Y -0.01fF
C20434 NAND2X1_LOC_807/B NAND2X1_LOC_288/A 0.14fF
C20435 NOR2X1_LOC_357/Y INVX1_LOC_270/A 0.12fF
C20436 NOR2X1_LOC_598/B INVX1_LOC_199/A 0.03fF
C20437 NOR2X1_LOC_168/A INVX1_LOC_33/A 0.01fF
C20438 NOR2X1_LOC_91/A NAND2X1_LOC_804/Y 0.12fF
C20439 NAND2X1_LOC_543/Y INVX1_LOC_41/Y 0.00fF
C20440 INVX1_LOC_32/A INVX1_LOC_131/Y 0.15fF
C20441 NAND2X1_LOC_579/A INPUT_0 0.10fF
C20442 NOR2X1_LOC_355/A INVX1_LOC_30/A 0.10fF
C20443 INVX1_LOC_136/A INVX1_LOC_10/A 5.43fF
C20444 NOR2X1_LOC_716/B INVX1_LOC_256/Y 0.57fF
C20445 INVX1_LOC_35/A NOR2X1_LOC_368/Y 0.01fF
C20446 INVX1_LOC_279/A NOR2X1_LOC_360/Y 0.15fF
C20447 INVX1_LOC_72/A INVX1_LOC_66/A 0.01fF
C20448 INVX1_LOC_36/A NOR2X1_LOC_246/A 0.07fF
C20449 INVX1_LOC_278/A NAND2X1_LOC_241/Y 0.04fF
C20450 NOR2X1_LOC_641/B INVX1_LOC_90/A 0.02fF
C20451 NAND2X1_LOC_784/A INVX1_LOC_37/A 0.07fF
C20452 INVX1_LOC_54/Y INVX1_LOC_104/A 0.03fF
C20453 NOR2X1_LOC_828/Y VDD 0.06fF
C20454 NOR2X1_LOC_369/Y INVX1_LOC_140/A 0.02fF
C20455 INVX1_LOC_38/A NOR2X1_LOC_693/Y 0.03fF
C20456 NAND2X1_LOC_725/B INVX1_LOC_309/A 0.03fF
C20457 INVX1_LOC_132/A NOR2X1_LOC_516/B 0.10fF
C20458 NOR2X1_LOC_52/B NAND2X1_LOC_660/A 0.09fF
C20459 INVX1_LOC_83/A NOR2X1_LOC_325/Y 0.00fF
C20460 INVX1_LOC_34/A NAND2X1_LOC_341/a_36_24# 0.00fF
C20461 INVX1_LOC_66/Y INVX1_LOC_270/A 0.03fF
C20462 NOR2X1_LOC_67/Y NOR2X1_LOC_721/B 0.06fF
C20463 INVX1_LOC_36/A INVX1_LOC_55/Y 0.03fF
C20464 INVX1_LOC_234/A NAND2X1_LOC_837/Y 0.01fF
C20465 INVX1_LOC_178/Y NOR2X1_LOC_660/Y 0.00fF
C20466 INVX1_LOC_35/A INVX1_LOC_46/A 0.47fF
C20467 NOR2X1_LOC_401/Y INVX1_LOC_168/A 0.04fF
C20468 NOR2X1_LOC_690/A INVX1_LOC_25/Y 0.00fF
C20469 NAND2X1_LOC_139/A INVX1_LOC_316/Y 0.02fF
C20470 NAND2X1_LOC_807/B INVX1_LOC_19/A 0.03fF
C20471 INVX1_LOC_286/Y INVX1_LOC_140/A 0.10fF
C20472 NOR2X1_LOC_364/A NAND2X1_LOC_454/Y 0.09fF
C20473 INVX1_LOC_18/A INPUT_1 0.03fF
C20474 NAND2X1_LOC_361/Y INVX1_LOC_30/Y 0.03fF
C20475 NOR2X1_LOC_67/A NOR2X1_LOC_709/A 0.03fF
C20476 NOR2X1_LOC_399/A NOR2X1_LOC_399/Y 0.00fF
C20477 INVX1_LOC_12/A NAND2X1_LOC_74/B 0.10fF
C20478 INVX1_LOC_24/A NAND2X1_LOC_861/Y 0.07fF
C20479 NAND2X1_LOC_783/A NOR2X1_LOC_152/Y 0.01fF
C20480 NOR2X1_LOC_671/a_36_216# NOR2X1_LOC_671/Y 0.02fF
C20481 INVX1_LOC_178/A NOR2X1_LOC_56/Y 0.11fF
C20482 NOR2X1_LOC_89/A INVX1_LOC_29/A 0.12fF
C20483 NAND2X1_LOC_552/A VDD 0.04fF
C20484 NOR2X1_LOC_48/B INVX1_LOC_19/A 0.07fF
C20485 INVX1_LOC_178/A NAND2X1_LOC_659/B 0.05fF
C20486 INVX1_LOC_5/A VDD 1.55fF
C20487 NAND2X1_LOC_741/B NOR2X1_LOC_380/Y 0.05fF
C20488 NAND2X1_LOC_347/B INVX1_LOC_93/Y 0.01fF
C20489 NOR2X1_LOC_152/Y NOR2X1_LOC_130/A 0.07fF
C20490 NAND2X1_LOC_84/Y INVX1_LOC_89/A 0.38fF
C20491 NOR2X1_LOC_380/A NAND2X1_LOC_866/A 0.04fF
C20492 NOR2X1_LOC_629/B NAND2X1_LOC_735/B 0.01fF
C20493 NOR2X1_LOC_632/Y NOR2X1_LOC_718/B 0.01fF
C20494 NAND2X1_LOC_725/B INVX1_LOC_11/Y 0.03fF
C20495 NOR2X1_LOC_84/Y INVX1_LOC_16/A 0.10fF
C20496 INVX1_LOC_57/Y NOR2X1_LOC_323/Y 0.16fF
C20497 NOR2X1_LOC_589/A NOR2X1_LOC_367/B 0.07fF
C20498 NAND2X1_LOC_291/B NAND2X1_LOC_233/a_36_24# 0.02fF
C20499 NOR2X1_LOC_231/B NOR2X1_LOC_9/Y 0.05fF
C20500 NOR2X1_LOC_208/Y INVX1_LOC_55/Y 0.07fF
C20501 INVX1_LOC_45/A NOR2X1_LOC_594/Y 0.07fF
C20502 INVX1_LOC_182/Y NOR2X1_LOC_360/Y 0.01fF
C20503 NOR2X1_LOC_482/Y INVX1_LOC_16/A 0.97fF
C20504 NAND2X1_LOC_551/A NOR2X1_LOC_237/Y 0.02fF
C20505 INVX1_LOC_178/A VDD 4.77fF
C20506 INVX1_LOC_49/A NAND2X1_LOC_105/a_36_24# 0.00fF
C20507 NAND2X1_LOC_3/B INVX1_LOC_19/A 0.03fF
C20508 NOR2X1_LOC_19/B NAND2X1_LOC_837/Y 0.01fF
C20509 NOR2X1_LOC_78/B NOR2X1_LOC_121/A 0.03fF
C20510 INVX1_LOC_64/A INVX1_LOC_9/A 0.08fF
C20511 NOR2X1_LOC_739/Y NOR2X1_LOC_833/Y 0.03fF
C20512 NOR2X1_LOC_623/B NOR2X1_LOC_633/A 0.34fF
C20513 NOR2X1_LOC_307/A NOR2X1_LOC_711/Y 0.01fF
C20514 NOR2X1_LOC_246/A NOR2X1_LOC_309/Y 0.02fF
C20515 NAND2X1_LOC_303/Y NAND2X1_LOC_453/A 0.03fF
C20516 NOR2X1_LOC_160/B NAND2X1_LOC_642/Y 0.06fF
C20517 NAND2X1_LOC_326/A INVX1_LOC_37/A 0.08fF
C20518 NOR2X1_LOC_640/Y INVX1_LOC_58/Y 0.00fF
C20519 NOR2X1_LOC_494/Y VDD 0.25fF
C20520 NAND2X1_LOC_680/a_36_24# NOR2X1_LOC_577/Y 0.02fF
C20521 NOR2X1_LOC_644/A NOR2X1_LOC_147/B 0.00fF
C20522 NOR2X1_LOC_654/A NOR2X1_LOC_697/Y 0.02fF
C20523 NOR2X1_LOC_589/A NOR2X1_LOC_131/a_36_216# 0.01fF
C20524 INVX1_LOC_186/Y NOR2X1_LOC_631/Y 0.21fF
C20525 INVX1_LOC_210/Y NOR2X1_LOC_78/A 0.01fF
C20526 INVX1_LOC_271/A NOR2X1_LOC_435/B 0.04fF
C20527 NOR2X1_LOC_576/B NOR2X1_LOC_822/Y 0.02fF
C20528 INVX1_LOC_33/A NOR2X1_LOC_163/Y 0.04fF
C20529 INVX1_LOC_201/Y NOR2X1_LOC_19/B 0.14fF
C20530 NAND2X1_LOC_735/B INVX1_LOC_22/A 0.03fF
C20531 NOR2X1_LOC_561/Y NOR2X1_LOC_131/Y 0.04fF
C20532 INVX1_LOC_84/Y NOR2X1_LOC_459/A 0.02fF
C20533 INVX1_LOC_47/A INVX1_LOC_149/A 0.01fF
C20534 NOR2X1_LOC_263/a_36_216# NAND2X1_LOC_842/B 0.00fF
C20535 INVX1_LOC_174/A INVX1_LOC_76/A 0.12fF
C20536 NOR2X1_LOC_706/Y NOR2X1_LOC_713/B 0.07fF
C20537 NAND2X1_LOC_337/B VDD 1.28fF
C20538 INPUT_5 INVX1_LOC_22/A 0.01fF
C20539 INVX1_LOC_305/Y INVX1_LOC_83/A 0.24fF
C20540 INVX1_LOC_34/Y INPUT_1 0.32fF
C20541 NOR2X1_LOC_816/A VDD 1.11fF
C20542 INVX1_LOC_45/Y NAND2X1_LOC_123/a_36_24# 0.00fF
C20543 INVX1_LOC_206/Y NOR2X1_LOC_303/Y 6.10fF
C20544 NOR2X1_LOC_843/B NAND2X1_LOC_63/Y 0.07fF
C20545 NOR2X1_LOC_142/Y INVX1_LOC_42/Y 0.54fF
C20546 INVX1_LOC_298/Y NOR2X1_LOC_89/A 12.65fF
C20547 NOR2X1_LOC_598/a_36_216# NOR2X1_LOC_78/A 0.00fF
C20548 NOR2X1_LOC_385/Y INVX1_LOC_240/A 0.05fF
C20549 INVX1_LOC_28/A NOR2X1_LOC_84/Y 0.34fF
C20550 INVX1_LOC_141/Y NOR2X1_LOC_305/a_36_216# 0.00fF
C20551 INVX1_LOC_1/A NOR2X1_LOC_652/a_36_216# 0.00fF
C20552 INVX1_LOC_19/A NOR2X1_LOC_836/A 0.00fF
C20553 NOR2X1_LOC_589/A NOR2X1_LOC_561/Y 0.07fF
C20554 NOR2X1_LOC_91/A NOR2X1_LOC_519/a_36_216# 0.00fF
C20555 NAND2X1_LOC_838/Y NAND2X1_LOC_560/A 0.02fF
C20556 INVX1_LOC_251/A INVX1_LOC_4/Y 0.04fF
C20557 INVX1_LOC_30/A INVX1_LOC_126/A 0.12fF
C20558 INVX1_LOC_285/Y INVX1_LOC_63/Y 0.09fF
C20559 INVX1_LOC_17/A NOR2X1_LOC_331/B 0.03fF
C20560 NOR2X1_LOC_191/A NOR2X1_LOC_153/a_36_216# 0.00fF
C20561 INVX1_LOC_255/Y INVX1_LOC_90/A 0.07fF
C20562 INVX1_LOC_30/A NOR2X1_LOC_111/A 0.10fF
C20563 NOR2X1_LOC_471/Y NOR2X1_LOC_331/B 0.00fF
C20564 INVX1_LOC_14/Y NOR2X1_LOC_274/B 0.00fF
C20565 INVX1_LOC_155/A NOR2X1_LOC_78/A 0.03fF
C20566 INVX1_LOC_18/A NOR2X1_LOC_586/Y 0.15fF
C20567 NOR2X1_LOC_160/B NOR2X1_LOC_271/Y 0.55fF
C20568 NAND2X1_LOC_773/Y NOR2X1_LOC_79/Y 0.05fF
C20569 INVX1_LOC_58/A INVX1_LOC_109/Y 0.12fF
C20570 INVX1_LOC_27/A NAND2X1_LOC_574/A 0.05fF
C20571 NOR2X1_LOC_726/Y INVX1_LOC_117/A 0.05fF
C20572 INVX1_LOC_161/Y INVX1_LOC_54/A 0.14fF
C20573 NOR2X1_LOC_137/A INVX1_LOC_150/A 0.50fF
C20574 NOR2X1_LOC_147/a_36_216# INVX1_LOC_23/A 0.00fF
C20575 NOR2X1_LOC_264/Y NOR2X1_LOC_78/A 0.52fF
C20576 INVX1_LOC_35/A NOR2X1_LOC_671/Y 0.03fF
C20577 INVX1_LOC_12/A NOR2X1_LOC_660/Y 0.12fF
C20578 NAND2X1_LOC_331/a_36_24# NOR2X1_LOC_106/A 0.00fF
C20579 NOR2X1_LOC_798/A NOR2X1_LOC_691/B 0.03fF
C20580 INPUT_0 INVX1_LOC_43/A 0.01fF
C20581 GATE_865 NOR2X1_LOC_380/Y 0.05fF
C20582 NOR2X1_LOC_208/Y NOR2X1_LOC_357/Y 1.13fF
C20583 INVX1_LOC_17/A NOR2X1_LOC_592/B 0.00fF
C20584 NAND2X1_LOC_218/B D_INPUT_3 0.67fF
C20585 INVX1_LOC_90/A NOR2X1_LOC_71/Y 0.03fF
C20586 INVX1_LOC_255/Y NAND2X1_LOC_348/A 2.34fF
C20587 INVX1_LOC_11/A NOR2X1_LOC_58/Y 0.07fF
C20588 NOR2X1_LOC_751/Y INVX1_LOC_38/A 0.05fF
C20589 INVX1_LOC_32/A NOR2X1_LOC_416/A 0.10fF
C20590 NOR2X1_LOC_92/Y NAND2X1_LOC_477/Y 0.01fF
C20591 INVX1_LOC_155/Y NOR2X1_LOC_137/a_36_216# 0.00fF
C20592 NOR2X1_LOC_655/B INVX1_LOC_125/Y 0.19fF
C20593 NOR2X1_LOC_619/A NOR2X1_LOC_188/A 0.06fF
C20594 NOR2X1_LOC_644/A INVX1_LOC_97/A 0.02fF
C20595 INVX1_LOC_64/A NOR2X1_LOC_861/Y 0.10fF
C20596 NOR2X1_LOC_577/Y INVX1_LOC_14/Y 0.10fF
C20597 NOR2X1_LOC_619/A NOR2X1_LOC_548/B 0.01fF
C20598 INVX1_LOC_65/A NOR2X1_LOC_175/A 0.11fF
C20599 INVX1_LOC_90/A NOR2X1_LOC_644/A 0.03fF
C20600 NAND2X1_LOC_562/B NAND2X1_LOC_659/B 0.02fF
C20601 NAND2X1_LOC_724/A NOR2X1_LOC_605/A 0.02fF
C20602 NOR2X1_LOC_249/Y NOR2X1_LOC_33/B 0.05fF
C20603 INVX1_LOC_18/A INVX1_LOC_118/A 0.08fF
C20604 NAND2X1_LOC_366/A VDD -0.00fF
C20605 NAND2X1_LOC_564/B INVX1_LOC_6/A 0.03fF
C20606 INVX1_LOC_254/Y INVX1_LOC_117/A 0.02fF
C20607 NOR2X1_LOC_152/Y NAND2X1_LOC_811/B 0.10fF
C20608 NAND2X1_LOC_466/Y NAND2X1_LOC_453/A 0.04fF
C20609 NOR2X1_LOC_377/Y VDD 0.12fF
C20610 INVX1_LOC_269/A NAND2X1_LOC_82/Y 0.03fF
C20611 NAND2X1_LOC_149/Y INVX1_LOC_114/Y 0.05fF
C20612 NAND2X1_LOC_562/B VDD 0.04fF
C20613 NOR2X1_LOC_482/Y NOR2X1_LOC_253/Y 0.02fF
C20614 INVX1_LOC_136/A INVX1_LOC_307/A 0.07fF
C20615 NAND2X1_LOC_711/B INVX1_LOC_118/A 0.24fF
C20616 NOR2X1_LOC_348/B INVX1_LOC_14/Y 0.01fF
C20617 NOR2X1_LOC_637/Y INVX1_LOC_118/A 0.09fF
C20618 NOR2X1_LOC_558/A NOR2X1_LOC_709/A 0.00fF
C20619 INVX1_LOC_90/A NOR2X1_LOC_751/A 0.04fF
C20620 INVX1_LOC_136/A NOR2X1_LOC_445/B 0.10fF
C20621 NOR2X1_LOC_437/Y INVX1_LOC_54/A 0.07fF
C20622 NOR2X1_LOC_643/A NAND2X1_LOC_207/Y 0.06fF
C20623 INVX1_LOC_224/A INVX1_LOC_29/A 0.01fF
C20624 INVX1_LOC_22/A NOR2X1_LOC_448/A 0.01fF
C20625 NOR2X1_LOC_383/B NOR2X1_LOC_748/A 0.03fF
C20626 INVX1_LOC_172/A INVX1_LOC_118/A 0.03fF
C20627 INVX1_LOC_64/A NOR2X1_LOC_825/a_36_216# 0.00fF
C20628 INVX1_LOC_24/A INVX1_LOC_291/A 0.03fF
C20629 NOR2X1_LOC_441/Y NOR2X1_LOC_653/Y 0.00fF
C20630 NAND2X1_LOC_350/A INVX1_LOC_19/A 0.07fF
C20631 INVX1_LOC_11/A INVX1_LOC_29/A 0.48fF
C20632 NAND2X1_LOC_337/B INVX1_LOC_133/A 0.03fF
C20633 INVX1_LOC_24/A NAND2X1_LOC_802/Y 0.11fF
C20634 INVX1_LOC_279/A NOR2X1_LOC_269/Y 0.90fF
C20635 NOR2X1_LOC_759/Y INVX1_LOC_92/A 0.03fF
C20636 NAND2X1_LOC_701/a_36_24# NAND2X1_LOC_782/B 0.01fF
C20637 INVX1_LOC_89/A INVX1_LOC_48/A 0.49fF
C20638 NAND2X1_LOC_175/Y NOR2X1_LOC_109/Y 0.07fF
C20639 INVX1_LOC_256/Y NAND2X1_LOC_633/Y 0.32fF
C20640 INVX1_LOC_22/A NAND2X1_LOC_212/Y 0.02fF
C20641 NAND2X1_LOC_149/Y NOR2X1_LOC_467/A 0.05fF
C20642 INVX1_LOC_202/A INVX1_LOC_92/A 0.04fF
C20643 INVX1_LOC_218/Y INVX1_LOC_19/A 0.04fF
C20644 NOR2X1_LOC_756/Y INPUT_0 0.05fF
C20645 NAND2X1_LOC_793/B INVX1_LOC_181/A 0.21fF
C20646 NOR2X1_LOC_773/Y VDD 3.27fF
C20647 NOR2X1_LOC_441/Y INVX1_LOC_19/A 0.05fF
C20648 NAND2X1_LOC_369/a_36_24# NOR2X1_LOC_188/A 0.01fF
C20649 NOR2X1_LOC_68/A INVX1_LOC_285/A 0.00fF
C20650 NOR2X1_LOC_68/A INVX1_LOC_265/Y 0.01fF
C20651 NOR2X1_LOC_550/B INVX1_LOC_92/A 0.07fF
C20652 INVX1_LOC_22/A NOR2X1_LOC_853/a_36_216# 0.00fF
C20653 NAND2X1_LOC_96/A NOR2X1_LOC_537/Y 0.07fF
C20654 INVX1_LOC_164/A INVX1_LOC_95/Y 0.07fF
C20655 NAND2X1_LOC_364/A NAND2X1_LOC_475/Y 0.02fF
C20656 NOR2X1_LOC_298/Y INVX1_LOC_11/Y 1.03fF
C20657 NAND2X1_LOC_338/B NAND2X1_LOC_96/A 2.04fF
C20658 INVX1_LOC_103/A NOR2X1_LOC_270/a_36_216# 0.02fF
C20659 NOR2X1_LOC_68/A NOR2X1_LOC_814/A 8.28fF
C20660 NOR2X1_LOC_589/A INVX1_LOC_76/A 0.26fF
C20661 NAND2X1_LOC_67/Y INVX1_LOC_4/A 0.03fF
C20662 INVX1_LOC_161/Y NOR2X1_LOC_48/B 0.03fF
C20663 NOR2X1_LOC_433/A NOR2X1_LOC_58/Y 0.01fF
C20664 INVX1_LOC_23/Y INVX1_LOC_306/Y 0.17fF
C20665 INVX1_LOC_14/Y INVX1_LOC_22/A 0.01fF
C20666 NOR2X1_LOC_369/Y INVX1_LOC_42/A 0.01fF
C20667 NOR2X1_LOC_419/Y NAND2X1_LOC_85/Y 0.02fF
C20668 NAND2X1_LOC_323/B NAND2X1_LOC_96/A 0.14fF
C20669 NOR2X1_LOC_561/Y INVX1_LOC_20/A 0.07fF
C20670 INVX1_LOC_7/A INVX1_LOC_20/A 0.12fF
C20671 NAND2X1_LOC_850/A INVX1_LOC_98/A 0.18fF
C20672 NOR2X1_LOC_372/A NAND2X1_LOC_254/Y 0.01fF
C20673 INVX1_LOC_41/A NOR2X1_LOC_216/B 0.01fF
C20674 INVX1_LOC_229/Y INVX1_LOC_76/A 0.03fF
C20675 NOR2X1_LOC_666/A INVX1_LOC_271/Y 0.07fF
C20676 NAND2X1_LOC_577/A INVX1_LOC_284/A 0.00fF
C20677 NOR2X1_LOC_346/B INVX1_LOC_230/A 0.08fF
C20678 NOR2X1_LOC_540/B INVX1_LOC_97/A 0.02fF
C20679 NOR2X1_LOC_793/Y NOR2X1_LOC_334/Y 1.49fF
C20680 NOR2X1_LOC_91/A INVX1_LOC_21/A 0.05fF
C20681 INVX1_LOC_21/A NOR2X1_LOC_668/Y 0.04fF
C20682 INVX1_LOC_35/A NAND2X1_LOC_9/Y 0.09fF
C20683 INVX1_LOC_249/Y INVX1_LOC_92/A 0.07fF
C20684 INVX1_LOC_286/Y INVX1_LOC_42/A 0.40fF
C20685 INVX1_LOC_50/A INVX1_LOC_50/Y 0.01fF
C20686 NOR2X1_LOC_470/B INVX1_LOC_78/A 0.15fF
C20687 NOR2X1_LOC_181/Y NOR2X1_LOC_155/A 0.01fF
C20688 INVX1_LOC_35/A INVX1_LOC_233/A 0.07fF
C20689 INVX1_LOC_136/A INVX1_LOC_12/A 1.89fF
C20690 INVX1_LOC_182/Y NOR2X1_LOC_269/Y 0.00fF
C20691 INVX1_LOC_17/Y NAND2X1_LOC_778/Y 0.06fF
C20692 NAND2X1_LOC_634/Y NOR2X1_LOC_89/A 0.31fF
C20693 NOR2X1_LOC_389/A D_INPUT_5 0.01fF
C20694 NOR2X1_LOC_237/Y NAND2X1_LOC_489/Y 0.06fF
C20695 NAND2X1_LOC_773/Y INVX1_LOC_26/A 0.01fF
C20696 NOR2X1_LOC_332/A VDD 2.64fF
C20697 NOR2X1_LOC_599/A NOR2X1_LOC_48/B 0.03fF
C20698 NAND2X1_LOC_796/B INVX1_LOC_57/A 0.01fF
C20699 NAND2X1_LOC_708/Y NOR2X1_LOC_53/Y 0.01fF
C20700 INVX1_LOC_21/A INVX1_LOC_23/A 2.90fF
C20701 INVX1_LOC_140/A NOR2X1_LOC_56/Y 0.05fF
C20702 NAND2X1_LOC_807/Y NOR2X1_LOC_279/Y 0.01fF
C20703 INVX1_LOC_298/Y INVX1_LOC_11/A 0.01fF
C20704 INVX1_LOC_266/A INVX1_LOC_50/A 0.07fF
C20705 INVX1_LOC_36/A INVX1_LOC_32/A 0.13fF
C20706 INVX1_LOC_11/A NOR2X1_LOC_281/Y 0.02fF
C20707 NOR2X1_LOC_91/A NOR2X1_LOC_469/a_36_216# 0.00fF
C20708 INVX1_LOC_35/A NOR2X1_LOC_798/A 0.09fF
C20709 NOR2X1_LOC_433/A INVX1_LOC_29/A 0.10fF
C20710 NAND2X1_LOC_559/Y NAND2X1_LOC_725/Y 0.05fF
C20711 INVX1_LOC_2/A NOR2X1_LOC_127/a_36_216# 0.02fF
C20712 INVX1_LOC_18/A INVX1_LOC_257/A 0.07fF
C20713 NOR2X1_LOC_169/B INVX1_LOC_4/A 0.02fF
C20714 NOR2X1_LOC_542/Y INVX1_LOC_117/A 0.07fF
C20715 NOR2X1_LOC_142/Y INVX1_LOC_19/A 0.00fF
C20716 NAND2X1_LOC_477/A NAND2X1_LOC_477/Y 0.07fF
C20717 INVX1_LOC_95/Y NOR2X1_LOC_368/A 0.01fF
C20718 INVX1_LOC_233/Y NOR2X1_LOC_496/Y 0.01fF
C20719 INVX1_LOC_36/A NOR2X1_LOC_329/Y 0.09fF
C20720 NOR2X1_LOC_710/B NOR2X1_LOC_383/B 0.01fF
C20721 NOR2X1_LOC_593/Y INVX1_LOC_29/A 0.02fF
C20722 INVX1_LOC_140/A VDD 3.33fF
C20723 INVX1_LOC_212/Y NOR2X1_LOC_340/A 0.05fF
C20724 INVX1_LOC_45/A INVX1_LOC_94/Y 0.45fF
C20725 NAND2X1_LOC_807/Y NAND2X1_LOC_804/Y 0.02fF
C20726 NAND2X1_LOC_35/Y NOR2X1_LOC_824/A 0.04fF
C20727 INVX1_LOC_140/A NAND2X1_LOC_800/A 0.03fF
C20728 NOR2X1_LOC_360/Y NOR2X1_LOC_38/B 0.03fF
C20729 INVX1_LOC_311/Y INVX1_LOC_117/A 0.05fF
C20730 NOR2X1_LOC_596/A D_INPUT_5 0.01fF
C20731 NAND2X1_LOC_291/a_36_24# INVX1_LOC_37/A 0.00fF
C20732 NAND2X1_LOC_660/Y NAND2X1_LOC_798/B 0.07fF
C20733 NOR2X1_LOC_332/A NOR2X1_LOC_846/a_36_216# 0.01fF
C20734 INVX1_LOC_36/A NAND2X1_LOC_175/Y 0.25fF
C20735 NAND2X1_LOC_35/Y INVX1_LOC_237/A 0.03fF
C20736 NAND2X1_LOC_391/Y INVX1_LOC_13/Y 0.07fF
C20737 NOR2X1_LOC_208/Y INVX1_LOC_32/A 0.03fF
C20738 NAND2X1_LOC_555/Y NAND2X1_LOC_222/a_36_24# 0.01fF
C20739 INVX1_LOC_14/A NOR2X1_LOC_392/Y 0.21fF
C20740 NAND2X1_LOC_463/B VDD 0.91fF
C20741 NOR2X1_LOC_590/A NOR2X1_LOC_831/a_36_216# 0.00fF
C20742 NOR2X1_LOC_74/a_36_216# INVX1_LOC_37/A 0.00fF
C20743 INVX1_LOC_91/A NAND2X1_LOC_655/A 0.01fF
C20744 INVX1_LOC_8/A NOR2X1_LOC_89/A 0.05fF
C20745 NOR2X1_LOC_644/A INVX1_LOC_38/A 0.03fF
C20746 NOR2X1_LOC_272/Y NOR2X1_LOC_791/Y 0.01fF
C20747 NAND2X1_LOC_783/A INVX1_LOC_291/A 0.17fF
C20748 NOR2X1_LOC_52/B INVX1_LOC_29/A 0.10fF
C20749 NOR2X1_LOC_527/Y INVX1_LOC_37/A 0.05fF
C20750 NOR2X1_LOC_130/A INVX1_LOC_291/A 0.46fF
C20751 INVX1_LOC_159/A INVX1_LOC_78/A 0.07fF
C20752 NOR2X1_LOC_655/B INVX1_LOC_19/A 0.08fF
C20753 INVX1_LOC_228/Y NOR2X1_LOC_660/Y 0.09fF
C20754 NAND2X1_LOC_800/Y NAND2X1_LOC_802/Y 0.07fF
C20755 INPUT_3 NOR2X1_LOC_416/A 0.07fF
C20756 NOR2X1_LOC_428/Y INVX1_LOC_23/A 0.07fF
C20757 NOR2X1_LOC_620/Y INVX1_LOC_15/A 0.02fF
C20758 NAND2X1_LOC_374/Y NAND2X1_LOC_500/B 0.04fF
C20759 NAND2X1_LOC_468/B INVX1_LOC_91/A 0.03fF
C20760 NOR2X1_LOC_91/Y NOR2X1_LOC_89/Y 0.08fF
C20761 NOR2X1_LOC_171/Y NOR2X1_LOC_331/B 0.06fF
C20762 INVX1_LOC_72/A NAND2X1_LOC_99/A 0.00fF
C20763 INVX1_LOC_90/A NAND2X1_LOC_243/Y 0.10fF
C20764 INVX1_LOC_45/A INVX1_LOC_296/A 0.04fF
C20765 INVX1_LOC_5/A NOR2X1_LOC_361/B 0.01fF
C20766 NOR2X1_LOC_191/B INVX1_LOC_78/A 0.01fF
C20767 INVX1_LOC_10/A NOR2X1_LOC_117/a_36_216# 0.00fF
C20768 INVX1_LOC_71/A INVX1_LOC_94/Y 0.01fF
C20769 NOR2X1_LOC_790/B INVX1_LOC_292/A 0.95fF
C20770 NOR2X1_LOC_595/Y NAND2X1_LOC_655/B 0.05fF
C20771 NOR2X1_LOC_837/A INVX1_LOC_37/A 0.01fF
C20772 NAND2X1_LOC_571/Y INVX1_LOC_237/A 0.02fF
C20773 NAND2X1_LOC_330/a_36_24# INVX1_LOC_94/Y 0.01fF
C20774 INVX1_LOC_13/A INVX1_LOC_63/A 0.14fF
C20775 INVX1_LOC_223/A INVX1_LOC_270/Y 0.14fF
C20776 INVX1_LOC_64/A NOR2X1_LOC_331/Y 0.05fF
C20777 NOR2X1_LOC_309/Y INVX1_LOC_32/A 0.01fF
C20778 INVX1_LOC_235/A INVX1_LOC_14/A 0.04fF
C20779 INVX1_LOC_235/Y INVX1_LOC_1/A 0.01fF
C20780 NOR2X1_LOC_724/Y NOR2X1_LOC_155/A 0.11fF
C20781 NOR2X1_LOC_570/a_36_216# NOR2X1_LOC_383/B 0.00fF
C20782 NOR2X1_LOC_285/Y NOR2X1_LOC_160/B 0.06fF
C20783 NAND2X1_LOC_149/Y INVX1_LOC_1/A 0.07fF
C20784 NOR2X1_LOC_594/Y NOR2X1_LOC_331/B 0.19fF
C20785 INVX1_LOC_22/A NOR2X1_LOC_831/Y 0.52fF
C20786 NAND2X1_LOC_354/Y INVX1_LOC_23/A 0.03fF
C20787 INVX1_LOC_71/A INVX1_LOC_181/A 0.75fF
C20788 NOR2X1_LOC_824/Y INVX1_LOC_20/A 0.08fF
C20789 INVX1_LOC_52/Y NOR2X1_LOC_205/Y -0.00fF
C20790 NAND2X1_LOC_30/Y D_INPUT_6 0.99fF
C20791 NOR2X1_LOC_510/Y NOR2X1_LOC_816/A 0.03fF
C20792 INVX1_LOC_295/A NOR2X1_LOC_450/B -0.03fF
C20793 INVX1_LOC_147/Y INVX1_LOC_76/A 0.01fF
C20794 NAND2X1_LOC_622/B NOR2X1_LOC_629/Y 0.02fF
C20795 NOR2X1_LOC_246/A INVX1_LOC_63/A 0.10fF
C20796 NAND2X1_LOC_577/A NOR2X1_LOC_663/A 0.06fF
C20797 NAND2X1_LOC_348/A NOR2X1_LOC_61/A 0.02fF
C20798 INVX1_LOC_208/A NAND2X1_LOC_792/B 0.01fF
C20799 INVX1_LOC_20/A INVX1_LOC_76/A 0.23fF
C20800 NOR2X1_LOC_516/Y NOR2X1_LOC_415/Y 0.09fF
C20801 NOR2X1_LOC_82/A NAND2X1_LOC_347/B 0.04fF
C20802 NOR2X1_LOC_99/B INVX1_LOC_19/A 0.07fF
C20803 NOR2X1_LOC_19/B NAND2X1_LOC_574/A 0.45fF
C20804 INVX1_LOC_133/Y NOR2X1_LOC_334/Y 0.02fF
C20805 INVX1_LOC_21/A INVX1_LOC_31/A 0.24fF
C20806 NAND2X1_LOC_640/Y NAND2X1_LOC_442/a_36_24# 0.00fF
C20807 NOR2X1_LOC_392/B INVX1_LOC_16/Y 0.10fF
C20808 NOR2X1_LOC_848/Y INVX1_LOC_17/A 2.07fF
C20809 NOR2X1_LOC_683/a_36_216# INVX1_LOC_117/A 0.01fF
C20810 INVX1_LOC_299/A NOR2X1_LOC_541/Y 0.01fF
C20811 NOR2X1_LOC_361/B NAND2X1_LOC_337/B 0.11fF
C20812 NOR2X1_LOC_272/Y INVX1_LOC_30/A 0.00fF
C20813 NOR2X1_LOC_91/A NAND2X1_LOC_785/Y 0.03fF
C20814 INVX1_LOC_186/A INVX1_LOC_274/A 0.07fF
C20815 NOR2X1_LOC_554/B INVX1_LOC_38/Y 0.63fF
C20816 INPUT_6 INVX1_LOC_77/A 0.23fF
C20817 NAND2X1_LOC_140/A NOR2X1_LOC_89/A 0.00fF
C20818 NOR2X1_LOC_550/B INVX1_LOC_53/A 0.15fF
C20819 NOR2X1_LOC_74/A INVX1_LOC_220/A 0.15fF
C20820 INVX1_LOC_27/A NOR2X1_LOC_723/a_36_216# 0.01fF
C20821 NOR2X1_LOC_647/A NOR2X1_LOC_818/Y 0.21fF
C20822 INVX1_LOC_224/Y NOR2X1_LOC_315/Y 0.79fF
C20823 INVX1_LOC_2/A NOR2X1_LOC_658/a_36_216# 0.00fF
C20824 NAND2X1_LOC_338/B NAND2X1_LOC_99/A 0.28fF
C20825 INVX1_LOC_299/A INVX1_LOC_45/A 0.03fF
C20826 NOR2X1_LOC_32/B INVX1_LOC_34/A 0.50fF
C20827 INVX1_LOC_103/A INVX1_LOC_81/Y 0.01fF
C20828 NOR2X1_LOC_493/B NOR2X1_LOC_383/B 0.01fF
C20829 NAND2X1_LOC_385/a_36_24# NOR2X1_LOC_593/Y 0.00fF
C20830 INVX1_LOC_217/Y NOR2X1_LOC_392/Y 0.02fF
C20831 NOR2X1_LOC_91/A NOR2X1_LOC_667/A 0.24fF
C20832 INVX1_LOC_299/A NOR2X1_LOC_568/A 0.08fF
C20833 NOR2X1_LOC_320/Y INVX1_LOC_63/A 0.03fF
C20834 INVX1_LOC_7/A INVX1_LOC_4/A 0.05fF
C20835 NOR2X1_LOC_91/A INVX1_LOC_248/A 0.01fF
C20836 INVX1_LOC_255/Y NAND2X1_LOC_223/A 0.07fF
C20837 NAND2X1_LOC_182/A NAND2X1_LOC_860/A 0.11fF
C20838 INVX1_LOC_10/A NAND2X1_LOC_647/B 0.02fF
C20839 INVX1_LOC_298/A INVX1_LOC_49/A 0.01fF
C20840 INVX1_LOC_31/Y NAND2X1_LOC_63/Y 0.09fF
C20841 D_INPUT_0 INVX1_LOC_47/Y 0.01fF
C20842 NOR2X1_LOC_441/Y INVX1_LOC_161/Y 0.02fF
C20843 INVX1_LOC_77/A NOR2X1_LOC_849/A 0.02fF
C20844 NOR2X1_LOC_799/a_36_216# INVX1_LOC_58/Y 0.01fF
C20845 NOR2X1_LOC_189/A NAND2X1_LOC_794/B 0.02fF
C20846 NOR2X1_LOC_486/Y INVX1_LOC_179/A 0.03fF
C20847 NOR2X1_LOC_657/B NOR2X1_LOC_155/A 0.05fF
C20848 NOR2X1_LOC_604/Y NOR2X1_LOC_423/Y 0.01fF
C20849 NOR2X1_LOC_315/Y NAND2X1_LOC_793/B 0.01fF
C20850 NAND2X1_LOC_721/B INVX1_LOC_11/A 0.00fF
C20851 NAND2X1_LOC_785/A NAND2X1_LOC_787/A 0.00fF
C20852 NOR2X1_LOC_296/Y INVX1_LOC_36/A 0.08fF
C20853 INVX1_LOC_5/A INVX1_LOC_153/Y 0.10fF
C20854 INVX1_LOC_64/A NOR2X1_LOC_367/B 0.15fF
C20855 NOR2X1_LOC_427/a_36_216# INVX1_LOC_72/A 0.00fF
C20856 NAND2X1_LOC_560/A NAND2X1_LOC_254/Y 0.02fF
C20857 NOR2X1_LOC_567/a_36_216# NOR2X1_LOC_640/Y 0.00fF
C20858 INVX1_LOC_41/A INVX1_LOC_93/A 0.07fF
C20859 NOR2X1_LOC_456/Y NOR2X1_LOC_78/B 0.16fF
C20860 NOR2X1_LOC_500/A INVX1_LOC_24/Y 0.23fF
C20861 NAND2X1_LOC_834/a_36_24# INVX1_LOC_57/A 0.01fF
C20862 INVX1_LOC_36/A INPUT_3 0.07fF
C20863 NOR2X1_LOC_598/B NOR2X1_LOC_778/B 0.03fF
C20864 INVX1_LOC_258/Y INVX1_LOC_237/Y 0.00fF
C20865 NOR2X1_LOC_321/Y INVX1_LOC_49/A 0.08fF
C20866 NAND2X1_LOC_803/B NOR2X1_LOC_68/A 0.01fF
C20867 NOR2X1_LOC_604/Y NOR2X1_LOC_222/Y 0.03fF
C20868 NAND2X1_LOC_358/Y INVX1_LOC_26/Y 0.06fF
C20869 NOR2X1_LOC_405/A NAND2X1_LOC_475/Y 0.01fF
C20870 NOR2X1_LOC_441/Y INVX1_LOC_312/A 0.06fF
C20871 NAND2X1_LOC_577/A NAND2X1_LOC_136/a_36_24# 0.01fF
C20872 INVX1_LOC_278/A NAND2X1_LOC_181/Y 0.01fF
C20873 INVX1_LOC_50/A INVX1_LOC_30/Y 0.17fF
C20874 INVX1_LOC_41/A NAND2X1_LOC_513/B 0.01fF
C20875 INVX1_LOC_5/A INVX1_LOC_177/A 0.03fF
C20876 INVX1_LOC_25/A INVX1_LOC_16/A 10.19fF
C20877 INVX1_LOC_97/Y NOR2X1_LOC_778/B 0.01fF
C20878 NOR2X1_LOC_309/Y INVX1_LOC_171/Y 0.01fF
C20879 INVX1_LOC_93/A NAND2X1_LOC_477/A 0.10fF
C20880 NOR2X1_LOC_470/B INVX1_LOC_113/Y 0.00fF
C20881 INVX1_LOC_64/A INVX1_LOC_179/Y 0.09fF
C20882 INVX1_LOC_136/A NAND2X1_LOC_733/Y 0.03fF
C20883 NOR2X1_LOC_112/a_36_216# NOR2X1_LOC_865/Y 0.00fF
C20884 INVX1_LOC_45/A NOR2X1_LOC_524/Y 0.17fF
C20885 NAND2X1_LOC_354/Y INVX1_LOC_31/A 0.00fF
C20886 NOR2X1_LOC_99/B INVX1_LOC_26/Y 0.12fF
C20887 NOR2X1_LOC_590/A NOR2X1_LOC_68/A 0.30fF
C20888 NOR2X1_LOC_824/A NOR2X1_LOC_234/Y 0.08fF
C20889 NOR2X1_LOC_521/Y INVX1_LOC_23/A 0.01fF
C20890 INVX1_LOC_5/A INVX1_LOC_280/Y 0.04fF
C20891 NOR2X1_LOC_122/A NOR2X1_LOC_142/Y 0.01fF
C20892 NOR2X1_LOC_731/Y INVX1_LOC_213/A 0.04fF
C20893 NOR2X1_LOC_706/a_36_216# NAND2X1_LOC_425/Y 0.01fF
C20894 INVX1_LOC_150/A NOR2X1_LOC_383/B 0.02fF
C20895 INPUT_0 NOR2X1_LOC_620/A 0.01fF
C20896 INVX1_LOC_21/A NOR2X1_LOC_290/Y 0.01fF
C20897 INVX1_LOC_39/A INVX1_LOC_34/Y 0.02fF
C20898 NOR2X1_LOC_205/Y INVX1_LOC_63/Y 0.01fF
C20899 NAND2X1_LOC_364/A INVX1_LOC_30/A 0.23fF
C20900 INVX1_LOC_2/A D_INPUT_6 0.01fF
C20901 INVX1_LOC_21/A INVX1_LOC_191/Y 0.11fF
C20902 INVX1_LOC_89/A NOR2X1_LOC_383/B 0.09fF
C20903 NAND2X1_LOC_642/Y NAND2X1_LOC_207/B 0.01fF
C20904 INVX1_LOC_224/A INVX1_LOC_8/A 0.03fF
C20905 INVX1_LOC_48/Y NOR2X1_LOC_84/Y 0.06fF
C20906 NOR2X1_LOC_356/A NAND2X1_LOC_72/a_36_24# 0.00fF
C20907 INVX1_LOC_136/A INVX1_LOC_217/A 0.17fF
C20908 NAND2X1_LOC_564/B NOR2X1_LOC_109/Y 0.00fF
C20909 NAND2X1_LOC_840/B NOR2X1_LOC_406/A 0.00fF
C20910 INVX1_LOC_2/A NOR2X1_LOC_321/Y 0.28fF
C20911 INVX1_LOC_11/A INVX1_LOC_8/A 0.07fF
C20912 INVX1_LOC_64/A NOR2X1_LOC_561/Y 0.22fF
C20913 INVX1_LOC_74/A INVX1_LOC_29/A 0.00fF
C20914 INVX1_LOC_286/Y NOR2X1_LOC_152/Y 0.11fF
C20915 NOR2X1_LOC_524/Y INVX1_LOC_71/A 0.02fF
C20916 D_INPUT_1 NOR2X1_LOC_76/A 1.05fF
C20917 NOR2X1_LOC_721/Y INVX1_LOC_78/A 0.03fF
C20918 INVX1_LOC_84/A INVX1_LOC_117/A 0.10fF
C20919 INVX1_LOC_14/Y INVX1_LOC_186/Y 0.10fF
C20920 INVX1_LOC_269/A NOR2X1_LOC_168/B 0.01fF
C20921 NOR2X1_LOC_103/Y NOR2X1_LOC_315/Y 0.00fF
C20922 NOR2X1_LOC_602/B NOR2X1_LOC_841/A 0.06fF
C20923 NAND2X1_LOC_725/B NAND2X1_LOC_374/Y 0.19fF
C20924 NAND2X1_LOC_348/A INVX1_LOC_16/Y 0.00fF
C20925 INVX1_LOC_62/Y NOR2X1_LOC_360/Y 0.07fF
C20926 INVX1_LOC_102/Y INVX1_LOC_181/A 0.00fF
C20927 INVX1_LOC_280/Y NOR2X1_LOC_494/Y 0.03fF
C20928 NOR2X1_LOC_56/Y INVX1_LOC_42/A 0.09fF
C20929 NOR2X1_LOC_9/Y NAND2X1_LOC_447/a_36_24# 0.00fF
C20930 INVX1_LOC_77/A INVX1_LOC_142/A 0.23fF
C20931 NOR2X1_LOC_859/A INVX1_LOC_77/A 0.03fF
C20932 NOR2X1_LOC_841/A INVX1_LOC_54/A 0.10fF
C20933 VDD INVX1_LOC_263/Y 0.41fF
C20934 NOR2X1_LOC_114/a_36_216# NOR2X1_LOC_814/A 0.00fF
C20935 NAND2X1_LOC_705/Y INVX1_LOC_22/A 0.01fF
C20936 NOR2X1_LOC_614/a_36_216# NOR2X1_LOC_542/Y 0.00fF
C20937 NOR2X1_LOC_361/B NOR2X1_LOC_773/Y 0.27fF
C20938 INVX1_LOC_159/A NOR2X1_LOC_152/Y 0.07fF
C20939 INVX1_LOC_35/A NAND2X1_LOC_842/B 0.01fF
C20940 INVX1_LOC_1/A INVX1_LOC_16/A 1.06fF
C20941 NOR2X1_LOC_723/Y INVX1_LOC_63/Y 0.11fF
C20942 NAND2X1_LOC_303/Y INVX1_LOC_22/A 0.16fF
C20943 INVX1_LOC_14/A INVX1_LOC_25/Y 0.44fF
C20944 NOR2X1_LOC_226/A NAND2X1_LOC_793/Y 0.10fF
C20945 D_INPUT_1 INVX1_LOC_73/A 0.07fF
C20946 NAND2X1_LOC_348/A NAND2X1_LOC_205/A 0.00fF
C20947 NAND2X1_LOC_193/a_36_24# INVX1_LOC_159/A 0.00fF
C20948 NOR2X1_LOC_815/Y INVX1_LOC_18/A 0.02fF
C20949 VDD INVX1_LOC_42/A 3.93fF
C20950 NAND2X1_LOC_571/Y INVX1_LOC_234/A 0.10fF
C20951 INVX1_LOC_144/A INVX1_LOC_271/A 0.01fF
C20952 NAND2X1_LOC_51/B INVX1_LOC_23/A 0.01fF
C20953 INVX1_LOC_280/Y NOR2X1_LOC_816/A 0.03fF
C20954 NAND2X1_LOC_800/A INVX1_LOC_42/A 0.06fF
C20955 NOR2X1_LOC_82/A NOR2X1_LOC_382/a_36_216# 0.00fF
C20956 INVX1_LOC_45/A NOR2X1_LOC_315/Y 0.08fF
C20957 NOR2X1_LOC_825/Y INVX1_LOC_3/Y 0.03fF
C20958 INVX1_LOC_58/A NOR2X1_LOC_335/B 0.05fF
C20959 NOR2X1_LOC_15/Y NAND2X1_LOC_319/A 0.00fF
C20960 NOR2X1_LOC_703/Y NOR2X1_LOC_383/B 0.29fF
C20961 INVX1_LOC_214/A INVX1_LOC_31/A 0.15fF
C20962 INVX1_LOC_21/A INVX1_LOC_313/A 0.24fF
C20963 INVX1_LOC_45/Y INVX1_LOC_33/A 0.01fF
C20964 NAND2X1_LOC_785/A INVX1_LOC_30/A 0.20fF
C20965 NOR2X1_LOC_106/Y NOR2X1_LOC_577/Y 0.02fF
C20966 NOR2X1_LOC_667/A INVX1_LOC_31/A 0.07fF
C20967 INVX1_LOC_76/A INVX1_LOC_4/A 0.09fF
C20968 NAND2X1_LOC_220/B INVX1_LOC_117/A 0.01fF
C20969 NAND2X1_LOC_854/B NAND2X1_LOC_537/Y 0.38fF
C20970 INVX1_LOC_304/Y INVX1_LOC_136/A 0.07fF
C20971 INVX1_LOC_47/Y NOR2X1_LOC_266/B 0.09fF
C20972 NOR2X1_LOC_52/B NAND2X1_LOC_634/Y 0.01fF
C20973 INVX1_LOC_248/A INVX1_LOC_31/A 0.07fF
C20974 INVX1_LOC_41/A NOR2X1_LOC_500/A 0.10fF
C20975 INVX1_LOC_102/A NOR2X1_LOC_536/A 0.07fF
C20976 INVX1_LOC_78/A NOR2X1_LOC_56/Y 0.03fF
C20977 NOR2X1_LOC_32/B INPUT_0 0.01fF
C20978 INVX1_LOC_269/A NAND2X1_LOC_656/Y 0.07fF
C20979 NOR2X1_LOC_329/B NOR2X1_LOC_674/Y 0.30fF
C20980 INVX1_LOC_283/Y INVX1_LOC_113/Y -0.00fF
C20981 INVX1_LOC_2/Y NAND2X1_LOC_296/a_36_24# 0.00fF
C20982 INVX1_LOC_50/A INVX1_LOC_96/A 0.06fF
C20983 NOR2X1_LOC_471/Y NAND2X1_LOC_479/Y 0.09fF
C20984 NAND2X1_LOC_11/Y INVX1_LOC_30/A 0.02fF
C20985 NOR2X1_LOC_89/A INVX1_LOC_118/Y 0.02fF
C20986 INVX1_LOC_98/A INVX1_LOC_57/A 0.07fF
C20987 INVX1_LOC_21/A NAND2X1_LOC_807/Y 0.07fF
C20988 INVX1_LOC_78/A NOR2X1_LOC_136/a_36_216# 0.00fF
C20989 NOR2X1_LOC_334/A INVX1_LOC_53/A 0.03fF
C20990 INVX1_LOC_117/A INVX1_LOC_15/A 0.29fF
C20991 NAND2X1_LOC_763/B NAND2X1_LOC_11/Y 0.16fF
C20992 NOR2X1_LOC_78/A INVX1_LOC_57/A 0.17fF
C20993 INVX1_LOC_73/A NOR2X1_LOC_652/Y 0.07fF
C20994 NOR2X1_LOC_91/A INVX1_LOC_304/A 0.07fF
C20995 INVX1_LOC_17/A INVX1_LOC_135/A 0.12fF
C20996 NAND2X1_LOC_337/B NAND2X1_LOC_573/A 0.01fF
C20997 INVX1_LOC_181/Y NOR2X1_LOC_709/A 0.01fF
C20998 NOR2X1_LOC_222/Y INVX1_LOC_72/A 0.03fF
C20999 INVX1_LOC_216/Y D_INPUT_0 0.01fF
C21000 INVX1_LOC_132/A NOR2X1_LOC_264/Y 0.02fF
C21001 INVX1_LOC_206/A INVX1_LOC_94/A 0.02fF
C21002 INVX1_LOC_136/A NOR2X1_LOC_566/Y 0.06fF
C21003 VDD INVX1_LOC_78/A 2.73fF
C21004 INVX1_LOC_13/A NOR2X1_LOC_606/a_36_216# 0.00fF
C21005 INVX1_LOC_201/Y NAND2X1_LOC_5/a_36_24# 0.01fF
C21006 INVX1_LOC_310/Y NOR2X1_LOC_285/B 0.02fF
C21007 INVX1_LOC_41/A NOR2X1_LOC_254/Y 0.03fF
C21008 INVX1_LOC_5/A INVX1_LOC_285/Y 0.07fF
C21009 INVX1_LOC_34/A NOR2X1_LOC_364/Y 0.01fF
C21010 NOR2X1_LOC_220/A NOR2X1_LOC_360/Y 0.01fF
C21011 NAND2X1_LOC_338/B NAND2X1_LOC_656/A 0.01fF
C21012 NOR2X1_LOC_273/Y NOR2X1_LOC_78/B 0.01fF
C21013 INVX1_LOC_30/A NOR2X1_LOC_86/A 0.01fF
C21014 NOR2X1_LOC_384/Y INVX1_LOC_16/A 0.42fF
C21015 NOR2X1_LOC_78/B NOR2X1_LOC_759/Y 0.03fF
C21016 INVX1_LOC_38/A INVX1_LOC_21/Y 0.03fF
C21017 NOR2X1_LOC_369/Y NAND2X1_LOC_861/Y 0.04fF
C21018 NAND2X1_LOC_555/Y INVX1_LOC_135/A 1.40fF
C21019 INVX1_LOC_288/A VDD 0.12fF
C21020 INVX1_LOC_226/Y NOR2X1_LOC_791/a_36_216# 0.00fF
C21021 INVX1_LOC_208/A NOR2X1_LOC_359/Y -0.03fF
C21022 NOR2X1_LOC_65/B VDD 1.34fF
C21023 INVX1_LOC_18/A NAND2X1_LOC_735/B 0.00fF
C21024 NOR2X1_LOC_52/B INVX1_LOC_8/A 0.02fF
C21025 INVX1_LOC_21/A INVX1_LOC_6/A 0.13fF
C21026 NOR2X1_LOC_772/B INVX1_LOC_91/A 0.05fF
C21027 NOR2X1_LOC_242/A NOR2X1_LOC_334/A 0.51fF
C21028 NOR2X1_LOC_78/B NOR2X1_LOC_550/B 0.03fF
C21029 NAND2X1_LOC_30/Y NOR2X1_LOC_163/a_36_216# 0.00fF
C21030 INVX1_LOC_14/A INVX1_LOC_75/A 0.28fF
C21031 NOR2X1_LOC_277/a_36_216# INVX1_LOC_304/A 0.01fF
C21032 INVX1_LOC_18/A NOR2X1_LOC_302/a_36_216# 0.00fF
C21033 INVX1_LOC_41/A INVX1_LOC_54/Y 0.00fF
C21034 NAND2X1_LOC_357/B INVX1_LOC_240/A 0.02fF
C21035 NOR2X1_LOC_681/Y NOR2X1_LOC_654/A 0.10fF
C21036 NOR2X1_LOC_843/A NOR2X1_LOC_175/A 0.01fF
C21037 INVX1_LOC_58/A NOR2X1_LOC_825/Y 0.01fF
C21038 INVX1_LOC_18/A INPUT_5 0.52fF
C21039 INVX1_LOC_32/A NOR2X1_LOC_435/A 0.03fF
C21040 INVX1_LOC_37/A NOR2X1_LOC_654/A 0.13fF
C21041 NOR2X1_LOC_334/Y NOR2X1_LOC_729/A 0.00fF
C21042 INVX1_LOC_26/A NOR2X1_LOC_98/B 0.01fF
C21043 NOR2X1_LOC_303/Y NOR2X1_LOC_211/A 0.08fF
C21044 INVX1_LOC_13/Y INVX1_LOC_91/A 0.25fF
C21045 NOR2X1_LOC_561/Y INVX1_LOC_130/Y 0.02fF
C21046 NOR2X1_LOC_632/Y INVX1_LOC_24/A 0.03fF
C21047 NOR2X1_LOC_433/A INVX1_LOC_151/Y 0.02fF
C21048 INVX1_LOC_136/A NAND2X1_LOC_808/A 0.00fF
C21049 NOR2X1_LOC_88/Y INVX1_LOC_3/Y 0.15fF
C21050 INVX1_LOC_269/A NAND2X1_LOC_622/B 0.01fF
C21051 INVX1_LOC_27/A NOR2X1_LOC_845/A 0.04fF
C21052 NOR2X1_LOC_197/A NOR2X1_LOC_197/Y 0.00fF
C21053 NOR2X1_LOC_520/B INVX1_LOC_218/A 0.04fF
C21054 NOR2X1_LOC_68/A NOR2X1_LOC_763/Y 0.01fF
C21055 NAND2X1_LOC_564/B NOR2X1_LOC_237/Y 0.01fF
C21056 NAND2X1_LOC_635/a_36_24# INVX1_LOC_296/A 0.00fF
C21057 NOR2X1_LOC_98/a_36_216# INVX1_LOC_57/A 0.00fF
C21058 INVX1_LOC_70/Y NAND2X1_LOC_474/Y 0.12fF
C21059 INVX1_LOC_64/A INVX1_LOC_76/A 0.31fF
C21060 NAND2X1_LOC_785/A NAND2X1_LOC_722/A 0.02fF
C21061 NOR2X1_LOC_843/B INVX1_LOC_230/A 1.16fF
C21062 INVX1_LOC_172/A NAND2X1_LOC_735/B 0.00fF
C21063 NOR2X1_LOC_78/B INVX1_LOC_249/Y 0.01fF
C21064 NOR2X1_LOC_89/A NOR2X1_LOC_258/Y 0.08fF
C21065 INVX1_LOC_280/Y NAND2X1_LOC_562/B 0.00fF
C21066 INVX1_LOC_37/A INVX1_LOC_58/Y 0.07fF
C21067 NOR2X1_LOC_218/A INPUT_0 0.11fF
C21068 INVX1_LOC_163/A INVX1_LOC_167/Y 0.17fF
C21069 INVX1_LOC_152/Y VDD 0.27fF
C21070 GATE_811 NAND2X1_LOC_853/Y 0.03fF
C21071 NAND2X1_LOC_812/a_36_24# NAND2X1_LOC_852/Y 0.07fF
C21072 INVX1_LOC_90/A NAND2X1_LOC_342/a_36_24# 0.00fF
C21073 INVX1_LOC_88/A NOR2X1_LOC_114/A 0.13fF
C21074 NOR2X1_LOC_261/Y INVX1_LOC_117/A 0.27fF
C21075 NOR2X1_LOC_690/A INVX1_LOC_22/A 0.04fF
C21076 INVX1_LOC_215/A NOR2X1_LOC_172/Y 0.04fF
C21077 NOR2X1_LOC_459/B NOR2X1_LOC_375/Y 0.11fF
C21078 INVX1_LOC_84/A INVX1_LOC_3/Y 0.35fF
C21079 NAND2X1_LOC_466/Y INVX1_LOC_22/A 0.01fF
C21080 NOR2X1_LOC_393/a_36_216# INVX1_LOC_30/A 0.00fF
C21081 NOR2X1_LOC_850/B INVX1_LOC_19/A 0.15fF
C21082 NOR2X1_LOC_52/B NOR2X1_LOC_315/a_36_216# 0.01fF
C21083 INVX1_LOC_32/A INVX1_LOC_63/A 0.26fF
C21084 INVX1_LOC_88/A INVX1_LOC_91/A 0.15fF
C21085 INVX1_LOC_26/Y NOR2X1_LOC_622/a_36_216# 0.00fF
C21086 NOR2X1_LOC_194/Y INVX1_LOC_22/A 0.20fF
C21087 NOR2X1_LOC_274/Y INVX1_LOC_171/A 0.02fF
C21088 NOR2X1_LOC_788/B INVX1_LOC_24/A 0.00fF
C21089 NAND2X1_LOC_564/B NOR2X1_LOC_309/Y 0.10fF
C21090 NAND2X1_LOC_254/Y INVX1_LOC_29/A 0.03fF
C21091 INVX1_LOC_83/A NOR2X1_LOC_550/B 0.01fF
C21092 INVX1_LOC_64/A NAND2X1_LOC_418/a_36_24# 0.00fF
C21093 NOR2X1_LOC_180/a_36_216# INVX1_LOC_30/A 0.02fF
C21094 NOR2X1_LOC_433/A NAND2X1_LOC_140/A 0.04fF
C21095 NOR2X1_LOC_68/A NOR2X1_LOC_703/A 0.18fF
C21096 INVX1_LOC_280/Y NOR2X1_LOC_773/Y 0.16fF
C21097 INVX1_LOC_54/Y NOR2X1_LOC_211/A 0.33fF
C21098 NAND2X1_LOC_374/a_36_24# INPUT_1 0.01fF
C21099 INVX1_LOC_154/A NOR2X1_LOC_345/A 0.04fF
C21100 INVX1_LOC_159/A NAND2X1_LOC_661/A 0.01fF
C21101 INVX1_LOC_33/A NOR2X1_LOC_71/Y 0.09fF
C21102 NOR2X1_LOC_215/A VDD 0.07fF
C21103 NOR2X1_LOC_865/Y NOR2X1_LOC_342/B 0.03fF
C21104 NOR2X1_LOC_175/B NAND2X1_LOC_173/a_36_24# 0.00fF
C21105 INVX1_LOC_1/A NOR2X1_LOC_35/Y 0.10fF
C21106 INVX1_LOC_179/A NOR2X1_LOC_748/A 0.07fF
C21107 NOR2X1_LOC_437/a_36_216# INVX1_LOC_182/Y 0.00fF
C21108 INVX1_LOC_161/Y INVX1_LOC_291/Y 0.99fF
C21109 INVX1_LOC_77/A NOR2X1_LOC_535/a_36_216# 0.00fF
C21110 INVX1_LOC_271/A NOR2X1_LOC_155/A 0.03fF
C21111 NOR2X1_LOC_389/A NOR2X1_LOC_269/Y 0.10fF
C21112 NAND2X1_LOC_175/Y INVX1_LOC_63/A 0.08fF
C21113 INVX1_LOC_49/A INVX1_LOC_148/A 0.07fF
C21114 INVX1_LOC_105/Y NOR2X1_LOC_155/A 0.01fF
C21115 NOR2X1_LOC_644/A INVX1_LOC_33/A 0.03fF
C21116 INVX1_LOC_90/A NOR2X1_LOC_570/B 0.08fF
C21117 INVX1_LOC_259/Y INVX1_LOC_92/A 0.02fF
C21118 NOR2X1_LOC_315/Y NOR2X1_LOC_123/B 0.01fF
C21119 INVX1_LOC_255/Y INVX1_LOC_40/A 0.09fF
C21120 NAND2X1_LOC_647/B INVX1_LOC_12/A 0.08fF
C21121 INVX1_LOC_58/A NOR2X1_LOC_88/Y 0.10fF
C21122 NOR2X1_LOC_503/Y NOR2X1_LOC_56/Y 0.03fF
C21123 NAND2X1_LOC_561/B INVX1_LOC_46/A 0.01fF
C21124 INVX1_LOC_78/A INVX1_LOC_133/A 0.00fF
C21125 NAND2X1_LOC_341/A INVX1_LOC_268/A 0.01fF
C21126 NOR2X1_LOC_828/B INVX1_LOC_33/A 0.07fF
C21127 NOR2X1_LOC_808/A NOR2X1_LOC_326/Y 0.01fF
C21128 INVX1_LOC_304/Y NAND2X1_LOC_862/Y 0.06fF
C21129 NOR2X1_LOC_500/B INVX1_LOC_91/A 0.02fF
C21130 INVX1_LOC_61/Y NOR2X1_LOC_124/A 0.02fF
C21131 NOR2X1_LOC_151/Y NOR2X1_LOC_730/a_36_216# 0.02fF
C21132 NOR2X1_LOC_757/A NOR2X1_LOC_757/Y 0.03fF
C21133 NOR2X1_LOC_773/Y NAND2X1_LOC_573/A 0.14fF
C21134 NOR2X1_LOC_794/B NOR2X1_LOC_35/Y 0.03fF
C21135 NOR2X1_LOC_785/A INVX1_LOC_143/Y 0.28fF
C21136 INVX1_LOC_35/A NOR2X1_LOC_146/a_36_216# 0.00fF
C21137 INVX1_LOC_30/A NOR2X1_LOC_405/A 0.25fF
C21138 INVX1_LOC_221/A INVX1_LOC_28/A 0.03fF
C21139 INVX1_LOC_89/A NOR2X1_LOC_168/A 0.01fF
C21140 INVX1_LOC_3/Y INVX1_LOC_15/A 0.55fF
C21141 INVX1_LOC_58/A INVX1_LOC_84/A 0.69fF
C21142 NOR2X1_LOC_624/A INVX1_LOC_31/Y 0.09fF
C21143 INVX1_LOC_31/A NOR2X1_LOC_670/Y 0.09fF
C21144 NOR2X1_LOC_503/Y VDD 0.44fF
C21145 NOR2X1_LOC_75/Y INVX1_LOC_37/A 0.01fF
C21146 INVX1_LOC_104/A NOR2X1_LOC_569/a_36_216# 0.00fF
C21147 NOR2X1_LOC_65/B INVX1_LOC_133/A 0.12fF
C21148 NOR2X1_LOC_622/A INVX1_LOC_63/A 0.08fF
C21149 NOR2X1_LOC_471/Y INVX1_LOC_139/Y 0.02fF
C21150 INVX1_LOC_227/A NOR2X1_LOC_570/Y 0.01fF
C21151 NOR2X1_LOC_170/a_36_216# INVX1_LOC_91/A 0.01fF
C21152 INVX1_LOC_36/A NOR2X1_LOC_279/Y 0.00fF
C21153 NAND2X1_LOC_799/a_36_24# INVX1_LOC_140/A 0.07fF
C21154 NOR2X1_LOC_103/Y NAND2X1_LOC_93/a_36_24# 0.00fF
C21155 INVX1_LOC_17/A INVX1_LOC_280/A 0.14fF
C21156 INVX1_LOC_36/A NOR2X1_LOC_173/a_36_216# 0.02fF
C21157 NOR2X1_LOC_667/A NAND2X1_LOC_807/Y 1.23fF
C21158 NOR2X1_LOC_720/B INPUT_0 0.00fF
C21159 INVX1_LOC_18/A NAND2X1_LOC_212/Y 0.02fF
C21160 INVX1_LOC_27/A NOR2X1_LOC_155/A 12.72fF
C21161 INVX1_LOC_30/A NOR2X1_LOC_857/A 0.09fF
C21162 NOR2X1_LOC_844/Y VDD 0.00fF
C21163 INVX1_LOC_303/A INVX1_LOC_91/A 0.07fF
C21164 D_INPUT_4 INVX1_LOC_192/Y 0.24fF
C21165 INVX1_LOC_162/Y INVX1_LOC_126/Y 0.42fF
C21166 NOR2X1_LOC_180/B NOR2X1_LOC_553/Y 0.16fF
C21167 INVX1_LOC_111/Y INVX1_LOC_75/A 0.04fF
C21168 NOR2X1_LOC_186/Y NAND2X1_LOC_286/a_36_24# 0.00fF
C21169 INVX1_LOC_237/Y INVX1_LOC_167/Y 0.19fF
C21170 NOR2X1_LOC_392/B INVX1_LOC_286/A 0.10fF
C21171 INVX1_LOC_191/Y NAND2X1_LOC_51/B 0.02fF
C21172 INVX1_LOC_53/A NAND2X1_LOC_74/B 0.03fF
C21173 NAND2X1_LOC_793/Y INVX1_LOC_118/A 0.01fF
C21174 NOR2X1_LOC_8/a_36_216# INVX1_LOC_59/Y 0.00fF
C21175 NOR2X1_LOC_721/A NOR2X1_LOC_721/Y 0.08fF
C21176 NOR2X1_LOC_554/B VDD 1.25fF
C21177 NOR2X1_LOC_92/Y INVX1_LOC_35/Y 0.07fF
C21178 NOR2X1_LOC_590/A NOR2X1_LOC_114/a_36_216# 0.00fF
C21179 INVX1_LOC_18/A INVX1_LOC_14/Y 0.31fF
C21180 NAND2X1_LOC_474/Y INVX1_LOC_285/A 0.17fF
C21181 INVX1_LOC_45/A NAND2X1_LOC_96/A 0.07fF
C21182 INVX1_LOC_62/A NOR2X1_LOC_99/B 0.04fF
C21183 INVX1_LOC_32/A NOR2X1_LOC_65/Y 0.00fF
C21184 INVX1_LOC_26/A NOR2X1_LOC_38/B 0.07fF
C21185 NAND2X1_LOC_594/a_36_24# NOR2X1_LOC_653/Y 0.00fF
C21186 NAND2X1_LOC_573/Y NAND2X1_LOC_286/a_36_24# 0.01fF
C21187 INVX1_LOC_300/Y INVX1_LOC_46/A 0.03fF
C21188 NOR2X1_LOC_616/Y NAND2X1_LOC_622/B 0.05fF
C21189 NOR2X1_LOC_273/Y INVX1_LOC_46/A 0.10fF
C21190 INPUT_2 NOR2X1_LOC_655/Y 0.15fF
C21191 INPUT_3 NOR2X1_LOC_656/Y 0.01fF
C21192 INVX1_LOC_35/A INVX1_LOC_284/A 0.07fF
C21193 INVX1_LOC_223/A NOR2X1_LOC_536/A 0.00fF
C21194 NAND2X1_LOC_850/Y NOR2X1_LOC_167/Y 0.01fF
C21195 NAND2X1_LOC_632/B NOR2X1_LOC_24/Y 0.32fF
C21196 NOR2X1_LOC_634/B NOR2X1_LOC_334/A 0.02fF
C21197 NOR2X1_LOC_264/Y NAND2X1_LOC_642/Y 0.03fF
C21198 NAND2X1_LOC_162/B INVX1_LOC_37/A 0.01fF
C21199 NOR2X1_LOC_78/B NOR2X1_LOC_334/A 0.35fF
C21200 INVX1_LOC_232/A NOR2X1_LOC_74/A 0.10fF
C21201 INVX1_LOC_58/A INVX1_LOC_15/A 0.13fF
C21202 NOR2X1_LOC_152/Y VDD 3.59fF
C21203 NOR2X1_LOC_188/A INVX1_LOC_16/A 0.00fF
C21204 NAND2X1_LOC_785/B INVX1_LOC_54/A 0.15fF
C21205 INVX1_LOC_300/Y NOR2X1_LOC_766/Y 0.05fF
C21206 NOR2X1_LOC_773/Y NOR2X1_LOC_183/a_36_216# -0.02fF
C21207 INVX1_LOC_113/Y VDD 0.98fF
C21208 NOR2X1_LOC_152/Y NAND2X1_LOC_800/A 0.06fF
C21209 INVX1_LOC_232/A NOR2X1_LOC_9/Y 0.10fF
C21210 NAND2X1_LOC_581/a_36_24# INVX1_LOC_15/A 0.00fF
C21211 NAND2X1_LOC_254/Y NOR2X1_LOC_291/a_36_216# 0.00fF
C21212 NAND2X1_LOC_350/A NOR2X1_LOC_841/A 0.10fF
C21213 NOR2X1_LOC_716/B INVX1_LOC_37/A 0.24fF
C21214 INVX1_LOC_10/A INVX1_LOC_67/Y 0.00fF
C21215 INVX1_LOC_286/Y NAND2X1_LOC_802/Y 0.07fF
C21216 NOR2X1_LOC_309/Y NOR2X1_LOC_279/Y 0.03fF
C21217 NOR2X1_LOC_554/B NOR2X1_LOC_846/a_36_216# 0.00fF
C21218 INVX1_LOC_223/A NAND2X1_LOC_93/B 0.68fF
C21219 INVX1_LOC_89/A NOR2X1_LOC_163/Y 0.12fF
C21220 NOR2X1_LOC_329/B INVX1_LOC_313/Y 0.02fF
C21221 NOR2X1_LOC_137/A INVX1_LOC_75/A 0.08fF
C21222 NOR2X1_LOC_383/Y NOR2X1_LOC_9/Y 0.02fF
C21223 NOR2X1_LOC_637/A INVX1_LOC_118/A 0.01fF
C21224 NOR2X1_LOC_441/Y NOR2X1_LOC_841/A 0.14fF
C21225 INPUT_2 INVX1_LOC_3/A 0.45fF
C21226 INVX1_LOC_136/A INVX1_LOC_92/A 0.17fF
C21227 INVX1_LOC_224/Y NAND2X1_LOC_99/A 0.07fF
C21228 NAND2X1_LOC_612/a_36_24# INVX1_LOC_3/A 0.00fF
C21229 NAND2X1_LOC_72/B INVX1_LOC_58/Y 0.11fF
C21230 INVX1_LOC_89/A NOR2X1_LOC_74/Y 0.01fF
C21231 INVX1_LOC_55/Y NOR2X1_LOC_742/A 0.07fF
C21232 INPUT_3 INVX1_LOC_63/A 0.15fF
C21233 NOR2X1_LOC_464/Y NOR2X1_LOC_678/A 0.01fF
C21234 NOR2X1_LOC_759/A INVX1_LOC_117/Y 0.01fF
C21235 NOR2X1_LOC_433/A INVX1_LOC_118/Y 0.08fF
C21236 INVX1_LOC_111/Y NOR2X1_LOC_309/a_36_216# 0.00fF
C21237 INVX1_LOC_44/Y INVX1_LOC_76/A 0.01fF
C21238 INVX1_LOC_5/A INVX1_LOC_4/Y 0.09fF
C21239 NAND2X1_LOC_850/Y INVX1_LOC_76/A 0.10fF
C21240 NOR2X1_LOC_721/A VDD 0.12fF
C21241 NOR2X1_LOC_570/B INVX1_LOC_38/A 0.02fF
C21242 NOR2X1_LOC_361/B INVX1_LOC_42/A 0.07fF
C21243 INVX1_LOC_271/A NOR2X1_LOC_125/Y 0.01fF
C21244 INVX1_LOC_28/A NOR2X1_LOC_188/A 0.05fF
C21245 NOR2X1_LOC_342/B NOR2X1_LOC_342/A 0.00fF
C21246 NOR2X1_LOC_307/B VDD 0.02fF
C21247 NOR2X1_LOC_172/Y INVX1_LOC_54/A 0.07fF
C21248 NAND2X1_LOC_768/a_36_24# NAND2X1_LOC_773/B 0.00fF
C21249 NOR2X1_LOC_16/Y INVX1_LOC_117/A 0.07fF
C21250 INVX1_LOC_90/A INVX1_LOC_286/A 0.07fF
C21251 INVX1_LOC_21/A NAND2X1_LOC_646/a_36_24# 0.00fF
C21252 NOR2X1_LOC_419/a_36_216# INVX1_LOC_46/Y 0.01fF
C21253 INVX1_LOC_249/A NOR2X1_LOC_155/A 0.02fF
C21254 NOR2X1_LOC_716/B NOR2X1_LOC_177/Y 0.04fF
C21255 NOR2X1_LOC_316/Y NOR2X1_LOC_536/A -0.01fF
C21256 INVX1_LOC_64/A NOR2X1_LOC_447/A 0.03fF
C21257 NOR2X1_LOC_510/Y INVX1_LOC_78/A 1.48fF
C21258 NOR2X1_LOC_389/B INVX1_LOC_286/A 0.01fF
C21259 INVX1_LOC_6/Y NOR2X1_LOC_155/A 0.01fF
C21260 NAND2X1_LOC_860/Y VDD 0.01fF
C21261 INVX1_LOC_49/A NAND2X1_LOC_798/B 0.07fF
C21262 NOR2X1_LOC_52/B INVX1_LOC_118/Y 0.04fF
C21263 NAND2X1_LOC_859/Y NOR2X1_LOC_670/Y 0.34fF
C21264 VDD NAND2X1_LOC_859/B 0.01fF
C21265 NOR2X1_LOC_392/B INVX1_LOC_54/A 0.10fF
C21266 NAND2X1_LOC_348/A INVX1_LOC_154/Y 0.09fF
C21267 NOR2X1_LOC_332/A INVX1_LOC_316/A -0.02fF
C21268 INVX1_LOC_58/A INVX1_LOC_278/A 0.08fF
C21269 INVX1_LOC_186/A NOR2X1_LOC_356/A 0.07fF
C21270 GATE_741 NOR2X1_LOC_829/A 0.42fF
C21271 INVX1_LOC_58/A NOR2X1_LOC_489/a_36_216# 0.02fF
C21272 INVX1_LOC_186/A NAND2X1_LOC_472/a_36_24# 0.01fF
C21273 INVX1_LOC_43/Y INVX1_LOC_127/Y 0.05fF
C21274 NAND2X1_LOC_715/B INVX1_LOC_271/A 0.00fF
C21275 INVX1_LOC_90/A INVX1_LOC_95/A 0.03fF
C21276 NOR2X1_LOC_470/A INVX1_LOC_37/A 0.18fF
C21277 NAND2X1_LOC_308/B INVX1_LOC_11/Y 0.01fF
C21278 INVX1_LOC_215/Y INVX1_LOC_15/A 0.07fF
C21279 NOR2X1_LOC_455/Y INVX1_LOC_64/A 0.00fF
C21280 INVX1_LOC_223/Y NOR2X1_LOC_383/B 0.00fF
C21281 NOR2X1_LOC_389/B INVX1_LOC_95/A 0.16fF
C21282 NOR2X1_LOC_361/B INVX1_LOC_78/A 0.04fF
C21283 NOR2X1_LOC_424/Y INVX1_LOC_37/A 0.14fF
C21284 NOR2X1_LOC_186/Y INVX1_LOC_57/A 0.23fF
C21285 NAND2X1_LOC_778/Y INVX1_LOC_50/A 0.09fF
C21286 NOR2X1_LOC_286/Y NOR2X1_LOC_334/Y 0.04fF
C21287 NOR2X1_LOC_644/A NOR2X1_LOC_486/Y 0.00fF
C21288 INVX1_LOC_1/Y INVX1_LOC_66/Y 0.02fF
C21289 NOR2X1_LOC_802/A NOR2X1_LOC_809/B 0.02fF
C21290 NAND2X1_LOC_850/A NAND2X1_LOC_642/Y 0.21fF
C21291 INVX1_LOC_311/A INVX1_LOC_6/A 0.49fF
C21292 INVX1_LOC_21/A INVX1_LOC_270/A 0.01fF
C21293 NOR2X1_LOC_411/A INVX1_LOC_64/A 0.18fF
C21294 NOR2X1_LOC_717/Y INVX1_LOC_283/A 0.01fF
C21295 NOR2X1_LOC_717/B INVX1_LOC_37/A 0.04fF
C21296 NOR2X1_LOC_203/a_36_216# INVX1_LOC_53/A 0.01fF
C21297 NOR2X1_LOC_468/Y INVX1_LOC_26/A 0.08fF
C21298 NOR2X1_LOC_356/A NAND2X1_LOC_447/Y 0.05fF
C21299 NAND2X1_LOC_214/B NOR2X1_LOC_598/B 0.01fF
C21300 NOR2X1_LOC_92/Y NAND2X1_LOC_286/B 0.03fF
C21301 NOR2X1_LOC_672/Y INVX1_LOC_203/A 0.11fF
C21302 NAND2X1_LOC_656/Y INVX1_LOC_12/Y 0.15fF
C21303 NAND2X1_LOC_315/a_36_24# INVX1_LOC_29/A 0.01fF
C21304 NAND2X1_LOC_861/Y VDD 0.62fF
C21305 NAND2X1_LOC_634/Y NAND2X1_LOC_254/Y 0.04fF
C21306 NOR2X1_LOC_68/A NOR2X1_LOC_67/Y 0.01fF
C21307 INVX1_LOC_27/A NOR2X1_LOC_125/Y 0.07fF
C21308 NAND2X1_LOC_116/A NOR2X1_LOC_243/B 0.07fF
C21309 INVX1_LOC_21/A NOR2X1_LOC_416/A 0.07fF
C21310 INVX1_LOC_215/A INVX1_LOC_38/A 0.07fF
C21311 NOR2X1_LOC_859/A NOR2X1_LOC_861/Y 0.03fF
C21312 NAND2X1_LOC_573/Y INVX1_LOC_57/A 0.01fF
C21313 NOR2X1_LOC_748/a_36_216# NOR2X1_LOC_641/Y 0.03fF
C21314 NOR2X1_LOC_226/A NAND2X1_LOC_798/B 0.19fF
C21315 D_INPUT_0 INVX1_LOC_33/Y 0.06fF
C21316 NOR2X1_LOC_65/B NOR2X1_LOC_361/B 0.25fF
C21317 INVX1_LOC_50/A NOR2X1_LOC_15/Y 3.58fF
C21318 NOR2X1_LOC_598/B INVX1_LOC_27/A 0.24fF
C21319 NOR2X1_LOC_828/A INVX1_LOC_37/A 0.01fF
C21320 INVX1_LOC_25/A INVX1_LOC_48/Y 0.02fF
C21321 NAND2X1_LOC_557/Y NAND2X1_LOC_579/A 0.03fF
C21322 NOR2X1_LOC_551/B INVX1_LOC_19/A 0.01fF
C21323 INVX1_LOC_77/A INVX1_LOC_69/A 0.05fF
C21324 NOR2X1_LOC_103/Y NAND2X1_LOC_99/A 2.91fF
C21325 NAND2X1_LOC_564/A NOR2X1_LOC_468/Y 0.01fF
C21326 INVX1_LOC_225/A NOR2X1_LOC_662/A 0.01fF
C21327 INVX1_LOC_156/A VDD 0.12fF
C21328 NAND2X1_LOC_860/A NOR2X1_LOC_92/Y 0.17fF
C21329 NOR2X1_LOC_74/A NAND2X1_LOC_447/Y 0.10fF
C21330 INVX1_LOC_21/A NOR2X1_LOC_109/Y 0.16fF
C21331 NAND2X1_LOC_740/B NOR2X1_LOC_305/Y 0.46fF
C21332 NOR2X1_LOC_824/A NAND2X1_LOC_725/A 0.10fF
C21333 NOR2X1_LOC_244/B NOR2X1_LOC_865/Y 0.05fF
C21334 NAND2X1_LOC_661/A VDD -0.00fF
C21335 INVX1_LOC_282/A INVX1_LOC_76/A 0.15fF
C21336 INVX1_LOC_304/A INVX1_LOC_6/A 0.07fF
C21337 NOR2X1_LOC_67/A NOR2X1_LOC_813/a_36_216# 0.00fF
C21338 NAND2X1_LOC_555/Y NAND2X1_LOC_416/a_36_24# 0.00fF
C21339 INVX1_LOC_208/Y NAND2X1_LOC_288/A 0.04fF
C21340 NOR2X1_LOC_188/A NOR2X1_LOC_35/Y 0.10fF
C21341 NOR2X1_LOC_9/Y NAND2X1_LOC_447/Y 0.01fF
C21342 INVX1_LOC_56/Y NOR2X1_LOC_179/a_36_216# 0.00fF
C21343 NAND2X1_LOC_725/A INVX1_LOC_237/A 0.18fF
C21344 NOR2X1_LOC_34/B NAND2X1_LOC_27/a_36_24# 0.02fF
C21345 NOR2X1_LOC_845/A NAND2X1_LOC_813/a_36_24# 0.02fF
C21346 NOR2X1_LOC_151/Y INVX1_LOC_37/A 0.07fF
C21347 INVX1_LOC_269/A NOR2X1_LOC_717/A 0.19fF
C21348 INVX1_LOC_201/Y NOR2X1_LOC_610/Y 0.06fF
C21349 INVX1_LOC_53/Y NAND2X1_LOC_572/B 0.07fF
C21350 INVX1_LOC_90/A NOR2X1_LOC_602/B 0.01fF
C21351 INVX1_LOC_153/Y INVX1_LOC_42/A 0.46fF
C21352 INVX1_LOC_10/A NOR2X1_LOC_364/A 0.14fF
C21353 VDD INVX1_LOC_158/Y 0.21fF
C21354 INVX1_LOC_8/A NAND2X1_LOC_254/Y 0.07fF
C21355 NOR2X1_LOC_763/Y NAND2X1_LOC_430/a_36_24# 0.01fF
C21356 INVX1_LOC_174/A INVX1_LOC_23/A 0.05fF
C21357 INVX1_LOC_83/A INVX1_LOC_75/Y 0.04fF
C21358 NOR2X1_LOC_274/Y INVX1_LOC_4/A 0.01fF
C21359 INVX1_LOC_45/A NAND2X1_LOC_99/A 0.08fF
C21360 INVX1_LOC_90/A INVX1_LOC_54/A 7.85fF
C21361 NOR2X1_LOC_791/A INVX1_LOC_23/Y -0.07fF
C21362 INVX1_LOC_5/A NOR2X1_LOC_205/Y 0.01fF
C21363 INVX1_LOC_89/A INVX1_LOC_179/A 0.03fF
C21364 NOR2X1_LOC_78/B NAND2X1_LOC_74/B 0.13fF
C21365 NAND2X1_LOC_30/Y NAND2X1_LOC_31/a_36_24# 0.00fF
C21366 NOR2X1_LOC_778/B INVX1_LOC_29/A 1.70fF
C21367 NOR2X1_LOC_152/a_36_216# INVX1_LOC_273/A 0.02fF
C21368 NOR2X1_LOC_773/Y NAND2X1_LOC_81/B 0.07fF
C21369 INVX1_LOC_62/Y INVX1_LOC_26/A 0.18fF
C21370 INVX1_LOC_177/A INVX1_LOC_42/A 0.03fF
C21371 INVX1_LOC_10/A INVX1_LOC_285/A 0.07fF
C21372 INVX1_LOC_208/Y INVX1_LOC_19/A 0.00fF
C21373 INVX1_LOC_24/A NAND2X1_LOC_61/Y 0.09fF
C21374 NOR2X1_LOC_91/Y NAND2X1_LOC_442/a_36_24# 0.00fF
C21375 INVX1_LOC_27/A NOR2X1_LOC_271/a_36_216# 0.01fF
C21376 NOR2X1_LOC_516/B NAND2X1_LOC_82/Y 0.01fF
C21377 NOR2X1_LOC_178/Y INVX1_LOC_43/Y 0.01fF
C21378 INVX1_LOC_48/Y INVX1_LOC_1/A 0.10fF
C21379 INVX1_LOC_280/Y INVX1_LOC_42/A 0.03fF
C21380 INVX1_LOC_286/A NOR2X1_LOC_561/A 0.02fF
C21381 INVX1_LOC_71/A NAND2X1_LOC_99/A 0.06fF
C21382 NOR2X1_LOC_458/Y INVX1_LOC_78/A 0.00fF
C21383 INVX1_LOC_153/Y INVX1_LOC_78/A 0.18fF
C21384 INVX1_LOC_136/A INVX1_LOC_53/A 0.11fF
C21385 INVX1_LOC_224/Y NAND2X1_LOC_656/A 0.11fF
C21386 NAND2X1_LOC_303/Y NOR2X1_LOC_536/Y 0.02fF
C21387 INVX1_LOC_2/A INVX1_LOC_47/Y 0.01fF
C21388 NAND2X1_LOC_764/a_36_24# INVX1_LOC_53/A 0.01fF
C21389 INVX1_LOC_290/A INVX1_LOC_261/Y 0.01fF
C21390 INVX1_LOC_35/A INVX1_LOC_72/A 0.10fF
C21391 NOR2X1_LOC_181/A INVX1_LOC_37/A 0.01fF
C21392 INVX1_LOC_49/A NAND2X1_LOC_211/a_36_24# 0.00fF
C21393 NAND2X1_LOC_392/Y NAND2X1_LOC_74/B 0.05fF
C21394 NOR2X1_LOC_226/A INVX1_LOC_47/Y 0.29fF
C21395 INVX1_LOC_77/A INVX1_LOC_270/Y 0.17fF
C21396 NOR2X1_LOC_457/B NOR2X1_LOC_678/A 0.01fF
C21397 NAND2X1_LOC_568/A NAND2X1_LOC_537/Y 0.02fF
C21398 NOR2X1_LOC_15/Y NAND2X1_LOC_227/Y 0.07fF
C21399 NOR2X1_LOC_357/Y INVX1_LOC_139/A 0.01fF
C21400 NAND2X1_LOC_660/a_36_24# INVX1_LOC_49/Y 0.00fF
C21401 NOR2X1_LOC_824/A NOR2X1_LOC_372/A 0.12fF
C21402 INVX1_LOC_132/A INVX1_LOC_57/A 0.07fF
C21403 INVX1_LOC_59/A INVX1_LOC_230/Y 0.14fF
C21404 INVX1_LOC_177/A INVX1_LOC_78/A 0.04fF
C21405 NAND2X1_LOC_799/a_36_24# INVX1_LOC_78/A 0.00fF
C21406 INVX1_LOC_83/A NAND2X1_LOC_207/Y 0.39fF
C21407 NOR2X1_LOC_481/A INVX1_LOC_57/A 0.00fF
C21408 INVX1_LOC_222/Y INVX1_LOC_45/A 0.93fF
C21409 INVX1_LOC_1/Y INVX1_LOC_32/A 0.03fF
C21410 INVX1_LOC_222/Y NOR2X1_LOC_568/A 0.01fF
C21411 INVX1_LOC_33/A NAND2X1_LOC_205/A 0.01fF
C21412 INVX1_LOC_21/A INVX1_LOC_36/A 13.40fF
C21413 NAND2X1_LOC_477/A NAND2X1_LOC_286/B 0.03fF
C21414 NOR2X1_LOC_454/Y NOR2X1_LOC_230/Y 0.06fF
C21415 INVX1_LOC_254/Y NAND2X1_LOC_363/B 0.00fF
C21416 INVX1_LOC_135/A NOR2X1_LOC_346/A 0.01fF
C21417 NOR2X1_LOC_561/a_36_216# INVX1_LOC_29/Y 0.00fF
C21418 INVX1_LOC_21/A NOR2X1_LOC_267/A 0.04fF
C21419 INVX1_LOC_225/A INVX1_LOC_57/A 3.56fF
C21420 NAND2X1_LOC_785/a_36_24# INVX1_LOC_41/Y 0.00fF
C21421 INVX1_LOC_41/A NAND2X1_LOC_860/A 0.07fF
C21422 NOR2X1_LOC_288/A INVX1_LOC_57/A 0.03fF
C21423 NAND2X1_LOC_162/A INVX1_LOC_78/A 0.01fF
C21424 INVX1_LOC_263/A NAND2X1_LOC_454/Y 0.04fF
C21425 INVX1_LOC_90/A NAND2X1_LOC_807/B 0.02fF
C21426 NAND2X1_LOC_571/B INVX1_LOC_34/A 0.01fF
C21427 INVX1_LOC_239/A INVX1_LOC_195/A 0.01fF
C21428 NAND2X1_LOC_714/a_36_24# INVX1_LOC_141/Y 0.00fF
C21429 INVX1_LOC_48/Y NOR2X1_LOC_384/Y 0.23fF
C21430 INVX1_LOC_64/A INVX1_LOC_237/Y 0.13fF
C21431 NAND2X1_LOC_53/Y NOR2X1_LOC_590/A 0.08fF
C21432 INVX1_LOC_124/A INVX1_LOC_270/Y 0.05fF
C21433 NOR2X1_LOC_389/B NAND2X1_LOC_807/B 0.22fF
C21434 INVX1_LOC_50/A INVX1_LOC_96/Y 0.69fF
C21435 INVX1_LOC_40/A INVX1_LOC_16/Y 1.49fF
C21436 NOR2X1_LOC_647/B NAND2X1_LOC_612/a_36_24# 0.02fF
C21437 INVX1_LOC_90/A NOR2X1_LOC_48/B 0.14fF
C21438 INVX1_LOC_25/A NOR2X1_LOC_84/Y 0.01fF
C21439 INVX1_LOC_21/A NOR2X1_LOC_208/Y 0.08fF
C21440 NAND2X1_LOC_860/A NAND2X1_LOC_477/A 0.10fF
C21441 NOR2X1_LOC_510/Y NOR2X1_LOC_152/Y 0.10fF
C21442 NAND2X1_LOC_725/Y NAND2X1_LOC_717/Y 0.17fF
C21443 INVX1_LOC_40/A NOR2X1_LOC_39/Y 0.07fF
C21444 NAND2X1_LOC_728/Y NAND2X1_LOC_303/Y 0.10fF
C21445 INVX1_LOC_80/Y NOR2X1_LOC_660/Y 0.02fF
C21446 INVX1_LOC_233/Y NAND2X1_LOC_562/B 0.01fF
C21447 INVX1_LOC_33/Y NAND2X1_LOC_848/A 0.01fF
C21448 INVX1_LOC_21/A NOR2X1_LOC_237/Y 2.14fF
C21449 NOR2X1_LOC_332/A INVX1_LOC_4/Y 0.03fF
C21450 NOR2X1_LOC_182/a_36_216# NOR2X1_LOC_678/A 0.00fF
C21451 INVX1_LOC_256/A INVX1_LOC_223/A 0.10fF
C21452 INPUT_1 INVX1_LOC_47/Y 0.01fF
C21453 NOR2X1_LOC_528/a_36_216# INVX1_LOC_78/A 0.00fF
C21454 NOR2X1_LOC_852/B NOR2X1_LOC_852/Y -0.01fF
C21455 D_INPUT_1 NAND2X1_LOC_181/Y 0.03fF
C21456 INVX1_LOC_135/A INVX1_LOC_94/Y 0.10fF
C21457 NAND2X1_LOC_633/Y NOR2X1_LOC_177/Y 0.06fF
C21458 NOR2X1_LOC_91/A NOR2X1_LOC_589/A 0.07fF
C21459 VDD INVX1_LOC_291/A 0.00fF
C21460 NAND2X1_LOC_218/B INVX1_LOC_14/A 0.12fF
C21461 INVX1_LOC_35/A NOR2X1_LOC_537/Y 0.00fF
C21462 INVX1_LOC_35/A NAND2X1_LOC_338/B 0.22fF
C21463 VDD NAND2X1_LOC_802/Y 0.38fF
C21464 NAND2X1_LOC_800/A INVX1_LOC_291/A 0.12fF
C21465 NAND2X1_LOC_89/a_36_24# NOR2X1_LOC_160/B 0.00fF
C21466 NOR2X1_LOC_91/A INVX1_LOC_229/Y 0.41fF
C21467 INVX1_LOC_305/A NAND2X1_LOC_171/a_36_24# 0.01fF
C21468 NOR2X1_LOC_742/A INVX1_LOC_32/A 0.07fF
C21469 NOR2X1_LOC_802/A INVX1_LOC_50/Y 0.09fF
C21470 INVX1_LOC_21/A NOR2X1_LOC_309/Y 0.14fF
C21471 INVX1_LOC_35/A NAND2X1_LOC_323/B 0.00fF
C21472 D_INPUT_0 INVX1_LOC_23/Y 0.08fF
C21473 NOR2X1_LOC_130/A NAND2X1_LOC_61/Y 0.03fF
C21474 NOR2X1_LOC_15/Y NOR2X1_LOC_679/B 0.07fF
C21475 INVX1_LOC_196/Y INVX1_LOC_271/Y -0.00fF
C21476 NOR2X1_LOC_319/B NOR2X1_LOC_856/A 0.11fF
C21477 NOR2X1_LOC_667/A NOR2X1_LOC_109/Y 0.14fF
C21478 INVX1_LOC_91/A INVX1_LOC_272/A 0.07fF
C21479 NOR2X1_LOC_589/A INVX1_LOC_23/A 0.24fF
C21480 INVX1_LOC_38/A INVX1_LOC_54/A 0.53fF
C21481 INVX1_LOC_248/A NOR2X1_LOC_109/Y 0.18fF
C21482 NOR2X1_LOC_459/B INVX1_LOC_163/A 0.06fF
C21483 NOR2X1_LOC_860/Y INVX1_LOC_230/A 0.03fF
C21484 NOR2X1_LOC_206/a_36_216# INVX1_LOC_96/Y 0.00fF
C21485 INVX1_LOC_27/A NOR2X1_LOC_156/B 0.02fF
C21486 INVX1_LOC_13/Y NAND2X1_LOC_374/Y 0.32fF
C21487 INVX1_LOC_223/Y NOR2X1_LOC_168/A 0.05fF
C21488 NOR2X1_LOC_363/Y NAND2X1_LOC_792/a_36_24# 0.00fF
C21489 NAND2X1_LOC_552/A NAND2X1_LOC_862/A 0.28fF
C21490 INVX1_LOC_36/A NAND2X1_LOC_354/Y 0.00fF
C21491 INVX1_LOC_6/A INVX1_LOC_19/Y 0.05fF
C21492 INVX1_LOC_272/Y NAND2X1_LOC_354/B 0.07fF
C21493 NOR2X1_LOC_3/a_36_216# INVX1_LOC_30/A 0.01fF
C21494 NOR2X1_LOC_445/Y NOR2X1_LOC_457/A 0.05fF
C21495 NOR2X1_LOC_51/A INVX1_LOC_54/A 0.25fF
C21496 NAND2X1_LOC_350/A NOR2X1_LOC_172/Y 0.00fF
C21497 INVX1_LOC_1/A NOR2X1_LOC_84/Y 0.10fF
C21498 INVX1_LOC_293/Y INVX1_LOC_46/A 0.06fF
C21499 NOR2X1_LOC_368/Y NAND2X1_LOC_74/B 0.01fF
C21500 INVX1_LOC_123/A INVX1_LOC_3/Y 0.19fF
C21501 NOR2X1_LOC_841/A NAND2X1_LOC_61/a_36_24# 0.06fF
C21502 NAND2X1_LOC_483/Y NAND2X1_LOC_550/A 0.03fF
C21503 NOR2X1_LOC_219/B NOR2X1_LOC_160/B 0.01fF
C21504 NAND2X1_LOC_798/B INVX1_LOC_118/A 0.14fF
C21505 INVX1_LOC_256/A INVX1_LOC_149/Y 0.03fF
C21506 NAND2X1_LOC_721/A NAND2X1_LOC_489/Y 0.41fF
C21507 NOR2X1_LOC_644/A NOR2X1_LOC_748/A 0.03fF
C21508 INVX1_LOC_1/A INVX1_LOC_216/A 0.02fF
C21509 NAND2X1_LOC_131/a_36_24# NOR2X1_LOC_84/Y 0.01fF
C21510 NOR2X1_LOC_318/B INVX1_LOC_32/A 0.03fF
C21511 NOR2X1_LOC_441/Y NOR2X1_LOC_172/Y 0.02fF
C21512 INVX1_LOC_314/Y NOR2X1_LOC_82/a_36_216# 0.00fF
C21513 NOR2X1_LOC_33/A NOR2X1_LOC_249/Y 0.01fF
C21514 NOR2X1_LOC_439/B NOR2X1_LOC_383/B 0.02fF
C21515 INVX1_LOC_46/A NAND2X1_LOC_74/B 1.24fF
C21516 INVX1_LOC_64/A NAND2X1_LOC_45/Y 0.01fF
C21517 INVX1_LOC_57/Y NOR2X1_LOC_373/a_36_216# 0.00fF
C21518 NOR2X1_LOC_92/Y INVX1_LOC_172/Y 0.03fF
C21519 NOR2X1_LOC_376/A INVX1_LOC_22/A 0.00fF
C21520 NOR2X1_LOC_98/A NAND2X1_LOC_74/B -0.03fF
C21521 INVX1_LOC_93/Y INVX1_LOC_32/A 0.10fF
C21522 NOR2X1_LOC_180/B NOR2X1_LOC_678/A 0.01fF
C21523 NOR2X1_LOC_454/a_36_216# INVX1_LOC_72/A 0.00fF
C21524 INVX1_LOC_75/A NOR2X1_LOC_383/B 0.11fF
C21525 INVX1_LOC_11/A NOR2X1_LOC_520/A 0.01fF
C21526 NAND2X1_LOC_799/a_36_24# NOR2X1_LOC_503/Y 0.00fF
C21527 NOR2X1_LOC_359/Y NOR2X1_LOC_363/a_36_216# 0.00fF
C21528 INVX1_LOC_2/A NOR2X1_LOC_679/Y 0.05fF
C21529 D_INPUT_6 INPUT_5 0.10fF
C21530 NAND2X1_LOC_348/A NAND2X1_LOC_215/A 0.00fF
C21531 NOR2X1_LOC_160/B NOR2X1_LOC_168/B 0.04fF
C21532 NOR2X1_LOC_412/a_36_216# NOR2X1_LOC_384/Y 0.01fF
C21533 INVX1_LOC_94/A NOR2X1_LOC_303/Y 0.10fF
C21534 INVX1_LOC_64/A NOR2X1_LOC_330/a_36_216# 0.02fF
C21535 INVX1_LOC_14/A INVX1_LOC_22/A 0.22fF
C21536 NOR2X1_LOC_817/Y INVX1_LOC_40/A 0.01fF
C21537 INVX1_LOC_1/A INVX1_LOC_290/A 0.17fF
C21538 INVX1_LOC_58/A NOR2X1_LOC_310/a_36_216# 0.10fF
C21539 NOR2X1_LOC_690/A INVX1_LOC_18/A 0.10fF
C21540 NOR2X1_LOC_716/B NAND2X1_LOC_198/B 0.24fF
C21541 NOR2X1_LOC_299/Y INVX1_LOC_242/A 0.03fF
C21542 NAND2X1_LOC_739/B NOR2X1_LOC_577/Y 0.06fF
C21543 INVX1_LOC_100/Y INVX1_LOC_26/A 0.01fF
C21544 INVX1_LOC_300/Y NAND2X1_LOC_812/A 0.05fF
C21545 NOR2X1_LOC_78/B NOR2X1_LOC_276/Y 0.03fF
C21546 NAND2X1_LOC_338/B NAND2X1_LOC_527/a_36_24# 0.01fF
C21547 INVX1_LOC_73/A NOR2X1_LOC_678/A 0.00fF
C21548 NAND2X1_LOC_182/a_36_24# NAND2X1_LOC_793/Y 0.01fF
C21549 INVX1_LOC_24/A NOR2X1_LOC_520/B 0.09fF
C21550 INVX1_LOC_11/A NOR2X1_LOC_748/Y 0.00fF
C21551 NOR2X1_LOC_194/Y INVX1_LOC_18/A 0.01fF
C21552 INVX1_LOC_24/A NAND2X1_LOC_325/Y 0.07fF
C21553 NOR2X1_LOC_68/A INVX1_LOC_104/A 0.10fF
C21554 INVX1_LOC_13/A NOR2X1_LOC_82/A 0.13fF
C21555 NOR2X1_LOC_690/A NAND2X1_LOC_711/B 0.39fF
C21556 VDD NOR2X1_LOC_609/Y 0.18fF
C21557 NOR2X1_LOC_590/A NOR2X1_LOC_500/Y 0.45fF
C21558 NOR2X1_LOC_445/B NOR2X1_LOC_814/A 0.01fF
C21559 INVX1_LOC_299/A INVX1_LOC_135/A 0.03fF
C21560 INVX1_LOC_36/A INVX1_LOC_214/A 0.03fF
C21561 NOR2X1_LOC_346/A INVX1_LOC_280/A 0.05fF
C21562 INVX1_LOC_226/Y NOR2X1_LOC_590/A 0.03fF
C21563 NAND2X1_LOC_860/A NOR2X1_LOC_71/a_36_216# 0.01fF
C21564 INVX1_LOC_36/A NOR2X1_LOC_667/A 0.18fF
C21565 INVX1_LOC_314/Y INVX1_LOC_8/A 0.10fF
C21566 INVX1_LOC_34/A NOR2X1_LOC_495/Y 0.02fF
C21567 NOR2X1_LOC_197/Y INVX1_LOC_50/Y 0.02fF
C21568 INVX1_LOC_36/A INVX1_LOC_248/A 0.98fF
C21569 NOR2X1_LOC_690/A INVX1_LOC_172/A 0.07fF
C21570 NOR2X1_LOC_712/Y NOR2X1_LOC_712/B 0.01fF
C21571 NOR2X1_LOC_48/B INVX1_LOC_38/A 0.63fF
C21572 NAND2X1_LOC_9/Y NOR2X1_LOC_334/A 0.01fF
C21573 INVX1_LOC_153/Y INVX1_LOC_113/Y 0.01fF
C21574 INVX1_LOC_136/A NOR2X1_LOC_78/B 0.16fF
C21575 NAND2X1_LOC_803/B INVX1_LOC_10/A 0.02fF
C21576 INVX1_LOC_247/Y NOR2X1_LOC_778/B 0.01fF
C21577 NOR2X1_LOC_418/a_36_216# INVX1_LOC_72/A 0.00fF
C21578 NOR2X1_LOC_824/A NAND2X1_LOC_560/A 0.01fF
C21579 NOR2X1_LOC_717/Y INVX1_LOC_22/A 0.03fF
C21580 INVX1_LOC_57/A NAND2X1_LOC_642/Y 0.11fF
C21581 INVX1_LOC_83/A NOR2X1_LOC_307/A 1.25fF
C21582 NAND2X1_LOC_326/A INVX1_LOC_28/A 0.29fF
C21583 NOR2X1_LOC_310/Y INVX1_LOC_77/A 0.02fF
C21584 INVX1_LOC_57/Y INVX1_LOC_25/Y 0.14fF
C21585 INVX1_LOC_224/A INVX1_LOC_65/Y 0.00fF
C21586 NOR2X1_LOC_294/Y NOR2X1_LOC_516/B 0.03fF
C21587 INVX1_LOC_121/Y INVX1_LOC_113/Y 0.16fF
C21588 INVX1_LOC_276/A INVX1_LOC_24/A 0.03fF
C21589 NOR2X1_LOC_89/A INVX1_LOC_70/A 0.10fF
C21590 NOR2X1_LOC_160/B NAND2X1_LOC_656/Y 0.07fF
C21591 NOR2X1_LOC_364/A INVX1_LOC_12/A 0.01fF
C21592 INVX1_LOC_293/A INVX1_LOC_135/A 0.01fF
C21593 NOR2X1_LOC_590/A INVX1_LOC_10/A 0.11fF
C21594 NOR2X1_LOC_91/A INVX1_LOC_20/A 1.20fF
C21595 NAND2X1_LOC_244/A NOR2X1_LOC_693/Y 0.00fF
C21596 NOR2X1_LOC_67/A INVX1_LOC_24/A 0.18fF
C21597 NOR2X1_LOC_540/B NOR2X1_LOC_748/A 0.01fF
C21598 INVX1_LOC_216/Y INPUT_1 0.01fF
C21599 INVX1_LOC_11/A D_GATE_366 0.07fF
C21600 INVX1_LOC_290/Y NAND2X1_LOC_93/B 0.07fF
C21601 INVX1_LOC_201/Y NOR2X1_LOC_516/Y 0.05fF
C21602 NAND2X1_LOC_149/Y NOR2X1_LOC_74/a_36_216# 0.01fF
C21603 NOR2X1_LOC_392/B NOR2X1_LOC_142/Y 0.33fF
C21604 INVX1_LOC_45/A INVX1_LOC_220/Y 0.12fF
C21605 NOR2X1_LOC_152/A INVX1_LOC_94/Y 0.05fF
C21606 INVX1_LOC_34/A INVX1_LOC_219/Y 0.04fF
C21607 NOR2X1_LOC_679/Y NAND2X1_LOC_648/A 0.03fF
C21608 INVX1_LOC_182/Y NOR2X1_LOC_359/a_36_216# 0.00fF
C21609 NOR2X1_LOC_222/Y INVX1_LOC_71/A 0.03fF
C21610 INVX1_LOC_147/Y INVX1_LOC_23/A 0.06fF
C21611 INVX1_LOC_111/Y NOR2X1_LOC_577/Y 0.01fF
C21612 NAND2X1_LOC_350/A INVX1_LOC_90/A 0.84fF
C21613 NOR2X1_LOC_626/Y INVX1_LOC_6/A 0.00fF
C21614 NOR2X1_LOC_691/A INVX1_LOC_19/A 0.01fF
C21615 NOR2X1_LOC_798/A NOR2X1_LOC_334/A 0.02fF
C21616 GATE_811 NAND2X1_LOC_812/a_36_24# 0.02fF
C21617 NOR2X1_LOC_360/Y NOR2X1_LOC_188/a_36_216# 0.12fF
C21618 NAND2X1_LOC_739/B INVX1_LOC_22/A 0.03fF
C21619 INVX1_LOC_98/A INVX1_LOC_306/Y 0.10fF
C21620 INVX1_LOC_12/A INVX1_LOC_285/A 0.72fF
C21621 INVX1_LOC_27/A INVX1_LOC_201/A 0.01fF
C21622 NAND2X1_LOC_574/A NOR2X1_LOC_610/Y 0.03fF
C21623 INVX1_LOC_23/A INVX1_LOC_20/A 0.29fF
C21624 INVX1_LOC_90/A INVX1_LOC_218/Y 0.03fF
C21625 INVX1_LOC_314/Y NOR2X1_LOC_315/a_36_216# 0.00fF
C21626 NOR2X1_LOC_468/Y NOR2X1_LOC_368/A 0.02fF
C21627 NOR2X1_LOC_91/A NOR2X1_LOC_765/Y 0.03fF
C21628 NOR2X1_LOC_401/a_36_216# NOR2X1_LOC_716/B 0.01fF
C21629 NOR2X1_LOC_78/A INVX1_LOC_306/Y 0.03fF
C21630 INVX1_LOC_32/A INVX1_LOC_117/Y 0.00fF
C21631 NAND2X1_LOC_84/Y INVX1_LOC_22/A 0.15fF
C21632 NAND2X1_LOC_558/a_36_24# INVX1_LOC_282/A 0.00fF
C21633 INVX1_LOC_90/A NOR2X1_LOC_441/Y 0.03fF
C21634 NOR2X1_LOC_641/B INVX1_LOC_89/A 0.08fF
C21635 INVX1_LOC_12/A NOR2X1_LOC_814/A 0.03fF
C21636 NAND2X1_LOC_848/A INVX1_LOC_23/Y 0.03fF
C21637 NOR2X1_LOC_658/Y NOR2X1_LOC_214/B 0.01fF
C21638 INVX1_LOC_269/A NOR2X1_LOC_337/A 0.03fF
C21639 INVX1_LOC_292/A NOR2X1_LOC_564/Y 0.01fF
C21640 NOR2X1_LOC_619/A NOR2X1_LOC_419/Y 0.02fF
C21641 INVX1_LOC_77/Y NOR2X1_LOC_654/A 0.02fF
C21642 NOR2X1_LOC_751/Y INVX1_LOC_89/A 0.03fF
C21643 NOR2X1_LOC_821/Y NOR2X1_LOC_822/Y 0.01fF
C21644 NOR2X1_LOC_716/B INVX1_LOC_53/Y 0.07fF
C21645 NOR2X1_LOC_667/A NOR2X1_LOC_309/Y 0.07fF
C21646 NOR2X1_LOC_457/A NOR2X1_LOC_335/B 0.13fF
C21647 D_INPUT_1 INVX1_LOC_117/A 0.03fF
C21648 INVX1_LOC_311/Y INVX1_LOC_30/A 0.03fF
C21649 INVX1_LOC_208/A INVX1_LOC_88/Y 0.44fF
C21650 INVX1_LOC_45/A NOR2X1_LOC_329/B 0.06fF
C21651 INVX1_LOC_91/A INVX1_LOC_198/A 0.01fF
C21652 NOR2X1_LOC_6/B NAND2X1_LOC_672/B 0.04fF
C21653 NOR2X1_LOC_121/Y INVX1_LOC_232/A 0.03fF
C21654 INVX1_LOC_215/A INVX1_LOC_33/A 0.07fF
C21655 NOR2X1_LOC_671/Y NAND2X1_LOC_74/B 0.00fF
C21656 INVX1_LOC_1/A INVX1_LOC_160/A 0.14fF
C21657 INVX1_LOC_171/A INVX1_LOC_111/A 0.01fF
C21658 INVX1_LOC_91/A NOR2X1_LOC_271/B 0.12fF
C21659 INVX1_LOC_57/A NOR2X1_LOC_271/Y 0.09fF
C21660 NAND2X1_LOC_475/Y INVX1_LOC_15/A 0.03fF
C21661 INVX1_LOC_45/A D_INPUT_4 0.01fF
C21662 NOR2X1_LOC_220/A INVX1_LOC_149/A 0.40fF
C21663 INVX1_LOC_270/Y INVX1_LOC_9/A 0.05fF
C21664 INVX1_LOC_180/A NOR2X1_LOC_130/A 0.02fF
C21665 NOR2X1_LOC_690/A NOR2X1_LOC_690/Y 0.28fF
C21666 INVX1_LOC_150/Y NOR2X1_LOC_114/A 0.02fF
C21667 NAND2X1_LOC_229/a_36_24# INVX1_LOC_143/A 0.01fF
C21668 INVX1_LOC_104/A NOR2X1_LOC_570/Y 0.03fF
C21669 INVX1_LOC_31/A INVX1_LOC_222/A 0.15fF
C21670 INVX1_LOC_23/Y INVX1_LOC_46/Y 0.14fF
C21671 INVX1_LOC_17/A NOR2X1_LOC_45/B 2.24fF
C21672 NAND2X1_LOC_92/a_36_24# NAND2X1_LOC_99/A 0.00fF
C21673 NOR2X1_LOC_89/A INVX1_LOC_102/A 0.07fF
C21674 NOR2X1_LOC_137/A NOR2X1_LOC_577/Y 0.01fF
C21675 NOR2X1_LOC_612/B INVX1_LOC_22/A 0.04fF
C21676 NOR2X1_LOC_516/B NOR2X1_LOC_168/B 0.03fF
C21677 NOR2X1_LOC_418/Y INVX1_LOC_191/Y 0.24fF
C21678 INVX1_LOC_2/A NOR2X1_LOC_328/Y 0.03fF
C21679 NOR2X1_LOC_246/A NAND2X1_LOC_316/a_36_24# 0.01fF
C21680 INVX1_LOC_150/Y INVX1_LOC_91/A 0.24fF
C21681 NOR2X1_LOC_278/A NAND2X1_LOC_392/Y 0.01fF
C21682 INVX1_LOC_47/Y NAND2X1_LOC_63/Y 0.23fF
C21683 NOR2X1_LOC_329/B INVX1_LOC_71/A 0.03fF
C21684 NOR2X1_LOC_599/A NOR2X1_LOC_387/A 0.03fF
C21685 NOR2X1_LOC_328/Y NOR2X1_LOC_226/A 0.05fF
C21686 NOR2X1_LOC_67/A NAND2X1_LOC_565/B 0.01fF
C21687 NOR2X1_LOC_392/B NOR2X1_LOC_99/B 0.00fF
C21688 NOR2X1_LOC_17/a_36_216# D_INPUT_5 0.00fF
C21689 INVX1_LOC_223/A INVX1_LOC_69/Y 0.01fF
C21690 NOR2X1_LOC_706/A NOR2X1_LOC_546/B 0.02fF
C21691 D_INPUT_0 NAND2X1_LOC_116/A 0.17fF
C21692 INVX1_LOC_41/A INVX1_LOC_85/Y 0.01fF
C21693 NOR2X1_LOC_238/Y NOR2X1_LOC_322/Y 0.01fF
C21694 INVX1_LOC_135/A NOR2X1_LOC_315/Y 0.01fF
C21695 NAND2X1_LOC_574/A NOR2X1_LOC_35/a_36_216# 0.01fF
C21696 INVX1_LOC_271/A NOR2X1_LOC_58/Y 0.01fF
C21697 INVX1_LOC_256/A INVX1_LOC_314/A 0.03fF
C21698 INVX1_LOC_114/Y NOR2X1_LOC_467/A 0.03fF
C21699 NOR2X1_LOC_289/Y NOR2X1_LOC_433/A 0.09fF
C21700 NOR2X1_LOC_757/Y NOR2X1_LOC_665/A 0.00fF
C21701 INVX1_LOC_296/Y INVX1_LOC_297/A 0.01fF
C21702 INVX1_LOC_276/A NAND2X1_LOC_783/A 0.15fF
C21703 NOR2X1_LOC_294/Y INVX1_LOC_315/Y 0.07fF
C21704 NOR2X1_LOC_471/Y INVX1_LOC_199/Y 0.04fF
C21705 NOR2X1_LOC_471/Y INVX1_LOC_247/A 0.01fF
C21706 INVX1_LOC_310/A INVX1_LOC_135/A 0.16fF
C21707 NAND2X1_LOC_395/a_36_24# INVX1_LOC_164/A 0.01fF
C21708 NAND2X1_LOC_787/A NOR2X1_LOC_88/Y 0.03fF
C21709 NOR2X1_LOC_657/Y NOR2X1_LOC_78/A 0.03fF
C21710 NOR2X1_LOC_590/A NOR2X1_LOC_799/B 0.01fF
C21711 NOR2X1_LOC_52/B D_GATE_366 0.01fF
C21712 NOR2X1_LOC_1/Y NOR2X1_LOC_30/Y 0.18fF
C21713 NOR2X1_LOC_706/A INVX1_LOC_275/A 0.67fF
C21714 NOR2X1_LOC_103/Y NAND2X1_LOC_611/a_36_24# 0.00fF
C21715 NOR2X1_LOC_67/A NOR2X1_LOC_130/A 0.07fF
C21716 INVX1_LOC_4/Y INVX1_LOC_42/A 0.17fF
C21717 INVX1_LOC_227/A NOR2X1_LOC_500/Y 0.08fF
C21718 NOR2X1_LOC_669/A NAND2X1_LOC_175/Y 0.05fF
C21719 INVX1_LOC_208/A NAND2X1_LOC_656/Y 0.07fF
C21720 NAND2X1_LOC_348/A NOR2X1_LOC_340/Y 0.04fF
C21721 INVX1_LOC_83/A NAND2X1_LOC_304/a_36_24# 0.00fF
C21722 INVX1_LOC_36/A INVX1_LOC_304/A 0.01fF
C21723 NAND2X1_LOC_361/Y INPUT_0 0.08fF
C21724 NAND2X1_LOC_35/Y INVX1_LOC_35/Y 0.01fF
C21725 INVX1_LOC_31/A INVX1_LOC_20/A 0.26fF
C21726 NOR2X1_LOC_655/B INVX1_LOC_90/A 0.03fF
C21727 INVX1_LOC_243/Y NOR2X1_LOC_48/Y 0.01fF
C21728 NOR2X1_LOC_464/B NOR2X1_LOC_331/B 0.01fF
C21729 NOR2X1_LOC_510/Y INVX1_LOC_291/A 0.02fF
C21730 INVX1_LOC_82/Y NOR2X1_LOC_6/B 0.06fF
C21731 NOR2X1_LOC_241/A INVX1_LOC_117/A 0.01fF
C21732 NAND2X1_LOC_787/A INVX1_LOC_84/A 0.04fF
C21733 NOR2X1_LOC_655/B NOR2X1_LOC_389/B 0.10fF
C21734 INVX1_LOC_50/A INVX1_LOC_49/Y 0.01fF
C21735 D_INPUT_0 INVX1_LOC_232/A 0.01fF
C21736 INVX1_LOC_279/Y VDD 0.41fF
C21737 INVX1_LOC_134/A NOR2X1_LOC_319/B 0.02fF
C21738 NOR2X1_LOC_584/Y NOR2X1_LOC_639/Y 0.02fF
C21739 NAND2X1_LOC_192/B NOR2X1_LOC_331/B 0.02fF
C21740 NAND2X1_LOC_9/Y INVX1_LOC_293/Y 0.04fF
C21741 INVX1_LOC_13/A INVX1_LOC_306/A 0.03fF
C21742 INVX1_LOC_33/A INVX1_LOC_286/A 0.07fF
C21743 NAND2X1_LOC_463/B NOR2X1_LOC_399/A 0.01fF
C21744 INVX1_LOC_271/A INVX1_LOC_29/A 1.72fF
C21745 INVX1_LOC_32/A INVX1_LOC_87/A 0.03fF
C21746 NOR2X1_LOC_763/Y NAND2X1_LOC_663/a_36_24# 0.06fF
C21747 NOR2X1_LOC_454/Y NAND2X1_LOC_93/B 0.01fF
C21748 INVX1_LOC_227/A INVX1_LOC_10/A 0.14fF
C21749 NAND2X1_LOC_556/a_36_24# INVX1_LOC_282/A 0.00fF
C21750 INVX1_LOC_142/A INVX1_LOC_76/A 0.94fF
C21751 INVX1_LOC_255/Y INVX1_LOC_89/A 0.21fF
C21752 INVX1_LOC_69/Y INVX1_LOC_149/Y 0.02fF
C21753 NOR2X1_LOC_589/A INVX1_LOC_313/A 0.03fF
C21754 NAND2X1_LOC_513/B NOR2X1_LOC_155/A 0.01fF
C21755 NOR2X1_LOC_168/A INVX1_LOC_75/A 0.01fF
C21756 NAND2X1_LOC_350/A INVX1_LOC_38/A 0.04fF
C21757 INVX1_LOC_32/A INVX1_LOC_175/A 0.03fF
C21758 INVX1_LOC_293/A INVX1_LOC_280/A 0.29fF
C21759 NOR2X1_LOC_655/B NAND2X1_LOC_348/A 0.01fF
C21760 NOR2X1_LOC_454/Y NAND2X1_LOC_425/Y 0.01fF
C21761 INVX1_LOC_136/A INVX1_LOC_46/A 2.88fF
C21762 NOR2X1_LOC_500/Y NOR2X1_LOC_703/A 0.02fF
C21763 INVX1_LOC_140/A NAND2X1_LOC_862/A 0.01fF
C21764 INVX1_LOC_78/A INVX1_LOC_4/Y 0.14fF
C21765 NAND2X1_LOC_9/Y NAND2X1_LOC_74/B 0.08fF
C21766 INVX1_LOC_34/A INVX1_LOC_159/Y 0.01fF
C21767 NOR2X1_LOC_557/A INVX1_LOC_8/A 0.02fF
C21768 INVX1_LOC_233/A NAND2X1_LOC_74/B 0.07fF
C21769 NOR2X1_LOC_770/B INVX1_LOC_91/A 0.00fF
C21770 NOR2X1_LOC_441/Y INVX1_LOC_38/A 0.06fF
C21771 NOR2X1_LOC_617/a_36_216# INVX1_LOC_20/A -0.00fF
C21772 INVX1_LOC_229/Y NAND2X1_LOC_866/B 0.10fF
C21773 INVX1_LOC_279/A INVX1_LOC_196/Y 0.22fF
C21774 NOR2X1_LOC_140/A NAND2X1_LOC_141/Y 0.01fF
C21775 INVX1_LOC_27/A NOR2X1_LOC_673/B 0.04fF
C21776 NAND2X1_LOC_860/A INVX1_LOC_168/Y 0.04fF
C21777 NAND2X1_LOC_569/a_36_24# NOR2X1_LOC_536/A 0.00fF
C21778 NOR2X1_LOC_34/A NOR2X1_LOC_814/A 0.04fF
C21779 INVX1_LOC_21/A INVX1_LOC_63/A 0.38fF
C21780 INVX1_LOC_135/A NAND2X1_LOC_624/A 0.03fF
C21781 NOR2X1_LOC_188/A NAND2X1_LOC_292/a_36_24# 0.00fF
C21782 INVX1_LOC_90/A NOR2X1_LOC_99/B 0.07fF
C21783 NAND2X1_LOC_593/Y INVX1_LOC_76/A 0.10fF
C21784 NOR2X1_LOC_179/Y NOR2X1_LOC_271/B 0.34fF
C21785 NAND2X1_LOC_35/Y NOR2X1_LOC_824/a_36_216# 0.01fF
C21786 NOR2X1_LOC_570/B NOR2X1_LOC_486/Y 0.10fF
C21787 NOR2X1_LOC_65/B INVX1_LOC_4/Y 0.10fF
C21788 D_INPUT_1 INVX1_LOC_3/Y 0.11fF
C21789 NAND2X1_LOC_553/A NAND2X1_LOC_74/B 0.01fF
C21790 INVX1_LOC_48/A NOR2X1_LOC_346/B 0.03fF
C21791 INVX1_LOC_233/Y INVX1_LOC_42/A 0.07fF
C21792 INVX1_LOC_11/A INVX1_LOC_123/Y 0.03fF
C21793 INVX1_LOC_239/A NOR2X1_LOC_662/A 0.37fF
C21794 NOR2X1_LOC_644/A INVX1_LOC_89/A 0.03fF
C21795 NOR2X1_LOC_131/Y INVX1_LOC_6/A 0.31fF
C21796 INVX1_LOC_23/A INVX1_LOC_4/A 0.03fF
C21797 NOR2X1_LOC_798/A NAND2X1_LOC_74/B 0.05fF
C21798 INVX1_LOC_227/A NAND2X1_LOC_132/a_36_24# 0.00fF
C21799 NAND2X1_LOC_787/A INVX1_LOC_15/A 0.03fF
C21800 NOR2X1_LOC_590/A INVX1_LOC_307/A 0.07fF
C21801 NOR2X1_LOC_298/Y NAND2X1_LOC_863/A 0.03fF
C21802 NOR2X1_LOC_643/A NOR2X1_LOC_814/A 0.07fF
C21803 NAND2X1_LOC_352/B NOR2X1_LOC_831/B 0.02fF
C21804 INVX1_LOC_27/A INVX1_LOC_29/A 7.67fF
C21805 NOR2X1_LOC_557/Y NOR2X1_LOC_558/A 0.01fF
C21806 NAND2X1_LOC_363/B INVX1_LOC_15/A 0.07fF
C21807 INVX1_LOC_53/A NAND2X1_LOC_647/B 0.01fF
C21808 INVX1_LOC_182/A INVX1_LOC_97/A 0.02fF
C21809 INVX1_LOC_77/A NAND2X1_LOC_639/A 0.07fF
C21810 NOR2X1_LOC_828/B INVX1_LOC_89/A 0.03fF
C21811 NOR2X1_LOC_590/A NOR2X1_LOC_445/B 0.12fF
C21812 NOR2X1_LOC_589/A INVX1_LOC_6/A 0.30fF
C21813 INVX1_LOC_206/Y NOR2X1_LOC_570/Y 0.00fF
C21814 NOR2X1_LOC_469/a_36_216# INVX1_LOC_63/A 0.00fF
C21815 INVX1_LOC_90/A INVX1_LOC_182/A 0.07fF
C21816 NOR2X1_LOC_87/B NOR2X1_LOC_35/Y 0.05fF
C21817 NOR2X1_LOC_6/B INVX1_LOC_2/Y 0.03fF
C21818 INVX1_LOC_77/A NOR2X1_LOC_536/A 0.06fF
C21819 INVX1_LOC_30/A NOR2X1_LOC_88/Y 0.07fF
C21820 NOR2X1_LOC_751/A INVX1_LOC_89/A 0.01fF
C21821 INVX1_LOC_289/A INVX1_LOC_187/A 0.02fF
C21822 NOR2X1_LOC_205/Y INVX1_LOC_263/Y 0.32fF
C21823 INVX1_LOC_18/A NOR2X1_LOC_88/a_36_216# 0.00fF
C21824 NOR2X1_LOC_348/Y INVX1_LOC_290/Y 0.04fF
C21825 NAND2X1_LOC_116/A NOR2X1_LOC_859/Y 0.01fF
C21826 NAND2X1_LOC_561/B INVX1_LOC_284/A 0.09fF
C21827 INVX1_LOC_31/A NOR2X1_LOC_68/a_36_216# 0.01fF
C21828 NAND2X1_LOC_420/a_36_24# INVX1_LOC_23/A 0.01fF
C21829 NOR2X1_LOC_154/a_36_216# INVX1_LOC_117/A 0.01fF
C21830 INVX1_LOC_30/A INVX1_LOC_84/A 0.18fF
C21831 INVX1_LOC_75/A NOR2X1_LOC_163/Y 0.07fF
C21832 NOR2X1_LOC_205/Y INVX1_LOC_42/A 0.03fF
C21833 NAND2X1_LOC_803/B INVX1_LOC_12/A 0.02fF
C21834 INVX1_LOC_33/A INVX1_LOC_54/A 2.27fF
C21835 INVX1_LOC_77/A NAND2X1_LOC_93/B 0.20fF
C21836 NAND2X1_LOC_392/A INVX1_LOC_126/A 0.01fF
C21837 INVX1_LOC_2/A INVX1_LOC_33/Y 0.42fF
C21838 NOR2X1_LOC_303/Y NOR2X1_LOC_155/A 0.03fF
C21839 NAND2X1_LOC_114/B NAND2X1_LOC_207/B 0.00fF
C21840 INVX1_LOC_45/A NOR2X1_LOC_691/B 0.07fF
C21841 NOR2X1_LOC_91/A INVX1_LOC_64/A 0.06fF
C21842 INVX1_LOC_35/A NOR2X1_LOC_400/B 0.01fF
C21843 INVX1_LOC_13/A INVX1_LOC_59/Y 0.09fF
C21844 INVX1_LOC_124/A NOR2X1_LOC_536/A 0.04fF
C21845 INVX1_LOC_58/A D_INPUT_1 0.05fF
C21846 NOR2X1_LOC_717/Y INVX1_LOC_186/Y 0.07fF
C21847 NOR2X1_LOC_644/A NOR2X1_LOC_703/Y 0.10fF
C21848 NOR2X1_LOC_52/B NOR2X1_LOC_142/a_36_216# 0.00fF
C21849 INVX1_LOC_1/A NOR2X1_LOC_467/A 0.08fF
C21850 NOR2X1_LOC_226/A INVX1_LOC_33/Y 0.03fF
C21851 INVX1_LOC_256/A INVX1_LOC_290/Y 0.10fF
C21852 INVX1_LOC_77/A NAND2X1_LOC_425/Y 0.10fF
C21853 NAND2X1_LOC_349/a_36_24# NAND2X1_LOC_211/Y 0.00fF
C21854 NOR2X1_LOC_620/B INVX1_LOC_117/A 0.03fF
C21855 NOR2X1_LOC_590/A INVX1_LOC_12/A 0.10fF
C21856 NOR2X1_LOC_286/a_36_216# INVX1_LOC_26/Y 0.00fF
C21857 NAND2X1_LOC_859/Y INVX1_LOC_20/A 0.03fF
C21858 INVX1_LOC_245/A VDD -0.00fF
C21859 NOR2X1_LOC_701/Y INVX1_LOC_46/A 0.01fF
C21860 INVX1_LOC_13/A INVX1_LOC_176/A 0.03fF
C21861 NOR2X1_LOC_19/B INVX1_LOC_201/A 0.04fF
C21862 INVX1_LOC_30/A NAND2X1_LOC_651/B 0.05fF
C21863 NOR2X1_LOC_454/Y NAND2X1_LOC_470/B 0.03fF
C21864 INVX1_LOC_217/Y NOR2X1_LOC_88/A 0.01fF
C21865 INVX1_LOC_41/A NOR2X1_LOC_461/A 0.01fF
C21866 NOR2X1_LOC_91/Y NOR2X1_LOC_662/A 0.19fF
C21867 INVX1_LOC_298/Y INVX1_LOC_27/A 0.07fF
C21868 NAND2X1_LOC_140/A NOR2X1_LOC_657/B 0.29fF
C21869 NOR2X1_LOC_78/A NOR2X1_LOC_356/A 0.09fF
C21870 NOR2X1_LOC_82/A INVX1_LOC_32/A 0.21fF
C21871 INVX1_LOC_64/A INVX1_LOC_23/A 0.53fF
C21872 NOR2X1_LOC_254/Y NOR2X1_LOC_155/A 0.03fF
C21873 NAND2X1_LOC_564/B NAND2X1_LOC_721/A 0.07fF
C21874 NOR2X1_LOC_457/A INVX1_LOC_15/A 0.01fF
C21875 NOR2X1_LOC_294/Y NAND2X1_LOC_207/B 0.03fF
C21876 INVX1_LOC_27/A NOR2X1_LOC_33/Y -0.00fF
C21877 INVX1_LOC_101/Y NOR2X1_LOC_334/Y 0.03fF
C21878 INVX1_LOC_278/A NAND2X1_LOC_787/A 0.04fF
C21879 INVX1_LOC_89/A NOR2X1_LOC_540/B 0.05fF
C21880 INVX1_LOC_49/A INVX1_LOC_220/A 0.44fF
C21881 INVX1_LOC_77/A INVX1_LOC_3/A 0.00fF
C21882 INVX1_LOC_223/A NOR2X1_LOC_89/A 0.07fF
C21883 NOR2X1_LOC_497/Y NAND2X1_LOC_623/B 0.03fF
C21884 NAND2X1_LOC_9/Y NAND2X1_LOC_358/B 0.01fF
C21885 NOR2X1_LOC_171/Y NOR2X1_LOC_45/B 0.09fF
C21886 NAND2X1_LOC_656/Y NAND2X1_LOC_211/Y 0.18fF
C21887 NAND2X1_LOC_35/Y NAND2X1_LOC_860/A 0.01fF
C21888 INVX1_LOC_124/A NAND2X1_LOC_93/B 0.03fF
C21889 NOR2X1_LOC_71/Y NAND2X1_LOC_244/A 0.27fF
C21890 NAND2X1_LOC_465/Y INVX1_LOC_35/Y 0.18fF
C21891 NOR2X1_LOC_234/Y INVX1_LOC_35/Y 0.04fF
C21892 NAND2X1_LOC_798/A INVX1_LOC_54/A 0.01fF
C21893 INVX1_LOC_299/A NOR2X1_LOC_541/B 0.02fF
C21894 INVX1_LOC_1/A INVX1_LOC_116/Y 0.03fF
C21895 NOR2X1_LOC_837/Y INVX1_LOC_19/A 0.01fF
C21896 NAND2X1_LOC_866/B INVX1_LOC_20/A 0.25fF
C21897 INVX1_LOC_230/Y NOR2X1_LOC_38/B 0.32fF
C21898 NOR2X1_LOC_760/a_36_216# NOR2X1_LOC_334/Y 0.00fF
C21899 INVX1_LOC_98/A NOR2X1_LOC_74/A -0.02fF
C21900 INVX1_LOC_31/A INVX1_LOC_4/A 3.70fF
C21901 NOR2X1_LOC_78/A NOR2X1_LOC_74/A 0.07fF
C21902 INVX1_LOC_97/Y INVX1_LOC_99/Y 0.11fF
C21903 NOR2X1_LOC_312/Y NOR2X1_LOC_111/A 0.01fF
C21904 INVX1_LOC_303/A INVX1_LOC_125/A 0.06fF
C21905 NOR2X1_LOC_788/B VDD 0.26fF
C21906 INVX1_LOC_30/A INVX1_LOC_15/A 8.93fF
C21907 NAND2X1_LOC_807/Y INVX1_LOC_20/A 0.52fF
C21908 INVX1_LOC_98/A NOR2X1_LOC_9/Y 0.12fF
C21909 INVX1_LOC_278/A NOR2X1_LOC_791/Y 0.08fF
C21910 INVX1_LOC_135/A NAND2X1_LOC_96/A 0.07fF
C21911 NOR2X1_LOC_228/a_36_216# NAND2X1_LOC_63/Y 0.00fF
C21912 NOR2X1_LOC_78/A NOR2X1_LOC_9/Y 0.11fF
C21913 NAND2X1_LOC_763/B INVX1_LOC_15/A 0.05fF
C21914 NAND2X1_LOC_357/A NAND2X1_LOC_288/B 0.01fF
C21915 INVX1_LOC_25/A INVX1_LOC_1/A 0.29fF
C21916 NOR2X1_LOC_99/B INVX1_LOC_38/A 0.08fF
C21917 NAND2X1_LOC_722/A INVX1_LOC_84/A 0.05fF
C21918 NAND2X1_LOC_564/a_36_24# INVX1_LOC_19/A -0.00fF
C21919 INVX1_LOC_232/A INVX1_LOC_46/Y 0.19fF
C21920 NOR2X1_LOC_135/Y VDD 0.53fF
C21921 NOR2X1_LOC_560/A NAND2X1_LOC_96/A -0.02fF
C21922 INVX1_LOC_36/A NOR2X1_LOC_248/A 0.01fF
C21923 NOR2X1_LOC_720/B INVX1_LOC_19/A 0.06fF
C21924 NOR2X1_LOC_134/Y INVX1_LOC_23/Y 0.02fF
C21925 NOR2X1_LOC_589/A INVX1_LOC_131/Y 0.07fF
C21926 NOR2X1_LOC_302/B INVX1_LOC_179/A 0.01fF
C21927 NOR2X1_LOC_516/B NOR2X1_LOC_820/a_36_216# 0.01fF
C21928 NOR2X1_LOC_554/B INVX1_LOC_4/Y 0.02fF
C21929 INVX1_LOC_136/A NOR2X1_LOC_282/a_36_216# 0.01fF
C21930 NOR2X1_LOC_233/a_36_216# NOR2X1_LOC_291/Y 0.01fF
C21931 NOR2X1_LOC_403/B INVX1_LOC_3/Y 0.02fF
C21932 D_INPUT_2 INVX1_LOC_3/Y 0.12fF
C21933 INVX1_LOC_295/A NAND2X1_LOC_427/a_36_24# 0.01fF
C21934 INVX1_LOC_111/A INVX1_LOC_4/A 0.02fF
C21935 NOR2X1_LOC_667/A INVX1_LOC_63/A 0.32fF
C21936 NOR2X1_LOC_780/B INVX1_LOC_213/A 0.00fF
C21937 NOR2X1_LOC_237/Y INVX1_LOC_19/Y 0.41fF
C21938 INVX1_LOC_16/A NAND2X1_LOC_572/B 0.07fF
C21939 INVX1_LOC_50/A INVX1_LOC_161/A 0.02fF
C21940 INVX1_LOC_248/A INVX1_LOC_63/A 0.06fF
C21941 INVX1_LOC_6/A INVX1_LOC_20/A 0.55fF
C21942 NOR2X1_LOC_763/Y NAND2X1_LOC_428/a_36_24# 0.00fF
C21943 NOR2X1_LOC_147/B NOR2X1_LOC_850/B 0.00fF
C21944 INVX1_LOC_206/A INVX1_LOC_29/A 0.03fF
C21945 INVX1_LOC_171/A NOR2X1_LOC_79/A 0.02fF
C21946 INVX1_LOC_43/Y INVX1_LOC_23/A 0.03fF
C21947 INVX1_LOC_22/A NOR2X1_LOC_127/Y 0.11fF
C21948 INVX1_LOC_35/A NOR2X1_LOC_103/Y 0.03fF
C21949 INVX1_LOC_182/A INVX1_LOC_38/A 0.07fF
C21950 NOR2X1_LOC_52/B INVX1_LOC_102/A 0.07fF
C21951 INVX1_LOC_89/A INVX1_LOC_89/Y 0.06fF
C21952 NOR2X1_LOC_147/A VDD 0.00fF
C21953 NAND2X1_LOC_332/Y INVX1_LOC_32/A 0.00fF
C21954 INVX1_LOC_77/A NAND2X1_LOC_470/B 0.01fF
C21955 INVX1_LOC_166/A INVX1_LOC_195/Y 0.03fF
C21956 NAND2X1_LOC_561/B NOR2X1_LOC_384/A 0.16fF
C21957 INVX1_LOC_249/A INVX1_LOC_298/Y 0.03fF
C21958 INVX1_LOC_50/A INVX1_LOC_79/Y 0.01fF
C21959 NAND2X1_LOC_808/A INVX1_LOC_285/A 0.02fF
C21960 NAND2X1_LOC_808/A INVX1_LOC_265/Y 0.00fF
C21961 INVX1_LOC_50/A NOR2X1_LOC_518/a_36_216# 0.00fF
C21962 INVX1_LOC_64/A INVX1_LOC_31/A 0.08fF
C21963 NOR2X1_LOC_837/Y INVX1_LOC_26/Y 0.06fF
C21964 NOR2X1_LOC_526/Y INVX1_LOC_42/A 0.03fF
C21965 NOR2X1_LOC_91/Y INVX1_LOC_57/A 0.03fF
C21966 NOR2X1_LOC_529/Y INVX1_LOC_3/Y 0.03fF
C21967 INVX1_LOC_278/A INVX1_LOC_30/A 0.56fF
C21968 NOR2X1_LOC_82/Y INVX1_LOC_12/A 0.02fF
C21969 INVX1_LOC_58/A NAND2X1_LOC_391/a_36_24# 0.00fF
C21970 INVX1_LOC_35/A INVX1_LOC_45/A 1.98fF
C21971 NOR2X1_LOC_439/B INVX1_LOC_179/A 0.25fF
C21972 NAND2X1_LOC_798/A NOR2X1_LOC_48/B 0.02fF
C21973 NAND2X1_LOC_9/Y INVX1_LOC_136/A 0.06fF
C21974 INVX1_LOC_119/A INVX1_LOC_21/Y 0.05fF
C21975 NAND2X1_LOC_862/A INVX1_LOC_42/A 0.00fF
C21976 INVX1_LOC_35/A NOR2X1_LOC_568/A 0.03fF
C21977 INVX1_LOC_177/A NOR2X1_LOC_609/Y 0.01fF
C21978 NOR2X1_LOC_309/Y NOR2X1_LOC_248/A 0.01fF
C21979 NOR2X1_LOC_703/A NOR2X1_LOC_445/B 0.02fF
C21980 NAND2X1_LOC_525/a_36_24# INVX1_LOC_92/A 0.01fF
C21981 INVX1_LOC_233/A INVX1_LOC_136/A 0.07fF
C21982 INVX1_LOC_75/A INVX1_LOC_179/A 0.03fF
C21983 NOR2X1_LOC_75/Y NAND2X1_LOC_149/Y 0.02fF
C21984 INVX1_LOC_88/A NAND2X1_LOC_538/Y 0.02fF
C21985 NOR2X1_LOC_167/Y INVX1_LOC_185/A 0.05fF
C21986 NOR2X1_LOC_577/Y NOR2X1_LOC_383/B 0.25fF
C21987 INVX1_LOC_234/A INVX1_LOC_29/A 0.19fF
C21988 NOR2X1_LOC_274/Y INVX1_LOC_129/A 0.11fF
C21989 INVX1_LOC_227/A INVX1_LOC_12/A 0.07fF
C21990 NOR2X1_LOC_500/A NOR2X1_LOC_598/B 0.10fF
C21991 NOR2X1_LOC_739/Y NOR2X1_LOC_740/Y 0.01fF
C21992 NOR2X1_LOC_598/B NOR2X1_LOC_303/Y 0.43fF
C21993 NAND2X1_LOC_462/B NAND2X1_LOC_410/a_36_24# 0.00fF
C21994 INVX1_LOC_298/Y INVX1_LOC_206/A 0.02fF
C21995 INVX1_LOC_34/A INVX1_LOC_50/A 4.21fF
C21996 INVX1_LOC_174/Y NOR2X1_LOC_460/a_36_216# 0.00fF
C21997 NAND2X1_LOC_144/a_36_24# INVX1_LOC_92/A 0.01fF
C21998 INVX1_LOC_35/A INVX1_LOC_71/A 0.20fF
C21999 INVX1_LOC_136/A NOR2X1_LOC_798/A 0.03fF
C22000 NOR2X1_LOC_544/A NOR2X1_LOC_334/Y 0.03fF
C22001 NOR2X1_LOC_479/B NAND2X1_LOC_618/Y 0.05fF
C22002 INVX1_LOC_211/Y INVX1_LOC_103/A 0.09fF
C22003 INVX1_LOC_35/A NOR2X1_LOC_707/a_36_216# 0.00fF
C22004 INVX1_LOC_2/A INVX1_LOC_23/Y 0.16fF
C22005 NOR2X1_LOC_708/Y NAND2X1_LOC_782/a_36_24# 0.00fF
C22006 NOR2X1_LOC_824/A NAND2X1_LOC_634/Y 0.10fF
C22007 NOR2X1_LOC_790/B NOR2X1_LOC_344/A 0.14fF
C22008 NOR2X1_LOC_772/A INVX1_LOC_29/A 0.00fF
C22009 NOR2X1_LOC_82/A INPUT_3 0.67fF
C22010 INVX1_LOC_116/A NOR2X1_LOC_220/B 0.04fF
C22011 NOR2X1_LOC_19/B INVX1_LOC_29/A 1.95fF
C22012 NOR2X1_LOC_91/A NAND2X1_LOC_850/Y 0.04fF
C22013 NAND2X1_LOC_860/A NOR2X1_LOC_234/Y -0.02fF
C22014 INVX1_LOC_50/A NAND2X1_LOC_231/Y 0.01fF
C22015 NOR2X1_LOC_92/Y NOR2X1_LOC_68/A 0.07fF
C22016 NOR2X1_LOC_78/A NOR2X1_LOC_865/Y 0.08fF
C22017 INVX1_LOC_97/Y NOR2X1_LOC_254/Y 0.15fF
C22018 NOR2X1_LOC_741/a_36_216# INVX1_LOC_12/A 0.00fF
C22019 INVX1_LOC_5/A INVX1_LOC_207/A 0.03fF
C22020 NOR2X1_LOC_454/Y NOR2X1_LOC_781/Y 0.04fF
C22021 NOR2X1_LOC_78/A NOR2X1_LOC_243/B 0.07fF
C22022 INVX1_LOC_14/A INVX1_LOC_18/A 0.08fF
C22023 INVX1_LOC_233/A NOR2X1_LOC_278/A 0.04fF
C22024 NAND2X1_LOC_149/Y NAND2X1_LOC_162/B 0.08fF
C22025 INVX1_LOC_11/A INVX1_LOC_223/A 0.03fF
C22026 NOR2X1_LOC_689/A INVX1_LOC_22/A 0.01fF
C22027 NOR2X1_LOC_598/B INVX1_LOC_54/Y 0.00fF
C22028 NAND2X1_LOC_850/Y INVX1_LOC_23/A 0.07fF
C22029 NOR2X1_LOC_658/Y NOR2X1_LOC_160/B 0.07fF
C22030 NAND2X1_LOC_342/Y INVX1_LOC_53/A 0.03fF
C22031 NAND2X1_LOC_363/B NOR2X1_LOC_16/Y 0.03fF
C22032 INVX1_LOC_40/A NAND2X1_LOC_215/A 0.46fF
C22033 NOR2X1_LOC_325/A NOR2X1_LOC_383/B 0.04fF
C22034 NAND2X1_LOC_208/B INVX1_LOC_61/Y 0.03fF
C22035 NOR2X1_LOC_516/B NOR2X1_LOC_105/a_36_216# 0.01fF
C22036 INVX1_LOC_190/A NAND2X1_LOC_470/B 0.07fF
C22037 NOR2X1_LOC_99/B NAND2X1_LOC_223/A 0.07fF
C22038 INVX1_LOC_22/A NOR2X1_LOC_383/B 0.13fF
C22039 NOR2X1_LOC_186/Y INVX1_LOC_294/Y 0.01fF
C22040 INVX1_LOC_151/Y INVX1_LOC_271/A 0.01fF
C22041 INVX1_LOC_33/Y INVX1_LOC_118/A 0.08fF
C22042 INVX1_LOC_224/Y NOR2X1_LOC_121/A 0.02fF
C22043 NOR2X1_LOC_845/A NOR2X1_LOC_721/B 0.01fF
C22044 NOR2X1_LOC_772/B NOR2X1_LOC_709/A 0.10fF
C22045 NAND2X1_LOC_810/B INVX1_LOC_20/A 0.03fF
C22046 NOR2X1_LOC_536/A INVX1_LOC_9/A 0.96fF
C22047 INVX1_LOC_27/A INVX1_LOC_8/A 0.15fF
C22048 INVX1_LOC_140/A D_INPUT_5 0.17fF
C22049 NOR2X1_LOC_816/Y INVX1_LOC_54/A 0.02fF
C22050 NOR2X1_LOC_91/A NOR2X1_LOC_700/a_36_216# 0.00fF
C22051 INVX1_LOC_208/A NOR2X1_LOC_717/A 0.10fF
C22052 NAND2X1_LOC_587/a_36_24# INVX1_LOC_174/A 0.01fF
C22053 INVX1_LOC_13/Y NOR2X1_LOC_709/A 0.17fF
C22054 NOR2X1_LOC_590/A NAND2X1_LOC_355/Y 0.02fF
C22055 INVX1_LOC_104/A NAND2X1_LOC_474/Y 0.01fF
C22056 INVX1_LOC_28/A NOR2X1_LOC_394/Y 0.01fF
C22057 INVX1_LOC_5/A NAND2X1_LOC_451/Y -0.04fF
C22058 INVX1_LOC_89/A INVX1_LOC_16/Y 0.56fF
C22059 NOR2X1_LOC_784/B NOR2X1_LOC_383/B 0.00fF
C22060 INVX1_LOC_256/A INVX1_LOC_77/A 0.16fF
C22061 D_INPUT_0 INVX1_LOC_112/Y 0.01fF
C22062 NOR2X1_LOC_438/a_36_216# NOR2X1_LOC_716/B 0.01fF
C22063 INVX1_LOC_255/Y NOR2X1_LOC_392/Y 2.37fF
C22064 INPUT_1 INVX1_LOC_23/Y 0.21fF
C22065 NOR2X1_LOC_138/a_36_216# NOR2X1_LOC_649/B 0.03fF
C22066 NAND2X1_LOC_51/B NAND2X1_LOC_452/Y 0.04fF
C22067 NAND2X1_LOC_140/A INVX1_LOC_271/A 0.02fF
C22068 NAND2X1_LOC_93/B INVX1_LOC_9/A 0.07fF
C22069 NAND2X1_LOC_364/Y NOR2X1_LOC_160/B 0.03fF
C22070 INVX1_LOC_64/A NAND2X1_LOC_859/Y 0.00fF
C22071 NOR2X1_LOC_795/Y INVX1_LOC_299/A 0.05fF
C22072 INVX1_LOC_161/Y INVX1_LOC_155/Y 0.03fF
C22073 NOR2X1_LOC_384/Y NOR2X1_LOC_522/a_36_216# 0.00fF
C22074 INVX1_LOC_89/A NAND2X1_LOC_205/A 0.03fF
C22075 INVX1_LOC_11/A INVX1_LOC_149/Y 0.02fF
C22076 INVX1_LOC_6/A INVX1_LOC_4/A 0.14fF
C22077 NOR2X1_LOC_516/B NOR2X1_LOC_649/Y 0.10fF
C22078 NOR2X1_LOC_391/a_36_216# NOR2X1_LOC_38/B 0.00fF
C22079 INVX1_LOC_24/A NAND2X1_LOC_311/a_36_24# 0.00fF
C22080 INVX1_LOC_11/A INVX1_LOC_162/Y 0.01fF
C22081 NAND2X1_LOC_794/B NOR2X1_LOC_165/Y 0.03fF
C22082 INVX1_LOC_18/A NOR2X1_LOC_522/Y 0.19fF
C22083 INVX1_LOC_11/A INVX1_LOC_85/A 0.05fF
C22084 NOR2X1_LOC_329/B NOR2X1_LOC_106/a_36_216# 0.01fF
C22085 INVX1_LOC_286/Y NOR2X1_LOC_753/Y 0.16fF
C22086 INVX1_LOC_72/A NOR2X1_LOC_759/Y 0.03fF
C22087 INVX1_LOC_14/A INVX1_LOC_34/Y 0.14fF
C22088 INVX1_LOC_28/A NOR2X1_LOC_654/A 0.10fF
C22089 NOR2X1_LOC_13/Y NAND2X1_LOC_195/Y 0.01fF
C22090 NOR2X1_LOC_792/B NAND2X1_LOC_337/B 0.02fF
C22091 NOR2X1_LOC_264/Y NAND2X1_LOC_114/B 0.08fF
C22092 INVX1_LOC_27/A NAND2X1_LOC_158/a_36_24# 0.00fF
C22093 INVX1_LOC_202/A INVX1_LOC_72/A 0.08fF
C22094 NOR2X1_LOC_441/Y INVX1_LOC_33/A 0.03fF
C22095 NAND2X1_LOC_350/A NAND2X1_LOC_466/A 0.03fF
C22096 NAND2X1_LOC_728/Y NAND2X1_LOC_739/B 0.05fF
C22097 NOR2X1_LOC_456/Y INVX1_LOC_313/Y 0.01fF
C22098 INVX1_LOC_90/A INVX1_LOC_308/A 0.02fF
C22099 NOR2X1_LOC_246/Y INVX1_LOC_53/A 0.01fF
C22100 INVX1_LOC_286/Y NAND2X1_LOC_325/Y 0.07fF
C22101 NOR2X1_LOC_91/A INVX1_LOC_282/A 0.01fF
C22102 NOR2X1_LOC_723/Y INVX1_LOC_113/Y 0.00fF
C22103 NOR2X1_LOC_763/A INVX1_LOC_22/A 0.01fF
C22104 INVX1_LOC_64/A INVX1_LOC_313/A 0.00fF
C22105 NAND2X1_LOC_357/B NAND2X1_LOC_352/B 0.30fF
C22106 NOR2X1_LOC_401/A INVX1_LOC_256/Y 0.11fF
C22107 INVX1_LOC_223/A NOR2X1_LOC_593/Y 0.17fF
C22108 INVX1_LOC_3/A INVX1_LOC_9/A 0.07fF
C22109 INVX1_LOC_299/A NOR2X1_LOC_614/Y 0.00fF
C22110 NOR2X1_LOC_78/A NOR2X1_LOC_855/A 1.72fF
C22111 INVX1_LOC_64/A NAND2X1_LOC_866/B 0.07fF
C22112 NOR2X1_LOC_598/B NOR2X1_LOC_112/Y 0.14fF
C22113 NAND2X1_LOC_344/a_36_24# INVX1_LOC_234/A 0.00fF
C22114 NAND2X1_LOC_763/B NAND2X1_LOC_21/Y 0.05fF
C22115 INVX1_LOC_30/A NAND2X1_LOC_464/Y 0.10fF
C22116 NAND2X1_LOC_172/a_36_24# INVX1_LOC_53/A 0.00fF
C22117 NOR2X1_LOC_45/B INVX1_LOC_94/Y 0.03fF
C22118 NOR2X1_LOC_139/Y NOR2X1_LOC_334/Y 0.04fF
C22119 INVX1_LOC_172/A NOR2X1_LOC_522/Y 0.06fF
C22120 NOR2X1_LOC_470/A NAND2X1_LOC_149/Y 0.06fF
C22121 INVX1_LOC_2/A NOR2X1_LOC_596/Y 0.01fF
C22122 INVX1_LOC_21/A NAND2X1_LOC_554/a_36_24# 0.00fF
C22123 INVX1_LOC_229/A GATE_865 0.06fF
C22124 INVX1_LOC_59/Y INVX1_LOC_32/A 0.11fF
C22125 NOR2X1_LOC_781/Y INVX1_LOC_77/A 0.26fF
C22126 INVX1_LOC_50/A INPUT_0 13.59fF
C22127 INVX1_LOC_112/A INVX1_LOC_32/A 0.01fF
C22128 NOR2X1_LOC_577/Y NOR2X1_LOC_512/Y 0.01fF
C22129 NOR2X1_LOC_609/Y NOR2X1_LOC_137/B 0.02fF
C22130 NAND2X1_LOC_149/Y NOR2X1_LOC_424/Y 0.06fF
C22131 INVX1_LOC_41/A NOR2X1_LOC_68/A 0.21fF
C22132 NOR2X1_LOC_488/Y INVX1_LOC_200/A 0.16fF
C22133 NOR2X1_LOC_595/Y INVX1_LOC_78/A 0.03fF
C22134 NAND2X1_LOC_350/A NAND2X1_LOC_798/A 0.03fF
C22135 NOR2X1_LOC_570/a_36_216# NOR2X1_LOC_570/B 0.00fF
C22136 NOR2X1_LOC_160/B INVX1_LOC_256/Y 0.03fF
C22137 INVX1_LOC_285/A INVX1_LOC_92/A 0.03fF
C22138 INVX1_LOC_35/A INVX1_LOC_102/Y 0.39fF
C22139 INVX1_LOC_27/A NAND2X1_LOC_140/A 0.01fF
C22140 INVX1_LOC_223/A NOR2X1_LOC_52/B 0.01fF
C22141 NOR2X1_LOC_635/A D_INPUT_7 0.00fF
C22142 NOR2X1_LOC_194/Y NAND2X1_LOC_16/Y 0.02fF
C22143 INVX1_LOC_67/Y INVX1_LOC_53/A 0.01fF
C22144 NOR2X1_LOC_607/a_36_216# NOR2X1_LOC_577/Y 0.01fF
C22145 INVX1_LOC_181/Y NOR2X1_LOC_557/Y 0.13fF
C22146 NOR2X1_LOC_226/A NAND2X1_LOC_543/a_36_24# 0.01fF
C22147 NOR2X1_LOC_16/Y INVX1_LOC_30/A 0.11fF
C22148 NOR2X1_LOC_814/A INVX1_LOC_92/A 7.24fF
C22149 INVX1_LOC_31/A NAND2X1_LOC_850/Y 0.05fF
C22150 NOR2X1_LOC_405/A NOR2X1_LOC_278/Y 0.07fF
C22151 NOR2X1_LOC_75/Y INVX1_LOC_16/A 0.00fF
C22152 NAND2X1_LOC_594/a_36_24# INVX1_LOC_90/A 0.00fF
C22153 NAND2X1_LOC_860/A NOR2X1_LOC_83/Y 0.03fF
C22154 NOR2X1_LOC_80/Y INVX1_LOC_20/A 0.01fF
C22155 NAND2X1_LOC_341/A NOR2X1_LOC_389/A 0.02fF
C22156 INVX1_LOC_41/A NOR2X1_LOC_545/A 0.01fF
C22157 INVX1_LOC_34/A INVX1_LOC_105/A 0.10fF
C22158 NOR2X1_LOC_510/Y NOR2X1_LOC_135/Y 0.00fF
C22159 INVX1_LOC_111/Y INVX1_LOC_18/A 0.09fF
C22160 INVX1_LOC_58/A NOR2X1_LOC_144/a_36_216# 0.12fF
C22161 NOR2X1_LOC_214/a_36_216# INVX1_LOC_63/Y 0.01fF
C22162 NAND2X1_LOC_579/A INVX1_LOC_90/A 0.02fF
C22163 NAND2X1_LOC_802/A NAND2X1_LOC_799/Y 0.10fF
C22164 NAND2X1_LOC_99/Y INVX1_LOC_8/A 0.03fF
C22165 INVX1_LOC_64/A INVX1_LOC_6/A 0.22fF
C22166 INVX1_LOC_50/A NAND2X1_LOC_649/B 0.01fF
C22167 INVX1_LOC_235/Y INVX1_LOC_135/Y 0.03fF
C22168 INVX1_LOC_21/A NOR2X1_LOC_742/A 0.07fF
C22169 INVX1_LOC_36/A NOR2X1_LOC_418/Y 0.02fF
C22170 INVX1_LOC_33/A NOR2X1_LOC_142/Y 0.06fF
C22171 NAND2X1_LOC_803/B NAND2X1_LOC_808/A 0.02fF
C22172 INVX1_LOC_49/A NAND2X1_LOC_116/A 0.03fF
C22173 INVX1_LOC_181/Y INVX1_LOC_143/A 0.00fF
C22174 NOR2X1_LOC_817/Y INVX1_LOC_89/A 0.43fF
C22175 NAND2X1_LOC_588/B NAND2X1_LOC_588/a_36_24# 0.01fF
C22176 NOR2X1_LOC_78/B NOR2X1_LOC_791/a_36_216# 0.00fF
C22177 NOR2X1_LOC_395/Y INVX1_LOC_46/A 0.05fF
C22178 NOR2X1_LOC_216/B INVX1_LOC_29/A 0.05fF
C22179 NOR2X1_LOC_593/Y INVX1_LOC_149/Y 0.01fF
C22180 NAND2X1_LOC_687/A INVX1_LOC_273/A 0.01fF
C22181 NAND2X1_LOC_36/A GATE_662 0.03fF
C22182 NOR2X1_LOC_593/Y INVX1_LOC_85/A 0.02fF
C22183 NOR2X1_LOC_794/a_36_216# INVX1_LOC_177/A 0.00fF
C22184 INVX1_LOC_45/A NOR2X1_LOC_188/Y 0.01fF
C22185 NAND2X1_LOC_57/a_36_24# INVX1_LOC_137/A 0.01fF
C22186 NOR2X1_LOC_78/A NOR2X1_LOC_342/A 0.09fF
C22187 VDD NAND2X1_LOC_61/Y 0.03fF
C22188 INVX1_LOC_36/A NOR2X1_LOC_589/A 0.13fF
C22189 NOR2X1_LOC_661/a_36_216# NOR2X1_LOC_662/A 0.02fF
C22190 NOR2X1_LOC_590/A NAND2X1_LOC_808/A 0.00fF
C22191 NOR2X1_LOC_186/Y NOR2X1_LOC_9/Y 0.16fF
C22192 NAND2X1_LOC_231/Y INVX1_LOC_105/A 0.02fF
C22193 INVX1_LOC_225/A INVX1_LOC_294/Y 0.01fF
C22194 NOR2X1_LOC_92/Y INVX1_LOC_147/A 0.10fF
C22195 INVX1_LOC_37/A NOR2X1_LOC_621/A 0.04fF
C22196 INVX1_LOC_290/A NOR2X1_LOC_194/a_36_216# 0.00fF
C22197 NOR2X1_LOC_267/A NOR2X1_LOC_589/A 0.08fF
C22198 INVX1_LOC_179/A INVX1_LOC_283/A 0.00fF
C22199 INVX1_LOC_5/A NAND2X1_LOC_677/a_36_24# 0.00fF
C22200 INVX1_LOC_315/Y NOR2X1_LOC_649/Y 0.03fF
C22201 NOR2X1_LOC_761/Y NAND2X1_LOC_809/A 0.18fF
C22202 INVX1_LOC_60/Y NOR2X1_LOC_6/B 0.44fF
C22203 INVX1_LOC_55/Y INVX1_LOC_292/A 0.06fF
C22204 INVX1_LOC_266/A NOR2X1_LOC_541/a_36_216# 0.00fF
C22205 NAND2X1_LOC_477/Y INVX1_LOC_29/A 0.03fF
C22206 NOR2X1_LOC_79/A INVX1_LOC_4/A 0.03fF
C22207 NOR2X1_LOC_666/Y NOR2X1_LOC_151/a_36_216# 0.02fF
C22208 NOR2X1_LOC_468/Y NOR2X1_LOC_292/Y 0.08fF
C22209 INVX1_LOC_177/Y INVX1_LOC_10/A 0.07fF
C22210 NOR2X1_LOC_360/A NOR2X1_LOC_416/A 0.01fF
C22211 INVX1_LOC_1/A NOR2X1_LOC_188/A 0.01fF
C22212 NOR2X1_LOC_68/A INVX1_LOC_121/A 0.02fF
C22213 NOR2X1_LOC_35/Y INVX1_LOC_58/Y 0.10fF
C22214 VDD NOR2X1_LOC_452/A 0.24fF
C22215 INVX1_LOC_145/A NOR2X1_LOC_589/A 0.01fF
C22216 INVX1_LOC_1/A NOR2X1_LOC_548/B 0.05fF
C22217 INVX1_LOC_21/A NOR2X1_LOC_318/B 0.11fF
C22218 NAND2X1_LOC_642/Y INVX1_LOC_306/Y 0.08fF
C22219 NAND2X1_LOC_588/B INVX1_LOC_83/A 0.22fF
C22220 INVX1_LOC_71/A NOR2X1_LOC_188/Y 0.01fF
C22221 NAND2X1_LOC_200/B INVX1_LOC_8/A 0.03fF
C22222 NOR2X1_LOC_137/A INVX1_LOC_18/A 0.03fF
C22223 INVX1_LOC_255/Y NOR2X1_LOC_554/a_36_216# 0.00fF
C22224 NOR2X1_LOC_716/B INVX1_LOC_16/A 0.07fF
C22225 INVX1_LOC_20/A NOR2X1_LOC_109/Y 0.08fF
C22226 INVX1_LOC_23/Y INVX1_LOC_118/A 0.09fF
C22227 INVX1_LOC_21/A INVX1_LOC_93/Y 0.07fF
C22228 NAND2X1_LOC_610/a_36_24# NOR2X1_LOC_709/A 0.00fF
C22229 NAND2X1_LOC_656/Y NOR2X1_LOC_363/a_36_216# 0.01fF
C22230 INVX1_LOC_135/A NAND2X1_LOC_656/A 0.05fF
C22231 NOR2X1_LOC_177/a_36_216# NOR2X1_LOC_438/Y 0.00fF
C22232 INVX1_LOC_136/A NAND2X1_LOC_842/B 0.05fF
C22233 NOR2X1_LOC_460/B INVX1_LOC_174/Y 0.01fF
C22234 NOR2X1_LOC_156/Y INVX1_LOC_78/A 0.01fF
C22235 NOR2X1_LOC_794/B NOR2X1_LOC_188/A 0.00fF
C22236 INVX1_LOC_104/A NOR2X1_LOC_500/Y 0.09fF
C22237 NOR2X1_LOC_632/Y INVX1_LOC_153/Y 0.03fF
C22238 NAND2X1_LOC_53/Y INVX1_LOC_206/Y 0.08fF
C22239 NOR2X1_LOC_15/Y NOR2X1_LOC_192/A 0.01fF
C22240 INVX1_LOC_8/A INVX1_LOC_137/A 0.00fF
C22241 NOR2X1_LOC_678/A INVX1_LOC_117/A 0.03fF
C22242 INVX1_LOC_284/A NAND2X1_LOC_74/B 0.03fF
C22243 INVX1_LOC_271/A INVX1_LOC_118/Y 0.00fF
C22244 INVX1_LOC_304/Y NOR2X1_LOC_488/Y 0.11fF
C22245 INVX1_LOC_209/Y NOR2X1_LOC_298/Y 0.05fF
C22246 NOR2X1_LOC_78/B NAND2X1_LOC_342/Y 0.05fF
C22247 NAND2X1_LOC_358/Y INVX1_LOC_33/A 0.01fF
C22248 INVX1_LOC_61/Y INPUT_0 0.07fF
C22249 NAND2X1_LOC_543/Y NOR2X1_LOC_52/B 0.02fF
C22250 INVX1_LOC_41/A NOR2X1_LOC_545/a_36_216# 0.00fF
C22251 NOR2X1_LOC_504/Y NAND2X1_LOC_853/Y 0.30fF
C22252 INVX1_LOC_43/Y INVX1_LOC_6/A 0.01fF
C22253 NOR2X1_LOC_764/Y INVX1_LOC_77/A 0.01fF
C22254 NAND2X1_LOC_180/a_36_24# NAND2X1_LOC_564/B 0.00fF
C22255 NOR2X1_LOC_589/A NOR2X1_LOC_309/Y 0.03fF
C22256 INVX1_LOC_45/A NOR2X1_LOC_534/a_36_216# 0.00fF
C22257 NOR2X1_LOC_655/B INVX1_LOC_40/A 0.05fF
C22258 INVX1_LOC_269/A NOR2X1_LOC_396/Y 0.22fF
C22259 NAND2X1_LOC_479/Y NOR2X1_LOC_423/Y 0.03fF
C22260 NOR2X1_LOC_89/A INVX1_LOC_290/Y 0.07fF
C22261 INVX1_LOC_234/A INVX1_LOC_8/A 0.45fF
C22262 INVX1_LOC_35/A NOR2X1_LOC_331/B 0.07fF
C22263 D_INPUT_0 NAND2X1_LOC_139/A 0.05fF
C22264 INVX1_LOC_313/Y NOR2X1_LOC_550/B 0.10fF
C22265 INVX1_LOC_104/A INVX1_LOC_10/A 1.05fF
C22266 INVX1_LOC_124/A NOR2X1_LOC_440/Y 0.18fF
C22267 NOR2X1_LOC_669/a_36_216# NOR2X1_LOC_305/Y 0.00fF
C22268 NOR2X1_LOC_757/Y INVX1_LOC_16/A 0.19fF
C22269 NOR2X1_LOC_222/Y NAND2X1_LOC_479/Y 0.12fF
C22270 NOR2X1_LOC_716/B INVX1_LOC_28/A 0.07fF
C22271 NOR2X1_LOC_309/Y INVX1_LOC_171/A 1.60fF
C22272 INVX1_LOC_124/Y INVX1_LOC_98/A 0.14fF
C22273 NOR2X1_LOC_836/Y NOR2X1_LOC_836/B 0.04fF
C22274 INVX1_LOC_306/Y NOR2X1_LOC_271/Y 0.07fF
C22275 NOR2X1_LOC_226/A NOR2X1_LOC_383/Y 0.00fF
C22276 NOR2X1_LOC_364/A INVX1_LOC_53/A 0.11fF
C22277 NOR2X1_LOC_772/B NOR2X1_LOC_489/A 0.01fF
C22278 INVX1_LOC_103/A NOR2X1_LOC_357/Y 0.10fF
C22279 INVX1_LOC_2/A NOR2X1_LOC_366/Y 0.02fF
C22280 NOR2X1_LOC_793/Y VDD 0.12fF
C22281 INVX1_LOC_269/A INVX1_LOC_37/A 0.14fF
C22282 INVX1_LOC_41/A NAND2X1_LOC_150/a_36_24# 0.00fF
C22283 INVX1_LOC_200/A NAND2X1_LOC_650/B 0.02fF
C22284 INPUT_3 INVX1_LOC_59/Y 0.02fF
C22285 INVX1_LOC_143/A INVX1_LOC_148/Y 0.01fF
C22286 NOR2X1_LOC_788/B INVX1_LOC_177/A 0.00fF
C22287 INVX1_LOC_122/Y NOR2X1_LOC_349/A 0.09fF
C22288 NOR2X1_LOC_328/Y INPUT_5 0.00fF
C22289 INVX1_LOC_57/A NOR2X1_LOC_661/a_36_216# 0.00fF
C22290 NAND2X1_LOC_579/A NAND2X1_LOC_849/B 0.12fF
C22291 D_INPUT_1 NAND2X1_LOC_475/Y 0.04fF
C22292 NOR2X1_LOC_383/B INVX1_LOC_186/Y 0.07fF
C22293 NOR2X1_LOC_667/Y INVX1_LOC_76/A 0.01fF
C22294 INVX1_LOC_53/A INVX1_LOC_285/A 0.03fF
C22295 NAND2X1_LOC_579/A INVX1_LOC_38/A 0.07fF
C22296 NOR2X1_LOC_380/Y GATE_811 0.03fF
C22297 INVX1_LOC_299/A INVX1_LOC_299/Y 0.04fF
C22298 NAND2X1_LOC_640/Y NOR2X1_LOC_74/A -0.00fF
C22299 INVX1_LOC_40/A NOR2X1_LOC_99/B 0.00fF
C22300 INVX1_LOC_69/Y INVX1_LOC_77/A 0.07fF
C22301 NAND2X1_LOC_654/B INVX1_LOC_266/Y 0.02fF
C22302 NOR2X1_LOC_222/Y INVX1_LOC_295/A 0.10fF
C22303 INVX1_LOC_132/A NOR2X1_LOC_9/Y 0.83fF
C22304 NOR2X1_LOC_78/B NOR2X1_LOC_246/Y 0.01fF
C22305 INVX1_LOC_53/A NOR2X1_LOC_814/A 0.09fF
C22306 NAND2X1_LOC_861/Y NAND2X1_LOC_862/A 0.01fF
C22307 NOR2X1_LOC_15/Y NAND2X1_LOC_276/a_36_24# 0.00fF
C22308 NOR2X1_LOC_717/B INVX1_LOC_16/A 0.00fF
C22309 NOR2X1_LOC_700/Y NOR2X1_LOC_701/Y 0.01fF
C22310 NOR2X1_LOC_71/Y INVX1_LOC_25/Y 0.10fF
C22311 NOR2X1_LOC_523/A NOR2X1_LOC_865/A 0.00fF
C22312 NOR2X1_LOC_383/B NOR2X1_LOC_777/B 0.09fF
C22313 NOR2X1_LOC_858/A INVX1_LOC_19/A 0.00fF
C22314 NOR2X1_LOC_202/Y NOR2X1_LOC_423/Y 0.06fF
C22315 D_INPUT_0 NAND2X1_LOC_112/Y 0.00fF
C22316 INVX1_LOC_36/A INVX1_LOC_20/A 1.90fF
C22317 NOR2X1_LOC_1/Y INVX1_LOC_296/A 0.07fF
C22318 INVX1_LOC_147/A NAND2X1_LOC_477/A 0.02fF
C22319 NAND2X1_LOC_651/a_36_24# NAND2X1_LOC_451/Y 0.00fF
C22320 NOR2X1_LOC_658/Y NAND2X1_LOC_211/Y 0.15fF
C22321 INVX1_LOC_78/A D_INPUT_5 0.03fF
C22322 INVX1_LOC_55/A INVX1_LOC_117/A 0.04fF
C22323 NOR2X1_LOC_824/A NAND2X1_LOC_244/a_36_24# 0.01fF
C22324 INVX1_LOC_77/A NOR2X1_LOC_725/A 0.20fF
C22325 INVX1_LOC_28/A NOR2X1_LOC_757/Y 0.04fF
C22326 INVX1_LOC_49/A INVX1_LOC_186/A 0.06fF
C22327 NOR2X1_LOC_80/Y INVX1_LOC_4/A 0.19fF
C22328 INVX1_LOC_13/A INVX1_LOC_120/A 0.03fF
C22329 INVX1_LOC_232/A INPUT_1 0.07fF
C22330 NOR2X1_LOC_244/a_36_216# NAND2X1_LOC_348/A 0.01fF
C22331 NOR2X1_LOC_772/B INVX1_LOC_294/A 0.05fF
C22332 INVX1_LOC_225/A NOR2X1_LOC_9/Y 0.12fF
C22333 NAND2X1_LOC_361/Y INVX1_LOC_125/Y 0.02fF
C22334 INVX1_LOC_256/A INVX1_LOC_9/A 0.18fF
C22335 NAND2X1_LOC_67/Y NAND2X1_LOC_93/B 0.07fF
C22336 NOR2X1_LOC_48/B NOR2X1_LOC_635/B 0.02fF
C22337 NOR2X1_LOC_222/Y NOR2X1_LOC_202/Y 0.01fF
C22338 INVX1_LOC_57/A NOR2X1_LOC_461/Y 0.05fF
C22339 NOR2X1_LOC_209/Y NOR2X1_LOC_74/A 0.10fF
C22340 NAND2X1_LOC_577/A NOR2X1_LOC_813/Y 0.02fF
C22341 NOR2X1_LOC_383/Y INPUT_1 0.46fF
C22342 INVX1_LOC_124/A INVX1_LOC_69/Y 0.14fF
C22343 INVX1_LOC_299/A NOR2X1_LOC_862/B 0.05fF
C22344 INVX1_LOC_180/A NOR2X1_LOC_56/Y 0.03fF
C22345 NOR2X1_LOC_238/Y NAND2X1_LOC_241/Y 0.21fF
C22346 INVX1_LOC_36/A NOR2X1_LOC_765/Y 0.08fF
C22347 NAND2X1_LOC_102/a_36_24# INVX1_LOC_40/A 0.00fF
C22348 INVX1_LOC_64/A NOR2X1_LOC_633/A 0.03fF
C22349 INVX1_LOC_271/Y NOR2X1_LOC_464/Y 0.04fF
C22350 NOR2X1_LOC_725/A NOR2X1_LOC_732/A 0.00fF
C22351 INVX1_LOC_24/A NAND2X1_LOC_254/a_36_24# 0.00fF
C22352 NAND2X1_LOC_577/A INVX1_LOC_280/A 0.03fF
C22353 NOR2X1_LOC_557/Y NOR2X1_LOC_675/A 0.37fF
C22354 NOR2X1_LOC_419/Y NOR2X1_LOC_35/Y 0.03fF
C22355 NOR2X1_LOC_146/Y NOR2X1_LOC_706/A 0.02fF
C22356 NOR2X1_LOC_151/Y INVX1_LOC_16/A 0.85fF
C22357 INVX1_LOC_305/A INVX1_LOC_117/A 0.08fF
C22358 INVX1_LOC_99/Y INVX1_LOC_29/A 0.26fF
C22359 NOR2X1_LOC_237/Y INVX1_LOC_20/A 0.12fF
C22360 NOR2X1_LOC_860/B INVX1_LOC_2/Y 0.18fF
C22361 NOR2X1_LOC_441/Y NOR2X1_LOC_351/Y 0.00fF
C22362 NOR2X1_LOC_315/Y NOR2X1_LOC_45/B 0.03fF
C22363 INVX1_LOC_255/Y INVX1_LOC_75/A 0.03fF
C22364 INVX1_LOC_6/A NAND2X1_LOC_850/Y 0.07fF
C22365 NOR2X1_LOC_401/B INVX1_LOC_286/A 0.01fF
C22366 INVX1_LOC_226/Y NOR2X1_LOC_394/a_36_216# 0.01fF
C22367 INVX1_LOC_270/A INVX1_LOC_4/A 0.03fF
C22368 NOR2X1_LOC_74/Y INVX1_LOC_22/A 0.13fF
C22369 NOR2X1_LOC_716/B NOR2X1_LOC_35/Y 0.03fF
C22370 INVX1_LOC_180/A VDD 0.12fF
C22371 NOR2X1_LOC_402/a_36_216# INVX1_LOC_286/A 0.01fF
C22372 NOR2X1_LOC_52/B NAND2X1_LOC_843/a_36_24# 0.00fF
C22373 NOR2X1_LOC_753/Y VDD 0.29fF
C22374 INVX1_LOC_93/A INVX1_LOC_29/A 0.08fF
C22375 INVX1_LOC_135/A NOR2X1_LOC_329/B 0.10fF
C22376 NOR2X1_LOC_590/A INVX1_LOC_92/A 0.03fF
C22377 NOR2X1_LOC_561/Y NOR2X1_LOC_313/a_36_216# 0.01fF
C22378 INVX1_LOC_206/Y NOR2X1_LOC_500/Y 0.01fF
C22379 NAND2X1_LOC_833/Y NOR2X1_LOC_305/Y 0.02fF
C22380 NOR2X1_LOC_419/Y NOR2X1_LOC_133/a_36_216# 0.01fF
C22381 NOR2X1_LOC_520/B VDD 0.02fF
C22382 NAND2X1_LOC_20/B INVX1_LOC_3/A 0.01fF
C22383 NAND2X1_LOC_325/Y VDD 0.03fF
C22384 NOR2X1_LOC_304/Y NOR2X1_LOC_48/B 0.04fF
C22385 NAND2X1_LOC_656/A INVX1_LOC_280/A 0.10fF
C22386 NOR2X1_LOC_309/Y INVX1_LOC_20/A 0.07fF
C22387 INVX1_LOC_75/A NOR2X1_LOC_71/Y 0.07fF
C22388 INVX1_LOC_295/A D_INPUT_4 0.04fF
C22389 INVX1_LOC_158/A INVX1_LOC_176/A 0.01fF
C22390 INVX1_LOC_2/A NAND2X1_LOC_447/Y 0.03fF
C22391 NOR2X1_LOC_668/Y NOR2X1_LOC_720/A 0.09fF
C22392 NOR2X1_LOC_239/a_36_216# INVX1_LOC_46/Y 0.00fF
C22393 NOR2X1_LOC_644/A NOR2X1_LOC_439/B 0.00fF
C22394 NOR2X1_LOC_794/A INVX1_LOC_220/Y 0.25fF
C22395 NOR2X1_LOC_201/A NAND2X1_LOC_65/a_36_24# 0.02fF
C22396 NOR2X1_LOC_533/Y INVX1_LOC_264/A 0.23fF
C22397 INVX1_LOC_136/A NAND2X1_LOC_243/B 0.05fF
C22398 INVX1_LOC_90/A NAND2X1_LOC_693/a_36_24# 0.00fF
C22399 NAND2X1_LOC_866/B INVX1_LOC_282/A 0.07fF
C22400 NOR2X1_LOC_644/A INVX1_LOC_75/A 0.03fF
C22401 INVX1_LOC_287/A NOR2X1_LOC_383/B 0.00fF
C22402 NOR2X1_LOC_678/a_36_216# INVX1_LOC_290/Y 0.00fF
C22403 INVX1_LOC_133/Y VDD 0.37fF
C22404 INVX1_LOC_303/A NOR2X1_LOC_489/A 0.04fF
C22405 NAND2X1_LOC_342/Y INVX1_LOC_46/A 0.02fF
C22406 INVX1_LOC_120/A NAND2X1_LOC_111/a_36_24# 0.00fF
C22407 INVX1_LOC_276/A VDD 0.12fF
C22408 INVX1_LOC_35/A NOR2X1_LOC_449/A 0.03fF
C22409 NOR2X1_LOC_669/Y NOR2X1_LOC_48/B 0.46fF
C22410 INVX1_LOC_70/Y NAND2X1_LOC_392/Y 0.11fF
C22411 NOR2X1_LOC_392/Y INVX1_LOC_16/Y 0.36fF
C22412 NOR2X1_LOC_828/B INVX1_LOC_75/A 0.00fF
C22413 NOR2X1_LOC_382/Y INVX1_LOC_84/A 0.08fF
C22414 INVX1_LOC_89/A INVX1_LOC_286/A 0.07fF
C22415 INVX1_LOC_276/A NAND2X1_LOC_800/A 0.15fF
C22416 NOR2X1_LOC_67/A VDD 2.13fF
C22417 INVX1_LOC_240/A NOR2X1_LOC_692/Y 0.11fF
C22418 INVX1_LOC_61/Y NOR2X1_LOC_84/B -0.03fF
C22419 D_INPUT_0 NOR2X1_LOC_78/A 0.07fF
C22420 NOR2X1_LOC_667/A NAND2X1_LOC_721/A 0.35fF
C22421 INVX1_LOC_11/A INVX1_LOC_290/Y 0.04fF
C22422 NAND2X1_LOC_634/Y NAND2X1_LOC_477/Y 0.02fF
C22423 INVX1_LOC_5/A INVX1_LOC_26/A 0.14fF
C22424 INVX1_LOC_23/A NOR2X1_LOC_629/A 0.00fF
C22425 INVX1_LOC_278/Y NAND2X1_LOC_804/Y 0.07fF
C22426 INVX1_LOC_64/A INVX1_LOC_270/A 0.01fF
C22427 NOR2X1_LOC_392/Y NAND2X1_LOC_205/A 0.00fF
C22428 INPUT_6 INVX1_LOC_23/A 0.01fF
C22429 NOR2X1_LOC_742/A INVX1_LOC_311/A 0.05fF
C22430 INVX1_LOC_58/A NOR2X1_LOC_678/A 0.03fF
C22431 INVX1_LOC_103/A INVX1_LOC_32/A 0.12fF
C22432 INVX1_LOC_206/Y NOR2X1_LOC_302/Y 0.21fF
C22433 INVX1_LOC_21/A INVX1_LOC_175/A 0.03fF
C22434 INVX1_LOC_119/A INVX1_LOC_54/A 0.03fF
C22435 NOR2X1_LOC_510/Y NAND2X1_LOC_61/Y 0.01fF
C22436 INVX1_LOC_222/Y NOR2X1_LOC_541/B 0.09fF
C22437 NAND2X1_LOC_354/B INVX1_LOC_92/A 0.49fF
C22438 NOR2X1_LOC_220/A INVX1_LOC_44/A 0.10fF
C22439 INVX1_LOC_39/A INVX1_LOC_23/Y 0.07fF
C22440 INVX1_LOC_52/A INVX1_LOC_281/A 0.02fF
C22441 NAND2X1_LOC_624/B INVX1_LOC_23/A 0.03fF
C22442 NOR2X1_LOC_201/A NOR2X1_LOC_849/A 0.02fF
C22443 NAND2X1_LOC_466/Y NAND2X1_LOC_798/B 0.05fF
C22444 INVX1_LOC_184/A NOR2X1_LOC_814/A 0.04fF
C22445 NOR2X1_LOC_717/B NOR2X1_LOC_35/Y 0.05fF
C22446 NOR2X1_LOC_598/B NOR2X1_LOC_634/Y 0.04fF
C22447 INVX1_LOC_8/A NOR2X1_LOC_216/B 0.07fF
C22448 INVX1_LOC_72/A NAND2X1_LOC_74/B 0.06fF
C22449 INVX1_LOC_88/A NOR2X1_LOC_334/Y 0.22fF
C22450 NAND2X1_LOC_711/Y NOR2X1_LOC_48/B 0.00fF
C22451 NOR2X1_LOC_188/A NOR2X1_LOC_548/B 0.14fF
C22452 INVX1_LOC_104/A INVX1_LOC_307/A 0.07fF
C22453 INVX1_LOC_269/A NAND2X1_LOC_72/B 0.01fF
C22454 INVX1_LOC_14/A NAND2X1_LOC_443/a_36_24# 0.00fF
C22455 INVX1_LOC_13/Y NAND2X1_LOC_464/B 0.50fF
C22456 INVX1_LOC_292/A INVX1_LOC_32/A 0.07fF
C22457 INVX1_LOC_136/A INVX1_LOC_284/A 0.18fF
C22458 INVX1_LOC_104/A NOR2X1_LOC_445/B 0.07fF
C22459 NAND2X1_LOC_660/Y NOR2X1_LOC_60/Y 0.11fF
C22460 INVX1_LOC_110/Y INVX1_LOC_15/A 0.17fF
C22461 D_INPUT_1 NOR2X1_LOC_791/Y 0.03fF
C22462 INVX1_LOC_310/A NOR2X1_LOC_862/B 0.10fF
C22463 NOR2X1_LOC_660/Y NOR2X1_LOC_663/A 0.00fF
C22464 INVX1_LOC_182/A NOR2X1_LOC_486/Y 0.01fF
C22465 INVX1_LOC_174/A NAND2X1_LOC_452/Y 0.02fF
C22466 NOR2X1_LOC_243/Y NOR2X1_LOC_243/B -0.01fF
C22467 NOR2X1_LOC_78/B NOR2X1_LOC_364/A 1.33fF
C22468 NOR2X1_LOC_561/Y NOR2X1_LOC_536/A 0.33fF
C22469 NOR2X1_LOC_303/Y INVX1_LOC_29/A 0.01fF
C22470 NOR2X1_LOC_360/Y INVX1_LOC_42/A 0.11fF
C22471 INVX1_LOC_7/A NOR2X1_LOC_536/A 0.05fF
C22472 NAND2X1_LOC_361/Y INVX1_LOC_19/A 0.14fF
C22473 NOR2X1_LOC_74/A NAND2X1_LOC_642/Y 0.07fF
C22474 INVX1_LOC_25/Y NAND2X1_LOC_243/Y 0.06fF
C22475 NAND2X1_LOC_19/a_36_24# NAND2X1_LOC_223/B 0.00fF
C22476 NOR2X1_LOC_516/B NOR2X1_LOC_640/Y 0.10fF
C22477 NOR2X1_LOC_810/A INVX1_LOC_9/A 0.03fF
C22478 INVX1_LOC_25/Y INVX1_LOC_89/Y 0.10fF
C22479 INVX1_LOC_36/A INVX1_LOC_4/A 0.62fF
C22480 INVX1_LOC_83/A NOR2X1_LOC_862/a_36_216# 0.02fF
C22481 NOR2X1_LOC_507/B INVX1_LOC_122/A 0.00fF
C22482 NOR2X1_LOC_598/B NAND2X1_LOC_473/A 2.12fF
C22483 INVX1_LOC_263/A INVX1_LOC_307/A 0.35fF
C22484 NOR2X1_LOC_15/Y INVX1_LOC_29/Y 0.36fF
C22485 INVX1_LOC_77/A NOR2X1_LOC_89/A 0.19fF
C22486 NOR2X1_LOC_151/Y NOR2X1_LOC_35/Y 0.03fF
C22487 NAND2X1_LOC_738/B NOR2X1_LOC_536/Y 0.26fF
C22488 NOR2X1_LOC_9/Y NAND2X1_LOC_642/Y 0.11fF
C22489 INVX1_LOC_22/A INVX1_LOC_179/A 0.24fF
C22490 NOR2X1_LOC_78/B INVX1_LOC_285/A 0.07fF
C22491 NOR2X1_LOC_68/A NOR2X1_LOC_687/a_36_216# 0.00fF
C22492 NOR2X1_LOC_254/Y INVX1_LOC_29/A 0.01fF
C22493 INVX1_LOC_7/A NOR2X1_LOC_655/Y 0.01fF
C22494 NOR2X1_LOC_433/A INVX1_LOC_290/Y 0.27fF
C22495 NOR2X1_LOC_791/Y NOR2X1_LOC_652/Y 0.00fF
C22496 INVX1_LOC_150/A INVX1_LOC_54/A 0.02fF
C22497 NOR2X1_LOC_547/B NOR2X1_LOC_814/A 0.08fF
C22498 INVX1_LOC_50/A INVX1_LOC_225/Y 2.01fF
C22499 NOR2X1_LOC_593/Y INVX1_LOC_290/Y 0.08fF
C22500 D_INPUT_1 NOR2X1_LOC_457/A 0.11fF
C22501 NAND2X1_LOC_338/B INVX1_LOC_293/Y 0.02fF
C22502 NOR2X1_LOC_329/B NOR2X1_LOC_152/A 0.03fF
C22503 INVX1_LOC_227/A INVX1_LOC_92/A 0.07fF
C22504 INVX1_LOC_31/A NOR2X1_LOC_720/A 0.01fF
C22505 NAND2X1_LOC_114/B INVX1_LOC_57/A 0.89fF
C22506 NOR2X1_LOC_152/Y D_INPUT_5 0.53fF
C22507 INVX1_LOC_104/A INVX1_LOC_12/A 0.07fF
C22508 NOR2X1_LOC_208/Y INVX1_LOC_4/A 0.03fF
C22509 INVX1_LOC_89/A INVX1_LOC_54/A 0.09fF
C22510 INVX1_LOC_311/A INVX1_LOC_139/A 0.01fF
C22511 INVX1_LOC_133/Y INVX1_LOC_133/A 0.03fF
C22512 NOR2X1_LOC_848/Y INVX1_LOC_35/A 0.15fF
C22513 NAND2X1_LOC_725/A NAND2X1_LOC_537/Y 0.10fF
C22514 NOR2X1_LOC_457/B INVX1_LOC_271/Y 0.05fF
C22515 NOR2X1_LOC_763/Y INVX1_LOC_92/A 0.65fF
C22516 NAND2X1_LOC_803/B INVX1_LOC_53/A 0.02fF
C22517 INVX1_LOC_72/A NOR2X1_LOC_45/a_36_216# 0.00fF
C22518 INVX1_LOC_54/Y INVX1_LOC_29/A 0.10fF
C22519 INVX1_LOC_16/A NOR2X1_LOC_666/a_36_216# 0.00fF
C22520 INVX1_LOC_124/A NOR2X1_LOC_89/A 0.02fF
C22521 INVX1_LOC_141/Y INVX1_LOC_57/A 0.03fF
C22522 NOR2X1_LOC_551/Y VDD 0.14fF
C22523 INVX1_LOC_36/A NAND2X1_LOC_420/a_36_24# 0.00fF
C22524 NOR2X1_LOC_537/Y NAND2X1_LOC_74/B 0.46fF
C22525 NAND2X1_LOC_859/a_36_24# INVX1_LOC_284/A 0.01fF
C22526 NAND2X1_LOC_338/B NAND2X1_LOC_74/B 0.21fF
C22527 NOR2X1_LOC_160/B NOR2X1_LOC_247/Y 0.15fF
C22528 NOR2X1_LOC_537/Y NAND2X1_LOC_207/Y 0.01fF
C22529 NOR2X1_LOC_514/A INVX1_LOC_23/A 0.78fF
C22530 INVX1_LOC_288/Y INVX1_LOC_72/A 0.03fF
C22531 NAND2X1_LOC_860/A NOR2X1_LOC_372/A 0.38fF
C22532 INVX1_LOC_61/A INVX1_LOC_23/Y 0.01fF
C22533 INVX1_LOC_119/A NOR2X1_LOC_48/B 0.43fF
C22534 NOR2X1_LOC_92/Y NAND2X1_LOC_474/Y 0.07fF
C22535 NOR2X1_LOC_590/A INVX1_LOC_53/A 0.15fF
C22536 NAND2X1_LOC_548/a_36_24# INVX1_LOC_29/A 0.00fF
C22537 INVX1_LOC_2/A NOR2X1_LOC_46/a_36_216# 0.01fF
C22538 INVX1_LOC_98/A NOR2X1_LOC_266/B 0.18fF
C22539 NOR2X1_LOC_589/A INVX1_LOC_63/A 5.65fF
C22540 INVX1_LOC_7/A NOR2X1_LOC_649/B 0.06fF
C22541 NOR2X1_LOC_65/B NOR2X1_LOC_360/Y 0.10fF
C22542 D_INPUT_1 INVX1_LOC_30/A 0.03fF
C22543 INVX1_LOC_18/A NOR2X1_LOC_383/B 0.17fF
C22544 INVX1_LOC_85/Y NOR2X1_LOC_155/A 0.03fF
C22545 INVX1_LOC_7/A INVX1_LOC_3/A 0.18fF
C22546 INVX1_LOC_248/A NOR2X1_LOC_669/A 0.01fF
C22547 NOR2X1_LOC_78/A NOR2X1_LOC_266/B 0.04fF
C22548 INVX1_LOC_232/A NAND2X1_LOC_63/Y 0.05fF
C22549 NOR2X1_LOC_91/A INVX1_LOC_41/Y 0.13fF
C22550 NOR2X1_LOC_309/Y INVX1_LOC_4/A 0.08fF
C22551 INVX1_LOC_83/A NOR2X1_LOC_814/A 0.15fF
C22552 NAND2X1_LOC_136/a_36_24# NOR2X1_LOC_660/Y 0.00fF
C22553 NAND2X1_LOC_862/Y INVX1_LOC_119/Y 0.04fF
C22554 INVX1_LOC_69/Y INVX1_LOC_9/A 0.07fF
C22555 INVX1_LOC_64/A INVX1_LOC_36/A 0.10fF
C22556 NOR2X1_LOC_454/Y INVX1_LOC_11/A 0.19fF
C22557 INVX1_LOC_272/Y NOR2X1_LOC_92/Y 0.10fF
C22558 NOR2X1_LOC_274/B NOR2X1_LOC_405/Y 0.04fF
C22559 INVX1_LOC_135/A NOR2X1_LOC_691/B 0.29fF
C22560 INVX1_LOC_171/A INVX1_LOC_63/A 0.02fF
C22561 NAND2X1_LOC_361/Y INVX1_LOC_26/Y 0.08fF
C22562 INVX1_LOC_31/A NOR2X1_LOC_849/A 0.03fF
C22563 NOR2X1_LOC_84/Y NOR2X1_LOC_394/Y 0.05fF
C22564 INVX1_LOC_187/A INVX1_LOC_77/Y 0.02fF
C22565 NAND2X1_LOC_214/B NOR2X1_LOC_414/a_36_216# 0.02fF
C22566 NOR2X1_LOC_242/A NOR2X1_LOC_590/A 0.06fF
C22567 NAND2X1_LOC_9/Y NOR2X1_LOC_791/a_36_216# 0.00fF
C22568 INVX1_LOC_240/A NAND2X1_LOC_175/Y 0.02fF
C22569 NOR2X1_LOC_182/a_36_216# INVX1_LOC_271/Y 0.01fF
C22570 NOR2X1_LOC_617/Y INVX1_LOC_23/A 0.02fF
C22571 INVX1_LOC_256/A NAND2X1_LOC_67/Y 0.07fF
C22572 NOR2X1_LOC_336/B INVX1_LOC_50/Y 0.05fF
C22573 NOR2X1_LOC_456/Y INVX1_LOC_71/A 0.07fF
C22574 NAND2X1_LOC_593/Y INVX1_LOC_23/A 0.01fF
C22575 INVX1_LOC_30/A NOR2X1_LOC_652/Y 0.02fF
C22576 NAND2X1_LOC_721/A NOR2X1_LOC_670/Y 0.22fF
C22577 INVX1_LOC_14/A NAND2X1_LOC_793/Y 2.26fF
C22578 INVX1_LOC_21/A NAND2X1_LOC_36/A 0.01fF
C22579 NOR2X1_LOC_272/Y NOR2X1_LOC_248/Y 0.02fF
C22580 INVX1_LOC_36/A NAND2X1_LOC_27/a_36_24# 0.00fF
C22581 NOR2X1_LOC_203/Y NOR2X1_LOC_334/Y 0.03fF
C22582 NAND2X1_LOC_357/B NOR2X1_LOC_282/Y 0.03fF
C22583 NAND2X1_LOC_451/Y INVX1_LOC_78/A 0.10fF
C22584 INVX1_LOC_64/A INVX1_LOC_145/A 0.23fF
C22585 NAND2X1_LOC_361/Y NAND2X1_LOC_265/a_36_24# 0.01fF
C22586 INVX1_LOC_206/Y INVX1_LOC_307/A 0.18fF
C22587 INVX1_LOC_50/A NAND2X1_LOC_811/Y 0.04fF
C22588 NAND2X1_LOC_364/A INVX1_LOC_50/Y 0.10fF
C22589 NOR2X1_LOC_811/A NOR2X1_LOC_812/A 0.00fF
C22590 NOR2X1_LOC_91/Y INVX1_LOC_306/Y 0.27fF
C22591 NOR2X1_LOC_279/a_36_216# NOR2X1_LOC_301/A 0.00fF
C22592 INVX1_LOC_251/Y NAND2X1_LOC_99/A 0.01fF
C22593 NOR2X1_LOC_536/A INVX1_LOC_76/A 0.30fF
C22594 INVX1_LOC_277/A INVX1_LOC_1/A 0.03fF
C22595 INVX1_LOC_21/A NAND2X1_LOC_514/Y 0.01fF
C22596 NAND2X1_LOC_740/Y NAND2X1_LOC_731/Y 0.00fF
C22597 INVX1_LOC_140/A NOR2X1_LOC_36/B 0.05fF
C22598 INVX1_LOC_114/A NAND2X1_LOC_220/a_36_24# 0.00fF
C22599 NAND2X1_LOC_354/B INVX1_LOC_53/A 0.07fF
C22600 INVX1_LOC_50/A INVX1_LOC_266/Y 0.03fF
C22601 NOR2X1_LOC_598/B NOR2X1_LOC_486/B 0.21fF
C22602 NOR2X1_LOC_78/A INVX1_LOC_46/Y 0.21fF
C22603 INVX1_LOC_64/A NOR2X1_LOC_804/B 0.07fF
C22604 NOR2X1_LOC_773/Y INVX1_LOC_26/A 0.02fF
C22605 NOR2X1_LOC_600/Y INVX1_LOC_307/A 0.21fF
C22606 INVX1_LOC_11/A NAND2X1_LOC_387/a_36_24# 0.00fF
C22607 NOR2X1_LOC_168/B INVX1_LOC_57/A 0.14fF
C22608 NOR2X1_LOC_167/Y NOR2X1_LOC_661/A 0.02fF
C22609 NOR2X1_LOC_536/A NAND2X1_LOC_84/a_36_24# 0.00fF
C22610 NAND2X1_LOC_560/A NOR2X1_LOC_824/a_36_216# 0.00fF
C22611 NAND2X1_LOC_866/B NOR2X1_LOC_496/a_36_216# 0.00fF
C22612 NOR2X1_LOC_561/Y NAND2X1_LOC_470/B 0.20fF
C22613 VDD NOR2X1_LOC_729/A 0.37fF
C22614 NOR2X1_LOC_649/a_36_216# NOR2X1_LOC_649/Y 0.01fF
C22615 INVX1_LOC_5/A INVX1_LOC_315/A 0.10fF
C22616 NAND2X1_LOC_93/B INVX1_LOC_76/A 0.07fF
C22617 INVX1_LOC_89/A NAND2X1_LOC_3/B 0.00fF
C22618 NAND2X1_LOC_725/B INVX1_LOC_24/A 0.11fF
C22619 NOR2X1_LOC_406/a_36_216# NAND2X1_LOC_357/B 0.00fF
C22620 INVX1_LOC_31/A NOR2X1_LOC_514/A 0.02fF
C22621 NOR2X1_LOC_454/Y NOR2X1_LOC_433/A 0.03fF
C22622 NOR2X1_LOC_425/Y INVX1_LOC_54/A 0.01fF
C22623 INVX1_LOC_36/A INVX1_LOC_43/Y 0.13fF
C22624 NAND2X1_LOC_385/a_36_24# INVX1_LOC_54/Y 0.00fF
C22625 INVX1_LOC_91/A NOR2X1_LOC_257/Y 0.00fF
C22626 INVX1_LOC_41/A NAND2X1_LOC_474/Y 0.02fF
C22627 NAND2X1_LOC_425/Y INVX1_LOC_76/A 0.01fF
C22628 INVX1_LOC_21/A NAND2X1_LOC_332/Y 0.02fF
C22629 NAND2X1_LOC_549/Y NAND2X1_LOC_549/B 0.12fF
C22630 NOR2X1_LOC_276/Y INVX1_LOC_72/A 0.00fF
C22631 NOR2X1_LOC_807/B NOR2X1_LOC_324/Y 0.01fF
C22632 NAND2X1_LOC_803/B NAND2X1_LOC_156/a_36_24# 0.01fF
C22633 INVX1_LOC_290/A NOR2X1_LOC_654/A 0.01fF
C22634 NAND2X1_LOC_363/B NOR2X1_LOC_620/B 0.05fF
C22635 NOR2X1_LOC_375/Y NOR2X1_LOC_476/B 0.00fF
C22636 INVX1_LOC_76/Y NOR2X1_LOC_460/Y 0.14fF
C22637 NOR2X1_LOC_180/B INVX1_LOC_271/Y 0.04fF
C22638 NAND2X1_LOC_13/a_36_24# INVX1_LOC_314/Y 0.00fF
C22639 INVX1_LOC_224/A INVX1_LOC_77/A 0.03fF
C22640 NAND2X1_LOC_358/B NAND2X1_LOC_323/B 0.07fF
C22641 NAND2X1_LOC_850/Y NOR2X1_LOC_109/Y 0.07fF
C22642 INVX1_LOC_61/Y INVX1_LOC_72/Y 0.14fF
C22643 INVX1_LOC_11/A INVX1_LOC_77/A 1.68fF
C22644 NOR2X1_LOC_510/Y INVX1_LOC_133/Y 0.41fF
C22645 INVX1_LOC_1/A NOR2X1_LOC_285/B 0.02fF
C22646 NOR2X1_LOC_817/Y NOR2X1_LOC_554/a_36_216# 0.00fF
C22647 INVX1_LOC_76/A INVX1_LOC_3/A 0.91fF
C22648 NAND2X1_LOC_96/A NOR2X1_LOC_862/B 0.10fF
C22649 INVX1_LOC_276/A NOR2X1_LOC_510/Y 0.02fF
C22650 NOR2X1_LOC_454/Y NOR2X1_LOC_52/B 0.04fF
C22651 NAND2X1_LOC_656/Y INVX1_LOC_57/A 0.00fF
C22652 NAND2X1_LOC_796/B INVX1_LOC_2/A 0.13fF
C22653 INVX1_LOC_46/A INVX1_LOC_285/A 0.15fF
C22654 INVX1_LOC_20/A INVX1_LOC_63/A 0.10fF
C22655 NAND2X1_LOC_363/Y NOR2X1_LOC_836/A 0.83fF
C22656 INVX1_LOC_31/A INVX1_LOC_41/Y 0.03fF
C22657 NOR2X1_LOC_666/Y INVX1_LOC_88/Y 0.31fF
C22658 INVX1_LOC_57/Y INVX1_LOC_18/A 0.07fF
C22659 INVX1_LOC_136/A INVX1_LOC_72/A 0.30fF
C22660 NOR2X1_LOC_590/A INVX1_LOC_184/A 0.01fF
C22661 NOR2X1_LOC_15/Y INVX1_LOC_60/Y 0.03fF
C22662 NOR2X1_LOC_357/Y NOR2X1_LOC_631/A 0.01fF
C22663 INVX1_LOC_36/A INVX1_LOC_130/Y 0.03fF
C22664 INVX1_LOC_41/A NAND2X1_LOC_53/Y 0.36fF
C22665 INVX1_LOC_46/A NOR2X1_LOC_814/A 0.07fF
C22666 INVX1_LOC_227/A INVX1_LOC_53/A 0.09fF
C22667 INVX1_LOC_1/A NOR2X1_LOC_300/Y 0.00fF
C22668 INVX1_LOC_132/Y INVX1_LOC_57/A 0.03fF
C22669 INVX1_LOC_89/A NAND2X1_LOC_215/A 0.07fF
C22670 INVX1_LOC_243/Y NAND2X1_LOC_638/Y 0.31fF
C22671 NAND2X1_LOC_447/Y NAND2X1_LOC_63/Y 0.01fF
C22672 NOR2X1_LOC_763/Y INVX1_LOC_53/A 0.02fF
C22673 INVX1_LOC_31/A NAND2X1_LOC_593/Y 0.46fF
C22674 INVX1_LOC_45/A NOR2X1_LOC_274/a_36_216# 0.01fF
C22675 INVX1_LOC_144/A NAND2X1_LOC_454/Y 0.06fF
C22676 NOR2X1_LOC_793/Y INVX1_LOC_177/A 0.00fF
C22677 NOR2X1_LOC_274/a_36_216# NOR2X1_LOC_568/A 0.01fF
C22678 INVX1_LOC_18/A NOR2X1_LOC_512/Y 0.00fF
C22679 INVX1_LOC_2/A NOR2X1_LOC_232/a_36_216# 0.00fF
C22680 INVX1_LOC_39/A INVX1_LOC_232/A 0.01fF
C22681 D_GATE_366 INVX1_LOC_105/Y 0.02fF
C22682 NOR2X1_LOC_361/B INVX1_LOC_133/Y 1.14fF
C22683 INVX1_LOC_100/A INVX1_LOC_165/A 0.02fF
C22684 NAND2X1_LOC_582/a_36_24# NAND2X1_LOC_30/Y 0.00fF
C22685 INVX1_LOC_35/A INVX1_LOC_135/A 0.33fF
C22686 NOR2X1_LOC_134/Y NAND2X1_LOC_139/A 0.09fF
C22687 INVX1_LOC_124/A INVX1_LOC_11/A 0.03fF
C22688 INVX1_LOC_182/A NOR2X1_LOC_748/A 0.10fF
C22689 NOR2X1_LOC_598/B INVX1_LOC_85/Y 0.11fF
C22690 NOR2X1_LOC_67/A NOR2X1_LOC_361/B 0.10fF
C22691 NOR2X1_LOC_32/B INVX1_LOC_90/A 0.02fF
C22692 NAND2X1_LOC_53/Y NOR2X1_LOC_207/A 0.01fF
C22693 INVX1_LOC_119/A NAND2X1_LOC_350/A 0.09fF
C22694 NOR2X1_LOC_384/Y NOR2X1_LOC_625/Y 0.01fF
C22695 NOR2X1_LOC_208/Y INVX1_LOC_130/Y 0.37fF
C22696 INVX1_LOC_28/A NOR2X1_LOC_591/A 0.06fF
C22697 NOR2X1_LOC_191/B INVX1_LOC_181/Y 0.01fF
C22698 NOR2X1_LOC_639/B INVX1_LOC_90/A 0.01fF
C22699 NOR2X1_LOC_289/Y INVX1_LOC_271/A 0.10fF
C22700 INVX1_LOC_24/A INVX1_LOC_309/Y 0.01fF
C22701 INVX1_LOC_18/A NAND2X1_LOC_632/B 0.13fF
C22702 NOR2X1_LOC_158/B INVX1_LOC_91/A 0.00fF
C22703 NOR2X1_LOC_273/Y INVX1_LOC_71/A 0.03fF
C22704 INVX1_LOC_50/A INVX1_LOC_42/Y 0.00fF
C22705 VDD NOR2X1_LOC_584/Y 0.08fF
C22706 NAND2X1_LOC_624/B NAND2X1_LOC_866/B 0.05fF
C22707 NOR2X1_LOC_328/Y NAND2X1_LOC_303/Y 0.10fF
C22708 NOR2X1_LOC_703/A INVX1_LOC_53/A 0.03fF
C22709 NOR2X1_LOC_790/B NOR2X1_LOC_564/Y 0.03fF
C22710 INVX1_LOC_33/Y NOR2X1_LOC_831/Y 0.25fF
C22711 NOR2X1_LOC_186/Y D_INPUT_0 0.07fF
C22712 NOR2X1_LOC_759/Y INVX1_LOC_71/A 0.94fF
C22713 NOR2X1_LOC_634/A NAND2X1_LOC_412/a_36_24# 0.02fF
C22714 INVX1_LOC_269/A INVX1_LOC_53/Y 0.07fF
C22715 NAND2X1_LOC_727/Y NAND2X1_LOC_724/A 0.01fF
C22716 NOR2X1_LOC_269/Y INVX1_LOC_78/A 1.75fF
C22717 INVX1_LOC_202/A INVX1_LOC_71/A 0.07fF
C22718 INVX1_LOC_256/A NOR2X1_LOC_131/a_36_216# 0.00fF
C22719 INVX1_LOC_45/Y NOR2X1_LOC_577/Y 0.08fF
C22720 INVX1_LOC_34/A NOR2X1_LOC_791/B 0.04fF
C22721 NAND2X1_LOC_555/Y NAND2X1_LOC_578/B 0.02fF
C22722 NOR2X1_LOC_92/Y INVX1_LOC_10/A 0.07fF
C22723 NOR2X1_LOC_632/Y NOR2X1_LOC_205/Y 0.00fF
C22724 NOR2X1_LOC_590/A NOR2X1_LOC_78/B 0.10fF
C22725 INVX1_LOC_242/Y INVX1_LOC_22/A 0.01fF
C22726 NAND2X1_LOC_573/Y D_INPUT_0 0.07fF
C22727 NAND2X1_LOC_214/B NOR2X1_LOC_750/A 0.01fF
C22728 NOR2X1_LOC_431/Y NOR2X1_LOC_172/Y 0.00fF
C22729 NAND2X1_LOC_364/A NOR2X1_LOC_6/B 0.07fF
C22730 NOR2X1_LOC_433/A INVX1_LOC_77/A 0.10fF
C22731 INVX1_LOC_27/A INVX1_LOC_65/Y 0.01fF
C22732 NOR2X1_LOC_798/A INVX1_LOC_87/Y 0.04fF
C22733 NOR2X1_LOC_45/B NAND2X1_LOC_99/A 0.04fF
C22734 INVX1_LOC_64/A NOR2X1_LOC_19/Y 0.27fF
C22735 NOR2X1_LOC_716/B NOR2X1_LOC_350/A 0.04fF
C22736 NOR2X1_LOC_75/Y INVX1_LOC_290/A 0.07fF
C22737 NOR2X1_LOC_15/Y NOR2X1_LOC_355/A 0.03fF
C22738 NOR2X1_LOC_593/Y INVX1_LOC_77/A 0.05fF
C22739 NOR2X1_LOC_89/A INVX1_LOC_9/A 0.12fF
C22740 NOR2X1_LOC_778/B INVX1_LOC_223/A 0.07fF
C22741 INVX1_LOC_179/A INVX1_LOC_186/Y 2.28fF
C22742 NOR2X1_LOC_769/A NAND2X1_LOC_451/Y 0.09fF
C22743 NAND2X1_LOC_470/B INVX1_LOC_76/A 0.47fF
C22744 NOR2X1_LOC_155/A NAND2X1_LOC_782/B 0.03fF
C22745 NOR2X1_LOC_644/B INVX1_LOC_16/A 0.01fF
C22746 NOR2X1_LOC_127/a_36_216# NOR2X1_LOC_127/Y 0.00fF
C22747 INVX1_LOC_11/A NAND2X1_LOC_796/Y 0.02fF
C22748 INVX1_LOC_36/A NAND2X1_LOC_850/Y 0.15fF
C22749 INVX1_LOC_136/A NAND2X1_LOC_338/B 0.17fF
C22750 INVX1_LOC_256/A NOR2X1_LOC_561/Y 0.18fF
C22751 NOR2X1_LOC_637/B NAND2X1_LOC_175/B 0.02fF
C22752 INVX1_LOC_275/A NAND2X1_LOC_686/a_36_24# 0.01fF
C22753 INVX1_LOC_202/Y INVX1_LOC_15/A 0.01fF
C22754 NOR2X1_LOC_267/A NAND2X1_LOC_850/Y 0.15fF
C22755 NOR2X1_LOC_626/Y NOR2X1_LOC_742/A 0.03fF
C22756 NAND2X1_LOC_213/A NOR2X1_LOC_156/A 0.03fF
C22757 NAND2X1_LOC_803/B INVX1_LOC_83/A 0.02fF
C22758 INVX1_LOC_77/A NOR2X1_LOC_52/B 0.34fF
C22759 INVX1_LOC_147/Y NOR2X1_LOC_65/Y 0.05fF
C22760 INVX1_LOC_35/Y INVX1_LOC_29/A 0.07fF
C22761 INVX1_LOC_105/A INVX1_LOC_266/Y 0.00fF
C22762 NOR2X1_LOC_742/a_36_216# INVX1_LOC_85/Y 0.00fF
C22763 NOR2X1_LOC_392/B INVX1_LOC_155/Y 0.00fF
C22764 NOR2X1_LOC_751/Y INVX1_LOC_22/A 0.02fF
C22765 INVX1_LOC_34/A NOR2X1_LOC_124/B 0.01fF
C22766 NAND2X1_LOC_39/a_36_24# NOR2X1_LOC_589/A 0.00fF
C22767 NOR2X1_LOC_673/B NOR2X1_LOC_721/B 0.01fF
C22768 NOR2X1_LOC_590/A INVX1_LOC_83/A 0.10fF
C22769 INVX1_LOC_233/A INVX1_LOC_70/Y 0.03fF
C22770 NOR2X1_LOC_606/Y INVX1_LOC_7/A 0.02fF
C22771 NOR2X1_LOC_301/A NOR2X1_LOC_653/a_36_216# 0.00fF
C22772 NOR2X1_LOC_716/B NOR2X1_LOC_84/Y 0.58fF
C22773 INVX1_LOC_124/A NOR2X1_LOC_593/Y 0.10fF
C22774 NOR2X1_LOC_152/Y NAND2X1_LOC_451/Y 0.00fF
C22775 INVX1_LOC_13/A NAND2X1_LOC_351/A 0.02fF
C22776 NAND2X1_LOC_741/B INPUT_5 0.01fF
C22777 INVX1_LOC_22/Y INVX1_LOC_83/A 0.03fF
C22778 NAND2X1_LOC_579/A NOR2X1_LOC_323/Y 0.34fF
C22779 INVX1_LOC_218/Y INVX1_LOC_89/A 0.05fF
C22780 NOR2X1_LOC_804/a_36_216# NOR2X1_LOC_551/B 0.00fF
C22781 NOR2X1_LOC_389/A NOR2X1_LOC_473/B 0.10fF
C22782 NAND2X1_LOC_638/a_36_24# NOR2X1_LOC_467/A 0.01fF
C22783 VDD NAND2X1_LOC_787/Y -0.00fF
C22784 NOR2X1_LOC_67/A NOR2X1_LOC_132/Y 0.01fF
C22785 INVX1_LOC_180/Y INVX1_LOC_15/A 0.04fF
C22786 INVX1_LOC_94/A NOR2X1_LOC_570/Y 0.00fF
C22787 INVX1_LOC_124/A NOR2X1_LOC_52/B 0.01fF
C22788 NOR2X1_LOC_817/Y INVX1_LOC_75/A 0.07fF
C22789 NOR2X1_LOC_349/A INVX1_LOC_50/Y 0.80fF
C22790 NOR2X1_LOC_721/B INVX1_LOC_29/A 0.01fF
C22791 NAND2X1_LOC_859/Y INVX1_LOC_41/Y 0.00fF
C22792 INVX1_LOC_33/A INVX1_LOC_43/A 0.00fF
C22793 INVX1_LOC_291/Y NOR2X1_LOC_304/Y 0.06fF
C22794 INVX1_LOC_269/A NOR2X1_LOC_113/B 0.01fF
C22795 INVX1_LOC_172/A NAND2X1_LOC_170/A 0.03fF
C22796 NOR2X1_LOC_820/A NOR2X1_LOC_332/A 0.03fF
C22797 INVX1_LOC_48/Y NOR2X1_LOC_392/a_36_216# 0.01fF
C22798 NOR2X1_LOC_778/B INVX1_LOC_149/Y 0.02fF
C22799 INVX1_LOC_208/Y INVX1_LOC_33/A 0.66fF
C22800 NOR2X1_LOC_309/Y NAND2X1_LOC_850/Y 0.10fF
C22801 INVX1_LOC_41/A INVX1_LOC_226/Y 0.01fF
C22802 INVX1_LOC_136/A INVX1_LOC_313/Y 0.12fF
C22803 NAND2X1_LOC_341/A INVX1_LOC_63/Y 0.02fF
C22804 INVX1_LOC_30/A NOR2X1_LOC_497/Y 0.03fF
C22805 NAND2X1_LOC_659/A INVX1_LOC_32/A 0.95fF
C22806 NOR2X1_LOC_646/A INVX1_LOC_34/A 0.06fF
C22807 NOR2X1_LOC_272/Y NOR2X1_LOC_124/A 0.21fF
C22808 NOR2X1_LOC_455/a_36_216# NOR2X1_LOC_500/Y 0.00fF
C22809 NOR2X1_LOC_607/A NOR2X1_LOC_137/A 0.38fF
C22810 NOR2X1_LOC_266/a_36_216# NAND2X1_LOC_842/B 0.00fF
C22811 NOR2X1_LOC_226/A NAND2X1_LOC_572/a_36_24# 0.01fF
C22812 VDD INVX1_LOC_68/A 0.12fF
C22813 NOR2X1_LOC_155/A NAND2X1_LOC_454/Y 0.52fF
C22814 NAND2X1_LOC_364/Y INVX1_LOC_160/Y 0.12fF
C22815 INVX1_LOC_29/A NOR2X1_LOC_610/Y 0.01fF
C22816 INVX1_LOC_223/A NAND2X1_LOC_123/Y 0.03fF
C22817 NAND2X1_LOC_11/a_36_24# NAND2X1_LOC_11/Y 0.02fF
C22818 NOR2X1_LOC_91/A INVX1_LOC_185/A 0.50fF
C22819 INVX1_LOC_35/A NOR2X1_LOC_813/Y 0.07fF
C22820 NOR2X1_LOC_454/Y INVX1_LOC_199/A 0.14fF
C22821 NOR2X1_LOC_631/A INVX1_LOC_32/A 0.09fF
C22822 INVX1_LOC_130/A INPUT_0 0.03fF
C22823 INVX1_LOC_266/A NOR2X1_LOC_405/A 0.00fF
C22824 INVX1_LOC_50/Y NOR2X1_LOC_857/A 0.10fF
C22825 NAND2X1_LOC_866/B INVX1_LOC_41/Y 0.00fF
C22826 NAND2X1_LOC_36/A NAND2X1_LOC_51/B 1.82fF
C22827 NOR2X1_LOC_373/Y NOR2X1_LOC_373/a_36_216# 0.00fF
C22828 INVX1_LOC_132/A D_INPUT_0 0.07fF
C22829 NOR2X1_LOC_431/Y INVX1_LOC_90/A 0.01fF
C22830 INVX1_LOC_41/A INVX1_LOC_10/A 0.03fF
C22831 NOR2X1_LOC_456/Y NOR2X1_LOC_331/B 0.45fF
C22832 INVX1_LOC_17/A INVX1_LOC_91/A 0.31fF
C22833 INVX1_LOC_21/A INVX1_LOC_176/A 0.58fF
C22834 INVX1_LOC_226/Y NOR2X1_LOC_398/Y 0.01fF
C22835 INVX1_LOC_4/A INVX1_LOC_63/A 0.04fF
C22836 INVX1_LOC_285/A NOR2X1_LOC_282/a_36_216# 0.00fF
C22837 NOR2X1_LOC_32/B INVX1_LOC_38/A 0.12fF
C22838 INVX1_LOC_36/A INVX1_LOC_282/A 0.07fF
C22839 NOR2X1_LOC_498/Y INVX1_LOC_10/A 0.06fF
C22840 INVX1_LOC_18/A NOR2X1_LOC_163/Y 0.01fF
C22841 NOR2X1_LOC_464/B INVX1_LOC_247/A 0.01fF
C22842 INVX1_LOC_35/A INVX1_LOC_280/A 0.14fF
C22843 NOR2X1_LOC_639/B INVX1_LOC_38/A 0.02fF
C22844 NOR2X1_LOC_65/B NOR2X1_LOC_79/Y 0.03fF
C22845 NOR2X1_LOC_142/Y INVX1_LOC_150/A 0.01fF
C22846 INVX1_LOC_64/A NOR2X1_LOC_865/A 0.02fF
C22847 NOR2X1_LOC_32/B NOR2X1_LOC_96/Y 0.56fF
C22848 NOR2X1_LOC_332/A INVX1_LOC_315/A 0.02fF
C22849 INVX1_LOC_2/A NAND2X1_LOC_112/Y 0.04fF
C22850 INVX1_LOC_299/A NAND2X1_LOC_280/a_36_24# 0.00fF
C22851 NOR2X1_LOC_15/Y INVX1_LOC_126/A 0.49fF
C22852 NAND2X1_LOC_357/A INVX1_LOC_95/A 0.45fF
C22853 INVX1_LOC_18/A NOR2X1_LOC_74/Y 0.02fF
C22854 INVX1_LOC_282/Y NAND2X1_LOC_866/a_36_24# 0.07fF
C22855 INVX1_LOC_89/A NOR2X1_LOC_340/Y 0.20fF
C22856 INVX1_LOC_225/A D_INPUT_0 0.03fF
C22857 NAND2X1_LOC_477/A INVX1_LOC_10/A 0.00fF
C22858 NOR2X1_LOC_82/A INVX1_LOC_304/A 0.07fF
C22859 NOR2X1_LOC_791/B INPUT_0 0.03fF
C22860 NOR2X1_LOC_68/A INVX1_LOC_144/A 0.07fF
C22861 NOR2X1_LOC_470/B INVX1_LOC_115/A 0.08fF
C22862 NOR2X1_LOC_169/B INVX1_LOC_69/Y 0.03fF
C22863 NOR2X1_LOC_328/Y NOR2X1_LOC_226/a_36_216# 0.00fF
C22864 NOR2X1_LOC_288/A D_INPUT_0 0.03fF
C22865 NOR2X1_LOC_91/Y NOR2X1_LOC_74/A 0.24fF
C22866 NAND2X1_LOC_214/Y VDD 0.00fF
C22867 NAND2X1_LOC_788/a_36_24# INVX1_LOC_33/Y 0.00fF
C22868 NOR2X1_LOC_186/Y NAND2X1_LOC_848/A 0.10fF
C22869 NOR2X1_LOC_590/A NOR2X1_LOC_311/Y 0.03fF
C22870 NAND2X1_LOC_139/A INPUT_1 0.04fF
C22871 NOR2X1_LOC_738/a_36_216# NOR2X1_LOC_687/Y 0.02fF
C22872 NOR2X1_LOC_334/Y INVX1_LOC_272/A 0.01fF
C22873 INVX1_LOC_225/A NOR2X1_LOC_389/a_36_216# 0.01fF
C22874 NOR2X1_LOC_720/B INVX1_LOC_90/A 0.01fF
C22875 NOR2X1_LOC_32/B NAND2X1_LOC_848/Y 0.03fF
C22876 INVX1_LOC_25/A NAND2X1_LOC_572/B 0.07fF
C22877 INVX1_LOC_256/A INVX1_LOC_76/A 0.20fF
C22878 NOR2X1_LOC_634/A NOR2X1_LOC_634/Y 0.08fF
C22879 NOR2X1_LOC_286/Y VDD 0.10fF
C22880 INVX1_LOC_124/Y NAND2X1_LOC_642/Y 0.05fF
C22881 NOR2X1_LOC_178/Y NAND2X1_LOC_93/B 0.45fF
C22882 NAND2X1_LOC_573/Y NAND2X1_LOC_848/A 0.10fF
C22883 NOR2X1_LOC_644/A NOR2X1_LOC_348/B 0.34fF
C22884 NOR2X1_LOC_255/a_36_216# INVX1_LOC_25/Y 0.02fF
C22885 NOR2X1_LOC_84/Y NOR2X1_LOC_130/Y 0.03fF
C22886 NOR2X1_LOC_757/A INVX1_LOC_208/A 0.01fF
C22887 NAND2X1_LOC_572/a_36_24# INPUT_1 0.00fF
C22888 INVX1_LOC_215/A NAND2X1_LOC_349/B 0.02fF
C22889 INVX1_LOC_88/A NAND2X1_LOC_472/Y 0.14fF
C22890 NOR2X1_LOC_433/A NAND2X1_LOC_832/Y 0.01fF
C22891 INVX1_LOC_224/Y INVX1_LOC_293/Y 0.19fF
C22892 NOR2X1_LOC_655/B INVX1_LOC_89/A 0.38fF
C22893 NOR2X1_LOC_134/Y NAND2X1_LOC_464/A 0.00fF
C22894 NOR2X1_LOC_391/A INVX1_LOC_16/A 0.03fF
C22895 NAND2X1_LOC_563/a_36_24# D_INPUT_3 0.01fF
C22896 NAND2X1_LOC_320/a_36_24# NOR2X1_LOC_356/A 0.00fF
C22897 NAND2X1_LOC_550/A INVX1_LOC_37/A 0.07fF
C22898 INVX1_LOC_135/A INVX1_LOC_84/Y 0.02fF
C22899 NOR2X1_LOC_596/A NOR2X1_LOC_355/B 0.05fF
C22900 NOR2X1_LOC_373/Y INVX1_LOC_25/Y 0.01fF
C22901 NAND2X1_LOC_286/B INVX1_LOC_29/A 0.09fF
C22902 NAND2X1_LOC_833/Y NAND2X1_LOC_858/B 0.02fF
C22903 NOR2X1_LOC_736/Y INVX1_LOC_96/Y 0.04fF
C22904 INVX1_LOC_50/A INVX1_LOC_19/A 2.34fF
C22905 NOR2X1_LOC_160/B INVX1_LOC_37/A 0.50fF
C22906 NAND2X1_LOC_558/a_36_24# NOR2X1_LOC_536/A 0.00fF
C22907 NAND2X1_LOC_9/Y NOR2X1_LOC_814/A 0.03fF
C22908 NOR2X1_LOC_606/Y INVX1_LOC_76/A 0.01fF
C22909 INVX1_LOC_292/Y NOR2X1_LOC_801/A 0.03fF
C22910 NOR2X1_LOC_590/A INVX1_LOC_46/A 0.11fF
C22911 INVX1_LOC_233/A INVX1_LOC_265/Y 0.00fF
C22912 NOR2X1_LOC_160/B NOR2X1_LOC_231/A 0.01fF
C22913 NOR2X1_LOC_717/B NOR2X1_LOC_374/B 0.00fF
C22914 NAND2X1_LOC_541/Y INPUT_1 0.01fF
C22915 INVX1_LOC_5/A INVX1_LOC_260/Y 0.01fF
C22916 NAND2X1_LOC_553/a_36_24# INVX1_LOC_89/A 0.00fF
C22917 NAND2X1_LOC_475/Y NOR2X1_LOC_678/A 0.00fF
C22918 NOR2X1_LOC_590/A NOR2X1_LOC_98/A 0.01fF
C22919 NOR2X1_LOC_219/Y NOR2X1_LOC_214/B 0.03fF
C22920 NOR2X1_LOC_71/Y INVX1_LOC_22/A 0.00fF
C22921 NAND2X1_LOC_214/B INVX1_LOC_123/Y 0.03fF
C22922 INVX1_LOC_24/A NAND2X1_LOC_655/A 0.01fF
C22923 INVX1_LOC_26/A INVX1_LOC_42/A 0.06fF
C22924 NOR2X1_LOC_124/B INPUT_0 0.01fF
C22925 NOR2X1_LOC_238/Y NAND2X1_LOC_623/B 0.00fF
C22926 NOR2X1_LOC_598/B NAND2X1_LOC_782/B 0.02fF
C22927 INVX1_LOC_224/Y NAND2X1_LOC_74/B 0.34fF
C22928 NOR2X1_LOC_38/a_36_216# INVX1_LOC_23/Y 0.01fF
C22929 INVX1_LOC_171/A INVX1_LOC_1/Y 0.08fF
C22930 INVX1_LOC_157/A NOR2X1_LOC_561/Y 0.03fF
C22931 NOR2X1_LOC_654/A INVX1_LOC_261/Y 0.01fF
C22932 INVX1_LOC_224/A INVX1_LOC_9/A -0.04fF
C22933 INVX1_LOC_64/A INVX1_LOC_63/A 0.07fF
C22934 NOR2X1_LOC_152/Y NOR2X1_LOC_269/Y 0.06fF
C22935 INVX1_LOC_311/Y INVX1_LOC_83/Y 0.01fF
C22936 NOR2X1_LOC_78/B NOR2X1_LOC_741/a_36_216# 0.00fF
C22937 INVX1_LOC_2/A NAND2X1_LOC_840/Y 0.02fF
C22938 NOR2X1_LOC_802/A INPUT_0 0.07fF
C22939 INVX1_LOC_49/A NOR2X1_LOC_78/A 0.15fF
C22940 INVX1_LOC_11/A INVX1_LOC_9/A 0.14fF
C22941 NOR2X1_LOC_188/A NOR2X1_LOC_87/B 0.03fF
C22942 INVX1_LOC_24/A NAND2X1_LOC_468/B 0.00fF
C22943 NOR2X1_LOC_644/A INVX1_LOC_22/A 0.06fF
C22944 NAND2X1_LOC_860/A INVX1_LOC_29/A 5.19fF
C22945 NAND2X1_LOC_35/Y NAND2X1_LOC_768/Y 0.03fF
C22946 INVX1_LOC_44/Y NOR2X1_LOC_208/A 0.24fF
C22947 NOR2X1_LOC_763/Y INVX1_LOC_83/A 0.10fF
C22948 NAND2X1_LOC_358/Y INVX1_LOC_89/A 0.03fF
C22949 NOR2X1_LOC_724/Y NOR2X1_LOC_730/Y 0.49fF
C22950 INVX1_LOC_24/Y INVX1_LOC_307/A 0.02fF
C22951 NOR2X1_LOC_798/A NOR2X1_LOC_814/A 0.06fF
C22952 NOR2X1_LOC_735/a_36_216# NOR2X1_LOC_357/Y 0.01fF
C22953 INVX1_LOC_279/A NOR2X1_LOC_180/B 1.01fF
C22954 NOR2X1_LOC_255/Y INVX1_LOC_42/A 0.02fF
C22955 INVX1_LOC_24/Y NOR2X1_LOC_445/B 0.10fF
C22956 NOR2X1_LOC_551/Y INVX1_LOC_177/A 0.01fF
C22957 NOR2X1_LOC_543/A NOR2X1_LOC_356/A 0.01fF
C22958 NAND2X1_LOC_27/a_36_24# INVX1_LOC_63/A 0.00fF
C22959 NAND2X1_LOC_703/Y INVX1_LOC_285/A 0.01fF
C22960 INVX1_LOC_89/A NOR2X1_LOC_99/B 0.21fF
C22961 INVX1_LOC_181/Y VDD 1.12fF
C22962 INVX1_LOC_13/Y NAND2X1_LOC_773/B 0.21fF
C22963 NOR2X1_LOC_233/a_36_216# NAND2X1_LOC_489/Y 0.00fF
C22964 INVX1_LOC_163/A NOR2X1_LOC_649/B 0.01fF
C22965 NAND2X1_LOC_110/a_36_24# INVX1_LOC_158/Y 0.00fF
C22966 NOR2X1_LOC_673/A NAND2X1_LOC_218/A 0.22fF
C22967 INVX1_LOC_78/A INVX1_LOC_26/A 0.47fF
C22968 INVX1_LOC_31/A INVX1_LOC_185/A 0.03fF
C22969 NAND2X1_LOC_508/A NOR2X1_LOC_99/B 0.03fF
C22970 INVX1_LOC_2/A NOR2X1_LOC_78/A 0.01fF
C22971 INVX1_LOC_279/A INVX1_LOC_73/A 0.02fF
C22972 NOR2X1_LOC_226/A INVX1_LOC_98/A 0.76fF
C22973 INVX1_LOC_286/A INVX1_LOC_25/Y 0.55fF
C22974 INVX1_LOC_21/A NOR2X1_LOC_340/A 0.13fF
C22975 NAND2X1_LOC_563/Y NAND2X1_LOC_659/B 0.02fF
C22976 NOR2X1_LOC_226/A NOR2X1_LOC_78/A 0.07fF
C22977 NOR2X1_LOC_474/A INVX1_LOC_194/Y 0.01fF
C22978 NOR2X1_LOC_596/A INVX1_LOC_281/Y 0.01fF
C22979 NOR2X1_LOC_281/Y NAND2X1_LOC_286/B 0.00fF
C22980 INVX1_LOC_89/A INVX1_LOC_182/A 0.07fF
C22981 INVX1_LOC_34/A INVX1_LOC_2/Y 0.07fF
C22982 NOR2X1_LOC_489/B INVX1_LOC_47/Y 0.01fF
C22983 NOR2X1_LOC_65/B INVX1_LOC_26/A 0.15fF
C22984 NOR2X1_LOC_220/A NOR2X1_LOC_562/B 0.06fF
C22985 INVX1_LOC_29/A NAND2X1_LOC_473/A 0.07fF
C22986 NOR2X1_LOC_759/Y NOR2X1_LOC_331/B 0.02fF
C22987 NOR2X1_LOC_317/B INVX1_LOC_37/A 0.01fF
C22988 NOR2X1_LOC_52/B NAND2X1_LOC_649/a_36_24# 0.00fF
C22989 INVX1_LOC_208/A NAND2X1_LOC_329/a_36_24# 0.01fF
C22990 NOR2X1_LOC_6/B NOR2X1_LOC_857/A 0.05fF
C22991 NOR2X1_LOC_561/Y INVX1_LOC_69/Y 0.01fF
C22992 NOR2X1_LOC_447/Y INVX1_LOC_38/A 0.03fF
C22993 INVX1_LOC_202/A NOR2X1_LOC_331/B 0.31fF
C22994 INVX1_LOC_50/A INVX1_LOC_26/Y 3.04fF
C22995 NOR2X1_LOC_92/Y INVX1_LOC_12/A 1.59fF
C22996 INVX1_LOC_136/A NOR2X1_LOC_79/a_36_216# 0.01fF
C22997 NOR2X1_LOC_218/Y NOR2X1_LOC_78/A 0.08fF
C22998 NAND2X1_LOC_563/Y VDD 0.92fF
C22999 NOR2X1_LOC_808/A NOR2X1_LOC_324/B 0.03fF
C23000 NOR2X1_LOC_689/A NAND2X1_LOC_724/Y 0.01fF
C23001 INVX1_LOC_34/A NOR2X1_LOC_363/Y 0.05fF
C23002 NAND2X1_LOC_181/Y INVX1_LOC_95/Y 0.04fF
C23003 INVX1_LOC_43/Y INVX1_LOC_63/A 0.03fF
C23004 INVX1_LOC_18/A INVX1_LOC_179/A 0.11fF
C23005 NAND2X1_LOC_67/Y NOR2X1_LOC_89/A 0.15fF
C23006 NOR2X1_LOC_71/Y INVX1_LOC_100/A 0.81fF
C23007 NOR2X1_LOC_589/A NOR2X1_LOC_318/B 0.03fF
C23008 NOR2X1_LOC_433/A INVX1_LOC_9/A 0.01fF
C23009 NAND2X1_LOC_634/Y INVX1_LOC_35/Y 0.18fF
C23010 INVX1_LOC_240/A NAND2X1_LOC_804/Y 0.12fF
C23011 NOR2X1_LOC_68/A NOR2X1_LOC_155/A 0.56fF
C23012 INVX1_LOC_13/Y NOR2X1_LOC_393/Y 0.03fF
C23013 NOR2X1_LOC_103/Y NAND2X1_LOC_74/B 0.07fF
C23014 INVX1_LOC_30/Y NOR2X1_LOC_405/A 0.00fF
C23015 NOR2X1_LOC_593/Y INVX1_LOC_9/A 0.14fF
C23016 INVX1_LOC_189/A INVX1_LOC_37/A 0.00fF
C23017 INVX1_LOC_35/A NOR2X1_LOC_541/B 0.01fF
C23018 INVX1_LOC_225/A NAND2X1_LOC_848/A 0.03fF
C23019 INVX1_LOC_182/Y INVX1_LOC_73/A 0.23fF
C23020 NOR2X1_LOC_589/A INVX1_LOC_93/Y 0.33fF
C23021 NAND2X1_LOC_724/Y NAND2X1_LOC_738/B 7.16fF
C23022 NAND2X1_LOC_357/A NAND2X1_LOC_807/B 0.07fF
C23023 INVX1_LOC_22/Y NOR2X1_LOC_68/Y 0.10fF
C23024 INVX1_LOC_144/Y NOR2X1_LOC_447/B 0.02fF
C23025 NOR2X1_LOC_720/B INVX1_LOC_38/A 0.01fF
C23026 INVX1_LOC_23/A INVX1_LOC_270/Y 0.17fF
C23027 NAND2X1_LOC_79/Y NOR2X1_LOC_216/B 0.02fF
C23028 NOR2X1_LOC_423/Y INVX1_LOC_281/A 0.01fF
C23029 INVX1_LOC_61/Y INVX1_LOC_19/A 0.52fF
C23030 NAND2X1_LOC_783/A NAND2X1_LOC_655/A 0.06fF
C23031 INVX1_LOC_2/A NOR2X1_LOC_60/Y 0.07fF
C23032 NAND2X1_LOC_556/a_36_24# NOR2X1_LOC_536/A 0.00fF
C23033 INVX1_LOC_196/A INVX1_LOC_117/A 0.03fF
C23034 INVX1_LOC_1/Y INVX1_LOC_20/A 0.03fF
C23035 NOR2X1_LOC_488/Y INVX1_LOC_46/A 0.00fF
C23036 NOR2X1_LOC_431/a_36_216# NOR2X1_LOC_697/Y 0.00fF
C23037 NOR2X1_LOC_736/Y NOR2X1_LOC_733/Y 0.15fF
C23038 INVX1_LOC_57/A NOR2X1_LOC_717/A 0.22fF
C23039 NOR2X1_LOC_52/B INVX1_LOC_9/A 0.03fF
C23040 NOR2X1_LOC_82/Y INVX1_LOC_46/A 0.03fF
C23041 INVX1_LOC_14/A INVX1_LOC_47/Y 0.19fF
C23042 NOR2X1_LOC_392/Y NAND2X1_LOC_215/A 0.18fF
C23043 NAND2X1_LOC_840/B NOR2X1_LOC_111/A 0.06fF
C23044 D_INPUT_0 NAND2X1_LOC_642/Y 0.10fF
C23045 INVX1_LOC_98/A INPUT_1 0.18fF
C23046 NOR2X1_LOC_769/a_36_216# INVX1_LOC_117/A 0.01fF
C23047 NOR2X1_LOC_320/a_36_216# INVX1_LOC_54/A 0.00fF
C23048 NOR2X1_LOC_516/B INVX1_LOC_37/A 0.02fF
C23049 NOR2X1_LOC_78/A INPUT_1 0.33fF
C23050 INVX1_LOC_32/Y VDD 0.21fF
C23051 INVX1_LOC_41/A INVX1_LOC_307/A 0.07fF
C23052 NOR2X1_LOC_222/Y INVX1_LOC_281/A 0.08fF
C23053 NOR2X1_LOC_589/A INVX1_LOC_139/A 0.01fF
C23054 INVX1_LOC_171/A INVX1_LOC_93/Y 0.08fF
C23055 INVX1_LOC_45/A NAND2X1_LOC_74/B 0.10fF
C23056 INVX1_LOC_53/Y INVX1_LOC_12/Y 0.01fF
C23057 INVX1_LOC_177/A NOR2X1_LOC_729/A 0.03fF
C23058 NOR2X1_LOC_130/A NAND2X1_LOC_468/B 0.03fF
C23059 NOR2X1_LOC_15/Y INVX1_LOC_253/A 0.03fF
C23060 INVX1_LOC_298/A NOR2X1_LOC_383/B 0.00fF
C23061 NOR2X1_LOC_568/A NAND2X1_LOC_74/B 0.11fF
C23062 INVX1_LOC_157/A INVX1_LOC_76/A 0.03fF
C23063 INVX1_LOC_41/A NOR2X1_LOC_445/B 0.07fF
C23064 INVX1_LOC_34/A NOR2X1_LOC_608/Y 0.00fF
C23065 NOR2X1_LOC_637/B NOR2X1_LOC_697/Y 0.26fF
C23066 NOR2X1_LOC_457/a_36_216# NOR2X1_LOC_464/Y 0.00fF
C23067 NOR2X1_LOC_175/A NOR2X1_LOC_641/Y 0.02fF
C23068 INVX1_LOC_286/A INVX1_LOC_75/A 0.08fF
C23069 INVX1_LOC_135/A NOR2X1_LOC_347/a_36_216# 0.00fF
C23070 INVX1_LOC_120/A NOR2X1_LOC_332/B 0.22fF
C23071 NOR2X1_LOC_329/B NOR2X1_LOC_45/B 0.23fF
C23072 INVX1_LOC_268/A INVX1_LOC_117/A 0.00fF
C23073 INVX1_LOC_104/A INVX1_LOC_92/A 0.07fF
C23074 INVX1_LOC_227/A INVX1_LOC_46/A 0.07fF
C23075 NAND2X1_LOC_391/Y INVX1_LOC_181/A 0.01fF
C23076 NAND2X1_LOC_622/B NAND2X1_LOC_621/a_36_24# 0.02fF
C23077 NAND2X1_LOC_562/B INVX1_LOC_260/Y 0.38fF
C23078 INVX1_LOC_221/Y INVX1_LOC_94/Y 0.01fF
C23079 NAND2X1_LOC_608/a_36_24# NOR2X1_LOC_717/A 0.07fF
C23080 NOR2X1_LOC_533/Y NAND2X1_LOC_175/Y 0.01fF
C23081 INVX1_LOC_33/A NOR2X1_LOC_691/A 0.01fF
C23082 VDD INVX1_LOC_148/Y 0.59fF
C23083 INVX1_LOC_6/A NOR2X1_LOC_368/a_36_216# 0.02fF
C23084 NOR2X1_LOC_68/A NOR2X1_LOC_833/B 0.03fF
C23085 INVX1_LOC_34/A NOR2X1_LOC_485/Y 0.05fF
C23086 INVX1_LOC_71/A NAND2X1_LOC_74/B 0.08fF
C23087 INVX1_LOC_25/Y INVX1_LOC_54/A 0.03fF
C23088 NOR2X1_LOC_678/A NOR2X1_LOC_840/A 0.15fF
C23089 NAND2X1_LOC_837/Y INVX1_LOC_12/A 0.08fF
C23090 NAND2X1_LOC_693/a_36_24# NOR2X1_LOC_486/Y 0.00fF
C23091 INVX1_LOC_122/Y INVX1_LOC_15/A 0.16fF
C23092 INVX1_LOC_163/A NOR2X1_LOC_476/B 0.01fF
C23093 NAND2X1_LOC_465/Y NAND2X1_LOC_768/Y 0.22fF
C23094 NAND2X1_LOC_832/Y INVX1_LOC_199/A 0.01fF
C23095 NOR2X1_LOC_500/B NAND2X1_LOC_615/a_36_24# 0.06fF
C23096 INVX1_LOC_41/A INVX1_LOC_12/A 0.10fF
C23097 INVX1_LOC_50/A INVX1_LOC_161/Y 0.08fF
C23098 NOR2X1_LOC_516/Y INVX1_LOC_29/A 0.13fF
C23099 NOR2X1_LOC_498/Y INVX1_LOC_12/A 0.07fF
C23100 INVX1_LOC_232/Y INVX1_LOC_84/A 0.00fF
C23101 NOR2X1_LOC_706/A INVX1_LOC_37/A 0.01fF
C23102 NAND2X1_LOC_162/B NOR2X1_LOC_467/A 0.06fF
C23103 NAND2X1_LOC_84/Y INVX1_LOC_47/Y 0.08fF
C23104 NAND2X1_LOC_850/Y INVX1_LOC_63/A 0.25fF
C23105 NOR2X1_LOC_332/A NOR2X1_LOC_660/a_36_216# 0.01fF
C23106 INVX1_LOC_182/Y NOR2X1_LOC_122/a_36_216# 0.00fF
C23107 NAND2X1_LOC_477/A INVX1_LOC_12/A 0.07fF
C23108 NOR2X1_LOC_457/A NOR2X1_LOC_678/A 0.00fF
C23109 INVX1_LOC_89/A NOR2X1_LOC_622/a_36_216# 0.00fF
C23110 NOR2X1_LOC_207/A INVX1_LOC_12/A 0.03fF
C23111 NOR2X1_LOC_763/A D_INPUT_6 0.10fF
C23112 INPUT_0 NOR2X1_LOC_363/Y 0.02fF
C23113 NOR2X1_LOC_67/A NAND2X1_LOC_81/B 0.02fF
C23114 NOR2X1_LOC_369/a_36_216# INVX1_LOC_42/A 0.00fF
C23115 INVX1_LOC_50/A NOR2X1_LOC_599/A 0.03fF
C23116 D_INPUT_6 NOR2X1_LOC_582/A 0.11fF
C23117 INVX1_LOC_18/A NOR2X1_LOC_693/Y 0.07fF
C23118 NOR2X1_LOC_577/Y INVX1_LOC_21/Y 0.34fF
C23119 NAND2X1_LOC_734/B NOR2X1_LOC_48/B 0.02fF
C23120 NOR2X1_LOC_272/Y NOR2X1_LOC_15/Y 0.03fF
C23121 NOR2X1_LOC_859/a_36_216# INVX1_LOC_5/A 0.02fF
C23122 NAND2X1_LOC_9/Y NOR2X1_LOC_590/A 0.11fF
C23123 NOR2X1_LOC_725/A INVX1_LOC_76/A 0.19fF
C23124 INVX1_LOC_10/A NOR2X1_LOC_435/B 0.03fF
C23125 NAND2X1_LOC_807/Y INVX1_LOC_185/A 0.00fF
C23126 NOR2X1_LOC_478/A NOR2X1_LOC_598/B 0.01fF
C23127 INVX1_LOC_136/A INVX1_LOC_224/Y 0.10fF
C23128 INVX1_LOC_21/A INVX1_LOC_103/A 0.07fF
C23129 INVX1_LOC_75/A INVX1_LOC_54/A 0.11fF
C23130 NOR2X1_LOC_778/B INVX1_LOC_290/Y 0.10fF
C23131 NOR2X1_LOC_706/B INVX1_LOC_91/A 0.00fF
C23132 INVX1_LOC_230/Y INVX1_LOC_5/A 0.14fF
C23133 NOR2X1_LOC_266/B NAND2X1_LOC_642/Y 0.02fF
C23134 INVX1_LOC_30/A NOR2X1_LOC_678/A 0.10fF
C23135 NOR2X1_LOC_612/B INVX1_LOC_47/Y 0.03fF
C23136 NAND2X1_LOC_860/A NOR2X1_LOC_82/a_36_216# 0.00fF
C23137 NOR2X1_LOC_769/B NOR2X1_LOC_68/A 0.01fF
C23138 NOR2X1_LOC_746/a_36_216# INVX1_LOC_117/A 0.01fF
C23139 NAND2X1_LOC_860/A NAND2X1_LOC_634/Y 0.18fF
C23140 NOR2X1_LOC_675/A VDD -0.00fF
C23141 INVX1_LOC_45/A NAND2X1_LOC_358/B 0.02fF
C23142 INVX1_LOC_172/A NOR2X1_LOC_693/Y 0.07fF
C23143 INVX1_LOC_74/Y D_INPUT_3 0.01fF
C23144 NOR2X1_LOC_453/Y INVX1_LOC_103/A 0.00fF
C23145 INVX1_LOC_177/Y INVX1_LOC_53/A 0.03fF
C23146 NAND2X1_LOC_109/a_36_24# INVX1_LOC_37/A 0.00fF
C23147 INVX1_LOC_50/A NOR2X1_LOC_437/Y 0.07fF
C23148 INVX1_LOC_27/A INPUT_2 0.23fF
C23149 NOR2X1_LOC_598/B NOR2X1_LOC_68/A 3.54fF
C23150 VDD NOR2X1_LOC_833/Y 0.39fF
C23151 INVX1_LOC_232/Y INVX1_LOC_15/A 0.03fF
C23152 INVX1_LOC_21/A INVX1_LOC_292/A 0.08fF
C23153 NOR2X1_LOC_590/A NOR2X1_LOC_798/A 0.05fF
C23154 INVX1_LOC_58/A NOR2X1_LOC_238/Y 0.01fF
C23155 INVX1_LOC_18/A NOR2X1_LOC_405/Y 0.01fF
C23156 INVX1_LOC_230/Y INVX1_LOC_178/A 0.03fF
C23157 NOR2X1_LOC_690/A INVX1_LOC_23/Y 0.15fF
C23158 NOR2X1_LOC_430/A INVX1_LOC_57/A 0.32fF
C23159 NOR2X1_LOC_636/A INVX1_LOC_262/A 0.00fF
C23160 INVX1_LOC_83/Y INVX1_LOC_15/A 0.01fF
C23161 VDD INVX1_LOC_115/A 0.00fF
C23162 NAND2X1_LOC_842/B NOR2X1_LOC_814/A 0.01fF
C23163 NOR2X1_LOC_561/Y NOR2X1_LOC_89/A 0.01fF
C23164 INVX1_LOC_121/A INVX1_LOC_12/A 0.04fF
C23165 INVX1_LOC_197/Y INVX1_LOC_15/A 0.00fF
C23166 INVX1_LOC_95/Y INVX1_LOC_117/A 0.04fF
C23167 NAND2X1_LOC_222/B NAND2X1_LOC_20/B 0.22fF
C23168 NOR2X1_LOC_75/Y INVX1_LOC_1/A 0.04fF
C23169 INVX1_LOC_149/A INVX1_LOC_78/A 0.07fF
C23170 NAND2X1_LOC_364/Y INVX1_LOC_57/A 0.03fF
C23171 NAND2X1_LOC_650/B INVX1_LOC_46/A 0.07fF
C23172 INVX1_LOC_78/Y INVX1_LOC_274/A 0.01fF
C23173 INVX1_LOC_98/A INVX1_LOC_118/A 0.02fF
C23174 NOR2X1_LOC_67/A INVX1_LOC_4/Y 0.10fF
C23175 INVX1_LOC_56/Y INVX1_LOC_32/A 0.01fF
C23176 NAND2X1_LOC_721/A INVX1_LOC_20/A 0.11fF
C23177 INVX1_LOC_25/A NOR2X1_LOC_716/B 0.07fF
C23178 NOR2X1_LOC_69/A INVX1_LOC_281/A 0.05fF
C23179 NOR2X1_LOC_92/Y NAND2X1_LOC_733/Y 0.10fF
C23180 INVX1_LOC_135/A NAND2X1_LOC_206/B 0.00fF
C23181 INVX1_LOC_1/Y INVX1_LOC_4/A 0.06fF
C23182 INVX1_LOC_34/A INVX1_LOC_29/Y 0.03fF
C23183 NOR2X1_LOC_860/B INVX1_LOC_138/Y 0.03fF
C23184 INVX1_LOC_36/A NOR2X1_LOC_440/B 0.01fF
C23185 NOR2X1_LOC_470/A NOR2X1_LOC_467/A 0.08fF
C23186 INVX1_LOC_233/Y NOR2X1_LOC_753/Y 0.01fF
C23187 NOR2X1_LOC_347/a_36_216# INVX1_LOC_280/A 0.01fF
C23188 INVX1_LOC_13/Y INVX1_LOC_24/A 0.14fF
C23189 NAND2X1_LOC_860/A INVX1_LOC_8/A 0.17fF
C23190 NAND2X1_LOC_303/Y NAND2X1_LOC_741/B 0.03fF
C23191 NOR2X1_LOC_563/a_36_216# NOR2X1_LOC_334/Y 0.01fF
C23192 NOR2X1_LOC_560/A NAND2X1_LOC_206/B 0.18fF
C23193 NAND2X1_LOC_755/a_36_24# NAND2X1_LOC_215/A 0.00fF
C23194 NOR2X1_LOC_391/Y INVX1_LOC_84/A 0.01fF
C23195 NOR2X1_LOC_92/Y INVX1_LOC_217/A 0.08fF
C23196 NOR2X1_LOC_719/B NOR2X1_LOC_38/B 0.01fF
C23197 INVX1_LOC_104/A INVX1_LOC_53/A 0.20fF
C23198 NAND2X1_LOC_642/Y INVX1_LOC_46/Y 0.02fF
C23199 NAND2X1_LOC_464/A INVX1_LOC_118/A 0.02fF
C23200 INVX1_LOC_254/Y INVX1_LOC_50/Y 0.05fF
C23201 NOR2X1_LOC_15/Y NAND2X1_LOC_364/A 0.03fF
C23202 NOR2X1_LOC_772/B NOR2X1_LOC_557/Y 0.42fF
C23203 NOR2X1_LOC_312/Y INVX1_LOC_15/A 0.07fF
C23204 D_INPUT_4 NOR2X1_LOC_1/Y 0.01fF
C23205 INVX1_LOC_71/A NAND2X1_LOC_793/a_36_24# 0.00fF
C23206 INVX1_LOC_25/Y NOR2X1_LOC_438/Y 0.07fF
C23207 NOR2X1_LOC_186/Y INVX1_LOC_49/A 0.07fF
C23208 INVX1_LOC_280/Y NAND2X1_LOC_787/Y 0.00fF
C23209 INVX1_LOC_17/A NOR2X1_LOC_372/Y 0.01fF
C23210 NOR2X1_LOC_667/Y INVX1_LOC_31/A 0.01fF
C23211 INVX1_LOC_45/A NOR2X1_LOC_307/A 0.03fF
C23212 INVX1_LOC_103/A NAND2X1_LOC_354/Y 0.02fF
C23213 INVX1_LOC_21/A NAND2X1_LOC_681/a_36_24# 0.00fF
C23214 NAND2X1_LOC_453/A INVX1_LOC_54/A 0.79fF
C23215 NAND2X1_LOC_123/Y INVX1_LOC_290/Y 0.21fF
C23216 INVX1_LOC_136/A NOR2X1_LOC_103/Y 0.24fF
C23217 INVX1_LOC_13/Y NOR2X1_LOC_557/Y 0.07fF
C23218 NOR2X1_LOC_586/a_36_216# NOR2X1_LOC_158/Y 0.01fF
C23219 NAND2X1_LOC_36/A INVX1_LOC_174/A 0.58fF
C23220 INVX1_LOC_58/A NAND2X1_LOC_54/a_36_24# 0.00fF
C23221 NAND2X1_LOC_377/Y INVX1_LOC_175/A 0.01fF
C23222 NAND2X1_LOC_87/a_36_24# NOR2X1_LOC_52/B 0.00fF
C23223 INVX1_LOC_21/A INVX1_LOC_67/A 0.02fF
C23224 NOR2X1_LOC_361/B INVX1_LOC_181/Y 0.42fF
C23225 NOR2X1_LOC_401/A NAND2X1_LOC_198/B 0.02fF
C23226 INVX1_LOC_58/A NAND2X1_LOC_841/A 0.03fF
C23227 INVX1_LOC_88/A INVX1_LOC_24/A 0.06fF
C23228 INVX1_LOC_313/Y NAND2X1_LOC_647/B 0.02fF
C23229 NOR2X1_LOC_655/B NOR2X1_LOC_392/Y 0.10fF
C23230 INVX1_LOC_39/A NAND2X1_LOC_139/A 0.01fF
C23231 NOR2X1_LOC_772/a_36_216# INVX1_LOC_29/Y 0.00fF
C23232 INVX1_LOC_171/A INVX1_LOC_87/A 0.04fF
C23233 INVX1_LOC_64/A NOR2X1_LOC_362/a_36_216# 0.00fF
C23234 INVX1_LOC_20/A NAND2X1_LOC_770/Y 0.01fF
C23235 NOR2X1_LOC_537/A INVX1_LOC_1/A 0.00fF
C23236 NOR2X1_LOC_71/a_36_216# INVX1_LOC_12/A 0.00fF
C23237 INVX1_LOC_58/A INVX1_LOC_268/A 0.02fF
C23238 NAND2X1_LOC_860/A NOR2X1_LOC_315/a_36_216# 0.01fF
C23239 NOR2X1_LOC_545/B NOR2X1_LOC_814/A 0.01fF
C23240 NOR2X1_LOC_772/B INVX1_LOC_143/A 0.01fF
C23241 INVX1_LOC_1/A NOR2X1_LOC_716/B 0.10fF
C23242 NAND2X1_LOC_391/Y NOR2X1_LOC_315/Y 0.02fF
C23243 NOR2X1_LOC_160/B NAND2X1_LOC_198/B 0.47fF
C23244 NAND2X1_LOC_778/Y NAND2X1_LOC_785/A 0.10fF
C23245 NOR2X1_LOC_78/A NAND2X1_LOC_63/Y 1.68fF
C23246 INVX1_LOC_2/A NOR2X1_LOC_186/Y 0.14fF
C23247 INVX1_LOC_256/A NOR2X1_LOC_274/Y 0.02fF
C23248 INVX1_LOC_233/A NOR2X1_LOC_82/Y 0.03fF
C23249 INVX1_LOC_45/A INVX1_LOC_136/A 0.06fF
C23250 INVX1_LOC_13/Y INVX1_LOC_143/A 0.07fF
C23251 INVX1_LOC_17/A NAND2X1_LOC_585/a_36_24# 0.00fF
C23252 INVX1_LOC_305/A INVX1_LOC_30/A 0.30fF
C23253 INVX1_LOC_136/A NOR2X1_LOC_568/A 0.10fF
C23254 NOR2X1_LOC_276/Y INVX1_LOC_71/A 0.03fF
C23255 NAND2X1_LOC_22/a_36_24# NAND2X1_LOC_30/Y 0.00fF
C23256 NAND2X1_LOC_715/a_36_24# INVX1_LOC_271/A 0.00fF
C23257 NAND2X1_LOC_35/Y INVX1_LOC_226/Y 0.23fF
C23258 NOR2X1_LOC_528/Y INVX1_LOC_102/A 0.10fF
C23259 INVX1_LOC_136/A NAND2X1_LOC_856/A 0.03fF
C23260 NOR2X1_LOC_765/Y NAND2X1_LOC_770/Y 0.00fF
C23261 NOR2X1_LOC_831/B INVX1_LOC_66/Y 0.03fF
C23262 NAND2X1_LOC_67/Y NOR2X1_LOC_52/B 0.10fF
C23263 NOR2X1_LOC_218/A INVX1_LOC_33/A 0.01fF
C23264 NAND2X1_LOC_341/A INVX1_LOC_5/A 0.68fF
C23265 INVX1_LOC_2/A NAND2X1_LOC_573/Y 0.62fF
C23266 INVX1_LOC_46/Y NOR2X1_LOC_271/Y 0.03fF
C23267 INVX1_LOC_39/A NAND2X1_LOC_541/Y 0.01fF
C23268 INVX1_LOC_313/A INVX1_LOC_270/Y 0.34fF
C23269 NAND2X1_LOC_785/A NOR2X1_LOC_15/Y 0.01fF
C23270 NOR2X1_LOC_820/A NOR2X1_LOC_554/B 0.02fF
C23271 NOR2X1_LOC_750/Y D_INPUT_0 0.01fF
C23272 NOR2X1_LOC_791/B INVX1_LOC_72/Y 0.02fF
C23273 INVX1_LOC_200/Y INVX1_LOC_90/A 0.04fF
C23274 NAND2X1_LOC_565/B INVX1_LOC_13/Y -0.02fF
C23275 NOR2X1_LOC_160/B INVX1_LOC_310/Y 0.03fF
C23276 NOR2X1_LOC_382/Y D_INPUT_2 0.29fF
C23277 NAND2X1_LOC_35/B NAND2X1_LOC_725/B 0.04fF
C23278 INVX1_LOC_2/A NAND2X1_LOC_724/A 0.01fF
C23279 NAND2X1_LOC_785/B NOR2X1_LOC_495/Y 0.10fF
C23280 VDD NAND2X1_LOC_500/B 0.01fF
C23281 INVX1_LOC_36/A NAND2X1_LOC_593/Y 0.07fF
C23282 VDD NOR2X1_LOC_509/A -0.00fF
C23283 INVX1_LOC_11/A NAND2X1_LOC_629/Y 0.00fF
C23284 INVX1_LOC_136/A INVX1_LOC_71/A 0.34fF
C23285 INVX1_LOC_217/A NAND2X1_LOC_837/Y 0.10fF
C23286 INVX1_LOC_215/Y NOR2X1_LOC_574/A 0.01fF
C23287 NOR2X1_LOC_829/Y NAND2X1_LOC_855/Y 0.06fF
C23288 NOR2X1_LOC_669/A INVX1_LOC_20/A 0.01fF
C23289 NAND2X1_LOC_862/Y NAND2X1_LOC_793/B 0.03fF
C23290 NOR2X1_LOC_498/Y NAND2X1_LOC_733/Y 0.07fF
C23291 NOR2X1_LOC_89/A INVX1_LOC_76/A 0.82fF
C23292 INVX1_LOC_25/A NOR2X1_LOC_120/a_36_216# 0.00fF
C23293 NOR2X1_LOC_598/B NOR2X1_LOC_163/A 0.00fF
C23294 NOR2X1_LOC_457/B NOR2X1_LOC_596/A 0.08fF
C23295 INVX1_LOC_230/Y NAND2X1_LOC_562/B 0.06fF
C23296 INVX1_LOC_2/A NOR2X1_LOC_215/a_36_216# 0.01fF
C23297 NOR2X1_LOC_331/Y NOR2X1_LOC_52/B 0.05fF
C23298 INVX1_LOC_199/Y NOR2X1_LOC_477/B 0.01fF
C23299 NOR2X1_LOC_446/a_36_216# NOR2X1_LOC_348/B 0.01fF
C23300 INVX1_LOC_17/A NAND2X1_LOC_374/Y 0.04fF
C23301 NOR2X1_LOC_634/A NOR2X1_LOC_461/A 0.01fF
C23302 NOR2X1_LOC_288/a_36_216# NOR2X1_LOC_634/B 0.00fF
C23303 INVX1_LOC_11/A INVX1_LOC_243/A 0.01fF
C23304 NAND2X1_LOC_213/A NAND2X1_LOC_160/a_36_24# 0.01fF
C23305 INVX1_LOC_95/Y INVX1_LOC_3/Y 0.20fF
C23306 NOR2X1_LOC_91/A INVX1_LOC_126/Y 0.01fF
C23307 INVX1_LOC_93/Y INVX1_LOC_4/A 0.20fF
C23308 INVX1_LOC_91/A INVX1_LOC_94/Y 0.00fF
C23309 INVX1_LOC_13/Y NOR2X1_LOC_130/A 0.07fF
C23310 INVX1_LOC_2/A NOR2X1_LOC_45/Y 0.00fF
C23311 INVX1_LOC_269/A INVX1_LOC_16/A 0.08fF
C23312 VDD NOR2X1_LOC_114/Y 0.41fF
C23313 NOR2X1_LOC_48/B NAND2X1_LOC_453/A 0.10fF
C23314 INVX1_LOC_303/A INVX1_LOC_24/A 0.07fF
C23315 NOR2X1_LOC_612/Y INVX1_LOC_294/A 0.01fF
C23316 NAND2X1_LOC_390/a_36_24# INVX1_LOC_14/A 0.00fF
C23317 NAND2X1_LOC_1/Y D_INPUT_5 0.02fF
C23318 NOR2X1_LOC_15/Y NOR2X1_LOC_86/A 0.08fF
C23319 NOR2X1_LOC_391/A INVX1_LOC_48/Y 0.07fF
C23320 INVX1_LOC_58/A NOR2X1_LOC_594/a_36_216# 0.00fF
C23321 NOR2X1_LOC_498/Y INVX1_LOC_217/A -0.00fF
C23322 NOR2X1_LOC_216/B INVX1_LOC_123/Y 0.21fF
C23323 NOR2X1_LOC_510/B NOR2X1_LOC_697/Y 0.10fF
C23324 NOR2X1_LOC_554/B INVX1_LOC_315/A 0.03fF
C23325 NOR2X1_LOC_401/a_36_216# NOR2X1_LOC_160/B 0.00fF
C23326 INPUT_0 INVX1_LOC_29/Y 0.03fF
C23327 INVX1_LOC_314/Y INVX1_LOC_77/A 0.07fF
C23328 INVX1_LOC_90/A NOR2X1_LOC_406/A 0.04fF
C23329 INVX1_LOC_21/A INVX1_LOC_120/A 0.09fF
C23330 NAND2X1_LOC_784/A NOR2X1_LOC_527/Y 0.02fF
C23331 NAND2X1_LOC_787/B NAND2X1_LOC_837/Y 0.12fF
C23332 INVX1_LOC_61/A NAND2X1_LOC_139/A 0.04fF
C23333 NOR2X1_LOC_331/B NAND2X1_LOC_74/B 0.07fF
C23334 NOR2X1_LOC_124/B INVX1_LOC_72/Y 0.05fF
C23335 NAND2X1_LOC_59/a_36_24# INVX1_LOC_174/A 0.00fF
C23336 INVX1_LOC_206/A INVX1_LOC_223/A 0.02fF
C23337 NAND2X1_LOC_287/B INVX1_LOC_15/A 0.02fF
C23338 NOR2X1_LOC_219/Y NOR2X1_LOC_160/B 0.17fF
C23339 NOR2X1_LOC_861/a_36_216# NAND2X1_LOC_206/Y 0.01fF
C23340 INVX1_LOC_1/A NOR2X1_LOC_326/Y 0.04fF
C23341 NOR2X1_LOC_717/B INVX1_LOC_1/A 0.03fF
C23342 NOR2X1_LOC_82/A NOR2X1_LOC_589/A 0.04fF
C23343 INVX1_LOC_132/A INVX1_LOC_49/A 0.06fF
C23344 NOR2X1_LOC_99/Y NAND2X1_LOC_773/B 0.07fF
C23345 NAND2X1_LOC_624/B NOR2X1_LOC_19/Y 0.10fF
C23346 NOR2X1_LOC_160/B INVX1_LOC_53/Y 0.03fF
C23347 INVX1_LOC_143/A NOR2X1_LOC_500/B 0.10fF
C23348 NAND2X1_LOC_481/a_36_24# NOR2X1_LOC_87/B 0.01fF
C23349 INVX1_LOC_219/A INVX1_LOC_14/A 0.00fF
C23350 NAND2X1_LOC_783/A INVX1_LOC_88/A 0.10fF
C23351 INVX1_LOC_280/A NAND2X1_LOC_206/B 0.02fF
C23352 INVX1_LOC_11/A NOR2X1_LOC_561/Y 0.07fF
C23353 INVX1_LOC_303/A NOR2X1_LOC_557/Y 0.35fF
C23354 NOR2X1_LOC_691/B NOR2X1_LOC_862/B 0.11fF
C23355 INVX1_LOC_91/A INVX1_LOC_296/A 0.09fF
C23356 NOR2X1_LOC_548/B INVX1_LOC_58/Y 0.10fF
C23357 NOR2X1_LOC_68/A NOR2X1_LOC_156/B 0.03fF
C23358 NOR2X1_LOC_309/Y INVX1_LOC_41/Y 0.01fF
C23359 NOR2X1_LOC_682/a_36_216# INVX1_LOC_273/A 0.00fF
C23360 INVX1_LOC_20/A INVX1_LOC_87/A 0.02fF
C23361 NAND2X1_LOC_579/A INVX1_LOC_89/A 0.09fF
C23362 INVX1_LOC_88/A NOR2X1_LOC_130/A 0.03fF
C23363 NOR2X1_LOC_219/a_36_216# INVX1_LOC_63/Y 0.01fF
C23364 NOR2X1_LOC_441/Y INVX1_LOC_25/Y 0.00fF
C23365 NOR2X1_LOC_468/Y NOR2X1_LOC_76/A 0.02fF
C23366 INVX1_LOC_206/Y INVX1_LOC_53/A 0.01fF
C23367 INVX1_LOC_119/Y INVX1_LOC_285/A 0.02fF
C23368 NOR2X1_LOC_498/Y NAND2X1_LOC_787/B 0.37fF
C23369 INVX1_LOC_249/A INVX1_LOC_85/A 0.49fF
C23370 NOR2X1_LOC_78/B INVX1_LOC_177/Y 0.10fF
C23371 INVX1_LOC_163/A INVX1_LOC_169/A 0.06fF
C23372 INVX1_LOC_225/A INVX1_LOC_49/A 0.08fF
C23373 NAND2X1_LOC_190/Y NOR2X1_LOC_180/B 0.07fF
C23374 NOR2X1_LOC_791/a_36_216# NAND2X1_LOC_338/B 0.00fF
C23375 INVX1_LOC_292/A NOR2X1_LOC_565/B 0.01fF
C23376 NAND2X1_LOC_114/a_36_24# NOR2X1_LOC_350/A 0.01fF
C23377 NOR2X1_LOC_717/B NOR2X1_LOC_794/B 0.00fF
C23378 NOR2X1_LOC_592/B NAND2X1_LOC_74/B 0.02fF
C23379 INVX1_LOC_5/A NOR2X1_LOC_391/a_36_216# 0.00fF
C23380 NAND2X1_LOC_350/B NAND2X1_LOC_198/B 0.04fF
C23381 INVX1_LOC_269/A INVX1_LOC_28/A 0.22fF
C23382 INVX1_LOC_271/Y INVX1_LOC_117/A 0.03fF
C23383 INVX1_LOC_35/A NOR2X1_LOC_45/B 0.10fF
C23384 NOR2X1_LOC_647/Y INVX1_LOC_255/Y -0.00fF
C23385 NAND2X1_LOC_733/Y NOR2X1_LOC_299/Y 0.03fF
C23386 INVX1_LOC_64/A NOR2X1_LOC_318/B 0.02fF
C23387 INVX1_LOC_58/A INVX1_LOC_187/Y 0.04fF
C23388 NOR2X1_LOC_246/A NAND2X1_LOC_352/B 0.02fF
C23389 INVX1_LOC_132/A INVX1_LOC_2/A 0.10fF
C23390 NOR2X1_LOC_570/B NOR2X1_LOC_348/B 1.03fF
C23391 NOR2X1_LOC_209/Y INVX1_LOC_49/A 0.07fF
C23392 INVX1_LOC_303/A INVX1_LOC_143/A 1.21fF
C23393 NOR2X1_LOC_778/B INVX1_LOC_77/A 0.03fF
C23394 NOR2X1_LOC_160/B NOR2X1_LOC_507/B 0.07fF
C23395 INVX1_LOC_202/A NOR2X1_LOC_366/B 0.30fF
C23396 NOR2X1_LOC_644/A NOR2X1_LOC_787/a_36_216# 0.00fF
C23397 INVX1_LOC_94/A NOR2X1_LOC_500/Y 0.21fF
C23398 INVX1_LOC_88/A NOR2X1_LOC_216/Y 0.14fF
C23399 INVX1_LOC_132/A NOR2X1_LOC_226/A 0.25fF
C23400 INVX1_LOC_260/Y INVX1_LOC_42/A 0.03fF
C23401 INVX1_LOC_33/A NOR2X1_LOC_131/A 0.01fF
C23402 NOR2X1_LOC_52/B NOR2X1_LOC_367/B 0.01fF
C23403 INVX1_LOC_58/A NOR2X1_LOC_305/Y 0.05fF
C23404 NOR2X1_LOC_809/B INVX1_LOC_15/A 0.15fF
C23405 NOR2X1_LOC_226/A NAND2X1_LOC_640/Y 0.02fF
C23406 NAND2X1_LOC_479/Y NOR2X1_LOC_759/Y 0.03fF
C23407 INPUT_2 NOR2X1_LOC_19/B 0.25fF
C23408 NOR2X1_LOC_590/A NAND2X1_LOC_842/B 0.00fF
C23409 INVX1_LOC_2/A INVX1_LOC_225/A 0.10fF
C23410 INVX1_LOC_202/A NAND2X1_LOC_479/Y 0.05fF
C23411 NOR2X1_LOC_831/B INVX1_LOC_32/A 0.03fF
C23412 NOR2X1_LOC_91/A NOR2X1_LOC_536/A 0.11fF
C23413 INVX1_LOC_136/A NOR2X1_LOC_123/B 0.94fF
C23414 INVX1_LOC_39/A NOR2X1_LOC_78/A 0.08fF
C23415 INVX1_LOC_181/Y NAND2X1_LOC_573/A 0.12fF
C23416 INVX1_LOC_18/A NOR2X1_LOC_71/Y 0.03fF
C23417 NOR2X1_LOC_226/A INVX1_LOC_225/A 0.07fF
C23418 D_INPUT_0 NOR2X1_LOC_91/Y 0.03fF
C23419 INVX1_LOC_103/A INVX1_LOC_311/A 0.01fF
C23420 NOR2X1_LOC_635/A NAND2X1_LOC_11/Y 0.22fF
C23421 INVX1_LOC_94/A INVX1_LOC_10/A 3.06fF
C23422 NOR2X1_LOC_78/B INVX1_LOC_104/A 2.20fF
C23423 NOR2X1_LOC_667/A INVX1_LOC_240/A 0.03fF
C23424 NAND2X1_LOC_731/Y NAND2X1_LOC_691/a_36_24# 0.01fF
C23425 NOR2X1_LOC_434/A NOR2X1_LOC_857/A 0.03fF
C23426 NAND2X1_LOC_639/A INVX1_LOC_23/A 0.12fF
C23427 INVX1_LOC_64/A INVX1_LOC_139/A 0.04fF
C23428 NOR2X1_LOC_635/a_36_216# INVX1_LOC_37/A 0.00fF
C23429 INVX1_LOC_301/A NAND2X1_LOC_782/a_36_24# 0.02fF
C23430 INVX1_LOC_215/A NOR2X1_LOC_577/Y 0.08fF
C23431 NOR2X1_LOC_570/B INVX1_LOC_22/A 0.12fF
C23432 NOR2X1_LOC_561/Y NOR2X1_LOC_433/A 0.14fF
C23433 INVX1_LOC_134/A NAND2X1_LOC_821/a_36_24# 0.00fF
C23434 NOR2X1_LOC_633/A INVX1_LOC_69/A 0.03fF
C23435 NOR2X1_LOC_536/A INVX1_LOC_23/A 0.07fF
C23436 NOR2X1_LOC_644/A INVX1_LOC_18/A 0.03fF
C23437 INVX1_LOC_226/Y NAND2X1_LOC_465/Y 0.01fF
C23438 INVX1_LOC_299/A INVX1_LOC_91/A 0.56fF
C23439 NOR2X1_LOC_160/B NOR2X1_LOC_113/B 0.03fF
C23440 INVX1_LOC_64/A NAND2X1_LOC_721/A 0.00fF
C23441 INVX1_LOC_41/A NOR2X1_LOC_730/A 0.02fF
C23442 INVX1_LOC_248/Y NOR2X1_LOC_305/Y 0.02fF
C23443 NOR2X1_LOC_15/Y NOR2X1_LOC_405/A 0.15fF
C23444 INVX1_LOC_136/A INVX1_LOC_102/Y 0.07fF
C23445 INVX1_LOC_116/A NOR2X1_LOC_389/B 0.01fF
C23446 NAND2X1_LOC_741/Y VDD 0.03fF
C23447 INVX1_LOC_21/A NOR2X1_LOC_137/Y 0.01fF
C23448 NAND2X1_LOC_182/A NAND2X1_LOC_392/Y 0.01fF
C23449 INVX1_LOC_34/A NOR2X1_LOC_355/A 0.07fF
C23450 INVX1_LOC_263/A NOR2X1_LOC_78/B 0.45fF
C23451 INVX1_LOC_35/A NOR2X1_LOC_499/B 0.04fF
C23452 INVX1_LOC_131/Y INVX1_LOC_270/Y 0.19fF
C23453 NOR2X1_LOC_61/B VDD -0.00fF
C23454 NOR2X1_LOC_561/Y NOR2X1_LOC_52/B 0.15fF
C23455 INVX1_LOC_5/A INVX1_LOC_44/A 0.04fF
C23456 NOR2X1_LOC_230/Y INVX1_LOC_6/A 0.34fF
C23457 NOR2X1_LOC_205/a_36_216# NOR2X1_LOC_500/Y 0.01fF
C23458 NAND2X1_LOC_361/Y INVX1_LOC_90/A 1.07fF
C23459 INVX1_LOC_289/Y INVX1_LOC_20/A 0.03fF
C23460 NAND2X1_LOC_579/A NAND2X1_LOC_244/A 0.04fF
C23461 INVX1_LOC_23/A NAND2X1_LOC_93/B 0.08fF
C23462 NOR2X1_LOC_778/B NOR2X1_LOC_687/Y 0.03fF
C23463 INVX1_LOC_269/A NOR2X1_LOC_35/Y 0.10fF
C23464 NAND2X1_LOC_640/Y INPUT_1 0.07fF
C23465 NOR2X1_LOC_202/Y NOR2X1_LOC_759/Y 0.01fF
C23466 NAND2X1_LOC_563/A INVX1_LOC_16/A 0.03fF
C23467 INVX1_LOC_77/A NAND2X1_LOC_123/Y 2.47fF
C23468 INVX1_LOC_50/A NOR2X1_LOC_841/A 0.01fF
C23469 NAND2X1_LOC_725/B VDD 0.25fF
C23470 NOR2X1_LOC_246/A NAND2X1_LOC_357/B 0.01fF
C23471 NOR2X1_LOC_865/A NOR2X1_LOC_849/A 0.11fF
C23472 INVX1_LOC_23/A NAND2X1_LOC_425/Y 0.02fF
C23473 INVX1_LOC_101/Y VDD 0.42fF
C23474 NAND2X1_LOC_861/Y NOR2X1_LOC_369/a_36_216# 0.01fF
C23475 NOR2X1_LOC_617/Y NOR2X1_LOC_19/Y 0.01fF
C23476 INVX1_LOC_90/A INVX1_LOC_219/Y 0.01fF
C23477 INVX1_LOC_11/A INVX1_LOC_76/A 0.46fF
C23478 NOR2X1_LOC_524/Y INVX1_LOC_91/A 0.10fF
C23479 NOR2X1_LOC_82/A INVX1_LOC_20/A 0.11fF
C23480 INVX1_LOC_57/A NOR2X1_LOC_697/Y 0.03fF
C23481 INVX1_LOC_185/A NOR2X1_LOC_109/Y 0.03fF
C23482 INVX1_LOC_34/A NOR2X1_LOC_736/Y 0.04fF
C23483 NAND2X1_LOC_454/Y INVX1_LOC_29/A 0.07fF
C23484 INVX1_LOC_5/A NOR2X1_LOC_641/Y 0.01fF
C23485 INVX1_LOC_208/A NOR2X1_LOC_665/A 0.45fF
C23486 NAND2X1_LOC_773/Y INVX1_LOC_117/A 0.01fF
C23487 INVX1_LOC_35/A NOR2X1_LOC_862/B 0.23fF
C23488 INVX1_LOC_64/A INVX1_LOC_117/Y 0.04fF
C23489 NOR2X1_LOC_186/Y INVX1_LOC_118/A 0.24fF
C23490 NOR2X1_LOC_244/a_36_216# INVX1_LOC_89/A 0.00fF
C23491 INVX1_LOC_215/A INVX1_LOC_22/A 0.15fF
C23492 INVX1_LOC_23/A NOR2X1_LOC_649/B 0.08fF
C23493 NAND2X1_LOC_550/A NAND2X1_LOC_242/a_36_24# 0.01fF
C23494 NOR2X1_LOC_419/Y NOR2X1_LOC_188/A 0.03fF
C23495 NOR2X1_LOC_570/A NOR2X1_LOC_570/Y 0.16fF
C23496 INVX1_LOC_181/Y NOR2X1_LOC_183/a_36_216# -0.00fF
C23497 NOR2X1_LOC_449/A NAND2X1_LOC_74/B 0.06fF
C23498 INVX1_LOC_23/A INVX1_LOC_3/A 0.09fF
C23499 NAND2X1_LOC_471/Y INVX1_LOC_42/A 0.01fF
C23500 NAND2X1_LOC_350/A NAND2X1_LOC_453/A 1.74fF
C23501 INVX1_LOC_103/A NOR2X1_LOC_506/a_36_216# 0.00fF
C23502 NOR2X1_LOC_142/Y INVX1_LOC_75/A 0.50fF
C23503 NOR2X1_LOC_419/Y NOR2X1_LOC_548/B 0.02fF
C23504 INVX1_LOC_129/A INVX1_LOC_63/A 0.01fF
C23505 NOR2X1_LOC_716/B NOR2X1_LOC_188/A 0.10fF
C23506 NOR2X1_LOC_168/B NOR2X1_LOC_356/A 0.00fF
C23507 NAND2X1_LOC_573/Y INVX1_LOC_118/A 0.17fF
C23508 INVX1_LOC_124/A NAND2X1_LOC_123/Y 0.06fF
C23509 NAND2X1_LOC_500/Y INVX1_LOC_20/A 0.11fF
C23510 NOR2X1_LOC_716/B NOR2X1_LOC_548/B 0.10fF
C23511 INVX1_LOC_1/A NOR2X1_LOC_709/B 0.04fF
C23512 INVX1_LOC_13/A NOR2X1_LOC_128/B 0.12fF
C23513 INVX1_LOC_88/Y NOR2X1_LOC_74/A 0.08fF
C23514 NOR2X1_LOC_220/A NOR2X1_LOC_180/B 0.96fF
C23515 INVX1_LOC_1/A NOR2X1_LOC_209/B 0.02fF
C23516 NOR2X1_LOC_441/Y NOR2X1_LOC_65/a_36_216# 0.02fF
C23517 NOR2X1_LOC_703/Y NOR2X1_LOC_551/B 0.29fF
C23518 NOR2X1_LOC_773/Y NOR2X1_LOC_153/a_36_216# 0.00fF
C23519 NOR2X1_LOC_92/Y INVX1_LOC_92/A 0.07fF
C23520 INVX1_LOC_87/A INVX1_LOC_4/A 0.10fF
C23521 NOR2X1_LOC_724/Y NOR2X1_LOC_687/Y 0.06fF
C23522 NOR2X1_LOC_655/B INVX1_LOC_75/A 0.99fF
C23523 NOR2X1_LOC_52/B NOR2X1_LOC_167/Y 0.03fF
C23524 NOR2X1_LOC_354/B VDD 0.50fF
C23525 NOR2X1_LOC_276/Y NOR2X1_LOC_331/B 0.12fF
C23526 INVX1_LOC_31/A NOR2X1_LOC_536/A 0.39fF
C23527 INVX1_LOC_49/A NAND2X1_LOC_642/Y 0.29fF
C23528 NOR2X1_LOC_34/A NAND2X1_LOC_574/A 0.06fF
C23529 INVX1_LOC_271/A INVX1_LOC_290/Y 0.00fF
C23530 NAND2X1_LOC_198/B NAND2X1_LOC_211/Y 0.10fF
C23531 NOR2X1_LOC_849/A INVX1_LOC_63/A 0.03fF
C23532 INVX1_LOC_90/A NAND2X1_LOC_319/A 0.74fF
C23533 NOR2X1_LOC_624/A NOR2X1_LOC_78/A 0.00fF
C23534 INVX1_LOC_47/Y NOR2X1_LOC_383/B 0.07fF
C23535 NOR2X1_LOC_720/B NAND2X1_LOC_490/a_36_24# 0.01fF
C23536 VDD INVX1_LOC_309/Y 0.27fF
C23537 INVX1_LOC_298/Y NAND2X1_LOC_454/Y 0.07fF
C23538 NOR2X1_LOC_315/Y INVX1_LOC_91/A 0.10fF
C23539 NAND2X1_LOC_53/Y NOR2X1_LOC_155/A 0.03fF
C23540 NAND2X1_LOC_35/Y INVX1_LOC_12/A 0.10fF
C23541 NOR2X1_LOC_433/A INVX1_LOC_76/A 0.38fF
C23542 NOR2X1_LOC_78/B INVX1_LOC_206/Y 0.03fF
C23543 INVX1_LOC_110/Y NOR2X1_LOC_61/Y 0.08fF
C23544 INVX1_LOC_31/A NOR2X1_LOC_655/Y 0.04fF
C23545 NOR2X1_LOC_643/A NAND2X1_LOC_574/A 0.04fF
C23546 NOR2X1_LOC_859/A NOR2X1_LOC_865/A 0.13fF
C23547 INVX1_LOC_170/A INVX1_LOC_118/A 0.07fF
C23548 NAND2X1_LOC_332/Y INVX1_LOC_147/Y 0.00fF
C23549 INVX1_LOC_136/A NOR2X1_LOC_331/B 0.17fF
C23550 NOR2X1_LOC_593/Y INVX1_LOC_76/A 0.02fF
C23551 NOR2X1_LOC_91/Y NAND2X1_LOC_848/A 0.71fF
C23552 NOR2X1_LOC_160/B NAND2X1_LOC_238/a_36_24# 0.01fF
C23553 NOR2X1_LOC_637/B INVX1_LOC_37/A 0.44fF
C23554 NOR2X1_LOC_569/A NOR2X1_LOC_548/Y 0.11fF
C23555 NOR2X1_LOC_395/Y NAND2X1_LOC_402/B 0.05fF
C23556 INVX1_LOC_2/A NAND2X1_LOC_642/Y 0.01fF
C23557 INVX1_LOC_151/A INVX1_LOC_76/A 0.01fF
C23558 INVX1_LOC_286/A INVX1_LOC_22/A 0.18fF
C23559 INVX1_LOC_93/A INVX1_LOC_102/A 0.14fF
C23560 NAND2X1_LOC_571/Y INVX1_LOC_12/A 0.07fF
C23561 INVX1_LOC_58/A INVX1_LOC_271/Y 0.10fF
C23562 NAND2X1_LOC_139/A D_INPUT_3 0.05fF
C23563 INVX1_LOC_144/A INVX1_LOC_10/A 0.19fF
C23564 NOR2X1_LOC_78/B NOR2X1_LOC_600/Y 0.12fF
C23565 NAND2X1_LOC_656/Y NOR2X1_LOC_74/A 0.07fF
C23566 NAND2X1_LOC_180/a_36_24# INVX1_LOC_20/A 0.01fF
C23567 NOR2X1_LOC_226/A NAND2X1_LOC_642/Y 0.36fF
C23568 NOR2X1_LOC_52/B INVX1_LOC_76/A 0.41fF
C23569 INVX1_LOC_93/Y NAND2X1_LOC_850/Y 0.03fF
C23570 NAND2X1_LOC_787/B NOR2X1_LOC_494/a_36_216# 0.01fF
C23571 NAND2X1_LOC_543/Y NOR2X1_LOC_528/Y 0.01fF
C23572 NOR2X1_LOC_788/B NOR2X1_LOC_567/B 0.14fF
C23573 NAND2X1_LOC_838/Y INVX1_LOC_76/A 0.09fF
C23574 INVX1_LOC_18/A NAND2X1_LOC_243/Y 0.07fF
C23575 NAND2X1_LOC_182/A INVX1_LOC_46/A 0.03fF
C23576 NOR2X1_LOC_355/A INPUT_0 0.03fF
C23577 INVX1_LOC_104/A INVX1_LOC_46/A 0.10fF
C23578 NOR2X1_LOC_495/Y INVX1_LOC_38/A 0.04fF
C23579 NAND2X1_LOC_702/a_36_24# INVX1_LOC_32/A 0.00fF
C23580 INVX1_LOC_249/Y INVX1_LOC_139/Y 0.01fF
C23581 INVX1_LOC_314/Y INVX1_LOC_9/A 0.13fF
C23582 NOR2X1_LOC_636/B INVX1_LOC_262/Y 0.06fF
C23583 INVX1_LOC_31/A NOR2X1_LOC_649/B 0.62fF
C23584 NAND2X1_LOC_231/Y INVX1_LOC_126/A 0.13fF
C23585 INVX1_LOC_17/A INVX1_LOC_125/A 0.07fF
C23586 INVX1_LOC_50/Y INVX1_LOC_15/A 0.38fF
C23587 INVX1_LOC_136/A NOR2X1_LOC_592/B 0.06fF
C23588 INVX1_LOC_31/A INVX1_LOC_3/A 0.14fF
C23589 NAND2X1_LOC_361/Y INVX1_LOC_38/A 0.07fF
C23590 INVX1_LOC_34/A NOR2X1_LOC_694/Y 0.03fF
C23591 INVX1_LOC_313/Y INVX1_LOC_67/Y 0.17fF
C23592 NOR2X1_LOC_803/A INVX1_LOC_75/A 0.19fF
C23593 INVX1_LOC_63/Y INVX1_LOC_281/Y 0.05fF
C23594 INVX1_LOC_182/A NOR2X1_LOC_439/B 0.02fF
C23595 INVX1_LOC_24/A NOR2X1_LOC_99/Y 0.21fF
C23596 NOR2X1_LOC_644/Y INVX1_LOC_14/Y 0.11fF
C23597 INVX1_LOC_134/Y VDD 0.62fF
C23598 NAND2X1_LOC_79/Y NOR2X1_LOC_78/Y 0.08fF
C23599 NOR2X1_LOC_376/a_36_216# NAND2X1_LOC_93/B 0.00fF
C23600 INVX1_LOC_182/A INVX1_LOC_75/A 0.07fF
C23601 INVX1_LOC_290/A INVX1_LOC_187/A 0.00fF
C23602 INVX1_LOC_83/A INVX1_LOC_86/Y 1.11fF
C23603 INVX1_LOC_31/A NOR2X1_LOC_814/a_36_216# 0.00fF
C23604 NOR2X1_LOC_577/Y INVX1_LOC_54/A 0.15fF
C23605 INVX1_LOC_59/A INVX1_LOC_3/Y 0.02fF
C23606 NAND2X1_LOC_89/a_36_24# NOR2X1_LOC_243/B 0.01fF
C23607 INVX1_LOC_72/A INVX1_LOC_285/A 0.24fF
C23608 NAND2X1_LOC_784/A NOR2X1_LOC_654/A 0.04fF
C23609 NAND2X1_LOC_641/a_36_24# NAND2X1_LOC_850/Y 0.01fF
C23610 NAND2X1_LOC_231/Y NOR2X1_LOC_111/A 0.15fF
C23611 NOR2X1_LOC_372/a_36_216# NAND2X1_LOC_489/Y 0.00fF
C23612 INVX1_LOC_21/A NOR2X1_LOC_227/A 0.01fF
C23613 NOR2X1_LOC_376/a_36_216# NAND2X1_LOC_425/Y 0.01fF
C23614 INVX1_LOC_94/A NOR2X1_LOC_445/B -0.01fF
C23615 INVX1_LOC_72/A NOR2X1_LOC_814/A 0.03fF
C23616 NAND2X1_LOC_493/a_36_24# INVX1_LOC_20/A 0.01fF
C23617 NAND2X1_LOC_721/A NAND2X1_LOC_850/Y 0.02fF
C23618 NOR2X1_LOC_219/Y NAND2X1_LOC_211/Y 0.01fF
C23619 NOR2X1_LOC_639/B NOR2X1_LOC_635/B 0.03fF
C23620 INVX1_LOC_191/Y NAND2X1_LOC_639/A 0.02fF
C23621 INVX1_LOC_263/A INVX1_LOC_46/A 0.07fF
C23622 INVX1_LOC_225/A INVX1_LOC_118/A 0.04fF
C23623 NOR2X1_LOC_278/Y NOR2X1_LOC_652/Y 0.07fF
C23624 INVX1_LOC_303/A NOR2X1_LOC_197/B 0.09fF
C23625 INVX1_LOC_241/A VDD -0.00fF
C23626 INVX1_LOC_71/A NOR2X1_LOC_117/a_36_216# 0.00fF
C23627 INVX1_LOC_41/A INVX1_LOC_92/A 0.03fF
C23628 NOR2X1_LOC_629/a_36_216# NOR2X1_LOC_629/Y 0.02fF
C23629 NOR2X1_LOC_309/Y INVX1_LOC_185/A 0.01fF
C23630 INVX1_LOC_230/Y INVX1_LOC_42/A 0.83fF
C23631 INVX1_LOC_16/A INVX1_LOC_12/Y 0.11fF
C23632 INVX1_LOC_41/Y INVX1_LOC_63/A 0.01fF
C23633 INPUT_1 NAND2X1_LOC_642/Y 0.09fF
C23634 NAND2X1_LOC_391/Y NAND2X1_LOC_99/A 0.03fF
C23635 NOR2X1_LOC_395/a_36_216# NOR2X1_LOC_396/Y 0.00fF
C23636 INVX1_LOC_306/A INVX1_LOC_20/A 0.07fF
C23637 NOR2X1_LOC_778/B INVX1_LOC_9/A 0.13fF
C23638 INVX1_LOC_145/Y NAND2X1_LOC_211/Y 0.03fF
C23639 NOR2X1_LOC_82/A INVX1_LOC_4/A 0.04fF
C23640 NOR2X1_LOC_298/Y VDD 5.69fF
C23641 NOR2X1_LOC_135/Y NOR2X1_LOC_269/Y 0.04fF
C23642 NAND2X1_LOC_352/B INVX1_LOC_32/A 0.10fF
C23643 NOR2X1_LOC_723/a_36_216# INVX1_LOC_12/A 0.00fF
C23644 NOR2X1_LOC_68/A INVX1_LOC_29/A 1.54fF
C23645 INVX1_LOC_8/A NOR2X1_LOC_49/a_36_216# 0.01fF
C23646 NOR2X1_LOC_74/A INVX1_LOC_78/Y 0.03fF
C23647 INVX1_LOC_6/A INVX1_LOC_126/Y 0.11fF
C23648 NOR2X1_LOC_593/a_36_216# INVX1_LOC_179/A 0.00fF
C23649 NAND2X1_LOC_852/Y INVX1_LOC_118/A 0.05fF
C23650 INVX1_LOC_181/Y NAND2X1_LOC_81/B 0.07fF
C23651 INVX1_LOC_286/A INVX1_LOC_100/A 0.07fF
C23652 INVX1_LOC_279/A INVX1_LOC_117/A 0.07fF
C23653 INVX1_LOC_24/A INVX1_LOC_272/A 0.07fF
C23654 INVX1_LOC_14/A INVX1_LOC_23/Y 0.20fF
C23655 NAND2X1_LOC_859/Y NOR2X1_LOC_536/A 0.08fF
C23656 INVX1_LOC_75/A NOR2X1_LOC_502/a_36_216# 0.00fF
C23657 INVX1_LOC_108/Y INVX1_LOC_50/Y 0.18fF
C23658 INVX1_LOC_94/A INVX1_LOC_12/A 0.03fF
C23659 INVX1_LOC_49/A NOR2X1_LOC_48/Y 0.03fF
C23660 NOR2X1_LOC_758/Y INVX1_LOC_63/A 0.01fF
C23661 NOR2X1_LOC_315/Y NOR2X1_LOC_179/Y 0.04fF
C23662 INVX1_LOC_58/A INVX1_LOC_59/A 0.25fF
C23663 INVX1_LOC_22/A INVX1_LOC_54/A 0.24fF
C23664 NOR2X1_LOC_454/Y INVX1_LOC_105/Y 0.02fF
C23665 NOR2X1_LOC_112/Y INVX1_LOC_36/Y 0.03fF
C23666 NOR2X1_LOC_6/B INVX1_LOC_84/A 0.08fF
C23667 NOR2X1_LOC_545/A INVX1_LOC_29/A 0.01fF
C23668 INVX1_LOC_132/A NAND2X1_LOC_63/Y 0.02fF
C23669 INVX1_LOC_45/A NAND2X1_LOC_647/B 0.02fF
C23670 NOR2X1_LOC_348/Y INVX1_LOC_23/A 0.67fF
C23671 NOR2X1_LOC_315/Y INVX1_LOC_203/A 0.01fF
C23672 NOR2X1_LOC_92/Y INVX1_LOC_53/A 0.07fF
C23673 INVX1_LOC_95/A INVX1_LOC_100/A 0.01fF
C23674 NOR2X1_LOC_329/B NOR2X1_LOC_139/a_36_216# 0.00fF
C23675 INVX1_LOC_28/A INVX1_LOC_12/Y 0.10fF
C23676 INVX1_LOC_24/Y INVX1_LOC_53/A 0.05fF
C23677 NAND2X1_LOC_866/B NOR2X1_LOC_536/A 0.07fF
C23678 INVX1_LOC_18/A INVX1_LOC_21/Y 0.04fF
C23679 INPUT_0 INVX1_LOC_126/A 0.04fF
C23680 NOR2X1_LOC_537/Y NOR2X1_LOC_814/A 0.07fF
C23681 NOR2X1_LOC_87/Y NAND2X1_LOC_206/Y 0.04fF
C23682 NAND2X1_LOC_338/B NOR2X1_LOC_814/A 0.07fF
C23683 NOR2X1_LOC_577/Y NOR2X1_LOC_48/B 0.09fF
C23684 NOR2X1_LOC_802/A INVX1_LOC_19/A 0.34fF
C23685 INPUT_1 NOR2X1_LOC_271/Y 0.04fF
C23686 INVX1_LOC_289/Y INVX1_LOC_64/A 0.03fF
C23687 INVX1_LOC_256/A INVX1_LOC_23/A 0.80fF
C23688 NAND2X1_LOC_573/a_36_24# INVX1_LOC_32/A 0.06fF
C23689 INVX1_LOC_121/A INVX1_LOC_92/A 0.03fF
C23690 NAND2X1_LOC_807/Y NOR2X1_LOC_536/A 0.45fF
C23691 NAND2X1_LOC_323/B NOR2X1_LOC_814/A 0.01fF
C23692 NOR2X1_LOC_488/Y INVX1_LOC_119/Y 0.03fF
C23693 INVX1_LOC_57/Y NOR2X1_LOC_693/a_36_216# 0.00fF
C23694 NAND2X1_LOC_53/Y NOR2X1_LOC_598/B 0.10fF
C23695 INVX1_LOC_71/A NAND2X1_LOC_647/B 0.03fF
C23696 INVX1_LOC_10/A NOR2X1_LOC_155/A 0.09fF
C23697 NOR2X1_LOC_478/A INVX1_LOC_204/A 0.20fF
C23698 NOR2X1_LOC_142/Y INVX1_LOC_283/A 0.00fF
C23699 INPUT_0 NOR2X1_LOC_111/A 0.05fF
C23700 INVX1_LOC_298/Y NOR2X1_LOC_68/A 0.02fF
C23701 INVX1_LOC_64/A NOR2X1_LOC_82/A 0.02fF
C23702 NOR2X1_LOC_454/Y INVX1_LOC_27/A 0.59fF
C23703 NAND2X1_LOC_740/Y NOR2X1_LOC_15/Y 0.01fF
C23704 NOR2X1_LOC_609/a_36_216# NOR2X1_LOC_334/Y 0.01fF
C23705 NAND2X1_LOC_123/Y INVX1_LOC_9/A 0.02fF
C23706 INVX1_LOC_206/Y INVX1_LOC_46/A 0.03fF
C23707 INVX1_LOC_30/Y INVX1_LOC_84/A 0.07fF
C23708 NOR2X1_LOC_178/Y INVX1_LOC_11/A 0.77fF
C23709 INVX1_LOC_96/Y INVX1_LOC_109/Y 0.18fF
C23710 INVX1_LOC_36/A INVX1_LOC_270/Y 0.24fF
C23711 NOR2X1_LOC_52/B INVX1_LOC_127/Y 0.08fF
C23712 NAND2X1_LOC_354/Y NOR2X1_LOC_677/Y 0.00fF
C23713 NAND2X1_LOC_468/B NOR2X1_LOC_56/Y 0.03fF
C23714 NOR2X1_LOC_122/Y INVX1_LOC_92/A 0.05fF
C23715 INVX1_LOC_204/A NOR2X1_LOC_68/A 0.03fF
C23716 NAND2X1_LOC_357/B INVX1_LOC_32/A 0.12fF
C23717 NOR2X1_LOC_836/B VDD -0.00fF
C23718 NAND2X1_LOC_66/a_36_24# INVX1_LOC_284/A 0.00fF
C23719 NOR2X1_LOC_823/Y NAND2X1_LOC_836/Y 0.00fF
C23720 NOR2X1_LOC_254/A INVX1_LOC_5/A 0.13fF
C23721 NOR2X1_LOC_139/Y VDD 0.36fF
C23722 NOR2X1_LOC_798/A NOR2X1_LOC_288/a_36_216# 0.00fF
C23723 INVX1_LOC_6/A NOR2X1_LOC_536/A 0.10fF
C23724 INVX1_LOC_289/Y NAND2X1_LOC_704/a_36_24# 0.06fF
C23725 INVX1_LOC_199/A INVX1_LOC_76/A 0.03fF
C23726 NOR2X1_LOC_619/A NAND2X1_LOC_207/B 0.05fF
C23727 INVX1_LOC_269/A INVX1_LOC_48/Y 0.10fF
C23728 NAND2X1_LOC_35/Y NAND2X1_LOC_733/Y 0.42fF
C23729 INVX1_LOC_244/Y INVX1_LOC_296/A 0.02fF
C23730 NOR2X1_LOC_570/Y INVX1_LOC_29/A 0.03fF
C23731 NAND2X1_LOC_800/A NAND2X1_LOC_655/A 0.04fF
C23732 INPUT_0 INVX1_LOC_127/A 0.01fF
C23733 NAND2X1_LOC_753/a_36_24# INVX1_LOC_223/A 0.00fF
C23734 INVX1_LOC_13/A NOR2X1_LOC_610/a_36_216# 0.00fF
C23735 VDD NAND2X1_LOC_468/B 0.01fF
C23736 VDD NOR2X1_LOC_683/Y 0.12fF
C23737 NOR2X1_LOC_459/B INVX1_LOC_175/A 0.05fF
C23738 INVX1_LOC_22/A NOR2X1_LOC_48/B 0.61fF
C23739 INVX1_LOC_77/A INVX1_LOC_271/A 0.07fF
C23740 NAND2X1_LOC_149/Y NOR2X1_LOC_160/B 0.07fF
C23741 D_INPUT_0 NAND2X1_LOC_82/Y 0.22fF
C23742 INVX1_LOC_147/A NOR2X1_LOC_58/Y 0.36fF
C23743 INVX1_LOC_64/A NAND2X1_LOC_514/Y 0.28fF
C23744 INVX1_LOC_17/A NAND2X1_LOC_538/Y 0.10fF
C23745 NAND2X1_LOC_35/Y INVX1_LOC_217/A 0.26fF
C23746 NAND2X1_LOC_787/A NOR2X1_LOC_238/Y 0.02fF
C23747 NOR2X1_LOC_130/A INVX1_LOC_272/A 0.07fF
C23748 NOR2X1_LOC_557/A INVX1_LOC_9/A 0.20fF
C23749 INVX1_LOC_135/A NAND2X1_LOC_74/B 0.02fF
C23750 INVX1_LOC_50/A NOR2X1_LOC_172/Y 0.01fF
C23751 INVX1_LOC_6/A NAND2X1_LOC_93/B 0.15fF
C23752 NAND2X1_LOC_807/Y NOR2X1_LOC_661/A 0.04fF
C23753 INVX1_LOC_135/A NAND2X1_LOC_207/Y 0.05fF
C23754 NOR2X1_LOC_665/A NAND2X1_LOC_791/a_36_24# 0.00fF
C23755 NAND2X1_LOC_555/Y NAND2X1_LOC_218/A 0.00fF
C23756 INVX1_LOC_17/A NOR2X1_LOC_250/A 0.02fF
C23757 NAND2X1_LOC_555/Y NOR2X1_LOC_140/A 0.07fF
C23758 INVX1_LOC_103/A INVX1_LOC_174/A 0.15fF
C23759 NAND2X1_LOC_642/Y INVX1_LOC_118/A 0.07fF
C23760 NAND2X1_LOC_849/A NAND2X1_LOC_489/Y 0.02fF
C23761 INVX1_LOC_58/A NOR2X1_LOC_144/Y 0.27fF
C23762 INVX1_LOC_41/A INVX1_LOC_53/A 8.25fF
C23763 NOR2X1_LOC_445/a_36_216# NOR2X1_LOC_457/A 0.00fF
C23764 NOR2X1_LOC_82/A INVX1_LOC_43/Y 0.05fF
C23765 NOR2X1_LOC_197/Y INVX1_LOC_19/A 0.01fF
C23766 INVX1_LOC_286/Y INVX1_LOC_88/A 0.00fF
C23767 NAND2X1_LOC_341/A INVX1_LOC_78/A 0.02fF
C23768 INVX1_LOC_188/A NOR2X1_LOC_457/A 0.06fF
C23769 NAND2X1_LOC_35/Y NAND2X1_LOC_787/B 0.17fF
C23770 NOR2X1_LOC_455/a_36_216# INVX1_LOC_53/A 0.01fF
C23771 INVX1_LOC_221/A NOR2X1_LOC_591/A 0.21fF
C23772 INVX1_LOC_6/A INVX1_LOC_3/A 0.05fF
C23773 NOR2X1_LOC_216/Y INVX1_LOC_272/A 0.03fF
C23774 INVX1_LOC_256/A INVX1_LOC_31/A 0.01fF
C23775 GATE_479 INVX1_LOC_78/A 0.03fF
C23776 INVX1_LOC_58/A NOR2X1_LOC_432/a_36_216# 0.00fF
C23777 INVX1_LOC_214/A NOR2X1_LOC_677/Y 0.00fF
C23778 INVX1_LOC_34/Y NAND2X1_LOC_205/A 0.76fF
C23779 NOR2X1_LOC_647/B INVX1_LOC_31/A 0.01fF
C23780 NAND2X1_LOC_477/A INVX1_LOC_53/A 0.01fF
C23781 NAND2X1_LOC_300/a_36_24# NOR2X1_LOC_109/Y 0.00fF
C23782 NAND2X1_LOC_182/A INVX1_LOC_233/A 0.04fF
C23783 NOR2X1_LOC_98/B INVX1_LOC_117/A 0.03fF
C23784 INVX1_LOC_27/A INVX1_LOC_77/A 0.30fF
C23785 NOR2X1_LOC_203/a_36_216# NOR2X1_LOC_388/Y 0.00fF
C23786 NAND2X1_LOC_451/Y NOR2X1_LOC_452/A 0.03fF
C23787 NOR2X1_LOC_612/a_36_216# INVX1_LOC_57/A 0.00fF
C23788 NOR2X1_LOC_647/Y NOR2X1_LOC_817/Y 0.09fF
C23789 INVX1_LOC_232/Y D_INPUT_1 0.31fF
C23790 INVX1_LOC_255/Y NOR2X1_LOC_647/A 0.02fF
C23791 INVX1_LOC_21/A NOR2X1_LOC_636/A 0.01fF
C23792 NOR2X1_LOC_178/Y NOR2X1_LOC_52/B 0.30fF
C23793 NOR2X1_LOC_256/Y INVX1_LOC_42/A 0.01fF
C23794 NAND2X1_LOC_803/B INVX1_LOC_72/A 0.03fF
C23795 INVX1_LOC_144/A INVX1_LOC_12/A 0.09fF
C23796 NOR2X1_LOC_561/a_36_216# NOR2X1_LOC_652/Y 0.11fF
C23797 NOR2X1_LOC_804/a_36_216# INVX1_LOC_292/Y 0.01fF
C23798 INVX1_LOC_41/A NOR2X1_LOC_242/A 0.07fF
C23799 NAND2X1_LOC_140/A NAND2X1_LOC_454/Y 0.01fF
C23800 NOR2X1_LOC_68/A NOR2X1_LOC_745/a_36_216# 0.00fF
C23801 NOR2X1_LOC_75/Y NOR2X1_LOC_194/a_36_216# 0.00fF
C23802 NOR2X1_LOC_83/Y INVX1_LOC_12/A 0.04fF
C23803 NAND2X1_LOC_363/B INVX1_LOC_196/A 0.01fF
C23804 D_INPUT_7 NOR2X1_LOC_22/a_36_216# -0.00fF
C23805 NOR2X1_LOC_667/Y INVX1_LOC_36/A 0.03fF
C23806 INVX1_LOC_163/A NOR2X1_LOC_474/A 0.12fF
C23807 INVX1_LOC_93/A INVX1_LOC_162/Y 0.02fF
C23808 NOR2X1_LOC_798/A INVX1_LOC_104/A 0.03fF
C23809 NOR2X1_LOC_590/A INVX1_LOC_72/A 0.03fF
C23810 NOR2X1_LOC_124/A INVX1_LOC_84/A 0.07fF
C23811 INVX1_LOC_1/Y INVX1_LOC_129/A -0.01fF
C23812 INVX1_LOC_256/A INVX1_LOC_111/A 0.01fF
C23813 INVX1_LOC_50/A NOR2X1_LOC_512/a_36_216# 0.02fF
C23814 NOR2X1_LOC_658/Y NOR2X1_LOC_657/Y 0.01fF
C23815 INVX1_LOC_118/A NOR2X1_LOC_271/Y 0.01fF
C23816 INVX1_LOC_258/Y INVX1_LOC_240/A 0.01fF
C23817 INVX1_LOC_64/A INVX1_LOC_278/Y 0.15fF
C23818 NOR2X1_LOC_246/A NOR2X1_LOC_282/Y 0.01fF
C23819 INVX1_LOC_226/Y INVX1_LOC_51/A 0.09fF
C23820 VDD NAND2X1_LOC_141/Y 0.80fF
C23821 NOR2X1_LOC_689/Y INVX1_LOC_10/A 0.37fF
C23822 NOR2X1_LOC_405/A INVX1_LOC_49/Y 0.10fF
C23823 NOR2X1_LOC_810/A INVX1_LOC_23/A 0.03fF
C23824 INVX1_LOC_25/A NOR2X1_LOC_391/A 0.04fF
C23825 INVX1_LOC_58/A INVX1_LOC_279/A 0.17fF
C23826 NOR2X1_LOC_536/A INVX1_LOC_131/Y 0.01fF
C23827 INVX1_LOC_256/Y INVX1_LOC_306/Y 0.01fF
C23828 INVX1_LOC_229/A NAND2X1_LOC_736/B 0.04fF
C23829 NOR2X1_LOC_242/A INVX1_LOC_64/Y 0.03fF
C23830 NOR2X1_LOC_441/Y NOR2X1_LOC_351/a_36_216# 0.00fF
C23831 NOR2X1_LOC_552/A NAND2X1_LOC_74/B 0.08fF
C23832 NAND2X1_LOC_63/Y NAND2X1_LOC_642/Y 0.02fF
C23833 VDD NOR2X1_LOC_66/Y 0.10fF
C23834 NAND2X1_LOC_721/B NOR2X1_LOC_68/A 0.14fF
C23835 VDD NOR2X1_LOC_820/B -0.00fF
C23836 NAND2X1_LOC_149/Y INVX1_LOC_189/A -0.08fF
C23837 INVX1_LOC_173/Y INVX1_LOC_173/A 0.01fF
C23838 INVX1_LOC_178/A INVX1_LOC_144/Y 0.01fF
C23839 INVX1_LOC_50/A INVX1_LOC_90/A 3.08fF
C23840 NAND2X1_LOC_739/B NAND2X1_LOC_741/B 0.01fF
C23841 INVX1_LOC_247/Y NOR2X1_LOC_68/A 0.36fF
C23842 NOR2X1_LOC_238/Y INVX1_LOC_30/A 0.03fF
C23843 INVX1_LOC_101/Y INVX1_LOC_177/A 0.04fF
C23844 INVX1_LOC_2/Y INVX1_LOC_19/A 0.03fF
C23845 NOR2X1_LOC_441/Y NOR2X1_LOC_577/Y 0.07fF
C23846 NOR2X1_LOC_92/Y NOR2X1_LOC_78/B 0.07fF
C23847 INVX1_LOC_223/A NOR2X1_LOC_303/Y 0.03fF
C23848 NAND2X1_LOC_725/A INVX1_LOC_10/A 0.14fF
C23849 INVX1_LOC_96/A INVX1_LOC_15/A 0.16fF
C23850 INVX1_LOC_21/A INVX1_LOC_56/Y 0.02fF
C23851 INVX1_LOC_135/A NOR2X1_LOC_660/Y 0.03fF
C23852 INVX1_LOC_269/A INVX1_LOC_216/A 0.14fF
C23853 NAND2X1_LOC_725/B INVX1_LOC_280/Y 0.03fF
C23854 NOR2X1_LOC_32/B INVX1_LOC_89/A 0.07fF
C23855 INVX1_LOC_24/Y NOR2X1_LOC_78/B 0.00fF
C23856 NAND2X1_LOC_563/A INVX1_LOC_48/Y 0.01fF
C23857 INVX1_LOC_6/A NAND2X1_LOC_470/B 0.03fF
C23858 NOR2X1_LOC_433/Y INVX1_LOC_179/A 0.01fF
C23859 NOR2X1_LOC_75/Y NOR2X1_LOC_300/Y 0.01fF
C23860 NOR2X1_LOC_468/Y NAND2X1_LOC_181/Y 0.03fF
C23861 NAND2X1_LOC_848/A NOR2X1_LOC_661/a_36_216# 0.12fF
C23862 INVX1_LOC_227/A NOR2X1_LOC_674/Y 0.18fF
C23863 NOR2X1_LOC_607/A INVX1_LOC_45/Y 0.07fF
C23864 NOR2X1_LOC_760/a_36_216# INVX1_LOC_177/A 0.00fF
C23865 INVX1_LOC_58/A INVX1_LOC_182/Y 0.01fF
C23866 INVX1_LOC_248/A NOR2X1_LOC_533/Y 0.14fF
C23867 INVX1_LOC_280/A INVX1_LOC_293/Y 0.01fF
C23868 NOR2X1_LOC_74/A NOR2X1_LOC_727/B 0.03fF
C23869 NAND2X1_LOC_717/Y NAND2X1_LOC_550/A 0.28fF
C23870 NAND2X1_LOC_171/a_36_24# NOR2X1_LOC_175/A 0.00fF
C23871 NOR2X1_LOC_82/A NAND2X1_LOC_850/Y 0.07fF
C23872 NOR2X1_LOC_286/a_36_216# INVX1_LOC_89/A 0.00fF
C23873 NOR2X1_LOC_813/Y NAND2X1_LOC_74/B 0.07fF
C23874 INVX1_LOC_14/A INVX1_LOC_232/A 0.18fF
C23875 INVX1_LOC_103/A NOR2X1_LOC_131/Y 0.01fF
C23876 NAND2X1_LOC_740/Y NOR2X1_LOC_576/B 0.03fF
C23877 INVX1_LOC_136/A NOR2X1_LOC_388/Y 0.01fF
C23878 INVX1_LOC_264/Y INVX1_LOC_273/A 0.02fF
C23879 NOR2X1_LOC_527/Y NOR2X1_LOC_654/A 0.06fF
C23880 NOR2X1_LOC_468/Y NAND2X1_LOC_390/A 0.02fF
C23881 INVX1_LOC_239/A NAND2X1_LOC_462/B 0.02fF
C23882 NAND2X1_LOC_658/a_36_24# INVX1_LOC_15/A 0.00fF
C23883 INVX1_LOC_185/A NOR2X1_LOC_654/a_36_216# 0.00fF
C23884 INVX1_LOC_34/A NAND2X1_LOC_364/A 0.03fF
C23885 NOR2X1_LOC_590/A NOR2X1_LOC_537/Y 0.03fF
C23886 NOR2X1_LOC_590/A NAND2X1_LOC_338/B 0.10fF
C23887 INVX1_LOC_185/A INVX1_LOC_63/A 0.03fF
C23888 INVX1_LOC_58/A NAND2X1_LOC_858/B 0.07fF
C23889 NOR2X1_LOC_383/Y INVX1_LOC_14/A 0.00fF
C23890 INVX1_LOC_280/A NAND2X1_LOC_74/B 0.14fF
C23891 INVX1_LOC_186/Y INVX1_LOC_54/A 0.08fF
C23892 NOR2X1_LOC_276/Y NOR2X1_LOC_366/B 0.01fF
C23893 NOR2X1_LOC_177/Y NOR2X1_LOC_662/A -0.00fF
C23894 INVX1_LOC_103/A NOR2X1_LOC_589/A 0.06fF
C23895 NOR2X1_LOC_590/A NAND2X1_LOC_323/B 0.03fF
C23896 NOR2X1_LOC_92/Y INVX1_LOC_83/A 0.10fF
C23897 NAND2X1_LOC_578/B NAND2X1_LOC_577/A 0.30fF
C23898 NAND2X1_LOC_9/Y NOR2X1_LOC_394/a_36_216# 0.00fF
C23899 INVX1_LOC_91/A NAND2X1_LOC_99/A 0.10fF
C23900 NAND2X1_LOC_550/A INVX1_LOC_16/A 0.07fF
C23901 VDD NOR2X1_LOC_685/Y 0.14fF
C23902 NOR2X1_LOC_74/A NOR2X1_LOC_717/A 0.61fF
C23903 NOR2X1_LOC_274/Y NOR2X1_LOC_593/Y 0.02fF
C23904 D_INPUT_0 NAND2X1_LOC_780/Y 0.01fF
C23905 INVX1_LOC_45/A NAND2X1_LOC_342/Y 0.05fF
C23906 INVX1_LOC_69/Y INVX1_LOC_23/A 0.01fF
C23907 NAND2X1_LOC_350/A INVX1_LOC_22/A 0.07fF
C23908 INVX1_LOC_307/Y INVX1_LOC_19/A 0.00fF
C23909 INVX1_LOC_24/Y INVX1_LOC_83/A 0.65fF
C23910 NOR2X1_LOC_160/B INVX1_LOC_16/A 0.10fF
C23911 INVX1_LOC_230/Y NAND2X1_LOC_859/B 0.00fF
C23912 NAND2X1_LOC_364/Y NAND2X1_LOC_367/A 0.10fF
C23913 NAND2X1_LOC_181/a_36_24# INVX1_LOC_43/Y 0.00fF
C23914 INVX1_LOC_30/A NOR2X1_LOC_769/a_36_216# 0.01fF
C23915 NOR2X1_LOC_655/B NOR2X1_LOC_274/B 0.07fF
C23916 NOR2X1_LOC_391/B NOR2X1_LOC_660/Y 0.03fF
C23917 NAND2X1_LOC_361/Y INVX1_LOC_33/A 0.07fF
C23918 INVX1_LOC_2/A NOR2X1_LOC_91/Y 0.03fF
C23919 NOR2X1_LOC_250/Y NAND2X1_LOC_656/Y 0.04fF
C23920 NOR2X1_LOC_142/Y NOR2X1_LOC_577/Y 0.10fF
C23921 NOR2X1_LOC_441/Y INVX1_LOC_22/A 0.05fF
C23922 NOR2X1_LOC_624/A INVX1_LOC_132/A 0.08fF
C23923 NOR2X1_LOC_523/A INVX1_LOC_120/A 0.03fF
C23924 INVX1_LOC_85/A NOR2X1_LOC_303/Y 0.02fF
C23925 NOR2X1_LOC_725/A INVX1_LOC_23/A 0.03fF
C23926 INVX1_LOC_17/A NOR2X1_LOC_106/A 0.01fF
C23927 NOR2X1_LOC_323/Y NOR2X1_LOC_406/A 0.01fF
C23928 NOR2X1_LOC_67/A NOR2X1_LOC_360/Y 0.07fF
C23929 NOR2X1_LOC_226/A NOR2X1_LOC_91/Y 0.23fF
C23930 NOR2X1_LOC_673/A NAND2X1_LOC_206/Y 0.07fF
C23931 INVX1_LOC_178/A NOR2X1_LOC_322/Y 0.28fF
C23932 INVX1_LOC_11/A NAND2X1_LOC_45/Y 0.03fF
C23933 INVX1_LOC_268/A INVX1_LOC_30/A 0.06fF
C23934 NOR2X1_LOC_781/Y INVX1_LOC_191/Y 0.00fF
C23935 INPUT_3 NOR2X1_LOC_128/B 0.01fF
C23936 INVX1_LOC_93/Y INVX1_LOC_129/A -0.03fF
C23937 INVX1_LOC_256/A INVX1_LOC_313/A 0.25fF
C23938 INVX1_LOC_12/A NOR2X1_LOC_155/A 0.14fF
C23939 NOR2X1_LOC_772/Y NOR2X1_LOC_773/a_36_216# 0.00fF
C23940 NAND2X1_LOC_342/Y INVX1_LOC_71/A 0.00fF
C23941 NOR2X1_LOC_272/Y INPUT_0 0.01fF
C23942 NAND2X1_LOC_714/a_36_24# INVX1_LOC_28/A 0.01fF
C23943 INVX1_LOC_312/Y NAND2X1_LOC_660/Y 0.01fF
C23944 INVX1_LOC_250/A NOR2X1_LOC_605/B 0.00fF
C23945 INVX1_LOC_232/Y D_INPUT_2 0.07fF
C23946 INVX1_LOC_27/A NAND2X1_LOC_832/Y 0.03fF
C23947 INVX1_LOC_90/A NAND2X1_LOC_227/Y 0.00fF
C23948 NAND2X1_LOC_860/A NOR2X1_LOC_80/a_36_216# 0.01fF
C23949 NOR2X1_LOC_479/B NOR2X1_LOC_480/A 0.01fF
C23950 NOR2X1_LOC_80/Y NOR2X1_LOC_536/A 0.28fF
C23951 INVX1_LOC_78/A INVX1_LOC_44/A 0.03fF
C23952 NAND2X1_LOC_569/a_36_24# INVX1_LOC_234/A 0.00fF
C23953 NOR2X1_LOC_456/Y INVX1_LOC_247/A 0.19fF
C23954 NOR2X1_LOC_598/B NOR2X1_LOC_799/B 0.01fF
C23955 INVX1_LOC_278/A NOR2X1_LOC_124/A 0.02fF
C23956 INVX1_LOC_243/Y INVX1_LOC_37/A 0.01fF
C23957 NOR2X1_LOC_703/B INVX1_LOC_220/Y 0.01fF
C23958 INVX1_LOC_227/A INVX1_LOC_72/A 0.07fF
C23959 INVX1_LOC_5/A NOR2X1_LOC_562/B 0.10fF
C23960 NOR2X1_LOC_111/Y INVX1_LOC_161/Y 0.04fF
C23961 NAND2X1_LOC_542/a_36_24# NOR2X1_LOC_45/B 0.01fF
C23962 NAND2X1_LOC_363/B INVX1_LOC_95/Y 0.01fF
C23963 NAND2X1_LOC_550/A INVX1_LOC_28/A 0.08fF
C23964 NOR2X1_LOC_681/Y INVX1_LOC_57/A 0.07fF
C23965 NOR2X1_LOC_15/Y NOR2X1_LOC_335/B 0.07fF
C23966 NAND2X1_LOC_84/Y INVX1_LOC_232/A 0.72fF
C23967 NOR2X1_LOC_590/A INVX1_LOC_313/Y 0.08fF
C23968 D_INPUT_0 INVX1_LOC_312/Y 0.09fF
C23969 NOR2X1_LOC_251/Y INVX1_LOC_77/A 0.04fF
C23970 NOR2X1_LOC_211/Y INVX1_LOC_93/Y 0.02fF
C23971 NOR2X1_LOC_160/B INVX1_LOC_28/A 0.07fF
C23972 NOR2X1_LOC_32/B NOR2X1_LOC_24/Y 0.02fF
C23973 INVX1_LOC_37/A INVX1_LOC_57/A 0.72fF
C23974 NAND2X1_LOC_338/B NAND2X1_LOC_518/a_36_24# 0.00fF
C23975 INVX1_LOC_41/A NOR2X1_LOC_78/B 0.07fF
C23976 NAND2X1_LOC_341/A NOR2X1_LOC_152/Y 0.01fF
C23977 INVX1_LOC_64/A INVX1_LOC_59/Y 0.05fF
C23978 NOR2X1_LOC_616/a_36_216# NOR2X1_LOC_413/Y 0.01fF
C23979 INVX1_LOC_136/A INVX1_LOC_135/A 0.10fF
C23980 INVX1_LOC_30/A NOR2X1_LOC_367/a_36_216# 0.00fF
C23981 NAND2X1_LOC_112/Y NOR2X1_LOC_106/Y 0.05fF
C23982 NAND2X1_LOC_361/Y INVX1_LOC_40/A 0.00fF
C23983 NAND2X1_LOC_228/a_36_24# INVX1_LOC_105/A 0.00fF
C23984 NOR2X1_LOC_510/Y NAND2X1_LOC_655/A 0.01fF
C23985 INVX1_LOC_83/A NOR2X1_LOC_798/a_36_216# 0.00fF
C23986 INVX1_LOC_47/A INVX1_LOC_30/A 1.01fF
C23987 INVX1_LOC_85/A NOR2X1_LOC_353/Y 0.01fF
C23988 INVX1_LOC_45/A NOR2X1_LOC_246/Y 0.06fF
C23989 NOR2X1_LOC_80/Y NAND2X1_LOC_93/B 0.12fF
C23990 INVX1_LOC_64/A INVX1_LOC_176/A 0.03fF
C23991 INVX1_LOC_259/Y INVX1_LOC_139/Y 0.55fF
C23992 NOR2X1_LOC_655/B NOR2X1_LOC_348/B 0.01fF
C23993 NOR2X1_LOC_536/A INVX1_LOC_270/A 0.10fF
C23994 NAND2X1_LOC_374/Y NOR2X1_LOC_315/Y 0.00fF
C23995 GATE_479 INVX1_LOC_113/Y 0.01fF
C23996 NOR2X1_LOC_791/Y INVX1_LOC_95/Y 0.03fF
C23997 NAND2X1_LOC_508/A NAND2X1_LOC_510/A 0.05fF
C23998 NOR2X1_LOC_78/B NAND2X1_LOC_477/A 1.45fF
C23999 INVX1_LOC_50/A INVX1_LOC_38/A 4.09fF
C24000 NOR2X1_LOC_510/Y NAND2X1_LOC_468/B 0.07fF
C24001 NAND2X1_LOC_777/a_36_24# INVX1_LOC_33/Y 0.00fF
C24002 NOR2X1_LOC_142/Y INVX1_LOC_22/A 0.07fF
C24003 INVX1_LOC_93/Y NOR2X1_LOC_440/B 0.01fF
C24004 NOR2X1_LOC_78/B NOR2X1_LOC_398/Y 0.04fF
C24005 NAND2X1_LOC_348/A INVX1_LOC_61/Y 0.01fF
C24006 INVX1_LOC_136/A NOR2X1_LOC_248/a_36_216# 0.00fF
C24007 NOR2X1_LOC_91/Y INPUT_1 0.65fF
C24008 NOR2X1_LOC_711/A NOR2X1_LOC_307/A 0.31fF
C24009 INVX1_LOC_256/A INVX1_LOC_6/A 0.14fF
C24010 NOR2X1_LOC_772/B VDD 0.74fF
C24011 NOR2X1_LOC_88/Y INVX1_LOC_273/A 0.03fF
C24012 NOR2X1_LOC_241/a_36_216# INVX1_LOC_143/Y 0.00fF
C24013 INVX1_LOC_136/A NOR2X1_LOC_490/Y 0.03fF
C24014 NAND2X1_LOC_563/A NOR2X1_LOC_84/Y 0.02fF
C24015 NAND2X1_LOC_561/B NOR2X1_LOC_45/B 0.07fF
C24016 NOR2X1_LOC_781/A INVX1_LOC_63/Y 0.01fF
C24017 INVX1_LOC_269/A INVX1_LOC_160/A 0.01fF
C24018 NOR2X1_LOC_78/B INVX1_LOC_64/Y 0.07fF
C24019 INVX1_LOC_34/A NOR2X1_LOC_86/A 0.16fF
C24020 INVX1_LOC_277/A NOR2X1_LOC_151/Y 0.01fF
C24021 NOR2X1_LOC_297/A NOR2X1_LOC_673/A 0.01fF
C24022 INVX1_LOC_202/Y NOR2X1_LOC_678/A 0.01fF
C24023 INVX1_LOC_41/A NAND2X1_LOC_392/Y 0.02fF
C24024 NOR2X1_LOC_598/B INVX1_LOC_114/A 0.03fF
C24025 INVX1_LOC_145/Y INVX1_LOC_155/A 0.12fF
C24026 NOR2X1_LOC_266/a_36_216# INVX1_LOC_102/Y -0.01fF
C24027 NOR2X1_LOC_599/Y NOR2X1_LOC_387/A 0.18fF
C24028 NOR2X1_LOC_742/A INVX1_LOC_142/A 0.06fF
C24029 NOR2X1_LOC_778/B INVX1_LOC_179/Y 0.01fF
C24030 INVX1_LOC_45/A INVX1_LOC_67/Y 0.00fF
C24031 NAND2X1_LOC_287/B NOR2X1_LOC_652/Y 0.03fF
C24032 INVX1_LOC_13/Y VDD 0.13fF
C24033 INVX1_LOC_90/A NAND2X1_LOC_845/a_36_24# 0.00fF
C24034 NOR2X1_LOC_92/Y NOR2X1_LOC_368/Y 0.08fF
C24035 INVX1_LOC_50/A NOR2X1_LOC_51/A 0.01fF
C24036 NOR2X1_LOC_761/Y INPUT_0 0.19fF
C24037 NAND2X1_LOC_364/A INVX1_LOC_131/A 0.09fF
C24038 NAND2X1_LOC_717/Y NAND2X1_LOC_853/Y 0.02fF
C24039 INVX1_LOC_201/Y NOR2X1_LOC_459/A 0.39fF
C24040 INVX1_LOC_41/A INVX1_LOC_83/A 0.34fF
C24041 NAND2X1_LOC_717/Y NAND2X1_LOC_705/a_36_24# 0.00fF
C24042 INVX1_LOC_270/A NAND2X1_LOC_93/B 0.07fF
C24043 INVX1_LOC_14/A INVX1_LOC_74/Y 0.04fF
C24044 INVX1_LOC_279/A NOR2X1_LOC_344/a_36_216# 0.00fF
C24045 INVX1_LOC_84/A INVX1_LOC_273/A 0.03fF
C24046 INVX1_LOC_57/A NOR2X1_LOC_743/Y 0.05fF
C24047 NOR2X1_LOC_536/A NOR2X1_LOC_109/Y 0.09fF
C24048 INVX1_LOC_36/Y NAND2X1_LOC_473/A 0.11fF
C24049 NAND2X1_LOC_308/Y INVX1_LOC_10/A 0.02fF
C24050 NAND2X1_LOC_477/A NAND2X1_LOC_392/Y 0.03fF
C24051 INVX1_LOC_30/Y NOR2X1_LOC_16/Y 0.47fF
C24052 NOR2X1_LOC_655/B INVX1_LOC_22/A 0.10fF
C24053 INVX1_LOC_36/A INVX1_LOC_126/Y 0.25fF
C24054 NOR2X1_LOC_91/A INVX1_LOC_297/A 0.03fF
C24055 NAND2X1_LOC_364/A INPUT_0 0.10fF
C24056 INVX1_LOC_2/A NOR2X1_LOC_543/A 0.07fF
C24057 NAND2X1_LOC_253/a_36_24# NOR2X1_LOC_833/B 0.00fF
C24058 NOR2X1_LOC_92/Y INVX1_LOC_46/A 0.06fF
C24059 NOR2X1_LOC_179/Y NAND2X1_LOC_99/A 0.02fF
C24060 NOR2X1_LOC_209/Y NOR2X1_LOC_302/a_36_216# 0.00fF
C24061 NAND2X1_LOC_860/A INVX1_LOC_70/A 0.07fF
C24062 GATE_741 NOR2X1_LOC_766/Y 0.04fF
C24063 INVX1_LOC_208/A INVX1_LOC_16/A 0.08fF
C24064 NAND2X1_LOC_740/B NOR2X1_LOC_152/Y 0.04fF
C24065 NAND2X1_LOC_740/Y NAND2X1_LOC_770/a_36_24# 0.01fF
C24066 INVX1_LOC_103/A INVX1_LOC_20/A 0.12fF
C24067 NAND2X1_LOC_214/B INVX1_LOC_9/A 0.00fF
C24068 NOR2X1_LOC_598/B INVX1_LOC_307/A 0.17fF
C24069 NAND2X1_LOC_400/a_36_24# NAND2X1_LOC_773/B 0.00fF
C24070 INVX1_LOC_48/Y INVX1_LOC_12/Y 0.77fF
C24071 INVX1_LOC_71/A INVX1_LOC_67/Y 0.08fF
C24072 NOR2X1_LOC_746/a_36_216# INVX1_LOC_30/A 0.00fF
C24073 INVX1_LOC_88/A VDD 1.93fF
C24074 NOR2X1_LOC_172/Y NAND2X1_LOC_652/Y 0.00fF
C24075 NOR2X1_LOC_383/B INVX1_LOC_220/A 0.01fF
C24076 INVX1_LOC_286/A INVX1_LOC_18/A 0.01fF
C24077 D_INPUT_0 NOR2X1_LOC_168/B 0.03fF
C24078 INVX1_LOC_208/Y NAND2X1_LOC_349/B 0.00fF
C24079 NAND2X1_LOC_550/A NOR2X1_LOC_253/Y 0.02fF
C24080 INVX1_LOC_39/A NOR2X1_LOC_271/Y 0.00fF
C24081 NOR2X1_LOC_6/B NOR2X1_LOC_5/a_36_216# 0.01fF
C24082 NOR2X1_LOC_142/Y NOR2X1_LOC_735/Y -0.01fF
C24083 NOR2X1_LOC_796/B VDD 0.48fF
C24084 NOR2X1_LOC_588/A INVX1_LOC_30/A 0.03fF
C24085 NOR2X1_LOC_570/A NOR2X1_LOC_500/Y 0.03fF
C24086 NOR2X1_LOC_598/B NOR2X1_LOC_445/B 0.12fF
C24087 INVX1_LOC_97/Y INVX1_LOC_307/A -0.01fF
C24088 NOR2X1_LOC_146/Y NAND2X1_LOC_149/B 0.18fF
C24089 NOR2X1_LOC_122/A NOR2X1_LOC_363/Y 0.07fF
C24090 NAND2X1_LOC_842/B INVX1_LOC_104/A 0.00fF
C24091 NAND2X1_LOC_150/a_36_24# INVX1_LOC_8/A 0.00fF
C24092 NOR2X1_LOC_160/B NOR2X1_LOC_35/Y 0.11fF
C24093 INVX1_LOC_27/A INVX1_LOC_9/A 0.28fF
C24094 INVX1_LOC_303/A NOR2X1_LOC_721/Y 0.08fF
C24095 NOR2X1_LOC_346/B NOR2X1_LOC_99/B 0.07fF
C24096 NAND2X1_LOC_848/A NAND2X1_LOC_780/Y 0.04fF
C24097 NOR2X1_LOC_416/A INVX1_LOC_3/A 0.42fF
C24098 INVX1_LOC_136/A NOR2X1_LOC_552/A 0.10fF
C24099 INVX1_LOC_53/A NOR2X1_LOC_435/B 0.03fF
C24100 INVX1_LOC_182/A NOR2X1_LOC_348/B 0.50fF
C24101 NOR2X1_LOC_38/B INVX1_LOC_3/Y 0.26fF
C24102 NOR2X1_LOC_736/Y INVX1_LOC_266/Y 0.07fF
C24103 INVX1_LOC_161/Y NAND2X1_LOC_687/A 0.01fF
C24104 NAND2X1_LOC_805/a_36_24# NAND2X1_LOC_287/B 0.00fF
C24105 NAND2X1_LOC_656/A INVX1_LOC_91/A 0.08fF
C24106 NAND2X1_LOC_780/a_36_24# NOR2X1_LOC_109/Y 0.01fF
C24107 INVX1_LOC_136/A NOR2X1_LOC_566/a_36_216# 0.00fF
C24108 NOR2X1_LOC_91/A NOR2X1_LOC_89/A 3.40fF
C24109 INVX1_LOC_19/A INVX1_LOC_29/Y 0.03fF
C24110 NAND2X1_LOC_656/Y NAND2X1_LOC_660/Y 0.03fF
C24111 NOR2X1_LOC_400/A NAND2X1_LOC_659/A 0.01fF
C24112 D_INPUT_0 NOR2X1_LOC_789/A 0.01fF
C24113 NOR2X1_LOC_106/Y NOR2X1_LOC_78/A 0.03fF
C24114 NAND2X1_LOC_778/Y NOR2X1_LOC_88/Y 0.12fF
C24115 NOR2X1_LOC_315/Y NOR2X1_LOC_184/a_36_216# 0.01fF
C24116 INVX1_LOC_21/A NOR2X1_LOC_831/B 0.49fF
C24117 NOR2X1_LOC_389/A INVX1_LOC_117/A 0.10fF
C24118 D_INPUT_6 NAND2X1_LOC_50/a_36_24# 0.00fF
C24119 NOR2X1_LOC_262/a_36_216# NOR2X1_LOC_89/A 0.00fF
C24120 NOR2X1_LOC_214/B INVX1_LOC_290/A 0.06fF
C24121 VDD NOR2X1_LOC_500/B 1.52fF
C24122 NOR2X1_LOC_160/B NAND2X1_LOC_236/a_36_24# 0.00fF
C24123 INVX1_LOC_121/A INVX1_LOC_83/A 0.02fF
C24124 INVX1_LOC_208/A INVX1_LOC_28/A 0.11fF
C24125 NAND2X1_LOC_785/A INPUT_0 0.02fF
C24126 INVX1_LOC_17/A NOR2X1_LOC_489/A 0.00fF
C24127 INVX1_LOC_11/Y NOR2X1_LOC_484/Y 0.01fF
C24128 NOR2X1_LOC_756/Y INVX1_LOC_25/Y 0.01fF
C24129 D_INPUT_0 NAND2X1_LOC_656/Y 0.12fF
C24130 NOR2X1_LOC_89/A INVX1_LOC_23/A 4.18fF
C24131 INVX1_LOC_233/Y NAND2X1_LOC_500/B 0.07fF
C24132 NOR2X1_LOC_773/Y NOR2X1_LOC_322/Y 0.45fF
C24133 NOR2X1_LOC_291/Y NAND2X1_LOC_489/Y 0.01fF
C24134 NAND2X1_LOC_778/Y INVX1_LOC_84/A 0.01fF
C24135 NOR2X1_LOC_598/B INVX1_LOC_12/A 0.09fF
C24136 NOR2X1_LOC_577/Y INVX1_LOC_291/Y 0.16fF
C24137 NOR2X1_LOC_6/B INVX1_LOC_123/A 0.05fF
C24138 INVX1_LOC_182/A INVX1_LOC_22/A 0.09fF
C24139 NOR2X1_LOC_15/Y NOR2X1_LOC_88/Y 0.20fF
C24140 NOR2X1_LOC_550/B INVX1_LOC_247/A 0.01fF
C24141 INVX1_LOC_227/A INVX1_LOC_313/Y 0.00fF
C24142 D_INPUT_0 INVX1_LOC_132/Y 0.03fF
C24143 INVX1_LOC_34/A NOR2X1_LOC_405/A 0.04fF
C24144 INVX1_LOC_136/A NOR2X1_LOC_813/Y 0.02fF
C24145 INVX1_LOC_312/Y NAND2X1_LOC_848/A 0.10fF
C24146 INVX1_LOC_256/A INVX1_LOC_131/Y 0.21fF
C24147 INVX1_LOC_36/A NOR2X1_LOC_536/A 0.31fF
C24148 NAND2X1_LOC_725/A INVX1_LOC_12/A 2.45fF
C24149 NAND2X1_LOC_837/Y INVX1_LOC_46/A 0.08fF
C24150 INVX1_LOC_282/A NAND2X1_LOC_493/a_36_24# 0.00fF
C24151 NOR2X1_LOC_170/A INVX1_LOC_23/A 0.02fF
C24152 INVX1_LOC_41/Y NAND2X1_LOC_721/A 0.12fF
C24153 NOR2X1_LOC_15/Y INVX1_LOC_84/A 0.40fF
C24154 INVX1_LOC_136/A INVX1_LOC_280/A 0.03fF
C24155 NOR2X1_LOC_561/Y NOR2X1_LOC_597/Y 0.04fF
C24156 INVX1_LOC_277/A NOR2X1_LOC_209/B 0.01fF
C24157 NOR2X1_LOC_186/Y NOR2X1_LOC_831/Y 0.02fF
C24158 INVX1_LOC_303/A VDD 0.02fF
C24159 INVX1_LOC_133/Y NOR2X1_LOC_269/Y 0.00fF
C24160 NOR2X1_LOC_596/A INVX1_LOC_117/A 0.14fF
C24161 NOR2X1_LOC_273/Y INVX1_LOC_281/A 0.94fF
C24162 NOR2X1_LOC_672/Y VDD 0.22fF
C24163 NOR2X1_LOC_693/a_36_216# NOR2X1_LOC_693/Y 0.01fF
C24164 NOR2X1_LOC_437/Y NOR2X1_LOC_363/Y 0.31fF
C24165 INVX1_LOC_36/A NOR2X1_LOC_655/Y 0.01fF
C24166 NAND2X1_LOC_474/Y INVX1_LOC_29/A 0.01fF
C24167 INVX1_LOC_232/A INVX1_LOC_48/A 0.46fF
C24168 NAND2X1_LOC_477/A NOR2X1_LOC_368/Y 0.12fF
C24169 INVX1_LOC_41/A INVX1_LOC_46/A 2.28fF
C24170 NOR2X1_LOC_222/Y INVX1_LOC_91/A 0.15fF
C24171 NAND2X1_LOC_231/Y NOR2X1_LOC_405/A 0.10fF
C24172 NAND2X1_LOC_59/B VDD 0.74fF
C24173 NAND2X1_LOC_573/Y NOR2X1_LOC_831/Y 0.12fF
C24174 NAND2X1_LOC_357/B NOR2X1_LOC_279/Y 0.04fF
C24175 INVX1_LOC_18/A INVX1_LOC_54/A 1.08fF
C24176 INVX1_LOC_240/A INVX1_LOC_20/A 0.20fF
C24177 NOR2X1_LOC_91/Y INVX1_LOC_118/A 0.04fF
C24178 INVX1_LOC_36/A NAND2X1_LOC_93/B 0.10fF
C24179 INVX1_LOC_129/A INVX1_LOC_87/A 0.02fF
C24180 NOR2X1_LOC_383/B INVX1_LOC_23/Y 0.02fF
C24181 NOR2X1_LOC_152/a_36_216# INVX1_LOC_38/A 0.00fF
C24182 NOR2X1_LOC_237/Y NOR2X1_LOC_536/A 0.07fF
C24183 NOR2X1_LOC_456/Y NOR2X1_LOC_465/Y 0.74fF
C24184 NOR2X1_LOC_544/A INVX1_LOC_65/A 0.01fF
C24185 NOR2X1_LOC_829/A INVX1_LOC_296/Y 0.00fF
C24186 INVX1_LOC_105/A INVX1_LOC_38/A 0.07fF
C24187 NOR2X1_LOC_92/Y NOR2X1_LOC_671/Y 0.01fF
C24188 INVX1_LOC_83/A NAND2X1_LOC_662/B 0.15fF
C24189 INVX1_LOC_27/A NOR2X1_LOC_861/Y 0.10fF
C24190 NAND2X1_LOC_477/A INVX1_LOC_46/A 0.01fF
C24191 INVX1_LOC_21/A NAND2X1_LOC_430/B 0.00fF
C24192 NOR2X1_LOC_637/Y INVX1_LOC_54/A 0.20fF
C24193 NAND2X1_LOC_722/A NOR2X1_LOC_305/Y 0.02fF
C24194 INVX1_LOC_168/A VDD 0.12fF
C24195 NOR2X1_LOC_207/A INVX1_LOC_46/A 0.01fF
C24196 NAND2X1_LOC_357/B NAND2X1_LOC_804/Y 0.01fF
C24197 INVX1_LOC_220/Y INVX1_LOC_91/A 0.32fF
C24198 INVX1_LOC_291/Y INVX1_LOC_22/A 0.03fF
C24199 INVX1_LOC_45/A INVX1_LOC_285/A 0.07fF
C24200 NAND2X1_LOC_798/a_36_24# INVX1_LOC_118/A 0.00fF
C24201 INVX1_LOC_36/A NAND2X1_LOC_780/a_36_24# 0.01fF
C24202 NOR2X1_LOC_756/Y INVX1_LOC_75/A 0.10fF
C24203 INVX1_LOC_172/A INVX1_LOC_54/A 0.07fF
C24204 NOR2X1_LOC_91/A NAND2X1_LOC_804/A 0.01fF
C24205 INVX1_LOC_94/A INVX1_LOC_92/A 0.07fF
C24206 NOR2X1_LOC_84/Y INVX1_LOC_12/Y 0.02fF
C24207 NOR2X1_LOC_208/Y NAND2X1_LOC_93/B 0.07fF
C24208 INVX1_LOC_36/A NOR2X1_LOC_649/B 0.04fF
C24209 NOR2X1_LOC_322/Y INVX1_LOC_140/A 0.10fF
C24210 NOR2X1_LOC_329/B INVX1_LOC_79/A 0.03fF
C24211 NAND2X1_LOC_577/A INVX1_LOC_203/A 0.07fF
C24212 INVX1_LOC_45/A NOR2X1_LOC_814/A 0.16fF
C24213 NOR2X1_LOC_356/A NOR2X1_LOC_337/A 0.14fF
C24214 NOR2X1_LOC_309/Y NOR2X1_LOC_536/A 0.10fF
C24215 INVX1_LOC_36/A INVX1_LOC_3/A 0.43fF
C24216 NOR2X1_LOC_203/Y VDD 0.03fF
C24217 INVX1_LOC_290/A NOR2X1_LOC_275/A 0.14fF
C24218 NOR2X1_LOC_516/B NOR2X1_LOC_35/Y 0.05fF
C24219 NOR2X1_LOC_561/Y NOR2X1_LOC_657/B 0.03fF
C24220 NOR2X1_LOC_557/Y NOR2X1_LOC_612/Y 0.03fF
C24221 NOR2X1_LOC_377/Y INVX1_LOC_193/A 0.19fF
C24222 NAND2X1_LOC_209/a_36_24# D_INPUT_5 0.01fF
C24223 NOR2X1_LOC_15/Y INVX1_LOC_15/A 0.17fF
C24224 INVX1_LOC_70/Y NOR2X1_LOC_123/B 0.05fF
C24225 NAND2X1_LOC_799/A NOR2X1_LOC_48/B 0.16fF
C24226 INVX1_LOC_77/A NOR2X1_LOC_216/B 0.07fF
C24227 INVX1_LOC_239/A NAND2X1_LOC_618/Y 0.00fF
C24228 INVX1_LOC_31/A NOR2X1_LOC_89/A 0.07fF
C24229 INVX1_LOC_24/A NOR2X1_LOC_673/A 0.00fF
C24230 INVX1_LOC_206/A INVX1_LOC_9/A 0.05fF
C24231 INVX1_LOC_87/A NOR2X1_LOC_440/B 0.50fF
C24232 INVX1_LOC_71/A INVX1_LOC_285/A 0.10fF
C24233 NAND2X1_LOC_364/Y NOR2X1_LOC_865/Y 0.09fF
C24234 NOR2X1_LOC_380/A INVX1_LOC_11/Y 0.00fF
C24235 NOR2X1_LOC_309/Y NAND2X1_LOC_93/B 0.03fF
C24236 NOR2X1_LOC_32/B NOR2X1_LOC_392/Y 0.01fF
C24237 INVX1_LOC_71/A NOR2X1_LOC_814/A 0.12fF
C24238 NOR2X1_LOC_428/Y NAND2X1_LOC_430/B 0.12fF
C24239 NOR2X1_LOC_329/B INVX1_LOC_91/A 3.98fF
C24240 NOR2X1_LOC_716/B NAND2X1_LOC_572/B 1.18fF
C24241 D_INPUT_7 INPUT_7 0.03fF
C24242 INVX1_LOC_80/A VDD 0.12fF
C24243 NAND2X1_LOC_538/Y INVX1_LOC_94/Y 0.02fF
C24244 NAND2X1_LOC_200/B INVX1_LOC_9/A 0.01fF
C24245 NOR2X1_LOC_299/Y INVX1_LOC_46/A 4.64fF
C24246 INVX1_LOC_143/A NOR2X1_LOC_612/Y 0.01fF
C24247 NAND2X1_LOC_842/B NAND2X1_LOC_674/a_36_24# 0.01fF
C24248 INVX1_LOC_62/A INVX1_LOC_2/Y 0.02fF
C24249 INVX1_LOC_131/A NOR2X1_LOC_113/A 0.04fF
C24250 INVX1_LOC_292/A INVX1_LOC_4/A 0.07fF
C24251 NOR2X1_LOC_250/A INVX1_LOC_94/Y 0.08fF
C24252 INVX1_LOC_131/A NOR2X1_LOC_405/A 0.03fF
C24253 NOR2X1_LOC_360/Y NOR2X1_LOC_327/a_36_216# 0.02fF
C24254 INVX1_LOC_124/A NOR2X1_LOC_216/B 0.05fF
C24255 NOR2X1_LOC_457/A INVX1_LOC_271/Y 0.02fF
C24256 INVX1_LOC_153/Y NOR2X1_LOC_66/Y 0.06fF
C24257 NOR2X1_LOC_81/a_36_216# NAND2X1_LOC_63/Y 0.00fF
C24258 INVX1_LOC_308/Y NOR2X1_LOC_301/A 0.06fF
C24259 NOR2X1_LOC_698/a_36_216# NOR2X1_LOC_748/A 0.01fF
C24260 INVX1_LOC_18/A NOR2X1_LOC_48/B 0.07fF
C24261 INVX1_LOC_298/Y NAND2X1_LOC_53/Y 0.07fF
C24262 NAND2X1_LOC_308/B VDD 0.03fF
C24263 INVX1_LOC_41/A NOR2X1_LOC_68/Y 0.01fF
C24264 NOR2X1_LOC_376/a_36_216# NOR2X1_LOC_89/A 0.00fF
C24265 NAND2X1_LOC_778/Y INVX1_LOC_278/A 0.10fF
C24266 INVX1_LOC_21/A NOR2X1_LOC_790/B 0.03fF
C24267 INPUT_0 NOR2X1_LOC_113/A 0.02fF
C24268 INVX1_LOC_224/A NOR2X1_LOC_668/Y 0.01fF
C24269 INPUT_0 NOR2X1_LOC_405/A 0.07fF
C24270 NOR2X1_LOC_647/A NOR2X1_LOC_817/Y 0.36fF
C24271 INVX1_LOC_244/A VDD 0.17fF
C24272 INVX1_LOC_28/A NAND2X1_LOC_211/Y 0.05fF
C24273 NOR2X1_LOC_309/Y NOR2X1_LOC_661/A 0.05fF
C24274 NOR2X1_LOC_91/A INVX1_LOC_11/A 2.48fF
C24275 INVX1_LOC_35/A NAND2X1_LOC_391/Y 4.60fF
C24276 INVX1_LOC_58/A NOR2X1_LOC_468/Y 0.00fF
C24277 NAND2X1_LOC_711/B NOR2X1_LOC_48/B 0.05fF
C24278 NOR2X1_LOC_303/Y INVX1_LOC_290/Y 0.10fF
C24279 NAND2X1_LOC_840/B NOR2X1_LOC_88/Y 0.03fF
C24280 INVX1_LOC_96/Y INVX1_LOC_84/A 0.10fF
C24281 INVX1_LOC_58/A NAND2X1_LOC_190/Y 0.10fF
C24282 NAND2X1_LOC_9/Y NOR2X1_LOC_92/Y 0.03fF
C24283 INVX1_LOC_25/A INVX1_LOC_269/A 0.29fF
C24284 NOR2X1_LOC_846/Y INVX1_LOC_5/A 0.32fF
C24285 NOR2X1_LOC_381/Y D_INPUT_1 0.04fF
C24286 INVX1_LOC_17/A NAND2X1_LOC_464/B 0.00fF
C24287 NOR2X1_LOC_440/Y NOR2X1_LOC_79/A 0.08fF
C24288 NAND2X1_LOC_361/Y INVX1_LOC_106/Y 0.00fF
C24289 INVX1_LOC_30/A INVX1_LOC_271/Y 0.07fF
C24290 NOR2X1_LOC_332/A NOR2X1_LOC_54/a_36_216# 0.01fF
C24291 INVX1_LOC_18/A NAND2X1_LOC_3/B 0.27fF
C24292 INVX1_LOC_233/A NOR2X1_LOC_92/Y 0.07fF
C24293 INVX1_LOC_256/A INVX1_LOC_270/A 3.12fF
C24294 NOR2X1_LOC_789/A INVX1_LOC_46/Y 0.02fF
C24295 NAND2X1_LOC_773/Y NAND2X1_LOC_363/B 0.01fF
C24296 INVX1_LOC_172/A NOR2X1_LOC_48/B 0.07fF
C24297 NOR2X1_LOC_602/A NAND2X1_LOC_175/Y 0.02fF
C24298 INVX1_LOC_278/A NOR2X1_LOC_15/Y 0.08fF
C24299 NOR2X1_LOC_598/B NOR2X1_LOC_643/A 0.01fF
C24300 INVX1_LOC_268/A INVX1_LOC_113/A 0.07fF
C24301 INVX1_LOC_11/A INVX1_LOC_23/A 0.17fF
C24302 NOR2X1_LOC_730/A NOR2X1_LOC_155/A 0.01fF
C24303 INVX1_LOC_233/Y NAND2X1_LOC_725/B 0.07fF
C24304 INVX1_LOC_34/A INVX1_LOC_109/Y 0.00fF
C24305 INPUT_0 NOR2X1_LOC_857/A 0.07fF
C24306 NOR2X1_LOC_860/B INVX1_LOC_15/A 0.15fF
C24307 NAND2X1_LOC_308/Y INVX1_LOC_12/A 0.03fF
C24308 INVX1_LOC_50/A NOR2X1_LOC_483/B 0.04fF
C24309 NOR2X1_LOC_68/A NOR2X1_LOC_158/a_36_216# 0.01fF
C24310 INVX1_LOC_224/Y NOR2X1_LOC_590/A 0.02fF
C24311 NOR2X1_LOC_411/a_36_216# NAND2X1_LOC_725/B 0.00fF
C24312 INVX1_LOC_57/Y INVX1_LOC_23/Y 0.01fF
C24313 NOR2X1_LOC_689/Y NAND2X1_LOC_733/Y 0.03fF
C24314 INVX1_LOC_64/A INVX1_LOC_103/A 0.27fF
C24315 NOR2X1_LOC_387/A NAND2X1_LOC_453/A 0.12fF
C24316 NAND2X1_LOC_652/Y INVX1_LOC_38/A 0.04fF
C24317 INVX1_LOC_58/A NOR2X1_LOC_389/A 0.10fF
C24318 INVX1_LOC_251/Y NAND2X1_LOC_74/B 0.06fF
C24319 INVX1_LOC_24/A NOR2X1_LOC_409/B 0.07fF
C24320 INVX1_LOC_315/Y NOR2X1_LOC_35/Y 0.03fF
C24321 NOR2X1_LOC_19/B INVX1_LOC_9/A 0.00fF
C24322 NOR2X1_LOC_798/A INVX1_LOC_24/Y 0.03fF
C24323 NAND2X1_LOC_377/Y NAND2X1_LOC_659/A -0.00fF
C24324 NOR2X1_LOC_852/B NOR2X1_LOC_839/B 0.00fF
C24325 INVX1_LOC_13/Y NOR2X1_LOC_361/B 0.10fF
C24326 NOR2X1_LOC_567/B NOR2X1_LOC_729/A 0.07fF
C24327 NOR2X1_LOC_510/Y INVX1_LOC_88/A 0.92fF
C24328 NOR2X1_LOC_537/Y NOR2X1_LOC_67/Y 0.02fF
C24329 INVX1_LOC_64/A INVX1_LOC_292/A 0.07fF
C24330 INVX1_LOC_279/A NAND2X1_LOC_475/Y 0.10fF
C24331 NAND2X1_LOC_738/B NAND2X1_LOC_741/B 0.03fF
C24332 NAND2X1_LOC_30/Y NAND2X1_LOC_18/a_36_24# 0.00fF
C24333 NOR2X1_LOC_544/A NOR2X1_LOC_830/Y 0.01fF
C24334 NOR2X1_LOC_388/Y NAND2X1_LOC_647/B 0.06fF
C24335 D_INPUT_1 NOR2X1_LOC_248/Y 0.01fF
C24336 NOR2X1_LOC_635/A INVX1_LOC_15/A 0.01fF
C24337 INVX1_LOC_83/A NOR2X1_LOC_435/B 0.21fF
C24338 NOR2X1_LOC_366/Y NOR2X1_LOC_127/Y 0.00fF
C24339 NOR2X1_LOC_500/Y INVX1_LOC_29/A 0.11fF
C24340 INPUT_6 NAND2X1_LOC_36/A 0.27fF
C24341 INVX1_LOC_226/Y INVX1_LOC_29/A 0.06fF
C24342 INVX1_LOC_27/A NAND2X1_LOC_20/B 0.04fF
C24343 NAND2X1_LOC_708/Y INVX1_LOC_286/Y 0.05fF
C24344 INVX1_LOC_21/A D_GATE_741 0.06fF
C24345 NAND2X1_LOC_198/B INVX1_LOC_57/A 0.02fF
C24346 NAND2X1_LOC_724/A NAND2X1_LOC_303/Y 0.01fF
C24347 INVX1_LOC_15/Y INVX1_LOC_15/A 0.00fF
C24348 NOR2X1_LOC_617/Y NOR2X1_LOC_19/a_36_216# 0.00fF
C24349 NOR2X1_LOC_91/A NOR2X1_LOC_433/A 0.03fF
C24350 INVX1_LOC_269/A INVX1_LOC_1/A 0.25fF
C24351 NOR2X1_LOC_749/a_36_216# INVX1_LOC_63/A 0.01fF
C24352 NOR2X1_LOC_303/a_36_216# INVX1_LOC_179/A 0.00fF
C24353 INVX1_LOC_21/A NAND2X1_LOC_352/B 0.15fF
C24354 INVX1_LOC_58/A NOR2X1_LOC_596/A 0.17fF
C24355 INVX1_LOC_101/Y NOR2X1_LOC_205/Y 0.00fF
C24356 NAND2X1_LOC_859/Y NOR2X1_LOC_89/A 0.02fF
C24357 NOR2X1_LOC_361/B INVX1_LOC_88/A 0.14fF
C24358 INVX1_LOC_10/A INVX1_LOC_29/A 0.75fF
C24359 D_INPUT_1 NAND2X1_LOC_187/a_36_24# 0.00fF
C24360 NAND2X1_LOC_725/A INVX1_LOC_217/A 0.10fF
C24361 INVX1_LOC_94/A INVX1_LOC_53/A 0.02fF
C24362 NOR2X1_LOC_669/a_36_216# NOR2X1_LOC_816/A 0.00fF
C24363 INVX1_LOC_48/Y NOR2X1_LOC_160/B 0.07fF
C24364 NOR2X1_LOC_248/Y NOR2X1_LOC_652/Y 0.01fF
C24365 INVX1_LOC_102/Y INVX1_LOC_285/A 1.24fF
C24366 INVX1_LOC_71/A NOR2X1_LOC_292/a_36_216# 0.12fF
C24367 INVX1_LOC_50/A INVX1_LOC_33/A 1.46fF
C24368 NOR2X1_LOC_433/A INVX1_LOC_23/A 3.85fF
C24369 NOR2X1_LOC_690/Y NOR2X1_LOC_48/B 0.05fF
C24370 NOR2X1_LOC_474/A INVX1_LOC_23/A 0.00fF
C24371 NOR2X1_LOC_718/B NOR2X1_LOC_302/A 0.03fF
C24372 INVX1_LOC_28/A NOR2X1_LOC_605/A 0.41fF
C24373 INVX1_LOC_162/Y NAND2X1_LOC_286/B 0.01fF
C24374 INVX1_LOC_182/Y NAND2X1_LOC_475/Y 0.03fF
C24375 INVX1_LOC_310/Y INVX1_LOC_57/A 0.07fF
C24376 INPUT_1 NAND2X1_LOC_82/Y 0.45fF
C24377 NOR2X1_LOC_91/A NOR2X1_LOC_52/B 0.06fF
C24378 NOR2X1_LOC_593/Y INVX1_LOC_23/A 0.02fF
C24379 NAND2X1_LOC_303/Y NAND2X1_LOC_389/a_36_24# 0.06fF
C24380 NOR2X1_LOC_537/A INVX1_LOC_58/Y 0.04fF
C24381 INVX1_LOC_313/A NOR2X1_LOC_89/A 0.37fF
C24382 INVX1_LOC_235/Y INVX1_LOC_195/A 0.05fF
C24383 NOR2X1_LOC_178/Y INVX1_LOC_314/Y 0.01fF
C24384 NAND2X1_LOC_866/B NOR2X1_LOC_89/A 0.02fF
C24385 NAND2X1_LOC_222/B INVX1_LOC_31/A 0.01fF
C24386 INVX1_LOC_151/A INVX1_LOC_23/A 0.01fF
C24387 INVX1_LOC_46/A NOR2X1_LOC_494/a_36_216# 0.00fF
C24388 NOR2X1_LOC_67/A INVX1_LOC_26/A 0.14fF
C24389 NAND2X1_LOC_9/Y INVX1_LOC_41/A 0.01fF
C24390 NAND2X1_LOC_773/Y INVX1_LOC_30/A 0.19fF
C24391 INVX1_LOC_224/A INVX1_LOC_31/A 0.03fF
C24392 D_INPUT_1 NOR2X1_LOC_6/B 0.26fF
C24393 NAND2X1_LOC_725/A NAND2X1_LOC_787/B 0.19fF
C24394 INVX1_LOC_11/A INVX1_LOC_31/A 0.27fF
C24395 NOR2X1_LOC_52/B INVX1_LOC_23/A 4.93fF
C24396 NOR2X1_LOC_795/a_36_216# INVX1_LOC_15/A 0.01fF
C24397 NAND2X1_LOC_72/Y INVX1_LOC_33/A 0.08fF
C24398 NOR2X1_LOC_590/A NOR2X1_LOC_541/Y 0.58fF
C24399 NAND2X1_LOC_807/Y NOR2X1_LOC_89/A 0.07fF
C24400 NAND2X1_LOC_381/Y INVX1_LOC_31/A 0.06fF
C24401 NOR2X1_LOC_82/A NOR2X1_LOC_514/A 0.01fF
C24402 NOR2X1_LOC_456/Y NOR2X1_LOC_180/Y 0.01fF
C24403 NAND2X1_LOC_560/A INVX1_LOC_12/A 0.03fF
C24404 NAND2X1_LOC_552/A NAND2X1_LOC_833/Y 0.52fF
C24405 NOR2X1_LOC_71/Y INVX1_LOC_47/Y 0.01fF
C24406 GATE_741 NAND2X1_LOC_866/A 0.01fF
C24407 NAND2X1_LOC_860/A NOR2X1_LOC_316/Y 0.03fF
C24408 NOR2X1_LOC_232/Y NOR2X1_LOC_384/Y 0.02fF
C24409 INVX1_LOC_45/A NAND2X1_LOC_803/B 0.02fF
C24410 INVX1_LOC_233/A NAND2X1_LOC_477/A 0.10fF
C24411 INVX1_LOC_64/A INVX1_LOC_240/A 0.07fF
C24412 INVX1_LOC_28/A NAND2X1_LOC_791/a_36_24# 0.01fF
C24413 NAND2X1_LOC_9/Y NOR2X1_LOC_398/Y 0.01fF
C24414 INVX1_LOC_256/A INVX1_LOC_36/A 0.19fF
C24415 NOR2X1_LOC_410/a_36_216# INVX1_LOC_11/A 0.02fF
C24416 NOR2X1_LOC_552/Y INVX1_LOC_19/A 0.01fF
C24417 NOR2X1_LOC_67/A NOR2X1_LOC_255/Y 0.04fF
C24418 NAND2X1_LOC_513/B INVX1_LOC_77/A 0.08fF
C24419 INVX1_LOC_103/A INVX1_LOC_130/Y 0.01fF
C24420 NAND2X1_LOC_9/Y INVX1_LOC_64/Y 0.40fF
C24421 INVX1_LOC_304/Y NAND2X1_LOC_725/A 0.23fF
C24422 NAND2X1_LOC_740/Y INVX1_LOC_34/A 0.03fF
C24423 INVX1_LOC_37/A INVX1_LOC_274/A 0.69fF
C24424 INVX1_LOC_41/A NOR2X1_LOC_798/A 0.03fF
C24425 INVX1_LOC_316/A NAND2X1_LOC_141/Y 0.15fF
C24426 NOR2X1_LOC_322/Y INVX1_LOC_42/A 0.08fF
C24427 NAND2X1_LOC_800/Y NOR2X1_LOC_409/B 0.00fF
C24428 INVX1_LOC_25/A NAND2X1_LOC_563/A 0.02fF
C24429 INVX1_LOC_21/A INVX1_LOC_212/Y 0.01fF
C24430 INVX1_LOC_17/A NOR2X1_LOC_523/B 0.02fF
C24431 INVX1_LOC_178/A NAND2X1_LOC_833/Y 0.01fF
C24432 INVX1_LOC_298/Y INVX1_LOC_10/A 0.03fF
C24433 INVX1_LOC_21/A NOR2X1_LOC_344/A 0.02fF
C24434 NOR2X1_LOC_106/A INVX1_LOC_94/Y 0.14fF
C24435 VDD NOR2X1_LOC_99/Y 0.49fF
C24436 INVX1_LOC_249/A NAND2X1_LOC_67/Y 1.52fF
C24437 NOR2X1_LOC_456/Y NOR2X1_LOC_458/B 0.01fF
C24438 INVX1_LOC_45/A NOR2X1_LOC_590/A 3.48fF
C24439 NOR2X1_LOC_231/B NOR2X1_LOC_641/B 0.00fF
C24440 NAND2X1_LOC_381/a_36_24# NOR2X1_LOC_554/B 0.01fF
C24441 NOR2X1_LOC_381/Y D_INPUT_2 0.11fF
C24442 NAND2X1_LOC_721/A INVX1_LOC_185/A 0.12fF
C24443 INVX1_LOC_53/Y INVX1_LOC_57/A 0.04fF
C24444 NOR2X1_LOC_205/a_36_216# INVX1_LOC_53/A 0.01fF
C24445 NAND2X1_LOC_350/A INVX1_LOC_18/A 0.07fF
C24446 INVX1_LOC_104/A NOR2X1_LOC_674/Y 0.09fF
C24447 INVX1_LOC_1/Y INVX1_LOC_270/Y 0.03fF
C24448 NOR2X1_LOC_590/A NOR2X1_LOC_568/A 0.11fF
C24449 NOR2X1_LOC_136/Y INVX1_LOC_53/A 0.04fF
C24450 NAND2X1_LOC_382/a_36_24# NOR2X1_LOC_554/B 0.01fF
C24451 NOR2X1_LOC_383/Y NOR2X1_LOC_383/B 0.80fF
C24452 NOR2X1_LOC_746/Y NAND2X1_LOC_782/B 0.01fF
C24453 NAND2X1_LOC_51/B NAND2X1_LOC_430/B 0.01fF
C24454 INVX1_LOC_93/A NAND2X1_LOC_650/a_36_24# 0.01fF
C24455 INVX1_LOC_6/A NOR2X1_LOC_89/A 1.41fF
C24456 INVX1_LOC_64/A NOR2X1_LOC_533/A 0.03fF
C24457 NOR2X1_LOC_473/B INVX1_LOC_78/A 0.15fF
C24458 NOR2X1_LOC_231/B NOR2X1_LOC_751/Y 0.04fF
C24459 INVX1_LOC_217/A NOR2X1_LOC_372/A 0.01fF
C24460 NOR2X1_LOC_323/a_36_216# INVX1_LOC_185/A 0.00fF
C24461 INVX1_LOC_21/A NAND2X1_LOC_357/B 0.14fF
C24462 INVX1_LOC_256/A INVX1_LOC_145/A 0.33fF
C24463 NOR2X1_LOC_488/Y NAND2X1_LOC_793/B 0.09fF
C24464 INVX1_LOC_48/A NAND2X1_LOC_263/a_36_24# 0.00fF
C24465 VDD INVX1_LOC_107/Y 0.37fF
C24466 INVX1_LOC_256/A NOR2X1_LOC_208/Y 0.56fF
C24467 INVX1_LOC_34/A NAND2X1_LOC_706/Y 0.03fF
C24468 NOR2X1_LOC_100/A NOR2X1_LOC_849/A 0.00fF
C24469 NOR2X1_LOC_99/B NOR2X1_LOC_843/B 0.07fF
C24470 NOR2X1_LOC_561/Y INVX1_LOC_271/A 0.10fF
C24471 NOR2X1_LOC_45/B NAND2X1_LOC_74/B 0.14fF
C24472 INVX1_LOC_27/A NAND2X1_LOC_629/Y 0.00fF
C24473 NOR2X1_LOC_637/Y NAND2X1_LOC_350/A 0.01fF
C24474 INVX1_LOC_233/Y INVX1_LOC_241/A 0.23fF
C24475 NAND2X1_LOC_554/a_36_24# INVX1_LOC_270/Y 0.05fF
C24476 INVX1_LOC_14/A NAND2X1_LOC_139/A 0.17fF
C24477 NOR2X1_LOC_355/B INVX1_LOC_42/A 2.51fF
C24478 NOR2X1_LOC_590/A INVX1_LOC_71/A 3.20fF
C24479 INVX1_LOC_135/A NOR2X1_LOC_414/Y 0.01fF
C24480 NAND2X1_LOC_625/a_36_24# INVX1_LOC_76/A 0.01fF
C24481 NOR2X1_LOC_65/B NOR2X1_LOC_473/B -0.01fF
C24482 NOR2X1_LOC_187/Y NOR2X1_LOC_348/B 0.03fF
C24483 NOR2X1_LOC_322/Y INVX1_LOC_78/A 0.03fF
C24484 NOR2X1_LOC_790/B NOR2X1_LOC_565/B 0.00fF
C24485 INVX1_LOC_126/A INVX1_LOC_19/A 0.06fF
C24486 NOR2X1_LOC_835/B NOR2X1_LOC_839/B 0.03fF
C24487 NOR2X1_LOC_160/B NOR2X1_LOC_6/a_36_216# 0.02fF
C24488 NOR2X1_LOC_816/A NAND2X1_LOC_833/Y 0.00fF
C24489 INVX1_LOC_36/A NOR2X1_LOC_781/Y 0.01fF
C24490 INVX1_LOC_2/A NAND2X1_LOC_780/Y 0.03fF
C24491 NOR2X1_LOC_15/Y NOR2X1_LOC_16/Y 0.01fF
C24492 NAND2X1_LOC_214/B NOR2X1_LOC_719/A 0.27fF
C24493 NOR2X1_LOC_433/A INVX1_LOC_31/A 0.11fF
C24494 NAND2X1_LOC_654/B NOR2X1_LOC_635/B 0.01fF
C24495 NOR2X1_LOC_798/A NOR2X1_LOC_211/A 0.00fF
C24496 NOR2X1_LOC_361/B INVX1_LOC_168/A 0.38fF
C24497 INVX1_LOC_233/Y NOR2X1_LOC_298/Y 0.10fF
C24498 INVX1_LOC_5/A NOR2X1_LOC_781/A 0.17fF
C24499 INVX1_LOC_88/A INVX1_LOC_177/A 0.01fF
C24500 NOR2X1_LOC_401/A NOR2X1_LOC_84/Y 0.03fF
C24501 INVX1_LOC_256/A NOR2X1_LOC_309/Y 0.14fF
C24502 NOR2X1_LOC_52/Y NOR2X1_LOC_759/Y 0.00fF
C24503 NAND2X1_LOC_209/a_36_24# NAND2X1_LOC_451/Y 0.00fF
C24504 NOR2X1_LOC_593/Y INVX1_LOC_31/A 0.10fF
C24505 NOR2X1_LOC_35/Y NAND2X1_LOC_207/B 1.79fF
C24506 NOR2X1_LOC_471/Y NOR2X1_LOC_718/B 0.02fF
C24507 NAND2X1_LOC_725/B NOR2X1_LOC_526/Y 0.03fF
C24508 NOR2X1_LOC_68/A NAND2X1_LOC_79/Y 0.02fF
C24509 NOR2X1_LOC_270/Y NOR2X1_LOC_759/Y 0.02fF
C24510 INVX1_LOC_5/A NOR2X1_LOC_719/B 0.01fF
C24511 NAND2X1_LOC_313/a_36_24# NOR2X1_LOC_317/B 0.02fF
C24512 VDD INVX1_LOC_272/A 0.92fF
C24513 NOR2X1_LOC_111/A INVX1_LOC_19/A 0.08fF
C24514 NAND2X1_LOC_214/B INVX1_LOC_7/A 1.75fF
C24515 INVX1_LOC_64/A INVX1_LOC_120/A 0.03fF
C24516 NAND2X1_LOC_563/A INVX1_LOC_1/A 1.44fF
C24517 INVX1_LOC_202/A NOR2X1_LOC_270/Y 0.00fF
C24518 NOR2X1_LOC_536/A INVX1_LOC_63/A 0.28fF
C24519 NOR2X1_LOC_155/A INVX1_LOC_92/A 0.15fF
C24520 NOR2X1_LOC_825/Y NOR2X1_LOC_672/a_36_216# 0.00fF
C24521 NAND2X1_LOC_733/Y NAND2X1_LOC_308/Y 0.03fF
C24522 NOR2X1_LOC_160/B NOR2X1_LOC_84/Y 0.05fF
C24523 NAND2X1_LOC_550/A NOR2X1_LOC_482/Y 0.01fF
C24524 INVX1_LOC_27/A NOR2X1_LOC_561/Y 0.07fF
C24525 INVX1_LOC_45/A NAND2X1_LOC_354/B 0.01fF
C24526 INVX1_LOC_50/A NOR2X1_LOC_323/Y 0.03fF
C24527 NOR2X1_LOC_656/Y NOR2X1_LOC_649/B 0.03fF
C24528 INVX1_LOC_31/A NOR2X1_LOC_52/B 0.19fF
C24529 NAND2X1_LOC_579/A INVX1_LOC_22/A 0.08fF
C24530 D_INPUT_0 NOR2X1_LOC_649/Y 0.07fF
C24531 NOR2X1_LOC_846/Y NOR2X1_LOC_332/A 0.04fF
C24532 INVX1_LOC_27/A INVX1_LOC_7/A 0.16fF
C24533 INVX1_LOC_215/A NOR2X1_LOC_321/Y 0.50fF
C24534 VDD NOR2X1_LOC_76/B -0.00fF
C24535 NOR2X1_LOC_694/Y NOR2X1_LOC_11/Y 0.01fF
C24536 NAND2X1_LOC_731/Y NAND2X1_LOC_738/a_36_24# 0.00fF
C24537 INVX1_LOC_69/Y INVX1_LOC_28/Y 0.01fF
C24538 INVX1_LOC_5/A NOR2X1_LOC_180/B 0.08fF
C24539 NOR2X1_LOC_500/A INVX1_LOC_77/A 0.03fF
C24540 INVX1_LOC_77/A NOR2X1_LOC_303/Y 0.01fF
C24541 NOR2X1_LOC_655/Y INVX1_LOC_63/A 0.01fF
C24542 INVX1_LOC_69/Y INVX1_LOC_270/A 0.01fF
C24543 INVX1_LOC_2/A INVX1_LOC_141/Y 3.29fF
C24544 INVX1_LOC_104/A INVX1_LOC_72/A 0.07fF
C24545 NOR2X1_LOC_593/Y INVX1_LOC_111/A 0.03fF
C24546 NOR2X1_LOC_791/B NOR2X1_LOC_392/B 0.13fF
C24547 INVX1_LOC_216/Y INVX1_LOC_255/Y 0.04fF
C24548 NAND2X1_LOC_85/Y NOR2X1_LOC_243/B 0.06fF
C24549 INVX1_LOC_144/A INVX1_LOC_53/A 0.10fF
C24550 NAND2X1_LOC_276/Y NAND2X1_LOC_656/A 0.15fF
C24551 NOR2X1_LOC_226/A INVX1_LOC_141/Y 0.03fF
C24552 INVX1_LOC_2/A INVX1_LOC_312/Y 0.06fF
C24553 NOR2X1_LOC_419/Y NOR2X1_LOC_716/B 0.04fF
C24554 INVX1_LOC_105/A INVX1_LOC_33/A 0.07fF
C24555 INVX1_LOC_186/A NOR2X1_LOC_383/B 0.03fF
C24556 NOR2X1_LOC_730/B INVX1_LOC_53/A 0.01fF
C24557 NOR2X1_LOC_642/a_36_216# NOR2X1_LOC_649/B 0.05fF
C24558 INVX1_LOC_279/A NOR2X1_LOC_457/A 0.36fF
C24559 INVX1_LOC_251/A INVX1_LOC_117/A 0.03fF
C24560 NOR2X1_LOC_318/B INVX1_LOC_270/Y 1.29fF
C24561 INVX1_LOC_1/A NOR2X1_LOC_214/B 0.11fF
C24562 NAND2X1_LOC_180/a_36_24# INVX1_LOC_41/Y 0.00fF
C24563 NOR2X1_LOC_6/B D_INPUT_2 0.18fF
C24564 INVX1_LOC_35/A NOR2X1_LOC_728/B 0.03fF
C24565 NOR2X1_LOC_78/B NOR2X1_LOC_723/a_36_216# 0.00fF
C24566 NOR2X1_LOC_655/B INVX1_LOC_18/A 0.11fF
C24567 NOR2X1_LOC_92/Y NAND2X1_LOC_842/B 0.01fF
C24568 INVX1_LOC_5/A NOR2X1_LOC_569/A 0.01fF
C24569 NOR2X1_LOC_89/A NOR2X1_LOC_79/A 0.20fF
C24570 INVX1_LOC_307/A INVX1_LOC_29/A 0.01fF
C24571 NOR2X1_LOC_703/Y INVX1_LOC_292/Y 0.23fF
C24572 NOR2X1_LOC_88/Y INVX1_LOC_49/Y 0.03fF
C24573 INVX1_LOC_35/A NOR2X1_LOC_114/A 0.01fF
C24574 NOR2X1_LOC_649/B INVX1_LOC_63/A 0.03fF
C24575 NAND2X1_LOC_568/a_36_24# NAND2X1_LOC_354/B 0.00fF
C24576 NOR2X1_LOC_355/A INVX1_LOC_161/Y 0.14fF
C24577 NAND2X1_LOC_740/Y INPUT_0 0.03fF
C24578 INVX1_LOC_50/A NOR2X1_LOC_486/Y 0.38fF
C24579 NOR2X1_LOC_89/A INVX1_LOC_131/Y 0.00fF
C24580 INVX1_LOC_3/A INVX1_LOC_63/A 0.03fF
C24581 NOR2X1_LOC_180/Y NOR2X1_LOC_550/B 0.09fF
C24582 NOR2X1_LOC_654/a_36_216# NOR2X1_LOC_661/A 0.02fF
C24583 NAND2X1_LOC_447/Y NOR2X1_LOC_383/B 0.03fF
C24584 INVX1_LOC_247/Y NOR2X1_LOC_500/Y 0.02fF
C24585 INVX1_LOC_29/A NOR2X1_LOC_445/B 0.20fF
C24586 NOR2X1_LOC_558/A INVX1_LOC_26/A 0.01fF
C24587 NOR2X1_LOC_635/A NAND2X1_LOC_21/Y 0.02fF
C24588 NOR2X1_LOC_78/B INVX1_LOC_94/A 0.39fF
C24589 INVX1_LOC_35/A INVX1_LOC_91/A 3.03fF
C24590 INVX1_LOC_12/A NOR2X1_LOC_58/Y 0.02fF
C24591 NAND2X1_LOC_287/B NOR2X1_LOC_318/A 0.02fF
C24592 D_INPUT_1 NOR2X1_LOC_124/A 0.05fF
C24593 INVX1_LOC_54/Y INVX1_LOC_77/A 0.07fF
C24594 D_INPUT_1 INVX1_LOC_188/Y 0.02fF
C24595 INVX1_LOC_290/A NAND2X1_LOC_195/Y -0.00fF
C24596 NAND2X1_LOC_559/Y NOR2X1_LOC_380/Y 0.04fF
C24597 NOR2X1_LOC_168/B INVX1_LOC_49/A 0.00fF
C24598 NAND2X1_LOC_796/a_36_24# NAND2X1_LOC_783/A 0.00fF
C24599 INVX1_LOC_36/A NOR2X1_LOC_440/Y 0.05fF
C24600 INVX1_LOC_279/A INVX1_LOC_30/A 0.26fF
C24601 NOR2X1_LOC_677/Y INVX1_LOC_20/A 0.05fF
C24602 INVX1_LOC_278/Y INVX1_LOC_41/Y 0.01fF
C24603 INVX1_LOC_58/A NAND2X1_LOC_469/B 0.03fF
C24604 INVX1_LOC_84/A INVX1_LOC_49/Y 0.03fF
C24605 INVX1_LOC_45/A INVX1_LOC_227/A 0.01fF
C24606 INVX1_LOC_11/A NAND2X1_LOC_807/Y 0.17fF
C24607 INVX1_LOC_271/A INVX1_LOC_76/A 2.02fF
C24608 INVX1_LOC_200/Y NAND2X1_LOC_244/A 0.03fF
C24609 INVX1_LOC_45/A NOR2X1_LOC_763/Y 0.04fF
C24610 INVX1_LOC_2/A NOR2X1_LOC_219/B 0.03fF
C24611 NAND2X1_LOC_571/B NOR2X1_LOC_24/Y 0.04fF
C24612 INVX1_LOC_39/Y INPUT_1 0.01fF
C24613 NOR2X1_LOC_23/a_36_216# NOR2X1_LOC_671/Y 0.00fF
C24614 NOR2X1_LOC_787/a_36_216# INVX1_LOC_182/A 0.01fF
C24615 INVX1_LOC_279/Y INVX1_LOC_196/Y 0.01fF
C24616 INVX1_LOC_2/A INVX1_LOC_88/Y 0.00fF
C24617 NOR2X1_LOC_773/Y NAND2X1_LOC_833/Y 0.01fF
C24618 INVX1_LOC_269/A NOR2X1_LOC_188/A 0.29fF
C24619 NOR2X1_LOC_218/A INVX1_LOC_75/A 0.04fF
C24620 NOR2X1_LOC_13/Y NAND2X1_LOC_660/Y 0.01fF
C24621 NOR2X1_LOC_567/a_36_216# INVX1_LOC_58/Y 0.01fF
C24622 NOR2X1_LOC_220/B NOR2X1_LOC_405/A 0.03fF
C24623 NOR2X1_LOC_818/Y NAND2X1_LOC_847/a_36_24# 0.00fF
C24624 INVX1_LOC_57/A INVX1_LOC_77/Y 0.07fF
C24625 INVX1_LOC_64/A NAND2X1_LOC_440/a_36_24# 0.00fF
C24626 INVX1_LOC_49/A NAND2X1_LOC_349/a_36_24# 0.00fF
C24627 INVX1_LOC_269/A NOR2X1_LOC_548/B 0.01fF
C24628 INVX1_LOC_104/A NOR2X1_LOC_537/Y 3.27fF
C24629 NOR2X1_LOC_599/A NAND2X1_LOC_644/a_36_24# 0.00fF
C24630 NOR2X1_LOC_266/B NOR2X1_LOC_717/A 0.00fF
C24631 INVX1_LOC_25/A INVX1_LOC_12/Y 0.10fF
C24632 INVX1_LOC_88/A INVX1_LOC_285/Y 0.01fF
C24633 INVX1_LOC_191/Y NOR2X1_LOC_52/B 0.01fF
C24634 NOR2X1_LOC_496/Y NAND2X1_LOC_623/B 0.18fF
C24635 INVX1_LOC_124/A INVX1_LOC_54/Y 0.47fF
C24636 NOR2X1_LOC_667/A NAND2X1_LOC_357/B 0.15fF
C24637 INVX1_LOC_227/A INVX1_LOC_71/A 0.69fF
C24638 INVX1_LOC_1/A NOR2X1_LOC_741/A 0.03fF
C24639 NAND2X1_LOC_470/B NOR2X1_LOC_435/A 0.02fF
C24640 NAND2X1_LOC_733/Y NAND2X1_LOC_560/A 0.13fF
C24641 NAND2X1_LOC_708/Y VDD 0.23fF
C24642 INVX1_LOC_226/Y INVX1_LOC_8/A 0.19fF
C24643 INVX1_LOC_45/A NOR2X1_LOC_703/A 0.03fF
C24644 INVX1_LOC_11/A INVX1_LOC_6/A 0.82fF
C24645 INVX1_LOC_177/Y INVX1_LOC_313/Y 0.92fF
C24646 NOR2X1_LOC_772/B NAND2X1_LOC_267/B 0.01fF
C24647 NAND2X1_LOC_569/A INVX1_LOC_16/A 0.01fF
C24648 INVX1_LOC_12/A INVX1_LOC_29/A 0.10fF
C24649 NAND2X1_LOC_214/B INVX1_LOC_76/A 0.00fF
C24650 NOR2X1_LOC_317/B NOR2X1_LOC_374/B 0.01fF
C24651 D_INPUT_0 NOR2X1_LOC_13/Y 0.01fF
C24652 NAND2X1_LOC_35/Y INVX1_LOC_46/A 0.20fF
C24653 NOR2X1_LOC_68/A D_GATE_366 0.07fF
C24654 NOR2X1_LOC_203/Y INVX1_LOC_177/A 0.01fF
C24655 NOR2X1_LOC_299/Y NAND2X1_LOC_866/A 0.15fF
C24656 INVX1_LOC_14/A INVX1_LOC_98/A 0.03fF
C24657 INVX1_LOC_182/Y INVX1_LOC_30/A 0.03fF
C24658 INVX1_LOC_280/A NOR2X1_LOC_414/Y 0.03fF
C24659 NOR2X1_LOC_798/A NOR2X1_LOC_538/a_36_216# 0.00fF
C24660 INVX1_LOC_298/Y INVX1_LOC_307/A 0.03fF
C24661 INVX1_LOC_286/A NAND2X1_LOC_793/Y 0.46fF
C24662 INVX1_LOC_176/A NOR2X1_LOC_849/A 0.03fF
C24663 INVX1_LOC_49/A NAND2X1_LOC_656/Y 0.05fF
C24664 INVX1_LOC_14/A NOR2X1_LOC_78/A 0.12fF
C24665 NOR2X1_LOC_824/A NOR2X1_LOC_824/Y 0.05fF
C24666 NOR2X1_LOC_68/A NOR2X1_LOC_750/A 0.32fF
C24667 INVX1_LOC_13/Y NAND2X1_LOC_267/B 0.09fF
C24668 INVX1_LOC_182/A INVX1_LOC_18/A 0.07fF
C24669 NAND2X1_LOC_510/A INVX1_LOC_75/A 0.04fF
C24670 NAND2X1_LOC_363/B NOR2X1_LOC_98/B 0.03fF
C24671 INVX1_LOC_27/A INVX1_LOC_76/A 0.16fF
C24672 NOR2X1_LOC_631/A INVX1_LOC_4/A 0.37fF
C24673 D_INPUT_0 NAND2X1_LOC_364/Y 0.07fF
C24674 NOR2X1_LOC_433/A INVX1_LOC_313/A 0.01fF
C24675 NOR2X1_LOC_78/B NOR2X1_LOC_136/Y 0.03fF
C24676 NOR2X1_LOC_440/Y NOR2X1_LOC_309/Y 0.03fF
C24677 NAND2X1_LOC_859/Y NOR2X1_LOC_52/B 2.58fF
C24678 NOR2X1_LOC_664/Y INVX1_LOC_7/A 0.05fF
C24679 INVX1_LOC_49/Y INVX1_LOC_15/A 0.03fF
C24680 NAND2X1_LOC_858/B INVX1_LOC_30/A 0.00fF
C24681 NOR2X1_LOC_791/B NAND2X1_LOC_348/A 0.00fF
C24682 NAND2X1_LOC_361/Y INVX1_LOC_89/A 0.25fF
C24683 NAND2X1_LOC_753/a_36_24# INVX1_LOC_9/A 0.01fF
C24684 NAND2X1_LOC_799/A INVX1_LOC_291/Y 0.03fF
C24685 INVX1_LOC_211/A NOR2X1_LOC_45/B 0.08fF
C24686 INVX1_LOC_49/A NAND2X1_LOC_638/Y 0.06fF
C24687 INVX1_LOC_239/A D_GATE_479 0.02fF
C24688 INVX1_LOC_77/A NOR2X1_LOC_112/Y 0.03fF
C24689 NOR2X1_LOC_769/B INVX1_LOC_92/A 0.01fF
C24690 INVX1_LOC_95/A NAND2X1_LOC_793/Y 0.06fF
C24691 INVX1_LOC_225/Y NOR2X1_LOC_405/A 0.19fF
C24692 NAND2X1_LOC_223/B INVX1_LOC_3/A 0.01fF
C24693 NAND2X1_LOC_618/Y NAND2X1_LOC_82/Y 0.15fF
C24694 VDD INVX1_LOC_198/A 0.02fF
C24695 VDD NOR2X1_LOC_271/B 0.08fF
C24696 NOR2X1_LOC_598/B INVX1_LOC_92/A 0.45fF
C24697 NOR2X1_LOC_13/Y NAND2X1_LOC_538/a_36_24# 0.00fF
C24698 NAND2X1_LOC_785/A NAND2X1_LOC_862/a_36_24# 0.00fF
C24699 INVX1_LOC_41/A NAND2X1_LOC_842/B 0.16fF
C24700 INVX1_LOC_28/A INVX1_LOC_155/A 0.09fF
C24701 INVX1_LOC_34/A NOR2X1_LOC_597/A 0.01fF
C24702 NOR2X1_LOC_111/Y NOR2X1_LOC_172/Y 0.06fF
C24703 NOR2X1_LOC_479/B INVX1_LOC_255/Y 0.02fF
C24704 INVX1_LOC_53/A NOR2X1_LOC_155/A 0.11fF
C24705 NOR2X1_LOC_52/B INVX1_LOC_313/A 0.08fF
C24706 NAND2X1_LOC_560/A NAND2X1_LOC_787/B 0.03fF
C24707 NAND2X1_LOC_222/a_36_24# NOR2X1_LOC_814/A 0.00fF
C24708 INVX1_LOC_208/A INVX1_LOC_290/A 0.02fF
C24709 NAND2X1_LOC_175/Y INVX1_LOC_264/A 0.10fF
C24710 INVX1_LOC_1/A INVX1_LOC_12/Y 0.19fF
C24711 NOR2X1_LOC_740/Y VDD 0.31fF
C24712 INVX1_LOC_104/A INVX1_LOC_313/Y 0.00fF
C24713 NAND2X1_LOC_833/Y INVX1_LOC_140/A 0.24fF
C24714 NAND2X1_LOC_838/Y NAND2X1_LOC_866/B 0.08fF
C24715 NOR2X1_LOC_278/a_36_216# INVX1_LOC_256/Y 0.00fF
C24716 NOR2X1_LOC_299/Y NOR2X1_LOC_505/Y 0.04fF
C24717 INVX1_LOC_136/A NOR2X1_LOC_45/B 0.20fF
C24718 INVX1_LOC_254/Y INPUT_0 0.22fF
C24719 NOR2X1_LOC_565/a_36_216# NOR2X1_LOC_550/B 0.02fF
C24720 INVX1_LOC_65/A NOR2X1_LOC_500/B 0.44fF
C24721 INVX1_LOC_31/A INVX1_LOC_74/A 0.03fF
C24722 NOR2X1_LOC_52/B NAND2X1_LOC_807/Y 0.07fF
C24723 INVX1_LOC_150/Y VDD 0.98fF
C24724 INVX1_LOC_298/Y INVX1_LOC_12/A 0.03fF
C24725 INVX1_LOC_161/Y NOR2X1_LOC_111/A 0.01fF
C24726 NOR2X1_LOC_68/A NOR2X1_LOC_746/Y 0.10fF
C24727 NOR2X1_LOC_218/Y NAND2X1_LOC_656/Y 0.02fF
C24728 NOR2X1_LOC_433/A INVX1_LOC_6/A 0.11fF
C24729 NOR2X1_LOC_173/Y INVX1_LOC_54/A 0.10fF
C24730 INVX1_LOC_7/A INVX1_LOC_137/A 0.01fF
C24731 NAND2X1_LOC_348/A NOR2X1_LOC_124/B 0.00fF
C24732 NOR2X1_LOC_321/Y INVX1_LOC_54/A 0.02fF
C24733 NOR2X1_LOC_82/Y NOR2X1_LOC_123/B 0.01fF
C24734 INVX1_LOC_136/A INVX1_LOC_247/A 0.03fF
C24735 NAND2X1_LOC_728/Y INVX1_LOC_291/Y 0.02fF
C24736 INVX1_LOC_240/A INVX1_LOC_282/A 0.10fF
C24737 INVX1_LOC_49/A INVX1_LOC_78/Y 0.03fF
C24738 NOR2X1_LOC_593/Y INVX1_LOC_6/A 0.01fF
C24739 NOR2X1_LOC_471/Y NAND2X1_LOC_472/Y 0.01fF
C24740 NAND2X1_LOC_84/Y NOR2X1_LOC_78/A 0.01fF
C24741 NOR2X1_LOC_646/a_36_216# INVX1_LOC_135/A 0.00fF
C24742 NOR2X1_LOC_91/A NAND2X1_LOC_254/Y 0.07fF
C24743 INVX1_LOC_263/A INVX1_LOC_313/Y 0.00fF
C24744 NOR2X1_LOC_89/A INVX1_LOC_270/A 0.03fF
C24745 NAND2X1_LOC_803/B NOR2X1_LOC_331/B 0.03fF
C24746 NOR2X1_LOC_562/B INVX1_LOC_113/Y 0.13fF
C24747 INVX1_LOC_312/A NOR2X1_LOC_111/A 0.03fF
C24748 INVX1_LOC_254/A NAND2X1_LOC_642/Y 0.15fF
C24749 NOR2X1_LOC_92/Y NAND2X1_LOC_243/B 0.05fF
C24750 NOR2X1_LOC_299/Y NOR2X1_LOC_700/Y 0.07fF
C24751 INVX1_LOC_303/A INVX1_LOC_65/A 0.03fF
C24752 NOR2X1_LOC_52/B INVX1_LOC_6/A 2.97fF
C24753 NAND2X1_LOC_452/Y NAND2X1_LOC_470/B 0.02fF
C24754 NAND2X1_LOC_140/A INVX1_LOC_10/A 0.02fF
C24755 NOR2X1_LOC_773/Y INVX1_LOC_73/A 0.46fF
C24756 INVX1_LOC_138/Y INVX1_LOC_19/A 0.07fF
C24757 NAND2X1_LOC_793/Y INVX1_LOC_54/A 0.01fF
C24758 NAND2X1_LOC_254/Y INVX1_LOC_23/A 0.11fF
C24759 NOR2X1_LOC_78/B INVX1_LOC_144/A 0.07fF
C24760 INVX1_LOC_229/Y INVX1_LOC_173/Y 0.32fF
C24761 INVX1_LOC_78/A NOR2X1_LOC_464/Y 0.04fF
C24762 INVX1_LOC_249/A INVX1_LOC_76/A 0.09fF
C24763 INVX1_LOC_32/A NOR2X1_LOC_646/B 0.01fF
C24764 INVX1_LOC_94/A INVX1_LOC_46/A 0.07fF
C24765 NOR2X1_LOC_646/A NAND2X1_LOC_348/A 0.09fF
C24766 NOR2X1_LOC_717/B NOR2X1_LOC_828/A 1.07fF
C24767 NOR2X1_LOC_431/Y NAND2X1_LOC_453/A 0.01fF
C24768 INVX1_LOC_41/A NOR2X1_LOC_545/B 0.01fF
C24769 INVX1_LOC_233/A INVX1_LOC_168/Y 0.01fF
C24770 INVX1_LOC_165/A INVX1_LOC_23/Y 0.03fF
C24771 INVX1_LOC_7/A NOR2X1_LOC_19/B 0.06fF
C24772 NOR2X1_LOC_89/A NOR2X1_LOC_109/Y 0.28fF
C24773 NOR2X1_LOC_521/Y NAND2X1_LOC_849/A 0.10fF
C24774 NOR2X1_LOC_272/Y INVX1_LOC_19/A 0.03fF
C24775 NAND2X1_LOC_803/B NOR2X1_LOC_592/B 0.02fF
C24776 D_INPUT_7 INVX1_LOC_38/A 0.01fF
C24777 INVX1_LOC_13/Y NAND2X1_LOC_81/B 0.04fF
C24778 NOR2X1_LOC_510/Y INVX1_LOC_272/A 0.07fF
C24779 INVX1_LOC_312/Y INVX1_LOC_118/A 0.10fF
C24780 NAND2X1_LOC_670/a_36_24# INVX1_LOC_9/A 0.00fF
C24781 INVX1_LOC_166/A INVX1_LOC_253/A 0.11fF
C24782 NOR2X1_LOC_716/B NAND2X1_LOC_633/Y 0.78fF
C24783 NOR2X1_LOC_264/Y NOR2X1_LOC_35/Y 0.10fF
C24784 NOR2X1_LOC_400/B NOR2X1_LOC_415/Y 0.01fF
C24785 INVX1_LOC_166/A INVX1_LOC_90/Y 0.02fF
C24786 INVX1_LOC_34/A NOR2X1_LOC_825/Y 0.10fF
C24787 NOR2X1_LOC_554/B NOR2X1_LOC_54/a_36_216# 0.00fF
C24788 NOR2X1_LOC_848/Y NOR2X1_LOC_814/A 0.00fF
C24789 NOR2X1_LOC_693/Y INVX1_LOC_23/Y 0.01fF
C24790 NAND2X1_LOC_16/Y INVX1_LOC_54/A 0.01fF
C24791 NOR2X1_LOC_717/B NOR2X1_LOC_151/Y 0.01fF
C24792 INVX1_LOC_17/A NAND2X1_LOC_206/Y 0.07fF
C24793 INVX1_LOC_140/A NOR2X1_LOC_76/A 0.29fF
C24794 D_INPUT_7 NOR2X1_LOC_51/A 0.33fF
C24795 NAND2X1_LOC_462/B NAND2X1_LOC_622/B 0.02fF
C24796 NOR2X1_LOC_322/Y NAND2X1_LOC_861/Y 0.10fF
C24797 INVX1_LOC_239/A INVX1_LOC_167/A 0.04fF
C24798 INVX1_LOC_83/A INVX1_LOC_144/A 0.10fF
C24799 NOR2X1_LOC_773/Y NAND2X1_LOC_729/B 0.04fF
C24800 INVX1_LOC_27/A NAND2X1_LOC_202/a_36_24# 0.00fF
C24801 NOR2X1_LOC_637/A INVX1_LOC_54/A 0.01fF
C24802 NOR2X1_LOC_500/A INVX1_LOC_9/A 0.01fF
C24803 INVX1_LOC_256/A INVX1_LOC_63/A 1.08fF
C24804 INVX1_LOC_113/Y INVX1_LOC_281/Y 0.01fF
C24805 NOR2X1_LOC_441/Y NOR2X1_LOC_127/a_36_216# 0.00fF
C24806 NOR2X1_LOC_303/Y INVX1_LOC_9/A 0.12fF
C24807 INVX1_LOC_63/Y INVX1_LOC_117/A 0.12fF
C24808 NOR2X1_LOC_92/Y INVX1_LOC_284/A 0.85fF
C24809 NOR2X1_LOC_647/B INVX1_LOC_63/A 0.00fF
C24810 NOR2X1_LOC_647/A NAND2X1_LOC_215/A 0.01fF
C24811 INVX1_LOC_247/Y INVX1_LOC_307/A 0.01fF
C24812 NOR2X1_LOC_828/A NOR2X1_LOC_151/Y 0.01fF
C24813 NOR2X1_LOC_361/B INVX1_LOC_272/A 0.04fF
C24814 INVX1_LOC_27/A INVX1_LOC_127/Y 0.02fF
C24815 NOR2X1_LOC_772/B INVX1_LOC_4/Y 0.07fF
C24816 NOR2X1_LOC_188/Y INVX1_LOC_91/A 0.05fF
C24817 INVX1_LOC_50/A NOR2X1_LOC_748/A 0.06fF
C24818 INVX1_LOC_200/A INVX1_LOC_29/A 0.01fF
C24819 VDD NOR2X1_LOC_87/Y 0.24fF
C24820 NAND2X1_LOC_364/A NAND2X1_LOC_288/A 0.10fF
C24821 NOR2X1_LOC_791/Y NOR2X1_LOC_38/B 0.03fF
C24822 INVX1_LOC_192/A INVX1_LOC_38/A 0.01fF
C24823 INVX1_LOC_13/Y INVX1_LOC_4/Y 0.95fF
C24824 INVX1_LOC_256/Y NOR2X1_LOC_266/B 0.01fF
C24825 NOR2X1_LOC_254/Y INVX1_LOC_9/A 0.05fF
C24826 NOR2X1_LOC_289/Y INVX1_LOC_147/A 0.01fF
C24827 NAND2X1_LOC_483/Y INVX1_LOC_118/A 0.05fF
C24828 INVX1_LOC_1/A NOR2X1_LOC_554/A 0.01fF
C24829 NAND2X1_LOC_793/Y NAND2X1_LOC_807/B 0.13fF
C24830 NOR2X1_LOC_433/A INVX1_LOC_131/Y 0.04fF
C24831 INVX1_LOC_77/A NAND2X1_LOC_656/B 0.01fF
C24832 INVX1_LOC_206/Y INVX1_LOC_313/Y 0.07fF
C24833 NOR2X1_LOC_593/Y NOR2X1_LOC_79/A 0.27fF
C24834 NOR2X1_LOC_99/B NAND2X1_LOC_86/Y 0.04fF
C24835 NOR2X1_LOC_716/B INVX1_LOC_71/Y 0.04fF
C24836 NOR2X1_LOC_336/B INVX1_LOC_19/A 0.01fF
C24837 INVX1_LOC_64/A NOR2X1_LOC_677/Y 0.05fF
C24838 INVX1_LOC_290/A NAND2X1_LOC_211/Y 0.44fF
C24839 NOR2X1_LOC_717/B NOR2X1_LOC_181/A 0.00fF
C24840 NOR2X1_LOC_561/Y NOR2X1_LOC_314/a_36_216# 0.01fF
C24841 NOR2X1_LOC_722/a_36_216# INVX1_LOC_179/A 0.00fF
C24842 NOR2X1_LOC_598/B INVX1_LOC_53/A 0.27fF
C24843 NOR2X1_LOC_353/Y INVX1_LOC_9/A 0.05fF
C24844 INVX1_LOC_31/A NAND2X1_LOC_254/Y 0.03fF
C24845 INVX1_LOC_174/A NAND2X1_LOC_430/B 0.05fF
C24846 INVX1_LOC_313/Y NOR2X1_LOC_600/Y 0.01fF
C24847 NAND2X1_LOC_364/A INVX1_LOC_19/A 0.12fF
C24848 INVX1_LOC_299/A NOR2X1_LOC_334/Y 0.11fF
C24849 INVX1_LOC_50/A NOR2X1_LOC_304/Y 0.01fF
C24850 NOR2X1_LOC_247/Y NOR2X1_LOC_342/A 0.01fF
C24851 NOR2X1_LOC_543/A INVX1_LOC_14/Y 0.25fF
C24852 INVX1_LOC_34/A NOR2X1_LOC_88/Y 0.01fF
C24853 INVX1_LOC_36/A NOR2X1_LOC_89/A 0.43fF
C24854 NOR2X1_LOC_82/a_36_216# INVX1_LOC_12/A 0.02fF
C24855 NAND2X1_LOC_9/Y NAND2X1_LOC_35/Y 0.60fF
C24856 INVX1_LOC_124/A NAND2X1_LOC_656/B 0.01fF
C24857 INVX1_LOC_57/Y NOR2X1_LOC_46/a_36_216# 0.00fF
C24858 NOR2X1_LOC_160/B NOR2X1_LOC_801/B 0.07fF
C24859 INVX1_LOC_1/Y NOR2X1_LOC_536/A 0.04fF
C24860 NOR2X1_LOC_156/B INVX1_LOC_92/A 0.15fF
C24861 NOR2X1_LOC_267/A NOR2X1_LOC_89/A 0.44fF
C24862 NOR2X1_LOC_632/Y INVX1_LOC_44/A 0.00fF
C24863 INVX1_LOC_243/Y NAND2X1_LOC_149/Y 0.05fF
C24864 NOR2X1_LOC_140/a_36_216# NAND2X1_LOC_574/A 0.01fF
C24865 INVX1_LOC_82/A NAND2X1_LOC_141/Y 0.03fF
C24866 NOR2X1_LOC_568/A NOR2X1_LOC_169/a_36_216# 0.01fF
C24867 NOR2X1_LOC_646/a_36_216# INVX1_LOC_280/A 0.00fF
C24868 INVX1_LOC_34/A INVX1_LOC_84/A 2.51fF
C24869 NOR2X1_LOC_67/A NOR2X1_LOC_235/Y 0.03fF
C24870 INVX1_LOC_90/A INVX1_LOC_2/Y 0.00fF
C24871 INVX1_LOC_50/Y NOR2X1_LOC_678/A 0.02fF
C24872 NOR2X1_LOC_295/Y NAND2X1_LOC_475/Y 0.08fF
C24873 INVX1_LOC_228/A INVX1_LOC_12/A 0.08fF
C24874 NOR2X1_LOC_68/A NAND2X1_LOC_295/a_36_24# 0.00fF
C24875 INVX1_LOC_55/Y NOR2X1_LOC_357/Y 0.07fF
C24876 NOR2X1_LOC_528/Y NOR2X1_LOC_167/Y 0.05fF
C24877 NOR2X1_LOC_457/B INVX1_LOC_42/A 0.01fF
C24878 NOR2X1_LOC_78/B NOR2X1_LOC_155/A 0.10fF
C24879 INVX1_LOC_145/A NOR2X1_LOC_89/A 0.31fF
C24880 NOR2X1_LOC_151/Y NOR2X1_LOC_181/A 0.05fF
C24881 NOR2X1_LOC_208/Y NOR2X1_LOC_89/A 0.07fF
C24882 INVX1_LOC_17/A NOR2X1_LOC_639/Y 0.04fF
C24883 NAND2X1_LOC_837/Y INVX1_LOC_284/A 0.08fF
C24884 NAND2X1_LOC_383/a_36_24# NAND2X1_LOC_725/B 0.01fF
C24885 NOR2X1_LOC_19/B INVX1_LOC_76/A 0.08fF
C24886 NAND2X1_LOC_148/a_36_24# INVX1_LOC_193/A 0.00fF
C24887 NOR2X1_LOC_385/Y INVX1_LOC_20/A 0.27fF
C24888 NOR2X1_LOC_356/A INVX1_LOC_37/A 0.07fF
C24889 NAND2X1_LOC_350/A NAND2X1_LOC_466/a_36_24# 0.01fF
C24890 NOR2X1_LOC_617/a_36_216# NAND2X1_LOC_254/Y 0.00fF
C24891 NOR2X1_LOC_78/A INVX1_LOC_48/A 0.74fF
C24892 INVX1_LOC_93/Y INVX1_LOC_126/Y 0.02fF
C24893 NAND2X1_LOC_725/Y INVX1_LOC_269/A 0.01fF
C24894 D_INPUT_1 NOR2X1_LOC_15/Y 0.07fF
C24895 NOR2X1_LOC_237/Y NOR2X1_LOC_89/A 0.29fF
C24896 INVX1_LOC_1/Y NAND2X1_LOC_93/B 6.73fF
C24897 INVX1_LOC_286/Y NOR2X1_LOC_409/B 0.03fF
C24898 NOR2X1_LOC_160/B INVX1_LOC_116/Y 0.01fF
C24899 NOR2X1_LOC_92/Y NAND2X1_LOC_627/a_36_24# 0.01fF
C24900 NOR2X1_LOC_178/Y INVX1_LOC_27/A 0.04fF
C24901 NAND2X1_LOC_656/Y INVX1_LOC_118/A 0.02fF
C24902 INVX1_LOC_71/A NOR2X1_LOC_169/a_36_216# 0.00fF
C24903 NAND2X1_LOC_858/a_36_24# NOR2X1_LOC_88/Y 0.01fF
C24904 NAND2X1_LOC_787/A NOR2X1_LOC_468/Y 0.04fF
C24905 NAND2X1_LOC_162/A INVX1_LOC_107/Y 0.02fF
C24906 NOR2X1_LOC_686/B INVX1_LOC_54/A 0.02fF
C24907 INVX1_LOC_199/A INVX1_LOC_6/A 0.01fF
C24908 NAND2X1_LOC_348/A INVX1_LOC_2/Y 0.08fF
C24909 NOR2X1_LOC_719/A NOR2X1_LOC_216/B 0.12fF
C24910 INVX1_LOC_21/A NOR2X1_LOC_291/Y 0.01fF
C24911 INVX1_LOC_8/A INVX1_LOC_12/A 0.07fF
C24912 NOR2X1_LOC_689/Y NAND2X1_LOC_727/a_36_24# 0.00fF
C24913 NOR2X1_LOC_589/A NOR2X1_LOC_831/B 0.07fF
C24914 INVX1_LOC_27/A NOR2X1_LOC_34/B 0.02fF
C24915 INVX1_LOC_144/A INVX1_LOC_46/A 0.23fF
C24916 INVX1_LOC_157/A NOR2X1_LOC_435/A 0.33fF
C24917 INVX1_LOC_168/A NAND2X1_LOC_81/B 0.03fF
C24918 NOR2X1_LOC_74/A INVX1_LOC_37/A 0.22fF
C24919 NOR2X1_LOC_595/Y NAND2X1_LOC_655/A 0.00fF
C24920 NOR2X1_LOC_561/Y NOR2X1_LOC_216/B 0.03fF
C24921 NOR2X1_LOC_336/B INVX1_LOC_26/Y 0.03fF
C24922 NOR2X1_LOC_309/Y NOR2X1_LOC_89/A 0.11fF
C24923 NOR2X1_LOC_83/Y INVX1_LOC_46/A 0.14fF
C24924 INVX1_LOC_25/A NOR2X1_LOC_160/B 0.24fF
C24925 NOR2X1_LOC_457/B INVX1_LOC_78/A 0.40fF
C24926 INVX1_LOC_50/A NAND2X1_LOC_711/Y 0.01fF
C24927 INVX1_LOC_64/A NOR2X1_LOC_533/Y 0.03fF
C24928 NOR2X1_LOC_112/Y INVX1_LOC_9/A 0.16fF
C24929 INVX1_LOC_83/A NOR2X1_LOC_155/A 0.06fF
C24930 NAND2X1_LOC_112/Y NOR2X1_LOC_127/Y 0.09fF
C24931 NOR2X1_LOC_9/Y INVX1_LOC_37/A 0.03fF
C24932 NOR2X1_LOC_15/Y NOR2X1_LOC_652/Y 0.06fF
C24933 NAND2X1_LOC_11/Y NOR2X1_LOC_11/Y 0.00fF
C24934 NOR2X1_LOC_836/Y NOR2X1_LOC_836/a_36_216# 0.03fF
C24935 NOR2X1_LOC_9/Y NOR2X1_LOC_231/A 0.01fF
C24936 INVX1_LOC_11/A NOR2X1_LOC_109/Y 0.07fF
C24937 INVX1_LOC_303/A INVX1_LOC_4/Y 0.10fF
C24938 NAND2X1_LOC_364/A INVX1_LOC_26/Y 0.04fF
C24939 INVX1_LOC_16/A NOR2X1_LOC_662/A 0.10fF
C24940 INVX1_LOC_34/A INVX1_LOC_15/A 0.29fF
C24941 NOR2X1_LOC_186/Y INVX1_LOC_14/A 0.08fF
C24942 D_INPUT_0 NAND2X1_LOC_94/a_36_24# 0.00fF
C24943 INVX1_LOC_181/Y INVX1_LOC_26/A 0.08fF
C24944 NOR2X1_LOC_290/Y NAND2X1_LOC_254/Y 0.01fF
C24945 INVX1_LOC_58/A NAND2X1_LOC_154/Y 0.01fF
C24946 NAND2X1_LOC_360/a_36_24# NOR2X1_LOC_160/B 0.00fF
C24947 INVX1_LOC_135/A INVX1_LOC_285/A 0.10fF
C24948 INVX1_LOC_24/A NOR2X1_LOC_302/A 0.01fF
C24949 INVX1_LOC_135/A INVX1_LOC_265/Y 0.61fF
C24950 NOR2X1_LOC_346/Y NOR2X1_LOC_35/Y 0.05fF
C24951 NOR2X1_LOC_315/a_36_216# INVX1_LOC_12/A 0.00fF
C24952 NAND2X1_LOC_573/Y INVX1_LOC_14/A 0.15fF
C24953 INVX1_LOC_135/A NOR2X1_LOC_814/A 9.37fF
C24954 NOR2X1_LOC_272/Y INVX1_LOC_161/Y 0.10fF
C24955 NAND2X1_LOC_569/B NAND2X1_LOC_577/A 0.03fF
C24956 INVX1_LOC_21/A NOR2X1_LOC_745/Y 0.01fF
C24957 NAND2X1_LOC_231/Y INVX1_LOC_15/A 0.01fF
C24958 INVX1_LOC_49/A NOR2X1_LOC_727/B 0.03fF
C24959 NOR2X1_LOC_318/B NOR2X1_LOC_536/A 0.05fF
C24960 NOR2X1_LOC_248/a_36_216# INVX1_LOC_285/A 0.00fF
C24961 NOR2X1_LOC_591/Y INVX1_LOC_273/A 0.02fF
C24962 NOR2X1_LOC_205/Y INVX1_LOC_88/A 0.03fF
C24963 NAND2X1_LOC_348/A NOR2X1_LOC_608/Y 0.00fF
C24964 NOR2X1_LOC_816/a_36_216# INVX1_LOC_31/A 0.00fF
C24965 INVX1_LOC_39/A INVX1_LOC_39/Y 0.01fF
C24966 NOR2X1_LOC_808/A NOR2X1_LOC_855/A 0.05fF
C24967 INVX1_LOC_2/A INVX1_LOC_128/Y 0.20fF
C24968 NAND2X1_LOC_859/Y NAND2X1_LOC_254/Y 0.03fF
C24969 INVX1_LOC_93/Y NOR2X1_LOC_536/A 0.07fF
C24970 NAND2X1_LOC_190/Y NOR2X1_LOC_457/A 0.10fF
C24971 NOR2X1_LOC_802/A INVX1_LOC_18/Y 0.09fF
C24972 INPUT_0 NOR2X1_LOC_88/Y 0.07fF
C24973 NOR2X1_LOC_250/a_36_216# NOR2X1_LOC_250/Y -0.00fF
C24974 INVX1_LOC_21/A NOR2X1_LOC_602/A 0.01fF
C24975 INVX1_LOC_236/A NAND2X1_LOC_175/Y 0.42fF
C24976 INVX1_LOC_28/A NOR2X1_LOC_662/A 0.10fF
C24977 NOR2X1_LOC_160/B INVX1_LOC_1/A 1.08fF
C24978 NAND2X1_LOC_796/B INVX1_LOC_57/Y 0.06fF
C24979 INVX1_LOC_305/A INVX1_LOC_50/Y 0.07fF
C24980 NOR2X1_LOC_846/Y NOR2X1_LOC_554/B 0.29fF
C24981 NOR2X1_LOC_772/Y INVX1_LOC_29/Y 0.00fF
C24982 INVX1_LOC_13/A INVX1_LOC_32/A 0.12fF
C24983 INVX1_LOC_58/A INVX1_LOC_63/Y 0.14fF
C24984 INVX1_LOC_77/A NOR2X1_LOC_634/Y 0.00fF
C24985 INVX1_LOC_59/A NOR2X1_LOC_382/Y 0.04fF
C24986 NOR2X1_LOC_709/A NAND2X1_LOC_99/A 0.17fF
C24987 INVX1_LOC_41/A NAND2X1_LOC_275/a_36_24# 0.00fF
C24988 NAND2X1_LOC_198/B INVX1_LOC_306/Y 0.10fF
C24989 NOR2X1_LOC_251/a_36_216# INVX1_LOC_45/A -0.00fF
C24990 NAND2X1_LOC_35/Y NAND2X1_LOC_866/A 1.98fF
C24991 NOR2X1_LOC_318/B NAND2X1_LOC_93/B 0.08fF
C24992 NOR2X1_LOC_52/B INVX1_LOC_270/A 1.97fF
C24993 NOR2X1_LOC_321/a_36_216# NOR2X1_LOC_334/Y 0.00fF
C24994 INVX1_LOC_21/A NOR2X1_LOC_546/A 0.38fF
C24995 INPUT_0 INVX1_LOC_84/A 0.24fF
C24996 NOR2X1_LOC_392/B INVX1_LOC_29/Y 0.01fF
C24997 NOR2X1_LOC_802/A NAND2X1_LOC_279/a_36_24# 0.00fF
C24998 NAND2X1_LOC_14/a_36_24# INVX1_LOC_32/A 0.00fF
C24999 NOR2X1_LOC_468/Y INVX1_LOC_30/A 0.61fF
C25000 NOR2X1_LOC_667/A NOR2X1_LOC_282/Y 0.01fF
C25001 NAND2X1_LOC_866/B NAND2X1_LOC_254/Y 0.07fF
C25002 NOR2X1_LOC_92/Y INVX1_LOC_72/A 0.17fF
C25003 NOR2X1_LOC_751/a_36_216# NAND2X1_LOC_364/A 0.00fF
C25004 INVX1_LOC_278/A INVX1_LOC_34/A 0.01fF
C25005 INVX1_LOC_93/Y NAND2X1_LOC_93/B 0.07fF
C25006 INVX1_LOC_2/Y INVX1_LOC_38/A 0.00fF
C25007 NAND2X1_LOC_222/B INVX1_LOC_36/A -0.00fF
C25008 NOR2X1_LOC_32/B NOR2X1_LOC_629/B 0.03fF
C25009 D_INPUT_1 NAND2X1_LOC_141/A 0.28fF
C25010 NAND2X1_LOC_579/A INVX1_LOC_18/A 0.78fF
C25011 NAND2X1_LOC_721/A NOR2X1_LOC_536/A 0.04fF
C25012 NOR2X1_LOC_246/A INVX1_LOC_32/A 0.10fF
C25013 INVX1_LOC_219/Y NOR2X1_LOC_392/Y 0.02fF
C25014 NOR2X1_LOC_689/A NAND2X1_LOC_724/a_36_24# 0.00fF
C25015 NAND2X1_LOC_182/A NAND2X1_LOC_793/B 0.14fF
C25016 NAND2X1_LOC_837/Y NOR2X1_LOC_384/A 0.07fF
C25017 INVX1_LOC_69/Y INVX1_LOC_63/A 0.07fF
C25018 NOR2X1_LOC_679/B NOR2X1_LOC_304/Y 0.03fF
C25019 INVX1_LOC_11/A INVX1_LOC_36/A 1.04fF
C25020 NAND2X1_LOC_656/A NAND2X1_LOC_218/A 0.06fF
C25021 NOR2X1_LOC_405/A NAND2X1_LOC_288/A 0.03fF
C25022 NAND2X1_LOC_577/A NOR2X1_LOC_530/Y 0.02fF
C25023 INVX1_LOC_201/Y NOR2X1_LOC_663/A 0.00fF
C25024 NOR2X1_LOC_78/B NOR2X1_LOC_125/Y 0.45fF
C25025 NOR2X1_LOC_174/B NOR2X1_LOC_623/B 0.03fF
C25026 NAND2X1_LOC_863/B NAND2X1_LOC_828/a_36_24# 0.01fF
C25027 NAND2X1_LOC_555/Y NAND2X1_LOC_37/a_36_24# 0.00fF
C25028 INVX1_LOC_238/A NAND2X1_LOC_733/Y 0.04fF
C25029 NOR2X1_LOC_778/B INVX1_LOC_23/A 0.07fF
C25030 NOR2X1_LOC_251/a_36_216# INVX1_LOC_71/A -0.02fF
C25031 VDD NOR2X1_LOC_612/Y 0.23fF
C25032 INVX1_LOC_200/A NAND2X1_LOC_634/Y 0.00fF
C25033 NOR2X1_LOC_52/B NOR2X1_LOC_109/Y 0.19fF
C25034 NAND2X1_LOC_785/A NAND2X1_LOC_790/a_36_24# 0.01fF
C25035 NAND2X1_LOC_740/Y NAND2X1_LOC_811/Y 0.15fF
C25036 NOR2X1_LOC_598/B NOR2X1_LOC_547/B 0.03fF
C25037 NOR2X1_LOC_598/B NOR2X1_LOC_78/B 0.13fF
C25038 NOR2X1_LOC_606/a_36_216# NOR2X1_LOC_606/Y 0.00fF
C25039 NOR2X1_LOC_389/A INVX1_LOC_30/A 0.01fF
C25040 INVX1_LOC_11/A NAND2X1_LOC_587/a_36_24# 0.00fF
C25041 NOR2X1_LOC_226/A NOR2X1_LOC_717/A 0.04fF
C25042 NOR2X1_LOC_216/B INVX1_LOC_76/A 0.07fF
C25043 INVX1_LOC_16/A INVX1_LOC_57/A 0.53fF
C25044 NOR2X1_LOC_749/a_36_216# INVX1_LOC_87/A 0.01fF
C25045 INVX1_LOC_172/A NAND2X1_LOC_579/A 0.07fF
C25046 INVX1_LOC_17/A INVX1_LOC_24/A 0.09fF
C25047 INVX1_LOC_37/A NOR2X1_LOC_650/a_36_216# 0.01fF
C25048 NOR2X1_LOC_373/Y NOR2X1_LOC_693/a_36_216# 0.00fF
C25049 NAND2X1_LOC_149/Y NAND2X1_LOC_686/a_36_24# 0.01fF
C25050 NOR2X1_LOC_76/A INVX1_LOC_78/A 0.11fF
C25051 INVX1_LOC_25/A NOR2X1_LOC_516/B 0.13fF
C25052 INVX1_LOC_237/Y INVX1_LOC_237/A 0.01fF
C25053 NOR2X1_LOC_246/A NAND2X1_LOC_175/Y 0.01fF
C25054 NAND2X1_LOC_734/B NOR2X1_LOC_406/A 0.10fF
C25055 NOR2X1_LOC_130/A NOR2X1_LOC_301/A 0.03fF
C25056 NAND2X1_LOC_199/B INVX1_LOC_30/A 0.04fF
C25057 NOR2X1_LOC_155/A INVX1_LOC_46/A 0.16fF
C25058 NAND2X1_LOC_767/a_36_24# NOR2X1_LOC_68/A 0.01fF
C25059 INVX1_LOC_97/Y NOR2X1_LOC_78/B 0.15fF
C25060 NOR2X1_LOC_761/Y NOR2X1_LOC_599/A 0.01fF
C25061 INVX1_LOC_58/A NAND2X1_LOC_848/a_36_24# 0.00fF
C25062 INVX1_LOC_11/A NOR2X1_LOC_208/Y 0.03fF
C25063 NOR2X1_LOC_637/A NAND2X1_LOC_350/A 0.09fF
C25064 NOR2X1_LOC_71/Y INVX1_LOC_23/Y 0.03fF
C25065 NAND2X1_LOC_797/a_36_24# NOR2X1_LOC_781/Y 0.00fF
C25066 INVX1_LOC_225/A NOR2X1_LOC_792/a_36_216# 0.00fF
C25067 NAND2X1_LOC_725/B INVX1_LOC_207/A 0.07fF
C25068 NAND2X1_LOC_569/A INVX1_LOC_48/Y 0.02fF
C25069 NOR2X1_LOC_356/A NAND2X1_LOC_72/B 0.00fF
C25070 NOR2X1_LOC_113/A INVX1_LOC_19/A 0.09fF
C25071 INVX1_LOC_37/A NOR2X1_LOC_865/Y 0.03fF
C25072 NOR2X1_LOC_471/Y INVX1_LOC_24/A 0.02fF
C25073 NOR2X1_LOC_405/A INVX1_LOC_19/A 0.09fF
C25074 INVX1_LOC_14/A NAND2X1_LOC_640/Y -0.02fF
C25075 INVX1_LOC_1/A NOR2X1_LOC_317/B 0.03fF
C25076 NAND2X1_LOC_541/a_36_24# INVX1_LOC_16/A 0.00fF
C25077 NOR2X1_LOC_570/A INVX1_LOC_53/A 0.03fF
C25078 NOR2X1_LOC_639/B INVX1_LOC_22/A 0.09fF
C25079 INPUT_0 INVX1_LOC_15/A 0.94fF
C25080 NOR2X1_LOC_111/A NOR2X1_LOC_841/A 0.10fF
C25081 INVX1_LOC_64/A INVX1_LOC_56/Y 0.00fF
C25082 NAND2X1_LOC_739/B NAND2X1_LOC_389/a_36_24# 0.00fF
C25083 INVX1_LOC_227/A NOR2X1_LOC_493/A 0.01fF
C25084 NOR2X1_LOC_401/a_36_216# INVX1_LOC_306/Y 0.00fF
C25085 NAND2X1_LOC_65/a_36_24# INVX1_LOC_120/A 0.00fF
C25086 INVX1_LOC_17/A NOR2X1_LOC_557/Y 0.00fF
C25087 VDD NOR2X1_LOC_673/A 0.08fF
C25088 INVX1_LOC_107/A INVX1_LOC_30/A 0.08fF
C25089 INVX1_LOC_35/A NOR2X1_LOC_209/a_36_216# 0.02fF
C25090 INVX1_LOC_225/A INVX1_LOC_14/A 0.13fF
C25091 NOR2X1_LOC_126/a_36_216# INVX1_LOC_76/A 0.00fF
C25092 INVX1_LOC_50/A INVX1_LOC_89/A 0.06fF
C25093 NOR2X1_LOC_637/B INVX1_LOC_246/A 0.05fF
C25094 INVX1_LOC_162/A INVX1_LOC_308/Y 0.10fF
C25095 INVX1_LOC_314/Y INVX1_LOC_31/A 0.10fF
C25096 NAND2X1_LOC_787/A NAND2X1_LOC_795/Y 0.01fF
C25097 INVX1_LOC_286/A INVX1_LOC_47/Y 0.19fF
C25098 NOR2X1_LOC_433/Y INVX1_LOC_54/A 0.11fF
C25099 NOR2X1_LOC_598/B INVX1_LOC_83/A 0.45fF
C25100 INVX1_LOC_11/A NOR2X1_LOC_309/Y -0.01fF
C25101 NOR2X1_LOC_92/Y NAND2X1_LOC_338/B 0.22fF
C25102 NOR2X1_LOC_857/A INVX1_LOC_19/A 0.15fF
C25103 INVX1_LOC_90/A INVX1_LOC_29/Y 0.03fF
C25104 NAND2X1_LOC_798/B INVX1_LOC_54/A 0.20fF
C25105 NOR2X1_LOC_169/B NOR2X1_LOC_303/Y 0.10fF
C25106 NOR2X1_LOC_724/Y INVX1_LOC_23/A 0.03fF
C25107 INVX1_LOC_72/A NAND2X1_LOC_837/Y 0.07fF
C25108 NOR2X1_LOC_91/A NOR2X1_LOC_597/Y 0.04fF
C25109 INVX1_LOC_130/A INVX1_LOC_33/A 0.01fF
C25110 D_INPUT_3 NAND2X1_LOC_82/Y 0.18fF
C25111 NOR2X1_LOC_541/Y INVX1_LOC_104/A 0.01fF
C25112 NOR2X1_LOC_389/B INVX1_LOC_29/Y 0.07fF
C25113 NAND2X1_LOC_508/A NOR2X1_LOC_105/Y 0.03fF
C25114 NOR2X1_LOC_590/A NOR2X1_LOC_388/Y 0.16fF
C25115 INVX1_LOC_28/A INVX1_LOC_57/A 7.77fF
C25116 NAND2X1_LOC_308/Y NAND2X1_LOC_727/a_36_24# 0.00fF
C25117 NOR2X1_LOC_65/B INVX1_LOC_73/A 0.07fF
C25118 INVX1_LOC_36/A NOR2X1_LOC_433/A 0.26fF
C25119 NAND2X1_LOC_35/Y NOR2X1_LOC_700/Y 0.16fF
C25120 INVX1_LOC_177/Y INVX1_LOC_71/A 0.07fF
C25121 INPUT_1 NOR2X1_LOC_717/A 0.16fF
C25122 INVX1_LOC_17/A INVX1_LOC_143/A 0.07fF
C25123 INVX1_LOC_280/A NOR2X1_LOC_814/A 0.03fF
C25124 INVX1_LOC_75/A NOR2X1_LOC_113/a_36_216# 0.12fF
C25125 NAND2X1_LOC_241/Y INVX1_LOC_42/A 0.01fF
C25126 NOR2X1_LOC_500/A NOR2X1_LOC_324/Y 0.04fF
C25127 NAND2X1_LOC_649/B INVX1_LOC_15/A 0.01fF
C25128 NOR2X1_LOC_625/a_36_216# NAND2X1_LOC_837/Y 0.01fF
C25129 INVX1_LOC_36/A NOR2X1_LOC_593/Y 0.03fF
C25130 NAND2X1_LOC_123/Y INVX1_LOC_23/A 0.03fF
C25131 NOR2X1_LOC_703/B NOR2X1_LOC_550/B 0.00fF
C25132 NOR2X1_LOC_516/B INVX1_LOC_1/A 0.14fF
C25133 NOR2X1_LOC_843/A NOR2X1_LOC_500/B 0.03fF
C25134 INVX1_LOC_41/A INVX1_LOC_72/A 0.10fF
C25135 NOR2X1_LOC_295/Y INVX1_LOC_30/A 1.29fF
C25136 NOR2X1_LOC_666/Y INVX1_LOC_16/A 0.24fF
C25137 NOR2X1_LOC_498/Y INVX1_LOC_72/A 0.07fF
C25138 NAND2X1_LOC_85/Y INVX1_LOC_46/Y 0.03fF
C25139 NOR2X1_LOC_791/B INVX1_LOC_33/A 0.03fF
C25140 NOR2X1_LOC_590/Y INVX1_LOC_89/A 0.05fF
C25141 NOR2X1_LOC_721/B INVX1_LOC_9/A 0.01fF
C25142 NOR2X1_LOC_2/Y INVX1_LOC_296/Y 0.05fF
C25143 NAND2X1_LOC_181/Y NOR2X1_LOC_786/a_36_216# 0.00fF
C25144 INVX1_LOC_120/A NOR2X1_LOC_849/A 0.60fF
C25145 INVX1_LOC_45/A INVX1_LOC_104/A 0.14fF
C25146 INVX1_LOC_145/A NOR2X1_LOC_433/A 0.05fF
C25147 INVX1_LOC_104/A NOR2X1_LOC_568/A 0.07fF
C25148 NOR2X1_LOC_208/Y NOR2X1_LOC_433/A 0.42fF
C25149 NOR2X1_LOC_13/Y INVX1_LOC_49/A 0.08fF
C25150 INVX1_LOC_36/A NOR2X1_LOC_52/B 0.30fF
C25151 INVX1_LOC_64/A NOR2X1_LOC_385/Y 0.04fF
C25152 NAND2X1_LOC_53/Y NAND2X1_LOC_831/a_36_24# 0.00fF
C25153 INVX1_LOC_41/A INVX1_LOC_198/Y 0.12fF
C25154 NOR2X1_LOC_357/Y INVX1_LOC_32/A 0.03fF
C25155 INVX1_LOC_2/A NOR2X1_LOC_658/Y 0.61fF
C25156 NOR2X1_LOC_208/Y NOR2X1_LOC_593/Y 0.12fF
C25157 NOR2X1_LOC_557/A NOR2X1_LOC_668/Y 0.03fF
C25158 INVX1_LOC_256/A INVX1_LOC_1/Y 0.25fF
C25159 NOR2X1_LOC_613/a_36_216# NAND2X1_LOC_866/B 0.03fF
C25160 INVX1_LOC_13/A NOR2X1_LOC_296/Y 0.10fF
C25161 INVX1_LOC_81/A INVX1_LOC_33/A 0.03fF
C25162 INVX1_LOC_43/Y INVX1_LOC_56/Y 0.00fF
C25163 NOR2X1_LOC_207/A INVX1_LOC_72/A 0.02fF
C25164 INVX1_LOC_278/A INPUT_0 0.79fF
C25165 NOR2X1_LOC_458/a_36_216# INVX1_LOC_206/Y 0.01fF
C25166 NAND2X1_LOC_778/Y NOR2X1_LOC_497/Y 0.01fF
C25167 NOR2X1_LOC_602/A INVX1_LOC_248/A 0.10fF
C25168 INVX1_LOC_78/A NAND2X1_LOC_241/Y 0.01fF
C25169 NOR2X1_LOC_78/A NOR2X1_LOC_383/B 0.11fF
C25170 INVX1_LOC_17/A NAND2X1_LOC_783/A 0.13fF
C25171 INVX1_LOC_37/A NOR2X1_LOC_855/A 0.01fF
C25172 NOR2X1_LOC_577/Y INVX1_LOC_155/Y 0.02fF
C25173 INVX1_LOC_13/A INPUT_3 1.63fF
C25174 NOR2X1_LOC_589/A NAND2X1_LOC_352/B 0.07fF
C25175 INVX1_LOC_25/A INVX1_LOC_315/Y 0.11fF
C25176 INVX1_LOC_145/A NOR2X1_LOC_52/B 0.02fF
C25177 NAND2X1_LOC_182/A INVX1_LOC_71/A 0.04fF
C25178 NOR2X1_LOC_264/Y NOR2X1_LOC_350/A 0.05fF
C25179 INVX1_LOC_104/A INVX1_LOC_71/A 0.27fF
C25180 INVX1_LOC_2/Y NAND2X1_LOC_223/A 0.03fF
C25181 NOR2X1_LOC_208/Y NOR2X1_LOC_52/B 0.02fF
C25182 INVX1_LOC_17/A NOR2X1_LOC_130/A 0.11fF
C25183 NAND2X1_LOC_656/A NOR2X1_LOC_709/A 0.18fF
C25184 INVX1_LOC_29/A INVX1_LOC_92/A 0.83fF
C25185 VDD NOR2X1_LOC_409/B 0.09fF
C25186 NOR2X1_LOC_658/Y NOR2X1_LOC_218/Y 0.04fF
C25187 NOR2X1_LOC_309/Y NOR2X1_LOC_433/A 0.03fF
C25188 NAND2X1_LOC_141/A D_INPUT_2 0.11fF
C25189 NOR2X1_LOC_456/Y INVX1_LOC_91/A 2.05fF
C25190 NOR2X1_LOC_280/Y NOR2X1_LOC_301/A 0.01fF
C25191 INVX1_LOC_163/A NOR2X1_LOC_19/B 0.00fF
C25192 NAND2X1_LOC_10/a_36_24# INVX1_LOC_123/A 0.01fF
C25193 INVX1_LOC_2/A NOR2X1_LOC_13/Y 0.10fF
C25194 NOR2X1_LOC_791/B INVX1_LOC_40/A 0.03fF
C25195 INVX1_LOC_96/A NOR2X1_LOC_678/A 0.72fF
C25196 NOR2X1_LOC_770/B INVX1_LOC_153/Y 0.13fF
C25197 INVX1_LOC_36/A NAND2X1_LOC_645/a_36_24# 0.00fF
C25198 INVX1_LOC_223/A NOR2X1_LOC_570/Y 0.32fF
C25199 NOR2X1_LOC_309/Y NOR2X1_LOC_593/Y 0.02fF
C25200 INVX1_LOC_26/Y NOR2X1_LOC_857/A 0.05fF
C25201 NOR2X1_LOC_657/B INVX1_LOC_23/A 0.55fF
C25202 NOR2X1_LOC_717/B NOR2X1_LOC_644/B 0.07fF
C25203 NAND2X1_LOC_53/Y D_GATE_366 0.03fF
C25204 NOR2X1_LOC_227/B INVX1_LOC_75/A 0.04fF
C25205 INVX1_LOC_93/A NOR2X1_LOC_167/Y 0.11fF
C25206 NOR2X1_LOC_590/A INVX1_LOC_135/A 0.05fF
C25207 NAND2X1_LOC_538/Y NOR2X1_LOC_329/B 0.07fF
C25208 INVX1_LOC_33/A NOR2X1_LOC_802/A 0.02fF
C25209 INVX1_LOC_57/A NOR2X1_LOC_35/Y 0.10fF
C25210 INVX1_LOC_84/A NOR2X1_LOC_84/B 0.02fF
C25211 NOR2X1_LOC_446/A NOR2X1_LOC_644/A 0.01fF
C25212 NOR2X1_LOC_536/A INVX1_LOC_87/A 0.02fF
C25213 NOR2X1_LOC_48/B NAND2X1_LOC_798/B 0.10fF
C25214 NOR2X1_LOC_68/A NAND2X1_LOC_662/Y 0.03fF
C25215 NOR2X1_LOC_445/Y INVX1_LOC_266/Y 0.09fF
C25216 NAND2X1_LOC_854/B NAND2X1_LOC_856/A 0.01fF
C25217 NOR2X1_LOC_613/a_36_216# INVX1_LOC_6/A 0.00fF
C25218 NOR2X1_LOC_250/A NOR2X1_LOC_329/B 0.08fF
C25219 INVX1_LOC_89/A INVX1_LOC_61/Y 0.03fF
C25220 INVX1_LOC_2/A NAND2X1_LOC_175/B 0.31fF
C25221 NOR2X1_LOC_689/Y INVX1_LOC_46/A 0.03fF
C25222 NOR2X1_LOC_309/Y NOR2X1_LOC_52/B 0.11fF
C25223 INVX1_LOC_17/A NOR2X1_LOC_216/Y 0.01fF
C25224 NOR2X1_LOC_252/Y INVX1_LOC_24/A 0.02fF
C25225 INVX1_LOC_41/A NOR2X1_LOC_537/Y 0.03fF
C25226 NOR2X1_LOC_590/A NOR2X1_LOC_560/A 0.02fF
C25227 NAND2X1_LOC_721/B NAND2X1_LOC_808/A 0.01fF
C25228 INVX1_LOC_41/A NAND2X1_LOC_338/B 0.12fF
C25229 NOR2X1_LOC_299/Y INVX1_LOC_72/A 0.19fF
C25230 NOR2X1_LOC_447/Y INVX1_LOC_22/A 0.01fF
C25231 INVX1_LOC_41/A NAND2X1_LOC_323/B 0.03fF
C25232 NAND2X1_LOC_659/a_36_24# INVX1_LOC_175/A 0.00fF
C25233 NOR2X1_LOC_89/A INVX1_LOC_63/A 0.01fF
C25234 NOR2X1_LOC_346/A NAND2X1_LOC_206/Y 0.03fF
C25235 NOR2X1_LOC_859/A INVX1_LOC_120/A 0.03fF
C25236 INVX1_LOC_178/A NAND2X1_LOC_623/B 0.01fF
C25237 NAND2X1_LOC_714/B INVX1_LOC_91/A 0.03fF
C25238 NOR2X1_LOC_831/B INVX1_LOC_4/A 0.14fF
C25239 NAND2X1_LOC_561/B INVX1_LOC_309/A 0.01fF
C25240 INVX1_LOC_207/A INVX1_LOC_241/A 0.02fF
C25241 NOR2X1_LOC_214/B NOR2X1_LOC_194/a_36_216# 0.00fF
C25242 NAND2X1_LOC_93/B INVX1_LOC_87/A 0.03fF
C25243 NAND2X1_LOC_470/B INVX1_LOC_117/Y 0.06fF
C25244 NOR2X1_LOC_82/A INVX1_LOC_126/Y 0.01fF
C25245 NOR2X1_LOC_644/B NOR2X1_LOC_151/Y 0.01fF
C25246 NOR2X1_LOC_561/A INVX1_LOC_29/Y 0.07fF
C25247 NAND2X1_LOC_338/B NOR2X1_LOC_398/Y 0.02fF
C25248 NAND2X1_LOC_725/A INVX1_LOC_46/A 0.08fF
C25249 NOR2X1_LOC_364/Y INVX1_LOC_22/A 0.05fF
C25250 NOR2X1_LOC_122/Y INVX1_LOC_72/A 0.03fF
C25251 NAND2X1_LOC_243/Y INVX1_LOC_23/Y 0.43fF
C25252 NOR2X1_LOC_160/B NOR2X1_LOC_188/A 0.10fF
C25253 NOR2X1_LOC_78/B NAND2X1_LOC_660/A 1.27fF
C25254 INVX1_LOC_273/Y NOR2X1_LOC_152/Y 0.03fF
C25255 NAND2X1_LOC_715/B INVX1_LOC_46/A 0.07fF
C25256 INVX1_LOC_298/Y INVX1_LOC_92/A 0.06fF
C25257 NOR2X1_LOC_602/a_36_216# NOR2X1_LOC_329/B 0.02fF
C25258 NOR2X1_LOC_160/B NOR2X1_LOC_548/B 0.10fF
C25259 NAND2X1_LOC_637/Y INVX1_LOC_296/A 0.01fF
C25260 NOR2X1_LOC_137/Y NOR2X1_LOC_674/a_36_216# 0.00fF
C25261 NAND2X1_LOC_81/B NOR2X1_LOC_76/B 0.01fF
C25262 NOR2X1_LOC_84/Y INVX1_LOC_316/Y 0.02fF
C25263 INVX1_LOC_207/A NOR2X1_LOC_298/Y 0.36fF
C25264 NOR2X1_LOC_789/B INVX1_LOC_20/A 0.01fF
C25265 NOR2X1_LOC_226/A INVX1_LOC_256/Y 0.01fF
C25266 NOR2X1_LOC_354/B NOR2X1_LOC_567/B 0.09fF
C25267 INVX1_LOC_227/A NOR2X1_LOC_388/Y 0.21fF
C25268 INVX1_LOC_14/A NAND2X1_LOC_642/Y 0.13fF
C25269 INVX1_LOC_13/A INVX1_LOC_158/A 0.04fF
C25270 NOR2X1_LOC_620/B INVX1_LOC_226/A 0.03fF
C25271 INVX1_LOC_256/A NOR2X1_LOC_318/B 0.12fF
C25272 NOR2X1_LOC_481/A NOR2X1_LOC_137/A 1.22fF
C25273 INVX1_LOC_226/Y NOR2X1_LOC_520/A 0.03fF
C25274 INVX1_LOC_77/A INVX1_LOC_85/Y 0.03fF
C25275 INVX1_LOC_5/A INVX1_LOC_117/A 0.29fF
C25276 NOR2X1_LOC_563/a_36_216# INVX1_LOC_177/A 0.00fF
C25277 NOR2X1_LOC_822/Y INVX1_LOC_22/A 0.02fF
C25278 INVX1_LOC_204/A INVX1_LOC_92/A 0.02fF
C25279 NOR2X1_LOC_211/A NOR2X1_LOC_537/Y 0.20fF
C25280 NAND2X1_LOC_367/A NAND2X1_LOC_367/B 0.19fF
C25281 NAND2X1_LOC_364/Y NAND2X1_LOC_366/a_36_24# 0.02fF
C25282 NAND2X1_LOC_833/Y NAND2X1_LOC_861/Y 0.20fF
C25283 INVX1_LOC_175/A NOR2X1_LOC_649/B 0.04fF
C25284 NOR2X1_LOC_532/Y INVX1_LOC_33/A 0.01fF
C25285 INVX1_LOC_290/A NAND2X1_LOC_661/B 0.03fF
C25286 INVX1_LOC_161/Y NOR2X1_LOC_405/A 0.01fF
C25287 NOR2X1_LOC_355/A NOR2X1_LOC_392/B 0.13fF
C25288 NAND2X1_LOC_779/a_36_24# NOR2X1_LOC_574/A 0.00fF
C25289 INVX1_LOC_31/A NOR2X1_LOC_557/A 0.17fF
C25290 NOR2X1_LOC_708/Y NOR2X1_LOC_708/B 0.38fF
C25291 NAND2X1_LOC_198/B NOR2X1_LOC_74/A 0.10fF
C25292 INVX1_LOC_289/A NAND2X1_LOC_752/a_36_24# 0.02fF
C25293 NAND2X1_LOC_722/A NAND2X1_LOC_795/Y 0.01fF
C25294 NOR2X1_LOC_32/B NOR2X1_LOC_88/A 0.02fF
C25295 NOR2X1_LOC_590/A NOR2X1_LOC_552/A 0.12fF
C25296 INVX1_LOC_53/A NOR2X1_LOC_634/A 0.01fF
C25297 INVX1_LOC_83/A NAND2X1_LOC_660/A 0.20fF
C25298 NOR2X1_LOC_300/Y NOR2X1_LOC_214/B 0.03fF
C25299 NOR2X1_LOC_229/Y INVX1_LOC_290/A 0.05fF
C25300 INVX1_LOC_161/Y NOR2X1_LOC_682/a_36_216# 0.00fF
C25301 NOR2X1_LOC_808/A D_INPUT_0 0.04fF
C25302 INVX1_LOC_35/A NAND2X1_LOC_647/a_36_24# 0.00fF
C25303 INVX1_LOC_312/A NOR2X1_LOC_405/A 0.02fF
C25304 INVX1_LOC_68/Y NOR2X1_LOC_199/B 0.03fF
C25305 NOR2X1_LOC_440/Y INVX1_LOC_1/Y 0.07fF
C25306 NOR2X1_LOC_178/Y NOR2X1_LOC_216/B 0.10fF
C25307 NAND2X1_LOC_195/Y NOR2X1_LOC_43/Y 0.02fF
C25308 INVX1_LOC_289/Y NOR2X1_LOC_536/A 0.00fF
C25309 INVX1_LOC_314/Y INVX1_LOC_6/A 0.06fF
C25310 INVX1_LOC_9/A NAND2X1_LOC_473/A 0.22fF
C25311 INVX1_LOC_245/Y INVX1_LOC_37/A 0.01fF
C25312 INVX1_LOC_36/A NOR2X1_LOC_601/Y 0.01fF
C25313 NAND2X1_LOC_454/Y INVX1_LOC_290/Y 0.03fF
C25314 INVX1_LOC_104/A INVX1_LOC_102/Y 0.00fF
C25315 NOR2X1_LOC_176/Y NAND2X1_LOC_793/Y 0.09fF
C25316 INVX1_LOC_256/Y INPUT_1 0.00fF
C25317 INVX1_LOC_45/A NOR2X1_LOC_840/a_36_216# 0.00fF
C25318 INVX1_LOC_236/Y NOR2X1_LOC_305/Y 0.01fF
C25319 INVX1_LOC_30/A NAND2X1_LOC_469/B 0.13fF
C25320 INVX1_LOC_14/A NOR2X1_LOC_271/Y 0.06fF
C25321 NOR2X1_LOC_756/Y INVX1_LOC_34/Y 0.07fF
C25322 NOR2X1_LOC_510/Y NOR2X1_LOC_58/a_36_216# 0.01fF
C25323 INVX1_LOC_314/Y NOR2X1_LOC_10/a_36_216# 0.00fF
C25324 NOR2X1_LOC_82/A NOR2X1_LOC_536/A 0.09fF
C25325 INVX1_LOC_300/Y INVX1_LOC_11/Y 0.01fF
C25326 NOR2X1_LOC_550/B INVX1_LOC_91/A 0.01fF
C25327 NOR2X1_LOC_383/Y NOR2X1_LOC_71/Y 0.15fF
C25328 INVX1_LOC_85/Y NOR2X1_LOC_687/Y 0.03fF
C25329 NAND2X1_LOC_564/B NAND2X1_LOC_551/A 0.00fF
C25330 NOR2X1_LOC_590/A NOR2X1_LOC_152/A 0.05fF
C25331 NOR2X1_LOC_91/A INVX1_LOC_170/Y 0.12fF
C25332 D_INPUT_1 NAND2X1_LOC_80/a_36_24# 0.01fF
C25333 NOR2X1_LOC_67/A NOR2X1_LOC_256/Y 0.04fF
C25334 NOR2X1_LOC_16/Y INPUT_0 0.01fF
C25335 INVX1_LOC_53/A INVX1_LOC_29/A 7.48fF
C25336 NAND2X1_LOC_63/Y NOR2X1_LOC_717/A 0.01fF
C25337 NOR2X1_LOC_763/Y INVX1_LOC_295/A 0.14fF
C25338 INVX1_LOC_302/A INVX1_LOC_22/A 0.02fF
C25339 NOR2X1_LOC_82/A NAND2X1_LOC_93/B 0.68fF
C25340 NOR2X1_LOC_303/Y INVX1_LOC_76/A 0.13fF
C25341 NAND2X1_LOC_363/B NAND2X1_LOC_200/a_36_24# 0.00fF
C25342 INVX1_LOC_17/A NOR2X1_LOC_197/B 0.91fF
C25343 NOR2X1_LOC_387/Y INVX1_LOC_20/A 0.03fF
C25344 INVX1_LOC_269/A NAND2X1_LOC_572/B 0.10fF
C25345 NOR2X1_LOC_294/Y INVX1_LOC_230/A 0.00fF
C25346 INVX1_LOC_208/A NOR2X1_LOC_188/A 0.01fF
C25347 INVX1_LOC_53/Y NOR2X1_LOC_74/A 0.07fF
C25348 NAND2X1_LOC_35/Y INVX1_LOC_284/A 0.10fF
C25349 NOR2X1_LOC_516/B NOR2X1_LOC_188/A 0.06fF
C25350 NAND2X1_LOC_350/A NAND2X1_LOC_798/B 2.81fF
C25351 NOR2X1_LOC_311/Y NAND2X1_LOC_660/A 0.10fF
C25352 NOR2X1_LOC_665/A NOR2X1_LOC_74/A 0.16fF
C25353 INVX1_LOC_53/Y NOR2X1_LOC_9/Y 0.09fF
C25354 NOR2X1_LOC_612/B NAND2X1_LOC_642/Y 0.02fF
C25355 NAND2X1_LOC_391/Y NAND2X1_LOC_74/B 0.16fF
C25356 NOR2X1_LOC_254/Y INVX1_LOC_76/A 0.01fF
C25357 NOR2X1_LOC_329/B NOR2X1_LOC_106/A 0.01fF
C25358 NOR2X1_LOC_635/a_36_216# NOR2X1_LOC_467/A 0.00fF
C25359 INVX1_LOC_275/A INVX1_LOC_14/Y 0.16fF
C25360 NAND2X1_LOC_363/B INVX1_LOC_251/A 0.01fF
C25361 INVX1_LOC_69/Y INVX1_LOC_1/Y 0.07fF
C25362 NAND2X1_LOC_222/B INVX1_LOC_63/A 0.00fF
C25363 NOR2X1_LOC_82/A NOR2X1_LOC_649/B 0.18fF
C25364 NAND2X1_LOC_36/A NAND2X1_LOC_93/B 0.01fF
C25365 NAND2X1_LOC_526/a_36_24# INVX1_LOC_91/A 0.01fF
C25366 NOR2X1_LOC_122/Y INVX1_LOC_313/Y 0.01fF
C25367 INVX1_LOC_224/A INVX1_LOC_63/A 0.03fF
C25368 NOR2X1_LOC_82/A INVX1_LOC_3/A 3.37fF
C25369 INVX1_LOC_23/Y NOR2X1_LOC_39/Y 0.05fF
C25370 NOR2X1_LOC_172/Y NOR2X1_LOC_111/A 0.16fF
C25371 NAND2X1_LOC_357/B INVX1_LOC_20/A 0.14fF
C25372 NAND2X1_LOC_721/B INVX1_LOC_92/A 0.03fF
C25373 NAND2X1_LOC_48/a_36_24# INVX1_LOC_9/A 0.00fF
C25374 INVX1_LOC_11/A INVX1_LOC_63/A 0.61fF
C25375 INVX1_LOC_5/A INVX1_LOC_3/Y 0.18fF
C25376 NAND2X1_LOC_36/A NAND2X1_LOC_425/Y 0.00fF
C25377 NAND2X1_LOC_369/a_36_24# NOR2X1_LOC_356/A 0.00fF
C25378 NAND2X1_LOC_381/Y INVX1_LOC_63/A 0.16fF
C25379 NAND2X1_LOC_366/A INVX1_LOC_117/A 0.10fF
C25380 NAND2X1_LOC_656/A NOR2X1_LOC_489/A 0.35fF
C25381 INVX1_LOC_23/Y NAND2X1_LOC_205/A 0.10fF
C25382 NAND2X1_LOC_464/B NAND2X1_LOC_99/A 0.07fF
C25383 INVX1_LOC_175/A NOR2X1_LOC_476/B 0.00fF
C25384 NOR2X1_LOC_353/Y INVX1_LOC_76/A 0.02fF
C25385 INVX1_LOC_297/Y INVX1_LOC_11/Y 0.02fF
C25386 INVX1_LOC_298/Y INVX1_LOC_53/A 0.49fF
C25387 INVX1_LOC_83/A INVX1_LOC_201/A 0.04fF
C25388 NAND2X1_LOC_549/B INVX1_LOC_20/A 0.01fF
C25389 NAND2X1_LOC_660/A INVX1_LOC_46/A 0.07fF
C25390 NOR2X1_LOC_377/Y INVX1_LOC_117/A 0.03fF
C25391 INVX1_LOC_178/A INVX1_LOC_3/Y 0.28fF
C25392 NOR2X1_LOC_860/B NOR2X1_LOC_61/Y 0.53fF
C25393 INVX1_LOC_160/Y INVX1_LOC_160/A 0.01fF
C25394 NOR2X1_LOC_748/Y NOR2X1_LOC_799/B 0.14fF
C25395 NOR2X1_LOC_440/Y INVX1_LOC_93/Y 0.10fF
C25396 NOR2X1_LOC_486/B INVX1_LOC_9/A 1.34fF
C25397 INVX1_LOC_271/A INVX1_LOC_23/A 0.17fF
C25398 INVX1_LOC_40/A INVX1_LOC_2/Y 0.03fF
C25399 INVX1_LOC_13/A NOR2X1_LOC_332/B 0.03fF
C25400 NOR2X1_LOC_596/A INVX1_LOC_113/A 0.35fF
C25401 NOR2X1_LOC_210/B VDD 0.01fF
C25402 NAND2X1_LOC_802/A NOR2X1_LOC_88/Y 0.01fF
C25403 NOR2X1_LOC_309/Y NOR2X1_LOC_675/a_36_216# 0.00fF
C25404 NOR2X1_LOC_644/A INVX1_LOC_186/A 0.03fF
C25405 NOR2X1_LOC_679/Y NOR2X1_LOC_48/B 0.07fF
C25406 NOR2X1_LOC_794/A NOR2X1_LOC_703/A 0.00fF
C25407 INVX1_LOC_218/A NAND2X1_LOC_96/A 0.07fF
C25408 INVX1_LOC_240/A INVX1_LOC_185/A 0.47fF
C25409 INVX1_LOC_49/A NAND2X1_LOC_85/Y 0.00fF
C25410 INVX1_LOC_299/A NAND2X1_LOC_615/a_36_24# 0.00fF
C25411 INVX1_LOC_8/A INVX1_LOC_92/A 0.05fF
C25412 NAND2X1_LOC_9/Y NOR2X1_LOC_598/B 0.05fF
C25413 NOR2X1_LOC_828/B NOR2X1_LOC_685/A 0.04fF
C25414 INVX1_LOC_246/A NAND2X1_LOC_419/a_36_24# 0.01fF
C25415 NAND2X1_LOC_9/Y INVX1_LOC_51/A 0.02fF
C25416 NAND2X1_LOC_319/A NAND2X1_LOC_453/A 0.02fF
C25417 NAND2X1_LOC_837/a_36_24# NAND2X1_LOC_859/B 0.00fF
C25418 INVX1_LOC_58/A NAND2X1_LOC_552/A 0.03fF
C25419 NOR2X1_LOC_186/Y NOR2X1_LOC_383/B 0.03fF
C25420 NAND2X1_LOC_802/A INVX1_LOC_84/A 0.00fF
C25421 NAND2X1_LOC_166/a_36_24# INVX1_LOC_29/A 0.01fF
C25422 INVX1_LOC_64/A NOR2X1_LOC_790/B 0.07fF
C25423 NOR2X1_LOC_91/A NOR2X1_LOC_824/A 0.07fF
C25424 NOR2X1_LOC_201/A INVX1_LOC_27/A -0.00fF
C25425 INVX1_LOC_58/A INVX1_LOC_5/A 0.22fF
C25426 NOR2X1_LOC_714/Y INVX1_LOC_307/Y 0.34fF
C25427 NOR2X1_LOC_246/A NOR2X1_LOC_279/Y 0.01fF
C25428 NOR2X1_LOC_234/Y NAND2X1_LOC_243/B 0.11fF
C25429 INVX1_LOC_7/Y INVX1_LOC_224/Y 0.01fF
C25430 INPUT_3 INVX1_LOC_32/A 1.02fF
C25431 NOR2X1_LOC_3/a_36_216# NOR2X1_LOC_11/Y 0.00fF
C25432 NOR2X1_LOC_552/A NOR2X1_LOC_703/A 0.01fF
C25433 NAND2X1_LOC_493/a_36_24# NOR2X1_LOC_536/A 0.00fF
C25434 INVX1_LOC_11/A NAND2X1_LOC_452/Y 0.03fF
C25435 INVX1_LOC_263/A NOR2X1_LOC_331/B -0.07fF
C25436 NOR2X1_LOC_433/A INVX1_LOC_63/A 0.14fF
C25437 NOR2X1_LOC_644/A NAND2X1_LOC_447/Y 0.17fF
C25438 INVX1_LOC_77/A NAND2X1_LOC_782/B 0.08fF
C25439 D_INPUT_0 INVX1_LOC_37/A 0.03fF
C25440 NOR2X1_LOC_160/Y INVX1_LOC_38/A 0.02fF
C25441 NOR2X1_LOC_151/Y NOR2X1_LOC_352/a_36_216# 0.00fF
C25442 NOR2X1_LOC_186/Y NAND2X1_LOC_777/a_36_24# 0.01fF
C25443 INVX1_LOC_49/A NAND2X1_LOC_249/a_36_24# 0.01fF
C25444 INVX1_LOC_196/A NOR2X1_LOC_809/B 0.07fF
C25445 NOR2X1_LOC_593/Y INVX1_LOC_63/A 0.00fF
C25446 NAND2X1_LOC_222/B NAND2X1_LOC_223/B 0.02fF
C25447 INVX1_LOC_58/A INVX1_LOC_178/A 0.03fF
C25448 INVX1_LOC_27/A INVX1_LOC_23/A 0.12fF
C25449 NOR2X1_LOC_689/A NAND2X1_LOC_724/A 0.17fF
C25450 NOR2X1_LOC_598/B NOR2X1_LOC_798/A 0.03fF
C25451 NOR2X1_LOC_412/a_36_216# NOR2X1_LOC_662/A 0.01fF
C25452 INVX1_LOC_20/Y VDD 0.21fF
C25453 INVX1_LOC_224/Y NOR2X1_LOC_92/Y 0.09fF
C25454 INVX1_LOC_48/Y INVX1_LOC_57/A 0.07fF
C25455 NOR2X1_LOC_447/Y INVX1_LOC_261/A 0.40fF
C25456 NOR2X1_LOC_328/Y INVX1_LOC_54/A 0.04fF
C25457 INVX1_LOC_90/A NOR2X1_LOC_111/A 0.10fF
C25458 INVX1_LOC_69/Y NOR2X1_LOC_318/B 0.29fF
C25459 INVX1_LOC_2/A NOR2X1_LOC_697/Y 0.03fF
C25460 NOR2X1_LOC_382/Y NOR2X1_LOC_38/B 0.11fF
C25461 NAND2X1_LOC_777/a_36_24# NAND2X1_LOC_573/Y 0.00fF
C25462 NOR2X1_LOC_732/A NAND2X1_LOC_782/B 0.05fF
C25463 NOR2X1_LOC_52/B INVX1_LOC_63/A 0.06fF
C25464 INVX1_LOC_266/Y INVX1_LOC_84/A 0.07fF
C25465 NAND2X1_LOC_849/A INVX1_LOC_20/A 0.01fF
C25466 NOR2X1_LOC_226/A NOR2X1_LOC_697/Y 0.07fF
C25467 NAND2X1_LOC_36/A NAND2X1_LOC_470/B 0.01fF
C25468 NAND2X1_LOC_560/A INVX1_LOC_46/A 0.03fF
C25469 NOR2X1_LOC_590/A NOR2X1_LOC_541/B 0.01fF
C25470 NOR2X1_LOC_810/A NOR2X1_LOC_856/A 0.02fF
C25471 NAND2X1_LOC_35/Y NOR2X1_LOC_384/A 0.01fF
C25472 NOR2X1_LOC_657/B INVX1_LOC_6/A 0.03fF
C25473 NOR2X1_LOC_741/a_36_216# INVX1_LOC_139/Y 0.00fF
C25474 INVX1_LOC_35/A NOR2X1_LOC_140/A 0.15fF
C25475 NOR2X1_LOC_15/Y NOR2X1_LOC_678/A 0.03fF
C25476 NOR2X1_LOC_591/Y INVX1_LOC_49/Y 0.08fF
C25477 INVX1_LOC_269/A INVX1_LOC_58/Y 0.02fF
C25478 NOR2X1_LOC_318/B NOR2X1_LOC_543/a_36_216# 0.00fF
C25479 NOR2X1_LOC_139/Y NOR2X1_LOC_269/Y 0.07fF
C25480 NOR2X1_LOC_664/Y NOR2X1_LOC_664/a_36_216# 0.03fF
C25481 INVX1_LOC_246/A INVX1_LOC_57/A 0.07fF
C25482 D_INPUT_0 NOR2X1_LOC_177/Y 0.03fF
C25483 INVX1_LOC_159/A NOR2X1_LOC_158/B 0.02fF
C25484 INVX1_LOC_50/A NOR2X1_LOC_599/Y 0.42fF
C25485 INVX1_LOC_58/A NOR2X1_LOC_816/A 0.05fF
C25486 INVX1_LOC_55/Y NOR2X1_LOC_261/A 0.01fF
C25487 INVX1_LOC_306/A NAND2X1_LOC_93/B 0.00fF
C25488 NOR2X1_LOC_234/Y INVX1_LOC_284/A 0.02fF
C25489 NAND2X1_LOC_634/a_36_24# NOR2X1_LOC_291/Y 0.01fF
C25490 INVX1_LOC_24/A INVX1_LOC_94/Y 0.07fF
C25491 INVX1_LOC_31/A INVX1_LOC_271/A 0.01fF
C25492 NAND2X1_LOC_468/B NOR2X1_LOC_269/Y 0.01fF
C25493 NAND2X1_LOC_451/Y NAND2X1_LOC_639/a_36_24# 0.00fF
C25494 NAND2X1_LOC_59/B D_INPUT_5 0.16fF
C25495 INVX1_LOC_83/A NOR2X1_LOC_58/Y 0.32fF
C25496 D_INPUT_1 NAND2X1_LOC_208/B 0.03fF
C25497 NOR2X1_LOC_78/B INVX1_LOC_29/A 0.14fF
C25498 NAND2X1_LOC_11/Y INPUT_7 0.18fF
C25499 NOR2X1_LOC_687/Y NAND2X1_LOC_782/B 0.01fF
C25500 INVX1_LOC_77/A NAND2X1_LOC_454/Y 0.07fF
C25501 INVX1_LOC_177/Y NOR2X1_LOC_106/a_36_216# 0.00fF
C25502 NOR2X1_LOC_236/a_36_216# INVX1_LOC_3/A 0.02fF
C25503 INVX1_LOC_17/A INVX1_LOC_38/Y 0.02fF
C25504 NAND2X1_LOC_562/B INVX1_LOC_3/Y 0.17fF
C25505 NAND2X1_LOC_367/B NOR2X1_LOC_865/Y 0.29fF
C25506 INVX1_LOC_306/A INVX1_LOC_3/A 0.02fF
C25507 INVX1_LOC_248/Y NOR2X1_LOC_816/A 0.03fF
C25508 NAND2X1_LOC_862/a_36_24# INVX1_LOC_84/A 0.00fF
C25509 NAND2X1_LOC_721/B INVX1_LOC_53/A 0.12fF
C25510 INVX1_LOC_266/Y INVX1_LOC_15/A 0.04fF
C25511 INVX1_LOC_24/A INVX1_LOC_296/A 0.07fF
C25512 INVX1_LOC_254/Y INVX1_LOC_26/Y 0.02fF
C25513 INVX1_LOC_58/A NOR2X1_LOC_273/a_36_216# 0.00fF
C25514 INVX1_LOC_247/Y INVX1_LOC_53/A 0.01fF
C25515 INVX1_LOC_137/Y NAND2X1_LOC_74/B 0.01fF
C25516 INVX1_LOC_206/Y NOR2X1_LOC_331/B 0.07fF
C25517 NAND2X1_LOC_214/B INVX1_LOC_31/A 0.14fF
C25518 INVX1_LOC_1/Y NOR2X1_LOC_89/A 0.02fF
C25519 NOR2X1_LOC_298/Y NOR2X1_LOC_36/B 0.12fF
C25520 NOR2X1_LOC_32/B INVX1_LOC_18/A 0.17fF
C25521 NOR2X1_LOC_433/A NOR2X1_LOC_65/Y 0.01fF
C25522 NOR2X1_LOC_655/B INVX1_LOC_47/Y 0.10fF
C25523 NAND2X1_LOC_392/Y INVX1_LOC_29/A 0.00fF
C25524 NAND2X1_LOC_506/a_36_24# NOR2X1_LOC_243/B 0.00fF
C25525 NOR2X1_LOC_92/Y NOR2X1_LOC_103/Y 0.00fF
C25526 INVX1_LOC_305/A NOR2X1_LOC_434/A 0.04fF
C25527 NAND2X1_LOC_593/Y NOR2X1_LOC_677/Y 0.04fF
C25528 NOR2X1_LOC_328/Y NOR2X1_LOC_48/B 0.05fF
C25529 NAND2X1_LOC_35/Y INVX1_LOC_72/A 0.07fF
C25530 NOR2X1_LOC_350/A INVX1_LOC_57/A 0.02fF
C25531 NOR2X1_LOC_374/A NOR2X1_LOC_383/B 0.03fF
C25532 NAND2X1_LOC_123/Y NOR2X1_LOC_117/Y 0.00fF
C25533 INVX1_LOC_95/Y INVX1_LOC_129/Y 0.02fF
C25534 INVX1_LOC_185/Y NOR2X1_LOC_301/A 0.02fF
C25535 INVX1_LOC_27/A INVX1_LOC_31/A 0.08fF
C25536 NOR2X1_LOC_481/A NOR2X1_LOC_383/B 0.07fF
C25537 NOR2X1_LOC_824/A INVX1_LOC_31/A 0.07fF
C25538 INVX1_LOC_83/A INVX1_LOC_29/A 0.07fF
C25539 NOR2X1_LOC_6/a_36_216# INVX1_LOC_57/A 0.00fF
C25540 NAND2X1_LOC_32/a_36_24# NAND2X1_LOC_555/Y 0.00fF
C25541 NOR2X1_LOC_128/B NOR2X1_LOC_128/A 0.02fF
C25542 NOR2X1_LOC_542/Y INVX1_LOC_19/A 0.56fF
C25543 NOR2X1_LOC_751/A NAND2X1_LOC_750/a_36_24# 0.02fF
C25544 INVX1_LOC_201/Y NOR2X1_LOC_400/B 0.05fF
C25545 INVX1_LOC_9/Y INVX1_LOC_32/A 0.26fF
C25546 NOR2X1_LOC_600/Y NOR2X1_LOC_331/B 0.01fF
C25547 NOR2X1_LOC_454/Y NOR2X1_LOC_478/A 0.01fF
C25548 NOR2X1_LOC_470/B NOR2X1_LOC_471/Y 0.08fF
C25549 NOR2X1_LOC_496/Y INVX1_LOC_30/A 0.01fF
C25550 INVX1_LOC_33/A INVX1_LOC_29/Y 0.03fF
C25551 INVX1_LOC_225/A NOR2X1_LOC_383/B 0.07fF
C25552 NOR2X1_LOC_32/B INVX1_LOC_172/A 0.02fF
C25553 NOR2X1_LOC_681/Y NOR2X1_LOC_682/Y 0.05fF
C25554 NOR2X1_LOC_849/a_36_216# INVX1_LOC_27/A 0.02fF
C25555 NOR2X1_LOC_536/A INVX1_LOC_59/Y 0.02fF
C25556 NOR2X1_LOC_737/a_36_216# INVX1_LOC_179/A 0.00fF
C25557 NOR2X1_LOC_288/A NOR2X1_LOC_383/B 0.03fF
C25558 INVX1_LOC_136/A NAND2X1_LOC_391/Y 0.01fF
C25559 INVX1_LOC_13/Y NOR2X1_LOC_360/Y 0.07fF
C25560 INVX1_LOC_311/Y INVX1_LOC_19/A 0.13fF
C25561 D_INPUT_1 INVX1_LOC_34/A 0.22fF
C25562 INVX1_LOC_1/Y INVX1_LOC_104/Y 0.01fF
C25563 INVX1_LOC_45/A NOR2X1_LOC_92/Y 0.10fF
C25564 INVX1_LOC_298/Y NOR2X1_LOC_78/B 0.03fF
C25565 INVX1_LOC_75/Y INVX1_LOC_91/A 0.01fF
C25566 D_GATE_366 INVX1_LOC_12/A 0.10fF
C25567 NAND2X1_LOC_595/a_36_24# NAND2X1_LOC_555/Y 0.00fF
C25568 INVX1_LOC_201/Y NAND2X1_LOC_38/a_36_24# 0.01fF
C25569 INVX1_LOC_58/A NAND2X1_LOC_562/B 0.01fF
C25570 INVX1_LOC_45/A INVX1_LOC_24/Y 2.14fF
C25571 NOR2X1_LOC_802/A NOR2X1_LOC_748/A 0.12fF
C25572 NOR2X1_LOC_560/A NOR2X1_LOC_67/Y 0.06fF
C25573 INVX1_LOC_215/Y NOR2X1_LOC_816/A 0.01fF
C25574 INVX1_LOC_104/A NOR2X1_LOC_493/A 0.06fF
C25575 NOR2X1_LOC_84/Y INVX1_LOC_57/A 0.07fF
C25576 NOR2X1_LOC_332/A INVX1_LOC_3/Y 0.07fF
C25577 INVX1_LOC_224/Y NOR2X1_LOC_398/Y 0.00fF
C25578 NOR2X1_LOC_454/Y NOR2X1_LOC_68/A 0.17fF
C25579 INVX1_LOC_17/A INVX1_LOC_286/Y 1.41fF
C25580 INVX1_LOC_64/A NOR2X1_LOC_344/A 0.16fF
C25581 INVX1_LOC_59/Y NOR2X1_LOC_655/Y 0.00fF
C25582 NAND2X1_LOC_200/B NOR2X1_LOC_668/Y 0.11fF
C25583 NOR2X1_LOC_689/A NAND2X1_LOC_852/Y 0.05fF
C25584 NAND2X1_LOC_463/B INVX1_LOC_163/Y 0.01fF
C25585 INVX1_LOC_206/A INVX1_LOC_23/A 0.02fF
C25586 NAND2X1_LOC_231/Y NAND2X1_LOC_231/a_36_24# 0.02fF
C25587 NOR2X1_LOC_145/Y INVX1_LOC_193/A 0.21fF
C25588 NOR2X1_LOC_289/Y INVX1_LOC_12/A 0.00fF
C25589 NOR2X1_LOC_692/Y NAND2X1_LOC_804/Y 0.00fF
C25590 NOR2X1_LOC_111/A INVX1_LOC_38/A 0.03fF
C25591 INVX1_LOC_232/A INVX1_LOC_16/Y 0.59fF
C25592 NOR2X1_LOC_440/Y INVX1_LOC_87/A 0.07fF
C25593 NAND2X1_LOC_570/Y INVX1_LOC_23/A 0.01fF
C25594 NOR2X1_LOC_742/A NOR2X1_LOC_89/A 0.07fF
C25595 NOR2X1_LOC_45/B INVX1_LOC_285/A 0.07fF
C25596 INVX1_LOC_14/A NOR2X1_LOC_91/Y 0.24fF
C25597 INVX1_LOC_64/A NAND2X1_LOC_357/B 0.07fF
C25598 NAND2X1_LOC_783/A INVX1_LOC_94/Y 0.03fF
C25599 INVX1_LOC_88/A NOR2X1_LOC_360/Y 0.01fF
C25600 INVX1_LOC_277/A NOR2X1_LOC_160/B 0.07fF
C25601 NOR2X1_LOC_92/Y INVX1_LOC_71/A 0.10fF
C25602 NOR2X1_LOC_456/Y NOR2X1_LOC_352/Y 0.01fF
C25603 INVX1_LOC_35/A NOR2X1_LOC_709/A 0.01fF
C25604 INVX1_LOC_33/Y NOR2X1_LOC_602/B 0.01fF
C25605 INVX1_LOC_34/A NOR2X1_LOC_652/Y 0.07fF
C25606 INVX1_LOC_299/A INVX1_LOC_24/A 0.27fF
C25607 INVX1_LOC_58/A NOR2X1_LOC_773/Y 0.31fF
C25608 NOR2X1_LOC_130/A INVX1_LOC_94/Y 0.03fF
C25609 NAND2X1_LOC_738/B NAND2X1_LOC_852/Y 0.03fF
C25610 NOR2X1_LOC_76/A NOR2X1_LOC_89/a_36_216# 0.01fF
C25611 NOR2X1_LOC_188/A NAND2X1_LOC_207/B 0.03fF
C25612 INVX1_LOC_14/A NOR2X1_LOC_81/a_36_216# 0.01fF
C25613 INVX1_LOC_17/Y INVX1_LOC_22/A 0.18fF
C25614 INVX1_LOC_211/Y NAND2X1_LOC_354/Y 0.14fF
C25615 INVX1_LOC_135/A NOR2X1_LOC_415/Y 0.09fF
C25616 INVX1_LOC_256/A NAND2X1_LOC_514/Y 0.03fF
C25617 INVX1_LOC_50/A NAND2X1_LOC_349/B 0.01fF
C25618 NOR2X1_LOC_538/B INVX1_LOC_24/A 0.02fF
C25619 INVX1_LOC_232/A NAND2X1_LOC_205/A 0.39fF
C25620 INVX1_LOC_33/Y INVX1_LOC_54/A 0.03fF
C25621 NOR2X1_LOC_15/Y NAND2X1_LOC_738/a_36_24# 0.00fF
C25622 INVX1_LOC_290/A INVX1_LOC_57/A 0.03fF
C25623 INVX1_LOC_90/A INVX1_LOC_90/Y 0.02fF
C25624 INVX1_LOC_64/A NAND2X1_LOC_549/B 0.01fF
C25625 NOR2X1_LOC_91/A INVX1_LOC_234/A 0.00fF
C25626 NOR2X1_LOC_373/Y INVX1_LOC_23/Y 0.00fF
C25627 INVX1_LOC_174/A NOR2X1_LOC_546/A 0.42fF
C25628 INVX1_LOC_225/Y NOR2X1_LOC_168/Y 0.02fF
C25629 NAND2X1_LOC_35/Y NAND2X1_LOC_338/B 0.01fF
C25630 NOR2X1_LOC_58/Y INVX1_LOC_46/A 0.17fF
C25631 NAND2X1_LOC_391/Y NOR2X1_LOC_278/A 0.04fF
C25632 INVX1_LOC_59/Y INVX1_LOC_3/A 0.03fF
C25633 NOR2X1_LOC_299/Y NAND2X1_LOC_402/B 0.00fF
C25634 NOR2X1_LOC_264/a_36_216# NOR2X1_LOC_716/B 0.00fF
C25635 NOR2X1_LOC_51/A NOR2X1_LOC_694/Y 0.43fF
C25636 INVX1_LOC_269/A NOR2X1_LOC_716/B 0.10fF
C25637 INVX1_LOC_293/A INVX1_LOC_24/A 0.00fF
C25638 NOR2X1_LOC_383/Y NAND2X1_LOC_205/A 0.25fF
C25639 INVX1_LOC_42/Y INVX1_LOC_15/A 0.01fF
C25640 NAND2X1_LOC_848/A NOR2X1_LOC_177/Y 0.27fF
C25641 NOR2X1_LOC_329/B NOR2X1_LOC_334/Y 0.02fF
C25642 INVX1_LOC_91/A NAND2X1_LOC_74/B 0.24fF
C25643 NOR2X1_LOC_130/A INVX1_LOC_181/A 0.07fF
C25644 NAND2X1_LOC_231/Y NOR2X1_LOC_652/Y 0.10fF
C25645 D_INPUT_0 NAND2X1_LOC_96/a_36_24# 0.00fF
C25646 INVX1_LOC_74/A INVX1_LOC_63/A 0.05fF
C25647 NOR2X1_LOC_264/Y INVX1_LOC_1/A 0.02fF
C25648 INVX1_LOC_234/A INVX1_LOC_23/A 0.21fF
C25649 NAND2X1_LOC_568/A NAND2X1_LOC_568/a_36_24# 0.00fF
C25650 NOR2X1_LOC_318/B NOR2X1_LOC_89/A 0.09fF
C25651 NOR2X1_LOC_824/A NOR2X1_LOC_290/Y 0.22fF
C25652 INVX1_LOC_254/A NAND2X1_LOC_114/B 0.09fF
C25653 INVX1_LOC_21/A INVX1_LOC_210/A 0.12fF
C25654 VDD NOR2X1_LOC_450/B -0.00fF
C25655 INVX1_LOC_64/A NOR2X1_LOC_540/a_36_216# 0.00fF
C25656 NOR2X1_LOC_216/Y INVX1_LOC_94/Y 0.03fF
C25657 INVX1_LOC_41/A NOR2X1_LOC_103/Y 0.12fF
C25658 NOR2X1_LOC_403/B NAND2X1_LOC_208/B 0.05fF
C25659 NAND2X1_LOC_551/A NAND2X1_LOC_97/a_36_24# 0.00fF
C25660 INVX1_LOC_93/Y NOR2X1_LOC_89/A 0.02fF
C25661 NOR2X1_LOC_461/A INVX1_LOC_9/A 0.03fF
C25662 VDD NOR2X1_LOC_257/Y 0.24fF
C25663 NOR2X1_LOC_478/A INVX1_LOC_77/A 0.00fF
C25664 NAND2X1_LOC_51/B NOR2X1_LOC_158/Y 0.05fF
C25665 NOR2X1_LOC_446/A NOR2X1_LOC_570/B 0.24fF
C25666 INVX1_LOC_16/A INVX1_LOC_306/Y 0.08fF
C25667 NAND2X1_LOC_140/A INVX1_LOC_53/A 0.01fF
C25668 NOR2X1_LOC_160/B NOR2X1_LOC_285/B 0.06fF
C25669 NAND2X1_LOC_53/Y INVX1_LOC_85/A 0.01fF
C25670 NOR2X1_LOC_589/Y INVX1_LOC_78/A 0.01fF
C25671 NOR2X1_LOC_552/A NOR2X1_LOC_169/a_36_216# 0.01fF
C25672 INVX1_LOC_36/A INVX1_LOC_314/Y 0.07fF
C25673 NOR2X1_LOC_103/Y NAND2X1_LOC_477/A 0.09fF
C25674 NOR2X1_LOC_15/Y NOR2X1_LOC_191/A 0.01fF
C25675 NAND2X1_LOC_23/a_36_24# INVX1_LOC_75/A 0.00fF
C25676 INVX1_LOC_46/A INVX1_LOC_29/A 0.30fF
C25677 INVX1_LOC_21/A INVX1_LOC_13/A 0.08fF
C25678 INVX1_LOC_118/A NOR2X1_LOC_697/Y 0.05fF
C25679 NOR2X1_LOC_538/B INVX1_LOC_143/A 0.01fF
C25680 NOR2X1_LOC_197/Y NOR2X1_LOC_748/A 0.15fF
C25681 NOR2X1_LOC_19/B INVX1_LOC_23/A 0.77fF
C25682 NOR2X1_LOC_664/Y INVX1_LOC_31/A 0.95fF
C25683 NOR2X1_LOC_160/B NOR2X1_LOC_87/B 0.00fF
C25684 INVX1_LOC_41/A INVX1_LOC_45/A 4.72fF
C25685 INVX1_LOC_50/A INVX1_LOC_75/A 0.09fF
C25686 NOR2X1_LOC_824/A NAND2X1_LOC_859/Y 0.10fF
C25687 INVX1_LOC_58/A INVX1_LOC_140/A 0.19fF
C25688 INVX1_LOC_110/Y NOR2X1_LOC_844/A 0.04fF
C25689 NOR2X1_LOC_68/A INVX1_LOC_77/A 3.49fF
C25690 NAND2X1_LOC_149/Y NAND2X1_LOC_149/B 0.11fF
C25691 INVX1_LOC_1/A INVX1_LOC_316/Y 0.00fF
C25692 INVX1_LOC_30/A INVX1_LOC_63/Y 0.78fF
C25693 NAND2X1_LOC_493/Y INVX1_LOC_22/A 0.00fF
C25694 INVX1_LOC_303/A NOR2X1_LOC_360/Y 0.07fF
C25695 NOR2X1_LOC_795/Y NOR2X1_LOC_590/A 0.00fF
C25696 NAND2X1_LOC_721/A NOR2X1_LOC_89/A 0.07fF
C25697 INVX1_LOC_64/A NOR2X1_LOC_702/Y 0.01fF
C25698 NOR2X1_LOC_160/B NAND2X1_LOC_360/B 0.09fF
C25699 NAND2X1_LOC_569/A NOR2X1_LOC_384/Y 0.15fF
C25700 NOR2X1_LOC_296/a_36_216# INVX1_LOC_226/Y 0.00fF
C25701 INVX1_LOC_7/A NAND2X1_LOC_473/A 0.07fF
C25702 NAND2X1_LOC_623/B INVX1_LOC_78/A 0.01fF
C25703 INVX1_LOC_45/A NAND2X1_LOC_477/A 0.01fF
C25704 INVX1_LOC_224/A INVX1_LOC_1/Y 0.00fF
C25705 INVX1_LOC_21/A NOR2X1_LOC_246/A 0.14fF
C25706 NAND2X1_LOC_724/Y NOR2X1_LOC_387/A 0.03fF
C25707 NOR2X1_LOC_250/Y INVX1_LOC_53/Y 0.23fF
C25708 D_INPUT_1 INPUT_0 0.17fF
C25709 NAND2X1_LOC_364/A NOR2X1_LOC_392/B 0.08fF
C25710 INVX1_LOC_27/A INVX1_LOC_313/A 0.03fF
C25711 NOR2X1_LOC_68/A NOR2X1_LOC_732/A 0.02fF
C25712 INVX1_LOC_11/A INVX1_LOC_1/Y 4.81fF
C25713 NOR2X1_LOC_545/A INVX1_LOC_77/A 0.09fF
C25714 INVX1_LOC_30/A NOR2X1_LOC_175/A 0.05fF
C25715 INVX1_LOC_117/A INVX1_LOC_42/A 0.11fF
C25716 NOR2X1_LOC_637/a_36_216# NOR2X1_LOC_637/Y 0.00fF
C25717 NOR2X1_LOC_91/A NOR2X1_LOC_528/Y 0.01fF
C25718 INVX1_LOC_6/A INVX1_LOC_271/A 0.05fF
C25719 NAND2X1_LOC_770/Y INVX1_LOC_297/A 0.07fF
C25720 NOR2X1_LOC_272/Y INVX1_LOC_90/A 0.05fF
C25721 NOR2X1_LOC_583/Y INVX1_LOC_38/A 0.01fF
C25722 INVX1_LOC_33/Y NOR2X1_LOC_48/B 0.07fF
C25723 NAND2X1_LOC_200/B INVX1_LOC_31/A 0.01fF
C25724 NOR2X1_LOC_862/B NOR2X1_LOC_814/A 0.10fF
C25725 NAND2X1_LOC_72/Y INVX1_LOC_75/A 0.12fF
C25726 NOR2X1_LOC_824/A NAND2X1_LOC_866/B 0.14fF
C25727 INVX1_LOC_41/A INVX1_LOC_71/A 0.07fF
C25728 NOR2X1_LOC_272/Y NOR2X1_LOC_389/B 0.10fF
C25729 NAND2X1_LOC_348/A INVX1_LOC_138/Y 0.01fF
C25730 INVX1_LOC_288/Y INVX1_LOC_91/A 0.01fF
C25731 INVX1_LOC_34/A D_INPUT_2 0.05fF
C25732 INVX1_LOC_269/A NOR2X1_LOC_326/Y 0.31fF
C25733 NAND2X1_LOC_348/A NOR2X1_LOC_860/a_36_216# 0.00fF
C25734 INVX1_LOC_45/A NOR2X1_LOC_405/a_36_216# 0.00fF
C25735 NAND2X1_LOC_521/a_36_24# NOR2X1_LOC_844/A 0.00fF
C25736 INVX1_LOC_61/Y INVX1_LOC_25/Y 0.08fF
C25737 NOR2X1_LOC_328/a_36_216# NOR2X1_LOC_25/Y 0.00fF
C25738 NAND2X1_LOC_78/a_36_24# NOR2X1_LOC_188/A 0.01fF
C25739 NOR2X1_LOC_810/A INVX1_LOC_134/A 0.02fF
C25740 INVX1_LOC_24/A NOR2X1_LOC_315/Y 0.01fF
C25741 NOR2X1_LOC_314/Y INVX1_LOC_78/A 0.01fF
C25742 INVX1_LOC_247/Y NOR2X1_LOC_78/B 0.01fF
C25743 NOR2X1_LOC_815/Y NAND2X1_LOC_175/B 0.04fF
C25744 NOR2X1_LOC_383/B NAND2X1_LOC_642/Y 0.16fF
C25745 NAND2X1_LOC_477/A INVX1_LOC_71/A 0.10fF
C25746 VDD NOR2X1_LOC_30/Y 0.24fF
C25747 INVX1_LOC_223/A NOR2X1_LOC_500/Y 0.01fF
C25748 NOR2X1_LOC_690/A NAND2X1_LOC_483/Y 0.07fF
C25749 NOR2X1_LOC_432/Y INVX1_LOC_24/A 0.01fF
C25750 INPUT_0 NOR2X1_LOC_652/Y 0.37fF
C25751 NOR2X1_LOC_609/a_36_216# INVX1_LOC_177/A 0.00fF
C25752 INVX1_LOC_298/Y INVX1_LOC_46/A 0.02fF
C25753 VDD NOR2X1_LOC_301/A 0.21fF
C25754 NOR2X1_LOC_281/Y INVX1_LOC_46/A 0.00fF
C25755 NOR2X1_LOC_274/Y INVX1_LOC_54/Y 0.02fF
C25756 INVX1_LOC_17/A NAND2X1_LOC_186/a_36_24# 0.00fF
C25757 NOR2X1_LOC_92/Y INVX1_LOC_102/Y 0.07fF
C25758 INVX1_LOC_234/A INVX1_LOC_31/A 0.46fF
C25759 NOR2X1_LOC_75/Y NOR2X1_LOC_214/B 0.00fF
C25760 INVX1_LOC_78/A INVX1_LOC_117/A 0.16fF
C25761 VDD NOR2X1_LOC_302/A -0.00fF
C25762 NOR2X1_LOC_388/Y INVX1_LOC_104/A 1.30fF
C25763 INVX1_LOC_12/A INVX1_LOC_123/Y 0.00fF
C25764 INVX1_LOC_84/A INVX1_LOC_19/A 0.59fF
C25765 INVX1_LOC_24/A INVX1_LOC_52/A 0.03fF
C25766 NOR2X1_LOC_68/A NOR2X1_LOC_687/Y 0.13fF
C25767 NAND2X1_LOC_149/Y NOR2X1_LOC_74/A 0.08fF
C25768 NOR2X1_LOC_808/A INVX1_LOC_49/A 1.52fF
C25769 NOR2X1_LOC_179/Y NAND2X1_LOC_74/B 0.01fF
C25770 NOR2X1_LOC_433/A NOR2X1_LOC_362/a_36_216# 0.01fF
C25771 INVX1_LOC_27/A INVX1_LOC_6/A 0.26fF
C25772 INVX1_LOC_139/Y NOR2X1_LOC_632/a_36_216# 0.00fF
C25773 INVX1_LOC_223/A INVX1_LOC_10/A 0.10fF
C25774 NAND2X1_LOC_757/a_36_24# INVX1_LOC_25/Y -0.00fF
C25775 INVX1_LOC_34/A NOR2X1_LOC_529/Y 0.03fF
C25776 INVX1_LOC_50/A NAND2X1_LOC_453/A 0.03fF
C25777 INVX1_LOC_270/Y NOR2X1_LOC_137/Y 0.01fF
C25778 NOR2X1_LOC_215/Y NAND2X1_LOC_479/Y 0.01fF
C25779 INVX1_LOC_116/A INVX1_LOC_22/A 0.02fF
C25780 NOR2X1_LOC_764/Y NAND2X1_LOC_36/A 0.01fF
C25781 INVX1_LOC_37/A NOR2X1_LOC_451/a_36_216# 0.00fF
C25782 NOR2X1_LOC_65/B INVX1_LOC_117/A 0.10fF
C25783 NAND2X1_LOC_860/A INVX1_LOC_76/A 0.09fF
C25784 INVX1_LOC_11/A NOR2X1_LOC_742/A 0.11fF
C25785 INVX1_LOC_103/A NOR2X1_LOC_313/a_36_216# 0.00fF
C25786 INVX1_LOC_27/A NOR2X1_LOC_10/a_36_216# 0.12fF
C25787 NOR2X1_LOC_495/Y INVX1_LOC_22/A 0.00fF
C25788 NAND2X1_LOC_549/Y INVX1_LOC_20/A 0.01fF
C25789 NOR2X1_LOC_289/a_36_216# NOR2X1_LOC_172/Y 0.00fF
C25790 NOR2X1_LOC_78/B INVX1_LOC_8/A 0.17fF
C25791 INVX1_LOC_17/A NOR2X1_LOC_721/Y 0.00fF
C25792 INVX1_LOC_107/Y D_INPUT_5 0.16fF
C25793 NAND2X1_LOC_338/B NAND2X1_LOC_465/Y 0.39fF
C25794 INVX1_LOC_31/A NOR2X1_LOC_19/B 0.16fF
C25795 INVX1_LOC_14/Y NOR2X1_LOC_717/A 0.08fF
C25796 NOR2X1_LOC_315/Y INVX1_LOC_143/A 0.08fF
C25797 NOR2X1_LOC_791/B INVX1_LOC_89/A 0.03fF
C25798 D_INPUT_0 NAND2X1_LOC_198/B 0.10fF
C25799 NOR2X1_LOC_593/Y INVX1_LOC_1/Y 0.01fF
C25800 NOR2X1_LOC_383/B NOR2X1_LOC_271/Y 0.02fF
C25801 INVX1_LOC_269/A NOR2X1_LOC_392/a_36_216# 0.12fF
C25802 NOR2X1_LOC_307/B NOR2X1_LOC_731/A 0.24fF
C25803 NOR2X1_LOC_430/A INPUT_5 0.04fF
C25804 NOR2X1_LOC_553/B NOR2X1_LOC_550/B 0.17fF
C25805 INVX1_LOC_90/A NAND2X1_LOC_364/A 0.09fF
C25806 INVX1_LOC_75/A INVX1_LOC_61/Y 0.07fF
C25807 INVX1_LOC_214/A INVX1_LOC_236/A 0.02fF
C25808 INVX1_LOC_310/A INVX1_LOC_143/A 0.00fF
C25809 NOR2X1_LOC_671/Y INVX1_LOC_29/A 0.03fF
C25810 INVX1_LOC_60/Y INVX1_LOC_40/A 0.92fF
C25811 INVX1_LOC_294/Y INVX1_LOC_16/A 0.04fF
C25812 INVX1_LOC_255/Y NAND2X1_LOC_139/A 0.02fF
C25813 NOR2X1_LOC_389/B NAND2X1_LOC_364/A 0.08fF
C25814 NOR2X1_LOC_653/Y INVX1_LOC_15/A 0.05fF
C25815 INVX1_LOC_163/Y INVX1_LOC_42/A 0.49fF
C25816 NOR2X1_LOC_419/a_36_216# NOR2X1_LOC_99/B 0.00fF
C25817 INVX1_LOC_90/A NAND2X1_LOC_100/a_36_24# 0.00fF
C25818 INVX1_LOC_54/A NOR2X1_LOC_686/a_36_216# 0.01fF
C25819 NOR2X1_LOC_567/B NOR2X1_LOC_500/B 0.11fF
C25820 INVX1_LOC_88/A NOR2X1_LOC_269/Y 0.10fF
C25821 INVX1_LOC_223/A NAND2X1_LOC_132/a_36_24# 0.00fF
C25822 NOR2X1_LOC_52/B INVX1_LOC_1/Y 0.07fF
C25823 NOR2X1_LOC_516/B NOR2X1_LOC_87/B 1.26fF
C25824 NAND2X1_LOC_332/a_36_24# NAND2X1_LOC_211/Y 0.01fF
C25825 INVX1_LOC_102/A INVX1_LOC_12/A 0.07fF
C25826 NOR2X1_LOC_75/Y NOR2X1_LOC_741/A 0.01fF
C25827 NAND2X1_LOC_660/a_36_24# NOR2X1_LOC_577/Y 0.00fF
C25828 INVX1_LOC_102/A NOR2X1_LOC_519/Y 0.05fF
C25829 NOR2X1_LOC_121/A NOR2X1_LOC_709/A 0.02fF
C25830 INVX1_LOC_181/Y NOR2X1_LOC_153/a_36_216# 0.00fF
C25831 NOR2X1_LOC_355/A INVX1_LOC_33/A 0.01fF
C25832 INVX1_LOC_19/A INVX1_LOC_15/A 0.30fF
C25833 NOR2X1_LOC_557/Y INVX1_LOC_66/A -0.03fF
C25834 INVX1_LOC_161/Y INVX1_LOC_264/Y 0.01fF
C25835 NAND2X1_LOC_803/B NOR2X1_LOC_45/B 0.03fF
C25836 INVX1_LOC_289/A NOR2X1_LOC_226/A 0.03fF
C25837 INVX1_LOC_77/A NOR2X1_LOC_163/A 0.01fF
C25838 INVX1_LOC_41/A NOR2X1_LOC_123/B 0.25fF
C25839 NAND2X1_LOC_347/B INVX1_LOC_20/A 0.13fF
C25840 INVX1_LOC_11/A INVX1_LOC_93/Y 0.07fF
C25841 NOR2X1_LOC_770/Y INVX1_LOC_49/A 0.05fF
C25842 INVX1_LOC_45/A NAND2X1_LOC_309/a_36_24# 0.00fF
C25843 NAND2X1_LOC_182/a_36_24# INVX1_LOC_256/Y 0.00fF
C25844 NOR2X1_LOC_202/Y NOR2X1_LOC_215/Y 0.17fF
C25845 INVX1_LOC_72/A NOR2X1_LOC_83/Y 0.02fF
C25846 INVX1_LOC_17/A NOR2X1_LOC_56/Y 0.08fF
C25847 INVX1_LOC_31/A NOR2X1_LOC_528/Y 2.03fF
C25848 INVX1_LOC_135/A INVX1_LOC_104/A 1.24fF
C25849 NOR2X1_LOC_590/A NOR2X1_LOC_45/B 0.03fF
C25850 NOR2X1_LOC_679/Y INVX1_LOC_291/Y 0.02fF
C25851 INVX1_LOC_111/Y NOR2X1_LOC_543/A 0.28fF
C25852 NAND2X1_LOC_866/A NAND2X1_LOC_560/A 0.03fF
C25853 NAND2X1_LOC_537/Y INVX1_LOC_76/A 0.20fF
C25854 INVX1_LOC_89/A NOR2X1_LOC_124/B 0.01fF
C25855 INVX1_LOC_159/A NOR2X1_LOC_594/Y 0.01fF
C25856 NOR2X1_LOC_315/Y NOR2X1_LOC_130/A 0.03fF
C25857 NOR2X1_LOC_216/B INVX1_LOC_23/A 0.07fF
C25858 INVX1_LOC_136/A INVX1_LOC_309/A 0.03fF
C25859 INVX1_LOC_3/Y INVX1_LOC_42/A 1.30fF
C25860 NOR2X1_LOC_292/Y INVX1_LOC_181/Y 0.07fF
C25861 NOR2X1_LOC_641/B NOR2X1_LOC_78/A 0.00fF
C25862 NOR2X1_LOC_647/B INVX1_LOC_59/Y 0.00fF
C25863 INVX1_LOC_17/A INVX1_LOC_146/Y 0.03fF
C25864 INVX1_LOC_89/A NOR2X1_LOC_802/A 0.06fF
C25865 INPUT_0 D_INPUT_2 0.03fF
C25866 NOR2X1_LOC_464/B NAND2X1_LOC_472/Y 0.03fF
C25867 INVX1_LOC_17/A VDD 1.37fF
C25868 NOR2X1_LOC_590/A INVX1_LOC_247/A 0.03fF
C25869 INVX1_LOC_166/A INVX1_LOC_84/A 0.01fF
C25870 NOR2X1_LOC_742/A NOR2X1_LOC_593/Y 0.02fF
C25871 INVX1_LOC_41/A INVX1_LOC_102/Y 0.06fF
C25872 NAND2X1_LOC_785/A INVX1_LOC_90/A 0.14fF
C25873 NAND2X1_LOC_99/A NAND2X1_LOC_773/B 0.74fF
C25874 NAND2X1_LOC_555/Y NAND2X1_LOC_659/B 0.50fF
C25875 INVX1_LOC_136/A INVX1_LOC_91/A 0.63fF
C25876 NAND2X1_LOC_227/Y NAND2X1_LOC_453/A 0.01fF
C25877 NOR2X1_LOC_2/Y NOR2X1_LOC_11/a_36_216# 0.00fF
C25878 NAND2X1_LOC_30/Y INVX1_LOC_37/A 0.05fF
C25879 NOR2X1_LOC_89/A INVX1_LOC_87/A 0.02fF
C25880 NOR2X1_LOC_473/B INVX1_LOC_133/Y 0.00fF
C25881 NOR2X1_LOC_322/Y NAND2X1_LOC_325/Y 0.00fF
C25882 NOR2X1_LOC_667/A NOR2X1_LOC_246/A 0.01fF
C25883 INVX1_LOC_249/A INVX1_LOC_6/A 0.13fF
C25884 INVX1_LOC_85/A NOR2X1_LOC_302/Y 0.00fF
C25885 NOR2X1_LOC_589/Y INVX1_LOC_113/Y 0.21fF
C25886 NAND2X1_LOC_213/A INVX1_LOC_38/A 0.03fF
C25887 NOR2X1_LOC_92/Y NOR2X1_LOC_331/B 0.03fF
C25888 INVX1_LOC_248/A NOR2X1_LOC_246/A 0.01fF
C25889 NOR2X1_LOC_471/Y VDD 1.25fF
C25890 INVX1_LOC_36/A NOR2X1_LOC_657/B 0.24fF
C25891 NOR2X1_LOC_658/Y NAND2X1_LOC_212/Y 0.01fF
C25892 NOR2X1_LOC_569/Y INVX1_LOC_220/Y 0.13fF
C25893 INVX1_LOC_136/A INVX1_LOC_11/Y 0.06fF
C25894 INVX1_LOC_21/A NOR2X1_LOC_451/A 0.42fF
C25895 NAND2X1_LOC_363/B INVX1_LOC_27/Y 0.41fF
C25896 NAND2X1_LOC_662/Y INVX1_LOC_10/A 0.04fF
C25897 INVX1_LOC_13/Y NOR2X1_LOC_79/Y 0.20fF
C25898 NAND2X1_LOC_555/Y VDD 0.00fF
C25899 D_INPUT_0 INVX1_LOC_53/Y 0.96fF
C25900 NOR2X1_LOC_251/Y INVX1_LOC_313/A 0.02fF
C25901 NOR2X1_LOC_619/A D_INPUT_0 0.02fF
C25902 INVX1_LOC_33/A NOR2X1_LOC_552/Y 0.01fF
C25903 NOR2X1_LOC_798/A NOR2X1_LOC_634/A 0.02fF
C25904 INVX1_LOC_234/A NAND2X1_LOC_859/Y 0.65fF
C25905 NOR2X1_LOC_264/Y NOR2X1_LOC_188/A 0.01fF
C25906 NOR2X1_LOC_413/Y NAND2X1_LOC_622/B 0.02fF
C25907 D_INPUT_1 NOR2X1_LOC_84/B 0.18fF
C25908 INVX1_LOC_84/A NAND2X1_LOC_790/a_36_24# 0.00fF
C25909 NOR2X1_LOC_264/Y NOR2X1_LOC_548/B 0.12fF
C25910 NOR2X1_LOC_471/Y NOR2X1_LOC_684/a_36_216# 0.00fF
C25911 INVX1_LOC_53/Y NOR2X1_LOC_389/a_36_216# 0.00fF
C25912 NOR2X1_LOC_433/A NOR2X1_LOC_318/B 0.01fF
C25913 INVX1_LOC_57/A INVX1_LOC_261/Y 0.03fF
C25914 INVX1_LOC_182/Y NOR2X1_LOC_757/a_36_216# 0.00fF
C25915 NOR2X1_LOC_388/Y INVX1_LOC_206/Y 0.00fF
C25916 NOR2X1_LOC_242/A NOR2X1_LOC_240/A 0.04fF
C25917 INVX1_LOC_278/A INVX1_LOC_19/A 0.08fF
C25918 NOR2X1_LOC_208/Y NOR2X1_LOC_657/B 0.00fF
C25919 NOR2X1_LOC_441/Y INVX1_LOC_33/Y 1.63fF
C25920 INVX1_LOC_30/Y INVX1_LOC_47/A 0.00fF
C25921 NOR2X1_LOC_593/Y NOR2X1_LOC_318/B 0.24fF
C25922 INVX1_LOC_104/Y INVX1_LOC_87/A 0.01fF
C25923 INVX1_LOC_90/A NOR2X1_LOC_86/A 0.13fF
C25924 NAND2X1_LOC_634/Y INVX1_LOC_46/A 0.03fF
C25925 NAND2X1_LOC_9/Y INVX1_LOC_29/A 0.03fF
C25926 NOR2X1_LOC_433/A INVX1_LOC_93/Y 0.02fF
C25927 NAND2X1_LOC_654/B INVX1_LOC_22/A 0.00fF
C25928 INVX1_LOC_50/A INVX1_LOC_283/A 0.03fF
C25929 NOR2X1_LOC_609/a_36_216# NOR2X1_LOC_137/B 0.00fF
C25930 NOR2X1_LOC_794/A INVX1_LOC_104/A 0.02fF
C25931 INVX1_LOC_26/Y INVX1_LOC_15/A 0.03fF
C25932 INVX1_LOC_58/A INVX1_LOC_42/A 8.07fF
C25933 INVX1_LOC_103/A NAND2X1_LOC_93/B 0.08fF
C25934 INVX1_LOC_136/A NOR2X1_LOC_653/a_36_216# 0.01fF
C25935 INVX1_LOC_233/A INVX1_LOC_29/A 0.07fF
C25936 INVX1_LOC_299/A NOR2X1_LOC_197/B 0.10fF
C25937 NAND2X1_LOC_198/B NOR2X1_LOC_266/B 0.02fF
C25938 NOR2X1_LOC_593/Y INVX1_LOC_93/Y 0.00fF
C25939 NOR2X1_LOC_620/B INPUT_0 0.00fF
C25940 NOR2X1_LOC_393/Y NAND2X1_LOC_99/A 0.03fF
C25941 NAND2X1_LOC_725/B INVX1_LOC_260/Y 0.03fF
C25942 NOR2X1_LOC_769/A INVX1_LOC_117/A 0.01fF
C25943 INVX1_LOC_243/Y NOR2X1_LOC_467/A 0.17fF
C25944 NAND2X1_LOC_72/B NAND2X1_LOC_71/a_36_24# 0.02fF
C25945 INVX1_LOC_49/A NOR2X1_LOC_631/B 0.04fF
C25946 INVX1_LOC_11/A INVX1_LOC_117/Y 0.03fF
C25947 INVX1_LOC_21/A NAND2X1_LOC_489/Y 0.07fF
C25948 INVX1_LOC_315/Y NOR2X1_LOC_87/B 0.07fF
C25949 INVX1_LOC_103/A NAND2X1_LOC_425/Y 0.01fF
C25950 NOR2X1_LOC_318/B NOR2X1_LOC_52/B 0.83fF
C25951 NOR2X1_LOC_392/B NOR2X1_LOC_405/A 0.05fF
C25952 NOR2X1_LOC_552/A INVX1_LOC_104/A 0.07fF
C25953 INVX1_LOC_174/Y NOR2X1_LOC_706/A 0.00fF
C25954 INVX1_LOC_217/A NOR2X1_LOC_692/a_36_216# 0.00fF
C25955 INVX1_LOC_16/A NOR2X1_LOC_74/A 0.10fF
C25956 NOR2X1_LOC_433/A INVX1_LOC_139/A 0.03fF
C25957 INVX1_LOC_292/A NAND2X1_LOC_93/B 0.03fF
C25958 INPUT_6 NAND2X1_LOC_430/B 0.01fF
C25959 INVX1_LOC_161/Y NOR2X1_LOC_88/Y 0.03fF
C25960 NOR2X1_LOC_52/B INVX1_LOC_93/Y 0.07fF
C25961 NAND2X1_LOC_364/A INVX1_LOC_38/A 0.07fF
C25962 INVX1_LOC_186/Y NOR2X1_LOC_698/a_36_216# 0.00fF
C25963 NOR2X1_LOC_798/A INVX1_LOC_29/A 0.03fF
C25964 NOR2X1_LOC_6/B INVX1_LOC_95/Y 0.00fF
C25965 INVX1_LOC_24/A NAND2X1_LOC_96/A 0.08fF
C25966 NAND2X1_LOC_741/B INVX1_LOC_54/A 0.12fF
C25967 INVX1_LOC_49/A INVX1_LOC_37/A 1.30fF
C25968 NAND2X1_LOC_45/Y NOR2X1_LOC_112/Y 0.14fF
C25969 INVX1_LOC_16/A NOR2X1_LOC_9/Y 0.07fF
C25970 NOR2X1_LOC_590/A NOR2X1_LOC_862/B 0.06fF
C25971 NOR2X1_LOC_68/A INVX1_LOC_9/A 3.74fF
C25972 NOR2X1_LOC_152/Y INVX1_LOC_117/A 0.03fF
C25973 INVX1_LOC_286/A INVX1_LOC_232/A 0.12fF
C25974 NAND2X1_LOC_849/a_36_24# INVX1_LOC_309/A 0.00fF
C25975 INVX1_LOC_6/A INVX1_LOC_137/A 0.00fF
C25976 INVX1_LOC_31/A NOR2X1_LOC_216/B 0.08fF
C25977 NAND2X1_LOC_748/a_36_24# NAND2X1_LOC_74/B 0.01fF
C25978 NOR2X1_LOC_160/B NAND2X1_LOC_572/B 0.44fF
C25979 INVX1_LOC_58/A INVX1_LOC_78/A 0.15fF
C25980 INVX1_LOC_33/A NOR2X1_LOC_111/A 0.09fF
C25981 NOR2X1_LOC_716/B INVX1_LOC_12/Y 0.40fF
C25982 INVX1_LOC_8/A INVX1_LOC_46/A 0.02fF
C25983 INVX1_LOC_161/Y INVX1_LOC_84/A 0.03fF
C25984 INVX1_LOC_82/Y INVX1_LOC_89/A 0.01fF
C25985 NOR2X1_LOC_488/Y NOR2X1_LOC_45/B 0.00fF
C25986 INVX1_LOC_8/A NOR2X1_LOC_98/A 0.01fF
C25987 INVX1_LOC_217/A NOR2X1_LOC_517/a_36_216# 0.00fF
C25988 INVX1_LOC_14/A NAND2X1_LOC_82/Y 0.02fF
C25989 NOR2X1_LOC_52/B INVX1_LOC_139/A 0.34fF
C25990 NAND2X1_LOC_787/B NOR2X1_LOC_692/a_36_216# 0.01fF
C25991 NOR2X1_LOC_52/Y NOR2X1_LOC_364/A 0.31fF
C25992 NOR2X1_LOC_798/Y NOR2X1_LOC_809/A 0.00fF
C25993 INVX1_LOC_35/A NOR2X1_LOC_334/Y 0.07fF
C25994 INVX1_LOC_72/A NOR2X1_LOC_155/A 0.11fF
C25995 INVX1_LOC_223/A NOR2X1_LOC_445/B 0.01fF
C25996 INVX1_LOC_17/A INVX1_LOC_133/A 0.07fF
C25997 NAND2X1_LOC_156/B INVX1_LOC_6/A 0.45fF
C25998 NAND2X1_LOC_859/Y NOR2X1_LOC_528/Y 0.24fF
C25999 INVX1_LOC_289/Y NOR2X1_LOC_89/A 0.05fF
C26000 NOR2X1_LOC_52/B NAND2X1_LOC_721/A 0.07fF
C26001 INVX1_LOC_21/A INVX1_LOC_32/A 0.06fF
C26002 NAND2X1_LOC_205/A INVX1_LOC_112/Y 0.02fF
C26003 INVX1_LOC_2/A INVX1_LOC_37/A 0.15fF
C26004 INVX1_LOC_271/A INVX1_LOC_270/A 0.10fF
C26005 INVX1_LOC_198/Y NOR2X1_LOC_155/A 0.12fF
C26006 INVX1_LOC_28/A NOR2X1_LOC_74/A 0.03fF
C26007 INVX1_LOC_11/A NOR2X1_LOC_669/A 0.01fF
C26008 INVX1_LOC_240/A NOR2X1_LOC_536/A 0.06fF
C26009 INVX1_LOC_55/Y INVX1_LOC_311/A 0.98fF
C26010 NOR2X1_LOC_226/A NOR2X1_LOC_681/Y 0.04fF
C26011 INVX1_LOC_33/A INVX1_LOC_127/A 0.07fF
C26012 NOR2X1_LOC_82/A NOR2X1_LOC_89/A 3.79fF
C26013 NOR2X1_LOC_226/A INVX1_LOC_37/A 0.15fF
C26014 INVX1_LOC_25/A INVX1_LOC_57/A 0.09fF
C26015 NAND2X1_LOC_837/Y NOR2X1_LOC_491/Y 0.12fF
C26016 INVX1_LOC_30/Y INVX1_LOC_95/Y 0.03fF
C26017 INVX1_LOC_50/Y INVX1_LOC_271/Y 0.02fF
C26018 INVX1_LOC_200/A INVX1_LOC_102/A 0.02fF
C26019 NOR2X1_LOC_772/B INVX1_LOC_26/A 0.01fF
C26020 INVX1_LOC_282/A NAND2X1_LOC_849/A 0.02fF
C26021 NOR2X1_LOC_78/A NOR2X1_LOC_71/Y 0.02fF
C26022 NOR2X1_LOC_636/B NOR2X1_LOC_48/B 0.01fF
C26023 NAND2X1_LOC_477/A NOR2X1_LOC_331/B 0.07fF
C26024 NOR2X1_LOC_122/A INVX1_LOC_15/A 0.01fF
C26025 NAND2X1_LOC_347/B INVX1_LOC_4/A 0.03fF
C26026 INVX1_LOC_136/A INVX1_LOC_203/A 0.10fF
C26027 NAND2X1_LOC_785/A INVX1_LOC_38/A 0.38fF
C26028 INVX1_LOC_53/Y NOR2X1_LOC_266/B 0.03fF
C26029 NOR2X1_LOC_384/Y NOR2X1_LOC_662/A 0.07fF
C26030 NOR2X1_LOC_307/B INVX1_LOC_117/A 0.14fF
C26031 INVX1_LOC_21/A NAND2X1_LOC_175/Y 0.08fF
C26032 INVX1_LOC_13/Y INVX1_LOC_26/A 0.11fF
C26033 NOR2X1_LOC_252/Y VDD 0.12fF
C26034 NOR2X1_LOC_644/A NOR2X1_LOC_78/A 0.04fF
C26035 NOR2X1_LOC_533/A NOR2X1_LOC_536/A 0.27fF
C26036 NOR2X1_LOC_667/A NOR2X1_LOC_692/Y 0.01fF
C26037 NOR2X1_LOC_186/Y NAND2X1_LOC_288/B 0.27fF
C26038 NOR2X1_LOC_91/A INVX1_LOC_93/A -0.02fF
C26039 NAND2X1_LOC_807/Y NOR2X1_LOC_528/Y -0.00fF
C26040 INVX1_LOC_90/A NOR2X1_LOC_405/A 0.04fF
C26041 INVX1_LOC_161/Y INVX1_LOC_15/A 0.07fF
C26042 INVX1_LOC_223/A INVX1_LOC_12/A 0.03fF
C26043 NOR2X1_LOC_78/B INVX1_LOC_118/Y 0.07fF
C26044 NOR2X1_LOC_758/Y NOR2X1_LOC_831/B 0.01fF
C26045 NOR2X1_LOC_389/B NOR2X1_LOC_405/A 0.11fF
C26046 INVX1_LOC_279/A NOR2X1_LOC_858/B 0.03fF
C26047 NOR2X1_LOC_199/B VDD 0.00fF
C26048 INVX1_LOC_314/Y INVX1_LOC_63/A 2.20fF
C26049 INVX1_LOC_149/Y NOR2X1_LOC_445/B 0.01fF
C26050 NOR2X1_LOC_71/Y NAND2X1_LOC_464/A 0.07fF
C26051 INVX1_LOC_64/A NAND2X1_LOC_549/Y 0.00fF
C26052 NAND2X1_LOC_214/B NOR2X1_LOC_416/A 0.08fF
C26053 INVX1_LOC_103/A NAND2X1_LOC_470/B 0.09fF
C26054 INVX1_LOC_21/A INVX1_LOC_262/A 0.01fF
C26055 INVX1_LOC_2/A NOR2X1_LOC_743/Y 0.02fF
C26056 NAND2X1_LOC_787/A NAND2X1_LOC_552/A 0.04fF
C26057 INVX1_LOC_224/A INVX1_LOC_87/A 0.00fF
C26058 NAND2X1_LOC_477/A NOR2X1_LOC_592/B 0.06fF
C26059 NOR2X1_LOC_226/A NOR2X1_LOC_177/Y 0.02fF
C26060 NAND2X1_LOC_849/B NOR2X1_LOC_86/A 0.01fF
C26061 INVX1_LOC_89/A INVX1_LOC_2/Y 0.03fF
C26062 NAND2X1_LOC_514/Y NOR2X1_LOC_89/A 0.06fF
C26063 INVX1_LOC_217/A INVX1_LOC_102/A 0.04fF
C26064 INVX1_LOC_36/A INVX1_LOC_170/Y 0.00fF
C26065 INVX1_LOC_85/Y INVX1_LOC_76/A 0.03fF
C26066 NAND2X1_LOC_363/B INVX1_LOC_5/A 0.07fF
C26067 NOR2X1_LOC_209/Y INVX1_LOC_179/A 0.10fF
C26068 INVX1_LOC_265/A INVX1_LOC_265/Y 0.30fF
C26069 NAND2X1_LOC_55/a_36_24# INVX1_LOC_3/A 0.00fF
C26070 NOR2X1_LOC_356/A NOR2X1_LOC_35/Y 0.10fF
C26071 NOR2X1_LOC_751/A NOR2X1_LOC_78/A 0.01fF
C26072 NOR2X1_LOC_570/Y INVX1_LOC_9/A 0.12fF
C26073 INVX1_LOC_215/Y INVX1_LOC_78/A 0.34fF
C26074 INVX1_LOC_198/Y NOR2X1_LOC_833/B 0.05fF
C26075 NOR2X1_LOC_68/A NOR2X1_LOC_861/Y 0.15fF
C26076 INPUT_1 INVX1_LOC_37/A 0.03fF
C26077 NAND2X1_LOC_787/A INVX1_LOC_178/A 0.01fF
C26078 NOR2X1_LOC_528/Y INVX1_LOC_6/A 0.22fF
C26079 NAND2X1_LOC_21/Y INVX1_LOC_19/A 0.06fF
C26080 INVX1_LOC_1/A INVX1_LOC_57/A 0.15fF
C26081 NOR2X1_LOC_554/B INVX1_LOC_3/Y 0.07fF
C26082 NAND2X1_LOC_361/Y NOR2X1_LOC_777/B 2.27fF
C26083 NAND2X1_LOC_855/Y INVX1_LOC_76/A 0.04fF
C26084 INVX1_LOC_136/A INVX1_LOC_231/A 0.04fF
C26085 INVX1_LOC_286/Y INVX1_LOC_94/Y 0.02fF
C26086 NAND2X1_LOC_652/Y NAND2X1_LOC_453/A 0.02fF
C26087 INVX1_LOC_120/A NOR2X1_LOC_536/A 0.10fF
C26088 INVX1_LOC_5/A NOR2X1_LOC_840/A 0.02fF
C26089 NOR2X1_LOC_171/Y VDD 0.12fF
C26090 NAND2X1_LOC_276/Y NAND2X1_LOC_74/B 7.55fF
C26091 NAND2X1_LOC_354/Y NOR2X1_LOC_329/Y 0.10fF
C26092 NAND2X1_LOC_316/a_36_24# NOR2X1_LOC_89/A 0.01fF
C26093 NOR2X1_LOC_74/A NOR2X1_LOC_35/Y 0.01fF
C26094 INVX1_LOC_76/Y INVX1_LOC_19/A 0.01fF
C26095 NOR2X1_LOC_140/a_36_216# INVX1_LOC_29/A 0.00fF
C26096 INVX1_LOC_286/A NAND2X1_LOC_447/Y 0.10fF
C26097 NOR2X1_LOC_778/B INVX1_LOC_63/A 0.03fF
C26098 NOR2X1_LOC_16/Y INVX1_LOC_19/A 0.05fF
C26099 NOR2X1_LOC_9/Y NOR2X1_LOC_35/Y 0.05fF
C26100 NAND2X1_LOC_364/A NAND2X1_LOC_223/A 0.01fF
C26101 NOR2X1_LOC_594/Y VDD 0.01fF
C26102 NAND2X1_LOC_354/Y NAND2X1_LOC_175/Y 0.04fF
C26103 NOR2X1_LOC_122/Y NOR2X1_LOC_331/B 0.02fF
C26104 NOR2X1_LOC_87/B NAND2X1_LOC_207/B 0.02fF
C26105 INVX1_LOC_48/Y INVX1_LOC_306/Y 0.82fF
C26106 NOR2X1_LOC_34/B NAND2X1_LOC_473/A 0.02fF
C26107 NOR2X1_LOC_316/Y INVX1_LOC_12/A -0.03fF
C26108 NOR2X1_LOC_299/Y NOR2X1_LOC_491/Y 0.02fF
C26109 NOR2X1_LOC_112/B NAND2X1_LOC_96/A 0.13fF
C26110 NAND2X1_LOC_35/Y NOR2X1_LOC_103/Y 0.03fF
C26111 INVX1_LOC_163/A INVX1_LOC_242/A 0.19fF
C26112 NOR2X1_LOC_516/B NAND2X1_LOC_219/B 0.23fF
C26113 INVX1_LOC_50/A NOR2X1_LOC_274/B 0.94fF
C26114 D_GATE_366 INVX1_LOC_92/A 0.03fF
C26115 INVX1_LOC_36/A INVX1_LOC_271/A 0.13fF
C26116 NOR2X1_LOC_689/Y INVX1_LOC_72/A 0.04fF
C26117 NOR2X1_LOC_45/B NAND2X1_LOC_650/B 0.07fF
C26118 INVX1_LOC_22/A INVX1_LOC_240/Y 0.00fF
C26119 NOR2X1_LOC_384/Y INVX1_LOC_57/A 0.03fF
C26120 INVX1_LOC_17/A NOR2X1_LOC_510/Y 0.03fF
C26121 INVX1_LOC_24/A NAND2X1_LOC_99/A 0.16fF
C26122 NOR2X1_LOC_11/a_36_216# NOR2X1_LOC_36/A 0.02fF
C26123 INVX1_LOC_200/Y INVX1_LOC_18/A 0.03fF
C26124 NAND2X1_LOC_714/B NAND2X1_LOC_538/Y 0.07fF
C26125 NOR2X1_LOC_791/Y NOR2X1_LOC_786/a_36_216# 0.00fF
C26126 NAND2X1_LOC_218/B NAND2X1_LOC_23/a_36_24# 0.00fF
C26127 INVX1_LOC_303/A INVX1_LOC_26/A 0.24fF
C26128 NOR2X1_LOC_703/A NOR2X1_LOC_862/B 0.59fF
C26129 INVX1_LOC_199/A INVX1_LOC_139/A 0.03fF
C26130 NAND2X1_LOC_559/Y INVX1_LOC_229/A 0.20fF
C26131 NAND2X1_LOC_571/B INVX1_LOC_18/A 0.03fF
C26132 INVX1_LOC_88/A NOR2X1_LOC_666/A 0.03fF
C26133 INVX1_LOC_103/A NOR2X1_LOC_348/Y 0.02fF
C26134 INPUT_0 NOR2X1_LOC_61/Y 0.18fF
C26135 NAND2X1_LOC_662/Y INVX1_LOC_12/A 0.11fF
C26136 INVX1_LOC_83/A NOR2X1_LOC_258/Y 0.03fF
C26137 NOR2X1_LOC_500/Y INVX1_LOC_290/Y 0.01fF
C26138 INVX1_LOC_45/A NAND2X1_LOC_35/Y 0.02fF
C26139 INVX1_LOC_249/A INVX1_LOC_270/A 0.03fF
C26140 NAND2X1_LOC_53/Y NOR2X1_LOC_454/Y 0.10fF
C26141 NOR2X1_LOC_791/B NOR2X1_LOC_392/Y 0.01fF
C26142 NOR2X1_LOC_208/Y INVX1_LOC_271/A 0.01fF
C26143 NAND2X1_LOC_552/A INVX1_LOC_30/A 0.02fF
C26144 INVX1_LOC_93/A INVX1_LOC_31/A 0.07fF
C26145 NAND2X1_LOC_207/a_36_24# INVX1_LOC_36/A 0.00fF
C26146 INVX1_LOC_245/Y NAND2X1_LOC_149/Y 0.11fF
C26147 NAND2X1_LOC_361/Y NOR2X1_LOC_843/B 0.07fF
C26148 INVX1_LOC_6/Y INVX1_LOC_270/A 0.02fF
C26149 NOR2X1_LOC_500/A INVX1_LOC_23/A 0.01fF
C26150 NAND2X1_LOC_725/A INVX1_LOC_72/A 0.17fF
C26151 INVX1_LOC_5/A INVX1_LOC_30/A 1.94fF
C26152 INVX1_LOC_17/Y INVX1_LOC_172/A 0.01fF
C26153 NOR2X1_LOC_817/a_36_216# INVX1_LOC_269/A 0.01fF
C26154 NOR2X1_LOC_303/Y INVX1_LOC_23/A 0.03fF
C26155 INVX1_LOC_50/A NOR2X1_LOC_577/Y 0.08fF
C26156 INVX1_LOC_17/A NOR2X1_LOC_361/B 0.10fF
C26157 NAND2X1_LOC_214/B INVX1_LOC_36/A 0.07fF
C26158 INVX1_LOC_232/Y NOR2X1_LOC_38/B 0.06fF
C26159 NOR2X1_LOC_703/Y INVX1_LOC_307/Y 0.11fF
C26160 INVX1_LOC_58/A NOR2X1_LOC_152/Y 0.03fF
C26161 INVX1_LOC_163/A NOR2X1_LOC_573/Y 0.05fF
C26162 NOR2X1_LOC_708/Y NAND2X1_LOC_782/B 0.07fF
C26163 D_INPUT_1 NOR2X1_LOC_643/Y 0.36fF
C26164 NAND2X1_LOC_859/B INVX1_LOC_3/Y 0.05fF
C26165 INVX1_LOC_58/A INVX1_LOC_113/Y 0.02fF
C26166 NOR2X1_LOC_405/A INVX1_LOC_38/A 0.03fF
C26167 INVX1_LOC_225/A NAND2X1_LOC_288/B 0.02fF
C26168 INVX1_LOC_256/A INVX1_LOC_103/A 0.14fF
C26169 INVX1_LOC_10/A INVX1_LOC_290/Y 0.07fF
C26170 INVX1_LOC_178/A INVX1_LOC_30/A 2.50fF
C26171 INVX1_LOC_37/Y NAND2X1_LOC_244/A 0.10fF
C26172 INVX1_LOC_36/A INVX1_LOC_27/A 0.15fF
C26173 INVX1_LOC_11/A NOR2X1_LOC_82/A 0.01fF
C26174 INVX1_LOC_6/A NOR2X1_LOC_216/B 0.01fF
C26175 NOR2X1_LOC_739/Y NOR2X1_LOC_307/A 0.30fF
C26176 INVX1_LOC_214/A NAND2X1_LOC_175/Y 0.03fF
C26177 NOR2X1_LOC_667/A NAND2X1_LOC_175/Y 0.12fF
C26178 NOR2X1_LOC_82/A NAND2X1_LOC_381/Y 0.04fF
C26179 NOR2X1_LOC_131/a_36_216# NAND2X1_LOC_454/Y 0.01fF
C26180 NOR2X1_LOC_254/Y INVX1_LOC_23/A 0.73fF
C26181 NAND2X1_LOC_610/a_36_24# INVX1_LOC_26/A 0.00fF
C26182 INVX1_LOC_248/A NAND2X1_LOC_175/Y 0.05fF
C26183 INVX1_LOC_206/A INVX1_LOC_28/Y 0.06fF
C26184 NAND2X1_LOC_721/B NAND2X1_LOC_703/Y -0.07fF
C26185 INVX1_LOC_50/A NOR2X1_LOC_348/B 0.07fF
C26186 NAND2X1_LOC_842/B INVX1_LOC_29/A 0.05fF
C26187 NOR2X1_LOC_655/B INVX1_LOC_23/Y 0.10fF
C26188 INVX1_LOC_221/A INVX1_LOC_57/A 0.01fF
C26189 NAND2X1_LOC_738/B GATE_811 0.04fF
C26190 NAND2X1_LOC_320/a_36_24# NOR2X1_LOC_383/B 0.01fF
C26191 NAND2X1_LOC_72/Y NOR2X1_LOC_577/Y 0.02fF
C26192 INVX1_LOC_256/A INVX1_LOC_292/A 0.01fF
C26193 NOR2X1_LOC_75/Y NOR2X1_LOC_160/B 0.03fF
C26194 NOR2X1_LOC_746/Y INVX1_LOC_92/A 0.15fF
C26195 NAND2X1_LOC_9/Y INVX1_LOC_8/A 0.10fF
C26196 NAND2X1_LOC_778/Y NOR2X1_LOC_238/Y 0.03fF
C26197 INVX1_LOC_222/Y INVX1_LOC_24/A 0.14fF
C26198 INVX1_LOC_34/A NOR2X1_LOC_678/A 0.03fF
C26199 INVX1_LOC_38/A NOR2X1_LOC_857/A 0.10fF
C26200 NOR2X1_LOC_513/Y INVX1_LOC_31/A 0.02fF
C26201 INVX1_LOC_233/A INVX1_LOC_8/A 0.03fF
C26202 NOR2X1_LOC_124/B NOR2X1_LOC_392/Y 0.00fF
C26203 D_INPUT_1 INVX1_LOC_266/Y 0.03fF
C26204 INVX1_LOC_62/A INVX1_LOC_15/A 0.07fF
C26205 INVX1_LOC_6/A NAND2X1_LOC_477/Y 0.76fF
C26206 NOR2X1_LOC_480/A INVX1_LOC_239/A 0.14fF
C26207 NOR2X1_LOC_589/A NOR2X1_LOC_158/Y 0.03fF
C26208 INVX1_LOC_11/A NAND2X1_LOC_36/A 0.34fF
C26209 INVX1_LOC_118/Y INVX1_LOC_46/A 4.86fF
C26210 INVX1_LOC_91/A NOR2X1_LOC_117/a_36_216# 0.01fF
C26211 INVX1_LOC_172/A NOR2X1_LOC_406/A 0.02fF
C26212 INVX1_LOC_54/Y INVX1_LOC_23/A 0.03fF
C26213 NAND2X1_LOC_551/A INVX1_LOC_19/Y 0.16fF
C26214 INVX1_LOC_50/A NOR2X1_LOC_175/B 0.07fF
C26215 NOR2X1_LOC_561/Y NAND2X1_LOC_454/Y 1.84fF
C26216 INVX1_LOC_36/A NAND2X1_LOC_151/a_36_24# 0.01fF
C26217 NAND2X1_LOC_337/B INVX1_LOC_30/A 0.10fF
C26218 INVX1_LOC_37/A INVX1_LOC_118/A 0.25fF
C26219 NOR2X1_LOC_184/a_36_216# NAND2X1_LOC_74/B 0.00fF
C26220 NOR2X1_LOC_220/a_36_216# INVX1_LOC_1/A 0.00fF
C26221 D_GATE_741 INVX1_LOC_142/A 0.05fF
C26222 NOR2X1_LOC_598/B NOR2X1_LOC_537/Y 0.08fF
C26223 INVX1_LOC_224/Y INVX1_LOC_56/A 0.03fF
C26224 NOR2X1_LOC_272/Y INVX1_LOC_33/A 0.49fF
C26225 NOR2X1_LOC_598/B NAND2X1_LOC_338/B 0.02fF
C26226 NOR2X1_LOC_557/A INVX1_LOC_63/A 0.07fF
C26227 INVX1_LOC_237/Y INVX1_LOC_242/A 0.03fF
C26228 INVX1_LOC_50/A INVX1_LOC_22/A 0.23fF
C26229 NOR2X1_LOC_595/a_36_216# INVX1_LOC_312/Y 0.01fF
C26230 INVX1_LOC_123/A INVX1_LOC_19/A 0.19fF
C26231 NOR2X1_LOC_437/a_36_216# INVX1_LOC_88/A 0.00fF
C26232 INVX1_LOC_51/A NAND2X1_LOC_338/B 0.05fF
C26233 INVX1_LOC_232/A NAND2X1_LOC_215/A 0.19fF
C26234 INVX1_LOC_315/Y NAND2X1_LOC_219/B 0.39fF
C26235 NOR2X1_LOC_75/Y NOR2X1_LOC_733/a_36_216# 0.00fF
C26236 NOR2X1_LOC_598/B NAND2X1_LOC_323/B 0.22fF
C26237 INVX1_LOC_58/A NAND2X1_LOC_859/B 0.18fF
C26238 INVX1_LOC_289/Y NOR2X1_LOC_433/A 0.03fF
C26239 NOR2X1_LOC_84/Y INVX1_LOC_306/Y 0.13fF
C26240 INVX1_LOC_27/A NOR2X1_LOC_309/Y 0.03fF
C26241 NAND2X1_LOC_213/A INVX1_LOC_33/A 0.30fF
C26242 NOR2X1_LOC_130/A NAND2X1_LOC_99/A 0.03fF
C26243 NOR2X1_LOC_646/A NOR2X1_LOC_392/Y 0.02fF
C26244 NOR2X1_LOC_269/Y INVX1_LOC_272/A 0.08fF
C26245 NAND2X1_LOC_53/Y INVX1_LOC_77/A 0.07fF
C26246 INVX1_LOC_59/A NOR2X1_LOC_6/B 0.03fF
C26247 NOR2X1_LOC_401/A NOR2X1_LOC_716/B 0.03fF
C26248 NOR2X1_LOC_224/Y INVX1_LOC_22/A 0.07fF
C26249 INVX1_LOC_124/A NAND2X1_LOC_474/Y 0.03fF
C26250 VDD NOR2X1_LOC_430/Y 0.13fF
C26251 INVX1_LOC_215/Y NOR2X1_LOC_152/Y 0.03fF
C26252 INVX1_LOC_311/A INVX1_LOC_32/A 0.72fF
C26253 NOR2X1_LOC_177/Y INVX1_LOC_118/A 0.03fF
C26254 INVX1_LOC_238/A NAND2X1_LOC_866/A 0.04fF
C26255 INVX1_LOC_57/Y NOR2X1_LOC_91/Y 0.21fF
C26256 NOR2X1_LOC_545/B INVX1_LOC_29/A 0.50fF
C26257 NOR2X1_LOC_743/Y INVX1_LOC_118/A 0.07fF
C26258 INVX1_LOC_30/A NOR2X1_LOC_759/a_36_216# 0.00fF
C26259 INVX1_LOC_58/A NAND2X1_LOC_861/Y 0.07fF
C26260 INVX1_LOC_45/A INVX1_LOC_94/A 0.49fF
C26261 NOR2X1_LOC_160/B NOR2X1_LOC_716/B 0.17fF
C26262 INVX1_LOC_20/A INVX1_LOC_264/A 0.00fF
C26263 NAND2X1_LOC_303/Y NOR2X1_LOC_504/Y 0.10fF
C26264 NOR2X1_LOC_391/Y NOR2X1_LOC_38/B 0.01fF
C26265 INVX1_LOC_89/A INVX1_LOC_29/Y 0.07fF
C26266 NAND2X1_LOC_799/A NAND2X1_LOC_799/Y 0.09fF
C26267 INVX1_LOC_94/A NOR2X1_LOC_568/A 0.01fF
C26268 NOR2X1_LOC_103/Y NAND2X1_LOC_465/Y 0.05fF
C26269 NOR2X1_LOC_471/Y INVX1_LOC_153/Y 0.03fF
C26270 NOR2X1_LOC_772/A INVX1_LOC_270/A 0.02fF
C26271 INVX1_LOC_249/A INVX1_LOC_36/A 0.00fF
C26272 INVX1_LOC_21/A INVX1_LOC_9/Y 0.01fF
C26273 NOR2X1_LOC_82/A NOR2X1_LOC_52/B 1.99fF
C26274 INVX1_LOC_50/A NOR2X1_LOC_735/Y 0.01fF
C26275 INVX1_LOC_132/A NOR2X1_LOC_641/B 0.02fF
C26276 INVX1_LOC_252/Y NOR2X1_LOC_6/B 0.03fF
C26277 INVX1_LOC_21/A NAND2X1_LOC_564/B 0.07fF
C26278 INVX1_LOC_6/Y INVX1_LOC_36/A 0.01fF
C26279 D_GATE_366 INVX1_LOC_53/A 0.03fF
C26280 NAND2X1_LOC_198/B NAND2X1_LOC_197/a_36_24# 0.02fF
C26281 NOR2X1_LOC_598/B INVX1_LOC_313/Y 0.01fF
C26282 NAND2X1_LOC_63/Y INVX1_LOC_37/A 0.02fF
C26283 INVX1_LOC_279/A INVX1_LOC_50/Y 0.07fF
C26284 INVX1_LOC_31/A NOR2X1_LOC_84/A 0.48fF
C26285 NOR2X1_LOC_336/B INVX1_LOC_33/A 0.03fF
C26286 NOR2X1_LOC_369/Y NOR2X1_LOC_315/Y 0.06fF
C26287 INVX1_LOC_24/A NAND2X1_LOC_656/A 0.03fF
C26288 NAND2X1_LOC_722/A NOR2X1_LOC_816/A 0.02fF
C26289 NOR2X1_LOC_590/A NOR2X1_LOC_180/Y 0.06fF
C26290 INVX1_LOC_58/A NAND2X1_LOC_661/A 0.01fF
C26291 NOR2X1_LOC_514/A NOR2X1_LOC_514/Y 0.04fF
C26292 NAND2X1_LOC_392/A NOR2X1_LOC_468/Y 0.00fF
C26293 INVX1_LOC_96/A INVX1_LOC_271/Y 0.22fF
C26294 INVX1_LOC_97/Y INVX1_LOC_313/Y -0.02fF
C26295 INVX1_LOC_94/A INVX1_LOC_71/A 0.02fF
C26296 INVX1_LOC_24/A NOR2X1_LOC_484/Y 0.05fF
C26297 INVX1_LOC_136/A NAND2X1_LOC_276/Y 0.26fF
C26298 NAND2X1_LOC_198/B INVX1_LOC_49/A 0.05fF
C26299 NAND2X1_LOC_364/A INVX1_LOC_33/A 0.03fF
C26300 NAND2X1_LOC_787/A INVX1_LOC_140/A 0.05fF
C26301 NAND2X1_LOC_773/Y INVX1_LOC_30/Y 0.05fF
C26302 INVX1_LOC_249/A NOR2X1_LOC_208/Y 0.08fF
C26303 INVX1_LOC_36/A NOR2X1_LOC_664/Y 0.03fF
C26304 NAND2X1_LOC_364/A NOR2X1_LOC_743/a_36_216# 0.00fF
C26305 NAND2X1_LOC_562/B INVX1_LOC_30/A 0.01fF
C26306 INVX1_LOC_11/A NAND2X1_LOC_59/a_36_24# 0.00fF
C26307 NOR2X1_LOC_103/Y INVX1_LOC_56/A 0.03fF
C26308 INVX1_LOC_64/A NOR2X1_LOC_564/Y 0.03fF
C26309 NAND2X1_LOC_721/A NAND2X1_LOC_254/Y 0.02fF
C26310 INVX1_LOC_123/A INVX1_LOC_26/Y 0.16fF
C26311 NOR2X1_LOC_188/A INVX1_LOC_57/A 0.25fF
C26312 INVX1_LOC_6/Y NOR2X1_LOC_208/Y 0.18fF
C26313 NAND2X1_LOC_308/Y INVX1_LOC_72/A 0.10fF
C26314 NAND2X1_LOC_321/a_36_24# INVX1_LOC_196/A 0.06fF
C26315 NOR2X1_LOC_481/A INVX1_LOC_45/Y 0.16fF
C26316 INVX1_LOC_223/Y NOR2X1_LOC_532/Y 0.00fF
C26317 NAND2X1_LOC_543/Y INVX1_LOC_200/A 0.07fF
C26318 NOR2X1_LOC_548/B INVX1_LOC_57/A 0.07fF
C26319 NAND2X1_LOC_58/a_36_24# INVX1_LOC_135/A 0.01fF
C26320 NOR2X1_LOC_435/B NOR2X1_LOC_592/B 0.01fF
C26321 NOR2X1_LOC_557/Y NAND2X1_LOC_656/A 0.02fF
C26322 NOR2X1_LOC_607/A INVX1_LOC_155/Y 0.00fF
C26323 NAND2X1_LOC_227/Y INVX1_LOC_22/A 0.06fF
C26324 NAND2X1_LOC_624/B NAND2X1_LOC_849/A 0.02fF
C26325 INVX1_LOC_37/A INVX1_LOC_257/A 0.00fF
C26326 NOR2X1_LOC_92/Y INVX1_LOC_135/A 0.10fF
C26327 INVX1_LOC_225/Y NOR2X1_LOC_553/Y 0.57fF
C26328 INVX1_LOC_38/A INVX1_LOC_109/Y 0.01fF
C26329 INPUT_0 NOR2X1_LOC_678/A -0.00fF
C26330 NAND2X1_LOC_514/Y NOR2X1_LOC_52/B 0.01fF
C26331 INVX1_LOC_14/A NAND2X1_LOC_656/Y 0.01fF
C26332 NOR2X1_LOC_13/Y NAND2X1_LOC_466/Y 0.02fF
C26333 NOR2X1_LOC_68/A NAND2X1_LOC_629/Y 0.01fF
C26334 INVX1_LOC_157/A INVX1_LOC_103/A 0.03fF
C26335 INVX1_LOC_250/A NAND2X1_LOC_718/a_36_24# 0.00fF
C26336 NOR2X1_LOC_753/Y NAND2X1_LOC_833/Y 0.69fF
C26337 NOR2X1_LOC_510/Y NOR2X1_LOC_171/Y 0.01fF
C26338 NOR2X1_LOC_773/Y INVX1_LOC_30/A 0.10fF
C26339 NAND2X1_LOC_454/Y INVX1_LOC_76/A 0.10fF
C26340 NOR2X1_LOC_631/B NOR2X1_LOC_631/Y 0.02fF
C26341 INVX1_LOC_136/A NAND2X1_LOC_374/Y 0.07fF
C26342 NOR2X1_LOC_433/A NAND2X1_LOC_332/Y 0.11fF
C26343 INVX1_LOC_24/A NOR2X1_LOC_423/Y 0.02fF
C26344 VDD INVX1_LOC_94/Y 0.27fF
C26345 NOR2X1_LOC_470/A NOR2X1_LOC_160/B 0.15fF
C26346 INVX1_LOC_2/A NAND2X1_LOC_198/B 0.08fF
C26347 NOR2X1_LOC_68/A INVX1_LOC_243/A 0.00fF
C26348 NOR2X1_LOC_15/Y INVX1_LOC_175/Y 0.12fF
C26349 INVX1_LOC_54/Y INVX1_LOC_111/A 0.05fF
C26350 NAND2X1_LOC_802/A NOR2X1_LOC_591/Y 0.02fF
C26351 NOR2X1_LOC_226/A NAND2X1_LOC_198/B 0.48fF
C26352 NAND2X1_LOC_794/B NOR2X1_LOC_74/A 0.02fF
C26353 NOR2X1_LOC_717/B NOR2X1_LOC_160/B 0.03fF
C26354 INVX1_LOC_36/A NOR2X1_LOC_695/Y 0.02fF
C26355 INVX1_LOC_36/A INVX1_LOC_137/A 0.05fF
C26356 NAND2X1_LOC_555/Y NAND2X1_LOC_378/a_36_24# 0.01fF
C26357 NOR2X1_LOC_455/a_36_216# NOR2X1_LOC_388/Y 0.00fF
C26358 INVX1_LOC_102/A INVX1_LOC_92/A 0.08fF
C26359 NAND2X1_LOC_468/B NAND2X1_LOC_201/a_36_24# 0.00fF
C26360 NAND2X1_LOC_332/Y INVX1_LOC_151/A 0.00fF
C26361 NOR2X1_LOC_791/B INVX1_LOC_25/Y 0.01fF
C26362 NOR2X1_LOC_222/Y INVX1_LOC_24/A 0.03fF
C26363 NOR2X1_LOC_340/Y NAND2X1_LOC_116/A 0.01fF
C26364 NOR2X1_LOC_426/Y INPUT_5 0.06fF
C26365 INVX1_LOC_290/Y INVX1_LOC_307/A 0.03fF
C26366 NOR2X1_LOC_528/Y NOR2X1_LOC_109/Y 0.46fF
C26367 NOR2X1_LOC_441/Y NOR2X1_LOC_366/Y 0.21fF
C26368 NOR2X1_LOC_68/A NOR2X1_LOC_719/A 0.06fF
C26369 VDD INVX1_LOC_181/A 0.00fF
C26370 NOR2X1_LOC_250/Y INVX1_LOC_28/A 0.03fF
C26371 NOR2X1_LOC_828/A NOR2X1_LOC_160/B 0.07fF
C26372 NOR2X1_LOC_811/B INVX1_LOC_49/A 0.01fF
C26373 VDD INVX1_LOC_296/A 0.34fF
C26374 NAND2X1_LOC_577/A NOR2X1_LOC_130/A 0.20fF
C26375 INVX1_LOC_108/A INVX1_LOC_15/A 0.27fF
C26376 NAND2X1_LOC_198/a_36_24# NOR2X1_LOC_71/Y 0.00fF
C26377 INVX1_LOC_170/A NOR2X1_LOC_71/Y 0.19fF
C26378 NOR2X1_LOC_68/A NOR2X1_LOC_561/Y 0.07fF
C26379 NOR2X1_LOC_446/A INVX1_LOC_182/A 0.20fF
C26380 INVX1_LOC_226/Y INVX1_LOC_77/A 0.07fF
C26381 NOR2X1_LOC_68/A INVX1_LOC_7/A 0.14fF
C26382 INVX1_LOC_314/Y INVX1_LOC_1/Y 0.07fF
C26383 INVX1_LOC_49/A INVX1_LOC_53/Y 0.03fF
C26384 NOR2X1_LOC_619/A INVX1_LOC_49/A 0.05fF
C26385 INVX1_LOC_2/Y NOR2X1_LOC_392/Y 0.08fF
C26386 NOR2X1_LOC_841/A INVX1_LOC_15/A 0.11fF
C26387 NOR2X1_LOC_679/B INVX1_LOC_22/A 0.02fF
C26388 NAND2X1_LOC_53/Y NAND2X1_LOC_832/Y 0.02fF
C26389 INVX1_LOC_17/A INVX1_LOC_285/Y 0.01fF
C26390 D_INPUT_0 NOR2X1_LOC_744/Y 0.06fF
C26391 INVX1_LOC_130/A INVX1_LOC_75/A 0.06fF
C26392 INVX1_LOC_135/A NAND2X1_LOC_837/Y 0.01fF
C26393 NOR2X1_LOC_121/Y INVX1_LOC_16/A 0.01fF
C26394 INVX1_LOC_77/A INVX1_LOC_10/A 0.25fF
C26395 INVX1_LOC_36/A NOR2X1_LOC_19/B 0.31fF
C26396 INVX1_LOC_30/A INVX1_LOC_140/A 0.17fF
C26397 INVX1_LOC_284/A INVX1_LOC_29/A 0.03fF
C26398 INVX1_LOC_145/Y INVX1_LOC_49/A 0.01fF
C26399 INVX1_LOC_238/Y INVX1_LOC_282/A 0.00fF
C26400 INVX1_LOC_18/A NAND2X1_LOC_654/B 0.03fF
C26401 INVX1_LOC_72/A NAND2X1_LOC_560/A 0.03fF
C26402 INVX1_LOC_304/Y NAND2X1_LOC_543/Y 0.12fF
C26403 INVX1_LOC_12/A INVX1_LOC_290/Y 0.07fF
C26404 INVX1_LOC_2/A NOR2X1_LOC_219/Y 0.50fF
C26405 NOR2X1_LOC_15/Y INVX1_LOC_95/Y 0.10fF
C26406 INVX1_LOC_45/A INVX1_LOC_144/A 0.08fF
C26407 NAND2X1_LOC_338/B NAND2X1_LOC_528/a_36_24# 0.00fF
C26408 INVX1_LOC_254/Y INVX1_LOC_90/A 0.00fF
C26409 INVX1_LOC_41/A INVX1_LOC_135/A 0.08fF
C26410 INVX1_LOC_24/A NOR2X1_LOC_329/B 0.13fF
C26411 NAND2X1_LOC_226/a_36_24# NOR2X1_LOC_814/A 0.01fF
C26412 NOR2X1_LOC_717/B NOR2X1_LOC_317/B 0.16fF
C26413 NOR2X1_LOC_490/Y NAND2X1_LOC_837/Y 0.01fF
C26414 NOR2X1_LOC_655/B INVX1_LOC_232/A 0.10fF
C26415 INVX1_LOC_201/Y INVX1_LOC_135/A 1.63fF
C26416 NOR2X1_LOC_226/A INVX1_LOC_53/Y 0.98fF
C26417 NOR2X1_LOC_67/A NOR2X1_LOC_62/a_36_216# 0.00fF
C26418 INVX1_LOC_208/A NOR2X1_LOC_757/Y 0.02fF
C26419 NOR2X1_LOC_46/a_36_216# NOR2X1_LOC_48/B 0.03fF
C26420 NOR2X1_LOC_216/B INVX1_LOC_270/A 0.01fF
C26421 NOR2X1_LOC_493/B INVX1_LOC_101/A 0.04fF
C26422 INVX1_LOC_305/A INPUT_0 0.07fF
C26423 INVX1_LOC_205/Y VDD 0.26fF
C26424 INVX1_LOC_256/A NOR2X1_LOC_141/a_36_216# 0.00fF
C26425 INVX1_LOC_2/A NOR2X1_LOC_665/A 0.17fF
C26426 INVX1_LOC_15/A INPUT_7 0.02fF
C26427 INVX1_LOC_58/A NAND2X1_LOC_802/Y 0.07fF
C26428 INVX1_LOC_124/A INVX1_LOC_10/A 0.93fF
C26429 INVX1_LOC_200/Y NAND2X1_LOC_489/a_36_24# 0.00fF
C26430 NAND2X1_LOC_116/A NOR2X1_LOC_99/B 0.07fF
C26431 NOR2X1_LOC_15/Y NOR2X1_LOC_305/Y 0.03fF
C26432 NOR2X1_LOC_831/B INVX1_LOC_270/Y 0.01fF
C26433 INVX1_LOC_11/A INVX1_LOC_59/Y 0.03fF
C26434 NOR2X1_LOC_458/a_36_216# NOR2X1_LOC_155/A -0.00fF
C26435 NOR2X1_LOC_202/a_36_216# NOR2X1_LOC_357/Y 0.00fF
C26436 NOR2X1_LOC_219/Y NOR2X1_LOC_218/Y 0.02fF
C26437 NOR2X1_LOC_701/a_36_216# INVX1_LOC_22/A 0.01fF
C26438 INVX1_LOC_133/A INVX1_LOC_94/Y 0.06fF
C26439 NOR2X1_LOC_82/A INVX1_LOC_74/A 0.02fF
C26440 NOR2X1_LOC_210/a_36_216# INVX1_LOC_37/A 0.00fF
C26441 NOR2X1_LOC_68/A NOR2X1_LOC_167/Y 0.02fF
C26442 NOR2X1_LOC_424/Y INVX1_LOC_189/A 0.09fF
C26443 INVX1_LOC_299/A VDD 0.33fF
C26444 INVX1_LOC_89/A INVX1_LOC_60/Y 0.68fF
C26445 NOR2X1_LOC_220/a_36_216# NOR2X1_LOC_188/A 0.12fF
C26446 INVX1_LOC_11/A INVX1_LOC_176/A 0.02fF
C26447 NOR2X1_LOC_355/A NOR2X1_LOC_493/B 0.00fF
C26448 NOR2X1_LOC_65/B NAND2X1_LOC_475/Y 0.18fF
C26449 INVX1_LOC_27/A NOR2X1_LOC_865/A 0.61fF
C26450 INVX1_LOC_144/A INVX1_LOC_71/A 0.02fF
C26451 NOR2X1_LOC_147/B INVX1_LOC_311/Y 0.02fF
C26452 NOR2X1_LOC_92/Y NOR2X1_LOC_813/Y 0.07fF
C26453 NOR2X1_LOC_538/B VDD 0.42fF
C26454 NOR2X1_LOC_392/Y NOR2X1_LOC_608/Y -0.03fF
C26455 NAND2X1_LOC_579/A INVX1_LOC_33/Y 0.02fF
C26456 NAND2X1_LOC_361/Y INVX1_LOC_31/Y 0.03fF
C26457 NOR2X1_LOC_83/Y INVX1_LOC_71/A 0.08fF
C26458 NOR2X1_LOC_309/Y NOR2X1_LOC_772/A 0.00fF
C26459 NOR2X1_LOC_500/Y NOR2X1_LOC_549/a_36_216# 0.00fF
C26460 INVX1_LOC_132/A NOR2X1_LOC_751/A 0.00fF
C26461 INVX1_LOC_215/A NAND2X1_LOC_112/Y 0.05fF
C26462 INVX1_LOC_271/A INVX1_LOC_63/A 0.03fF
C26463 NAND2X1_LOC_796/B INVX1_LOC_54/A 0.01fF
C26464 NOR2X1_LOC_92/Y INVX1_LOC_280/A 0.03fF
C26465 INVX1_LOC_293/A VDD -0.00fF
C26466 NOR2X1_LOC_92/Y NOR2X1_LOC_94/Y 0.08fF
C26467 INVX1_LOC_50/A INVX1_LOC_186/Y 0.04fF
C26468 NOR2X1_LOC_717/B NOR2X1_LOC_516/B 0.05fF
C26469 NOR2X1_LOC_78/B D_GATE_366 0.03fF
C26470 INVX1_LOC_232/A NOR2X1_LOC_99/B 0.17fF
C26471 INVX1_LOC_5/A INVX1_LOC_113/A 0.07fF
C26472 NOR2X1_LOC_533/Y NOR2X1_LOC_536/A 0.08fF
C26473 D_INPUT_0 INVX1_LOC_16/A 0.18fF
C26474 NOR2X1_LOC_544/A INVX1_LOC_196/Y 0.05fF
C26475 NOR2X1_LOC_209/Y NOR2X1_LOC_828/B 0.03fF
C26476 D_INPUT_1 INVX1_LOC_19/A 0.03fF
C26477 NAND2X1_LOC_214/B NAND2X1_LOC_609/a_36_24# 0.00fF
C26478 INVX1_LOC_222/Y NOR2X1_LOC_197/B 0.03fF
C26479 INVX1_LOC_24/A INPUT_4 0.05fF
C26480 NOR2X1_LOC_524/Y VDD 0.20fF
C26481 NOR2X1_LOC_246/A NOR2X1_LOC_589/A 0.06fF
C26482 NAND2X1_LOC_53/Y INVX1_LOC_9/A 0.07fF
C26483 INVX1_LOC_314/Y INVX1_LOC_93/Y 0.01fF
C26484 INVX1_LOC_35/A NAND2X1_LOC_773/B 0.04fF
C26485 NAND2X1_LOC_207/a_36_24# INVX1_LOC_63/A 0.00fF
C26486 NOR2X1_LOC_68/A INVX1_LOC_76/A 0.31fF
C26487 INVX1_LOC_49/Y NAND2X1_LOC_590/a_36_24# 0.00fF
C26488 NOR2X1_LOC_160/B NOR2X1_LOC_707/A 0.22fF
C26489 INVX1_LOC_190/A INVX1_LOC_10/A 0.02fF
C26490 NAND2X1_LOC_214/B INVX1_LOC_63/A 0.10fF
C26491 INVX1_LOC_64/A INVX1_LOC_264/A 0.00fF
C26492 NOR2X1_LOC_653/Y NOR2X1_LOC_652/Y 0.00fF
C26493 NAND2X1_LOC_727/Y INVX1_LOC_28/A 0.02fF
C26494 INVX1_LOC_77/A NOR2X1_LOC_799/B 0.01fF
C26495 INVX1_LOC_75/A NAND2X1_LOC_672/B 0.06fF
C26496 INVX1_LOC_33/A NOR2X1_LOC_405/A 0.10fF
C26497 NOR2X1_LOC_160/B NOR2X1_LOC_209/B 0.03fF
C26498 NOR2X1_LOC_590/Y INVX1_LOC_186/Y 0.02fF
C26499 INVX1_LOC_28/A NAND2X1_LOC_660/Y 1.01fF
C26500 NOR2X1_LOC_743/a_36_216# NOR2X1_LOC_405/A 0.01fF
C26501 NOR2X1_LOC_309/Y NOR2X1_LOC_528/Y -0.04fF
C26502 NAND2X1_LOC_191/a_36_24# INVX1_LOC_307/A 0.00fF
C26503 NAND2X1_LOC_569/B NAND2X1_LOC_74/B 0.13fF
C26504 NOR2X1_LOC_516/B NOR2X1_LOC_151/Y 0.02fF
C26505 INVX1_LOC_27/A INVX1_LOC_63/A 5.76fF
C26506 NAND2X1_LOC_352/a_36_24# NOR2X1_LOC_743/Y 0.00fF
C26507 NAND2X1_LOC_787/A INVX1_LOC_42/A 1.51fF
C26508 INVX1_LOC_215/Y INVX1_LOC_291/A 0.01fF
C26509 INVX1_LOC_83/A D_GATE_366 0.07fF
C26510 NAND2X1_LOC_363/B INVX1_LOC_42/A 0.03fF
C26511 NAND2X1_LOC_519/a_36_24# INVX1_LOC_226/A 0.00fF
C26512 NAND2X1_LOC_783/A NOR2X1_LOC_329/B 0.10fF
C26513 INVX1_LOC_245/A NOR2X1_LOC_589/Y 0.07fF
C26514 D_INPUT_0 INVX1_LOC_28/A 0.16fF
C26515 NAND2X1_LOC_51/B GATE_662 0.03fF
C26516 INVX1_LOC_78/A NOR2X1_LOC_135/a_36_216# 0.00fF
C26517 INVX1_LOC_31/A NOR2X1_LOC_78/Y 0.01fF
C26518 NOR2X1_LOC_215/Y INVX1_LOC_281/A 0.02fF
C26519 NAND2X1_LOC_342/Y INVX1_LOC_91/A 0.11fF
C26520 NOR2X1_LOC_329/B NOR2X1_LOC_130/A 0.12fF
C26521 INVX1_LOC_33/A NOR2X1_LOC_857/A 0.07fF
C26522 INVX1_LOC_90/A NOR2X1_LOC_597/A 0.02fF
C26523 INVX1_LOC_174/Y INVX1_LOC_86/A 0.00fF
C26524 INVX1_LOC_265/A NAND2X1_LOC_650/B 0.18fF
C26525 NOR2X1_LOC_789/A INVX1_LOC_48/A 0.03fF
C26526 INVX1_LOC_162/A VDD 0.25fF
C26527 NOR2X1_LOC_400/A INVX1_LOC_32/A 0.02fF
C26528 NAND2X1_LOC_837/Y INVX1_LOC_280/A 0.01fF
C26529 NOR2X1_LOC_456/Y NOR2X1_LOC_334/Y 0.02fF
C26530 NOR2X1_LOC_624/A INVX1_LOC_37/A 0.22fF
C26531 INVX1_LOC_223/A INVX1_LOC_92/A 0.07fF
C26532 NAND2X1_LOC_198/B INVX1_LOC_118/A 0.24fF
C26533 INVX1_LOC_45/A NOR2X1_LOC_155/A 0.24fF
C26534 NOR2X1_LOC_454/Y INVX1_LOC_12/A 0.19fF
C26535 NOR2X1_LOC_532/Y INVX1_LOC_75/A 0.01fF
C26536 INVX1_LOC_36/A NOR2X1_LOC_216/B 0.01fF
C26537 NAND2X1_LOC_787/A INVX1_LOC_78/A 0.03fF
C26538 NAND2X1_LOC_796/B NOR2X1_LOC_48/B 0.03fF
C26539 INVX1_LOC_1/Y NOR2X1_LOC_557/A 0.07fF
C26540 NOR2X1_LOC_315/Y VDD 1.44fF
C26541 NAND2X1_LOC_363/B INVX1_LOC_78/A 0.07fF
C26542 NOR2X1_LOC_667/A NOR2X1_LOC_279/Y 0.01fF
C26543 NAND2X1_LOC_785/Y NAND2X1_LOC_804/Y -0.01fF
C26544 NOR2X1_LOC_843/B NOR2X1_LOC_105/Y 0.12fF
C26545 INVX1_LOC_271/A NOR2X1_LOC_65/Y 0.03fF
C26546 NOR2X1_LOC_140/A NOR2X1_LOC_847/B 0.03fF
C26547 NOR2X1_LOC_335/B NOR2X1_LOC_355/a_36_216# 0.00fF
C26548 NOR2X1_LOC_626/Y INVX1_LOC_32/A 0.03fF
C26549 INVX1_LOC_112/Y NAND2X1_LOC_215/A 0.24fF
C26550 NOR2X1_LOC_216/Y NOR2X1_LOC_329/B 0.09fF
C26551 NOR2X1_LOC_392/B NOR2X1_LOC_440/a_36_216# 0.12fF
C26552 INVX1_LOC_310/A VDD 0.12fF
C26553 INVX1_LOC_263/A INVX1_LOC_247/A 0.05fF
C26554 NOR2X1_LOC_250/A NAND2X1_LOC_74/B 0.03fF
C26555 NOR2X1_LOC_432/Y VDD 0.12fF
C26556 NOR2X1_LOC_91/A NAND2X1_LOC_860/A 0.07fF
C26557 INVX1_LOC_103/A NOR2X1_LOC_89/A 0.01fF
C26558 NAND2X1_LOC_785/B INVX1_LOC_84/A 0.12fF
C26559 NAND2X1_LOC_564/B INVX1_LOC_304/A 0.07fF
C26560 NAND2X1_LOC_717/Y NAND2X1_LOC_839/a_36_24# 0.00fF
C26561 NAND2X1_LOC_721/B INVX1_LOC_119/Y 0.02fF
C26562 NOR2X1_LOC_396/Y NAND2X1_LOC_735/B 0.00fF
C26563 INVX1_LOC_82/Y INVX1_LOC_75/A 0.03fF
C26564 NOR2X1_LOC_431/Y NAND2X1_LOC_798/B 0.01fF
C26565 INVX1_LOC_13/Y NAND2X1_LOC_471/Y 0.07fF
C26566 INVX1_LOC_2/A INVX1_LOC_77/Y 0.07fF
C26567 NAND2X1_LOC_784/A INVX1_LOC_57/A 0.00fF
C26568 INVX1_LOC_71/A NOR2X1_LOC_155/A 0.13fF
C26569 NAND2X1_LOC_840/B NOR2X1_LOC_305/Y 0.06fF
C26570 NOR2X1_LOC_65/B NAND2X1_LOC_363/B 0.01fF
C26571 INVX1_LOC_77/A INVX1_LOC_307/A 0.07fF
C26572 INVX1_LOC_197/A INVX1_LOC_194/Y 0.00fF
C26573 INVX1_LOC_52/A VDD 0.12fF
C26574 NOR2X1_LOC_82/A NAND2X1_LOC_254/Y 0.22fF
C26575 NOR2X1_LOC_667/A NAND2X1_LOC_804/Y 0.38fF
C26576 NOR2X1_LOC_33/A NOR2X1_LOC_35/Y 0.42fF
C26577 NAND2X1_LOC_725/A NAND2X1_LOC_402/B 0.00fF
C26578 INVX1_LOC_279/A INVX1_LOC_188/Y 0.01fF
C26579 NOR2X1_LOC_360/Y NOR2X1_LOC_673/A 0.20fF
C26580 INVX1_LOC_292/A NOR2X1_LOC_89/A 0.03fF
C26581 INVX1_LOC_13/A INVX1_LOC_20/A 0.03fF
C26582 NAND2X1_LOC_860/A INVX1_LOC_23/A 0.09fF
C26583 INVX1_LOC_77/A NOR2X1_LOC_445/B 0.16fF
C26584 INVX1_LOC_207/Y INVX1_LOC_167/Y 0.12fF
C26585 INVX1_LOC_268/Y VDD 0.21fF
C26586 NOR2X1_LOC_589/A NOR2X1_LOC_357/Y 1.19fF
C26587 NOR2X1_LOC_810/A INVX1_LOC_143/Y 0.00fF
C26588 NOR2X1_LOC_381/Y NOR2X1_LOC_38/B 0.60fF
C26589 NAND2X1_LOC_239/a_36_24# INVX1_LOC_118/A 0.00fF
C26590 NAND2X1_LOC_357/B INVX1_LOC_185/A 0.02fF
C26591 INVX1_LOC_27/A NAND2X1_LOC_223/B 0.04fF
C26592 NAND2X1_LOC_860/A NOR2X1_LOC_277/a_36_216# 0.00fF
C26593 NOR2X1_LOC_15/Y INVX1_LOC_271/Y 0.08fF
C26594 NOR2X1_LOC_781/B NOR2X1_LOC_586/Y 0.02fF
C26595 NOR2X1_LOC_781/A NAND2X1_LOC_637/a_36_24# 0.01fF
C26596 INVX1_LOC_245/A INVX1_LOC_117/A 0.05fF
C26597 INVX1_LOC_72/A INVX1_LOC_29/A 0.18fF
C26598 NAND2X1_LOC_500/Y NAND2X1_LOC_254/Y 0.07fF
C26599 D_INPUT_0 NOR2X1_LOC_35/Y 0.03fF
C26600 NAND2X1_LOC_123/Y NOR2X1_LOC_318/B 0.01fF
C26601 INVX1_LOC_85/A INVX1_LOC_92/A 0.00fF
C26602 NOR2X1_LOC_361/B INVX1_LOC_94/Y 0.04fF
C26603 INVX1_LOC_45/A NOR2X1_LOC_833/B 0.21fF
C26604 INVX1_LOC_174/A INVX1_LOC_32/A 0.02fF
C26605 INVX1_LOC_17/A INVX1_LOC_4/Y 0.26fF
C26606 INVX1_LOC_104/A NOR2X1_LOC_862/B 0.02fF
C26607 INVX1_LOC_83/A INVX1_LOC_36/Y 0.03fF
C26608 NOR2X1_LOC_309/Y NOR2X1_LOC_216/B 0.01fF
C26609 NOR2X1_LOC_616/Y NOR2X1_LOC_629/Y 0.00fF
C26610 NOR2X1_LOC_246/A INVX1_LOC_20/A 0.10fF
C26611 INVX1_LOC_54/Y NOR2X1_LOC_79/A 0.01fF
C26612 NOR2X1_LOC_237/Y NAND2X1_LOC_477/Y 1.68fF
C26613 NAND2X1_LOC_848/A INVX1_LOC_16/A 0.07fF
C26614 INVX1_LOC_30/A INVX1_LOC_42/A 0.13fF
C26615 INVX1_LOC_25/A INVX1_LOC_306/Y 0.03fF
C26616 VDD INVX1_LOC_66/A 0.12fF
C26617 D_INPUT_2 INVX1_LOC_19/A 0.04fF
C26618 NOR2X1_LOC_500/Y INVX1_LOC_9/A 0.14fF
C26619 INVX1_LOC_226/Y INVX1_LOC_9/A 0.07fF
C26620 NAND2X1_LOC_551/A INVX1_LOC_20/A 0.20fF
C26621 INVX1_LOC_67/Y INVX1_LOC_91/A 0.01fF
C26622 NOR2X1_LOC_457/A INVX1_LOC_78/A 6.96fF
C26623 INVX1_LOC_90/A NOR2X1_LOC_825/Y 0.13fF
C26624 NOR2X1_LOC_163/A INVX1_LOC_76/A 0.06fF
C26625 NOR2X1_LOC_111/A NOR2X1_LOC_110/a_36_216# 0.05fF
C26626 INVX1_LOC_280/Y NOR2X1_LOC_630/a_36_216# 0.00fF
C26627 NOR2X1_LOC_290/Y INVX1_LOC_35/Y 0.06fF
C26628 INVX1_LOC_32/Y INVX1_LOC_193/A 0.01fF
C26629 INVX1_LOC_53/Y INVX1_LOC_118/A 0.02fF
C26630 NOR2X1_LOC_91/A NAND2X1_LOC_537/Y 0.07fF
C26631 VDD NAND2X1_LOC_624/A 0.00fF
C26632 INVX1_LOC_182/Y INVX1_LOC_188/Y 0.01fF
C26633 NOR2X1_LOC_468/Y NOR2X1_LOC_72/Y 0.00fF
C26634 NOR2X1_LOC_256/a_36_216# INVX1_LOC_284/A 0.01fF
C26635 D_GATE_366 INVX1_LOC_46/A 0.03fF
C26636 NOR2X1_LOC_419/Y NAND2X1_LOC_207/B 0.03fF
C26637 NAND2X1_LOC_323/B NOR2X1_LOC_634/A 0.05fF
C26638 INVX1_LOC_286/A INVX1_LOC_98/A 0.07fF
C26639 VDD NOR2X1_LOC_166/Y 0.14fF
C26640 INVX1_LOC_77/A INVX1_LOC_12/A 0.10fF
C26641 INVX1_LOC_56/Y NAND2X1_LOC_93/B 0.05fF
C26642 INVX1_LOC_93/A NOR2X1_LOC_109/Y 0.00fF
C26643 INVX1_LOC_286/A NOR2X1_LOC_78/A 0.07fF
C26644 INVX1_LOC_10/A INVX1_LOC_9/A 0.10fF
C26645 NOR2X1_LOC_708/B INVX1_LOC_301/A 0.01fF
C26646 D_INPUT_1 NOR2X1_LOC_122/A 0.48fF
C26647 NOR2X1_LOC_210/B NOR2X1_LOC_156/Y 0.00fF
C26648 NOR2X1_LOC_279/a_36_216# INVX1_LOC_285/A 0.01fF
C26649 NAND2X1_LOC_21/Y INPUT_7 0.04fF
C26650 NOR2X1_LOC_687/Y INVX1_LOC_307/A 0.07fF
C26651 NOR2X1_LOC_71/Y NOR2X1_LOC_271/Y 0.07fF
C26652 INVX1_LOC_147/A INVX1_LOC_76/A 0.01fF
C26653 NAND2X1_LOC_662/Y INVX1_LOC_92/A 0.00fF
C26654 NOR2X1_LOC_709/A INVX1_LOC_293/Y 1.49fF
C26655 NOR2X1_LOC_585/a_36_216# NOR2X1_LOC_158/Y 0.01fF
C26656 INVX1_LOC_30/A INVX1_LOC_78/A 1.42fF
C26657 NOR2X1_LOC_140/A NOR2X1_LOC_660/Y 0.03fF
C26658 INVX1_LOC_33/A INVX1_LOC_109/Y 0.01fF
C26659 NAND2X1_LOC_392/Y INVX1_LOC_70/A 0.01fF
C26660 INVX1_LOC_14/A NOR2X1_LOC_717/A 0.14fF
C26661 NAND2X1_LOC_807/A INVX1_LOC_57/A 0.01fF
C26662 INVX1_LOC_206/Y INVX1_LOC_247/A 0.03fF
C26663 INVX1_LOC_75/A NAND2X1_LOC_129/a_36_24# 0.01fF
C26664 INVX1_LOC_8/A INVX1_LOC_284/A 0.07fF
C26665 D_INPUT_1 INVX1_LOC_161/Y 0.07fF
C26666 INVX1_LOC_143/A NOR2X1_LOC_691/B 0.03fF
C26667 INVX1_LOC_28/A NAND2X1_LOC_848/A 0.17fF
C26668 INVX1_LOC_239/A INVX1_LOC_253/Y 0.20fF
C26669 NOR2X1_LOC_207/a_36_216# INVX1_LOC_54/A 0.00fF
C26670 INVX1_LOC_95/A INVX1_LOC_98/A 0.00fF
C26671 NAND2X1_LOC_352/B INVX1_LOC_270/Y 0.02fF
C26672 NOR2X1_LOC_456/a_36_216# INVX1_LOC_50/Y 0.01fF
C26673 INVX1_LOC_75/A NOR2X1_LOC_363/Y 0.05fF
C26674 NOR2X1_LOC_709/A NAND2X1_LOC_74/B 0.07fF
C26675 NAND2X1_LOC_567/Y INVX1_LOC_231/A 0.09fF
C26676 NOR2X1_LOC_598/B NOR2X1_LOC_541/Y 0.02fF
C26677 INVX1_LOC_124/A INVX1_LOC_12/A 2.27fF
C26678 NOR2X1_LOC_65/B INVX1_LOC_30/A 0.17fF
C26679 NOR2X1_LOC_172/Y INVX1_LOC_15/A 0.03fF
C26680 INVX1_LOC_1/A INVX1_LOC_306/Y 0.10fF
C26681 NOR2X1_LOC_537/Y INVX1_LOC_29/A 0.03fF
C26682 NOR2X1_LOC_302/Y INVX1_LOC_9/A 0.04fF
C26683 NAND2X1_LOC_338/B INVX1_LOC_29/A 0.14fF
C26684 NOR2X1_LOC_721/Y NAND2X1_LOC_96/A 0.00fF
C26685 NOR2X1_LOC_600/Y INVX1_LOC_247/A 0.11fF
C26686 NOR2X1_LOC_147/B INVX1_LOC_15/A 0.17fF
C26687 INVX1_LOC_314/Y INVX1_LOC_87/A 0.08fF
C26688 NOR2X1_LOC_550/B NOR2X1_LOC_334/Y 0.10fF
C26689 NAND2X1_LOC_132/a_36_24# INVX1_LOC_9/A 0.01fF
C26690 NAND2X1_LOC_777/a_36_24# INVX1_LOC_141/Y 0.00fF
C26691 NOR2X1_LOC_147/A INVX1_LOC_117/A 0.03fF
C26692 NOR2X1_LOC_415/a_36_216# NAND2X1_LOC_141/Y 0.08fF
C26693 INVX1_LOC_135/A NAND2X1_LOC_574/A 0.12fF
C26694 INVX1_LOC_144/A NOR2X1_LOC_331/B 0.17fF
C26695 INVX1_LOC_50/A INVX1_LOC_18/A 0.13fF
C26696 NAND2X1_LOC_656/Y NOR2X1_LOC_127/Y 0.01fF
C26697 INVX1_LOC_90/A NOR2X1_LOC_88/Y 0.28fF
C26698 NAND2X1_LOC_728/Y INVX1_LOC_50/A 0.07fF
C26699 NOR2X1_LOC_124/a_36_216# INVX1_LOC_74/A 0.02fF
C26700 INVX1_LOC_45/A NOR2X1_LOC_598/B 2.81fF
C26701 NOR2X1_LOC_403/a_36_216# INVX1_LOC_26/A 0.00fF
C26702 INVX1_LOC_223/A INVX1_LOC_53/A 0.05fF
C26703 INVX1_LOC_303/A NAND2X1_LOC_616/a_36_24# 0.00fF
C26704 INVX1_LOC_74/A INVX1_LOC_59/Y 0.03fF
C26705 NOR2X1_LOC_598/B NOR2X1_LOC_568/A 0.38fF
C26706 NOR2X1_LOC_6/B NOR2X1_LOC_38/B 0.09fF
C26707 NAND2X1_LOC_773/Y NOR2X1_LOC_15/Y 0.01fF
C26708 NOR2X1_LOC_80/a_36_216# INVX1_LOC_46/A 0.00fF
C26709 INVX1_LOC_50/A NAND2X1_LOC_711/B 0.10fF
C26710 NOR2X1_LOC_152/Y NOR2X1_LOC_135/a_36_216# 0.01fF
C26711 NOR2X1_LOC_355/a_36_216# INVX1_LOC_84/A 0.00fF
C26712 NOR2X1_LOC_160/B NOR2X1_LOC_343/B 0.01fF
C26713 INVX1_LOC_13/A NOR2X1_LOC_128/A 0.01fF
C26714 INVX1_LOC_90/A INVX1_LOC_84/A 0.41fF
C26715 INVX1_LOC_88/A NOR2X1_LOC_359/a_36_216# 0.00fF
C26716 NAND2X1_LOC_834/a_36_24# NOR2X1_LOC_48/B 0.00fF
C26717 INVX1_LOC_94/A NOR2X1_LOC_493/A 0.04fF
C26718 INVX1_LOC_37/A NAND2X1_LOC_212/Y 0.02fF
C26719 NAND2X1_LOC_725/A NAND2X1_LOC_856/A 0.11fF
C26720 NOR2X1_LOC_382/Y INVX1_LOC_5/A 0.07fF
C26721 NOR2X1_LOC_389/B INVX1_LOC_84/A 0.07fF
C26722 INVX1_LOC_50/A INVX1_LOC_172/A 0.03fF
C26723 INVX1_LOC_200/Y NAND2X1_LOC_374/a_36_24# 0.00fF
C26724 INVX1_LOC_136/A NAND2X1_LOC_569/B 0.20fF
C26725 INVX1_LOC_16/A NOR2X1_LOC_754/A 0.04fF
C26726 NOR2X1_LOC_585/Y NOR2X1_LOC_586/Y 0.13fF
C26727 D_INPUT_1 NOR2X1_LOC_437/Y 0.16fF
C26728 NAND2X1_LOC_796/B NOR2X1_LOC_441/Y 0.91fF
C26729 INVX1_LOC_64/A NOR2X1_LOC_759/A 0.03fF
C26730 INVX1_LOC_27/A NOR2X1_LOC_606/a_36_216# 0.02fF
C26731 INVX1_LOC_144/A NOR2X1_LOC_592/B 0.21fF
C26732 NOR2X1_LOC_598/B INVX1_LOC_71/A 0.07fF
C26733 INVX1_LOC_36/A INVX1_LOC_93/A 0.46fF
C26734 INVX1_LOC_11/A INVX1_LOC_103/A 0.19fF
C26735 INVX1_LOC_35/A INVX1_LOC_24/A 0.15fF
C26736 INVX1_LOC_27/A NOR2X1_LOC_688/Y 0.01fF
C26737 INVX1_LOC_31/A NAND2X1_LOC_473/A 0.18fF
C26738 NAND2X1_LOC_661/a_36_24# INVX1_LOC_117/Y 0.00fF
C26739 NOR2X1_LOC_590/Y INVX1_LOC_18/A 0.18fF
C26740 NOR2X1_LOC_19/B INVX1_LOC_63/A 0.04fF
C26741 INVX1_LOC_88/Y NOR2X1_LOC_383/B 0.14fF
C26742 INVX1_LOC_14/Y INVX1_LOC_37/A 0.04fF
C26743 NAND2X1_LOC_348/A INVX1_LOC_84/A 0.05fF
C26744 NOR2X1_LOC_589/A INVX1_LOC_32/A 0.10fF
C26745 INVX1_LOC_313/Y INVX1_LOC_29/A 0.11fF
C26746 NOR2X1_LOC_486/B INVX1_LOC_23/A 0.06fF
C26747 NAND2X1_LOC_537/Y INVX1_LOC_31/A 0.07fF
C26748 NAND2X1_LOC_866/B NOR2X1_LOC_824/a_36_216# 0.00fF
C26749 INVX1_LOC_25/A INVX1_LOC_294/Y 0.03fF
C26750 NAND2X1_LOC_377/Y INVX1_LOC_32/A 0.07fF
C26751 NOR2X1_LOC_244/a_36_216# NOR2X1_LOC_342/B 0.03fF
C26752 INVX1_LOC_13/A INVX1_LOC_4/A 0.12fF
C26753 NOR2X1_LOC_516/Y INVX1_LOC_23/A 0.03fF
C26754 VDD NAND2X1_LOC_96/A 0.01fF
C26755 INVX1_LOC_263/A NOR2X1_LOC_465/Y 0.75fF
C26756 INVX1_LOC_11/A INVX1_LOC_292/A 0.07fF
C26757 NOR2X1_LOC_349/A NAND2X1_LOC_258/a_36_24# 0.00fF
C26758 NOR2X1_LOC_168/B NOR2X1_LOC_383/B 0.10fF
C26759 NAND2X1_LOC_465/A INVX1_LOC_118/A 0.03fF
C26760 NOR2X1_LOC_473/B NOR2X1_LOC_114/Y 0.11fF
C26761 NOR2X1_LOC_425/Y NOR2X1_LOC_694/Y 0.07fF
C26762 NAND2X1_LOC_11/Y NOR2X1_LOC_635/B 0.13fF
C26763 NOR2X1_LOC_96/Y NOR2X1_LOC_825/Y 0.17fF
C26764 NOR2X1_LOC_211/A NOR2X1_LOC_541/B 0.07fF
C26765 INVX1_LOC_171/A INVX1_LOC_32/A 3.34fF
C26766 NOR2X1_LOC_114/A NOR2X1_LOC_814/A 0.02fF
C26767 NAND2X1_LOC_860/A NOR2X1_LOC_290/Y 0.32fF
C26768 INVX1_LOC_91/A INVX1_LOC_285/A 0.10fF
C26769 NOR2X1_LOC_612/B NOR2X1_LOC_717/A 0.03fF
C26770 INVX1_LOC_90/A INVX1_LOC_15/A 0.17fF
C26771 INVX1_LOC_266/Y NOR2X1_LOC_678/A 0.05fF
C26772 NOR2X1_LOC_528/Y NOR2X1_LOC_654/a_36_216# 0.00fF
C26773 INVX1_LOC_136/A NOR2X1_LOC_250/A 0.03fF
C26774 NOR2X1_LOC_35/Y INVX1_LOC_46/Y 0.10fF
C26775 INVX1_LOC_111/Y NOR2X1_LOC_717/A 0.02fF
C26776 INVX1_LOC_91/A NOR2X1_LOC_814/A 0.16fF
C26777 INVX1_LOC_229/Y NAND2X1_LOC_175/Y 0.51fF
C26778 NAND2X1_LOC_9/Y NOR2X1_LOC_520/A 0.04fF
C26779 NAND2X1_LOC_149/Y INVX1_LOC_49/A 0.14fF
C26780 NAND2X1_LOC_714/B INVX1_LOC_209/Y 0.00fF
C26781 NAND2X1_LOC_832/Y INVX1_LOC_12/A 0.01fF
C26782 INVX1_LOC_77/Y INVX1_LOC_118/A 0.07fF
C26783 NOR2X1_LOC_825/Y NAND2X1_LOC_848/Y 0.00fF
C26784 INVX1_LOC_136/A NOR2X1_LOC_530/Y 0.01fF
C26785 INVX1_LOC_55/Y INVX1_LOC_4/A 0.07fF
C26786 INVX1_LOC_35/A INVX1_LOC_143/A 0.07fF
C26787 INVX1_LOC_89/A INVX1_LOC_90/Y 0.01fF
C26788 INVX1_LOC_172/Y INVX1_LOC_23/A 0.03fF
C26789 INVX1_LOC_25/Y INVX1_LOC_29/Y 0.02fF
C26790 NOR2X1_LOC_368/A NOR2X1_LOC_76/B 0.03fF
C26791 INVX1_LOC_93/A NOR2X1_LOC_309/Y 0.10fF
C26792 NOR2X1_LOC_9/Y NOR2X1_LOC_641/a_36_216# 0.00fF
C26793 NOR2X1_LOC_590/A NOR2X1_LOC_703/B 0.03fF
C26794 INVX1_LOC_50/A NOR2X1_LOC_690/Y 0.09fF
C26795 NAND2X1_LOC_787/A NAND2X1_LOC_860/Y 0.01fF
C26796 INVX1_LOC_58/A NOR2X1_LOC_632/Y 0.03fF
C26797 INVX1_LOC_103/A NOR2X1_LOC_433/A 0.22fF
C26798 INVX1_LOC_35/A INVX1_LOC_68/Y 0.27fF
C26799 NAND2X1_LOC_348/A INVX1_LOC_15/A 0.08fF
C26800 NOR2X1_LOC_82/A INVX1_LOC_314/Y 0.02fF
C26801 INVX1_LOC_48/Y NOR2X1_LOC_121/Y 0.03fF
C26802 NAND2X1_LOC_656/Y NOR2X1_LOC_383/B 0.03fF
C26803 INVX1_LOC_298/Y INVX1_LOC_313/Y 0.05fF
C26804 NOR2X1_LOC_769/A INVX1_LOC_30/A 0.17fF
C26805 NOR2X1_LOC_607/Y INVX1_LOC_161/Y 0.07fF
C26806 NOR2X1_LOC_347/a_36_216# NAND2X1_LOC_206/Y 0.01fF
C26807 NOR2X1_LOC_730/Y INVX1_LOC_53/A 0.11fF
C26808 INVX1_LOC_1/A INVX1_LOC_294/Y 0.02fF
C26809 INVX1_LOC_222/A INVX1_LOC_32/A 0.10fF
C26810 INVX1_LOC_20/A NAND2X1_LOC_489/Y 0.07fF
C26811 NOR2X1_LOC_361/B INVX1_LOC_162/A 0.10fF
C26812 INVX1_LOC_21/A INVX1_LOC_214/A 0.12fF
C26813 INVX1_LOC_132/Y NOR2X1_LOC_383/B 0.03fF
C26814 NOR2X1_LOC_653/a_36_216# INVX1_LOC_285/A 0.01fF
C26815 INVX1_LOC_13/A INVX1_LOC_64/A 0.10fF
C26816 INVX1_LOC_2/A NAND2X1_LOC_149/Y 0.09fF
C26817 INVX1_LOC_21/A NOR2X1_LOC_667/A 0.43fF
C26818 NOR2X1_LOC_831/B NOR2X1_LOC_536/A 0.07fF
C26819 NAND2X1_LOC_849/B NOR2X1_LOC_88/Y 0.71fF
C26820 NOR2X1_LOC_756/Y INVX1_LOC_23/Y 0.03fF
C26821 INVX1_LOC_312/Y NOR2X1_LOC_512/Y 0.02fF
C26822 INVX1_LOC_21/A INVX1_LOC_248/A 0.09fF
C26823 NOR2X1_LOC_155/A NOR2X1_LOC_331/B 0.07fF
C26824 INVX1_LOC_307/A INVX1_LOC_9/A 0.07fF
C26825 NOR2X1_LOC_88/Y INVX1_LOC_38/A 0.03fF
C26826 NOR2X1_LOC_361/B NOR2X1_LOC_315/Y 0.10fF
C26827 INVX1_LOC_230/Y NOR2X1_LOC_672/Y 0.24fF
C26828 NAND2X1_LOC_807/Y NAND2X1_LOC_286/B 0.15fF
C26829 NOR2X1_LOC_32/B INVX1_LOC_219/A 0.03fF
C26830 INVX1_LOC_292/A NOR2X1_LOC_593/Y 0.07fF
C26831 INVX1_LOC_103/A NOR2X1_LOC_52/B 0.17fF
C26832 INVX1_LOC_9/A NOR2X1_LOC_445/B 0.07fF
C26833 NAND2X1_LOC_62/a_36_24# INVX1_LOC_92/A 0.00fF
C26834 INVX1_LOC_85/Y INVX1_LOC_23/A 0.06fF
C26835 INVX1_LOC_36/A NOR2X1_LOC_303/Y 0.03fF
C26836 NAND2X1_LOC_787/A NAND2X1_LOC_861/Y 0.10fF
C26837 INVX1_LOC_30/A NOR2X1_LOC_152/Y 0.10fF
C26838 NAND2X1_LOC_559/Y NAND2X1_LOC_733/B 0.18fF
C26839 NOR2X1_LOC_420/Y INVX1_LOC_30/Y 0.01fF
C26840 INVX1_LOC_35/A NOR2X1_LOC_130/A 17.88fF
C26841 NOR2X1_LOC_216/B NOR2X1_LOC_656/Y 0.05fF
C26842 NOR2X1_LOC_798/A NOR2X1_LOC_748/Y 0.01fF
C26843 NOR2X1_LOC_164/Y INVX1_LOC_102/A 0.02fF
C26844 NOR2X1_LOC_261/Y INVX1_LOC_90/A 0.15fF
C26845 NAND2X1_LOC_584/a_36_24# INVX1_LOC_11/A 0.01fF
C26846 NOR2X1_LOC_772/B NOR2X1_LOC_468/a_36_216# 0.00fF
C26847 INVX1_LOC_27/A INVX1_LOC_1/Y 0.07fF
C26848 NOR2X1_LOC_591/Y INVX1_LOC_161/Y 0.02fF
C26849 INVX1_LOC_144/A NOR2X1_LOC_449/A 0.08fF
C26850 NAND2X1_LOC_53/Y NAND2X1_LOC_629/Y 0.00fF
C26851 NAND2X1_LOC_849/B INVX1_LOC_84/A 0.47fF
C26852 INVX1_LOC_266/A NOR2X1_LOC_220/A 0.10fF
C26853 INVX1_LOC_269/A NOR2X1_LOC_616/Y 0.01fF
C26854 INVX1_LOC_14/A INVX1_LOC_256/Y 0.07fF
C26855 NAND2X1_LOC_35/Y INVX1_LOC_135/A 0.10fF
C26856 NOR2X1_LOC_453/Y NOR2X1_LOC_223/a_36_216# -0.02fF
C26857 INVX1_LOC_84/A INVX1_LOC_38/A 0.12fF
C26858 INVX1_LOC_303/A NAND2X1_LOC_689/a_36_24# 0.01fF
C26859 INVX1_LOC_31/A NOR2X1_LOC_516/Y 0.02fF
C26860 INVX1_LOC_278/A INVX1_LOC_90/A 0.16fF
C26861 NAND2X1_LOC_555/Y INVX1_LOC_82/A 0.14fF
C26862 INVX1_LOC_105/A INVX1_LOC_18/A 0.01fF
C26863 INVX1_LOC_269/A NAND2X1_LOC_563/A 0.15fF
C26864 NOR2X1_LOC_614/Y INVX1_LOC_24/Y 0.13fF
C26865 NOR2X1_LOC_296/a_36_216# NOR2X1_LOC_78/B 0.02fF
C26866 NOR2X1_LOC_831/B NAND2X1_LOC_93/B 0.07fF
C26867 NOR2X1_LOC_754/A NOR2X1_LOC_253/Y 0.01fF
C26868 NAND2X1_LOC_725/Y NOR2X1_LOC_380/Y 0.03fF
C26869 INVX1_LOC_255/Y INVX1_LOC_239/A 0.01fF
C26870 NOR2X1_LOC_9/Y INVX1_LOC_116/Y 0.02fF
C26871 NOR2X1_LOC_96/Y INVX1_LOC_84/A 0.18fF
C26872 INVX1_LOC_64/A INVX1_LOC_207/Y 0.25fF
C26873 NOR2X1_LOC_561/Y NAND2X1_LOC_474/Y 0.01fF
C26874 INVX1_LOC_102/A INVX1_LOC_46/A 0.08fF
C26875 INVX1_LOC_64/A INVX1_LOC_55/Y 0.07fF
C26876 INVX1_LOC_75/A INVX1_LOC_29/Y 0.07fF
C26877 INVX1_LOC_235/Y NAND2X1_LOC_462/B 0.31fF
C26878 INVX1_LOC_147/Y INVX1_LOC_32/A 0.29fF
C26879 NOR2X1_LOC_557/A INVX1_LOC_87/A 0.12fF
C26880 NOR2X1_LOC_124/A NOR2X1_LOC_38/B 0.00fF
C26881 NOR2X1_LOC_208/Y NOR2X1_LOC_303/Y 0.03fF
C26882 NOR2X1_LOC_468/Y INVX1_LOC_30/Y 0.21fF
C26883 INVX1_LOC_72/A INVX1_LOC_8/A 0.01fF
C26884 NOR2X1_LOC_311/a_36_216# NAND2X1_LOC_175/Y 0.00fF
C26885 NOR2X1_LOC_527/Y INVX1_LOC_57/A 0.01fF
C26886 NOR2X1_LOC_436/a_36_216# NOR2X1_LOC_174/B 0.00fF
C26887 NOR2X1_LOC_817/a_36_216# NOR2X1_LOC_516/B 0.00fF
C26888 INVX1_LOC_25/A NOR2X1_LOC_74/A 0.07fF
C26889 INVX1_LOC_32/A INVX1_LOC_20/A 0.10fF
C26890 NAND2X1_LOC_308/Y NAND2X1_LOC_856/A 0.24fF
C26891 INVX1_LOC_171/A INVX1_LOC_171/Y 0.05fF
C26892 NOR2X1_LOC_15/Y INVX1_LOC_279/A 0.07fF
C26893 NOR2X1_LOC_272/Y INVX1_LOC_89/A 0.00fF
C26894 NAND2X1_LOC_733/A NOR2X1_LOC_822/Y 0.04fF
C26895 INVX1_LOC_284/Y NAND2X1_LOC_839/A 0.12fF
C26896 INVX1_LOC_42/Y NOR2X1_LOC_678/A 0.03fF
C26897 NAND2X1_LOC_848/Y INVX1_LOC_84/A 0.03fF
C26898 D_INPUT_0 INVX1_LOC_48/Y 0.77fF
C26899 NOR2X1_LOC_357/Y INVX1_LOC_4/A 0.10fF
C26900 INVX1_LOC_25/A NOR2X1_LOC_9/Y 0.69fF
C26901 NOR2X1_LOC_837/A INVX1_LOC_57/A 0.02fF
C26902 INVX1_LOC_35/A NOR2X1_LOC_112/B 0.03fF
C26903 INVX1_LOC_36/A INVX1_LOC_54/Y 0.29fF
C26904 INVX1_LOC_34/A NOR2X1_LOC_238/Y 0.00fF
C26905 INVX1_LOC_136/A NOR2X1_LOC_709/A 0.10fF
C26906 INVX1_LOC_12/A INVX1_LOC_9/A 0.07fF
C26907 NAND2X1_LOC_639/A NAND2X1_LOC_430/B 0.05fF
C26908 NOR2X1_LOC_553/Y NOR2X1_LOC_553/a_36_216# 0.00fF
C26909 INVX1_LOC_62/Y NOR2X1_LOC_6/B 0.36fF
C26910 NOR2X1_LOC_216/B INVX1_LOC_63/A 0.12fF
C26911 NOR2X1_LOC_134/Y INVX1_LOC_16/A 0.06fF
C26912 NAND2X1_LOC_860/A INVX1_LOC_6/A 0.16fF
C26913 INVX1_LOC_129/Y INVX1_LOC_251/A 0.03fF
C26914 NOR2X1_LOC_78/B INVX1_LOC_223/A 0.03fF
C26915 NAND2X1_LOC_213/A INVX1_LOC_89/A 0.38fF
C26916 NAND2X1_LOC_57/a_36_24# NAND2X1_LOC_338/B 0.00fF
C26917 INVX1_LOC_278/Y NAND2X1_LOC_185/a_36_24# 0.00fF
C26918 NAND2X1_LOC_642/Y NOR2X1_LOC_39/Y 0.00fF
C26919 INVX1_LOC_174/A GATE_662 0.17fF
C26920 NOR2X1_LOC_160/B NAND2X1_LOC_41/Y 0.01fF
C26921 NAND2X1_LOC_483/Y NAND2X1_LOC_632/B -0.00fF
C26922 NAND2X1_LOC_175/Y INVX1_LOC_20/A 0.16fF
C26923 NOR2X1_LOC_831/Y NOR2X1_LOC_743/Y 0.07fF
C26924 NOR2X1_LOC_78/A NAND2X1_LOC_215/A 0.17fF
C26925 NOR2X1_LOC_772/B NOR2X1_LOC_292/Y 0.02fF
C26926 NOR2X1_LOC_565/A NOR2X1_LOC_500/Y 0.03fF
C26927 NAND2X1_LOC_860/Y INVX1_LOC_30/A 0.05fF
C26928 INVX1_LOC_135/A NAND2X1_LOC_377/a_36_24# 0.00fF
C26929 NAND2X1_LOC_112/Y NOR2X1_LOC_441/Y 1.68fF
C26930 NOR2X1_LOC_445/Y INVX1_LOC_33/A 0.04fF
C26931 NOR2X1_LOC_391/A NOR2X1_LOC_160/B 0.18fF
C26932 NOR2X1_LOC_15/Y NOR2X1_LOC_166/a_36_216# 0.00fF
C26933 NAND2X1_LOC_860/A NOR2X1_LOC_10/a_36_216# 0.00fF
C26934 INVX1_LOC_27/A NOR2X1_LOC_742/A 0.59fF
C26935 INVX1_LOC_2/A NOR2X1_LOC_744/Y 0.01fF
C26936 NOR2X1_LOC_264/Y NOR2X1_LOC_716/B 0.21fF
C26937 INVX1_LOC_30/A NAND2X1_LOC_859/B 0.01fF
C26938 NOR2X1_LOC_718/B NOR2X1_LOC_550/B 0.10fF
C26939 INVX1_LOC_11/A INVX1_LOC_120/A 0.03fF
C26940 INVX1_LOC_38/A INVX1_LOC_15/A 0.21fF
C26941 INVX1_LOC_21/A NAND2X1_LOC_51/B 0.01fF
C26942 INVX1_LOC_163/A NAND2X1_LOC_462/a_36_24# 0.00fF
C26943 NOR2X1_LOC_208/Y NOR2X1_LOC_353/Y 0.01fF
C26944 D_INPUT_7 INVX1_LOC_22/A 0.01fF
C26945 INVX1_LOC_51/Y INVX1_LOC_50/Y 0.05fF
C26946 NOR2X1_LOC_15/Y INVX1_LOC_182/Y 0.03fF
C26947 INVX1_LOC_290/Y INVX1_LOC_92/A 0.09fF
C26948 INVX1_LOC_21/A INVX1_LOC_311/A 0.12fF
C26949 INVX1_LOC_223/Y NOR2X1_LOC_552/Y 0.02fF
C26950 NAND2X1_LOC_115/a_36_24# INVX1_LOC_104/A 0.06fF
C26951 NAND2X1_LOC_175/Y NOR2X1_LOC_765/Y 0.05fF
C26952 NOR2X1_LOC_186/Y INVX1_LOC_286/A 0.04fF
C26953 NAND2X1_LOC_218/B NAND2X1_LOC_672/B 0.01fF
C26954 NOR2X1_LOC_718/B INVX1_LOC_249/Y 0.11fF
C26955 NOR2X1_LOC_857/A NOR2X1_LOC_748/A 0.21fF
C26956 INVX1_LOC_24/A NOR2X1_LOC_121/A 1.32fF
C26957 INVX1_LOC_77/A NOR2X1_LOC_566/Y 0.04fF
C26958 INVX1_LOC_251/Y INVX1_LOC_41/A 0.03fF
C26959 NOR2X1_LOC_382/Y NOR2X1_LOC_332/A 0.03fF
C26960 INVX1_LOC_46/A INVX1_LOC_296/Y 0.05fF
C26961 INVX1_LOC_1/A NOR2X1_LOC_74/A 0.29fF
C26962 INVX1_LOC_35/A NOR2X1_LOC_209/A 0.07fF
C26963 NOR2X1_LOC_454/Y NAND2X1_LOC_841/a_36_24# 0.00fF
C26964 NOR2X1_LOC_144/Y INVX1_LOC_96/Y 0.01fF
C26965 NOR2X1_LOC_239/a_36_216# NOR2X1_LOC_99/B 0.01fF
C26966 INVX1_LOC_58/A NAND2X1_LOC_39/Y 0.03fF
C26967 NOR2X1_LOC_15/Y NAND2X1_LOC_858/B 0.07fF
C26968 NOR2X1_LOC_447/Y NOR2X1_LOC_328/Y 0.01fF
C26969 INVX1_LOC_30/A NAND2X1_LOC_861/Y 1.47fF
C26970 INVX1_LOC_8/A NOR2X1_LOC_537/Y 0.07fF
C26971 NOR2X1_LOC_483/B INVX1_LOC_311/Y 0.01fF
C26972 NOR2X1_LOC_134/Y INVX1_LOC_28/A 0.02fF
C26973 NAND2X1_LOC_338/B INVX1_LOC_8/A 0.36fF
C26974 INVX1_LOC_54/Y NOR2X1_LOC_309/Y 0.05fF
C26975 INVX1_LOC_278/A NOR2X1_LOC_92/a_36_216# 0.00fF
C26976 NAND2X1_LOC_364/A INVX1_LOC_150/A 0.02fF
C26977 INVX1_LOC_1/A NOR2X1_LOC_9/Y 0.18fF
C26978 INVX1_LOC_27/A NOR2X1_LOC_318/B 0.07fF
C26979 NOR2X1_LOC_205/a_36_216# NOR2X1_LOC_388/Y 0.00fF
C26980 INVX1_LOC_49/A INVX1_LOC_16/A 0.03fF
C26981 NAND2X1_LOC_206/B NAND2X1_LOC_206/Y 0.02fF
C26982 INVX1_LOC_41/A NOR2X1_LOC_614/Y 0.01fF
C26983 NAND2X1_LOC_785/Y NOR2X1_LOC_667/A 0.00fF
C26984 NOR2X1_LOC_91/Y NOR2X1_LOC_71/Y 0.00fF
C26985 INVX1_LOC_286/Y NOR2X1_LOC_329/B 0.17fF
C26986 INVX1_LOC_64/A NOR2X1_LOC_357/Y 0.13fF
C26987 NAND2X1_LOC_343/a_36_24# INVX1_LOC_49/A 0.00fF
C26988 INVX1_LOC_89/A NAND2X1_LOC_364/A 0.08fF
C26989 NOR2X1_LOC_569/Y NOR2X1_LOC_550/B 0.01fF
C26990 INVX1_LOC_27/A INVX1_LOC_93/Y 0.10fF
C26991 NOR2X1_LOC_456/Y NAND2X1_LOC_472/Y 1.11fF
C26992 NOR2X1_LOC_794/B NOR2X1_LOC_74/A 0.00fF
C26993 NOR2X1_LOC_612/Y INVX1_LOC_26/A 0.01fF
C26994 NOR2X1_LOC_92/Y NOR2X1_LOC_45/B 0.78fF
C26995 INVX1_LOC_247/Y INVX1_LOC_313/Y 0.04fF
C26996 INVX1_LOC_21/A INVX1_LOC_304/A 0.14fF
C26997 INVX1_LOC_268/A INVX1_LOC_34/A 0.03fF
C26998 NOR2X1_LOC_644/Y NOR2X1_LOC_655/B 0.04fF
C26999 INVX1_LOC_104/A NOR2X1_LOC_388/a_36_216# 0.00fF
C27000 INVX1_LOC_90/A NOR2X1_LOC_168/Y 0.03fF
C27001 NAND2X1_LOC_205/A NOR2X1_LOC_271/Y 0.02fF
C27002 NOR2X1_LOC_331/B NOR2X1_LOC_125/Y 0.03fF
C27003 D_INPUT_0 NOR2X1_LOC_350/A 0.04fF
C27004 NOR2X1_LOC_703/B NOR2X1_LOC_703/A 0.49fF
C27005 NOR2X1_LOC_155/A NOR2X1_LOC_449/A 0.01fF
C27006 NAND2X1_LOC_499/a_36_24# NAND2X1_LOC_254/Y 0.00fF
C27007 INVX1_LOC_35/A NOR2X1_LOC_115/a_36_216# 0.00fF
C27008 INVX1_LOC_299/A INVX1_LOC_65/A 0.05fF
C27009 NOR2X1_LOC_468/Y NOR2X1_LOC_124/A 0.02fF
C27010 NOR2X1_LOC_667/A INVX1_LOC_248/A 0.13fF
C27011 NAND2X1_LOC_474/Y INVX1_LOC_76/A 0.10fF
C27012 INVX1_LOC_243/Y NAND2X1_LOC_638/a_36_24# 0.00fF
C27013 NOR2X1_LOC_829/A NAND2X1_LOC_810/B 0.00fF
C27014 INVX1_LOC_136/A NAND2X1_LOC_863/A 0.01fF
C27015 NAND2X1_LOC_35/Y NOR2X1_LOC_813/Y 0.02fF
C27016 INVX1_LOC_162/A NAND2X1_LOC_573/A 0.01fF
C27017 NOR2X1_LOC_596/A NOR2X1_LOC_156/A 0.08fF
C27018 INVX1_LOC_27/A INVX1_LOC_139/A 0.01fF
C27019 INVX1_LOC_17/A NOR2X1_LOC_595/Y 0.01fF
C27020 INVX1_LOC_206/A INVX1_LOC_1/Y 0.13fF
C27021 INVX1_LOC_222/Y VDD 0.42fF
C27022 NAND2X1_LOC_803/B INVX1_LOC_91/A 0.02fF
C27023 NOR2X1_LOC_412/a_36_216# D_INPUT_0 0.00fF
C27024 INVX1_LOC_2/A INVX1_LOC_16/A 0.17fF
C27025 NAND2X1_LOC_190/Y INVX1_LOC_188/Y 0.01fF
C27026 NOR2X1_LOC_590/A NOR2X1_LOC_114/A 0.01fF
C27027 NOR2X1_LOC_615/Y INVX1_LOC_91/A 0.06fF
C27028 NOR2X1_LOC_500/Y INVX1_LOC_179/Y 0.02fF
C27029 NAND2X1_LOC_33/Y NAND2X1_LOC_461/a_36_24# 0.00fF
C27030 INVX1_LOC_181/Y INVX1_LOC_73/A 0.03fF
C27031 NOR2X1_LOC_226/A INVX1_LOC_16/A 0.07fF
C27032 NOR2X1_LOC_582/Y NAND2X1_LOC_51/B 0.02fF
C27033 INVX1_LOC_33/A NOR2X1_LOC_542/Y 0.54fF
C27034 NOR2X1_LOC_223/B INVX1_LOC_38/A 0.04fF
C27035 NOR2X1_LOC_824/A NAND2X1_LOC_721/A 0.07fF
C27036 INVX1_LOC_26/A NOR2X1_LOC_673/A 0.15fF
C27037 NAND2X1_LOC_715/B NOR2X1_LOC_331/B 0.00fF
C27038 NOR2X1_LOC_590/A INVX1_LOC_91/A 0.34fF
C27039 INVX1_LOC_23/A NOR2X1_LOC_461/A 0.05fF
C27040 INVX1_LOC_49/A INVX1_LOC_28/A 2.40fF
C27041 NAND2X1_LOC_200/B INVX1_LOC_1/Y 0.12fF
C27042 NOR2X1_LOC_464/B VDD 0.02fF
C27043 NOR2X1_LOC_111/Y NOR2X1_LOC_577/Y 0.04fF
C27044 INVX1_LOC_249/A NOR2X1_LOC_742/A 0.01fF
C27045 NAND2X1_LOC_9/Y INVX1_LOC_70/A 0.17fF
C27046 NOR2X1_LOC_441/Y NOR2X1_LOC_78/A 0.01fF
C27047 NAND2X1_LOC_361/Y INVX1_LOC_148/A 0.01fF
C27048 D_INPUT_0 NOR2X1_LOC_84/Y 0.15fF
C27049 NAND2X1_LOC_774/a_36_24# INVX1_LOC_46/A 0.01fF
C27050 INVX1_LOC_233/A INVX1_LOC_70/A 0.01fF
C27051 NOR2X1_LOC_186/Y NOR2X1_LOC_602/B 0.01fF
C27052 NAND2X1_LOC_53/Y INVX1_LOC_76/A 0.23fF
C27053 NOR2X1_LOC_406/a_36_216# INVX1_LOC_185/A 0.00fF
C27054 NAND2X1_LOC_192/B VDD 0.01fF
C27055 D_INPUT_0 INVX1_LOC_216/A 0.05fF
C27056 NOR2X1_LOC_596/A NAND2X1_LOC_328/a_36_24# 0.02fF
C27057 INVX1_LOC_284/Y NOR2X1_LOC_823/Y 0.08fF
C27058 INVX1_LOC_35/A NOR2X1_LOC_197/B 0.03fF
C27059 NOR2X1_LOC_186/Y INVX1_LOC_54/A 0.07fF
C27060 INVX1_LOC_64/A INVX1_LOC_260/A 0.00fF
C27061 NOR2X1_LOC_318/A INVX1_LOC_19/A 0.03fF
C27062 INPUT_3 INVX1_LOC_20/A 0.09fF
C27063 NOR2X1_LOC_687/Y NOR2X1_LOC_730/A 0.02fF
C27064 NOR2X1_LOC_15/Y NOR2X1_LOC_98/B 0.03fF
C27065 INVX1_LOC_226/Y INVX1_LOC_7/A 0.09fF
C27066 NAND2X1_LOC_573/Y NOR2X1_LOC_602/B 0.02fF
C27067 NOR2X1_LOC_667/A NAND2X1_LOC_804/a_36_24# 0.00fF
C27068 NAND2X1_LOC_577/A NAND2X1_LOC_659/B 0.39fF
C27069 NOR2X1_LOC_763/Y NAND2X1_LOC_451/a_36_24# 0.01fF
C27070 INVX1_LOC_32/A INVX1_LOC_4/A 0.22fF
C27071 NAND2X1_LOC_573/Y INVX1_LOC_54/A 0.07fF
C27072 NOR2X1_LOC_400/B INVX1_LOC_29/A 0.07fF
C27073 INVX1_LOC_23/A NAND2X1_LOC_782/B 0.04fF
C27074 INVX1_LOC_2/A INVX1_LOC_28/A 0.41fF
C27075 INVX1_LOC_98/Y NAND2X1_LOC_850/A 0.05fF
C27076 NOR2X1_LOC_45/B NAND2X1_LOC_837/Y 0.07fF
C27077 NAND2X1_LOC_553/A INVX1_LOC_123/Y 0.00fF
C27078 NOR2X1_LOC_355/A NAND2X1_LOC_349/B 0.20fF
C27079 NOR2X1_LOC_160/B INVX1_LOC_122/A 0.09fF
C27080 NOR2X1_LOC_226/A INVX1_LOC_28/A 0.27fF
C27081 NAND2X1_LOC_577/A VDD 0.05fF
C27082 NOR2X1_LOC_561/Y INVX1_LOC_10/A 0.10fF
C27083 NOR2X1_LOC_565/a_36_216# INVX1_LOC_104/A 0.00fF
C27084 NOR2X1_LOC_552/A INVX1_LOC_94/A 0.02fF
C27085 INVX1_LOC_279/A NAND2X1_LOC_130/a_36_24# 0.00fF
C27086 NOR2X1_LOC_30/Y D_INPUT_5 0.02fF
C27087 INVX1_LOC_16/A NAND2X1_LOC_648/A 0.03fF
C27088 NOR2X1_LOC_454/Y INVX1_LOC_92/A 0.08fF
C27089 NOR2X1_LOC_710/A INVX1_LOC_117/A 0.00fF
C27090 INVX1_LOC_16/A INPUT_1 0.48fF
C27091 INVX1_LOC_223/A INVX1_LOC_46/A 0.03fF
C27092 INVX1_LOC_89/A NOR2X1_LOC_86/A 0.16fF
C27093 INVX1_LOC_19/A NOR2X1_LOC_678/A 0.03fF
C27094 NAND2X1_LOC_352/B NOR2X1_LOC_536/A 0.03fF
C27095 INVX1_LOC_48/Y INVX1_LOC_46/Y 0.64fF
C27096 NOR2X1_LOC_561/Y NOR2X1_LOC_504/a_36_216# 0.01fF
C27097 INVX1_LOC_186/A NOR2X1_LOC_551/B 0.03fF
C27098 INVX1_LOC_94/Y INVX1_LOC_4/Y 0.32fF
C27099 NOR2X1_LOC_392/B INVX1_LOC_123/A 0.02fF
C27100 NOR2X1_LOC_772/A INVX1_LOC_1/Y 0.01fF
C27101 INVX1_LOC_24/Y NOR2X1_LOC_862/B 0.01fF
C27102 NOR2X1_LOC_723/a_36_216# INVX1_LOC_139/Y 0.00fF
C27103 NOR2X1_LOC_113/A NAND2X1_LOC_283/a_36_24# 0.00fF
C27104 NOR2X1_LOC_111/Y INVX1_LOC_22/A 0.05fF
C27105 NAND2X1_LOC_354/B INVX1_LOC_91/A 0.02fF
C27106 NOR2X1_LOC_773/Y NOR2X1_LOC_527/a_36_216# 0.01fF
C27107 NOR2X1_LOC_789/B INVX1_LOC_3/A 0.03fF
C27108 INVX1_LOC_93/A INVX1_LOC_63/A 0.00fF
C27109 INVX1_LOC_213/Y INVX1_LOC_186/A 0.03fF
C27110 NOR2X1_LOC_45/Y INVX1_LOC_54/A 0.02fF
C27111 NAND2X1_LOC_656/A VDD 0.79fF
C27112 INVX1_LOC_53/A INVX1_LOC_290/Y 0.01fF
C27113 NOR2X1_LOC_744/a_36_216# NOR2X1_LOC_111/A 0.00fF
C27114 INVX1_LOC_249/A INVX1_LOC_139/A 0.15fF
C27115 INVX1_LOC_49/A NOR2X1_LOC_35/Y 0.28fF
C27116 INVX1_LOC_41/A INVX1_LOC_247/A 0.00fF
C27117 NOR2X1_LOC_45/B NAND2X1_LOC_477/A 0.28fF
C27118 VDD NOR2X1_LOC_484/Y -0.00fF
C27119 INVX1_LOC_34/A INVX1_LOC_95/Y 0.07fF
C27120 INVX1_LOC_206/A NOR2X1_LOC_318/B 0.03fF
C27121 INVX1_LOC_225/A INVX1_LOC_95/A 0.05fF
C27122 D_GATE_741 NAND2X1_LOC_425/Y 0.02fF
C27123 INVX1_LOC_256/A NOR2X1_LOC_831/B 0.20fF
C27124 NOR2X1_LOC_458/B INVX1_LOC_206/Y 0.03fF
C27125 NOR2X1_LOC_759/Y NAND2X1_LOC_472/Y 0.02fF
C27126 NAND2X1_LOC_146/a_36_24# NOR2X1_LOC_148/Y 0.00fF
C27127 NOR2X1_LOC_655/B NOR2X1_LOC_78/A 0.05fF
C27128 NOR2X1_LOC_168/Y INVX1_LOC_38/A 0.03fF
C27129 NOR2X1_LOC_493/B NOR2X1_LOC_405/A 0.25fF
C27130 NOR2X1_LOC_465/a_36_216# INVX1_LOC_32/A 0.01fF
C27131 NOR2X1_LOC_186/Y NAND2X1_LOC_807/B 0.01fF
C27132 NOR2X1_LOC_220/A INVX1_LOC_96/A 0.01fF
C27133 NOR2X1_LOC_577/Y NAND2X1_LOC_687/A 0.04fF
C27134 INVX1_LOC_136/A NOR2X1_LOC_489/A 0.21fF
C27135 INVX1_LOC_30/A INVX1_LOC_291/A 0.07fF
C27136 INVX1_LOC_28/A INPUT_1 0.10fF
C27137 NOR2X1_LOC_355/A INVX1_LOC_75/A 0.05fF
C27138 INVX1_LOC_64/A INVX1_LOC_32/A 0.07fF
C27139 NOR2X1_LOC_550/B NAND2X1_LOC_472/Y 0.10fF
C27140 INVX1_LOC_36/A NOR2X1_LOC_78/Y 0.06fF
C27141 NAND2X1_LOC_454/Y INVX1_LOC_23/A 0.08fF
C27142 NOR2X1_LOC_577/Y NOR2X1_LOC_363/Y 0.00fF
C27143 NAND2X1_LOC_573/a_36_24# NOR2X1_LOC_536/A 0.00fF
C27144 NOR2X1_LOC_690/A INVX1_LOC_37/A 0.00fF
C27145 NOR2X1_LOC_251/Y NOR2X1_LOC_318/B -0.01fF
C27146 INVX1_LOC_196/A NOR2X1_LOC_324/A 0.49fF
C27147 INVX1_LOC_45/A NOR2X1_LOC_634/A 0.02fF
C27148 INVX1_LOC_64/A NOR2X1_LOC_623/B 0.00fF
C27149 NAND2X1_LOC_860/A NOR2X1_LOC_80/Y 0.04fF
C27150 NAND2X1_LOC_740/B NAND2X1_LOC_308/B 0.01fF
C27151 INVX1_LOC_64/A NOR2X1_LOC_329/Y 0.04fF
C27152 NOR2X1_LOC_169/B NOR2X1_LOC_445/B 0.01fF
C27153 NAND2X1_LOC_67/Y INVX1_LOC_12/A 0.07fF
C27154 INVX1_LOC_104/A NOR2X1_LOC_139/a_36_216# 0.00fF
C27155 NOR2X1_LOC_84/Y NOR2X1_LOC_266/B 0.01fF
C27156 NOR2X1_LOC_316/Y INVX1_LOC_46/A 0.01fF
C27157 NOR2X1_LOC_423/Y VDD 0.33fF
C27158 INVX1_LOC_21/A INVX1_LOC_19/Y 0.01fF
C27159 NOR2X1_LOC_412/a_36_216# NAND2X1_LOC_848/A 0.02fF
C27160 INVX1_LOC_141/Y INVX1_LOC_250/Y 0.04fF
C27161 NAND2X1_LOC_21/Y INVX1_LOC_38/A 0.02fF
C27162 INVX1_LOC_45/A NAND2X1_LOC_606/a_36_24# 0.00fF
C27163 NAND2X1_LOC_573/Y NOR2X1_LOC_48/B 0.22fF
C27164 NOR2X1_LOC_234/Y NOR2X1_LOC_813/Y 0.01fF
C27165 NOR2X1_LOC_562/A NOR2X1_LOC_352/Y 0.03fF
C27166 INVX1_LOC_64/A NAND2X1_LOC_175/Y 0.07fF
C27167 NOR2X1_LOC_219/Y NAND2X1_LOC_212/Y 0.00fF
C27168 NOR2X1_LOC_203/a_36_216# NOR2X1_LOC_334/Y 0.01fF
C27169 INVX1_LOC_57/A NOR2X1_LOC_654/A 0.14fF
C27170 NAND2X1_LOC_358/Y NOR2X1_LOC_78/A 0.05fF
C27171 NOR2X1_LOC_533/Y NOR2X1_LOC_89/A 0.03fF
C27172 INVX1_LOC_41/A NOR2X1_LOC_499/B 0.09fF
C27173 NAND2X1_LOC_149/Y INVX1_LOC_257/A 0.02fF
C27174 INVX1_LOC_2/Y NOR2X1_LOC_346/B 0.07fF
C27175 NOR2X1_LOC_356/A NOR2X1_LOC_188/A 0.11fF
C27176 NAND2X1_LOC_357/B NOR2X1_LOC_536/A 0.14fF
C27177 NOR2X1_LOC_470/B NOR2X1_LOC_477/B 0.18fF
C27178 NOR2X1_LOC_763/Y INVX1_LOC_91/A 0.01fF
C27179 NOR2X1_LOC_222/Y VDD 0.43fF
C27180 NAND2X1_LOC_640/Y INVX1_LOC_54/A 0.00fF
C27181 NOR2X1_LOC_356/A NOR2X1_LOC_548/B 0.01fF
C27182 INVX1_LOC_226/Y INVX1_LOC_76/A 0.10fF
C27183 INVX1_LOC_77/A INVX1_LOC_92/A 0.21fF
C27184 INVX1_LOC_269/A NOR2X1_LOC_554/A 0.01fF
C27185 NOR2X1_LOC_78/A NOR2X1_LOC_99/B 0.09fF
C27186 NOR2X1_LOC_383/B NOR2X1_LOC_717/A 0.11fF
C27187 INVX1_LOC_136/A INVX1_LOC_294/A 0.03fF
C27188 NAND2X1_LOC_21/Y NOR2X1_LOC_51/A 0.03fF
C27189 NAND2X1_LOC_564/B INVX1_LOC_20/A 0.10fF
C27190 NOR2X1_LOC_405/A INVX1_LOC_150/A 0.02fF
C27191 INVX1_LOC_225/A INVX1_LOC_54/A 0.03fF
C27192 NOR2X1_LOC_405/A NOR2X1_LOC_110/a_36_216# 0.00fF
C27193 INVX1_LOC_89/A NOR2X1_LOC_349/A 0.09fF
C27194 NAND2X1_LOC_563/A INVX1_LOC_12/Y 0.01fF
C27195 INVX1_LOC_41/A NOR2X1_LOC_676/Y 0.04fF
C27196 INVX1_LOC_17/A D_INPUT_5 0.01fF
C27197 NOR2X1_LOC_473/B NOR2X1_LOC_139/Y 0.06fF
C27198 INVX1_LOC_89/A NOR2X1_LOC_405/A 0.10fF
C27199 INVX1_LOC_41/A NOR2X1_LOC_862/B 0.24fF
C27200 INVX1_LOC_45/A INVX1_LOC_29/A 3.26fF
C27201 INVX1_LOC_299/A INVX1_LOC_4/Y 0.07fF
C27202 INVX1_LOC_305/A INVX1_LOC_19/A 0.07fF
C27203 NAND2X1_LOC_708/Y NOR2X1_LOC_696/Y 0.22fF
C27204 NOR2X1_LOC_188/A NOR2X1_LOC_74/A 2.52fF
C27205 NOR2X1_LOC_568/A INVX1_LOC_29/A 0.00fF
C27206 INVX1_LOC_10/A INVX1_LOC_76/A 4.82fF
C27207 INVX1_LOC_22/A INVX1_LOC_37/Y 0.01fF
C27208 NOR2X1_LOC_770/a_36_216# NAND2X1_LOC_93/B 0.00fF
C27209 VDD INVX1_LOC_220/Y 0.02fF
C27210 NAND2X1_LOC_508/A NOR2X1_LOC_349/A 0.05fF
C27211 NAND2X1_LOC_717/Y INVX1_LOC_118/A 0.05fF
C27212 NOR2X1_LOC_703/A INVX1_LOC_91/A 0.05fF
C27213 NOR2X1_LOC_188/A NOR2X1_LOC_9/Y 0.03fF
C27214 NOR2X1_LOC_399/a_36_216# NOR2X1_LOC_629/Y 0.00fF
C27215 NOR2X1_LOC_770/a_36_216# NAND2X1_LOC_425/Y 0.01fF
C27216 NOR2X1_LOC_548/B NOR2X1_LOC_9/Y 0.05fF
C27217 INVX1_LOC_138/Y NOR2X1_LOC_392/Y 0.01fF
C27218 NAND2X1_LOC_198/B NOR2X1_LOC_831/Y 0.47fF
C27219 INVX1_LOC_234/A NAND2X1_LOC_721/A 0.08fF
C27220 INPUT_5 INVX1_LOC_77/Y 0.34fF
C27221 INPUT_3 INVX1_LOC_4/A 0.10fF
C27222 INVX1_LOC_33/A INVX1_LOC_84/A 0.08fF
C27223 INVX1_LOC_89/A NOR2X1_LOC_857/A 0.08fF
C27224 NOR2X1_LOC_380/A VDD 0.33fF
C27225 INVX1_LOC_183/Y NAND2X1_LOC_650/B 0.01fF
C27226 NOR2X1_LOC_593/Y NOR2X1_LOC_631/A 0.14fF
C27227 NOR2X1_LOC_329/B NOR2X1_LOC_56/Y 0.98fF
C27228 INVX1_LOC_25/Y INVX1_LOC_127/A 0.01fF
C27229 INVX1_LOC_50/A NOR2X1_LOC_321/Y 0.10fF
C27230 NOR2X1_LOC_514/Y NOR2X1_LOC_649/B 0.03fF
C27231 INVX1_LOC_71/A INVX1_LOC_29/A 0.30fF
C27232 INVX1_LOC_73/A NOR2X1_LOC_675/A 0.05fF
C27233 INVX1_LOC_16/A INVX1_LOC_118/A 1.05fF
C27234 NOR2X1_LOC_361/B NAND2X1_LOC_99/A 0.10fF
C27235 NOR2X1_LOC_572/a_36_216# INVX1_LOC_280/A 0.01fF
C27236 NOR2X1_LOC_254/Y INVX1_LOC_63/A 0.06fF
C27237 INVX1_LOC_179/Y INVX1_LOC_307/A 0.02fF
C27238 NAND2X1_LOC_79/Y INVX1_LOC_284/A 0.11fF
C27239 NAND2X1_LOC_337/B NOR2X1_LOC_278/Y 0.07fF
C27240 NOR2X1_LOC_329/B NOR2X1_LOC_136/a_36_216# 0.01fF
C27241 NOR2X1_LOC_366/B NOR2X1_LOC_155/A 0.05fF
C27242 INVX1_LOC_121/A NOR2X1_LOC_378/Y 0.01fF
C27243 INVX1_LOC_49/A INVX1_LOC_109/A 0.01fF
C27244 NAND2X1_LOC_798/A NOR2X1_LOC_88/Y 0.02fF
C27245 NAND2X1_LOC_357/B NOR2X1_LOC_661/A 0.08fF
C27246 NOR2X1_LOC_329/B INVX1_LOC_146/Y 0.01fF
C27247 NOR2X1_LOC_454/Y INVX1_LOC_53/A 0.07fF
C27248 INVX1_LOC_95/Y INPUT_0 0.13fF
C27249 NOR2X1_LOC_329/B VDD 1.89fF
C27250 NAND2X1_LOC_369/a_36_24# INVX1_LOC_14/Y 0.00fF
C27251 NOR2X1_LOC_713/a_36_216# INVX1_LOC_91/A 0.00fF
C27252 INVX1_LOC_286/A NAND2X1_LOC_642/Y 0.19fF
C27253 D_GATE_579 INVX1_LOC_241/Y 0.05fF
C27254 INVX1_LOC_162/A NAND2X1_LOC_81/B 0.36fF
C27255 D_INPUT_4 VDD 0.75fF
C27256 INVX1_LOC_1/Y NOR2X1_LOC_216/B 0.54fF
C27257 NAND2X1_LOC_479/Y NOR2X1_LOC_155/A 0.01fF
C27258 INVX1_LOC_54/Y INVX1_LOC_63/A 0.00fF
C27259 INVX1_LOC_136/A NOR2X1_LOC_334/Y 0.10fF
C27260 NOR2X1_LOC_122/A NOR2X1_LOC_678/A 0.00fF
C27261 INVX1_LOC_72/A NOR2X1_LOC_158/a_36_216# 0.00fF
C27262 INVX1_LOC_298/Y INVX1_LOC_45/A 0.02fF
C27263 NOR2X1_LOC_848/Y NOR2X1_LOC_598/B 0.25fF
C27264 NOR2X1_LOC_315/Y NAND2X1_LOC_81/B 0.07fF
C27265 NAND2X1_LOC_9/Y NOR2X1_LOC_296/a_36_216# 0.00fF
C27266 INVX1_LOC_40/A INVX1_LOC_84/A 0.43fF
C27267 INVX1_LOC_225/A NAND2X1_LOC_807/B 0.89fF
C27268 NOR2X1_LOC_367/B INVX1_LOC_12/A 0.48fF
C27269 NAND2X1_LOC_156/B INVX1_LOC_117/Y 0.16fF
C27270 NOR2X1_LOC_639/B NOR2X1_LOC_636/B 0.02fF
C27271 INVX1_LOC_45/A NOR2X1_LOC_318/a_36_216# 0.00fF
C27272 INVX1_LOC_36/A NAND2X1_LOC_286/B 0.01fF
C27273 INVX1_LOC_22/A NOR2X1_LOC_485/Y 0.00fF
C27274 NAND2X1_LOC_849/A NOR2X1_LOC_536/A 0.05fF
C27275 INVX1_LOC_2/A INVX1_LOC_109/A 0.01fF
C27276 INVX1_LOC_95/A NAND2X1_LOC_642/Y 0.03fF
C27277 INVX1_LOC_33/A INVX1_LOC_15/A 3.18fF
C27278 INVX1_LOC_28/A INVX1_LOC_118/A 0.23fF
C27279 INVX1_LOC_305/A INVX1_LOC_26/Y 0.35fF
C27280 NAND2X1_LOC_796/B NAND2X1_LOC_579/A 0.02fF
C27281 NOR2X1_LOC_68/A NOR2X1_LOC_668/Y 0.04fF
C27282 NOR2X1_LOC_201/A NOR2X1_LOC_68/A 0.00fF
C27283 NAND2X1_LOC_354/B INVX1_LOC_231/A 0.17fF
C27284 NAND2X1_LOC_214/B NOR2X1_LOC_82/A 0.07fF
C27285 NAND2X1_LOC_387/a_36_24# INVX1_LOC_53/A 0.00fF
C27286 INVX1_LOC_298/Y INVX1_LOC_71/A 0.02fF
C27287 NOR2X1_LOC_128/B NOR2X1_LOC_649/B 0.03fF
C27288 NOR2X1_LOC_551/Y INVX1_LOC_117/A 0.02fF
C27289 NAND2X1_LOC_149/Y NOR2X1_LOC_210/a_36_216# -0.00fF
C27290 NAND2X1_LOC_466/A INVX1_LOC_15/A 0.00fF
C27291 INVX1_LOC_58/A NAND2X1_LOC_726/a_36_24# 0.01fF
C27292 NOR2X1_LOC_128/B INVX1_LOC_3/A 0.08fF
C27293 NOR2X1_LOC_482/Y NOR2X1_LOC_754/A 0.01fF
C27294 NOR2X1_LOC_197/A INVX1_LOC_5/A 0.01fF
C27295 INVX1_LOC_16/A NAND2X1_LOC_63/Y 0.03fF
C27296 NAND2X1_LOC_721/A NOR2X1_LOC_528/Y 0.03fF
C27297 NOR2X1_LOC_457/a_36_216# NOR2X1_LOC_15/Y 0.00fF
C27298 INVX1_LOC_36/A NAND2X1_LOC_860/A 0.15fF
C27299 INVX1_LOC_255/Y NAND2X1_LOC_82/Y 0.05fF
C27300 NOR2X1_LOC_78/B INVX1_LOC_290/Y 0.08fF
C27301 NOR2X1_LOC_68/A INVX1_LOC_23/A 2.67fF
C27302 NOR2X1_LOC_609/A INVX1_LOC_57/A 0.03fF
C27303 NOR2X1_LOC_15/Y NOR2X1_LOC_468/Y 0.04fF
C27304 INVX1_LOC_27/A NOR2X1_LOC_82/A 0.32fF
C27305 VDD INPUT_4 0.17fF
C27306 NOR2X1_LOC_714/Y INVX1_LOC_15/A 0.01fF
C27307 INVX1_LOC_71/A NOR2X1_LOC_318/a_36_216# 0.00fF
C27308 NOR2X1_LOC_92/Y INVX1_LOC_258/A 0.15fF
C27309 NOR2X1_LOC_94/a_36_216# NOR2X1_LOC_671/Y 0.00fF
C27310 INVX1_LOC_269/A NOR2X1_LOC_793/A 0.27fF
C27311 NOR2X1_LOC_528/Y NOR2X1_LOC_323/a_36_216# 0.01fF
C27312 NAND2X1_LOC_141/A NOR2X1_LOC_38/B 0.04fF
C27313 NAND2X1_LOC_634/Y NAND2X1_LOC_793/B 0.04fF
C27314 NOR2X1_LOC_67/A INVX1_LOC_3/Y 0.28fF
C27315 INVX1_LOC_21/A INVX1_LOC_174/A 0.15fF
C27316 NAND2X1_LOC_563/A NOR2X1_LOC_554/A 0.01fF
C27317 NAND2X1_LOC_850/Y INVX1_LOC_32/A 0.10fF
C27318 NOR2X1_LOC_186/Y NOR2X1_LOC_441/Y 0.04fF
C27319 NAND2X1_LOC_364/Y NOR2X1_LOC_383/B 0.06fF
C27320 NOR2X1_LOC_456/Y INVX1_LOC_24/A 0.07fF
C27321 NOR2X1_LOC_561/Y INVX1_LOC_12/A 0.22fF
C27322 NOR2X1_LOC_433/A NOR2X1_LOC_677/Y 0.03fF
C27323 NAND2X1_LOC_483/Y NOR2X1_LOC_693/Y 0.00fF
C27324 NOR2X1_LOC_419/Y INVX1_LOC_57/A 0.18fF
C27325 INVX1_LOC_35/A INVX1_LOC_159/A 0.07fF
C27326 NOR2X1_LOC_323/Y NOR2X1_LOC_88/Y 0.03fF
C27327 NOR2X1_LOC_276/a_36_216# NOR2X1_LOC_678/A 0.00fF
C27328 INVX1_LOC_279/A INVX1_LOC_99/A 0.14fF
C27329 INVX1_LOC_6/A NOR2X1_LOC_487/Y 0.02fF
C27330 NOR2X1_LOC_643/A NAND2X1_LOC_20/B 0.01fF
C27331 NOR2X1_LOC_453/Y INVX1_LOC_174/A 0.02fF
C27332 NOR2X1_LOC_16/Y NAND2X1_LOC_223/A 0.04fF
C27333 NOR2X1_LOC_716/B INVX1_LOC_57/A 0.21fF
C27334 INVX1_LOC_58/A NOR2X1_LOC_753/Y 0.03fF
C27335 INVX1_LOC_245/Y INVX1_LOC_1/A 0.03fF
C27336 INVX1_LOC_103/A NAND2X1_LOC_192/a_36_24# 0.02fF
C27337 INVX1_LOC_223/Y NOR2X1_LOC_336/B 0.00fF
C27338 NOR2X1_LOC_134/Y INVX1_LOC_48/Y 0.03fF
C27339 NOR2X1_LOC_577/Y INVX1_LOC_29/Y 0.08fF
C27340 INVX1_LOC_11/A NOR2X1_LOC_533/Y 0.03fF
C27341 NOR2X1_LOC_824/A NAND2X1_LOC_500/Y 0.03fF
C27342 NAND2X1_LOC_860/A NOR2X1_LOC_237/Y 0.07fF
C27343 NOR2X1_LOC_711/A NOR2X1_LOC_155/A 0.01fF
C27344 INVX1_LOC_77/A INVX1_LOC_53/A 0.27fF
C27345 NOR2X1_LOC_437/Y NOR2X1_LOC_678/A 0.06fF
C27346 NOR2X1_LOC_309/Y NAND2X1_LOC_286/B 0.01fF
C27347 NOR2X1_LOC_602/B NAND2X1_LOC_642/Y 0.02fF
C27348 INVX1_LOC_269/A NOR2X1_LOC_160/B 0.24fF
C27349 INVX1_LOC_85/Y INVX1_LOC_301/A 0.03fF
C27350 INVX1_LOC_224/Y INVX1_LOC_8/A 2.36fF
C27351 NAND2X1_LOC_332/Y INVX1_LOC_271/A 0.02fF
C27352 NOR2X1_LOC_609/A NAND2X1_LOC_608/a_36_24# 0.02fF
C27353 D_INPUT_1 NOR2X1_LOC_772/Y 0.02fF
C27354 INVX1_LOC_58/A NAND2X1_LOC_325/Y 0.01fF
C27355 INVX1_LOC_224/Y NAND2X1_LOC_399/a_36_24# 0.01fF
C27356 INVX1_LOC_78/Y INVX1_LOC_179/A 0.03fF
C27357 NAND2X1_LOC_200/B INVX1_LOC_87/A 0.00fF
C27358 INVX1_LOC_284/Y NOR2X1_LOC_494/Y 0.20fF
C27359 INVX1_LOC_36/A NAND2X1_LOC_473/A 0.01fF
C27360 NOR2X1_LOC_78/A NOR2X1_LOC_622/a_36_216# 0.00fF
C27361 NOR2X1_LOC_329/B INVX1_LOC_133/A 0.01fF
C27362 INVX1_LOC_48/A NAND2X1_LOC_85/Y 0.01fF
C27363 NAND2X1_LOC_7/a_36_24# INVX1_LOC_125/A 0.00fF
C27364 NOR2X1_LOC_773/Y NOR2X1_LOC_278/Y 0.07fF
C27365 INVX1_LOC_256/A NAND2X1_LOC_352/B 0.02fF
C27366 INVX1_LOC_27/A NAND2X1_LOC_153/a_36_24# 0.06fF
C27367 INVX1_LOC_5/A NAND2X1_LOC_7/Y 0.04fF
C27368 NOR2X1_LOC_318/B NOR2X1_LOC_216/B 0.07fF
C27369 NOR2X1_LOC_309/Y NOR2X1_LOC_15/a_36_216# 0.00fF
C27370 INVX1_LOC_259/Y NOR2X1_LOC_718/B 0.00fF
C27371 INVX1_LOC_36/A NAND2X1_LOC_537/Y 0.17fF
C27372 NOR2X1_LOC_774/a_36_216# NAND2X1_LOC_175/Y 0.00fF
C27373 INVX1_LOC_102/Y INVX1_LOC_29/A 0.07fF
C27374 NAND2X1_LOC_473/a_36_24# NOR2X1_LOC_649/B 0.01fF
C27375 NAND2X1_LOC_714/B INVX1_LOC_24/A 0.03fF
C27376 NAND2X1_LOC_738/B NOR2X1_LOC_504/Y 0.08fF
C27377 INVX1_LOC_256/A INVX1_LOC_81/Y 0.01fF
C27378 INVX1_LOC_58/A INVX1_LOC_133/Y 0.03fF
C27379 D_INPUT_0 NOR2X1_LOC_801/B 0.18fF
C27380 INVX1_LOC_236/Y NOR2X1_LOC_816/A 0.03fF
C27381 INVX1_LOC_93/Y NOR2X1_LOC_216/B 0.10fF
C27382 INVX1_LOC_124/A INVX1_LOC_53/A 0.02fF
C27383 INVX1_LOC_136/A INVX1_LOC_308/Y 0.03fF
C27384 NOR2X1_LOC_441/Y NOR2X1_LOC_45/Y 0.00fF
C27385 NAND2X1_LOC_57/a_36_24# NOR2X1_LOC_103/Y 0.00fF
C27386 INVX1_LOC_58/A NOR2X1_LOC_67/A 0.08fF
C27387 D_INPUT_1 NAND2X1_LOC_294/a_36_24# 0.01fF
C27388 INVX1_LOC_64/A INVX1_LOC_158/A 0.00fF
C27389 INVX1_LOC_11/A NAND2X1_LOC_351/A 0.00fF
C27390 NOR2X1_LOC_430/A NOR2X1_LOC_763/A 0.02fF
C27391 NOR2X1_LOC_15/Y NOR2X1_LOC_596/A 0.08fF
C27392 NOR2X1_LOC_366/B NOR2X1_LOC_125/Y 0.01fF
C27393 NAND2X1_LOC_357/A NAND2X1_LOC_364/A 0.40fF
C27394 INVX1_LOC_17/A NOR2X1_LOC_360/Y 0.11fF
C27395 NOR2X1_LOC_430/A NOR2X1_LOC_582/A 0.10fF
C27396 NOR2X1_LOC_599/Y NOR2X1_LOC_761/Y 0.07fF
C27397 INVX1_LOC_13/A NOR2X1_LOC_720/A 0.01fF
C27398 NOR2X1_LOC_392/B NOR2X1_LOC_652/Y 0.10fF
C27399 NAND2X1_LOC_35/Y NAND2X1_LOC_839/Y 0.08fF
C27400 INVX1_LOC_22/A INVX1_LOC_29/Y 0.19fF
C27401 NOR2X1_LOC_331/Y NAND2X1_LOC_355/Y 0.06fF
C27402 NOR2X1_LOC_68/A NAND2X1_LOC_179/a_36_24# 0.01fF
C27403 INVX1_LOC_59/A INVX1_LOC_34/A 0.00fF
C27404 NOR2X1_LOC_455/Y NOR2X1_LOC_500/Y -0.02fF
C27405 NOR2X1_LOC_175/A INVX1_LOC_50/Y 0.05fF
C27406 NOR2X1_LOC_687/Y INVX1_LOC_53/A 2.50fF
C27407 NOR2X1_LOC_68/A INVX1_LOC_31/A 0.83fF
C27408 INVX1_LOC_232/Y INVX1_LOC_5/A 0.00fF
C27409 NOR2X1_LOC_189/A NAND2X1_LOC_787/a_36_24# 0.00fF
C27410 NAND2X1_LOC_751/a_36_24# INVX1_LOC_232/A 0.00fF
C27411 NOR2X1_LOC_598/B NAND2X1_LOC_479/Y 0.01fF
C27412 NAND2X1_LOC_360/B INVX1_LOC_306/Y 0.04fF
C27413 INVX1_LOC_307/A NAND2X1_LOC_418/a_36_24# 0.00fF
C27414 INVX1_LOC_2/A NAND2X1_LOC_794/B 0.01fF
C27415 NOR2X1_LOC_295/Y NOR2X1_LOC_15/Y 0.02fF
C27416 NOR2X1_LOC_100/A INVX1_LOC_27/A 0.03fF
C27417 NOR2X1_LOC_636/A INVX1_LOC_11/A 0.08fF
C27418 INVX1_LOC_10/Y NOR2X1_LOC_155/A 0.56fF
C27419 NOR2X1_LOC_549/a_36_216# INVX1_LOC_53/A 0.01fF
C27420 NOR2X1_LOC_19/B INVX1_LOC_175/A 0.03fF
C27421 D_INPUT_7 INVX1_LOC_18/A 0.05fF
C27422 INVX1_LOC_25/A D_INPUT_0 0.49fF
C27423 INVX1_LOC_9/A INVX1_LOC_92/A 0.10fF
C27424 INVX1_LOC_256/A NOR2X1_LOC_344/A 0.01fF
C27425 NOR2X1_LOC_103/Y INVX1_LOC_8/A 0.11fF
C27426 NOR2X1_LOC_78/A NOR2X1_LOC_850/B 0.02fF
C27427 NOR2X1_LOC_331/B NOR2X1_LOC_58/Y 0.07fF
C27428 NOR2X1_LOC_169/a_36_216# INVX1_LOC_91/A 0.01fF
C27429 VDD NOR2X1_LOC_691/B 0.03fF
C27430 NAND2X1_LOC_63/Y NOR2X1_LOC_35/Y 0.01fF
C27431 NOR2X1_LOC_454/Y NOR2X1_LOC_78/B 0.01fF
C27432 INVX1_LOC_190/A INVX1_LOC_53/A 0.01fF
C27433 NOR2X1_LOC_598/B INVX1_LOC_135/A 0.17fF
C27434 INPUT_0 INVX1_LOC_271/Y 0.00fF
C27435 INVX1_LOC_199/A NAND2X1_LOC_469/a_36_24# 0.02fF
C27436 NAND2X1_LOC_585/a_36_24# NOR2X1_LOC_590/A 0.01fF
C27437 NOR2X1_LOC_510/Y NOR2X1_LOC_269/a_36_216# 0.00fF
C27438 NOR2X1_LOC_272/Y INVX1_LOC_25/Y 0.03fF
C27439 INVX1_LOC_163/A INVX1_LOC_197/A 0.01fF
C27440 D_INPUT_1 INVX1_LOC_90/A 0.30fF
C27441 INVX1_LOC_39/A INVX1_LOC_16/A 0.11fF
C27442 NOR2X1_LOC_590/A NAND2X1_LOC_276/Y 0.03fF
C27443 INVX1_LOC_269/A NOR2X1_LOC_399/a_36_216# 0.00fF
C27444 INVX1_LOC_37/A INVX1_LOC_262/Y 0.02fF
C27445 D_INPUT_1 NOR2X1_LOC_389/B 0.08fF
C27446 NAND2X1_LOC_634/Y INVX1_LOC_71/A 0.00fF
C27447 INVX1_LOC_12/A INVX1_LOC_76/A 0.43fF
C27448 INVX1_LOC_6/A NAND2X1_LOC_454/Y 0.16fF
C27449 NOR2X1_LOC_15/Y NOR2X1_LOC_220/A 0.10fF
C27450 INVX1_LOC_21/A NOR2X1_LOC_589/A 0.10fF
C27451 NOR2X1_LOC_273/Y INVX1_LOC_24/A 0.05fF
C27452 INVX1_LOC_45/A NAND2X1_LOC_310/a_36_24# 0.00fF
C27453 INVX1_LOC_123/A NAND2X1_LOC_223/A 0.07fF
C27454 INVX1_LOC_225/A NOR2X1_LOC_441/Y 0.03fF
C27455 NAND2X1_LOC_552/A NOR2X1_LOC_312/Y 0.01fF
C27456 INVX1_LOC_24/A NOR2X1_LOC_759/Y 0.00fF
C27457 INVX1_LOC_269/A INVX1_LOC_208/A 0.00fF
C27458 INVX1_LOC_45/A INVX1_LOC_8/A 0.07fF
C27459 NOR2X1_LOC_486/Y INVX1_LOC_15/A 0.07fF
C27460 NOR2X1_LOC_205/Y INVX1_LOC_52/A 0.01fF
C27461 NOR2X1_LOC_425/a_36_216# INVX1_LOC_286/Y 0.00fF
C27462 INVX1_LOC_276/A INVX1_LOC_215/Y 0.03fF
C27463 INVX1_LOC_188/A INVX1_LOC_266/Y 0.00fF
C27464 INVX1_LOC_269/A NOR2X1_LOC_516/B 0.41fF
C27465 NOR2X1_LOC_615/Y NAND2X1_LOC_374/Y 0.04fF
C27466 INVX1_LOC_290/Y INVX1_LOC_46/A 0.07fF
C27467 D_INPUT_1 NAND2X1_LOC_348/A 0.03fF
C27468 NAND2X1_LOC_253/a_36_24# INVX1_LOC_76/A 0.00fF
C27469 INVX1_LOC_147/A INVX1_LOC_23/A 0.26fF
C27470 INVX1_LOC_27/A INVX1_LOC_306/A 0.01fF
C27471 NOR2X1_LOC_595/Y INVX1_LOC_94/Y 0.01fF
C27472 NOR2X1_LOC_226/A INVX1_LOC_246/A 0.20fF
C27473 INVX1_LOC_33/A NOR2X1_LOC_168/Y 0.64fF
C27474 VDD NOR2X1_LOC_477/B 0.00fF
C27475 NOR2X1_LOC_778/B INVX1_LOC_292/A 0.07fF
C27476 INVX1_LOC_11/A INVX1_LOC_56/Y 0.03fF
C27477 INVX1_LOC_90/A NOR2X1_LOC_652/Y 0.11fF
C27478 NOR2X1_LOC_454/Y INVX1_LOC_83/A 0.10fF
C27479 NOR2X1_LOC_331/B INVX1_LOC_29/A 0.07fF
C27480 NOR2X1_LOC_703/B INVX1_LOC_104/A 0.08fF
C27481 NOR2X1_LOC_389/B NOR2X1_LOC_652/Y 0.11fF
C27482 NOR2X1_LOC_82/A INVX1_LOC_137/A 0.00fF
C27483 INVX1_LOC_49/A NOR2X1_LOC_350/A 0.00fF
C27484 NOR2X1_LOC_48/Y INVX1_LOC_54/A 0.01fF
C27485 NOR2X1_LOC_802/A INVX1_LOC_18/A 0.10fF
C27486 D_INPUT_0 INVX1_LOC_1/A 0.23fF
C27487 NAND2X1_LOC_642/a_36_24# INVX1_LOC_15/A 0.01fF
C27488 NOR2X1_LOC_510/Y NOR2X1_LOC_329/B 0.07fF
C27489 INVX1_LOC_71/A INVX1_LOC_8/A 0.01fF
C27490 INVX1_LOC_24/A INVX1_LOC_249/Y 0.01fF
C27491 NAND2X1_LOC_854/B INVX1_LOC_221/Y 0.17fF
C27492 NAND2X1_LOC_35/Y INVX1_LOC_91/Y 0.02fF
C27493 NOR2X1_LOC_791/B INVX1_LOC_34/Y 0.16fF
C27494 INVX1_LOC_48/Y INPUT_1 0.25fF
C27495 NOR2X1_LOC_82/A INVX1_LOC_234/A 0.17fF
C27496 NOR2X1_LOC_655/Y NOR2X1_LOC_610/a_36_216# 0.00fF
C27497 INVX1_LOC_91/A NOR2X1_LOC_441/a_36_216# 0.01fF
C27498 NOR2X1_LOC_607/Y NOR2X1_LOC_392/B 0.05fF
C27499 NOR2X1_LOC_860/B NOR2X1_LOC_844/A 0.06fF
C27500 NOR2X1_LOC_481/A NOR2X1_LOC_142/Y 0.10fF
C27501 NOR2X1_LOC_590/A NOR2X1_LOC_553/B 0.03fF
C27502 NAND2X1_LOC_564/B NAND2X1_LOC_860/a_36_24# 0.01fF
C27503 NOR2X1_LOC_596/A INVX1_LOC_96/Y 0.01fF
C27504 NAND2X1_LOC_622/B INVX1_LOC_253/Y 0.15fF
C27505 NOR2X1_LOC_272/Y INVX1_LOC_75/A 0.07fF
C27506 INVX1_LOC_88/A NOR2X1_LOC_473/B 0.02fF
C27507 NAND2X1_LOC_779/a_36_24# NOR2X1_LOC_816/A 0.00fF
C27508 NAND2X1_LOC_733/Y NOR2X1_LOC_561/Y 0.10fF
C27509 INVX1_LOC_5/A NOR2X1_LOC_391/Y 0.01fF
C27510 NOR2X1_LOC_312/Y NAND2X1_LOC_337/B 0.14fF
C27511 INVX1_LOC_210/Y NAND2X1_LOC_41/Y 0.10fF
C27512 INVX1_LOC_34/A NOR2X1_LOC_144/Y 0.01fF
C27513 NAND2X1_LOC_731/Y NOR2X1_LOC_773/Y 0.01fF
C27514 NOR2X1_LOC_518/Y NAND2X1_LOC_170/A 0.06fF
C27515 NOR2X1_LOC_351/Y INVX1_LOC_15/A 0.01fF
C27516 INVX1_LOC_135/A NOR2X1_LOC_372/A 0.07fF
C27517 NOR2X1_LOC_361/B NOR2X1_LOC_329/B 0.17fF
C27518 NOR2X1_LOC_626/Y INVX1_LOC_311/A 0.04fF
C27519 INVX1_LOC_41/A NOR2X1_LOC_180/Y 0.01fF
C27520 NOR2X1_LOC_89/A NOR2X1_LOC_831/B 0.08fF
C27521 INVX1_LOC_21/A INVX1_LOC_222/A 0.04fF
C27522 NAND2X1_LOC_213/A INVX1_LOC_75/A 0.03fF
C27523 NOR2X1_LOC_86/Y NOR2X1_LOC_86/A 0.13fF
C27524 INVX1_LOC_61/A INVX1_LOC_16/A 0.02fF
C27525 NOR2X1_LOC_78/B INVX1_LOC_77/A 0.13fF
C27526 INVX1_LOC_59/A INPUT_0 0.03fF
C27527 NAND2X1_LOC_35/Y NOR2X1_LOC_45/B 0.17fF
C27528 INVX1_LOC_132/A NOR2X1_LOC_655/B 0.10fF
C27529 INVX1_LOC_284/A INVX1_LOC_123/Y 0.04fF
C27530 INVX1_LOC_293/Y NAND2X1_LOC_773/B 0.16fF
C27531 NOR2X1_LOC_151/Y NOR2X1_LOC_666/Y 0.02fF
C27532 INVX1_LOC_125/A NOR2X1_LOC_814/A 0.01fF
C27533 INVX1_LOC_90/A NAND2X1_LOC_805/a_36_24# 0.00fF
C27534 NOR2X1_LOC_82/A NOR2X1_LOC_19/B 0.19fF
C27535 NOR2X1_LOC_432/a_36_216# INVX1_LOC_34/A 0.02fF
C27536 NAND2X1_LOC_773/Y INPUT_0 0.05fF
C27537 NOR2X1_LOC_420/a_36_216# NOR2X1_LOC_78/A 0.00fF
C27538 INVX1_LOC_35/A NOR2X1_LOC_56/Y 0.07fF
C27539 NAND2X1_LOC_703/Y NAND2X1_LOC_851/a_36_24# 0.00fF
C27540 NAND2X1_LOC_782/B INVX1_LOC_301/A 0.08fF
C27541 NOR2X1_LOC_6/B NOR2X1_LOC_175/A 0.02fF
C27542 INVX1_LOC_254/A NOR2X1_LOC_619/A 0.08fF
C27543 INVX1_LOC_298/Y NOR2X1_LOC_331/B 0.07fF
C27544 INVX1_LOC_64/A NOR2X1_LOC_332/B 0.02fF
C27545 NOR2X1_LOC_536/A NOR2X1_LOC_282/Y 0.03fF
C27546 D_INPUT_0 NOR2X1_LOC_384/Y 1.07fF
C27547 NOR2X1_LOC_261/a_36_216# INVX1_LOC_37/A 0.00fF
C27548 INVX1_LOC_292/A NAND2X1_LOC_123/Y 0.07fF
C27549 NOR2X1_LOC_760/a_36_216# INVX1_LOC_73/A 0.02fF
C27550 INVX1_LOC_21/A NOR2X1_LOC_311/a_36_216# 0.00fF
C27551 NOR2X1_LOC_655/B INVX1_LOC_225/A 0.10fF
C27552 INVX1_LOC_36/A NAND2X1_LOC_128/a_36_24# 0.01fF
C27553 NOR2X1_LOC_788/B INVX1_LOC_30/A 0.71fF
C27554 NOR2X1_LOC_773/Y NOR2X1_LOC_561/a_36_216# 0.00fF
C27555 INVX1_LOC_49/A NOR2X1_LOC_374/B 0.00fF
C27556 NAND2X1_LOC_571/Y NOR2X1_LOC_45/B 0.28fF
C27557 NAND2X1_LOC_477/A NAND2X1_LOC_470/a_36_24# 0.02fF
C27558 INVX1_LOC_290/A INVX1_LOC_49/A 0.07fF
C27559 INVX1_LOC_45/Y NAND2X1_LOC_656/Y 0.08fF
C27560 NOR2X1_LOC_220/B INVX1_LOC_95/Y 0.10fF
C27561 NAND2X1_LOC_214/B INVX1_LOC_59/Y 0.04fF
C27562 NOR2X1_LOC_532/Y INVX1_LOC_18/A 0.03fF
C27563 INVX1_LOC_174/A NAND2X1_LOC_51/B 0.25fF
C27564 INVX1_LOC_35/A VDD 2.12fF
C27565 NOR2X1_LOC_15/Y INVX1_LOC_100/Y 0.01fF
C27566 INVX1_LOC_72/A D_GATE_366 0.07fF
C27567 NOR2X1_LOC_577/Y INVX1_LOC_101/A 0.01fF
C27568 NOR2X1_LOC_731/a_36_216# NOR2X1_LOC_738/A 0.03fF
C27569 NOR2X1_LOC_251/a_36_216# INVX1_LOC_91/A -0.01fF
C27570 INVX1_LOC_200/A NOR2X1_LOC_167/Y 0.01fF
C27571 NOR2X1_LOC_226/A NOR2X1_LOC_84/Y 0.01fF
C27572 NOR2X1_LOC_388/Y NOR2X1_LOC_570/A 0.02fF
C27573 NAND2X1_LOC_338/B NOR2X1_LOC_520/A 0.00fF
C27574 INVX1_LOC_64/A NAND2X1_LOC_804/Y 0.07fF
C27575 NAND2X1_LOC_717/Y NAND2X1_LOC_733/B 0.03fF
C27576 INVX1_LOC_83/A INVX1_LOC_77/A 1.99fF
C27577 INVX1_LOC_36/A NAND2X1_LOC_855/Y 0.07fF
C27578 NOR2X1_LOC_709/B INVX1_LOC_57/A 0.02fF
C27579 NOR2X1_LOC_52/B INVX1_LOC_56/Y 0.01fF
C27580 NAND2X1_LOC_841/A INVX1_LOC_266/Y 0.02fF
C27581 INVX1_LOC_27/A NOR2X1_LOC_300/a_36_216# 0.01fF
C27582 NOR2X1_LOC_48/B NOR2X1_LOC_48/Y 0.01fF
C27583 NOR2X1_LOC_336/B INVX1_LOC_75/A 0.00fF
C27584 NOR2X1_LOC_68/A NAND2X1_LOC_807/Y 0.10fF
C27585 NAND2X1_LOC_149/Y NAND2X1_LOC_212/Y 0.05fF
C27586 INVX1_LOC_5/A NOR2X1_LOC_168/a_36_216# 0.02fF
C27587 INVX1_LOC_21/A INVX1_LOC_20/A 1.38fF
C27588 INVX1_LOC_34/A INVX1_LOC_279/A 0.11fF
C27589 NOR2X1_LOC_598/B INVX1_LOC_280/A 0.03fF
C27590 INVX1_LOC_27/A INVX1_LOC_176/A 0.03fF
C27591 INVX1_LOC_93/A NAND2X1_LOC_641/a_36_24# 0.01fF
C27592 NAND2X1_LOC_549/Y NOR2X1_LOC_536/A 0.02fF
C27593 NOR2X1_LOC_361/Y INVX1_LOC_22/A 0.04fF
C27594 INVX1_LOC_254/Y INVX1_LOC_89/A 0.02fF
C27595 NOR2X1_LOC_533/A NAND2X1_LOC_532/a_36_24# 0.00fF
C27596 D_GATE_741 NOR2X1_LOC_725/A 0.24fF
C27597 NOR2X1_LOC_627/a_36_216# INVX1_LOC_16/A 0.02fF
C27598 INVX1_LOC_53/A INVX1_LOC_9/A 0.52fF
C27599 INVX1_LOC_179/A NOR2X1_LOC_727/B 0.03fF
C27600 NAND2X1_LOC_364/A INVX1_LOC_75/A 0.08fF
C27601 INVX1_LOC_93/A NAND2X1_LOC_721/A 0.02fF
C27602 INVX1_LOC_54/Y INVX1_LOC_1/Y 0.54fF
C27603 INVX1_LOC_235/Y D_GATE_479 0.03fF
C27604 INVX1_LOC_103/A NOR2X1_LOC_657/B 0.02fF
C27605 INVX1_LOC_177/Y INVX1_LOC_79/A 0.01fF
C27606 INVX1_LOC_2/A INVX1_LOC_290/A 0.10fF
C27607 INVX1_LOC_269/A NOR2X1_LOC_324/B 0.02fF
C27608 INVX1_LOC_33/Y NOR2X1_LOC_406/A 0.02fF
C27609 NOR2X1_LOC_454/Y INVX1_LOC_46/A 0.02fF
C27610 INVX1_LOC_177/A INVX1_LOC_220/Y 0.01fF
C27611 NOR2X1_LOC_748/Y NOR2X1_LOC_537/Y 0.26fF
C27612 NOR2X1_LOC_123/B INVX1_LOC_8/A 0.00fF
C27613 NOR2X1_LOC_78/B NOR2X1_LOC_687/Y 0.03fF
C27614 NAND2X1_LOC_149/Y INVX1_LOC_14/Y 0.12fF
C27615 INVX1_LOC_163/A INVX1_LOC_178/Y 0.01fF
C27616 NAND2X1_LOC_564/B NAND2X1_LOC_850/Y 0.38fF
C27617 NOR2X1_LOC_561/A NOR2X1_LOC_652/Y 0.01fF
C27618 NAND2X1_LOC_563/A NOR2X1_LOC_516/B 0.01fF
C27619 NOR2X1_LOC_749/Y INVX1_LOC_8/A 0.03fF
C27620 INVX1_LOC_25/A INVX1_LOC_46/Y 0.09fF
C27621 INVX1_LOC_1/A NOR2X1_LOC_266/B 0.03fF
C27622 INVX1_LOC_202/A NOR2X1_LOC_216/Y 0.27fF
C27623 NOR2X1_LOC_742/A NOR2X1_LOC_303/Y 0.02fF
C27624 NAND2X1_LOC_222/A INVX1_LOC_3/A 0.05fF
C27625 NOR2X1_LOC_455/Y INVX1_LOC_307/A 0.00fF
C27626 INVX1_LOC_218/Y NAND2X1_LOC_642/Y 0.22fF
C27627 NOR2X1_LOC_68/A INVX1_LOC_6/A 0.03fF
C27628 NOR2X1_LOC_456/Y NOR2X1_LOC_197/B 0.10fF
C27629 INVX1_LOC_14/A INVX1_LOC_37/A 0.19fF
C27630 INVX1_LOC_194/A NAND2X1_LOC_624/A 0.03fF
C27631 NOR2X1_LOC_441/Y NAND2X1_LOC_642/Y 0.03fF
C27632 NAND2X1_LOC_286/B INVX1_LOC_63/A 0.04fF
C27633 INVX1_LOC_286/A NOR2X1_LOC_91/Y 0.05fF
C27634 NOR2X1_LOC_218/Y INVX1_LOC_290/A 0.66fF
C27635 INVX1_LOC_16/A NOR2X1_LOC_85/a_36_216# 0.01fF
C27636 INVX1_LOC_25/Y NOR2X1_LOC_86/A 0.45fF
C27637 INVX1_LOC_232/Y NOR2X1_LOC_332/A 0.09fF
C27638 NOR2X1_LOC_242/A INVX1_LOC_9/A 0.03fF
C27639 NAND2X1_LOC_347/B NOR2X1_LOC_536/A 0.02fF
C27640 NOR2X1_LOC_84/Y INPUT_1 0.13fF
C27641 INVX1_LOC_34/A INVX1_LOC_182/Y 0.04fF
C27642 NOR2X1_LOC_596/A NOR2X1_LOC_733/Y 0.05fF
C27643 NOR2X1_LOC_449/A INVX1_LOC_29/A 0.03fF
C27644 NOR2X1_LOC_502/Y VDD 0.38fF
C27645 NOR2X1_LOC_444/a_36_216# NOR2X1_LOC_814/A 0.01fF
C27646 INVX1_LOC_16/A INPUT_5 0.06fF
C27647 INVX1_LOC_193/Y NOR2X1_LOC_546/a_36_216# 0.00fF
C27648 D_GATE_366 INVX1_LOC_192/Y 0.45fF
C27649 INVX1_LOC_216/A INPUT_1 0.18fF
C27650 NAND2X1_LOC_581/Y D_INPUT_4 0.01fF
C27651 NOR2X1_LOC_312/Y NOR2X1_LOC_773/Y 0.04fF
C27652 NOR2X1_LOC_286/Y INVX1_LOC_117/A 0.03fF
C27653 NAND2X1_LOC_81/B NAND2X1_LOC_99/A 0.03fF
C27654 NAND2X1_LOC_733/Y INVX1_LOC_76/A 0.17fF
C27655 NAND2X1_LOC_651/B NOR2X1_LOC_635/B 0.63fF
C27656 NOR2X1_LOC_329/B INVX1_LOC_177/A 0.56fF
C27657 INVX1_LOC_217/A NOR2X1_LOC_164/a_36_216# 0.00fF
C27658 NOR2X1_LOC_781/a_36_216# INVX1_LOC_290/A 0.01fF
C27659 NAND2X1_LOC_860/A INVX1_LOC_63/A 0.04fF
C27660 INVX1_LOC_83/A NOR2X1_LOC_687/Y 0.03fF
C27661 NOR2X1_LOC_746/Y INVX1_LOC_198/Y 0.31fF
C27662 NOR2X1_LOC_544/A NOR2X1_LOC_180/B 0.28fF
C27663 NOR2X1_LOC_576/B NAND2X1_LOC_863/B 0.69fF
C27664 INVX1_LOC_104/A INVX1_LOC_79/A 0.02fF
C27665 NOR2X1_LOC_160/B INVX1_LOC_12/Y 0.11fF
C27666 NOR2X1_LOC_516/B NOR2X1_LOC_814/Y 0.01fF
C27667 INVX1_LOC_72/Y INVX1_LOC_95/Y 0.01fF
C27668 INVX1_LOC_33/A NOR2X1_LOC_548/a_36_216# 0.00fF
C27669 NAND2X1_LOC_647/B NOR2X1_LOC_334/Y 0.01fF
C27670 INVX1_LOC_90/A NOR2X1_LOC_553/Y 0.05fF
C27671 NAND2X1_LOC_354/Y INVX1_LOC_20/A 0.00fF
C27672 NAND2X1_LOC_347/B NAND2X1_LOC_93/B 0.11fF
C27673 NAND2X1_LOC_624/B NAND2X1_LOC_489/Y 0.01fF
C27674 INVX1_LOC_217/A INVX1_LOC_76/A 0.07fF
C27675 INVX1_LOC_93/Y NOR2X1_LOC_303/Y 0.09fF
C27676 INVX1_LOC_73/Y INVX1_LOC_54/A 0.01fF
C27677 INVX1_LOC_104/A NOR2X1_LOC_728/B 0.06fF
C27678 NAND2X1_LOC_67/Y INVX1_LOC_92/A 0.96fF
C27679 INVX1_LOC_14/A NOR2X1_LOC_743/Y 0.02fF
C27680 INVX1_LOC_58/A NOR2X1_LOC_584/Y 0.02fF
C27681 INVX1_LOC_35/A INVX1_LOC_133/A 0.26fF
C27682 NOR2X1_LOC_551/B NOR2X1_LOC_78/A 0.03fF
C27683 NOR2X1_LOC_168/A NOR2X1_LOC_337/A 0.01fF
C27684 INVX1_LOC_246/A INVX1_LOC_118/A 0.03fF
C27685 NOR2X1_LOC_635/B INVX1_LOC_15/A 0.03fF
C27686 NOR2X1_LOC_78/B NAND2X1_LOC_832/Y 0.17fF
C27687 INVX1_LOC_136/A NAND2X1_LOC_472/Y 0.07fF
C27688 INVX1_LOC_197/Y NAND2X1_LOC_463/B 0.09fF
C27689 NOR2X1_LOC_411/A INVX1_LOC_12/A 0.18fF
C27690 NOR2X1_LOC_704/a_36_216# NOR2X1_LOC_78/A 0.00fF
C27691 NOR2X1_LOC_602/A NOR2X1_LOC_536/A 0.39fF
C27692 NOR2X1_LOC_45/B NAND2X1_LOC_465/Y 0.15fF
C27693 INVX1_LOC_296/A D_INPUT_5 0.22fF
C27694 INVX1_LOC_15/A INVX1_LOC_275/Y 0.00fF
C27695 INVX1_LOC_104/A INVX1_LOC_91/A 0.42fF
C27696 INVX1_LOC_15/A NOR2X1_LOC_748/A 0.17fF
C27697 INVX1_LOC_4/Y NAND2X1_LOC_99/A 0.10fF
C27698 NOR2X1_LOC_165/Y NOR2X1_LOC_74/A 0.15fF
C27699 NOR2X1_LOC_178/Y INVX1_LOC_12/A 0.07fF
C27700 NOR2X1_LOC_384/Y NAND2X1_LOC_848/A 0.07fF
C27701 NOR2X1_LOC_82/A NOR2X1_LOC_216/B 0.41fF
C27702 INVX1_LOC_45/A INVX1_LOC_118/Y 0.06fF
C27703 INVX1_LOC_63/A NAND2X1_LOC_473/A 0.33fF
C27704 NOR2X1_LOC_814/A NAND2X1_LOC_218/A 0.01fF
C27705 NAND2X1_LOC_787/B INVX1_LOC_76/A 0.06fF
C27706 INVX1_LOC_77/A INVX1_LOC_46/A 0.19fF
C27707 NOR2X1_LOC_589/A NAND2X1_LOC_51/B 0.00fF
C27708 NOR2X1_LOC_666/Y NOR2X1_LOC_666/a_36_216# 0.01fF
C27709 INVX1_LOC_304/Y NOR2X1_LOC_164/a_36_216# 0.01fF
C27710 NOR2X1_LOC_664/Y INVX1_LOC_59/Y 0.02fF
C27711 INVX1_LOC_40/A INVX1_LOC_123/A 0.19fF
C27712 NAND2X1_LOC_454/Y INVX1_LOC_270/A 0.07fF
C27713 NOR2X1_LOC_577/Y NOR2X1_LOC_111/A 0.07fF
C27714 INVX1_LOC_136/A NAND2X1_LOC_637/Y 0.06fF
C27715 NOR2X1_LOC_65/B NOR2X1_LOC_278/Y 0.00fF
C27716 NOR2X1_LOC_824/A NAND2X1_LOC_499/a_36_24# 0.01fF
C27717 NOR2X1_LOC_589/A INVX1_LOC_311/A 0.07fF
C27718 INVX1_LOC_54/Y INVX1_LOC_93/Y 0.11fF
C27719 INVX1_LOC_279/A INPUT_0 0.08fF
C27720 NOR2X1_LOC_655/B NAND2X1_LOC_642/Y 0.10fF
C27721 INVX1_LOC_53/A INVX1_LOC_274/Y 0.13fF
C27722 NOR2X1_LOC_91/Y INVX1_LOC_54/A 0.25fF
C27723 INVX1_LOC_299/A NOR2X1_LOC_856/B 0.01fF
C27724 INVX1_LOC_13/Y NAND2X1_LOC_456/a_36_24# 0.01fF
C27725 NOR2X1_LOC_233/a_36_216# NAND2X1_LOC_254/Y 0.00fF
C27726 INVX1_LOC_96/Y NAND2X1_LOC_469/B 0.00fF
C27727 NOR2X1_LOC_335/B INVX1_LOC_150/A 0.03fF
C27728 NOR2X1_LOC_736/Y NOR2X1_LOC_735/Y 0.09fF
C27729 INVX1_LOC_71/A INVX1_LOC_118/Y 0.06fF
C27730 INVX1_LOC_230/Y NOR2X1_LOC_673/A 0.07fF
C27731 D_INPUT_0 NOR2X1_LOC_188/A 0.03fF
C27732 NOR2X1_LOC_707/B NAND2X1_LOC_425/Y 0.03fF
C27733 INVX1_LOC_257/Y VDD -0.00fF
C27734 INVX1_LOC_28/A NAND2X1_LOC_680/a_36_24# 0.00fF
C27735 INVX1_LOC_57/A NOR2X1_LOC_39/a_36_216# 0.00fF
C27736 NAND2X1_LOC_808/A NOR2X1_LOC_167/Y 0.00fF
C27737 INVX1_LOC_124/A INVX1_LOC_46/A 0.12fF
C27738 D_INPUT_0 NOR2X1_LOC_548/B 0.01fF
C27739 NOR2X1_LOC_490/Y NAND2X1_LOC_560/A 0.03fF
C27740 NOR2X1_LOC_667/A INVX1_LOC_20/A 0.12fF
C27741 NOR2X1_LOC_598/B NOR2X1_LOC_541/B 0.02fF
C27742 NOR2X1_LOC_189/A INVX1_LOC_118/A 0.05fF
C27743 INVX1_LOC_24/A INVX1_LOC_75/Y 0.03fF
C27744 INVX1_LOC_248/A INVX1_LOC_20/A 0.29fF
C27745 NOR2X1_LOC_546/A NAND2X1_LOC_425/Y -0.01fF
C27746 NAND2X1_LOC_660/Y NOR2X1_LOC_43/Y 0.08fF
C27747 NOR2X1_LOC_82/A NAND2X1_LOC_82/a_36_24# 0.01fF
C27748 INVX1_LOC_21/A INVX1_LOC_4/A 0.03fF
C27749 NOR2X1_LOC_392/B NOR2X1_LOC_99/a_36_216# 0.01fF
C27750 NOR2X1_LOC_237/Y NOR2X1_LOC_487/Y 0.01fF
C27751 INVX1_LOC_90/A NAND2X1_LOC_814/a_36_24# 0.00fF
C27752 NOR2X1_LOC_773/Y NAND2X1_LOC_287/B 0.01fF
C27753 INVX1_LOC_305/Y VDD 0.28fF
C27754 INVX1_LOC_84/Y VDD 0.21fF
C27755 NOR2X1_LOC_750/Y NAND2X1_LOC_215/A -0.03fF
C27756 NOR2X1_LOC_561/Y NOR2X1_LOC_56/a_36_216# 0.01fF
C27757 NOR2X1_LOC_591/Y INVX1_LOC_38/A 2.47fF
C27758 NOR2X1_LOC_15/Y INVX1_LOC_251/A 0.01fF
C27759 NOR2X1_LOC_679/a_36_216# INVX1_LOC_42/A 0.00fF
C27760 NOR2X1_LOC_74/a_36_216# NOR2X1_LOC_74/A 0.02fF
C27761 VDD NOR2X1_LOC_121/A 0.41fF
C27762 NOR2X1_LOC_571/a_36_216# INPUT_4 0.00fF
C27763 INVX1_LOC_11/A NAND2X1_LOC_430/B 0.03fF
C27764 NOR2X1_LOC_433/A NOR2X1_LOC_831/B 0.09fF
C27765 NOR2X1_LOC_550/B NOR2X1_LOC_197/B 0.16fF
C27766 INVX1_LOC_136/A NAND2X1_LOC_773/B 0.03fF
C27767 INVX1_LOC_234/A INVX1_LOC_59/Y 0.08fF
C27768 INVX1_LOC_16/A INVX1_LOC_14/Y 0.01fF
C27769 INVX1_LOC_290/A NOR2X1_LOC_586/Y 0.06fF
C27770 INVX1_LOC_208/A INVX1_LOC_12/Y 0.11fF
C27771 NOR2X1_LOC_84/Y INVX1_LOC_118/A 0.19fF
C27772 NOR2X1_LOC_655/B NOR2X1_LOC_271/Y 0.03fF
C27773 VDD NOR2X1_LOC_188/Y 0.28fF
C27774 INVX1_LOC_236/Y INVX1_LOC_42/A 0.02fF
C27775 NAND2X1_LOC_858/B INPUT_0 0.01fF
C27776 NOR2X1_LOC_634/B INVX1_LOC_9/A 0.07fF
C27777 INVX1_LOC_24/A INVX1_LOC_293/Y -0.00fF
C27778 NOR2X1_LOC_78/B INVX1_LOC_9/A 0.19fF
C27779 NOR2X1_LOC_91/A NAND2X1_LOC_474/Y 0.51fF
C27780 NOR2X1_LOC_617/Y NAND2X1_LOC_489/Y 0.01fF
C27781 NOR2X1_LOC_68/A NOR2X1_LOC_633/A 0.05fF
C27782 NAND2X1_LOC_629/Y INVX1_LOC_92/A 0.01fF
C27783 INVX1_LOC_151/Y NOR2X1_LOC_331/B 0.03fF
C27784 NOR2X1_LOC_52/B NOR2X1_LOC_831/B 0.05fF
C27785 INVX1_LOC_161/Y NOR2X1_LOC_681/a_36_216# 0.00fF
C27786 INVX1_LOC_119/A NOR2X1_LOC_88/Y 0.11fF
C27787 NOR2X1_LOC_65/B NAND2X1_LOC_475/a_36_24# 0.00fF
C27788 INVX1_LOC_89/A NOR2X1_LOC_825/Y 0.10fF
C27789 INVX1_LOC_75/A NOR2X1_LOC_349/A 0.05fF
C27790 INVX1_LOC_24/A NAND2X1_LOC_74/B 0.39fF
C27791 INVX1_LOC_75/A NOR2X1_LOC_113/A 0.03fF
C27792 NOR2X1_LOC_45/B INVX1_LOC_144/A 1.18fF
C27793 INVX1_LOC_75/A NOR2X1_LOC_405/A 0.20fF
C27794 NAND2X1_LOC_159/a_36_24# NOR2X1_LOC_536/A 0.00fF
C27795 NOR2X1_LOC_229/a_36_216# INVX1_LOC_54/A 0.00fF
C27796 INVX1_LOC_243/A INVX1_LOC_92/A 0.01fF
C27797 NAND2X1_LOC_474/Y INVX1_LOC_23/A 0.07fF
C27798 NOR2X1_LOC_19/B INVX1_LOC_59/Y 0.03fF
C27799 INVX1_LOC_17/A INVX1_LOC_26/A 0.00fF
C27800 NAND2X1_LOC_208/B NOR2X1_LOC_38/B 0.04fF
C27801 NOR2X1_LOC_6/B INVX1_LOC_27/Y 0.03fF
C27802 NOR2X1_LOC_350/A NAND2X1_LOC_63/Y 0.03fF
C27803 INVX1_LOC_290/A INVX1_LOC_118/A 0.03fF
C27804 NOR2X1_LOC_91/Y NOR2X1_LOC_48/B 0.01fF
C27805 NOR2X1_LOC_91/A INVX1_LOC_272/Y 0.06fF
C27806 INVX1_LOC_35/A NOR2X1_LOC_510/Y 0.07fF
C27807 INVX1_LOC_303/A INVX1_LOC_106/A -0.03fF
C27808 INVX1_LOC_21/A INVX1_LOC_64/A 0.18fF
C27809 NAND2X1_LOC_123/Y NOR2X1_LOC_137/Y 0.03fF
C27810 INVX1_LOC_5/A INVX1_LOC_50/Y 0.07fF
C27811 NOR2X1_LOC_709/A NOR2X1_LOC_814/A 0.01fF
C27812 INVX1_LOC_86/Y INVX1_LOC_91/A 0.21fF
C27813 INVX1_LOC_103/A INVX1_LOC_271/A 0.00fF
C27814 NAND2X1_LOC_451/Y NOR2X1_LOC_430/Y 0.01fF
C27815 INVX1_LOC_83/A INVX1_LOC_9/A 0.07fF
C27816 NOR2X1_LOC_208/a_36_216# NOR2X1_LOC_197/B 0.00fF
C27817 NAND2X1_LOC_140/A NOR2X1_LOC_331/B 0.04fF
C27818 NOR2X1_LOC_388/Y INVX1_LOC_29/A 0.05fF
C27819 NOR2X1_LOC_230/Y NOR2X1_LOC_158/Y 0.06fF
C27820 INVX1_LOC_36/A NAND2X1_LOC_454/Y 0.03fF
C27821 INVX1_LOC_272/Y INVX1_LOC_23/A 0.05fF
C27822 INVX1_LOC_255/Y NOR2X1_LOC_820/a_36_216# 0.00fF
C27823 NAND2X1_LOC_53/Y INVX1_LOC_23/A 1.02fF
C27824 NOR2X1_LOC_717/B INVX1_LOC_274/A 0.00fF
C27825 NOR2X1_LOC_561/Y INVX1_LOC_92/A 0.17fF
C27826 INVX1_LOC_35/A NOR2X1_LOC_361/B 0.05fF
C27827 NAND2X1_LOC_778/Y NOR2X1_LOC_496/Y 0.03fF
C27828 INVX1_LOC_30/A NAND2X1_LOC_61/Y 0.07fF
C27829 INVX1_LOC_95/Y INVX1_LOC_125/Y 0.10fF
C27830 NOR2X1_LOC_770/a_36_216# NOR2X1_LOC_89/A 0.00fF
C27831 NOR2X1_LOC_790/B INVX1_LOC_11/A 0.06fF
C27832 INVX1_LOC_196/A INVX1_LOC_19/A 0.05fF
C27833 INVX1_LOC_224/A NAND2X1_LOC_69/a_36_24# 0.00fF
C27834 INVX1_LOC_135/A INVX1_LOC_152/A 0.12fF
C27835 NAND2X1_LOC_357/B NOR2X1_LOC_89/A 0.15fF
C27836 INVX1_LOC_49/A NOR2X1_LOC_467/A 0.07fF
C27837 NAND2X1_LOC_556/a_36_24# INVX1_LOC_12/A 0.01fF
C27838 INVX1_LOC_49/A NOR2X1_LOC_801/B 0.03fF
C27839 NOR2X1_LOC_828/A INVX1_LOC_274/A 0.03fF
C27840 NAND2X1_LOC_261/a_36_24# NOR2X1_LOC_342/A 0.00fF
C27841 INVX1_LOC_39/A INVX1_LOC_48/Y 0.54fF
C27842 INVX1_LOC_143/A NAND2X1_LOC_74/B 0.10fF
C27843 NOR2X1_LOC_208/Y NAND2X1_LOC_454/Y 0.10fF
C27844 NAND2X1_LOC_391/Y NOR2X1_LOC_92/Y 0.03fF
C27845 NOR2X1_LOC_91/Y NOR2X1_LOC_438/Y 0.01fF
C27846 INPUT_0 NOR2X1_LOC_98/B 0.00fF
C27847 NAND2X1_LOC_102/a_36_24# NOR2X1_LOC_271/Y 0.00fF
C27848 INVX1_LOC_89/A NOR2X1_LOC_88/Y 0.00fF
C27849 INVX1_LOC_30/A NOR2X1_LOC_452/A 0.06fF
C27850 INVX1_LOC_34/A NOR2X1_LOC_38/B 0.09fF
C27851 NAND2X1_LOC_593/Y NAND2X1_LOC_175/Y 0.02fF
C27852 NAND2X1_LOC_573/Y NAND2X1_LOC_579/A 0.09fF
C27853 NOR2X1_LOC_405/A NOR2X1_LOC_309/a_36_216# 0.00fF
C27854 INVX1_LOC_27/A INVX1_LOC_103/A 0.17fF
C27855 NOR2X1_LOC_565/A INVX1_LOC_53/A 0.03fF
C27856 NOR2X1_LOC_92/Y NAND2X1_LOC_576/a_36_24# 0.01fF
C27857 INVX1_LOC_150/A INVX1_LOC_84/A 0.01fF
C27858 INVX1_LOC_304/A INVX1_LOC_20/A 0.08fF
C27859 NOR2X1_LOC_151/Y INVX1_LOC_274/A 0.78fF
C27860 NAND2X1_LOC_545/a_36_24# INVX1_LOC_23/A 0.00fF
C27861 NAND2X1_LOC_565/B NAND2X1_LOC_74/B 0.06fF
C27862 INVX1_LOC_18/A INVX1_LOC_29/Y 0.27fF
C27863 NOR2X1_LOC_168/Y NOR2X1_LOC_748/A 0.13fF
C27864 NAND2X1_LOC_348/A NOR2X1_LOC_61/Y -0.02fF
C27865 NAND2X1_LOC_652/Y NAND2X1_LOC_798/B 0.03fF
C27866 NOR2X1_LOC_68/A NOR2X1_LOC_416/A 0.20fF
C27867 INVX1_LOC_22/A NOR2X1_LOC_583/Y 0.07fF
C27868 INVX1_LOC_89/A INVX1_LOC_84/A 0.24fF
C27869 NOR2X1_LOC_275/A NAND2X1_LOC_211/Y 0.06fF
C27870 NOR2X1_LOC_292/Y NOR2X1_LOC_612/Y 0.05fF
C27871 INVX1_LOC_298/Y NOR2X1_LOC_388/Y 0.07fF
C27872 INVX1_LOC_64/A NAND2X1_LOC_354/Y 0.07fF
C27873 INVX1_LOC_259/Y INVX1_LOC_24/A 0.00fF
C27874 NAND2X1_LOC_30/Y INVX1_LOC_1/A 0.56fF
C27875 NAND2X1_LOC_192/B NOR2X1_LOC_205/Y 0.01fF
C27876 INVX1_LOC_266/Y INVX1_LOC_271/Y 0.10fF
C27877 NOR2X1_LOC_516/B NOR2X1_LOC_554/A 0.00fF
C27878 NOR2X1_LOC_68/A NOR2X1_LOC_109/Y 0.14fF
C27879 INVX1_LOC_135/A INVX1_LOC_29/A 0.31fF
C27880 INVX1_LOC_223/A NOR2X1_LOC_674/Y 0.02fF
C27881 NOR2X1_LOC_167/Y INVX1_LOC_92/A 0.05fF
C27882 NOR2X1_LOC_264/Y NOR2X1_LOC_621/A 0.00fF
C27883 NOR2X1_LOC_130/A NAND2X1_LOC_74/B 20.44fF
C27884 INVX1_LOC_25/A INVX1_LOC_49/A 0.07fF
C27885 NAND2X1_LOC_803/B NAND2X1_LOC_538/Y 0.04fF
C27886 NOR2X1_LOC_793/A NOR2X1_LOC_160/B 0.03fF
C27887 NAND2X1_LOC_714/B INVX1_LOC_286/Y 0.07fF
C27888 INVX1_LOC_115/A INVX1_LOC_117/A 0.02fF
C27889 NAND2X1_LOC_9/Y INVX1_LOC_77/A 0.37fF
C27890 INVX1_LOC_11/A D_GATE_741 0.02fF
C27891 NOR2X1_LOC_736/Y INVX1_LOC_186/Y 0.03fF
C27892 NOR2X1_LOC_473/B INVX1_LOC_272/A 0.03fF
C27893 NAND2X1_LOC_787/A NOR2X1_LOC_753/Y 0.00fF
C27894 D_INPUT_1 INVX1_LOC_33/A 0.19fF
C27895 NOR2X1_LOC_401/A NOR2X1_LOC_160/B 0.13fF
C27896 NOR2X1_LOC_560/A INVX1_LOC_29/A 0.02fF
C27897 D_INPUT_7 D_INPUT_6 0.01fF
C27898 NOR2X1_LOC_468/Y NAND2X1_LOC_208/B 0.01fF
C27899 NOR2X1_LOC_590/A NAND2X1_LOC_538/Y 0.07fF
C27900 INVX1_LOC_83/A NOR2X1_LOC_861/Y 0.43fF
C27901 NOR2X1_LOC_312/Y INVX1_LOC_42/A 0.25fF
C27902 NOR2X1_LOC_9/Y NAND2X1_LOC_572/B 0.04fF
C27903 INVX1_LOC_196/A INVX1_LOC_26/Y 0.16fF
C27904 NOR2X1_LOC_35/Y INVX1_LOC_230/A 0.10fF
C27905 INVX1_LOC_17/A INVX1_LOC_141/A 0.02fF
C27906 INVX1_LOC_11/A NAND2X1_LOC_352/B 0.23fF
C27907 INVX1_LOC_89/A NAND2X1_LOC_220/B 0.13fF
C27908 INVX1_LOC_272/Y INVX1_LOC_31/A 0.31fF
C27909 NOR2X1_LOC_32/B NAND2X1_LOC_139/A 0.03fF
C27910 NOR2X1_LOC_181/A INVX1_LOC_274/A 0.03fF
C27911 NOR2X1_LOC_147/B NOR2X1_LOC_678/A 0.03fF
C27912 NOR2X1_LOC_808/A NOR2X1_LOC_383/B 0.04fF
C27913 INVX1_LOC_225/A INVX1_LOC_308/A 0.01fF
C27914 NAND2X1_LOC_451/Y INVX1_LOC_296/A 0.66fF
C27915 NOR2X1_LOC_210/A INVX1_LOC_78/A 0.22fF
C27916 INVX1_LOC_24/Y NOR2X1_LOC_703/B 0.03fF
C27917 INVX1_LOC_48/Y INVX1_LOC_61/A 0.02fF
C27918 NOR2X1_LOC_798/A INVX1_LOC_77/A 0.06fF
C27919 NAND2X1_LOC_103/a_36_24# NAND2X1_LOC_475/Y 0.06fF
C27920 INVX1_LOC_46/A INVX1_LOC_9/A 0.11fF
C27921 NOR2X1_LOC_795/Y NOR2X1_LOC_598/B 0.10fF
C27922 INVX1_LOC_25/A NOR2X1_LOC_818/Y 0.07fF
C27923 INVX1_LOC_89/A INVX1_LOC_15/A 0.48fF
C27924 NOR2X1_LOC_716/B INVX1_LOC_306/Y 0.53fF
C27925 NOR2X1_LOC_91/A INVX1_LOC_226/Y 0.11fF
C27926 NOR2X1_LOC_646/A NOR2X1_LOC_647/A 0.04fF
C27927 INVX1_LOC_233/A NAND2X1_LOC_650/a_36_24# 0.00fF
C27928 NAND2X1_LOC_785/Y INVX1_LOC_64/A 0.03fF
C27929 INVX1_LOC_247/A NOR2X1_LOC_155/A 0.01fF
C27930 NOR2X1_LOC_272/Y NOR2X1_LOC_577/Y 0.03fF
C27931 INVX1_LOC_33/A NOR2X1_LOC_652/Y 0.07fF
C27932 INVX1_LOC_2/Y NOR2X1_LOC_860/Y 0.02fF
C27933 INVX1_LOC_25/A NOR2X1_LOC_226/A 0.07fF
C27934 NOR2X1_LOC_852/B NOR2X1_LOC_242/A 0.04fF
C27935 INVX1_LOC_75/A INVX1_LOC_109/Y 0.10fF
C27936 INVX1_LOC_88/A NOR2X1_LOC_457/B 0.01fF
C27937 INVX1_LOC_40/A NAND2X1_LOC_90/a_36_24# 0.00fF
C27938 NOR2X1_LOC_750/Y NOR2X1_LOC_655/B 0.13fF
C27939 NOR2X1_LOC_216/B INVX1_LOC_59/Y 0.03fF
C27940 INVX1_LOC_35/A INVX1_LOC_177/A 2.49fF
C27941 INVX1_LOC_112/A NOR2X1_LOC_216/B 0.05fF
C27942 INVX1_LOC_76/A INVX1_LOC_92/A 0.25fF
C27943 NAND2X1_LOC_508/A INVX1_LOC_15/A 0.06fF
C27944 INVX1_LOC_27/A INVX1_LOC_67/A 0.03fF
C27945 INVX1_LOC_5/A NOR2X1_LOC_6/B 0.30fF
C27946 NOR2X1_LOC_328/Y INVX1_LOC_50/A 0.78fF
C27947 D_INPUT_1 INVX1_LOC_40/A 1.05fF
C27948 INVX1_LOC_179/Y INVX1_LOC_53/A 0.01fF
C27949 NOR2X1_LOC_312/Y INVX1_LOC_78/A 0.75fF
C27950 INVX1_LOC_278/A NOR2X1_LOC_401/B 0.00fF
C27951 NOR2X1_LOC_500/Y INVX1_LOC_23/A 0.04fF
C27952 D_INPUT_1 INVX1_LOC_165/Y 0.01fF
C27953 INVX1_LOC_226/Y INVX1_LOC_23/A 0.03fF
C27954 NOR2X1_LOC_602/a_36_216# NOR2X1_LOC_590/A 0.00fF
C27955 NOR2X1_LOC_226/A NAND2X1_LOC_370/a_36_24# 0.01fF
C27956 NOR2X1_LOC_488/a_36_216# NAND2X1_LOC_787/A 0.00fF
C27957 INVX1_LOC_278/A NOR2X1_LOC_402/a_36_216# 0.00fF
C27958 NOR2X1_LOC_91/A INVX1_LOC_10/A 0.29fF
C27959 INVX1_LOC_1/A INVX1_LOC_49/A 0.56fF
C27960 NOR2X1_LOC_794/A INVX1_LOC_29/A 0.05fF
C27961 INVX1_LOC_64/A NOR2X1_LOC_667/A 0.07fF
C27962 NOR2X1_LOC_331/B INVX1_LOC_118/Y 0.01fF
C27963 NOR2X1_LOC_598/B NOR2X1_LOC_614/Y 0.03fF
C27964 NOR2X1_LOC_346/B INVX1_LOC_138/Y 0.02fF
C27965 NAND2X1_LOC_39/Y INVX1_LOC_113/A 0.04fF
C27966 INVX1_LOC_124/A NOR2X1_LOC_798/A 0.02fF
C27967 INVX1_LOC_6/Y INVX1_LOC_103/A 0.01fF
C27968 NOR2X1_LOC_824/A INVX1_LOC_240/A 0.10fF
C27969 INVX1_LOC_85/Y NOR2X1_LOC_307/Y 0.01fF
C27970 NOR2X1_LOC_588/A NOR2X1_LOC_11/Y 0.10fF
C27971 NAND2X1_LOC_860/A INVX1_LOC_1/Y 0.00fF
C27972 NOR2X1_LOC_391/Y INVX1_LOC_42/A 0.00fF
C27973 INVX1_LOC_39/A NOR2X1_LOC_84/Y 0.08fF
C27974 INVX1_LOC_269/A INVX1_LOC_155/A 0.16fF
C27975 NOR2X1_LOC_753/a_36_216# NAND2X1_LOC_799/A 0.00fF
C27976 INVX1_LOC_34/A NOR2X1_LOC_468/Y 0.03fF
C27977 NOR2X1_LOC_328/Y NOR2X1_LOC_224/Y 0.01fF
C27978 NOR2X1_LOC_441/Y NOR2X1_LOC_91/Y 0.14fF
C27979 INVX1_LOC_237/A INVX1_LOC_240/A 0.03fF
C27980 INVX1_LOC_223/A INVX1_LOC_72/A 0.07fF
C27981 NOR2X1_LOC_264/a_36_216# NOR2X1_LOC_264/Y 0.00fF
C27982 INVX1_LOC_90/A NOR2X1_LOC_318/A 0.01fF
C27983 INVX1_LOC_47/A INVX1_LOC_26/Y 0.00fF
C27984 INVX1_LOC_10/A INVX1_LOC_23/A 0.31fF
C27985 NOR2X1_LOC_552/A INVX1_LOC_29/A 0.09fF
C27986 INVX1_LOC_152/A INVX1_LOC_280/A 0.01fF
C27987 NAND2X1_LOC_537/Y NAND2X1_LOC_326/a_36_24# 0.00fF
C27988 NAND2X1_LOC_538/Y NAND2X1_LOC_354/B 0.03fF
C27989 NOR2X1_LOC_561/Y INVX1_LOC_53/A 0.25fF
C27990 INVX1_LOC_36/A NOR2X1_LOC_68/A 0.17fF
C27991 NAND2X1_LOC_798/a_36_24# NAND2X1_LOC_350/A 0.00fF
C27992 INVX1_LOC_11/A NOR2X1_LOC_344/A 0.02fF
C27993 INVX1_LOC_73/Y NOR2X1_LOC_142/Y 0.39fF
C27994 INPUT_0 NOR2X1_LOC_38/B 0.28fF
C27995 INVX1_LOC_49/Y NAND2X1_LOC_655/B 0.01fF
C27996 NOR2X1_LOC_433/A NAND2X1_LOC_352/B 0.31fF
C27997 INVX1_LOC_21/A NAND2X1_LOC_850/Y 0.14fF
C27998 INVX1_LOC_52/Y INVX1_LOC_96/Y -0.01fF
C27999 INVX1_LOC_67/Y NOR2X1_LOC_334/Y 0.01fF
C28000 INVX1_LOC_64/A NOR2X1_LOC_521/Y 0.00fF
C28001 NOR2X1_LOC_703/Y INVX1_LOC_15/A 0.07fF
C28002 INVX1_LOC_42/Y INVX1_LOC_271/Y 0.01fF
C28003 NAND2X1_LOC_717/Y NAND2X1_LOC_705/Y 0.35fF
C28004 NOR2X1_LOC_155/A NOR2X1_LOC_499/B 0.00fF
C28005 NOR2X1_LOC_770/Y NOR2X1_LOC_383/B 0.01fF
C28006 NOR2X1_LOC_82/A NOR2X1_LOC_84/A 0.27fF
C28007 INVX1_LOC_35/A NAND2X1_LOC_573/A 0.00fF
C28008 NOR2X1_LOC_186/Y INVX1_LOC_208/Y 0.04fF
C28009 INVX1_LOC_166/A INVX1_LOC_175/Y 0.03fF
C28010 INVX1_LOC_2/A INVX1_LOC_1/A 0.08fF
C28011 NOR2X1_LOC_205/Y NOR2X1_LOC_423/Y 0.01fF
C28012 INVX1_LOC_135/A NOR2X1_LOC_416/a_36_216# 0.00fF
C28013 INVX1_LOC_255/Y NOR2X1_LOC_649/Y 0.06fF
C28014 NOR2X1_LOC_261/Y INVX1_LOC_89/A 0.07fF
C28015 INVX1_LOC_136/A INVX1_LOC_24/A 0.17fF
C28016 INVX1_LOC_11/A NAND2X1_LOC_357/B 0.24fF
C28017 NOR2X1_LOC_93/Y INVX1_LOC_316/Y 0.01fF
C28018 NOR2X1_LOC_722/Y NOR2X1_LOC_596/A 0.00fF
C28019 INVX1_LOC_25/A INPUT_1 0.44fF
C28020 NOR2X1_LOC_785/a_36_216# INVX1_LOC_26/Y 0.00fF
C28021 NOR2X1_LOC_272/Y INVX1_LOC_22/A 0.10fF
C28022 INVX1_LOC_161/Y NOR2X1_LOC_574/A 0.04fF
C28023 NOR2X1_LOC_226/A INVX1_LOC_1/A 0.13fF
C28024 INVX1_LOC_34/A NOR2X1_LOC_389/A 0.01fF
C28025 NAND2X1_LOC_573/Y INVX1_LOC_208/Y 0.08fF
C28026 INVX1_LOC_159/A NOR2X1_LOC_759/Y 0.01fF
C28027 INVX1_LOC_90/A NOR2X1_LOC_678/A 0.03fF
C28028 INVX1_LOC_34/A NAND2X1_LOC_199/B 0.04fF
C28029 NOR2X1_LOC_155/A NOR2X1_LOC_676/Y 0.01fF
C28030 NOR2X1_LOC_222/Y NOR2X1_LOC_205/Y 0.16fF
C28031 NOR2X1_LOC_356/A INVX1_LOC_58/Y 0.01fF
C28032 NOR2X1_LOC_469/a_36_216# NAND2X1_LOC_850/Y 0.00fF
C28033 INVX1_LOC_108/Y NAND2X1_LOC_508/A 0.16fF
C28034 NOR2X1_LOC_235/a_36_216# INVX1_LOC_25/Y 0.00fF
C28035 NOR2X1_LOC_332/A INVX1_LOC_50/Y 0.07fF
C28036 INVX1_LOC_206/A INVX1_LOC_292/A 0.07fF
C28037 NAND2X1_LOC_303/Y INVX1_LOC_16/A 0.10fF
C28038 INVX1_LOC_269/A INVX1_LOC_316/Y 0.01fF
C28039 VDD NAND2X1_LOC_206/B 0.08fF
C28040 INVX1_LOC_136/A NOR2X1_LOC_557/Y 0.28fF
C28041 NOR2X1_LOC_536/A INVX1_LOC_264/A 0.02fF
C28042 NOR2X1_LOC_454/Y NOR2X1_LOC_583/a_36_216# 0.01fF
C28043 NOR2X1_LOC_813/Y INVX1_LOC_29/A 0.07fF
C28044 NOR2X1_LOC_590/A NOR2X1_LOC_709/A 0.03fF
C28045 INVX1_LOC_14/A INVX1_LOC_53/Y 0.02fF
C28046 NOR2X1_LOC_68/A NOR2X1_LOC_804/B 0.10fF
C28047 NOR2X1_LOC_778/A INVX1_LOC_33/A 0.17fF
C28048 INVX1_LOC_41/A NOR2X1_LOC_703/B 0.03fF
C28049 NAND2X1_LOC_326/A NAND2X1_LOC_660/Y 0.03fF
C28050 NOR2X1_LOC_15/Y NOR2X1_LOC_188/a_36_216# 0.01fF
C28051 NOR2X1_LOC_489/A NOR2X1_LOC_814/A 0.03fF
C28052 INVX1_LOC_20/A INVX1_LOC_19/Y 0.27fF
C28053 INVX1_LOC_5/A NOR2X1_LOC_156/A 0.06fF
C28054 INVX1_LOC_280/A INVX1_LOC_29/A 0.11fF
C28055 INVX1_LOC_27/A INVX1_LOC_120/A 2.09fF
C28056 INVX1_LOC_223/Y NOR2X1_LOC_542/Y 0.00fF
C28057 NOR2X1_LOC_328/Y NAND2X1_LOC_227/Y 0.01fF
C28058 INVX1_LOC_208/A NOR2X1_LOC_160/B 0.07fF
C28059 NOR2X1_LOC_316/Y INVX1_LOC_72/A 0.09fF
C28060 INVX1_LOC_34/A NOR2X1_LOC_596/A 0.06fF
C28061 D_INPUT_0 NAND2X1_LOC_326/A 0.08fF
C28062 NOR2X1_LOC_835/B INVX1_LOC_53/A 0.02fF
C28063 INVX1_LOC_152/Y NOR2X1_LOC_97/A 0.22fF
C28064 NOR2X1_LOC_516/B NOR2X1_LOC_160/B 0.13fF
C28065 NOR2X1_LOC_381/Y NOR2X1_LOC_332/A 0.05fF
C28066 INVX1_LOC_2/A NOR2X1_LOC_384/Y 0.41fF
C28067 NOR2X1_LOC_67/A INVX1_LOC_30/A 0.19fF
C28068 NOR2X1_LOC_78/B NOR2X1_LOC_169/B 0.04fF
C28069 INVX1_LOC_226/Y INVX1_LOC_31/A 0.03fF
C28070 INVX1_LOC_136/A INVX1_LOC_143/A 0.10fF
C28071 NOR2X1_LOC_374/A NOR2X1_LOC_551/B 0.01fF
C28072 INVX1_LOC_35/A INVX1_LOC_285/Y 0.01fF
C28073 NAND2X1_LOC_659/A NAND2X1_LOC_657/a_36_24# 0.01fF
C28074 NOR2X1_LOC_41/Y INVX1_LOC_159/A 0.01fF
C28075 NOR2X1_LOC_456/Y NOR2X1_LOC_337/Y 0.01fF
C28076 INVX1_LOC_294/A INVX1_LOC_285/A 0.01fF
C28077 INVX1_LOC_78/A NAND2X1_LOC_287/B 0.68fF
C28078 NOR2X1_LOC_593/Y NOR2X1_LOC_344/A 0.03fF
C28079 INVX1_LOC_1/A INPUT_1 0.48fF
C28080 NOR2X1_LOC_374/A NOR2X1_LOC_704/a_36_216# 0.00fF
C28081 NOR2X1_LOC_335/A NOR2X1_LOC_392/B 0.01fF
C28082 INVX1_LOC_269/A NOR2X1_LOC_395/a_36_216# 0.00fF
C28083 NOR2X1_LOC_111/Y NOR2X1_LOC_321/Y 0.09fF
C28084 NOR2X1_LOC_336/B INVX1_LOC_22/A 0.00fF
C28085 NAND2X1_LOC_357/B NOR2X1_LOC_433/A 0.39fF
C28086 NOR2X1_LOC_598/B NOR2X1_LOC_45/B 0.03fF
C28087 NAND2X1_LOC_303/Y INVX1_LOC_28/A 0.30fF
C28088 INVX1_LOC_298/Y INVX1_LOC_139/Y 0.03fF
C28089 INVX1_LOC_136/A NAND2X1_LOC_565/B 0.01fF
C28090 NOR2X1_LOC_647/A INVX1_LOC_2/Y 0.01fF
C28091 NAND2X1_LOC_722/A NOR2X1_LOC_753/Y 0.15fF
C28092 INVX1_LOC_72/A NAND2X1_LOC_662/Y 0.07fF
C28093 NAND2X1_LOC_364/A INVX1_LOC_22/A 0.17fF
C28094 INVX1_LOC_299/A NOR2X1_LOC_567/B 0.04fF
C28095 NOR2X1_LOC_792/B INVX1_LOC_162/A 0.04fF
C28096 NAND2X1_LOC_725/A NOR2X1_LOC_45/B 0.05fF
C28097 INVX1_LOC_135/A NOR2X1_LOC_703/a_36_216# 0.01fF
C28098 NAND2X1_LOC_538/a_36_24# NAND2X1_LOC_326/A 0.01fF
C28099 NAND2X1_LOC_440/a_36_24# INVX1_LOC_271/A 0.00fF
C28100 NOR2X1_LOC_392/a_36_216# INVX1_LOC_306/Y 0.01fF
C28101 INVX1_LOC_35/A INVX1_LOC_65/A 0.12fF
C28102 INVX1_LOC_5/A INVX1_LOC_96/A 0.03fF
C28103 NOR2X1_LOC_598/B INVX1_LOC_199/Y 0.02fF
C28104 INVX1_LOC_88/A INVX1_LOC_73/A 0.04fF
C28105 INVX1_LOC_6/A NAND2X1_LOC_474/Y 0.09fF
C28106 INVX1_LOC_63/Y INVX1_LOC_96/Y 0.02fF
C28107 INVX1_LOC_37/A NOR2X1_LOC_383/B 0.15fF
C28108 NOR2X1_LOC_286/a_36_216# NOR2X1_LOC_78/A 0.00fF
C28109 INVX1_LOC_121/Y INVX1_LOC_257/Y 1.22fF
C28110 NAND2X1_LOC_357/B NOR2X1_LOC_52/B 0.07fF
C28111 NOR2X1_LOC_216/B NOR2X1_LOC_116/a_36_216# 0.01fF
C28112 NAND2X1_LOC_564/B INVX1_LOC_41/Y 0.45fF
C28113 NOR2X1_LOC_468/Y INPUT_0 0.53fF
C28114 NOR2X1_LOC_690/A NAND2X1_LOC_717/Y 0.04fF
C28115 INVX1_LOC_45/A NOR2X1_LOC_333/A 0.01fF
C28116 NOR2X1_LOC_620/B INVX1_LOC_33/A 0.03fF
C28117 INVX1_LOC_7/Y INVX1_LOC_91/A 0.01fF
C28118 INVX1_LOC_53/A INVX1_LOC_76/A 0.69fF
C28119 NAND2X1_LOC_563/Y NOR2X1_LOC_515/a_36_216# 0.01fF
C28120 INVX1_LOC_178/Y INVX1_LOC_23/A 0.01fF
C28121 INVX1_LOC_136/A NAND2X1_LOC_800/Y 0.03fF
C28122 NOR2X1_LOC_92/Y INVX1_LOC_309/A 0.03fF
C28123 INVX1_LOC_136/A NOR2X1_LOC_130/A 0.13fF
C28124 INVX1_LOC_5/A NOR2X1_LOC_124/A 0.00fF
C28125 INVX1_LOC_64/A NOR2X1_LOC_670/Y 0.00fF
C28126 INVX1_LOC_38/A NOR2X1_LOC_318/A 0.03fF
C28127 INVX1_LOC_278/A NAND2X1_LOC_244/A 0.02fF
C28128 INVX1_LOC_50/A INVX1_LOC_33/Y 0.03fF
C28129 NOR2X1_LOC_825/Y NOR2X1_LOC_392/Y 0.02fF
C28130 INVX1_LOC_34/A NOR2X1_LOC_399/Y 0.06fF
C28131 NAND2X1_LOC_260/a_36_24# INVX1_LOC_78/A 0.00fF
C28132 NOR2X1_LOC_456/Y VDD 0.22fF
C28133 NOR2X1_LOC_52/B NAND2X1_LOC_655/a_36_24# 0.00fF
C28134 INVX1_LOC_245/Y NOR2X1_LOC_74/a_36_216# 0.00fF
C28135 NOR2X1_LOC_432/a_36_216# INVX1_LOC_266/Y 0.00fF
C28136 NOR2X1_LOC_216/Y NOR2X1_LOC_276/Y 0.00fF
C28137 INVX1_LOC_223/A INVX1_LOC_313/Y 0.00fF
C28138 NOR2X1_LOC_226/A INVX1_LOC_221/A 0.01fF
C28139 NOR2X1_LOC_75/Y NOR2X1_LOC_74/A 0.03fF
C28140 NOR2X1_LOC_78/B NOR2X1_LOC_367/B 0.46fF
C28141 NOR2X1_LOC_210/A INVX1_LOC_113/Y 0.01fF
C28142 NOR2X1_LOC_384/Y INPUT_1 0.57fF
C28143 NAND2X1_LOC_454/Y NOR2X1_LOC_435/A 0.04fF
C28144 NOR2X1_LOC_114/a_36_216# INVX1_LOC_270/A 0.00fF
C28145 NAND2X1_LOC_773/Y INVX1_LOC_125/Y 0.05fF
C28146 NOR2X1_LOC_92/Y INVX1_LOC_91/A 0.22fF
C28147 INVX1_LOC_89/A NOR2X1_LOC_168/Y 0.01fF
C28148 GATE_741 INVX1_LOC_11/Y 0.33fF
C28149 INVX1_LOC_164/Y INVX1_LOC_168/A 0.00fF
C28150 NOR2X1_LOC_690/A INVX1_LOC_16/A 0.02fF
C28151 INVX1_LOC_135/A INVX1_LOC_228/A 0.23fF
C28152 INVX1_LOC_163/Y NAND2X1_LOC_402/a_36_24# 0.00fF
C28153 NOR2X1_LOC_155/A NOR2X1_LOC_465/Y 0.00fF
C28154 NAND2X1_LOC_53/Y INVX1_LOC_6/A 0.24fF
C28155 NAND2X1_LOC_745/a_36_24# INVX1_LOC_91/A 0.01fF
C28156 NAND2X1_LOC_79/a_36_24# NOR2X1_LOC_719/B 0.00fF
C28157 INVX1_LOC_45/A NOR2X1_LOC_289/Y 0.03fF
C28158 INVX1_LOC_24/A NAND2X1_LOC_862/Y 0.07fF
C28159 NAND2X1_LOC_714/B NOR2X1_LOC_56/Y 0.01fF
C28160 INVX1_LOC_178/A NAND2X1_LOC_658/a_36_24# 0.00fF
C28161 NOR2X1_LOC_92/Y INVX1_LOC_11/Y 0.46fF
C28162 NAND2X1_LOC_633/Y INVX1_LOC_306/Y 0.02fF
C28163 NOR2X1_LOC_262/Y INVX1_LOC_89/A 0.03fF
C28164 NOR2X1_LOC_78/B INVX1_LOC_179/Y 0.01fF
C28165 NOR2X1_LOC_667/A NAND2X1_LOC_850/Y 0.02fF
C28166 NOR2X1_LOC_447/A INVX1_LOC_92/A 0.03fF
C28167 NOR2X1_LOC_82/Y NOR2X1_LOC_709/A 0.03fF
C28168 INVX1_LOC_258/Y INVX1_LOC_20/A 0.14fF
C28169 NOR2X1_LOC_629/a_36_216# NAND2X1_LOC_735/B 0.00fF
C28170 NOR2X1_LOC_416/a_36_216# INVX1_LOC_280/A 0.01fF
C28171 INVX1_LOC_38/A NOR2X1_LOC_678/A 0.03fF
C28172 INVX1_LOC_290/Y NOR2X1_LOC_755/Y 0.06fF
C28173 NOR2X1_LOC_553/B INVX1_LOC_104/A 0.00fF
C28174 INVX1_LOC_34/A NAND2X1_LOC_795/Y 0.12fF
C28175 NAND2X1_LOC_9/Y INVX1_LOC_9/A 0.41fF
C28176 INVX1_LOC_36/A NOR2X1_LOC_2/Y 0.01fF
C28177 INVX1_LOC_38/A INVX1_LOC_295/Y 0.04fF
C28178 NOR2X1_LOC_829/A NAND2X1_LOC_770/Y 0.03fF
C28179 NOR2X1_LOC_231/a_36_216# NOR2X1_LOC_9/Y 0.00fF
C28180 NOR2X1_LOC_92/Y NOR2X1_LOC_421/Y 0.09fF
C28181 NAND2X1_LOC_714/B VDD 0.16fF
C28182 NOR2X1_LOC_84/B NOR2X1_LOC_38/B 0.00fF
C28183 INVX1_LOC_268/Y NAND2X1_LOC_451/Y 0.03fF
C28184 NAND2X1_LOC_11/Y INVX1_LOC_22/A 0.00fF
C28185 NOR2X1_LOC_6/B NOR2X1_LOC_332/A 0.02fF
C28186 INVX1_LOC_279/A INVX1_LOC_266/Y 0.10fF
C28187 NAND2X1_LOC_714/B NAND2X1_LOC_800/A 0.03fF
C28188 NAND2X1_LOC_563/A INVX1_LOC_316/Y 0.11fF
C28189 NOR2X1_LOC_205/Y NOR2X1_LOC_69/A 0.01fF
C28190 NOR2X1_LOC_763/A INVX1_LOC_37/A 0.07fF
C28191 INVX1_LOC_23/A INVX1_LOC_307/A 0.09fF
C28192 INVX1_LOC_103/A NOR2X1_LOC_314/a_36_216# 0.02fF
C28193 NOR2X1_LOC_609/A NOR2X1_LOC_74/A 0.03fF
C28194 NOR2X1_LOC_623/B INVX1_LOC_69/A 0.01fF
C28195 INVX1_LOC_271/Y INVX1_LOC_19/A 0.17fF
C28196 INVX1_LOC_224/Y INVX1_LOC_123/Y 0.02fF
C28197 NOR2X1_LOC_307/A NOR2X1_LOC_209/A 0.02fF
C28198 NOR2X1_LOC_92/Y NOR2X1_LOC_653/a_36_216# 0.03fF
C28199 NAND2X1_LOC_361/Y NOR2X1_LOC_775/Y 0.01fF
C28200 INVX1_LOC_23/A NOR2X1_LOC_445/B 0.41fF
C28201 NOR2X1_LOC_650/a_36_216# INVX1_LOC_58/Y 0.01fF
C28202 NAND2X1_LOC_561/B VDD 0.03fF
C28203 NOR2X1_LOC_78/B NOR2X1_LOC_561/Y 0.07fF
C28204 NAND2X1_LOC_344/a_36_24# INVX1_LOC_280/A 0.01fF
C28205 INVX1_LOC_1/A NAND2X1_LOC_605/a_36_24# 0.00fF
C28206 NOR2X1_LOC_598/B NOR2X1_LOC_862/B 0.21fF
C28207 NOR2X1_LOC_78/B INVX1_LOC_7/A 0.07fF
C28208 INVX1_LOC_247/Y NOR2X1_LOC_794/A 0.16fF
C28209 NOR2X1_LOC_690/A INVX1_LOC_28/A 0.03fF
C28210 NOR2X1_LOC_589/A NOR2X1_LOC_131/Y 0.05fF
C28211 NOR2X1_LOC_798/A INVX1_LOC_9/A 0.10fF
C28212 NAND2X1_LOC_510/A NOR2X1_LOC_78/A 0.04fF
C28213 NOR2X1_LOC_725/A NOR2X1_LOC_707/B 0.22fF
C28214 INVX1_LOC_243/A INVX1_LOC_83/A 0.01fF
C28215 NAND2X1_LOC_564/B NAND2X1_LOC_861/a_36_24# 0.01fF
C28216 NOR2X1_LOC_576/B NAND2X1_LOC_839/A 0.52fF
C28217 NOR2X1_LOC_671/Y NOR2X1_LOC_825/a_36_216# 0.00fF
C28218 NAND2X1_LOC_326/A NAND2X1_LOC_848/A 0.10fF
C28219 NAND2X1_LOC_837/Y INVX1_LOC_309/A 0.00fF
C28220 NOR2X1_LOC_375/Y NOR2X1_LOC_459/A 0.01fF
C28221 NOR2X1_LOC_445/Y INVX1_LOC_75/A 0.05fF
C28222 INVX1_LOC_124/A NAND2X1_LOC_842/B 0.26fF
C28223 INVX1_LOC_49/A NOR2X1_LOC_188/A 0.03fF
C28224 NOR2X1_LOC_414/Y NAND2X1_LOC_206/Y 0.04fF
C28225 NOR2X1_LOC_405/A NOR2X1_LOC_274/B 0.12fF
C28226 INVX1_LOC_88/A NOR2X1_LOC_122/a_36_216# 0.00fF
C28227 NOR2X1_LOC_419/Y NOR2X1_LOC_9/Y 0.01fF
C28228 INVX1_LOC_290/A INPUT_5 0.03fF
C28229 NOR2X1_LOC_36/B INVX1_LOC_296/A 0.13fF
C28230 NOR2X1_LOC_52/B NAND2X1_LOC_849/A 0.06fF
C28231 NOR2X1_LOC_91/A INVX1_LOC_12/A 0.13fF
C28232 NOR2X1_LOC_716/B NOR2X1_LOC_9/Y 0.23fF
C28233 NOR2X1_LOC_392/Y INVX1_LOC_84/A 0.22fF
C28234 INVX1_LOC_182/Y INVX1_LOC_266/Y 0.03fF
C28235 NAND2X1_LOC_839/Y NAND2X1_LOC_560/A 0.01fF
C28236 NAND2X1_LOC_837/Y INVX1_LOC_91/A 0.07fF
C28237 NOR2X1_LOC_91/A NOR2X1_LOC_519/Y 0.03fF
C28238 INVX1_LOC_1/A INVX1_LOC_118/A 0.10fF
C28239 INVX1_LOC_215/A NAND2X1_LOC_656/Y 0.50fF
C28240 INVX1_LOC_111/Y NAND2X1_LOC_369/a_36_24# 0.01fF
C28241 INVX1_LOC_304/Y NOR2X1_LOC_716/a_36_216# 0.00fF
C28242 INVX1_LOC_41/A NOR2X1_LOC_728/B 0.00fF
C28243 NAND2X1_LOC_11/a_36_24# INVX1_LOC_140/A 0.05fF
C28244 NOR2X1_LOC_337/Y NOR2X1_LOC_550/B 0.18fF
C28245 INVX1_LOC_25/A NAND2X1_LOC_63/Y 0.03fF
C28246 NOR2X1_LOC_844/A INPUT_0 0.03fF
C28247 NOR2X1_LOC_561/Y INVX1_LOC_83/A 0.10fF
C28248 INVX1_LOC_11/Y NAND2X1_LOC_837/Y 0.07fF
C28249 INVX1_LOC_7/A INVX1_LOC_83/A 0.05fF
C28250 INVX1_LOC_57/Y INVX1_LOC_37/A 0.07fF
C28251 INVX1_LOC_12/A INVX1_LOC_23/A 0.44fF
C28252 INVX1_LOC_49/A NOR2X1_LOC_43/Y 0.08fF
C28253 INVX1_LOC_41/A INVX1_LOC_91/A 0.11fF
C28254 NOR2X1_LOC_577/Y NOR2X1_LOC_405/A 0.08fF
C28255 INVX1_LOC_98/Y NOR2X1_LOC_74/A 0.10fF
C28256 INVX1_LOC_2/A NOR2X1_LOC_188/A 0.07fF
C28257 INVX1_LOC_313/A INVX1_LOC_10/A 0.07fF
C28258 INVX1_LOC_27/A NAND2X1_LOC_659/A 0.04fF
C28259 INVX1_LOC_299/A NOR2X1_LOC_79/Y 0.00fF
C28260 NOR2X1_LOC_731/a_36_216# INVX1_LOC_117/A 0.00fF
C28261 NOR2X1_LOC_158/Y NAND2X1_LOC_470/B 0.03fF
C28262 INVX1_LOC_18/A NOR2X1_LOC_111/A 0.07fF
C28263 NOR2X1_LOC_78/B NOR2X1_LOC_835/B 0.01fF
C28264 INVX1_LOC_300/Y VDD 0.28fF
C28265 NOR2X1_LOC_273/Y VDD 0.61fF
C28266 INVX1_LOC_136/A NAND2X1_LOC_811/B 0.18fF
C28267 NOR2X1_LOC_759/Y NOR2X1_LOC_69/a_36_216# 0.00fF
C28268 NOR2X1_LOC_759/Y VDD 0.58fF
C28269 NOR2X1_LOC_173/a_36_216# NAND2X1_LOC_593/Y 0.01fF
C28270 NOR2X1_LOC_91/Y NOR2X1_LOC_176/Y 0.00fF
C28271 NOR2X1_LOC_498/Y INVX1_LOC_11/Y 0.07fF
C28272 INVX1_LOC_83/A NOR2X1_LOC_708/Y 0.03fF
C28273 NAND2X1_LOC_303/B INVX1_LOC_173/Y 0.02fF
C28274 NOR2X1_LOC_679/a_36_216# NAND2X1_LOC_802/Y 0.00fF
C28275 NOR2X1_LOC_798/A NOR2X1_LOC_691/a_36_216# 0.00fF
C28276 NAND2X1_LOC_361/Y NAND2X1_LOC_447/Y 0.01fF
C28277 NAND2X1_LOC_477/A INVX1_LOC_91/A 0.11fF
C28278 INVX1_LOC_202/A VDD 0.50fF
C28279 NOR2X1_LOC_577/Y NOR2X1_LOC_682/a_36_216# 0.00fF
C28280 NOR2X1_LOC_387/A NAND2X1_LOC_852/Y 0.05fF
C28281 NOR2X1_LOC_78/A NOR2X1_LOC_174/a_36_216# 0.02fF
C28282 NOR2X1_LOC_406/a_36_216# NOR2X1_LOC_89/A 0.00fF
C28283 INVX1_LOC_141/Y INVX1_LOC_54/A 2.72fF
C28284 INVX1_LOC_41/Y NAND2X1_LOC_804/Y 0.04fF
C28285 NOR2X1_LOC_398/Y INVX1_LOC_91/A 0.01fF
C28286 NOR2X1_LOC_92/Y INVX1_LOC_203/A 0.10fF
C28287 NOR2X1_LOC_717/B NAND2X1_LOC_472/a_36_24# 0.00fF
C28288 NOR2X1_LOC_256/a_36_216# NOR2X1_LOC_813/Y 0.01fF
C28289 NOR2X1_LOC_84/A INVX1_LOC_59/Y 0.03fF
C28290 NOR2X1_LOC_550/B VDD 1.76fF
C28291 NOR2X1_LOC_68/A NOR2X1_LOC_865/A 0.03fF
C28292 INVX1_LOC_308/Y INVX1_LOC_285/A 0.04fF
C28293 INVX1_LOC_312/Y INVX1_LOC_54/A 0.07fF
C28294 NAND2X1_LOC_149/Y INVX1_LOC_262/Y 0.05fF
C28295 NOR2X1_LOC_78/A NOR2X1_LOC_131/A 0.01fF
C28296 NOR2X1_LOC_392/Y INVX1_LOC_15/A 0.07fF
C28297 INVX1_LOC_269/A NOR2X1_LOC_662/A 0.47fF
C28298 NOR2X1_LOC_638/a_36_216# INVX1_LOC_77/Y -0.01fF
C28299 NOR2X1_LOC_232/Y NOR2X1_LOC_662/A 0.01fF
C28300 NAND2X1_LOC_773/Y INVX1_LOC_19/A 0.03fF
C28301 INVX1_LOC_26/A INVX1_LOC_181/A 0.31fF
C28302 INVX1_LOC_155/A INVX1_LOC_12/Y 0.01fF
C28303 INVX1_LOC_34/A NAND2X1_LOC_212/a_36_24# 0.00fF
C28304 NOR2X1_LOC_717/B NOR2X1_LOC_74/A 0.03fF
C28305 NOR2X1_LOC_516/B INVX1_LOC_315/Y 1.14fF
C28306 INVX1_LOC_1/A NAND2X1_LOC_63/Y 0.10fF
C28307 INVX1_LOC_43/A NAND2X1_LOC_642/Y 0.03fF
C28308 INVX1_LOC_35/A INVX1_LOC_4/Y 0.03fF
C28309 NAND2X1_LOC_860/A INVX1_LOC_87/A 0.01fF
C28310 NOR2X1_LOC_742/A INVX1_LOC_85/Y 0.13fF
C28311 INVX1_LOC_10/A INVX1_LOC_6/A 8.16fF
C28312 NOR2X1_LOC_52/Y NOR2X1_LOC_155/A 0.50fF
C28313 NAND2X1_LOC_710/a_36_24# INVX1_LOC_118/A 0.00fF
C28314 NOR2X1_LOC_113/B NOR2X1_LOC_137/A 0.00fF
C28315 NOR2X1_LOC_813/Y INVX1_LOC_8/A 0.08fF
C28316 INVX1_LOC_171/A INVX1_LOC_222/A 0.06fF
C28317 NOR2X1_LOC_405/A INVX1_LOC_22/A 0.15fF
C28318 INVX1_LOC_83/A NAND2X1_LOC_251/a_36_24# 0.00fF
C28319 NOR2X1_LOC_270/Y NOR2X1_LOC_155/A 0.58fF
C28320 NOR2X1_LOC_78/B INVX1_LOC_76/A 0.31fF
C28321 NAND2X1_LOC_555/Y NAND2X1_LOC_225/a_36_24# 0.01fF
C28322 NOR2X1_LOC_41/Y VDD 0.12fF
C28323 INVX1_LOC_216/A D_INPUT_3 0.05fF
C28324 INVX1_LOC_22/A NAND2X1_LOC_422/a_36_24# 0.00fF
C28325 NOR2X1_LOC_677/Y INVX1_LOC_271/A 0.11fF
C28326 INVX1_LOC_121/A INVX1_LOC_91/A 0.01fF
C28327 INVX1_LOC_8/A INVX1_LOC_280/A 0.11fF
C28328 INVX1_LOC_71/A INVX1_LOC_70/A 0.01fF
C28329 INVX1_LOC_53/A NOR2X1_LOC_447/A 0.00fF
C28330 NOR2X1_LOC_68/A NAND2X1_LOC_609/a_36_24# 0.00fF
C28331 INVX1_LOC_89/A INVX1_LOC_123/A 0.10fF
C28332 NOR2X1_LOC_219/B INVX1_LOC_54/A 0.01fF
C28333 INVX1_LOC_91/Y NAND2X1_LOC_560/A 0.01fF
C28334 INVX1_LOC_134/Y INVX1_LOC_117/A 0.02fF
C28335 NAND2X1_LOC_72/Y NAND2X1_LOC_72/a_36_24# 0.03fF
C28336 INVX1_LOC_208/A NAND2X1_LOC_211/Y 0.19fF
C28337 NAND2X1_LOC_793/B NAND2X1_LOC_439/a_36_24# 0.01fF
C28338 INVX1_LOC_297/Y VDD -0.00fF
C28339 NOR2X1_LOC_210/a_36_216# NOR2X1_LOC_467/A -0.00fF
C28340 NAND2X1_LOC_787/A NAND2X1_LOC_787/Y 0.01fF
C28341 INVX1_LOC_236/A NOR2X1_LOC_536/A 0.06fF
C28342 NOR2X1_LOC_151/Y NOR2X1_LOC_74/A 0.10fF
C28343 INVX1_LOC_316/Y NOR2X1_LOC_37/a_36_216# 0.02fF
C28344 INVX1_LOC_22/A NOR2X1_LOC_857/A 0.01fF
C28345 INVX1_LOC_178/A INVX1_LOC_273/A 0.05fF
C28346 NOR2X1_LOC_78/B NAND2X1_LOC_418/a_36_24# 0.00fF
C28347 INVX1_LOC_75/A NOR2X1_LOC_335/B 0.03fF
C28348 NOR2X1_LOC_788/a_36_216# NOR2X1_LOC_564/Y 0.00fF
C28349 NOR2X1_LOC_299/Y INVX1_LOC_11/Y 3.02fF
C28350 NOR2X1_LOC_544/A INVX1_LOC_117/A 0.07fF
C28351 NOR2X1_LOC_68/A INVX1_LOC_63/A 0.24fF
C28352 INVX1_LOC_31/A INVX1_LOC_12/A 0.09fF
C28353 INVX1_LOC_1/A NAND2X1_LOC_618/Y 0.07fF
C28354 NOR2X1_LOC_419/Y NOR2X1_LOC_243/B 0.00fF
C28355 NAND2X1_LOC_110/a_36_24# NAND2X1_LOC_96/A 0.00fF
C28356 NOR2X1_LOC_455/Y INVX1_LOC_53/A -0.03fF
C28357 NAND2X1_LOC_568/A INVX1_LOC_231/A 0.04fF
C28358 INVX1_LOC_229/Y INVX1_LOC_20/A 0.08fF
C28359 NAND2X1_LOC_361/Y NAND2X1_LOC_750/a_36_24# 0.00fF
C28360 INVX1_LOC_266/A INVX1_LOC_78/A 0.07fF
C28361 NOR2X1_LOC_348/a_36_216# INVX1_LOC_290/Y 0.01fF
C28362 NOR2X1_LOC_561/Y INVX1_LOC_46/A 2.99fF
C28363 NOR2X1_LOC_791/a_36_216# NAND2X1_LOC_773/B 0.01fF
C28364 INVX1_LOC_43/A NOR2X1_LOC_271/Y 0.25fF
C28365 INVX1_LOC_83/A INVX1_LOC_76/A 0.50fF
C28366 INVX1_LOC_40/A NOR2X1_LOC_99/a_36_216# 0.00fF
C28367 NOR2X1_LOC_45/B NAND2X1_LOC_560/A 0.03fF
C28368 INVX1_LOC_141/Y NOR2X1_LOC_48/B 0.71fF
C28369 NOR2X1_LOC_372/a_36_216# NAND2X1_LOC_254/Y 0.00fF
C28370 NOR2X1_LOC_180/Y NOR2X1_LOC_155/A 0.01fF
C28371 NOR2X1_LOC_795/Y NOR2X1_LOC_634/A 0.57fF
C28372 INVX1_LOC_1/A NOR2X1_LOC_631/Y 0.20fF
C28373 INVX1_LOC_159/A NAND2X1_LOC_74/B 0.00fF
C28374 NAND2X1_LOC_474/Y INVX1_LOC_270/A 0.00fF
C28375 INVX1_LOC_13/A NOR2X1_LOC_536/A 0.03fF
C28376 NOR2X1_LOC_434/Y INVX1_LOC_53/A 0.01fF
C28377 INVX1_LOC_72/A INVX1_LOC_290/Y 0.07fF
C28378 INVX1_LOC_25/A INVX1_LOC_39/A 0.06fF
C28379 INVX1_LOC_212/A NOR2X1_LOC_340/A 0.06fF
C28380 NAND2X1_LOC_360/B INVX1_LOC_46/Y 0.02fF
C28381 NOR2X1_LOC_816/A INVX1_LOC_273/A 0.12fF
C28382 INVX1_LOC_201/Y INVX1_LOC_203/A 0.18fF
C28383 NOR2X1_LOC_261/a_36_216# NAND2X1_LOC_149/Y 0.01fF
C28384 INVX1_LOC_21/A INPUT_6 0.01fF
C28385 NOR2X1_LOC_590/A NOR2X1_LOC_334/Y 0.09fF
C28386 NOR2X1_LOC_597/A NAND2X1_LOC_453/A 0.01fF
C28387 INVX1_LOC_141/A INVX1_LOC_94/Y 0.07fF
C28388 NOR2X1_LOC_458/B NOR2X1_LOC_155/A 0.00fF
C28389 NOR2X1_LOC_288/A NOR2X1_LOC_691/A 0.06fF
C28390 INVX1_LOC_11/A NOR2X1_LOC_282/Y 0.01fF
C28391 NOR2X1_LOC_91/A INVX1_LOC_200/A 0.01fF
C28392 INVX1_LOC_229/A NAND2X1_LOC_725/Y 0.03fF
C28393 INVX1_LOC_13/A NOR2X1_LOC_655/Y 0.30fF
C28394 NAND2X1_LOC_755/a_36_24# INVX1_LOC_84/A 0.00fF
C28395 INVX1_LOC_269/A INVX1_LOC_57/A 0.23fF
C28396 NOR2X1_LOC_667/Y NAND2X1_LOC_175/Y 0.05fF
C28397 NOR2X1_LOC_246/A NOR2X1_LOC_536/A 0.02fF
C28398 NAND2X1_LOC_35/Y NAND2X1_LOC_391/Y 0.07fF
C28399 INVX1_LOC_13/A NAND2X1_LOC_93/B 0.01fF
C28400 NOR2X1_LOC_86/A NOR2X1_LOC_88/A 0.01fF
C28401 NAND2X1_LOC_551/A NOR2X1_LOC_536/A 0.19fF
C28402 NOR2X1_LOC_163/Y INVX1_LOC_37/A 0.03fF
C28403 NAND2X1_LOC_656/Y INVX1_LOC_54/A 0.07fF
C28404 INVX1_LOC_31/A NOR2X1_LOC_686/A 0.00fF
C28405 INVX1_LOC_72/Y NOR2X1_LOC_38/B 0.04fF
C28406 NOR2X1_LOC_91/A NAND2X1_LOC_733/Y 0.22fF
C28407 NAND2X1_LOC_796/B NOR2X1_LOC_406/A 0.41fF
C28408 NOR2X1_LOC_627/Y INVX1_LOC_186/Y 0.01fF
C28409 NAND2X1_LOC_794/B NAND2X1_LOC_788/a_36_24# 0.02fF
C28410 NOR2X1_LOC_74/Y INVX1_LOC_37/A 0.02fF
C28411 NAND2X1_LOC_779/a_36_24# INVX1_LOC_291/A 0.01fF
C28412 NAND2X1_LOC_860/A NOR2X1_LOC_82/A 0.27fF
C28413 NOR2X1_LOC_15/Y NAND2X1_LOC_552/A 0.02fF
C28414 INVX1_LOC_64/A NOR2X1_LOC_523/A 0.02fF
C28415 NOR2X1_LOC_15/Y INVX1_LOC_5/A 0.10fF
C28416 NOR2X1_LOC_606/Y NOR2X1_LOC_646/B 0.06fF
C28417 NAND2X1_LOC_141/A NAND2X1_LOC_83/a_36_24# 0.00fF
C28418 NAND2X1_LOC_809/A NAND2X1_LOC_802/Y 0.04fF
C28419 NOR2X1_LOC_6/B INVX1_LOC_42/A 1.17fF
C28420 INVX1_LOC_13/A NOR2X1_LOC_649/B 0.07fF
C28421 NOR2X1_LOC_781/Y NOR2X1_LOC_158/Y 0.04fF
C28422 INVX1_LOC_135/A NAND2X1_LOC_244/a_36_24# 0.06fF
C28423 NOR2X1_LOC_334/A VDD 0.33fF
C28424 NOR2X1_LOC_289/Y NOR2X1_LOC_331/B 0.04fF
C28425 INVX1_LOC_13/A INVX1_LOC_3/A 0.47fF
C28426 INVX1_LOC_50/A NAND2X1_LOC_741/B 0.05fF
C28427 NOR2X1_LOC_91/A INVX1_LOC_217/A 0.10fF
C28428 NOR2X1_LOC_311/a_36_216# INVX1_LOC_20/A 0.01fF
C28429 INVX1_LOC_10/A NOR2X1_LOC_117/Y 0.01fF
C28430 INVX1_LOC_39/A INVX1_LOC_1/A 0.03fF
C28431 NAND2X1_LOC_753/a_36_24# INVX1_LOC_292/A 0.00fF
C28432 NAND2X1_LOC_364/A NOR2X1_LOC_843/B 0.01fF
C28433 NOR2X1_LOC_15/Y INVX1_LOC_178/A 0.12fF
C28434 INVX1_LOC_234/Y INVX1_LOC_237/A 0.11fF
C28435 D_INPUT_0 NAND2X1_LOC_572/B 0.01fF
C28436 INVX1_LOC_235/Y INVX1_LOC_14/A 0.19fF
C28437 NOR2X1_LOC_732/a_36_216# NOR2X1_LOC_155/A 0.01fF
C28438 NOR2X1_LOC_398/a_36_216# INVX1_LOC_3/Y 0.00fF
C28439 NOR2X1_LOC_709/B NOR2X1_LOC_74/A 0.02fF
C28440 NOR2X1_LOC_516/B NAND2X1_LOC_207/B 0.02fF
C28441 INVX1_LOC_217/A INVX1_LOC_23/A 0.00fF
C28442 NAND2X1_LOC_824/a_36_24# NOR2X1_LOC_865/Y 0.01fF
C28443 INVX1_LOC_269/A NOR2X1_LOC_475/A 0.01fF
C28444 INVX1_LOC_279/A INVX1_LOC_19/A 0.09fF
C28445 INVX1_LOC_71/A NAND2X1_LOC_439/a_36_24# 0.00fF
C28446 INVX1_LOC_289/Y NAND2X1_LOC_537/Y 0.14fF
C28447 NOR2X1_LOC_246/A NOR2X1_LOC_661/A 0.00fF
C28448 NOR2X1_LOC_91/A NAND2X1_LOC_787/B 0.05fF
C28449 INVX1_LOC_33/A NOR2X1_LOC_318/A 0.03fF
C28450 NAND2X1_LOC_316/a_36_24# NAND2X1_LOC_286/B 0.00fF
C28451 NOR2X1_LOC_333/a_36_216# NOR2X1_LOC_814/A 0.01fF
C28452 INVX1_LOC_56/Y INVX1_LOC_170/Y 0.09fF
C28453 NAND2X1_LOC_577/a_36_24# INVX1_LOC_15/A 0.00fF
C28454 NOR2X1_LOC_783/A NOR2X1_LOC_779/Y 0.00fF
C28455 INVX1_LOC_30/Y INVX1_LOC_42/A 0.03fF
C28456 NOR2X1_LOC_216/Y NOR2X1_LOC_117/a_36_216# 0.00fF
C28457 INVX1_LOC_76/A INVX1_LOC_46/A 0.33fF
C28458 NOR2X1_LOC_334/a_36_216# INVX1_LOC_9/A 0.02fF
C28459 INVX1_LOC_310/Y NOR2X1_LOC_383/B 0.07fF
C28460 NOR2X1_LOC_15/Y NOR2X1_LOC_816/A 0.88fF
C28461 INVX1_LOC_25/Y INVX1_LOC_15/A 0.14fF
C28462 NOR2X1_LOC_315/Y INVX1_LOC_26/A 0.03fF
C28463 NOR2X1_LOC_683/Y INVX1_LOC_117/A 0.06fF
C28464 NOR2X1_LOC_168/A NAND2X1_LOC_72/B 0.01fF
C28465 INVX1_LOC_2/A NOR2X1_LOC_338/a_36_216# 0.00fF
C28466 NOR2X1_LOC_554/B INVX1_LOC_50/Y 0.07fF
C28467 INVX1_LOC_20/A NOR2X1_LOC_765/Y 0.02fF
C28468 INVX1_LOC_36/A NAND2X1_LOC_474/Y 0.10fF
C28469 NOR2X1_LOC_91/A INVX1_LOC_304/Y 0.09fF
C28470 INVX1_LOC_75/A INVX1_LOC_84/A 0.21fF
C28471 INVX1_LOC_39/A NOR2X1_LOC_384/Y 0.11fF
C28472 NOR2X1_LOC_827/a_36_216# INVX1_LOC_26/Y 0.00fF
C28473 NAND2X1_LOC_866/B INVX1_LOC_12/A 0.07fF
C28474 INVX1_LOC_278/A NOR2X1_LOC_373/a_36_216# 0.01fF
C28475 NOR2X1_LOC_121/A INVX1_LOC_4/Y 0.03fF
C28476 NOR2X1_LOC_458/Y NOR2X1_LOC_456/Y -0.10fF
C28477 NOR2X1_LOC_267/A NAND2X1_LOC_474/Y 0.05fF
C28478 INVX1_LOC_147/A INVX1_LOC_63/A 0.06fF
C28479 NOR2X1_LOC_643/A INVX1_LOC_31/A 0.02fF
C28480 INVX1_LOC_223/Y NOR2X1_LOC_168/Y 0.01fF
C28481 NOR2X1_LOC_75/Y INVX1_LOC_245/Y 0.02fF
C28482 NOR2X1_LOC_76/A NOR2X1_LOC_76/B 0.04fF
C28483 INVX1_LOC_41/A NOR2X1_LOC_668/a_36_216# 0.00fF
C28484 NOR2X1_LOC_791/Y INVX1_LOC_181/Y 0.02fF
C28485 INVX1_LOC_5/A NOR2X1_LOC_860/B 0.14fF
C28486 NOR2X1_LOC_454/Y INVX1_LOC_72/A 0.06fF
C28487 INVX1_LOC_33/A NOR2X1_LOC_678/A 0.03fF
C28488 INVX1_LOC_228/Y INVX1_LOC_31/A 0.05fF
C28489 NAND2X1_LOC_564/A NOR2X1_LOC_315/Y 0.01fF
C28490 INVX1_LOC_200/A INVX1_LOC_31/A 0.10fF
C28491 NOR2X1_LOC_510/Y NOR2X1_LOC_759/Y 0.00fF
C28492 NOR2X1_LOC_188/Y INVX1_LOC_4/Y 0.03fF
C28493 INVX1_LOC_21/A INVX1_LOC_41/Y 0.03fF
C28494 INVX1_LOC_313/Y INVX1_LOC_290/Y 0.50fF
C28495 NAND2X1_LOC_722/A NAND2X1_LOC_787/Y 0.01fF
C28496 INVX1_LOC_58/A NOR2X1_LOC_200/a_36_216# 0.00fF
C28497 INVX1_LOC_35/A NOR2X1_LOC_843/A 0.04fF
C28498 INVX1_LOC_77/A NOR2X1_LOC_674/Y 0.06fF
C28499 INVX1_LOC_30/Y INVX1_LOC_78/A 0.03fF
C28500 NOR2X1_LOC_598/B NOR2X1_LOC_180/Y 0.03fF
C28501 NAND2X1_LOC_638/Y NOR2X1_LOC_48/B 0.04fF
C28502 NAND2X1_LOC_740/Y NOR2X1_LOC_577/Y 0.18fF
C28503 INVX1_LOC_35/A INVX1_LOC_82/A 0.01fF
C28504 NAND2X1_LOC_579/A NOR2X1_LOC_91/Y 0.12fF
C28505 INVX1_LOC_227/A NOR2X1_LOC_334/Y 0.02fF
C28506 INVX1_LOC_2/A NAND2X1_LOC_784/A 0.08fF
C28507 INVX1_LOC_21/A NAND2X1_LOC_593/Y 0.07fF
C28508 NOR2X1_LOC_78/Y INVX1_LOC_59/Y 0.01fF
C28509 NAND2X1_LOC_30/Y NAND2X1_LOC_3/a_36_24# 0.00fF
C28510 NOR2X1_LOC_631/B INVX1_LOC_179/A 0.07fF
C28511 INVX1_LOC_171/A INVX1_LOC_4/A 0.11fF
C28512 INVX1_LOC_102/Y INVX1_LOC_102/A 0.02fF
C28513 INVX1_LOC_223/A NOR2X1_LOC_541/Y 0.16fF
C28514 NOR2X1_LOC_188/A NAND2X1_LOC_63/Y 0.07fF
C28515 NOR2X1_LOC_721/Y NAND2X1_LOC_74/B 0.01fF
C28516 NAND2X1_LOC_563/A INVX1_LOC_57/A 0.16fF
C28517 NOR2X1_LOC_536/A INVX1_LOC_66/Y 0.09fF
C28518 NOR2X1_LOC_160/B INVX1_LOC_210/Y 0.06fF
C28519 NAND2X1_LOC_849/A NAND2X1_LOC_254/Y 0.01fF
C28520 NOR2X1_LOC_548/B NAND2X1_LOC_63/Y 0.01fF
C28521 NOR2X1_LOC_357/Y NAND2X1_LOC_93/B 0.03fF
C28522 NOR2X1_LOC_536/A NOR2X1_LOC_692/Y 0.04fF
C28523 INVX1_LOC_75/A NAND2X1_LOC_220/B 0.08fF
C28524 INVX1_LOC_11/A NOR2X1_LOC_546/A 0.01fF
C28525 NOR2X1_LOC_790/B NOR2X1_LOC_778/B 0.05fF
C28526 NOR2X1_LOC_65/B INVX1_LOC_30/Y 0.03fF
C28527 NOR2X1_LOC_455/Y NOR2X1_LOC_78/B 0.00fF
C28528 INVX1_LOC_21/A NOR2X1_LOC_758/Y 0.02fF
C28529 INVX1_LOC_34/A NOR2X1_LOC_496/Y 0.02fF
C28530 INVX1_LOC_185/A NAND2X1_LOC_804/Y 0.02fF
C28531 NOR2X1_LOC_665/A NOR2X1_LOC_383/B 0.01fF
C28532 INVX1_LOC_6/A INVX1_LOC_12/A 3.62fF
C28533 NOR2X1_LOC_163/A NAND2X1_LOC_452/Y 0.01fF
C28534 NOR2X1_LOC_439/B INVX1_LOC_15/A 0.01fF
C28535 NOR2X1_LOC_441/Y INVX1_LOC_312/Y 0.24fF
C28536 INVX1_LOC_37/A INVX1_LOC_179/A 0.05fF
C28537 NAND2X1_LOC_391/Y NAND2X1_LOC_465/Y 0.19fF
C28538 NOR2X1_LOC_789/A NAND2X1_LOC_215/A 0.01fF
C28539 INVX1_LOC_5/A INVX1_LOC_96/Y 0.92fF
C28540 D_INPUT_4 D_INPUT_5 6.66fF
C28541 INVX1_LOC_15/Y INVX1_LOC_5/A 0.09fF
C28542 NOR2X1_LOC_88/Y NAND2X1_LOC_453/A 0.07fF
C28543 NOR2X1_LOC_451/A NAND2X1_LOC_639/A 0.04fF
C28544 INVX1_LOC_34/A INVX1_LOC_52/Y -0.01fF
C28545 NOR2X1_LOC_309/Y NAND2X1_LOC_474/Y 0.28fF
C28546 INVX1_LOC_75/A INVX1_LOC_15/A 0.19fF
C28547 INVX1_LOC_136/A INVX1_LOC_286/Y 0.10fF
C28548 INVX1_LOC_45/A INVX1_LOC_223/A 0.02fF
C28549 INVX1_LOC_278/A INVX1_LOC_25/Y 0.75fF
C28550 INVX1_LOC_315/Y NAND2X1_LOC_207/B 0.02fF
C28551 NOR2X1_LOC_156/A INVX1_LOC_78/A 0.01fF
C28552 INVX1_LOC_10/A INVX1_LOC_270/A 0.04fF
C28553 NAND2X1_LOC_543/Y NAND2X1_LOC_793/B 0.03fF
C28554 NOR2X1_LOC_266/B NAND2X1_LOC_572/B 0.02fF
C28555 NOR2X1_LOC_45/B INVX1_LOC_29/A 0.25fF
C28556 NOR2X1_LOC_624/A INVX1_LOC_1/A 0.00fF
C28557 NOR2X1_LOC_588/A INPUT_7 0.12fF
C28558 INPUT_0 INVX1_LOC_251/A 0.01fF
C28559 NOR2X1_LOC_336/B INVX1_LOC_18/A 0.00fF
C28560 INVX1_LOC_5/A INVX1_LOC_226/A 0.00fF
C28561 INVX1_LOC_15/Y INVX1_LOC_178/A 0.40fF
C28562 INVX1_LOC_292/A NOR2X1_LOC_303/Y 0.10fF
C28563 INVX1_LOC_140/A INVX1_LOC_273/A 0.03fF
C28564 NOR2X1_LOC_15/Y NAND2X1_LOC_562/B 0.07fF
C28565 NAND2X1_LOC_799/a_36_24# NAND2X1_LOC_714/B 0.01fF
C28566 INVX1_LOC_41/A NOR2X1_LOC_739/Y 0.01fF
C28567 NOR2X1_LOC_220/B NOR2X1_LOC_220/A 0.08fF
C28568 INVX1_LOC_84/A NAND2X1_LOC_453/A 0.03fF
C28569 NOR2X1_LOC_798/A INVX1_LOC_179/Y 0.00fF
C28570 INVX1_LOC_8/Y NOR2X1_LOC_160/B 0.03fF
C28571 INVX1_LOC_222/A INVX1_LOC_4/A 0.13fF
C28572 INVX1_LOC_64/A NOR2X1_LOC_589/A 0.10fF
C28573 NAND2X1_LOC_778/Y NOR2X1_LOC_773/Y 0.17fF
C28574 NAND2X1_LOC_9/Y INVX1_LOC_7/A 0.04fF
C28575 NAND2X1_LOC_749/a_36_24# INVX1_LOC_232/A 0.00fF
C28576 INVX1_LOC_181/Y INVX1_LOC_30/A 0.05fF
C28577 NAND2X1_LOC_624/B NOR2X1_LOC_521/Y 0.48fF
C28578 NOR2X1_LOC_56/Y NAND2X1_LOC_74/B 0.07fF
C28579 INVX1_LOC_247/A INVX1_LOC_29/A 0.00fF
C28580 NAND2X1_LOC_364/A INVX1_LOC_18/A 0.07fF
C28581 VDD INVX1_LOC_293/Y 0.75fF
C28582 INVX1_LOC_61/A NOR2X1_LOC_384/Y 0.18fF
C28583 INVX1_LOC_136/A INVX1_LOC_159/A 0.10fF
C28584 INVX1_LOC_2/A NAND2X1_LOC_326/A 0.07fF
C28585 NOR2X1_LOC_160/B INVX1_LOC_155/A 0.03fF
C28586 NOR2X1_LOC_82/A NOR2X1_LOC_516/Y 0.01fF
C28587 D_INPUT_1 INVX1_LOC_89/A 0.13fF
C28588 INVX1_LOC_299/A INVX1_LOC_149/A 0.04fF
C28589 NAND2X1_LOC_190/Y INVX1_LOC_266/Y 0.03fF
C28590 NOR2X1_LOC_541/Y INVX1_LOC_149/Y 0.11fF
C28591 INVX1_LOC_223/A INVX1_LOC_71/A 0.13fF
C28592 INVX1_LOC_136/A NOR2X1_LOC_191/B 0.04fF
C28593 INVX1_LOC_27/A INVX1_LOC_56/Y 0.01fF
C28594 NOR2X1_LOC_857/A NOR2X1_LOC_777/B 0.44fF
C28595 NAND2X1_LOC_363/B INVX1_LOC_148/Y 0.02fF
C28596 NOR2X1_LOC_617/a_36_216# INVX1_LOC_217/A 0.11fF
C28597 NAND2X1_LOC_656/A NOR2X1_LOC_360/Y 0.10fF
C28598 NOR2X1_LOC_391/A INVX1_LOC_306/Y 0.07fF
C28599 INVX1_LOC_280/Y NAND2X1_LOC_561/B 0.03fF
C28600 NOR2X1_LOC_15/Y NOR2X1_LOC_773/Y 0.19fF
C28601 NOR2X1_LOC_620/Y NOR2X1_LOC_500/B 0.20fF
C28602 VDD NAND2X1_LOC_74/B 3.21fF
C28603 INVX1_LOC_77/A INVX1_LOC_72/A 4.85fF
C28604 NAND2X1_LOC_354/Y NAND2X1_LOC_593/Y 0.01fF
C28605 NOR2X1_LOC_536/A NAND2X1_LOC_489/Y 0.02fF
C28606 NOR2X1_LOC_590/A NOR2X1_LOC_718/B 0.14fF
C28607 INPUT_4 D_INPUT_5 0.09fF
C28608 NOR2X1_LOC_434/Y INVX1_LOC_83/A 0.03fF
C28609 INVX1_LOC_249/A NOR2X1_LOC_735/a_36_216# 0.00fF
C28610 INVX1_LOC_21/A NAND2X1_LOC_692/a_36_24# 0.00fF
C28611 INVX1_LOC_304/Y INVX1_LOC_31/A 0.43fF
C28612 NOR2X1_LOC_34/B INVX1_LOC_83/A 0.04fF
C28613 INVX1_LOC_96/A INVX1_LOC_78/A 0.05fF
C28614 INVX1_LOC_77/A INVX1_LOC_198/Y 0.05fF
C28615 NOR2X1_LOC_389/A INVX1_LOC_266/Y 0.10fF
C28616 VDD NOR2X1_LOC_847/B -0.00fF
C28617 INVX1_LOC_45/A INVX1_LOC_149/Y 0.39fF
C28618 INVX1_LOC_305/A INVX1_LOC_33/A 0.50fF
C28619 NOR2X1_LOC_722/Y INVX1_LOC_63/Y 0.01fF
C28620 INVX1_LOC_14/A INVX1_LOC_16/A 0.13fF
C28621 NAND2X1_LOC_212/Y NOR2X1_LOC_467/A 0.01fF
C28622 NOR2X1_LOC_568/A INVX1_LOC_149/Y 0.03fF
C28623 NAND2X1_LOC_199/B INVX1_LOC_266/Y 0.01fF
C28624 NAND2X1_LOC_572/B INVX1_LOC_46/Y -0.01fF
C28625 NOR2X1_LOC_220/A INVX1_LOC_225/Y 0.03fF
C28626 INVX1_LOC_163/A NOR2X1_LOC_459/A 0.12fF
C28627 INVX1_LOC_254/A NOR2X1_LOC_350/A 0.00fF
C28628 NOR2X1_LOC_242/A NAND2X1_LOC_45/Y 0.10fF
C28629 NOR2X1_LOC_816/A NAND2X1_LOC_840/B 0.17fF
C28630 INVX1_LOC_278/A INVX1_LOC_75/A 0.46fF
C28631 INPUT_6 NAND2X1_LOC_51/B 0.10fF
C28632 INVX1_LOC_279/A NOR2X1_LOC_122/A 0.01fF
C28633 INVX1_LOC_20/A INVX1_LOC_4/A 0.47fF
C28634 NOR2X1_LOC_6/B NOR2X1_LOC_554/B 0.02fF
C28635 NAND2X1_LOC_453/A INVX1_LOC_15/A 0.08fF
C28636 INVX1_LOC_214/Y INVX1_LOC_31/A 0.03fF
C28637 NAND2X1_LOC_775/a_36_24# INVX1_LOC_30/A 0.00fF
C28638 INVX1_LOC_14/A NAND2X1_LOC_388/a_36_24# 0.00fF
C28639 INVX1_LOC_124/Y INVX1_LOC_98/Y 0.06fF
C28640 NAND2X1_LOC_854/B NAND2X1_LOC_538/Y 0.05fF
C28641 INVX1_LOC_124/A INVX1_LOC_72/A 0.08fF
C28642 NOR2X1_LOC_620/Y INVX1_LOC_303/A 0.02fF
C28643 NOR2X1_LOC_349/A NOR2X1_LOC_843/B 0.21fF
C28644 NOR2X1_LOC_67/A NOR2X1_LOC_382/Y 0.01fF
C28645 NAND2X1_LOC_650/B NAND2X1_LOC_444/B 0.03fF
C28646 INVX1_LOC_13/A NOR2X1_LOC_647/B 0.03fF
C28647 NOR2X1_LOC_718/Y INVX1_LOC_113/Y 0.01fF
C28648 INVX1_LOC_107/A INVX1_LOC_266/Y 0.01fF
C28649 INVX1_LOC_225/Y NOR2X1_LOC_548/Y 0.02fF
C28650 INVX1_LOC_71/A INVX1_LOC_149/Y 0.03fF
C28651 NOR2X1_LOC_471/Y GATE_479 0.01fF
C28652 NAND2X1_LOC_785/Y INVX1_LOC_41/Y 0.01fF
C28653 NOR2X1_LOC_189/A NOR2X1_LOC_690/A 0.01fF
C28654 INVX1_LOC_162/Y INVX1_LOC_71/A 0.10fF
C28655 INVX1_LOC_61/Y INVX1_LOC_232/A 0.05fF
C28656 NAND2X1_LOC_778/Y INVX1_LOC_140/A 0.10fF
C28657 NOR2X1_LOC_445/Y NOR2X1_LOC_577/Y 0.01fF
C28658 INVX1_LOC_233/A NOR2X1_LOC_167/Y 0.01fF
C28659 INVX1_LOC_49/A NOR2X1_LOC_285/B 0.01fF
C28660 NOR2X1_LOC_78/A NOR2X1_LOC_858/A 0.00fF
C28661 INVX1_LOC_222/Y NOR2X1_LOC_567/B 0.10fF
C28662 INVX1_LOC_286/A NOR2X1_LOC_717/A 0.20fF
C28663 INVX1_LOC_85/A INVX1_LOC_71/A 0.01fF
C28664 NOR2X1_LOC_590/A NOR2X1_LOC_569/Y 0.72fF
C28665 NAND2X1_LOC_11/Y INVX1_LOC_18/A 0.28fF
C28666 NAND2X1_LOC_840/Y NOR2X1_LOC_406/A 0.02fF
C28667 NOR2X1_LOC_596/A INVX1_LOC_266/Y 0.14fF
C28668 NOR2X1_LOC_536/A INVX1_LOC_32/A 0.07fF
C28669 NOR2X1_LOC_717/Y INVX1_LOC_16/A 0.01fF
C28670 NOR2X1_LOC_412/a_36_216# NOR2X1_LOC_690/A 0.00fF
C28671 INVX1_LOC_226/Y INVX1_LOC_36/A 0.04fF
C28672 NOR2X1_LOC_219/B NOR2X1_LOC_142/Y 0.03fF
C28673 NAND2X1_LOC_163/a_36_24# INVX1_LOC_49/A 0.02fF
C28674 INVX1_LOC_136/A NOR2X1_LOC_568/a_36_216# 0.06fF
C28675 INVX1_LOC_29/A NOR2X1_LOC_862/B 1.80fF
C28676 INVX1_LOC_13/A NOR2X1_LOC_606/Y 0.44fF
C28677 NAND2X1_LOC_35/Y INVX1_LOC_309/A 0.03fF
C28678 INVX1_LOC_34/A INVX1_LOC_63/Y 0.08fF
C28679 INVX1_LOC_256/A NOR2X1_LOC_246/A 0.01fF
C28680 NAND2X1_LOC_785/A INVX1_LOC_172/A 0.07fF
C28681 INVX1_LOC_14/A INVX1_LOC_28/A 0.07fF
C28682 NAND2X1_LOC_338/B NAND2X1_LOC_101/a_36_24# 0.00fF
C28683 NOR2X1_LOC_15/Y INVX1_LOC_140/A 0.11fF
C28684 INVX1_LOC_153/Y INVX1_LOC_249/Y 0.12fF
C28685 INVX1_LOC_77/A INVX1_LOC_192/Y 0.06fF
C28686 INVX1_LOC_177/A NOR2X1_LOC_550/B 0.03fF
C28687 NOR2X1_LOC_384/Y NOR2X1_LOC_85/a_36_216# 0.01fF
C28688 INVX1_LOC_58/A NAND2X1_LOC_468/B 0.03fF
C28689 NOR2X1_LOC_122/A INVX1_LOC_182/Y 0.00fF
C28690 NOR2X1_LOC_441/Y NAND2X1_LOC_656/Y 0.27fF
C28691 INVX1_LOC_31/A NAND2X1_LOC_808/A 0.07fF
C28692 INVX1_LOC_37/A NOR2X1_LOC_693/Y 0.07fF
C28693 NAND2X1_LOC_338/B INVX1_LOC_77/A 0.14fF
C28694 NAND2X1_LOC_35/Y INVX1_LOC_91/A 0.08fF
C28695 INVX1_LOC_288/Y VDD -0.00fF
C28696 INVX1_LOC_18/A NOR2X1_LOC_86/A 0.01fF
C28697 INVX1_LOC_78/A NOR2X1_LOC_684/Y 0.04fF
C28698 NOR2X1_LOC_15/Y NAND2X1_LOC_463/B 0.00fF
C28699 INVX1_LOC_36/A INVX1_LOC_10/A 1.17fF
C28700 INVX1_LOC_208/A NOR2X1_LOC_363/a_36_216# 0.01fF
C28701 NOR2X1_LOC_536/A NAND2X1_LOC_175/Y 0.04fF
C28702 NOR2X1_LOC_486/Y NOR2X1_LOC_678/A 0.03fF
C28703 NAND2X1_LOC_739/B INVX1_LOC_16/A 0.03fF
C28704 NAND2X1_LOC_323/B INVX1_LOC_77/A 0.23fF
C28705 NOR2X1_LOC_420/Y INVX1_LOC_125/Y 0.02fF
C28706 NAND2X1_LOC_96/A INVX1_LOC_26/A 0.01fF
C28707 NOR2X1_LOC_414/a_36_216# INVX1_LOC_135/A 0.00fF
C28708 INVX1_LOC_32/A NAND2X1_LOC_93/B 0.02fF
C28709 NAND2X1_LOC_703/Y NOR2X1_LOC_167/Y 0.00fF
C28710 NAND2X1_LOC_624/B INVX1_LOC_255/A 0.00fF
C28711 NAND2X1_LOC_231/Y INVX1_LOC_63/Y 0.01fF
C28712 NAND2X1_LOC_35/Y INVX1_LOC_11/Y 0.07fF
C28713 INVX1_LOC_25/A D_INPUT_3 0.02fF
C28714 NAND2X1_LOC_659/B NOR2X1_LOC_660/Y 0.12fF
C28715 INVX1_LOC_182/Y INVX1_LOC_161/Y -0.01fF
C28716 NOR2X1_LOC_778/B NOR2X1_LOC_344/A 0.11fF
C28717 NAND2X1_LOC_731/a_36_24# NAND2X1_LOC_731/Y 0.00fF
C28718 NOR2X1_LOC_498/Y NAND2X1_LOC_374/Y 0.62fF
C28719 NAND2X1_LOC_9/Y INVX1_LOC_76/A 0.17fF
C28720 INVX1_LOC_215/A NOR2X1_LOC_13/Y 0.10fF
C28721 INVX1_LOC_15/Y NAND2X1_LOC_562/B 0.08fF
C28722 NAND2X1_LOC_72/Y NAND2X1_LOC_447/Y 0.44fF
C28723 INVX1_LOC_150/Y INVX1_LOC_73/A 0.07fF
C28724 INVX1_LOC_12/Y INVX1_LOC_57/A 0.08fF
C28725 INVX1_LOC_32/A NAND2X1_LOC_425/Y 0.01fF
C28726 INVX1_LOC_233/A INVX1_LOC_76/A 0.10fF
C28727 INVX1_LOC_259/Y VDD 0.42fF
C28728 NOR2X1_LOC_804/B NOR2X1_LOC_500/Y 0.02fF
C28729 INVX1_LOC_208/A INVX1_LOC_155/A 0.00fF
C28730 INVX1_LOC_64/A INVX1_LOC_20/A 0.21fF
C28731 INVX1_LOC_177/Y NOR2X1_LOC_106/A 0.00fF
C28732 NOR2X1_LOC_649/a_36_216# NOR2X1_LOC_516/B 0.00fF
C28733 INVX1_LOC_109/Y INVX1_LOC_186/Y 0.02fF
C28734 NOR2X1_LOC_437/Y INVX1_LOC_279/A 0.68fF
C28735 VDD NOR2X1_LOC_660/Y 0.36fF
C28736 NOR2X1_LOC_208/Y INVX1_LOC_10/A 0.01fF
C28737 INVX1_LOC_229/Y NAND2X1_LOC_863/Y 0.67fF
C28738 NOR2X1_LOC_607/A NOR2X1_LOC_355/A 0.00fF
C28739 INVX1_LOC_217/A NAND2X1_LOC_866/B 0.03fF
C28740 NOR2X1_LOC_227/B NOR2X1_LOC_78/A 0.01fF
C28741 NOR2X1_LOC_833/Y NOR2X1_LOC_840/A 0.07fF
C28742 NAND2X1_LOC_358/B VDD 0.01fF
C28743 INVX1_LOC_135/A NAND2X1_LOC_79/Y 0.02fF
C28744 INVX1_LOC_32/A NOR2X1_LOC_649/B 0.07fF
C28745 NAND2X1_LOC_553/A INVX1_LOC_76/A 0.01fF
C28746 NAND2X1_LOC_811/Y NAND2X1_LOC_863/B 0.44fF
C28747 INVX1_LOC_32/A INVX1_LOC_3/A 0.16fF
C28748 NOR2X1_LOC_860/B NOR2X1_LOC_332/A 0.09fF
C28749 NAND2X1_LOC_181/Y INVX1_LOC_168/A 0.02fF
C28750 INVX1_LOC_203/Y NOR2X1_LOC_459/A 0.01fF
C28751 NAND2X1_LOC_35/Y NOR2X1_LOC_290/a_36_216# 0.01fF
C28752 D_INPUT_0 NOR2X1_LOC_419/Y 0.01fF
C28753 INVX1_LOC_89/A D_INPUT_2 0.02fF
C28754 NOR2X1_LOC_822/Y NAND2X1_LOC_852/Y 0.05fF
C28755 NAND2X1_LOC_288/B NOR2X1_LOC_743/Y 0.40fF
C28756 INVX1_LOC_26/Y NOR2X1_LOC_624/B 0.01fF
C28757 NOR2X1_LOC_194/Y INVX1_LOC_290/A 0.06fF
C28758 NOR2X1_LOC_91/A INVX1_LOC_92/A 0.03fF
C28759 NOR2X1_LOC_278/a_36_216# NOR2X1_LOC_716/B 0.01fF
C28760 INVX1_LOC_234/A NAND2X1_LOC_673/a_36_24# 0.01fF
C28761 D_INPUT_0 NOR2X1_LOC_716/B 0.14fF
C28762 INVX1_LOC_16/A NOR2X1_LOC_612/B 0.05fF
C28763 NOR2X1_LOC_142/Y NAND2X1_LOC_656/Y 0.10fF
C28764 NOR2X1_LOC_68/A NOR2X1_LOC_742/A 0.03fF
C28765 INVX1_LOC_304/Y NAND2X1_LOC_859/Y 0.01fF
C28766 INVX1_LOC_77/A INVX1_LOC_313/Y 0.05fF
C28767 INVX1_LOC_33/A NOR2X1_LOC_354/a_36_216# 0.00fF
C28768 NOR2X1_LOC_309/Y INVX1_LOC_10/A 0.03fF
C28769 NAND2X1_LOC_866/B NAND2X1_LOC_787/B 0.10fF
C28770 INVX1_LOC_75/A NOR2X1_LOC_168/Y 0.01fF
C28771 INVX1_LOC_13/Y INVX1_LOC_117/A 0.04fF
C28772 INVX1_LOC_215/Y NAND2X1_LOC_655/A 0.02fF
C28773 NAND2X1_LOC_703/Y NAND2X1_LOC_405/a_36_24# 0.00fF
C28774 NOR2X1_LOC_655/B NOR2X1_LOC_789/A 0.17fF
C28775 NOR2X1_LOC_778/B NOR2X1_LOC_540/a_36_216# 0.00fF
C28776 INVX1_LOC_23/A INVX1_LOC_92/A 0.19fF
C28777 NOR2X1_LOC_437/Y INVX1_LOC_182/Y 0.02fF
C28778 INVX1_LOC_50/A NAND2X1_LOC_750/a_36_24# 0.01fF
C28779 INVX1_LOC_1/A D_INPUT_3 0.37fF
C28780 NOR2X1_LOC_596/A INVX1_LOC_42/Y 0.04fF
C28781 NOR2X1_LOC_321/Y NOR2X1_LOC_111/A 0.02fF
C28782 NOR2X1_LOC_589/A NAND2X1_LOC_850/Y 0.03fF
C28783 NOR2X1_LOC_557/Y INVX1_LOC_87/Y 0.01fF
C28784 INVX1_LOC_1/A INVX1_LOC_14/Y 0.10fF
C28785 NOR2X1_LOC_332/A NAND2X1_LOC_141/A 0.00fF
C28786 NOR2X1_LOC_516/B INVX1_LOC_316/Y 0.11fF
C28787 INVX1_LOC_217/A INVX1_LOC_6/A 0.05fF
C28788 INVX1_LOC_138/Y NOR2X1_LOC_860/Y 0.01fF
C28789 NOR2X1_LOC_848/Y INVX1_LOC_36/Y 0.04fF
C28790 INVX1_LOC_1/A NAND2X1_LOC_618/a_36_24# 0.00fF
C28791 NAND2X1_LOC_355/Y INVX1_LOC_6/A 0.01fF
C28792 NAND2X1_LOC_646/a_36_24# INVX1_LOC_12/A 0.01fF
C28793 NOR2X1_LOC_674/Y INVX1_LOC_9/A 0.01fF
C28794 INVX1_LOC_12/A NOR2X1_LOC_80/Y 0.81fF
C28795 NAND2X1_LOC_79/Y NOR2X1_LOC_391/B 0.06fF
C28796 INVX1_LOC_304/Y NAND2X1_LOC_866/B 0.01fF
C28797 INVX1_LOC_256/A NOR2X1_LOC_357/Y 0.03fF
C28798 INVX1_LOC_81/Y NOR2X1_LOC_657/B 0.10fF
C28799 NOR2X1_LOC_45/B NAND2X1_LOC_634/Y 0.56fF
C28800 INVX1_LOC_58/A NOR2X1_LOC_66/Y 0.03fF
C28801 NOR2X1_LOC_601/a_36_216# NOR2X1_LOC_155/A 0.00fF
C28802 INVX1_LOC_162/Y INVX1_LOC_102/Y 0.13fF
C28803 INVX1_LOC_211/A VDD -0.00fF
C28804 INVX1_LOC_273/A INVX1_LOC_42/A 0.04fF
C28805 INVX1_LOC_18/A NOR2X1_LOC_113/A 0.02fF
C28806 INVX1_LOC_21/A INVX1_LOC_185/A 0.03fF
C28807 NOR2X1_LOC_276/Y VDD 0.12fF
C28808 INVX1_LOC_18/A NOR2X1_LOC_405/A 0.17fF
C28809 INVX1_LOC_143/A INVX1_LOC_87/Y 0.01fF
C28810 NAND2X1_LOC_49/a_36_24# NOR2X1_LOC_130/A 0.01fF
C28811 INVX1_LOC_227/A NOR2X1_LOC_569/Y 0.17fF
C28812 NAND2X1_LOC_326/A INVX1_LOC_118/A 0.10fF
C28813 INVX1_LOC_94/A INVX1_LOC_91/A 0.17fF
C28814 INVX1_LOC_136/A NOR2X1_LOC_56/Y 0.10fF
C28815 INVX1_LOC_75/A INVX1_LOC_76/Y 0.03fF
C28816 NOR2X1_LOC_137/A INVX1_LOC_16/A 0.07fF
C28817 INVX1_LOC_85/Y NOR2X1_LOC_731/Y 0.01fF
C28818 NOR2X1_LOC_789/A NOR2X1_LOC_99/B 0.01fF
C28819 INVX1_LOC_32/A NAND2X1_LOC_470/B 0.06fF
C28820 INVX1_LOC_12/A INVX1_LOC_270/A 0.07fF
C28821 NOR2X1_LOC_315/Y NOR2X1_LOC_368/A 0.04fF
C28822 NOR2X1_LOC_590/A NAND2X1_LOC_472/Y 0.07fF
C28823 INVX1_LOC_27/A NOR2X1_LOC_831/B 0.07fF
C28824 INVX1_LOC_229/Y NOR2X1_LOC_700/a_36_216# 0.02fF
C28825 NOR2X1_LOC_641/B INVX1_LOC_37/A 0.08fF
C28826 D_INPUT_4 NAND2X1_LOC_451/Y 0.00fF
C28827 INVX1_LOC_41/Y INVX1_LOC_304/A 0.00fF
C28828 NOR2X1_LOC_641/B NOR2X1_LOC_231/A 0.01fF
C28829 NOR2X1_LOC_577/Y INVX1_LOC_264/Y 0.01fF
C28830 NAND2X1_LOC_35/Y INVX1_LOC_203/A 0.10fF
C28831 INPUT_3 NOR2X1_LOC_536/A 0.03fF
C28832 NOR2X1_LOC_500/A NOR2X1_LOC_542/B 0.02fF
C28833 NAND2X1_LOC_783/Y NAND2X1_LOC_848/A 0.37fF
C28834 INPUT_0 NOR2X1_LOC_175/A 0.03fF
C28835 NOR2X1_LOC_617/Y INVX1_LOC_255/A 0.01fF
C28836 INVX1_LOC_136/A VDD 8.22fF
C28837 NAND2X1_LOC_361/Y NOR2X1_LOC_78/A 0.11fF
C28838 NOR2X1_LOC_751/Y INVX1_LOC_37/A 0.03fF
C28839 NAND2X1_LOC_358/Y INVX1_LOC_132/Y 0.00fF
C28840 NAND2X1_LOC_807/A INVX1_LOC_118/A 0.03fF
C28841 NOR2X1_LOC_751/Y NOR2X1_LOC_231/A 0.01fF
C28842 INVX1_LOC_136/A NAND2X1_LOC_800/A 0.03fF
C28843 NOR2X1_LOC_500/B INVX1_LOC_117/A 0.07fF
C28844 NOR2X1_LOC_136/Y INVX1_LOC_79/A 0.16fF
C28845 INVX1_LOC_135/A NOR2X1_LOC_333/A 0.01fF
C28846 NOR2X1_LOC_226/A NOR2X1_LOC_815/A 0.01fF
C28847 NOR2X1_LOC_561/Y NAND2X1_LOC_842/B 0.07fF
C28848 NOR2X1_LOC_68/A NAND2X1_LOC_721/A 0.26fF
C28849 NAND2X1_LOC_803/B NAND2X1_LOC_434/Y 0.06fF
C28850 NAND2X1_LOC_832/a_36_24# INVX1_LOC_6/A 0.01fF
C28851 NAND2X1_LOC_866/A INVX1_LOC_76/A 0.18fF
C28852 NAND2X1_LOC_474/Y INVX1_LOC_63/A 0.07fF
C28853 NOR2X1_LOC_414/a_36_216# INVX1_LOC_280/A 0.01fF
C28854 INPUT_3 NOR2X1_LOC_655/Y 0.05fF
C28855 INVX1_LOC_13/A NAND2X1_LOC_293/a_36_24# 0.00fF
C28856 D_INPUT_0 NOR2X1_LOC_130/Y 0.01fF
C28857 INVX1_LOC_124/Y NOR2X1_LOC_709/B 0.23fF
C28858 NOR2X1_LOC_274/Y INVX1_LOC_46/A 0.01fF
C28859 NOR2X1_LOC_720/B NAND2X1_LOC_642/Y 0.01fF
C28860 NAND2X1_LOC_87/a_36_24# INVX1_LOC_284/A 0.01fF
C28861 INVX1_LOC_256/Y INVX1_LOC_286/A 0.10fF
C28862 INVX1_LOC_47/Y INVX1_LOC_29/Y 0.35fF
C28863 INVX1_LOC_135/A NOR2X1_LOC_750/A 0.04fF
C28864 NAND2X1_LOC_807/Y NAND2X1_LOC_808/A 0.98fF
C28865 INVX1_LOC_295/A D_GATE_366 0.04fF
C28866 NOR2X1_LOC_392/B INVX1_LOC_95/Y 0.10fF
C28867 INVX1_LOC_5/A INVX1_LOC_99/A 0.45fF
C28868 NOR2X1_LOC_658/Y INVX1_LOC_54/A 0.07fF
C28869 NOR2X1_LOC_510/Y NAND2X1_LOC_74/B 0.07fF
C28870 INVX1_LOC_178/A INVX1_LOC_49/Y 0.03fF
C28871 INVX1_LOC_90/A INVX1_LOC_47/A 0.04fF
C28872 INVX1_LOC_72/A INVX1_LOC_9/A 0.07fF
C28873 INVX1_LOC_28/A NOR2X1_LOC_137/A 0.07fF
C28874 INVX1_LOC_120/A NOR2X1_LOC_112/Y 0.04fF
C28875 NOR2X1_LOC_716/B NOR2X1_LOC_266/B 0.03fF
C28876 INVX1_LOC_135/A NOR2X1_LOC_750/a_36_216# 0.00fF
C28877 INVX1_LOC_155/A NAND2X1_LOC_211/Y 0.02fF
C28878 NOR2X1_LOC_389/B INVX1_LOC_47/A 0.08fF
C28879 INVX1_LOC_31/A INVX1_LOC_92/A 0.47fF
C28880 INVX1_LOC_35/A D_INPUT_5 0.01fF
C28881 INVX1_LOC_229/Y INVX1_LOC_282/A 0.03fF
C28882 INVX1_LOC_26/A NAND2X1_LOC_99/A 0.03fF
C28883 NAND2X1_LOC_254/Y NOR2X1_LOC_291/Y 0.17fF
C28884 INVX1_LOC_303/A INVX1_LOC_117/A 0.07fF
C28885 NOR2X1_LOC_296/Y INVX1_LOC_3/A 0.12fF
C28886 NOR2X1_LOC_468/Y INVX1_LOC_19/A 0.03fF
C28887 NAND2X1_LOC_79/Y INVX1_LOC_280/A 0.03fF
C28888 NOR2X1_LOC_238/Y INVX1_LOC_38/A 0.03fF
C28889 NOR2X1_LOC_706/Y INVX1_LOC_174/Y 0.01fF
C28890 NOR2X1_LOC_340/A NAND2X1_LOC_473/A 0.07fF
C28891 NAND2X1_LOC_778/Y INVX1_LOC_42/A 0.01fF
C28892 INVX1_LOC_64/A INVX1_LOC_4/A 0.03fF
C28893 INVX1_LOC_256/Y INVX1_LOC_95/A 0.01fF
C28894 INPUT_3 NOR2X1_LOC_649/B 0.23fF
C28895 NAND2X1_LOC_586/a_36_24# INVX1_LOC_118/A 0.00fF
C28896 VDD NOR2X1_LOC_278/A 0.48fF
C28897 INPUT_3 INVX1_LOC_3/A 2.46fF
C28898 NOR2X1_LOC_269/a_36_216# NOR2X1_LOC_269/Y 0.01fF
C28899 NAND2X1_LOC_550/A NOR2X1_LOC_662/A 0.10fF
C28900 INVX1_LOC_13/Y INVX1_LOC_3/Y 0.03fF
C28901 NOR2X1_LOC_716/B NAND2X1_LOC_848/A 0.10fF
C28902 NOR2X1_LOC_361/B NAND2X1_LOC_74/B 0.03fF
C28903 NOR2X1_LOC_68/A INVX1_LOC_117/Y 0.05fF
C28904 INVX1_LOC_11/A INVX1_LOC_264/A 0.01fF
C28905 NAND2X1_LOC_72/B NOR2X1_LOC_405/Y 0.02fF
C28906 NAND2X1_LOC_37/a_36_24# NOR2X1_LOC_814/A 0.00fF
C28907 NOR2X1_LOC_471/a_36_216# NOR2X1_LOC_678/A 0.00fF
C28908 NAND2X1_LOC_850/Y INVX1_LOC_20/A 0.10fF
C28909 NOR2X1_LOC_15/Y INVX1_LOC_42/A 0.19fF
C28910 INVX1_LOC_98/Y NOR2X1_LOC_266/B 0.18fF
C28911 INVX1_LOC_111/A INVX1_LOC_92/A 0.02fF
C28912 NOR2X1_LOC_816/A INVX1_LOC_49/Y 0.03fF
C28913 NOR2X1_LOC_590/a_36_216# NOR2X1_LOC_742/A 0.01fF
C28914 NOR2X1_LOC_590/A NAND2X1_LOC_773/B 0.15fF
C28915 NOR2X1_LOC_389/A INVX1_LOC_19/A 0.01fF
C28916 INVX1_LOC_180/A INVX1_LOC_180/Y 0.06fF
C28917 NAND2X1_LOC_175/B INVX1_LOC_54/A 0.09fF
C28918 NOR2X1_LOC_216/Y INVX1_LOC_67/Y 0.13fF
C28919 NOR2X1_LOC_419/Y INVX1_LOC_46/Y 0.67fF
C28920 NAND2X1_LOC_778/Y INVX1_LOC_78/A 0.03fF
C28921 NOR2X1_LOC_678/A NOR2X1_LOC_748/A 0.05fF
C28922 INVX1_LOC_53/A INVX1_LOC_23/A 0.40fF
C28923 INVX1_LOC_24/A INVX1_LOC_285/A 0.42fF
C28924 NOR2X1_LOC_716/B INVX1_LOC_46/Y -0.01fF
C28925 NOR2X1_LOC_706/A INVX1_LOC_86/A 0.21fF
C28926 NOR2X1_LOC_701/Y VDD 0.18fF
C28927 NOR2X1_LOC_577/Y NOR2X1_LOC_88/Y 0.07fF
C28928 D_INPUT_1 NOR2X1_LOC_392/Y 0.14fF
C28929 INVX1_LOC_24/A NOR2X1_LOC_814/A 0.07fF
C28930 NOR2X1_LOC_408/a_36_216# D_INPUT_5 0.00fF
C28931 NOR2X1_LOC_537/Y INVX1_LOC_9/A 0.13fF
C28932 INVX1_LOC_256/A INVX1_LOC_32/A 0.07fF
C28933 NAND2X1_LOC_338/B INVX1_LOC_9/A 0.07fF
C28934 NOR2X1_LOC_774/a_36_216# NOR2X1_LOC_765/Y 0.00fF
C28935 INVX1_LOC_36/A INVX1_LOC_12/A 0.32fF
C28936 NOR2X1_LOC_15/Y INVX1_LOC_78/A 0.38fF
C28937 INVX1_LOC_58/A NOR2X1_LOC_772/B 1.51fF
C28938 NOR2X1_LOC_52/Y INVX1_LOC_29/A 0.06fF
C28939 NAND2X1_LOC_702/a_36_24# INVX1_LOC_271/A 0.00fF
C28940 INVX1_LOC_90/A INVX1_LOC_95/Y 0.02fF
C28941 NOR2X1_LOC_303/Y NOR2X1_LOC_631/A 0.08fF
C28942 INVX1_LOC_62/Y INVX1_LOC_19/A 0.08fF
C28943 NOR2X1_LOC_577/Y INVX1_LOC_84/A 0.14fF
C28944 NOR2X1_LOC_389/B INVX1_LOC_95/Y 0.02fF
C28945 NOR2X1_LOC_557/Y INVX1_LOC_285/A 0.15fF
C28946 INVX1_LOC_256/Y INVX1_LOC_54/A 0.54fF
C28947 NAND2X1_LOC_564/B NOR2X1_LOC_536/A 2.79fF
C28948 INVX1_LOC_58/A INVX1_LOC_13/Y 0.03fF
C28949 NAND2X1_LOC_796/B INVX1_LOC_50/A 0.00fF
C28950 NOR2X1_LOC_653/B INVX1_LOC_57/A 0.06fF
C28951 D_INPUT_0 NAND2X1_LOC_633/Y 0.07fF
C28952 INVX1_LOC_268/A INVX1_LOC_38/A 0.03fF
C28953 NOR2X1_LOC_667/A INVX1_LOC_185/A 0.08fF
C28954 NOR2X1_LOC_734/a_36_216# NOR2X1_LOC_9/Y 0.00fF
C28955 NAND2X1_LOC_149/Y NOR2X1_LOC_383/B 0.07fF
C28956 INVX1_LOC_11/A NOR2X1_LOC_158/Y 0.07fF
C28957 INVX1_LOC_191/Y INVX1_LOC_92/A 0.05fF
C28958 NOR2X1_LOC_557/Y NOR2X1_LOC_814/A 0.07fF
C28959 NOR2X1_LOC_71/Y INVX1_LOC_37/A 0.03fF
C28960 NOR2X1_LOC_242/A INVX1_LOC_23/A 0.03fF
C28961 NOR2X1_LOC_810/A NOR2X1_LOC_319/B 0.37fF
C28962 INVX1_LOC_144/A INVX1_LOC_91/A 0.09fF
C28963 NAND2X1_LOC_862/Y VDD 0.23fF
C28964 INVX1_LOC_90/A NOR2X1_LOC_305/Y 0.19fF
C28965 NOR2X1_LOC_65/B NOR2X1_LOC_15/Y 0.06fF
C28966 NOR2X1_LOC_91/A NOR2X1_LOC_267/a_36_216# 0.00fF
C28967 NAND2X1_LOC_842/B INVX1_LOC_76/A 0.10fF
C28968 NOR2X1_LOC_518/Y NOR2X1_LOC_48/B 0.03fF
C28969 NOR2X1_LOC_208/Y INVX1_LOC_12/A 0.07fF
C28970 NOR2X1_LOC_178/Y NAND2X1_LOC_553/A 0.08fF
C28971 NOR2X1_LOC_348/B INVX1_LOC_84/A 0.03fF
C28972 NOR2X1_LOC_441/Y INVX1_LOC_128/Y 0.00fF
C28973 NOR2X1_LOC_644/A INVX1_LOC_37/A 0.03fF
C28974 NOR2X1_LOC_712/Y INVX1_LOC_19/A 0.01fF
C28975 NAND2X1_LOC_715/a_36_24# NOR2X1_LOC_331/B 0.00fF
C28976 INVX1_LOC_41/A INVX1_LOC_125/A 0.02fF
C28977 INVX1_LOC_71/A INVX1_LOC_290/Y 0.11fF
C28978 NOR2X1_LOC_295/Y INVX1_LOC_19/A 0.02fF
C28979 INVX1_LOC_11/A NAND2X1_LOC_299/a_36_24# 0.01fF
C28980 NOR2X1_LOC_226/A NAND2X1_LOC_572/B 0.03fF
C28981 NOR2X1_LOC_828/B INVX1_LOC_37/A 0.03fF
C28982 INVX1_LOC_58/A INVX1_LOC_88/A 0.52fF
C28983 INVX1_LOC_282/A INVX1_LOC_20/A 0.10fF
C28984 INVX1_LOC_56/Y NOR2X1_LOC_216/B 0.05fF
C28985 NOR2X1_LOC_434/Y NOR2X1_LOC_798/A 0.01fF
C28986 NOR2X1_LOC_763/Y NAND2X1_LOC_637/Y 0.01fF
C28987 NOR2X1_LOC_430/A NOR2X1_LOC_48/B 0.02fF
C28988 INVX1_LOC_22/A NOR2X1_LOC_88/Y 0.03fF
C28989 INVX1_LOC_143/A NOR2X1_LOC_814/A 0.03fF
C28990 NAND2X1_LOC_662/Y NOR2X1_LOC_592/B 0.03fF
C28991 NAND2X1_LOC_550/A INVX1_LOC_57/A 0.07fF
C28992 INVX1_LOC_177/Y NOR2X1_LOC_334/Y 0.02fF
C28993 INVX1_LOC_10/A NOR2X1_LOC_435/A -0.00fF
C28994 NOR2X1_LOC_160/B INVX1_LOC_57/A 0.35fF
C28995 NOR2X1_LOC_309/Y INVX1_LOC_12/A 0.03fF
C28996 INVX1_LOC_233/Y NAND2X1_LOC_561/B 0.10fF
C28997 INVX1_LOC_313/Y INVX1_LOC_9/A 0.08fF
C28998 NOR2X1_LOC_750/A INVX1_LOC_280/A 0.03fF
C28999 NOR2X1_LOC_423/a_36_216# NOR2X1_LOC_205/Y 0.03fF
C29000 INVX1_LOC_48/A NOR2X1_LOC_35/Y 0.03fF
C29001 INVX1_LOC_68/Y NOR2X1_LOC_814/A 0.06fF
C29002 NOR2X1_LOC_188/A INVX1_LOC_14/Y 0.15fF
C29003 INVX1_LOC_27/A NOR2X1_LOC_789/B 0.01fF
C29004 NAND2X1_LOC_573/Y NOR2X1_LOC_406/A 0.11fF
C29005 NOR2X1_LOC_577/Y INVX1_LOC_15/A 0.07fF
C29006 NOR2X1_LOC_672/Y INVX1_LOC_3/Y 0.04fF
C29007 NOR2X1_LOC_500/Y INVX1_LOC_63/A 0.03fF
C29008 INVX1_LOC_22/A INVX1_LOC_84/A 0.42fF
C29009 NOR2X1_LOC_750/a_36_216# INVX1_LOC_280/A 0.01fF
C29010 INVX1_LOC_230/Y NAND2X1_LOC_205/a_36_24# 0.04fF
C29011 INVX1_LOC_226/Y INVX1_LOC_63/A 0.07fF
C29012 NOR2X1_LOC_220/A INVX1_LOC_19/A 0.04fF
C29013 INPUT_6 INVX1_LOC_174/A 0.08fF
C29014 NOR2X1_LOC_791/B INVX1_LOC_23/Y 0.08fF
C29015 INVX1_LOC_269/A INVX1_LOC_306/Y 0.10fF
C29016 NAND2X1_LOC_740/Y NOR2X1_LOC_536/Y 0.03fF
C29017 NAND2X1_LOC_724/A NOR2X1_LOC_406/A 0.07fF
C29018 INVX1_LOC_31/A INVX1_LOC_53/A 0.12fF
C29019 NOR2X1_LOC_458/B INVX1_LOC_29/A 0.01fF
C29020 NOR2X1_LOC_152/Y INVX1_LOC_273/A 0.38fF
C29021 NAND2X1_LOC_656/A INVX1_LOC_26/A 0.02fF
C29022 INVX1_LOC_62/Y INVX1_LOC_26/Y 0.08fF
C29023 INVX1_LOC_64/A INVX1_LOC_43/Y 0.28fF
C29024 NAND2X1_LOC_357/A NOR2X1_LOC_652/Y 0.03fF
C29025 INVX1_LOC_215/A NAND2X1_LOC_249/a_36_24# 0.00fF
C29026 NAND2X1_LOC_807/Y INVX1_LOC_92/A 0.07fF
C29027 NOR2X1_LOC_188/A INVX1_LOC_230/A 0.03fF
C29028 NOR2X1_LOC_130/A INVX1_LOC_285/A 0.07fF
C29029 INVX1_LOC_69/Y INVX1_LOC_66/Y 0.10fF
C29030 INVX1_LOC_10/A INVX1_LOC_63/A 0.02fF
C29031 NOR2X1_LOC_120/a_36_216# INVX1_LOC_46/Y 0.00fF
C29032 INVX1_LOC_48/Y INVX1_LOC_14/A 0.13fF
C29033 NOR2X1_LOC_772/A NOR2X1_LOC_831/B 0.02fF
C29034 INPUT_1 NAND2X1_LOC_572/B 0.46fF
C29035 NOR2X1_LOC_147/B INVX1_LOC_271/Y 0.03fF
C29036 NAND2X1_LOC_840/B INVX1_LOC_42/A 0.34fF
C29037 NOR2X1_LOC_815/A INVX1_LOC_118/A 0.03fF
C29038 INVX1_LOC_104/A NOR2X1_LOC_334/Y 0.07fF
C29039 NOR2X1_LOC_719/A INVX1_LOC_284/A 0.00fF
C29040 NOR2X1_LOC_315/Y NAND2X1_LOC_471/Y 0.00fF
C29041 NOR2X1_LOC_92/Y NOR2X1_LOC_250/A 0.03fF
C29042 NOR2X1_LOC_540/B INVX1_LOC_37/A 0.02fF
C29043 INVX1_LOC_27/A NAND2X1_LOC_352/B 0.02fF
C29044 INVX1_LOC_120/A NOR2X1_LOC_721/B 0.00fF
C29045 INVX1_LOC_79/A NOR2X1_LOC_155/A 0.01fF
C29046 NAND2X1_LOC_35/Y NOR2X1_LOC_372/Y 0.03fF
C29047 INVX1_LOC_224/Y INVX1_LOC_77/A 0.01fF
C29048 NOR2X1_LOC_198/a_36_216# NOR2X1_LOC_197/B 0.00fF
C29049 INVX1_LOC_35/A NOR2X1_LOC_360/Y 0.01fF
C29050 NOR2X1_LOC_588/A INVX1_LOC_38/A 0.03fF
C29051 INVX1_LOC_58/A INVX1_LOC_303/A 0.07fF
C29052 NAND2X1_LOC_765/a_36_24# INVX1_LOC_78/A 0.00fF
C29053 INVX1_LOC_96/Y INVX1_LOC_78/A 0.07fF
C29054 INVX1_LOC_6/A INVX1_LOC_92/A 2.06fF
C29055 NOR2X1_LOC_325/A INVX1_LOC_15/A 0.06fF
C29056 D_INPUT_2 NOR2X1_LOC_392/Y 0.01fF
C29057 INVX1_LOC_58/A NOR2X1_LOC_672/Y 0.01fF
C29058 INVX1_LOC_22/A INVX1_LOC_15/A 0.14fF
C29059 NOR2X1_LOC_728/B NOR2X1_LOC_155/A -0.00fF
C29060 INVX1_LOC_152/Y NOR2X1_LOC_860/B 0.02fF
C29061 INVX1_LOC_73/Y NOR2X1_LOC_218/A 0.24fF
C29062 NOR2X1_LOC_510/Y INVX1_LOC_136/A 0.10fF
C29063 INVX1_LOC_135/A INVX1_LOC_102/A 0.10fF
C29064 NOR2X1_LOC_246/A NOR2X1_LOC_89/A 0.07fF
C29065 NOR2X1_LOC_588/A NOR2X1_LOC_51/A 0.03fF
C29066 INVX1_LOC_187/Y INVX1_LOC_38/A 0.01fF
C29067 INVX1_LOC_45/A NOR2X1_LOC_454/Y 0.07fF
C29068 NAND2X1_LOC_579/A INVX1_LOC_141/Y 0.03fF
C29069 NAND2X1_LOC_840/B INVX1_LOC_78/A 0.00fF
C29070 NOR2X1_LOC_557/Y NOR2X1_LOC_292/a_36_216# 0.00fF
C29071 NAND2X1_LOC_551/A NOR2X1_LOC_89/A 0.42fF
C29072 NOR2X1_LOC_826/a_36_216# INVX1_LOC_217/Y 0.00fF
C29073 NOR2X1_LOC_689/A NAND2X1_LOC_717/Y 0.05fF
C29074 INVX1_LOC_140/A INVX1_LOC_49/Y 0.03fF
C29075 NOR2X1_LOC_155/A INVX1_LOC_91/A 0.10fF
C29076 INVX1_LOC_55/Y NOR2X1_LOC_89/A 0.04fF
C29077 NAND2X1_LOC_160/a_36_24# INVX1_LOC_78/A 0.00fF
C29078 NOR2X1_LOC_167/Y INVX1_LOC_119/Y 0.26fF
C29079 NAND2X1_LOC_633/Y NAND2X1_LOC_848/A 0.10fF
C29080 INVX1_LOC_239/A INVX1_LOC_195/Y 0.03fF
C29081 INVX1_LOC_80/Y INVX1_LOC_23/A 0.00fF
C29082 NOR2X1_LOC_305/Y INVX1_LOC_38/A 0.07fF
C29083 NOR2X1_LOC_415/A INVX1_LOC_32/A 0.04fF
C29084 NOR2X1_LOC_91/A NOR2X1_LOC_78/B 0.02fF
C29085 NOR2X1_LOC_389/A INVX1_LOC_161/Y 0.10fF
C29086 INVX1_LOC_2/A NOR2X1_LOC_654/A 0.08fF
C29087 INVX1_LOC_235/Y NOR2X1_LOC_480/A 0.03fF
C29088 NOR2X1_LOC_647/B INPUT_3 0.00fF
C29089 INVX1_LOC_230/Y INVX1_LOC_293/A 0.02fF
C29090 NOR2X1_LOC_274/Y NOR2X1_LOC_798/A 0.02fF
C29091 NOR2X1_LOC_643/A INVX1_LOC_36/A 0.03fF
C29092 INVX1_LOC_250/A NAND2X1_LOC_724/A 0.03fF
C29093 INVX1_LOC_136/A NOR2X1_LOC_361/B 0.13fF
C29094 INVX1_LOC_35/A NOR2X1_LOC_792/B 0.01fF
C29095 NAND2X1_LOC_53/Y NAND2X1_LOC_39/a_36_24# 0.00fF
C29096 NAND2X1_LOC_725/Y NAND2X1_LOC_733/B 0.08fF
C29097 NOR2X1_LOC_634/B INVX1_LOC_23/A 0.12fF
C29098 INVX1_LOC_34/A INVX1_LOC_5/A 4.28fF
C29099 NAND2X1_LOC_729/Y NAND2X1_LOC_303/Y 0.05fF
C29100 NOR2X1_LOC_454/Y INVX1_LOC_71/A 0.07fF
C29101 INVX1_LOC_53/Y NAND2X1_LOC_288/B 0.00fF
C29102 INVX1_LOC_58/A NOR2X1_LOC_203/Y 0.01fF
C29103 NOR2X1_LOC_529/Y NOR2X1_LOC_392/Y 0.01fF
C29104 NOR2X1_LOC_78/B INVX1_LOC_23/A 1.00fF
C29105 INVX1_LOC_88/A NOR2X1_LOC_338/Y 0.00fF
C29106 NAND2X1_LOC_347/B INVX1_LOC_314/Y 0.06fF
C29107 INVX1_LOC_16/A NOR2X1_LOC_383/B 0.06fF
C29108 INVX1_LOC_176/A NOR2X1_LOC_461/A 0.14fF
C29109 NOR2X1_LOC_655/B NOR2X1_LOC_717/A 0.08fF
C29110 NOR2X1_LOC_82/A NOR2X1_LOC_68/A 0.05fF
C29111 NAND2X1_LOC_695/a_36_24# INVX1_LOC_19/A 0.00fF
C29112 INVX1_LOC_37/A NAND2X1_LOC_243/Y 0.01fF
C29113 NOR2X1_LOC_516/B INVX1_LOC_57/A 0.13fF
C29114 NOR2X1_LOC_15/Y NOR2X1_LOC_152/Y 0.32fF
C29115 INVX1_LOC_35/A NAND2X1_LOC_451/Y 0.07fF
C29116 NOR2X1_LOC_205/Y NOR2X1_LOC_759/Y 0.18fF
C29117 NOR2X1_LOC_91/A NAND2X1_LOC_392/Y 0.00fF
C29118 INVX1_LOC_34/A INVX1_LOC_178/A 0.14fF
C29119 INVX1_LOC_50/A NAND2X1_LOC_112/Y 0.03fF
C29120 D_INPUT_1 INVX1_LOC_25/Y 0.04fF
C29121 INVX1_LOC_36/A NAND2X1_LOC_733/Y 0.10fF
C29122 NOR2X1_LOC_816/A NOR2X1_LOC_518/a_36_216# 0.00fF
C29123 NOR2X1_LOC_15/Y INVX1_LOC_113/Y 0.03fF
C29124 NOR2X1_LOC_203/a_36_216# INVX1_LOC_177/A 0.00fF
C29125 NAND2X1_LOC_687/a_36_24# INVX1_LOC_291/A 0.01fF
C29126 INVX1_LOC_90/A INVX1_LOC_271/Y 0.07fF
C29127 NOR2X1_LOC_298/Y NAND2X1_LOC_828/a_36_24# 0.09fF
C29128 INVX1_LOC_47/A NAND2X1_LOC_223/A 0.01fF
C29129 NAND2X1_LOC_803/B INVX1_LOC_24/A 0.05fF
C29130 NAND2X1_LOC_35/Y NAND2X1_LOC_374/Y 0.02fF
C29131 NOR2X1_LOC_261/Y INVX1_LOC_22/A 0.07fF
C29132 INVX1_LOC_37/A NAND2X1_LOC_50/a_36_24# 0.00fF
C29133 NOR2X1_LOC_99/Y INVX1_LOC_117/A 0.09fF
C29134 INVX1_LOC_5/A NAND2X1_LOC_231/Y 0.19fF
C29135 NOR2X1_LOC_15/Y NAND2X1_LOC_676/a_36_24# 0.01fF
C29136 NAND2X1_LOC_579/A NAND2X1_LOC_483/Y 0.16fF
C29137 NOR2X1_LOC_103/Y INVX1_LOC_77/A 0.07fF
C29138 NAND2X1_LOC_350/A NOR2X1_LOC_13/Y 0.10fF
C29139 INVX1_LOC_201/Y NOR2X1_LOC_140/A 0.16fF
C29140 INVX1_LOC_41/A NAND2X1_LOC_346/a_36_24# 0.00fF
C29141 INVX1_LOC_119/Y INVX1_LOC_76/A 0.02fF
C29142 NOR2X1_LOC_280/Y INVX1_LOC_285/A 0.02fF
C29143 INPUT_4 NOR2X1_LOC_36/B 0.03fF
C29144 INVX1_LOC_77/A NOR2X1_LOC_541/Y 0.01fF
C29145 NOR2X1_LOC_590/A INVX1_LOC_24/A 0.63fF
C29146 NOR2X1_LOC_215/A INVX1_LOC_96/Y 0.02fF
C29147 INVX1_LOC_36/A INVX1_LOC_217/A 0.07fF
C29148 INVX1_LOC_5/A NAND2X1_LOC_195/a_36_24# 0.00fF
C29149 INVX1_LOC_36/A NAND2X1_LOC_355/Y 0.01fF
C29150 INVX1_LOC_69/Y INVX1_LOC_32/A 0.07fF
C29151 INVX1_LOC_83/A INVX1_LOC_23/A 3.18fF
C29152 NAND2X1_LOC_537/Y INVX1_LOC_240/A 0.04fF
C29153 NOR2X1_LOC_223/B INVX1_LOC_22/A 0.01fF
C29154 NAND2X1_LOC_725/A NAND2X1_LOC_712/A 0.09fF
C29155 NAND2X1_LOC_11/Y D_INPUT_6 0.35fF
C29156 NOR2X1_LOC_346/Y NAND2X1_LOC_207/B 0.02fF
C29157 INVX1_LOC_25/Y NOR2X1_LOC_652/Y 0.01fF
C29158 NOR2X1_LOC_445/a_36_216# INVX1_LOC_33/A 0.00fF
C29159 NOR2X1_LOC_740/Y NOR2X1_LOC_731/A 0.02fF
C29160 INVX1_LOC_34/A NOR2X1_LOC_816/A 0.03fF
C29161 INVX1_LOC_146/A NOR2X1_LOC_447/A 0.01fF
C29162 INVX1_LOC_286/Y NAND2X1_LOC_567/Y 0.01fF
C29163 INVX1_LOC_200/A NOR2X1_LOC_309/Y 0.02fF
C29164 INVX1_LOC_280/A INVX1_LOC_123/Y 0.02fF
C29165 INVX1_LOC_28/A NOR2X1_LOC_383/B 0.10fF
C29166 INVX1_LOC_58/A NAND2X1_LOC_308/B 0.08fF
C29167 INVX1_LOC_316/A NOR2X1_LOC_847/B 0.01fF
C29168 INVX1_LOC_45/A INVX1_LOC_77/A 1.26fF
C29169 INVX1_LOC_313/A INVX1_LOC_53/A 0.94fF
C29170 NOR2X1_LOC_250/A NAND2X1_LOC_477/A 0.03fF
C29171 INVX1_LOC_77/A NOR2X1_LOC_568/A 0.66fF
C29172 INVX1_LOC_1/Y NAND2X1_LOC_474/Y 0.07fF
C29173 INVX1_LOC_89/A NOR2X1_LOC_678/A 0.03fF
C29174 INVX1_LOC_206/Y NOR2X1_LOC_334/Y 0.16fF
C29175 NAND2X1_LOC_181/Y NOR2X1_LOC_271/B 0.00fF
C29176 NAND2X1_LOC_808/A NOR2X1_LOC_109/Y 0.09fF
C29177 NOR2X1_LOC_533/A NAND2X1_LOC_537/Y 0.01fF
C29178 INVX1_LOC_76/A INVX1_LOC_284/A 0.17fF
C29179 NOR2X1_LOC_561/Y NOR2X1_LOC_674/Y 0.16fF
C29180 NOR2X1_LOC_357/Y NOR2X1_LOC_89/A 0.25fF
C29181 NOR2X1_LOC_368/A NAND2X1_LOC_99/A 0.02fF
C29182 NOR2X1_LOC_211/Y INVX1_LOC_171/A 0.01fF
C29183 INVX1_LOC_54/A NOR2X1_LOC_697/Y 0.04fF
C29184 NAND2X1_LOC_375/a_36_24# INVX1_LOC_22/A 0.00fF
C29185 NOR2X1_LOC_88/A NOR2X1_LOC_88/Y 0.09fF
C29186 NOR2X1_LOC_658/Y NOR2X1_LOC_142/Y 0.13fF
C29187 NAND2X1_LOC_807/Y INVX1_LOC_53/A 0.09fF
C29188 NOR2X1_LOC_15/Y NAND2X1_LOC_859/B 0.03fF
C29189 INVX1_LOC_31/A INVX1_LOC_80/Y 0.02fF
C29190 NAND2X1_LOC_231/Y NAND2X1_LOC_337/B 0.10fF
C29191 INVX1_LOC_136/A NOR2X1_LOC_132/Y 0.02fF
C29192 INVX1_LOC_223/A NOR2X1_LOC_388/Y 0.01fF
C29193 INVX1_LOC_193/A NOR2X1_LOC_257/Y 0.02fF
C29194 NOR2X1_LOC_216/B NOR2X1_LOC_831/B 0.10fF
C29195 INVX1_LOC_2/A NAND2X1_LOC_783/Y 0.03fF
C29196 NOR2X1_LOC_724/Y INVX1_LOC_213/A 0.07fF
C29197 INVX1_LOC_27/A NOR2X1_LOC_128/B 0.08fF
C29198 D_INPUT_1 INVX1_LOC_75/A 0.26fF
C29199 NOR2X1_LOC_690/A NOR2X1_LOC_384/Y 0.05fF
C29200 INVX1_LOC_20/A NOR2X1_LOC_496/a_36_216# 0.00fF
C29201 NOR2X1_LOC_600/Y NOR2X1_LOC_334/Y 0.07fF
C29202 NAND2X1_LOC_563/Y NOR2X1_LOC_382/Y 0.02fF
C29203 NAND2X1_LOC_778/Y NAND2X1_LOC_861/Y 0.10fF
C29204 INVX1_LOC_77/A INVX1_LOC_71/A 0.19fF
C29205 INVX1_LOC_276/A INVX1_LOC_236/Y 0.00fF
C29206 NAND2X1_LOC_739/B INVX1_LOC_231/Y 0.09fF
C29207 INVX1_LOC_35/A NOR2X1_LOC_567/B 0.07fF
C29208 NOR2X1_LOC_590/A INVX1_LOC_143/A 0.08fF
C29209 INVX1_LOC_45/A INVX1_LOC_124/A 0.10fF
C29210 NOR2X1_LOC_833/B NOR2X1_LOC_698/Y 0.01fF
C29211 NOR2X1_LOC_667/Y INVX1_LOC_248/A 0.02fF
C29212 NOR2X1_LOC_78/B INVX1_LOC_31/A 5.21fF
C29213 NOR2X1_LOC_359/Y INVX1_LOC_155/Y 0.06fF
C29214 NAND2X1_LOC_541/Y INVX1_LOC_61/Y 0.01fF
C29215 NOR2X1_LOC_419/Y INVX1_LOC_49/A 0.00fF
C29216 INVX1_LOC_13/A INVX1_LOC_11/A 0.34fF
C29217 INVX1_LOC_24/A NAND2X1_LOC_354/B 0.03fF
C29218 INVX1_LOC_307/A INVX1_LOC_63/A 0.07fF
C29219 INVX1_LOC_64/A INVX1_LOC_282/A 0.07fF
C29220 INVX1_LOC_136/A INVX1_LOC_177/A 0.03fF
C29221 NOR2X1_LOC_197/B NOR2X1_LOC_814/A 0.14fF
C29222 VDD NAND2X1_LOC_647/B 0.34fF
C29223 INVX1_LOC_59/A INVX1_LOC_90/A 0.01fF
C29224 INVX1_LOC_132/A NAND2X1_LOC_361/Y 1.78fF
C29225 NOR2X1_LOC_15/Y NAND2X1_LOC_861/Y 0.19fF
C29226 NOR2X1_LOC_681/Y INVX1_LOC_21/Y 0.23fF
C29227 INVX1_LOC_6/A INVX1_LOC_53/A 2.62fF
C29228 INVX1_LOC_278/A INVX1_LOC_100/A 0.08fF
C29229 INVX1_LOC_36/A INVX1_LOC_214/Y 0.03fF
C29230 NOR2X1_LOC_445/B INVX1_LOC_63/A 0.07fF
C29231 NOR2X1_LOC_100/A NOR2X1_LOC_68/A 0.03fF
C29232 INVX1_LOC_37/A INVX1_LOC_21/Y 0.03fF
C29233 NOR2X1_LOC_331/B INVX1_LOC_290/Y 0.03fF
C29234 INVX1_LOC_50/A NOR2X1_LOC_78/A 0.06fF
C29235 INVX1_LOC_75/A NOR2X1_LOC_108/a_36_216# 0.00fF
C29236 NAND2X1_LOC_773/Y INVX1_LOC_90/A 0.01fF
C29237 NAND2X1_LOC_552/A INPUT_0 0.02fF
C29238 INVX1_LOC_75/A NOR2X1_LOC_652/Y 0.07fF
C29239 NAND2X1_LOC_803/B NAND2X1_LOC_783/A 0.01fF
C29240 INVX1_LOC_5/A INPUT_0 0.18fF
C29241 NOR2X1_LOC_91/A NOR2X1_LOC_164/Y 0.06fF
C29242 NOR2X1_LOC_419/Y INVX1_LOC_60/A 0.04fF
C29243 NAND2X1_LOC_773/Y NOR2X1_LOC_389/B 0.10fF
C29244 INVX1_LOC_124/A INVX1_LOC_71/A 0.69fF
C29245 INVX1_LOC_12/A NOR2X1_LOC_435/A 0.03fF
C29246 NAND2X1_LOC_725/A INVX1_LOC_309/A 0.05fF
C29247 NOR2X1_LOC_599/A NAND2X1_LOC_863/B 0.01fF
C29248 INVX1_LOC_11/A NOR2X1_LOC_246/A 0.09fF
C29249 NAND2X1_LOC_803/B NOR2X1_LOC_130/A 0.02fF
C29250 NOR2X1_LOC_689/Y INVX1_LOC_11/Y 0.03fF
C29251 INVX1_LOC_45/A NOR2X1_LOC_687/Y 0.03fF
C29252 NOR2X1_LOC_824/A NAND2X1_LOC_849/A 0.02fF
C29253 NOR2X1_LOC_598/B INVX1_LOC_91/A 0.07fF
C29254 NAND2X1_LOC_149/Y NOR2X1_LOC_163/Y 0.19fF
C29255 VDD NOR2X1_LOC_395/Y 0.12fF
C29256 NOR2X1_LOC_379/Y INVX1_LOC_76/Y 0.36fF
C29257 INVX1_LOC_269/A NOR2X1_LOC_356/A 0.62fF
C29258 INPUT_3 NOR2X1_LOC_415/A 0.00fF
C29259 INVX1_LOC_17/A NOR2X1_LOC_473/B 0.03fF
C29260 NOR2X1_LOC_590/A NAND2X1_LOC_783/A 0.03fF
C29261 NAND2X1_LOC_363/B NOR2X1_LOC_836/B 0.01fF
C29262 INVX1_LOC_178/A INPUT_0 0.10fF
C29263 NOR2X1_LOC_433/A INVX1_LOC_236/A 0.39fF
C29264 INVX1_LOC_84/A INVX1_LOC_186/Y 0.07fF
C29265 NOR2X1_LOC_383/B NOR2X1_LOC_35/Y 0.01fF
C29266 NOR2X1_LOC_791/B INVX1_LOC_232/A 0.07fF
C29267 NAND2X1_LOC_63/Y NAND2X1_LOC_572/B 0.03fF
C29268 INVX1_LOC_34/A NAND2X1_LOC_562/B 0.07fF
C29269 INVX1_LOC_11/A INVX1_LOC_55/Y 0.04fF
C29270 NOR2X1_LOC_91/A INVX1_LOC_46/A 9.08fF
C29271 NAND2X1_LOC_149/Y NOR2X1_LOC_74/Y 0.03fF
C29272 NOR2X1_LOC_590/A NOR2X1_LOC_130/A 0.15fF
C29273 INVX1_LOC_83/A INVX1_LOC_31/A 0.10fF
C29274 INVX1_LOC_55/A INVX1_LOC_89/A 0.01fF
C29275 NOR2X1_LOC_703/B NOR2X1_LOC_570/A 0.05fF
C29276 NOR2X1_LOC_168/Y INVX1_LOC_22/A 0.03fF
C29277 INVX1_LOC_2/A NOR2X1_LOC_716/B 0.17fF
C29278 NOR2X1_LOC_488/Y INVX1_LOC_24/A 0.03fF
C29279 INVX1_LOC_41/A NOR2X1_LOC_709/A 0.15fF
C29280 INVX1_LOC_63/Y INVX1_LOC_266/Y 0.10fF
C29281 NAND2X1_LOC_340/a_36_24# INVX1_LOC_90/A 0.00fF
C29282 NOR2X1_LOC_99/Y INVX1_LOC_3/Y 0.07fF
C29283 INVX1_LOC_38/A INVX1_LOC_271/Y 0.08fF
C29284 NOR2X1_LOC_111/A NAND2X1_LOC_211/a_36_24# 0.01fF
C29285 NOR2X1_LOC_561/Y INVX1_LOC_72/A 0.36fF
C29286 INVX1_LOC_84/A INVX1_LOC_261/A 0.05fF
C29287 INVX1_LOC_109/A NOR2X1_LOC_127/Y 0.02fF
C29288 INVX1_LOC_136/A NAND2X1_LOC_573/A 0.10fF
C29289 INVX1_LOC_33/A INVX1_LOC_196/A 0.03fF
C29290 INVX1_LOC_316/A NOR2X1_LOC_660/Y 0.10fF
C29291 NOR2X1_LOC_542/B NOR2X1_LOC_634/Y 0.01fF
C29292 NOR2X1_LOC_403/B INVX1_LOC_25/Y 0.04fF
C29293 NOR2X1_LOC_222/Y NOR2X1_LOC_214/a_36_216# 0.00fF
C29294 NAND2X1_LOC_840/B NOR2X1_LOC_152/Y 0.03fF
C29295 NOR2X1_LOC_360/Y NOR2X1_LOC_188/Y 0.27fF
C29296 NOR2X1_LOC_226/A NOR2X1_LOC_716/B 0.41fF
C29297 INVX1_LOC_304/Y NOR2X1_LOC_309/Y 0.07fF
C29298 INVX1_LOC_17/A NOR2X1_LOC_322/Y 0.77fF
C29299 INVX1_LOC_269/A NOR2X1_LOC_74/A 0.18fF
C29300 NAND2X1_LOC_725/A INVX1_LOC_11/Y 0.12fF
C29301 NOR2X1_LOC_607/a_36_216# INVX1_LOC_16/A 0.01fF
C29302 VDD NOR2X1_LOC_414/Y 0.13fF
C29303 NAND2X1_LOC_53/Y NOR2X1_LOC_742/A 0.12fF
C29304 INVX1_LOC_23/A INVX1_LOC_46/A 0.18fF
C29305 NOR2X1_LOC_91/A NOR2X1_LOC_766/Y 0.03fF
C29306 NAND2X1_LOC_337/B INVX1_LOC_131/A 0.21fF
C29307 NOR2X1_LOC_262/Y INVX1_LOC_22/A 0.01fF
C29308 INVX1_LOC_12/A INVX1_LOC_63/A 0.10fF
C29309 NOR2X1_LOC_48/B NOR2X1_LOC_697/Y 0.03fF
C29310 NOR2X1_LOC_89/A NAND2X1_LOC_489/Y 0.01fF
C29311 INVX1_LOC_159/A NAND2X1_LOC_662/a_36_24# 0.00fF
C29312 NAND2X1_LOC_36/A NOR2X1_LOC_163/A 0.07fF
C29313 INVX1_LOC_34/A NOR2X1_LOC_773/Y 0.32fF
C29314 INVX1_LOC_269/A NOR2X1_LOC_9/Y 0.10fF
C29315 NOR2X1_LOC_592/A INVX1_LOC_144/A -0.00fF
C29316 NOR2X1_LOC_267/a_36_216# INVX1_LOC_6/A 0.00fF
C29317 NAND2X1_LOC_456/Y INVX1_LOC_42/A 0.01fF
C29318 NOR2X1_LOC_638/a_36_216# INVX1_LOC_290/A 0.00fF
C29319 NAND2X1_LOC_624/B INVX1_LOC_20/A 0.00fF
C29320 INVX1_LOC_83/A NAND2X1_LOC_106/a_36_24# 0.00fF
C29321 INVX1_LOC_291/A INVX1_LOC_273/A 0.13fF
C29322 NAND2X1_LOC_21/Y INVX1_LOC_22/A 0.02fF
C29323 INVX1_LOC_268/A INVX1_LOC_33/A 0.05fF
C29324 NOR2X1_LOC_590/A NOR2X1_LOC_216/Y 0.31fF
C29325 NAND2X1_LOC_198/B NOR2X1_LOC_71/Y 0.07fF
C29326 NOR2X1_LOC_309/Y NOR2X1_LOC_566/Y 0.36fF
C29327 NAND2X1_LOC_81/B NAND2X1_LOC_74/B 0.03fF
C29328 NOR2X1_LOC_284/B NOR2X1_LOC_802/A 0.07fF
C29329 INVX1_LOC_93/Y NAND2X1_LOC_474/Y 0.08fF
C29330 NOR2X1_LOC_816/A INPUT_0 0.02fF
C29331 INVX1_LOC_57/Y INVX1_LOC_28/A 0.01fF
C29332 VDD NOR2X1_LOC_665/Y 0.07fF
C29333 INVX1_LOC_81/A NOR2X1_LOC_366/Y 0.66fF
C29334 NAND2X1_LOC_358/Y NAND2X1_LOC_364/Y 0.01fF
C29335 NOR2X1_LOC_124/B INVX1_LOC_232/A 0.01fF
C29336 NOR2X1_LOC_321/Y NOR2X1_LOC_405/A 0.01fF
C29337 INVX1_LOC_224/Y INVX1_LOC_9/A 0.05fF
C29338 INVX1_LOC_49/Y INVX1_LOC_42/A 0.07fF
C29339 INVX1_LOC_17/A NOR2X1_LOC_355/B 1.52fF
C29340 NOR2X1_LOC_654/A INVX1_LOC_118/A 0.02fF
C29341 NAND2X1_LOC_476/Y INVX1_LOC_15/A 0.01fF
C29342 INVX1_LOC_311/Y INVX1_LOC_18/A 0.01fF
C29343 INVX1_LOC_49/A NOR2X1_LOC_326/Y 0.01fF
C29344 NAND2X1_LOC_364/A INVX1_LOC_148/A 0.02fF
C29345 NOR2X1_LOC_717/B INVX1_LOC_49/A 0.03fF
C29346 NOR2X1_LOC_335/A INVX1_LOC_150/A 0.00fF
C29347 NAND2X1_LOC_231/Y NOR2X1_LOC_773/Y 0.10fF
C29348 NOR2X1_LOC_246/A NOR2X1_LOC_433/A 0.07fF
C29349 INVX1_LOC_186/Y INVX1_LOC_15/A 0.03fF
C29350 INVX1_LOC_279/A NOR2X1_LOC_147/B 0.01fF
C29351 NOR2X1_LOC_433/A NOR2X1_LOC_503/a_36_216# 0.00fF
C29352 INVX1_LOC_28/A NOR2X1_LOC_512/Y 0.00fF
C29353 INVX1_LOC_104/A NOR2X1_LOC_569/Y 0.80fF
C29354 NAND2X1_LOC_799/A INVX1_LOC_264/Y 0.02fF
C29355 NAND2X1_LOC_175/Y INVX1_LOC_297/A 0.09fF
C29356 INVX1_LOC_20/A NOR2X1_LOC_440/B 0.01fF
C29357 NOR2X1_LOC_349/A NOR2X1_LOC_345/A 0.30fF
C29358 INVX1_LOC_262/Y NOR2X1_LOC_467/A 0.02fF
C29359 INVX1_LOC_12/Y INVX1_LOC_306/Y 0.21fF
C29360 INVX1_LOC_270/A INVX1_LOC_92/A 0.08fF
C29361 INVX1_LOC_293/Y INVX1_LOC_4/Y 0.10fF
C29362 NOR2X1_LOC_716/B INPUT_1 0.16fF
C29363 INVX1_LOC_280/Y NOR2X1_LOC_701/Y 0.01fF
C29364 INVX1_LOC_21/A NAND2X1_LOC_639/A 0.14fF
C29365 INVX1_LOC_55/Y NOR2X1_LOC_593/Y 0.03fF
C29366 NOR2X1_LOC_89/A INVX1_LOC_32/A 0.07fF
C29367 INVX1_LOC_62/A NOR2X1_LOC_844/A 0.19fF
C29368 NAND2X1_LOC_722/A NOR2X1_LOC_298/Y 0.10fF
C29369 INVX1_LOC_53/A INVX1_LOC_131/Y 0.19fF
C29370 INVX1_LOC_75/A D_INPUT_2 0.12fF
C29371 NOR2X1_LOC_246/A NOR2X1_LOC_52/B 0.03fF
C29372 INVX1_LOC_7/A NOR2X1_LOC_537/Y 0.21fF
C29373 NAND2X1_LOC_74/B INVX1_LOC_4/Y 0.72fF
C29374 INVX1_LOC_58/A INVX1_LOC_107/Y 0.02fF
C29375 NOR2X1_LOC_646/A INVX1_LOC_232/A -0.08fF
C29376 INVX1_LOC_78/A INVX1_LOC_49/Y 0.04fF
C29377 INVX1_LOC_21/A NOR2X1_LOC_536/A 0.13fF
C29378 NAND2X1_LOC_338/B INVX1_LOC_7/A 0.01fF
C29379 INVX1_LOC_2/A NOR2X1_LOC_717/B 0.03fF
C29380 NAND2X1_LOC_549/B INVX1_LOC_234/A 0.01fF
C29381 INVX1_LOC_276/A NAND2X1_LOC_779/a_36_24# 0.00fF
C29382 NOR2X1_LOC_151/Y INVX1_LOC_49/A 0.07fF
C29383 INVX1_LOC_11/A NOR2X1_LOC_357/Y 0.08fF
C29384 INVX1_LOC_117/A INVX1_LOC_198/A -0.01fF
C29385 NAND2X1_LOC_53/Y INVX1_LOC_139/A 0.04fF
C29386 NAND2X1_LOC_693/a_36_24# INVX1_LOC_275/A 0.00fF
C29387 INVX1_LOC_223/A NOR2X1_LOC_552/A 0.01fF
C29388 NOR2X1_LOC_19/B NOR2X1_LOC_514/Y 0.03fF
C29389 NOR2X1_LOC_78/B INVX1_LOC_313/A 0.03fF
C29390 NOR2X1_LOC_89/A NAND2X1_LOC_175/Y 0.07fF
C29391 NOR2X1_LOC_740/Y INVX1_LOC_117/A 0.18fF
C29392 NOR2X1_LOC_65/B INVX1_LOC_49/Y 0.68fF
C29393 INVX1_LOC_98/Y INPUT_1 0.16fF
C29394 INVX1_LOC_59/A NOR2X1_LOC_96/Y 0.12fF
C29395 INVX1_LOC_30/A NAND2X1_LOC_468/B 0.05fF
C29396 INVX1_LOC_1/Y INVX1_LOC_10/A 0.20fF
C29397 INVX1_LOC_240/A NAND2X1_LOC_855/Y 0.00fF
C29398 NAND2X1_LOC_35/Y NOR2X1_LOC_103/a_36_216# 0.01fF
C29399 NOR2X1_LOC_801/B NAND2X1_LOC_761/a_36_24# 0.00fF
C29400 INVX1_LOC_21/A NAND2X1_LOC_93/B 0.03fF
C29401 NOR2X1_LOC_733/Y INVX1_LOC_113/Y 0.00fF
C29402 INVX1_LOC_313/Y INVX1_LOC_179/Y 0.02fF
C29403 INVX1_LOC_31/A INVX1_LOC_46/A 0.03fF
C29404 NOR2X1_LOC_71/Y INVX1_LOC_53/Y 0.05fF
C29405 INVX1_LOC_47/A INVX1_LOC_40/A 0.09fF
C29406 INVX1_LOC_226/Y NOR2X1_LOC_559/a_36_216# 0.00fF
C29407 NOR2X1_LOC_554/B NAND2X1_LOC_819/a_36_24# 0.01fF
C29408 INVX1_LOC_18/A NOR2X1_LOC_683/a_36_216# 0.02fF
C29409 NOR2X1_LOC_584/Y NOR2X1_LOC_638/Y 0.00fF
C29410 NAND2X1_LOC_191/a_36_24# NOR2X1_LOC_331/B 0.01fF
C29411 NOR2X1_LOC_68/A INVX1_LOC_59/Y 0.08fF
C29412 NOR2X1_LOC_428/Y NAND2X1_LOC_639/A 0.04fF
C29413 INVX1_LOC_21/A NAND2X1_LOC_425/Y 0.01fF
C29414 INVX1_LOC_58/A INVX1_LOC_272/A 0.07fF
C29415 INVX1_LOC_299/A NOR2X1_LOC_641/Y 0.03fF
C29416 INVX1_LOC_57/A NAND2X1_LOC_207/B 0.02fF
C29417 NOR2X1_LOC_233/a_36_216# INVX1_LOC_35/Y 0.01fF
C29418 INVX1_LOC_72/A INVX1_LOC_76/A 0.26fF
C29419 INVX1_LOC_40/Y VDD 0.41fF
C29420 NOR2X1_LOC_68/A INVX1_LOC_112/A 0.01fF
C29421 INVX1_LOC_2/A NOR2X1_LOC_151/Y 0.03fF
C29422 NOR2X1_LOC_453/Y NAND2X1_LOC_93/B 0.18fF
C29423 NAND2X1_LOC_554/a_36_24# INVX1_LOC_10/A 0.01fF
C29424 NOR2X1_LOC_103/Y INVX1_LOC_9/A 0.07fF
C29425 NOR2X1_LOC_391/A D_INPUT_0 0.09fF
C29426 INVX1_LOC_23/A NOR2X1_LOC_671/Y 0.03fF
C29427 INVX1_LOC_69/Y NOR2X1_LOC_337/a_36_216# 0.01fF
C29428 NOR2X1_LOC_541/Y INVX1_LOC_9/A 0.01fF
C29429 NOR2X1_LOC_68/A INVX1_LOC_176/A 0.13fF
C29430 INVX1_LOC_53/A NOR2X1_LOC_633/A 0.06fF
C29431 NOR2X1_LOC_15/Y NAND2X1_LOC_802/Y 0.07fF
C29432 NAND2X1_LOC_767/a_36_24# INVX1_LOC_280/A 0.00fF
C29433 NOR2X1_LOC_718/B INVX1_LOC_206/Y 0.06fF
C29434 INVX1_LOC_279/A INVX1_LOC_97/A 0.05fF
C29435 INVX1_LOC_305/Y NOR2X1_LOC_567/B 0.01fF
C29436 INVX1_LOC_28/A NAND2X1_LOC_170/A 0.08fF
C29437 INVX1_LOC_38/Y NOR2X1_LOC_814/A 0.01fF
C29438 NOR2X1_LOC_453/Y NAND2X1_LOC_425/Y 0.17fF
C29439 INVX1_LOC_198/Y INVX1_LOC_76/A 0.52fF
C29440 INVX1_LOC_213/Y INVX1_LOC_78/Y 0.00fF
C29441 INVX1_LOC_21/A NOR2X1_LOC_649/B 0.07fF
C29442 NOR2X1_LOC_793/Y NOR2X1_LOC_809/B 0.02fF
C29443 NAND2X1_LOC_588/B VDD 0.01fF
C29444 INVX1_LOC_90/A INVX1_LOC_279/A 0.08fF
C29445 INVX1_LOC_41/Y INVX1_LOC_20/A 0.04fF
C29446 NOR2X1_LOC_204/a_36_216# INVX1_LOC_59/Y 0.00fF
C29447 NOR2X1_LOC_843/B INVX1_LOC_15/A 0.04fF
C29448 NOR2X1_LOC_561/Y INVX1_LOC_313/Y 0.01fF
C29449 NAND2X1_LOC_783/Y INVX1_LOC_118/A 0.06fF
C29450 NAND2X1_LOC_574/A NOR2X1_LOC_611/a_36_216# 0.01fF
C29451 NAND2X1_LOC_574/A NAND2X1_LOC_218/A 0.01fF
C29452 INVX1_LOC_5/A NOR2X1_LOC_84/B 0.02fF
C29453 NAND2X1_LOC_550/A NAND2X1_LOC_241/a_36_24# 0.00fF
C29454 NOR2X1_LOC_617/Y INVX1_LOC_20/A -0.00fF
C29455 NOR2X1_LOC_773/Y INPUT_0 0.21fF
C29456 INVX1_LOC_111/A INVX1_LOC_46/A 0.02fF
C29457 NAND2X1_LOC_357/B NOR2X1_LOC_528/Y 0.27fF
C29458 NOR2X1_LOC_140/A NAND2X1_LOC_574/A 0.01fF
C29459 NOR2X1_LOC_739/Y NOR2X1_LOC_155/A 0.01fF
C29460 INVX1_LOC_226/A INVX1_LOC_158/Y 0.34fF
C29461 NAND2X1_LOC_593/Y INVX1_LOC_20/A 0.06fF
C29462 INVX1_LOC_33/A INVX1_LOC_95/Y 0.09fF
C29463 NOR2X1_LOC_67/A NOR2X1_LOC_391/Y -0.02fF
C29464 NOR2X1_LOC_552/A INVX1_LOC_149/Y 0.02fF
C29465 NOR2X1_LOC_78/B INVX1_LOC_6/A 0.10fF
C29466 NOR2X1_LOC_802/A INVX1_LOC_186/A 0.07fF
C29467 INVX1_LOC_135/A NAND2X1_LOC_622/a_36_24# 0.00fF
C29468 NOR2X1_LOC_582/Y NAND2X1_LOC_639/A 0.04fF
C29469 NAND2X1_LOC_471/Y NAND2X1_LOC_99/A 0.03fF
C29470 NOR2X1_LOC_433/A NOR2X1_LOC_357/Y 0.07fF
C29471 NAND2X1_LOC_45/Y NOR2X1_LOC_702/a_36_216# 0.02fF
C29472 NOR2X1_LOC_570/B NOR2X1_LOC_631/B 0.01fF
C29473 INVX1_LOC_45/A INVX1_LOC_9/A 0.10fF
C29474 NOR2X1_LOC_568/A INVX1_LOC_9/A 0.07fF
C29475 NOR2X1_LOC_128/B NOR2X1_LOC_19/B 0.00fF
C29476 NAND2X1_LOC_567/Y VDD 0.03fF
C29477 NAND2X1_LOC_308/Y INVX1_LOC_11/Y 0.04fF
C29478 NAND2X1_LOC_660/A INVX1_LOC_91/A 0.16fF
C29479 NOR2X1_LOC_426/Y INVX1_LOC_54/A 0.19fF
C29480 NOR2X1_LOC_763/a_36_216# INVX1_LOC_37/A 0.00fF
C29481 INVX1_LOC_227/A NOR2X1_LOC_216/Y 0.23fF
C29482 NAND2X1_LOC_578/a_36_24# NOR2X1_LOC_662/A 0.01fF
C29483 NOR2X1_LOC_593/Y NOR2X1_LOC_357/Y 0.02fF
C29484 NAND2X1_LOC_567/Y NAND2X1_LOC_800/A 0.03fF
C29485 INVX1_LOC_88/A NAND2X1_LOC_475/Y 0.05fF
C29486 NOR2X1_LOC_299/Y NAND2X1_LOC_863/A 0.05fF
C29487 NOR2X1_LOC_590/A NOR2X1_LOC_197/B 0.08fF
C29488 NAND2X1_LOC_595/a_36_24# NOR2X1_LOC_814/A 0.01fF
C29489 NOR2X1_LOC_643/A INVX1_LOC_63/A 0.00fF
C29490 NOR2X1_LOC_300/Y NAND2X1_LOC_212/Y 0.20fF
C29491 NAND2X1_LOC_799/A INVX1_LOC_84/A 3.53fF
C29492 NAND2X1_LOC_350/A NOR2X1_LOC_697/Y 0.01fF
C29493 NOR2X1_LOC_503/A NAND2X1_LOC_648/A 0.01fF
C29494 NOR2X1_LOC_495/Y NOR2X1_LOC_495/a_36_216# 0.00fF
C29495 INVX1_LOC_36/A INVX1_LOC_92/A 0.20fF
C29496 INVX1_LOC_200/A INVX1_LOC_63/A 0.01fF
C29497 INVX1_LOC_206/Y NOR2X1_LOC_569/Y 0.00fF
C29498 NOR2X1_LOC_318/B NOR2X1_LOC_500/Y 0.01fF
C29499 INVX1_LOC_6/A NAND2X1_LOC_392/Y 0.03fF
C29500 NOR2X1_LOC_332/A INPUT_0 0.35fF
C29501 NOR2X1_LOC_52/B NOR2X1_LOC_357/Y 0.04fF
C29502 INVX1_LOC_71/A INVX1_LOC_9/A 0.33fF
C29503 INVX1_LOC_77/A NOR2X1_LOC_331/B 0.07fF
C29504 INVX1_LOC_85/A INVX1_LOC_139/Y 0.00fF
C29505 NOR2X1_LOC_770/B INVX1_LOC_117/A 0.02fF
C29506 NOR2X1_LOC_384/Y NOR2X1_LOC_88/a_36_216# 0.02fF
C29507 INVX1_LOC_83/A INVX1_LOC_6/A 0.03fF
C29508 INVX1_LOC_286/Y INVX1_LOC_285/A 0.48fF
C29509 INVX1_LOC_40/A INVX1_LOC_95/Y 0.38fF
C29510 NAND2X1_LOC_338/B INVX1_LOC_76/A 0.11fF
C29511 INVX1_LOC_49/A NOR2X1_LOC_709/B 0.03fF
C29512 INVX1_LOC_18/A NOR2X1_LOC_88/Y 0.10fF
C29513 NOR2X1_LOC_742/A NOR2X1_LOC_302/Y 0.04fF
C29514 NAND2X1_LOC_840/a_36_24# INVX1_LOC_33/Y 0.00fF
C29515 NOR2X1_LOC_19/B NAND2X1_LOC_849/A 1.50fF
C29516 INVX1_LOC_90/A NAND2X1_LOC_858/B 0.01fF
C29517 NOR2X1_LOC_503/Y INVX1_LOC_49/Y 0.13fF
C29518 NAND2X1_LOC_342/Y VDD 0.28fF
C29519 NOR2X1_LOC_520/a_36_216# INVX1_LOC_176/A 0.00fF
C29520 NOR2X1_LOC_716/B INVX1_LOC_118/A 0.07fF
C29521 INVX1_LOC_31/A NOR2X1_LOC_68/Y 0.03fF
C29522 NOR2X1_LOC_91/A NAND2X1_LOC_9/Y 0.03fF
C29523 NOR2X1_LOC_318/B INVX1_LOC_10/A 0.20fF
C29524 NOR2X1_LOC_226/A NAND2X1_LOC_633/Y 0.04fF
C29525 NOR2X1_LOC_208/Y INVX1_LOC_92/A 0.07fF
C29526 INVX1_LOC_108/Y NOR2X1_LOC_843/B 0.11fF
C29527 NOR2X1_LOC_739/Y NOR2X1_LOC_833/B 0.06fF
C29528 NOR2X1_LOC_91/A INVX1_LOC_233/A 0.14fF
C29529 NOR2X1_LOC_440/B INVX1_LOC_4/A 0.02fF
C29530 INVX1_LOC_53/A INVX1_LOC_270/A 0.10fF
C29531 INVX1_LOC_41/A NOR2X1_LOC_489/A 0.05fF
C29532 INPUT_0 INVX1_LOC_140/A 0.10fF
C29533 INVX1_LOC_93/Y INVX1_LOC_10/A 0.07fF
C29534 INVX1_LOC_13/A INVX1_LOC_74/A 0.02fF
C29535 INVX1_LOC_18/A INVX1_LOC_84/A 0.18fF
C29536 NOR2X1_LOC_87/B INVX1_LOC_230/A 0.02fF
C29537 INVX1_LOC_2/Y INVX1_LOC_232/A 0.01fF
C29538 NAND2X1_LOC_9/Y INVX1_LOC_23/A 0.19fF
C29539 INVX1_LOC_31/A NOR2X1_LOC_671/Y 0.03fF
C29540 NOR2X1_LOC_191/B INVX1_LOC_285/A 0.18fF
C29541 INVX1_LOC_224/A INVX1_LOC_32/A 0.03fF
C29542 NAND2X1_LOC_560/A INVX1_LOC_309/A 0.00fF
C29543 NAND2X1_LOC_591/a_36_24# INVX1_LOC_186/Y 0.01fF
C29544 NOR2X1_LOC_667/A NOR2X1_LOC_536/A 0.19fF
C29545 INVX1_LOC_233/A INVX1_LOC_23/A 0.08fF
C29546 NOR2X1_LOC_174/A INVX1_LOC_186/A 0.01fF
C29547 INVX1_LOC_11/A INVX1_LOC_32/A 0.20fF
C29548 INVX1_LOC_58/A NAND2X1_LOC_708/Y 0.03fF
C29549 INVX1_LOC_263/A NAND2X1_LOC_472/Y 0.09fF
C29550 INVX1_LOC_248/A NOR2X1_LOC_536/A 0.60fF
C29551 NAND2X1_LOC_859/Y INVX1_LOC_46/A 0.03fF
C29552 INVX1_LOC_24/Y NOR2X1_LOC_334/Y 0.01fF
C29553 INVX1_LOC_64/A NOR2X1_LOC_629/A 0.01fF
C29554 INVX1_LOC_136/A NAND2X1_LOC_81/B 0.28fF
C29555 NOR2X1_LOC_309/Y INVX1_LOC_92/A 0.03fF
C29556 INVX1_LOC_18/A NAND2X1_LOC_651/B 0.03fF
C29557 NAND2X1_LOC_208/B INVX1_LOC_42/A 0.01fF
C29558 NOR2X1_LOC_71/Y NAND2X1_LOC_465/A 0.05fF
C29559 NOR2X1_LOC_703/B INVX1_LOC_29/A 0.03fF
C29560 INVX1_LOC_172/A INVX1_LOC_84/A 0.03fF
C29561 NAND2X1_LOC_740/Y NAND2X1_LOC_724/Y 0.03fF
C29562 NOR2X1_LOC_186/Y INVX1_LOC_50/A 0.07fF
C29563 NAND2X1_LOC_222/A INVX1_LOC_27/A 0.02fF
C29564 NOR2X1_LOC_328/Y NOR2X1_LOC_694/Y 0.00fF
C29565 NAND2X1_LOC_560/A INVX1_LOC_91/A 0.03fF
C29566 NAND2X1_LOC_553/A INVX1_LOC_23/A 0.00fF
C29567 NOR2X1_LOC_338/Y INVX1_LOC_272/A 0.03fF
C29568 NOR2X1_LOC_68/A NOR2X1_LOC_340/A 0.12fF
C29569 INVX1_LOC_103/A NAND2X1_LOC_454/Y 0.07fF
C29570 NOR2X1_LOC_443/Y INVX1_LOC_27/A 0.13fF
C29571 NOR2X1_LOC_741/A NOR2X1_LOC_74/A 0.01fF
C29572 NOR2X1_LOC_798/A INVX1_LOC_23/A 3.27fF
C29573 INVX1_LOC_64/A NAND2X1_LOC_624/B 0.03fF
C29574 NOR2X1_LOC_94/a_36_216# INVX1_LOC_280/A 0.00fF
C29575 NAND2X1_LOC_681/a_36_24# NAND2X1_LOC_782/B 0.01fF
C29576 INVX1_LOC_232/A NAND2X1_LOC_276/a_36_24# 0.06fF
C29577 NOR2X1_LOC_521/Y NOR2X1_LOC_536/A 0.02fF
C29578 NAND2X1_LOC_560/A INVX1_LOC_11/Y 0.03fF
C29579 NOR2X1_LOC_516/Y NAND2X1_LOC_659/A 0.08fF
C29580 NOR2X1_LOC_78/B INVX1_LOC_131/Y 0.07fF
C29581 INVX1_LOC_50/A NAND2X1_LOC_573/Y 0.07fF
C29582 INVX1_LOC_11/A NAND2X1_LOC_175/Y 0.08fF
C29583 NOR2X1_LOC_152/Y INVX1_LOC_49/Y 0.13fF
C29584 NOR2X1_LOC_542/a_36_216# NOR2X1_LOC_814/A 0.00fF
C29585 NOR2X1_LOC_226/A INVX1_LOC_71/Y 0.02fF
C29586 NOR2X1_LOC_363/Y NOR2X1_LOC_366/Y 0.00fF
C29587 INVX1_LOC_54/Y NOR2X1_LOC_831/B 0.16fF
C29588 NAND2X1_LOC_866/B INVX1_LOC_46/A 0.09fF
C29589 NOR2X1_LOC_352/Y NOR2X1_LOC_155/A 0.01fF
C29590 INVX1_LOC_72/A INVX1_LOC_127/Y 0.02fF
C29591 NOR2X1_LOC_92/Y NAND2X1_LOC_464/B 0.07fF
C29592 NOR2X1_LOC_419/Y NAND2X1_LOC_63/Y 0.02fF
C29593 NAND2X1_LOC_840/B INVX1_LOC_291/A 0.02fF
C29594 NOR2X1_LOC_246/Y VDD 0.12fF
C29595 INVX1_LOC_24/A NOR2X1_LOC_67/Y 0.19fF
C29596 INVX1_LOC_279/A INVX1_LOC_38/A 0.43fF
C29597 NOR2X1_LOC_471/Y NOR2X1_LOC_464/Y 0.01fF
C29598 NOR2X1_LOC_516/B INVX1_LOC_274/A 0.04fF
C29599 INVX1_LOC_50/A NAND2X1_LOC_724/A 0.07fF
C29600 INVX1_LOC_87/Y VDD 0.41fF
C29601 INVX1_LOC_64/A NOR2X1_LOC_849/A 0.03fF
C29602 NOR2X1_LOC_638/a_36_216# INVX1_LOC_261/Y 0.00fF
C29603 NOR2X1_LOC_716/B NAND2X1_LOC_63/Y 0.09fF
C29604 NAND2X1_LOC_807/Y INVX1_LOC_46/A 0.03fF
C29605 INVX1_LOC_63/Y INVX1_LOC_19/A 0.03fF
C29606 NAND2X1_LOC_762/a_36_24# INVX1_LOC_15/A 0.00fF
C29607 NOR2X1_LOC_52/B NAND2X1_LOC_489/Y 0.03fF
C29608 INVX1_LOC_18/A INVX1_LOC_15/A 0.14fF
C29609 NAND2X1_LOC_364/A INVX1_LOC_47/Y 0.01fF
C29610 NOR2X1_LOC_561/Y NOR2X1_LOC_506/Y 0.02fF
C29611 NOR2X1_LOC_223/a_36_216# NAND2X1_LOC_425/Y -0.01fF
C29612 INVX1_LOC_25/A INVX1_LOC_14/A 2.92fF
C29613 INVX1_LOC_16/A INVX1_LOC_179/A 0.08fF
C29614 NAND2X1_LOC_12/a_36_24# INVX1_LOC_15/A 0.00fF
C29615 INVX1_LOC_232/A NOR2X1_LOC_608/Y 0.01fF
C29616 INVX1_LOC_136/A INVX1_LOC_4/Y 0.34fF
C29617 NAND2X1_LOC_169/Y INVX1_LOC_93/A 0.05fF
C29618 INVX1_LOC_13/Y NOR2X1_LOC_791/Y 0.01fF
C29619 INVX1_LOC_6/A NOR2X1_LOC_368/Y 0.08fF
C29620 INVX1_LOC_235/Y INVX1_LOC_253/Y 0.63fF
C29621 NOR2X1_LOC_516/B NOR2X1_LOC_820/Y 0.05fF
C29622 INVX1_LOC_11/A NOR2X1_LOC_622/A 0.05fF
C29623 NOR2X1_LOC_749/Y INVX1_LOC_9/A 0.01fF
C29624 NOR2X1_LOC_448/B INVX1_LOC_295/Y 0.05fF
C29625 VDD INVX1_LOC_67/Y 0.21fF
C29626 NOR2X1_LOC_667/A NOR2X1_LOC_661/A 0.07fF
C29627 NOR2X1_LOC_824/A NOR2X1_LOC_291/Y 0.37fF
C29628 NOR2X1_LOC_175/A INVX1_LOC_19/A 0.07fF
C29629 INVX1_LOC_163/A NOR2X1_LOC_663/A 0.03fF
C29630 INVX1_LOC_10/A INVX1_LOC_117/Y 0.01fF
C29631 INVX1_LOC_79/Y INVX1_LOC_78/A 0.06fF
C29632 INVX1_LOC_34/A INVX1_LOC_42/A 0.24fF
C29633 NOR2X1_LOC_433/A INVX1_LOC_32/A 0.02fF
C29634 NAND2X1_LOC_342/Y INVX1_LOC_133/A 0.52fF
C29635 NAND2X1_LOC_6/a_36_24# INVX1_LOC_3/A 0.00fF
C29636 NOR2X1_LOC_74/A INVX1_LOC_12/Y 0.10fF
C29637 NAND2X1_LOC_814/a_36_24# NAND2X1_LOC_453/A 0.00fF
C29638 INVX1_LOC_6/A INVX1_LOC_46/A 0.22fF
C29639 NOR2X1_LOC_593/Y INVX1_LOC_32/A 1.44fF
C29640 NAND2X1_LOC_556/a_36_24# INVX1_LOC_284/A 0.00fF
C29641 INVX1_LOC_316/Y NOR2X1_LOC_662/A 0.03fF
C29642 INVX1_LOC_190/A NOR2X1_LOC_592/B 0.01fF
C29643 NOR2X1_LOC_97/a_36_216# NOR2X1_LOC_865/Y 0.00fF
C29644 INVX1_LOC_181/Y NOR2X1_LOC_278/Y 0.07fF
C29645 INVX1_LOC_27/A NAND2X1_LOC_347/B 0.01fF
C29646 INVX1_LOC_12/Y NOR2X1_LOC_9/Y 0.30fF
C29647 INPUT_1 INVX1_LOC_71/Y 0.09fF
C29648 INVX1_LOC_90/A NOR2X1_LOC_624/B 0.01fF
C29649 NOR2X1_LOC_401/A INVX1_LOC_306/Y 0.01fF
C29650 NOR2X1_LOC_99/B NAND2X1_LOC_85/Y 0.13fF
C29651 INVX1_LOC_151/A INVX1_LOC_32/A 0.01fF
C29652 NAND2X1_LOC_9/Y INVX1_LOC_31/A 0.11fF
C29653 NOR2X1_LOC_846/Y INVX1_LOC_17/A 0.01fF
C29654 INVX1_LOC_233/A INVX1_LOC_31/A 0.07fF
C29655 INVX1_LOC_206/Y NAND2X1_LOC_472/Y 0.07fF
C29656 NOR2X1_LOC_52/B INVX1_LOC_32/A 0.12fF
C29657 NOR2X1_LOC_433/A NAND2X1_LOC_175/Y 1.06fF
C29658 INVX1_LOC_41/A NOR2X1_LOC_334/Y 0.07fF
C29659 INVX1_LOC_70/Y VDD 0.21fF
C29660 INVX1_LOC_33/A INVX1_LOC_271/Y 0.03fF
C29661 INVX1_LOC_36/A INVX1_LOC_53/A 0.20fF
C29662 INVX1_LOC_200/Y NOR2X1_LOC_91/Y 0.00fF
C29663 NOR2X1_LOC_91/A NAND2X1_LOC_866/A 0.02fF
C29664 NOR2X1_LOC_160/B INVX1_LOC_306/Y 0.49fF
C29665 NOR2X1_LOC_357/Y INVX1_LOC_199/A 0.03fF
C29666 INVX1_LOC_21/A INVX1_LOC_256/A 0.12fF
C29667 NAND2X1_LOC_9/Y NOR2X1_LOC_410/a_36_216# 0.00fF
C29668 NAND2X1_LOC_363/B NOR2X1_LOC_500/B 0.07fF
C29669 INVX1_LOC_34/A INVX1_LOC_78/A 0.11fF
C29670 NOR2X1_LOC_455/a_36_216# NOR2X1_LOC_334/Y 0.00fF
C29671 INVX1_LOC_1/Y INVX1_LOC_12/A 0.07fF
C29672 NOR2X1_LOC_261/Y INVX1_LOC_18/A 0.36fF
C29673 INVX1_LOC_1/A INVX1_LOC_14/A 0.91fF
C29674 NOR2X1_LOC_92/Y INVX1_LOC_308/Y 0.03fF
C29675 NAND2X1_LOC_564/B NOR2X1_LOC_89/A 0.00fF
C29676 INVX1_LOC_177/A NAND2X1_LOC_647/B 0.01fF
C29677 NOR2X1_LOC_600/Y NAND2X1_LOC_472/Y 0.23fF
C29678 INVX1_LOC_278/A INVX1_LOC_18/A 0.07fF
C29679 NOR2X1_LOC_91/A NAND2X1_LOC_812/A 0.15fF
C29680 INVX1_LOC_121/A NAND2X1_LOC_259/a_36_24# 0.00fF
C29681 NOR2X1_LOC_772/B INVX1_LOC_30/A 0.01fF
C29682 INVX1_LOC_272/Y INVX1_LOC_289/Y 0.15fF
C29683 NOR2X1_LOC_859/A INVX1_LOC_64/A 0.03fF
C29684 INVX1_LOC_233/Y INVX1_LOC_136/A 2.64fF
C29685 NOR2X1_LOC_798/A INVX1_LOC_31/A 0.05fF
C29686 NAND2X1_LOC_218/B D_INPUT_1 0.08fF
C29687 NOR2X1_LOC_533/Y NAND2X1_LOC_537/Y 0.28fF
C29688 NOR2X1_LOC_178/Y INVX1_LOC_72/A 0.73fF
C29689 INVX1_LOC_132/A INVX1_LOC_50/A 0.07fF
C29690 INVX1_LOC_149/Y NOR2X1_LOC_541/B 0.00fF
C29691 INVX1_LOC_311/A NAND2X1_LOC_93/B 0.07fF
C29692 NOR2X1_LOC_52/B NAND2X1_LOC_175/Y 0.07fF
C29693 INVX1_LOC_83/A NOR2X1_LOC_633/A 0.07fF
C29694 INVX1_LOC_13/Y INVX1_LOC_30/A 0.15fF
C29695 NOR2X1_LOC_65/B INVX1_LOC_34/A 0.15fF
C29696 NOR2X1_LOC_500/A NOR2X1_LOC_790/B 0.32fF
C29697 D_INPUT_1 NOR2X1_LOC_577/Y 0.07fF
C29698 NAND2X1_LOC_703/Y INVX1_LOC_31/A 0.07fF
C29699 NOR2X1_LOC_738/Y NOR2X1_LOC_740/Y 0.04fF
C29700 INVX1_LOC_304/A NOR2X1_LOC_536/A 0.07fF
C29701 INVX1_LOC_60/Y INVX1_LOC_23/Y 0.16fF
C29702 NAND2X1_LOC_231/Y INVX1_LOC_78/A 0.03fF
C29703 NOR2X1_LOC_124/B INVX1_LOC_112/Y 0.03fF
C29704 INVX1_LOC_183/Y INVX1_LOC_29/A 0.01fF
C29705 INVX1_LOC_278/A INVX1_LOC_172/A 0.03fF
C29706 INVX1_LOC_64/A NOR2X1_LOC_617/Y 0.02fF
C29707 NAND2X1_LOC_222/B INPUT_3 0.01fF
C29708 INVX1_LOC_50/A INVX1_LOC_225/A 0.01fF
C29709 NOR2X1_LOC_264/Y INVX1_LOC_57/A 0.21fF
C29710 NOR2X1_LOC_175/A INVX1_LOC_26/Y 0.02fF
C29711 NOR2X1_LOC_536/A NOR2X1_LOC_670/Y 0.02fF
C29712 NOR2X1_LOC_209/Y NOR2X1_LOC_306/a_36_216# 0.00fF
C29713 NOR2X1_LOC_804/B INVX1_LOC_53/A 0.09fF
C29714 INVX1_LOC_64/A NAND2X1_LOC_593/Y 0.03fF
C29715 INVX1_LOC_35/A NOR2X1_LOC_712/B 0.08fF
C29716 INVX1_LOC_11/A INPUT_3 0.06fF
C29717 INVX1_LOC_1/A NOR2X1_LOC_717/Y 0.10fF
C29718 NOR2X1_LOC_721/Y NOR2X1_LOC_814/A 0.02fF
C29719 NOR2X1_LOC_798/A INVX1_LOC_111/A 0.00fF
C29720 NOR2X1_LOC_65/B NAND2X1_LOC_231/Y 0.10fF
C29721 NAND2X1_LOC_381/Y INPUT_3 0.01fF
C29722 INVX1_LOC_33/Y NOR2X1_LOC_111/A 0.05fF
C29723 D_INPUT_1 NOR2X1_LOC_348/B 0.01fF
C29724 NOR2X1_LOC_643/Y INVX1_LOC_5/A 0.01fF
C29725 NOR2X1_LOC_285/Y NAND2X1_LOC_361/Y 0.03fF
C29726 INVX1_LOC_88/A INVX1_LOC_30/A 0.08fF
C29727 INVX1_LOC_95/A NOR2X1_LOC_743/Y 0.00fF
C29728 NOR2X1_LOC_309/Y INVX1_LOC_53/A 0.01fF
C29729 INVX1_LOC_25/A NOR2X1_LOC_612/B 0.42fF
C29730 NOR2X1_LOC_742/A INVX1_LOC_12/A 0.14fF
C29731 NAND2X1_LOC_633/Y INVX1_LOC_118/A 0.07fF
C29732 NAND2X1_LOC_802/A INVX1_LOC_178/A 0.24fF
C29733 INVX1_LOC_16/A NOR2X1_LOC_693/Y 0.07fF
C29734 NOR2X1_LOC_520/B INVX1_LOC_50/Y 0.07fF
C29735 NAND2X1_LOC_149/Y NAND2X1_LOC_161/a_36_24# 0.01fF
C29736 INVX1_LOC_303/A NAND2X1_LOC_63/a_36_24# 0.00fF
C29737 INVX1_LOC_230/Y NAND2X1_LOC_577/A 0.07fF
C29738 NOR2X1_LOC_68/A INVX1_LOC_103/A 0.17fF
C29739 INVX1_LOC_37/A INVX1_LOC_54/A 0.09fF
C29740 NOR2X1_LOC_590/A INVX1_LOC_286/Y 0.10fF
C29741 NOR2X1_LOC_226/A NOR2X1_LOC_591/A 0.03fF
C29742 INVX1_LOC_35/A INVX1_LOC_149/A 0.04fF
C29743 NAND2X1_LOC_567/a_36_24# INVX1_LOC_94/Y 0.00fF
C29744 NAND2X1_LOC_84/Y INVX1_LOC_1/A 0.12fF
C29745 INVX1_LOC_131/Y INVX1_LOC_46/A 0.01fF
C29746 INPUT_0 NOR2X1_LOC_847/A 0.60fF
C29747 NOR2X1_LOC_421/a_36_216# NOR2X1_LOC_561/Y 0.01fF
C29748 INVX1_LOC_224/Y NOR2X1_LOC_719/A 0.01fF
C29749 VDD NOR2X1_LOC_364/A 0.53fF
C29750 NAND2X1_LOC_803/B INVX1_LOC_159/A 0.02fF
C29751 NOR2X1_LOC_92/Y INVX1_LOC_209/Y 0.00fF
C29752 INVX1_LOC_34/A NOR2X1_LOC_215/A 0.02fF
C29753 INVX1_LOC_38/A NOR2X1_LOC_450/A 0.01fF
C29754 INVX1_LOC_5/A INVX1_LOC_266/Y 0.20fF
C29755 NAND2X1_LOC_188/a_36_24# INVX1_LOC_72/A 0.01fF
C29756 INPUT_0 INVX1_LOC_42/A 0.14fF
C29757 NOR2X1_LOC_372/A NOR2X1_LOC_372/Y 0.10fF
C29758 INVX1_LOC_190/A NOR2X1_LOC_449/A 0.15fF
C29759 NOR2X1_LOC_473/B INVX1_LOC_94/Y 0.01fF
C29760 D_INPUT_1 INVX1_LOC_22/A 1.12fF
C29761 NOR2X1_LOC_68/A INVX1_LOC_292/A 0.10fF
C29762 NOR2X1_LOC_471/Y NOR2X1_LOC_457/B 0.07fF
C29763 NOR2X1_LOC_178/Y NAND2X1_LOC_338/B 0.02fF
C29764 NOR2X1_LOC_331/B INVX1_LOC_9/A 0.03fF
C29765 NOR2X1_LOC_589/A INVX1_LOC_270/Y 1.57fF
C29766 NOR2X1_LOC_78/B NOR2X1_LOC_109/Y 0.04fF
C29767 NOR2X1_LOC_91/A NOR2X1_LOC_700/Y 0.07fF
C29768 NOR2X1_LOC_791/Y INVX1_LOC_168/A 0.23fF
C29769 INVX1_LOC_30/A NOR2X1_LOC_500/B 0.01fF
C29770 NOR2X1_LOC_209/Y NOR2X1_LOC_590/Y 0.05fF
C29771 NOR2X1_LOC_231/B NAND2X1_LOC_364/A 0.02fF
C29772 NOR2X1_LOC_590/A INVX1_LOC_159/A 0.01fF
C29773 INVX1_LOC_91/A INVX1_LOC_29/A 0.33fF
C29774 INVX1_LOC_28/A INVX1_LOC_165/A 0.03fF
C29775 INVX1_LOC_224/Y INVX1_LOC_7/A 0.04fF
C29776 NOR2X1_LOC_169/B NOR2X1_LOC_568/A 0.01fF
C29777 INVX1_LOC_230/Y NAND2X1_LOC_656/A 0.10fF
C29778 INVX1_LOC_37/A NOR2X1_LOC_430/a_36_216# 0.00fF
C29779 NOR2X1_LOC_318/B INVX1_LOC_12/A 0.07fF
C29780 NAND2X1_LOC_348/A NOR2X1_LOC_38/B 0.79fF
C29781 VDD INVX1_LOC_285/A 2.58fF
C29782 NOR2X1_LOC_84/Y NAND2X1_LOC_75/a_36_24# 0.06fF
C29783 NOR2X1_LOC_468/Y NOR2X1_LOC_392/B 0.01fF
C29784 INVX1_LOC_269/Y INVX1_LOC_33/A 0.08fF
C29785 VDD INVX1_LOC_265/Y 0.28fF
C29786 NOR2X1_LOC_9/a_36_216# INVX1_LOC_63/A 0.02fF
C29787 INVX1_LOC_131/A INVX1_LOC_78/A 0.39fF
C29788 NOR2X1_LOC_602/B NOR2X1_LOC_743/Y 0.03fF
C29789 NOR2X1_LOC_45/B INVX1_LOC_102/A 0.07fF
C29790 INVX1_LOC_105/A NOR2X1_LOC_45/Y 1.04fF
C29791 VDD NOR2X1_LOC_814/A 2.53fF
C29792 NAND2X1_LOC_96/A NOR2X1_LOC_461/B 0.06fF
C29793 INVX1_LOC_93/Y INVX1_LOC_12/A 0.07fF
C29794 INVX1_LOC_247/Y NOR2X1_LOC_703/B 0.00fF
C29795 NOR2X1_LOC_177/Y INVX1_LOC_54/A 0.45fF
C29796 INVX1_LOC_28/A NOR2X1_LOC_693/Y 0.07fF
C29797 NAND2X1_LOC_51/B NAND2X1_LOC_470/B 0.91fF
C29798 INVX1_LOC_99/Y NOR2X1_LOC_540/a_36_216# 0.00fF
C29799 INVX1_LOC_285/Y NAND2X1_LOC_647/B 0.27fF
C29800 NAND2X1_LOC_549/Y INVX1_LOC_234/A 0.01fF
C29801 NOR2X1_LOC_384/Y NOR2X1_LOC_522/Y 0.01fF
C29802 INVX1_LOC_75/A NOR2X1_LOC_34/Y 0.03fF
C29803 INVX1_LOC_22/A NOR2X1_LOC_652/Y 0.26fF
C29804 D_INPUT_3 NAND2X1_LOC_219/B 0.50fF
C29805 INVX1_LOC_11/A NOR2X1_LOC_337/a_36_216# 0.00fF
C29806 NAND2X1_LOC_794/B NAND2X1_LOC_170/A 0.05fF
C29807 INPUT_0 INVX1_LOC_78/A 10.15fF
C29808 NOR2X1_LOC_169/B INVX1_LOC_71/A 0.01fF
C29809 INVX1_LOC_11/A INVX1_LOC_158/A 0.30fF
C29810 INVX1_LOC_303/A INVX1_LOC_30/A 0.02fF
C29811 NAND2X1_LOC_842/B INVX1_LOC_23/A 0.07fF
C29812 NOR2X1_LOC_720/B NAND2X1_LOC_114/B 0.00fF
C29813 NAND2X1_LOC_350/A NAND2X1_LOC_453/a_36_24# 0.01fF
C29814 NAND2X1_LOC_729/Y NAND2X1_LOC_739/B 0.45fF
C29815 INVX1_LOC_12/A INVX1_LOC_139/A 0.19fF
C29816 NOR2X1_LOC_455/Y INVX1_LOC_313/Y 0.00fF
C29817 NAND2X1_LOC_773/Y INVX1_LOC_40/A 0.78fF
C29818 INVX1_LOC_286/Y NAND2X1_LOC_354/B 0.03fF
C29819 NOR2X1_LOC_405/A INVX1_LOC_47/Y 0.10fF
C29820 NOR2X1_LOC_722/Y INVX1_LOC_113/Y 0.00fF
C29821 INVX1_LOC_27/A NAND2X1_LOC_159/a_36_24# 0.00fF
C29822 NOR2X1_LOC_65/B INPUT_0 0.10fF
C29823 NOR2X1_LOC_831/B NAND2X1_LOC_656/B 0.01fF
C29824 INVX1_LOC_237/Y INVX1_LOC_72/A 1.33fF
C29825 NAND2X1_LOC_763/B NAND2X1_LOC_59/B 0.23fF
C29826 NAND2X1_LOC_21/Y INVX1_LOC_18/A 0.51fF
C29827 NAND2X1_LOC_287/B NAND2X1_LOC_807/a_36_24# 0.00fF
C29828 INVX1_LOC_74/A INVX1_LOC_32/A 0.48fF
C29829 NOR2X1_LOC_89/A NAND2X1_LOC_804/Y 0.02fF
C29830 INVX1_LOC_2/A NOR2X1_LOC_644/B 0.02fF
C29831 NOR2X1_LOC_439/B NOR2X1_LOC_678/A 0.01fF
C29832 NOR2X1_LOC_681/Y NOR2X1_LOC_48/B 0.05fF
C29833 INVX1_LOC_37/A NOR2X1_LOC_48/B 0.30fF
C29834 NAND2X1_LOC_647/B NOR2X1_LOC_137/B 0.00fF
C29835 INVX1_LOC_226/Y NOR2X1_LOC_82/A 0.13fF
C29836 INVX1_LOC_298/Y INVX1_LOC_91/A 0.02fF
C29837 NOR2X1_LOC_420/Y INVX1_LOC_90/A 0.01fF
C29838 NOR2X1_LOC_141/a_36_216# NAND2X1_LOC_454/Y 0.01fF
C29839 NAND2X1_LOC_374/Y NOR2X1_LOC_372/A -0.03fF
C29840 INVX1_LOC_75/A NOR2X1_LOC_678/A 0.03fF
C29841 INVX1_LOC_289/Y INVX1_LOC_10/A 0.10fF
C29842 D_INPUT_1 INVX1_LOC_100/A 0.12fF
C29843 NOR2X1_LOC_486/Y INVX1_LOC_271/Y 0.07fF
C29844 NOR2X1_LOC_607/Y NOR2X1_LOC_577/Y 0.03fF
C29845 INVX1_LOC_181/Y NOR2X1_LOC_561/a_36_216# 0.00fF
C29846 INVX1_LOC_41/Y NAND2X1_LOC_833/a_36_24# 0.00fF
C29847 NOR2X1_LOC_488/Y NOR2X1_LOC_369/Y 0.05fF
C29848 INVX1_LOC_63/A INVX1_LOC_92/A 0.09fF
C29849 INVX1_LOC_11/A GATE_662 0.07fF
C29850 NOR2X1_LOC_559/B NOR2X1_LOC_520/B 0.19fF
C29851 NOR2X1_LOC_454/Y INVX1_LOC_295/A 0.11fF
C29852 INVX1_LOC_91/A NOR2X1_LOC_318/a_36_216# 0.01fF
C29853 INVX1_LOC_152/Y INPUT_0 0.01fF
C29854 INVX1_LOC_25/A INVX1_LOC_48/A 0.08fF
C29855 INVX1_LOC_45/A INVX1_LOC_179/Y 0.04fF
C29856 INVX1_LOC_39/A NOR2X1_LOC_120/a_36_216# 0.01fF
C29857 INVX1_LOC_269/A D_INPUT_0 0.24fF
C29858 INVX1_LOC_49/Y INVX1_LOC_291/A 0.16fF
C29859 INVX1_LOC_36/A NOR2X1_LOC_78/B 2.89fF
C29860 INVX1_LOC_34/A NOR2X1_LOC_152/Y 0.03fF
C29861 INVX1_LOC_24/A INVX1_LOC_104/A 0.07fF
C29862 INVX1_LOC_292/A NOR2X1_LOC_570/Y 0.05fF
C29863 NOR2X1_LOC_232/Y D_INPUT_0 0.16fF
C29864 NOR2X1_LOC_45/B INVX1_LOC_296/Y 0.03fF
C29865 INVX1_LOC_5/A INVX1_LOC_42/Y 0.01fF
C29866 NOR2X1_LOC_273/a_36_216# INVX1_LOC_266/Y 0.01fF
C29867 INVX1_LOC_34/A NAND2X1_LOC_193/a_36_24# 0.00fF
C29868 INVX1_LOC_49/Y NAND2X1_LOC_802/Y 0.12fF
C29869 NOR2X1_LOC_80/Y INVX1_LOC_46/A 0.01fF
C29870 INVX1_LOC_233/A INVX1_LOC_6/A 0.14fF
C29871 INVX1_LOC_34/A INVX1_LOC_113/Y 0.03fF
C29872 NOR2X1_LOC_468/Y INVX1_LOC_90/A 0.06fF
C29873 NOR2X1_LOC_218/A NAND2X1_LOC_656/Y 0.01fF
C29874 NAND2X1_LOC_703/Y NAND2X1_LOC_807/Y 0.02fF
C29875 INVX1_LOC_50/A NAND2X1_LOC_642/Y 0.07fF
C29876 NOR2X1_LOC_829/Y INVX1_LOC_11/Y 0.00fF
C29877 NAND2X1_LOC_190/Y INVX1_LOC_90/A 0.01fF
C29878 NOR2X1_LOC_693/Y NOR2X1_LOC_253/Y 0.06fF
C29879 NOR2X1_LOC_793/A NOR2X1_LOC_356/A 0.03fF
C29880 INVX1_LOC_12/A INVX1_LOC_117/Y 0.03fF
C29881 NAND2X1_LOC_807/B NOR2X1_LOC_743/Y 0.14fF
C29882 NOR2X1_LOC_295/Y NOR2X1_LOC_772/Y 0.25fF
C29883 NOR2X1_LOC_591/Y NOR2X1_LOC_577/Y 0.03fF
C29884 NOR2X1_LOC_83/Y NOR2X1_LOC_81/Y 0.12fF
C29885 NOR2X1_LOC_230/Y NOR2X1_LOC_589/A 0.01fF
C29886 NOR2X1_LOC_520/B NOR2X1_LOC_6/B 0.05fF
C29887 INVX1_LOC_41/A NOR2X1_LOC_718/B 0.02fF
C29888 INVX1_LOC_41/Y NAND2X1_LOC_850/Y 0.02fF
C29889 NAND2X1_LOC_557/a_36_24# INVX1_LOC_309/A 0.00fF
C29890 NOR2X1_LOC_78/B NOR2X1_LOC_208/Y 0.07fF
C29891 NAND2X1_LOC_231/Y NOR2X1_LOC_152/Y 0.10fF
C29892 INVX1_LOC_45/A NOR2X1_LOC_561/Y 0.08fF
C29893 INVX1_LOC_36/A NAND2X1_LOC_392/Y 0.03fF
C29894 INVX1_LOC_224/Y INVX1_LOC_76/A 0.07fF
C29895 INVX1_LOC_21/A INVX1_LOC_69/Y 0.07fF
C29896 NOR2X1_LOC_311/Y NOR2X1_LOC_109/Y 0.02fF
C29897 INVX1_LOC_270/A INVX1_LOC_46/A 0.28fF
C29898 INVX1_LOC_45/Y INVX1_LOC_16/A 4.20fF
C29899 NOR2X1_LOC_267/A NAND2X1_LOC_392/Y 0.37fF
C29900 INVX1_LOC_90/A NOR2X1_LOC_389/A 0.04fF
C29901 INVX1_LOC_39/A NOR2X1_LOC_392/a_36_216# 0.00fF
C29902 NOR2X1_LOC_160/B NOR2X1_LOC_356/A 0.07fF
C29903 INVX1_LOC_37/A NOR2X1_LOC_836/A 0.10fF
C29904 NAND2X1_LOC_557/a_36_24# INVX1_LOC_91/A 0.01fF
C29905 INVX1_LOC_215/A NAND2X1_LOC_198/B 0.10fF
C29906 INVX1_LOC_17/A INVX1_LOC_73/A 0.03fF
C29907 INVX1_LOC_295/A NAND2X1_LOC_387/a_36_24# 0.01fF
C29908 INVX1_LOC_36/A INVX1_LOC_83/A 0.30fF
C29909 NOR2X1_LOC_389/B NOR2X1_LOC_389/A 0.33fF
C29910 INVX1_LOC_14/A NOR2X1_LOC_188/A 0.06fF
C29911 NOR2X1_LOC_524/Y NOR2X1_LOC_473/B 0.08fF
C29912 NOR2X1_LOC_773/Y NAND2X1_LOC_811/Y 0.02fF
C29913 INVX1_LOC_143/A INVX1_LOC_104/A 0.00fF
C29914 NOR2X1_LOC_78/B NOR2X1_LOC_309/Y 0.03fF
C29915 NOR2X1_LOC_67/A NOR2X1_LOC_6/B 0.07fF
C29916 NOR2X1_LOC_561/Y INVX1_LOC_71/A 0.17fF
C29917 INVX1_LOC_232/Y NAND2X1_LOC_563/Y 0.19fF
C29918 NAND2X1_LOC_254/Y NAND2X1_LOC_489/Y 3.04fF
C29919 NOR2X1_LOC_68/A INVX1_LOC_120/A 0.22fF
C29920 INVX1_LOC_30/A INVX1_LOC_244/A 0.06fF
C29921 INVX1_LOC_7/A INVX1_LOC_71/A 0.02fF
C29922 INVX1_LOC_34/A NAND2X1_LOC_859/B 0.01fF
C29923 NOR2X1_LOC_160/B NOR2X1_LOC_74/A 0.29fF
C29924 INVX1_LOC_46/A NOR2X1_LOC_109/Y 0.10fF
C29925 NOR2X1_LOC_177/Y NOR2X1_LOC_438/Y 0.02fF
C29926 NOR2X1_LOC_84/B INVX1_LOC_42/A 0.02fF
C29927 NOR2X1_LOC_304/Y NOR2X1_LOC_305/Y 0.02fF
C29928 INVX1_LOC_279/A INVX1_LOC_33/A 0.07fF
C29929 INVX1_LOC_135/A INVX1_LOC_77/A 0.10fF
C29930 NOR2X1_LOC_643/Y NOR2X1_LOC_332/A 0.03fF
C29931 NOR2X1_LOC_160/B NOR2X1_LOC_9/Y 0.26fF
C29932 INVX1_LOC_60/Y INVX1_LOC_232/A 0.03fF
C29933 INVX1_LOC_209/Y NOR2X1_LOC_299/Y 0.03fF
C29934 NOR2X1_LOC_493/A INVX1_LOC_9/A 0.04fF
C29935 NAND2X1_LOC_564/B NOR2X1_LOC_52/B 0.07fF
C29936 INVX1_LOC_295/A INVX1_LOC_77/A 0.06fF
C29937 NAND2X1_LOC_656/Y INVX1_LOC_155/Y 0.01fF
C29938 NAND2X1_LOC_866/A NAND2X1_LOC_866/B 0.02fF
C29939 INVX1_LOC_177/Y NOR2X1_LOC_216/Y 0.27fF
C29940 INVX1_LOC_45/Y INVX1_LOC_28/A 0.05fF
C29941 NOR2X1_LOC_831/B NAND2X1_LOC_286/B 0.01fF
C29942 NOR2X1_LOC_632/Y INVX1_LOC_96/Y 0.24fF
C29943 NOR2X1_LOC_590/A NOR2X1_LOC_337/Y 0.04fF
C29944 INVX1_LOC_45/A INVX1_LOC_303/Y 0.01fF
C29945 NOR2X1_LOC_701/a_36_216# NAND2X1_LOC_852/Y 0.16fF
C29946 NOR2X1_LOC_468/Y NOR2X1_LOC_92/a_36_216# 0.00fF
C29947 INPUT_0 NOR2X1_LOC_554/B 0.16fF
C29948 NAND2X1_LOC_341/A NOR2X1_LOC_222/Y 0.01fF
C29949 INVX1_LOC_191/Y NOR2X1_LOC_583/a_36_216# 0.00fF
C29950 INVX1_LOC_227/Y NOR2X1_LOC_188/A 0.01fF
C29951 NOR2X1_LOC_669/Y NOR2X1_LOC_305/Y 0.13fF
C29952 NAND2X1_LOC_802/A INVX1_LOC_140/A 0.09fF
C29953 NOR2X1_LOC_91/A INVX1_LOC_119/Y 0.02fF
C29954 NAND2X1_LOC_803/B NOR2X1_LOC_56/Y 0.02fF
C29955 NOR2X1_LOC_647/A INVX1_LOC_84/A 0.20fF
C29956 INVX1_LOC_41/Y INVX1_LOC_282/A 0.00fF
C29957 INVX1_LOC_53/A NOR2X1_LOC_435/A 0.01fF
C29958 NOR2X1_LOC_168/Y NOR2X1_LOC_548/A 0.01fF
C29959 NOR2X1_LOC_75/Y NAND2X1_LOC_212/Y 0.02fF
C29960 INVX1_LOC_269/A NOR2X1_LOC_266/B 0.01fF
C29961 INVX1_LOC_64/A INVX1_LOC_185/A 0.03fF
C29962 INVX1_LOC_32/A NAND2X1_LOC_254/Y 2.90fF
C29963 NOR2X1_LOC_202/Y INVX1_LOC_77/A 0.01fF
C29964 NOR2X1_LOC_295/Y NOR2X1_LOC_389/B 0.02fF
C29965 NOR2X1_LOC_103/Y INVX1_LOC_76/A 0.09fF
C29966 NOR2X1_LOC_553/Y INVX1_LOC_22/A 0.03fF
C29967 INVX1_LOC_33/A INVX1_LOC_182/Y 0.03fF
C29968 INPUT_3 INVX1_LOC_74/A 0.44fF
C29969 NAND2X1_LOC_198/B INVX1_LOC_286/A 0.10fF
C29970 NOR2X1_LOC_590/A NOR2X1_LOC_56/Y 0.08fF
C29971 INVX1_LOC_36/A NOR2X1_LOC_311/Y 0.07fF
C29972 NOR2X1_LOC_82/A INVX1_LOC_178/Y 0.02fF
C29973 INVX1_LOC_247/Y INVX1_LOC_91/A 0.02fF
C29974 INVX1_LOC_226/Y NOR2X1_LOC_236/a_36_216# 0.00fF
C29975 INVX1_LOC_89/A INVX1_LOC_196/A 0.03fF
C29976 INVX1_LOC_24/A INVX1_LOC_206/Y 0.03fF
C29977 NAND2X1_LOC_803/B VDD 0.61fF
C29978 INVX1_LOC_222/Y NOR2X1_LOC_641/Y 0.00fF
C29979 NOR2X1_LOC_667/Y INVX1_LOC_20/A 0.04fF
C29980 INVX1_LOC_200/A NAND2X1_LOC_721/A 0.07fF
C29981 NOR2X1_LOC_791/B NOR2X1_LOC_78/A 0.03fF
C29982 NOR2X1_LOC_615/Y VDD 0.12fF
C29983 NAND2X1_LOC_563/A D_INPUT_0 0.02fF
C29984 INVX1_LOC_57/A NOR2X1_LOC_662/A 0.01fF
C29985 NOR2X1_LOC_798/A NOR2X1_LOC_79/A 0.01fF
C29986 INVX1_LOC_24/A INVX1_LOC_86/Y 0.53fF
C29987 NAND2X1_LOC_350/A INVX1_LOC_37/A 0.04fF
C29988 NOR2X1_LOC_136/Y NOR2X1_LOC_106/A 0.00fF
C29989 NOR2X1_LOC_232/Y NAND2X1_LOC_848/A 0.01fF
C29990 NOR2X1_LOC_216/Y INVX1_LOC_104/A 0.42fF
C29991 NOR2X1_LOC_590/A INVX1_LOC_146/Y 0.02fF
C29992 NAND2X1_LOC_190/Y INVX1_LOC_38/A 0.01fF
C29993 NOR2X1_LOC_590/A VDD 3.46fF
C29994 NOR2X1_LOC_510/Y NOR2X1_LOC_364/A 0.15fF
C29995 INVX1_LOC_90/A NOR2X1_LOC_220/A 0.55fF
C29996 INVX1_LOC_53/A INVX1_LOC_63/A 0.43fF
C29997 NAND2X1_LOC_348/A NOR2X1_LOC_844/A 0.05fF
C29998 INVX1_LOC_286/Y NAND2X1_LOC_650/B -0.02fF
C29999 NOR2X1_LOC_322/Y NOR2X1_LOC_315/Y 0.00fF
C30000 INVX1_LOC_45/A INVX1_LOC_76/A 0.33fF
C30001 NAND2X1_LOC_745/a_36_24# NAND2X1_LOC_637/Y 0.00fF
C30002 NOR2X1_LOC_71/Y INVX1_LOC_16/A 0.03fF
C30003 NOR2X1_LOC_91/A INVX1_LOC_284/A 0.04fF
C30004 INVX1_LOC_22/Y VDD 0.50fF
C30005 NOR2X1_LOC_220/A NOR2X1_LOC_389/B 0.06fF
C30006 INVX1_LOC_174/A NAND2X1_LOC_639/A 0.80fF
C30007 INVX1_LOC_183/A INVX1_LOC_42/A 0.01fF
C30008 NAND2X1_LOC_198/B INVX1_LOC_95/A 0.01fF
C30009 INVX1_LOC_81/A NOR2X1_LOC_78/A 0.03fF
C30010 INVX1_LOC_202/A NOR2X1_LOC_269/Y 0.01fF
C30011 NAND2X1_LOC_647/B INVX1_LOC_4/Y 0.02fF
C30012 NOR2X1_LOC_848/Y INVX1_LOC_9/A 0.04fF
C30013 NOR2X1_LOC_751/Y NOR2X1_LOC_35/Y 0.20fF
C30014 NOR2X1_LOC_89/A NAND2X1_LOC_97/a_36_24# 0.00fF
C30015 NAND2X1_LOC_856/A INVX1_LOC_76/A 0.06fF
C30016 INVX1_LOC_11/A NOR2X1_LOC_261/A 0.02fF
C30017 NAND2X1_LOC_374/Y NAND2X1_LOC_560/A 0.02fF
C30018 INVX1_LOC_36/A INVX1_LOC_46/A 0.24fF
C30019 NAND2X1_LOC_223/A NOR2X1_LOC_38/B 0.03fF
C30020 NOR2X1_LOC_516/B NOR2X1_LOC_356/A 0.12fF
C30021 INVX1_LOC_90/A NOR2X1_LOC_548/Y 0.98fF
C30022 NOR2X1_LOC_128/B NAND2X1_LOC_125/a_36_24# 0.02fF
C30023 NOR2X1_LOC_83/Y NOR2X1_LOC_709/A 0.01fF
C30024 NOR2X1_LOC_331/Y NOR2X1_LOC_331/B 0.07fF
C30025 INVX1_LOC_23/A INVX1_LOC_284/A 0.07fF
C30026 INVX1_LOC_203/A NOR2X1_LOC_291/a_36_216# 0.01fF
C30027 NOR2X1_LOC_497/Y INVX1_LOC_22/A 0.80fF
C30028 NOR2X1_LOC_389/A INVX1_LOC_38/A 0.01fF
C30029 INVX1_LOC_111/Y NOR2X1_LOC_188/A 0.02fF
C30030 NOR2X1_LOC_391/A INPUT_1 0.03fF
C30031 NOR2X1_LOC_504/Y NOR2X1_LOC_387/A 0.00fF
C30032 INVX1_LOC_8/A INVX1_LOC_91/A 0.19fF
C30033 NAND2X1_LOC_112/Y NOR2X1_LOC_111/Y 0.10fF
C30034 NOR2X1_LOC_238/Y NAND2X1_LOC_244/A 0.01fF
C30035 NOR2X1_LOC_237/Y NOR2X1_LOC_368/Y 0.05fF
C30036 NOR2X1_LOC_791/A INVX1_LOC_12/Y 0.21fF
C30037 NAND2X1_LOC_399/a_36_24# INVX1_LOC_91/A 0.01fF
C30038 INVX1_LOC_5/A INVX1_LOC_19/A 1.23fF
C30039 INVX1_LOC_71/A INVX1_LOC_76/A 0.24fF
C30040 INVX1_LOC_271/Y NOR2X1_LOC_471/a_36_216# 0.01fF
C30041 NOR2X1_LOC_383/B NOR2X1_LOC_801/B 0.01fF
C30042 NAND2X1_LOC_569/a_36_24# INVX1_LOC_280/A 0.01fF
C30043 INVX1_LOC_208/A NOR2X1_LOC_74/A 0.02fF
C30044 INVX1_LOC_290/A NOR2X1_LOC_163/Y 0.05fF
C30045 INVX1_LOC_196/A NOR2X1_LOC_703/Y 0.01fF
C30046 NOR2X1_LOC_557/Y NAND2X1_LOC_674/a_36_24# 0.06fF
C30047 NOR2X1_LOC_208/Y INVX1_LOC_46/A 0.08fF
C30048 NOR2X1_LOC_802/A NOR2X1_LOC_78/A 0.07fF
C30049 INVX1_LOC_174/A NAND2X1_LOC_93/B 0.12fF
C30050 INVX1_LOC_47/A INVX1_LOC_89/A 0.01fF
C30051 NOR2X1_LOC_401/a_36_216# INVX1_LOC_286/A 0.00fF
C30052 NOR2X1_LOC_361/B INVX1_LOC_285/A 0.17fF
C30053 INVX1_LOC_134/A NOR2X1_LOC_445/B 0.17fF
C30054 NOR2X1_LOC_237/Y INVX1_LOC_46/A 0.29fF
C30055 INVX1_LOC_269/A INVX1_LOC_5/Y 0.01fF
C30056 NOR2X1_LOC_798/A NOR2X1_LOC_633/A 0.02fF
C30057 NAND2X1_LOC_832/Y NAND2X1_LOC_479/Y 0.03fF
C30058 INVX1_LOC_28/A NOR2X1_LOC_71/Y 0.07fF
C30059 NOR2X1_LOC_441/Y NOR2X1_LOC_743/Y 0.02fF
C30060 NOR2X1_LOC_780/B NAND2X1_LOC_782/B 0.10fF
C30061 INVX1_LOC_174/A NAND2X1_LOC_425/Y 0.79fF
C30062 NAND2X1_LOC_337/B NAND2X1_LOC_288/A 0.04fF
C30063 NOR2X1_LOC_160/B NOR2X1_LOC_865/Y 0.09fF
C30064 INVX1_LOC_62/Y INVX1_LOC_38/A 0.15fF
C30065 INPUT_5 NOR2X1_LOC_21/a_36_216# 0.00fF
C30066 INVX1_LOC_31/A NAND2X1_LOC_243/B 0.02fF
C30067 INVX1_LOC_286/A INVX1_LOC_53/Y 0.07fF
C30068 INVX1_LOC_271/Y NOR2X1_LOC_748/A 0.10fF
C30069 NOR2X1_LOC_589/A INVX1_LOC_126/Y 0.04fF
C30070 INVX1_LOC_21/A NOR2X1_LOC_89/A 2.21fF
C30071 NOR2X1_LOC_160/B NOR2X1_LOC_243/B 0.18fF
C30072 NOR2X1_LOC_596/A INVX1_LOC_38/A 0.12fF
C30073 NOR2X1_LOC_791/Y NOR2X1_LOC_76/B 0.06fF
C30074 INVX1_LOC_58/A NOR2X1_LOC_409/B 0.01fF
C30075 NAND2X1_LOC_354/B VDD 0.18fF
C30076 INVX1_LOC_185/Y NAND2X1_LOC_650/B 0.01fF
C30077 INVX1_LOC_53/A NAND2X1_LOC_452/Y 0.01fF
C30078 INVX1_LOC_150/Y NAND2X1_LOC_475/Y 0.22fF
C30079 NOR2X1_LOC_226/A INVX1_LOC_187/A 0.02fF
C30080 INVX1_LOC_89/A NOR2X1_LOC_785/a_36_216# 0.00fF
C30081 NOR2X1_LOC_67/A NOR2X1_LOC_124/A 0.02fF
C30082 NAND2X1_LOC_354/B NAND2X1_LOC_800/A 1.06fF
C30083 NOR2X1_LOC_764/Y NAND2X1_LOC_51/B 0.01fF
C30084 NOR2X1_LOC_309/Y INVX1_LOC_46/A 0.12fF
C30085 INVX1_LOC_93/Y NOR2X1_LOC_566/Y 0.30fF
C30086 NOR2X1_LOC_646/A NOR2X1_LOC_78/A 0.06fF
C30087 INVX1_LOC_41/A NAND2X1_LOC_472/Y 0.03fF
C30088 NOR2X1_LOC_97/A INVX1_LOC_148/Y 0.17fF
C30089 INVX1_LOC_289/Y INVX1_LOC_12/A 0.05fF
C30090 INVX1_LOC_13/A NOR2X1_LOC_557/A 0.00fF
C30091 NOR2X1_LOC_45/B NAND2X1_LOC_662/Y 0.10fF
C30092 INVX1_LOC_31/A INVX1_LOC_119/Y 0.01fF
C30093 INVX1_LOC_21/A NOR2X1_LOC_170/A 0.01fF
C30094 INVX1_LOC_304/Y NAND2X1_LOC_721/A 0.03fF
C30095 NAND2X1_LOC_739/a_36_24# INVX1_LOC_231/A 0.00fF
C30096 NAND2X1_LOC_337/B INVX1_LOC_19/A 0.07fF
C30097 INVX1_LOC_95/A INVX1_LOC_53/Y 0.27fF
C30098 NOR2X1_LOC_840/Y NOR2X1_LOC_858/A 0.12fF
C30099 NOR2X1_LOC_538/B INVX1_LOC_106/A 0.00fF
C30100 D_INPUT_6 INVX1_LOC_15/A 0.26fF
C30101 INVX1_LOC_226/Y INVX1_LOC_59/Y 0.09fF
C30102 INVX1_LOC_276/Y VDD 0.26fF
C30103 INVX1_LOC_70/Y NAND2X1_LOC_573/A 0.38fF
C30104 NOR2X1_LOC_82/A INVX1_LOC_12/A 0.10fF
C30105 NOR2X1_LOC_388/Y INVX1_LOC_9/A 0.02fF
C30106 INVX1_LOC_276/A NAND2X1_LOC_687/a_36_24# 0.00fF
C30107 INVX1_LOC_276/Y NAND2X1_LOC_800/A 0.20fF
C30108 NOR2X1_LOC_265/a_36_216# NAND2X1_LOC_650/B 0.01fF
C30109 NAND2X1_LOC_819/Y VDD 0.01fF
C30110 NOR2X1_LOC_590/A INVX1_LOC_133/A 0.03fF
C30111 INVX1_LOC_226/Y INVX1_LOC_176/A 0.03fF
C30112 NOR2X1_LOC_848/Y NOR2X1_LOC_861/Y 0.01fF
C30113 NAND2X1_LOC_842/B INVX1_LOC_6/A 0.74fF
C30114 INVX1_LOC_230/Y NOR2X1_LOC_671/a_36_216# 0.02fF
C30115 INVX1_LOC_279/A NOR2X1_LOC_486/Y 0.01fF
C30116 NOR2X1_LOC_488/Y VDD 0.48fF
C30117 NOR2X1_LOC_210/A INVX1_LOC_115/A 0.02fF
C30118 INVX1_LOC_5/A INVX1_LOC_26/Y 0.12fF
C30119 NOR2X1_LOC_103/Y INVX1_LOC_127/Y 0.00fF
C30120 INVX1_LOC_31/A INVX1_LOC_284/A 0.07fF
C30121 INVX1_LOC_30/A INVX1_LOC_272/A 0.08fF
C30122 NAND2X1_LOC_812/A NAND2X1_LOC_810/B 0.01fF
C30123 INVX1_LOC_34/A NAND2X1_LOC_802/Y 0.07fF
C30124 NAND2X1_LOC_35/Y NAND2X1_LOC_464/B 0.03fF
C30125 NOR2X1_LOC_272/Y INVX1_LOC_23/Y 0.10fF
C30126 NOR2X1_LOC_210/B INVX1_LOC_117/A 0.03fF
C30127 INVX1_LOC_189/Y INVX1_LOC_38/A 0.01fF
C30128 INVX1_LOC_40/A NOR2X1_LOC_98/B 0.07fF
C30129 INVX1_LOC_89/A INVX1_LOC_95/Y 0.08fF
C30130 INVX1_LOC_122/Y NOR2X1_LOC_509/A 0.03fF
C30131 NAND2X1_LOC_214/B NOR2X1_LOC_646/B 0.08fF
C30132 NOR2X1_LOC_220/A INVX1_LOC_38/A 0.03fF
C30133 NAND2X1_LOC_65/a_36_24# NOR2X1_LOC_849/A 0.00fF
C30134 INVX1_LOC_31/A NOR2X1_LOC_643/a_36_216# 0.01fF
C30135 INVX1_LOC_184/Y NOR2X1_LOC_814/A 0.05fF
C30136 INVX1_LOC_23/A NOR2X1_LOC_663/A 0.01fF
C30137 INVX1_LOC_227/A VDD 0.05fF
C30138 NOR2X1_LOC_91/A NOR2X1_LOC_384/A 0.00fF
C30139 NOR2X1_LOC_123/B INVX1_LOC_76/A 0.10fF
C30140 NOR2X1_LOC_763/Y VDD 0.12fF
C30141 NOR2X1_LOC_360/Y NAND2X1_LOC_74/B 0.07fF
C30142 INVX1_LOC_104/A NOR2X1_LOC_197/B 0.10fF
C30143 NOR2X1_LOC_188/A INVX1_LOC_48/A 0.03fF
C30144 NOR2X1_LOC_717/B INVX1_LOC_14/Y 0.01fF
C30145 INVX1_LOC_233/A NOR2X1_LOC_109/Y 0.00fF
C30146 NOR2X1_LOC_356/A NOR2X1_LOC_324/B 0.23fF
C30147 NAND2X1_LOC_850/Y INVX1_LOC_185/A 0.01fF
C30148 INVX1_LOC_8/A NOR2X1_LOC_179/Y 0.06fF
C30149 NOR2X1_LOC_589/A NOR2X1_LOC_536/A 0.03fF
C30150 INVX1_LOC_301/Y INVX1_LOC_301/A 0.01fF
C30151 NOR2X1_LOC_644/A NOR2X1_LOC_35/Y 0.03fF
C30152 NAND2X1_LOC_721/A NAND2X1_LOC_808/A 0.02fF
C30153 NOR2X1_LOC_548/Y INVX1_LOC_38/A 0.07fF
C30154 INVX1_LOC_135/A INVX1_LOC_194/Y 0.01fF
C30155 NAND2X1_LOC_198/B NAND2X1_LOC_807/B 0.01fF
C30156 NOR2X1_LOC_219/Y INVX1_LOC_54/A 0.04fF
C30157 D_INPUT_0 INVX1_LOC_12/Y 0.03fF
C30158 INVX1_LOC_72/Y INVX1_LOC_42/A 0.02fF
C30159 INVX1_LOC_225/Y INVX1_LOC_78/A 0.07fF
C30160 INVX1_LOC_174/A NAND2X1_LOC_470/B 0.05fF
C30161 INVX1_LOC_1/A NOR2X1_LOC_383/B 0.35fF
C30162 INVX1_LOC_229/Y NOR2X1_LOC_536/A 0.10fF
C30163 INVX1_LOC_90/A NOR2X1_LOC_447/B 0.03fF
C30164 NOR2X1_LOC_561/Y NOR2X1_LOC_331/B 0.17fF
C30165 INVX1_LOC_41/A NAND2X1_LOC_773/B 0.02fF
C30166 INVX1_LOC_246/Y INVX1_LOC_42/A 0.00fF
C30167 NAND2X1_LOC_795/Y INVX1_LOC_38/A 0.01fF
C30168 INVX1_LOC_16/A NAND2X1_LOC_243/Y 0.10fF
C30169 INVX1_LOC_102/Y INVX1_LOC_76/A 0.10fF
C30170 INVX1_LOC_205/A INVX1_LOC_15/A 0.00fF
C30171 INVX1_LOC_83/A NOR2X1_LOC_865/A 0.05fF
C30172 INVX1_LOC_16/A INVX1_LOC_89/Y 0.01fF
C30173 NOR2X1_LOC_784/Y NOR2X1_LOC_383/B 0.04fF
C30174 INVX1_LOC_50/A INVX1_LOC_73/Y 0.02fF
C30175 VDD NOR2X1_LOC_703/A 0.00fF
C30176 NOR2X1_LOC_598/B NAND2X1_LOC_218/A 0.00fF
C30177 INVX1_LOC_1/Y INVX1_LOC_92/A 0.10fF
C30178 NAND2X1_LOC_462/B NOR2X1_LOC_629/Y 0.00fF
C30179 INVX1_LOC_177/A NOR2X1_LOC_814/A 0.03fF
C30180 NAND2X1_LOC_802/A INVX1_LOC_42/A 0.00fF
C30181 INVX1_LOC_182/A INVX1_LOC_37/A 0.12fF
C30182 INVX1_LOC_135/A INVX1_LOC_9/A 0.03fF
C30183 NAND2X1_LOC_352/B NAND2X1_LOC_286/B 0.01fF
C30184 NAND2X1_LOC_703/Y NOR2X1_LOC_109/Y 0.36fF
C30185 NOR2X1_LOC_794/B NOR2X1_LOC_383/B 0.02fF
C30186 NOR2X1_LOC_151/Y INVX1_LOC_14/Y 0.03fF
C30187 NOR2X1_LOC_398/Y NAND2X1_LOC_773/B 0.03fF
C30188 NOR2X1_LOC_516/B NOR2X1_LOC_243/B 0.10fF
C30189 INVX1_LOC_314/Y INVX1_LOC_32/A 0.07fF
C30190 NOR2X1_LOC_78/B INVX1_LOC_63/A 0.34fF
C30191 INVX1_LOC_265/A INVX1_LOC_102/A 0.02fF
C30192 NOR2X1_LOC_561/Y NOR2X1_LOC_592/B 0.05fF
C30193 NAND2X1_LOC_123/Y INVX1_LOC_66/Y 0.05fF
C30194 NOR2X1_LOC_6/B NOR2X1_LOC_67/a_36_216# 0.00fF
C30195 NOR2X1_LOC_225/a_36_216# INVX1_LOC_29/Y 0.00fF
C30196 INVX1_LOC_62/Y NAND2X1_LOC_223/A 0.07fF
C30197 INVX1_LOC_171/A NAND2X1_LOC_93/B 0.03fF
C30198 NAND2X1_LOC_738/B NOR2X1_LOC_766/a_36_216# 0.00fF
C30199 INVX1_LOC_246/Y INVX1_LOC_78/A 0.00fF
C30200 NOR2X1_LOC_773/Y INVX1_LOC_19/A 0.07fF
C30201 NOR2X1_LOC_91/A INVX1_LOC_72/A 0.13fF
C30202 NAND2X1_LOC_859/Y INVX1_LOC_119/Y 0.31fF
C30203 NOR2X1_LOC_791/Y NOR2X1_LOC_271/B 0.02fF
C30204 NOR2X1_LOC_178/Y NOR2X1_LOC_103/Y 0.02fF
C30205 NOR2X1_LOC_160/B NOR2X1_LOC_342/A 0.17fF
C30206 NAND2X1_LOC_573/A INVX1_LOC_285/A 0.10fF
C30207 INVX1_LOC_35/A INVX1_LOC_230/Y 0.07fF
C30208 NAND2X1_LOC_802/A INVX1_LOC_78/A 0.06fF
C30209 INVX1_LOC_28/A NAND2X1_LOC_243/Y 0.01fF
C30210 NOR2X1_LOC_667/A NOR2X1_LOC_89/A 0.12fF
C30211 INVX1_LOC_2/Y NOR2X1_LOC_78/A 0.01fF
C30212 INVX1_LOC_21/A INVX1_LOC_224/A 0.05fF
C30213 NOR2X1_LOC_317/B NOR2X1_LOC_855/A 0.10fF
C30214 INVX1_LOC_72/A INVX1_LOC_23/A 5.44fF
C30215 INVX1_LOC_50/A NOR2X1_LOC_91/Y 0.09fF
C30216 INVX1_LOC_278/Y NOR2X1_LOC_519/Y 0.02fF
C30217 INVX1_LOC_77/A NOR2X1_LOC_541/B 0.20fF
C30218 NOR2X1_LOC_510/Y NAND2X1_LOC_803/B 0.02fF
C30219 INVX1_LOC_21/A INVX1_LOC_11/A 1.20fF
C30220 NAND2X1_LOC_9/Y INVX1_LOC_36/A 0.04fF
C30221 D_INPUT_1 INVX1_LOC_18/A 0.14fF
C30222 NOR2X1_LOC_310/Y INVX1_LOC_4/A 0.04fF
C30223 INVX1_LOC_83/A INVX1_LOC_63/A 0.41fF
C30224 INVX1_LOC_233/A INVX1_LOC_36/A 0.08fF
C30225 INVX1_LOC_178/A INVX1_LOC_161/Y 0.05fF
C30226 NOR2X1_LOC_742/A INVX1_LOC_92/A 0.09fF
C30227 INVX1_LOC_53/Y NAND2X1_LOC_807/B 0.01fF
C30228 INVX1_LOC_286/A NOR2X1_LOC_652/a_36_216# 0.01fF
C30229 NOR2X1_LOC_78/A NOR2X1_LOC_363/Y 0.01fF
C30230 NAND2X1_LOC_729/Y NAND2X1_LOC_738/B 0.01fF
C30231 INVX1_LOC_108/Y INVX1_LOC_205/A 0.05fF
C30232 INVX1_LOC_198/Y INVX1_LOC_23/A 0.01fF
C30233 NOR2X1_LOC_553/B INVX1_LOC_29/A 0.01fF
C30234 NOR2X1_LOC_113/B INVX1_LOC_54/A 0.04fF
C30235 NOR2X1_LOC_309/Y NOR2X1_LOC_282/a_36_216# 0.01fF
C30236 INVX1_LOC_30/Y NOR2X1_LOC_327/a_36_216# 0.00fF
C30237 NOR2X1_LOC_510/Y NOR2X1_LOC_590/A 0.03fF
C30238 NOR2X1_LOC_453/Y INVX1_LOC_11/A 0.01fF
C30239 NOR2X1_LOC_332/A INVX1_LOC_19/A 0.19fF
C30240 NOR2X1_LOC_405/A INVX1_LOC_33/Y 0.02fF
C30241 INVX1_LOC_49/A NAND2X1_LOC_64/a_36_24# 0.02fF
C30242 INVX1_LOC_141/Y NOR2X1_LOC_406/A 0.03fF
C30243 NAND2X1_LOC_859/Y INVX1_LOC_284/A 0.62fF
C30244 INPUT_0 NAND2X1_LOC_802/Y 0.14fF
C30245 INVX1_LOC_266/Y INVX1_LOC_78/A 0.02fF
C30246 INVX1_LOC_118/Y INVX1_LOC_91/A 0.04fF
C30247 NAND2X1_LOC_650/B VDD 0.48fF
C30248 INVX1_LOC_136/A NOR2X1_LOC_212/a_36_216# 0.01fF
C30249 NAND2X1_LOC_53/Y INVX1_LOC_103/A 0.10fF
C30250 INVX1_LOC_276/A INVX1_LOC_273/A 0.42fF
C30251 INVX1_LOC_14/A NAND2X1_LOC_807/A 0.01fF
C30252 INVX1_LOC_40/A NOR2X1_LOC_38/B 0.03fF
C30253 NAND2X1_LOC_326/A NOR2X1_LOC_595/a_36_216# 0.00fF
C30254 INVX1_LOC_228/Y NOR2X1_LOC_82/A 0.01fF
C30255 NOR2X1_LOC_859/A NOR2X1_LOC_849/A 0.14fF
C30256 NOR2X1_LOC_552/A INVX1_LOC_9/A 0.07fF
C30257 NOR2X1_LOC_205/a_36_216# NOR2X1_LOC_334/Y 0.01fF
C30258 NAND2X1_LOC_357/B NAND2X1_LOC_286/B 0.00fF
C30259 INVX1_LOC_18/A NOR2X1_LOC_652/Y 0.07fF
C30260 NOR2X1_LOC_136/Y NOR2X1_LOC_334/Y 0.02fF
C30261 INVX1_LOC_12/Y NOR2X1_LOC_266/B 0.05fF
C30262 NOR2X1_LOC_78/A INVX1_LOC_307/Y 0.01fF
C30263 NOR2X1_LOC_617/Y NAND2X1_LOC_624/B 0.06fF
C30264 INVX1_LOC_38/A NAND2X1_LOC_655/B 0.01fF
C30265 INVX1_LOC_10/A NOR2X1_LOC_116/a_36_216# 0.00fF
C30266 NOR2X1_LOC_590/A NOR2X1_LOC_361/B 0.06fF
C30267 NOR2X1_LOC_78/A NOR2X1_LOC_358/a_36_216# 0.00fF
C30268 NOR2X1_LOC_234/Y NAND2X1_LOC_464/B -0.03fF
C30269 INVX1_LOC_38/A NAND2X1_LOC_469/B 0.03fF
C30270 NOR2X1_LOC_536/A INVX1_LOC_20/A 0.49fF
C30271 NOR2X1_LOC_482/Y NOR2X1_LOC_693/Y 0.25fF
C30272 INVX1_LOC_135/A NOR2X1_LOC_861/Y 0.86fF
C30273 NOR2X1_LOC_318/B INVX1_LOC_92/A 0.07fF
C30274 INVX1_LOC_30/A INVX1_LOC_198/A 0.00fF
C30275 NOR2X1_LOC_816/A INVX1_LOC_161/Y 0.05fF
C30276 NOR2X1_LOC_91/A NAND2X1_LOC_338/B 0.07fF
C30277 INVX1_LOC_7/Y INVX1_LOC_24/A 0.02fF
C30278 INVX1_LOC_277/Y INVX1_LOC_1/A 0.03fF
C30279 NOR2X1_LOC_331/B INVX1_LOC_76/A 0.08fF
C30280 INVX1_LOC_140/A NOR2X1_LOC_11/Y 0.03fF
C30281 NOR2X1_LOC_686/B INVX1_LOC_15/A 0.01fF
C30282 INVX1_LOC_124/Y NOR2X1_LOC_401/A 0.02fF
C30283 INVX1_LOC_6/A INVX1_LOC_119/Y 0.13fF
C30284 NOR2X1_LOC_193/a_36_216# INVX1_LOC_63/A 0.01fF
C30285 NOR2X1_LOC_78/B NOR2X1_LOC_65/Y 0.00fF
C30286 INVX1_LOC_93/Y INVX1_LOC_92/A 0.07fF
C30287 INVX1_LOC_285/Y NOR2X1_LOC_814/A 0.01fF
C30288 NOR2X1_LOC_589/A NAND2X1_LOC_470/B 0.03fF
C30289 NOR2X1_LOC_560/A NOR2X1_LOC_861/Y 0.01fF
C30290 INVX1_LOC_233/A NOR2X1_LOC_309/Y 0.10fF
C30291 NOR2X1_LOC_655/Y INVX1_LOC_20/A 0.01fF
C30292 INVX1_LOC_16/A INVX1_LOC_16/Y 0.33fF
C30293 INVX1_LOC_22/A NOR2X1_LOC_318/A 2.96fF
C30294 NAND2X1_LOC_337/B INVX1_LOC_312/A -0.01fF
C30295 INVX1_LOC_21/A NOR2X1_LOC_433/A 0.12fF
C30296 NOR2X1_LOC_92/Y INVX1_LOC_24/A 0.89fF
C30297 NAND2X1_LOC_338/B INVX1_LOC_23/A 0.29fF
C30298 INVX1_LOC_150/Y INVX1_LOC_30/A 0.29fF
C30299 NAND2X1_LOC_93/B INVX1_LOC_20/A 0.08fF
C30300 INVX1_LOC_83/A NAND2X1_LOC_452/Y 0.03fF
C30301 NOR2X1_LOC_666/A NOR2X1_LOC_759/Y 0.28fF
C30302 INVX1_LOC_24/Y INVX1_LOC_24/A 0.02fF
C30303 NOR2X1_LOC_561/Y NOR2X1_LOC_449/A 0.11fF
C30304 NAND2X1_LOC_323/B INVX1_LOC_23/A 0.00fF
C30305 NAND2X1_LOC_778/Y NAND2X1_LOC_325/Y 0.01fF
C30306 INVX1_LOC_21/A NOR2X1_LOC_593/Y 0.10fF
C30307 NOR2X1_LOC_667/A NAND2X1_LOC_804/A 0.02fF
C30308 NAND2X1_LOC_713/a_36_24# INVX1_LOC_24/A 0.01fF
C30309 NAND2X1_LOC_21/Y D_INPUT_6 0.37fF
C30310 INVX1_LOC_139/A INVX1_LOC_92/A 0.06fF
C30311 INVX1_LOC_42/Y INVX1_LOC_42/A 0.01fF
C30312 INVX1_LOC_148/A INVX1_LOC_15/A 0.03fF
C30313 NOR2X1_LOC_491/Y INVX1_LOC_76/A 0.11fF
C30314 INVX1_LOC_83/A NOR2X1_LOC_307/Y 0.03fF
C30315 INVX1_LOC_77/Y INVX1_LOC_54/A 0.04fF
C30316 INVX1_LOC_311/A NOR2X1_LOC_89/A 0.08fF
C30317 INVX1_LOC_89/A INVX1_LOC_271/Y 0.09fF
C30318 INVX1_LOC_91/A NOR2X1_LOC_258/Y 0.01fF
C30319 INVX1_LOC_16/A NAND2X1_LOC_205/A 0.03fF
C30320 INVX1_LOC_65/A NOR2X1_LOC_814/A 0.00fF
C30321 NOR2X1_LOC_798/A NOR2X1_LOC_309/Y 1.47fF
C30322 NOR2X1_LOC_15/Y NOR2X1_LOC_753/Y 0.03fF
C30323 INVX1_LOC_280/A INVX1_LOC_9/A 0.10fF
C30324 NAND2X1_LOC_721/A INVX1_LOC_92/A 0.03fF
C30325 NOR2X1_LOC_163/Y NOR2X1_LOC_467/A 0.30fF
C30326 INVX1_LOC_269/A INVX1_LOC_49/A 0.07fF
C30327 NAND2X1_LOC_741/B NOR2X1_LOC_761/Y 0.06fF
C30328 NOR2X1_LOC_468/Y INVX1_LOC_33/A 2.28fF
C30329 INVX1_LOC_21/A NOR2X1_LOC_52/B 19.48fF
C30330 INVX1_LOC_250/A INVX1_LOC_141/Y 0.01fF
C30331 INVX1_LOC_279/A NOR2X1_LOC_748/A 0.10fF
C30332 INVX1_LOC_1/Y INVX1_LOC_53/A 0.03fF
C30333 NAND2X1_LOC_374/Y NOR2X1_LOC_291/a_36_216# 0.00fF
C30334 INVX1_LOC_20/A NOR2X1_LOC_649/B 0.02fF
C30335 NAND2X1_LOC_190/Y INVX1_LOC_33/A 0.03fF
C30336 NAND2X1_LOC_703/Y NOR2X1_LOC_309/Y 0.02fF
C30337 INVX1_LOC_70/Y NAND2X1_LOC_81/B 0.91fF
C30338 INVX1_LOC_20/A INVX1_LOC_3/A 0.10fF
C30339 NOR2X1_LOC_340/a_36_216# NOR2X1_LOC_340/A 0.02fF
C30340 INVX1_LOC_22/A NOR2X1_LOC_678/A 0.03fF
C30341 INVX1_LOC_22/A INVX1_LOC_295/Y 0.01fF
C30342 NOR2X1_LOC_441/Y NAND2X1_LOC_198/B 0.03fF
C30343 NAND2X1_LOC_802/A NOR2X1_LOC_503/Y 0.02fF
C30344 NOR2X1_LOC_76/A INVX1_LOC_181/A 0.00fF
C30345 INVX1_LOC_125/Y INVX1_LOC_42/A 0.07fF
C30346 INVX1_LOC_73/A INVX1_LOC_94/Y 0.03fF
C30347 NOR2X1_LOC_590/A INVX1_LOC_184/Y 0.02fF
C30348 NAND2X1_LOC_563/Y NOR2X1_LOC_381/Y 0.04fF
C30349 INVX1_LOC_46/A INVX1_LOC_63/A 13.30fF
C30350 INVX1_LOC_136/A NOR2X1_LOC_360/Y 0.07fF
C30351 INVX1_LOC_304/A NOR2X1_LOC_89/A 0.08fF
C30352 NOR2X1_LOC_393/a_36_216# INVX1_LOC_23/Y 0.01fF
C30353 NAND2X1_LOC_842/B INVX1_LOC_270/A 0.02fF
C30354 INVX1_LOC_13/A NAND2X1_LOC_214/B 0.07fF
C30355 INVX1_LOC_45/A NOR2X1_LOC_274/Y 0.01fF
C30356 INVX1_LOC_12/A INVX1_LOC_59/Y 0.03fF
C30357 NOR2X1_LOC_389/A INVX1_LOC_33/A 0.10fF
C30358 INVX1_LOC_2/A INVX1_LOC_269/A 0.07fF
C30359 INVX1_LOC_313/Y INVX1_LOC_23/A 0.15fF
C30360 INVX1_LOC_24/Y INVX1_LOC_143/A 0.10fF
C30361 NOR2X1_LOC_557/A INVX1_LOC_32/A 0.07fF
C30362 NOR2X1_LOC_78/a_36_216# NOR2X1_LOC_78/Y 0.01fF
C30363 NOR2X1_LOC_160/B NOR2X1_LOC_121/Y 0.05fF
C30364 NOR2X1_LOC_272/Y INVX1_LOC_232/A 0.01fF
C30365 NOR2X1_LOC_389/A NOR2X1_LOC_743/a_36_216# 0.00fF
C30366 NOR2X1_LOC_274/Y NOR2X1_LOC_568/A 0.47fF
C30367 NOR2X1_LOC_75/Y NOR2X1_LOC_194/Y 0.01fF
C30368 NOR2X1_LOC_67/A NOR2X1_LOC_15/Y 0.08fF
C30369 INVX1_LOC_2/A NOR2X1_LOC_232/Y 0.20fF
C30370 INVX1_LOC_14/A NAND2X1_LOC_360/B 0.16fF
C30371 INVX1_LOC_117/A NOR2X1_LOC_257/Y 0.02fF
C30372 INVX1_LOC_191/A INVX1_LOC_78/A 0.14fF
C30373 NAND2X1_LOC_387/B INVX1_LOC_77/A 0.03fF
C30374 NOR2X1_LOC_226/A INVX1_LOC_269/A 0.70fF
C30375 NOR2X1_LOC_250/A NAND2X1_LOC_660/A 0.01fF
C30376 INVX1_LOC_13/A INVX1_LOC_27/A 0.28fF
C30377 NAND2X1_LOC_239/a_36_24# NAND2X1_LOC_350/A 0.01fF
C30378 NOR2X1_LOC_384/Y NAND2X1_LOC_632/B 0.01fF
C30379 NOR2X1_LOC_643/Y NOR2X1_LOC_554/B 0.03fF
C30380 NAND2X1_LOC_354/Y NOR2X1_LOC_433/A 0.01fF
C30381 NOR2X1_LOC_689/Y NAND2X1_LOC_863/A 0.03fF
C30382 NOR2X1_LOC_636/B NAND2X1_LOC_11/Y 0.15fF
C30383 INVX1_LOC_39/A NOR2X1_LOC_391/A 0.04fF
C30384 INVX1_LOC_35/A INVX1_LOC_196/Y 0.03fF
C30385 NOR2X1_LOC_20/Y NOR2X1_LOC_399/Y 0.15fF
C30386 NOR2X1_LOC_658/Y NOR2X1_LOC_364/Y -0.02fF
C30387 INVX1_LOC_24/A NAND2X1_LOC_837/Y 0.07fF
C30388 INVX1_LOC_11/A NOR2X1_LOC_667/A 0.25fF
C30389 INVX1_LOC_166/A NAND2X1_LOC_463/B 0.01fF
C30390 VDD NOR2X1_LOC_67/Y 0.18fF
C30391 NOR2X1_LOC_636/A NOR2X1_LOC_68/A 0.01fF
C30392 INVX1_LOC_11/A INVX1_LOC_248/A 0.43fF
C30393 NOR2X1_LOC_158/a_36_216# INVX1_LOC_91/A 0.00fF
C30394 NOR2X1_LOC_88/Y NAND2X1_LOC_798/B 0.47fF
C30395 NAND2X1_LOC_623/a_36_24# NAND2X1_LOC_866/B 0.02fF
C30396 INVX1_LOC_6/A NOR2X1_LOC_134/a_36_216# 0.00fF
C30397 NOR2X1_LOC_272/Y NOR2X1_LOC_366/Y 0.03fF
C30398 NOR2X1_LOC_590/A INVX1_LOC_177/A 0.03fF
C30399 NOR2X1_LOC_188/A NOR2X1_LOC_383/B 0.00fF
C30400 INVX1_LOC_140/Y INVX1_LOC_173/A 0.04fF
C30401 NOR2X1_LOC_214/a_36_216# NOR2X1_LOC_759/Y 0.00fF
C30402 INVX1_LOC_107/Y INVX1_LOC_113/A 0.00fF
C30403 INVX1_LOC_256/A NOR2X1_LOC_131/Y 0.03fF
C30404 INVX1_LOC_31/A NOR2X1_LOC_537/Y 0.12fF
C30405 INVX1_LOC_136/A NOR2X1_LOC_792/B 0.00fF
C30406 INVX1_LOC_254/A NOR2X1_LOC_419/Y 0.00fF
C30407 NAND2X1_LOC_338/B INVX1_LOC_31/A 0.07fF
C30408 NOR2X1_LOC_716/a_36_216# NAND2X1_LOC_793/B 0.02fF
C30409 NOR2X1_LOC_837/Y NAND2X1_LOC_364/Y 0.03fF
C30410 INVX1_LOC_33/A NOR2X1_LOC_596/A 0.03fF
C30411 INVX1_LOC_41/A INVX1_LOC_24/A 0.03fF
C30412 NOR2X1_LOC_65/B INVX1_LOC_125/Y 0.10fF
C30413 NOR2X1_LOC_48/B INVX1_LOC_77/Y 0.10fF
C30414 GATE_579 INVX1_LOC_22/A 0.03fF
C30415 INVX1_LOC_269/A NAND2X1_LOC_462/B 0.01fF
C30416 NOR2X1_LOC_92/Y NAND2X1_LOC_800/Y 0.01fF
C30417 NOR2X1_LOC_498/Y INVX1_LOC_24/A 0.09fF
C30418 INVX1_LOC_292/A NOR2X1_LOC_500/Y 1.20fF
C30419 NOR2X1_LOC_92/Y NOR2X1_LOC_130/A 0.10fF
C30420 INVX1_LOC_78/Y NOR2X1_LOC_858/A 0.65fF
C30421 NOR2X1_LOC_793/A D_INPUT_0 0.03fF
C30422 INVX1_LOC_27/A INVX1_LOC_55/Y 0.30fF
C30423 INVX1_LOC_256/A NOR2X1_LOC_589/A 0.22fF
C30424 INVX1_LOC_103/A INVX1_LOC_10/A 0.26fF
C30425 INVX1_LOC_55/A INVX1_LOC_22/A 0.04fF
C30426 NOR2X1_LOC_604/Y INVX1_LOC_6/A 0.01fF
C30427 INVX1_LOC_191/Y INVX1_LOC_72/A 0.03fF
C30428 INVX1_LOC_88/A NOR2X1_LOC_60/a_36_216# 0.00fF
C30429 NAND2X1_LOC_483/Y NOR2X1_LOC_495/Y 0.87fF
C30430 NAND2X1_LOC_773/Y INVX1_LOC_89/A 0.01fF
C30431 NOR2X1_LOC_33/A NOR2X1_LOC_160/B 0.01fF
C30432 NOR2X1_LOC_619/A INVX1_LOC_218/Y 0.22fF
C30433 NOR2X1_LOC_191/B INVX1_LOC_104/A 0.05fF
C30434 INVX1_LOC_280/A NOR2X1_LOC_861/Y 0.02fF
C30435 NAND2X1_LOC_435/a_36_24# INVX1_LOC_186/Y 0.01fF
C30436 NAND2X1_LOC_811/Y NOR2X1_LOC_152/Y 0.06fF
C30437 INVX1_LOC_24/A NAND2X1_LOC_477/A 0.03fF
C30438 NAND2X1_LOC_764/a_36_24# NAND2X1_LOC_451/Y 0.00fF
C30439 INVX1_LOC_98/A INVX1_LOC_29/Y 0.00fF
C30440 NAND2X1_LOC_374/Y NAND2X1_LOC_634/Y 0.18fF
C30441 INVX1_LOC_47/Y NOR2X1_LOC_440/a_36_216# 0.01fF
C30442 INVX1_LOC_41/A NOR2X1_LOC_557/Y 0.10fF
C30443 NOR2X1_LOC_449/A INVX1_LOC_76/A 0.03fF
C30444 INVX1_LOC_269/A INPUT_1 0.21fF
C30445 INVX1_LOC_292/A INVX1_LOC_10/A 0.03fF
C30446 VDD NOR2X1_LOC_415/Y 0.35fF
C30447 D_INPUT_0 NAND2X1_LOC_550/A 0.07fF
C30448 NOR2X1_LOC_318/B INVX1_LOC_53/A 0.04fF
C30449 NOR2X1_LOC_795/Y INVX1_LOC_77/A 0.05fF
C30450 INVX1_LOC_278/Y INVX1_LOC_217/A 0.03fF
C30451 NAND2X1_LOC_276/Y INVX1_LOC_8/A 0.07fF
C30452 NOR2X1_LOC_590/A NAND2X1_LOC_573/A 0.00fF
C30453 NOR2X1_LOC_669/A INVX1_LOC_92/A 0.02fF
C30454 NOR2X1_LOC_536/A INVX1_LOC_4/A 0.48fF
C30455 NOR2X1_LOC_403/B INVX1_LOC_34/Y 0.05fF
C30456 NOR2X1_LOC_152/Y INVX1_LOC_266/Y 0.30fF
C30457 INVX1_LOC_256/A INVX1_LOC_171/A 0.01fF
C30458 NOR2X1_LOC_590/A NOR2X1_LOC_785/Y 0.04fF
C30459 D_INPUT_0 NOR2X1_LOC_160/B 10.43fF
C30460 INVX1_LOC_286/Y NAND2X1_LOC_854/B 0.05fF
C30461 INVX1_LOC_113/Y INVX1_LOC_266/Y 0.23fF
C30462 NOR2X1_LOC_764/Y INVX1_LOC_174/A 0.03fF
C30463 INVX1_LOC_284/Y NOR2X1_LOC_298/Y 0.40fF
C30464 D_GATE_741 INVX1_LOC_85/Y 0.00fF
C30465 NAND2X1_LOC_364/A INVX1_LOC_232/A 0.11fF
C30466 INVX1_LOC_305/A INVX1_LOC_22/A 0.01fF
C30467 NAND2X1_LOC_833/Y NOR2X1_LOC_315/Y 0.08fF
C30468 INVX1_LOC_62/Y INVX1_LOC_40/A 0.01fF
C30469 INVX1_LOC_76/Y NOR2X1_LOC_379/a_36_216# 0.00fF
C30470 INVX1_LOC_1/A NOR2X1_LOC_163/Y 0.09fF
C30471 INVX1_LOC_46/A NOR2X1_LOC_65/Y 0.00fF
C30472 NAND2X1_LOC_81/B INVX1_LOC_285/A 0.09fF
C30473 INVX1_LOC_214/A NOR2X1_LOC_433/A 0.12fF
C30474 NAND2X1_LOC_563/Y NOR2X1_LOC_6/B 0.06fF
C30475 NOR2X1_LOC_294/a_36_216# NOR2X1_LOC_332/A 0.01fF
C30476 NOR2X1_LOC_222/Y NOR2X1_LOC_219/a_36_216# 0.00fF
C30477 NOR2X1_LOC_655/Y INVX1_LOC_4/A 0.01fF
C30478 INVX1_LOC_280/A NOR2X1_LOC_825/a_36_216# 0.00fF
C30479 NOR2X1_LOC_808/A NOR2X1_LOC_551/B 0.01fF
C30480 INVX1_LOC_41/A INVX1_LOC_143/A 0.41fF
C30481 NOR2X1_LOC_614/Y INVX1_LOC_77/A 0.47fF
C30482 INVX1_LOC_161/Y INVX1_LOC_140/A 0.03fF
C30483 NOR2X1_LOC_128/A INVX1_LOC_3/A 0.03fF
C30484 NAND2X1_LOC_798/B INVX1_LOC_15/A 0.23fF
C30485 NAND2X1_LOC_93/B INVX1_LOC_4/A 3.04fF
C30486 INVX1_LOC_94/A NOR2X1_LOC_569/Y 0.00fF
C30487 NOR2X1_LOC_220/A INVX1_LOC_33/A 0.03fF
C30488 INVX1_LOC_78/Y NOR2X1_LOC_698/a_36_216# 0.00fF
C30489 INVX1_LOC_196/A INVX1_LOC_176/Y 0.25fF
C30490 INVX1_LOC_11/A NAND2X1_LOC_51/B 0.08fF
C30491 NAND2X1_LOC_325/Y NAND2X1_LOC_840/B 0.00fF
C30492 NOR2X1_LOC_541/B INVX1_LOC_9/A 0.05fF
C30493 NOR2X1_LOC_778/B NOR2X1_LOC_337/a_36_216# 0.02fF
C30494 INVX1_LOC_214/A NOR2X1_LOC_52/B 0.03fF
C30495 INVX1_LOC_72/A NAND2X1_LOC_866/B 0.07fF
C30496 NAND2X1_LOC_99/Y INVX1_LOC_13/A 0.02fF
C30497 INVX1_LOC_36/A NAND2X1_LOC_842/B 1.35fF
C30498 NOR2X1_LOC_219/Y NOR2X1_LOC_142/Y 0.22fF
C30499 INVX1_LOC_11/A INVX1_LOC_311/A 1.05fF
C30500 NOR2X1_LOC_454/Y NOR2X1_LOC_45/B 0.13fF
C30501 NOR2X1_LOC_667/A NOR2X1_LOC_52/B 0.07fF
C30502 NAND2X1_LOC_721/A INVX1_LOC_53/A 0.42fF
C30503 INVX1_LOC_24/A NOR2X1_LOC_299/Y 0.13fF
C30504 NOR2X1_LOC_382/a_36_216# NOR2X1_LOC_84/A 0.00fF
C30505 NOR2X1_LOC_155/A NOR2X1_LOC_334/Y 0.07fF
C30506 INVX1_LOC_248/A NOR2X1_LOC_52/B 0.07fF
C30507 INVX1_LOC_87/A INVX1_LOC_92/A 0.13fF
C30508 INVX1_LOC_256/A INVX1_LOC_222/A 0.03fF
C30509 NOR2X1_LOC_290/Y NAND2X1_LOC_338/B 0.02fF
C30510 INVX1_LOC_33/A NOR2X1_LOC_548/Y 0.01fF
C30511 NAND2X1_LOC_657/a_36_24# INVX1_LOC_32/A 0.00fF
C30512 INVX1_LOC_36/A INVX1_LOC_146/A 0.01fF
C30513 NOR2X1_LOC_471/Y NOR2X1_LOC_589/Y 0.04fF
C30514 NOR2X1_LOC_267/A NAND2X1_LOC_842/B 0.05fF
C30515 INVX1_LOC_19/A INVX1_LOC_42/A 2.05fF
C30516 INVX1_LOC_47/Y INVX1_LOC_84/A 0.07fF
C30517 NAND2X1_LOC_367/A INVX1_LOC_160/Y 0.01fF
C30518 NOR2X1_LOC_649/B INVX1_LOC_4/A 0.04fF
C30519 NOR2X1_LOC_632/Y INVX1_LOC_34/A 2.05fF
C30520 INVX1_LOC_3/A INVX1_LOC_4/A 0.04fF
C30521 NOR2X1_LOC_142/Y NOR2X1_LOC_665/A 0.10fF
C30522 INVX1_LOC_67/A INVX1_LOC_10/A 0.03fF
C30523 NOR2X1_LOC_454/Y INVX1_LOC_199/Y 0.10fF
C30524 NAND2X1_LOC_865/a_36_24# INVX1_LOC_41/Y 0.00fF
C30525 INVX1_LOC_276/A NAND2X1_LOC_840/B 0.03fF
C30526 NOR2X1_LOC_196/A NOR2X1_LOC_112/Y 0.07fF
C30527 INVX1_LOC_41/A NOR2X1_LOC_739/a_36_216# 0.00fF
C30528 NOR2X1_LOC_590/A INVX1_LOC_285/Y 0.19fF
C30529 NOR2X1_LOC_267/a_36_216# INVX1_LOC_93/Y 0.00fF
C30530 INVX1_LOC_27/A NOR2X1_LOC_357/Y 0.07fF
C30531 NOR2X1_LOC_238/a_36_216# INVX1_LOC_28/A 0.01fF
C30532 INVX1_LOC_4/Y NOR2X1_LOC_814/A 0.10fF
C30533 NOR2X1_LOC_626/a_36_216# INVX1_LOC_139/Y 0.00fF
C30534 INVX1_LOC_64/A NOR2X1_LOC_536/A 0.07fF
C30535 NOR2X1_LOC_521/Y NOR2X1_LOC_52/B 0.05fF
C30536 INVX1_LOC_249/A INVX1_LOC_55/Y 0.03fF
C30537 INVX1_LOC_41/A NOR2X1_LOC_130/A 0.03fF
C30538 NAND2X1_LOC_190/Y NOR2X1_LOC_486/Y 0.01fF
C30539 INVX1_LOC_78/A NOR2X1_LOC_653/Y 0.12fF
C30540 NAND2X1_LOC_361/Y INVX1_LOC_132/Y 0.03fF
C30541 INVX1_LOC_240/A INVX1_LOC_10/A 0.02fF
C30542 INVX1_LOC_255/Y INVX1_LOC_216/A -0.01fF
C30543 NAND2X1_LOC_796/B NOR2X1_LOC_111/A 0.06fF
C30544 NOR2X1_LOC_15/Y NAND2X1_LOC_855/a_36_24# 0.00fF
C30545 NOR2X1_LOC_78/B INVX1_LOC_1/Y 0.01fF
C30546 NOR2X1_LOC_89/A INVX1_LOC_19/Y 0.01fF
C30547 NOR2X1_LOC_276/Y NOR2X1_LOC_269/Y 0.37fF
C30548 INVX1_LOC_172/A NOR2X1_LOC_497/Y 0.03fF
C30549 INVX1_LOC_35/A NOR2X1_LOC_641/Y 0.02fF
C30550 INVX1_LOC_90/A INVX1_LOC_63/Y 0.04fF
C30551 INVX1_LOC_227/A INVX1_LOC_177/A 0.03fF
C30552 INVX1_LOC_72/A INVX1_LOC_6/A 0.44fF
C30553 INVX1_LOC_308/A NOR2X1_LOC_743/Y 0.01fF
C30554 INVX1_LOC_53/A INVX1_LOC_117/Y 0.03fF
C30555 NAND2X1_LOC_477/A NOR2X1_LOC_130/A 0.45fF
C30556 INVX1_LOC_78/A INVX1_LOC_19/A 0.18fF
C30557 NOR2X1_LOC_616/Y NAND2X1_LOC_462/B 0.00fF
C30558 NOR2X1_LOC_590/A INVX1_LOC_65/A 1.39fF
C30559 NOR2X1_LOC_71/Y NOR2X1_LOC_84/Y 0.19fF
C30560 NOR2X1_LOC_315/Y NOR2X1_LOC_76/A 0.70fF
C30561 NOR2X1_LOC_401/A NOR2X1_LOC_266/B 0.05fF
C30562 INVX1_LOC_64/A NAND2X1_LOC_93/B 1.75fF
C30563 INVX1_LOC_256/A INVX1_LOC_20/A 0.00fF
C30564 NOR2X1_LOC_68/A NOR2X1_LOC_377/a_36_216# 0.00fF
C30565 INVX1_LOC_22/Y INVX1_LOC_65/A 0.00fF
C30566 NOR2X1_LOC_827/a_36_216# INVX1_LOC_89/A 0.00fF
C30567 NOR2X1_LOC_250/Y NAND2X1_LOC_211/Y 0.01fF
C30568 NOR2X1_LOC_309/Y NAND2X1_LOC_842/B 0.02fF
C30569 INVX1_LOC_5/A INVX1_LOC_108/A 0.01fF
C30570 NOR2X1_LOC_169/B NOR2X1_LOC_552/A 0.01fF
C30571 NAND2X1_LOC_364/A INVX1_LOC_186/A 0.14fF
C30572 INVX1_LOC_13/A INVX1_LOC_137/A 0.00fF
C30573 INVX1_LOC_206/A INVX1_LOC_55/Y 0.00fF
C30574 INVX1_LOC_26/A NAND2X1_LOC_74/B 0.10fF
C30575 NOR2X1_LOC_65/B INVX1_LOC_19/A 0.06fF
C30576 NOR2X1_LOC_433/A INVX1_LOC_311/A 0.14fF
C30577 INVX1_LOC_17/A INVX1_LOC_117/A 0.07fF
C30578 INVX1_LOC_290/Y NOR2X1_LOC_465/Y 0.27fF
C30579 NOR2X1_LOC_160/B NOR2X1_LOC_266/B 0.03fF
C30580 NAND2X1_LOC_63/Y NOR2X1_LOC_621/A 0.04fF
C30581 INVX1_LOC_8/Y NOR2X1_LOC_9/Y 0.01fF
C30582 NAND2X1_LOC_308/Y NAND2X1_LOC_863/A 0.09fF
C30583 INVX1_LOC_135/A NOR2X1_LOC_375/Y 0.02fF
C30584 NOR2X1_LOC_593/Y INVX1_LOC_311/A 0.03fF
C30585 NAND2X1_LOC_327/a_36_24# NOR2X1_LOC_52/B 0.00fF
C30586 D_INPUT_0 NOR2X1_LOC_516/B 0.08fF
C30587 INVX1_LOC_177/A NOR2X1_LOC_703/A 0.01fF
C30588 INVX1_LOC_35/Y NOR2X1_LOC_291/Y 0.02fF
C30589 NOR2X1_LOC_644/B INVX1_LOC_14/Y 0.18fF
C30590 INVX1_LOC_135/A NOR2X1_LOC_719/A 0.01fF
C30591 NAND2X1_LOC_454/Y NOR2X1_LOC_270/a_36_216# 0.01fF
C30592 NOR2X1_LOC_113/B NOR2X1_LOC_142/Y 0.02fF
C30593 NAND2X1_LOC_9/Y INVX1_LOC_63/A 0.11fF
C30594 NAND2X1_LOC_563/A INPUT_1 0.03fF
C30595 INVX1_LOC_64/A INVX1_LOC_3/A 0.03fF
C30596 NAND2X1_LOC_476/Y NOR2X1_LOC_678/A 0.01fF
C30597 NOR2X1_LOC_471/Y INVX1_LOC_117/A 0.08fF
C30598 NAND2X1_LOC_364/A NAND2X1_LOC_447/Y 0.10fF
C30599 INVX1_LOC_233/A INVX1_LOC_63/A 0.08fF
C30600 NOR2X1_LOC_809/a_36_216# INVX1_LOC_83/A 0.00fF
C30601 NAND2X1_LOC_564/A NAND2X1_LOC_74/B 0.01fF
C30602 NAND2X1_LOC_550/A NAND2X1_LOC_848/A 0.12fF
C30603 INVX1_LOC_48/Y INVX1_LOC_89/Y 0.01fF
C30604 NOR2X1_LOC_52/B INVX1_LOC_311/A 0.01fF
C30605 NAND2X1_LOC_456/a_36_24# NAND2X1_LOC_99/A 0.00fF
C30606 INVX1_LOC_135/A INVX1_LOC_7/A 0.06fF
C30607 NOR2X1_LOC_328/Y NOR2X1_LOC_597/A 0.06fF
C30608 NOR2X1_LOC_78/B NOR2X1_LOC_742/A 0.10fF
C30609 NOR2X1_LOC_440/Y INVX1_LOC_171/A 0.02fF
C30610 INVX1_LOC_237/A INVX1_LOC_260/A 0.01fF
C30611 INVX1_LOC_279/A INVX1_LOC_89/A 0.07fF
C30612 INVX1_LOC_1/A INVX1_LOC_179/A 0.10fF
C30613 NAND2X1_LOC_35/Y NAND2X1_LOC_773/B 0.03fF
C30614 INVX1_LOC_177/Y VDD 0.09fF
C30615 INVX1_LOC_24/A NOR2X1_LOC_538/a_36_216# 0.02fF
C30616 INVX1_LOC_104/A NOR2X1_LOC_337/Y 0.02fF
C30617 INVX1_LOC_77/A INVX1_LOC_199/Y 0.05fF
C30618 INVX1_LOC_75/A NAND2X1_LOC_841/A 0.11fF
C30619 INVX1_LOC_103/A INVX1_LOC_307/A 0.11fF
C30620 INVX1_LOC_215/A INVX1_LOC_28/A 0.07fF
C30621 NOR2X1_LOC_798/A INVX1_LOC_63/A 0.05fF
C30622 INVX1_LOC_13/A NOR2X1_LOC_19/B 1.51fF
C30623 NOR2X1_LOC_215/Y VDD -0.00fF
C30624 NOR2X1_LOC_564/a_36_216# INVX1_LOC_177/A 0.00fF
C30625 NOR2X1_LOC_503/Y NOR2X1_LOC_508/a_36_216# 0.02fF
C30626 NAND2X1_LOC_850/Y INVX1_LOC_126/Y 0.03fF
C30627 INVX1_LOC_249/A NOR2X1_LOC_357/Y 0.80fF
C30628 INVX1_LOC_268/A INVX1_LOC_75/A 0.00fF
C30629 INVX1_LOC_13/Y NAND2X1_LOC_772/a_36_24# 0.00fF
C30630 NOR2X1_LOC_824/A NAND2X1_LOC_489/Y 0.05fF
C30631 INVX1_LOC_271/A INVX1_LOC_32/A 0.73fF
C30632 INVX1_LOC_14/A NAND2X1_LOC_572/B 0.27fF
C30633 INVX1_LOC_50/Y NOR2X1_LOC_509/A 0.02fF
C30634 INVX1_LOC_33/A NAND2X1_LOC_469/B 0.03fF
C30635 INVX1_LOC_43/Y NAND2X1_LOC_93/B 0.01fF
C30636 NOR2X1_LOC_52/B INVX1_LOC_304/A 0.18fF
C30637 NAND2X1_LOC_337/B NOR2X1_LOC_841/A 0.10fF
C30638 NOR2X1_LOC_78/B NOR2X1_LOC_318/B 0.03fF
C30639 INVX1_LOC_58/A NOR2X1_LOC_158/B 0.00fF
C30640 NOR2X1_LOC_742/A INVX1_LOC_83/A 0.76fF
C30641 INVX1_LOC_286/A INVX1_LOC_16/A 0.07fF
C30642 NOR2X1_LOC_52/B NOR2X1_LOC_670/Y 0.19fF
C30643 NOR2X1_LOC_473/B NOR2X1_LOC_329/B 0.01fF
C30644 NOR2X1_LOC_282/Y NAND2X1_LOC_286/B 0.07fF
C30645 INVX1_LOC_77/A INVX1_LOC_281/A 0.07fF
C30646 NOR2X1_LOC_315/Y NAND2X1_LOC_241/Y 0.05fF
C30647 NAND2X1_LOC_638/Y NAND2X1_LOC_654/B 0.00fF
C30648 INVX1_LOC_271/A NAND2X1_LOC_175/Y 0.01fF
C30649 NOR2X1_LOC_489/a_36_216# INVX1_LOC_47/Y 0.00fF
C30650 NOR2X1_LOC_78/B INVX1_LOC_93/Y 0.07fF
C30651 INVX1_LOC_15/A NAND2X1_LOC_31/a_36_24# 0.00fF
C30652 INVX1_LOC_21/A NAND2X1_LOC_254/Y 0.03fF
C30653 NOR2X1_LOC_598/B NOR2X1_LOC_334/Y 0.10fF
C30654 NOR2X1_LOC_140/A INVX1_LOC_29/A 0.00fF
C30655 NOR2X1_LOC_264/a_36_216# NAND2X1_LOC_63/Y 0.00fF
C30656 NAND2X1_LOC_35/Y NOR2X1_LOC_393/Y 0.05fF
C30657 INVX1_LOC_227/A INVX1_LOC_285/Y 0.10fF
C30658 NAND2X1_LOC_214/B INVX1_LOC_32/A 0.07fF
C30659 INVX1_LOC_213/Y INVX1_LOC_37/A 0.54fF
C30660 INVX1_LOC_104/A VDD 2.29fF
C30661 INVX1_LOC_90/A INVX1_LOC_302/Y 0.10fF
C30662 NOR2X1_LOC_91/A INVX1_LOC_224/Y 0.07fF
C30663 INVX1_LOC_136/A NOR2X1_LOC_79/Y 0.03fF
C30664 NOR2X1_LOC_220/A NOR2X1_LOC_486/Y 1.40fF
C30665 INVX1_LOC_135/A NOR2X1_LOC_167/Y 0.01fF
C30666 INVX1_LOC_97/Y NOR2X1_LOC_334/Y -0.03fF
C30667 INVX1_LOC_64/A NAND2X1_LOC_470/B 0.07fF
C30668 NAND2X1_LOC_149/Y NOR2X1_LOC_48/B 0.01fF
C30669 NAND2X1_LOC_156/a_36_24# INVX1_LOC_117/Y 0.00fF
C30670 NAND2X1_LOC_629/Y INVX1_LOC_139/Y 0.02fF
C30671 INVX1_LOC_95/Y INVX1_LOC_25/Y 0.03fF
C30672 INVX1_LOC_27/A INVX1_LOC_32/A 0.80fF
C30673 INVX1_LOC_103/A INVX1_LOC_12/A 0.41fF
C30674 NAND2X1_LOC_715/B NOR2X1_LOC_334/Y 0.65fF
C30675 INVX1_LOC_278/A NOR2X1_LOC_693/a_36_216# 0.01fF
C30676 INVX1_LOC_63/Y INVX1_LOC_38/A 0.03fF
C30677 NOR2X1_LOC_78/B INVX1_LOC_139/A 0.01fF
C30678 NOR2X1_LOC_218/Y NOR2X1_LOC_275/A 0.00fF
C30679 NAND2X1_LOC_850/A NOR2X1_LOC_74/A 0.17fF
C30680 INVX1_LOC_224/Y INVX1_LOC_23/A 0.10fF
C30681 NOR2X1_LOC_91/A NAND2X1_LOC_793/B 0.01fF
C30682 NOR2X1_LOC_530/Y INVX1_LOC_29/A 0.03fF
C30683 NOR2X1_LOC_374/A INVX1_LOC_307/Y 0.01fF
C30684 INVX1_LOC_93/Y NAND2X1_LOC_392/Y 0.00fF
C30685 NOR2X1_LOC_355/A NOR2X1_LOC_78/A 0.03fF
C30686 NOR2X1_LOC_544/A NOR2X1_LOC_858/B 0.04fF
C30687 NOR2X1_LOC_61/a_36_216# INVX1_LOC_280/A 0.00fF
C30688 INVX1_LOC_77/A NOR2X1_LOC_862/B 0.13fF
C30689 NOR2X1_LOC_226/A INVX1_LOC_12/Y 0.10fF
C30690 INVX1_LOC_292/A INVX1_LOC_12/A 0.03fF
C30691 INVX1_LOC_174/A NOR2X1_LOC_89/A 0.09fF
C30692 INVX1_LOC_263/A VDD 0.03fF
C30693 INVX1_LOC_161/Y INVX1_LOC_42/A 0.03fF
C30694 NAND2X1_LOC_479/Y INVX1_LOC_76/A 0.07fF
C30695 NOR2X1_LOC_175/A INVX1_LOC_38/A 0.07fF
C30696 NOR2X1_LOC_431/Y NOR2X1_LOC_697/Y 0.01fF
C30697 INVX1_LOC_227/A NOR2X1_LOC_137/B 0.02fF
C30698 NAND2X1_LOC_84/Y NAND2X1_LOC_572/B 0.01fF
C30699 INVX1_LOC_1/Y INVX1_LOC_46/A 0.14fF
C30700 NAND2X1_LOC_550/A NOR2X1_LOC_754/A 0.08fF
C30701 INVX1_LOC_17/A INVX1_LOC_3/Y 0.00fF
C30702 NAND2X1_LOC_850/Y NOR2X1_LOC_536/A 0.07fF
C30703 NOR2X1_LOC_218/Y INVX1_LOC_12/Y 0.14fF
C30704 NOR2X1_LOC_554/B INVX1_LOC_19/A 0.15fF
C30705 NOR2X1_LOC_516/B NOR2X1_LOC_859/Y 0.06fF
C30706 INVX1_LOC_269/A NAND2X1_LOC_618/Y 0.02fF
C30707 INVX1_LOC_41/A NOR2X1_LOC_197/B 0.03fF
C30708 NAND2X1_LOC_112/Y NOR2X1_LOC_111/A 0.05fF
C30709 INVX1_LOC_177/Y INVX1_LOC_133/A 0.00fF
C30710 NAND2X1_LOC_854/B VDD 0.06fF
C30711 NOR2X1_LOC_637/a_36_216# NOR2X1_LOC_697/Y 0.00fF
C30712 NOR2X1_LOC_464/B NOR2X1_LOC_464/Y 0.01fF
C30713 INVX1_LOC_10/A NOR2X1_LOC_137/Y 0.03fF
C30714 INVX1_LOC_57/A INVX1_LOC_306/Y 0.07fF
C30715 INVX1_LOC_135/A INVX1_LOC_76/A 0.19fF
C30716 INVX1_LOC_256/A INVX1_LOC_4/A 0.37fF
C30717 INVX1_LOC_63/Y NOR2X1_LOC_697/a_36_216# 0.00fF
C30718 NOR2X1_LOC_751/Y NOR2X1_LOC_641/a_36_216# 0.00fF
C30719 INVX1_LOC_48/Y INVX1_LOC_16/Y 0.03fF
C30720 NOR2X1_LOC_599/A INVX1_LOC_42/A 0.07fF
C30721 NAND2X1_LOC_555/Y INVX1_LOC_3/Y 0.17fF
C30722 D_INPUT_0 NAND2X1_LOC_211/Y 0.03fF
C30723 INVX1_LOC_11/A NOR2X1_LOC_248/A 0.08fF
C30724 INVX1_LOC_10/A NOR2X1_LOC_822/a_36_216# 0.00fF
C30725 INVX1_LOC_65/A NOR2X1_LOC_703/A 0.01fF
C30726 INVX1_LOC_295/A INVX1_LOC_76/A 0.04fF
C30727 NOR2X1_LOC_720/B NAND2X1_LOC_85/Y 0.02fF
C30728 NOR2X1_LOC_231/B INVX1_LOC_15/A 0.03fF
C30729 NAND2X1_LOC_860/A NOR2X1_LOC_291/Y 0.18fF
C30730 NAND2X1_LOC_549/a_36_24# INVX1_LOC_84/A 0.00fF
C30731 NOR2X1_LOC_719/A INVX1_LOC_280/A 0.01fF
C30732 NOR2X1_LOC_152/Y INVX1_LOC_19/A 0.07fF
C30733 INVX1_LOC_161/Y INVX1_LOC_78/A 0.28fF
C30734 NAND2X1_LOC_181/Y NOR2X1_LOC_118/a_36_216# 0.00fF
C30735 NOR2X1_LOC_843/A NOR2X1_LOC_814/A 0.14fF
C30736 NOR2X1_LOC_606/Y INVX1_LOC_4/A 0.03fF
C30737 NOR2X1_LOC_753/Y INVX1_LOC_49/Y 0.00fF
C30738 NOR2X1_LOC_590/A INVX1_LOC_4/Y 0.17fF
C30739 INVX1_LOC_50/A NAND2X1_LOC_780/Y 0.02fF
C30740 NOR2X1_LOC_438/a_36_216# NOR2X1_LOC_438/Y 0.00fF
C30741 NAND2X1_LOC_374/Y NAND2X1_LOC_244/a_36_24# 0.00fF
C30742 INVX1_LOC_16/A INVX1_LOC_54/A 0.99fF
C30743 INVX1_LOC_48/Y NAND2X1_LOC_205/A 0.10fF
C30744 INVX1_LOC_75/A INVX1_LOC_95/Y 0.07fF
C30745 INVX1_LOC_7/A INVX1_LOC_280/A 0.06fF
C30746 NOR2X1_LOC_552/Y NOR2X1_LOC_78/A 0.04fF
C30747 NAND2X1_LOC_735/B NOR2X1_LOC_629/Y 0.05fF
C30748 NOR2X1_LOC_91/A NOR2X1_LOC_103/Y 0.03fF
C30749 NAND2X1_LOC_325/Y INVX1_LOC_49/Y 0.00fF
C30750 INVX1_LOC_12/Y INPUT_1 0.09fF
C30751 INVX1_LOC_75/A NOR2X1_LOC_33/a_36_216# -0.02fF
C30752 INVX1_LOC_81/Y NAND2X1_LOC_454/Y 0.01fF
C30753 NOR2X1_LOC_202/Y INVX1_LOC_76/A 0.03fF
C30754 NAND2X1_LOC_588/B D_INPUT_5 0.01fF
C30755 INVX1_LOC_59/A NOR2X1_LOC_392/Y 0.01fF
C30756 INVX1_LOC_272/Y NOR2X1_LOC_677/Y 0.02fF
C30757 NAND2X1_LOC_465/Y NAND2X1_LOC_773/B 0.02fF
C30758 NOR2X1_LOC_65/B INVX1_LOC_161/Y 0.00fF
C30759 INVX1_LOC_311/A INVX1_LOC_199/A 0.12fF
C30760 INVX1_LOC_8/A INVX1_LOC_125/A 0.05fF
C30761 NOR2X1_LOC_754/a_36_216# NOR2X1_LOC_253/Y 0.00fF
C30762 NOR2X1_LOC_211/A NOR2X1_LOC_197/B 0.03fF
C30763 INVX1_LOC_58/A INVX1_LOC_17/A 0.13fF
C30764 INVX1_LOC_72/A NOR2X1_LOC_80/Y 0.29fF
C30765 INVX1_LOC_104/A INVX1_LOC_133/A 0.10fF
C30766 INVX1_LOC_64/A NOR2X1_LOC_348/Y 0.02fF
C30767 NOR2X1_LOC_103/Y INVX1_LOC_23/A 0.07fF
C30768 INVX1_LOC_50/A NAND2X1_LOC_114/B 0.07fF
C30769 NOR2X1_LOC_541/Y INVX1_LOC_23/A 0.07fF
C30770 NAND2X1_LOC_161/a_36_24# NOR2X1_LOC_467/A 0.01fF
C30771 NAND2X1_LOC_840/Y NOR2X1_LOC_111/A 0.06fF
C30772 NOR2X1_LOC_262/Y INVX1_LOC_47/Y 0.04fF
C30773 NOR2X1_LOC_332/A INVX1_LOC_108/A 0.03fF
C30774 NOR2X1_LOC_721/A INVX1_LOC_19/A 0.01fF
C30775 NOR2X1_LOC_479/B INVX1_LOC_84/A 0.00fF
C30776 NOR2X1_LOC_192/A NAND2X1_LOC_642/Y 0.01fF
C30777 INVX1_LOC_276/A INVX1_LOC_49/Y 0.30fF
C30778 NOR2X1_LOC_91/A INVX1_LOC_45/A 0.01fF
C30779 INVX1_LOC_134/A INVX1_LOC_53/A 0.01fF
C30780 INVX1_LOC_224/Y INVX1_LOC_31/A 0.07fF
C30781 INVX1_LOC_83/A INVX1_LOC_117/Y 0.05fF
C30782 INVX1_LOC_136/A INVX1_LOC_26/A 0.37fF
C30783 NOR2X1_LOC_328/Y INVX1_LOC_84/A 0.03fF
C30784 INVX1_LOC_277/A NOR2X1_LOC_383/B 0.00fF
C30785 NOR2X1_LOC_307/B INVX1_LOC_19/A 0.03fF
C30786 NAND2X1_LOC_306/a_36_24# INVX1_LOC_94/Y 0.00fF
C30787 INVX1_LOC_89/A NOR2X1_LOC_624/B 0.01fF
C30788 INVX1_LOC_206/Y VDD 0.60fF
C30789 NOR2X1_LOC_460/Y INVX1_LOC_198/A 0.21fF
C30790 INVX1_LOC_256/A INVX1_LOC_64/A 0.21fF
C30791 INVX1_LOC_50/A INVX1_LOC_312/Y 0.07fF
C30792 INVX1_LOC_28/A INVX1_LOC_54/A 0.31fF
C30793 INVX1_LOC_282/A NOR2X1_LOC_536/A 0.37fF
C30794 NOR2X1_LOC_405/A NAND2X1_LOC_447/Y 0.01fF
C30795 NOR2X1_LOC_577/Y NOR2X1_LOC_681/a_36_216# 0.01fF
C30796 NOR2X1_LOC_758/a_36_216# NOR2X1_LOC_278/Y 0.01fF
C30797 INVX1_LOC_86/Y VDD 0.25fF
C30798 INVX1_LOC_186/A NOR2X1_LOC_857/A 0.07fF
C30799 INVX1_LOC_72/A INVX1_LOC_270/A 2.54fF
C30800 INVX1_LOC_39/A INVX1_LOC_269/A 0.01fF
C30801 NOR2X1_LOC_664/Y INVX1_LOC_32/A 0.02fF
C30802 INVX1_LOC_45/A INVX1_LOC_23/A 0.29fF
C30803 NAND2X1_LOC_9/Y NOR2X1_LOC_606/a_36_216# 0.00fF
C30804 INVX1_LOC_31/A NAND2X1_LOC_793/B 0.07fF
C30805 NOR2X1_LOC_173/Y NAND2X1_LOC_175/a_36_24# 0.00fF
C30806 NOR2X1_LOC_318/B INVX1_LOC_46/A 0.10fF
C30807 NAND2X1_LOC_36/A INVX1_LOC_53/A 0.01fF
C30808 INVX1_LOC_57/Y NAND2X1_LOC_784/A 0.06fF
C30809 NOR2X1_LOC_130/A NOR2X1_LOC_435/B 0.01fF
C30810 NAND2X1_LOC_793/Y NOR2X1_LOC_652/Y 0.02fF
C30811 INVX1_LOC_219/A INVX1_LOC_84/A 0.04fF
C30812 NOR2X1_LOC_626/Y INVX1_LOC_11/A 0.61fF
C30813 NOR2X1_LOC_91/A INVX1_LOC_71/A 0.03fF
C30814 VDD NOR2X1_LOC_600/Y 0.24fF
C30815 NAND2X1_LOC_214/B INPUT_3 0.07fF
C30816 NOR2X1_LOC_458/B INVX1_LOC_290/Y 0.04fF
C30817 INVX1_LOC_93/Y INVX1_LOC_46/A 0.07fF
C30818 NOR2X1_LOC_706/a_36_216# INVX1_LOC_91/A 0.00fF
C30819 NOR2X1_LOC_251/a_36_216# NOR2X1_LOC_361/B 0.02fF
C30820 NOR2X1_LOC_237/Y NOR2X1_LOC_134/a_36_216# 0.00fF
C30821 D_INPUT_1 NOR2X1_LOC_607/A 0.01fF
C30822 NOR2X1_LOC_790/B NOR2X1_LOC_68/A 0.10fF
C30823 NAND2X1_LOC_514/Y INVX1_LOC_53/A 0.02fF
C30824 INVX1_LOC_18/A NOR2X1_LOC_678/A 0.03fF
C30825 INVX1_LOC_144/A NAND2X1_LOC_434/Y 0.02fF
C30826 INVX1_LOC_27/A INPUT_3 0.34fF
C30827 NOR2X1_LOC_589/A NOR2X1_LOC_89/A 0.39fF
C30828 NAND2X1_LOC_153/a_36_24# INVX1_LOC_53/A 0.00fF
C30829 NAND2X1_LOC_551/A NAND2X1_LOC_477/Y 0.03fF
C30830 INVX1_LOC_71/A INVX1_LOC_23/A 0.16fF
C30831 INVX1_LOC_16/A NOR2X1_LOC_48/B 0.29fF
C30832 NOR2X1_LOC_60/a_36_216# INVX1_LOC_272/A 0.01fF
C30833 INVX1_LOC_41/Y NOR2X1_LOC_754/Y 0.00fF
C30834 INVX1_LOC_40/A INVX1_LOC_251/A 0.03fF
C30835 NOR2X1_LOC_251/Y INVX1_LOC_32/A -0.00fF
C30836 NOR2X1_LOC_624/A NOR2X1_LOC_621/A 0.29fF
C30837 NAND2X1_LOC_842/B INVX1_LOC_63/A 0.07fF
C30838 NOR2X1_LOC_479/B INVX1_LOC_15/A 0.00fF
C30839 NAND2X1_LOC_740/Y NAND2X1_LOC_741/B 0.00fF
C30840 NOR2X1_LOC_278/A INVX1_LOC_26/A 0.03fF
C30841 D_INPUT_0 NAND2X1_LOC_207/B 0.05fF
C30842 NAND2X1_LOC_222/B NAND2X1_LOC_19/a_36_24# 0.01fF
C30843 INVX1_LOC_50/A NOR2X1_LOC_219/B 0.03fF
C30844 INVX1_LOC_168/A NOR2X1_LOC_278/Y 0.04fF
C30845 INVX1_LOC_50/A NAND2X1_LOC_483/Y 0.00fF
C30846 NOR2X1_LOC_366/Y INVX1_LOC_109/Y 0.05fF
C30847 NAND2X1_LOC_35/Y INVX1_LOC_24/A 0.08fF
C30848 NAND2X1_LOC_721/A INVX1_LOC_46/A 0.03fF
C30849 NOR2X1_LOC_813/Y INVX1_LOC_76/A 0.49fF
C30850 NOR2X1_LOC_92/Y INVX1_LOC_286/Y 0.07fF
C30851 INVX1_LOC_17/A INVX1_LOC_215/Y 0.69fF
C30852 INVX1_LOC_294/Y INVX1_LOC_57/A 0.03fF
C30853 INVX1_LOC_171/A NOR2X1_LOC_89/A 0.04fF
C30854 NOR2X1_LOC_152/A INVX1_LOC_76/A 0.01fF
C30855 INVX1_LOC_247/A INVX1_LOC_9/A 0.03fF
C30856 INVX1_LOC_11/A INVX1_LOC_174/A 0.72fF
C30857 NAND2X1_LOC_231/Y NAND2X1_LOC_61/Y 0.15fF
C30858 INVX1_LOC_225/A INVX1_LOC_29/Y 0.07fF
C30859 INVX1_LOC_183/Y INVX1_LOC_102/A 0.02fF
C30860 NOR2X1_LOC_641/B INVX1_LOC_1/A 0.07fF
C30861 NOR2X1_LOC_459/B NOR2X1_LOC_476/B 0.19fF
C30862 INVX1_LOC_234/A INVX1_LOC_32/A 0.04fF
C30863 NOR2X1_LOC_455/Y NOR2X1_LOC_388/Y 0.05fF
C30864 NOR2X1_LOC_687/Y NOR2X1_LOC_685/B 0.01fF
C30865 NOR2X1_LOC_706/B INVX1_LOC_117/A 0.00fF
C30866 NAND2X1_LOC_725/A INVX1_LOC_209/Y 0.02fF
C30867 NOR2X1_LOC_74/A NOR2X1_LOC_662/A 0.02fF
C30868 NOR2X1_LOC_351/Y NAND2X1_LOC_469/B 0.00fF
C30869 NAND2X1_LOC_568/A INVX1_LOC_286/Y 0.02fF
C30870 NOR2X1_LOC_134/Y NAND2X1_LOC_550/A 0.01fF
C30871 NOR2X1_LOC_570/A NOR2X1_LOC_334/Y 0.04fF
C30872 NOR2X1_LOC_84/Y NAND2X1_LOC_205/A 0.18fF
C30873 NAND2X1_LOC_21/Y NAND2X1_LOC_31/a_36_24# 0.00fF
C30874 NOR2X1_LOC_751/Y INVX1_LOC_1/A 0.00fF
C30875 INVX1_LOC_140/A INPUT_7 0.44fF
C30876 NOR2X1_LOC_597/a_36_216# INVX1_LOC_12/A 0.00fF
C30877 NAND2X1_LOC_181/Y INVX1_LOC_181/A 0.01fF
C30878 NOR2X1_LOC_719/a_36_216# NOR2X1_LOC_38/B 0.00fF
C30879 INVX1_LOC_21/A INVX1_LOC_314/Y 0.07fF
C30880 INVX1_LOC_64/Y NOR2X1_LOC_260/Y 0.20fF
C30881 NAND2X1_LOC_326/A NOR2X1_LOC_512/Y 0.05fF
C30882 INVX1_LOC_28/A NOR2X1_LOC_48/B 0.14fF
C30883 NOR2X1_LOC_755/a_36_216# INVX1_LOC_290/Y -0.00fF
C30884 NOR2X1_LOC_537/Y NOR2X1_LOC_416/A 0.07fF
C30885 INVX1_LOC_5/A NOR2X1_LOC_147/B 0.03fF
C30886 NOR2X1_LOC_15/Y INVX1_LOC_181/Y 0.26fF
C30887 NOR2X1_LOC_542/B NOR2X1_LOC_445/B 0.01fF
C30888 NOR2X1_LOC_368/A NAND2X1_LOC_74/B 0.02fF
C30889 INVX1_LOC_39/Y INVX1_LOC_61/Y 0.03fF
C30890 INVX1_LOC_228/A NOR2X1_LOC_140/A 0.46fF
C30891 NOR2X1_LOC_232/Y INVX1_LOC_61/A 0.07fF
C30892 INVX1_LOC_89/A NOR2X1_LOC_38/B 0.10fF
C30893 NOR2X1_LOC_626/Y NOR2X1_LOC_593/Y 0.01fF
C30894 NOR2X1_LOC_361/B NAND2X1_LOC_357/a_36_24# 0.01fF
C30895 INVX1_LOC_12/Y INVX1_LOC_118/A 0.10fF
C30896 NOR2X1_LOC_459/A INVX1_LOC_175/A 1.25fF
C30897 NOR2X1_LOC_644/A NOR2X1_LOC_801/B 0.00fF
C30898 NOR2X1_LOC_68/A D_GATE_741 0.11fF
C30899 INVX1_LOC_143/Y NOR2X1_LOC_445/B 0.02fF
C30900 NOR2X1_LOC_19/B INVX1_LOC_32/A 0.24fF
C30901 INVX1_LOC_256/A INVX1_LOC_130/Y 0.01fF
C30902 INVX1_LOC_45/A INVX1_LOC_31/A 0.18fF
C30903 INVX1_LOC_46/A INVX1_LOC_117/Y 0.03fF
C30904 INVX1_LOC_55/A INVX1_LOC_18/A 0.04fF
C30905 INVX1_LOC_20/A INVX1_LOC_297/A 0.12fF
C30906 INVX1_LOC_255/Y INVX1_LOC_25/A 0.21fF
C30907 NOR2X1_LOC_819/a_36_216# INVX1_LOC_31/A 0.01fF
C30908 NAND2X1_LOC_354/a_36_24# NAND2X1_LOC_354/Y 0.02fF
C30909 NOR2X1_LOC_276/B NOR2X1_LOC_276/Y -0.00fF
C30910 NOR2X1_LOC_230/a_36_216# INVX1_LOC_72/A 0.00fF
C30911 INVX1_LOC_14/A NOR2X1_LOC_716/B 0.14fF
C30912 INVX1_LOC_46/A NAND2X1_LOC_770/Y 1.98fF
C30913 NOR2X1_LOC_196/Y INVX1_LOC_15/A 0.01fF
C30914 NAND2X1_LOC_472/Y NOR2X1_LOC_155/A 0.01fF
C30915 INVX1_LOC_50/A NAND2X1_LOC_656/Y 0.30fF
C30916 NAND2X1_LOC_573/Y NAND2X1_LOC_840/a_36_24# 0.00fF
C30917 INVX1_LOC_161/Y NOR2X1_LOC_152/Y 1.98fF
C30918 NOR2X1_LOC_76/A NAND2X1_LOC_99/A 0.04fF
C30919 NOR2X1_LOC_294/a_36_216# NOR2X1_LOC_554/B 0.00fF
C30920 INVX1_LOC_36/A INVX1_LOC_72/A 1.04fF
C30921 INVX1_LOC_233/A INVX1_LOC_1/Y 0.03fF
C30922 INVX1_LOC_33/Y NOR2X1_LOC_88/Y 0.03fF
C30923 NOR2X1_LOC_439/B INVX1_LOC_271/Y 0.04fF
C30924 INVX1_LOC_223/A NOR2X1_LOC_703/B 0.94fF
C30925 NOR2X1_LOC_15/Y NOR2X1_LOC_192/a_36_216# 0.00fF
C30926 NAND2X1_LOC_562/Y INVX1_LOC_269/A 0.02fF
C30927 NAND2X1_LOC_303/B INVX1_LOC_173/A 0.03fF
C30928 NAND2X1_LOC_859/Y NAND2X1_LOC_793/B 0.01fF
C30929 INVX1_LOC_102/A INVX1_LOC_91/A 0.07fF
C30930 NAND2X1_LOC_35/Y NAND2X1_LOC_565/B 0.01fF
C30931 INVX1_LOC_21/A NOR2X1_LOC_778/B 0.07fF
C30932 INVX1_LOC_31/A INVX1_LOC_71/A 0.01fF
C30933 INVX1_LOC_75/A INVX1_LOC_271/Y 0.07fF
C30934 NOR2X1_LOC_160/B INVX1_LOC_49/A 0.27fF
C30935 NOR2X1_LOC_272/Y NAND2X1_LOC_541/Y 0.16fF
C30936 NOR2X1_LOC_766/Y NAND2X1_LOC_770/Y 0.07fF
C30937 NOR2X1_LOC_765/Y INVX1_LOC_297/A 0.17fF
C30938 NOR2X1_LOC_123/B INVX1_LOC_23/A 0.07fF
C30939 NAND2X1_LOC_228/a_36_24# INVX1_LOC_5/A 0.00fF
C30940 INVX1_LOC_39/A NAND2X1_LOC_563/A 0.01fF
C30941 INVX1_LOC_313/Y INVX1_LOC_270/A 0.03fF
C30942 INVX1_LOC_69/Y INVX1_LOC_4/A 0.07fF
C30943 NAND2X1_LOC_550/a_36_24# INVX1_LOC_13/Y 0.00fF
C30944 NOR2X1_LOC_82/A INVX1_LOC_80/Y 0.02fF
C30945 NOR2X1_LOC_356/A INVX1_LOC_57/A 0.02fF
C30946 NOR2X1_LOC_91/A INVX1_LOC_102/Y 0.02fF
C30947 NOR2X1_LOC_798/A INVX1_LOC_1/Y 0.05fF
C30948 NOR2X1_LOC_208/Y INVX1_LOC_72/A 0.01fF
C30949 NAND2X1_LOC_9/Y NOR2X1_LOC_559/a_36_216# 0.01fF
C30950 NOR2X1_LOC_664/Y INPUT_3 0.53fF
C30951 NOR2X1_LOC_843/A NOR2X1_LOC_590/A 0.03fF
C30952 NOR2X1_LOC_89/A INVX1_LOC_20/A 0.30fF
C30953 INVX1_LOC_59/A INVX1_LOC_25/Y 0.01fF
C30954 INVX1_LOC_88/A NOR2X1_LOC_757/a_36_216# 0.00fF
C30955 NOR2X1_LOC_196/A NAND2X1_LOC_48/a_36_24# 0.00fF
C30956 NAND2X1_LOC_35/Y NOR2X1_LOC_130/A 0.07fF
C30957 NAND2X1_LOC_866/B NAND2X1_LOC_793/B 0.01fF
C30958 NOR2X1_LOC_226/A NOR2X1_LOC_401/A 0.04fF
C30959 INVX1_LOC_188/A NOR2X1_LOC_348/B 0.02fF
C30960 INVX1_LOC_2/A NAND2X1_LOC_550/A 0.07fF
C30961 NAND2X1_LOC_733/Y INVX1_LOC_240/A 0.26fF
C30962 INVX1_LOC_102/Y INVX1_LOC_23/A 0.07fF
C30963 INVX1_LOC_174/Y NOR2X1_LOC_463/a_36_216# 0.00fF
C30964 INVX1_LOC_134/A NOR2X1_LOC_634/B 0.02fF
C30965 NOR2X1_LOC_82/A NOR2X1_LOC_78/B 0.03fF
C30966 INVX1_LOC_5/A INVX1_LOC_97/A 0.02fF
C30967 INVX1_LOC_2/A NOR2X1_LOC_160/B 0.17fF
C30968 INVX1_LOC_134/A NOR2X1_LOC_78/B 0.05fF
C30969 INVX1_LOC_85/Y INVX1_LOC_213/A 0.04fF
C30970 INVX1_LOC_256/A NAND2X1_LOC_850/Y 0.02fF
C30971 INVX1_LOC_255/Y INVX1_LOC_1/A 0.07fF
C30972 NOR2X1_LOC_255/a_36_216# INVX1_LOC_48/Y 0.00fF
C30973 NAND2X1_LOC_552/A INVX1_LOC_90/A 0.00fF
C30974 INVX1_LOC_37/A NOR2X1_LOC_470/a_36_216# 0.00fF
C30975 NOR2X1_LOC_74/A INVX1_LOC_57/A 0.24fF
C30976 NOR2X1_LOC_420/Y INVX1_LOC_89/A 0.01fF
C30977 INVX1_LOC_5/A INVX1_LOC_90/A 0.18fF
C30978 NOR2X1_LOC_226/A NOR2X1_LOC_160/B 0.20fF
C30979 INVX1_LOC_269/A NAND2X1_LOC_735/B 0.02fF
C30980 INVX1_LOC_58/A NOR2X1_LOC_594/Y 0.27fF
C30981 NOR2X1_LOC_309/Y INVX1_LOC_72/A 0.01fF
C30982 NAND2X1_LOC_817/a_36_24# NOR2X1_LOC_649/B -0.01fF
C30983 NOR2X1_LOC_102/a_36_216# INVX1_LOC_284/A 0.01fF
C30984 NOR2X1_LOC_9/Y INVX1_LOC_57/A 0.13fF
C30985 INVX1_LOC_224/Y INVX1_LOC_6/A 0.17fF
C30986 INVX1_LOC_303/A NAND2X1_LOC_7/Y 0.02fF
C30987 NAND2X1_LOC_84/Y NOR2X1_LOC_716/B 0.00fF
C30988 INVX1_LOC_217/A INVX1_LOC_240/A 0.15fF
C30989 INVX1_LOC_61/A NAND2X1_LOC_137/a_36_24# 0.00fF
C30990 NOR2X1_LOC_363/Y NAND2X1_LOC_792/B 0.15fF
C30991 NOR2X1_LOC_296/Y INVX1_LOC_137/A 0.03fF
C30992 INVX1_LOC_135/A INVX1_LOC_163/A 0.96fF
C30993 NOR2X1_LOC_67/A NAND2X1_LOC_208/B 0.03fF
C30994 INVX1_LOC_41/A NOR2X1_LOC_191/B 0.00fF
C30995 NOR2X1_LOC_625/Y NAND2X1_LOC_632/B 0.12fF
C30996 INVX1_LOC_50/A INVX1_LOC_78/Y 0.01fF
C30997 INVX1_LOC_36/A NAND2X1_LOC_633/a_36_24# 0.00fF
C30998 INVX1_LOC_11/A NOR2X1_LOC_589/A 0.07fF
C30999 INVX1_LOC_90/A INVX1_LOC_178/A 0.06fF
C31000 NOR2X1_LOC_68/A NAND2X1_LOC_357/B 1.11fF
C31001 INVX1_LOC_136/A INVX1_LOC_149/A 0.10fF
C31002 INVX1_LOC_44/A NOR2X1_LOC_631/a_36_216# 0.00fF
C31003 INVX1_LOC_227/A NOR2X1_LOC_205/Y 0.02fF
C31004 INVX1_LOC_36/A NOR2X1_LOC_537/Y 0.03fF
C31005 NOR2X1_LOC_772/A INVX1_LOC_171/Y 0.11fF
C31006 INVX1_LOC_36/A NAND2X1_LOC_338/B 0.15fF
C31007 INVX1_LOC_1/A NOR2X1_LOC_71/Y 0.10fF
C31008 NOR2X1_LOC_82/A NAND2X1_LOC_392/Y 0.03fF
C31009 INVX1_LOC_291/A INVX1_LOC_19/A 0.07fF
C31010 INVX1_LOC_177/Y INVX1_LOC_177/A 0.14fF
C31011 INVX1_LOC_24/A NAND2X1_LOC_465/Y 0.45fF
C31012 NAND2X1_LOC_361/Y NAND2X1_LOC_364/Y 0.56fF
C31013 NOR2X1_LOC_234/Y INVX1_LOC_24/A 0.00fF
C31014 INVX1_LOC_188/A INVX1_LOC_22/A 0.01fF
C31015 INVX1_LOC_5/A NAND2X1_LOC_348/A 0.15fF
C31016 NAND2X1_LOC_656/a_36_24# INVX1_LOC_14/A 0.00fF
C31017 INVX1_LOC_33/Y INVX1_LOC_15/A 0.03fF
C31018 INVX1_LOC_21/A NAND2X1_LOC_123/Y 0.05fF
C31019 INVX1_LOC_64/A INVX1_LOC_69/Y 0.07fF
C31020 INVX1_LOC_87/A INVX1_LOC_46/A 0.03fF
C31021 INVX1_LOC_33/A INVX1_LOC_63/Y 0.03fF
C31022 NOR2X1_LOC_498/Y NAND2X1_LOC_486/a_36_24# 0.00fF
C31023 NOR2X1_LOC_78/B NAND2X1_LOC_514/Y 0.02fF
C31024 INVX1_LOC_163/A INVX1_LOC_169/Y 0.07fF
C31025 NOR2X1_LOC_596/A NOR2X1_LOC_493/B 0.07fF
C31026 NAND2X1_LOC_207/B INVX1_LOC_46/Y 0.07fF
C31027 NOR2X1_LOC_574/A NOR2X1_LOC_577/Y 0.04fF
C31028 NAND2X1_LOC_642/Y INVX1_LOC_29/Y 0.02fF
C31029 INVX1_LOC_240/A NAND2X1_LOC_787/B 0.60fF
C31030 INVX1_LOC_14/A NOR2X1_LOC_120/a_36_216# 0.01fF
C31031 NOR2X1_LOC_828/B INVX1_LOC_1/A 0.07fF
C31032 INVX1_LOC_90/A NAND2X1_LOC_337/B 0.11fF
C31033 INVX1_LOC_49/A INVX1_LOC_189/A 0.00fF
C31034 NAND2X1_LOC_550/A INPUT_1 0.19fF
C31035 NOR2X1_LOC_421/Y INVX1_LOC_296/Y 0.03fF
C31036 INVX1_LOC_90/A NOR2X1_LOC_816/A 0.07fF
C31037 NAND2X1_LOC_773/Y INVX1_LOC_75/A 0.16fF
C31038 NOR2X1_LOC_618/a_36_216# INVX1_LOC_62/Y 0.01fF
C31039 NOR2X1_LOC_389/A INVX1_LOC_89/A 0.15fF
C31040 NAND2X1_LOC_786/a_36_24# INVX1_LOC_143/A 0.01fF
C31041 NOR2X1_LOC_160/B INPUT_1 0.21fF
C31042 NOR2X1_LOC_717/B NOR2X1_LOC_717/Y 0.03fF
C31043 NAND2X1_LOC_36/A INVX1_LOC_83/A 1.35fF
C31044 NOR2X1_LOC_644/A NOR2X1_LOC_794/B 0.67fF
C31045 INVX1_LOC_8/A NOR2X1_LOC_709/A 0.17fF
C31046 NAND2X1_LOC_341/A NOR2X1_LOC_759/Y 0.01fF
C31047 INVX1_LOC_88/A NOR2X1_LOC_218/a_36_216# 0.00fF
C31048 INVX1_LOC_1/A NOR2X1_LOC_751/A 0.04fF
C31049 NAND2X1_LOC_350/A INVX1_LOC_28/A 0.98fF
C31050 NOR2X1_LOC_666/Y NOR2X1_LOC_74/A 1.75fF
C31051 NOR2X1_LOC_272/Y INVX1_LOC_98/A 0.10fF
C31052 NAND2X1_LOC_563/Y NAND2X1_LOC_141/A 0.11fF
C31053 INVX1_LOC_208/A INVX1_LOC_49/A 0.03fF
C31054 INVX1_LOC_45/A INVX1_LOC_313/A 0.99fF
C31055 INVX1_LOC_104/A INVX1_LOC_177/A 0.06fF
C31056 NOR2X1_LOC_216/B INVX1_LOC_32/A 0.07fF
C31057 NOR2X1_LOC_67/A INVX1_LOC_34/A 0.26fF
C31058 INPUT_3 NOR2X1_LOC_19/B 0.19fF
C31059 NOR2X1_LOC_750/Y INVX1_LOC_2/Y 0.41fF
C31060 INVX1_LOC_117/A INVX1_LOC_296/A 0.36fF
C31061 NOR2X1_LOC_78/B NAND2X1_LOC_332/Y 0.02fF
C31062 NOR2X1_LOC_772/Y NOR2X1_LOC_773/Y 0.01fF
C31063 INVX1_LOC_21/A NOR2X1_LOC_557/A 0.06fF
C31064 NOR2X1_LOC_272/Y NOR2X1_LOC_78/A 0.03fF
C31065 NOR2X1_LOC_516/B INVX1_LOC_49/A 0.04fF
C31066 INVX1_LOC_284/A INVX1_LOC_63/A 0.07fF
C31067 INVX1_LOC_118/A NOR2X1_LOC_89/Y 0.06fF
C31068 INVX1_LOC_252/Y INVX1_LOC_75/A 0.01fF
C31069 NOR2X1_LOC_441/Y INVX1_LOC_28/A 0.03fF
C31070 NOR2X1_LOC_798/A INVX1_LOC_93/Y 0.07fF
C31071 NOR2X1_LOC_589/A NOR2X1_LOC_433/A 0.18fF
C31072 INVX1_LOC_11/A INVX1_LOC_222/A 0.01fF
C31073 INVX1_LOC_124/Y NAND2X1_LOC_850/A 0.06fF
C31074 NOR2X1_LOC_643/a_36_216# INVX1_LOC_63/A 0.00fF
C31075 INVX1_LOC_13/A NAND2X1_LOC_5/a_36_24# 0.00fF
C31076 NOR2X1_LOC_639/B INVX1_LOC_37/A 0.01fF
C31077 NAND2X1_LOC_181/Y NOR2X1_LOC_315/Y 0.02fF
C31078 NOR2X1_LOC_142/Y INVX1_LOC_16/A 0.15fF
C31079 NOR2X1_LOC_103/Y INVX1_LOC_6/A 0.01fF
C31080 NOR2X1_LOC_598/B NAND2X1_LOC_472/Y 0.10fF
C31081 NOR2X1_LOC_536/A INVX1_LOC_129/A 0.02fF
C31082 INVX1_LOC_233/A NAND2X1_LOC_721/A 0.14fF
C31083 INVX1_LOC_89/A INVX1_LOC_62/Y 0.44fF
C31084 NOR2X1_LOC_13/Y NAND2X1_LOC_660/a_36_24# 0.00fF
C31085 INVX1_LOC_89/A NOR2X1_LOC_596/A 0.06fF
C31086 NOR2X1_LOC_331/B INVX1_LOC_23/A 0.08fF
C31087 INVX1_LOC_13/A NOR2X1_LOC_84/A 0.01fF
C31088 NOR2X1_LOC_151/Y NOR2X1_LOC_717/Y 0.01fF
C31089 NAND2X1_LOC_360/B NAND2X1_LOC_347/a_36_24# 0.02fF
C31090 INVX1_LOC_313/A INVX1_LOC_71/A 0.60fF
C31091 INVX1_LOC_78/A NOR2X1_LOC_841/A 0.01fF
C31092 INVX1_LOC_203/Y INVX1_LOC_135/A 0.03fF
C31093 NOR2X1_LOC_15/Y NOR2X1_LOC_675/A 0.00fF
C31094 INVX1_LOC_2/A INVX1_LOC_208/A 0.30fF
C31095 INVX1_LOC_7/Y VDD 0.21fF
C31096 NOR2X1_LOC_481/A NOR2X1_LOC_355/A 0.17fF
C31097 NOR2X1_LOC_589/A NOR2X1_LOC_52/B 0.10fF
C31098 NAND2X1_LOC_624/B NOR2X1_LOC_536/A 0.02fF
C31099 NOR2X1_LOC_516/B NOR2X1_LOC_818/Y 0.03fF
C31100 GATE_741 VDD 0.33fF
C31101 NOR2X1_LOC_793/Y NOR2X1_LOC_324/A 0.04fF
C31102 NOR2X1_LOC_186/Y NOR2X1_LOC_111/A 0.08fF
C31103 INVX1_LOC_196/A NOR2X1_LOC_325/A 0.01fF
C31104 NOR2X1_LOC_632/Y INVX1_LOC_266/Y 0.05fF
C31105 INVX1_LOC_171/A NOR2X1_LOC_593/Y 0.04fF
C31106 INVX1_LOC_35/A INVX1_LOC_193/A 0.00fF
C31107 NAND2X1_LOC_569/A D_INPUT_0 0.02fF
C31108 INVX1_LOC_136/A NOR2X1_LOC_368/A 0.72fF
C31109 NAND2X1_LOC_803/B NOR2X1_LOC_595/Y 0.02fF
C31110 INVX1_LOC_45/A INVX1_LOC_6/A 0.10fF
C31111 NOR2X1_LOC_331/Y NOR2X1_LOC_45/B 0.01fF
C31112 INVX1_LOC_39/A INVX1_LOC_12/Y 0.03fF
C31113 NOR2X1_LOC_65/B NOR2X1_LOC_841/A 0.10fF
C31114 NOR2X1_LOC_488/Y NAND2X1_LOC_862/A 0.00fF
C31115 NAND2X1_LOC_465/Y NOR2X1_LOC_130/A 0.07fF
C31116 NAND2X1_LOC_660/Y NAND2X1_LOC_661/B 0.14fF
C31117 INVX1_LOC_5/A INVX1_LOC_38/A 0.18fF
C31118 NOR2X1_LOC_92/Y VDD 0.61fF
C31119 NOR2X1_LOC_82/A NOR2X1_LOC_368/Y 0.01fF
C31120 INVX1_LOC_84/A INVX1_LOC_23/Y 0.07fF
C31121 NAND2X1_LOC_222/B INVX1_LOC_20/A 0.01fF
C31122 NAND2X1_LOC_573/Y NOR2X1_LOC_111/A 0.07fF
C31123 NAND2X1_LOC_841/A INVX1_LOC_22/A 0.01fF
C31124 NOR2X1_LOC_218/Y INVX1_LOC_208/A 0.02fF
C31125 NOR2X1_LOC_590/A NOR2X1_LOC_595/Y 0.53fF
C31126 NOR2X1_LOC_383/B NAND2X1_LOC_572/B 0.07fF
C31127 NAND2X1_LOC_553/a_36_24# INVX1_LOC_16/A 0.00fF
C31128 INVX1_LOC_159/A NAND2X1_LOC_662/B 0.01fF
C31129 INVX1_LOC_24/Y VDD 1.64fF
C31130 NOR2X1_LOC_165/Y NAND2X1_LOC_170/A 0.01fF
C31131 NOR2X1_LOC_89/A INVX1_LOC_4/A 1.15fF
C31132 NAND2X1_LOC_444/B INVX1_LOC_29/A 0.01fF
C31133 NOR2X1_LOC_77/a_36_216# INVX1_LOC_4/Y 0.13fF
C31134 INVX1_LOC_208/Y INVX1_LOC_53/Y 1.00fF
C31135 INVX1_LOC_269/A D_INPUT_3 0.15fF
C31136 INVX1_LOC_5/A NOR2X1_LOC_96/Y 0.11fF
C31137 NOR2X1_LOC_216/a_36_216# INVX1_LOC_155/A 0.00fF
C31138 INVX1_LOC_14/A NAND2X1_LOC_633/Y 0.00fF
C31139 NAND2X1_LOC_276/Y NOR2X1_LOC_750/A 0.03fF
C31140 NOR2X1_LOC_334/Y INVX1_LOC_29/A 0.18fF
C31141 INVX1_LOC_11/A INVX1_LOC_20/A 2.40fF
C31142 NOR2X1_LOC_748/a_36_216# INVX1_LOC_22/A 0.00fF
C31143 NAND2X1_LOC_471/Y NAND2X1_LOC_74/B 0.00fF
C31144 INVX1_LOC_269/A INVX1_LOC_14/Y 0.07fF
C31145 NOR2X1_LOC_658/Y INVX1_LOC_159/Y 0.01fF
C31146 INVX1_LOC_90/A NOR2X1_LOC_377/Y 0.00fF
C31147 NOR2X1_LOC_794/B NOR2X1_LOC_540/B 0.00fF
C31148 NOR2X1_LOC_329/B NAND2X1_LOC_833/Y 0.01fF
C31149 INVX1_LOC_232/Y INVX1_LOC_80/A 0.02fF
C31150 INVX1_LOC_28/A NOR2X1_LOC_142/Y 0.10fF
C31151 INVX1_LOC_178/A INVX1_LOC_38/A 0.03fF
C31152 INVX1_LOC_223/A INVX1_LOC_91/A 0.02fF
C31153 NOR2X1_LOC_536/A NOR2X1_LOC_440/B 0.17fF
C31154 INVX1_LOC_57/A NOR2X1_LOC_461/a_36_216# 0.00fF
C31155 INVX1_LOC_299/A INVX1_LOC_117/A 0.03fF
C31156 NOR2X1_LOC_653/B INVX1_LOC_118/A 0.02fF
C31157 NOR2X1_LOC_82/A INVX1_LOC_46/A 0.02fF
C31158 NAND2X1_LOC_508/A NOR2X1_LOC_844/A 0.05fF
C31159 NAND2X1_LOC_568/A NAND2X1_LOC_800/A 0.02fF
C31160 NAND2X1_LOC_67/Y INVX1_LOC_281/A 0.00fF
C31161 NOR2X1_LOC_753/Y INPUT_0 0.07fF
C31162 INVX1_LOC_83/A NAND2X1_LOC_684/a_36_24# 0.07fF
C31163 INVX1_LOC_71/A INVX1_LOC_6/A 2.81fF
C31164 INVX1_LOC_83/A NOR2X1_LOC_731/Y 0.01fF
C31165 NOR2X1_LOC_570/A NOR2X1_LOC_569/Y 0.01fF
C31166 NAND2X1_LOC_364/A NOR2X1_LOC_78/A 0.11fF
C31167 INVX1_LOC_145/Y INVX1_LOC_208/Y 0.00fF
C31168 INVX1_LOC_5/A NAND2X1_LOC_848/Y 0.07fF
C31169 NAND2X1_LOC_340/a_36_24# NAND2X1_LOC_453/A 0.01fF
C31170 INVX1_LOC_41/A NOR2X1_LOC_721/Y 0.02fF
C31171 D_INPUT_0 INVX1_LOC_316/Y 0.11fF
C31172 NOR2X1_LOC_419/Y INVX1_LOC_48/A 0.02fF
C31173 NOR2X1_LOC_593/Y INVX1_LOC_222/A 0.42fF
C31174 INVX1_LOC_90/A NOR2X1_LOC_773/Y 0.10fF
C31175 NOR2X1_LOC_389/B NOR2X1_LOC_773/Y 0.00fF
C31176 NAND2X1_LOC_93/B NOR2X1_LOC_440/B 0.07fF
C31177 NAND2X1_LOC_464/B INVX1_LOC_29/A 0.98fF
C31178 NOR2X1_LOC_662/a_36_216# NOR2X1_LOC_649/B 0.01fF
C31179 NOR2X1_LOC_742/A NOR2X1_LOC_718/a_36_216# 0.01fF
C31180 NAND2X1_LOC_500/Y INVX1_LOC_46/A 0.01fF
C31181 NAND2X1_LOC_201/a_36_24# NAND2X1_LOC_74/B 0.01fF
C31182 NAND2X1_LOC_733/Y NOR2X1_LOC_822/a_36_216# 0.00fF
C31183 NOR2X1_LOC_458/Y INVX1_LOC_206/Y 0.00fF
C31184 NOR2X1_LOC_474/A INVX1_LOC_167/Y 0.08fF
C31185 NOR2X1_LOC_516/B INPUT_1 0.04fF
C31186 INVX1_LOC_47/A INVX1_LOC_22/A 0.03fF
C31187 INVX1_LOC_174/A NOR2X1_LOC_376/Y 0.04fF
C31188 NOR2X1_LOC_816/A INVX1_LOC_38/A 0.11fF
C31189 INVX1_LOC_104/A INVX1_LOC_285/Y 0.10fF
C31190 NAND2X1_LOC_842/B INVX1_LOC_1/Y 0.05fF
C31191 NOR2X1_LOC_754/a_36_216# NOR2X1_LOC_482/Y 0.01fF
C31192 INVX1_LOC_23/Y INVX1_LOC_15/A 0.03fF
C31193 NAND2X1_LOC_359/Y INVX1_LOC_154/Y 0.12fF
C31194 INVX1_LOC_213/A NAND2X1_LOC_782/B 0.04fF
C31195 INVX1_LOC_206/Y INVX1_LOC_121/Y 0.37fF
C31196 NAND2X1_LOC_550/A INVX1_LOC_118/A 0.09fF
C31197 NAND2X1_LOC_95/a_36_24# INVX1_LOC_296/A 0.00fF
C31198 INVX1_LOC_13/A NOR2X1_LOC_112/Y 0.24fF
C31199 NOR2X1_LOC_67/A INPUT_0 0.08fF
C31200 INVX1_LOC_286/A NOR2X1_LOC_84/Y 0.19fF
C31201 INVX1_LOC_103/A INVX1_LOC_92/A 0.25fF
C31202 INVX1_LOC_143/A NOR2X1_LOC_83/Y 0.06fF
C31203 NOR2X1_LOC_160/B INVX1_LOC_118/A 0.01fF
C31204 INVX1_LOC_149/Y INVX1_LOC_91/A 0.02fF
C31205 INVX1_LOC_90/A NAND2X1_LOC_317/a_36_24# 0.00fF
C31206 INVX1_LOC_246/A INVX1_LOC_54/A 0.01fF
C31207 INVX1_LOC_298/Y NOR2X1_LOC_334/Y 0.07fF
C31208 NOR2X1_LOC_433/A INVX1_LOC_147/Y 0.02fF
C31209 INVX1_LOC_206/Y INVX1_LOC_177/A 0.89fF
C31210 INVX1_LOC_161/Y INVX1_LOC_291/A -0.09fF
C31211 INVX1_LOC_49/A NOR2X1_LOC_324/B 0.02fF
C31212 NOR2X1_LOC_357/Y NOR2X1_LOC_303/Y 0.10fF
C31213 INVX1_LOC_64/A NOR2X1_LOC_89/A 1.54fF
C31214 NOR2X1_LOC_433/A INVX1_LOC_20/A 0.03fF
C31215 VDD NAND2X1_LOC_837/Y 1.09fF
C31216 NAND2X1_LOC_85/a_36_24# INVX1_LOC_63/A 0.01fF
C31217 NOR2X1_LOC_445/Y NAND2X1_LOC_447/Y 0.08fF
C31218 NOR2X1_LOC_837/Y INVX1_LOC_37/A 0.01fF
C31219 INVX1_LOC_104/A INVX1_LOC_65/A 0.10fF
C31220 D_INPUT_1 INVX1_LOC_47/Y 0.03fF
C31221 NOR2X1_LOC_632/Y INVX1_LOC_42/Y 0.00fF
C31222 INVX1_LOC_292/A INVX1_LOC_92/A 0.03fF
C31223 NOR2X1_LOC_359/Y NOR2X1_LOC_363/Y 0.03fF
C31224 INVX1_LOC_49/A NAND2X1_LOC_211/Y 0.60fF
C31225 INVX1_LOC_201/Y NAND2X1_LOC_659/B 0.03fF
C31226 INVX1_LOC_151/A INVX1_LOC_147/Y 0.02fF
C31227 INVX1_LOC_279/A INVX1_LOC_75/A 0.17fF
C31228 INPUT_3 NOR2X1_LOC_216/B 0.03fF
C31229 INVX1_LOC_104/A NOR2X1_LOC_137/B 0.07fF
C31230 NAND2X1_LOC_477/A NOR2X1_LOC_56/Y 0.00fF
C31231 NOR2X1_LOC_569/A INVX1_LOC_220/Y 0.01fF
C31232 INVX1_LOC_17/A NAND2X1_LOC_475/Y 0.03fF
C31233 INVX1_LOC_41/A VDD 1.20fF
C31234 INVX1_LOC_34/A NOR2X1_LOC_558/A 0.04fF
C31235 INVX1_LOC_45/A INVX1_LOC_131/Y 0.07fF
C31236 NAND2X1_LOC_348/A NOR2X1_LOC_332/A 0.02fF
C31237 NOR2X1_LOC_730/Y NOR2X1_LOC_728/B 0.11fF
C31238 NAND2X1_LOC_332/Y INVX1_LOC_46/A 0.01fF
C31239 NOR2X1_LOC_498/Y VDD 0.29fF
C31240 NOR2X1_LOC_617/Y NOR2X1_LOC_536/A 0.02fF
C31241 INVX1_LOC_201/Y VDD 0.21fF
C31242 NOR2X1_LOC_392/Y NOR2X1_LOC_38/B 0.05fF
C31243 NOR2X1_LOC_599/A NAND2X1_LOC_802/Y 0.09fF
C31244 NOR2X1_LOC_52/B INVX1_LOC_20/A 0.09fF
C31245 NOR2X1_LOC_384/Y NAND2X1_LOC_243/Y 0.02fF
C31246 INVX1_LOC_90/A INVX1_LOC_140/A 0.07fF
C31247 NAND2X1_LOC_537/Y INVX1_LOC_264/A 0.06fF
C31248 NAND2X1_LOC_703/Y NOR2X1_LOC_669/A 0.04fF
C31249 NAND2X1_LOC_794/B NOR2X1_LOC_48/B 0.89fF
C31250 NOR2X1_LOC_554/B INVX1_LOC_108/A 0.05fF
C31251 INVX1_LOC_144/A NOR2X1_LOC_130/A 0.04fF
C31252 NAND2X1_LOC_564/B NOR2X1_LOC_528/Y 0.01fF
C31253 INVX1_LOC_136/A NOR2X1_LOC_235/Y 0.03fF
C31254 NAND2X1_LOC_839/Y INVX1_LOC_76/A 0.01fF
C31255 NOR2X1_LOC_588/A INVX1_LOC_22/A 0.03fF
C31256 NOR2X1_LOC_78/B INVX1_LOC_59/Y 0.07fF
C31257 INVX1_LOC_25/A INVX1_LOC_16/Y 0.02fF
C31258 NAND2X1_LOC_477/A VDD 1.60fF
C31259 NAND2X1_LOC_662/Y INVX1_LOC_91/A 0.46fF
C31260 NOR2X1_LOC_745/Y NAND2X1_LOC_782/B 0.00fF
C31261 NAND2X1_LOC_39/Y INVX1_LOC_266/Y 0.02fF
C31262 INVX1_LOC_50/A NOR2X1_LOC_727/B 0.03fF
C31263 NOR2X1_LOC_636/B NAND2X1_LOC_651/B 0.05fF
C31264 INVX1_LOC_47/Y NOR2X1_LOC_652/Y 0.01fF
C31265 NAND2X1_LOC_543/a_36_24# INVX1_LOC_84/A 0.00fF
C31266 NOR2X1_LOC_514/A NOR2X1_LOC_649/B 0.05fF
C31267 NOR2X1_LOC_78/B NOR2X1_LOC_300/a_36_216# 0.00fF
C31268 NOR2X1_LOC_249/Y INVX1_LOC_15/A 0.46fF
C31269 INVX1_LOC_2/A NAND2X1_LOC_211/Y 0.04fF
C31270 INVX1_LOC_136/A NOR2X1_LOC_832/a_36_216# 0.12fF
C31271 INVX1_LOC_45/A NOR2X1_LOC_117/Y 0.01fF
C31272 NAND2X1_LOC_787/A NOR2X1_LOC_301/A 0.00fF
C31273 NOR2X1_LOC_398/Y VDD 0.18fF
C31274 NOR2X1_LOC_207/A VDD 0.24fF
C31275 INVX1_LOC_278/Y NOR2X1_LOC_164/Y 0.02fF
C31276 NOR2X1_LOC_123/B INVX1_LOC_6/A 0.07fF
C31277 INVX1_LOC_291/Y INVX1_LOC_16/A 0.01fF
C31278 NOR2X1_LOC_547/B INVX1_LOC_176/A 0.01fF
C31279 NOR2X1_LOC_758/Y NOR2X1_LOC_536/A 0.01fF
C31280 INVX1_LOC_89/A INVX1_LOC_51/Y 0.03fF
C31281 NOR2X1_LOC_533/Y INVX1_LOC_12/A 0.08fF
C31282 NOR2X1_LOC_189/A INVX1_LOC_54/A 0.02fF
C31283 INVX1_LOC_64/Y VDD 0.36fF
C31284 NOR2X1_LOC_561/Y NOR2X1_LOC_45/B 0.19fF
C31285 NOR2X1_LOC_315/Y INVX1_LOC_117/A 0.00fF
C31286 INVX1_LOC_95/Y INVX1_LOC_22/A 0.02fF
C31287 INVX1_LOC_278/A INVX1_LOC_23/Y 0.01fF
C31288 INVX1_LOC_5/A NAND2X1_LOC_223/A 0.03fF
C31289 INVX1_LOC_24/A NOR2X1_LOC_155/A 0.03fF
C31290 NOR2X1_LOC_160/B NAND2X1_LOC_63/Y 0.04fF
C31291 NOR2X1_LOC_589/A INVX1_LOC_199/A 0.03fF
C31292 NOR2X1_LOC_377/Y INVX1_LOC_38/A 0.00fF
C31293 NAND2X1_LOC_115/a_36_24# INVX1_LOC_9/A 0.00fF
C31294 INVX1_LOC_310/A INVX1_LOC_117/A 0.07fF
C31295 INVX1_LOC_25/A NAND2X1_LOC_205/A 0.05fF
C31296 INVX1_LOC_279/Y INVX1_LOC_19/A 0.01fF
C31297 NAND2X1_LOC_563/A D_INPUT_3 0.28fF
C31298 INVX1_LOC_230/Y NAND2X1_LOC_74/B 0.34fF
C31299 INVX1_LOC_278/Y INVX1_LOC_46/A 0.07fF
C31300 NOR2X1_LOC_798/A INVX1_LOC_87/A 0.06fF
C31301 NOR2X1_LOC_218/Y NAND2X1_LOC_211/Y 0.20fF
C31302 NOR2X1_LOC_413/Y NOR2X1_LOC_629/Y 0.00fF
C31303 INVX1_LOC_22/A NOR2X1_LOC_305/Y 0.03fF
C31304 NOR2X1_LOC_542/Y INVX1_LOC_186/A 0.03fF
C31305 VDD NOR2X1_LOC_211/A 0.24fF
C31306 NOR2X1_LOC_360/Y NOR2X1_LOC_814/A 0.17fF
C31307 NOR2X1_LOC_152/Y NOR2X1_LOC_841/A 0.10fF
C31308 INVX1_LOC_71/A NOR2X1_LOC_117/Y 0.03fF
C31309 INVX1_LOC_102/Y INVX1_LOC_6/A 0.03fF
C31310 INVX1_LOC_45/A NOR2X1_LOC_633/A 0.03fF
C31311 NOR2X1_LOC_636/B INVX1_LOC_15/A 0.07fF
C31312 INVX1_LOC_246/A NOR2X1_LOC_48/B 0.10fF
C31313 NOR2X1_LOC_706/Y NOR2X1_LOC_706/A 0.00fF
C31314 NOR2X1_LOC_773/Y NOR2X1_LOC_561/A 0.01fF
C31315 NOR2X1_LOC_590/Y NOR2X1_LOC_727/B 0.01fF
C31316 INVX1_LOC_311/Y INVX1_LOC_186/A 0.07fF
C31317 NOR2X1_LOC_751/A NOR2X1_LOC_548/B 0.03fF
C31318 NOR2X1_LOC_773/Y INVX1_LOC_38/A 0.07fF
C31319 NOR2X1_LOC_309/Y NOR2X1_LOC_79/a_36_216# 0.00fF
C31320 NOR2X1_LOC_99/B NOR2X1_LOC_35/Y 0.10fF
C31321 INVX1_LOC_268/Y INVX1_LOC_117/A 0.01fF
C31322 NOR2X1_LOC_482/Y INVX1_LOC_54/A 0.01fF
C31323 NOR2X1_LOC_214/B NAND2X1_LOC_212/Y 0.02fF
C31324 INVX1_LOC_83/A INVX1_LOC_176/A 0.03fF
C31325 NAND2X1_LOC_562/B NAND2X1_LOC_848/Y 0.08fF
C31326 NAND2X1_LOC_842/B INVX1_LOC_93/Y 0.08fF
C31327 NAND2X1_LOC_848/A INVX1_LOC_316/Y 0.00fF
C31328 NAND2X1_LOC_500/a_36_24# INVX1_LOC_118/A 0.00fF
C31329 INVX1_LOC_36/A NOR2X1_LOC_226/Y 0.00fF
C31330 NOR2X1_LOC_596/Y INVX1_LOC_15/A 0.01fF
C31331 NOR2X1_LOC_299/Y VDD 0.64fF
C31332 INVX1_LOC_306/A INVX1_LOC_46/A 0.23fF
C31333 NOR2X1_LOC_523/B INVX1_LOC_29/A 0.08fF
C31334 INVX1_LOC_89/A NAND2X1_LOC_414/a_36_24# 0.00fF
C31335 INVX1_LOC_21/A INVX1_LOC_271/A 0.07fF
C31336 NOR2X1_LOC_6/B NAND2X1_LOC_141/Y 0.08fF
C31337 NOR2X1_LOC_703/B INVX1_LOC_290/Y 0.00fF
C31338 NAND2X1_LOC_705/a_36_24# INVX1_LOC_118/A 0.00fF
C31339 INVX1_LOC_298/A INVX1_LOC_295/Y 0.00fF
C31340 NOR2X1_LOC_792/B INVX1_LOC_285/A 0.01fF
C31341 INVX1_LOC_108/Y NOR2X1_LOC_846/A 0.01fF
C31342 INVX1_LOC_182/A NOR2X1_LOC_35/Y 0.10fF
C31343 NOR2X1_LOC_45/B NOR2X1_LOC_167/Y 0.03fF
C31344 INVX1_LOC_290/A INVX1_LOC_54/A 0.05fF
C31345 NOR2X1_LOC_122/Y VDD 0.12fF
C31346 NAND2X1_LOC_319/a_36_24# NOR2X1_LOC_510/B 0.00fF
C31347 NAND2X1_LOC_850/A NOR2X1_LOC_266/B 0.39fF
C31348 INVX1_LOC_58/A INVX1_LOC_299/A 0.27fF
C31349 INVX1_LOC_13/A NOR2X1_LOC_78/Y 0.03fF
C31350 NOR2X1_LOC_189/A NOR2X1_LOC_48/B 0.08fF
C31351 INVX1_LOC_25/A NOR2X1_LOC_817/Y 0.06fF
C31352 NOR2X1_LOC_537/Y INVX1_LOC_63/A 0.10fF
C31353 INVX1_LOC_247/Y NOR2X1_LOC_334/Y 0.02fF
C31354 NOR2X1_LOC_78/A NOR2X1_LOC_349/A 0.12fF
C31355 NAND2X1_LOC_338/B INVX1_LOC_63/A 0.11fF
C31356 NOR2X1_LOC_272/Y NOR2X1_LOC_186/Y 0.10fF
C31357 INVX1_LOC_103/A INVX1_LOC_53/A 0.11fF
C31358 INVX1_LOC_30/A NOR2X1_LOC_301/A 0.06fF
C31359 NOR2X1_LOC_303/Y INVX1_LOC_32/A 0.07fF
C31360 INVX1_LOC_17/A NAND2X1_LOC_787/A 0.05fF
C31361 NOR2X1_LOC_78/A NOR2X1_LOC_113/A 0.06fF
C31362 NOR2X1_LOC_78/A NOR2X1_LOC_405/A 0.09fF
C31363 INVX1_LOC_17/A NAND2X1_LOC_363/B 0.07fF
C31364 NAND2X1_LOC_662/B VDD 0.03fF
C31365 INVX1_LOC_21/A INVX1_LOC_27/A 0.40fF
C31366 NAND2X1_LOC_9/Y NOR2X1_LOC_82/A 0.10fF
C31367 NOR2X1_LOC_739/a_36_216# NOR2X1_LOC_155/A 0.00fF
C31368 INVX1_LOC_64/A INVX1_LOC_224/A 0.03fF
C31369 INVX1_LOC_21/A NOR2X1_LOC_824/A 0.05fF
C31370 INVX1_LOC_45/A INVX1_LOC_28/Y 0.01fF
C31371 INVX1_LOC_10/A NOR2X1_LOC_831/B 0.07fF
C31372 INVX1_LOC_232/A INVX1_LOC_84/A 0.10fF
C31373 NOR2X1_LOC_392/B INVX1_LOC_42/A 0.00fF
C31374 NOR2X1_LOC_67/A NOR2X1_LOC_84/B 0.00fF
C31375 INVX1_LOC_233/A NOR2X1_LOC_82/A 0.10fF
C31376 INVX1_LOC_140/A INVX1_LOC_38/A 1.30fF
C31377 INVX1_LOC_64/A INVX1_LOC_11/A 0.19fF
C31378 NOR2X1_LOC_510/Y NOR2X1_LOC_92/Y 0.09fF
C31379 NAND2X1_LOC_841/A INVX1_LOC_186/Y 0.00fF
C31380 INVX1_LOC_124/Y INVX1_LOC_57/A 0.03fF
C31381 INVX1_LOC_45/A INVX1_LOC_270/A 0.03fF
C31382 NOR2X1_LOC_658/Y INVX1_LOC_50/A 0.09fF
C31383 INVX1_LOC_292/A INVX1_LOC_53/A 0.47fF
C31384 NAND2X1_LOC_564/B NAND2X1_LOC_477/Y 0.00fF
C31385 NAND2X1_LOC_319/A NOR2X1_LOC_697/Y 0.01fF
C31386 NOR2X1_LOC_593/Y INVX1_LOC_4/A 0.13fF
C31387 INVX1_LOC_224/Y INVX1_LOC_36/A 0.10fF
C31388 NOR2X1_LOC_45/B INVX1_LOC_76/A 0.32fF
C31389 NOR2X1_LOC_802/A NOR2X1_LOC_640/B 0.03fF
C31390 NAND2X1_LOC_472/a_36_24# INVX1_LOC_274/A 0.00fF
C31391 INVX1_LOC_13/A NOR2X1_LOC_721/B 0.01fF
C31392 NAND2X1_LOC_850/Y NOR2X1_LOC_89/A 0.07fF
C31393 NOR2X1_LOC_78/A NOR2X1_LOC_857/A 0.07fF
C31394 INVX1_LOC_126/A NAND2X1_LOC_642/Y 0.04fF
C31395 NAND2X1_LOC_634/Y NAND2X1_LOC_464/B 0.07fF
C31396 NAND2X1_LOC_231/Y NAND2X1_LOC_807/a_36_24# 0.06fF
C31397 INVX1_LOC_50/A NOR2X1_LOC_518/Y 0.07fF
C31398 NAND2X1_LOC_116/A INVX1_LOC_15/A 0.10fF
C31399 INVX1_LOC_140/A NOR2X1_LOC_51/A 0.33fF
C31400 NAND2X1_LOC_354/Y INVX1_LOC_271/A 0.19fF
C31401 NOR2X1_LOC_806/Y NOR2X1_LOC_812/A 0.56fF
C31402 NOR2X1_LOC_172/Y INVX1_LOC_78/A 0.71fF
C31403 NOR2X1_LOC_632/Y INVX1_LOC_19/A 0.00fF
C31404 NOR2X1_LOC_609/A NOR2X1_LOC_383/B 0.01fF
C31405 NOR2X1_LOC_483/B INVX1_LOC_5/A 0.04fF
C31406 NOR2X1_LOC_798/A INVX1_LOC_134/A 0.04fF
C31407 INVX1_LOC_56/Y INVX1_LOC_12/A 0.03fF
C31408 INVX1_LOC_71/A INVX1_LOC_28/Y 0.01fF
C31409 INVX1_LOC_6/A NOR2X1_LOC_331/B 0.18fF
C31410 NOR2X1_LOC_92/Y NOR2X1_LOC_361/B 0.07fF
C31411 INVX1_LOC_54/Y INVX1_LOC_32/A 2.69fF
C31412 NOR2X1_LOC_74/A INVX1_LOC_274/A 0.10fF
C31413 INVX1_LOC_104/A INVX1_LOC_4/Y 0.07fF
C31414 NAND2X1_LOC_800/A NAND2X1_LOC_648/a_36_24# 0.00fF
C31415 NOR2X1_LOC_569/Y INVX1_LOC_29/A 0.01fF
C31416 INVX1_LOC_50/A NOR2X1_LOC_13/Y 0.00fF
C31417 D_INPUT_0 NOR2X1_LOC_662/A 0.03fF
C31418 NOR2X1_LOC_111/A NAND2X1_LOC_642/Y 0.07fF
C31419 INVX1_LOC_71/A INVX1_LOC_270/A 0.10fF
C31420 INVX1_LOC_39/A NOR2X1_LOC_160/B 0.03fF
C31421 INVX1_LOC_45/A NOR2X1_LOC_109/Y 0.03fF
C31422 INVX1_LOC_13/A NOR2X1_LOC_610/Y 0.05fF
C31423 NOR2X1_LOC_195/A NAND2X1_LOC_473/A 0.03fF
C31424 NOR2X1_LOC_52/a_36_216# NAND2X1_LOC_469/B 0.00fF
C31425 NAND2X1_LOC_464/Y INVX1_LOC_23/Y 0.01fF
C31426 NOR2X1_LOC_817/Y INVX1_LOC_1/A 0.43fF
C31427 NOR2X1_LOC_65/B NOR2X1_LOC_172/Y 0.03fF
C31428 INVX1_LOC_224/Y NOR2X1_LOC_237/Y 0.50fF
C31429 INVX1_LOC_313/Y INVX1_LOC_63/A 0.07fF
C31430 NOR2X1_LOC_716/B NOR2X1_LOC_383/B 0.07fF
C31431 NOR2X1_LOC_65/B NOR2X1_LOC_772/Y 0.01fF
C31432 NOR2X1_LOC_598/B INVX1_LOC_24/A 0.15fF
C31433 INVX1_LOC_290/A NOR2X1_LOC_48/B 0.05fF
C31434 NOR2X1_LOC_391/Y NOR2X1_LOC_99/Y -0.00fF
C31435 INVX1_LOC_83/A NOR2X1_LOC_340/A 0.26fF
C31436 NOR2X1_LOC_68/A INVX1_LOC_213/A 0.03fF
C31437 INVX1_LOC_135/A NOR2X1_LOC_664/a_36_216# 0.01fF
C31438 NOR2X1_LOC_658/Y NOR2X1_LOC_206/a_36_216# 0.01fF
C31439 NOR2X1_LOC_788/B INVX1_LOC_19/A 0.00fF
C31440 D_INPUT_3 NOR2X1_LOC_37/a_36_216# 0.00fF
C31441 NOR2X1_LOC_65/B NOR2X1_LOC_392/B 0.03fF
C31442 NOR2X1_LOC_567/B NOR2X1_LOC_814/A 0.07fF
C31443 NAND2X1_LOC_814/a_36_24# NAND2X1_LOC_798/B 0.00fF
C31444 NAND2X1_LOC_725/A INVX1_LOC_24/A 0.04fF
C31445 INVX1_LOC_6/A NOR2X1_LOC_592/B 0.02fF
C31446 INVX1_LOC_25/Y NOR2X1_LOC_38/B 0.90fF
C31447 NOR2X1_LOC_186/Y NAND2X1_LOC_364/A 0.51fF
C31448 NAND2X1_LOC_53/Y D_GATE_741 0.02fF
C31449 NOR2X1_LOC_828/Y INVX1_LOC_33/A 0.07fF
C31450 NOR2X1_LOC_388/Y INVX1_LOC_23/A 0.07fF
C31451 INVX1_LOC_281/A INVX1_LOC_76/A 1.87fF
C31452 NOR2X1_LOC_683/Y NOR2X1_LOC_684/Y 0.03fF
C31453 INVX1_LOC_71/A NOR2X1_LOC_109/Y 0.03fF
C31454 INVX1_LOC_67/A INVX1_LOC_53/A 0.03fF
C31455 NOR2X1_LOC_324/A NOR2X1_LOC_729/A 0.03fF
C31456 INVX1_LOC_11/A INVX1_LOC_43/Y 0.03fF
C31457 INVX1_LOC_64/A NOR2X1_LOC_433/A 0.10fF
C31458 NOR2X1_LOC_334/A NOR2X1_LOC_461/B 0.01fF
C31459 NOR2X1_LOC_848/Y INVX1_LOC_31/A 1.03fF
C31460 INVX1_LOC_22/A INVX1_LOC_271/Y 0.07fF
C31461 NOR2X1_LOC_355/a_36_216# INVX1_LOC_42/A 0.01fF
C31462 INVX1_LOC_64/A NOR2X1_LOC_593/Y 0.03fF
C31463 INVX1_LOC_90/A INVX1_LOC_42/A 0.35fF
C31464 INVX1_LOC_50/A NOR2X1_LOC_504/Y 0.17fF
C31465 NOR2X1_LOC_763/Y D_INPUT_5 0.00fF
C31466 NAND2X1_LOC_350/A INVX1_LOC_246/A 0.10fF
C31467 INVX1_LOC_58/A NOR2X1_LOC_315/Y 0.10fF
C31468 NOR2X1_LOC_84/Y NAND2X1_LOC_215/A 0.09fF
C31469 NOR2X1_LOC_175/A NOR2X1_LOC_748/A 0.41fF
C31470 NAND2X1_LOC_181/Y NAND2X1_LOC_99/A 0.00fF
C31471 NOR2X1_LOC_389/B INVX1_LOC_42/A 0.42fF
C31472 INVX1_LOC_303/A INVX1_LOC_50/Y 0.10fF
C31473 INVX1_LOC_108/Y NAND2X1_LOC_116/A 0.08fF
C31474 NOR2X1_LOC_218/a_36_216# INVX1_LOC_272/A 0.00fF
C31475 NOR2X1_LOC_385/Y INVX1_LOC_12/A 0.09fF
C31476 INVX1_LOC_17/A INVX1_LOC_30/A 1.45fF
C31477 NOR2X1_LOC_309/Y NAND2X1_LOC_793/B 0.01fF
C31478 INVX1_LOC_5/A INVX1_LOC_33/A 0.06fF
C31479 NAND2X1_LOC_480/a_36_24# INVX1_LOC_78/A 0.00fF
C31480 INVX1_LOC_89/A INVX1_LOC_251/A 0.02fF
C31481 NAND2X1_LOC_624/A INVX1_LOC_3/Y 0.05fF
C31482 INVX1_LOC_58/A NOR2X1_LOC_432/Y 0.02fF
C31483 INVX1_LOC_36/A NOR2X1_LOC_103/Y 0.14fF
C31484 NOR2X1_LOC_647/a_36_216# INVX1_LOC_31/A 0.01fF
C31485 NOR2X1_LOC_61/B NOR2X1_LOC_860/B 0.03fF
C31486 INVX1_LOC_64/A NOR2X1_LOC_52/B 0.25fF
C31487 NOR2X1_LOC_598/B INVX1_LOC_143/A 0.17fF
C31488 NOR2X1_LOC_448/B NOR2X1_LOC_596/A 0.05fF
C31489 NOR2X1_LOC_332/A NAND2X1_LOC_223/A 0.07fF
C31490 NOR2X1_LOC_366/B INVX1_LOC_23/A 0.05fF
C31491 NAND2X1_LOC_140/A NOR2X1_LOC_334/Y 0.03fF
C31492 NAND2X1_LOC_348/A INVX1_LOC_42/A 0.01fF
C31493 NOR2X1_LOC_205/Y NOR2X1_LOC_215/Y 0.04fF
C31494 NOR2X1_LOC_808/A INVX1_LOC_292/Y 0.16fF
C31495 NOR2X1_LOC_68/A NOR2X1_LOC_745/Y 0.04fF
C31496 INVX1_LOC_230/Y INVX1_LOC_136/A 0.01fF
C31497 NOR2X1_LOC_435/B NOR2X1_LOC_56/Y 0.03fF
C31498 INPUT_0 NAND2X1_LOC_807/a_36_24# 0.01fF
C31499 NOR2X1_LOC_272/Y INVX1_LOC_225/A 0.10fF
C31500 NAND2X1_LOC_35/B NAND2X1_LOC_35/Y 0.01fF
C31501 NOR2X1_LOC_598/B INVX1_LOC_68/Y 0.03fF
C31502 INVX1_LOC_90/A INVX1_LOC_78/A 0.31fF
C31503 NOR2X1_LOC_510/Y NAND2X1_LOC_477/A 0.07fF
C31504 NOR2X1_LOC_790/B NOR2X1_LOC_500/Y 0.03fF
C31505 INVX1_LOC_233/A INVX1_LOC_278/Y 0.01fF
C31506 INVX1_LOC_127/A NOR2X1_LOC_271/Y 0.07fF
C31507 NOR2X1_LOC_91/A INVX1_LOC_135/A 0.01fF
C31508 INVX1_LOC_45/A INVX1_LOC_36/A 3.95fF
C31509 NOR2X1_LOC_389/B INVX1_LOC_78/A 0.12fF
C31510 NOR2X1_LOC_590/A NOR2X1_LOC_360/Y 0.06fF
C31511 NAND2X1_LOC_218/B INVX1_LOC_252/Y 0.02fF
C31512 NOR2X1_LOC_201/A INVX1_LOC_135/A 0.00fF
C31513 NOR2X1_LOC_658/Y NOR2X1_LOC_659/a_36_216# 0.02fF
C31514 NOR2X1_LOC_237/Y NOR2X1_LOC_103/Y 0.03fF
C31515 INVX1_LOC_21/A INVX1_LOC_206/A 0.02fF
C31516 NOR2X1_LOC_717/B NOR2X1_LOC_383/B 0.06fF
C31517 NOR2X1_LOC_246/A NAND2X1_LOC_286/B 0.13fF
C31518 INVX1_LOC_75/A NOR2X1_LOC_38/B 0.06fF
C31519 VDD NAND2X1_LOC_574/A 3.16fF
C31520 NAND2X1_LOC_39/a_36_24# INVX1_LOC_72/A 0.01fF
C31521 INVX1_LOC_41/A NOR2X1_LOC_361/B 0.17fF
C31522 VDD NOR2X1_LOC_435/B -0.00fF
C31523 INVX1_LOC_40/Y NOR2X1_LOC_820/A 0.00fF
C31524 NOR2X1_LOC_690/A NOR2X1_LOC_232/Y 0.18fF
C31525 INVX1_LOC_5/A INVX1_LOC_40/A 0.09fF
C31526 INVX1_LOC_87/Y INVX1_LOC_26/A 0.02fF
C31527 INVX1_LOC_269/A NOR2X1_LOC_413/Y 0.25fF
C31528 D_INPUT_0 INVX1_LOC_57/A 0.31fF
C31529 NOR2X1_LOC_78/A INVX1_LOC_109/Y 0.01fF
C31530 NOR2X1_LOC_65/B INVX1_LOC_90/A 0.26fF
C31531 NAND2X1_LOC_9/Y NOR2X1_LOC_236/a_36_216# 0.00fF
C31532 NOR2X1_LOC_68/A INVX1_LOC_110/A 0.01fF
C31533 VDD INVX1_LOC_136/Y 0.09fF
C31534 INPUT_1 NAND2X1_LOC_442/a_36_24# 0.01fF
C31535 INVX1_LOC_135/A INVX1_LOC_23/A 0.05fF
C31536 NAND2X1_LOC_721/A INVX1_LOC_119/Y 0.02fF
C31537 NAND2X1_LOC_337/B INVX1_LOC_33/A 0.01fF
C31538 NOR2X1_LOC_65/B NOR2X1_LOC_389/B 0.07fF
C31539 INVX1_LOC_178/A NAND2X1_LOC_798/A 0.08fF
C31540 NOR2X1_LOC_205/Y INVX1_LOC_104/A 0.05fF
C31541 NAND2X1_LOC_337/B NOR2X1_LOC_743/a_36_216# 0.01fF
C31542 INVX1_LOC_45/A INVX1_LOC_145/A 0.01fF
C31543 NAND2X1_LOC_9/Y INVX1_LOC_306/A 0.02fF
C31544 INVX1_LOC_24/Y INVX1_LOC_177/A 0.12fF
C31545 INPUT_3 NAND2X1_LOC_5/a_36_24# 0.01fF
C31546 NOR2X1_LOC_389/a_36_216# INVX1_LOC_57/A 0.00fF
C31547 NOR2X1_LOC_561/Y NOR2X1_LOC_53/Y 0.05fF
C31548 NAND2X1_LOC_537/Y INVX1_LOC_236/A 0.44fF
C31549 INVX1_LOC_36/A INVX1_LOC_71/A 0.35fF
C31550 NOR2X1_LOC_624/A NOR2X1_LOC_160/B 0.01fF
C31551 NOR2X1_LOC_92/Y INVX1_LOC_280/Y 0.09fF
C31552 INVX1_LOC_269/A NAND2X1_LOC_675/a_36_24# 0.02fF
C31553 INVX1_LOC_186/A INVX1_LOC_15/A 0.11fF
C31554 NAND2X1_LOC_569/A NOR2X1_LOC_134/Y 0.02fF
C31555 INVX1_LOC_13/Y INVX1_LOC_30/Y 0.24fF
C31556 INPUT_3 NOR2X1_LOC_84/A 0.03fF
C31557 NAND2X1_LOC_860/A NAND2X1_LOC_551/A 0.03fF
C31558 NAND2X1_LOC_725/A NAND2X1_LOC_800/Y 0.03fF
C31559 INVX1_LOC_223/Y NOR2X1_LOC_548/Y 0.02fF
C31560 INVX1_LOC_304/A INVX1_LOC_170/Y 0.01fF
C31561 INVX1_LOC_35/A NOR2X1_LOC_76/A 0.07fF
C31562 INVX1_LOC_45/A NOR2X1_LOC_804/B 0.07fF
C31563 NOR2X1_LOC_703/B INVX1_LOC_77/A 0.05fF
C31564 INVX1_LOC_43/Y NOR2X1_LOC_52/B 0.32fF
C31565 INVX1_LOC_57/Y NOR2X1_LOC_716/B 0.10fF
C31566 INVX1_LOC_103/A NOR2X1_LOC_78/B 0.08fF
C31567 NOR2X1_LOC_151/Y NOR2X1_LOC_383/B 0.06fF
C31568 NOR2X1_LOC_590/A NOR2X1_LOC_792/B 0.00fF
C31569 NAND2X1_LOC_848/A NOR2X1_LOC_662/A 3.40fF
C31570 NAND2X1_LOC_254/Y INVX1_LOC_20/A 2.05fF
C31571 NOR2X1_LOC_468/Y INVX1_LOC_25/Y 2.74fF
C31572 INVX1_LOC_291/A NOR2X1_LOC_841/A 0.10fF
C31573 NAND2X1_LOC_773/Y INVX1_LOC_22/A 0.45fF
C31574 NAND2X1_LOC_579/A INVX1_LOC_16/A 0.10fF
C31575 NOR2X1_LOC_433/A INVX1_LOC_130/Y 0.03fF
C31576 NOR2X1_LOC_188/A NOR2X1_LOC_39/Y 0.12fF
C31577 INVX1_LOC_21/A INVX1_LOC_234/A 0.07fF
C31578 NOR2X1_LOC_440/Y NOR2X1_LOC_440/B 0.04fF
C31579 NOR2X1_LOC_155/A NOR2X1_LOC_197/B 0.03fF
C31580 INVX1_LOC_145/A INVX1_LOC_71/A 0.01fF
C31581 VDD INVX1_LOC_168/Y 0.21fF
C31582 INVX1_LOC_263/A NOR2X1_LOC_205/Y 0.33fF
C31583 NOR2X1_LOC_208/Y INVX1_LOC_71/A 0.03fF
C31584 NAND2X1_LOC_726/a_36_24# NAND2X1_LOC_811/Y 0.00fF
C31585 NAND2X1_LOC_721/A INVX1_LOC_284/A 0.03fF
C31586 INVX1_LOC_45/A NOR2X1_LOC_309/Y 0.03fF
C31587 INPUT_0 NAND2X1_LOC_787/Y 0.08fF
C31588 INVX1_LOC_172/A NOR2X1_LOC_238/Y 0.03fF
C31589 NOR2X1_LOC_13/Y INVX1_LOC_105/A 0.03fF
C31590 NAND2X1_LOC_741/Y NOR2X1_LOC_576/B 0.03fF
C31591 NAND2X1_LOC_655/A INVX1_LOC_273/A 0.08fF
C31592 NOR2X1_LOC_219/a_36_216# NOR2X1_LOC_759/Y 0.00fF
C31593 NAND2X1_LOC_800/a_36_24# INVX1_LOC_231/A 0.00fF
C31594 NOR2X1_LOC_309/Y NOR2X1_LOC_568/A 0.04fF
C31595 NOR2X1_LOC_78/B INVX1_LOC_292/A 0.07fF
C31596 NOR2X1_LOC_92/Y NAND2X1_LOC_573/A 0.19fF
C31597 D_INPUT_3 NOR2X1_LOC_554/A 0.01fF
C31598 INVX1_LOC_185/A NOR2X1_LOC_661/A 0.64fF
C31599 NOR2X1_LOC_242/A INVX1_LOC_120/A 0.34fF
C31600 INVX1_LOC_35/A INVX1_LOC_73/A 0.03fF
C31601 INVX1_LOC_225/A NAND2X1_LOC_364/A 0.20fF
C31602 INVX1_LOC_152/Y NAND2X1_LOC_348/A 0.02fF
C31603 INVX1_LOC_34/A INVX1_LOC_181/Y 0.04fF
C31604 INVX1_LOC_280/A NOR2X1_LOC_664/a_36_216# 0.00fF
C31605 NOR2X1_LOC_739/Y NOR2X1_LOC_730/Y 0.04fF
C31606 NOR2X1_LOC_574/A INVX1_LOC_18/A 0.04fF
C31607 INVX1_LOC_48/Y NOR2X1_LOC_99/B 0.01fF
C31608 NAND2X1_LOC_30/Y NOR2X1_LOC_764/a_36_216# 0.00fF
C31609 NOR2X1_LOC_531/a_36_216# INVX1_LOC_104/A 0.00fF
C31610 NOR2X1_LOC_45/B NOR2X1_LOC_447/A 0.58fF
C31611 NAND2X1_LOC_849/B INVX1_LOC_42/A 0.14fF
C31612 NOR2X1_LOC_172/Y NOR2X1_LOC_152/Y 0.02fF
C31613 INVX1_LOC_25/A INVX1_LOC_286/A 0.07fF
C31614 INVX1_LOC_207/Y INVX1_LOC_242/A 0.52fF
C31615 NAND2X1_LOC_637/Y INVX1_LOC_29/A 0.01fF
C31616 NOR2X1_LOC_794/A INVX1_LOC_23/A 0.00fF
C31617 INVX1_LOC_49/A INVX1_LOC_155/A 0.05fF
C31618 INVX1_LOC_38/A INVX1_LOC_42/A 7.76fF
C31619 INVX1_LOC_35/Y NAND2X1_LOC_489/Y 0.14fF
C31620 INVX1_LOC_21/A NOR2X1_LOC_19/B 0.07fF
C31621 INVX1_LOC_103/A INVX1_LOC_83/A 0.10fF
C31622 NOR2X1_LOC_309/Y INVX1_LOC_71/A 0.11fF
C31623 INVX1_LOC_303/A NOR2X1_LOC_6/B 0.10fF
C31624 NAND2X1_LOC_522/a_36_24# INVX1_LOC_120/A 0.00fF
C31625 NOR2X1_LOC_67/A INVX1_LOC_72/Y 0.06fF
C31626 NAND2X1_LOC_699/a_36_24# INVX1_LOC_4/A 0.01fF
C31627 NAND2X1_LOC_579/A INVX1_LOC_28/A 0.10fF
C31628 NOR2X1_LOC_552/A INVX1_LOC_23/A 0.25fF
C31629 INVX1_LOC_18/A NAND2X1_LOC_841/A 0.03fF
C31630 NAND2X1_LOC_175/B NAND2X1_LOC_174/a_36_24# 0.01fF
C31631 NOR2X1_LOC_431/a_36_216# NOR2X1_LOC_226/A 0.00fF
C31632 INVX1_LOC_72/A INVX1_LOC_1/Y 0.07fF
C31633 NOR2X1_LOC_9/Y INVX1_LOC_306/Y 0.03fF
C31634 INVX1_LOC_12/A NOR2X1_LOC_831/B 0.95fF
C31635 INVX1_LOC_81/Y INVX1_LOC_10/A 0.01fF
C31636 INVX1_LOC_280/Y NAND2X1_LOC_837/Y 0.07fF
C31637 INVX1_LOC_268/A INVX1_LOC_18/A 0.02fF
C31638 INVX1_LOC_223/A NOR2X1_LOC_553/B 0.00fF
C31639 INVX1_LOC_90/A NOR2X1_LOC_503/Y 0.03fF
C31640 INVX1_LOC_135/A INVX1_LOC_31/A 0.46fF
C31641 INVX1_LOC_27/A INVX1_LOC_311/A 0.04fF
C31642 NOR2X1_LOC_468/Y INVX1_LOC_75/A 0.07fF
C31643 INVX1_LOC_298/Y NAND2X1_LOC_472/Y 0.07fF
C31644 INVX1_LOC_41/A INVX1_LOC_177/A 0.03fF
C31645 INVX1_LOC_195/A NAND2X1_LOC_462/B 0.06fF
C31646 NOR2X1_LOC_433/A NAND2X1_LOC_850/Y 0.01fF
C31647 NOR2X1_LOC_334/Y INVX1_LOC_118/Y 1.30fF
C31648 NOR2X1_LOC_52/Y NOR2X1_LOC_561/Y 0.03fF
C31649 INVX1_LOC_78/A INVX1_LOC_38/A 8.20fF
C31650 NOR2X1_LOC_456/Y NAND2X1_LOC_602/a_36_24# 0.01fF
C31651 NAND2X1_LOC_190/Y INVX1_LOC_75/A 0.02fF
C31652 NOR2X1_LOC_266/B INVX1_LOC_57/A 0.03fF
C31653 NOR2X1_LOC_78/Y INVX1_LOC_32/A 0.03fF
C31654 INVX1_LOC_117/A NAND2X1_LOC_99/A 0.02fF
C31655 INVX1_LOC_64/A INVX1_LOC_199/A 0.02fF
C31656 NOR2X1_LOC_135/Y INVX1_LOC_161/Y 0.01fF
C31657 NOR2X1_LOC_455/a_36_216# INVX1_LOC_177/A 0.00fF
C31658 NOR2X1_LOC_78/B INVX1_LOC_67/A 0.03fF
C31659 NOR2X1_LOC_669/A INVX1_LOC_119/Y 0.07fF
C31660 INVX1_LOC_53/A INVX1_LOC_143/Y 0.13fF
C31661 NOR2X1_LOC_91/A NOR2X1_LOC_813/Y 0.03fF
C31662 INVX1_LOC_49/A NAND2X1_LOC_452/a_36_24# 0.01fF
C31663 INVX1_LOC_37/A NOR2X1_LOC_858/A 0.02fF
C31664 INVX1_LOC_200/Y INVX1_LOC_37/A 0.03fF
C31665 INVX1_LOC_193/Y INVX1_LOC_198/A 0.11fF
C31666 INVX1_LOC_36/A NOR2X1_LOC_123/B 0.33fF
C31667 INVX1_LOC_227/A NOR2X1_LOC_360/Y 0.10fF
C31668 NOR2X1_LOC_773/Y INVX1_LOC_33/A 0.07fF
C31669 NOR2X1_LOC_75/Y NOR2X1_LOC_163/Y 0.02fF
C31670 NAND2X1_LOC_9/Y INVX1_LOC_176/A 1.42fF
C31671 NOR2X1_LOC_498/Y INVX1_LOC_280/Y 0.07fF
C31672 NOR2X1_LOC_229/Y INVX1_LOC_49/A 0.46fF
C31673 NOR2X1_LOC_186/Y NOR2X1_LOC_113/A 0.00fF
C31674 NOR2X1_LOC_616/Y NOR2X1_LOC_413/Y 0.01fF
C31675 INVX1_LOC_53/A NOR2X1_LOC_137/Y 0.14fF
C31676 INVX1_LOC_5/A NOR2X1_LOC_486/Y 0.09fF
C31677 NOR2X1_LOC_186/Y NOR2X1_LOC_405/A 0.10fF
C31678 NOR2X1_LOC_589/A INVX1_LOC_314/Y 0.01fF
C31679 NOR2X1_LOC_51/A INVX1_LOC_78/A 0.47fF
C31680 NOR2X1_LOC_168/B NOR2X1_LOC_802/A 0.34fF
C31681 INVX1_LOC_1/A INVX1_LOC_286/A 0.10fF
C31682 NOR2X1_LOC_91/A INVX1_LOC_280/A 0.03fF
C31683 INVX1_LOC_85/A NOR2X1_LOC_352/Y 0.01fF
C31684 INVX1_LOC_13/Y NOR2X1_LOC_124/A 0.02fF
C31685 NOR2X1_LOC_201/A INVX1_LOC_280/A 0.01fF
C31686 NOR2X1_LOC_65/B INVX1_LOC_38/A 0.21fF
C31687 NOR2X1_LOC_590/A NOR2X1_LOC_567/B 0.08fF
C31688 NOR2X1_LOC_272/Y NAND2X1_LOC_642/Y 0.03fF
C31689 NOR2X1_LOC_454/Y INVX1_LOC_91/A 0.17fF
C31690 NOR2X1_LOC_813/Y INVX1_LOC_23/A 0.07fF
C31691 NAND2X1_LOC_733/Y NOR2X1_LOC_385/Y 0.08fF
C31692 NOR2X1_LOC_52/B NAND2X1_LOC_850/Y 0.07fF
C31693 NOR2X1_LOC_536/A INVX1_LOC_270/Y 0.01fF
C31694 NOR2X1_LOC_389/A INVX1_LOC_75/A 0.10fF
C31695 NAND2X1_LOC_848/A INVX1_LOC_57/A 0.03fF
C31696 NOR2X1_LOC_331/B INVX1_LOC_270/A 0.10fF
C31697 INVX1_LOC_277/A NOR2X1_LOC_828/B 0.05fF
C31698 INVX1_LOC_49/A INVX1_LOC_160/Y 0.06fF
C31699 NOR2X1_LOC_249/a_36_216# INVX1_LOC_75/A 0.00fF
C31700 NAND2X1_LOC_736/Y NAND2X1_LOC_863/B 0.04fF
C31701 NOR2X1_LOC_171/Y INVX1_LOC_30/A 0.04fF
C31702 NAND2X1_LOC_573/Y NOR2X1_LOC_405/A 0.03fF
C31703 NAND2X1_LOC_35/Y VDD 2.22fF
C31704 NOR2X1_LOC_478/a_36_216# INVX1_LOC_113/Y 0.00fF
C31705 INVX1_LOC_155/Y NOR2X1_LOC_665/A 0.06fF
C31706 NOR2X1_LOC_720/B NOR2X1_LOC_619/A 0.00fF
C31707 INVX1_LOC_23/A INVX1_LOC_280/A 0.09fF
C31708 NOR2X1_LOC_383/B NOR2X1_LOC_209/B 0.43fF
C31709 NOR2X1_LOC_639/B INVX1_LOC_77/Y 0.04fF
C31710 INVX1_LOC_36/A INVX1_LOC_102/Y 0.10fF
C31711 NAND2X1_LOC_520/a_36_24# INVX1_LOC_90/A 0.00fF
C31712 NOR2X1_LOC_242/A INVX1_LOC_143/Y 0.01fF
C31713 INVX1_LOC_24/Y INVX1_LOC_65/A 0.10fF
C31714 NOR2X1_LOC_68/A NOR2X1_LOC_564/Y 0.03fF
C31715 INVX1_LOC_41/A NAND2X1_LOC_573/A 0.02fF
C31716 INVX1_LOC_32/A NOR2X1_LOC_721/B 0.11fF
C31717 NOR2X1_LOC_391/B INVX1_LOC_31/A 0.09fF
C31718 NOR2X1_LOC_267/A INVX1_LOC_102/Y 0.02fF
C31719 INVX1_LOC_202/A NOR2X1_LOC_473/B 0.17fF
C31720 INVX1_LOC_255/Y NOR2X1_LOC_87/B 0.07fF
C31721 INVX1_LOC_90/A NOR2X1_LOC_152/Y 0.07fF
C31722 NOR2X1_LOC_48/B INVX1_LOC_261/Y 0.03fF
C31723 NOR2X1_LOC_432/a_36_216# INVX1_LOC_22/A 0.00fF
C31724 NAND2X1_LOC_475/Y INVX1_LOC_94/Y 0.03fF
C31725 NAND2X1_LOC_37/a_36_24# INVX1_LOC_201/A 0.00fF
C31726 INVX1_LOC_80/A NOR2X1_LOC_6/B 0.11fF
C31727 NOR2X1_LOC_677/Y INVX1_LOC_92/A 0.08fF
C31728 INVX1_LOC_279/A NOR2X1_LOC_348/B 0.15fF
C31729 INVX1_LOC_1/Y NOR2X1_LOC_537/Y 0.03fF
C31730 INVX1_LOC_33/Y NOR2X1_LOC_652/Y 0.06fF
C31731 INVX1_LOC_24/A NAND2X1_LOC_560/A 0.03fF
C31732 NOR2X1_LOC_160/B NOR2X1_LOC_343/a_36_216# 0.00fF
C31733 NAND2X1_LOC_357/B INVX1_LOC_10/A 0.04fF
C31734 NAND2X1_LOC_726/Y NOR2X1_LOC_773/Y 0.01fF
C31735 INVX1_LOC_89/A INVX1_LOC_63/Y 0.13fF
C31736 NAND2X1_LOC_162/B NOR2X1_LOC_163/Y 0.02fF
C31737 NOR2X1_LOC_596/A INVX1_LOC_75/A 0.08fF
C31738 NOR2X1_LOC_605/B NOR2X1_LOC_773/Y 0.02fF
C31739 INVX1_LOC_26/A NOR2X1_LOC_814/A 0.02fF
C31740 NAND2X1_LOC_569/A INPUT_1 0.02fF
C31741 NAND2X1_LOC_725/B NOR2X1_LOC_27/a_36_216# 0.00fF
C31742 INVX1_LOC_181/Y INPUT_0 0.03fF
C31743 NOR2X1_LOC_194/Y NOR2X1_LOC_214/B 0.01fF
C31744 INVX1_LOC_182/Y NOR2X1_LOC_577/Y -0.01fF
C31745 NOR2X1_LOC_598/B NOR2X1_LOC_197/B 0.10fF
C31746 INVX1_LOC_103/A INVX1_LOC_46/A 0.07fF
C31747 INVX1_LOC_84/A INVX1_LOC_112/Y -0.03fF
C31748 NOR2X1_LOC_48/B NOR2X1_LOC_467/A 0.14fF
C31749 NAND2X1_LOC_195/Y NOR2X1_LOC_7/Y 0.01fF
C31750 NOR2X1_LOC_763/Y NAND2X1_LOC_451/Y 0.71fF
C31751 NOR2X1_LOC_790/B NOR2X1_LOC_445/B 0.02fF
C31752 INVX1_LOC_89/A NOR2X1_LOC_175/A 0.09fF
C31753 NAND2X1_LOC_61/Y INVX1_LOC_19/A 0.02fF
C31754 NOR2X1_LOC_318/B INVX1_LOC_72/A 0.15fF
C31755 INVX1_LOC_249/A INVX1_LOC_311/A 0.15fF
C31756 INVX1_LOC_97/Y NOR2X1_LOC_197/B 0.03fF
C31757 INVX1_LOC_224/Y INVX1_LOC_63/A 0.07fF
C31758 INVX1_LOC_75/A NOR2X1_LOC_712/Y 0.03fF
C31759 NOR2X1_LOC_332/A INVX1_LOC_40/A 0.11fF
C31760 INVX1_LOC_279/A INVX1_LOC_22/A 0.26fF
C31761 NAND2X1_LOC_223/A INVX1_LOC_42/A 0.03fF
C31762 NOR2X1_LOC_224/Y NOR2X1_LOC_697/Y 0.01fF
C31763 INVX1_LOC_72/A INVX1_LOC_93/Y 0.10fF
C31764 NOR2X1_LOC_160/B D_INPUT_3 0.01fF
C31765 NOR2X1_LOC_295/Y INVX1_LOC_75/A 0.02fF
C31766 INVX1_LOC_292/A INVX1_LOC_46/A 0.07fF
C31767 NOR2X1_LOC_434/Y NOR2X1_LOC_862/B 0.46fF
C31768 INVX1_LOC_182/Y NOR2X1_LOC_348/B 0.01fF
C31769 NOR2X1_LOC_481/a_36_216# INVX1_LOC_29/A 0.00fF
C31770 NAND2X1_LOC_860/A NAND2X1_LOC_489/Y 0.01fF
C31771 NOR2X1_LOC_570/B NOR2X1_LOC_188/A 0.00fF
C31772 INVX1_LOC_241/A NOR2X1_LOC_576/B 0.03fF
C31773 NOR2X1_LOC_521/Y INVX1_LOC_234/A 0.01fF
C31774 NOR2X1_LOC_416/a_36_216# NAND2X1_LOC_206/Y 0.01fF
C31775 NOR2X1_LOC_816/A NOR2X1_LOC_816/Y 0.02fF
C31776 INVX1_LOC_1/A INVX1_LOC_54/A 0.13fF
C31777 NAND2X1_LOC_838/Y INVX1_LOC_282/A 0.05fF
C31778 INVX1_LOC_135/A NAND2X1_LOC_859/Y 0.03fF
C31779 NAND2X1_LOC_563/Y INPUT_0 1.01fF
C31780 INPUT_1 INVX1_LOC_316/Y 0.03fF
C31781 INVX1_LOC_265/A NOR2X1_LOC_167/Y 0.15fF
C31782 INVX1_LOC_77/A INVX1_LOC_91/A 1.94fF
C31783 NAND2X1_LOC_796/B NOR2X1_LOC_88/Y 0.04fF
C31784 NOR2X1_LOC_294/Y INVX1_LOC_2/Y 0.04fF
C31785 NOR2X1_LOC_52/Y INVX1_LOC_76/A 0.03fF
C31786 INVX1_LOC_254/Y NOR2X1_LOC_78/A 0.02fF
C31787 INVX1_LOC_30/A NOR2X1_LOC_706/B 0.06fF
C31788 NOR2X1_LOC_589/Y NOR2X1_LOC_423/Y 0.06fF
C31789 NOR2X1_LOC_667/Y NOR2X1_LOC_536/A 0.01fF
C31790 INVX1_LOC_208/Y INVX1_LOC_28/A 0.02fF
C31791 NOR2X1_LOC_89/A INVX1_LOC_129/A 0.00fF
C31792 INVX1_LOC_237/Y NOR2X1_LOC_45/B 0.01fF
C31793 INVX1_LOC_18/A NOR2X1_LOC_305/Y 0.23fF
C31794 NOR2X1_LOC_576/B NOR2X1_LOC_298/Y 3.85fF
C31795 INVX1_LOC_132/A NOR2X1_LOC_405/A 0.00fF
C31796 NOR2X1_LOC_394/Y INVX1_LOC_165/A 0.00fF
C31797 INVX1_LOC_3/Y NAND2X1_LOC_99/A 0.00fF
C31798 NOR2X1_LOC_220/A INVX1_LOC_75/A 0.03fF
C31799 NOR2X1_LOC_773/Y NOR2X1_LOC_323/Y 0.04fF
C31800 INVX1_LOC_31/A INVX1_LOC_280/A 0.19fF
C31801 INVX1_LOC_78/A NAND2X1_LOC_223/A 0.07fF
C31802 INVX1_LOC_83/A INVX1_LOC_120/A 0.03fF
C31803 INVX1_LOC_182/Y INVX1_LOC_22/A 0.01fF
C31804 INVX1_LOC_21/A NAND2X1_LOC_477/Y 0.07fF
C31805 NOR2X1_LOC_232/a_36_216# NOR2X1_LOC_88/Y 0.03fF
C31806 INVX1_LOC_314/Y INVX1_LOC_20/A 0.09fF
C31807 NOR2X1_LOC_521/Y NOR2X1_LOC_19/B 0.10fF
C31808 INVX1_LOC_94/A VDD 0.10fF
C31809 INVX1_LOC_225/A NOR2X1_LOC_113/A 0.02fF
C31810 INVX1_LOC_34/A NOR2X1_LOC_675/A -0.01fF
C31811 INVX1_LOC_225/A NOR2X1_LOC_405/A 0.08fF
C31812 INVX1_LOC_124/A INVX1_LOC_91/A 0.54fF
C31813 INVX1_LOC_36/A NOR2X1_LOC_331/B 0.37fF
C31814 NOR2X1_LOC_75/Y INVX1_LOC_179/A 0.00fF
C31815 INVX1_LOC_90/A NAND2X1_LOC_861/Y 0.37fF
C31816 NOR2X1_LOC_366/B INVX1_LOC_6/A 0.03fF
C31817 INVX1_LOC_75/A NOR2X1_LOC_548/Y 0.13fF
C31818 INVX1_LOC_64/A NAND2X1_LOC_254/Y 0.09fF
C31819 INVX1_LOC_135/A NAND2X1_LOC_807/Y 0.10fF
C31820 NAND2X1_LOC_860/A INVX1_LOC_32/A 0.10fF
C31821 INVX1_LOC_277/Y NOR2X1_LOC_209/B 0.04fF
C31822 NOR2X1_LOC_27/Y INVX1_LOC_11/Y 0.06fF
C31823 NAND2X1_LOC_350/B NOR2X1_LOC_7/Y 0.10fF
C31824 NOR2X1_LOC_703/B INVX1_LOC_9/A 0.12fF
C31825 NOR2X1_LOC_667/A NOR2X1_LOC_528/Y 0.00fF
C31826 NOR2X1_LOC_785/A NOR2X1_LOC_445/B 0.03fF
C31827 INVX1_LOC_30/Y NOR2X1_LOC_83/a_36_216# 0.00fF
C31828 NOR2X1_LOC_447/Y INVX1_LOC_77/Y 0.01fF
C31829 INVX1_LOC_41/A NAND2X1_LOC_267/B 0.02fF
C31830 NOR2X1_LOC_687/Y NOR2X1_LOC_728/B 0.06fF
C31831 NAND2X1_LOC_227/Y NOR2X1_LOC_697/Y 0.02fF
C31832 INVX1_LOC_168/A NOR2X1_LOC_124/A 0.13fF
C31833 NAND2X1_LOC_361/Y INVX1_LOC_37/A 0.21fF
C31834 NAND2X1_LOC_479/Y INVX1_LOC_6/A 3.56fF
C31835 INVX1_LOC_77/A NOR2X1_LOC_698/Y 0.21fF
C31836 INVX1_LOC_232/A INVX1_LOC_123/A 0.20fF
C31837 NAND2X1_LOC_850/A INPUT_1 0.02fF
C31838 NOR2X1_LOC_92/Y NAND2X1_LOC_81/B 0.01fF
C31839 INVX1_LOC_95/Y INVX1_LOC_34/Y 0.38fF
C31840 NOR2X1_LOC_103/Y INVX1_LOC_63/A 0.07fF
C31841 INVX1_LOC_57/Y INVX1_LOC_71/Y 0.14fF
C31842 NOR2X1_LOC_288/A NOR2X1_LOC_857/A 0.08fF
C31843 NAND2X1_LOC_275/a_36_24# INVX1_LOC_87/A 0.00fF
C31844 NAND2X1_LOC_840/B NAND2X1_LOC_655/A 0.00fF
C31845 NAND2X1_LOC_465/Y VDD 0.08fF
C31846 INVX1_LOC_36/A NOR2X1_LOC_491/Y 0.03fF
C31847 INVX1_LOC_240/A INVX1_LOC_46/A 0.07fF
C31848 NOR2X1_LOC_152/Y INVX1_LOC_38/A 0.10fF
C31849 NOR2X1_LOC_234/Y VDD 0.35fF
C31850 INVX1_LOC_36/A NOR2X1_LOC_592/B 0.03fF
C31851 NOR2X1_LOC_456/Y NOR2X1_LOC_464/Y 0.02fF
C31852 NOR2X1_LOC_455/Y NOR2X1_LOC_465/Y 0.09fF
C31853 INPUT_0 INVX1_LOC_148/Y 0.02fF
C31854 NAND2X1_LOC_16/a_36_24# INVX1_LOC_113/A 0.01fF
C31855 NAND2X1_LOC_149/Y NOR2X1_LOC_470/a_36_216# 0.01fF
C31856 INVX1_LOC_113/Y INVX1_LOC_38/A 0.03fF
C31857 D_INPUT_1 INVX1_LOC_23/Y 0.19fF
C31858 NOR2X1_LOC_657/B NOR2X1_LOC_131/Y 0.05fF
C31859 INVX1_LOC_135/A INVX1_LOC_6/A 0.03fF
C31860 NOR2X1_LOC_78/B INVX1_LOC_143/Y 0.03fF
C31861 INVX1_LOC_58/A NAND2X1_LOC_99/A 0.02fF
C31862 INVX1_LOC_190/Y INVX1_LOC_144/A 0.01fF
C31863 INVX1_LOC_269/Y NOR2X1_LOC_777/B 0.01fF
C31864 NOR2X1_LOC_401/Y INVX1_LOC_76/A 0.07fF
C31865 INPUT_3 NOR2X1_LOC_721/B 0.03fF
C31866 NAND2X1_LOC_300/a_36_24# NOR2X1_LOC_536/A 0.00fF
C31867 NOR2X1_LOC_637/B INVX1_LOC_118/A 0.08fF
C31868 INVX1_LOC_159/A NOR2X1_LOC_155/A 0.17fF
C31869 NOR2X1_LOC_356/A NOR2X1_LOC_74/A 0.01fF
C31870 INVX1_LOC_30/A NOR2X1_LOC_430/Y 0.05fF
C31871 NOR2X1_LOC_423/Y INVX1_LOC_117/A 0.11fF
C31872 NOR2X1_LOC_589/A NOR2X1_LOC_657/B 0.03fF
C31873 NAND2X1_LOC_130/a_36_24# NOR2X1_LOC_139/Y 0.01fF
C31874 NAND2X1_LOC_787/A INVX1_LOC_181/A 0.01fF
C31875 NOR2X1_LOC_82/A INVX1_LOC_284/A 0.14fF
C31876 INVX1_LOC_25/A NAND2X1_LOC_215/A 0.14fF
C31877 INVX1_LOC_45/A INVX1_LOC_63/A 0.14fF
C31878 NOR2X1_LOC_663/A INVX1_LOC_175/A 0.02fF
C31879 INVX1_LOC_290/A NAND2X1_LOC_274/a_36_24# 0.00fF
C31880 NOR2X1_LOC_136/Y VDD 0.26fF
C31881 NAND2X1_LOC_569/A INVX1_LOC_118/A -0.02fF
C31882 NOR2X1_LOC_677/Y INVX1_LOC_53/A 0.03fF
C31883 NOR2X1_LOC_636/A INVX1_LOC_92/A 0.01fF
C31884 VDD INVX1_LOC_56/A 0.12fF
C31885 NOR2X1_LOC_383/a_36_216# INVX1_LOC_95/Y 0.11fF
C31886 NOR2X1_LOC_819/a_36_216# INVX1_LOC_63/A 0.00fF
C31887 NAND2X1_LOC_381/a_36_24# NOR2X1_LOC_847/B 0.00fF
C31888 NOR2X1_LOC_516/B D_INPUT_3 0.12fF
C31889 NOR2X1_LOC_222/Y INVX1_LOC_117/A 0.07fF
C31890 NAND2X1_LOC_130/a_36_24# NAND2X1_LOC_468/B 0.00fF
C31891 NOR2X1_LOC_542/Y NOR2X1_LOC_78/A 0.38fF
C31892 INVX1_LOC_239/A INVX1_LOC_253/A 0.02fF
C31893 NOR2X1_LOC_789/A INVX1_LOC_2/Y 0.01fF
C31894 INVX1_LOC_1/A NAND2X1_LOC_3/B 0.23fF
C31895 INVX1_LOC_83/A NOR2X1_LOC_542/B 0.02fF
C31896 NOR2X1_LOC_344/A INVX1_LOC_307/A 0.01fF
C31897 INVX1_LOC_5/A NOR2X1_LOC_635/B 0.00fF
C31898 INVX1_LOC_234/A NOR2X1_LOC_670/Y 0.32fF
C31899 NOR2X1_LOC_202/Y INVX1_LOC_6/A 0.04fF
C31900 INVX1_LOC_24/A NOR2X1_LOC_673/B 0.02fF
C31901 NOR2X1_LOC_197/Y INVX1_LOC_78/Y 0.01fF
C31902 NAND2X1_LOC_367/A NOR2X1_LOC_865/Y 0.24fF
C31903 INVX1_LOC_5/A NOR2X1_LOC_748/A 0.17fF
C31904 INVX1_LOC_83/A INVX1_LOC_143/Y 0.00fF
C31905 NOR2X1_LOC_74/A NOR2X1_LOC_9/Y 0.34fF
C31906 INVX1_LOC_58/Y NOR2X1_LOC_405/Y 0.04fF
C31907 INVX1_LOC_71/A INVX1_LOC_63/A 0.12fF
C31908 NAND2X1_LOC_537/Y NAND2X1_LOC_175/Y 0.08fF
C31909 INVX1_LOC_286/A NOR2X1_LOC_188/A 0.01fF
C31910 INVX1_LOC_2/A NAND2X1_LOC_487/a_36_24# 0.06fF
C31911 NOR2X1_LOC_19/B INVX1_LOC_255/A 0.07fF
C31912 NAND2X1_LOC_577/A INVX1_LOC_3/Y 0.07fF
C31913 NOR2X1_LOC_112/Y NOR2X1_LOC_332/B 0.09fF
C31914 INVX1_LOC_24/A INVX1_LOC_29/A 0.52fF
C31915 NOR2X1_LOC_598/B INVX1_LOC_38/Y 0.74fF
C31916 NOR2X1_LOC_360/Y NOR2X1_LOC_67/Y 0.03fF
C31917 NAND2X1_LOC_656/Y NOR2X1_LOC_363/Y 0.04fF
C31918 NAND2X1_LOC_859/Y INVX1_LOC_280/A 0.01fF
C31919 INVX1_LOC_143/A NOR2X1_LOC_634/A 0.48fF
C31920 NOR2X1_LOC_226/A NOR2X1_LOC_510/B 0.46fF
C31921 INVX1_LOC_41/Y NOR2X1_LOC_89/A 0.03fF
C31922 NAND2X1_LOC_141/A NAND2X1_LOC_141/Y 0.06fF
C31923 NOR2X1_LOC_520/B INVX1_LOC_19/A 0.07fF
C31924 INVX1_LOC_224/A NOR2X1_LOC_720/A 0.02fF
C31925 INVX1_LOC_8/A NAND2X1_LOC_773/B 0.83fF
C31926 INVX1_LOC_34/A NAND2X1_LOC_500/B 0.02fF
C31927 INVX1_LOC_96/Y NOR2X1_LOC_66/Y 0.09fF
C31928 NAND2X1_LOC_654/B INVX1_LOC_37/A 0.01fF
C31929 INVX1_LOC_144/A NOR2X1_LOC_56/Y 0.20fF
C31930 INVX1_LOC_41/A NAND2X1_LOC_81/B 0.03fF
C31931 NOR2X1_LOC_644/Y INVX1_LOC_84/A 0.08fF
C31932 NOR2X1_LOC_250/a_36_216# INVX1_LOC_50/A 0.00fF
C31933 INVX1_LOC_22/A NOR2X1_LOC_624/B 0.04fF
C31934 NOR2X1_LOC_557/Y INVX1_LOC_29/A 0.02fF
C31935 INVX1_LOC_30/Y NOR2X1_LOC_99/Y 0.00fF
C31936 INVX1_LOC_30/A INVX1_LOC_94/Y 0.30fF
C31937 NOR2X1_LOC_590/A INVX1_LOC_26/A 0.07fF
C31938 INVX1_LOC_21/A INVX1_LOC_99/Y 0.00fF
C31939 NOR2X1_LOC_264/Y NAND2X1_LOC_63/Y 0.05fF
C31940 INVX1_LOC_17/A NAND2X1_LOC_458/a_36_24# 0.01fF
C31941 NOR2X1_LOC_470/B NOR2X1_LOC_598/B 0.20fF
C31942 NOR2X1_LOC_706/A INVX1_LOC_14/Y 0.00fF
C31943 INVX1_LOC_256/A INVX1_LOC_270/Y 0.34fF
C31944 INVX1_LOC_233/Y NOR2X1_LOC_92/Y 1.66fF
C31945 NOR2X1_LOC_758/Y NOR2X1_LOC_89/A 0.46fF
C31946 INVX1_LOC_33/A INVX1_LOC_42/A 0.04fF
C31947 INVX1_LOC_21/A INVX1_LOC_93/A 0.07fF
C31948 NOR2X1_LOC_554/B NAND2X1_LOC_223/A 0.07fF
C31949 INVX1_LOC_18/A INVX1_LOC_271/Y 0.07fF
C31950 INVX1_LOC_144/A VDD 1.44fF
C31951 D_INPUT_1 NOR2X1_LOC_446/A 0.04fF
C31952 NAND2X1_LOC_357/B INVX1_LOC_12/A 0.07fF
C31953 D_INPUT_1 NAND2X1_LOC_563/a_36_24# 0.00fF
C31954 INVX1_LOC_50/A NOR2X1_LOC_254/a_36_216# 0.00fF
C31955 NOR2X1_LOC_626/Y INVX1_LOC_27/A 0.01fF
C31956 NOR2X1_LOC_68/A NOR2X1_LOC_158/Y 0.48fF
C31957 INVX1_LOC_11/A INPUT_6 0.02fF
C31958 NOR2X1_LOC_772/B NOR2X1_LOC_15/Y 0.22fF
C31959 INVX1_LOC_314/Y INVX1_LOC_4/A 0.10fF
C31960 NOR2X1_LOC_83/Y VDD 0.35fF
C31961 INVX1_LOC_230/Y NOR2X1_LOC_414/Y 0.04fF
C31962 NOR2X1_LOC_717/B INVX1_LOC_179/A 0.02fF
C31963 NAND2X1_LOC_35/Y NOR2X1_LOC_361/B 0.01fF
C31964 NOR2X1_LOC_67/A INVX1_LOC_19/A 0.07fF
C31965 NOR2X1_LOC_411/Y NAND2X1_LOC_725/B 0.15fF
C31966 INVX1_LOC_30/A INVX1_LOC_181/A 0.10fF
C31967 NOR2X1_LOC_730/B VDD 0.02fF
C31968 NOR2X1_LOC_387/A NAND2X1_LOC_448/a_36_24# 0.00fF
C31969 NOR2X1_LOC_15/Y INVX1_LOC_13/Y 0.13fF
C31970 INVX1_LOC_143/A INVX1_LOC_29/A 0.07fF
C31971 INVX1_LOC_6/A INVX1_LOC_139/Y 0.01fF
C31972 INVX1_LOC_30/A INVX1_LOC_296/A 0.05fF
C31973 INVX1_LOC_221/A NOR2X1_LOC_48/B 0.03fF
C31974 INVX1_LOC_90/A INVX1_LOC_291/A 0.07fF
C31975 NAND2X1_LOC_381/a_36_24# NOR2X1_LOC_660/Y 0.00fF
C31976 NOR2X1_LOC_824/A NAND2X1_LOC_778/a_36_24# 0.00fF
C31977 INVX1_LOC_258/Y INVX1_LOC_237/A 0.24fF
C31978 INVX1_LOC_58/A NAND2X1_LOC_577/A 0.03fF
C31979 INVX1_LOC_298/Y INVX1_LOC_24/A 0.03fF
C31980 NAND2X1_LOC_382/a_36_24# NOR2X1_LOC_660/Y 0.00fF
C31981 NOR2X1_LOC_459/A NAND2X1_LOC_659/A 0.09fF
C31982 NAND2X1_LOC_763/B INVX1_LOC_296/A 0.05fF
C31983 NOR2X1_LOC_824/A NAND2X1_LOC_634/a_36_24# 0.00fF
C31984 NOR2X1_LOC_516/Y INVX1_LOC_32/A 0.07fF
C31985 INVX1_LOC_315/Y D_INPUT_3 0.03fF
C31986 INVX1_LOC_8/A NOR2X1_LOC_393/Y 0.01fF
C31987 INVX1_LOC_255/Y NAND2X1_LOC_219/B 0.82fF
C31988 INVX1_LOC_79/A INVX1_LOC_9/A 0.01fF
C31989 NOR2X1_LOC_71/Y NAND2X1_LOC_572/B -0.02fF
C31990 INVX1_LOC_27/A NOR2X1_LOC_523/A -0.00fF
C31991 NOR2X1_LOC_68/A NOR2X1_LOC_646/B 0.02fF
C31992 NOR2X1_LOC_544/A INVX1_LOC_99/A 0.01fF
C31993 INVX1_LOC_24/Y NOR2X1_LOC_790/A 0.02fF
C31994 INVX1_LOC_41/A INVX1_LOC_4/Y 0.09fF
C31995 NOR2X1_LOC_403/B INVX1_LOC_23/Y 0.02fF
C31996 NAND2X1_LOC_582/a_36_24# INVX1_LOC_15/A 0.00fF
C31997 INVX1_LOC_33/A INVX1_LOC_78/A 0.19fF
C31998 NAND2X1_LOC_565/B INVX1_LOC_29/A 0.05fF
C31999 INVX1_LOC_40/A NOR2X1_LOC_847/A 0.01fF
C32000 INVX1_LOC_89/A INVX1_LOC_27/Y 0.03fF
C32001 NAND2X1_LOC_725/A INVX1_LOC_286/Y 0.37fF
C32002 NOR2X1_LOC_84/a_36_216# NOR2X1_LOC_38/B 0.00fF
C32003 INVX1_LOC_40/A INVX1_LOC_42/A 0.68fF
C32004 NOR2X1_LOC_123/B INVX1_LOC_63/A 0.07fF
C32005 NOR2X1_LOC_15/Y INVX1_LOC_88/A 0.05fF
C32006 NAND2X1_LOC_212/Y NAND2X1_LOC_211/Y 0.04fF
C32007 INVX1_LOC_269/A INVX1_LOC_14/A 0.11fF
C32008 INVX1_LOC_58/A NAND2X1_LOC_656/A 0.04fF
C32009 NOR2X1_LOC_749/Y INVX1_LOC_63/A 0.03fF
C32010 INVX1_LOC_243/Y INVX1_LOC_49/A 0.06fF
C32011 NAND2X1_LOC_463/B INVX1_LOC_241/Y 0.00fF
C32012 NAND2X1_LOC_705/Y NAND2X1_LOC_550/A 0.02fF
C32013 NOR2X1_LOC_65/B INVX1_LOC_33/A 0.13fF
C32014 INPUT_1 NOR2X1_LOC_662/A 0.01fF
C32015 INVX1_LOC_49/A INVX1_LOC_57/A 0.17fF
C32016 INPUT_3 NAND2X1_LOC_473/A 0.02fF
C32017 INVX1_LOC_91/A INVX1_LOC_9/A 0.11fF
C32018 NOR2X1_LOC_669/Y NOR2X1_LOC_816/A 0.04fF
C32019 NOR2X1_LOC_130/A INVX1_LOC_29/A 0.03fF
C32020 NAND2X1_LOC_573/A INVX1_LOC_168/Y 0.00fF
C32021 NOR2X1_LOC_447/B NAND2X1_LOC_453/A 0.03fF
C32022 NOR2X1_LOC_537/Y INVX1_LOC_87/A 0.06fF
C32023 INVX1_LOC_28/A NAND2X1_LOC_604/a_36_24# 0.00fF
C32024 INVX1_LOC_233/Y NAND2X1_LOC_837/Y 0.10fF
C32025 INVX1_LOC_102/Y INVX1_LOC_63/A 0.07fF
C32026 NAND2X1_LOC_798/A INVX1_LOC_78/A 0.22fF
C32027 NOR2X1_LOC_857/A NOR2X1_LOC_863/A 0.00fF
C32028 NOR2X1_LOC_43/Y INVX1_LOC_54/A 0.46fF
C32029 NOR2X1_LOC_132/a_36_216# INVX1_LOC_284/A 0.01fF
C32030 NOR2X1_LOC_211/A INVX1_LOC_4/Y 0.00fF
C32031 NOR2X1_LOC_337/Y NOR2X1_LOC_155/A 0.00fF
C32032 INVX1_LOC_60/A INVX1_LOC_57/A 0.01fF
C32033 INVX1_LOC_35/A NOR2X1_LOC_620/Y 0.03fF
C32034 INVX1_LOC_235/Y INVX1_LOC_195/Y 0.04fF
C32035 NOR2X1_LOC_753/Y NAND2X1_LOC_790/a_36_24# 0.01fF
C32036 INVX1_LOC_17/A INVX1_LOC_110/Y 0.06fF
C32037 INVX1_LOC_152/Y INVX1_LOC_33/A 0.03fF
C32038 INVX1_LOC_299/A INVX1_LOC_30/A 0.14fF
C32039 NOR2X1_LOC_795/Y INVX1_LOC_23/A 0.01fF
C32040 INVX1_LOC_21/A INVX1_LOC_212/A 0.01fF
C32041 INVX1_LOC_58/A NOR2X1_LOC_423/Y 0.02fF
C32042 NOR2X1_LOC_211/Y NOR2X1_LOC_593/Y 0.02fF
C32043 INVX1_LOC_2/A INVX1_LOC_57/A 0.20fF
C32044 NAND2X1_LOC_773/Y INVX1_LOC_18/A 0.07fF
C32045 NOR2X1_LOC_538/B INVX1_LOC_30/A 0.01fF
C32046 NAND2X1_LOC_773/a_36_24# INVX1_LOC_40/A 0.00fF
C32047 NOR2X1_LOC_848/Y INVX1_LOC_36/A 0.01fF
C32048 INVX1_LOC_21/A NOR2X1_LOC_303/Y 0.03fF
C32049 NAND2X1_LOC_711/Y NOR2X1_LOC_816/A 0.01fF
C32050 NAND2X1_LOC_787/A NOR2X1_LOC_315/Y 0.04fF
C32051 INVX1_LOC_244/Y NOR2X1_LOC_454/Y 0.04fF
C32052 NOR2X1_LOC_65/B INVX1_LOC_40/A 0.03fF
C32053 NOR2X1_LOC_181/A INVX1_LOC_179/A 0.01fF
C32054 NOR2X1_LOC_226/A INVX1_LOC_57/A 0.25fF
C32055 NOR2X1_LOC_67/A NAND2X1_LOC_557/Y 0.02fF
C32056 NOR2X1_LOC_656/a_36_216# INVX1_LOC_269/A 0.01fF
C32057 INVX1_LOC_25/A NOR2X1_LOC_655/B 2.03fF
C32058 INVX1_LOC_131/A NOR2X1_LOC_114/Y 0.10fF
C32059 NOR2X1_LOC_82/A INVX1_LOC_72/A 1.08fF
C32060 INVX1_LOC_58/A NOR2X1_LOC_222/Y 0.07fF
C32061 NOR2X1_LOC_410/Y INVX1_LOC_11/A 0.03fF
C32062 NOR2X1_LOC_78/A INVX1_LOC_84/A 0.57fF
C32063 NOR2X1_LOC_121/Y INVX1_LOC_306/Y 0.03fF
C32064 NAND2X1_LOC_512/a_36_24# INVX1_LOC_77/A 0.01fF
C32065 INVX1_LOC_282/A NAND2X1_LOC_254/Y 0.03fF
C32066 NAND2X1_LOC_809/A NOR2X1_LOC_409/B 0.01fF
C32067 NOR2X1_LOC_791/Y INVX1_LOC_162/A 0.02fF
C32068 NAND2X1_LOC_214/Y NOR2X1_LOC_643/Y 0.01fF
C32069 NOR2X1_LOC_614/Y INVX1_LOC_23/A 0.01fF
C32070 INVX1_LOC_39/A NAND2X1_LOC_569/A 0.02fF
C32071 INVX1_LOC_21/A NOR2X1_LOC_254/Y 0.03fF
C32072 NOR2X1_LOC_433/a_36_216# INVX1_LOC_27/A 0.01fF
C32073 NAND2X1_LOC_35/B NAND2X1_LOC_725/A 0.00fF
C32074 INVX1_LOC_41/A NOR2X1_LOC_790/A 0.08fF
C32075 D_INPUT_1 INVX1_LOC_232/A 0.01fF
C32076 INPUT_0 NOR2X1_LOC_114/Y 0.03fF
C32077 VDD NOR2X1_LOC_155/A 2.03fF
C32078 INVX1_LOC_35/A NAND2X1_LOC_181/Y 0.03fF
C32079 INVX1_LOC_64/A NOR2X1_LOC_778/B 0.04fF
C32080 NOR2X1_LOC_791/Y NOR2X1_LOC_315/Y 0.11fF
C32081 NOR2X1_LOC_666/Y INVX1_LOC_49/A 0.00fF
C32082 NOR2X1_LOC_589/A INVX1_LOC_271/A 0.03fF
C32083 NAND2X1_LOC_35/Y INVX1_LOC_280/Y 0.10fF
C32084 INVX1_LOC_55/Y NAND2X1_LOC_454/Y 0.07fF
C32085 NOR2X1_LOC_589/A INVX1_LOC_105/Y 0.04fF
C32086 NOR2X1_LOC_477/a_36_216# NOR2X1_LOC_68/A 0.00fF
C32087 NOR2X1_LOC_231/a_36_216# NOR2X1_LOC_751/Y 0.03fF
C32088 NAND2X1_LOC_564/B NAND2X1_LOC_860/A 0.07fF
C32089 NAND2X1_LOC_655/A INVX1_LOC_49/Y 0.02fF
C32090 INVX1_LOC_34/A NAND2X1_LOC_725/B 0.00fF
C32091 NOR2X1_LOC_87/Y INVX1_LOC_50/Y 0.05fF
C32092 NOR2X1_LOC_843/A INVX1_LOC_24/Y 0.03fF
C32093 NOR2X1_LOC_536/A NAND2X1_LOC_93/B 0.06fF
C32094 NOR2X1_LOC_565/A NOR2X1_LOC_703/B 0.01fF
C32095 INVX1_LOC_269/A INVX1_LOC_217/Y 0.02fF
C32096 INVX1_LOC_38/A INVX1_LOC_291/A 0.16fF
C32097 INVX1_LOC_21/A INVX1_LOC_54/Y 0.02fF
C32098 NOR2X1_LOC_15/Y NOR2X1_LOC_234/a_36_216# 0.00fF
C32099 INVX1_LOC_43/Y INVX1_LOC_314/Y 0.00fF
C32100 NOR2X1_LOC_667/A INVX1_LOC_93/A 0.02fF
C32101 NAND2X1_LOC_656/Y INVX1_LOC_29/Y 5.11fF
C32102 NAND2X1_LOC_740/Y NAND2X1_LOC_852/Y 0.03fF
C32103 INVX1_LOC_75/Y INVX1_LOC_193/A 0.22fF
C32104 NAND2X1_LOC_855/Y NAND2X1_LOC_175/Y 0.04fF
C32105 INVX1_LOC_25/A NOR2X1_LOC_99/B 1.60fF
C32106 INVX1_LOC_135/A NOR2X1_LOC_416/A 0.01fF
C32107 NAND2X1_LOC_190/Y NOR2X1_LOC_348/B 0.10fF
C32108 INVX1_LOC_280/Y NAND2X1_LOC_571/Y 0.01fF
C32109 NOR2X1_LOC_389/A NOR2X1_LOC_577/Y 0.03fF
C32110 NAND2X1_LOC_721/B INVX1_LOC_24/A 0.68fF
C32111 NOR2X1_LOC_690/A NAND2X1_LOC_550/A 0.01fF
C32112 NOR2X1_LOC_510/B INVX1_LOC_118/A 0.01fF
C32113 INPUT_1 INVX1_LOC_57/A 0.06fF
C32114 INVX1_LOC_39/A INVX1_LOC_316/Y 0.00fF
C32115 NAND2X1_LOC_214/B NAND2X1_LOC_666/a_36_24# 0.01fF
C32116 INVX1_LOC_2/A NOR2X1_LOC_666/Y 0.00fF
C32117 NAND2X1_LOC_1/Y INPUT_7 0.17fF
C32118 NAND2X1_LOC_651/a_36_24# NOR2X1_LOC_635/B 0.00fF
C32119 NOR2X1_LOC_728/B INVX1_LOC_274/Y 0.22fF
C32120 INVX1_LOC_24/A NAND2X1_LOC_634/Y 0.10fF
C32121 NOR2X1_LOC_655/B INVX1_LOC_1/A 0.01fF
C32122 INVX1_LOC_233/Y NOR2X1_LOC_299/Y 0.07fF
C32123 INVX1_LOC_269/A INVX1_LOC_111/Y 0.02fF
C32124 NAND2X1_LOC_9/Y INVX1_LOC_120/A 0.00fF
C32125 INVX1_LOC_59/Y INVX1_LOC_284/A 0.24fF
C32126 NAND2X1_LOC_298/a_36_24# INVX1_LOC_186/Y 0.00fF
C32127 INVX1_LOC_112/A INVX1_LOC_284/A 0.03fF
C32128 NOR2X1_LOC_2/Y NOR2X1_LOC_25/Y 0.47fF
C32129 INVX1_LOC_256/A NOR2X1_LOC_310/Y 0.03fF
C32130 NOR2X1_LOC_536/A INVX1_LOC_3/A 0.51fF
C32131 NOR2X1_LOC_78/A INVX1_LOC_15/A 0.34fF
C32132 NAND2X1_LOC_26/a_36_24# INVX1_LOC_174/A 0.00fF
C32133 NOR2X1_LOC_456/Y NOR2X1_LOC_180/B 0.07fF
C32134 NOR2X1_LOC_691/B INVX1_LOC_117/A 0.06fF
C32135 INVX1_LOC_135/A NOR2X1_LOC_109/Y 0.10fF
C32136 INVX1_LOC_5/A NOR2X1_LOC_719/a_36_216# 0.00fF
C32137 INVX1_LOC_27/A NOR2X1_LOC_589/A 0.11fF
C32138 INVX1_LOC_161/Y INVX1_LOC_133/Y 0.03fF
C32139 NOR2X1_LOC_435/A NOR2X1_LOC_592/B 0.01fF
C32140 NAND2X1_LOC_44/a_36_24# INVX1_LOC_49/A 0.00fF
C32141 NAND2X1_LOC_93/B NAND2X1_LOC_425/Y 1.49fF
C32142 NOR2X1_LOC_361/B NOR2X1_LOC_136/Y 0.06fF
C32143 NOR2X1_LOC_82/A NAND2X1_LOC_338/B 0.17fF
C32144 INVX1_LOC_276/A INVX1_LOC_161/Y 0.03fF
C32145 NOR2X1_LOC_278/a_36_216# INVX1_LOC_306/Y 0.00fF
C32146 NOR2X1_LOC_331/B INVX1_LOC_63/A 0.07fF
C32147 NOR2X1_LOC_831/B INVX1_LOC_92/A 0.07fF
C32148 NAND2X1_LOC_733/Y NAND2X1_LOC_357/B 0.01fF
C32149 INVX1_LOC_20/A INVX1_LOC_170/Y 0.00fF
C32150 VDD NOR2X1_LOC_833/B 0.05fF
C32151 NAND2X1_LOC_840/a_36_24# INVX1_LOC_141/Y 0.00fF
C32152 NOR2X1_LOC_468/Y INVX1_LOC_22/A 0.38fF
C32153 INVX1_LOC_5/A INVX1_LOC_89/A 14.90fF
C32154 NOR2X1_LOC_655/Y NOR2X1_LOC_649/B 0.13fF
C32155 NOR2X1_LOC_848/a_36_216# NOR2X1_LOC_332/A 0.01fF
C32156 NOR2X1_LOC_590/A INVX1_LOC_149/A 0.01fF
C32157 NOR2X1_LOC_655/Y INVX1_LOC_3/A 0.21fF
C32158 NAND2X1_LOC_190/Y INVX1_LOC_22/A 0.90fF
C32159 NAND2X1_LOC_208/B NOR2X1_LOC_398/a_36_216# 0.15fF
C32160 NOR2X1_LOC_662/A INVX1_LOC_118/A 0.10fF
C32161 NOR2X1_LOC_315/Y INVX1_LOC_30/A 0.03fF
C32162 NOR2X1_LOC_596/A NOR2X1_LOC_577/Y 0.08fF
C32163 INVX1_LOC_289/A NAND2X1_LOC_227/Y 0.03fF
C32164 INVX1_LOC_64/A NAND2X1_LOC_123/Y 0.00fF
C32165 NAND2X1_LOC_93/B INVX1_LOC_3/A 0.02fF
C32166 INVX1_LOC_5/A NAND2X1_LOC_508/A 0.03fF
C32167 NAND2X1_LOC_569/A INVX1_LOC_61/A 0.01fF
C32168 NOR2X1_LOC_729/A INVX1_LOC_19/A 0.49fF
C32169 NOR2X1_LOC_42/a_36_216# INVX1_LOC_3/Y 0.01fF
C32170 NOR2X1_LOC_103/Y INVX1_LOC_1/Y 0.00fF
C32171 NAND2X1_LOC_207/B INVX1_LOC_230/A 0.02fF
C32172 NOR2X1_LOC_865/Y NOR2X1_LOC_243/B 0.02fF
C32173 NAND2X1_LOC_36/A INVX1_LOC_192/Y 0.86fF
C32174 NOR2X1_LOC_433/A NAND2X1_LOC_593/Y 1.01fF
C32175 NOR2X1_LOC_486/Y INVX1_LOC_78/A 0.03fF
C32176 NOR2X1_LOC_209/Y NOR2X1_LOC_726/Y 0.33fF
C32177 INVX1_LOC_254/Y INVX1_LOC_132/A 0.01fF
C32178 NOR2X1_LOC_91/A NOR2X1_LOC_45/B 0.04fF
C32179 NAND2X1_LOC_711/Y NOR2X1_LOC_773/Y 0.01fF
C32180 INVX1_LOC_104/A NOR2X1_LOC_360/Y 0.10fF
C32181 NOR2X1_LOC_477/B INVX1_LOC_117/A 0.02fF
C32182 INVX1_LOC_24/A INVX1_LOC_8/A 0.23fF
C32183 INVX1_LOC_125/A NAND2X1_LOC_62/a_36_24# 0.00fF
C32184 NAND2X1_LOC_49/a_36_24# INVX1_LOC_230/Y 0.01fF
C32185 NOR2X1_LOC_592/B INVX1_LOC_63/A 0.00fF
C32186 INVX1_LOC_21/A NOR2X1_LOC_112/Y 0.65fF
C32187 NAND2X1_LOC_785/A NOR2X1_LOC_91/Y 1.51fF
C32188 NOR2X1_LOC_389/A INVX1_LOC_22/A 0.01fF
C32189 INVX1_LOC_269/A NOR2X1_LOC_137/A 0.07fF
C32190 NOR2X1_LOC_790/a_36_216# NOR2X1_LOC_542/Y 0.00fF
C32191 NOR2X1_LOC_52/B INVX1_LOC_41/Y 0.03fF
C32192 INVX1_LOC_279/A NOR2X1_LOC_787/a_36_216# 0.00fF
C32193 INVX1_LOC_226/A NOR2X1_LOC_500/B 0.12fF
C32194 NOR2X1_LOC_649/B INVX1_LOC_3/A 0.07fF
C32195 NOR2X1_LOC_15/Y NAND2X1_LOC_308/B 0.02fF
C32196 NAND2X1_LOC_361/Y INVX1_LOC_310/Y 0.31fF
C32197 NOR2X1_LOC_703/B INVX1_LOC_179/Y 0.02fF
C32198 NOR2X1_LOC_220/A NOR2X1_LOC_274/B 0.07fF
C32199 NOR2X1_LOC_617/Y NOR2X1_LOC_52/B 0.02fF
C32200 NOR2X1_LOC_45/B INVX1_LOC_23/A 0.13fF
C32201 NOR2X1_LOC_155/A INVX1_LOC_133/A 0.45fF
C32202 NOR2X1_LOC_89/A INVX1_LOC_185/A 1.40fF
C32203 NOR2X1_LOC_52/B NAND2X1_LOC_593/Y 0.07fF
C32204 INVX1_LOC_45/A INVX1_LOC_1/Y 0.00fF
C32205 INVX1_LOC_41/A NOR2X1_LOC_843/A 0.03fF
C32206 INVX1_LOC_40/A NOR2X1_LOC_554/B 0.20fF
C32207 INVX1_LOC_30/A INVX1_LOC_268/Y 0.11fF
C32208 NAND2X1_LOC_337/B NOR2X1_LOC_110/a_36_216# 0.00fF
C32209 NOR2X1_LOC_197/B INVX1_LOC_29/A 0.01fF
C32210 INVX1_LOC_278/A INVX1_LOC_98/A 0.35fF
C32211 NOR2X1_LOC_510/Y INVX1_LOC_144/A 0.07fF
C32212 INVX1_LOC_62/Y NOR2X1_LOC_346/B 0.07fF
C32213 INVX1_LOC_97/Y NOR2X1_LOC_337/Y 0.10fF
C32214 INVX1_LOC_108/Y NOR2X1_LOC_78/A 0.05fF
C32215 INVX1_LOC_50/A NOR2X1_LOC_631/B 0.68fF
C32216 INVX1_LOC_36/A NAND2X1_LOC_479/Y 0.01fF
C32217 NAND2X1_LOC_225/a_36_24# NOR2X1_LOC_814/A 0.01fF
C32218 NOR2X1_LOC_182/a_36_216# NOR2X1_LOC_550/B 0.13fF
C32219 INVX1_LOC_278/A NOR2X1_LOC_78/A 0.06fF
C32220 NOR2X1_LOC_784/Y NOR2X1_LOC_803/A 0.29fF
C32221 NOR2X1_LOC_816/Y INVX1_LOC_78/A 0.01fF
C32222 INVX1_LOC_147/Y INVX1_LOC_271/A 0.24fF
C32223 INVX1_LOC_45/Y NOR2X1_LOC_757/Y 0.14fF
C32224 INVX1_LOC_201/Y INVX1_LOC_82/A 0.04fF
C32225 NAND2X1_LOC_563/Y NOR2X1_LOC_514/a_36_216# 0.01fF
C32226 NOR2X1_LOC_61/B INPUT_0 0.28fF
C32227 INVX1_LOC_241/Y INVX1_LOC_42/A 0.03fF
C32228 INVX1_LOC_314/Y NAND2X1_LOC_850/Y 0.22fF
C32229 D_INPUT_1 NAND2X1_LOC_447/Y 0.00fF
C32230 INVX1_LOC_229/A NOR2X1_LOC_380/Y 0.07fF
C32231 NAND2X1_LOC_564/B NAND2X1_LOC_640/a_36_24# 0.00fF
C32232 INVX1_LOC_13/A NOR2X1_LOC_68/A 0.22fF
C32233 NAND2X1_LOC_430/B INVX1_LOC_92/A 0.09fF
C32234 NAND2X1_LOC_287/B NAND2X1_LOC_287/a_36_24# 0.00fF
C32235 NOR2X1_LOC_473/B NOR2X1_LOC_276/Y 0.02fF
C32236 INVX1_LOC_200/Y NAND2X1_LOC_242/a_36_24# 0.00fF
C32237 INVX1_LOC_208/A NOR2X1_LOC_106/Y 0.02fF
C32238 NOR2X1_LOC_689/Y VDD 0.12fF
C32239 INVX1_LOC_95/A NOR2X1_LOC_129/a_36_216# 0.00fF
C32240 NOR2X1_LOC_596/A INVX1_LOC_22/A 0.12fF
C32241 INVX1_LOC_279/A INVX1_LOC_18/A 0.07fF
C32242 INVX1_LOC_50/A INVX1_LOC_37/A 0.10fF
C32243 INVX1_LOC_64/A NOR2X1_LOC_657/B 0.28fF
C32244 NAND2X1_LOC_141/Y NOR2X1_LOC_128/a_36_216# 0.01fF
C32245 INVX1_LOC_36/A INVX1_LOC_135/A 0.11fF
C32246 VDD NOR2X1_LOC_125/Y 0.24fF
C32247 INVX1_LOC_215/Y NOR2X1_LOC_329/B 0.08fF
C32248 INVX1_LOC_1/Y INVX1_LOC_71/A 0.17fF
C32249 NOR2X1_LOC_711/Y INVX1_LOC_213/A 0.06fF
C32250 NOR2X1_LOC_769/B VDD -0.00fF
C32251 NOR2X1_LOC_351/Y INVX1_LOC_78/A 0.02fF
C32252 NOR2X1_LOC_208/Y NAND2X1_LOC_479/Y 0.03fF
C32253 NOR2X1_LOC_794/B INVX1_LOC_182/A 0.02fF
C32254 NOR2X1_LOC_468/Y INVX1_LOC_100/A 0.08fF
C32255 INVX1_LOC_143/A INVX1_LOC_8/A 0.10fF
C32256 NOR2X1_LOC_413/Y NOR2X1_LOC_399/a_36_216# 0.01fF
C32257 INVX1_LOC_278/A NAND2X1_LOC_464/A 0.03fF
C32258 NOR2X1_LOC_498/Y NOR2X1_LOC_526/Y 0.00fF
C32259 NOR2X1_LOC_316/Y NOR2X1_LOC_709/A 0.02fF
C32260 NOR2X1_LOC_598/B VDD 4.57fF
C32261 D_INPUT_6 NOR2X1_LOC_588/A 0.17fF
C32262 NOR2X1_LOC_246/A NOR2X1_LOC_68/A 0.03fF
C32263 NOR2X1_LOC_331/B NOR2X1_LOC_65/Y 0.00fF
C32264 INVX1_LOC_51/A VDD -0.00fF
C32265 INVX1_LOC_5/A NOR2X1_LOC_24/Y 0.00fF
C32266 INVX1_LOC_30/A NOR2X1_LOC_166/Y 0.02fF
C32267 INVX1_LOC_245/Y NOR2X1_LOC_74/A 0.20fF
C32268 INVX1_LOC_155/Y INVX1_LOC_16/A 0.03fF
C32269 NAND2X1_LOC_721/A NAND2X1_LOC_793/B 0.07fF
C32270 NOR2X1_LOC_220/A NOR2X1_LOC_348/B 0.30fF
C32271 INVX1_LOC_97/Y VDD 0.21fF
C32272 NAND2X1_LOC_214/B INVX1_LOC_20/A 0.03fF
C32273 NAND2X1_LOC_477/Y INVX1_LOC_19/Y 0.19fF
C32274 NAND2X1_LOC_725/A VDD 4.64fF
C32275 NAND2X1_LOC_717/Y NOR2X1_LOC_822/Y 0.06fF
C32276 NOR2X1_LOC_295/Y INVX1_LOC_22/A 0.00fF
C32277 NOR2X1_LOC_68/A INVX1_LOC_55/Y 0.08fF
C32278 NAND2X1_LOC_725/A NAND2X1_LOC_800/A 0.03fF
C32279 NOR2X1_LOC_449/A NOR2X1_LOC_435/A 0.37fF
C32280 NAND2X1_LOC_715/B VDD 0.71fF
C32281 NOR2X1_LOC_205/a_36_216# INVX1_LOC_177/A 0.00fF
C32282 NOR2X1_LOC_298/Y NAND2X1_LOC_864/a_36_24# 0.09fF
C32283 INVX1_LOC_45/A NOR2X1_LOC_742/A 0.03fF
C32284 INVX1_LOC_280/A NOR2X1_LOC_416/A 0.04fF
C32285 INVX1_LOC_35/A INVX1_LOC_117/A 0.41fF
C32286 NAND2X1_LOC_445/a_36_24# INVX1_LOC_19/A 0.00fF
C32287 INVX1_LOC_218/Y NOR2X1_LOC_188/A 0.13fF
C32288 INVX1_LOC_135/A NOR2X1_LOC_237/Y 0.03fF
C32289 INVX1_LOC_23/A NOR2X1_LOC_499/B 0.01fF
C32290 INVX1_LOC_57/A INVX1_LOC_118/A 0.23fF
C32291 NOR2X1_LOC_266/B INVX1_LOC_306/Y 0.00fF
C32292 INVX1_LOC_27/A INVX1_LOC_20/A 0.11fF
C32293 NOR2X1_LOC_93/a_36_216# INVX1_LOC_316/Y 0.00fF
C32294 NOR2X1_LOC_590/Y INVX1_LOC_37/A 0.04fF
C32295 NOR2X1_LOC_636/A INVX1_LOC_83/A 0.07fF
C32296 INVX1_LOC_13/Y NAND2X1_LOC_266/a_36_24# 0.01fF
C32297 INVX1_LOC_124/Y NOR2X1_LOC_74/A 0.59fF
C32298 NOR2X1_LOC_520/A INVX1_LOC_218/A 0.00fF
C32299 NOR2X1_LOC_824/A INVX1_LOC_20/A 0.02fF
C32300 NAND2X1_LOC_363/B NAND2X1_LOC_93/a_36_24# 0.00fF
C32301 NOR2X1_LOC_843/B NOR2X1_LOC_624/B 0.01fF
C32302 INVX1_LOC_135/A NOR2X1_LOC_804/B 0.07fF
C32303 NOR2X1_LOC_716/B NOR2X1_LOC_71/Y -0.02fF
C32304 NOR2X1_LOC_148/A INVX1_LOC_75/A 0.01fF
C32305 NOR2X1_LOC_662/A NAND2X1_LOC_618/Y 0.02fF
C32306 NOR2X1_LOC_841/A NAND2X1_LOC_61/Y 0.41fF
C32307 INVX1_LOC_124/Y NOR2X1_LOC_9/Y 0.04fF
C32308 NOR2X1_LOC_180/B NOR2X1_LOC_550/B 0.10fF
C32309 NOR2X1_LOC_78/B INVX1_LOC_56/Y 0.03fF
C32310 INVX1_LOC_33/A NOR2X1_LOC_150/a_36_216# 0.01fF
C32311 NOR2X1_LOC_130/A INVX1_LOC_8/A 0.13fF
C32312 NOR2X1_LOC_671/a_36_216# INVX1_LOC_3/Y 0.01fF
C32313 INVX1_LOC_189/Y INVX1_LOC_22/A 0.01fF
C32314 NAND2X1_LOC_509/a_36_24# NOR2X1_LOC_45/B 0.00fF
C32315 INVX1_LOC_135/A NOR2X1_LOC_309/Y 0.10fF
C32316 NAND2X1_LOC_858/B INVX1_LOC_18/A 0.08fF
C32317 INVX1_LOC_80/A NAND2X1_LOC_141/A 0.01fF
C32318 NAND2X1_LOC_357/B NAND2X1_LOC_808/A 0.01fF
C32319 NOR2X1_LOC_220/A INVX1_LOC_22/A 0.07fF
C32320 INVX1_LOC_23/A NOR2X1_LOC_862/B 0.01fF
C32321 NOR2X1_LOC_621/B INVX1_LOC_63/A 0.01fF
C32322 NAND2X1_LOC_254/Y NOR2X1_LOC_496/a_36_216# 0.00fF
C32323 NOR2X1_LOC_742/A INVX1_LOC_71/A 0.02fF
C32324 NOR2X1_LOC_361/Y NAND2X1_LOC_656/Y 0.01fF
C32325 INVX1_LOC_31/A NOR2X1_LOC_45/B 0.58fF
C32326 INVX1_LOC_202/A INVX1_LOC_73/A 0.03fF
C32327 INVX1_LOC_89/A NOR2X1_LOC_377/Y 0.01fF
C32328 NOR2X1_LOC_111/A NAND2X1_LOC_780/Y 0.03fF
C32329 INVX1_LOC_28/A INVX1_LOC_155/Y 0.03fF
C32330 INVX1_LOC_45/A NOR2X1_LOC_318/B 0.23fF
C32331 NAND2X1_LOC_863/B INVX1_LOC_22/A 0.08fF
C32332 INVX1_LOC_53/A NOR2X1_LOC_831/B 0.43fF
C32333 INVX1_LOC_221/Y INVX1_LOC_76/A 0.07fF
C32334 NOR2X1_LOC_169/B INVX1_LOC_91/A 0.05fF
C32335 NAND2X1_LOC_338/B INVX1_LOC_306/A 0.03fF
C32336 NOR2X1_LOC_318/B NOR2X1_LOC_568/A -0.03fF
C32337 INVX1_LOC_94/A INVX1_LOC_285/Y 0.22fF
C32338 INVX1_LOC_14/A INVX1_LOC_12/Y 0.39fF
C32339 NOR2X1_LOC_548/Y INVX1_LOC_22/A 0.07fF
C32340 INVX1_LOC_102/A NAND2X1_LOC_444/B 0.03fF
C32341 NOR2X1_LOC_248/a_36_216# NOR2X1_LOC_309/Y 0.00fF
C32342 INVX1_LOC_311/A NOR2X1_LOC_303/Y 0.01fF
C32343 NAND2X1_LOC_839/Y NAND2X1_LOC_866/B 0.03fF
C32344 INVX1_LOC_45/A INVX1_LOC_93/Y 0.07fF
C32345 NOR2X1_LOC_716/B NOR2X1_LOC_751/A 0.02fF
C32346 INVX1_LOC_75/A INVX1_LOC_63/Y 0.10fF
C32347 NOR2X1_LOC_569/A NOR2X1_LOC_550/B 0.10fF
C32348 INVX1_LOC_164/A NOR2X1_LOC_82/Y 0.03fF
C32349 NOR2X1_LOC_481/A NOR2X1_LOC_335/B 0.01fF
C32350 INVX1_LOC_33/A INVX1_LOC_158/Y 0.00fF
C32351 INVX1_LOC_46/Y INVX1_LOC_306/Y 0.02fF
C32352 NOR2X1_LOC_372/A VDD 0.12fF
C32353 NOR2X1_LOC_67/Y INVX1_LOC_26/A 0.27fF
C32354 NOR2X1_LOC_209/Y INVX1_LOC_311/Y 0.04fF
C32355 NOR2X1_LOC_355/A NAND2X1_LOC_349/a_36_24# 0.00fF
C32356 NOR2X1_LOC_510/Y NOR2X1_LOC_155/A 0.00fF
C32357 NAND2X1_LOC_326/A INVX1_LOC_54/A 0.08fF
C32358 INVX1_LOC_130/Y NOR2X1_LOC_657/B 0.09fF
C32359 NAND2X1_LOC_656/Y INVX1_LOC_101/A 0.06fF
C32360 NOR2X1_LOC_318/B INVX1_LOC_71/A 0.10fF
C32361 INVX1_LOC_1/Y NOR2X1_LOC_123/B 0.07fF
C32362 NAND2X1_LOC_63/Y INVX1_LOC_57/A 0.13fF
C32363 NOR2X1_LOC_827/a_36_216# INVX1_LOC_31/Y 0.00fF
C32364 INVX1_LOC_256/A NOR2X1_LOC_536/A 0.03fF
C32365 NAND2X1_LOC_330/a_36_24# NOR2X1_LOC_318/B 0.00fF
C32366 NOR2X1_LOC_804/B NOR2X1_LOC_794/A 0.11fF
C32367 INVX1_LOC_21/A INVX1_LOC_35/Y 0.51fF
C32368 INVX1_LOC_141/Y NOR2X1_LOC_111/A 0.10fF
C32369 INVX1_LOC_63/Y NOR2X1_LOC_7/a_36_216# 0.00fF
C32370 INVX1_LOC_93/Y INVX1_LOC_71/A 0.10fF
C32371 INVX1_LOC_94/A NOR2X1_LOC_137/B 0.05fF
C32372 NOR2X1_LOC_500/Y NOR2X1_LOC_564/Y 0.02fF
C32373 INVX1_LOC_312/Y NOR2X1_LOC_111/A -0.00fF
C32374 INVX1_LOC_254/Y NAND2X1_LOC_642/Y 0.40fF
C32375 NOR2X1_LOC_355/A NAND2X1_LOC_656/Y 0.07fF
C32376 NOR2X1_LOC_186/Y INVX1_LOC_84/A 0.09fF
C32377 INVX1_LOC_13/Y NAND2X1_LOC_456/Y 0.03fF
C32378 INVX1_LOC_11/A INVX1_LOC_185/A 0.00fF
C32379 INVX1_LOC_36/A NOR2X1_LOC_558/a_36_216# 0.00fF
C32380 NOR2X1_LOC_655/B NOR2X1_LOC_188/A 0.10fF
C32381 NOR2X1_LOC_361/B NOR2X1_LOC_155/A 0.03fF
C32382 INVX1_LOC_89/A NOR2X1_LOC_332/A 0.22fF
C32383 INVX1_LOC_36/A NOR2X1_LOC_152/A 0.04fF
C32384 INVX1_LOC_251/Y INVX1_LOC_6/A 0.01fF
C32385 NAND2X1_LOC_784/A NOR2X1_LOC_48/B 0.07fF
C32386 NOR2X1_LOC_647/B NOR2X1_LOC_655/Y 0.01fF
C32387 INVX1_LOC_128/A NAND2X1_LOC_61/Y 0.01fF
C32388 NAND2X1_LOC_35/Y NAND2X1_LOC_81/B 0.03fF
C32389 NOR2X1_LOC_544/A INPUT_0 0.46fF
C32390 INVX1_LOC_36/A INVX1_LOC_10/Y 0.01fF
C32391 NOR2X1_LOC_577/Y NAND2X1_LOC_655/B 0.01fF
C32392 INVX1_LOC_256/A NAND2X1_LOC_93/B 3.89fF
C32393 D_GATE_741 INVX1_LOC_92/A 0.07fF
C32394 INVX1_LOC_71/A INVX1_LOC_139/A 0.06fF
C32395 INVX1_LOC_21/A NOR2X1_LOC_721/B 0.03fF
C32396 NOR2X1_LOC_781/B NAND2X1_LOC_654/B 0.10fF
C32397 NOR2X1_LOC_106/Y NAND2X1_LOC_211/Y 0.13fF
C32398 INVX1_LOC_36/A INVX1_LOC_280/A 0.03fF
C32399 NOR2X1_LOC_717/B NOR2X1_LOC_644/A 0.00fF
C32400 NOR2X1_LOC_25/Y NOR2X1_LOC_36/A 0.02fF
C32401 NAND2X1_LOC_508/A NOR2X1_LOC_332/A 0.07fF
C32402 D_INPUT_0 NOR2X1_LOC_356/A 0.07fF
C32403 INVX1_LOC_35/A NOR2X1_LOC_460/A 0.01fF
C32404 NAND2X1_LOC_624/B NAND2X1_LOC_254/Y 0.00fF
C32405 NAND2X1_LOC_724/A INVX1_LOC_84/A 0.08fF
C32406 INVX1_LOC_13/Y NAND2X1_LOC_80/a_36_24# 0.01fF
C32407 NOR2X1_LOC_717/B NOR2X1_LOC_828/B 0.00fF
C32408 NOR2X1_LOC_309/Y NOR2X1_LOC_566/a_36_216# 0.02fF
C32409 NOR2X1_LOC_246/a_36_216# NOR2X1_LOC_389/B 0.01fF
C32410 NAND2X1_LOC_464/Y NAND2X1_LOC_464/A 0.15fF
C32411 NOR2X1_LOC_304/Y INVX1_LOC_42/A 0.29fF
C32412 INVX1_LOC_35/A INVX1_LOC_3/Y 0.07fF
C32413 INVX1_LOC_50/A NAND2X1_LOC_72/B 0.03fF
C32414 NOR2X1_LOC_208/Y NOR2X1_LOC_57/a_36_216# 0.00fF
C32415 NOR2X1_LOC_828/A NOR2X1_LOC_644/A 0.10fF
C32416 NOR2X1_LOC_606/Y NAND2X1_LOC_93/B 0.02fF
C32417 INVX1_LOC_179/Y INVX1_LOC_91/A 0.03fF
C32418 NOR2X1_LOC_400/a_36_216# NOR2X1_LOC_415/Y 0.00fF
C32419 NAND2X1_LOC_562/B NOR2X1_LOC_24/Y 0.01fF
C32420 NOR2X1_LOC_720/B NOR2X1_LOC_35/Y 0.04fF
C32421 INVX1_LOC_202/A NOR2X1_LOC_122/a_36_216# 0.00fF
C32422 INVX1_LOC_63/Y NAND2X1_LOC_453/A 0.01fF
C32423 NOR2X1_LOC_152/Y NOR2X1_LOC_816/Y 0.03fF
C32424 INVX1_LOC_27/A NOR2X1_LOC_128/A 0.03fF
C32425 NOR2X1_LOC_848/Y INVX1_LOC_63/A 0.05fF
C32426 INVX1_LOC_23/A NOR2X1_LOC_685/B 0.07fF
C32427 NOR2X1_LOC_194/a_36_216# INVX1_LOC_54/A 0.00fF
C32428 INVX1_LOC_45/A INVX1_LOC_117/Y 0.03fF
C32429 INVX1_LOC_135/A NOR2X1_LOC_19/Y 0.03fF
C32430 NOR2X1_LOC_647/B NOR2X1_LOC_649/B 0.01fF
C32431 NOR2X1_LOC_647/B INVX1_LOC_3/A 0.03fF
C32432 NAND2X1_LOC_462/B NAND2X1_LOC_621/a_36_24# 0.00fF
C32433 NAND2X1_LOC_231/Y NAND2X1_LOC_468/B 0.05fF
C32434 NAND2X1_LOC_308/Y VDD 0.04fF
C32435 D_INPUT_0 NOR2X1_LOC_74/A 0.09fF
C32436 INVX1_LOC_88/A INVX1_LOC_49/Y 0.02fF
C32437 NAND2X1_LOC_347/B INVX1_LOC_12/A 0.00fF
C32438 NOR2X1_LOC_188/A NOR2X1_LOC_99/B 0.07fF
C32439 NOR2X1_LOC_286/Y INVX1_LOC_19/A 0.03fF
C32440 NOR2X1_LOC_353/a_36_216# INVX1_LOC_9/A 0.02fF
C32441 NAND2X1_LOC_214/B INVX1_LOC_4/A 0.03fF
C32442 NOR2X1_LOC_186/Y INVX1_LOC_15/A 0.07fF
C32443 NOR2X1_LOC_647/a_36_216# INVX1_LOC_63/A 0.00fF
C32444 D_INPUT_0 NOR2X1_LOC_9/Y 0.07fF
C32445 INVX1_LOC_91/Y NAND2X1_LOC_866/B 0.01fF
C32446 NOR2X1_LOC_152/Y NOR2X1_LOC_351/Y 0.65fF
C32447 VDD NOR2X1_LOC_156/B 0.28fF
C32448 NAND2X1_LOC_859/Y NOR2X1_LOC_45/B 0.03fF
C32449 NAND2X1_LOC_338/B INVX1_LOC_176/A 0.01fF
C32450 VDD NAND2X1_LOC_660/A 0.06fF
C32451 NAND2X1_LOC_72/Y NAND2X1_LOC_72/B 0.03fF
C32452 NOR2X1_LOC_606/Y INVX1_LOC_3/A 0.01fF
C32453 NOR2X1_LOC_561/Y INVX1_LOC_91/A 0.17fF
C32454 INVX1_LOC_183/Y NOR2X1_LOC_167/Y 0.01fF
C32455 INVX1_LOC_257/Y INVX1_LOC_117/A 0.01fF
C32456 NOR2X1_LOC_828/B NOR2X1_LOC_151/Y 0.00fF
C32457 INVX1_LOC_7/A INVX1_LOC_91/A 0.44fF
C32458 NOR2X1_LOC_292/Y INVX1_LOC_87/Y 0.09fF
C32459 NAND2X1_LOC_323/B INVX1_LOC_176/A 0.08fF
C32460 INVX1_LOC_49/A INVX1_LOC_274/A 0.07fF
C32461 NAND2X1_LOC_276/Y INVX1_LOC_9/A 0.03fF
C32462 INVX1_LOC_27/A INVX1_LOC_4/A 0.09fF
C32463 NOR2X1_LOC_414/a_36_216# NAND2X1_LOC_206/Y 0.01fF
C32464 NAND2X1_LOC_573/Y INVX1_LOC_15/A 0.07fF
C32465 INVX1_LOC_90/A NOR2X1_LOC_147/A 0.01fF
C32466 NOR2X1_LOC_392/B NAND2X1_LOC_297/a_36_24# 0.06fF
C32467 NAND2X1_LOC_363/B NAND2X1_LOC_99/A 0.07fF
C32468 INVX1_LOC_22/A NAND2X1_LOC_469/B 0.02fF
C32469 INVX1_LOC_14/A NOR2X1_LOC_554/A 0.04fF
C32470 NAND2X1_LOC_807/A NAND2X1_LOC_807/B 0.02fF
C32471 NOR2X1_LOC_695/Y INVX1_LOC_20/A 0.02fF
C32472 NOR2X1_LOC_91/A NOR2X1_LOC_53/Y 0.04fF
C32473 D_INPUT_3 INVX1_LOC_316/Y 0.28fF
C32474 NOR2X1_LOC_99/B NOR2X1_LOC_100/a_36_216# 0.01fF
C32475 NOR2X1_LOC_249/Y NOR2X1_LOC_34/Y 0.02fF
C32476 NOR2X1_LOC_717/A INVX1_LOC_29/Y 0.40fF
C32477 INVX1_LOC_286/Y INVX1_LOC_29/A 0.00fF
C32478 NOR2X1_LOC_45/B NAND2X1_LOC_866/B 0.09fF
C32479 INVX1_LOC_93/Y NOR2X1_LOC_123/B 0.01fF
C32480 NOR2X1_LOC_447/B INVX1_LOC_22/A 0.00fF
C32481 NAND2X1_LOC_618/Y NOR2X1_LOC_475/A 0.07fF
C32482 INVX1_LOC_58/A INVX1_LOC_35/A 0.29fF
C32483 INVX1_LOC_64/A INVX1_LOC_271/A 0.54fF
C32484 NOR2X1_LOC_717/B NOR2X1_LOC_540/B 0.02fF
C32485 INVX1_LOC_61/A NOR2X1_LOC_662/A 0.04fF
C32486 NAND2X1_LOC_116/A NOR2X1_LOC_61/Y 0.00fF
C32487 NOR2X1_LOC_561/Y NOR2X1_LOC_421/Y 0.05fF
C32488 NOR2X1_LOC_300/Y INVX1_LOC_54/A 0.03fF
C32489 NOR2X1_LOC_458/Y NOR2X1_LOC_155/A 0.01fF
C32490 NOR2X1_LOC_570/A VDD 0.24fF
C32491 NOR2X1_LOC_790/B INVX1_LOC_53/A 0.01fF
C32492 INVX1_LOC_153/Y NOR2X1_LOC_155/A 0.01fF
C32493 NOR2X1_LOC_52/B INVX1_LOC_185/A 0.03fF
C32494 INVX1_LOC_234/A INVX1_LOC_20/A 0.07fF
C32495 NOR2X1_LOC_45/B NAND2X1_LOC_807/Y 0.07fF
C32496 NOR2X1_LOC_352/Y INVX1_LOC_9/A 0.05fF
C32497 INVX1_LOC_21/A NAND2X1_LOC_286/B 0.03fF
C32498 NAND2X1_LOC_357/B INVX1_LOC_92/A 0.07fF
C32499 NOR2X1_LOC_802/A NOR2X1_LOC_640/Y 0.07fF
C32500 NOR2X1_LOC_596/A INVX1_LOC_186/Y 0.35fF
C32501 NOR2X1_LOC_45/Y INVX1_LOC_15/A 0.03fF
C32502 INVX1_LOC_159/A INVX1_LOC_29/A 0.07fF
C32503 INVX1_LOC_39/A INVX1_LOC_57/A 0.03fF
C32504 NOR2X1_LOC_481/A INVX1_LOC_84/A 0.00fF
C32505 INVX1_LOC_124/A NAND2X1_LOC_647/a_36_24# 0.00fF
C32506 NAND2X1_LOC_656/Y NOR2X1_LOC_111/A 0.07fF
C32507 INVX1_LOC_93/Y INVX1_LOC_102/Y 0.09fF
C32508 INVX1_LOC_233/Y NAND2X1_LOC_35/Y 0.17fF
C32509 INVX1_LOC_5/A NOR2X1_LOC_392/Y 0.11fF
C32510 INVX1_LOC_34/A NOR2X1_LOC_66/Y 0.01fF
C32511 NAND2X1_LOC_53/Y NOR2X1_LOC_158/Y 0.02fF
C32512 INVX1_LOC_82/A NAND2X1_LOC_574/A 0.03fF
C32513 NOR2X1_LOC_191/B INVX1_LOC_29/A 0.02fF
C32514 INVX1_LOC_17/A NOR2X1_LOC_278/Y 0.01fF
C32515 INVX1_LOC_225/A INVX1_LOC_84/A 0.07fF
C32516 INVX1_LOC_21/A NAND2X1_LOC_860/A 0.10fF
C32517 INVX1_LOC_64/A NAND2X1_LOC_214/B 0.27fF
C32518 NOR2X1_LOC_6/B NOR2X1_LOC_673/A 0.05fF
C32519 NOR2X1_LOC_286/Y INVX1_LOC_26/Y 0.01fF
C32520 NOR2X1_LOC_19/B INVX1_LOC_20/A 0.02fF
C32521 NOR2X1_LOC_818/Y NOR2X1_LOC_820/Y 0.01fF
C32522 NAND2X1_LOC_654/B NOR2X1_LOC_585/Y 0.01fF
C32523 NOR2X1_LOC_553/B INVX1_LOC_9/A 0.06fF
C32524 NOR2X1_LOC_78/B NOR2X1_LOC_831/B 0.07fF
C32525 INVX1_LOC_269/A NOR2X1_LOC_383/B 0.14fF
C32526 NAND2X1_LOC_562/Y NOR2X1_LOC_662/A 0.07fF
C32527 NOR2X1_LOC_470/B INVX1_LOC_204/A 0.04fF
C32528 NOR2X1_LOC_151/Y NOR2X1_LOC_540/B 0.03fF
C32529 INVX1_LOC_178/A NOR2X1_LOC_392/Y 0.01fF
C32530 NOR2X1_LOC_45/B INVX1_LOC_6/A 2.11fF
C32531 INVX1_LOC_64/A INVX1_LOC_27/A 0.15fF
C32532 INVX1_LOC_135/A NOR2X1_LOC_865/A 0.03fF
C32533 NOR2X1_LOC_68/A INVX1_LOC_32/A 0.12fF
C32534 NOR2X1_LOC_617/Y NAND2X1_LOC_254/Y 0.01fF
C32535 NAND2X1_LOC_341/A NOR2X1_LOC_364/A 0.02fF
C32536 NOR2X1_LOC_78/A INVX1_LOC_123/A 0.10fF
C32537 INPUT_0 NAND2X1_LOC_468/B 0.05fF
C32538 INVX1_LOC_64/A NOR2X1_LOC_824/A 0.07fF
C32539 NOR2X1_LOC_510/Y NAND2X1_LOC_715/B 0.02fF
C32540 INVX1_LOC_233/Y NAND2X1_LOC_571/Y 0.05fF
C32541 INVX1_LOC_223/Y INVX1_LOC_5/A 0.03fF
C32542 NOR2X1_LOC_441/Y NOR2X1_LOC_338/a_36_216# 0.00fF
C32543 NAND2X1_LOC_560/A VDD 0.83fF
C32544 INVX1_LOC_79/A INVX1_LOC_76/A 0.10fF
C32545 INVX1_LOC_224/Y NOR2X1_LOC_82/A 1.48fF
C32546 NAND2X1_LOC_563/Y INVX1_LOC_19/A 0.03fF
C32547 INVX1_LOC_64/A INVX1_LOC_237/A 0.03fF
C32548 NOR2X1_LOC_440/Y NAND2X1_LOC_93/B 0.07fF
C32549 INVX1_LOC_185/Y INVX1_LOC_29/A 0.02fF
C32550 NOR2X1_LOC_604/Y INVX1_LOC_103/A 0.06fF
C32551 NOR2X1_LOC_74/A NOR2X1_LOC_266/B 0.03fF
C32552 INVX1_LOC_136/A NOR2X1_LOC_464/Y 0.02fF
C32553 NAND2X1_LOC_861/Y NOR2X1_LOC_177/a_36_216# 0.01fF
C32554 NAND2X1_LOC_534/a_36_24# INVX1_LOC_49/Y 0.00fF
C32555 INVX1_LOC_249/A INVX1_LOC_4/A 0.00fF
C32556 NAND2X1_LOC_350/a_36_24# NOR2X1_LOC_435/A 0.00fF
C32557 INVX1_LOC_94/A INVX1_LOC_4/Y 0.10fF
C32558 INVX1_LOC_30/A NAND2X1_LOC_99/A 0.05fF
C32559 INVX1_LOC_309/A INVX1_LOC_76/A 0.00fF
C32560 NOR2X1_LOC_68/A NAND2X1_LOC_175/Y 0.07fF
C32561 INVX1_LOC_132/A INVX1_LOC_15/A 0.18fF
C32562 NOR2X1_LOC_374/A INVX1_LOC_15/A 0.03fF
C32563 NOR2X1_LOC_9/Y NOR2X1_LOC_266/B 0.04fF
C32564 NOR2X1_LOC_220/A INVX1_LOC_186/Y 0.10fF
C32565 INVX1_LOC_21/A NAND2X1_LOC_473/A 0.07fF
C32566 NOR2X1_LOC_375/Y INVX1_LOC_203/A 0.00fF
C32567 NOR2X1_LOC_361/B NAND2X1_LOC_715/B 0.20fF
C32568 INVX1_LOC_119/A INVX1_LOC_42/A 0.00fF
C32569 NAND2X1_LOC_352/B INVX1_LOC_53/A 0.14fF
C32570 NOR2X1_LOC_62/a_36_216# INVX1_LOC_293/Y 0.01fF
C32571 INVX1_LOC_71/A INVX1_LOC_87/A 0.01fF
C32572 NOR2X1_LOC_551/B NOR2X1_LOC_801/B 0.01fF
C32573 NOR2X1_LOC_596/Y NOR2X1_LOC_678/A 0.01fF
C32574 INVX1_LOC_91/A INVX1_LOC_76/A 0.37fF
C32575 NAND2X1_LOC_848/A NOR2X1_LOC_74/A 0.10fF
C32576 INVX1_LOC_21/A NAND2X1_LOC_537/Y 0.07fF
C32577 INVX1_LOC_11/Y NOR2X1_LOC_824/Y 0.05fF
C32578 INVX1_LOC_225/A INVX1_LOC_15/A 0.03fF
C32579 NOR2X1_LOC_778/Y INVX1_LOC_23/A 0.06fF
C32580 NOR2X1_LOC_68/A INVX1_LOC_262/A 0.02fF
C32581 INVX1_LOC_6/A INVX1_LOC_281/A 0.37fF
C32582 NOR2X1_LOC_664/Y INVX1_LOC_4/A 0.03fF
C32583 INVX1_LOC_69/Y NOR2X1_LOC_536/A 0.02fF
C32584 INVX1_LOC_11/Y INVX1_LOC_76/A 5.07fF
C32585 INVX1_LOC_50/A NAND2X1_LOC_198/B 0.03fF
C32586 INVX1_LOC_278/A INVX1_LOC_170/A 0.01fF
C32587 NOR2X1_LOC_270/Y INVX1_LOC_23/A 0.01fF
C32588 INVX1_LOC_135/A INVX1_LOC_63/A 0.15fF
C32589 INVX1_LOC_292/A NOR2X1_LOC_674/Y 0.02fF
C32590 NOR2X1_LOC_225/a_36_216# NOR2X1_LOC_652/Y 0.01fF
C32591 NAND2X1_LOC_9/Y NAND2X1_LOC_351/A 0.00fF
C32592 NOR2X1_LOC_209/Y INVX1_LOC_15/A 0.07fF
C32593 NOR2X1_LOC_419/Y NOR2X1_LOC_39/Y 0.10fF
C32594 NOR2X1_LOC_815/A INVX1_LOC_54/A 0.05fF
C32595 NOR2X1_LOC_391/B NOR2X1_LOC_656/Y 0.01fF
C32596 NOR2X1_LOC_172/Y NAND2X1_LOC_61/Y 0.01fF
C32597 NOR2X1_LOC_165/Y NOR2X1_LOC_48/B 0.04fF
C32598 INVX1_LOC_27/A INVX1_LOC_43/Y 0.02fF
C32599 INVX1_LOC_34/Y NOR2X1_LOC_38/B 0.09fF
C32600 INVX1_LOC_13/Y NAND2X1_LOC_208/B 0.15fF
C32601 INVX1_LOC_119/A INVX1_LOC_78/A 0.03fF
C32602 INVX1_LOC_256/A NOR2X1_LOC_348/Y 0.10fF
C32603 NOR2X1_LOC_464/B NOR2X1_LOC_457/A 0.01fF
C32604 INVX1_LOC_314/Y INVX1_LOC_129/A 0.01fF
C32605 NOR2X1_LOC_433/A INVX1_LOC_270/Y 0.07fF
C32606 INVX1_LOC_209/Y INVX1_LOC_296/Y 0.03fF
C32607 NOR2X1_LOC_91/A INVX1_LOC_265/A 0.01fF
C32608 NAND2X1_LOC_363/B NAND2X1_LOC_656/A 0.02fF
C32609 INVX1_LOC_69/Y NAND2X1_LOC_93/B 0.07fF
C32610 INVX1_LOC_104/A INVX1_LOC_26/A 0.00fF
C32611 NOR2X1_LOC_121/A INVX1_LOC_3/Y 0.01fF
C32612 NAND2X1_LOC_190/Y NOR2X1_LOC_787/a_36_216# 0.00fF
C32613 NAND2X1_LOC_293/a_36_24# INVX1_LOC_3/A 0.02fF
C32614 NOR2X1_LOC_9/Y INVX1_LOC_46/Y -0.01fF
C32615 INVX1_LOC_285/Y NOR2X1_LOC_155/A 0.03fF
C32616 NOR2X1_LOC_76/A NAND2X1_LOC_74/B 0.12fF
C32617 NOR2X1_LOC_844/A NOR2X1_LOC_843/B 0.03fF
C32618 INPUT_0 NAND2X1_LOC_141/Y 0.11fF
C32619 NOR2X1_LOC_160/B INVX1_LOC_14/A 0.22fF
C32620 NOR2X1_LOC_82/A NOR2X1_LOC_103/Y 0.18fF
C32621 NOR2X1_LOC_346/Y INVX1_LOC_230/A 0.05fF
C32622 INVX1_LOC_76/A NOR2X1_LOC_698/Y 0.01fF
C32623 NOR2X1_LOC_848/a_36_216# NOR2X1_LOC_554/B 0.00fF
C32624 INVX1_LOC_137/A INVX1_LOC_4/A 0.03fF
C32625 NOR2X1_LOC_52/B INVX1_LOC_270/Y 0.33fF
C32626 INVX1_LOC_89/A INVX1_LOC_42/A 10.90fF
C32627 NOR2X1_LOC_562/A INVX1_LOC_44/A 0.02fF
C32628 NOR2X1_LOC_598/B INVX1_LOC_153/Y 0.11fF
C32629 NOR2X1_LOC_667/Y INVX1_LOC_11/A 0.04fF
C32630 NOR2X1_LOC_91/A NAND2X1_LOC_596/a_36_24# 0.01fF
C32631 NOR2X1_LOC_180/Y INVX1_LOC_23/A 0.05fF
C32632 NOR2X1_LOC_152/Y NOR2X1_LOC_304/Y 0.42fF
C32633 NOR2X1_LOC_667/A NAND2X1_LOC_286/B 0.11fF
C32634 NOR2X1_LOC_725/A NAND2X1_LOC_425/Y 0.04fF
C32635 NAND2X1_LOC_579/A NOR2X1_LOC_384/Y 0.09fF
C32636 NOR2X1_LOC_598/B INVX1_LOC_121/Y 0.02fF
C32637 NOR2X1_LOC_145/Y INVX1_LOC_38/A 0.05fF
C32638 NOR2X1_LOC_19/B NOR2X1_LOC_128/A 0.01fF
C32639 NOR2X1_LOC_391/B INVX1_LOC_63/A 0.09fF
C32640 NAND2X1_LOC_357/B INVX1_LOC_53/A 0.01fF
C32641 NAND2X1_LOC_562/B NOR2X1_LOC_392/Y 0.07fF
C32642 NAND2X1_LOC_219/a_36_24# INVX1_LOC_36/A 0.00fF
C32643 D_INPUT_1 NOR2X1_LOC_644/Y 0.01fF
C32644 NOR2X1_LOC_813/Y NOR2X1_LOC_102/a_36_216# 0.01fF
C32645 NOR2X1_LOC_689/Y INVX1_LOC_280/Y 0.08fF
C32646 INVX1_LOC_103/A INVX1_LOC_72/A 0.07fF
C32647 NOR2X1_LOC_401/Y INVX1_LOC_23/A 0.06fF
C32648 NOR2X1_LOC_598/B INVX1_LOC_177/A 0.05fF
C32649 INVX1_LOC_314/Y NOR2X1_LOC_440/B 0.01fF
C32650 INVX1_LOC_157/A NAND2X1_LOC_470/B 0.01fF
C32651 NOR2X1_LOC_428/a_36_216# INVX1_LOC_30/A 0.01fF
C32652 INVX1_LOC_50/A NOR2X1_LOC_219/Y 0.08fF
C32653 INVX1_LOC_34/A INVX1_LOC_13/Y 0.08fF
C32654 INVX1_LOC_50/A INVX1_LOC_53/Y 0.00fF
C32655 INVX1_LOC_295/A NAND2X1_LOC_452/Y 0.05fF
C32656 NOR2X1_LOC_216/B INVX1_LOC_20/A 0.01fF
C32657 VDD INVX1_LOC_152/A 0.24fF
C32658 NAND2X1_LOC_740/Y GATE_811 0.25fF
C32659 NOR2X1_LOC_205/Y INVX1_LOC_94/A 0.01fF
C32660 INVX1_LOC_17/Y INVX1_LOC_16/A 0.02fF
C32661 INVX1_LOC_84/A NAND2X1_LOC_642/Y 0.07fF
C32662 INVX1_LOC_126/Y NOR2X1_LOC_89/A 0.12fF
C32663 INVX1_LOC_292/A INVX1_LOC_72/A 0.03fF
C32664 INVX1_LOC_21/A NOR2X1_LOC_486/B 1.25fF
C32665 INVX1_LOC_89/A INVX1_LOC_78/A 0.09fF
C32666 NOR2X1_LOC_552/A INVX1_LOC_63/A 0.07fF
C32667 VDD NOR2X1_LOC_634/A 0.53fF
C32668 NOR2X1_LOC_749/Y INVX1_LOC_87/A 0.04fF
C32669 NAND2X1_LOC_345/a_36_24# INVX1_LOC_78/A 0.00fF
C32670 NOR2X1_LOC_19/B INVX1_LOC_4/A 0.01fF
C32671 NAND2X1_LOC_735/B INVX1_LOC_57/A 0.00fF
C32672 INVX1_LOC_50/A NOR2X1_LOC_665/A 0.15fF
C32673 INPUT_3 NOR2X1_LOC_68/A 0.03fF
C32674 NAND2X1_LOC_555/Y INVX1_LOC_122/Y 0.00fF
C32675 NOR2X1_LOC_92/Y INVX1_LOC_207/A 0.08fF
C32676 NOR2X1_LOC_598/B NAND2X1_LOC_162/A 0.04fF
C32677 INVX1_LOC_45/A NAND2X1_LOC_36/A 0.02fF
C32678 NAND2X1_LOC_721/a_36_24# NOR2X1_LOC_406/A 0.00fF
C32679 NOR2X1_LOC_831/B INVX1_LOC_46/A 0.63fF
C32680 NOR2X1_LOC_389/A INVX1_LOC_18/A 0.10fF
C32681 NOR2X1_LOC_337/Y INVX1_LOC_29/A 0.02fF
C32682 VDD NOR2X1_LOC_58/Y -0.00fF
C32683 NOR2X1_LOC_527/Y NOR2X1_LOC_48/B 0.15fF
C32684 NAND2X1_LOC_725/A INVX1_LOC_280/Y 0.05fF
C32685 NOR2X1_LOC_82/A INVX1_LOC_71/A 0.49fF
C32686 NOR2X1_LOC_816/Y INVX1_LOC_291/A 0.02fF
C32687 NAND2X1_LOC_734/B INVX1_LOC_178/A 0.02fF
C32688 NAND2X1_LOC_586/a_36_24# NAND2X1_LOC_350/A 0.01fF
C32689 INVX1_LOC_147/A INVX1_LOC_32/A 0.03fF
C32690 INVX1_LOC_17/A NAND2X1_LOC_7/Y 0.07fF
C32691 NAND2X1_LOC_35/Y NOR2X1_LOC_526/Y 0.02fF
C32692 INVX1_LOC_148/Y INVX1_LOC_26/Y 0.03fF
C32693 NOR2X1_LOC_201/a_36_216# NOR2X1_LOC_68/A 0.00fF
C32694 NAND2X1_LOC_199/B INVX1_LOC_18/A 0.03fF
C32695 NOR2X1_LOC_582/a_36_216# INVX1_LOC_30/A 0.01fF
C32696 NOR2X1_LOC_92/Y NOR2X1_LOC_792/B 0.01fF
C32697 NOR2X1_LOC_226/A INVX1_LOC_306/Y 0.01fF
C32698 NAND2X1_LOC_477/Y INVX1_LOC_20/A 0.07fF
C32699 INVX1_LOC_224/Y INVX1_LOC_306/A 0.01fF
C32700 INVX1_LOC_34/A INVX1_LOC_88/A 0.04fF
C32701 NOR2X1_LOC_65/B INVX1_LOC_89/A 3.94fF
C32702 INVX1_LOC_101/A NOR2X1_LOC_717/A 0.01fF
C32703 NOR2X1_LOC_639/B INVX1_LOC_290/A 0.07fF
C32704 NOR2X1_LOC_859/Y NOR2X1_LOC_243/B 0.00fF
C32705 NAND2X1_LOC_199/a_36_24# INVX1_LOC_30/A 0.01fF
C32706 VDD NOR2X1_LOC_673/B -0.00fF
C32707 NOR2X1_LOC_598/B NOR2X1_LOC_785/Y 0.03fF
C32708 NAND2X1_LOC_553/A INVX1_LOC_56/Y 0.01fF
C32709 INVX1_LOC_5/A NAND2X1_LOC_716/a_36_24# 0.00fF
C32710 INVX1_LOC_162/Y INVX1_LOC_308/Y 0.09fF
C32711 NAND2X1_LOC_656/A INVX1_LOC_30/A 0.01fF
C32712 INVX1_LOC_136/A NOR2X1_LOC_457/B 0.42fF
C32713 NAND2X1_LOC_577/a_36_24# INVX1_LOC_178/A 0.00fF
C32714 INVX1_LOC_107/A INVX1_LOC_18/A 0.01fF
C32715 INVX1_LOC_64/A INVX1_LOC_234/A 0.11fF
C32716 NOR2X1_LOC_355/A NOR2X1_LOC_717/A 0.10fF
C32717 NOR2X1_LOC_329/B NOR2X1_LOC_135/a_36_216# 0.01fF
C32718 INVX1_LOC_64/A NAND2X1_LOC_156/B 0.05fF
C32719 NOR2X1_LOC_302/Y NAND2X1_LOC_299/a_36_24# 0.00fF
C32720 INVX1_LOC_269/A NOR2X1_LOC_168/A 0.03fF
C32721 NAND2X1_LOC_785/B NOR2X1_LOC_753/Y 0.01fF
C32722 INVX1_LOC_17/Y INVX1_LOC_28/A 0.08fF
C32723 NOR2X1_LOC_596/A INVX1_LOC_18/A 0.14fF
C32724 NOR2X1_LOC_496/Y INVX1_LOC_22/A 0.11fF
C32725 NAND2X1_LOC_231/Y INVX1_LOC_88/A 0.01fF
C32726 NOR2X1_LOC_667/A NAND2X1_LOC_537/Y 0.01fF
C32727 NOR2X1_LOC_394/a_36_216# INVX1_LOC_26/A 0.00fF
C32728 VDD INVX1_LOC_29/A 1.93fF
C32729 INVX1_LOC_84/A NOR2X1_LOC_271/Y 0.03fF
C32730 NAND2X1_LOC_179/a_36_24# NOR2X1_LOC_180/Y 0.00fF
C32731 NAND2X1_LOC_642/Y INVX1_LOC_15/A 1.64fF
C32732 INVX1_LOC_280/A INVX1_LOC_63/A 0.14fF
C32733 NOR2X1_LOC_592/B INVX1_LOC_117/Y 0.00fF
C32734 NAND2X1_LOC_244/A INVX1_LOC_42/A 0.06fF
C32735 INVX1_LOC_136/A NAND2X1_LOC_833/Y 0.07fF
C32736 INVX1_LOC_95/Y INVX1_LOC_47/Y 0.03fF
C32737 NOR2X1_LOC_272/Y NAND2X1_LOC_656/Y 0.10fF
C32738 NOR2X1_LOC_516/B INVX1_LOC_14/A 0.10fF
C32739 INVX1_LOC_51/Y NOR2X1_LOC_843/B 0.04fF
C32740 NOR2X1_LOC_641/Y NOR2X1_LOC_814/A 0.02fF
C32741 INVX1_LOC_41/A NOR2X1_LOC_360/Y 0.03fF
C32742 NOR2X1_LOC_78/B NAND2X1_LOC_352/B 0.72fF
C32743 INVX1_LOC_64/A NOR2X1_LOC_19/B 0.15fF
C32744 INPUT_1 INVX1_LOC_306/Y 0.05fF
C32745 NOR2X1_LOC_295/Y INVX1_LOC_18/A 0.02fF
C32746 INVX1_LOC_72/A INVX1_LOC_240/A 5.36fF
C32747 INVX1_LOC_255/Y NOR2X1_LOC_817/a_36_216# 0.00fF
C32748 INVX1_LOC_76/A INVX1_LOC_231/A 0.03fF
C32749 INVX1_LOC_125/A INVX1_LOC_9/A 0.05fF
C32750 NOR2X1_LOC_89/A NOR2X1_LOC_536/A 0.14fF
C32751 NOR2X1_LOC_336/B NOR2X1_LOC_168/B 0.04fF
C32752 NAND2X1_LOC_181/a_36_24# NOR2X1_LOC_103/Y 0.00fF
C32753 INVX1_LOC_207/A NAND2X1_LOC_837/Y 0.07fF
C32754 INVX1_LOC_120/A NAND2X1_LOC_85/a_36_24# 0.01fF
C32755 INVX1_LOC_28/A NOR2X1_LOC_406/A 0.20fF
C32756 NOR2X1_LOC_613/Y NAND2X1_LOC_866/B 0.20fF
C32757 NOR2X1_LOC_592/A NOR2X1_LOC_561/Y 0.00fF
C32758 NOR2X1_LOC_222/Y INVX1_LOC_30/A 0.16fF
C32759 INVX1_LOC_5/A INVX1_LOC_75/A 0.38fF
C32760 INVX1_LOC_78/A NAND2X1_LOC_244/A 0.01fF
C32761 D_INPUT_1 INVX1_LOC_98/A 0.07fF
C32762 INVX1_LOC_45/A NAND2X1_LOC_59/a_36_24# 0.02fF
C32763 NOR2X1_LOC_103/Y INVX1_LOC_306/A 0.00fF
C32764 NAND2X1_LOC_149/Y NAND2X1_LOC_654/B 0.04fF
C32765 NAND2X1_LOC_180/a_36_24# INVX1_LOC_71/A 0.00fF
C32766 NOR2X1_LOC_90/a_36_216# INVX1_LOC_25/Y 0.00fF
C32767 NOR2X1_LOC_250/Y D_INPUT_0 0.26fF
C32768 INVX1_LOC_17/A NOR2X1_LOC_312/Y 0.01fF
C32769 D_INPUT_1 NOR2X1_LOC_78/A 0.10fF
C32770 INVX1_LOC_83/A D_GATE_741 0.01fF
C32771 INVX1_LOC_211/Y INVX1_LOC_10/A 0.08fF
C32772 NOR2X1_LOC_498/Y INVX1_LOC_207/A 0.08fF
C32773 INVX1_LOC_119/A NOR2X1_LOC_152/Y 0.10fF
C32774 NOR2X1_LOC_220/A INVX1_LOC_18/A 0.12fF
C32775 NOR2X1_LOC_82/A NOR2X1_LOC_123/B 0.00fF
C32776 NOR2X1_LOC_658/Y NOR2X1_LOC_222/a_36_216# 0.01fF
C32777 NOR2X1_LOC_89/A NAND2X1_LOC_93/B 0.24fF
C32778 INVX1_LOC_13/Y INPUT_0 0.17fF
C32779 INVX1_LOC_1/A NOR2X1_LOC_756/Y 0.01fF
C32780 INVX1_LOC_186/A NOR2X1_LOC_678/A 0.17fF
C32781 INVX1_LOC_298/Y VDD 0.24fF
C32782 NAND2X1_LOC_287/B NOR2X1_LOC_301/A 0.08fF
C32783 INVX1_LOC_77/A NOR2X1_LOC_709/A 0.01fF
C32784 NOR2X1_LOC_824/A INVX1_LOC_282/A 0.07fF
C32785 NOR2X1_LOC_860/B NOR2X1_LOC_87/Y 0.04fF
C32786 INVX1_LOC_224/Y INVX1_LOC_59/Y 0.00fF
C32787 VDD NOR2X1_LOC_33/Y 0.14fF
C32788 INVX1_LOC_223/A NOR2X1_LOC_569/Y 0.00fF
C32789 NOR2X1_LOC_565/A NOR2X1_LOC_553/B 0.01fF
C32790 INVX1_LOC_30/A INVX1_LOC_220/Y 0.03fF
C32791 NOR2X1_LOC_89/A NAND2X1_LOC_425/Y 0.10fF
C32792 NOR2X1_LOC_598/B INVX1_LOC_65/A 0.30fF
C32793 INVX1_LOC_24/Y NOR2X1_LOC_567/B 0.37fF
C32794 NAND2X1_LOC_489/Y NAND2X1_LOC_768/Y 0.23fF
C32795 NAND2X1_LOC_53/Y INVX1_LOC_55/Y 0.07fF
C32796 NOR2X1_LOC_656/a_36_216# NOR2X1_LOC_516/B 0.00fF
C32797 NOR2X1_LOC_360/Y NOR2X1_LOC_211/A 0.01fF
C32798 NOR2X1_LOC_227/a_36_216# INVX1_LOC_75/A 0.00fF
C32799 NAND2X1_LOC_860/A INVX1_LOC_304/A 1.18fF
C32800 INVX1_LOC_136/A NOR2X1_LOC_781/A 0.12fF
C32801 NOR2X1_LOC_45/B NOR2X1_LOC_109/Y 0.23fF
C32802 INVX1_LOC_278/A NAND2X1_LOC_642/Y 0.01fF
C32803 NOR2X1_LOC_829/Y VDD 0.51fF
C32804 INVX1_LOC_155/A NAND2X1_LOC_675/a_36_24# 0.00fF
C32805 NOR2X1_LOC_738/A NOR2X1_LOC_307/A 0.06fF
C32806 NOR2X1_LOC_718/B INVX1_LOC_85/A 0.04fF
C32807 INVX1_LOC_204/A VDD 0.24fF
C32808 NOR2X1_LOC_68/A GATE_662 0.01fF
C32809 INVX1_LOC_292/A INVX1_LOC_313/Y 0.30fF
C32810 NOR2X1_LOC_613/Y INVX1_LOC_6/A 0.06fF
C32811 NAND2X1_LOC_765/a_36_24# NOR2X1_LOC_770/B 0.02fF
C32812 NOR2X1_LOC_860/Y NOR2X1_LOC_38/B 0.00fF
C32813 INVX1_LOC_98/A NOR2X1_LOC_652/Y 0.05fF
C32814 NOR2X1_LOC_422/a_36_216# INVX1_LOC_209/Y 0.00fF
C32815 INVX1_LOC_24/A NOR2X1_LOC_748/Y 0.03fF
C32816 NOR2X1_LOC_82/A INVX1_LOC_102/Y 0.00fF
C32817 NOR2X1_LOC_78/B NOR2X1_LOC_344/A 0.03fF
C32818 NOR2X1_LOC_78/A NOR2X1_LOC_652/Y 0.07fF
C32819 NAND2X1_LOC_55/a_36_24# NAND2X1_LOC_338/B 0.00fF
C32820 INVX1_LOC_88/A INPUT_0 0.03fF
C32821 INVX1_LOC_149/A INVX1_LOC_104/A 0.07fF
C32822 NAND2X1_LOC_364/A NAND2X1_LOC_656/Y 0.03fF
C32823 NOR2X1_LOC_495/Y INVX1_LOC_16/A 0.03fF
C32824 NOR2X1_LOC_447/Y INVX1_LOC_290/A 0.00fF
C32825 NAND2X1_LOC_337/B INVX1_LOC_75/A 0.06fF
C32826 NOR2X1_LOC_200/a_36_216# INVX1_LOC_266/Y 0.00fF
C32827 INVX1_LOC_124/A NOR2X1_LOC_709/A 0.06fF
C32828 NOR2X1_LOC_67/A NOR2X1_LOC_392/B 0.53fF
C32829 INVX1_LOC_136/A NOR2X1_LOC_76/A 0.07fF
C32830 INVX1_LOC_270/A INVX1_LOC_281/A 0.00fF
C32831 INVX1_LOC_89/A NOR2X1_LOC_554/B 0.07fF
C32832 INVX1_LOC_73/A NOR2X1_LOC_276/Y 0.02fF
C32833 NAND2X1_LOC_558/a_36_24# INVX1_LOC_309/A 0.00fF
C32834 NAND2X1_LOC_364/A INVX1_LOC_132/Y 0.11fF
C32835 NAND2X1_LOC_363/B NAND2X1_LOC_611/a_36_24# 0.00fF
C32836 INVX1_LOC_63/Y INVX1_LOC_22/A 0.08fF
C32837 NAND2X1_LOC_734/B NOR2X1_LOC_773/Y 0.02fF
C32838 NOR2X1_LOC_329/B INVX1_LOC_30/A 0.07fF
C32839 NAND2X1_LOC_350/A NOR2X1_LOC_815/A 0.04fF
C32840 INVX1_LOC_256/A INVX1_LOC_69/Y 0.10fF
C32841 INVX1_LOC_250/A INVX1_LOC_28/A 0.01fF
C32842 NOR2X1_LOC_114/Y INVX1_LOC_19/A 0.00fF
C32843 NAND2X1_LOC_508/A NOR2X1_LOC_554/B 0.46fF
C32844 NOR2X1_LOC_175/B NOR2X1_LOC_175/A 0.01fF
C32845 INVX1_LOC_93/A INVX1_LOC_20/A 0.08fF
C32846 D_INPUT_4 INVX1_LOC_30/A 0.00fF
C32847 NOR2X1_LOC_445/Y NOR2X1_LOC_543/A 0.01fF
C32848 NOR2X1_LOC_332/A NOR2X1_LOC_554/a_36_216# 0.01fF
C32849 INVX1_LOC_171/A NOR2X1_LOC_303/Y 0.15fF
C32850 NOR2X1_LOC_654/A INVX1_LOC_54/A 0.02fF
C32851 NOR2X1_LOC_137/Y NOR2X1_LOC_674/Y 0.01fF
C32852 INVX1_LOC_77/A NOR2X1_LOC_106/A 0.03fF
C32853 NAND2X1_LOC_276/Y INVX1_LOC_7/A 0.03fF
C32854 NAND2X1_LOC_763/B D_INPUT_4 0.02fF
C32855 INVX1_LOC_207/A NOR2X1_LOC_299/Y 0.07fF
C32856 INVX1_LOC_136/A INVX1_LOC_73/A 0.03fF
C32857 NOR2X1_LOC_175/A INVX1_LOC_22/A 0.39fF
C32858 NOR2X1_LOC_619/A NOR2X1_LOC_720/a_36_216# 0.00fF
C32859 NAND2X1_LOC_739/a_36_24# NAND2X1_LOC_800/A 0.00fF
C32860 NOR2X1_LOC_717/B NOR2X1_LOC_570/B 0.35fF
C32861 INVX1_LOC_178/A NAND2X1_LOC_453/A 0.10fF
C32862 INPUT_0 NOR2X1_LOC_500/B 0.15fF
C32863 D_INPUT_3 INVX1_LOC_252/A 0.01fF
C32864 INVX1_LOC_90/A NOR2X1_LOC_753/Y 0.03fF
C32865 NOR2X1_LOC_570/A INVX1_LOC_177/A 0.01fF
C32866 NAND2X1_LOC_367/A NAND2X1_LOC_366/a_36_24# 0.00fF
C32867 NAND2X1_LOC_833/Y NAND2X1_LOC_862/Y 0.05fF
C32868 INVX1_LOC_49/A NOR2X1_LOC_356/A 0.08fF
C32869 NOR2X1_LOC_773/Y INVX1_LOC_25/Y 0.10fF
C32870 INVX1_LOC_90/A NOR2X1_LOC_520/B 0.07fF
C32871 NOR2X1_LOC_788/B INVX1_LOC_33/A 0.03fF
C32872 INVX1_LOC_90/A NAND2X1_LOC_325/Y 0.03fF
C32873 NAND2X1_LOC_255/a_36_24# NOR2X1_LOC_748/A 0.00fF
C32874 INVX1_LOC_2/A NOR2X1_LOC_171/a_36_216# 0.00fF
C32875 NOR2X1_LOC_52/Y INVX1_LOC_6/A 0.00fF
C32876 NOR2X1_LOC_708/Y NAND2X1_LOC_696/a_36_24# 0.00fF
C32877 INVX1_LOC_124/Y NOR2X1_LOC_191/a_36_216# 0.00fF
C32878 NOR2X1_LOC_270/Y INVX1_LOC_6/A 0.04fF
C32879 NOR2X1_LOC_735/Y INVX1_LOC_63/Y 0.01fF
C32880 INVX1_LOC_118/A INVX1_LOC_306/Y 0.27fF
C32881 INVX1_LOC_13/A INVX1_LOC_226/Y 1.83fF
C32882 NAND2X1_LOC_722/A NOR2X1_LOC_380/A 0.39fF
C32883 NOR2X1_LOC_846/B NOR2X1_LOC_87/B 0.00fF
C32884 INVX1_LOC_36/A NOR2X1_LOC_45/B 3.78fF
C32885 NOR2X1_LOC_521/Y INVX1_LOC_172/Y 0.24fF
C32886 INVX1_LOC_41/A NOR2X1_LOC_567/B 0.07fF
C32887 INVX1_LOC_54/Y INVX1_LOC_171/A 0.03fF
C32888 INVX1_LOC_222/A NOR2X1_LOC_303/Y 0.10fF
C32889 INVX1_LOC_12/A NOR2X1_LOC_158/Y 0.07fF
C32890 INVX1_LOC_303/A INPUT_0 0.07fF
C32891 INVX1_LOC_305/A INVX1_LOC_186/A 0.07fF
C32892 INVX1_LOC_49/A NOR2X1_LOC_74/A 1.03fF
C32893 NAND2X1_LOC_740/B NAND2X1_LOC_354/B 0.55fF
C32894 NOR2X1_LOC_334/Y INVX1_LOC_290/Y 0.01fF
C32895 NOR2X1_LOC_151/Y NOR2X1_LOC_570/B 0.02fF
C32896 INVX1_LOC_276/A INVX1_LOC_90/A 0.72fF
C32897 NOR2X1_LOC_304/Y NAND2X1_LOC_802/Y 0.02fF
C32898 INVX1_LOC_136/A NAND2X1_LOC_729/B 0.01fF
C32899 INVX1_LOC_2/A NOR2X1_LOC_356/A 0.03fF
C32900 NAND2X1_LOC_323/B INVX1_LOC_120/A 0.00fF
C32901 NAND2X1_LOC_352/B INVX1_LOC_46/A 0.03fF
C32902 INVX1_LOC_49/A NOR2X1_LOC_9/Y 0.07fF
C32903 INVX1_LOC_173/Y NOR2X1_LOC_505/Y 0.08fF
C32904 INVX1_LOC_36/A INVX1_LOC_247/A 0.96fF
C32905 NOR2X1_LOC_67/A INVX1_LOC_90/A 0.07fF
C32906 NAND2X1_LOC_219/B NAND2X1_LOC_215/A 0.01fF
C32907 INVX1_LOC_238/A VDD 0.19fF
C32908 NOR2X1_LOC_721/Y INVX1_LOC_8/A 0.46fF
C32909 NOR2X1_LOC_488/a_36_216# INVX1_LOC_90/A 0.00fF
C32910 NOR2X1_LOC_716/B INVX1_LOC_286/A 0.19fF
C32911 INVX1_LOC_45/A INVX1_LOC_176/A 0.03fF
C32912 INVX1_LOC_35/A NAND2X1_LOC_475/Y 0.01fF
C32913 INVX1_LOC_33/A NOR2X1_LOC_147/A 0.04fF
C32914 INVX1_LOC_11/A NOR2X1_LOC_536/A 0.40fF
C32915 NOR2X1_LOC_510/Y NOR2X1_LOC_58/Y 0.01fF
C32916 INVX1_LOC_124/Y NOR2X1_LOC_266/B 0.19fF
C32917 INVX1_LOC_89/A NAND2X1_LOC_859/B 0.01fF
C32918 NOR2X1_LOC_15/Y NOR2X1_LOC_612/Y 0.02fF
C32919 D_INPUT_0 NAND2X1_LOC_660/Y 0.01fF
C32920 INVX1_LOC_55/Y NOR2X1_LOC_500/Y 0.08fF
C32921 NOR2X1_LOC_237/Y NOR2X1_LOC_45/B 0.19fF
C32922 INVX1_LOC_280/Y NAND2X1_LOC_560/A 0.03fF
C32923 NAND2X1_LOC_733/B NOR2X1_LOC_380/Y 0.17fF
C32924 INVX1_LOC_282/Y NAND2X1_LOC_463/B 3.76fF
C32925 NAND2X1_LOC_721/B VDD 0.13fF
C32926 INVX1_LOC_103/A NOR2X1_LOC_506/Y 0.02fF
C32927 INVX1_LOC_72/A NOR2X1_LOC_137/Y 0.03fF
C32928 NOR2X1_LOC_391/A NOR2X1_LOC_71/Y 0.16fF
C32929 NOR2X1_LOC_690/A NOR2X1_LOC_526/a_36_216# 0.01fF
C32930 NOR2X1_LOC_590/A INVX1_LOC_44/A 0.39fF
C32931 INVX1_LOC_2/A NOR2X1_LOC_74/A 0.32fF
C32932 NOR2X1_LOC_67/A NAND2X1_LOC_348/A 0.00fF
C32933 NAND2X1_LOC_634/Y VDD 0.82fF
C32934 NOR2X1_LOC_561/Y NOR2X1_LOC_510/a_36_216# 0.01fF
C32935 D_INPUT_7 INVX1_LOC_37/A 0.01fF
C32936 INVX1_LOC_247/Y VDD 0.47fF
C32937 NOR2X1_LOC_598/B NOR2X1_LOC_830/Y 0.04fF
C32938 NOR2X1_LOC_48/B NOR2X1_LOC_654/A 0.11fF
C32939 INVX1_LOC_54/Y INVX1_LOC_222/A 0.01fF
C32940 NOR2X1_LOC_773/Y INVX1_LOC_75/A 0.07fF
C32941 INVX1_LOC_140/A INVX1_LOC_25/Y 0.07fF
C32942 NOR2X1_LOC_75/Y INVX1_LOC_54/A 0.04fF
C32943 NOR2X1_LOC_226/A NOR2X1_LOC_74/A 0.50fF
C32944 NAND2X1_LOC_556/a_36_24# INVX1_LOC_309/A 0.00fF
C32945 INVX1_LOC_2/A NOR2X1_LOC_9/Y 0.10fF
C32946 NOR2X1_LOC_716/B INVX1_LOC_95/A 0.02fF
C32947 NOR2X1_LOC_205/Y NOR2X1_LOC_155/A 0.03fF
C32948 NOR2X1_LOC_647/A NOR2X1_LOC_38/B 0.00fF
C32949 INVX1_LOC_11/A NAND2X1_LOC_93/B 0.06fF
C32950 NOR2X1_LOC_278/Y INVX1_LOC_94/Y 0.00fF
C32951 NOR2X1_LOC_309/Y NOR2X1_LOC_45/B 0.07fF
C32952 INVX1_LOC_302/Y INVX1_LOC_22/A 0.01fF
C32953 NOR2X1_LOC_220/A NOR2X1_LOC_548/A 0.03fF
C32954 INVX1_LOC_228/A VDD 0.12fF
C32955 INVX1_LOC_290/A INVX1_LOC_302/A 0.03fF
C32956 NOR2X1_LOC_226/A NOR2X1_LOC_9/Y 0.51fF
C32957 INVX1_LOC_239/A INVX1_LOC_84/A 0.01fF
C32958 INVX1_LOC_21/A NAND2X1_LOC_782/B 0.25fF
C32959 NOR2X1_LOC_590/A NOR2X1_LOC_641/Y 0.00fF
C32960 NOR2X1_LOC_392/Y INVX1_LOC_42/A 0.01fF
C32961 INVX1_LOC_11/A NAND2X1_LOC_425/Y 0.14fF
C32962 NAND2X1_LOC_573/a_36_24# INVX1_LOC_46/A 0.00fF
C32963 NAND2X1_LOC_361/Y NOR2X1_LOC_35/Y 0.10fF
C32964 NOR2X1_LOC_559/a_36_216# NOR2X1_LOC_560/A 0.02fF
C32965 INVX1_LOC_163/A INVX1_LOC_203/A 0.03fF
C32966 NOR2X1_LOC_510/Y INVX1_LOC_29/A 0.07fF
C32967 NAND2X1_LOC_350/A NAND2X1_LOC_436/a_36_24# 0.02fF
C32968 INVX1_LOC_43/Y NOR2X1_LOC_216/B 0.01fF
C32969 NAND2X1_LOC_276/Y INVX1_LOC_76/A 0.07fF
C32970 NAND2X1_LOC_222/B INVX1_LOC_3/A 0.11fF
C32971 NOR2X1_LOC_528/Y NAND2X1_LOC_850/Y 0.06fF
C32972 NOR2X1_LOC_16/Y NAND2X1_LOC_642/Y 0.01fF
C32973 NOR2X1_LOC_68/A NOR2X1_LOC_261/A 0.03fF
C32974 NOR2X1_LOC_548/A NOR2X1_LOC_548/Y 0.12fF
C32975 INVX1_LOC_11/A NOR2X1_LOC_649/B 0.00fF
C32976 NOR2X1_LOC_208/Y INVX1_LOC_281/A 0.00fF
C32977 NOR2X1_LOC_543/A NOR2X1_LOC_335/B 0.01fF
C32978 INVX1_LOC_5/A INVX1_LOC_283/A 0.04fF
C32979 NOR2X1_LOC_639/B NOR2X1_LOC_467/A 0.04fF
C32980 NOR2X1_LOC_332/A INVX1_LOC_75/A 0.07fF
C32981 NAND2X1_LOC_381/Y NOR2X1_LOC_649/B 0.02fF
C32982 INVX1_LOC_80/A INPUT_0 0.01fF
C32983 INVX1_LOC_98/Y INVX1_LOC_95/A 0.01fF
C32984 NOR2X1_LOC_550/B INVX1_LOC_117/A 0.10fF
C32985 VDD INVX1_LOC_8/A 1.71fF
C32986 NOR2X1_LOC_433/A NOR2X1_LOC_536/A 0.06fF
C32987 NOR2X1_LOC_296/a_36_216# NAND2X1_LOC_773/B 0.01fF
C32988 NAND2X1_LOC_357/B INVX1_LOC_46/A 0.07fF
C32989 NOR2X1_LOC_348/Y NOR2X1_LOC_89/A 0.16fF
C32990 NOR2X1_LOC_753/Y INVX1_LOC_38/A 0.07fF
C32991 NOR2X1_LOC_361/B INVX1_LOC_29/A 0.07fF
C32992 NOR2X1_LOC_473/B INVX1_LOC_67/Y 0.49fF
C32993 NOR2X1_LOC_168/B NOR2X1_LOC_857/A 0.06fF
C32994 INVX1_LOC_172/Y INVX1_LOC_255/A 0.01fF
C32995 NOR2X1_LOC_352/Y INVX1_LOC_76/A 0.01fF
C32996 NOR2X1_LOC_74/A INPUT_1 0.10fF
C32997 NOR2X1_LOC_520/B INVX1_LOC_38/A 0.03fF
C32998 NAND2X1_LOC_323/B INVX1_LOC_143/Y 0.03fF
C32999 NAND2X1_LOC_325/Y INVX1_LOC_38/A 0.12fF
C33000 NOR2X1_LOC_823/Y INVX1_LOC_22/A 0.01fF
C33001 INVX1_LOC_83/A NAND2X1_LOC_473/a_36_24# 0.01fF
C33002 NAND2X1_LOC_133/a_36_24# INVX1_LOC_48/A 0.01fF
C33003 NAND2X1_LOC_474/Y INVX1_LOC_32/A 0.10fF
C33004 NOR2X1_LOC_91/Y NOR2X1_LOC_88/Y 0.03fF
C33005 INVX1_LOC_311/A INVX1_LOC_85/Y 0.02fF
C33006 NAND2X1_LOC_332/Y NOR2X1_LOC_331/B 0.00fF
C33007 INVX1_LOC_61/A NAND2X1_LOC_243/a_36_24# 0.01fF
C33008 INPUT_1 NOR2X1_LOC_9/Y 0.33fF
C33009 NOR2X1_LOC_716/B INVX1_LOC_54/A 0.03fF
C33010 INVX1_LOC_239/A INVX1_LOC_15/A 0.01fF
C33011 NOR2X1_LOC_52/B NOR2X1_LOC_536/A 0.12fF
C33012 NOR2X1_LOC_852/Y NOR2X1_LOC_839/B 0.36fF
C33013 INVX1_LOC_68/Y INVX1_LOC_36/Y 0.26fF
C33014 INVX1_LOC_256/A NOR2X1_LOC_89/A 0.50fF
C33015 NAND2X1_LOC_838/Y NOR2X1_LOC_536/A 0.01fF
C33016 INVX1_LOC_211/Y INVX1_LOC_12/A 0.03fF
C33017 INVX1_LOC_24/A INVX1_LOC_123/Y 0.12fF
C33018 NAND2X1_LOC_773/Y INVX1_LOC_47/Y 0.10fF
C33019 NAND2X1_LOC_656/Y NOR2X1_LOC_405/A 0.08fF
C33020 INVX1_LOC_151/Y VDD 0.41fF
C33021 NOR2X1_LOC_91/Y INVX1_LOC_84/A 0.04fF
C33022 NAND2X1_LOC_479/Y INVX1_LOC_139/A 0.03fF
C33023 INVX1_LOC_34/A NOR2X1_LOC_99/Y 0.07fF
C33024 NOR2X1_LOC_804/B NOR2X1_LOC_862/B 0.02fF
C33025 INVX1_LOC_276/A INVX1_LOC_38/A 0.16fF
C33026 NOR2X1_LOC_709/A INVX1_LOC_9/A 0.03fF
C33027 INVX1_LOC_73/Y INVX1_LOC_15/A 0.04fF
C33028 NOR2X1_LOC_67/A NAND2X1_LOC_849/B 0.25fF
C33029 NAND2X1_LOC_53/Y INVX1_LOC_32/A 0.07fF
C33030 NOR2X1_LOC_122/Y NOR2X1_LOC_269/Y 0.00fF
C33031 INVX1_LOC_119/A INVX1_LOC_291/A 0.10fF
C33032 NOR2X1_LOC_828/B NAND2X1_LOC_682/a_36_24# 0.00fF
C33033 NOR2X1_LOC_717/B NAND2X1_LOC_454/a_36_24# 0.00fF
C33034 INVX1_LOC_21/A NOR2X1_LOC_831/a_36_216# 0.00fF
C33035 NAND2X1_LOC_317/a_36_24# NAND2X1_LOC_453/A 0.00fF
C33036 INVX1_LOC_40/A NAND2X1_LOC_297/a_36_24# 0.00fF
C33037 INVX1_LOC_35/A NAND2X1_LOC_363/B 0.03fF
C33038 NOR2X1_LOC_92/Y INVX1_LOC_26/A 0.06fF
C33039 NAND2X1_LOC_65/a_36_24# INVX1_LOC_27/A 0.00fF
C33040 NOR2X1_LOC_808/A INVX1_LOC_307/Y 0.23fF
C33041 NOR2X1_LOC_186/Y D_INPUT_1 0.03fF
C33042 INVX1_LOC_11/A NAND2X1_LOC_470/B 0.02fF
C33043 NOR2X1_LOC_757/A NOR2X1_LOC_363/Y 0.15fF
C33044 NOR2X1_LOC_188/A NOR2X1_LOC_501/B 0.03fF
C33045 INVX1_LOC_233/Y NAND2X1_LOC_725/A 0.10fF
C33046 NAND2X1_LOC_140/A VDD 0.29fF
C33047 INVX1_LOC_45/A NOR2X1_LOC_116/a_36_216# -0.00fF
C33048 INVX1_LOC_77/A NAND2X1_LOC_781/a_36_24# 0.01fF
C33049 INVX1_LOC_135/A NAND2X1_LOC_721/A 0.01fF
C33050 INVX1_LOC_64/A INVX1_LOC_99/Y 0.05fF
C33051 NOR2X1_LOC_604/a_36_216# INVX1_LOC_27/A 0.01fF
C33052 NOR2X1_LOC_68/A NOR2X1_LOC_147/a_36_216# 0.00fF
C33053 INVX1_LOC_233/A NAND2X1_LOC_169/Y 0.01fF
C33054 NOR2X1_LOC_631/B NOR2X1_LOC_197/Y 0.03fF
C33055 INVX1_LOC_313/Y NOR2X1_LOC_137/Y 0.11fF
C33056 INVX1_LOC_35/A NOR2X1_LOC_840/A 0.04fF
C33057 INVX1_LOC_14/A NAND2X1_LOC_442/a_36_24# 0.00fF
C33058 NOR2X1_LOC_690/A NOR2X1_LOC_662/A 0.08fF
C33059 INVX1_LOC_24/A INVX1_LOC_102/A 0.07fF
C33060 NAND2X1_LOC_9/Y NOR2X1_LOC_789/B 0.04fF
C33061 NOR2X1_LOC_447/Y INVX1_LOC_261/Y 0.00fF
C33062 NAND2X1_LOC_564/A NOR2X1_LOC_92/Y 0.02fF
C33063 NAND2X1_LOC_662/Y NAND2X1_LOC_637/Y 0.07fF
C33064 INVX1_LOC_63/Y INVX1_LOC_186/Y 0.10fF
C33065 INVX1_LOC_236/Y INVX1_LOC_94/Y 0.00fF
C33066 INVX1_LOC_51/Y NAND2X1_LOC_86/Y 0.04fF
C33067 INVX1_LOC_266/Y NOR2X1_LOC_66/Y 0.00fF
C33068 D_INPUT_0 NAND2X1_LOC_848/A 0.13fF
C33069 INVX1_LOC_69/Y NOR2X1_LOC_543/a_36_216# 0.01fF
C33070 NAND2X1_LOC_784/A NAND2X1_LOC_579/A 0.02fF
C33071 NOR2X1_LOC_655/B NAND2X1_LOC_572/B 0.03fF
C33072 NAND2X1_LOC_860/A NAND2X1_LOC_634/a_36_24# 0.00fF
C33073 NOR2X1_LOC_91/Y INVX1_LOC_15/A 0.03fF
C33074 INVX1_LOC_140/A NAND2X1_LOC_453/A 0.10fF
C33075 NOR2X1_LOC_202/Y INVX1_LOC_139/A 0.01fF
C33076 NOR2X1_LOC_824/A NAND2X1_LOC_624/B 0.03fF
C33077 NAND2X1_LOC_733/Y NOR2X1_LOC_25/Y 0.05fF
C33078 NOR2X1_LOC_473/B NOR2X1_LOC_366/a_36_216# 0.00fF
C33079 INVX1_LOC_13/Y NOR2X1_LOC_220/B 0.03fF
C33080 INVX1_LOC_71/A NOR2X1_LOC_116/a_36_216# 0.01fF
C33081 NOR2X1_LOC_186/Y NOR2X1_LOC_652/Y 1.21fF
C33082 INVX1_LOC_36/A NOR2X1_LOC_465/Y 0.03fF
C33083 NOR2X1_LOC_106/A INVX1_LOC_9/A 0.33fF
C33084 INVX1_LOC_39/A INVX1_LOC_306/Y 0.04fF
C33085 NOR2X1_LOC_219/B INVX1_LOC_109/Y 0.03fF
C33086 NOR2X1_LOC_742/A INVX1_LOC_139/Y 0.02fF
C33087 NAND2X1_LOC_350/A NOR2X1_LOC_654/A 0.04fF
C33088 NOR2X1_LOC_160/B NOR2X1_LOC_383/B 0.13fF
C33089 INVX1_LOC_27/A NOR2X1_LOC_849/A 0.06fF
C33090 INVX1_LOC_248/Y NAND2X1_LOC_714/B 0.01fF
C33091 NOR2X1_LOC_318/B NOR2X1_LOC_552/A 0.04fF
C33092 INVX1_LOC_208/A NOR2X1_LOC_127/Y 0.02fF
C33093 INVX1_LOC_6/A NOR2X1_LOC_603/Y 0.02fF
C33094 NOR2X1_LOC_785/Y NOR2X1_LOC_634/A 0.31fF
C33095 NOR2X1_LOC_303/Y INVX1_LOC_4/A 0.17fF
C33096 INVX1_LOC_177/A INVX1_LOC_29/A 0.09fF
C33097 NAND2X1_LOC_33/Y INVX1_LOC_42/A 0.03fF
C33098 NAND2X1_LOC_231/Y INVX1_LOC_272/A 0.10fF
C33099 D_INPUT_0 INVX1_LOC_46/Y 0.19fF
C33100 INVX1_LOC_226/Y NAND2X1_LOC_489/Y 0.02fF
C33101 NOR2X1_LOC_544/A INVX1_LOC_19/A 0.08fF
C33102 INVX1_LOC_193/Y NOR2X1_LOC_706/B 0.00fF
C33103 INVX1_LOC_286/A NAND2X1_LOC_633/Y 0.10fF
C33104 INVX1_LOC_6/A NOR2X1_LOC_139/a_36_216# 0.00fF
C33105 INVX1_LOC_49/A NOR2X1_LOC_855/A 0.03fF
C33106 INVX1_LOC_77/A NOR2X1_LOC_334/Y 0.14fF
C33107 NOR2X1_LOC_135/Y NOR2X1_LOC_351/Y 0.01fF
C33108 NAND2X1_LOC_549/B NOR2X1_LOC_671/Y 0.01fF
C33109 NOR2X1_LOC_543/A INVX1_LOC_84/A 0.06fF
C33110 NAND2X1_LOC_181/Y NAND2X1_LOC_74/B 0.04fF
C33111 NOR2X1_LOC_596/a_36_216# NAND2X1_LOC_454/Y 0.03fF
C33112 D_INPUT_1 INVX1_LOC_170/A 0.06fF
C33113 INVX1_LOC_17/A INVX1_LOC_50/Y 0.07fF
C33114 INVX1_LOC_55/Y INVX1_LOC_307/A 0.07fF
C33115 NOR2X1_LOC_334/A INVX1_LOC_117/A 0.02fF
C33116 NOR2X1_LOC_562/B NOR2X1_LOC_562/A 0.12fF
C33117 NOR2X1_LOC_270/Y INVX1_LOC_270/A 0.19fF
C33118 NAND2X1_LOC_366/a_36_24# NOR2X1_LOC_865/Y 0.00fF
C33119 NOR2X1_LOC_373/a_36_216# INVX1_LOC_78/A 0.00fF
C33120 NOR2X1_LOC_703/B INVX1_LOC_23/A 0.03fF
C33121 NAND2X1_LOC_842/B NOR2X1_LOC_831/B 0.07fF
C33122 NOR2X1_LOC_74/A INVX1_LOC_118/A 0.07fF
C33123 INVX1_LOC_35/A INVX1_LOC_30/A 1.16fF
C33124 INVX1_LOC_95/A NAND2X1_LOC_633/Y 0.00fF
C33125 INVX1_LOC_24/A INVX1_LOC_296/Y 0.03fF
C33126 INVX1_LOC_49/A NAND2X1_LOC_425/a_36_24# 0.01fF
C33127 NOR2X1_LOC_716/B NOR2X1_LOC_438/Y 0.04fF
C33128 INVX1_LOC_25/Y INVX1_LOC_42/A 0.26fF
C33129 INVX1_LOC_58/A NOR2X1_LOC_273/Y 0.03fF
C33130 NAND2X1_LOC_364/A NOR2X1_LOC_717/A 0.05fF
C33131 INVX1_LOC_54/Y INVX1_LOC_4/A 0.10fF
C33132 NOR2X1_LOC_320/a_36_216# INVX1_LOC_78/A 0.00fF
C33133 NAND2X1_LOC_357/B NOR2X1_LOC_282/a_36_216# 0.00fF
C33134 INVX1_LOC_286/A NOR2X1_LOC_709/B 0.03fF
C33135 INVX1_LOC_36/A NOR2X1_LOC_53/Y 0.01fF
C33136 INVX1_LOC_41/A INVX1_LOC_26/A 4.82fF
C33137 INVX1_LOC_58/A NOR2X1_LOC_759/Y 0.17fF
C33138 NOR2X1_LOC_299/Y NOR2X1_LOC_36/B 0.01fF
C33139 INVX1_LOC_162/A NOR2X1_LOC_278/Y 0.07fF
C33140 NAND2X1_LOC_573/A INVX1_LOC_29/A 0.10fF
C33141 INVX1_LOC_93/Y NOR2X1_LOC_558/a_36_216# 0.01fF
C33142 INVX1_LOC_254/A INVX1_LOC_57/A 0.02fF
C33143 INVX1_LOC_278/A NOR2X1_LOC_91/Y 0.06fF
C33144 INVX1_LOC_305/A NAND2X1_LOC_431/a_36_24# 0.01fF
C33145 NOR2X1_LOC_440/Y NOR2X1_LOC_89/A 0.01fF
C33146 NAND2X1_LOC_593/Y INVX1_LOC_271/A 0.01fF
C33147 NOR2X1_LOC_802/A NAND2X1_LOC_72/B 0.01fF
C33148 NOR2X1_LOC_468/Y NAND2X1_LOC_793/Y 0.02fF
C33149 NOR2X1_LOC_569/Y INVX1_LOC_290/Y 0.01fF
C33150 NOR2X1_LOC_500/Y INVX1_LOC_32/A 0.07fF
C33151 INVX1_LOC_226/Y INVX1_LOC_32/A 0.14fF
C33152 NOR2X1_LOC_837/B NAND2X1_LOC_363/B 0.02fF
C33153 INVX1_LOC_35/A NOR2X1_LOC_705/a_36_216# 0.00fF
C33154 NOR2X1_LOC_317/B NOR2X1_LOC_383/B 0.03fF
C33155 NOR2X1_LOC_322/Y INVX1_LOC_285/A 0.29fF
C33156 NOR2X1_LOC_332/A NAND2X1_LOC_291/B 0.11fF
C33157 INVX1_LOC_298/Y INVX1_LOC_177/A 0.03fF
C33158 NOR2X1_LOC_474/A NOR2X1_LOC_476/B 0.48fF
C33159 INVX1_LOC_240/A NAND2X1_LOC_402/B 0.04fF
C33160 NOR2X1_LOC_67/A NAND2X1_LOC_223/A 0.12fF
C33161 NOR2X1_LOC_481/A D_INPUT_1 0.08fF
C33162 NOR2X1_LOC_690/A INVX1_LOC_57/A 3.91fF
C33163 INVX1_LOC_256/A INVX1_LOC_11/A 0.22fF
C33164 NOR2X1_LOC_130/A INVX1_LOC_102/A 0.07fF
C33165 INVX1_LOC_64/A NOR2X1_LOC_303/Y 0.03fF
C33166 INVX1_LOC_42/Y NOR2X1_LOC_66/Y 0.02fF
C33167 INVX1_LOC_13/Y INVX1_LOC_72/Y 0.02fF
C33168 NOR2X1_LOC_859/A INVX1_LOC_27/A 0.03fF
C33169 NOR2X1_LOC_413/Y INVX1_LOC_57/A 0.01fF
C33170 NOR2X1_LOC_741/A INVX1_LOC_179/A 0.01fF
C33171 INVX1_LOC_33/Y NOR2X1_LOC_305/Y 0.00fF
C33172 INVX1_LOC_36/Y NOR2X1_LOC_115/a_36_216# 0.00fF
C33173 INVX1_LOC_85/Y NOR2X1_LOC_307/a_36_216# 0.00fF
C33174 NOR2X1_LOC_760/a_36_216# INVX1_LOC_161/Y 0.01fF
C33175 NAND2X1_LOC_218/B INVX1_LOC_5/A 0.03fF
C33176 INVX1_LOC_21/A NOR2X1_LOC_68/A 0.38fF
C33177 NOR2X1_LOC_45/B NOR2X1_LOC_435/A 0.03fF
C33178 D_INPUT_1 INVX1_LOC_225/A 0.56fF
C33179 INVX1_LOC_55/Y INVX1_LOC_12/A 0.03fF
C33180 NOR2X1_LOC_558/A NOR2X1_LOC_561/A 0.08fF
C33181 INVX1_LOC_58/A INVX1_LOC_249/Y 0.04fF
C33182 NOR2X1_LOC_687/Y NOR2X1_LOC_334/Y 0.07fF
C33183 INVX1_LOC_10/A INVX1_LOC_32/A 0.07fF
C33184 INVX1_LOC_25/Y INVX1_LOC_78/A 0.12fF
C33185 INVX1_LOC_292/A NOR2X1_LOC_541/Y 0.01fF
C33186 INVX1_LOC_90/A NAND2X1_LOC_807/a_36_24# 0.00fF
C33187 NAND2X1_LOC_721/A NOR2X1_LOC_813/Y 0.00fF
C33188 NOR2X1_LOC_446/A INVX1_LOC_188/A 0.11fF
C33189 INVX1_LOC_45/A INVX1_LOC_103/A 0.07fF
C33190 NOR2X1_LOC_464/a_36_216# NOR2X1_LOC_678/A 0.00fF
C33191 NAND2X1_LOC_35/Y INVX1_LOC_207/A 0.08fF
C33192 INVX1_LOC_64/A NOR2X1_LOC_254/Y 0.04fF
C33193 NAND2X1_LOC_200/B NOR2X1_LOC_720/A 0.01fF
C33194 NOR2X1_LOC_689/A NAND2X1_LOC_853/Y 0.12fF
C33195 VDD INVX1_LOC_118/Y 0.58fF
C33196 INVX1_LOC_58/A NOR2X1_LOC_41/Y 0.01fF
C33197 NAND2X1_LOC_721/A INVX1_LOC_280/A 0.02fF
C33198 NOR2X1_LOC_617/Y NOR2X1_LOC_824/A -0.11fF
C33199 NOR2X1_LOC_533/Y INVX1_LOC_72/A 0.42fF
C33200 NOR2X1_LOC_74/A NAND2X1_LOC_63/Y 0.01fF
C33201 NOR2X1_LOC_496/Y INVX1_LOC_172/A 0.01fF
C33202 NAND2X1_LOC_578/B INVX1_LOC_23/A 0.04fF
C33203 NAND2X1_LOC_363/B NAND2X1_LOC_667/a_36_24# 0.00fF
C33204 INPUT_0 INVX1_LOC_272/A 0.07fF
C33205 NOR2X1_LOC_65/B INVX1_LOC_25/Y 0.01fF
C33206 NAND2X1_LOC_633/Y INVX1_LOC_54/A 0.34fF
C33207 INVX1_LOC_208/A NOR2X1_LOC_383/B 2.00fF
C33208 NOR2X1_LOC_644/B NAND2X1_LOC_597/a_36_24# 0.02fF
C33209 NOR2X1_LOC_503/A NOR2X1_LOC_48/B 0.01fF
C33210 NAND2X1_LOC_392/A INVX1_LOC_181/A 0.01fF
C33211 INVX1_LOC_75/A NOR2X1_LOC_847/A 0.05fF
C33212 INVX1_LOC_178/A NOR2X1_LOC_577/Y 0.10fF
C33213 INVX1_LOC_57/Y NAND2X1_LOC_550/A -0.02fF
C33214 INVX1_LOC_10/A NAND2X1_LOC_175/Y 0.07fF
C33215 NOR2X1_LOC_516/B NOR2X1_LOC_383/B 0.03fF
C33216 INVX1_LOC_5/A NOR2X1_LOC_629/B 0.02fF
C33217 INVX1_LOC_45/A INVX1_LOC_292/A 0.08fF
C33218 NOR2X1_LOC_65/B NAND2X1_LOC_349/B 0.25fF
C33219 INVX1_LOC_269/A INVX1_LOC_45/Y 0.13fF
C33220 INVX1_LOC_75/A INVX1_LOC_42/A 0.14fF
C33221 NOR2X1_LOC_9/Y NAND2X1_LOC_63/Y 0.08fF
C33222 INVX1_LOC_10/A NOR2X1_LOC_821/a_36_216# 0.00fF
C33223 NOR2X1_LOC_391/A INVX1_LOC_16/Y 0.10fF
C33224 INVX1_LOC_33/Y NAND2X1_LOC_600/a_36_24# 0.00fF
C33225 NOR2X1_LOC_45/B INVX1_LOC_63/A 0.10fF
C33226 NAND2X1_LOC_738/B NAND2X1_LOC_853/Y 0.07fF
C33227 INVX1_LOC_285/Y INVX1_LOC_29/A 0.02fF
C33228 NAND2X1_LOC_724/Y NAND2X1_LOC_863/B 0.27fF
C33229 INVX1_LOC_50/A INVX1_LOC_16/A 0.22fF
C33230 NOR2X1_LOC_576/B NOR2X1_LOC_409/B 0.02fF
C33231 INVX1_LOC_229/Y NOR2X1_LOC_829/A 0.23fF
C33232 INVX1_LOC_225/A NOR2X1_LOC_652/Y 0.11fF
C33233 INVX1_LOC_35/Y INVX1_LOC_20/A 0.02fF
C33234 NAND2X1_LOC_579/A NOR2X1_LOC_625/Y 0.05fF
C33235 INPUT_0 NOR2X1_LOC_76/B 0.00fF
C33236 INVX1_LOC_135/A INVX1_LOC_175/A 0.09fF
C33237 NOR2X1_LOC_532/Y NAND2X1_LOC_72/B 0.07fF
C33238 INVX1_LOC_59/A NAND2X1_LOC_549/a_36_24# 0.00fF
C33239 INVX1_LOC_48/A NAND2X1_LOC_207/B 0.03fF
C33240 INVX1_LOC_103/A INVX1_LOC_71/A 0.07fF
C33241 INVX1_LOC_69/Y NOR2X1_LOC_89/A 0.07fF
C33242 INVX1_LOC_74/A NOR2X1_LOC_649/B 0.02fF
C33243 NAND2X1_LOC_725/A NOR2X1_LOC_526/Y 0.04fF
C33244 INVX1_LOC_74/A INVX1_LOC_3/A 0.14fF
C33245 INVX1_LOC_247/A INVX1_LOC_63/A 0.03fF
C33246 NAND2X1_LOC_859/B NOR2X1_LOC_392/Y 0.00fF
C33247 NOR2X1_LOC_793/Y INVX1_LOC_33/A 0.01fF
C33248 INVX1_LOC_5/A NOR2X1_LOC_346/B 4.83fF
C33249 NOR2X1_LOC_224/Y INVX1_LOC_16/A 0.06fF
C33250 NOR2X1_LOC_250/Y INVX1_LOC_49/A 0.09fF
C33251 NAND2X1_LOC_703/Y NAND2X1_LOC_357/B 0.03fF
C33252 NAND2X1_LOC_93/B NOR2X1_LOC_376/Y 0.08fF
C33253 INVX1_LOC_256/A NOR2X1_LOC_433/A 0.30fF
C33254 NOR2X1_LOC_91/A INVX1_LOC_183/Y 0.01fF
C33255 INVX1_LOC_292/A INVX1_LOC_71/A 0.07fF
C33256 NAND2X1_LOC_468/B INVX1_LOC_19/A 0.03fF
C33257 NOR2X1_LOC_361/B INVX1_LOC_8/A 0.10fF
C33258 INVX1_LOC_65/A INVX1_LOC_29/A 0.30fF
C33259 INVX1_LOC_93/A NAND2X1_LOC_850/Y 0.87fF
C33260 INVX1_LOC_245/Y INVX1_LOC_49/A 0.05fF
C33261 INVX1_LOC_36/A NOR2X1_LOC_270/Y 0.01fF
C33262 INVX1_LOC_13/Y NAND2X1_LOC_334/a_36_24# 0.00fF
C33263 INVX1_LOC_254/Y NAND2X1_LOC_114/B 0.01fF
C33264 INVX1_LOC_234/A NOR2X1_LOC_629/A 0.04fF
C33265 INVX1_LOC_69/Y NOR2X1_LOC_170/A 0.03fF
C33266 NOR2X1_LOC_816/A NOR2X1_LOC_577/Y 0.64fF
C33267 NOR2X1_LOC_865/A NOR2X1_LOC_862/B 0.32fF
C33268 INVX1_LOC_256/A NOR2X1_LOC_593/Y 0.01fF
C33269 INVX1_LOC_75/A INVX1_LOC_78/A 0.19fF
C33270 INVX1_LOC_218/Y NOR2X1_LOC_419/Y 0.01fF
C33271 INVX1_LOC_5/A INVX1_LOC_22/A 0.17fF
C33272 NOR2X1_LOC_376/Y NAND2X1_LOC_425/Y 0.03fF
C33273 INVX1_LOC_223/A INVX1_LOC_24/A 0.03fF
C33274 INVX1_LOC_34/A INVX1_LOC_150/Y 0.07fF
C33275 NOR2X1_LOC_510/Y INVX1_LOC_151/Y 0.01fF
C33276 NOR2X1_LOC_403/B INVX1_LOC_170/A 0.00fF
C33277 INVX1_LOC_17/A NOR2X1_LOC_6/B 0.02fF
C33278 VDD NOR2X1_LOC_258/Y 0.11fF
C33279 INVX1_LOC_71/Y INVX1_LOC_54/A 0.11fF
C33280 NAND2X1_LOC_624/B INVX1_LOC_234/A 0.07fF
C33281 NOR2X1_LOC_710/A INVX1_LOC_33/A 0.01fF
C33282 NOR2X1_LOC_596/A NAND2X1_LOC_16/Y -0.00fF
C33283 NOR2X1_LOC_211/a_36_216# INVX1_LOC_171/A 0.00fF
C33284 INVX1_LOC_50/A INVX1_LOC_28/A 0.14fF
C33285 INVX1_LOC_124/Y INVX1_LOC_49/A 0.01fF
C33286 NAND2X1_LOC_550/A NAND2X1_LOC_706/a_36_24# 0.00fF
C33287 INVX1_LOC_256/A NOR2X1_LOC_52/B 1.93fF
C33288 INVX1_LOC_20/A NOR2X1_LOC_824/a_36_216# 0.02fF
C33289 INVX1_LOC_178/A INVX1_LOC_22/A 0.54fF
C33290 NOR2X1_LOC_307/A NOR2X1_LOC_731/A 0.00fF
C33291 INVX1_LOC_94/A NOR2X1_LOC_360/Y 0.01fF
C33292 NOR2X1_LOC_357/Y INVX1_LOC_12/A 0.46fF
C33293 NOR2X1_LOC_65/B INVX1_LOC_75/A 0.19fF
C33294 INVX1_LOC_83/A INVX1_LOC_213/A 0.10fF
C33295 NOR2X1_LOC_208/Y NOR2X1_LOC_270/Y 0.44fF
C33296 NAND2X1_LOC_555/Y NOR2X1_LOC_6/B 0.05fF
C33297 NOR2X1_LOC_684/Y NOR2X1_LOC_257/Y 0.01fF
C33298 NAND2X1_LOC_13/a_36_24# INVX1_LOC_143/A 0.01fF
C33299 INVX1_LOC_2/A INVX1_LOC_245/Y 0.03fF
C33300 NOR2X1_LOC_564/Y INVX1_LOC_53/A 0.00fF
C33301 INVX1_LOC_14/A INVX1_LOC_316/Y 0.02fF
C33302 NAND2X1_LOC_453/A INVX1_LOC_42/A 0.02fF
C33303 NOR2X1_LOC_2/Y INVX1_LOC_173/A 0.01fF
C33304 NAND2X1_LOC_74/B INVX1_LOC_117/A 0.17fF
C33305 INVX1_LOC_277/A INVX1_LOC_213/Y 0.02fF
C33306 INVX1_LOC_30/A NOR2X1_LOC_365/a_36_216# 0.00fF
C33307 NOR2X1_LOC_91/A INVX1_LOC_309/A 0.00fF
C33308 INVX1_LOC_79/A INVX1_LOC_23/A 0.07fF
C33309 INVX1_LOC_64/A NOR2X1_LOC_112/Y 0.02fF
C33310 INVX1_LOC_255/Y INVX1_LOC_269/A 3.16fF
C33311 INVX1_LOC_18/A INVX1_LOC_63/Y 0.09fF
C33312 NOR2X1_LOC_703/a_36_216# INVX1_LOC_177/A 0.00fF
C33313 NOR2X1_LOC_160/B NAND2X1_LOC_347/a_36_24# 0.00fF
C33314 NOR2X1_LOC_296/Y INVX1_LOC_226/Y 0.01fF
C33315 NAND2X1_LOC_624/B NOR2X1_LOC_19/B 0.03fF
C33316 INVX1_LOC_59/A INVX1_LOC_219/A 0.01fF
C33317 INVX1_LOC_233/Y NAND2X1_LOC_560/A 0.01fF
C33318 NOR2X1_LOC_147/A INVX1_LOC_275/Y 0.15fF
C33319 NOR2X1_LOC_772/Y INVX1_LOC_181/Y 0.20fF
C33320 NAND2X1_LOC_725/Y NOR2X1_LOC_387/A 0.03fF
C33321 INVX1_LOC_5/A NOR2X1_LOC_735/Y -0.01fF
C33322 INVX1_LOC_12/A NOR2X1_LOC_692/Y 0.01fF
C33323 INVX1_LOC_13/A INVX1_LOC_228/Y 0.00fF
C33324 NAND2X1_LOC_227/Y INVX1_LOC_16/A 0.01fF
C33325 INVX1_LOC_11/A NOR2X1_LOC_397/a_36_216# 0.02fF
C33326 NAND2X1_LOC_337/B INVX1_LOC_22/A 0.07fF
C33327 INVX1_LOC_67/A INVX1_LOC_71/A 0.00fF
C33328 NOR2X1_LOC_91/A INVX1_LOC_91/A 0.17fF
C33329 NOR2X1_LOC_226/A INVX1_LOC_124/Y 0.21fF
C33330 NOR2X1_LOC_295/Y NOR2X1_LOC_607/A 0.01fF
C33331 INVX1_LOC_226/Y INPUT_3 0.09fF
C33332 NOR2X1_LOC_584/Y INVX1_LOC_38/A 0.00fF
C33333 NOR2X1_LOC_536/A NAND2X1_LOC_254/Y 0.02fF
C33334 NOR2X1_LOC_45/B NOR2X1_LOC_65/Y 0.01fF
C33335 NAND2X1_LOC_361/Y NOR2X1_LOC_350/A 0.00fF
C33336 NAND2X1_LOC_812/A NOR2X1_LOC_387/Y 0.01fF
C33337 NOR2X1_LOC_602/A NOR2X1_LOC_78/B 0.00fF
C33338 INVX1_LOC_247/Y INVX1_LOC_177/A 0.02fF
C33339 NOR2X1_LOC_162/Y INVX1_LOC_77/A 0.28fF
C33340 INVX1_LOC_95/Y INVX1_LOC_23/Y 0.19fF
C33341 INVX1_LOC_24/A INVX1_LOC_85/A 1.57fF
C33342 INVX1_LOC_269/A NOR2X1_LOC_71/Y 0.19fF
C33343 NAND2X1_LOC_338/B NAND2X1_LOC_351/A 0.05fF
C33344 INVX1_LOC_61/Y INVX1_LOC_16/A 0.08fF
C33345 INVX1_LOC_36/A NOR2X1_LOC_458/B 0.02fF
C33346 NOR2X1_LOC_533/A NAND2X1_LOC_856/A 0.02fF
C33347 NOR2X1_LOC_91/A INVX1_LOC_11/Y 0.10fF
C33348 INVX1_LOC_136/A NAND2X1_LOC_181/Y 0.03fF
C33349 NOR2X1_LOC_320/a_36_216# NOR2X1_LOC_152/Y 0.01fF
C33350 INVX1_LOC_78/A NAND2X1_LOC_453/A 0.03fF
C33351 NAND2X1_LOC_323/B NAND2X1_LOC_351/A 0.09fF
C33352 INVX1_LOC_91/A INVX1_LOC_23/A 0.25fF
C33353 NOR2X1_LOC_667/A NOR2X1_LOC_68/A 0.07fF
C33354 NOR2X1_LOC_82/A INVX1_LOC_135/A 0.18fF
C33355 NOR2X1_LOC_829/A INVX1_LOC_20/A 0.03fF
C33356 NOR2X1_LOC_65/a_36_216# INVX1_LOC_78/A 0.00fF
C33357 INVX1_LOC_248/A NOR2X1_LOC_68/A 0.07fF
C33358 INVX1_LOC_72/A INVX1_LOC_56/Y 0.02fF
C33359 D_INPUT_1 NAND2X1_LOC_642/Y 0.16fF
C33360 NOR2X1_LOC_324/B NOR2X1_LOC_383/B 0.04fF
C33361 NAND2X1_LOC_633/Y NOR2X1_LOC_438/Y 0.06fF
C33362 NAND2X1_LOC_63/Y NOR2X1_LOC_243/B 0.00fF
C33363 NOR2X1_LOC_495/Y NOR2X1_LOC_482/Y 0.02fF
C33364 INVX1_LOC_50/A NOR2X1_LOC_253/Y 0.03fF
C33365 INVX1_LOC_50/A NOR2X1_LOC_35/Y 0.00fF
C33366 NOR2X1_LOC_66/Y INVX1_LOC_19/A 0.07fF
C33367 NOR2X1_LOC_405/A NOR2X1_LOC_717/A 0.05fF
C33368 INVX1_LOC_265/A NOR2X1_LOC_309/Y 0.14fF
C33369 NAND2X1_LOC_11/Y NOR2X1_LOC_430/A 0.03fF
C33370 NAND2X1_LOC_391/Y INVX1_LOC_6/A 0.17fF
C33371 NOR2X1_LOC_298/Y NOR2X1_LOC_599/A 0.04fF
C33372 NOR2X1_LOC_273/a_36_216# INVX1_LOC_22/A 0.00fF
C33373 NOR2X1_LOC_629/B NAND2X1_LOC_562/B 0.02fF
C33374 NOR2X1_LOC_92/Y NOR2X1_LOC_368/A 0.22fF
C33375 NOR2X1_LOC_655/B NOR2X1_LOC_716/B 0.10fF
C33376 NOR2X1_LOC_334/Y INVX1_LOC_9/A 3.95fF
C33377 NOR2X1_LOC_219/Y INVX1_LOC_81/A 0.00fF
C33378 INPUT_0 NOR2X1_LOC_271/B 0.04fF
C33379 INVX1_LOC_32/A INVX1_LOC_307/A 0.07fF
C33380 NOR2X1_LOC_67/A INVX1_LOC_33/A 0.08fF
C33381 NAND2X1_LOC_860/A INVX1_LOC_20/A 0.10fF
C33382 INVX1_LOC_45/A INVX1_LOC_120/A 0.01fF
C33383 INVX1_LOC_295/A NAND2X1_LOC_36/A 0.05fF
C33384 INVX1_LOC_150/Y INVX1_LOC_131/A 0.12fF
C33385 INVX1_LOC_124/Y INPUT_1 0.30fF
C33386 INVX1_LOC_32/A NOR2X1_LOC_445/B 1.24fF
C33387 NAND2X1_LOC_254/Y INVX1_LOC_3/A 0.01fF
C33388 INVX1_LOC_167/Y INVX1_LOC_242/A 0.08fF
C33389 NOR2X1_LOC_142/Y NOR2X1_LOC_757/Y 0.10fF
C33390 INVX1_LOC_83/A NOR2X1_LOC_546/A 0.01fF
C33391 NOR2X1_LOC_605/B NOR2X1_LOC_753/Y 0.01fF
C33392 NAND2X1_LOC_361/Y NAND2X1_LOC_282/a_36_24# 0.00fF
C33393 NOR2X1_LOC_514/A NOR2X1_LOC_19/B 0.25fF
C33394 NAND2X1_LOC_81/B INVX1_LOC_29/A 2.82fF
C33395 INVX1_LOC_150/Y INPUT_0 0.07fF
C33396 NOR2X1_LOC_315/Y NAND2X1_LOC_318/a_36_24# 0.00fF
C33397 NAND2X1_LOC_181/Y NOR2X1_LOC_278/A 0.03fF
C33398 NOR2X1_LOC_316/Y INVX1_LOC_143/A 0.09fF
C33399 NOR2X1_LOC_617/Y INVX1_LOC_234/A 0.02fF
C33400 NOR2X1_LOC_82/A NOR2X1_LOC_391/B 0.19fF
C33401 INVX1_LOC_11/A INVX1_LOC_69/Y 0.07fF
C33402 INVX1_LOC_259/Y INVX1_LOC_117/A 0.03fF
C33403 INVX1_LOC_38/A NAND2X1_LOC_787/Y 0.01fF
C33404 NAND2X1_LOC_90/a_36_24# NOR2X1_LOC_271/Y 0.00fF
C33405 INVX1_LOC_159/A D_GATE_366 0.05fF
C33406 NOR2X1_LOC_249/Y NOR2X1_LOC_33/a_36_216# -0.00fF
C33407 D_INPUT_1 NOR2X1_LOC_271/Y 0.03fF
C33408 INVX1_LOC_90/A INVX1_LOC_181/Y 0.03fF
C33409 INVX1_LOC_314/Y NOR2X1_LOC_749/a_36_216# 0.01fF
C33410 NOR2X1_LOC_419/Y NOR2X1_LOC_99/B 0.23fF
C33411 INVX1_LOC_223/A NOR2X1_LOC_216/Y 0.10fF
C33412 D_INPUT_0 INVX1_LOC_49/A 2.63fF
C33413 NOR2X1_LOC_389/B INVX1_LOC_181/Y 0.02fF
C33414 NAND2X1_LOC_360/B INVX1_LOC_43/A 0.09fF
C33415 NOR2X1_LOC_769/A INVX1_LOC_75/A 0.02fF
C33416 INVX1_LOC_11/A NOR2X1_LOC_725/A 0.28fF
C33417 NOR2X1_LOC_67/A INVX1_LOC_40/A 0.07fF
C33418 INVX1_LOC_20/A NAND2X1_LOC_473/A 0.21fF
C33419 INVX1_LOC_75/A NOR2X1_LOC_554/B 0.07fF
C33420 NOR2X1_LOC_336/B NOR2X1_LOC_337/A 0.04fF
C33421 NOR2X1_LOC_284/B NOR2X1_LOC_287/A 0.00fF
C33422 INVX1_LOC_251/Y INVX1_LOC_1/Y 0.00fF
C33423 NAND2X1_LOC_82/Y INVX1_LOC_15/A 0.03fF
C33424 INVX1_LOC_161/Y NOR2X1_LOC_139/Y 0.03fF
C33425 NAND2X1_LOC_74/B INVX1_LOC_3/Y 0.01fF
C33426 INVX1_LOC_161/Y NAND2X1_LOC_655/A 0.01fF
C33427 NOR2X1_LOC_573/Y INVX1_LOC_167/Y 0.01fF
C33428 NOR2X1_LOC_68/A NAND2X1_LOC_51/B 0.05fF
C33429 INVX1_LOC_41/A NAND2X1_LOC_117/a_36_24# 0.00fF
C33430 INVX1_LOC_2/A NAND2X1_LOC_660/Y 0.12fF
C33431 NOR2X1_LOC_617/Y NOR2X1_LOC_19/B 0.51fF
C33432 INVX1_LOC_12/A INVX1_LOC_32/A 0.06fF
C33433 INVX1_LOC_162/Y NOR2X1_LOC_130/A 0.01fF
C33434 NOR2X1_LOC_561/Y NOR2X1_LOC_709/A 0.01fF
C33435 NAND2X1_LOC_537/Y INVX1_LOC_20/A 0.07fF
C33436 NAND2X1_LOC_347/B INVX1_LOC_46/A 0.02fF
C33437 D_INPUT_0 INVX1_LOC_60/A 0.02fF
C33438 INVX1_LOC_7/A NOR2X1_LOC_709/A 0.07fF
C33439 NOR2X1_LOC_773/Y INVX1_LOC_22/A 0.41fF
C33440 NOR2X1_LOC_474/A INVX1_LOC_169/A 0.01fF
C33441 INVX1_LOC_31/A INVX1_LOC_91/A 0.09fF
C33442 INVX1_LOC_58/A NOR2X1_LOC_13/a_36_216# 0.00fF
C33443 NAND2X1_LOC_538/Y INVX1_LOC_76/A 0.16fF
C33444 NOR2X1_LOC_400/B NAND2X1_LOC_659/A 0.03fF
C33445 INVX1_LOC_255/Y NAND2X1_LOC_563/A 0.10fF
C33446 NOR2X1_LOC_121/Y INPUT_1 0.01fF
C33447 NOR2X1_LOC_577/Y INVX1_LOC_140/A 0.10fF
C33448 INVX1_LOC_29/A INVX1_LOC_4/Y 0.18fF
C33449 NOR2X1_LOC_598/B NOR2X1_LOC_156/Y 0.03fF
C33450 NOR2X1_LOC_100/A INVX1_LOC_135/A 0.01fF
C33451 INVX1_LOC_75/A NOR2X1_LOC_152/Y 0.13fF
C33452 INVX1_LOC_2/A D_INPUT_0 0.15fF
C33453 NAND2X1_LOC_563/Y INVX1_LOC_90/A 0.04fF
C33454 INVX1_LOC_300/A NAND2X1_LOC_863/B 0.03fF
C33455 NOR2X1_LOC_510/Y INVX1_LOC_118/Y 0.07fF
C33456 NAND2X1_LOC_273/a_36_24# INVX1_LOC_23/A 0.01fF
C33457 INVX1_LOC_75/A INVX1_LOC_113/Y 0.05fF
C33458 NOR2X1_LOC_647/a_36_216# INVX1_LOC_59/Y 0.00fF
C33459 INVX1_LOC_104/A INVX1_LOC_196/Y 0.12fF
C33460 NAND2X1_LOC_364/a_36_24# INVX1_LOC_143/A 0.00fF
C33461 NOR2X1_LOC_179/Y INVX1_LOC_23/A 0.18fF
C33462 NOR2X1_LOC_226/A D_INPUT_0 0.07fF
C33463 NAND2X1_LOC_99/A NAND2X1_LOC_772/a_36_24# 0.00fF
C33464 INVX1_LOC_5/A NOR2X1_LOC_88/A 0.01fF
C33465 INVX1_LOC_305/A NOR2X1_LOC_78/A 0.07fF
C33466 NOR2X1_LOC_100/A NOR2X1_LOC_560/A 0.03fF
C33467 INVX1_LOC_12/A NAND2X1_LOC_175/Y 0.10fF
C33468 NOR2X1_LOC_503/Y NAND2X1_LOC_453/A 0.07fF
C33469 INVX1_LOC_203/A INVX1_LOC_23/A 0.05fF
C33470 INVX1_LOC_41/Y NOR2X1_LOC_528/Y 0.03fF
C33471 NOR2X1_LOC_454/Y NAND2X1_LOC_637/Y 0.09fF
C33472 GATE_662 NAND2X1_LOC_663/a_36_24# 0.02fF
C33473 NOR2X1_LOC_569/Y NOR2X1_LOC_549/a_36_216# 0.00fF
C33474 NOR2X1_LOC_82/A NOR2X1_LOC_813/Y 0.15fF
C33475 INVX1_LOC_21/A NAND2X1_LOC_430/a_36_24# 0.00fF
C33476 NOR2X1_LOC_279/a_36_216# NAND2X1_LOC_807/Y 0.00fF
C33477 NAND2X1_LOC_861/Y INVX1_LOC_25/Y 0.07fF
C33478 INVX1_LOC_197/Y NAND2X1_LOC_624/A 0.06fF
C33479 NOR2X1_LOC_307/A INVX1_LOC_117/A 0.00fF
C33480 NOR2X1_LOC_376/a_36_216# INVX1_LOC_91/A 0.00fF
C33481 INVX1_LOC_103/A NOR2X1_LOC_331/B 0.10fF
C33482 INVX1_LOC_245/A INVX1_LOC_89/A 0.01fF
C33483 NOR2X1_LOC_391/A NAND2X1_LOC_384/a_36_24# 0.00fF
C33484 NOR2X1_LOC_720/B NOR2X1_LOC_188/A 0.01fF
C33485 NOR2X1_LOC_1/a_36_216# D_INPUT_4 0.00fF
C33486 NOR2X1_LOC_82/A INVX1_LOC_280/A 0.14fF
C33487 INVX1_LOC_58/A NAND2X1_LOC_74/B 0.06fF
C33488 NOR2X1_LOC_828/Y NOR2X1_LOC_777/B 0.07fF
C33489 NOR2X1_LOC_471/Y NOR2X1_LOC_684/Y -0.00fF
C33490 INVX1_LOC_228/A INVX1_LOC_316/A 0.18fF
C33491 INVX1_LOC_90/A INVX1_LOC_32/Y 0.01fF
C33492 NOR2X1_LOC_526/Y NAND2X1_LOC_560/A 0.01fF
C33493 NOR2X1_LOC_250/Y INVX1_LOC_118/A 0.25fF
C33494 INVX1_LOC_299/A NOR2X1_LOC_809/B 0.00fF
C33495 NOR2X1_LOC_437/Y NAND2X1_LOC_468/B 0.02fF
C33496 NOR2X1_LOC_520/B NAND2X1_LOC_490/a_36_24# 0.00fF
C33497 INVX1_LOC_63/Y NOR2X1_LOC_43/a_36_216# 0.00fF
C33498 INVX1_LOC_5/A INVX1_LOC_186/Y 0.24fF
C33499 NOR2X1_LOC_92/Y INVX1_LOC_260/Y 0.08fF
C33500 NOR2X1_LOC_246/A NAND2X1_LOC_808/A 0.43fF
C33501 INVX1_LOC_290/A NAND2X1_LOC_654/B 0.05fF
C33502 INVX1_LOC_140/A INVX1_LOC_22/A 0.04fF
C33503 INVX1_LOC_227/A NOR2X1_LOC_473/B 0.02fF
C33504 NOR2X1_LOC_488/Y NOR2X1_LOC_322/Y 0.02fF
C33505 INVX1_LOC_298/Y INVX1_LOC_4/Y 0.03fF
C33506 NAND2X1_LOC_549/Y NOR2X1_LOC_671/Y 0.01fF
C33507 D_INPUT_1 NAND2X1_LOC_792/B 0.23fF
C33508 INVX1_LOC_136/A INVX1_LOC_117/A 0.10fF
C33509 NAND2X1_LOC_79/Y VDD 0.02fF
C33510 INVX1_LOC_103/A NOR2X1_LOC_592/B 0.03fF
C33511 INVX1_LOC_13/Y INVX1_LOC_19/A 0.10fF
C33512 INVX1_LOC_71/A NOR2X1_LOC_137/Y 0.03fF
C33513 NOR2X1_LOC_773/Y INVX1_LOC_100/A 0.02fF
C33514 D_INPUT_0 INPUT_1 1.18fF
C33515 NAND2X1_LOC_463/B INVX1_LOC_22/A 0.00fF
C33516 NAND2X1_LOC_854/B NAND2X1_LOC_740/B 0.04fF
C33517 INVX1_LOC_217/A NOR2X1_LOC_692/Y 0.03fF
C33518 NOR2X1_LOC_120/a_36_216# NOR2X1_LOC_99/B 0.01fF
C33519 NOR2X1_LOC_152/Y NOR2X1_LOC_65/a_36_216# 0.00fF
C33520 INVX1_LOC_191/Y INVX1_LOC_91/A 0.02fF
C33521 NOR2X1_LOC_598/B D_INPUT_5 0.07fF
C33522 NOR2X1_LOC_717/B INVX1_LOC_182/A 0.00fF
C33523 NOR2X1_LOC_599/Y NAND2X1_LOC_802/Y 0.18fF
C33524 INVX1_LOC_181/Y NOR2X1_LOC_561/A 0.01fF
C33525 NOR2X1_LOC_595/Y NAND2X1_LOC_660/A 0.10fF
C33526 INVX1_LOC_175/A NAND2X1_LOC_416/a_36_24# 0.02fF
C33527 NOR2X1_LOC_191/A INVX1_LOC_98/A 0.01fF
C33528 INVX1_LOC_33/A NOR2X1_LOC_558/A 0.06fF
C33529 NAND2X1_LOC_860/A INVX1_LOC_4/A 0.08fF
C33530 INVX1_LOC_77/A NAND2X1_LOC_472/Y 0.07fF
C33531 INVX1_LOC_14/A NOR2X1_LOC_662/A 0.02fF
C33532 NOR2X1_LOC_336/B NOR2X1_LOC_640/Y 0.02fF
C33533 INVX1_LOC_251/Y INVX1_LOC_93/Y 0.01fF
C33534 NOR2X1_LOC_64/a_36_216# INVX1_LOC_20/A 0.00fF
C33535 INVX1_LOC_292/Y NOR2X1_LOC_801/B 0.01fF
C33536 INVX1_LOC_162/A NAND2X1_LOC_287/B 0.36fF
C33537 INVX1_LOC_314/Y NOR2X1_LOC_536/A 0.09fF
C33538 NOR2X1_LOC_688/Y NOR2X1_LOC_862/B 0.13fF
C33539 INVX1_LOC_6/A INVX1_LOC_137/Y 0.02fF
C33540 NOR2X1_LOC_716/B NOR2X1_LOC_176/Y 0.01fF
C33541 NAND2X1_LOC_656/Y NOR2X1_LOC_335/B 0.07fF
C33542 INVX1_LOC_141/Y NOR2X1_LOC_88/Y 0.03fF
C33543 INVX1_LOC_88/A INVX1_LOC_19/A 0.05fF
C33544 INVX1_LOC_143/A INVX1_LOC_314/A 0.04fF
C33545 NOR2X1_LOC_52/Y NOR2X1_LOC_435/A 0.01fF
C33546 INVX1_LOC_53/A NOR2X1_LOC_158/Y 0.07fF
C33547 NOR2X1_LOC_709/A INVX1_LOC_76/A 0.01fF
C33548 INVX1_LOC_223/A NOR2X1_LOC_197/B 0.03fF
C33549 INVX1_LOC_72/Y NOR2X1_LOC_99/Y 0.08fF
C33550 INVX1_LOC_28/A NAND2X1_LOC_652/Y 0.01fF
C33551 NAND2X1_LOC_787/B NOR2X1_LOC_692/Y 0.11fF
C33552 INVX1_LOC_72/A NOR2X1_LOC_831/B 0.03fF
C33553 NAND2X1_LOC_51/B NOR2X1_LOC_163/A 0.00fF
C33554 NOR2X1_LOC_733/a_36_216# INVX1_LOC_179/A 0.00fF
C33555 NOR2X1_LOC_848/Y NOR2X1_LOC_340/A 0.19fF
C33556 INVX1_LOC_227/A NOR2X1_LOC_355/B 0.01fF
C33557 INVX1_LOC_141/Y INVX1_LOC_84/A 0.03fF
C33558 NOR2X1_LOC_596/A NOR2X1_LOC_433/Y 0.01fF
C33559 INVX1_LOC_31/A INVX1_LOC_203/A 0.10fF
C33560 NOR2X1_LOC_635/B NOR2X1_LOC_452/A 0.02fF
C33561 INVX1_LOC_95/Y INVX1_LOC_232/A 0.10fF
C33562 INVX1_LOC_224/A NOR2X1_LOC_89/A 0.03fF
C33563 INVX1_LOC_89/A NOR2X1_LOC_147/A 0.01fF
C33564 NOR2X1_LOC_226/A NOR2X1_LOC_266/B 0.13fF
C33565 INVX1_LOC_314/Y NAND2X1_LOC_93/B 0.10fF
C33566 INVX1_LOC_33/A NOR2X1_LOC_729/A 0.13fF
C33567 INVX1_LOC_11/A NOR2X1_LOC_89/A 0.63fF
C33568 NOR2X1_LOC_226/A NOR2X1_LOC_682/Y 0.01fF
C33569 INVX1_LOC_33/A NAND2X1_LOC_268/a_36_24# 0.01fF
C33570 NAND2X1_LOC_35/Y INVX1_LOC_26/A 0.02fF
C33571 NOR2X1_LOC_383/Y INVX1_LOC_95/Y 0.65fF
C33572 INVX1_LOC_276/A NOR2X1_LOC_816/Y 0.01fF
C33573 NOR2X1_LOC_718/B INVX1_LOC_9/A 0.07fF
C33574 INPUT_3 INVX1_LOC_12/A 0.03fF
C33575 NOR2X1_LOC_468/Y INVX1_LOC_47/Y 0.02fF
C33576 INVX1_LOC_313/A INVX1_LOC_91/A 0.09fF
C33577 INVX1_LOC_2/A NAND2X1_LOC_848/A 0.10fF
C33578 INVX1_LOC_217/A NAND2X1_LOC_489/Y 0.03fF
C33579 NOR2X1_LOC_100/A INVX1_LOC_280/A -0.01fF
C33580 NOR2X1_LOC_500/B INVX1_LOC_19/A 0.17fF
C33581 NAND2X1_LOC_866/B INVX1_LOC_91/A 0.08fF
C33582 INVX1_LOC_5/A NOR2X1_LOC_843/B 0.04fF
C33583 NOR2X1_LOC_489/B INVX1_LOC_57/A 0.06fF
C33584 NOR2X1_LOC_717/a_36_216# NOR2X1_LOC_155/A 0.00fF
C33585 NOR2X1_LOC_748/Y VDD 0.28fF
C33586 NOR2X1_LOC_186/Y NOR2X1_LOC_318/A 0.07fF
C33587 INVX1_LOC_228/Y INVX1_LOC_32/A 0.03fF
C33588 NOR2X1_LOC_226/A NAND2X1_LOC_848/A 0.10fF
C33589 INVX1_LOC_11/A NOR2X1_LOC_170/A 0.00fF
C33590 NOR2X1_LOC_92/Y NAND2X1_LOC_471/Y 0.02fF
C33591 INVX1_LOC_135/A NOR2X1_LOC_124/a_36_216# 0.00fF
C33592 NOR2X1_LOC_714/Y NOR2X1_LOC_729/A 0.05fF
C33593 INVX1_LOC_135/A INVX1_LOC_59/Y 0.27fF
C33594 NOR2X1_LOC_382/Y NOR2X1_LOC_671/a_36_216# 0.00fF
C33595 INVX1_LOC_135/A INVX1_LOC_112/A 0.03fF
C33596 INVX1_LOC_79/A INVX1_LOC_6/A 0.00fF
C33597 NAND2X1_LOC_807/Y INVX1_LOC_91/A 0.08fF
C33598 INVX1_LOC_202/A NAND2X1_LOC_475/Y 0.66fF
C33599 NAND2X1_LOC_562/B NOR2X1_LOC_88/A 0.02fF
C33600 INVX1_LOC_286/Y INVX1_LOC_102/A 0.25fF
C33601 INVX1_LOC_90/A NOR2X1_LOC_675/A 0.01fF
C33602 NAND2X1_LOC_866/B INVX1_LOC_11/Y 0.07fF
C33603 NAND2X1_LOC_35/Y NOR2X1_LOC_255/Y 0.12fF
C33604 NOR2X1_LOC_658/Y INVX1_LOC_109/Y 0.10fF
C33605 INVX1_LOC_135/A INVX1_LOC_176/A 0.04fF
C33606 NOR2X1_LOC_389/B NOR2X1_LOC_675/A -0.01fF
C33607 NAND2X1_LOC_114/B INVX1_LOC_15/A 0.07fF
C33608 NAND2X1_LOC_573/Y NOR2X1_LOC_318/A 0.07fF
C33609 INVX1_LOC_50/A NAND2X1_LOC_794/B 0.04fF
C33610 NAND2X1_LOC_833/Y INVX1_LOC_285/A 0.02fF
C33611 NOR2X1_LOC_742/A NOR2X1_LOC_555/a_36_216# 0.01fF
C33612 NOR2X1_LOC_106/A INVX1_LOC_76/A 0.06fF
C33613 NOR2X1_LOC_363/Y NOR2X1_LOC_665/A 0.14fF
C33614 NOR2X1_LOC_15/Y NOR2X1_LOC_301/A 0.03fF
C33615 NOR2X1_LOC_454/Y NOR2X1_LOC_639/Y 0.05fF
C33616 NAND2X1_LOC_833/Y INVX1_LOC_265/Y 0.43fF
C33617 NOR2X1_LOC_71/Y NAND2X1_LOC_457/a_36_24# 0.01fF
C33618 NAND2X1_LOC_773/Y INVX1_LOC_23/Y 0.02fF
C33619 NOR2X1_LOC_156/B NOR2X1_LOC_156/Y 0.08fF
C33620 INVX1_LOC_27/A INVX1_LOC_270/Y 0.07fF
C33621 INVX1_LOC_32/Y INVX1_LOC_38/A 0.02fF
C33622 NAND2X1_LOC_319/a_36_24# INVX1_LOC_118/A 0.00fF
C33623 NAND2X1_LOC_470/a_36_24# NOR2X1_LOC_435/A 0.00fF
C33624 INVX1_LOC_298/Y NOR2X1_LOC_205/Y 0.03fF
C33625 INVX1_LOC_34/A NOR2X1_LOC_673/A 0.03fF
C33626 INVX1_LOC_2/A INVX1_LOC_46/Y 0.10fF
C33627 INVX1_LOC_269/A INVX1_LOC_16/Y 0.20fF
C33628 INVX1_LOC_303/A INVX1_LOC_19/A 0.07fF
C33629 INVX1_LOC_103/A NOR2X1_LOC_449/A 0.19fF
C33630 NOR2X1_LOC_792/a_36_216# INVX1_LOC_57/A 0.00fF
C33631 INVX1_LOC_176/A NOR2X1_LOC_560/A 0.03fF
C33632 INVX1_LOC_266/Y INVX1_LOC_107/Y 0.10fF
C33633 INVX1_LOC_65/Y VDD 0.36fF
C33634 NOR2X1_LOC_213/a_36_216# INVX1_LOC_179/A 0.00fF
C33635 INPUT_1 NOR2X1_LOC_266/B 1.04fF
C33636 NOR2X1_LOC_71/Y INVX1_LOC_12/Y 0.10fF
C33637 NOR2X1_LOC_226/A INVX1_LOC_46/Y -0.01fF
C33638 INVX1_LOC_312/Y INVX1_LOC_15/A 0.07fF
C33639 NOR2X1_LOC_569/Y INVX1_LOC_9/A 0.08fF
C33640 NAND2X1_LOC_357/B INVX1_LOC_119/Y 0.02fF
C33641 NOR2X1_LOC_596/Y INVX1_LOC_271/Y 0.05fF
C33642 D_GATE_366 VDD 0.18fF
C33643 NAND2X1_LOC_579/A NOR2X1_LOC_654/A 0.03fF
C33644 NOR2X1_LOC_523/B NOR2X1_LOC_861/Y 0.06fF
C33645 INVX1_LOC_136/A INVX1_LOC_3/Y 0.20fF
C33646 INVX1_LOC_35/A NOR2X1_LOC_460/Y 0.02fF
C33647 INVX1_LOC_6/A INVX1_LOC_91/A 0.15fF
C33648 NOR2X1_LOC_356/A INVX1_LOC_14/Y 0.03fF
C33649 NAND2X1_LOC_59/B INVX1_LOC_19/A 0.02fF
C33650 NOR2X1_LOC_813/Y NOR2X1_LOC_132/a_36_216# 0.01fF
C33651 INVX1_LOC_14/A INVX1_LOC_57/A 0.09fF
C33652 NOR2X1_LOC_180/Y INVX1_LOC_63/A 0.03fF
C33653 NOR2X1_LOC_433/A NOR2X1_LOC_89/A 0.14fF
C33654 NAND2X1_LOC_550/A NOR2X1_LOC_693/Y 0.01fF
C33655 NAND2X1_LOC_863/A INVX1_LOC_76/A 0.10fF
C33656 NAND2X1_LOC_733/Y NAND2X1_LOC_175/Y 0.10fF
C33657 NAND2X1_LOC_807/Y NOR2X1_LOC_653/a_36_216# 0.00fF
C33658 NAND2X1_LOC_733/Y NOR2X1_LOC_821/a_36_216# 0.00fF
C33659 INVX1_LOC_8/A NAND2X1_LOC_81/B 0.03fF
C33660 NOR2X1_LOC_289/Y VDD 0.13fF
C33661 NOR2X1_LOC_593/Y NOR2X1_LOC_89/A 0.02fF
C33662 NOR2X1_LOC_843/A INVX1_LOC_29/A 0.05fF
C33663 NAND2X1_LOC_848/A INPUT_1 0.03fF
C33664 NOR2X1_LOC_577/Y INVX1_LOC_42/A 0.15fF
C33665 NOR2X1_LOC_391/B INVX1_LOC_59/Y 0.07fF
C33666 NAND2X1_LOC_355/Y NOR2X1_LOC_329/Y 0.03fF
C33667 D_INPUT_0 INVX1_LOC_118/A 0.16fF
C33668 NOR2X1_LOC_274/B INVX1_LOC_78/A 0.07fF
C33669 INVX1_LOC_82/A INVX1_LOC_29/A 0.02fF
C33670 INVX1_LOC_113/Y INVX1_LOC_283/A 0.00fF
C33671 NOR2X1_LOC_348/B INVX1_LOC_263/Y 0.01fF
C33672 NOR2X1_LOC_86/a_36_216# INVX1_LOC_20/A 0.00fF
C33673 NOR2X1_LOC_456/Y NOR2X1_LOC_457/A 0.41fF
C33674 INVX1_LOC_298/Y NOR2X1_LOC_723/Y 0.01fF
C33675 NOR2X1_LOC_74/A INVX1_LOC_14/Y 0.01fF
C33676 INVX1_LOC_64/A NAND2X1_LOC_537/Y 0.07fF
C33677 NOR2X1_LOC_500/B INVX1_LOC_26/Y 0.06fF
C33678 INVX1_LOC_21/A NAND2X1_LOC_474/Y 0.07fF
C33679 NOR2X1_LOC_742/A INVX1_LOC_281/A 0.01fF
C33680 INVX1_LOC_58/A NOR2X1_LOC_276/Y 0.01fF
C33681 NOR2X1_LOC_52/B NOR2X1_LOC_89/A 0.16fF
C33682 INVX1_LOC_292/A NOR2X1_LOC_493/A 0.14fF
C33683 INVX1_LOC_185/Y INVX1_LOC_102/A 0.01fF
C33684 NAND2X1_LOC_361/a_36_24# INVX1_LOC_42/A 0.01fF
C33685 NAND2X1_LOC_124/a_36_24# NOR2X1_LOC_363/Y 0.00fF
C33686 NOR2X1_LOC_803/A NOR2X1_LOC_209/B 0.00fF
C33687 NOR2X1_LOC_348/B INVX1_LOC_42/A 0.03fF
C33688 NOR2X1_LOC_97/A NAND2X1_LOC_96/A 0.05fF
C33689 INVX1_LOC_299/A INVX1_LOC_50/Y 0.10fF
C33690 NAND2X1_LOC_858/B INVX1_LOC_33/Y 0.02fF
C33691 NOR2X1_LOC_668/a_36_216# INVX1_LOC_31/A 0.01fF
C33692 INPUT_1 INVX1_LOC_46/Y 0.07fF
C33693 INVX1_LOC_88/Y INVX1_LOC_15/A 0.03fF
C33694 NOR2X1_LOC_295/Y INVX1_LOC_47/Y 0.01fF
C33695 INVX1_LOC_55/Y INVX1_LOC_92/A 0.03fF
C33696 INVX1_LOC_35/A INVX1_LOC_110/Y 0.07fF
C33697 INVX1_LOC_95/Y NAND2X1_LOC_447/Y 0.19fF
C33698 INVX1_LOC_14/A INVX1_LOC_252/A 0.04fF
C33699 NOR2X1_LOC_577/Y INVX1_LOC_78/A 1.72fF
C33700 INVX1_LOC_238/A INVX1_LOC_233/Y 0.00fF
C33701 NAND2X1_LOC_656/Y INVX1_LOC_84/A 0.22fF
C33702 INVX1_LOC_58/A INVX1_LOC_136/A 0.43fF
C33703 NOR2X1_LOC_746/Y VDD 0.13fF
C33704 INVX1_LOC_8/A INVX1_LOC_4/Y 0.17fF
C33705 INVX1_LOC_206/Y INVX1_LOC_44/A 0.07fF
C33706 NOR2X1_LOC_45/B NAND2X1_LOC_721/A 0.03fF
C33707 NOR2X1_LOC_294/Y INVX1_LOC_108/Y 0.04fF
C33708 INVX1_LOC_21/A NAND2X1_LOC_53/Y 0.14fF
C33709 INVX1_LOC_22/A INVX1_LOC_263/Y 0.01fF
C33710 NOR2X1_LOC_265/a_36_216# INVX1_LOC_102/A 0.01fF
C33711 NAND2X1_LOC_571/B NOR2X1_LOC_384/Y 0.01fF
C33712 INVX1_LOC_34/A NOR2X1_LOC_409/B 0.03fF
C33713 INVX1_LOC_266/A INVX1_LOC_299/A 0.00fF
C33714 NAND2X1_LOC_786/a_36_24# INVX1_LOC_26/A 0.00fF
C33715 INVX1_LOC_303/A INVX1_LOC_26/Y 0.14fF
C33716 NOR2X1_LOC_168/B INVX1_LOC_15/A 0.02fF
C33717 INVX1_LOC_88/A NOR2X1_LOC_122/A 0.03fF
C33718 NAND2X1_LOC_84/Y INVX1_LOC_57/A 0.03fF
C33719 D_INPUT_1 NOR2X1_LOC_359/Y 0.01fF
C33720 NOR2X1_LOC_65/B NOR2X1_LOC_577/Y 0.00fF
C33721 NAND2X1_LOC_477/A NAND2X1_LOC_471/Y 0.02fF
C33722 INVX1_LOC_17/A NOR2X1_LOC_15/Y 0.06fF
C33723 INVX1_LOC_22/A INVX1_LOC_42/A 0.22fF
C33724 NOR2X1_LOC_348/B INVX1_LOC_78/A 0.07fF
C33725 NOR2X1_LOC_189/A INVX1_LOC_50/A 0.04fF
C33726 D_INPUT_0 NAND2X1_LOC_63/Y 0.06fF
C33727 NOR2X1_LOC_817/Y INVX1_LOC_269/A 0.02fF
C33728 NOR2X1_LOC_658/a_36_216# INVX1_LOC_63/Y 0.01fF
C33729 NAND2X1_LOC_465/Y INVX1_LOC_26/A 0.07fF
C33730 INVX1_LOC_36/Y VDD 0.50fF
C33731 INVX1_LOC_225/A NOR2X1_LOC_318/A 0.01fF
C33732 NAND2X1_LOC_552/A INVX1_LOC_18/A 0.03fF
C33733 INVX1_LOC_224/A INVX1_LOC_11/A 0.03fF
C33734 NOR2X1_LOC_471/Y NOR2X1_LOC_15/Y 0.03fF
C33735 INVX1_LOC_230/Y NOR2X1_LOC_92/Y 0.04fF
C33736 INVX1_LOC_135/A NOR2X1_LOC_340/A 0.03fF
C33737 INVX1_LOC_255/Y NOR2X1_LOC_554/A 0.00fF
C33738 INVX1_LOC_251/Y INVX1_LOC_87/A 0.05fF
C33739 INVX1_LOC_88/A INVX1_LOC_161/Y 0.11fF
C33740 INVX1_LOC_73/A INVX1_LOC_285/A 0.07fF
C33741 INVX1_LOC_5/A INVX1_LOC_18/A 4.56fF
C33742 NOR2X1_LOC_813/Y INVX1_LOC_59/Y 0.11fF
C33743 INVX1_LOC_179/Y NOR2X1_LOC_334/Y 0.01fF
C33744 INVX1_LOC_48/Y INVX1_LOC_61/Y 0.55fF
C33745 NOR2X1_LOC_528/Y INVX1_LOC_185/A 0.01fF
C33746 INVX1_LOC_37/Y NAND2X1_LOC_242/a_36_24# 0.00fF
C33747 INVX1_LOC_73/A NOR2X1_LOC_814/A 0.03fF
C33748 INVX1_LOC_11/A NAND2X1_LOC_381/Y 0.24fF
C33749 NOR2X1_LOC_643/A INPUT_3 0.02fF
C33750 NOR2X1_LOC_124/a_36_216# INVX1_LOC_280/A 0.00fF
C33751 NOR2X1_LOC_738/Y NOR2X1_LOC_307/A 0.01fF
C33752 NOR2X1_LOC_111/A INVX1_LOC_37/A 0.07fF
C33753 INVX1_LOC_301/Y INVX1_LOC_213/A 0.02fF
C33754 NAND2X1_LOC_633/Y NOR2X1_LOC_176/Y 0.01fF
C33755 INVX1_LOC_25/Y NOR2X1_LOC_89/a_36_216# 0.01fF
C33756 NOR2X1_LOC_315/Y NOR2X1_LOC_72/Y 0.00fF
C33757 INVX1_LOC_59/Y INVX1_LOC_280/A 0.20fF
C33758 INVX1_LOC_112/A INVX1_LOC_280/A 0.05fF
C33759 NAND2X1_LOC_799/A NOR2X1_LOC_816/A 0.44fF
C33760 NOR2X1_LOC_211/Y NOR2X1_LOC_303/Y 0.04fF
C33761 INVX1_LOC_228/Y INPUT_3 0.01fF
C33762 INVX1_LOC_178/A INVX1_LOC_18/A 0.10fF
C33763 NOR2X1_LOC_131/Y NAND2X1_LOC_454/Y 0.03fF
C33764 INVX1_LOC_139/A INVX1_LOC_281/A 0.35fF
C33765 NAND2X1_LOC_513/B INVX1_LOC_142/A 0.21fF
C33766 NOR2X1_LOC_710/B NOR2X1_LOC_710/A 0.02fF
C33767 NAND2X1_LOC_720/a_36_24# NAND2X1_LOC_703/Y -0.02fF
C33768 INVX1_LOC_38/A INVX1_LOC_115/A 0.00fF
C33769 NOR2X1_LOC_843/A NOR2X1_LOC_843/a_36_216# 0.02fF
C33770 NOR2X1_LOC_45/B INVX1_LOC_117/Y 0.03fF
C33771 NAND2X1_LOC_440/a_36_24# NOR2X1_LOC_331/B 0.00fF
C33772 INVX1_LOC_176/A INVX1_LOC_280/A 0.04fF
C33773 NOR2X1_LOC_666/Y NOR2X1_LOC_717/Y 0.21fF
C33774 INVX1_LOC_93/A INVX1_LOC_41/Y 0.02fF
C33775 NOR2X1_LOC_91/A NAND2X1_LOC_374/Y 0.07fF
C33776 NAND2X1_LOC_561/B INVX1_LOC_30/A 0.09fF
C33777 NOR2X1_LOC_269/Y NOR2X1_LOC_155/A 0.07fF
C33778 INVX1_LOC_22/A INVX1_LOC_78/A 0.36fF
C33779 NOR2X1_LOC_612/B INVX1_LOC_57/A 0.00fF
C33780 INVX1_LOC_172/A INVX1_LOC_5/A 0.00fF
C33781 INVX1_LOC_50/A NOR2X1_LOC_482/Y 0.13fF
C33782 NAND2X1_LOC_725/A INVX1_LOC_207/A 0.22fF
C33783 NOR2X1_LOC_644/A NOR2X1_LOC_842/a_36_216# 0.00fF
C33784 INVX1_LOC_58/A NAND2X1_LOC_859/a_36_24# 0.00fF
C33785 NOR2X1_LOC_589/A NAND2X1_LOC_454/Y 0.05fF
C33786 INVX1_LOC_13/Y NAND2X1_LOC_119/a_36_24# 0.01fF
C33787 NOR2X1_LOC_561/Y NOR2X1_LOC_334/Y 0.10fF
C33788 NOR2X1_LOC_78/B NOR2X1_LOC_646/B 0.01fF
C33789 NOR2X1_LOC_420/a_36_216# NOR2X1_LOC_716/B 0.00fF
C33790 INVX1_LOC_6/A INVX1_LOC_203/A 0.00fF
C33791 NOR2X1_LOC_454/Y INVX1_LOC_24/A 0.07fF
C33792 INVX1_LOC_91/A NOR2X1_LOC_117/Y 0.04fF
C33793 NOR2X1_LOC_533/Y NAND2X1_LOC_856/A 0.03fF
C33794 INVX1_LOC_64/A NOR2X1_LOC_143/a_36_216# 0.00fF
C33795 NOR2X1_LOC_769/B NAND2X1_LOC_451/Y 0.04fF
C33796 INVX1_LOC_272/Y NAND2X1_LOC_354/Y 0.04fF
C33797 NOR2X1_LOC_68/A NOR2X1_LOC_523/A 0.07fF
C33798 INVX1_LOC_172/A INVX1_LOC_178/A 0.14fF
C33799 INVX1_LOC_288/A INVX1_LOC_22/A 0.01fF
C33800 NOR2X1_LOC_641/B NOR2X1_LOC_160/B 0.08fF
C33801 NOR2X1_LOC_130/a_36_216# NOR2X1_LOC_38/B 0.00fF
C33802 NOR2X1_LOC_65/B INVX1_LOC_22/A 1.01fF
C33803 NOR2X1_LOC_216/Y INVX1_LOC_290/Y 0.03fF
C33804 INVX1_LOC_116/A INVX1_LOC_1/A 0.01fF
C33805 NAND2X1_LOC_472/Y INVX1_LOC_9/A 0.07fF
C33806 NOR2X1_LOC_598/B NAND2X1_LOC_451/Y 0.63fF
C33807 INVX1_LOC_224/Y NOR2X1_LOC_121/a_36_216# 0.00fF
C33808 INVX1_LOC_83/A NOR2X1_LOC_158/Y 0.10fF
C33809 NOR2X1_LOC_357/Y INVX1_LOC_92/A 0.07fF
C33810 NAND2X1_LOC_468/B NOR2X1_LOC_841/A 0.03fF
C33811 INVX1_LOC_224/Y INVX1_LOC_56/Y 0.00fF
C33812 INVX1_LOC_136/A INVX1_LOC_215/Y 0.03fF
C33813 NOR2X1_LOC_678/a_36_216# NOR2X1_LOC_433/A 0.01fF
C33814 NAND2X1_LOC_654/B NOR2X1_LOC_467/A 0.02fF
C33815 NAND2X1_LOC_808/A NAND2X1_LOC_175/Y 0.03fF
C33816 VDD INVX1_LOC_70/A 0.34fF
C33817 NOR2X1_LOC_448/Y INVX1_LOC_49/A 0.01fF
C33818 NOR2X1_LOC_751/Y NOR2X1_LOC_160/B 0.11fF
C33819 INVX1_LOC_39/A NOR2X1_LOC_121/Y 0.01fF
C33820 NOR2X1_LOC_816/A INVX1_LOC_18/A 5.17fF
C33821 NOR2X1_LOC_437/Y INVX1_LOC_88/A 0.02fF
C33822 NOR2X1_LOC_211/Y INVX1_LOC_54/Y 0.01fF
C33823 INVX1_LOC_53/Y INVX1_LOC_29/Y 0.03fF
C33824 D_GATE_741 INVX1_LOC_198/Y 0.04fF
C33825 NOR2X1_LOC_111/A NOR2X1_LOC_743/Y 0.04fF
C33826 NOR2X1_LOC_71/Y NOR2X1_LOC_89/Y -0.00fF
C33827 NAND2X1_LOC_848/A INVX1_LOC_118/A 0.17fF
C33828 NOR2X1_LOC_447/B NAND2X1_LOC_798/B 0.01fF
C33829 NAND2X1_LOC_579/A NOR2X1_LOC_716/B 0.10fF
C33830 INVX1_LOC_17/A NOR2X1_LOC_860/B 0.16fF
C33831 INVX1_LOC_37/A NOR2X1_LOC_600/a_36_216# 0.00fF
C33832 INVX1_LOC_100/A INVX1_LOC_42/A -0.04fF
C33833 NAND2X1_LOC_361/Y INVX1_LOC_1/A 0.08fF
C33834 INVX1_LOC_81/Y INVX1_LOC_72/A 0.03fF
C33835 NOR2X1_LOC_332/A NOR2X1_LOC_843/B 0.08fF
C33836 NAND2X1_LOC_36/A NAND2X1_LOC_387/B 0.17fF
C33837 NOR2X1_LOC_669/Y NAND2X1_LOC_325/Y 0.01fF
C33838 VDD INVX1_LOC_123/Y 0.23fF
C33839 NOR2X1_LOC_391/A NAND2X1_LOC_215/A 0.12fF
C33840 INVX1_LOC_45/Y NOR2X1_LOC_160/B 0.12fF
C33841 INVX1_LOC_256/A INVX1_LOC_314/Y 0.16fF
C33842 NAND2X1_LOC_711/B NOR2X1_LOC_816/A 0.00fF
C33843 INVX1_LOC_11/A NOR2X1_LOC_433/A 0.14fF
C33844 INVX1_LOC_64/A INVX1_LOC_172/Y 0.88fF
C33845 INVX1_LOC_25/A NOR2X1_LOC_789/a_36_216# 0.00fF
C33846 INVX1_LOC_45/A NAND2X1_LOC_351/A 0.08fF
C33847 NAND2X1_LOC_30/Y INVX1_LOC_49/A -0.02fF
C33848 INVX1_LOC_230/Y NAND2X1_LOC_837/Y 0.00fF
C33849 INVX1_LOC_11/A NOR2X1_LOC_593/Y 0.47fF
C33850 NAND2X1_LOC_677/a_36_24# NOR2X1_LOC_833/B 0.00fF
C33851 NOR2X1_LOC_137/A INVX1_LOC_57/A 0.00fF
C33852 INVX1_LOC_299/A NOR2X1_LOC_6/B -0.04fF
C33853 NOR2X1_LOC_273/Y INVX1_LOC_30/A 0.03fF
C33854 INVX1_LOC_30/A NOR2X1_LOC_759/Y 0.03fF
C33855 INVX1_LOC_78/Y INVX1_LOC_15/A 0.05fF
C33856 INPUT_0 NOR2X1_LOC_409/B 0.05fF
C33857 INVX1_LOC_311/Y NOR2X1_LOC_727/B 0.02fF
C33858 INVX1_LOC_202/A INVX1_LOC_30/A 0.18fF
C33859 INVX1_LOC_21/A NOR2X1_LOC_500/Y 0.07fF
C33860 NOR2X1_LOC_167/Y NAND2X1_LOC_444/B 0.01fF
C33861 INVX1_LOC_21/A INVX1_LOC_226/Y 0.98fF
C33862 NOR2X1_LOC_246/A INVX1_LOC_53/A 0.44fF
C33863 INVX1_LOC_11/A NOR2X1_LOC_52/B 0.06fF
C33864 INVX1_LOC_292/A NOR2X1_LOC_388/Y 0.08fF
C33865 NOR2X1_LOC_590/A NAND2X1_LOC_833/Y 0.00fF
C33866 NOR2X1_LOC_174/B INVX1_LOC_53/A 0.00fF
C33867 INVX1_LOC_70/Y NAND2X1_LOC_404/a_36_24# 0.00fF
C33868 NOR2X1_LOC_451/A INVX1_LOC_92/A 0.10fF
C33869 NAND2X1_LOC_276/Y INVX1_LOC_31/A 0.17fF
C33870 NOR2X1_LOC_266/B NAND2X1_LOC_63/Y 0.35fF
C33871 NOR2X1_LOC_83/Y NOR2X1_LOC_316/a_36_216# 0.00fF
C33872 INVX1_LOC_55/Y INVX1_LOC_53/A 0.08fF
C33873 NOR2X1_LOC_583/Y INVX1_LOC_37/A 0.01fF
C33874 INVX1_LOC_9/A NAND2X1_LOC_206/Y 0.07fF
C33875 NOR2X1_LOC_471/Y INVX1_LOC_96/Y 0.02fF
C33876 INVX1_LOC_21/A INVX1_LOC_10/A 0.13fF
C33877 INVX1_LOC_186/A INVX1_LOC_271/Y 0.03fF
C33878 NOR2X1_LOC_590/A NOR2X1_LOC_182/a_36_216# 0.02fF
C33879 NOR2X1_LOC_804/B NOR2X1_LOC_703/B 0.05fF
C33880 VDD INVX1_LOC_102/A 1.41fF
C33881 NAND2X1_LOC_51/a_36_24# INPUT_7 0.00fF
C33882 INVX1_LOC_12/A NAND2X1_LOC_804/Y 0.07fF
C33883 NAND2X1_LOC_555/Y NAND2X1_LOC_141/A 0.03fF
C33884 NOR2X1_LOC_68/A INVX1_LOC_153/A 0.01fF
C33885 INVX1_LOC_61/Y NOR2X1_LOC_84/Y 0.24fF
C33886 NOR2X1_LOC_817/Y NAND2X1_LOC_563/A 0.15fF
C33887 INVX1_LOC_24/A INVX1_LOC_77/A 0.11fF
C33888 NOR2X1_LOC_598/B NOR2X1_LOC_567/B 0.12fF
C33889 INVX1_LOC_39/A D_INPUT_0 0.01fF
C33890 NOR2X1_LOC_103/Y INVX1_LOC_56/Y 0.01fF
C33891 INVX1_LOC_181/Y INVX1_LOC_33/A 0.03fF
C33892 INVX1_LOC_103/A NAND2X1_LOC_479/Y 0.02fF
C33893 NAND2X1_LOC_468/B INVX1_LOC_128/A -0.00fF
C33894 NAND2X1_LOC_357/B INVX1_LOC_72/A 0.03fF
C33895 NAND2X1_LOC_374/Y INVX1_LOC_31/A 0.07fF
C33896 NOR2X1_LOC_340/A INVX1_LOC_280/A 0.08fF
C33897 INVX1_LOC_18/A NOR2X1_LOC_377/Y 0.01fF
C33898 INVX1_LOC_223/Y NOR2X1_LOC_788/B 0.16fF
C33899 NOR2X1_LOC_288/A INVX1_LOC_305/A 0.30fF
C33900 NAND2X1_LOC_564/B INVX1_LOC_200/A 0.00fF
C33901 NAND2X1_LOC_562/B INVX1_LOC_18/A 0.01fF
C33902 NOR2X1_LOC_577/Y NOR2X1_LOC_152/Y 0.34fF
C33903 NOR2X1_LOC_41/Y INVX1_LOC_30/A 0.07fF
C33904 NOR2X1_LOC_89/A NOR2X1_LOC_376/Y 0.01fF
C33905 NOR2X1_LOC_114/A INVX1_LOC_270/A 0.20fF
C33906 INVX1_LOC_232/Y NAND2X1_LOC_577/A 0.05fF
C33907 NOR2X1_LOC_503/Y INVX1_LOC_22/A 0.00fF
C33908 INVX1_LOC_91/A INVX1_LOC_28/Y 0.01fF
C33909 NOR2X1_LOC_335/B NOR2X1_LOC_717/A 0.10fF
C33910 NAND2X1_LOC_543/Y NOR2X1_LOC_369/Y 0.05fF
C33911 NOR2X1_LOC_334/Y INVX1_LOC_76/A 0.37fF
C33912 NOR2X1_LOC_557/Y INVX1_LOC_77/A 0.03fF
C33913 INVX1_LOC_255/Y NOR2X1_LOC_160/B 0.03fF
C33914 NOR2X1_LOC_481/A NOR2X1_LOC_335/A 0.02fF
C33915 INVX1_LOC_91/A INVX1_LOC_270/A 0.10fF
C33916 NOR2X1_LOC_68/A INVX1_LOC_259/A 0.03fF
C33917 NOR2X1_LOC_816/A NOR2X1_LOC_690/Y 0.16fF
C33918 NOR2X1_LOC_510/Y NOR2X1_LOC_289/Y 0.01fF
C33919 NOR2X1_LOC_446/A INVX1_LOC_279/A 0.01fF
C33920 NAND2X1_LOC_363/B NOR2X1_LOC_334/A 0.07fF
C33921 INVX1_LOC_239/A NOR2X1_LOC_575/Y 0.13fF
C33922 NOR2X1_LOC_433/A INVX1_LOC_151/A 0.05fF
C33923 NOR2X1_LOC_269/Y NOR2X1_LOC_125/Y 0.02fF
C33924 NOR2X1_LOC_158/Y INVX1_LOC_46/A 0.03fF
C33925 NAND2X1_LOC_63/Y INVX1_LOC_46/Y 0.02fF
C33926 INVX1_LOC_45/A INVX1_LOC_56/Y 0.23fF
C33927 NOR2X1_LOC_195/A INVX1_LOC_83/A 0.04fF
C33928 INVX1_LOC_172/A NAND2X1_LOC_562/B 0.01fF
C33929 NOR2X1_LOC_478/A NOR2X1_LOC_589/A 0.07fF
C33930 INVX1_LOC_103/A INVX1_LOC_295/A 0.08fF
C33931 INVX1_LOC_21/A NAND2X1_LOC_132/a_36_24# 0.00fF
C33932 NOR2X1_LOC_773/Y INVX1_LOC_18/A 0.14fF
C33933 NOR2X1_LOC_754/A INVX1_LOC_118/A 0.03fF
C33934 INVX1_LOC_244/Y INVX1_LOC_191/Y 0.02fF
C33935 NOR2X1_LOC_433/A NOR2X1_LOC_52/B 0.47fF
C33936 NAND2X1_LOC_550/A NOR2X1_LOC_71/Y 0.01fF
C33937 NOR2X1_LOC_25/Y INVX1_LOC_46/A 0.43fF
C33938 NOR2X1_LOC_61/B NAND2X1_LOC_348/A 0.03fF
C33939 NOR2X1_LOC_565/A NOR2X1_LOC_569/Y 0.01fF
C33940 INVX1_LOC_36/A NAND2X1_LOC_712/A 0.06fF
C33941 NOR2X1_LOC_88/A INVX1_LOC_42/A 0.47fF
C33942 NOR2X1_LOC_160/B NOR2X1_LOC_71/Y 0.35fF
C33943 NAND2X1_LOC_47/a_36_24# INVX1_LOC_89/A 0.00fF
C33944 NOR2X1_LOC_791/B INVX1_LOC_16/A 0.09fF
C33945 INVX1_LOC_2/A INVX1_LOC_49/A 0.78fF
C33946 INVX1_LOC_119/A NAND2X1_LOC_325/Y 0.00fF
C33947 INVX1_LOC_77/A INVX1_LOC_143/A 0.14fF
C33948 INVX1_LOC_45/Y INVX1_LOC_208/A 0.08fF
C33949 INVX1_LOC_124/A NOR2X1_LOC_557/Y -0.00fF
C33950 INVX1_LOC_91/A NOR2X1_LOC_109/Y 0.07fF
C33951 NOR2X1_LOC_710/A INVX1_LOC_89/A 0.01fF
C33952 INVX1_LOC_174/A NOR2X1_LOC_163/A 0.04fF
C33953 NOR2X1_LOC_68/A NOR2X1_LOC_589/A 0.08fF
C33954 NOR2X1_LOC_134/Y INPUT_1 0.06fF
C33955 INVX1_LOC_159/A NAND2X1_LOC_662/Y 0.73fF
C33956 NAND2X1_LOC_715/B NOR2X1_LOC_269/Y 0.05fF
C33957 INVX1_LOC_103/A NOR2X1_LOC_202/Y 0.01fF
C33958 NOR2X1_LOC_644/A NOR2X1_LOC_160/B 0.07fF
C33959 INVX1_LOC_172/A NOR2X1_LOC_773/Y 0.05fF
C33960 NOR2X1_LOC_586/a_36_216# INVX1_LOC_72/A 0.00fF
C33961 VDD INVX1_LOC_296/Y 0.19fF
C33962 NAND2X1_LOC_569/a_36_24# NOR2X1_LOC_130/A 0.01fF
C33963 NOR2X1_LOC_590/A NOR2X1_LOC_180/B 0.07fF
C33964 INVX1_LOC_32/A INVX1_LOC_92/A 0.10fF
C33965 NOR2X1_LOC_718/B NAND2X1_LOC_629/Y 0.01fF
C33966 NOR2X1_LOC_647/Y NOR2X1_LOC_332/A -0.02fF
C33967 NOR2X1_LOC_828/B NOR2X1_LOC_160/B 0.03fF
C33968 NOR2X1_LOC_152/Y INVX1_LOC_22/A 2.61fF
C33969 INVX1_LOC_314/Y NOR2X1_LOC_397/a_36_216# 0.00fF
C33970 NOR2X1_LOC_288/A NAND2X1_LOC_690/a_36_24# 0.01fF
C33971 NOR2X1_LOC_279/a_36_216# NOR2X1_LOC_309/Y 0.01fF
C33972 INVX1_LOC_272/A INVX1_LOC_19/A 0.07fF
C33973 INVX1_LOC_49/A NOR2X1_LOC_161/Y 0.01fF
C33974 INVX1_LOC_113/Y INVX1_LOC_22/A 0.09fF
C33975 INVX1_LOC_105/A INVX1_LOC_290/A 0.02fF
C33976 NOR2X1_LOC_544/A NOR2X1_LOC_147/B 0.09fF
C33977 NOR2X1_LOC_488/Y NAND2X1_LOC_833/Y 0.01fF
C33978 INVX1_LOC_276/A INVX1_LOC_119/A 0.01fF
C33979 D_INPUT_0 INVX1_LOC_61/A 0.12fF
C33980 INVX1_LOC_269/A INVX1_LOC_286/A 0.10fF
C33981 NOR2X1_LOC_861/Y NAND2X1_LOC_206/Y 0.05fF
C33982 NOR2X1_LOC_590/A INVX1_LOC_73/A 0.03fF
C33983 NAND2X1_LOC_53/Y INVX1_LOC_311/A 0.98fF
C33984 INVX1_LOC_124/A INVX1_LOC_143/A 0.00fF
C33985 NOR2X1_LOC_473/B INVX1_LOC_177/Y 0.10fF
C33986 NOR2X1_LOC_160/B NOR2X1_LOC_751/A 0.01fF
C33987 NAND2X1_LOC_175/Y INVX1_LOC_92/A 0.08fF
C33988 INVX1_LOC_209/Y NOR2X1_LOC_561/Y 0.11fF
C33989 INVX1_LOC_289/Y NOR2X1_LOC_45/B 0.01fF
C33990 NOR2X1_LOC_525/Y NOR2X1_LOC_484/Y 0.00fF
C33991 NOR2X1_LOC_124/B INVX1_LOC_16/A 0.03fF
C33992 INVX1_LOC_2/A NOR2X1_LOC_226/A 0.09fF
C33993 NAND2X1_LOC_529/a_36_24# NOR2X1_LOC_548/B 0.02fF
C33994 NOR2X1_LOC_717/A NOR2X1_LOC_440/a_36_216# 0.00fF
C33995 NOR2X1_LOC_721/A NOR2X1_LOC_346/B 0.01fF
C33996 NOR2X1_LOC_590/A NOR2X1_LOC_569/A 0.04fF
C33997 NAND2X1_LOC_113/a_36_24# NOR2X1_LOC_188/A 0.00fF
C33998 NAND2X1_LOC_500/Y INVX1_LOC_91/Y 0.07fF
C33999 NOR2X1_LOC_773/Y NOR2X1_LOC_709/a_36_216# 0.00fF
C34000 INVX1_LOC_18/A INVX1_LOC_140/A 0.12fF
C34001 INVX1_LOC_304/Y NAND2X1_LOC_564/B -0.01fF
C34002 INVX1_LOC_36/A INVX1_LOC_79/A 0.13fF
C34003 INVX1_LOC_292/A NOR2X1_LOC_794/A 0.03fF
C34004 INVX1_LOC_30/Y NOR2X1_LOC_315/Y 0.10fF
C34005 INVX1_LOC_21/A INVX1_LOC_178/Y 0.03fF
C34006 INVX1_LOC_273/Y NAND2X1_LOC_354/B 0.01fF
C34007 NOR2X1_LOC_250/a_36_216# NOR2X1_LOC_405/A 0.02fF
C34008 INVX1_LOC_262/A INVX1_LOC_92/A 0.03fF
C34009 NOR2X1_LOC_767/a_36_216# INVX1_LOC_16/A 0.00fF
C34010 NOR2X1_LOC_89/A NOR2X1_LOC_159/a_36_216# 0.00fF
C34011 INVX1_LOC_89/A NOR2X1_LOC_520/B 0.16fF
C34012 INVX1_LOC_29/A D_INPUT_5 0.00fF
C34013 NOR2X1_LOC_667/a_36_216# INVX1_LOC_91/A 0.01fF
C34014 NAND2X1_LOC_96/A INVX1_LOC_50/Y 0.07fF
C34015 NOR2X1_LOC_109/Y NAND2X1_LOC_783/a_36_24# 0.01fF
C34016 INVX1_LOC_11/A NOR2X1_LOC_601/Y 0.03fF
C34017 INVX1_LOC_213/Y NOR2X1_LOC_717/B 0.00fF
C34018 INVX1_LOC_36/A INVX1_LOC_309/A 0.03fF
C34019 INVX1_LOC_256/A NOR2X1_LOC_657/B 0.04fF
C34020 NOR2X1_LOC_828/A NOR2X1_LOC_551/B 0.00fF
C34021 INVX1_LOC_13/A NOR2X1_LOC_547/B 0.03fF
C34022 INVX1_LOC_78/A INVX1_LOC_186/Y 0.07fF
C34023 INVX1_LOC_313/Y NOR2X1_LOC_344/A 0.03fF
C34024 INVX1_LOC_13/A NOR2X1_LOC_78/B 0.42fF
C34025 NAND2X1_LOC_374/Y NAND2X1_LOC_859/Y 0.10fF
C34026 INVX1_LOC_41/A INVX1_LOC_196/Y 0.03fF
C34027 INVX1_LOC_172/A INVX1_LOC_140/A 0.07fF
C34028 INVX1_LOC_11/A INVX1_LOC_74/A 0.19fF
C34029 NAND2X1_LOC_213/A INVX1_LOC_37/A 0.01fF
C34030 INVX1_LOC_224/Y NOR2X1_LOC_179/a_36_216# 0.01fF
C34031 NAND2X1_LOC_500/Y NOR2X1_LOC_45/B 0.01fF
C34032 INVX1_LOC_223/A NOR2X1_LOC_337/Y 0.34fF
C34033 NOR2X1_LOC_216/Y INVX1_LOC_77/A 0.12fF
C34034 NAND2X1_LOC_381/Y INVX1_LOC_74/A 0.28fF
C34035 INVX1_LOC_27/A NOR2X1_LOC_536/A 0.29fF
C34036 INVX1_LOC_24/A NAND2X1_LOC_832/Y 0.06fF
C34037 NOR2X1_LOC_773/Y NOR2X1_LOC_690/Y 0.02fF
C34038 INVX1_LOC_251/Y INVX1_LOC_306/A 0.01fF
C34039 INVX1_LOC_213/Y NOR2X1_LOC_828/A 0.00fF
C34040 NOR2X1_LOC_824/A NOR2X1_LOC_536/A 0.07fF
C34041 NOR2X1_LOC_667/A INVX1_LOC_10/A 0.03fF
C34042 NOR2X1_LOC_473/B INVX1_LOC_104/A 0.10fF
C34043 INVX1_LOC_116/A NOR2X1_LOC_188/A 0.27fF
C34044 INVX1_LOC_255/Y NOR2X1_LOC_516/B 2.51fF
C34045 INVX1_LOC_36/A INVX1_LOC_91/A 0.39fF
C34046 NOR2X1_LOC_112/B INVX1_LOC_77/A 0.02fF
C34047 INVX1_LOC_207/A NAND2X1_LOC_560/A 0.04fF
C34048 NAND2X1_LOC_575/a_36_24# INVX1_LOC_33/Y 0.00fF
C34049 INVX1_LOC_2/A NAND2X1_LOC_648/A 0.03fF
C34050 NOR2X1_LOC_500/Y NOR2X1_LOC_565/B 0.02fF
C34051 INVX1_LOC_93/A INVX1_LOC_185/A 0.03fF
C34052 INVX1_LOC_2/A INPUT_1 0.04fF
C34053 NOR2X1_LOC_67/A INVX1_LOC_89/A 0.18fF
C34054 INPUT_2 VDD 0.20fF
C34055 INVX1_LOC_245/Y INVX1_LOC_14/Y 0.03fF
C34056 INVX1_LOC_36/A INVX1_LOC_11/Y 0.06fF
C34057 NOR2X1_LOC_837/Y NOR2X1_LOC_837/A 0.00fF
C34058 INVX1_LOC_27/A NOR2X1_LOC_655/Y 0.10fF
C34059 NAND2X1_LOC_361/Y NOR2X1_LOC_188/A 0.03fF
C34060 NAND2X1_LOC_374/Y NAND2X1_LOC_866/B 0.04fF
C34061 NAND2X1_LOC_35/Y INVX1_LOC_260/Y 0.01fF
C34062 NOR2X1_LOC_226/A INPUT_1 0.80fF
C34063 INVX1_LOC_213/Y NOR2X1_LOC_151/Y 0.35fF
C34064 INVX1_LOC_41/A NOR2X1_LOC_292/Y 0.01fF
C34065 INVX1_LOC_84/A NOR2X1_LOC_717/A 0.10fF
C34066 NAND2X1_LOC_361/Y NOR2X1_LOC_548/B 0.10fF
C34067 NOR2X1_LOC_78/B INVX1_LOC_55/Y 0.04fF
C34068 NOR2X1_LOC_717/B NAND2X1_LOC_513/a_36_24# 0.00fF
C34069 INVX1_LOC_145/A INVX1_LOC_91/A 0.03fF
C34070 INVX1_LOC_27/A NAND2X1_LOC_93/B 0.95fF
C34071 INVX1_LOC_124/A NOR2X1_LOC_216/Y 0.13fF
C34072 INVX1_LOC_21/A INVX1_LOC_307/A 0.07fF
C34073 INVX1_LOC_39/A INVX1_LOC_46/Y 0.04fF
C34074 D_INPUT_0 NOR2X1_LOC_85/a_36_216# 0.00fF
C34075 INVX1_LOC_13/A INVX1_LOC_83/A 0.07fF
C34076 INVX1_LOC_268/A NOR2X1_LOC_207/a_36_216# 0.01fF
C34077 NAND2X1_LOC_276/Y INVX1_LOC_6/A 0.04fF
C34078 D_INPUT_1 NAND2X1_LOC_82/Y 0.11fF
C34079 INVX1_LOC_269/A INVX1_LOC_54/A 0.10fF
C34080 INVX1_LOC_21/A NOR2X1_LOC_445/B 0.12fF
C34081 NAND2X1_LOC_733/Y NAND2X1_LOC_804/Y 0.43fF
C34082 NAND2X1_LOC_783/A NAND2X1_LOC_796/Y 0.05fF
C34083 NOR2X1_LOC_644/A NOR2X1_LOC_516/B 0.03fF
C34084 NAND2X1_LOC_214/B INVX1_LOC_3/A 0.06fF
C34085 NOR2X1_LOC_68/A INVX1_LOC_20/A 0.06fF
C34086 NOR2X1_LOC_540/a_36_216# INVX1_LOC_313/Y 0.00fF
C34087 INVX1_LOC_145/Y NOR2X1_LOC_355/A 0.06fF
C34088 NOR2X1_LOC_804/B INVX1_LOC_91/A 0.09fF
C34089 NAND2X1_LOC_571/Y INVX1_LOC_260/Y 0.03fF
C34090 NOR2X1_LOC_68/A NOR2X1_LOC_360/A 0.01fF
C34091 NOR2X1_LOC_666/A NOR2X1_LOC_155/A 0.21fF
C34092 NAND2X1_LOC_787/A NAND2X1_LOC_74/B 0.02fF
C34093 NOR2X1_LOC_337/Y INVX1_LOC_149/Y 0.11fF
C34094 NAND2X1_LOC_758/a_36_24# INVX1_LOC_76/A 0.01fF
C34095 INVX1_LOC_190/A NOR2X1_LOC_130/A 0.02fF
C34096 NAND2X1_LOC_332/Y NOR2X1_LOC_45/B 0.07fF
C34097 INVX1_LOC_94/Y INVX1_LOC_273/A 0.02fF
C34098 NAND2X1_LOC_364/A INVX1_LOC_37/A 0.12fF
C34099 NAND2X1_LOC_363/B NAND2X1_LOC_74/B 0.07fF
C34100 NAND2X1_LOC_364/A NOR2X1_LOC_231/A 0.03fF
C34101 INVX1_LOC_27/A INVX1_LOC_3/A 1.50fF
C34102 NOR2X1_LOC_38/B INVX1_LOC_23/Y 0.10fF
C34103 NOR2X1_LOC_355/B INVX1_LOC_104/A 0.03fF
C34104 INVX1_LOC_135/A INVX1_LOC_120/A 0.03fF
C34105 NOR2X1_LOC_78/B NOR2X1_LOC_320/Y 0.02fF
C34106 NOR2X1_LOC_598/B NOR2X1_LOC_633/a_36_216# 0.01fF
C34107 INVX1_LOC_217/A NAND2X1_LOC_804/Y 0.73fF
C34108 NOR2X1_LOC_134/Y INVX1_LOC_118/A 0.08fF
C34109 NOR2X1_LOC_727/B INVX1_LOC_15/A 0.03fF
C34110 INVX1_LOC_83/A NOR2X1_LOC_174/B 0.03fF
C34111 INVX1_LOC_75/A NAND2X1_LOC_671/a_36_24# 0.00fF
C34112 INVX1_LOC_73/A NOR2X1_LOC_82/Y 0.03fF
C34113 NOR2X1_LOC_721/B NOR2X1_LOC_849/A 0.03fF
C34114 NOR2X1_LOC_309/Y INVX1_LOC_91/A 0.03fF
C34115 NAND2X1_LOC_549/Y INVX1_LOC_284/A 0.00fF
C34116 NOR2X1_LOC_172/Y NAND2X1_LOC_468/B 0.00fF
C34117 NAND2X1_LOC_374/Y INVX1_LOC_6/A 0.07fF
C34118 NOR2X1_LOC_778/B INVX1_LOC_69/Y 0.08fF
C34119 NOR2X1_LOC_368/A INVX1_LOC_56/A 0.01fF
C34120 INVX1_LOC_88/A NOR2X1_LOC_841/A 0.01fF
C34121 NAND2X1_LOC_3/B NAND2X1_LOC_64/a_36_24# -0.00fF
C34122 NAND2X1_LOC_656/A INVX1_LOC_129/Y 0.52fF
C34123 INVX1_LOC_209/Y INVX1_LOC_76/A 0.06fF
C34124 INVX1_LOC_120/A NOR2X1_LOC_560/A 0.02fF
C34125 NOR2X1_LOC_791/Y NAND2X1_LOC_74/B 1.28fF
C34126 INVX1_LOC_61/A NAND2X1_LOC_848/A 0.04fF
C34127 INVX1_LOC_227/A INVX1_LOC_73/A 0.07fF
C34128 INVX1_LOC_53/A INVX1_LOC_32/A 0.21fF
C34129 NOR2X1_LOC_315/Y NOR2X1_LOC_124/A 0.03fF
C34130 INVX1_LOC_196/A NOR2X1_LOC_78/A 0.54fF
C34131 NOR2X1_LOC_52/B INVX1_LOC_199/A 0.01fF
C34132 NAND2X1_LOC_833/Y NAND2X1_LOC_650/B 0.10fF
C34133 NOR2X1_LOC_717/A INVX1_LOC_15/A 0.00fF
C34134 NOR2X1_LOC_312/Y NOR2X1_LOC_329/B 0.01fF
C34135 NOR2X1_LOC_559/B NAND2X1_LOC_96/A 0.02fF
C34136 INVX1_LOC_21/A INVX1_LOC_12/A 0.10fF
C34137 D_INPUT_6 NOR2X1_LOC_17/a_36_216# 0.00fF
C34138 NAND2X1_LOC_787/B NAND2X1_LOC_804/Y 0.01fF
C34139 NOR2X1_LOC_613/a_36_216# NOR2X1_LOC_89/A 0.00fF
C34140 NAND2X1_LOC_181/Y INVX1_LOC_70/Y 0.01fF
C34141 INVX1_LOC_24/A INVX1_LOC_9/A 20.95fF
C34142 VDD INVX1_LOC_149/Y 0.34fF
C34143 NOR2X1_LOC_191/A NAND2X1_LOC_642/Y 0.17fF
C34144 NOR2X1_LOC_789/A INVX1_LOC_123/A 0.03fF
C34145 INVX1_LOC_162/Y VDD 0.47fF
C34146 NAND2X1_LOC_394/a_36_24# INVX1_LOC_32/A 0.00fF
C34147 NOR2X1_LOC_455/Y NOR2X1_LOC_334/Y -0.04fF
C34148 INVX1_LOC_45/A NOR2X1_LOC_831/B 0.11fF
C34149 NOR2X1_LOC_740/Y INVX1_LOC_19/A 0.07fF
C34150 INVX1_LOC_255/Y INVX1_LOC_315/Y 0.01fF
C34151 NOR2X1_LOC_52/Y INVX1_LOC_117/Y 0.00fF
C34152 NAND2X1_LOC_364/A NOR2X1_LOC_743/Y 0.10fF
C34153 INVX1_LOC_265/A NAND2X1_LOC_721/A 0.44fF
C34154 INVX1_LOC_230/Y NOR2X1_LOC_23/a_36_216# 0.01fF
C34155 INVX1_LOC_85/A VDD 0.00fF
C34156 NOR2X1_LOC_788/B INVX1_LOC_75/A 0.07fF
C34157 NOR2X1_LOC_568/A NOR2X1_LOC_831/B 0.00fF
C34158 INVX1_LOC_53/A NAND2X1_LOC_175/Y 0.07fF
C34159 INVX1_LOC_17/A INVX1_LOC_49/Y 0.08fF
C34160 NOR2X1_LOC_309/Y NOR2X1_LOC_653/a_36_216# 0.01fF
C34161 NOR2X1_LOC_316/Y VDD 0.11fF
C34162 INPUT_0 NOR2X1_LOC_72/a_36_216# 0.00fF
C34163 INVX1_LOC_64/A NAND2X1_LOC_454/Y 0.17fF
C34164 NAND2X1_LOC_35/Y NAND2X1_LOC_471/Y 0.01fF
C34165 INVX1_LOC_150/Y INVX1_LOC_19/A 0.05fF
C34166 NOR2X1_LOC_276/B NOR2X1_LOC_155/A 0.01fF
C34167 INVX1_LOC_57/A NOR2X1_LOC_383/B 10.16fF
C34168 INVX1_LOC_304/Y NAND2X1_LOC_804/Y 0.00fF
C34169 INVX1_LOC_279/A INVX1_LOC_186/A 0.07fF
C34170 INVX1_LOC_214/Y NOR2X1_LOC_173/a_36_216# 0.00fF
C34171 INVX1_LOC_49/A INVX1_LOC_118/A 0.03fF
C34172 NOR2X1_LOC_6/B NAND2X1_LOC_96/A 0.01fF
C34173 NOR2X1_LOC_78/B NOR2X1_LOC_357/Y 0.07fF
C34174 INVX1_LOC_35/A NOR2X1_LOC_278/Y 0.03fF
C34175 INVX1_LOC_249/A NAND2X1_LOC_93/B 0.03fF
C34176 NOR2X1_LOC_488/Y NAND2X1_LOC_241/Y 0.04fF
C34177 NAND2X1_LOC_11/Y INVX1_LOC_37/A 0.09fF
C34178 NOR2X1_LOC_577/Y INVX1_LOC_291/A 0.13fF
C34179 INVX1_LOC_136/A NAND2X1_LOC_475/Y 1.01fF
C34180 INVX1_LOC_41/A NOR2X1_LOC_641/Y 0.02fF
C34181 INVX1_LOC_31/A INVX1_LOC_125/A 0.10fF
C34182 INVX1_LOC_71/A NOR2X1_LOC_831/B 0.07fF
C34183 NAND2X1_LOC_799/A INVX1_LOC_42/A 0.03fF
C34184 INVX1_LOC_57/Y NOR2X1_LOC_662/A 0.10fF
C34185 INVX1_LOC_311/A NOR2X1_LOC_302/Y 0.05fF
C34186 NOR2X1_LOC_703/B INVX1_LOC_63/A 0.03fF
C34187 INVX1_LOC_77/A NOR2X1_LOC_197/B 0.01fF
C34188 NOR2X1_LOC_103/Y NAND2X1_LOC_74/a_36_24# 0.00fF
C34189 NOR2X1_LOC_647/A INVX1_LOC_5/A 0.32fF
C34190 NAND2X1_LOC_24/a_36_24# NOR2X1_LOC_35/Y 0.01fF
C34191 INVX1_LOC_279/A NAND2X1_LOC_447/Y 0.01fF
C34192 NOR2X1_LOC_360/Y NOR2X1_LOC_673/B 0.01fF
C34193 INVX1_LOC_69/Y NAND2X1_LOC_123/Y 0.09fF
C34194 NAND2X1_LOC_543/Y VDD 0.01fF
C34195 NOR2X1_LOC_817/Y NOR2X1_LOC_554/A 0.02fF
C34196 NOR2X1_LOC_78/B NOR2X1_LOC_319/B 6.65fF
C34197 NOR2X1_LOC_328/Y NOR2X1_LOC_447/B 0.03fF
C34198 INVX1_LOC_47/A NOR2X1_LOC_78/A 0.01fF
C34199 INVX1_LOC_135/A NOR2X1_LOC_542/B 0.02fF
C34200 INVX1_LOC_90/A NAND2X1_LOC_655/A 0.07fF
C34201 INVX1_LOC_110/Y NAND2X1_LOC_206/B 0.10fF
C34202 NAND2X1_LOC_662/Y VDD 0.22fF
C34203 INVX1_LOC_13/A INVX1_LOC_46/A 0.00fF
C34204 NOR2X1_LOC_589/A NOR2X1_LOC_364/a_36_216# 0.02fF
C34205 INVX1_LOC_63/Y NAND2X1_LOC_798/B 0.02fF
C34206 INVX1_LOC_30/A NAND2X1_LOC_74/B 6.47fF
C34207 NOR2X1_LOC_730/Y VDD 0.24fF
C34208 INVX1_LOC_13/A NOR2X1_LOC_98/A 0.01fF
C34209 INVX1_LOC_16/A INVX1_LOC_37/Y 0.02fF
C34210 INVX1_LOC_88/A INVX1_LOC_128/A 0.01fF
C34211 INVX1_LOC_2/A INVX1_LOC_118/A 0.37fF
C34212 INVX1_LOC_143/A INVX1_LOC_9/A 0.08fF
C34213 NOR2X1_LOC_363/Y INVX1_LOC_16/A 0.07fF
C34214 NOR2X1_LOC_806/Y NOR2X1_LOC_856/A 0.02fF
C34215 NOR2X1_LOC_643/Y NOR2X1_LOC_673/A 0.03fF
C34216 NOR2X1_LOC_430/A INVX1_LOC_84/A 0.13fF
C34217 INVX1_LOC_41/A NOR2X1_LOC_461/B 0.14fF
C34218 NOR2X1_LOC_226/A INVX1_LOC_118/A 0.18fF
C34219 NAND2X1_LOC_551/A NOR2X1_LOC_368/Y 0.05fF
C34220 NAND2X1_LOC_99/Y INVX1_LOC_3/A 0.02fF
C34221 NAND2X1_LOC_354/Y INVX1_LOC_12/A 0.12fF
C34222 INVX1_LOC_206/A NAND2X1_LOC_93/B 0.04fF
C34223 NOR2X1_LOC_360/Y INVX1_LOC_29/A 0.01fF
C34224 NOR2X1_LOC_647/Y NOR2X1_LOC_847/A 0.27fF
C34225 INVX1_LOC_90/A NOR2X1_LOC_683/Y 0.02fF
C34226 NOR2X1_LOC_620/Y NOR2X1_LOC_814/A 0.01fF
C34227 NOR2X1_LOC_237/Y INVX1_LOC_203/A 0.00fF
C34228 INVX1_LOC_68/Y INVX1_LOC_9/A 0.01fF
C34229 D_INPUT_0 D_INPUT_3 2.63fF
C34230 NOR2X1_LOC_785/a_36_216# NOR2X1_LOC_78/A 0.00fF
C34231 NOR2X1_LOC_384/a_36_216# INVX1_LOC_42/A 0.02fF
C34232 INVX1_LOC_224/Y NOR2X1_LOC_789/B 0.01fF
C34233 NAND2X1_LOC_784/A NOR2X1_LOC_406/A 0.08fF
C34234 NOR2X1_LOC_246/A INVX1_LOC_46/A 0.07fF
C34235 NAND2X1_LOC_799/A INVX1_LOC_78/A 0.00fF
C34236 D_INPUT_2 NAND2X1_LOC_82/Y 0.02fF
C34237 INVX1_LOC_113/Y INVX1_LOC_186/Y 0.00fF
C34238 INVX1_LOC_18/A INVX1_LOC_42/A 0.28fF
C34239 INVX1_LOC_40/Y INVX1_LOC_3/Y 0.26fF
C34240 NOR2X1_LOC_763/A INVX1_LOC_57/A 0.02fF
C34241 NOR2X1_LOC_437/Y INVX1_LOC_272/A 0.05fF
C34242 NOR2X1_LOC_15/Y INVX1_LOC_181/A 0.03fF
C34243 NAND2X1_LOC_551/A INVX1_LOC_46/A 0.01fF
C34244 INVX1_LOC_234/A NOR2X1_LOC_536/A 0.01fF
C34245 INVX1_LOC_182/Y NAND2X1_LOC_447/Y 0.03fF
C34246 INVX1_LOC_49/A NAND2X1_LOC_63/Y 0.01fF
C34247 NOR2X1_LOC_666/Y NOR2X1_LOC_383/B 0.65fF
C34248 INVX1_LOC_50/A INVX1_LOC_1/A 0.10fF
C34249 INVX1_LOC_174/A NOR2X1_LOC_36/A 0.10fF
C34250 INVX1_LOC_55/Y INVX1_LOC_46/A 0.11fF
C34251 INVX1_LOC_83/A NOR2X1_LOC_319/B 0.00fF
C34252 INVX1_LOC_314/Y NOR2X1_LOC_89/A 0.14fF
C34253 NAND2X1_LOC_860/A NOR2X1_LOC_440/B 0.01fF
C34254 NAND2X1_LOC_859/B NOR2X1_LOC_88/A 0.12fF
C34255 INVX1_LOC_269/A NAND2X1_LOC_215/A 0.01fF
C34256 NOR2X1_LOC_860/B NOR2X1_LOC_346/A 0.03fF
C34257 NAND2X1_LOC_570/Y NOR2X1_LOC_649/B 0.03fF
C34258 INVX1_LOC_22/A NAND2X1_LOC_802/Y 0.07fF
C34259 NOR2X1_LOC_708/B NAND2X1_LOC_782/a_36_24# 0.00fF
C34260 INVX1_LOC_137/A NAND2X1_LOC_93/B 0.49fF
C34261 NOR2X1_LOC_791/a_36_216# INVX1_LOC_3/Y 0.00fF
C34262 NOR2X1_LOC_68/A INVX1_LOC_4/A 0.07fF
C34263 NOR2X1_LOC_336/B NAND2X1_LOC_72/B 0.02fF
C34264 NAND2X1_LOC_717/Y NOR2X1_LOC_485/Y 0.02fF
C34265 INVX1_LOC_172/A INVX1_LOC_42/A 0.18fF
C34266 INVX1_LOC_28/A INVX1_LOC_37/Y 0.01fF
C34267 NAND2X1_LOC_840/Y NOR2X1_LOC_305/Y 0.03fF
C34268 INVX1_LOC_28/A NOR2X1_LOC_363/Y 0.07fF
C34269 GATE_662 INVX1_LOC_92/A 0.01fF
C34270 NOR2X1_LOC_561/Y NAND2X1_LOC_434/Y 0.05fF
C34271 INVX1_LOC_222/Y INVX1_LOC_50/Y 0.03fF
C34272 INVX1_LOC_256/A INVX1_LOC_271/A 0.04fF
C34273 NOR2X1_LOC_13/Y INVX1_LOC_15/A 0.10fF
C34274 NOR2X1_LOC_792/B INVX1_LOC_29/A 0.01fF
C34275 INVX1_LOC_33/A NOR2X1_LOC_114/Y 0.31fF
C34276 INVX1_LOC_18/A INVX1_LOC_78/A 6.83fF
C34277 INVX1_LOC_184/A NOR2X1_LOC_623/B 0.02fF
C34278 NAND2X1_LOC_785/Y INVX1_LOC_12/A 0.06fF
C34279 INVX1_LOC_130/Y NAND2X1_LOC_454/Y 0.01fF
C34280 INVX1_LOC_73/Y NOR2X1_LOC_678/A 0.00fF
C34281 NOR2X1_LOC_214/B INVX1_LOC_54/A 0.04fF
C34282 NOR2X1_LOC_320/Y INVX1_LOC_46/A 0.05fF
C34283 NOR2X1_LOC_160/B NAND2X1_LOC_205/A 1.11fF
C34284 NOR2X1_LOC_19/B NOR2X1_LOC_536/A 0.03fF
C34285 INPUT_1 INVX1_LOC_118/A 0.08fF
C34286 INVX1_LOC_95/Y INVX1_LOC_98/A 0.15fF
C34287 INVX1_LOC_2/A NAND2X1_LOC_63/Y 0.03fF
C34288 INVX1_LOC_21/A NOR2X1_LOC_34/A 0.04fF
C34289 NOR2X1_LOC_790/B NOR2X1_LOC_541/Y 0.10fF
C34290 INVX1_LOC_95/Y NOR2X1_LOC_78/A 0.08fF
C34291 NOR2X1_LOC_590/Y INVX1_LOC_1/A 0.00fF
C34292 NOR2X1_LOC_577/Y NOR2X1_LOC_609/Y 0.03fF
C34293 INVX1_LOC_137/A INVX1_LOC_3/A 0.06fF
C34294 NOR2X1_LOC_52/B NAND2X1_LOC_254/Y 0.03fF
C34295 NAND2X1_LOC_451/Y INVX1_LOC_29/A 0.05fF
C34296 NOR2X1_LOC_226/A NAND2X1_LOC_63/Y 0.02fF
C34297 INVX1_LOC_14/A INVX1_LOC_306/Y 0.32fF
C34298 INVX1_LOC_222/Y INVX1_LOC_266/A 0.01fF
C34299 INVX1_LOC_277/A NOR2X1_LOC_858/A 0.01fF
C34300 NOR2X1_LOC_554/B NOR2X1_LOC_843/B 0.09fF
C34301 NOR2X1_LOC_216/Y INVX1_LOC_9/A 0.10fF
C34302 NOR2X1_LOC_65/B INVX1_LOC_18/A 0.10fF
C34303 NOR2X1_LOC_600/Y NAND2X1_LOC_602/a_36_24# 0.00fF
C34304 INVX1_LOC_62/Y INVX1_LOC_23/Y 0.30fF
C34305 NOR2X1_LOC_667/A INVX1_LOC_12/A 5.10fF
C34306 NAND2X1_LOC_591/a_36_24# NOR2X1_LOC_727/B 0.00fF
C34307 INVX1_LOC_57/Y INVX1_LOC_57/A 0.27fF
C34308 INVX1_LOC_286/A INVX1_LOC_12/Y 0.10fF
C34309 NOR2X1_LOC_19/B NOR2X1_LOC_655/Y 0.80fF
C34310 INVX1_LOC_172/A INVX1_LOC_78/A 0.03fF
C34311 INVX1_LOC_34/Y INVX1_LOC_42/A 0.01fF
C34312 INVX1_LOC_234/A INVX1_LOC_3/A 0.03fF
C34313 INVX1_LOC_7/A NAND2X1_LOC_206/Y 0.04fF
C34314 NOR2X1_LOC_415/a_36_216# NAND2X1_LOC_574/A 0.01fF
C34315 INVX1_LOC_135/A NAND2X1_LOC_659/A 0.15fF
C34316 INVX1_LOC_280/Y INVX1_LOC_102/A 0.38fF
C34317 INVX1_LOC_45/A NOR2X1_LOC_790/B 0.07fF
C34318 NOR2X1_LOC_454/Y NOR2X1_LOC_470/B 0.14fF
C34319 NOR2X1_LOC_67/A NOR2X1_LOC_490/a_36_216# 0.00fF
C34320 NAND2X1_LOC_569/B INVX1_LOC_31/A 0.09fF
C34321 NAND2X1_LOC_729/Y INVX1_LOC_50/A 0.03fF
C34322 INVX1_LOC_21/A INVX1_LOC_200/A 0.03fF
C34323 NAND2X1_LOC_53/Y NOR2X1_LOC_626/Y 0.02fF
C34324 INVX1_LOC_49/A NOR2X1_LOC_631/Y 0.02fF
C34325 INVX1_LOC_7/A NAND2X1_LOC_773/B 0.18fF
C34326 INVX1_LOC_136/A NAND2X1_LOC_787/A 0.03fF
C34327 INVX1_LOC_256/A INVX1_LOC_27/A 0.72fF
C34328 INVX1_LOC_34/A NOR2X1_LOC_30/Y 0.00fF
C34329 NAND2X1_LOC_465/Y NAND2X1_LOC_471/Y 0.05fF
C34330 NOR2X1_LOC_464/a_36_216# INVX1_LOC_271/Y 0.00fF
C34331 INVX1_LOC_136/A NAND2X1_LOC_363/B 0.01fF
C34332 NOR2X1_LOC_647/B INVX1_LOC_27/A 0.03fF
C34333 INVX1_LOC_314/A VDD 0.12fF
C34334 NAND2X1_LOC_214/B NOR2X1_LOC_606/Y 0.01fF
C34335 NOR2X1_LOC_78/B INVX1_LOC_32/A 0.79fF
C34336 INVX1_LOC_39/A NOR2X1_LOC_134/Y 0.02fF
C34337 NOR2X1_LOC_173/Y NOR2X1_LOC_816/A 0.09fF
C34338 NOR2X1_LOC_703/Y NOR2X1_LOC_729/A 3.05fF
C34339 INVX1_LOC_183/Y INVX1_LOC_63/A 0.01fF
C34340 INVX1_LOC_2/Y NOR2X1_LOC_35/Y 0.38fF
C34341 INVX1_LOC_86/Y INVX1_LOC_193/A -0.01fF
C34342 NAND2X1_LOC_813/a_36_24# NOR2X1_LOC_536/A 0.00fF
C34343 NAND2X1_LOC_800/a_36_24# NAND2X1_LOC_800/A 0.00fF
C34344 INVX1_LOC_304/A NOR2X1_LOC_301/a_36_216# 0.01fF
C34345 INVX1_LOC_64/A NOR2X1_LOC_68/A 0.20fF
C34346 INVX1_LOC_136/A NAND2X1_LOC_565/a_36_24# 0.01fF
C34347 NOR2X1_LOC_19/B NOR2X1_LOC_649/B 0.24fF
C34348 INVX1_LOC_195/A INVX1_LOC_253/Y 0.00fF
C34349 NOR2X1_LOC_758/Y NAND2X1_LOC_286/B 0.04fF
C34350 NAND2X1_LOC_655/A INVX1_LOC_38/A 0.21fF
C34351 NOR2X1_LOC_19/B INVX1_LOC_3/A 0.22fF
C34352 NOR2X1_LOC_357/Y INVX1_LOC_46/A 0.19fF
C34353 NOR2X1_LOC_632/Y INVX1_LOC_283/A 0.02fF
C34354 INVX1_LOC_27/A NOR2X1_LOC_606/Y 0.08fF
C34355 INVX1_LOC_5/A INVX1_LOC_205/A 0.00fF
C34356 INVX1_LOC_144/A NOR2X1_LOC_832/a_36_216# 0.01fF
C34357 NOR2X1_LOC_790/B INVX1_LOC_71/A 0.01fF
C34358 NOR2X1_LOC_446/A NAND2X1_LOC_190/Y 0.05fF
C34359 INVX1_LOC_37/A NOR2X1_LOC_857/A 0.98fF
C34360 INVX1_LOC_31/A NAND2X1_LOC_218/A 0.01fF
C34361 INVX1_LOC_136/A NOR2X1_LOC_791/Y 0.11fF
C34362 NOR2X1_LOC_140/A INVX1_LOC_31/A 0.07fF
C34363 NAND2X1_LOC_1/a_36_24# INPUT_7 0.00fF
C34364 INVX1_LOC_1/A INVX1_LOC_61/Y 0.10fF
C34365 INVX1_LOC_232/A NOR2X1_LOC_38/B 0.07fF
C34366 NAND2X1_LOC_468/B INVX1_LOC_38/A 0.10fF
C34367 NAND2X1_LOC_231/Y NOR2X1_LOC_301/A 0.01fF
C34368 NOR2X1_LOC_635/A INVX1_LOC_296/A 0.01fF
C34369 NOR2X1_LOC_78/B NAND2X1_LOC_175/Y 0.08fF
C34370 NAND2X1_LOC_840/B INVX1_LOC_94/Y 0.07fF
C34371 NOR2X1_LOC_570/Y INVX1_LOC_4/A 0.03fF
C34372 NAND2X1_LOC_799/A NOR2X1_LOC_503/Y 0.01fF
C34373 INVX1_LOC_64/A NOR2X1_LOC_545/A 0.01fF
C34374 NOR2X1_LOC_817/Y NOR2X1_LOC_160/B 0.06fF
C34375 INVX1_LOC_91/A NOR2X1_LOC_435/A 0.03fF
C34376 NAND2X1_LOC_538/Y INVX1_LOC_31/A 0.09fF
C34377 NOR2X1_LOC_459/A INVX1_LOC_32/A 0.00fF
C34378 INVX1_LOC_25/A NOR2X1_LOC_773/a_36_216# 0.01fF
C34379 NOR2X1_LOC_833/Y NOR2X1_LOC_833/a_36_216# 0.00fF
C34380 INVX1_LOC_66/Y INVX1_LOC_46/A 0.01fF
C34381 NAND2X1_LOC_347/B INVX1_LOC_72/A 0.08fF
C34382 NOR2X1_LOC_405/A NOR2X1_LOC_743/Y 0.02fF
C34383 INVX1_LOC_7/A NOR2X1_LOC_297/A 0.01fF
C34384 INVX1_LOC_83/A INVX1_LOC_32/A 0.01fF
C34385 NOR2X1_LOC_567/B INVX1_LOC_29/A 0.16fF
C34386 NAND2X1_LOC_725/B NAND2X1_LOC_501/a_36_24# 0.01fF
C34387 INVX1_LOC_83/A NOR2X1_LOC_623/B 3.76fF
C34388 NAND2X1_LOC_123/Y NOR2X1_LOC_89/A 0.03fF
C34389 NOR2X1_LOC_772/B NOR2X1_LOC_772/Y 0.02fF
C34390 INVX1_LOC_77/Y NOR2X1_LOC_694/Y 0.04fF
C34391 NOR2X1_LOC_530/Y INVX1_LOC_31/A 2.05fF
C34392 INVX1_LOC_10/A NOR2X1_LOC_248/A 0.07fF
C34393 INVX1_LOC_36/A NOR2X1_LOC_592/A 0.07fF
C34394 NOR2X1_LOC_417/a_36_216# INVX1_LOC_178/A 0.02fF
C34395 NAND2X1_LOC_724/Y NOR2X1_LOC_773/Y 0.36fF
C34396 NOR2X1_LOC_598/B INVX1_LOC_149/A 0.01fF
C34397 NOR2X1_LOC_772/B NOR2X1_LOC_392/B 0.60fF
C34398 NAND2X1_LOC_51/B INVX1_LOC_12/A 0.01fF
C34399 INVX1_LOC_136/A NOR2X1_LOC_457/A 0.10fF
C34400 NAND2X1_LOC_67/Y INVX1_LOC_24/A 0.01fF
C34401 INVX1_LOC_20/A NOR2X1_LOC_695/a_36_216# 0.00fF
C34402 NOR2X1_LOC_528/Y NOR2X1_LOC_661/A 0.01fF
C34403 INVX1_LOC_45/A NAND2X1_LOC_352/B 0.72fF
C34404 NOR2X1_LOC_276/Y INVX1_LOC_30/A 0.00fF
C34405 INVX1_LOC_122/Y NOR2X1_LOC_502/Y 0.02fF
C34406 INVX1_LOC_91/A INVX1_LOC_63/A 5.59fF
C34407 INVX1_LOC_176/A NOR2X1_LOC_862/B 0.03fF
C34408 INVX1_LOC_13/Y NOR2X1_LOC_392/B 0.10fF
C34409 INVX1_LOC_311/A INVX1_LOC_12/A 0.66fF
C34410 NOR2X1_LOC_67/A NOR2X1_LOC_392/Y 0.03fF
C34411 INVX1_LOC_278/A INVX1_LOC_256/Y 0.10fF
C34412 INVX1_LOC_232/Y INVX1_LOC_35/A 0.03fF
C34413 NOR2X1_LOC_470/B INVX1_LOC_77/A 0.07fF
C34414 NAND2X1_LOC_858/B NOR2X1_LOC_46/a_36_216# 0.01fF
C34415 INVX1_LOC_16/A INVX1_LOC_29/Y 0.06fF
C34416 INVX1_LOC_222/Y NOR2X1_LOC_6/B -0.00fF
C34417 INVX1_LOC_59/A NAND2X1_LOC_139/A 0.01fF
C34418 NOR2X1_LOC_647/A NOR2X1_LOC_332/A 0.02fF
C34419 INVX1_LOC_11/A INVX1_LOC_314/Y 0.20fF
C34420 NAND2X1_LOC_799/A NOR2X1_LOC_152/Y 0.07fF
C34421 INVX1_LOC_249/A INVX1_LOC_256/A 0.03fF
C34422 INVX1_LOC_88/A NOR2X1_LOC_172/Y 0.28fF
C34423 NOR2X1_LOC_45/B NAND2X1_LOC_499/a_36_24# 0.01fF
C34424 NAND2X1_LOC_338/B NOR2X1_LOC_291/Y 0.09fF
C34425 INVX1_LOC_48/Y NOR2X1_LOC_124/B 0.03fF
C34426 NAND2X1_LOC_624/B INVX1_LOC_172/Y 0.00fF
C34427 NOR2X1_LOC_596/Y NOR2X1_LOC_596/A 0.01fF
C34428 INVX1_LOC_136/A INVX1_LOC_30/A 1.99fF
C34429 INVX1_LOC_6/Y INVX1_LOC_256/A 0.09fF
C34430 NAND2X1_LOC_9/Y INVX1_LOC_13/A 0.22fF
C34431 INVX1_LOC_269/A NOR2X1_LOC_142/Y 0.19fF
C34432 GATE_662 INVX1_LOC_53/A 0.03fF
C34433 INVX1_LOC_1/A NOR2X1_LOC_773/a_36_216# 0.01fF
C34434 D_INPUT_1 NAND2X1_LOC_656/Y 0.07fF
C34435 INVX1_LOC_17/A INVX1_LOC_34/A 0.03fF
C34436 NOR2X1_LOC_216/B NOR2X1_LOC_536/A 0.03fF
C34437 NOR2X1_LOC_15/Y NOR2X1_LOC_315/Y 0.03fF
C34438 NOR2X1_LOC_647/Y NOR2X1_LOC_554/B 0.23fF
C34439 INVX1_LOC_46/Y INVX1_LOC_230/A 0.03fF
C34440 NOR2X1_LOC_517/Y INVX1_LOC_217/A 0.05fF
C34441 INVX1_LOC_21/A INVX1_LOC_214/Y 0.03fF
C34442 NOR2X1_LOC_541/Y NOR2X1_LOC_344/A 0.67fF
C34443 INVX1_LOC_46/A NAND2X1_LOC_489/Y 0.01fF
C34444 INVX1_LOC_76/A NAND2X1_LOC_773/B 0.12fF
C34445 NOR2X1_LOC_106/A INVX1_LOC_23/A 0.05fF
C34446 INVX1_LOC_41/A NOR2X1_LOC_254/A 0.19fF
C34447 NOR2X1_LOC_620/Y NOR2X1_LOC_590/A 0.00fF
C34448 NOR2X1_LOC_197/B INVX1_LOC_9/A 0.19fF
C34449 NOR2X1_LOC_826/Y D_INPUT_0 0.01fF
C34450 NOR2X1_LOC_471/Y INVX1_LOC_34/A 0.10fF
C34451 NOR2X1_LOC_620/Y INVX1_LOC_22/Y 0.02fF
C34452 INVX1_LOC_117/A NOR2X1_LOC_814/A 0.33fF
C34453 NOR2X1_LOC_272/Y INVX1_LOC_53/Y 0.01fF
C34454 NOR2X1_LOC_91/A NAND2X1_LOC_863/A 0.07fF
C34455 NAND2X1_LOC_787/A NAND2X1_LOC_862/Y 0.20fF
C34456 NOR2X1_LOC_655/B INVX1_LOC_269/A 0.10fF
C34457 INVX1_LOC_229/A NAND2X1_LOC_733/B 0.28fF
C34458 INPUT_0 NOR2X1_LOC_301/A 0.10fF
C34459 INVX1_LOC_220/Y INVX1_LOC_50/Y 0.03fF
C34460 INVX1_LOC_136/Y INVX1_LOC_44/A 0.24fF
C34461 NAND2X1_LOC_640/a_36_24# INVX1_LOC_41/Y 0.00fF
C34462 NOR2X1_LOC_536/A NAND2X1_LOC_477/Y 0.03fF
C34463 INVX1_LOC_256/A INVX1_LOC_206/A 0.10fF
C34464 INVX1_LOC_17/A NAND2X1_LOC_231/Y 0.10fF
C34465 NOR2X1_LOC_806/Y INVX1_LOC_134/A 0.12fF
C34466 INVX1_LOC_18/A NOR2X1_LOC_152/Y 0.33fF
C34467 NOR2X1_LOC_453/Y D_GATE_222 -0.02fF
C34468 NOR2X1_LOC_589/A NAND2X1_LOC_474/Y 0.00fF
C34469 NOR2X1_LOC_852/A NAND2X1_LOC_361/Y 0.03fF
C34470 NOR2X1_LOC_216/B NAND2X1_LOC_93/B 0.10fF
C34471 INVX1_LOC_45/A NOR2X1_LOC_344/A 0.03fF
C34472 NAND2X1_LOC_728/Y NOR2X1_LOC_152/Y 0.11fF
C34473 INVX1_LOC_36/A NAND2X1_LOC_276/Y 0.00fF
C34474 INVX1_LOC_18/A INVX1_LOC_113/Y 0.14fF
C34475 INVX1_LOC_11/A NOR2X1_LOC_778/B 0.29fF
C34476 NOR2X1_LOC_568/A NOR2X1_LOC_344/A 0.02fF
C34477 NOR2X1_LOC_641/B NOR2X1_LOC_264/Y 0.00fF
C34478 NOR2X1_LOC_296/Y NOR2X1_LOC_78/B 0.19fF
C34479 NAND2X1_LOC_725/Y NOR2X1_LOC_409/Y 0.59fF
C34480 INVX1_LOC_33/A NOR2X1_LOC_354/B 0.02fF
C34481 VDD INVX1_LOC_290/Y 2.03fF
C34482 NOR2X1_LOC_591/Y INVX1_LOC_141/Y 0.03fF
C34483 INVX1_LOC_27/A NOR2X1_LOC_415/A 0.01fF
C34484 NOR2X1_LOC_773/Y NAND2X1_LOC_793/Y 0.07fF
C34485 NOR2X1_LOC_583/Y INVX1_LOC_77/Y 0.03fF
C34486 NOR2X1_LOC_506/a_36_216# INVX1_LOC_12/A 0.00fF
C34487 INVX1_LOC_21/A NAND2X1_LOC_808/A 0.00fF
C34488 INVX1_LOC_50/A NOR2X1_LOC_188/A 0.04fF
C34489 NOR2X1_LOC_772/B NOR2X1_LOC_389/B 0.08fF
C34490 INVX1_LOC_229/A NAND2X1_LOC_735/B 0.00fF
C34491 NOR2X1_LOC_208/Y NOR2X1_LOC_353/a_36_216# 0.00fF
C34492 NOR2X1_LOC_468/Y NOR2X1_LOC_383/Y 0.08fF
C34493 INVX1_LOC_50/A NOR2X1_LOC_548/B 1.36fF
C34494 NOR2X1_LOC_798/A NOR2X1_LOC_174/B 0.82fF
C34495 NOR2X1_LOC_405/A NAND2X1_LOC_72/B 0.03fF
C34496 NOR2X1_LOC_311/Y NAND2X1_LOC_175/Y 0.05fF
C34497 INVX1_LOC_13/Y INVX1_LOC_90/A 0.03fF
C34498 NOR2X1_LOC_817/Y NOR2X1_LOC_516/B 0.03fF
C34499 NOR2X1_LOC_609/A INVX1_LOC_155/Y 0.00fF
C34500 INVX1_LOC_45/Y INVX1_LOC_155/A 0.04fF
C34501 NOR2X1_LOC_360/Y INVX1_LOC_8/A 0.07fF
C34502 NOR2X1_LOC_88/Y NOR2X1_LOC_697/Y 0.00fF
C34503 NOR2X1_LOC_667/A NAND2X1_LOC_733/Y 0.03fF
C34504 INVX1_LOC_32/A INVX1_LOC_46/A 0.04fF
C34505 NOR2X1_LOC_216/B NOR2X1_LOC_649/B 0.00fF
C34506 INVX1_LOC_13/Y NOR2X1_LOC_389/B 1.40fF
C34507 NAND2X1_LOC_785/Y INVX1_LOC_217/A 0.06fF
C34508 INVX1_LOC_223/A INVX1_LOC_177/A 0.00fF
C34509 INVX1_LOC_39/A INPUT_1 2.88fF
C34510 NAND2X1_LOC_77/a_36_24# INVX1_LOC_89/A 0.00fF
C34511 NOR2X1_LOC_614/Y INVX1_LOC_292/A 0.00fF
C34512 NOR2X1_LOC_246/A NAND2X1_LOC_703/Y 0.18fF
C34513 NOR2X1_LOC_151/a_36_216# NOR2X1_LOC_678/A 0.00fF
C34514 NOR2X1_LOC_612/Y INVX1_LOC_19/A 0.03fF
C34515 NOR2X1_LOC_344/A INVX1_LOC_71/A 0.04fF
C34516 NAND2X1_LOC_53/Y NOR2X1_LOC_589/A 1.65fF
C34517 INVX1_LOC_136/A NAND2X1_LOC_722/A 0.98fF
C34518 INVX1_LOC_35/A NOR2X1_LOC_97/A 0.02fF
C34519 NOR2X1_LOC_489/B NOR2X1_LOC_74/A 0.02fF
C34520 NAND2X1_LOC_656/A NOR2X1_LOC_6/B 0.13fF
C34521 NAND2X1_LOC_30/Y INPUT_5 0.15fF
C34522 NAND2X1_LOC_315/a_36_24# NOR2X1_LOC_52/B 0.00fF
C34523 INVX1_LOC_35/A INVX1_LOC_193/Y 0.03fF
C34524 NOR2X1_LOC_124/A NAND2X1_LOC_99/A 0.02fF
C34525 NAND2X1_LOC_72/Y NOR2X1_LOC_188/A 0.21fF
C34526 NOR2X1_LOC_15/Y NAND2X1_LOC_624/A 0.01fF
C34527 INVX1_LOC_84/A NOR2X1_LOC_697/Y 0.04fF
C34528 NOR2X1_LOC_36/A INVX1_LOC_20/A 0.00fF
C34529 NOR2X1_LOC_67/A NOR2X1_LOC_86/Y 0.02fF
C34530 NAND2X1_LOC_455/B INVX1_LOC_118/A 0.20fF
C34531 NAND2X1_LOC_357/B INVX1_LOC_71/A 0.10fF
C34532 INVX1_LOC_24/A NAND2X1_LOC_629/Y 0.05fF
C34533 INVX1_LOC_124/A NOR2X1_LOC_191/B 0.01fF
C34534 NOR2X1_LOC_667/A INVX1_LOC_217/A 0.02fF
C34535 NOR2X1_LOC_720/B NOR2X1_LOC_419/Y 0.00fF
C34536 INVX1_LOC_314/Y NOR2X1_LOC_52/B 0.03fF
C34537 D_INPUT_6 INVX1_LOC_140/A 0.14fF
C34538 NAND2X1_LOC_361/Y NOR2X1_LOC_285/B 0.01fF
C34539 NOR2X1_LOC_179/Y INVX1_LOC_63/A 0.06fF
C34540 INVX1_LOC_90/A INVX1_LOC_88/A 0.04fF
C34541 NAND2X1_LOC_175/Y INVX1_LOC_46/A 0.23fF
C34542 NOR2X1_LOC_286/Y INVX1_LOC_89/A 0.01fF
C34543 NOR2X1_LOC_373/Y NAND2X1_LOC_550/A 0.04fF
C34544 NAND2X1_LOC_384/a_36_24# NOR2X1_LOC_160/B 0.00fF
C34545 NAND2X1_LOC_741/B NAND2X1_LOC_863/B 0.03fF
C34546 NOR2X1_LOC_15/Y NOR2X1_LOC_166/Y 0.01fF
C34547 NOR2X1_LOC_527/Y NOR2X1_LOC_406/A 0.01fF
C34548 NOR2X1_LOC_389/B INVX1_LOC_88/A 0.03fF
C34549 INPUT_3 INVX1_LOC_83/A 0.00fF
C34550 NOR2X1_LOC_841/A INVX1_LOC_272/A 0.10fF
C34551 NOR2X1_LOC_208/Y NOR2X1_LOC_352/Y 0.02fF
C34552 NOR2X1_LOC_389/A NOR2X1_LOC_366/Y 0.28fF
C34553 INVX1_LOC_93/A INVX1_LOC_126/Y 0.12fF
C34554 INVX1_LOC_18/A NAND2X1_LOC_859/B 0.02fF
C34555 NAND2X1_LOC_364/A INVX1_LOC_53/Y 0.07fF
C34556 NAND2X1_LOC_796/B NAND2X1_LOC_858/B 0.25fF
C34557 INVX1_LOC_263/A NOR2X1_LOC_457/B 0.02fF
C34558 INVX1_LOC_269/A NOR2X1_LOC_381/a_36_216# 0.01fF
C34559 INVX1_LOC_223/Y NOR2X1_LOC_551/Y 0.01fF
C34560 NOR2X1_LOC_237/Y NAND2X1_LOC_374/Y 0.02fF
C34561 NOR2X1_LOC_815/Y INVX1_LOC_2/A 0.14fF
C34562 NAND2X1_LOC_82/a_36_24# NOR2X1_LOC_649/B 0.00fF
C34563 NAND2X1_LOC_733/Y NAND2X1_LOC_804/a_36_24# 0.06fF
C34564 NAND2X1_LOC_218/B NAND2X1_LOC_671/a_36_24# 0.00fF
C34565 NAND2X1_LOC_116/A NOR2X1_LOC_844/A 0.03fF
C34566 INVX1_LOC_85/A INVX1_LOC_121/Y 0.00fF
C34567 INVX1_LOC_294/Y NOR2X1_LOC_612/B 0.01fF
C34568 NOR2X1_LOC_667/A NAND2X1_LOC_787/B 0.00fF
C34569 NOR2X1_LOC_617/Y INVX1_LOC_172/Y 0.02fF
C34570 INVX1_LOC_24/A NOR2X1_LOC_719/A 0.00fF
C34571 NOR2X1_LOC_124/B NOR2X1_LOC_84/Y 0.01fF
C34572 NAND2X1_LOC_785/Y INVX1_LOC_304/Y -0.01fF
C34573 INVX1_LOC_14/A NOR2X1_LOC_74/A 0.16fF
C34574 INVX1_LOC_30/Y NAND2X1_LOC_656/A 0.02fF
C34575 NOR2X1_LOC_647/B NOR2X1_LOC_19/B 0.02fF
C34576 NOR2X1_LOC_220/A NOR2X1_LOC_562/a_36_216# 0.13fF
C34577 INVX1_LOC_30/A NAND2X1_LOC_862/Y 0.05fF
C34578 NOR2X1_LOC_332/A INVX1_LOC_205/A 0.01fF
C34579 INVX1_LOC_81/A INVX1_LOC_290/A 0.04fF
C34580 INVX1_LOC_24/A NOR2X1_LOC_561/Y 0.07fF
C34581 INVX1_LOC_17/A INPUT_0 0.91fF
C34582 INVX1_LOC_14/A NOR2X1_LOC_9/Y 0.23fF
C34583 INVX1_LOC_90/A NOR2X1_LOC_500/B 0.13fF
C34584 INVX1_LOC_24/A INVX1_LOC_7/A 0.04fF
C34585 NAND2X1_LOC_85/Y INVX1_LOC_15/A 0.10fF
C34586 INVX1_LOC_18/A NAND2X1_LOC_861/Y 0.07fF
C34587 INVX1_LOC_142/A INVX1_LOC_85/Y 0.01fF
C34588 INVX1_LOC_35/A NAND2X1_LOC_287/B 0.07fF
C34589 INVX1_LOC_255/Y NOR2X1_LOC_649/a_36_216# 0.01fF
C34590 INVX1_LOC_304/Y NOR2X1_LOC_667/A 0.00fF
C34591 NOR2X1_LOC_420/Y NAND2X1_LOC_447/Y 0.11fF
C34592 NOR2X1_LOC_464/B INVX1_LOC_96/A 0.01fF
C34593 NOR2X1_LOC_401/A INVX1_LOC_286/A 0.02fF
C34594 NOR2X1_LOC_287/A NOR2X1_LOC_288/A 0.00fF
C34595 NOR2X1_LOC_252/Y INVX1_LOC_34/A 0.02fF
C34596 NAND2X1_LOC_773/Y NOR2X1_LOC_78/A 0.01fF
C34597 NOR2X1_LOC_648/a_36_216# NOR2X1_LOC_655/B 0.02fF
C34598 INVX1_LOC_61/A INPUT_1 0.19fF
C34599 INVX1_LOC_254/A D_INPUT_0 0.03fF
C34600 NOR2X1_LOC_448/Y NOR2X1_LOC_448/A 0.07fF
C34601 NAND2X1_LOC_555/Y INPUT_0 0.09fF
C34602 NOR2X1_LOC_644/A NOR2X1_LOC_598/a_36_216# 0.00fF
C34603 INVX1_LOC_224/A NOR2X1_LOC_557/A 0.32fF
C34604 NOR2X1_LOC_561/Y NOR2X1_LOC_557/Y 0.26fF
C34605 INVX1_LOC_96/Y INVX1_LOC_52/A 0.03fF
C34606 INVX1_LOC_214/A INVX1_LOC_214/Y 0.01fF
C34607 INVX1_LOC_103/A NOR2X1_LOC_45/B 0.14fF
C34608 INVX1_LOC_274/A NOR2X1_LOC_383/B 0.01fF
C34609 NOR2X1_LOC_186/Y NOR2X1_LOC_305/Y 0.13fF
C34610 NOR2X1_LOC_65/B NAND2X1_LOC_488/a_36_24# 0.01fF
C34611 INVX1_LOC_172/A NAND2X1_LOC_861/Y 0.91fF
C34612 NOR2X1_LOC_160/B INVX1_LOC_286/A 0.11fF
C34613 INVX1_LOC_303/A INVX1_LOC_90/A 0.09fF
C34614 NOR2X1_LOC_643/Y INVX1_LOC_20/Y 0.03fF
C34615 INVX1_LOC_17/A NAND2X1_LOC_649/B 0.01fF
C34616 INVX1_LOC_132/A INVX1_LOC_47/A 0.00fF
C34617 NOR2X1_LOC_690/A D_INPUT_0 0.02fF
C34618 NOR2X1_LOC_67/A INVX1_LOC_25/Y 1.25fF
C34619 NAND2X1_LOC_190/Y NAND2X1_LOC_447/Y 0.20fF
C34620 INVX1_LOC_9/Y NOR2X1_LOC_78/B 0.02fF
C34621 NAND2X1_LOC_573/Y NOR2X1_LOC_305/Y 0.01fF
C34622 NOR2X1_LOC_226/A NAND2X1_LOC_182/a_36_24# 0.01fF
C34623 INVX1_LOC_90/A NOR2X1_LOC_672/Y 0.12fF
C34624 NAND2X1_LOC_569/A NOR2X1_LOC_71/Y 0.05fF
C34625 NOR2X1_LOC_615/Y NAND2X1_LOC_623/B 0.09fF
C34626 NOR2X1_LOC_413/Y D_INPUT_0 0.01fF
C34627 INVX1_LOC_223/A INVX1_LOC_285/Y 0.01fF
C34628 NOR2X1_LOC_454/Y VDD 2.80fF
C34629 INVX1_LOC_227/Y NOR2X1_LOC_74/A 0.01fF
C34630 INVX1_LOC_200/A INVX1_LOC_304/A 0.06fF
C34631 INVX1_LOC_58/A NOR2X1_LOC_364/A 0.07fF
C34632 INVX1_LOC_33/A NOR2X1_LOC_552/a_36_216# 0.00fF
C34633 NOR2X1_LOC_644/Y INVX1_LOC_279/A 0.08fF
C34634 NAND2X1_LOC_364/A NOR2X1_LOC_113/B 0.02fF
C34635 NOR2X1_LOC_773/Y INVX1_LOC_300/A 0.14fF
C34636 NOR2X1_LOC_223/a_36_216# D_GATE_222 0.02fF
C34637 INVX1_LOC_93/A NOR2X1_LOC_536/A 0.07fF
C34638 NAND2X1_LOC_702/a_36_24# NOR2X1_LOC_331/B 0.01fF
C34639 INVX1_LOC_128/A INVX1_LOC_272/A 0.03fF
C34640 NAND2X1_LOC_724/A NOR2X1_LOC_305/Y 0.00fF
C34641 INVX1_LOC_272/Y INVX1_LOC_20/A 0.12fF
C34642 NOR2X1_LOC_168/Y NOR2X1_LOC_337/A 0.01fF
C34643 NOR2X1_LOC_381/Y NOR2X1_LOC_42/a_36_216# 0.00fF
C34644 NOR2X1_LOC_135/Y NOR2X1_LOC_577/Y 0.03fF
C34645 INVX1_LOC_49/Y INVX1_LOC_94/Y 2.29fF
C34646 NAND2X1_LOC_563/Y INVX1_LOC_89/A 0.07fF
C34647 INVX1_LOC_38/Y INVX1_LOC_9/A 0.06fF
C34648 NAND2X1_LOC_68/a_36_24# INVX1_LOC_281/A 0.03fF
C34649 INVX1_LOC_255/Y INVX1_LOC_316/Y 0.03fF
C34650 NAND2X1_LOC_84/Y NOR2X1_LOC_74/A 0.08fF
C34651 NOR2X1_LOC_180/B INVX1_LOC_104/A 0.08fF
C34652 NOR2X1_LOC_186/Y NAND2X1_LOC_600/a_36_24# 0.00fF
C34653 INVX1_LOC_24/A NOR2X1_LOC_167/Y 0.03fF
C34654 INVX1_LOC_62/A NOR2X1_LOC_87/Y -0.01fF
C34655 INVX1_LOC_8/Y NOR2X1_LOC_751/A 0.02fF
C34656 NOR2X1_LOC_632/Y INVX1_LOC_22/A 0.03fF
C34657 NOR2X1_LOC_667/A NAND2X1_LOC_808/A 0.27fF
C34658 INVX1_LOC_58/A INVX1_LOC_285/A 0.33fF
C34659 INVX1_LOC_248/A NAND2X1_LOC_808/A 0.00fF
C34660 NAND2X1_LOC_84/Y NOR2X1_LOC_9/Y 0.00fF
C34661 NAND2X1_LOC_15/a_36_24# NAND2X1_LOC_96/A 0.00fF
C34662 INVX1_LOC_10/A NOR2X1_LOC_131/Y 0.03fF
C34663 NOR2X1_LOC_598/B NOR2X1_LOC_800/a_36_216# 0.15fF
C34664 INVX1_LOC_58/A NOR2X1_LOC_814/A 0.07fF
C34665 NAND2X1_LOC_564/B NAND2X1_LOC_392/Y 0.04fF
C34666 INVX1_LOC_26/A INVX1_LOC_29/A 0.02fF
C34667 NOR2X1_LOC_15/Y NAND2X1_LOC_93/a_36_24# 0.00fF
C34668 NAND2X1_LOC_573/Y NAND2X1_LOC_600/a_36_24# 0.00fF
C34669 NAND2X1_LOC_112/Y INVX1_LOC_279/A 0.00fF
C34670 INVX1_LOC_103/A INVX1_LOC_281/A 0.10fF
C34671 INVX1_LOC_111/Y NOR2X1_LOC_356/A 0.03fF
C34672 NAND2X1_LOC_462/B NAND2X1_LOC_735/B 0.00fF
C34673 INVX1_LOC_223/A NOR2X1_LOC_137/B 0.01fF
C34674 INVX1_LOC_73/A INVX1_LOC_104/A 0.07fF
C34675 NOR2X1_LOC_264/Y NOR2X1_LOC_751/A 0.01fF
C34676 NAND2X1_LOC_725/Y INVX1_LOC_240/Y 0.12fF
C34677 NOR2X1_LOC_589/A INVX1_LOC_10/A 0.06fF
C34678 INVX1_LOC_88/A INVX1_LOC_38/A 0.06fF
C34679 NOR2X1_LOC_355/A INVX1_LOC_16/A 0.07fF
C34680 NAND2X1_LOC_364/A NOR2X1_LOC_557/a_36_216# 0.00fF
C34681 NOR2X1_LOC_647/A NOR2X1_LOC_847/A 0.35fF
C34682 INVX1_LOC_21/A INVX1_LOC_92/A 0.61fF
C34683 INVX1_LOC_299/A NAND2X1_LOC_204/a_36_24# 0.00fF
C34684 NAND2X1_LOC_198/B NOR2X1_LOC_405/A 0.36fF
C34685 NOR2X1_LOC_644/Y INVX1_LOC_182/Y 0.01fF
C34686 NAND2X1_LOC_331/a_36_24# NAND2X1_LOC_349/B 0.06fF
C34687 INVX1_LOC_83/A GATE_662 0.07fF
C34688 INVX1_LOC_178/A NAND2X1_LOC_798/B 0.03fF
C34689 INVX1_LOC_217/A NOR2X1_LOC_670/Y 0.18fF
C34690 NOR2X1_LOC_569/A INVX1_LOC_104/A 0.03fF
C34691 NOR2X1_LOC_590/A INVX1_LOC_117/A 0.19fF
C34692 NOR2X1_LOC_612/B NOR2X1_LOC_74/A 0.08fF
C34693 NOR2X1_LOC_561/Y NOR2X1_LOC_130/A 0.04fF
C34694 INVX1_LOC_22/Y INVX1_LOC_117/A 0.03fF
C34695 INVX1_LOC_24/A NOR2X1_LOC_824/Y 0.05fF
C34696 NOR2X1_LOC_67/A INVX1_LOC_75/A 0.07fF
C34697 NAND2X1_LOC_337/a_36_24# NOR2X1_LOC_536/A 0.00fF
C34698 INVX1_LOC_111/Y NOR2X1_LOC_74/A 0.00fF
C34699 NAND2X1_LOC_725/B INVX1_LOC_241/Y 0.02fF
C34700 INVX1_LOC_49/A NOR2X1_LOC_448/A 0.01fF
C34701 NOR2X1_LOC_97/a_36_216# NOR2X1_LOC_99/B 0.04fF
C34702 INVX1_LOC_33/A NOR2X1_LOC_139/Y 0.06fF
C34703 INVX1_LOC_24/A INVX1_LOC_76/A 2.28fF
C34704 INVX1_LOC_206/A INVX1_LOC_69/Y 0.90fF
C34705 INVX1_LOC_6/A NOR2X1_LOC_709/A 0.17fF
C34706 NOR2X1_LOC_135/Y INVX1_LOC_22/A 0.00fF
C34707 NAND2X1_LOC_722/A NOR2X1_LOC_165/a_36_216# 0.03fF
C34708 INVX1_LOC_132/A INVX1_LOC_95/Y 0.10fF
C34709 NOR2X1_LOC_632/Y NOR2X1_LOC_735/Y 0.15fF
C34710 INVX1_LOC_311/A NAND2X1_LOC_832/a_36_24# 0.00fF
C34711 NOR2X1_LOC_160/B INVX1_LOC_54/A 0.03fF
C34712 NAND2X1_LOC_799/A NAND2X1_LOC_802/Y 0.05fF
C34713 NOR2X1_LOC_45/B INVX1_LOC_240/A 0.03fF
C34714 NOR2X1_LOC_106/A INVX1_LOC_313/A 0.01fF
C34715 INVX1_LOC_89/A INVX1_LOC_148/Y 0.01fF
C34716 INVX1_LOC_190/A INVX1_LOC_190/Y 0.09fF
C34717 NAND2X1_LOC_670/a_36_24# NOR2X1_LOC_536/A 0.00fF
C34718 INVX1_LOC_33/A NAND2X1_LOC_468/B 0.03fF
C34719 NOR2X1_LOC_91/A NAND2X1_LOC_444/B 0.01fF
C34720 NOR2X1_LOC_38/B INVX1_LOC_112/Y 0.02fF
C34721 NOR2X1_LOC_744/Y NOR2X1_LOC_111/A 0.03fF
C34722 NOR2X1_LOC_814/Y NOR2X1_LOC_846/B 0.05fF
C34723 INVX1_LOC_2/A NOR2X1_LOC_7/Y 0.11fF
C34724 INVX1_LOC_180/A NAND2X1_LOC_453/A 0.01fF
C34725 NOR2X1_LOC_827/a_36_216# NOR2X1_LOC_78/A 0.00fF
C34726 INVX1_LOC_77/A VDD 3.64fF
C34727 NOR2X1_LOC_415/A NOR2X1_LOC_19/B 0.06fF
C34728 NOR2X1_LOC_355/A INVX1_LOC_28/A 0.09fF
C34729 INVX1_LOC_225/A INVX1_LOC_95/Y 0.01fF
C34730 NOR2X1_LOC_428/Y INVX1_LOC_92/A 0.12fF
C34731 INVX1_LOC_254/Y INVX1_LOC_37/A 0.04fF
C34732 INVX1_LOC_292/A NOR2X1_LOC_862/B 0.34fF
C34733 INVX1_LOC_284/A NOR2X1_LOC_293/a_36_216# 0.01fF
C34734 NAND2X1_LOC_372/a_36_24# INVX1_LOC_206/Y 0.01fF
C34735 NAND2X1_LOC_9/Y INVX1_LOC_32/A 0.06fF
C34736 INVX1_LOC_49/A INVX1_LOC_14/Y 0.05fF
C34737 INVX1_LOC_15/A NOR2X1_LOC_247/Y 0.21fF
C34738 NOR2X1_LOC_391/Y NOR2X1_LOC_121/A -0.00fF
C34739 INVX1_LOC_233/A INVX1_LOC_32/A 0.10fF
C34740 NAND2X1_LOC_195/Y INVX1_LOC_54/A 0.00fF
C34741 NOR2X1_LOC_334/Y INVX1_LOC_23/A 0.25fF
C34742 NOR2X1_LOC_186/Y NAND2X1_LOC_806/a_36_24# 0.00fF
C34743 INVX1_LOC_27/A NOR2X1_LOC_89/A 0.10fF
C34744 INVX1_LOC_1/Y NOR2X1_LOC_114/A 0.01fF
C34745 INVX1_LOC_38/Y NOR2X1_LOC_861/Y 0.01fF
C34746 INVX1_LOC_2/A NAND2X1_LOC_212/Y 0.00fF
C34747 INVX1_LOC_18/A INVX1_LOC_291/A 0.07fF
C34748 NOR2X1_LOC_565/A NOR2X1_LOC_197/B 0.28fF
C34749 INVX1_LOC_303/A INVX1_LOC_38/A 0.07fF
C34750 INVX1_LOC_1/Y INVX1_LOC_91/A 0.27fF
C34751 NAND2X1_LOC_354/Y INVX1_LOC_92/A 0.03fF
C34752 INVX1_LOC_57/A NOR2X1_LOC_693/Y 0.07fF
C34753 NOR2X1_LOC_27/Y VDD 0.12fF
C34754 NAND2X1_LOC_303/B INVX1_LOC_140/Y 0.12fF
C34755 INVX1_LOC_124/A VDD 1.64fF
C34756 INVX1_LOC_57/A NAND2X1_LOC_288/B 0.00fF
C34757 NOR2X1_LOC_582/Y INVX1_LOC_92/A 1.01fF
C34758 NOR2X1_LOC_405/A INVX1_LOC_53/Y 0.07fF
C34759 NOR2X1_LOC_798/A INVX1_LOC_32/A 0.03fF
C34760 NOR2X1_LOC_690/A NAND2X1_LOC_848/A 0.08fF
C34761 NAND2X1_LOC_129/a_36_24# NOR2X1_LOC_84/Y 0.01fF
C34762 NOR2X1_LOC_798/A NOR2X1_LOC_623/B 0.03fF
C34763 INVX1_LOC_2/A INVX1_LOC_14/Y 0.12fF
C34764 INVX1_LOC_279/A NOR2X1_LOC_78/A 0.22fF
C34765 NOR2X1_LOC_815/Y INVX1_LOC_118/A 0.03fF
C34766 INVX1_LOC_298/A INVX1_LOC_78/A 0.02fF
C34767 INVX1_LOC_50/A NAND2X1_LOC_784/A 0.13fF
C34768 NAND2X1_LOC_474/Y INVX1_LOC_4/A -0.02fF
C34769 NOR2X1_LOC_80/Y NOR2X1_LOC_81/Y 0.11fF
C34770 NAND2X1_LOC_564/B NOR2X1_LOC_368/Y 0.03fF
C34771 NAND2X1_LOC_672/a_36_24# NOR2X1_LOC_673/A 0.02fF
C34772 NOR2X1_LOC_226/A INVX1_LOC_14/Y 0.00fF
C34773 INVX1_LOC_226/Y INVX1_LOC_20/A 0.07fF
C34774 NOR2X1_LOC_730/B INVX1_LOC_196/Y 0.03fF
C34775 NOR2X1_LOC_840/Y NOR2X1_LOC_678/A -0.01fF
C34776 NAND2X1_LOC_140/A NOR2X1_LOC_269/Y 0.03fF
C34777 NOR2X1_LOC_558/A INVX1_LOC_25/Y 0.46fF
C34778 INVX1_LOC_235/Y INVX1_LOC_253/A 0.04fF
C34779 INVX1_LOC_9/Y INVX1_LOC_46/A 0.04fF
C34780 INVX1_LOC_54/Y NOR2X1_LOC_536/A 1.12fF
C34781 NOR2X1_LOC_672/Y NAND2X1_LOC_848/Y 0.11fF
C34782 NAND2X1_LOC_39/Y INVX1_LOC_22/A 0.14fF
C34783 INVX1_LOC_235/Y INVX1_LOC_90/Y 0.02fF
C34784 D_INPUT_1 NOR2X1_LOC_717/A 0.02fF
C34785 NAND2X1_LOC_564/B INVX1_LOC_46/A 0.07fF
C34786 INVX1_LOC_269/A NOR2X1_LOC_28/a_36_216# 0.01fF
C34787 NOR2X1_LOC_687/Y VDD 0.69fF
C34788 NOR2X1_LOC_507/B NOR2X1_LOC_349/A -0.00fF
C34789 NAND2X1_LOC_840/Y NAND2X1_LOC_858/B 0.09fF
C34790 NAND2X1_LOC_390/A NAND2X1_LOC_650/B 0.37fF
C34791 INVX1_LOC_215/A NAND2X1_LOC_211/Y 0.23fF
C34792 INVX1_LOC_226/A NAND2X1_LOC_96/A 0.03fF
C34793 NOR2X1_LOC_399/Y INVX1_LOC_166/Y 0.09fF
C34794 INVX1_LOC_190/A NOR2X1_LOC_56/Y 0.03fF
C34795 NOR2X1_LOC_321/Y INVX1_LOC_78/A 0.19fF
C34796 NOR2X1_LOC_392/B NOR2X1_LOC_99/Y 0.82fF
C34797 INVX1_LOC_10/A INVX1_LOC_20/A 0.04fF
C34798 NOR2X1_LOC_180/B NOR2X1_LOC_600/Y 0.01fF
C34799 NAND2X1_LOC_703/Y NAND2X1_LOC_175/Y 0.02fF
C34800 NAND2X1_LOC_783/A INVX1_LOC_76/A 0.10fF
C34801 NOR2X1_LOC_383/B INVX1_LOC_306/Y 0.02fF
C34802 NOR2X1_LOC_709/A NOR2X1_LOC_79/A 0.10fF
C34803 VDD NAND2X1_LOC_796/Y 0.00fF
C34804 INVX1_LOC_290/A NOR2X1_LOC_363/Y 0.01fF
C34805 NOR2X1_LOC_654/A NOR2X1_LOC_406/A 0.14fF
C34806 NOR2X1_LOC_130/A INVX1_LOC_76/A 0.07fF
C34807 INVX1_LOC_16/A NOR2X1_LOC_694/Y 0.20fF
C34808 INVX1_LOC_298/Y NOR2X1_LOC_666/A 0.02fF
C34809 NOR2X1_LOC_742/A INVX1_LOC_91/A 0.07fF
C34810 INVX1_LOC_89/A INVX1_LOC_115/A 0.01fF
C34811 INVX1_LOC_54/Y NAND2X1_LOC_93/B 0.03fF
C34812 D_INPUT_1 NOR2X1_LOC_649/Y 0.09fF
C34813 INVX1_LOC_190/A VDD 0.12fF
C34814 INPUT_5 NOR2X1_LOC_694/a_36_216# 0.00fF
C34815 NOR2X1_LOC_15/Y NAND2X1_LOC_99/A 0.22fF
C34816 NOR2X1_LOC_84/A NOR2X1_LOC_649/B 0.01fF
C34817 INVX1_LOC_208/A INVX1_LOC_54/A 0.07fF
C34818 INVX1_LOC_214/A INVX1_LOC_92/A 0.18fF
C34819 NAND2X1_LOC_118/a_36_24# NOR2X1_LOC_862/B 0.06fF
C34820 NOR2X1_LOC_667/A INVX1_LOC_92/A 0.07fF
C34821 NOR2X1_LOC_763/Y INVX1_LOC_117/A 0.00fF
C34822 NOR2X1_LOC_778/B NOR2X1_LOC_858/a_36_216# 0.00fF
C34823 NOR2X1_LOC_717/A NOR2X1_LOC_652/Y 0.27fF
C34824 NAND2X1_LOC_276/Y INVX1_LOC_63/A 0.18fF
C34825 D_INPUT_3 INPUT_1 0.49fF
C34826 INVX1_LOC_248/A INVX1_LOC_92/A 0.29fF
C34827 INVX1_LOC_35/A INVX1_LOC_50/Y 0.04fF
C34828 INVX1_LOC_21/A INVX1_LOC_53/A 0.17fF
C34829 INVX1_LOC_73/A NAND2X1_LOC_674/a_36_24# 0.01fF
C34830 INVX1_LOC_17/A INVX1_LOC_183/A 0.02fF
C34831 INVX1_LOC_249/A NOR2X1_LOC_89/A 0.03fF
C34832 NOR2X1_LOC_113/B NOR2X1_LOC_405/A 0.05fF
C34833 INVX1_LOC_121/A INVX1_LOC_193/A 0.02fF
C34834 NOR2X1_LOC_172/Y INVX1_LOC_272/A 0.01fF
C34835 INVX1_LOC_28/A NOR2X1_LOC_111/A 0.07fF
C34836 INVX1_LOC_241/A INVX1_LOC_241/Y 0.01fF
C34837 INVX1_LOC_153/A INVX1_LOC_12/A 0.01fF
C34838 NAND2X1_LOC_341/A NOR2X1_LOC_155/A 0.03fF
C34839 NOR2X1_LOC_624/A NAND2X1_LOC_63/Y 0.02fF
C34840 INVX1_LOC_314/Y NOR2X1_LOC_159/a_36_216# 0.01fF
C34841 INVX1_LOC_41/A INVX1_LOC_106/A 0.03fF
C34842 NOR2X1_LOC_599/A NOR2X1_LOC_409/B 0.75fF
C34843 INVX1_LOC_11/A INVX1_LOC_271/A 0.03fF
C34844 NOR2X1_LOC_318/B INVX1_LOC_91/A 0.03fF
C34845 NAND2X1_LOC_842/B INVX1_LOC_66/Y 0.04fF
C34846 NOR2X1_LOC_703/A INVX1_LOC_117/A 0.01fF
C34847 NOR2X1_LOC_500/B INVX1_LOC_18/Y 0.20fF
C34848 INVX1_LOC_72/A NOR2X1_LOC_158/Y 1.42fF
C34849 INVX1_LOC_58/A NAND2X1_LOC_803/B 0.02fF
C34850 INVX1_LOC_93/Y INVX1_LOC_91/A 2.45fF
C34851 NOR2X1_LOC_160/B NAND2X1_LOC_215/A 0.03fF
C34852 NAND2X1_LOC_832/Y VDD 0.20fF
C34853 INVX1_LOC_153/Y INVX1_LOC_290/Y 0.02fF
C34854 INVX1_LOC_289/A INVX1_LOC_84/A 0.01fF
C34855 NOR2X1_LOC_261/a_36_216# INVX1_LOC_245/Y 0.00fF
C34856 NAND2X1_LOC_9/Y NOR2X1_LOC_296/Y 0.01fF
C34857 INVX1_LOC_40/A NOR2X1_LOC_820/B 0.01fF
C34858 NOR2X1_LOC_690/A NOR2X1_LOC_754/A -0.01fF
C34859 INVX1_LOC_272/Y INVX1_LOC_64/A 0.07fF
C34860 INVX1_LOC_58/A NOR2X1_LOC_590/A 0.03fF
C34861 INVX1_LOC_206/A NOR2X1_LOC_89/A 0.07fF
C34862 INVX1_LOC_45/A NOR2X1_LOC_443/Y 0.02fF
C34863 NOR2X1_LOC_647/A NOR2X1_LOC_554/B 0.05fF
C34864 INVX1_LOC_33/A NOR2X1_LOC_685/Y 0.03fF
C34865 NOR2X1_LOC_769/a_36_216# NOR2X1_LOC_48/Y 0.00fF
C34866 NAND2X1_LOC_214/B NAND2X1_LOC_222/B 0.01fF
C34867 INVX1_LOC_90/A NOR2X1_LOC_99/Y 0.00fF
C34868 NAND2X1_LOC_9/Y INPUT_3 0.36fF
C34869 INVX1_LOC_95/Y NAND2X1_LOC_642/Y 0.27fF
C34870 INVX1_LOC_120/A NOR2X1_LOC_862/B 0.00fF
C34871 NAND2X1_LOC_789/a_36_24# INVX1_LOC_26/Y 0.00fF
C34872 INVX1_LOC_255/Y NOR2X1_LOC_662/A 0.09fF
C34873 INVX1_LOC_177/A INVX1_LOC_290/Y 0.05fF
C34874 NAND2X1_LOC_214/B INVX1_LOC_11/A 0.07fF
C34875 INVX1_LOC_303/A NAND2X1_LOC_223/A 0.03fF
C34876 NAND2X1_LOC_866/A NAND2X1_LOC_175/Y 0.12fF
C34877 NAND2X1_LOC_149/Y NAND2X1_LOC_213/A 0.03fF
C34878 INVX1_LOC_196/Y NOR2X1_LOC_155/A 0.00fF
C34879 NAND2X1_LOC_222/B INVX1_LOC_27/A 0.04fF
C34880 NOR2X1_LOC_632/Y INVX1_LOC_186/Y 0.02fF
C34881 NAND2X1_LOC_200/B NOR2X1_LOC_89/A 0.22fF
C34882 NAND2X1_LOC_125/a_36_24# NOR2X1_LOC_649/B 0.00fF
C34883 NOR2X1_LOC_131/Y INVX1_LOC_12/A 0.03fF
C34884 NOR2X1_LOC_721/Y INVX1_LOC_9/A 0.02fF
C34885 NOR2X1_LOC_502/Y INVX1_LOC_50/Y 0.00fF
C34886 NAND2X1_LOC_562/Y NAND2X1_LOC_618/Y 0.27fF
C34887 INVX1_LOC_34/A INVX1_LOC_94/Y 0.03fF
C34888 INVX1_LOC_11/A INVX1_LOC_27/A 0.47fF
C34889 NOR2X1_LOC_464/B NOR2X1_LOC_15/Y 0.01fF
C34890 INVX1_LOC_149/Y INVX1_LOC_4/Y 0.02fF
C34891 INVX1_LOC_25/A NOR2X1_LOC_791/B 0.08fF
C34892 NAND2X1_LOC_862/A INVX1_LOC_102/A 0.01fF
C34893 NOR2X1_LOC_382/Y NOR2X1_LOC_660/Y 0.01fF
C34894 NOR2X1_LOC_219/Y INVX1_LOC_109/Y 0.02fF
C34895 NAND2X1_LOC_354/Y INVX1_LOC_53/A 0.05fF
C34896 NOR2X1_LOC_808/A INVX1_LOC_15/A 0.03fF
C34897 NOR2X1_LOC_71/Y NOR2X1_LOC_662/A 0.01fF
C34898 NOR2X1_LOC_91/A INVX1_LOC_209/Y 0.01fF
C34899 INVX1_LOC_45/A INVX1_LOC_213/A 0.08fF
C34900 NOR2X1_LOC_589/A INVX1_LOC_12/A 3.39fF
C34901 NAND2X1_LOC_51/B INVX1_LOC_92/A 0.06fF
C34902 NOR2X1_LOC_816/Y NAND2X1_LOC_655/A 0.04fF
C34903 NAND2X1_LOC_347/B NOR2X1_LOC_103/Y 0.01fF
C34904 NAND2X1_LOC_348/A NOR2X1_LOC_861/a_36_216# 0.00fF
C34905 INVX1_LOC_37/A NOR2X1_LOC_683/a_36_216# 0.00fF
C34906 NOR2X1_LOC_337/Y INVX1_LOC_9/A 0.01fF
C34907 NOR2X1_LOC_709/A NOR2X1_LOC_80/Y 0.68fF
C34908 INVX1_LOC_8/A INVX1_LOC_26/A 0.76fF
C34909 NOR2X1_LOC_653/B NOR2X1_LOC_441/Y 0.01fF
C34910 NOR2X1_LOC_164/Y NAND2X1_LOC_804/Y 0.05fF
C34911 NOR2X1_LOC_433/A INVX1_LOC_271/A 0.21fF
C34912 INVX1_LOC_311/A INVX1_LOC_92/A 0.46fF
C34913 NOR2X1_LOC_269/Y INVX1_LOC_118/Y 0.27fF
C34914 NAND2X1_LOC_595/a_36_24# NAND2X1_LOC_20/B 0.00fF
C34915 INVX1_LOC_200/Y NOR2X1_LOC_716/B 0.00fF
C34916 NAND2X1_LOC_231/Y INVX1_LOC_94/Y 0.01fF
C34917 INVX1_LOC_232/A INVX1_LOC_251/A 0.01fF
C34918 INVX1_LOC_34/A INVX1_LOC_296/A 0.03fF
C34919 NOR2X1_LOC_500/Y INVX1_LOC_4/A 0.07fF
C34920 INVX1_LOC_226/Y INVX1_LOC_4/A 0.07fF
C34921 INVX1_LOC_294/Y NOR2X1_LOC_383/B 0.03fF
C34922 INVX1_LOC_24/Y NAND2X1_LOC_171/a_36_24# 0.07fF
C34923 INVX1_LOC_90/A INVX1_LOC_272/A 0.07fF
C34924 INVX1_LOC_171/A INVX1_LOC_12/A 0.07fF
C34925 INVX1_LOC_95/Y NOR2X1_LOC_271/Y 0.08fF
C34926 NOR2X1_LOC_68/A NOR2X1_LOC_849/A 0.03fF
C34927 VDD INVX1_LOC_194/Y 0.21fF
C34928 NOR2X1_LOC_667/Y NAND2X1_LOC_537/Y 0.01fF
C34929 NOR2X1_LOC_667/a_36_216# NAND2X1_LOC_538/Y 0.01fF
C34930 NAND2X1_LOC_804/Y INVX1_LOC_46/A 0.07fF
C34931 NAND2X1_LOC_578/B INVX1_LOC_175/A 0.03fF
C34932 INVX1_LOC_151/A INVX1_LOC_271/A 0.01fF
C34933 INVX1_LOC_284/Y NAND2X1_LOC_561/B 0.16fF
C34934 NAND2X1_LOC_803/B INVX1_LOC_215/Y 0.04fF
C34935 INVX1_LOC_25/A NOR2X1_LOC_124/B 0.13fF
C34936 INVX1_LOC_39/A INVX1_LOC_61/A 0.09fF
C34937 INVX1_LOC_91/A INVX1_LOC_117/Y 0.05fF
C34938 INVX1_LOC_36/A NAND2X1_LOC_218/A 0.01fF
C34939 NAND2X1_LOC_468/B NOR2X1_LOC_351/Y 0.11fF
C34940 NOR2X1_LOC_78/A NOR2X1_LOC_624/B 0.01fF
C34941 NOR2X1_LOC_52/B INVX1_LOC_271/A 0.14fF
C34942 NOR2X1_LOC_290/Y NAND2X1_LOC_464/B 0.01fF
C34943 D_INPUT_7 INVX1_LOC_1/A 0.02fF
C34944 INVX1_LOC_88/Y NOR2X1_LOC_678/A 0.41fF
C34945 INVX1_LOC_223/A NOR2X1_LOC_205/Y 0.01fF
C34946 INVX1_LOC_36/A NAND2X1_LOC_538/Y 0.01fF
C34947 NOR2X1_LOC_791/A INVX1_LOC_14/A -0.02fF
C34948 NOR2X1_LOC_791/B INVX1_LOC_1/A 0.56fF
C34949 NAND2X1_LOC_9/Y INVX1_LOC_158/A 0.06fF
C34950 VDD INVX1_LOC_9/A 1.19fF
C34951 NAND2X1_LOC_725/Y INVX1_LOC_209/A 0.05fF
C34952 INVX1_LOC_35/A NOR2X1_LOC_6/B 0.04fF
C34953 D_INPUT_0 NAND2X1_LOC_761/a_36_24# 0.01fF
C34954 INVX1_LOC_201/A NAND2X1_LOC_225/a_36_24# 0.00fF
C34955 INVX1_LOC_22/A NAND2X1_LOC_61/Y 0.26fF
C34956 INVX1_LOC_103/A NOR2X1_LOC_52/Y 0.03fF
C34957 INVX1_LOC_13/Y INVX1_LOC_33/A 0.07fF
C34958 INVX1_LOC_27/A NOR2X1_LOC_433/A 0.09fF
C34959 D_GATE_366 D_INPUT_5 0.03fF
C34960 NOR2X1_LOC_15/Y NAND2X1_LOC_656/A 0.92fF
C34961 INVX1_LOC_103/A NOR2X1_LOC_270/Y 0.06fF
C34962 NOR2X1_LOC_686/B INVX1_LOC_78/A 0.01fF
C34963 NAND2X1_LOC_347/B INVX1_LOC_71/A 0.11fF
C34964 INVX1_LOC_11/Y NAND2X1_LOC_770/Y 0.05fF
C34965 NAND2X1_LOC_842/B INVX1_LOC_32/A 0.01fF
C34966 INVX1_LOC_50/A NOR2X1_LOC_165/Y 0.44fF
C34967 NOR2X1_LOC_321/Y NOR2X1_LOC_152/Y 0.02fF
C34968 INVX1_LOC_214/A INVX1_LOC_53/A 0.05fF
C34969 NAND2X1_LOC_326/A NOR2X1_LOC_152/a_36_216# 0.00fF
C34970 INVX1_LOC_27/A NOR2X1_LOC_593/Y 0.01fF
C34971 NOR2X1_LOC_667/A INVX1_LOC_53/A 0.08fF
C34972 INVX1_LOC_313/A NOR2X1_LOC_334/Y 0.02fF
C34973 NOR2X1_LOC_700/Y NAND2X1_LOC_175/Y 0.04fF
C34974 INVX1_LOC_248/A INVX1_LOC_53/A 0.07fF
C34975 INVX1_LOC_58/A NOR2X1_LOC_488/Y 0.03fF
C34976 INVX1_LOC_76/A NOR2X1_LOC_197/B 0.00fF
C34977 INVX1_LOC_132/A NAND2X1_LOC_773/Y 0.06fF
C34978 INVX1_LOC_25/A NOR2X1_LOC_646/A 0.38fF
C34979 INVX1_LOC_255/Y INVX1_LOC_57/A 0.15fF
C34980 NAND2X1_LOC_656/Y NOR2X1_LOC_318/A 0.08fF
C34981 NOR2X1_LOC_285/Y INVX1_LOC_196/A 0.06fF
C34982 NAND2X1_LOC_667/a_36_24# INVX1_LOC_50/Y 0.01fF
C34983 NOR2X1_LOC_361/B INVX1_LOC_77/A 0.10fF
C34984 NOR2X1_LOC_807/B NOR2X1_LOC_500/A 0.03fF
C34985 NOR2X1_LOC_602/A INVX1_LOC_45/A 0.01fF
C34986 NOR2X1_LOC_681/Y NOR2X1_LOC_88/Y 0.07fF
C34987 NOR2X1_LOC_331/Y INVX1_LOC_159/A 0.01fF
C34988 INVX1_LOC_249/A INVX1_LOC_11/A 0.00fF
C34989 INVX1_LOC_27/A NOR2X1_LOC_52/B 0.18fF
C34990 INVX1_LOC_285/Y INVX1_LOC_290/Y 0.10fF
C34991 NOR2X1_LOC_824/A NOR2X1_LOC_52/B 0.07fF
C34992 INVX1_LOC_256/A NOR2X1_LOC_303/Y 0.10fF
C34993 INVX1_LOC_64/A NOR2X1_LOC_500/Y 0.03fF
C34994 INVX1_LOC_88/A INVX1_LOC_33/A 0.51fF
C34995 INVX1_LOC_64/A INVX1_LOC_226/Y 0.03fF
C34996 INVX1_LOC_136/A NOR2X1_LOC_382/Y 0.04fF
C34997 NOR2X1_LOC_329/B INVX1_LOC_273/A 0.09fF
C34998 NOR2X1_LOC_598/B GATE_479 0.02fF
C34999 NOR2X1_LOC_528/Y NOR2X1_LOC_89/A 0.11fF
C35000 NAND2X1_LOC_773/Y INVX1_LOC_225/A 0.10fF
C35001 INVX1_LOC_58/A INVX1_LOC_227/A 0.10fF
C35002 INVX1_LOC_233/A NAND2X1_LOC_564/B 1.12fF
C35003 INVX1_LOC_14/A NOR2X1_LOC_121/Y 0.06fF
C35004 NOR2X1_LOC_717/B NOR2X1_LOC_858/A 0.02fF
C35005 NOR2X1_LOC_71/Y INVX1_LOC_57/A 0.12fF
C35006 NOR2X1_LOC_603/a_36_216# INVX1_LOC_27/A 0.01fF
C35007 INVX1_LOC_21/A NOR2X1_LOC_78/B 0.13fF
C35008 NOR2X1_LOC_263/a_36_216# NOR2X1_LOC_15/Y 0.00fF
C35009 INVX1_LOC_117/A NOR2X1_LOC_688/a_36_216# 0.02fF
C35010 NOR2X1_LOC_68/A INVX1_LOC_142/A 0.03fF
C35011 INVX1_LOC_37/A INVX1_LOC_84/A 0.06fF
C35012 INVX1_LOC_13/Y INVX1_LOC_40/A 0.26fF
C35013 NOR2X1_LOC_536/A INVX1_LOC_35/Y 0.05fF
C35014 NOR2X1_LOC_565/B INVX1_LOC_53/A 0.03fF
C35015 NOR2X1_LOC_554/B INVX1_LOC_205/A 0.00fF
C35016 NOR2X1_LOC_859/A NOR2X1_LOC_68/A 0.00fF
C35017 NAND2X1_LOC_763/B NAND2X1_LOC_588/B 0.01fF
C35018 NAND2X1_LOC_850/Y NAND2X1_LOC_474/Y 0.73fF
C35019 INVX1_LOC_13/Y INVX1_LOC_165/Y 0.03fF
C35020 NOR2X1_LOC_107/Y INVX1_LOC_8/A 0.00fF
C35021 INVX1_LOC_107/Y INVX1_LOC_38/A 0.03fF
C35022 INPUT_0 INVX1_LOC_94/Y 0.03fF
C35023 NAND2X1_LOC_656/Y NOR2X1_LOC_678/A 0.02fF
C35024 NOR2X1_LOC_356/A NOR2X1_LOC_383/B 0.19fF
C35025 NOR2X1_LOC_828/A NOR2X1_LOC_858/A 0.33fF
C35026 INVX1_LOC_34/A INVX1_LOC_293/A 0.01fF
C35027 INVX1_LOC_11/A NAND2X1_LOC_26/a_36_24# 0.00fF
C35028 INVX1_LOC_64/A INVX1_LOC_10/A 1.98fF
C35029 INVX1_LOC_147/Y INVX1_LOC_12/A 0.01fF
C35030 INVX1_LOC_1/A NOR2X1_LOC_767/a_36_216# 0.00fF
C35031 NAND2X1_LOC_721/A INVX1_LOC_203/A 0.34fF
C35032 NOR2X1_LOC_479/B INVX1_LOC_178/A 0.01fF
C35033 NOR2X1_LOC_644/Y NAND2X1_LOC_190/Y 0.07fF
C35034 NOR2X1_LOC_392/B INVX1_LOC_150/Y 0.02fF
C35035 INVX1_LOC_6/A NOR2X1_LOC_334/Y 0.07fF
C35036 NOR2X1_LOC_272/Y INVX1_LOC_16/A 0.00fF
C35037 NAND2X1_LOC_151/a_36_24# NOR2X1_LOC_52/B 0.00fF
C35038 NOR2X1_LOC_328/Y INVX1_LOC_178/A 0.06fF
C35039 INVX1_LOC_12/A INVX1_LOC_20/A 0.15fF
C35040 INVX1_LOC_37/A NAND2X1_LOC_651/B 0.01fF
C35041 NOR2X1_LOC_598/B INVX1_LOC_196/Y 1.80fF
C35042 INPUT_4 NOR2X1_LOC_59/a_36_216# 0.00fF
C35043 INVX1_LOC_219/A INVX1_LOC_5/A 0.03fF
C35044 NOR2X1_LOC_78/A NOR2X1_LOC_38/B 0.00fF
C35045 INVX1_LOC_256/A INVX1_LOC_54/Y 0.07fF
C35046 INVX1_LOC_33/A NOR2X1_LOC_500/B 0.02fF
C35047 NOR2X1_LOC_471/Y INVX1_LOC_266/Y 1.03fF
C35048 NOR2X1_LOC_68/A NAND2X1_LOC_593/Y 0.07fF
C35049 NOR2X1_LOC_536/A NOR2X1_LOC_721/B 0.01fF
C35050 INVX1_LOC_58/A NOR2X1_LOC_741/a_36_216# 0.00fF
C35051 INVX1_LOC_224/A NAND2X1_LOC_200/B 0.05fF
C35052 INPUT_0 INVX1_LOC_181/A 0.68fF
C35053 INVX1_LOC_21/A NOR2X1_LOC_459/A 0.03fF
C35054 NOR2X1_LOC_74/A NOR2X1_LOC_383/B 0.26fF
C35055 INVX1_LOC_255/Y NOR2X1_LOC_475/A 0.03fF
C35056 INVX1_LOC_5/A NOR2X1_LOC_130/a_36_216# 0.00fF
C35057 NOR2X1_LOC_793/Y NOR2X1_LOC_325/A 0.04fF
C35058 NAND2X1_LOC_208/B NOR2X1_LOC_315/Y 0.03fF
C35059 INVX1_LOC_91/A INVX1_LOC_87/A 0.03fF
C35060 INVX1_LOC_50/A NOR2X1_LOC_527/Y 0.15fF
C35061 NOR2X1_LOC_655/B NOR2X1_LOC_160/B 0.10fF
C35062 NAND2X1_LOC_745/a_36_24# NOR2X1_LOC_781/A 0.00fF
C35063 INVX1_LOC_21/A INVX1_LOC_83/A 1.59fF
C35064 NOR2X1_LOC_623/a_36_216# NAND2X1_LOC_364/A 0.00fF
C35065 VDD NOR2X1_LOC_861/Y 0.31fF
C35066 INVX1_LOC_37/A NAND2X1_LOC_220/B 0.10fF
C35067 NOR2X1_LOC_79/A INVX1_LOC_294/A 0.00fF
C35068 NOR2X1_LOC_9/Y NOR2X1_LOC_383/B 0.07fF
C35069 NAND2X1_LOC_577/A NAND2X1_LOC_141/A 0.08fF
C35070 NAND2X1_LOC_649/B INVX1_LOC_94/Y 0.20fF
C35071 NAND2X1_LOC_860/Y NAND2X1_LOC_793/Y 0.01fF
C35072 INVX1_LOC_38/A INVX1_LOC_272/A 0.17fF
C35073 INVX1_LOC_33/A NOR2X1_LOC_170/a_36_216# 0.00fF
C35074 NAND2X1_LOC_51/B INVX1_LOC_53/A 0.04fF
C35075 INVX1_LOC_281/A NAND2X1_LOC_469/a_36_24# 0.00fF
C35076 INVX1_LOC_133/A INVX1_LOC_9/A 0.22fF
C35077 VDD NOR2X1_LOC_812/A 0.24fF
C35078 NOR2X1_LOC_662/A NAND2X1_LOC_243/Y 0.01fF
C35079 INVX1_LOC_254/A INVX1_LOC_49/A 0.01fF
C35080 INVX1_LOC_14/Y INVX1_LOC_257/A 0.00fF
C35081 INVX1_LOC_36/A NOR2X1_LOC_709/A 8.77fF
C35082 NOR2X1_LOC_453/Y INVX1_LOC_83/A 0.03fF
C35083 INVX1_LOC_249/A NOR2X1_LOC_593/Y 0.19fF
C35084 D_GATE_222 INVX1_LOC_174/A -0.03fF
C35085 INVX1_LOC_37/A INVX1_LOC_15/A 0.28fF
C35086 NOR2X1_LOC_82/A INVX1_LOC_137/Y 0.01fF
C35087 NOR2X1_LOC_274/Y NOR2X1_LOC_557/Y 0.02fF
C35088 NAND2X1_LOC_361/Y NOR2X1_LOC_419/Y 0.02fF
C35089 NOR2X1_LOC_231/A INVX1_LOC_15/A 0.03fF
C35090 NOR2X1_LOC_92/Y NOR2X1_LOC_76/A 0.09fF
C35091 NOR2X1_LOC_441/Y INVX1_LOC_208/A 0.27fF
C35092 NOR2X1_LOC_272/Y INVX1_LOC_28/A 0.10fF
C35093 D_INPUT_0 INVX1_LOC_14/A 0.23fF
C35094 INVX1_LOC_305/A NOR2X1_LOC_168/B 0.12fF
C35095 NAND2X1_LOC_361/Y NOR2X1_LOC_716/B 0.03fF
C35096 INVX1_LOC_239/A INVX1_LOC_175/Y 0.38fF
C35097 VDD INVX1_LOC_274/Y 0.13fF
C35098 INVX1_LOC_90/A INVX1_LOC_198/A 0.02fF
C35099 INVX1_LOC_5/A NOR2X1_LOC_196/Y 0.01fF
C35100 NAND2X1_LOC_581/Y INVX1_LOC_77/A 0.01fF
C35101 NOR2X1_LOC_790/B NOR2X1_LOC_794/A 0.02fF
C35102 INVX1_LOC_49/A NAND2X1_LOC_466/Y 0.01fF
C35103 NOR2X1_LOC_655/Y NOR2X1_LOC_610/Y 0.01fF
C35104 NAND2X1_LOC_475/Y INVX1_LOC_285/A 0.01fF
C35105 INVX1_LOC_249/A NOR2X1_LOC_52/B 0.03fF
C35106 INVX1_LOC_78/Y NOR2X1_LOC_678/A 2.07fF
C35107 NAND2X1_LOC_475/Y NOR2X1_LOC_814/A 0.01fF
C35108 NAND2X1_LOC_861/Y NAND2X1_LOC_793/Y 0.01fF
C35109 NOR2X1_LOC_186/Y NAND2X1_LOC_858/B 0.03fF
C35110 INVX1_LOC_77/A INVX1_LOC_177/A 0.06fF
C35111 NOR2X1_LOC_593/a_36_216# INVX1_LOC_113/Y 0.00fF
C35112 NAND2X1_LOC_733/Y INVX1_LOC_229/Y 0.03fF
C35113 INVX1_LOC_286/Y NOR2X1_LOC_561/Y 0.07fF
C35114 NOR2X1_LOC_312/Y NAND2X1_LOC_336/a_36_24# 0.06fF
C35115 NAND2X1_LOC_510/A NAND2X1_LOC_41/Y 0.07fF
C35116 INVX1_LOC_245/A INVX1_LOC_18/A 0.11fF
C35117 NOR2X1_LOC_274/Y INVX1_LOC_143/A -0.03fF
C35118 INVX1_LOC_133/Y NOR2X1_LOC_577/Y 0.20fF
C35119 NAND2X1_LOC_364/A INVX1_LOC_16/A 0.09fF
C35120 INVX1_LOC_157/Y INVX1_LOC_15/A -0.01fF
C35121 INVX1_LOC_34/A NOR2X1_LOC_315/Y 0.10fF
C35122 INVX1_LOC_276/A NOR2X1_LOC_577/Y 0.62fF
C35123 INVX1_LOC_181/Y INVX1_LOC_25/Y 0.02fF
C35124 NOR2X1_LOC_177/Y INVX1_LOC_15/A 0.06fF
C35125 NAND2X1_LOC_573/Y NAND2X1_LOC_858/B -0.00fF
C35126 INVX1_LOC_2/A NOR2X1_LOC_690/A 0.03fF
C35127 NOR2X1_LOC_743/Y INVX1_LOC_15/A 0.06fF
C35128 INVX1_LOC_125/A INVX1_LOC_63/A 0.03fF
C35129 NOR2X1_LOC_432/Y INVX1_LOC_34/A 0.04fF
C35130 INVX1_LOC_299/A INPUT_0 0.03fF
C35131 INVX1_LOC_25/A INVX1_LOC_2/Y 0.10fF
C35132 INVX1_LOC_217/A INVX1_LOC_229/Y 0.07fF
C35133 NOR2X1_LOC_420/Y NOR2X1_LOC_78/A 0.01fF
C35134 NOR2X1_LOC_309/Y NOR2X1_LOC_709/A 0.01fF
C35135 INVX1_LOC_3/A NOR2X1_LOC_610/Y 0.01fF
C35136 NOR2X1_LOC_89/A NAND2X1_LOC_477/Y 0.11fF
C35137 NOR2X1_LOC_791/Y INVX1_LOC_70/Y 0.02fF
C35138 INVX1_LOC_307/A INVX1_LOC_4/A 0.07fF
C35139 NAND2X1_LOC_33/Y NAND2X1_LOC_35/a_36_24# 0.00fF
C35140 NOR2X1_LOC_536/A NAND2X1_LOC_286/B 0.08fF
C35141 NOR2X1_LOC_261/Y INVX1_LOC_37/A 0.17fF
C35142 INVX1_LOC_21/A NOR2X1_LOC_311/Y 0.02fF
C35143 NOR2X1_LOC_423/Y INVX1_LOC_96/Y 0.01fF
C35144 INVX1_LOC_34/A INVX1_LOC_52/A 0.01fF
C35145 NOR2X1_LOC_445/B INVX1_LOC_4/A 0.07fF
C35146 NAND2X1_LOC_472/Y INVX1_LOC_23/A 0.11fF
C35147 NAND2X1_LOC_35/Y NAND2X1_LOC_836/Y -0.01fF
C35148 INVX1_LOC_208/A NOR2X1_LOC_142/Y 0.12fF
C35149 INVX1_LOC_234/Y NOR2X1_LOC_45/B 0.01fF
C35150 INVX1_LOC_278/A INVX1_LOC_37/A 0.07fF
C35151 INVX1_LOC_269/A NOR2X1_LOC_501/B 0.01fF
C35152 INVX1_LOC_45/A NOR2X1_LOC_564/Y 0.03fF
C35153 NOR2X1_LOC_788/B INVX1_LOC_18/A 0.01fF
C35154 NOR2X1_LOC_468/Y INVX1_LOC_98/A 0.07fF
C35155 INVX1_LOC_27/A INVX1_LOC_199/A 0.07fF
C35156 NOR2X1_LOC_506/a_36_216# INVX1_LOC_53/A 0.02fF
C35157 NAND2X1_LOC_84/Y D_INPUT_0 0.05fF
C35158 NOR2X1_LOC_686/B NOR2X1_LOC_152/Y 0.03fF
C35159 INVX1_LOC_279/A NOR2X1_LOC_374/A 0.05fF
C35160 NOR2X1_LOC_468/Y NOR2X1_LOC_78/A 0.03fF
C35161 NOR2X1_LOC_251/Y NOR2X1_LOC_52/B 0.00fF
C35162 INVX1_LOC_145/A NOR2X1_LOC_106/A 0.12fF
C35163 NOR2X1_LOC_222/Y INVX1_LOC_96/Y 0.07fF
C35164 NAND2X1_LOC_156/B NOR2X1_LOC_433/A 0.07fF
C35165 NAND2X1_LOC_860/A NOR2X1_LOC_536/A 0.07fF
C35166 INVX1_LOC_27/A INVX1_LOC_74/A 0.01fF
C35167 NAND2X1_LOC_773/Y NAND2X1_LOC_642/Y 0.10fF
C35168 NOR2X1_LOC_657/a_36_216# NAND2X1_LOC_469/B 0.00fF
C35169 INVX1_LOC_36/A NAND2X1_LOC_863/A 0.07fF
C35170 NOR2X1_LOC_68/A NOR2X1_LOC_535/a_36_216# 0.14fF
C35171 NOR2X1_LOC_299/Y NAND2X1_LOC_838/a_36_24# 0.01fF
C35172 NAND2X1_LOC_785/A INVX1_LOC_16/A 0.10fF
C35173 NOR2X1_LOC_82/A INVX1_LOC_91/A 0.00fF
C35174 INVX1_LOC_164/A INVX1_LOC_8/A 0.03fF
C35175 NOR2X1_LOC_413/Y NAND2X1_LOC_462/B 0.06fF
C35176 INVX1_LOC_63/Y NOR2X1_LOC_366/Y 0.05fF
C35177 INVX1_LOC_177/A NOR2X1_LOC_687/Y 0.03fF
C35178 INVX1_LOC_21/A INVX1_LOC_46/A 0.59fF
C35179 INVX1_LOC_57/Y NOR2X1_LOC_74/A 0.11fF
C35180 INVX1_LOC_286/Y NOR2X1_LOC_167/Y 0.00fF
C35181 INVX1_LOC_34/A INVX1_LOC_66/A 0.01fF
C35182 NOR2X1_LOC_627/Y INVX1_LOC_16/A 0.05fF
C35183 NOR2X1_LOC_655/B NOR2X1_LOC_516/B 0.12fF
C35184 INVX1_LOC_217/Y D_INPUT_0 -0.00fF
C35185 INVX1_LOC_119/Y NAND2X1_LOC_175/Y 0.02fF
C35186 NOR2X1_LOC_778/B NOR2X1_LOC_439/a_36_216# 0.00fF
C35187 NOR2X1_LOC_32/B NOR2X1_LOC_629/Y 0.06fF
C35188 NOR2X1_LOC_598/B NOR2X1_LOC_641/Y 0.01fF
C35189 INVX1_LOC_234/A NOR2X1_LOC_52/B 0.19fF
C35190 NAND2X1_LOC_514/Y INVX1_LOC_79/A 0.01fF
C35191 INVX1_LOC_13/A NOR2X1_LOC_537/Y 0.07fF
C35192 NOR2X1_LOC_680/a_36_216# NOR2X1_LOC_678/A 0.00fF
C35193 INVX1_LOC_181/Y INVX1_LOC_75/A 0.12fF
C35194 INVX1_LOC_177/A NOR2X1_LOC_549/a_36_216# 0.00fF
C35195 NOR2X1_LOC_440/Y INVX1_LOC_54/Y -0.00fF
C35196 NOR2X1_LOC_748/Y NOR2X1_LOC_539/a_36_216# 0.00fF
C35197 INVX1_LOC_13/A NAND2X1_LOC_338/B 0.30fF
C35198 NOR2X1_LOC_389/A NOR2X1_LOC_78/A 0.01fF
C35199 NOR2X1_LOC_301/A NOR2X1_LOC_653/Y 0.01fF
C35200 INVX1_LOC_27/Y INVX1_LOC_23/Y 0.04fF
C35201 INVX1_LOC_135/A NAND2X1_LOC_357/B 0.10fF
C35202 INVX1_LOC_32/A INVX1_LOC_284/A 0.14fF
C35203 NOR2X1_LOC_643/A INVX1_LOC_20/A 0.15fF
C35204 INVX1_LOC_41/A NOR2X1_LOC_180/B 0.01fF
C35205 NAND2X1_LOC_860/A NAND2X1_LOC_93/B 0.21fF
C35206 INVX1_LOC_178/A INVX1_LOC_33/Y 0.05fF
C35207 NOR2X1_LOC_160/B NOR2X1_LOC_502/a_36_216# 0.00fF
C35208 NAND2X1_LOC_543/Y NAND2X1_LOC_862/A 0.01fF
C35209 NOR2X1_LOC_690/A INPUT_1 0.01fF
C35210 INVX1_LOC_90/A NOR2X1_LOC_770/B 0.02fF
C35211 INVX1_LOC_203/A INVX1_LOC_175/A 0.02fF
C35212 NOR2X1_LOC_474/A NOR2X1_LOC_19/B 0.00fF
C35213 NAND2X1_LOC_67/Y NOR2X1_LOC_69/a_36_216# 0.01fF
C35214 NAND2X1_LOC_67/Y VDD 0.24fF
C35215 NOR2X1_LOC_565/A NOR2X1_LOC_337/Y 0.20fF
C35216 INVX1_LOC_12/A INVX1_LOC_4/A 2.18fF
C35217 NOR2X1_LOC_15/Y NAND2X1_LOC_611/a_36_24# 0.00fF
C35218 INVX1_LOC_14/A NOR2X1_LOC_266/B 0.33fF
C35219 NAND2X1_LOC_500/Y INVX1_LOC_91/A 0.01fF
C35220 NAND2X1_LOC_456/Y NAND2X1_LOC_99/A 0.01fF
C35221 INVX1_LOC_13/A NAND2X1_LOC_323/B 0.26fF
C35222 NAND2X1_LOC_708/Y NOR2X1_LOC_51/A 0.00fF
C35223 NOR2X1_LOC_468/Y NOR2X1_LOC_176/a_36_216# 0.00fF
C35224 INVX1_LOC_47/Y INVX1_LOC_42/A 0.42fF
C35225 NAND2X1_LOC_477/A NOR2X1_LOC_76/A 0.12fF
C35226 NAND2X1_LOC_218/a_36_24# INVX1_LOC_3/A 0.01fF
C35227 NOR2X1_LOC_30/Y NOR2X1_LOC_11/Y 0.00fF
C35228 INVX1_LOC_147/A NAND2X1_LOC_593/Y 0.01fF
C35229 NOR2X1_LOC_340/A NAND2X1_LOC_226/a_36_24# 0.00fF
C35230 INVX1_LOC_194/A NAND2X1_LOC_622/a_36_24# 0.00fF
C35231 NOR2X1_LOC_301/A INVX1_LOC_19/A 0.04fF
C35232 NOR2X1_LOC_92/Y NAND2X1_LOC_837/a_36_24# 0.00fF
C35233 NAND2X1_LOC_20/B VDD 0.01fF
C35234 INVX1_LOC_64/A INVX1_LOC_307/A 0.22fF
C35235 NAND2X1_LOC_579/A NOR2X1_LOC_492/Y 0.03fF
C35236 NOR2X1_LOC_91/A NAND2X1_LOC_773/B 0.03fF
C35237 INVX1_LOC_16/A NOR2X1_LOC_86/A 0.59fF
C35238 INVX1_LOC_41/A INVX1_LOC_73/A 0.03fF
C35239 NOR2X1_LOC_500/A INVX1_LOC_69/Y 0.02fF
C35240 INVX1_LOC_64/A NOR2X1_LOC_445/B 0.07fF
C35241 INVX1_LOC_69/Y NOR2X1_LOC_303/Y 0.10fF
C35242 NOR2X1_LOC_317/A NOR2X1_LOC_78/A 0.02fF
C35243 NOR2X1_LOC_331/Y INVX1_LOC_146/Y 0.02fF
C35244 INVX1_LOC_77/A INVX1_LOC_285/Y 0.01fF
C35245 NAND2X1_LOC_785/A INVX1_LOC_28/A 0.07fF
C35246 NAND2X1_LOC_308/Y NAND2X1_LOC_740/B 0.00fF
C35247 NAND2X1_LOC_551/A NAND2X1_LOC_338/B 0.12fF
C35248 NAND2X1_LOC_733/Y INVX1_LOC_20/A 0.07fF
C35249 NOR2X1_LOC_48/a_36_216# INVX1_LOC_296/A 0.01fF
C35250 NAND2X1_LOC_537/Y NOR2X1_LOC_536/A 0.32fF
C35251 NAND2X1_LOC_773/Y NOR2X1_LOC_271/Y 0.03fF
C35252 INVX1_LOC_14/A NAND2X1_LOC_848/A 0.10fF
C35253 NOR2X1_LOC_355/B INVX1_LOC_94/A 0.07fF
C35254 NOR2X1_LOC_331/Y VDD 0.17fF
C35255 INVX1_LOC_193/Y NOR2X1_LOC_550/B 0.00fF
C35256 INVX1_LOC_171/A NOR2X1_LOC_566/Y 0.01fF
C35257 NOR2X1_LOC_635/A D_INPUT_4 0.01fF
C35258 NAND2X1_LOC_705/Y INVX1_LOC_118/A 0.14fF
C35259 NAND2X1_LOC_80/a_36_24# NAND2X1_LOC_99/A 0.00fF
C35260 NOR2X1_LOC_168/A NOR2X1_LOC_356/A 0.02fF
C35261 NAND2X1_LOC_858/B NAND2X1_LOC_640/Y -0.00fF
C35262 NOR2X1_LOC_778/B NOR2X1_LOC_724/Y 0.45fF
C35263 NOR2X1_LOC_516/B NOR2X1_LOC_99/B 0.10fF
C35264 NAND2X1_LOC_639/a_36_24# NOR2X1_LOC_635/B 0.00fF
C35265 INVX1_LOC_286/Y INVX1_LOC_76/A 0.09fF
C35266 NOR2X1_LOC_626/Y INVX1_LOC_92/A 0.04fF
C35267 NOR2X1_LOC_441/Y NAND2X1_LOC_211/Y 0.21fF
C35268 INVX1_LOC_23/A NAND2X1_LOC_773/B 1.28fF
C35269 NOR2X1_LOC_368/A INVX1_LOC_8/A 0.35fF
C35270 NAND2X1_LOC_337/B INVX1_LOC_33/Y 0.03fF
C35271 NAND2X1_LOC_363/B NOR2X1_LOC_814/A 0.07fF
C35272 INVX1_LOC_314/Y NOR2X1_LOC_557/A 0.07fF
C35273 INVX1_LOC_5/A NAND2X1_LOC_52/a_36_24# 0.00fF
C35274 NOR2X1_LOC_361/B INVX1_LOC_9/A 0.05fF
C35275 INVX1_LOC_2/A NOR2X1_LOC_736/a_36_216# 0.00fF
C35276 NAND2X1_LOC_179/a_36_24# NAND2X1_LOC_472/Y 0.00fF
C35277 NAND2X1_LOC_162/a_36_24# NAND2X1_LOC_451/Y 0.01fF
C35278 NOR2X1_LOC_321/Y INVX1_LOC_291/A -0.01fF
C35279 INVX1_LOC_225/A NAND2X1_LOC_858/B 0.09fF
C35280 NOR2X1_LOC_530/a_36_216# NOR2X1_LOC_536/A 0.00fF
C35281 NOR2X1_LOC_516/B NOR2X1_LOC_846/B 0.01fF
C35282 INVX1_LOC_88/A NOR2X1_LOC_351/Y 0.01fF
C35283 INVX1_LOC_18/A NAND2X1_LOC_1/Y 0.33fF
C35284 NOR2X1_LOC_565/A VDD 0.24fF
C35285 NOR2X1_LOC_315/Y INPUT_0 0.32fF
C35286 INVX1_LOC_217/A INVX1_LOC_20/A 0.05fF
C35287 NAND2X1_LOC_364/A NOR2X1_LOC_35/Y 0.10fF
C35288 NOR2X1_LOC_289/a_36_216# INVX1_LOC_28/A 0.00fF
C35289 INVX1_LOC_185/Y NOR2X1_LOC_167/Y 0.01fF
C35290 INVX1_LOC_72/A NOR2X1_LOC_357/Y 0.07fF
C35291 NOR2X1_LOC_169/B VDD -0.00fF
C35292 NAND2X1_LOC_348/A NOR2X1_LOC_87/Y -0.01fF
C35293 NOR2X1_LOC_718/B INVX1_LOC_6/A 0.28fF
C35294 NOR2X1_LOC_329/B NAND2X1_LOC_840/B 0.39fF
C35295 NAND2X1_LOC_12/a_36_24# NAND2X1_LOC_1/Y 0.00fF
C35296 NOR2X1_LOC_791/Y INVX1_LOC_285/A 0.03fF
C35297 INVX1_LOC_90/A NAND2X1_LOC_168/a_36_24# 0.00fF
C35298 INVX1_LOC_77/A INVX1_LOC_65/A 0.08fF
C35299 INVX1_LOC_159/A INVX1_LOC_76/A 0.54fF
C35300 INVX1_LOC_18/A NAND2X1_LOC_39/Y 0.02fF
C35301 INVX1_LOC_124/A INVX1_LOC_285/Y 0.02fF
C35302 INVX1_LOC_14/A INVX1_LOC_46/Y 0.10fF
C35303 INVX1_LOC_190/Y NOR2X1_LOC_561/Y 0.04fF
C35304 INVX1_LOC_144/Y INVX1_LOC_144/A 0.10fF
C35305 NOR2X1_LOC_328/Y INVX1_LOC_140/A 0.05fF
C35306 NOR2X1_LOC_516/B NOR2X1_LOC_381/a_36_216# 0.00fF
C35307 INVX1_LOC_77/A NOR2X1_LOC_137/B 0.09fF
C35308 INVX1_LOC_211/Y NOR2X1_LOC_506/Y 0.13fF
C35309 NOR2X1_LOC_65/B INVX1_LOC_47/Y 0.09fF
C35310 NOR2X1_LOC_91/A NOR2X1_LOC_393/Y 0.03fF
C35311 VDD NOR2X1_LOC_324/Y 0.02fF
C35312 INVX1_LOC_54/Y INVX1_LOC_69/Y 0.01fF
C35313 NOR2X1_LOC_168/Y INVX1_LOC_37/A 0.03fF
C35314 INVX1_LOC_124/A NOR2X1_LOC_183/a_36_216# 0.00fF
C35315 NOR2X1_LOC_78/B INVX1_LOC_311/A 0.08fF
C35316 NOR2X1_LOC_649/B NAND2X1_LOC_473/A 0.17fF
C35317 INVX1_LOC_64/A INVX1_LOC_12/A 4.59fF
C35318 INVX1_LOC_3/A NAND2X1_LOC_473/A 0.91fF
C35319 INVX1_LOC_64/A NOR2X1_LOC_519/Y 0.03fF
C35320 INVX1_LOC_78/A NOR2X1_LOC_693/a_36_216# 0.00fF
C35321 INVX1_LOC_72/A INVX1_LOC_66/Y 0.08fF
C35322 INVX1_LOC_72/A NOR2X1_LOC_692/Y 0.08fF
C35323 INVX1_LOC_119/A NAND2X1_LOC_655/A 0.10fF
C35324 NAND2X1_LOC_787/B INVX1_LOC_20/A 0.03fF
C35325 NOR2X1_LOC_635/a_36_216# NOR2X1_LOC_48/B 0.00fF
C35326 NAND2X1_LOC_170/A NOR2X1_LOC_74/A 0.04fF
C35327 NOR2X1_LOC_843/A INVX1_LOC_314/A 0.05fF
C35328 INVX1_LOC_62/Y NOR2X1_LOC_98/a_36_216# 0.00fF
C35329 INVX1_LOC_63/A NAND2X1_LOC_218/A 0.01fF
C35330 NOR2X1_LOC_393/Y INVX1_LOC_23/A 0.01fF
C35331 NOR2X1_LOC_334/Y INVX1_LOC_270/A 0.10fF
C35332 NOR2X1_LOC_852/B VDD 0.14fF
C35333 NAND2X1_LOC_395/a_36_24# INVX1_LOC_98/A 0.00fF
C35334 NAND2X1_LOC_785/Y NOR2X1_LOC_164/Y 0.01fF
C35335 INVX1_LOC_55/Y INVX1_LOC_313/Y 0.07fF
C35336 NAND2X1_LOC_493/a_36_24# INVX1_LOC_309/A 0.00fF
C35337 INVX1_LOC_21/A NOR2X1_LOC_671/Y 0.03fF
C35338 INVX1_LOC_50/Y NAND2X1_LOC_206/B 0.01fF
C35339 NAND2X1_LOC_21/Y INVX1_LOC_37/A 0.01fF
C35340 INVX1_LOC_248/A NOR2X1_LOC_311/Y 0.01fF
C35341 INVX1_LOC_278/Y INVX1_LOC_91/A 0.07fF
C35342 INVX1_LOC_83/A NAND2X1_LOC_51/B 0.10fF
C35343 NOR2X1_LOC_332/A NOR2X1_LOC_196/Y 0.01fF
C35344 INVX1_LOC_30/A NOR2X1_LOC_364/A 0.02fF
C35345 INVX1_LOC_53/A NOR2X1_LOC_248/A 0.01fF
C35346 INVX1_LOC_96/Y NOR2X1_LOC_69/A 0.10fF
C35347 NOR2X1_LOC_250/A INVX1_LOC_63/A 0.06fF
C35348 NOR2X1_LOC_65/B NAND2X1_LOC_211/a_36_24# 0.00fF
C35349 NOR2X1_LOC_68/A INVX1_LOC_185/A 0.00fF
C35350 NAND2X1_LOC_785/Y INVX1_LOC_46/A 0.03fF
C35351 NOR2X1_LOC_824/A NAND2X1_LOC_254/Y 0.09fF
C35352 INVX1_LOC_17/A INVX1_LOC_19/A 2.13fF
C35353 INVX1_LOC_124/A NAND2X1_LOC_267/B 0.18fF
C35354 INVX1_LOC_83/A INVX1_LOC_311/A 0.06fF
C35355 INPUT_6 NOR2X1_LOC_36/A 0.05fF
C35356 NAND2X1_LOC_629/Y VDD 0.40fF
C35357 NOR2X1_LOC_590/A NAND2X1_LOC_475/Y 0.05fF
C35358 INVX1_LOC_57/A NOR2X1_LOC_39/Y 0.19fF
C35359 NOR2X1_LOC_122/Y INVX1_LOC_73/A 0.01fF
C35360 NOR2X1_LOC_405/A INVX1_LOC_16/A 0.03fF
C35361 NOR2X1_LOC_490/Y NAND2X1_LOC_849/A 0.01fF
C35362 INVX1_LOC_50/A NOR2X1_LOC_654/A 0.00fF
C35363 INVX1_LOC_224/Y NOR2X1_LOC_646/B 0.10fF
C35364 D_INPUT_0 INVX1_LOC_48/A 0.50fF
C35365 INVX1_LOC_30/A INVX1_LOC_285/A 0.66fF
C35366 INVX1_LOC_104/A INVX1_LOC_117/A 0.48fF
C35367 NOR2X1_LOC_471/Y INVX1_LOC_19/A 0.02fF
C35368 INVX1_LOC_30/A INVX1_LOC_265/Y 0.01fF
C35369 NOR2X1_LOC_770/B INVX1_LOC_38/A 0.04fF
C35370 NOR2X1_LOC_637/B INVX1_LOC_54/A 0.07fF
C35371 INVX1_LOC_64/A NOR2X1_LOC_29/a_36_216# 0.00fF
C35372 NOR2X1_LOC_667/A INVX1_LOC_46/A 0.17fF
C35373 INPUT_0 NOR2X1_LOC_166/Y 0.04fF
C35374 INVX1_LOC_179/Y VDD 0.20fF
C35375 INVX1_LOC_30/A NOR2X1_LOC_814/A 0.32fF
C35376 INVX1_LOC_31/A NAND2X1_LOC_773/B 0.07fF
C35377 INVX1_LOC_248/A INVX1_LOC_46/A 0.03fF
C35378 NOR2X1_LOC_205/Y INVX1_LOC_290/Y 0.02fF
C35379 NAND2X1_LOC_84/Y INVX1_LOC_46/Y -0.00fF
C35380 INVX1_LOC_155/A INVX1_LOC_54/A 2.51fF
C35381 NOR2X1_LOC_690/A INVX1_LOC_118/A 0.32fF
C35382 NAND2X1_LOC_374/Y NAND2X1_LOC_721/A 0.07fF
C35383 INVX1_LOC_257/Y NOR2X1_LOC_684/Y -0.01fF
C35384 INVX1_LOC_304/A NAND2X1_LOC_392/Y 0.02fF
C35385 NAND2X1_LOC_363/Y NOR2X1_LOC_836/B 0.03fF
C35386 INVX1_LOC_25/A INVX1_LOC_29/Y 0.94fF
C35387 INVX1_LOC_230/Y INVX1_LOC_29/A 0.09fF
C35388 INVX1_LOC_43/Y INVX1_LOC_12/A 0.05fF
C35389 INVX1_LOC_50/A INVX1_LOC_58/Y 0.07fF
C35390 NOR2X1_LOC_647/B NOR2X1_LOC_610/Y 0.00fF
C35391 INVX1_LOC_132/A NOR2X1_LOC_624/B 0.04fF
C35392 INVX1_LOC_33/A NOR2X1_LOC_99/Y 1.05fF
C35393 NOR2X1_LOC_561/Y NOR2X1_LOC_56/Y 0.02fF
C35394 NOR2X1_LOC_375/Y VDD 0.40fF
C35395 NOR2X1_LOC_558/A INVX1_LOC_22/A 0.01fF
C35396 NOR2X1_LOC_254/A NOR2X1_LOC_833/B 0.11fF
C35397 NOR2X1_LOC_679/Y INVX1_LOC_42/A 0.02fF
C35398 NOR2X1_LOC_773/Y INVX1_LOC_33/Y 0.02fF
C35399 NOR2X1_LOC_74/Y NOR2X1_LOC_74/A 0.00fF
C35400 INVX1_LOC_234/A INVX1_LOC_74/A 0.05fF
C35401 NOR2X1_LOC_576/B INPUT_4 0.01fF
C35402 NOR2X1_LOC_172/Y NOR2X1_LOC_58/a_36_216# 0.00fF
C35403 INVX1_LOC_177/A INVX1_LOC_9/A 0.04fF
C35404 INPUT_3 NOR2X1_LOC_643/a_36_216# 0.01fF
C35405 NAND2X1_LOC_549/B INVX1_LOC_280/A 0.10fF
C35406 INVX1_LOC_33/A INVX1_LOC_107/Y 0.03fF
C35407 NOR2X1_LOC_717/A NOR2X1_LOC_678/A 0.00fF
C35408 NOR2X1_LOC_561/Y VDD 4.38fF
C35409 NAND2X1_LOC_808/A INVX1_LOC_20/A 0.01fF
C35410 INVX1_LOC_7/A VDD 0.93fF
C35411 INVX1_LOC_89/A NOR2X1_LOC_683/Y 0.01fF
C35412 INVX1_LOC_28/A NOR2X1_LOC_405/A 0.03fF
C35413 INVX1_LOC_35/A NOR2X1_LOC_434/A 0.01fF
C35414 NOR2X1_LOC_52/B NOR2X1_LOC_216/B 0.18fF
C35415 INVX1_LOC_259/A INVX1_LOC_92/A 0.03fF
C35416 NAND2X1_LOC_850/A INVX1_LOC_95/A 0.00fF
C35417 NOR2X1_LOC_456/Y INVX1_LOC_50/Y 0.16fF
C35418 NAND2X1_LOC_717/a_36_24# INVX1_LOC_118/A 0.00fF
C35419 NOR2X1_LOC_325/A NOR2X1_LOC_729/A 0.03fF
C35420 NOR2X1_LOC_516/Y NOR2X1_LOC_649/B 0.02fF
C35421 NOR2X1_LOC_67/A NOR2X1_LOC_88/A 0.01fF
C35422 NOR2X1_LOC_679/Y INVX1_LOC_78/A 0.05fF
C35423 NOR2X1_LOC_19/B INVX1_LOC_74/A 0.00fF
C35424 NOR2X1_LOC_229/Y INVX1_LOC_54/A 0.02fF
C35425 NOR2X1_LOC_708/Y VDD 0.12fF
C35426 INVX1_LOC_40/A NOR2X1_LOC_99/Y 0.02fF
C35427 INVX1_LOC_17/A INVX1_LOC_26/Y 0.09fF
C35428 NAND2X1_LOC_9/Y INVX1_LOC_21/A 0.09fF
C35429 NOR2X1_LOC_309/Y INVX1_LOC_294/A 0.01fF
C35430 NOR2X1_LOC_32/B NOR2X1_LOC_93/Y 0.04fF
C35431 INVX1_LOC_77/A NOR2X1_LOC_830/Y 0.01fF
C35432 INVX1_LOC_170/A NOR2X1_LOC_38/B 0.04fF
C35433 INVX1_LOC_21/A INVX1_LOC_233/A 0.14fF
C35434 INVX1_LOC_303/A INVX1_LOC_106/Y 0.00fF
C35435 INVX1_LOC_33/A INVX1_LOC_272/A 0.07fF
C35436 INVX1_LOC_1/A INVX1_LOC_29/Y 0.03fF
C35437 NOR2X1_LOC_250/A NOR2X1_LOC_65/Y 0.00fF
C35438 INVX1_LOC_75/A INVX1_LOC_115/A 0.05fF
C35439 INVX1_LOC_36/A NOR2X1_LOC_334/Y 0.07fF
C35440 NAND2X1_LOC_198/B INVX1_LOC_15/A 0.01fF
C35441 NOR2X1_LOC_756/Y INVX1_LOC_12/Y 0.22fF
C35442 INVX1_LOC_45/A NOR2X1_LOC_158/Y 0.07fF
C35443 INVX1_LOC_5/A NOR2X1_LOC_846/A 0.01fF
C35444 NOR2X1_LOC_817/Y INVX1_LOC_57/A 0.09fF
C35445 NOR2X1_LOC_589/A INVX1_LOC_92/A 0.56fF
C35446 INVX1_LOC_245/Y NOR2X1_LOC_383/B 0.03fF
C35447 INVX1_LOC_35/A NOR2X1_LOC_15/Y 0.06fF
C35448 NOR2X1_LOC_303/Y NOR2X1_LOC_170/A 0.35fF
C35449 NAND2X1_LOC_338/B NAND2X1_LOC_489/Y 0.02fF
C35450 NOR2X1_LOC_686/B INVX1_LOC_291/A 0.05fF
C35451 NAND2X1_LOC_807/Y NAND2X1_LOC_603/a_36_24# 0.01fF
C35452 NAND2X1_LOC_208/B NAND2X1_LOC_99/A 0.02fF
C35453 INVX1_LOC_21/A NOR2X1_LOC_798/A 0.03fF
C35454 NAND2X1_LOC_783/Y INVX1_LOC_50/A 0.02fF
C35455 INVX1_LOC_255/Y NOR2X1_LOC_820/Y 0.03fF
C35456 INVX1_LOC_72/A NAND2X1_LOC_175/Y 0.10fF
C35457 INVX1_LOC_2/Y NOR2X1_LOC_188/A 0.03fF
C35458 NOR2X1_LOC_702/Y INVX1_LOC_280/A 0.08fF
C35459 INVX1_LOC_135/A NOR2X1_LOC_78/a_36_216# 0.00fF
C35460 INVX1_LOC_287/A NOR2X1_LOC_710/A 0.01fF
C35461 INVX1_LOC_166/A NAND2X1_LOC_555/Y 0.01fF
C35462 INVX1_LOC_136/A NOR2X1_LOC_278/Y 0.08fF
C35463 NOR2X1_LOC_835/B VDD 0.15fF
C35464 INVX1_LOC_256/A NAND2X1_LOC_860/A 0.02fF
C35465 INVX1_LOC_232/A INVX1_LOC_27/Y 0.08fF
C35466 NOR2X1_LOC_168/Y NAND2X1_LOC_72/B 0.01fF
C35467 NAND2X1_LOC_753/a_36_24# INVX1_LOC_11/A 0.01fF
C35468 VDD NOR2X1_LOC_167/Y 0.67fF
C35469 INVX1_LOC_303/Y VDD 0.41fF
C35470 NOR2X1_LOC_598/B NOR2X1_LOC_254/A 0.10fF
C35471 INVX1_LOC_174/A INVX1_LOC_53/A 0.86fF
C35472 INVX1_LOC_171/A INVX1_LOC_92/A 0.03fF
C35473 INVX1_LOC_299/A NOR2X1_LOC_220/B 0.03fF
C35474 NOR2X1_LOC_272/Y INVX1_LOC_48/Y 0.47fF
C35475 NOR2X1_LOC_78/A NAND2X1_LOC_469/B 0.16fF
C35476 INVX1_LOC_77/A INVX1_LOC_4/Y 6.60fF
C35477 INPUT_0 NAND2X1_LOC_96/A 0.07fF
C35478 INVX1_LOC_54/Y NOR2X1_LOC_89/A 0.05fF
C35479 INVX1_LOC_6/A NAND2X1_LOC_472/Y 0.13fF
C35480 NOR2X1_LOC_473/B NOR2X1_LOC_155/A 0.19fF
C35481 NAND2X1_LOC_363/B NOR2X1_LOC_590/A 0.07fF
C35482 NAND2X1_LOC_763/B NAND2X1_LOC_40/a_36_24# 0.00fF
C35483 INVX1_LOC_196/A NOR2X1_LOC_461/Y 0.08fF
C35484 INVX1_LOC_227/A NAND2X1_LOC_475/Y 0.10fF
C35485 INVX1_LOC_89/A NAND2X1_LOC_141/Y 0.15fF
C35486 NOR2X1_LOC_297/a_36_216# NOR2X1_LOC_38/B 0.00fF
C35487 NOR2X1_LOC_91/A INVX1_LOC_24/A 3.98fF
C35488 NAND2X1_LOC_363/B INVX1_LOC_22/Y 0.02fF
C35489 INVX1_LOC_1/Y INVX1_LOC_125/A 0.07fF
C35490 NAND2X1_LOC_392/A NAND2X1_LOC_74/B 0.11fF
C35491 NOR2X1_LOC_56/Y INVX1_LOC_76/A 0.03fF
C35492 NAND2X1_LOC_552/A NAND2X1_LOC_543/a_36_24# 0.00fF
C35493 NOR2X1_LOC_373/Y NOR2X1_LOC_662/A 0.02fF
C35494 INVX1_LOC_285/Y INVX1_LOC_9/A 0.10fF
C35495 INVX1_LOC_304/A INVX1_LOC_46/A 0.07fF
C35496 NOR2X1_LOC_537/Y INVX1_LOC_32/A 0.07fF
C35497 INVX1_LOC_22/A NOR2X1_LOC_584/Y 0.03fF
C35498 NOR2X1_LOC_186/Y NOR2X1_LOC_389/A 0.10fF
C35499 NAND2X1_LOC_338/B INVX1_LOC_32/A 0.17fF
C35500 INVX1_LOC_290/A NOR2X1_LOC_583/Y 0.01fF
C35501 NAND2X1_LOC_274/a_36_24# NAND2X1_LOC_211/Y 0.01fF
C35502 NOR2X1_LOC_344/A NOR2X1_LOC_541/B 0.00fF
C35503 VDD NOR2X1_LOC_824/Y 0.20fF
C35504 INVX1_LOC_24/A INVX1_LOC_23/A 0.84fF
C35505 INVX1_LOC_124/A INVX1_LOC_4/Y 0.01fF
C35506 NOR2X1_LOC_516/B NOR2X1_LOC_850/B 0.05fF
C35507 INVX1_LOC_220/Y INVX1_LOC_99/A 0.12fF
C35508 NOR2X1_LOC_35/Y NOR2X1_LOC_857/A 0.01fF
C35509 INVX1_LOC_64/A INVX1_LOC_217/A 0.07fF
C35510 NOR2X1_LOC_74/A INVX1_LOC_179/A 0.03fF
C35511 INVX1_LOC_278/A NAND2X1_LOC_198/B 0.01fF
C35512 INVX1_LOC_64/A NAND2X1_LOC_355/Y 0.06fF
C35513 NAND2X1_LOC_642/Y NOR2X1_LOC_98/B 0.01fF
C35514 INVX1_LOC_34/A NAND2X1_LOC_99/A 0.07fF
C35515 VDD INVX1_LOC_76/A 9.57fF
C35516 NOR2X1_LOC_278/A NOR2X1_LOC_278/Y 0.16fF
C35517 INVX1_LOC_50/A NOR2X1_LOC_716/B 0.19fF
C35518 NAND2X1_LOC_579/A NAND2X1_LOC_550/A 0.10fF
C35519 INVX1_LOC_193/Y INVX1_LOC_75/Y 0.92fF
C35520 NAND2X1_LOC_191/a_36_24# NOR2X1_LOC_205/Y 0.00fF
C35521 NOR2X1_LOC_99/B NAND2X1_LOC_207/B 0.07fF
C35522 NAND2X1_LOC_800/A INVX1_LOC_76/A 0.04fF
C35523 NOR2X1_LOC_415/a_36_216# INVX1_LOC_29/A 0.00fF
C35524 INVX1_LOC_299/A INVX1_LOC_225/Y 0.37fF
C35525 INVX1_LOC_234/A NAND2X1_LOC_254/Y 0.00fF
C35526 INVX1_LOC_279/A NAND2X1_LOC_792/B 0.01fF
C35527 INVX1_LOC_35/A NOR2X1_LOC_860/B 0.07fF
C35528 NOR2X1_LOC_516/B NOR2X1_LOC_28/a_36_216# 0.00fF
C35529 INVX1_LOC_17/A INVX1_LOC_161/Y 0.21fF
C35530 INVX1_LOC_48/A INVX1_LOC_46/Y 0.25fF
C35531 NOR2X1_LOC_134/Y INVX1_LOC_14/A 0.09fF
C35532 NAND2X1_LOC_348/A NOR2X1_LOC_673/A 0.03fF
C35533 INVX1_LOC_72/A INVX1_LOC_171/Y 0.36fF
C35534 NOR2X1_LOC_665/A INVX1_LOC_15/A 0.06fF
C35535 NOR2X1_LOC_329/B INVX1_LOC_49/Y 0.09fF
C35536 NOR2X1_LOC_137/B INVX1_LOC_9/A 0.04fF
C35537 INVX1_LOC_191/Y NOR2X1_LOC_639/Y 0.01fF
C35538 NOR2X1_LOC_468/Y INVX1_LOC_170/A 0.00fF
C35539 INVX1_LOC_64/A NAND2X1_LOC_787/B 0.07fF
C35540 INVX1_LOC_58/A INVX1_LOC_104/A 0.10fF
C35541 NOR2X1_LOC_328/Y INVX1_LOC_78/A 0.03fF
C35542 NOR2X1_LOC_540/B INVX1_LOC_274/A 0.03fF
C35543 INVX1_LOC_75/A NOR2X1_LOC_509/A 0.03fF
C35544 NOR2X1_LOC_420/Y INVX1_LOC_132/A 0.01fF
C35545 INVX1_LOC_27/A INVX1_LOC_314/Y 0.01fF
C35546 NOR2X1_LOC_848/Y INVX1_LOC_110/A 0.03fF
C35547 NOR2X1_LOC_19/B NAND2X1_LOC_254/Y 0.18fF
C35548 INVX1_LOC_89/A NOR2X1_LOC_685/Y 0.02fF
C35549 NAND2X1_LOC_803/B INVX1_LOC_30/A 0.06fF
C35550 INVX1_LOC_226/Y NOR2X1_LOC_720/A 0.01fF
C35551 INVX1_LOC_313/Y INVX1_LOC_32/A 0.07fF
C35552 NAND2X1_LOC_53/Y INVX1_LOC_142/A 0.09fF
C35553 NOR2X1_LOC_45/Y NAND2X1_LOC_199/B 0.14fF
C35554 NOR2X1_LOC_615/Y INVX1_LOC_30/A 0.02fF
C35555 INVX1_LOC_282/A INVX1_LOC_12/A 0.09fF
C35556 INVX1_LOC_304/Y INVX1_LOC_64/A 0.07fF
C35557 INVX1_LOC_35/A NAND2X1_LOC_141/A 0.06fF
C35558 INVX1_LOC_182/Y NAND2X1_LOC_792/B 0.01fF
C35559 INVX1_LOC_20/A INVX1_LOC_92/A 0.10fF
C35560 INVX1_LOC_5/A NAND2X1_LOC_116/A 0.05fF
C35561 INVX1_LOC_75/A NOR2X1_LOC_114/Y 0.04fF
C35562 NOR2X1_LOC_295/Y NOR2X1_LOC_186/Y 0.02fF
C35563 NAND2X1_LOC_35/B NOR2X1_LOC_411/A 0.26fF
C35564 NAND2X1_LOC_736/Y NAND2X1_LOC_741/Y 0.01fF
C35565 INVX1_LOC_2/A NOR2X1_LOC_489/B 0.39fF
C35566 NOR2X1_LOC_590/A INVX1_LOC_30/A 0.22fF
C35567 INVX1_LOC_58/A INVX1_LOC_263/A 0.10fF
C35568 INVX1_LOC_232/Y NOR2X1_LOC_660/Y 0.15fF
C35569 INVX1_LOC_278/A NOR2X1_LOC_401/a_36_216# 0.00fF
C35570 NAND2X1_LOC_555/Y NAND2X1_LOC_672/a_36_24# 0.01fF
C35571 INVX1_LOC_292/A NOR2X1_LOC_703/B 0.05fF
C35572 NOR2X1_LOC_71/Y NAND2X1_LOC_477/a_36_24# 0.00fF
C35573 INVX1_LOC_13/A INVX1_LOC_224/Y 0.11fF
C35574 INVX1_LOC_93/A NOR2X1_LOC_52/B 0.07fF
C35575 NOR2X1_LOC_790/B NOR2X1_LOC_614/Y 0.00fF
C35576 NOR2X1_LOC_488/Y NAND2X1_LOC_787/A 0.62fF
C35577 INVX1_LOC_35/A INVX1_LOC_226/A 0.03fF
C35578 INVX1_LOC_33/A INVX1_LOC_198/A -0.00fF
C35579 INVX1_LOC_11/A NOR2X1_LOC_303/Y 0.04fF
C35580 INVX1_LOC_272/Y NAND2X1_LOC_593/Y 0.24fF
C35581 NOR2X1_LOC_91/A NOR2X1_LOC_130/A 0.03fF
C35582 NAND2X1_LOC_499/a_36_24# INVX1_LOC_91/A 0.00fF
C35583 NAND2X1_LOC_67/Y INVX1_LOC_153/Y 0.39fF
C35584 NAND2X1_LOC_860/A NOR2X1_LOC_397/a_36_216# 0.00fF
C35585 INVX1_LOC_13/A NAND2X1_LOC_38/a_36_24# 0.00fF
C35586 NOR2X1_LOC_753/Y NAND2X1_LOC_799/A 0.02fF
C35587 NOR2X1_LOC_589/A INVX1_LOC_53/A 0.17fF
C35588 INVX1_LOC_50/A NOR2X1_LOC_717/B 0.03fF
C35589 NOR2X1_LOC_75/Y INVX1_LOC_105/A 0.00fF
C35590 D_INPUT_1 NOR2X1_LOC_757/A 0.00fF
C35591 D_INPUT_0 NOR2X1_LOC_383/B 0.00fF
C35592 NOR2X1_LOC_443/Y INVX1_LOC_135/A 0.03fF
C35593 NOR2X1_LOC_679/Y NOR2X1_LOC_152/Y 0.02fF
C35594 INVX1_LOC_24/A INVX1_LOC_31/A 0.58fF
C35595 NAND2X1_LOC_33/Y NAND2X1_LOC_725/B 0.00fF
C35596 NOR2X1_LOC_612/a_36_216# NOR2X1_LOC_652/Y 0.00fF
C35597 NOR2X1_LOC_637/B NAND2X1_LOC_350/A 0.02fF
C35598 INVX1_LOC_223/A NOR2X1_LOC_360/Y 0.10fF
C35599 NOR2X1_LOC_15/Y INVX1_LOC_257/Y 0.05fF
C35600 NOR2X1_LOC_82/A NAND2X1_LOC_276/Y 0.03fF
C35601 NOR2X1_LOC_130/A INVX1_LOC_23/A 0.13fF
C35602 INVX1_LOC_33/A INVX1_LOC_150/Y 0.07fF
C35603 INVX1_LOC_5/A INVX1_LOC_232/A 0.01fF
C35604 INVX1_LOC_90/A NAND2X1_LOC_287/a_36_24# 0.00fF
C35605 INVX1_LOC_35/A NOR2X1_LOC_97/B 0.28fF
C35606 NOR2X1_LOC_309/Y INVX1_LOC_308/Y 0.03fF
C35607 NOR2X1_LOC_151/a_36_216# INVX1_LOC_271/Y 0.01fF
C35608 NOR2X1_LOC_667/A NAND2X1_LOC_703/Y 0.09fF
C35609 INVX1_LOC_84/A INVX1_LOC_77/Y 0.07fF
C35610 NOR2X1_LOC_160/B NOR2X1_LOC_551/B 0.06fF
C35611 INVX1_LOC_91/A NOR2X1_LOC_116/a_36_216# -0.01fF
C35612 NAND2X1_LOC_740/Y INVX1_LOC_16/A 0.02fF
C35613 NOR2X1_LOC_510/B INVX1_LOC_54/A 0.15fF
C35614 NOR2X1_LOC_473/B NOR2X1_LOC_125/Y 0.01fF
C35615 INVX1_LOC_136/A NAND2X1_LOC_731/Y 0.19fF
C35616 INVX1_LOC_248/A NAND2X1_LOC_703/Y 0.02fF
C35617 INVX1_LOC_2/A INVX1_LOC_14/A 0.16fF
C35618 INVX1_LOC_14/A NOR2X1_LOC_818/Y 0.07fF
C35619 NOR2X1_LOC_92/Y NAND2X1_LOC_181/Y 0.03fF
C35620 INVX1_LOC_49/A NOR2X1_LOC_717/Y 0.06fF
C35621 INVX1_LOC_230/Y INVX1_LOC_8/A 0.07fF
C35622 NOR2X1_LOC_441/Y INVX1_LOC_155/A 0.00fF
C35623 NOR2X1_LOC_68/A NOR2X1_LOC_257/a_36_216# 0.00fF
C35624 NOR2X1_LOC_272/Y INVX1_LOC_290/A 0.08fF
C35625 NOR2X1_LOC_226/A INVX1_LOC_14/A 0.15fF
C35626 NAND2X1_LOC_287/B NAND2X1_LOC_74/B 0.07fF
C35627 INVX1_LOC_36/A INVX1_LOC_209/Y 0.03fF
C35628 INVX1_LOC_11/A INVX1_LOC_54/Y 0.00fF
C35629 INVX1_LOC_225/A NOR2X1_LOC_389/A 0.01fF
C35630 INVX1_LOC_5/A NOR2X1_LOC_366/Y 0.07fF
C35631 INVX1_LOC_180/A INVX1_LOC_18/A 0.02fF
C35632 NOR2X1_LOC_548/a_36_216# NAND2X1_LOC_72/B 0.00fF
C35633 INVX1_LOC_34/A NAND2X1_LOC_577/A 0.07fF
C35634 NOR2X1_LOC_510/Y NOR2X1_LOC_561/Y 0.03fF
C35635 INPUT_0 NAND2X1_LOC_99/A 1.24fF
C35636 NOR2X1_LOC_296/Y NAND2X1_LOC_338/B 0.16fF
C35637 INVX1_LOC_50/A NOR2X1_LOC_151/Y 0.03fF
C35638 NOR2X1_LOC_187/Y INVX1_LOC_208/A 0.00fF
C35639 NOR2X1_LOC_788/B NAND2X1_LOC_533/a_36_24# 0.02fF
C35640 NOR2X1_LOC_772/B INVX1_LOC_89/A 0.09fF
C35641 INVX1_LOC_200/A NAND2X1_LOC_850/Y 0.14fF
C35642 NOR2X1_LOC_216/Y INVX1_LOC_23/A 0.10fF
C35643 NOR2X1_LOC_71/Y INVX1_LOC_306/Y 0.10fF
C35644 NOR2X1_LOC_332/A NOR2X1_LOC_846/A 0.02fF
C35645 INPUT_3 NOR2X1_LOC_537/Y 0.09fF
C35646 NOR2X1_LOC_489/A INVX1_LOC_63/A 0.03fF
C35647 INVX1_LOC_13/Y INVX1_LOC_89/A 0.03fF
C35648 NAND2X1_LOC_308/B NOR2X1_LOC_304/Y 0.03fF
C35649 INPUT_3 NAND2X1_LOC_338/B 0.02fF
C35650 NAND2X1_LOC_324/a_36_24# NAND2X1_LOC_660/Y 0.00fF
C35651 NOR2X1_LOC_15/Y NOR2X1_LOC_188/Y 0.05fF
C35652 NOR2X1_LOC_662/A INVX1_LOC_54/A 0.20fF
C35653 VDD INVX1_LOC_127/Y 0.26fF
C35654 NAND2X1_LOC_588/a_36_24# INVX1_LOC_174/A 0.00fF
C35655 INVX1_LOC_19/Y INVX1_LOC_46/A 0.01fF
C35656 NOR2X1_LOC_690/A INVX1_LOC_61/A 0.01fF
C35657 INVX1_LOC_31/A INVX1_LOC_143/A 0.10fF
C35658 NOR2X1_LOC_188/A INVX1_LOC_29/Y 2.89fF
C35659 NAND2X1_LOC_303/Y INPUT_5 0.23fF
C35660 NOR2X1_LOC_160/B INVX1_LOC_43/A 0.03fF
C35661 INVX1_LOC_33/Y INVX1_LOC_42/A 0.03fF
C35662 NOR2X1_LOC_565/A INVX1_LOC_177/A 0.01fF
C35663 INVX1_LOC_2/A NOR2X1_LOC_717/Y 0.03fF
C35664 INVX1_LOC_45/A INVX1_LOC_236/A 0.00fF
C35665 INVX1_LOC_34/A NAND2X1_LOC_656/A 0.03fF
C35666 INVX1_LOC_286/A INVX1_LOC_57/A 0.08fF
C35667 NOR2X1_LOC_328/Y NOR2X1_LOC_503/Y 0.02fF
C35668 NAND2X1_LOC_483/Y NOR2X1_LOC_238/Y 0.00fF
C35669 NAND2X1_LOC_500/Y NAND2X1_LOC_374/Y 0.03fF
C35670 NOR2X1_LOC_777/B NOR2X1_LOC_729/A 0.03fF
C35671 NOR2X1_LOC_351/Y INVX1_LOC_272/A 0.37fF
C35672 NOR2X1_LOC_593/Y NOR2X1_LOC_303/Y 0.35fF
C35673 INVX1_LOC_21/A NAND2X1_LOC_842/B 0.03fF
C35674 INVX1_LOC_58/A INVX1_LOC_206/Y 0.39fF
C35675 NAND2X1_LOC_821/a_36_24# INVX1_LOC_53/A 0.00fF
C35676 NAND2X1_LOC_358/B NOR2X1_LOC_97/A 0.04fF
C35677 NOR2X1_LOC_843/A INVX1_LOC_77/A 0.03fF
C35678 INVX1_LOC_276/A INVX1_LOC_18/A 0.08fF
C35679 NAND2X1_LOC_740/B NAND2X1_LOC_739/a_36_24# 0.02fF
C35680 INVX1_LOC_227/A NOR2X1_LOC_457/A 0.06fF
C35681 NOR2X1_LOC_620/Y INVX1_LOC_41/A 0.01fF
C35682 INVX1_LOC_177/A NOR2X1_LOC_324/Y 0.01fF
C35683 NOR2X1_LOC_67/A INVX1_LOC_18/A 1.55fF
C35684 INVX1_LOC_33/A NAND2X1_LOC_494/a_36_24# 0.01fF
C35685 NOR2X1_LOC_456/Y INVX1_LOC_96/A 0.02fF
C35686 INVX1_LOC_24/A NOR2X1_LOC_290/Y 0.01fF
C35687 INVX1_LOC_14/A INPUT_1 0.61fF
C35688 NOR2X1_LOC_711/A INVX1_LOC_213/A 0.05fF
C35689 NOR2X1_LOC_481/A NOR2X1_LOC_295/Y 0.05fF
C35690 NOR2X1_LOC_135/Y NOR2X1_LOC_321/Y 0.11fF
C35691 INVX1_LOC_95/A INVX1_LOC_57/A 0.07fF
C35692 INVX1_LOC_1/A NOR2X1_LOC_736/Y 0.06fF
C35693 INVX1_LOC_174/A INVX1_LOC_83/A 0.47fF
C35694 INVX1_LOC_45/A INVX1_LOC_13/A 0.10fF
C35695 NOR2X1_LOC_718/Y INVX1_LOC_249/Y 0.33fF
C35696 NAND2X1_LOC_551/A NOR2X1_LOC_103/Y 0.20fF
C35697 NOR2X1_LOC_419/Y NOR2X1_LOC_720/a_36_216# 0.00fF
C35698 NAND2X1_LOC_783/A INVX1_LOC_31/A 0.02fF
C35699 INVX1_LOC_33/Y INVX1_LOC_78/A 0.03fF
C35700 NAND2X1_LOC_116/a_36_24# NOR2X1_LOC_554/B 0.00fF
C35701 NOR2X1_LOC_226/A NAND2X1_LOC_84/Y 0.18fF
C35702 NOR2X1_LOC_209/A INVX1_LOC_23/A 0.01fF
C35703 INVX1_LOC_146/Y NOR2X1_LOC_447/A 0.30fF
C35704 NOR2X1_LOC_295/Y INVX1_LOC_225/A 0.02fF
C35705 INVX1_LOC_227/A INVX1_LOC_30/A 0.10fF
C35706 NAND2X1_LOC_9/Y INVX1_LOC_304/A 0.08fF
C35707 NOR2X1_LOC_67/A INVX1_LOC_172/A 0.07fF
C35708 INVX1_LOC_5/A INVX1_LOC_186/A 0.37fF
C35709 INVX1_LOC_34/A NOR2X1_LOC_423/Y 0.04fF
C35710 NAND2X1_LOC_712/a_36_24# NOR2X1_LOC_45/B 0.00fF
C35711 INVX1_LOC_54/Y NOR2X1_LOC_593/Y 1.21fF
C35712 NAND2X1_LOC_35/B INVX1_LOC_237/Y 0.26fF
C35713 INVX1_LOC_9/A INVX1_LOC_4/Y 0.12fF
C35714 INVX1_LOC_181/Y INVX1_LOC_22/A 0.02fF
C35715 NAND2X1_LOC_574/A NOR2X1_LOC_14/a_36_216# 0.01fF
C35716 NOR2X1_LOC_763/Y INVX1_LOC_30/A 0.04fF
C35717 INVX1_LOC_233/A INVX1_LOC_304/A 0.00fF
C35718 INVX1_LOC_57/Y D_INPUT_0 0.07fF
C35719 NAND2X1_LOC_763/B NOR2X1_LOC_763/Y 0.07fF
C35720 NOR2X1_LOC_91/A NAND2X1_LOC_811/B 0.03fF
C35721 INVX1_LOC_53/A INVX1_LOC_20/A 0.06fF
C35722 INVX1_LOC_278/A NAND2X1_LOC_465/A 0.03fF
C35723 INVX1_LOC_135/A INVX1_LOC_110/A 0.00fF
C35724 INVX1_LOC_45/A NOR2X1_LOC_174/B 0.14fF
C35725 INVX1_LOC_24/A NAND2X1_LOC_859/Y 0.13fF
C35726 NOR2X1_LOC_433/a_36_216# NOR2X1_LOC_78/B 0.00fF
C35727 INVX1_LOC_4/A INVX1_LOC_92/A 0.11fF
C35728 INVX1_LOC_314/Y INVX1_LOC_137/A 0.00fF
C35729 INVX1_LOC_89/A NOR2X1_LOC_500/B 0.03fF
C35730 NAND2X1_LOC_472/Y INVX1_LOC_270/A 0.01fF
C35731 NAND2X1_LOC_67/Y INVX1_LOC_285/Y 0.07fF
C35732 INVX1_LOC_13/A INVX1_LOC_71/A 0.05fF
C35733 INVX1_LOC_34/A NOR2X1_LOC_222/Y 0.09fF
C35734 INVX1_LOC_119/A NAND2X1_LOC_534/a_36_24# 0.00fF
C35735 INVX1_LOC_279/A NOR2X1_LOC_359/Y 0.02fF
C35736 NOR2X1_LOC_455/Y VDD 0.19fF
C35737 NAND2X1_LOC_338/B INVX1_LOC_158/A 0.04fF
C35738 INVX1_LOC_94/A NOR2X1_LOC_335/a_36_216# 0.00fF
C35739 NAND2X1_LOC_454/Y NAND2X1_LOC_93/B 0.07fF
C35740 NOR2X1_LOC_411/A VDD 0.00fF
C35741 INVX1_LOC_245/Y NOR2X1_LOC_74/Y 0.01fF
C35742 NOR2X1_LOC_432/Y INVX1_LOC_266/Y 0.02fF
C35743 D_INPUT_0 NOR2X1_LOC_512/Y 0.00fF
C35744 NOR2X1_LOC_467/a_36_216# INVX1_LOC_113/Y 0.00fF
C35745 NOR2X1_LOC_401/B INVX1_LOC_168/A 0.14fF
C35746 INVX1_LOC_27/A NOR2X1_LOC_657/B 0.42fF
C35747 INVX1_LOC_30/A NOR2X1_LOC_703/A 0.05fF
C35748 INVX1_LOC_178/Y NOR2X1_LOC_662/a_36_216# 0.00fF
C35749 NOR2X1_LOC_424/a_36_216# INVX1_LOC_113/Y 0.00fF
C35750 NAND2X1_LOC_322/a_36_24# NOR2X1_LOC_374/A 0.00fF
C35751 NOR2X1_LOC_178/Y VDD 0.24fF
C35752 INVX1_LOC_177/A INVX1_LOC_179/Y 0.02fF
C35753 INVX1_LOC_41/A NAND2X1_LOC_390/A 0.31fF
C35754 NOR2X1_LOC_155/A NOR2X1_LOC_464/Y 0.01fF
C35755 NOR2X1_LOC_226/A INVX1_LOC_111/Y 0.03fF
C35756 INVX1_LOC_26/A INVX1_LOC_70/A 0.03fF
C35757 NOR2X1_LOC_246/A INVX1_LOC_71/A 0.10fF
C35758 INVX1_LOC_23/A NOR2X1_LOC_148/Y 0.00fF
C35759 NOR2X1_LOC_584/Y INVX1_LOC_261/A 0.01fF
C35760 NOR2X1_LOC_583/Y INVX1_LOC_261/Y 0.01fF
C35761 NAND2X1_LOC_549/Y NOR2X1_LOC_813/Y 0.01fF
C35762 NOR2X1_LOC_510/Y INVX1_LOC_76/A 0.37fF
C35763 NOR2X1_LOC_413/Y NAND2X1_LOC_735/B 0.55fF
C35764 INVX1_LOC_24/A NAND2X1_LOC_866/B 0.09fF
C35765 NOR2X1_LOC_434/Y VDD 0.12fF
C35766 NOR2X1_LOC_209/Y NOR2X1_LOC_220/A 0.51fF
C35767 NOR2X1_LOC_329/B INVX1_LOC_79/Y 0.01fF
C35768 NOR2X1_LOC_468/Y NAND2X1_LOC_642/Y 0.11fF
C35769 NAND2X1_LOC_149/Y NOR2X1_LOC_683/a_36_216# 0.01fF
C35770 D_INPUT_6 NAND2X1_LOC_1/Y 0.18fF
C35771 INVX1_LOC_103/A INVX1_LOC_91/A 0.07fF
C35772 INVX1_LOC_57/A INVX1_LOC_54/A 0.15fF
C35773 NOR2X1_LOC_287/A NOR2X1_LOC_168/B 0.03fF
C35774 NAND2X1_LOC_577/A INPUT_0 0.05fF
C35775 INVX1_LOC_163/A NAND2X1_LOC_659/B 0.14fF
C35776 INVX1_LOC_303/A INVX1_LOC_89/A 0.13fF
C35777 INVX1_LOC_1/Y NOR2X1_LOC_709/A 0.08fF
C35778 NAND2X1_LOC_549/Y INVX1_LOC_280/A 0.00fF
C35779 NAND2X1_LOC_390/A NAND2X1_LOC_477/A 0.03fF
C35780 INVX1_LOC_24/A NAND2X1_LOC_807/Y 0.07fF
C35781 NAND2X1_LOC_444/B INVX1_LOC_63/A 0.02fF
C35782 NOR2X1_LOC_78/B NOR2X1_LOC_131/Y 0.01fF
C35783 INVX1_LOC_217/A INVX1_LOC_282/A 0.12fF
C35784 NOR2X1_LOC_334/Y INVX1_LOC_63/A 0.07fF
C35785 NOR2X1_LOC_829/A INVX1_LOC_297/A 0.02fF
C35786 NOR2X1_LOC_641/B NOR2X1_LOC_9/Y 0.01fF
C35787 NOR2X1_LOC_554/B NOR2X1_LOC_196/Y 0.22fF
C35788 INVX1_LOC_182/Y NOR2X1_LOC_359/Y -0.00fF
C35789 NAND2X1_LOC_59/B INVX1_LOC_89/A 0.25fF
C35790 NOR2X1_LOC_92/Y NOR2X1_LOC_422/Y 0.02fF
C35791 INVX1_LOC_292/A INVX1_LOC_91/A 0.07fF
C35792 NAND2X1_LOC_662/Y NAND2X1_LOC_451/Y 0.00fF
C35793 NOR2X1_LOC_561/Y INVX1_LOC_177/A 0.01fF
C35794 INVX1_LOC_163/A VDD -0.00fF
C35795 NAND2X1_LOC_116/A NOR2X1_LOC_332/A 0.02fF
C35796 NAND2X1_LOC_852/Y NAND2X1_LOC_863/B 0.59fF
C35797 NOR2X1_LOC_751/Y NOR2X1_LOC_9/Y 0.23fF
C35798 NOR2X1_LOC_78/B NOR2X1_LOC_589/A 10.59fF
C35799 INVX1_LOC_208/A INVX1_LOC_208/Y 0.02fF
C35800 INVX1_LOC_94/Y INVX1_LOC_19/A 0.03fF
C35801 NOR2X1_LOC_361/B INVX1_LOC_76/A 0.39fF
C35802 NAND2X1_LOC_858/B NOR2X1_LOC_91/Y 0.01fF
C35803 INVX1_LOC_23/A NOR2X1_LOC_197/B 0.01fF
C35804 NAND2X1_LOC_656/A INPUT_0 0.02fF
C35805 INVX1_LOC_57/A NOR2X1_LOC_430/a_36_216# 0.02fF
C35806 INVX1_LOC_87/A INVX1_LOC_125/A 0.21fF
C35807 NOR2X1_LOC_662/A NOR2X1_LOC_438/Y 0.16fF
C35808 NAND2X1_LOC_103/a_36_24# INVX1_LOC_18/A 0.00fF
C35809 INVX1_LOC_181/Y INVX1_LOC_100/A 0.04fF
C35810 NOR2X1_LOC_255/Y INVX1_LOC_123/Y 0.07fF
C35811 NOR2X1_LOC_608/a_36_216# INVX1_LOC_7/A 0.00fF
C35812 INVX1_LOC_113/Y NOR2X1_LOC_303/a_36_216# 0.00fF
C35813 INVX1_LOC_64/A INVX1_LOC_92/A 0.21fF
C35814 INVX1_LOC_163/A NAND2X1_LOC_463/a_36_24# 0.00fF
C35815 NOR2X1_LOC_45/Y NAND2X1_LOC_469/B 0.03fF
C35816 INVX1_LOC_24/Y INVX1_LOC_117/A 0.11fF
C35817 INVX1_LOC_24/A INVX1_LOC_6/A 0.08fF
C35818 NOR2X1_LOC_30/Y INPUT_7 0.10fF
C35819 NOR2X1_LOC_220/a_36_216# INVX1_LOC_286/A 0.00fF
C35820 NOR2X1_LOC_241/A INVX1_LOC_37/A 0.01fF
C35821 INVX1_LOC_282/A NAND2X1_LOC_787/B 0.00fF
C35822 INVX1_LOC_271/A NAND2X1_LOC_432/a_36_24# 0.00fF
C35823 INVX1_LOC_67/A INVX1_LOC_79/A 0.00fF
C35824 INVX1_LOC_196/A INVX1_LOC_132/Y 0.01fF
C35825 NAND2X1_LOC_735/B NOR2X1_LOC_32/a_36_216# 0.00fF
C35826 INVX1_LOC_19/A INVX1_LOC_181/A 0.07fF
C35827 NOR2X1_LOC_743/Y NOR2X1_LOC_652/Y 0.20fF
C35828 NOR2X1_LOC_416/A NAND2X1_LOC_206/Y 0.02fF
C35829 INVX1_LOC_19/A INVX1_LOC_296/A 0.02fF
C35830 NOR2X1_LOC_218/A INVX1_LOC_12/Y 0.01fF
C35831 NOR2X1_LOC_589/A NAND2X1_LOC_392/Y 0.03fF
C35832 NOR2X1_LOC_468/Y NOR2X1_LOC_271/Y 0.03fF
C35833 NOR2X1_LOC_36/B INVX1_LOC_296/Y 0.03fF
C35834 NOR2X1_LOC_11/Y INVX1_LOC_296/A 0.16fF
C35835 NAND2X1_LOC_74/B NOR2X1_LOC_72/Y 0.00fF
C35836 INVX1_LOC_56/A NOR2X1_LOC_76/A 0.20fF
C35837 INVX1_LOC_141/Y NOR2X1_LOC_305/Y 0.27fF
C35838 NOR2X1_LOC_89/A NAND2X1_LOC_286/B 0.23fF
C35839 NAND2X1_LOC_231/Y NOR2X1_LOC_329/B 0.10fF
C35840 NAND2X1_LOC_377/Y NOR2X1_LOC_459/A 0.01fF
C35841 INVX1_LOC_23/Y INVX1_LOC_42/A 0.13fF
C35842 INVX1_LOC_304/Y INVX1_LOC_282/A 0.11fF
C35843 INVX1_LOC_14/A INVX1_LOC_118/A 0.28fF
C35844 NOR2X1_LOC_205/Y INVX1_LOC_9/A 0.04fF
C35845 INVX1_LOC_30/A NAND2X1_LOC_650/B 0.35fF
C35846 INVX1_LOC_312/Y NOR2X1_LOC_305/Y 0.14fF
C35847 INVX1_LOC_96/A NOR2X1_LOC_550/B 0.28fF
C35848 NOR2X1_LOC_263/a_36_216# INPUT_0 0.01fF
C35849 NAND2X1_LOC_807/B INVX1_LOC_57/A 0.29fF
C35850 NOR2X1_LOC_227/A NAND2X1_LOC_226/a_36_24# 0.02fF
C35851 NAND2X1_LOC_39/Y NAND2X1_LOC_16/Y 0.15fF
C35852 INVX1_LOC_243/Y NOR2X1_LOC_48/B 0.01fF
C35853 INVX1_LOC_136/A NAND2X1_LOC_287/B 0.10fF
C35854 INVX1_LOC_240/A INVX1_LOC_309/A 0.03fF
C35855 NOR2X1_LOC_604/a_36_216# INVX1_LOC_12/A 0.00fF
C35856 NOR2X1_LOC_48/B INVX1_LOC_57/A 0.15fF
C35857 NAND2X1_LOC_454/Y NAND2X1_LOC_470/B 0.36fF
C35858 INVX1_LOC_36/A NAND2X1_LOC_472/Y 0.04fF
C35859 NOR2X1_LOC_778/A INVX1_LOC_37/A 0.01fF
C35860 NAND2X1_LOC_860/A NOR2X1_LOC_89/A 0.11fF
C35861 INVX1_LOC_72/A NAND2X1_LOC_804/Y 0.03fF
C35862 NOR2X1_LOC_400/B INVX1_LOC_32/A 0.04fF
C35863 INVX1_LOC_235/Y INVX1_LOC_84/A 0.44fF
C35864 INVX1_LOC_2/A INVX1_LOC_48/A 0.10fF
C35865 NOR2X1_LOC_357/Y INVX1_LOC_71/A 0.12fF
C35866 INVX1_LOC_224/Y INVX1_LOC_32/A 0.10fF
C35867 NAND2X1_LOC_357/B NOR2X1_LOC_45/B 0.07fF
C35868 NAND2X1_LOC_149/Y INVX1_LOC_84/A 0.07fF
C35869 INVX1_LOC_57/Y NAND2X1_LOC_848/A 0.10fF
C35870 NOR2X1_LOC_68/A NAND2X1_LOC_639/A 0.04fF
C35871 GATE_865 NAND2X1_LOC_463/B 0.03fF
C35872 NOR2X1_LOC_679/Y NAND2X1_LOC_802/Y 0.08fF
C35873 NAND2X1_LOC_866/a_36_24# NOR2X1_LOC_380/Y 0.01fF
C35874 NOR2X1_LOC_274/Y VDD 0.60fF
C35875 INVX1_LOC_78/A INVX1_LOC_23/Y 0.00fF
C35876 INVX1_LOC_110/A INVX1_LOC_280/A -0.02fF
C35877 INVX1_LOC_17/A NOR2X1_LOC_841/A 0.10fF
C35878 INVX1_LOC_245/Y INVX1_LOC_179/A 0.02fF
C35879 NAND2X1_LOC_350/A NOR2X1_LOC_510/B 0.15fF
C35880 NOR2X1_LOC_68/A NOR2X1_LOC_536/A 0.03fF
C35881 NOR2X1_LOC_817/Y NOR2X1_LOC_820/Y 0.02fF
C35882 NOR2X1_LOC_387/A NAND2X1_LOC_853/Y 0.03fF
C35883 INVX1_LOC_34/A NOR2X1_LOC_69/A 0.01fF
C35884 NOR2X1_LOC_78/A NOR2X1_LOC_175/A 0.10fF
C35885 INVX1_LOC_50/Y NAND2X1_LOC_74/B 0.02fF
C35886 NAND2X1_LOC_807/Y NOR2X1_LOC_130/A 0.07fF
C35887 INVX1_LOC_240/A INVX1_LOC_11/Y 2.36fF
C35888 INVX1_LOC_203/Y VDD 0.00fF
C35889 NOR2X1_LOC_297/A NOR2X1_LOC_416/A 0.04fF
C35890 INVX1_LOC_36/A NAND2X1_LOC_637/Y 0.07fF
C35891 NOR2X1_LOC_208/Y NAND2X1_LOC_472/Y 0.01fF
C35892 INVX1_LOC_78/A NOR2X1_LOC_686/a_36_216# 0.00fF
C35893 INVX1_LOC_153/Y INVX1_LOC_76/A 0.10fF
C35894 NOR2X1_LOC_512/Y NAND2X1_LOC_848/A 0.06fF
C35895 INVX1_LOC_93/Y NOR2X1_LOC_709/A 0.10fF
C35896 INVX1_LOC_237/Y VDD 0.45fF
C35897 INVX1_LOC_101/A NOR2X1_LOC_188/A 0.02fF
C35898 INVX1_LOC_53/A INVX1_LOC_4/A 0.07fF
C35899 NOR2X1_LOC_750/Y NOR2X1_LOC_38/B 0.06fF
C35900 NAND2X1_LOC_149/Y NAND2X1_LOC_651/B 0.04fF
C35901 INVX1_LOC_208/A NOR2X1_LOC_501/B 0.03fF
C35902 NAND2X1_LOC_200/B NOR2X1_LOC_557/A 0.07fF
C35903 INVX1_LOC_71/A INVX1_LOC_66/Y 0.03fF
C35904 NOR2X1_LOC_65/B INVX1_LOC_23/Y 0.07fF
C35905 INVX1_LOC_21/A INVX1_LOC_284/A 0.03fF
C35906 INVX1_LOC_12/A NOR2X1_LOC_440/B 0.76fF
C35907 NOR2X1_LOC_499/a_36_216# NOR2X1_LOC_499/B 0.00fF
C35908 INVX1_LOC_299/A INVX1_LOC_19/A 0.27fF
C35909 NOR2X1_LOC_799/B NOR2X1_LOC_538/Y 0.15fF
C35910 NOR2X1_LOC_216/Y INVX1_LOC_313/A 0.11fF
C35911 INVX1_LOC_65/A INVX1_LOC_179/Y 0.01fF
C35912 NOR2X1_LOC_103/Y NAND2X1_LOC_489/Y 0.01fF
C35913 NOR2X1_LOC_538/B INVX1_LOC_19/A 0.00fF
C35914 INVX1_LOC_14/A NAND2X1_LOC_63/Y 0.09fF
C35915 NOR2X1_LOC_355/A NOR2X1_LOC_188/A 0.01fF
C35916 INVX1_LOC_41/A INVX1_LOC_117/A 7.43fF
C35917 INVX1_LOC_26/Y NOR2X1_LOC_621/a_36_216# 0.00fF
C35918 INVX1_LOC_2/Y NOR2X1_LOC_87/B 0.04fF
C35919 NOR2X1_LOC_68/A NAND2X1_LOC_93/B 0.07fF
C35920 NOR2X1_LOC_154/a_36_216# INVX1_LOC_37/A 0.00fF
C35921 NAND2X1_LOC_149/Y NAND2X1_LOC_220/B 0.04fF
C35922 NAND2X1_LOC_323/B NOR2X1_LOC_332/B 0.05fF
C35923 NOR2X1_LOC_78/B INVX1_LOC_20/A 0.03fF
C35924 NAND2X1_LOC_537/Y NOR2X1_LOC_89/A 0.07fF
C35925 NOR2X1_LOC_130/A INVX1_LOC_6/A 0.03fF
C35926 NOR2X1_LOC_71/Y NOR2X1_LOC_9/Y 0.01fF
C35927 INVX1_LOC_280/Y INVX1_LOC_76/A 0.03fF
C35928 NOR2X1_LOC_644/A NOR2X1_LOC_74/A 0.05fF
C35929 NOR2X1_LOC_457/B NOR2X1_LOC_155/A 0.01fF
C35930 INVX1_LOC_17/A INPUT_7 0.03fF
C35931 NOR2X1_LOC_441/Y NOR2X1_LOC_662/A 0.16fF
C35932 NAND2X1_LOC_149/Y INVX1_LOC_15/A 0.07fF
C35933 NOR2X1_LOC_454/Y D_INPUT_5 0.04fF
C35934 INVX1_LOC_28/A NOR2X1_LOC_335/B 0.02fF
C35935 NOR2X1_LOC_92/Y INVX1_LOC_3/Y 0.10fF
C35936 INVX1_LOC_24/A NAND2X1_LOC_810/B 0.02fF
C35937 NAND2X1_LOC_162/A INVX1_LOC_76/A 0.08fF
C35938 NOR2X1_LOC_329/B INPUT_0 0.03fF
C35939 NAND2X1_LOC_715/a_36_24# NOR2X1_LOC_269/Y 0.00fF
C35940 INVX1_LOC_48/A INPUT_1 0.05fF
C35941 INVX1_LOC_87/A NOR2X1_LOC_81/Y 0.04fF
C35942 INVX1_LOC_314/Y NOR2X1_LOC_216/B 0.01fF
C35943 NAND2X1_LOC_213/A NOR2X1_LOC_467/A 0.26fF
C35944 NOR2X1_LOC_318/B NOR2X1_LOC_106/A 0.25fF
C35945 NOR2X1_LOC_68/A INVX1_LOC_3/A 0.06fF
C35946 NAND2X1_LOC_199/B NOR2X1_LOC_48/Y 0.08fF
C35947 INVX1_LOC_208/Y NAND2X1_LOC_211/Y 0.06fF
C35948 INVX1_LOC_36/A NAND2X1_LOC_773/B 0.11fF
C35949 NOR2X1_LOC_68/A NOR2X1_LOC_661/A 0.06fF
C35950 INVX1_LOC_16/Y INVX1_LOC_306/Y 0.27fF
C35951 NAND2X1_LOC_714/B INVX1_LOC_273/A 0.03fF
C35952 NOR2X1_LOC_794/A NOR2X1_LOC_564/Y 0.01fF
C35953 NAND2X1_LOC_392/Y INVX1_LOC_20/A 0.43fF
C35954 NOR2X1_LOC_216/Y INVX1_LOC_6/A 1.16fF
C35955 NOR2X1_LOC_103/Y INVX1_LOC_32/A 0.17fF
C35956 INVX1_LOC_5/A INVX1_LOC_112/Y 0.02fF
C35957 NOR2X1_LOC_589/A INVX1_LOC_46/A 0.27fF
C35958 INVX1_LOC_103/A INVX1_LOC_231/A 0.00fF
C35959 INVX1_LOC_14/A NAND2X1_LOC_618/Y 0.28fF
C35960 NOR2X1_LOC_751/A NOR2X1_LOC_9/Y 0.00fF
C35961 INVX1_LOC_83/A INVX1_LOC_20/A 0.10fF
C35962 INVX1_LOC_64/A INVX1_LOC_53/A 6.28fF
C35963 INVX1_LOC_229/Y INVX1_LOC_46/A 0.78fF
C35964 NAND2X1_LOC_205/A INVX1_LOC_306/Y 0.10fF
C35965 NOR2X1_LOC_182/a_36_216# NOR2X1_LOC_155/A 0.00fF
C35966 NAND2X1_LOC_364/A NOR2X1_LOC_641/a_36_216# 0.00fF
C35967 INVX1_LOC_27/A INVX1_LOC_271/A 0.03fF
C35968 NAND2X1_LOC_45/Y VDD 0.20fF
C35969 INVX1_LOC_121/A INVX1_LOC_117/A 0.04fF
C35970 NOR2X1_LOC_272/Y INVX1_LOC_25/A 0.35fF
C35971 INVX1_LOC_256/A NAND2X1_LOC_454/Y 0.68fF
C35972 NAND2X1_LOC_84/Y NAND2X1_LOC_63/Y 0.01fF
C35973 NOR2X1_LOC_446/A INVX1_LOC_78/A 0.01fF
C35974 NOR2X1_LOC_846/Y NOR2X1_LOC_598/B 0.12fF
C35975 INVX1_LOC_229/Y NOR2X1_LOC_766/Y 0.06fF
C35976 INVX1_LOC_45/A INVX1_LOC_32/A 0.10fF
C35977 INVX1_LOC_275/Y INVX1_LOC_198/A 0.02fF
C35978 NOR2X1_LOC_360/Y INVX1_LOC_290/Y 0.12fF
C35979 NOR2X1_LOC_538/B INVX1_LOC_26/Y 0.00fF
C35980 NOR2X1_LOC_568/A INVX1_LOC_32/A 0.07fF
C35981 INVX1_LOC_1/Y NOR2X1_LOC_489/A 0.01fF
C35982 INVX1_LOC_45/A NOR2X1_LOC_623/B -0.01fF
C35983 INVX1_LOC_75/A NAND2X1_LOC_468/B 0.02fF
C35984 INVX1_LOC_104/A NAND2X1_LOC_475/Y 0.10fF
C35985 NAND2X1_LOC_807/Y NOR2X1_LOC_280/Y 0.04fF
C35986 NOR2X1_LOC_637/Y NOR2X1_LOC_584/Y 0.00fF
C35987 NOR2X1_LOC_261/Y NAND2X1_LOC_149/Y 0.19fF
C35988 INVX1_LOC_58/A NOR2X1_LOC_92/Y 0.30fF
C35989 NAND2X1_LOC_593/Y INVX1_LOC_12/A 0.00fF
C35990 NAND2X1_LOC_560/A NAND2X1_LOC_836/Y 0.01fF
C35991 INVX1_LOC_11/A NAND2X1_LOC_286/B 0.01fF
C35992 NOR2X1_LOC_860/B NAND2X1_LOC_206/B 0.08fF
C35993 INVX1_LOC_2/A NOR2X1_LOC_127/Y 0.57fF
C35994 NOR2X1_LOC_169/B INVX1_LOC_4/Y 0.02fF
C35995 NOR2X1_LOC_456/Y NOR2X1_LOC_15/Y 0.01fF
C35996 NAND2X1_LOC_796/B NAND2X1_LOC_552/A 0.00fF
C35997 NOR2X1_LOC_296/Y INVX1_LOC_224/Y 0.00fF
C35998 INVX1_LOC_16/A NOR2X1_LOC_88/Y 0.07fF
C35999 INVX1_LOC_10/A INVX1_LOC_185/A 0.01fF
C36000 NOR2X1_LOC_315/Y INVX1_LOC_19/A 0.04fF
C36001 INVX1_LOC_248/A INVX1_LOC_119/Y 0.01fF
C36002 INVX1_LOC_45/A NAND2X1_LOC_175/Y 0.41fF
C36003 NAND2X1_LOC_214/B INVX1_LOC_27/A 0.25fF
C36004 NAND2X1_LOC_837/Y INVX1_LOC_3/Y 0.08fF
C36005 NAND2X1_LOC_807/Y NAND2X1_LOC_811/B 0.12fF
C36006 INVX1_LOC_100/Y NAND2X1_LOC_642/Y 0.01fF
C36007 INVX1_LOC_21/A NOR2X1_LOC_674/Y 0.15fF
C36008 NOR2X1_LOC_311/a_36_216# NOR2X1_LOC_311/Y 0.02fF
C36009 NOR2X1_LOC_6/B NAND2X1_LOC_74/B 0.14fF
C36010 INVX1_LOC_71/A INVX1_LOC_32/A 0.10fF
C36011 NOR2X1_LOC_199/B INVX1_LOC_108/A 0.22fF
C36012 NAND2X1_LOC_350/A INVX1_LOC_57/A 0.07fF
C36013 NOR2X1_LOC_381/Y NOR2X1_LOC_660/Y 0.05fF
C36014 NAND2X1_LOC_856/A NAND2X1_LOC_175/Y 0.04fF
C36015 INVX1_LOC_55/Y NOR2X1_LOC_331/B 0.07fF
C36016 NOR2X1_LOC_68/A NAND2X1_LOC_470/B 0.03fF
C36017 INVX1_LOC_11/A NAND2X1_LOC_860/A 0.03fF
C36018 NAND2X1_LOC_784/a_36_24# NOR2X1_LOC_406/A -0.00fF
C36019 NOR2X1_LOC_91/A INVX1_LOC_286/Y 0.17fF
C36020 INVX1_LOC_285/Y INVX1_LOC_76/A 0.07fF
C36021 INVX1_LOC_77/A D_INPUT_5 0.11fF
C36022 INVX1_LOC_218/A INVX1_LOC_63/A 0.03fF
C36023 INVX1_LOC_16/A INVX1_LOC_84/A 0.31fF
C36024 NOR2X1_LOC_441/Y INVX1_LOC_57/A 0.03fF
C36025 INVX1_LOC_89/A NOR2X1_LOC_99/Y 0.15fF
C36026 INVX1_LOC_1/Y INVX1_LOC_294/A 0.05fF
C36027 INPUT_0 NOR2X1_LOC_107/a_36_216# 0.00fF
C36028 NAND2X1_LOC_364/A INVX1_LOC_116/Y 0.02fF
C36029 INVX1_LOC_41/A INVX1_LOC_3/Y 0.01fF
C36030 NAND2X1_LOC_463/B INVX1_LOC_166/Y 0.15fF
C36031 NOR2X1_LOC_623/a_36_216# INVX1_LOC_15/A 0.01fF
C36032 NAND2X1_LOC_374/Y NAND2X1_LOC_499/a_36_24# 0.00fF
C36033 INVX1_LOC_201/Y INVX1_LOC_3/Y 0.05fF
C36034 INVX1_LOC_72/Y NAND2X1_LOC_99/A 0.01fF
C36035 NOR2X1_LOC_272/Y INVX1_LOC_1/A 0.40fF
C36036 NAND2X1_LOC_642/Y NAND2X1_LOC_655/B 0.09fF
C36037 NOR2X1_LOC_311/Y INVX1_LOC_20/A 0.18fF
C36038 INVX1_LOC_39/A INVX1_LOC_14/A 0.14fF
C36039 INVX1_LOC_160/A NOR2X1_LOC_857/A 0.10fF
C36040 NOR2X1_LOC_180/B NOR2X1_LOC_155/A 0.01fF
C36041 INVX1_LOC_22/A NAND2X1_LOC_500/B 0.01fF
C36042 INVX1_LOC_217/Y NAND2X1_LOC_618/Y 0.01fF
C36043 NOR2X1_LOC_738/A NOR2X1_LOC_155/A 0.08fF
C36044 NAND2X1_LOC_181/Y INVX1_LOC_168/Y 0.01fF
C36045 NOR2X1_LOC_398/Y INVX1_LOC_3/Y 0.03fF
C36046 NAND2X1_LOC_213/A INVX1_LOC_1/A 0.07fF
C36047 NAND2X1_LOC_222/B NAND2X1_LOC_473/A 0.02fF
C36048 INVX1_LOC_28/A NOR2X1_LOC_88/Y 7.28fF
C36049 INVX1_LOC_30/Y NAND2X1_LOC_74/B 0.02fF
C36050 INVX1_LOC_88/Y INVX1_LOC_271/Y 0.05fF
C36051 NAND2X1_LOC_711/B NAND2X1_LOC_787/Y 0.04fF
C36052 D_INPUT_1 NAND2X1_LOC_198/B 0.34fF
C36053 NOR2X1_LOC_152/Y NOR2X1_LOC_686/a_36_216# 0.01fF
C36054 INVX1_LOC_31/A INVX1_LOC_38/Y 0.26fF
C36055 NAND2X1_LOC_67/Y NOR2X1_LOC_205/Y 0.00fF
C36056 INVX1_LOC_73/A NOR2X1_LOC_155/A 0.00fF
C36057 INVX1_LOC_232/A INVX1_LOC_42/A 0.44fF
C36058 INVX1_LOC_290/A INVX1_LOC_109/Y 0.10fF
C36059 NOR2X1_LOC_299/Y INVX1_LOC_163/Y 0.01fF
C36060 NAND2X1_LOC_11/Y NOR2X1_LOC_467/A 0.05fF
C36061 NAND2X1_LOC_361/Y NOR2X1_LOC_621/A 0.18fF
C36062 INVX1_LOC_66/A INVX1_LOC_19/A 0.02fF
C36063 INVX1_LOC_58/A NAND2X1_LOC_837/Y 1.26fF
C36064 NOR2X1_LOC_82/A NOR2X1_LOC_140/A 0.07fF
C36065 INVX1_LOC_49/A NOR2X1_LOC_383/B 4.36fF
C36066 NOR2X1_LOC_521/Y INVX1_LOC_284/A 0.00fF
C36067 NOR2X1_LOC_78/B INVX1_LOC_4/A 0.17fF
C36068 INVX1_LOC_90/A NOR2X1_LOC_257/Y 0.03fF
C36069 INVX1_LOC_20/A INVX1_LOC_46/A 2.11fF
C36070 INVX1_LOC_28/A INVX1_LOC_84/A 0.25fF
C36071 INVX1_LOC_162/Y INVX1_LOC_26/A 0.02fF
C36072 NOR2X1_LOC_709/A INVX1_LOC_87/A 0.03fF
C36073 INVX1_LOC_75/A NAND2X1_LOC_141/Y 0.22fF
C36074 NOR2X1_LOC_216/Y NOR2X1_LOC_117/Y 0.05fF
C36075 NOR2X1_LOC_383/Y INVX1_LOC_42/A 0.01fF
C36076 INVX1_LOC_103/A NOR2X1_LOC_592/A -0.01fF
C36077 NOR2X1_LOC_557/Y INVX1_LOC_270/A 0.21fF
C36078 INVX1_LOC_143/A NOR2X1_LOC_80/Y 0.32fF
C36079 INVX1_LOC_223/Y NOR2X1_LOC_500/B 0.00fF
C36080 NOR2X1_LOC_511/a_36_216# INVX1_LOC_78/A 0.00fF
C36081 NOR2X1_LOC_91/A INVX1_LOC_185/Y 0.01fF
C36082 NOR2X1_LOC_848/Y NOR2X1_LOC_195/A 0.06fF
C36083 INVX1_LOC_16/A INVX1_LOC_15/A 0.06fF
C36084 INVX1_LOC_233/A NAND2X1_LOC_169/a_36_24# 0.00fF
C36085 NOR2X1_LOC_527/a_36_216# INVX1_LOC_285/A 0.00fF
C36086 INVX1_LOC_64/A INVX1_LOC_184/A 0.04fF
C36087 INVX1_LOC_58/A INVX1_LOC_41/A 0.03fF
C36088 INVX1_LOC_21/A INVX1_LOC_72/A 0.10fF
C36089 NAND2X1_LOC_79/a_36_24# NOR2X1_LOC_392/Y 0.00fF
C36090 INVX1_LOC_20/A NOR2X1_LOC_766/Y 0.51fF
C36091 NOR2X1_LOC_554/B NOR2X1_LOC_846/A 0.01fF
C36092 INVX1_LOC_310/A INVX1_LOC_26/Y 0.01fF
C36093 NAND2X1_LOC_198/B NOR2X1_LOC_652/Y 0.10fF
C36094 NOR2X1_LOC_672/Y NOR2X1_LOC_392/Y 0.02fF
C36095 INVX1_LOC_93/Y NOR2X1_LOC_489/A 0.04fF
C36096 INVX1_LOC_46/A NOR2X1_LOC_765/Y 0.03fF
C36097 NOR2X1_LOC_160/B NOR2X1_LOC_218/A 0.02fF
C36098 INVX1_LOC_21/A INVX1_LOC_198/Y 0.01fF
C36099 INVX1_LOC_2/A NOR2X1_LOC_383/B 0.12fF
C36100 INVX1_LOC_35/A INVX1_LOC_34/A 0.13fF
C36101 INVX1_LOC_266/A INVX1_LOC_136/A 0.37fF
C36102 NOR2X1_LOC_52/B NOR2X1_LOC_15/a_36_216# 0.01fF
C36103 NOR2X1_LOC_809/a_36_216# NOR2X1_LOC_334/Y 0.02fF
C36104 NAND2X1_LOC_182/A NAND2X1_LOC_787/A 0.01fF
C36105 NAND2X1_LOC_860/A NOR2X1_LOC_52/B 0.05fF
C36106 NOR2X1_LOC_123/B INVX1_LOC_32/A 0.10fF
C36107 NOR2X1_LOC_226/A NOR2X1_LOC_383/B 0.07fF
C36108 INVX1_LOC_58/A NOR2X1_LOC_207/A 0.02fF
C36109 NOR2X1_LOC_91/A NOR2X1_LOC_265/a_36_216# 0.00fF
C36110 INVX1_LOC_7/A INVX1_LOC_4/Y 0.03fF
C36111 INVX1_LOC_83/A INVX1_LOC_4/A 0.10fF
C36112 INVX1_LOC_1/A NAND2X1_LOC_364/A 0.18fF
C36113 NOR2X1_LOC_655/B INVX1_LOC_57/A 0.05fF
C36114 INVX1_LOC_249/A INVX1_LOC_27/A 0.03fF
C36115 NOR2X1_LOC_765/Y NOR2X1_LOC_766/Y 0.02fF
C36116 NOR2X1_LOC_6/B NOR2X1_LOC_660/Y 0.09fF
C36117 NOR2X1_LOC_802/A INVX1_LOC_58/Y 0.02fF
C36118 INVX1_LOC_14/A INVX1_LOC_61/A 0.07fF
C36119 NOR2X1_LOC_455/Y INVX1_LOC_177/A 0.02fF
C36120 INVX1_LOC_157/A NAND2X1_LOC_454/Y 0.04fF
C36121 NOR2X1_LOC_65/B INVX1_LOC_232/A 0.10fF
C36122 INVX1_LOC_230/Y NOR2X1_LOC_414/a_36_216# 0.00fF
C36123 NOR2X1_LOC_160/B NAND2X1_LOC_510/A 0.02fF
C36124 NOR2X1_LOC_423/a_36_216# INVX1_LOC_96/Y 0.00fF
C36125 INVX1_LOC_286/Y INVX1_LOC_31/A 0.07fF
C36126 INVX1_LOC_28/A INVX1_LOC_15/A 0.14fF
C36127 INVX1_LOC_256/A NOR2X1_LOC_68/A 0.07fF
C36128 INVX1_LOC_35/A NAND2X1_LOC_231/Y 0.12fF
C36129 INVX1_LOC_57/Y NOR2X1_LOC_134/Y 0.03fF
C36130 NOR2X1_LOC_819/a_36_216# INPUT_3 0.00fF
C36131 INVX1_LOC_102/Y INVX1_LOC_32/A 0.10fF
C36132 D_INPUT_1 INVX1_LOC_53/Y 0.03fF
C36133 INVX1_LOC_200/A INVX1_LOC_41/Y 0.71fF
C36134 INVX1_LOC_64/A NOR2X1_LOC_78/B 2.46fF
C36135 INVX1_LOC_20/Y NAND2X1_LOC_223/A 0.03fF
C36136 INVX1_LOC_101/Y NOR2X1_LOC_577/Y 0.00fF
C36137 NOR2X1_LOC_690/A NAND2X1_LOC_705/Y 0.02fF
C36138 NOR2X1_LOC_355/B INVX1_LOC_29/A 0.05fF
C36139 NOR2X1_LOC_690/Y NAND2X1_LOC_787/Y 0.02fF
C36140 NOR2X1_LOC_296/Y INVX1_LOC_71/A 0.41fF
C36141 NAND2X1_LOC_430/a_36_24# NAND2X1_LOC_639/A 0.01fF
C36142 NAND2X1_LOC_358/Y INVX1_LOC_57/A 0.07fF
C36143 INVX1_LOC_99/Y NOR2X1_LOC_778/B 0.01fF
C36144 D_INPUT_1 NOR2X1_LOC_665/A 0.08fF
C36145 INVX1_LOC_90/A NOR2X1_LOC_301/A 0.03fF
C36146 INVX1_LOC_10/A INVX1_LOC_270/Y 0.89fF
C36147 INVX1_LOC_230/Y NAND2X1_LOC_79/Y 0.02fF
C36148 INVX1_LOC_136/A NOR2X1_LOC_248/Y 0.01fF
C36149 NAND2X1_LOC_564/B NAND2X1_LOC_793/B -0.09fF
C36150 NOR2X1_LOC_666/Y NOR2X1_LOC_142/Y 0.01fF
C36151 INVX1_LOC_21/A NOR2X1_LOC_537/Y 0.07fF
C36152 NOR2X1_LOC_760/a_36_216# NOR2X1_LOC_577/Y 0.01fF
C36153 INPUT_0 NOR2X1_LOC_620/a_36_216# 0.00fF
C36154 INVX1_LOC_21/A NAND2X1_LOC_338/B 0.07fF
C36155 NOR2X1_LOC_124/A NAND2X1_LOC_74/B 0.02fF
C36156 NOR2X1_LOC_215/a_36_216# INVX1_LOC_63/Y 0.01fF
C36157 NOR2X1_LOC_474/A NOR2X1_LOC_573/Y 0.16fF
C36158 INVX1_LOC_166/A NAND2X1_LOC_624/A 0.04fF
C36159 NOR2X1_LOC_269/Y INVX1_LOC_290/Y 0.00fF
C36160 NAND2X1_LOC_537/Y NOR2X1_LOC_52/B 0.39fF
C36161 INPUT_1 NOR2X1_LOC_383/B 0.01fF
C36162 INVX1_LOC_17/A NOR2X1_LOC_392/B 0.03fF
C36163 INVX1_LOC_21/A NAND2X1_LOC_323/B 0.06fF
C36164 NAND2X1_LOC_796/B NOR2X1_LOC_773/Y -0.08fF
C36165 INVX1_LOC_13/Y INVX1_LOC_25/Y 0.14fF
C36166 INVX1_LOC_36/A INVX1_LOC_24/A 5.76fF
C36167 INVX1_LOC_2/Y NAND2X1_LOC_219/B 0.19fF
C36168 INVX1_LOC_53/Y NOR2X1_LOC_652/Y 0.65fF
C36169 NOR2X1_LOC_627/Y INVX1_LOC_1/A 0.00fF
C36170 NOR2X1_LOC_457/A INVX1_LOC_104/A 0.07fF
C36171 NOR2X1_LOC_45/Y INVX1_LOC_63/Y 0.03fF
C36172 INVX1_LOC_239/A NOR2X1_LOC_399/Y 0.03fF
C36173 INVX1_LOC_181/Y INVX1_LOC_18/A 0.03fF
C36174 NAND2X1_LOC_472/Y INVX1_LOC_63/A 0.07fF
C36175 INVX1_LOC_217/A INVX1_LOC_41/Y 0.07fF
C36176 D_INPUT_1 NOR2X1_LOC_76/a_36_216# 0.00fF
C36177 NOR2X1_LOC_68/A NOR2X1_LOC_781/Y 0.05fF
C36178 INVX1_LOC_64/A INVX1_LOC_83/A 11.93fF
C36179 NAND2X1_LOC_11/Y INVX1_LOC_1/A 0.03fF
C36180 INVX1_LOC_55/Y NOR2X1_LOC_493/A 0.03fF
C36181 NAND2X1_LOC_783/A NOR2X1_LOC_109/Y 0.10fF
C36182 NOR2X1_LOC_670/Y INVX1_LOC_284/A 0.16fF
C36183 NOR2X1_LOC_671/Y INVX1_LOC_20/A 0.01fF
C36184 INVX1_LOC_38/A NOR2X1_LOC_450/B 0.02fF
C36185 NAND2X1_LOC_719/a_36_24# INVX1_LOC_96/Y 0.00fF
C36186 INVX1_LOC_27/A INVX1_LOC_137/A 0.01fF
C36187 NOR2X1_LOC_82/A NOR2X1_LOC_709/A 0.12fF
C36188 NOR2X1_LOC_598/B NOR2X1_LOC_180/B 0.26fF
C36189 NAND2X1_LOC_705/Y NAND2X1_LOC_717/a_36_24# 0.01fF
C36190 NOR2X1_LOC_617/Y INVX1_LOC_217/A 0.57fF
C36191 NOR2X1_LOC_130/A NOR2X1_LOC_109/Y 0.07fF
C36192 INVX1_LOC_215/Y NAND2X1_LOC_477/A 0.24fF
C36193 NOR2X1_LOC_551/a_36_216# NOR2X1_LOC_383/B 0.00fF
C36194 NAND2X1_LOC_642/Y INVX1_LOC_251/A 0.01fF
C36195 INVX1_LOC_31/A NOR2X1_LOC_4/a_36_216# 0.01fF
C36196 INVX1_LOC_78/Y INVX1_LOC_271/Y 0.03fF
C36197 INVX1_LOC_17/A NAND2X1_LOC_294/a_36_24# 0.00fF
C36198 NAND2X1_LOC_96/A INVX1_LOC_19/A 0.07fF
C36199 NOR2X1_LOC_598/B NOR2X1_LOC_738/A 0.15fF
C36200 INVX1_LOC_36/A NOR2X1_LOC_557/Y 0.18fF
C36201 INVX1_LOC_77/A NOR2X1_LOC_360/Y 0.08fF
C36202 INVX1_LOC_38/A NOR2X1_LOC_257/Y 0.00fF
C36203 NOR2X1_LOC_208/Y INVX1_LOC_24/A 0.03fF
C36204 NOR2X1_LOC_61/A NOR2X1_LOC_865/Y 0.02fF
C36205 INVX1_LOC_97/Y NOR2X1_LOC_180/B -0.01fF
C36206 NAND2X1_LOC_725/B INVX1_LOC_22/A 0.06fF
C36207 INVX1_LOC_278/A INVX1_LOC_28/A 0.07fF
C36208 INVX1_LOC_163/A NAND2X1_LOC_376/a_36_24# 0.00fF
C36209 INVX1_LOC_88/A INVX1_LOC_25/Y 0.01fF
C36210 NAND2X1_LOC_27/a_36_24# INVX1_LOC_83/A 0.00fF
C36211 NOR2X1_LOC_61/A NOR2X1_LOC_243/B 0.05fF
C36212 NAND2X1_LOC_182/A INVX1_LOC_30/A 0.03fF
C36213 NOR2X1_LOC_643/Y NAND2X1_LOC_656/A 0.04fF
C36214 NOR2X1_LOC_237/Y INVX1_LOC_24/A 0.00fF
C36215 INVX1_LOC_30/A INVX1_LOC_104/A 0.31fF
C36216 NOR2X1_LOC_798/A INVX1_LOC_171/A 0.03fF
C36217 NOR2X1_LOC_78/B INVX1_LOC_43/Y 0.06fF
C36218 NOR2X1_LOC_35/Y INVX1_LOC_15/A 0.47fF
C36219 NOR2X1_LOC_148/Y INVX1_LOC_301/A 0.00fF
C36220 INVX1_LOC_208/A NOR2X1_LOC_218/A 0.02fF
C36221 INVX1_LOC_35/A INVX1_LOC_131/A 0.22fF
C36222 INVX1_LOC_58/A NAND2X1_LOC_662/B 0.13fF
C36223 NOR2X1_LOC_225/a_36_216# NOR2X1_LOC_773/Y 0.00fF
C36224 INVX1_LOC_70/Y NOR2X1_LOC_278/Y 0.11fF
C36225 INVX1_LOC_161/Y NOR2X1_LOC_321/a_36_216# 0.01fF
C36226 D_INPUT_1 NOR2X1_LOC_113/B 0.03fF
C36227 INVX1_LOC_254/Y NOR2X1_LOC_350/A 0.20fF
C36228 NAND2X1_LOC_564/B NOR2X1_LOC_103/Y 0.00fF
C36229 NAND2X1_LOC_116/A NOR2X1_LOC_554/B 0.00fF
C36230 NAND2X1_LOC_214/B NOR2X1_LOC_19/B 0.02fF
C36231 INVX1_LOC_21/A INVX1_LOC_313/Y 0.08fF
C36232 INVX1_LOC_2/A INVX1_LOC_57/Y 0.07fF
C36233 NOR2X1_LOC_604/Y INVX1_LOC_311/A 0.11fF
C36234 INVX1_LOC_76/A INVX1_LOC_4/Y 0.10fF
C36235 INVX1_LOC_46/A INVX1_LOC_4/A 0.44fF
C36236 INVX1_LOC_36/A INVX1_LOC_143/A 0.03fF
C36237 INVX1_LOC_35/A INPUT_0 7.57fF
C36238 INVX1_LOC_47/Y NAND2X1_LOC_262/a_36_24# 0.01fF
C36239 INVX1_LOC_124/A NOR2X1_LOC_360/Y 0.16fF
C36240 INVX1_LOC_89/A INVX1_LOC_198/A 0.00fF
C36241 INVX1_LOC_57/Y NOR2X1_LOC_226/A 0.10fF
C36242 NOR2X1_LOC_337/Y INVX1_LOC_23/A 0.02fF
C36243 INVX1_LOC_13/A NOR2X1_LOC_647/a_36_216# 0.02fF
C36244 NOR2X1_LOC_722/a_36_216# INVX1_LOC_113/Y 0.00fF
C36245 INVX1_LOC_27/A NOR2X1_LOC_19/B 0.92fF
C36246 NOR2X1_LOC_667/A INVX1_LOC_72/A 0.04fF
C36247 INVX1_LOC_304/Y INVX1_LOC_41/Y 0.01fF
C36248 INVX1_LOC_13/Y INVX1_LOC_75/A 0.07fF
C36249 INVX1_LOC_12/A INVX1_LOC_185/A 0.03fF
C36250 INVX1_LOC_292/A NOR2X1_LOC_553/B 0.01fF
C36251 NOR2X1_LOC_577/Y NOR2X1_LOC_578/a_36_216# 0.02fF
C36252 NOR2X1_LOC_91/A NOR2X1_LOC_56/Y 0.02fF
C36253 NOR2X1_LOC_273/Y INVX1_LOC_96/Y 0.00fF
C36254 NOR2X1_LOC_689/Y NAND2X1_LOC_729/B 0.03fF
C36255 NOR2X1_LOC_471/Y NOR2X1_LOC_478/a_36_216# 0.00fF
C36256 NOR2X1_LOC_89/A NOR2X1_LOC_487/Y 0.04fF
C36257 INVX1_LOC_103/A NOR2X1_LOC_510/a_36_216# 0.01fF
C36258 INVX1_LOC_268/A NOR2X1_LOC_658/Y 0.03fF
C36259 INVX1_LOC_150/Y INVX1_LOC_150/A 0.04fF
C36260 INVX1_LOC_181/Y NOR2X1_LOC_709/a_36_216# 0.00fF
C36261 INVX1_LOC_251/A NOR2X1_LOC_271/Y 0.07fF
C36262 NOR2X1_LOC_331/B INVX1_LOC_32/A 0.30fF
C36263 INVX1_LOC_25/A NOR2X1_LOC_405/A 0.18fF
C36264 INVX1_LOC_17/A INVX1_LOC_90/A 0.28fF
C36265 NAND2X1_LOC_206/Y INVX1_LOC_63/A 0.07fF
C36266 NOR2X1_LOC_354/B NOR2X1_LOC_325/A 0.02fF
C36267 NOR2X1_LOC_309/Y NOR2X1_LOC_557/Y 0.14fF
C36268 NOR2X1_LOC_500/A NOR2X1_LOC_778/B 0.03fF
C36269 INVX1_LOC_17/A NOR2X1_LOC_389/B 0.54fF
C36270 NOR2X1_LOC_27/Y INVX1_LOC_207/A 0.02fF
C36271 NOR2X1_LOC_181/Y NOR2X1_LOC_254/Y 0.09fF
C36272 NOR2X1_LOC_511/a_36_216# NOR2X1_LOC_152/Y 0.01fF
C36273 NOR2X1_LOC_56/Y INVX1_LOC_23/A 0.07fF
C36274 NOR2X1_LOC_91/A VDD 2.59fF
C36275 INVX1_LOC_286/A INVX1_LOC_306/Y 0.11fF
C36276 VDD NOR2X1_LOC_668/Y 0.24fF
C36277 INVX1_LOC_136/A INVX1_LOC_30/Y 0.03fF
C36278 NAND2X1_LOC_659/B INVX1_LOC_23/A 0.02fF
C36279 INVX1_LOC_77/A NAND2X1_LOC_451/Y 0.10fF
C36280 NAND2X1_LOC_734/B NAND2X1_LOC_734/a_36_24# 0.00fF
C36281 NOR2X1_LOC_384/Y NOR2X1_LOC_86/A 0.24fF
C36282 NOR2X1_LOC_471/Y INVX1_LOC_90/A 0.00fF
C36283 INVX1_LOC_63/A NAND2X1_LOC_773/B 0.07fF
C36284 NOR2X1_LOC_91/A NAND2X1_LOC_800/A 0.03fF
C36285 NAND2X1_LOC_364/Y INVX1_LOC_196/A 0.03fF
C36286 INVX1_LOC_35/Y NAND2X1_LOC_254/Y 0.24fF
C36287 NAND2X1_LOC_35/Y NAND2X1_LOC_623/B 0.13fF
C36288 INVX1_LOC_39/A INVX1_LOC_48/A 0.02fF
C36289 INVX1_LOC_36/A NAND2X1_LOC_783/A 0.14fF
C36290 INVX1_LOC_88/A INVX1_LOC_75/A 0.14fF
C36291 INVX1_LOC_38/A NOR2X1_LOC_30/Y 0.04fF
C36292 NAND2X1_LOC_725/A NAND2X1_LOC_729/B 0.20fF
C36293 INVX1_LOC_36/A NOR2X1_LOC_525/a_36_216# 0.02fF
C36294 INVX1_LOC_5/A NOR2X1_LOC_78/A 0.08fF
C36295 NAND2X1_LOC_555/Y INVX1_LOC_90/A 0.07fF
C36296 INVX1_LOC_298/Y INVX1_LOC_281/Y 0.09fF
C36297 NAND2X1_LOC_96/A INVX1_LOC_26/Y 0.07fF
C36298 INVX1_LOC_146/Y INVX1_LOC_23/A 0.05fF
C36299 NAND2X1_LOC_30/Y NOR2X1_LOC_163/Y 0.03fF
C36300 INVX1_LOC_36/A NOR2X1_LOC_130/A 0.08fF
C36301 INVX1_LOC_230/Y NOR2X1_LOC_750/A 0.03fF
C36302 INVX1_LOC_17/A NAND2X1_LOC_348/A 0.06fF
C36303 INVX1_LOC_64/A NOR2X1_LOC_164/Y 0.00fF
C36304 INVX1_LOC_108/Y NOR2X1_LOC_35/Y 0.25fF
C36305 NOR2X1_LOC_658/Y NOR2X1_LOC_367/a_36_216# 0.01fF
C36306 NAND2X1_LOC_564/B INVX1_LOC_71/A 0.07fF
C36307 NAND2X1_LOC_9/Y INVX1_LOC_20/A 0.09fF
C36308 VDD INVX1_LOC_23/A 1.59fF
C36309 NOR2X1_LOC_680/a_36_216# INVX1_LOC_271/Y 0.01fF
C36310 INVX1_LOC_32/A NOR2X1_LOC_592/B 0.09fF
C36311 NOR2X1_LOC_474/A INVX1_LOC_172/Y 0.00fF
C36312 NOR2X1_LOC_778/B NOR2X1_LOC_254/Y 0.01fF
C36313 NOR2X1_LOC_434/Y INVX1_LOC_65/A 0.00fF
C36314 NOR2X1_LOC_843/A INVX1_LOC_179/Y 0.00fF
C36315 NOR2X1_LOC_489/A INVX1_LOC_87/A 0.30fF
C36316 INVX1_LOC_233/A INVX1_LOC_20/A 0.37fF
C36317 INVX1_LOC_230/Y NOR2X1_LOC_750/a_36_216# 0.00fF
C36318 NOR2X1_LOC_423/Y INVX1_LOC_266/Y 0.09fF
C36319 NAND2X1_LOC_784/A NOR2X1_LOC_111/A 0.20fF
C36320 INVX1_LOC_95/A INVX1_LOC_306/Y 0.01fF
C36321 INVX1_LOC_286/Y NAND2X1_LOC_807/Y 0.10fF
C36322 INVX1_LOC_27/A NAND2X1_LOC_813/a_36_24# 0.00fF
C36323 NAND2X1_LOC_1/Y NAND2X1_LOC_31/a_36_24# 0.01fF
C36324 INVX1_LOC_208/A INVX1_LOC_155/Y 0.07fF
C36325 NOR2X1_LOC_816/A NAND2X1_LOC_840/Y 0.01fF
C36326 INVX1_LOC_208/Y INVX1_LOC_155/A 0.22fF
C36327 INVX1_LOC_57/Y INPUT_1 0.09fF
C36328 NAND2X1_LOC_574/A INVX1_LOC_3/Y 0.03fF
C36329 NAND2X1_LOC_514/Y NOR2X1_LOC_106/A 0.00fF
C36330 INVX1_LOC_37/A NOR2X1_LOC_678/A 0.03fF
C36331 INVX1_LOC_64/A INVX1_LOC_46/A 0.17fF
C36332 INVX1_LOC_280/A NOR2X1_LOC_646/B 0.07fF
C36333 NOR2X1_LOC_576/B INVX1_LOC_300/Y 0.06fF
C36334 INVX1_LOC_229/Y NAND2X1_LOC_866/A 0.78fF
C36335 INVX1_LOC_26/A NAND2X1_LOC_62/a_36_24# 0.01fF
C36336 NOR2X1_LOC_23/a_36_216# INVX1_LOC_3/Y 0.01fF
C36337 NOR2X1_LOC_222/Y INVX1_LOC_266/Y 0.07fF
C36338 GATE_811 NAND2X1_LOC_863/B 0.27fF
C36339 NOR2X1_LOC_457/A INVX1_LOC_206/Y 0.10fF
C36340 INVX1_LOC_17/A NAND2X1_LOC_123/a_36_24# 0.00fF
C36341 NOR2X1_LOC_318/A NOR2X1_LOC_743/Y 0.07fF
C36342 INVX1_LOC_94/Y NOR2X1_LOC_841/A 0.01fF
C36343 INVX1_LOC_259/Y NOR2X1_LOC_684/Y 0.04fF
C36344 NOR2X1_LOC_237/Y NOR2X1_LOC_130/A 0.07fF
C36345 INVX1_LOC_1/A NOR2X1_LOC_405/A 0.04fF
C36346 NAND2X1_LOC_721/B NOR2X1_LOC_322/Y 0.24fF
C36347 NAND2X1_LOC_858/B INVX1_LOC_141/Y 0.02fF
C36348 NOR2X1_LOC_459/B NOR2X1_LOC_459/A 0.15fF
C36349 NOR2X1_LOC_140/A INVX1_LOC_59/Y 0.01fF
C36350 NAND2X1_LOC_51/B INVX1_LOC_72/A 0.10fF
C36351 NAND2X1_LOC_703/Y INVX1_LOC_20/A 0.01fF
C36352 NAND2X1_LOC_858/B INVX1_LOC_312/Y 0.06fF
C36353 NOR2X1_LOC_813/Y NOR2X1_LOC_293/a_36_216# 0.01fF
C36354 NOR2X1_LOC_443/Y NOR2X1_LOC_862/B 0.09fF
C36355 NOR2X1_LOC_457/A NOR2X1_LOC_600/Y 0.00fF
C36356 NAND2X1_LOC_724/a_36_24# NOR2X1_LOC_773/Y 0.01fF
C36357 INVX1_LOC_87/A INVX1_LOC_294/A 0.13fF
C36358 NOR2X1_LOC_278/Y INVX1_LOC_285/A 0.07fF
C36359 NOR2X1_LOC_175/B NOR2X1_LOC_175/a_36_216# 0.01fF
C36360 INVX1_LOC_159/A NAND2X1_LOC_653/a_36_24# 0.00fF
C36361 INVX1_LOC_33/A NOR2X1_LOC_72/a_36_216# 0.00fF
C36362 NOR2X1_LOC_38/B NAND2X1_LOC_82/Y 0.25fF
C36363 INVX1_LOC_109/A INVX1_LOC_15/A 0.01fF
C36364 INVX1_LOC_129/A INVX1_LOC_92/A 0.10fF
C36365 NAND2X1_LOC_227/Y INVX1_LOC_187/A 0.06fF
C36366 NOR2X1_LOC_770/B INVX1_LOC_89/A 0.01fF
C36367 NAND2X1_LOC_364/A NOR2X1_LOC_188/A 0.13fF
C36368 NOR2X1_LOC_309/Y NOR2X1_LOC_130/A 0.07fF
C36369 INVX1_LOC_1/A NOR2X1_LOC_857/A 0.07fF
C36370 NAND2X1_LOC_364/A NOR2X1_LOC_548/B 0.10fF
C36371 NOR2X1_LOC_205/Y INVX1_LOC_76/A 0.01fF
C36372 INVX1_LOC_77/A NOR2X1_LOC_567/B 0.09fF
C36373 INVX1_LOC_306/A NOR2X1_LOC_709/A 0.31fF
C36374 INVX1_LOC_55/Y NOR2X1_LOC_388/Y 0.01fF
C36375 NOR2X1_LOC_175/a_36_216# INVX1_LOC_22/A 0.01fF
C36376 NOR2X1_LOC_392/Y NOR2X1_LOC_99/Y 0.01fF
C36377 INVX1_LOC_14/A D_INPUT_3 0.62fF
C36378 NOR2X1_LOC_68/A INVX1_LOC_69/Y 0.10fF
C36379 INVX1_LOC_239/Y D_GATE_579 0.25fF
C36380 INVX1_LOC_276/A NOR2X1_LOC_686/B 0.04fF
C36381 NAND2X1_LOC_850/Y NAND2X1_LOC_392/Y 0.02fF
C36382 INVX1_LOC_49/A NOR2X1_LOC_163/Y 0.03fF
C36383 INVX1_LOC_14/A INVX1_LOC_14/Y 0.04fF
C36384 INVX1_LOC_241/A INVX1_LOC_22/A 0.27fF
C36385 NAND2X1_LOC_474/Y NOR2X1_LOC_536/A 0.03fF
C36386 NOR2X1_LOC_171/Y NOR2X1_LOC_172/Y 0.22fF
C36387 INVX1_LOC_14/A NAND2X1_LOC_618/a_36_24# 0.01fF
C36388 NOR2X1_LOC_392/Y NOR2X1_LOC_861/a_36_216# 0.00fF
C36389 INVX1_LOC_159/A INVX1_LOC_6/A 0.18fF
C36390 INVX1_LOC_28/A NAND2X1_LOC_464/Y 0.02fF
C36391 NAND2X1_LOC_493/Y NOR2X1_LOC_492/Y 0.17fF
C36392 INVX1_LOC_229/Y NOR2X1_LOC_505/Y 0.06fF
C36393 INVX1_LOC_54/A INVX1_LOC_306/Y 0.03fF
C36394 NOR2X1_LOC_191/B INVX1_LOC_6/A 0.33fF
C36395 NOR2X1_LOC_89/A NAND2X1_LOC_454/Y 0.07fF
C36396 INVX1_LOC_19/A NAND2X1_LOC_99/A 0.16fF
C36397 NOR2X1_LOC_763/A INVX1_LOC_118/A 0.25fF
C36398 NOR2X1_LOC_298/Y INVX1_LOC_22/A 0.02fF
C36399 INVX1_LOC_45/A NOR2X1_LOC_332/B 0.01fF
C36400 NOR2X1_LOC_742/A NOR2X1_LOC_718/B 0.03fF
C36401 NAND2X1_LOC_214/B NOR2X1_LOC_216/B 0.08fF
C36402 INVX1_LOC_55/A INVX1_LOC_37/A 0.01fF
C36403 NOR2X1_LOC_570/B NOR2X1_LOC_74/A 0.00fF
C36404 INVX1_LOC_136/A NOR2X1_LOC_124/A 0.01fF
C36405 INVX1_LOC_283/Y INVX1_LOC_6/A 0.00fF
C36406 NAND2X1_LOC_63/Y NOR2X1_LOC_383/B 0.03fF
C36407 INVX1_LOC_31/A VDD 5.21fF
C36408 NAND2X1_LOC_570/Y NOR2X1_LOC_19/B 0.04fF
C36409 INVX1_LOC_255/Y D_INPUT_0 0.14fF
C36410 INVX1_LOC_17/A INVX1_LOC_38/A 6.34fF
C36411 INVX1_LOC_296/A INPUT_7 0.06fF
C36412 INVX1_LOC_133/A INVX1_LOC_23/A 0.07fF
C36413 INVX1_LOC_13/A INVX1_LOC_135/A 0.13fF
C36414 INVX1_LOC_85/Y NOR2X1_LOC_738/a_36_216# 0.00fF
C36415 INVX1_LOC_27/A NOR2X1_LOC_216/B 0.10fF
C36416 NOR2X1_LOC_430/A NOR2X1_LOC_588/A 0.18fF
C36417 INVX1_LOC_36/A NOR2X1_LOC_280/Y 0.04fF
C36418 INVX1_LOC_77/A NOR2X1_LOC_269/Y 0.42fF
C36419 NOR2X1_LOC_754/A NOR2X1_LOC_693/Y 0.04fF
C36420 NAND2X1_LOC_341/A D_GATE_366 0.01fF
C36421 INVX1_LOC_229/Y NOR2X1_LOC_700/Y 0.04fF
C36422 NAND2X1_LOC_51/B INVX1_LOC_192/Y 0.13fF
C36423 NOR2X1_LOC_577/Y NOR2X1_LOC_139/Y 0.31fF
C36424 NOR2X1_LOC_134/a_36_216# INVX1_LOC_19/Y 0.00fF
C36425 NOR2X1_LOC_168/Y NOR2X1_LOC_35/Y 0.01fF
C36426 NOR2X1_LOC_577/Y NAND2X1_LOC_655/A 0.12fF
C36427 INVX1_LOC_13/A NOR2X1_LOC_560/A -0.02fF
C36428 NAND2X1_LOC_794/B INVX1_LOC_84/A 0.07fF
C36429 NOR2X1_LOC_456/Y INVX1_LOC_99/A 0.42fF
C36430 INVX1_LOC_200/A INVX1_LOC_185/A 0.01fF
C36431 NOR2X1_LOC_589/A NAND2X1_LOC_842/B 0.34fF
C36432 D_INPUT_0 NOR2X1_LOC_71/Y 0.03fF
C36433 NAND2X1_LOC_53/Y NAND2X1_LOC_93/B 0.07fF
C36434 NAND2X1_LOC_860/A NAND2X1_LOC_254/Y 0.01fF
C36435 INVX1_LOC_111/A VDD 0.00fF
C36436 INVX1_LOC_64/A NOR2X1_LOC_671/Y 1.92fF
C36437 NOR2X1_LOC_561/Y NAND2X1_LOC_830/a_36_24# 0.00fF
C36438 NOR2X1_LOC_473/B NAND2X1_LOC_140/A 0.26fF
C36439 NAND2X1_LOC_308/Y NAND2X1_LOC_729/B 0.22fF
C36440 INVX1_LOC_48/Y INVX1_LOC_84/A 0.52fF
C36441 INVX1_LOC_31/A NOR2X1_LOC_846/a_36_216# 0.00fF
C36442 D_INPUT_0 NOR2X1_LOC_644/A 0.00fF
C36443 INVX1_LOC_222/Y INVX1_LOC_19/A 0.07fF
C36444 INVX1_LOC_234/A NOR2X1_LOC_19/B 0.11fF
C36445 NAND2X1_LOC_812/A INVX1_LOC_20/A 0.00fF
C36446 INVX1_LOC_28/A NAND2X1_LOC_691/a_36_24# 0.00fF
C36447 NAND2X1_LOC_862/A NOR2X1_LOC_167/Y 0.01fF
C36448 NAND2X1_LOC_733/Y INVX1_LOC_185/A 0.23fF
C36449 INVX1_LOC_57/Y INVX1_LOC_118/A 0.82fF
C36450 INVX1_LOC_182/Y NAND2X1_LOC_656/Y 0.09fF
C36451 NAND2X1_LOC_714/B INVX1_LOC_49/Y 0.03fF
C36452 INVX1_LOC_246/A NOR2X1_LOC_88/Y 0.07fF
C36453 NOR2X1_LOC_307/B INVX1_LOC_186/A 0.03fF
C36454 NOR2X1_LOC_773/Y INVX1_LOC_98/A 0.02fF
C36455 INVX1_LOC_13/A NOR2X1_LOC_391/B 2.40fF
C36456 NAND2X1_LOC_9/Y INVX1_LOC_4/A 0.03fF
C36457 NOR2X1_LOC_360/Y INVX1_LOC_9/A 1.01fF
C36458 NOR2X1_LOC_773/Y NOR2X1_LOC_78/A 0.07fF
C36459 INVX1_LOC_123/A INVX1_LOC_16/A 0.51fF
C36460 NAND2X1_LOC_35/Y INVX1_LOC_3/Y 0.04fF
C36461 INVX1_LOC_90/A NOR2X1_LOC_171/Y 0.01fF
C36462 NAND2X1_LOC_741/B NAND2X1_LOC_802/Y 0.15fF
C36463 INVX1_LOC_269/A INVX1_LOC_240/Y 0.01fF
C36464 NOR2X1_LOC_309/Y NOR2X1_LOC_280/Y 0.04fF
C36465 NOR2X1_LOC_512/Y INVX1_LOC_118/A 0.28fF
C36466 NAND2X1_LOC_796/B INVX1_LOC_42/A 0.15fF
C36467 NOR2X1_LOC_178/Y NAND2X1_LOC_269/a_36_24# 0.00fF
C36468 NOR2X1_LOC_147/B NOR2X1_LOC_706/B 0.11fF
C36469 INVX1_LOC_56/Y INVX1_LOC_91/A 0.01fF
C36470 NOR2X1_LOC_15/Y NAND2X1_LOC_74/B 0.10fF
C36471 INVX1_LOC_256/Y INVX1_LOC_95/Y 0.13fF
C36472 INVX1_LOC_271/Y NOR2X1_LOC_717/A 0.01fF
C36473 INVX1_LOC_14/A NOR2X1_LOC_831/Y 0.01fF
C36474 NOR2X1_LOC_290/Y VDD 0.12fF
C36475 INVX1_LOC_90/A NOR2X1_LOC_594/Y 0.33fF
C36476 NOR2X1_LOC_798/A INVX1_LOC_4/A 0.06fF
C36477 NAND2X1_LOC_758/a_36_24# INVX1_LOC_117/Y 0.00fF
C36478 INVX1_LOC_191/Y VDD 0.45fF
C36479 INVX1_LOC_111/Y INVX1_LOC_14/Y 0.62fF
C36480 NOR2X1_LOC_505/a_36_216# INVX1_LOC_46/A 0.01fF
C36481 NAND2X1_LOC_468/B INVX1_LOC_22/A 0.05fF
C36482 NAND2X1_LOC_850/Y INVX1_LOC_46/A 0.07fF
C36483 NOR2X1_LOC_304/Y NOR2X1_LOC_409/B 0.10fF
C36484 NOR2X1_LOC_606/a_36_216# NAND2X1_LOC_773/B 0.00fF
C36485 NAND2X1_LOC_593/Y INVX1_LOC_92/A 0.03fF
C36486 NOR2X1_LOC_332/A NOR2X1_LOC_78/A 0.05fF
C36487 NOR2X1_LOC_208/Y NOR2X1_LOC_197/B 0.16fF
C36488 INVX1_LOC_180/A NAND2X1_LOC_798/B 0.35fF
C36489 INVX1_LOC_236/A NOR2X1_LOC_152/A 0.21fF
C36490 INVX1_LOC_122/Y NOR2X1_LOC_814/A 0.55fF
C36491 INVX1_LOC_308/A INVX1_LOC_57/A 0.01fF
C36492 INVX1_LOC_49/A INVX1_LOC_179/A 0.06fF
C36493 NAND2X1_LOC_218/B NAND2X1_LOC_141/Y -0.01fF
C36494 NAND2X1_LOC_479/Y NOR2X1_LOC_357/Y 0.07fF
C36495 NOR2X1_LOC_757/Y NOR2X1_LOC_363/Y 0.03fF
C36496 NAND2X1_LOC_859/Y VDD 0.82fF
C36497 NOR2X1_LOC_230/Y INVX1_LOC_12/A 0.14fF
C36498 INVX1_LOC_24/A INVX1_LOC_63/A 5.31fF
C36499 INVX1_LOC_58/A NAND2X1_LOC_35/Y 0.16fF
C36500 NAND2X1_LOC_742/a_36_24# NOR2X1_LOC_829/A 0.01fF
C36501 NAND2X1_LOC_9/Y INVX1_LOC_64/A 0.17fF
C36502 NOR2X1_LOC_635/a_36_216# NOR2X1_LOC_639/B 0.02fF
C36503 INVX1_LOC_226/Y NOR2X1_LOC_536/A 0.09fF
C36504 INVX1_LOC_286/A NOR2X1_LOC_74/A 1.57fF
C36505 INVX1_LOC_39/A NOR2X1_LOC_383/B 0.03fF
C36506 NOR2X1_LOC_731/A NOR2X1_LOC_155/A 0.03fF
C36507 NAND2X1_LOC_656/A INVX1_LOC_19/A 0.72fF
C36508 INVX1_LOC_38/Y NOR2X1_LOC_416/A 0.02fF
C36509 INVX1_LOC_17/A NAND2X1_LOC_223/A 0.00fF
C36510 INVX1_LOC_21/A INVX1_LOC_224/Y 0.02fF
C36511 NOR2X1_LOC_68/A NOR2X1_LOC_89/A 0.09fF
C36512 NAND2X1_LOC_53/Y NAND2X1_LOC_470/B 0.32fF
C36513 NOR2X1_LOC_510/Y INVX1_LOC_23/A 0.11fF
C36514 INVX1_LOC_53/A NOR2X1_LOC_674/a_36_216# 0.01fF
C36515 INVX1_LOC_134/A NOR2X1_LOC_334/Y 0.02fF
C36516 NOR2X1_LOC_252/Y INVX1_LOC_38/A 0.04fF
C36517 INVX1_LOC_2/A INVX1_LOC_179/A 0.03fF
C36518 INVX1_LOC_286/A NOR2X1_LOC_9/Y 0.13fF
C36519 INVX1_LOC_313/A VDD 0.11fF
C36520 INVX1_LOC_13/A INVX1_LOC_280/A 0.20fF
C36521 NOR2X1_LOC_557/Y INVX1_LOC_63/A 0.07fF
C36522 NOR2X1_LOC_574/A NOR2X1_LOC_697/Y 0.00fF
C36523 INVX1_LOC_18/A NOR2X1_LOC_114/Y 0.00fF
C36524 NAND2X1_LOC_67/a_36_24# INVX1_LOC_50/A 0.00fF
C36525 NOR2X1_LOC_91/A NOR2X1_LOC_361/B 0.08fF
C36526 NAND2X1_LOC_866/B VDD 0.87fF
C36527 INVX1_LOC_10/A NOR2X1_LOC_536/A 0.56fF
C36528 NOR2X1_LOC_360/Y NOR2X1_LOC_861/Y 0.03fF
C36529 INVX1_LOC_21/A NAND2X1_LOC_793/B 0.03fF
C36530 NAND2X1_LOC_579/A INVX1_LOC_57/A 0.09fF
C36531 INVX1_LOC_90/A NOR2X1_LOC_706/B 0.03fF
C36532 NOR2X1_LOC_748/Y NOR2X1_LOC_641/Y 0.20fF
C36533 INVX1_LOC_95/A NOR2X1_LOC_74/A 0.07fF
C36534 NOR2X1_LOC_405/A NOR2X1_LOC_188/A 2.05fF
C36535 INVX1_LOC_50/A INVX1_LOC_269/A 0.07fF
C36536 INVX1_LOC_55/Y INVX1_LOC_139/Y 0.03fF
C36537 INVX1_LOC_64/A NOR2X1_LOC_798/A 0.03fF
C36538 NAND2X1_LOC_555/Y NAND2X1_LOC_223/A 0.09fF
C36539 NOR2X1_LOC_178/Y NAND2X1_LOC_540/a_36_24# 0.00fF
C36540 INVX1_LOC_226/Y NAND2X1_LOC_93/B 0.00fF
C36541 NOR2X1_LOC_437/a_36_216# INVX1_LOC_290/Y 0.01fF
C36542 NAND2X1_LOC_807/Y VDD 0.58fF
C36543 NOR2X1_LOC_84/Y INVX1_LOC_84/A 0.72fF
C36544 NOR2X1_LOC_71/Y NAND2X1_LOC_848/A 0.03fF
C36545 INVX1_LOC_2/A INVX1_LOC_250/Y 0.19fF
C36546 INVX1_LOC_77/A NOR2X1_LOC_633/a_36_216# 0.00fF
C36547 NOR2X1_LOC_590/A NOR2X1_LOC_278/Y 0.12fF
C36548 NAND2X1_LOC_787/A NOR2X1_LOC_92/Y 0.00fF
C36549 NOR2X1_LOC_202/Y NOR2X1_LOC_357/Y 0.04fF
C36550 NOR2X1_LOC_482/Y INVX1_LOC_84/A 0.00fF
C36551 NOR2X1_LOC_361/B INVX1_LOC_23/A 0.18fF
C36552 NOR2X1_LOC_226/A NAND2X1_LOC_267/a_36_24# 0.01fF
C36553 NOR2X1_LOC_436/a_36_216# NOR2X1_LOC_798/A 0.00fF
C36554 INVX1_LOC_55/Y INVX1_LOC_10/Y 0.03fF
C36555 NAND2X1_LOC_363/B INVX1_LOC_24/Y 0.00fF
C36556 INVX1_LOC_143/A INVX1_LOC_63/A 0.14fF
C36557 INVX1_LOC_282/A INVX1_LOC_46/A 0.18fF
C36558 INVX1_LOC_200/Y NAND2X1_LOC_550/A 0.02fF
C36559 NOR2X1_LOC_720/B NAND2X1_LOC_207/B 0.01fF
C36560 INVX1_LOC_10/A NAND2X1_LOC_93/B 0.55fF
C36561 NAND2X1_LOC_692/a_36_24# INVX1_LOC_92/A 0.01fF
C36562 NAND2X1_LOC_808/A INVX1_LOC_185/A 0.00fF
C36563 NAND2X1_LOC_514/Y NOR2X1_LOC_334/Y 0.01fF
C36564 INVX1_LOC_56/Y NOR2X1_LOC_179/Y 0.01fF
C36565 NOR2X1_LOC_590/A NOR2X1_LOC_844/a_36_216# 0.00fF
C36566 D_INPUT_0 NAND2X1_LOC_243/Y 0.05fF
C36567 NOR2X1_LOC_350/A INVX1_LOC_15/A 0.03fF
C36568 INVX1_LOC_269/A NAND2X1_LOC_72/Y 0.03fF
C36569 INVX1_LOC_226/Y INVX1_LOC_3/A 0.23fF
C36570 INVX1_LOC_22/A NOR2X1_LOC_66/Y 0.03fF
C36571 INVX1_LOC_123/A NOR2X1_LOC_35/Y 0.03fF
C36572 NOR2X1_LOC_130/A NOR2X1_LOC_435/A 0.04fF
C36573 INVX1_LOC_134/Y NOR2X1_LOC_777/B 0.01fF
C36574 INVX1_LOC_146/Y INVX1_LOC_6/A 0.01fF
C36575 NOR2X1_LOC_644/Y INVX1_LOC_263/Y 0.01fF
C36576 NOR2X1_LOC_111/A NOR2X1_LOC_527/Y 0.08fF
C36577 NOR2X1_LOC_92/Y NOR2X1_LOC_791/Y 0.13fF
C36578 VDD INVX1_LOC_6/A 1.52fF
C36579 NOR2X1_LOC_828/A INVX1_LOC_307/Y 0.00fF
C36580 INVX1_LOC_298/Y NOR2X1_LOC_457/B 0.07fF
C36581 INVX1_LOC_290/A INVX1_LOC_84/A 0.03fF
C36582 NOR2X1_LOC_388/Y INVX1_LOC_32/A 0.03fF
C36583 INVX1_LOC_35/A INVX1_LOC_225/Y 0.01fF
C36584 NOR2X1_LOC_567/B INVX1_LOC_9/A 0.07fF
C36585 NOR2X1_LOC_160/B INVX1_LOC_292/Y 0.07fF
C36586 NOR2X1_LOC_644/Y INVX1_LOC_42/A 0.05fF
C36587 NAND2X1_LOC_198/B NOR2X1_LOC_318/A 0.37fF
C36588 NOR2X1_LOC_433/A NAND2X1_LOC_454/Y 0.07fF
C36589 NOR2X1_LOC_595/Y INVX1_LOC_76/A 0.17fF
C36590 NOR2X1_LOC_172/Y INVX1_LOC_94/Y 0.17fF
C36591 NOR2X1_LOC_593/Y NAND2X1_LOC_454/Y 1.94fF
C36592 INVX1_LOC_58/A NOR2X1_LOC_723/a_36_216# 0.00fF
C36593 INVX1_LOC_24/A NOR2X1_LOC_65/Y 0.03fF
C36594 NOR2X1_LOC_312/Y INVX1_LOC_285/A 0.02fF
C36595 INVX1_LOC_5/A NOR2X1_LOC_45/Y 0.03fF
C36596 INVX1_LOC_77/A INVX1_LOC_26/A 0.03fF
C36597 NOR2X1_LOC_186/Y NAND2X1_LOC_337/B 0.09fF
C36598 INVX1_LOC_21/A NOR2X1_LOC_103/Y 0.00fF
C36599 NAND2X1_LOC_553/A INVX1_LOC_43/Y 0.02fF
C36600 NAND2X1_LOC_541/Y INVX1_LOC_42/A 0.03fF
C36601 NOR2X1_LOC_186/Y NOR2X1_LOC_816/A 0.92fF
C36602 NOR2X1_LOC_74/A INVX1_LOC_54/A 0.07fF
C36603 INVX1_LOC_286/Y NOR2X1_LOC_109/Y 0.10fF
C36604 INVX1_LOC_135/A NAND2X1_LOC_489/Y 0.03fF
C36605 INVX1_LOC_21/A NOR2X1_LOC_541/Y 0.71fF
C36606 INVX1_LOC_89/A NOR2X1_LOC_673/A 0.06fF
C36607 NAND2X1_LOC_132/a_36_24# NAND2X1_LOC_93/B 0.01fF
C36608 NAND2X1_LOC_338/B INVX1_LOC_19/Y 0.01fF
C36609 NOR2X1_LOC_130/A INVX1_LOC_63/A 0.08fF
C36610 NAND2X1_LOC_119/a_36_24# NAND2X1_LOC_99/A 0.01fF
C36611 NOR2X1_LOC_788/B INVX1_LOC_220/A 0.18fF
C36612 NOR2X1_LOC_781/A INVX1_LOC_29/A 0.00fF
C36613 NOR2X1_LOC_609/A INVX1_LOC_29/Y 0.18fF
C36614 NOR2X1_LOC_790/B NOR2X1_LOC_703/B 0.15fF
C36615 INVX1_LOC_217/A NOR2X1_LOC_754/Y 0.03fF
C36616 INVX1_LOC_243/A D_INPUT_5 0.01fF
C36617 INVX1_LOC_58/A INVX1_LOC_94/A 0.10fF
C36618 NOR2X1_LOC_91/A NOR2X1_LOC_132/Y 0.06fF
C36619 NOR2X1_LOC_52/B NAND2X1_LOC_454/Y 0.08fF
C36620 NOR2X1_LOC_510/Y INVX1_LOC_31/A 0.05fF
C36621 NAND2X1_LOC_573/Y NAND2X1_LOC_337/B 0.02fF
C36622 NAND2X1_LOC_573/Y NOR2X1_LOC_816/A 0.00fF
C36623 NOR2X1_LOC_335/a_36_216# INVX1_LOC_29/A 0.00fF
C36624 NAND2X1_LOC_550/A NAND2X1_LOC_493/Y 0.04fF
C36625 NOR2X1_LOC_208/A NOR2X1_LOC_197/B 0.09fF
C36626 NOR2X1_LOC_227/B NOR2X1_LOC_160/B 0.04fF
C36627 INVX1_LOC_36/A INVX1_LOC_38/Y 0.00fF
C36628 NAND2X1_LOC_860/A INVX1_LOC_314/Y 1.43fF
C36629 INVX1_LOC_313/A INVX1_LOC_133/A 0.02fF
C36630 NAND2X1_LOC_724/A NOR2X1_LOC_816/A 0.08fF
C36631 NOR2X1_LOC_490/Y NAND2X1_LOC_489/Y 0.02fF
C36632 INVX1_LOC_21/A INVX1_LOC_45/A 0.47fF
C36633 NAND2X1_LOC_593/Y INVX1_LOC_53/A 0.03fF
C36634 NOR2X1_LOC_76/A INVX1_LOC_29/A 0.42fF
C36635 INVX1_LOC_124/A INVX1_LOC_26/A 0.01fF
C36636 INVX1_LOC_21/A NOR2X1_LOC_568/A 0.23fF
C36637 NOR2X1_LOC_132/Y INVX1_LOC_23/A 0.05fF
C36638 INVX1_LOC_290/A INVX1_LOC_15/A 0.09fF
C36639 INVX1_LOC_27/A NAND2X1_LOC_670/a_36_24# 0.00fF
C36640 NOR2X1_LOC_180/B INVX1_LOC_29/A 0.04fF
C36641 NOR2X1_LOC_410/Y NOR2X1_LOC_242/A 0.04fF
C36642 NOR2X1_LOC_329/B INVX1_LOC_19/A 1.24fF
C36643 INVX1_LOC_258/Y INVX1_LOC_72/A 0.03fF
C36644 NOR2X1_LOC_357/Y NOR2X1_LOC_57/a_36_216# 0.00fF
C36645 NAND2X1_LOC_840/a_36_24# NOR2X1_LOC_654/A 0.00fF
C36646 NAND2X1_LOC_729/Y NAND2X1_LOC_740/Y 0.04fF
C36647 INVX1_LOC_2/A NOR2X1_LOC_693/Y 0.07fF
C36648 NOR2X1_LOC_831/B NOR2X1_LOC_114/A 0.09fF
C36649 NOR2X1_LOC_789/A NOR2X1_LOC_38/B 0.01fF
C36650 NOR2X1_LOC_92/Y INVX1_LOC_30/A 0.34fF
C36651 NAND2X1_LOC_575/a_36_24# INVX1_LOC_141/Y 0.00fF
C36652 NOR2X1_LOC_6/B NOR2X1_LOC_414/Y 0.10fF
C36653 INVX1_LOC_1/A NOR2X1_LOC_726/Y 0.01fF
C36654 INVX1_LOC_58/A NAND2X1_LOC_465/Y 0.01fF
C36655 INVX1_LOC_24/Y INVX1_LOC_30/A 0.53fF
C36656 D_INPUT_4 INVX1_LOC_19/A 0.01fF
C36657 NOR2X1_LOC_826/Y INVX1_LOC_217/Y 0.01fF
C36658 INVX1_LOC_41/A NAND2X1_LOC_363/B 0.04fF
C36659 INVX1_LOC_233/Y INVX1_LOC_237/Y 0.00fF
C36660 NOR2X1_LOC_91/A INVX1_LOC_280/Y 0.06fF
C36661 NOR2X1_LOC_831/B INVX1_LOC_91/A 0.10fF
C36662 INVX1_LOC_136/A NOR2X1_LOC_15/Y 0.44fF
C36663 INVX1_LOC_132/A INVX1_LOC_5/A 0.08fF
C36664 INVX1_LOC_135/A INVX1_LOC_32/A 0.92fF
C36665 INVX1_LOC_90/A NOR2X1_LOC_157/a_36_216# 0.01fF
C36666 NAND2X1_LOC_112/Y INVX1_LOC_78/A 0.06fF
C36667 NOR2X1_LOC_235/a_36_216# NOR2X1_LOC_384/Y 0.01fF
C36668 NOR2X1_LOC_647/a_36_216# INPUT_3 0.00fF
C36669 INVX1_LOC_230/Y NAND2X1_LOC_767/a_36_24# 0.00fF
C36670 INVX1_LOC_73/A INVX1_LOC_29/A 0.03fF
C36671 NOR2X1_LOC_598/B NOR2X1_LOC_731/A 0.01fF
C36672 INVX1_LOC_75/A INVX1_LOC_272/A 0.31fF
C36673 INVX1_LOC_21/A INVX1_LOC_71/A 0.28fF
C36674 INVX1_LOC_177/A INVX1_LOC_23/A 0.07fF
C36675 NAND2X1_LOC_552/A NAND2X1_LOC_640/Y 0.17fF
C36676 INVX1_LOC_304/Y NOR2X1_LOC_754/Y 0.01fF
C36677 INVX1_LOC_27/A NOR2X1_LOC_303/Y 0.00fF
C36678 INVX1_LOC_53/Y NOR2X1_LOC_318/A 0.08fF
C36679 INVX1_LOC_10/A NAND2X1_LOC_470/B 0.69fF
C36680 NOR2X1_LOC_667/a_36_216# INVX1_LOC_286/Y 0.00fF
C36681 INVX1_LOC_278/A NOR2X1_LOC_84/Y 0.12fF
C36682 NOR2X1_LOC_313/a_36_216# INVX1_LOC_12/A 0.00fF
C36683 NAND2X1_LOC_739/B NAND2X1_LOC_303/Y 0.03fF
C36684 INVX1_LOC_225/A NAND2X1_LOC_552/A 0.01fF
C36685 NOR2X1_LOC_843/A NOR2X1_LOC_434/Y 0.01fF
C36686 INVX1_LOC_224/A NOR2X1_LOC_68/A 0.63fF
C36687 INVX1_LOC_35/A INVX1_LOC_266/Y 0.03fF
C36688 NAND2X1_LOC_141/A NOR2X1_LOC_660/Y 0.56fF
C36689 INVX1_LOC_1/Y NOR2X1_LOC_481/a_36_216# 0.01fF
C36690 INVX1_LOC_41/A NOR2X1_LOC_791/Y 0.02fF
C36691 NOR2X1_LOC_604/a_36_216# NOR2X1_LOC_78/B 0.00fF
C36692 INVX1_LOC_88/A NOR2X1_LOC_351/a_36_216# 0.00fF
C36693 INVX1_LOC_6/A INVX1_LOC_133/A 0.00fF
C36694 NAND2X1_LOC_348/A NOR2X1_LOC_346/A 0.01fF
C36695 INVX1_LOC_11/A NOR2X1_LOC_68/A 0.32fF
C36696 NAND2X1_LOC_243/B INVX1_LOC_20/A 0.01fF
C36697 VDD INVX1_LOC_131/Y 0.25fF
C36698 INVX1_LOC_135/A NAND2X1_LOC_175/Y 0.10fF
C36699 INVX1_LOC_41/A NAND2X1_LOC_63/a_36_24# 0.00fF
C36700 INVX1_LOC_233/A NAND2X1_LOC_850/Y 0.00fF
C36701 NOR2X1_LOC_91/A NAND2X1_LOC_573/A 0.02fF
C36702 INVX1_LOC_90/A INVX1_LOC_94/Y 0.03fF
C36703 INVX1_LOC_181/Y NAND2X1_LOC_793/Y 0.10fF
C36704 NOR2X1_LOC_74/A NOR2X1_LOC_48/B 0.14fF
C36705 D_INPUT_1 INVX1_LOC_16/A 0.20fF
C36706 INVX1_LOC_289/Y INVX1_LOC_209/Y 0.02fF
C36707 D_INPUT_0 INVX1_LOC_16/Y 0.03fF
C36708 INVX1_LOC_36/A INVX1_LOC_286/Y 0.03fF
C36709 VDD NAND2X1_LOC_810/B 0.08fF
C36710 INVX1_LOC_224/A NOR2X1_LOC_545/A 0.01fF
C36711 INVX1_LOC_210/Y NAND2X1_LOC_510/A 0.03fF
C36712 NOR2X1_LOC_32/B INVX1_LOC_316/Y 0.02fF
C36713 INVX1_LOC_88/A NOR2X1_LOC_577/Y 0.10fF
C36714 D_INPUT_0 NOR2X1_LOC_39/Y 0.20fF
C36715 INVX1_LOC_119/Y INVX1_LOC_20/A 0.03fF
C36716 NAND2X1_LOC_848/A NAND2X1_LOC_243/Y 0.46fF
C36717 NOR2X1_LOC_130/A NOR2X1_LOC_65/Y 0.05fF
C36718 NOR2X1_LOC_155/A INVX1_LOC_117/A 0.57fF
C36719 NAND2X1_LOC_149/Y NOR2X1_LOC_154/a_36_216# 0.01fF
C36720 INVX1_LOC_34/A NAND2X1_LOC_561/B 0.16fF
C36721 NAND2X1_LOC_550/A NOR2X1_LOC_495/Y 0.15fF
C36722 NAND2X1_LOC_287/B INVX1_LOC_285/A 0.01fF
C36723 INVX1_LOC_17/A INVX1_LOC_33/A 0.07fF
C36724 INVX1_LOC_194/A INVX1_LOC_163/A 0.04fF
C36725 INPUT_4 NOR2X1_LOC_11/Y 0.06fF
C36726 INPUT_1 NOR2X1_LOC_693/Y 0.07fF
C36727 INVX1_LOC_178/Y NOR2X1_LOC_649/B 0.04fF
C36728 NOR2X1_LOC_391/B INVX1_LOC_32/A 0.02fF
C36729 INVX1_LOC_13/Y NOR2X1_LOC_175/B 0.04fF
C36730 NAND2X1_LOC_9/Y NOR2X1_LOC_721/a_36_216# 0.01fF
C36731 NOR2X1_LOC_665/A NOR2X1_LOC_678/A 0.03fF
C36732 INVX1_LOC_163/A NOR2X1_LOC_399/A 0.04fF
C36733 INVX1_LOC_223/Y NAND2X1_LOC_165/a_36_24# 0.01fF
C36734 NOR2X1_LOC_186/Y NOR2X1_LOC_773/Y 0.01fF
C36735 D_INPUT_0 NAND2X1_LOC_205/A 0.54fF
C36736 NOR2X1_LOC_772/B INVX1_LOC_22/A 0.19fF
C36737 INVX1_LOC_34/A NAND2X1_LOC_719/a_36_24# 0.00fF
C36738 INVX1_LOC_36/A INVX1_LOC_159/A 0.04fF
C36739 NOR2X1_LOC_78/B NOR2X1_LOC_852/Y 0.04fF
C36740 NOR2X1_LOC_78/A INVX1_LOC_42/A 0.07fF
C36741 INVX1_LOC_90/A INVX1_LOC_296/A 0.03fF
C36742 NAND2X1_LOC_361/Y NOR2X1_LOC_160/B 0.10fF
C36743 INVX1_LOC_36/A NOR2X1_LOC_191/B 0.19fF
C36744 INVX1_LOC_30/A NAND2X1_LOC_837/Y 0.10fF
C36745 INVX1_LOC_13/Y INVX1_LOC_22/A 0.03fF
C36746 NAND2X1_LOC_637/Y INVX1_LOC_117/Y 0.31fF
C36747 INVX1_LOC_16/A NOR2X1_LOC_652/Y 0.07fF
C36748 INVX1_LOC_225/A NAND2X1_LOC_337/B 0.01fF
C36749 INVX1_LOC_185/A INVX1_LOC_92/A 0.03fF
C36750 INVX1_LOC_58/A NAND2X1_LOC_307/a_36_24# 0.01fF
C36751 NAND2X1_LOC_462/B INVX1_LOC_253/Y 0.03fF
C36752 VDD INVX1_LOC_301/A 0.12fF
C36753 INVX1_LOC_236/Y NAND2X1_LOC_354/B 0.04fF
C36754 NOR2X1_LOC_369/Y NOR2X1_LOC_309/Y 0.04fF
C36755 NAND2X1_LOC_93/B INVX1_LOC_307/A 0.03fF
C36756 INVX1_LOC_27/Y NOR2X1_LOC_271/Y 0.13fF
C36757 INVX1_LOC_20/A INVX1_LOC_284/A 1.03fF
C36758 VDD NOR2X1_LOC_633/A 0.03fF
C36759 NOR2X1_LOC_552/A INVX1_LOC_32/A 0.07fF
C36760 D_INPUT_1 INVX1_LOC_28/A 0.17fF
C36761 NAND2X1_LOC_724/A NOR2X1_LOC_773/Y 0.00fF
C36762 NAND2X1_LOC_803/a_36_24# NOR2X1_LOC_109/Y 0.01fF
C36763 INVX1_LOC_41/A INVX1_LOC_30/A 0.40fF
C36764 NAND2X1_LOC_464/A INVX1_LOC_42/A 0.00fF
C36765 NOR2X1_LOC_68/A NOR2X1_LOC_433/A 0.07fF
C36766 NOR2X1_LOC_276/B INVX1_LOC_77/A 0.02fF
C36767 INVX1_LOC_286/Y NOR2X1_LOC_309/Y 0.10fF
C36768 INVX1_LOC_11/A NOR2X1_LOC_520/a_36_216# 0.00fF
C36769 INVX1_LOC_98/A INVX1_LOC_78/A 0.18fF
C36770 INVX1_LOC_83/A NOR2X1_LOC_849/A 0.03fF
C36771 NOR2X1_LOC_514/A INVX1_LOC_80/Y 0.01fF
C36772 INVX1_LOC_174/A INVX1_LOC_192/Y 0.10fF
C36773 NOR2X1_LOC_268/a_36_216# INVX1_LOC_49/A 0.01fF
C36774 NOR2X1_LOC_763/A INPUT_5 0.19fF
C36775 NOR2X1_LOC_703/B NOR2X1_LOC_344/A 0.02fF
C36776 INVX1_LOC_40/Y NOR2X1_LOC_6/B 0.01fF
C36777 NOR2X1_LOC_45/B NOR2X1_LOC_158/Y 0.89fF
C36778 NOR2X1_LOC_78/A INVX1_LOC_78/A 0.10fF
C36779 NOR2X1_LOC_582/A INPUT_5 0.03fF
C36780 INVX1_LOC_193/A NOR2X1_LOC_258/Y 0.01fF
C36781 INVX1_LOC_88/A INVX1_LOC_22/A 0.03fF
C36782 NAND2X1_LOC_863/Y NAND2X1_LOC_866/A 0.36fF
C36783 INVX1_LOC_182/Y NOR2X1_LOC_717/A 0.03fF
C36784 INVX1_LOC_21/A NOR2X1_LOC_123/B 0.03fF
C36785 INVX1_LOC_64/A INVX1_LOC_146/A 0.03fF
C36786 NOR2X1_LOC_815/Y NOR2X1_LOC_512/Y 0.06fF
C36787 INVX1_LOC_30/A NAND2X1_LOC_477/A 0.13fF
C36788 INVX1_LOC_76/A D_INPUT_5 0.07fF
C36789 NOR2X1_LOC_833/B INVX1_LOC_117/A 0.03fF
C36790 NOR2X1_LOC_45/B NOR2X1_LOC_25/Y 0.18fF
C36791 INVX1_LOC_256/A NOR2X1_LOC_500/Y 0.13fF
C36792 NAND2X1_LOC_778/Y NAND2X1_LOC_862/Y 0.04fF
C36793 INVX1_LOC_12/A NOR2X1_LOC_536/A 0.25fF
C36794 NOR2X1_LOC_558/A INVX1_LOC_47/Y 0.00fF
C36795 NOR2X1_LOC_273/Y INVX1_LOC_34/A 0.03fF
C36796 INVX1_LOC_285/Y INVX1_LOC_23/A 0.10fF
C36797 NOR2X1_LOC_688/Y INVX1_LOC_143/A 0.01fF
C36798 INVX1_LOC_139/Y INVX1_LOC_32/A 0.03fF
C36799 NOR2X1_LOC_68/A NOR2X1_LOC_52/B 6.39fF
C36800 INVX1_LOC_34/A NOR2X1_LOC_759/Y 0.04fF
C36801 NOR2X1_LOC_598/B NOR2X1_LOC_589/Y 0.02fF
C36802 NOR2X1_LOC_318/B NOR2X1_LOC_481/a_36_216# 0.00fF
C36803 NOR2X1_LOC_541/a_36_216# INVX1_LOC_58/Y 0.01fF
C36804 NOR2X1_LOC_248/Y NAND2X1_LOC_342/Y 0.08fF
C36805 NAND2X1_LOC_563/A INVX1_LOC_61/Y 0.01fF
C36806 NOR2X1_LOC_65/B NOR2X1_LOC_78/A 0.08fF
C36807 INVX1_LOC_136/A INVX1_LOC_96/Y 0.02fF
C36808 NOR2X1_LOC_637/B NOR2X1_LOC_637/a_36_216# 0.00fF
C36809 NOR2X1_LOC_596/A INVX1_LOC_88/Y 0.05fF
C36810 INVX1_LOC_202/A INVX1_LOC_34/A 0.17fF
C36811 INVX1_LOC_45/A NOR2X1_LOC_667/A 0.04fF
C36812 NOR2X1_LOC_346/A INVX1_LOC_38/A 0.01fF
C36813 INVX1_LOC_45/A INVX1_LOC_248/A 0.01fF
C36814 NOR2X1_LOC_197/B INVX1_LOC_63/A 0.01fF
C36815 INVX1_LOC_230/Y NOR2X1_LOC_94/a_36_216# 0.01fF
C36816 NOR2X1_LOC_309/Y NOR2X1_LOC_191/B 0.10fF
C36817 INVX1_LOC_133/A INVX1_LOC_131/Y 0.03fF
C36818 NOR2X1_LOC_813/Y INVX1_LOC_32/A 0.07fF
C36819 INVX1_LOC_235/Y NOR2X1_LOC_575/Y 0.10fF
C36820 INVX1_LOC_226/Y NOR2X1_LOC_606/Y 0.00fF
C36821 NOR2X1_LOC_486/Y NOR2X1_LOC_302/A 0.01fF
C36822 INVX1_LOC_256/A INVX1_LOC_10/A 0.43fF
C36823 INVX1_LOC_2/A NOR2X1_LOC_268/a_36_216# -0.02fF
C36824 NOR2X1_LOC_410/Y NOR2X1_LOC_78/B 0.05fF
C36825 NOR2X1_LOC_361/B INVX1_LOC_313/A 0.05fF
C36826 INVX1_LOC_21/A INVX1_LOC_102/Y 0.07fF
C36827 INVX1_LOC_299/A INVX1_LOC_90/A 0.07fF
C36828 INVX1_LOC_12/A NAND2X1_LOC_93/B 0.03fF
C36829 NOR2X1_LOC_419/Y INVX1_LOC_60/Y 0.10fF
C36830 INVX1_LOC_299/A NOR2X1_LOC_389/B 0.01fF
C36831 INVX1_LOC_32/A INVX1_LOC_280/A 0.27fF
C36832 NOR2X1_LOC_418/Y INVX1_LOC_72/A 0.05fF
C36833 NOR2X1_LOC_538/B INVX1_LOC_90/A 0.02fF
C36834 NOR2X1_LOC_690/A INVX1_LOC_217/Y 0.11fF
C36835 INVX1_LOC_1/A INVX1_LOC_311/Y 0.02fF
C36836 NOR2X1_LOC_790/B INVX1_LOC_91/A 0.08fF
C36837 INVX1_LOC_65/A INVX1_LOC_23/A 0.01fF
C36838 NOR2X1_LOC_389/A NAND2X1_LOC_656/Y 0.10fF
C36839 INVX1_LOC_149/A INVX1_LOC_77/A 0.01fF
C36840 INVX1_LOC_13/Y INVX1_LOC_100/A 0.06fF
C36841 INPUT_3 INVX1_LOC_135/A 0.10fF
C36842 NAND2X1_LOC_569/A NAND2X1_LOC_564/a_36_24# 0.02fF
C36843 INVX1_LOC_11/A NOR2X1_LOC_163/A 0.04fF
C36844 NOR2X1_LOC_134/Y NOR2X1_LOC_71/Y 0.02fF
C36845 NAND2X1_LOC_724/A INVX1_LOC_140/A 0.10fF
C36846 NAND2X1_LOC_363/B NAND2X1_LOC_823/a_36_24# 0.00fF
C36847 NOR2X1_LOC_264/Y NOR2X1_LOC_720/B 0.07fF
C36848 NOR2X1_LOC_589/A INVX1_LOC_72/A 0.96fF
C36849 INVX1_LOC_75/A INVX1_LOC_198/A 0.03fF
C36850 VDD INVX1_LOC_28/Y 0.44fF
C36851 INVX1_LOC_135/A NOR2X1_LOC_201/a_36_216# 0.00fF
C36852 NOR2X1_LOC_590/A NOR2X1_LOC_312/Y 0.00fF
C36853 NOR2X1_LOC_152/A NAND2X1_LOC_175/Y 0.05fF
C36854 INVX1_LOC_75/A NOR2X1_LOC_271/B 0.05fF
C36855 INVX1_LOC_38/A INVX1_LOC_94/Y 0.40fF
C36856 INVX1_LOC_304/A NAND2X1_LOC_793/B 0.98fF
C36857 NOR2X1_LOC_203/Y NOR2X1_LOC_577/Y 0.04fF
C36858 INVX1_LOC_14/Y NOR2X1_LOC_383/B 0.01fF
C36859 VDD INVX1_LOC_270/A 1.53fF
C36860 INVX1_LOC_12/A NOR2X1_LOC_649/B 0.02fF
C36861 NAND2X1_LOC_298/a_36_24# NOR2X1_LOC_727/B 0.00fF
C36862 NOR2X1_LOC_75/Y NOR2X1_LOC_736/Y 0.08fF
C36863 NOR2X1_LOC_498/Y NAND2X1_LOC_722/A 0.00fF
C36864 INVX1_LOC_161/Y NOR2X1_LOC_329/B 0.97fF
C36865 NOR2X1_LOC_391/A NOR2X1_LOC_791/B 0.03fF
C36866 INVX1_LOC_93/A NOR2X1_LOC_528/Y 0.10fF
C36867 NOR2X1_LOC_403/B INVX1_LOC_16/A 0.03fF
C36868 INVX1_LOC_83/A INVX1_LOC_142/A 0.38fF
C36869 NOR2X1_LOC_111/A NOR2X1_LOC_654/A 0.25fF
C36870 INVX1_LOC_5/A NAND2X1_LOC_642/Y 0.08fF
C36871 INVX1_LOC_50/A INVX1_LOC_12/Y 0.03fF
C36872 NOR2X1_LOC_607/Y INVX1_LOC_16/A 0.19fF
C36873 INVX1_LOC_11/A INVX1_LOC_147/A 1.20fF
C36874 NOR2X1_LOC_15/Y NOR2X1_LOC_165/a_36_216# 0.00fF
C36875 INVX1_LOC_303/A INVX1_LOC_22/A 0.07fF
C36876 NAND2X1_LOC_112/Y NOR2X1_LOC_152/Y 0.03fF
C36877 INVX1_LOC_150/Y INVX1_LOC_75/A 0.30fF
C36878 INVX1_LOC_48/Y INVX1_LOC_123/A 0.01fF
C36879 D_INPUT_4 NOR2X1_LOC_22/a_36_216# 0.00fF
C36880 NOR2X1_LOC_279/a_36_216# NAND2X1_LOC_357/B 0.00fF
C36881 NOR2X1_LOC_246/Y NOR2X1_LOC_248/Y 0.09fF
C36882 INVX1_LOC_26/A INVX1_LOC_9/A 4.87fF
C36883 NAND2X1_LOC_361/Y NOR2X1_LOC_516/B 0.10fF
C36884 INVX1_LOC_49/Y NAND2X1_LOC_74/B 0.03fF
C36885 INVX1_LOC_293/A NAND2X1_LOC_348/A 0.00fF
C36886 NOR2X1_LOC_361/B INVX1_LOC_6/A 0.07fF
C36887 NAND2X1_LOC_632/B NAND2X1_LOC_735/B 0.28fF
C36888 NOR2X1_LOC_609/A NOR2X1_LOC_355/A 0.13fF
C36889 INVX1_LOC_225/A NOR2X1_LOC_773/Y 0.02fF
C36890 NAND2X1_LOC_494/a_36_24# INVX1_LOC_25/Y 0.01fF
C36891 NOR2X1_LOC_769/B INVX1_LOC_117/A 0.03fF
C36892 INVX1_LOC_225/Y NOR2X1_LOC_534/a_36_216# 0.01fF
C36893 INVX1_LOC_38/A INVX1_LOC_296/A 0.07fF
C36894 NOR2X1_LOC_557/Y INVX1_LOC_1/Y 0.01fF
C36895 INVX1_LOC_247/Y NOR2X1_LOC_180/B 0.00fF
C36896 NOR2X1_LOC_309/Y NOR2X1_LOC_568/a_36_216# 0.00fF
C36897 NAND2X1_LOC_231/Y NOR2X1_LOC_41/Y 0.08fF
C36898 NOR2X1_LOC_598/B INVX1_LOC_117/A 0.30fF
C36899 VDD NOR2X1_LOC_109/Y 0.14fF
C36900 NOR2X1_LOC_808/A INVX1_LOC_196/A 0.00fF
C36901 INVX1_LOC_243/A NAND2X1_LOC_451/Y 0.03fF
C36902 INVX1_LOC_51/A INVX1_LOC_117/A 0.03fF
C36903 INPUT_3 NOR2X1_LOC_391/B 0.04fF
C36904 INVX1_LOC_179/A NOR2X1_LOC_631/Y 0.00fF
C36905 NOR2X1_LOC_441/Y NOR2X1_LOC_74/A 0.10fF
C36906 NOR2X1_LOC_505/a_36_216# NOR2X1_LOC_505/Y 0.03fF
C36907 INVX1_LOC_45/A NAND2X1_LOC_51/B 0.01fF
C36908 NOR2X1_LOC_51/A INVX1_LOC_296/A 0.07fF
C36909 D_GATE_741 INVX1_LOC_91/A 0.02fF
C36910 INVX1_LOC_114/Y NAND2X1_LOC_220/B 0.21fF
C36911 NAND2X1_LOC_799/A NAND2X1_LOC_655/A 0.07fF
C36912 NOR2X1_LOC_773/Y NAND2X1_LOC_852/Y 0.54fF
C36913 NOR2X1_LOC_403/B INVX1_LOC_28/A 0.19fF
C36914 NAND2X1_LOC_651/B NOR2X1_LOC_467/A 0.26fF
C36915 INVX1_LOC_255/Y NOR2X1_LOC_818/Y 0.01fF
C36916 INVX1_LOC_211/Y NOR2X1_LOC_45/B 0.01fF
C36917 INVX1_LOC_46/A NOR2X1_LOC_440/B 0.01fF
C36918 INVX1_LOC_143/A INVX1_LOC_1/Y 0.09fF
C36919 NOR2X1_LOC_644/A INVX1_LOC_49/A 0.03fF
C36920 INVX1_LOC_124/Y INVX1_LOC_286/A 0.10fF
C36921 INVX1_LOC_24/A NOR2X1_LOC_742/A 0.09fF
C36922 INVX1_LOC_53/A INVX1_LOC_185/A 0.00fF
C36923 NAND2X1_LOC_337/B NAND2X1_LOC_642/Y 0.08fF
C36924 INVX1_LOC_8/A NOR2X1_LOC_76/A 0.24fF
C36925 NOR2X1_LOC_385/a_36_216# NOR2X1_LOC_577/Y 0.01fF
C36926 NOR2X1_LOC_865/Y NOR2X1_LOC_836/A 0.10fF
C36927 INVX1_LOC_58/A NOR2X1_LOC_155/A 0.11fF
C36928 INVX1_LOC_256/A NOR2X1_LOC_799/B 0.01fF
C36929 INVX1_LOC_90/A INVX1_LOC_162/A 0.09fF
C36930 NAND2X1_LOC_722/A NOR2X1_LOC_299/Y 0.46fF
C36931 NAND2X1_LOC_220/B NOR2X1_LOC_467/A 0.03fF
C36932 NOR2X1_LOC_389/B INVX1_LOC_162/A 0.05fF
C36933 NOR2X1_LOC_759/Y INPUT_0 0.00fF
C36934 NAND2X1_LOC_640/Y INVX1_LOC_140/A 0.01fF
C36935 INVX1_LOC_202/A INPUT_0 0.07fF
C36936 INVX1_LOC_2/A NOR2X1_LOC_71/Y 0.03fF
C36937 INVX1_LOC_21/A NOR2X1_LOC_331/B 0.16fF
C36938 INVX1_LOC_147/A NOR2X1_LOC_433/A 0.17fF
C36939 INVX1_LOC_90/A NOR2X1_LOC_315/Y 0.22fF
C36940 INVX1_LOC_26/Y NOR2X1_LOC_691/B 0.01fF
C36941 INVX1_LOC_12/A NAND2X1_LOC_470/B 0.09fF
C36942 INVX1_LOC_72/A INVX1_LOC_167/Y 0.18fF
C36943 INVX1_LOC_31/A INVX1_LOC_316/A -0.01fF
C36944 NOR2X1_LOC_477/a_36_216# INVX1_LOC_199/Y 0.00fF
C36945 INVX1_LOC_311/A INVX1_LOC_71/A 0.10fF
C36946 NOR2X1_LOC_19/B NOR2X1_LOC_84/A 0.31fF
C36947 INVX1_LOC_124/Y INVX1_LOC_95/A 0.00fF
C36948 NOR2X1_LOC_226/A NOR2X1_LOC_71/Y 0.01fF
C36949 NOR2X1_LOC_554/B NOR2X1_LOC_78/A 0.02fF
C36950 INVX1_LOC_25/A INVX1_LOC_84/A 0.14fF
C36951 INVX1_LOC_35/A NAND2X1_LOC_288/A 0.01fF
C36952 NOR2X1_LOC_591/Y INVX1_LOC_28/A 0.04fF
C36953 INVX1_LOC_15/A NOR2X1_LOC_467/A 0.05fF
C36954 INVX1_LOC_18/A NAND2X1_LOC_655/A 0.07fF
C36955 INVX1_LOC_215/A NAND2X1_LOC_660/Y 0.10fF
C36956 INVX1_LOC_15/A NOR2X1_LOC_801/B 0.07fF
C36957 INVX1_LOC_2/A NOR2X1_LOC_644/A 0.07fF
C36958 INVX1_LOC_17/A NOR2X1_LOC_816/Y 0.05fF
C36959 INVX1_LOC_280/Y NAND2X1_LOC_866/B 0.07fF
C36960 INVX1_LOC_299/A INVX1_LOC_38/A 0.07fF
C36961 INVX1_LOC_36/A NOR2X1_LOC_56/Y 0.07fF
C36962 INVX1_LOC_54/Y NOR2X1_LOC_772/A 0.01fF
C36963 NAND2X1_LOC_98/a_36_24# NOR2X1_LOC_96/Y 0.00fF
C36964 INVX1_LOC_312/Y NAND2X1_LOC_655/B 0.01fF
C36965 NOR2X1_LOC_392/Y NOR2X1_LOC_673/A 0.07fF
C36966 NOR2X1_LOC_142/Y NOR2X1_LOC_74/A 0.47fF
C36967 INVX1_LOC_240/A NAND2X1_LOC_863/A 0.42fF
C36968 NOR2X1_LOC_445/Y NOR2X1_LOC_188/A 0.15fF
C36969 NOR2X1_LOC_655/B NOR2X1_LOC_356/A 0.18fF
C36970 NAND2X1_LOC_783/Y NOR2X1_LOC_111/A 0.04fF
C36971 NAND2X1_LOC_842/B NAND2X1_LOC_850/Y 0.03fF
C36972 NOR2X1_LOC_776/a_36_216# INVX1_LOC_117/A 0.00fF
C36973 NAND2X1_LOC_859/Y NOR2X1_LOC_528/a_36_216# 0.00fF
C36974 INVX1_LOC_35/A NOR2X1_LOC_653/Y 0.01fF
C36975 NAND2X1_LOC_564/B INVX1_LOC_135/A 0.10fF
C36976 NAND2X1_LOC_370/a_36_24# INVX1_LOC_84/A 0.00fF
C36977 NOR2X1_LOC_68/A INVX1_LOC_199/A 0.02fF
C36978 INVX1_LOC_89/A NOR2X1_LOC_210/B 0.30fF
C36979 INVX1_LOC_147/A NOR2X1_LOC_52/B 0.18fF
C36980 NOR2X1_LOC_32/B NOR2X1_LOC_662/A 0.07fF
C36981 INVX1_LOC_18/A NAND2X1_LOC_468/B 0.14fF
C36982 INVX1_LOC_153/Y INVX1_LOC_6/A 0.01fF
C36983 INVX1_LOC_215/A D_INPUT_0 0.02fF
C36984 INVX1_LOC_21/A NOR2X1_LOC_592/B 0.03fF
C36985 INVX1_LOC_72/A INVX1_LOC_20/A 0.15fF
C36986 INVX1_LOC_18/A NOR2X1_LOC_683/Y 0.10fF
C36987 NOR2X1_LOC_68/A INVX1_LOC_74/A 0.01fF
C36988 NOR2X1_LOC_584/Y NOR2X1_LOC_651/a_36_216# 0.00fF
C36989 NOR2X1_LOC_78/A NOR2X1_LOC_152/Y 0.14fF
C36990 INVX1_LOC_23/A NAND2X1_LOC_81/B 0.01fF
C36991 INVX1_LOC_61/Y INVX1_LOC_12/Y 0.16fF
C36992 INVX1_LOC_36/A INVX1_LOC_146/Y 0.15fF
C36993 INVX1_LOC_157/A INVX1_LOC_10/A 0.03fF
C36994 INVX1_LOC_36/A VDD 1.77fF
C36995 NOR2X1_LOC_824/A INVX1_LOC_35/Y 0.02fF
C36996 NOR2X1_LOC_567/B INVX1_LOC_179/Y 0.02fF
C36997 NOR2X1_LOC_348/Y INVX1_LOC_307/A 0.00fF
C36998 INVX1_LOC_255/Y INPUT_1 0.08fF
C36999 INVX1_LOC_41/Y NOR2X1_LOC_164/Y 0.10fF
C37000 INVX1_LOC_304/A INVX1_LOC_71/A 0.04fF
C37001 INVX1_LOC_35/A INVX1_LOC_19/A 3.91fF
C37002 NOR2X1_LOC_360/Y INVX1_LOC_76/A 0.39fF
C37003 INVX1_LOC_100/A INVX1_LOC_168/A 0.10fF
C37004 INPUT_3 INVX1_LOC_280/A 0.07fF
C37005 NAND2X1_LOC_165/a_36_24# INVX1_LOC_75/A 0.00fF
C37006 NOR2X1_LOC_267/A VDD 0.09fF
C37007 NOR2X1_LOC_361/B INVX1_LOC_131/Y 0.14fF
C37008 D_INPUT_0 NOR2X1_LOC_373/Y 0.01fF
C37009 NOR2X1_LOC_730/Y INVX1_LOC_196/Y 0.22fF
C37010 NAND2X1_LOC_733/Y NOR2X1_LOC_536/A 0.01fF
C37011 NOR2X1_LOC_497/Y INVX1_LOC_16/A 0.64fF
C37012 NOR2X1_LOC_655/B NOR2X1_LOC_74/A 0.16fF
C37013 INVX1_LOC_50/Y NOR2X1_LOC_814/A 0.12fF
C37014 INVX1_LOC_32/A NAND2X1_LOC_416/a_36_24# 0.00fF
C37015 INVX1_LOC_38/Y INVX1_LOC_63/A 0.07fF
C37016 NOR2X1_LOC_466/a_36_216# NAND2X1_LOC_425/Y 0.01fF
C37017 NOR2X1_LOC_480/A D_GATE_479 0.01fF
C37018 NOR2X1_LOC_201/a_36_216# INVX1_LOC_280/A 0.01fF
C37019 INVX1_LOC_24/A INVX1_LOC_139/A 0.08fF
C37020 NOR2X1_LOC_557/Y INVX1_LOC_93/Y 0.19fF
C37021 NOR2X1_LOC_254/Y NOR2X1_LOC_197/a_36_216# 0.02fF
C37022 NOR2X1_LOC_770/a_36_216# INVX1_LOC_91/A 0.00fF
C37023 NOR2X1_LOC_655/B NOR2X1_LOC_9/Y 0.10fF
C37024 INVX1_LOC_41/Y INVX1_LOC_46/A 0.06fF
C37025 INVX1_LOC_64/A NOR2X1_LOC_755/Y -0.01fF
C37026 INVX1_LOC_145/A VDD -0.00fF
C37027 NAND2X1_LOC_357/B INVX1_LOC_91/A 0.23fF
C37028 INVX1_LOC_57/A NOR2X1_LOC_620/A 0.05fF
C37029 INVX1_LOC_64/A INVX1_LOC_284/A 0.09fF
C37030 INVX1_LOC_256/A INVX1_LOC_307/A 0.03fF
C37031 NOR2X1_LOC_738/Y NOR2X1_LOC_155/A 0.00fF
C37032 INVX1_LOC_27/A NOR2X1_LOC_721/B 0.02fF
C37033 NAND2X1_LOC_860/A INVX1_LOC_170/Y 0.04fF
C37034 NOR2X1_LOC_668/Y INVX1_LOC_4/Y 0.01fF
C37035 NOR2X1_LOC_208/Y VDD 1.99fF
C37036 INVX1_LOC_207/A NOR2X1_LOC_824/Y 0.04fF
C37037 NAND2X1_LOC_30/Y NAND2X1_LOC_50/a_36_24# 0.00fF
C37038 NOR2X1_LOC_552/A NOR2X1_LOC_337/a_36_216# 0.01fF
C37039 NOR2X1_LOC_71/Y INPUT_1 0.11fF
C37040 NOR2X1_LOC_184/a_36_216# INVX1_LOC_56/Y 0.00fF
C37041 INVX1_LOC_24/A NAND2X1_LOC_721/A 0.06fF
C37042 INVX1_LOC_217/A NOR2X1_LOC_536/A 0.03fF
C37043 NAND2X1_LOC_757/a_36_24# INVX1_LOC_12/Y 0.05fF
C37044 INVX1_LOC_1/A INVX1_LOC_84/A 0.58fF
C37045 NOR2X1_LOC_237/Y VDD 0.94fF
C37046 NAND2X1_LOC_357/B INVX1_LOC_11/Y 0.03fF
C37047 INVX1_LOC_69/Y NOR2X1_LOC_500/Y 0.15fF
C37048 NOR2X1_LOC_724/Y INVX1_LOC_85/Y 0.03fF
C37049 NOR2X1_LOC_788/a_36_216# NOR2X1_LOC_500/Y 0.00fF
C37050 INVX1_LOC_228/Y NOR2X1_LOC_649/B 0.01fF
C37051 NAND2X1_LOC_131/a_36_24# INVX1_LOC_84/A 0.00fF
C37052 INVX1_LOC_23/A INVX1_LOC_4/Y 0.27fF
C37053 INVX1_LOC_90/A NOR2X1_LOC_166/Y 0.01fF
C37054 INVX1_LOC_27/A NOR2X1_LOC_610/Y 0.06fF
C37055 NOR2X1_LOC_186/Y INVX1_LOC_42/A 0.10fF
C37056 NOR2X1_LOC_758/Y INVX1_LOC_46/A 0.04fF
C37057 NOR2X1_LOC_791/Y INVX1_LOC_168/Y 0.34fF
C37058 INVX1_LOC_33/A NOR2X1_LOC_706/B 0.03fF
C37059 NOR2X1_LOC_315/Y NOR2X1_LOC_92/a_36_216# 0.00fF
C37060 NOR2X1_LOC_773/Y NAND2X1_LOC_642/Y 0.07fF
C37061 INVX1_LOC_206/Y NOR2X1_LOC_577/a_36_216# 0.00fF
C37062 NOR2X1_LOC_309/Y VDD 1.99fF
C37063 INVX1_LOC_6/A NAND2X1_LOC_573/A 0.12fF
C37064 NAND2X1_LOC_325/Y INVX1_LOC_33/Y 0.17fF
C37065 NOR2X1_LOC_52/B NOR2X1_LOC_364/a_36_216# 0.00fF
C37066 INVX1_LOC_69/Y INVX1_LOC_10/A 0.03fF
C37067 NAND2X1_LOC_787/B NOR2X1_LOC_536/A 0.50fF
C37068 INVX1_LOC_6/A NOR2X1_LOC_528/a_36_216# 0.00fF
C37069 NOR2X1_LOC_574/A INVX1_LOC_37/A 0.03fF
C37070 NOR2X1_LOC_82/A NAND2X1_LOC_773/B 0.17fF
C37071 NAND2X1_LOC_573/Y INVX1_LOC_42/A 0.07fF
C37072 NAND2X1_LOC_338/B INVX1_LOC_20/A 0.14fF
C37073 NAND2X1_LOC_357/B NOR2X1_LOC_653/a_36_216# 0.00fF
C37074 NOR2X1_LOC_384/Y NOR2X1_LOC_88/Y 0.80fF
C37075 NAND2X1_LOC_451/Y INVX1_LOC_76/A 0.11fF
C37076 NOR2X1_LOC_278/a_36_216# INVX1_LOC_286/A 0.01fF
C37077 D_INPUT_0 INVX1_LOC_286/A 0.03fF
C37078 INVX1_LOC_289/A INVX1_LOC_187/Y 0.05fF
C37079 NOR2X1_LOC_248/Y INVX1_LOC_285/A 0.01fF
C37080 INVX1_LOC_272/Y NOR2X1_LOC_89/A 0.00fF
C37081 NOR2X1_LOC_561/Y NOR2X1_LOC_269/Y 0.04fF
C37082 NOR2X1_LOC_359/a_36_216# INVX1_LOC_290/Y 0.01fF
C37083 INVX1_LOC_196/A INVX1_LOC_37/A 0.03fF
C37084 INVX1_LOC_286/Y INVX1_LOC_63/A 0.00fF
C37085 INVX1_LOC_218/A INVX1_LOC_176/A 0.01fF
C37086 INVX1_LOC_85/A INVX1_LOC_44/A 0.03fF
C37087 NAND2X1_LOC_53/Y NOR2X1_LOC_89/A 0.72fF
C37088 INVX1_LOC_256/A INVX1_LOC_12/A 0.14fF
C37089 NOR2X1_LOC_156/B INVX1_LOC_117/A 0.03fF
C37090 INVX1_LOC_35/A INVX1_LOC_26/Y 1.17fF
C37091 NAND2X1_LOC_9/Y NOR2X1_LOC_720/A 0.02fF
C37092 INVX1_LOC_182/A NOR2X1_LOC_74/A 0.19fF
C37093 INVX1_LOC_58/A NOR2X1_LOC_125/Y 0.10fF
C37094 NOR2X1_LOC_384/Y INVX1_LOC_84/A 0.72fF
C37095 NOR2X1_LOC_553/Y NOR2X1_LOC_35/Y 0.01fF
C37096 NOR2X1_LOC_769/a_36_216# INVX1_LOC_37/A 0.00fF
C37097 NOR2X1_LOC_186/Y INVX1_LOC_78/A 0.19fF
C37098 NOR2X1_LOC_246/A NOR2X1_LOC_45/B 0.03fF
C37099 INVX1_LOC_1/A INVX1_LOC_15/A 0.35fF
C37100 NOR2X1_LOC_32/B INVX1_LOC_57/A 0.23fF
C37101 INVX1_LOC_250/A NOR2X1_LOC_605/A 0.07fF
C37102 INVX1_LOC_35/A INVX1_LOC_166/A 0.77fF
C37103 NOR2X1_LOC_748/a_36_216# INVX1_LOC_37/A 0.01fF
C37104 NAND2X1_LOC_208/B NAND2X1_LOC_74/B 0.01fF
C37105 NOR2X1_LOC_641/B NAND2X1_LOC_63/Y 0.02fF
C37106 NAND2X1_LOC_551/A NOR2X1_LOC_45/B 0.44fF
C37107 INVX1_LOC_36/A INVX1_LOC_133/A 1.82fF
C37108 NOR2X1_LOC_387/A NOR2X1_LOC_380/Y 0.74fF
C37109 INVX1_LOC_268/A INVX1_LOC_37/A 0.66fF
C37110 INVX1_LOC_213/Y INVX1_LOC_274/A 0.03fF
C37111 NOR2X1_LOC_123/B INVX1_LOC_304/A 0.00fF
C37112 NAND2X1_LOC_573/Y INVX1_LOC_78/A 0.07fF
C37113 NAND2X1_LOC_849/A INVX1_LOC_309/A 0.08fF
C37114 INVX1_LOC_136/A INVX1_LOC_49/Y 0.01fF
C37115 NOR2X1_LOC_664/Y NOR2X1_LOC_78/Y 0.54fF
C37116 NOR2X1_LOC_335/B NOR2X1_LOC_188/A 0.23fF
C37117 NOR2X1_LOC_65/B NOR2X1_LOC_186/Y 1.54fF
C37118 INVX1_LOC_289/A NAND2X1_LOC_446/a_36_24# 0.00fF
C37119 INVX1_LOC_58/A NAND2X1_LOC_715/B 0.03fF
C37120 NOR2X1_LOC_71/Y NAND2X1_LOC_455/a_36_24# 0.00fF
C37121 INVX1_LOC_299/A INVX1_LOC_18/Y 0.01fF
C37122 NOR2X1_LOC_321/a_36_216# INVX1_LOC_38/A 0.02fF
C37123 NOR2X1_LOC_216/Y NOR2X1_LOC_318/B 0.11fF
C37124 NAND2X1_LOC_849/A INVX1_LOC_91/A 0.06fF
C37125 NOR2X1_LOC_372/A INVX1_LOC_3/Y 0.00fF
C37126 NAND2X1_LOC_560/A NAND2X1_LOC_623/B 0.10fF
C37127 NOR2X1_LOC_837/B INVX1_LOC_19/A 0.27fF
C37128 INVX1_LOC_285/Y INVX1_LOC_6/A 0.17fF
C37129 INVX1_LOC_145/A INVX1_LOC_133/A 0.02fF
C37130 NOR2X1_LOC_627/a_36_216# INVX1_LOC_179/A 0.00fF
C37131 INVX1_LOC_299/A NAND2X1_LOC_256/a_36_24# 0.00fF
C37132 NOR2X1_LOC_183/a_36_216# INVX1_LOC_6/A 0.00fF
C37133 INVX1_LOC_193/Y NOR2X1_LOC_713/a_36_216# 0.00fF
C37134 INVX1_LOC_1/Y NOR2X1_LOC_16/a_36_216# 0.02fF
C37135 NOR2X1_LOC_207/A INVX1_LOC_113/A 0.03fF
C37136 INVX1_LOC_292/A NOR2X1_LOC_334/Y 0.02fF
C37137 NOR2X1_LOC_320/Y NOR2X1_LOC_45/B 0.01fF
C37138 INVX1_LOC_24/A NOR2X1_LOC_669/A 0.07fF
C37139 NOR2X1_LOC_790/A INVX1_LOC_23/A 0.01fF
C37140 NAND2X1_LOC_860/A INVX1_LOC_27/A 0.04fF
C37141 INVX1_LOC_31/A INVX1_LOC_4/Y 0.06fF
C37142 NAND2X1_LOC_860/A NOR2X1_LOC_824/A 0.67fF
C37143 INVX1_LOC_299/A NAND2X1_LOC_279/a_36_24# 0.00fF
C37144 NOR2X1_LOC_6/B NOR2X1_LOC_814/A 0.10fF
C37145 NAND2X1_LOC_834/a_36_24# INVX1_LOC_291/A 0.00fF
C37146 D_INPUT_1 INVX1_LOC_48/Y 0.03fF
C37147 NOR2X1_LOC_599/Y NOR2X1_LOC_409/B 0.46fF
C37148 NAND2X1_LOC_513/a_36_24# INVX1_LOC_274/A 0.00fF
C37149 NOR2X1_LOC_384/Y INVX1_LOC_15/A 0.07fF
C37150 INVX1_LOC_185/Y INVX1_LOC_63/A 0.01fF
C37151 NOR2X1_LOC_373/Y NAND2X1_LOC_848/A 0.29fF
C37152 D_GATE_222 NAND2X1_LOC_93/B -0.01fF
C37153 NOR2X1_LOC_620/Y INVX1_LOC_29/A 0.01fF
C37154 NAND2X1_LOC_660/Y INVX1_LOC_54/A 0.02fF
C37155 NAND2X1_LOC_738/B NAND2X1_LOC_303/Y 0.03fF
C37156 NOR2X1_LOC_798/A NOR2X1_LOC_211/Y 0.01fF
C37157 INVX1_LOC_72/A INVX1_LOC_4/A 0.10fF
C37158 INVX1_LOC_90/A NAND2X1_LOC_96/A 0.07fF
C37159 NOR2X1_LOC_100/A NAND2X1_LOC_206/Y -0.03fF
C37160 INVX1_LOC_305/A NAND2X1_LOC_278/a_36_24# 0.00fF
C37161 INVX1_LOC_34/A NAND2X1_LOC_74/B 0.14fF
C37162 D_GATE_222 NAND2X1_LOC_425/Y 0.02fF
C37163 NOR2X1_LOC_205/Y INVX1_LOC_23/A 0.08fF
C37164 INVX1_LOC_132/A INVX1_LOC_42/A 0.07fF
C37165 NAND2X1_LOC_23/a_36_24# NOR2X1_LOC_160/B 0.02fF
C37166 INVX1_LOC_181/Y INVX1_LOC_47/Y 0.06fF
C37167 NOR2X1_LOC_468/Y NOR2X1_LOC_717/A 0.02fF
C37168 INVX1_LOC_1/Y NOR2X1_LOC_197/B 0.31fF
C37169 INVX1_LOC_13/A NOR2X1_LOC_862/B 0.10fF
C37170 INVX1_LOC_278/A INVX1_LOC_1/A 0.10fF
C37171 INVX1_LOC_50/A NAND2X1_LOC_550/A 0.00fF
C37172 NOR2X1_LOC_2/Y NOR2X1_LOC_40/a_36_216# 0.00fF
C37173 NOR2X1_LOC_71/Y INVX1_LOC_118/A 0.28fF
C37174 D_INPUT_0 INVX1_LOC_54/A 0.03fF
C37175 NAND2X1_LOC_190/Y NOR2X1_LOC_717/A 0.14fF
C37176 NOR2X1_LOC_302/a_36_216# INVX1_LOC_179/A 0.00fF
C37177 NAND2X1_LOC_573/A INVX1_LOC_131/Y 0.03fF
C37178 NAND2X1_LOC_640/Y INVX1_LOC_42/A 0.02fF
C37179 INVX1_LOC_50/A NOR2X1_LOC_160/B 8.53fF
C37180 NAND2X1_LOC_214/B NAND2X1_LOC_473/A 0.01fF
C37181 NOR2X1_LOC_448/a_36_216# INVX1_LOC_295/Y 0.00fF
C37182 NOR2X1_LOC_166/Y INVX1_LOC_38/A 0.05fF
C37183 NOR2X1_LOC_798/A NOR2X1_LOC_440/B 0.01fF
C37184 INVX1_LOC_225/A INVX1_LOC_42/A 0.11fF
C37185 INVX1_LOC_70/Y NOR2X1_LOC_124/A 0.02fF
C37186 NOR2X1_LOC_74/A NOR2X1_LOC_176/Y 0.01fF
C37187 INVX1_LOC_58/A NOR2X1_LOC_372/A 0.03fF
C37188 INVX1_LOC_35/A INVX1_LOC_161/Y 0.07fF
C37189 NAND2X1_LOC_231/Y NAND2X1_LOC_74/B 0.04fF
C37190 INVX1_LOC_27/A NAND2X1_LOC_473/A 0.07fF
C37191 INVX1_LOC_171/A NOR2X1_LOC_79/a_36_216# 0.00fF
C37192 INVX1_LOC_286/A NOR2X1_LOC_266/B 0.03fF
C37193 INPUT_1 NAND2X1_LOC_243/Y 0.00fF
C37194 NAND2X1_LOC_544/a_36_24# NAND2X1_LOC_550/A 0.00fF
C37195 INVX1_LOC_190/Y NOR2X1_LOC_435/A 0.01fF
C37196 INVX1_LOC_89/Y INPUT_1 0.01fF
C37197 NOR2X1_LOC_174/B NOR2X1_LOC_862/B 0.05fF
C37198 NOR2X1_LOC_99/B NOR2X1_LOC_865/Y 0.06fF
C37199 NOR2X1_LOC_269/Y INVX1_LOC_76/A 0.19fF
C37200 NOR2X1_LOC_99/B NOR2X1_LOC_243/B 0.05fF
C37201 NAND2X1_LOC_339/a_36_24# INVX1_LOC_32/A 0.00fF
C37202 INVX1_LOC_132/A INVX1_LOC_78/A 0.07fF
C37203 INVX1_LOC_67/A NOR2X1_LOC_334/Y 0.03fF
C37204 INVX1_LOC_33/A INVX1_LOC_94/Y 0.07fF
C37205 INVX1_LOC_22/A INVX1_LOC_272/A 0.08fF
C37206 INVX1_LOC_64/A NOR2X1_LOC_348/a_36_216# 0.01fF
C37207 NOR2X1_LOC_336/B INVX1_LOC_58/Y 0.22fF
C37208 INVX1_LOC_75/A NOR2X1_LOC_612/Y 0.01fF
C37209 INVX1_LOC_89/A NAND2X1_LOC_73/a_36_24# 0.00fF
C37210 INVX1_LOC_64/A NOR2X1_LOC_361/a_36_216# 0.00fF
C37211 INVX1_LOC_35/A INVX1_LOC_312/A 0.01fF
C37212 NOR2X1_LOC_557/Y INVX1_LOC_87/A 0.08fF
C37213 INVX1_LOC_11/A NAND2X1_LOC_474/Y 0.07fF
C37214 NAND2X1_LOC_808/A NOR2X1_LOC_661/A 0.01fF
C37215 INVX1_LOC_95/A NOR2X1_LOC_266/B 0.00fF
C37216 NOR2X1_LOC_838/a_36_216# INVX1_LOC_26/Y 0.00fF
C37217 NOR2X1_LOC_561/Y NOR2X1_LOC_36/B 0.18fF
C37218 NAND2X1_LOC_390/A INVX1_LOC_29/A 0.04fF
C37219 INVX1_LOC_303/A NOR2X1_LOC_843/B 0.07fF
C37220 NAND2X1_LOC_9/Y NOR2X1_LOC_410/Y 0.01fF
C37221 NOR2X1_LOC_590/A INVX1_LOC_50/Y 0.78fF
C37222 INVX1_LOC_225/A INVX1_LOC_78/A 0.54fF
C37223 INVX1_LOC_306/A NAND2X1_LOC_773/B 0.14fF
C37224 NOR2X1_LOC_329/B NOR2X1_LOC_841/A 0.51fF
C37225 NAND2X1_LOC_35/Y INVX1_LOC_30/A 0.09fF
C37226 INVX1_LOC_132/A NOR2X1_LOC_65/B 0.10fF
C37227 INVX1_LOC_64/A INVX1_LOC_72/A 0.25fF
C37228 INVX1_LOC_89/A NOR2X1_LOC_257/Y 0.01fF
C37229 NOR2X1_LOC_440/Y INVX1_LOC_12/A 0.94fF
C37230 NAND2X1_LOC_338/B INVX1_LOC_4/A 0.07fF
C37231 INVX1_LOC_55/A NAND2X1_LOC_149/Y 0.02fF
C37232 NOR2X1_LOC_533/Y NAND2X1_LOC_538/Y 0.12fF
C37233 NOR2X1_LOC_71/Y NAND2X1_LOC_63/Y 0.43fF
C37234 INVX1_LOC_10/A NOR2X1_LOC_89/A 0.10fF
C37235 NOR2X1_LOC_724/Y NAND2X1_LOC_782/B 0.02fF
C37236 NOR2X1_LOC_596/A NOR2X1_LOC_717/A 0.08fF
C37237 NAND2X1_LOC_151/a_36_24# NAND2X1_LOC_537/Y 0.01fF
C37238 NOR2X1_LOC_392/B NAND2X1_LOC_99/A 0.10fF
C37239 INVX1_LOC_246/A NAND2X1_LOC_175/a_36_24# 0.01fF
C37240 INVX1_LOC_83/A INVX1_LOC_69/A 0.04fF
C37241 INVX1_LOC_233/A INVX1_LOC_41/Y 0.08fF
C37242 NOR2X1_LOC_510/Y INVX1_LOC_36/A 0.03fF
C37243 NOR2X1_LOC_305/Y INVX1_LOC_37/A 0.07fF
C37244 NOR2X1_LOC_614/Y NOR2X1_LOC_623/B 0.06fF
C37245 NAND2X1_LOC_552/A NOR2X1_LOC_91/Y 0.33fF
C37246 NOR2X1_LOC_65/B INVX1_LOC_225/A 0.15fF
C37247 INVX1_LOC_155/Y INVX1_LOC_57/A 0.00fF
C37248 INVX1_LOC_143/A INVX1_LOC_87/A 0.36fF
C37249 INVX1_LOC_60/A NOR2X1_LOC_39/Y 0.01fF
C37250 NAND2X1_LOC_53/Y INVX1_LOC_11/A 0.10fF
C37251 INVX1_LOC_266/A NOR2X1_LOC_590/A 0.31fF
C37252 INVX1_LOC_75/A NOR2X1_LOC_673/A 0.03fF
C37253 INVX1_LOC_69/Y NOR2X1_LOC_445/B 0.07fF
C37254 NOR2X1_LOC_227/B INVX1_LOC_210/Y 0.01fF
C37255 NOR2X1_LOC_332/B INVX1_LOC_280/A 0.00fF
C37256 NOR2X1_LOC_71/Y NAND2X1_LOC_455/B 0.16fF
C37257 NOR2X1_LOC_720/B INVX1_LOC_57/A 0.01fF
C37258 NOR2X1_LOC_357/Y INVX1_LOC_281/A 0.02fF
C37259 NOR2X1_LOC_389/a_36_216# NAND2X1_LOC_807/B 0.00fF
C37260 INVX1_LOC_58/A NAND2X1_LOC_308/Y 0.03fF
C37261 INVX1_LOC_255/Y NAND2X1_LOC_618/Y 0.02fF
C37262 INVX1_LOC_2/A NOR2X1_LOC_39/Y 0.10fF
C37263 NOR2X1_LOC_67/A INVX1_LOC_23/Y 0.05fF
C37264 INVX1_LOC_178/A NOR2X1_LOC_91/Y 0.01fF
C37265 NOR2X1_LOC_188/A INVX1_LOC_84/A 0.14fF
C37266 INVX1_LOC_177/A INVX1_LOC_270/A 0.03fF
C37267 NOR2X1_LOC_45/B INVX1_LOC_260/A 0.02fF
C37268 NOR2X1_LOC_91/A NOR2X1_LOC_526/Y 0.03fF
C37269 NOR2X1_LOC_689/Y NAND2X1_LOC_353/a_36_24# 0.00fF
C37270 NOR2X1_LOC_15/Y NOR2X1_LOC_266/a_36_216# 0.00fF
C37271 NOR2X1_LOC_295/Y NOR2X1_LOC_717/A 0.01fF
C37272 VDD NOR2X1_LOC_865/A 0.12fF
C37273 INVX1_LOC_36/A NOR2X1_LOC_361/B 0.03fF
C37274 D_INPUT_1 NOR2X1_LOC_84/Y 0.20fF
C37275 NOR2X1_LOC_19/B NOR2X1_LOC_610/Y 0.02fF
C37276 NAND2X1_LOC_591/a_36_24# INVX1_LOC_1/A 0.00fF
C37277 D_INPUT_4 INPUT_7 0.04fF
C37278 NOR2X1_LOC_91/A NAND2X1_LOC_862/A 0.01fF
C37279 NOR2X1_LOC_56/Y NOR2X1_LOC_435/A -0.00fF
C37280 INVX1_LOC_269/A NOR2X1_LOC_791/B 0.01fF
C37281 NOR2X1_LOC_267/A NOR2X1_LOC_361/B 1.34fF
C37282 NOR2X1_LOC_78/B INVX1_LOC_270/Y 3.57fF
C37283 NOR2X1_LOC_751/A NAND2X1_LOC_63/Y 0.10fF
C37284 INVX1_LOC_88/A INVX1_LOC_18/A 0.17fF
C37285 INVX1_LOC_99/Y NOR2X1_LOC_254/Y 0.26fF
C37286 NOR2X1_LOC_656/a_36_216# INVX1_LOC_14/A 0.03fF
C37287 VDD NOR2X1_LOC_656/Y 0.12fF
C37288 NAND2X1_LOC_802/A NAND2X1_LOC_714/B 0.05fF
C37289 NAND2X1_LOC_798/a_36_24# INVX1_LOC_178/A 0.06fF
C37290 NOR2X1_LOC_433/A NAND2X1_LOC_474/Y 0.01fF
C37291 NAND2X1_LOC_96/A INVX1_LOC_38/A 0.07fF
C37292 INPUT_0 NAND2X1_LOC_74/B 5.36fF
C37293 NOR2X1_LOC_322/Y INVX1_LOC_102/A 0.10fF
C37294 INVX1_LOC_289/Y INVX1_LOC_24/A 0.03fF
C37295 NOR2X1_LOC_272/Y NOR2X1_LOC_716/B 0.10fF
C37296 INVX1_LOC_166/A INVX1_LOC_84/Y 0.05fF
C37297 INVX1_LOC_50/A INVX1_LOC_208/A 0.09fF
C37298 INVX1_LOC_45/A INVX1_LOC_174/A 0.03fF
C37299 NAND2X1_LOC_213/A NAND2X1_LOC_162/B 0.01fF
C37300 INVX1_LOC_37/A NAND2X1_LOC_289/a_36_24# 0.00fF
C37301 INVX1_LOC_282/A INVX1_LOC_284/A 0.18fF
C37302 INVX1_LOC_313/Y INVX1_LOC_4/A 0.07fF
C37303 NAND2X1_LOC_284/a_36_24# INVX1_LOC_118/A 0.00fF
C37304 NOR2X1_LOC_658/Y NOR2X1_LOC_389/A 0.10fF
C37305 INVX1_LOC_35/A NAND2X1_LOC_335/a_36_24# 0.00fF
C37306 NOR2X1_LOC_561/Y INVX1_LOC_26/A 0.00fF
C37307 INVX1_LOC_6/A NAND2X1_LOC_81/B 0.03fF
C37308 NOR2X1_LOC_45/B NAND2X1_LOC_489/Y 0.07fF
C37309 NOR2X1_LOC_361/B INVX1_LOC_145/A 0.02fF
C37310 INVX1_LOC_21/A NOR2X1_LOC_388/Y 0.02fF
C37311 NAND2X1_LOC_84/Y INVX1_LOC_14/A 0.13fF
C37312 INVX1_LOC_96/Y NOR2X1_LOC_665/Y 0.29fF
C37313 VDD NOR2X1_LOC_435/A -0.00fF
C37314 INVX1_LOC_43/Y INVX1_LOC_72/A 0.29fF
C37315 NAND2X1_LOC_35/Y NAND2X1_LOC_722/A 0.07fF
C37316 NOR2X1_LOC_516/B NOR2X1_LOC_105/Y 0.04fF
C37317 INPUT_0 NOR2X1_LOC_847/B 0.09fF
C37318 NAND2X1_LOC_724/A NOR2X1_LOC_152/Y 0.09fF
C37319 INVX1_LOC_136/A INVX1_LOC_161/A 0.51fF
C37320 INVX1_LOC_64/A NAND2X1_LOC_338/B 0.34fF
C37321 INVX1_LOC_69/Y INVX1_LOC_12/A 0.15fF
C37322 INVX1_LOC_14/Y INVX1_LOC_179/A 0.03fF
C37323 INVX1_LOC_27/A NOR2X1_LOC_516/Y 0.03fF
C37324 NOR2X1_LOC_74/A NOR2X1_LOC_850/B 0.11fF
C37325 NOR2X1_LOC_82/A INVX1_LOC_24/A 0.07fF
C37326 INVX1_LOC_47/A NAND2X1_LOC_72/B 0.03fF
C37327 NOR2X1_LOC_457/A INVX1_LOC_94/A 0.07fF
C37328 NAND2X1_LOC_794/B NOR2X1_LOC_591/Y 0.05fF
C37329 D_INPUT_0 NOR2X1_LOC_438/Y 0.04fF
C37330 NAND2X1_LOC_848/A INVX1_LOC_54/A 0.02fF
C37331 NAND2X1_LOC_21/Y INVX1_LOC_1/A 0.06fF
C37332 NOR2X1_LOC_52/B NAND2X1_LOC_474/Y 0.07fF
C37333 NAND2X1_LOC_639/A INVX1_LOC_92/A 0.10fF
C37334 NOR2X1_LOC_56/Y INVX1_LOC_63/A 0.01fF
C37335 INVX1_LOC_272/Y NOR2X1_LOC_433/A 0.01fF
C37336 INVX1_LOC_299/A INVX1_LOC_33/A 0.11fF
C37337 INVX1_LOC_13/Y INVX1_LOC_34/Y 0.03fF
C37338 INVX1_LOC_103/A INVX1_LOC_209/Y 0.20fF
C37339 NOR2X1_LOC_231/a_36_216# NAND2X1_LOC_364/A 0.00fF
C37340 NOR2X1_LOC_634/A INVX1_LOC_117/A 0.02fF
C37341 INVX1_LOC_16/A NOR2X1_LOC_678/A 0.07fF
C37342 NOR2X1_LOC_585/a_36_216# INVX1_LOC_72/A 0.00fF
C37343 NOR2X1_LOC_798/A NOR2X1_LOC_538/Y 0.01fF
C37344 NAND2X1_LOC_53/Y NOR2X1_LOC_433/A 0.16fF
C37345 INVX1_LOC_174/A INVX1_LOC_71/A 0.03fF
C37346 INVX1_LOC_215/Y NOR2X1_LOC_513/a_36_216# 0.00fF
C37347 NOR2X1_LOC_536/A INVX1_LOC_92/A 0.26fF
C37348 INVX1_LOC_176/A NAND2X1_LOC_206/Y 0.02fF
C37349 NAND2X1_LOC_708/Y INVX1_LOC_22/A 0.04fF
C37350 NOR2X1_LOC_790/B NOR2X1_LOC_553/B 0.42fF
C37351 INVX1_LOC_65/A NOR2X1_LOC_633/A 0.03fF
C37352 INVX1_LOC_43/A INVX1_LOC_306/Y 0.23fF
C37353 D_INPUT_0 NAND2X1_LOC_215/A 0.08fF
C37354 NAND2X1_LOC_53/Y NOR2X1_LOC_593/Y 0.02fF
C37355 INVX1_LOC_10/A NAND2X1_LOC_804/A 0.12fF
C37356 NOR2X1_LOC_361/B NOR2X1_LOC_309/Y 0.08fF
C37357 NAND2X1_LOC_193/a_36_24# NOR2X1_LOC_45/Y 0.01fF
C37358 INVX1_LOC_28/A NOR2X1_LOC_318/A 0.01fF
C37359 VDD INVX1_LOC_63/A 2.53fF
C37360 INVX1_LOC_130/Y INVX1_LOC_72/A 0.03fF
C37361 NOR2X1_LOC_759/A NOR2X1_LOC_52/Y 0.05fF
C37362 NOR2X1_LOC_791/Y INVX1_LOC_56/A 0.01fF
C37363 NAND2X1_LOC_128/a_36_24# INVX1_LOC_271/A 0.00fF
C37364 INVX1_LOC_14/A NOR2X1_LOC_612/B 0.45fF
C37365 NAND2X1_LOC_642/Y INVX1_LOC_42/A 0.16fF
C37366 INPUT_1 NAND2X1_LOC_205/A 0.50fF
C37367 INVX1_LOC_216/Y NAND2X1_LOC_563/Y 0.03fF
C37368 INVX1_LOC_17/A INVX1_LOC_119/A 0.17fF
C37369 NAND2X1_LOC_665/a_36_24# NAND2X1_LOC_215/A 0.00fF
C37370 INVX1_LOC_6/A INVX1_LOC_4/Y 0.18fF
C37371 NAND2X1_LOC_53/Y NOR2X1_LOC_52/B 0.02fF
C37372 NOR2X1_LOC_45/B INVX1_LOC_32/A 0.03fF
C37373 NOR2X1_LOC_468/Y INVX1_LOC_256/Y 0.00fF
C37374 NAND2X1_LOC_93/B INVX1_LOC_92/A 0.06fF
C37375 INVX1_LOC_105/A NAND2X1_LOC_195/Y 0.39fF
C37376 NOR2X1_LOC_68/A INVX1_LOC_314/Y 0.07fF
C37377 NOR2X1_LOC_817/Y NOR2X1_LOC_818/Y 0.17fF
C37378 NOR2X1_LOC_524/Y INVX1_LOC_33/A 0.01fF
C37379 NOR2X1_LOC_45/B NOR2X1_LOC_329/Y 0.01fF
C37380 NOR2X1_LOC_465/a_36_216# INVX1_LOC_313/Y 0.00fF
C37381 NOR2X1_LOC_590/A NOR2X1_LOC_6/B 0.05fF
C37382 INVX1_LOC_233/Y NAND2X1_LOC_866/B 0.10fF
C37383 NOR2X1_LOC_458/Y INVX1_LOC_36/A 0.02fF
C37384 INVX1_LOC_36/A INVX1_LOC_153/Y 0.01fF
C37385 INVX1_LOC_64/A INVX1_LOC_313/Y 0.35fF
C37386 INVX1_LOC_247/A INVX1_LOC_32/A 0.03fF
C37387 INVX1_LOC_28/A NOR2X1_LOC_678/A 0.00fF
C37388 INVX1_LOC_117/A INVX1_LOC_29/A 0.39fF
C37389 INVX1_LOC_267/A NAND2X1_LOC_555/Y 0.02fF
C37390 INVX1_LOC_136/A INVX1_LOC_34/A 7.30fF
C37391 INVX1_LOC_30/A NAND2X1_LOC_465/Y 0.05fF
C37392 NAND2X1_LOC_59/B INVX1_LOC_18/A 0.01fF
C37393 NAND2X1_LOC_338/B INVX1_LOC_43/Y 0.04fF
C37394 INVX1_LOC_21/A INVX1_LOC_135/A 0.11fF
C37395 INVX1_LOC_201/Y NOR2X1_LOC_476/Y 0.00fF
C37396 INVX1_LOC_11/A NOR2X1_LOC_500/Y 0.07fF
C37397 NOR2X1_LOC_45/B NAND2X1_LOC_175/Y 0.07fF
C37398 NOR2X1_LOC_846/a_36_216# INVX1_LOC_63/A 0.01fF
C37399 INVX1_LOC_226/Y INVX1_LOC_11/A 0.29fF
C37400 INVX1_LOC_285/Y INVX1_LOC_270/A 0.10fF
C37401 NOR2X1_LOC_682/Y NOR2X1_LOC_48/B 0.04fF
C37402 INVX1_LOC_78/A NAND2X1_LOC_642/Y 0.13fF
C37403 INVX1_LOC_266/A INVX1_LOC_227/A 0.21fF
C37404 NOR2X1_LOC_657/B NAND2X1_LOC_454/Y 0.03fF
C37405 NAND2X1_LOC_350/A NAND2X1_LOC_319/a_36_24# 0.01fF
C37406 NAND2X1_LOC_545/a_36_24# NOR2X1_LOC_52/B 0.00fF
C37407 INVX1_LOC_300/Y NAND2X1_LOC_811/Y 0.03fF
C37408 NOR2X1_LOC_155/A NAND2X1_LOC_475/Y 0.00fF
C37409 NOR2X1_LOC_208/Y INVX1_LOC_153/Y 0.10fF
C37410 INVX1_LOC_108/Y NOR2X1_LOC_188/A 0.00fF
C37411 INPUT_0 NOR2X1_LOC_660/Y 0.66fF
C37412 NOR2X1_LOC_91/A NOR2X1_LOC_595/Y 0.21fF
C37413 NOR2X1_LOC_453/Y INVX1_LOC_295/A 0.02fF
C37414 NOR2X1_LOC_196/Y INVX1_LOC_68/A 0.01fF
C37415 INVX1_LOC_25/A INVX1_LOC_123/A 0.15fF
C37416 INVX1_LOC_42/A NOR2X1_LOC_271/Y 0.02fF
C37417 INVX1_LOC_136/A NAND2X1_LOC_231/Y 0.10fF
C37418 INVX1_LOC_36/A INVX1_LOC_280/Y 0.03fF
C37419 NAND2X1_LOC_350/A NAND2X1_LOC_660/Y 0.07fF
C37420 INVX1_LOC_11/A INVX1_LOC_10/A 0.08fF
C37421 NOR2X1_LOC_65/B NAND2X1_LOC_642/Y 0.10fF
C37422 NOR2X1_LOC_334/Y NOR2X1_LOC_137/Y 0.02fF
C37423 INVX1_LOC_49/A NOR2X1_LOC_570/B 0.01fF
C37424 VDD NAND2X1_LOC_452/Y 0.22fF
C37425 NOR2X1_LOC_390/a_36_216# INVX1_LOC_77/A 0.00fF
C37426 INVX1_LOC_17/A INVX1_LOC_150/A 0.01fF
C37427 INVX1_LOC_292/A NOR2X1_LOC_569/Y 0.67fF
C37428 NOR2X1_LOC_34/Y NOR2X1_LOC_35/Y 0.03fF
C37429 INVX1_LOC_237/Y INVX1_LOC_207/A 0.14fF
C37430 NOR2X1_LOC_273/Y INVX1_LOC_266/Y 0.01fF
C37431 INVX1_LOC_269/A NOR2X1_LOC_532/Y 0.01fF
C37432 NOR2X1_LOC_778/B NOR2X1_LOC_68/A 0.01fF
C37433 INVX1_LOC_37/A INVX1_LOC_271/Y 0.07fF
C37434 NOR2X1_LOC_403/B NOR2X1_LOC_84/Y 0.05fF
C37435 NOR2X1_LOC_82/A NOR2X1_LOC_130/A 0.09fF
C37436 NOR2X1_LOC_219/B INVX1_LOC_63/Y 0.02fF
C37437 INVX1_LOC_17/A INVX1_LOC_89/A 0.03fF
C37438 NOR2X1_LOC_264/Y NAND2X1_LOC_361/Y 0.17fF
C37439 VDD NOR2X1_LOC_307/Y 0.24fF
C37440 INVX1_LOC_26/A INVX1_LOC_76/A 0.07fF
C37441 INVX1_LOC_136/A NOR2X1_LOC_772/a_36_216# 0.01fF
C37442 NOR2X1_LOC_137/B INVX1_LOC_270/A 0.01fF
C37443 NOR2X1_LOC_89/A INVX1_LOC_307/A 0.04fF
C37444 NAND2X1_LOC_806/a_36_24# NOR2X1_LOC_743/Y 0.00fF
C37445 INVX1_LOC_54/Y NOR2X1_LOC_303/Y 0.03fF
C37446 INVX1_LOC_282/A NOR2X1_LOC_384/A 0.15fF
C37447 INVX1_LOC_45/A NOR2X1_LOC_589/A 8.20fF
C37448 NOR2X1_LOC_303/Y NOR2X1_LOC_353/Y 0.02fF
C37449 NOR2X1_LOC_134/Y NOR2X1_LOC_373/Y 0.06fF
C37450 VDD NAND2X1_LOC_223/B 0.01fF
C37451 NOR2X1_LOC_817/Y INPUT_1 0.04fF
C37452 NAND2X1_LOC_96/A NAND2X1_LOC_223/A 0.42fF
C37453 INVX1_LOC_33/A NOR2X1_LOC_315/Y 0.10fF
C37454 INVX1_LOC_17/A NAND2X1_LOC_508/A 0.07fF
C37455 NOR2X1_LOC_471/Y INVX1_LOC_89/A 0.03fF
C37456 NAND2X1_LOC_785/A NOR2X1_LOC_716/B 0.02fF
C37457 D_INPUT_0 INVX1_LOC_218/Y 0.03fF
C37458 INVX1_LOC_239/A NAND2X1_LOC_463/B 0.00fF
C37459 NOR2X1_LOC_405/A INVX1_LOC_58/Y 0.13fF
C37460 INVX1_LOC_224/Y INVX1_LOC_20/A 0.03fF
C37461 NOR2X1_LOC_78/A NAND2X1_LOC_248/a_36_24# 0.01fF
C37462 VDD NOR2X1_LOC_65/Y 0.49fF
C37463 NOR2X1_LOC_804/B INVX1_LOC_177/A 0.08fF
C37464 D_INPUT_0 NOR2X1_LOC_441/Y 0.04fF
C37465 INVX1_LOC_298/Y INVX1_LOC_117/A 0.03fF
C37466 NOR2X1_LOC_406/a_36_216# INVX1_LOC_91/A 0.00fF
C37467 INVX1_LOC_36/A NAND2X1_LOC_573/A 0.01fF
C37468 NAND2X1_LOC_555/Y INVX1_LOC_89/A 0.22fF
C37469 NAND2X1_LOC_350/B INVX1_LOC_105/A 0.01fF
C37470 INVX1_LOC_50/A NAND2X1_LOC_211/Y 0.04fF
C37471 INVX1_LOC_11/A NOR2X1_LOC_302/Y 0.04fF
C37472 NAND2X1_LOC_579/A NOR2X1_LOC_74/A 0.15fF
C37473 NOR2X1_LOC_474/A INVX1_LOC_197/A 0.15fF
C37474 INVX1_LOC_133/A INVX1_LOC_63/A 0.02fF
C37475 NOR2X1_LOC_255/Y INVX1_LOC_76/A 0.33fF
C37476 INVX1_LOC_270/Y INVX1_LOC_46/A 0.01fF
C37477 INVX1_LOC_310/Y INVX1_LOC_196/A 0.15fF
C37478 NOR2X1_LOC_191/B INVX1_LOC_1/Y 0.98fF
C37479 NOR2X1_LOC_267/A NAND2X1_LOC_573/A 0.05fF
C37480 NOR2X1_LOC_706/B INVX1_LOC_275/Y 0.02fF
C37481 INVX1_LOC_36/A NAND2X1_LOC_143/a_36_24# 0.00fF
C37482 NOR2X1_LOC_276/B NOR2X1_LOC_561/Y 0.01fF
C37483 INVX1_LOC_249/Y INVX1_LOC_266/Y 0.01fF
C37484 INVX1_LOC_45/A INVX1_LOC_171/A 0.01fF
C37485 NAND2X1_LOC_848/A NOR2X1_LOC_438/Y 0.02fF
C37486 NOR2X1_LOC_35/Y NOR2X1_LOC_678/A 0.05fF
C37487 INVX1_LOC_90/A NAND2X1_LOC_577/A 3.57fF
C37488 NOR2X1_LOC_170/A NOR2X1_LOC_445/B 0.03fF
C37489 INVX1_LOC_20/A NAND2X1_LOC_793/B 0.04fF
C37490 INVX1_LOC_171/A NOR2X1_LOC_568/A 0.00fF
C37491 NOR2X1_LOC_267/a_36_216# INVX1_LOC_126/Y 0.01fF
C37492 INVX1_LOC_204/A INVX1_LOC_117/A 0.04fF
C37493 NOR2X1_LOC_589/A INVX1_LOC_71/A 0.69fF
C37494 INVX1_LOC_46/A NOR2X1_LOC_754/Y 0.01fF
C37495 NAND2X1_LOC_773/a_36_24# NOR2X1_LOC_271/Y 0.00fF
C37496 NOR2X1_LOC_593/Y NOR2X1_LOC_500/Y 0.07fF
C37497 NAND2X1_LOC_181/Y INVX1_LOC_8/A 0.02fF
C37498 INVX1_LOC_223/A NOR2X1_LOC_473/B 0.05fF
C37499 NAND2X1_LOC_79/Y NOR2X1_LOC_719/B 0.22fF
C37500 INVX1_LOC_21/A NOR2X1_LOC_552/A 0.06fF
C37501 INVX1_LOC_14/A INVX1_LOC_48/A 0.07fF
C37502 NOR2X1_LOC_205/Y INVX1_LOC_6/A 0.31fF
C37503 NAND2X1_LOC_470/B INVX1_LOC_92/A 0.02fF
C37504 NAND2X1_LOC_563/A NOR2X1_LOC_124/B 0.03fF
C37505 INVX1_LOC_277/A INVX1_LOC_311/Y 0.15fF
C37506 INVX1_LOC_215/A INVX1_LOC_49/A 0.09fF
C37507 NAND2X1_LOC_254/Y NAND2X1_LOC_768/Y 0.01fF
C37508 INVX1_LOC_24/A INVX1_LOC_306/A 0.01fF
C37509 NOR2X1_LOC_541/Y INVX1_LOC_222/A 0.01fF
C37510 INVX1_LOC_34/A NOR2X1_LOC_701/Y 0.04fF
C37511 NOR2X1_LOC_770/B INVX1_LOC_22/A 0.48fF
C37512 NOR2X1_LOC_68/A NOR2X1_LOC_724/Y 0.12fF
C37513 NOR2X1_LOC_433/A INVX1_LOC_10/A 0.14fF
C37514 NOR2X1_LOC_276/Y INPUT_0 0.10fF
C37515 INVX1_LOC_219/Y INVX1_LOC_316/Y 0.01fF
C37516 NAND2X1_LOC_361/Y INVX1_LOC_160/Y 0.12fF
C37517 NAND2X1_LOC_562/Y INVX1_LOC_255/Y 0.03fF
C37518 INVX1_LOC_226/Y NOR2X1_LOC_52/B 0.01fF
C37519 INVX1_LOC_171/A INVX1_LOC_71/A 0.01fF
C37520 NOR2X1_LOC_703/B NOR2X1_LOC_564/Y 0.05fF
C37521 INVX1_LOC_53/A NOR2X1_LOC_536/A 0.06fF
C37522 NOR2X1_LOC_89/A INVX1_LOC_12/A 0.06fF
C37523 INVX1_LOC_90/A NAND2X1_LOC_656/A 0.02fF
C37524 NOR2X1_LOC_209/Y NOR2X1_LOC_307/B 0.43fF
C37525 INVX1_LOC_31/Y NOR2X1_LOC_500/B 0.05fF
C37526 NOR2X1_LOC_389/B NAND2X1_LOC_656/A 0.26fF
C37527 INVX1_LOC_30/A INVX1_LOC_144/A 0.07fF
C37528 NOR2X1_LOC_504/Y NAND2X1_LOC_863/B 0.08fF
C37529 NOR2X1_LOC_91/Y INVX1_LOC_140/A 0.14fF
C37530 INVX1_LOC_72/A INVX1_LOC_282/A 0.07fF
C37531 INVX1_LOC_45/A INVX1_LOC_222/A 0.01fF
C37532 D_INPUT_0 NOR2X1_LOC_340/Y 0.00fF
C37533 NOR2X1_LOC_309/Y NAND2X1_LOC_573/A 0.10fF
C37534 NAND2X1_LOC_640/Y NAND2X1_LOC_861/Y 0.03fF
C37535 INVX1_LOC_3/Y INVX1_LOC_29/A 0.08fF
C37536 INVX1_LOC_222/A NOR2X1_LOC_568/A 0.01fF
C37537 NOR2X1_LOC_67/A INVX1_LOC_232/A 0.10fF
C37538 INVX1_LOC_136/A INPUT_0 0.39fF
C37539 NOR2X1_LOC_52/B INVX1_LOC_10/A 0.26fF
C37540 INVX1_LOC_2/A INVX1_LOC_215/A 0.15fF
C37541 INVX1_LOC_36/A INVX1_LOC_285/Y 0.03fF
C37542 INVX1_LOC_46/Y NAND2X1_LOC_215/A 0.21fF
C37543 NOR2X1_LOC_590/A INVX1_LOC_96/A 0.04fF
C37544 NAND2X1_LOC_53/Y INVX1_LOC_199/A 0.12fF
C37545 NOR2X1_LOC_723/Y INVX1_LOC_6/A 0.01fF
C37546 D_INPUT_6 NAND2X1_LOC_51/a_36_24# 0.00fF
C37547 INVX1_LOC_21/A NOR2X1_LOC_813/Y 0.07fF
C37548 NAND2X1_LOC_348/A NAND2X1_LOC_656/A 0.03fF
C37549 NOR2X1_LOC_15/Y NOR2X1_LOC_562/A 0.03fF
C37550 NOR2X1_LOC_335/A INVX1_LOC_28/A 0.04fF
C37551 INVX1_LOC_64/A NOR2X1_LOC_506/Y 0.00fF
C37552 INVX1_LOC_53/A NAND2X1_LOC_93/B 0.36fF
C37553 INVX1_LOC_233/A INVX1_LOC_185/A 0.01fF
C37554 INVX1_LOC_279/Y NOR2X1_LOC_78/A 0.01fF
C37555 INVX1_LOC_21/A NOR2X1_LOC_152/A 0.01fF
C37556 INVX1_LOC_36/A NOR2X1_LOC_183/a_36_216# -0.00fF
C37557 INVX1_LOC_35/A INVX1_LOC_108/A 0.02fF
C37558 NOR2X1_LOC_647/A NOR2X1_LOC_820/B 0.24fF
C37559 NAND2X1_LOC_784/A NOR2X1_LOC_88/Y 0.05fF
C37560 INVX1_LOC_17/A NAND2X1_LOC_244/A 0.02fF
C37561 NOR2X1_LOC_172/Y NOR2X1_LOC_329/B 0.03fF
C37562 NOR2X1_LOC_103/Y INVX1_LOC_20/A 0.07fF
C37563 INVX1_LOC_209/Y NOR2X1_LOC_597/a_36_216# 0.00fF
C37564 INVX1_LOC_223/A NOR2X1_LOC_355/B 0.09fF
C37565 INVX1_LOC_303/A INVX1_LOC_31/Y 0.03fF
C37566 NOR2X1_LOC_168/Y NOR2X1_LOC_548/B 0.35fF
C37567 INVX1_LOC_222/Y INVX1_LOC_38/A 0.03fF
C37568 NAND2X1_LOC_860/A NOR2X1_LOC_216/B 0.03fF
C37569 INVX1_LOC_45/A NOR2X1_LOC_311/a_36_216# 0.00fF
C37570 INVX1_LOC_21/A INVX1_LOC_280/A 0.19fF
C37571 INVX1_LOC_53/A NAND2X1_LOC_425/Y 0.20fF
C37572 NOR2X1_LOC_742/A INVX1_LOC_283/Y -0.06fF
C37573 INVX1_LOC_21/A NOR2X1_LOC_94/Y 0.06fF
C37574 INVX1_LOC_89/A NOR2X1_LOC_507/a_36_216# 0.00fF
C37575 INVX1_LOC_30/Y NOR2X1_LOC_82/Y 0.10fF
C37576 NOR2X1_LOC_655/B D_INPUT_0 0.03fF
C37577 INVX1_LOC_214/A INVX1_LOC_135/A 0.10fF
C37578 INVX1_LOC_130/A NOR2X1_LOC_275/A 0.00fF
C37579 NOR2X1_LOC_19/B NOR2X1_LOC_516/Y 0.00fF
C37580 NOR2X1_LOC_667/A INVX1_LOC_135/A 0.45fF
C37581 NOR2X1_LOC_208/Y INVX1_LOC_285/Y 0.10fF
C37582 INVX1_LOC_248/A INVX1_LOC_135/A 0.10fF
C37583 NOR2X1_LOC_68/A NOR2X1_LOC_557/A 3.76fF
C37584 INVX1_LOC_234/A INVX1_LOC_172/Y 0.02fF
C37585 NOR2X1_LOC_540/a_36_216# NOR2X1_LOC_553/B 0.02fF
C37586 INVX1_LOC_48/Y NOR2X1_LOC_99/a_36_216# 0.01fF
C37587 INVX1_LOC_103/A NAND2X1_LOC_472/Y 0.13fF
C37588 INVX1_LOC_35/A NOR2X1_LOC_841/A 0.78fF
C37589 NOR2X1_LOC_546/A INVX1_LOC_91/A 0.04fF
C37590 INVX1_LOC_141/A INVX1_LOC_76/A 0.02fF
C37591 NOR2X1_LOC_328/Y NOR2X1_LOC_53/a_36_216# 0.00fF
C37592 NAND2X1_LOC_860/A NAND2X1_LOC_477/Y 0.03fF
C37593 NOR2X1_LOC_658/Y NAND2X1_LOC_469/B 0.14fF
C37594 NOR2X1_LOC_526/Y NAND2X1_LOC_866/B 0.05fF
C37595 INVX1_LOC_39/A INVX1_LOC_89/Y 0.01fF
C37596 NAND2X1_LOC_463/B GATE_811 0.03fF
C37597 NOR2X1_LOC_369/Y NAND2X1_LOC_721/A 0.04fF
C37598 INVX1_LOC_49/A INVX1_LOC_286/A 0.01fF
C37599 INVX1_LOC_45/A INVX1_LOC_20/A 0.10fF
C37600 NAND2X1_LOC_656/Y NOR2X1_LOC_188/a_36_216# 0.02fF
C37601 NAND2X1_LOC_703/Y INVX1_LOC_185/A 0.00fF
C37602 INVX1_LOC_290/A NOR2X1_LOC_747/a_36_216# 0.00fF
C37603 NOR2X1_LOC_757/A INVX1_LOC_279/A 0.01fF
C37604 INVX1_LOC_32/A NOR2X1_LOC_465/Y 1.18fF
C37605 NOR2X1_LOC_688/Y VDD 0.18fF
C37606 INVX1_LOC_135/A NOR2X1_LOC_521/Y 0.02fF
C37607 INPUT_0 NOR2X1_LOC_278/A 0.04fF
C37608 NOR2X1_LOC_191/B INVX1_LOC_93/Y 0.36fF
C37609 INVX1_LOC_58/A INVX1_LOC_29/A 0.07fF
C37610 NAND2X1_LOC_854/a_36_24# INVX1_LOC_76/A 0.01fF
C37611 D_INPUT_0 NAND2X1_LOC_358/Y 2.73fF
C37612 NOR2X1_LOC_348/Y INVX1_LOC_92/A 0.15fF
C37613 NAND2X1_LOC_374/Y NAND2X1_LOC_849/A 0.02fF
C37614 INVX1_LOC_196/Y NOR2X1_LOC_687/Y 3.79fF
C37615 INVX1_LOC_24/A INVX1_LOC_59/Y 0.00fF
C37616 NAND2X1_LOC_778/Y INVX1_LOC_285/A 0.26fF
C37617 INVX1_LOC_172/Y NOR2X1_LOC_19/B 0.06fF
C37618 NOR2X1_LOC_16/Y NOR2X1_LOC_188/A 0.02fF
C37619 NOR2X1_LOC_13/Y NAND2X1_LOC_655/B 0.01fF
C37620 NOR2X1_LOC_255/a_36_216# INPUT_1 0.00fF
C37621 INVX1_LOC_103/A NAND2X1_LOC_434/Y 0.03fF
C37622 NOR2X1_LOC_48/B NOR2X1_LOC_451/a_36_216# 0.00fF
C37623 INVX1_LOC_203/A NOR2X1_LOC_291/Y 0.14fF
C37624 NOR2X1_LOC_629/A INVX1_LOC_284/A 0.07fF
C37625 NOR2X1_LOC_441/Y NAND2X1_LOC_848/A 0.03fF
C37626 D_INPUT_0 NOR2X1_LOC_99/B 0.07fF
C37627 NOR2X1_LOC_716/B NOR2X1_LOC_405/A 0.03fF
C37628 NOR2X1_LOC_804/B INVX1_LOC_65/A 0.10fF
C37629 INVX1_LOC_24/A INVX1_LOC_176/A 0.01fF
C37630 NOR2X1_LOC_510/Y INVX1_LOC_63/A 0.07fF
C37631 NAND2X1_LOC_57/a_36_24# INVX1_LOC_117/A 0.00fF
C37632 INVX1_LOC_71/A INVX1_LOC_20/A 0.08fF
C37633 NAND2X1_LOC_112/Y NOR2X1_LOC_135/Y 0.02fF
C37634 NOR2X1_LOC_521/Y NOR2X1_LOC_490/Y 0.00fF
C37635 NOR2X1_LOC_791/B INVX1_LOC_12/Y 0.03fF
C37636 NOR2X1_LOC_210/B INVX1_LOC_75/A 0.16fF
C37637 INVX1_LOC_2/A INVX1_LOC_286/A 0.10fF
C37638 INVX1_LOC_11/A INVX1_LOC_307/A 0.07fF
C37639 NOR2X1_LOC_373/Y INPUT_1 0.02fF
C37640 INVX1_LOC_256/A INVX1_LOC_92/A 0.13fF
C37641 NAND2X1_LOC_508/A NOR2X1_LOC_199/B 0.10fF
C37642 INVX1_LOC_85/A NOR2X1_LOC_562/B 0.02fF
C37643 NOR2X1_LOC_589/A INVX1_LOC_102/Y 0.08fF
C37644 NAND2X1_LOC_624/B INVX1_LOC_284/A 0.07fF
C37645 NOR2X1_LOC_457/A NOR2X1_LOC_155/A 0.00fF
C37646 INVX1_LOC_28/Y INVX1_LOC_4/Y 0.04fF
C37647 NOR2X1_LOC_15/Y INVX1_LOC_285/A 0.04fF
C37648 INVX1_LOC_224/Y INVX1_LOC_4/A 0.03fF
C37649 INVX1_LOC_11/A NOR2X1_LOC_445/B 0.07fF
C37650 INVX1_LOC_23/A D_INPUT_5 0.01fF
C37651 INVX1_LOC_88/A NOR2X1_LOC_127/a_36_216# 0.00fF
C37652 NOR2X1_LOC_15/Y INVX1_LOC_265/Y 0.01fF
C37653 NOR2X1_LOC_226/A INVX1_LOC_286/A 0.29fF
C37654 NOR2X1_LOC_757/A INVX1_LOC_182/Y 0.01fF
C37655 NOR2X1_LOC_721/Y INVX1_LOC_1/Y 0.03fF
C37656 NOR2X1_LOC_15/Y NOR2X1_LOC_814/A 0.03fF
C37657 INVX1_LOC_311/A NAND2X1_LOC_479/Y 0.03fF
C37658 NOR2X1_LOC_548/Y NOR2X1_LOC_337/A 0.18fF
C37659 INVX1_LOC_50/Y NOR2X1_LOC_67/Y -0.00fF
C37660 NOR2X1_LOC_361/B INVX1_LOC_63/A 0.11fF
C37661 NOR2X1_LOC_840/A NOR2X1_LOC_833/B 0.01fF
C37662 INVX1_LOC_271/A NAND2X1_LOC_454/Y 0.01fF
C37663 NOR2X1_LOC_561/Y NOR2X1_LOC_313/Y 0.04fF
C37664 INVX1_LOC_90/A NOR2X1_LOC_329/B 0.35fF
C37665 INVX1_LOC_30/A NOR2X1_LOC_155/A 0.50fF
C37666 NOR2X1_LOC_226/A INVX1_LOC_95/A 0.02fF
C37667 INVX1_LOC_53/A NAND2X1_LOC_470/B 0.04fF
C37668 NAND2X1_LOC_354/B NAND2X1_LOC_687/a_36_24# 0.00fF
C37669 INVX1_LOC_33/A NAND2X1_LOC_96/A 0.09fF
C37670 INVX1_LOC_58/A INVX1_LOC_298/Y 0.07fF
C37671 INVX1_LOC_295/A NAND2X1_LOC_51/B 0.06fF
C37672 NOR2X1_LOC_310/Y INVX1_LOC_46/A 0.01fF
C37673 INVX1_LOC_61/A NAND2X1_LOC_243/Y 0.03fF
C37674 INVX1_LOC_75/A INVX1_LOC_20/Y 0.02fF
C37675 NAND2X1_LOC_564/B NOR2X1_LOC_45/B 0.08fF
C37676 INVX1_LOC_296/A NOR2X1_LOC_635/B 0.48fF
C37677 INVX1_LOC_8/A INVX1_LOC_117/A 0.07fF
C37678 INVX1_LOC_239/A INVX1_LOC_42/A 0.09fF
C37679 INVX1_LOC_159/A INVX1_LOC_117/Y 0.85fF
C37680 INVX1_LOC_221/Y INVX1_LOC_264/A 0.06fF
C37681 INVX1_LOC_136/A NAND2X1_LOC_240/a_36_24# 0.00fF
C37682 NAND2X1_LOC_159/a_36_24# INVX1_LOC_91/A 0.02fF
C37683 INVX1_LOC_18/A INVX1_LOC_107/Y 0.04fF
C37684 INVX1_LOC_77/A NOR2X1_LOC_641/Y 0.00fF
C37685 INVX1_LOC_95/Y INVX1_LOC_53/Y 0.33fF
C37686 INVX1_LOC_17/Y INVX1_LOC_57/A 0.01fF
C37687 NOR2X1_LOC_851/a_36_216# NOR2X1_LOC_858/A 0.02fF
C37688 INVX1_LOC_49/A INVX1_LOC_54/A 0.03fF
C37689 INVX1_LOC_11/A INVX1_LOC_12/A 0.39fF
C37690 INVX1_LOC_200/A NOR2X1_LOC_89/A 0.47fF
C37691 INVX1_LOC_204/Y INVX1_LOC_78/A 0.25fF
C37692 INVX1_LOC_303/A NAND2X1_LOC_488/a_36_24# 0.00fF
C37693 NOR2X1_LOC_686/B NAND2X1_LOC_655/A 0.08fF
C37694 INVX1_LOC_62/Y NAND2X1_LOC_85/Y 0.40fF
C37695 INVX1_LOC_286/A INPUT_1 0.03fF
C37696 NAND2X1_LOC_326/A INVX1_LOC_15/A 0.07fF
C37697 NOR2X1_LOC_151/Y NOR2X1_LOC_180/a_36_216# 0.00fF
C37698 INVX1_LOC_25/A D_INPUT_1 0.30fF
C37699 INVX1_LOC_129/A NAND2X1_LOC_275/a_36_24# 0.02fF
C37700 INVX1_LOC_27/A NAND2X1_LOC_454/Y 0.07fF
C37701 NOR2X1_LOC_593/Y INVX1_LOC_307/A 0.07fF
C37702 NOR2X1_LOC_667/A NOR2X1_LOC_152/A 0.08fF
C37703 INVX1_LOC_1/Y VDD 0.65fF
C37704 INVX1_LOC_64/A INVX1_LOC_224/Y 0.01fF
C37705 INVX1_LOC_255/Y D_INPUT_3 0.17fF
C37706 INVX1_LOC_41/Y INVX1_LOC_119/Y 0.06fF
C37707 INVX1_LOC_2/A NOR2X1_LOC_602/B 0.02fF
C37708 NOR2X1_LOC_78/B NOR2X1_LOC_536/A 0.10fF
C37709 INVX1_LOC_36/A NAND2X1_LOC_81/B 0.03fF
C37710 NAND2X1_LOC_218/B NOR2X1_LOC_673/A 0.06fF
C37711 INVX1_LOC_5/A NOR2X1_LOC_840/Y 0.00fF
C37712 NOR2X1_LOC_769/A NOR2X1_LOC_48/Y 0.00fF
C37713 INVX1_LOC_40/A NAND2X1_LOC_96/A 0.04fF
C37714 INVX1_LOC_39/A INVX1_LOC_16/Y 0.10fF
C37715 NOR2X1_LOC_593/Y NOR2X1_LOC_445/B 0.37fF
C37716 NOR2X1_LOC_130/A INVX1_LOC_59/Y 0.10fF
C37717 NOR2X1_LOC_598/B NAND2X1_LOC_363/B 0.10fF
C37718 INVX1_LOC_135/A NOR2X1_LOC_670/Y 0.10fF
C37719 INVX1_LOC_90/A INPUT_4 0.03fF
C37720 NOR2X1_LOC_222/Y INVX1_LOC_38/A 0.20fF
C37721 NOR2X1_LOC_510/Y NOR2X1_LOC_65/Y 0.00fF
C37722 NOR2X1_LOC_860/B NOR2X1_LOC_814/A 0.07fF
C37723 NOR2X1_LOC_564/Y INVX1_LOC_91/A 0.62fF
C37724 NOR2X1_LOC_103/Y INVX1_LOC_4/A 0.07fF
C37725 INVX1_LOC_40/A NAND2X1_LOC_93/a_36_24# 0.00fF
C37726 NOR2X1_LOC_267/A NAND2X1_LOC_81/B 0.04fF
C37727 INVX1_LOC_2/A INVX1_LOC_54/A 0.41fF
C37728 INVX1_LOC_95/A INPUT_1 0.00fF
C37729 INVX1_LOC_18/A INVX1_LOC_272/A 0.08fF
C37730 NOR2X1_LOC_92/Y NOR2X1_LOC_278/Y 4.05fF
C37731 NAND2X1_LOC_30/Y NAND2X1_LOC_3/B 1.50fF
C37732 INVX1_LOC_279/A INVX1_LOC_37/A 0.14fF
C37733 INVX1_LOC_51/A NAND2X1_LOC_363/B 0.03fF
C37734 INVX1_LOC_30/A NOR2X1_LOC_833/B 0.03fF
C37735 NOR2X1_LOC_123/B INVX1_LOC_20/A 0.23fF
C37736 NAND2X1_LOC_787/A NAND2X1_LOC_725/A 0.01fF
C37737 NOR2X1_LOC_598/B NOR2X1_LOC_640/a_36_216# 0.01fF
C37738 INVX1_LOC_57/A NOR2X1_LOC_406/A 0.03fF
C37739 NOR2X1_LOC_226/A INVX1_LOC_54/A 0.44fF
C37740 NAND2X1_LOC_705/Y NOR2X1_LOC_693/Y 0.00fF
C37741 INVX1_LOC_34/Y NOR2X1_LOC_99/Y 0.31fF
C37742 INVX1_LOC_25/A NOR2X1_LOC_652/Y 0.17fF
C37743 INVX1_LOC_217/A NOR2X1_LOC_89/A 0.09fF
C37744 INVX1_LOC_39/A NAND2X1_LOC_205/A 0.03fF
C37745 INVX1_LOC_2/Y NOR2X1_LOC_814/Y 0.16fF
C37746 INVX1_LOC_255/Y INVX1_LOC_230/A 0.00fF
C37747 NOR2X1_LOC_709/A NOR2X1_LOC_831/B 0.02fF
C37748 NOR2X1_LOC_78/B NAND2X1_LOC_93/B 0.03fF
C37749 INVX1_LOC_299/A NOR2X1_LOC_798/Y 0.01fF
C37750 INVX1_LOC_193/Y INVX1_LOC_86/Y 0.02fF
C37751 NAND2X1_LOC_392/Y NOR2X1_LOC_536/A 0.03fF
C37752 NOR2X1_LOC_589/A NOR2X1_LOC_331/B 0.07fF
C37753 NOR2X1_LOC_655/B INVX1_LOC_46/Y 0.10fF
C37754 NOR2X1_LOC_521/Y INVX1_LOC_280/A 0.01fF
C37755 NAND2X1_LOC_567/Y INVX1_LOC_49/Y 0.15fF
C37756 NOR2X1_LOC_550/B INVX1_LOC_19/A 0.01fF
C37757 NOR2X1_LOC_91/Y INVX1_LOC_42/A 0.03fF
C37758 NOR2X1_LOC_99/B NOR2X1_LOC_859/Y 0.02fF
C37759 INVX1_LOC_89/A NOR2X1_LOC_706/B 0.00fF
C37760 INVX1_LOC_80/Y NOR2X1_LOC_649/B 0.01fF
C37761 NAND2X1_LOC_3/a_36_24# INVX1_LOC_15/A 0.00fF
C37762 INVX1_LOC_174/A NAND2X1_LOC_467/a_36_24# 0.00fF
C37763 INVX1_LOC_22/A NOR2X1_LOC_612/Y 0.01fF
C37764 INVX1_LOC_230/Y NOR2X1_LOC_825/a_36_216# 0.00fF
C37765 INVX1_LOC_45/A INVX1_LOC_4/A 0.03fF
C37766 NOR2X1_LOC_590/A INVX1_LOC_273/A 0.03fF
C37767 INVX1_LOC_299/A NOR2X1_LOC_748/A 0.10fF
C37768 NOR2X1_LOC_643/Y NAND2X1_LOC_207/Y 0.02fF
C37769 INVX1_LOC_83/A NOR2X1_LOC_536/A 0.01fF
C37770 NOR2X1_LOC_568/A INVX1_LOC_4/A 0.14fF
C37771 NOR2X1_LOC_459/A NAND2X1_LOC_659/a_36_24# 0.00fF
C37772 NOR2X1_LOC_205/Y INVX1_LOC_270/A 0.03fF
C37773 NOR2X1_LOC_433/A INVX1_LOC_12/A 0.09fF
C37774 NOR2X1_LOC_85/a_36_216# NAND2X1_LOC_243/Y 0.01fF
C37775 D_INPUT_1 INVX1_LOC_1/A 0.13fF
C37776 INVX1_LOC_269/A INVX1_LOC_29/Y 0.10fF
C37777 INVX1_LOC_36/A INVX1_LOC_4/Y 0.01fF
C37778 NOR2X1_LOC_674/a_36_216# NOR2X1_LOC_674/Y 0.00fF
C37779 NOR2X1_LOC_538/B NOR2X1_LOC_748/A 0.02fF
C37780 NAND2X1_LOC_504/a_36_24# INVX1_LOC_122/A 0.00fF
C37781 INVX1_LOC_279/A INVX1_LOC_157/Y 0.02fF
C37782 INVX1_LOC_50/A NOR2X1_LOC_217/a_36_216# 0.01fF
C37783 INVX1_LOC_177/A INVX1_LOC_63/A 0.03fF
C37784 NAND2X1_LOC_360/B INVX1_LOC_84/A 1.16fF
C37785 NOR2X1_LOC_742/A VDD 1.18fF
C37786 NOR2X1_LOC_843/A NOR2X1_LOC_633/A 0.01fF
C37787 NOR2X1_LOC_373/Y INVX1_LOC_118/A 0.10fF
C37788 NOR2X1_LOC_256/a_36_216# INVX1_LOC_3/Y 0.01fF
C37789 NOR2X1_LOC_112/B INVX1_LOC_176/A 0.18fF
C37790 NOR2X1_LOC_78/B INVX1_LOC_3/A 0.00fF
C37791 NOR2X1_LOC_368/A INVX1_LOC_76/A 0.03fF
C37792 NAND2X1_LOC_833/Y INVX1_LOC_102/A 0.02fF
C37793 NOR2X1_LOC_309/Y NAND2X1_LOC_81/B 0.08fF
C37794 NOR2X1_LOC_344/a_36_216# INVX1_LOC_29/A 0.00fF
C37795 INVX1_LOC_83/A NOR2X1_LOC_655/Y 0.03fF
C37796 NAND2X1_LOC_319/A NOR2X1_LOC_510/B 0.05fF
C37797 INVX1_LOC_224/Y INVX1_LOC_43/Y -0.01fF
C37798 NOR2X1_LOC_773/Y NOR2X1_LOC_661/a_36_216# 0.00fF
C37799 INVX1_LOC_71/A INVX1_LOC_4/A 0.36fF
C37800 NOR2X1_LOC_91/Y INVX1_LOC_78/A 0.03fF
C37801 NOR2X1_LOC_52/B INVX1_LOC_12/A 1.41fF
C37802 INVX1_LOC_83/A NAND2X1_LOC_93/B 2.16fF
C37803 INVX1_LOC_256/A INVX1_LOC_53/A 0.22fF
C37804 NAND2X1_LOC_858/B INVX1_LOC_37/A 0.07fF
C37805 NOR2X1_LOC_561/Y NOR2X1_LOC_832/a_36_216# 0.01fF
C37806 NOR2X1_LOC_329/B INVX1_LOC_38/A 3.90fF
C37807 NOR2X1_LOC_6/B NOR2X1_LOC_67/Y 0.00fF
C37808 INPUT_1 INVX1_LOC_54/A 0.07fF
C37809 INVX1_LOC_304/Y NOR2X1_LOC_89/A 0.07fF
C37810 INVX1_LOC_311/A INVX1_LOC_139/Y 0.01fF
C37811 NOR2X1_LOC_852/Y NOR2X1_LOC_857/a_36_216# 0.00fF
C37812 NOR2X1_LOC_99/B INVX1_LOC_46/Y 3.12fF
C37813 INVX1_LOC_64/A NOR2X1_LOC_103/Y 0.02fF
C37814 D_INPUT_4 INVX1_LOC_38/A 0.03fF
C37815 INVX1_LOC_49/A NAND2X1_LOC_3/B 0.30fF
C37816 INVX1_LOC_83/A NAND2X1_LOC_425/Y 0.14fF
C37817 INVX1_LOC_1/A NOR2X1_LOC_652/Y 0.30fF
C37818 INVX1_LOC_35/A NOR2X1_LOC_705/B 0.00fF
C37819 INVX1_LOC_8/A INVX1_LOC_3/Y 1.24fF
C37820 NAND2X1_LOC_733/Y NAND2X1_LOC_804/A 0.03fF
C37821 NOR2X1_LOC_791/Y NOR2X1_LOC_271/a_36_216# 0.00fF
C37822 NOR2X1_LOC_603/a_36_216# INVX1_LOC_12/A 0.00fF
C37823 INVX1_LOC_6/Y NAND2X1_LOC_454/Y 0.01fF
C37824 NOR2X1_LOC_769/B INVX1_LOC_30/A 0.06fF
C37825 INVX1_LOC_227/Y NOR2X1_LOC_383/B 0.01fF
C37826 INVX1_LOC_58/A NAND2X1_LOC_721/B 0.48fF
C37827 NOR2X1_LOC_318/B VDD 1.02fF
C37828 INVX1_LOC_2/A NOR2X1_LOC_48/B 1.92fF
C37829 INVX1_LOC_83/A NOR2X1_LOC_649/B 0.52fF
C37830 NAND2X1_LOC_763/B NOR2X1_LOC_769/B 0.15fF
C37831 NAND2X1_LOC_573/A INVX1_LOC_63/A 0.01fF
C37832 NOR2X1_LOC_274/Y INVX1_LOC_26/A -0.00fF
C37833 INVX1_LOC_83/A INVX1_LOC_3/A 0.07fF
C37834 INVX1_LOC_5/A NAND2X1_LOC_114/B 0.07fF
C37835 NOR2X1_LOC_598/B INVX1_LOC_30/A 2.67fF
C37836 INVX1_LOC_88/A NOR2X1_LOC_173/Y 0.11fF
C37837 NOR2X1_LOC_68/A INVX1_LOC_271/A 0.03fF
C37838 NOR2X1_LOC_87/B INVX1_LOC_15/A 0.08fF
C37839 D_INPUT_4 NOR2X1_LOC_51/A 0.01fF
C37840 NOR2X1_LOC_226/A NOR2X1_LOC_48/B 4.79fF
C37841 NAND2X1_LOC_763/B NOR2X1_LOC_598/B 0.19fF
C37842 INVX1_LOC_93/Y VDD 1.66fF
C37843 NOR2X1_LOC_309/Y INVX1_LOC_4/Y 0.08fF
C37844 NOR2X1_LOC_360/Y INVX1_LOC_23/A 0.10fF
C37845 NAND2X1_LOC_354/B INVX1_LOC_273/A 0.06fF
C37846 INVX1_LOC_217/A NAND2X1_LOC_804/A 0.02fF
C37847 INVX1_LOC_45/A INVX1_LOC_64/A 7.12fF
C37848 INVX1_LOC_41/A NOR2X1_LOC_278/Y 0.03fF
C37849 INVX1_LOC_226/Y NAND2X1_LOC_254/Y 0.10fF
C37850 INVX1_LOC_233/Y INVX1_LOC_36/A 0.09fF
C37851 NAND2X1_LOC_714/B INVX1_LOC_161/Y 0.03fF
C37852 NAND2X1_LOC_490/a_36_24# NAND2X1_LOC_96/A 0.00fF
C37853 INVX1_LOC_64/A NAND2X1_LOC_856/A 0.03fF
C37854 INVX1_LOC_108/Y NAND2X1_LOC_481/a_36_24# 0.00fF
C37855 NOR2X1_LOC_570/B NOR2X1_LOC_631/Y 0.00fF
C37856 INVX1_LOC_119/A INVX1_LOC_94/Y 0.01fF
C37857 INVX1_LOC_33/A NAND2X1_LOC_99/A 0.07fF
C37858 INVX1_LOC_286/A INVX1_LOC_118/A 0.03fF
C37859 NOR2X1_LOC_91/A INVX1_LOC_207/A 0.13fF
C37860 NOR2X1_LOC_6/B NOR2X1_LOC_415/Y 0.07fF
C37861 NOR2X1_LOC_332/A NAND2X1_LOC_82/Y 0.01fF
C37862 NOR2X1_LOC_311/Y NOR2X1_LOC_536/A 0.01fF
C37863 INVX1_LOC_1/A NOR2X1_LOC_241/A 0.02fF
C37864 NOR2X1_LOC_294/Y INVX1_LOC_5/A 0.68fF
C37865 INVX1_LOC_235/A NAND2X1_LOC_555/Y 0.04fF
C37866 INVX1_LOC_187/Y INVX1_LOC_77/Y 0.02fF
C37867 NOR2X1_LOC_513/Y NAND2X1_LOC_537/Y 0.00fF
C37868 NOR2X1_LOC_667/Y NAND2X1_LOC_703/Y 0.01fF
C37869 INVX1_LOC_178/A INVX1_LOC_141/Y 0.01fF
C37870 VDD INVX1_LOC_139/A 0.01fF
C37871 INVX1_LOC_50/A INVX1_LOC_155/A 0.00fF
C37872 NOR2X1_LOC_372/Y NOR2X1_LOC_291/Y 0.14fF
C37873 NAND2X1_LOC_361/Y INVX1_LOC_57/A 0.10fF
C37874 INVX1_LOC_69/Y INVX1_LOC_92/A 0.07fF
C37875 NOR2X1_LOC_52/B NOR2X1_LOC_686/A 0.03fF
C37876 NAND2X1_LOC_555/Y NAND2X1_LOC_393/a_36_24# 0.01fF
C37877 INVX1_LOC_136/A NOR2X1_LOC_220/B 0.03fF
C37878 NAND2X1_LOC_808/A NOR2X1_LOC_89/A 0.07fF
C37879 NAND2X1_LOC_214/B NOR2X1_LOC_68/A 1.17fF
C37880 INVX1_LOC_276/Y INVX1_LOC_273/A 0.02fF
C37881 NOR2X1_LOC_536/A NOR2X1_LOC_368/Y 0.01fF
C37882 INVX1_LOC_266/Y NOR2X1_LOC_45/a_36_216# 0.00fF
C37883 NOR2X1_LOC_15/Y NOR2X1_LOC_590/A 0.03fF
C37884 INVX1_LOC_50/A NOR2X1_LOC_264/Y 0.07fF
C37885 NAND2X1_LOC_787/B NAND2X1_LOC_804/A 0.00fF
C37886 INVX1_LOC_64/A INVX1_LOC_71/A 0.14fF
C37887 NAND2X1_LOC_721/A VDD 0.32fF
C37888 INVX1_LOC_34/A NOR2X1_LOC_414/Y 0.12fF
C37889 INVX1_LOC_62/A NAND2X1_LOC_206/B 0.52fF
C37890 INVX1_LOC_51/Y NAND2X1_LOC_85/Y 0.00fF
C37891 NOR2X1_LOC_658/Y INVX1_LOC_52/Y 0.01fF
C37892 INVX1_LOC_147/Y NOR2X1_LOC_331/B 0.05fF
C37893 INVX1_LOC_58/A INVX1_LOC_8/A 0.15fF
C37894 INVX1_LOC_289/Y INVX1_LOC_286/Y 0.00fF
C37895 NOR2X1_LOC_670/Y INVX1_LOC_280/A 0.01fF
C37896 INVX1_LOC_43/Y NOR2X1_LOC_103/Y 0.24fF
C37897 INVX1_LOC_72/A NOR2X1_LOC_440/B 0.32fF
C37898 INVX1_LOC_27/A NOR2X1_LOC_68/A 0.19fF
C37899 NOR2X1_LOC_612/B NOR2X1_LOC_383/B 0.46fF
C37900 NOR2X1_LOC_226/A NOR2X1_LOC_438/Y 0.03fF
C37901 NOR2X1_LOC_51/A INPUT_4 0.01fF
C37902 NOR2X1_LOC_536/A INVX1_LOC_46/A 9.04fF
C37903 NOR2X1_LOC_363/Y INVX1_LOC_12/Y 0.07fF
C37904 INVX1_LOC_111/Y NOR2X1_LOC_383/B 0.00fF
C37905 NAND2X1_LOC_338/B NOR2X1_LOC_720/A 0.04fF
C37906 NAND2X1_LOC_642/a_36_24# NAND2X1_LOC_96/A 0.00fF
C37907 NAND2X1_LOC_648/A NOR2X1_LOC_48/B 0.00fF
C37908 INVX1_LOC_57/Y INVX1_LOC_14/A 0.11fF
C37909 INVX1_LOC_204/Y INVX1_LOC_113/Y 0.01fF
C37910 INPUT_1 NOR2X1_LOC_48/B 0.05fF
C37911 INVX1_LOC_36/A NOR2X1_LOC_205/Y 0.03fF
C37912 INVX1_LOC_2/A NAND2X1_LOC_215/A 0.12fF
C37913 NOR2X1_LOC_665/A INVX1_LOC_271/Y 0.07fF
C37914 INVX1_LOC_40/A NAND2X1_LOC_99/A 0.07fF
C37915 INVX1_LOC_35/A NOR2X1_LOC_392/B 0.03fF
C37916 D_INPUT_0 NOR2X1_LOC_28/a_36_216# 0.00fF
C37917 INVX1_LOC_34/A NOR2X1_LOC_665/Y 0.01fF
C37918 NOR2X1_LOC_778/A INVX1_LOC_1/A 0.24fF
C37919 INVX1_LOC_165/Y NAND2X1_LOC_99/A 0.02fF
C37920 INVX1_LOC_5/A NOR2X1_LOC_219/B 0.04fF
C37921 NOR2X1_LOC_442/a_36_216# NAND2X1_LOC_364/A 0.00fF
C37922 NOR2X1_LOC_816/A INVX1_LOC_141/Y 0.03fF
C37923 INVX1_LOC_108/Y NOR2X1_LOC_87/B 0.03fF
C37924 NOR2X1_LOC_123/B INVX1_LOC_4/A -0.01fF
C37925 NOR2X1_LOC_586/Y INVX1_LOC_54/A 0.11fF
C37926 NAND2X1_LOC_337/B INVX1_LOC_312/Y 0.00fF
C37927 VDD NOR2X1_LOC_856/A 0.23fF
C37928 INVX1_LOC_83/A NAND2X1_LOC_470/B 0.00fF
C37929 NOR2X1_LOC_78/A NAND2X1_LOC_42/a_36_24# 0.00fF
C37930 NOR2X1_LOC_334/A INVX1_LOC_19/A 0.02fF
C37931 INVX1_LOC_1/A D_INPUT_2 0.07fF
C37932 INVX1_LOC_136/A INVX1_LOC_225/Y 0.10fF
C37933 INVX1_LOC_202/A NOR2X1_LOC_122/A 0.04fF
C37934 NAND2X1_LOC_796/B NAND2X1_LOC_325/Y 0.10fF
C37935 INVX1_LOC_150/Y INVX1_LOC_18/A 0.02fF
C37936 NAND2X1_LOC_93/B INVX1_LOC_46/A 0.16fF
C37937 NAND2X1_LOC_725/A NAND2X1_LOC_722/A 0.10fF
C37938 INVX1_LOC_44/A INVX1_LOC_9/A 0.07fF
C37939 INVX1_LOC_103/A INVX1_LOC_24/A 0.04fF
C37940 NOR2X1_LOC_589/A NOR2X1_LOC_106/a_36_216# 0.01fF
C37941 INVX1_LOC_286/A NAND2X1_LOC_63/Y 0.03fF
C37942 VDD INVX1_LOC_117/Y 0.21fF
C37943 NOR2X1_LOC_208/Y NOR2X1_LOC_205/Y 0.14fF
C37944 INVX1_LOC_104/A INVX1_LOC_50/Y 0.07fF
C37945 INVX1_LOC_196/Y INVX1_LOC_274/Y 0.19fF
C37946 INVX1_LOC_37/A NOR2X1_LOC_624/B 0.02fF
C37947 NOR2X1_LOC_791/B NOR2X1_LOC_160/B 0.03fF
C37948 INVX1_LOC_5/A NOR2X1_LOC_168/B 0.03fF
C37949 NOR2X1_LOC_318/B INVX1_LOC_133/A 0.03fF
C37950 VDD NAND2X1_LOC_770/Y 0.01fF
C37951 INVX1_LOC_292/A INVX1_LOC_24/A 0.07fF
C37952 NAND2X1_LOC_374/Y NOR2X1_LOC_291/Y 0.12fF
C37953 NOR2X1_LOC_789/B NOR2X1_LOC_709/A 0.06fF
C37954 NOR2X1_LOC_447/B NOR2X1_LOC_697/Y 0.02fF
C37955 NOR2X1_LOC_137/A NOR2X1_LOC_383/B 0.10fF
C37956 INVX1_LOC_54/A INVX1_LOC_118/A 0.38fF
C37957 NOR2X1_LOC_510/Y NOR2X1_LOC_362/a_36_216# 0.02fF
C37958 NOR2X1_LOC_459/A NOR2X1_LOC_476/B 0.37fF
C37959 NOR2X1_LOC_254/A INVX1_LOC_77/A 0.18fF
C37960 INVX1_LOC_266/A INVX1_LOC_104/A 0.39fF
C37961 NAND2X1_LOC_350/A INVX1_LOC_49/A 0.07fF
C37962 INVX1_LOC_89/A INVX1_LOC_296/A 0.72fF
C37963 INVX1_LOC_284/Y NAND2X1_LOC_837/Y 0.15fF
C37964 INVX1_LOC_89/A NOR2X1_LOC_621/a_36_216# 0.00fF
C37965 INVX1_LOC_157/A INVX1_LOC_53/A 0.49fF
C37966 NAND2X1_LOC_391/a_36_24# NOR2X1_LOC_384/Y 0.01fF
C37967 NAND2X1_LOC_860/a_36_24# INVX1_LOC_71/A 0.00fF
C37968 INVX1_LOC_199/A INVX1_LOC_12/A 0.07fF
C37969 NOR2X1_LOC_209/a_36_216# INVX1_LOC_213/A 0.01fF
C37970 INVX1_LOC_218/Y INVX1_LOC_49/A 0.03fF
C37971 INVX1_LOC_142/A INVX1_LOC_198/Y 0.44fF
C37972 NAND2X1_LOC_778/Y NOR2X1_LOC_488/Y 0.01fF
C37973 INVX1_LOC_41/A NOR2X1_LOC_197/A 0.01fF
C37974 NOR2X1_LOC_82/A NOR2X1_LOC_4/a_36_216# 0.00fF
C37975 INPUT_1 NAND2X1_LOC_215/A 0.09fF
C37976 NAND2X1_LOC_149/Y NOR2X1_LOC_769/a_36_216# 0.00fF
C37977 INVX1_LOC_243/Y NAND2X1_LOC_654/B 0.12fF
C37978 INVX1_LOC_279/Y NOR2X1_LOC_374/A 0.01fF
C37979 NOR2X1_LOC_441/Y INVX1_LOC_49/A 0.03fF
C37980 NOR2X1_LOC_721/Y INVX1_LOC_87/A 0.19fF
C37981 INVX1_LOC_12/A INVX1_LOC_74/A 0.24fF
C37982 NOR2X1_LOC_764/Y INVX1_LOC_53/A 0.03fF
C37983 INVX1_LOC_200/A NOR2X1_LOC_52/B 0.17fF
C37984 NOR2X1_LOC_805/a_36_216# INVX1_LOC_177/A 0.00fF
C37985 NOR2X1_LOC_360/Y INVX1_LOC_111/A 0.00fF
C37986 NOR2X1_LOC_67/A NOR2X1_LOC_232/a_36_216# 0.01fF
C37987 NOR2X1_LOC_361/B NOR2X1_LOC_362/a_36_216# 0.00fF
C37988 INVX1_LOC_100/A NAND2X1_LOC_400/a_36_24# 0.01fF
C37989 INVX1_LOC_14/A NAND2X1_LOC_347/a_36_24# 0.01fF
C37990 NOR2X1_LOC_400/A INVX1_LOC_135/A 0.03fF
C37991 INVX1_LOC_268/A NAND2X1_LOC_149/Y 0.09fF
C37992 INVX1_LOC_39/A NOR2X1_LOC_255/a_36_216# 0.00fF
C37993 INVX1_LOC_35/A INVX1_LOC_90/A 1.88fF
C37994 NOR2X1_LOC_160/B NOR2X1_LOC_802/A 0.07fF
C37995 NOR2X1_LOC_658/Y INVX1_LOC_63/Y 1.18fF
C37996 VDD NOR2X1_LOC_669/A 0.00fF
C37997 NOR2X1_LOC_567/B INVX1_LOC_23/A 0.07fF
C37998 NAND2X1_LOC_583/a_36_24# NAND2X1_LOC_11/Y 0.00fF
C37999 NAND2X1_LOC_204/a_36_24# NOR2X1_LOC_814/A 0.01fF
C38000 INVX1_LOC_28/A NAND2X1_LOC_590/a_36_24# 0.01fF
C38001 INVX1_LOC_256/A NOR2X1_LOC_78/B 3.84fF
C38002 INVX1_LOC_147/A INVX1_LOC_271/A 0.07fF
C38003 NOR2X1_LOC_334/A INVX1_LOC_26/Y 0.03fF
C38004 NOR2X1_LOC_155/A INVX1_LOC_113/A 0.07fF
C38005 INVX1_LOC_185/A INVX1_LOC_119/Y 0.02fF
C38006 NOR2X1_LOC_158/Y INVX1_LOC_91/A 0.22fF
C38007 NAND2X1_LOC_549/B NOR2X1_LOC_530/Y 0.22fF
C38008 NOR2X1_LOC_226/A NAND2X1_LOC_350/A 0.51fF
C38009 INVX1_LOC_202/A NOR2X1_LOC_437/Y 0.11fF
C38010 INVX1_LOC_136/A NAND2X1_LOC_811/Y 0.02fF
C38011 NOR2X1_LOC_248/Y INVX1_LOC_104/A 0.08fF
C38012 NOR2X1_LOC_216/B NOR2X1_LOC_49/a_36_216# 0.01fF
C38013 NOR2X1_LOC_770/B INVX1_LOC_18/A 0.03fF
C38014 INVX1_LOC_313/Y NOR2X1_LOC_674/a_36_216# 0.00fF
C38015 INVX1_LOC_11/A D_GATE_222 0.00fF
C38016 INVX1_LOC_2/A NOR2X1_LOC_441/Y 0.07fF
C38017 INVX1_LOC_269/A INVX1_LOC_101/A 0.00fF
C38018 INVX1_LOC_17/A NAND2X1_LOC_349/B 0.11fF
C38019 NOR2X1_LOC_609/a_36_216# NOR2X1_LOC_577/Y 0.01fF
C38020 NOR2X1_LOC_664/Y NOR2X1_LOC_68/A 0.02fF
C38021 NOR2X1_LOC_15/Y INVX1_LOC_227/A 0.13fF
C38022 INVX1_LOC_282/A NAND2X1_LOC_793/B 0.04fF
C38023 INVX1_LOC_30/A NAND2X1_LOC_660/A 1.25fF
C38024 NAND2X1_LOC_391/Y NAND2X1_LOC_551/A 0.46fF
C38025 INVX1_LOC_35/A NAND2X1_LOC_348/A 0.07fF
C38026 NOR2X1_LOC_590/A INVX1_LOC_226/A 0.03fF
C38027 INVX1_LOC_217/A NOR2X1_LOC_52/B 0.05fF
C38028 NOR2X1_LOC_590/A NAND2X1_LOC_840/B 0.05fF
C38029 NOR2X1_LOC_13/Y INVX1_LOC_63/Y 0.13fF
C38030 INVX1_LOC_136/A INVX1_LOC_266/Y 0.00fF
C38031 NOR2X1_LOC_92/Y NAND2X1_LOC_809/A 0.03fF
C38032 NOR2X1_LOC_794/B NOR2X1_LOC_553/Y 0.00fF
C38033 INVX1_LOC_235/Y INVX1_LOC_175/Y 0.16fF
C38034 INVX1_LOC_269/A NOR2X1_LOC_355/A 0.33fF
C38035 INVX1_LOC_69/Y INVX1_LOC_53/A 0.01fF
C38036 INVX1_LOC_41/A NAND2X1_LOC_7/Y 0.01fF
C38037 INVX1_LOC_24/A INVX1_LOC_240/A 0.03fF
C38038 NAND2X1_LOC_659/B NAND2X1_LOC_619/a_36_24# 0.01fF
C38039 INVX1_LOC_230/Y NOR2X1_LOC_719/A 0.01fF
C38040 INVX1_LOC_84/A NAND2X1_LOC_572/B 0.07fF
C38041 NAND2X1_LOC_659/B INVX1_LOC_175/A 0.05fF
C38042 INVX1_LOC_135/A NOR2X1_LOC_523/A 0.00fF
C38043 NOR2X1_LOC_788/a_36_216# INVX1_LOC_53/A 0.01fF
C38044 NAND2X1_LOC_807/B INVX1_LOC_118/A 0.09fF
C38045 INVX1_LOC_49/A NOR2X1_LOC_340/Y 0.00fF
C38046 INVX1_LOC_299/A INVX1_LOC_89/A 0.07fF
C38047 INVX1_LOC_49/A NOR2X1_LOC_142/Y 0.17fF
C38048 INVX1_LOC_103/A NOR2X1_LOC_130/A 0.05fF
C38049 NAND2X1_LOC_470/B INVX1_LOC_46/A 3.76fF
C38050 INVX1_LOC_11/A NAND2X1_LOC_808/A 0.06fF
C38051 NOR2X1_LOC_807/B INVX1_LOC_83/A 0.19fF
C38052 NOR2X1_LOC_269/Y INVX1_LOC_23/A 0.11fF
C38053 VDD INVX1_LOC_87/A 0.39fF
C38054 NOR2X1_LOC_538/B INVX1_LOC_89/A 0.09fF
C38055 NOR2X1_LOC_48/B INVX1_LOC_118/A 0.12fF
C38056 INVX1_LOC_230/Y INVX1_LOC_7/A 0.57fF
C38057 NOR2X1_LOC_68/A NAND2X1_LOC_200/B 0.01fF
C38058 NOR2X1_LOC_89/A INVX1_LOC_92/A 0.20fF
C38059 NOR2X1_LOC_331/B INVX1_LOC_4/A 0.07fF
C38060 NAND2X1_LOC_860/Y NOR2X1_LOC_91/Y 0.01fF
C38061 INVX1_LOC_293/A INVX1_LOC_89/A 0.03fF
C38062 INVX1_LOC_5/A INVX1_LOC_78/Y 0.03fF
C38063 INVX1_LOC_71/A NAND2X1_LOC_850/Y 0.10fF
C38064 INVX1_LOC_295/A INVX1_LOC_174/A 0.25fF
C38065 INVX1_LOC_284/Y NOR2X1_LOC_299/Y 0.01fF
C38066 NAND2X1_LOC_733/A NOR2X1_LOC_298/Y 0.04fF
C38067 NOR2X1_LOC_536/A NOR2X1_LOC_282/a_36_216# 0.02fF
C38068 NAND2X1_LOC_656/A INVX1_LOC_40/A 0.34fF
C38069 NOR2X1_LOC_653/Y NAND2X1_LOC_74/B 0.01fF
C38070 INVX1_LOC_76/A NOR2X1_LOC_696/Y 0.50fF
C38071 NAND2X1_LOC_61/Y NOR2X1_LOC_60/Y 0.21fF
C38072 NAND2X1_LOC_475/Y INVX1_LOC_29/A 0.10fF
C38073 NOR2X1_LOC_238/Y INVX1_LOC_16/A 0.05fF
C38074 NOR2X1_LOC_294/Y NOR2X1_LOC_332/A 0.06fF
C38075 INVX1_LOC_2/A NOR2X1_LOC_142/Y 0.45fF
C38076 INVX1_LOC_221/A NOR2X1_LOC_591/Y 0.00fF
C38077 NOR2X1_LOC_36/a_36_216# D_INPUT_5 0.00fF
C38078 INVX1_LOC_304/Y NOR2X1_LOC_52/B 0.30fF
C38079 INVX1_LOC_17/A INVX1_LOC_75/A 0.18fF
C38080 NOR2X1_LOC_68/A INVX1_LOC_234/A 0.03fF
C38081 NOR2X1_LOC_593/Y NOR2X1_LOC_566/Y 0.01fF
C38082 NOR2X1_LOC_68/A NAND2X1_LOC_156/B 0.03fF
C38083 NOR2X1_LOC_67/A NAND2X1_LOC_139/A 0.02fF
C38084 INVX1_LOC_21/A NOR2X1_LOC_45/B 0.13fF
C38085 NOR2X1_LOC_349/A NOR2X1_LOC_343/B -0.00fF
C38086 INVX1_LOC_266/A INVX1_LOC_206/Y 0.00fF
C38087 INVX1_LOC_269/A NOR2X1_LOC_552/Y 0.01fF
C38088 INVX1_LOC_19/A NAND2X1_LOC_74/B 0.38fF
C38089 INVX1_LOC_12/Y INVX1_LOC_29/Y 0.01fF
C38090 INVX1_LOC_19/A NAND2X1_LOC_207/Y 0.02fF
C38091 INVX1_LOC_292/A NOR2X1_LOC_216/Y 0.14fF
C38092 INVX1_LOC_223/A NOR2X1_LOC_180/B 0.00fF
C38093 NAND2X1_LOC_354/B NAND2X1_LOC_840/B 0.28fF
C38094 NAND2X1_LOC_543/Y NAND2X1_LOC_833/Y 0.17fF
C38095 INVX1_LOC_41/A NAND2X1_LOC_392/A 0.01fF
C38096 NOR2X1_LOC_91/Y NAND2X1_LOC_861/Y 0.05fF
C38097 INVX1_LOC_118/A NOR2X1_LOC_438/Y 0.05fF
C38098 INVX1_LOC_214/Y NOR2X1_LOC_52/B 0.03fF
C38099 INVX1_LOC_141/Y INVX1_LOC_140/A 0.05fF
C38100 INVX1_LOC_314/Y INVX1_LOC_10/A 0.01fF
C38101 NAND2X1_LOC_555/Y INVX1_LOC_75/A 0.13fF
C38102 INVX1_LOC_21/A INVX1_LOC_247/A 0.03fF
C38103 NOR2X1_LOC_392/B NOR2X1_LOC_121/A 0.10fF
C38104 INVX1_LOC_191/Y NAND2X1_LOC_451/Y 0.01fF
C38105 INVX1_LOC_30/A NAND2X1_LOC_560/A 0.07fF
C38106 INVX1_LOC_176/A INVX1_LOC_38/Y 0.24fF
C38107 NOR2X1_LOC_791/A NOR2X1_LOC_756/Y 0.10fF
C38108 NOR2X1_LOC_361/B NOR2X1_LOC_318/B 0.05fF
C38109 NAND2X1_LOC_341/A NOR2X1_LOC_367/B 0.25fF
C38110 NAND2X1_LOC_9/Y NOR2X1_LOC_536/A 0.03fF
C38111 NOR2X1_LOC_226/A NOR2X1_LOC_655/B 0.02fF
C38112 INVX1_LOC_223/A INVX1_LOC_73/A 0.07fF
C38113 NOR2X1_LOC_516/B NOR2X1_LOC_802/A 0.10fF
C38114 NOR2X1_LOC_68/A NOR2X1_LOC_19/B 0.03fF
C38115 INVX1_LOC_233/A NOR2X1_LOC_536/A 0.07fF
C38116 NOR2X1_LOC_67/A NAND2X1_LOC_541/Y 0.06fF
C38117 INVX1_LOC_174/Y INVX1_LOC_76/Y 0.27fF
C38118 INVX1_LOC_276/A NAND2X1_LOC_834/a_36_24# 0.00fF
C38119 NOR2X1_LOC_361/B INVX1_LOC_93/Y 0.18fF
C38120 INVX1_LOC_35/A INVX1_LOC_38/A 0.06fF
C38121 INVX1_LOC_289/Y NOR2X1_LOC_56/Y 0.17fF
C38122 INVX1_LOC_200/Y NAND2X1_LOC_241/a_36_24# 0.00fF
C38123 INVX1_LOC_4/Y INVX1_LOC_63/A 0.17fF
C38124 D_INPUT_0 NOR2X1_LOC_551/B 0.00fF
C38125 NOR2X1_LOC_473/B INVX1_LOC_77/A 0.03fF
C38126 NOR2X1_LOC_238/Y INVX1_LOC_28/A 0.06fF
C38127 NOR2X1_LOC_626/Y INVX1_LOC_139/Y 0.01fF
C38128 NOR2X1_LOC_778/B NOR2X1_LOC_500/Y 0.07fF
C38129 INVX1_LOC_209/Y INVX1_LOC_173/Y 0.02fF
C38130 NAND2X1_LOC_112/Y INVX1_LOC_133/Y 0.03fF
C38131 NOR2X1_LOC_620/Y INVX1_LOC_65/Y 0.12fF
C38132 NOR2X1_LOC_498/Y NOR2X1_LOC_525/Y 0.00fF
C38133 INVX1_LOC_64/A NOR2X1_LOC_331/B 0.39fF
C38134 NOR2X1_LOC_690/A NOR2X1_LOC_71/Y 0.01fF
C38135 NOR2X1_LOC_68/A NOR2X1_LOC_589/a_36_216# 0.00fF
C38136 NOR2X1_LOC_635/A NOR2X1_LOC_763/Y 0.03fF
C38137 INVX1_LOC_89/A NAND2X1_LOC_157/a_36_24# 0.00fF
C38138 INVX1_LOC_303/A INVX1_LOC_148/A 0.00fF
C38139 INVX1_LOC_207/A NAND2X1_LOC_866/B 0.08fF
C38140 NOR2X1_LOC_92/Y NAND2X1_LOC_287/B 0.08fF
C38141 NOR2X1_LOC_88/Y NOR2X1_LOC_654/A 0.30fF
C38142 NOR2X1_LOC_15/Y NAND2X1_LOC_650/B 0.11fF
C38143 NAND2X1_LOC_9/Y NAND2X1_LOC_93/B 0.01fF
C38144 INVX1_LOC_49/A INVX1_LOC_182/A 0.22fF
C38145 INVX1_LOC_289/Y VDD 0.87fF
C38146 INVX1_LOC_225/A NOR2X1_LOC_246/a_36_216# 0.09fF
C38147 NOR2X1_LOC_589/A NOR2X1_LOC_366/B 0.03fF
C38148 NAND2X1_LOC_364/A NOR2X1_LOC_734/a_36_216# 0.00fF
C38149 NOR2X1_LOC_810/A NOR2X1_LOC_78/B 0.03fF
C38150 INVX1_LOC_17/A NOR2X1_LOC_309/a_36_216# 0.01fF
C38151 INVX1_LOC_289/Y NAND2X1_LOC_800/A 0.03fF
C38152 INVX1_LOC_33/A NOR2X1_LOC_329/B 0.07fF
C38153 NAND2X1_LOC_190/Y INVX1_LOC_37/A 0.36fF
C38154 NAND2X1_LOC_860/A INVX1_LOC_35/Y 0.00fF
C38155 INVX1_LOC_2/A NOR2X1_LOC_99/B 0.10fF
C38156 INVX1_LOC_136/A INVX1_LOC_125/Y 0.10fF
C38157 INVX1_LOC_90/A INVX1_LOC_257/Y 0.30fF
C38158 INVX1_LOC_17/A NAND2X1_LOC_453/A 0.16fF
C38159 NAND2X1_LOC_363/B NOR2X1_LOC_634/A 0.01fF
C38160 INVX1_LOC_33/A D_INPUT_4 0.01fF
C38161 NOR2X1_LOC_216/Y INVX1_LOC_67/A 0.08fF
C38162 INVX1_LOC_124/A NOR2X1_LOC_473/B 0.01fF
C38163 INVX1_LOC_310/A INVX1_LOC_89/A 0.32fF
C38164 INVX1_LOC_36/A NOR2X1_LOC_595/Y 0.04fF
C38165 NOR2X1_LOC_82/A VDD 1.38fF
C38166 INVX1_LOC_64/A NOR2X1_LOC_592/B 0.03fF
C38167 INVX1_LOC_256/A INVX1_LOC_46/A 0.09fF
C38168 NOR2X1_LOC_742/A INVX1_LOC_153/Y 0.10fF
C38169 NAND2X1_LOC_354/Y NOR2X1_LOC_45/B 0.00fF
C38170 NOR2X1_LOC_589/A NAND2X1_LOC_479/Y 0.00fF
C38171 INVX1_LOC_134/A VDD 0.11fF
C38172 NOR2X1_LOC_68/A NOR2X1_LOC_528/Y -0.01fF
C38173 NOR2X1_LOC_123/B NAND2X1_LOC_850/Y 0.29fF
C38174 NOR2X1_LOC_781/A NAND2X1_LOC_662/Y 0.16fF
C38175 INVX1_LOC_26/Y NAND2X1_LOC_74/B 0.15fF
C38176 INVX1_LOC_41/A NOR2X1_LOC_97/A 0.01fF
C38177 NOR2X1_LOC_798/A NAND2X1_LOC_93/B 0.03fF
C38178 NOR2X1_LOC_742/A INVX1_LOC_121/Y 0.20fF
C38179 NAND2X1_LOC_9/Y INVX1_LOC_3/A 0.18fF
C38180 NOR2X1_LOC_278/Y INVX1_LOC_168/Y 0.01fF
C38181 NAND2X1_LOC_550/A INVX1_LOC_37/Y 0.08fF
C38182 INVX1_LOC_279/A NOR2X1_LOC_665/A 0.01fF
C38183 NAND2X1_LOC_357/B NAND2X1_LOC_863/A 0.01fF
C38184 NOR2X1_LOC_389/A INVX1_LOC_37/A 0.01fF
C38185 NOR2X1_LOC_523/A INVX1_LOC_280/A 0.00fF
C38186 NAND2X1_LOC_722/A NAND2X1_LOC_560/A 0.15fF
C38187 NAND2X1_LOC_652/Y NAND2X1_LOC_661/B 0.00fF
C38188 NOR2X1_LOC_160/B NOR2X1_LOC_363/Y 0.01fF
C38189 NAND2X1_LOC_500/Y VDD 0.11fF
C38190 NAND2X1_LOC_36/A VDD 0.43fF
C38191 INVX1_LOC_135/A NAND2X1_LOC_377/Y 0.03fF
C38192 NOR2X1_LOC_810/A INVX1_LOC_83/A 0.00fF
C38193 INVX1_LOC_102/Y NAND2X1_LOC_850/Y -0.02fF
C38194 NOR2X1_LOC_174/A NOR2X1_LOC_516/B 0.01fF
C38195 NOR2X1_LOC_660/Y INVX1_LOC_19/A -0.00fF
C38196 NOR2X1_LOC_30/a_36_216# INPUT_5 0.00fF
C38197 NAND2X1_LOC_787/A INVX1_LOC_29/A 0.03fF
C38198 NOR2X1_LOC_238/Y NOR2X1_LOC_253/Y 0.01fF
C38199 NOR2X1_LOC_160/B NAND2X1_LOC_276/a_36_24# 0.00fF
C38200 INVX1_LOC_1/A NAND2X1_LOC_435/a_36_24# 0.00fF
C38201 NAND2X1_LOC_350/A INVX1_LOC_118/A 0.48fF
C38202 NAND2X1_LOC_514/Y VDD 0.03fF
C38203 NAND2X1_LOC_363/B INVX1_LOC_29/A 0.11fF
C38204 INVX1_LOC_53/A NOR2X1_LOC_89/A 0.18fF
C38205 NOR2X1_LOC_764/Y INVX1_LOC_83/A 0.00fF
C38206 NAND2X1_LOC_391/Y NAND2X1_LOC_489/Y 0.03fF
C38207 INVX1_LOC_11/A INVX1_LOC_92/A 0.37fF
C38208 NAND2X1_LOC_192/a_36_24# INVX1_LOC_307/A 0.00fF
C38209 NOR2X1_LOC_160/B INVX1_LOC_307/Y 0.05fF
C38210 NOR2X1_LOC_99/B INPUT_1 0.07fF
C38211 NOR2X1_LOC_78/B INVX1_LOC_69/Y 0.01fF
C38212 NOR2X1_LOC_596/A INVX1_LOC_37/A 0.06fF
C38213 NAND2X1_LOC_227/Y NOR2X1_LOC_510/B 0.04fF
C38214 NOR2X1_LOC_441/Y INVX1_LOC_118/A 0.69fF
C38215 INVX1_LOC_182/Y NOR2X1_LOC_665/A 0.00fF
C38216 NAND2X1_LOC_703/Y NOR2X1_LOC_661/A 0.01fF
C38217 NAND2X1_LOC_123/Y INVX1_LOC_10/A 0.01fF
C38218 NOR2X1_LOC_726/Y NOR2X1_LOC_209/B 0.11fF
C38219 INVX1_LOC_236/A INVX1_LOC_91/A 0.02fF
C38220 NOR2X1_LOC_389/A NOR2X1_LOC_743/Y 0.03fF
C38221 NOR2X1_LOC_553/Y NOR2X1_LOC_188/A 0.31fF
C38222 NOR2X1_LOC_791/Y INVX1_LOC_29/A 0.02fF
C38223 NOR2X1_LOC_597/Y INVX1_LOC_10/A 0.01fF
C38224 INVX1_LOC_292/A NOR2X1_LOC_197/B 0.10fF
C38225 INVX1_LOC_285/Y INVX1_LOC_1/Y 0.53fF
C38226 NOR2X1_LOC_501/a_36_216# NOR2X1_LOC_335/B 0.01fF
C38227 NOR2X1_LOC_667/A NOR2X1_LOC_45/B 0.07fF
C38228 NOR2X1_LOC_67/A NOR2X1_LOC_78/A 0.09fF
C38229 NOR2X1_LOC_173/Y INVX1_LOC_272/A 0.18fF
C38230 NOR2X1_LOC_91/A INVX1_LOC_26/A 0.22fF
C38231 INVX1_LOC_2/A INVX1_LOC_291/Y 0.03fF
C38232 INVX1_LOC_248/A NOR2X1_LOC_45/B 0.07fF
C38233 NAND2X1_LOC_672/B INVX1_LOC_315/Y 0.01fF
C38234 INVX1_LOC_72/A INVX1_LOC_185/A 0.03fF
C38235 NAND2X1_LOC_332/Y VDD 0.16fF
C38236 NAND2X1_LOC_570/a_36_24# NAND2X1_LOC_659/B 0.01fF
C38237 NOR2X1_LOC_717/Y INVX1_LOC_179/A 0.00fF
C38238 INVX1_LOC_18/A NOR2X1_LOC_612/Y 0.01fF
C38239 INVX1_LOC_226/Y NOR2X1_LOC_557/A 0.05fF
C38240 NAND2X1_LOC_550/A NOR2X1_LOC_485/Y 0.26fF
C38241 NOR2X1_LOC_790/B NOR2X1_LOC_334/Y 0.03fF
C38242 NOR2X1_LOC_772/B INVX1_LOC_47/Y 0.04fF
C38243 NAND2X1_LOC_515/a_36_24# INVX1_LOC_9/A 0.00fF
C38244 NOR2X1_LOC_112/B INVX1_LOC_120/A 0.00fF
C38245 INVX1_LOC_30/A NOR2X1_LOC_58/Y 0.28fF
C38246 NOR2X1_LOC_360/Y NOR2X1_LOC_79/A 0.02fF
C38247 INVX1_LOC_83/A NOR2X1_LOC_710/a_36_216# 0.02fF
C38248 NOR2X1_LOC_285/A INVX1_LOC_26/Y 0.01fF
C38249 NAND2X1_LOC_477/A NAND2X1_LOC_287/B 0.10fF
C38250 INVX1_LOC_26/A INVX1_LOC_23/A 1.49fF
C38251 NOR2X1_LOC_468/Y NOR2X1_LOC_178/a_36_216# 0.02fF
C38252 INVX1_LOC_143/A INVX1_LOC_143/Y 0.09fF
C38253 INVX1_LOC_13/Y INVX1_LOC_47/Y 0.07fF
C38254 INVX1_LOC_13/A INVX1_LOC_91/A 0.03fF
C38255 NOR2X1_LOC_220/A NOR2X1_LOC_631/B 0.10fF
C38256 NOR2X1_LOC_100/A VDD -0.00fF
C38257 NOR2X1_LOC_68/A NOR2X1_LOC_216/B 0.17fF
C38258 NAND2X1_LOC_803/B INVX1_LOC_49/Y 0.02fF
C38259 NOR2X1_LOC_349/A NAND2X1_LOC_41/Y 0.05fF
C38260 INVX1_LOC_263/A INVX1_LOC_188/Y 0.01fF
C38261 NOR2X1_LOC_778/B NOR2X1_LOC_850/a_36_216# 0.00fF
C38262 INVX1_LOC_50/A INVX1_LOC_57/A 0.22fF
C38263 NOR2X1_LOC_457/A INVX1_LOC_29/A 5.28fF
C38264 INVX1_LOC_95/Y INVX1_LOC_16/A 0.07fF
C38265 INVX1_LOC_161/Y NAND2X1_LOC_74/B 0.07fF
C38266 INVX1_LOC_111/A NOR2X1_LOC_79/Y 0.00fF
C38267 INVX1_LOC_122/Y NAND2X1_LOC_574/A 0.04fF
C38268 NOR2X1_LOC_218/Y NAND2X1_LOC_274/a_36_24# 0.01fF
C38269 NOR2X1_LOC_380/Y NOR2X1_LOC_409/Y 2.50fF
C38270 NOR2X1_LOC_815/Y INVX1_LOC_54/A 0.04fF
C38271 NOR2X1_LOC_590/A INVX1_LOC_49/Y 0.05fF
C38272 NOR2X1_LOC_731/Y VDD 0.26fF
C38273 INVX1_LOC_93/Y NAND2X1_LOC_573/A 0.18fF
C38274 NOR2X1_LOC_220/A INVX1_LOC_37/A 0.01fF
C38275 NAND2X1_LOC_341/A INVX1_LOC_76/A 0.04fF
C38276 INVX1_LOC_136/A NOR2X1_LOC_653/Y 0.03fF
C38277 NOR2X1_LOC_433/A INVX1_LOC_92/A 0.03fF
C38278 INVX1_LOC_257/Y INVX1_LOC_38/A 0.03fF
C38279 INVX1_LOC_278/Y VDD 0.45fF
C38280 INPUT_2 NOR2X1_LOC_14/a_36_216# 0.04fF
C38281 NOR2X1_LOC_204/a_36_216# NOR2X1_LOC_216/B 0.02fF
C38282 INVX1_LOC_21/A NOR2X1_LOC_685/B 0.11fF
C38283 NOR2X1_LOC_226/A NOR2X1_LOC_176/Y 0.01fF
C38284 INVX1_LOC_10/A NOR2X1_LOC_657/B 0.10fF
C38285 NOR2X1_LOC_516/B INVX1_LOC_2/Y 0.04fF
C38286 INVX1_LOC_1/Y NAND2X1_LOC_267/B 0.00fF
C38287 INVX1_LOC_26/Y NOR2X1_LOC_845/a_36_216# 0.00fF
C38288 NOR2X1_LOC_690/A NAND2X1_LOC_243/Y 0.72fF
C38289 NOR2X1_LOC_593/Y INVX1_LOC_92/A 0.03fF
C38290 INPUT_0 INVX1_LOC_67/Y 0.03fF
C38291 NAND2X1_LOC_84/Y NAND2X1_LOC_267/a_36_24# 0.00fF
C38292 NOR2X1_LOC_716/B NOR2X1_LOC_88/Y 0.07fF
C38293 NAND2X1_LOC_463/B NAND2X1_LOC_622/B 0.01fF
C38294 INVX1_LOC_136/A INVX1_LOC_19/A 0.18fF
C38295 INVX1_LOC_5/A NOR2X1_LOC_727/B 0.03fF
C38296 NAND2X1_LOC_550/A NAND2X1_LOC_614/a_36_24# 0.01fF
C38297 INVX1_LOC_34/A NOR2X1_LOC_364/A 0.00fF
C38298 INVX1_LOC_208/A NOR2X1_LOC_363/Y 0.01fF
C38299 NAND2X1_LOC_116/A NAND2X1_LOC_86/a_36_24# 0.01fF
C38300 INVX1_LOC_30/A INVX1_LOC_29/A 6.32fF
C38301 NAND2X1_LOC_555/Y GATE_222 0.02fF
C38302 NOR2X1_LOC_548/Y INVX1_LOC_37/A 1.82fF
C38303 INVX1_LOC_291/Y NAND2X1_LOC_648/A 0.02fF
C38304 INVX1_LOC_171/A NOR2X1_LOC_566/a_36_216# 0.00fF
C38305 INVX1_LOC_269/A INVX1_LOC_253/A 0.01fF
C38306 NAND2X1_LOC_763/B INVX1_LOC_29/A 0.04fF
C38307 INVX1_LOC_141/Y INVX1_LOC_42/A 0.03fF
C38308 INVX1_LOC_135/A INVX1_LOC_20/A 0.67fF
C38309 NOR2X1_LOC_52/B INVX1_LOC_92/A 0.21fF
C38310 INVX1_LOC_157/A INVX1_LOC_46/A 0.05fF
C38311 INVX1_LOC_312/Y INVX1_LOC_42/A 0.19fF
C38312 INVX1_LOC_135/A NOR2X1_LOC_360/A 0.01fF
C38313 INVX1_LOC_63/Y NOR2X1_LOC_697/Y 0.06fF
C38314 INVX1_LOC_222/Y NOR2X1_LOC_748/A 0.03fF
C38315 NOR2X1_LOC_716/B INVX1_LOC_84/A 0.14fF
C38316 VDD INVX1_LOC_306/A 0.19fF
C38317 NAND2X1_LOC_549/Y NAND2X1_LOC_569/B 0.01fF
C38318 NOR2X1_LOC_378/a_36_216# NAND2X1_LOC_93/B 0.00fF
C38319 INVX1_LOC_34/A INVX1_LOC_285/A 0.07fF
C38320 INVX1_LOC_36/A NAND2X1_LOC_214/a_36_24# 0.00fF
C38321 NAND2X1_LOC_222/A NAND2X1_LOC_218/A 0.01fF
C38322 NAND2X1_LOC_51/B NOR2X1_LOC_45/B 0.00fF
C38323 NOR2X1_LOC_231/a_36_216# INVX1_LOC_15/A 0.01fF
C38324 INVX1_LOC_217/A NAND2X1_LOC_254/Y 0.05fF
C38325 INVX1_LOC_34/A NOR2X1_LOC_814/A 0.03fF
C38326 NOR2X1_LOC_355/A INVX1_LOC_12/Y 0.01fF
C38327 NOR2X1_LOC_378/a_36_216# NAND2X1_LOC_425/Y 0.01fF
C38328 NOR2X1_LOC_778/B INVX1_LOC_307/A 0.14fF
C38329 NAND2X1_LOC_181/Y INVX1_LOC_70/A 0.03fF
C38330 NOR2X1_LOC_708/B NAND2X1_LOC_782/B 0.20fF
C38331 INVX1_LOC_314/Y INVX1_LOC_12/A 0.03fF
C38332 NOR2X1_LOC_318/B INVX1_LOC_285/Y 0.10fF
C38333 NOR2X1_LOC_333/A INVX1_LOC_117/A 0.01fF
C38334 INVX1_LOC_28/A NOR2X1_LOC_305/Y 0.07fF
C38335 INVX1_LOC_50/A NOR2X1_LOC_666/Y 0.00fF
C38336 NOR2X1_LOC_778/B NOR2X1_LOC_445/B 0.08fF
C38337 INVX1_LOC_206/Y INVX1_LOC_96/A 0.03fF
C38338 INVX1_LOC_6/A NOR2X1_LOC_269/Y 0.07fF
C38339 NOR2X1_LOC_666/A INVX1_LOC_23/A 0.01fF
C38340 NOR2X1_LOC_111/Y NAND2X1_LOC_211/Y 0.05fF
C38341 INVX1_LOC_89/A NAND2X1_LOC_96/A 0.14fF
C38342 NOR2X1_LOC_551/Y NOR2X1_LOC_78/A 0.02fF
C38343 INVX1_LOC_65/Y INVX1_LOC_117/A 0.04fF
C38344 NAND2X1_LOC_740/B INVX1_LOC_76/A 0.13fF
C38345 NAND2X1_LOC_231/Y INVX1_LOC_285/A 0.10fF
C38346 INVX1_LOC_5/A NOR2X1_LOC_649/Y 0.12fF
C38347 NAND2X1_LOC_354/B INVX1_LOC_49/Y 0.06fF
C38348 NOR2X1_LOC_256/Y INVX1_LOC_76/A 0.06fF
C38349 D_GATE_366 INVX1_LOC_117/A 0.07fF
C38350 NAND2X1_LOC_348/A NOR2X1_LOC_347/a_36_216# 0.00fF
C38351 INPUT_5 INVX1_LOC_54/A 0.43fF
C38352 INVX1_LOC_272/Y INVX1_LOC_271/A 0.02fF
C38353 NOR2X1_LOC_216/Y NOR2X1_LOC_137/Y 0.03fF
C38354 NAND2X1_LOC_841/a_36_24# INVX1_LOC_199/A 0.01fF
C38355 INVX1_LOC_312/Y INVX1_LOC_78/A 0.07fF
C38356 INVX1_LOC_93/Y NOR2X1_LOC_183/a_36_216# -0.01fF
C38357 NAND2X1_LOC_53/Y INVX1_LOC_105/Y 0.01fF
C38358 INVX1_LOC_96/A NOR2X1_LOC_600/Y 0.00fF
C38359 NAND2X1_LOC_842/B NOR2X1_LOC_536/A 0.01fF
C38360 INVX1_LOC_75/A NOR2X1_LOC_706/B 0.03fF
C38361 NOR2X1_LOC_473/B INVX1_LOC_9/A 0.09fF
C38362 NOR2X1_LOC_772/a_36_216# INVX1_LOC_285/A 0.13fF
C38363 NAND2X1_LOC_483/Y INVX1_LOC_42/A 0.00fF
C38364 INVX1_LOC_11/A INVX1_LOC_53/A 0.51fF
C38365 NOR2X1_LOC_419/Y INVX1_LOC_15/A 0.03fF
C38366 INVX1_LOC_303/A INVX1_LOC_47/Y 0.04fF
C38367 NOR2X1_LOC_160/B INVX1_LOC_29/Y 0.03fF
C38368 INVX1_LOC_285/Y INVX1_LOC_139/A 0.12fF
C38369 INVX1_LOC_27/A NAND2X1_LOC_474/Y 0.10fF
C38370 NOR2X1_LOC_848/Y INVX1_LOC_64/A 0.00fF
C38371 NOR2X1_LOC_45/B INVX1_LOC_304/A 0.12fF
C38372 INVX1_LOC_61/Y INVX1_LOC_57/A 0.07fF
C38373 NAND2X1_LOC_347/B NOR2X1_LOC_81/Y 0.07fF
C38374 INVX1_LOC_69/Y INVX1_LOC_46/A 0.07fF
C38375 NOR2X1_LOC_716/B INVX1_LOC_15/A 0.07fF
C38376 NOR2X1_LOC_65/B INVX1_LOC_312/Y 0.00fF
C38377 NOR2X1_LOC_655/B NAND2X1_LOC_63/Y 0.05fF
C38378 INVX1_LOC_233/A INVX1_LOC_256/A 0.01fF
C38379 INVX1_LOC_293/A NOR2X1_LOC_392/Y 0.01fF
C38380 INVX1_LOC_277/Y NOR2X1_LOC_383/B 0.02fF
C38381 NOR2X1_LOC_332/A NOR2X1_LOC_820/a_36_216# 0.01fF
C38382 NAND2X1_LOC_549/Y NOR2X1_LOC_530/Y 0.27fF
C38383 NOR2X1_LOC_501/a_36_216# INVX1_LOC_84/A 0.00fF
C38384 NOR2X1_LOC_763/A NOR2X1_LOC_582/A 0.06fF
C38385 INVX1_LOC_2/Y INVX1_LOC_315/Y 0.44fF
C38386 NOR2X1_LOC_388/Y INVX1_LOC_4/A 0.03fF
C38387 INVX1_LOC_311/A INVX1_LOC_281/A 0.08fF
C38388 NOR2X1_LOC_724/Y INVX1_LOC_307/A 0.02fF
C38389 NOR2X1_LOC_360/Y INVX1_LOC_28/Y 0.06fF
C38390 NOR2X1_LOC_78/B NOR2X1_LOC_89/A 0.19fF
C38391 NOR2X1_LOC_78/A NOR2X1_LOC_558/A 0.01fF
C38392 NAND2X1_LOC_9/Y NOR2X1_LOC_606/Y 0.28fF
C38393 INVX1_LOC_136/A NAND2X1_LOC_557/Y -0.00fF
C38394 INVX1_LOC_30/A NOR2X1_LOC_843/a_36_216# 0.00fF
C38395 NOR2X1_LOC_344/A NOR2X1_LOC_334/Y 0.01fF
C38396 NOR2X1_LOC_717/B INVX1_LOC_84/A 0.03fF
C38397 INVX1_LOC_45/A INPUT_6 0.01fF
C38398 INVX1_LOC_93/Y NAND2X1_LOC_267/B 0.03fF
C38399 INVX1_LOC_256/A NOR2X1_LOC_798/A 0.03fF
C38400 NAND2X1_LOC_807/A NOR2X1_LOC_652/Y 0.04fF
C38401 NOR2X1_LOC_242/A INVX1_LOC_11/A 3.45fF
C38402 NAND2X1_LOC_531/a_36_24# INVX1_LOC_84/A 0.00fF
C38403 NAND2X1_LOC_35/Y INVX1_LOC_284/Y 2.86fF
C38404 NAND2X1_LOC_53/Y INVX1_LOC_27/A 1.77fF
C38405 D_INPUT_0 NOR2X1_LOC_691/A 0.04fF
C38406 INVX1_LOC_24/A NOR2X1_LOC_677/Y 0.01fF
C38407 INVX1_LOC_229/A NAND2X1_LOC_579/A 0.00fF
C38408 NOR2X1_LOC_360/Y NOR2X1_LOC_416/A 0.02fF
C38409 NAND2X1_LOC_787/A NAND2X1_LOC_634/Y 0.02fF
C38410 INVX1_LOC_92/Y INVX1_LOC_9/A 0.01fF
C38411 NOR2X1_LOC_349/A INVX1_LOC_122/A 0.09fF
C38412 NOR2X1_LOC_78/B NOR2X1_LOC_170/A 0.02fF
C38413 NOR2X1_LOC_130/Y INVX1_LOC_84/A 0.01fF
C38414 NOR2X1_LOC_746/Y INVX1_LOC_117/A 0.02fF
C38415 VDD INVX1_LOC_59/Y 1.39fF
C38416 INVX1_LOC_112/A VDD 0.24fF
C38417 NOR2X1_LOC_658/Y INVX1_LOC_5/A 0.04fF
C38418 INVX1_LOC_144/A INVX1_LOC_180/Y 0.01fF
C38419 INVX1_LOC_282/A NOR2X1_LOC_491/Y 0.03fF
C38420 NOR2X1_LOC_272/a_36_216# NOR2X1_LOC_441/Y 0.00fF
C38421 NAND2X1_LOC_390/A INVX1_LOC_102/A 0.02fF
C38422 NOR2X1_LOC_789/A INVX1_LOC_42/A 0.00fF
C38423 NOR2X1_LOC_355/B INVX1_LOC_9/A 0.15fF
C38424 NAND2X1_LOC_392/Y NOR2X1_LOC_89/A 0.35fF
C38425 NOR2X1_LOC_99/B NAND2X1_LOC_63/Y 0.14fF
C38426 INVX1_LOC_176/A VDD 0.44fF
C38427 INVX1_LOC_41/Y NAND2X1_LOC_793/B 0.30fF
C38428 NOR2X1_LOC_503/A INVX1_LOC_84/A 0.09fF
C38429 NAND2X1_LOC_741/Y NAND2X1_LOC_741/B 0.02fF
C38430 NOR2X1_LOC_78/A NOR2X1_LOC_729/A 0.03fF
C38431 INVX1_LOC_83/A NOR2X1_LOC_89/A 0.12fF
C38432 INVX1_LOC_131/A NOR2X1_LOC_814/A 0.02fF
C38433 NOR2X1_LOC_398/a_36_216# INVX1_LOC_23/Y 0.01fF
C38434 NOR2X1_LOC_433/A INVX1_LOC_53/A 1.19fF
C38435 NOR2X1_LOC_447/B INVX1_LOC_37/A 0.00fF
C38436 NOR2X1_LOC_813/Y INVX1_LOC_20/A 0.42fF
C38437 NOR2X1_LOC_151/Y INVX1_LOC_84/A 0.03fF
C38438 NOR2X1_LOC_220/A NAND2X1_LOC_72/B 0.33fF
C38439 INPUT_0 INVX1_LOC_285/A 0.14fF
C38440 NOR2X1_LOC_363/Y NAND2X1_LOC_211/Y 0.01fF
C38441 NOR2X1_LOC_451/A INVX1_LOC_91/A 0.14fF
C38442 NOR2X1_LOC_593/Y INVX1_LOC_53/A 0.07fF
C38443 INVX1_LOC_44/A INVX1_LOC_76/A 0.02fF
C38444 NOR2X1_LOC_773/a_36_216# INVX1_LOC_57/A 0.00fF
C38445 NOR2X1_LOC_613/a_36_216# INVX1_LOC_217/A 0.01fF
C38446 INPUT_0 INVX1_LOC_265/Y 0.00fF
C38447 INVX1_LOC_278/A NOR2X1_LOC_716/B 0.17fF
C38448 INVX1_LOC_5/A NOR2X1_LOC_13/Y 0.01fF
C38449 INVX1_LOC_22/A NOR2X1_LOC_158/B 0.02fF
C38450 INVX1_LOC_1/Y INVX1_LOC_4/Y 0.06fF
C38451 INVX1_LOC_280/A INVX1_LOC_20/A 0.10fF
C38452 INPUT_0 NOR2X1_LOC_814/A 0.17fF
C38453 NOR2X1_LOC_94/Y INVX1_LOC_20/A 0.24fF
C38454 INVX1_LOC_35/A INVX1_LOC_33/A 0.50fF
C38455 NOR2X1_LOC_540/a_36_216# NOR2X1_LOC_334/Y 0.01fF
C38456 INVX1_LOC_16/A INVX1_LOC_271/Y 0.09fF
C38457 NOR2X1_LOC_459/a_36_216# NOR2X1_LOC_476/B 0.00fF
C38458 NAND2X1_LOC_349/B INVX1_LOC_94/Y 0.47fF
C38459 INVX1_LOC_269/A NOR2X1_LOC_336/B 0.01fF
C38460 INVX1_LOC_35/A NOR2X1_LOC_743/a_36_216# 0.00fF
C38461 NAND2X1_LOC_212/Y INVX1_LOC_54/A 0.02fF
C38462 NOR2X1_LOC_360/A INVX1_LOC_280/A 0.06fF
C38463 INVX1_LOC_22/A NOR2X1_LOC_30/Y 0.12fF
C38464 NOR2X1_LOC_180/B INVX1_LOC_290/Y 0.03fF
C38465 NOR2X1_LOC_717/B INVX1_LOC_15/A 0.06fF
C38466 NAND2X1_LOC_363/B INVX1_LOC_8/A 0.07fF
C38467 INVX1_LOC_157/Y NAND2X1_LOC_469/B 0.00fF
C38468 NOR2X1_LOC_567/B NOR2X1_LOC_633/A 0.02fF
C38469 NOR2X1_LOC_548/Y NAND2X1_LOC_72/B 0.01fF
C38470 NOR2X1_LOC_324/B INVX1_LOC_307/Y 0.15fF
C38471 NOR2X1_LOC_52/B INVX1_LOC_53/A 6.59fF
C38472 INVX1_LOC_199/A INVX1_LOC_92/A 0.02fF
C38473 INVX1_LOC_135/A INVX1_LOC_4/A 0.07fF
C38474 NOR2X1_LOC_597/Y INVX1_LOC_12/A 0.01fF
C38475 INVX1_LOC_309/A NAND2X1_LOC_489/Y 0.00fF
C38476 INVX1_LOC_269/A NAND2X1_LOC_364/A 0.05fF
C38477 INVX1_LOC_71/A NOR2X1_LOC_440/B 0.10fF
C38478 NOR2X1_LOC_745/a_36_216# INVX1_LOC_30/A 0.00fF
C38479 NAND2X1_LOC_376/a_36_24# INVX1_LOC_175/A 0.00fF
C38480 NOR2X1_LOC_468/Y NAND2X1_LOC_198/B 0.10fF
C38481 INVX1_LOC_25/Y INVX1_LOC_181/A 0.07fF
C38482 NOR2X1_LOC_828/A INVX1_LOC_15/A 0.05fF
C38483 NOR2X1_LOC_361/B NAND2X1_LOC_514/Y 0.05fF
C38484 INVX1_LOC_41/A INVX1_LOC_50/Y 0.14fF
C38485 NAND2X1_LOC_656/Y INVX1_LOC_78/A 0.03fF
C38486 INVX1_LOC_136/A INVX1_LOC_161/Y 0.10fF
C38487 NAND2X1_LOC_348/A NAND2X1_LOC_206/B 0.09fF
C38488 INVX1_LOC_73/A INVX1_LOC_290/Y 0.07fF
C38489 NAND2X1_LOC_387/B INVX1_LOC_174/A 0.04fF
C38490 NOR2X1_LOC_510/Y NAND2X1_LOC_332/Y 0.02fF
C38491 NOR2X1_LOC_791/Y INVX1_LOC_8/A 0.05fF
C38492 INVX1_LOC_208/A INVX1_LOC_29/Y 0.08fF
C38493 NAND2X1_LOC_378/a_36_24# INVX1_LOC_175/A 0.00fF
C38494 NOR2X1_LOC_219/B NOR2X1_LOC_215/A 0.18fF
C38495 INVX1_LOC_21/A NAND2X1_LOC_115/a_36_24# 0.00fF
C38496 NOR2X1_LOC_518/Y NOR2X1_LOC_816/A 0.01fF
C38497 NAND2X1_LOC_297/a_36_24# NOR2X1_LOC_271/Y 0.00fF
C38498 INVX1_LOC_35/A INVX1_LOC_120/Y 0.02fF
C38499 NOR2X1_LOC_773/Y NOR2X1_LOC_717/A 0.00fF
C38500 NAND2X1_LOC_724/A NOR2X1_LOC_753/Y 0.07fF
C38501 NAND2X1_LOC_76/a_36_24# INVX1_LOC_18/A 0.00fF
C38502 INVX1_LOC_220/Y NOR2X1_LOC_748/A 0.11fF
C38503 NOR2X1_LOC_151/Y INVX1_LOC_15/A 0.08fF
C38504 INVX1_LOC_64/A NOR2X1_LOC_366/B 0.29fF
C38505 NOR2X1_LOC_65/B NAND2X1_LOC_656/Y 0.01fF
C38506 INVX1_LOC_249/A NAND2X1_LOC_53/Y 0.10fF
C38507 NOR2X1_LOC_820/A INVX1_LOC_31/A 0.05fF
C38508 NOR2X1_LOC_225/a_36_216# INVX1_LOC_181/Y 0.00fF
C38509 INVX1_LOC_79/A INVX1_LOC_32/A 0.01fF
C38510 INVX1_LOC_45/A INVX1_LOC_142/A 0.06fF
C38511 NOR2X1_LOC_230/Y INVX1_LOC_72/A 0.04fF
C38512 INVX1_LOC_17/A NOR2X1_LOC_577/Y 0.09fF
C38513 INVX1_LOC_46/A INVX1_LOC_297/A 3.66fF
C38514 NOR2X1_LOC_332/A NOR2X1_LOC_105/a_36_216# 0.01fF
C38515 INVX1_LOC_136/A NOR2X1_LOC_599/A 0.06fF
C38516 INVX1_LOC_10/A INVX1_LOC_271/A 0.44fF
C38517 INVX1_LOC_202/Y NOR2X1_LOC_155/A 0.01fF
C38518 NOR2X1_LOC_790/B NOR2X1_LOC_569/Y 0.13fF
C38519 NOR2X1_LOC_78/A NOR2X1_LOC_327/a_36_216# 0.00fF
C38520 INVX1_LOC_93/Y NAND2X1_LOC_81/B 0.07fF
C38521 NOR2X1_LOC_294/Y NOR2X1_LOC_554/B 0.20fF
C38522 NOR2X1_LOC_437/Y NOR2X1_LOC_276/Y 0.00fF
C38523 NAND2X1_LOC_182/A NOR2X1_LOC_15/Y 0.03fF
C38524 NAND2X1_LOC_218/B NAND2X1_LOC_555/Y 0.14fF
C38525 NAND2X1_LOC_243/B NOR2X1_LOC_536/A 0.05fF
C38526 NOR2X1_LOC_15/Y INVX1_LOC_104/A 0.08fF
C38527 NOR2X1_LOC_82/A NOR2X1_LOC_132/Y 0.03fF
C38528 INVX1_LOC_75/A INVX1_LOC_94/Y 0.03fF
C38529 NAND2X1_LOC_347/B NOR2X1_LOC_709/A 0.07fF
C38530 NAND2X1_LOC_357/A INVX1_LOC_162/A 0.16fF
C38531 NOR2X1_LOC_657/B INVX1_LOC_12/A 0.28fF
C38532 NOR2X1_LOC_766/Y INVX1_LOC_297/A 0.03fF
C38533 NOR2X1_LOC_290/a_36_216# NAND2X1_LOC_489/Y 0.00fF
C38534 NAND2X1_LOC_175/B NOR2X1_LOC_816/A 0.16fF
C38535 INVX1_LOC_2/A NAND2X1_LOC_579/A 0.01fF
C38536 NAND2X1_LOC_357/B INVX1_LOC_308/Y 0.03fF
C38537 NOR2X1_LOC_32/B D_INPUT_0 0.48fF
C38538 NOR2X1_LOC_456/Y INVX1_LOC_97/A 0.04fF
C38539 NOR2X1_LOC_45/B INVX1_LOC_19/Y 0.03fF
C38540 NOR2X1_LOC_89/A NOR2X1_LOC_368/Y 0.13fF
C38541 INVX1_LOC_226/Y INVX1_LOC_27/A 0.08fF
C38542 INVX1_LOC_58/A D_GATE_366 0.07fF
C38543 INVX1_LOC_45/A NAND2X1_LOC_593/Y 0.05fF
C38544 NOR2X1_LOC_226/A NAND2X1_LOC_579/A 0.10fF
C38545 INVX1_LOC_32/A INVX1_LOC_91/A 3.25fF
C38546 NOR2X1_LOC_536/A INVX1_LOC_119/Y 0.09fF
C38547 INVX1_LOC_266/A NOR2X1_LOC_405/a_36_216# 0.00fF
C38548 NOR2X1_LOC_456/Y INVX1_LOC_90/A 0.07fF
C38549 INVX1_LOC_34/A NOR2X1_LOC_590/A 0.03fF
C38550 NAND2X1_LOC_391/Y NAND2X1_LOC_564/B 0.37fF
C38551 INVX1_LOC_64/A INVX1_LOC_135/A 0.22fF
C38552 INVX1_LOC_2/Y NAND2X1_LOC_207/B 0.74fF
C38553 NAND2X1_LOC_35/Y NOR2X1_LOC_525/Y 0.01fF
C38554 INVX1_LOC_31/A INVX1_LOC_315/A 0.07fF
C38555 NOR2X1_LOC_440/Y NOR2X1_LOC_798/A 0.00fF
C38556 VDD NOR2X1_LOC_340/A 0.18fF
C38557 INVX1_LOC_222/A NOR2X1_LOC_541/B 0.07fF
C38558 INVX1_LOC_59/A INVX1_LOC_16/A 0.01fF
C38559 INVX1_LOC_161/Y NOR2X1_LOC_111/a_36_216# 0.01fF
C38560 NOR2X1_LOC_810/A NOR2X1_LOC_798/A 0.03fF
C38561 NOR2X1_LOC_91/A NOR2X1_LOC_368/A 0.46fF
C38562 INVX1_LOC_78/Y INVX1_LOC_78/A 0.01fF
C38563 INVX1_LOC_36/A INVX1_LOC_207/A 0.14fF
C38564 NOR2X1_LOC_15/Y INVX1_LOC_263/A 0.02fF
C38565 NOR2X1_LOC_552/A INVX1_LOC_4/A 0.07fF
C38566 INVX1_LOC_17/A NOR2X1_LOC_346/B 0.38fF
C38567 NOR2X1_LOC_91/A NOR2X1_LOC_313/Y 0.05fF
C38568 NOR2X1_LOC_318/B INVX1_LOC_4/Y 1.25fF
C38569 NOR2X1_LOC_89/A INVX1_LOC_46/A 0.25fF
C38570 INVX1_LOC_11/A NOR2X1_LOC_547/B 0.01fF
C38571 INVX1_LOC_11/A NOR2X1_LOC_78/B 0.39fF
C38572 NOR2X1_LOC_332/A NOR2X1_LOC_649/Y 0.03fF
C38573 NOR2X1_LOC_181/A INVX1_LOC_15/A 0.01fF
C38574 INVX1_LOC_6/A INVX1_LOC_26/A 5.09fF
C38575 NOR2X1_LOC_468/Y INVX1_LOC_53/Y 1.29fF
C38576 NOR2X1_LOC_454/Y NOR2X1_LOC_781/A 0.01fF
C38577 NAND2X1_LOC_581/Y NAND2X1_LOC_36/A 0.04fF
C38578 INVX1_LOC_41/Y INVX1_LOC_71/A 0.00fF
C38579 INVX1_LOC_30/A INVX1_LOC_8/A 0.12fF
C38580 INVX1_LOC_27/A INVX1_LOC_10/A 0.47fF
C38581 INVX1_LOC_11/A NAND2X1_LOC_588/a_36_24# 0.00fF
C38582 NOR2X1_LOC_146/a_36_216# NAND2X1_LOC_425/Y 0.01fF
C38583 INVX1_LOC_93/Y INVX1_LOC_4/Y 0.26fF
C38584 INVX1_LOC_39/A NOR2X1_LOC_99/B -0.00fF
C38585 INVX1_LOC_255/Y INVX1_LOC_14/A 0.16fF
C38586 INVX1_LOC_33/A NOR2X1_LOC_325/Y 0.02fF
C38587 INVX1_LOC_91/A NAND2X1_LOC_175/Y 0.15fF
C38588 NOR2X1_LOC_590/A NAND2X1_LOC_231/Y 0.03fF
C38589 INVX1_LOC_17/A INVX1_LOC_22/A 0.18fF
C38590 NOR2X1_LOC_368/A INVX1_LOC_23/A 0.04fF
C38591 INVX1_LOC_222/Y INVX1_LOC_89/A 0.03fF
C38592 NOR2X1_LOC_15/Y NAND2X1_LOC_854/B 0.05fF
C38593 INVX1_LOC_71/Y INVX1_LOC_84/A 0.05fF
C38594 NOR2X1_LOC_232/Y NOR2X1_LOC_86/A 0.15fF
C38595 NOR2X1_LOC_837/B INVX1_LOC_33/A 0.00fF
C38596 NOR2X1_LOC_536/A INVX1_LOC_284/A 0.22fF
C38597 NAND2X1_LOC_633/Y INVX1_LOC_15/A 0.07fF
C38598 INVX1_LOC_224/Y NOR2X1_LOC_368/a_36_216# 0.01fF
C38599 NAND2X1_LOC_564/A INVX1_LOC_6/A 0.01fF
C38600 NOR2X1_LOC_361/B NOR2X1_LOC_236/a_36_216# 0.13fF
C38601 NOR2X1_LOC_363/Y NAND2X1_LOC_791/a_36_24# 0.00fF
C38602 NOR2X1_LOC_122/a_36_216# INVX1_LOC_290/Y 0.01fF
C38603 INVX1_LOC_11/Y NAND2X1_LOC_175/Y 1.23fF
C38604 NOR2X1_LOC_533/A INVX1_LOC_286/Y 0.03fF
C38605 INVX1_LOC_106/A INVX1_LOC_9/A 0.01fF
C38606 NOR2X1_LOC_471/Y INVX1_LOC_22/A 0.11fF
C38607 NOR2X1_LOC_219/Y NOR2X1_LOC_389/A 0.06fF
C38608 INVX1_LOC_90/A NAND2X1_LOC_714/B 0.01fF
C38609 INVX1_LOC_41/A NOR2X1_LOC_559/B 0.01fF
C38610 INVX1_LOC_36/A NAND2X1_LOC_451/Y 0.03fF
C38611 NOR2X1_LOC_35/Y INVX1_LOC_271/Y 0.10fF
C38612 NOR2X1_LOC_160/B NOR2X1_LOC_160/Y 0.18fF
C38613 NOR2X1_LOC_389/A INVX1_LOC_53/Y 0.09fF
C38614 NAND2X1_LOC_222/B INVX1_LOC_83/A -0.00fF
C38615 INVX1_LOC_216/Y INVX1_LOC_80/A 0.10fF
C38616 INVX1_LOC_14/A NOR2X1_LOC_71/Y 0.14fF
C38617 INVX1_LOC_49/A NOR2X1_LOC_551/B 0.18fF
C38618 NAND2X1_LOC_366/A NAND2X1_LOC_364/Y 0.06fF
C38619 INVX1_LOC_224/A INVX1_LOC_83/A 0.11fF
C38620 NOR2X1_LOC_340/A NAND2X1_LOC_41/a_36_24# 0.00fF
C38621 NAND2X1_LOC_63/Y NOR2X1_LOC_622/a_36_216# 0.01fF
C38622 INVX1_LOC_27/A NOR2X1_LOC_302/Y 0.02fF
C38623 NAND2X1_LOC_267/B INVX1_LOC_87/A 0.02fF
C38624 INVX1_LOC_11/A INVX1_LOC_83/A 0.59fF
C38625 NOR2X1_LOC_215/Y INVX1_LOC_96/Y 0.01fF
C38626 NOR2X1_LOC_468/Y NOR2X1_LOC_76/a_36_216# 0.01fF
C38627 NOR2X1_LOC_57/a_36_216# INVX1_LOC_4/A 0.02fF
C38628 INVX1_LOC_5/A NOR2X1_LOC_337/A 0.03fF
C38629 NOR2X1_LOC_238/Y NOR2X1_LOC_482/Y 0.03fF
C38630 INVX1_LOC_103/A INVX1_LOC_190/Y 0.03fF
C38631 NOR2X1_LOC_315/Y NOR2X1_LOC_373/a_36_216# 0.00fF
C38632 NOR2X1_LOC_355/A NOR2X1_LOC_160/B 0.03fF
C38633 INVX1_LOC_240/A NAND2X1_LOC_486/a_36_24# 0.06fF
C38634 INVX1_LOC_280/A INVX1_LOC_4/A 0.01fF
C38635 INVX1_LOC_203/A NAND2X1_LOC_489/Y 0.15fF
C38636 NOR2X1_LOC_841/A NAND2X1_LOC_74/B 0.07fF
C38637 INVX1_LOC_41/A NOR2X1_LOC_6/B 1.81fF
C38638 INVX1_LOC_205/Y INVX1_LOC_75/A 0.04fF
C38639 NAND2X1_LOC_833/Y NAND2X1_LOC_650/a_36_24# 0.01fF
C38640 INVX1_LOC_201/Y NOR2X1_LOC_6/B 0.06fF
C38641 NAND2X1_LOC_563/Y NAND2X1_LOC_139/A 0.02fF
C38642 NOR2X1_LOC_656/a_36_216# INVX1_LOC_255/Y 0.00fF
C38643 INVX1_LOC_299/A INVX1_LOC_75/A 0.16fF
C38644 INVX1_LOC_64/A NOR2X1_LOC_552/A 0.07fF
C38645 NAND2X1_LOC_741/B NOR2X1_LOC_298/Y 0.03fF
C38646 NOR2X1_LOC_78/B NOR2X1_LOC_433/A 3.41fF
C38647 NOR2X1_LOC_792/B NOR2X1_LOC_309/Y 0.00fF
C38648 NOR2X1_LOC_619/A INVX1_LOC_62/Y 0.11fF
C38649 NOR2X1_LOC_422/Y INVX1_LOC_296/Y 0.01fF
C38650 INVX1_LOC_24/A INVX1_LOC_56/Y 0.01fF
C38651 D_INPUT_3 NAND2X1_LOC_215/A 0.06fF
C38652 NOR2X1_LOC_78/B NOR2X1_LOC_593/Y 0.03fF
C38653 NAND2X1_LOC_577/A INVX1_LOC_89/A 0.07fF
C38654 INVX1_LOC_284/A INVX1_LOC_3/A 0.07fF
C38655 NOR2X1_LOC_570/Y NOR2X1_LOC_303/Y 0.09fF
C38656 NOR2X1_LOC_596/A NOR2X1_LOC_665/A 0.06fF
C38657 NOR2X1_LOC_666/A INVX1_LOC_6/A 0.01fF
C38658 NAND2X1_LOC_861/a_36_24# INVX1_LOC_71/A 0.00fF
C38659 NAND2X1_LOC_99/Y INVX1_LOC_226/Y 0.03fF
C38660 INVX1_LOC_208/Y INVX1_LOC_49/A 0.00fF
C38661 INVX1_LOC_305/Y INVX1_LOC_33/A 0.02fF
C38662 INVX1_LOC_46/A NAND2X1_LOC_804/A 0.01fF
C38663 INVX1_LOC_215/A NOR2X1_LOC_106/Y 0.17fF
C38664 NAND2X1_LOC_35/B INVX1_LOC_240/A 0.41fF
C38665 NOR2X1_LOC_15/Y INVX1_LOC_206/Y 5.39fF
C38666 INVX1_LOC_258/Y NOR2X1_LOC_45/B 0.03fF
C38667 NOR2X1_LOC_590/A INVX1_LOC_131/A 0.00fF
C38668 NOR2X1_LOC_78/B NOR2X1_LOC_52/B 0.29fF
C38669 INVX1_LOC_54/Y NAND2X1_LOC_134/a_36_24# 0.00fF
C38670 INVX1_LOC_34/A NOR2X1_LOC_82/Y 0.03fF
C38671 INVX1_LOC_45/A NOR2X1_LOC_535/a_36_216# 0.00fF
C38672 INVX1_LOC_45/Y NOR2X1_LOC_137/A 0.06fF
C38673 INVX1_LOC_6/Y INVX1_LOC_10/A 0.04fF
C38674 NOR2X1_LOC_569/Y NOR2X1_LOC_344/A 0.02fF
C38675 INVX1_LOC_13/A NAND2X1_LOC_276/Y 0.03fF
C38676 INVX1_LOC_255/Y INVX1_LOC_217/Y 0.01fF
C38677 NOR2X1_LOC_459/A NOR2X1_LOC_474/A 0.09fF
C38678 INVX1_LOC_89/A NAND2X1_LOC_656/A 0.20fF
C38679 NOR2X1_LOC_6/B NOR2X1_LOC_211/A 0.04fF
C38680 NOR2X1_LOC_590/A INPUT_0 10.72fF
C38681 NOR2X1_LOC_315/Y INVX1_LOC_25/Y 0.20fF
C38682 INVX1_LOC_83/A NOR2X1_LOC_433/A 0.10fF
C38683 NOR2X1_LOC_15/Y NOR2X1_LOC_600/Y 0.01fF
C38684 NOR2X1_LOC_603/a_36_216# NOR2X1_LOC_78/B 0.00fF
C38685 NOR2X1_LOC_456/Y INVX1_LOC_38/A 0.08fF
C38686 INVX1_LOC_64/A NOR2X1_LOC_813/Y 0.02fF
C38687 NOR2X1_LOC_32/B NAND2X1_LOC_848/A 0.03fF
C38688 NOR2X1_LOC_742/A NOR2X1_LOC_723/Y 0.03fF
C38689 INVX1_LOC_206/A NOR2X1_LOC_500/Y 0.01fF
C38690 INVX1_LOC_22/Y INPUT_0 0.82fF
C38691 NAND2X1_LOC_794/B NOR2X1_LOC_305/Y 0.00fF
C38692 INVX1_LOC_269/A NOR2X1_LOC_405/A 0.07fF
C38693 NOR2X1_LOC_286/Y NOR2X1_LOC_78/A 0.01fF
C38694 INVX1_LOC_34/A INVX1_LOC_227/A 0.07fF
C38695 NOR2X1_LOC_550/B INVX1_LOC_97/A 0.09fF
C38696 INVX1_LOC_11/A NOR2X1_LOC_311/Y 0.02fF
C38697 NOR2X1_LOC_383/B INVX1_LOC_179/A 0.03fF
C38698 INVX1_LOC_64/A INVX1_LOC_280/A 0.08fF
C38699 INVX1_LOC_308/A INVX1_LOC_118/A 0.03fF
C38700 NOR2X1_LOC_468/Y NAND2X1_LOC_465/A 0.01fF
C38701 INVX1_LOC_90/A NOR2X1_LOC_550/B 0.06fF
C38702 INVX1_LOC_64/A NOR2X1_LOC_94/Y 0.01fF
C38703 INVX1_LOC_120/A NAND2X1_LOC_135/a_36_24# 0.00fF
C38704 INVX1_LOC_278/A NOR2X1_LOC_709/B 0.00fF
C38705 NAND2X1_LOC_647/B INVX1_LOC_19/A 0.00fF
C38706 INVX1_LOC_135/A NOR2X1_LOC_459/B 0.04fF
C38707 NOR2X1_LOC_361/B INVX1_LOC_59/Y 0.00fF
C38708 INVX1_LOC_103/A NOR2X1_LOC_56/Y -0.01fF
C38709 INVX1_LOC_271/A INVX1_LOC_307/A 0.10fF
C38710 INVX1_LOC_35/A NOR2X1_LOC_351/Y 0.39fF
C38711 INVX1_LOC_174/A NAND2X1_LOC_149/a_36_24# 0.00fF
C38712 NAND2X1_LOC_803/B NAND2X1_LOC_649/B 0.32fF
C38713 NOR2X1_LOC_272/Y INVX1_LOC_12/Y 0.26fF
C38714 NOR2X1_LOC_720/B D_INPUT_0 0.06fF
C38715 NOR2X1_LOC_82/A INVX1_LOC_316/A 0.02fF
C38716 INVX1_LOC_83/A NOR2X1_LOC_52/B 0.08fF
C38717 INVX1_LOC_206/A INVX1_LOC_10/A 0.05fF
C38718 INVX1_LOC_229/Y NAND2X1_LOC_839/Y 0.45fF
C38719 INVX1_LOC_40/A NOR2X1_LOC_121/A 0.03fF
C38720 NOR2X1_LOC_430/A INVX1_LOC_140/A 0.07fF
C38721 NOR2X1_LOC_778/B NOR2X1_LOC_730/A 0.01fF
C38722 INVX1_LOC_53/A NOR2X1_LOC_858/a_36_216# 0.00fF
C38723 NOR2X1_LOC_205/Y INVX1_LOC_139/A 0.00fF
C38724 INVX1_LOC_77/A INVX1_LOC_73/A 0.07fF
C38725 NOR2X1_LOC_561/Y INVX1_LOC_144/Y -0.03fF
C38726 INVX1_LOC_226/Y INVX1_LOC_137/A 0.01fF
C38727 NOR2X1_LOC_536/A NOR2X1_LOC_384/A 0.16fF
C38728 NOR2X1_LOC_846/Y INVX1_LOC_9/A 0.01fF
C38729 NOR2X1_LOC_657/Y INVX1_LOC_159/Y 0.04fF
C38730 INVX1_LOC_89/A NOR2X1_LOC_423/Y 0.06fF
C38731 INVX1_LOC_103/A VDD 4.44fF
C38732 NOR2X1_LOC_738/A NOR2X1_LOC_732/A 0.01fF
C38733 INVX1_LOC_36/A NOR2X1_LOC_269/Y 0.09fF
C38734 NOR2X1_LOC_312/Y NOR2X1_LOC_312/a_36_216# 0.00fF
C38735 INVX1_LOC_268/A INVX1_LOC_290/A 0.02fF
C38736 NAND2X1_LOC_714/B INVX1_LOC_38/A 0.03fF
C38737 INVX1_LOC_11/A INVX1_LOC_46/A 0.03fF
C38738 INVX1_LOC_186/Y NOR2X1_LOC_302/A 0.04fF
C38739 INVX1_LOC_103/A NAND2X1_LOC_800/A 0.00fF
C38740 INVX1_LOC_5/A NOR2X1_LOC_640/Y 0.42fF
C38741 NOR2X1_LOC_254/A INVX1_LOC_76/A 0.61fF
C38742 INVX1_LOC_135/A NAND2X1_LOC_850/Y 0.10fF
C38743 INVX1_LOC_279/A INVX1_LOC_16/A 0.07fF
C38744 INVX1_LOC_119/A NOR2X1_LOC_329/B 0.46fF
C38745 INVX1_LOC_181/Y INVX1_LOC_98/A 0.02fF
C38746 NOR2X1_LOC_222/Y INVX1_LOC_89/A 0.03fF
C38747 NOR2X1_LOC_355/A INVX1_LOC_208/A 0.18fF
C38748 INVX1_LOC_292/A VDD 0.30fF
C38749 NAND2X1_LOC_561/B INVX1_LOC_38/A 0.15fF
C38750 INVX1_LOC_181/Y NOR2X1_LOC_78/A 0.03fF
C38751 NOR2X1_LOC_419/Y INVX1_LOC_123/A 0.01fF
C38752 NAND2X1_LOC_361/Y NOR2X1_LOC_9/Y 0.02fF
C38753 NAND2X1_LOC_452/Y D_INPUT_5 0.16fF
C38754 NAND2X1_LOC_579/A INVX1_LOC_118/A 0.10fF
C38755 NOR2X1_LOC_315/Y INVX1_LOC_75/A 0.07fF
C38756 INVX1_LOC_124/A INVX1_LOC_73/A 0.94fF
C38757 NOR2X1_LOC_208/Y NOR2X1_LOC_269/Y 0.02fF
C38758 NAND2X1_LOC_303/Y INVX1_LOC_54/A 0.03fF
C38759 NOR2X1_LOC_295/Y NOR2X1_LOC_113/B 0.04fF
C38760 NOR2X1_LOC_663/A NOR2X1_LOC_649/B 0.02fF
C38761 NAND2X1_LOC_474/Y NOR2X1_LOC_216/B 0.10fF
C38762 INVX1_LOC_50/Y NAND2X1_LOC_574/A 0.03fF
C38763 INVX1_LOC_271/A INVX1_LOC_12/A 0.25fF
C38764 INVX1_LOC_105/Y INVX1_LOC_12/A 0.11fF
C38765 NAND2X1_LOC_198/B NAND2X1_LOC_469/B 0.01fF
C38766 INVX1_LOC_89/A INVX1_LOC_220/Y 0.02fF
C38767 INVX1_LOC_174/A NOR2X1_LOC_378/Y 0.01fF
C38768 NOR2X1_LOC_738/A NOR2X1_LOC_687/Y 0.01fF
C38769 INVX1_LOC_178/A NOR2X1_LOC_697/Y 0.05fF
C38770 NOR2X1_LOC_724/Y NOR2X1_LOC_730/A 0.01fF
C38771 INVX1_LOC_87/A INVX1_LOC_4/Y 0.02fF
C38772 INVX1_LOC_58/A INVX1_LOC_102/A 0.26fF
C38773 NOR2X1_LOC_717/A INVX1_LOC_263/Y 0.07fF
C38774 NAND2X1_LOC_9/Y NOR2X1_LOC_89/A 0.00fF
C38775 NOR2X1_LOC_160/B INVX1_LOC_127/A 0.01fF
C38776 NOR2X1_LOC_520/B NAND2X1_LOC_642/Y 0.00fF
C38777 INVX1_LOC_182/Y INVX1_LOC_16/A 0.03fF
C38778 INVX1_LOC_95/Y NOR2X1_LOC_6/a_36_216# 0.01fF
C38779 NAND2X1_LOC_364/A INVX1_LOC_12/Y 0.01fF
C38780 INVX1_LOC_314/Y NOR2X1_LOC_9/a_36_216# 0.00fF
C38781 NOR2X1_LOC_337/a_36_216# INVX1_LOC_91/A 0.01fF
C38782 INVX1_LOC_233/A NOR2X1_LOC_89/A 0.15fF
C38783 NOR2X1_LOC_717/A INVX1_LOC_42/A 0.03fF
C38784 INVX1_LOC_279/A INVX1_LOC_28/A 0.07fF
C38785 INVX1_LOC_9/Y INVX1_LOC_79/A 0.02fF
C38786 NOR2X1_LOC_420/a_36_216# NAND2X1_LOC_63/Y 0.00fF
C38787 INVX1_LOC_72/A NOR2X1_LOC_536/A 0.21fF
C38788 NOR2X1_LOC_52/B NOR2X1_LOC_311/Y 0.00fF
C38789 NOR2X1_LOC_82/Y INPUT_0 0.03fF
C38790 NAND2X1_LOC_214/B INVX1_LOC_12/A 0.02fF
C38791 NOR2X1_LOC_433/A INVX1_LOC_46/A 0.32fF
C38792 INVX1_LOC_31/A NOR2X1_LOC_660/a_36_216# 0.01fF
C38793 NAND2X1_LOC_339/a_36_24# INVX1_LOC_147/Y 0.00fF
C38794 INVX1_LOC_31/A NOR2X1_LOC_235/Y 0.02fF
C38795 NAND2X1_LOC_794/B NOR2X1_LOC_189/a_36_216# 0.01fF
C38796 NOR2X1_LOC_593/Y INVX1_LOC_46/A 0.14fF
C38797 NAND2X1_LOC_724/Y NOR2X1_LOC_409/B 0.03fF
C38798 NOR2X1_LOC_798/A NOR2X1_LOC_89/A 0.46fF
C38799 NOR2X1_LOC_544/A INVX1_LOC_186/A 0.07fF
C38800 INVX1_LOC_27/A INVX1_LOC_12/A 0.29fF
C38801 D_INPUT_1 NOR2X1_LOC_394/Y 0.02fF
C38802 NOR2X1_LOC_816/A NOR2X1_LOC_697/Y 0.00fF
C38803 NOR2X1_LOC_824/A INVX1_LOC_12/A 0.07fF
C38804 INVX1_LOC_75/A INVX1_LOC_66/A 0.02fF
C38805 INVX1_LOC_227/A INPUT_0 0.72fF
C38806 NOR2X1_LOC_759/Y INVX1_LOC_38/A 0.00fF
C38807 INVX1_LOC_63/Y INVX1_LOC_37/A 0.01fF
C38808 INVX1_LOC_89/A D_INPUT_4 0.01fF
C38809 INVX1_LOC_224/A NOR2X1_LOC_68/Y 0.01fF
C38810 NOR2X1_LOC_418/Y NOR2X1_LOC_45/B 0.02fF
C38811 INVX1_LOC_72/A NAND2X1_LOC_93/B 0.10fF
C38812 INVX1_LOC_11/A NOR2X1_LOC_68/Y 0.03fF
C38813 NOR2X1_LOC_78/B INVX1_LOC_199/A 0.03fF
C38814 NAND2X1_LOC_538/Y INVX1_LOC_264/A 0.02fF
C38815 INVX1_LOC_240/A VDD 2.14fF
C38816 NAND2X1_LOC_703/Y NAND2X1_LOC_668/a_36_24# 0.00fF
C38817 NOR2X1_LOC_52/B INVX1_LOC_46/A 0.13fF
C38818 NAND2X1_LOC_593/Y NOR2X1_LOC_331/B 0.02fF
C38819 NOR2X1_LOC_68/A NOR2X1_LOC_78/Y 0.03fF
C38820 INVX1_LOC_251/Y INVX1_LOC_20/A 0.12fF
C38821 INVX1_LOC_240/A NAND2X1_LOC_800/A 0.33fF
C38822 INVX1_LOC_182/Y INVX1_LOC_28/A 0.03fF
C38823 NOR2X1_LOC_644/B INVX1_LOC_84/A 0.03fF
C38824 NOR2X1_LOC_589/A NOR2X1_LOC_45/B 0.18fF
C38825 NOR2X1_LOC_471/Y INVX1_LOC_186/Y 0.02fF
C38826 NOR2X1_LOC_636/B NAND2X1_LOC_639/a_36_24# 0.01fF
C38827 NAND2X1_LOC_231/Y NAND2X1_LOC_650/B 0.13fF
C38828 NOR2X1_LOC_175/A INVX1_LOC_37/A 0.07fF
C38829 NOR2X1_LOC_554/B NOR2X1_LOC_820/a_36_216# 0.01fF
C38830 NOR2X1_LOC_343/B INVX1_LOC_15/A 0.02fF
C38831 NOR2X1_LOC_357/Y NOR2X1_LOC_352/Y 0.10fF
C38832 INVX1_LOC_136/A NOR2X1_LOC_841/A 0.39fF
C38833 NAND2X1_LOC_363/B NAND2X1_LOC_91/a_36_24# 0.00fF
C38834 NOR2X1_LOC_374/A NOR2X1_LOC_729/A 0.03fF
C38835 NOR2X1_LOC_547/a_36_216# INVX1_LOC_176/A 0.00fF
C38836 NOR2X1_LOC_219/Y NAND2X1_LOC_469/B 0.01fF
C38837 NOR2X1_LOC_655/B INVX1_LOC_14/Y 0.01fF
C38838 INVX1_LOC_314/Y INVX1_LOC_92/A 0.04fF
C38839 NOR2X1_LOC_65/B NOR2X1_LOC_717/A 0.01fF
C38840 INVX1_LOC_290/A INVX1_LOC_187/Y 0.01fF
C38841 INPUT_0 NOR2X1_LOC_703/A 0.03fF
C38842 NOR2X1_LOC_139/Y NOR2X1_LOC_366/Y 0.03fF
C38843 NOR2X1_LOC_589/A INVX1_LOC_199/Y 0.01fF
C38844 NOR2X1_LOC_690/A INVX1_LOC_54/A 0.10fF
C38845 NOR2X1_LOC_78/A INVX1_LOC_148/Y 0.03fF
C38846 NOR2X1_LOC_372/Y NAND2X1_LOC_489/Y 0.01fF
C38847 INVX1_LOC_230/Y NOR2X1_LOC_664/a_36_216# 0.00fF
C38848 NAND2X1_LOC_466/Y INVX1_LOC_54/A 0.01fF
C38849 NOR2X1_LOC_288/A NOR2X1_LOC_729/A 0.08fF
C38850 NOR2X1_LOC_442/a_36_216# INVX1_LOC_15/A 0.01fF
C38851 INVX1_LOC_35/A NOR2X1_LOC_748/A 0.05fF
C38852 NOR2X1_LOC_537/Y NOR2X1_LOC_536/A 0.03fF
C38853 INVX1_LOC_18/A NOR2X1_LOC_257/Y 0.03fF
C38854 NOR2X1_LOC_151/Y NOR2X1_LOC_728/a_36_216# 0.00fF
C38855 NOR2X1_LOC_194/Y INVX1_LOC_54/A 0.01fF
C38856 NAND2X1_LOC_338/B NOR2X1_LOC_536/A 0.24fF
C38857 INVX1_LOC_13/Y INVX1_LOC_23/Y 0.03fF
C38858 NOR2X1_LOC_296/a_36_216# INVX1_LOC_3/Y 0.00fF
C38859 NOR2X1_LOC_366/Y NAND2X1_LOC_468/B 0.02fF
C38860 NOR2X1_LOC_360/Y INVX1_LOC_63/A 0.08fF
C38861 NOR2X1_LOC_322/Y NOR2X1_LOC_167/Y 0.05fF
C38862 INVX1_LOC_279/A NOR2X1_LOC_35/Y 0.10fF
C38863 INVX1_LOC_303/A NAND2X1_LOC_52/a_36_24# 0.07fF
C38864 NOR2X1_LOC_382/Y INVX1_LOC_29/A 1.16fF
C38865 NOR2X1_LOC_557/Y NOR2X1_LOC_831/B 0.08fF
C38866 NOR2X1_LOC_754/Y NAND2X1_LOC_793/B 0.06fF
C38867 NAND2X1_LOC_812/A INVX1_LOC_297/A 0.02fF
C38868 NAND2X1_LOC_464/B NOR2X1_LOC_291/Y 0.53fF
C38869 NOR2X1_LOC_309/Y NOR2X1_LOC_79/Y 0.01fF
C38870 NAND2X1_LOC_662/Y INVX1_LOC_117/A 0.14fF
C38871 NOR2X1_LOC_355/A NAND2X1_LOC_211/Y 0.18fF
C38872 NOR2X1_LOC_584/a_36_216# NOR2X1_LOC_584/Y 0.00fF
C38873 NOR2X1_LOC_82/A INVX1_LOC_4/Y 0.08fF
C38874 NOR2X1_LOC_644/B INVX1_LOC_15/A 0.01fF
C38875 INVX1_LOC_192/Y NAND2X1_LOC_93/B 0.02fF
C38876 NAND2X1_LOC_521/a_36_24# INVX1_LOC_29/A 0.01fF
C38877 INVX1_LOC_120/A VDD 0.00fF
C38878 NOR2X1_LOC_62/a_36_216# INVX1_LOC_9/A 0.00fF
C38879 NOR2X1_LOC_6/B NAND2X1_LOC_574/A 2.81fF
C38880 INVX1_LOC_192/Y NAND2X1_LOC_425/Y 0.09fF
C38881 NOR2X1_LOC_666/A INVX1_LOC_270/A 0.02fF
C38882 INVX1_LOC_121/A NOR2X1_LOC_684/Y 0.01fF
C38883 INVX1_LOC_249/A INVX1_LOC_12/A 0.13fF
C38884 INVX1_LOC_17/A NOR2X1_LOC_843/B 0.09fF
C38885 INVX1_LOC_108/Y NAND2X1_LOC_816/a_36_24# 0.00fF
C38886 INVX1_LOC_67/A INVX1_LOC_133/A -0.02fF
C38887 NOR2X1_LOC_792/B INVX1_LOC_63/A 0.02fF
C38888 INVX1_LOC_83/A NOR2X1_LOC_376/Y 0.02fF
C38889 INVX1_LOC_14/A NAND2X1_LOC_205/A 0.01fF
C38890 NOR2X1_LOC_172/Y NAND2X1_LOC_74/B 0.03fF
C38891 NOR2X1_LOC_19/B INVX1_LOC_178/Y 0.04fF
C38892 NOR2X1_LOC_359/a_36_216# INVX1_LOC_23/A 0.02fF
C38893 INVX1_LOC_226/Y NOR2X1_LOC_216/B 0.03fF
C38894 NAND2X1_LOC_338/B INVX1_LOC_3/A 1.41fF
C38895 INVX1_LOC_91/Y INVX1_LOC_20/A 0.00fF
C38896 NOR2X1_LOC_392/B NAND2X1_LOC_74/B 0.01fF
C38897 INVX1_LOC_72/A NAND2X1_LOC_470/B 0.02fF
C38898 INVX1_LOC_311/A NOR2X1_LOC_603/Y 0.03fF
C38899 NAND2X1_LOC_374/Y NAND2X1_LOC_489/Y 0.00fF
C38900 INPUT_0 NAND2X1_LOC_650/B 0.03fF
C38901 NOR2X1_LOC_180/B INVX1_LOC_9/A 0.08fF
C38902 INVX1_LOC_36/A INVX1_LOC_26/A 0.25fF
C38903 NAND2X1_LOC_9/Y INVX1_LOC_11/A 0.09fF
C38904 INVX1_LOC_104/A INVX1_LOC_99/A 0.07fF
C38905 NAND2X1_LOC_342/Y INVX1_LOC_19/A 0.02fF
C38906 INVX1_LOC_22/A NOR2X1_LOC_430/Y 0.00fF
C38907 INVX1_LOC_10/A NOR2X1_LOC_216/B 0.03fF
C38908 INVX1_LOC_233/A INVX1_LOC_11/A 0.07fF
C38909 NOR2X1_LOC_34/A INVX1_LOC_27/A 0.01fF
C38910 INVX1_LOC_230/Y INVX1_LOC_23/A 1.41fF
C38911 INVX1_LOC_57/Y NOR2X1_LOC_693/Y 0.49fF
C38912 NOR2X1_LOC_267/A INVX1_LOC_26/A 0.18fF
C38913 NOR2X1_LOC_403/B NOR2X1_LOC_394/Y 0.14fF
C38914 NOR2X1_LOC_45/B INVX1_LOC_147/Y 0.01fF
C38915 NAND2X1_LOC_276/Y INVX1_LOC_32/A 0.07fF
C38916 NOR2X1_LOC_13/Y INVX1_LOC_78/A 0.08fF
C38917 NOR2X1_LOC_152/Y INVX1_LOC_128/Y 0.01fF
C38918 INVX1_LOC_18/A NOR2X1_LOC_302/A 0.01fF
C38919 NOR2X1_LOC_378/a_36_216# NOR2X1_LOC_89/A 0.00fF
C38920 INVX1_LOC_45/A INVX1_LOC_270/Y 0.13fF
C38921 INVX1_LOC_313/Y NAND2X1_LOC_93/B 0.01fF
C38922 NOR2X1_LOC_45/B INVX1_LOC_20/A 0.18fF
C38923 INVX1_LOC_73/A INVX1_LOC_9/A 0.07fF
C38924 NOR2X1_LOC_562/B INVX1_LOC_76/A 0.10fF
C38925 NOR2X1_LOC_391/A INVX1_LOC_84/A 0.16fF
C38926 INVX1_LOC_59/A INVX1_LOC_48/Y 0.00fF
C38927 NOR2X1_LOC_430/A INVX1_LOC_78/A 0.00fF
C38928 NAND2X1_LOC_553/A INVX1_LOC_11/A 0.04fF
C38929 NOR2X1_LOC_554/B NOR2X1_LOC_105/a_36_216# 0.00fF
C38930 NOR2X1_LOC_577/Y INVX1_LOC_94/Y 0.00fF
C38931 INVX1_LOC_58/A INVX1_LOC_223/A 0.01fF
C38932 NOR2X1_LOC_510/Y INVX1_LOC_103/A 0.03fF
C38933 NOR2X1_LOC_643/A INVX1_LOC_27/A 0.01fF
C38934 INVX1_LOC_11/A NOR2X1_LOC_798/A 0.03fF
C38935 NAND2X1_LOC_577/A NOR2X1_LOC_392/Y 0.07fF
C38936 INVX1_LOC_258/Y INVX1_LOC_258/A 0.09fF
C38937 NOR2X1_LOC_15/Y NOR2X1_LOC_92/Y 0.31fF
C38938 INVX1_LOC_277/A NOR2X1_LOC_678/A 0.05fF
C38939 NAND2X1_LOC_354/Y NAND2X1_LOC_678/a_36_24# 0.00fF
C38940 NOR2X1_LOC_558/A NAND2X1_LOC_642/Y 0.00fF
C38941 INVX1_LOC_284/Y NAND2X1_LOC_725/A 0.01fF
C38942 NOR2X1_LOC_65/B NOR2X1_LOC_13/Y 0.38fF
C38943 INVX1_LOC_233/Y NAND2X1_LOC_500/Y 0.04fF
C38944 INVX1_LOC_45/Y NOR2X1_LOC_383/B 2.25fF
C38945 NOR2X1_LOC_824/Y NAND2X1_LOC_836/Y 0.14fF
C38946 NOR2X1_LOC_689/Y NAND2X1_LOC_731/Y 0.16fF
C38947 INVX1_LOC_2/Y NOR2X1_LOC_346/Y 0.08fF
C38948 NOR2X1_LOC_437/a_36_216# INVX1_LOC_270/A 0.12fF
C38949 NAND2X1_LOC_854/B INVX1_LOC_49/Y 0.01fF
C38950 INVX1_LOC_254/Y NOR2X1_LOC_621/A 0.00fF
C38951 NOR2X1_LOC_542/B VDD 0.07fF
C38952 NOR2X1_LOC_113/A INVX1_LOC_12/Y 0.01fF
C38953 INVX1_LOC_11/A NAND2X1_LOC_703/Y 0.06fF
C38954 INVX1_LOC_61/Y INVX1_LOC_306/Y 0.35fF
C38955 NOR2X1_LOC_405/A INVX1_LOC_12/Y 0.10fF
C38956 NOR2X1_LOC_272/Y NOR2X1_LOC_160/B 0.01fF
C38957 INVX1_LOC_251/Y INVX1_LOC_4/A 0.07fF
C38958 INVX1_LOC_71/A INVX1_LOC_270/Y 0.46fF
C38959 NAND2X1_LOC_836/Y INVX1_LOC_76/A 0.01fF
C38960 NOR2X1_LOC_424/Y NAND2X1_LOC_449/a_36_24# 0.00fF
C38961 INVX1_LOC_11/Y NAND2X1_LOC_804/Y 0.08fF
C38962 INVX1_LOC_279/A INVX1_LOC_109/A 0.45fF
C38963 INVX1_LOC_89/A NOR2X1_LOC_691/B 0.01fF
C38964 VDD INVX1_LOC_143/Y 0.13fF
C38965 INVX1_LOC_140/A NOR2X1_LOC_697/Y 0.03fF
C38966 NOR2X1_LOC_817/Y INVX1_LOC_14/A 0.42fF
C38967 NOR2X1_LOC_790/B INVX1_LOC_24/A 0.03fF
C38968 INVX1_LOC_234/A INVX1_LOC_12/A 1.27fF
C38969 NAND2X1_LOC_564/A NOR2X1_LOC_237/Y 0.11fF
C38970 NOR2X1_LOC_234/a_36_216# INVX1_LOC_23/Y 0.00fF
C38971 NAND2X1_LOC_149/Y NOR2X1_LOC_389/A 0.10fF
C38972 NAND2X1_LOC_656/A NOR2X1_LOC_392/Y 0.10fF
C38973 NAND2X1_LOC_451/Y NAND2X1_LOC_452/Y 0.06fF
C38974 VDD NOR2X1_LOC_137/Y 0.15fF
C38975 NOR2X1_LOC_94/a_36_216# INVX1_LOC_3/Y 0.01fF
C38976 D_INPUT_1 NOR2X1_LOC_716/B 0.07fF
C38977 NAND2X1_LOC_725/A NAND2X1_LOC_731/Y 0.02fF
C38978 NOR2X1_LOC_658/Y NOR2X1_LOC_215/A 0.03fF
C38979 INVX1_LOC_268/A NOR2X1_LOC_467/A 0.32fF
C38980 NOR2X1_LOC_554/B NOR2X1_LOC_649/Y 0.24fF
C38981 NOR2X1_LOC_111/A NAND2X1_LOC_211/Y 0.43fF
C38982 NOR2X1_LOC_567/B INVX1_LOC_63/A 0.03fF
C38983 INVX1_LOC_90/A NAND2X1_LOC_74/B 1.09fF
C38984 INVX1_LOC_16/A NOR2X1_LOC_38/B 0.06fF
C38985 NAND2X1_LOC_41/Y INVX1_LOC_15/A 0.04fF
C38986 INVX1_LOC_21/A NOR2X1_LOC_703/B 0.03fF
C38987 NOR2X1_LOC_214/B INVX1_LOC_109/Y 0.02fF
C38988 NOR2X1_LOC_557/A INVX1_LOC_92/A 0.09fF
C38989 NOR2X1_LOC_824/A INVX1_LOC_217/A 0.10fF
C38990 NOR2X1_LOC_186/Y INVX1_LOC_181/Y 0.00fF
C38991 INVX1_LOC_36/A NOR2X1_LOC_666/A 0.04fF
C38992 INVX1_LOC_22/A INVX1_LOC_94/Y 0.42fF
C38993 NAND2X1_LOC_699/a_36_24# INVX1_LOC_46/A 0.00fF
C38994 NOR2X1_LOC_709/A NOR2X1_LOC_646/B 0.01fF
C38995 INVX1_LOC_58/A INVX1_LOC_85/A 0.01fF
C38996 NOR2X1_LOC_802/A INVX1_LOC_57/A 0.07fF
C38997 INVX1_LOC_41/A NOR2X1_LOC_434/A 0.02fF
C38998 INVX1_LOC_89/A NOR2X1_LOC_477/B 0.02fF
C38999 INVX1_LOC_286/Y NOR2X1_LOC_533/Y 0.06fF
C39000 NOR2X1_LOC_789/B INVX1_LOC_24/A 0.02fF
C39001 INVX1_LOC_299/A NOR2X1_LOC_274/B 1.31fF
C39002 NOR2X1_LOC_590/A INVX1_LOC_225/Y 0.03fF
C39003 NOR2X1_LOC_307/B NOR2X1_LOC_727/B 0.02fF
C39004 INVX1_LOC_221/A NAND2X1_LOC_590/a_36_24# 0.00fF
C39005 NAND2X1_LOC_9/Y NOR2X1_LOC_52/B 0.01fF
C39006 INVX1_LOC_88/Y NOR2X1_LOC_665/a_36_216# 0.00fF
C39007 NAND2X1_LOC_149/Y NOR2X1_LOC_596/A 0.14fF
C39008 NAND2X1_LOC_348/A NAND2X1_LOC_74/B 0.01fF
C39009 NAND2X1_LOC_785/a_36_24# NAND2X1_LOC_833/Y 0.00fF
C39010 INVX1_LOC_25/Y NAND2X1_LOC_99/A 0.19fF
C39011 INVX1_LOC_233/A NOR2X1_LOC_52/B 0.14fF
C39012 NOR2X1_LOC_68/A NAND2X1_LOC_537/Y 0.03fF
C39013 INVX1_LOC_230/Y INVX1_LOC_31/A 0.46fF
C39014 INVX1_LOC_306/A INVX1_LOC_4/Y 0.01fF
C39015 INVX1_LOC_17/A INVX1_LOC_18/A 1.63fF
C39016 INVX1_LOC_266/A INVX1_LOC_94/A 0.10fF
C39017 NOR2X1_LOC_798/A NOR2X1_LOC_593/Y 0.00fF
C39018 INPUT_0 NOR2X1_LOC_77/a_36_216# 0.00fF
C39019 INVX1_LOC_256/A INVX1_LOC_72/A 0.22fF
C39020 NOR2X1_LOC_208/Y NOR2X1_LOC_666/A 0.09fF
C39021 NOR2X1_LOC_824/A NAND2X1_LOC_787/B 0.10fF
C39022 NOR2X1_LOC_15/Y NAND2X1_LOC_837/Y 0.45fF
C39023 INVX1_LOC_74/Y NAND2X1_LOC_141/Y 0.03fF
C39024 D_INPUT_1 NOR2X1_LOC_757/Y 0.01fF
C39025 INVX1_LOC_22/A INVX1_LOC_296/A 0.09fF
C39026 NOR2X1_LOC_778/B INVX1_LOC_53/A 0.16fF
C39027 NOR2X1_LOC_667/Y INVX1_LOC_45/A 0.01fF
C39028 INVX1_LOC_36/A INVX1_LOC_141/A 0.01fF
C39029 INVX1_LOC_187/A INVX1_LOC_84/A 0.00fF
C39030 NOR2X1_LOC_471/Y INVX1_LOC_18/A 0.09fF
C39031 NAND2X1_LOC_341/A INVX1_LOC_23/A 0.03fF
C39032 NOR2X1_LOC_160/B NAND2X1_LOC_364/A 2.08fF
C39033 INVX1_LOC_28/A NOR2X1_LOC_38/B 0.16fF
C39034 INVX1_LOC_17/A NOR2X1_LOC_637/Y 0.02fF
C39035 INVX1_LOC_58/A NAND2X1_LOC_662/Y 0.01fF
C39036 NOR2X1_LOC_439/a_36_216# INVX1_LOC_53/A 0.00fF
C39037 NOR2X1_LOC_78/A NOR2X1_LOC_509/A 0.01fF
C39038 NAND2X1_LOC_53/Y NOR2X1_LOC_303/Y 0.00fF
C39039 INVX1_LOC_41/A NOR2X1_LOC_15/Y 0.03fF
C39040 NAND2X1_LOC_268/a_36_24# NOR2X1_LOC_271/Y 0.00fF
C39041 NOR2X1_LOC_598/B NOR2X1_LOC_210/A 0.02fF
C39042 NOR2X1_LOC_445/Y INVX1_LOC_269/A 0.03fF
C39043 INVX1_LOC_47/A INVX1_LOC_116/Y 0.00fF
C39044 NAND2X1_LOC_567/Y INVX1_LOC_161/Y 0.00fF
C39045 NOR2X1_LOC_328/Y NAND2X1_LOC_708/Y 0.63fF
C39046 NOR2X1_LOC_246/A NAND2X1_LOC_285/a_36_24# 0.01fF
C39047 INVX1_LOC_108/Y NAND2X1_LOC_41/Y 0.10fF
C39048 INVX1_LOC_54/Y NAND2X1_LOC_474/Y 0.01fF
C39049 INVX1_LOC_21/A NAND2X1_LOC_578/B 0.91fF
C39050 INVX1_LOC_36/A NOR2X1_LOC_820/A 0.10fF
C39051 INVX1_LOC_58/A NAND2X1_LOC_715/a_36_24# 0.01fF
C39052 NOR2X1_LOC_772/B INVX1_LOC_232/A 0.10fF
C39053 INVX1_LOC_36/A NOR2X1_LOC_276/B 0.01fF
C39054 D_INPUT_1 NOR2X1_LOC_717/B 0.00fF
C39055 INVX1_LOC_254/A INVX1_LOC_218/Y 0.30fF
C39056 NOR2X1_LOC_15/Y NAND2X1_LOC_477/A 0.03fF
C39057 NOR2X1_LOC_441/Y NOR2X1_LOC_106/Y 0.02fF
C39058 VDD NOR2X1_LOC_631/A 0.11fF
C39059 INVX1_LOC_15/Y NOR2X1_LOC_92/Y 0.02fF
C39060 INVX1_LOC_135/A NOR2X1_LOC_629/A 0.01fF
C39061 INVX1_LOC_177/Y INVX1_LOC_79/Y 0.24fF
C39062 NOR2X1_LOC_644/A NOR2X1_LOC_383/B 0.05fF
C39063 INVX1_LOC_235/Y NOR2X1_LOC_399/Y 0.03fF
C39064 INVX1_LOC_13/Y INVX1_LOC_232/A 0.03fF
C39065 INVX1_LOC_50/A NOR2X1_LOC_356/A 0.07fF
C39066 NOR2X1_LOC_781/Y INVX1_LOC_72/A 0.07fF
C39067 NOR2X1_LOC_562/A INVX1_LOC_19/A 0.06fF
C39068 INPUT_3 NAND2X1_LOC_276/Y 0.09fF
C39069 INVX1_LOC_289/A INVX1_LOC_178/A 0.06fF
C39070 INVX1_LOC_1/A INVX1_LOC_196/A 0.10fF
C39071 NOR2X1_LOC_685/A NOR2X1_LOC_685/Y 0.02fF
C39072 NAND2X1_LOC_350/A NAND2X1_LOC_466/Y 0.03fF
C39073 INVX1_LOC_35/A INVX1_LOC_150/A 0.06fF
C39074 NOR2X1_LOC_92/a_36_216# NAND2X1_LOC_74/B 0.00fF
C39075 NOR2X1_LOC_561/Y NOR2X1_LOC_304/a_36_216# 0.01fF
C39076 NOR2X1_LOC_314/a_36_216# INVX1_LOC_12/A 0.00fF
C39077 NAND2X1_LOC_538/Y INVX1_LOC_236/A 0.02fF
C39078 INVX1_LOC_35/A NOR2X1_LOC_110/a_36_216# 0.00fF
C39079 INVX1_LOC_6/A NAND2X1_LOC_471/Y 0.04fF
C39080 NOR2X1_LOC_828/B NOR2X1_LOC_383/B 0.04fF
C39081 D_INPUT_0 INVX1_LOC_292/Y 0.01fF
C39082 INVX1_LOC_75/A NAND2X1_LOC_99/A 0.07fF
C39083 NAND2X1_LOC_624/B INVX1_LOC_135/A 0.07fF
C39084 INVX1_LOC_259/Y INVX1_LOC_90/A 0.01fF
C39085 NAND2X1_LOC_492/a_36_24# NOR2X1_LOC_717/A 0.00fF
C39086 NOR2X1_LOC_724/Y INVX1_LOC_53/A 0.03fF
C39087 INVX1_LOC_35/A INVX1_LOC_89/A 3.10fF
C39088 NAND2X1_LOC_363/B INVX1_LOC_65/Y 0.00fF
C39089 NOR2X1_LOC_276/B NOR2X1_LOC_208/Y 0.03fF
C39090 INVX1_LOC_1/A NAND2X1_LOC_841/A 0.04fF
C39091 INVX1_LOC_90/A NOR2X1_LOC_660/Y 0.15fF
C39092 INVX1_LOC_136/A NOR2X1_LOC_172/Y 0.01fF
C39093 INVX1_LOC_13/A NOR2X1_LOC_611/a_36_216# 0.00fF
C39094 NOR2X1_LOC_382/Y INVX1_LOC_8/A 0.01fF
C39095 INVX1_LOC_292/A INVX1_LOC_177/A 0.01fF
C39096 NOR2X1_LOC_468/Y INVX1_LOC_16/A 3.02fF
C39097 INVX1_LOC_136/A NOR2X1_LOC_772/Y 0.10fF
C39098 NAND2X1_LOC_123/Y INVX1_LOC_53/A 0.07fF
C39099 NAND2X1_LOC_254/Y INVX1_LOC_46/A 0.01fF
C39100 INVX1_LOC_299/A INVX1_LOC_22/A 0.07fF
C39101 INVX1_LOC_36/A INVX1_LOC_315/A 0.36fF
C39102 INVX1_LOC_50/A NOR2X1_LOC_74/A 0.15fF
C39103 INVX1_LOC_13/A NOR2X1_LOC_140/A 0.18fF
C39104 NOR2X1_LOC_785/A INVX1_LOC_143/A 0.42fF
C39105 NAND2X1_LOC_72/Y NOR2X1_LOC_356/A 0.18fF
C39106 NAND2X1_LOC_717/Y NAND2X1_LOC_546/a_36_24# 0.00fF
C39107 INVX1_LOC_90/A NOR2X1_LOC_845/a_36_216# 0.01fF
C39108 INVX1_LOC_247/A INVX1_LOC_4/A 0.03fF
C39109 NOR2X1_LOC_13/Y NOR2X1_LOC_152/Y 0.10fF
C39110 INVX1_LOC_24/A NOR2X1_LOC_387/Y 0.01fF
C39111 NAND2X1_LOC_624/B NOR2X1_LOC_490/Y 0.02fF
C39112 INVX1_LOC_45/A NOR2X1_LOC_310/Y 0.01fF
C39113 NOR2X1_LOC_538/B INVX1_LOC_22/A 0.02fF
C39114 INVX1_LOC_136/A NOR2X1_LOC_392/B 0.10fF
C39115 GATE_741 NOR2X1_LOC_576/B 0.36fF
C39116 INVX1_LOC_50/A NOR2X1_LOC_9/Y 0.03fF
C39117 NOR2X1_LOC_68/A NOR2X1_LOC_486/B 0.08fF
C39118 NOR2X1_LOC_310/Y NOR2X1_LOC_568/A 0.04fF
C39119 NAND2X1_LOC_171/a_36_24# INVX1_LOC_179/Y 0.01fF
C39120 NOR2X1_LOC_273/Y INVX1_LOC_33/A 0.00fF
C39121 INVX1_LOC_38/A NAND2X1_LOC_74/B 3.68fF
C39122 NOR2X1_LOC_560/A NOR2X1_LOC_849/A 0.02fF
C39123 INVX1_LOC_269/A NOR2X1_LOC_32/Y 0.02fF
C39124 NOR2X1_LOC_71/Y NAND2X1_LOC_75/a_36_24# 0.01fF
C39125 NOR2X1_LOC_218/Y NOR2X1_LOC_218/A 0.31fF
C39126 INVX1_LOC_33/A NOR2X1_LOC_759/Y 0.02fF
C39127 INVX1_LOC_24/A NOR2X1_LOC_344/A 0.04fF
C39128 INVX1_LOC_34/A NOR2X1_LOC_215/Y 0.01fF
C39129 NOR2X1_LOC_598/B NOR2X1_LOC_97/A 0.54fF
C39130 INVX1_LOC_104/A INVX1_LOC_79/Y 0.01fF
C39131 NAND2X1_LOC_794/B NOR2X1_LOC_166/a_36_216# 0.04fF
C39132 NOR2X1_LOC_620/Y INVX1_LOC_77/A 0.03fF
C39133 INVX1_LOC_202/A INVX1_LOC_33/A 0.00fF
C39134 INVX1_LOC_225/A INVX1_LOC_181/Y 0.01fF
C39135 NAND2X1_LOC_500/Y NOR2X1_LOC_526/Y 0.07fF
C39136 NOR2X1_LOC_45/B NAND2X1_LOC_420/a_36_24# 0.00fF
C39137 NAND2X1_LOC_308/Y NAND2X1_LOC_731/Y 0.02fF
C39138 INVX1_LOC_88/A NOR2X1_LOC_366/Y 0.01fF
C39139 NAND2X1_LOC_72/Y NOR2X1_LOC_74/A 0.18fF
C39140 INVX1_LOC_122/A INVX1_LOC_15/A 0.02fF
C39141 NAND2X1_LOC_357/B INVX1_LOC_24/A 0.07fF
C39142 NAND2X1_LOC_802/A NAND2X1_LOC_354/B 0.03fF
C39143 NOR2X1_LOC_103/a_36_216# NAND2X1_LOC_489/Y 0.00fF
C39144 INVX1_LOC_313/Y NOR2X1_LOC_348/Y 0.01fF
C39145 NAND2X1_LOC_577/A INVX1_LOC_25/Y 0.00fF
C39146 INVX1_LOC_230/Y NAND2X1_LOC_859/Y 0.00fF
C39147 NAND2X1_LOC_733/Y NOR2X1_LOC_695/Y 0.07fF
C39148 INVX1_LOC_47/A INVX1_LOC_1/A 0.07fF
C39149 NAND2X1_LOC_364/Y NAND2X1_LOC_365/a_36_24# 0.01fF
C39150 NOR2X1_LOC_653/Y INVX1_LOC_285/A 0.02fF
C39151 INVX1_LOC_35/A NOR2X1_LOC_703/Y 0.68fF
C39152 INVX1_LOC_269/A NOR2X1_LOC_542/Y -0.00fF
C39153 NOR2X1_LOC_720/B INVX1_LOC_49/A 0.08fF
C39154 INVX1_LOC_281/A INVX1_LOC_4/A 0.01fF
C39155 INVX1_LOC_21/A INVX1_LOC_79/A 0.47fF
C39156 D_INPUT_0 NAND2X1_LOC_529/a_36_24# 0.00fF
C39157 NAND2X1_LOC_650/B INVX1_LOC_183/A 0.03fF
C39158 NOR2X1_LOC_216/B INVX1_LOC_12/A 0.10fF
C39159 NOR2X1_LOC_860/B INVX1_LOC_64/Y 0.02fF
C39160 NOR2X1_LOC_431/Y NOR2X1_LOC_226/A 0.02fF
C39161 INVX1_LOC_19/A INVX1_LOC_285/A 0.07fF
C39162 NOR2X1_LOC_516/B NAND2X1_LOC_364/A 0.10fF
C39163 INVX1_LOC_25/A INVX1_LOC_95/Y 0.02fF
C39164 INVX1_LOC_256/A INVX1_LOC_313/Y 0.01fF
C39165 NOR2X1_LOC_78/B INVX1_LOC_314/Y 0.03fF
C39166 INVX1_LOC_34/A INVX1_LOC_104/A 0.07fF
C39167 INVX1_LOC_11/A NAND2X1_LOC_842/B 0.03fF
C39168 INVX1_LOC_64/A NOR2X1_LOC_45/B 0.18fF
C39169 NOR2X1_LOC_447/Y NOR2X1_LOC_226/A 0.01fF
C39170 NOR2X1_LOC_456/Y NOR2X1_LOC_486/Y 0.07fF
C39171 INVX1_LOC_19/A NOR2X1_LOC_814/A 0.97fF
C39172 NOR2X1_LOC_360/Y INVX1_LOC_1/Y 0.04fF
C39173 INVX1_LOC_47/Y NOR2X1_LOC_612/Y 0.02fF
C39174 INVX1_LOC_228/Y NOR2X1_LOC_19/B 0.03fF
C39175 NOR2X1_LOC_440/Y INVX1_LOC_72/A 0.06fF
C39176 NOR2X1_LOC_500/A NOR2X1_LOC_500/Y 0.03fF
C39177 INVX1_LOC_201/Y NAND2X1_LOC_141/A 0.01fF
C39178 VDD NOR2X1_LOC_677/Y 0.43fF
C39179 NOR2X1_LOC_500/Y NOR2X1_LOC_303/Y 0.10fF
C39180 NOR2X1_LOC_596/A INVX1_LOC_16/A 0.07fF
C39181 NOR2X1_LOC_102/a_36_216# INVX1_LOC_26/A 0.03fF
C39182 INVX1_LOC_2/A NOR2X1_LOC_364/Y -0.02fF
C39183 NOR2X1_LOC_703/B NOR2X1_LOC_565/B 0.01fF
C39184 INVX1_LOC_217/A INVX1_LOC_234/A 0.01fF
C39185 NOR2X1_LOC_89/A INVX1_LOC_119/Y 0.02fF
C39186 INVX1_LOC_64/A INVX1_LOC_247/A 0.01fF
C39187 NAND2X1_LOC_35/Y NOR2X1_LOC_124/A 0.06fF
C39188 INVX1_LOC_269/A NOR2X1_LOC_335/B 0.03fF
C39189 NOR2X1_LOC_859/A INVX1_LOC_135/A 0.00fF
C39190 INVX1_LOC_303/A INVX1_LOC_232/A 0.10fF
C39191 NOR2X1_LOC_389/A INVX1_LOC_28/A 0.10fF
C39192 NOR2X1_LOC_778/A NOR2X1_LOC_717/B 0.01fF
C39193 NOR2X1_LOC_577/Y NOR2X1_LOC_321/a_36_216# 0.00fF
C39194 INVX1_LOC_21/A INVX1_LOC_91/A 0.26fF
C39195 NAND2X1_LOC_79/a_36_24# INVX1_LOC_232/A 0.01fF
C39196 NOR2X1_LOC_828/Y INVX1_LOC_37/A 0.23fF
C39197 NOR2X1_LOC_772/B NAND2X1_LOC_447/Y 0.09fF
C39198 NOR2X1_LOC_186/Y NAND2X1_LOC_107/a_36_24# 0.00fF
C39199 INVX1_LOC_30/A D_GATE_366 0.01fF
C39200 INVX1_LOC_161/Y INVX1_LOC_67/Y 0.02fF
C39201 NOR2X1_LOC_598/B NOR2X1_LOC_858/B 0.03fF
C39202 NOR2X1_LOC_42/a_36_216# NOR2X1_LOC_392/Y 0.00fF
C39203 INVX1_LOC_5/A NOR2X1_LOC_631/B 0.98fF
C39204 NOR2X1_LOC_186/Y NOR2X1_LOC_675/A 0.00fF
C39205 NOR2X1_LOC_53/Y INVX1_LOC_20/A 0.01fF
C39206 INVX1_LOC_103/A INVX1_LOC_285/Y 0.12fF
C39207 INVX1_LOC_280/Y INVX1_LOC_240/A 0.02fF
C39208 NOR2X1_LOC_219/Y INVX1_LOC_63/Y 0.04fF
C39209 NOR2X1_LOC_320/Y NOR2X1_LOC_250/A 0.02fF
C39210 NAND2X1_LOC_164/a_36_24# NOR2X1_LOC_802/A 0.00fF
C39211 INVX1_LOC_14/A INVX1_LOC_286/A 0.43fF
C39212 INVX1_LOC_136/A INVX1_LOC_90/A 1.89fF
C39213 INVX1_LOC_224/Y NOR2X1_LOC_536/A 0.03fF
C39214 INVX1_LOC_284/Y NAND2X1_LOC_560/A 0.03fF
C39215 INVX1_LOC_13/Y NAND2X1_LOC_447/Y 0.03fF
C39216 NOR2X1_LOC_453/Y INVX1_LOC_91/A 0.63fF
C39217 INVX1_LOC_135/A INVX1_LOC_41/Y 0.01fF
C39218 NAND2X1_LOC_391/Y INVX1_LOC_304/A 0.01fF
C39219 INVX1_LOC_136/A NOR2X1_LOC_389/B 0.10fF
C39220 NOR2X1_LOC_68/A INVX1_LOC_85/Y 0.03fF
C39221 NOR2X1_LOC_295/Y INVX1_LOC_16/A 0.10fF
C39222 NOR2X1_LOC_617/Y INVX1_LOC_135/A 0.02fF
C39223 NOR2X1_LOC_99/Y INVX1_LOC_23/Y 0.07fF
C39224 NOR2X1_LOC_289/Y INVX1_LOC_30/A 0.01fF
C39225 INVX1_LOC_63/Y NOR2X1_LOC_665/A 0.12fF
C39226 NAND2X1_LOC_552/A INVX1_LOC_37/A 0.05fF
C39227 NOR2X1_LOC_48/B INVX1_LOC_262/Y 0.03fF
C39228 INVX1_LOC_135/A NAND2X1_LOC_593/Y 0.04fF
C39229 NOR2X1_LOC_263/a_36_216# INVX1_LOC_25/Y 0.02fF
C39230 NAND2X1_LOC_787/A NOR2X1_LOC_692/a_36_216# 0.00fF
C39231 NOR2X1_LOC_629/A INVX1_LOC_280/A 0.01fF
C39232 INVX1_LOC_5/A INVX1_LOC_37/A 0.20fF
C39233 NOR2X1_LOC_89/A NOR2X1_LOC_755/Y 0.00fF
C39234 INVX1_LOC_292/A INVX1_LOC_285/Y 0.03fF
C39235 NOR2X1_LOC_711/A NAND2X1_LOC_305/a_36_24# 0.00fF
C39236 NOR2X1_LOC_731/A NOR2X1_LOC_687/Y 0.03fF
C39237 NOR2X1_LOC_778/B NOR2X1_LOC_78/B 0.05fF
C39238 NOR2X1_LOC_315/Y INVX1_LOC_22/A 0.06fF
C39239 INVX1_LOC_200/A NOR2X1_LOC_528/Y 0.12fF
C39240 D_INPUT_1 NOR2X1_LOC_709/B 0.05fF
C39241 INVX1_LOC_5/A NOR2X1_LOC_231/A 0.08fF
C39242 INVX1_LOC_64/A INVX1_LOC_281/A 0.17fF
C39243 INVX1_LOC_78/A NOR2X1_LOC_697/Y 0.05fF
C39244 NAND2X1_LOC_361/Y D_INPUT_0 0.07fF
C39245 NOR2X1_LOC_272/Y NAND2X1_LOC_211/Y 0.04fF
C39246 INVX1_LOC_14/A INVX1_LOC_95/A 0.10fF
C39247 NOR2X1_LOC_355/A INVX1_LOC_155/A 0.20fF
C39248 NOR2X1_LOC_744/a_36_216# NOR2X1_LOC_329/B 0.01fF
C39249 INVX1_LOC_1/A INVX1_LOC_95/Y 0.12fF
C39250 INVX1_LOC_136/A NAND2X1_LOC_348/A 0.00fF
C39251 INVX1_LOC_36/A NOR2X1_LOC_368/A 0.03fF
C39252 INVX1_LOC_32/A INVX1_LOC_125/A 0.19fF
C39253 NAND2X1_LOC_717/Y NAND2X1_LOC_863/B 0.03fF
C39254 NOR2X1_LOC_432/Y INVX1_LOC_22/A 0.01fF
C39255 INVX1_LOC_13/A NOR2X1_LOC_709/A 0.09fF
C39256 NAND2X1_LOC_624/B INVX1_LOC_280/A 0.03fF
C39257 INVX1_LOC_271/A INVX1_LOC_92/A 0.73fF
C39258 NOR2X1_LOC_500/A NAND2X1_LOC_323/a_36_24# 0.01fF
C39259 INVX1_LOC_234/Y VDD 0.33fF
C39260 NOR2X1_LOC_433/A NAND2X1_LOC_842/B 0.00fF
C39261 NOR2X1_LOC_303/Y NOR2X1_LOC_302/Y 0.04fF
C39262 NAND2X1_LOC_736/Y NOR2X1_LOC_380/A 6.69fF
C39263 INVX1_LOC_177/Y INPUT_0 0.46fF
C39264 NOR2X1_LOC_160/B NOR2X1_LOC_349/A 0.14fF
C39265 NOR2X1_LOC_639/B INVX1_LOC_118/A 0.02fF
C39266 NAND2X1_LOC_190/Y NOR2X1_LOC_35/Y 0.03fF
C39267 INVX1_LOC_227/A INVX1_LOC_266/Y 0.00fF
C39268 NAND2X1_LOC_656/A INVX1_LOC_75/A 0.02fF
C39269 NOR2X1_LOC_160/B NOR2X1_LOC_405/A 0.14fF
C39270 NAND2X1_LOC_357/B NOR2X1_LOC_130/A 0.07fF
C39271 INVX1_LOC_69/Y INVX1_LOC_72/A 0.14fF
C39272 INVX1_LOC_292/A INVX1_LOC_65/A 0.10fF
C39273 INVX1_LOC_26/A INVX1_LOC_63/A 0.13fF
C39274 NOR2X1_LOC_605/a_36_216# NOR2X1_LOC_773/Y 0.01fF
C39275 INVX1_LOC_26/Y NOR2X1_LOC_814/A 0.04fF
C39276 NOR2X1_LOC_454/Y INVX1_LOC_117/A 0.17fF
C39277 INVX1_LOC_89/A INVX1_LOC_257/Y 0.00fF
C39278 NOR2X1_LOC_790/B NOR2X1_LOC_197/B 0.01fF
C39279 NAND2X1_LOC_223/A NAND2X1_LOC_74/B 0.07fF
C39280 INVX1_LOC_292/A NOR2X1_LOC_137/B 0.93fF
C39281 NOR2X1_LOC_533/Y VDD 0.67fF
C39282 NAND2X1_LOC_223/A NAND2X1_LOC_207/Y 0.39fF
C39283 NOR2X1_LOC_295/Y INVX1_LOC_28/A 0.01fF
C39284 INVX1_LOC_224/Y INVX1_LOC_3/A 0.07fF
C39285 NOR2X1_LOC_746/Y INVX1_LOC_30/A 0.05fF
C39286 INVX1_LOC_314/Y NOR2X1_LOC_193/a_36_216# 0.02fF
C39287 INVX1_LOC_71/A INVX1_LOC_126/Y 0.10fF
C39288 NOR2X1_LOC_778/B INVX1_LOC_83/A 0.03fF
C39289 INVX1_LOC_64/A NOR2X1_LOC_862/B 0.02fF
C39290 NOR2X1_LOC_52/B NAND2X1_LOC_842/B 0.03fF
C39291 NOR2X1_LOC_533/Y NAND2X1_LOC_800/A 0.02fF
C39292 INVX1_LOC_217/A NOR2X1_LOC_528/Y 0.28fF
C39293 NOR2X1_LOC_278/Y INVX1_LOC_29/A 1.31fF
C39294 INVX1_LOC_99/Y INVX1_LOC_307/A 0.02fF
C39295 NOR2X1_LOC_788/B NOR2X1_LOC_168/B 0.00fF
C39296 INVX1_LOC_160/Y NOR2X1_LOC_835/A 0.00fF
C39297 NAND2X1_LOC_84/Y INVX1_LOC_286/A 0.08fF
C39298 NOR2X1_LOC_318/B NOR2X1_LOC_360/Y 0.10fF
C39299 NOR2X1_LOC_160/B NOR2X1_LOC_857/A 0.08fF
C39300 NOR2X1_LOC_816/A INVX1_LOC_37/A 0.07fF
C39301 NAND2X1_LOC_38/a_36_24# INVX1_LOC_3/A 0.00fF
C39302 INVX1_LOC_16/A NAND2X1_LOC_795/Y 0.26fF
C39303 NOR2X1_LOC_78/B NOR2X1_LOC_724/Y 0.01fF
C39304 INVX1_LOC_50/Y NOR2X1_LOC_155/A 0.02fF
C39305 NOR2X1_LOC_180/B INVX1_LOC_179/Y 0.00fF
C39306 INVX1_LOC_102/A NOR2X1_LOC_167/a_36_216# 0.01fF
C39307 NAND2X1_LOC_833/Y NOR2X1_LOC_167/Y 0.02fF
C39308 NOR2X1_LOC_741/a_36_216# INVX1_LOC_266/Y 0.01fF
C39309 NOR2X1_LOC_147/A INVX1_LOC_275/A 0.12fF
C39310 INVX1_LOC_93/Y NOR2X1_LOC_360/Y 0.08fF
C39311 INVX1_LOC_27/A INVX1_LOC_92/A 0.61fF
C39312 NOR2X1_LOC_103/Y NOR2X1_LOC_536/A 0.12fF
C39313 INVX1_LOC_181/Y NAND2X1_LOC_642/Y 0.01fF
C39314 INVX1_LOC_89/A NOR2X1_LOC_121/A 0.12fF
C39315 INVX1_LOC_33/A NOR2X1_LOC_334/A 0.01fF
C39316 NAND2X1_LOC_358/Y NAND2X1_LOC_358/a_36_24# 0.02fF
C39317 INVX1_LOC_104/A INPUT_0 0.14fF
C39318 INVX1_LOC_14/A INVX1_LOC_54/A 0.10fF
C39319 NAND2X1_LOC_660/a_36_24# NAND2X1_LOC_660/Y 0.02fF
C39320 NOR2X1_LOC_315/Y INVX1_LOC_100/A 0.74fF
C39321 INVX1_LOC_62/Y NOR2X1_LOC_35/Y 0.10fF
C39322 NOR2X1_LOC_222/Y INVX1_LOC_75/A 0.03fF
C39323 INVX1_LOC_289/A INVX1_LOC_140/A 0.05fF
C39324 NOR2X1_LOC_576/B NOR2X1_LOC_299/Y 1.24fF
C39325 INVX1_LOC_45/A NAND2X1_LOC_639/A 1.18fF
C39326 INVX1_LOC_58/A INVX1_LOC_290/Y 0.10fF
C39327 NOR2X1_LOC_392/Y NOR2X1_LOC_671/a_36_216# 0.01fF
C39328 NOR2X1_LOC_486/Y NOR2X1_LOC_550/B 0.12fF
C39329 INVX1_LOC_286/A NOR2X1_LOC_612/B 0.03fF
C39330 NOR2X1_LOC_93/Y INVX1_LOC_84/A 0.02fF
C39331 NOR2X1_LOC_569/Y NOR2X1_LOC_564/Y 0.08fF
C39332 NOR2X1_LOC_103/Y NAND2X1_LOC_93/B 0.01fF
C39333 NOR2X1_LOC_6/B NOR2X1_LOC_845/A 0.00fF
C39334 INVX1_LOC_45/A NOR2X1_LOC_536/A 1.80fF
C39335 NOR2X1_LOC_232/Y NOR2X1_LOC_88/Y 0.04fF
C39336 NAND2X1_LOC_9/Y NAND2X1_LOC_254/Y 0.35fF
C39337 INVX1_LOC_304/Y NOR2X1_LOC_528/Y 0.10fF
C39338 NAND2X1_LOC_337/B NOR2X1_LOC_743/Y 0.30fF
C39339 INVX1_LOC_83/A NOR2X1_LOC_724/Y 0.03fF
C39340 NAND2X1_LOC_856/A NOR2X1_LOC_536/A 0.00fF
C39341 NOR2X1_LOC_751/a_36_216# NOR2X1_LOC_814/A 0.00fF
C39342 INVX1_LOC_62/Y NOR2X1_LOC_133/a_36_216# 0.01fF
C39343 INVX1_LOC_314/Y INVX1_LOC_46/A 0.07fF
C39344 INVX1_LOC_225/A NAND2X1_LOC_107/a_36_24# 0.01fF
C39345 INVX1_LOC_136/A NAND2X1_LOC_849/B 0.03fF
C39346 INVX1_LOC_225/A NOR2X1_LOC_675/A -0.01fF
C39347 NOR2X1_LOC_859/A INVX1_LOC_280/A 0.01fF
C39348 INVX1_LOC_136/A INVX1_LOC_38/A 0.11fF
C39349 NAND2X1_LOC_837/Y NOR2X1_LOC_492/a_36_216# 0.00fF
C39350 INVX1_LOC_90/A NAND2X1_LOC_862/Y 0.04fF
C39351 NOR2X1_LOC_713/B NOR2X1_LOC_706/B 0.04fF
C39352 NOR2X1_LOC_561/Y INVX1_LOC_73/A 2.02fF
C39353 INVX1_LOC_269/A INVX1_LOC_84/A 0.20fF
C39354 NOR2X1_LOC_636/A VDD -0.00fF
C39355 NOR2X1_LOC_232/Y INVX1_LOC_84/A 0.01fF
C39356 NAND2X1_LOC_341/A INVX1_LOC_6/A 1.54fF
C39357 NAND2X1_LOC_560/A NOR2X1_LOC_525/Y 0.00fF
C39358 NOR2X1_LOC_667/A INVX1_LOC_91/A 0.09fF
C39359 INVX1_LOC_30/Y NOR2X1_LOC_83/Y 0.01fF
C39360 INVX1_LOC_248/A INVX1_LOC_91/A 0.68fF
C39361 NOR2X1_LOC_45/B NAND2X1_LOC_850/Y 0.07fF
C39362 INVX1_LOC_11/A INVX1_LOC_119/Y 0.02fF
C39363 INVX1_LOC_41/A NAND2X1_LOC_266/a_36_24# 0.00fF
C39364 NOR2X1_LOC_503/Y NOR2X1_LOC_697/Y 0.12fF
C39365 INVX1_LOC_77/A INVX1_LOC_117/A 0.42fF
C39366 NOR2X1_LOC_103/Y INVX1_LOC_3/A 0.09fF
C39367 INVX1_LOC_45/A NAND2X1_LOC_93/B 0.03fF
C39368 NOR2X1_LOC_92/Y INVX1_LOC_49/Y 0.05fF
C39369 NOR2X1_LOC_544/A NOR2X1_LOC_78/A 0.01fF
C39370 INVX1_LOC_71/A NOR2X1_LOC_536/A 0.33fF
C39371 NOR2X1_LOC_590/A NAND2X1_LOC_288/A 0.01fF
C39372 NOR2X1_LOC_223/a_36_216# INVX1_LOC_91/A 0.00fF
C39373 NOR2X1_LOC_521/Y INVX1_LOC_309/A 0.22fF
C39374 NOR2X1_LOC_667/A INVX1_LOC_11/Y 0.03fF
C39375 NOR2X1_LOC_78/B NOR2X1_LOC_657/B 0.03fF
C39376 NOR2X1_LOC_617/Y INVX1_LOC_280/A 0.02fF
C39377 NAND2X1_LOC_357/B NOR2X1_LOC_280/Y 0.04fF
C39378 NOR2X1_LOC_792/a_36_216# NAND2X1_LOC_807/B 0.00fF
C39379 NOR2X1_LOC_248/Y NOR2X1_LOC_155/A 0.06fF
C39380 INVX1_LOC_299/A NOR2X1_LOC_777/B 0.03fF
C39381 NOR2X1_LOC_377/Y INVX1_LOC_37/A 0.01fF
C39382 NOR2X1_LOC_431/Y INVX1_LOC_118/A 0.05fF
C39383 INVX1_LOC_208/A NOR2X1_LOC_405/A 0.48fF
C39384 NOR2X1_LOC_203/Y NAND2X1_LOC_447/Y 0.37fF
C39385 NOR2X1_LOC_465/a_36_216# NOR2X1_LOC_465/Y 0.01fF
C39386 NAND2X1_LOC_568/A INVX1_LOC_49/Y 0.03fF
C39387 NOR2X1_LOC_401/Y INVX1_LOC_20/A 0.01fF
C39388 INVX1_LOC_177/A NOR2X1_LOC_137/Y 0.73fF
C39389 INVX1_LOC_64/A NOR2X1_LOC_465/Y 0.09fF
C39390 INVX1_LOC_14/A NAND2X1_LOC_807/B 0.03fF
C39391 INVX1_LOC_134/A NOR2X1_LOC_856/B 0.06fF
C39392 INVX1_LOC_47/A NOR2X1_LOC_188/A 0.01fF
C39393 NOR2X1_LOC_93/Y INVX1_LOC_15/A 0.00fF
C39394 NOR2X1_LOC_329/B INVX1_LOC_75/A 0.03fF
C39395 NOR2X1_LOC_13/Y INVX1_LOC_291/A 0.10fF
C39396 INVX1_LOC_45/A INVX1_LOC_3/A 0.03fF
C39397 NOR2X1_LOC_637/a_36_216# INVX1_LOC_118/A 0.02fF
C39398 NAND2X1_LOC_357/B NAND2X1_LOC_811/B 0.03fF
C39399 INVX1_LOC_47/A NOR2X1_LOC_548/B 0.03fF
C39400 INVX1_LOC_71/A NAND2X1_LOC_93/B 4.28fF
C39401 INVX1_LOC_5/A NAND2X1_LOC_72/B 0.03fF
C39402 NOR2X1_LOC_528/Y NAND2X1_LOC_808/A 0.01fF
C39403 INVX1_LOC_11/A INVX1_LOC_284/A 0.07fF
C39404 INVX1_LOC_223/A NAND2X1_LOC_475/Y 0.29fF
C39405 INVX1_LOC_249/A INVX1_LOC_92/A 0.16fF
C39406 NOR2X1_LOC_590/A INVX1_LOC_19/A 0.18fF
C39407 INVX1_LOC_14/A NOR2X1_LOC_48/B 0.02fF
C39408 INVX1_LOC_57/A INVX1_LOC_29/Y 0.73fF
C39409 NOR2X1_LOC_303/Y INVX1_LOC_307/A 0.07fF
C39410 NAND2X1_LOC_672/a_36_24# NOR2X1_LOC_814/A 0.00fF
C39411 NOR2X1_LOC_773/Y INVX1_LOC_37/A 0.07fF
C39412 NOR2X1_LOC_456/Y NOR2X1_LOC_748/A 0.10fF
C39413 NOR2X1_LOC_140/A INVX1_LOC_32/A 0.02fF
C39414 NOR2X1_LOC_500/A NOR2X1_LOC_445/B 0.04fF
C39415 INVX1_LOC_71/A NAND2X1_LOC_425/Y 0.06fF
C39416 NOR2X1_LOC_303/Y NOR2X1_LOC_445/B 0.10fF
C39417 INVX1_LOC_271/A INVX1_LOC_53/A 0.03fF
C39418 NOR2X1_LOC_153/a_36_216# INVX1_LOC_6/A 0.00fF
C39419 INVX1_LOC_48/Y NOR2X1_LOC_38/B 0.07fF
C39420 NOR2X1_LOC_516/B NOR2X1_LOC_857/A 0.10fF
C39421 NOR2X1_LOC_548/Y NOR2X1_LOC_35/Y 0.10fF
C39422 NOR2X1_LOC_160/B INVX1_LOC_109/Y 0.07fF
C39423 INVX1_LOC_269/A INVX1_LOC_15/A 0.14fF
C39424 INVX1_LOC_102/Y INVX1_LOC_126/Y 0.01fF
C39425 VDD INVX1_LOC_56/Y 0.44fF
C39426 NOR2X1_LOC_346/B NAND2X1_LOC_96/A 0.07fF
C39427 NOR2X1_LOC_820/A INVX1_LOC_63/A 0.03fF
C39428 D_INPUT_6 NOR2X1_LOC_30/Y 0.55fF
C39429 NOR2X1_LOC_68/A NAND2X1_LOC_782/B 0.04fF
C39430 NOR2X1_LOC_785/Y INVX1_LOC_143/Y 0.00fF
C39431 NOR2X1_LOC_254/Y INVX1_LOC_307/A 0.09fF
C39432 NOR2X1_LOC_152/Y NOR2X1_LOC_697/Y 0.01fF
C39433 INVX1_LOC_11/Y NAND2X1_LOC_804/a_36_24# 0.01fF
C39434 NOR2X1_LOC_344/A NOR2X1_LOC_197/B 0.02fF
C39435 INVX1_LOC_71/A INVX1_LOC_3/A 0.29fF
C39436 NAND2X1_LOC_437/a_36_24# NOR2X1_LOC_440/B 0.02fF
C39437 NOR2X1_LOC_687/Y INVX1_LOC_117/A 0.03fF
C39438 INVX1_LOC_122/Y INVX1_LOC_29/A 0.08fF
C39439 INVX1_LOC_35/A NOR2X1_LOC_392/Y 0.07fF
C39440 INVX1_LOC_75/A NAND2X1_LOC_4/a_36_24# 0.00fF
C39441 NAND2X1_LOC_608/a_36_24# INVX1_LOC_29/Y 0.00fF
C39442 INVX1_LOC_30/A INVX1_LOC_102/A 0.33fF
C39443 NOR2X1_LOC_510/Y NOR2X1_LOC_677/Y 0.22fF
C39444 INVX1_LOC_72/A NOR2X1_LOC_89/A 0.04fF
C39445 INVX1_LOC_206/A INVX1_LOC_92/A 0.07fF
C39446 NOR2X1_LOC_76/A INVX1_LOC_76/A 0.03fF
C39447 NAND2X1_LOC_538/Y NAND2X1_LOC_175/Y 0.07fF
C39448 NAND2X1_LOC_799/A INVX1_LOC_94/Y 0.05fF
C39449 NOR2X1_LOC_45/B INVX1_LOC_282/A 0.14fF
C39450 NOR2X1_LOC_598/B INVX1_LOC_50/Y 0.14fF
C39451 NAND2X1_LOC_36/A D_INPUT_5 0.55fF
C39452 INVX1_LOC_173/Y VDD 0.63fF
C39453 NAND2X1_LOC_514/a_36_24# INVX1_LOC_9/A 0.00fF
C39454 INVX1_LOC_54/Y NOR2X1_LOC_445/B 0.34fF
C39455 INVX1_LOC_311/A INVX1_LOC_91/A 0.03fF
C39456 INVX1_LOC_27/A INVX1_LOC_53/A 0.15fF
C39457 INVX1_LOC_315/A INVX1_LOC_63/A 0.01fF
C39458 NOR2X1_LOC_32/B INVX1_LOC_39/A 0.08fF
C39459 INVX1_LOC_58/A NOR2X1_LOC_454/Y 0.19fF
C39460 NAND2X1_LOC_793/Y NOR2X1_LOC_301/A 0.03fF
C39461 NAND2X1_LOC_141/A NAND2X1_LOC_574/A 0.01fF
C39462 INVX1_LOC_232/A NOR2X1_LOC_99/Y 0.15fF
C39463 INVX1_LOC_35/A INVX1_LOC_235/A 0.01fF
C39464 NOR2X1_LOC_329/B NAND2X1_LOC_453/A 0.07fF
C39465 INVX1_LOC_14/A NAND2X1_LOC_215/A 0.17fF
C39466 NOR2X1_LOC_123/B NOR2X1_LOC_536/A 0.13fF
C39467 NAND2X1_LOC_778/Y NAND2X1_LOC_35/Y 0.04fF
C39468 INVX1_LOC_33/A NAND2X1_LOC_74/B 0.16fF
C39469 NOR2X1_LOC_329/B NOR2X1_LOC_65/a_36_216# 0.01fF
C39470 INVX1_LOC_96/Y INVX1_LOC_136/Y 0.01fF
C39471 NOR2X1_LOC_385/Y VDD 0.00fF
C39472 NOR2X1_LOC_250/Y INVX1_LOC_50/A 0.01fF
C39473 INVX1_LOC_266/A NOR2X1_LOC_598/B 0.02fF
C39474 INVX1_LOC_226/Y INVX1_LOC_35/Y 0.00fF
C39475 INVX1_LOC_140/A INVX1_LOC_37/A 0.07fF
C39476 INVX1_LOC_1/Y NOR2X1_LOC_79/Y 0.28fF
C39477 NOR2X1_LOC_383/Y NOR2X1_LOC_99/Y 0.03fF
C39478 INVX1_LOC_77/A NOR2X1_LOC_460/A 0.01fF
C39479 NOR2X1_LOC_590/A INVX1_LOC_26/Y 0.92fF
C39480 NAND2X1_LOC_477/A INVX1_LOC_49/Y 0.01fF
C39481 NOR2X1_LOC_78/A NOR2X1_LOC_139/Y 0.36fF
C39482 INVX1_LOC_22/Y INVX1_LOC_26/Y 0.50fF
C39483 INVX1_LOC_18/A INVX1_LOC_94/Y 0.07fF
C39484 NOR2X1_LOC_137/A INVX1_LOC_54/A 0.01fF
C39485 NOR2X1_LOC_789/a_36_216# INVX1_LOC_46/Y 0.01fF
C39486 NAND2X1_LOC_563/A INVX1_LOC_84/A 0.03fF
C39487 INVX1_LOC_135/A INVX1_LOC_185/A 0.01fF
C39488 NOR2X1_LOC_432/Y INVX1_LOC_186/Y 0.01fF
C39489 NOR2X1_LOC_602/a_36_216# NAND2X1_LOC_175/Y 0.01fF
C39490 NAND2X1_LOC_35/Y NOR2X1_LOC_15/Y 0.08fF
C39491 NOR2X1_LOC_254/A INVX1_LOC_23/A 0.16fF
C39492 NOR2X1_LOC_360/Y INVX1_LOC_87/A 0.03fF
C39493 INVX1_LOC_40/A INVX1_LOC_293/Y 0.00fF
C39494 NOR2X1_LOC_52/B INVX1_LOC_284/A 0.68fF
C39495 INVX1_LOC_230/Y NOR2X1_LOC_416/A 0.04fF
C39496 NOR2X1_LOC_78/A NAND2X1_LOC_468/B 0.03fF
C39497 D_INPUT_1 NOR2X1_LOC_644/B 0.02fF
C39498 NOR2X1_LOC_285/Y NOR2X1_LOC_286/Y 0.00fF
C39499 INVX1_LOC_224/Y NOR2X1_LOC_606/Y 0.02fF
C39500 INVX1_LOC_54/Y INVX1_LOC_12/A 0.07fF
C39501 INVX1_LOC_226/Y NOR2X1_LOC_721/B 0.02fF
C39502 INVX1_LOC_232/Y INVX1_LOC_29/A 0.03fF
C39503 NAND2X1_LOC_722/A INVX1_LOC_102/A 0.03fF
C39504 NOR2X1_LOC_237/Y NAND2X1_LOC_471/Y 0.01fF
C39505 NOR2X1_LOC_537/Y NOR2X1_LOC_89/A 0.03fF
C39506 NAND2X1_LOC_338/B NOR2X1_LOC_89/A 0.19fF
C39507 INVX1_LOC_58/A NAND2X1_LOC_569/a_36_24# 0.00fF
C39508 INVX1_LOC_18/A INVX1_LOC_296/A 0.12fF
C39509 INVX1_LOC_40/A NAND2X1_LOC_74/B 0.06fF
C39510 INVX1_LOC_36/A NOR2X1_LOC_696/Y 0.07fF
C39511 NOR2X1_LOC_644/A INVX1_LOC_179/A 0.00fF
C39512 NAND2X1_LOC_729/B INVX1_LOC_76/A 0.01fF
C39513 INVX1_LOC_140/A NOR2X1_LOC_177/Y 0.16fF
C39514 INVX1_LOC_200/A INVX1_LOC_93/A 0.08fF
C39515 NOR2X1_LOC_156/A NOR2X1_LOC_155/A 0.07fF
C39516 NAND2X1_LOC_138/a_36_24# INVX1_LOC_9/A 0.00fF
C39517 INVX1_LOC_164/A INVX1_LOC_63/A 1.69fF
C39518 INPUT_0 NOR2X1_LOC_119/a_36_216# 0.00fF
C39519 INVX1_LOC_27/A NAND2X1_LOC_522/a_36_24# -0.00fF
C39520 NOR2X1_LOC_471/Y INVX1_LOC_298/A 0.02fF
C39521 NAND2X1_LOC_392/A INVX1_LOC_29/A 0.01fF
C39522 NOR2X1_LOC_403/a_36_216# INVX1_LOC_23/Y 0.01fF
C39523 D_GATE_366 INVX1_LOC_113/A 0.07fF
C39524 INVX1_LOC_17/A D_INPUT_6 0.26fF
C39525 INVX1_LOC_21/A NOR2X1_LOC_592/A 0.01fF
C39526 INVX1_LOC_233/A NAND2X1_LOC_185/a_36_24# 0.01fF
C39527 INVX1_LOC_17/A NOR2X1_LOC_173/Y 0.23fF
C39528 NAND2X1_LOC_773/Y INVX1_LOC_1/A 0.21fF
C39529 NOR2X1_LOC_175/A NAND2X1_LOC_278/a_36_24# 0.00fF
C39530 NOR2X1_LOC_84/Y NOR2X1_LOC_38/B 0.16fF
C39531 NOR2X1_LOC_137/B NOR2X1_LOC_137/Y 0.02fF
C39532 NOR2X1_LOC_763/Y INVX1_LOC_19/A 0.02fF
C39533 INVX1_LOC_64/A NOR2X1_LOC_52/Y 0.01fF
C39534 NOR2X1_LOC_366/Y INVX1_LOC_272/A 0.02fF
C39535 NOR2X1_LOC_537/Y INVX1_LOC_104/Y 0.09fF
C39536 INVX1_LOC_103/A NOR2X1_LOC_205/Y 2.61fF
C39537 NOR2X1_LOC_790/A INVX1_LOC_292/A 0.01fF
C39538 NAND2X1_LOC_706/Y NAND2X1_LOC_550/A 0.01fF
C39539 INVX1_LOC_58/A INVX1_LOC_77/A 7.33fF
C39540 INPUT_3 NAND2X1_LOC_218/A 0.01fF
C39541 NAND2X1_LOC_468/B NOR2X1_LOC_60/Y 0.00fF
C39542 INPUT_3 NOR2X1_LOC_140/A 0.03fF
C39543 NOR2X1_LOC_570/B NOR2X1_LOC_383/B 0.23fF
C39544 NOR2X1_LOC_791/B INVX1_LOC_306/Y 0.11fF
C39545 INVX1_LOC_233/A INVX1_LOC_314/Y 0.07fF
C39546 NOR2X1_LOC_718/B NAND2X1_LOC_299/a_36_24# 0.01fF
C39547 NOR2X1_LOC_205/Y INVX1_LOC_292/A 0.05fF
C39548 NAND2X1_LOC_803/B INVX1_LOC_161/Y 0.03fF
C39549 INVX1_LOC_256/A NOR2X1_LOC_541/Y 0.04fF
C39550 NOR2X1_LOC_614/a_36_216# INVX1_LOC_77/A 0.00fF
C39551 NOR2X1_LOC_703/A INVX1_LOC_19/A 0.03fF
C39552 INVX1_LOC_49/A INVX1_LOC_292/Y 0.13fF
C39553 INVX1_LOC_24/A NOR2X1_LOC_291/Y 0.28fF
C39554 INVX1_LOC_289/A INVX1_LOC_78/A 0.01fF
C39555 INVX1_LOC_313/Y NOR2X1_LOC_89/A 0.01fF
C39556 INVX1_LOC_96/A NOR2X1_LOC_155/A 0.74fF
C39557 INVX1_LOC_60/Y INVX1_LOC_57/A 0.08fF
C39558 NOR2X1_LOC_75/Y INVX1_LOC_55/A 0.06fF
C39559 NOR2X1_LOC_690/A NAND2X1_LOC_827/a_36_24# 0.00fF
C39560 NAND2X1_LOC_358/B INVX1_LOC_33/A 0.01fF
C39561 NOR2X1_LOC_590/A INVX1_LOC_161/Y 0.03fF
C39562 NOR2X1_LOC_443/Y INVX1_LOC_143/A 0.03fF
C39563 NOR2X1_LOC_591/Y NOR2X1_LOC_591/A 0.09fF
C39564 NOR2X1_LOC_598/B NOR2X1_LOC_6/B 0.01fF
C39565 INVX1_LOC_200/Y INVX1_LOC_2/A 0.03fF
C39566 NOR2X1_LOC_106/A INVX1_LOC_32/A 0.05fF
C39567 NAND2X1_LOC_639/A NAND2X1_LOC_635/a_36_24# 0.03fF
C39568 INVX1_LOC_299/A INVX1_LOC_18/A 1.08fF
C39569 NOR2X1_LOC_814/Y INVX1_LOC_15/A 0.05fF
C39570 INVX1_LOC_1/Y INVX1_LOC_26/A 0.03fF
C39571 INVX1_LOC_256/A INVX1_LOC_45/A 0.87fF
C39572 NOR2X1_LOC_78/B INVX1_LOC_271/A 0.03fF
C39573 INVX1_LOC_206/A INVX1_LOC_53/A 0.01fF
C39574 INVX1_LOC_200/Y NOR2X1_LOC_226/A 0.01fF
C39575 INVX1_LOC_223/A NOR2X1_LOC_457/A 0.03fF
C39576 INVX1_LOC_233/Y INVX1_LOC_240/A 0.10fF
C39577 NOR2X1_LOC_540/B INVX1_LOC_179/A 0.01fF
C39578 INVX1_LOC_11/A INVX1_LOC_72/A 0.07fF
C39579 INVX1_LOC_17/A INVX1_LOC_205/A 0.02fF
C39580 INVX1_LOC_269/A NOR2X1_LOC_168/Y 0.01fF
C39581 INVX1_LOC_256/A NOR2X1_LOC_568/A 0.16fF
C39582 NOR2X1_LOC_15/Y INVX1_LOC_94/A 0.03fF
C39583 NOR2X1_LOC_160/B NOR2X1_LOC_726/Y 0.04fF
C39584 NOR2X1_LOC_272/Y INVX1_LOC_155/A 0.00fF
C39585 INVX1_LOC_117/A INVX1_LOC_9/A 0.19fF
C39586 NOR2X1_LOC_590/A INVX1_LOC_312/A 0.01fF
C39587 NOR2X1_LOC_124/B INVX1_LOC_306/Y 0.02fF
C39588 INVX1_LOC_230/Y INVX1_LOC_36/A 0.03fF
C39589 INVX1_LOC_17/A NOR2X1_LOC_607/A 0.01fF
C39590 NAND2X1_LOC_801/a_36_24# NOR2X1_LOC_409/B 0.00fF
C39591 NAND2X1_LOC_105/a_36_24# INVX1_LOC_94/Y 0.00fF
C39592 NAND2X1_LOC_198/B NAND2X1_LOC_337/B 0.10fF
C39593 NAND2X1_LOC_149/Y INVX1_LOC_63/Y 0.10fF
C39594 INVX1_LOC_50/A NAND2X1_LOC_660/Y 0.01fF
C39595 INVX1_LOC_226/Y NAND2X1_LOC_860/A 0.01fF
C39596 INVX1_LOC_55/Y NOR2X1_LOC_334/Y 0.08fF
C39597 NAND2X1_LOC_555/Y INVX1_LOC_205/A 0.39fF
C39598 VDD NOR2X1_LOC_831/B 0.39fF
C39599 NAND2X1_LOC_347/B NOR2X1_LOC_557/Y 0.01fF
C39600 INVX1_LOC_64/A NOR2X1_LOC_458/B 0.03fF
C39601 NAND2X1_LOC_787/A NAND2X1_LOC_543/Y 0.01fF
C39602 INVX1_LOC_34/A NOR2X1_LOC_92/Y 0.20fF
C39603 INVX1_LOC_223/A INVX1_LOC_30/A 0.01fF
C39604 INVX1_LOC_256/A INVX1_LOC_71/A 0.54fF
C39605 NOR2X1_LOC_690/A NAND2X1_LOC_579/A 0.08fF
C39606 NOR2X1_LOC_478/A NOR2X1_LOC_68/A 0.02fF
C39607 NOR2X1_LOC_91/A NAND2X1_LOC_567/a_36_24# 0.01fF
C39608 INVX1_LOC_2/A NOR2X1_LOC_406/A 0.07fF
C39609 NOR2X1_LOC_641/B NOR2X1_LOC_751/Y 0.03fF
C39610 INVX1_LOC_35/A INVX1_LOC_25/Y 1.57fF
C39611 NOR2X1_LOC_121/A NOR2X1_LOC_392/Y 0.10fF
C39612 NAND2X1_LOC_214/B NOR2X1_LOC_78/B 0.07fF
C39613 NOR2X1_LOC_135/Y INVX1_LOC_128/Y 0.00fF
C39614 INVX1_LOC_256/A NAND2X1_LOC_330/a_36_24# 0.06fF
C39615 NAND2X1_LOC_563/Y INVX1_LOC_239/A 0.01fF
C39616 NOR2X1_LOC_32/B NAND2X1_LOC_735/B 0.01fF
C39617 NOR2X1_LOC_226/A NOR2X1_LOC_406/A 0.03fF
C39618 INVX1_LOC_50/A D_INPUT_0 0.09fF
C39619 INVX1_LOC_83/A INVX1_LOC_271/A 0.03fF
C39620 NOR2X1_LOC_355/A INVX1_LOC_57/A 0.07fF
C39621 NOR2X1_LOC_15/Y NOR2X1_LOC_234/Y -0.03fF
C39622 NOR2X1_LOC_331/B NAND2X1_LOC_93/B 0.07fF
C39623 NOR2X1_LOC_536/A NOR2X1_LOC_491/Y 0.01fF
C39624 NOR2X1_LOC_219/Y INVX1_LOC_5/A 0.22fF
C39625 INVX1_LOC_251/Y NOR2X1_LOC_440/B 0.09fF
C39626 NAND2X1_LOC_860/A INVX1_LOC_10/A 0.01fF
C39627 INVX1_LOC_27/A NOR2X1_LOC_78/B 0.34fF
C39628 NAND2X1_LOC_740/Y NAND2X1_LOC_853/Y 0.03fF
C39629 INVX1_LOC_228/Y NOR2X1_LOC_84/A 0.07fF
C39630 INVX1_LOC_5/A NOR2X1_LOC_619/A 0.03fF
C39631 INVX1_LOC_45/A NOR2X1_LOC_781/Y 0.03fF
C39632 NOR2X1_LOC_468/Y NOR2X1_LOC_84/Y 0.19fF
C39633 NAND2X1_LOC_863/A NAND2X1_LOC_175/Y 0.16fF
C39634 NOR2X1_LOC_606/Y INVX1_LOC_71/A 0.00fF
C39635 NAND2X1_LOC_354/B INVX1_LOC_161/Y 0.03fF
C39636 INVX1_LOC_12/Y INVX1_LOC_84/A 0.02fF
C39637 NOR2X1_LOC_92/Y NAND2X1_LOC_231/Y 0.10fF
C39638 INVX1_LOC_280/Y INVX1_LOC_234/Y 0.15fF
C39639 INVX1_LOC_200/Y INPUT_1 0.05fF
C39640 INVX1_LOC_33/A NOR2X1_LOC_276/Y 0.01fF
C39641 NAND2X1_LOC_650/B INVX1_LOC_19/A 0.99fF
C39642 NAND2X1_LOC_347/B INVX1_LOC_143/A 0.00fF
C39643 NOR2X1_LOC_717/B NOR2X1_LOC_678/A 0.00fF
C39644 NOR2X1_LOC_753/Y INVX1_LOC_141/Y 0.03fF
C39645 NAND2X1_LOC_469/B INVX1_LOC_109/A 0.00fF
C39646 INVX1_LOC_5/A NOR2X1_LOC_665/A 0.04fF
C39647 NOR2X1_LOC_433/A NOR2X1_LOC_361/a_36_216# 0.01fF
C39648 NOR2X1_LOC_456/Y INVX1_LOC_89/A 0.08fF
C39649 NOR2X1_LOC_473/B INVX1_LOC_23/A 0.00fF
C39650 INVX1_LOC_108/Y NOR2X1_LOC_814/Y 0.02fF
C39651 NOR2X1_LOC_496/Y INVX1_LOC_16/A 0.05fF
C39652 NOR2X1_LOC_655/B INVX1_LOC_14/A 0.03fF
C39653 INVX1_LOC_5/A NOR2X1_LOC_781/B 0.07fF
C39654 NOR2X1_LOC_91/A NOR2X1_LOC_322/Y 0.03fF
C39655 INVX1_LOC_244/Y NOR2X1_LOC_582/Y 0.01fF
C39656 INVX1_LOC_225/Y INVX1_LOC_104/A 0.12fF
C39657 NOR2X1_LOC_296/Y NOR2X1_LOC_709/A 1.02fF
C39658 NOR2X1_LOC_2/Y NOR2X1_LOC_47/a_36_216# 0.00fF
C39659 NAND2X1_LOC_287/B INVX1_LOC_29/A 0.13fF
C39660 INVX1_LOC_224/A NOR2X1_LOC_537/Y 0.03fF
C39661 NAND2X1_LOC_325/Y INVX1_LOC_141/Y 0.03fF
C39662 NAND2X1_LOC_207/a_36_24# INVX1_LOC_83/A 0.01fF
C39663 NOR2X1_LOC_433/A INVX1_LOC_72/A 0.07fF
C39664 INVX1_LOC_11/A INVX1_LOC_192/Y 0.02fF
C39665 INVX1_LOC_21/A NOR2X1_LOC_553/B 0.03fF
C39666 NAND2X1_LOC_35/Y NOR2X1_LOC_576/B 2.12fF
C39667 INVX1_LOC_11/A NOR2X1_LOC_537/Y 0.46fF
C39668 NOR2X1_LOC_598/B NOR2X1_LOC_156/A 0.03fF
C39669 INVX1_LOC_11/A NAND2X1_LOC_338/B 0.10fF
C39670 NAND2X1_LOC_214/B INVX1_LOC_83/A 0.01fF
C39671 NOR2X1_LOC_355/A NAND2X1_LOC_608/a_36_24# 0.00fF
C39672 INVX1_LOC_8/Y NAND2X1_LOC_364/A 0.02fF
C39673 NOR2X1_LOC_717/Y NOR2X1_LOC_142/Y 0.07fF
C39674 INVX1_LOC_109/Y NAND2X1_LOC_211/Y 0.09fF
C39675 INVX1_LOC_100/A NAND2X1_LOC_99/A 0.07fF
C39676 INVX1_LOC_136/A INVX1_LOC_33/A 0.06fF
C39677 NOR2X1_LOC_275/A INVX1_LOC_15/A 0.04fF
C39678 INVX1_LOC_276/Y INVX1_LOC_161/Y 0.01fF
C39679 INVX1_LOC_214/Y NOR2X1_LOC_513/Y 0.15fF
C39680 NAND2X1_LOC_96/A NOR2X1_LOC_777/B 1.04fF
C39681 INVX1_LOC_286/Y NAND2X1_LOC_357/B 0.10fF
C39682 NAND2X1_LOC_348/A NOR2X1_LOC_414/Y 0.01fF
C39683 INVX1_LOC_11/A NAND2X1_LOC_323/B 0.08fF
C39684 NOR2X1_LOC_361/B INVX1_LOC_56/Y 0.03fF
C39685 INVX1_LOC_291/A NOR2X1_LOC_697/Y 0.00fF
C39686 NAND2X1_LOC_550/A NAND2X1_LOC_483/a_36_24# 0.00fF
C39687 INVX1_LOC_37/A INVX1_LOC_42/A 0.12fF
C39688 INVX1_LOC_27/A INVX1_LOC_83/A 0.13fF
C39689 NAND2X1_LOC_208/B NOR2X1_LOC_398/Y 0.30fF
C39690 NAND2X1_LOC_112/Y INVX1_LOC_88/A 0.02fF
C39691 VDD NAND2X1_LOC_430/B 0.02fF
C39692 INVX1_LOC_58/A NAND2X1_LOC_832/Y 0.05fF
C39693 INVX1_LOC_108/A NOR2X1_LOC_814/A 0.03fF
C39694 INVX1_LOC_286/A NOR2X1_LOC_383/B 0.07fF
C39695 NOR2X1_LOC_67/A INVX1_LOC_39/Y 0.05fF
C39696 NOR2X1_LOC_151/Y NOR2X1_LOC_678/A 0.00fF
C39697 INVX1_LOC_289/A NOR2X1_LOC_503/Y 0.00fF
C39698 NOR2X1_LOC_738/Y NOR2X1_LOC_687/Y 0.05fF
C39699 NOR2X1_LOC_52/B INVX1_LOC_72/A 0.13fF
C39700 NAND2X1_LOC_92/a_36_24# INVX1_LOC_3/A 0.00fF
C39701 NOR2X1_LOC_660/a_36_216# INVX1_LOC_63/A 0.00fF
C39702 INVX1_LOC_35/A INVX1_LOC_75/A 4.24fF
C39703 NAND2X1_LOC_337/B INVX1_LOC_53/Y 0.07fF
C39704 NOR2X1_LOC_315/Y INVX1_LOC_18/A 0.03fF
C39705 NAND2X1_LOC_537/Y INVX1_LOC_10/A 0.07fF
C39706 NAND2X1_LOC_36/A NAND2X1_LOC_451/Y 0.03fF
C39707 INVX1_LOC_34/A NAND2X1_LOC_837/Y 0.08fF
C39708 INVX1_LOC_93/Y INVX1_LOC_26/A 0.01fF
C39709 NAND2X1_LOC_361/a_36_24# NAND2X1_LOC_656/A 0.01fF
C39710 INVX1_LOC_250/A INVX1_LOC_2/A 0.01fF
C39711 NAND2X1_LOC_361/Y INVX1_LOC_49/A 0.07fF
C39712 NOR2X1_LOC_537/A NAND2X1_LOC_536/a_36_24# 0.00fF
C39713 INVX1_LOC_14/A NOR2X1_LOC_99/B 0.07fF
C39714 NOR2X1_LOC_432/Y INVX1_LOC_18/A 0.01fF
C39715 NOR2X1_LOC_355/B INVX1_LOC_23/A 0.03fF
C39716 NOR2X1_LOC_389/A INVX1_LOC_290/A 0.10fF
C39717 INVX1_LOC_227/A INVX1_LOC_161/Y 0.10fF
C39718 NOR2X1_LOC_793/A NOR2X1_LOC_542/Y 0.02fF
C39719 INVX1_LOC_279/A NOR2X1_LOC_794/B 0.02fF
C39720 NOR2X1_LOC_246/A INVX1_LOC_308/Y 0.03fF
C39721 NOR2X1_LOC_790/B NOR2X1_LOC_337/Y 0.02fF
C39722 NOR2X1_LOC_681/Y INVX1_LOC_78/A 0.00fF
C39723 NOR2X1_LOC_15/Y NAND2X1_LOC_307/a_36_24# 0.00fF
C39724 INVX1_LOC_78/A INVX1_LOC_37/A 0.15fF
C39725 NOR2X1_LOC_831/B INVX1_LOC_133/A 0.02fF
C39726 NOR2X1_LOC_220/A NAND2X1_LOC_272/a_36_24# 0.00fF
C39727 NAND2X1_LOC_199/B INVX1_LOC_290/A 0.06fF
C39728 INVX1_LOC_136/A INVX1_LOC_40/A 0.08fF
C39729 INVX1_LOC_41/A INVX1_LOC_34/A 0.03fF
C39730 INVX1_LOC_256/A NOR2X1_LOC_123/B 0.00fF
C39731 NAND2X1_LOC_9/Y NOR2X1_LOC_557/A 0.02fF
C39732 INVX1_LOC_136/A NAND2X1_LOC_726/Y 0.02fF
C39733 NOR2X1_LOC_89/A NOR2X1_LOC_79/a_36_216# 0.03fF
C39734 NOR2X1_LOC_498/Y INVX1_LOC_34/A 0.02fF
C39735 INVX1_LOC_30/A NAND2X1_LOC_662/Y 0.11fF
C39736 NAND2X1_LOC_198/B NOR2X1_LOC_773/Y 0.10fF
C39737 NAND2X1_LOC_287/B NOR2X1_LOC_281/Y 0.03fF
C39738 INVX1_LOC_232/Y INVX1_LOC_228/A 0.01fF
C39739 NAND2X1_LOC_84/Y NOR2X1_LOC_655/B 0.06fF
C39740 INVX1_LOC_11/A INVX1_LOC_313/Y 0.07fF
C39741 NAND2X1_LOC_53/Y INVX1_LOC_85/Y 0.02fF
C39742 INVX1_LOC_136/A NOR2X1_LOC_605/B 0.00fF
C39743 INVX1_LOC_249/A NOR2X1_LOC_78/B 0.04fF
C39744 NOR2X1_LOC_590/A INVX1_LOC_62/A 0.02fF
C39745 INVX1_LOC_2/A NAND2X1_LOC_361/Y 0.03fF
C39746 NAND2X1_LOC_45/a_36_24# INVX1_LOC_64/Y 0.00fF
C39747 INVX1_LOC_290/A INVX1_LOC_107/A 0.05fF
C39748 NAND2X1_LOC_560/a_36_24# NOR2X1_LOC_380/Y 0.01fF
C39749 NOR2X1_LOC_181/A NOR2X1_LOC_678/A 0.01fF
C39750 NOR2X1_LOC_92/Y INPUT_0 0.17fF
C39751 NAND2X1_LOC_656/A INVX1_LOC_22/A 0.10fF
C39752 INVX1_LOC_258/Y INVX1_LOC_309/A 0.36fF
C39753 INVX1_LOC_41/A NAND2X1_LOC_231/Y 0.00fF
C39754 INVX1_LOC_57/Y NOR2X1_LOC_373/Y 0.20fF
C39755 INVX1_LOC_271/A INVX1_LOC_46/A 0.07fF
C39756 INVX1_LOC_24/Y INPUT_0 0.26fF
C39757 NAND2X1_LOC_784/A NOR2X1_LOC_305/Y 0.09fF
C39758 NAND2X1_LOC_96/A NOR2X1_LOC_843/B 0.07fF
C39759 INVX1_LOC_13/Y NOR2X1_LOC_78/A 1.27fF
C39760 INVX1_LOC_290/A NOR2X1_LOC_596/A 0.10fF
C39761 INVX1_LOC_232/Y NOR2X1_LOC_516/a_36_216# 0.00fF
C39762 INVX1_LOC_105/Y INVX1_LOC_46/A 0.24fF
C39763 INVX1_LOC_256/A INVX1_LOC_102/Y 0.57fF
C39764 INVX1_LOC_104/A INVX1_LOC_266/Y 0.02fF
C39765 NAND2X1_LOC_574/A NOR2X1_LOC_128/a_36_216# 0.01fF
C39766 NOR2X1_LOC_111/A INVX1_LOC_57/A 0.01fF
C39767 NOR2X1_LOC_158/Y NAND2X1_LOC_637/Y 0.09fF
C39768 NOR2X1_LOC_209/A INVX1_LOC_213/A 0.01fF
C39769 INVX1_LOC_18/A INVX1_LOC_66/A 0.01fF
C39770 NOR2X1_LOC_502/Y INVX1_LOC_75/A 0.05fF
C39771 INVX1_LOC_265/A NAND2X1_LOC_850/Y 0.09fF
C39772 INVX1_LOC_290/Y NAND2X1_LOC_475/Y 0.10fF
C39773 NOR2X1_LOC_664/Y NOR2X1_LOC_78/B 0.01fF
C39774 NOR2X1_LOC_440/Y INVX1_LOC_71/A 0.10fF
C39775 NOR2X1_LOC_177/Y INVX1_LOC_78/A 0.03fF
C39776 NOR2X1_LOC_32/B D_INPUT_3 0.06fF
C39777 NAND2X1_LOC_231/Y NAND2X1_LOC_477/A 0.19fF
C39778 NAND2X1_LOC_338/B NOR2X1_LOC_52/B 0.01fF
C39779 INVX1_LOC_78/A NOR2X1_LOC_743/Y 0.01fF
C39780 INVX1_LOC_50/A NAND2X1_LOC_848/A 0.01fF
C39781 INVX1_LOC_152/Y INVX1_LOC_37/A 0.01fF
C39782 INVX1_LOC_63/Y INVX1_LOC_16/A 0.07fF
C39783 NOR2X1_LOC_322/Y INVX1_LOC_31/A 0.07fF
C39784 NOR2X1_LOC_67/Y INVX1_LOC_19/A 0.19fF
C39785 NAND2X1_LOC_154/Y INVX1_LOC_28/A 0.01fF
C39786 INVX1_LOC_36/A NOR2X1_LOC_153/a_36_216# 0.01fF
C39787 NAND2X1_LOC_470/B NOR2X1_LOC_592/B 0.35fF
C39788 INVX1_LOC_5/A NOR2X1_LOC_585/Y 0.09fF
C39789 NOR2X1_LOC_68/A NOR2X1_LOC_163/A 0.01fF
C39790 NOR2X1_LOC_655/B INVX1_LOC_111/Y 0.02fF
C39791 NOR2X1_LOC_300/Y NAND2X1_LOC_841/A 0.15fF
C39792 NOR2X1_LOC_189/A NAND2X1_LOC_795/Y 0.00fF
C39793 NAND2X1_LOC_717/Y NAND2X1_LOC_839/A 0.03fF
C39794 INVX1_LOC_106/Y NAND2X1_LOC_74/B 0.11fF
C39795 INVX1_LOC_13/Y NAND2X1_LOC_464/A 0.05fF
C39796 INVX1_LOC_17/Y INVX1_LOC_118/A 0.01fF
C39797 INVX1_LOC_88/A NOR2X1_LOC_78/A 0.03fF
C39798 NOR2X1_LOC_383/B INVX1_LOC_54/A 0.07fF
C39799 NOR2X1_LOC_740/Y INVX1_LOC_186/A 0.01fF
C39800 INVX1_LOC_54/Y NOR2X1_LOC_566/Y 0.01fF
C39801 INVX1_LOC_98/Y NOR2X1_LOC_191/A 0.25fF
C39802 INVX1_LOC_58/A INVX1_LOC_9/A 0.10fF
C39803 NOR2X1_LOC_598/B NOR2X1_LOC_684/Y 0.48fF
C39804 NAND2X1_LOC_391/Y INVX1_LOC_20/A 0.00fF
C39805 INVX1_LOC_263/A INVX1_LOC_266/Y 0.11fF
C39806 NAND2X1_LOC_169/Y VDD 0.01fF
C39807 NOR2X1_LOC_263/a_36_216# INVX1_LOC_22/A 0.00fF
C39808 NOR2X1_LOC_423/Y INVX1_LOC_22/A 0.05fF
C39809 INVX1_LOC_80/A NAND2X1_LOC_139/A 0.08fF
C39810 INVX1_LOC_92/Y INVX1_LOC_31/A 0.02fF
C39811 NAND2X1_LOC_254/Y INVX1_LOC_284/A 0.08fF
C39812 INVX1_LOC_89/A NOR2X1_LOC_550/B 0.03fF
C39813 NOR2X1_LOC_789/B VDD -0.00fF
C39814 INVX1_LOC_27/A INVX1_LOC_46/A 0.19fF
C39815 NOR2X1_LOC_824/A INVX1_LOC_46/A 0.07fF
C39816 INVX1_LOC_36/A NOR2X1_LOC_292/Y 0.03fF
C39817 INVX1_LOC_174/A INVX1_LOC_91/A 0.00fF
C39818 NAND2X1_LOC_366/A NAND2X1_LOC_367/B 0.05fF
C39819 NOR2X1_LOC_142/Y NOR2X1_LOC_137/A 0.10fF
C39820 NOR2X1_LOC_383/a_36_216# NOR2X1_LOC_315/Y 0.01fF
C39821 INVX1_LOC_26/Y NOR2X1_LOC_688/a_36_216# 0.00fF
C39822 INVX1_LOC_45/A INVX1_LOC_69/Y 0.14fF
C39823 NOR2X1_LOC_148/Y INVX1_LOC_213/A 0.02fF
C39824 NOR2X1_LOC_773/Y INVX1_LOC_53/Y 0.03fF
C39825 NOR2X1_LOC_593/Y INVX1_LOC_313/Y 0.07fF
C39826 NOR2X1_LOC_222/Y INVX1_LOC_22/A 0.03fF
C39827 NOR2X1_LOC_67/A NOR2X1_LOC_789/A 0.01fF
C39828 INVX1_LOC_2/A NAND2X1_LOC_319/A 0.03fF
C39829 NOR2X1_LOC_329/B NOR2X1_LOC_577/Y 0.63fF
C39830 NOR2X1_LOC_717/B NAND2X1_LOC_177/a_36_24# 0.00fF
C39831 INVX1_LOC_133/Y NAND2X1_LOC_656/Y 0.18fF
C39832 INVX1_LOC_13/A INVX1_LOC_218/A 0.02fF
C39833 INVX1_LOC_1/A NAND2X1_LOC_298/a_36_24# 0.00fF
C39834 INVX1_LOC_34/A NOR2X1_LOC_122/Y 0.11fF
C39835 INVX1_LOC_28/A INVX1_LOC_63/Y 0.03fF
C39836 INVX1_LOC_53/A NOR2X1_LOC_216/B 0.03fF
C39837 NOR2X1_LOC_45/Y NAND2X1_LOC_468/B 0.03fF
C39838 INVX1_LOC_210/Y NOR2X1_LOC_349/A 0.03fF
C39839 NOR2X1_LOC_78/A NOR2X1_LOC_500/B 2.53fF
C39840 NOR2X1_LOC_543/a_36_216# NOR2X1_LOC_568/A 0.01fF
C39841 INVX1_LOC_14/A NOR2X1_LOC_176/Y 0.02fF
C39842 NOR2X1_LOC_634/Y NOR2X1_LOC_445/B 0.25fF
C39843 NOR2X1_LOC_41/Y INVX1_LOC_89/A 0.05fF
C39844 D_GATE_741 VDD 0.35fF
C39845 INVX1_LOC_69/Y INVX1_LOC_71/A 0.29fF
C39846 NAND2X1_LOC_464/B NAND2X1_LOC_489/Y 0.05fF
C39847 INVX1_LOC_88/A NOR2X1_LOC_60/Y 0.01fF
C39848 NOR2X1_LOC_19/B INVX1_LOC_80/Y 0.01fF
C39849 NOR2X1_LOC_348/Y NOR2X1_LOC_331/B 0.07fF
C39850 NOR2X1_LOC_156/B NOR2X1_LOC_156/A 0.09fF
C39851 INVX1_LOC_90/A NAND2X1_LOC_342/Y 0.03fF
C39852 INVX1_LOC_30/A INVX1_LOC_314/A 0.01fF
C39853 NAND2X1_LOC_218/B NAND2X1_LOC_4/a_36_24# 0.00fF
C39854 INVX1_LOC_246/A NOR2X1_LOC_447/B 0.02fF
C39855 NAND2X1_LOC_352/B VDD 0.23fF
C39856 INVX1_LOC_41/A INPUT_0 0.23fF
C39857 NOR2X1_LOC_389/B NAND2X1_LOC_342/Y 0.00fF
C39858 INVX1_LOC_93/A INVX1_LOC_92/A 0.19fF
C39859 NOR2X1_LOC_849/A NOR2X1_LOC_862/B 0.01fF
C39860 NOR2X1_LOC_45/B INVX1_LOC_41/Y 0.03fF
C39861 NAND2X1_LOC_493/Y INVX1_LOC_118/A 0.00fF
C39862 INVX1_LOC_201/Y INPUT_0 0.08fF
C39863 NOR2X1_LOC_678/A NOR2X1_LOC_666/a_36_216# 0.00fF
C39864 NOR2X1_LOC_67/Y INVX1_LOC_26/Y 0.23fF
C39865 NOR2X1_LOC_334/Y INVX1_LOC_32/A 0.08fF
C39866 NOR2X1_LOC_553/B NOR2X1_LOC_565/B 0.04fF
C39867 INVX1_LOC_81/Y VDD 0.21fF
C39868 NAND2X1_LOC_74/B NOR2X1_LOC_748/A 0.36fF
C39869 INVX1_LOC_3/Y NOR2X1_LOC_825/a_36_216# 0.01fF
C39870 NOR2X1_LOC_543/a_36_216# INVX1_LOC_71/A 0.00fF
C39871 NOR2X1_LOC_78/B NOR2X1_LOC_19/B 0.57fF
C39872 NOR2X1_LOC_516/B NOR2X1_LOC_542/Y 0.15fF
C39873 NAND2X1_LOC_739/B INVX1_LOC_291/Y 0.00fF
C39874 INVX1_LOC_310/A INVX1_LOC_31/Y 0.14fF
C39875 NOR2X1_LOC_45/B NAND2X1_LOC_593/Y 0.07fF
C39876 INVX1_LOC_303/A NOR2X1_LOC_78/A 0.07fF
C39877 NAND2X1_LOC_35/Y NAND2X1_LOC_456/Y 0.02fF
C39878 INPUT_0 NAND2X1_LOC_477/A 0.10fF
C39879 INVX1_LOC_256/A NOR2X1_LOC_331/B 0.22fF
C39880 INVX1_LOC_224/Y NOR2X1_LOC_89/A 0.08fF
C39881 NOR2X1_LOC_667/Y NOR2X1_LOC_152/A 0.06fF
C39882 NOR2X1_LOC_337/Y NOR2X1_LOC_344/A 0.08fF
C39883 NAND2X1_LOC_796/a_36_24# INVX1_LOC_33/Y 0.00fF
C39884 NOR2X1_LOC_6/B INVX1_LOC_201/A 0.01fF
C39885 NOR2X1_LOC_769/A INVX1_LOC_37/A 0.01fF
C39886 NOR2X1_LOC_500/Y NOR2X1_LOC_569/a_36_216# 0.00fF
C39887 NOR2X1_LOC_15/Y NOR2X1_LOC_155/A 0.03fF
C39888 INPUT_6 NOR2X1_LOC_1/Y 0.46fF
C39889 NAND2X1_LOC_860/A INVX1_LOC_12/A 0.02fF
C39890 INVX1_LOC_50/A NOR2X1_LOC_754/A 0.01fF
C39891 NOR2X1_LOC_329/B INVX1_LOC_22/A 0.08fF
C39892 INVX1_LOC_78/A NAND2X1_LOC_72/B 0.03fF
C39893 INVX1_LOC_171/Y INVX1_LOC_294/A 0.27fF
C39894 NOR2X1_LOC_89/A NAND2X1_LOC_793/B 0.07fF
C39895 INVX1_LOC_206/Y INVX1_LOC_266/Y 0.04fF
C39896 NOR2X1_LOC_361/B NOR2X1_LOC_831/B 0.16fF
C39897 INVX1_LOC_35/A NAND2X1_LOC_291/B 0.03fF
C39898 D_INPUT_4 INVX1_LOC_22/A 0.04fF
C39899 INVX1_LOC_17/A NAND2X1_LOC_798/B 0.08fF
C39900 NAND2X1_LOC_456/a_36_24# INVX1_LOC_23/A 0.00fF
C39901 INVX1_LOC_31/A NOR2X1_LOC_54/a_36_216# 0.00fF
C39902 NOR2X1_LOC_759/Y NOR2X1_LOC_52/a_36_216# 0.00fF
C39903 NAND2X1_LOC_470/B NOR2X1_LOC_449/A 0.12fF
C39904 INVX1_LOC_128/Y NAND2X1_LOC_61/Y 0.15fF
C39905 INVX1_LOC_98/A INVX1_LOC_168/A 0.26fF
C39906 NOR2X1_LOC_655/B INVX1_LOC_48/A 0.10fF
C39907 INVX1_LOC_208/A NOR2X1_LOC_335/B 0.03fF
C39908 INVX1_LOC_249/A INVX1_LOC_46/A 0.03fF
C39909 NOR2X1_LOC_781/a_36_216# NAND2X1_LOC_654/B 0.00fF
C39910 INVX1_LOC_26/A INVX1_LOC_87/A 0.09fF
C39911 NOR2X1_LOC_646/a_36_216# NAND2X1_LOC_348/A 0.00fF
C39912 NOR2X1_LOC_322/Y NAND2X1_LOC_859/Y 0.10fF
C39913 NOR2X1_LOC_473/B INVX1_LOC_313/A 0.10fF
C39914 NOR2X1_LOC_681/Y NOR2X1_LOC_152/Y 0.04fF
C39915 NOR2X1_LOC_589/A INVX1_LOC_79/A 0.42fF
C39916 INVX1_LOC_50/Y INVX1_LOC_29/A 0.06fF
C39917 INVX1_LOC_2/A INVX1_LOC_159/Y 0.00fF
C39918 INVX1_LOC_233/A INVX1_LOC_170/Y 0.01fF
C39919 NOR2X1_LOC_152/Y INVX1_LOC_37/A 0.10fF
C39920 NOR2X1_LOC_387/Y VDD 0.26fF
C39921 NAND2X1_LOC_550/A NOR2X1_LOC_88/Y 0.07fF
C39922 INVX1_LOC_21/A INVX1_LOC_125/A 0.06fF
C39923 INVX1_LOC_83/A NOR2X1_LOC_19/B 0.60fF
C39924 INVX1_LOC_25/A NOR2X1_LOC_38/B 0.26fF
C39925 INVX1_LOC_90/A NOR2X1_LOC_246/Y 0.01fF
C39926 NOR2X1_LOC_532/Y NOR2X1_LOC_356/A 0.01fF
C39927 INVX1_LOC_57/Y INVX1_LOC_54/A 0.10fF
C39928 NOR2X1_LOC_246/Y NOR2X1_LOC_389/B 0.03fF
C39929 INVX1_LOC_212/Y VDD 0.32fF
C39930 NOR2X1_LOC_344/A VDD 0.61fF
C39931 NAND2X1_LOC_390/A NOR2X1_LOC_167/Y 0.10fF
C39932 NOR2X1_LOC_208/Y INVX1_LOC_44/A 0.01fF
C39933 INVX1_LOC_166/A NOR2X1_LOC_415/Y 0.01fF
C39934 INVX1_LOC_90/A NAND2X1_LOC_7/a_36_24# 0.00fF
C39935 NAND2X1_LOC_717/Y NOR2X1_LOC_823/Y 0.01fF
C39936 NOR2X1_LOC_848/Y NOR2X1_LOC_814/a_36_216# 0.00fF
C39937 INVX1_LOC_230/Y NAND2X1_LOC_609/a_36_24# 0.00fF
C39938 INVX1_LOC_23/A NOR2X1_LOC_685/a_36_216# 0.00fF
C39939 NOR2X1_LOC_590/A NOR2X1_LOC_841/A 0.03fF
C39940 NAND2X1_LOC_550/A INVX1_LOC_84/A 0.07fF
C39941 NOR2X1_LOC_717/B NAND2X1_LOC_496/a_36_24# 0.00fF
C39942 NAND2X1_LOC_360/B INVX1_LOC_95/Y 0.03fF
C39943 NOR2X1_LOC_514/Y VDD 0.24fF
C39944 INVX1_LOC_266/A INVX1_LOC_29/A 0.07fF
C39945 NOR2X1_LOC_512/Y INVX1_LOC_54/A 0.00fF
C39946 NOR2X1_LOC_175/A NOR2X1_LOC_35/Y 0.11fF
C39947 NOR2X1_LOC_160/B INVX1_LOC_84/A 0.14fF
C39948 NAND2X1_LOC_357/B VDD 1.59fF
C39949 INVX1_LOC_90/A NAND2X1_LOC_525/a_36_24# 0.00fF
C39950 NOR2X1_LOC_859/A NOR2X1_LOC_862/B 0.08fF
C39951 INVX1_LOC_230/Y INVX1_LOC_63/A 0.07fF
C39952 NOR2X1_LOC_589/A INVX1_LOC_91/A 0.07fF
C39953 NOR2X1_LOC_763/A NOR2X1_LOC_48/B 0.02fF
C39954 NOR2X1_LOC_441/Y NOR2X1_LOC_127/Y 0.08fF
C39955 NAND2X1_LOC_537/Y INVX1_LOC_12/A 0.14fF
C39956 NOR2X1_LOC_495/Y INVX1_LOC_118/A 0.02fF
C39957 NOR2X1_LOC_322/Y NAND2X1_LOC_807/Y 0.04fF
C39958 INVX1_LOC_278/A NOR2X1_LOC_89/Y 0.01fF
C39959 INVX1_LOC_48/A NOR2X1_LOC_99/B 0.08fF
C39960 NAND2X1_LOC_181/Y INVX1_LOC_76/A 0.07fF
C39961 NAND2X1_LOC_549/B VDD 0.01fF
C39962 NAND2X1_LOC_629/Y INVX1_LOC_117/A 0.01fF
C39963 INVX1_LOC_89/A NOR2X1_LOC_334/A 0.61fF
C39964 NOR2X1_LOC_103/Y NOR2X1_LOC_89/A 0.24fF
C39965 NOR2X1_LOC_473/B INVX1_LOC_6/A 0.26fF
C39966 INVX1_LOC_90/A NAND2X1_LOC_144/a_36_24# 0.00fF
C39967 INVX1_LOC_290/A NAND2X1_LOC_469/B 0.26fF
C39968 NOR2X1_LOC_251/Y INVX1_LOC_46/A 0.01fF
C39969 INVX1_LOC_171/A INVX1_LOC_91/A 0.03fF
C39970 NOR2X1_LOC_457/A INVX1_LOC_290/Y 0.07fF
C39971 INVX1_LOC_229/Y INVX1_LOC_11/Y 0.10fF
C39972 NAND2X1_LOC_712/A INVX1_LOC_20/A 0.01fF
C39973 NOR2X1_LOC_388/Y NAND2X1_LOC_93/B 0.07fF
C39974 INVX1_LOC_1/A NOR2X1_LOC_38/B 0.11fF
C39975 NOR2X1_LOC_389/A INVX1_LOC_114/Y 0.06fF
C39976 INVX1_LOC_17/A INVX1_LOC_47/Y 0.74fF
C39977 NOR2X1_LOC_248/Y INVX1_LOC_29/A 0.01fF
C39978 NOR2X1_LOC_322/Y INVX1_LOC_6/A 0.18fF
C39979 NOR2X1_LOC_561/Y NOR2X1_LOC_314/Y 0.04fF
C39980 NOR2X1_LOC_561/Y NOR2X1_LOC_422/Y 0.05fF
C39981 INVX1_LOC_160/Y NOR2X1_LOC_857/A 0.00fF
C39982 NOR2X1_LOC_826/Y NOR2X1_LOC_32/B 0.02fF
C39983 INVX1_LOC_45/A NOR2X1_LOC_89/A 0.07fF
C39984 NAND2X1_LOC_550/A INVX1_LOC_15/A 0.07fF
C39985 NOR2X1_LOC_711/Y INVX1_LOC_85/Y 0.01fF
C39986 INVX1_LOC_77/A NAND2X1_LOC_475/Y 0.19fF
C39987 INVX1_LOC_174/A NAND2X1_LOC_429/a_36_24# 0.01fF
C39988 NOR2X1_LOC_160/B INVX1_LOC_15/A 0.43fF
C39989 INVX1_LOC_30/A INVX1_LOC_290/Y 0.10fF
C39990 NOR2X1_LOC_772/Y INVX1_LOC_285/A 0.32fF
C39991 NOR2X1_LOC_389/A NOR2X1_LOC_467/A 0.10fF
C39992 D_INPUT_6 INVX1_LOC_296/A 0.06fF
C39993 NOR2X1_LOC_272/Y INVX1_LOC_57/A 0.10fF
C39994 INVX1_LOC_58/A NOR2X1_LOC_626/a_36_216# 0.01fF
C39995 INVX1_LOC_54/Y INVX1_LOC_92/A 0.03fF
C39996 NOR2X1_LOC_70/a_36_216# INPUT_4 0.00fF
C39997 NAND2X1_LOC_866/B NAND2X1_LOC_836/Y 0.10fF
C39998 INVX1_LOC_57/Y NOR2X1_LOC_48/B 0.04fF
C39999 NOR2X1_LOC_392/B INVX1_LOC_285/A 0.10fF
C40000 NAND2X1_LOC_861/Y INVX1_LOC_37/A 0.07fF
C40001 NOR2X1_LOC_107/Y INVX1_LOC_87/A 0.01fF
C40002 INVX1_LOC_90/A NOR2X1_LOC_562/A 0.01fF
C40003 INVX1_LOC_34/A INVX1_LOC_136/Y 0.01fF
C40004 NOR2X1_LOC_192/A NOR2X1_LOC_74/A 0.02fF
C40005 NOR2X1_LOC_78/A NOR2X1_LOC_83/a_36_216# 0.00fF
C40006 NOR2X1_LOC_568/A NOR2X1_LOC_170/A 0.01fF
C40007 NOR2X1_LOC_392/B NOR2X1_LOC_814/A 0.01fF
C40008 NAND2X1_LOC_465/Y NAND2X1_LOC_456/Y 0.07fF
C40009 NOR2X1_LOC_78/B NOR2X1_LOC_216/B 0.03fF
C40010 NOR2X1_LOC_411/Y NAND2X1_LOC_35/Y 0.05fF
C40011 INVX1_LOC_64/A NAND2X1_LOC_208/a_36_24# 0.00fF
C40012 NOR2X1_LOC_82/A INVX1_LOC_26/A 0.11fF
C40013 NAND2X1_LOC_9/Y INVX1_LOC_27/A 0.07fF
C40014 INVX1_LOC_71/A NOR2X1_LOC_89/A 0.07fF
C40015 NOR2X1_LOC_6/B NOR2X1_LOC_673/B 0.01fF
C40016 NOR2X1_LOC_702/Y VDD 0.12fF
C40017 NAND2X1_LOC_654/B NOR2X1_LOC_586/Y 0.04fF
C40018 NOR2X1_LOC_772/A INVX1_LOC_46/A 0.04fF
C40019 INVX1_LOC_135/A NOR2X1_LOC_536/A 0.02fF
C40020 INVX1_LOC_233/A INVX1_LOC_27/A 0.10fF
C40021 NAND2X1_LOC_330/a_36_24# NOR2X1_LOC_89/A 0.01fF
C40022 NAND2X1_LOC_361/Y NAND2X1_LOC_63/Y 0.04fF
C40023 INVX1_LOC_25/A NOR2X1_LOC_468/Y 0.10fF
C40024 INVX1_LOC_124/A NAND2X1_LOC_475/Y 0.10fF
C40025 NAND2X1_LOC_214/B NAND2X1_LOC_553/A 0.01fF
C40026 NOR2X1_LOC_186/Y NOR2X1_LOC_772/B 0.00fF
C40027 NAND2X1_LOC_319/A INVX1_LOC_118/A 0.01fF
C40028 INVX1_LOC_224/A INVX1_LOC_224/Y 0.14fF
C40029 NAND2X1_LOC_793/Y INVX1_LOC_181/A 0.20fF
C40030 INVX1_LOC_55/Y NAND2X1_LOC_472/Y 0.07fF
C40031 D_INPUT_1 INVX1_LOC_269/A 0.25fF
C40032 INVX1_LOC_50/A NAND2X1_LOC_787/a_36_24# 0.01fF
C40033 INVX1_LOC_224/Y INVX1_LOC_11/A 1.20fF
C40034 NAND2X1_LOC_182/A INVX1_LOC_19/A 0.03fF
C40035 INVX1_LOC_135/A NAND2X1_LOC_659/a_36_24# 0.01fF
C40036 NOR2X1_LOC_598/B NOR2X1_LOC_15/Y 0.05fF
C40037 INVX1_LOC_233/Y INVX1_LOC_234/Y 0.05fF
C40038 INVX1_LOC_104/A INVX1_LOC_19/A 0.15fF
C40039 NAND2X1_LOC_849/A VDD 0.13fF
C40040 NAND2X1_LOC_741/B NOR2X1_LOC_409/B 0.06fF
C40041 NOR2X1_LOC_423/Y INVX1_LOC_186/Y 0.00fF
C40042 NAND2X1_LOC_563/Y NAND2X1_LOC_82/Y 0.25fF
C40043 NAND2X1_LOC_553/A INVX1_LOC_27/A 0.01fF
C40044 INVX1_LOC_226/Y NOR2X1_LOC_49/a_36_216# 0.00fF
C40045 NOR2X1_LOC_596/A NOR2X1_LOC_467/A 0.07fF
C40046 INVX1_LOC_71/A NOR2X1_LOC_170/A 0.01fF
C40047 INVX1_LOC_140/A INVX1_LOC_77/Y 0.10fF
C40048 NOR2X1_LOC_6/B INVX1_LOC_29/A 4.17fF
C40049 NAND2X1_LOC_149/Y INVX1_LOC_5/A 0.12fF
C40050 NOR2X1_LOC_15/Y NAND2X1_LOC_725/A 0.05fF
C40051 INVX1_LOC_278/A NOR2X1_LOC_401/A 0.01fF
C40052 NOR2X1_LOC_490/Y NOR2X1_LOC_536/A 0.01fF
C40053 INVX1_LOC_167/Y INVX1_LOC_11/Y 0.26fF
C40054 INVX1_LOC_309/A INVX1_LOC_20/A 0.03fF
C40055 INVX1_LOC_136/A NOR2X1_LOC_471/a_36_216# 0.02fF
C40056 INVX1_LOC_208/A INVX1_LOC_84/A 0.01fF
C40057 NAND2X1_LOC_820/a_36_24# NOR2X1_LOC_649/B 0.01fF
C40058 INVX1_LOC_31/A NOR2X1_LOC_699/a_36_216# 0.15fF
C40059 NOR2X1_LOC_71/Y NAND2X1_LOC_243/Y 0.00fF
C40060 INVX1_LOC_58/A NOR2X1_LOC_331/Y 0.03fF
C40061 NAND2X1_LOC_861/Y NOR2X1_LOC_177/Y 0.04fF
C40062 NAND2X1_LOC_655/A NAND2X1_LOC_642/Y 0.15fF
C40063 NAND2X1_LOC_573/A NOR2X1_LOC_831/B 0.23fF
C40064 NAND2X1_LOC_198/B INVX1_LOC_78/A 0.05fF
C40065 NOR2X1_LOC_516/B INVX1_LOC_84/A 0.09fF
C40066 NOR2X1_LOC_222/Y INVX1_LOC_186/Y 0.07fF
C40067 NOR2X1_LOC_607/A INVX1_LOC_94/Y 0.01fF
C40068 INVX1_LOC_295/A NAND2X1_LOC_93/B 0.41fF
C40069 NOR2X1_LOC_788/B NOR2X1_LOC_640/Y 0.02fF
C40070 NOR2X1_LOC_208/A INVX1_LOC_44/A 0.16fF
C40071 NOR2X1_LOC_835/B INVX1_LOC_117/A 0.26fF
C40072 INVX1_LOC_278/A NOR2X1_LOC_160/B 0.50fF
C40073 INVX1_LOC_269/A NOR2X1_LOC_652/Y 0.37fF
C40074 INVX1_LOC_91/A INVX1_LOC_20/A 0.19fF
C40075 INVX1_LOC_24/A NOR2X1_LOC_25/Y 0.03fF
C40076 NOR2X1_LOC_186/Y INVX1_LOC_88/A 0.26fF
C40077 INVX1_LOC_303/Y INVX1_LOC_117/A 0.01fF
C40078 NOR2X1_LOC_644/B NOR2X1_LOC_678/A 0.00fF
C40079 INVX1_LOC_295/A NAND2X1_LOC_425/Y 0.19fF
C40080 NOR2X1_LOC_86/A NOR2X1_LOC_662/A 0.99fF
C40081 NOR2X1_LOC_528/Y INVX1_LOC_46/A 0.08fF
C40082 NOR2X1_LOC_718/B INVX1_LOC_32/A 0.03fF
C40083 NOR2X1_LOC_238/a_36_216# NOR2X1_LOC_693/Y -0.01fF
C40084 NOR2X1_LOC_163/Y INVX1_LOC_54/A 0.01fF
C40085 INVX1_LOC_21/A NAND2X1_LOC_538/Y 0.07fF
C40086 NOR2X1_LOC_65/B NAND2X1_LOC_198/B 0.03fF
C40087 NOR2X1_LOC_13/Y NAND2X1_LOC_61/Y 0.10fF
C40088 NAND2X1_LOC_338/B NAND2X1_LOC_254/Y 0.01fF
C40089 INVX1_LOC_13/A NAND2X1_LOC_773/B 0.11fF
C40090 INVX1_LOC_56/Y NAND2X1_LOC_81/B 0.03fF
C40091 INVX1_LOC_135/A NOR2X1_LOC_649/B 0.10fF
C40092 NAND2X1_LOC_364/A INVX1_LOC_57/A 0.11fF
C40093 NOR2X1_LOC_614/Y INVX1_LOC_69/A 0.00fF
C40094 NOR2X1_LOC_618/a_36_216# NAND2X1_LOC_74/B 0.00fF
C40095 INVX1_LOC_6/A INVX1_LOC_281/Y 0.01fF
C40096 INVX1_LOC_11/Y INVX1_LOC_20/A 8.49fF
C40097 INVX1_LOC_135/A INVX1_LOC_3/A 0.57fF
C40098 NOR2X1_LOC_828/A NAND2X1_LOC_438/a_36_24# 0.00fF
C40099 NOR2X1_LOC_643/A NAND2X1_LOC_473/A 0.02fF
C40100 INVX1_LOC_24/A NAND2X1_LOC_299/a_36_24# 0.00fF
C40101 NAND2X1_LOC_112/Y INVX1_LOC_272/A 0.03fF
C40102 NOR2X1_LOC_468/Y INVX1_LOC_1/A 0.10fF
C40103 INVX1_LOC_24/A NOR2X1_LOC_646/B 0.00fF
C40104 INVX1_LOC_135/A NOR2X1_LOC_661/A 0.07fF
C40105 NOR2X1_LOC_457/B INVX1_LOC_23/A 0.19fF
C40106 INVX1_LOC_90/A INVX1_LOC_285/A 0.09fF
C40107 INVX1_LOC_35/A NOR2X1_LOC_274/B 0.23fF
C40108 NOR2X1_LOC_389/B INVX1_LOC_285/A 0.10fF
C40109 INVX1_LOC_20/A NOR2X1_LOC_421/Y 0.03fF
C40110 NOR2X1_LOC_846/Y INVX1_LOC_31/A 0.24fF
C40111 NAND2X1_LOC_778/Y NOR2X1_LOC_372/A 0.14fF
C40112 INVX1_LOC_90/A NOR2X1_LOC_814/A 0.07fF
C40113 NOR2X1_LOC_391/B NOR2X1_LOC_655/Y 0.72fF
C40114 INVX1_LOC_89/A INVX1_LOC_293/Y 0.00fF
C40115 INVX1_LOC_64/A NOR2X1_LOC_703/B 0.03fF
C40116 NAND2X1_LOC_350/B INVX1_LOC_15/A 0.09fF
C40117 NOR2X1_LOC_456/a_36_216# NOR2X1_LOC_794/B 0.00fF
C40118 NAND2X1_LOC_170/A NOR2X1_LOC_48/B 0.03fF
C40119 NOR2X1_LOC_91/A NAND2X1_LOC_833/Y 0.09fF
C40120 NOR2X1_LOC_314/Y INVX1_LOC_76/A 0.04fF
C40121 NOR2X1_LOC_389/B NOR2X1_LOC_814/A 0.07fF
C40122 INVX1_LOC_50/A INVX1_LOC_49/A 0.55fF
C40123 INVX1_LOC_11/Y NOR2X1_LOC_765/Y 0.01fF
C40124 INVX1_LOC_13/Y INVX1_LOC_170/A 0.01fF
C40125 INVX1_LOC_234/A NOR2X1_LOC_671/Y 0.03fF
C40126 NOR2X1_LOC_500/A INVX1_LOC_53/A 0.08fF
C40127 INVX1_LOC_208/A INVX1_LOC_15/A 0.01fF
C40128 INVX1_LOC_149/A INVX1_LOC_87/A 0.02fF
C40129 NOR2X1_LOC_303/Y INVX1_LOC_53/A 0.10fF
C40130 NOR2X1_LOC_598/B NOR2X1_LOC_860/B 0.07fF
C40131 INVX1_LOC_224/A NOR2X1_LOC_103/Y 0.07fF
C40132 NOR2X1_LOC_142/Y NOR2X1_LOC_383/B 0.17fF
C40133 NOR2X1_LOC_516/B INVX1_LOC_15/A 0.16fF
C40134 INVX1_LOC_35/A NAND2X1_LOC_218/B 0.01fF
C40135 INVX1_LOC_11/A NOR2X1_LOC_103/Y 0.07fF
C40136 NAND2X1_LOC_190/Y NOR2X1_LOC_794/B 0.04fF
C40137 INVX1_LOC_89/A NAND2X1_LOC_74/B 2.67fF
C40138 NOR2X1_LOC_389/A INVX1_LOC_1/A 0.29fF
C40139 INVX1_LOC_285/Y NOR2X1_LOC_831/B 0.00fF
C40140 NOR2X1_LOC_15/Y NOR2X1_LOC_372/A 0.00fF
C40141 INVX1_LOC_76/A INVX1_LOC_117/A 0.55fF
C40142 INVX1_LOC_21/A NOR2X1_LOC_602/a_36_216# 0.00fF
C40143 NAND2X1_LOC_9/Y NAND2X1_LOC_99/Y 0.01fF
C40144 NOR2X1_LOC_45/B INVX1_LOC_185/A 0.03fF
C40145 INVX1_LOC_11/A NOR2X1_LOC_541/Y 0.07fF
C40146 NOR2X1_LOC_361/B NAND2X1_LOC_352/B 0.17fF
C40147 INPUT_0 NAND2X1_LOC_574/A 0.02fF
C40148 INVX1_LOC_62/A NOR2X1_LOC_67/Y 0.02fF
C40149 INVX1_LOC_88/A NOR2X1_LOC_45/Y 0.00fF
C40150 NAND2X1_LOC_363/B INVX1_LOC_77/A 0.10fF
C40151 NOR2X1_LOC_454/Y INVX1_LOC_30/A 0.07fF
C40152 NAND2X1_LOC_348/A NOR2X1_LOC_814/A 0.07fF
C40153 INVX1_LOC_222/Y INVX1_LOC_18/A 0.01fF
C40154 INVX1_LOC_35/A NOR2X1_LOC_577/Y 2.53fF
C40155 NAND2X1_LOC_733/Y NAND2X1_LOC_537/Y 0.20fF
C40156 INVX1_LOC_294/Y INVX1_LOC_29/Y 0.36fF
C40157 INVX1_LOC_35/A NOR2X1_LOC_379/Y 0.04fF
C40158 INVX1_LOC_25/A NOR2X1_LOC_295/Y 0.01fF
C40159 INVX1_LOC_34/Y NAND2X1_LOC_99/A 0.01fF
C40160 INVX1_LOC_9/Y NOR2X1_LOC_334/Y 0.01fF
C40161 INVX1_LOC_77/A NOR2X1_LOC_640/a_36_216# 0.00fF
C40162 INVX1_LOC_224/Y NOR2X1_LOC_52/B 0.04fF
C40163 NOR2X1_LOC_391/B NOR2X1_LOC_649/B 0.01fF
C40164 NOR2X1_LOC_32/B NOR2X1_LOC_690/A 0.01fF
C40165 INVX1_LOC_205/Y INVX1_LOC_205/A 0.01fF
C40166 INVX1_LOC_53/Y INVX1_LOC_78/A 0.03fF
C40167 NAND2X1_LOC_785/A INVX1_LOC_57/A 0.07fF
C40168 NAND2X1_LOC_624/a_36_24# INVX1_LOC_255/A 0.00fF
C40169 NOR2X1_LOC_220/A INVX1_LOC_116/Y 0.20fF
C40170 NAND2X1_LOC_555/a_36_24# NOR2X1_LOC_249/Y 0.00fF
C40171 NOR2X1_LOC_32/B NOR2X1_LOC_413/Y 0.02fF
C40172 INVX1_LOC_2/A INVX1_LOC_50/A 1.13fF
C40173 NOR2X1_LOC_655/B NOR2X1_LOC_383/B 0.02fF
C40174 NOR2X1_LOC_667/A NAND2X1_LOC_285/a_36_24# 0.01fF
C40175 NOR2X1_LOC_705/B NOR2X1_LOC_590/A 0.03fF
C40176 NAND2X1_LOC_35/Y INVX1_LOC_34/A 0.07fF
C40177 NOR2X1_LOC_226/A INVX1_LOC_50/A 0.03fF
C40178 INVX1_LOC_45/A INVX1_LOC_11/A 0.22fF
C40179 INVX1_LOC_102/Y NOR2X1_LOC_89/A 0.07fF
C40180 NOR2X1_LOC_52/B NAND2X1_LOC_793/B 0.18fF
C40181 NAND2X1_LOC_11/Y INVX1_LOC_57/A 0.08fF
C40182 INVX1_LOC_11/A NOR2X1_LOC_568/A 0.03fF
C40183 NOR2X1_LOC_813/Y NOR2X1_LOC_536/A 0.04fF
C40184 NAND2X1_LOC_579/A NOR2X1_LOC_522/Y 0.11fF
C40185 INVX1_LOC_246/Y NOR2X1_LOC_92/Y 0.01fF
C40186 NOR2X1_LOC_790/B INVX1_LOC_177/A 0.01fF
C40187 INVX1_LOC_10/A NAND2X1_LOC_454/Y 0.02fF
C40188 NOR2X1_LOC_152/A NOR2X1_LOC_536/A 0.29fF
C40189 NOR2X1_LOC_772/B INVX1_LOC_225/A 0.14fF
C40190 NOR2X1_LOC_65/B INVX1_LOC_53/Y 0.01fF
C40191 NAND2X1_LOC_656/A NAND2X1_LOC_216/a_36_24# 0.01fF
C40192 INVX1_LOC_1/A NOR2X1_LOC_596/A 0.08fF
C40193 INVX1_LOC_206/Y INVX1_LOC_19/A 0.03fF
C40194 NAND2X1_LOC_53/Y NOR2X1_LOC_68/A 0.07fF
C40195 D_INPUT_1 NAND2X1_LOC_563/A 0.10fF
C40196 NOR2X1_LOC_381/Y INVX1_LOC_228/A 0.03fF
C40197 NAND2X1_LOC_802/A NOR2X1_LOC_92/Y 0.05fF
C40198 NOR2X1_LOC_236/a_36_216# INVX1_LOC_26/A 0.00fF
C40199 NOR2X1_LOC_536/A INVX1_LOC_280/A 0.08fF
C40200 INVX1_LOC_177/Y INVX1_LOC_161/Y 0.04fF
C40201 NOR2X1_LOC_681/Y INVX1_LOC_291/A 0.01fF
C40202 INVX1_LOC_157/A NOR2X1_LOC_449/A 0.02fF
C40203 INVX1_LOC_37/A INVX1_LOC_291/A 0.07fF
C40204 INVX1_LOC_269/A D_INPUT_2 0.07fF
C40205 INVX1_LOC_139/Y NAND2X1_LOC_93/B 0.03fF
C40206 INVX1_LOC_295/A NAND2X1_LOC_470/B 0.03fF
C40207 NAND2X1_LOC_740/Y NAND2X1_LOC_812/a_36_24# 0.00fF
C40208 NOR2X1_LOC_598/B INVX1_LOC_226/A 0.02fF
C40209 INVX1_LOC_34/A NAND2X1_LOC_571/Y 0.19fF
C40210 NAND2X1_LOC_573/a_36_24# NOR2X1_LOC_361/B 0.01fF
C40211 NOR2X1_LOC_216/B INVX1_LOC_46/A 0.01fF
C40212 INVX1_LOC_35/A NOR2X1_LOC_175/B 0.16fF
C40213 NOR2X1_LOC_86/A INVX1_LOC_57/A 0.03fF
C40214 NOR2X1_LOC_91/A INVX1_LOC_273/Y 0.01fF
C40215 NOR2X1_LOC_65/B INVX1_LOC_145/Y 0.01fF
C40216 INVX1_LOC_136/A NAND2X1_LOC_711/Y 0.03fF
C40217 NOR2X1_LOC_373/Y NOR2X1_LOC_693/Y 0.05fF
C40218 INVX1_LOC_292/A NOR2X1_LOC_360/Y 0.01fF
C40219 INVX1_LOC_50/A NAND2X1_LOC_664/a_36_24# 0.00fF
C40220 INVX1_LOC_11/A INVX1_LOC_71/A 13.15fF
C40221 NAND2X1_LOC_477/Y NOR2X1_LOC_368/Y 0.07fF
C40222 INVX1_LOC_108/Y NOR2X1_LOC_516/B 0.00fF
C40223 INVX1_LOC_99/Y NOR2X1_LOC_78/B 0.01fF
C40224 NOR2X1_LOC_78/A INVX1_LOC_272/A 0.03fF
C40225 NAND2X1_LOC_149/Y NOR2X1_LOC_377/Y 0.03fF
C40226 NAND2X1_LOC_571/B NAND2X1_LOC_735/B 0.00fF
C40227 NAND2X1_LOC_9/Y INVX1_LOC_137/A 0.01fF
C40228 INVX1_LOC_58/A NOR2X1_LOC_561/Y 0.14fF
C40229 NAND2X1_LOC_725/B NAND2X1_LOC_736/B 0.07fF
C40230 NOR2X1_LOC_91/A NOR2X1_LOC_76/A 0.07fF
C40231 INVX1_LOC_35/A INVX1_LOC_22/A 0.12fF
C40232 NOR2X1_LOC_818/a_36_216# NOR2X1_LOC_516/B 0.02fF
C40233 INVX1_LOC_2/A NOR2X1_LOC_206/a_36_216# 0.00fF
C40234 NOR2X1_LOC_381/Y INVX1_LOC_8/A 0.01fF
C40235 INVX1_LOC_203/A INVX1_LOC_20/A 0.03fF
C40236 NOR2X1_LOC_15/Y NAND2X1_LOC_308/Y 0.08fF
C40237 NOR2X1_LOC_689/Y NOR2X1_LOC_576/B 0.22fF
C40238 NOR2X1_LOC_598/B NOR2X1_LOC_97/B 0.06fF
C40239 NOR2X1_LOC_722/Y NOR2X1_LOC_723/a_36_216# 0.00fF
C40240 NOR2X1_LOC_364/A INVX1_LOC_38/A 0.22fF
C40241 NAND2X1_LOC_803/B NOR2X1_LOC_172/Y 0.34fF
C40242 INVX1_LOC_225/A INVX1_LOC_88/A 0.00fF
C40243 NAND2X1_LOC_477/Y INVX1_LOC_46/A 0.12fF
C40244 NOR2X1_LOC_593/Y NOR2X1_LOC_541/Y 0.04fF
C40245 NOR2X1_LOC_71/Y NAND2X1_LOC_205/A 0.04fF
C40246 NOR2X1_LOC_285/A INVX1_LOC_89/A 0.06fF
C40247 NOR2X1_LOC_791/A NOR2X1_LOC_791/B 0.00fF
C40248 INVX1_LOC_5/A INVX1_LOC_16/A 0.14fF
C40249 INVX1_LOC_256/A NOR2X1_LOC_388/Y 0.10fF
C40250 INVX1_LOC_135/A NOR2X1_LOC_476/B 0.01fF
C40251 NOR2X1_LOC_361/B NAND2X1_LOC_357/B 0.47fF
C40252 NOR2X1_LOC_220/B NOR2X1_LOC_211/A 0.04fF
C40253 NOR2X1_LOC_76/A INVX1_LOC_23/A 0.29fF
C40254 NAND2X1_LOC_778/a_36_24# NAND2X1_LOC_374/Y 0.00fF
C40255 NOR2X1_LOC_813/Y INVX1_LOC_3/A 0.07fF
C40256 INVX1_LOC_179/A INVX1_LOC_54/A 0.01fF
C40257 NOR2X1_LOC_2/Y NOR2X1_LOC_36/A 0.61fF
C40258 NOR2X1_LOC_180/B INVX1_LOC_23/A 0.07fF
C40259 NOR2X1_LOC_219/Y NOR2X1_LOC_215/A 0.10fF
C40260 INVX1_LOC_259/Y INVX1_LOC_89/A 0.01fF
C40261 NAND2X1_LOC_833/Y INVX1_LOC_31/A 0.01fF
C40262 INVX1_LOC_77/A INVX1_LOC_30/A 0.45fF
C40263 INVX1_LOC_161/Y INVX1_LOC_104/A 0.08fF
C40264 NAND2X1_LOC_656/A INVX1_LOC_18/A 0.73fF
C40265 INVX1_LOC_45/A NOR2X1_LOC_433/A 3.22fF
C40266 NOR2X1_LOC_92/Y NAND2X1_LOC_334/a_36_24# 0.01fF
C40267 INVX1_LOC_182/A NOR2X1_LOC_383/B 0.18fF
C40268 INVX1_LOC_178/A INVX1_LOC_16/A 0.10fF
C40269 INVX1_LOC_314/Y INVX1_LOC_72/A 0.08fF
C40270 INVX1_LOC_132/A NOR2X1_LOC_500/B 0.10fF
C40271 INVX1_LOC_89/A NOR2X1_LOC_660/Y 0.03fF
C40272 NOR2X1_LOC_220/A INVX1_LOC_1/A 0.10fF
C40273 NAND2X1_LOC_763/B INVX1_LOC_77/A 0.01fF
C40274 INVX1_LOC_214/Y NAND2X1_LOC_537/Y 0.00fF
C40275 INVX1_LOC_280/A INVX1_LOC_3/A 0.82fF
C40276 INVX1_LOC_93/A NAND2X1_LOC_392/Y 0.03fF
C40277 NOR2X1_LOC_321/Y NOR2X1_LOC_321/a_36_216# 0.00fF
C40278 NOR2X1_LOC_553/a_36_216# INVX1_LOC_104/A 0.00fF
C40279 INVX1_LOC_91/A INVX1_LOC_4/A 0.12fF
C40280 NAND2X1_LOC_465/A INVX1_LOC_42/A 0.00fF
C40281 NOR2X1_LOC_590/A NOR2X1_LOC_392/B 0.03fF
C40282 INVX1_LOC_38/A NOR2X1_LOC_814/A 0.07fF
C40283 NOR2X1_LOC_667/A NAND2X1_LOC_538/Y 0.04fF
C40284 INVX1_LOC_45/A NOR2X1_LOC_593/Y 0.02fF
C40285 NOR2X1_LOC_754/a_36_216# NOR2X1_LOC_693/Y 0.00fF
C40286 INVX1_LOC_14/A INVX1_LOC_43/A 0.04fF
C40287 INVX1_LOC_2/A NAND2X1_LOC_227/Y 0.44fF
C40288 NOR2X1_LOC_593/Y NOR2X1_LOC_568/A 0.02fF
C40289 NAND2X1_LOC_475/Y INVX1_LOC_9/A 0.10fF
C40290 NAND2X1_LOC_198/B NOR2X1_LOC_152/Y 0.10fF
C40291 NOR2X1_LOC_65/B NOR2X1_LOC_113/B 0.01fF
C40292 NAND2X1_LOC_9/Y NOR2X1_LOC_19/B 0.08fF
C40293 NOR2X1_LOC_226/A NAND2X1_LOC_227/Y 0.19fF
C40294 INVX1_LOC_73/A INVX1_LOC_23/A 0.07fF
C40295 NOR2X1_LOC_60/Y INVX1_LOC_272/A 0.03fF
C40296 INVX1_LOC_45/A NOR2X1_LOC_52/B 0.10fF
C40297 INVX1_LOC_76/A INVX1_LOC_3/Y 0.17fF
C40298 NOR2X1_LOC_456/Y INVX1_LOC_75/A 0.07fF
C40299 NOR2X1_LOC_259/B NAND2X1_LOC_257/a_36_24# 0.02fF
C40300 INVX1_LOC_30/A NAND2X1_LOC_650/a_36_24# 0.00fF
C40301 NOR2X1_LOC_74/A INVX1_LOC_29/Y 0.26fF
C40302 NOR2X1_LOC_220/A NOR2X1_LOC_794/B 0.01fF
C40303 NOR2X1_LOC_75/Y NAND2X1_LOC_841/A 0.19fF
C40304 INVX1_LOC_21/A NOR2X1_LOC_106/A 0.03fF
C40305 NOR2X1_LOC_433/A INVX1_LOC_71/A 0.19fF
C40306 INVX1_LOC_124/A INVX1_LOC_30/A 0.15fF
C40307 NAND2X1_LOC_552/A INVX1_LOC_28/A 0.03fF
C40308 INVX1_LOC_20/A INVX1_LOC_231/A 0.00fF
C40309 NAND2X1_LOC_784/A NAND2X1_LOC_858/B 0.40fF
C40310 NAND2X1_LOC_211/Y INVX1_LOC_15/A 0.07fF
C40311 INVX1_LOC_255/Y NOR2X1_LOC_817/Y 0.03fF
C40312 INVX1_LOC_58/A NOR2X1_LOC_167/Y 0.03fF
C40313 NOR2X1_LOC_593/Y INVX1_LOC_71/A 0.02fF
C40314 NOR2X1_LOC_9/Y INVX1_LOC_29/Y 0.01fF
C40315 NOR2X1_LOC_75/Y INVX1_LOC_268/A 0.16fF
C40316 INVX1_LOC_132/A INVX1_LOC_303/A 0.02fF
C40317 INVX1_LOC_256/A NAND2X1_LOC_479/Y 0.03fF
C40318 NAND2X1_LOC_311/a_36_24# NOR2X1_LOC_168/B 0.00fF
C40319 NOR2X1_LOC_816/A INVX1_LOC_16/A 0.03fF
C40320 NOR2X1_LOC_89/A NOR2X1_LOC_331/B 0.07fF
C40321 INVX1_LOC_2/A NOR2X1_LOC_659/a_36_216# 0.00fF
C40322 INVX1_LOC_18/A NOR2X1_LOC_423/Y 0.53fF
C40323 NAND2X1_LOC_123/Y NOR2X1_LOC_674/Y 0.30fF
C40324 INVX1_LOC_27/A NAND2X1_LOC_842/B 0.38fF
C40325 NAND2X1_LOC_472/Y INVX1_LOC_32/A 0.07fF
C40326 INVX1_LOC_178/A INVX1_LOC_28/A 0.22fF
C40327 INVX1_LOC_40/Y INVX1_LOC_40/A 0.09fF
C40328 INVX1_LOC_254/Y NOR2X1_LOC_264/Y 0.25fF
C40329 INVX1_LOC_26/A INVX1_LOC_59/Y 0.05fF
C40330 NOR2X1_LOC_471/Y NOR2X1_LOC_424/a_36_216# 0.00fF
C40331 NOR2X1_LOC_52/B INVX1_LOC_71/A 0.27fF
C40332 NOR2X1_LOC_624/A NAND2X1_LOC_361/Y 0.08fF
C40333 INVX1_LOC_64/A INVX1_LOC_309/A 0.03fF
C40334 NOR2X1_LOC_222/Y INVX1_LOC_18/A 0.07fF
C40335 INVX1_LOC_11/A NOR2X1_LOC_123/B 0.07fF
C40336 INVX1_LOC_24/A INVX1_LOC_236/A 0.04fF
C40337 NAND2X1_LOC_330/a_36_24# NOR2X1_LOC_52/B 0.00fF
C40338 NOR2X1_LOC_405/A INVX1_LOC_57/A 0.12fF
C40339 NOR2X1_LOC_785/Y NOR2X1_LOC_785/A 0.27fF
C40340 NOR2X1_LOC_286/Y INVX1_LOC_132/Y 0.19fF
C40341 INVX1_LOC_108/Y INVX1_LOC_315/Y 0.01fF
C40342 NOR2X1_LOC_840/Y NOR2X1_LOC_833/Y 0.13fF
C40343 NOR2X1_LOC_45/B NOR2X1_LOC_754/Y 0.01fF
C40344 NOR2X1_LOC_862/B INVX1_LOC_69/A 0.46fF
C40345 INVX1_LOC_233/A NOR2X1_LOC_528/Y 0.10fF
C40346 INVX1_LOC_78/A INVX1_LOC_77/Y 0.02fF
C40347 INVX1_LOC_14/A NOR2X1_LOC_756/Y 0.11fF
C40348 NOR2X1_LOC_68/A NOR2X1_LOC_500/Y 0.03fF
C40349 INVX1_LOC_207/A INVX1_LOC_240/A 0.04fF
C40350 INVX1_LOC_235/Y NAND2X1_LOC_463/B -0.01fF
C40351 INVX1_LOC_314/Y NOR2X1_LOC_537/Y 0.07fF
C40352 NOR2X1_LOC_500/A NOR2X1_LOC_78/B 0.03fF
C40353 INVX1_LOC_226/Y NOR2X1_LOC_68/A 0.03fF
C40354 INVX1_LOC_2/A INVX1_LOC_105/A 0.01fF
C40355 INVX1_LOC_188/A NOR2X1_LOC_717/B 0.00fF
C40356 NOR2X1_LOC_121/Y NOR2X1_LOC_124/B 0.14fF
C40357 NOR2X1_LOC_352/a_36_216# NOR2X1_LOC_678/A 0.00fF
C40358 VDD NOR2X1_LOC_282/Y 0.18fF
C40359 INVX1_LOC_64/A INVX1_LOC_91/A 0.25fF
C40360 NAND2X1_LOC_803/B INVX1_LOC_90/A 0.11fF
C40361 INVX1_LOC_34/A NOR2X1_LOC_234/Y 0.00fF
C40362 NOR2X1_LOC_790/B INVX1_LOC_65/A 0.10fF
C40363 NOR2X1_LOC_78/B NOR2X1_LOC_303/Y 0.12fF
C40364 NOR2X1_LOC_325/A NOR2X1_LOC_325/Y 0.18fF
C40365 NOR2X1_LOC_6/B INVX1_LOC_8/A 0.12fF
C40366 NAND2X1_LOC_222/A VDD -0.00fF
C40367 NAND2X1_LOC_489/Y NAND2X1_LOC_773/B 0.01fF
C40368 NOR2X1_LOC_590/A INVX1_LOC_97/A 0.05fF
C40369 INVX1_LOC_33/Y NOR2X1_LOC_301/A 0.00fF
C40370 NOR2X1_LOC_305/Y NOR2X1_LOC_654/A 0.10fF
C40371 INVX1_LOC_177/A NOR2X1_LOC_344/A 0.02fF
C40372 NOR2X1_LOC_443/Y VDD 0.36fF
C40373 INVX1_LOC_57/A NOR2X1_LOC_857/A 0.07fF
C40374 INVX1_LOC_58/A INVX1_LOC_76/A 0.34fF
C40375 INVX1_LOC_33/A NAND2X1_LOC_342/Y 0.22fF
C40376 NOR2X1_LOC_590/A INVX1_LOC_90/A 0.16fF
C40377 NOR2X1_LOC_446/a_36_216# NOR2X1_LOC_644/A 0.00fF
C40378 NOR2X1_LOC_536/A NAND2X1_LOC_437/a_36_24# 0.00fF
C40379 INVX1_LOC_64/A INVX1_LOC_11/Y 0.06fF
C40380 NOR2X1_LOC_816/A INVX1_LOC_28/A 0.17fF
C40381 NOR2X1_LOC_455/a_36_216# INVX1_LOC_266/Y 0.01fF
C40382 INVX1_LOC_268/A NAND2X1_LOC_162/B 0.01fF
C40383 INVX1_LOC_61/Y INPUT_1 0.16fF
C40384 NAND2X1_LOC_860/A NOR2X1_LOC_9/a_36_216# 0.00fF
C40385 INVX1_LOC_22/Y INVX1_LOC_90/A 0.00fF
C40386 INVX1_LOC_13/A INVX1_LOC_24/A 0.14fF
C40387 NOR2X1_LOC_68/A INVX1_LOC_10/A 0.07fF
C40388 NOR2X1_LOC_78/B NOR2X1_LOC_254/Y 0.06fF
C40389 INVX1_LOC_13/Y NAND2X1_LOC_642/Y 0.07fF
C40390 D_INPUT_0 NOR2X1_LOC_791/B 0.00fF
C40391 NOR2X1_LOC_619/a_36_216# INVX1_LOC_176/A 0.01fF
C40392 INVX1_LOC_36/A NOR2X1_LOC_473/B 0.99fF
C40393 INVX1_LOC_136/A INVX1_LOC_89/A 2.84fF
C40394 D_INPUT_1 INVX1_LOC_12/Y 0.10fF
C40395 NOR2X1_LOC_207/A INVX1_LOC_266/Y 0.01fF
C40396 NAND2X1_LOC_549/Y VDD 0.00fF
C40397 NAND2X1_LOC_733/Y NAND2X1_LOC_855/Y 0.02fF
C40398 NAND2X1_LOC_584/a_36_24# NAND2X1_LOC_451/Y 0.00fF
C40399 NAND2X1_LOC_573/a_36_24# NAND2X1_LOC_573/A 0.01fF
C40400 INVX1_LOC_5/A NOR2X1_LOC_35/Y 0.05fF
C40401 INVX1_LOC_90/A NAND2X1_LOC_589/a_36_24# 0.00fF
C40402 NAND2X1_LOC_454/Y INVX1_LOC_307/A 0.03fF
C40403 INVX1_LOC_98/A NOR2X1_LOC_271/B 0.01fF
C40404 NAND2X1_LOC_736/B INVX1_LOC_241/A 0.00fF
C40405 INVX1_LOC_27/A NOR2X1_LOC_545/B 0.03fF
C40406 NOR2X1_LOC_278/Y INVX1_LOC_70/A 0.02fF
C40407 INVX1_LOC_290/A INVX1_LOC_63/Y 0.10fF
C40408 VDD INVX1_LOC_213/A 0.60fF
C40409 NAND2X1_LOC_833/Y NAND2X1_LOC_859/Y 0.00fF
C40410 INVX1_LOC_32/A NAND2X1_LOC_206/Y 0.03fF
C40411 NOR2X1_LOC_395/Y INVX1_LOC_241/Y 0.10fF
C40412 INVX1_LOC_50/A INVX1_LOC_118/A 0.13fF
C40413 INVX1_LOC_30/Y INVX1_LOC_8/A 0.03fF
C40414 NOR2X1_LOC_329/B INVX1_LOC_18/A 0.07fF
C40415 VDD NOR2X1_LOC_291/Y 0.45fF
C40416 INVX1_LOC_103/A NOR2X1_LOC_269/Y 0.00fF
C40417 INVX1_LOC_55/Y INVX1_LOC_24/A 0.03fF
C40418 INVX1_LOC_93/A INVX1_LOC_46/A 0.07fF
C40419 INVX1_LOC_32/A NAND2X1_LOC_773/B 0.01fF
C40420 INVX1_LOC_83/A NOR2X1_LOC_708/B 0.16fF
C40421 D_INPUT_4 INVX1_LOC_18/A 0.03fF
C40422 NAND2X1_LOC_736/B NOR2X1_LOC_298/Y 0.05fF
C40423 INVX1_LOC_227/A NOR2X1_LOC_392/B 0.00fF
C40424 NOR2X1_LOC_619/A NOR2X1_LOC_721/A 0.02fF
C40425 NOR2X1_LOC_298/Y GATE_811 0.02fF
C40426 INVX1_LOC_12/Y NOR2X1_LOC_652/Y 0.10fF
C40427 INVX1_LOC_150/Y NOR2X1_LOC_78/A 0.08fF
C40428 NAND2X1_LOC_357/B NAND2X1_LOC_573/A 0.10fF
C40429 NAND2X1_LOC_363/B INVX1_LOC_9/A 0.14fF
C40430 NAND2X1_LOC_714/B NAND2X1_LOC_453/A 0.17fF
C40431 NAND2X1_LOC_223/A NOR2X1_LOC_814/A 0.10fF
C40432 NAND2X1_LOC_528/a_36_24# INVX1_LOC_226/A 0.00fF
C40433 INVX1_LOC_43/Y INVX1_LOC_91/A 0.01fF
C40434 NOR2X1_LOC_637/Y NOR2X1_LOC_329/B 0.03fF
C40435 NOR2X1_LOC_679/B NAND2X1_LOC_648/A 0.01fF
C40436 INVX1_LOC_47/A NOR2X1_LOC_716/B 0.02fF
C40437 INVX1_LOC_226/Y NOR2X1_LOC_520/a_36_216# 0.00fF
C40438 D_INPUT_0 NOR2X1_LOC_124/B 0.22fF
C40439 NOR2X1_LOC_653/Y NOR2X1_LOC_281/a_36_216# 0.01fF
C40440 NAND2X1_LOC_833/Y NAND2X1_LOC_866/B 0.04fF
C40441 NOR2X1_LOC_273/Y INVX1_LOC_75/A 0.03fF
C40442 NOR2X1_LOC_773/Y INVX1_LOC_16/A 0.07fF
C40443 NAND2X1_LOC_347/B VDD 0.40fF
C40444 INVX1_LOC_75/A NOR2X1_LOC_759/Y 0.03fF
C40445 NOR2X1_LOC_274/a_36_216# INVX1_LOC_75/A 0.00fF
C40446 NOR2X1_LOC_52/B NOR2X1_LOC_123/B 0.07fF
C40447 NOR2X1_LOC_644/A NOR2X1_LOC_570/B 0.03fF
C40448 INVX1_LOC_202/A INVX1_LOC_75/A 0.10fF
C40449 D_INPUT_0 NOR2X1_LOC_802/A 0.07fF
C40450 INVX1_LOC_13/Y NOR2X1_LOC_271/Y 0.03fF
C40451 INVX1_LOC_62/Y NOR2X1_LOC_188/A 0.12fF
C40452 NOR2X1_LOC_433/A INVX1_LOC_102/Y 0.08fF
C40453 NOR2X1_LOC_570/Y NOR2X1_LOC_500/Y 0.03fF
C40454 NOR2X1_LOC_230/Y NOR2X1_LOC_45/B 0.20fF
C40455 NOR2X1_LOC_585/a_36_216# INVX1_LOC_91/A 0.00fF
C40456 INVX1_LOC_24/A NOR2X1_LOC_320/Y 0.04fF
C40457 INVX1_LOC_124/Y NOR2X1_LOC_192/A 0.06fF
C40458 NOR2X1_LOC_237/Y NOR2X1_LOC_322/Y 0.03fF
C40459 NAND2X1_LOC_9/Y NOR2X1_LOC_216/B 0.03fF
C40460 INVX1_LOC_62/Y NOR2X1_LOC_548/B 0.03fF
C40461 INVX1_LOC_75/A NOR2X1_LOC_550/B 0.06fF
C40462 INVX1_LOC_233/A NOR2X1_LOC_216/B 0.10fF
C40463 INVX1_LOC_12/A NAND2X1_LOC_454/Y 0.14fF
C40464 INVX1_LOC_215/Y INVX1_LOC_76/A 0.10fF
C40465 NOR2X1_LOC_19/B NOR2X1_LOC_140/a_36_216# 0.00fF
C40466 NOR2X1_LOC_68/A NOR2X1_LOC_340/a_36_216# 0.00fF
C40467 NOR2X1_LOC_745/Y VDD 0.12fF
C40468 INVX1_LOC_33/A INVX1_LOC_67/Y 0.00fF
C40469 INVX1_LOC_17/A INVX1_LOC_33/Y 0.03fF
C40470 NAND2X1_LOC_116/a_36_24# NOR2X1_LOC_199/B 0.00fF
C40471 INVX1_LOC_32/A NOR2X1_LOC_297/A 0.15fF
C40472 INVX1_LOC_183/Y NAND2X1_LOC_850/Y 0.01fF
C40473 INVX1_LOC_72/A NOR2X1_LOC_657/B 0.30fF
C40474 NOR2X1_LOC_778/B INVX1_LOC_313/Y 0.11fF
C40475 INVX1_LOC_310/A INVX1_LOC_148/A 0.00fF
C40476 NAND2X1_LOC_337/a_36_24# INVX1_LOC_46/A 0.00fF
C40477 NOR2X1_LOC_646/A D_INPUT_0 0.03fF
C40478 INVX1_LOC_36/A NAND2X1_LOC_602/a_36_24# 0.00fF
C40479 NAND2X1_LOC_66/a_36_24# INVX1_LOC_90/A 0.00fF
C40480 NAND2X1_LOC_215/a_36_24# NAND2X1_LOC_215/A 0.01fF
C40481 INVX1_LOC_50/A NAND2X1_LOC_63/Y 0.03fF
C40482 INVX1_LOC_230/Y NAND2X1_LOC_721/A 0.01fF
C40483 INVX1_LOC_2/A NAND2X1_LOC_652/Y 0.02fF
C40484 INVX1_LOC_238/Y VDD 0.17fF
C40485 NAND2X1_LOC_807/B NAND2X1_LOC_288/B 0.05fF
C40486 NOR2X1_LOC_208/Y NOR2X1_LOC_562/B 0.00fF
C40487 NOR2X1_LOC_220/a_36_216# NOR2X1_LOC_405/A 0.01fF
C40488 NOR2X1_LOC_150/a_36_216# INVX1_LOC_53/Y 0.00fF
C40489 NOR2X1_LOC_488/Y INVX1_LOC_90/A 0.65fF
C40490 INVX1_LOC_13/A NOR2X1_LOC_130/A 0.00fF
C40491 INVX1_LOC_11/A NOR2X1_LOC_331/B 0.14fF
C40492 NOR2X1_LOC_226/A NAND2X1_LOC_652/Y 0.02fF
C40493 NOR2X1_LOC_773/Y INVX1_LOC_28/A 0.16fF
C40494 INVX1_LOC_90/A NOR2X1_LOC_82/Y 0.09fF
C40495 INVX1_LOC_64/A INVX1_LOC_203/A 0.03fF
C40496 NAND2X1_LOC_803/B INVX1_LOC_38/A 0.02fF
C40497 NOR2X1_LOC_256/a_36_216# NOR2X1_LOC_124/A 0.00fF
C40498 NOR2X1_LOC_439/a_36_216# INVX1_LOC_313/Y 0.00fF
C40499 NOR2X1_LOC_707/B VDD -0.00fF
C40500 INVX1_LOC_271/A NOR2X1_LOC_755/Y -0.00fF
C40501 NOR2X1_LOC_457/A INVX1_LOC_9/A 0.07fF
C40502 INVX1_LOC_110/A VDD -0.00fF
C40503 INVX1_LOC_199/A INVX1_LOC_71/A 0.02fF
C40504 NOR2X1_LOC_383/Y NOR2X1_LOC_72/a_36_216# 0.01fF
C40505 NAND2X1_LOC_227/Y INVX1_LOC_118/A 0.00fF
C40506 NOR2X1_LOC_338/Y INVX1_LOC_76/A -0.02fF
C40507 NOR2X1_LOC_415/A INVX1_LOC_135/A 0.01fF
C40508 NOR2X1_LOC_454/Y INVX1_LOC_113/A 0.02fF
C40509 NAND2X1_LOC_537/Y INVX1_LOC_92/A 0.07fF
C40510 NAND2X1_LOC_231/Y INVX1_LOC_144/A 0.10fF
C40511 INVX1_LOC_108/Y NAND2X1_LOC_207/B 0.01fF
C40512 INVX1_LOC_35/A NOR2X1_LOC_777/B 0.03fF
C40513 NOR2X1_LOC_590/A INVX1_LOC_38/A 11.04fF
C40514 NOR2X1_LOC_392/Y NAND2X1_LOC_74/B 0.01fF
C40515 NOR2X1_LOC_419/Y INVX1_LOC_95/Y 0.31fF
C40516 INVX1_LOC_63/Y NOR2X1_LOC_41/a_36_216# 0.00fF
C40517 NOR2X1_LOC_546/A VDD -0.00fF
C40518 NOR2X1_LOC_598/B INVX1_LOC_99/A 0.02fF
C40519 NOR2X1_LOC_246/A NOR2X1_LOC_130/A 0.07fF
C40520 NOR2X1_LOC_196/A VDD 0.00fF
C40521 INVX1_LOC_24/A NOR2X1_LOC_357/Y 0.01fF
C40522 NOR2X1_LOC_716/B INVX1_LOC_95/Y 0.17fF
C40523 NOR2X1_LOC_208/a_36_216# INVX1_LOC_75/A 0.02fF
C40524 NAND2X1_LOC_409/a_36_24# INVX1_LOC_19/A -0.00fF
C40525 NAND2X1_LOC_773/Y NAND2X1_LOC_572/B 0.23fF
C40526 NOR2X1_LOC_220/A NOR2X1_LOC_188/A 0.08fF
C40527 NOR2X1_LOC_764/Y INVX1_LOC_295/A 0.12fF
C40528 INVX1_LOC_132/Y INVX1_LOC_148/Y 0.00fF
C40529 NAND2X1_LOC_551/A NOR2X1_LOC_130/A 0.07fF
C40530 D_INPUT_1 NOR2X1_LOC_554/A 0.02fF
C40531 INPUT_0 INVX1_LOC_56/A 0.01fF
C40532 INVX1_LOC_11/A NOR2X1_LOC_592/B 0.03fF
C40533 NOR2X1_LOC_220/A NOR2X1_LOC_548/B 0.10fF
C40534 INVX1_LOC_8/A NOR2X1_LOC_124/A 0.01fF
C40535 D_INPUT_2 NOR2X1_LOC_37/a_36_216# 0.00fF
C40536 INVX1_LOC_290/A INVX1_LOC_302/Y 0.16fF
C40537 INVX1_LOC_21/A NAND2X1_LOC_781/a_36_24# 0.00fF
C40538 NOR2X1_LOC_92/Y NOR2X1_LOC_653/Y 0.05fF
C40539 NOR2X1_LOC_355/A NOR2X1_LOC_356/A -0.01fF
C40540 INVX1_LOC_30/A INVX1_LOC_9/A 0.18fF
C40541 INVX1_LOC_13/A NOR2X1_LOC_112/B 0.05fF
C40542 NOR2X1_LOC_68/A INVX1_LOC_114/A 0.00fF
C40543 NOR2X1_LOC_292/Y INVX1_LOC_1/Y 0.01fF
C40544 NOR2X1_LOC_557/A NOR2X1_LOC_537/Y 0.07fF
C40545 NAND2X1_LOC_276/Y INVX1_LOC_20/A 0.00fF
C40546 NAND2X1_LOC_214/B INVX1_LOC_284/A 0.54fF
C40547 INVX1_LOC_223/Y NAND2X1_LOC_74/B 0.01fF
C40548 NAND2X1_LOC_338/B NOR2X1_LOC_557/A 0.02fF
C40549 INVX1_LOC_101/A NOR2X1_LOC_74/A 0.00fF
C40550 NOR2X1_LOC_500/A NAND2X1_LOC_417/a_36_24# 0.00fF
C40551 INVX1_LOC_135/A NAND2X1_LOC_293/a_36_24# 0.06fF
C40552 INVX1_LOC_163/A INVX1_LOC_163/Y 0.08fF
C40553 INVX1_LOC_24/A NOR2X1_LOC_692/Y 0.00fF
C40554 NOR2X1_LOC_92/Y INVX1_LOC_19/A 1.77fF
C40555 NOR2X1_LOC_576/B NAND2X1_LOC_560/A 0.02fF
C40556 NAND2X1_LOC_610/a_36_24# NAND2X1_LOC_642/Y 0.01fF
C40557 NOR2X1_LOC_548/B NOR2X1_LOC_548/Y 0.02fF
C40558 INVX1_LOC_24/Y INVX1_LOC_19/A 0.17fF
C40559 NOR2X1_LOC_781/A INVX1_LOC_6/A 0.01fF
C40560 INVX1_LOC_50/A NOR2X1_LOC_631/Y 0.03fF
C40561 INVX1_LOC_64/A INVX1_LOC_231/A 0.04fF
C40562 INVX1_LOC_43/Y NOR2X1_LOC_179/Y 0.01fF
C40563 NAND2X1_LOC_123/Y INVX1_LOC_313/Y 0.05fF
C40564 NOR2X1_LOC_190/a_36_216# INVX1_LOC_95/A 0.00fF
C40565 NOR2X1_LOC_355/A NOR2X1_LOC_74/A 0.01fF
C40566 NOR2X1_LOC_15/Y INVX1_LOC_29/A 3.08fF
C40567 INVX1_LOC_235/Y INVX1_LOC_42/A 0.00fF
C40568 INVX1_LOC_45/Y INVX1_LOC_54/A 0.06fF
C40569 NOR2X1_LOC_296/Y NAND2X1_LOC_773/B 0.03fF
C40570 INPUT_3 NAND2X1_LOC_206/Y 0.07fF
C40571 NOR2X1_LOC_433/A NOR2X1_LOC_331/B 0.17fF
C40572 INVX1_LOC_28/A INVX1_LOC_140/A 0.10fF
C40573 NOR2X1_LOC_68/A INVX1_LOC_307/A 0.10fF
C40574 NOR2X1_LOC_557/Y INVX1_LOC_66/Y 0.00fF
C40575 NAND2X1_LOC_374/Y INVX1_LOC_20/A 0.00fF
C40576 NOR2X1_LOC_593/Y NOR2X1_LOC_331/B 0.07fF
C40577 INVX1_LOC_54/Y INVX1_LOC_46/A 0.49fF
C40578 NOR2X1_LOC_68/A NOR2X1_LOC_445/B 0.10fF
C40579 NAND2X1_LOC_354/B INVX1_LOC_38/A 0.01fF
C40580 INVX1_LOC_6/A NOR2X1_LOC_76/A 0.07fF
C40581 NAND2X1_LOC_133/a_36_24# INVX1_LOC_123/A 0.00fF
C40582 NOR2X1_LOC_860/B INVX1_LOC_152/A 0.03fF
C40583 NOR2X1_LOC_736/Y NOR2X1_LOC_74/A 0.09fF
C40584 INVX1_LOC_151/A NOR2X1_LOC_331/B 0.03fF
C40585 INVX1_LOC_88/A NAND2X1_LOC_792/B 0.01fF
C40586 NAND2X1_LOC_352/B NAND2X1_LOC_81/B 0.05fF
C40587 NOR2X1_LOC_45/Y INVX1_LOC_272/A 0.01fF
C40588 NOR2X1_LOC_552/Y NOR2X1_LOC_356/A 0.01fF
C40589 NOR2X1_LOC_825/Y INVX1_LOC_316/Y 0.03fF
C40590 NAND2X1_LOC_578/a_36_24# INVX1_LOC_15/A 0.00fF
C40591 NAND2X1_LOC_171/a_36_24# NOR2X1_LOC_633/A 0.00fF
C40592 NOR2X1_LOC_103/Y NAND2X1_LOC_254/Y 0.01fF
C40593 INVX1_LOC_21/A NOR2X1_LOC_334/Y 0.09fF
C40594 INVX1_LOC_286/Y INVX1_LOC_264/A 0.02fF
C40595 NOR2X1_LOC_52/B NOR2X1_LOC_331/B 5.04fF
C40596 NOR2X1_LOC_468/a_36_216# INVX1_LOC_93/Y 0.01fF
C40597 INVX1_LOC_251/Y NOR2X1_LOC_536/A 0.03fF
C40598 NOR2X1_LOC_433/A NOR2X1_LOC_592/B 0.03fF
C40599 NAND2X1_LOC_859/Y NAND2X1_LOC_241/Y 0.01fF
C40600 INVX1_LOC_33/A NOR2X1_LOC_364/A 0.14fF
C40601 INVX1_LOC_245/A INVX1_LOC_37/A 0.01fF
C40602 NAND2X1_LOC_149/Y INVX1_LOC_78/A 0.68fF
C40603 NOR2X1_LOC_591/A NAND2X1_LOC_590/a_36_24# 0.02fF
C40604 NOR2X1_LOC_486/B INVX1_LOC_92/A -0.02fF
C40605 INVX1_LOC_34/A NOR2X1_LOC_155/A 0.06fF
C40606 INVX1_LOC_24/A NAND2X1_LOC_489/Y 0.06fF
C40607 INVX1_LOC_53/A NOR2X1_LOC_634/Y 0.01fF
C40608 NOR2X1_LOC_332/A NOR2X1_LOC_35/Y 0.10fF
C40609 NOR2X1_LOC_520/B NAND2X1_LOC_85/Y 0.00fF
C40610 INVX1_LOC_282/A INVX1_LOC_309/A 0.07fF
C40611 INVX1_LOC_170/A NOR2X1_LOC_76/B 0.02fF
C40612 INVX1_LOC_45/A NAND2X1_LOC_254/Y 0.27fF
C40613 INVX1_LOC_33/A INVX1_LOC_285/A 0.07fF
C40614 INVX1_LOC_298/Y NOR2X1_LOC_15/Y 0.07fF
C40615 INVX1_LOC_93/Y NOR2X1_LOC_153/a_36_216# 0.01fF
C40616 NOR2X1_LOC_52/B NOR2X1_LOC_592/B 0.03fF
C40617 D_INPUT_0 INVX1_LOC_2/Y 0.15fF
C40618 NAND2X1_LOC_838/Y NOR2X1_LOC_491/Y 0.05fF
C40619 NAND2X1_LOC_859/Y NAND2X1_LOC_837/a_36_24# 0.01fF
C40620 INVX1_LOC_21/A NAND2X1_LOC_464/B 0.07fF
C40621 NOR2X1_LOC_432/Y NOR2X1_LOC_433/Y 0.03fF
C40622 NOR2X1_LOC_68/A INVX1_LOC_12/A 0.18fF
C40623 NOR2X1_LOC_246/A NOR2X1_LOC_280/Y 0.29fF
C40624 INVX1_LOC_251/Y NAND2X1_LOC_93/B 0.02fF
C40625 INVX1_LOC_282/A INVX1_LOC_91/A 0.07fF
C40626 INVX1_LOC_33/A NOR2X1_LOC_814/A 0.28fF
C40627 INVX1_LOC_24/Y INVX1_LOC_26/Y 0.06fF
C40628 NOR2X1_LOC_837/B NOR2X1_LOC_777/B 0.42fF
C40629 INVX1_LOC_11/A NAND2X1_LOC_467/a_36_24# 0.00fF
C40630 NAND2X1_LOC_645/a_36_24# NOR2X1_LOC_331/B 0.00fF
C40631 NOR2X1_LOC_188/A NAND2X1_LOC_498/a_36_24# 0.01fF
C40632 NOR2X1_LOC_78/B NOR2X1_LOC_78/Y 0.03fF
C40633 NOR2X1_LOC_567/B NOR2X1_LOC_542/B 0.02fF
C40634 NOR2X1_LOC_860/B INVX1_LOC_29/A 0.07fF
C40635 INVX1_LOC_210/Y INVX1_LOC_15/A 0.00fF
C40636 NOR2X1_LOC_829/Y NOR2X1_LOC_15/Y 0.00fF
C40637 NOR2X1_LOC_533/a_36_216# INVX1_LOC_76/A 0.01fF
C40638 NOR2X1_LOC_604/Y INVX1_LOC_27/A 0.03fF
C40639 INVX1_LOC_233/A INVX1_LOC_93/A 1.14fF
C40640 NAND2X1_LOC_525/a_36_24# NOR2X1_LOC_486/Y 0.00fF
C40641 INVX1_LOC_282/A INVX1_LOC_11/Y 0.07fF
C40642 INVX1_LOC_256/A NOR2X1_LOC_541/B 0.01fF
C40643 NOR2X1_LOC_567/B INVX1_LOC_143/Y 0.01fF
C40644 NOR2X1_LOC_590/A NAND2X1_LOC_223/A 0.12fF
C40645 INVX1_LOC_41/A INVX1_LOC_19/A 0.34fF
C40646 NAND2X1_LOC_477/A NOR2X1_LOC_653/Y 0.02fF
C40647 NOR2X1_LOC_292/Y INVX1_LOC_93/Y 0.03fF
C40648 NOR2X1_LOC_564/Y VDD 0.35fF
C40649 INVX1_LOC_51/Y NOR2X1_LOC_100/a_36_216# 0.02fF
C40650 NAND2X1_LOC_341/A INVX1_LOC_117/Y 0.03fF
C40651 INVX1_LOC_69/Y NOR2X1_LOC_552/A 1.56fF
C40652 NOR2X1_LOC_590/A INVX1_LOC_18/Y 0.06fF
C40653 NOR2X1_LOC_646/A INVX1_LOC_46/Y 0.06fF
C40654 INVX1_LOC_126/A NOR2X1_LOC_74/A 0.03fF
C40655 NOR2X1_LOC_824/A NAND2X1_LOC_623/a_36_24# 0.00fF
C40656 NAND2X1_LOC_537/Y INVX1_LOC_53/A 0.07fF
C40657 INVX1_LOC_286/Y NOR2X1_LOC_25/Y 0.02fF
C40658 INVX1_LOC_24/A INVX1_LOC_32/A 0.15fF
C40659 NAND2X1_LOC_477/A INVX1_LOC_19/A 4.38fF
C40660 NOR2X1_LOC_272/Y INVX1_LOC_306/Y 0.10fF
C40661 NOR2X1_LOC_388/Y NOR2X1_LOC_89/A 0.07fF
C40662 INVX1_LOC_36/A NOR2X1_LOC_464/Y 0.01fF
C40663 NOR2X1_LOC_32/B INVX1_LOC_14/A 0.45fF
C40664 NAND2X1_LOC_357/B NAND2X1_LOC_81/B 0.10fF
C40665 INVX1_LOC_6/A NAND2X1_LOC_241/Y 0.02fF
C40666 NAND2X1_LOC_660/A INVX1_LOC_49/Y 0.13fF
C40667 NOR2X1_LOC_543/a_36_216# NOR2X1_LOC_552/A 0.01fF
C40668 NAND2X1_LOC_141/A INVX1_LOC_29/A 0.03fF
C40669 INVX1_LOC_316/Y INVX1_LOC_84/A 0.01fF
C40670 D_INPUT_1 NOR2X1_LOC_160/B 0.17fF
C40671 NOR2X1_LOC_15/Y NOR2X1_LOC_291/a_36_216# 0.00fF
C40672 NOR2X1_LOC_216/Y INVX1_LOC_66/Y 0.19fF
C40673 INVX1_LOC_27/A NAND2X1_LOC_85/a_36_24# 0.00fF
C40674 D_INPUT_0 NOR2X1_LOC_608/Y 0.00fF
C40675 NAND2X1_LOC_565/B NAND2X1_LOC_489/Y 0.01fF
C40676 INVX1_LOC_226/Y NAND2X1_LOC_768/Y 0.01fF
C40677 INVX1_LOC_249/Y INVX1_LOC_283/A 0.15fF
C40678 INVX1_LOC_24/A NAND2X1_LOC_175/Y 0.19fF
C40679 INVX1_LOC_193/Y NOR2X1_LOC_706/a_36_216# 0.00fF
C40680 NAND2X1_LOC_440/a_36_24# NOR2X1_LOC_269/Y 0.00fF
C40681 NOR2X1_LOC_264/Y INVX1_LOC_15/A 0.03fF
C40682 INVX1_LOC_226/A INVX1_LOC_29/A 0.03fF
C40683 INVX1_LOC_72/A INVX1_LOC_271/A 0.16fF
C40684 NAND2X1_LOC_705/Y NAND2X1_LOC_493/Y 0.02fF
C40685 NOR2X1_LOC_344/A INVX1_LOC_4/Y 0.07fF
C40686 INVX1_LOC_17/A NOR2X1_LOC_249/Y 0.00fF
C40687 NAND2X1_LOC_725/A INVX1_LOC_161/A 0.10fF
C40688 INVX1_LOC_72/A INVX1_LOC_105/Y 0.03fF
C40689 NOR2X1_LOC_366/B NOR2X1_LOC_89/A 0.06fF
C40690 INVX1_LOC_25/Y NAND2X1_LOC_74/B 0.17fF
C40691 INVX1_LOC_17/A NOR2X1_LOC_846/A 0.06fF
C40692 NAND2X1_LOC_842/B NOR2X1_LOC_216/B 0.01fF
C40693 NOR2X1_LOC_186/Y INVX1_LOC_150/Y 0.12fF
C40694 INVX1_LOC_182/A INVX1_LOC_179/A 0.02fF
C40695 NAND2X1_LOC_830/a_36_24# NOR2X1_LOC_831/B 0.00fF
C40696 NAND2X1_LOC_794/B NOR2X1_LOC_816/A 0.22fF
C40697 NOR2X1_LOC_160/B NOR2X1_LOC_652/Y 0.46fF
C40698 NOR2X1_LOC_486/Y NOR2X1_LOC_562/A 0.13fF
C40699 NOR2X1_LOC_130/A NAND2X1_LOC_489/Y 0.03fF
C40700 NOR2X1_LOC_87/B NOR2X1_LOC_38/B 0.24fF
C40701 INVX1_LOC_75/A INVX1_LOC_75/Y 0.04fF
C40702 INVX1_LOC_131/A NOR2X1_LOC_155/A 0.02fF
C40703 INVX1_LOC_136/A NOR2X1_LOC_392/Y 0.00fF
C40704 NAND2X1_LOC_661/B INVX1_LOC_15/A 0.08fF
C40705 NAND2X1_LOC_392/A INVX1_LOC_102/A 0.05fF
C40706 INVX1_LOC_143/A INVX1_LOC_32/A 0.07fF
C40707 INVX1_LOC_103/A NOR2X1_LOC_666/A 0.02fF
C40708 NOR2X1_LOC_443/Y INVX1_LOC_184/Y 0.00fF
C40709 INVX1_LOC_35/A NOR2X1_LOC_647/Y 0.18fF
C40710 NAND2X1_LOC_557/Y NAND2X1_LOC_837/Y 0.03fF
C40711 INVX1_LOC_178/A INVX1_LOC_246/A 0.10fF
C40712 NAND2X1_LOC_555/Y NOR2X1_LOC_249/Y 0.05fF
C40713 INVX1_LOC_16/A INVX1_LOC_42/A 0.43fF
C40714 NOR2X1_LOC_45/B NOR2X1_LOC_536/A 0.17fF
C40715 INVX1_LOC_35/A INVX1_LOC_18/A 0.24fF
C40716 INVX1_LOC_143/A NOR2X1_LOC_623/B -0.02fF
C40717 INVX1_LOC_41/A INVX1_LOC_26/Y 0.13fF
C40718 NOR2X1_LOC_92/Y INVX1_LOC_161/Y 0.07fF
C40719 INVX1_LOC_39/A INVX1_LOC_61/Y 0.25fF
C40720 INVX1_LOC_254/Y INVX1_LOC_57/A 0.02fF
C40721 NAND2X1_LOC_1/Y INVX1_LOC_37/A 0.00fF
C40722 INVX1_LOC_181/Y NOR2X1_LOC_717/A 0.01fF
C40723 INPUT_0 NOR2X1_LOC_155/A 0.00fF
C40724 INVX1_LOC_234/A INVX1_LOC_284/A 0.17fF
C40725 NOR2X1_LOC_551/B NOR2X1_LOC_383/B 0.02fF
C40726 INVX1_LOC_73/A NOR2X1_LOC_117/Y 0.01fF
C40727 NOR2X1_LOC_315/Y NOR2X1_LOC_693/a_36_216# 0.00fF
C40728 INVX1_LOC_316/Y INVX1_LOC_15/A 0.03fF
C40729 NOR2X1_LOC_846/Y INVX1_LOC_36/A 0.01fF
C40730 INVX1_LOC_249/A NOR2X1_LOC_604/Y 0.15fF
C40731 NAND2X1_LOC_778/Y NAND2X1_LOC_721/B 0.03fF
C40732 INVX1_LOC_135/A NOR2X1_LOC_89/A 0.10fF
C40733 NOR2X1_LOC_689/Y INVX1_LOC_34/A 0.03fF
C40734 INVX1_LOC_17/Y NOR2X1_LOC_690/A 0.02fF
C40735 INVX1_LOC_298/Y INVX1_LOC_96/Y 0.01fF
C40736 INVX1_LOC_35/A NOR2X1_LOC_713/B 0.01fF
C40737 NAND2X1_LOC_568/A INVX1_LOC_161/Y 0.00fF
C40738 NOR2X1_LOC_323/Y INVX1_LOC_285/A 0.01fF
C40739 INVX1_LOC_201/Y INVX1_LOC_166/A 0.59fF
C40740 NOR2X1_LOC_601/Y NOR2X1_LOC_331/B 0.03fF
C40741 INVX1_LOC_240/A NAND2X1_LOC_401/a_36_24# 0.00fF
C40742 INVX1_LOC_27/A INVX1_LOC_72/A 0.19fF
C40743 NOR2X1_LOC_824/A INVX1_LOC_72/A 0.07fF
C40744 INVX1_LOC_48/Y NOR2X1_LOC_90/a_36_216# 0.00fF
C40745 NOR2X1_LOC_92/Y INVX1_LOC_312/A 0.03fF
C40746 NOR2X1_LOC_554/a_36_216# NOR2X1_LOC_660/Y 0.00fF
C40747 NOR2X1_LOC_391/Y INVX1_LOC_123/Y 0.00fF
C40748 NOR2X1_LOC_682/Y NAND2X1_LOC_687/A 0.08fF
C40749 NOR2X1_LOC_92/Y NOR2X1_LOC_599/A 0.06fF
C40750 NOR2X1_LOC_160/B NOR2X1_LOC_241/A 0.14fF
C40751 NOR2X1_LOC_769/A NAND2X1_LOC_149/Y 0.03fF
C40752 INVX1_LOC_230/Y NOR2X1_LOC_82/A 0.12fF
C40753 NOR2X1_LOC_598/B INVX1_LOC_34/A 0.03fF
C40754 INVX1_LOC_90/A NOR2X1_LOC_67/Y 0.03fF
C40755 INVX1_LOC_237/A INVX1_LOC_72/A 0.03fF
C40756 INVX1_LOC_57/Y NAND2X1_LOC_579/A 0.16fF
C40757 NOR2X1_LOC_32/B INVX1_LOC_217/Y 0.00fF
C40758 NOR2X1_LOC_731/A INVX1_LOC_23/A 0.03fF
C40759 INVX1_LOC_16/A INVX1_LOC_78/A 0.03fF
C40760 INVX1_LOC_278/A NAND2X1_LOC_569/A -0.02fF
C40761 NOR2X1_LOC_91/A NAND2X1_LOC_181/Y 0.03fF
C40762 NOR2X1_LOC_130/A INVX1_LOC_32/A 0.17fF
C40763 NOR2X1_LOC_456/Y NOR2X1_LOC_348/B 0.26fF
C40764 NAND2X1_LOC_833/Y NOR2X1_LOC_109/Y 0.01fF
C40765 NOR2X1_LOC_798/A NOR2X1_LOC_303/Y 0.00fF
C40766 NOR2X1_LOC_15/Y NAND2X1_LOC_634/Y 0.13fF
C40767 NOR2X1_LOC_19/B INVX1_LOC_284/A 0.07fF
C40768 INVX1_LOC_92/Y INVX1_LOC_63/A 0.04fF
C40769 INVX1_LOC_34/A NAND2X1_LOC_725/A 0.40fF
C40770 INVX1_LOC_77/A NOR2X1_LOC_460/Y 0.04fF
C40771 INVX1_LOC_28/A INVX1_LOC_42/A 0.15fF
C40772 INVX1_LOC_75/A NAND2X1_LOC_74/B 0.03fF
C40773 INVX1_LOC_150/A NAND2X1_LOC_647/B 0.01fF
C40774 INVX1_LOC_59/Y NOR2X1_LOC_660/a_36_216# 0.00fF
C40775 NOR2X1_LOC_550/a_36_216# NOR2X1_LOC_794/B 0.00fF
C40776 NOR2X1_LOC_211/A INVX1_LOC_26/Y 0.21fF
C40777 INVX1_LOC_43/A NOR2X1_LOC_383/B 0.29fF
C40778 NOR2X1_LOC_169/B NOR2X1_LOC_457/A 0.01fF
C40779 NOR2X1_LOC_528/Y INVX1_LOC_119/Y 0.16fF
C40780 INVX1_LOC_147/A INVX1_LOC_12/A 0.11fF
C40781 INVX1_LOC_136/A NAND2X1_LOC_357/A 0.07fF
C40782 NOR2X1_LOC_784/Y NOR2X1_LOC_148/A 0.02fF
C40783 NAND2X1_LOC_30/Y D_INPUT_7 0.95fF
C40784 NAND2X1_LOC_149/Y NOR2X1_LOC_152/Y 0.02fF
C40785 NOR2X1_LOC_65/B INVX1_LOC_16/A 0.07fF
C40786 NOR2X1_LOC_717/B INVX1_LOC_271/Y 0.01fF
C40787 NOR2X1_LOC_276/B INVX1_LOC_103/A 0.01fF
C40788 NOR2X1_LOC_2/Y INVX1_LOC_12/A 0.01fF
C40789 NAND2X1_LOC_181/Y INVX1_LOC_23/A 0.33fF
C40790 NAND2X1_LOC_714/B NOR2X1_LOC_577/Y 0.07fF
C40791 INVX1_LOC_75/A NOR2X1_LOC_847/B 0.03fF
C40792 NAND2X1_LOC_35/Y NOR2X1_LOC_821/Y 0.01fF
C40793 NAND2X1_LOC_860/A NOR2X1_LOC_78/B 0.07fF
C40794 NAND2X1_LOC_783/A NAND2X1_LOC_175/Y 0.12fF
C40795 NOR2X1_LOC_91/A NAND2X1_LOC_390/A -0.00fF
C40796 INVX1_LOC_88/A NOR2X1_LOC_359/Y 0.00fF
C40797 NOR2X1_LOC_45/B NOR2X1_LOC_661/A 0.03fF
C40798 NAND2X1_LOC_848/A NAND2X1_LOC_846/a_36_24# 0.02fF
C40799 NOR2X1_LOC_634/B NOR2X1_LOC_634/Y 0.01fF
C40800 D_INPUT_1 INVX1_LOC_208/A 0.08fF
C40801 NOR2X1_LOC_130/A NAND2X1_LOC_175/Y 0.19fF
C40802 INVX1_LOC_2/Y INVX1_LOC_46/Y 0.01fF
C40803 NAND2X1_LOC_724/Y NAND2X1_LOC_857/a_36_24# 0.01fF
C40804 NAND2X1_LOC_725/Y NAND2X1_LOC_863/B 0.06fF
C40805 NAND2X1_LOC_656/B INVX1_LOC_46/A 0.02fF
C40806 NOR2X1_LOC_188/A NAND2X1_LOC_200/a_36_24# 0.00fF
C40807 INVX1_LOC_5/A NOR2X1_LOC_84/Y -0.03fF
C40808 NAND2X1_LOC_579/A NAND2X1_LOC_632/B 0.02fF
C40809 INVX1_LOC_64/A NAND2X1_LOC_374/Y 0.10fF
C40810 D_INPUT_1 NOR2X1_LOC_516/B 0.08fF
C40811 INVX1_LOC_136/A NOR2X1_LOC_599/Y 0.11fF
C40812 NOR2X1_LOC_277/a_36_216# NAND2X1_LOC_181/Y 0.00fF
C40813 NAND2X1_LOC_773/Y NOR2X1_LOC_716/B 0.10fF
C40814 NOR2X1_LOC_828/A INVX1_LOC_271/Y 0.00fF
C40815 INVX1_LOC_21/A NOR2X1_LOC_718/B 0.07fF
C40816 NOR2X1_LOC_788/B NAND2X1_LOC_72/B 0.03fF
C40817 NAND2X1_LOC_785/a_36_24# NAND2X1_LOC_722/A 0.00fF
C40818 INVX1_LOC_123/A NAND2X1_LOC_207/B 0.01fF
C40819 NOR2X1_LOC_334/A NAND2X1_LOC_291/B 0.01fF
C40820 NAND2X1_LOC_514/a_36_24# INVX1_LOC_23/A 0.01fF
C40821 INVX1_LOC_269/A NOR2X1_LOC_335/A 0.03fF
C40822 NOR2X1_LOC_456/Y INVX1_LOC_22/A 0.05fF
C40823 INVX1_LOC_90/A NOR2X1_LOC_415/Y 0.00fF
C40824 NOR2X1_LOC_690/A NAND2X1_LOC_493/Y 0.15fF
C40825 INVX1_LOC_225/Y INVX1_LOC_94/A 0.25fF
C40826 INVX1_LOC_281/A NAND2X1_LOC_93/B 0.07fF
C40827 INVX1_LOC_1/A INVX1_LOC_63/Y 0.10fF
C40828 INPUT_3 INVX1_LOC_24/A 0.03fF
C40829 INVX1_LOC_28/A INVX1_LOC_78/A 0.31fF
C40830 NOR2X1_LOC_798/A INVX1_LOC_54/Y 0.00fF
C40831 NOR2X1_LOC_286/Y NAND2X1_LOC_364/Y 0.01fF
C40832 NOR2X1_LOC_99/Y NOR2X1_LOC_271/Y 0.06fF
C40833 NAND2X1_LOC_860/A NAND2X1_LOC_392/Y 0.04fF
C40834 NOR2X1_LOC_189/A NOR2X1_LOC_816/A 0.03fF
C40835 INVX1_LOC_27/A NOR2X1_LOC_537/Y 0.07fF
C40836 INVX1_LOC_103/A INVX1_LOC_103/Y 0.11fF
C40837 NAND2X1_LOC_93/B NOR2X1_LOC_378/Y 0.06fF
C40838 INVX1_LOC_27/A NAND2X1_LOC_338/B 1.46fF
C40839 INVX1_LOC_136/A NOR2X1_LOC_86/Y 0.02fF
C40840 NOR2X1_LOC_825/Y NOR2X1_LOC_662/A 0.07fF
C40841 NAND2X1_LOC_108/a_36_24# INVX1_LOC_29/A 0.01fF
C40842 NAND2X1_LOC_794/B NOR2X1_LOC_773/Y 0.07fF
C40843 NOR2X1_LOC_151/Y INVX1_LOC_271/Y 0.05fF
C40844 INVX1_LOC_36/A NOR2X1_LOC_457/B 0.09fF
C40845 D_INPUT_1 NAND2X1_LOC_133/a_36_24# 0.01fF
C40846 INVX1_LOC_64/A NOR2X1_LOC_553/B 0.04fF
C40847 NOR2X1_LOC_378/Y NAND2X1_LOC_425/Y -0.02fF
C40848 INVX1_LOC_5/A INVX1_LOC_290/A 0.24fF
C40849 INVX1_LOC_17/A NAND2X1_LOC_116/A 0.03fF
C40850 NOR2X1_LOC_65/B INVX1_LOC_28/A 0.50fF
C40851 INVX1_LOC_45/A INVX1_LOC_314/Y 0.03fF
C40852 NOR2X1_LOC_620/Y INVX1_LOC_31/A 0.16fF
C40853 NOR2X1_LOC_748/Y INVX1_LOC_50/Y 0.05fF
C40854 NOR2X1_LOC_759/A INVX1_LOC_159/A 0.15fF
C40855 NOR2X1_LOC_590/A INVX1_LOC_33/A 0.16fF
C40856 INVX1_LOC_83/A NOR2X1_LOC_634/Y 0.00fF
C40857 INVX1_LOC_225/A INVX1_LOC_150/Y 0.30fF
C40858 NOR2X1_LOC_292/Y INVX1_LOC_87/A 0.04fF
C40859 VDD INVX1_LOC_264/A 0.30fF
C40860 NOR2X1_LOC_590/A NOR2X1_LOC_743/a_36_216# 0.00fF
C40861 NOR2X1_LOC_808/A NOR2X1_LOC_793/Y 0.00fF
C40862 INVX1_LOC_161/Y NAND2X1_LOC_477/A 0.07fF
C40863 NAND2X1_LOC_800/A INVX1_LOC_264/A 0.02fF
C40864 NAND2X1_LOC_453/A NAND2X1_LOC_74/B 0.68fF
C40865 NOR2X1_LOC_209/Y NOR2X1_LOC_740/Y 0.32fF
C40866 NOR2X1_LOC_552/A NOR2X1_LOC_170/A 0.03fF
C40867 NOR2X1_LOC_786/a_36_216# NOR2X1_LOC_84/Y 0.00fF
C40868 INVX1_LOC_21/A NOR2X1_LOC_569/Y 0.07fF
C40869 NOR2X1_LOC_65/a_36_216# NAND2X1_LOC_74/B 0.01fF
C40870 NOR2X1_LOC_253/Y INVX1_LOC_42/A 0.08fF
C40871 INVX1_LOC_73/A INVX1_LOC_270/A 0.07fF
C40872 NOR2X1_LOC_75/Y NOR2X1_LOC_432/a_36_216# 0.00fF
C40873 NOR2X1_LOC_167/a_36_216# NOR2X1_LOC_167/Y 0.00fF
C40874 INVX1_LOC_46/Y NOR2X1_LOC_608/Y 0.02fF
C40875 NOR2X1_LOC_89/A INVX1_LOC_139/Y 0.03fF
C40876 NOR2X1_LOC_88/Y NOR2X1_LOC_510/B 0.34fF
C40877 NOR2X1_LOC_45/B NAND2X1_LOC_470/B 0.09fF
C40878 INVX1_LOC_10/A NAND2X1_LOC_474/Y 0.07fF
C40879 NOR2X1_LOC_569/a_36_216# INVX1_LOC_53/A 0.01fF
C40880 NOR2X1_LOC_778/B NOR2X1_LOC_541/Y 0.06fF
C40881 NOR2X1_LOC_54/a_36_216# INVX1_LOC_63/A 0.00fF
C40882 NOR2X1_LOC_689/Y INPUT_0 0.03fF
C40883 INVX1_LOC_314/Y INVX1_LOC_71/A 0.10fF
C40884 NOR2X1_LOC_335/B INVX1_LOC_57/A 0.07fF
C40885 NAND2X1_LOC_858/B NOR2X1_LOC_654/A 0.00fF
C40886 INVX1_LOC_30/A NOR2X1_LOC_367/B 0.01fF
C40887 INVX1_LOC_17/A INVX1_LOC_232/A 0.07fF
C40888 NOR2X1_LOC_778/A NOR2X1_LOC_317/B 0.04fF
C40889 INVX1_LOC_286/Y INVX1_LOC_236/A 0.00fF
C40890 INVX1_LOC_83/A NAND2X1_LOC_473/A 0.09fF
C40891 INVX1_LOC_59/A NAND2X1_LOC_531/a_36_24# 0.00fF
C40892 INVX1_LOC_75/A NOR2X1_LOC_660/Y 0.05fF
C40893 NOR2X1_LOC_19/B NOR2X1_LOC_663/A 0.01fF
C40894 NOR2X1_LOC_181/A INVX1_LOC_271/Y 0.03fF
C40895 NAND2X1_LOC_738/B NOR2X1_LOC_387/A 0.11fF
C40896 NOR2X1_LOC_598/B INPUT_0 0.20fF
C40897 INVX1_LOC_45/Y NOR2X1_LOC_142/Y 0.07fF
C40898 INVX1_LOC_18/A INVX1_LOC_257/Y 0.14fF
C40899 INVX1_LOC_101/Y NAND2X1_LOC_656/Y 0.03fF
C40900 NOR2X1_LOC_590/A INVX1_LOC_40/A 0.41fF
C40901 NAND2X1_LOC_524/a_36_24# INVX1_LOC_77/A 0.01fF
C40902 NOR2X1_LOC_67/Y INVX1_LOC_38/A 0.12fF
C40903 NOR2X1_LOC_723/a_36_216# INVX1_LOC_266/Y 0.01fF
C40904 INVX1_LOC_243/A INVX1_LOC_30/A 0.02fF
C40905 INVX1_LOC_51/A INPUT_0 0.00fF
C40906 INVX1_LOC_45/A NOR2X1_LOC_778/B 0.03fF
C40907 INVX1_LOC_297/A NAND2X1_LOC_771/a_36_24# 0.02fF
C40908 INVX1_LOC_83/A NAND2X1_LOC_537/Y 0.01fF
C40909 INVX1_LOC_30/A INVX1_LOC_179/Y 0.73fF
C40910 NOR2X1_LOC_690/A NOR2X1_LOC_495/Y 0.01fF
C40911 NAND2X1_LOC_763/B INVX1_LOC_243/A 0.02fF
C40912 NAND2X1_LOC_794/B INVX1_LOC_140/A 0.10fF
C40913 NAND2X1_LOC_725/A INPUT_0 0.19fF
C40914 D_INPUT_1 INVX1_LOC_315/Y 0.02fF
C40915 NAND2X1_LOC_33/a_36_24# NAND2X1_LOC_462/B -0.00fF
C40916 NOR2X1_LOC_300/Y NOR2X1_LOC_596/A 0.01fF
C40917 NAND2X1_LOC_338/B NAND2X1_LOC_338/a_36_24# 0.01fF
C40918 INVX1_LOC_192/A INVX1_LOC_49/A 0.04fF
C40919 INVX1_LOC_11/A INVX1_LOC_135/A 0.11fF
C40920 INVX1_LOC_94/A INVX1_LOC_266/Y 0.00fF
C40921 NOR2X1_LOC_388/Y NOR2X1_LOC_593/Y 0.07fF
C40922 NOR2X1_LOC_438/a_36_216# NAND2X1_LOC_861/Y 0.01fF
C40923 VDD NOR2X1_LOC_158/Y 0.86fF
C40924 NAND2X1_LOC_624/B INVX1_LOC_309/A 0.05fF
C40925 D_INPUT_6 D_INPUT_4 0.01fF
C40926 NOR2X1_LOC_321/Y NOR2X1_LOC_329/B 1.03fF
C40927 INVX1_LOC_11/A INVX1_LOC_295/A 4.74fF
C40928 VDD NOR2X1_LOC_25/Y 0.60fF
C40929 INVX1_LOC_136/A INVX1_LOC_25/Y 0.05fF
C40930 NOR2X1_LOC_272/Y NOR2X1_LOC_74/A 0.10fF
C40931 INVX1_LOC_84/A NOR2X1_LOC_662/A 0.07fF
C40932 NOR2X1_LOC_829/A INVX1_LOC_46/A 0.03fF
C40933 INVX1_LOC_49/A NOR2X1_LOC_802/A 0.07fF
C40934 NOR2X1_LOC_309/Y NAND2X1_LOC_833/Y 0.03fF
C40935 INPUT_3 NOR2X1_LOC_130/A 0.01fF
C40936 NOR2X1_LOC_91/A NOR2X1_LOC_314/Y 0.01fF
C40937 NOR2X1_LOC_216/B INVX1_LOC_284/A 1.77fF
C40938 INVX1_LOC_36/A NOR2X1_LOC_781/A 0.00fF
C40939 INVX1_LOC_34/A NAND2X1_LOC_308/Y 0.04fF
C40940 NOR2X1_LOC_778/B INVX1_LOC_71/A 3.92fF
C40941 NOR2X1_LOC_561/Y INVX1_LOC_30/A 0.22fF
C40942 NAND2X1_LOC_286/B INVX1_LOC_46/A 0.02fF
C40943 NAND2X1_LOC_787/A NOR2X1_LOC_164/a_36_216# 0.00fF
C40944 INVX1_LOC_136/Y INVX1_LOC_19/A 0.01fF
C40945 INVX1_LOC_238/A NOR2X1_LOC_576/B 0.04fF
C40946 NOR2X1_LOC_272/Y NOR2X1_LOC_9/Y 0.10fF
C40947 NAND2X1_LOC_99/Y NAND2X1_LOC_338/B 0.04fF
C40948 NOR2X1_LOC_636/A NAND2X1_LOC_451/Y 0.04fF
C40949 NOR2X1_LOC_392/B INVX1_LOC_104/A 0.00fF
C40950 NAND2X1_LOC_53/Y NOR2X1_LOC_302/Y 0.05fF
C40951 NOR2X1_LOC_273/Y INVX1_LOC_22/A 0.01fF
C40952 NOR2X1_LOC_246/A INVX1_LOC_286/Y 0.28fF
C40953 INVX1_LOC_50/A INVX1_LOC_14/Y 0.03fF
C40954 NOR2X1_LOC_433/A NOR2X1_LOC_366/B 0.02fF
C40955 NOR2X1_LOC_759/Y INVX1_LOC_22/A 0.02fF
C40956 NOR2X1_LOC_668/Y INVX1_LOC_117/A 0.02fF
C40957 NOR2X1_LOC_516/B D_INPUT_2 0.12fF
C40958 NOR2X1_LOC_218/Y INVX1_LOC_81/A 0.80fF
C40959 INPUT_0 NOR2X1_LOC_271/a_36_216# 0.00fF
C40960 NAND2X1_LOC_787/A INVX1_LOC_76/A 0.03fF
C40961 INVX1_LOC_106/A INVX1_LOC_63/A 0.01fF
C40962 INVX1_LOC_37/A NOR2X1_LOC_452/A 0.01fF
C40963 INVX1_LOC_36/A NOR2X1_LOC_76/A 1.20fF
C40964 INVX1_LOC_103/A NOR2X1_LOC_313/Y 0.02fF
C40965 NOR2X1_LOC_68/A NAND2X1_LOC_808/A 0.01fF
C40966 NAND2X1_LOC_860/A INVX1_LOC_46/A 0.10fF
C40967 INVX1_LOC_113/Y INVX1_LOC_16/A 0.03fF
C40968 INVX1_LOC_45/A NOR2X1_LOC_724/Y 0.03fF
C40969 INVX1_LOC_33/A NOR2X1_LOC_82/Y 0.03fF
C40970 NOR2X1_LOC_336/B NOR2X1_LOC_356/A 0.00fF
C40971 INVX1_LOC_23/A INVX1_LOC_117/A 0.39fF
C40972 NOR2X1_LOC_276/Y INVX1_LOC_75/A 0.05fF
C40973 NAND2X1_LOC_338/B NAND2X1_LOC_471/a_36_24# 0.00fF
C40974 NAND2X1_LOC_454/Y INVX1_LOC_92/A 0.07fF
C40975 NOR2X1_LOC_68/A NOR2X1_LOC_155/a_36_216# 0.00fF
C40976 D_INPUT_6 INPUT_4 0.29fF
C40977 NOR2X1_LOC_791/B INPUT_1 0.88fF
C40978 NAND2X1_LOC_381/Y NOR2X1_LOC_391/B 0.00fF
C40979 INVX1_LOC_45/A NAND2X1_LOC_123/Y 0.03fF
C40980 INVX1_LOC_38/A NOR2X1_LOC_441/a_36_216# 0.00fF
C40981 NOR2X1_LOC_772/A INVX1_LOC_72/A 0.00fF
C40982 NAND2X1_LOC_392/A INVX1_LOC_162/Y 0.03fF
C40983 INVX1_LOC_99/A INVX1_LOC_29/A 0.07fF
C40984 INVX1_LOC_20/A NOR2X1_LOC_81/Y 0.01fF
C40985 INVX1_LOC_90/A NAND2X1_LOC_357/a_36_24# 0.00fF
C40986 INVX1_LOC_25/Y NOR2X1_LOC_278/A 0.06fF
C40987 NAND2X1_LOC_364/A NOR2X1_LOC_73/a_36_216# 0.00fF
C40988 NOR2X1_LOC_791/Y INVX1_LOC_76/A 0.03fF
C40989 INVX1_LOC_249/Y INVX1_LOC_22/A 0.01fF
C40990 NAND2X1_LOC_733/Y NOR2X1_LOC_2/Y 0.14fF
C40991 INVX1_LOC_227/A INVX1_LOC_33/A 0.07fF
C40992 INVX1_LOC_36/A INVX1_LOC_73/A 0.06fF
C40993 INVX1_LOC_135/A NOR2X1_LOC_433/A 0.01fF
C40994 NOR2X1_LOC_662/A INVX1_LOC_15/A 0.05fF
C40995 NAND2X1_LOC_200/B NOR2X1_LOC_537/Y 0.09fF
C40996 NOR2X1_LOC_6/B NOR2X1_LOC_748/Y 0.05fF
C40997 INVX1_LOC_314/Y NOR2X1_LOC_749/Y 0.03fF
C40998 NOR2X1_LOC_128/a_36_216# INVX1_LOC_29/A 0.00fF
C40999 INVX1_LOC_135/A NOR2X1_LOC_474/A 0.07fF
C41000 NOR2X1_LOC_52/B NAND2X1_LOC_479/Y 0.03fF
C41001 NAND2X1_LOC_364/Y INVX1_LOC_148/Y 0.04fF
C41002 NOR2X1_LOC_237/Y NOR2X1_LOC_76/A 0.70fF
C41003 INVX1_LOC_136/A INVX1_LOC_75/A 0.15fF
C41004 NOR2X1_LOC_705/B INVX1_LOC_86/Y 0.02fF
C41005 NOR2X1_LOC_637/A NOR2X1_LOC_329/B 0.01fF
C41006 NAND2X1_LOC_326/A NAND2X1_LOC_655/B 0.07fF
C41007 INVX1_LOC_11/A NOR2X1_LOC_552/A 0.07fF
C41008 NOR2X1_LOC_437/Y NOR2X1_LOC_122/Y 0.11fF
C41009 INVX1_LOC_20/A NAND2X1_LOC_218/A 0.01fF
C41010 NOR2X1_LOC_38/B NAND2X1_LOC_219/B 0.01fF
C41011 INVX1_LOC_271/Y NOR2X1_LOC_666/a_36_216# 0.01fF
C41012 NAND2X1_LOC_819/Y INVX1_LOC_40/A 0.15fF
C41013 NOR2X1_LOC_137/A INVX1_LOC_155/Y 0.00fF
C41014 INVX1_LOC_30/A NOR2X1_LOC_167/Y 0.01fF
C41015 NAND2X1_LOC_116/A NOR2X1_LOC_199/B 0.00fF
C41016 INVX1_LOC_255/Y NOR2X1_LOC_655/B 0.12fF
C41017 INVX1_LOC_28/A NOR2X1_LOC_152/Y 0.24fF
C41018 NAND2X1_LOC_123/Y INVX1_LOC_71/A 0.01fF
C41019 NAND2X1_LOC_364/A NOR2X1_LOC_74/A 0.03fF
C41020 NAND2X1_LOC_338/B INVX1_LOC_137/A 0.10fF
C41021 INVX1_LOC_17/A NAND2X1_LOC_447/Y 0.01fF
C41022 INVX1_LOC_21/A NAND2X1_LOC_472/Y 0.07fF
C41023 INVX1_LOC_314/Y INVX1_LOC_102/Y 0.02fF
C41024 NOR2X1_LOC_88/Y INVX1_LOC_57/A 0.10fF
C41025 NAND2X1_LOC_538/Y INVX1_LOC_20/A 0.07fF
C41026 INVX1_LOC_135/A NOR2X1_LOC_52/B 0.11fF
C41027 NOR2X1_LOC_208/Y INVX1_LOC_73/A 0.00fF
C41028 D_INPUT_0 INVX1_LOC_60/Y 0.07fF
C41029 NOR2X1_LOC_474/A INVX1_LOC_169/Y 0.01fF
C41030 NAND2X1_LOC_364/A NOR2X1_LOC_9/Y 0.02fF
C41031 NOR2X1_LOC_134/a_36_216# NAND2X1_LOC_477/Y 0.01fF
C41032 INVX1_LOC_49/A NOR2X1_LOC_197/Y 0.01fF
C41033 NOR2X1_LOC_328/Y NOR2X1_LOC_447/a_36_216# 0.00fF
C41034 INVX1_LOC_211/Y NOR2X1_LOC_56/Y 0.03fF
C41035 NOR2X1_LOC_124/B INPUT_1 0.00fF
C41036 INVX1_LOC_89/A NAND2X1_LOC_122/a_36_24# 0.00fF
C41037 INVX1_LOC_33/A NOR2X1_LOC_703/A 0.01fF
C41038 INVX1_LOC_90/A INVX1_LOC_104/A 0.10fF
C41039 INVX1_LOC_171/A NOR2X1_LOC_709/A 0.01fF
C41040 NAND2X1_LOC_555/Y INVX1_LOC_74/Y 0.04fF
C41041 NOR2X1_LOC_590/A NOR2X1_LOC_486/Y 0.05fF
C41042 NAND2X1_LOC_430/B D_INPUT_5 0.01fF
C41043 INVX1_LOC_279/A NOR2X1_LOC_757/Y 0.22fF
C41044 INVX1_LOC_230/Y INVX1_LOC_59/Y 0.19fF
C41045 NOR2X1_LOC_389/B INVX1_LOC_104/A 0.18fF
C41046 INVX1_LOC_78/A INVX1_LOC_109/A 0.01fF
C41047 INVX1_LOC_230/Y INVX1_LOC_112/A 0.03fF
C41048 NOR2X1_LOC_530/Y INVX1_LOC_20/A 0.03fF
C41049 INVX1_LOC_312/Y NAND2X1_LOC_655/A 0.00fF
C41050 INVX1_LOC_84/A INVX1_LOC_57/A 0.14fF
C41051 INVX1_LOC_34/A NAND2X1_LOC_560/A 0.04fF
C41052 INVX1_LOC_11/A INVX1_LOC_139/Y 0.05fF
C41053 NOR2X1_LOC_195/A VDD -0.00fF
C41054 NOR2X1_LOC_250/Y NOR2X1_LOC_111/A 0.42fF
C41055 NOR2X1_LOC_251/a_36_216# INVX1_LOC_38/A 0.00fF
C41056 NOR2X1_LOC_617/Y INVX1_LOC_309/A 0.27fF
C41057 NAND2X1_LOC_88/a_36_24# NOR2X1_LOC_560/A 0.01fF
C41058 INVX1_LOC_211/Y VDD 0.03fF
C41059 NOR2X1_LOC_632/Y NOR2X1_LOC_665/A 0.01fF
C41060 NAND2X1_LOC_35/B INVX1_LOC_207/Y 0.01fF
C41061 NOR2X1_LOC_271/B NOR2X1_LOC_271/Y 0.06fF
C41062 INVX1_LOC_243/Y NAND2X1_LOC_651/B 0.26fF
C41063 NOR2X1_LOC_309/Y INVX1_LOC_73/A 0.03fF
C41064 INVX1_LOC_177/A NOR2X1_LOC_564/Y 0.01fF
C41065 NOR2X1_LOC_202/Y NOR2X1_LOC_52/B 0.13fF
C41066 INVX1_LOC_41/Y INVX1_LOC_91/A 0.03fF
C41067 NOR2X1_LOC_569/Y NOR2X1_LOC_565/B 0.02fF
C41068 NAND2X1_LOC_803/B NOR2X1_LOC_816/Y 0.02fF
C41069 INVX1_LOC_256/A INVX1_LOC_281/A 0.02fF
C41070 NAND2X1_LOC_564/B NOR2X1_LOC_130/A 0.03fF
C41071 INVX1_LOC_30/A INVX1_LOC_76/A 0.17fF
C41072 INVX1_LOC_105/A NOR2X1_LOC_7/Y 0.01fF
C41073 INVX1_LOC_197/Y NAND2X1_LOC_622/a_36_24# 0.00fF
C41074 NAND2X1_LOC_308/Y INPUT_0 0.07fF
C41075 NAND2X1_LOC_9/Y NOR2X1_LOC_721/B 0.04fF
C41076 NOR2X1_LOC_843/B NAND2X1_LOC_206/B 0.03fF
C41077 INVX1_LOC_11/A INVX1_LOC_280/A 0.07fF
C41078 INVX1_LOC_278/A NOR2X1_LOC_662/A 0.10fF
C41079 NAND2X1_LOC_192/a_36_24# NOR2X1_LOC_331/B 0.00fF
C41080 NOR2X1_LOC_246/a_36_216# INVX1_LOC_53/Y 0.00fF
C41081 NOR2X1_LOC_646/A INPUT_1 0.04fF
C41082 NOR2X1_LOC_718/B INVX1_LOC_311/A 0.89fF
C41083 NOR2X1_LOC_394/Y NOR2X1_LOC_38/B 0.14fF
C41084 NOR2X1_LOC_554/B NOR2X1_LOC_35/Y 0.10fF
C41085 NOR2X1_LOC_441/Y NAND2X1_LOC_284/a_36_24# 0.00fF
C41086 INVX1_LOC_31/A INVX1_LOC_117/A 0.07fF
C41087 NAND2X1_LOC_785/A NOR2X1_LOC_74/A 0.02fF
C41088 INVX1_LOC_71/A NOR2X1_LOC_657/B 0.07fF
C41089 INVX1_LOC_136/A NAND2X1_LOC_453/A 0.10fF
C41090 INVX1_LOC_182/Y NOR2X1_LOC_757/Y 0.01fF
C41091 INVX1_LOC_93/A INVX1_LOC_119/Y 0.06fF
C41092 NAND2X1_LOC_374/Y INVX1_LOC_282/A 0.07fF
C41093 NAND2X1_LOC_35/Y INVX1_LOC_19/A 0.07fF
C41094 INVX1_LOC_224/Y INVX1_LOC_170/Y 0.01fF
C41095 NOR2X1_LOC_593/Y NOR2X1_LOC_552/A 0.02fF
C41096 NOR2X1_LOC_759/A VDD 0.02fF
C41097 NOR2X1_LOC_828/A INVX1_LOC_279/A 0.04fF
C41098 NOR2X1_LOC_92/Y NOR2X1_LOC_841/A 0.74fF
C41099 NOR2X1_LOC_846/Y INVX1_LOC_63/A 0.46fF
C41100 NAND2X1_LOC_189/a_36_24# NAND2X1_LOC_656/Y 0.01fF
C41101 INVX1_LOC_63/Y NOR2X1_LOC_43/Y 0.01fF
C41102 INVX1_LOC_21/A NAND2X1_LOC_206/Y 0.07fF
C41103 INVX1_LOC_142/A NOR2X1_LOC_698/Y 0.26fF
C41104 INVX1_LOC_255/Y NOR2X1_LOC_381/a_36_216# 0.00fF
C41105 NAND2X1_LOC_554/a_36_24# NOR2X1_LOC_473/B 0.00fF
C41106 INVX1_LOC_290/A INVX1_LOC_140/A 0.03fF
C41107 INVX1_LOC_239/Y NAND2X1_LOC_463/B 0.01fF
C41108 NOR2X1_LOC_468/Y NAND2X1_LOC_572/B 0.07fF
C41109 INVX1_LOC_83/A INVX1_LOC_85/Y 0.97fF
C41110 INVX1_LOC_57/A INVX1_LOC_15/A 0.17fF
C41111 INVX1_LOC_103/A NOR2X1_LOC_832/a_36_216# 0.00fF
C41112 INVX1_LOC_275/A NOR2X1_LOC_683/Y 0.01fF
C41113 NAND2X1_LOC_181/Y INVX1_LOC_6/A 0.03fF
C41114 INVX1_LOC_23/A INVX1_LOC_3/Y 0.24fF
C41115 NAND2X1_LOC_28/a_36_24# INVX1_LOC_89/A 0.00fF
C41116 INVX1_LOC_24/A NAND2X1_LOC_804/Y 0.01fF
C41117 INVX1_LOC_13/A NOR2X1_LOC_721/Y 0.00fF
C41118 INVX1_LOC_28/A NAND2X1_LOC_861/Y 0.07fF
C41119 INVX1_LOC_229/Y NAND2X1_LOC_863/A 0.14fF
C41120 NOR2X1_LOC_717/B INVX1_LOC_182/Y 0.00fF
C41121 NOR2X1_LOC_478/A INVX1_LOC_92/A 0.04fF
C41122 NAND2X1_LOC_181/Y NOR2X1_LOC_10/a_36_216# 0.00fF
C41123 INVX1_LOC_89/A NAND2X1_LOC_7/a_36_24# 0.00fF
C41124 D_GATE_366 NOR2X1_LOC_156/A 0.01fF
C41125 NOR2X1_LOC_593/Y INVX1_LOC_139/Y 0.01fF
C41126 NOR2X1_LOC_419/Y NOR2X1_LOC_98/B 0.01fF
C41127 INVX1_LOC_162/Y NAND2X1_LOC_287/B 0.02fF
C41128 NOR2X1_LOC_644/A INVX1_LOC_182/A 0.01fF
C41129 INVX1_LOC_82/Y INPUT_1 0.01fF
C41130 INVX1_LOC_53/A NAND2X1_LOC_454/Y 0.06fF
C41131 NOR2X1_LOC_709/A INVX1_LOC_20/A 1.06fF
C41132 INVX1_LOC_16/Y NAND2X1_LOC_215/A 0.02fF
C41133 INVX1_LOC_5/A NOR2X1_LOC_467/A 0.02fF
C41134 NOR2X1_LOC_270/Y NAND2X1_LOC_93/B 0.07fF
C41135 NAND2X1_LOC_722/A INVX1_LOC_76/A 0.07fF
C41136 NOR2X1_LOC_721/A NOR2X1_LOC_35/Y 0.06fF
C41137 INVX1_LOC_72/A NOR2X1_LOC_216/B 0.10fF
C41138 INVX1_LOC_1/A NAND2X1_LOC_83/a_36_24# 0.00fF
C41139 NOR2X1_LOC_68/A INVX1_LOC_92/A 0.30fF
C41140 INVX1_LOC_48/Y INVX1_LOC_42/A 0.04fF
C41141 INVX1_LOC_58/A NOR2X1_LOC_91/A 0.31fF
C41142 INVX1_LOC_2/A INVX1_LOC_2/Y 0.23fF
C41143 D_INPUT_4 NOR2X1_LOC_163/a_36_216# 0.00fF
C41144 INVX1_LOC_236/A VDD 0.36fF
C41145 NOR2X1_LOC_81/Y INVX1_LOC_4/A 0.03fF
C41146 INVX1_LOC_272/Y INVX1_LOC_12/A 0.12fF
C41147 NOR2X1_LOC_360/Y NOR2X1_LOC_831/B 0.10fF
C41148 VDD INVX1_LOC_210/A 0.12fF
C41149 INVX1_LOC_276/A NOR2X1_LOC_681/Y 0.01fF
C41150 INVX1_LOC_276/A INVX1_LOC_37/A 0.07fF
C41151 INVX1_LOC_30/Y NOR2X1_LOC_80/a_36_216# 0.00fF
C41152 NOR2X1_LOC_52/B NOR2X1_LOC_152/A 0.00fF
C41153 NAND2X1_LOC_53/Y INVX1_LOC_12/A 0.26fF
C41154 NAND2X1_LOC_205/A NAND2X1_LOC_215/A 0.16fF
C41155 INVX1_LOC_174/A NAND2X1_LOC_259/a_36_24# 0.01fF
C41156 INVX1_LOC_35/A NOR2X1_LOC_647/A 0.06fF
C41157 INVX1_LOC_49/A INVX1_LOC_307/Y 0.00fF
C41158 NAND2X1_LOC_656/Y NOR2X1_LOC_139/Y 0.25fF
C41159 INVX1_LOC_104/A INVX1_LOC_38/A 0.07fF
C41160 INVX1_LOC_58/A INVX1_LOC_23/A 0.21fF
C41161 NOR2X1_LOC_52/B INVX1_LOC_280/A 0.01fF
C41162 INVX1_LOC_15/A NOR2X1_LOC_475/A 0.07fF
C41163 NOR2X1_LOC_391/A INVX1_LOC_95/Y 0.07fF
C41164 NOR2X1_LOC_749/Y NOR2X1_LOC_557/A 0.01fF
C41165 NOR2X1_LOC_666/Y INVX1_LOC_15/A 0.00fF
C41166 NOR2X1_LOC_172/a_36_216# NOR2X1_LOC_536/A 0.02fF
C41167 NOR2X1_LOC_103/Y INVX1_LOC_170/Y 0.00fF
C41168 INVX1_LOC_278/A INVX1_LOC_57/A 0.14fF
C41169 INVX1_LOC_225/A NOR2X1_LOC_612/Y 0.02fF
C41170 NOR2X1_LOC_392/Y NOR2X1_LOC_414/Y 0.02fF
C41171 NOR2X1_LOC_92/Y INVX1_LOC_128/A 0.18fF
C41172 NOR2X1_LOC_473/B NOR2X1_LOC_318/B -0.03fF
C41173 NAND2X1_LOC_347/B INVX1_LOC_4/Y 0.01fF
C41174 NAND2X1_LOC_656/Y NAND2X1_LOC_468/B 0.02fF
C41175 NOR2X1_LOC_667/A NAND2X1_LOC_603/a_36_24# 0.00fF
C41176 NAND2X1_LOC_804/A NAND2X1_LOC_794/a_36_24# 0.02fF
C41177 NAND2X1_LOC_866/B NAND2X1_LOC_623/B 0.03fF
C41178 NOR2X1_LOC_489/a_36_216# INVX1_LOC_57/A 0.00fF
C41179 NAND2X1_LOC_9/Y NAND2X1_LOC_860/A 0.09fF
C41180 INVX1_LOC_13/A VDD 0.96fF
C41181 INVX1_LOC_90/A NOR2X1_LOC_600/Y 0.52fF
C41182 NOR2X1_LOC_433/A NOR2X1_LOC_473/a_36_216# 0.01fF
C41183 INVX1_LOC_135/A INVX1_LOC_74/A 0.12fF
C41184 NOR2X1_LOC_218/Y NOR2X1_LOC_363/Y 0.21fF
C41185 INVX1_LOC_233/A NAND2X1_LOC_860/A 0.39fF
C41186 NOR2X1_LOC_808/A NOR2X1_LOC_729/A 0.03fF
C41187 INVX1_LOC_110/Y NOR2X1_LOC_861/Y 0.93fF
C41188 NOR2X1_LOC_273/Y INVX1_LOC_186/Y 0.01fF
C41189 INVX1_LOC_202/A NAND2X1_LOC_476/Y 0.01fF
C41190 INVX1_LOC_90/A NAND2X1_LOC_674/a_36_24# 0.00fF
C41191 INVX1_LOC_25/A INVX1_LOC_5/A 0.80fF
C41192 NOR2X1_LOC_657/Y INVX1_LOC_109/Y 0.03fF
C41193 NOR2X1_LOC_759/Y INVX1_LOC_186/Y 0.00fF
C41194 NOR2X1_LOC_792/B NOR2X1_LOC_831/B 0.02fF
C41195 NOR2X1_LOC_564/Y INVX1_LOC_65/A 0.03fF
C41196 NOR2X1_LOC_742/A NOR2X1_LOC_562/B 0.20fF
C41197 INVX1_LOC_247/Y INVX1_LOC_99/A 0.01fF
C41198 INVX1_LOC_34/A NAND2X1_LOC_606/a_36_24# 0.01fF
C41199 INVX1_LOC_31/A INVX1_LOC_3/Y 0.75fF
C41200 NOR2X1_LOC_454/Y NOR2X1_LOC_638/Y 0.05fF
C41201 INVX1_LOC_224/Y INVX1_LOC_27/A 0.06fF
C41202 INVX1_LOC_266/Y NOR2X1_LOC_155/A 0.12fF
C41203 NAND2X1_LOC_579/A NOR2X1_LOC_693/Y 0.10fF
C41204 NAND2X1_LOC_214/B NAND2X1_LOC_415/a_36_24# 0.00fF
C41205 NOR2X1_LOC_246/A VDD 0.00fF
C41206 NAND2X1_LOC_370/a_36_24# NAND2X1_LOC_552/A 0.01fF
C41207 D_INPUT_0 NOR2X1_LOC_111/A 0.20fF
C41208 NOR2X1_LOC_550/B INVX1_LOC_186/Y 0.10fF
C41209 NAND2X1_LOC_477/A NOR2X1_LOC_841/A 0.12fF
C41210 NOR2X1_LOC_639/a_36_216# INVX1_LOC_77/Y 0.01fF
C41211 NOR2X1_LOC_174/B VDD 0.34fF
C41212 INVX1_LOC_50/A NAND2X1_LOC_705/Y 0.00fF
C41213 INVX1_LOC_182/A NOR2X1_LOC_540/B 0.01fF
C41214 INVX1_LOC_2/Y INPUT_1 0.00fF
C41215 NOR2X1_LOC_810/A INVX1_LOC_299/Y 0.09fF
C41216 NOR2X1_LOC_798/A NOR2X1_LOC_211/a_36_216# 0.00fF
C41217 INVX1_LOC_36/A NAND2X1_LOC_404/a_36_24# 0.00fF
C41218 NAND2X1_LOC_338/B NOR2X1_LOC_216/B 0.03fF
C41219 INVX1_LOC_27/A NAND2X1_LOC_38/a_36_24# 0.02fF
C41220 INVX1_LOC_246/A INVX1_LOC_78/A 0.15fF
C41221 NAND2X1_LOC_634/a_36_24# NAND2X1_LOC_464/B 0.01fF
C41222 INVX1_LOC_207/Y VDD -0.00fF
C41223 NOR2X1_LOC_405/A NOR2X1_LOC_74/A 6.15fF
C41224 NOR2X1_LOC_516/B NOR2X1_LOC_61/Y 0.10fF
C41225 INVX1_LOC_55/Y VDD 0.18fF
C41226 INVX1_LOC_50/A NAND2X1_LOC_303/Y 0.18fF
C41227 NOR2X1_LOC_798/A NOR2X1_LOC_634/Y 0.00fF
C41228 NOR2X1_LOC_152/Y INVX1_LOC_109/A 0.01fF
C41229 NOR2X1_LOC_644/B INVX1_LOC_271/Y 0.04fF
C41230 NAND2X1_LOC_575/a_36_24# NOR2X1_LOC_654/A 0.00fF
C41231 NOR2X1_LOC_577/Y NAND2X1_LOC_74/B 0.07fF
C41232 NAND2X1_LOC_521/a_36_24# NOR2X1_LOC_861/Y 0.00fF
C41233 INVX1_LOC_215/A INVX1_LOC_54/A 0.02fF
C41234 NOR2X1_LOC_112/B NOR2X1_LOC_332/B 0.00fF
C41235 NAND2X1_LOC_623/B INVX1_LOC_6/A 0.01fF
C41236 NOR2X1_LOC_78/B NOR2X1_LOC_49/a_36_216# 0.00fF
C41237 NOR2X1_LOC_405/A NOR2X1_LOC_9/Y 0.21fF
C41238 NOR2X1_LOC_636/B INVX1_LOC_296/A 0.31fF
C41239 INVX1_LOC_16/A NAND2X1_LOC_802/Y 0.07fF
C41240 INVX1_LOC_249/Y INVX1_LOC_186/Y 0.02fF
C41241 NOR2X1_LOC_828/Y INVX1_LOC_1/A 0.07fF
C41242 INVX1_LOC_159/A INVX1_LOC_32/A 0.02fF
C41243 NOR2X1_LOC_91/A INVX1_LOC_215/Y 0.00fF
C41244 NOR2X1_LOC_318/B NOR2X1_LOC_355/B 0.07fF
C41245 NOR2X1_LOC_500/Y NOR2X1_LOC_445/B 0.00fF
C41246 INVX1_LOC_35/A NOR2X1_LOC_321/Y 0.07fF
C41247 INVX1_LOC_286/Y NAND2X1_LOC_175/Y 0.17fF
C41248 INVX1_LOC_166/A NAND2X1_LOC_377/a_36_24# 0.01fF
C41249 INVX1_LOC_34/A INVX1_LOC_29/A 0.16fF
C41250 NOR2X1_LOC_763/a_36_216# NOR2X1_LOC_48/B 0.00fF
C41251 INVX1_LOC_286/A INVX1_LOC_95/A 0.01fF
C41252 NAND2X1_LOC_656/A INVX1_LOC_47/Y 0.23fF
C41253 INVX1_LOC_101/Y NOR2X1_LOC_717/A 0.00fF
C41254 NOR2X1_LOC_738/Y INVX1_LOC_23/A 0.01fF
C41255 INVX1_LOC_159/A NOR2X1_LOC_329/Y 0.08fF
C41256 NOR2X1_LOC_52/Y NAND2X1_LOC_470/B 0.11fF
C41257 INVX1_LOC_164/Y INVX1_LOC_63/A 0.08fF
C41258 NOR2X1_LOC_322/Y NAND2X1_LOC_721/A 0.08fF
C41259 INVX1_LOC_10/A INVX1_LOC_307/A 0.07fF
C41260 INVX1_LOC_33/A NOR2X1_LOC_169/a_36_216# 0.00fF
C41261 NOR2X1_LOC_320/Y VDD 0.12fF
C41262 NOR2X1_LOC_590/A NOR2X1_LOC_748/A 0.05fF
C41263 INVX1_LOC_298/Y NOR2X1_LOC_722/Y 0.01fF
C41264 NOR2X1_LOC_9/Y NOR2X1_LOC_857/A 0.01fF
C41265 NOR2X1_LOC_99/B NOR2X1_LOC_61/A 0.04fF
C41266 INVX1_LOC_5/A INVX1_LOC_1/A 0.20fF
C41267 INVX1_LOC_205/Y NOR2X1_LOC_249/Y 0.01fF
C41268 NOR2X1_LOC_742/A INVX1_LOC_281/Y 0.01fF
C41269 NOR2X1_LOC_419/Y NOR2X1_LOC_38/B 0.16fF
C41270 INVX1_LOC_35/A NAND2X1_LOC_793/Y 0.03fF
C41271 INVX1_LOC_58/A INVX1_LOC_31/A 0.13fF
C41272 NAND2X1_LOC_231/Y INVX1_LOC_29/A 0.77fF
C41273 NAND2X1_LOC_741/B INVX1_LOC_296/A 0.03fF
C41274 INVX1_LOC_251/Y NOR2X1_LOC_89/A 0.12fF
C41275 NOR2X1_LOC_160/B NOR2X1_LOC_678/A 3.01fF
C41276 NOR2X1_LOC_346/B NAND2X1_LOC_74/B 0.15fF
C41277 INVX1_LOC_45/A INVX1_LOC_271/A 0.03fF
C41278 NOR2X1_LOC_84/Y INVX1_LOC_42/A 0.20fF
C41279 INVX1_LOC_64/A NOR2X1_LOC_530/Y 0.00fF
C41280 NOR2X1_LOC_163/A INVX1_LOC_92/A 0.01fF
C41281 INVX1_LOC_6/A INVX1_LOC_117/A 1.70fF
C41282 NOR2X1_LOC_482/Y INVX1_LOC_42/A 0.39fF
C41283 INVX1_LOC_28/A INVX1_LOC_291/A 0.07fF
C41284 INVX1_LOC_40/A NOR2X1_LOC_77/a_36_216# 0.00fF
C41285 INVX1_LOC_5/A NOR2X1_LOC_794/B 0.03fF
C41286 NOR2X1_LOC_757/a_36_216# INVX1_LOC_290/Y 0.01fF
C41287 INVX1_LOC_77/A NOR2X1_LOC_278/Y 0.02fF
C41288 INVX1_LOC_17/A NAND2X1_LOC_796/B 0.07fF
C41289 INVX1_LOC_22/A NAND2X1_LOC_74/B 0.05fF
C41290 INVX1_LOC_226/Y INVX1_LOC_12/A 0.03fF
C41291 INVX1_LOC_150/A NOR2X1_LOC_814/A 0.02fF
C41292 NOR2X1_LOC_329/B NAND2X1_LOC_798/B 0.07fF
C41293 INVX1_LOC_27/A NOR2X1_LOC_103/Y 0.14fF
C41294 NAND2X1_LOC_451/Y NAND2X1_LOC_430/B 0.33fF
C41295 INVX1_LOC_211/Y NOR2X1_LOC_510/Y 0.16fF
C41296 INVX1_LOC_206/Y INVX1_LOC_38/A 0.03fF
C41297 NAND2X1_LOC_714/B NAND2X1_LOC_799/A 0.00fF
C41298 NOR2X1_LOC_338/Y INVX1_LOC_23/A 0.01fF
C41299 NAND2X1_LOC_812/A NOR2X1_LOC_829/A 0.02fF
C41300 INVX1_LOC_171/A INVX1_LOC_294/A 0.03fF
C41301 NOR2X1_LOC_709/A INVX1_LOC_4/A 1.52fF
C41302 INVX1_LOC_83/A NAND2X1_LOC_782/B 0.07fF
C41303 INVX1_LOC_239/Y INVX1_LOC_42/A 0.01fF
C41304 INVX1_LOC_89/A NOR2X1_LOC_814/A 0.31fF
C41305 NOR2X1_LOC_593/Y NOR2X1_LOC_541/B 0.06fF
C41306 NOR2X1_LOC_68/A INVX1_LOC_53/A 0.62fF
C41307 INVX1_LOC_80/A NAND2X1_LOC_82/Y 0.03fF
C41308 INVX1_LOC_50/A NOR2X1_LOC_106/Y 0.16fF
C41309 INVX1_LOC_298/Y INVX1_LOC_34/A 0.03fF
C41310 INVX1_LOC_71/A INVX1_LOC_271/A 0.68fF
C41311 INVX1_LOC_77/A NOR2X1_LOC_844/a_36_216# 0.01fF
C41312 NOR2X1_LOC_305/a_36_216# NOR2X1_LOC_305/Y 0.00fF
C41313 NOR2X1_LOC_262/Y INVX1_LOC_57/A 0.03fF
C41314 INPUT_0 INVX1_LOC_152/A 0.01fF
C41315 INVX1_LOC_42/Y NOR2X1_LOC_155/A 0.03fF
C41316 INVX1_LOC_45/A NAND2X1_LOC_214/B 0.00fF
C41317 NAND2X1_LOC_796/a_36_24# NOR2X1_LOC_186/Y 0.00fF
C41318 NOR2X1_LOC_180/B INVX1_LOC_63/A 0.07fF
C41319 INVX1_LOC_286/A INVX1_LOC_54/A 0.02fF
C41320 NAND2X1_LOC_222/B NAND2X1_LOC_219/a_36_24# 0.02fF
C41321 INPUT_0 NOR2X1_LOC_634/A 0.20fF
C41322 NAND2X1_LOC_508/A NOR2X1_LOC_814/A 0.02fF
C41323 INVX1_LOC_10/A INVX1_LOC_12/A 4.44fF
C41324 NOR2X1_LOC_357/Y NOR2X1_LOC_69/a_36_216# 0.01fF
C41325 NOR2X1_LOC_272/Y INVX1_LOC_124/Y 0.34fF
C41326 NOR2X1_LOC_357/Y VDD 1.40fF
C41327 NOR2X1_LOC_600/Y INVX1_LOC_38/A 0.00fF
C41328 INVX1_LOC_173/Y NOR2X1_LOC_36/B 0.06fF
C41329 INVX1_LOC_187/A NAND2X1_LOC_446/a_36_24# 0.02fF
C41330 INVX1_LOC_155/Y NOR2X1_LOC_383/B 0.00fF
C41331 NOR2X1_LOC_482/Y INVX1_LOC_78/A 0.13fF
C41332 NOR2X1_LOC_315/Y INVX1_LOC_23/Y 0.00fF
C41333 NAND2X1_LOC_218/B NOR2X1_LOC_660/Y 0.03fF
C41334 INVX1_LOC_45/A INVX1_LOC_27/A 0.03fF
C41335 NOR2X1_LOC_690/A INVX1_LOC_50/A 0.03fF
C41336 INVX1_LOC_204/A INVX1_LOC_34/A 0.01fF
C41337 NOR2X1_LOC_504/a_36_216# INVX1_LOC_12/A 0.00fF
C41338 INVX1_LOC_148/A NOR2X1_LOC_691/B 0.00fF
C41339 NOR2X1_LOC_598/B NOR2X1_LOC_643/Y 0.02fF
C41340 NOR2X1_LOC_78/B NAND2X1_LOC_454/Y 0.16fF
C41341 NAND2X1_LOC_859/Y INVX1_LOC_3/Y 0.13fF
C41342 NOR2X1_LOC_32/B NAND2X1_LOC_632/B 0.05fF
C41343 INVX1_LOC_185/A INVX1_LOC_91/A 0.03fF
C41344 INVX1_LOC_135/A NAND2X1_LOC_254/Y 0.03fF
C41345 INVX1_LOC_255/Y NOR2X1_LOC_28/a_36_216# 0.01fF
C41346 NAND2X1_LOC_852/Y NOR2X1_LOC_409/B 0.01fF
C41347 INVX1_LOC_178/A NOR2X1_LOC_384/Y 0.03fF
C41348 INVX1_LOC_39/A NOR2X1_LOC_791/B 0.04fF
C41349 INVX1_LOC_74/A INVX1_LOC_280/A 0.04fF
C41350 INVX1_LOC_95/A INVX1_LOC_54/A 0.01fF
C41351 VDD NOR2X1_LOC_319/B 0.31fF
C41352 NOR2X1_LOC_710/B NAND2X1_LOC_701/a_36_24# 0.00fF
C41353 INVX1_LOC_266/A INVX1_LOC_223/A 0.02fF
C41354 VDD INVX1_LOC_66/Y 0.73fF
C41355 INVX1_LOC_11/Y INVX1_LOC_185/A 0.06fF
C41356 INVX1_LOC_35/A NOR2X1_LOC_379/a_36_216# 0.00fF
C41357 VDD NOR2X1_LOC_692/Y 0.26fF
C41358 NOR2X1_LOC_589/A NOR2X1_LOC_334/Y 0.07fF
C41359 NOR2X1_LOC_75/Y NOR2X1_LOC_389/A 0.01fF
C41360 INVX1_LOC_21/A INVX1_LOC_24/A 0.21fF
C41361 NOR2X1_LOC_16/Y INVX1_LOC_57/A 0.03fF
C41362 NOR2X1_LOC_203/a_36_216# NOR2X1_LOC_577/Y 0.01fF
C41363 NAND2X1_LOC_804/Y NAND2X1_LOC_811/B 0.04fF
C41364 INVX1_LOC_290/A INVX1_LOC_78/A 0.04fF
C41365 NOR2X1_LOC_111/A NAND2X1_LOC_848/A 0.10fF
C41366 NAND2X1_LOC_513/B INVX1_LOC_198/Y 0.01fF
C41367 NOR2X1_LOC_644/A NOR2X1_LOC_850/B 0.01fF
C41368 INVX1_LOC_144/A INVX1_LOC_19/A 0.07fF
C41369 INVX1_LOC_27/A INVX1_LOC_71/A 0.41fF
C41370 INVX1_LOC_215/Y INVX1_LOC_31/A 0.41fF
C41371 NAND2X1_LOC_796/B NAND2X1_LOC_547/a_36_24# 0.01fF
C41372 NAND2X1_LOC_725/A NAND2X1_LOC_811/Y 0.05fF
C41373 INVX1_LOC_58/A INVX1_LOC_191/Y 0.01fF
C41374 NOR2X1_LOC_420/Y NOR2X1_LOC_716/B 0.08fF
C41375 INVX1_LOC_11/A NAND2X1_LOC_387/B 0.03fF
C41376 INVX1_LOC_37/A NOR2X1_LOC_729/A 0.00fF
C41377 NOR2X1_LOC_226/A INVX1_LOC_29/Y 0.01fF
C41378 NAND2X1_LOC_763/a_36_24# NAND2X1_LOC_451/Y 0.00fF
C41379 INPUT_0 INVX1_LOC_29/A 2.20fF
C41380 NOR2X1_LOC_68/A NAND2X1_LOC_522/a_36_24# 0.01fF
C41381 INVX1_LOC_288/Y INVX1_LOC_22/A 0.01fF
C41382 NOR2X1_LOC_124/A INVX1_LOC_123/Y 0.02fF
C41383 INVX1_LOC_288/A INVX1_LOC_290/A 0.01fF
C41384 INVX1_LOC_256/A NOR2X1_LOC_52/Y 0.15fF
C41385 INVX1_LOC_25/A NOR2X1_LOC_773/Y 0.02fF
C41386 NOR2X1_LOC_487/Y INVX1_LOC_46/A 0.02fF
C41387 INVX1_LOC_37/Y INVX1_LOC_118/A 0.05fF
C41388 NOR2X1_LOC_130/Y NOR2X1_LOC_38/B 0.00fF
C41389 INVX1_LOC_100/A NAND2X1_LOC_74/B 0.04fF
C41390 NOR2X1_LOC_218/a_36_216# INVX1_LOC_290/Y 0.00fF
C41391 INVX1_LOC_256/A NOR2X1_LOC_270/Y 0.15fF
C41392 NOR2X1_LOC_35/Y NAND2X1_LOC_255/a_36_24# 0.07fF
C41393 INVX1_LOC_28/A NOR2X1_LOC_609/Y 0.01fF
C41394 D_INPUT_1 INVX1_LOC_316/Y 0.08fF
C41395 NAND2X1_LOC_651/a_36_24# NOR2X1_LOC_467/A 0.01fF
C41396 INVX1_LOC_224/Y INVX1_LOC_137/A 0.00fF
C41397 NOR2X1_LOC_637/B NAND2X1_LOC_175/a_36_24# 0.00fF
C41398 NOR2X1_LOC_220/A INVX1_LOC_58/Y 0.10fF
C41399 INVX1_LOC_305/A NOR2X1_LOC_160/B 0.08fF
C41400 INVX1_LOC_39/A NOR2X1_LOC_124/B 0.01fF
C41401 VDD INVX1_LOC_260/A -0.00fF
C41402 NOR2X1_LOC_626/Y NOR2X1_LOC_718/B 0.06fF
C41403 NOR2X1_LOC_92/Y NOR2X1_LOC_172/Y 0.13fF
C41404 NOR2X1_LOC_251/a_36_216# INVX1_LOC_33/A -0.00fF
C41405 NAND2X1_LOC_624/B NAND2X1_LOC_374/Y 0.02fF
C41406 NOR2X1_LOC_99/B INVX1_LOC_16/Y 0.31fF
C41407 NOR2X1_LOC_468/Y NOR2X1_LOC_716/B 0.09fF
C41408 INVX1_LOC_178/A INVX1_LOC_221/A 0.01fF
C41409 NOR2X1_LOC_75/Y NOR2X1_LOC_596/A 0.08fF
C41410 INVX1_LOC_208/A NOR2X1_LOC_678/A 0.05fF
C41411 NOR2X1_LOC_763/Y NOR2X1_LOC_635/B 0.07fF
C41412 INVX1_LOC_58/A NAND2X1_LOC_859/Y 0.19fF
C41413 NOR2X1_LOC_516/B NOR2X1_LOC_678/A 0.00fF
C41414 NOR2X1_LOC_510/Y INVX1_LOC_236/A 0.26fF
C41415 NOR2X1_LOC_570/Y INVX1_LOC_53/A 0.03fF
C41416 INVX1_LOC_75/A NAND2X1_LOC_647/B 0.06fF
C41417 INVX1_LOC_266/A INVX1_LOC_149/Y 0.02fF
C41418 NOR2X1_LOC_646/a_36_216# NOR2X1_LOC_392/Y 0.00fF
C41419 NOR2X1_LOC_45/B NOR2X1_LOC_89/A 0.22fF
C41420 INVX1_LOC_136/A NOR2X1_LOC_274/B 0.10fF
C41421 INVX1_LOC_21/A INVX1_LOC_143/A 0.07fF
C41422 INVX1_LOC_25/A NOR2X1_LOC_332/A 0.21fF
C41423 INVX1_LOC_219/Y INVX1_LOC_14/A 0.00fF
C41424 VDD NAND2X1_LOC_489/Y 0.62fF
C41425 INVX1_LOC_95/A NAND2X1_LOC_807/B 0.23fF
C41426 INVX1_LOC_174/A NOR2X1_LOC_162/Y 0.01fF
C41427 NOR2X1_LOC_274/Y INVX1_LOC_30/A 0.03fF
C41428 INPUT_1 INVX1_LOC_29/Y 0.00fF
C41429 NOR2X1_LOC_273/Y INVX1_LOC_18/A 0.15fF
C41430 INVX1_LOC_24/A NAND2X1_LOC_354/Y 0.01fF
C41431 INVX1_LOC_269/A INVX1_LOC_196/A 0.10fF
C41432 NAND2X1_LOC_728/Y INVX1_LOC_300/Y 0.27fF
C41433 INVX1_LOC_292/A NOR2X1_LOC_390/a_36_216# 0.00fF
C41434 NOR2X1_LOC_284/B INVX1_LOC_299/A 0.01fF
C41435 INVX1_LOC_92/Y INVX1_LOC_87/A 0.14fF
C41436 INPUT_2 NOR2X1_LOC_6/B 0.10fF
C41437 INVX1_LOC_224/Y NOR2X1_LOC_19/B 0.00fF
C41438 NOR2X1_LOC_163/A INVX1_LOC_53/A 0.04fF
C41439 INVX1_LOC_64/A NOR2X1_LOC_106/A 0.05fF
C41440 INVX1_LOC_58/A NAND2X1_LOC_807/Y -0.02fF
C41441 INVX1_LOC_1/A NOR2X1_LOC_773/Y 0.12fF
C41442 INVX1_LOC_245/A NAND2X1_LOC_149/Y 0.04fF
C41443 NAND2X1_LOC_208/B INVX1_LOC_8/A 0.03fF
C41444 INVX1_LOC_136/A NOR2X1_LOC_577/Y 0.35fF
C41445 NAND2X1_LOC_53/Y NAND2X1_LOC_832/a_36_24# 0.01fF
C41446 INVX1_LOC_18/A NOR2X1_LOC_550/B 0.01fF
C41447 INVX1_LOC_119/A NOR2X1_LOC_590/A 0.60fF
C41448 INVX1_LOC_117/A INVX1_LOC_301/A 0.02fF
C41449 INVX1_LOC_118/A NOR2X1_LOC_485/Y 0.02fF
C41450 NOR2X1_LOC_584/Y INVX1_LOC_37/A 0.03fF
C41451 NOR2X1_LOC_419/Y INVX1_LOC_62/Y 0.79fF
C41452 NOR2X1_LOC_56/Y INVX1_LOC_32/A 0.07fF
C41453 INVX1_LOC_79/A INVX1_LOC_270/Y 0.02fF
C41454 NOR2X1_LOC_829/Y INPUT_0 0.03fF
C41455 INVX1_LOC_299/A INVX1_LOC_232/A 0.01fF
C41456 NAND2X1_LOC_200/B NOR2X1_LOC_103/Y 0.13fF
C41457 INVX1_LOC_21/A NAND2X1_LOC_783/A 0.11fF
C41458 NOR2X1_LOC_352/a_36_216# INVX1_LOC_271/Y 0.01fF
C41459 INVX1_LOC_99/Y INVX1_LOC_313/Y 0.01fF
C41460 NOR2X1_LOC_590/A NOR2X1_LOC_493/B 0.10fF
C41461 NOR2X1_LOC_155/A NAND2X1_LOC_288/A 0.09fF
C41462 INVX1_LOC_21/A NOR2X1_LOC_130/A 0.09fF
C41463 NOR2X1_LOC_136/Y INVX1_LOC_161/Y 0.04fF
C41464 INVX1_LOC_27/A NOR2X1_LOC_123/B 0.10fF
C41465 NAND2X1_LOC_787/A NOR2X1_LOC_716/a_36_216# 0.00fF
C41466 NOR2X1_LOC_819/a_36_216# NOR2X1_LOC_664/Y 0.00fF
C41467 NAND2X1_LOC_562/B NOR2X1_LOC_384/Y 0.01fF
C41468 INVX1_LOC_45/A INVX1_LOC_206/A 0.08fF
C41469 INVX1_LOC_136/A NOR2X1_LOC_348/B 0.07fF
C41470 NOR2X1_LOC_845/A INVX1_LOC_26/Y 0.01fF
C41471 NAND2X1_LOC_468/B INVX1_LOC_128/Y 0.00fF
C41472 NOR2X1_LOC_813/Y NAND2X1_LOC_254/Y 0.08fF
C41473 NOR2X1_LOC_103/Y INVX1_LOC_137/A 0.00fF
C41474 VDD INVX1_LOC_32/A 2.27fF
C41475 NOR2X1_LOC_168/B NOR2X1_LOC_500/B 0.04fF
C41476 INVX1_LOC_293/A INVX1_LOC_232/A 0.01fF
C41477 INVX1_LOC_58/A INVX1_LOC_6/A 1.37fF
C41478 INVX1_LOC_1/A NOR2X1_LOC_332/A 0.08fF
C41479 NOR2X1_LOC_89/A NOR2X1_LOC_378/Y 0.00fF
C41480 NOR2X1_LOC_607/a_36_216# INVX1_LOC_155/Y 0.00fF
C41481 VDD NOR2X1_LOC_623/B 0.08fF
C41482 INVX1_LOC_211/A INVX1_LOC_22/A 0.01fF
C41483 INVX1_LOC_54/Y INVX1_LOC_72/A 0.42fF
C41484 NAND2X1_LOC_579/A NOR2X1_LOC_71/Y 0.01fF
C41485 INVX1_LOC_146/Y NOR2X1_LOC_329/Y 0.11fF
C41486 INVX1_LOC_88/A NAND2X1_LOC_656/Y 0.17fF
C41487 INVX1_LOC_84/A NOR2X1_LOC_820/Y 0.05fF
C41488 NAND2X1_LOC_254/Y INVX1_LOC_280/A 0.02fF
C41489 NOR2X1_LOC_717/B NAND2X1_LOC_190/Y 0.00fF
C41490 NAND2X1_LOC_564/B NOR2X1_LOC_369/Y 0.01fF
C41491 VDD NOR2X1_LOC_329/Y 0.13fF
C41492 NAND2X1_LOC_785/Y INVX1_LOC_24/A 0.06fF
C41493 INVX1_LOC_91/A INVX1_LOC_270/Y 0.71fF
C41494 INVX1_LOC_36/A NAND2X1_LOC_181/Y 0.03fF
C41495 NOR2X1_LOC_92/Y INVX1_LOC_90/A 0.31fF
C41496 NOR2X1_LOC_246/A NOR2X1_LOC_361/B 0.08fF
C41497 INVX1_LOC_45/A NOR2X1_LOC_251/Y 0.23fF
C41498 NOR2X1_LOC_155/A INVX1_LOC_19/A 0.07fF
C41499 INVX1_LOC_24/Y INVX1_LOC_90/A 0.03fF
C41500 NAND2X1_LOC_454/Y INVX1_LOC_46/A 2.10fF
C41501 NOR2X1_LOC_68/A NOR2X1_LOC_547/B 0.01fF
C41502 INVX1_LOC_21/A NOR2X1_LOC_216/Y 0.01fF
C41503 NOR2X1_LOC_68/A NOR2X1_LOC_78/B 0.14fF
C41504 INVX1_LOC_5/A NOR2X1_LOC_188/A 0.07fF
C41505 NOR2X1_LOC_784/B NOR2X1_LOC_307/A 0.01fF
C41506 NAND2X1_LOC_468/B NAND2X1_LOC_424/a_36_24# 0.00fF
C41507 INVX1_LOC_215/A NOR2X1_LOC_441/Y 0.02fF
C41508 VDD NAND2X1_LOC_175/Y 2.32fF
C41509 INVX1_LOC_206/A INVX1_LOC_71/A 0.19fF
C41510 INVX1_LOC_41/A NOR2X1_LOC_147/B 0.03fF
C41511 NAND2X1_LOC_43/a_36_24# INVX1_LOC_83/A 0.01fF
C41512 NOR2X1_LOC_78/Y INVX1_LOC_284/A 0.08fF
C41513 NOR2X1_LOC_644/B INVX1_LOC_279/A 0.01fF
C41514 NOR2X1_LOC_48/B INVX1_LOC_54/A 0.04fF
C41515 INVX1_LOC_91/A NOR2X1_LOC_754/Y 0.02fF
C41516 NOR2X1_LOC_528/Y NAND2X1_LOC_793/B 0.10fF
C41517 NOR2X1_LOC_476/Y NOR2X1_LOC_375/Y 0.01fF
C41518 INVX1_LOC_214/A INVX1_LOC_24/A 1.09fF
C41519 INVX1_LOC_21/A NOR2X1_LOC_112/B 0.07fF
C41520 INVX1_LOC_34/A INVX1_LOC_8/A 0.11fF
C41521 INVX1_LOC_41/A NOR2X1_LOC_392/B 0.01fF
C41522 NOR2X1_LOC_667/A INVX1_LOC_24/A 0.07fF
C41523 INVX1_LOC_33/A INVX1_LOC_104/A 0.13fF
C41524 NAND2X1_LOC_733/Y INVX1_LOC_10/A 0.30fF
C41525 INVX1_LOC_136/A INVX1_LOC_22/A 1.47fF
C41526 INVX1_LOC_305/A NOR2X1_LOC_516/B 0.10fF
C41527 INVX1_LOC_248/A INVX1_LOC_24/A 0.07fF
C41528 NAND2X1_LOC_58/a_36_24# NAND2X1_LOC_348/A 0.01fF
C41529 NOR2X1_LOC_303/Y NOR2X1_LOC_537/Y 0.16fF
C41530 NOR2X1_LOC_172/Y NAND2X1_LOC_477/A 0.03fF
C41531 NOR2X1_LOC_743/a_36_216# INVX1_LOC_104/A 0.12fF
C41532 NOR2X1_LOC_590/A INVX1_LOC_150/A 0.16fF
C41533 NOR2X1_LOC_457/a_36_216# NOR2X1_LOC_151/Y 0.00fF
C41534 NOR2X1_LOC_617/Y NAND2X1_LOC_374/Y -0.04fF
C41535 NOR2X1_LOC_590/A NOR2X1_LOC_110/a_36_216# 0.00fF
C41536 NAND2X1_LOC_308/Y NAND2X1_LOC_811/Y 0.38fF
C41537 NOR2X1_LOC_500/A NAND2X1_LOC_323/B 0.01fF
C41538 NAND2X1_LOC_526/a_36_24# NOR2X1_LOC_713/B -0.02fF
C41539 NAND2X1_LOC_464/B INVX1_LOC_20/A 0.00fF
C41540 INVX1_LOC_45/A INVX1_LOC_234/A 0.00fF
C41541 INVX1_LOC_119/A NAND2X1_LOC_354/B 0.04fF
C41542 INVX1_LOC_274/A INVX1_LOC_15/A 1.61fF
C41543 NAND2X1_LOC_733/Y NOR2X1_LOC_504/a_36_216# 0.15fF
C41544 NOR2X1_LOC_590/A INVX1_LOC_89/A 8.03fF
C41545 VDD INVX1_LOC_262/A 0.12fF
C41546 D_INPUT_7 INPUT_5 0.30fF
C41547 NOR2X1_LOC_251/Y INVX1_LOC_71/A 0.03fF
C41548 NOR2X1_LOC_792/B NAND2X1_LOC_357/B 0.05fF
C41549 INVX1_LOC_60/A INVX1_LOC_60/Y 0.08fF
C41550 D_INPUT_2 INVX1_LOC_316/Y 0.46fF
C41551 NOR2X1_LOC_220/A NOR2X1_LOC_537/A 0.04fF
C41552 INVX1_LOC_22/Y INVX1_LOC_89/A 0.02fF
C41553 INVX1_LOC_157/A NOR2X1_LOC_52/Y 0.02fF
C41554 INVX1_LOC_217/A INVX1_LOC_10/A 0.07fF
C41555 INVX1_LOC_5/A NOR2X1_LOC_43/Y 0.08fF
C41556 NOR2X1_LOC_48/B NOR2X1_LOC_430/a_36_216# 0.00fF
C41557 VDD NOR2X1_LOC_622/A 0.12fF
C41558 INVX1_LOC_71/A INVX1_LOC_137/A 0.14fF
C41559 NOR2X1_LOC_590/A NAND2X1_LOC_508/A 0.06fF
C41560 NOR2X1_LOC_446/a_36_216# INVX1_LOC_182/A 0.00fF
C41561 NAND2X1_LOC_354/Y NOR2X1_LOC_130/A 0.02fF
C41562 INVX1_LOC_2/A INVX1_LOC_60/Y 0.10fF
C41563 NOR2X1_LOC_68/A INVX1_LOC_83/A 0.31fF
C41564 INVX1_LOC_290/A NOR2X1_LOC_152/Y 0.07fF
C41565 INVX1_LOC_49/A NOR2X1_LOC_835/A 0.10fF
C41566 NOR2X1_LOC_210/A INVX1_LOC_77/A 0.01fF
C41567 INVX1_LOC_263/A INVX1_LOC_33/A 0.73fF
C41568 INVX1_LOC_49/A NOR2X1_LOC_160/Y 0.02fF
C41569 NOR2X1_LOC_644/B INVX1_LOC_182/Y 0.00fF
C41570 INVX1_LOC_161/Y INVX1_LOC_144/A 0.07fF
C41571 INVX1_LOC_290/A INVX1_LOC_113/Y 0.03fF
C41572 INVX1_LOC_2/Y INVX1_LOC_138/A 0.02fF
C41573 NOR2X1_LOC_619/A NOR2X1_LOC_520/B 0.02fF
C41574 NOR2X1_LOC_717/B NOR2X1_LOC_596/A 0.06fF
C41575 INVX1_LOC_54/A NOR2X1_LOC_438/Y 0.06fF
C41576 INVX1_LOC_45/A NOR2X1_LOC_19/B 0.12fF
C41577 NAND2X1_LOC_53/Y NAND2X1_LOC_841/a_36_24# 0.00fF
C41578 INVX1_LOC_19/A NOR2X1_LOC_833/B 0.04fF
C41579 INVX1_LOC_54/Y NOR2X1_LOC_537/Y 0.00fF
C41580 INVX1_LOC_299/A INVX1_LOC_186/A 0.03fF
C41581 INPUT_3 NOR2X1_LOC_721/Y 0.01fF
C41582 INVX1_LOC_271/A NOR2X1_LOC_331/B 1.26fF
C41583 INVX1_LOC_209/Y INVX1_LOC_229/Y 0.03fF
C41584 INVX1_LOC_10/A NAND2X1_LOC_787/B 0.03fF
C41585 INVX1_LOC_40/Y INVX1_LOC_75/A 0.03fF
C41586 INVX1_LOC_76/A NOR2X1_LOC_460/Y 0.36fF
C41587 NOR2X1_LOC_355/A INVX1_LOC_49/A 0.01fF
C41588 NOR2X1_LOC_529/Y INVX1_LOC_316/Y 0.01fF
C41589 NOR2X1_LOC_531/a_36_216# NOR2X1_LOC_564/Y 0.00fF
C41590 NOR2X1_LOC_520/A INVX1_LOC_226/A 0.03fF
C41591 INVX1_LOC_17/A NOR2X1_LOC_78/A 0.13fF
C41592 INVX1_LOC_21/A NOR2X1_LOC_280/Y 0.03fF
C41593 INVX1_LOC_11/A NOR2X1_LOC_45/B 0.11fF
C41594 INVX1_LOC_303/A INVX1_LOC_132/Y 0.09fF
C41595 INVX1_LOC_313/Y NOR2X1_LOC_303/Y 0.10fF
C41596 NOR2X1_LOC_272/Y NOR2X1_LOC_266/B 0.01fF
C41597 INVX1_LOC_11/A NAND2X1_LOC_149/a_36_24# 0.01fF
C41598 VDD INVX1_LOC_171/Y 0.27fF
C41599 INVX1_LOC_269/A INVX1_LOC_95/Y 0.10fF
C41600 NOR2X1_LOC_383/Y NOR2X1_LOC_315/Y 0.43fF
C41601 INVX1_LOC_30/Y NOR2X1_LOC_316/Y 0.02fF
C41602 INVX1_LOC_299/A NAND2X1_LOC_447/Y 0.10fF
C41603 INVX1_LOC_2/A NOR2X1_LOC_222/a_36_216# 0.00fF
C41604 NOR2X1_LOC_250/Y NOR2X1_LOC_405/A 0.06fF
C41605 NOR2X1_LOC_92/Y NOR2X1_LOC_92/a_36_216# 0.02fF
C41606 NAND2X1_LOC_349/B NAND2X1_LOC_342/Y 0.00fF
C41607 INVX1_LOC_224/Y NOR2X1_LOC_216/B 1.72fF
C41608 NOR2X1_LOC_78/B NOR2X1_LOC_570/Y 0.05fF
C41609 NOR2X1_LOC_667/Y INVX1_LOC_91/A 0.02fF
C41610 INVX1_LOC_15/A NOR2X1_LOC_33/B 0.01fF
C41611 INVX1_LOC_41/A INVX1_LOC_90/A 0.13fF
C41612 INVX1_LOC_11/A INVX1_LOC_247/A 0.03fF
C41613 NOR2X1_LOC_151/Y NOR2X1_LOC_596/A 0.04fF
C41614 NOR2X1_LOC_468/Y NAND2X1_LOC_633/Y 0.02fF
C41615 NOR2X1_LOC_298/Y NOR2X1_LOC_504/Y 0.05fF
C41616 INVX1_LOC_227/A NOR2X1_LOC_493/B 0.02fF
C41617 NOR2X1_LOC_644/A NOR2X1_LOC_551/B 0.03fF
C41618 INVX1_LOC_201/Y INVX1_LOC_90/A 0.01fF
C41619 INVX1_LOC_313/Y NOR2X1_LOC_254/Y 0.01fF
C41620 INVX1_LOC_21/A NOR2X1_LOC_115/a_36_216# 0.02fF
C41621 INVX1_LOC_55/Y INVX1_LOC_153/Y 1.53fF
C41622 NOR2X1_LOC_445/Y NOR2X1_LOC_356/A 0.20fF
C41623 NAND2X1_LOC_391/Y NOR2X1_LOC_536/A 0.01fF
C41624 INVX1_LOC_228/A INPUT_0 0.01fF
C41625 NOR2X1_LOC_424/a_36_216# NOR2X1_LOC_222/Y 0.01fF
C41626 INVX1_LOC_214/A NAND2X1_LOC_783/A 0.10fF
C41627 NOR2X1_LOC_701/Y INVX1_LOC_22/A 0.30fF
C41628 INVX1_LOC_24/A INVX1_LOC_311/A 0.95fF
C41629 INVX1_LOC_27/A NOR2X1_LOC_331/B 0.07fF
C41630 INVX1_LOC_90/A NAND2X1_LOC_477/A 0.03fF
C41631 INVX1_LOC_182/A NOR2X1_LOC_570/B 0.07fF
C41632 NOR2X1_LOC_286/Y INVX1_LOC_37/A 0.03fF
C41633 INVX1_LOC_64/A NOR2X1_LOC_104/a_36_216# 0.03fF
C41634 INVX1_LOC_248/A NAND2X1_LOC_783/A 0.10fF
C41635 NOR2X1_LOC_632/Y INVX1_LOC_16/A 0.03fF
C41636 NOR2X1_LOC_97/A INVX1_LOC_77/A 0.01fF
C41637 NOR2X1_LOC_296/Y VDD 0.02fF
C41638 NOR2X1_LOC_778/B INVX1_LOC_135/A 0.02fF
C41639 NAND2X1_LOC_9/Y NOR2X1_LOC_49/a_36_216# 0.00fF
C41640 NOR2X1_LOC_717/B NOR2X1_LOC_220/A 0.03fF
C41641 INVX1_LOC_78/A INVX1_LOC_114/Y 0.01fF
C41642 NOR2X1_LOC_92/Y INVX1_LOC_38/A 0.18fF
C41643 INVX1_LOC_23/A NAND2X1_LOC_475/Y 0.10fF
C41644 INVX1_LOC_55/Y INVX1_LOC_177/A 0.03fF
C41645 NOR2X1_LOC_419/Y INVX1_LOC_51/Y 0.02fF
C41646 INVX1_LOC_93/A NAND2X1_LOC_444/a_36_24# 0.01fF
C41647 INVX1_LOC_183/A INVX1_LOC_29/A 0.01fF
C41648 NOR2X1_LOC_445/Y NOR2X1_LOC_74/A 0.17fF
C41649 INVX1_LOC_49/A NOR2X1_LOC_552/Y 0.00fF
C41650 INPUT_3 VDD 2.08fF
C41651 NOR2X1_LOC_92/Y NOR2X1_LOC_96/Y 0.03fF
C41652 INVX1_LOC_2/A NOR2X1_LOC_736/Y 0.13fF
C41653 NOR2X1_LOC_214/B NAND2X1_LOC_841/A 0.04fF
C41654 INPUT_0 INVX1_LOC_8/A 0.17fF
C41655 INVX1_LOC_259/Y INVX1_LOC_186/Y 0.00fF
C41656 NOR2X1_LOC_13/Y NAND2X1_LOC_655/A 0.01fF
C41657 INVX1_LOC_221/Y NOR2X1_LOC_536/A 0.01fF
C41658 INVX1_LOC_33/A INVX1_LOC_206/Y 0.03fF
C41659 D_INPUT_0 NOR2X1_LOC_86/A 1.45fF
C41660 INVX1_LOC_268/A NOR2X1_LOC_214/B 0.27fF
C41661 NOR2X1_LOC_334/Y INVX1_LOC_4/A 0.07fF
C41662 INVX1_LOC_78/A NOR2X1_LOC_467/A 0.12fF
C41663 INVX1_LOC_21/A NOR2X1_LOC_197/B 3.71fF
C41664 NAND2X1_LOC_63/Y INVX1_LOC_29/Y 0.00fF
C41665 NAND2X1_LOC_323/B NOR2X1_LOC_112/Y 0.04fF
C41666 INVX1_LOC_90/A NOR2X1_LOC_211/A 0.23fF
C41667 NOR2X1_LOC_598/B INVX1_LOC_19/A 0.53fF
C41668 NOR2X1_LOC_433/A NOR2X1_LOC_45/B 4.13fF
C41669 INVX1_LOC_83/A NOR2X1_LOC_545/a_36_216# 0.02fF
C41670 NAND2X1_LOC_348/A INVX1_LOC_64/Y 0.05fF
C41671 NOR2X1_LOC_389/B NOR2X1_LOC_211/A 0.01fF
C41672 NOR2X1_LOC_92/Y NAND2X1_LOC_848/Y 0.02fF
C41673 NOR2X1_LOC_246/A NAND2X1_LOC_573/A 0.10fF
C41674 NOR2X1_LOC_13/Y NAND2X1_LOC_468/B 0.05fF
C41675 INVX1_LOC_84/A INVX1_LOC_306/Y 1.72fF
C41676 INVX1_LOC_25/A NOR2X1_LOC_847/A 0.07fF
C41677 INVX1_LOC_234/Y INVX1_LOC_260/Y 0.15fF
C41678 NOR2X1_LOC_220/A NOR2X1_LOC_151/Y 0.03fF
C41679 NOR2X1_LOC_122/A NOR2X1_LOC_155/A 0.01fF
C41680 INVX1_LOC_36/A INVX1_LOC_117/A 0.14fF
C41681 INVX1_LOC_25/A INVX1_LOC_42/A 0.14fF
C41682 INVX1_LOC_272/Y INVX1_LOC_92/A 0.07fF
C41683 NOR2X1_LOC_763/Y INVX1_LOC_89/A 0.06fF
C41684 INVX1_LOC_90/A INVX1_LOC_121/A 0.23fF
C41685 NAND2X1_LOC_350/A INVX1_LOC_54/A 0.15fF
C41686 INVX1_LOC_151/A NOR2X1_LOC_45/B 0.01fF
C41687 NAND2X1_LOC_731/a_36_24# INVX1_LOC_28/A 0.00fF
C41688 NAND2X1_LOC_53/Y INVX1_LOC_92/A 0.19fF
C41689 INVX1_LOC_73/A INVX1_LOC_1/Y 0.07fF
C41690 INVX1_LOC_11/A NOR2X1_LOC_862/B 0.03fF
C41691 NOR2X1_LOC_310/Y INVX1_LOC_91/A 0.05fF
C41692 NOR2X1_LOC_52/B NOR2X1_LOC_45/B 0.24fF
C41693 INVX1_LOC_83/A NOR2X1_LOC_163/A 0.01fF
C41694 NOR2X1_LOC_655/B INVX1_LOC_286/A 0.10fF
C41695 NOR2X1_LOC_103/Y NOR2X1_LOC_216/B 0.10fF
C41696 INVX1_LOC_209/Y INVX1_LOC_20/A 0.06fF
C41697 NOR2X1_LOC_441/Y INVX1_LOC_54/A 4.34fF
C41698 INVX1_LOC_161/Y NOR2X1_LOC_155/A 0.07fF
C41699 NOR2X1_LOC_368/A INVX1_LOC_56/Y 0.08fF
C41700 NAND2X1_LOC_537/Y INVX1_LOC_119/Y 0.00fF
C41701 INVX1_LOC_122/Y INVX1_LOC_9/A 0.03fF
C41702 NAND2X1_LOC_357/A INVX1_LOC_285/A 0.11fF
C41703 NOR2X1_LOC_542/Y NOR2X1_LOC_356/A -0.03fF
C41704 INVX1_LOC_153/Y NOR2X1_LOC_357/Y 0.10fF
C41705 INVX1_LOC_49/A NOR2X1_LOC_111/A 0.03fF
C41706 NOR2X1_LOC_91/A NOR2X1_LOC_167/a_36_216# 0.00fF
C41707 INVX1_LOC_23/Y NAND2X1_LOC_99/A 0.02fF
C41708 NAND2X1_LOC_849/B NAND2X1_LOC_837/Y 0.38fF
C41709 INVX1_LOC_147/A INVX1_LOC_83/A 0.39fF
C41710 NAND2X1_LOC_778/Y INVX1_LOC_102/A 0.10fF
C41711 NOR2X1_LOC_778/B NOR2X1_LOC_552/A 0.08fF
C41712 NAND2X1_LOC_833/Y NAND2X1_LOC_721/A 0.13fF
C41713 NOR2X1_LOC_103/Y NAND2X1_LOC_477/Y 0.01fF
C41714 NAND2X1_LOC_837/Y INVX1_LOC_38/A 0.07fF
C41715 INVX1_LOC_25/A INVX1_LOC_78/A 0.07fF
C41716 NOR2X1_LOC_613/Y NOR2X1_LOC_89/A 0.01fF
C41717 NOR2X1_LOC_433/A INVX1_LOC_281/A 0.07fF
C41718 NOR2X1_LOC_804/B INVX1_LOC_117/A 0.41fF
C41719 INVX1_LOC_45/A NOR2X1_LOC_216/B 0.27fF
C41720 INVX1_LOC_136/A NOR2X1_LOC_88/A 0.04fF
C41721 NOR2X1_LOC_332/A NOR2X1_LOC_188/A 0.14fF
C41722 INVX1_LOC_158/A VDD 0.25fF
C41723 INVX1_LOC_64/A NOR2X1_LOC_334/Y 0.57fF
C41724 INVX1_LOC_41/A NOR2X1_LOC_561/A 0.05fF
C41725 NAND2X1_LOC_7/Y INVX1_LOC_9/A 0.41fF
C41726 NOR2X1_LOC_510/Y INVX1_LOC_32/A 0.00fF
C41727 INVX1_LOC_1/A NOR2X1_LOC_847/A 0.07fF
C41728 NAND2X1_LOC_134/a_36_24# INVX1_LOC_46/A 0.01fF
C41729 INVX1_LOC_294/Y NOR2X1_LOC_440/a_36_216# 0.01fF
C41730 NOR2X1_LOC_328/Y INPUT_4 0.01fF
C41731 NOR2X1_LOC_15/Y INVX1_LOC_102/A 0.16fF
C41732 INVX1_LOC_41/A INVX1_LOC_38/A 0.03fF
C41733 NOR2X1_LOC_712/Y NOR2X1_LOC_707/A 0.01fF
C41734 INVX1_LOC_1/A INVX1_LOC_42/A 0.13fF
C41735 NAND2X1_LOC_116/A NAND2X1_LOC_96/A 0.07fF
C41736 INVX1_LOC_33/A NOR2X1_LOC_119/a_36_216# 0.00fF
C41737 NOR2X1_LOC_598/B INVX1_LOC_26/Y 0.03fF
C41738 NOR2X1_LOC_276/a_36_216# NOR2X1_LOC_155/A 0.00fF
C41739 NOR2X1_LOC_667/A NOR2X1_LOC_280/Y 0.08fF
C41740 NOR2X1_LOC_498/Y INVX1_LOC_38/A 0.07fF
C41741 NOR2X1_LOC_307/A NOR2X1_LOC_777/B 0.00fF
C41742 INVX1_LOC_173/A NAND2X1_LOC_408/a_36_24# 0.02fF
C41743 NOR2X1_LOC_335/B NOR2X1_LOC_356/A 0.01fF
C41744 NOR2X1_LOC_91/A NAND2X1_LOC_787/A 0.03fF
C41745 NOR2X1_LOC_52/B INVX1_LOC_281/A 0.06fF
C41746 INVX1_LOC_2/A NOR2X1_LOC_111/A 2.41fF
C41747 INVX1_LOC_311/Y NOR2X1_LOC_74/A 0.03fF
C41748 NOR2X1_LOC_318/B NOR2X1_LOC_335/a_36_216# 0.00fF
C41749 INVX1_LOC_13/A INVX1_LOC_316/A 0.04fF
C41750 NOR2X1_LOC_666/A NOR2X1_LOC_270/a_36_216# 0.00fF
C41751 D_INPUT_1 INVX1_LOC_57/A 7.50fF
C41752 NAND2X1_LOC_776/a_36_24# INVX1_LOC_84/A 0.00fF
C41753 NOR2X1_LOC_488/Y NAND2X1_LOC_244/A 0.00fF
C41754 NAND2X1_LOC_363/B NOR2X1_LOC_668/Y 0.01fF
C41755 INVX1_LOC_62/A NOR2X1_LOC_845/A 0.19fF
C41756 NAND2X1_LOC_525/a_36_24# INVX1_LOC_75/A 0.00fF
C41757 INVX1_LOC_9/Y NOR2X1_LOC_136/a_36_216# 0.00fF
C41758 NAND2X1_LOC_672/B D_INPUT_3 0.01fF
C41759 INVX1_LOC_71/A NOR2X1_LOC_216/B 1.51fF
C41760 NOR2X1_LOC_530/a_36_216# INVX1_LOC_284/A 0.00fF
C41761 NAND2X1_LOC_477/A INVX1_LOC_38/A 0.03fF
C41762 NOR2X1_LOC_142/Y INVX1_LOC_54/A 1.51fF
C41763 D_INPUT_0 NOR2X1_LOC_405/A 0.07fF
C41764 NOR2X1_LOC_510/Y NAND2X1_LOC_175/Y 0.64fF
C41765 INVX1_LOC_9/Y VDD 0.24fF
C41766 NOR2X1_LOC_383/B INVX1_LOC_292/Y 0.10fF
C41767 NOR2X1_LOC_361/B INVX1_LOC_32/A 1.69fF
C41768 NOR2X1_LOC_667/A NAND2X1_LOC_811/B 0.03fF
C41769 NOR2X1_LOC_186/Y NOR2X1_LOC_301/A 0.09fF
C41770 NAND2X1_LOC_733/Y INVX1_LOC_12/A 0.03fF
C41771 NAND2X1_LOC_564/B VDD 0.19fF
C41772 NAND2X1_LOC_350/A NOR2X1_LOC_48/B 0.10fF
C41773 INVX1_LOC_304/A NOR2X1_LOC_130/A 0.07fF
C41774 NAND2X1_LOC_363/B INVX1_LOC_23/A 0.07fF
C41775 INVX1_LOC_280/Y NOR2X1_LOC_692/Y 0.08fF
C41776 NOR2X1_LOC_174/B INVX1_LOC_65/A 0.12fF
C41777 GATE_662 VDD 0.07fF
C41778 NAND2X1_LOC_451/a_36_24# NAND2X1_LOC_639/A 0.01fF
C41779 INVX1_LOC_58/A NOR2X1_LOC_109/Y 2.02fF
C41780 INVX1_LOC_1/A INVX1_LOC_78/A 0.21fF
C41781 INVX1_LOC_88/A INVX1_LOC_128/Y 0.13fF
C41782 NAND2X1_LOC_573/Y NOR2X1_LOC_301/A 0.20fF
C41783 NOR2X1_LOC_60/a_36_216# INVX1_LOC_76/A 0.01fF
C41784 INVX1_LOC_18/A NAND2X1_LOC_74/B 0.10fF
C41785 INVX1_LOC_24/Y INVX1_LOC_18/Y 0.09fF
C41786 INVX1_LOC_57/A NOR2X1_LOC_652/Y 0.71fF
C41787 INVX1_LOC_217/A INVX1_LOC_12/A 0.07fF
C41788 D_INPUT_0 NOR2X1_LOC_857/A 0.16fF
C41789 NOR2X1_LOC_211/A INVX1_LOC_38/A 0.01fF
C41790 INVX1_LOC_73/A NOR2X1_LOC_318/B 0.07fF
C41791 NOR2X1_LOC_772/B NOR2X1_LOC_717/A 0.10fF
C41792 INVX1_LOC_217/A NOR2X1_LOC_519/Y 0.11fF
C41793 INVX1_LOC_69/Y NOR2X1_LOC_500/a_36_216# 0.14fF
C41794 NOR2X1_LOC_791/Y INVX1_LOC_23/A 0.05fF
C41795 NOR2X1_LOC_384/Y INVX1_LOC_42/A 0.09fF
C41796 NAND2X1_LOC_848/A NOR2X1_LOC_86/A 0.07fF
C41797 INVX1_LOC_16/A NOR2X1_LOC_186/a_36_216# 0.00fF
C41798 INVX1_LOC_73/A INVX1_LOC_93/Y 0.07fF
C41799 INVX1_LOC_13/Y NOR2X1_LOC_717/A 0.67fF
C41800 NOR2X1_LOC_65/B INVX1_LOC_1/A 0.03fF
C41801 INVX1_LOC_278/A INVX1_LOC_306/Y 0.10fF
C41802 D_INPUT_1 INVX1_LOC_252/A 0.01fF
C41803 NAND2X1_LOC_734/B INVX1_LOC_285/A 0.14fF
C41804 INVX1_LOC_280/Y INVX1_LOC_260/A 0.00fF
C41805 NOR2X1_LOC_657/Y INVX1_LOC_15/A 0.02fF
C41806 NAND2X1_LOC_338/B INVX1_LOC_35/Y 0.04fF
C41807 INVX1_LOC_121/A INVX1_LOC_38/A 0.07fF
C41808 NOR2X1_LOC_589/A NAND2X1_LOC_637/Y 0.60fF
C41809 NOR2X1_LOC_769/A NOR2X1_LOC_467/A 0.33fF
C41810 NOR2X1_LOC_500/Y INVX1_LOC_92/A 0.16fF
C41811 NAND2X1_LOC_156/B NOR2X1_LOC_331/B 0.15fF
C41812 INVX1_LOC_174/A NAND2X1_LOC_70/a_36_24# 0.01fF
C41813 NAND2X1_LOC_787/B INVX1_LOC_12/A 0.09fF
C41814 INVX1_LOC_113/Y INVX1_LOC_114/Y 0.01fF
C41815 INVX1_LOC_82/Y D_INPUT_3 0.01fF
C41816 NAND2X1_LOC_578/B NOR2X1_LOC_649/B 0.03fF
C41817 INVX1_LOC_137/Y NAND2X1_LOC_93/B 0.01fF
C41818 INVX1_LOC_137/A NAND2X1_LOC_92/a_36_24# 0.01fF
C41819 NOR2X1_LOC_781/A INVX1_LOC_117/Y 0.29fF
C41820 INVX1_LOC_147/A INVX1_LOC_46/A 0.29fF
C41821 NOR2X1_LOC_329/B INVX1_LOC_33/Y 0.00fF
C41822 NOR2X1_LOC_775/Y NAND2X1_LOC_96/A 0.03fF
C41823 NOR2X1_LOC_561/Y INVX1_LOC_180/Y 0.04fF
C41824 NOR2X1_LOC_457/A INVX1_LOC_23/A 0.16fF
C41825 NOR2X1_LOC_537/Y NOR2X1_LOC_721/B 0.03fF
C41826 INVX1_LOC_272/Y INVX1_LOC_53/A 0.07fF
C41827 NAND2X1_LOC_338/B NOR2X1_LOC_721/B 0.01fF
C41828 INVX1_LOC_10/A INVX1_LOC_92/A 0.10fF
C41829 NAND2X1_LOC_660/A INVX1_LOC_19/A 0.13fF
C41830 INVX1_LOC_25/Y INVX1_LOC_285/A 0.08fF
C41831 INVX1_LOC_50/A NOR2X1_LOC_595/a_36_216# 0.00fF
C41832 NAND2X1_LOC_181/Y INVX1_LOC_63/A 0.72fF
C41833 NOR2X1_LOC_152/Y NOR2X1_LOC_467/A 0.01fF
C41834 INVX1_LOC_285/Y NOR2X1_LOC_357/Y 0.03fF
C41835 INVX1_LOC_304/Y INVX1_LOC_12/A 0.07fF
C41836 INVX1_LOC_266/Y INVX1_LOC_29/A 0.05fF
C41837 NOR2X1_LOC_217/a_36_216# NOR2X1_LOC_678/A 0.00fF
C41838 NOR2X1_LOC_91/A INVX1_LOC_30/A 0.26fF
C41839 INVX1_LOC_113/Y NOR2X1_LOC_467/A 0.00fF
C41840 INVX1_LOC_221/A INVX1_LOC_42/A 0.04fF
C41841 NOR2X1_LOC_93/Y INVX1_LOC_59/A 0.07fF
C41842 INVX1_LOC_50/A NOR2X1_LOC_717/Y 0.03fF
C41843 NOR2X1_LOC_486/Y NOR2X1_LOC_600/Y 0.12fF
C41844 NOR2X1_LOC_577/Y NAND2X1_LOC_647/B 0.00fF
C41845 INVX1_LOC_220/Y INVX1_LOC_220/A 0.19fF
C41846 NOR2X1_LOC_123/B NOR2X1_LOC_216/B 0.10fF
C41847 NAND2X1_LOC_787/A INVX1_LOC_31/A 0.03fF
C41848 NAND2X1_LOC_390/A INVX1_LOC_63/A 0.31fF
C41849 NOR2X1_LOC_601/Y INVX1_LOC_247/A 0.06fF
C41850 INVX1_LOC_200/Y INVX1_LOC_57/Y 0.03fF
C41851 INVX1_LOC_30/A INVX1_LOC_23/A 2.79fF
C41852 NAND2X1_LOC_656/A INVX1_LOC_23/Y 0.04fF
C41853 INVX1_LOC_62/Y NOR2X1_LOC_39/a_36_216# 0.01fF
C41854 INVX1_LOC_286/A NOR2X1_LOC_176/Y 0.03fF
C41855 INVX1_LOC_199/A INVX1_LOC_199/Y 0.04fF
C41856 INVX1_LOC_58/A INVX1_LOC_36/A 1.06fF
C41857 INVX1_LOC_17/A NOR2X1_LOC_186/Y 0.22fF
C41858 NAND2X1_LOC_363/B INVX1_LOC_31/A 0.07fF
C41859 INVX1_LOC_89/A NOR2X1_LOC_688/a_36_216# 0.00fF
C41860 NOR2X1_LOC_848/Y INVX1_LOC_27/A 0.03fF
C41861 INVX1_LOC_135/A NAND2X1_LOC_657/a_36_24# 0.00fF
C41862 INVX1_LOC_309/A NOR2X1_LOC_536/A 1.88fF
C41863 INVX1_LOC_25/A NOR2X1_LOC_554/B 0.21fF
C41864 NOR2X1_LOC_453/Y NOR2X1_LOC_470/B 0.01fF
C41865 INVX1_LOC_41/A NAND2X1_LOC_223/A 0.03fF
C41866 INVX1_LOC_177/A INVX1_LOC_32/A 0.03fF
C41867 NAND2X1_LOC_860/A INVX1_LOC_72/A 0.09fF
C41868 NAND2X1_LOC_724/Y INVX1_LOC_300/Y 0.13fF
C41869 INVX1_LOC_172/Y INVX1_LOC_284/A 0.02fF
C41870 NAND2X1_LOC_565/a_36_24# INVX1_LOC_31/A 0.00fF
C41871 NAND2X1_LOC_739/B INVX1_LOC_50/A 0.03fF
C41872 NOR2X1_LOC_114/A NOR2X1_LOC_536/A 0.03fF
C41873 INVX1_LOC_17/A NAND2X1_LOC_573/Y 0.98fF
C41874 NAND2X1_LOC_639/A INVX1_LOC_91/A 0.02fF
C41875 INVX1_LOC_259/Y INVX1_LOC_18/A 0.02fF
C41876 NAND2X1_LOC_725/A NOR2X1_LOC_599/A 0.03fF
C41877 NAND2X1_LOC_9/Y NOR2X1_LOC_68/A 0.10fF
C41878 NOR2X1_LOC_647/Y NOR2X1_LOC_660/Y 0.19fF
C41879 INVX1_LOC_277/A INVX1_LOC_5/A 0.02fF
C41880 INVX1_LOC_223/Y NOR2X1_LOC_590/A 0.05fF
C41881 NOR2X1_LOC_536/A INVX1_LOC_91/A 0.42fF
C41882 NOR2X1_LOC_383/a_36_216# NAND2X1_LOC_74/B 0.00fF
C41883 INVX1_LOC_58/A NOR2X1_LOC_208/Y 0.10fF
C41884 INVX1_LOC_95/Y INVX1_LOC_12/Y 0.10fF
C41885 NAND2X1_LOC_656/Y INVX1_LOC_272/A 0.53fF
C41886 NOR2X1_LOC_714/a_36_216# NOR2X1_LOC_729/A 0.02fF
C41887 NOR2X1_LOC_356/A INVX1_LOC_84/A 0.04fF
C41888 VDD NOR2X1_LOC_279/Y 0.00fF
C41889 INVX1_LOC_225/A NOR2X1_LOC_301/A 1.61fF
C41890 NOR2X1_LOC_731/A NOR2X1_LOC_307/Y 0.07fF
C41891 NAND2X1_LOC_361/Y NOR2X1_LOC_383/B 0.07fF
C41892 NAND2X1_LOC_555/Y NAND2X1_LOC_574/a_36_24# 0.01fF
C41893 NAND2X1_LOC_326/A NOR2X1_LOC_816/A 0.07fF
C41894 INVX1_LOC_37/A INVX1_LOC_115/A 0.04fF
C41895 INVX1_LOC_21/A INVX1_LOC_286/Y 0.08fF
C41896 INVX1_LOC_64/A NOR2X1_LOC_523/B 0.01fF
C41897 NOR2X1_LOC_74/A NOR2X1_LOC_88/Y 0.07fF
C41898 INVX1_LOC_195/Y INVX1_LOC_253/Y 0.01fF
C41899 INVX1_LOC_199/A INVX1_LOC_281/A 0.01fF
C41900 NOR2X1_LOC_682/Y NOR2X1_LOC_682/a_36_216# 0.01fF
C41901 INVX1_LOC_2/Y D_INPUT_3 0.00fF
C41902 INVX1_LOC_57/Y NOR2X1_LOC_406/A 0.00fF
C41903 NOR2X1_LOC_246/A NAND2X1_LOC_81/B 0.00fF
C41904 INVX1_LOC_11/Y NOR2X1_LOC_536/A 0.06fF
C41905 NOR2X1_LOC_585/Y NAND2X1_LOC_637/a_36_24# 0.00fF
C41906 NAND2X1_LOC_850/Y NAND2X1_LOC_444/B 0.03fF
C41907 INVX1_LOC_298/Y INVX1_LOC_266/Y 0.07fF
C41908 INVX1_LOC_144/A NOR2X1_LOC_841/A 0.02fF
C41909 NOR2X1_LOC_829/Y NAND2X1_LOC_811/Y 0.02fF
C41910 INVX1_LOC_75/A INVX1_LOC_285/A 0.08fF
C41911 INVX1_LOC_75/A NOR2X1_LOC_814/A 2.05fF
C41912 VDD NAND2X1_LOC_804/Y 0.26fF
C41913 NOR2X1_LOC_798/A NOR2X1_LOC_68/A 0.05fF
C41914 NOR2X1_LOC_644/B NAND2X1_LOC_190/Y 0.00fF
C41915 INVX1_LOC_72/A INVX1_LOC_242/A 0.02fF
C41916 NOR2X1_LOC_91/A NAND2X1_LOC_722/A 0.09fF
C41917 INVX1_LOC_91/A NAND2X1_LOC_93/B 0.39fF
C41918 INVX1_LOC_104/A NOR2X1_LOC_748/A 0.10fF
C41919 NOR2X1_LOC_74/A INVX1_LOC_84/A 0.13fF
C41920 NOR2X1_LOC_569/Y INVX1_LOC_4/A 0.02fF
C41921 NOR2X1_LOC_209/Y NOR2X1_LOC_302/A 0.01fF
C41922 NAND2X1_LOC_573/A INVX1_LOC_32/A 0.34fF
C41923 INVX1_LOC_21/A INVX1_LOC_159/A 0.03fF
C41924 INVX1_LOC_58/A NOR2X1_LOC_309/Y 0.04fF
C41925 NOR2X1_LOC_15/Y INVX1_LOC_223/A 0.07fF
C41926 INVX1_LOC_13/A INVX1_LOC_4/Y 0.03fF
C41927 NOR2X1_LOC_476/Y INVX1_LOC_163/A 0.07fF
C41928 NOR2X1_LOC_391/A NOR2X1_LOC_38/B 0.00fF
C41929 NOR2X1_LOC_626/Y INVX1_LOC_24/A 0.02fF
C41930 NOR2X1_LOC_68/A NAND2X1_LOC_703/Y 0.02fF
C41931 NAND2X1_LOC_721/A NAND2X1_LOC_837/a_36_24# 0.01fF
C41932 INVX1_LOC_91/A NAND2X1_LOC_425/Y 0.64fF
C41933 NOR2X1_LOC_9/Y INVX1_LOC_84/A 0.07fF
C41934 INVX1_LOC_2/Y INVX1_LOC_230/A 0.21fF
C41935 NOR2X1_LOC_135/Y INVX1_LOC_109/A 0.01fF
C41936 INVX1_LOC_77/A INVX1_LOC_50/Y 0.03fF
C41937 NAND2X1_LOC_537/Y INVX1_LOC_72/A 0.10fF
C41938 INVX1_LOC_1/A NOR2X1_LOC_554/B 0.29fF
C41939 INVX1_LOC_22/A NOR2X1_LOC_395/Y 0.05fF
C41940 NOR2X1_LOC_655/B NAND2X1_LOC_215/A 0.10fF
C41941 NOR2X1_LOC_620/B INVX1_LOC_57/A 0.00fF
C41942 INVX1_LOC_10/A NAND2X1_LOC_247/a_36_24# 0.00fF
C41943 NOR2X1_LOC_272/Y INVX1_LOC_49/A 0.01fF
C41944 NAND2X1_LOC_655/A NOR2X1_LOC_697/Y 0.01fF
C41945 NOR2X1_LOC_185/a_36_216# NAND2X1_LOC_74/B 0.01fF
C41946 NOR2X1_LOC_366/B INVX1_LOC_271/A 0.01fF
C41947 INVX1_LOC_91/A INVX1_LOC_3/A 0.77fF
C41948 NOR2X1_LOC_111/A INVX1_LOC_118/A 0.10fF
C41949 NAND2X1_LOC_860/A NAND2X1_LOC_338/B 1.20fF
C41950 NOR2X1_LOC_356/A INVX1_LOC_15/A 0.07fF
C41951 NAND2X1_LOC_784/A NOR2X1_LOC_773/Y 0.01fF
C41952 NAND2X1_LOC_757/a_36_24# INVX1_LOC_14/A -0.02fF
C41953 NOR2X1_LOC_176/Y INVX1_LOC_54/A 0.03fF
C41954 NOR2X1_LOC_13/Y INVX1_LOC_88/A 0.01fF
C41955 INVX1_LOC_266/A INVX1_LOC_77/A 0.01fF
C41956 NAND2X1_LOC_9/Y NOR2X1_LOC_520/a_36_216# 0.01fF
C41957 INVX1_LOC_5/A NOR2X1_LOC_87/B 0.07fF
C41958 INVX1_LOC_31/A INVX1_LOC_30/A 0.39fF
C41959 NOR2X1_LOC_188/A INVX1_LOC_42/A 0.07fF
C41960 INVX1_LOC_1/A INVX1_LOC_113/Y 0.05fF
C41961 NOR2X1_LOC_86/a_36_216# INVX1_LOC_284/A 0.00fF
C41962 NOR2X1_LOC_500/Y INVX1_LOC_53/A 1.38fF
C41963 INVX1_LOC_89/A NOR2X1_LOC_415/Y 0.01fF
C41964 NOR2X1_LOC_773/Y NOR2X1_LOC_129/a_36_216# 0.01fF
C41965 NOR2X1_LOC_19/Y INVX1_LOC_3/Y 0.18fF
C41966 NAND2X1_LOC_733/Y INVX1_LOC_217/A 0.10fF
C41967 INVX1_LOC_24/Y INVX1_LOC_33/A 0.03fF
C41968 NAND2X1_LOC_550/A NOR2X1_LOC_238/Y -0.03fF
C41969 INVX1_LOC_174/A INVX1_LOC_24/A 0.08fF
C41970 INVX1_LOC_17/A INVX1_LOC_132/A 0.07fF
C41971 INVX1_LOC_161/Y NOR2X1_LOC_513/a_36_216# 0.01fF
C41972 NOR2X1_LOC_590/A NOR2X1_LOC_744/a_36_216# 0.00fF
C41973 NOR2X1_LOC_74/A INVX1_LOC_15/A 0.20fF
C41974 INVX1_LOC_88/A NAND2X1_LOC_175/B 0.05fF
C41975 NAND2X1_LOC_656/Y NOR2X1_LOC_125/a_36_216# 0.00fF
C41976 INVX1_LOC_17/A NOR2X1_LOC_481/A 0.10fF
C41977 INVX1_LOC_17/A NAND2X1_LOC_640/Y 0.01fF
C41978 NOR2X1_LOC_644/B NOR2X1_LOC_596/A 0.07fF
C41979 NOR2X1_LOC_15/Y INVX1_LOC_162/Y 0.03fF
C41980 NAND2X1_LOC_787/A NAND2X1_LOC_859/Y 0.02fF
C41981 INVX1_LOC_114/A INVX1_LOC_92/A 0.04fF
C41982 NOR2X1_LOC_709/A NOR2X1_LOC_440/B 0.00fF
C41983 NOR2X1_LOC_286/Y INVX1_LOC_310/Y 0.11fF
C41984 NOR2X1_LOC_360/A NAND2X1_LOC_206/Y 0.06fF
C41985 INVX1_LOC_135/A INVX1_LOC_271/A 0.01fF
C41986 NOR2X1_LOC_15/Y INVX1_LOC_85/A 0.03fF
C41987 NOR2X1_LOC_272/Y NOR2X1_LOC_226/A 0.10fF
C41988 INVX1_LOC_136/A INVX1_LOC_18/A 0.54fF
C41989 INVX1_LOC_10/A INVX1_LOC_53/A 0.35fF
C41990 NOR2X1_LOC_45/B NAND2X1_LOC_254/Y 1.83fF
C41991 NOR2X1_LOC_78/B NAND2X1_LOC_474/Y 0.07fF
C41992 INVX1_LOC_20/A NAND2X1_LOC_773/B 0.47fF
C41993 NAND2X1_LOC_728/Y INVX1_LOC_136/A 0.07fF
C41994 INVX1_LOC_17/A INVX1_LOC_225/A 0.10fF
C41995 NOR2X1_LOC_537/Y NAND2X1_LOC_473/A 0.14fF
C41996 INVX1_LOC_12/A NOR2X1_LOC_56/a_36_216# 0.00fF
C41997 INVX1_LOC_30/A INVX1_LOC_111/A 0.01fF
C41998 INVX1_LOC_27/A NOR2X1_LOC_366/B 0.01fF
C41999 NAND2X1_LOC_218/B INVX1_LOC_40/Y 0.03fF
C42000 NAND2X1_LOC_273/a_36_24# NOR2X1_LOC_536/A 0.00fF
C42001 INVX1_LOC_25/A NOR2X1_LOC_150/a_36_216# 0.00fF
C42002 INVX1_LOC_45/A NOR2X1_LOC_303/Y 0.03fF
C42003 NAND2X1_LOC_733/Y NAND2X1_LOC_787/B 0.03fF
C42004 INVX1_LOC_41/A NOR2X1_LOC_483/B 0.06fF
C42005 NOR2X1_LOC_188/A INVX1_LOC_78/A 0.10fF
C42006 NOR2X1_LOC_568/A NOR2X1_LOC_303/Y 0.10fF
C42007 NOR2X1_LOC_272/Y NOR2X1_LOC_218/Y 0.06fF
C42008 INVX1_LOC_304/Y INVX1_LOC_200/A 0.22fF
C42009 INVX1_LOC_117/A INVX1_LOC_63/A 0.07fF
C42010 NOR2X1_LOC_92/Y NAND2X1_LOC_798/A 0.03fF
C42011 NAND2X1_LOC_854/B NOR2X1_LOC_304/Y 0.04fF
C42012 INVX1_LOC_188/Y INVX1_LOC_290/Y 0.01fF
C42013 NAND2X1_LOC_198/B INVX1_LOC_181/Y 0.10fF
C42014 INVX1_LOC_27/A NAND2X1_LOC_479/Y 0.07fF
C42015 INVX1_LOC_1/A NOR2X1_LOC_307/B 0.05fF
C42016 NAND2X1_LOC_787/A NAND2X1_LOC_866/B 0.01fF
C42017 NOR2X1_LOC_631/A INVX1_LOC_44/A 0.40fF
C42018 NAND2X1_LOC_560/a_36_24# NAND2X1_LOC_733/B 0.01fF
C42019 INVX1_LOC_136/A INVX1_LOC_172/A 0.07fF
C42020 INVX1_LOC_307/A INVX1_LOC_92/A 0.01fF
C42021 NOR2X1_LOC_536/A INVX1_LOC_203/A 0.03fF
C42022 INVX1_LOC_103/A INVX1_LOC_144/Y -0.02fF
C42023 NOR2X1_LOC_858/a_36_216# NOR2X1_LOC_862/B 0.02fF
C42024 NAND2X1_LOC_214/B INVX1_LOC_135/A 0.06fF
C42025 NAND2X1_LOC_364/A INVX1_LOC_49/A 0.09fF
C42026 NAND2X1_LOC_392/Y NAND2X1_LOC_474/Y 0.14fF
C42027 NAND2X1_LOC_53/Y NOR2X1_LOC_78/B 0.12fF
C42028 NAND2X1_LOC_30/Y NAND2X1_LOC_11/Y 0.13fF
C42029 INVX1_LOC_217/A NAND2X1_LOC_787/B 0.23fF
C42030 NOR2X1_LOC_65/B NOR2X1_LOC_188/A 0.45fF
C42031 NAND2X1_LOC_35/Y INVX1_LOC_90/A 0.07fF
C42032 NOR2X1_LOC_240/a_36_216# NAND2X1_LOC_359/Y 0.00fF
C42033 INVX1_LOC_91/A NAND2X1_LOC_470/B 0.06fF
C42034 NAND2X1_LOC_754/a_36_24# INVX1_LOC_24/Y 0.00fF
C42035 NOR2X1_LOC_78/A INVX1_LOC_94/Y 0.03fF
C42036 INVX1_LOC_9/Y NOR2X1_LOC_361/B 0.08fF
C42037 NOR2X1_LOC_160/B INVX1_LOC_196/A 0.21fF
C42038 NOR2X1_LOC_303/Y INVX1_LOC_71/A 0.07fF
C42039 INVX1_LOC_27/A INVX1_LOC_135/A 0.68fF
C42040 NOR2X1_LOC_735/Y NOR2X1_LOC_665/Y 0.02fF
C42041 NOR2X1_LOC_584/Y INVX1_LOC_77/Y 0.29fF
C42042 NOR2X1_LOC_824/A INVX1_LOC_135/A 0.10fF
C42043 NOR2X1_LOC_468/Y NOR2X1_LOC_391/A 0.03fF
C42044 INVX1_LOC_72/Y INVX1_LOC_8/A 0.02fF
C42045 NOR2X1_LOC_52/Y NOR2X1_LOC_52/B 0.19fF
C42046 INVX1_LOC_45/Y INVX1_LOC_155/Y 0.03fF
C42047 NOR2X1_LOC_816/A NOR2X1_LOC_165/Y 0.05fF
C42048 INVX1_LOC_45/A INVX1_LOC_54/Y 0.03fF
C42049 NOR2X1_LOC_287/A NOR2X1_LOC_160/B 0.01fF
C42050 NAND2X1_LOC_567/Y NOR2X1_LOC_577/Y 0.01fF
C42051 NOR2X1_LOC_570/a_36_216# INVX1_LOC_104/A 0.00fF
C42052 NOR2X1_LOC_272/Y INPUT_1 0.04fF
C42053 INVX1_LOC_34/A NAND2X1_LOC_79/Y 0.03fF
C42054 NOR2X1_LOC_667/A INVX1_LOC_286/Y 0.10fF
C42055 INVX1_LOC_36/A NAND2X1_LOC_353/a_36_24# 0.01fF
C42056 INVX1_LOC_304/Y INVX1_LOC_217/A 0.11fF
C42057 NAND2X1_LOC_642/Y NOR2X1_LOC_301/A 0.03fF
C42058 INVX1_LOC_27/A NOR2X1_LOC_560/A 0.02fF
C42059 INVX1_LOC_35/A NOR2X1_LOC_196/Y 0.01fF
C42060 INVX1_LOC_191/Y INVX1_LOC_30/A 0.05fF
C42061 INVX1_LOC_54/Y NOR2X1_LOC_568/A 0.18fF
C42062 INVX1_LOC_278/A NOR2X1_LOC_74/A 0.00fF
C42063 INVX1_LOC_284/Y NAND2X1_LOC_835/a_36_24# 0.01fF
C42064 INVX1_LOC_248/A INVX1_LOC_286/Y 0.10fF
C42065 D_INPUT_0 NOR2X1_LOC_235/a_36_216# 0.00fF
C42066 NOR2X1_LOC_392/B INVX1_LOC_94/A 0.07fF
C42067 INVX1_LOC_223/Y NOR2X1_LOC_703/A 0.99fF
C42068 NAND2X1_LOC_787/A INVX1_LOC_6/A 0.03fF
C42069 INVX1_LOC_2/A NAND2X1_LOC_364/A 0.10fF
C42070 INVX1_LOC_93/A INVX1_LOC_102/Y -0.09fF
C42071 INVX1_LOC_1/A NOR2X1_LOC_150/a_36_216# 0.01fF
C42072 INVX1_LOC_278/A NOR2X1_LOC_9/Y 0.24fF
C42073 NOR2X1_LOC_78/A NOR2X1_LOC_621/a_36_216# 0.00fF
C42074 NOR2X1_LOC_634/A INVX1_LOC_19/A 0.02fF
C42075 NAND2X1_LOC_363/B INVX1_LOC_6/A 0.04fF
C42076 NAND2X1_LOC_472/Y INVX1_LOC_4/A 0.07fF
C42077 NOR2X1_LOC_15/Y NAND2X1_LOC_622/a_36_24# 0.00fF
C42078 NOR2X1_LOC_226/A NAND2X1_LOC_364/A 2.79fF
C42079 INVX1_LOC_41/A INVX1_LOC_33/A 0.13fF
C42080 NAND2X1_LOC_53/Y INVX1_LOC_83/A 0.24fF
C42081 INVX1_LOC_77/A NOR2X1_LOC_6/B 0.00fF
C42082 INVX1_LOC_203/A NOR2X1_LOC_649/B 0.10fF
C42083 INVX1_LOC_12/A INVX1_LOC_92/A 0.12fF
C42084 NOR2X1_LOC_82/A NOR2X1_LOC_76/A 0.07fF
C42085 INVX1_LOC_54/Y INVX1_LOC_71/A 0.15fF
C42086 INVX1_LOC_251/Y INVX1_LOC_314/Y 0.09fF
C42087 INVX1_LOC_55/Y NOR2X1_LOC_205/Y 0.06fF
C42088 NOR2X1_LOC_384/Y NAND2X1_LOC_859/B 0.01fF
C42089 INVX1_LOC_304/Y NAND2X1_LOC_787/B 0.32fF
C42090 NAND2X1_LOC_859/Y INVX1_LOC_30/A 0.01fF
C42091 NOR2X1_LOC_208/Y NOR2X1_LOC_357/a_36_216# 0.00fF
C42092 NOR2X1_LOC_791/Y INVX1_LOC_6/A 0.02fF
C42093 NOR2X1_LOC_307/Y INVX1_LOC_117/A 0.02fF
C42094 INVX1_LOC_269/A INVX1_LOC_182/Y 0.00fF
C42095 INVX1_LOC_123/A INVX1_LOC_306/Y 0.01fF
C42096 INVX1_LOC_136/A NOR2X1_LOC_690/Y 0.01fF
C42097 INVX1_LOC_47/A NOR2X1_LOC_160/B 0.02fF
C42098 INVX1_LOC_181/Y INVX1_LOC_53/Y 1.28fF
C42099 NOR2X1_LOC_176/Y NOR2X1_LOC_438/Y 0.00fF
C42100 INVX1_LOC_206/A NOR2X1_LOC_388/Y 0.01fF
C42101 NAND2X1_LOC_656/A INVX1_LOC_232/A 0.10fF
C42102 VDD INVX1_LOC_173/A -0.00fF
C42103 INVX1_LOC_300/A INVX1_LOC_300/Y 0.09fF
C42104 INVX1_LOC_33/A INVX1_LOC_64/Y 1.44fF
C42105 NOR2X1_LOC_533/Y NAND2X1_LOC_740/B 0.02fF
C42106 NAND2X1_LOC_711/B NOR2X1_LOC_701/Y 0.07fF
C42107 INVX1_LOC_21/A NOR2X1_LOC_337/Y 0.17fF
C42108 INVX1_LOC_24/A NOR2X1_LOC_589/A 0.16fF
C42109 INVX1_LOC_53/A NOR2X1_LOC_850/a_36_216# 0.00fF
C42110 INVX1_LOC_14/Y INVX1_LOC_29/Y 0.01fF
C42111 INVX1_LOC_85/A INVX1_LOC_96/Y 0.00fF
C42112 INVX1_LOC_104/A NOR2X1_LOC_493/B 0.07fF
C42113 INVX1_LOC_30/A NAND2X1_LOC_866/B 1.35fF
C42114 INVX1_LOC_256/A INVX1_LOC_79/A 0.10fF
C42115 GATE_222 NOR2X1_LOC_814/A 0.02fF
C42116 INVX1_LOC_19/A INVX1_LOC_29/A 0.73fF
C42117 INVX1_LOC_30/Y INVX1_LOC_77/A 0.03fF
C42118 INVX1_LOC_45/A NOR2X1_LOC_112/Y 0.01fF
C42119 INVX1_LOC_30/A NAND2X1_LOC_807/Y 0.10fF
C42120 INVX1_LOC_142/Y INVX1_LOC_85/Y 0.01fF
C42121 INVX1_LOC_41/A NAND2X1_LOC_754/a_36_24# 0.01fF
C42122 NOR2X1_LOC_590/A INVX1_LOC_75/A 0.11fF
C42123 NOR2X1_LOC_443/a_36_216# INPUT_0 0.00fF
C42124 NOR2X1_LOC_226/A NAND2X1_LOC_785/A 0.52fF
C42125 INVX1_LOC_256/Y INVX1_LOC_168/A 0.37fF
C42126 NAND2X1_LOC_726/a_36_24# INVX1_LOC_28/A 0.00fF
C42127 INVX1_LOC_21/A NOR2X1_LOC_56/Y 0.07fF
C42128 INVX1_LOC_21/A NAND2X1_LOC_659/B 0.07fF
C42129 INVX1_LOC_299/A NOR2X1_LOC_78/A 0.03fF
C42130 INVX1_LOC_17/A NAND2X1_LOC_669/a_36_24# 0.01fF
C42131 INVX1_LOC_3/Y INVX1_LOC_63/A 0.14fF
C42132 INVX1_LOC_198/Y INVX1_LOC_85/Y 0.05fF
C42133 NOR2X1_LOC_510/Y NOR2X1_LOC_173/a_36_216# 0.00fF
C42134 INVX1_LOC_35/A INVX1_LOC_33/Y 0.04fF
C42135 NOR2X1_LOC_168/Y NOR2X1_LOC_356/A 0.01fF
C42136 INVX1_LOC_2/A NOR2X1_LOC_289/a_36_216# 0.00fF
C42137 INVX1_LOC_13/A INVX1_LOC_82/A 0.36fF
C42138 NAND2X1_LOC_725/B NOR2X1_LOC_396/Y 0.21fF
C42139 NOR2X1_LOC_621/A NOR2X1_LOC_624/B 0.05fF
C42140 NOR2X1_LOC_538/B NOR2X1_LOC_78/A 0.00fF
C42141 NAND2X1_LOC_574/A NAND2X1_LOC_223/A 0.02fF
C42142 INVX1_LOC_26/Y NOR2X1_LOC_634/A 0.38fF
C42143 NAND2X1_LOC_167/a_36_24# NOR2X1_LOC_703/A 0.00fF
C42144 NOR2X1_LOC_489/A INVX1_LOC_129/A 0.06fF
C42145 INVX1_LOC_21/A INVX1_LOC_146/Y 0.01fF
C42146 INVX1_LOC_172/A NAND2X1_LOC_862/Y 0.06fF
C42147 INVX1_LOC_256/A INVX1_LOC_91/A 0.47fF
C42148 INVX1_LOC_21/A VDD 2.24fF
C42149 INVX1_LOC_4/A NAND2X1_LOC_773/B 0.07fF
C42150 NOR2X1_LOC_340/Y NOR2X1_LOC_99/B 0.02fF
C42151 NAND2X1_LOC_474/Y INVX1_LOC_46/A 1.46fF
C42152 NOR2X1_LOC_78/B NOR2X1_LOC_500/Y 0.07fF
C42153 INVX1_LOC_292/A NOR2X1_LOC_355/B 0.09fF
C42154 INVX1_LOC_17/A NAND2X1_LOC_642/Y 0.06fF
C42155 NAND2X1_LOC_214/B NOR2X1_LOC_813/Y 0.02fF
C42156 INVX1_LOC_27/A INVX1_LOC_139/Y 0.05fF
C42157 INVX1_LOC_32/A NAND2X1_LOC_81/B 0.16fF
C42158 INVX1_LOC_226/Y NOR2X1_LOC_78/B 0.03fF
C42159 INVX1_LOC_293/A NOR2X1_LOC_78/A 0.03fF
C42160 NOR2X1_LOC_430/A INVX1_LOC_244/A 0.22fF
C42161 NAND2X1_LOC_35/Y INVX1_LOC_38/A 0.07fF
C42162 INVX1_LOC_2/A NOR2X1_LOC_86/A 0.09fF
C42163 NOR2X1_LOC_67/A INVX1_LOC_16/A 1.52fF
C42164 NOR2X1_LOC_664/Y INVX1_LOC_135/A 0.27fF
C42165 INVX1_LOC_30/A INVX1_LOC_6/A 1.21fF
C42166 NOR2X1_LOC_473/B INVX1_LOC_67/A 0.03fF
C42167 NAND2X1_LOC_564/a_36_24# NOR2X1_LOC_71/Y -0.01fF
C42168 NOR2X1_LOC_479/B INVX1_LOC_84/Y 0.02fF
C42169 NOR2X1_LOC_554/B NOR2X1_LOC_188/A 0.03fF
C42170 NOR2X1_LOC_753/Y INVX1_LOC_28/A 0.03fF
C42171 NOR2X1_LOC_453/Y VDD 0.28fF
C42172 NOR2X1_LOC_843/A NOR2X1_LOC_174/B 0.76fF
C42173 NAND2X1_LOC_214/B INVX1_LOC_280/A 0.12fF
C42174 NOR2X1_LOC_598/B INVX1_LOC_108/A 0.02fF
C42175 NOR2X1_LOC_281/Y NOR2X1_LOC_653/Y 0.05fF
C42176 NOR2X1_LOC_332/A NOR2X1_LOC_87/B 0.09fF
C42177 INVX1_LOC_34/A D_GATE_366 0.50fF
C42178 INVX1_LOC_297/Y INVX1_LOC_300/A 0.24fF
C42179 INVX1_LOC_69/Y NOR2X1_LOC_703/B 0.01fF
C42180 NOR2X1_LOC_82/Y INVX1_LOC_25/Y 0.02fF
C42181 INVX1_LOC_89/A INVX1_LOC_104/A 0.07fF
C42182 NOR2X1_LOC_205/Y NOR2X1_LOC_357/Y 0.10fF
C42183 INVX1_LOC_53/A INVX1_LOC_307/A 0.14fF
C42184 INVX1_LOC_128/Y INVX1_LOC_272/A 0.28fF
C42185 NOR2X1_LOC_160/B INVX1_LOC_95/Y 0.34fF
C42186 INPUT_3 INVX1_LOC_316/A 0.08fF
C42187 INVX1_LOC_34/A NOR2X1_LOC_750/A 0.01fF
C42188 INVX1_LOC_50/Y INVX1_LOC_9/A 0.03fF
C42189 NOR2X1_LOC_78/B INVX1_LOC_10/A 0.07fF
C42190 INVX1_LOC_24/A INVX1_LOC_222/A 0.05fF
C42191 NAND2X1_LOC_112/Y NOR2X1_LOC_321/a_36_216# 0.00fF
C42192 NOR2X1_LOC_524/Y NOR2X1_LOC_78/A 0.05fF
C42193 INVX1_LOC_53/A NOR2X1_LOC_445/B 0.23fF
C42194 INVX1_LOC_27/A INVX1_LOC_280/A 0.07fF
C42195 INVX1_LOC_298/Y INVX1_LOC_19/A 0.03fF
C42196 INVX1_LOC_54/Y NOR2X1_LOC_123/B 0.01fF
C42197 NOR2X1_LOC_262/Y NOR2X1_LOC_74/A 0.02fF
C42198 NAND2X1_LOC_571/Y INVX1_LOC_38/A 0.07fF
C42199 NAND2X1_LOC_475/Y INVX1_LOC_270/A 0.10fF
C42200 NOR2X1_LOC_655/B NOR2X1_LOC_99/B 0.10fF
C42201 NOR2X1_LOC_577/Y INVX1_LOC_67/Y 0.00fF
C42202 NOR2X1_LOC_197/A INVX1_LOC_76/A 0.02fF
C42203 NAND2X1_LOC_53/Y INVX1_LOC_46/A 0.26fF
C42204 NAND2X1_LOC_729/a_36_24# INVX1_LOC_240/A 0.01fF
C42205 INVX1_LOC_233/Y INVX1_LOC_260/A 0.04fF
C42206 NAND2X1_LOC_803/B NAND2X1_LOC_453/A 0.02fF
C42207 NOR2X1_LOC_272/Y INVX1_LOC_118/A 0.10fF
C42208 INVX1_LOC_257/A NAND2X1_LOC_628/a_36_24# 0.02fF
C42209 INVX1_LOC_83/A NOR2X1_LOC_374/a_36_216# 0.00fF
C42210 INVX1_LOC_171/A INVX1_LOC_143/A 0.00fF
C42211 INVX1_LOC_284/Y NOR2X1_LOC_824/Y 0.03fF
C42212 NAND2X1_LOC_741/B INPUT_4 0.14fF
C42213 NOR2X1_LOC_598/B NOR2X1_LOC_801/A 0.40fF
C42214 NOR2X1_LOC_172/Y INVX1_LOC_144/A 0.01fF
C42215 INVX1_LOC_283/Y INVX1_LOC_311/A 0.01fF
C42216 INVX1_LOC_109/A NAND2X1_LOC_61/Y 0.04fF
C42217 INVX1_LOC_236/Y INVX1_LOC_76/A 0.00fF
C42218 NOR2X1_LOC_590/A NOR2X1_LOC_309/a_36_216# 0.00fF
C42219 INVX1_LOC_26/Y INVX1_LOC_29/A 0.07fF
C42220 INVX1_LOC_58/A INVX1_LOC_63/A 0.00fF
C42221 NOR2X1_LOC_240/Y NOR2X1_LOC_240/A 0.01fF
C42222 INVX1_LOC_284/Y INVX1_LOC_76/A 2.54fF
C42223 NOR2X1_LOC_428/Y VDD 0.12fF
C42224 NAND2X1_LOC_555/Y D_GATE_662 0.01fF
C42225 NOR2X1_LOC_781/Y INVX1_LOC_91/A 0.01fF
C42226 NOR2X1_LOC_590/A NAND2X1_LOC_453/A 0.08fF
C42227 INVX1_LOC_266/A INVX1_LOC_9/A 0.19fF
C42228 INVX1_LOC_276/A INVX1_LOC_28/A 0.07fF
C42229 INVX1_LOC_32/A INVX1_LOC_4/Y 0.29fF
C42230 NOR2X1_LOC_639/a_36_216# INVX1_LOC_290/A 0.00fF
C42231 NOR2X1_LOC_68/A NOR2X1_LOC_545/B 0.02fF
C42232 NAND2X1_LOC_579/A INVX1_LOC_54/A 0.10fF
C42233 INVX1_LOC_166/A INVX1_LOC_29/A 0.05fF
C42234 NOR2X1_LOC_158/Y D_INPUT_5 0.04fF
C42235 NOR2X1_LOC_648/a_36_216# INVX1_LOC_182/Y 0.00fF
C42236 NOR2X1_LOC_392/B NOR2X1_LOC_83/Y 0.04fF
C42237 NOR2X1_LOC_191/A NAND2X1_LOC_850/A 0.13fF
C42238 NOR2X1_LOC_242/A NOR2X1_LOC_445/B 0.00fF
C42239 NOR2X1_LOC_738/A NOR2X1_LOC_731/Y 0.18fF
C42240 INVX1_LOC_83/A INVX1_LOC_10/A 0.10fF
C42241 INVX1_LOC_135/A INVX1_LOC_234/A 1.33fF
C42242 INVX1_LOC_87/Y INVX1_LOC_22/A 0.01fF
C42243 NAND2X1_LOC_354/Y INVX1_LOC_146/Y 0.00fF
C42244 INVX1_LOC_24/A INVX1_LOC_147/Y 0.20fF
C42245 NOR2X1_LOC_517/Y VDD 0.12fF
C42246 NAND2X1_LOC_589/a_36_24# NAND2X1_LOC_453/A 0.00fF
C42247 NOR2X1_LOC_688/Y INVX1_LOC_117/A 0.04fF
C42248 NAND2X1_LOC_354/Y VDD 0.19fF
C42249 INVX1_LOC_104/A NOR2X1_LOC_703/Y 0.08fF
C42250 INVX1_LOC_49/A NOR2X1_LOC_405/A 0.08fF
C42251 NOR2X1_LOC_520/A INPUT_0 0.01fF
C42252 INVX1_LOC_53/A INVX1_LOC_12/A 0.33fF
C42253 INVX1_LOC_24/A INVX1_LOC_20/A 0.18fF
C42254 NOR2X1_LOC_582/Y VDD 0.26fF
C42255 INVX1_LOC_5/A NAND2X1_LOC_219/B -0.00fF
C42256 INVX1_LOC_308/A NAND2X1_LOC_807/B 0.01fF
C42257 NOR2X1_LOC_160/B NAND2X1_LOC_289/a_36_24# 0.00fF
C42258 NOR2X1_LOC_773/Y NOR2X1_LOC_527/Y 0.04fF
C42259 NOR2X1_LOC_315/Y INVX1_LOC_98/A 0.02fF
C42260 NOR2X1_LOC_315/Y NOR2X1_LOC_78/A 0.04fF
C42261 NOR2X1_LOC_103/Y INVX1_LOC_35/Y 0.28fF
C42262 INVX1_LOC_88/A NOR2X1_LOC_697/Y 1.18fF
C42263 INVX1_LOC_249/A INVX1_LOC_139/Y 0.00fF
C42264 INVX1_LOC_49/A NOR2X1_LOC_857/A 0.07fF
C42265 NAND2X1_LOC_348/A NOR2X1_LOC_572/a_36_216# 0.00fF
C42266 INVX1_LOC_21/A INVX1_LOC_133/A 0.03fF
C42267 INVX1_LOC_310/A NOR2X1_LOC_78/A 0.01fF
C42268 INVX1_LOC_135/A NOR2X1_LOC_19/B 0.66fF
C42269 NOR2X1_LOC_181/Y INVX1_LOC_247/A 0.01fF
C42270 NAND2X1_LOC_331/a_36_24# INVX1_LOC_28/A 0.01fF
C42271 INVX1_LOC_227/A INVX1_LOC_75/A 0.17fF
C42272 INVX1_LOC_2/A NOR2X1_LOC_405/A 0.05fF
C42273 INVX1_LOC_15/A NOR2X1_LOC_342/A 0.01fF
C42274 INVX1_LOC_30/A NOR2X1_LOC_79/A 0.04fF
C42275 NOR2X1_LOC_391/Y NOR2X1_LOC_719/A 0.15fF
C42276 NAND2X1_LOC_391/Y NOR2X1_LOC_89/A 0.03fF
C42277 NOR2X1_LOC_500/B NOR2X1_LOC_640/Y 0.13fF
C42278 NOR2X1_LOC_321/Y NAND2X1_LOC_74/B 0.07fF
C42279 NOR2X1_LOC_52/B NOR2X1_LOC_603/Y 0.04fF
C42280 NOR2X1_LOC_226/A NOR2X1_LOC_405/A 0.00fF
C42281 INVX1_LOC_50/Y NOR2X1_LOC_861/Y 0.07fF
C42282 NOR2X1_LOC_315/Y NAND2X1_LOC_464/A 0.01fF
C42283 INVX1_LOC_245/Y INVX1_LOC_84/A 0.03fF
C42284 NOR2X1_LOC_303/Y NOR2X1_LOC_331/B 0.07fF
C42285 NOR2X1_LOC_577/Y NOR2X1_LOC_366/a_36_216# 0.00fF
C42286 NOR2X1_LOC_690/A INVX1_LOC_37/Y 0.01fF
C42287 NAND2X1_LOC_785/Y VDD 0.09fF
C42288 NOR2X1_LOC_778/B INVX1_LOC_247/A 0.00fF
C42289 INVX1_LOC_57/A NOR2X1_LOC_318/A 0.01fF
C42290 INVX1_LOC_215/Y INVX1_LOC_63/A 0.15fF
C42291 NOR2X1_LOC_490/Y NOR2X1_LOC_19/B 0.01fF
C42292 NOR2X1_LOC_68/A NOR2X1_LOC_156/a_36_216# 0.00fF
C42293 INVX1_LOC_200/Y NOR2X1_LOC_693/Y 0.01fF
C42294 INVX1_LOC_143/A INVX1_LOC_20/A 0.00fF
C42295 INVX1_LOC_50/A NOR2X1_LOC_383/B 0.06fF
C42296 NOR2X1_LOC_273/Y NOR2X1_LOC_433/Y 0.05fF
C42297 NAND2X1_LOC_276/Y NOR2X1_LOC_536/A 0.00fF
C42298 INPUT_0 INVX1_LOC_65/Y 0.12fF
C42299 INVX1_LOC_90/A INVX1_LOC_144/A 0.10fF
C42300 NAND2X1_LOC_326/A INVX1_LOC_42/A 0.01fF
C42301 NOR2X1_LOC_675/A INVX1_LOC_53/Y 0.00fF
C42302 NOR2X1_LOC_15/Y INVX1_LOC_290/Y 0.07fF
C42303 INVX1_LOC_90/A NOR2X1_LOC_83/Y 0.14fF
C42304 INVX1_LOC_75/A NOR2X1_LOC_703/A 0.02fF
C42305 NAND2X1_LOC_579/A NOR2X1_LOC_48/B 0.01fF
C42306 NAND2X1_LOC_793/Y NAND2X1_LOC_74/B 0.03fF
C42307 NOR2X1_LOC_334/Y NOR2X1_LOC_674/a_36_216# 0.00fF
C42308 INVX1_LOC_214/A VDD -0.00fF
C42309 INVX1_LOC_161/Y INVX1_LOC_29/A 0.07fF
C42310 INVX1_LOC_50/A NAND2X1_LOC_738/B 0.04fF
C42311 INVX1_LOC_35/A INVX1_LOC_23/Y 0.03fF
C42312 NOR2X1_LOC_667/A VDD 0.84fF
C42313 INVX1_LOC_71/A NAND2X1_LOC_656/B 0.06fF
C42314 NOR2X1_LOC_664/Y INVX1_LOC_280/A 0.16fF
C42315 INVX1_LOC_36/A NAND2X1_LOC_475/Y 0.11fF
C42316 INVX1_LOC_250/A INVX1_LOC_250/Y 0.01fF
C42317 INVX1_LOC_135/A NOR2X1_LOC_528/Y 0.01fF
C42318 INVX1_LOC_248/A VDD 0.12fF
C42319 INVX1_LOC_35/A NOR2X1_LOC_342/B 0.01fF
C42320 NOR2X1_LOC_186/Y INVX1_LOC_94/Y 0.26fF
C42321 NAND2X1_LOC_650/B INVX1_LOC_25/Y 0.07fF
C42322 INVX1_LOC_280/Y NAND2X1_LOC_804/Y 0.46fF
C42323 NOR2X1_LOC_68/A INVX1_LOC_119/Y 0.02fF
C42324 NAND2X1_LOC_276/Y NOR2X1_LOC_655/Y 0.00fF
C42325 NOR2X1_LOC_500/Y INVX1_LOC_46/A 0.07fF
C42326 NOR2X1_LOC_6/B INVX1_LOC_9/A 0.17fF
C42327 INVX1_LOC_279/A NOR2X1_LOC_275/A 0.02fF
C42328 INVX1_LOC_226/Y INVX1_LOC_46/A 0.01fF
C42329 INVX1_LOC_90/A NOR2X1_LOC_845/A 0.19fF
C42330 INVX1_LOC_226/Y NOR2X1_LOC_98/A -0.01fF
C42331 NAND2X1_LOC_72/Y NOR2X1_LOC_383/B 0.00fF
C42332 NAND2X1_LOC_276/Y NAND2X1_LOC_93/B 0.04fF
C42333 NOR2X1_LOC_719/B INVX1_LOC_59/Y 0.01fF
C42334 INVX1_LOC_83/A NOR2X1_LOC_711/Y 0.23fF
C42335 INVX1_LOC_235/A NOR2X1_LOC_415/Y 0.01fF
C42336 INVX1_LOC_290/A NAND2X1_LOC_39/Y 0.03fF
C42337 INVX1_LOC_269/A NOR2X1_LOC_38/B 0.05fF
C42338 NAND2X1_LOC_390/A NAND2X1_LOC_641/a_36_24# 0.00fF
C42339 INVX1_LOC_30/A NOR2X1_LOC_633/A 0.00fF
C42340 NOR2X1_LOC_525/Y NOR2X1_LOC_824/Y 0.04fF
C42341 NOR2X1_LOC_521/Y VDD 0.00fF
C42342 NOR2X1_LOC_130/A INVX1_LOC_147/Y 0.06fF
C42343 NOR2X1_LOC_147/B NOR2X1_LOC_155/A 0.03fF
C42344 NAND2X1_LOC_218/B NOR2X1_LOC_814/A 0.77fF
C42345 NOR2X1_LOC_208/Y NAND2X1_LOC_475/Y 0.02fF
C42346 NAND2X1_LOC_326/A INVX1_LOC_78/A 0.04fF
C42347 NAND2X1_LOC_783/A INVX1_LOC_20/A 0.01fF
C42348 NOR2X1_LOC_778/B NOR2X1_LOC_499/B 0.00fF
C42349 NOR2X1_LOC_419/Y INVX1_LOC_27/Y 0.04fF
C42350 NAND2X1_LOC_800/Y INVX1_LOC_20/A 0.01fF
C42351 NOR2X1_LOC_341/a_36_216# INVX1_LOC_63/A 0.01fF
C42352 INVX1_LOC_1/Y INVX1_LOC_117/A 0.01fF
C42353 NOR2X1_LOC_136/Y INVX1_LOC_38/A 0.03fF
C42354 NAND2X1_LOC_364/A NAND2X1_LOC_63/Y 0.01fF
C42355 NAND2X1_LOC_347/B NOR2X1_LOC_316/a_36_216# 0.00fF
C42356 INVX1_LOC_10/A INVX1_LOC_46/A 0.13fF
C42357 NOR2X1_LOC_525/Y INVX1_LOC_76/A 0.03fF
C42358 VDD NOR2X1_LOC_565/B 0.26fF
C42359 NOR2X1_LOC_130/A INVX1_LOC_20/A 0.05fF
C42360 INVX1_LOC_34/A INVX1_LOC_123/Y 0.01fF
C42361 NAND2X1_LOC_402/B INVX1_LOC_242/A 0.02fF
C42362 NAND2X1_LOC_11/Y INVX1_LOC_118/A 0.03fF
C42363 D_INPUT_0 NOR2X1_LOC_825/Y 0.03fF
C42364 NAND2X1_LOC_347/B INVX1_LOC_26/A 0.01fF
C42365 D_INPUT_1 INVX1_LOC_306/Y 1.01fF
C42366 NOR2X1_LOC_399/Y NOR2X1_LOC_629/Y 0.00fF
C42367 NAND2X1_LOC_276/Y NOR2X1_LOC_649/B 0.01fF
C42368 INVX1_LOC_5/A INVX1_LOC_58/Y 0.07fF
C42369 NOR2X1_LOC_68/A INVX1_LOC_284/A 0.26fF
C42370 NAND2X1_LOC_276/Y INVX1_LOC_3/A 4.09fF
C42371 NOR2X1_LOC_65/B NAND2X1_LOC_326/A 0.14fF
C42372 NOR2X1_LOC_13/Y INVX1_LOC_272/A 0.10fF
C42373 NOR2X1_LOC_690/A NOR2X1_LOC_485/Y 0.01fF
C42374 INPUT_5 NOR2X1_LOC_694/Y 0.01fF
C42375 NOR2X1_LOC_518/a_36_216# INVX1_LOC_102/A 0.01fF
C42376 INPUT_3 INVX1_LOC_4/Y 0.06fF
C42377 NOR2X1_LOC_78/B INVX1_LOC_307/A 0.13fF
C42378 NOR2X1_LOC_473/B NOR2X1_LOC_137/Y 0.16fF
C42379 NOR2X1_LOC_778/B NOR2X1_LOC_862/B 0.01fF
C42380 INVX1_LOC_30/Y INVX1_LOC_9/A 0.05fF
C42381 NOR2X1_LOC_634/B NOR2X1_LOC_445/B 0.16fF
C42382 NAND2X1_LOC_660/A NOR2X1_LOC_841/A 0.10fF
C42383 NOR2X1_LOC_309/Y NAND2X1_LOC_475/Y 0.01fF
C42384 INVX1_LOC_70/Y INVX1_LOC_100/A 0.97fF
C42385 NAND2X1_LOC_323/B NOR2X1_LOC_461/A 0.07fF
C42386 INVX1_LOC_234/A INVX1_LOC_280/A 0.80fF
C42387 NOR2X1_LOC_703/B NOR2X1_LOC_170/A 0.14fF
C42388 INVX1_LOC_69/Y INVX1_LOC_91/A 1.61fF
C42389 NOR2X1_LOC_78/B NOR2X1_LOC_445/B 0.01fF
C42390 INVX1_LOC_234/A NOR2X1_LOC_94/Y 0.05fF
C42391 NOR2X1_LOC_740/Y NOR2X1_LOC_727/B 0.04fF
C42392 NOR2X1_LOC_788/a_36_216# INVX1_LOC_91/A 0.00fF
C42393 NAND2X1_LOC_338/B NOR2X1_LOC_49/a_36_216# 0.00fF
C42394 INVX1_LOC_8/A INVX1_LOC_19/A 0.06fF
C42395 INVX1_LOC_121/A NAND2X1_LOC_459/a_36_24# 0.00fF
C42396 NAND2X1_LOC_175/B INVX1_LOC_272/A 0.03fF
C42397 NOR2X1_LOC_364/A INVX1_LOC_22/A 1.15fF
C42398 NOR2X1_LOC_725/A INVX1_LOC_91/A 0.02fF
C42399 NOR2X1_LOC_816/A NOR2X1_LOC_654/A 0.10fF
C42400 NOR2X1_LOC_666/Y NOR2X1_LOC_678/A 0.12fF
C42401 INVX1_LOC_72/A NAND2X1_LOC_454/Y 0.08fF
C42402 NAND2X1_LOC_51/B VDD 0.99fF
C42403 NOR2X1_LOC_543/a_36_216# INVX1_LOC_91/A 0.01fF
C42404 NOR2X1_LOC_19/B NOR2X1_LOC_813/Y 0.00fF
C42405 NOR2X1_LOC_201/A INVX1_LOC_110/Y 0.11fF
C42406 INVX1_LOC_24/A INVX1_LOC_4/A 0.03fF
C42407 INVX1_LOC_21/A NOR2X1_LOC_510/Y 0.03fF
C42408 INVX1_LOC_154/A NOR2X1_LOC_349/A 0.12fF
C42409 INVX1_LOC_34/A INVX1_LOC_102/A 0.09fF
C42410 NOR2X1_LOC_147/B NOR2X1_LOC_833/B 0.03fF
C42411 NOR2X1_LOC_724/Y NOR2X1_LOC_499/B 0.05fF
C42412 NAND2X1_LOC_860/A NOR2X1_LOC_103/Y 0.02fF
C42413 NOR2X1_LOC_272/Y INVX1_LOC_39/A 0.02fF
C42414 NOR2X1_LOC_391/Y INVX1_LOC_76/A -0.01fF
C42415 NAND2X1_LOC_808/A INVX1_LOC_92/A 0.07fF
C42416 NOR2X1_LOC_261/Y INVX1_LOC_245/Y 0.16fF
C42417 NOR2X1_LOC_19/B INVX1_LOC_280/A 0.12fF
C42418 NOR2X1_LOC_191/B NOR2X1_LOC_248/A 0.13fF
C42419 INVX1_LOC_22/A NOR2X1_LOC_814/A 0.07fF
C42420 NOR2X1_LOC_705/B NOR2X1_LOC_598/B 0.03fF
C42421 NOR2X1_LOC_91/Y NOR2X1_LOC_301/A 0.00fF
C42422 INVX1_LOC_135/A NOR2X1_LOC_216/B 0.07fF
C42423 INVX1_LOC_30/A INVX1_LOC_270/A 0.10fF
C42424 INVX1_LOC_83/A NOR2X1_LOC_445/B 0.05fF
C42425 INVX1_LOC_304/A NOR2X1_LOC_123/a_36_216# 0.00fF
C42426 INVX1_LOC_57/Y INVX1_LOC_50/A 0.08fF
C42427 NOR2X1_LOC_557/Y INVX1_LOC_4/A 0.15fF
C42428 NOR2X1_LOC_78/B INVX1_LOC_12/A 1.67fF
C42429 NOR2X1_LOC_382/Y INVX1_LOC_23/A 0.03fF
C42430 NOR2X1_LOC_843/A NOR2X1_LOC_623/B 0.03fF
C42431 INVX1_LOC_90/A NOR2X1_LOC_155/A 0.05fF
C42432 NAND2X1_LOC_231/Y INVX1_LOC_102/A 0.06fF
C42433 INVX1_LOC_255/A NAND2X1_LOC_659/B 0.05fF
C42434 INVX1_LOC_144/A INVX1_LOC_38/A 0.08fF
C42435 NOR2X1_LOC_75/Y INVX1_LOC_5/A 0.03fF
C42436 INVX1_LOC_21/A NOR2X1_LOC_361/B 0.15fF
C42437 INVX1_LOC_303/A NAND2X1_LOC_221/a_36_24# 0.00fF
C42438 NOR2X1_LOC_481/A INVX1_LOC_94/Y 0.14fF
C42439 NOR2X1_LOC_389/B NOR2X1_LOC_155/A 0.00fF
C42440 INVX1_LOC_45/A NAND2X1_LOC_860/A 0.09fF
C42441 NOR2X1_LOC_836/B INVX1_LOC_37/A 0.18fF
C42442 INVX1_LOC_278/A INVX1_LOC_124/Y 0.28fF
C42443 NOR2X1_LOC_471/Y INVX1_LOC_204/Y 0.04fF
C42444 NOR2X1_LOC_681/Y NAND2X1_LOC_655/A 0.39fF
C42445 NAND2X1_LOC_863/A INVX1_LOC_185/A 0.01fF
C42446 D_INPUT_0 INVX1_LOC_84/A 0.81fF
C42447 NAND2X1_LOC_787/A INVX1_LOC_36/A 0.07fF
C42448 INVX1_LOC_37/A NAND2X1_LOC_655/A 0.07fF
C42449 INVX1_LOC_71/A NAND2X1_LOC_286/B 0.03fF
C42450 INVX1_LOC_50/A NOR2X1_LOC_512/Y 0.01fF
C42451 NOR2X1_LOC_495/Y NOR2X1_LOC_693/Y 0.02fF
C42452 NAND2X1_LOC_793/Y NAND2X1_LOC_793/a_36_24# 0.02fF
C42453 VDD INVX1_LOC_255/A 0.00fF
C42454 INVX1_LOC_269/A NOR2X1_LOC_468/Y 0.55fF
C42455 NOR2X1_LOC_218/Y INVX1_LOC_109/Y 0.04fF
C42456 INVX1_LOC_304/A VDD 0.80fF
C42457 NOR2X1_LOC_78/A NAND2X1_LOC_96/A 0.07fF
C42458 NOR2X1_LOC_332/A NAND2X1_LOC_219/B 0.21fF
C42459 INVX1_LOC_30/A NOR2X1_LOC_109/Y 0.10fF
C42460 INVX1_LOC_45/A NOR2X1_LOC_834/a_36_216# 0.00fF
C42461 NOR2X1_LOC_280/Y INVX1_LOC_20/A 0.20fF
C42462 INPUT_0 INVX1_LOC_70/A 0.31fF
C42463 NOR2X1_LOC_845/A INVX1_LOC_38/A -0.01fF
C42464 NAND2X1_LOC_665/a_36_24# INVX1_LOC_84/A 0.01fF
C42465 INVX1_LOC_143/A INVX1_LOC_4/A 0.32fF
C42466 VDD NOR2X1_LOC_670/Y 0.12fF
C42467 INVX1_LOC_37/A NOR2X1_LOC_683/Y 0.02fF
C42468 INVX1_LOC_96/A INVX1_LOC_9/A 0.05fF
C42469 INVX1_LOC_8/A INVX1_LOC_26/Y 0.99fF
C42470 NOR2X1_LOC_836/Y NOR2X1_LOC_852/Y 0.23fF
C42471 NOR2X1_LOC_335/A INVX1_LOC_57/A 0.00fF
C42472 NAND2X1_LOC_594/a_36_24# NOR2X1_LOC_441/Y 0.00fF
C42473 NOR2X1_LOC_506/a_36_216# NOR2X1_LOC_56/Y 0.00fF
C42474 NAND2X1_LOC_860/A INVX1_LOC_71/A 0.24fF
C42475 INVX1_LOC_62/A INVX1_LOC_29/A 0.01fF
C42476 NAND2X1_LOC_555/Y INVX1_LOC_239/A 0.67fF
C42477 NAND2X1_LOC_563/A NOR2X1_LOC_38/B 0.05fF
C42478 INVX1_LOC_36/A NOR2X1_LOC_791/Y 0.05fF
C42479 INVX1_LOC_83/A INVX1_LOC_12/A 0.10fF
C42480 NAND2X1_LOC_773/Y NOR2X1_LOC_160/B 0.10fF
C42481 INVX1_LOC_279/A NOR2X1_LOC_842/a_36_216# 0.00fF
C42482 INVX1_LOC_222/A NOR2X1_LOC_197/B 0.02fF
C42483 NOR2X1_LOC_391/B NOR2X1_LOC_216/B 0.00fF
C42484 NOR2X1_LOC_470/B INVX1_LOC_174/A 0.11fF
C42485 INVX1_LOC_41/A NOR2X1_LOC_748/A 0.31fF
C42486 INVX1_LOC_64/A INVX1_LOC_24/A 6.06fF
C42487 INPUT_0 INVX1_LOC_123/Y 0.03fF
C42488 NAND2X1_LOC_787/A NOR2X1_LOC_237/Y 0.01fF
C42489 NOR2X1_LOC_510/Y NAND2X1_LOC_354/Y 0.02fF
C42490 NOR2X1_LOC_267/A NOR2X1_LOC_791/Y 0.01fF
C42491 NOR2X1_LOC_33/A INVX1_LOC_15/A 0.01fF
C42492 NOR2X1_LOC_405/A INVX1_LOC_118/A 0.07fF
C42493 NAND2X1_LOC_660/Y INVX1_LOC_15/A 0.03fF
C42494 INVX1_LOC_37/A NAND2X1_LOC_51/a_36_24# 0.02fF
C42495 NOR2X1_LOC_667/Y NAND2X1_LOC_538/Y 0.13fF
C42496 INVX1_LOC_208/A INVX1_LOC_271/Y 0.10fF
C42497 D_INPUT_1 INVX1_LOC_294/Y 0.01fF
C42498 NAND2X1_LOC_848/A NOR2X1_LOC_825/Y 0.01fF
C42499 NOR2X1_LOC_78/B NOR2X1_LOC_686/A 0.04fF
C42500 NOR2X1_LOC_516/B INVX1_LOC_271/Y 0.01fF
C42501 NOR2X1_LOC_598/B NOR2X1_LOC_147/B 0.09fF
C42502 INVX1_LOC_266/A NOR2X1_LOC_169/B 0.03fF
C42503 NAND2X1_LOC_468/B INVX1_LOC_157/Y -0.00fF
C42504 INVX1_LOC_5/A NOR2X1_LOC_419/Y 0.03fF
C42505 INVX1_LOC_45/A NAND2X1_LOC_537/Y 0.01fF
C42506 NAND2X1_LOC_787/A NOR2X1_LOC_309/Y 0.10fF
C42507 NAND2X1_LOC_552/A NOR2X1_LOC_716/B 0.01fF
C42508 D_INPUT_0 INVX1_LOC_15/A 0.21fF
C42509 NAND2X1_LOC_537/Y NAND2X1_LOC_856/A 0.00fF
C42510 INVX1_LOC_5/A NOR2X1_LOC_716/B 0.06fF
C42511 NAND2X1_LOC_794/B NOR2X1_LOC_753/Y 0.07fF
C42512 INVX1_LOC_35/A NAND2X1_LOC_116/A 0.05fF
C42513 NOR2X1_LOC_791/B INVX1_LOC_14/A 0.02fF
C42514 INVX1_LOC_36/A NOR2X1_LOC_457/A 0.03fF
C42515 INVX1_LOC_58/A NOR2X1_LOC_362/a_36_216# 0.00fF
C42516 NOR2X1_LOC_773/Y NOR2X1_LOC_654/A 0.02fF
C42517 INVX1_LOC_110/Y INVX1_LOC_31/A 0.07fF
C42518 INVX1_LOC_182/A NOR2X1_LOC_850/B 0.02fF
C42519 INVX1_LOC_11/A NOR2X1_LOC_703/B 0.03fF
C42520 INVX1_LOC_136/A NAND2X1_LOC_793/Y 0.08fF
C42521 INVX1_LOC_178/A NOR2X1_LOC_716/B 0.10fF
C42522 INVX1_LOC_17/A NOR2X1_LOC_91/Y 0.03fF
C42523 INVX1_LOC_103/A NOR2X1_LOC_457/B 0.08fF
C42524 INVX1_LOC_11/Y INVX1_LOC_297/A 0.03fF
C42525 INVX1_LOC_50/A NAND2X1_LOC_170/A 0.03fF
C42526 INVX1_LOC_294/Y NOR2X1_LOC_652/Y 0.05fF
C42527 NAND2X1_LOC_326/A NOR2X1_LOC_152/Y 0.04fF
C42528 NOR2X1_LOC_211/A NOR2X1_LOC_748/A 0.56fF
C42529 NOR2X1_LOC_15/Y INVX1_LOC_77/A 0.06fF
C42530 INVX1_LOC_46/A INVX1_LOC_307/A 0.07fF
C42531 NOR2X1_LOC_382/Y INVX1_LOC_31/A 0.02fF
C42532 INPUT_0 INVX1_LOC_102/A 0.10fF
C42533 NOR2X1_LOC_791/Y NOR2X1_LOC_309/Y 0.02fF
C42534 INVX1_LOC_64/A INVX1_LOC_143/A 0.09fF
C42535 NOR2X1_LOC_75/Y NOR2X1_LOC_273/a_36_216# 0.00fF
C42536 NOR2X1_LOC_590/A NOR2X1_LOC_274/B 0.02fF
C42537 INVX1_LOC_58/A INVX1_LOC_1/Y 0.03fF
C42538 INVX1_LOC_223/Y INVX1_LOC_104/A 0.02fF
C42539 INVX1_LOC_83/A NOR2X1_LOC_686/A 0.40fF
C42540 INVX1_LOC_313/Y NAND2X1_LOC_454/Y 0.01fF
C42541 NOR2X1_LOC_113/B NOR2X1_LOC_114/Y 0.01fF
C42542 NAND2X1_LOC_9/Y INVX1_LOC_226/Y 2.36fF
C42543 INVX1_LOC_35/A NOR2X1_LOC_244/B 0.01fF
C42544 INVX1_LOC_22/A NOR2X1_LOC_292/a_36_216# 0.00fF
C42545 INVX1_LOC_117/Y INVX1_LOC_117/A 0.25fF
C42546 INVX1_LOC_36/A INVX1_LOC_30/A 0.14fF
C42547 NOR2X1_LOC_612/a_36_216# NOR2X1_LOC_772/B 0.01fF
C42548 INVX1_LOC_132/A NOR2X1_LOC_538/B 0.01fF
C42549 NAND2X1_LOC_567/Y NAND2X1_LOC_799/A 0.00fF
C42550 INVX1_LOC_24/A INVX1_LOC_43/Y 0.03fF
C42551 INVX1_LOC_21/A INVX1_LOC_177/A 0.06fF
C42552 NOR2X1_LOC_730/A INVX1_LOC_53/A 0.01fF
C42553 NOR2X1_LOC_405/A NAND2X1_LOC_63/Y 0.01fF
C42554 NAND2X1_LOC_35/Y INVX1_LOC_165/Y 0.04fF
C42555 NOR2X1_LOC_510/Y INVX1_LOC_214/A 0.00fF
C42556 INVX1_LOC_251/Y INVX1_LOC_27/A 0.01fF
C42557 NAND2X1_LOC_803/B NOR2X1_LOC_577/Y 0.02fF
C42558 NOR2X1_LOC_89/A INVX1_LOC_91/A 1.94fF
C42559 INVX1_LOC_119/A NOR2X1_LOC_92/Y 0.10fF
C42560 NOR2X1_LOC_295/Y INVX1_LOC_269/A 0.00fF
C42561 INVX1_LOC_299/A INVX1_LOC_225/A 0.45fF
C42562 NOR2X1_LOC_716/B NOR2X1_LOC_786/a_36_216# 0.01fF
C42563 INVX1_LOC_17/Y NOR2X1_LOC_71/Y 0.01fF
C42564 INVX1_LOC_14/A NOR2X1_LOC_124/B 0.62fF
C42565 NOR2X1_LOC_321/Y NOR2X1_LOC_111/a_36_216# 0.00fF
C42566 INVX1_LOC_226/Y NAND2X1_LOC_553/A 0.02fF
C42567 NOR2X1_LOC_155/A INVX1_LOC_38/A 0.07fF
C42568 NOR2X1_LOC_68/A INVX1_LOC_72/A 0.07fF
C42569 NOR2X1_LOC_828/Y NOR2X1_LOC_717/B 0.00fF
C42570 INVX1_LOC_124/A NOR2X1_LOC_15/Y 0.17fF
C42571 NOR2X1_LOC_216/B INVX1_LOC_280/A 0.07fF
C42572 NAND2X1_LOC_763/B NAND2X1_LOC_587/a_36_24# 0.00fF
C42573 INVX1_LOC_75/A NOR2X1_LOC_415/Y 0.01fF
C42574 NAND2X1_LOC_588/B INVX1_LOC_18/A 0.02fF
C42575 NOR2X1_LOC_590/A NOR2X1_LOC_577/Y 0.08fF
C42576 NAND2X1_LOC_808/A INVX1_LOC_53/A 0.09fF
C42577 INVX1_LOC_233/A INVX1_LOC_10/A 0.00fF
C42578 NOR2X1_LOC_208/Y INVX1_LOC_30/A 0.32fF
C42579 INVX1_LOC_232/Y INVX1_LOC_163/A 0.01fF
C42580 INVX1_LOC_136/A NOR2X1_LOC_607/A 0.01fF
C42581 NOR2X1_LOC_67/A INVX1_LOC_48/Y 0.01fF
C42582 INVX1_LOC_278/A D_INPUT_0 0.07fF
C42583 NOR2X1_LOC_644/A NOR2X1_LOC_858/A 0.00fF
C42584 NOR2X1_LOC_170/A INVX1_LOC_91/A 0.04fF
C42585 NOR2X1_LOC_68/A INVX1_LOC_198/Y 0.00fF
C42586 NOR2X1_LOC_278/A NAND2X1_LOC_793/Y 0.01fF
C42587 NOR2X1_LOC_648/a_36_216# NAND2X1_LOC_190/Y 0.00fF
C42588 NOR2X1_LOC_237/Y INVX1_LOC_30/A 0.10fF
C42589 INVX1_LOC_64/A NAND2X1_LOC_800/Y 0.04fF
C42590 INVX1_LOC_61/A NAND2X1_LOC_100/a_36_24# 0.09fF
C42591 NOR2X1_LOC_828/Y NOR2X1_LOC_828/A 0.00fF
C42592 INVX1_LOC_163/A INVX1_LOC_197/Y 0.05fF
C42593 INVX1_LOC_64/A NOR2X1_LOC_130/A 0.06fF
C42594 NAND2X1_LOC_848/A INVX1_LOC_84/A 0.02fF
C42595 NOR2X1_LOC_598/B INVX1_LOC_90/A 0.17fF
C42596 NOR2X1_LOC_641/B NAND2X1_LOC_361/Y 0.02fF
C42597 INVX1_LOC_269/A NOR2X1_LOC_399/Y 0.01fF
C42598 NOR2X1_LOC_804/B INVX1_LOC_30/A 0.15fF
C42599 NOR2X1_LOC_717/B INVX1_LOC_5/A 0.03fF
C42600 INVX1_LOC_269/A NOR2X1_LOC_220/A 0.10fF
C42601 INVX1_LOC_12/A INVX1_LOC_46/A 0.76fF
C42602 NAND2X1_LOC_640/a_36_24# INVX1_LOC_71/A 0.00fF
C42603 NAND2X1_LOC_577/A NAND2X1_LOC_139/A 0.03fF
C42604 NOR2X1_LOC_111/A NOR2X1_LOC_831/Y 0.09fF
C42605 NOR2X1_LOC_519/Y INVX1_LOC_46/A 0.02fF
C42606 NAND2X1_LOC_728/Y NAND2X1_LOC_567/Y 0.09fF
C42607 INVX1_LOC_21/A NAND2X1_LOC_573/A 0.07fF
C42608 NAND2X1_LOC_725/A INVX1_LOC_90/A 0.03fF
C42609 INVX1_LOC_34/A INVX1_LOC_223/A 0.07fF
C42610 INVX1_LOC_58/A NOR2X1_LOC_742/A 0.05fF
C42611 NOR2X1_LOC_644/A INVX1_LOC_292/Y 0.01fF
C42612 VDD NOR2X1_LOC_240/B -0.00fF
C42613 NOR2X1_LOC_319/B NOR2X1_LOC_856/B 0.01fF
C42614 INVX1_LOC_135/A INVX1_LOC_93/A 0.10fF
C42615 NOR2X1_LOC_82/A NAND2X1_LOC_181/Y 0.03fF
C42616 NOR2X1_LOC_646/A INVX1_LOC_14/A 0.07fF
C42617 INVX1_LOC_5/A NOR2X1_LOC_130/Y 0.02fF
C42618 NOR2X1_LOC_309/Y INVX1_LOC_30/A 0.21fF
C42619 NOR2X1_LOC_632/Y INVX1_LOC_1/A 0.05fF
C42620 INVX1_LOC_170/A NOR2X1_LOC_315/Y 0.00fF
C42621 NOR2X1_LOC_470/B NOR2X1_LOC_589/A 0.49fF
C42622 INVX1_LOC_230/Y NAND2X1_LOC_549/B 0.03fF
C42623 INVX1_LOC_7/Y INVX1_LOC_89/A 0.00fF
C42624 NAND2X1_LOC_642/Y INVX1_LOC_94/Y 0.12fF
C42625 INVX1_LOC_118/Y INVX1_LOC_19/A 0.03fF
C42626 NOR2X1_LOC_624/A NAND2X1_LOC_364/A -0.03fF
C42627 NOR2X1_LOC_860/B INVX1_LOC_77/A 0.07fF
C42628 INVX1_LOC_269/A NOR2X1_LOC_548/Y 0.21fF
C42629 D_INPUT_1 NOR2X1_LOC_74/A 0.10fF
C42630 INVX1_LOC_101/Y NOR2X1_LOC_665/A 0.02fF
C42631 NOR2X1_LOC_598/B NAND2X1_LOC_348/A 0.07fF
C42632 NAND2X1_LOC_577/A NAND2X1_LOC_139/a_36_24# 0.02fF
C42633 NAND2X1_LOC_643/a_36_24# INVX1_LOC_94/Y 0.00fF
C42634 VDD INVX1_LOC_19/Y 0.44fF
C42635 NOR2X1_LOC_590/A NOR2X1_LOC_346/B 0.03fF
C42636 INVX1_LOC_33/A INVX1_LOC_94/A 0.08fF
C42637 INVX1_LOC_98/A NAND2X1_LOC_99/A 0.01fF
C42638 NAND2X1_LOC_559/Y NOR2X1_LOC_298/Y 0.06fF
C42639 INVX1_LOC_84/A INVX1_LOC_46/Y 0.09fF
C42640 NAND2X1_LOC_803/B INVX1_LOC_22/A 0.01fF
C42641 INVX1_LOC_36/A NAND2X1_LOC_722/A 0.07fF
C42642 NOR2X1_LOC_757/A INVX1_LOC_88/A 0.16fF
C42643 NOR2X1_LOC_78/A NAND2X1_LOC_99/A 0.07fF
C42644 D_INPUT_1 NOR2X1_LOC_9/Y 0.16fF
C42645 NOR2X1_LOC_615/Y INVX1_LOC_22/A 0.01fF
C42646 NOR2X1_LOC_554/B NOR2X1_LOC_87/B 0.09fF
C42647 NAND2X1_LOC_721/A INVX1_LOC_3/Y 0.34fF
C42648 NOR2X1_LOC_388/Y NOR2X1_LOC_303/Y 0.05fF
C42649 NOR2X1_LOC_92/Y INVX1_LOC_89/A 0.07fF
C42650 NAND2X1_LOC_842/B NAND2X1_LOC_474/Y 0.63fF
C42651 INVX1_LOC_5/A NOR2X1_LOC_151/Y 0.07fF
C42652 NOR2X1_LOC_643/A INVX1_LOC_83/A 0.02fF
C42653 NOR2X1_LOC_778/B NOR2X1_LOC_778/Y -0.01fF
C42654 NOR2X1_LOC_859/Y INVX1_LOC_15/A 0.01fF
C42655 NOR2X1_LOC_590/A INVX1_LOC_22/A 0.08fF
C42656 INVX1_LOC_24/Y INVX1_LOC_89/A 0.08fF
C42657 NAND2X1_LOC_796/B NOR2X1_LOC_329/B 0.01fF
C42658 NAND2X1_LOC_642/Y INVX1_LOC_181/A 0.00fF
C42659 NOR2X1_LOC_45/B INVX1_LOC_271/A 0.45fF
C42660 INVX1_LOC_41/A NAND2X1_LOC_850/a_36_24# 0.00fF
C42661 NOR2X1_LOC_68/A NOR2X1_LOC_537/Y 0.03fF
C42662 NAND2X1_LOC_354/B NOR2X1_LOC_577/Y 0.07fF
C42663 INVX1_LOC_108/A INVX1_LOC_29/A 0.00fF
C42664 INVX1_LOC_12/Y NOR2X1_LOC_38/B 0.18fF
C42665 INVX1_LOC_22/Y INVX1_LOC_22/A 0.10fF
C42666 NOR2X1_LOC_68/A NAND2X1_LOC_338/B 0.14fF
C42667 INVX1_LOC_58/A NOR2X1_LOC_318/B 0.10fF
C42668 NOR2X1_LOC_635/A INVX1_LOC_77/A 0.05fF
C42669 INVX1_LOC_279/A NOR2X1_LOC_160/B 0.71fF
C42670 NAND2X1_LOC_798/B NAND2X1_LOC_74/B 0.07fF
C42671 NOR2X1_LOC_68/A NAND2X1_LOC_323/B 0.00fF
C42672 INVX1_LOC_161/Y NAND2X1_LOC_140/A 0.01fF
C42673 INVX1_LOC_58/A INVX1_LOC_93/Y 0.30fF
C42674 INVX1_LOC_35/A NOR2X1_LOC_685/A 0.01fF
C42675 NAND2X1_LOC_464/A NAND2X1_LOC_99/A 0.02fF
C42676 INVX1_LOC_35/A INVX1_LOC_186/A 0.03fF
C42677 INVX1_LOC_77/A INVX1_LOC_96/Y 0.03fF
C42678 NOR2X1_LOC_824/A INVX1_LOC_91/Y 0.01fF
C42679 NOR2X1_LOC_9/Y NOR2X1_LOC_652/Y 0.27fF
C42680 INVX1_LOC_87/A INVX1_LOC_117/A 0.01fF
C42681 INVX1_LOC_225/A INVX1_LOC_162/A 0.03fF
C42682 INVX1_LOC_11/Y NAND2X1_LOC_804/A 0.02fF
C42683 INVX1_LOC_132/A INVX1_LOC_310/A 0.29fF
C42684 INVX1_LOC_34/A INVX1_LOC_85/A 0.03fF
C42685 NAND2X1_LOC_592/a_36_24# INVX1_LOC_18/A 0.00fF
C42686 NAND2X1_LOC_349/B INVX1_LOC_177/Y 0.02fF
C42687 INVX1_LOC_21/A INVX1_LOC_285/Y 0.01fF
C42688 INVX1_LOC_14/A INVX1_LOC_82/Y 0.04fF
C42689 NOR2X1_LOC_389/A NOR2X1_LOC_214/B 0.01fF
C42690 INVX1_LOC_276/Y NOR2X1_LOC_577/Y 0.06fF
C42691 INVX1_LOC_181/Y INVX1_LOC_16/A 0.03fF
C42692 INVX1_LOC_13/A NOR2X1_LOC_360/Y 0.03fF
C42693 INVX1_LOC_292/A NOR2X1_LOC_180/B 0.03fF
C42694 INVX1_LOC_77/A INVX1_LOC_226/A 0.03fF
C42695 NOR2X1_LOC_181/Y NOR2X1_LOC_180/Y 0.29fF
C42696 INVX1_LOC_61/A NOR2X1_LOC_86/A 0.21fF
C42697 INVX1_LOC_90/A NOR2X1_LOC_372/A 0.03fF
C42698 INVX1_LOC_35/A INVX1_LOC_74/Y 0.02fF
C42699 INVX1_LOC_103/A INVX1_LOC_73/A 0.00fF
C42700 INVX1_LOC_201/Y INVX1_LOC_267/A 0.01fF
C42701 INVX1_LOC_58/A INVX1_LOC_139/A 0.01fF
C42702 NOR2X1_LOC_67/A NOR2X1_LOC_412/a_36_216# 0.00fF
C42703 INVX1_LOC_35/A NAND2X1_LOC_447/Y 0.03fF
C42704 INVX1_LOC_18/A NAND2X1_LOC_662/a_36_24# 0.01fF
C42705 NAND2X1_LOC_444/B INVX1_LOC_185/A 0.09fF
C42706 NOR2X1_LOC_136/Y INVX1_LOC_33/A 0.03fF
C42707 NAND2X1_LOC_231/Y INVX1_LOC_162/Y 0.11fF
C42708 INVX1_LOC_24/A NOR2X1_LOC_721/a_36_216# 0.00fF
C42709 NOR2X1_LOC_89/A INVX1_LOC_203/A 0.01fF
C42710 INVX1_LOC_45/A INVX1_LOC_85/Y 0.07fF
C42711 INVX1_LOC_58/A NAND2X1_LOC_721/A 0.44fF
C42712 NOR2X1_LOC_824/A NOR2X1_LOC_45/B 0.07fF
C42713 INVX1_LOC_278/A NOR2X1_LOC_266/B 0.03fF
C42714 INVX1_LOC_292/A INVX1_LOC_73/A 0.06fF
C42715 INVX1_LOC_195/A INVX1_LOC_175/Y 0.02fF
C42716 INVX1_LOC_58/A NOR2X1_LOC_323/a_36_216# 0.00fF
C42717 NOR2X1_LOC_798/A NOR2X1_LOC_799/B 0.00fF
C42718 INVX1_LOC_237/A NOR2X1_LOC_45/B 0.68fF
C42719 INVX1_LOC_77/A NOR2X1_LOC_97/B 0.03fF
C42720 NOR2X1_LOC_67/A NOR2X1_LOC_84/Y 0.17fF
C42721 NOR2X1_LOC_500/A INVX1_LOC_135/A 0.07fF
C42722 NOR2X1_LOC_731/A NOR2X1_LOC_731/Y 0.02fF
C42723 NOR2X1_LOC_68/A INVX1_LOC_313/Y 0.03fF
C42724 NOR2X1_LOC_400/A VDD 0.00fF
C42725 INVX1_LOC_21/A NOR2X1_LOC_137/B 0.02fF
C42726 INVX1_LOC_34/A NAND2X1_LOC_662/Y 0.08fF
C42727 INVX1_LOC_227/A NOR2X1_LOC_577/Y 0.01fF
C42728 INVX1_LOC_292/A NOR2X1_LOC_569/A 0.03fF
C42729 NAND2X1_LOC_338/B NAND2X1_LOC_464/a_36_24# 0.00fF
C42730 NOR2X1_LOC_214/B NOR2X1_LOC_596/A 0.06fF
C42731 INVX1_LOC_50/Y INVX1_LOC_76/A 0.17fF
C42732 INVX1_LOC_279/A NOR2X1_LOC_544/a_36_216# 0.00fF
C42733 INVX1_LOC_89/A NAND2X1_LOC_837/Y 0.05fF
C42734 NAND2X1_LOC_349/B INVX1_LOC_104/A 0.05fF
C42735 NOR2X1_LOC_773/Y INVX1_LOC_98/Y 0.02fF
C42736 NOR2X1_LOC_667/A INVX1_LOC_280/Y 0.03fF
C42737 NAND2X1_LOC_733/B NAND2X1_LOC_723/a_36_24# 0.02fF
C42738 NOR2X1_LOC_598/B INVX1_LOC_38/A 0.21fF
C42739 INVX1_LOC_278/A NAND2X1_LOC_848/A 0.10fF
C42740 INVX1_LOC_11/A INVX1_LOC_91/A 0.55fF
C42741 NOR2X1_LOC_626/Y VDD 0.18fF
C42742 NAND2X1_LOC_149/Y INVX1_LOC_115/A 0.04fF
C42743 INVX1_LOC_8/Y INVX1_LOC_47/A 0.01fF
C42744 NOR2X1_LOC_92/Y NOR2X1_LOC_24/Y 0.02fF
C42745 NAND2X1_LOC_569/B NOR2X1_LOC_536/A 0.30fF
C42746 INVX1_LOC_223/A INPUT_0 0.03fF
C42747 INVX1_LOC_177/Y INVX1_LOC_75/A 0.68fF
C42748 INVX1_LOC_97/Y INVX1_LOC_38/A 0.05fF
C42749 INVX1_LOC_258/Y VDD 0.21fF
C42750 INVX1_LOC_7/A NOR2X1_LOC_6/B 0.08fF
C42751 NAND2X1_LOC_725/A INVX1_LOC_38/A 0.03fF
C42752 INVX1_LOC_50/A INVX1_LOC_179/A 0.03fF
C42753 INVX1_LOC_138/Y INVX1_LOC_230/A 0.01fF
C42754 INVX1_LOC_1/A NAND2X1_LOC_1/Y 0.02fF
C42755 INVX1_LOC_41/A INVX1_LOC_89/A 0.18fF
C42756 NAND2X1_LOC_231/Y NAND2X1_LOC_662/Y 0.03fF
C42757 INVX1_LOC_58/A INVX1_LOC_117/Y 0.08fF
C42758 INVX1_LOC_5/A NAND2X1_LOC_423/a_36_24# 0.00fF
C42759 NAND2X1_LOC_715/B INVX1_LOC_38/A 0.06fF
C42760 NOR2X1_LOC_612/Y NOR2X1_LOC_717/A 0.02fF
C42761 INVX1_LOC_201/Y INVX1_LOC_89/A 0.83fF
C42762 INVX1_LOC_274/A NOR2X1_LOC_678/A 0.00fF
C42763 NOR2X1_LOC_536/A NOR2X1_LOC_81/Y 0.01fF
C42764 NOR2X1_LOC_65/B NAND2X1_LOC_572/B 0.03fF
C42765 INVX1_LOC_49/A INVX1_LOC_311/Y 0.03fF
C42766 INVX1_LOC_177/A NOR2X1_LOC_565/B 0.01fF
C42767 NOR2X1_LOC_246/A NOR2X1_LOC_792/B 0.02fF
C42768 INVX1_LOC_24/A INVX1_LOC_282/A 0.15fF
C42769 INVX1_LOC_1/A NAND2X1_LOC_39/Y 0.02fF
C42770 NOR2X1_LOC_99/a_36_216# INVX1_LOC_306/Y 0.00fF
C42771 INVX1_LOC_53/A INVX1_LOC_92/A 0.20fF
C42772 INVX1_LOC_27/A INVX1_LOC_281/A 0.01fF
C42773 INVX1_LOC_14/A INVX1_LOC_2/Y 0.03fF
C42774 NAND2X1_LOC_714/B INVX1_LOC_33/Y 0.00fF
C42775 NAND2X1_LOC_564/B NAND2X1_LOC_862/A 0.23fF
C42776 NAND2X1_LOC_11/Y INPUT_5 1.01fF
C42777 INVX1_LOC_232/A NOR2X1_LOC_121/A 0.31fF
C42778 NOR2X1_LOC_82/Y INVX1_LOC_22/A 0.08fF
C42779 NOR2X1_LOC_15/Y INVX1_LOC_194/Y 0.01fF
C42780 NAND2X1_LOC_195/a_36_24# NAND2X1_LOC_662/Y 0.02fF
C42781 NAND2X1_LOC_725/A NOR2X1_LOC_51/A 0.04fF
C42782 NOR2X1_LOC_843/B NOR2X1_LOC_814/A 0.13fF
C42783 NOR2X1_LOC_716/B INVX1_LOC_140/A 0.37fF
C42784 NOR2X1_LOC_468/Y INVX1_LOC_12/Y 0.10fF
C42785 NOR2X1_LOC_355/A NAND2X1_LOC_675/a_36_24# 0.00fF
C42786 NOR2X1_LOC_433/A INVX1_LOC_79/A 0.07fF
C42787 NOR2X1_LOC_25/Y NOR2X1_LOC_36/B 0.24fF
C42788 INVX1_LOC_113/Y NOR2X1_LOC_74/a_36_216# 0.00fF
C42789 INVX1_LOC_279/A INVX1_LOC_208/A 0.10fF
C42790 INVX1_LOC_89/A INVX1_LOC_64/Y 0.07fF
C42791 NAND2X1_LOC_552/A INVX1_LOC_71/Y 0.19fF
C42792 NOR2X1_LOC_130/A NAND2X1_LOC_850/Y 0.07fF
C42793 D_GATE_366 INVX1_LOC_266/Y 0.07fF
C42794 INVX1_LOC_64/A NOR2X1_LOC_197/B 0.01fF
C42795 NOR2X1_LOC_394/Y INVX1_LOC_42/A 0.00fF
C42796 INVX1_LOC_279/A NOR2X1_LOC_516/B 0.07fF
C42797 NAND2X1_LOC_361/Y NOR2X1_LOC_751/A 0.01fF
C42798 NAND2X1_LOC_363/a_36_24# NAND2X1_LOC_363/Y 0.02fF
C42799 NOR2X1_LOC_596/A NOR2X1_LOC_741/A 0.01fF
C42800 INVX1_LOC_174/A VDD 0.22fF
C42801 INVX1_LOC_33/A INVX1_LOC_144/A 0.01fF
C42802 NAND2X1_LOC_93/B NOR2X1_LOC_81/Y 0.02fF
C42803 NOR2X1_LOC_590/Y INVX1_LOC_179/A 0.01fF
C42804 D_GATE_222 INVX1_LOC_83/A -0.01fF
C42805 INVX1_LOC_286/Y INVX1_LOC_20/A 0.15fF
C42806 NAND2X1_LOC_708/Y NOR2X1_LOC_697/Y 0.06fF
C42807 NOR2X1_LOC_48/Y INVX1_LOC_296/A 0.18fF
C42808 NAND2X1_LOC_538/Y NOR2X1_LOC_536/A 0.03fF
C42809 INVX1_LOC_171/A NOR2X1_LOC_568/a_36_216# 0.00fF
C42810 NOR2X1_LOC_82/A INVX1_LOC_117/A 0.05fF
C42811 NAND2X1_LOC_581/Y NAND2X1_LOC_51/B 0.02fF
C42812 NOR2X1_LOC_15/Y INVX1_LOC_9/A 0.09fF
C42813 NAND2X1_LOC_656/A NOR2X1_LOC_78/A 0.02fF
C42814 INVX1_LOC_75/A INVX1_LOC_104/A 0.33fF
C42815 INVX1_LOC_1/A NOR2X1_LOC_186/a_36_216# 0.00fF
C42816 NAND2X1_LOC_733/Y INVX1_LOC_46/A 0.03fF
C42817 INVX1_LOC_311/A INVX1_LOC_153/Y 0.10fF
C42818 NOR2X1_LOC_655/Y NOR2X1_LOC_611/a_36_216# 0.00fF
C42819 INVX1_LOC_183/A INVX1_LOC_102/A 0.03fF
C42820 NAND2X1_LOC_270/a_36_24# INVX1_LOC_8/A 0.00fF
C42821 NOR2X1_LOC_250/A NOR2X1_LOC_536/A 0.01fF
C42822 NOR2X1_LOC_52/B INVX1_LOC_79/A 0.07fF
C42823 NAND2X1_LOC_336/a_36_24# INVX1_LOC_33/Y 0.00fF
C42824 INVX1_LOC_89/A NOR2X1_LOC_211/A 0.01fF
C42825 INVX1_LOC_162/Y INPUT_0 0.19fF
C42826 INVX1_LOC_217/A NOR2X1_LOC_164/Y 0.08fF
C42827 NOR2X1_LOC_798/A NOR2X1_LOC_445/B 0.02fF
C42828 NAND2X1_LOC_363/B INVX1_LOC_63/A 0.07fF
C42829 INVX1_LOC_144/A NAND2X1_LOC_466/A 0.03fF
C42830 INVX1_LOC_27/A NOR2X1_LOC_862/B 0.21fF
C42831 NOR2X1_LOC_500/A NOR2X1_LOC_552/A 0.22fF
C42832 NOR2X1_LOC_433/A INVX1_LOC_91/A 0.22fF
C42833 NAND2X1_LOC_326/A INVX1_LOC_291/A 0.02fF
C42834 NOR2X1_LOC_530/Y NOR2X1_LOC_536/A 0.01fF
C42835 NOR2X1_LOC_552/A NOR2X1_LOC_303/Y 0.10fF
C42836 INVX1_LOC_311/A INVX1_LOC_121/Y 0.00fF
C42837 NAND2X1_LOC_198/B NAND2X1_LOC_468/B 0.05fF
C42838 NOR2X1_LOC_500/B INVX1_LOC_37/A 0.01fF
C42839 INVX1_LOC_161/Y INVX1_LOC_118/Y 0.07fF
C42840 NOR2X1_LOC_593/Y INVX1_LOC_91/A 0.06fF
C42841 NOR2X1_LOC_654/A INVX1_LOC_42/A 0.01fF
C42842 INVX1_LOC_2/A NOR2X1_LOC_335/B 0.06fF
C42843 INVX1_LOC_217/A INVX1_LOC_46/A 1.82fF
C42844 NOR2X1_LOC_218/A INVX1_LOC_54/A 0.03fF
C42845 INVX1_LOC_89/A INVX1_LOC_121/A 0.01fF
C42846 INVX1_LOC_208/A INVX1_LOC_182/Y 0.22fF
C42847 NAND2X1_LOC_364/A INVX1_LOC_14/Y 0.08fF
C42848 NAND2X1_LOC_9/Y INVX1_LOC_12/A 0.03fF
C42849 NOR2X1_LOC_52/B NOR2X1_LOC_114/A 0.05fF
C42850 INVX1_LOC_58/A NAND2X1_LOC_636/a_36_24# 0.00fF
C42851 NOR2X1_LOC_791/Y INVX1_LOC_63/A 0.05fF
C42852 INVX1_LOC_142/A NAND2X1_LOC_472/Y 0.00fF
C42853 NAND2X1_LOC_112/Y NOR2X1_LOC_329/B 0.02fF
C42854 INVX1_LOC_233/A INVX1_LOC_12/A 0.39fF
C42855 INVX1_LOC_77/A NOR2X1_LOC_137/a_36_216# 0.00fF
C42856 NAND2X1_LOC_165/a_36_24# NOR2X1_LOC_337/A 0.00fF
C42857 NAND2X1_LOC_842/B INVX1_LOC_10/A 0.19fF
C42858 NAND2X1_LOC_303/B NAND2X1_LOC_302/a_36_24# 0.02fF
C42859 NOR2X1_LOC_52/B INVX1_LOC_91/A 0.18fF
C42860 NOR2X1_LOC_140/A NOR2X1_LOC_649/B 0.07fF
C42861 INVX1_LOC_3/A NAND2X1_LOC_218/A 0.05fF
C42862 NOR2X1_LOC_140/A INVX1_LOC_3/A 0.08fF
C42863 INVX1_LOC_240/A NAND2X1_LOC_729/B 0.52fF
C42864 NOR2X1_LOC_553/Y NOR2X1_LOC_74/A 0.00fF
C42865 NOR2X1_LOC_303/Y INVX1_LOC_139/Y 0.09fF
C42866 NAND2X1_LOC_553/A INVX1_LOC_12/A 0.03fF
C42867 NOR2X1_LOC_639/B NOR2X1_LOC_48/B 0.03fF
C42868 NOR2X1_LOC_315/Y NAND2X1_LOC_642/Y 0.01fF
C42869 INVX1_LOC_303/A INVX1_LOC_37/A 0.26fF
C42870 NAND2X1_LOC_787/B INVX1_LOC_46/A 0.07fF
C42871 INVX1_LOC_21/A NAND2X1_LOC_81/B 4.02fF
C42872 NOR2X1_LOC_91/A NOR2X1_LOC_278/Y 0.03fF
C42873 INVX1_LOC_153/A VDD -0.00fF
C42874 NOR2X1_LOC_798/A INVX1_LOC_12/A 0.02fF
C42875 INVX1_LOC_54/Y NOR2X1_LOC_552/A 0.04fF
C42876 INVX1_LOC_78/A NOR2X1_LOC_654/A 0.03fF
C42877 INVX1_LOC_304/Y NOR2X1_LOC_164/Y 0.03fF
C42878 INVX1_LOC_249/A INVX1_LOC_281/A 0.17fF
C42879 INVX1_LOC_30/A NOR2X1_LOC_435/A 0.03fF
C42880 NOR2X1_LOC_6/B INVX1_LOC_76/A 0.12fF
C42881 INVX1_LOC_58/A INVX1_LOC_87/A 0.03fF
C42882 NAND2X1_LOC_391/Y NAND2X1_LOC_254/Y 0.03fF
C42883 INVX1_LOC_53/A NAND2X1_LOC_247/a_36_24# 0.00fF
C42884 NOR2X1_LOC_598/B NAND2X1_LOC_223/A 0.07fF
C42885 INVX1_LOC_50/A NOR2X1_LOC_693/Y 0.02fF
C42886 NOR2X1_LOC_860/B INVX1_LOC_9/A 0.47fF
C42887 INVX1_LOC_304/Y INVX1_LOC_46/A 0.07fF
C42888 INVX1_LOC_136/A NAND2X1_LOC_798/B 0.10fF
C42889 INVX1_LOC_78/A INVX1_LOC_58/Y 0.07fF
C42890 NOR2X1_LOC_695/Y NOR2X1_LOC_45/B 0.01fF
C42891 INVX1_LOC_242/Y INVX1_LOC_240/Y 0.10fF
C42892 NOR2X1_LOC_598/B INVX1_LOC_18/Y 0.02fF
C42893 NOR2X1_LOC_736/Y NOR2X1_LOC_736/a_36_216# 0.02fF
C42894 INVX1_LOC_259/A VDD -0.00fF
C42895 D_INPUT_0 INVX1_LOC_123/A 0.07fF
C42896 NOR2X1_LOC_329/B NAND2X1_LOC_840/Y 0.01fF
C42897 NOR2X1_LOC_590/A INVX1_LOC_186/Y 0.07fF
C42898 INVX1_LOC_72/Y INVX1_LOC_123/Y 0.01fF
C42899 INVX1_LOC_234/A NOR2X1_LOC_45/B 0.25fF
C42900 INVX1_LOC_135/Y NAND2X1_LOC_463/B 0.15fF
C42901 NAND2X1_LOC_156/B NOR2X1_LOC_45/B 0.09fF
C42902 INVX1_LOC_18/A INVX1_LOC_285/A 0.15fF
C42903 INVX1_LOC_30/A INVX1_LOC_63/A 0.18fF
C42904 INVX1_LOC_21/A INVX1_LOC_4/Y 0.35fF
C42905 NAND2X1_LOC_308/Y NAND2X1_LOC_264/a_36_24# 0.00fF
C42906 INVX1_LOC_13/Y NAND2X1_LOC_72/B 0.01fF
C42907 INVX1_LOC_45/A NAND2X1_LOC_782/B 0.01fF
C42908 NOR2X1_LOC_709/A NOR2X1_LOC_536/A 0.13fF
C42909 NAND2X1_LOC_629/Y NOR2X1_LOC_684/Y 0.02fF
C42910 NOR2X1_LOC_315/Y NOR2X1_LOC_271/Y 0.02fF
C42911 VDD NOR2X1_LOC_131/Y 0.01fF
C42912 INVX1_LOC_304/A NAND2X1_LOC_573/A 0.02fF
C42913 NOR2X1_LOC_418/Y VDD 0.09fF
C42914 INVX1_LOC_18/A NOR2X1_LOC_814/A 0.08fF
C42915 NAND2X1_LOC_751/a_36_24# NAND2X1_LOC_215/A 0.01fF
C42916 NOR2X1_LOC_178/Y NOR2X1_LOC_72/Y 0.02fF
C42917 NAND2X1_LOC_660/A INVX1_LOC_38/A 0.19fF
C42918 NOR2X1_LOC_731/Y INVX1_LOC_117/A 0.01fF
C42919 INVX1_LOC_33/A NOR2X1_LOC_155/A 0.17fF
C42920 NOR2X1_LOC_554/B NAND2X1_LOC_219/B 0.01fF
C42921 NOR2X1_LOC_773/Y NOR2X1_LOC_322/a_36_216# 0.01fF
C42922 NOR2X1_LOC_82/A INVX1_LOC_3/Y 1.62fF
C42923 INVX1_LOC_11/A NAND2X1_LOC_429/a_36_24# 0.00fF
C42924 NOR2X1_LOC_172/Y NOR2X1_LOC_58/Y 0.01fF
C42925 NOR2X1_LOC_433/A NAND2X1_LOC_273/a_36_24# 0.01fF
C42926 NOR2X1_LOC_743/a_36_216# NOR2X1_LOC_155/A 0.00fF
C42927 NOR2X1_LOC_589/A VDD 0.63fF
C42928 NAND2X1_LOC_30/Y INVX1_LOC_15/A 0.34fF
C42929 INVX1_LOC_279/A NAND2X1_LOC_211/Y 0.07fF
C42930 NAND2X1_LOC_377/Y VDD 0.02fF
C42931 NOR2X1_LOC_329/B NOR2X1_LOC_78/A 0.03fF
C42932 NOR2X1_LOC_822/Y INVX1_LOC_54/A 0.09fF
C42933 INVX1_LOC_229/Y VDD 2.19fF
C42934 INVX1_LOC_75/A INVX1_LOC_86/Y 0.06fF
C42935 INVX1_LOC_49/A INVX1_LOC_84/A 0.20fF
C42936 INVX1_LOC_311/A INVX1_LOC_285/Y 0.08fF
C42937 NOR2X1_LOC_214/B NAND2X1_LOC_469/B 0.01fF
C42938 NOR2X1_LOC_773/Y NOR2X1_LOC_709/B 0.01fF
C42939 NOR2X1_LOC_709/A NAND2X1_LOC_93/B 0.08fF
C42940 NOR2X1_LOC_134/Y INVX1_LOC_15/A 0.03fF
C42941 NOR2X1_LOC_451/A NAND2X1_LOC_451/Y 0.07fF
C42942 NOR2X1_LOC_63/a_36_216# INVX1_LOC_46/Y 0.00fF
C42943 NOR2X1_LOC_160/B NOR2X1_LOC_38/B 0.03fF
C42944 INVX1_LOC_171/A VDD 0.26fF
C42945 NOR2X1_LOC_75/Y INVX1_LOC_78/A 0.06fF
C42946 NOR2X1_LOC_78/B INVX1_LOC_92/A 0.05fF
C42947 INVX1_LOC_306/A INVX1_LOC_117/A 0.03fF
C42948 INVX1_LOC_2/A NOR2X1_LOC_88/Y 0.20fF
C42949 INVX1_LOC_178/A NOR2X1_LOC_591/A 0.01fF
C42950 INVX1_LOC_44/Y NOR2X1_LOC_197/B 0.02fF
C42951 INVX1_LOC_254/Y NAND2X1_LOC_63/Y 0.05fF
C42952 NOR2X1_LOC_226/A NOR2X1_LOC_88/Y 0.14fF
C42953 NOR2X1_LOC_97/B INVX1_LOC_9/A 0.05fF
C42954 INVX1_LOC_136/A INVX1_LOC_47/Y 0.03fF
C42955 INVX1_LOC_244/A INVX1_LOC_37/A 0.12fF
C42956 NOR2X1_LOC_709/A INVX1_LOC_3/A 0.11fF
C42957 NAND2X1_LOC_837/Y NOR2X1_LOC_490/a_36_216# 0.01fF
C42958 NOR2X1_LOC_360/Y INVX1_LOC_32/A 13.92fF
C42959 NOR2X1_LOC_772/Y INVX1_LOC_29/A 0.05fF
C42960 INVX1_LOC_14/A INVX1_LOC_29/Y 4.87fF
C42961 INVX1_LOC_2/A INVX1_LOC_84/A 0.36fF
C42962 NAND2X1_LOC_633/Y INVX1_LOC_140/A 0.62fF
C42963 NOR2X1_LOC_860/B NOR2X1_LOC_861/Y 1.72fF
C42964 NOR2X1_LOC_92/Y NOR2X1_LOC_392/Y 0.00fF
C42965 INVX1_LOC_73/A NOR2X1_LOC_137/Y 0.03fF
C42966 NOR2X1_LOC_500/B NAND2X1_LOC_72/B 0.04fF
C42967 NOR2X1_LOC_45/B NOR2X1_LOC_528/Y 0.27fF
C42968 NOR2X1_LOC_226/A INVX1_LOC_84/A 1.32fF
C42969 NAND2X1_LOC_276/Y NOR2X1_LOC_89/A 0.45fF
C42970 NOR2X1_LOC_392/B INVX1_LOC_29/A 0.03fF
C42971 NOR2X1_LOC_716/B INVX1_LOC_42/A 0.14fF
C42972 NAND2X1_LOC_128/a_36_24# NOR2X1_LOC_331/B 0.01fF
C42973 NOR2X1_LOC_590/A NOR2X1_LOC_843/B 0.03fF
C42974 INVX1_LOC_58/A NOR2X1_LOC_82/A 0.09fF
C42975 NAND2X1_LOC_338/B NAND2X1_LOC_768/Y 0.12fF
C42976 INVX1_LOC_22/Y NOR2X1_LOC_843/B 0.00fF
C42977 NAND2X1_LOC_683/a_36_24# INVX1_LOC_291/A 0.01fF
C42978 INVX1_LOC_75/A NAND2X1_LOC_8/a_36_24# 0.00fF
C42979 NOR2X1_LOC_647/A INVX1_LOC_40/Y 0.01fF
C42980 NAND2X1_LOC_53/Y NOR2X1_LOC_604/Y 0.02fF
C42981 INVX1_LOC_34/A INVX1_LOC_290/Y 0.11fF
C42982 NOR2X1_LOC_112/Y INVX1_LOC_280/A 0.03fF
C42983 NOR2X1_LOC_567/B NOR2X1_LOC_319/B 0.13fF
C42984 INVX1_LOC_170/A NAND2X1_LOC_99/A 0.01fF
C42985 INVX1_LOC_222/A VDD 0.12fF
C42986 INVX1_LOC_135/A NOR2X1_LOC_78/Y 0.30fF
C42987 INVX1_LOC_287/A NAND2X1_LOC_701/a_36_24# 0.00fF
C42988 NOR2X1_LOC_456/Y NOR2X1_LOC_446/A 0.02fF
C42989 INVX1_LOC_49/A INVX1_LOC_15/A 17.35fF
C42990 INVX1_LOC_83/A INVX1_LOC_92/A 0.17fF
C42991 INVX1_LOC_216/Y NOR2X1_LOC_660/Y 0.04fF
C42992 INVX1_LOC_233/A INVX1_LOC_200/A 0.18fF
C42993 INVX1_LOC_30/A NOR2X1_LOC_65/Y 0.04fF
C42994 NOR2X1_LOC_170/a_36_216# NAND2X1_LOC_72/B 0.00fF
C42995 INVX1_LOC_1/Y NAND2X1_LOC_475/Y 0.10fF
C42996 NAND2X1_LOC_560/A INVX1_LOC_38/A 0.03fF
C42997 NAND2X1_LOC_162/B INVX1_LOC_78/A 0.01fF
C42998 INVX1_LOC_71/A NAND2X1_LOC_454/Y 0.07fF
C42999 INVX1_LOC_96/A INVX1_LOC_76/A 0.01fF
C43000 D_INPUT_1 INVX1_LOC_124/Y 0.03fF
C43001 INVX1_LOC_230/Y NAND2X1_LOC_549/Y 0.01fF
C43002 INVX1_LOC_278/A NOR2X1_LOC_134/Y 0.02fF
C43003 NAND2X1_LOC_374/Y NOR2X1_LOC_89/A 0.05fF
C43004 NOR2X1_LOC_419/Y INVX1_LOC_78/A 0.02fF
C43005 NOR2X1_LOC_91/Y INVX1_LOC_181/A 0.01fF
C43006 INVX1_LOC_6/A INVX1_LOC_202/Y 0.01fF
C43007 NOR2X1_LOC_346/B NOR2X1_LOC_67/Y 0.07fF
C43008 NOR2X1_LOC_748/Y INVX1_LOC_19/A 0.05fF
C43009 NOR2X1_LOC_275/A NAND2X1_LOC_469/B 0.01fF
C43010 NOR2X1_LOC_716/B INVX1_LOC_78/A 0.15fF
C43011 INVX1_LOC_89/A NAND2X1_LOC_574/A 0.01fF
C43012 NOR2X1_LOC_270/Y INVX1_LOC_271/A 0.01fF
C43013 INVX1_LOC_24/A NOR2X1_LOC_720/A 0.00fF
C43014 NOR2X1_LOC_124/A INVX1_LOC_76/A 0.01fF
C43015 INVX1_LOC_140/A INVX1_LOC_71/Y 0.03fF
C43016 NOR2X1_LOC_589/A INVX1_LOC_133/A 1.72fF
C43017 INVX1_LOC_64/A INVX1_LOC_286/Y 0.15fF
C43018 NOR2X1_LOC_245/a_36_216# NOR2X1_LOC_653/Y 0.00fF
C43019 NAND2X1_LOC_390/a_36_24# NAND2X1_LOC_74/B 0.01fF
C43020 NOR2X1_LOC_848/Y NAND2X1_LOC_473/A 0.04fF
C43021 NOR2X1_LOC_405/A INVX1_LOC_14/Y 0.54fF
C43022 NOR2X1_LOC_420/Y NOR2X1_LOC_160/B 0.01fF
C43023 INVX1_LOC_2/A INVX1_LOC_15/A 0.59fF
C43024 NAND2X1_LOC_348/A INVX1_LOC_152/A 0.25fF
C43025 NOR2X1_LOC_238/Y INVX1_LOC_57/A 0.10fF
C43026 NAND2X1_LOC_648/A INVX1_LOC_84/A 0.00fF
C43027 NOR2X1_LOC_68/A NAND2X1_LOC_415/a_36_24# 0.00fF
C43028 VDD INVX1_LOC_147/Y 0.25fF
C43029 INPUT_1 INVX1_LOC_84/A 11.14fF
C43030 INVX1_LOC_290/A NOR2X1_LOC_584/Y 0.01fF
C43031 NOR2X1_LOC_226/A INVX1_LOC_15/A 0.38fF
C43032 NOR2X1_LOC_152/Y NOR2X1_LOC_654/A 0.10fF
C43033 NOR2X1_LOC_65/B NOR2X1_LOC_716/B 0.10fF
C43034 INVX1_LOC_91/A NOR2X1_LOC_376/Y 0.01fF
C43035 NAND2X1_LOC_96/A NAND2X1_LOC_642/Y 0.01fF
C43036 NOR2X1_LOC_189/A NAND2X1_LOC_787/Y 0.01fF
C43037 VDD INVX1_LOC_20/A 1.64fF
C43038 NOR2X1_LOC_391/B NOR2X1_LOC_78/Y 0.11fF
C43039 INVX1_LOC_219/A NAND2X1_LOC_74/B 0.01fF
C43040 INVX1_LOC_64/A INVX1_LOC_159/A 0.04fF
C43041 NAND2X1_LOC_800/A INVX1_LOC_20/A 0.01fF
C43042 VDD NOR2X1_LOC_360/A 0.24fF
C43043 NAND2X1_LOC_837/Y NOR2X1_LOC_392/Y 0.01fF
C43044 INVX1_LOC_160/A NOR2X1_LOC_729/A 0.01fF
C43045 NOR2X1_LOC_92/Y NOR2X1_LOC_599/Y 0.14fF
C43046 NOR2X1_LOC_468/Y NOR2X1_LOC_160/B 0.35fF
C43047 INVX1_LOC_97/A INVX1_LOC_29/A 0.04fF
C43048 NOR2X1_LOC_261/Y INVX1_LOC_49/A 0.19fF
C43049 NOR2X1_LOC_557/Y INVX1_LOC_129/A -0.02fF
C43050 NOR2X1_LOC_355/a_36_216# INVX1_LOC_29/A 0.00fF
C43051 NOR2X1_LOC_516/B NOR2X1_LOC_38/B 0.06fF
C43052 INVX1_LOC_90/A INVX1_LOC_29/A 2.75fF
C43053 GATE_662 D_INPUT_5 0.03fF
C43054 INVX1_LOC_123/A INVX1_LOC_46/Y 0.15fF
C43055 INVX1_LOC_17/A NAND2X1_LOC_114/B 0.07fF
C43056 INVX1_LOC_72/A NAND2X1_LOC_474/Y 0.00fF
C43057 NOR2X1_LOC_598/B INVX1_LOC_33/A 4.81fF
C43058 NOR2X1_LOC_389/B INVX1_LOC_29/A 0.04fF
C43059 NOR2X1_LOC_236/a_36_216# INVX1_LOC_3/Y 0.00fF
C43060 VDD NOR2X1_LOC_765/Y 0.39fF
C43061 NOR2X1_LOC_802/A NOR2X1_LOC_383/B 0.07fF
C43062 NAND2X1_LOC_303/Y NOR2X1_LOC_761/Y 0.05fF
C43063 NAND2X1_LOC_462/B INVX1_LOC_15/A 0.00fF
C43064 INVX1_LOC_191/Y NOR2X1_LOC_638/Y 0.01fF
C43065 NOR2X1_LOC_223/B INVX1_LOC_49/A 0.06fF
C43066 INVX1_LOC_17/A INVX1_LOC_141/Y 0.05fF
C43067 INVX1_LOC_35/A NAND2X1_LOC_139/A 0.01fF
C43068 NAND2X1_LOC_451/Y INVX1_LOC_262/A 0.03fF
C43069 NOR2X1_LOC_612/B INVX1_LOC_29/Y 0.30fF
C43070 NOR2X1_LOC_272/Y NOR2X1_LOC_106/Y 0.27fF
C43071 NAND2X1_LOC_715/B INVX1_LOC_33/A 0.72fF
C43072 INVX1_LOC_17/A INVX1_LOC_312/Y 0.70fF
C43073 INVX1_LOC_196/A INVX1_LOC_57/A 0.03fF
C43074 INVX1_LOC_17/A NOR2X1_LOC_294/Y 0.98fF
C43075 NAND2X1_LOC_348/A INVX1_LOC_29/A 0.07fF
C43076 NOR2X1_LOC_160/B NOR2X1_LOC_249/a_36_216# 0.00fF
C43077 INVX1_LOC_28/A NOR2X1_LOC_114/Y 0.01fF
C43078 NOR2X1_LOC_470/A INVX1_LOC_78/A 0.15fF
C43079 NOR2X1_LOC_486/Y NOR2X1_LOC_155/A 0.03fF
C43080 NOR2X1_LOC_503/A INVX1_LOC_42/A 0.01fF
C43081 INVX1_LOC_143/A INVX1_LOC_129/A 0.01fF
C43082 NOR2X1_LOC_261/Y INVX1_LOC_2/A 0.18fF
C43083 NOR2X1_LOC_91/A NAND2X1_LOC_392/A 0.01fF
C43084 INVX1_LOC_304/Y INVX1_LOC_233/A 0.01fF
C43085 INPUT_1 INVX1_LOC_15/A 0.03fF
C43086 INVX1_LOC_232/Y INVX1_LOC_23/A 0.07fF
C43087 NOR2X1_LOC_67/A INVX1_LOC_25/A 0.15fF
C43088 NOR2X1_LOC_424/Y INVX1_LOC_78/A 0.09fF
C43089 INVX1_LOC_13/A INVX1_LOC_26/A 0.03fF
C43090 NAND2X1_LOC_53/Y INVX1_LOC_72/A 0.21fF
C43091 INVX1_LOC_236/Y INVX1_LOC_31/A 0.05fF
C43092 NOR2X1_LOC_748/Y INVX1_LOC_26/Y 0.01fF
C43093 NOR2X1_LOC_646/a_36_216# NOR2X1_LOC_647/A 0.02fF
C43094 NOR2X1_LOC_318/B NAND2X1_LOC_475/Y 0.10fF
C43095 INVX1_LOC_88/A NAND2X1_LOC_198/B 0.05fF
C43096 INVX1_LOC_223/A INVX1_LOC_225/Y 0.03fF
C43097 NOR2X1_LOC_634/B INVX1_LOC_53/A 0.02fF
C43098 INVX1_LOC_2/A INVX1_LOC_278/A 0.07fF
C43099 NOR2X1_LOC_717/B INVX1_LOC_78/A 0.03fF
C43100 NOR2X1_LOC_689/Y NAND2X1_LOC_726/Y 0.07fF
C43101 NOR2X1_LOC_151/Y INVX1_LOC_42/A 0.00fF
C43102 NOR2X1_LOC_45/B NAND2X1_LOC_477/Y 0.10fF
C43103 NOR2X1_LOC_78/B INVX1_LOC_53/A 0.31fF
C43104 NAND2X1_LOC_803/B INVX1_LOC_18/A 0.02fF
C43105 NAND2X1_LOC_736/Y GATE_741 0.03fF
C43106 INVX1_LOC_46/A INVX1_LOC_92/A 0.07fF
C43107 NAND2X1_LOC_35/B INVX1_LOC_64/A 0.36fF
C43108 INVX1_LOC_278/A NOR2X1_LOC_226/A 1.09fF
C43109 NAND2X1_LOC_53/Y INVX1_LOC_198/Y 0.24fF
C43110 NOR2X1_LOC_78/A NOR2X1_LOC_691/B 0.01fF
C43111 INVX1_LOC_201/Y INVX1_LOC_235/A 0.05fF
C43112 INPUT_0 INVX1_LOC_290/Y 0.03fF
C43113 NOR2X1_LOC_598/B INVX1_LOC_40/A 0.22fF
C43114 NOR2X1_LOC_454/Y INVX1_LOC_34/A 0.02fF
C43115 NOR2X1_LOC_536/A NOR2X1_LOC_489/A 0.25fF
C43116 INPUT_3 NOR2X1_LOC_360/Y 0.03fF
C43117 NOR2X1_LOC_590/A INVX1_LOC_18/A 0.11fF
C43118 INVX1_LOC_313/A NOR2X1_LOC_278/Y 0.19fF
C43119 NOR2X1_LOC_567/B NOR2X1_LOC_623/B 0.02fF
C43120 NOR2X1_LOC_746/Y INVX1_LOC_19/A 0.01fF
C43121 NAND2X1_LOC_199/B NAND2X1_LOC_195/Y 0.02fF
C43122 INVX1_LOC_201/Y NAND2X1_LOC_393/a_36_24# 0.03fF
C43123 NOR2X1_LOC_431/Y NAND2X1_LOC_350/A 0.03fF
C43124 NOR2X1_LOC_160/B NOR2X1_LOC_596/A 0.03fF
C43125 INVX1_LOC_65/Y INVX1_LOC_26/Y 0.03fF
C43126 NAND2X1_LOC_363/B INVX1_LOC_1/Y 0.01fF
C43127 NOR2X1_LOC_392/a_36_216# INVX1_LOC_42/A 0.00fF
C43128 NAND2X1_LOC_726/Y NAND2X1_LOC_725/A 0.05fF
C43129 GATE_741 INVX1_LOC_282/Y 0.00fF
C43130 NOR2X1_LOC_503/A INVX1_LOC_78/A 0.02fF
C43131 NOR2X1_LOC_405/A NOR2X1_LOC_831/Y 0.04fF
C43132 NOR2X1_LOC_615/Y INVX1_LOC_172/A 0.01fF
C43133 INVX1_LOC_35/A NAND2X1_LOC_112/Y 0.03fF
C43134 INVX1_LOC_45/A NOR2X1_LOC_68/A 0.31fF
C43135 INVX1_LOC_200/Y NOR2X1_LOC_373/Y 0.01fF
C43136 NOR2X1_LOC_78/Y INVX1_LOC_280/A 0.46fF
C43137 NOR2X1_LOC_75/Y INVX1_LOC_113/Y 0.09fF
C43138 NAND2X1_LOC_30/Y NAND2X1_LOC_21/Y 2.28fF
C43139 NOR2X1_LOC_637/Y NOR2X1_LOC_590/A 0.04fF
C43140 INVX1_LOC_304/A NAND2X1_LOC_81/B 0.03fF
C43141 NOR2X1_LOC_242/A NOR2X1_LOC_78/B 0.10fF
C43142 INVX1_LOC_91/A NAND2X1_LOC_254/Y 0.15fF
C43143 NOR2X1_LOC_798/A NOR2X1_LOC_566/Y 0.01fF
C43144 NOR2X1_LOC_151/Y INVX1_LOC_78/A 0.03fF
C43145 D_INPUT_1 D_INPUT_0 0.23fF
C43146 NAND2X1_LOC_733/Y NAND2X1_LOC_866/A 0.02fF
C43147 NAND2X1_LOC_799/A NAND2X1_LOC_354/B 0.03fF
C43148 NAND2X1_LOC_741/B INVX1_LOC_300/Y 0.00fF
C43149 INVX1_LOC_143/A NOR2X1_LOC_440/B 0.07fF
C43150 INVX1_LOC_258/Y INVX1_LOC_280/Y 0.03fF
C43151 NOR2X1_LOC_454/Y NAND2X1_LOC_231/Y 0.04fF
C43152 NOR2X1_LOC_178/Y INVX1_LOC_30/Y 0.05fF
C43153 NOR2X1_LOC_218/A NOR2X1_LOC_142/Y 0.06fF
C43154 INVX1_LOC_83/A INVX1_LOC_53/A 0.17fF
C43155 NAND2X1_LOC_860/A INVX1_LOC_135/A 0.37fF
C43156 NAND2X1_LOC_67/Y INVX1_LOC_96/Y 0.08fF
C43157 NOR2X1_LOC_363/Y NOR2X1_LOC_127/Y 0.01fF
C43158 INVX1_LOC_49/Y NAND2X1_LOC_649/a_36_24# 0.00fF
C43159 INVX1_LOC_50/A NOR2X1_LOC_644/A 0.03fF
C43160 NAND2X1_LOC_564/A NAND2X1_LOC_551/A 0.15fF
C43161 INVX1_LOC_5/A NAND2X1_LOC_41/Y 0.03fF
C43162 NOR2X1_LOC_351/Y NOR2X1_LOC_155/A 0.00fF
C43163 NOR2X1_LOC_160/B NOR2X1_LOC_712/Y 0.00fF
C43164 NOR2X1_LOC_592/A NOR2X1_LOC_52/B 0.01fF
C43165 INVX1_LOC_135/A NOR2X1_LOC_634/Y 0.03fF
C43166 NAND2X1_LOC_212/Y INVX1_LOC_109/Y 0.01fF
C43167 NOR2X1_LOC_88/Y INVX1_LOC_118/A 0.07fF
C43168 NOR2X1_LOC_134/Y NAND2X1_LOC_464/Y 0.01fF
C43169 NOR2X1_LOC_67/A INVX1_LOC_1/A 0.10fF
C43170 INVX1_LOC_5/A NOR2X1_LOC_391/A 0.00fF
C43171 NAND2X1_LOC_581/Y INVX1_LOC_174/A 0.03fF
C43172 NOR2X1_LOC_269/Y INVX1_LOC_32/A 0.04fF
C43173 NOR2X1_LOC_82/A NOR2X1_LOC_515/a_36_216# 0.00fF
C43174 INVX1_LOC_59/A INVX1_LOC_316/Y 0.01fF
C43175 INVX1_LOC_315/Y NOR2X1_LOC_38/B 0.02fF
C43176 INVX1_LOC_37/A INVX1_LOC_272/A 0.07fF
C43177 NOR2X1_LOC_68/A INVX1_LOC_71/A 0.07fF
C43178 INVX1_LOC_161/Y NOR2X1_LOC_574/a_36_216# 0.00fF
C43179 NAND2X1_LOC_198/B NOR2X1_LOC_758/a_36_216# 0.10fF
C43180 INVX1_LOC_217/A NAND2X1_LOC_866/A 0.12fF
C43181 NOR2X1_LOC_92/Y INVX1_LOC_25/Y 0.07fF
C43182 INVX1_LOC_278/A INPUT_1 0.34fF
C43183 INVX1_LOC_6/A NOR2X1_LOC_278/Y 0.03fF
C43184 INVX1_LOC_24/A INVX1_LOC_41/Y 0.03fF
C43185 INVX1_LOC_11/A NOR2X1_LOC_352/Y 0.04fF
C43186 INVX1_LOC_6/Y NOR2X1_LOC_270/Y 0.03fF
C43187 NOR2X1_LOC_785/a_36_216# INVX1_LOC_57/A 0.02fF
C43188 INVX1_LOC_177/Y NOR2X1_LOC_577/Y 0.02fF
C43189 NAND2X1_LOC_190/Y INVX1_LOC_208/A 0.10fF
C43190 INVX1_LOC_84/A INVX1_LOC_118/A 0.10fF
C43191 INVX1_LOC_59/Y INVX1_LOC_3/Y 0.71fF
C43192 NOR2X1_LOC_222/Y NOR2X1_LOC_215/a_36_216# 0.00fF
C43193 INVX1_LOC_50/A NOR2X1_LOC_751/A 0.09fF
C43194 INVX1_LOC_33/Y NAND2X1_LOC_74/B 0.03fF
C43195 INVX1_LOC_24/A NAND2X1_LOC_593/Y 0.04fF
C43196 INVX1_LOC_88/A INVX1_LOC_53/Y 0.00fF
C43197 NAND2X1_LOC_254/Y NOR2X1_LOC_290/a_36_216# 0.00fF
C43198 NOR2X1_LOC_606/Y NOR2X1_LOC_709/A 0.01fF
C43199 INVX1_LOC_104/A NOR2X1_LOC_274/B 0.07fF
C43200 NOR2X1_LOC_15/Y NOR2X1_LOC_561/Y 0.25fF
C43201 NAND2X1_LOC_728/Y NAND2X1_LOC_354/B 0.12fF
C43202 NOR2X1_LOC_361/B NOR2X1_LOC_589/A 0.65fF
C43203 INVX1_LOC_38/A INVX1_LOC_29/A 0.17fF
C43204 NOR2X1_LOC_441/Y NOR2X1_LOC_131/A 0.00fF
C43205 NAND2X1_LOC_332/Y NOR2X1_LOC_338/Y 0.03fF
C43206 INVX1_LOC_88/A NOR2X1_LOC_665/A 0.91fF
C43207 NAND2X1_LOC_703/Y NAND2X1_LOC_808/A 0.28fF
C43208 NAND2X1_LOC_93/B INVX1_LOC_294/A 0.05fF
C43209 INVX1_LOC_135/A NAND2X1_LOC_473/A 0.04fF
C43210 INVX1_LOC_232/Y INVX1_LOC_31/A 0.41fF
C43211 INVX1_LOC_223/A INVX1_LOC_266/Y 0.00fF
C43212 NOR2X1_LOC_74/A NOR2X1_LOC_678/A 0.06fF
C43213 INVX1_LOC_286/Y NAND2X1_LOC_850/Y -0.02fF
C43214 NOR2X1_LOC_328/Y INVX1_LOC_211/A 0.01fF
C43215 INVX1_LOC_208/A NOR2X1_LOC_389/A 0.45fF
C43216 VDD INVX1_LOC_4/A 1.39fF
C43217 NOR2X1_LOC_315/Y NOR2X1_LOC_91/Y 0.02fF
C43218 INVX1_LOC_225/A NAND2X1_LOC_656/A 0.10fF
C43219 NOR2X1_LOC_186/Y NOR2X1_LOC_329/B 0.07fF
C43220 INVX1_LOC_5/A NAND2X1_LOC_709/a_36_24# 0.00fF
C43221 INVX1_LOC_239/A NAND2X1_LOC_624/A 0.02fF
C43222 INVX1_LOC_135/A NAND2X1_LOC_537/Y 0.10fF
C43223 NAND2X1_LOC_21/Y INVX1_LOC_49/A 0.05fF
C43224 INVX1_LOC_95/Y NOR2X1_LOC_55/a_36_216# 0.00fF
C43225 INVX1_LOC_34/A INVX1_LOC_77/A 0.17fF
C43226 INVX1_LOC_244/Y NOR2X1_LOC_52/B 0.00fF
C43227 INVX1_LOC_76/A INVX1_LOC_273/A 0.00fF
C43228 INVX1_LOC_17/A NAND2X1_LOC_656/Y 0.14fF
C43229 NAND2X1_LOC_198/B INVX1_LOC_168/A 0.05fF
C43230 NOR2X1_LOC_817/a_36_216# NOR2X1_LOC_332/A 0.01fF
C43231 NOR2X1_LOC_67/A NOR2X1_LOC_384/Y 1.94fF
C43232 NOR2X1_LOC_778/B NOR2X1_LOC_703/B 0.03fF
C43233 NOR2X1_LOC_795/Y NOR2X1_LOC_500/A 0.10fF
C43234 NAND2X1_LOC_633/Y INVX1_LOC_78/A 0.07fF
C43235 NAND2X1_LOC_573/Y NOR2X1_LOC_329/B 0.50fF
C43236 NOR2X1_LOC_67/A NOR2X1_LOC_522/a_36_216# 0.01fF
C43237 INVX1_LOC_94/A NOR2X1_LOC_493/B 0.00fF
C43238 INVX1_LOC_24/A NOR2X1_LOC_538/Y 0.06fF
C43239 NOR2X1_LOC_142/Y INVX1_LOC_155/Y 0.03fF
C43240 INVX1_LOC_104/A NOR2X1_LOC_577/Y 0.50fF
C43241 INVX1_LOC_30/A INVX1_LOC_1/Y 0.26fF
C43242 NAND2X1_LOC_377/a_36_24# INVX1_LOC_89/A 0.00fF
C43243 INVX1_LOC_256/A NOR2X1_LOC_106/A 0.04fF
C43244 INVX1_LOC_226/Y INVX1_LOC_72/A 0.00fF
C43245 INVX1_LOC_64/A NOR2X1_LOC_337/Y 0.02fF
C43246 INVX1_LOC_95/Y INVX1_LOC_57/A 0.15fF
C43247 INVX1_LOC_41/A INVX1_LOC_176/Y 0.01fF
C43248 INVX1_LOC_71/Y INVX1_LOC_42/A 0.01fF
C43249 INVX1_LOC_118/A INVX1_LOC_15/A 0.17fF
C43250 INVX1_LOC_35/A NOR2X1_LOC_78/A 0.19fF
C43251 NOR2X1_LOC_419/Y NOR2X1_LOC_721/A 0.01fF
C43252 NOR2X1_LOC_91/A NAND2X1_LOC_287/B 0.10fF
C43253 NOR2X1_LOC_392/B INVX1_LOC_8/A 0.10fF
C43254 NAND2X1_LOC_778/Y NOR2X1_LOC_167/Y 0.30fF
C43255 NOR2X1_LOC_226/A NOR2X1_LOC_262/Y 0.01fF
C43256 INVX1_LOC_146/Y NAND2X1_LOC_420/a_36_24# 0.01fF
C43257 NOR2X1_LOC_598/B NOR2X1_LOC_486/Y 0.07fF
C43258 INVX1_LOC_58/A NOR2X1_LOC_300/a_36_216# 0.00fF
C43259 INVX1_LOC_208/A NOR2X1_LOC_596/A 0.01fF
C43260 INVX1_LOC_124/A INVX1_LOC_34/A 0.07fF
C43261 NOR2X1_LOC_500/A NOR2X1_LOC_614/Y 0.02fF
C43262 NAND2X1_LOC_63/Y INVX1_LOC_84/A 0.03fF
C43263 NOR2X1_LOC_455/Y INVX1_LOC_188/Y 0.04fF
C43264 NOR2X1_LOC_331/B NAND2X1_LOC_454/Y 0.07fF
C43265 NOR2X1_LOC_305/Y INVX1_LOC_57/A 0.07fF
C43266 INVX1_LOC_72/A INVX1_LOC_10/A 0.34fF
C43267 INVX1_LOC_284/Y NAND2X1_LOC_866/B 0.07fF
C43268 NOR2X1_LOC_503/A NOR2X1_LOC_503/Y 0.04fF
C43269 D_INPUT_1 NOR2X1_LOC_266/B 0.03fF
C43270 INVX1_LOC_64/A NOR2X1_LOC_56/Y 0.03fF
C43271 INVX1_LOC_93/A NOR2X1_LOC_45/B 0.07fF
C43272 INVX1_LOC_279/A NOR2X1_LOC_598/a_36_216# 0.00fF
C43273 INVX1_LOC_85/A INVX1_LOC_266/Y 0.03fF
C43274 NOR2X1_LOC_15/Y NOR2X1_LOC_167/Y 2.28fF
C43275 NOR2X1_LOC_763/Y INVX1_LOC_18/A 0.07fF
C43276 NAND2X1_LOC_552/a_36_24# INVX1_LOC_41/Y 0.00fF
C43277 INVX1_LOC_88/A NOR2X1_LOC_113/B 0.01fF
C43278 NOR2X1_LOC_716/B NAND2X1_LOC_860/Y 0.03fF
C43279 NOR2X1_LOC_613/Y NOR2X1_LOC_528/Y 0.00fF
C43280 INVX1_LOC_276/A INVX1_LOC_221/A 0.66fF
C43281 INVX1_LOC_314/Y INVX1_LOC_137/Y 0.02fF
C43282 INVX1_LOC_53/A INVX1_LOC_46/A 0.13fF
C43283 NAND2X1_LOC_563/Y INVX1_LOC_216/A 0.04fF
C43284 INVX1_LOC_202/Y INVX1_LOC_270/A 0.01fF
C43285 NAND2X1_LOC_99/A NOR2X1_LOC_271/Y 0.24fF
C43286 NOR2X1_LOC_334/Y NAND2X1_LOC_93/B 0.07fF
C43287 NAND2X1_LOC_721/B INVX1_LOC_90/A 0.03fF
C43288 INVX1_LOC_247/Y INVX1_LOC_97/A 0.14fF
C43289 INVX1_LOC_185/Y NAND2X1_LOC_850/Y 0.00fF
C43290 NAND2X1_LOC_374/Y NOR2X1_LOC_52/B 0.07fF
C43291 INVX1_LOC_203/A NAND2X1_LOC_254/Y 0.11fF
C43292 INVX1_LOC_38/A NOR2X1_LOC_318/a_36_216# 0.00fF
C43293 INVX1_LOC_41/A INVX1_LOC_25/Y 0.23fF
C43294 NAND2X1_LOC_35/Y NAND2X1_LOC_244/A 0.01fF
C43295 INVX1_LOC_64/A INVX1_LOC_146/Y -0.00fF
C43296 NAND2X1_LOC_787/A NAND2X1_LOC_721/A 0.11fF
C43297 NOR2X1_LOC_759/Y NOR2X1_LOC_366/Y 0.02fF
C43298 INVX1_LOC_94/A INVX1_LOC_150/A 0.01fF
C43299 INVX1_LOC_64/A VDD 4.31fF
C43300 INVX1_LOC_178/A INVX1_LOC_187/A 0.01fF
C43301 NOR2X1_LOC_252/Y NAND2X1_LOC_483/Y 0.05fF
C43302 INVX1_LOC_102/A INVX1_LOC_19/A 0.07fF
C43303 NOR2X1_LOC_470/A INVX1_LOC_113/Y 0.01fF
C43304 INVX1_LOC_202/A NOR2X1_LOC_366/Y 0.14fF
C43305 NOR2X1_LOC_510/Y INVX1_LOC_147/Y 0.01fF
C43306 INVX1_LOC_83/A INVX1_LOC_184/A 0.04fF
C43307 INVX1_LOC_22/Y INVX1_LOC_31/Y 0.34fF
C43308 INVX1_LOC_13/Y NAND2X1_LOC_465/A 0.01fF
C43309 NAND2X1_LOC_726/Y NAND2X1_LOC_308/Y 0.01fF
C43310 D_INPUT_0 D_INPUT_2 0.64fF
C43311 INVX1_LOC_64/A NAND2X1_LOC_800/A 0.04fF
C43312 INVX1_LOC_178/Y NOR2X1_LOC_663/A 0.01fF
C43313 NOR2X1_LOC_424/Y INVX1_LOC_113/Y 0.01fF
C43314 INVX1_LOC_263/A NOR2X1_LOC_348/B 0.00fF
C43315 NOR2X1_LOC_690/A NOR2X1_LOC_86/A 0.03fF
C43316 NOR2X1_LOC_155/A NOR2X1_LOC_471/a_36_216# 0.00fF
C43317 NOR2X1_LOC_510/Y INVX1_LOC_20/A 0.18fF
C43318 NOR2X1_LOC_516/B NOR2X1_LOC_844/A 0.03fF
C43319 NOR2X1_LOC_742/A INVX1_LOC_30/A 0.03fF
C43320 NOR2X1_LOC_78/B NOR2X1_LOC_634/B 0.16fF
C43321 INVX1_LOC_104/A INVX1_LOC_22/A 0.14fF
C43322 NAND2X1_LOC_477/A INVX1_LOC_25/Y 0.10fF
C43323 NOR2X1_LOC_584/Y INVX1_LOC_261/Y 0.80fF
C43324 NOR2X1_LOC_590/A NOR2X1_LOC_548/A 0.00fF
C43325 INVX1_LOC_12/A INVX1_LOC_284/A 0.14fF
C43326 INVX1_LOC_45/A INVX1_LOC_147/A 0.42fF
C43327 INVX1_LOC_18/A NOR2X1_LOC_703/A 0.03fF
C43328 INVX1_LOC_27/A NOR2X1_LOC_603/Y 0.03fF
C43329 NAND2X1_LOC_571/Y NOR2X1_LOC_24/Y 0.01fF
C43330 NAND2X1_LOC_322/a_36_24# NOR2X1_LOC_317/B 0.00fF
C43331 INVX1_LOC_307/Y NOR2X1_LOC_383/B 0.08fF
C43332 INVX1_LOC_84/A NAND2X1_LOC_618/Y 0.07fF
C43333 NAND2X1_LOC_149/Y NOR2X1_LOC_683/Y 0.06fF
C43334 NOR2X1_LOC_213/a_36_216# NOR2X1_LOC_220/A 0.01fF
C43335 INVX1_LOC_200/Y INVX1_LOC_54/A 0.00fF
C43336 NOR2X1_LOC_398/Y INVX1_LOC_25/Y 0.04fF
C43337 NOR2X1_LOC_160/B NAND2X1_LOC_695/a_36_24# 0.01fF
C43338 NOR2X1_LOC_453/Y INVX1_LOC_115/Y 0.01fF
C43339 NOR2X1_LOC_513/Y NOR2X1_LOC_45/B 0.01fF
C43340 NOR2X1_LOC_457/A NOR2X1_LOC_318/B 0.46fF
C43341 INVX1_LOC_291/A NOR2X1_LOC_654/A 0.10fF
C43342 NAND2X1_LOC_397/a_36_24# NAND2X1_LOC_659/B 0.00fF
C43343 INVX1_LOC_226/Y NOR2X1_LOC_537/Y 0.07fF
C43344 NOR2X1_LOC_716/B NAND2X1_LOC_861/Y 0.10fF
C43345 NAND2X1_LOC_662/Y INVX1_LOC_266/Y 0.03fF
C43346 NAND2X1_LOC_736/Y NOR2X1_LOC_299/Y 10.63fF
C43347 INVX1_LOC_226/Y NAND2X1_LOC_338/B 1.59fF
C43348 NOR2X1_LOC_502/Y NOR2X1_LOC_78/A 0.01fF
C43349 NAND2X1_LOC_223/A NOR2X1_LOC_673/B 0.02fF
C43350 NAND2X1_LOC_63/Y INVX1_LOC_15/A 0.09fF
C43351 INVX1_LOC_278/A INVX1_LOC_118/A 0.64fF
C43352 INVX1_LOC_135/A NOR2X1_LOC_516/Y 0.09fF
C43353 NOR2X1_LOC_723/Y INVX1_LOC_311/A 0.04fF
C43354 NOR2X1_LOC_829/A NAND2X1_LOC_771/a_36_24# 0.00fF
C43355 NOR2X1_LOC_440/Y NOR2X1_LOC_709/A 0.01fF
C43356 NOR2X1_LOC_155/A NOR2X1_LOC_748/A 0.05fF
C43357 NOR2X1_LOC_15/Y INVX1_LOC_76/A 8.80fF
C43358 NOR2X1_LOC_214/B INVX1_LOC_63/Y 0.01fF
C43359 INVX1_LOC_182/Y NOR2X1_LOC_363/a_36_216# 0.00fF
C43360 INVX1_LOC_14/A INVX1_LOC_126/A 0.03fF
C43361 INVX1_LOC_23/A NOR2X1_LOC_809/B 0.02fF
C43362 NOR2X1_LOC_92/Y NAND2X1_LOC_453/A 0.08fF
C43363 GATE_662 NAND2X1_LOC_451/Y 0.05fF
C43364 NOR2X1_LOC_361/B INVX1_LOC_20/A 0.03fF
C43365 D_INPUT_1 INVX1_LOC_46/Y 0.08fF
C43366 NAND2X1_LOC_853/Y NAND2X1_LOC_863/B 0.83fF
C43367 NOR2X1_LOC_590/A NAND2X1_LOC_86/Y 0.01fF
C43368 INVX1_LOC_305/A NOR2X1_LOC_9/Y 0.00fF
C43369 INVX1_LOC_90/A INVX1_LOC_8/A 0.02fF
C43370 NOR2X1_LOC_770/B NOR2X1_LOC_770/Y 0.00fF
C43371 NOR2X1_LOC_234/Y INVX1_LOC_89/A 0.01fF
C43372 NAND2X1_LOC_715/B NOR2X1_LOC_351/Y 0.09fF
C43373 INVX1_LOC_263/A INVX1_LOC_22/A 0.08fF
C43374 INVX1_LOC_13/Y NOR2X1_LOC_652/a_36_216# 0.01fF
C43375 NAND2X1_LOC_717/Y NOR2X1_LOC_298/Y 3.48fF
C43376 NAND2X1_LOC_615/a_36_24# INVX1_LOC_69/A 0.00fF
C43377 INVX1_LOC_293/Y INVX1_LOC_23/Y 0.09fF
C43378 D_INPUT_0 NOR2X1_LOC_529/Y 0.02fF
C43379 INVX1_LOC_103/A NOR2X1_LOC_314/Y 0.06fF
C43380 INVX1_LOC_5/A NOR2X1_LOC_629/Y 0.03fF
C43381 INVX1_LOC_233/A INVX1_LOC_92/A 0.02fF
C43382 NOR2X1_LOC_318/B INVX1_LOC_30/A 0.10fF
C43383 NOR2X1_LOC_355/A INVX1_LOC_111/Y 0.00fF
C43384 INVX1_LOC_182/Y INVX1_LOC_155/A 0.00fF
C43385 INVX1_LOC_14/A NOR2X1_LOC_111/A 0.02fF
C43386 INVX1_LOC_41/A NOR2X1_LOC_439/B 0.03fF
C43387 NOR2X1_LOC_653/Y NOR2X1_LOC_280/a_36_216# 0.00fF
C43388 NOR2X1_LOC_78/B INVX1_LOC_83/A 0.13fF
C43389 INVX1_LOC_209/Y NOR2X1_LOC_313/a_36_216# 0.00fF
C43390 INVX1_LOC_77/A INPUT_0 0.17fF
C43391 NAND2X1_LOC_725/A INVX1_LOC_241/Y 0.02fF
C43392 D_INPUT_0 NOR2X1_LOC_620/B 0.02fF
C43393 INVX1_LOC_30/A INVX1_LOC_93/Y 2.25fF
C43394 INVX1_LOC_41/A INVX1_LOC_75/A 0.09fF
C43395 NAND2X1_LOC_588/a_36_24# INVX1_LOC_83/A 0.00fF
C43396 INVX1_LOC_116/A INVX1_LOC_286/A 0.01fF
C43397 NAND2X1_LOC_537/Y NOR2X1_LOC_152/A 0.04fF
C43398 INVX1_LOC_103/A INVX1_LOC_117/A 0.10fF
C43399 INVX1_LOC_23/Y NAND2X1_LOC_74/B 0.17fF
C43400 INVX1_LOC_201/Y INVX1_LOC_75/A 0.35fF
C43401 NAND2X1_LOC_735/B NOR2X1_LOC_32/Y 0.03fF
C43402 INVX1_LOC_135/A INVX1_LOC_172/Y 0.02fF
C43403 NOR2X1_LOC_389/A NAND2X1_LOC_211/Y 0.01fF
C43404 NOR2X1_LOC_520/B NOR2X1_LOC_188/A 0.72fF
C43405 NOR2X1_LOC_798/A INVX1_LOC_92/A 0.03fF
C43406 NOR2X1_LOC_589/A NAND2X1_LOC_573/A 0.02fF
C43407 INVX1_LOC_34/A NAND2X1_LOC_832/Y 0.03fF
C43408 NOR2X1_LOC_392/Y NOR2X1_LOC_23/a_36_216# 0.00fF
C43409 INVX1_LOC_124/A INVX1_LOC_131/A 0.23fF
C43410 NAND2X1_LOC_357/B NOR2X1_LOC_322/Y 0.44fF
C43411 NAND2X1_LOC_618/Y INVX1_LOC_15/A 0.03fF
C43412 INVX1_LOC_206/Y NOR2X1_LOC_577/Y 0.01fF
C43413 NOR2X1_LOC_530/a_36_216# NOR2X1_LOC_813/Y 0.01fF
C43414 INVX1_LOC_1/A NOR2X1_LOC_729/A 0.03fF
C43415 NOR2X1_LOC_11/Y INVX1_LOC_296/Y 0.41fF
C43416 INVX1_LOC_56/Y NOR2X1_LOC_76/A 0.04fF
C43417 INVX1_LOC_314/Y INVX1_LOC_91/A 0.08fF
C43418 NOR2X1_LOC_332/A NAND2X1_LOC_41/Y 0.01fF
C43419 INVX1_LOC_292/A INVX1_LOC_117/A 0.01fF
C43420 INVX1_LOC_313/Y NOR2X1_LOC_500/Y 0.67fF
C43421 INVX1_LOC_89/A NOR2X1_LOC_507/A 0.01fF
C43422 INVX1_LOC_119/A INVX1_LOC_144/A 0.01fF
C43423 NAND2X1_LOC_703/Y INVX1_LOC_92/A 0.23fF
C43424 INVX1_LOC_124/A INPUT_0 0.07fF
C43425 INVX1_LOC_30/A NAND2X1_LOC_721/A 0.11fF
C43426 NOR2X1_LOC_833/B NOR2X1_LOC_748/A 0.01fF
C43427 INVX1_LOC_18/A NAND2X1_LOC_650/B 0.44fF
C43428 INVX1_LOC_26/A INVX1_LOC_32/A 0.13fF
C43429 INVX1_LOC_235/A NAND2X1_LOC_574/A 0.00fF
C43430 INVX1_LOC_206/Y NOR2X1_LOC_348/B 0.17fF
C43431 NOR2X1_LOC_303/Y INVX1_LOC_247/A 0.03fF
C43432 NOR2X1_LOC_604/Y INVX1_LOC_12/A 0.04fF
C43433 INVX1_LOC_130/Y VDD 0.47fF
C43434 INVX1_LOC_39/A INVX1_LOC_84/A 0.10fF
C43435 NOR2X1_LOC_355/A NOR2X1_LOC_137/A 0.14fF
C43436 NOR2X1_LOC_191/A NOR2X1_LOC_74/A 0.11fF
C43437 INVX1_LOC_36/A INVX1_LOC_202/Y 0.01fF
C43438 NOR2X1_LOC_591/A INVX1_LOC_42/A 0.02fF
C43439 INVX1_LOC_313/Y INVX1_LOC_10/A 0.01fF
C43440 INVX1_LOC_136/A INVX1_LOC_33/Y 0.01fF
C43441 D_INPUT_5 INVX1_LOC_173/A 0.01fF
C43442 NOR2X1_LOC_710/B NOR2X1_LOC_155/A 0.03fF
C43443 NAND2X1_LOC_866/B NOR2X1_LOC_525/Y 0.01fF
C43444 NAND2X1_LOC_454/Y NOR2X1_LOC_449/A 0.01fF
C43445 INVX1_LOC_278/A NAND2X1_LOC_455/B 0.34fF
C43446 INVX1_LOC_2/A INVX1_LOC_123/A 0.10fF
C43447 NAND2X1_LOC_863/Y VDD 0.01fF
C43448 NOR2X1_LOC_348/B NOR2X1_LOC_600/Y 0.63fF
C43449 NOR2X1_LOC_254/Y INVX1_LOC_247/A 0.69fF
C43450 NOR2X1_LOC_214/a_36_216# NOR2X1_LOC_357/Y 0.01fF
C43451 NAND2X1_LOC_218/B NAND2X1_LOC_8/a_36_24# 0.00fF
C43452 INVX1_LOC_40/A INVX1_LOC_201/A 0.02fF
C43453 INVX1_LOC_61/Y INVX1_LOC_89/Y 0.02fF
C43454 NOR2X1_LOC_312/Y NAND2X1_LOC_807/Y 0.04fF
C43455 NOR2X1_LOC_68/A NOR2X1_LOC_331/B 0.07fF
C43456 NAND2X1_LOC_296/a_36_24# NOR2X1_LOC_416/A 0.00fF
C43457 NOR2X1_LOC_208/Y INVX1_LOC_202/Y 0.03fF
C43458 INVX1_LOC_79/Y INVX1_LOC_9/A 0.01fF
C43459 NOR2X1_LOC_778/B INVX1_LOC_91/A 0.12fF
C43460 NAND2X1_LOC_793/Y INVX1_LOC_285/A 0.09fF
C43461 INVX1_LOC_206/Y INVX1_LOC_22/A 0.03fF
C43462 INVX1_LOC_12/A NOR2X1_LOC_384/A 0.01fF
C43463 INVX1_LOC_30/A INVX1_LOC_117/Y 0.04fF
C43464 NOR2X1_LOC_459/B VDD -0.00fF
C43465 NOR2X1_LOC_770/B INVX1_LOC_37/A 0.01fF
C43466 NOR2X1_LOC_48/B NOR2X1_LOC_406/A 0.08fF
C43467 NOR2X1_LOC_799/B NOR2X1_LOC_537/Y 0.01fF
C43468 NOR2X1_LOC_500/A NOR2X1_LOC_499/B 0.12fF
C43469 NOR2X1_LOC_78/A NOR2X1_LOC_121/A 0.01fF
C43470 INVX1_LOC_96/Y INVX1_LOC_76/A 0.18fF
C43471 NAND2X1_LOC_477/A NAND2X1_LOC_453/A 0.14fF
C43472 INVX1_LOC_24/A INVX1_LOC_185/A 0.03fF
C43473 NAND2X1_LOC_363/B INVX1_LOC_87/A 0.01fF
C43474 INVX1_LOC_22/A NOR2X1_LOC_600/Y 0.15fF
C43475 NAND2X1_LOC_350/B NAND2X1_LOC_469/B 0.11fF
C43476 INVX1_LOC_280/Y INVX1_LOC_20/A 0.03fF
C43477 NOR2X1_LOC_68/A NOR2X1_LOC_592/B 0.03fF
C43478 INVX1_LOC_21/A D_INPUT_5 0.01fF
C43479 NOR2X1_LOC_495/Y INVX1_LOC_54/A 0.01fF
C43480 VDD INVX1_LOC_44/Y 0.00fF
C43481 INVX1_LOC_61/A NOR2X1_LOC_88/Y 0.12fF
C43482 NOR2X1_LOC_383/B INVX1_LOC_29/Y 1.01fF
C43483 NOR2X1_LOC_78/B INVX1_LOC_46/A 0.44fF
C43484 INVX1_LOC_299/A NOR2X1_LOC_640/B 0.01fF
C43485 NAND2X1_LOC_840/B INVX1_LOC_76/A 0.07fF
C43486 NOR2X1_LOC_711/A INVX1_LOC_85/Y 0.06fF
C43487 NOR2X1_LOC_500/A NOR2X1_LOC_862/B 0.10fF
C43488 INVX1_LOC_34/A INVX1_LOC_9/A 0.07fF
C43489 VDD NAND2X1_LOC_850/Y 0.53fF
C43490 INVX1_LOC_271/A NAND2X1_LOC_678/a_36_24# 0.02fF
C43491 INVX1_LOC_217/A INVX1_LOC_119/Y 0.04fF
C43492 INVX1_LOC_24/A NAND2X1_LOC_809/a_36_24# 0.01fF
C43493 NOR2X1_LOC_598/B INVX1_LOC_275/Y 0.02fF
C43494 INVX1_LOC_83/A NOR2X1_LOC_311/Y 0.01fF
C43495 INVX1_LOC_123/A INPUT_1 0.07fF
C43496 NOR2X1_LOC_598/B NOR2X1_LOC_748/A 0.19fF
C43497 NAND2X1_LOC_860/Y NAND2X1_LOC_633/Y 0.04fF
C43498 INVX1_LOC_205/A NOR2X1_LOC_814/A 0.01fF
C43499 NAND2X1_LOC_209/a_36_24# NOR2X1_LOC_467/A 0.00fF
C43500 NAND2X1_LOC_562/B NOR2X1_LOC_629/Y 0.01fF
C43501 NOR2X1_LOC_162/Y NAND2X1_LOC_93/B 0.02fF
C43502 INVX1_LOC_225/Y INVX1_LOC_290/Y 0.05fF
C43503 INVX1_LOC_33/A NOR2X1_LOC_634/A 0.08fF
C43504 NAND2X1_LOC_573/A INVX1_LOC_20/A 0.01fF
C43505 INVX1_LOC_50/Y NOR2X1_LOC_668/Y 0.01fF
C43506 NOR2X1_LOC_264/Y NOR2X1_LOC_624/B 0.01fF
C43507 NOR2X1_LOC_201/A INVX1_LOC_50/Y 0.08fF
C43508 NOR2X1_LOC_162/Y NAND2X1_LOC_425/Y 0.13fF
C43509 NAND2X1_LOC_392/Y INVX1_LOC_46/A 0.05fF
C43510 INVX1_LOC_156/Y VDD 0.26fF
C43511 INVX1_LOC_28/A NAND2X1_LOC_655/A 0.07fF
C43512 INVX1_LOC_14/A INVX1_LOC_90/Y 0.01fF
C43513 NOR2X1_LOC_666/Y INVX1_LOC_271/Y 0.11fF
C43514 NAND2X1_LOC_123/Y INVX1_LOC_91/A 0.02fF
C43515 NOR2X1_LOC_708/Y NOR2X1_LOC_708/A 0.04fF
C43516 INVX1_LOC_72/A INVX1_LOC_12/A 1.55fF
C43517 NOR2X1_LOC_160/B INVX1_LOC_251/A 0.05fF
C43518 NOR2X1_LOC_576/B INVX1_LOC_76/A 0.02fF
C43519 INVX1_LOC_172/Y INVX1_LOC_280/A 0.01fF
C43520 NOR2X1_LOC_294/Y NOR2X1_LOC_346/A 0.06fF
C43521 NOR2X1_LOC_329/B NAND2X1_LOC_642/Y 1.06fF
C43522 NAND2X1_LOC_198/B INVX1_LOC_272/A 0.33fF
C43523 INVX1_LOC_50/Y INVX1_LOC_23/A 0.03fF
C43524 NOR2X1_LOC_372/Y NAND2X1_LOC_254/Y 0.01fF
C43525 INVX1_LOC_217/A INVX1_LOC_284/A 0.03fF
C43526 INVX1_LOC_256/A NOR2X1_LOC_334/Y 0.19fF
C43527 INVX1_LOC_62/Y NAND2X1_LOC_207/B 0.07fF
C43528 INVX1_LOC_187/A INVX1_LOC_140/A 0.05fF
C43529 INVX1_LOC_28/A NAND2X1_LOC_468/B 0.01fF
C43530 NAND2X1_LOC_861/Y NAND2X1_LOC_633/Y 0.04fF
C43531 INVX1_LOC_132/A NOR2X1_LOC_691/B 0.50fF
C43532 NOR2X1_LOC_434/Y NOR2X1_LOC_434/A 0.00fF
C43533 NOR2X1_LOC_798/A INVX1_LOC_53/A 0.04fF
C43534 NAND2X1_LOC_9/Y NOR2X1_LOC_242/A 0.03fF
C43535 INVX1_LOC_35/A NOR2X1_LOC_186/Y 0.10fF
C43536 NAND2X1_LOC_773/Y INVX1_LOC_57/A 0.03fF
C43537 INVX1_LOC_304/Y INVX1_LOC_119/Y 0.07fF
C43538 NOR2X1_LOC_250/Y NOR2X1_LOC_318/A 0.09fF
C43539 NOR2X1_LOC_510/Y INVX1_LOC_64/A 2.27fF
C43540 NOR2X1_LOC_386/a_36_216# INPUT_4 0.00fF
C43541 NOR2X1_LOC_361/Y NOR2X1_LOC_127/Y 0.01fF
C43542 NAND2X1_LOC_807/Y NAND2X1_LOC_287/B 0.24fF
C43543 NAND2X1_LOC_703/Y INVX1_LOC_53/A 0.07fF
C43544 INVX1_LOC_266/A INVX1_LOC_23/A 0.01fF
C43545 NAND2X1_LOC_323/B NOR2X1_LOC_445/B 0.14fF
C43546 INVX1_LOC_141/Y INVX1_LOC_94/Y 0.00fF
C43547 NOR2X1_LOC_288/A NOR2X1_LOC_691/B 0.11fF
C43548 INVX1_LOC_33/A INVX1_LOC_29/A 0.58fF
C43549 INVX1_LOC_233/Y INVX1_LOC_258/Y 0.07fF
C43550 INVX1_LOC_149/Y INVX1_LOC_19/A 0.00fF
C43551 INPUT_3 INVX1_LOC_26/A 0.19fF
C43552 INVX1_LOC_61/A INVX1_LOC_15/A 0.04fF
C43553 NAND2X1_LOC_319/A INVX1_LOC_54/A 0.63fF
C43554 INVX1_LOC_35/A NAND2X1_LOC_573/Y 0.07fF
C43555 NAND2X1_LOC_787/B INVX1_LOC_284/A 0.00fF
C43556 INVX1_LOC_10/A NOR2X1_LOC_506/Y 0.34fF
C43557 INVX1_LOC_58/A INVX1_LOC_103/A 0.17fF
C43558 INVX1_LOC_30/A INVX1_LOC_87/A 0.03fF
C43559 NOR2X1_LOC_93/Y INVX1_LOC_5/A 0.01fF
C43560 INVX1_LOC_282/A VDD 0.43fF
C43561 NAND2X1_LOC_807/Y NAND2X1_LOC_808/a_36_24# 0.01fF
C43562 INVX1_LOC_230/Y NOR2X1_LOC_646/B 0.03fF
C43563 INVX1_LOC_36/A NOR2X1_LOC_278/Y 0.51fF
C43564 NAND2X1_LOC_67/a_36_24# INVX1_LOC_5/A 0.00fF
C43565 INVX1_LOC_17/A NOR2X1_LOC_717/A 0.01fF
C43566 INVX1_LOC_135/A NOR2X1_LOC_487/Y 0.04fF
C43567 NOR2X1_LOC_335/B INVX1_LOC_14/Y 0.02fF
C43568 INVX1_LOC_64/A NOR2X1_LOC_361/B 0.49fF
C43569 INVX1_LOC_58/A INVX1_LOC_292/A 0.10fF
C43570 NOR2X1_LOC_267/A NOR2X1_LOC_278/Y 0.04fF
C43571 INVX1_LOC_136/A INVX1_LOC_23/Y 0.17fF
C43572 INVX1_LOC_269/A INVX1_LOC_5/A 0.10fF
C43573 INVX1_LOC_136/A NAND2X1_LOC_72/a_36_24# 0.06fF
C43574 NAND2X1_LOC_861/Y INVX1_LOC_71/Y 0.02fF
C43575 NOR2X1_LOC_709/A NOR2X1_LOC_89/A 0.49fF
C43576 NAND2X1_LOC_799/Y NOR2X1_LOC_48/B 0.01fF
C43577 NAND2X1_LOC_740/Y NAND2X1_LOC_303/Y 0.10fF
C43578 INVX1_LOC_232/A INVX1_LOC_293/Y -0.02fF
C43579 NAND2X1_LOC_563/a_36_24# NOR2X1_LOC_660/Y -0.03fF
C43580 INVX1_LOC_64/Y NAND2X1_LOC_291/B 0.03fF
C43581 NOR2X1_LOC_599/A INVX1_LOC_296/Y 0.03fF
C43582 NAND2X1_LOC_809/A NAND2X1_LOC_810/B 0.09fF
C43583 INVX1_LOC_272/Y NAND2X1_LOC_502/a_36_24# 0.00fF
C43584 NAND2X1_LOC_338/B INVX1_LOC_12/A 0.03fF
C43585 INVX1_LOC_89/A NOR2X1_LOC_155/A 0.07fF
C43586 NOR2X1_LOC_624/A INVX1_LOC_15/A -0.02fF
C43587 INVX1_LOC_266/Y INVX1_LOC_290/Y 0.17fF
C43588 NOR2X1_LOC_91/Y NAND2X1_LOC_99/A 0.06fF
C43589 INVX1_LOC_6/A INVX1_LOC_129/Y 0.00fF
C43590 INVX1_LOC_35/A NOR2X1_LOC_45/Y 0.03fF
C43591 NAND2X1_LOC_562/Y INVX1_LOC_15/A 0.02fF
C43592 INVX1_LOC_147/A NOR2X1_LOC_331/B 0.42fF
C43593 NOR2X1_LOC_440/Y INVX1_LOC_294/A 0.01fF
C43594 INVX1_LOC_153/Y INVX1_LOC_4/A 0.10fF
C43595 INVX1_LOC_313/Y INVX1_LOC_307/A 0.02fF
C43596 NOR2X1_LOC_813/Y NOR2X1_LOC_86/a_36_216# 0.01fF
C43597 INVX1_LOC_179/Y INVX1_LOC_99/A 0.01fF
C43598 INVX1_LOC_269/A INVX1_LOC_178/A 0.05fF
C43599 NAND2X1_LOC_705/Y NAND2X1_LOC_706/Y 0.18fF
C43600 NAND2X1_LOC_374/Y NAND2X1_LOC_254/Y 0.57fF
C43601 NAND2X1_LOC_808/A INVX1_LOC_119/Y 0.02fF
C43602 NAND2X1_LOC_662/Y INVX1_LOC_19/A 0.07fF
C43603 NOR2X1_LOC_15/Y INVX1_LOC_163/A 0.24fF
C43604 INVX1_LOC_232/A NAND2X1_LOC_74/B 0.26fF
C43605 INPUT_0 INVX1_LOC_9/A 0.22fF
C43606 NOR2X1_LOC_503/A NAND2X1_LOC_802/Y 0.05fF
C43607 INVX1_LOC_149/A INVX1_LOC_32/A 0.07fF
C43608 NOR2X1_LOC_60/a_36_216# INVX1_LOC_63/A 0.01fF
C43609 NOR2X1_LOC_589/A NAND2X1_LOC_81/B 0.08fF
C43610 INVX1_LOC_8/A NAND2X1_LOC_223/A 0.46fF
C43611 INVX1_LOC_298/Y INVX1_LOC_33/A 0.03fF
C43612 INVX1_LOC_177/A INVX1_LOC_4/A 0.03fF
C43613 INVX1_LOC_25/A INVX1_LOC_181/Y 0.03fF
C43614 NOR2X1_LOC_383/Y NAND2X1_LOC_74/B 0.03fF
C43615 NOR2X1_LOC_164/Y INVX1_LOC_46/A 0.03fF
C43616 INVX1_LOC_31/A INVX1_LOC_50/Y 0.18fF
C43617 NAND2X1_LOC_469/B NAND2X1_LOC_211/Y 2.08fF
C43618 NAND2X1_LOC_642/Y NOR2X1_LOC_107/a_36_216# 0.00fF
C43619 NOR2X1_LOC_286/Y INVX1_LOC_1/A 0.07fF
C43620 NOR2X1_LOC_202/a_36_216# NOR2X1_LOC_205/Y 0.00fF
C43621 INVX1_LOC_73/A NOR2X1_LOC_831/B 0.03fF
C43622 NAND2X1_LOC_267/B INVX1_LOC_20/A 0.02fF
C43623 NOR2X1_LOC_750/Y NAND2X1_LOC_656/A 0.16fF
C43624 NOR2X1_LOC_489/B NAND2X1_LOC_364/A 0.01fF
C43625 INVX1_LOC_33/A NOR2X1_LOC_318/a_36_216# 0.00fF
C43626 NOR2X1_LOC_309/Y NOR2X1_LOC_278/Y 0.09fF
C43627 INVX1_LOC_24/A NOR2X1_LOC_754/Y 0.01fF
C43628 NOR2X1_LOC_542/B INVX1_LOC_117/A 0.15fF
C43629 NOR2X1_LOC_590/A NOR2X1_LOC_173/Y 0.03fF
C43630 INVX1_LOC_90/A NOR2X1_LOC_258/Y 0.02fF
C43631 INVX1_LOC_148/A NOR2X1_LOC_814/A 0.02fF
C43632 NOR2X1_LOC_783/A NOR2X1_LOC_796/B 0.01fF
C43633 D_INPUT_1 INVX1_LOC_49/A 0.10fF
C43634 NOR2X1_LOC_391/A INVX1_LOC_42/A 0.03fF
C43635 INVX1_LOC_75/A NAND2X1_LOC_574/A -0.04fF
C43636 NOR2X1_LOC_6/B NOR2X1_LOC_668/Y 0.01fF
C43637 INVX1_LOC_50/A NOR2X1_LOC_570/B 0.09fF
C43638 INVX1_LOC_45/A NAND2X1_LOC_474/Y 0.07fF
C43639 INVX1_LOC_143/Y INVX1_LOC_117/A 0.01fF
C43640 INVX1_LOC_316/Y NOR2X1_LOC_38/B 0.03fF
C43641 INVX1_LOC_239/A NAND2X1_LOC_577/A 0.08fF
C43642 NOR2X1_LOC_106/A NOR2X1_LOC_89/A 0.03fF
C43643 INVX1_LOC_266/A INVX1_LOC_31/A 0.00fF
C43644 NAND2X1_LOC_735/B INVX1_LOC_15/A 0.00fF
C43645 NOR2X1_LOC_324/A INVX1_LOC_9/A 0.00fF
C43646 NOR2X1_LOC_381/Y INVX1_LOC_31/A 0.10fF
C43647 INVX1_LOC_35/A INVX1_LOC_132/A 0.07fF
C43648 INVX1_LOC_313/Y INVX1_LOC_12/A 0.01fF
C43649 INVX1_LOC_46/A NOR2X1_LOC_766/Y 0.03fF
C43650 INVX1_LOC_21/A NOR2X1_LOC_360/Y 0.01fF
C43651 NOR2X1_LOC_6/B INVX1_LOC_23/A 0.07fF
C43652 INVX1_LOC_55/A INVX1_LOC_245/Y 0.01fF
C43653 NOR2X1_LOC_647/A NAND2X1_LOC_819/Y 0.01fF
C43654 NAND2X1_LOC_479/Y NAND2X1_LOC_454/Y 0.02fF
C43655 INVX1_LOC_64/A INVX1_LOC_153/Y 0.01fF
C43656 NOR2X1_LOC_657/a_36_216# NOR2X1_LOC_759/Y 0.00fF
C43657 INVX1_LOC_35/A INVX1_LOC_225/A 0.06fF
C43658 NOR2X1_LOC_810/A NOR2X1_LOC_334/Y 0.10fF
C43659 INVX1_LOC_49/A NOR2X1_LOC_652/Y 0.07fF
C43660 INVX1_LOC_2/A D_INPUT_1 0.47fF
C43661 INVX1_LOC_45/A NAND2X1_LOC_53/Y 0.09fF
C43662 NOR2X1_LOC_33/A NOR2X1_LOC_34/Y 0.01fF
C43663 NOR2X1_LOC_82/A INVX1_LOC_30/A 0.07fF
C43664 NOR2X1_LOC_711/A NAND2X1_LOC_782/B 0.01fF
C43665 INVX1_LOC_14/A NAND2X1_LOC_364/A 0.00fF
C43666 NAND2X1_LOC_654/B NOR2X1_LOC_48/B 0.02fF
C43667 NOR2X1_LOC_497/Y NOR2X1_LOC_754/A 0.03fF
C43668 NOR2X1_LOC_795/Y NOR2X1_LOC_634/Y 0.01fF
C43669 INVX1_LOC_251/Y NAND2X1_LOC_860/A 0.29fF
C43670 INVX1_LOC_223/A INVX1_LOC_161/Y 0.25fF
C43671 NOR2X1_LOC_280/Y INVX1_LOC_185/A 0.00fF
C43672 INVX1_LOC_1/A INVX1_LOC_181/Y 0.01fF
C43673 NAND2X1_LOC_656/Y INVX1_LOC_94/Y 0.11fF
C43674 NOR2X1_LOC_226/A D_INPUT_1 0.07fF
C43675 NAND2X1_LOC_35/Y NAND2X1_LOC_33/Y 0.01fF
C43676 NOR2X1_LOC_848/Y NOR2X1_LOC_68/A 0.02fF
C43677 INVX1_LOC_58/A NOR2X1_LOC_533/A 0.25fF
C43678 INVX1_LOC_36/Y INVX1_LOC_108/A 0.01fF
C43679 INVX1_LOC_206/Y INVX1_LOC_186/Y 0.07fF
C43680 NAND2X1_LOC_787/B NOR2X1_LOC_384/A 0.06fF
C43681 INVX1_LOC_171/A INVX1_LOC_4/Y 0.18fF
C43682 INVX1_LOC_87/Y INVX1_LOC_47/Y 0.03fF
C43683 INVX1_LOC_226/Y INVX1_LOC_224/Y 0.03fF
C43684 INVX1_LOC_64/A INVX1_LOC_177/A 0.03fF
C43685 NAND2X1_LOC_9/Y NOR2X1_LOC_547/B 0.01fF
C43686 INVX1_LOC_35/A NOR2X1_LOC_209/Y 0.04fF
C43687 INVX1_LOC_265/A INVX1_LOC_93/A 0.03fF
C43688 NAND2X1_LOC_9/Y NOR2X1_LOC_78/B 0.15fF
C43689 NOR2X1_LOC_92/Y NOR2X1_LOC_577/Y 0.07fF
C43690 INVX1_LOC_233/A NOR2X1_LOC_78/B 0.07fF
C43691 NOR2X1_LOC_61/Y NOR2X1_LOC_859/Y 0.00fF
C43692 NAND2X1_LOC_551/A NAND2X1_LOC_471/Y 0.02fF
C43693 NOR2X1_LOC_52/a_36_216# NOR2X1_LOC_155/A 0.00fF
C43694 INVX1_LOC_101/A NOR2X1_LOC_383/B 0.00fF
C43695 INVX1_LOC_36/A INVX1_LOC_284/Y 2.53fF
C43696 INVX1_LOC_50/A INVX1_LOC_215/A 0.04fF
C43697 INVX1_LOC_17/A NOR2X1_LOC_13/Y 0.51fF
C43698 INVX1_LOC_118/Y INVX1_LOC_38/A 0.03fF
C43699 INVX1_LOC_64/A INVX1_LOC_280/Y 0.03fF
C43700 NOR2X1_LOC_820/A INPUT_3 0.01fF
C43701 INVX1_LOC_21/A NOR2X1_LOC_792/B 0.01fF
C43702 INVX1_LOC_185/A NAND2X1_LOC_811/B 0.01fF
C43703 INPUT_0 NOR2X1_LOC_861/Y 0.07fF
C43704 NAND2X1_LOC_36/A INVX1_LOC_30/A 0.03fF
C43705 D_INPUT_0 NOR2X1_LOC_318/A 0.09fF
C43706 NAND2X1_LOC_326/A NAND2X1_LOC_325/Y 0.10fF
C43707 NAND2X1_LOC_472/Y NAND2X1_LOC_93/B 0.07fF
C43708 NAND2X1_LOC_53/Y INVX1_LOC_71/A 0.17fF
C43709 NOR2X1_LOC_815/a_36_216# INVX1_LOC_88/A 0.00fF
C43710 NAND2X1_LOC_51/B D_INPUT_5 2.77fF
C43711 NAND2X1_LOC_763/B NAND2X1_LOC_36/A 0.02fF
C43712 NAND2X1_LOC_568/A NOR2X1_LOC_577/Y 0.01fF
C43713 NOR2X1_LOC_369/Y INVX1_LOC_41/Y 0.01fF
C43714 NAND2X1_LOC_553/A NOR2X1_LOC_78/B 0.02fF
C43715 INVX1_LOC_34/A NAND2X1_LOC_67/Y 0.01fF
C43716 NOR2X1_LOC_368/A INVX1_LOC_32/A 0.01fF
C43717 NOR2X1_LOC_241/A INVX1_LOC_49/A 0.15fF
C43718 NOR2X1_LOC_435/B NAND2X1_LOC_453/A 0.03fF
C43719 NOR2X1_LOC_355/A NOR2X1_LOC_383/B 0.07fF
C43720 NOR2X1_LOC_92/Y NOR2X1_LOC_629/B 0.01fF
C43721 NOR2X1_LOC_798/A NOR2X1_LOC_634/B 0.03fF
C43722 NAND2X1_LOC_563/A INVX1_LOC_5/A 0.02fF
C43723 NOR2X1_LOC_679/Y NAND2X1_LOC_567/Y 0.04fF
C43724 NOR2X1_LOC_226/A NOR2X1_LOC_652/Y 0.00fF
C43725 NAND2X1_LOC_35/Y INVX1_LOC_25/Y 0.09fF
C43726 INVX1_LOC_225/Y INVX1_LOC_77/A 0.13fF
C43727 INVX1_LOC_17/A NAND2X1_LOC_175/B 0.09fF
C43728 NOR2X1_LOC_798/A NOR2X1_LOC_78/B 0.03fF
C43729 D_INPUT_3 INVX1_LOC_84/A 0.05fF
C43730 NOR2X1_LOC_454/Y INVX1_LOC_266/Y 0.13fF
C43731 INVX1_LOC_21/A NAND2X1_LOC_451/Y 0.21fF
C43732 NAND2X1_LOC_9/Y NAND2X1_LOC_392/Y 0.00fF
C43733 NAND2X1_LOC_563/Y INVX1_LOC_1/A 0.05fF
C43734 NOR2X1_LOC_572/a_36_216# NOR2X1_LOC_392/Y 0.01fF
C43735 INVX1_LOC_217/A INVX1_LOC_72/A 0.07fF
C43736 INVX1_LOC_14/Y INVX1_LOC_84/A 5.48fF
C43737 NOR2X1_LOC_772/B INVX1_LOC_16/A 0.03fF
C43738 INVX1_LOC_269/A NAND2X1_LOC_562/B 0.04fF
C43739 NOR2X1_LOC_486/Y INVX1_LOC_29/A 0.00fF
C43740 INVX1_LOC_233/A NAND2X1_LOC_392/Y 0.01fF
C43741 NOR2X1_LOC_559/B INVX1_LOC_31/A 0.04fF
C43742 INVX1_LOC_285/Y INVX1_LOC_4/A 0.06fF
C43743 INVX1_LOC_166/A NAND2X1_LOC_622/a_36_24# 0.01fF
C43744 NAND2X1_LOC_638/Y INVX1_LOC_296/A 0.06fF
C43745 NAND2X1_LOC_468/B INVX1_LOC_109/A 0.03fF
C43746 NAND2X1_LOC_538/Y NOR2X1_LOC_52/B 0.19fF
C43747 NAND2X1_LOC_9/Y INVX1_LOC_83/A 0.03fF
C43748 NOR2X1_LOC_769/B INVX1_LOC_89/A 0.02fF
C43749 INVX1_LOC_276/A NAND2X1_LOC_326/A 0.00fF
C43750 INVX1_LOC_49/Y INVX1_LOC_76/A 0.01fF
C43751 INVX1_LOC_13/Y INVX1_LOC_16/A 0.51fF
C43752 INVX1_LOC_299/A NOR2X1_LOC_168/B 2.04fF
C43753 INVX1_LOC_233/Y INVX1_LOC_229/Y 0.10fF
C43754 NOR2X1_LOC_389/A INVX1_LOC_155/A 0.02fF
C43755 NOR2X1_LOC_160/B INVX1_LOC_63/Y 0.07fF
C43756 NAND2X1_LOC_81/B INVX1_LOC_20/A 0.03fF
C43757 NAND2X1_LOC_363/B INVX1_LOC_306/A 0.11fF
C43758 INVX1_LOC_2/Y NAND2X1_LOC_215/a_36_24# 0.00fF
C43759 NOR2X1_LOC_250/A NOR2X1_LOC_52/B 0.95fF
C43760 D_INPUT_1 INPUT_1 0.45fF
C43761 NOR2X1_LOC_598/B INVX1_LOC_89/A 0.78fF
C43762 NAND2X1_LOC_181/a_36_24# NOR2X1_LOC_791/Y 0.01fF
C43763 INPUT_3 INVX1_LOC_315/A 0.20fF
C43764 INVX1_LOC_11/A NOR2X1_LOC_709/A 0.13fF
C43765 NAND2X1_LOC_84/Y NAND2X1_LOC_364/A 0.07fF
C43766 INVX1_LOC_51/A INVX1_LOC_89/A 0.00fF
C43767 NAND2X1_LOC_212/Y NAND2X1_LOC_220/B 0.00fF
C43768 NOR2X1_LOC_788/B INVX1_LOC_58/Y 0.01fF
C43769 NOR2X1_LOC_361/B NAND2X1_LOC_850/Y 0.29fF
C43770 INVX1_LOC_27/A INVX1_LOC_137/Y 0.11fF
C43771 INVX1_LOC_269/A NOR2X1_LOC_773/Y 0.03fF
C43772 NAND2X1_LOC_842/B INVX1_LOC_53/A 0.23fF
C43773 NOR2X1_LOC_312/Y NOR2X1_LOC_109/Y 0.10fF
C43774 NOR2X1_LOC_598/B NAND2X1_LOC_508/A 0.07fF
C43775 NAND2X1_LOC_711/Y NAND2X1_LOC_308/Y 0.00fF
C43776 INVX1_LOC_72/A NAND2X1_LOC_787/B 0.70fF
C43777 INVX1_LOC_31/A NOR2X1_LOC_6/B 0.18fF
C43778 NOR2X1_LOC_92/Y INVX1_LOC_22/A 0.78fF
C43779 NAND2X1_LOC_332/Y INVX1_LOC_30/A 0.01fF
C43780 NOR2X1_LOC_160/B NOR2X1_LOC_175/A 0.00fF
C43781 NAND2X1_LOC_391/Y INVX1_LOC_234/A 0.00fF
C43782 INVX1_LOC_146/A INVX1_LOC_53/A 0.17fF
C43783 INVX1_LOC_36/A NOR2X1_LOC_561/a_36_216# 0.00fF
C43784 INVX1_LOC_2/A NOR2X1_LOC_371/a_36_216# 0.01fF
C43785 INVX1_LOC_113/A INVX1_LOC_117/Y 0.06fF
C43786 INVX1_LOC_5/A NOR2X1_LOC_814/Y 0.21fF
C43787 INVX1_LOC_38/A NOR2X1_LOC_258/Y 0.02fF
C43788 INVX1_LOC_5/A NOR2X1_LOC_214/B 0.20fF
C43789 NOR2X1_LOC_798/A INVX1_LOC_83/A 0.03fF
C43790 NAND2X1_LOC_195/Y INVX1_LOC_63/Y 0.01fF
C43791 INVX1_LOC_260/Y INVX1_LOC_260/A 0.09fF
C43792 INVX1_LOC_88/A INVX1_LOC_16/A 0.07fF
C43793 NAND2X1_LOC_60/a_36_24# NOR2X1_LOC_243/B 0.00fF
C43794 NOR2X1_LOC_428/Y NAND2X1_LOC_451/Y 0.11fF
C43795 INVX1_LOC_6/A NOR2X1_LOC_72/Y 0.02fF
C43796 NAND2X1_LOC_858/B INVX1_LOC_57/A 0.68fF
C43797 INVX1_LOC_115/A NOR2X1_LOC_467/A 0.04fF
C43798 NOR2X1_LOC_552/Y NOR2X1_LOC_383/B 0.00fF
C43799 INVX1_LOC_226/Y NOR2X1_LOC_103/Y 0.01fF
C43800 INVX1_LOC_119/Y INVX1_LOC_92/A 0.15fF
C43801 NOR2X1_LOC_541/Y NOR2X1_LOC_500/Y 0.01fF
C43802 INPUT_1 NOR2X1_LOC_652/Y 0.00fF
C43803 INVX1_LOC_187/A INVX1_LOC_78/A 0.00fF
C43804 INVX1_LOC_104/A INVX1_LOC_18/A 0.14fF
C43805 NAND2X1_LOC_267/B INVX1_LOC_4/A 0.03fF
C43806 INVX1_LOC_14/Y INVX1_LOC_15/A 0.01fF
C43807 INVX1_LOC_20/A INVX1_LOC_4/Y 0.07fF
C43808 NOR2X1_LOC_790/B NOR2X1_LOC_569/A 0.07fF
C43809 INVX1_LOC_13/Y INVX1_LOC_28/A 0.04fF
C43810 NOR2X1_LOC_351/Y INVX1_LOC_29/A 0.07fF
C43811 NOR2X1_LOC_406/a_36_216# NOR2X1_LOC_322/Y 0.02fF
C43812 INVX1_LOC_124/Y NOR2X1_LOC_191/A 0.04fF
C43813 NAND2X1_LOC_276/Y INVX1_LOC_314/Y 0.01fF
C43814 NAND2X1_LOC_218/B INVX1_LOC_201/Y 0.64fF
C43815 NAND2X1_LOC_93/B NAND2X1_LOC_773/B 0.01fF
C43816 INVX1_LOC_269/A NOR2X1_LOC_332/A 1.39fF
C43817 NAND2X1_LOC_854/B NAND2X1_LOC_799/A 0.24fF
C43818 INVX1_LOC_12/A NOR2X1_LOC_506/Y 0.12fF
C43819 NOR2X1_LOC_598/B NOR2X1_LOC_703/Y 0.10fF
C43820 INVX1_LOC_271/A INVX1_LOC_91/A 0.03fF
C43821 INVX1_LOC_230/Y INVX1_LOC_13/A 0.09fF
C43822 INVX1_LOC_278/Y INVX1_LOC_30/A 0.12fF
C43823 INVX1_LOC_64/A INVX1_LOC_285/Y 0.54fF
C43824 NAND2X1_LOC_350/A NAND2X1_LOC_319/A 0.14fF
C43825 INVX1_LOC_45/A NOR2X1_LOC_500/Y 0.06fF
C43826 INVX1_LOC_117/A NOR2X1_LOC_835/a_36_216# 0.00fF
C43827 INVX1_LOC_45/A INVX1_LOC_226/Y 0.72fF
C43828 NOR2X1_LOC_629/Y INVX1_LOC_42/A 0.03fF
C43829 NOR2X1_LOC_455/a_36_216# NOR2X1_LOC_577/Y 0.00fF
C43830 INVX1_LOC_102/Y NAND2X1_LOC_474/Y 0.11fF
C43831 INVX1_LOC_30/Y INVX1_LOC_31/A 0.15fF
C43832 NOR2X1_LOC_255/a_36_216# INVX1_LOC_61/Y 0.00fF
C43833 INVX1_LOC_33/A INVX1_LOC_8/A 0.07fF
C43834 INVX1_LOC_3/A NAND2X1_LOC_206/Y 0.17fF
C43835 NAND2X1_LOC_763/B NAND2X1_LOC_59/a_36_24# 0.00fF
C43836 NAND2X1_LOC_860/A NOR2X1_LOC_45/B 0.07fF
C43837 INVX1_LOC_230/A INVX1_LOC_15/A 0.17fF
C43838 NOR2X1_LOC_755/Y INVX1_LOC_92/A 0.02fF
C43839 INVX1_LOC_268/A NOR2X1_LOC_657/Y 0.00fF
C43840 INVX1_LOC_27/A INVX1_LOC_79/A 0.01fF
C43841 INVX1_LOC_77/A INVX1_LOC_266/Y 0.07fF
C43842 NOR2X1_LOC_577/Y NAND2X1_LOC_477/A 0.10fF
C43843 NOR2X1_LOC_276/Y NOR2X1_LOC_366/Y 0.21fF
C43844 INVX1_LOC_25/A NOR2X1_LOC_675/A -0.00fF
C43845 INVX1_LOC_136/A INVX1_LOC_232/A 0.16fF
C43846 NOR2X1_LOC_124/A INVX1_LOC_23/A 0.02fF
C43847 INVX1_LOC_88/A INVX1_LOC_28/A 0.18fF
C43848 INVX1_LOC_3/A NAND2X1_LOC_773/B 0.08fF
C43849 NAND2X1_LOC_341/A NOR2X1_LOC_759/A 0.27fF
C43850 INVX1_LOC_10/Y NAND2X1_LOC_454/Y 0.03fF
C43851 INVX1_LOC_34/A NOR2X1_LOC_367/B 0.13fF
C43852 NOR2X1_LOC_180/Y NOR2X1_LOC_254/Y 0.03fF
C43853 NOR2X1_LOC_593/Y NOR2X1_LOC_709/A 0.01fF
C43854 NOR2X1_LOC_68/A NAND2X1_LOC_479/Y 0.03fF
C43855 NOR2X1_LOC_458/B NOR2X1_LOC_303/Y 0.08fF
C43856 INVX1_LOC_45/A INVX1_LOC_10/A 0.56fF
C43857 VDD NOR2X1_LOC_720/A -0.00fF
C43858 NOR2X1_LOC_67/A NOR2X1_LOC_625/Y 0.02fF
C43859 NOR2X1_LOC_554/B NAND2X1_LOC_41/Y 0.02fF
C43860 INVX1_LOC_35/A NAND2X1_LOC_642/Y 0.03fF
C43861 INVX1_LOC_64/A INVX1_LOC_65/A 0.01fF
C43862 INVX1_LOC_37/Y NOR2X1_LOC_693/Y 0.01fF
C43863 NOR2X1_LOC_103/a_36_216# NAND2X1_LOC_254/Y 0.00fF
C43864 NOR2X1_LOC_620/B INVX1_LOC_49/A 0.01fF
C43865 NAND2X1_LOC_856/A INVX1_LOC_10/A 0.03fF
C43866 NOR2X1_LOC_500/Y INVX1_LOC_71/A 0.07fF
C43867 NAND2X1_LOC_214/B INVX1_LOC_91/A 0.02fF
C43868 INVX1_LOC_226/Y INVX1_LOC_71/A 0.16fF
C43869 INVX1_LOC_39/A INVX1_LOC_123/A -0.02fF
C43870 INVX1_LOC_36/A NAND2X1_LOC_779/a_36_24# 0.01fF
C43871 INVX1_LOC_22/A NAND2X1_LOC_837/Y 0.14fF
C43872 NOR2X1_LOC_92/Y INVX1_LOC_100/A 0.03fF
C43873 INVX1_LOC_36/A NOR2X1_LOC_525/Y 0.09fF
C43874 INVX1_LOC_279/Y NOR2X1_LOC_828/A 0.06fF
C43875 NAND2X1_LOC_574/A GATE_222 0.07fF
C43876 INVX1_LOC_36/A NAND2X1_LOC_809/A 0.01fF
C43877 VDD INVX1_LOC_129/A -0.00fF
C43878 INVX1_LOC_36/A NOR2X1_LOC_312/Y 0.08fF
C43879 INVX1_LOC_136/A NAND2X1_LOC_523/a_36_24# 0.01fF
C43880 NOR2X1_LOC_753/Y NOR2X1_LOC_165/Y 0.05fF
C43881 NOR2X1_LOC_52/B NOR2X1_LOC_709/A 0.07fF
C43882 NAND2X1_LOC_350/B INVX1_LOC_63/Y 0.03fF
C43883 NOR2X1_LOC_590/A INVX1_LOC_148/A 0.01fF
C43884 INVX1_LOC_305/A D_INPUT_0 0.09fF
C43885 INVX1_LOC_27/A INVX1_LOC_91/A 0.30fF
C43886 INVX1_LOC_274/A INVX1_LOC_271/Y -0.01fF
C43887 NOR2X1_LOC_261/Y INVX1_LOC_14/Y 1.03fF
C43888 NAND2X1_LOC_363/B INVX1_LOC_176/A 0.05fF
C43889 INVX1_LOC_233/Y INVX1_LOC_20/A 0.08fF
C43890 NOR2X1_LOC_607/A INVX1_LOC_227/A 0.01fF
C43891 INVX1_LOC_2/A NOR2X1_LOC_591/Y 0.34fF
C43892 NOR2X1_LOC_824/A INVX1_LOC_91/A 0.38fF
C43893 INVX1_LOC_135/A NOR2X1_LOC_68/A 8.37fF
C43894 NAND2X1_LOC_9/Y INVX1_LOC_46/A 0.00fF
C43895 INPUT_6 VDD 0.83fF
C43896 NAND2X1_LOC_364/A NOR2X1_LOC_137/A 0.04fF
C43897 INVX1_LOC_208/A INVX1_LOC_63/Y 0.10fF
C43898 NOR2X1_LOC_203/a_36_216# NAND2X1_LOC_447/Y 0.12fF
C43899 NAND2X1_LOC_9/Y NOR2X1_LOC_98/A 0.01fF
C43900 INVX1_LOC_95/Y INVX1_LOC_306/Y 0.19fF
C43901 INVX1_LOC_233/A INVX1_LOC_46/A 0.07fF
C43902 INVX1_LOC_57/A NOR2X1_LOC_98/B 0.02fF
C43903 INVX1_LOC_40/A INVX1_LOC_8/A 0.04fF
C43904 INVX1_LOC_10/A INVX1_LOC_71/A 0.12fF
C43905 INVX1_LOC_41/A INVX1_LOC_22/A 0.05fF
C43906 INVX1_LOC_47/Y INVX1_LOC_285/A 0.00fF
C43907 INVX1_LOC_150/Y NOR2X1_LOC_113/B 0.05fF
C43908 NOR2X1_LOC_445/a_36_216# NOR2X1_LOC_74/A 0.01fF
C43909 NOR2X1_LOC_498/Y INVX1_LOC_22/A 0.00fF
C43910 NAND2X1_LOC_624/B VDD 0.17fF
C43911 NOR2X1_LOC_68/A NOR2X1_LOC_560/A 0.00fF
C43912 INVX1_LOC_34/A NOR2X1_LOC_719/A 0.19fF
C43913 NOR2X1_LOC_78/B NOR2X1_LOC_718/a_36_216# 0.00fF
C43914 NOR2X1_LOC_388/Y NOR2X1_LOC_570/Y 0.04fF
C43915 NOR2X1_LOC_211/Y VDD 0.24fF
C43916 NOR2X1_LOC_824/A INVX1_LOC_11/Y 0.17fF
C43917 NAND2X1_LOC_570/Y NAND2X1_LOC_578/B 0.04fF
C43918 NOR2X1_LOC_234/Y INVX1_LOC_25/Y 0.03fF
C43919 INVX1_LOC_135/A NOR2X1_LOC_204/a_36_216# 0.01fF
C43920 INVX1_LOC_47/Y NOR2X1_LOC_814/A 0.20fF
C43921 NAND2X1_LOC_537/Y NOR2X1_LOC_45/B 0.07fF
C43922 NAND2X1_LOC_21/Y INPUT_5 0.19fF
C43923 NOR2X1_LOC_860/B NAND2X1_LOC_45/Y 0.22fF
C43924 INVX1_LOC_278/Y NAND2X1_LOC_722/A 0.02fF
C43925 NOR2X1_LOC_414/a_36_216# NAND2X1_LOC_348/A 0.00fF
C43926 INVX1_LOC_50/A INVX1_LOC_54/A 8.76fF
C43927 INVX1_LOC_34/A NOR2X1_LOC_561/Y 3.00fF
C43928 INVX1_LOC_14/A NOR2X1_LOC_405/A 0.02fF
C43929 INVX1_LOC_1/A NOR2X1_LOC_675/A -0.00fF
C43930 VDD NOR2X1_LOC_849/A 0.29fF
C43931 D_INPUT_2 INPUT_1 1.09fF
C43932 INVX1_LOC_34/A INVX1_LOC_7/A 1.91fF
C43933 NAND2X1_LOC_721/B NOR2X1_LOC_323/Y 0.18fF
C43934 D_INPUT_1 INVX1_LOC_118/A 0.60fF
C43935 INVX1_LOC_5/A INVX1_LOC_12/Y 0.00fF
C43936 NAND2X1_LOC_287/a_36_24# NOR2X1_LOC_743/Y 0.00fF
C43937 NOR2X1_LOC_200/a_36_216# INVX1_LOC_290/A 0.01fF
C43938 NOR2X1_LOC_140/A INVX1_LOC_74/A 0.01fF
C43939 INVX1_LOC_33/A NAND2X1_LOC_140/A 0.00fF
C43940 VDD NOR2X1_LOC_852/Y 0.51fF
C43941 NAND2X1_LOC_471/Y NAND2X1_LOC_489/Y 0.01fF
C43942 VDD NOR2X1_LOC_440/B 0.02fF
C43943 INVX1_LOC_71/A NOR2X1_LOC_302/Y 0.08fF
C43944 NOR2X1_LOC_175/B NOR2X1_LOC_211/A 0.19fF
C43945 NAND2X1_LOC_181/Y INVX1_LOC_56/Y 0.00fF
C43946 NOR2X1_LOC_224/Y INVX1_LOC_54/A 0.01fF
C43947 NOR2X1_LOC_180/B NOR2X1_LOC_344/A 0.02fF
C43948 NOR2X1_LOC_380/A GATE_811 0.00fF
C43949 INVX1_LOC_75/A INVX1_LOC_94/A 0.13fF
C43950 NAND2X1_LOC_79/Y NAND2X1_LOC_348/A 0.01fF
C43951 NOR2X1_LOC_312/Y NOR2X1_LOC_309/Y 0.04fF
C43952 NOR2X1_LOC_278/Y INVX1_LOC_63/A 0.07fF
C43953 NAND2X1_LOC_231/Y NOR2X1_LOC_561/Y 0.10fF
C43954 NOR2X1_LOC_68/A NOR2X1_LOC_391/B 0.01fF
C43955 NOR2X1_LOC_778/B NOR2X1_LOC_553/B 0.01fF
C43956 NAND2X1_LOC_349/B NOR2X1_LOC_136/Y 0.03fF
C43957 NOR2X1_LOC_604/Y INVX1_LOC_92/A 0.03fF
C43958 NOR2X1_LOC_52/B NOR2X1_LOC_106/A 0.32fF
C43959 NOR2X1_LOC_211/A INVX1_LOC_22/A 0.15fF
C43960 NOR2X1_LOC_780/B INVX1_LOC_117/A 0.01fF
C43961 INVX1_LOC_276/A NAND2X1_LOC_683/a_36_24# 0.01fF
C43962 INVX1_LOC_174/A INVX1_LOC_115/Y 0.02fF
C43963 NOR2X1_LOC_68/A NOR2X1_LOC_794/A 0.02fF
C43964 NOR2X1_LOC_171/Y NAND2X1_LOC_175/B 0.00fF
C43965 NOR2X1_LOC_289/Y NOR2X1_LOC_172/Y 0.01fF
C43966 NAND2X1_LOC_599/a_36_24# INVX1_LOC_307/A 0.00fF
C43967 INVX1_LOC_118/A NOR2X1_LOC_652/Y 0.08fF
C43968 NOR2X1_LOC_89/A NOR2X1_LOC_334/Y 0.14fF
C43969 NOR2X1_LOC_695/Y NAND2X1_LOC_712/A 0.09fF
C43970 INVX1_LOC_310/A INVX1_LOC_132/Y 0.02fF
C43971 NOR2X1_LOC_354/B INVX1_LOC_160/A 0.74fF
C43972 NOR2X1_LOC_75/Y NAND2X1_LOC_39/Y 0.01fF
C43973 NAND2X1_LOC_563/A NOR2X1_LOC_332/A 0.10fF
C43974 INVX1_LOC_45/A NOR2X1_LOC_799/B 0.01fF
C43975 NAND2X1_LOC_656/Y NOR2X1_LOC_321/a_36_216# 0.00fF
C43976 NOR2X1_LOC_45/B NAND2X1_LOC_640/a_36_24# 0.01fF
C43977 NOR2X1_LOC_372/A NAND2X1_LOC_244/A 0.03fF
C43978 INVX1_LOC_53/A INVX1_LOC_119/Y 0.02fF
C43979 NOR2X1_LOC_32/a_36_216# NOR2X1_LOC_32/Y 0.03fF
C43980 NOR2X1_LOC_799/B NOR2X1_LOC_568/A 0.04fF
C43981 NOR2X1_LOC_68/A NOR2X1_LOC_552/A 0.10fF
C43982 NAND2X1_LOC_534/a_36_24# INVX1_LOC_28/A 0.00fF
C43983 INVX1_LOC_196/A NOR2X1_LOC_356/A 0.10fF
C43984 NAND2X1_LOC_208/B INVX1_LOC_76/A 0.01fF
C43985 INVX1_LOC_86/Y NOR2X1_LOC_713/B 0.19fF
C43986 NOR2X1_LOC_299/Y INVX1_LOC_22/A 0.06fF
C43987 NOR2X1_LOC_421/a_36_216# INVX1_LOC_12/A 0.00fF
C43988 INVX1_LOC_256/A NAND2X1_LOC_472/Y 0.10fF
C43989 INVX1_LOC_29/A NOR2X1_LOC_635/B 0.03fF
C43990 NOR2X1_LOC_78/B NAND2X1_LOC_842/B 0.07fF
C43991 INVX1_LOC_41/A INVX1_LOC_100/A 0.05fF
C43992 NOR2X1_LOC_718/Y INVX1_LOC_6/A 0.06fF
C43993 INVX1_LOC_136/A NAND2X1_LOC_447/Y 0.10fF
C43994 INVX1_LOC_77/A INVX1_LOC_125/Y 0.07fF
C43995 NOR2X1_LOC_514/A VDD 0.02fF
C43996 INVX1_LOC_202/A NOR2X1_LOC_78/A 0.07fF
C43997 INVX1_LOC_29/A NOR2X1_LOC_748/A 0.03fF
C43998 NAND2X1_LOC_578/B NOR2X1_LOC_19/B 0.10fF
C43999 INVX1_LOC_4/A INVX1_LOC_4/Y 4.70fF
C44000 NOR2X1_LOC_324/A NOR2X1_LOC_324/Y 0.01fF
C44001 INVX1_LOC_224/Y INVX1_LOC_12/A 0.03fF
C44002 NOR2X1_LOC_89/A NAND2X1_LOC_464/B 0.12fF
C44003 INVX1_LOC_36/A NAND2X1_LOC_287/B 0.15fF
C44004 NOR2X1_LOC_789/a_36_216# NOR2X1_LOC_99/B 0.01fF
C44005 NOR2X1_LOC_92/Y NOR2X1_LOC_88/A 0.03fF
C44006 INVX1_LOC_142/A VDD 0.42fF
C44007 NAND2X1_LOC_832/Y INVX1_LOC_266/Y 0.01fF
C44008 NOR2X1_LOC_6/B INVX1_LOC_6/A 0.04fF
C44009 NAND2X1_LOC_51/B NAND2X1_LOC_451/Y 0.11fF
C44010 NOR2X1_LOC_123/B INVX1_LOC_10/A 0.01fF
C44011 INVX1_LOC_35/A NOR2X1_LOC_48/Y 0.08fF
C44012 NAND2X1_LOC_149/Y INVX1_LOC_107/Y 0.00fF
C44013 NOR2X1_LOC_641/B NAND2X1_LOC_230/a_36_24# 0.00fF
C44014 NOR2X1_LOC_410/Y VDD 0.24fF
C44015 INVX1_LOC_225/Y INVX1_LOC_9/A 0.08fF
C44016 INVX1_LOC_50/A NOR2X1_LOC_48/B 0.34fF
C44017 INVX1_LOC_27/A NOR2X1_LOC_179/Y 0.01fF
C44018 INVX1_LOC_280/Y INVX1_LOC_282/A 0.07fF
C44019 NAND2X1_LOC_227/Y INVX1_LOC_54/A 0.00fF
C44020 NOR2X1_LOC_617/Y NAND2X1_LOC_659/B 0.01fF
C44021 NOR2X1_LOC_272/Y NOR2X1_LOC_127/Y 0.10fF
C44022 INVX1_LOC_64/A NAND2X1_LOC_81/B 0.00fF
C44023 INVX1_LOC_200/A NAND2X1_LOC_444/a_36_24# 0.00fF
C44024 NAND2X1_LOC_391/Y NAND2X1_LOC_477/Y 0.10fF
C44025 INVX1_LOC_197/Y NOR2X1_LOC_19/Y 0.01fF
C44026 NOR2X1_LOC_332/A NOR2X1_LOC_814/Y 0.03fF
C44027 INVX1_LOC_303/A NOR2X1_LOC_35/Y 0.10fF
C44028 INVX1_LOC_41/Y VDD 0.41fF
C44029 NOR2X1_LOC_576/B NOR2X1_LOC_576/a_36_216# 0.00fF
C44030 NOR2X1_LOC_824/A INVX1_LOC_203/A 0.03fF
C44031 INVX1_LOC_32/A NAND2X1_LOC_201/a_36_24# 0.00fF
C44032 NAND2X1_LOC_803/B NAND2X1_LOC_798/B 0.03fF
C44033 NAND2X1_LOC_866/A INVX1_LOC_46/A 0.02fF
C44034 NOR2X1_LOC_617/Y VDD 0.77fF
C44035 INPUT_3 NOR2X1_LOC_660/a_36_216# 0.00fF
C44036 INVX1_LOC_206/A INVX1_LOC_91/A 0.29fF
C44037 INVX1_LOC_2/A NOR2X1_LOC_144/a_36_216# 0.02fF
C44038 NAND2X1_LOC_357/B NAND2X1_LOC_729/B 0.02fF
C44039 NAND2X1_LOC_63/Y NOR2X1_LOC_652/Y 0.00fF
C44040 NAND2X1_LOC_593/Y VDD 0.51fF
C44041 INVX1_LOC_57/A NOR2X1_LOC_38/B 0.14fF
C44042 INVX1_LOC_295/A NOR2X1_LOC_163/A 0.10fF
C44043 INVX1_LOC_45/Y NOR2X1_LOC_363/Y 0.04fF
C44044 INVX1_LOC_90/A INVX1_LOC_65/Y 0.00fF
C44045 INVX1_LOC_10/A INVX1_LOC_102/Y 0.05fF
C44046 INVX1_LOC_17/A NOR2X1_LOC_697/Y 0.05fF
C44047 INVX1_LOC_286/Y INVX1_LOC_185/A 0.20fF
C44048 NOR2X1_LOC_634/B NOR2X1_LOC_334/a_36_216# 0.00fF
C44049 NOR2X1_LOC_68/A INVX1_LOC_280/A 0.53fF
C44050 INVX1_LOC_47/Y NOR2X1_LOC_292/a_36_216# 0.01fF
C44051 NOR2X1_LOC_454/Y INVX1_LOC_19/A 0.07fF
C44052 NOR2X1_LOC_590/A NAND2X1_LOC_798/B 0.07fF
C44053 INVX1_LOC_34/A INVX1_LOC_76/A 0.64fF
C44054 INVX1_LOC_135/A NAND2X1_LOC_462/a_36_24# 0.00fF
C44055 INVX1_LOC_103/A NAND2X1_LOC_475/Y 0.00fF
C44056 INVX1_LOC_111/Y NOR2X1_LOC_405/A 0.05fF
C44057 INVX1_LOC_24/A NOR2X1_LOC_536/A 0.23fF
C44058 INVX1_LOC_63/Y NAND2X1_LOC_211/Y 0.08fF
C44059 NOR2X1_LOC_561/Y INPUT_0 0.01fF
C44060 NOR2X1_LOC_758/Y VDD 0.40fF
C44061 INVX1_LOC_30/Y INVX1_LOC_6/A 0.03fF
C44062 INVX1_LOC_45/A INVX1_LOC_307/A 0.07fF
C44063 NOR2X1_LOC_251/Y INVX1_LOC_91/A 0.04fF
C44064 NOR2X1_LOC_204/a_36_216# INVX1_LOC_280/A 0.01fF
C44065 NOR2X1_LOC_309/Y NAND2X1_LOC_287/B 0.02fF
C44066 INVX1_LOC_72/A INVX1_LOC_92/A 0.15fF
C44067 NAND2X1_LOC_812/A NOR2X1_LOC_766/Y 0.00fF
C44068 INVX1_LOC_45/A NOR2X1_LOC_445/B 0.07fF
C44069 INVX1_LOC_292/A NAND2X1_LOC_475/Y 0.03fF
C44070 NOR2X1_LOC_768/a_36_216# INVX1_LOC_75/A 0.00fF
C44071 NOR2X1_LOC_403/B INVX1_LOC_118/A 0.01fF
C44072 NOR2X1_LOC_568/A NOR2X1_LOC_445/B 0.00fF
C44073 NAND2X1_LOC_589/a_36_24# NAND2X1_LOC_798/B 0.00fF
C44074 NOR2X1_LOC_557/Y NOR2X1_LOC_536/A 0.03fF
C44075 NAND2X1_LOC_231/Y INVX1_LOC_76/A 0.10fF
C44076 INVX1_LOC_88/A INVX1_LOC_109/A 0.01fF
C44077 INVX1_LOC_290/A NOR2X1_LOC_139/Y 0.05fF
C44078 NOR2X1_LOC_231/B NOR2X1_LOC_814/A 0.03fF
C44079 INVX1_LOC_198/Y INVX1_LOC_92/A 0.01fF
C44080 INVX1_LOC_24/A NAND2X1_LOC_93/B 0.03fF
C44081 NAND2X1_LOC_622/B NAND2X1_LOC_624/A 0.01fF
C44082 NOR2X1_LOC_750/A NAND2X1_LOC_348/A 0.01fF
C44083 INVX1_LOC_269/A NOR2X1_LOC_847/A 0.01fF
C44084 INVX1_LOC_105/A INVX1_LOC_54/A 0.00fF
C44085 VDD NOR2X1_LOC_538/Y 0.24fF
C44086 NOR2X1_LOC_526/Y INVX1_LOC_20/A 0.62fF
C44087 NOR2X1_LOC_122/A INVX1_LOC_290/Y 0.02fF
C44088 INVX1_LOC_33/A INVX1_LOC_118/Y 0.03fF
C44089 INVX1_LOC_308/Y NOR2X1_LOC_89/A 0.04fF
C44090 NAND2X1_LOC_837/Y NOR2X1_LOC_88/A 0.11fF
C44091 NOR2X1_LOC_103/Y INVX1_LOC_12/A 0.07fF
C44092 INVX1_LOC_269/A INVX1_LOC_42/A 0.11fF
C44093 INVX1_LOC_234/A INVX1_LOC_91/A 0.03fF
C44094 INVX1_LOC_47/A NOR2X1_LOC_9/Y 0.23fF
C44095 NOR2X1_LOC_750/a_36_216# NAND2X1_LOC_348/A 0.00fF
C44096 NOR2X1_LOC_191/A NOR2X1_LOC_266/B 0.03fF
C44097 INVX1_LOC_71/A INVX1_LOC_307/A 0.07fF
C44098 NOR2X1_LOC_505/Y INVX1_LOC_46/A 0.14fF
C44099 INVX1_LOC_24/A NAND2X1_LOC_425/Y 0.01fF
C44100 INVX1_LOC_290/A NAND2X1_LOC_468/B 0.02fF
C44101 NOR2X1_LOC_538/a_36_216# INVX1_LOC_22/A 0.00fF
C44102 NOR2X1_LOC_606/Y NAND2X1_LOC_773/B 0.01fF
C44103 NAND2X1_LOC_699/a_36_24# NOR2X1_LOC_709/A 0.02fF
C44104 INVX1_LOC_71/A NOR2X1_LOC_445/B 0.10fF
C44105 NAND2X1_LOC_341/A NOR2X1_LOC_357/Y 0.09fF
C44106 NOR2X1_LOC_773/Y INVX1_LOC_12/Y 0.10fF
C44107 NAND2X1_LOC_577/A NAND2X1_LOC_82/Y 0.08fF
C44108 NOR2X1_LOC_574/a_36_216# INVX1_LOC_38/A 0.01fF
C44109 NOR2X1_LOC_557/Y NAND2X1_LOC_93/B 0.07fF
C44110 NOR2X1_LOC_210/B INVX1_LOC_37/A 0.04fF
C44111 NOR2X1_LOC_19/B INVX1_LOC_309/A 0.03fF
C44112 NAND2X1_LOC_218/B NAND2X1_LOC_574/A -0.07fF
C44113 NOR2X1_LOC_137/A NOR2X1_LOC_405/A 0.04fF
C44114 INVX1_LOC_255/Y INVX1_LOC_2/Y 0.00fF
C44115 INVX1_LOC_143/A NOR2X1_LOC_536/A 0.03fF
C44116 INVX1_LOC_83/A NOR2X1_LOC_545/B 0.02fF
C44117 INVX1_LOC_266/Y INVX1_LOC_9/A 0.02fF
C44118 INVX1_LOC_24/A INVX1_LOC_3/A 0.61fF
C44119 NAND2X1_LOC_850/A INVX1_LOC_100/Y 0.01fF
C44120 NOR2X1_LOC_205/Y INVX1_LOC_4/A 0.00fF
C44121 INVX1_LOC_90/A NOR2X1_LOC_746/Y 0.02fF
C44122 INVX1_LOC_21/A INVX1_LOC_26/A 0.03fF
C44123 NOR2X1_LOC_91/A NAND2X1_LOC_778/Y 0.01fF
C44124 INVX1_LOC_45/A INVX1_LOC_12/A 0.25fF
C44125 NOR2X1_LOC_160/B NOR2X1_LOC_462/a_36_216# 0.02fF
C44126 NOR2X1_LOC_690/A NOR2X1_LOC_88/Y 1.99fF
C44127 NAND2X1_LOC_9/Y INVX1_LOC_233/A 0.03fF
C44128 NAND2X1_LOC_749/a_36_24# NAND2X1_LOC_215/A 0.01fF
C44129 INPUT_0 NOR2X1_LOC_167/Y 0.08fF
C44130 NOR2X1_LOC_264/a_36_216# INVX1_LOC_78/A 0.01fF
C44131 NAND2X1_LOC_856/A INVX1_LOC_12/A 0.03fF
C44132 INVX1_LOC_174/A D_INPUT_5 0.09fF
C44133 INVX1_LOC_269/A INVX1_LOC_78/A 0.07fF
C44134 NOR2X1_LOC_420/Y INVX1_LOC_57/A 0.00fF
C44135 INVX1_LOC_230/Y INVX1_LOC_32/A 1.18fF
C44136 NAND2X1_LOC_565/B NOR2X1_LOC_536/A 0.00fF
C44137 NOR2X1_LOC_700/Y INVX1_LOC_46/A 0.25fF
C44138 NAND2X1_LOC_7/Y INVX1_LOC_63/A 0.01fF
C44139 INVX1_LOC_43/Y NAND2X1_LOC_269/a_36_24# 0.00fF
C44140 INVX1_LOC_11/A NOR2X1_LOC_334/Y 0.38fF
C44141 NOR2X1_LOC_392/B INVX1_LOC_123/Y 0.22fF
C44142 INVX1_LOC_233/Y INVX1_LOC_64/A 0.07fF
C44143 NAND2X1_LOC_9/Y NAND2X1_LOC_553/A 0.02fF
C44144 INVX1_LOC_143/A NAND2X1_LOC_93/B 0.07fF
C44145 INVX1_LOC_256/Y NOR2X1_LOC_118/a_36_216# 0.00fF
C44146 NOR2X1_LOC_690/A INVX1_LOC_84/A 0.03fF
C44147 NOR2X1_LOC_537/Y INVX1_LOC_92/A 0.07fF
C44148 NOR2X1_LOC_91/A NOR2X1_LOC_15/Y 5.20fF
C44149 INVX1_LOC_39/A D_INPUT_1 0.05fF
C44150 INVX1_LOC_53/A NOR2X1_LOC_674/Y 0.03fF
C44151 INVX1_LOC_77/A INVX1_LOC_19/A 14.25fF
C44152 INVX1_LOC_314/Y INVX1_LOC_125/A 0.04fF
C44153 NOR2X1_LOC_411/A NOR2X1_LOC_411/Y 0.12fF
C44154 NOR2X1_LOC_71/Y INVX1_LOC_37/Y 0.24fF
C44155 NOR2X1_LOC_5/a_36_216# D_INPUT_3 0.00fF
C44156 NOR2X1_LOC_65/B INVX1_LOC_269/A 0.10fF
C44157 INVX1_LOC_71/A INVX1_LOC_12/A 0.14fF
C44158 NAND2X1_LOC_783/A NOR2X1_LOC_536/A 0.03fF
C44159 INVX1_LOC_41/A INVX1_LOC_186/Y 0.04fF
C44160 NAND2X1_LOC_842/B INVX1_LOC_46/A 0.03fF
C44161 INVX1_LOC_200/Y NAND2X1_LOC_579/A 0.03fF
C44162 NOR2X1_LOC_815/a_36_216# INVX1_LOC_272/A 0.01fF
C44163 NOR2X1_LOC_468/Y INVX1_LOC_57/A 0.13fF
C44164 INVX1_LOC_10/A NOR2X1_LOC_331/B 0.21fF
C44165 NOR2X1_LOC_130/A NOR2X1_LOC_536/A 0.10fF
C44166 INVX1_LOC_31/A INVX1_LOC_273/A 1.32fF
C44167 INVX1_LOC_16/A NOR2X1_LOC_99/Y 0.03fF
C44168 INVX1_LOC_95/Y NOR2X1_LOC_74/A 0.22fF
C44169 NOR2X1_LOC_15/Y INVX1_LOC_23/A 5.79fF
C44170 NOR2X1_LOC_437/Y INVX1_LOC_290/Y 0.04fF
C44171 NOR2X1_LOC_732/A INVX1_LOC_19/A 0.03fF
C44172 NAND2X1_LOC_571/B NAND2X1_LOC_579/A 0.03fF
C44173 INVX1_LOC_95/Y NOR2X1_LOC_9/Y 0.10fF
C44174 NOR2X1_LOC_448/Y INVX1_LOC_295/Y 0.07fF
C44175 INVX1_LOC_58/A NOR2X1_LOC_533/Y 0.04fF
C44176 NAND2X1_LOC_570/Y INVX1_LOC_203/A 0.02fF
C44177 INPUT_0 INVX1_LOC_76/A 2.52fF
C44178 INVX1_LOC_124/A INVX1_LOC_19/A 0.05fF
C44179 D_GATE_366 INVX1_LOC_38/A 0.03fF
C44180 INVX1_LOC_144/A NAND2X1_LOC_453/A 0.01fF
C44181 NOR2X1_LOC_679/B NOR2X1_LOC_48/B 0.04fF
C44182 INVX1_LOC_90/A NAND2X1_LOC_617/a_36_24# 0.00fF
C44183 NOR2X1_LOC_476/Y INVX1_LOC_175/A 0.01fF
C44184 NOR2X1_LOC_389/A INVX1_LOC_57/A 0.00fF
C44185 INVX1_LOC_200/A NAND2X1_LOC_793/B 0.15fF
C44186 INVX1_LOC_10/A NOR2X1_LOC_592/B 0.11fF
C44187 INVX1_LOC_50/A NOR2X1_LOC_441/Y 0.11fF
C44188 NAND2X1_LOC_773/Y INVX1_LOC_306/Y 0.03fF
C44189 NAND2X1_LOC_579/A NOR2X1_LOC_406/A 0.02fF
C44190 INVX1_LOC_27/A NAND2X1_LOC_748/a_36_24# 0.00fF
C44191 NOR2X1_LOC_289/Y INVX1_LOC_38/A 0.04fF
C44192 NOR2X1_LOC_13/Y INVX1_LOC_94/Y 0.55fF
C44193 NOR2X1_LOC_791/B INVX1_LOC_16/Y 1.45fF
C44194 NOR2X1_LOC_497/Y INVX1_LOC_118/A 0.69fF
C44195 NAND2X1_LOC_850/Y NAND2X1_LOC_81/B 0.07fF
C44196 INVX1_LOC_89/A NOR2X1_LOC_634/A 0.01fF
C44197 NOR2X1_LOC_433/A NOR2X1_LOC_334/Y 0.19fF
C44198 NOR2X1_LOC_791/a_36_216# INVX1_LOC_23/Y 0.01fF
C44199 INVX1_LOC_313/Y INVX1_LOC_92/A 0.03fF
C44200 NAND2X1_LOC_466/Y INVX1_LOC_15/A 0.10fF
C44201 NOR2X1_LOC_413/Y INVX1_LOC_15/A 0.01fF
C44202 NOR2X1_LOC_595/Y INVX1_LOC_20/A 0.03fF
C44203 NAND2X1_LOC_364/A NOR2X1_LOC_383/B 0.03fF
C44204 NOR2X1_LOC_687/Y INVX1_LOC_19/A 0.03fF
C44205 NOR2X1_LOC_593/Y NOR2X1_LOC_334/Y 0.07fF
C44206 NOR2X1_LOC_377/a_36_216# INVX1_LOC_117/A 0.01fF
C44207 NAND2X1_LOC_649/B INVX1_LOC_76/A 0.01fF
C44208 NAND2X1_LOC_725/A NOR2X1_LOC_599/Y 0.06fF
C44209 NOR2X1_LOC_791/B NAND2X1_LOC_205/A 0.03fF
C44210 INVX1_LOC_234/A INVX1_LOC_203/A 0.10fF
C44211 NAND2X1_LOC_563/A NOR2X1_LOC_847/A 0.21fF
C44212 NOR2X1_LOC_736/Y INVX1_LOC_179/A 0.05fF
C44213 NAND2X1_LOC_352/a_36_24# NOR2X1_LOC_652/Y 0.01fF
C44214 INVX1_LOC_5/A NOR2X1_LOC_160/B 0.19fF
C44215 NAND2X1_LOC_579/A NAND2X1_LOC_493/Y 0.04fF
C44216 NOR2X1_LOC_130/A INVX1_LOC_3/A 0.03fF
C44217 INVX1_LOC_77/A INVX1_LOC_26/Y 0.03fF
C44218 INVX1_LOC_72/A INVX1_LOC_53/A 0.14fF
C44219 NOR2X1_LOC_201/A NOR2X1_LOC_860/B 0.01fF
C44220 NOR2X1_LOC_186/Y NAND2X1_LOC_336/a_36_24# 0.00fF
C44221 NAND2X1_LOC_540/a_36_24# INVX1_LOC_43/Y 0.00fF
C44222 NAND2X1_LOC_563/A INVX1_LOC_42/A 0.04fF
C44223 INVX1_LOC_62/Y INVX1_LOC_57/A 0.01fF
C44224 NOR2X1_LOC_439/B NOR2X1_LOC_155/A 0.01fF
C44225 INVX1_LOC_49/A NOR2X1_LOC_318/A 0.06fF
C44226 INVX1_LOC_33/A NAND2X1_LOC_91/a_36_24# 0.01fF
C44227 INVX1_LOC_178/A NAND2X1_LOC_550/A 0.10fF
C44228 NOR2X1_LOC_312/Y INVX1_LOC_63/A 0.30fF
C44229 NOR2X1_LOC_52/B NOR2X1_LOC_334/Y 0.07fF
C44230 NAND2X1_LOC_753/a_36_24# NOR2X1_LOC_703/B 0.00fF
C44231 NAND2X1_LOC_814/a_36_24# INVX1_LOC_118/A 0.00fF
C44232 INVX1_LOC_75/A NOR2X1_LOC_155/A 0.15fF
C44233 NOR2X1_LOC_430/A INVX1_LOC_296/A 0.04fF
C44234 NOR2X1_LOC_92/Y NAND2X1_LOC_799/A 0.03fF
C44235 NAND2X1_LOC_573/Y NAND2X1_LOC_336/a_36_24# 0.00fF
C44236 INVX1_LOC_41/A NOR2X1_LOC_843/B 0.03fF
C44237 INVX1_LOC_150/A INVX1_LOC_29/A 0.01fF
C44238 INVX1_LOC_5/A NAND2X1_LOC_195/Y 0.05fF
C44239 INVX1_LOC_36/A INVX1_LOC_50/Y 0.03fF
C44240 NAND2X1_LOC_585/a_36_24# INVX1_LOC_271/A 0.00fF
C44241 INVX1_LOC_11/A INVX1_LOC_308/Y 0.49fF
C44242 NAND2X1_LOC_325/Y NOR2X1_LOC_654/A 1.05fF
C44243 NOR2X1_LOC_82/Y INVX1_LOC_47/Y 0.23fF
C44244 NOR2X1_LOC_19/B INVX1_LOC_203/A 0.10fF
C44245 INVX1_LOC_89/A INVX1_LOC_29/A 0.13fF
C44246 INVX1_LOC_50/A NOR2X1_LOC_142/Y 0.03fF
C44247 INVX1_LOC_298/Y NOR2X1_LOC_493/B 0.10fF
C44248 NOR2X1_LOC_594/Y NOR2X1_LOC_697/Y 0.05fF
C44249 NOR2X1_LOC_589/A D_INPUT_5 0.02fF
C44250 NOR2X1_LOC_15/Y INVX1_LOC_31/A 0.11fF
C44251 INVX1_LOC_58/A NAND2X1_LOC_673/a_36_24# 0.00fF
C44252 NOR2X1_LOC_295/Y INVX1_LOC_57/A 0.02fF
C44253 INVX1_LOC_49/A NOR2X1_LOC_678/A 0.03fF
C44254 NOR2X1_LOC_45/B NOR2X1_LOC_487/Y 0.05fF
C44255 NOR2X1_LOC_824/A NOR2X1_LOC_372/Y 0.04fF
C44256 NOR2X1_LOC_124/B NAND2X1_LOC_205/A 0.35fF
C44257 INVX1_LOC_49/A INVX1_LOC_295/Y 0.01fF
C44258 INVX1_LOC_213/Y NOR2X1_LOC_858/A 0.02fF
C44259 NAND2X1_LOC_508/A INVX1_LOC_29/A 0.01fF
C44260 NOR2X1_LOC_357/Y INVX1_LOC_44/A 0.03fF
C44261 NOR2X1_LOC_828/Y NOR2X1_LOC_317/B 0.06fF
C44262 INVX1_LOC_28/A INVX1_LOC_272/A 0.07fF
C44263 INVX1_LOC_292/A NOR2X1_LOC_457/A 0.07fF
C44264 NOR2X1_LOC_332/A NOR2X1_LOC_554/A 0.01fF
C44265 NOR2X1_LOC_669/Y NAND2X1_LOC_721/B 0.08fF
C44266 INVX1_LOC_90/A INVX1_LOC_102/A 0.09fF
C44267 NAND2X1_LOC_564/B NAND2X1_LOC_471/Y 0.00fF
C44268 NOR2X1_LOC_6/B NOR2X1_LOC_416/A 0.03fF
C44269 NOR2X1_LOC_551/B INVX1_LOC_292/Y 0.16fF
C44270 NOR2X1_LOC_216/B INVX1_LOC_91/A 0.12fF
C44271 NAND2X1_LOC_581/Y INPUT_6 0.01fF
C44272 INVX1_LOC_30/Y NOR2X1_LOC_80/Y 0.06fF
C44273 NAND2X1_LOC_139/A NOR2X1_LOC_660/Y 0.00fF
C44274 NOR2X1_LOC_92/Y INVX1_LOC_18/A 0.17fF
C44275 INVX1_LOC_256/Y INVX1_LOC_181/A 0.08fF
C44276 INVX1_LOC_276/A NOR2X1_LOC_654/A 0.03fF
C44277 NAND2X1_LOC_787/A INVX1_LOC_240/A 0.03fF
C44278 NAND2X1_LOC_141/A INVX1_LOC_23/A 0.00fF
C44279 INVX1_LOC_1/A NOR2X1_LOC_354/B 0.01fF
C44280 INVX1_LOC_64/A NOR2X1_LOC_843/A 2.54fF
C44281 INVX1_LOC_230/Y INPUT_3 0.00fF
C44282 NOR2X1_LOC_510/Y NAND2X1_LOC_593/Y 0.02fF
C44283 INVX1_LOC_24/Y INVX1_LOC_18/A 0.11fF
C44284 INVX1_LOC_34/A NOR2X1_LOC_178/Y 0.07fF
C44285 NOR2X1_LOC_411/Y INVX1_LOC_237/Y 0.03fF
C44286 INVX1_LOC_15/Y INVX1_LOC_23/A 0.03fF
C44287 INVX1_LOC_269/A NOR2X1_LOC_554/B 0.01fF
C44288 NOR2X1_LOC_382/Y NOR2X1_LOC_82/A 0.01fF
C44289 INVX1_LOC_304/Y NAND2X1_LOC_793/B 0.07fF
C44290 NAND2X1_LOC_214/B NAND2X1_LOC_276/Y 0.03fF
C44291 INVX1_LOC_192/Y INVX1_LOC_53/A 0.01fF
C44292 INVX1_LOC_225/Y NOR2X1_LOC_565/A 0.00fF
C44293 NOR2X1_LOC_667/Y INVX1_LOC_286/Y 0.03fF
C44294 NOR2X1_LOC_401/Y NAND2X1_LOC_860/A 0.03fF
C44295 INVX1_LOC_64/A NOR2X1_LOC_399/A 0.02fF
C44296 INVX1_LOC_225/Y NOR2X1_LOC_169/B 0.03fF
C44297 NAND2X1_LOC_290/a_36_24# INVX1_LOC_23/A 0.01fF
C44298 VDD INVX1_LOC_185/A 0.76fF
C44299 INVX1_LOC_2/A NOR2X1_LOC_678/A 0.03fF
C44300 NAND2X1_LOC_728/Y NAND2X1_LOC_568/A 0.01fF
C44301 NOR2X1_LOC_843/A NOR2X1_LOC_436/a_36_216# 0.00fF
C44302 NOR2X1_LOC_666/Y NOR2X1_LOC_596/A 0.07fF
C44303 NAND2X1_LOC_139/a_36_24# NOR2X1_LOC_660/Y 0.00fF
C44304 NOR2X1_LOC_130/A NAND2X1_LOC_470/B 0.12fF
C44305 INVX1_LOC_292/A INVX1_LOC_30/A 0.11fF
C44306 NOR2X1_LOC_604/Y NOR2X1_LOC_78/B 0.01fF
C44307 INVX1_LOC_10/A NOR2X1_LOC_449/A 0.13fF
C44308 INVX1_LOC_27/A NAND2X1_LOC_276/Y 0.03fF
C44309 INVX1_LOC_258/Y INVX1_LOC_207/A 0.05fF
C44310 NOR2X1_LOC_92/Y INVX1_LOC_172/A 0.17fF
C44311 NOR2X1_LOC_500/Y NOR2X1_LOC_493/A 0.02fF
C44312 NOR2X1_LOC_78/A INVX1_LOC_293/Y 0.10fF
C44313 NAND2X1_LOC_323/B INVX1_LOC_53/A 0.03fF
C44314 INVX1_LOC_58/A INVX1_LOC_56/Y 0.00fF
C44315 NOR2X1_LOC_215/a_36_216# NOR2X1_LOC_759/Y 0.00fF
C44316 INVX1_LOC_177/A NOR2X1_LOC_674/a_36_216# 0.00fF
C44317 INVX1_LOC_100/A INVX1_LOC_168/Y 0.00fF
C44318 INVX1_LOC_256/A INVX1_LOC_24/A 0.10fF
C44319 INVX1_LOC_64/A NOR2X1_LOC_526/Y 0.01fF
C44320 NAND2X1_LOC_149/Y NOR2X1_LOC_770/B 0.02fF
C44321 INVX1_LOC_13/Y NOR2X1_LOC_84/Y 0.19fF
C44322 INVX1_LOC_200/A INVX1_LOC_71/A 0.25fF
C44323 NOR2X1_LOC_557/A INVX1_LOC_125/A 0.52fF
C44324 INVX1_LOC_298/Y INVX1_LOC_89/A 0.04fF
C44325 NOR2X1_LOC_626/a_36_216# INVX1_LOC_266/Y 0.00fF
C44326 NOR2X1_LOC_453/Y INVX1_LOC_103/Y 0.01fF
C44327 INVX1_LOC_98/A NAND2X1_LOC_74/B 0.02fF
C44328 INPUT_0 INVX1_LOC_127/Y 0.01fF
C44329 INVX1_LOC_36/A NOR2X1_LOC_248/Y 0.01fF
C44330 NOR2X1_LOC_351/Y INVX1_LOC_118/Y 0.02fF
C44331 NOR2X1_LOC_91/A NOR2X1_LOC_576/B 0.05fF
C44332 NOR2X1_LOC_78/A NAND2X1_LOC_74/B 0.18fF
C44333 INVX1_LOC_5/A NAND2X1_LOC_350/B 0.01fF
C44334 INVX1_LOC_222/Y NOR2X1_LOC_168/B 0.03fF
C44335 INVX1_LOC_161/Y INVX1_LOC_77/A 0.15fF
C44336 NAND2X1_LOC_708/Y INVX1_LOC_16/A 0.04fF
C44337 INVX1_LOC_119/Y INVX1_LOC_46/A 0.03fF
C44338 INVX1_LOC_5/A INVX1_LOC_208/A 0.01fF
C44339 NOR2X1_LOC_770/A INVX1_LOC_174/A 0.02fF
C44340 NAND2X1_LOC_475/Y NOR2X1_LOC_137/Y 0.34fF
C44341 NOR2X1_LOC_280/Y NOR2X1_LOC_661/A 0.06fF
C44342 NAND2X1_LOC_35/Y INVX1_LOC_22/A 0.13fF
C44343 NOR2X1_LOC_590/A NOR2X1_LOC_419/a_36_216# 0.00fF
C44344 NOR2X1_LOC_606/Y INVX1_LOC_24/A 0.00fF
C44345 INVX1_LOC_204/A INVX1_LOC_89/A 0.01fF
C44346 INVX1_LOC_11/A NOR2X1_LOC_162/Y 0.01fF
C44347 NOR2X1_LOC_331/B INVX1_LOC_307/A 0.07fF
C44348 NOR2X1_LOC_860/B INVX1_LOC_31/A 0.07fF
C44349 NOR2X1_LOC_599/Y NOR2X1_LOC_387/a_36_216# 0.00fF
C44350 INVX1_LOC_5/A NOR2X1_LOC_516/B 0.11fF
C44351 NAND2X1_LOC_740/B NAND2X1_LOC_175/Y 0.05fF
C44352 NOR2X1_LOC_653/B NOR2X1_LOC_773/Y 0.13fF
C44353 NOR2X1_LOC_824/A NAND2X1_LOC_374/Y 1.64fF
C44354 NAND2X1_LOC_287/B INVX1_LOC_63/A 0.07fF
C44355 INVX1_LOC_36/A NAND2X1_LOC_356/a_36_24# 0.00fF
C44356 NOR2X1_LOC_78/B NOR2X1_LOC_857/a_36_216# 0.00fF
C44357 INVX1_LOC_33/Y INVX1_LOC_285/A 0.02fF
C44358 NAND2X1_LOC_11/Y NOR2X1_LOC_763/A 0.34fF
C44359 NOR2X1_LOC_15/Y NOR2X1_LOC_290/Y 0.35fF
C44360 NOR2X1_LOC_74/A INVX1_LOC_271/Y 0.17fF
C44361 INVX1_LOC_37/A NOR2X1_LOC_257/Y 0.01fF
C44362 INVX1_LOC_11/A NOR2X1_LOC_718/B 0.18fF
C44363 NAND2X1_LOC_11/Y NOR2X1_LOC_582/A 0.14fF
C44364 NOR2X1_LOC_679/Y NAND2X1_LOC_354/B 0.15fF
C44365 NOR2X1_LOC_15/Y INVX1_LOC_191/Y 0.14fF
C44366 INVX1_LOC_129/Y INVX1_LOC_63/A 0.07fF
C44367 NOR2X1_LOC_384/a_36_216# NAND2X1_LOC_837/Y 0.01fF
C44368 NAND2X1_LOC_391/a_36_24# INVX1_LOC_61/A 0.01fF
C44369 NAND2X1_LOC_182/A NAND2X1_LOC_793/Y 0.50fF
C44370 NAND2X1_LOC_464/A NAND2X1_LOC_74/B 0.06fF
C44371 NOR2X1_LOC_459/A NOR2X1_LOC_663/A 0.02fF
C44372 INVX1_LOC_18/A NAND2X1_LOC_837/Y 0.10fF
C44373 INVX1_LOC_50/A INVX1_LOC_182/A 0.07fF
C44374 INVX1_LOC_239/A INVX1_LOC_84/Y 0.01fF
C44375 INVX1_LOC_313/Y INVX1_LOC_53/A 0.15fF
C44376 NAND2X1_LOC_778/Y NAND2X1_LOC_859/Y 0.28fF
C44377 VDD INVX1_LOC_69/A -0.00fF
C44378 INVX1_LOC_46/A INVX1_LOC_284/A 0.00fF
C44379 INVX1_LOC_256/A INVX1_LOC_143/A 0.03fF
C44380 INVX1_LOC_183/A NOR2X1_LOC_167/Y 0.01fF
C44381 NOR2X1_LOC_276/a_36_216# INVX1_LOC_77/A 0.02fF
C44382 NOR2X1_LOC_212/a_36_216# INVX1_LOC_171/A 0.00fF
C44383 NOR2X1_LOC_98/a_36_216# NAND2X1_LOC_74/B 0.00fF
C44384 NOR2X1_LOC_45/B NAND2X1_LOC_454/Y 0.68fF
C44385 NOR2X1_LOC_598/B NOR2X1_LOC_439/B 0.21fF
C44386 INVX1_LOC_11/A INVX1_LOC_218/A 0.06fF
C44387 NOR2X1_LOC_88/a_36_216# NOR2X1_LOC_88/Y 0.00fF
C44388 INVX1_LOC_31/A NAND2X1_LOC_141/A 0.00fF
C44389 INVX1_LOC_110/Y NOR2X1_LOC_100/A 0.26fF
C44390 INVX1_LOC_174/A NAND2X1_LOC_451/Y 0.14fF
C44391 INVX1_LOC_136/A NAND2X1_LOC_139/A 0.01fF
C44392 INVX1_LOC_211/Y INVX1_LOC_144/Y 0.03fF
C44393 INVX1_LOC_41/A INVX1_LOC_18/A 0.09fF
C44394 INVX1_LOC_223/A NOR2X1_LOC_392/B 0.17fF
C44395 INVX1_LOC_69/Y NOR2X1_LOC_481/a_36_216# 0.01fF
C44396 NOR2X1_LOC_248/Y NOR2X1_LOC_309/Y 0.01fF
C44397 NOR2X1_LOC_89/A NAND2X1_LOC_472/Y 0.07fF
C44398 NOR2X1_LOC_15/Y NAND2X1_LOC_859/Y 0.98fF
C44399 INVX1_LOC_36/A NOR2X1_LOC_6/B 0.02fF
C44400 INVX1_LOC_172/A NAND2X1_LOC_837/Y 0.07fF
C44401 INVX1_LOC_94/A NOR2X1_LOC_577/Y 0.01fF
C44402 NOR2X1_LOC_437/Y INVX1_LOC_77/A 0.07fF
C44403 NOR2X1_LOC_598/B INVX1_LOC_75/A 1.39fF
C44404 INVX1_LOC_88/A INVX1_LOC_290/A 0.00fF
C44405 INVX1_LOC_93/A INVX1_LOC_183/Y 0.01fF
C44406 NOR2X1_LOC_738/A INVX1_LOC_213/A 0.04fF
C44407 NOR2X1_LOC_318/B NOR2X1_LOC_278/Y 0.00fF
C44408 INVX1_LOC_19/A INVX1_LOC_9/A 0.50fF
C44409 INVX1_LOC_12/Y INVX1_LOC_42/A 0.37fF
C44410 NOR2X1_LOC_160/B NOR2X1_LOC_773/Y 0.07fF
C44411 NOR2X1_LOC_639/B INVX1_LOC_302/A 0.02fF
C44412 NOR2X1_LOC_89/A NAND2X1_LOC_603/a_36_24# 0.01fF
C44413 INVX1_LOC_303/A NOR2X1_LOC_350/A 0.01fF
C44414 INVX1_LOC_57/Y NAND2X1_LOC_785/A 0.01fF
C44415 NAND2X1_LOC_53/Y NAND2X1_LOC_479/Y 0.07fF
C44416 INVX1_LOC_150/Y INVX1_LOC_16/A 0.68fF
C44417 INVX1_LOC_11/A NOR2X1_LOC_569/Y 0.07fF
C44418 INVX1_LOC_93/Y NOR2X1_LOC_278/Y 0.07fF
C44419 INVX1_LOC_97/Y INVX1_LOC_75/A 0.05fF
C44420 INVX1_LOC_12/A NOR2X1_LOC_331/B 1.29fF
C44421 INVX1_LOC_31/A INVX1_LOC_226/A 0.03fF
C44422 INVX1_LOC_233/Y INVX1_LOC_282/A 0.10fF
C44423 INVX1_LOC_31/A NAND2X1_LOC_840/B 2.25fF
C44424 INVX1_LOC_102/A INVX1_LOC_38/A 0.08fF
C44425 NOR2X1_LOC_716/B NOR2X1_LOC_753/Y 0.06fF
C44426 NOR2X1_LOC_419/Y NOR2X1_LOC_520/B 0.01fF
C44427 INVX1_LOC_223/A NAND2X1_LOC_294/a_36_24# 0.00fF
C44428 INVX1_LOC_304/A INVX1_LOC_26/A 0.07fF
C44429 NOR2X1_LOC_207/A INVX1_LOC_18/A 0.01fF
C44430 NOR2X1_LOC_607/A INVX1_LOC_104/A 0.02fF
C44431 NAND2X1_LOC_295/a_36_24# INVX1_LOC_38/A 0.00fF
C44432 INVX1_LOC_182/Y NOR2X1_LOC_644/a_36_216# 0.00fF
C44433 NAND2X1_LOC_99/Y NAND2X1_LOC_276/Y 0.08fF
C44434 NOR2X1_LOC_658/Y INVX1_LOC_52/A 0.01fF
C44435 NOR2X1_LOC_78/B INVX1_LOC_72/A 0.09fF
C44436 NOR2X1_LOC_178/Y INPUT_0 0.09fF
C44437 NOR2X1_LOC_405/A NOR2X1_LOC_383/B 0.03fF
C44438 NAND2X1_LOC_35/Y INVX1_LOC_100/A -0.00fF
C44439 NOR2X1_LOC_434/Y INPUT_0 0.02fF
C44440 NAND2X1_LOC_563/A NOR2X1_LOC_554/B 0.09fF
C44441 INVX1_LOC_314/Y NOR2X1_LOC_709/A 0.17fF
C44442 NOR2X1_LOC_329/B NAND2X1_LOC_780/Y 0.01fF
C44443 NOR2X1_LOC_160/B NOR2X1_LOC_332/A 0.11fF
C44444 NOR2X1_LOC_718/B NOR2X1_LOC_593/Y 0.01fF
C44445 INVX1_LOC_12/Y INVX1_LOC_78/A 1.04fF
C44446 INVX1_LOC_12/A NOR2X1_LOC_592/B 0.07fF
C44447 NOR2X1_LOC_824/A NAND2X1_LOC_844/a_36_24# 0.01fF
C44448 NAND2X1_LOC_477/Y INVX1_LOC_203/A 0.06fF
C44449 INVX1_LOC_21/A NOR2X1_LOC_368/A 0.03fF
C44450 INVX1_LOC_300/Y NAND2X1_LOC_852/Y 0.01fF
C44451 INVX1_LOC_36/A INVX1_LOC_30/Y 0.07fF
C44452 NOR2X1_LOC_220/a_36_216# NOR2X1_LOC_220/A 0.00fF
C44453 NAND2X1_LOC_213/A NOR2X1_LOC_163/Y 0.23fF
C44454 NOR2X1_LOC_533/Y NOR2X1_LOC_533/a_36_216# 0.00fF
C44455 INVX1_LOC_310/A NAND2X1_LOC_364/Y 0.15fF
C44456 NOR2X1_LOC_209/Y NOR2X1_LOC_550/B 0.10fF
C44457 NAND2X1_LOC_778/Y INVX1_LOC_6/A 0.05fF
C44458 NOR2X1_LOC_383/B NOR2X1_LOC_857/A 0.07fF
C44459 INVX1_LOC_72/Y NOR2X1_LOC_719/A 0.02fF
C44460 NOR2X1_LOC_657/Y INVX1_LOC_279/A 0.01fF
C44461 INVX1_LOC_5/A INVX1_LOC_315/Y 0.10fF
C44462 NAND2X1_LOC_67/Y INVX1_LOC_42/Y 0.04fF
C44463 NAND2X1_LOC_773/Y NOR2X1_LOC_74/A 0.10fF
C44464 INVX1_LOC_41/A INVX1_LOC_34/Y 0.03fF
C44465 NOR2X1_LOC_392/B NOR2X1_LOC_316/Y 0.01fF
C44466 NOR2X1_LOC_65/B INVX1_LOC_12/Y 0.10fF
C44467 NOR2X1_LOC_205/a_36_216# NOR2X1_LOC_577/Y 0.01fF
C44468 VDD INVX1_LOC_270/Y 1.14fF
C44469 INVX1_LOC_63/Y NAND2X1_LOC_661/B 0.00fF
C44470 INVX1_LOC_121/A INVX1_LOC_18/A 0.02fF
C44471 NOR2X1_LOC_136/Y NOR2X1_LOC_577/Y 0.01fF
C44472 NOR2X1_LOC_798/A NOR2X1_LOC_334/a_36_216# 0.00fF
C44473 INVX1_LOC_83/A INVX1_LOC_72/A 0.10fF
C44474 NAND2X1_LOC_350/A NAND2X1_LOC_652/Y 0.02fF
C44475 D_INPUT_1 D_INPUT_3 0.76fF
C44476 INVX1_LOC_166/A INVX1_LOC_194/Y 0.03fF
C44477 NOR2X1_LOC_222/Y NOR2X1_LOC_219/B 0.01fF
C44478 NOR2X1_LOC_488/a_36_216# NOR2X1_LOC_716/B 0.01fF
C44479 NAND2X1_LOC_722/A INVX1_LOC_240/A 0.07fF
C44480 NAND2X1_LOC_773/Y NOR2X1_LOC_9/Y 0.29fF
C44481 D_INPUT_1 INVX1_LOC_14/Y 0.03fF
C44482 INVX1_LOC_83/A INVX1_LOC_142/Y 0.01fF
C44483 INVX1_LOC_262/Y NAND2X1_LOC_651/B 0.21fF
C44484 NOR2X1_LOC_15/Y INVX1_LOC_6/A 0.09fF
C44485 NOR2X1_LOC_197/A NOR2X1_LOC_742/A 0.02fF
C44486 NOR2X1_LOC_84/Y INVX1_LOC_168/A 0.03fF
C44487 VDD NOR2X1_LOC_754/Y 0.44fF
C44488 INVX1_LOC_90/A INVX1_LOC_223/A 0.03fF
C44489 NOR2X1_LOC_554/B NOR2X1_LOC_814/Y 0.12fF
C44490 INVX1_LOC_83/A INVX1_LOC_198/Y 0.03fF
C44491 INVX1_LOC_26/Y INVX1_LOC_9/A 0.10fF
C44492 NOR2X1_LOC_388/Y NOR2X1_LOC_500/Y 0.09fF
C44493 NOR2X1_LOC_334/Y NOR2X1_LOC_858/a_36_216# 0.01fF
C44494 NOR2X1_LOC_329/B INVX1_LOC_141/Y 0.07fF
C44495 NOR2X1_LOC_318/A INVX1_LOC_118/A 0.00fF
C44496 INVX1_LOC_171/A NOR2X1_LOC_360/Y 0.03fF
C44497 NOR2X1_LOC_592/a_36_216# INVX1_LOC_144/A 0.01fF
C44498 NAND2X1_LOC_802/A NOR2X1_LOC_561/Y 0.01fF
C44499 INVX1_LOC_109/A INVX1_LOC_272/A 0.01fF
C44500 INVX1_LOC_45/Y NOR2X1_LOC_355/A 0.40fF
C44501 NOR2X1_LOC_177/Y NOR2X1_LOC_301/A 0.10fF
C44502 NOR2X1_LOC_618/a_36_216# INVX1_LOC_8/A 0.01fF
C44503 NAND2X1_LOC_725/A NAND2X1_LOC_453/A 0.03fF
C44504 NOR2X1_LOC_329/B INVX1_LOC_312/Y 0.20fF
C44505 NOR2X1_LOC_643/Y INVX1_LOC_7/A 0.00fF
C44506 NOR2X1_LOC_301/A NOR2X1_LOC_743/Y 0.04fF
C44507 NOR2X1_LOC_700/Y NAND2X1_LOC_866/A 0.02fF
C44508 INVX1_LOC_228/A INVX1_LOC_89/A 0.43fF
C44509 NOR2X1_LOC_440/Y NOR2X1_LOC_557/Y 0.02fF
C44510 NOR2X1_LOC_861/Y INVX1_LOC_19/A 0.07fF
C44511 NAND2X1_LOC_338/B NOR2X1_LOC_547/B 0.03fF
C44512 NOR2X1_LOC_78/B NAND2X1_LOC_338/B 1.30fF
C44513 INVX1_LOC_207/A INVX1_LOC_229/Y 0.07fF
C44514 NAND2X1_LOC_323/B NOR2X1_LOC_634/B 0.03fF
C44515 NOR2X1_LOC_388/Y INVX1_LOC_10/A 0.07fF
C44516 NOR2X1_LOC_758/Y NAND2X1_LOC_573/A 0.00fF
C44517 NAND2X1_LOC_323/B NOR2X1_LOC_547/B -0.00fF
C44518 INVX1_LOC_262/Y INVX1_LOC_15/A 0.01fF
C44519 NOR2X1_LOC_214/B INVX1_LOC_113/Y 0.01fF
C44520 NAND2X1_LOC_267/B NOR2X1_LOC_440/B 0.14fF
C44521 NAND2X1_LOC_112/Y NOR2X1_LOC_111/a_36_216# 0.00fF
C44522 INVX1_LOC_46/A NOR2X1_LOC_384/A 0.01fF
C44523 NAND2X1_LOC_799/A NAND2X1_LOC_648/a_36_24# 0.00fF
C44524 INVX1_LOC_53/A NOR2X1_LOC_506/Y 0.06fF
C44525 NAND2X1_LOC_639/a_36_24# NOR2X1_LOC_467/A 0.01fF
C44526 NOR2X1_LOC_554/A NOR2X1_LOC_847/A 0.19fF
C44527 NOR2X1_LOC_685/B NAND2X1_LOC_782/B 0.04fF
C44528 NOR2X1_LOC_276/Y NOR2X1_LOC_78/A 0.03fF
C44529 NAND2X1_LOC_633/a_36_24# NAND2X1_LOC_392/Y 0.00fF
C44530 INVX1_LOC_18/A NAND2X1_LOC_662/B 0.76fF
C44531 INVX1_LOC_89/A INVX1_LOC_8/A 0.10fF
C44532 NAND2X1_LOC_574/A NOR2X1_LOC_843/B 0.07fF
C44533 NOR2X1_LOC_440/Y INVX1_LOC_143/A 0.01fF
C44534 NOR2X1_LOC_385/a_36_216# INVX1_LOC_231/Y 0.00fF
C44535 INVX1_LOC_90/A INVX1_LOC_149/Y 0.03fF
C44536 INVX1_LOC_80/A INVX1_LOC_216/A 0.19fF
C44537 INVX1_LOC_223/A NAND2X1_LOC_123/a_36_24# 0.00fF
C44538 INVX1_LOC_90/A INVX1_LOC_162/Y 0.01fF
C44539 INVX1_LOC_39/A NOR2X1_LOC_99/a_36_216# 0.00fF
C44540 INVX1_LOC_36/A INVX1_LOC_96/A 0.00fF
C44541 NAND2X1_LOC_162/a_36_24# INVX1_LOC_33/A 0.01fF
C44542 INVX1_LOC_83/A INVX1_LOC_192/Y 0.34fF
C44543 INVX1_LOC_90/A INVX1_LOC_85/A 0.03fF
C44544 NAND2X1_LOC_213/a_36_24# NOR2X1_LOC_467/A 0.01fF
C44545 INVX1_LOC_83/A NOR2X1_LOC_537/Y 0.02fF
C44546 NAND2X1_LOC_338/B INVX1_LOC_83/A 0.07fF
C44547 INVX1_LOC_17/A INVX1_LOC_37/A 0.45fF
C44548 INVX1_LOC_24/A INVX1_LOC_69/Y 0.07fF
C44549 INVX1_LOC_90/A NOR2X1_LOC_316/Y 0.01fF
C44550 NAND2X1_LOC_736/Y NAND2X1_LOC_560/A 0.20fF
C44551 INVX1_LOC_136/A NOR2X1_LOC_78/A 0.04fF
C44552 INVX1_LOC_135/A INVX1_LOC_197/A 0.15fF
C44553 NOR2X1_LOC_478/A INVX1_LOC_199/Y 0.12fF
C44554 NOR2X1_LOC_577/Y INVX1_LOC_144/A 0.03fF
C44555 NAND2X1_LOC_53/Y INVX1_LOC_139/Y 0.01fF
C44556 INVX1_LOC_124/Y INVX1_LOC_95/Y 0.98fF
C44557 NAND2X1_LOC_323/B INVX1_LOC_83/A 0.04fF
C44558 NOR2X1_LOC_91/A INVX1_LOC_49/Y 0.06fF
C44559 NOR2X1_LOC_68/A NOR2X1_LOC_45/B 3.57fF
C44560 NAND2X1_LOC_456/Y INVX1_LOC_23/A 0.01fF
C44561 INVX1_LOC_12/A NOR2X1_LOC_449/A 0.03fF
C44562 INVX1_LOC_277/A NOR2X1_LOC_833/Y 0.38fF
C44563 INVX1_LOC_36/A NOR2X1_LOC_124/A 0.00fF
C44564 NOR2X1_LOC_287/A D_INPUT_0 0.04fF
C44565 INVX1_LOC_11/A NAND2X1_LOC_472/Y 0.07fF
C44566 NOR2X1_LOC_471/Y INVX1_LOC_37/A 0.03fF
C44567 INVX1_LOC_226/Y INVX1_LOC_135/A 0.10fF
C44568 D_GATE_741 INVX1_LOC_117/A 0.02fF
C44569 NOR2X1_LOC_516/B NOR2X1_LOC_332/A 1.58fF
C44570 NOR2X1_LOC_78/B INVX1_LOC_313/Y 0.13fF
C44571 NOR2X1_LOC_667/Y VDD 0.08fF
C44572 INVX1_LOC_233/A INVX1_LOC_119/Y 0.12fF
C44573 NOR2X1_LOC_191/A INPUT_1 0.01fF
C44574 NOR2X1_LOC_208/Y INVX1_LOC_96/A 0.02fF
C44575 NAND2X1_LOC_803/B INVX1_LOC_33/Y 0.00fF
C44576 NOR2X1_LOC_791/A INVX1_LOC_95/Y 0.01fF
C44577 INVX1_LOC_133/A INVX1_LOC_270/Y 0.96fF
C44578 NOR2X1_LOC_500/A INVX1_LOC_91/A 0.05fF
C44579 NAND2X1_LOC_114/B NOR2X1_LOC_107/a_36_216# 0.01fF
C44580 NOR2X1_LOC_303/Y INVX1_LOC_91/A 0.28fF
C44581 NOR2X1_LOC_67/A NOR2X1_LOC_120/a_36_216# 0.00fF
C44582 NOR2X1_LOC_785/A INVX1_LOC_117/A 0.01fF
C44583 NOR2X1_LOC_68/A INVX1_LOC_199/Y 0.00fF
C44584 INVX1_LOC_75/A NOR2X1_LOC_156/B 0.12fF
C44585 NOR2X1_LOC_72/a_36_216# INVX1_LOC_53/Y 0.01fF
C44586 INVX1_LOC_48/Y NOR2X1_LOC_99/Y 0.02fF
C44587 NOR2X1_LOC_230/Y VDD 0.13fF
C44588 INVX1_LOC_226/Y NOR2X1_LOC_560/A 0.01fF
C44589 NAND2X1_LOC_543/Y INVX1_LOC_90/A 0.18fF
C44590 NOR2X1_LOC_590/A INVX1_LOC_33/Y 0.01fF
C44591 NOR2X1_LOC_15/Y NOR2X1_LOC_79/A 0.21fF
C44592 NOR2X1_LOC_584/Y NOR2X1_LOC_654/A 0.27fF
C44593 INVX1_LOC_23/A NAND2X1_LOC_80/a_36_24# 0.00fF
C44594 INVX1_LOC_90/A NOR2X1_LOC_94/a_36_216# 0.00fF
C44595 INVX1_LOC_299/A NOR2X1_LOC_640/Y 0.01fF
C44596 INVX1_LOC_72/Y INVX1_LOC_76/A 0.02fF
C44597 INVX1_LOC_72/A INVX1_LOC_46/A 0.35fF
C44598 INVX1_LOC_161/Y INVX1_LOC_9/A 0.09fF
C44599 INVX1_LOC_11/A NAND2X1_LOC_637/Y 0.07fF
C44600 NOR2X1_LOC_470/B NAND2X1_LOC_93/B 0.01fF
C44601 INVX1_LOC_23/A INVX1_LOC_99/A 0.04fF
C44602 NAND2X1_LOC_254/Y NAND2X1_LOC_464/B 0.03fF
C44603 INVX1_LOC_35/A NAND2X1_LOC_82/Y 0.07fF
C44604 INVX1_LOC_111/Y NOR2X1_LOC_335/B 0.02fF
C44605 NOR2X1_LOC_742/A INVX1_LOC_83/Y 0.01fF
C44606 NOR2X1_LOC_360/Y NOR2X1_LOC_360/A 0.00fF
C44607 NOR2X1_LOC_392/Y INVX1_LOC_29/A 0.07fF
C44608 INVX1_LOC_33/A NOR2X1_LOC_746/Y 0.15fF
C44609 NOR2X1_LOC_254/Y INVX1_LOC_91/A 0.72fF
C44610 INVX1_LOC_50/Y INVX1_LOC_63/A 10.58fF
C44611 NOR2X1_LOC_249/Y NOR2X1_LOC_814/A 0.11fF
C44612 NOR2X1_LOC_471/Y NAND2X1_LOC_629/a_36_24# 0.01fF
C44613 INVX1_LOC_286/Y NOR2X1_LOC_536/A 0.03fF
C44614 INVX1_LOC_96/Y INVX1_LOC_6/A 0.78fF
C44615 NOR2X1_LOC_470/B NAND2X1_LOC_425/Y 0.02fF
C44616 INVX1_LOC_215/A NOR2X1_LOC_111/Y 0.04fF
C44617 INVX1_LOC_136/A NOR2X1_LOC_60/Y 0.00fF
C44618 INVX1_LOC_1/A NAND2X1_LOC_141/Y 0.01fF
C44619 NOR2X1_LOC_561/a_36_216# INVX1_LOC_93/Y 0.01fF
C44620 NOR2X1_LOC_767/a_36_216# INVX1_LOC_286/A 0.01fF
C44621 NOR2X1_LOC_376/A INVX1_LOC_84/A 0.06fF
C44622 NOR2X1_LOC_248/a_36_216# INVX1_LOC_10/A 0.00fF
C44623 INVX1_LOC_223/A INVX1_LOC_38/A 0.03fF
C44624 D_INPUT_2 D_INPUT_3 2.94fF
C44625 NOR2X1_LOC_576/B NAND2X1_LOC_866/B 0.02fF
C44626 INVX1_LOC_5/A NAND2X1_LOC_207/B 4.55fF
C44627 NOR2X1_LOC_219/a_36_216# NOR2X1_LOC_357/Y 0.00fF
C44628 NOR2X1_LOC_720/A INVX1_LOC_4/Y 0.00fF
C44629 INVX1_LOC_256/A NOR2X1_LOC_197/B 0.10fF
C44630 NOR2X1_LOC_67/A NOR2X1_LOC_392/a_36_216# 0.00fF
C44631 INVX1_LOC_144/A INVX1_LOC_22/A 0.20fF
C44632 NOR2X1_LOC_329/B NAND2X1_LOC_656/Y 0.33fF
C44633 INVX1_LOC_54/Y INVX1_LOC_91/A 0.16fF
C44634 NOR2X1_LOC_186/Y NAND2X1_LOC_74/B 1.81fF
C44635 INVX1_LOC_207/A INVX1_LOC_20/A 8.35fF
C44636 INVX1_LOC_223/Y INVX1_LOC_29/A 0.09fF
C44637 NAND2X1_LOC_553/A INVX1_LOC_284/A 0.01fF
C44638 INVX1_LOC_14/A INVX1_LOC_84/A 0.92fF
C44639 NOR2X1_LOC_570/B NOR2X1_LOC_556/a_36_216# 0.00fF
C44640 NOR2X1_LOC_716/B NOR2X1_LOC_558/A 0.04fF
C44641 NAND2X1_LOC_355/Y NOR2X1_LOC_331/B 0.07fF
C44642 INVX1_LOC_284/Y NOR2X1_LOC_823/a_36_216# 0.02fF
C44643 INVX1_LOC_235/A INVX1_LOC_29/A 0.01fF
C44644 NAND2X1_LOC_811/Y INVX1_LOC_76/A 0.03fF
C44645 INVX1_LOC_217/Y NOR2X1_LOC_825/Y 0.00fF
C44646 NOR2X1_LOC_794/A NOR2X1_LOC_500/Y 0.01fF
C44647 INVX1_LOC_279/A NOR2X1_LOC_74/A 0.17fF
C44648 NAND2X1_LOC_573/Y NAND2X1_LOC_74/B 0.07fF
C44649 INVX1_LOC_45/A INVX1_LOC_92/A 0.11fF
C44650 INVX1_LOC_111/A NAND2X1_LOC_204/a_36_24# 0.02fF
C44651 NOR2X1_LOC_593/Y NAND2X1_LOC_472/Y 0.07fF
C44652 INVX1_LOC_266/Y INVX1_LOC_76/A 0.28fF
C44653 INVX1_LOC_11/A NAND2X1_LOC_773/B 0.07fF
C44654 NOR2X1_LOC_552/A NOR2X1_LOC_500/Y 0.12fF
C44655 NOR2X1_LOC_310/Y VDD 0.18fF
C44656 NOR2X1_LOC_721/Y NOR2X1_LOC_749/a_36_216# 0.03fF
C44657 NOR2X1_LOC_816/A NOR2X1_LOC_605/A 0.07fF
C44658 NOR2X1_LOC_529/Y D_INPUT_3 0.06fF
C44659 NOR2X1_LOC_211/Y INVX1_LOC_4/Y 0.00fF
C44660 D_INPUT_0 NAND2X1_LOC_519/a_36_24# 0.00fF
C44661 NOR2X1_LOC_589/A NOR2X1_LOC_269/Y 0.07fF
C44662 NAND2X1_LOC_189/a_36_24# NOR2X1_LOC_188/A 0.01fF
C44663 NAND2X1_LOC_357/A INVX1_LOC_29/A 0.08fF
C44664 NOR2X1_LOC_38/B INVX1_LOC_306/Y 0.10fF
C44665 INVX1_LOC_253/A INVX1_LOC_253/Y 0.14fF
C44666 INVX1_LOC_286/Y NOR2X1_LOC_661/A 0.01fF
C44667 NAND2X1_LOC_338/B INVX1_LOC_46/A 0.22fF
C44668 NOR2X1_LOC_332/A INVX1_LOC_315/Y 0.23fF
C44669 NAND2X1_LOC_338/B NOR2X1_LOC_98/A 0.01fF
C44670 INVX1_LOC_71/A INVX1_LOC_92/A 0.06fF
C44671 INVX1_LOC_246/A INVX1_LOC_272/A 0.01fF
C44672 INVX1_LOC_135/A NOR2X1_LOC_340/a_36_216# 0.00fF
C44673 INVX1_LOC_85/A INVX1_LOC_38/A 0.03fF
C44674 INVX1_LOC_31/A INVX1_LOC_49/Y 0.03fF
C44675 INVX1_LOC_182/Y NOR2X1_LOC_74/A 0.03fF
C44676 INVX1_LOC_110/Y NOR2X1_LOC_340/A 0.01fF
C44677 NOR2X1_LOC_261/a_36_216# NOR2X1_LOC_261/Y 0.15fF
C44678 INVX1_LOC_41/A NAND2X1_LOC_488/a_36_24# 0.00fF
C44679 NOR2X1_LOC_577/Y NOR2X1_LOC_155/A 0.05fF
C44680 NOR2X1_LOC_160/B NOR2X1_LOC_847/A 0.07fF
C44681 INVX1_LOC_14/A INVX1_LOC_15/A 0.07fF
C44682 NAND2X1_LOC_550/A INVX1_LOC_42/A 0.16fF
C44683 INVX1_LOC_13/Y INVX1_LOC_116/Y 0.00fF
C44684 NOR2X1_LOC_160/B INVX1_LOC_42/A 0.14fF
C44685 NOR2X1_LOC_45/B NOR2X1_LOC_163/A 0.01fF
C44686 D_INPUT_0 INVX1_LOC_95/Y 0.07fF
C44687 NOR2X1_LOC_387/A NOR2X1_LOC_409/Y 0.03fF
C44688 INVX1_LOC_170/A NAND2X1_LOC_74/B 0.02fF
C44689 NOR2X1_LOC_32/B NAND2X1_LOC_571/B 0.08fF
C44690 NAND2X1_LOC_858/B NOR2X1_LOC_74/A 0.14fF
C44691 INVX1_LOC_75/A INVX1_LOC_201/A 0.72fF
C44692 INVX1_LOC_214/Y NOR2X1_LOC_331/B 0.02fF
C44693 INVX1_LOC_33/A INVX1_LOC_123/Y 0.13fF
C44694 NAND2X1_LOC_645/a_36_24# NAND2X1_LOC_472/Y 0.00fF
C44695 NOR2X1_LOC_349/B VDD 0.12fF
C44696 NAND2X1_LOC_741/Y NAND2X1_LOC_725/Y 0.01fF
C44697 NAND2X1_LOC_740/Y NAND2X1_LOC_738/B 0.13fF
C44698 INVX1_LOC_25/A INVX1_LOC_13/Y 0.18fF
C44699 INVX1_LOC_280/Y INVX1_LOC_185/A 0.31fF
C44700 NOR2X1_LOC_733/Y INVX1_LOC_6/A 0.21fF
C44701 NOR2X1_LOC_627/Y INVX1_LOC_179/A 0.01fF
C44702 NOR2X1_LOC_15/Y INVX1_LOC_28/Y 0.02fF
C44703 NOR2X1_LOC_4/a_36_216# NOR2X1_LOC_649/B 0.01fF
C44704 NOR2X1_LOC_778/B NOR2X1_LOC_830/a_36_216# 0.00fF
C44705 NAND2X1_LOC_550/A INVX1_LOC_78/A 0.04fF
C44706 NOR2X1_LOC_717/Y INVX1_LOC_15/A 0.01fF
C44707 INVX1_LOC_11/A NAND2X1_LOC_70/a_36_24# 0.00fF
C44708 INVX1_LOC_24/A NOR2X1_LOC_89/A 0.16fF
C44709 NAND2X1_LOC_391/Y NAND2X1_LOC_860/A 0.04fF
C44710 INVX1_LOC_313/Y INVX1_LOC_46/A 0.07fF
C44711 INVX1_LOC_50/A NAND2X1_LOC_579/A 1.52fF
C44712 NOR2X1_LOC_160/B INVX1_LOC_78/A 0.10fF
C44713 NOR2X1_LOC_667/a_36_216# INVX1_LOC_273/A 0.00fF
C44714 INVX1_LOC_24/A NAND2X1_LOC_668/a_36_24# 0.01fF
C44715 NOR2X1_LOC_15/Y INVX1_LOC_270/A 0.65fF
C44716 INVX1_LOC_16/A NOR2X1_LOC_612/Y 0.02fF
C44717 INVX1_LOC_132/A NAND2X1_LOC_74/B 0.10fF
C44718 NOR2X1_LOC_6/B INVX1_LOC_63/A 0.11fF
C44719 NOR2X1_LOC_313/a_36_216# NOR2X1_LOC_56/Y 0.00fF
C44720 NOR2X1_LOC_612/B INVX1_LOC_84/A 0.07fF
C44721 NOR2X1_LOC_759/Y NAND2X1_LOC_792/B 0.07fF
C44722 NOR2X1_LOC_238/Y NOR2X1_LOC_754/A 0.01fF
C44723 INVX1_LOC_286/A NOR2X1_LOC_192/A 0.14fF
C44724 D_INPUT_7 NAND2X1_LOC_3/B 0.04fF
C44725 NOR2X1_LOC_716/B NOR2X1_LOC_327/a_36_216# 0.00fF
C44726 INVX1_LOC_111/Y INVX1_LOC_84/A 0.02fF
C44727 INVX1_LOC_25/A INVX1_LOC_88/A 0.02fF
C44728 INVX1_LOC_22/A NOR2X1_LOC_155/A 0.42fF
C44729 INVX1_LOC_42/Y INVX1_LOC_76/A 0.01fF
C44730 NOR2X1_LOC_326/Y NOR2X1_LOC_729/A 0.02fF
C44731 NOR2X1_LOC_52/B NAND2X1_LOC_773/B 0.02fF
C44732 NOR2X1_LOC_717/B NOR2X1_LOC_729/A 0.03fF
C44733 NOR2X1_LOC_590/A INVX1_LOC_23/Y 0.15fF
C44734 NOR2X1_LOC_360/Y INVX1_LOC_4/A 0.14fF
C44735 NOR2X1_LOC_557/Y NOR2X1_LOC_89/A 0.03fF
C44736 NOR2X1_LOC_65/B NOR2X1_LOC_160/B 1.70fF
C44737 NOR2X1_LOC_388/Y INVX1_LOC_12/A 0.05fF
C44738 NOR2X1_LOC_561/Y NOR2X1_LOC_508/a_36_216# 0.01fF
C44739 INVX1_LOC_36/A INVX1_LOC_273/A 0.17fF
C44740 INVX1_LOC_225/A NAND2X1_LOC_74/B 0.03fF
C44741 NAND2X1_LOC_374/Y NAND2X1_LOC_477/Y 0.11fF
C44742 NOR2X1_LOC_71/Y INVX1_LOC_127/A 0.03fF
C44743 INVX1_LOC_278/A INVX1_LOC_14/A 0.07fF
C44744 NOR2X1_LOC_52/Y NAND2X1_LOC_454/Y 0.16fF
C44745 NOR2X1_LOC_68/A NOR2X1_LOC_685/B 0.03fF
C44746 INVX1_LOC_290/A INVX1_LOC_107/Y 0.11fF
C44747 NOR2X1_LOC_270/Y NAND2X1_LOC_454/Y 0.41fF
C44748 NOR2X1_LOC_15/Y NOR2X1_LOC_109/Y 0.03fF
C44749 NOR2X1_LOC_772/B INVX1_LOC_1/A 0.07fF
C44750 INVX1_LOC_159/A NAND2X1_LOC_470/B 0.07fF
C44751 NOR2X1_LOC_828/A NOR2X1_LOC_729/A 0.18fF
C44752 NOR2X1_LOC_773/Y NOR2X1_LOC_605/A 0.02fF
C44753 NOR2X1_LOC_687/Y NOR2X1_LOC_801/A 0.02fF
C44754 NOR2X1_LOC_541/Y INVX1_LOC_53/A 0.01fF
C44755 VDD INVX1_LOC_126/Y 0.37fF
C44756 NOR2X1_LOC_191/a_36_216# INVX1_LOC_95/Y 0.00fF
C44757 INVX1_LOC_135/A INVX1_LOC_307/A 0.00fF
C44758 INVX1_LOC_179/Y INVX1_LOC_19/A 0.03fF
C44759 INVX1_LOC_232/A NOR2X1_LOC_814/A 0.07fF
C44760 NOR2X1_LOC_468/Y INVX1_LOC_306/Y 0.11fF
C44761 INVX1_LOC_13/Y INVX1_LOC_1/A 0.15fF
C44762 NOR2X1_LOC_749/Y INVX1_LOC_92/A 0.01fF
C44763 INVX1_LOC_135/A NOR2X1_LOC_445/B 0.07fF
C44764 INVX1_LOC_27/A NAND2X1_LOC_218/A 0.03fF
C44765 INVX1_LOC_171/A NOR2X1_LOC_79/Y 0.01fF
C44766 NAND2X1_LOC_208/B INVX1_LOC_23/A 0.01fF
C44767 INVX1_LOC_27/A NOR2X1_LOC_140/A 0.01fF
C44768 INVX1_LOC_217/Y INVX1_LOC_15/A 0.03fF
C44769 NAND2X1_LOC_190/Y NOR2X1_LOC_644/a_36_216# 0.00fF
C44770 NAND2X1_LOC_364/A NAND2X1_LOC_288/B 0.13fF
C44771 NOR2X1_LOC_91/A NOR2X1_LOC_518/a_36_216# 0.01fF
C44772 INVX1_LOC_143/A NOR2X1_LOC_89/A 0.02fF
C44773 NOR2X1_LOC_92/Y NOR2X1_LOC_173/Y 0.03fF
C44774 INVX1_LOC_30/Y INVX1_LOC_63/A 0.02fF
C44775 NOR2X1_LOC_562/B NOR2X1_LOC_357/Y 0.03fF
C44776 NOR2X1_LOC_92/Y NOR2X1_LOC_321/Y 0.07fF
C44777 NOR2X1_LOC_644/A NOR2X1_LOC_600/a_36_216# 0.00fF
C44778 INVX1_LOC_45/A INVX1_LOC_53/A 5.02fF
C44779 INVX1_LOC_25/Y INVX1_LOC_29/A 0.18fF
C44780 NOR2X1_LOC_791/B NAND2X1_LOC_215/A 0.01fF
C44781 INVX1_LOC_28/A NOR2X1_LOC_58/a_36_216# 0.00fF
C44782 INVX1_LOC_303/A INVX1_LOC_116/Y 0.00fF
C44783 INVX1_LOC_290/A INVX1_LOC_272/A 0.00fF
C44784 NOR2X1_LOC_598/B NOR2X1_LOC_274/B 0.17fF
C44785 NOR2X1_LOC_561/Y INVX1_LOC_19/A 0.08fF
C44786 INVX1_LOC_35/A INVX1_LOC_312/Y 0.09fF
C44787 NAND2X1_LOC_9/Y INVX1_LOC_72/A 0.00fF
C44788 NAND2X1_LOC_479/Y INVX1_LOC_12/A 0.07fF
C44789 INVX1_LOC_95/Y NOR2X1_LOC_266/B 0.03fF
C44790 NOR2X1_LOC_516/B NOR2X1_LOC_847/A 0.03fF
C44791 NOR2X1_LOC_852/B INVX1_LOC_26/Y 0.01fF
C44792 NAND2X1_LOC_549/B INVX1_LOC_3/Y 0.02fF
C44793 INVX1_LOC_229/Y NOR2X1_LOC_36/B 0.18fF
C44794 INVX1_LOC_88/A INVX1_LOC_1/A 0.02fF
C44795 NAND2X1_LOC_363/B NAND2X1_LOC_351/A 0.04fF
C44796 NOR2X1_LOC_588/a_36_216# INVX1_LOC_84/A 0.02fF
C44797 INVX1_LOC_21/A INVX1_LOC_230/Y 0.03fF
C44798 NOR2X1_LOC_92/Y NAND2X1_LOC_793/Y 0.08fF
C44799 NOR2X1_LOC_340/a_36_216# INVX1_LOC_280/A 0.01fF
C44800 INVX1_LOC_132/Y NOR2X1_LOC_691/B 0.04fF
C44801 NOR2X1_LOC_860/B NOR2X1_LOC_416/A 0.47fF
C44802 NOR2X1_LOC_601/Y NAND2X1_LOC_472/Y 0.03fF
C44803 INVX1_LOC_143/A INVX1_LOC_104/Y 0.01fF
C44804 NOR2X1_LOC_91/A INVX1_LOC_34/A 1.92fF
C44805 NOR2X1_LOC_703/A INVX1_LOC_220/A 0.01fF
C44806 NAND2X1_LOC_656/A NOR2X1_LOC_717/A 0.10fF
C44807 NAND2X1_LOC_35/Y INVX1_LOC_18/A 0.07fF
C44808 NOR2X1_LOC_796/B NOR2X1_LOC_784/Y 0.00fF
C44809 INVX1_LOC_64/A NOR2X1_LOC_360/Y 0.10fF
C44810 NAND2X1_LOC_218/B NOR2X1_LOC_598/B 0.06fF
C44811 NOR2X1_LOC_6/B NAND2X1_LOC_223/B 0.07fF
C44812 NOR2X1_LOC_332/A NAND2X1_LOC_207/B 0.02fF
C44813 INVX1_LOC_221/Y NAND2X1_LOC_537/Y 0.03fF
C44814 INVX1_LOC_71/A INVX1_LOC_53/A 0.22fF
C44815 NOR2X1_LOC_445/Y NOR2X1_LOC_383/B 0.00fF
C44816 INVX1_LOC_189/A INVX1_LOC_78/A 0.03fF
C44817 INVX1_LOC_35/A NOR2X1_LOC_546/B 0.00fF
C44818 INVX1_LOC_135/A INVX1_LOC_12/A 0.03fF
C44819 NOR2X1_LOC_778/B NOR2X1_LOC_334/Y 0.28fF
C44820 NOR2X1_LOC_708/Y INVX1_LOC_19/A 0.17fF
C44821 INVX1_LOC_233/Y INVX1_LOC_41/Y 0.00fF
C44822 INVX1_LOC_136/A NOR2X1_LOC_186/Y 0.16fF
C44823 NOR2X1_LOC_130/A NOR2X1_LOC_89/A 0.03fF
C44824 NOR2X1_LOC_52/B NOR2X1_LOC_639/Y 0.04fF
C44825 INVX1_LOC_69/Y NOR2X1_LOC_197/B 0.10fF
C44826 NOR2X1_LOC_740/a_36_216# NOR2X1_LOC_740/Y 0.04fF
C44827 INVX1_LOC_60/Y NOR2X1_LOC_39/Y 0.10fF
C44828 INVX1_LOC_34/A INVX1_LOC_23/A 0.23fF
C44829 NOR2X1_LOC_124/B NAND2X1_LOC_215/A 0.10fF
C44830 NOR2X1_LOC_322/Y NAND2X1_LOC_489/Y 0.00fF
C44831 NOR2X1_LOC_227/a_36_216# INVX1_LOC_210/Y 0.00fF
C44832 NOR2X1_LOC_439/a_36_216# NOR2X1_LOC_334/Y 0.01fF
C44833 INVX1_LOC_208/A INVX1_LOC_78/A 0.27fF
C44834 NAND2X1_LOC_656/A NOR2X1_LOC_649/Y 0.10fF
C44835 NAND2X1_LOC_571/Y INVX1_LOC_18/A 0.11fF
C44836 NAND2X1_LOC_35/Y INVX1_LOC_172/A 0.07fF
C44837 INVX1_LOC_136/A NAND2X1_LOC_573/Y 0.10fF
C44838 NOR2X1_LOC_91/A NAND2X1_LOC_231/Y 0.03fF
C44839 NAND2X1_LOC_725/A NOR2X1_LOC_577/Y 0.10fF
C44840 INVX1_LOC_1/A NOR2X1_LOC_500/B 0.10fF
C44841 INVX1_LOC_58/A NAND2X1_LOC_357/B 0.07fF
C44842 INVX1_LOC_255/Y INVX1_LOC_253/A 0.01fF
C44843 INVX1_LOC_36/A NOR2X1_LOC_15/Y 1.64fF
C44844 INVX1_LOC_16/A NOR2X1_LOC_409/B 0.03fF
C44845 INVX1_LOC_96/Y INVX1_LOC_270/A 0.00fF
C44846 VDD NOR2X1_LOC_536/A 1.38fF
C44847 INVX1_LOC_90/A INVX1_LOC_290/Y 0.68fF
C44848 INVX1_LOC_64/A INVX1_LOC_207/A 0.03fF
C44849 INVX1_LOC_8/A NOR2X1_LOC_392/Y -0.02fF
C44850 NAND2X1_LOC_800/A NOR2X1_LOC_536/A 0.00fF
C44851 NOR2X1_LOC_32/B INVX1_LOC_219/Y 0.03fF
C44852 INVX1_LOC_136/A NAND2X1_LOC_724/A 0.07fF
C44853 NOR2X1_LOC_15/Y NOR2X1_LOC_267/A 0.13fF
C44854 NOR2X1_LOC_781/A NOR2X1_LOC_158/Y 0.01fF
C44855 INVX1_LOC_75/A INVX1_LOC_29/A 0.75fF
C44856 NOR2X1_LOC_552/A NOR2X1_LOC_445/B 0.19fF
C44857 INVX1_LOC_224/Y NOR2X1_LOC_78/B 0.70fF
C44858 INVX1_LOC_95/Y INVX1_LOC_46/Y 0.02fF
C44859 NAND2X1_LOC_231/Y INVX1_LOC_23/A 0.03fF
C44860 NOR2X1_LOC_216/Y NOR2X1_LOC_89/A 0.20fF
C44861 NOR2X1_LOC_65/B INVX1_LOC_208/A 0.01fF
C44862 NOR2X1_LOC_455/Y INVX1_LOC_266/Y 0.03fF
C44863 NOR2X1_LOC_2/Y NOR2X1_LOC_1/Y 0.00fF
C44864 NOR2X1_LOC_589/A INVX1_LOC_26/A 0.02fF
C44865 NOR2X1_LOC_264/Y INVX1_LOC_5/A 0.11fF
C44866 VDD NOR2X1_LOC_655/Y 0.37fF
C44867 INVX1_LOC_186/A NOR2X1_LOC_814/A 0.04fF
C44868 NAND2X1_LOC_9/Y NOR2X1_LOC_537/Y 0.03fF
C44869 NOR2X1_LOC_731/A INVX1_LOC_213/A 0.07fF
C44870 NOR2X1_LOC_15/Y NOR2X1_LOC_208/Y 0.03fF
C44871 INVX1_LOC_166/A NOR2X1_LOC_375/Y 0.02fF
C44872 NAND2X1_LOC_213/A NAND2X1_LOC_161/a_36_24# 0.00fF
C44873 INVX1_LOC_35/A NOR2X1_LOC_168/B 0.02fF
C44874 NAND2X1_LOC_9/Y NAND2X1_LOC_338/B 0.09fF
C44875 INVX1_LOC_17/A NAND2X1_LOC_198/B 0.10fF
C44876 VDD NAND2X1_LOC_93/B 2.59fF
C44877 NOR2X1_LOC_689/Y INVX1_LOC_22/A 0.00fF
C44878 INVX1_LOC_224/A INVX1_LOC_24/A 0.03fF
C44879 NOR2X1_LOC_646/A NAND2X1_LOC_215/A -0.03fF
C44880 NOR2X1_LOC_363/Y INVX1_LOC_54/A 0.05fF
C44881 NOR2X1_LOC_45/B NAND2X1_LOC_768/Y 0.03fF
C44882 NOR2X1_LOC_15/Y NOR2X1_LOC_237/Y 0.07fF
C44883 INVX1_LOC_303/A INVX1_LOC_1/A 0.08fF
C44884 NAND2X1_LOC_9/Y NAND2X1_LOC_323/B 0.08fF
C44885 NOR2X1_LOC_160/B NOR2X1_LOC_554/B 0.07fF
C44886 NOR2X1_LOC_748/Y NOR2X1_LOC_748/A 0.13fF
C44887 INVX1_LOC_11/A INVX1_LOC_24/A 0.44fF
C44888 INVX1_LOC_190/Y NAND2X1_LOC_470/B 0.08fF
C44889 NOR2X1_LOC_78/B NAND2X1_LOC_599/a_36_24# 0.00fF
C44890 NOR2X1_LOC_724/Y NOR2X1_LOC_334/Y -0.02fF
C44891 NAND2X1_LOC_288/A INVX1_LOC_76/A 0.10fF
C44892 NAND2X1_LOC_659/B NOR2X1_LOC_649/B 0.01fF
C44893 VDD NAND2X1_LOC_425/Y 2.53fF
C44894 INVX1_LOC_36/A NAND2X1_LOC_355/a_36_24# 0.00fF
C44895 INVX1_LOC_256/A NOR2X1_LOC_191/B 0.06fF
C44896 NOR2X1_LOC_124/A INVX1_LOC_63/A 0.08fF
C44897 INVX1_LOC_35/Y NOR2X1_LOC_290/a_36_216# 0.01fF
C44898 NAND2X1_LOC_447/Y NOR2X1_LOC_814/A 0.12fF
C44899 NOR2X1_LOC_598/B INVX1_LOC_22/A 0.26fF
C44900 NAND2X1_LOC_553/A NAND2X1_LOC_338/B 0.02fF
C44901 NAND2X1_LOC_59/B INVX1_LOC_1/A 0.13fF
C44902 NAND2X1_LOC_123/Y NOR2X1_LOC_334/Y 0.07fF
C44903 INVX1_LOC_136/A INVX1_LOC_170/A 0.11fF
C44904 INVX1_LOC_27/A NOR2X1_LOC_709/A 0.25fF
C44905 NAND2X1_LOC_840/B NOR2X1_LOC_109/Y 0.00fF
C44906 NAND2X1_LOC_725/Y NOR2X1_LOC_298/Y 0.93fF
C44907 NOR2X1_LOC_641/B NAND2X1_LOC_364/A 0.03fF
C44908 NOR2X1_LOC_798/A NOR2X1_LOC_537/Y 0.04fF
C44909 NOR2X1_LOC_321/Y NAND2X1_LOC_477/A 0.46fF
C44910 VDD NOR2X1_LOC_649/B 1.00fF
C44911 INVX1_LOC_37/A NOR2X1_LOC_430/Y 0.01fF
C44912 NOR2X1_LOC_15/Y NOR2X1_LOC_309/Y 0.11fF
C44913 NAND2X1_LOC_642/Y NAND2X1_LOC_74/B 0.14fF
C44914 NAND2X1_LOC_725/A INVX1_LOC_22/A 0.13fF
C44915 NAND2X1_LOC_96/A NAND2X1_LOC_94/a_36_24# 0.02fF
C44916 VDD INVX1_LOC_3/A 0.51fF
C44917 INVX1_LOC_108/A INVX1_LOC_9/A 0.39fF
C44918 INVX1_LOC_5/A INVX1_LOC_316/Y 0.15fF
C44919 INVX1_LOC_255/Y INVX1_LOC_138/Y 0.00fF
C44920 NOR2X1_LOC_331/B INVX1_LOC_92/A 0.08fF
C44921 INVX1_LOC_65/A INVX1_LOC_69/A 0.11fF
C44922 NOR2X1_LOC_798/A NAND2X1_LOC_323/B 0.03fF
C44923 NOR2X1_LOC_751/Y NAND2X1_LOC_364/A 0.06fF
C44924 NOR2X1_LOC_160/B INVX1_LOC_113/Y 0.03fF
C44925 INVX1_LOC_41/A NAND2X1_LOC_793/Y 0.02fF
C44926 NAND2X1_LOC_715/B INVX1_LOC_22/A 0.01fF
C44927 VDD NOR2X1_LOC_661/A 0.33fF
C44928 INVX1_LOC_10/A NAND2X1_LOC_794/a_36_24# 0.01fF
C44929 NOR2X1_LOC_441/Y INVX1_LOC_81/A 0.04fF
C44930 INVX1_LOC_48/A INVX1_LOC_15/A 0.21fF
C44931 INVX1_LOC_76/A INVX1_LOC_19/A 0.09fF
C44932 INVX1_LOC_45/A INVX1_LOC_184/A 0.03fF
C44933 NOR2X1_LOC_791/Y INVX1_LOC_56/Y 0.03fF
C44934 INVX1_LOC_99/Y NOR2X1_LOC_553/B 0.25fF
C44935 INVX1_LOC_35/A NAND2X1_LOC_656/Y 0.08fF
C44936 INVX1_LOC_298/Y INVX1_LOC_75/A 0.02fF
C44937 NOR2X1_LOC_690/A NOR2X1_LOC_371/a_36_216# 0.00fF
C44938 INVX1_LOC_174/A INVX1_LOC_103/Y 0.02fF
C44939 NAND2X1_LOC_569/B INVX1_LOC_234/A 0.41fF
C44940 INVX1_LOC_75/A NOR2X1_LOC_33/Y -0.02fF
C44941 NAND2X1_LOC_477/A NAND2X1_LOC_793/Y 0.03fF
C44942 NOR2X1_LOC_516/B NOR2X1_LOC_655/a_36_216# 0.00fF
C44943 INVX1_LOC_238/A NAND2X1_LOC_736/Y 0.65fF
C44944 NAND2X1_LOC_149/Y NOR2X1_LOC_210/B 0.06fF
C44945 NOR2X1_LOC_636/A INVX1_LOC_30/A 0.05fF
C44946 INVX1_LOC_34/A INVX1_LOC_31/A 0.20fF
C44947 NAND2X1_LOC_193/a_36_24# NAND2X1_LOC_195/Y 0.00fF
C44948 INVX1_LOC_132/A INVX1_LOC_136/A 0.10fF
C44949 INVX1_LOC_223/A INVX1_LOC_33/A 0.04fF
C44950 NOR2X1_LOC_91/A INPUT_0 0.24fF
C44951 INVX1_LOC_11/A INVX1_LOC_143/A 0.09fF
C44952 INPUT_0 NOR2X1_LOC_668/Y 0.01fF
C44953 NOR2X1_LOC_590/A NAND2X1_LOC_116/A 0.10fF
C44954 NOR2X1_LOC_78/B NOR2X1_LOC_103/Y 0.07fF
C44955 NOR2X1_LOC_201/A INPUT_0 0.00fF
C44956 NOR2X1_LOC_209/Y NOR2X1_LOC_307/A 0.01fF
C44957 INVX1_LOC_12/A INVX1_LOC_139/Y 0.04fF
C44958 INVX1_LOC_293/Y NOR2X1_LOC_271/Y 0.00fF
C44959 INVX1_LOC_232/Y NOR2X1_LOC_82/A 1.97fF
C44960 NOR2X1_LOC_481/A INVX1_LOC_136/A 0.06fF
C44961 NAND2X1_LOC_383/a_36_24# INVX1_LOC_282/A 0.00fF
C44962 NAND2X1_LOC_67/a_36_24# NOR2X1_LOC_632/Y 0.00fF
C44963 NOR2X1_LOC_453/Y GATE_479 0.03fF
C44964 INVX1_LOC_133/A NOR2X1_LOC_536/A 0.02fF
C44965 NAND2X1_LOC_84/Y NOR2X1_LOC_262/Y 0.00fF
C44966 INVX1_LOC_238/A INVX1_LOC_282/Y 0.54fF
C44967 NOR2X1_LOC_813/Y INVX1_LOC_12/A 0.09fF
C44968 NOR2X1_LOC_45/B NOR2X1_LOC_36/A 0.02fF
C44969 INVX1_LOC_24/A NOR2X1_LOC_433/A 0.10fF
C44970 NOR2X1_LOC_559/a_36_216# INVX1_LOC_50/Y 0.01fF
C44971 INVX1_LOC_267/Y NAND2X1_LOC_555/Y 0.02fF
C44972 NOR2X1_LOC_272/Y NOR2X1_LOC_71/Y 0.10fF
C44973 INVX1_LOC_17/A INVX1_LOC_53/Y 0.02fF
C44974 INVX1_LOC_136/A INVX1_LOC_225/A 0.24fF
C44975 INVX1_LOC_17/A NOR2X1_LOC_619/A 0.02fF
C44976 NAND2X1_LOC_721/B NAND2X1_LOC_734/B 0.03fF
C44977 NOR2X1_LOC_89/A NAND2X1_LOC_811/B 0.01fF
C44978 NOR2X1_LOC_658/Y NOR2X1_LOC_423/Y 0.02fF
C44979 INPUT_0 INVX1_LOC_23/A 1.18fF
C44980 INVX1_LOC_64/A NOR2X1_LOC_567/B 0.07fF
C44981 INVX1_LOC_24/A NOR2X1_LOC_593/Y 0.08fF
C44982 NAND2X1_LOC_74/B NOR2X1_LOC_271/Y 0.07fF
C44983 INVX1_LOC_59/A D_INPUT_0 0.04fF
C44984 INVX1_LOC_1/A INVX1_LOC_80/A 0.06fF
C44985 NOR2X1_LOC_837/Y NAND2X1_LOC_361/Y 0.03fF
C44986 INVX1_LOC_12/A INVX1_LOC_280/A 0.07fF
C44987 NOR2X1_LOC_56/Y NAND2X1_LOC_470/B 0.14fF
C44988 NOR2X1_LOC_68/A NOR2X1_LOC_180/Y 0.46fF
C44989 INVX1_LOC_300/Y GATE_811 0.05fF
C44990 NOR2X1_LOC_831/B NAND2X1_LOC_475/Y 0.01fF
C44991 NOR2X1_LOC_155/A NAND2X1_LOC_476/Y 0.01fF
C44992 INVX1_LOC_286/A INVX1_LOC_29/Y 0.11fF
C44993 INVX1_LOC_45/A NOR2X1_LOC_78/B 0.21fF
C44994 NOR2X1_LOC_658/Y NOR2X1_LOC_222/Y 0.48fF
C44995 NOR2X1_LOC_454/Y INVX1_LOC_90/A 0.02fF
C44996 INVX1_LOC_17/A INVX1_LOC_145/Y 0.01fF
C44997 NOR2X1_LOC_590/A INVX1_LOC_232/A 0.01fF
C44998 NOR2X1_LOC_405/A NAND2X1_LOC_288/B 0.02fF
C44999 NOR2X1_LOC_78/B NOR2X1_LOC_568/A 0.00fF
C45000 NOR2X1_LOC_372/A INVX1_LOC_22/A 0.32fF
C45001 NOR2X1_LOC_561/Y INVX1_LOC_161/Y 0.10fF
C45002 NOR2X1_LOC_147/B INVX1_LOC_77/A 0.20fF
C45003 INVX1_LOC_24/A NOR2X1_LOC_52/B 0.37fF
C45004 NOR2X1_LOC_742/A INVX1_LOC_50/Y 0.01fF
C45005 NOR2X1_LOC_636/B NOR2X1_LOC_763/Y 0.92fF
C45006 INVX1_LOC_11/A NAND2X1_LOC_783/A 0.24fF
C45007 INVX1_LOC_24/A NAND2X1_LOC_838/Y 1.16fF
C45008 NOR2X1_LOC_746/Y INVX1_LOC_275/Y 0.01fF
C45009 INVX1_LOC_230/Y NOR2X1_LOC_521/Y 0.01fF
C45010 VDD NAND2X1_LOC_470/B 0.62fF
C45011 INVX1_LOC_78/A NAND2X1_LOC_211/Y 0.27fF
C45012 NOR2X1_LOC_392/B INVX1_LOC_77/A 0.17fF
C45013 INVX1_LOC_200/A INVX1_LOC_135/A 0.10fF
C45014 INVX1_LOC_37/A INVX1_LOC_94/Y 0.08fF
C45015 INVX1_LOC_234/A NOR2X1_LOC_530/Y 0.12fF
C45016 INVX1_LOC_11/A NOR2X1_LOC_130/A 0.06fF
C45017 INVX1_LOC_269/A NOR2X1_LOC_788/B 0.05fF
C45018 INVX1_LOC_26/A INVX1_LOC_20/A 0.03fF
C45019 INVX1_LOC_181/Y INVX1_LOC_98/Y 0.04fF
C45020 NAND2X1_LOC_860/A INVX1_LOC_91/A 0.03fF
C45021 NOR2X1_LOC_208/Y INVX1_LOC_96/Y 0.05fF
C45022 INVX1_LOC_33/A INVX1_LOC_149/Y 0.02fF
C45023 INVX1_LOC_13/Y NOR2X1_LOC_188/A 0.03fF
C45024 NOR2X1_LOC_140/A NOR2X1_LOC_19/B 0.00fF
C45025 INVX1_LOC_32/A INVX1_LOC_193/A 0.03fF
C45026 INVX1_LOC_224/Y NOR2X1_LOC_368/Y 0.03fF
C45027 NAND2X1_LOC_243/B INVX1_LOC_284/A 0.01fF
C45028 INVX1_LOC_13/Y NOR2X1_LOC_548/B 0.05fF
C45029 NOR2X1_LOC_516/B NOR2X1_LOC_554/B 0.08fF
C45030 NOR2X1_LOC_324/A INVX1_LOC_23/A 0.01fF
C45031 NOR2X1_LOC_420/Y NOR2X1_LOC_9/Y 0.00fF
C45032 NOR2X1_LOC_303/Y NOR2X1_LOC_352/Y 0.19fF
C45033 NOR2X1_LOC_295/Y INVX1_LOC_294/Y 0.02fF
C45034 NOR2X1_LOC_557/Y NOR2X1_LOC_52/B 0.91fF
C45035 NOR2X1_LOC_78/B INVX1_LOC_71/A 0.14fF
C45036 NOR2X1_LOC_577/Y NAND2X1_LOC_660/A 0.33fF
C45037 NOR2X1_LOC_65/B NAND2X1_LOC_211/Y 0.01fF
C45038 INVX1_LOC_64/A NOR2X1_LOC_269/Y 0.10fF
C45039 NOR2X1_LOC_267/a_36_216# INVX1_LOC_102/Y 0.01fF
C45040 INVX1_LOC_189/A INVX1_LOC_113/Y 0.00fF
C45041 INVX1_LOC_41/Y NAND2X1_LOC_862/A 0.02fF
C45042 NOR2X1_LOC_583/a_36_216# INVX1_LOC_72/A 0.00fF
C45043 INVX1_LOC_49/A INVX1_LOC_196/A 0.15fF
C45044 NOR2X1_LOC_405/A NOR2X1_LOC_405/Y 0.04fF
C45045 NOR2X1_LOC_78/a_36_216# INVX1_LOC_3/Y 0.09fF
C45046 NOR2X1_LOC_448/A INVX1_LOC_295/Y 0.01fF
C45047 NOR2X1_LOC_256/a_36_216# INVX1_LOC_25/Y 0.00fF
C45048 NAND2X1_LOC_341/a_36_24# INVX1_LOC_105/A 0.00fF
C45049 INVX1_LOC_45/A INVX1_LOC_83/A 0.24fF
C45050 INVX1_LOC_37/A INVX1_LOC_296/A 0.20fF
C45051 NOR2X1_LOC_468/Y NOR2X1_LOC_74/A 0.01fF
C45052 INVX1_LOC_2/Y NAND2X1_LOC_215/A 0.14fF
C45053 INVX1_LOC_124/A NOR2X1_LOC_392/B 0.39fF
C45054 NAND2X1_LOC_190/Y NOR2X1_LOC_74/A 0.07fF
C45055 NOR2X1_LOC_276/a_36_216# NOR2X1_LOC_561/Y 0.01fF
C45056 INVX1_LOC_221/A NAND2X1_LOC_534/a_36_24# 0.02fF
C45057 NOR2X1_LOC_443/Y INVX1_LOC_117/A 0.09fF
C45058 NOR2X1_LOC_468/Y NOR2X1_LOC_9/Y 0.07fF
C45059 VDD NOR2X1_LOC_476/B 0.07fF
C45060 INVX1_LOC_135/A INVX1_LOC_217/A 0.01fF
C45061 INVX1_LOC_11/A NOR2X1_LOC_112/B 0.01fF
C45062 NOR2X1_LOC_791/B NOR2X1_LOC_99/B 0.01fF
C45063 NOR2X1_LOC_361/B INVX1_LOC_126/Y 0.06fF
C45064 NOR2X1_LOC_441/Y NOR2X1_LOC_111/Y 0.01fF
C45065 INVX1_LOC_71/A NAND2X1_LOC_392/Y 0.04fF
C45066 NOR2X1_LOC_437/Y NOR2X1_LOC_561/Y 0.10fF
C45067 INVX1_LOC_313/A INVX1_LOC_79/Y 0.01fF
C45068 INVX1_LOC_14/Y NOR2X1_LOC_678/A 0.03fF
C45069 INVX1_LOC_14/A INVX1_LOC_123/A 0.07fF
C45070 INVX1_LOC_186/Y NOR2X1_LOC_833/B 0.01fF
C45071 INVX1_LOC_25/Y INVX1_LOC_8/A 1.79fF
C45072 NAND2X1_LOC_254/Y NAND2X1_LOC_773/B 0.01fF
C45073 NAND2X1_LOC_399/a_36_24# INVX1_LOC_25/Y 0.00fF
C45074 INVX1_LOC_11/Y INVX1_LOC_242/A 0.08fF
C45075 INVX1_LOC_83/A INVX1_LOC_71/A 0.15fF
C45076 NOR2X1_LOC_353/Y NOR2X1_LOC_352/Y 0.00fF
C45077 NAND2X1_LOC_326/A NAND2X1_LOC_655/A 0.03fF
C45078 NAND2X1_LOC_562/B INVX1_LOC_316/Y 0.04fF
C45079 NOR2X1_LOC_68/A NOR2X1_LOC_732/a_36_216# 0.00fF
C45080 NAND2X1_LOC_537/Y INVX1_LOC_91/A 0.01fF
C45081 NAND2X1_LOC_308/Y INVX1_LOC_22/A 0.06fF
C45082 INVX1_LOC_55/Y NOR2X1_LOC_457/B 0.07fF
C45083 NAND2X1_LOC_366/A INVX1_LOC_160/Y 0.00fF
C45084 INVX1_LOC_34/A NAND2X1_LOC_859/Y 0.01fF
C45085 NOR2X1_LOC_553/B NOR2X1_LOC_254/Y 0.01fF
C45086 INVX1_LOC_31/A INPUT_0 0.66fF
C45087 NOR2X1_LOC_177/Y INVX1_LOC_181/A 0.09fF
C45088 INVX1_LOC_305/Y NOR2X1_LOC_168/B 0.14fF
C45089 NOR2X1_LOC_433/A NOR2X1_LOC_130/A 0.10fF
C45090 INVX1_LOC_53/A NOR2X1_LOC_331/B 0.10fF
C45091 NOR2X1_LOC_649/a_36_216# NOR2X1_LOC_332/A 0.01fF
C45092 INVX1_LOC_21/A NOR2X1_LOC_331/a_36_216# 0.02fF
C45093 INVX1_LOC_213/A INVX1_LOC_117/A 0.20fF
C45094 NAND2X1_LOC_53/Y NOR2X1_LOC_45/B 0.01fF
C45095 INVX1_LOC_90/A INVX1_LOC_77/A 0.12fF
C45096 NAND2X1_LOC_757/a_36_24# NOR2X1_LOC_756/Y 0.00fF
C45097 NOR2X1_LOC_709/A INVX1_LOC_137/A 0.02fF
C45098 INVX1_LOC_2/A INVX1_LOC_268/A 0.03fF
C45099 NOR2X1_LOC_389/B INVX1_LOC_77/A 0.03fF
C45100 NOR2X1_LOC_13/Y NOR2X1_LOC_329/B 0.20fF
C45101 INVX1_LOC_17/A NOR2X1_LOC_557/a_36_216# 0.00fF
C45102 INVX1_LOC_25/A NOR2X1_LOC_99/Y 0.08fF
C45103 INVX1_LOC_287/A NOR2X1_LOC_155/A 0.03fF
C45104 NOR2X1_LOC_751/A NAND2X1_LOC_364/A 0.02fF
C45105 INVX1_LOC_18/A INVX1_LOC_144/A 0.07fF
C45106 NAND2X1_LOC_783/A NOR2X1_LOC_52/B 0.06fF
C45107 NOR2X1_LOC_590/A INVX1_LOC_186/A 0.01fF
C45108 NOR2X1_LOC_608/Y NAND2X1_LOC_215/A 0.02fF
C45109 VDD NOR2X1_LOC_348/Y 0.31fF
C45110 NOR2X1_LOC_103/Y NOR2X1_LOC_368/Y 0.00fF
C45111 NOR2X1_LOC_701/Y NAND2X1_LOC_852/Y 0.31fF
C45112 NOR2X1_LOC_778/B NOR2X1_LOC_569/Y 0.07fF
C45113 INVX1_LOC_34/A NAND2X1_LOC_866/B 0.10fF
C45114 INVX1_LOC_304/Y INVX1_LOC_135/A 0.03fF
C45115 NOR2X1_LOC_722/Y INVX1_LOC_6/A 0.01fF
C45116 NOR2X1_LOC_52/B NOR2X1_LOC_130/A 0.09fF
C45117 INVX1_LOC_21/A INVX1_LOC_44/A 0.07fF
C45118 INVX1_LOC_233/A NAND2X1_LOC_444/a_36_24# 0.01fF
C45119 INVX1_LOC_6/A INVX1_LOC_79/Y 0.01fF
C45120 NOR2X1_LOC_67/A NOR2X1_LOC_391/A 0.07fF
C45121 INVX1_LOC_299/A INVX1_LOC_37/A 0.07fF
C45122 NOR2X1_LOC_596/A NOR2X1_LOC_74/A 0.17fF
C45123 NOR2X1_LOC_216/Y NOR2X1_LOC_433/A 0.07fF
C45124 INVX1_LOC_41/A INVX1_LOC_148/A 0.04fF
C45125 INVX1_LOC_85/Y NOR2X1_LOC_727/a_36_216# 0.00fF
C45126 INVX1_LOC_53/A NOR2X1_LOC_592/B 0.01fF
C45127 NOR2X1_LOC_393/Y NAND2X1_LOC_254/Y 0.03fF
C45128 NAND2X1_LOC_348/A INVX1_LOC_77/A 0.07fF
C45129 NOR2X1_LOC_637/Y INVX1_LOC_144/A 0.05fF
C45130 INVX1_LOC_209/Y NOR2X1_LOC_597/Y 0.00fF
C45131 NAND2X1_LOC_347/B INVX1_LOC_117/A 0.00fF
C45132 NOR2X1_LOC_690/A NOR2X1_LOC_497/Y 0.04fF
C45133 INVX1_LOC_84/A NOR2X1_LOC_383/B 0.03fF
C45134 NOR2X1_LOC_170/a_36_216# NOR2X1_LOC_548/B 0.00fF
C45135 INVX1_LOC_161/Y INVX1_LOC_76/A 0.22fF
C45136 INVX1_LOC_149/A INVX1_LOC_171/A 0.03fF
C45137 INVX1_LOC_45/A NOR2X1_LOC_311/Y 0.02fF
C45138 NOR2X1_LOC_742/A NOR2X1_LOC_718/Y 0.03fF
C45139 NOR2X1_LOC_538/B INVX1_LOC_37/A 0.00fF
C45140 INVX1_LOC_57/A INVX1_LOC_27/Y 0.05fF
C45141 NOR2X1_LOC_103/Y INVX1_LOC_46/A 0.12fF
C45142 NOR2X1_LOC_590/A NAND2X1_LOC_447/Y 0.03fF
C45143 INVX1_LOC_124/A INVX1_LOC_90/A 0.02fF
C45144 NOR2X1_LOC_554/B INVX1_LOC_315/Y 0.11fF
C45145 INVX1_LOC_230/Y NOR2X1_LOC_670/Y 0.00fF
C45146 NOR2X1_LOC_1/Y NOR2X1_LOC_36/A 0.07fF
C45147 NOR2X1_LOC_538/B NOR2X1_LOC_231/A 0.04fF
C45148 INVX1_LOC_2/A NOR2X1_LOC_367/a_36_216# 0.00fF
C45149 NOR2X1_LOC_383/Y NOR2X1_LOC_82/Y 0.00fF
C45150 INVX1_LOC_30/Y INVX1_LOC_1/Y 0.11fF
C45151 INVX1_LOC_214/Y INVX1_LOC_135/A 0.05fF
C45152 NOR2X1_LOC_78/B NOR2X1_LOC_123/B 0.07fF
C45153 INVX1_LOC_303/A NOR2X1_LOC_188/A 0.10fF
C45154 INVX1_LOC_256/A VDD 3.45fF
C45155 NOR2X1_LOC_454/Y INVX1_LOC_38/A 0.10fF
C45156 INVX1_LOC_89/A NOR2X1_LOC_520/A 0.00fF
C45157 INVX1_LOC_207/A INVX1_LOC_282/A 0.07fF
C45158 NAND2X1_LOC_218/B INVX1_LOC_201/A 0.03fF
C45159 INVX1_LOC_17/A INVX1_LOC_77/Y 0.07fF
C45160 INVX1_LOC_21/A NOR2X1_LOC_641/Y 0.00fF
C45161 NOR2X1_LOC_318/A NOR2X1_LOC_831/Y 0.07fF
C45162 INVX1_LOC_303/A NOR2X1_LOC_548/B 0.10fF
C45163 INVX1_LOC_75/A INVX1_LOC_8/A 0.07fF
C45164 INVX1_LOC_130/Y NOR2X1_LOC_269/Y 0.00fF
C45165 INVX1_LOC_136/A NAND2X1_LOC_642/Y 0.29fF
C45166 INVX1_LOC_103/A INVX1_LOC_202/Y 0.01fF
C45167 NOR2X1_LOC_361/B NOR2X1_LOC_536/A 0.03fF
C45168 NOR2X1_LOC_332/A INVX1_LOC_316/Y 0.01fF
C45169 NOR2X1_LOC_658/Y NOR2X1_LOC_69/A 0.01fF
C45170 INVX1_LOC_222/Y NOR2X1_LOC_640/Y 0.04fF
C45171 NOR2X1_LOC_19/B NOR2X1_LOC_709/A 0.01fF
C45172 INVX1_LOC_13/A NOR2X1_LOC_719/B 0.03fF
C45173 NOR2X1_LOC_216/Y NOR2X1_LOC_52/B 0.09fF
C45174 NOR2X1_LOC_798/A NOR2X1_LOC_79/a_36_216# 0.00fF
C45175 NAND2X1_LOC_860/A INVX1_LOC_203/A 0.03fF
C45176 NOR2X1_LOC_657/Y NAND2X1_LOC_469/B 0.03fF
C45177 NAND2X1_LOC_53/Y INVX1_LOC_281/A 0.08fF
C45178 NAND2X1_LOC_231/Y NAND2X1_LOC_807/Y 0.39fF
C45179 NOR2X1_LOC_295/Y NOR2X1_LOC_74/A 0.01fF
C45180 INVX1_LOC_229/Y NAND2X1_LOC_863/a_36_24# 0.01fF
C45181 D_GATE_222 INVX1_LOC_295/A -0.01fF
C45182 NAND2X1_LOC_656/Y NOR2X1_LOC_188/Y 0.14fF
C45183 INVX1_LOC_178/A NOR2X1_LOC_510/B 0.06fF
C45184 NOR2X1_LOC_220/A NOR2X1_LOC_356/A 0.10fF
C45185 NOR2X1_LOC_606/Y VDD 0.39fF
C45186 NOR2X1_LOC_598/B INVX1_LOC_186/Y 0.03fF
C45187 INVX1_LOC_34/A INVX1_LOC_6/A 0.63fF
C45188 INVX1_LOC_45/A INVX1_LOC_46/A 0.13fF
C45189 NOR2X1_LOC_791/Y NOR2X1_LOC_179/a_36_216# 0.00fF
C45190 INVX1_LOC_89/A NOR2X1_LOC_748/Y 0.14fF
C45191 NOR2X1_LOC_773/Y NAND2X1_LOC_850/A 0.01fF
C45192 NOR2X1_LOC_78/B INVX1_LOC_102/Y 2.49fF
C45193 NOR2X1_LOC_568/A INVX1_LOC_46/A 1.31fF
C45194 INVX1_LOC_15/Y NOR2X1_LOC_19/Y 0.25fF
C45195 NOR2X1_LOC_441/Y NOR2X1_LOC_363/Y 0.05fF
C45196 NOR2X1_LOC_751/Y NOR2X1_LOC_857/A 0.01fF
C45197 NAND2X1_LOC_141/a_36_24# NAND2X1_LOC_141/Y 0.02fF
C45198 INVX1_LOC_149/A INVX1_LOC_222/A 0.00fF
C45199 INVX1_LOC_5/A NOR2X1_LOC_662/A 0.07fF
C45200 NAND2X1_LOC_796/B INVX1_LOC_285/A -0.03fF
C45201 INVX1_LOC_135/A NAND2X1_LOC_808/A 0.10fF
C45202 NOR2X1_LOC_356/A NOR2X1_LOC_548/Y 0.09fF
C45203 NAND2X1_LOC_796/B INVX1_LOC_265/Y 0.00fF
C45204 INVX1_LOC_26/A INVX1_LOC_4/A 0.06fF
C45205 INPUT_3 NOR2X1_LOC_54/a_36_216# 0.00fF
C45206 INVX1_LOC_103/A INVX1_LOC_180/Y 0.03fF
C45207 INVX1_LOC_90/A NAND2X1_LOC_796/Y 0.01fF
C45208 NAND2X1_LOC_627/a_36_24# INVX1_LOC_284/A 0.00fF
C45209 NAND2X1_LOC_462/B INVX1_LOC_175/Y 0.04fF
C45210 INVX1_LOC_57/A NOR2X1_LOC_462/a_36_216# 0.00fF
C45211 NAND2X1_LOC_560/A INVX1_LOC_22/A 0.07fF
C45212 NOR2X1_LOC_220/A NOR2X1_LOC_74/A 0.05fF
C45213 INVX1_LOC_209/A NOR2X1_LOC_387/A 0.01fF
C45214 NAND2X1_LOC_231/Y INVX1_LOC_6/A 0.01fF
C45215 NOR2X1_LOC_781/Y VDD 0.12fF
C45216 NOR2X1_LOC_383/B INVX1_LOC_15/A 0.33fF
C45217 NOR2X1_LOC_763/A INVX1_LOC_84/A 0.01fF
C45218 NOR2X1_LOC_34/B INVX1_LOC_19/A 0.03fF
C45219 INVX1_LOC_71/A INVX1_LOC_46/A 0.37fF
C45220 INVX1_LOC_11/A NOR2X1_LOC_197/B 0.01fF
C45221 INVX1_LOC_89/A INVX1_LOC_65/Y 0.01fF
C45222 NAND2X1_LOC_149/Y NOR2X1_LOC_257/Y 0.03fF
C45223 INVX1_LOC_102/Y NAND2X1_LOC_392/Y 0.00fF
C45224 NAND2X1_LOC_551/A NOR2X1_LOC_76/A 0.03fF
C45225 NOR2X1_LOC_516/B INVX1_LOC_158/Y 0.37fF
C45226 INVX1_LOC_89/A D_GATE_366 0.03fF
C45227 INVX1_LOC_217/A INVX1_LOC_280/A 0.00fF
C45228 INVX1_LOC_2/A NOR2X1_LOC_588/A 0.01fF
C45229 NOR2X1_LOC_548/Y NOR2X1_LOC_74/A 0.03fF
C45230 INVX1_LOC_85/A NOR2X1_LOC_486/Y 0.10fF
C45231 NOR2X1_LOC_361/B INVX1_LOC_3/A 2.03fF
C45232 INPUT_6 D_INPUT_5 3.03fF
C45233 NOR2X1_LOC_15/Y INVX1_LOC_63/A 0.10fF
C45234 NAND2X1_LOC_549/Y INVX1_LOC_3/Y 0.02fF
C45235 NAND2X1_LOC_316/a_36_24# NAND2X1_LOC_287/B 0.00fF
C45236 INVX1_LOC_271/A NOR2X1_LOC_334/Y 0.06fF
C45237 INVX1_LOC_161/A NAND2X1_LOC_810/B 0.12fF
C45238 NOR2X1_LOC_91/A INVX1_LOC_183/A 0.01fF
C45239 INVX1_LOC_2/A INVX1_LOC_95/Y 0.10fF
C45240 INVX1_LOC_181/Y NOR2X1_LOC_709/B 0.00fF
C45241 INVX1_LOC_284/A NOR2X1_LOC_384/A 0.02fF
C45242 INVX1_LOC_31/A NAND2X1_LOC_240/a_36_24# 0.00fF
C45243 INVX1_LOC_226/Y NOR2X1_LOC_45/B 0.03fF
C45244 NOR2X1_LOC_52/B NOR2X1_LOC_280/Y 0.03fF
C45245 NOR2X1_LOC_226/A INVX1_LOC_95/Y 0.07fF
C45246 INVX1_LOC_77/A INVX1_LOC_38/A 1.35fF
C45247 INVX1_LOC_30/A NOR2X1_LOC_831/B 0.03fF
C45248 INVX1_LOC_35/A INVX1_LOC_128/Y 0.69fF
C45249 INVX1_LOC_53/A NAND2X1_LOC_467/a_36_24# 0.00fF
C45250 NOR2X1_LOC_142/Y NOR2X1_LOC_363/Y 0.10fF
C45251 INVX1_LOC_251/A INVX1_LOC_306/Y 0.11fF
C45252 INVX1_LOC_57/Y NOR2X1_LOC_88/Y 0.26fF
C45253 INVX1_LOC_232/Y INVX1_LOC_59/Y 0.01fF
C45254 NOR2X1_LOC_315/Y INVX1_LOC_37/A 0.03fF
C45255 NOR2X1_LOC_132/Y NOR2X1_LOC_536/A 0.01fF
C45256 INVX1_LOC_18/A NOR2X1_LOC_155/A 0.10fF
C45257 INVX1_LOC_53/A NOR2X1_LOC_449/A 0.06fF
C45258 INVX1_LOC_2/A NOR2X1_LOC_305/Y 0.43fF
C45259 NOR2X1_LOC_181/Y NAND2X1_LOC_472/Y 0.03fF
C45260 INVX1_LOC_256/A INVX1_LOC_133/A 0.12fF
C45261 NOR2X1_LOC_655/B INVX1_LOC_2/Y 0.03fF
C45262 NOR2X1_LOC_226/A NOR2X1_LOC_305/Y 0.10fF
C45263 NOR2X1_LOC_45/B INVX1_LOC_10/A 0.14fF
C45264 NOR2X1_LOC_598/B NOR2X1_LOC_843/B 0.08fF
C45265 INVX1_LOC_205/A NAND2X1_LOC_574/A 0.02fF
C45266 INPUT_0 NAND2X1_LOC_807/Y 0.11fF
C45267 INVX1_LOC_57/Y INVX1_LOC_84/A 0.74fF
C45268 INVX1_LOC_53/A NOR2X1_LOC_106/a_36_216# 0.01fF
C45269 INVX1_LOC_64/A INVX1_LOC_26/A 0.06fF
C45270 NOR2X1_LOC_557/Y NOR2X1_LOC_675/a_36_216# 0.04fF
C45271 NAND2X1_LOC_683/a_36_24# NAND2X1_LOC_655/A 0.00fF
C45272 NOR2X1_LOC_392/B INVX1_LOC_9/A 0.01fF
C45273 INVX1_LOC_27/A NOR2X1_LOC_334/Y 0.07fF
C45274 NOR2X1_LOC_65/B NAND2X1_LOC_78/a_36_24# 0.00fF
C45275 NAND2X1_LOC_9/Y INVX1_LOC_224/Y 0.73fF
C45276 INVX1_LOC_53/A NOR2X1_LOC_493/A 0.02fF
C45277 INVX1_LOC_227/A NAND2X1_LOC_447/Y 0.10fF
C45278 INVX1_LOC_157/A NOR2X1_LOC_56/Y 0.02fF
C45279 INVX1_LOC_85/Y INVX1_LOC_91/A 0.03fF
C45280 INVX1_LOC_89/A NOR2X1_LOC_746/Y 0.32fF
C45281 INVX1_LOC_131/A INVX1_LOC_6/A 0.07fF
C45282 INVX1_LOC_58/A NAND2X1_LOC_549/Y 0.02fF
C45283 NOR2X1_LOC_470/A INVX1_LOC_115/A 0.10fF
C45284 INVX1_LOC_36/A INVX1_LOC_49/Y 0.19fF
C45285 NOR2X1_LOC_388/Y INVX1_LOC_92/A 0.07fF
C45286 INVX1_LOC_268/Y INVX1_LOC_37/A 0.01fF
C45287 INVX1_LOC_162/A NOR2X1_LOC_743/Y 0.14fF
C45288 INVX1_LOC_280/Y NOR2X1_LOC_536/A 5.61fF
C45289 NOR2X1_LOC_226/A NAND2X1_LOC_446/a_36_24# 0.00fF
C45290 INVX1_LOC_243/Y INVX1_LOC_5/A 0.04fF
C45291 NOR2X1_LOC_285/A NOR2X1_LOC_285/Y 0.00fF
C45292 NOR2X1_LOC_593/Y NOR2X1_LOC_197/B 0.27fF
C45293 INVX1_LOC_164/A INVX1_LOC_20/A 0.32fF
C45294 INVX1_LOC_286/Y NOR2X1_LOC_89/A 0.07fF
C45295 NAND2X1_LOC_711/Y INVX1_LOC_102/A 0.07fF
C45296 NOR2X1_LOC_78/B NOR2X1_LOC_331/B 0.14fF
C45297 INVX1_LOC_64/A NOR2X1_LOC_255/Y 0.12fF
C45298 NAND2X1_LOC_552/A INVX1_LOC_57/A 0.06fF
C45299 NOR2X1_LOC_130/A INVX1_LOC_74/A 0.14fF
C45300 NOR2X1_LOC_440/Y VDD 0.96fF
C45301 INVX1_LOC_224/Y NAND2X1_LOC_553/A 0.03fF
C45302 INVX1_LOC_5/A INVX1_LOC_57/A 0.11fF
C45303 INVX1_LOC_186/A NOR2X1_LOC_703/A 0.05fF
C45304 NOR2X1_LOC_669/a_36_216# NAND2X1_LOC_175/Y 0.01fF
C45305 INVX1_LOC_58/A NOR2X1_LOC_406/a_36_216# 0.00fF
C45306 INVX1_LOC_215/A NOR2X1_LOC_111/A 0.01fF
C45307 NOR2X1_LOC_810/A VDD 0.12fF
C45308 INVX1_LOC_35/A NOR2X1_LOC_717/A 0.03fF
C45309 INVX1_LOC_299/A NAND2X1_LOC_72/B 0.07fF
C45310 INVX1_LOC_233/A NAND2X1_LOC_793/B 0.07fF
C45311 INVX1_LOC_233/Y NOR2X1_LOC_754/Y 0.29fF
C45312 NOR2X1_LOC_860/B INVX1_LOC_63/A 0.07fF
C45313 INVX1_LOC_122/Y NOR2X1_LOC_340/A 0.64fF
C45314 NAND2X1_LOC_214/B NAND2X1_LOC_607/a_36_24# 0.00fF
C45315 INPUT_0 INVX1_LOC_6/A 1.49fF
C45316 INVX1_LOC_95/Y INPUT_1 0.08fF
C45317 NOR2X1_LOC_554/B NAND2X1_LOC_207/B 0.05fF
C45318 INVX1_LOC_157/A VDD -0.00fF
C45319 NAND2X1_LOC_69/a_36_24# NAND2X1_LOC_363/B 0.01fF
C45320 INVX1_LOC_177/A NAND2X1_LOC_93/B 0.03fF
C45321 NAND2X1_LOC_477/A NAND2X1_LOC_798/B 0.03fF
C45322 INVX1_LOC_88/A NOR2X1_LOC_338/a_36_216# 0.00fF
C45323 INVX1_LOC_100/Y NOR2X1_LOC_74/A 0.02fF
C45324 NAND2X1_LOC_706/Y NOR2X1_LOC_693/Y 0.06fF
C45325 NOR2X1_LOC_123/B INVX1_LOC_46/A 0.14fF
C45326 INVX1_LOC_178/A INVX1_LOC_57/A 0.03fF
C45327 NOR2X1_LOC_795/Y NOR2X1_LOC_445/B 1.23fF
C45328 NOR2X1_LOC_274/Y INVX1_LOC_19/A 0.04fF
C45329 INVX1_LOC_299/A NOR2X1_LOC_863/B 0.02fF
C45330 NOR2X1_LOC_824/A NAND2X1_LOC_464/B 0.09fF
C45331 NOR2X1_LOC_709/A NOR2X1_LOC_216/B 0.10fF
C45332 INVX1_LOC_18/A NOR2X1_LOC_833/B 0.06fF
C45333 INVX1_LOC_30/A NAND2X1_LOC_430/B 0.02fF
C45334 NOR2X1_LOC_764/Y VDD 0.18fF
C45335 NAND2X1_LOC_364/Y NOR2X1_LOC_691/B 0.10fF
C45336 NOR2X1_LOC_214/B NAND2X1_LOC_39/Y 0.01fF
C45337 NOR2X1_LOC_844/A NOR2X1_LOC_243/B 0.05fF
C45338 NAND2X1_LOC_855/Y INVX1_LOC_11/Y 0.01fF
C45339 NAND2X1_LOC_218/B INVX1_LOC_29/A 0.01fF
C45340 NAND2X1_LOC_349/B INVX1_LOC_118/Y 0.04fF
C45341 INVX1_LOC_166/A INVX1_LOC_163/A 1.17fF
C45342 NAND2X1_LOC_206/a_36_24# INVX1_LOC_15/A 0.00fF
C45343 INVX1_LOC_104/A INVX1_LOC_220/A 0.03fF
C45344 INVX1_LOC_69/Y NOR2X1_LOC_337/Y 0.02fF
C45345 NAND2X1_LOC_573/A NOR2X1_LOC_536/A 0.15fF
C45346 INVX1_LOC_48/A INVX1_LOC_123/A 1.30fF
C45347 NAND2X1_LOC_508/A INVX1_LOC_36/Y 0.13fF
C45348 NOR2X1_LOC_151/Y NOR2X1_LOC_833/Y 0.00fF
C45349 INVX1_LOC_24/A NAND2X1_LOC_254/Y 0.39fF
C45350 D_INPUT_0 NOR2X1_LOC_98/B 0.02fF
C45351 VDD INVX1_LOC_169/A -0.00fF
C45352 NOR2X1_LOC_577/Y INVX1_LOC_29/A 0.07fF
C45353 INVX1_LOC_83/A NOR2X1_LOC_331/B 0.10fF
C45354 NOR2X1_LOC_82/A NOR2X1_LOC_72/Y 0.00fF
C45355 NOR2X1_LOC_86/A NAND2X1_LOC_243/Y 0.02fF
C45356 NOR2X1_LOC_457/B INVX1_LOC_32/A 0.07fF
C45357 NOR2X1_LOC_614/Y NOR2X1_LOC_445/B 0.02fF
C45358 D_INPUT_1 INVX1_LOC_14/A 0.20fF
C45359 NOR2X1_LOC_791/A NOR2X1_LOC_38/B 0.01fF
C45360 NAND2X1_LOC_479/Y INVX1_LOC_92/A 0.00fF
C45361 NOR2X1_LOC_389/A NAND2X1_LOC_425/a_36_24# 0.00fF
C45362 INVX1_LOC_50/A NOR2X1_LOC_218/A 0.06fF
C45363 NOR2X1_LOC_8/a_36_216# INVX1_LOC_3/Y 0.02fF
C45364 NOR2X1_LOC_317/A NOR2X1_LOC_855/A 0.02fF
C45365 NOR2X1_LOC_97/A INVX1_LOC_176/A 0.02fF
C45366 INVX1_LOC_11/A NOR2X1_LOC_260/Y 0.04fF
C45367 NOR2X1_LOC_355/A INVX1_LOC_54/A 0.05fF
C45368 NAND2X1_LOC_337/B INVX1_LOC_57/A 0.01fF
C45369 INVX1_LOC_33/A INVX1_LOC_290/Y 0.07fF
C45370 NOR2X1_LOC_816/A INVX1_LOC_57/A 0.07fF
C45371 NOR2X1_LOC_50/a_36_216# D_INPUT_5 0.00fF
C45372 NOR2X1_LOC_348/B INVX1_LOC_29/A 0.17fF
C45373 INVX1_LOC_90/A INVX1_LOC_9/A 0.77fF
C45374 INVX1_LOC_25/A INVX1_LOC_150/Y 0.00fF
C45375 INVX1_LOC_225/Y INVX1_LOC_23/A 0.01fF
C45376 NAND2X1_LOC_9/Y NOR2X1_LOC_103/Y 0.03fF
C45377 NAND2X1_LOC_725/A NOR2X1_LOC_536/Y 0.12fF
C45378 NAND2X1_LOC_198/B INVX1_LOC_94/Y 0.10fF
C45379 NOR2X1_LOC_773/Y NOR2X1_LOC_662/A 0.07fF
C45380 NOR2X1_LOC_315/Y NOR2X1_LOC_178/a_36_216# 0.00fF
C45381 NAND2X1_LOC_170/A INVX1_LOC_84/A 0.03fF
C45382 INVX1_LOC_73/A INVX1_LOC_66/Y 0.03fF
C45383 NOR2X1_LOC_561/Y NOR2X1_LOC_841/A 0.03fF
C45384 INVX1_LOC_69/Y VDD 1.61fF
C45385 INVX1_LOC_83/A NOR2X1_LOC_592/B 0.03fF
C45386 INVX1_LOC_163/A NAND2X1_LOC_398/a_36_24# 0.00fF
C45387 NOR2X1_LOC_721/A NAND2X1_LOC_207/B 0.03fF
C45388 INVX1_LOC_41/A INVX1_LOC_47/Y 0.49fF
C45389 INVX1_LOC_14/A NOR2X1_LOC_652/Y 0.11fF
C45390 NOR2X1_LOC_738/Y INVX1_LOC_213/A 0.06fF
C45391 NOR2X1_LOC_346/B INVX1_LOC_29/A 0.03fF
C45392 NOR2X1_LOC_481/A NAND2X1_LOC_647/B 0.25fF
C45393 NAND2X1_LOC_593/a_36_24# INVX1_LOC_78/A 0.00fF
C45394 INVX1_LOC_178/A NOR2X1_LOC_475/A 0.05fF
C45395 NAND2X1_LOC_553/A NOR2X1_LOC_103/Y 0.01fF
C45396 NAND2X1_LOC_348/A INVX1_LOC_9/A 0.10fF
C45397 INVX1_LOC_49/A INVX1_LOC_271/Y 0.07fF
C45398 INVX1_LOC_315/A INVX1_LOC_4/A 0.32fF
C45399 INVX1_LOC_89/A INVX1_LOC_123/Y 0.10fF
C45400 INVX1_LOC_77/A INVX1_LOC_18/Y 0.07fF
C45401 INVX1_LOC_95/A INVX1_LOC_126/A 0.03fF
C45402 NAND2X1_LOC_9/Y INVX1_LOC_45/A 0.06fF
C45403 NAND2X1_LOC_143/a_36_24# NOR2X1_LOC_649/B 0.00fF
C45404 NOR2X1_LOC_790/B INVX1_LOC_30/A 0.10fF
C45405 INVX1_LOC_155/A INVX1_LOC_78/A 0.03fF
C45406 NOR2X1_LOC_414/a_36_216# NOR2X1_LOC_392/Y 0.00fF
C45407 INVX1_LOC_22/A INVX1_LOC_29/A 0.17fF
C45408 NAND2X1_LOC_763/B NAND2X1_LOC_763/a_36_24# 0.08fF
C45409 NOR2X1_LOC_510/Y INVX1_LOC_256/A 0.10fF
C45410 INVX1_LOC_298/Y NOR2X1_LOC_577/Y 0.07fF
C45411 INVX1_LOC_131/A INVX1_LOC_131/Y 0.09fF
C45412 NAND2X1_LOC_860/A NOR2X1_LOC_372/Y 0.10fF
C45413 NOR2X1_LOC_750/Y INVX1_LOC_136/A 0.01fF
C45414 INVX1_LOC_233/A INVX1_LOC_45/A 0.08fF
C45415 INVX1_LOC_1/A NOR2X1_LOC_271/B 0.03fF
C45416 NAND2X1_LOC_833/Y NAND2X1_LOC_175/Y 0.01fF
C45417 NAND2X1_LOC_796/B NAND2X1_LOC_803/B 0.07fF
C45418 INVX1_LOC_57/Y INVX1_LOC_278/A 0.09fF
C45419 INVX1_LOC_88/A NAND2X1_LOC_326/A 0.01fF
C45420 NOR2X1_LOC_202/Y INVX1_LOC_92/A 0.03fF
C45421 NOR2X1_LOC_264/Y INVX1_LOC_78/A 0.07fF
C45422 NOR2X1_LOC_598/B INVX1_LOC_18/A 2.50fF
C45423 INVX1_LOC_149/A INVX1_LOC_4/A 0.07fF
C45424 NOR2X1_LOC_310/Y INVX1_LOC_4/Y 0.01fF
C45425 NOR2X1_LOC_793/Y INVX1_LOC_269/A 0.29fF
C45426 INVX1_LOC_13/A NOR2X1_LOC_14/a_36_216# 0.00fF
C45427 NAND2X1_LOC_565/B NAND2X1_LOC_254/Y 0.01fF
C45428 INVX1_LOC_1/A NOR2X1_LOC_740/Y 0.00fF
C45429 NOR2X1_LOC_329/B NOR2X1_LOC_697/Y 0.03fF
C45430 NOR2X1_LOC_471/Y NAND2X1_LOC_149/Y 0.09fF
C45431 INVX1_LOC_206/A NOR2X1_LOC_334/Y 0.02fF
C45432 NAND2X1_LOC_796/B NOR2X1_LOC_590/A 0.00fF
C45433 NOR2X1_LOC_65/B INVX1_LOC_155/A 0.02fF
C45434 INVX1_LOC_166/A INVX1_LOC_203/Y 0.04fF
C45435 NOR2X1_LOC_470/B INVX1_LOC_11/A 0.01fF
C45436 NOR2X1_LOC_679/Y NOR2X1_LOC_92/Y 0.02fF
C45437 NAND2X1_LOC_169/Y INVX1_LOC_30/A 0.01fF
C45438 NOR2X1_LOC_381/Y NOR2X1_LOC_82/A 0.06fF
C45439 INVX1_LOC_235/Y NAND2X1_LOC_555/Y 0.18fF
C45440 NOR2X1_LOC_91/A NAND2X1_LOC_811/Y 0.03fF
C45441 INVX1_LOC_285/Y NAND2X1_LOC_93/B 4.22fF
C45442 INVX1_LOC_45/A NOR2X1_LOC_798/A 0.03fF
C45443 NAND2X1_LOC_728/Y NAND2X1_LOC_725/A 0.10fF
C45444 INVX1_LOC_2/A INVX1_LOC_271/Y 0.07fF
C45445 NAND2X1_LOC_79/Y NOR2X1_LOC_392/Y 0.01fF
C45446 INPUT_0 NAND2X1_LOC_810/B 0.12fF
C45447 NOR2X1_LOC_211/Y NOR2X1_LOC_360/Y 0.03fF
C45448 NAND2X1_LOC_9/Y INVX1_LOC_71/A 0.01fF
C45449 INVX1_LOC_256/A NOR2X1_LOC_361/B 0.19fF
C45450 INVX1_LOC_72/A NOR2X1_LOC_674/Y 0.15fF
C45451 NAND2X1_LOC_714/B INVX1_LOC_141/Y 0.35fF
C45452 NOR2X1_LOC_798/A NOR2X1_LOC_568/A 0.00fF
C45453 INVX1_LOC_35/A NOR2X1_LOC_13/Y 0.03fF
C45454 INVX1_LOC_34/A INVX1_LOC_270/A 0.11fF
C45455 INVX1_LOC_233/A INVX1_LOC_71/A 0.10fF
C45456 INVX1_LOC_47/A NAND2X1_LOC_63/Y 0.09fF
C45457 NAND2X1_LOC_849/B NOR2X1_LOC_670/a_36_216# 0.01fF
C45458 NAND2X1_LOC_711/B NAND2X1_LOC_725/A 0.05fF
C45459 NOR2X1_LOC_679/Y NAND2X1_LOC_568/A 0.25fF
C45460 INVX1_LOC_140/A NOR2X1_LOC_662/A 0.02fF
C45461 NOR2X1_LOC_130/A NAND2X1_LOC_254/Y 0.03fF
C45462 INVX1_LOC_34/A NOR2X1_LOC_416/A 0.16fF
C45463 NAND2X1_LOC_562/B INVX1_LOC_57/A 0.01fF
C45464 INVX1_LOC_95/Y INVX1_LOC_118/A 0.10fF
C45465 NOR2X1_LOC_388/Y INVX1_LOC_53/A 0.10fF
C45466 NOR2X1_LOC_719/B INVX1_LOC_32/A 0.05fF
C45467 INVX1_LOC_53/Y INVX1_LOC_94/Y 0.10fF
C45468 NAND2X1_LOC_850/Y INVX1_LOC_26/A 0.21fF
C45469 NOR2X1_LOC_536/A NAND2X1_LOC_267/B 0.02fF
C45470 NAND2X1_LOC_96/A INVX1_LOC_37/A 0.07fF
C45471 NOR2X1_LOC_78/A NOR2X1_LOC_364/A 0.16fF
C45472 NOR2X1_LOC_798/A INVX1_LOC_71/A 0.03fF
C45473 INVX1_LOC_50/A NOR2X1_LOC_822/Y 0.01fF
C45474 INVX1_LOC_11/A INVX1_LOC_286/Y 0.01fF
C45475 INVX1_LOC_90/A NOR2X1_LOC_861/Y 0.17fF
C45476 NOR2X1_LOC_331/B INVX1_LOC_46/A 0.15fF
C45477 INVX1_LOC_21/A NAND2X1_LOC_515/a_36_24# 0.00fF
C45478 NAND2X1_LOC_740/Y NAND2X1_LOC_740/A 0.10fF
C45479 INVX1_LOC_266/Y INVX1_LOC_23/A 0.00fF
C45480 INVX1_LOC_124/Y NAND2X1_LOC_396/a_36_24# 0.01fF
C45481 INVX1_LOC_30/Y INVX1_LOC_87/A 0.07fF
C45482 NOR2X1_LOC_137/B NAND2X1_LOC_93/B 0.11fF
C45483 NOR2X1_LOC_76/A INVX1_LOC_32/A 0.10fF
C45484 INVX1_LOC_279/Y NOR2X1_LOC_160/B 0.01fF
C45485 D_INPUT_0 NOR2X1_LOC_38/B 0.19fF
C45486 D_GATE_741 INVX1_LOC_30/A 0.02fF
C45487 INVX1_LOC_247/A INVX1_LOC_307/A 0.01fF
C45488 NOR2X1_LOC_111/A NOR2X1_LOC_602/B 0.01fF
C45489 INVX1_LOC_145/Y INVX1_LOC_94/Y 0.01fF
C45490 NOR2X1_LOC_78/A INVX1_LOC_285/A 0.07fF
C45491 INVX1_LOC_101/Y NOR2X1_LOC_609/A 0.12fF
C45492 NOR2X1_LOC_773/Y INVX1_LOC_57/A 0.15fF
C45493 INPUT_0 NOR2X1_LOC_633/A 0.03fF
C45494 NOR2X1_LOC_235/Y INVX1_LOC_20/A 0.01fF
C45495 INVX1_LOC_22/A NOR2X1_LOC_318/a_36_216# 0.02fF
C45496 NAND2X1_LOC_860/A NAND2X1_LOC_374/Y 0.12fF
C45497 NOR2X1_LOC_111/A INVX1_LOC_54/A 0.07fF
C45498 NOR2X1_LOC_78/A NOR2X1_LOC_814/A 0.16fF
C45499 INVX1_LOC_100/A INVX1_LOC_29/A 0.01fF
C45500 NOR2X1_LOC_721/Y NOR2X1_LOC_89/A 0.06fF
C45501 INVX1_LOC_36/A INVX1_LOC_161/A 0.03fF
C45502 INVX1_LOC_11/A INVX1_LOC_159/A 0.19fF
C45503 INVX1_LOC_14/A D_INPUT_2 0.07fF
C45504 NAND2X1_LOC_348/A NOR2X1_LOC_861/Y 0.74fF
C45505 NOR2X1_LOC_590/A NOR2X1_LOC_239/a_36_216# 0.00fF
C45506 NAND2X1_LOC_784/a_36_24# NAND2X1_LOC_325/Y -0.00fF
C45507 INVX1_LOC_316/A NOR2X1_LOC_649/B 0.42fF
C45508 NOR2X1_LOC_454/Y INVX1_LOC_33/A 0.07fF
C45509 INVX1_LOC_35/A INVX1_LOC_256/Y 0.03fF
C45510 INVX1_LOC_139/Y INVX1_LOC_92/A 0.04fF
C45511 NOR2X1_LOC_491/Y INVX1_LOC_46/A 0.37fF
C45512 INVX1_LOC_316/A INVX1_LOC_3/A 0.46fF
C45513 INVX1_LOC_81/Y INVX1_LOC_30/A 0.00fF
C45514 NOR2X1_LOC_841/A INVX1_LOC_76/A 0.10fF
C45515 INVX1_LOC_38/A INVX1_LOC_9/A 18.14fF
C45516 NAND2X1_LOC_231/Y NOR2X1_LOC_109/Y 1.43fF
C45517 INVX1_LOC_11/A NOR2X1_LOC_191/B 0.49fF
C45518 NOR2X1_LOC_694/Y INVX1_LOC_54/A 0.01fF
C45519 INVX1_LOC_222/Y NOR2X1_LOC_799/a_36_216# 0.00fF
C45520 NOR2X1_LOC_791/Y NAND2X1_LOC_357/B 0.02fF
C45521 INVX1_LOC_90/A NOR2X1_LOC_825/a_36_216# 0.00fF
C45522 INVX1_LOC_27/A NOR2X1_LOC_718/B 0.08fF
C45523 NOR2X1_LOC_689/Y NOR2X1_LOC_690/Y 0.00fF
C45524 NOR2X1_LOC_372/A INVX1_LOC_18/A 0.03fF
C45525 NOR2X1_LOC_612/B NOR2X1_LOC_652/Y 0.02fF
C45526 INVX1_LOC_153/Y NOR2X1_LOC_348/Y 0.03fF
C45527 NOR2X1_LOC_100/A INVX1_LOC_50/Y 0.05fF
C45528 INVX1_LOC_245/Y NOR2X1_LOC_596/A 0.03fF
C45529 NOR2X1_LOC_334/A NOR2X1_LOC_461/Y 0.01fF
C45530 INVX1_LOC_278/A NAND2X1_LOC_170/A 0.00fF
C45531 VDD INVX1_LOC_297/A 0.05fF
C45532 INVX1_LOC_13/Y NAND2X1_LOC_360/B 0.07fF
C45533 NOR2X1_LOC_645/a_36_216# INVX1_LOC_141/Y 0.00fF
C45534 NAND2X1_LOC_483/Y NAND2X1_LOC_561/B 0.19fF
C45535 INVX1_LOC_35/A NOR2X1_LOC_146/Y 0.24fF
C45536 NOR2X1_LOC_45/B INVX1_LOC_12/A 0.38fF
C45537 NOR2X1_LOC_332/A INVX1_LOC_57/A 0.08fF
C45538 NOR2X1_LOC_188/Y NOR2X1_LOC_717/A 0.08fF
C45539 INVX1_LOC_95/Y NAND2X1_LOC_63/Y 0.03fF
C45540 NOR2X1_LOC_68/A NOR2X1_LOC_703/B 0.01fF
C45541 NOR2X1_LOC_643/Y INVX1_LOC_31/A 0.05fF
C45542 NAND2X1_LOC_725/A NOR2X1_LOC_690/Y 0.50fF
C45543 INVX1_LOC_135/A INVX1_LOC_53/A 0.05fF
C45544 INVX1_LOC_14/A NOR2X1_LOC_529/Y -0.00fF
C45545 NOR2X1_LOC_82/A NOR2X1_LOC_6/B 0.51fF
C45546 INVX1_LOC_1/A NAND2X1_LOC_301/a_36_24# 0.00fF
C45547 INVX1_LOC_10/A NOR2X1_LOC_53/Y 0.12fF
C45548 INVX1_LOC_243/Y NAND2X1_LOC_651/a_36_24# 0.00fF
C45549 NAND2X1_LOC_773/Y NOR2X1_LOC_226/A 0.18fF
C45550 INVX1_LOC_295/A INVX1_LOC_53/A 1.36fF
C45551 NOR2X1_LOC_486/Y INVX1_LOC_290/Y 0.00fF
C45552 NOR2X1_LOC_136/Y NOR2X1_LOC_321/Y 0.31fF
C45553 INVX1_LOC_233/A NOR2X1_LOC_123/B 0.03fF
C45554 NOR2X1_LOC_67/A INVX1_LOC_269/A 0.10fF
C45555 NOR2X1_LOC_807/B INVX1_LOC_177/A 0.00fF
C45556 INVX1_LOC_131/A INVX1_LOC_270/A 0.07fF
C45557 NOR2X1_LOC_394/a_36_216# INVX1_LOC_23/Y 0.01fF
C45558 NOR2X1_LOC_75/Y NOR2X1_LOC_200/a_36_216# 0.00fF
C45559 INVX1_LOC_18/A NOR2X1_LOC_513/a_36_216# 0.00fF
C45560 NOR2X1_LOC_67/A NOR2X1_LOC_232/Y 0.14fF
C45561 INVX1_LOC_140/A INVX1_LOC_57/A 0.07fF
C45562 INVX1_LOC_256/A INVX1_LOC_177/A 0.03fF
C45563 NOR2X1_LOC_369/Y NOR2X1_LOC_52/B 0.08fF
C45564 NAND2X1_LOC_394/a_36_24# INVX1_LOC_135/A 0.01fF
C45565 INVX1_LOC_307/A NOR2X1_LOC_862/B 0.02fF
C45566 VDD NOR2X1_LOC_89/A 3.36fF
C45567 INVX1_LOC_284/Y INVX1_LOC_240/A 0.01fF
C45568 NOR2X1_LOC_657/Y INVX1_LOC_63/Y 0.02fF
C45569 INVX1_LOC_34/A INVX1_LOC_36/A 0.16fF
C45570 NOR2X1_LOC_750/A NOR2X1_LOC_392/Y 0.02fF
C45571 NAND2X1_LOC_800/A NOR2X1_LOC_89/A 0.03fF
C45572 INVX1_LOC_24/A INVX1_LOC_314/Y 0.03fF
C45573 NOR2X1_LOC_445/B NOR2X1_LOC_862/B 0.10fF
C45574 NOR2X1_LOC_649/a_36_216# NOR2X1_LOC_554/B 0.00fF
C45575 INVX1_LOC_159/A NOR2X1_LOC_433/A 0.00fF
C45576 NOR2X1_LOC_15/Y INVX1_LOC_1/Y 0.16fF
C45577 INPUT_0 INVX1_LOC_270/A 0.05fF
C45578 NOR2X1_LOC_658/Y NOR2X1_LOC_365/a_36_216# 0.01fF
C45579 INVX1_LOC_286/Y NOR2X1_LOC_52/B 0.50fF
C45580 NOR2X1_LOC_441/Y NOR2X1_LOC_361/Y 0.05fF
C45581 NOR2X1_LOC_750/a_36_216# NOR2X1_LOC_392/Y 0.01fF
C45582 NOR2X1_LOC_636/a_36_216# NOR2X1_LOC_68/A 0.00fF
C45583 NAND2X1_LOC_357/B INVX1_LOC_30/A 0.10fF
C45584 NOR2X1_LOC_546/B NOR2X1_LOC_550/B 0.23fF
C45585 INVX1_LOC_12/A INVX1_LOC_281/A 0.13fF
C45586 INVX1_LOC_17/A INVX1_LOC_16/A 0.04fF
C45587 NOR2X1_LOC_435/B NAND2X1_LOC_798/B 0.08fF
C45588 INVX1_LOC_313/Y NOR2X1_LOC_674/Y 0.01fF
C45589 NOR2X1_LOC_111/A NOR2X1_LOC_48/B 0.15fF
C45590 NOR2X1_LOC_45/B NOR2X1_LOC_686/A 0.01fF
C45591 NAND2X1_LOC_729/B NAND2X1_LOC_175/Y 0.05fF
C45592 VDD NOR2X1_LOC_170/A 0.12fF
C45593 INVX1_LOC_84/A INVX1_LOC_179/A 0.03fF
C45594 NAND2X1_LOC_198/B INVX1_LOC_162/A 0.10fF
C45595 NOR2X1_LOC_219/B NOR2X1_LOC_759/Y 0.01fF
C45596 INVX1_LOC_21/A NOR2X1_LOC_473/B 0.01fF
C45597 NAND2X1_LOC_562/a_36_24# NAND2X1_LOC_578/B 0.00fF
C45598 NOR2X1_LOC_82/A INVX1_LOC_30/Y 0.06fF
C45599 NOR2X1_LOC_471/Y INVX1_LOC_16/A 0.03fF
C45600 INVX1_LOC_128/A INVX1_LOC_76/A 0.03fF
C45601 INVX1_LOC_36/A NAND2X1_LOC_231/Y 0.04fF
C45602 INVX1_LOC_34/A NOR2X1_LOC_208/Y 0.08fF
C45603 D_INPUT_1 INVX1_LOC_48/A 0.46fF
C45604 INVX1_LOC_159/A NOR2X1_LOC_52/B 0.04fF
C45605 INVX1_LOC_33/A INVX1_LOC_77/A 0.25fF
C45606 NOR2X1_LOC_550/B INVX1_LOC_275/A 0.09fF
C45607 VDD INVX1_LOC_104/Y 0.21fF
C45608 NAND2X1_LOC_198/B NOR2X1_LOC_315/Y 0.10fF
C45609 INVX1_LOC_64/A NOR2X1_LOC_368/A 0.02fF
C45610 INVX1_LOC_59/A INPUT_1 0.00fF
C45611 INVX1_LOC_174/A GATE_479 0.30fF
C45612 NAND2X1_LOC_338/B INVX1_LOC_72/A 0.01fF
C45613 NOR2X1_LOC_848/Y INVX1_LOC_83/A 1.97fF
C45614 INVX1_LOC_38/A NOR2X1_LOC_861/Y 0.02fF
C45615 NOR2X1_LOC_456/Y INVX1_LOC_78/Y 0.02fF
C45616 INPUT_0 NOR2X1_LOC_109/Y 0.19fF
C45617 INVX1_LOC_249/A NOR2X1_LOC_718/B 0.03fF
C45618 NAND2X1_LOC_655/A NOR2X1_LOC_654/A 0.10fF
C45619 NOR2X1_LOC_794/A INVX1_LOC_53/A 0.06fF
C45620 INVX1_LOC_49/A NOR2X1_LOC_144/Y 0.01fF
C45621 NOR2X1_LOC_168/A NOR2X1_LOC_168/Y 0.06fF
C45622 NAND2X1_LOC_54/a_36_24# INVX1_LOC_61/A 0.01fF
C45623 INVX1_LOC_33/A NOR2X1_LOC_732/A 0.02fF
C45624 NOR2X1_LOC_449/A INVX1_LOC_46/A 0.11fF
C45625 NOR2X1_LOC_739/Y INVX1_LOC_85/Y 0.00fF
C45626 NOR2X1_LOC_778/B INVX1_LOC_24/A 5.90fF
C45627 NOR2X1_LOC_82/a_36_216# INVX1_LOC_22/A 0.00fF
C45628 NOR2X1_LOC_158/Y INVX1_LOC_117/A 0.07fF
C45629 NOR2X1_LOC_536/A INVX1_LOC_4/Y 0.08fF
C45630 INVX1_LOC_314/Y INVX1_LOC_143/A 0.08fF
C45631 INVX1_LOC_34/A NOR2X1_LOC_309/Y 0.03fF
C45632 NOR2X1_LOC_758/Y NOR2X1_LOC_792/B 0.07fF
C45633 NOR2X1_LOC_693/Y NOR2X1_LOC_482/a_36_216# 0.01fF
C45634 NOR2X1_LOC_703/B NOR2X1_LOC_570/Y 0.13fF
C45635 INVX1_LOC_124/A INVX1_LOC_33/A 0.04fF
C45636 NOR2X1_LOC_15/Y NOR2X1_LOC_742/A 0.07fF
C45637 INVX1_LOC_17/A INVX1_LOC_28/A 0.85fF
C45638 NAND2X1_LOC_291/B NOR2X1_LOC_240/A 0.03fF
C45639 NOR2X1_LOC_441/Y NOR2X1_LOC_355/A 0.02fF
C45640 NAND2X1_LOC_733/A NOR2X1_LOC_299/Y 0.13fF
C45641 NOR2X1_LOC_321/Y INVX1_LOC_144/A 0.07fF
C45642 NAND2X1_LOC_81/B INVX1_LOC_3/A 0.02fF
C45643 INVX1_LOC_310/A INVX1_LOC_310/Y 0.19fF
C45644 NOR2X1_LOC_272/Y INVX1_LOC_286/A 0.10fF
C45645 INVX1_LOC_49/Y INVX1_LOC_63/A 0.03fF
C45646 INVX1_LOC_20/A NOR2X1_LOC_696/Y 0.11fF
C45647 INVX1_LOC_77/A INVX1_LOC_40/A 0.03fF
C45648 NOR2X1_LOC_52/Y INVX1_LOC_10/A 0.01fF
C45649 NAND2X1_LOC_223/A INVX1_LOC_9/A 0.16fF
C45650 INVX1_LOC_2/A NOR2X1_LOC_144/Y 0.06fF
C45651 INVX1_LOC_313/Y NOR2X1_LOC_348/a_36_216# 0.01fF
C45652 INVX1_LOC_21/A NOR2X1_LOC_355/B 0.07fF
C45653 NOR2X1_LOC_270/Y INVX1_LOC_10/A 0.02fF
C45654 NOR2X1_LOC_354/B NOR2X1_LOC_326/Y 0.10fF
C45655 NOR2X1_LOC_78/B NOR2X1_LOC_388/Y 0.03fF
C45656 INVX1_LOC_266/Y NOR2X1_LOC_75/a_36_216# 0.01fF
C45657 INVX1_LOC_224/A NOR2X1_LOC_721/Y 0.02fF
C45658 INVX1_LOC_225/A NAND2X1_LOC_342/Y 0.11fF
C45659 NAND2X1_LOC_357/B NAND2X1_LOC_722/A 0.02fF
C45660 INVX1_LOC_99/A INVX1_LOC_63/A 0.05fF
C45661 INVX1_LOC_88/A NOR2X1_LOC_815/A 0.00fF
C45662 NAND2X1_LOC_231/Y NOR2X1_LOC_309/Y 0.10fF
C45663 NOR2X1_LOC_38/B INVX1_LOC_46/Y 0.07fF
C45664 NAND2X1_LOC_863/a_36_24# NAND2X1_LOC_863/Y 0.02fF
C45665 NAND2X1_LOC_93/B INVX1_LOC_4/Y 0.42fF
C45666 INVX1_LOC_271/A NAND2X1_LOC_472/Y 0.14fF
C45667 INVX1_LOC_45/A NAND2X1_LOC_842/B 0.07fF
C45668 INVX1_LOC_54/Y NOR2X1_LOC_709/A 0.12fF
C45669 D_INPUT_0 INVX1_LOC_62/Y 0.19fF
C45670 INVX1_LOC_72/A INVX1_LOC_313/Y 0.03fF
C45671 NOR2X1_LOC_662/A INVX1_LOC_42/A 0.10fF
C45672 INVX1_LOC_33/A NOR2X1_LOC_687/Y 0.19fF
C45673 NAND2X1_LOC_656/Y NOR2X1_LOC_759/Y 0.01fF
C45674 NAND2X1_LOC_354/B NAND2X1_LOC_834/a_36_24# 0.00fF
C45675 NAND2X1_LOC_326/a_36_24# NAND2X1_LOC_840/B 0.00fF
C45676 NOR2X1_LOC_465/Y INVX1_LOC_307/A 0.10fF
C45677 NAND2X1_LOC_564/B NAND2X1_LOC_833/Y 0.03fF
C45678 INVX1_LOC_41/A NAND2X1_LOC_390/a_36_24# 0.00fF
C45679 NOR2X1_LOC_91/Y NAND2X1_LOC_862/Y 0.01fF
C45680 NOR2X1_LOC_828/B NOR2X1_LOC_726/Y 0.02fF
C45681 INVX1_LOC_202/A NAND2X1_LOC_656/Y 0.42fF
C45682 NOR2X1_LOC_590/A NAND2X1_LOC_840/Y 0.01fF
C45683 INVX1_LOC_39/A INVX1_LOC_95/Y 0.00fF
C45684 INVX1_LOC_162/A INVX1_LOC_53/Y 0.10fF
C45685 INVX1_LOC_43/Y NOR2X1_LOC_368/A 0.28fF
C45686 INVX1_LOC_279/A INVX1_LOC_49/A 0.07fF
C45687 INVX1_LOC_256/A INVX1_LOC_285/Y 0.10fF
C45688 NOR2X1_LOC_15/Y NOR2X1_LOC_318/B 0.07fF
C45689 NAND2X1_LOC_555/Y NAND2X1_LOC_126/a_36_24# -0.01fF
C45690 INVX1_LOC_12/A NOR2X1_LOC_1/Y 0.01fF
C45691 NOR2X1_LOC_772/a_36_216# NOR2X1_LOC_309/Y 0.00fF
C45692 NAND2X1_LOC_338/B NOR2X1_LOC_537/Y 0.07fF
C45693 INVX1_LOC_36/A INVX1_LOC_131/A 0.07fF
C45694 NOR2X1_LOC_172/Y NOR2X1_LOC_561/Y 0.02fF
C45695 NOR2X1_LOC_290/Y NAND2X1_LOC_334/a_36_24# 0.00fF
C45696 INVX1_LOC_176/A INVX1_LOC_50/Y 0.03fF
C45697 NOR2X1_LOC_392/B NOR2X1_LOC_719/A 0.04fF
C45698 INVX1_LOC_30/A NAND2X1_LOC_849/A 0.07fF
C45699 NOR2X1_LOC_446/A INVX1_LOC_206/Y 0.01fF
C45700 INVX1_LOC_11/A NOR2X1_LOC_337/Y 0.01fF
C45701 NOR2X1_LOC_791/B NOR2X1_LOC_756/Y 0.03fF
C45702 NOR2X1_LOC_315/Y INVX1_LOC_53/Y 0.03fF
C45703 NOR2X1_LOC_15/Y INVX1_LOC_93/Y 0.26fF
C45704 NOR2X1_LOC_649/B INVX1_LOC_4/Y 0.03fF
C45705 NAND2X1_LOC_572/a_36_24# NOR2X1_LOC_82/Y 0.00fF
C45706 INVX1_LOC_3/A INVX1_LOC_4/Y 0.01fF
C45707 NAND2X1_LOC_338/B NAND2X1_LOC_323/B 0.02fF
C45708 NOR2X1_LOC_577/Y NAND2X1_LOC_140/A 0.01fF
C45709 INVX1_LOC_18/A NAND2X1_LOC_560/A 0.00fF
C45710 INVX1_LOC_200/A NOR2X1_LOC_45/B 0.15fF
C45711 NOR2X1_LOC_78/B NOR2X1_LOC_366/B 0.03fF
C45712 NAND2X1_LOC_308/Y NOR2X1_LOC_690/Y 0.00fF
C45713 NOR2X1_LOC_67/A NAND2X1_LOC_563/A 0.02fF
C45714 INVX1_LOC_233/Y NOR2X1_LOC_536/A 0.01fF
C45715 INVX1_LOC_222/Y INVX1_LOC_37/A 0.03fF
C45716 NOR2X1_LOC_88/Y NOR2X1_LOC_693/Y 0.07fF
C45717 NOR2X1_LOC_583/Y NOR2X1_LOC_48/B 0.12fF
C45718 INVX1_LOC_36/A INPUT_0 7.45fF
C45719 NOR2X1_LOC_355/A NOR2X1_LOC_142/Y 0.10fF
C45720 INVX1_LOC_271/A NAND2X1_LOC_434/Y 0.01fF
C45721 NAND2X1_LOC_778/Y NAND2X1_LOC_721/A 0.00fF
C45722 INVX1_LOC_24/A NOR2X1_LOC_597/Y 0.03fF
C45723 NOR2X1_LOC_667/A NAND2X1_LOC_711/a_36_24# 0.01fF
C45724 INVX1_LOC_78/A NOR2X1_LOC_662/A 0.01fF
C45725 NOR2X1_LOC_78/B NAND2X1_LOC_479/Y 0.03fF
C45726 INVX1_LOC_11/A NOR2X1_LOC_56/Y 0.07fF
C45727 NOR2X1_LOC_500/Y NOR2X1_LOC_388/a_36_216# 0.01fF
C45728 INVX1_LOC_240/A NOR2X1_LOC_525/Y 0.04fF
C45729 NOR2X1_LOC_590/A NOR2X1_LOC_78/A 0.13fF
C45730 NAND2X1_LOC_733/a_36_24# NAND2X1_LOC_560/A 0.01fF
C45731 INVX1_LOC_2/A INVX1_LOC_279/A 0.07fF
C45732 NAND2X1_LOC_733/Y NOR2X1_LOC_45/B 0.03fF
C45733 NOR2X1_LOC_637/A INVX1_LOC_144/A 0.03fF
C45734 INVX1_LOC_84/A NOR2X1_LOC_693/Y 0.07fF
C45735 INVX1_LOC_17/A NOR2X1_LOC_35/Y 0.98fF
C45736 INVX1_LOC_22/A NOR2X1_LOC_315/a_36_216# 0.00fF
C45737 INVX1_LOC_22/Y NOR2X1_LOC_78/A 0.02fF
C45738 INVX1_LOC_172/A NAND2X1_LOC_560/A 0.05fF
C45739 INVX1_LOC_151/Y INVX1_LOC_22/A 0.01fF
C45740 NOR2X1_LOC_91/A NOR2X1_LOC_653/Y 0.01fF
C45741 INVX1_LOC_89/A INVX1_LOC_85/A 0.03fF
C45742 INVX1_LOC_298/Y INVX1_LOC_186/Y 0.15fF
C45743 NAND2X1_LOC_53/Y NOR2X1_LOC_603/Y 0.02fF
C45744 INVX1_LOC_225/A NOR2X1_LOC_246/Y 0.24fF
C45745 NAND2X1_LOC_288/A INVX1_LOC_23/A 0.08fF
C45746 NAND2X1_LOC_222/B VDD 0.04fF
C45747 NAND2X1_LOC_596/a_36_24# INVX1_LOC_10/A 0.01fF
C45748 NOR2X1_LOC_449/a_36_216# INVX1_LOC_144/A 0.01fF
C45749 NAND2X1_LOC_364/A INVX1_LOC_286/A 0.08fF
C45750 NOR2X1_LOC_15/Y NAND2X1_LOC_721/A 0.31fF
C45751 NOR2X1_LOC_632/Y INVX1_LOC_208/A 0.00fF
C45752 NOR2X1_LOC_92/Y INVX1_LOC_33/Y 0.03fF
C45753 NOR2X1_LOC_736/Y NOR2X1_LOC_142/Y 0.08fF
C45754 NAND2X1_LOC_579/A INVX1_LOC_37/Y 0.43fF
C45755 INVX1_LOC_5/A INVX1_LOC_274/A 0.07fF
C45756 NAND2X1_LOC_341/A NOR2X1_LOC_589/A 0.03fF
C45757 INVX1_LOC_21/A INVX1_LOC_193/A 0.05fF
C45758 NAND2X1_LOC_396/a_36_24# NOR2X1_LOC_266/B 0.00fF
C45759 NOR2X1_LOC_315/Y NOR2X1_LOC_76/a_36_216# 0.01fF
C45760 INVX1_LOC_11/A VDD 1.74fF
C45761 INVX1_LOC_90/A NAND2X1_LOC_629/Y 0.01fF
C45762 INVX1_LOC_135/A NOR2X1_LOC_78/B 0.50fF
C45763 NOR2X1_LOC_237/Y INPUT_0 0.00fF
C45764 NOR2X1_LOC_91/A INVX1_LOC_19/A 0.06fF
C45765 INVX1_LOC_230/Y INVX1_LOC_20/A 0.11fF
C45766 NOR2X1_LOC_392/Y INVX1_LOC_123/Y 0.15fF
C45767 NOR2X1_LOC_668/Y INVX1_LOC_19/A 0.08fF
C45768 NAND2X1_LOC_381/Y VDD 0.06fF
C45769 INVX1_LOC_36/A NAND2X1_LOC_649/B 0.00fF
C45770 INVX1_LOC_217/A NOR2X1_LOC_45/B 0.05fF
C45771 NAND2X1_LOC_555/Y NOR2X1_LOC_35/Y 0.12fF
C45772 NAND2X1_LOC_355/Y NOR2X1_LOC_45/B 0.01fF
C45773 NOR2X1_LOC_589/A GATE_479 0.01fF
C45774 NOR2X1_LOC_68/A INVX1_LOC_91/A 1.29fF
C45775 NOR2X1_LOC_428/a_36_216# INVX1_LOC_37/A 0.00fF
C45776 INVX1_LOC_49/Y NOR2X1_LOC_65/Y 0.01fF
C45777 NOR2X1_LOC_804/B INPUT_0 0.07fF
C45778 INVX1_LOC_63/Y NOR2X1_LOC_74/A 0.10fF
C45779 INVX1_LOC_119/Y NAND2X1_LOC_793/B 0.07fF
C45780 NOR2X1_LOC_843/B INVX1_LOC_29/A 0.03fF
C45781 INVX1_LOC_24/A NOR2X1_LOC_557/A 0.01fF
C45782 NAND2X1_LOC_364/A INVX1_LOC_95/A 0.09fF
C45783 NOR2X1_LOC_828/A NOR2X1_LOC_544/A 0.32fF
C45784 INVX1_LOC_5/A NOR2X1_LOC_820/Y 0.39fF
C45785 NOR2X1_LOC_55/a_36_216# INVX1_LOC_42/A 0.03fF
C45786 NOR2X1_LOC_550/B INVX1_LOC_78/Y 0.03fF
C45787 INVX1_LOC_23/A INVX1_LOC_19/A 1.49fF
C45788 NAND2X1_LOC_715/B NOR2X1_LOC_127/a_36_216# 0.00fF
C45789 INVX1_LOC_2/A INVX1_LOC_182/Y 0.03fF
C45790 INVX1_LOC_100/A INVX1_LOC_8/A 1.98fF
C45791 NOR2X1_LOC_309/Y INPUT_0 0.20fF
C45792 INVX1_LOC_269/A NOR2X1_LOC_729/A 0.07fF
C45793 INVX1_LOC_1/A NOR2X1_LOC_612/Y 0.02fF
C45794 NAND2X1_LOC_661/A NAND2X1_LOC_661/B 0.07fF
C45795 NOR2X1_LOC_441/Y NOR2X1_LOC_111/A 0.00fF
C45796 NAND2X1_LOC_564/B NOR2X1_LOC_76/A 0.01fF
C45797 INVX1_LOC_13/Y NAND2X1_LOC_572/B 0.07fF
C45798 NOR2X1_LOC_477/a_36_216# INVX1_LOC_117/A 0.01fF
C45799 INVX1_LOC_89/A NAND2X1_LOC_662/Y 0.07fF
C45800 NOR2X1_LOC_590/A NOR2X1_LOC_98/a_36_216# 0.00fF
C45801 INVX1_LOC_135/A NOR2X1_LOC_459/A 0.22fF
C45802 NOR2X1_LOC_186/Y INVX1_LOC_285/A 0.08fF
C45803 INVX1_LOC_57/A NOR2X1_LOC_847/A 0.28fF
C45804 NOR2X1_LOC_667/A NOR2X1_LOC_322/Y 0.02fF
C45805 NAND2X1_LOC_214/B NAND2X1_LOC_206/Y 0.07fF
C45806 NOR2X1_LOC_209/a_36_216# INVX1_LOC_85/Y 0.00fF
C45807 NOR2X1_LOC_660/Y NAND2X1_LOC_82/Y 0.12fF
C45808 INVX1_LOC_57/A INVX1_LOC_42/A 0.20fF
C45809 INVX1_LOC_135/A INVX1_LOC_83/A 0.07fF
C45810 INVX1_LOC_2/A NAND2X1_LOC_858/B 0.09fF
C45811 NOR2X1_LOC_205/Y NAND2X1_LOC_93/B 0.03fF
C45812 NOR2X1_LOC_186/Y NOR2X1_LOC_814/A 0.00fF
C45813 INVX1_LOC_90/A NOR2X1_LOC_561/Y 0.19fF
C45814 INVX1_LOC_266/Y INVX1_LOC_6/A 0.03fF
C45815 NOR2X1_LOC_175/A NOR2X1_LOC_9/Y 0.00fF
C45816 NOR2X1_LOC_433/A NOR2X1_LOC_56/Y 0.07fF
C45817 NAND2X1_LOC_340/a_36_24# INVX1_LOC_118/A 0.00fF
C45818 NOR2X1_LOC_788/a_36_216# INVX1_LOC_177/A 0.00fF
C45819 NOR2X1_LOC_389/B NOR2X1_LOC_561/Y 0.07fF
C45820 INVX1_LOC_295/A INVX1_LOC_83/A 0.79fF
C45821 INVX1_LOC_27/A NAND2X1_LOC_206/Y 0.07fF
C45822 INVX1_LOC_104/A INVX1_LOC_186/A 0.07fF
C45823 NOR2X1_LOC_474/A NAND2X1_LOC_659/B 0.05fF
C45824 NOR2X1_LOC_559/B INVX1_LOC_176/A -0.00fF
C45825 NOR2X1_LOC_565/a_36_216# NOR2X1_LOC_500/Y 0.02fF
C45826 NAND2X1_LOC_391/Y NAND2X1_LOC_768/Y 0.01fF
C45827 NOR2X1_LOC_53/Y INVX1_LOC_12/A 0.23fF
C45828 NOR2X1_LOC_68/A NOR2X1_LOC_698/Y 0.03fF
C45829 NAND2X1_LOC_541/a_36_24# INVX1_LOC_42/A 0.00fF
C45830 NAND2X1_LOC_348/A NOR2X1_LOC_719/A 0.00fF
C45831 INVX1_LOC_209/Y NOR2X1_LOC_314/a_36_216# 0.00fF
C45832 INVX1_LOC_27/A NAND2X1_LOC_773/B 0.07fF
C45833 NOR2X1_LOC_503/Y NOR2X1_LOC_510/B 1.53fF
C45834 NOR2X1_LOC_172/Y INVX1_LOC_76/A 0.01fF
C45835 NOR2X1_LOC_433/A VDD 2.09fF
C45836 INVX1_LOC_50/Y NOR2X1_LOC_340/A 0.13fF
C45837 NOR2X1_LOC_474/A VDD 0.24fF
C45838 INVX1_LOC_143/A NOR2X1_LOC_557/A 0.02fF
C45839 NOR2X1_LOC_68/A NAND2X1_LOC_783/a_36_24# 0.01fF
C45840 NAND2X1_LOC_348/A INVX1_LOC_7/A 0.04fF
C45841 INVX1_LOC_249/A NAND2X1_LOC_472/Y 0.01fF
C45842 INVX1_LOC_104/A NAND2X1_LOC_447/Y 0.10fF
C45843 NOR2X1_LOC_52/B NOR2X1_LOC_56/Y 0.07fF
C45844 NOR2X1_LOC_147/B INVX1_LOC_76/A 0.03fF
C45845 NOR2X1_LOC_593/Y VDD 0.40fF
C45846 NOR2X1_LOC_597/Y NAND2X1_LOC_800/Y 0.00fF
C45847 NOR2X1_LOC_510/Y NOR2X1_LOC_89/A 1.53fF
C45848 INVX1_LOC_21/A INVX1_LOC_106/A 0.01fF
C45849 INVX1_LOC_214/Y NOR2X1_LOC_45/B 0.03fF
C45850 NOR2X1_LOC_208/a_36_216# INVX1_LOC_78/Y 0.00fF
C45851 INVX1_LOC_6/Y NAND2X1_LOC_472/Y 0.04fF
C45852 INVX1_LOC_78/A INVX1_LOC_57/A 0.20fF
C45853 NOR2X1_LOC_388/Y INVX1_LOC_46/A 0.07fF
C45854 NOR2X1_LOC_392/B INVX1_LOC_76/A 0.03fF
C45855 NOR2X1_LOC_315/Y NAND2X1_LOC_465/A 0.01fF
C45856 NAND2X1_LOC_364/A INVX1_LOC_54/A 0.03fF
C45857 NOR2X1_LOC_78/B NOR2X1_LOC_552/A 0.01fF
C45858 NAND2X1_LOC_671/a_36_24# INVX1_LOC_315/Y 0.00fF
C45859 INVX1_LOC_151/A VDD -0.00fF
C45860 NOR2X1_LOC_82/Y INVX1_LOC_98/A 0.13fF
C45861 NAND2X1_LOC_773/Y NAND2X1_LOC_63/Y 0.05fF
C45862 NOR2X1_LOC_52/B INVX1_LOC_146/Y 0.01fF
C45863 NOR2X1_LOC_82/Y NOR2X1_LOC_78/A 0.03fF
C45864 NOR2X1_LOC_52/B VDD 1.21fF
C45865 NOR2X1_LOC_113/B INVX1_LOC_66/A 0.01fF
C45866 NAND2X1_LOC_842/B INVX1_LOC_102/Y 0.10fF
C45867 INVX1_LOC_26/A INVX1_LOC_129/A -0.00fF
C45868 NOR2X1_LOC_97/A INVX1_LOC_120/A 0.00fF
C45869 INVX1_LOC_75/A D_GATE_366 0.07fF
C45870 NAND2X1_LOC_838/Y VDD 0.16fF
C45871 INVX1_LOC_83/A NOR2X1_LOC_711/A 0.10fF
C45872 D_INPUT_0 INVX1_LOC_51/Y 0.00fF
C45873 INVX1_LOC_96/Y INVX1_LOC_139/A 0.00fF
C45874 INVX1_LOC_49/A NOR2X1_LOC_450/A 0.03fF
C45875 INVX1_LOC_26/Y INVX1_LOC_23/A 0.03fF
C45876 NOR2X1_LOC_65/B INVX1_LOC_57/A 0.07fF
C45877 NOR2X1_LOC_577/Y INVX1_LOC_118/Y 0.03fF
C45878 NOR2X1_LOC_423/Y INVX1_LOC_37/A 0.06fF
C45879 NOR2X1_LOC_383/B NAND2X1_LOC_90/a_36_24# 0.02fF
C45880 NOR2X1_LOC_844/A NOR2X1_LOC_859/Y 0.02fF
C45881 INVX1_LOC_18/A NOR2X1_LOC_58/Y 0.10fF
C45882 NOR2X1_LOC_689/Y NAND2X1_LOC_724/Y 0.12fF
C45883 NOR2X1_LOC_361/B NOR2X1_LOC_89/A 1.07fF
C45884 INVX1_LOC_99/Y NOR2X1_LOC_334/Y 0.01fF
C45885 INVX1_LOC_62/Y INVX1_LOC_46/Y 0.11fF
C45886 NOR2X1_LOC_588/A INPUT_5 0.07fF
C45887 NAND2X1_LOC_858/B INPUT_1 0.00fF
C45888 INVX1_LOC_215/A NOR2X1_LOC_405/A 0.14fF
C45889 INVX1_LOC_33/A INVX1_LOC_9/A 0.20fF
C45890 INVX1_LOC_60/A NOR2X1_LOC_98/B 0.03fF
C45891 INVX1_LOC_90/A NOR2X1_LOC_167/Y 0.03fF
C45892 NAND2X1_LOC_477/A INVX1_LOC_33/Y 0.03fF
C45893 D_INPUT_1 NOR2X1_LOC_383/B 0.20fF
C45894 INVX1_LOC_227/A NOR2X1_LOC_78/A 0.02fF
C45895 NOR2X1_LOC_787/a_36_216# INVX1_LOC_29/A 0.00fF
C45896 INVX1_LOC_93/A NAND2X1_LOC_444/B 0.03fF
C45897 NAND2X1_LOC_395/a_36_24# NOR2X1_LOC_266/B 0.00fF
C45898 INVX1_LOC_278/A NOR2X1_LOC_693/Y 0.09fF
C45899 INVX1_LOC_13/Y NOR2X1_LOC_394/Y 0.01fF
C45900 NOR2X1_LOC_594/Y INVX1_LOC_28/A 0.02fF
C45901 NOR2X1_LOC_78/B INVX1_LOC_139/Y 0.04fF
C45902 NOR2X1_LOC_380/Y NAND2X1_LOC_463/B 0.19fF
C45903 NOR2X1_LOC_45/B NAND2X1_LOC_808/A 0.08fF
C45904 INVX1_LOC_31/A INVX1_LOC_19/A 0.33fF
C45905 NAND2X1_LOC_114/B NAND2X1_LOC_74/B 0.26fF
C45906 NOR2X1_LOC_222/Y INVX1_LOC_37/A 0.03fF
C45907 NOR2X1_LOC_67/A INVX1_LOC_12/Y 0.08fF
C45908 INVX1_LOC_314/Y NOR2X1_LOC_197/B 0.01fF
C45909 NOR2X1_LOC_443/Y NAND2X1_LOC_363/B 0.01fF
C45910 NAND2X1_LOC_228/a_36_24# INVX1_LOC_76/A 0.01fF
C45911 INVX1_LOC_144/Y NOR2X1_LOC_506/a_36_216# 0.00fF
C45912 INVX1_LOC_187/Y INPUT_5 0.29fF
C45913 NOR2X1_LOC_78/B INVX1_LOC_10/Y 0.03fF
C45914 NOR2X1_LOC_512/a_36_216# INVX1_LOC_76/A 0.00fF
C45915 NOR2X1_LOC_742/A NOR2X1_LOC_733/Y 0.27fF
C45916 NOR2X1_LOC_147/A NOR2X1_LOC_706/A 0.06fF
C45917 NOR2X1_LOC_526/Y NOR2X1_LOC_536/A 0.01fF
C45918 INVX1_LOC_312/Y NAND2X1_LOC_74/B 0.14fF
C45919 NOR2X1_LOC_78/B INVX1_LOC_280/A 1.57fF
C45920 D_INPUT_0 NAND2X1_LOC_655/B 0.03fF
C45921 NAND2X1_LOC_785/A INVX1_LOC_54/A 0.76fF
C45922 NOR2X1_LOC_294/Y NAND2X1_LOC_207/Y 0.72fF
C45923 NOR2X1_LOC_383/B NOR2X1_LOC_652/Y 0.08fF
C45924 INVX1_LOC_289/Y INVX1_LOC_273/A 0.03fF
C45925 INVX1_LOC_45/A INVX1_LOC_284/A 0.72fF
C45926 NOR2X1_LOC_15/Y INVX1_LOC_87/A 0.16fF
C45927 INVX1_LOC_26/A NOR2X1_LOC_440/B 0.28fF
C45928 NOR2X1_LOC_619/A NAND2X1_LOC_96/A 0.03fF
C45929 NOR2X1_LOC_78/A NOR2X1_LOC_703/A 0.03fF
C45930 INVX1_LOC_50/A NOR2X1_LOC_406/A 0.00fF
C45931 INVX1_LOC_41/A NAND2X1_LOC_52/a_36_24# 0.00fF
C45932 INVX1_LOC_18/A INVX1_LOC_29/A 0.25fF
C45933 NOR2X1_LOC_724/Y NOR2X1_LOC_209/A 0.06fF
C45934 INVX1_LOC_111/A INVX1_LOC_19/A 0.00fF
C45935 NOR2X1_LOC_92/Y INVX1_LOC_23/Y 0.03fF
C45936 INVX1_LOC_40/A INVX1_LOC_9/A 1.76fF
C45937 NOR2X1_LOC_270/Y INVX1_LOC_12/A 0.07fF
C45938 INVX1_LOC_256/A INVX1_LOC_4/Y 0.17fF
C45939 INVX1_LOC_69/Y INVX1_LOC_285/Y 0.10fF
C45940 INVX1_LOC_135/A INVX1_LOC_46/A 0.03fF
C45941 INVX1_LOC_147/A INVX1_LOC_91/A 0.01fF
C45942 INVX1_LOC_230/Y INVX1_LOC_4/A 0.06fF
C45943 NAND2X1_LOC_20/B NAND2X1_LOC_223/A 0.29fF
C45944 NOR2X1_LOC_598/B INVX1_LOC_298/A 0.01fF
C45945 NAND2X1_LOC_364/A NAND2X1_LOC_807/B 0.09fF
C45946 NAND2X1_LOC_231/Y NOR2X1_LOC_435/A 0.03fF
C45947 NAND2X1_LOC_149/Y INVX1_LOC_296/A 0.18fF
C45948 INVX1_LOC_90/A INVX1_LOC_76/A 0.26fF
C45949 NAND2X1_LOC_860/A NOR2X1_LOC_81/Y 0.03fF
C45950 INVX1_LOC_22/A INVX1_LOC_118/Y 0.03fF
C45951 NAND2X1_LOC_218/a_36_24# NAND2X1_LOC_218/A 0.00fF
C45952 INVX1_LOC_225/A INVX1_LOC_285/A 0.10fF
C45953 NOR2X1_LOC_561/Y NOR2X1_LOC_561/A 0.06fF
C45954 NOR2X1_LOC_641/B INVX1_LOC_15/A 0.06fF
C45955 INVX1_LOC_34/A INVX1_LOC_63/A 0.07fF
C45956 NOR2X1_LOC_433/A INVX1_LOC_133/A 0.69fF
C45957 INVX1_LOC_82/A INVX1_LOC_3/A 0.05fF
C45958 NOR2X1_LOC_561/Y INVX1_LOC_38/A 0.15fF
C45959 NOR2X1_LOC_458/B INVX1_LOC_307/A 0.01fF
C45960 NAND2X1_LOC_535/a_36_24# INVX1_LOC_94/Y 0.00fF
C45961 INVX1_LOC_225/A NOR2X1_LOC_814/A 0.07fF
C45962 INVX1_LOC_311/A NOR2X1_LOC_562/B 0.02fF
C45963 NOR2X1_LOC_778/B NOR2X1_LOC_197/B 0.04fF
C45964 NOR2X1_LOC_751/Y INVX1_LOC_15/A 0.06fF
C45965 NOR2X1_LOC_606/Y INVX1_LOC_4/Y 0.22fF
C45966 NOR2X1_LOC_174/B INVX1_LOC_117/A 0.10fF
C45967 NAND2X1_LOC_740/B INVX1_LOC_20/A 0.01fF
C45968 INVX1_LOC_83/A INVX1_LOC_280/A 0.07fF
C45969 NOR2X1_LOC_91/A INVX1_LOC_161/Y 0.04fF
C45970 NOR2X1_LOC_187/Y INVX1_LOC_29/Y 0.14fF
C45971 NOR2X1_LOC_135/Y NAND2X1_LOC_211/Y 0.07fF
C45972 NOR2X1_LOC_329/B NOR2X1_LOC_681/Y 0.05fF
C45973 NOR2X1_LOC_564/a_36_216# NOR2X1_LOC_78/A 0.01fF
C45974 NOR2X1_LOC_329/B INVX1_LOC_37/A 0.10fF
C45975 INVX1_LOC_55/Y INVX1_LOC_117/A 0.09fF
C45976 NAND2X1_LOC_326/a_36_24# INVX1_LOC_49/Y 0.00fF
C45977 INVX1_LOC_54/Y INVX1_LOC_294/A 0.00fF
C45978 INVX1_LOC_286/A NOR2X1_LOC_405/A 0.03fF
C45979 INVX1_LOC_122/Y NOR2X1_LOC_227/A 0.01fF
C45980 D_INPUT_4 INVX1_LOC_37/A 0.01fF
C45981 NAND2X1_LOC_231/Y INVX1_LOC_63/A 0.10fF
C45982 NOR2X1_LOC_52/B INVX1_LOC_133/A 0.07fF
C45983 INVX1_LOC_31/A INVX1_LOC_26/Y 0.18fF
C45984 INVX1_LOC_161/Y INVX1_LOC_23/A 0.07fF
C45985 INVX1_LOC_206/Y NAND2X1_LOC_447/Y 0.03fF
C45986 NAND2X1_LOC_830/a_36_24# NOR2X1_LOC_536/A 0.00fF
C45987 INVX1_LOC_64/A NOR2X1_LOC_359/a_36_216# 0.01fF
C45988 NOR2X1_LOC_599/Y INVX1_LOC_296/Y 0.46fF
C45989 INVX1_LOC_89/A NAND2X1_LOC_62/a_36_24# 0.00fF
C45990 INVX1_LOC_140/Y VDD 0.21fF
C45991 INVX1_LOC_298/Y INVX1_LOC_18/A 0.03fF
C45992 NOR2X1_LOC_500/A NOR2X1_LOC_334/Y 0.07fF
C45993 INVX1_LOC_59/A INVX1_LOC_39/A 0.02fF
C45994 INVX1_LOC_255/Y INVX1_LOC_84/A 0.11fF
C45995 NOR2X1_LOC_303/Y NOR2X1_LOC_334/Y 0.10fF
C45996 INVX1_LOC_177/A NOR2X1_LOC_89/A 0.03fF
C45997 NOR2X1_LOC_71/Y NOR2X1_LOC_88/Y 0.03fF
C45998 NOR2X1_LOC_332/A NOR2X1_LOC_820/Y 0.03fF
C45999 NAND2X1_LOC_473/A NAND2X1_LOC_218/A 0.00fF
C46000 NOR2X1_LOC_576/B NAND2X1_LOC_770/Y 0.26fF
C46001 NAND2X1_LOC_198/B NAND2X1_LOC_99/A 0.08fF
C46002 INVX1_LOC_224/Y INVX1_LOC_72/A 0.00fF
C46003 INVX1_LOC_230/Y INVX1_LOC_64/A 0.08fF
C46004 NOR2X1_LOC_778/A NOR2X1_LOC_383/B 0.01fF
C46005 INVX1_LOC_137/A NAND2X1_LOC_773/B 0.01fF
C46006 NOR2X1_LOC_124/A INVX1_LOC_59/Y 0.00fF
C46007 INVX1_LOC_311/A INVX1_LOC_281/Y 0.04fF
C46008 NOR2X1_LOC_554/B INVX1_LOC_57/A 0.73fF
C46009 NOR2X1_LOC_329/B NOR2X1_LOC_743/Y 0.04fF
C46010 NOR2X1_LOC_786/a_36_216# INVX1_LOC_306/Y 0.00fF
C46011 NOR2X1_LOC_510/Y INVX1_LOC_11/A 0.07fF
C46012 NAND2X1_LOC_803/B NOR2X1_LOC_186/Y 0.00fF
C46013 NOR2X1_LOC_552/A INVX1_LOC_46/A 0.12fF
C46014 NOR2X1_LOC_717/Y NOR2X1_LOC_678/A 0.22fF
C46015 D_GATE_741 NOR2X1_LOC_460/Y 0.00fF
C46016 NOR2X1_LOC_254/Y NOR2X1_LOC_334/Y 0.01fF
C46017 NAND2X1_LOC_11/Y NOR2X1_LOC_48/B 0.00fF
C46018 NAND2X1_LOC_387/B INVX1_LOC_53/A 0.01fF
C46019 NOR2X1_LOC_71/Y INVX1_LOC_84/A 0.03fF
C46020 INVX1_LOC_289/Y NOR2X1_LOC_15/Y 0.36fF
C46021 NOR2X1_LOC_658/Y NOR2X1_LOC_423/a_36_216# 0.01fF
C46022 INVX1_LOC_58/A NOR2X1_LOC_759/A 0.24fF
C46023 NOR2X1_LOC_789/A NAND2X1_LOC_74/B 0.24fF
C46024 NOR2X1_LOC_210/B INVX1_LOC_114/Y 0.02fF
C46025 INVX1_LOC_182/A NOR2X1_LOC_600/a_36_216# 0.01fF
C46026 INVX1_LOC_292/A INVX1_LOC_50/Y 0.07fF
C46027 NOR2X1_LOC_205/Y NOR2X1_LOC_348/Y 0.01fF
C46028 INVX1_LOC_25/Y INVX1_LOC_102/A 0.07fF
C46029 NOR2X1_LOC_598/B INVX1_LOC_205/A 0.00fF
C46030 VDD NOR2X1_LOC_601/Y 0.24fF
C46031 INVX1_LOC_199/A VDD 0.14fF
C46032 INVX1_LOC_24/A INVX1_LOC_271/A 0.06fF
C46033 INVX1_LOC_77/A NOR2X1_LOC_635/B 0.03fF
C46034 NOR2X1_LOC_188/A NOR2X1_LOC_612/Y 0.02fF
C46035 NOR2X1_LOC_186/Y NOR2X1_LOC_590/A 0.06fF
C46036 NOR2X1_LOC_607/Y NOR2X1_LOC_383/B 0.05fF
C46037 NAND2X1_LOC_861/Y NOR2X1_LOC_662/A 0.07fF
C46038 INVX1_LOC_2/A NOR2X1_LOC_38/B 0.00fF
C46039 NAND2X1_LOC_803/B NAND2X1_LOC_573/Y 0.01fF
C46040 INVX1_LOC_41/A INVX1_LOC_23/Y 0.02fF
C46041 INVX1_LOC_77/A INVX1_LOC_275/Y 0.03fF
C46042 INVX1_LOC_50/A NOR2X1_LOC_495/Y 0.02fF
C46043 NOR2X1_LOC_550/B NOR2X1_LOC_727/B 0.01fF
C46044 VDD INVX1_LOC_74/A 0.29fF
C46045 NAND2X1_LOC_537/Y NAND2X1_LOC_538/Y 0.04fF
C46046 NAND2X1_LOC_181/Y INVX1_LOC_32/A 0.03fF
C46047 NOR2X1_LOC_152/Y INVX1_LOC_57/A 0.07fF
C46048 INVX1_LOC_77/A NOR2X1_LOC_748/A 0.12fF
C46049 NOR2X1_LOC_657/Y INVX1_LOC_5/A 0.00fF
C46050 NOR2X1_LOC_15/Y NOR2X1_LOC_82/A 0.07fF
C46051 NAND2X1_LOC_656/Y NAND2X1_LOC_74/B 0.19fF
C46052 INVX1_LOC_144/A NAND2X1_LOC_798/B 0.16fF
C46053 NOR2X1_LOC_595/Y NOR2X1_LOC_536/A 0.01fF
C46054 NOR2X1_LOC_272/Y NOR2X1_LOC_441/Y 0.24fF
C46055 NAND2X1_LOC_11/Y NAND2X1_LOC_3/B 0.06fF
C46056 INVX1_LOC_75/A INVX1_LOC_123/Y 0.03fF
C46057 NAND2X1_LOC_573/A NOR2X1_LOC_89/A 0.00fF
C46058 NAND2X1_LOC_807/Y NOR2X1_LOC_653/Y 0.10fF
C46059 INVX1_LOC_50/A NAND2X1_LOC_361/Y 0.07fF
C46060 INVX1_LOC_11/A NOR2X1_LOC_361/B 0.17fF
C46061 NOR2X1_LOC_528/a_36_216# NOR2X1_LOC_89/A 0.00fF
C46062 NOR2X1_LOC_590/A NAND2X1_LOC_573/Y 0.00fF
C46063 NOR2X1_LOC_210/B NOR2X1_LOC_467/A 0.48fF
C46064 NAND2X1_LOC_650/B NOR2X1_LOC_176/a_36_216# 0.01fF
C46065 INVX1_LOC_223/Y INVX1_LOC_223/A 0.04fF
C46066 INVX1_LOC_256/A NOR2X1_LOC_205/Y 0.12fF
C46067 INVX1_LOC_266/A INVX1_LOC_292/A 0.12fF
C46068 GATE_741 NAND2X1_LOC_741/B 0.00fF
C46069 INVX1_LOC_255/Y INVX1_LOC_15/A 0.08fF
C46070 INVX1_LOC_13/A INVX1_LOC_3/Y 0.17fF
C46071 NOR2X1_LOC_83/a_36_216# NAND2X1_LOC_572/B 0.01fF
C46072 NOR2X1_LOC_398/Y INVX1_LOC_23/Y 0.03fF
C46073 NOR2X1_LOC_558/A INVX1_LOC_12/Y 0.10fF
C46074 NAND2X1_LOC_807/Y INVX1_LOC_19/A 0.20fF
C46075 NOR2X1_LOC_824/Y INVX1_LOC_38/A 0.09fF
C46076 INVX1_LOC_17/A INVX1_LOC_246/A 0.07fF
C46077 NOR2X1_LOC_486/Y INVX1_LOC_9/A 0.26fF
C46078 NOR2X1_LOC_405/A INVX1_LOC_54/A 0.14fF
C46079 INVX1_LOC_179/Y INVX1_LOC_18/Y 0.31fF
C46080 NOR2X1_LOC_92/Y NAND2X1_LOC_741/B 0.07fF
C46081 NOR2X1_LOC_613/Y INVX1_LOC_217/A 0.05fF
C46082 NOR2X1_LOC_45/B INVX1_LOC_92/A 0.37fF
C46083 INVX1_LOC_64/Y NOR2X1_LOC_342/B 0.02fF
C46084 INVX1_LOC_15/Y NOR2X1_LOC_19/a_36_216# 0.00fF
C46085 INVX1_LOC_38/A INVX1_LOC_76/A 1.44fF
C46086 INVX1_LOC_16/A INVX1_LOC_94/Y 0.03fF
C46087 INVX1_LOC_290/A NOR2X1_LOC_158/B 0.00fF
C46088 INPUT_0 INVX1_LOC_63/A 0.35fF
C46089 VDD NOR2X1_LOC_376/Y 0.12fF
C46090 D_INPUT_0 INVX1_LOC_251/A 0.00fF
C46091 INVX1_LOC_194/A NOR2X1_LOC_476/B 0.02fF
C46092 INVX1_LOC_59/A INVX1_LOC_61/A 0.10fF
C46093 INVX1_LOC_27/A INVX1_LOC_24/A 0.13fF
C46094 NAND2X1_LOC_343/a_36_24# INVX1_LOC_94/Y 0.00fF
C46095 INVX1_LOC_161/Y INVX1_LOC_31/A 0.05fF
C46096 NOR2X1_LOC_824/A INVX1_LOC_24/A 0.03fF
C46097 NOR2X1_LOC_71/Y INVX1_LOC_15/A 0.03fF
C46098 NOR2X1_LOC_567/B INVX1_LOC_69/A 0.08fF
C46099 INVX1_LOC_224/Y NAND2X1_LOC_338/B 0.05fF
C46100 INVX1_LOC_13/Y NOR2X1_LOC_537/A 0.00fF
C46101 NOR2X1_LOC_795/Y INVX1_LOC_53/A 0.01fF
C46102 NOR2X1_LOC_78/A NOR2X1_LOC_688/a_36_216# 0.00fF
C46103 NOR2X1_LOC_510/Y NOR2X1_LOC_433/A 0.95fF
C46104 NAND2X1_LOC_860/A NOR2X1_LOC_709/A 0.07fF
C46105 INVX1_LOC_199/Y INVX1_LOC_92/A 0.01fF
C46106 INVX1_LOC_115/Y NAND2X1_LOC_93/B 0.01fF
C46107 INVX1_LOC_13/Y NOR2X1_LOC_716/B 0.07fF
C46108 INVX1_LOC_7/A NAND2X1_LOC_223/A 0.03fF
C46109 NOR2X1_LOC_448/Y NOR2X1_LOC_596/A 0.05fF
C46110 NOR2X1_LOC_745/Y INVX1_LOC_30/A 0.06fF
C46111 NOR2X1_LOC_103/Y INVX1_LOC_72/A 0.13fF
C46112 NOR2X1_LOC_815/A INVX1_LOC_272/A 0.01fF
C46113 INVX1_LOC_6/A INVX1_LOC_19/A 0.10fF
C46114 INVX1_LOC_269/A INVX1_LOC_181/Y 0.01fF
C46115 INVX1_LOC_115/Y NAND2X1_LOC_425/Y 0.01fF
C46116 NAND2X1_LOC_642/Y INVX1_LOC_285/A 0.07fF
C46117 NOR2X1_LOC_553/Y NOR2X1_LOC_383/B 0.01fF
C46118 INVX1_LOC_280/Y NAND2X1_LOC_804/A 0.00fF
C46119 INPUT_1 NOR2X1_LOC_38/B 0.04fF
C46120 NAND2X1_LOC_859/B INVX1_LOC_57/A 0.46fF
C46121 NOR2X1_LOC_294/a_36_216# INVX1_LOC_31/A 0.01fF
C46122 NOR2X1_LOC_510/Y INVX1_LOC_151/A 0.03fF
C46123 NAND2X1_LOC_623/B NAND2X1_LOC_489/Y 0.08fF
C46124 NOR2X1_LOC_828/B INVX1_LOC_15/A 0.01fF
C46125 INVX1_LOC_285/Y NOR2X1_LOC_89/A 0.01fF
C46126 NOR2X1_LOC_614/Y INVX1_LOC_53/A 0.06fF
C46127 INVX1_LOC_136/A INVX1_LOC_39/Y 0.01fF
C46128 NOR2X1_LOC_510/Y NOR2X1_LOC_52/B 0.18fF
C46129 NOR2X1_LOC_361/B NOR2X1_LOC_433/A 0.31fF
C46130 NOR2X1_LOC_602/A INVX1_LOC_30/A 0.05fF
C46131 INVX1_LOC_50/A NAND2X1_LOC_319/A 0.04fF
C46132 NOR2X1_LOC_420/Y INVX1_LOC_2/A 0.07fF
C46133 INVX1_LOC_28/A INVX1_LOC_94/Y 2.03fF
C46134 INVX1_LOC_45/A INVX1_LOC_72/A 0.10fF
C46135 INVX1_LOC_281/A INVX1_LOC_92/A 0.13fF
C46136 INVX1_LOC_136/A INVX1_LOC_312/Y 0.10fF
C46137 NOR2X1_LOC_94/a_36_216# NOR2X1_LOC_392/Y 0.01fF
C46138 INVX1_LOC_46/A NAND2X1_LOC_771/a_36_24# 0.01fF
C46139 NAND2X1_LOC_86/Y INVX1_LOC_29/A 0.01fF
C46140 NAND2X1_LOC_341/A INVX1_LOC_64/A 0.09fF
C46141 INVX1_LOC_72/A NAND2X1_LOC_856/A 0.03fF
C46142 INVX1_LOC_255/Y NOR2X1_LOC_818/a_36_216# 0.00fF
C46143 NOR2X1_LOC_130/A INVX1_LOC_271/A 0.03fF
C46144 INVX1_LOC_27/A INVX1_LOC_143/A 0.00fF
C46145 NAND2X1_LOC_217/a_36_24# NAND2X1_LOC_555/Y 0.01fF
C46146 INVX1_LOC_11/A INVX1_LOC_153/Y 0.01fF
C46147 NAND2X1_LOC_861/Y INVX1_LOC_57/A 0.07fF
C46148 INVX1_LOC_45/A INVX1_LOC_198/Y 0.03fF
C46149 NAND2X1_LOC_563/Y INVX1_LOC_269/A -0.02fF
C46150 NOR2X1_LOC_405/A NAND2X1_LOC_807/B 0.01fF
C46151 NOR2X1_LOC_150/a_36_216# INVX1_LOC_57/A 0.00fF
C46152 NOR2X1_LOC_361/B NOR2X1_LOC_52/B 0.18fF
C46153 NOR2X1_LOC_658/Y NOR2X1_LOC_759/Y 0.56fF
C46154 NOR2X1_LOC_389/A INVX1_LOC_49/A 0.21fF
C46155 INVX1_LOC_256/A NOR2X1_LOC_843/A 0.05fF
C46156 INVX1_LOC_132/A NOR2X1_LOC_590/A 0.07fF
C46157 NAND2X1_LOC_581/Y INVX1_LOC_11/A 0.01fF
C46158 INVX1_LOC_245/Y INVX1_LOC_63/Y 0.01fF
C46159 NAND2X1_LOC_770/a_36_24# NAND2X1_LOC_770/Y 0.00fF
C46160 INVX1_LOC_37/A NOR2X1_LOC_691/B 0.03fF
C46161 NAND2X1_LOC_9/Y INVX1_LOC_135/A 0.06fF
C46162 INVX1_LOC_11/A INVX1_LOC_121/Y 0.09fF
C46163 INVX1_LOC_226/Y NAND2X1_LOC_391/Y 0.12fF
C46164 INVX1_LOC_132/A INVX1_LOC_22/Y 0.03fF
C46165 INVX1_LOC_69/Y INVX1_LOC_4/Y 0.08fF
C46166 INVX1_LOC_2/A NAND2X1_LOC_190/Y 0.07fF
C46167 INVX1_LOC_233/A INVX1_LOC_135/A 0.10fF
C46168 NOR2X1_LOC_226/A NOR2X1_LOC_468/Y 0.09fF
C46169 INVX1_LOC_58/A INVX1_LOC_55/Y 0.08fF
C46170 INVX1_LOC_72/A INVX1_LOC_71/A 0.16fF
C46171 INVX1_LOC_12/A NOR2X1_LOC_603/Y 0.08fF
C46172 INVX1_LOC_36/A NOR2X1_LOC_643/Y 0.73fF
C46173 NAND2X1_LOC_721/B INVX1_LOC_172/A 0.32fF
C46174 INVX1_LOC_11/A INVX1_LOC_177/A 0.03fF
C46175 NOR2X1_LOC_82/A NAND2X1_LOC_141/A 0.08fF
C46176 NAND2X1_LOC_9/Y NOR2X1_LOC_560/A 0.04fF
C46177 INVX1_LOC_225/A NOR2X1_LOC_590/A 0.00fF
C46178 NOR2X1_LOC_15/Y INVX1_LOC_278/Y 0.10fF
C46179 NOR2X1_LOC_89/A NAND2X1_LOC_267/B 0.34fF
C46180 NAND2X1_LOC_149/Y INVX1_LOC_268/Y 0.03fF
C46181 NOR2X1_LOC_103/Y NOR2X1_LOC_537/Y 0.01fF
C46182 INVX1_LOC_88/A NOR2X1_LOC_757/Y 0.09fF
C46183 INVX1_LOC_33/A NOR2X1_LOC_169/B 0.01fF
C46184 NAND2X1_LOC_338/B NOR2X1_LOC_103/Y 0.75fF
C46185 NOR2X1_LOC_216/Y INVX1_LOC_271/A 0.00fF
C46186 INVX1_LOC_1/A NOR2X1_LOC_210/B 0.65fF
C46187 NOR2X1_LOC_317/A INVX1_LOC_49/A 0.07fF
C46188 INVX1_LOC_131/Y NAND2X1_LOC_288/A 0.02fF
C46189 NOR2X1_LOC_226/A NAND2X1_LOC_396/a_36_24# 0.00fF
C46190 INVX1_LOC_11/A NOR2X1_LOC_547/a_36_216# 0.00fF
C46191 INVX1_LOC_249/A INVX1_LOC_24/A 0.07fF
C46192 NOR2X1_LOC_178/Y INVX1_LOC_90/A 0.18fF
C46193 INVX1_LOC_36/A NAND2X1_LOC_811/Y 0.03fF
C46194 NOR2X1_LOC_540/B INVX1_LOC_15/A 0.03fF
C46195 VDD NAND2X1_LOC_254/Y 0.72fF
C46196 NOR2X1_LOC_798/A INVX1_LOC_135/A 0.03fF
C46197 NOR2X1_LOC_635/A NAND2X1_LOC_36/A 0.01fF
C46198 INVX1_LOC_174/Y INVX1_LOC_198/A 0.01fF
C46199 INVX1_LOC_134/A NAND2X1_LOC_290/a_36_24# 0.00fF
C46200 INVX1_LOC_49/A INVX1_LOC_62/Y 0.02fF
C46201 INVX1_LOC_2/A NOR2X1_LOC_389/A 0.10fF
C46202 INVX1_LOC_120/A INVX1_LOC_50/Y 0.15fF
C46203 NOR2X1_LOC_67/A NOR2X1_LOC_160/B 0.07fF
C46204 NAND2X1_LOC_276/Y NOR2X1_LOC_68/A 0.03fF
C46205 NOR2X1_LOC_590/A NOR2X1_LOC_209/Y 0.08fF
C46206 INVX1_LOC_84/A NAND2X1_LOC_243/Y 0.03fF
C46207 NOR2X1_LOC_230/a_36_216# INVX1_LOC_266/Y 0.00fF
C46208 INVX1_LOC_49/A NOR2X1_LOC_596/A 1.50fF
C46209 NAND2X1_LOC_364/A NOR2X1_LOC_142/Y 0.06fF
C46210 INVX1_LOC_37/A NOR2X1_LOC_477/B 0.01fF
C46211 NAND2X1_LOC_229/a_36_24# NOR2X1_LOC_160/B 0.00fF
C46212 INVX1_LOC_5/A NOR2X1_LOC_356/A 0.07fF
C46213 INVX1_LOC_21/A NOR2X1_LOC_76/A 0.05fF
C46214 INVX1_LOC_135/A NAND2X1_LOC_703/Y 0.10fF
C46215 INVX1_LOC_17/A INVX1_LOC_290/A 0.03fF
C46216 INVX1_LOC_64/A NAND2X1_LOC_740/B 0.04fF
C46217 INVX1_LOC_36/A INVX1_LOC_266/Y 0.06fF
C46218 NAND2X1_LOC_192/B NOR2X1_LOC_665/A 0.01fF
C46219 INVX1_LOC_64/A NOR2X1_LOC_256/Y 0.01fF
C46220 INVX1_LOC_280/A NOR2X1_LOC_671/Y 0.02fF
C46221 NOR2X1_LOC_94/Y NOR2X1_LOC_671/Y 0.01fF
C46222 INVX1_LOC_21/A NOR2X1_LOC_180/B 0.07fF
C46223 NOR2X1_LOC_331/B NOR2X1_LOC_755/Y -0.10fF
C46224 INVX1_LOC_235/Y NAND2X1_LOC_624/A 0.02fF
C46225 NOR2X1_LOC_15/Y INVX1_LOC_306/A 0.02fF
C46226 NOR2X1_LOC_454/Y INVX1_LOC_89/A 0.08fF
C46227 INVX1_LOC_303/A NOR2X1_LOC_716/B 0.02fF
C46228 INVX1_LOC_45/A NAND2X1_LOC_338/B 2.03fF
C46229 INVX1_LOC_62/Y INVX1_LOC_60/A 0.05fF
C46230 NAND2X1_LOC_632/B NAND2X1_LOC_631/a_36_24# 0.02fF
C46231 INVX1_LOC_106/Y INVX1_LOC_9/A 0.01fF
C46232 NAND2X1_LOC_559/Y NOR2X1_LOC_380/A 0.03fF
C46233 INVX1_LOC_131/Y INVX1_LOC_19/A 0.04fF
C46234 INVX1_LOC_11/A NAND2X1_LOC_573/A 0.03fF
C46235 INVX1_LOC_45/A NAND2X1_LOC_323/B 3.14fF
C46236 INVX1_LOC_32/A INVX1_LOC_117/A 0.30fF
C46237 NOR2X1_LOC_216/B NAND2X1_LOC_773/B 0.07fF
C46238 NAND2X1_LOC_219/a_36_24# INVX1_LOC_83/A 0.00fF
C46239 NOR2X1_LOC_718/B NOR2X1_LOC_303/Y 0.01fF
C46240 NOR2X1_LOC_655/B NAND2X1_LOC_364/A 0.10fF
C46241 NAND2X1_LOC_366/A NAND2X1_LOC_367/A 0.02fF
C46242 INVX1_LOC_109/Y INVX1_LOC_54/A 0.07fF
C46243 NOR2X1_LOC_468/Y INPUT_1 1.97fF
C46244 INVX1_LOC_5/A NOR2X1_LOC_74/A 0.52fF
C46245 NOR2X1_LOC_808/A NOR2X1_LOC_325/Y 0.01fF
C46246 NAND2X1_LOC_63/Y NOR2X1_LOC_624/B 0.06fF
C46247 INVX1_LOC_2/A INVX1_LOC_62/Y 0.10fF
C46248 NAND2X1_LOC_266/a_36_24# INVX1_LOC_87/A 0.00fF
C46249 INVX1_LOC_14/Y INVX1_LOC_271/Y 0.10fF
C46250 INVX1_LOC_21/A INVX1_LOC_73/A 0.03fF
C46251 NOR2X1_LOC_208/Y INVX1_LOC_266/Y 0.10fF
C46252 NAND2X1_LOC_465/A NAND2X1_LOC_99/A 0.02fF
C46253 INVX1_LOC_2/A NOR2X1_LOC_596/A 0.06fF
C46254 INVX1_LOC_44/A INVX1_LOC_4/A 0.08fF
C46255 NOR2X1_LOC_100/A NOR2X1_LOC_860/B 0.05fF
C46256 NOR2X1_LOC_13/Y NOR2X1_LOC_41/Y 0.04fF
C46257 NOR2X1_LOC_45/B INVX1_LOC_53/A 0.10fF
C46258 INVX1_LOC_71/A NAND2X1_LOC_633/a_36_24# 0.00fF
C46259 NOR2X1_LOC_276/Y NAND2X1_LOC_656/Y 0.03fF
C46260 NOR2X1_LOC_703/B NOR2X1_LOC_500/Y 0.32fF
C46261 INVX1_LOC_5/A NOR2X1_LOC_9/Y 0.03fF
C46262 INVX1_LOC_161/Y INVX1_LOC_313/A 0.02fF
C46263 NAND2X1_LOC_785/Y NAND2X1_LOC_833/Y 0.04fF
C46264 INVX1_LOC_178/A NOR2X1_LOC_74/A 0.03fF
C46265 NOR2X1_LOC_574/a_36_216# NOR2X1_LOC_577/Y 0.01fF
C46266 NAND2X1_LOC_338/B INVX1_LOC_71/A 0.78fF
C46267 INVX1_LOC_41/A NAND2X1_LOC_116/A 0.00fF
C46268 NOR2X1_LOC_716/B INVX1_LOC_168/A 0.04fF
C46269 NAND2X1_LOC_112/Y INVX1_LOC_177/Y 0.16fF
C46270 NOR2X1_LOC_593/Y INVX1_LOC_177/A 0.03fF
C46271 NOR2X1_LOC_38/B INVX1_LOC_118/A 0.09fF
C46272 NAND2X1_LOC_85/Y NAND2X1_LOC_206/B 0.01fF
C46273 NAND2X1_LOC_243/Y INVX1_LOC_15/A 0.05fF
C46274 INVX1_LOC_49/A INVX1_LOC_189/Y 0.01fF
C46275 INVX1_LOC_77/A NOR2X1_LOC_524/a_36_216# 0.00fF
C46276 NAND2X1_LOC_741/B NOR2X1_LOC_299/Y 0.03fF
C46277 NAND2X1_LOC_453/A INVX1_LOC_296/Y 0.09fF
C46278 NAND2X1_LOC_93/B D_INPUT_5 0.08fF
C46279 INVX1_LOC_58/A NOR2X1_LOC_357/Y 0.10fF
C46280 NOR2X1_LOC_220/A INVX1_LOC_49/A 0.03fF
C46281 INVX1_LOC_24/A NOR2X1_LOC_695/Y 0.06fF
C46282 NAND2X1_LOC_387/a_36_24# INVX1_LOC_89/A 0.00fF
C46283 NAND2X1_LOC_387/B INVX1_LOC_83/A 0.03fF
C46284 NOR2X1_LOC_667/A NAND2X1_LOC_833/Y 0.02fF
C46285 INVX1_LOC_8/A INVX1_LOC_34/Y 0.43fF
C46286 INVX1_LOC_33/A INVX1_LOC_179/Y 0.02fF
C46287 INVX1_LOC_248/A NAND2X1_LOC_833/Y 0.01fF
C46288 NAND2X1_LOC_425/Y D_INPUT_5 0.04fF
C46289 NOR2X1_LOC_569/Y NOR2X1_LOC_303/Y 0.23fF
C46290 NOR2X1_LOC_596/A NAND2X1_LOC_664/a_36_24# 0.01fF
C46291 NOR2X1_LOC_122/A INVX1_LOC_6/A 0.03fF
C46292 NAND2X1_LOC_474/Y INVX1_LOC_91/A 0.10fF
C46293 INVX1_LOC_45/A INVX1_LOC_313/Y 0.03fF
C46294 NOR2X1_LOC_793/a_36_216# INVX1_LOC_33/A 0.00fF
C46295 INPUT_2 INVX1_LOC_75/A 0.09fF
C46296 NAND2X1_LOC_34/a_36_24# INVX1_LOC_240/A 0.01fF
C46297 INVX1_LOC_294/Y NOR2X1_LOC_773/Y 0.52fF
C46298 INVX1_LOC_64/A NOR2X1_LOC_331/a_36_216# 0.01fF
C46299 NAND2X1_LOC_383/a_36_24# NOR2X1_LOC_536/A 0.00fF
C46300 INVX1_LOC_41/A INVX1_LOC_232/A 0.03fF
C46301 NAND2X1_LOC_612/a_36_24# INVX1_LOC_75/A 0.00fF
C46302 NOR2X1_LOC_524/Y INVX1_LOC_28/A 0.01fF
C46303 INVX1_LOC_33/A NOR2X1_LOC_719/A 0.00fF
C46304 NOR2X1_LOC_816/A NOR2X1_LOC_74/A 0.11fF
C46305 INVX1_LOC_35/A INVX1_LOC_37/A 0.13fF
C46306 NOR2X1_LOC_798/A NOR2X1_LOC_566/a_36_216# 0.00fF
C46307 INVX1_LOC_30/A NOR2X1_LOC_564/Y 0.07fF
C46308 INVX1_LOC_34/A INVX1_LOC_1/Y 0.07fF
C46309 INVX1_LOC_24/Y INVX1_LOC_186/A 0.03fF
C46310 INVX1_LOC_215/Y NOR2X1_LOC_320/Y 0.01fF
C46311 NOR2X1_LOC_89/A NAND2X1_LOC_81/B 0.04fF
C46312 INVX1_LOC_161/Y INVX1_LOC_6/A 0.21fF
C46313 INVX1_LOC_9/A NOR2X1_LOC_748/A 0.03fF
C46314 INVX1_LOC_3/Y NAND2X1_LOC_489/Y 0.39fF
C46315 INVX1_LOC_41/A NOR2X1_LOC_383/Y 0.72fF
C46316 NAND2X1_LOC_660/Y INVX1_LOC_63/Y 0.03fF
C46317 INVX1_LOC_77/A INVX1_LOC_150/A 0.16fF
C46318 NOR2X1_LOC_561/Y INVX1_LOC_33/A 0.18fF
C46319 NOR2X1_LOC_831/B NOR2X1_LOC_278/Y 0.07fF
C46320 NOR2X1_LOC_315/Y INVX1_LOC_16/A 0.04fF
C46321 NAND2X1_LOC_112/Y INVX1_LOC_104/A 0.03fF
C46322 INVX1_LOC_223/A INVX1_LOC_75/A 0.17fF
C46323 NOR2X1_LOC_644/Y INVX1_LOC_263/A 0.04fF
C46324 NOR2X1_LOC_226/A NAND2X1_LOC_395/a_36_24# 0.01fF
C46325 NOR2X1_LOC_742/A NOR2X1_LOC_722/Y 0.03fF
C46326 INVX1_LOC_89/A INVX1_LOC_77/A 5.97fF
C46327 INVX1_LOC_36/A INVX1_LOC_42/Y 0.01fF
C46328 INVX1_LOC_313/Y INVX1_LOC_71/A 0.07fF
C46329 NAND2X1_LOC_53/Y INVX1_LOC_91/A 0.51fF
C46330 INVX1_LOC_53/A NOR2X1_LOC_499/B 0.00fF
C46331 NAND2X1_LOC_198/B NOR2X1_LOC_329/B 0.10fF
C46332 INVX1_LOC_269/A NOR2X1_LOC_675/A 0.04fF
C46333 NOR2X1_LOC_411/A INVX1_LOC_38/A 0.01fF
C46334 NOR2X1_LOC_274/Y NOR2X1_LOC_389/B 0.06fF
C46335 INVX1_LOC_57/A INVX1_LOC_291/A 0.07fF
C46336 NOR2X1_LOC_561/Y NAND2X1_LOC_466/A 0.05fF
C46337 INVX1_LOC_24/A NOR2X1_LOC_19/B 0.00fF
C46338 NOR2X1_LOC_432/Y INVX1_LOC_16/A 0.09fF
C46339 NOR2X1_LOC_252/Y NOR2X1_LOC_482/Y 0.01fF
C46340 NOR2X1_LOC_97/A NAND2X1_LOC_351/A 0.21fF
C46341 NOR2X1_LOC_219/Y NOR2X1_LOC_222/Y 0.05fF
C46342 INVX1_LOC_64/A NOR2X1_LOC_96/a_36_216# 0.00fF
C46343 INVX1_LOC_59/A D_INPUT_3 0.01fF
C46344 INVX1_LOC_299/A NOR2X1_LOC_35/Y 0.10fF
C46345 NAND2X1_LOC_803/B NAND2X1_LOC_643/a_36_24# 0.01fF
C46346 INVX1_LOC_35/Y NAND2X1_LOC_464/B 0.19fF
C46347 INVX1_LOC_84/A INVX1_LOC_16/Y 0.01fF
C46348 NAND2X1_LOC_564/B NAND2X1_LOC_181/Y 0.06fF
C46349 INVX1_LOC_89/A NOR2X1_LOC_732/A 0.00fF
C46350 NOR2X1_LOC_795/Y INVX1_LOC_83/A 0.03fF
C46351 INVX1_LOC_124/A INVX1_LOC_150/A 0.06fF
C46352 NAND2X1_LOC_773/Y INVX1_LOC_14/Y 0.00fF
C46353 INVX1_LOC_120/A NOR2X1_LOC_6/B -0.00fF
C46354 NAND2X1_LOC_513/B NAND2X1_LOC_472/Y 0.01fF
C46355 NOR2X1_LOC_208/Y INVX1_LOC_42/Y 0.00fF
C46356 NOR2X1_LOC_590/A NAND2X1_LOC_642/Y 0.12fF
C46357 INVX1_LOC_35/A NOR2X1_LOC_743/Y 0.18fF
C46358 NAND2X1_LOC_579/A NOR2X1_LOC_111/A 0.04fF
C46359 INVX1_LOC_53/A NOR2X1_LOC_862/B 0.45fF
C46360 INVX1_LOC_183/A INVX1_LOC_63/A 0.00fF
C46361 INVX1_LOC_41/A NOR2X1_LOC_775/Y 0.02fF
C46362 INVX1_LOC_23/A NOR2X1_LOC_841/A 0.01fF
C46363 NOR2X1_LOC_561/Y NAND2X1_LOC_798/A 0.02fF
C46364 INVX1_LOC_159/A NAND2X1_LOC_661/a_36_24# 0.00fF
C46365 NOR2X1_LOC_441/Y NOR2X1_LOC_405/A 0.00fF
C46366 NOR2X1_LOC_399/Y NAND2X1_LOC_462/B 0.02fF
C46367 NOR2X1_LOC_89/A INVX1_LOC_4/Y 0.39fF
C46368 NOR2X1_LOC_748/Y INVX1_LOC_22/A 0.01fF
C46369 INVX1_LOC_7/A INVX1_LOC_40/A 0.07fF
C46370 INVX1_LOC_32/A INVX1_LOC_3/Y 0.22fF
C46371 INVX1_LOC_84/A NAND2X1_LOC_205/A 0.22fF
C46372 NOR2X1_LOC_483/B INVX1_LOC_76/A 0.02fF
C46373 INVX1_LOC_177/Y NOR2X1_LOC_78/A 0.07fF
C46374 INVX1_LOC_252/Y D_INPUT_3 0.01fF
C46375 NOR2X1_LOC_160/B NOR2X1_LOC_558/A 0.01fF
C46376 NOR2X1_LOC_716/B NOR2X1_LOC_83/a_36_216# 0.01fF
C46377 INVX1_LOC_82/A NAND2X1_LOC_293/a_36_24# 0.00fF
C46378 INVX1_LOC_58/A NAND2X1_LOC_489/Y 0.03fF
C46379 NOR2X1_LOC_427/a_36_216# INVX1_LOC_77/Y 0.01fF
C46380 INVX1_LOC_26/Y NOR2X1_LOC_633/A 0.01fF
C46381 INVX1_LOC_49/A INVX1_LOC_51/Y 0.00fF
C46382 INVX1_LOC_75/A INVX1_LOC_149/Y 0.00fF
C46383 INVX1_LOC_270/A INVX1_LOC_19/A 0.07fF
C46384 INVX1_LOC_24/A NOR2X1_LOC_528/Y 0.16fF
C46385 NOR2X1_LOC_355/A INVX1_LOC_208/Y 0.01fF
C46386 NOR2X1_LOC_218/A NOR2X1_LOC_363/Y 0.12fF
C46387 NOR2X1_LOC_170/A INVX1_LOC_4/Y 0.02fF
C46388 NAND2X1_LOC_395/a_36_24# INPUT_1 0.00fF
C46389 INVX1_LOC_85/A INVX1_LOC_75/A 0.03fF
C46390 NAND2X1_LOC_364/Y NOR2X1_LOC_334/A 0.03fF
C46391 NOR2X1_LOC_468/Y INVX1_LOC_118/A 0.00fF
C46392 NAND2X1_LOC_357/B NOR2X1_LOC_527/a_36_216# 0.00fF
C46393 NAND2X1_LOC_725/B NOR2X1_LOC_629/Y 0.03fF
C46394 INVX1_LOC_5/A NOR2X1_LOC_243/B 0.07fF
C46395 NOR2X1_LOC_416/A INVX1_LOC_19/A 0.07fF
C46396 NAND2X1_LOC_470/B D_INPUT_5 0.62fF
C46397 INVX1_LOC_89/A NOR2X1_LOC_687/Y 0.40fF
C46398 D_GATE_366 INVX1_LOC_22/A 0.02fF
C46399 INVX1_LOC_209/A NOR2X1_LOC_409/Y 0.01fF
C46400 NOR2X1_LOC_249/Y NAND2X1_LOC_574/A 0.08fF
C46401 INVX1_LOC_234/A NOR2X1_LOC_130/A 0.16fF
C46402 INVX1_LOC_41/A INVX1_LOC_186/A 0.03fF
C46403 INVX1_LOC_89/A NOR2X1_LOC_549/a_36_216# 0.02fF
C46404 INVX1_LOC_174/A INVX1_LOC_193/A -0.03fF
C46405 INVX1_LOC_34/A NOR2X1_LOC_318/B 0.07fF
C46406 NAND2X1_LOC_714/B NOR2X1_LOC_697/Y 0.01fF
C46407 INVX1_LOC_19/A NOR2X1_LOC_109/Y 0.11fF
C46408 NOR2X1_LOC_590/A NOR2X1_LOC_271/Y 0.01fF
C46409 NAND2X1_LOC_359/Y NAND2X1_LOC_359/A 0.61fF
C46410 NOR2X1_LOC_160/B NOR2X1_LOC_729/A 0.05fF
C46411 NAND2X1_LOC_546/a_36_24# INVX1_LOC_118/A 0.00fF
C46412 NOR2X1_LOC_773/Y NOR2X1_LOC_74/A 0.29fF
C46413 INVX1_LOC_131/A INVX1_LOC_1/Y 0.16fF
C46414 NOR2X1_LOC_860/B INVX1_LOC_176/A 0.01fF
C46415 NOR2X1_LOC_142/Y NOR2X1_LOC_405/A 0.11fF
C46416 NOR2X1_LOC_160/B NAND2X1_LOC_268/a_36_24# 0.00fF
C46417 INVX1_LOC_34/A INVX1_LOC_93/Y 0.07fF
C46418 INVX1_LOC_104/A NOR2X1_LOC_78/A 0.17fF
C46419 NOR2X1_LOC_837/B INVX1_LOC_37/A 0.02fF
C46420 NOR2X1_LOC_596/A NAND2X1_LOC_605/a_36_24# 0.00fF
C46421 INVX1_LOC_41/A NAND2X1_LOC_447/Y 0.02fF
C46422 NOR2X1_LOC_773/Y NOR2X1_LOC_9/Y 0.10fF
C46423 INVX1_LOC_181/Y INVX1_LOC_12/Y 0.01fF
C46424 INVX1_LOC_58/A INVX1_LOC_32/A 0.54fF
C46425 INVX1_LOC_314/Y VDD 1.66fF
C46426 NOR2X1_LOC_420/Y NAND2X1_LOC_63/Y 0.01fF
C46427 INVX1_LOC_201/Y INVX1_LOC_74/Y 0.01fF
C46428 INVX1_LOC_72/A NOR2X1_LOC_331/B 0.07fF
C46429 INVX1_LOC_1/Y INPUT_0 0.11fF
C46430 NOR2X1_LOC_360/Y NOR2X1_LOC_536/A 0.03fF
C46431 INVX1_LOC_33/A INVX1_LOC_76/A 1.02fF
C46432 NOR2X1_LOC_778/B NOR2X1_LOC_337/Y 0.23fF
C46433 NAND2X1_LOC_208/a_36_24# INVX1_LOC_12/A 0.01fF
C46434 NOR2X1_LOC_75/Y INVX1_LOC_107/Y 0.33fF
C46435 NOR2X1_LOC_19/B NOR2X1_LOC_130/A 0.46fF
C46436 NAND2X1_LOC_640/Y NAND2X1_LOC_650/B -0.01fF
C46437 NOR2X1_LOC_303/Y NAND2X1_LOC_472/Y 0.07fF
C46438 INVX1_LOC_128/A INVX1_LOC_23/A 0.02fF
C46439 NOR2X1_LOC_78/B NOR2X1_LOC_45/B 0.80fF
C46440 NOR2X1_LOC_516/B NOR2X1_LOC_551/Y 0.01fF
C46441 INVX1_LOC_34/A INVX1_LOC_139/A 1.84fF
C46442 INVX1_LOC_306/Y INVX1_LOC_42/A 0.11fF
C46443 NAND2X1_LOC_725/Y NOR2X1_LOC_409/B 0.03fF
C46444 NOR2X1_LOC_817/Y INVX1_LOC_84/A 0.00fF
C46445 NOR2X1_LOC_828/Y NOR2X1_LOC_855/A 0.03fF
C46446 NOR2X1_LOC_703/Y NOR2X1_LOC_687/Y 0.16fF
C46447 NOR2X1_LOC_655/B NOR2X1_LOC_405/A 0.05fF
C46448 NAND2X1_LOC_231/Y INVX1_LOC_93/Y 0.21fF
C46449 D_INPUT_1 INVX1_LOC_165/A 0.01fF
C46450 NOR2X1_LOC_321/Y INVX1_LOC_29/A 0.07fF
C46451 NOR2X1_LOC_569/A NOR2X1_LOC_565/B 0.23fF
C46452 INVX1_LOC_289/Y INVX1_LOC_49/Y 0.17fF
C46453 NOR2X1_LOC_500/Y INVX1_LOC_91/A 0.19fF
C46454 NOR2X1_LOC_468/Y NAND2X1_LOC_63/Y 0.03fF
C46455 INVX1_LOC_58/A NAND2X1_LOC_175/Y 0.07fF
C46456 INVX1_LOC_138/A NOR2X1_LOC_38/B 0.01fF
C46457 NOR2X1_LOC_144/Y INVX1_LOC_14/Y 0.07fF
C46458 INVX1_LOC_226/Y INVX1_LOC_91/A 0.07fF
C46459 NAND2X1_LOC_348/A NAND2X1_LOC_45/Y 0.02fF
C46460 INVX1_LOC_34/A NAND2X1_LOC_721/A 0.05fF
C46461 NOR2X1_LOC_181/Y VDD 0.12fF
C46462 INVX1_LOC_2/A NAND2X1_LOC_469/B 0.05fF
C46463 NOR2X1_LOC_599/A NAND2X1_LOC_810/B 0.01fF
C46464 NOR2X1_LOC_78/B INVX1_LOC_247/A 0.03fF
C46465 NOR2X1_LOC_496/Y NOR2X1_LOC_754/A -0.00fF
C46466 NOR2X1_LOC_254/Y NAND2X1_LOC_472/Y 0.21fF
C46467 NOR2X1_LOC_270/Y INVX1_LOC_92/A 0.15fF
C46468 INVX1_LOC_257/Y INVX1_LOC_37/A 0.01fF
C46469 INVX1_LOC_35/A NAND2X1_LOC_72/B 0.03fF
C46470 INVX1_LOC_207/A NOR2X1_LOC_536/A 0.06fF
C46471 NOR2X1_LOC_703/B NOR2X1_LOC_445/B 0.01fF
C46472 INVX1_LOC_251/Y INVX1_LOC_46/A 0.04fF
C46473 INVX1_LOC_11/A NAND2X1_LOC_81/B 0.00fF
C46474 NOR2X1_LOC_468/Y NAND2X1_LOC_455/B 0.01fF
C46475 NOR2X1_LOC_718/a_36_216# INVX1_LOC_139/Y 0.00fF
C46476 NOR2X1_LOC_205/Y NOR2X1_LOC_89/A 0.03fF
C46477 NOR2X1_LOC_554/B NOR2X1_LOC_820/Y 0.70fF
C46478 NAND2X1_LOC_793/Y INVX1_LOC_29/A 0.06fF
C46479 NAND2X1_LOC_578/B INVX1_LOC_178/Y 0.02fF
C46480 NOR2X1_LOC_355/A NOR2X1_LOC_501/B 0.01fF
C46481 INVX1_LOC_10/A INVX1_LOC_91/A 0.17fF
C46482 INVX1_LOC_39/A NOR2X1_LOC_38/B 0.03fF
C46483 NAND2X1_LOC_855/Y NAND2X1_LOC_863/A 0.03fF
C46484 NOR2X1_LOC_792/B NOR2X1_LOC_536/A 0.01fF
C46485 INVX1_LOC_226/A INVX1_LOC_176/A 0.01fF
C46486 INVX1_LOC_40/A INVX1_LOC_76/A 0.07fF
C46487 NOR2X1_LOC_778/B VDD 0.47fF
C46488 INVX1_LOC_24/A NOR2X1_LOC_216/B 0.04fF
C46489 NOR2X1_LOC_226/A NOR2X1_LOC_447/B 0.01fF
C46490 INVX1_LOC_36/A NOR2X1_LOC_653/Y 0.39fF
C46491 NOR2X1_LOC_13/Y NOR2X1_LOC_13/a_36_216# 0.02fF
C46492 NOR2X1_LOC_770/A NAND2X1_LOC_93/B 0.05fF
C46493 INVX1_LOC_83/A NOR2X1_LOC_45/B 0.11fF
C46494 INVX1_LOC_140/A NOR2X1_LOC_74/A 0.03fF
C46495 INVX1_LOC_248/Y NAND2X1_LOC_175/Y 0.04fF
C46496 NAND2X1_LOC_860/A NAND2X1_LOC_464/B 0.11fF
C46497 NAND2X1_LOC_35/Y INVX1_LOC_23/Y 0.62fF
C46498 NOR2X1_LOC_383/B NOR2X1_LOC_678/A 0.03fF
C46499 NAND2X1_LOC_162/B INVX1_LOC_107/Y 0.01fF
C46500 NAND2X1_LOC_451/Y NAND2X1_LOC_639/A 0.10fF
C46501 NOR2X1_LOC_91/Y INVX1_LOC_265/Y 0.00fF
C46502 INVX1_LOC_10/A INVX1_LOC_11/Y 8.23fF
C46503 NOR2X1_LOC_383/B INVX1_LOC_295/Y 0.10fF
C46504 NOR2X1_LOC_607/A NAND2X1_LOC_606/a_36_24# 0.02fF
C46505 NOR2X1_LOC_770/A NAND2X1_LOC_425/Y 0.03fF
C46506 INVX1_LOC_36/A INVX1_LOC_19/A 0.10fF
C46507 NOR2X1_LOC_78/B INVX1_LOC_281/A 0.00fF
C46508 NOR2X1_LOC_798/A NOR2X1_LOC_541/B 0.00fF
C46509 INVX1_LOC_135/A NOR2X1_LOC_545/B 0.03fF
C46510 INVX1_LOC_34/A INVX1_LOC_117/Y 1.01fF
C46511 INVX1_LOC_36/A NOR2X1_LOC_11/Y 1.74fF
C46512 NOR2X1_LOC_296/Y INVX1_LOC_3/Y 0.03fF
C46513 NOR2X1_LOC_493/B INVX1_LOC_9/A 0.11fF
C46514 NOR2X1_LOC_557/Y NOR2X1_LOC_216/B 0.10fF
C46515 INVX1_LOC_229/Y NAND2X1_LOC_836/Y 0.03fF
C46516 INVX1_LOC_24/A NAND2X1_LOC_477/Y 0.01fF
C46517 NAND2X1_LOC_288/B NOR2X1_LOC_652/Y 0.08fF
C46518 INVX1_LOC_304/A NOR2X1_LOC_76/A 0.02fF
C46519 NAND2X1_LOC_366/A NOR2X1_LOC_865/Y 0.05fF
C46520 INVX1_LOC_279/A INVX1_LOC_14/Y 0.10fF
C46521 NOR2X1_LOC_68/A INVX1_LOC_125/A 0.18fF
C46522 INVX1_LOC_224/A INVX1_LOC_4/Y -0.01fF
C46523 INPUT_3 INVX1_LOC_3/Y 0.04fF
C46524 NOR2X1_LOC_723/Y NOR2X1_LOC_89/A 0.04fF
C46525 INVX1_LOC_11/A INVX1_LOC_4/Y 0.72fF
C46526 NAND2X1_LOC_200/B NOR2X1_LOC_16/a_36_216# 0.00fF
C46527 GATE_662 INVX1_LOC_117/A 0.02fF
C46528 NOR2X1_LOC_643/Y INVX1_LOC_63/A 0.02fF
C46529 NOR2X1_LOC_753/Y NOR2X1_LOC_605/A 0.03fF
C46530 NOR2X1_LOC_208/Y INVX1_LOC_19/A 0.03fF
C46531 INVX1_LOC_36/A NAND2X1_LOC_227/a_36_24# 0.00fF
C46532 NAND2X1_LOC_303/B VDD 0.04fF
C46533 INVX1_LOC_1/A NOR2X1_LOC_302/A 0.03fF
C46534 NAND2X1_LOC_231/Y INVX1_LOC_117/Y 0.02fF
C46535 NOR2X1_LOC_318/B INPUT_0 0.07fF
C46536 NOR2X1_LOC_13/Y NAND2X1_LOC_74/B 0.07fF
C46537 NOR2X1_LOC_237/Y INVX1_LOC_19/A 0.16fF
C46538 NOR2X1_LOC_6/B NAND2X1_LOC_659/A 0.11fF
C46539 INVX1_LOC_17/A INVX1_LOC_116/Y 0.02fF
C46540 NOR2X1_LOC_860/B NOR2X1_LOC_340/A 0.01fF
C46541 NOR2X1_LOC_724/Y VDD 0.31fF
C46542 NOR2X1_LOC_78/B NOR2X1_LOC_862/B 0.01fF
C46543 NOR2X1_LOC_804/B INVX1_LOC_19/A 0.07fF
C46544 NOR2X1_LOC_122/A INVX1_LOC_270/A 0.03fF
C46545 NOR2X1_LOC_309/Y NOR2X1_LOC_653/Y 0.03fF
C46546 INVX1_LOC_308/Y NAND2X1_LOC_286/B 0.01fF
C46547 INVX1_LOC_93/Y INPUT_0 0.18fF
C46548 NAND2X1_LOC_195/a_36_24# INVX1_LOC_117/Y 0.00fF
C46549 NAND2X1_LOC_352/B NOR2X1_LOC_278/Y 0.00fF
C46550 NOR2X1_LOC_561/Y NOR2X1_LOC_351/Y 0.01fF
C46551 INVX1_LOC_83/A NOR2X1_LOC_378/Y 0.03fF
C46552 NOR2X1_LOC_146/Y INVX1_LOC_75/Y 0.02fF
C46553 NAND2X1_LOC_123/Y VDD 0.08fF
C46554 NOR2X1_LOC_338/Y INVX1_LOC_32/A 0.01fF
C46555 NAND2X1_LOC_842/B NOR2X1_LOC_558/a_36_216# 0.00fF
C46556 INVX1_LOC_224/Y NOR2X1_LOC_103/Y 0.30fF
C46557 INVX1_LOC_182/Y INVX1_LOC_14/Y 0.01fF
C46558 NOR2X1_LOC_597/Y VDD 0.24fF
C46559 NOR2X1_LOC_309/Y INVX1_LOC_19/A 0.13fF
C46560 INVX1_LOC_161/Y INVX1_LOC_270/A 0.01fF
C46561 INVX1_LOC_30/A NOR2X1_LOC_158/Y 0.07fF
C46562 INVX1_LOC_89/A INVX1_LOC_9/A 0.64fF
C46563 INVX1_LOC_27/A INVX1_LOC_38/Y 0.22fF
C46564 NOR2X1_LOC_142/Y INVX1_LOC_109/Y 0.14fF
C46565 NOR2X1_LOC_705/B INVX1_LOC_23/A 0.01fF
C46566 NAND2X1_LOC_508/A INVX1_LOC_9/A 0.03fF
C46567 INPUT_0 NAND2X1_LOC_721/A 0.02fF
C46568 NOR2X1_LOC_224/Y NAND2X1_LOC_227/Y 0.00fF
C46569 NOR2X1_LOC_45/B NOR2X1_LOC_368/Y 0.03fF
C46570 INVX1_LOC_83/A NOR2X1_LOC_862/B 0.08fF
C46571 INVX1_LOC_25/A NAND2X1_LOC_555/Y 0.24fF
C46572 INVX1_LOC_230/Y NOR2X1_LOC_629/A 0.01fF
C46573 NOR2X1_LOC_403/a_36_216# NOR2X1_LOC_394/Y 0.00fF
C46574 INVX1_LOC_45/A INVX1_LOC_224/Y 0.08fF
C46575 INVX1_LOC_256/Y NAND2X1_LOC_74/B 0.03fF
C46576 NOR2X1_LOC_332/A NOR2X1_LOC_865/Y 0.02fF
C46577 INVX1_LOC_161/Y NOR2X1_LOC_109/Y 0.01fF
C46578 NOR2X1_LOC_332/A NOR2X1_LOC_243/B 0.02fF
C46579 NOR2X1_LOC_593/Y INVX1_LOC_4/Y 0.45fF
C46580 INVX1_LOC_230/Y NAND2X1_LOC_624/B 0.03fF
C46581 NOR2X1_LOC_557/A VDD 0.09fF
C46582 NOR2X1_LOC_45/B INVX1_LOC_46/A 2.24fF
C46583 NOR2X1_LOC_373/Y INVX1_LOC_84/A 0.03fF
C46584 D_INPUT_0 INVX1_LOC_27/Y 0.10fF
C46585 NOR2X1_LOC_755/a_36_216# INVX1_LOC_92/A 0.00fF
C46586 NAND2X1_LOC_650/B NAND2X1_LOC_642/Y 0.08fF
C46587 NOR2X1_LOC_778/Y INVX1_LOC_53/A 0.01fF
C46588 NOR2X1_LOC_486/Y INVX1_LOC_76/A 0.22fF
C46589 NOR2X1_LOC_52/Y INVX1_LOC_53/A 0.49fF
C46590 NOR2X1_LOC_657/B VDD 0.12fF
C46591 INVX1_LOC_136/A NOR2X1_LOC_717/A 0.10fF
C46592 INVX1_LOC_269/A NAND2X1_LOC_725/B 0.03fF
C46593 NOR2X1_LOC_810/A NOR2X1_LOC_856/B 0.02fF
C46594 INVX1_LOC_312/A NOR2X1_LOC_109/Y -0.08fF
C46595 NOR2X1_LOC_437/Y INVX1_LOC_270/A 0.68fF
C46596 NOR2X1_LOC_15/Y INVX1_LOC_103/A 0.24fF
C46597 D_INPUT_1 INVX1_LOC_45/Y 0.04fF
C46598 NOR2X1_LOC_216/Y NOR2X1_LOC_216/B 0.01fF
C46599 INVX1_LOC_17/A INVX1_LOC_1/A 0.13fF
C46600 NOR2X1_LOC_763/Y NOR2X1_LOC_48/Y 0.02fF
C46601 NOR2X1_LOC_335/A NOR2X1_LOC_383/B 0.08fF
C46602 INVX1_LOC_293/A INVX1_LOC_48/Y 0.01fF
C46603 INVX1_LOC_35/A NAND2X1_LOC_198/B 0.01fF
C46604 NAND2X1_LOC_357/B NOR2X1_LOC_278/Y 0.08fF
C46605 NOR2X1_LOC_285/A NAND2X1_LOC_364/Y 0.02fF
C46606 INVX1_LOC_278/A NOR2X1_LOC_238/a_36_216# -0.01fF
C46607 NAND2X1_LOC_465/Y INVX1_LOC_23/Y 0.02fF
C46608 NOR2X1_LOC_234/Y INVX1_LOC_23/Y 0.03fF
C46609 NOR2X1_LOC_471/Y INVX1_LOC_1/A 0.02fF
C46610 NOR2X1_LOC_65/B INVX1_LOC_294/Y 0.01fF
C46611 INVX1_LOC_71/A NAND2X1_LOC_793/B 0.08fF
C46612 NOR2X1_LOC_15/Y INVX1_LOC_292/A 0.03fF
C46613 NOR2X1_LOC_392/a_36_216# NOR2X1_LOC_99/Y 0.03fF
C46614 INVX1_LOC_135/A INVX1_LOC_284/A 0.16fF
C46615 NOR2X1_LOC_78/B NOR2X1_LOC_465/Y 0.02fF
C46616 NOR2X1_LOC_172/Y INVX1_LOC_23/A 0.02fF
C46617 NAND2X1_LOC_96/A NOR2X1_LOC_35/Y 0.10fF
C46618 NAND2X1_LOC_555/Y INVX1_LOC_1/A 0.11fF
C46619 NOR2X1_LOC_816/Y INVX1_LOC_76/A 0.11fF
C46620 NOR2X1_LOC_286/Y NOR2X1_LOC_160/B 0.07fF
C46621 NOR2X1_LOC_147/B INVX1_LOC_23/A 0.01fF
C46622 NOR2X1_LOC_455/Y INVX1_LOC_33/A 0.03fF
C46623 NOR2X1_LOC_392/B INVX1_LOC_23/A 0.07fF
C46624 INVX1_LOC_91/A INVX1_LOC_307/A 0.07fF
C46625 INVX1_LOC_93/A INVX1_LOC_24/A 0.07fF
C46626 NAND2X1_LOC_16/a_36_24# INVX1_LOC_1/A 0.01fF
C46627 NOR2X1_LOC_520/A NOR2X1_LOC_843/B 0.02fF
C46628 NOR2X1_LOC_324/B NOR2X1_LOC_729/A 0.01fF
C46629 INVX1_LOC_36/A NOR2X1_LOC_122/A 0.01fF
C46630 INVX1_LOC_243/A NOR2X1_LOC_635/B 0.02fF
C46631 NOR2X1_LOC_373/Y INVX1_LOC_15/A 0.01fF
C46632 INVX1_LOC_91/A NOR2X1_LOC_445/B 0.08fF
C46633 INVX1_LOC_27/A NOR2X1_LOC_191/B 0.10fF
C46634 NOR2X1_LOC_178/Y INVX1_LOC_33/A 0.19fF
C46635 NOR2X1_LOC_208/A INVX1_LOC_19/A 0.01fF
C46636 NOR2X1_LOC_351/Y INVX1_LOC_76/A 0.12fF
C46637 NOR2X1_LOC_356/A INVX1_LOC_42/A 0.05fF
C46638 NOR2X1_LOC_76/A INVX1_LOC_19/Y 0.29fF
C46639 INVX1_LOC_286/A INVX1_LOC_84/A 0.07fF
C46640 NOR2X1_LOC_180/Y INVX1_LOC_53/A 0.03fF
C46641 NOR2X1_LOC_68/A NOR2X1_LOC_140/A 0.01fF
C46642 NOR2X1_LOC_764/Y D_INPUT_5 0.01fF
C46643 NOR2X1_LOC_84/Y NAND2X1_LOC_205/a_36_24# 0.01fF
C46644 INVX1_LOC_299/A NAND2X1_LOC_272/a_36_24# 0.00fF
C46645 INVX1_LOC_223/Y INVX1_LOC_77/A 0.03fF
C46646 INVX1_LOC_269/A NOR2X1_LOC_354/B 0.01fF
C46647 INVX1_LOC_45/A NOR2X1_LOC_103/Y 0.09fF
C46648 NAND2X1_LOC_508/A NOR2X1_LOC_861/Y 0.07fF
C46649 NAND2X1_LOC_304/a_36_24# NOR2X1_LOC_727/B 0.00fF
C46650 INVX1_LOC_88/Y NOR2X1_LOC_665/Y 0.01fF
C46651 NAND2X1_LOC_348/A NOR2X1_LOC_664/a_36_216# 0.00fF
C46652 INVX1_LOC_45/A NOR2X1_LOC_541/Y 0.04fF
C46653 NOR2X1_LOC_447/B INVX1_LOC_118/A 0.02fF
C46654 NAND2X1_LOC_294/a_36_24# INVX1_LOC_23/A 0.00fF
C46655 INVX1_LOC_16/A NAND2X1_LOC_99/A 0.08fF
C46656 NOR2X1_LOC_68/A NAND2X1_LOC_538/Y 0.07fF
C46657 INVX1_LOC_36/A INVX1_LOC_161/Y 0.22fF
C46658 NOR2X1_LOC_541/Y NOR2X1_LOC_568/A 0.04fF
C46659 INVX1_LOC_27/A INVX1_LOC_283/Y -0.01fF
C46660 NOR2X1_LOC_603/Y INVX1_LOC_92/A 0.01fF
C46661 NOR2X1_LOC_261/A INVX1_LOC_117/A 0.05fF
C46662 NOR2X1_LOC_337/A NAND2X1_LOC_74/B 0.00fF
C46663 INVX1_LOC_125/Y INVX1_LOC_63/A 0.09fF
C46664 INVX1_LOC_96/A NOR2X1_LOC_631/A 0.49fF
C46665 INVX1_LOC_75/A INVX1_LOC_290/Y 0.03fF
C46666 NOR2X1_LOC_208/Y NOR2X1_LOC_122/A 0.02fF
C46667 INVX1_LOC_74/Y NAND2X1_LOC_574/A 0.03fF
C46668 NOR2X1_LOC_74/A INVX1_LOC_42/A 0.17fF
C46669 NOR2X1_LOC_186/Y INVX1_LOC_104/A 0.10fF
C46670 INVX1_LOC_89/A NOR2X1_LOC_825/a_36_216# 0.01fF
C46671 INVX1_LOC_110/Y INVX1_LOC_110/A 0.38fF
C46672 INVX1_LOC_12/A INVX1_LOC_309/A 0.03fF
C46673 INVX1_LOC_64/A INVX1_LOC_144/Y 0.03fF
C46674 NOR2X1_LOC_388/a_36_216# INVX1_LOC_53/A 0.01fF
C46675 INVX1_LOC_24/A NOR2X1_LOC_513/Y 0.01fF
C46676 INVX1_LOC_58/A NAND2X1_LOC_564/B 0.46fF
C46677 NOR2X1_LOC_795/Y NOR2X1_LOC_798/A 0.02fF
C46678 NOR2X1_LOC_103/Y INVX1_LOC_71/A 0.10fF
C46679 INVX1_LOC_255/Y D_INPUT_1 0.15fF
C46680 NOR2X1_LOC_711/a_36_216# INVX1_LOC_213/A 0.01fF
C46681 NOR2X1_LOC_9/Y INVX1_LOC_42/A 0.07fF
C46682 INVX1_LOC_36/A NOR2X1_LOC_599/A 0.03fF
C46683 NOR2X1_LOC_160/B INVX1_LOC_181/Y 0.03fF
C46684 NOR2X1_LOC_356/A INVX1_LOC_78/A 0.07fF
C46685 INVX1_LOC_45/A NOR2X1_LOC_568/A 0.07fF
C46686 NOR2X1_LOC_541/Y INVX1_LOC_71/A 0.13fF
C46687 NAND2X1_LOC_218/B INPUT_2 0.05fF
C46688 INVX1_LOC_35/A INVX1_LOC_53/Y 0.10fF
C46689 NOR2X1_LOC_813/Y NAND2X1_LOC_243/B 0.02fF
C46690 INVX1_LOC_12/A INVX1_LOC_91/A 0.14fF
C46691 NOR2X1_LOC_45/B NOR2X1_LOC_671/Y 0.01fF
C46692 NAND2X1_LOC_218/B NAND2X1_LOC_612/a_36_24# 0.00fF
C46693 NAND2X1_LOC_149/Y NOR2X1_LOC_423/Y 0.12fF
C46694 NOR2X1_LOC_86/A NAND2X1_LOC_827/a_36_24# -0.00fF
C46695 INVX1_LOC_90/A NOR2X1_LOC_668/Y 0.01fF
C46696 INVX1_LOC_230/Y NOR2X1_LOC_617/Y 0.02fF
C46697 NOR2X1_LOC_91/A INVX1_LOC_90/A 0.34fF
C46698 NOR2X1_LOC_328/Y NAND2X1_LOC_725/A 0.53fF
C46699 NOR2X1_LOC_15/Y INVX1_LOC_240/A 0.21fF
C46700 INVX1_LOC_108/Y NOR2X1_LOC_195/a_36_216# 0.01fF
C46701 NOR2X1_LOC_759/A INVX1_LOC_30/A 0.72fF
C46702 NAND2X1_LOC_68/a_36_24# INVX1_LOC_96/Y 0.00fF
C46703 NOR2X1_LOC_77/a_36_216# NAND2X1_LOC_642/Y 0.00fF
C46704 NAND2X1_LOC_860/Y INVX1_LOC_306/Y 0.01fF
C46705 INVX1_LOC_21/A NAND2X1_LOC_181/Y 0.03fF
C46706 INVX1_LOC_34/A NOR2X1_LOC_82/A 0.19fF
C46707 INVX1_LOC_2/A INVX1_LOC_52/Y 0.01fF
C46708 NAND2X1_LOC_785/A NAND2X1_LOC_579/A 0.71fF
C46709 D_INPUT_1 NOR2X1_LOC_71/Y 0.23fF
C46710 INVX1_LOC_286/A INVX1_LOC_15/A 0.03fF
C46711 INVX1_LOC_11/Y INVX1_LOC_12/A 0.03fF
C46712 INVX1_LOC_178/Y INVX1_LOC_203/A 0.05fF
C46713 INVX1_LOC_62/A NOR2X1_LOC_416/A 0.02fF
C46714 INVX1_LOC_28/A NAND2X1_LOC_99/A 0.02fF
C46715 NOR2X1_LOC_246/a_36_216# INVX1_LOC_57/A 0.00fF
C46716 NOR2X1_LOC_205/Y NOR2X1_LOC_52/B 0.00fF
C46717 INVX1_LOC_97/A INVX1_LOC_23/A 0.13fF
C46718 NOR2X1_LOC_74/A INVX1_LOC_78/A 0.18fF
C46719 INVX1_LOC_45/A INVX1_LOC_71/A 0.22fF
C46720 NAND2X1_LOC_149/Y NOR2X1_LOC_222/Y 0.19fF
C46721 INVX1_LOC_278/A NOR2X1_LOC_373/Y 0.04fF
C46722 NAND2X1_LOC_186/a_36_24# INVX1_LOC_271/A 0.00fF
C46723 INPUT_0 INVX1_LOC_87/A 0.04fF
C46724 NOR2X1_LOC_272/Y INVX1_LOC_208/Y 0.01fF
C46725 NOR2X1_LOC_568/A INVX1_LOC_71/A 0.15fF
C46726 INVX1_LOC_90/A INVX1_LOC_23/A 0.17fF
C46727 INVX1_LOC_136/A NOR2X1_LOC_13/Y 0.10fF
C46728 INVX1_LOC_103/A INVX1_LOC_96/Y 0.10fF
C46729 INVX1_LOC_245/Y NOR2X1_LOC_377/Y 0.01fF
C46730 INVX1_LOC_12/A NOR2X1_LOC_421/Y 0.08fF
C46731 NOR2X1_LOC_561/Y NOR2X1_LOC_304/Y 0.03fF
C46732 NOR2X1_LOC_88/Y INVX1_LOC_54/A 0.22fF
C46733 D_INPUT_1 NOR2X1_LOC_644/A 0.02fF
C46734 NOR2X1_LOC_9/Y INVX1_LOC_78/A 1.06fF
C46735 INVX1_LOC_21/A NAND2X1_LOC_514/a_36_24# 0.00fF
C46736 NAND2X1_LOC_787/A NAND2X1_LOC_551/A 0.01fF
C46737 INVX1_LOC_223/A NOR2X1_LOC_577/Y 0.00fF
C46738 INVX1_LOC_13/Y NOR2X1_LOC_391/A 0.07fF
C46739 NOR2X1_LOC_201/A NAND2X1_LOC_348/A 0.06fF
C46740 INVX1_LOC_34/A NAND2X1_LOC_500/Y 0.01fF
C46741 INVX1_LOC_135/A NOR2X1_LOC_663/A 0.02fF
C46742 NOR2X1_LOC_392/B INVX1_LOC_31/A 0.07fF
C46743 INVX1_LOC_126/Y INVX1_LOC_26/A 0.01fF
C46744 NAND2X1_LOC_214/Y NOR2X1_LOC_516/B 0.02fF
C46745 NOR2X1_LOC_276/a_36_216# NOR2X1_LOC_208/Y 0.00fF
C46746 INVX1_LOC_5/A D_INPUT_0 1.49fF
C46747 NOR2X1_LOC_65/B NOR2X1_LOC_74/A 0.08fF
C46748 INVX1_LOC_64/A NOR2X1_LOC_473/B 0.19fF
C46749 INVX1_LOC_24/A NOR2X1_LOC_303/Y 0.04fF
C46750 INVX1_LOC_212/Y INVX1_LOC_122/Y 0.03fF
C46751 INVX1_LOC_84/A INVX1_LOC_54/A 0.66fF
C46752 NOR2X1_LOC_607/Y INVX1_LOC_45/Y 0.29fF
C46753 INVX1_LOC_93/A NOR2X1_LOC_130/A 0.07fF
C46754 NAND2X1_LOC_861/Y INVX1_LOC_306/Y 0.32fF
C46755 NOR2X1_LOC_65/B NOR2X1_LOC_9/Y 0.10fF
C46756 NAND2X1_LOC_579/A NOR2X1_LOC_86/A 0.12fF
C46757 INVX1_LOC_123/A INVX1_LOC_16/Y 0.05fF
C46758 NOR2X1_LOC_246/A NOR2X1_LOC_791/Y 0.01fF
C46759 NOR2X1_LOC_274/B INVX1_LOC_149/Y 0.14fF
C46760 VDD INVX1_LOC_170/Y 0.39fF
C46761 NOR2X1_LOC_632/Y NOR2X1_LOC_666/Y 0.00fF
C46762 NOR2X1_LOC_813/Y INVX1_LOC_284/A 1.53fF
C46763 INVX1_LOC_12/Y NOR2X1_LOC_114/Y 0.16fF
C46764 NOR2X1_LOC_598/B NOR2X1_LOC_196/Y 0.01fF
C46765 NOR2X1_LOC_565/a_36_216# INVX1_LOC_53/A 0.01fF
C46766 NOR2X1_LOC_147/a_36_216# INVX1_LOC_117/A 0.01fF
C46767 INVX1_LOC_24/A NOR2X1_LOC_254/Y 0.02fF
C46768 INVX1_LOC_269/A NOR2X1_LOC_298/Y 0.05fF
C46769 NAND2X1_LOC_794/B NOR2X1_LOC_166/Y 0.04fF
C46770 INVX1_LOC_280/A INVX1_LOC_284/A 0.25fF
C46771 D_INPUT_3 NOR2X1_LOC_38/B 0.09fF
C46772 NOR2X1_LOC_361/a_36_216# NOR2X1_LOC_366/B 0.01fF
C46773 INVX1_LOC_124/Y NOR2X1_LOC_773/Y 0.48fF
C46774 VDD NOR2X1_LOC_839/B 0.12fF
C46775 INVX1_LOC_35/A NOR2X1_LOC_113/B 0.08fF
C46776 NAND2X1_LOC_357/B NAND2X1_LOC_731/Y 0.01fF
C46777 NOR2X1_LOC_435/A INVX1_LOC_19/A 0.03fF
C46778 NOR2X1_LOC_592/A INVX1_LOC_10/A -0.01fF
C46779 NAND2X1_LOC_123/a_36_24# INVX1_LOC_23/A 0.00fF
C46780 INVX1_LOC_49/A INVX1_LOC_63/Y 0.15fF
C46781 NAND2X1_LOC_288/A INVX1_LOC_63/A 0.14fF
C46782 INVX1_LOC_136/A INVX1_LOC_256/Y 0.07fF
C46783 NAND2X1_LOC_783/A NOR2X1_LOC_513/Y 0.00fF
C46784 NOR2X1_LOC_640/Y NAND2X1_LOC_74/B 0.11fF
C46785 INVX1_LOC_278/A INVX1_LOC_286/A 0.20fF
C46786 NAND2X1_LOC_577/A INVX1_LOC_16/A 0.00fF
C46787 NAND2X1_LOC_733/Y NAND2X1_LOC_712/A 0.03fF
C46788 NAND2X1_LOC_367/A NAND2X1_LOC_365/a_36_24# 0.02fF
C46789 NOR2X1_LOC_661/a_36_216# INVX1_LOC_285/A 0.00fF
C46790 INVX1_LOC_24/A NOR2X1_LOC_353/Y 0.04fF
C46791 INVX1_LOC_223/A INVX1_LOC_22/A 0.03fF
C46792 INVX1_LOC_194/A NOR2X1_LOC_474/A 0.62fF
C46793 INVX1_LOC_200/A INVX1_LOC_183/Y 0.00fF
C46794 NOR2X1_LOC_653/Y INVX1_LOC_63/A 0.01fF
C46795 INVX1_LOC_21/A NAND2X1_LOC_138/a_36_24# 0.00fF
C46796 NAND2X1_LOC_325/a_36_24# NOR2X1_LOC_406/A 0.00fF
C46797 NOR2X1_LOC_474/A NOR2X1_LOC_399/A 0.01fF
C46798 INVX1_LOC_233/A NOR2X1_LOC_45/B 0.07fF
C46799 NOR2X1_LOC_454/Y INVX1_LOC_75/A 0.10fF
C46800 INVX1_LOC_208/Y NAND2X1_LOC_364/A 0.56fF
C46801 NOR2X1_LOC_488/Y NOR2X1_LOC_91/Y 0.01fF
C46802 NOR2X1_LOC_38/B INVX1_LOC_230/A 0.68fF
C46803 INVX1_LOC_72/A NAND2X1_LOC_479/Y 0.03fF
C46804 INVX1_LOC_54/A INVX1_LOC_15/A 0.21fF
C46805 INVX1_LOC_76/A INVX1_LOC_275/Y 0.03fF
C46806 INVX1_LOC_76/A NOR2X1_LOC_748/A 0.01fF
C46807 NOR2X1_LOC_292/Y NOR2X1_LOC_440/B 0.12fF
C46808 INVX1_LOC_225/A INVX1_LOC_104/A 0.10fF
C46809 INVX1_LOC_19/A INVX1_LOC_63/A 0.21fF
C46810 INVX1_LOC_54/Y NOR2X1_LOC_557/Y 0.16fF
C46811 NOR2X1_LOC_88/Y NOR2X1_LOC_48/B 0.19fF
C46812 INVX1_LOC_2/A INVX1_LOC_63/Y 0.05fF
C46813 VDD INVX1_LOC_271/A 0.15fF
C46814 INVX1_LOC_90/A INVX1_LOC_31/A 3.24fF
C46815 NOR2X1_LOC_440/Y NOR2X1_LOC_360/Y 0.15fF
C46816 INVX1_LOC_45/A NOR2X1_LOC_123/B 0.07fF
C46817 NOR2X1_LOC_536/A INVX1_LOC_26/A 0.37fF
C46818 NOR2X1_LOC_246/A INVX1_LOC_30/A 0.10fF
C46819 VDD INVX1_LOC_105/Y 0.02fF
C46820 INVX1_LOC_256/A NOR2X1_LOC_567/B 0.04fF
C46821 INVX1_LOC_255/Y D_INPUT_2 0.04fF
C46822 NOR2X1_LOC_226/A INVX1_LOC_63/Y 0.12fF
C46823 NOR2X1_LOC_315/Y NOR2X1_LOC_84/Y 0.19fF
C46824 NAND2X1_LOC_236/a_36_24# NAND2X1_LOC_99/A 0.01fF
C46825 NOR2X1_LOC_67/A NAND2X1_LOC_569/A 0.01fF
C46826 INVX1_LOC_17/Y INVX1_LOC_37/Y 0.09fF
C46827 NOR2X1_LOC_78/B NAND2X1_LOC_115/a_36_24# 0.01fF
C46828 NOR2X1_LOC_310/Y INVX1_LOC_149/A 0.06fF
C46829 INVX1_LOC_200/Y INVX1_LOC_37/Y 0.05fF
C46830 NAND2X1_LOC_551/A INVX1_LOC_30/A 0.05fF
C46831 INVX1_LOC_159/A NAND2X1_LOC_156/B 0.01fF
C46832 NAND2X1_LOC_349/B INVX1_LOC_77/A 0.03fF
C46833 NOR2X1_LOC_220/B INVX1_LOC_93/Y 0.12fF
C46834 NOR2X1_LOC_456/Y INVX1_LOC_37/A 0.07fF
C46835 NOR2X1_LOC_668/Y INVX1_LOC_38/A 0.03fF
C46836 INVX1_LOC_232/Y NOR2X1_LOC_514/Y 0.01fF
C46837 INVX1_LOC_17/A NOR2X1_LOC_188/A 0.25fF
C46838 INVX1_LOC_58/A NAND2X1_LOC_804/Y 0.02fF
C46839 NOR2X1_LOC_91/A INVX1_LOC_38/A 3.41fF
C46840 INVX1_LOC_84/A NOR2X1_LOC_48/B 0.43fF
C46841 NOR2X1_LOC_82/A INPUT_0 0.50fF
C46842 INVX1_LOC_226/Y NAND2X1_LOC_276/Y 0.07fF
C46843 INVX1_LOC_202/A NOR2X1_LOC_757/A 0.03fF
C46844 INVX1_LOC_256/Y NOR2X1_LOC_278/A 0.10fF
C46845 INVX1_LOC_17/A NOR2X1_LOC_548/B 0.03fF
C46846 NAND2X1_LOC_214/Y INVX1_LOC_315/Y 0.02fF
C46847 INVX1_LOC_53/A NOR2X1_LOC_139/a_36_216# 0.01fF
C46848 NOR2X1_LOC_186/Y NAND2X1_LOC_674/a_36_24# 0.00fF
C46849 NOR2X1_LOC_218/Y INVX1_LOC_63/Y 0.04fF
C46850 INVX1_LOC_55/A NOR2X1_LOC_74/Y 0.00fF
C46851 D_GATE_741 INVX1_LOC_193/Y 0.56fF
C46852 INVX1_LOC_18/A D_GATE_366 0.07fF
C46853 NOR2X1_LOC_806/Y NOR2X1_LOC_78/B 0.07fF
C46854 NOR2X1_LOC_778/B INVX1_LOC_177/A 0.03fF
C46855 NAND2X1_LOC_348/A INVX1_LOC_31/A 0.11fF
C46856 NOR2X1_LOC_466/a_36_216# INVX1_LOC_91/A 0.00fF
C46857 NOR2X1_LOC_304/Y INVX1_LOC_76/A 0.11fF
C46858 INVX1_LOC_22/A INVX1_LOC_149/Y 0.03fF
C46859 INVX1_LOC_299/A INVX1_LOC_160/A 0.02fF
C46860 INVX1_LOC_45/A INVX1_LOC_102/Y 2.53fF
C46861 INVX1_LOC_24/Y NOR2X1_LOC_78/A 2.91fF
C46862 INVX1_LOC_26/A NAND2X1_LOC_93/B 0.03fF
C46863 INVX1_LOC_38/A INVX1_LOC_23/A 0.13fF
C46864 NAND2X1_LOC_563/Y NOR2X1_LOC_516/B 0.08fF
C46865 NAND2X1_LOC_254/Y NAND2X1_LOC_81/B 0.00fF
C46866 NAND2X1_LOC_214/B VDD 0.14fF
C46867 INVX1_LOC_124/A INVX1_LOC_25/Y 0.25fF
C46868 NOR2X1_LOC_48/B NAND2X1_LOC_651/B 0.04fF
C46869 NAND2X1_LOC_787/A NOR2X1_LOC_692/Y 0.21fF
C46870 NOR2X1_LOC_389/B INVX1_LOC_111/A 0.00fF
C46871 NOR2X1_LOC_423/Y INVX1_LOC_16/A 0.06fF
C46872 NOR2X1_LOC_458/B NOR2X1_LOC_78/B 0.01fF
C46873 D_INPUT_1 NAND2X1_LOC_698/a_36_24# 0.01fF
C46874 INVX1_LOC_5/A NOR2X1_LOC_859/Y 0.07fF
C46875 INVX1_LOC_41/A NAND2X1_LOC_474/a_36_24# 0.00fF
C46876 INVX1_LOC_256/A NOR2X1_LOC_269/Y 0.10fF
C46877 INVX1_LOC_27/A VDD 2.86fF
C46878 NOR2X1_LOC_355/A INVX1_LOC_155/Y 0.02fF
C46879 INVX1_LOC_11/A NOR2X1_LOC_595/Y 0.08fF
C46880 NOR2X1_LOC_744/Y NOR2X1_LOC_329/B 0.03fF
C46881 INVX1_LOC_14/A INVX1_LOC_95/Y 0.36fF
C46882 NOR2X1_LOC_669/a_36_216# INVX1_LOC_20/A 0.02fF
C46883 NOR2X1_LOC_613/Y INVX1_LOC_46/A 0.01fF
C46884 INVX1_LOC_119/A NOR2X1_LOC_561/Y 0.02fF
C46885 NOR2X1_LOC_92/Y NAND2X1_LOC_464/A 0.01fF
C46886 NAND2X1_LOC_733/B NAND2X1_LOC_863/B 0.04fF
C46887 INVX1_LOC_178/A NOR2X1_LOC_682/Y 0.12fF
C46888 NOR2X1_LOC_84/A NOR2X1_LOC_130/A 0.02fF
C46889 INVX1_LOC_5/A NAND2X1_LOC_848/A 0.00fF
C46890 INVX1_LOC_47/Y INVX1_LOC_29/A 0.02fF
C46891 INVX1_LOC_278/A INVX1_LOC_54/A 0.07fF
C46892 NOR2X1_LOC_222/Y INVX1_LOC_16/A 3.53fF
C46893 INVX1_LOC_237/A VDD -0.00fF
C46894 INVX1_LOC_71/A INVX1_LOC_102/Y 0.10fF
C46895 D_INPUT_0 NAND2X1_LOC_562/B 0.03fF
C46896 INVX1_LOC_21/A INVX1_LOC_117/A 0.16fF
C46897 NAND2X1_LOC_736/Y NAND2X1_LOC_379/a_36_24# 0.01fF
C46898 INVX1_LOC_26/A INVX1_LOC_3/A 0.03fF
C46899 NAND2X1_LOC_727/Y NOR2X1_LOC_773/Y 0.02fF
C46900 NOR2X1_LOC_667/A NAND2X1_LOC_390/A 0.06fF
C46901 INVX1_LOC_11/A INVX1_LOC_115/Y 0.02fF
C46902 NOR2X1_LOC_388/Y INVX1_LOC_313/Y 0.01fF
C46903 NOR2X1_LOC_312/Y NAND2X1_LOC_357/B 0.12fF
C46904 INVX1_LOC_217/A INVX1_LOC_309/A 0.17fF
C46905 NAND2X1_LOC_9/Y NOR2X1_LOC_862/B 0.03fF
C46906 INVX1_LOC_2/A NOR2X1_LOC_370/a_36_216# 0.01fF
C46907 INVX1_LOC_26/Y INVX1_LOC_63/A 0.18fF
C46908 INVX1_LOC_69/Y NOR2X1_LOC_360/Y 0.10fF
C46909 NAND2X1_LOC_190/Y INVX1_LOC_14/Y 0.10fF
C46910 NOR2X1_LOC_718/B INVX1_LOC_85/Y 0.18fF
C46911 INVX1_LOC_77/A INVX1_LOC_75/A 1.06fF
C46912 NOR2X1_LOC_48/B INVX1_LOC_15/A 0.07fF
C46913 INVX1_LOC_179/A NOR2X1_LOC_678/A 0.40fF
C46914 INVX1_LOC_89/A NAND2X1_LOC_629/Y 0.00fF
C46915 NOR2X1_LOC_200/a_36_216# NOR2X1_LOC_214/B 0.00fF
C46916 NOR2X1_LOC_92/Y NOR2X1_LOC_60/Y 0.01fF
C46917 NAND2X1_LOC_733/Y INVX1_LOC_11/Y 2.98fF
C46918 INVX1_LOC_135/A NOR2X1_LOC_537/Y 0.03fF
C46919 NOR2X1_LOC_553/B NOR2X1_LOC_500/Y 0.02fF
C46920 NAND2X1_LOC_662/Y INVX1_LOC_22/A 0.07fF
C46921 INVX1_LOC_292/A NOR2X1_LOC_137/a_36_216# 0.00fF
C46922 INVX1_LOC_135/A NAND2X1_LOC_338/B 0.10fF
C46923 NAND2X1_LOC_525/a_36_24# INVX1_LOC_275/A 0.00fF
C46924 NAND2X1_LOC_717/Y NOR2X1_LOC_380/A 0.01fF
C46925 NOR2X1_LOC_160/B INVX1_LOC_115/A 0.46fF
C46926 INVX1_LOC_84/A NAND2X1_LOC_215/A 0.13fF
C46927 INVX1_LOC_295/A INVX1_LOC_192/Y 0.03fF
C46928 INVX1_LOC_217/A INVX1_LOC_91/A 0.07fF
C46929 INVX1_LOC_152/Y NOR2X1_LOC_865/Y 0.03fF
C46930 INVX1_LOC_113/Y NOR2X1_LOC_74/A 0.03fF
C46931 NOR2X1_LOC_496/Y INVX1_LOC_118/A 0.01fF
C46932 NAND2X1_LOC_550/A NAND2X1_LOC_254/a_36_24# 0.00fF
C46933 D_INPUT_0 NAND2X1_LOC_9/a_36_24# 0.00fF
C46934 D_INPUT_0 NOR2X1_LOC_773/Y 0.07fF
C46935 INVX1_LOC_135/A NAND2X1_LOC_323/B 0.00fF
C46936 NOR2X1_LOC_255/Y INVX1_LOC_3/A 0.17fF
C46937 NOR2X1_LOC_321/Y INVX1_LOC_118/Y 0.07fF
C46938 INVX1_LOC_152/Y NOR2X1_LOC_243/B 0.02fF
C46939 INVX1_LOC_5/A INVX1_LOC_46/Y 0.07fF
C46940 NOR2X1_LOC_781/A NOR2X1_LOC_589/A 0.09fF
C46941 INVX1_LOC_99/Y NOR2X1_LOC_197/B 0.03fF
C46942 NAND2X1_LOC_352/B NAND2X1_LOC_287/B 0.07fF
C46943 INVX1_LOC_75/A NOR2X1_LOC_732/A 0.01fF
C46944 NAND2X1_LOC_338/B NOR2X1_LOC_560/A -0.09fF
C46945 NAND2X1_LOC_3/B INVX1_LOC_15/A 0.20fF
C46946 NOR2X1_LOC_841/A NOR2X1_LOC_109/Y 0.13fF
C46947 NAND2X1_LOC_123/Y INVX1_LOC_177/A 0.03fF
C46948 INVX1_LOC_217/A INVX1_LOC_11/Y 0.07fF
C46949 NAND2X1_LOC_787/B INVX1_LOC_309/A 0.00fF
C46950 NOR2X1_LOC_798/A NOR2X1_LOC_862/B 0.05fF
C46951 NAND2X1_LOC_85/Y NOR2X1_LOC_845/a_36_216# 0.00fF
C46952 NOR2X1_LOC_375/Y INVX1_LOC_89/A 0.02fF
C46953 NOR2X1_LOC_742/A INVX1_LOC_266/Y 0.06fF
C46954 NAND2X1_LOC_144/a_36_24# INVX1_LOC_275/A 0.00fF
C46955 INVX1_LOC_124/A INVX1_LOC_75/A 0.10fF
C46956 INVX1_LOC_30/A NOR2X1_LOC_357/Y 0.00fF
C46957 INVX1_LOC_89/A NOR2X1_LOC_719/A 0.01fF
C46958 NOR2X1_LOC_816/A NAND2X1_LOC_848/A 0.24fF
C46959 NOR2X1_LOC_666/A NAND2X1_LOC_93/B 0.03fF
C46960 INVX1_LOC_5/A INVX1_LOC_5/Y 0.03fF
C46961 NOR2X1_LOC_392/B INVX1_LOC_6/A 0.01fF
C46962 NOR2X1_LOC_464/Y INVX1_LOC_4/A 0.03fF
C46963 NOR2X1_LOC_100/A INPUT_0 0.04fF
C46964 INVX1_LOC_41/A INVX1_LOC_98/A 0.03fF
C46965 INVX1_LOC_94/A NAND2X1_LOC_447/Y 0.10fF
C46966 NOR2X1_LOC_52/Y INVX1_LOC_46/A 0.03fF
C46967 NOR2X1_LOC_596/A NAND2X1_LOC_212/Y 0.02fF
C46968 INVX1_LOC_120/A NOR2X1_LOC_97/B 0.15fF
C46969 INVX1_LOC_141/A NOR2X1_LOC_536/A 0.01fF
C46970 NOR2X1_LOC_438/Y INVX1_LOC_15/A 0.03fF
C46971 INVX1_LOC_90/A NAND2X1_LOC_859/Y 0.12fF
C46972 NOR2X1_LOC_91/Y NAND2X1_LOC_650/B 0.19fF
C46973 INVX1_LOC_31/A NAND2X1_LOC_849/B 0.10fF
C46974 INVX1_LOC_41/A NOR2X1_LOC_78/A 0.19fF
C46975 D_INPUT_0 NOR2X1_LOC_332/A 0.09fF
C46976 INVX1_LOC_89/A INVX1_LOC_7/A 1.82fF
C46977 NOR2X1_LOC_655/B NOR2X1_LOC_335/B 0.03fF
C46978 INVX1_LOC_31/A INVX1_LOC_38/A 0.28fF
C46979 INVX1_LOC_171/Y NAND2X1_LOC_475/Y 0.01fF
C46980 INVX1_LOC_11/Y NAND2X1_LOC_787/B 0.15fF
C46981 NAND2X1_LOC_200/B NOR2X1_LOC_721/Y 0.02fF
C46982 NOR2X1_LOC_631/B NOR2X1_LOC_550/B 0.10fF
C46983 INVX1_LOC_296/A NOR2X1_LOC_467/A 1.13fF
C46984 NOR2X1_LOC_569/Y NOR2X1_LOC_569/a_36_216# 0.00fF
C46985 INVX1_LOC_278/Y INPUT_0 0.72fF
C46986 NOR2X1_LOC_596/A INVX1_LOC_14/Y 0.03fF
C46987 INVX1_LOC_314/Y NAND2X1_LOC_267/B 0.02fF
C46988 INVX1_LOC_304/Y INVX1_LOC_91/A 0.07fF
C46989 INVX1_LOC_45/A NOR2X1_LOC_331/B 0.07fF
C46990 INVX1_LOC_77/A NOR2X1_LOC_309/a_36_216# 0.00fF
C46991 INVX1_LOC_249/A NOR2X1_LOC_69/a_36_216# 0.00fF
C46992 INVX1_LOC_249/A VDD 0.41fF
C46993 NOR2X1_LOC_52/B NOR2X1_LOC_595/Y 0.01fF
C46994 NAND2X1_LOC_493/Y NOR2X1_LOC_485/Y 0.00fF
C46995 INVX1_LOC_233/Y NAND2X1_LOC_254/Y 0.01fF
C46996 NOR2X1_LOC_392/Y NOR2X1_LOC_861/Y 0.24fF
C46997 NOR2X1_LOC_810/A NOR2X1_LOC_567/B 0.13fF
C46998 INVX1_LOC_278/A NOR2X1_LOC_48/B -0.01fF
C46999 INVX1_LOC_104/A NAND2X1_LOC_642/Y 0.00fF
C47000 INVX1_LOC_34/A INVX1_LOC_59/Y 0.10fF
C47001 INVX1_LOC_34/A INVX1_LOC_112/A 0.01fF
C47002 INVX1_LOC_6/Y VDD 0.21fF
C47003 NAND2X1_LOC_833/Y INVX1_LOC_20/A 0.00fF
C47004 NOR2X1_LOC_596/Y NOR2X1_LOC_155/A 0.01fF
C47005 NAND2X1_LOC_350/A NOR2X1_LOC_88/Y 0.05fF
C47006 NOR2X1_LOC_550/B INVX1_LOC_37/A 0.43fF
C47007 D_INPUT_0 INVX1_LOC_140/A 0.07fF
C47008 NAND2X1_LOC_363/B INVX1_LOC_32/A 0.07fF
C47009 NOR2X1_LOC_677/Y INVX1_LOC_273/A 0.03fF
C47010 INVX1_LOC_30/A NOR2X1_LOC_451/A 0.05fF
C47011 NOR2X1_LOC_247/a_36_216# INVX1_LOC_36/Y 0.00fF
C47012 INVX1_LOC_90/A NAND2X1_LOC_807/Y 0.43fF
C47013 NOR2X1_LOC_773/Y NOR2X1_LOC_191/a_36_216# 0.01fF
C47014 NOR2X1_LOC_350/A NAND2X1_LOC_96/A 0.03fF
C47015 NOR2X1_LOC_454/a_36_216# INVX1_LOC_77/Y 0.00fF
C47016 NOR2X1_LOC_778/B INVX1_LOC_65/A 0.01fF
C47017 NOR2X1_LOC_664/Y VDD 0.88fF
C47018 INVX1_LOC_119/A INVX1_LOC_76/A 0.02fF
C47019 INVX1_LOC_71/A NOR2X1_LOC_331/B 0.26fF
C47020 NAND2X1_LOC_477/A NAND2X1_LOC_464/A 0.27fF
C47021 INPUT_0 INVX1_LOC_306/A 0.00fF
C47022 INVX1_LOC_45/A NOR2X1_LOC_592/B 0.03fF
C47023 NAND2X1_LOC_570/Y NAND2X1_LOC_659/B 0.02fF
C47024 D_GATE_222 INVX1_LOC_91/A 0.01fF
C47025 INVX1_LOC_161/Y INVX1_LOC_63/A 0.07fF
C47026 NAND2X1_LOC_357/B NAND2X1_LOC_287/B 0.15fF
C47027 NOR2X1_LOC_329/B INVX1_LOC_28/A 0.11fF
C47028 NAND2X1_LOC_181/Y INVX1_LOC_304/A 0.02fF
C47029 INVX1_LOC_266/Y INVX1_LOC_139/A 0.02fF
C47030 NOR2X1_LOC_392/Y NOR2X1_LOC_825/a_36_216# 0.00fF
C47031 NOR2X1_LOC_844/Y NOR2X1_LOC_243/B 0.04fF
C47032 NOR2X1_LOC_759/Y INVX1_LOC_157/Y 0.00fF
C47033 INVX1_LOC_208/Y NOR2X1_LOC_405/A 0.08fF
C47034 NOR2X1_LOC_791/Y INVX1_LOC_32/A 0.03fF
C47035 NOR2X1_LOC_82/A NOR2X1_LOC_84/B 0.00fF
C47036 INVX1_LOC_206/A VDD 0.57fF
C47037 INVX1_LOC_21/A INVX1_LOC_3/Y 0.07fF
C47038 NOR2X1_LOC_78/B NOR2X1_LOC_603/Y 0.01fF
C47039 NAND2X1_LOC_149/Y NOR2X1_LOC_477/B 0.04fF
C47040 INVX1_LOC_164/Y INVX1_LOC_20/A 0.07fF
C47041 NOR2X1_LOC_401/B INVX1_LOC_76/A 0.06fF
C47042 INVX1_LOC_56/Y NOR2X1_LOC_124/A 0.02fF
C47043 INVX1_LOC_16/A INPUT_4 0.01fF
C47044 NAND2X1_LOC_570/Y VDD 0.03fF
C47045 D_INPUT_1 NOR2X1_LOC_39/Y 0.04fF
C47046 NOR2X1_LOC_410/Y NOR2X1_LOC_461/B 0.12fF
C47047 NOR2X1_LOC_112/B NOR2X1_LOC_112/Y 0.11fF
C47048 NOR2X1_LOC_759/A INVX1_LOC_113/A 0.03fF
C47049 INVX1_LOC_314/A INVX1_LOC_22/A 0.04fF
C47050 INVX1_LOC_278/A NOR2X1_LOC_438/Y 0.01fF
C47051 NOR2X1_LOC_160/B NOR2X1_LOC_509/A 0.01fF
C47052 INVX1_LOC_90/A INVX1_LOC_6/A 0.13fF
C47053 INVX1_LOC_312/A INVX1_LOC_63/A -0.00fF
C47054 NOR2X1_LOC_191/B NOR2X1_LOC_216/B 0.02fF
C47055 NOR2X1_LOC_773/Y NOR2X1_LOC_266/B 0.01fF
C47056 INVX1_LOC_24/A INVX1_LOC_35/Y 0.58fF
C47057 INVX1_LOC_63/Y INVX1_LOC_118/A 0.00fF
C47058 NAND2X1_LOC_808/A INVX1_LOC_91/A 0.08fF
C47059 NAND2X1_LOC_200/B VDD 0.16fF
C47060 INVX1_LOC_30/A NAND2X1_LOC_489/Y 0.06fF
C47061 NOR2X1_LOC_389/B INVX1_LOC_6/A 0.01fF
C47062 NOR2X1_LOC_844/A INVX1_LOC_230/A 0.05fF
C47063 INVX1_LOC_176/Y INVX1_LOC_9/A 0.01fF
C47064 NOR2X1_LOC_820/A NOR2X1_LOC_649/B 0.03fF
C47065 NOR2X1_LOC_251/Y VDD 0.13fF
C47066 NOR2X1_LOC_500/A NAND2X1_LOC_237/a_36_24# 0.01fF
C47067 NAND2X1_LOC_722/A NOR2X1_LOC_692/Y 0.01fF
C47068 NOR2X1_LOC_418/a_36_216# INVX1_LOC_77/Y 0.01fF
C47069 NOR2X1_LOC_695/Y VDD 0.34fF
C47070 INVX1_LOC_103/Y NAND2X1_LOC_93/B 0.04fF
C47071 INVX1_LOC_69/Y NOR2X1_LOC_567/B 0.00fF
C47072 NOR2X1_LOC_160/B NOR2X1_LOC_114/Y 0.03fF
C47073 INVX1_LOC_191/Y INVX1_LOC_38/A 0.01fF
C47074 NOR2X1_LOC_537/Y INVX1_LOC_280/A 0.07fF
C47075 INVX1_LOC_11/A D_INPUT_5 0.09fF
C47076 NOR2X1_LOC_457/A INVX1_LOC_32/A 0.07fF
C47077 NOR2X1_LOC_773/Y NAND2X1_LOC_848/A 0.10fF
C47078 NOR2X1_LOC_561/Y NOR2X1_LOC_52/a_36_216# 0.01fF
C47079 INVX1_LOC_273/Y INVX1_LOC_20/A 0.01fF
C47080 NOR2X1_LOC_254/Y NOR2X1_LOC_197/B 0.04fF
C47081 INVX1_LOC_103/Y NAND2X1_LOC_425/Y 0.03fF
C47082 INVX1_LOC_24/A NOR2X1_LOC_721/B 0.06fF
C47083 INVX1_LOC_146/A NOR2X1_LOC_45/B 0.01fF
C47084 NOR2X1_LOC_198/a_36_216# INVX1_LOC_78/Y 0.00fF
C47085 NAND2X1_LOC_350/A INVX1_LOC_15/A 0.08fF
C47086 INVX1_LOC_234/A VDD 0.61fF
C47087 NAND2X1_LOC_156/B VDD 0.10fF
C47088 NAND2X1_LOC_811/Y NAND2X1_LOC_770/Y 0.01fF
C47089 NOR2X1_LOC_76/A INVX1_LOC_20/A 0.03fF
C47090 NOR2X1_LOC_510/Y INVX1_LOC_271/A 0.04fF
C47091 INVX1_LOC_89/A INVX1_LOC_76/A 0.18fF
C47092 INVX1_LOC_190/A NAND2X1_LOC_453/A 0.05fF
C47093 NAND2X1_LOC_177/a_36_24# INVX1_LOC_179/A 0.01fF
C47094 INVX1_LOC_218/Y INVX1_LOC_15/A 0.01fF
C47095 NOR2X1_LOC_441/Y INVX1_LOC_15/A 0.03fF
C47096 NAND2X1_LOC_859/Y NAND2X1_LOC_849/B 0.10fF
C47097 INVX1_LOC_18/A INVX1_LOC_102/A 0.07fF
C47098 NOR2X1_LOC_360/Y NOR2X1_LOC_89/A 0.05fF
C47099 NAND2X1_LOC_539/a_36_24# INVX1_LOC_94/Y 0.00fF
C47100 INVX1_LOC_58/A INVX1_LOC_21/A 0.07fF
C47101 INVX1_LOC_315/A NOR2X1_LOC_649/B 0.15fF
C47102 NOR2X1_LOC_142/Y INVX1_LOC_84/A 0.47fF
C47103 NAND2X1_LOC_139/A NOR2X1_LOC_23/a_36_216# 0.03fF
C47104 NOR2X1_LOC_790/B INVX1_LOC_50/Y 0.07fF
C47105 NAND2X1_LOC_349/B INVX1_LOC_9/A 0.20fF
C47106 NOR2X1_LOC_19/B NAND2X1_LOC_659/B 0.01fF
C47107 NOR2X1_LOC_302/B INVX1_LOC_9/A 0.01fF
C47108 INVX1_LOC_245/Y INVX1_LOC_78/A 0.01fF
C47109 INVX1_LOC_30/A INVX1_LOC_32/A 0.93fF
C47110 NOR2X1_LOC_598/B NOR2X1_LOC_846/A 0.02fF
C47111 NAND2X1_LOC_656/Y NOR2X1_LOC_366/a_36_216# 0.01fF
C47112 INVX1_LOC_30/A NOR2X1_LOC_623/B 0.20fF
C47113 INVX1_LOC_143/A NAND2X1_LOC_412/a_36_24# 0.00fF
C47114 INVX1_LOC_256/A INVX1_LOC_26/A 0.02fF
C47115 NAND2X1_LOC_711/B INVX1_LOC_102/A 0.07fF
C47116 NAND2X1_LOC_807/A NOR2X1_LOC_301/A 0.01fF
C47117 NOR2X1_LOC_624/a_36_216# INVX1_LOC_26/Y 0.00fF
C47118 NOR2X1_LOC_582/Y NAND2X1_LOC_95/a_36_24# 0.00fF
C47119 NOR2X1_LOC_772/A VDD 0.12fF
C47120 NOR2X1_LOC_71/a_36_216# NOR2X1_LOC_78/A 0.00fF
C47121 INVX1_LOC_31/A NAND2X1_LOC_223/A 0.07fF
C47122 INVX1_LOC_77/A NAND2X1_LOC_291/B 0.16fF
C47123 NOR2X1_LOC_770/A NOR2X1_LOC_89/A 0.01fF
C47124 NOR2X1_LOC_250/Y NOR2X1_LOC_65/B 0.68fF
C47125 NOR2X1_LOC_793/Y INVX1_LOC_57/A 0.21fF
C47126 INVX1_LOC_73/A INVX1_LOC_20/A 0.09fF
C47127 INVX1_LOC_2/A INVX1_LOC_27/Y 0.01fF
C47128 INVX1_LOC_35/A INVX1_LOC_235/Y 0.04fF
C47129 NOR2X1_LOC_19/B VDD 0.98fF
C47130 NOR2X1_LOC_361/B INVX1_LOC_271/A 0.00fF
C47131 INVX1_LOC_161/Y NOR2X1_LOC_65/Y 0.02fF
C47132 NAND2X1_LOC_549/a_36_24# INVX1_LOC_29/A 0.00fF
C47133 INVX1_LOC_35/A NAND2X1_LOC_149/Y 0.08fF
C47134 INVX1_LOC_172/A INVX1_LOC_102/A 0.07fF
C47135 NAND2X1_LOC_585/a_36_24# INVX1_LOC_12/A 0.00fF
C47136 INPUT_0 INVX1_LOC_59/Y 0.03fF
C47137 NOR2X1_LOC_168/B NOR2X1_LOC_814/A 0.03fF
C47138 NOR2X1_LOC_717/Y INVX1_LOC_271/Y 0.03fF
C47139 INVX1_LOC_85/A INVX1_LOC_186/Y 0.14fF
C47140 INVX1_LOC_96/Y NOR2X1_LOC_631/A 0.31fF
C47141 INVX1_LOC_313/A INVX1_LOC_38/A 0.01fF
C47142 NOR2X1_LOC_655/B INVX1_LOC_84/A 0.01fF
C47143 NAND2X1_LOC_565/B INVX1_LOC_35/Y 0.00fF
C47144 INVX1_LOC_226/Y NOR2X1_LOC_103/a_36_216# 0.00fF
C47145 NOR2X1_LOC_457/B INVX1_LOC_4/A 0.02fF
C47146 NOR2X1_LOC_391/A NOR2X1_LOC_99/Y 3.30fF
C47147 NAND2X1_LOC_866/B INVX1_LOC_38/A 0.07fF
C47148 INVX1_LOC_30/A NAND2X1_LOC_175/Y 0.10fF
C47149 NOR2X1_LOC_553/B INVX1_LOC_307/A 0.02fF
C47150 INPUT_0 INVX1_LOC_176/A 0.03fF
C47151 NOR2X1_LOC_817/Y D_INPUT_1 0.11fF
C47152 INVX1_LOC_21/A NAND2X1_LOC_190/a_36_24# 0.01fF
C47153 NOR2X1_LOC_799/a_36_216# NAND2X1_LOC_74/B 0.02fF
C47154 NOR2X1_LOC_68/A NOR2X1_LOC_334/Y 0.10fF
C47155 NOR2X1_LOC_67/A NOR2X1_LOC_662/A 0.07fF
C47156 NOR2X1_LOC_688/Y INVX1_LOC_26/Y 0.01fF
C47157 INVX1_LOC_25/A INVX1_LOC_293/A 0.05fF
C47158 NOR2X1_LOC_637/Y NOR2X1_LOC_329/a_36_216# 0.00fF
C47159 NOR2X1_LOC_792/B NOR2X1_LOC_89/A 0.29fF
C47160 NAND2X1_LOC_807/Y INVX1_LOC_38/A 0.07fF
C47161 INVX1_LOC_291/Y INVX1_LOC_264/Y 0.02fF
C47162 NOR2X1_LOC_121/Y INVX1_LOC_42/A 0.15fF
C47163 INVX1_LOC_140/A NAND2X1_LOC_848/A 0.10fF
C47164 NOR2X1_LOC_483/B INVX1_LOC_23/A 0.03fF
C47165 NAND2X1_LOC_51/B INVX1_LOC_117/A 0.02fF
C47166 NOR2X1_LOC_366/Y NOR2X1_LOC_155/A 0.04fF
C47167 NOR2X1_LOC_186/Y NOR2X1_LOC_92/Y 0.07fF
C47168 INVX1_LOC_314/Y INVX1_LOC_4/Y 0.10fF
C47169 INVX1_LOC_30/A INVX1_LOC_262/A 0.06fF
C47170 NOR2X1_LOC_348/B INVX1_LOC_290/Y 0.51fF
C47171 NOR2X1_LOC_91/A NAND2X1_LOC_501/a_36_24# 0.01fF
C47172 NOR2X1_LOC_340/Y INVX1_LOC_15/A 0.03fF
C47173 NOR2X1_LOC_334/A INVX1_LOC_37/A 0.25fF
C47174 NOR2X1_LOC_130/A INVX1_LOC_35/Y 0.09fF
C47175 INVX1_LOC_269/A INVX1_LOC_13/Y 0.10fF
C47176 NOR2X1_LOC_389/B NOR2X1_LOC_79/A 0.03fF
C47177 NOR2X1_LOC_142/Y INVX1_LOC_15/A 0.12fF
C47178 NOR2X1_LOC_15/Y NOR2X1_LOC_233/a_36_216# 0.00fF
C47179 NAND2X1_LOC_21/Y NAND2X1_LOC_3/B 0.65fF
C47180 NOR2X1_LOC_778/B NOR2X1_LOC_830/Y 0.01fF
C47181 INVX1_LOC_45/A NOR2X1_LOC_493/A 0.18fF
C47182 INVX1_LOC_75/A INVX1_LOC_9/A 0.29fF
C47183 NOR2X1_LOC_92/Y NAND2X1_LOC_573/Y 0.07fF
C47184 NOR2X1_LOC_528/Y VDD 1.21fF
C47185 NAND2X1_LOC_468/B NOR2X1_LOC_275/A 0.01fF
C47186 INVX1_LOC_1/Y INVX1_LOC_19/A 0.28fF
C47187 NAND2X1_LOC_656/Y NOR2X1_LOC_814/A 0.01fF
C47188 NOR2X1_LOC_526/Y NAND2X1_LOC_254/Y 0.05fF
C47189 INVX1_LOC_59/A INVX1_LOC_14/A 0.05fF
C47190 NOR2X1_LOC_99/B INVX1_LOC_84/A 0.07fF
C47191 NOR2X1_LOC_314/a_36_216# NOR2X1_LOC_56/Y 0.00fF
C47192 INVX1_LOC_6/A INVX1_LOC_38/A 0.03fF
C47193 NOR2X1_LOC_349/A NAND2X1_LOC_224/a_36_24# 0.01fF
C47194 INVX1_LOC_299/A INVX1_LOC_1/A 0.03fF
C47195 NAND2X1_LOC_773/Y INVX1_LOC_14/A 0.01fF
C47196 NOR2X1_LOC_703/B INVX1_LOC_53/A 0.03fF
C47197 NOR2X1_LOC_392/B NOR2X1_LOC_80/Y 0.15fF
C47198 INVX1_LOC_303/A NOR2X1_LOC_621/A 0.04fF
C47199 INVX1_LOC_62/A INVX1_LOC_63/A 0.07fF
C47200 INVX1_LOC_132/Y NOR2X1_LOC_814/A 0.13fF
C47201 INVX1_LOC_221/A INVX1_LOC_94/Y 0.03fF
C47202 INVX1_LOC_17/A NAND2X1_LOC_326/A 0.45fF
C47203 NOR2X1_LOC_15/Y NOR2X1_LOC_533/Y 0.03fF
C47204 NOR2X1_LOC_538/B INVX1_LOC_1/A 0.02fF
C47205 INVX1_LOC_22/A INVX1_LOC_290/Y 0.03fF
C47206 INVX1_LOC_225/A NOR2X1_LOC_281/a_36_216# 0.00fF
C47207 NAND2X1_LOC_555/Y NAND2X1_LOC_141/a_36_24# 0.01fF
C47208 INVX1_LOC_256/A NOR2X1_LOC_666/A 0.09fF
C47209 NAND2X1_LOC_803/B NAND2X1_LOC_780/Y 0.19fF
C47210 INVX1_LOC_93/A INVX1_LOC_286/Y -0.09fF
C47211 NAND2X1_LOC_860/A INVX1_LOC_24/A 0.06fF
C47212 NOR2X1_LOC_690/Y INVX1_LOC_102/A 0.09fF
C47213 NAND2X1_LOC_784/A NAND2X1_LOC_547/a_36_24# 0.00fF
C47214 INVX1_LOC_219/A INVX1_LOC_29/A 0.02fF
C47215 NAND2X1_LOC_192/a_36_24# NOR2X1_LOC_205/Y 0.00fF
C47216 NAND2X1_LOC_725/B NAND2X1_LOC_550/A 0.02fF
C47217 NOR2X1_LOC_778/B INVX1_LOC_4/Y 0.68fF
C47218 NOR2X1_LOC_772/Y INVX1_LOC_270/A 0.05fF
C47219 INVX1_LOC_252/Y INVX1_LOC_14/A 0.04fF
C47220 NAND2X1_LOC_722/A NAND2X1_LOC_175/Y 0.04fF
C47221 INVX1_LOC_30/A INVX1_LOC_171/Y 0.08fF
C47222 NAND2X1_LOC_325/Y INVX1_LOC_57/A 4.05fF
C47223 NOR2X1_LOC_590/A NAND2X1_LOC_780/Y 0.01fF
C47224 INVX1_LOC_268/Y NOR2X1_LOC_467/A 0.21fF
C47225 NAND2X1_LOC_642/Y NOR2X1_LOC_119/a_36_216# 0.01fF
C47226 INVX1_LOC_33/A INVX1_LOC_23/A 0.28fF
C47227 NAND2X1_LOC_342/a_36_24# NOR2X1_LOC_652/Y 0.00fF
C47228 NAND2X1_LOC_573/A INVX1_LOC_170/Y 0.09fF
C47229 NOR2X1_LOC_510/a_36_216# INVX1_LOC_12/A 0.00fF
C47230 INVX1_LOC_48/Y NAND2X1_LOC_577/A 0.01fF
C47231 NOR2X1_LOC_84/Y NAND2X1_LOC_99/A 0.19fF
C47232 INVX1_LOC_242/Y GATE_579 0.32fF
C47233 D_INPUT_0 INVX1_LOC_42/A 7.04fF
C47234 NOR2X1_LOC_537/Y NOR2X1_LOC_541/B 0.02fF
C47235 NOR2X1_LOC_823/Y INVX1_LOC_118/A 0.05fF
C47236 NOR2X1_LOC_92/Y INVX1_LOC_170/A 0.40fF
C47237 INPUT_1 NAND2X1_LOC_83/a_36_24# 0.00fF
C47238 INVX1_LOC_91/A INVX1_LOC_92/A 0.33fF
C47239 INVX1_LOC_186/A NOR2X1_LOC_155/A 0.03fF
C47240 NOR2X1_LOC_570/Y NOR2X1_LOC_334/Y 0.02fF
C47241 INVX1_LOC_35/A NOR2X1_LOC_623/a_36_216# 0.02fF
C47242 INVX1_LOC_25/A NOR2X1_LOC_315/Y 2.81fF
C47243 INVX1_LOC_269/A NOR2X1_LOC_500/B 0.01fF
C47244 INVX1_LOC_5/A INVX1_LOC_49/A 0.23fF
C47245 INVX1_LOC_196/A NOR2X1_LOC_383/B 0.03fF
C47246 INVX1_LOC_265/A INVX1_LOC_233/A 0.03fF
C47247 NOR2X1_LOC_99/B INVX1_LOC_15/A 0.08fF
C47248 NOR2X1_LOC_598/B NAND2X1_LOC_116/A 0.02fF
C47249 INVX1_LOC_276/A INVX1_LOC_57/A 0.05fF
C47250 NAND2X1_LOC_660/Y INVX1_LOC_78/A 0.02fF
C47251 NAND2X1_LOC_803/B INVX1_LOC_141/Y 0.01fF
C47252 NOR2X1_LOC_590/A NAND2X1_LOC_114/B 0.01fF
C47253 NOR2X1_LOC_521/a_36_216# INVX1_LOC_23/A 0.00fF
C47254 NOR2X1_LOC_67/A INVX1_LOC_57/A 0.14fF
C47255 NOR2X1_LOC_545/B NOR2X1_LOC_862/B 0.03fF
C47256 NAND2X1_LOC_774/a_36_24# INVX1_LOC_18/A 0.00fF
C47257 INVX1_LOC_22/Y NAND2X1_LOC_114/B 0.06fF
C47258 NOR2X1_LOC_846/B INVX1_LOC_15/A 0.02fF
C47259 NAND2X1_LOC_803/B INVX1_LOC_312/Y 0.03fF
C47260 INVX1_LOC_1/Y INVX1_LOC_26/Y 0.65fF
C47261 INVX1_LOC_212/Y INVX1_LOC_50/Y 0.01fF
C47262 INVX1_LOC_58/A NOR2X1_LOC_667/A 0.10fF
C47263 NAND2X1_LOC_840/B NOR2X1_LOC_677/Y 0.03fF
C47264 NOR2X1_LOC_45/B INVX1_LOC_119/Y 0.09fF
C47265 NOR2X1_LOC_590/A INVX1_LOC_141/Y 0.06fF
C47266 INVX1_LOC_224/A NOR2X1_LOC_360/Y 0.03fF
C47267 INVX1_LOC_17/A NAND2X1_LOC_481/a_36_24# 0.00fF
C47268 INPUT_0 NOR2X1_LOC_340/A 0.11fF
C47269 NAND2X1_LOC_860/A INVX1_LOC_143/A 0.01fF
C47270 NAND2X1_LOC_773/Y NAND2X1_LOC_84/Y 0.01fF
C47271 NOR2X1_LOC_440/Y INVX1_LOC_26/A 0.03fF
C47272 INVX1_LOC_24/A NAND2X1_LOC_537/Y 0.02fF
C47273 D_INPUT_0 INVX1_LOC_78/A 0.14fF
C47274 NOR2X1_LOC_284/B NOR2X1_LOC_598/B 0.03fF
C47275 NOR2X1_LOC_82/A INVX1_LOC_72/Y 0.07fF
C47276 NOR2X1_LOC_254/A INVX1_LOC_142/A 0.05fF
C47277 INVX1_LOC_233/A NOR2X1_LOC_401/Y 0.01fF
C47278 INVX1_LOC_27/A INVX1_LOC_153/Y 0.10fF
C47279 NOR2X1_LOC_65/B NAND2X1_LOC_660/Y 0.01fF
C47280 NOR2X1_LOC_590/A INVX1_LOC_312/Y 0.45fF
C47281 INVX1_LOC_165/Y INVX1_LOC_23/A 0.02fF
C47282 INVX1_LOC_256/A NOR2X1_LOC_276/B 0.01fF
C47283 INVX1_LOC_291/Y INVX1_LOC_84/A 0.03fF
C47284 INVX1_LOC_93/A INVX1_LOC_185/Y 0.01fF
C47285 NOR2X1_LOC_639/B NAND2X1_LOC_11/Y 0.01fF
C47286 INVX1_LOC_90/A NOR2X1_LOC_80/Y 0.10fF
C47287 INVX1_LOC_2/A NAND2X1_LOC_552/A 0.03fF
C47288 INVX1_LOC_132/A INVX1_LOC_24/Y 0.10fF
C47289 INVX1_LOC_201/Y NAND2X1_LOC_574/a_36_24# 0.03fF
C47290 NAND2X1_LOC_68/a_36_24# INVX1_LOC_34/A 0.00fF
C47291 NOR2X1_LOC_186/Y NAND2X1_LOC_477/A 0.10fF
C47292 VDD NOR2X1_LOC_216/B 1.97fF
C47293 INVX1_LOC_2/A INVX1_LOC_5/A 0.08fF
C47294 INVX1_LOC_5/A NOR2X1_LOC_818/Y 0.11fF
C47295 INVX1_LOC_27/A INVX1_LOC_121/Y 0.14fF
C47296 NAND2X1_LOC_565/B NAND2X1_LOC_860/A 0.00fF
C47297 INVX1_LOC_266/A NOR2X1_LOC_344/A 0.01fF
C47298 INVX1_LOC_64/A NAND2X1_LOC_372/a_36_24# 0.00fF
C47299 NOR2X1_LOC_226/A NAND2X1_LOC_552/A 0.05fF
C47300 INVX1_LOC_73/A INVX1_LOC_4/A 0.10fF
C47301 NOR2X1_LOC_130/A NAND2X1_LOC_286/B 0.03fF
C47302 NOR2X1_LOC_400/B INVX1_LOC_135/A 0.05fF
C47303 NOR2X1_LOC_65/B D_INPUT_0 1.68fF
C47304 NAND2X1_LOC_787/A NAND2X1_LOC_564/B 0.00fF
C47305 INVX1_LOC_225/A NOR2X1_LOC_92/Y 0.03fF
C47306 INVX1_LOC_35/A INVX1_LOC_16/A 0.10fF
C47307 NOR2X1_LOC_719/A NOR2X1_LOC_392/Y 0.20fF
C47308 NAND2X1_LOC_149/Y INVX1_LOC_257/Y -0.02fF
C47309 NOR2X1_LOC_709/A NAND2X1_LOC_474/Y 0.45fF
C47310 INVX1_LOC_248/Y INVX1_LOC_248/A 0.01fF
C47311 NOR2X1_LOC_536/A NOR2X1_LOC_235/Y 0.01fF
C47312 NAND2X1_LOC_573/Y NAND2X1_LOC_477/A 0.10fF
C47313 INVX1_LOC_2/A INVX1_LOC_178/A 0.01fF
C47314 NAND2X1_LOC_337/B INVX1_LOC_49/A 0.88fF
C47315 NOR2X1_LOC_45/B INVX1_LOC_284/A 0.14fF
C47316 INVX1_LOC_186/A NOR2X1_LOC_833/B 0.34fF
C47317 NOR2X1_LOC_366/Y NOR2X1_LOC_125/Y 0.00fF
C47318 INVX1_LOC_34/A INVX1_LOC_103/A 0.15fF
C47319 NOR2X1_LOC_691/A NOR2X1_LOC_857/A 0.03fF
C47320 NOR2X1_LOC_389/A NOR2X1_LOC_106/Y 0.03fF
C47321 INVX1_LOC_223/Y INVX1_LOC_179/Y 0.02fF
C47322 INVX1_LOC_245/Y INVX1_LOC_113/Y 0.45fF
C47323 NOR2X1_LOC_751/Y INVX1_LOC_305/A 0.08fF
C47324 INVX1_LOC_1/A NOR2X1_LOC_315/Y 0.10fF
C47325 INVX1_LOC_59/Y NOR2X1_LOC_84/B 0.00fF
C47326 VDD NAND2X1_LOC_477/Y 0.41fF
C47327 INVX1_LOC_64/A NOR2X1_LOC_781/A 0.03fF
C47328 NOR2X1_LOC_218/Y INVX1_LOC_5/A 0.02fF
C47329 NOR2X1_LOC_226/A INVX1_LOC_178/A 2.81fF
C47330 NOR2X1_LOC_82/A NOR2X1_LOC_514/a_36_216# 0.00fF
C47331 NOR2X1_LOC_824/A INVX1_LOC_280/Y 0.07fF
C47332 INVX1_LOC_7/A NOR2X1_LOC_392/Y 0.00fF
C47333 INVX1_LOC_90/A INVX1_LOC_270/A 0.06fF
C47334 NOR2X1_LOC_331/B NOR2X1_LOC_592/B 0.05fF
C47335 NAND2X1_LOC_860/A NOR2X1_LOC_130/A 0.07fF
C47336 INVX1_LOC_11/A NOR2X1_LOC_792/B 0.02fF
C47337 NOR2X1_LOC_389/B INVX1_LOC_270/A 0.01fF
C47338 INVX1_LOC_135/A NAND2X1_LOC_793/B 0.10fF
C47339 NOR2X1_LOC_68/A NOR2X1_LOC_523/B 0.05fF
C47340 INVX1_LOC_280/Y INVX1_LOC_237/A 0.04fF
C47341 NOR2X1_LOC_432/Y INVX1_LOC_1/A 0.01fF
C47342 INVX1_LOC_17/A NOR2X1_LOC_87/B 3.67fF
C47343 NOR2X1_LOC_61/Y NOR2X1_LOC_61/A 0.01fF
C47344 INVX1_LOC_34/A INVX1_LOC_292/A 0.03fF
C47345 INVX1_LOC_235/Y INVX1_LOC_84/Y 0.06fF
C47346 INVX1_LOC_90/A NOR2X1_LOC_416/A 0.19fF
C47347 INVX1_LOC_64/A INVX1_LOC_273/Y 0.01fF
C47348 INVX1_LOC_5/A NAND2X1_LOC_664/a_36_24# 0.00fF
C47349 INVX1_LOC_68/Y NAND2X1_LOC_473/A 0.16fF
C47350 INVX1_LOC_108/Y NOR2X1_LOC_846/B 0.01fF
C47351 INVX1_LOC_103/A NAND2X1_LOC_231/Y 0.10fF
C47352 INVX1_LOC_77/A NOR2X1_LOC_274/B 0.06fF
C47353 INVX1_LOC_50/A NOR2X1_LOC_197/Y 0.02fF
C47354 INVX1_LOC_256/A INVX1_LOC_149/A 0.02fF
C47355 INVX1_LOC_37/A NAND2X1_LOC_74/B 0.03fF
C47356 NOR2X1_LOC_454/Y INVX1_LOC_22/A 0.12fF
C47357 INVX1_LOC_161/A INVX1_LOC_240/A 0.05fF
C47358 NOR2X1_LOC_751/a_36_216# INVX1_LOC_1/Y 0.00fF
C47359 INVX1_LOC_255/A INVX1_LOC_3/Y 0.06fF
C47360 INVX1_LOC_11/A NAND2X1_LOC_451/Y 0.09fF
C47361 NOR2X1_LOC_557/A INVX1_LOC_4/Y 0.07fF
C47362 INVX1_LOC_87/Y NOR2X1_LOC_717/A 0.01fF
C47363 NAND2X1_LOC_391/Y NAND2X1_LOC_392/Y 0.20fF
C47364 INVX1_LOC_101/Y INVX1_LOC_208/A 0.00fF
C47365 INVX1_LOC_45/A NOR2X1_LOC_388/Y 0.02fF
C47366 INVX1_LOC_2/A NAND2X1_LOC_337/B 0.00fF
C47367 INVX1_LOC_2/A NOR2X1_LOC_816/A 0.06fF
C47368 INVX1_LOC_64/A NOR2X1_LOC_180/B 0.08fF
C47369 NOR2X1_LOC_361/B NOR2X1_LOC_251/Y 0.13fF
C47370 NOR2X1_LOC_598/B NOR2X1_LOC_775/Y 0.03fF
C47371 INVX1_LOC_125/Y INVX1_LOC_87/A 0.34fF
C47372 NAND2X1_LOC_555/Y NOR2X1_LOC_87/B 0.09fF
C47373 INVX1_LOC_90/A NOR2X1_LOC_109/Y 0.07fF
C47374 NOR2X1_LOC_443/Y NOR2X1_LOC_97/A 0.03fF
C47375 NOR2X1_LOC_435/A NOR2X1_LOC_841/A 0.03fF
C47376 INVX1_LOC_35/A INVX1_LOC_28/A 0.15fF
C47377 NOR2X1_LOC_670/Y INVX1_LOC_3/Y 0.12fF
C47378 INVX1_LOC_67/A INVX1_LOC_79/Y 0.01fF
C47379 NAND2X1_LOC_552/A INPUT_1 0.05fF
C47380 NOR2X1_LOC_226/A NOR2X1_LOC_816/A 0.10fF
C47381 INVX1_LOC_36/A NOR2X1_LOC_392/B 2.46fF
C47382 NAND2X1_LOC_348/A NOR2X1_LOC_416/A 0.19fF
C47383 INVX1_LOC_58/A NAND2X1_LOC_51/B 0.01fF
C47384 NOR2X1_LOC_590/A NOR2X1_LOC_168/B 0.09fF
C47385 INVX1_LOC_5/A INPUT_1 0.15fF
C47386 NOR2X1_LOC_307/a_36_216# INVX1_LOC_117/A 0.00fF
C47387 NOR2X1_LOC_593/Y NOR2X1_LOC_360/Y 0.01fF
C47388 INVX1_LOC_45/Y NOR2X1_LOC_335/A 0.00fF
C47389 NOR2X1_LOC_544/A NOR2X1_LOC_160/B 0.01fF
C47390 INVX1_LOC_79/A INVX1_LOC_53/A 0.08fF
C47391 INVX1_LOC_18/A INVX1_LOC_149/Y 0.00fF
C47392 INVX1_LOC_77/A NOR2X1_LOC_160/a_36_216# 0.00fF
C47393 INVX1_LOC_58/A INVX1_LOC_311/A 0.33fF
C47394 NAND2X1_LOC_577/A INVX1_LOC_216/A 0.07fF
C47395 INVX1_LOC_289/A INVX1_LOC_211/A 0.00fF
C47396 INVX1_LOC_64/A INVX1_LOC_73/A 0.01fF
C47397 INVX1_LOC_77/A NOR2X1_LOC_577/Y 0.45fF
C47398 INVX1_LOC_85/A INVX1_LOC_18/A 0.00fF
C47399 NOR2X1_LOC_379/Y INVX1_LOC_77/A 0.05fF
C47400 INVX1_LOC_269/A INVX1_LOC_80/A 0.04fF
C47401 NAND2X1_LOC_182/A NOR2X1_LOC_91/Y 0.00fF
C47402 NAND2X1_LOC_783/A NAND2X1_LOC_537/Y 0.29fF
C47403 NOR2X1_LOC_361/B INVX1_LOC_234/A 0.30fF
C47404 INVX1_LOC_123/A NAND2X1_LOC_215/A 1.27fF
C47405 NAND2X1_LOC_848/A INVX1_LOC_42/A 0.07fF
C47406 INVX1_LOC_31/A INVX1_LOC_40/A 0.44fF
C47407 NAND2X1_LOC_387/B INVX1_LOC_192/Y 0.03fF
C47408 INVX1_LOC_249/A INVX1_LOC_153/Y 0.03fF
C47409 D_INPUT_1 INVX1_LOC_286/A 0.07fF
C47410 INVX1_LOC_163/A INVX1_LOC_89/A 0.19fF
C47411 NAND2X1_LOC_291/B INVX1_LOC_9/A 0.04fF
C47412 INVX1_LOC_53/A NOR2X1_LOC_728/B 0.05fF
C47413 NOR2X1_LOC_194/Y NOR2X1_LOC_596/A 0.00fF
C47414 INVX1_LOC_132/A INVX1_LOC_41/A 0.10fF
C47415 INVX1_LOC_19/A INVX1_LOC_117/Y 0.03fF
C47416 NOR2X1_LOC_841/A INVX1_LOC_63/A 0.36fF
C47417 INVX1_LOC_256/A INVX1_LOC_164/A 0.23fF
C47418 NAND2X1_LOC_374/Y INVX1_LOC_217/A 0.10fF
C47419 NOR2X1_LOC_78/B NOR2X1_LOC_703/B 0.06fF
C47420 NOR2X1_LOC_743/Y NAND2X1_LOC_74/B 0.03fF
C47421 INVX1_LOC_78/A NOR2X1_LOC_266/B 0.15fF
C47422 INVX1_LOC_314/A NOR2X1_LOC_843/B 0.02fF
C47423 NAND2X1_LOC_833/Y NAND2X1_LOC_833/a_36_24# 0.00fF
C47424 INVX1_LOC_2/A NOR2X1_LOC_759/a_36_216# 0.00fF
C47425 NOR2X1_LOC_49/a_36_216# NAND2X1_LOC_773/B 0.01fF
C47426 NOR2X1_LOC_598/B INVX1_LOC_186/A 0.14fF
C47427 NOR2X1_LOC_682/Y INVX1_LOC_78/A 0.01fF
C47428 INVX1_LOC_95/Y NOR2X1_LOC_383/B 0.13fF
C47429 INVX1_LOC_53/A INVX1_LOC_91/A 0.30fF
C47430 NAND2X1_LOC_564/B INVX1_LOC_30/A 0.35fF
C47431 NOR2X1_LOC_68/A INVX1_LOC_218/A 0.03fF
C47432 NAND2X1_LOC_472/Y NAND2X1_LOC_454/Y 0.13fF
C47433 NOR2X1_LOC_89/A NOR2X1_LOC_79/Y 0.24fF
C47434 NOR2X1_LOC_590/A NAND2X1_LOC_656/Y 0.02fF
C47435 NOR2X1_LOC_772/Y NOR2X1_LOC_309/Y 0.21fF
C47436 INVX1_LOC_30/A GATE_662 0.04fF
C47437 NAND2X1_LOC_287/B NOR2X1_LOC_282/Y 0.03fF
C47438 NOR2X1_LOC_486/Y INVX1_LOC_23/A 0.01fF
C47439 INVX1_LOC_34/A INVX1_LOC_240/A 0.02fF
C47440 INVX1_LOC_50/A NOR2X1_LOC_556/a_36_216# 0.02fF
C47441 INVX1_LOC_99/Y NOR2X1_LOC_337/Y 0.06fF
C47442 NOR2X1_LOC_536/A NAND2X1_LOC_471/Y 0.14fF
C47443 INVX1_LOC_46/Y INVX1_LOC_42/A 0.14fF
C47444 INVX1_LOC_136/A NOR2X1_LOC_605/a_36_216# 0.00fF
C47445 NAND2X1_LOC_763/B GATE_662 0.06fF
C47446 INVX1_LOC_36/A NOR2X1_LOC_512/a_36_216# 0.00fF
C47447 INVX1_LOC_286/A NOR2X1_LOC_652/Y -0.01fF
C47448 NOR2X1_LOC_273/Y NOR2X1_LOC_219/Y 0.07fF
C47449 INVX1_LOC_18/A NAND2X1_LOC_662/Y 0.57fF
C47450 NOR2X1_LOC_309/Y NOR2X1_LOC_392/B 0.01fF
C47451 INVX1_LOC_27/A INVX1_LOC_285/Y 0.01fF
C47452 NAND2X1_LOC_848/A INVX1_LOC_78/A 0.02fF
C47453 INVX1_LOC_58/A NOR2X1_LOC_670/Y 0.09fF
C47454 INVX1_LOC_29/A INVX1_LOC_220/A 0.12fF
C47455 NOR2X1_LOC_219/Y NOR2X1_LOC_759/Y 0.10fF
C47456 INVX1_LOC_229/A NAND2X1_LOC_463/B 0.21fF
C47457 INVX1_LOC_225/A NAND2X1_LOC_477/A 0.03fF
C47458 INVX1_LOC_45/A INVX1_LOC_135/A 1.40fF
C47459 INVX1_LOC_41/A NOR2X1_LOC_209/Y 0.03fF
C47460 NAND2X1_LOC_30/Y INVX1_LOC_140/A 0.95fF
C47461 NOR2X1_LOC_773/Y INVX1_LOC_49/A 0.07fF
C47462 NOR2X1_LOC_540/B NOR2X1_LOC_678/A 0.01fF
C47463 INVX1_LOC_299/A NOR2X1_LOC_188/A 0.10fF
C47464 INVX1_LOC_246/A NOR2X1_LOC_329/B 0.07fF
C47465 NAND2X1_LOC_20/B INVX1_LOC_75/A 0.04fF
C47466 NOR2X1_LOC_99/a_36_216# INVX1_LOC_16/Y 0.01fF
C47467 INVX1_LOC_14/A NAND2X1_LOC_858/B 0.01fF
C47468 INVX1_LOC_77/A INVX1_LOC_22/A 0.81fF
C47469 NOR2X1_LOC_759/Y NOR2X1_LOC_665/A 0.02fF
C47470 INVX1_LOC_35/A NOR2X1_LOC_35/Y 0.05fF
C47471 INVX1_LOC_50/A NOR2X1_LOC_363/Y 0.01fF
C47472 INVX1_LOC_299/A NOR2X1_LOC_548/B 0.10fF
C47473 NAND2X1_LOC_141/Y NOR2X1_LOC_554/A 0.03fF
C47474 NOR2X1_LOC_392/Y INVX1_LOC_76/A 0.00fF
C47475 INVX1_LOC_103/A INPUT_0 0.01fF
C47476 NOR2X1_LOC_90/a_36_216# INPUT_1 0.00fF
C47477 INVX1_LOC_36/A INVX1_LOC_90/A 0.29fF
C47478 INVX1_LOC_259/Y INVX1_LOC_37/A 0.01fF
C47479 NOR2X1_LOC_413/Y NOR2X1_LOC_399/Y 0.03fF
C47480 NOR2X1_LOC_243/Y INVX1_LOC_64/Y 0.24fF
C47481 INVX1_LOC_17/A NOR2X1_LOC_815/A 0.45fF
C47482 INVX1_LOC_206/A INVX1_LOC_177/A 0.00fF
C47483 INVX1_LOC_95/A NOR2X1_LOC_652/Y 0.01fF
C47484 NAND2X1_LOC_660/Y NOR2X1_LOC_152/Y 0.02fF
C47485 NOR2X1_LOC_471/Y NOR2X1_LOC_74/a_36_216# 0.00fF
C47486 NOR2X1_LOC_763/A NOR2X1_LOC_588/A 0.04fF
C47487 INVX1_LOC_36/A NOR2X1_LOC_389/B 0.07fF
C47488 NAND2X1_LOC_35/Y NAND2X1_LOC_464/A 0.01fF
C47489 NOR2X1_LOC_582/A NOR2X1_LOC_588/A 0.03fF
C47490 INVX1_LOC_27/A INVX1_LOC_65/A 0.00fF
C47491 NOR2X1_LOC_570/B NOR2X1_LOC_553/Y 0.03fF
C47492 NAND2X1_LOC_787/A NAND2X1_LOC_804/Y 0.01fF
C47493 NAND2X1_LOC_358/B INVX1_LOC_37/A 0.00fF
C47494 NAND2X1_LOC_391/Y NOR2X1_LOC_368/Y 0.01fF
C47495 INVX1_LOC_292/A INPUT_0 0.07fF
C47496 NOR2X1_LOC_323/Y INVX1_LOC_31/A 0.08fF
C47497 NOR2X1_LOC_178/a_36_216# NAND2X1_LOC_74/B 0.00fF
C47498 INVX1_LOC_5/A NOR2X1_LOC_586/Y 0.41fF
C47499 INVX1_LOC_99/Y VDD 0.05fF
C47500 NOR2X1_LOC_92/Y NAND2X1_LOC_642/Y 0.03fF
C47501 INVX1_LOC_38/A NOR2X1_LOC_416/A 0.06fF
C47502 INVX1_LOC_2/A NOR2X1_LOC_773/Y 0.07fF
C47503 INVX1_LOC_57/A NOR2X1_LOC_729/A 0.07fF
C47504 INVX1_LOC_295/A INVX1_LOC_71/A 0.08fF
C47505 NOR2X1_LOC_565/A INVX1_LOC_75/A 0.04fF
C47506 NOR2X1_LOC_449/A NOR2X1_LOC_592/B 0.08fF
C47507 INVX1_LOC_226/Y NOR2X1_LOC_709/A 0.13fF
C47508 NOR2X1_LOC_780/B NOR2X1_LOC_708/A 0.23fF
C47509 NOR2X1_LOC_169/B INVX1_LOC_75/A 0.01fF
C47510 INVX1_LOC_36/A NAND2X1_LOC_348/A 0.03fF
C47511 INVX1_LOC_90/A NOR2X1_LOC_208/Y 0.03fF
C47512 NOR2X1_LOC_351/Y INVX1_LOC_23/A 0.04fF
C47513 INVX1_LOC_93/A VDD 0.00fF
C47514 INVX1_LOC_124/A INVX1_LOC_22/A 0.11fF
C47515 NOR2X1_LOC_226/A NOR2X1_LOC_773/Y 0.09fF
C47516 INVX1_LOC_181/Y NAND2X1_LOC_850/A 0.05fF
C47517 D_INPUT_1 INVX1_LOC_54/A 0.07fF
C47518 NOR2X1_LOC_65/B INVX1_LOC_46/Y 0.13fF
C47519 NOR2X1_LOC_111/A NOR2X1_LOC_406/A 0.24fF
C47520 INVX1_LOC_90/A NOR2X1_LOC_237/Y 0.03fF
C47521 NAND2X1_LOC_45/a_36_24# INVX1_LOC_120/A 0.00fF
C47522 INVX1_LOC_13/Y INVX1_LOC_12/Y 0.10fF
C47523 NOR2X1_LOC_590/A INVX1_LOC_78/Y 0.03fF
C47524 INVX1_LOC_73/A INVX1_LOC_130/Y 0.16fF
C47525 INVX1_LOC_33/A INVX1_LOC_313/A 0.42fF
C47526 INVX1_LOC_38/A NOR2X1_LOC_109/Y 0.03fF
C47527 NOR2X1_LOC_128/B NOR2X1_LOC_6/B 0.02fF
C47528 NAND2X1_LOC_513/B VDD 0.01fF
C47529 NOR2X1_LOC_241/a_36_216# INVX1_LOC_117/A 0.00fF
C47530 NOR2X1_LOC_754/A INVX1_LOC_42/A 0.02fF
C47531 NOR2X1_LOC_544/A NOR2X1_LOC_516/B 0.07fF
C47532 NOR2X1_LOC_322/Y INVX1_LOC_41/Y 0.03fF
C47533 NOR2X1_LOC_48/B NOR2X1_LOC_677/a_36_216# 0.01fF
C47534 NOR2X1_LOC_222/Y INVX1_LOC_290/A 0.08fF
C47535 NAND2X1_LOC_112/Y NOR2X1_LOC_136/Y 0.01fF
C47536 NOR2X1_LOC_863/Y NOR2X1_LOC_852/Y 0.03fF
C47537 INVX1_LOC_87/A INVX1_LOC_19/A 0.00fF
C47538 INVX1_LOC_193/Y NOR2X1_LOC_546/A 0.00fF
C47539 NOR2X1_LOC_63/a_36_216# NOR2X1_LOC_99/B 0.01fF
C47540 INVX1_LOC_16/A NOR2X1_LOC_121/A 0.04fF
C47541 INVX1_LOC_90/A NOR2X1_LOC_309/Y 0.04fF
C47542 NOR2X1_LOC_160/B NAND2X1_LOC_468/B 0.03fF
C47543 NOR2X1_LOC_332/A NOR2X1_LOC_818/Y 0.03fF
C47544 INVX1_LOC_280/Y INVX1_LOC_234/A 0.01fF
C47545 NAND2X1_LOC_72/B NAND2X1_LOC_74/B 0.03fF
C47546 D_INPUT_0 NOR2X1_LOC_721/A 0.02fF
C47547 NOR2X1_LOC_389/B NOR2X1_LOC_309/Y 0.03fF
C47548 NAND2X1_LOC_510/A NOR2X1_LOC_349/A 0.29fF
C47549 INVX1_LOC_50/A NOR2X1_LOC_485/Y 0.01fF
C47550 INVX1_LOC_45/A NOR2X1_LOC_552/A 0.07fF
C47551 INVX1_LOC_34/A NOR2X1_LOC_597/a_36_216# 0.02fF
C47552 INVX1_LOC_72/A NOR2X1_LOC_45/B 0.09fF
C47553 NOR2X1_LOC_513/Y VDD 0.12fF
C47554 INVX1_LOC_88/A INVX1_LOC_12/Y 0.03fF
C47555 INVX1_LOC_282/A NAND2X1_LOC_838/a_36_24# 0.00fF
C47556 NOR2X1_LOC_570/Y NOR2X1_LOC_569/Y 0.03fF
C47557 NOR2X1_LOC_552/A NOR2X1_LOC_568/A 0.01fF
C47558 NOR2X1_LOC_561/Y INVX1_LOC_25/Y 0.15fF
C47559 NOR2X1_LOC_298/Y NAND2X1_LOC_853/Y 0.04fF
C47560 INVX1_LOC_249/A INVX1_LOC_285/Y 0.03fF
C47561 INVX1_LOC_178/A INVX1_LOC_118/A 0.05fF
C47562 NAND2X1_LOC_833/Y INVX1_LOC_282/A 0.01fF
C47563 INVX1_LOC_23/Y INVX1_LOC_29/A 0.03fF
C47564 NOR2X1_LOC_89/A INVX1_LOC_26/A 3.89fF
C47565 INVX1_LOC_78/A NOR2X1_LOC_754/A 0.01fF
C47566 D_INPUT_0 NAND2X1_LOC_859/B 0.02fF
C47567 NOR2X1_LOC_717/A NOR2X1_LOC_814/A 0.05fF
C47568 NOR2X1_LOC_773/Y INPUT_1 0.00fF
C47569 INVX1_LOC_106/Y NOR2X1_LOC_668/Y 0.06fF
C47570 INVX1_LOC_33/A INVX1_LOC_6/A 0.38fF
C47571 INVX1_LOC_2/A INVX1_LOC_140/A 0.10fF
C47572 INVX1_LOC_310/Y NOR2X1_LOC_334/A 0.03fF
C47573 INVX1_LOC_240/A INPUT_0 0.02fF
C47574 NOR2X1_LOC_657/a_36_216# NOR2X1_LOC_155/A 0.00fF
C47575 NOR2X1_LOC_552/A INVX1_LOC_71/A 0.10fF
C47576 INVX1_LOC_227/A NAND2X1_LOC_656/Y 0.07fF
C47577 NOR2X1_LOC_226/A INVX1_LOC_140/A 0.11fF
C47578 NOR2X1_LOC_439/B INVX1_LOC_179/Y 0.09fF
C47579 NOR2X1_LOC_433/A NOR2X1_LOC_269/Y 0.10fF
C47580 INVX1_LOC_31/A NOR2X1_LOC_816/Y 0.05fF
C47581 NOR2X1_LOC_584/Y INVX1_LOC_57/A 0.03fF
C47582 NAND2X1_LOC_564/A NOR2X1_LOC_89/A 0.01fF
C47583 NOR2X1_LOC_337/Y NOR2X1_LOC_254/Y 0.02fF
C47584 INVX1_LOC_269/A NOR2X1_LOC_99/Y 0.14fF
C47585 INVX1_LOC_63/Y NOR2X1_LOC_7/Y 0.01fF
C47586 NOR2X1_LOC_855/A NAND2X1_LOC_829/a_36_24# 0.02fF
C47587 NOR2X1_LOC_667/a_36_216# INVX1_LOC_38/A 0.00fF
C47588 INVX1_LOC_75/A INVX1_LOC_179/Y 0.14fF
C47589 NOR2X1_LOC_78/B INVX1_LOC_79/A 0.68fF
C47590 NAND2X1_LOC_337/B INVX1_LOC_118/A 0.07fF
C47591 NOR2X1_LOC_816/A INVX1_LOC_118/A 0.01fF
C47592 INVX1_LOC_206/A INVX1_LOC_285/Y 0.08fF
C47593 NOR2X1_LOC_605/B NAND2X1_LOC_807/Y 0.03fF
C47594 INVX1_LOC_45/A NOR2X1_LOC_813/Y 0.08fF
C47595 NOR2X1_LOC_15/Y NOR2X1_LOC_831/B 0.07fF
C47596 NAND2X1_LOC_579/A NOR2X1_LOC_88/Y 0.03fF
C47597 INVX1_LOC_45/A NOR2X1_LOC_152/A 0.01fF
C47598 NAND2X1_LOC_721/B INVX1_LOC_33/Y 0.02fF
C47599 INVX1_LOC_21/A NAND2X1_LOC_475/Y 0.03fF
C47600 INVX1_LOC_35/A INVX1_LOC_109/A 0.03fF
C47601 INVX1_LOC_13/Y NAND2X1_LOC_465/a_36_24# 0.01fF
C47602 D_INPUT_0 NAND2X1_LOC_861/Y 0.07fF
C47603 NOR2X1_LOC_2/Y NOR2X1_LOC_44/a_36_216# 0.00fF
C47604 INVX1_LOC_41/A NAND2X1_LOC_642/Y 4.13fF
C47605 INVX1_LOC_268/A NOR2X1_LOC_163/Y 0.17fF
C47606 INVX1_LOC_36/A NOR2X1_LOC_561/A 0.01fF
C47607 INVX1_LOC_212/A VDD 0.12fF
C47608 NAND2X1_LOC_793/Y INVX1_LOC_70/A 0.01fF
C47609 NOR2X1_LOC_332/A INPUT_1 0.02fF
C47610 INVX1_LOC_45/A INVX1_LOC_280/A 0.02fF
C47611 NOR2X1_LOC_68/A NAND2X1_LOC_472/Y 0.10fF
C47612 INVX1_LOC_5/A NAND2X1_LOC_63/Y 0.05fF
C47613 INVX1_LOC_89/A NAND2X1_LOC_45/Y 3.09fF
C47614 NOR2X1_LOC_576/B INVX1_LOC_173/Y 0.04fF
C47615 NOR2X1_LOC_763/Y NAND2X1_LOC_638/Y 0.08fF
C47616 NOR2X1_LOC_500/A VDD 0.07fF
C47617 NOR2X1_LOC_52/B NOR2X1_LOC_269/Y 0.07fF
C47618 INVX1_LOC_36/A INVX1_LOC_38/A 1.50fF
C47619 INVX1_LOC_128/A NOR2X1_LOC_65/Y 0.08fF
C47620 NOR2X1_LOC_303/Y VDD 1.18fF
C47621 NOR2X1_LOC_577/Y NAND2X1_LOC_649/a_36_24# 0.00fF
C47622 NOR2X1_LOC_655/B INVX1_LOC_123/A 0.10fF
C47623 INVX1_LOC_63/Y NAND2X1_LOC_212/Y 0.01fF
C47624 NAND2X1_LOC_579/A INVX1_LOC_84/A 0.01fF
C47625 INVX1_LOC_26/Y INVX1_LOC_87/A 0.06fF
C47626 NAND2X1_LOC_832/Y INVX1_LOC_22/A 0.03fF
C47627 INVX1_LOC_40/A INVX1_LOC_6/A 0.11fF
C47628 NAND2X1_LOC_477/A NAND2X1_LOC_642/Y 0.03fF
C47629 INVX1_LOC_25/Y NOR2X1_LOC_167/Y 0.03fF
C47630 NAND2X1_LOC_112/Y INVX1_LOC_144/A 0.03fF
C47631 NOR2X1_LOC_454/Y INVX1_LOC_186/Y 0.08fF
C47632 NOR2X1_LOC_682/Y NOR2X1_LOC_152/Y 0.03fF
C47633 NOR2X1_LOC_561/Y INVX1_LOC_75/A 0.19fF
C47634 NOR2X1_LOC_632/Y NOR2X1_LOC_74/A 0.04fF
C47635 INVX1_LOC_10/A NAND2X1_LOC_863/A 0.13fF
C47636 NOR2X1_LOC_333/A INVX1_LOC_148/A 0.20fF
C47637 NAND2X1_LOC_338/B NOR2X1_LOC_45/B 0.07fF
C47638 INVX1_LOC_7/A INVX1_LOC_75/A 0.01fF
C47639 NOR2X1_LOC_383/B INVX1_LOC_271/Y 0.09fF
C47640 INVX1_LOC_35/A NOR2X1_LOC_460/a_36_216# 0.00fF
C47641 NOR2X1_LOC_78/B INVX1_LOC_91/A 0.27fF
C47642 NAND2X1_LOC_807/B NOR2X1_LOC_652/Y 0.01fF
C47643 NOR2X1_LOC_788/B NOR2X1_LOC_356/A 0.03fF
C47644 INVX1_LOC_36/A NOR2X1_LOC_51/A 0.06fF
C47645 INVX1_LOC_256/Y INVX1_LOC_70/Y 0.22fF
C47646 INVX1_LOC_34/A NOR2X1_LOC_137/Y 0.03fF
C47647 NAND2X1_LOC_465/Y NAND2X1_LOC_464/A 0.12fF
C47648 INVX1_LOC_201/Y D_GATE_662 0.01fF
C47649 NOR2X1_LOC_254/Y VDD 0.18fF
C47650 NOR2X1_LOC_68/A NAND2X1_LOC_637/Y 0.03fF
C47651 NOR2X1_LOC_454/Y INVX1_LOC_261/A 0.04fF
C47652 NOR2X1_LOC_658/Y NOR2X1_LOC_364/A 0.01fF
C47653 NOR2X1_LOC_84/A VDD 0.27fF
C47654 NOR2X1_LOC_208/Y INVX1_LOC_38/A 0.03fF
C47655 NAND2X1_LOC_223/A NOR2X1_LOC_416/A 0.07fF
C47656 INVX1_LOC_166/A INVX1_LOC_175/A 0.22fF
C47657 INVX1_LOC_153/A INVX1_LOC_117/A 0.03fF
C47658 INVX1_LOC_136/A NOR2X1_LOC_743/Y 0.01fF
C47659 INVX1_LOC_140/A INPUT_1 0.07fF
C47660 NOR2X1_LOC_300/a_36_216# INVX1_LOC_266/Y 0.00fF
C47661 NOR2X1_LOC_152/Y NAND2X1_LOC_848/A 0.01fF
C47662 D_INPUT_0 INVX1_LOC_158/Y 0.41fF
C47663 INVX1_LOC_230/Y INVX1_LOC_3/A 0.14fF
C47664 NOR2X1_LOC_68/A NAND2X1_LOC_434/Y 0.08fF
C47665 NOR2X1_LOC_666/A NOR2X1_LOC_89/A 0.01fF
C47666 NOR2X1_LOC_507/A NOR2X1_LOC_78/A 0.07fF
C47667 INVX1_LOC_120/A INPUT_0 0.02fF
C47668 NOR2X1_LOC_708/Y INVX1_LOC_75/A 0.01fF
C47669 NAND2X1_LOC_350/B NAND2X1_LOC_468/B 0.00fF
C47670 NOR2X1_LOC_533/Y INVX1_LOC_49/Y 0.00fF
C47671 NOR2X1_LOC_82/A INVX1_LOC_19/A 0.10fF
C47672 INVX1_LOC_134/A INVX1_LOC_19/A 0.01fF
C47673 INVX1_LOC_24/A NOR2X1_LOC_487/Y 0.01fF
C47674 INVX1_LOC_25/A NAND2X1_LOC_99/A 0.09fF
C47675 NOR2X1_LOC_788/B NOR2X1_LOC_74/A 0.02fF
C47676 INVX1_LOC_23/A NOR2X1_LOC_798/Y 0.01fF
C47677 NOR2X1_LOC_577/Y INVX1_LOC_9/A 0.01fF
C47678 INVX1_LOC_208/A NAND2X1_LOC_468/B 0.01fF
C47679 INVX1_LOC_54/Y VDD 0.77fF
C47680 NAND2X1_LOC_214/B INVX1_LOC_4/Y 0.01fF
C47681 VDD NOR2X1_LOC_353/Y 0.24fF
C47682 INVX1_LOC_244/Y INVX1_LOC_92/A 0.02fF
C47683 NAND2X1_LOC_724/Y INVX1_LOC_296/Y 0.05fF
C47684 NAND2X1_LOC_181/Y INVX1_LOC_20/A 0.92fF
C47685 INVX1_LOC_41/A NOR2X1_LOC_271/Y 0.11fF
C47686 NOR2X1_LOC_323/Y NAND2X1_LOC_807/Y 0.03fF
C47687 NOR2X1_LOC_528/Y NOR2X1_LOC_528/a_36_216# 0.00fF
C47688 INVX1_LOC_123/A NOR2X1_LOC_99/B 0.07fF
C47689 NAND2X1_LOC_67/Y INVX1_LOC_283/A 0.11fF
C47690 INVX1_LOC_23/A INVX1_LOC_275/Y 0.05fF
C47691 NOR2X1_LOC_446/A INVX1_LOC_29/A 0.01fF
C47692 NAND2X1_LOC_722/A NAND2X1_LOC_804/Y 0.36fF
C47693 INVX1_LOC_23/A NOR2X1_LOC_748/A 0.10fF
C47694 INVX1_LOC_259/A INVX1_LOC_117/A 0.03fF
C47695 D_INPUT_1 NAND2X1_LOC_215/A 0.07fF
C47696 NOR2X1_LOC_375/Y NOR2X1_LOC_480/a_36_216# 0.00fF
C47697 INVX1_LOC_83/A INVX1_LOC_91/A 6.67fF
C47698 NOR2X1_LOC_15/Y NOR2X1_LOC_270/a_36_216# 0.00fF
C47699 NOR2X1_LOC_107/Y NOR2X1_LOC_89/A 0.01fF
C47700 INVX1_LOC_25/Y INVX1_LOC_76/A 0.03fF
C47701 NAND2X1_LOC_20/B GATE_222 0.01fF
C47702 INVX1_LOC_178/A NAND2X1_LOC_618/Y 0.01fF
C47703 INVX1_LOC_27/A INVX1_LOC_4/Y 0.67fF
C47704 INVX1_LOC_5/A NOR2X1_LOC_631/Y 0.10fF
C47705 NAND2X1_LOC_716/a_36_24# INVX1_LOC_76/A 0.01fF
C47706 NAND2X1_LOC_360/a_36_24# NAND2X1_LOC_99/A 0.01fF
C47707 NAND2X1_LOC_349/B INVX1_LOC_76/A 0.10fF
C47708 NAND2X1_LOC_36/A INVX1_LOC_19/A 0.01fF
C47709 NOR2X1_LOC_348/B INVX1_LOC_9/A 0.03fF
C47710 NOR2X1_LOC_68/A NAND2X1_LOC_206/Y 0.05fF
C47711 NOR2X1_LOC_787/a_36_216# INVX1_LOC_290/Y 0.00fF
C47712 NAND2X1_LOC_390/A INVX1_LOC_20/A 0.12fF
C47713 NOR2X1_LOC_743/a_36_216# INVX1_LOC_131/Y 0.00fF
C47714 NOR2X1_LOC_91/A NOR2X1_LOC_304/Y 0.04fF
C47715 NOR2X1_LOC_593/Y NOR2X1_LOC_79/Y 0.03fF
C47716 NAND2X1_LOC_276/Y INVX1_LOC_92/A 0.00fF
C47717 INVX1_LOC_31/A INVX1_LOC_106/Y 0.01fF
C47718 INVX1_LOC_14/A NOR2X1_LOC_38/B 0.23fF
C47719 NOR2X1_LOC_134/Y INVX1_LOC_42/A 0.00fF
C47720 NOR2X1_LOC_249/Y NOR2X1_LOC_33/Y 0.00fF
C47721 NAND2X1_LOC_326/A INVX1_LOC_94/Y 0.64fF
C47722 NOR2X1_LOC_717/A NOR2X1_LOC_292/a_36_216# 0.01fF
C47723 NOR2X1_LOC_561/Y NAND2X1_LOC_453/A 0.05fF
C47724 NOR2X1_LOC_464/a_36_216# NOR2X1_LOC_155/A 0.00fF
C47725 INVX1_LOC_174/Y NOR2X1_LOC_706/B 0.00fF
C47726 NOR2X1_LOC_366/B NOR2X1_LOC_331/B 0.03fF
C47727 INVX1_LOC_33/A NOR2X1_LOC_117/Y 0.01fF
C47728 NOR2X1_LOC_209/A INVX1_LOC_85/Y 0.00fF
C47729 NOR2X1_LOC_589/A INVX1_LOC_117/A 0.15fF
C47730 INVX1_LOC_313/Y INVX1_LOC_247/A 0.02fF
C47731 NOR2X1_LOC_773/Y INVX1_LOC_118/A 0.10fF
C47732 NOR2X1_LOC_335/B NOR2X1_LOC_501/B 0.02fF
C47733 NAND2X1_LOC_198/B NAND2X1_LOC_74/B 0.01fF
C47734 INVX1_LOC_41/A NAND2X1_LOC_252/a_36_24# 0.01fF
C47735 NOR2X1_LOC_19/B INVX1_LOC_316/A 0.00fF
C47736 INVX1_LOC_77/A INVX1_LOC_186/Y 0.24fF
C47737 INVX1_LOC_58/A NOR2X1_LOC_626/Y 0.36fF
C47738 NOR2X1_LOC_325/A INVX1_LOC_9/A 0.00fF
C47739 INVX1_LOC_1/A NAND2X1_LOC_99/A 0.10fF
C47740 NOR2X1_LOC_172/Y INVX1_LOC_63/A 0.03fF
C47741 INVX1_LOC_22/A INVX1_LOC_9/A 0.10fF
C47742 NAND2X1_LOC_338/B NOR2X1_LOC_862/B 0.10fF
C47743 INVX1_LOC_34/A NOR2X1_LOC_631/A 0.02fF
C47744 NOR2X1_LOC_78/A NOR2X1_LOC_83/Y 0.12fF
C47745 INVX1_LOC_11/A INVX1_LOC_26/A 0.03fF
C47746 INVX1_LOC_21/A NAND2X1_LOC_787/A 0.03fF
C47747 NOR2X1_LOC_134/Y INVX1_LOC_78/A 0.00fF
C47748 NOR2X1_LOC_541/Y NOR2X1_LOC_541/B 0.03fF
C47749 INVX1_LOC_21/A NAND2X1_LOC_363/B 0.07fF
C47750 INVX1_LOC_233/A NAND2X1_LOC_391/Y 0.01fF
C47751 NOR2X1_LOC_6/B NOR2X1_LOC_673/a_36_216# 0.00fF
C47752 NOR2X1_LOC_112/Y VDD 0.14fF
C47753 INVX1_LOC_33/A INVX1_LOC_301/A 0.05fF
C47754 NAND2X1_LOC_563/Y NOR2X1_LOC_662/A 0.15fF
C47755 NAND2X1_LOC_861/Y NAND2X1_LOC_848/A 0.10fF
C47756 INVX1_LOC_233/Y NOR2X1_LOC_824/A 0.10fF
C47757 NAND2X1_LOC_317/a_36_24# INVX1_LOC_118/A 0.00fF
C47758 INVX1_LOC_75/A INVX1_LOC_76/A 0.87fF
C47759 NAND2X1_LOC_660/Y INVX1_LOC_291/A 0.06fF
C47760 GATE_479 NAND2X1_LOC_93/B 0.07fF
C47761 INVX1_LOC_35/A INVX1_LOC_48/Y 0.03fF
C47762 INVX1_LOC_39/A INVX1_LOC_5/A 0.01fF
C47763 NOR2X1_LOC_68/A NOR2X1_LOC_297/A 0.01fF
C47764 INVX1_LOC_278/A NAND2X1_LOC_579/A 0.10fF
C47765 INVX1_LOC_36/A NAND2X1_LOC_223/A 0.03fF
C47766 INVX1_LOC_233/Y INVX1_LOC_237/A 0.05fF
C47767 NOR2X1_LOC_311/Y INVX1_LOC_91/A 0.01fF
C47768 INVX1_LOC_34/A NAND2X1_LOC_469/a_36_24# 0.00fF
C47769 INVX1_LOC_136/A NAND2X1_LOC_72/B 0.04fF
C47770 NOR2X1_LOC_91/A NAND2X1_LOC_711/Y 0.15fF
C47771 GATE_479 NAND2X1_LOC_425/Y 0.07fF
C47772 NOR2X1_LOC_364/Y INVX1_LOC_109/Y -0.01fF
C47773 INVX1_LOC_155/A NOR2X1_LOC_114/Y 0.02fF
C47774 INVX1_LOC_43/A INVX1_LOC_84/A 0.07fF
C47775 NAND2X1_LOC_116/A INVX1_LOC_29/A 0.07fF
C47776 INVX1_LOC_21/A NOR2X1_LOC_791/Y 0.13fF
C47777 NOR2X1_LOC_590/A NOR2X1_LOC_727/B 0.06fF
C47778 INVX1_LOC_45/A NOR2X1_LOC_541/B 0.00fF
C47779 INPUT_0 NOR2X1_LOC_137/Y 0.03fF
C47780 NOR2X1_LOC_6/B NOR2X1_LOC_610/a_36_216# 0.01fF
C47781 NOR2X1_LOC_592/A INVX1_LOC_53/A 0.01fF
C47782 NOR2X1_LOC_568/A NOR2X1_LOC_541/B 0.11fF
C47783 INVX1_LOC_38/Y NAND2X1_LOC_473/A 0.06fF
C47784 INVX1_LOC_31/A NOR2X1_LOC_748/A 0.35fF
C47785 NAND2X1_LOC_740/B NOR2X1_LOC_536/A 0.02fF
C47786 NOR2X1_LOC_709/A INVX1_LOC_12/A 0.09fF
C47787 NAND2X1_LOC_634/Y INVX1_LOC_23/Y 0.45fF
C47788 NOR2X1_LOC_15/Y NAND2X1_LOC_169/Y 0.01fF
C47789 NOR2X1_LOC_516/B NOR2X1_LOC_820/B 0.05fF
C47790 INVX1_LOC_309/A INVX1_LOC_46/A 0.01fF
C47791 NOR2X1_LOC_354/Y VDD 0.00fF
C47792 NAND2X1_LOC_581/a_36_24# INVX1_LOC_174/A 0.01fF
C47793 NOR2X1_LOC_114/A INVX1_LOC_46/A 0.05fF
C47794 NOR2X1_LOC_188/A NAND2X1_LOC_96/A 0.07fF
C47795 NOR2X1_LOC_591/Y NOR2X1_LOC_48/B 0.02fF
C47796 NOR2X1_LOC_773/Y NAND2X1_LOC_63/Y 0.00fF
C47797 INVX1_LOC_140/A INVX1_LOC_118/A 1.51fF
C47798 INVX1_LOC_312/Y NOR2X1_LOC_441/a_36_216# 0.00fF
C47799 NOR2X1_LOC_590/A NOR2X1_LOC_717/A 0.12fF
C47800 INVX1_LOC_279/A NOR2X1_LOC_127/Y -0.02fF
C47801 NAND2X1_LOC_623/B INVX1_LOC_20/A 0.04fF
C47802 NOR2X1_LOC_548/B NAND2X1_LOC_96/A 0.03fF
C47803 INVX1_LOC_2/A INVX1_LOC_42/A 0.22fF
C47804 NAND2X1_LOC_364/A NOR2X1_LOC_113/a_36_216# 0.00fF
C47805 NOR2X1_LOC_214/B INVX1_LOC_107/Y 0.03fF
C47806 INVX1_LOC_213/Y INVX1_LOC_15/A 0.47fF
C47807 INVX1_LOC_49/A INVX1_LOC_78/A 0.47fF
C47808 INVX1_LOC_91/A INVX1_LOC_46/A 2.86fF
C47809 NOR2X1_LOC_772/B NOR2X1_LOC_160/B 0.01fF
C47810 NOR2X1_LOC_238/Y NOR2X1_LOC_693/Y 0.03fF
C47811 NOR2X1_LOC_459/A INVX1_LOC_203/A 0.02fF
C47812 NOR2X1_LOC_226/A INVX1_LOC_42/A 0.09fF
C47813 INVX1_LOC_53/Y NAND2X1_LOC_74/B 0.03fF
C47814 NOR2X1_LOC_322/Y INVX1_LOC_185/A 0.02fF
C47815 NOR2X1_LOC_775/Y NOR2X1_LOC_634/A 0.54fF
C47816 INVX1_LOC_13/Y NAND2X1_LOC_550/A 0.34fF
C47817 NOR2X1_LOC_619/A NAND2X1_LOC_74/B 0.12fF
C47818 NOR2X1_LOC_664/Y INVX1_LOC_4/Y 1.08fF
C47819 INVX1_LOC_21/A NOR2X1_LOC_457/A 0.04fF
C47820 NOR2X1_LOC_433/A INVX1_LOC_26/A 0.01fF
C47821 NOR2X1_LOC_346/B NOR2X1_LOC_861/Y 0.15fF
C47822 INVX1_LOC_13/Y NOR2X1_LOC_160/B 0.14fF
C47823 NAND2X1_LOC_562/B NAND2X1_LOC_618/Y 0.18fF
C47824 INVX1_LOC_181/Y INVX1_LOC_57/A 0.05fF
C47825 NOR2X1_LOC_716/B NOR2X1_LOC_301/A 0.01fF
C47826 INVX1_LOC_11/Y INVX1_LOC_46/A 0.10fF
C47827 NOR2X1_LOC_468/Y INVX1_LOC_14/A 0.14fF
C47828 NAND2X1_LOC_468/B NAND2X1_LOC_211/Y 0.03fF
C47829 NAND2X1_LOC_35/Y INVX1_LOC_170/A 0.05fF
C47830 INVX1_LOC_97/A INVX1_LOC_63/A 0.03fF
C47831 NOR2X1_LOC_65/B INVX1_LOC_49/A 1.43fF
C47832 NAND2X1_LOC_547/a_36_24# NOR2X1_LOC_654/A 0.00fF
C47833 INVX1_LOC_20/A NOR2X1_LOC_422/Y 0.01fF
C47834 INVX1_LOC_234/A NAND2X1_LOC_81/B 0.01fF
C47835 INVX1_LOC_206/A INVX1_LOC_4/Y 0.70fF
C47836 INPUT_5 NOR2X1_LOC_17/a_36_216# 0.00fF
C47837 NOR2X1_LOC_848/a_36_216# INVX1_LOC_31/A 0.00fF
C47838 INVX1_LOC_72/A NOR2X1_LOC_53/Y 0.26fF
C47839 NOR2X1_LOC_172/Y NOR2X1_LOC_65/Y 0.02fF
C47840 INVX1_LOC_90/A INVX1_LOC_63/A 0.27fF
C47841 NOR2X1_LOC_292/Y NAND2X1_LOC_93/B 0.05fF
C47842 INVX1_LOC_8/A INVX1_LOC_23/Y 2.17fF
C47843 NAND2X1_LOC_453/A INVX1_LOC_76/A 0.03fF
C47844 INVX1_LOC_289/Y INVX1_LOC_161/Y 0.03fF
C47845 NOR2X1_LOC_389/B INVX1_LOC_63/A 0.08fF
C47846 INVX1_LOC_11/Y NOR2X1_LOC_766/Y 0.06fF
C47847 INVX1_LOC_33/A INVX1_LOC_270/A 0.10fF
C47848 INVX1_LOC_2/A INVX1_LOC_78/A 8.66fF
C47849 NOR2X1_LOC_52/B INVX1_LOC_26/A 0.07fF
C47850 INVX1_LOC_269/A INVX1_LOC_150/Y 0.10fF
C47851 INVX1_LOC_39/A NOR2X1_LOC_90/a_36_216# 0.00fF
C47852 NAND2X1_LOC_462/B INVX1_LOC_42/A 0.06fF
C47853 INVX1_LOC_21/A INVX1_LOC_30/A 0.22fF
C47854 NOR2X1_LOC_285/A INVX1_LOC_310/Y 0.05fF
C47855 INVX1_LOC_224/A NOR2X1_LOC_107/Y 0.01fF
C47856 NAND2X1_LOC_200/B INVX1_LOC_4/Y 0.01fF
C47857 INVX1_LOC_20/A INVX1_LOC_117/A 0.03fF
C47858 NAND2X1_LOC_222/A NOR2X1_LOC_6/B 0.02fF
C47859 NOR2X1_LOC_226/A INVX1_LOC_78/A 0.11fF
C47860 NOR2X1_LOC_334/A NAND2X1_LOC_238/a_36_24# 0.01fF
C47861 INVX1_LOC_27/A NOR2X1_LOC_723/Y 0.03fF
C47862 INVX1_LOC_88/A NOR2X1_LOC_160/B 0.06fF
C47863 NOR2X1_LOC_388/Y NOR2X1_LOC_493/A 0.04fF
C47864 INVX1_LOC_58/A NOR2X1_LOC_433/a_36_216# 0.00fF
C47865 NOR2X1_LOC_76/a_36_216# NAND2X1_LOC_74/B 0.00fF
C47866 D_INPUT_1 NOR2X1_LOC_142/Y 0.10fF
C47867 NOR2X1_LOC_500/Y NOR2X1_LOC_334/Y 1.01fF
C47868 NAND2X1_LOC_577/A INVX1_LOC_1/A 0.28fF
C47869 NAND2X1_LOC_348/A INVX1_LOC_63/A 0.10fF
C47870 INVX1_LOC_286/Y NAND2X1_LOC_537/Y 0.09fF
C47871 NOR2X1_LOC_15/Y NOR2X1_LOC_372/a_36_216# 0.00fF
C47872 NAND2X1_LOC_341/A NAND2X1_LOC_470/B 0.01fF
C47873 NOR2X1_LOC_75/Y NOR2X1_LOC_471/Y 0.05fF
C47874 INVX1_LOC_35/A NOR2X1_LOC_460/B 0.01fF
C47875 NOR2X1_LOC_620/Y INVX1_LOC_64/A 0.03fF
C47876 INVX1_LOC_137/A INVX1_LOC_4/Y 0.07fF
C47877 NAND2X1_LOC_648/A INVX1_LOC_42/A 0.85fF
C47878 NOR2X1_LOC_570/B NOR2X1_LOC_678/A 0.27fF
C47879 NOR2X1_LOC_78/A NOR2X1_LOC_155/A 0.19fF
C47880 NOR2X1_LOC_454/Y INVX1_LOC_18/A 0.83fF
C47881 INVX1_LOC_191/Y NOR2X1_LOC_635/B 0.04fF
C47882 INVX1_LOC_119/A INVX1_LOC_23/A 0.10fF
C47883 INVX1_LOC_200/Y NAND2X1_LOC_785/A 0.00fF
C47884 INPUT_1 INVX1_LOC_42/A 0.18fF
C47885 INVX1_LOC_292/A INVX1_LOC_225/Y 0.06fF
C47886 NOR2X1_LOC_721/Y NOR2X1_LOC_721/B 0.11fF
C47887 NOR2X1_LOC_65/B NOR2X1_LOC_226/A 0.07fF
C47888 INVX1_LOC_33/A NOR2X1_LOC_109/Y 0.04fF
C47889 NAND2X1_LOC_785/Y NAND2X1_LOC_787/A 0.81fF
C47890 NAND2X1_LOC_832/Y INVX1_LOC_186/Y 0.01fF
C47891 NOR2X1_LOC_411/A NAND2X1_LOC_33/Y 0.29fF
C47892 NOR2X1_LOC_501/B INVX1_LOC_84/A 0.01fF
C47893 INVX1_LOC_10/A NOR2X1_LOC_334/Y 0.14fF
C47894 NOR2X1_LOC_252/a_36_216# NOR2X1_LOC_693/Y 0.00fF
C47895 NOR2X1_LOC_454/Y NOR2X1_LOC_637/Y 0.02fF
C47896 D_INPUT_1 NOR2X1_LOC_655/B 0.13fF
C47897 NOR2X1_LOC_401/B INVX1_LOC_23/A 0.02fF
C47898 NOR2X1_LOC_689/Y NAND2X1_LOC_724/a_36_24# 0.00fF
C47899 INVX1_LOC_1/A NAND2X1_LOC_656/A 0.03fF
C47900 NOR2X1_LOC_142/Y NOR2X1_LOC_108/a_36_216# 0.01fF
C47901 NOR2X1_LOC_160/B NOR2X1_LOC_500/B 0.10fF
C47902 INVX1_LOC_35/A NAND2X1_LOC_359/Y 0.06fF
C47903 INVX1_LOC_226/Y NAND2X1_LOC_464/B 0.11fF
C47904 NOR2X1_LOC_381/Y NOR2X1_LOC_8/a_36_216# 0.00fF
C47905 NOR2X1_LOC_428/Y INVX1_LOC_30/A 0.07fF
C47906 INVX1_LOC_10/Y NOR2X1_LOC_331/B 0.05fF
C47907 NAND2X1_LOC_30/Y NAND2X1_LOC_36/a_36_24# 0.00fF
C47908 NAND2X1_LOC_787/A NOR2X1_LOC_667/A 0.00fF
C47909 INVX1_LOC_35/A INVX1_LOC_216/A 0.03fF
C47910 VDD NOR2X1_LOC_78/Y 0.42fF
C47911 INVX1_LOC_58/A NOR2X1_LOC_418/Y 0.06fF
C47912 NOR2X1_LOC_690/A NOR2X1_LOC_496/Y 0.06fF
C47913 NAND2X1_LOC_514/Y INVX1_LOC_161/Y 0.02fF
C47914 NOR2X1_LOC_682/Y INVX1_LOC_291/A 0.02fF
C47915 VDD NAND2X1_LOC_656/B 0.01fF
C47916 INVX1_LOC_249/A NOR2X1_LOC_205/Y 0.70fF
C47917 NAND2X1_LOC_562/Y INVX1_LOC_178/A 0.58fF
C47918 INVX1_LOC_295/A NAND2X1_LOC_467/a_36_24# 0.01fF
C47919 GATE_741 GATE_811 0.02fF
C47920 INVX1_LOC_167/Y INVX1_LOC_163/Y 0.35fF
C47921 NAND2X1_LOC_648/A INVX1_LOC_78/A 0.00fF
C47922 NOR2X1_LOC_246/A NOR2X1_LOC_278/Y 0.11fF
C47923 NAND2X1_LOC_778/Y NAND2X1_LOC_357/B 0.01fF
C47924 INVX1_LOC_27/A INVX1_LOC_82/A 0.03fF
C47925 INVX1_LOC_313/Y NOR2X1_LOC_465/Y 0.03fF
C47926 INPUT_1 INVX1_LOC_78/A 0.06fF
C47927 VDD INVX1_LOC_35/Y 0.21fF
C47928 INVX1_LOC_279/A NOR2X1_LOC_383/B 0.14fF
C47929 NAND2X1_LOC_802/A INVX1_LOC_103/A 0.01fF
C47930 INVX1_LOC_17/A NOR2X1_LOC_419/Y 0.02fF
C47931 INVX1_LOC_201/Y INVX1_LOC_239/A 0.04fF
C47932 INVX1_LOC_58/A NOR2X1_LOC_589/A 0.18fF
C47933 NAND2X1_LOC_577/A NOR2X1_LOC_384/Y 0.01fF
C47934 NAND2X1_LOC_273/a_36_24# INVX1_LOC_46/A 0.00fF
C47935 NAND2X1_LOC_35/Y NAND2X1_LOC_852/Y 0.03fF
C47936 NAND2X1_LOC_848/A INVX1_LOC_291/A 0.14fF
C47937 INVX1_LOC_17/A NOR2X1_LOC_716/B 0.10fF
C47938 INVX1_LOC_89/A NOR2X1_LOC_668/Y 0.07fF
C47939 NOR2X1_LOC_305/Y INVX1_LOC_250/Y 0.22fF
C47940 NAND2X1_LOC_656/Y NOR2X1_LOC_441/a_36_216# 0.01fF
C47941 NAND2X1_LOC_385/a_36_24# INVX1_LOC_232/A 0.00fF
C47942 INVX1_LOC_50/A NOR2X1_LOC_355/A 0.00fF
C47943 NOR2X1_LOC_553/B INVX1_LOC_53/A 0.02fF
C47944 NOR2X1_LOC_178/Y INVX1_LOC_25/Y 0.07fF
C47945 INVX1_LOC_35/A INVX1_LOC_290/A 0.07fF
C47946 INVX1_LOC_2/A NOR2X1_LOC_215/A 0.04fF
C47947 NOR2X1_LOC_32/B NOR2X1_LOC_32/Y 0.04fF
C47948 NOR2X1_LOC_582/Y INVX1_LOC_30/A 0.06fF
C47949 NOR2X1_LOC_15/Y NAND2X1_LOC_357/B 0.07fF
C47950 INVX1_LOC_64/A NAND2X1_LOC_514/a_36_24# 0.01fF
C47951 INVX1_LOC_303/A NOR2X1_LOC_160/B 1.11fF
C47952 INVX1_LOC_59/Y INVX1_LOC_19/A 0.07fF
C47953 NOR2X1_LOC_45/B NOR2X1_LOC_226/Y 0.01fF
C47954 INVX1_LOC_150/A INVX1_LOC_23/A 0.00fF
C47955 INVX1_LOC_148/Y INVX1_LOC_57/A 0.12fF
C47956 D_INPUT_1 NOR2X1_LOC_99/B 0.07fF
C47957 INVX1_LOC_74/Y INVX1_LOC_29/A 0.01fF
C47958 INVX1_LOC_11/A INVX1_LOC_103/Y 0.01fF
C47959 NOR2X1_LOC_270/Y INVX1_LOC_72/A 0.02fF
C47960 NOR2X1_LOC_815/Y NOR2X1_LOC_816/A 0.00fF
C47961 INVX1_LOC_227/A NOR2X1_LOC_717/A 0.36fF
C47962 NOR2X1_LOC_596/A NOR2X1_LOC_717/Y 0.02fF
C47963 INVX1_LOC_1/A NOR2X1_LOC_423/Y 0.01fF
C47964 NOR2X1_LOC_468/Y NOR2X1_LOC_612/B 0.26fF
C47965 INVX1_LOC_203/A INVX1_LOC_46/A 0.04fF
C47966 INVX1_LOC_58/A INVX1_LOC_171/A 0.03fF
C47967 NOR2X1_LOC_201/A NAND2X1_LOC_508/A 0.10fF
C47968 NAND2X1_LOC_447/Y INVX1_LOC_29/A 0.03fF
C47969 NAND2X1_LOC_715/B NAND2X1_LOC_112/Y 0.06fF
C47970 NOR2X1_LOC_607/A INVX1_LOC_223/A 0.03fF
C47971 NOR2X1_LOC_824/A NOR2X1_LOC_526/Y 0.06fF
C47972 INVX1_LOC_161/Y NAND2X1_LOC_332/Y 0.02fF
C47973 VDD NOR2X1_LOC_721/B 0.40fF
C47974 INVX1_LOC_136/A NAND2X1_LOC_198/B 0.17fF
C47975 NOR2X1_LOC_473/B INVX1_LOC_270/Y 0.28fF
C47976 INVX1_LOC_89/A INVX1_LOC_23/A 4.97fF
C47977 NOR2X1_LOC_590/A NAND2X1_LOC_364/Y 0.02fF
C47978 INVX1_LOC_5/A NAND2X1_LOC_735/B 1.11fF
C47979 NAND2X1_LOC_465/A NAND2X1_LOC_74/B 0.01fF
C47980 NAND2X1_LOC_53/Y NOR2X1_LOC_718/B 0.06fF
C47981 INVX1_LOC_233/Y INVX1_LOC_234/A 0.12fF
C47982 INVX1_LOC_162/Y NAND2X1_LOC_793/Y 0.03fF
C47983 INVX1_LOC_48/A NOR2X1_LOC_38/B 0.07fF
C47984 NOR2X1_LOC_401/A INVX1_LOC_168/A 0.16fF
C47985 INVX1_LOC_103/A INVX1_LOC_266/Y 0.10fF
C47986 NOR2X1_LOC_590/A NAND2X1_LOC_175/B 0.07fF
C47987 INVX1_LOC_50/A NOR2X1_LOC_736/Y 0.04fF
C47988 NOR2X1_LOC_68/A INVX1_LOC_24/A 0.29fF
C47989 INVX1_LOC_182/Y NOR2X1_LOC_383/B 0.03fF
C47990 NOR2X1_LOC_222/Y INVX1_LOC_1/A 0.07fF
C47991 INVX1_LOC_269/A NAND2X1_LOC_165/a_36_24# 0.00fF
C47992 INVX1_LOC_233/A INVX1_LOC_183/Y 0.01fF
C47993 INVX1_LOC_251/Y NOR2X1_LOC_103/Y 0.00fF
C47994 INVX1_LOC_178/A NAND2X1_LOC_735/B 0.05fF
C47995 INVX1_LOC_314/Y NOR2X1_LOC_360/Y 0.07fF
C47996 INVX1_LOC_77/A INVX1_LOC_18/A 1.10fF
C47997 INVX1_LOC_48/Y NOR2X1_LOC_121/A 0.02fF
C47998 INVX1_LOC_36/A INVX1_LOC_33/A 0.13fF
C47999 D_INPUT_1 INVX1_LOC_182/A 0.03fF
C48000 INVX1_LOC_38/A INVX1_LOC_63/A 0.10fF
C48001 VDD NOR2X1_LOC_610/Y 0.12fF
C48002 INVX1_LOC_12/Y INVX1_LOC_272/A 0.22fF
C48003 INVX1_LOC_141/A NOR2X1_LOC_52/B 0.01fF
C48004 NOR2X1_LOC_160/B INVX1_LOC_168/A 0.02fF
C48005 INVX1_LOC_2/A NOR2X1_LOC_503/Y 0.07fF
C48006 INVX1_LOC_292/A INVX1_LOC_266/Y 0.00fF
C48007 INVX1_LOC_208/A INVX1_LOC_88/A 0.10fF
C48008 INVX1_LOC_119/A INVX1_LOC_31/A 1.31fF
C48009 INVX1_LOC_76/A INVX1_LOC_283/A 0.04fF
C48010 INVX1_LOC_30/Y NAND2X1_LOC_347/B 0.17fF
C48011 NAND2X1_LOC_361/Y NAND2X1_LOC_364/A 0.05fF
C48012 INVX1_LOC_186/Y INVX1_LOC_9/A 0.07fF
C48013 INVX1_LOC_236/Y INVX1_LOC_236/A 0.10fF
C48014 INVX1_LOC_20/A INVX1_LOC_3/Y 0.42fF
C48015 INVX1_LOC_175/Y INVX1_LOC_253/Y 0.21fF
C48016 NOR2X1_LOC_795/Y INVX1_LOC_45/A 0.00fF
C48017 NAND2X1_LOC_181/Y INVX1_LOC_43/Y 0.00fF
C48018 INVX1_LOC_239/A NOR2X1_LOC_299/Y 0.02fF
C48019 NOR2X1_LOC_481/A INVX1_LOC_94/A 0.06fF
C48020 INVX1_LOC_58/A INVX1_LOC_222/A 0.07fF
C48021 NOR2X1_LOC_31/a_36_216# D_INPUT_5 0.00fF
C48022 NAND2X1_LOC_833/Y INVX1_LOC_41/Y 0.34fF
C48023 INVX1_LOC_145/A INVX1_LOC_33/A 0.01fF
C48024 INVX1_LOC_49/A NOR2X1_LOC_152/Y 0.08fF
C48025 NOR2X1_LOC_396/Y NOR2X1_LOC_395/Y 0.09fF
C48026 INVX1_LOC_49/A INVX1_LOC_113/Y 0.03fF
C48027 NOR2X1_LOC_458/Y NOR2X1_LOC_303/Y 0.03fF
C48028 NOR2X1_LOC_564/Y INVX1_LOC_50/Y 0.06fF
C48029 INVX1_LOC_124/A INVX1_LOC_18/A 0.19fF
C48030 NAND2X1_LOC_722/A NOR2X1_LOC_517/Y 0.05fF
C48031 NOR2X1_LOC_667/A INVX1_LOC_30/A 0.42fF
C48032 NOR2X1_LOC_607/Y NOR2X1_LOC_142/Y 0.01fF
C48033 NOR2X1_LOC_334/Y NOR2X1_LOC_850/a_36_216# 0.01fF
C48034 INVX1_LOC_11/A INVX1_LOC_164/A 0.06fF
C48035 INVX1_LOC_122/Y INVX1_LOC_210/A 0.48fF
C48036 NOR2X1_LOC_818/Y NOR2X1_LOC_554/B 0.30fF
C48037 INVX1_LOC_238/A GATE_865 0.22fF
C48038 NOR2X1_LOC_848/Y INVX1_LOC_135/A 0.06fF
C48039 NOR2X1_LOC_794/B INVX1_LOC_220/Y 0.03fF
C48040 NAND2X1_LOC_208/B INVX1_LOC_56/Y 0.01fF
C48041 NOR2X1_LOC_592/a_36_216# NOR2X1_LOC_561/Y 0.01fF
C48042 NOR2X1_LOC_739/Y INVX1_LOC_83/A 0.03fF
C48043 NOR2X1_LOC_405/A NOR2X1_LOC_113/a_36_216# 0.01fF
C48044 NAND2X1_LOC_714/B INVX1_LOC_28/A 0.01fF
C48045 INVX1_LOC_125/A INVX1_LOC_92/A 0.85fF
C48046 INVX1_LOC_36/A INVX1_LOC_40/A 0.06fF
C48047 NAND2X1_LOC_725/B NOR2X1_LOC_395/a_36_216# -0.00fF
C48048 NOR2X1_LOC_78/A NOR2X1_LOC_125/Y 0.05fF
C48049 NOR2X1_LOC_68/A INVX1_LOC_143/A 0.14fF
C48050 INVX1_LOC_118/A INVX1_LOC_42/A 0.55fF
C48051 INVX1_LOC_117/A INVX1_LOC_4/A 0.05fF
C48052 NOR2X1_LOC_471/Y NOR2X1_LOC_424/Y 0.04fF
C48053 NOR2X1_LOC_500/A INVX1_LOC_177/A 0.13fF
C48054 NOR2X1_LOC_516/B NOR2X1_LOC_500/B 0.01fF
C48055 NOR2X1_LOC_675/A INVX1_LOC_57/A 0.00fF
C48056 NOR2X1_LOC_303/Y INVX1_LOC_177/A 0.29fF
C48057 INVX1_LOC_176/A INVX1_LOC_26/Y 0.06fF
C48058 NAND2X1_LOC_67/Y NOR2X1_LOC_735/Y 0.01fF
C48059 NOR2X1_LOC_214/a_36_216# NOR2X1_LOC_52/B 0.00fF
C48060 NOR2X1_LOC_598/B NOR2X1_LOC_78/A 0.19fF
C48061 NOR2X1_LOC_793/Y NOR2X1_LOC_356/A 0.10fF
C48062 NAND2X1_LOC_633/Y NOR2X1_LOC_301/A 0.01fF
C48063 NAND2X1_LOC_9/Y INVX1_LOC_91/A 0.06fF
C48064 NOR2X1_LOC_309/Y INVX1_LOC_33/A 0.03fF
C48065 VDD NOR2X1_LOC_829/A 0.04fF
C48066 INVX1_LOC_136/A INVX1_LOC_53/Y 0.01fF
C48067 NOR2X1_LOC_45/B NAND2X1_LOC_793/B 0.09fF
C48068 INVX1_LOC_233/A INVX1_LOC_91/A 1.11fF
C48069 INVX1_LOC_2/A NOR2X1_LOC_152/Y 0.52fF
C48070 NOR2X1_LOC_521/Y INVX1_LOC_30/A 0.00fF
C48071 NAND2X1_LOC_860/A NOR2X1_LOC_123/a_36_216# 0.00fF
C48072 NOR2X1_LOC_503/Y NAND2X1_LOC_648/A 0.01fF
C48073 INVX1_LOC_2/A INVX1_LOC_113/Y 0.03fF
C48074 INVX1_LOC_1/A D_INPUT_4 0.07fF
C48075 VDD NAND2X1_LOC_286/B 0.01fF
C48076 INVX1_LOC_240/A NAND2X1_LOC_811/Y 0.02fF
C48077 NAND2X1_LOC_562/Y NAND2X1_LOC_562/B 0.19fF
C48078 NOR2X1_LOC_226/A NOR2X1_LOC_152/Y 0.10fF
C48079 INVX1_LOC_5/A NOR2X1_LOC_7/Y 0.01fF
C48080 INVX1_LOC_38/A NAND2X1_LOC_452/Y 0.01fF
C48081 INVX1_LOC_149/A NOR2X1_LOC_593/Y 0.09fF
C48082 NAND2X1_LOC_787/A INVX1_LOC_304/A 0.39fF
C48083 NOR2X1_LOC_374/B NOR2X1_LOC_325/Y 0.11fF
C48084 NAND2X1_LOC_768/Y NAND2X1_LOC_773/B 0.34fF
C48085 INVX1_LOC_58/A INVX1_LOC_20/A 0.10fF
C48086 INVX1_LOC_89/A INVX1_LOC_31/A 0.49fF
C48087 INVX1_LOC_136/A NOR2X1_LOC_781/B 0.28fF
C48088 NOR2X1_LOC_295/Y NOR2X1_LOC_612/B 0.03fF
C48089 NOR2X1_LOC_456/Y NOR2X1_LOC_35/Y 0.10fF
C48090 NOR2X1_LOC_759/Y INVX1_LOC_16/A 0.05fF
C48091 INVX1_LOC_188/A NOR2X1_LOC_644/A 0.01fF
C48092 NOR2X1_LOC_52/B NOR2X1_LOC_369/a_36_216# 0.00fF
C48093 INVX1_LOC_12/A INVX1_LOC_294/A 0.03fF
C48094 INVX1_LOC_50/A NOR2X1_LOC_111/A 0.11fF
C48095 NOR2X1_LOC_798/A INVX1_LOC_91/A 0.03fF
C48096 INVX1_LOC_78/A INVX1_LOC_118/A 0.58fF
C48097 NOR2X1_LOC_816/A NAND2X1_LOC_680/a_36_24# 0.01fF
C48098 INVX1_LOC_225/A NOR2X1_LOC_312/a_36_216# 0.00fF
C48099 INVX1_LOC_303/A NOR2X1_LOC_516/B 0.10fF
C48100 NAND2X1_LOC_783/A NOR2X1_LOC_68/A 0.03fF
C48101 NAND2X1_LOC_785/Y NAND2X1_LOC_722/A 0.01fF
C48102 NAND2X1_LOC_508/A INVX1_LOC_31/A 3.27fF
C48103 NOR2X1_LOC_32/B NOR2X1_LOC_825/Y 0.14fF
C48104 NAND2X1_LOC_860/A VDD 1.57fF
C48105 NOR2X1_LOC_68/A NOR2X1_LOC_130/A 0.95fF
C48106 INVX1_LOC_161/A NOR2X1_LOC_385/Y 0.22fF
C48107 INVX1_LOC_5/A NAND2X1_LOC_212/Y 0.13fF
C48108 NOR2X1_LOC_471/Y NOR2X1_LOC_151/Y 0.01fF
C48109 NAND2X1_LOC_218/B INVX1_LOC_7/A 0.03fF
C48110 NOR2X1_LOC_454/a_36_216# INVX1_LOC_290/A 0.00fF
C48111 NOR2X1_LOC_334/Y INVX1_LOC_307/A 0.02fF
C48112 VDD NOR2X1_LOC_634/Y 0.24fF
C48113 NOR2X1_LOC_791/Y INVX1_LOC_304/A 0.26fF
C48114 NOR2X1_LOC_843/B INVX1_LOC_9/A 0.04fF
C48115 INVX1_LOC_34/A INVX1_LOC_56/Y 0.01fF
C48116 INVX1_LOC_179/A INVX1_LOC_271/Y 0.14fF
C48117 NAND2X1_LOC_733/Y NAND2X1_LOC_863/A 0.10fF
C48118 NOR2X1_LOC_227/B NOR2X1_LOC_349/A 0.06fF
C48119 NAND2X1_LOC_124/a_36_24# NOR2X1_LOC_276/Y 0.00fF
C48120 INVX1_LOC_232/A INVX1_LOC_8/A 0.10fF
C48121 NOR2X1_LOC_561/Y NOR2X1_LOC_577/Y 0.10fF
C48122 NOR2X1_LOC_65/B INVX1_LOC_118/A 0.02fF
C48123 NOR2X1_LOC_667/A NAND2X1_LOC_722/A 0.07fF
C48124 NAND2X1_LOC_735/a_36_24# INVX1_LOC_241/A 0.00fF
C48125 INVX1_LOC_41/Y NOR2X1_LOC_76/A 0.00fF
C48126 NOR2X1_LOC_392/B INVX1_LOC_1/Y 0.10fF
C48127 INVX1_LOC_5/A D_INPUT_3 0.73fF
C48128 INVX1_LOC_209/Y INVX1_LOC_10/A 0.08fF
C48129 NAND2X1_LOC_63/Y INVX1_LOC_42/A 0.03fF
C48130 INVX1_LOC_5/A INVX1_LOC_14/Y 0.10fF
C48131 NOR2X1_LOC_590/A NOR2X1_LOC_337/A 0.03fF
C48132 NAND2X1_LOC_350/A NAND2X1_LOC_814/a_36_24# 0.01fF
C48133 NOR2X1_LOC_367/B INVX1_LOC_22/A 0.08fF
C48134 INVX1_LOC_64/A INVX1_LOC_117/A 0.08fF
C48135 NAND2X1_LOC_508/A NAND2X1_LOC_106/a_36_24# 0.00fF
C48136 NAND2X1_LOC_51/B INVX1_LOC_30/A 0.05fF
C48137 NAND2X1_LOC_562/B NAND2X1_LOC_735/B 0.06fF
C48138 NOR2X1_LOC_103/Y NOR2X1_LOC_45/B 0.03fF
C48139 INVX1_LOC_209/Y NOR2X1_LOC_504/a_36_216# 0.00fF
C48140 NOR2X1_LOC_152/Y NAND2X1_LOC_648/A 0.02fF
C48141 NAND2X1_LOC_276/Y INVX1_LOC_83/A 0.01fF
C48142 NAND2X1_LOC_763/B NAND2X1_LOC_51/B 0.04fF
C48143 NOR2X1_LOC_860/B NOR2X1_LOC_702/Y 0.03fF
C48144 INVX1_LOC_28/A NOR2X1_LOC_759/Y 0.06fF
C48145 NOR2X1_LOC_226/A NAND2X1_LOC_860/Y 0.03fF
C48146 VDD INVX1_LOC_242/A 0.14fF
C48147 INVX1_LOC_57/Y NAND2X1_LOC_858/B 0.21fF
C48148 NOR2X1_LOC_299/Y GATE_811 0.03fF
C48149 NAND2X1_LOC_351/A INPUT_0 0.00fF
C48150 INVX1_LOC_104/A NAND2X1_LOC_656/Y 0.07fF
C48151 NAND2X1_LOC_223/A INVX1_LOC_63/A 0.03fF
C48152 VDD NAND2X1_LOC_473/A 0.20fF
C48153 NOR2X1_LOC_295/Y NOR2X1_LOC_137/A 0.02fF
C48154 INVX1_LOC_136/A NOR2X1_LOC_113/B 0.11fF
C48155 INVX1_LOC_226/Y INVX1_LOC_218/A 0.01fF
C48156 INVX1_LOC_54/A NOR2X1_LOC_678/A 0.03fF
C48157 NAND2X1_LOC_832/Y INVX1_LOC_18/A 0.11fF
C48158 INVX1_LOC_5/A INVX1_LOC_230/A 0.07fF
C48159 INVX1_LOC_232/Y INVX1_LOC_13/A 0.18fF
C48160 NAND2X1_LOC_833/Y NAND2X1_LOC_865/a_36_24# 0.01fF
C48161 INVX1_LOC_160/Y INVX1_LOC_134/Y 0.02fF
C48162 NOR2X1_LOC_131/a_36_216# INVX1_LOC_22/A 0.02fF
C48163 NAND2X1_LOC_390/A NAND2X1_LOC_850/Y 0.09fF
C48164 NOR2X1_LOC_418/a_36_216# INVX1_LOC_290/A 0.00fF
C48165 NOR2X1_LOC_78/B NOR2X1_LOC_553/B 0.01fF
C48166 INVX1_LOC_24/A NOR2X1_LOC_2/Y 0.03fF
C48167 NOR2X1_LOC_274/Y INVX1_LOC_75/A 0.04fF
C48168 INVX1_LOC_88/A NAND2X1_LOC_211/Y 0.03fF
C48169 NAND2X1_LOC_537/Y VDD -0.00fF
C48170 INVX1_LOC_77/A INVX1_LOC_31/Y 0.12fF
C48171 INVX1_LOC_78/A NAND2X1_LOC_63/Y 0.03fF
C48172 INVX1_LOC_45/A NOR2X1_LOC_45/B 0.10fF
C48173 NOR2X1_LOC_100/A INVX1_LOC_62/A 0.18fF
C48174 INVX1_LOC_12/Y NOR2X1_LOC_271/B 0.06fF
C48175 NOR2X1_LOC_569/Y NOR2X1_LOC_500/Y 0.01fF
C48176 NAND2X1_LOC_537/Y NAND2X1_LOC_800/A 0.06fF
C48177 INVX1_LOC_12/A NOR2X1_LOC_334/Y 0.15fF
C48178 NAND2X1_LOC_722/A NAND2X1_LOC_804/a_36_24# 0.00fF
C48179 NOR2X1_LOC_89/A NAND2X1_LOC_471/Y 0.02fF
C48180 INVX1_LOC_2/A NAND2X1_LOC_861/Y 0.07fF
C48181 INVX1_LOC_62/Y INVX1_LOC_48/A 0.01fF
C48182 NOR2X1_LOC_736/a_36_216# INVX1_LOC_63/Y 0.01fF
C48183 INVX1_LOC_34/A NOR2X1_LOC_385/Y 0.07fF
C48184 NOR2X1_LOC_753/Y NOR2X1_LOC_74/A 0.06fF
C48185 NAND2X1_LOC_301/a_36_24# NOR2X1_LOC_214/B 0.01fF
C48186 NOR2X1_LOC_19/B INVX1_LOC_82/A 0.01fF
C48187 NOR2X1_LOC_718/B NOR2X1_LOC_302/Y 0.05fF
C48188 INVX1_LOC_49/A INVX1_LOC_158/Y 0.07fF
C48189 NOR2X1_LOC_147/B NOR2X1_LOC_742/A 0.05fF
C48190 NOR2X1_LOC_226/A NAND2X1_LOC_861/Y 0.03fF
C48191 NOR2X1_LOC_360/Y NOR2X1_LOC_557/A 0.07fF
C48192 INVX1_LOC_30/A INVX1_LOC_304/A 0.10fF
C48193 NOR2X1_LOC_561/Y INVX1_LOC_22/A 0.15fF
C48194 NOR2X1_LOC_516/B INVX1_LOC_80/A 0.12fF
C48195 INVX1_LOC_86/Y NOR2X1_LOC_546/B 0.02fF
C48196 INVX1_LOC_36/A NOR2X1_LOC_486/Y 0.05fF
C48197 NOR2X1_LOC_573/Y VDD 0.00fF
C48198 INVX1_LOC_313/A NOR2X1_LOC_524/a_36_216# 0.01fF
C48199 NOR2X1_LOC_65/B NAND2X1_LOC_63/Y 0.03fF
C48200 INVX1_LOC_150/Y INVX1_LOC_12/Y 0.10fF
C48201 NOR2X1_LOC_32/B INVX1_LOC_84/A 0.89fF
C48202 INVX1_LOC_30/A NOR2X1_LOC_670/Y 0.00fF
C48203 NOR2X1_LOC_186/Y NOR2X1_LOC_155/A 0.15fF
C48204 NOR2X1_LOC_458/B INVX1_LOC_313/Y 0.02fF
C48205 NAND2X1_LOC_807/B NOR2X1_LOC_318/A 0.01fF
C48206 NOR2X1_LOC_848/Y INVX1_LOC_280/A 0.02fF
C48207 INVX1_LOC_26/A NAND2X1_LOC_254/Y 0.14fF
C48208 INVX1_LOC_27/A NOR2X1_LOC_156/Y 0.01fF
C48209 NOR2X1_LOC_440/Y NOR2X1_LOC_468/a_36_216# 0.00fF
C48210 NOR2X1_LOC_45/B INVX1_LOC_71/A 0.17fF
C48211 NAND2X1_LOC_150/a_36_24# INVX1_LOC_143/A -0.02fF
C48212 INVX1_LOC_43/Y INVX1_LOC_117/A 0.01fF
C48213 INVX1_LOC_18/A NOR2X1_LOC_670/a_36_216# 0.00fF
C48214 INVX1_LOC_213/Y NOR2X1_LOC_728/a_36_216# 0.02fF
C48215 INVX1_LOC_116/A NOR2X1_LOC_405/A 0.04fF
C48216 INVX1_LOC_21/Y NOR2X1_LOC_681/a_36_216# 0.00fF
C48217 NOR2X1_LOC_500/A INVX1_LOC_65/A 0.03fF
C48218 NOR2X1_LOC_338/Y INVX1_LOC_147/Y 0.15fF
C48219 INVX1_LOC_90/A INVX1_LOC_1/Y 0.10fF
C48220 INVX1_LOC_136/A NOR2X1_LOC_585/Y 0.09fF
C48221 NAND2X1_LOC_170/A NOR2X1_LOC_166/a_36_216# 0.00fF
C48222 NOR2X1_LOC_843/B NOR2X1_LOC_861/Y 0.07fF
C48223 INVX1_LOC_89/A NAND2X1_LOC_859/Y 0.03fF
C48224 NOR2X1_LOC_208/Y NOR2X1_LOC_486/Y 0.03fF
C48225 NOR2X1_LOC_389/B INVX1_LOC_1/Y 0.16fF
C48226 NAND2X1_LOC_866/A INVX1_LOC_11/Y 0.05fF
C48227 NOR2X1_LOC_68/A NOR2X1_LOC_280/Y 0.08fF
C48228 INVX1_LOC_71/A INVX1_LOC_247/A 0.03fF
C48229 NOR2X1_LOC_791/B INVX1_LOC_2/Y 0.01fF
C48230 INVX1_LOC_103/A NOR2X1_LOC_508/a_36_216# 0.00fF
C48231 NOR2X1_LOC_503/Y INVX1_LOC_118/A 0.03fF
C48232 NOR2X1_LOC_351/a_36_216# INVX1_LOC_76/A 0.01fF
C48233 NAND2X1_LOC_140/A NOR2X1_LOC_366/Y 0.27fF
C48234 INVX1_LOC_256/A NOR2X1_LOC_641/Y 0.01fF
C48235 NAND2X1_LOC_361/Y NOR2X1_LOC_405/A 0.01fF
C48236 NAND2X1_LOC_538/Y INVX1_LOC_92/A 0.07fF
C48237 NOR2X1_LOC_790/B INVX1_LOC_99/A 0.18fF
C48238 NOR2X1_LOC_392/Y NOR2X1_LOC_664/a_36_216# 0.00fF
C48239 INVX1_LOC_54/Y INVX1_LOC_285/Y 0.01fF
C48240 NOR2X1_LOC_392/B NOR2X1_LOC_318/B 0.07fF
C48241 NOR2X1_LOC_246/A NOR2X1_LOC_312/Y 0.11fF
C48242 NOR2X1_LOC_202/Y NAND2X1_LOC_479/Y 0.01fF
C48243 NOR2X1_LOC_690/A NOR2X1_LOC_823/Y 0.04fF
C48244 INVX1_LOC_78/A NOR2X1_LOC_631/Y 1.16fF
C48245 INVX1_LOC_135/A NOR2X1_LOC_560/A 0.00fF
C48246 NOR2X1_LOC_160/B NOR2X1_LOC_99/Y 0.19fF
C48247 NAND2X1_LOC_223/A NAND2X1_LOC_223/B 0.02fF
C48248 INVX1_LOC_45/A NOR2X1_LOC_499/B 0.03fF
C48249 NOR2X1_LOC_577/Y INVX1_LOC_76/A 0.18fF
C48250 NOR2X1_LOC_392/B INVX1_LOC_93/Y 0.10fF
C48251 NAND2X1_LOC_861/Y INPUT_1 0.07fF
C48252 INVX1_LOC_140/A INPUT_5 1.35fF
C48253 INPUT_0 INVX1_LOC_56/Y 0.04fF
C48254 NOR2X1_LOC_590/A NOR2X1_LOC_640/Y 0.13fF
C48255 INVX1_LOC_136/A NOR2X1_LOC_652/a_36_216# 0.01fF
C48256 NOR2X1_LOC_378/a_36_216# INVX1_LOC_91/A 0.00fF
C48257 NOR2X1_LOC_591/Y INVX1_LOC_291/Y 0.04fF
C48258 INVX1_LOC_58/A INVX1_LOC_4/A 0.25fF
C48259 INVX1_LOC_13/A NOR2X1_LOC_97/A 0.03fF
C48260 INVX1_LOC_135/A NOR2X1_LOC_346/a_36_216# 0.00fF
C48261 NOR2X1_LOC_32/B INVX1_LOC_15/A 0.42fF
C48262 INVX1_LOC_94/Y NOR2X1_LOC_654/A 0.10fF
C48263 INVX1_LOC_18/A INVX1_LOC_9/A 0.10fF
C48264 INVX1_LOC_1/A NOR2X1_LOC_691/B 0.07fF
C48265 INVX1_LOC_71/A INVX1_LOC_281/A 0.98fF
C48266 INVX1_LOC_35/A NOR2X1_LOC_467/A 0.12fF
C48267 INVX1_LOC_64/A INVX1_LOC_3/Y 0.98fF
C48268 NOR2X1_LOC_440/Y NOR2X1_LOC_292/Y 0.01fF
C48269 INVX1_LOC_35/A NOR2X1_LOC_801/B 0.02fF
C48270 NAND2X1_LOC_391/Y INVX1_LOC_284/A 0.00fF
C48271 NAND2X1_LOC_381/a_36_24# NOR2X1_LOC_649/B 0.00fF
C48272 NOR2X1_LOC_590/A NAND2X1_LOC_85/Y 0.62fF
C48273 VDD NOR2X1_LOC_486/B 0.00fF
C48274 VDD NOR2X1_LOC_516/Y 0.35fF
C48275 INVX1_LOC_45/A NOR2X1_LOC_862/B 0.10fF
C48276 INVX1_LOC_39/A INVX1_LOC_42/A 1.49fF
C48277 NAND2X1_LOC_382/a_36_24# NOR2X1_LOC_649/B 0.01fF
C48278 NOR2X1_LOC_590/A NOR2X1_LOC_697/Y 0.03fF
C48279 NOR2X1_LOC_191/A INVX1_LOC_95/A 0.00fF
C48280 INVX1_LOC_103/A INVX1_LOC_19/A 0.07fF
C48281 INVX1_LOC_90/A NOR2X1_LOC_742/A 0.07fF
C48282 NOR2X1_LOC_377/Y INVX1_LOC_14/Y 0.01fF
C48283 NOR2X1_LOC_389/A NOR2X1_LOC_127/Y 0.10fF
C48284 INVX1_LOC_135/A NOR2X1_LOC_391/B 0.14fF
C48285 INVX1_LOC_47/A NOR2X1_LOC_751/A 0.00fF
C48286 NOR2X1_LOC_152/Y INVX1_LOC_118/A 0.10fF
C48287 NOR2X1_LOC_68/A NOR2X1_LOC_197/B 0.37fF
C48288 INVX1_LOC_172/Y NAND2X1_LOC_659/B 0.02fF
C48289 INVX1_LOC_24/A NOR2X1_LOC_695/a_36_216# 0.02fF
C48290 INVX1_LOC_89/A INVX1_LOC_6/A 0.49fF
C48291 NOR2X1_LOC_348/B NAND2X1_LOC_418/a_36_24# 0.00fF
C48292 INVX1_LOC_292/A INVX1_LOC_19/A 0.07fF
C48293 NAND2X1_LOC_337/B NOR2X1_LOC_831/Y 0.34fF
C48294 NAND2X1_LOC_374/Y INVX1_LOC_46/A 0.10fF
C48295 NOR2X1_LOC_368/a_36_216# NOR2X1_LOC_76/A 0.01fF
C48296 NOR2X1_LOC_824/Y INVX1_LOC_22/A 0.40fF
C48297 NAND2X1_LOC_339/a_36_24# NOR2X1_LOC_331/B 0.01fF
C48298 INVX1_LOC_49/A INVX1_LOC_291/A 0.02fF
C48299 NOR2X1_LOC_703/A NOR2X1_LOC_337/A 0.14fF
C48300 NAND2X1_LOC_833/Y INVX1_LOC_185/A 0.02fF
C48301 NOR2X1_LOC_716/B NOR2X1_LOC_118/a_36_216# 0.01fF
C48302 INVX1_LOC_22/A INVX1_LOC_76/A 0.90fF
C48303 NOR2X1_LOC_385/Y INPUT_0 0.03fF
C48304 NOR2X1_LOC_340/Y NOR2X1_LOC_61/Y 0.03fF
C48305 INVX1_LOC_172/Y VDD 0.19fF
C48306 NOR2X1_LOC_646/A INVX1_LOC_2/Y 0.21fF
C48307 INVX1_LOC_14/A INVX1_LOC_251/A 0.07fF
C48308 NOR2X1_LOC_318/B NOR2X1_LOC_355/a_36_216# 0.00fF
C48309 NAND2X1_LOC_859/Y NAND2X1_LOC_244/A 0.07fF
C48310 NOR2X1_LOC_392/Y INVX1_LOC_23/A 0.07fF
C48311 INVX1_LOC_35/A INVX1_LOC_25/A 0.02fF
C48312 NAND2X1_LOC_842/B INVX1_LOC_91/A 0.13fF
C48313 INVX1_LOC_95/Y NOR2X1_LOC_71/Y 0.10fF
C48314 NAND2X1_LOC_36/A INPUT_7 0.44fF
C48315 INVX1_LOC_58/A INVX1_LOC_64/A 10.09fF
C48316 NAND2X1_LOC_484/a_36_24# INVX1_LOC_92/A 0.01fF
C48317 INVX1_LOC_90/A INVX1_LOC_93/Y 0.07fF
C48318 NOR2X1_LOC_218/A INVX1_LOC_15/A 0.04fF
C48319 INVX1_LOC_69/Y NOR2X1_LOC_336/a_36_216# 0.01fF
C48320 NOR2X1_LOC_447/Y INVX1_LOC_84/A 0.03fF
C48321 INVX1_LOC_34/A NOR2X1_LOC_831/B 0.03fF
C48322 NAND2X1_LOC_466/A NOR2X1_LOC_435/A 0.01fF
C48323 INVX1_LOC_24/A NAND2X1_LOC_768/Y 0.03fF
C48324 INVX1_LOC_225/A NOR2X1_LOC_155/A 0.07fF
C48325 INVX1_LOC_154/A INVX1_LOC_156/A 0.05fF
C48326 NOR2X1_LOC_389/B INVX1_LOC_93/Y 0.05fF
C48327 NAND2X1_LOC_123/Y NOR2X1_LOC_269/Y 0.00fF
C48328 INVX1_LOC_62/A INVX1_LOC_176/A 0.04fF
C48329 INVX1_LOC_200/A NAND2X1_LOC_444/B 0.01fF
C48330 NOR2X1_LOC_272/Y INVX1_LOC_50/A 0.03fF
C48331 INVX1_LOC_2/A INVX1_LOC_291/A 0.07fF
C48332 NOR2X1_LOC_332/A D_INPUT_3 0.14fF
C48333 NAND2X1_LOC_342/Y NOR2X1_LOC_743/Y 0.02fF
C48334 INVX1_LOC_2/A NAND2X1_LOC_802/Y 0.07fF
C48335 NOR2X1_LOC_826/Y INVX1_LOC_5/A 0.02fF
C48336 INVX1_LOC_223/Y INVX1_LOC_23/A 0.68fF
C48337 NOR2X1_LOC_246/A NAND2X1_LOC_287/B 1.21fF
C48338 INVX1_LOC_10/A NAND2X1_LOC_472/Y 0.29fF
C48339 NOR2X1_LOC_226/A INVX1_LOC_291/A 0.10fF
C48340 INVX1_LOC_33/A INVX1_LOC_63/A 0.04fF
C48341 NOR2X1_LOC_209/Y NOR2X1_LOC_155/A 0.03fF
C48342 INVX1_LOC_308/A NOR2X1_LOC_652/Y 0.01fF
C48343 NOR2X1_LOC_759/Y INVX1_LOC_109/A 0.00fF
C48344 NAND2X1_LOC_756/a_36_24# NOR2X1_LOC_363/Y 0.00fF
C48345 NOR2X1_LOC_315/Y NAND2X1_LOC_572/B 0.08fF
C48346 INVX1_LOC_85/Y VDD 0.44fF
C48347 NOR2X1_LOC_468/Y NOR2X1_LOC_383/B 0.03fF
C48348 INVX1_LOC_135/A NOR2X1_LOC_813/Y 0.10fF
C48349 NOR2X1_LOC_735/Y INVX1_LOC_76/A -0.02fF
C48350 INVX1_LOC_64/A NAND2X1_LOC_190/a_36_24# 0.00fF
C48351 INVX1_LOC_135/A NOR2X1_LOC_152/A 0.01fF
C48352 NAND2X1_LOC_190/Y NOR2X1_LOC_383/B 0.17fF
C48353 NOR2X1_LOC_689/Y NAND2X1_LOC_724/A 0.01fF
C48354 INVX1_LOC_233/A NAND2X1_LOC_170/a_36_24# 0.00fF
C48355 INVX1_LOC_90/A NAND2X1_LOC_721/A 5.65fF
C48356 NAND2X1_LOC_149/Y INVX1_LOC_259/Y 0.07fF
C48357 NOR2X1_LOC_83/Y NAND2X1_LOC_642/Y 0.06fF
C48358 INVX1_LOC_235/Y NOR2X1_LOC_660/Y 0.14fF
C48359 INVX1_LOC_135/A INVX1_LOC_280/A 1.11fF
C48360 INVX1_LOC_209/Y INVX1_LOC_12/A 0.07fF
C48361 D_INPUT_1 NOR2X1_LOC_187/Y 0.02fF
C48362 INVX1_LOC_236/Y NAND2X1_LOC_175/Y 0.04fF
C48363 NAND2X1_LOC_228/a_36_24# INVX1_LOC_117/Y 0.00fF
C48364 INVX1_LOC_266/Y NOR2X1_LOC_631/A 0.30fF
C48365 NAND2X1_LOC_855/Y VDD 0.03fF
C48366 NOR2X1_LOC_646/A NOR2X1_LOC_608/Y 0.13fF
C48367 NAND2X1_LOC_139/A INVX1_LOC_29/A 0.03fF
C48368 NOR2X1_LOC_366/B NOR2X1_LOC_473/a_36_216# 0.00fF
C48369 INVX1_LOC_36/Y NOR2X1_LOC_196/Y 0.00fF
C48370 NAND2X1_LOC_629/Y INVX1_LOC_186/Y 0.01fF
C48371 NAND2X1_LOC_860/A NOR2X1_LOC_361/B 0.10fF
C48372 INVX1_LOC_299/A INVX1_LOC_58/Y 0.08fF
C48373 NAND2X1_LOC_538/Y INVX1_LOC_53/A 0.07fF
C48374 INVX1_LOC_35/A INVX1_LOC_1/A 0.28fF
C48375 NAND2X1_LOC_861/Y INVX1_LOC_118/A 0.07fF
C48376 NOR2X1_LOC_560/A INVX1_LOC_280/A 0.02fF
C48377 INVX1_LOC_10/A NAND2X1_LOC_434/Y 0.01fF
C48378 NOR2X1_LOC_558/A NOR2X1_LOC_74/A 0.01fF
C48379 INVX1_LOC_41/A NOR2X1_LOC_461/Y 0.01fF
C48380 INVX1_LOC_279/A INVX1_LOC_179/A 0.01fF
C48381 NAND2X1_LOC_725/A NAND2X1_LOC_724/A 0.10fF
C48382 INVX1_LOC_41/A NOR2X1_LOC_640/B 0.06fF
C48383 INVX1_LOC_6/A NAND2X1_LOC_244/A 0.01fF
C48384 NAND2X1_LOC_291/a_36_24# NAND2X1_LOC_96/A 0.00fF
C48385 NAND2X1_LOC_794/B NAND2X1_LOC_714/B 0.01fF
C48386 NAND2X1_LOC_655/a_36_24# INVX1_LOC_49/Y 0.00fF
C48387 INVX1_LOC_40/A INVX1_LOC_63/A 0.39fF
C48388 INVX1_LOC_89/A NOR2X1_LOC_79/A 0.05fF
C48389 NOR2X1_LOC_558/A NOR2X1_LOC_9/Y 0.02fF
C48390 NOR2X1_LOC_346/a_36_216# INVX1_LOC_280/A 0.01fF
C48391 NOR2X1_LOC_356/A NOR2X1_LOC_729/A 0.07fF
C48392 NOR2X1_LOC_15/Y NOR2X1_LOC_291/Y 0.18fF
C48393 NOR2X1_LOC_303/Y INVX1_LOC_4/Y 0.21fF
C48394 INVX1_LOC_50/A NOR2X1_LOC_761/Y 0.05fF
C48395 INVX1_LOC_55/Y NAND2X1_LOC_260/a_36_24# 0.00fF
C48396 NOR2X1_LOC_742/A INVX1_LOC_38/A 0.07fF
C48397 INVX1_LOC_24/A NOR2X1_LOC_36/A 2.58fF
C48398 NAND2X1_LOC_731/Y NAND2X1_LOC_175/Y 0.01fF
C48399 INVX1_LOC_226/Y NAND2X1_LOC_773/B 0.40fF
C48400 NAND2X1_LOC_648/A NAND2X1_LOC_802/Y 0.02fF
C48401 NOR2X1_LOC_548/B NOR2X1_LOC_107/a_36_216# 0.03fF
C48402 INVX1_LOC_31/A NOR2X1_LOC_392/Y 0.15fF
C48403 INVX1_LOC_208/A INVX1_LOC_272/A 0.02fF
C48404 INVX1_LOC_50/A NAND2X1_LOC_364/A 0.07fF
C48405 INVX1_LOC_33/A NAND2X1_LOC_452/Y 0.02fF
C48406 INVX1_LOC_314/Y INVX1_LOC_26/A 0.09fF
C48407 NOR2X1_LOC_815/Y INVX1_LOC_78/A 0.02fF
C48408 NAND2X1_LOC_715/B NOR2X1_LOC_45/Y 0.01fF
C48409 NOR2X1_LOC_15/Y NAND2X1_LOC_347/B 0.07fF
C48410 NOR2X1_LOC_391/B INVX1_LOC_280/A 0.01fF
C48411 INVX1_LOC_17/A NAND2X1_LOC_816/a_36_24# 0.00fF
C48412 INVX1_LOC_16/A NAND2X1_LOC_74/B 0.11fF
C48413 INVX1_LOC_113/Y NOR2X1_LOC_631/Y 0.00fF
C48414 NAND2X1_LOC_112/Y INVX1_LOC_29/A 0.03fF
C48415 NOR2X1_LOC_596/A NOR2X1_LOC_383/B 0.07fF
C48416 NOR2X1_LOC_574/A INVX1_LOC_21/Y 0.01fF
C48417 NOR2X1_LOC_631/B NOR2X1_LOC_562/A 0.03fF
C48418 NOR2X1_LOC_131/A INVX1_LOC_15/A 0.02fF
C48419 INVX1_LOC_35/A NOR2X1_LOC_384/Y 0.07fF
C48420 INVX1_LOC_131/A NOR2X1_LOC_831/B 0.04fF
C48421 INVX1_LOC_232/Y INVX1_LOC_32/A 0.08fF
C48422 NAND2X1_LOC_654/a_36_24# INVX1_LOC_15/A 0.01fF
C48423 INVX1_LOC_103/A NOR2X1_LOC_122/A 0.01fF
C48424 NOR2X1_LOC_716/B INVX1_LOC_181/A 0.00fF
C48425 NOR2X1_LOC_318/B INVX1_LOC_38/A 0.05fF
C48426 INVX1_LOC_54/Y INVX1_LOC_4/Y 0.04fF
C48427 NOR2X1_LOC_272/Y INVX1_LOC_61/Y 0.10fF
C48428 NAND2X1_LOC_735/B INVX1_LOC_42/A 0.03fF
C48429 NOR2X1_LOC_45/B NOR2X1_LOC_331/B 0.20fF
C48430 NOR2X1_LOC_91/A NAND2X1_LOC_736/Y 0.03fF
C48431 INVX1_LOC_93/Y NOR2X1_LOC_561/A 0.03fF
C48432 NAND2X1_LOC_283/a_36_24# INVX1_LOC_270/A 0.00fF
C48433 NOR2X1_LOC_634/a_36_216# NOR2X1_LOC_383/B 0.02fF
C48434 INPUT_0 NOR2X1_LOC_831/B 0.03fF
C48435 NAND2X1_LOC_198/B NOR2X1_LOC_109/a_36_216# 0.01fF
C48436 INVX1_LOC_89/A INVX1_LOC_301/A 0.02fF
C48437 NOR2X1_LOC_160/B NOR2X1_LOC_271/B 0.01fF
C48438 INVX1_LOC_24/Y NAND2X1_LOC_114/B 0.24fF
C48439 INVX1_LOC_226/Y NOR2X1_LOC_393/Y 0.01fF
C48440 INVX1_LOC_103/A INVX1_LOC_161/Y 0.03fF
C48441 INPUT_0 NOR2X1_LOC_179/a_36_216# 0.00fF
C48442 NAND2X1_LOC_796/B NAND2X1_LOC_721/B 0.18fF
C48443 NOR2X1_LOC_266/B NAND2X1_LOC_262/a_36_24# 0.02fF
C48444 NOR2X1_LOC_68/A INVX1_LOC_38/Y 0.01fF
C48445 NOR2X1_LOC_497/a_36_216# NOR2X1_LOC_690/A 0.01fF
C48446 NOR2X1_LOC_332/A NAND2X1_LOC_233/a_36_24# 0.00fF
C48447 NOR2X1_LOC_598/B NOR2X1_LOC_374/A 0.12fF
C48448 NOR2X1_LOC_455/Y NOR2X1_LOC_577/Y -0.02fF
C48449 NAND2X1_LOC_45/Y NAND2X1_LOC_291/B 0.01fF
C48450 INVX1_LOC_247/A NOR2X1_LOC_331/B 0.42fF
C48451 NOR2X1_LOC_470/B NOR2X1_LOC_478/A 0.02fF
C48452 NAND2X1_LOC_833/Y NOR2X1_LOC_754/Y 0.00fF
C48453 INVX1_LOC_90/A NOR2X1_LOC_669/A 0.01fF
C48454 NAND2X1_LOC_729/B INVX1_LOC_185/A 0.00fF
C48455 INVX1_LOC_230/Y INVX1_LOC_11/A 0.07fF
C48456 NAND2X1_LOC_9/Y NAND2X1_LOC_276/Y 0.04fF
C48457 INVX1_LOC_28/A NAND2X1_LOC_74/B 0.10fF
C48458 INVX1_LOC_27/A NOR2X1_LOC_360/Y 0.07fF
C48459 NOR2X1_LOC_454/Y NAND2X1_LOC_16/Y 0.01fF
C48460 NOR2X1_LOC_802/A NOR2X1_LOC_809/A 0.20fF
C48461 NAND2X1_LOC_360/B NAND2X1_LOC_99/A 0.05fF
C48462 NAND2X1_LOC_785/A INVX1_LOC_50/A 0.05fF
C48463 NOR2X1_LOC_160/B INVX1_LOC_150/Y 0.07fF
C48464 INVX1_LOC_292/A INVX1_LOC_161/Y 0.05fF
C48465 NOR2X1_LOC_78/A NOR2X1_LOC_634/A 0.01fF
C48466 NOR2X1_LOC_45/B NOR2X1_LOC_592/B 0.03fF
C48467 NOR2X1_LOC_142/Y NOR2X1_LOC_678/A 0.04fF
C48468 INVX1_LOC_1/Y NAND2X1_LOC_223/A 0.84fF
C48469 NOR2X1_LOC_146/a_36_216# INVX1_LOC_91/A 0.00fF
C48470 NOR2X1_LOC_598/B NOR2X1_LOC_288/A 0.03fF
C48471 NAND2X1_LOC_721/A NAND2X1_LOC_849/B 0.02fF
C48472 NOR2X1_LOC_826/Y NAND2X1_LOC_562/B 0.01fF
C48473 NOR2X1_LOC_455/Y NOR2X1_LOC_348/B 0.05fF
C48474 INVX1_LOC_104/A NOR2X1_LOC_717/A 0.08fF
C48475 NOR2X1_LOC_220/A NOR2X1_LOC_383/B 0.01fF
C48476 NOR2X1_LOC_500/A NOR2X1_LOC_790/A 0.04fF
C48477 NOR2X1_LOC_91/A INVX1_LOC_25/Y 0.19fF
C48478 INPUT_5 INVX1_LOC_78/A 0.03fF
C48479 NOR2X1_LOC_690/A INVX1_LOC_5/A 0.00fF
C48480 NOR2X1_LOC_689/Y NAND2X1_LOC_852/Y 0.05fF
C48481 NAND2X1_LOC_463/B INVX1_LOC_167/A 0.01fF
C48482 NOR2X1_LOC_689/A NAND2X1_LOC_863/B 0.02fF
C48483 NOR2X1_LOC_689/a_36_216# NAND2X1_LOC_853/Y 0.03fF
C48484 INVX1_LOC_58/A NAND2X1_LOC_850/Y 0.74fF
C48485 INVX1_LOC_91/A INVX1_LOC_119/Y 0.02fF
C48486 INVX1_LOC_22/A NOR2X1_LOC_447/A 0.26fF
C48487 NOR2X1_LOC_598/B NOR2X1_LOC_209/Y 0.15fF
C48488 NOR2X1_LOC_413/Y INVX1_LOC_5/A 0.01fF
C48489 NOR2X1_LOC_784/Y NAND2X1_LOC_146/a_36_24# 0.00fF
C48490 INVX1_LOC_13/Y NAND2X1_LOC_569/A 0.02fF
C48491 VDD NOR2X1_LOC_487/Y 0.12fF
C48492 D_INPUT_1 INVX1_LOC_43/A 0.03fF
C48493 NOR2X1_LOC_276/a_36_216# INVX1_LOC_103/A 0.00fF
C48494 NOR2X1_LOC_194/Y INVX1_LOC_5/A 0.01fF
C48495 NAND2X1_LOC_763/B INVX1_LOC_174/A 0.64fF
C48496 NOR2X1_LOC_557/Y NAND2X1_LOC_474/Y 0.11fF
C48497 NOR2X1_LOC_824/A INVX1_LOC_207/A 0.03fF
C48498 INVX1_LOC_88/A NOR2X1_LOC_363/a_36_216# 0.00fF
C48499 NOR2X1_LOC_690/A INVX1_LOC_178/A 0.10fF
C48500 INVX1_LOC_272/Y INVX1_LOC_24/A 0.11fF
C48501 INVX1_LOC_25/Y INVX1_LOC_23/A 0.10fF
C48502 NOR2X1_LOC_94/Y INVX1_LOC_280/A 0.04fF
C48503 NOR2X1_LOC_548/Y NOR2X1_LOC_383/B 0.00fF
C48504 VDD NOR2X1_LOC_461/A -0.00fF
C48505 NOR2X1_LOC_312/Y NAND2X1_LOC_175/Y 0.01fF
C48506 NAND2X1_LOC_647/a_36_24# INVX1_LOC_46/A 0.00fF
C48507 NAND2X1_LOC_738/B NAND2X1_LOC_863/B 6.26fF
C48508 NAND2X1_LOC_573/A NAND2X1_LOC_286/B 0.06fF
C48509 INVX1_LOC_2/Y NOR2X1_LOC_608/Y 0.00fF
C48510 INVX1_LOC_25/A NOR2X1_LOC_121/A 0.63fF
C48511 NOR2X1_LOC_210/a_36_216# INVX1_LOC_113/Y 0.00fF
C48512 NOR2X1_LOC_413/Y INVX1_LOC_178/A 0.10fF
C48513 NAND2X1_LOC_53/Y INVX1_LOC_24/A 0.31fF
C48514 INVX1_LOC_299/A NOR2X1_LOC_537/A 0.01fF
C48515 INVX1_LOC_207/A INVX1_LOC_237/A 0.07fF
C48516 INVX1_LOC_10/A NOR2X1_LOC_481/a_36_216# 0.01fF
C48517 NAND2X1_LOC_349/B INVX1_LOC_23/A 0.17fF
C48518 INVX1_LOC_90/A INVX1_LOC_87/A 0.05fF
C48519 INVX1_LOC_309/A INVX1_LOC_284/A 0.16fF
C48520 NOR2X1_LOC_86/Y INVX1_LOC_31/A 0.01fF
C48521 INVX1_LOC_263/A NOR2X1_LOC_717/A 0.18fF
C48522 INVX1_LOC_135/A NAND2X1_LOC_416/a_36_24# 0.00fF
C48523 NAND2X1_LOC_721/A NAND2X1_LOC_848/Y 0.09fF
C48524 NAND2X1_LOC_472/Y INVX1_LOC_307/A 0.96fF
C48525 NOR2X1_LOC_389/B INVX1_LOC_87/A 0.08fF
C48526 NOR2X1_LOC_455/Y INVX1_LOC_22/A 0.04fF
C48527 INVX1_LOC_120/A INVX1_LOC_26/Y 0.00fF
C48528 INVX1_LOC_88/A INVX1_LOC_155/A 0.01fF
C48529 NOR2X1_LOC_78/A INVX1_LOC_29/A 0.10fF
C48530 NOR2X1_LOC_68/A INVX1_LOC_286/Y 0.10fF
C48531 NOR2X1_LOC_538/B NOR2X1_LOC_716/B 0.00fF
C48532 NOR2X1_LOC_860/Y INVX1_LOC_9/A 0.04fF
C48533 NOR2X1_LOC_542/B INVX1_LOC_19/A 0.03fF
C48534 INVX1_LOC_37/A INVX1_LOC_285/A 0.07fF
C48535 INVX1_LOC_159/Y INVX1_LOC_109/Y 0.02fF
C48536 NOR2X1_LOC_58/Y NOR2X1_LOC_60/Y 0.07fF
C48537 INVX1_LOC_91/A INVX1_LOC_284/A 0.07fF
C48538 NAND2X1_LOC_391/Y NAND2X1_LOC_338/B 0.07fF
C48539 INVX1_LOC_38/A INVX1_LOC_117/Y 0.03fF
C48540 NAND2X1_LOC_859/Y NOR2X1_LOC_392/Y 0.01fF
C48541 NAND2X1_LOC_724/A NAND2X1_LOC_308/Y 0.02fF
C48542 INVX1_LOC_37/A INVX1_LOC_265/Y 0.12fF
C48543 NAND2X1_LOC_860/A NAND2X1_LOC_573/A 0.04fF
C48544 NOR2X1_LOC_391/Y INVX1_LOC_32/A 0.01fF
C48545 NAND2X1_LOC_93/B INVX1_LOC_193/A 0.03fF
C48546 INVX1_LOC_161/Y INVX1_LOC_67/A 0.05fF
C48547 NOR2X1_LOC_533/Y NAND2X1_LOC_811/Y 0.09fF
C48548 NOR2X1_LOC_658/Y NOR2X1_LOC_215/Y 0.03fF
C48549 NAND2X1_LOC_725/Y NOR2X1_LOC_380/A 0.81fF
C48550 INVX1_LOC_291/A INVX1_LOC_118/A 0.10fF
C48551 INVX1_LOC_143/Y INVX1_LOC_19/A 0.03fF
C48552 INVX1_LOC_186/Y INVX1_LOC_76/A 0.13fF
C48553 INVX1_LOC_37/A NOR2X1_LOC_814/A 0.12fF
C48554 INVX1_LOC_161/A NOR2X1_LOC_387/Y 0.06fF
C48555 INVX1_LOC_93/A NAND2X1_LOC_862/A 0.03fF
C48556 NOR2X1_LOC_231/A NOR2X1_LOC_814/A 0.02fF
C48557 NOR2X1_LOC_665/A NOR2X1_LOC_665/Y 0.03fF
C48558 INVX1_LOC_287/A NOR2X1_LOC_708/Y 0.02fF
C48559 INVX1_LOC_31/A NOR2X1_LOC_554/a_36_216# 0.01fF
C48560 VDD NAND2X1_LOC_782/B 0.01fF
C48561 NOR2X1_LOC_82/A NOR2X1_LOC_392/B 0.03fF
C48562 INVX1_LOC_193/A NAND2X1_LOC_425/Y 0.01fF
C48563 INVX1_LOC_24/Y NOR2X1_LOC_168/B 0.03fF
C48564 NOR2X1_LOC_489/A INVX1_LOC_92/A 0.17fF
C48565 INVX1_LOC_41/A NAND2X1_LOC_114/B 0.15fF
C48566 NOR2X1_LOC_51/a_36_216# D_INPUT_5 0.00fF
C48567 NAND2X1_LOC_169/a_36_24# INVX1_LOC_30/A 0.00fF
C48568 NOR2X1_LOC_160/B NAND2X1_LOC_494/a_36_24# 0.00fF
C48569 NAND2X1_LOC_733/Y INVX1_LOC_209/Y 0.05fF
C48570 NOR2X1_LOC_68/A INVX1_LOC_159/A 0.03fF
C48571 INVX1_LOC_157/Y NOR2X1_LOC_364/A 0.03fF
C48572 NOR2X1_LOC_106/A INVX1_LOC_53/A 0.04fF
C48573 NOR2X1_LOC_35/Y NAND2X1_LOC_74/B 0.10fF
C48574 NOR2X1_LOC_35/Y NAND2X1_LOC_207/Y 0.16fF
C48575 INVX1_LOC_13/A INVX1_LOC_50/Y 0.07fF
C48576 NOR2X1_LOC_860/B INVX1_LOC_110/A 0.02fF
C48577 NAND2X1_LOC_211/Y INVX1_LOC_272/A 0.03fF
C48578 NOR2X1_LOC_274/Y NOR2X1_LOC_274/B 0.00fF
C48579 NAND2X1_LOC_303/Y NOR2X1_LOC_773/Y 0.02fF
C48580 NOR2X1_LOC_209/Y NOR2X1_LOC_742/a_36_216# 0.00fF
C48581 INVX1_LOC_230/Y NOR2X1_LOC_52/B 0.09fF
C48582 NOR2X1_LOC_590/A NOR2X1_LOC_799/a_36_216# 0.00fF
C48583 NAND2X1_LOC_784/A NOR2X1_LOC_329/B 0.02fF
C48584 NOR2X1_LOC_238/a_36_216# NOR2X1_LOC_238/Y 0.00fF
C48585 NOR2X1_LOC_54/a_36_216# INVX1_LOC_3/A 0.02fF
C48586 NOR2X1_LOC_75/Y NOR2X1_LOC_432/Y 0.01fF
C48587 NOR2X1_LOC_133/a_36_216# NAND2X1_LOC_74/B 0.00fF
C48588 NOR2X1_LOC_78/B NOR2X1_LOC_250/A 0.04fF
C48589 NAND2X1_LOC_755/a_36_24# INVX1_LOC_31/A 0.00fF
C48590 NOR2X1_LOC_607/A INVX1_LOC_77/A 0.01fF
C48591 INVX1_LOC_75/A INVX1_LOC_23/A 0.23fF
C48592 INVX1_LOC_14/Y INVX1_LOC_42/A 0.05fF
C48593 INVX1_LOC_12/A NAND2X1_LOC_472/Y 0.07fF
C48594 NAND2X1_LOC_206/a_36_24# NOR2X1_LOC_844/A 0.00fF
C48595 INVX1_LOC_45/A NOR2X1_LOC_180/Y 0.03fF
C48596 NOR2X1_LOC_843/B NAND2X1_LOC_251/a_36_24# 0.03fF
C48597 INVX1_LOC_232/Y INPUT_3 0.10fF
C48598 NOR2X1_LOC_381/Y INVX1_LOC_13/A 0.09fF
C48599 INVX1_LOC_312/Y NAND2X1_LOC_477/A 0.10fF
C48600 NOR2X1_LOC_45/B NOR2X1_LOC_449/A 0.03fF
C48601 NOR2X1_LOC_557/A INVX1_LOC_26/A 0.25fF
C48602 NOR2X1_LOC_92/Y NAND2X1_LOC_656/Y 0.07fF
C48603 INVX1_LOC_303/A INVX1_LOC_8/Y 0.05fF
C48604 INVX1_LOC_83/A NAND2X1_LOC_218/A 0.04fF
C48605 NOR2X1_LOC_790/B INPUT_0 0.07fF
C48606 INVX1_LOC_11/A GATE_479 0.03fF
C48607 NOR2X1_LOC_540/B INVX1_LOC_271/Y 0.05fF
C48608 NOR2X1_LOC_56/Y NAND2X1_LOC_454/Y -0.02fF
C48609 INVX1_LOC_294/Y INVX1_LOC_181/Y 0.54fF
C48610 INVX1_LOC_78/A NAND2X1_LOC_212/Y 0.00fF
C48611 NAND2X1_LOC_483/Y NAND2X1_LOC_837/Y 0.11fF
C48612 NOR2X1_LOC_815/Y NOR2X1_LOC_152/Y 0.01fF
C48613 INVX1_LOC_299/A NOR2X1_LOC_326/Y 0.00fF
C48614 INVX1_LOC_18/A NAND2X1_LOC_629/Y 0.00fF
C48615 INVX1_LOC_254/Y NAND2X1_LOC_361/Y 0.01fF
C48616 INVX1_LOC_35/A NOR2X1_LOC_188/A 0.04fF
C48617 NAND2X1_LOC_636/a_36_24# INVX1_LOC_38/A 0.00fF
C48618 NOR2X1_LOC_532/a_36_216# INVX1_LOC_179/Y 0.03fF
C48619 INVX1_LOC_31/A INVX1_LOC_25/Y 0.04fF
C48620 INVX1_LOC_206/A NOR2X1_LOC_360/Y 0.10fF
C48621 INVX1_LOC_83/A NAND2X1_LOC_538/Y 0.02fF
C48622 INVX1_LOC_35/A NOR2X1_LOC_548/B 0.01fF
C48623 INVX1_LOC_124/A NOR2X1_LOC_607/A 0.01fF
C48624 NOR2X1_LOC_335/A NOR2X1_LOC_142/Y 0.01fF
C48625 INVX1_LOC_243/A INVX1_LOC_18/A 0.02fF
C48626 NOR2X1_LOC_269/Y INVX1_LOC_271/A 0.23fF
C48627 NAND2X1_LOC_741/Y NOR2X1_LOC_380/Y 0.02fF
C48628 INVX1_LOC_289/Y INVX1_LOC_90/A 0.01fF
C48629 INVX1_LOC_57/A NAND2X1_LOC_655/A 0.07fF
C48630 INVX1_LOC_50/A NOR2X1_LOC_405/A 0.03fF
C48631 VDD NAND2X1_LOC_454/Y 1.44fF
C48632 INVX1_LOC_18/A INVX1_LOC_179/Y 1.31fF
C48633 INVX1_LOC_14/Y INVX1_LOC_78/A 0.45fF
C48634 NOR2X1_LOC_172/Y NAND2X1_LOC_332/Y 0.09fF
C48635 NAND2X1_LOC_169/Y INPUT_0 0.02fF
C48636 NAND2X1_LOC_326/A NOR2X1_LOC_329/B 0.68fF
C48637 NAND2X1_LOC_200/B NOR2X1_LOC_360/Y 0.08fF
C48638 NOR2X1_LOC_860/Y NOR2X1_LOC_861/Y 0.25fF
C48639 NOR2X1_LOC_172/a_36_216# INVX1_LOC_71/A 0.00fF
C48640 NOR2X1_LOC_589/A INVX1_LOC_30/A 0.10fF
C48641 INVX1_LOC_136/A INVX1_LOC_16/A 0.44fF
C48642 NOR2X1_LOC_716/B NOR2X1_LOC_315/Y 0.50fF
C48643 INVX1_LOC_95/Y NAND2X1_LOC_205/A 0.10fF
C48644 NOR2X1_LOC_82/A INVX1_LOC_90/A 0.07fF
C48645 NOR2X1_LOC_690/A NAND2X1_LOC_562/B 0.01fF
C48646 NOR2X1_LOC_91/A NAND2X1_LOC_453/A 0.23fF
C48647 NOR2X1_LOC_627/a_36_216# INVX1_LOC_113/Y 0.00fF
C48648 INVX1_LOC_34/A NAND2X1_LOC_357/B 0.90fF
C48649 INVX1_LOC_35/A NOR2X1_LOC_43/Y 0.06fF
C48650 NAND2X1_LOC_633/Y INVX1_LOC_181/A 0.02fF
C48651 NOR2X1_LOC_413/Y NAND2X1_LOC_562/B 0.01fF
C48652 NOR2X1_LOC_495/Y NAND2X1_LOC_483/a_36_24# 0.01fF
C48653 INVX1_LOC_24/A NOR2X1_LOC_500/Y 0.07fF
C48654 NAND2X1_LOC_624/B NAND2X1_LOC_623/B 0.08fF
C48655 INVX1_LOC_226/Y INVX1_LOC_24/A 0.49fF
C48656 NOR2X1_LOC_67/Y NAND2X1_LOC_85/Y 0.12fF
C48657 NOR2X1_LOC_631/A INVX1_LOC_19/A 0.06fF
C48658 INVX1_LOC_41/A NOR2X1_LOC_168/B 0.03fF
C48659 NOR2X1_LOC_331/B NOR2X1_LOC_465/Y 0.01fF
C48660 NAND2X1_LOC_99/a_36_24# NAND2X1_LOC_338/B 0.00fF
C48661 INVX1_LOC_309/A NOR2X1_LOC_384/A 0.01fF
C48662 NAND2X1_LOC_79/Y INVX1_LOC_232/A 0.00fF
C48663 NOR2X1_LOC_561/Y INVX1_LOC_18/A 0.34fF
C48664 INVX1_LOC_290/A NOR2X1_LOC_759/Y 0.01fF
C48665 INVX1_LOC_23/A NAND2X1_LOC_453/A 0.07fF
C48666 NAND2X1_LOC_787/A INVX1_LOC_20/A 0.03fF
C48667 INVX1_LOC_171/A INVX1_LOC_30/A 0.09fF
C48668 NAND2X1_LOC_390/A INVX1_LOC_41/Y 0.02fF
C48669 NOR2X1_LOC_720/A INVX1_LOC_117/A 0.00fF
C48670 INVX1_LOC_34/A NAND2X1_LOC_549/B 0.01fF
C48671 NOR2X1_LOC_222/a_36_216# INVX1_LOC_81/A 0.00fF
C48672 NOR2X1_LOC_708/A INVX1_LOC_213/A 0.00fF
C48673 INVX1_LOC_36/A INVX1_LOC_89/A 0.06fF
C48674 NAND2X1_LOC_363/B INVX1_LOC_20/A 0.03fF
C48675 NOR2X1_LOC_82/A NAND2X1_LOC_348/A 0.20fF
C48676 NOR2X1_LOC_67/A NOR2X1_LOC_121/Y 0.04fF
C48677 INVX1_LOC_202/A INVX1_LOC_290/A 0.06fF
C48678 INVX1_LOC_106/Y INVX1_LOC_63/A 0.00fF
C48679 NOR2X1_LOC_672/Y INVX1_LOC_316/Y 0.12fF
C48680 INVX1_LOC_295/A NAND2X1_LOC_387/B 0.05fF
C48681 INVX1_LOC_45/Y INVX1_LOC_279/A 0.04fF
C48682 INVX1_LOC_13/A NOR2X1_LOC_559/B 0.03fF
C48683 INVX1_LOC_203/A INVX1_LOC_284/A 0.10fF
C48684 NOR2X1_LOC_124/A NOR2X1_LOC_293/a_36_216# 0.00fF
C48685 INVX1_LOC_27/A NOR2X1_LOC_269/Y 0.07fF
C48686 NOR2X1_LOC_520/A NAND2X1_LOC_116/A 0.01fF
C48687 NAND2X1_LOC_352/B INVX1_LOC_131/A 0.13fF
C48688 INVX1_LOC_12/A NAND2X1_LOC_773/B 0.07fF
C48689 NAND2X1_LOC_231/Y NAND2X1_LOC_357/B 0.10fF
C48690 INVX1_LOC_24/A INVX1_LOC_10/A 0.04fF
C48691 NOR2X1_LOC_637/Y NOR2X1_LOC_561/Y 0.04fF
C48692 NOR2X1_LOC_483/B NOR2X1_LOC_742/A 0.03fF
C48693 NAND2X1_LOC_182/A INVX1_LOC_256/Y 0.36fF
C48694 NOR2X1_LOC_334/Y INVX1_LOC_92/A 0.07fF
C48695 INVX1_LOC_237/Y INVX1_LOC_22/A 0.09fF
C48696 NOR2X1_LOC_632/Y INVX1_LOC_49/A 0.03fF
C48697 INVX1_LOC_33/A INVX1_LOC_1/Y 0.07fF
C48698 INVX1_LOC_314/Y INVX1_LOC_164/A 0.01fF
C48699 INVX1_LOC_17/A NOR2X1_LOC_734/a_36_216# 0.00fF
C48700 INVX1_LOC_109/A NAND2X1_LOC_74/B 0.07fF
C48701 INVX1_LOC_31/A INVX1_LOC_75/A 0.07fF
C48702 INVX1_LOC_136/A INVX1_LOC_28/A 0.17fF
C48703 INVX1_LOC_90/A NAND2X1_LOC_153/a_36_24# 0.00fF
C48704 NOR2X1_LOC_791/Y INVX1_LOC_20/A 0.02fF
C48705 NAND2X1_LOC_341/A NOR2X1_LOC_52/B 0.00fF
C48706 INVX1_LOC_286/Y NOR2X1_LOC_2/Y 0.01fF
C48707 INVX1_LOC_46/A NOR2X1_LOC_81/Y 0.07fF
C48708 NAND2X1_LOC_538/Y NOR2X1_LOC_311/Y 0.10fF
C48709 INVX1_LOC_256/A NOR2X1_LOC_355/B 0.38fF
C48710 INVX1_LOC_13/A NOR2X1_LOC_6/B 0.13fF
C48711 NOR2X1_LOC_290/Y INVX1_LOC_25/Y 0.03fF
C48712 INVX1_LOC_167/A INVX1_LOC_42/A 0.01fF
C48713 D_INPUT_0 NOR2X1_LOC_520/B 0.30fF
C48714 INVX1_LOC_24/A NOR2X1_LOC_302/Y 0.17fF
C48715 NAND2X1_LOC_342/Y INVX1_LOC_53/Y 0.00fF
C48716 INVX1_LOC_45/Y INVX1_LOC_182/Y 0.04fF
C48717 INVX1_LOC_2/A NOR2X1_LOC_632/Y 0.04fF
C48718 INVX1_LOC_90/A NAND2X1_LOC_316/a_36_24# 0.00fF
C48719 NAND2X1_LOC_656/Y NAND2X1_LOC_477/A 0.03fF
C48720 NOR2X1_LOC_536/Y INVX1_LOC_76/A 0.14fF
C48721 INVX1_LOC_75/A INVX1_LOC_111/A 0.02fF
C48722 NOR2X1_LOC_433/A NOR2X1_LOC_153/a_36_216# 0.01fF
C48723 NAND2X1_LOC_338/B INVX1_LOC_137/Y 0.02fF
C48724 INVX1_LOC_17/Y NOR2X1_LOC_88/Y 0.01fF
C48725 INVX1_LOC_55/Y NOR2X1_LOC_718/Y 0.00fF
C48726 INVX1_LOC_117/A NOR2X1_LOC_852/Y 0.02fF
C48727 NAND2X1_LOC_722/A INVX1_LOC_229/Y 0.10fF
C48728 NAND2X1_LOC_736/Y NAND2X1_LOC_866/B 0.02fF
C48729 INVX1_LOC_72/A INVX1_LOC_309/A 0.03fF
C48730 INVX1_LOC_18/A NOR2X1_LOC_167/Y 0.03fF
C48731 INVX1_LOC_181/Y NOR2X1_LOC_74/A 0.01fF
C48732 INVX1_LOC_89/A NOR2X1_LOC_309/Y 0.03fF
C48733 INVX1_LOC_53/A NOR2X1_LOC_830/a_36_216# 0.00fF
C48734 INVX1_LOC_273/A INVX1_LOC_264/A 0.00fF
C48735 INVX1_LOC_226/Y NAND2X1_LOC_565/B 0.40fF
C48736 NAND2X1_LOC_30/Y NAND2X1_LOC_1/Y 1.20fF
C48737 INVX1_LOC_145/Y NAND2X1_LOC_342/Y 0.09fF
C48738 NOR2X1_LOC_238/Y NOR2X1_LOC_754/a_36_216# 0.00fF
C48739 NAND2X1_LOC_799/A INVX1_LOC_76/A 0.23fF
C48740 INVX1_LOC_166/A NAND2X1_LOC_659/A 0.38fF
C48741 INVX1_LOC_181/Y NOR2X1_LOC_9/Y 0.01fF
C48742 NOR2X1_LOC_590/A NOR2X1_LOC_631/B 0.07fF
C48743 INVX1_LOC_230/Y INVX1_LOC_74/A 0.03fF
C48744 NOR2X1_LOC_401/Y NOR2X1_LOC_123/B 0.01fF
C48745 INVX1_LOC_72/A INVX1_LOC_91/A 0.25fF
C48746 NOR2X1_LOC_250/A INVX1_LOC_46/A 0.04fF
C48747 NOR2X1_LOC_67/A D_INPUT_0 0.31fF
C48748 INVX1_LOC_200/Y INVX1_LOC_84/A 0.04fF
C48749 NOR2X1_LOC_82/a_36_216# NOR2X1_LOC_78/A 0.00fF
C48750 INVX1_LOC_161/Y NOR2X1_LOC_137/Y 0.02fF
C48751 INPUT_0 NOR2X1_LOC_387/Y 0.01fF
C48752 NOR2X1_LOC_385/Y NAND2X1_LOC_811/Y 0.00fF
C48753 NOR2X1_LOC_78/B NOR2X1_LOC_106/A 0.01fF
C48754 NAND2X1_LOC_734/B NAND2X1_LOC_807/Y 0.03fF
C48755 INVX1_LOC_282/Y NAND2X1_LOC_866/B 0.23fF
C48756 NAND2X1_LOC_471/Y NAND2X1_LOC_254/Y 0.01fF
C48757 INVX1_LOC_34/A NAND2X1_LOC_849/A 0.06fF
C48758 INVX1_LOC_172/A NOR2X1_LOC_167/Y 0.01fF
C48759 NOR2X1_LOC_321/Y INVX1_LOC_9/A 0.03fF
C48760 NAND2X1_LOC_562/a_36_24# NAND2X1_LOC_659/B 0.01fF
C48761 NAND2X1_LOC_286/B NAND2X1_LOC_81/B 0.00fF
C48762 NOR2X1_LOC_632/Y NAND2X1_LOC_664/a_36_24# 0.00fF
C48763 INVX1_LOC_72/A INVX1_LOC_11/Y 0.03fF
C48764 INVX1_LOC_30/A INVX1_LOC_147/Y 0.06fF
C48765 INVX1_LOC_226/Y NOR2X1_LOC_130/A 0.03fF
C48766 NAND2X1_LOC_198/B INVX1_LOC_70/Y 0.10fF
C48767 NOR2X1_LOC_373/a_36_216# INVX1_LOC_6/A 0.00fF
C48768 INVX1_LOC_11/A INVX1_LOC_44/A 0.07fF
C48769 NAND2X1_LOC_41/Y NOR2X1_LOC_199/B 0.17fF
C48770 NOR2X1_LOC_590/A INVX1_LOC_37/A 9.27fF
C48771 INVX1_LOC_177/A NOR2X1_LOC_569/a_36_216# 0.00fF
C48772 INVX1_LOC_30/A INVX1_LOC_20/A 0.35fF
C48773 NOR2X1_LOC_7/Y NOR2X1_LOC_152/Y 0.11fF
C48774 INVX1_LOC_2/A NOR2X1_LOC_135/Y 0.03fF
C48775 INVX1_LOC_278/Y INVX1_LOC_90/A 0.21fF
C48776 NOR2X1_LOC_88/Y NOR2X1_LOC_406/A 0.03fF
C48777 NOR2X1_LOC_804/B NOR2X1_LOC_703/Y 0.29fF
C48778 INPUT_0 NOR2X1_LOC_514/Y 0.05fF
C48779 INVX1_LOC_64/A NAND2X1_LOC_475/Y 0.01fF
C48780 NOR2X1_LOC_68/A NOR2X1_LOC_56/Y 0.07fF
C48781 INVX1_LOC_136/A NOR2X1_LOC_253/Y 0.01fF
C48782 NOR2X1_LOC_454/Y NOR2X1_LOC_433/Y 0.01fF
C48783 NOR2X1_LOC_769/B NOR2X1_LOC_48/Y 0.01fF
C48784 NAND2X1_LOC_357/B INPUT_0 0.10fF
C48785 NAND2X1_LOC_349/B INVX1_LOC_313/A 0.03fF
C48786 NOR2X1_LOC_100/A NAND2X1_LOC_348/A 0.04fF
C48787 NOR2X1_LOC_25/Y NOR2X1_LOC_59/a_36_216# 0.00fF
C48788 INVX1_LOC_41/A INVX1_LOC_78/Y 0.05fF
C48789 NOR2X1_LOC_246/Y INVX1_LOC_53/Y 0.01fF
C48790 INVX1_LOC_50/A INVX1_LOC_109/Y 0.09fF
C48791 NOR2X1_LOC_598/B NOR2X1_LOC_48/Y 0.00fF
C48792 INVX1_LOC_10/A NOR2X1_LOC_525/a_36_216# 0.00fF
C48793 INVX1_LOC_18/A INVX1_LOC_76/A 0.30fF
C48794 INVX1_LOC_24/A NOR2X1_LOC_799/B 0.03fF
C48795 NAND2X1_LOC_667/a_36_24# NOR2X1_LOC_188/A 0.02fF
C48796 INVX1_LOC_10/A NAND2X1_LOC_800/Y 0.03fF
C48797 NAND2X1_LOC_860/A NAND2X1_LOC_81/B 0.07fF
C48798 NAND2X1_LOC_728/Y INVX1_LOC_76/A 0.07fF
C48799 INVX1_LOC_10/A NOR2X1_LOC_130/A 0.09fF
C48800 NAND2X1_LOC_807/Y INVX1_LOC_25/Y 0.08fF
C48801 NAND2X1_LOC_560/A NAND2X1_LOC_852/Y 0.01fF
C48802 NOR2X1_LOC_750/A INVX1_LOC_232/A 0.12fF
C48803 INVX1_LOC_33/A NOR2X1_LOC_318/B 1.01fF
C48804 NOR2X1_LOC_554/B D_INPUT_3 0.07fF
C48805 INVX1_LOC_11/A NOR2X1_LOC_641/Y 0.04fF
C48806 INVX1_LOC_98/A INVX1_LOC_8/A 0.01fF
C48807 NOR2X1_LOC_68/A VDD 5.64fF
C48808 NOR2X1_LOC_78/A INVX1_LOC_8/A 0.14fF
C48809 NAND2X1_LOC_711/B INVX1_LOC_76/A 0.09fF
C48810 INVX1_LOC_13/Y NOR2X1_LOC_662/A 0.01fF
C48811 INVX1_LOC_209/Y NOR2X1_LOC_56/a_36_216# 0.00fF
C48812 NAND2X1_LOC_223/A INVX1_LOC_87/A 0.02fF
C48813 INVX1_LOC_33/A INVX1_LOC_93/Y 0.07fF
C48814 INVX1_LOC_142/A INVX1_LOC_117/A 0.07fF
C48815 NAND2X1_LOC_500/Y INVX1_LOC_38/A 0.01fF
C48816 NOR2X1_LOC_644/A INVX1_LOC_279/A 0.03fF
C48817 INVX1_LOC_120/A INVX1_LOC_62/A 0.15fF
C48818 INVX1_LOC_113/Y NAND2X1_LOC_212/Y 0.02fF
C48819 INVX1_LOC_73/Y NOR2X1_LOC_155/A 0.01fF
C48820 NAND2X1_LOC_36/A INVX1_LOC_38/A 0.46fF
C48821 NOR2X1_LOC_580/a_36_216# NAND2X1_LOC_463/B 0.00fF
C48822 NOR2X1_LOC_122/Y NAND2X1_LOC_656/Y 0.04fF
C48823 NOR2X1_LOC_237/Y NAND2X1_LOC_244/A 0.00fF
C48824 INVX1_LOC_103/A NOR2X1_LOC_841/A 0.02fF
C48825 NOR2X1_LOC_68/A NOR2X1_LOC_684/a_36_216# 0.00fF
C48826 NOR2X1_LOC_545/A VDD -0.00fF
C48827 INVX1_LOC_198/Y NOR2X1_LOC_698/Y 0.05fF
C48828 NOR2X1_LOC_666/Y NOR2X1_LOC_66/Y 0.25fF
C48829 NOR2X1_LOC_590/A NOR2X1_LOC_743/Y 0.57fF
C48830 NOR2X1_LOC_186/Y INVX1_LOC_29/A 0.13fF
C48831 INVX1_LOC_11/A NOR2X1_LOC_461/B 0.00fF
C48832 INVX1_LOC_48/Y INVX1_LOC_293/Y -0.01fF
C48833 NOR2X1_LOC_216/Y INVX1_LOC_10/A 0.02fF
C48834 NOR2X1_LOC_298/Y NOR2X1_LOC_380/Y 0.14fF
C48835 INVX1_LOC_25/Y INVX1_LOC_6/A 0.06fF
C48836 INVX1_LOC_113/Y INVX1_LOC_14/Y 0.03fF
C48837 NOR2X1_LOC_392/B INVX1_LOC_59/Y 0.01fF
C48838 NAND2X1_LOC_338/B INVX1_LOC_91/A 0.07fF
C48839 INVX1_LOC_205/A INVX1_LOC_9/A 0.00fF
C48840 NOR2X1_LOC_599/Y NAND2X1_LOC_810/B 0.01fF
C48841 NOR2X1_LOC_188/A NOR2X1_LOC_188/Y 0.01fF
C48842 NAND2X1_LOC_624/B INVX1_LOC_3/Y 0.00fF
C48843 NOR2X1_LOC_419/Y NAND2X1_LOC_96/A 0.04fF
C48844 NAND2X1_LOC_573/Y INVX1_LOC_29/A 0.08fF
C48845 NAND2X1_LOC_860/A INVX1_LOC_4/Y 0.01fF
C48846 NAND2X1_LOC_363/B INVX1_LOC_4/A 0.00fF
C48847 NAND2X1_LOC_354/B NOR2X1_LOC_681/Y 0.01fF
C48848 INVX1_LOC_48/Y NAND2X1_LOC_74/B 0.03fF
C48849 NOR2X1_LOC_128/B INPUT_0 0.00fF
C48850 NAND2X1_LOC_116/A INVX1_LOC_36/Y 0.02fF
C48851 NOR2X1_LOC_146/Y INVX1_LOC_86/Y 0.25fF
C48852 INVX1_LOC_94/Y NOR2X1_LOC_591/A 0.07fF
C48853 NOR2X1_LOC_607/A INVX1_LOC_9/A 0.01fF
C48854 INVX1_LOC_53/A NOR2X1_LOC_334/Y 0.23fF
C48855 NOR2X1_LOC_78/A NOR2X1_LOC_315/a_36_216# 0.00fF
C48856 NOR2X1_LOC_644/A INVX1_LOC_182/Y 0.56fF
C48857 INVX1_LOC_89/A NOR2X1_LOC_208/A 0.07fF
C48858 NAND2X1_LOC_838/a_36_24# NOR2X1_LOC_536/A 0.00fF
C48859 NOR2X1_LOC_238/Y INVX1_LOC_54/A 0.01fF
C48860 INVX1_LOC_8/A NOR2X1_LOC_98/a_36_216# 0.01fF
C48861 NOR2X1_LOC_709/A INVX1_LOC_46/A 0.13fF
C48862 INVX1_LOC_72/Y NOR2X1_LOC_101/a_36_216# 0.03fF
C48863 INVX1_LOC_24/A INVX1_LOC_307/A 0.07fF
C48864 NOR2X1_LOC_596/A INVX1_LOC_179/A 0.04fF
C48865 INVX1_LOC_276/A NOR2X1_LOC_682/Y 0.01fF
C48866 INVX1_LOC_77/A NOR2X1_LOC_433/Y 0.03fF
C48867 NOR2X1_LOC_698/a_36_216# INVX1_LOC_15/A 0.02fF
C48868 INVX1_LOC_47/A INVX1_LOC_286/A 0.01fF
C48869 INVX1_LOC_24/A NOR2X1_LOC_445/B 0.07fF
C48870 NOR2X1_LOC_593/Y NOR2X1_LOC_641/Y 0.04fF
C48871 NOR2X1_LOC_226/A NAND2X1_LOC_262/a_36_24# 0.00fF
C48872 INVX1_LOC_303/A NAND2X1_LOC_487/a_36_24# 0.00fF
C48873 NOR2X1_LOC_45/Y INVX1_LOC_29/A 0.03fF
C48874 INVX1_LOC_135/A NOR2X1_LOC_45/B 0.01fF
C48875 NOR2X1_LOC_530/Y NOR2X1_LOC_671/Y 0.00fF
C48876 INVX1_LOC_266/A INVX1_LOC_32/A 0.39fF
C48877 NOR2X1_LOC_510/Y NAND2X1_LOC_454/Y 0.01fF
C48878 NOR2X1_LOC_180/Y NOR2X1_LOC_331/B 0.10fF
C48879 NAND2X1_LOC_140/A NOR2X1_LOC_78/A 0.05fF
C48880 INVX1_LOC_58/A NOR2X1_LOC_604/a_36_216# 0.00fF
C48881 NOR2X1_LOC_815/Y INVX1_LOC_291/A 0.01fF
C48882 NAND2X1_LOC_198/B INVX1_LOC_285/A 0.10fF
C48883 NAND2X1_LOC_656/A NAND2X1_LOC_572/B 0.20fF
C48884 NOR2X1_LOC_381/Y INVX1_LOC_32/A 0.04fF
C48885 INVX1_LOC_200/Y INVX1_LOC_278/A 0.01fF
C48886 INVX1_LOC_33/A INVX1_LOC_117/Y 0.03fF
C48887 INVX1_LOC_276/A NAND2X1_LOC_848/A 0.22fF
C48888 NOR2X1_LOC_690/Y INVX1_LOC_76/A 0.08fF
C48889 INVX1_LOC_313/Y INVX1_LOC_91/A 0.19fF
C48890 NOR2X1_LOC_67/A NAND2X1_LOC_848/A 0.07fF
C48891 NOR2X1_LOC_92/Y INVX1_LOC_128/Y 1.53fF
C48892 NOR2X1_LOC_392/Y NOR2X1_LOC_416/A 0.04fF
C48893 INVX1_LOC_21/A NOR2X1_LOC_278/Y 0.10fF
C48894 INVX1_LOC_75/A INVX1_LOC_6/A 0.16fF
C48895 INVX1_LOC_27/A INVX1_LOC_26/A 0.05fF
C48896 NOR2X1_LOC_772/B INVX1_LOC_57/A 0.43fF
C48897 NOR2X1_LOC_718/B INVX1_LOC_92/A 0.14fF
C48898 NOR2X1_LOC_458/B NOR2X1_LOC_331/B 0.01fF
C48899 NOR2X1_LOC_457/A INVX1_LOC_4/A 1.74fF
C48900 NOR2X1_LOC_495/Y INVX1_LOC_84/A 0.01fF
C48901 INVX1_LOC_64/A NAND2X1_LOC_787/A 0.03fF
C48902 NAND2X1_LOC_740/Y INVX1_LOC_50/A 0.04fF
C48903 NOR2X1_LOC_312/Y NOR2X1_LOC_279/Y 0.19fF
C48904 NOR2X1_LOC_288/A NOR2X1_LOC_634/A 0.01fF
C48905 INVX1_LOC_278/Y INVX1_LOC_38/A 1.35fF
C48906 NAND2X1_LOC_656/A NAND2X1_LOC_219/B 0.21fF
C48907 INVX1_LOC_13/Y INVX1_LOC_57/A 0.10fF
C48908 NAND2X1_LOC_479/Y INVX1_LOC_281/A 0.07fF
C48909 INVX1_LOC_64/A NAND2X1_LOC_363/B 0.07fF
C48910 NAND2X1_LOC_214/B NOR2X1_LOC_255/Y 0.02fF
C48911 NOR2X1_LOC_659/a_36_216# INVX1_LOC_109/Y 0.01fF
C48912 NOR2X1_LOC_763/Y INVX1_LOC_37/A 0.01fF
C48913 INVX1_LOC_50/Y NOR2X1_LOC_622/A 0.11fF
C48914 NOR2X1_LOC_598/B INVX1_LOC_204/Y 0.03fF
C48915 NOR2X1_LOC_454/Y NOR2X1_LOC_651/a_36_216# 0.01fF
C48916 NAND2X1_LOC_833/Y NOR2X1_LOC_661/A 0.03fF
C48917 NAND2X1_LOC_841/A INVX1_LOC_54/A 0.01fF
C48918 NAND2X1_LOC_112/Y INVX1_LOC_118/Y 0.03fF
C48919 NOR2X1_LOC_658/a_36_216# NAND2X1_LOC_67/Y 0.01fF
C48920 INVX1_LOC_24/A INVX1_LOC_12/A 0.70fF
C48921 INVX1_LOC_50/A NAND2X1_LOC_706/Y 0.28fF
C48922 NOR2X1_LOC_296/a_36_216# INVX1_LOC_23/Y 0.01fF
C48923 NOR2X1_LOC_67/A INVX1_LOC_46/Y 0.15fF
C48924 NOR2X1_LOC_742/A NOR2X1_LOC_486/Y 0.07fF
C48925 NAND2X1_LOC_799/Y INVX1_LOC_84/A 0.15fF
C48926 INVX1_LOC_69/Y NOR2X1_LOC_355/B 0.00fF
C48927 INVX1_LOC_268/A INVX1_LOC_54/A 0.32fF
C48928 INVX1_LOC_222/Y INVX1_LOC_58/Y 0.12fF
C48929 INVX1_LOC_219/Y INVX1_LOC_84/A 0.03fF
C48930 NOR2X1_LOC_350/A NAND2X1_LOC_74/B 0.06fF
C48931 NOR2X1_LOC_220/A INVX1_LOC_179/A 0.18fF
C48932 NOR2X1_LOC_666/A INVX1_LOC_271/A 0.00fF
C48933 NOR2X1_LOC_637/B INVX1_LOC_272/A 0.02fF
C48934 NAND2X1_LOC_808/A NAND2X1_LOC_603/a_36_24# 0.00fF
C48935 INVX1_LOC_30/A INVX1_LOC_4/A 0.11fF
C48936 INVX1_LOC_132/A INVX1_LOC_29/A 0.07fF
C48937 NAND2X1_LOC_348/A NOR2X1_LOC_124/a_36_216# 0.00fF
C48938 NOR2X1_LOC_590/A NAND2X1_LOC_72/B 0.44fF
C48939 INVX1_LOC_64/A NOR2X1_LOC_791/Y 0.00fF
C48940 NAND2X1_LOC_348/A INVX1_LOC_59/Y 0.86fF
C48941 INVX1_LOC_72/A INVX1_LOC_231/A 0.05fF
C48942 NAND2X1_LOC_348/A INVX1_LOC_112/A 0.01fF
C48943 NOR2X1_LOC_481/A INVX1_LOC_29/A 0.01fF
C48944 INVX1_LOC_88/A INVX1_LOC_57/A 0.01fF
C48945 NAND2X1_LOC_640/Y INVX1_LOC_29/A 0.15fF
C48946 NOR2X1_LOC_500/Y NOR2X1_LOC_197/B 0.10fF
C48947 NOR2X1_LOC_76/A NOR2X1_LOC_536/A 0.07fF
C48948 NAND2X1_LOC_348/A INVX1_LOC_176/A 0.03fF
C48949 NOR2X1_LOC_111/Y NOR2X1_LOC_111/A 0.02fF
C48950 NOR2X1_LOC_557/Y INVX1_LOC_12/A 0.07fF
C48951 NOR2X1_LOC_639/a_36_216# INVX1_LOC_118/A 0.02fF
C48952 NAND2X1_LOC_863/A INVX1_LOC_46/A 0.19fF
C48953 INVX1_LOC_161/Y NOR2X1_LOC_677/Y 0.02fF
C48954 D_INPUT_0 NOR2X1_LOC_729/A 0.05fF
C48955 INVX1_LOC_225/A INVX1_LOC_29/A 0.22fF
C48956 NOR2X1_LOC_389/A NAND2X1_LOC_288/B 0.03fF
C48957 INVX1_LOC_286/A INVX1_LOC_95/Y 0.09fF
C48958 INVX1_LOC_232/A INVX1_LOC_123/Y 0.05fF
C48959 NOR2X1_LOC_617/Y INVX1_LOC_3/Y 0.00fF
C48960 NOR2X1_LOC_401/B INVX1_LOC_63/A 0.08fF
C48961 NOR2X1_LOC_2/Y VDD 0.51fF
C48962 NOR2X1_LOC_589/A INVX1_LOC_113/A 0.14fF
C48963 NOR2X1_LOC_323/Y NAND2X1_LOC_721/A 0.01fF
C48964 NOR2X1_LOC_690/A INVX1_LOC_42/A 0.13fF
C48965 INVX1_LOC_53/Y INVX1_LOC_285/A 0.21fF
C48966 INVX1_LOC_77/A INVX1_LOC_47/Y 0.03fF
C48967 NOR2X1_LOC_84/Y NAND2X1_LOC_74/B 0.06fF
C48968 NOR2X1_LOC_516/B NOR2X1_LOC_673/A 0.03fF
C48969 NOR2X1_LOC_413/Y INVX1_LOC_42/A 0.06fF
C48970 NOR2X1_LOC_52/Y NOR2X1_LOC_449/A 0.01fF
C48971 NOR2X1_LOC_202/Y INVX1_LOC_281/A 0.02fF
C48972 NAND2X1_LOC_319/A NOR2X1_LOC_88/Y 0.49fF
C48973 NOR2X1_LOC_550/a_36_216# NOR2X1_LOC_383/B 0.00fF
C48974 NOR2X1_LOC_62/a_36_216# INVX1_LOC_3/A 0.02fF
C48975 NOR2X1_LOC_456/Y NOR2X1_LOC_794/B 0.00fF
C48976 INVX1_LOC_73/A NOR2X1_LOC_536/A 0.03fF
C48977 INVX1_LOC_5/A INVX1_LOC_14/A 0.31fF
C48978 INVX1_LOC_190/A NAND2X1_LOC_798/B 0.02fF
C48979 NOR2X1_LOC_790/B INVX1_LOC_225/Y 0.24fF
C48980 NAND2X1_LOC_361/Y INVX1_LOC_15/A 0.09fF
C48981 INVX1_LOC_64/A NOR2X1_LOC_457/A 0.03fF
C48982 INVX1_LOC_292/A NOR2X1_LOC_493/a_36_216# 0.00fF
C48983 INVX1_LOC_96/A NOR2X1_LOC_357/Y 0.02fF
C48984 NAND2X1_LOC_737/a_36_24# INVX1_LOC_296/A 0.00fF
C48985 NOR2X1_LOC_106/Y INVX1_LOC_78/A 0.04fF
C48986 NAND2X1_LOC_741/B INVX1_LOC_296/Y 0.03fF
C48987 INVX1_LOC_95/A INVX1_LOC_95/Y 0.29fF
C48988 INVX1_LOC_143/A INVX1_LOC_12/A 0.15fF
C48989 NOR2X1_LOC_500/B INVX1_LOC_57/A 0.07fF
C48990 NAND2X1_LOC_319/A INVX1_LOC_84/A 0.03fF
C48991 INVX1_LOC_24/A NOR2X1_LOC_686/A 0.01fF
C48992 NAND2X1_LOC_851/a_36_24# INVX1_LOC_33/Y 0.00fF
C48993 NOR2X1_LOC_6/B INVX1_LOC_32/A 0.13fF
C48994 NAND2X1_LOC_391/Y NOR2X1_LOC_103/Y 0.03fF
C48995 NOR2X1_LOC_637/Y NOR2X1_LOC_447/A 0.06fF
C48996 INVX1_LOC_35/A INVX1_LOC_277/A 0.42fF
C48997 INVX1_LOC_124/A INVX1_LOC_47/Y -0.03fF
C48998 INVX1_LOC_153/Y NAND2X1_LOC_454/Y 0.10fF
C48999 INVX1_LOC_36/A NOR2X1_LOC_392/Y 0.07fF
C49000 INVX1_LOC_49/A NAND2X1_LOC_61/Y 0.05fF
C49001 INVX1_LOC_64/A INVX1_LOC_30/A 0.97fF
C49002 NOR2X1_LOC_791/Y INVX1_LOC_43/Y 0.02fF
C49003 NOR2X1_LOC_45/B NOR2X1_LOC_813/Y 0.07fF
C49004 NOR2X1_LOC_91/A NOR2X1_LOC_577/Y 0.14fF
C49005 NAND2X1_LOC_810/a_36_24# NOR2X1_LOC_829/A 0.00fF
C49006 INVX1_LOC_58/A INVX1_LOC_41/Y 0.03fF
C49007 INVX1_LOC_89/A INVX1_LOC_63/A 5.21fF
C49008 INPUT_1 NAND2X1_LOC_42/a_36_24# 0.00fF
C49009 INVX1_LOC_5/A NOR2X1_LOC_717/Y 0.07fF
C49010 NAND2X1_LOC_832/Y NOR2X1_LOC_433/Y 0.40fF
C49011 NOR2X1_LOC_279/Y NAND2X1_LOC_287/B 0.03fF
C49012 INVX1_LOC_17/A INVX1_LOC_269/A 0.13fF
C49013 INVX1_LOC_303/A INVX1_LOC_57/A 0.20fF
C49014 NOR2X1_LOC_45/B INVX1_LOC_280/A 0.30fF
C49015 NOR2X1_LOC_151/a_36_216# NOR2X1_LOC_155/A 0.00fF
C49016 INVX1_LOC_225/A NOR2X1_LOC_281/Y 0.01fF
C49017 INVX1_LOC_41/A NOR2X1_LOC_727/B 0.04fF
C49018 INVX1_LOC_236/A INVX1_LOC_273/A 0.01fF
C49019 NOR2X1_LOC_634/B NOR2X1_LOC_334/Y 0.02fF
C49020 NOR2X1_LOC_558/A NOR2X1_LOC_266/B 0.02fF
C49021 NOR2X1_LOC_577/Y INVX1_LOC_23/A 0.10fF
C49022 INVX1_LOC_63/Y NOR2X1_LOC_383/B 0.07fF
C49023 NAND2X1_LOC_800/Y INVX1_LOC_12/A 0.03fF
C49024 NOR2X1_LOC_32/B D_INPUT_2 0.14fF
C49025 INVX1_LOC_14/A NAND2X1_LOC_337/B 0.01fF
C49026 NOR2X1_LOC_78/B NOR2X1_LOC_334/Y 0.14fF
C49027 NOR2X1_LOC_130/A INVX1_LOC_12/A 2.56fF
C49028 INVX1_LOC_136/A NAND2X1_LOC_794/B 0.07fF
C49029 NOR2X1_LOC_381/Y INPUT_3 0.08fF
C49030 INVX1_LOC_251/Y NAND2X1_LOC_437/a_36_24# 0.01fF
C49031 INVX1_LOC_30/Y INVX1_LOC_32/A 0.03fF
C49032 D_INPUT_1 INVX1_LOC_155/Y 0.05fF
C49033 NOR2X1_LOC_510/Y NOR2X1_LOC_68/A 0.03fF
C49034 INVX1_LOC_21/A INVX1_LOC_122/Y 0.55fF
C49035 NAND2X1_LOC_555/Y INVX1_LOC_269/A 0.01fF
C49036 INVX1_LOC_2/A NAND2X1_LOC_61/Y 0.09fF
C49037 INVX1_LOC_255/Y NOR2X1_LOC_38/B 0.68fF
C49038 NAND2X1_LOC_853/Y NOR2X1_LOC_409/B 0.03fF
C49039 NOR2X1_LOC_473/B NOR2X1_LOC_89/A 0.12fF
C49040 NOR2X1_LOC_629/B INVX1_LOC_23/A 0.01fF
C49041 INVX1_LOC_41/A NOR2X1_LOC_717/A 0.00fF
C49042 INVX1_LOC_136/A INVX1_LOC_48/Y 0.02fF
C49043 INVX1_LOC_139/Y INVX1_LOC_281/A 0.00fF
C49044 NOR2X1_LOC_113/B NOR2X1_LOC_814/A 0.76fF
C49045 INVX1_LOC_34/A NAND2X1_LOC_549/Y 0.00fF
C49046 NOR2X1_LOC_564/Y INVX1_LOC_99/A 0.06fF
C49047 NOR2X1_LOC_445/Y NAND2X1_LOC_72/Y 0.14fF
C49048 NOR2X1_LOC_191/B NAND2X1_LOC_474/Y 0.01fF
C49049 INVX1_LOC_75/A INVX1_LOC_301/A 0.04fF
C49050 NAND2X1_LOC_561/B NOR2X1_LOC_384/Y 0.04fF
C49051 NAND2X1_LOC_35/Y NAND2X1_LOC_483/Y 0.07fF
C49052 INVX1_LOC_213/Y NOR2X1_LOC_678/A 0.00fF
C49053 NOR2X1_LOC_272/Y INVX1_LOC_81/A 0.03fF
C49054 NAND2X1_LOC_725/A NAND2X1_LOC_736/B 0.00fF
C49055 INVX1_LOC_225/A NAND2X1_LOC_385/a_36_24# 0.01fF
C49056 INVX1_LOC_21/A NAND2X1_LOC_7/Y 0.05fF
C49057 NAND2X1_LOC_348/A NOR2X1_LOC_340/A 0.02fF
C49058 INVX1_LOC_315/Y NOR2X1_LOC_673/A 2.77fF
C49059 NAND2X1_LOC_9/Y NOR2X1_LOC_709/A 0.08fF
C49060 NOR2X1_LOC_32/B NOR2X1_LOC_529/Y 0.03fF
C49061 INVX1_LOC_5/A INVX1_LOC_217/Y 0.00fF
C49062 NOR2X1_LOC_361/B NOR2X1_LOC_68/A 0.11fF
C49063 NOR2X1_LOC_632/Y NOR2X1_LOC_631/Y 0.03fF
C49064 INVX1_LOC_290/A NOR2X1_LOC_45/a_36_216# 0.01fF
C49065 NOR2X1_LOC_322/Y NOR2X1_LOC_89/A 0.14fF
C49066 NOR2X1_LOC_91/A INVX1_LOC_22/A 0.15fF
C49067 NOR2X1_LOC_92/Y NOR2X1_LOC_13/Y 0.10fF
C49068 INVX1_LOC_83/A NOR2X1_LOC_334/Y 0.03fF
C49069 NOR2X1_LOC_273/Y INVX1_LOC_1/A 0.04fF
C49070 INVX1_LOC_223/Y NOR2X1_LOC_804/B 0.01fF
C49071 NOR2X1_LOC_703/B NOR2X1_LOC_541/Y 0.02fF
C49072 INVX1_LOC_64/A NAND2X1_LOC_722/A 0.07fF
C49073 INVX1_LOC_288/Y INVX1_LOC_290/A 0.01fF
C49074 INVX1_LOC_89/A NAND2X1_LOC_452/Y 0.01fF
C49075 INVX1_LOC_216/A NOR2X1_LOC_660/Y 0.01fF
C49076 NAND2X1_LOC_654/B INVX1_LOC_15/A 0.02fF
C49077 NOR2X1_LOC_262/a_36_216# INVX1_LOC_22/A 0.00fF
C49078 INVX1_LOC_36/A NOR2X1_LOC_599/Y 0.03fF
C49079 INVX1_LOC_234/A INVX1_LOC_26/A 0.00fF
C49080 INVX1_LOC_6/Y NOR2X1_LOC_666/A 0.06fF
C49081 NAND2X1_LOC_303/Y NOR2X1_LOC_152/Y 0.10fF
C49082 INVX1_LOC_217/Y INVX1_LOC_178/A 0.01fF
C49083 INVX1_LOC_256/A NOR2X1_LOC_457/B 0.38fF
C49084 NOR2X1_LOC_325/A INVX1_LOC_23/A 0.37fF
C49085 INVX1_LOC_200/A INVX1_LOC_24/A 3.50fF
C49086 INVX1_LOC_28/A NAND2X1_LOC_647/B 0.04fF
C49087 INVX1_LOC_1/A NOR2X1_LOC_550/B 0.10fF
C49088 INVX1_LOC_22/A INVX1_LOC_23/A 1.79fF
C49089 NOR2X1_LOC_557/a_36_216# NOR2X1_LOC_814/A 0.01fF
C49090 NOR2X1_LOC_220/A NOR2X1_LOC_405/Y 0.02fF
C49091 INVX1_LOC_31/A NOR2X1_LOC_274/B 0.04fF
C49092 NOR2X1_LOC_368/A INVX1_LOC_170/Y 0.00fF
C49093 NOR2X1_LOC_92/Y NAND2X1_LOC_175/B 0.12fF
C49094 NOR2X1_LOC_793/Y INVX1_LOC_49/A 0.08fF
C49095 NAND2X1_LOC_623/a_36_24# NAND2X1_LOC_374/Y 0.00fF
C49096 NOR2X1_LOC_127/a_36_216# INVX1_LOC_76/A 0.01fF
C49097 NAND2X1_LOC_472/Y INVX1_LOC_92/A 0.18fF
C49098 NOR2X1_LOC_798/A NOR2X1_LOC_709/A 0.03fF
C49099 INVX1_LOC_101/A INVX1_LOC_29/Y 0.05fF
C49100 NOR2X1_LOC_826/Y NAND2X1_LOC_859/B 0.01fF
C49101 NOR2X1_LOC_590/A NAND2X1_LOC_198/B 0.03fF
C49102 INVX1_LOC_6/A INVX1_LOC_283/A 0.00fF
C49103 INVX1_LOC_45/A NOR2X1_LOC_703/B 0.03fF
C49104 INVX1_LOC_103/A NOR2X1_LOC_172/Y 0.02fF
C49105 NOR2X1_LOC_569/Y INVX1_LOC_53/A 0.02fF
C49106 NOR2X1_LOC_703/A NAND2X1_LOC_72/B 0.00fF
C49107 NAND2X1_LOC_53/Y INVX1_LOC_283/Y -0.01fF
C49108 NAND2X1_LOC_711/B NAND2X1_LOC_188/a_36_24# 0.00fF
C49109 NOR2X1_LOC_703/B NOR2X1_LOC_568/A 0.00fF
C49110 NAND2X1_LOC_642/Y INVX1_LOC_29/A 1.72fF
C49111 NOR2X1_LOC_255/Y INVX1_LOC_234/A 0.00fF
C49112 NAND2X1_LOC_733/Y INVX1_LOC_24/A 0.20fF
C49113 INVX1_LOC_36/A NOR2X1_LOC_765/a_36_216# 0.04fF
C49114 NOR2X1_LOC_791/Y NAND2X1_LOC_850/Y 0.02fF
C49115 INVX1_LOC_1/A INVX1_LOC_249/Y 0.02fF
C49116 INVX1_LOC_130/Y INVX1_LOC_30/A 0.03fF
C49117 NOR2X1_LOC_784/B INVX1_LOC_23/A 0.01fF
C49118 NAND2X1_LOC_47/a_36_24# INVX1_LOC_49/A 0.00fF
C49119 INVX1_LOC_35/A INVX1_LOC_174/Y 0.02fF
C49120 INVX1_LOC_124/Y INVX1_LOC_181/Y 0.02fF
C49121 NOR2X1_LOC_82/A INVX1_LOC_33/A 1.32fF
C49122 NOR2X1_LOC_794/B NOR2X1_LOC_550/B 0.01fF
C49123 INVX1_LOC_311/Y NOR2X1_LOC_306/a_36_216# 0.00fF
C49124 NOR2X1_LOC_355/A INVX1_LOC_29/Y 0.08fF
C49125 NAND2X1_LOC_670/a_36_24# NOR2X1_LOC_360/Y 0.00fF
C49126 NOR2X1_LOC_92/Y NOR2X1_LOC_504/Y 0.01fF
C49127 INVX1_LOC_225/Y NOR2X1_LOC_344/A 0.10fF
C49128 VDD NAND2X1_LOC_768/Y 0.00fF
C49129 NAND2X1_LOC_357/A NOR2X1_LOC_309/Y 0.12fF
C49130 INVX1_LOC_31/A NOR2X1_LOC_577/Y 0.49fF
C49131 NAND2X1_LOC_637/Y INVX1_LOC_92/A 0.02fF
C49132 INVX1_LOC_244/Y INVX1_LOC_72/A 0.02fF
C49133 INVX1_LOC_50/A NOR2X1_LOC_597/A 0.01fF
C49134 INVX1_LOC_95/Y NAND2X1_LOC_807/B 0.01fF
C49135 NOR2X1_LOC_92/Y INVX1_LOC_256/Y 0.07fF
C49136 INVX1_LOC_244/A INVX1_LOC_57/A 0.03fF
C49137 NOR2X1_LOC_590/A INVX1_LOC_310/Y 0.36fF
C49138 INVX1_LOC_24/A INVX1_LOC_217/A 0.24fF
C49139 INVX1_LOC_285/Y NAND2X1_LOC_454/Y 0.10fF
C49140 NOR2X1_LOC_329/B NOR2X1_LOC_654/A 0.00fF
C49141 NOR2X1_LOC_703/B INVX1_LOC_71/A 0.03fF
C49142 INVX1_LOC_292/A NOR2X1_LOC_392/B 0.01fF
C49143 INPUT_3 NOR2X1_LOC_6/B 0.12fF
C49144 NOR2X1_LOC_75/Y NOR2X1_LOC_423/Y 0.31fF
C49145 NAND2X1_LOC_36/A INVX1_LOC_33/A 0.02fF
C49146 NOR2X1_LOC_274/Y INVX1_LOC_18/A 0.00fF
C49147 NOR2X1_LOC_174/B NOR2X1_LOC_434/A 0.00fF
C49148 INVX1_LOC_14/A NOR2X1_LOC_773/Y 0.09fF
C49149 NOR2X1_LOC_360/Y NOR2X1_LOC_303/Y 0.01fF
C49150 INVX1_LOC_75/A INVX1_LOC_270/A 0.16fF
C49151 NOR2X1_LOC_124/A INVX1_LOC_32/A 0.04fF
C49152 NAND2X1_LOC_198/a_36_24# INVX1_LOC_8/A 0.00fF
C49153 INVX1_LOC_307/A NOR2X1_LOC_197/B 0.10fF
C49154 NOR2X1_LOC_243/B NAND2X1_LOC_86/a_36_24# 0.00fF
C49155 INVX1_LOC_136/A INVX1_LOC_231/Y 0.09fF
C49156 INVX1_LOC_170/A INVX1_LOC_8/A 0.20fF
C49157 INVX1_LOC_27/A INVX1_LOC_164/A 0.01fF
C49158 NOR2X1_LOC_91/A INVX1_LOC_100/A 0.05fF
C49159 NAND2X1_LOC_555/Y NAND2X1_LOC_127/a_36_24# 0.01fF
C49160 NAND2X1_LOC_239/a_36_24# NOR2X1_LOC_590/A 0.01fF
C49161 NAND2X1_LOC_640/Y NAND2X1_LOC_634/Y 0.01fF
C49162 NOR2X1_LOC_443/Y INPUT_0 0.55fF
C49163 NOR2X1_LOC_305/Y NOR2X1_LOC_48/B 0.08fF
C49164 NAND2X1_LOC_200/B NOR2X1_LOC_107/Y 0.01fF
C49165 NOR2X1_LOC_75/Y NOR2X1_LOC_222/Y 0.03fF
C49166 NOR2X1_LOC_197/B NOR2X1_LOC_445/B 0.10fF
C49167 NOR2X1_LOC_82/A INVX1_LOC_40/A 0.03fF
C49168 NOR2X1_LOC_831/B NAND2X1_LOC_288/A 0.27fF
C49169 NOR2X1_LOC_68/A INVX1_LOC_153/Y 0.11fF
C49170 NOR2X1_LOC_590/A NAND2X1_LOC_491/a_36_24# 0.01fF
C49171 NOR2X1_LOC_67/A NOR2X1_LOC_134/Y 0.01fF
C49172 INVX1_LOC_21/A NOR2X1_LOC_312/Y 0.24fF
C49173 INVX1_LOC_24/A NAND2X1_LOC_787/B 0.14fF
C49174 NOR2X1_LOC_716/B NAND2X1_LOC_656/A 0.02fF
C49175 NOR2X1_LOC_336/B NOR2X1_LOC_802/A 0.36fF
C49176 NAND2X1_LOC_787/A INVX1_LOC_282/A 0.01fF
C49177 NOR2X1_LOC_820/A NOR2X1_LOC_664/Y 0.01fF
C49178 NOR2X1_LOC_89/A INVX1_LOC_281/Y 0.01fF
C49179 NOR2X1_LOC_145/Y INVX1_LOC_257/A 0.07fF
C49180 INVX1_LOC_100/A INVX1_LOC_23/A 0.28fF
C49181 INVX1_LOC_236/Y INVX1_LOC_248/A 0.01fF
C49182 NOR2X1_LOC_836/Y NOR2X1_LOC_78/B 0.09fF
C49183 INVX1_LOC_31/A NOR2X1_LOC_346/B 0.01fF
C49184 NOR2X1_LOC_175/B INVX1_LOC_31/A 0.10fF
C49185 NOR2X1_LOC_68/A INVX1_LOC_121/Y 0.02fF
C49186 NOR2X1_LOC_103/Y INVX1_LOC_137/Y 0.01fF
C49187 NOR2X1_LOC_237/Y NOR2X1_LOC_373/a_36_216# 0.01fF
C49188 INVX1_LOC_136/A NOR2X1_LOC_84/Y 0.39fF
C49189 NOR2X1_LOC_295/Y INVX1_LOC_45/Y 0.04fF
C49190 NOR2X1_LOC_281/Y NAND2X1_LOC_642/Y 0.01fF
C49191 INVX1_LOC_304/A NOR2X1_LOC_278/Y 0.02fF
C49192 NOR2X1_LOC_89/A INVX1_LOC_193/A 0.24fF
C49193 INVX1_LOC_14/A NOR2X1_LOC_332/A 0.14fF
C49194 INVX1_LOC_136/A NOR2X1_LOC_482/Y 0.94fF
C49195 NOR2X1_LOC_607/Y INVX1_LOC_155/Y 0.01fF
C49196 NOR2X1_LOC_468/Y NOR2X1_LOC_71/Y 0.61fF
C49197 INVX1_LOC_30/A NAND2X1_LOC_850/Y 0.13fF
C49198 NOR2X1_LOC_68/A INVX1_LOC_177/A 0.03fF
C49199 NOR2X1_LOC_590/A INVX1_LOC_53/Y 0.12fF
C49200 INVX1_LOC_49/A NOR2X1_LOC_520/B 0.13fF
C49201 NOR2X1_LOC_820/B NOR2X1_LOC_820/Y 0.03fF
C49202 NOR2X1_LOC_456/a_36_216# NOR2X1_LOC_644/A 0.00fF
C49203 INVX1_LOC_224/Y INVX1_LOC_91/A 0.14fF
C49204 INVX1_LOC_290/A NOR2X1_LOC_276/Y 0.02fF
C49205 NAND2X1_LOC_11/Y D_INPUT_7 0.29fF
C49206 INVX1_LOC_304/Y INVX1_LOC_24/A 0.14fF
C49207 INVX1_LOC_31/A INVX1_LOC_22/A 0.16fF
C49208 NOR2X1_LOC_334/Y INVX1_LOC_46/A 0.14fF
C49209 INVX1_LOC_54/Y NOR2X1_LOC_360/Y 0.03fF
C49210 NOR2X1_LOC_481/A NAND2X1_LOC_310/a_36_24# 0.00fF
C49211 NOR2X1_LOC_15/Y NAND2X1_LOC_551/A 0.02fF
C49212 NOR2X1_LOC_14/a_36_216# NOR2X1_LOC_655/Y 0.00fF
C49213 NOR2X1_LOC_13/Y NAND2X1_LOC_477/A 0.10fF
C49214 NOR2X1_LOC_404/a_36_216# NAND2X1_LOC_463/B 0.00fF
C49215 INVX1_LOC_132/A INVX1_LOC_8/A 0.02fF
C49216 NOR2X1_LOC_831/B INVX1_LOC_19/A 1.15fF
C49217 NAND2X1_LOC_188/a_36_24# NOR2X1_LOC_690/Y 0.00fF
C49218 NOR2X1_LOC_15/Y INVX1_LOC_55/Y 0.07fF
C49219 NOR2X1_LOC_510/Y INVX1_LOC_147/A 0.01fF
C49220 INVX1_LOC_17/A NOR2X1_LOC_814/Y 0.01fF
C49221 INVX1_LOC_32/A NOR2X1_LOC_684/Y 0.03fF
C49222 INVX1_LOC_36/A INVX1_LOC_25/Y 0.03fF
C49223 VDD NOR2X1_LOC_36/A 0.30fF
C49224 INVX1_LOC_103/A INVX1_LOC_90/A 0.10fF
C49225 NAND2X1_LOC_190/Y NOR2X1_LOC_644/A 0.04fF
C49226 NOR2X1_LOC_624/a_36_216# INVX1_LOC_89/A 0.00fF
C49227 INVX1_LOC_24/A NAND2X1_LOC_832/a_36_24# 0.00fF
C49228 INVX1_LOC_36/A NAND2X1_LOC_349/B 0.03fF
C49229 INVX1_LOC_91/A NAND2X1_LOC_793/B 0.01fF
C49230 NOR2X1_LOC_67/a_36_216# INVX1_LOC_46/Y 0.00fF
C49231 NOR2X1_LOC_68/A NAND2X1_LOC_162/A 0.01fF
C49232 INVX1_LOC_214/Y INVX1_LOC_24/A 0.04fF
C49233 INVX1_LOC_21/A NOR2X1_LOC_97/A 0.03fF
C49234 INVX1_LOC_5/A INVX1_LOC_48/A 0.03fF
C49235 INVX1_LOC_27/A NOR2X1_LOC_368/A 0.01fF
C49236 INVX1_LOC_286/Y INVX1_LOC_10/A 9.09fF
C49237 NAND2X1_LOC_733/Y NOR2X1_LOC_525/a_36_216# 0.00fF
C49238 INVX1_LOC_2/A NOR2X1_LOC_753/Y 0.03fF
C49239 INVX1_LOC_217/Y NAND2X1_LOC_562/B -0.01fF
C49240 INVX1_LOC_136/A INVX1_LOC_290/A 0.02fF
C49241 NAND2X1_LOC_794/B NOR2X1_LOC_165/a_36_216# 0.01fF
C49242 INVX1_LOC_36/A NAND2X1_LOC_707/a_36_24# 0.00fF
C49243 INVX1_LOC_21/A INVX1_LOC_193/Y 0.03fF
C49244 NOR2X1_LOC_226/A INVX1_LOC_180/A 0.02fF
C49245 NOR2X1_LOC_464/B NOR2X1_LOC_151/Y 0.01fF
C49246 NOR2X1_LOC_270/Y NAND2X1_LOC_479/Y 0.05fF
C49247 NAND2X1_LOC_357/B NAND2X1_LOC_811/Y 0.02fF
C49248 INVX1_LOC_90/A INVX1_LOC_292/A 0.07fF
C49249 INVX1_LOC_119/A NAND2X1_LOC_326/a_36_24# 0.01fF
C49250 NAND2X1_LOC_722/A NAND2X1_LOC_833/a_36_24# 0.00fF
C49251 NAND2X1_LOC_347/B INPUT_0 0.53fF
C49252 INVX1_LOC_2/A NAND2X1_LOC_325/Y 0.03fF
C49253 INVX1_LOC_111/A INVX1_LOC_22/A 0.02fF
C49254 INVX1_LOC_101/Y NOR2X1_LOC_74/A 0.09fF
C49255 NAND2X1_LOC_276/Y NAND2X1_LOC_338/B 0.07fF
C49256 INVX1_LOC_145/A NAND2X1_LOC_349/B 0.10fF
C49257 NOR2X1_LOC_688/Y INVX1_LOC_89/A 0.02fF
C49258 NOR2X1_LOC_781/A NOR2X1_LOC_781/Y 0.16fF
C49259 NOR2X1_LOC_237/Y INVX1_LOC_25/Y 0.07fF
C49260 INVX1_LOC_256/A INVX1_LOC_73/A 0.00fF
C49261 NOR2X1_LOC_637/A NOR2X1_LOC_561/Y 0.02fF
C49262 NAND2X1_LOC_783/Y NOR2X1_LOC_329/B 0.01fF
C49263 INVX1_LOC_49/Y INVX1_LOC_264/A 0.16fF
C49264 INVX1_LOC_108/A NOR2X1_LOC_227/A 0.18fF
C49265 INVX1_LOC_159/A INVX1_LOC_10/A 0.01fF
C49266 NOR2X1_LOC_98/B NOR2X1_LOC_39/Y 0.01fF
C49267 INVX1_LOC_13/A NOR2X1_LOC_860/B 0.09fF
C49268 NOR2X1_LOC_607/A NOR2X1_LOC_561/Y 0.40fF
C49269 NAND2X1_LOC_773/Y INVX1_LOC_286/A 0.10fF
C49270 NOR2X1_LOC_656/a_36_216# NOR2X1_LOC_332/A 0.01fF
C49271 INVX1_LOC_188/A INVX1_LOC_182/A 0.05fF
C49272 INVX1_LOC_1/A NOR2X1_LOC_334/A 0.02fF
C49273 NOR2X1_LOC_449/a_36_216# NOR2X1_LOC_561/Y 0.01fF
C49274 NOR2X1_LOC_78/B NOR2X1_LOC_718/B 0.02fF
C49275 NOR2X1_LOC_48/Y INVX1_LOC_29/A 0.01fF
C49276 NOR2X1_LOC_191/B INVX1_LOC_10/A 0.72fF
C49277 INVX1_LOC_224/A INVX1_LOC_92/Y 0.00fF
C49278 INVX1_LOC_94/A NAND2X1_LOC_656/Y 0.72fF
C49279 INVX1_LOC_256/Y NAND2X1_LOC_477/A 0.03fF
C49280 INVX1_LOC_24/A NAND2X1_LOC_808/A 0.07fF
C49281 NOR2X1_LOC_690/A NAND2X1_LOC_859/B 0.17fF
C49282 INVX1_LOC_2/Y INVX1_LOC_138/Y 0.03fF
C49283 INVX1_LOC_276/A INVX1_LOC_2/A 0.07fF
C49284 INVX1_LOC_53/A NAND2X1_LOC_472/Y 0.07fF
C49285 NOR2X1_LOC_413/Y NAND2X1_LOC_859/B 0.02fF
C49286 NOR2X1_LOC_197/A INVX1_LOC_311/A 0.03fF
C49287 NOR2X1_LOC_309/Y INVX1_LOC_25/Y 0.10fF
C49288 INVX1_LOC_2/A NOR2X1_LOC_67/A 0.24fF
C49289 INVX1_LOC_276/A NOR2X1_LOC_226/A 0.01fF
C49290 NOR2X1_LOC_590/A NOR2X1_LOC_113/B 0.05fF
C49291 INVX1_LOC_236/A NAND2X1_LOC_840/B 0.18fF
C49292 NAND2X1_LOC_122/a_36_24# INVX1_LOC_16/A 0.00fF
C49293 INVX1_LOC_279/A NOR2X1_LOC_570/B 0.07fF
C49294 INVX1_LOC_222/Y NOR2X1_LOC_567/a_36_216# 0.00fF
C49295 INVX1_LOC_36/A INVX1_LOC_75/A 0.20fF
C49296 INVX1_LOC_30/A INVX1_LOC_282/A 0.05fF
C49297 NOR2X1_LOC_216/B INVX1_LOC_26/A 0.10fF
C49298 NOR2X1_LOC_103/Y INVX1_LOC_91/A 0.17fF
C49299 NAND2X1_LOC_331/a_36_24# INVX1_LOC_49/A 0.00fF
C49300 INVX1_LOC_11/A NOR2X1_LOC_562/B 0.02fF
C49301 INVX1_LOC_313/A NOR2X1_LOC_577/Y 0.01fF
C49302 INVX1_LOC_21/A NAND2X1_LOC_287/B 0.07fF
C49303 INVX1_LOC_102/A NOR2X1_LOC_46/a_36_216# 0.01fF
C49304 NOR2X1_LOC_189/a_36_216# NOR2X1_LOC_48/B 0.00fF
C49305 NOR2X1_LOC_162/Y INVX1_LOC_83/A 0.03fF
C49306 NOR2X1_LOC_570/Y INVX1_LOC_177/A 0.01fF
C49307 INVX1_LOC_58/A INVX1_LOC_185/A 0.05fF
C49308 INVX1_LOC_13/A NAND2X1_LOC_141/A 0.26fF
C49309 NOR2X1_LOC_473/B NOR2X1_LOC_433/A 0.10fF
C49310 VDD NAND2X1_LOC_474/Y 0.33fF
C49311 INVX1_LOC_110/A INPUT_0 0.05fF
C49312 INVX1_LOC_191/Y INVX1_LOC_22/A 0.02fF
C49313 NOR2X1_LOC_391/A NOR2X1_LOC_315/Y 0.01fF
C49314 INVX1_LOC_265/A INVX1_LOC_135/A 0.06fF
C49315 NAND2X1_LOC_728/a_36_24# NAND2X1_LOC_354/B 0.00fF
C49316 INVX1_LOC_50/A NOR2X1_LOC_88/Y 0.03fF
C49317 NOR2X1_LOC_15/Y NOR2X1_LOC_357/Y 0.03fF
C49318 NOR2X1_LOC_247/a_36_216# NAND2X1_LOC_45/Y 0.00fF
C49319 NOR2X1_LOC_424/Y NOR2X1_LOC_423/Y 1.19fF
C49320 NAND2X1_LOC_563/Y D_INPUT_0 0.72fF
C49321 NOR2X1_LOC_586/a_36_216# INVX1_LOC_266/Y 0.00fF
C49322 NOR2X1_LOC_78/B NOR2X1_LOC_569/Y 0.07fF
C49323 INVX1_LOC_53/A NAND2X1_LOC_434/Y 0.01fF
C49324 NOR2X1_LOC_208/Y INVX1_LOC_75/A 0.05fF
C49325 NAND2X1_LOC_866/A NAND2X1_LOC_863/A 0.31fF
C49326 INVX1_LOC_13/A INVX1_LOC_226/A 0.04fF
C49327 NOR2X1_LOC_82/Y INVX1_LOC_53/Y 0.09fF
C49328 NAND2X1_LOC_381/a_36_24# INVX1_LOC_74/A 0.01fF
C49329 INVX1_LOC_45/A INVX1_LOC_91/A 0.44fF
C49330 NOR2X1_LOC_186/Y INVX1_LOC_118/Y 0.02fF
C49331 INVX1_LOC_224/Y NOR2X1_LOC_179/Y 0.06fF
C49332 NOR2X1_LOC_828/B NOR2X1_LOC_712/Y 0.01fF
C49333 INVX1_LOC_272/Y VDD 0.55fF
C49334 NOR2X1_LOC_473/B NOR2X1_LOC_52/B 0.30fF
C49335 NOR2X1_LOC_568/A INVX1_LOC_91/A 0.71fF
C49336 NOR2X1_LOC_424/Y NOR2X1_LOC_222/Y 0.07fF
C49337 INVX1_LOC_50/A INVX1_LOC_84/A 0.09fF
C49338 NOR2X1_LOC_19/B INVX1_LOC_315/A 0.52fF
C49339 NAND2X1_LOC_53/Y VDD -0.00fF
C49340 NAND2X1_LOC_859/Y INVX1_LOC_22/A 0.01fF
C49341 NOR2X1_LOC_136/Y NAND2X1_LOC_656/Y 0.02fF
C49342 NOR2X1_LOC_667/A NOR2X1_LOC_312/Y 0.54fF
C49343 INVX1_LOC_17/A INVX1_LOC_12/Y 0.01fF
C49344 NAND2X1_LOC_765/a_36_24# INVX1_LOC_55/Y 0.01fF
C49345 INVX1_LOC_248/A NOR2X1_LOC_312/Y 0.01fF
C49346 NAND2X1_LOC_842/B NOR2X1_LOC_709/A 0.18fF
C49347 INVX1_LOC_40/A INVX1_LOC_306/A 0.03fF
C49348 INVX1_LOC_55/Y INVX1_LOC_96/Y 0.72fF
C49349 NAND2X1_LOC_573/Y INVX1_LOC_118/Y 0.02fF
C49350 NAND2X1_LOC_856/A INVX1_LOC_11/Y 0.02fF
C49351 INVX1_LOC_13/A NOR2X1_LOC_97/B 0.03fF
C49352 NOR2X1_LOC_657/Y NAND2X1_LOC_468/B 0.00fF
C49353 INVX1_LOC_181/Y NOR2X1_LOC_191/a_36_216# 0.01fF
C49354 INVX1_LOC_25/A INVX1_LOC_293/Y 0.23fF
C49355 NOR2X1_LOC_67/A INPUT_1 0.26fF
C49356 NOR2X1_LOC_577/Y INVX1_LOC_6/A 0.31fF
C49357 INVX1_LOC_223/A NAND2X1_LOC_447/Y 0.01fF
C49358 NOR2X1_LOC_169/a_36_216# NAND2X1_LOC_72/B 0.00fF
C49359 NOR2X1_LOC_778/B INVX1_LOC_196/Y 0.03fF
C49360 INVX1_LOC_49/A NOR2X1_LOC_551/Y 0.05fF
C49361 NOR2X1_LOC_309/Y INVX1_LOC_75/A 0.12fF
C49362 NOR2X1_LOC_224/Y INVX1_LOC_84/A 0.02fF
C49363 INVX1_LOC_1/Y INVX1_LOC_150/A 0.02fF
C49364 NOR2X1_LOC_322/Y NOR2X1_LOC_52/B 0.07fF
C49365 INVX1_LOC_23/A INVX1_LOC_186/Y 0.03fF
C49366 NAND2X1_LOC_342/Y INVX1_LOC_28/A 0.01fF
C49367 INVX1_LOC_103/A INVX1_LOC_38/A 0.15fF
C49368 INVX1_LOC_71/A INVX1_LOC_91/A 0.38fF
C49369 NOR2X1_LOC_220/A NOR2X1_LOC_644/A 0.03fF
C49370 NOR2X1_LOC_392/Y INVX1_LOC_63/A 0.07fF
C49371 NAND2X1_LOC_162/A NOR2X1_LOC_163/A 0.00fF
C49372 NOR2X1_LOC_355/A INVX1_LOC_101/A 0.03fF
C49373 INVX1_LOC_89/A INVX1_LOC_1/Y 0.07fF
C49374 INVX1_LOC_23/A NOR2X1_LOC_777/B 0.37fF
C49375 NOR2X1_LOC_516/B INVX1_LOC_20/Y 0.01fF
C49376 NAND2X1_LOC_866/B INVX1_LOC_22/A 0.10fF
C49377 INVX1_LOC_36/A NAND2X1_LOC_453/A 0.10fF
C49378 INVX1_LOC_25/A NAND2X1_LOC_74/B 1.84fF
C49379 NOR2X1_LOC_840/Y NOR2X1_LOC_833/B 0.00fF
C49380 INVX1_LOC_11/A INVX1_LOC_193/A 0.34fF
C49381 NOR2X1_LOC_790/B INVX1_LOC_19/A 0.10fF
C49382 INVX1_LOC_24/Y NOR2X1_LOC_640/Y 0.13fF
C49383 INVX1_LOC_292/A INVX1_LOC_38/A 0.07fF
C49384 NAND2X1_LOC_303/Y NAND2X1_LOC_802/Y 0.05fF
C49385 NOR2X1_LOC_553/B INVX1_LOC_313/Y 0.03fF
C49386 INVX1_LOC_45/A NOR2X1_LOC_698/Y 0.25fF
C49387 NOR2X1_LOC_798/A INVX1_LOC_294/A 0.00fF
C49388 INVX1_LOC_237/A INVX1_LOC_260/Y 0.30fF
C49389 INVX1_LOC_16/Y NOR2X1_LOC_38/B 0.00fF
C49390 D_INPUT_0 INVX1_LOC_148/Y 0.03fF
C49391 INVX1_LOC_190/Y INVX1_LOC_10/A 0.01fF
C49392 INVX1_LOC_223/Y INVX1_LOC_63/A 0.03fF
C49393 NAND2X1_LOC_778/Y NAND2X1_LOC_489/Y 0.01fF
C49394 NOR2X1_LOC_544/A NOR2X1_LOC_74/A 0.23fF
C49395 NAND2X1_LOC_175/Y INVX1_LOC_273/A 0.03fF
C49396 INVX1_LOC_50/A INVX1_LOC_15/A 0.20fF
C49397 INVX1_LOC_8/A NAND2X1_LOC_642/Y 0.03fF
C49398 NOR2X1_LOC_598/B NOR2X1_LOC_640/B 0.03fF
C49399 NAND2X1_LOC_569/B INVX1_LOC_284/A 0.54fF
C49400 INVX1_LOC_226/Y NOR2X1_LOC_721/Y 0.02fF
C49401 INVX1_LOC_90/A INVX1_LOC_120/A 0.03fF
C49402 INVX1_LOC_77/A NOR2X1_LOC_112/a_36_216# 0.01fF
C49403 NAND2X1_LOC_227/Y NOR2X1_LOC_88/Y 0.02fF
C49404 NOR2X1_LOC_257/a_36_216# INVX1_LOC_117/A 0.01fF
C49405 NOR2X1_LOC_38/B NAND2X1_LOC_205/A 0.01fF
C49406 INVX1_LOC_33/A INVX1_LOC_176/A 0.02fF
C49407 INVX1_LOC_209/Y INVX1_LOC_46/A 0.03fF
C49408 NAND2X1_LOC_538/Y INVX1_LOC_119/Y 0.04fF
C49409 NOR2X1_LOC_15/Y NAND2X1_LOC_489/Y 0.06fF
C49410 INVX1_LOC_31/A NOR2X1_LOC_88/A 0.01fF
C49411 NOR2X1_LOC_103/Y NOR2X1_LOC_179/Y 0.01fF
C49412 NOR2X1_LOC_41/Y NOR2X1_LOC_43/Y 0.03fF
C49413 INVX1_LOC_6/A INVX1_LOC_22/A 2.83fF
C49414 INVX1_LOC_87/A NOR2X1_LOC_748/A 0.04fF
C49415 NOR2X1_LOC_318/B NOR2X1_LOC_524/a_36_216# 0.00fF
C49416 NAND2X1_LOC_227/Y INVX1_LOC_84/A 0.08fF
C49417 NOR2X1_LOC_309/Y NOR2X1_LOC_309/a_36_216# 0.00fF
C49418 NAND2X1_LOC_656/Y INVX1_LOC_144/A 0.02fF
C49419 INVX1_LOC_89/A NOR2X1_LOC_742/A 0.07fF
C49420 NAND2X1_LOC_838/Y NAND2X1_LOC_836/Y 0.17fF
C49421 NOR2X1_LOC_655/B INVX1_LOC_95/Y 0.10fF
C49422 NAND2X1_LOC_111/a_36_24# NOR2X1_LOC_97/B 0.00fF
C49423 INVX1_LOC_233/A NAND2X1_LOC_444/B 0.02fF
C49424 INVX1_LOC_1/A NAND2X1_LOC_74/B 0.11fF
C49425 INVX1_LOC_104/A INVX1_LOC_37/A 0.19fF
C49426 INVX1_LOC_69/Y NOR2X1_LOC_335/a_36_216# 0.01fF
C49427 NOR2X1_LOC_669/Y NOR2X1_LOC_669/A 0.02fF
C49428 NOR2X1_LOC_357/Y INVX1_LOC_96/Y 0.46fF
C49429 NAND2X1_LOC_357/a_36_24# NOR2X1_LOC_743/Y 0.00fF
C49430 NOR2X1_LOC_360/Y NAND2X1_LOC_656/B 0.03fF
C49431 INVX1_LOC_53/A NAND2X1_LOC_70/a_36_24# 0.00fF
C49432 INVX1_LOC_14/A NOR2X1_LOC_847/A 0.07fF
C49433 INVX1_LOC_49/A NOR2X1_LOC_729/A 0.10fF
C49434 INVX1_LOC_1/A NOR2X1_LOC_847/B 0.11fF
C49435 NAND2X1_LOC_392/A INVX1_LOC_304/A 0.01fF
C49436 INVX1_LOC_40/A INVX1_LOC_59/Y 2.08fF
C49437 INVX1_LOC_24/A INVX1_LOC_92/A 7.76fF
C49438 INVX1_LOC_28/A INVX1_LOC_67/Y 0.02fF
C49439 INVX1_LOC_14/A INVX1_LOC_42/A 0.23fF
C49440 NAND2X1_LOC_352/B INVX1_LOC_19/A 0.03fF
C49441 NOR2X1_LOC_226/A NOR2X1_LOC_558/A 0.02fF
C49442 NOR2X1_LOC_667/A NAND2X1_LOC_287/B 0.33fF
C49443 NAND2X1_LOC_795/a_36_24# NAND2X1_LOC_804/Y 0.01fF
C49444 INVX1_LOC_197/A VDD -0.00fF
C49445 NOR2X1_LOC_828/Y NOR2X1_LOC_383/B 0.71fF
C49446 INPUT_0 NOR2X1_LOC_564/Y 0.03fF
C49447 NOR2X1_LOC_318/B INVX1_LOC_150/A 0.03fF
C49448 NOR2X1_LOC_798/A NOR2X1_LOC_334/Y 0.00fF
C49449 INVX1_LOC_240/A INVX1_LOC_38/A 0.03fF
C49450 NAND2X1_LOC_332/Y NOR2X1_LOC_351/Y 0.01fF
C49451 NAND2X1_LOC_363/B NOR2X1_LOC_720/A 0.05fF
C49452 NOR2X1_LOC_123/B INVX1_LOC_91/A 0.10fF
C49453 NOR2X1_LOC_15/Y INVX1_LOC_32/A 0.11fF
C49454 NOR2X1_LOC_530/Y INVX1_LOC_284/A 0.01fF
C49455 INVX1_LOC_75/A NOR2X1_LOC_208/A 0.05fF
C49456 NOR2X1_LOC_500/Y VDD 0.76fF
C49457 INVX1_LOC_278/A INVX1_LOC_50/A 0.00fF
C49458 NOR2X1_LOC_78/B NAND2X1_LOC_472/Y 0.07fF
C49459 INVX1_LOC_305/A NOR2X1_LOC_691/A 0.04fF
C49460 INVX1_LOC_226/Y VDD 1.15fF
C49461 INVX1_LOC_108/Y NOR2X1_LOC_105/Y 0.04fF
C49462 INVX1_LOC_20/Y INVX1_LOC_315/Y 0.01fF
C49463 NOR2X1_LOC_446/A INVX1_LOC_290/Y 0.03fF
C49464 INVX1_LOC_41/A NOR2X1_LOC_640/Y 0.08fF
C49465 NAND2X1_LOC_573/a_36_24# NAND2X1_LOC_288/A 0.01fF
C49466 INVX1_LOC_10/A NOR2X1_LOC_56/Y 1.91fF
C49467 NOR2X1_LOC_78/A INVX1_LOC_65/Y 0.01fF
C49468 NOR2X1_LOC_557/Y INVX1_LOC_92/A 0.07fF
C49469 NOR2X1_LOC_667/A NAND2X1_LOC_808/a_36_24# 0.00fF
C49470 NOR2X1_LOC_653/B NOR2X1_LOC_301/A 0.01fF
C49471 INVX1_LOC_25/A NOR2X1_LOC_660/Y 0.06fF
C49472 INVX1_LOC_286/Y INVX1_LOC_12/A 8.07fF
C49473 INVX1_LOC_89/A INVX1_LOC_93/Y 0.09fF
C49474 NAND2X1_LOC_182/A NOR2X1_LOC_177/Y 0.02fF
C49475 INVX1_LOC_63/Y INVX1_LOC_179/A 0.01fF
C49476 NOR2X1_LOC_360/Y NOR2X1_LOC_721/B 0.00fF
C49477 INVX1_LOC_5/A NOR2X1_LOC_383/B 0.10fF
C49478 NOR2X1_LOC_632/Y INVX1_LOC_14/Y 0.05fF
C49479 NAND2X1_LOC_181/Y NOR2X1_LOC_536/A 0.01fF
C49480 INVX1_LOC_204/A INVX1_LOC_204/Y 0.09fF
C49481 INVX1_LOC_104/A NOR2X1_LOC_743/Y 0.28fF
C49482 INVX1_LOC_276/A INVX1_LOC_118/A 0.10fF
C49483 NOR2X1_LOC_432/a_36_216# INVX1_LOC_54/A 0.00fF
C49484 NOR2X1_LOC_384/Y NAND2X1_LOC_74/B 0.04fF
C49485 INVX1_LOC_25/Y NOR2X1_LOC_102/a_36_216# 0.00fF
C49486 INVX1_LOC_88/Y NOR2X1_LOC_155/A 0.03fF
C49487 INVX1_LOC_269/A INVX1_LOC_94/Y 0.08fF
C49488 INVX1_LOC_35/A INVX1_LOC_58/Y 0.01fF
C49489 NAND2X1_LOC_555/Y NOR2X1_LOC_554/A 0.06fF
C49490 INVX1_LOC_10/A VDD 1.03fF
C49491 NOR2X1_LOC_15/Y NAND2X1_LOC_175/Y 0.09fF
C49492 INVX1_LOC_14/A INVX1_LOC_78/A 0.30fF
C49493 NOR2X1_LOC_205/Y NAND2X1_LOC_454/Y 0.07fF
C49494 NOR2X1_LOC_91/Y INVX1_LOC_29/A 0.10fF
C49495 INVX1_LOC_10/A NAND2X1_LOC_800/A 0.03fF
C49496 INVX1_LOC_100/A INVX1_LOC_6/A 0.01fF
C49497 NAND2X1_LOC_390/A NOR2X1_LOC_536/A 0.05fF
C49498 INVX1_LOC_45/A NOR2X1_LOC_483/a_36_216# 0.02fF
C49499 INVX1_LOC_159/A INVX1_LOC_12/A 0.01fF
C49500 INVX1_LOC_33/Y NAND2X1_LOC_796/Y 0.01fF
C49501 NOR2X1_LOC_457/B NOR2X1_LOC_89/A 0.07fF
C49502 INVX1_LOC_54/Y NOR2X1_LOC_79/Y 0.00fF
C49503 NOR2X1_LOC_623/a_36_216# NOR2X1_LOC_814/A 0.01fF
C49504 INVX1_LOC_143/A INVX1_LOC_92/A 0.07fF
C49505 NAND2X1_LOC_116/a_36_24# INVX1_LOC_9/A 0.00fF
C49506 NOR2X1_LOC_558/A INPUT_1 0.01fF
C49507 NOR2X1_LOC_65/B INVX1_LOC_14/A 0.04fF
C49508 INVX1_LOC_89/A NAND2X1_LOC_721/A 0.02fF
C49509 INVX1_LOC_134/A NOR2X1_LOC_856/a_36_216# 0.00fF
C49510 NOR2X1_LOC_174/A NOR2X1_LOC_857/A 0.03fF
C49511 NAND2X1_LOC_357/B NOR2X1_LOC_653/Y 0.05fF
C49512 INVX1_LOC_57/A NOR2X1_LOC_271/B 0.02fF
C49513 NOR2X1_LOC_320/a_36_216# INVX1_LOC_63/A 0.01fF
C49514 NOR2X1_LOC_344/A INVX1_LOC_19/A 0.01fF
C49515 INVX1_LOC_81/A INVX1_LOC_109/Y 0.08fF
C49516 NOR2X1_LOC_91/A NAND2X1_LOC_799/A 0.08fF
C49517 NOR2X1_LOC_468/Y NAND2X1_LOC_205/A 0.03fF
C49518 NOR2X1_LOC_614/Y NOR2X1_LOC_862/B 0.05fF
C49519 NAND2X1_LOC_764/a_36_24# NOR2X1_LOC_467/A 0.00fF
C49520 VDD NOR2X1_LOC_302/Y 0.12fF
C49521 NAND2X1_LOC_541/Y INVX1_LOC_123/Y 0.01fF
C49522 INVX1_LOC_283/Y INVX1_LOC_12/A 0.03fF
C49523 INVX1_LOC_279/A INVX1_LOC_54/A 0.07fF
C49524 NOR2X1_LOC_208/Y INVX1_LOC_283/A 0.01fF
C49525 NOR2X1_LOC_785/A INVX1_LOC_26/Y 0.00fF
C49526 INVX1_LOC_13/Y INVX1_LOC_306/Y 0.20fF
C49527 INVX1_LOC_120/A INVX1_LOC_38/A 0.08fF
C49528 INVX1_LOC_259/Y INVX1_LOC_1/A 0.01fF
C49529 NAND2X1_LOC_357/B INVX1_LOC_19/A 0.07fF
C49530 NAND2X1_LOC_833/Y NOR2X1_LOC_89/A 0.07fF
C49531 NAND2X1_LOC_690/a_36_24# NOR2X1_LOC_691/A 0.00fF
C49532 NAND2X1_LOC_859/Y NOR2X1_LOC_88/A 0.13fF
C49533 INVX1_LOC_83/A NAND2X1_LOC_637/Y 0.40fF
C49534 INVX1_LOC_1/A NOR2X1_LOC_660/Y 0.86fF
C49535 NOR2X1_LOC_68/A INVX1_LOC_4/Y 0.19fF
C49536 INVX1_LOC_21/A INVX1_LOC_50/Y 0.00fF
C49537 INVX1_LOC_31/A NOR2X1_LOC_843/B 0.11fF
C49538 INVX1_LOC_206/Y NOR2X1_LOC_631/B 0.00fF
C49539 NOR2X1_LOC_561/Y NAND2X1_LOC_798/B 0.07fF
C49540 INVX1_LOC_227/Y INVX1_LOC_78/A 0.08fF
C49541 INVX1_LOC_217/Y INVX1_LOC_42/A 0.00fF
C49542 INVX1_LOC_236/A INVX1_LOC_49/Y 0.25fF
C49543 NOR2X1_LOC_80/a_36_216# NOR2X1_LOC_78/A 0.00fF
C49544 INVX1_LOC_16/A INVX1_LOC_285/A 0.12fF
C49545 INVX1_LOC_33/A NOR2X1_LOC_116/a_36_216# 0.00fF
C49546 NOR2X1_LOC_78/B NAND2X1_LOC_773/B 0.21fF
C49547 NAND2X1_LOC_656/Y NOR2X1_LOC_155/A 0.07fF
C49548 NOR2X1_LOC_537/Y INVX1_LOC_125/A 0.07fF
C49549 NOR2X1_LOC_218/A NOR2X1_LOC_678/A 0.09fF
C49550 NOR2X1_LOC_160/B NAND2X1_LOC_203/a_36_24# 0.00fF
C49551 INVX1_LOC_16/A NOR2X1_LOC_814/A 0.03fF
C49552 INVX1_LOC_25/Y INVX1_LOC_63/A 0.07fF
C49553 INVX1_LOC_191/Y INVX1_LOC_261/A 0.01fF
C49554 INVX1_LOC_234/A INVX1_LOC_260/Y 0.11fF
C49555 NOR2X1_LOC_34/A NAND2X1_LOC_32/a_36_24# 0.02fF
C49556 INVX1_LOC_89/A INVX1_LOC_117/Y 0.12fF
C49557 NOR2X1_LOC_91/A INVX1_LOC_18/A 0.03fF
C49558 INVX1_LOC_51/A NAND2X1_LOC_114/B 0.01fF
C49559 INVX1_LOC_21/A INVX1_LOC_266/A 0.47fF
C49560 NOR2X1_LOC_15/Y INVX1_LOC_171/Y 0.01fF
C49561 NOR2X1_LOC_91/A NAND2X1_LOC_728/Y 0.26fF
C49562 INVX1_LOC_111/Y INVX1_LOC_42/A 0.01fF
C49563 INVX1_LOC_182/Y INVX1_LOC_54/A 0.02fF
C49564 NOR2X1_LOC_510/Y INVX1_LOC_272/Y 0.02fF
C49565 INVX1_LOC_62/Y NOR2X1_LOC_39/Y 0.03fF
C49566 INVX1_LOC_110/Y INVX1_LOC_64/A 0.18fF
C49567 NOR2X1_LOC_196/Y INVX1_LOC_9/A 0.23fF
C49568 NOR2X1_LOC_361/B NAND2X1_LOC_474/Y 0.46fF
C49569 INVX1_LOC_256/Y INVX1_LOC_168/Y 0.04fF
C49570 NOR2X1_LOC_91/A NAND2X1_LOC_711/B 0.01fF
C49571 INVX1_LOC_25/A INVX1_LOC_136/A 0.14fF
C49572 INVX1_LOC_50/A NOR2X1_LOC_168/Y 0.01fF
C49573 NOR2X1_LOC_294/Y NOR2X1_LOC_598/B 0.10fF
C49574 INVX1_LOC_22/A NOR2X1_LOC_633/A 0.00fF
C49575 NAND2X1_LOC_364/A INVX1_LOC_29/Y 0.03fF
C49576 NAND2X1_LOC_141/A INVX1_LOC_32/A 0.52fF
C49577 INVX1_LOC_77/A INVX1_LOC_23/Y 0.07fF
C49578 INVX1_LOC_18/A INVX1_LOC_23/A 0.17fF
C49579 INVX1_LOC_230/Y NAND2X1_LOC_214/B 0.36fF
C49580 NOR2X1_LOC_65/B NAND2X1_LOC_84/Y 0.24fF
C49581 INVX1_LOC_96/Y INVX1_LOC_32/A 0.07fF
C49582 NOR2X1_LOC_600/Y INVX1_LOC_37/A 0.01fF
C49583 NAND2X1_LOC_763/B INPUT_6 0.01fF
C49584 INVX1_LOC_34/A NOR2X1_LOC_158/Y 0.02fF
C49585 INVX1_LOC_41/A NAND2X1_LOC_221/a_36_24# 0.00fF
C49586 NOR2X1_LOC_711/Y VDD 0.00fF
C49587 NOR2X1_LOC_91/A INVX1_LOC_172/A 0.03fF
C49588 INVX1_LOC_90/A NAND2X1_LOC_659/A 0.01fF
C49589 INVX1_LOC_64/A NOR2X1_LOC_382/Y 0.05fF
C49590 NAND2X1_LOC_624/B INVX1_LOC_30/A 0.02fF
C49591 NOR2X1_LOC_78/A NOR2X1_LOC_317/a_36_216# 0.00fF
C49592 NOR2X1_LOC_799/B VDD 0.26fF
C49593 NOR2X1_LOC_211/Y INVX1_LOC_30/A 0.04fF
C49594 NOR2X1_LOC_543/A INVX1_LOC_29/A 0.01fF
C49595 INVX1_LOC_34/A NOR2X1_LOC_25/Y 0.03fF
C49596 INVX1_LOC_104/A NAND2X1_LOC_72/B 0.03fF
C49597 INVX1_LOC_178/Y NAND2X1_LOC_659/B 0.01fF
C49598 NOR2X1_LOC_211/a_36_216# NOR2X1_LOC_360/Y 0.01fF
C49599 INVX1_LOC_57/Y NAND2X1_LOC_552/A 0.05fF
C49600 NOR2X1_LOC_637/Y INVX1_LOC_23/A 0.03fF
C49601 NOR2X1_LOC_577/Y INVX1_LOC_270/A 0.10fF
C49602 NOR2X1_LOC_84/A INVX1_LOC_26/A 0.74fF
C49603 INVX1_LOC_24/A INVX1_LOC_53/A 5.71fF
C49604 NOR2X1_LOC_331/B INVX1_LOC_91/A 0.07fF
C49605 NOR2X1_LOC_598/B NOR2X1_LOC_546/B 0.02fF
C49606 NAND2X1_LOC_787/A INVX1_LOC_41/Y 0.00fF
C49607 INVX1_LOC_1/A NOR2X1_LOC_307/A 0.06fF
C49608 INVX1_LOC_94/A NOR2X1_LOC_717/A 0.29fF
C49609 INVX1_LOC_172/A INVX1_LOC_23/A 0.00fF
C49610 INVX1_LOC_64/A NAND2X1_LOC_521/a_36_24# 0.00fF
C49611 NAND2X1_LOC_721/A NAND2X1_LOC_244/A 0.03fF
C49612 INVX1_LOC_178/Y VDD 0.41fF
C49613 INVX1_LOC_224/Y NAND2X1_LOC_276/Y 0.03fF
C49614 INVX1_LOC_34/A NOR2X1_LOC_646/B 0.03fF
C49615 NAND2X1_LOC_231/Y NOR2X1_LOC_158/Y 0.03fF
C49616 NOR2X1_LOC_792/B NAND2X1_LOC_286/B 0.02fF
C49617 INVX1_LOC_267/A INVX1_LOC_175/A 0.01fF
C49618 INVX1_LOC_309/A NOR2X1_LOC_491/Y 0.01fF
C49619 INVX1_LOC_17/A NAND2X1_LOC_550/A 0.07fF
C49620 NOR2X1_LOC_446/a_36_216# NAND2X1_LOC_190/Y 0.00fF
C49621 INVX1_LOC_78/Y NOR2X1_LOC_155/A 0.05fF
C49622 NOR2X1_LOC_598/B INVX1_LOC_275/A 0.01fF
C49623 NOR2X1_LOC_76/A NOR2X1_LOC_89/A 0.08fF
C49624 INVX1_LOC_35/A NOR2X1_LOC_537/A 0.04fF
C49625 INVX1_LOC_17/A NOR2X1_LOC_160/B 0.11fF
C49626 NAND2X1_LOC_472/Y INVX1_LOC_46/A 0.07fF
C49627 INVX1_LOC_190/Y INVX1_LOC_12/A 0.10fF
C49628 INVX1_LOC_75/A INVX1_LOC_63/A 12.69fF
C49629 NAND2X1_LOC_186/a_36_24# INVX1_LOC_12/A 0.00fF
C49630 INVX1_LOC_200/A NOR2X1_LOC_369/Y 0.04fF
C49631 INVX1_LOC_35/A NOR2X1_LOC_716/B 0.07fF
C49632 NOR2X1_LOC_561/Y INVX1_LOC_47/Y 0.63fF
C49633 NOR2X1_LOC_577/a_36_216# INVX1_LOC_4/A 0.01fF
C49634 NAND2X1_LOC_840/B NAND2X1_LOC_175/Y 0.09fF
C49635 NOR2X1_LOC_337/Y NOR2X1_LOC_445/B 0.00fF
C49636 NOR2X1_LOC_577/Y NOR2X1_LOC_109/Y 0.07fF
C49637 INVX1_LOC_58/A NOR2X1_LOC_310/Y 0.08fF
C49638 INVX1_LOC_91/A NOR2X1_LOC_592/B 0.06fF
C49639 VDD INVX1_LOC_114/A 0.12fF
C49640 INVX1_LOC_5/A NAND2X1_LOC_632/B 0.03fF
C49641 NOR2X1_LOC_689/A NOR2X1_LOC_773/Y 0.06fF
C49642 INVX1_LOC_136/A INVX1_LOC_1/A 0.54fF
C49643 INVX1_LOC_200/A INVX1_LOC_286/Y -0.00fF
C49644 NOR2X1_LOC_836/B NOR2X1_LOC_865/Y 0.13fF
C49645 INVX1_LOC_45/A NOR2X1_LOC_739/Y 0.02fF
C49646 INVX1_LOC_6/A NAND2X1_LOC_476/Y 0.03fF
C49647 NOR2X1_LOC_166/a_36_216# NOR2X1_LOC_48/B 0.00fF
C49648 NAND2X1_LOC_555/Y NOR2X1_LOC_160/B 0.07fF
C49649 INVX1_LOC_14/A NOR2X1_LOC_554/B 0.14fF
C49650 INVX1_LOC_11/Y NOR2X1_LOC_491/Y 0.06fF
C49651 NOR2X1_LOC_536/A INVX1_LOC_117/A 0.07fF
C49652 NOR2X1_LOC_589/A NOR2X1_LOC_278/Y 0.07fF
C49653 INVX1_LOC_73/A NOR2X1_LOC_89/A 0.01fF
C49654 NOR2X1_LOC_772/B INVX1_LOC_294/Y 0.18fF
C49655 INVX1_LOC_6/A INVX1_LOC_186/Y 0.08fF
C49656 NOR2X1_LOC_598/B NOR2X1_LOC_168/B 0.44fF
C49657 NAND2X1_LOC_579/A NOR2X1_LOC_238/Y 0.03fF
C49658 NOR2X1_LOC_346/B NOR2X1_LOC_416/A 0.08fF
C49659 NOR2X1_LOC_188/A NAND2X1_LOC_74/B 0.23fF
C49660 NAND2X1_LOC_733/Y INVX1_LOC_286/Y 0.50fF
C49661 NOR2X1_LOC_548/B NAND2X1_LOC_74/B 0.03fF
C49662 NOR2X1_LOC_435/A NAND2X1_LOC_453/A 0.27fF
C49663 NOR2X1_LOC_91/A NOR2X1_LOC_690/Y 0.03fF
C49664 NOR2X1_LOC_391/A NAND2X1_LOC_99/A 0.07fF
C49665 NAND2X1_LOC_652/Y INVX1_LOC_15/A 1.14fF
C49666 NOR2X1_LOC_576/B NAND2X1_LOC_175/Y 0.53fF
C49667 INVX1_LOC_89/A INVX1_LOC_87/A 0.05fF
C49668 NAND2X1_LOC_9/Y INVX1_LOC_218/A 0.08fF
C49669 NAND2X1_LOC_561/B NOR2X1_LOC_625/Y 0.08fF
C49670 INVX1_LOC_168/A INVX1_LOC_306/Y 0.03fF
C49671 NOR2X1_LOC_647/Y INVX1_LOC_31/A 0.01fF
C49672 NAND2X1_LOC_803/B NOR2X1_LOC_744/Y 0.08fF
C49673 INVX1_LOC_21/A NOR2X1_LOC_6/B 3.34fF
C49674 NOR2X1_LOC_816/A NOR2X1_LOC_512/Y 0.02fF
C49675 VDD NOR2X1_LOC_445/B 0.63fF
C49676 INVX1_LOC_89/A INVX1_LOC_175/A 0.05fF
C49677 NAND2X1_LOC_858/B NOR2X1_LOC_48/B 0.02fF
C49678 INVX1_LOC_31/A INVX1_LOC_18/A 0.32fF
C49679 NAND2X1_LOC_93/B INVX1_LOC_117/A 0.12fF
C49680 NOR2X1_LOC_636/B INVX1_LOC_77/A 0.46fF
C49681 NOR2X1_LOC_272/Y NOR2X1_LOC_361/Y 0.15fF
C49682 NOR2X1_LOC_286/Y INVX1_LOC_49/A 2.81fF
C49683 INVX1_LOC_48/A INVX1_LOC_42/A 0.23fF
C49684 INVX1_LOC_78/Y NOR2X1_LOC_833/B 0.00fF
C49685 INVX1_LOC_30/A INVX1_LOC_142/A 0.10fF
C49686 NOR2X1_LOC_35/Y NOR2X1_LOC_814/A 0.12fF
C49687 NAND2X1_LOC_190/Y NOR2X1_LOC_570/B 0.03fF
C49688 INVX1_LOC_103/A INVX1_LOC_33/A 0.12fF
C49689 NOR2X1_LOC_590/A NOR2X1_LOC_744/Y 0.01fF
C49690 NOR2X1_LOC_43/Y NAND2X1_LOC_74/B 0.03fF
C49691 NAND2X1_LOC_656/Y NOR2X1_LOC_125/Y 0.03fF
C49692 NAND2X1_LOC_597/a_36_24# NOR2X1_LOC_596/A 0.00fF
C49693 INVX1_LOC_11/A NAND2X1_LOC_833/Y 0.03fF
C49694 INVX1_LOC_136/A NOR2X1_LOC_384/Y 0.26fF
C49695 INVX1_LOC_22/A NOR2X1_LOC_109/Y 0.00fF
C49696 NOR2X1_LOC_67/A INVX1_LOC_39/A 0.03fF
C49697 NAND2X1_LOC_276/Y NOR2X1_LOC_103/Y 0.08fF
C49698 NAND2X1_LOC_53/Y INVX1_LOC_153/Y 0.10fF
C49699 NAND2X1_LOC_453/A INVX1_LOC_63/A 0.09fF
C49700 INVX1_LOC_144/A INVX1_LOC_128/Y 0.10fF
C49701 INVX1_LOC_269/A NOR2X1_LOC_315/Y 0.01fF
C49702 INVX1_LOC_103/A NAND2X1_LOC_466/A 0.02fF
C49703 INVX1_LOC_30/A INVX1_LOC_41/Y 0.06fF
C49704 INVX1_LOC_12/A NOR2X1_LOC_56/Y 2.90fF
C49705 INVX1_LOC_292/A INVX1_LOC_33/A 0.07fF
C49706 NOR2X1_LOC_130/A INVX1_LOC_53/A 0.04fF
C49707 INVX1_LOC_200/A INVX1_LOC_185/Y 0.24fF
C49708 INVX1_LOC_117/A INVX1_LOC_3/A 0.08fF
C49709 INVX1_LOC_46/A NAND2X1_LOC_773/B 0.01fF
C49710 NOR2X1_LOC_617/Y INVX1_LOC_30/A 0.16fF
C49711 NAND2X1_LOC_53/Y INVX1_LOC_121/Y 0.01fF
C49712 NAND2X1_LOC_355/Y INVX1_LOC_159/A 0.00fF
C49713 NAND2X1_LOC_105/a_36_24# INVX1_LOC_23/A 0.00fF
C49714 INVX1_LOC_35/A NOR2X1_LOC_717/B 0.03fF
C49715 NAND2X1_LOC_773/Y NOR2X1_LOC_655/B 0.03fF
C49716 NOR2X1_LOC_155/A NOR2X1_LOC_680/a_36_216# 0.00fF
C49717 INVX1_LOC_75/A NAND2X1_LOC_223/B 0.09fF
C49718 NAND2X1_LOC_341/A INVX1_LOC_27/A 0.03fF
C49719 INVX1_LOC_30/A NAND2X1_LOC_593/Y 0.02fF
C49720 INVX1_LOC_18/A INVX1_LOC_111/A 0.01fF
C49721 NOR2X1_LOC_598/B INVX1_LOC_132/Y 0.03fF
C49722 INVX1_LOC_178/A NAND2X1_LOC_170/A 0.05fF
C49723 INVX1_LOC_17/Y NOR2X1_LOC_497/Y 0.05fF
C49724 NOR2X1_LOC_599/A NOR2X1_LOC_387/Y 0.01fF
C49725 NOR2X1_LOC_717/Y INVX1_LOC_113/Y 0.00fF
C49726 INVX1_LOC_35/A NAND2X1_LOC_656/a_36_24# 0.00fF
C49727 NAND2X1_LOC_52/a_36_24# INVX1_LOC_9/A 0.01fF
C49728 NOR2X1_LOC_89/A NAND2X1_LOC_241/Y 0.03fF
C49729 INVX1_LOC_230/Y NOR2X1_LOC_664/Y 0.21fF
C49730 NAND2X1_LOC_447/Y INVX1_LOC_290/Y 0.14fF
C49731 INVX1_LOC_36/A NOR2X1_LOC_577/Y 1.31fF
C49732 INVX1_LOC_1/A NAND2X1_LOC_304/a_36_24# 0.00fF
C49733 INVX1_LOC_304/Y NOR2X1_LOC_369/Y 0.05fF
C49734 VDD INVX1_LOC_12/A 2.01fF
C49735 NOR2X1_LOC_251/a_36_216# INVX1_LOC_53/Y -0.02fF
C49736 NOR2X1_LOC_185/a_36_216# NOR2X1_LOC_668/Y 0.01fF
C49737 INVX1_LOC_35/A NOR2X1_LOC_828/A 0.03fF
C49738 NOR2X1_LOC_631/A INVX1_LOC_38/A 0.45fF
C49739 INVX1_LOC_103/A NAND2X1_LOC_798/A 0.03fF
C49740 NOR2X1_LOC_510/Y INVX1_LOC_10/A 0.02fF
C49741 VDD NOR2X1_LOC_519/Y 0.23fF
C49742 NAND2X1_LOC_557/Y NAND2X1_LOC_849/A 0.01fF
C49743 NAND2X1_LOC_800/A INVX1_LOC_12/A 0.08fF
C49744 NOR2X1_LOC_471/Y INVX1_LOC_189/A -0.03fF
C49745 NAND2X1_LOC_573/A NAND2X1_LOC_474/Y 0.26fF
C49746 NOR2X1_LOC_15/Y NAND2X1_LOC_564/B 0.07fF
C49747 INVX1_LOC_226/Y NOR2X1_LOC_361/B 0.10fF
C49748 NAND2X1_LOC_739/B NOR2X1_LOC_152/Y 0.04fF
C49749 NOR2X1_LOC_176/a_36_216# INVX1_LOC_102/A 0.00fF
C49750 INVX1_LOC_224/Y NOR2X1_LOC_184/a_36_216# 0.01fF
C49751 INVX1_LOC_17/A INVX1_LOC_208/A 0.04fF
C49752 INVX1_LOC_256/A NAND2X1_LOC_181/Y 0.00fF
C49753 NOR2X1_LOC_388/Y NOR2X1_LOC_703/B 0.04fF
C49754 INVX1_LOC_181/Y INVX1_LOC_49/A 0.03fF
C49755 NOR2X1_LOC_272/Y NOR2X1_LOC_355/A 0.03fF
C49756 NOR2X1_LOC_216/Y INVX1_LOC_53/A 0.07fF
C49757 NOR2X1_LOC_457/B NOR2X1_LOC_593/Y 0.07fF
C49758 INVX1_LOC_17/A NOR2X1_LOC_516/B 0.12fF
C49759 NOR2X1_LOC_411/Y INVX1_LOC_207/Y 0.24fF
C49760 INVX1_LOC_31/A INVX1_LOC_34/Y 0.15fF
C49761 NOR2X1_LOC_65/B INVX1_LOC_48/A -0.10fF
C49762 NOR2X1_LOC_567/B NOR2X1_LOC_634/Y 0.09fF
C49763 INVX1_LOC_34/A NOR2X1_LOC_759/A 0.09fF
C49764 NOR2X1_LOC_309/Y NOR2X1_LOC_274/B 0.19fF
C49765 NOR2X1_LOC_843/A NOR2X1_LOC_68/A 0.52fF
C49766 NOR2X1_LOC_548/A INVX1_LOC_23/A 0.15fF
C49767 INVX1_LOC_35/A NOR2X1_LOC_151/Y 0.07fF
C49768 INVX1_LOC_250/A NOR2X1_LOC_591/Y 0.01fF
C49769 INVX1_LOC_312/Y NAND2X1_LOC_660/A 0.03fF
C49770 INVX1_LOC_247/A NOR2X1_LOC_465/Y 0.25fF
C49771 INVX1_LOC_88/A NOR2X1_LOC_171/a_36_216# 0.00fF
C49772 NOR2X1_LOC_816/A NAND2X1_LOC_170/A 0.04fF
C49773 NOR2X1_LOC_615/Y INVX1_LOC_16/A 0.02fF
C49774 INVX1_LOC_11/A NOR2X1_LOC_781/A 0.07fF
C49775 INVX1_LOC_72/A NOR2X1_LOC_709/A 2.54fF
C49776 NOR2X1_LOC_252/Y NAND2X1_LOC_550/A 0.04fF
C49777 NOR2X1_LOC_751/Y NOR2X1_LOC_175/A 0.00fF
C49778 INVX1_LOC_278/Y NAND2X1_LOC_711/Y 0.00fF
C49779 NAND2X1_LOC_754/a_36_24# INVX1_LOC_292/A 0.00fF
C49780 INVX1_LOC_269/A INVX1_LOC_66/A 0.11fF
C49781 NOR2X1_LOC_210/A INVX1_LOC_174/A 0.02fF
C49782 NOR2X1_LOC_590/A INVX1_LOC_16/A 0.03fF
C49783 NAND2X1_LOC_787/B NAND2X1_LOC_486/a_36_24# 0.00fF
C49784 NOR2X1_LOC_273/Y NOR2X1_LOC_300/Y 0.02fF
C49785 INVX1_LOC_41/A NOR2X1_LOC_730/a_36_216# 0.00fF
C49786 NOR2X1_LOC_584/Y INVX1_LOC_118/A 0.03fF
C49787 NOR2X1_LOC_772/B NOR2X1_LOC_74/A 0.17fF
C49788 INVX1_LOC_57/Y NOR2X1_LOC_773/Y 0.02fF
C49789 NOR2X1_LOC_598/B INVX1_LOC_78/Y 0.03fF
C49790 NOR2X1_LOC_536/A INVX1_LOC_3/Y 0.01fF
C49791 INVX1_LOC_269/A NAND2X1_LOC_624/A 0.00fF
C49792 NOR2X1_LOC_278/Y INVX1_LOC_20/A 0.48fF
C49793 NAND2X1_LOC_722/A INVX1_LOC_41/Y 0.07fF
C49794 NOR2X1_LOC_67/A INVX1_LOC_61/A 0.08fF
C49795 INVX1_LOC_13/Y NOR2X1_LOC_74/A 0.10fF
C49796 NOR2X1_LOC_763/A INVX1_LOC_140/A 0.10fF
C49797 NOR2X1_LOC_364/A INVX1_LOC_109/A 0.01fF
C49798 NAND2X1_LOC_562/B NAND2X1_LOC_632/B 0.04fF
C49799 INVX1_LOC_230/Y INVX1_LOC_234/A 0.56fF
C49800 NOR2X1_LOC_405/A INVX1_LOC_29/Y 0.11fF
C49801 INVX1_LOC_149/A NOR2X1_LOC_303/Y 0.10fF
C49802 INVX1_LOC_12/Y INVX1_LOC_94/Y 0.03fF
C49803 NOR2X1_LOC_582/A INVX1_LOC_140/A 0.01fF
C49804 INVX1_LOC_36/A INVX1_LOC_22/A 4.48fF
C49805 NOR2X1_LOC_82/A INVX1_LOC_89/A 0.15fF
C49806 NOR2X1_LOC_226/A INVX1_LOC_181/Y 0.00fF
C49807 NAND2X1_LOC_861/a_36_24# INVX1_LOC_30/A 0.06fF
C49808 INVX1_LOC_311/A INVX1_LOC_50/Y 0.06fF
C49809 NOR2X1_LOC_78/B INVX1_LOC_24/A 0.31fF
C49810 NOR2X1_LOC_637/Y INVX1_LOC_191/Y 0.00fF
C49811 INVX1_LOC_279/A NOR2X1_LOC_441/Y 0.07fF
C49812 INVX1_LOC_184/A INVX1_LOC_143/A 0.03fF
C49813 VDD NOR2X1_LOC_686/A 0.00fF
C49814 INVX1_LOC_284/Y INVX1_LOC_229/Y 0.10fF
C49815 INVX1_LOC_11/A NOR2X1_LOC_180/B 0.07fF
C49816 INVX1_LOC_71/A NOR2X1_LOC_352/Y 0.05fF
C49817 INVX1_LOC_13/Y NOR2X1_LOC_9/Y 0.07fF
C49818 NOR2X1_LOC_655/Y INVX1_LOC_3/Y 0.01fF
C49819 NOR2X1_LOC_45/B NOR2X1_LOC_53/Y 0.01fF
C49820 NOR2X1_LOC_284/B INVX1_LOC_77/A 0.04fF
C49821 INVX1_LOC_286/Y NAND2X1_LOC_808/A 0.01fF
C49822 NAND2X1_LOC_859/Y INVX1_LOC_18/A 0.10fF
C49823 NOR2X1_LOC_815/Y INVX1_LOC_276/A 0.02fF
C49824 NAND2X1_LOC_803/B INVX1_LOC_28/A 0.96fF
C49825 NAND2X1_LOC_425/Y NOR2X1_LOC_460/A -0.00fF
C49826 INVX1_LOC_209/Y NOR2X1_LOC_505/Y 0.11fF
C49827 NOR2X1_LOC_208/Y INVX1_LOC_22/A 0.07fF
C49828 NAND2X1_LOC_36/A INVX1_LOC_89/A 0.02fF
C49829 INVX1_LOC_21/A INVX1_LOC_96/A 0.03fF
C49830 NOR2X1_LOC_590/A INVX1_LOC_28/A 0.07fF
C49831 INVX1_LOC_230/Y NOR2X1_LOC_19/B 1.14fF
C49832 INVX1_LOC_135/A NOR2X1_LOC_703/B 0.05fF
C49833 NOR2X1_LOC_220/A NOR2X1_LOC_570/B 0.30fF
C49834 NOR2X1_LOC_326/Y NOR2X1_LOC_325/Y 0.08fF
C49835 NOR2X1_LOC_468/Y INVX1_LOC_286/A 1.58fF
C49836 NOR2X1_LOC_613/Y NOR2X1_LOC_45/B 0.01fF
C49837 NAND2X1_LOC_82/Y INVX1_LOC_29/A 0.07fF
C49838 INVX1_LOC_35/A NAND2X1_LOC_633/Y 0.07fF
C49839 NOR2X1_LOC_356/A NOR2X1_LOC_500/B 0.00fF
C49840 INVX1_LOC_54/Y INVX1_LOC_149/A 0.57fF
C49841 INVX1_LOC_24/A INVX1_LOC_83/A 0.17fF
C49842 NAND2X1_LOC_338/B NOR2X1_LOC_709/A 0.17fF
C49843 NOR2X1_LOC_649/B INVX1_LOC_3/Y 0.07fF
C49844 INVX1_LOC_31/A INVX1_LOC_31/Y 0.04fF
C49845 INVX1_LOC_217/Y NAND2X1_LOC_859/B 0.00fF
C49846 NAND2X1_LOC_53/Y INVX1_LOC_285/Y 0.08fF
C49847 NAND2X1_LOC_63/Y NOR2X1_LOC_327/a_36_216# 0.00fF
C49848 NAND2X1_LOC_721/A NOR2X1_LOC_392/Y 0.01fF
C49849 INVX1_LOC_3/A INVX1_LOC_3/Y 6.25fF
C49850 INVX1_LOC_58/A NOR2X1_LOC_536/A 2.27fF
C49851 INVX1_LOC_158/A INVX1_LOC_226/A 0.00fF
C49852 NAND2X1_LOC_795/a_36_24# NOR2X1_LOC_667/A 0.00fF
C49853 INVX1_LOC_13/A INVX1_LOC_34/A 0.05fF
C49854 INVX1_LOC_57/Y INVX1_LOC_140/A 0.10fF
C49855 INVX1_LOC_174/A INVX1_LOC_193/Y 0.01fF
C49856 NOR2X1_LOC_309/Y INVX1_LOC_22/A 0.03fF
C49857 INVX1_LOC_104/A INVX1_LOC_53/Y 0.06fF
C49858 INVX1_LOC_18/A NAND2X1_LOC_807/Y 0.07fF
C49859 INVX1_LOC_181/Y INPUT_1 0.00fF
C49860 INVX1_LOC_31/A NOR2X1_LOC_185/a_36_216# 0.01fF
C49861 INVX1_LOC_17/A INVX1_LOC_315/Y 0.05fF
C49862 INVX1_LOC_258/A NOR2X1_LOC_45/B 0.02fF
C49863 NOR2X1_LOC_500/Y INVX1_LOC_177/A 1.39fF
C49864 INVX1_LOC_279/A NOR2X1_LOC_142/Y 0.10fF
C49865 NOR2X1_LOC_468/Y INVX1_LOC_95/A 0.00fF
C49866 INVX1_LOC_72/A NAND2X1_LOC_863/A 0.55fF
C49867 NOR2X1_LOC_612/Y INVX1_LOC_57/A 0.01fF
C49868 INVX1_LOC_35/A NOR2X1_LOC_707/A 0.07fF
C49869 INVX1_LOC_78/A NOR2X1_LOC_127/Y 0.08fF
C49870 INVX1_LOC_172/A NAND2X1_LOC_866/B 1.25fF
C49871 INVX1_LOC_132/A INVX1_LOC_65/Y 0.01fF
C49872 NAND2X1_LOC_471/Y NAND2X1_LOC_477/Y 0.00fF
C49873 INVX1_LOC_120/A INVX1_LOC_33/A 0.00fF
C49874 NOR2X1_LOC_208/Y NOR2X1_LOC_735/Y -0.01fF
C49875 INVX1_LOC_36/A INVX1_LOC_100/A 0.23fF
C49876 INVX1_LOC_58/A NAND2X1_LOC_93/B 0.07fF
C49877 NAND2X1_LOC_455/B NAND2X1_LOC_445/a_36_24# 0.01fF
C49878 INVX1_LOC_32/A NAND2X1_LOC_80/a_36_24# 0.06fF
C49879 NAND2X1_LOC_555/Y INVX1_LOC_315/Y 0.22fF
C49880 NAND2X1_LOC_767/a_36_24# NOR2X1_LOC_78/A 0.00fF
C49881 INVX1_LOC_136/A NOR2X1_LOC_188/A 0.13fF
C49882 INVX1_LOC_35/A NOR2X1_LOC_209/B 0.03fF
C49883 INVX1_LOC_225/A NOR2X1_LOC_245/a_36_216# 0.00fF
C49884 INVX1_LOC_172/A NAND2X1_LOC_807/Y 0.03fF
C49885 NAND2X1_LOC_579/A NOR2X1_LOC_305/Y 0.02fF
C49886 NOR2X1_LOC_267/A INVX1_LOC_100/A 0.10fF
C49887 NAND2X1_LOC_391/Y NOR2X1_LOC_813/Y 0.01fF
C49888 INVX1_LOC_177/A INVX1_LOC_10/A 0.03fF
C49889 NOR2X1_LOC_92/Y INVX1_LOC_37/A 0.07fF
C49890 NOR2X1_LOC_479/B NOR2X1_LOC_375/Y 0.20fF
C49891 NOR2X1_LOC_282/Y NOR2X1_LOC_653/Y 0.05fF
C49892 INVX1_LOC_34/A INVX1_LOC_55/Y 0.03fF
C49893 INVX1_LOC_18/A INVX1_LOC_6/A 0.73fF
C49894 NOR2X1_LOC_655/B INVX1_LOC_279/A 0.01fF
C49895 NAND2X1_LOC_656/Y NAND2X1_LOC_660/A 0.03fF
C49896 INVX1_LOC_24/Y INVX1_LOC_37/A 0.66fF
C49897 NOR2X1_LOC_13/Y INVX1_LOC_144/A 0.10fF
C49898 NOR2X1_LOC_703/B NOR2X1_LOC_794/A 0.01fF
C49899 NOR2X1_LOC_389/A INVX1_LOC_95/A 0.04fF
C49900 INVX1_LOC_26/A NOR2X1_LOC_721/B 0.44fF
C49901 INVX1_LOC_53/A NOR2X1_LOC_197/B 0.10fF
C49902 NOR2X1_LOC_15/Y NAND2X1_LOC_804/Y 0.02fF
C49903 INVX1_LOC_280/Y INVX1_LOC_10/A 0.03fF
C49904 INVX1_LOC_49/Y NAND2X1_LOC_175/Y 0.03fF
C49905 NAND2X1_LOC_563/Y INPUT_1 0.05fF
C49906 NAND2X1_LOC_391/Y INVX1_LOC_280/A 0.01fF
C49907 NOR2X1_LOC_155/A NOR2X1_LOC_717/A 0.00fF
C49908 NAND2X1_LOC_354/B INVX1_LOC_28/A 0.02fF
C49909 INVX1_LOC_17/A NAND2X1_LOC_211/Y 0.00fF
C49910 INVX1_LOC_83/A INVX1_LOC_143/A 0.07fF
C49911 INVX1_LOC_228/Y VDD 0.26fF
C49912 INVX1_LOC_223/A NOR2X1_LOC_78/A 0.07fF
C49913 NAND2X1_LOC_483/Y NAND2X1_LOC_560/A 0.03fF
C49914 NOR2X1_LOC_846/A INVX1_LOC_9/A 0.01fF
C49915 INVX1_LOC_303/A NOR2X1_LOC_74/A 0.08fF
C49916 INVX1_LOC_200/A VDD 0.42fF
C49917 NOR2X1_LOC_246/A NAND2X1_LOC_231/Y 0.10fF
C49918 NAND2X1_LOC_476/Y INVX1_LOC_270/A 0.08fF
C49919 NOR2X1_LOC_282/Y INVX1_LOC_19/A 0.01fF
C49920 NOR2X1_LOC_78/B NOR2X1_LOC_130/A 0.07fF
C49921 INVX1_LOC_182/Y NOR2X1_LOC_142/Y 0.03fF
C49922 INVX1_LOC_314/Y INVX1_LOC_92/Y 0.04fF
C49923 NOR2X1_LOC_328/Y NOR2X1_LOC_561/Y 0.13fF
C49924 INVX1_LOC_121/Y NOR2X1_LOC_302/Y 0.01fF
C49925 NOR2X1_LOC_590/A NOR2X1_LOC_35/Y 0.06fF
C49926 NOR2X1_LOC_99/Y INVX1_LOC_306/Y 0.27fF
C49927 INVX1_LOC_136/A NOR2X1_LOC_43/Y 0.07fF
C49928 INVX1_LOC_5/A INVX1_LOC_179/A 0.13fF
C49929 INVX1_LOC_236/Y INVX1_LOC_20/A 0.00fF
C49930 INVX1_LOC_227/A INVX1_LOC_16/A 0.08fF
C49931 NOR2X1_LOC_703/B NOR2X1_LOC_552/A 0.01fF
C49932 INVX1_LOC_303/A NOR2X1_LOC_9/Y 0.03fF
C49933 INVX1_LOC_284/Y INVX1_LOC_20/A 0.03fF
C49934 INVX1_LOC_172/A INVX1_LOC_6/A 0.07fF
C49935 INVX1_LOC_194/A NAND2X1_LOC_462/a_36_24# 0.00fF
C49936 NOR2X1_LOC_718/Y INVX1_LOC_311/A 0.05fF
C49937 NAND2X1_LOC_733/Y VDD 5.14fF
C49938 NAND2X1_LOC_223/B GATE_222 0.05fF
C49939 INVX1_LOC_77/A NOR2X1_LOC_685/A 0.01fF
C49940 NOR2X1_LOC_468/Y INVX1_LOC_54/A 0.02fF
C49941 INVX1_LOC_77/A INVX1_LOC_186/A 0.10fF
C49942 NAND2X1_LOC_9/Y NAND2X1_LOC_773/B 0.23fF
C49943 NOR2X1_LOC_334/A NOR2X1_LOC_285/B 0.03fF
C49944 NOR2X1_LOC_655/B INVX1_LOC_182/Y 0.02fF
C49945 NOR2X1_LOC_92/Y NOR2X1_LOC_743/Y 0.03fF
C49946 NOR2X1_LOC_727/B NOR2X1_LOC_833/B 0.81fF
C49947 INVX1_LOC_103/A NOR2X1_LOC_351/Y 0.02fF
C49948 NOR2X1_LOC_130/A NAND2X1_LOC_392/Y 0.06fF
C49949 NOR2X1_LOC_488/Y INVX1_LOC_28/A 0.03fF
C49950 NOR2X1_LOC_295/Y INVX1_LOC_286/A 0.02fF
C49951 NOR2X1_LOC_383/B INVX1_LOC_42/A 0.03fF
C49952 INVX1_LOC_24/A NOR2X1_LOC_164/Y 0.06fF
C49953 NAND2X1_LOC_783/A INVX1_LOC_83/A 0.23fF
C49954 NOR2X1_LOC_120/a_36_216# NOR2X1_LOC_121/A 0.00fF
C49955 NOR2X1_LOC_470/B INVX1_LOC_92/A 0.16fF
C49956 NAND2X1_LOC_355/Y INVX1_LOC_146/Y 0.06fF
C49957 INVX1_LOC_217/A VDD 1.58fF
C49958 NOR2X1_LOC_860/B NOR2X1_LOC_332/B 0.00fF
C49959 INVX1_LOC_83/A NOR2X1_LOC_130/A 0.05fF
C49960 NAND2X1_LOC_355/Y VDD 0.03fF
C49961 NAND2X1_LOC_170/A INVX1_LOC_140/A 0.03fF
C49962 NOR2X1_LOC_203/Y NOR2X1_LOC_74/A 0.01fF
C49963 INVX1_LOC_77/A NAND2X1_LOC_447/Y 0.01fF
C49964 INVX1_LOC_89/A INVX1_LOC_306/A 0.01fF
C49965 NOR2X1_LOC_757/A NOR2X1_LOC_122/Y 0.18fF
C49966 INVX1_LOC_6/A NOR2X1_LOC_709/a_36_216# 0.00fF
C49967 INVX1_LOC_24/A INVX1_LOC_46/A 2.47fF
C49968 INVX1_LOC_33/A NOR2X1_LOC_542/B 0.02fF
C49969 NOR2X1_LOC_389/A INVX1_LOC_54/A 0.01fF
C49970 INVX1_LOC_75/A INVX1_LOC_1/Y 1.27fF
C49971 NOR2X1_LOC_742/A NOR2X1_LOC_302/B 0.03fF
C49972 INVX1_LOC_227/A INVX1_LOC_28/A 0.07fF
C49973 NOR2X1_LOC_592/A NOR2X1_LOC_592/B 0.01fF
C49974 INVX1_LOC_49/A INVX1_LOC_115/A 0.00fF
C49975 INVX1_LOC_41/A NOR2X1_LOC_631/B 0.04fF
C49976 INVX1_LOC_279/A INVX1_LOC_182/A 1.26fF
C49977 NOR2X1_LOC_316/Y NOR2X1_LOC_78/A 0.01fF
C49978 NAND2X1_LOC_725/B INVX1_LOC_5/Y 0.01fF
C49979 NAND2X1_LOC_199/B INVX1_LOC_54/A 0.04fF
C49980 INVX1_LOC_33/A INVX1_LOC_143/Y 0.13fF
C49981 NOR2X1_LOC_220/A INVX1_LOC_286/A 0.00fF
C49982 NOR2X1_LOC_38/B NAND2X1_LOC_215/A 0.08fF
C49983 INVX1_LOC_13/A INPUT_0 0.14fF
C49984 NOR2X1_LOC_256/Y INVX1_LOC_234/A 0.01fF
C49985 VDD NAND2X1_LOC_787/B 1.30fF
C49986 NAND2X1_LOC_708/a_36_24# INVX1_LOC_54/A 0.01fF
C49987 NAND2X1_LOC_2/a_36_24# GATE_662 0.00fF
C49988 INVX1_LOC_78/A NOR2X1_LOC_383/B 0.06fF
C49989 INVX1_LOC_230/Y NOR2X1_LOC_216/B 0.07fF
C49990 NAND2X1_LOC_474/Y NAND2X1_LOC_81/B 0.07fF
C49991 NOR2X1_LOC_510/Y INVX1_LOC_12/A 0.02fF
C49992 NOR2X1_LOC_180/Y INVX1_LOC_247/A 0.53fF
C49993 INVX1_LOC_30/A INVX1_LOC_185/A 0.01fF
C49994 NAND2X1_LOC_9/Y NOR2X1_LOC_393/Y 0.01fF
C49995 INVX1_LOC_286/Y INVX1_LOC_92/A 0.07fF
C49996 NOR2X1_LOC_557/Y INVX1_LOC_46/A 0.03fF
C49997 INVX1_LOC_34/A NOR2X1_LOC_357/Y 0.10fF
C49998 INVX1_LOC_58/A NAND2X1_LOC_470/B 0.03fF
C49999 INVX1_LOC_41/A INVX1_LOC_37/A 3.29fF
C50000 NOR2X1_LOC_52/B NAND2X1_LOC_241/Y 0.01fF
C50001 INVX1_LOC_107/A INVX1_LOC_54/A 0.01fF
C50002 NOR2X1_LOC_658/Y NOR2X1_LOC_155/A 0.07fF
C50003 NOR2X1_LOC_443/Y INVX1_LOC_26/Y 0.55fF
C50004 NOR2X1_LOC_685/A NOR2X1_LOC_687/Y 0.06fF
C50005 NOR2X1_LOC_194/Y NAND2X1_LOC_39/Y 0.00fF
C50006 INVX1_LOC_285/Y INVX1_LOC_10/A 0.10fF
C50007 NOR2X1_LOC_65/B NOR2X1_LOC_383/B 0.03fF
C50008 NOR2X1_LOC_246/A INPUT_0 0.07fF
C50009 NOR2X1_LOC_596/A INVX1_LOC_54/A 0.07fF
C50010 NAND2X1_LOC_349/B NOR2X1_LOC_318/B 0.06fF
C50011 INVX1_LOC_304/Y VDD 1.38fF
C50012 INVX1_LOC_95/Y INVX1_LOC_43/A 0.03fF
C50013 NOR2X1_LOC_458/B INVX1_LOC_247/A 0.02fF
C50014 NAND2X1_LOC_860/A NOR2X1_LOC_316/a_36_216# 0.01fF
C50015 INPUT_0 NOR2X1_LOC_174/B 0.06fF
C50016 NOR2X1_LOC_68/A NOR2X1_LOC_156/Y 0.08fF
C50017 INVX1_LOC_93/Y INVX1_LOC_25/Y 0.01fF
C50018 NAND2X1_LOC_734/B NAND2X1_LOC_721/A 0.10fF
C50019 NOR2X1_LOC_361/B INVX1_LOC_12/A 0.91fF
C50020 NAND2X1_LOC_860/A INVX1_LOC_26/A 0.07fF
C50021 NOR2X1_LOC_500/B NOR2X1_LOC_243/B 0.02fF
C50022 INVX1_LOC_182/A INVX1_LOC_182/Y 0.03fF
C50023 NOR2X1_LOC_315/Y INVX1_LOC_12/Y 0.33fF
C50024 INVX1_LOC_17/A NAND2X1_LOC_207/B 0.04fF
C50025 NAND2X1_LOC_715/B INVX1_LOC_128/Y 0.12fF
C50026 INVX1_LOC_34/A NOR2X1_LOC_692/Y 0.25fF
C50027 NAND2X1_LOC_728/Y NAND2X1_LOC_810/B 0.00fF
C50028 INVX1_LOC_143/A INVX1_LOC_46/A 0.01fF
C50029 NOR2X1_LOC_334/Y NOR2X1_LOC_674/Y 0.01fF
C50030 NAND2X1_LOC_575/a_36_24# NOR2X1_LOC_48/B 0.00fF
C50031 INVX1_LOC_214/Y VDD 0.17fF
C50032 NOR2X1_LOC_598/B NOR2X1_LOC_727/B 0.03fF
C50033 NOR2X1_LOC_742/A INVX1_LOC_75/A 0.07fF
C50034 NAND2X1_LOC_114/B INVX1_LOC_29/A 0.09fF
C50035 INVX1_LOC_135/A INVX1_LOC_91/A 0.10fF
C50036 INVX1_LOC_36/A NAND2X1_LOC_476/Y 0.01fF
C50037 NOR2X1_LOC_566/Y VDD 0.03fF
C50038 NAND2X1_LOC_392/A INVX1_LOC_20/A 0.00fF
C50039 NOR2X1_LOC_92/a_36_216# INVX1_LOC_56/Y 0.00fF
C50040 INVX1_LOC_72/A INVX1_LOC_294/A 0.02fF
C50041 NAND2X1_LOC_660/Y NAND2X1_LOC_468/B 0.03fF
C50042 NOR2X1_LOC_328/Y INVX1_LOC_76/A 0.02fF
C50043 NOR2X1_LOC_791/B INVX1_LOC_84/A 0.01fF
C50044 D_INPUT_0 NAND2X1_LOC_655/A 0.01fF
C50045 NAND2X1_LOC_116/A INVX1_LOC_9/A 0.00fF
C50046 INVX1_LOC_283/Y INVX1_LOC_92/A 0.06fF
C50047 NOR2X1_LOC_295/Y INVX1_LOC_54/A 0.02fF
C50048 INVX1_LOC_295/A INVX1_LOC_91/A 0.01fF
C50049 NOR2X1_LOC_602/A INVX1_LOC_19/A 0.06fF
C50050 NOR2X1_LOC_490/Y INVX1_LOC_309/A 0.01fF
C50051 NOR2X1_LOC_355/A NOR2X1_LOC_405/A 0.02fF
C50052 NOR2X1_LOC_299/Y NOR2X1_LOC_396/Y 0.03fF
C50053 D_GATE_222 VDD 0.16fF
C50054 NOR2X1_LOC_97/B NOR2X1_LOC_332/B 0.36fF
C50055 NOR2X1_LOC_858/A NOR2X1_LOC_678/A 0.01fF
C50056 INVX1_LOC_279/A NAND2X1_LOC_274/a_36_24# 0.00fF
C50057 INVX1_LOC_10/A NOR2X1_LOC_137/B 0.03fF
C50058 NOR2X1_LOC_707/B INVX1_LOC_19/A 0.29fF
C50059 NAND2X1_LOC_128/a_36_24# NOR2X1_LOC_269/Y 0.00fF
C50060 NOR2X1_LOC_389/A NAND2X1_LOC_807/B 0.57fF
C50061 INVX1_LOC_83/A NOR2X1_LOC_209/A 0.23fF
C50062 NOR2X1_LOC_763/A INVX1_LOC_78/A 0.01fF
C50063 NOR2X1_LOC_719/a_36_216# INVX1_LOC_59/Y 0.01fF
C50064 INVX1_LOC_153/Y INVX1_LOC_307/A 0.27fF
C50065 INVX1_LOC_235/Y NOR2X1_LOC_415/Y 0.02fF
C50066 NAND2X1_LOC_787/A NOR2X1_LOC_754/Y 0.02fF
C50067 NOR2X1_LOC_130/A NOR2X1_LOC_368/Y 0.01fF
C50068 NOR2X1_LOC_352/Y NOR2X1_LOC_331/B 0.01fF
C50069 NOR2X1_LOC_730/A VDD 0.24fF
C50070 NAND2X1_LOC_291/a_36_24# NOR2X1_LOC_334/A 0.01fF
C50071 NAND2X1_LOC_504/a_36_24# NOR2X1_LOC_349/A 0.01fF
C50072 NOR2X1_LOC_490/Y INVX1_LOC_91/A 0.04fF
C50073 INVX1_LOC_178/A NOR2X1_LOC_693/Y 0.10fF
C50074 NOR2X1_LOC_208/Y NAND2X1_LOC_476/Y 0.09fF
C50075 INVX1_LOC_24/Y NAND2X1_LOC_72/B 0.15fF
C50076 NAND2X1_LOC_477/A NOR2X1_LOC_743/Y 0.01fF
C50077 NOR2X1_LOC_525/Y INVX1_LOC_20/A 0.06fF
C50078 NAND2X1_LOC_722/A INVX1_LOC_185/A 0.02fF
C50079 INVX1_LOC_89/A INVX1_LOC_59/Y 0.06fF
C50080 INVX1_LOC_240/A INVX1_LOC_241/Y 0.08fF
C50081 INVX1_LOC_177/A NOR2X1_LOC_801/a_36_216# 0.00fF
C50082 NOR2X1_LOC_392/B NOR2X1_LOC_831/B 0.42fF
C50083 INVX1_LOC_121/A INVX1_LOC_37/A 0.01fF
C50084 NOR2X1_LOC_312/Y INVX1_LOC_20/A 0.13fF
C50085 VDD NAND2X1_LOC_808/A -0.00fF
C50086 INVX1_LOC_57/Y INVX1_LOC_42/A 0.03fF
C50087 INVX1_LOC_181/Y NAND2X1_LOC_63/Y 0.00fF
C50088 NOR2X1_LOC_577/Y INVX1_LOC_63/A 0.07fF
C50089 NOR2X1_LOC_130/A INVX1_LOC_46/A 0.03fF
C50090 INVX1_LOC_177/A INVX1_LOC_307/A 0.00fF
C50091 NOR2X1_LOC_318/B INVX1_LOC_75/A 0.25fF
C50092 INVX1_LOC_89/A INVX1_LOC_176/A 0.02fF
C50093 INVX1_LOC_130/A INVX1_LOC_15/A 0.05fF
C50094 NOR2X1_LOC_756/Y INVX1_LOC_95/Y 0.02fF
C50095 NOR2X1_LOC_168/B NOR2X1_LOC_634/A 0.73fF
C50096 INVX1_LOC_232/A INVX1_LOC_9/A 0.02fF
C50097 NOR2X1_LOC_598/B NOR2X1_LOC_649/Y 0.22fF
C50098 NOR2X1_LOC_811/A NOR2X1_LOC_808/B 0.05fF
C50099 INVX1_LOC_177/A NOR2X1_LOC_445/B 0.00fF
C50100 INVX1_LOC_269/A NAND2X1_LOC_99/A 0.10fF
C50101 INVX1_LOC_75/A INVX1_LOC_93/Y 0.08fF
C50102 NOR2X1_LOC_160/B INVX1_LOC_94/Y 0.05fF
C50103 NOR2X1_LOC_124/B INVX1_LOC_84/A 0.02fF
C50104 NOR2X1_LOC_173/Y INVX1_LOC_23/A 0.66fF
C50105 INVX1_LOC_34/A NAND2X1_LOC_489/Y 0.03fF
C50106 INVX1_LOC_314/Y INVX1_LOC_106/A -0.01fF
C50107 INVX1_LOC_92/Y NOR2X1_LOC_557/A 0.02fF
C50108 NOR2X1_LOC_78/B NOR2X1_LOC_197/B 0.03fF
C50109 D_INPUT_7 INVX1_LOC_15/A 0.01fF
C50110 NAND2X1_LOC_323/B NAND2X1_LOC_413/a_36_24# 0.01fF
C50111 NOR2X1_LOC_515/a_36_216# NOR2X1_LOC_649/B 0.01fF
C50112 NOR2X1_LOC_91/A NAND2X1_LOC_793/Y 0.03fF
C50113 NOR2X1_LOC_516/a_36_216# NAND2X1_LOC_82/Y 0.00fF
C50114 NOR2X1_LOC_68/A D_INPUT_5 0.03fF
C50115 NOR2X1_LOC_794/A INVX1_LOC_91/A 0.02fF
C50116 INVX1_LOC_22/A NOR2X1_LOC_435/A 0.03fF
C50117 NAND2X1_LOC_337/B NAND2X1_LOC_288/B 0.01fF
C50118 NOR2X1_LOC_248/Y NOR2X1_LOC_248/A 0.00fF
C50119 INVX1_LOC_75/A INVX1_LOC_139/A 0.01fF
C50120 INVX1_LOC_179/Y INVX1_LOC_220/A 0.36fF
C50121 NAND2X1_LOC_795/Y INVX1_LOC_54/A 0.01fF
C50122 INVX1_LOC_72/A NOR2X1_LOC_334/Y 0.07fF
C50123 INVX1_LOC_153/Y INVX1_LOC_12/A 0.12fF
C50124 INVX1_LOC_57/Y INVX1_LOC_78/A 0.96fF
C50125 NOR2X1_LOC_647/A INVX1_LOC_31/A 0.05fF
C50126 NOR2X1_LOC_332/A NOR2X1_LOC_332/Y 0.15fF
C50127 NAND2X1_LOC_640/Y INVX1_LOC_102/A -0.01fF
C50128 NOR2X1_LOC_599/a_36_216# NOR2X1_LOC_409/B 0.00fF
C50129 INVX1_LOC_58/A INVX1_LOC_256/A 0.39fF
C50130 INVX1_LOC_95/A INVX1_LOC_100/Y 0.01fF
C50131 INVX1_LOC_81/A INVX1_LOC_15/A 0.03fF
C50132 NOR2X1_LOC_552/A INVX1_LOC_91/A 2.95fF
C50133 NOR2X1_LOC_274/Y INVX1_LOC_47/Y 0.02fF
C50134 INVX1_LOC_292/A NOR2X1_LOC_748/A 0.10fF
C50135 NOR2X1_LOC_87/B NAND2X1_LOC_207/Y 0.03fF
C50136 NOR2X1_LOC_646/A INVX1_LOC_84/A 0.65fF
C50137 NOR2X1_LOC_82/A NOR2X1_LOC_392/Y 0.16fF
C50138 NOR2X1_LOC_168/B INVX1_LOC_29/A 0.03fF
C50139 NOR2X1_LOC_512/Y INVX1_LOC_78/A 0.00fF
C50140 INVX1_LOC_36/A NOR2X1_LOC_843/B 0.05fF
C50141 INVX1_LOC_177/A INVX1_LOC_12/A 0.10fF
C50142 NOR2X1_LOC_591/a_36_216# INVX1_LOC_42/A 0.00fF
C50143 INVX1_LOC_306/Y NOR2X1_LOC_271/B 0.39fF
C50144 NAND2X1_LOC_360/B NAND2X1_LOC_74/B 0.01fF
C50145 D_INPUT_1 INVX1_LOC_61/Y 0.08fF
C50146 INVX1_LOC_22/A INVX1_LOC_63/A 0.24fF
C50147 NAND2X1_LOC_116/A NOR2X1_LOC_861/Y 0.07fF
C50148 INVX1_LOC_34/A INVX1_LOC_32/A 1.15fF
C50149 NOR2X1_LOC_710/a_36_216# INVX1_LOC_117/A 0.00fF
C50150 INVX1_LOC_132/Y NOR2X1_LOC_634/A 0.02fF
C50151 INVX1_LOC_304/A NOR2X1_LOC_124/A 0.06fF
C50152 INVX1_LOC_21/A NOR2X1_LOC_15/Y 0.25fF
C50153 INVX1_LOC_280/Y INVX1_LOC_12/A 0.03fF
C50154 D_INPUT_0 NAND2X1_LOC_141/Y 0.11fF
C50155 NOR2X1_LOC_644/Y INVX1_LOC_290/Y 0.03fF
C50156 NOR2X1_LOC_56/a_36_216# NOR2X1_LOC_56/Y 0.00fF
C50157 INVX1_LOC_286/Y INVX1_LOC_53/A 0.07fF
C50158 INVX1_LOC_18/A INVX1_LOC_270/A 0.15fF
C50159 NAND2X1_LOC_181/Y NOR2X1_LOC_89/A 0.03fF
C50160 INVX1_LOC_226/Y NAND2X1_LOC_81/B 0.01fF
C50161 NAND2X1_LOC_20/B NOR2X1_LOC_249/Y 0.03fF
C50162 NOR2X1_LOC_717/a_36_216# NAND2X1_LOC_454/Y 0.01fF
C50163 NOR2X1_LOC_802/A INVX1_LOC_15/A 0.04fF
C50164 NAND2X1_LOC_823/a_36_24# INVX1_LOC_37/A 0.00fF
C50165 NAND2X1_LOC_194/a_36_24# NOR2X1_LOC_89/A 0.00fF
C50166 NOR2X1_LOC_682/Y NAND2X1_LOC_655/A 0.03fF
C50167 NAND2X1_LOC_563/Y NAND2X1_LOC_618/Y 0.43fF
C50168 INVX1_LOC_135/A INVX1_LOC_203/A 0.02fF
C50169 NOR2X1_LOC_405/A NOR2X1_LOC_111/A 0.28fF
C50170 NAND2X1_LOC_231/Y INVX1_LOC_32/A 0.03fF
C50171 INVX1_LOC_34/A NAND2X1_LOC_175/Y 0.07fF
C50172 NOR2X1_LOC_637/A INVX1_LOC_23/A 0.01fF
C50173 NOR2X1_LOC_152/A INVX1_LOC_91/A 0.06fF
C50174 INVX1_LOC_213/Y INVX1_LOC_271/Y 0.01fF
C50175 NOR2X1_LOC_222/a_36_216# INVX1_LOC_109/Y 0.01fF
C50176 NOR2X1_LOC_607/A INVX1_LOC_23/A 0.01fF
C50177 NOR2X1_LOC_171/a_36_216# INVX1_LOC_272/A 0.01fF
C50178 NOR2X1_LOC_15/Y NOR2X1_LOC_469/a_36_216# 0.00fF
C50179 NOR2X1_LOC_641/B INVX1_LOC_5/A 0.02fF
C50180 INVX1_LOC_159/A INVX1_LOC_53/A 0.07fF
C50181 INVX1_LOC_113/Y NOR2X1_LOC_383/B 0.68fF
C50182 NOR2X1_LOC_721/Y INVX1_LOC_92/A 0.09fF
C50183 INVX1_LOC_298/Y INVX1_LOC_88/Y 0.03fF
C50184 NOR2X1_LOC_655/B NOR2X1_LOC_38/B 0.01fF
C50185 INVX1_LOC_91/A INVX1_LOC_280/A -0.01fF
C50186 NAND2X1_LOC_287/B INVX1_LOC_20/A 0.11fF
C50187 NAND2X1_LOC_656/Y INVX1_LOC_29/A 0.10fF
C50188 NAND2X1_LOC_848/A NAND2X1_LOC_655/A 0.02fF
C50189 INVX1_LOC_205/Y NOR2X1_LOC_160/B 0.02fF
C50190 NOR2X1_LOC_191/B INVX1_LOC_53/A 0.01fF
C50191 NAND2X1_LOC_9/Y INVX1_LOC_24/A 0.22fF
C50192 INVX1_LOC_18/A NOR2X1_LOC_109/Y 0.07fF
C50193 INVX1_LOC_266/Y NOR2X1_LOC_158/Y 0.01fF
C50194 NOR2X1_LOC_315/Y NOR2X1_LOC_89/Y 0.01fF
C50195 NOR2X1_LOC_751/Y INVX1_LOC_5/A 0.06fF
C50196 INVX1_LOC_233/A INVX1_LOC_24/A 0.07fF
C50197 INVX1_LOC_285/Y INVX1_LOC_307/A 0.12fF
C50198 NOR2X1_LOC_749/Y INVX1_LOC_125/A 0.01fF
C50199 NOR2X1_LOC_130/A NOR2X1_LOC_671/Y 0.02fF
C50200 INVX1_LOC_299/A NOR2X1_LOC_160/B 0.03fF
C50201 INVX1_LOC_13/Y NOR2X1_LOC_791/A 0.03fF
C50202 INVX1_LOC_279/A NOR2X1_LOC_850/B 0.01fF
C50203 INVX1_LOC_214/A INVX1_LOC_273/A 0.05fF
C50204 NOR2X1_LOC_285/A NOR2X1_LOC_285/B 0.07fF
C50205 NOR2X1_LOC_667/A INVX1_LOC_273/A 0.02fF
C50206 NAND2X1_LOC_231/Y NAND2X1_LOC_175/Y 0.28fF
C50207 INVX1_LOC_144/A NOR2X1_LOC_697/Y 0.09fF
C50208 INVX1_LOC_33/Y INVX1_LOC_76/A 0.03fF
C50209 NOR2X1_LOC_598/B NAND2X1_LOC_364/Y 0.01fF
C50210 INVX1_LOC_225/A NOR2X1_LOC_280/a_36_216# 0.00fF
C50211 NAND2X1_LOC_537/Y INVX1_LOC_141/A 0.02fF
C50212 NOR2X1_LOC_500/Y INVX1_LOC_4/Y 0.01fF
C50213 NAND2X1_LOC_795/Y NOR2X1_LOC_48/B 0.06fF
C50214 INVX1_LOC_226/Y INVX1_LOC_4/Y 0.10fF
C50215 NOR2X1_LOC_538/B NOR2X1_LOC_160/B 0.02fF
C50216 NOR2X1_LOC_564/Y INVX1_LOC_19/A 0.03fF
C50217 NAND2X1_LOC_638/Y INVX1_LOC_29/A 0.01fF
C50218 NOR2X1_LOC_272/Y NAND2X1_LOC_364/A 0.03fF
C50219 NAND2X1_LOC_553/A INVX1_LOC_24/A 0.02fF
C50220 NAND2X1_LOC_584/a_36_24# NOR2X1_LOC_635/B 0.00fF
C50221 INVX1_LOC_208/A INVX1_LOC_94/Y 0.00fF
C50222 NAND2X1_LOC_850/Y NOR2X1_LOC_278/Y 0.07fF
C50223 INVX1_LOC_33/Y NAND2X1_LOC_405/a_36_24# 0.00fF
C50224 NAND2X1_LOC_447/Y INVX1_LOC_9/A 0.10fF
C50225 INVX1_LOC_269/A NAND2X1_LOC_577/A 0.22fF
C50226 NAND2X1_LOC_508/A NOR2X1_LOC_340/A 4.15fF
C50227 NOR2X1_LOC_211/A NAND2X1_LOC_72/B 0.03fF
C50228 NOR2X1_LOC_798/A INVX1_LOC_24/A 0.03fF
C50229 INVX1_LOC_71/A NOR2X1_LOC_81/Y 0.06fF
C50230 INVX1_LOC_224/Y NOR2X1_LOC_709/A 0.17fF
C50231 INVX1_LOC_136/A NAND2X1_LOC_326/A 0.03fF
C50232 INVX1_LOC_36/A NAND2X1_LOC_216/a_36_24# 0.00fF
C50233 INVX1_LOC_36/A NOR2X1_LOC_536/Y 0.01fF
C50234 INVX1_LOC_45/A NAND2X1_LOC_538/Y 0.13fF
C50235 INVX1_LOC_65/A INVX1_LOC_307/A 0.02fF
C50236 NOR2X1_LOC_845/A NAND2X1_LOC_85/Y 0.05fF
C50237 NOR2X1_LOC_590/A INVX1_LOC_246/A 0.07fF
C50238 INVX1_LOC_21/A NOR2X1_LOC_860/B 0.14fF
C50239 NAND2X1_LOC_338/B NAND2X1_LOC_464/B 0.16fF
C50240 INVX1_LOC_10/A INVX1_LOC_4/Y 0.07fF
C50241 NOR2X1_LOC_92/Y NAND2X1_LOC_198/B 0.17fF
C50242 NAND2X1_LOC_703/Y INVX1_LOC_24/A 0.07fF
C50243 NAND2X1_LOC_588/B INVX1_LOC_1/A 0.06fF
C50244 NOR2X1_LOC_56/Y INVX1_LOC_92/A 0.03fF
C50245 INVX1_LOC_65/A NOR2X1_LOC_445/B 0.10fF
C50246 NOR2X1_LOC_99/B NOR2X1_LOC_38/B 0.07fF
C50247 INVX1_LOC_277/A NOR2X1_LOC_307/A 0.02fF
C50248 INVX1_LOC_25/A NAND2X1_LOC_342/Y 0.04fF
C50249 NAND2X1_LOC_53/Y NOR2X1_LOC_723/Y 0.05fF
C50250 NAND2X1_LOC_852/Y INVX1_LOC_296/Y 0.41fF
C50251 NOR2X1_LOC_328/Y NOR2X1_LOC_447/A 0.01fF
C50252 NOR2X1_LOC_163/A D_INPUT_5 0.00fF
C50253 NOR2X1_LOC_441/Y NOR2X1_LOC_389/A 0.03fF
C50254 NOR2X1_LOC_91/A INVX1_LOC_300/A 0.04fF
C50255 NOR2X1_LOC_447/B INVX1_LOC_54/A 0.02fF
C50256 INVX1_LOC_136/A NAND2X1_LOC_807/A 0.03fF
C50257 INVX1_LOC_50/A NOR2X1_LOC_553/Y 0.03fF
C50258 NOR2X1_LOC_742/A INVX1_LOC_283/A 0.01fF
C50259 INVX1_LOC_146/Y INVX1_LOC_92/A 0.07fF
C50260 NOR2X1_LOC_589/Y NOR2X1_LOC_89/A 0.01fF
C50261 INVX1_LOC_7/A INVX1_LOC_23/Y 0.11fF
C50262 VDD INVX1_LOC_92/A 1.12fF
C50263 INVX1_LOC_285/Y INVX1_LOC_12/A 0.09fF
C50264 NOR2X1_LOC_15/Y NOR2X1_LOC_596/a_36_216# 0.00fF
C50265 INVX1_LOC_313/Y NOR2X1_LOC_334/Y 1.47fF
C50266 NOR2X1_LOC_780/B INVX1_LOC_33/A 0.02fF
C50267 NAND2X1_LOC_721/B INVX1_LOC_141/Y 0.03fF
C50268 NOR2X1_LOC_75/Y NOR2X1_LOC_273/Y 0.03fF
C50269 INVX1_LOC_21/A NOR2X1_LOC_635/A 0.30fF
C50270 INVX1_LOC_31/A INVX1_LOC_205/A 0.00fF
C50271 INVX1_LOC_25/A NOR2X1_LOC_646/a_36_216# 0.00fF
C50272 NAND2X1_LOC_656/Y NOR2X1_LOC_318/a_36_216# 0.01fF
C50273 NOR2X1_LOC_286/a_36_216# INVX1_LOC_196/A 0.01fF
C50274 INVX1_LOC_17/A INVX1_LOC_8/Y 0.01fF
C50275 INVX1_LOC_17/A NOR2X1_LOC_637/B 0.30fF
C50276 NOR2X1_LOC_602/a_36_216# INVX1_LOC_45/A 0.00fF
C50277 NOR2X1_LOC_620/Y INVX1_LOC_224/A 0.03fF
C50278 NOR2X1_LOC_2/Y D_INPUT_5 0.07fF
C50279 NOR2X1_LOC_533/A NOR2X1_LOC_304/Y 0.24fF
C50280 NOR2X1_LOC_88/Y INVX1_LOC_37/Y 0.08fF
C50281 INPUT_0 INVX1_LOC_32/A 0.16fF
C50282 INVX1_LOC_17/A INVX1_LOC_155/A 0.04fF
C50283 NOR2X1_LOC_798/A INVX1_LOC_143/A 0.00fF
C50284 INVX1_LOC_211/Y NAND2X1_LOC_802/A 0.08fF
C50285 INVX1_LOC_2/Y INVX1_LOC_84/A 0.04fF
C50286 INVX1_LOC_36/A INVX1_LOC_18/A 0.33fF
C50287 NOR2X1_LOC_510/Y INVX1_LOC_214/Y 0.47fF
C50288 NOR2X1_LOC_163/Y INVX1_LOC_78/A 0.03fF
C50289 INVX1_LOC_35/A NAND2X1_LOC_41/Y 0.00fF
C50290 NOR2X1_LOC_380/Y NOR2X1_LOC_409/B 0.06fF
C50291 NAND2X1_LOC_623/B NOR2X1_LOC_89/A 0.01fF
C50292 NAND2X1_LOC_860/A INVX1_LOC_164/A 0.01fF
C50293 NAND2X1_LOC_728/Y INVX1_LOC_36/A 0.07fF
C50294 INVX1_LOC_17/A NOR2X1_LOC_264/Y 0.07fF
C50295 NOR2X1_LOC_590/A NOR2X1_LOC_350/A 0.08fF
C50296 NAND2X1_LOC_129/a_36_24# INVX1_LOC_84/A 0.00fF
C50297 NOR2X1_LOC_456/Y NOR2X1_LOC_717/B 0.07fF
C50298 NOR2X1_LOC_615/a_36_216# NOR2X1_LOC_690/A 0.01fF
C50299 INVX1_LOC_316/A INVX1_LOC_12/A 0.01fF
C50300 NOR2X1_LOC_725/A NOR2X1_LOC_460/A -0.00fF
C50301 INVX1_LOC_255/Y INVX1_LOC_5/A 0.03fF
C50302 INVX1_LOC_102/A NAND2X1_LOC_642/Y 0.11fF
C50303 NOR2X1_LOC_74/Y INVX1_LOC_78/A 0.01fF
C50304 INVX1_LOC_22/Y NOR2X1_LOC_350/A 0.26fF
C50305 NAND2X1_LOC_711/B INVX1_LOC_36/A 0.07fF
C50306 INVX1_LOC_119/A INVX1_LOC_103/A 0.02fF
C50307 NOR2X1_LOC_473/B INVX1_LOC_271/A 0.00fF
C50308 INVX1_LOC_12/A NOR2X1_LOC_137/B 0.03fF
C50309 NOR2X1_LOC_68/A NOR2X1_LOC_360/Y 0.03fF
C50310 INVX1_LOC_36/A NOR2X1_LOC_637/Y 0.03fF
C50311 INVX1_LOC_25/A NOR2X1_LOC_246/Y 0.03fF
C50312 NAND2X1_LOC_114/B INVX1_LOC_8/A 0.07fF
C50313 INVX1_LOC_34/A INPUT_3 0.02fF
C50314 INPUT_0 NAND2X1_LOC_175/Y 0.07fF
C50315 INVX1_LOC_233/A NOR2X1_LOC_130/A 0.07fF
C50316 INVX1_LOC_159/A NAND2X1_LOC_156/a_36_24# 0.00fF
C50317 NOR2X1_LOC_667/A NOR2X1_LOC_15/Y 0.09fF
C50318 NOR2X1_LOC_813/Y INVX1_LOC_203/A 0.03fF
C50319 INVX1_LOC_230/Y NOR2X1_LOC_84/A 0.00fF
C50320 NOR2X1_LOC_103/Y NOR2X1_LOC_709/A 0.17fF
C50321 INVX1_LOC_190/Y INVX1_LOC_53/A 0.01fF
C50322 NOR2X1_LOC_655/B NAND2X1_LOC_190/Y 0.03fF
C50323 NOR2X1_LOC_479/B INVX1_LOC_163/A 0.09fF
C50324 INVX1_LOC_255/Y INVX1_LOC_178/A 0.04fF
C50325 INVX1_LOC_39/Y INVX1_LOC_8/A 0.33fF
C50326 NOR2X1_LOC_67/Y NOR2X1_LOC_35/Y 0.10fF
C50327 INVX1_LOC_136/A NOR2X1_LOC_625/Y 0.06fF
C50328 NOR2X1_LOC_772/B D_INPUT_0 0.00fF
C50329 NOR2X1_LOC_160/B NOR2X1_LOC_315/Y 0.51fF
C50330 NOR2X1_LOC_750/Y NOR2X1_LOC_750/A 0.01fF
C50331 NOR2X1_LOC_481/A INVX1_LOC_223/A 0.01fF
C50332 INVX1_LOC_209/Y INVX1_LOC_72/A 0.05fF
C50333 NOR2X1_LOC_237/Y INVX1_LOC_18/A 0.15fF
C50334 INVX1_LOC_203/A INVX1_LOC_280/A 0.10fF
C50335 INVX1_LOC_21/A NOR2X1_LOC_97/B 0.29fF
C50336 NOR2X1_LOC_111/A NOR2X1_LOC_841/a_36_216# 0.01fF
C50337 INVX1_LOC_83/A INVX1_LOC_38/Y 0.02fF
C50338 NOR2X1_LOC_828/Y NOR2X1_LOC_828/B 0.12fF
C50339 NAND2X1_LOC_21/Y D_INPUT_7 0.41fF
C50340 NAND2X1_LOC_796/B NAND2X1_LOC_796/Y 0.05fF
C50341 INVX1_LOC_33/A NAND2X1_LOC_351/A 0.06fF
C50342 INVX1_LOC_13/Y D_INPUT_0 0.03fF
C50343 INVX1_LOC_299/A NOR2X1_LOC_516/B 0.03fF
C50344 NAND2X1_LOC_11/a_36_24# INVX1_LOC_174/A 0.00fF
C50345 NOR2X1_LOC_512/Y NOR2X1_LOC_152/Y 0.01fF
C50346 INVX1_LOC_229/A INVX1_LOC_241/A 0.24fF
C50347 NOR2X1_LOC_804/B INVX1_LOC_18/A 0.07fF
C50348 NOR2X1_LOC_205/Y NOR2X1_LOC_500/Y 0.02fF
C50349 INVX1_LOC_292/A NOR2X1_LOC_493/B 0.01fF
C50350 INVX1_LOC_224/A NAND2X1_LOC_194/a_36_24# 0.00fF
C50351 NOR2X1_LOC_269/Y NAND2X1_LOC_454/Y 0.01fF
C50352 NOR2X1_LOC_89/A INVX1_LOC_117/A 0.10fF
C50353 INVX1_LOC_124/Y INVX1_LOC_168/A 0.09fF
C50354 NOR2X1_LOC_447/B NOR2X1_LOC_48/B 0.05fF
C50355 NOR2X1_LOC_310/Y INVX1_LOC_30/A 0.01fF
C50356 INVX1_LOC_5/A NOR2X1_LOC_644/A 0.03fF
C50357 NAND2X1_LOC_169/Y INVX1_LOC_90/A 0.06fF
C50358 NOR2X1_LOC_335/B INVX1_LOC_29/Y 0.07fF
C50359 NOR2X1_LOC_82/A INVX1_LOC_25/Y 0.13fF
C50360 INVX1_LOC_41/A NAND2X1_LOC_198/B 0.01fF
C50361 NAND2X1_LOC_745/a_36_24# NOR2X1_LOC_781/B 0.00fF
C50362 INVX1_LOC_88/A NAND2X1_LOC_660/Y 0.02fF
C50363 NOR2X1_LOC_187/Y INVX1_LOC_279/A 0.02fF
C50364 NAND2X1_LOC_9/Y NOR2X1_LOC_112/B 0.01fF
C50365 INVX1_LOC_2/Y INVX1_LOC_15/A 0.03fF
C50366 NOR2X1_LOC_309/Y INVX1_LOC_18/A 0.25fF
C50367 NAND2X1_LOC_500/B INVX1_LOC_118/A 0.01fF
C50368 INVX1_LOC_280/Y NAND2X1_LOC_733/Y 0.03fF
C50369 INVX1_LOC_58/A INVX1_LOC_69/Y 0.10fF
C50370 INVX1_LOC_27/A NOR2X1_LOC_473/B 0.07fF
C50371 INVX1_LOC_229/A NOR2X1_LOC_298/Y 0.05fF
C50372 NAND2X1_LOC_559/Y NOR2X1_LOC_299/Y 0.03fF
C50373 NOR2X1_LOC_454/Y NOR2X1_LOC_207/a_36_216# 0.00fF
C50374 NOR2X1_LOC_596/A NOR2X1_LOC_142/Y 0.07fF
C50375 NAND2X1_LOC_803/B INVX1_LOC_290/A 0.04fF
C50376 INVX1_LOC_254/A NOR2X1_LOC_520/B 0.00fF
C50377 NOR2X1_LOC_205/Y INVX1_LOC_10/A 0.03fF
C50378 INVX1_LOC_36/A NOR2X1_LOC_709/a_36_216# 0.00fF
C50379 NOR2X1_LOC_470/B INVX1_LOC_83/A 0.02fF
C50380 INVX1_LOC_266/A INVX1_LOC_171/A 0.03fF
C50381 NOR2X1_LOC_45/Y NAND2X1_LOC_662/Y 0.03fF
C50382 NAND2X1_LOC_306/a_36_24# NOR2X1_LOC_52/B 0.00fF
C50383 INVX1_LOC_94/Y NAND2X1_LOC_211/Y 0.27fF
C50384 INVX1_LOC_280/Y INVX1_LOC_217/A 0.07fF
C50385 INVX1_LOC_103/A INVX1_LOC_89/A 0.03fF
C50386 NOR2X1_LOC_456/a_36_216# INVX1_LOC_182/A 0.01fF
C50387 INVX1_LOC_71/A NOR2X1_LOC_709/A 0.07fF
C50388 NAND2X1_LOC_582/a_36_24# INVX1_LOC_77/A 0.01fF
C50389 NOR2X1_LOC_830/Y INVX1_LOC_307/A 0.04fF
C50390 INVX1_LOC_76/A INVX1_LOC_23/Y 0.10fF
C50391 NOR2X1_LOC_13/Y NAND2X1_LOC_660/A 0.48fF
C50392 INVX1_LOC_136/A NOR2X1_LOC_165/Y 0.04fF
C50393 INVX1_LOC_133/Y NOR2X1_LOC_106/Y 0.11fF
C50394 NOR2X1_LOC_632/Y NOR2X1_LOC_717/Y 0.03fF
C50395 NOR2X1_LOC_78/B NOR2X1_LOC_191/B 0.05fF
C50396 NOR2X1_LOC_531/a_36_216# NOR2X1_LOC_500/Y 0.00fF
C50397 INVX1_LOC_31/A NOR2X1_LOC_686/B 0.02fF
C50398 INVX1_LOC_90/A D_GATE_741 0.03fF
C50399 NOR2X1_LOC_340/Y NOR2X1_LOC_844/A 0.02fF
C50400 NOR2X1_LOC_187/Y INVX1_LOC_182/Y 0.01fF
C50401 NAND2X1_LOC_190/Y INVX1_LOC_182/A 0.22fF
C50402 INVX1_LOC_36/A NOR2X1_LOC_690/Y 0.11fF
C50403 INVX1_LOC_164/Y INVX1_LOC_314/Y 0.09fF
C50404 INVX1_LOC_201/A NOR2X1_LOC_649/Y 0.20fF
C50405 INVX1_LOC_292/A INVX1_LOC_89/A 0.07fF
C50406 NAND2X1_LOC_741/B NOR2X1_LOC_561/Y 0.03fF
C50407 NOR2X1_LOC_456/Y NOR2X1_LOC_181/A 0.04fF
C50408 INVX1_LOC_225/A INVX1_LOC_162/Y 0.01fF
C50409 NAND2X1_LOC_562/Y NAND2X1_LOC_563/Y 0.03fF
C50410 INVX1_LOC_34/A NAND2X1_LOC_147/a_36_24# 0.00fF
C50411 INVX1_LOC_202/A NOR2X1_LOC_757/Y 0.17fF
C50412 NAND2X1_LOC_349/B NAND2X1_LOC_514/Y 0.03fF
C50413 INVX1_LOC_53/A NOR2X1_LOC_56/Y 0.29fF
C50414 NAND2X1_LOC_807/Y NAND2X1_LOC_793/Y 0.10fF
C50415 INVX1_LOC_90/A NAND2X1_LOC_352/B 0.11fF
C50416 INVX1_LOC_12/Y NAND2X1_LOC_99/A 0.48fF
C50417 NOR2X1_LOC_74/A INVX1_LOC_198/A -0.01fF
C50418 NOR2X1_LOC_78/B INVX1_LOC_283/Y 0.01fF
C50419 INVX1_LOC_280/Y NAND2X1_LOC_787/B 0.14fF
C50420 NOR2X1_LOC_392/Y NOR2X1_LOC_124/a_36_216# 0.00fF
C50421 NOR2X1_LOC_544/A INVX1_LOC_49/A 0.44fF
C50422 NOR2X1_LOC_389/B NAND2X1_LOC_352/B 0.55fF
C50423 D_INPUT_0 NOR2X1_LOC_500/B 0.11fF
C50424 NOR2X1_LOC_392/Y INVX1_LOC_59/Y 0.61fF
C50425 NAND2X1_LOC_579/A NAND2X1_LOC_858/B 0.12fF
C50426 INVX1_LOC_112/A NOR2X1_LOC_392/Y 0.02fF
C50427 INVX1_LOC_45/A NOR2X1_LOC_106/A 0.01fF
C50428 INVX1_LOC_266/A INVX1_LOC_222/A 0.00fF
C50429 NAND2X1_LOC_573/Y NAND2X1_LOC_851/a_36_24# 0.00fF
C50430 INVX1_LOC_201/Y INVX1_LOC_267/Y 0.01fF
C50431 INVX1_LOC_217/A NOR2X1_LOC_528/a_36_216# 0.01fF
C50432 NOR2X1_LOC_15/Y INVX1_LOC_311/A 0.03fF
C50433 NOR2X1_LOC_641/a_36_216# NOR2X1_LOC_814/A 0.01fF
C50434 NOR2X1_LOC_67/A NOR2X1_LOC_690/A 0.09fF
C50435 INVX1_LOC_57/Y NAND2X1_LOC_861/Y 0.10fF
C50436 NOR2X1_LOC_82/A INVX1_LOC_75/A 0.11fF
C50437 NAND2X1_LOC_391/Y NOR2X1_LOC_45/B 0.07fF
C50438 INVX1_LOC_242/Y NAND2X1_LOC_463/B 0.01fF
C50439 INVX1_LOC_108/Y INVX1_LOC_2/Y 0.16fF
C50440 NOR2X1_LOC_209/Y INVX1_LOC_85/A 0.01fF
C50441 INVX1_LOC_27/A NOR2X1_LOC_562/B 0.10fF
C50442 VDD INVX1_LOC_53/A 2.81fF
C50443 INVX1_LOC_159/A INVX1_LOC_83/A 0.19fF
C50444 INVX1_LOC_33/A INVX1_LOC_56/Y 0.04fF
C50445 NOR2X1_LOC_272/Y NOR2X1_LOC_405/A 0.10fF
C50446 INVX1_LOC_62/Y NOR2X1_LOC_99/B 0.01fF
C50447 INVX1_LOC_41/A INVX1_LOC_53/Y 4.84fF
C50448 INVX1_LOC_304/Y INVX1_LOC_280/Y 0.51fF
C50449 NOR2X1_LOC_445/B INVX1_LOC_4/Y 0.75fF
C50450 INVX1_LOC_78/A INVX1_LOC_179/A 0.03fF
C50451 NAND2X1_LOC_471/Y INVX1_LOC_35/Y 0.01fF
C50452 NAND2X1_LOC_576/a_36_24# NOR2X1_LOC_45/B 0.00fF
C50453 INVX1_LOC_278/A INVX1_LOC_37/Y 0.01fF
C50454 INPUT_3 INPUT_0 0.10fF
C50455 NAND2X1_LOC_35/Y INVX1_LOC_37/A 0.01fF
C50456 INVX1_LOC_174/A NAND2X1_LOC_328/a_36_24# 0.00fF
C50457 INVX1_LOC_284/Y INVX1_LOC_282/A 0.02fF
C50458 NOR2X1_LOC_106/A INVX1_LOC_71/A 0.01fF
C50459 INVX1_LOC_104/A INVX1_LOC_16/A 0.14fF
C50460 INVX1_LOC_303/A D_INPUT_0 0.78fF
C50461 NOR2X1_LOC_717/B NOR2X1_LOC_550/B 0.03fF
C50462 INVX1_LOC_279/A NOR2X1_LOC_551/B 0.10fF
C50463 INVX1_LOC_145/A NAND2X1_LOC_105/a_36_24# 0.00fF
C50464 INVX1_LOC_255/Y NAND2X1_LOC_562/B 0.09fF
C50465 NAND2X1_LOC_856/A NAND2X1_LOC_863/A 0.01fF
C50466 NOR2X1_LOC_790/B INVX1_LOC_38/A 0.03fF
C50467 NAND2X1_LOC_363/B NOR2X1_LOC_536/A 0.42fF
C50468 NOR2X1_LOC_15/Y INVX1_LOC_304/A 0.07fF
C50469 NOR2X1_LOC_773/Y NOR2X1_LOC_190/a_36_216# 0.01fF
C50470 NAND2X1_LOC_338/B INVX1_LOC_218/A 0.15fF
C50471 D_INPUT_0 NOR2X1_LOC_672/Y 0.04fF
C50472 INVX1_LOC_214/A NAND2X1_LOC_840/B 0.01fF
C50473 NOR2X1_LOC_68/A NOR2X1_LOC_567/B 0.38fF
C50474 INVX1_LOC_310/A NOR2X1_LOC_516/B 0.09fF
C50475 NOR2X1_LOC_667/A NAND2X1_LOC_840/B 0.01fF
C50476 NOR2X1_LOC_242/A VDD 0.39fF
C50477 NOR2X1_LOC_92/Y NAND2X1_LOC_465/A 0.01fF
C50478 NAND2X1_LOC_276/Y INVX1_LOC_135/A 0.03fF
C50479 NOR2X1_LOC_860/Y NOR2X1_LOC_416/A 0.02fF
C50480 INVX1_LOC_248/A NAND2X1_LOC_840/B 0.01fF
C50481 NOR2X1_LOC_15/Y NOR2X1_LOC_670/Y 0.09fF
C50482 NAND2X1_LOC_565/a_36_24# NOR2X1_LOC_536/A 0.00fF
C50483 INVX1_LOC_228/Y INVX1_LOC_316/A 0.19fF
C50484 INVX1_LOC_17/A NOR2X1_LOC_346/Y 0.03fF
C50485 NAND2X1_LOC_392/A NAND2X1_LOC_850/Y 0.04fF
C50486 INVX1_LOC_15/Y NOR2X1_LOC_521/Y 0.03fF
C50487 NOR2X1_LOC_598/B NOR2X1_LOC_640/Y 0.76fF
C50488 NOR2X1_LOC_844/A NOR2X1_LOC_99/B 0.02fF
C50489 INVX1_LOC_23/A NAND2X1_LOC_798/B 0.07fF
C50490 INVX1_LOC_13/Y NAND2X1_LOC_848/A 0.03fF
C50491 INVX1_LOC_289/Y NAND2X1_LOC_453/A 0.05fF
C50492 NOR2X1_LOC_557/Y NAND2X1_LOC_842/B 0.43fF
C50493 INVX1_LOC_116/Y NOR2X1_LOC_814/A 0.08fF
C50494 INVX1_LOC_314/Y INVX1_LOC_73/A 0.00fF
C50495 NOR2X1_LOC_158/Y INVX1_LOC_19/A 0.07fF
C50496 INVX1_LOC_27/Y NOR2X1_LOC_39/Y 0.17fF
C50497 INVX1_LOC_263/A INVX1_LOC_16/A 0.01fF
C50498 INVX1_LOC_128/Y INVX1_LOC_29/A 0.01fF
C50499 INVX1_LOC_27/A INVX1_LOC_281/Y 0.01fF
C50500 NAND2X1_LOC_564/B NAND2X1_LOC_858/a_36_24# 0.00fF
C50501 NAND2X1_LOC_363/B NAND2X1_LOC_93/B 0.01fF
C50502 INVX1_LOC_12/A INVX1_LOC_4/Y 0.07fF
C50503 NOR2X1_LOC_123/B NOR2X1_LOC_709/A 0.76fF
C50504 INVX1_LOC_103/A NOR2X1_LOC_52/a_36_216# 0.01fF
C50505 INVX1_LOC_1/Y INVX1_LOC_22/A 0.69fF
C50506 INVX1_LOC_232/A NOR2X1_LOC_719/A 0.28fF
C50507 NAND2X1_LOC_350/A NAND2X1_LOC_469/B 0.03fF
C50508 INVX1_LOC_90/A NAND2X1_LOC_357/B 0.09fF
C50509 NOR2X1_LOC_791/B INVX1_LOC_123/A 0.12fF
C50510 NOR2X1_LOC_151/Y NOR2X1_LOC_550/B 0.10fF
C50511 NOR2X1_LOC_843/B INVX1_LOC_63/A 0.10fF
C50512 NOR2X1_LOC_468/Y NOR2X1_LOC_176/Y 0.01fF
C50513 NAND2X1_LOC_465/a_36_24# NAND2X1_LOC_99/A 0.00fF
C50514 INVX1_LOC_135/A NAND2X1_LOC_374/Y 0.10fF
C50515 NOR2X1_LOC_25/Y NOR2X1_LOC_11/Y 0.61fF
C50516 INVX1_LOC_25/A INVX1_LOC_285/A 0.07fF
C50517 INVX1_LOC_147/A NAND2X1_LOC_652/a_36_24# 0.01fF
C50518 INVX1_LOC_113/Y NOR2X1_LOC_74/Y 0.01fF
C50519 INVX1_LOC_28/A INVX1_LOC_104/A 0.17fF
C50520 INVX1_LOC_84/A INVX1_LOC_29/Y 0.06fF
C50521 INVX1_LOC_64/A NAND2X1_LOC_792/a_36_24# 0.00fF
C50522 NOR2X1_LOC_391/A NOR2X1_LOC_121/A 0.69fF
C50523 INVX1_LOC_55/Y INVX1_LOC_266/Y 0.09fF
C50524 INVX1_LOC_25/A NOR2X1_LOC_814/A 0.04fF
C50525 INVX1_LOC_7/A INVX1_LOC_232/A 0.52fF
C50526 INVX1_LOC_224/A INVX1_LOC_117/A 0.01fF
C50527 INVX1_LOC_165/A INVX1_LOC_42/A 0.01fF
C50528 NAND2X1_LOC_30/Y NAND2X1_LOC_51/a_36_24# 0.00fF
C50529 NAND2X1_LOC_350/A NOR2X1_LOC_447/B 0.01fF
C50530 NAND2X1_LOC_364/A NOR2X1_LOC_113/A 0.01fF
C50531 INVX1_LOC_90/A NAND2X1_LOC_549/B 0.01fF
C50532 NOR2X1_LOC_222/Y NOR2X1_LOC_214/B 0.00fF
C50533 INVX1_LOC_11/A INVX1_LOC_117/A 0.20fF
C50534 NOR2X1_LOC_163/A NAND2X1_LOC_451/Y 0.04fF
C50535 NAND2X1_LOC_364/A NOR2X1_LOC_405/A 2.21fF
C50536 NOR2X1_LOC_778/B NOR2X1_LOC_180/B 0.03fF
C50537 NOR2X1_LOC_510/Y INVX1_LOC_92/A 0.03fF
C50538 INVX1_LOC_13/Y INVX1_LOC_46/Y 1.01fF
C50539 NOR2X1_LOC_28/a_36_216# NOR2X1_LOC_38/B 0.03fF
C50540 NAND2X1_LOC_363/B INVX1_LOC_3/A 0.02fF
C50541 INVX1_LOC_255/Y NOR2X1_LOC_332/A 0.65fF
C50542 INVX1_LOC_25/Y NOR2X1_LOC_132/a_36_216# 0.00fF
C50543 NOR2X1_LOC_635/A NAND2X1_LOC_51/B 0.01fF
C50544 NAND2X1_LOC_165/a_36_24# NOR2X1_LOC_356/A 0.00fF
C50545 NAND2X1_LOC_725/B INVX1_LOC_118/A 3.11fF
C50546 NOR2X1_LOC_798/A NOR2X1_LOC_197/B 0.03fF
C50547 NOR2X1_LOC_160/B NAND2X1_LOC_96/A 0.07fF
C50548 NOR2X1_LOC_524/Y NAND2X1_LOC_211/Y 0.02fF
C50549 NOR2X1_LOC_336/B NOR2X1_LOC_857/A 0.01fF
C50550 NOR2X1_LOC_693/Y INVX1_LOC_42/A 0.34fF
C50551 NOR2X1_LOC_36/A D_INPUT_5 0.03fF
C50552 NOR2X1_LOC_561/Y NOR2X1_LOC_366/Y 0.03fF
C50553 INVX1_LOC_77/A NOR2X1_LOC_78/A 21.89fF
C50554 NOR2X1_LOC_220/A INVX1_LOC_182/A 0.10fF
C50555 INVX1_LOC_53/A INVX1_LOC_133/A 0.01fF
C50556 NAND2X1_LOC_324/a_36_24# INVX1_LOC_291/A 0.01fF
C50557 NAND2X1_LOC_197/a_36_24# NAND2X1_LOC_468/B 0.00fF
C50558 D_INPUT_0 INVX1_LOC_80/A 0.02fF
C50559 NOR2X1_LOC_328/Y NOR2X1_LOC_330/a_36_216# 0.00fF
C50560 NOR2X1_LOC_790/A NOR2X1_LOC_445/B 0.01fF
C50561 INVX1_LOC_58/A NOR2X1_LOC_89/A 1.63fF
C50562 NAND2X1_LOC_74/B INVX1_LOC_58/Y 0.07fF
C50563 NOR2X1_LOC_717/A INVX1_LOC_29/A 0.03fF
C50564 NOR2X1_LOC_594/Y NAND2X1_LOC_661/B 0.00fF
C50565 NAND2X1_LOC_656/Y NAND2X1_LOC_140/A 0.04fF
C50566 NOR2X1_LOC_500/B NOR2X1_LOC_859/Y 0.01fF
C50567 INVX1_LOC_30/A NAND2X1_LOC_639/A 0.06fF
C50568 NOR2X1_LOC_205/Y INVX1_LOC_307/A 0.73fF
C50569 INVX1_LOC_159/A INVX1_LOC_46/A 0.07fF
C50570 INVX1_LOC_72/A NAND2X1_LOC_472/Y 0.33fF
C50571 INVX1_LOC_49/A NAND2X1_LOC_468/B 0.03fF
C50572 INVX1_LOC_30/A NOR2X1_LOC_536/A 0.25fF
C50573 NOR2X1_LOC_742/A INVX1_LOC_22/A 0.07fF
C50574 INVX1_LOC_233/Y INVX1_LOC_12/A 0.04fF
C50575 NOR2X1_LOC_262/a_36_216# INVX1_LOC_47/Y 0.01fF
C50576 INVX1_LOC_89/A INVX1_LOC_120/A 0.03fF
C50577 NOR2X1_LOC_609/Y NOR2X1_LOC_383/B 0.01fF
C50578 INVX1_LOC_206/A NOR2X1_LOC_355/B 0.05fF
C50579 INVX1_LOC_124/A INVX1_LOC_98/A 0.04fF
C50580 INVX1_LOC_184/A VDD 0.12fF
C50581 INVX1_LOC_1/A INVX1_LOC_285/A 0.19fF
C50582 INVX1_LOC_162/Y NAND2X1_LOC_642/Y 0.00fF
C50583 NAND2X1_LOC_200/B INVX1_LOC_92/Y 0.03fF
C50584 INVX1_LOC_124/A NOR2X1_LOC_78/A 0.23fF
C50585 INVX1_LOC_230/Y NOR2X1_LOC_78/Y 0.03fF
C50586 INVX1_LOC_78/A NOR2X1_LOC_693/Y 0.24fF
C50587 INVX1_LOC_21/A INVX1_LOC_49/Y 0.03fF
C50588 NOR2X1_LOC_78/B NOR2X1_LOC_337/Y 0.02fF
C50589 INVX1_LOC_1/A NOR2X1_LOC_814/A 0.18fF
C50590 INVX1_LOC_120/A NAND2X1_LOC_508/A 0.08fF
C50591 NOR2X1_LOC_89/Y NAND2X1_LOC_99/A 0.01fF
C50592 INVX1_LOC_2/A NAND2X1_LOC_655/A 0.07fF
C50593 NOR2X1_LOC_335/B INVX1_LOC_101/A 0.00fF
C50594 NOR2X1_LOC_71/a_36_216# INVX1_LOC_53/Y 0.02fF
C50595 INVX1_LOC_72/A NAND2X1_LOC_637/Y 0.10fF
C50596 NOR2X1_LOC_647/Y NOR2X1_LOC_656/Y 0.18fF
C50597 NOR2X1_LOC_226/A NAND2X1_LOC_655/A 0.10fF
C50598 NOR2X1_LOC_724/Y NOR2X1_LOC_738/A 0.05fF
C50599 INVX1_LOC_30/A NAND2X1_LOC_93/B 0.07fF
C50600 INVX1_LOC_104/A NOR2X1_LOC_35/Y 0.10fF
C50601 NOR2X1_LOC_6/B INVX1_LOC_20/A 0.02fF
C50602 NOR2X1_LOC_303/Y INVX1_LOC_44/A 0.17fF
C50603 INVX1_LOC_256/A NAND2X1_LOC_475/Y 0.00fF
C50604 INVX1_LOC_2/A NAND2X1_LOC_468/B 0.04fF
C50605 INVX1_LOC_57/A NOR2X1_LOC_301/A 0.03fF
C50606 INVX1_LOC_34/A NAND2X1_LOC_804/Y 0.07fF
C50607 INVX1_LOC_50/A NOR2X1_LOC_318/A 0.03fF
C50608 NAND2X1_LOC_563/Y D_INPUT_3 1.11fF
C50609 NOR2X1_LOC_355/A NOR2X1_LOC_335/B 0.01fF
C50610 NAND2X1_LOC_45/Y NOR2X1_LOC_196/Y 0.02fF
C50611 NOR2X1_LOC_332/A NOR2X1_LOC_199/a_36_216# 0.01fF
C50612 INVX1_LOC_80/Y VDD 0.26fF
C50613 NOR2X1_LOC_318/B INVX1_LOC_22/A 0.02fF
C50614 NOR2X1_LOC_226/A NAND2X1_LOC_468/B 0.06fF
C50615 NOR2X1_LOC_357/Y INVX1_LOC_266/Y 0.05fF
C50616 NOR2X1_LOC_78/A NOR2X1_LOC_687/Y 0.03fF
C50617 INVX1_LOC_18/A NOR2X1_LOC_435/A 0.01fF
C50618 NOR2X1_LOC_672/Y NAND2X1_LOC_848/A 0.01fF
C50619 NOR2X1_LOC_602/A NOR2X1_LOC_841/A 0.02fF
C50620 NOR2X1_LOC_253/a_36_216# NOR2X1_LOC_693/Y 0.01fF
C50621 NOR2X1_LOC_703/B NOR2X1_LOC_862/B 0.02fF
C50622 INVX1_LOC_168/A NOR2X1_LOC_266/B 0.18fF
C50623 INVX1_LOC_78/A NOR2X1_LOC_405/Y 0.06fF
C50624 INVX1_LOC_51/Y NOR2X1_LOC_99/B 0.04fF
C50625 NAND2X1_LOC_712/A NOR2X1_LOC_45/B 0.01fF
C50626 NOR2X1_LOC_512/Y INVX1_LOC_291/A 0.01fF
C50627 GATE_579 INVX1_LOC_240/Y 0.01fF
C50628 NAND2X1_LOC_348/A NOR2X1_LOC_702/Y 0.03fF
C50629 INVX1_LOC_55/Y INVX1_LOC_42/Y 0.09fF
C50630 INVX1_LOC_161/Y INVX1_LOC_264/A 0.00fF
C50631 NOR2X1_LOC_205/Y INVX1_LOC_12/A 0.03fF
C50632 INVX1_LOC_298/Y NOR2X1_LOC_717/A 0.02fF
C50633 INVX1_LOC_93/Y INVX1_LOC_22/A 0.14fF
C50634 NOR2X1_LOC_344/A INVX1_LOC_38/A 0.08fF
C50635 NAND2X1_LOC_276/Y INVX1_LOC_280/A 0.07fF
C50636 NAND2X1_LOC_555/Y NOR2X1_LOC_662/A 0.00fF
C50637 NAND2X1_LOC_123/Y INVX1_LOC_73/A 1.71fF
C50638 NOR2X1_LOC_634/B VDD 0.05fF
C50639 NOR2X1_LOC_218/Y NAND2X1_LOC_468/B 0.16fF
C50640 INVX1_LOC_25/Y INVX1_LOC_59/Y 0.09fF
C50641 NOR2X1_LOC_542/Y NOR2X1_LOC_552/Y 0.09fF
C50642 NOR2X1_LOC_547/B VDD -0.00fF
C50643 NOR2X1_LOC_78/B VDD 1.52fF
C50644 NOR2X1_LOC_15/Y INVX1_LOC_19/Y 0.03fF
C50645 NOR2X1_LOC_705/a_36_216# NAND2X1_LOC_425/Y 0.01fF
C50646 NAND2X1_LOC_357/B INVX1_LOC_38/A 0.07fF
C50647 INVX1_LOC_232/A INVX1_LOC_76/A 1.27fF
C50648 INVX1_LOC_63/Y INVX1_LOC_54/A 0.31fF
C50649 INVX1_LOC_242/Y INVX1_LOC_42/A 0.01fF
C50650 INVX1_LOC_50/A NOR2X1_LOC_678/A 0.06fF
C50651 NOR2X1_LOC_647/Y INVX1_LOC_63/A 0.02fF
C50652 INVX1_LOC_5/A INVX1_LOC_16/Y 0.00fF
C50653 NOR2X1_LOC_353/Y INVX1_LOC_44/A 0.01fF
C50654 INVX1_LOC_113/Y INVX1_LOC_179/A 0.02fF
C50655 INVX1_LOC_259/A NOR2X1_LOC_684/Y 0.04fF
C50656 INVX1_LOC_22/A INVX1_LOC_139/A 0.01fF
C50657 INVX1_LOC_266/A INVX1_LOC_4/A 1.10fF
C50658 NOR2X1_LOC_730/a_36_216# NOR2X1_LOC_155/A 0.00fF
C50659 NAND2X1_LOC_364/Y NOR2X1_LOC_634/A 0.01fF
C50660 INVX1_LOC_30/Y INVX1_LOC_20/A 0.06fF
C50661 INVX1_LOC_18/A INVX1_LOC_63/A 3.87fF
C50662 INVX1_LOC_183/Y NOR2X1_LOC_45/B 0.07fF
C50663 NOR2X1_LOC_459/A NAND2X1_LOC_659/B 0.03fF
C50664 INVX1_LOC_72/A NAND2X1_LOC_773/B 0.01fF
C50665 NOR2X1_LOC_121/Y NOR2X1_LOC_99/Y 0.11fF
C50666 INVX1_LOC_24/A INVX1_LOC_119/Y 2.78fF
C50667 INVX1_LOC_153/Y INVX1_LOC_92/A 0.07fF
C50668 INVX1_LOC_83/A NOR2X1_LOC_56/Y 0.10fF
C50669 INVX1_LOC_11/A INVX1_LOC_3/Y 0.07fF
C50670 NOR2X1_LOC_738/a_36_216# INVX1_LOC_117/A 0.00fF
C50671 NAND2X1_LOC_721/A INVX1_LOC_22/A 0.10fF
C50672 INVX1_LOC_33/A NOR2X1_LOC_831/B 0.01fF
C50673 NAND2X1_LOC_53/Y D_INPUT_5 0.02fF
C50674 NOR2X1_LOC_666/A NAND2X1_LOC_454/Y 0.03fF
C50675 INVX1_LOC_71/A INVX1_LOC_294/A 0.27fF
C50676 VDD NAND2X1_LOC_392/Y 0.06fF
C50677 NOR2X1_LOC_516/B NAND2X1_LOC_96/A 0.10fF
C50678 NOR2X1_LOC_366/Y INVX1_LOC_76/A 0.01fF
C50679 INVX1_LOC_121/Y INVX1_LOC_92/A 0.02fF
C50680 INVX1_LOC_5/A NAND2X1_LOC_205/A 0.00fF
C50681 NOR2X1_LOC_723/Y INVX1_LOC_12/A 0.01fF
C50682 INVX1_LOC_225/Y INVX1_LOC_32/A 0.07fF
C50683 INVX1_LOC_49/A NOR2X1_LOC_66/Y 0.01fF
C50684 NOR2X1_LOC_322/Y NOR2X1_LOC_528/Y 0.27fF
C50685 INVX1_LOC_177/A INVX1_LOC_92/A 0.03fF
C50686 INVX1_LOC_311/A NOR2X1_LOC_733/Y 0.03fF
C50687 INVX1_LOC_83/A VDD 2.84fF
C50688 NOR2X1_LOC_816/A INVX1_LOC_21/Y 0.14fF
C50689 NAND2X1_LOC_430/a_36_24# NAND2X1_LOC_451/Y 0.00fF
C50690 INVX1_LOC_91/Y INVX1_LOC_91/A 0.01fF
C50691 NAND2X1_LOC_630/a_36_24# INVX1_LOC_92/A 0.00fF
C50692 NOR2X1_LOC_91/Y INVX1_LOC_102/A 0.02fF
C50693 NOR2X1_LOC_510/Y INVX1_LOC_53/A 0.10fF
C50694 NAND2X1_LOC_112/Y INVX1_LOC_9/A 0.01fF
C50695 NAND2X1_LOC_198/B INVX1_LOC_168/Y 0.01fF
C50696 NOR2X1_LOC_67/A NOR2X1_LOC_88/a_36_216# 0.01fF
C50697 NOR2X1_LOC_419/Y NAND2X1_LOC_74/B 0.10fF
C50698 INVX1_LOC_64/A INVX1_LOC_50/Y 0.07fF
C50699 INVX1_LOC_1/A NAND2X1_LOC_40/a_36_24# 0.00fF
C50700 INVX1_LOC_75/A INVX1_LOC_59/Y 0.05fF
C50701 NOR2X1_LOC_45/B INVX1_LOC_309/A 0.03fF
C50702 NAND2X1_LOC_162/A INVX1_LOC_92/A 0.02fF
C50703 INVX1_LOC_267/A NAND2X1_LOC_659/A 0.00fF
C50704 INVX1_LOC_93/Y INVX1_LOC_100/A 0.02fF
C50705 NOR2X1_LOC_716/B NAND2X1_LOC_74/B 0.20fF
C50706 NOR2X1_LOC_32/B INVX1_LOC_59/A 0.02fF
C50707 NAND2X1_LOC_656/Y INVX1_LOC_118/Y 0.04fF
C50708 INVX1_LOC_22/A INVX1_LOC_117/Y 0.03fF
C50709 INVX1_LOC_2/A NOR2X1_LOC_66/Y 0.03fF
C50710 INVX1_LOC_45/A NOR2X1_LOC_334/Y 0.09fF
C50711 INPUT_0 NOR2X1_LOC_332/B 0.06fF
C50712 INVX1_LOC_17/A INVX1_LOC_57/A 0.14fF
C50713 INVX1_LOC_30/A NAND2X1_LOC_470/B 0.10fF
C50714 NOR2X1_LOC_160/B NAND2X1_LOC_99/A 0.44fF
C50715 NOR2X1_LOC_818/Y NOR2X1_LOC_820/B 0.04fF
C50716 NOR2X1_LOC_537/Y NAND2X1_LOC_206/Y 0.07fF
C50717 NOR2X1_LOC_329/B INVX1_LOC_12/Y 0.03fF
C50718 INVX1_LOC_136/A NOR2X1_LOC_394/Y 0.03fF
C50719 NOR2X1_LOC_357/Y INVX1_LOC_42/Y 0.04fF
C50720 INVX1_LOC_34/Y INVX1_LOC_63/A 0.15fF
C50721 NOR2X1_LOC_45/B INVX1_LOC_91/A 0.24fF
C50722 INVX1_LOC_43/Y NOR2X1_LOC_72/Y 0.02fF
C50723 NOR2X1_LOC_361/B INVX1_LOC_53/A 0.58fF
C50724 NOR2X1_LOC_34/B NOR2X1_LOC_249/Y 0.00fF
C50725 INVX1_LOC_216/Y INVX1_LOC_23/A 0.00fF
C50726 INVX1_LOC_58/A INVX1_LOC_11/A 0.19fF
C50727 NOR2X1_LOC_321/Y NOR2X1_LOC_109/Y 0.02fF
C50728 NOR2X1_LOC_846/Y INVX1_LOC_27/A 0.03fF
C50729 INVX1_LOC_35/A INVX1_LOC_269/A 0.11fF
C50730 NOR2X1_LOC_381/Y INVX1_LOC_64/A 0.13fF
C50731 NAND2X1_LOC_559/Y NAND2X1_LOC_35/Y 0.07fF
C50732 NOR2X1_LOC_6/B NOR2X1_LOC_128/A 0.06fF
C50733 INVX1_LOC_144/A INVX1_LOC_37/A 0.05fF
C50734 NAND2X1_LOC_338/B NAND2X1_LOC_773/B 0.11fF
C50735 NAND2X1_LOC_581/a_36_24# INVX1_LOC_11/A 0.00fF
C50736 NOR2X1_LOC_276/B NAND2X1_LOC_454/Y 0.02fF
C50737 NOR2X1_LOC_45/B INVX1_LOC_11/Y 0.03fF
C50738 NOR2X1_LOC_474/A INVX1_LOC_3/Y 0.01fF
C50739 NOR2X1_LOC_113/A NOR2X1_LOC_405/A 0.02fF
C50740 NOR2X1_LOC_647/A INVX1_LOC_36/A 0.33fF
C50741 INVX1_LOC_247/A INVX1_LOC_91/A 0.05fF
C50742 INPUT_0 NAND2X1_LOC_804/Y 0.07fF
C50743 NOR2X1_LOC_78/B INVX1_LOC_133/A 0.07fF
C50744 NOR2X1_LOC_667/A INVX1_LOC_49/Y 0.00fF
C50745 NAND2X1_LOC_778/Y NAND2X1_LOC_778/a_36_24# 0.02fF
C50746 INVX1_LOC_71/A NOR2X1_LOC_334/Y 0.14fF
C50747 INVX1_LOC_72/A NOR2X1_LOC_639/Y 0.02fF
C50748 NOR2X1_LOC_730/B INVX1_LOC_37/A 0.02fF
C50749 INVX1_LOC_94/A NAND2X1_LOC_72/B 0.01fF
C50750 NOR2X1_LOC_68/A INVX1_LOC_26/A 0.04fF
C50751 INVX1_LOC_186/A INVX1_LOC_76/A 0.05fF
C50752 INVX1_LOC_101/A INVX1_LOC_84/A 0.01fF
C50753 NOR2X1_LOC_533/Y NOR2X1_LOC_304/Y 0.02fF
C50754 NAND2X1_LOC_161/a_36_24# INVX1_LOC_78/A 0.00fF
C50755 NOR2X1_LOC_817/Y INVX1_LOC_5/A 0.02fF
C50756 INVX1_LOC_11/A INVX1_LOC_248/Y 0.01fF
C50757 NOR2X1_LOC_526/Y INVX1_LOC_12/A 0.02fF
C50758 NOR2X1_LOC_473/B NOR2X1_LOC_216/B 0.01fF
C50759 NOR2X1_LOC_52/B INVX1_LOC_3/Y 0.01fF
C50760 INVX1_LOC_155/A INVX1_LOC_94/Y 0.04fF
C50761 NOR2X1_LOC_65/B INVX1_LOC_45/Y 0.30fF
C50762 NOR2X1_LOC_311/Y VDD 0.34fF
C50763 INVX1_LOC_233/A INVX1_LOC_286/Y -0.04fF
C50764 INVX1_LOC_13/A INVX1_LOC_19/A 0.28fF
C50765 NAND2X1_LOC_662/Y NOR2X1_LOC_48/Y 0.03fF
C50766 NOR2X1_LOC_6/B INVX1_LOC_4/A 0.02fF
C50767 NOR2X1_LOC_124/A INVX1_LOC_20/A 0.00fF
C50768 NOR2X1_LOC_355/A INVX1_LOC_84/A 0.00fF
C50769 INPUT_1 NAND2X1_LOC_141/Y 0.12fF
C50770 INVX1_LOC_266/Y INVX1_LOC_32/A 0.13fF
C50771 INVX1_LOC_89/A NAND2X1_LOC_659/A 0.20fF
C50772 NOR2X1_LOC_658/a_36_216# NOR2X1_LOC_208/Y 0.01fF
C50773 NOR2X1_LOC_527/a_36_216# INVX1_LOC_185/A 0.00fF
C50774 NAND2X1_LOC_579/A NAND2X1_LOC_575/a_36_24# 0.02fF
C50775 NAND2X1_LOC_348/A NOR2X1_LOC_78/a_36_216# 0.00fF
C50776 NOR2X1_LOC_246/A NOR2X1_LOC_653/Y 0.11fF
C50777 NOR2X1_LOC_74/A NOR2X1_LOC_612/Y 0.01fF
C50778 INVX1_LOC_136/A INVX1_LOC_58/Y 0.36fF
C50779 INVX1_LOC_13/Y NOR2X1_LOC_134/Y 0.41fF
C50780 NAND2X1_LOC_565/B INVX1_LOC_284/A 0.02fF
C50781 NOR2X1_LOC_655/B INVX1_LOC_251/A 0.06fF
C50782 NOR2X1_LOC_421/a_36_216# INVX1_LOC_209/Y 0.00fF
C50783 NOR2X1_LOC_187/Y NAND2X1_LOC_190/Y 0.05fF
C50784 INVX1_LOC_223/Y INVX1_LOC_292/A 0.00fF
C50785 INVX1_LOC_200/Y NOR2X1_LOC_238/Y 0.02fF
C50786 NAND2X1_LOC_811/Y NAND2X1_LOC_175/Y 0.07fF
C50787 VDD NOR2X1_LOC_164/Y 0.12fF
C50788 VDD NOR2X1_LOC_368/Y 0.12fF
C50789 INVX1_LOC_255/Y NOR2X1_LOC_847/A 0.02fF
C50790 NOR2X1_LOC_758/Y NOR2X1_LOC_278/Y 0.09fF
C50791 NOR2X1_LOC_636/A NOR2X1_LOC_635/B 0.01fF
C50792 NOR2X1_LOC_794/a_36_216# NOR2X1_LOC_383/B 0.00fF
C50793 NAND2X1_LOC_338/B NOR2X1_LOC_393/Y 0.02fF
C50794 INVX1_LOC_233/Y INVX1_LOC_217/A 0.10fF
C50795 NOR2X1_LOC_246/A INVX1_LOC_19/A 0.07fF
C50796 NAND2X1_LOC_555/Y INVX1_LOC_252/A 0.03fF
C50797 NOR2X1_LOC_604/Y INVX1_LOC_24/A 0.01fF
C50798 NOR2X1_LOC_262/Y INVX1_LOC_29/Y 0.09fF
C50799 INVX1_LOC_199/A INVX1_LOC_117/A 0.05fF
C50800 INVX1_LOC_91/A NOR2X1_LOC_378/Y 0.00fF
C50801 NOR2X1_LOC_454/Y NOR2X1_LOC_45/Y 0.06fF
C50802 NAND2X1_LOC_109/a_36_24# NAND2X1_LOC_96/A 0.00fF
C50803 INVX1_LOC_6/A NOR2X1_LOC_433/Y 0.01fF
C50804 NOR2X1_LOC_391/a_36_216# NOR2X1_LOC_78/Y 0.00fF
C50805 INVX1_LOC_58/A NOR2X1_LOC_433/A 0.21fF
C50806 INVX1_LOC_285/Y INVX1_LOC_92/A 0.07fF
C50807 NOR2X1_LOC_78/A INVX1_LOC_9/A 4.77fF
C50808 NAND2X1_LOC_551/A INVX1_LOC_19/A 0.14fF
C50809 VDD INVX1_LOC_46/A 1.47fF
C50810 NOR2X1_LOC_120/a_36_216# INVX1_LOC_293/Y 0.00fF
C50811 NOR2X1_LOC_566/Y INVX1_LOC_4/Y 0.06fF
C50812 NAND2X1_LOC_703/Y INVX1_LOC_286/Y 0.04fF
C50813 INVX1_LOC_58/A NOR2X1_LOC_593/Y 0.27fF
C50814 NAND2X1_LOC_655/A INVX1_LOC_118/A 0.10fF
C50815 NOR2X1_LOC_130/A INVX1_LOC_284/A 0.07fF
C50816 NOR2X1_LOC_590/A INVX1_LOC_1/A 0.79fF
C50817 INVX1_LOC_36/A D_INPUT_6 0.01fF
C50818 NOR2X1_LOC_264/Y NOR2X1_LOC_621/a_36_216# 0.00fF
C50819 NOR2X1_LOC_346/B INVX1_LOC_87/A 0.01fF
C50820 INVX1_LOC_36/A NOR2X1_LOC_173/Y 0.10fF
C50821 NOR2X1_LOC_175/B INVX1_LOC_87/A 0.01fF
C50822 INVX1_LOC_151/Y INVX1_LOC_128/Y 0.05fF
C50823 INVX1_LOC_11/A INVX1_LOC_215/Y 0.21fF
C50824 NOR2X1_LOC_71/Y INVX1_LOC_42/A 0.03fF
C50825 INVX1_LOC_21/A INVX1_LOC_79/Y 0.01fF
C50826 NOR2X1_LOC_790/B INVX1_LOC_33/A 0.00fF
C50827 INVX1_LOC_30/Y INVX1_LOC_4/A 0.12fF
C50828 NOR2X1_LOC_742/A INVX1_LOC_186/Y 0.01fF
C50829 NOR2X1_LOC_454/Y NOR2X1_LOC_584/a_36_216# 0.01fF
C50830 VDD NOR2X1_LOC_766/Y 0.32fF
C50831 NOR2X1_LOC_188/A NOR2X1_LOC_814/A 0.14fF
C50832 INVX1_LOC_216/Y INVX1_LOC_31/A 0.01fF
C50833 INVX1_LOC_58/A NOR2X1_LOC_52/B 0.54fF
C50834 NAND2X1_LOC_327/a_36_24# INVX1_LOC_49/Y 0.00fF
C50835 INVX1_LOC_22/A INVX1_LOC_87/A 0.06fF
C50836 NOR2X1_LOC_76/A INVX1_LOC_170/Y 0.00fF
C50837 INVX1_LOC_191/Y NOR2X1_LOC_651/a_36_216# 0.00fF
C50838 NOR2X1_LOC_763/Y NOR2X1_LOC_467/A 0.91fF
C50839 NOR2X1_LOC_548/B NOR2X1_LOC_814/A 0.10fF
C50840 INVX1_LOC_69/Y NAND2X1_LOC_475/Y 0.03fF
C50841 NOR2X1_LOC_68/A NOR2X1_LOC_560/a_36_216# 0.00fF
C50842 NOR2X1_LOC_598/B NOR2X1_LOC_799/a_36_216# 0.01fF
C50843 NOR2X1_LOC_590/A NOR2X1_LOC_794/B 0.03fF
C50844 NOR2X1_LOC_186/Y INVX1_LOC_77/A 0.08fF
C50845 NOR2X1_LOC_2/Y NOR2X1_LOC_36/B 0.40fF
C50846 INVX1_LOC_233/A INVX1_LOC_185/Y 0.01fF
C50847 INVX1_LOC_75/A NOR2X1_LOC_340/A 0.10fF
C50848 INVX1_LOC_64/A NOR2X1_LOC_6/B 0.41fF
C50849 INVX1_LOC_5/A NOR2X1_LOC_570/B 0.00fF
C50850 INVX1_LOC_177/A INVX1_LOC_53/A 0.09fF
C50851 INVX1_LOC_256/A INVX1_LOC_30/A 0.20fF
C50852 NOR2X1_LOC_91/A NOR2X1_LOC_328/Y 0.01fF
C50853 INVX1_LOC_58/A NOR2X1_LOC_603/a_36_216# 0.00fF
C50854 INVX1_LOC_36/A NAND2X1_LOC_793/Y 0.11fF
C50855 INVX1_LOC_143/A NAND2X1_LOC_275/a_36_24# 0.00fF
C50856 INVX1_LOC_304/Y INVX1_LOC_233/Y 0.07fF
C50857 NOR2X1_LOC_808/A NOR2X1_LOC_598/B 0.02fF
C50858 INVX1_LOC_13/A INVX1_LOC_26/Y 0.07fF
C50859 NOR2X1_LOC_187/Y NOR2X1_LOC_596/A 0.06fF
C50860 NOR2X1_LOC_45/Y NAND2X1_LOC_196/a_36_24# 0.00fF
C50861 D_INPUT_1 NAND2X1_LOC_672/B 0.02fF
C50862 NOR2X1_LOC_45/B INVX1_LOC_203/A 0.08fF
C50863 INVX1_LOC_21/A INVX1_LOC_34/A 0.06fF
C50864 NOR2X1_LOC_479/B INVX1_LOC_23/A 0.01fF
C50865 NOR2X1_LOC_632/Y NOR2X1_LOC_383/B 0.03fF
C50866 NOR2X1_LOC_523/A NOR2X1_LOC_860/B 0.01fF
C50867 INVX1_LOC_2/A NOR2X1_LOC_772/B 0.01fF
C50868 NAND2X1_LOC_34/a_36_24# INVX1_LOC_64/A 0.00fF
C50869 INVX1_LOC_289/Y NOR2X1_LOC_577/Y 0.07fF
C50870 NOR2X1_LOC_705/B NOR2X1_LOC_546/A 0.02fF
C50871 NOR2X1_LOC_756/Y NOR2X1_LOC_38/B 0.38fF
C50872 INVX1_LOC_201/Y INVX1_LOC_235/Y 0.17fF
C50873 NOR2X1_LOC_155/A INVX1_LOC_37/A 0.07fF
C50874 NOR2X1_LOC_167/Y NOR2X1_LOC_46/a_36_216# 0.00fF
C50875 INVX1_LOC_124/A NOR2X1_LOC_186/Y 0.04fF
C50876 NAND2X1_LOC_218/B NOR2X1_LOC_82/A 0.01fF
C50877 INVX1_LOC_232/Y NOR2X1_LOC_662/a_36_216# 0.00fF
C50878 INVX1_LOC_88/A INVX1_LOC_49/A 0.03fF
C50879 INVX1_LOC_52/Y NOR2X1_LOC_142/Y -0.00fF
C50880 INVX1_LOC_292/A NAND2X1_LOC_167/a_36_24# 0.00fF
C50881 NOR2X1_LOC_226/A NOR2X1_LOC_772/B 0.07fF
C50882 NOR2X1_LOC_644/A INVX1_LOC_78/A 0.03fF
C50883 INVX1_LOC_2/A INVX1_LOC_13/Y 0.03fF
C50884 NOR2X1_LOC_160/B NAND2X1_LOC_656/A 0.02fF
C50885 NAND2X1_LOC_347/B NOR2X1_LOC_392/B 0.03fF
C50886 NOR2X1_LOC_226/A INVX1_LOC_13/Y 0.10fF
C50887 INVX1_LOC_90/A NOR2X1_LOC_282/Y 0.03fF
C50888 INVX1_LOC_36/A INVX1_LOC_205/A 0.01fF
C50889 INVX1_LOC_85/Y NOR2X1_LOC_308/a_36_216# 0.00fF
C50890 INVX1_LOC_21/A NAND2X1_LOC_231/Y 0.01fF
C50891 GATE_741 NAND2X1_LOC_717/Y 0.03fF
C50892 NOR2X1_LOC_405/A NOR2X1_LOC_841/a_36_216# 0.01fF
C50893 D_GATE_741 INVX1_LOC_33/A 0.12fF
C50894 NAND2X1_LOC_573/A INVX1_LOC_53/A 0.71fF
C50895 NOR2X1_LOC_643/Y INPUT_3 0.04fF
C50896 NAND2X1_LOC_30/Y NAND2X1_LOC_59/B 2.34fF
C50897 NOR2X1_LOC_538/B NOR2X1_LOC_264/Y 0.02fF
C50898 NOR2X1_LOC_788/B NOR2X1_LOC_383/B 0.00fF
C50899 NOR2X1_LOC_798/A NOR2X1_LOC_568/a_36_216# 0.00fF
C50900 NAND2X1_LOC_623/B NAND2X1_LOC_254/Y 0.09fF
C50901 INVX1_LOC_139/A INVX1_LOC_186/Y 0.19fF
C50902 VDD NOR2X1_LOC_68/Y 0.13fF
C50903 NOR2X1_LOC_178/Y NOR2X1_LOC_383/Y 0.16fF
C50904 NOR2X1_LOC_357/Y INVX1_LOC_19/A 0.01fF
C50905 NAND2X1_LOC_350/A INVX1_LOC_63/Y 0.27fF
C50906 INVX1_LOC_245/Y NOR2X1_LOC_770/B 0.01fF
C50907 INVX1_LOC_24/A INVX1_LOC_72/A 0.06fF
C50908 NOR2X1_LOC_202/a_36_216# INVX1_LOC_96/Y 0.00fF
C50909 NOR2X1_LOC_254/A NOR2X1_LOC_254/Y 0.02fF
C50910 NOR2X1_LOC_743/a_36_216# NAND2X1_LOC_352/B 0.02fF
C50911 NOR2X1_LOC_309/Y NAND2X1_LOC_793/Y 0.08fF
C50912 NOR2X1_LOC_346/Y NOR2X1_LOC_346/A 0.00fF
C50913 INVX1_LOC_157/Y NOR2X1_LOC_155/A -0.00fF
C50914 INVX1_LOC_2/A INVX1_LOC_88/A 0.10fF
C50915 INVX1_LOC_133/A INVX1_LOC_46/A 0.01fF
C50916 NOR2X1_LOC_82/A NOR2X1_LOC_84/a_36_216# 0.00fF
C50917 INVX1_LOC_33/A INVX1_LOC_81/Y 0.01fF
C50918 NOR2X1_LOC_67/A INVX1_LOC_14/A 0.24fF
C50919 NOR2X1_LOC_635/A INVX1_LOC_174/A 0.05fF
C50920 INVX1_LOC_49/A NOR2X1_LOC_500/B 0.02fF
C50921 INVX1_LOC_215/Y NOR2X1_LOC_52/B 0.07fF
C50922 NAND2X1_LOC_633/Y NAND2X1_LOC_74/B 0.07fF
C50923 NOR2X1_LOC_361/B NOR2X1_LOC_78/B 0.22fF
C50924 INVX1_LOC_255/Y NOR2X1_LOC_655/a_36_216# 0.01fF
C50925 NOR2X1_LOC_226/A INVX1_LOC_88/A 0.00fF
C50926 NOR2X1_LOC_524/Y INVX1_LOC_155/A 0.15fF
C50927 NOR2X1_LOC_155/A NOR2X1_LOC_743/Y 0.01fF
C50928 NAND2X1_LOC_549/Y INVX1_LOC_90/A 0.01fF
C50929 VDD NOR2X1_LOC_671/Y 0.60fF
C50930 INVX1_LOC_161/Y INVX1_LOC_236/A 0.12fF
C50931 NOR2X1_LOC_186/Y NAND2X1_LOC_796/Y 0.02fF
C50932 INVX1_LOC_249/A NOR2X1_LOC_457/B -0.01fF
C50933 INVX1_LOC_269/A INVX1_LOC_305/Y 0.02fF
C50934 INVX1_LOC_6/A NOR2X1_LOC_693/a_36_216# 0.00fF
C50935 NOR2X1_LOC_92/Y INVX1_LOC_16/A 3.63fF
C50936 INVX1_LOC_136/A NOR2X1_LOC_716/B 0.17fF
C50937 INVX1_LOC_73/A INVX1_LOC_271/A 0.03fF
C50938 NOR2X1_LOC_657/a_36_216# NOR2X1_LOC_561/Y 0.01fF
C50939 INVX1_LOC_66/Y INVX1_LOC_19/A 0.01fF
C50940 NOR2X1_LOC_557/Y INVX1_LOC_72/A 0.31fF
C50941 INVX1_LOC_289/Y INVX1_LOC_22/A 0.01fF
C50942 NOR2X1_LOC_433/A NOR2X1_LOC_338/Y -0.01fF
C50943 NAND2X1_LOC_514/Y NOR2X1_LOC_577/Y 0.01fF
C50944 NOR2X1_LOC_510/Y INVX1_LOC_83/A 0.10fF
C50945 NAND2X1_LOC_192/B INVX1_LOC_208/A 0.06fF
C50946 INVX1_LOC_269/A NOR2X1_LOC_121/A 0.10fF
C50947 NOR2X1_LOC_218/Y INVX1_LOC_88/A 0.01fF
C50948 NAND2X1_LOC_96/A NAND2X1_LOC_207/B 0.02fF
C50949 NAND2X1_LOC_725/B NAND2X1_LOC_735/B 0.03fF
C50950 INVX1_LOC_200/A NAND2X1_LOC_862/A 0.04fF
C50951 NOR2X1_LOC_238/Y NOR2X1_LOC_495/Y 0.05fF
C50952 NAND2X1_LOC_149/Y INVX1_LOC_121/A 0.04fF
C50953 NOR2X1_LOC_15/Y NOR2X1_LOC_589/A 0.04fF
C50954 NAND2X1_LOC_573/Y NAND2X1_LOC_796/Y 0.01fF
C50955 NOR2X1_LOC_222/Y NOR2X1_LOC_160/B 0.03fF
C50956 INVX1_LOC_269/A NOR2X1_LOC_188/Y 0.03fF
C50957 INVX1_LOC_13/Y INPUT_1 0.09fF
C50958 NOR2X1_LOC_82/A INVX1_LOC_22/A 0.02fF
C50959 NAND2X1_LOC_332/Y NOR2X1_LOC_351/a_36_216# 0.00fF
C50960 NOR2X1_LOC_361/B NAND2X1_LOC_392/Y 0.05fF
C50961 INVX1_LOC_132/A INVX1_LOC_77/A 0.14fF
C50962 INVX1_LOC_232/Y NOR2X1_LOC_514/A 0.24fF
C50963 INVX1_LOC_303/A INVX1_LOC_49/A 0.07fF
C50964 NAND2X1_LOC_9/Y NOR2X1_LOC_721/Y 0.03fF
C50965 INVX1_LOC_135/A NOR2X1_LOC_140/A 0.07fF
C50966 INVX1_LOC_230/Y INVX1_LOC_172/Y 0.01fF
C50967 NOR2X1_LOC_763/Y INVX1_LOC_1/A 0.03fF
C50968 NOR2X1_LOC_481/A INVX1_LOC_77/A 0.20fF
C50969 NOR2X1_LOC_111/A INVX1_LOC_15/A 0.07fF
C50970 NOR2X1_LOC_541/Y NOR2X1_LOC_569/Y 0.01fF
C50971 INVX1_LOC_285/Y INVX1_LOC_53/A 0.10fF
C50972 NOR2X1_LOC_780/B INVX1_LOC_89/A 0.01fF
C50973 INVX1_LOC_208/Y NOR2X1_LOC_389/A 0.13fF
C50974 INVX1_LOC_20/A INVX1_LOC_273/A 0.92fF
C50975 NOR2X1_LOC_15/Y INVX1_LOC_171/A 0.06fF
C50976 INVX1_LOC_136/A INVX1_LOC_98/Y 0.05fF
C50977 INVX1_LOC_143/A INVX1_LOC_72/A 0.05fF
C50978 INVX1_LOC_135/A NAND2X1_LOC_538/Y 0.10fF
C50979 INVX1_LOC_90/A NAND2X1_LOC_347/B 0.64fF
C50980 NAND2X1_LOC_59/B INVX1_LOC_49/A 0.12fF
C50981 NOR2X1_LOC_216/Y NOR2X1_LOC_674/Y 0.33fF
C50982 INVX1_LOC_30/Y INVX1_LOC_43/Y 0.00fF
C50983 NOR2X1_LOC_718/B INVX1_LOC_71/A 0.07fF
C50984 NOR2X1_LOC_640/Y INVX1_LOC_29/A 0.07fF
C50985 NAND2X1_LOC_332/Y NOR2X1_LOC_577/Y 0.03fF
C50986 INVX1_LOC_93/A NOR2X1_LOC_322/Y 0.10fF
C50987 NOR2X1_LOC_817/Y NOR2X1_LOC_332/A 0.03fF
C50988 INVX1_LOC_225/A INVX1_LOC_77/A 0.07fF
C50989 INVX1_LOC_33/A NOR2X1_LOC_344/A 0.02fF
C50990 INVX1_LOC_83/Y INVX1_LOC_142/A 0.01fF
C50991 NAND2X1_LOC_500/Y INVX1_LOC_22/A 0.04fF
C50992 NOR2X1_LOC_92/Y INVX1_LOC_28/A 2.12fF
C50993 NOR2X1_LOC_67/A NOR2X1_LOC_522/Y 0.04fF
C50994 INVX1_LOC_24/A NOR2X1_LOC_537/Y 0.03fF
C50995 NOR2X1_LOC_142/Y INVX1_LOC_63/Y 0.31fF
C50996 NAND2X1_LOC_30/Y NAND2X1_LOC_1/a_36_24# 0.00fF
C50997 INVX1_LOC_24/A NAND2X1_LOC_338/B 0.19fF
C50998 NAND2X1_LOC_243/Y INVX1_LOC_42/A 0.19fF
C50999 NOR2X1_LOC_716/B NOR2X1_LOC_278/A 0.04fF
C51000 INVX1_LOC_78/A NAND2X1_LOC_284/a_36_24# 0.00fF
C51001 INVX1_LOC_89/Y INVX1_LOC_42/A 0.02fF
C51002 NOR2X1_LOC_295/a_36_216# NOR2X1_LOC_295/Y 0.03fF
C51003 INVX1_LOC_58/A INVX1_LOC_199/A 0.07fF
C51004 NAND2X1_LOC_85/Y INVX1_LOC_29/A 0.43fF
C51005 NOR2X1_LOC_136/Y NAND2X1_LOC_198/B 0.05fF
C51006 INVX1_LOC_21/A INPUT_0 0.23fF
C51007 INVX1_LOC_2/A INVX1_LOC_303/A 0.10fF
C51008 NOR2X1_LOC_209/Y INVX1_LOC_77/A 0.03fF
C51009 INVX1_LOC_226/Y NOR2X1_LOC_360/Y 0.07fF
C51010 INVX1_LOC_65/A INVX1_LOC_53/A 0.09fF
C51011 NOR2X1_LOC_440/Y INVX1_LOC_30/A -0.01fF
C51012 INVX1_LOC_18/A INVX1_LOC_1/Y 1.73fF
C51013 NOR2X1_LOC_481/A INVX1_LOC_124/A 0.02fF
C51014 NAND2X1_LOC_198/B INVX1_LOC_56/A 0.02fF
C51015 INVX1_LOC_255/Y NOR2X1_LOC_554/B 0.01fF
C51016 INVX1_LOC_221/A NAND2X1_LOC_354/B 0.02fF
C51017 INVX1_LOC_223/A NOR2X1_LOC_543/A 0.01fF
C51018 NAND2X1_LOC_543/Y NOR2X1_LOC_91/Y 0.15fF
C51019 NAND2X1_LOC_796/B NOR2X1_LOC_167/Y 0.07fF
C51020 NAND2X1_LOC_181/Y INVX1_LOC_314/Y 0.04fF
C51021 NAND2X1_LOC_569/A NOR2X1_LOC_315/Y 0.00fF
C51022 NOR2X1_LOC_226/A INVX1_LOC_303/A 1.22fF
C51023 NOR2X1_LOC_334/Y NOR2X1_LOC_331/B 0.01fF
C51024 INVX1_LOC_128/Y INVX1_LOC_118/Y 0.01fF
C51025 INVX1_LOC_53/A NOR2X1_LOC_137/B 0.01fF
C51026 NAND2X1_LOC_361/Y INVX1_LOC_196/A 0.07fF
C51027 NOR2X1_LOC_617/Y INVX1_LOC_197/Y 0.00fF
C51028 NOR2X1_LOC_516/B NAND2X1_LOC_656/A 0.03fF
C51029 NOR2X1_LOC_434/Y INVX1_LOC_186/A 0.07fF
C51030 INVX1_LOC_124/A INVX1_LOC_225/A 0.03fF
C51031 NOR2X1_LOC_526/Y NAND2X1_LOC_787/B 0.07fF
C51032 INVX1_LOC_64/A NOR2X1_LOC_124/A 0.02fF
C51033 INVX1_LOC_103/A INVX1_LOC_75/A 0.10fF
C51034 NOR2X1_LOC_91/A INVX1_LOC_33/Y 0.01fF
C51035 NAND2X1_LOC_725/A NOR2X1_LOC_396/Y 0.01fF
C51036 INVX1_LOC_64/A INVX1_LOC_188/Y 0.01fF
C51037 NOR2X1_LOC_498/Y NAND2X1_LOC_717/Y 0.05fF
C51038 D_INPUT_1 INVX1_LOC_2/Y 0.03fF
C51039 NOR2X1_LOC_274/Y INVX1_LOC_232/A 0.21fF
C51040 INVX1_LOC_72/A NAND2X1_LOC_800/Y 0.05fF
C51041 INVX1_LOC_136/A NOR2X1_LOC_717/B 0.03fF
C51042 NOR2X1_LOC_89/A NAND2X1_LOC_475/Y 0.01fF
C51043 NOR2X1_LOC_78/B INVX1_LOC_153/Y 0.90fF
C51044 NOR2X1_LOC_160/B NOR2X1_LOC_329/B 0.10fF
C51045 INVX1_LOC_34/A NOR2X1_LOC_667/A 0.03fF
C51046 NOR2X1_LOC_769/B INVX1_LOC_37/A 0.01fF
C51047 NOR2X1_LOC_226/A NAND2X1_LOC_734/a_36_24# 0.01fF
C51048 NOR2X1_LOC_569/Y INVX1_LOC_71/A 0.07fF
C51049 NOR2X1_LOC_602/A INVX1_LOC_90/A 0.09fF
C51050 INVX1_LOC_256/Y INVX1_LOC_8/A 0.04fF
C51051 INVX1_LOC_32/A NAND2X1_LOC_288/A 0.10fF
C51052 INVX1_LOC_129/Y INVX1_LOC_129/A 0.02fF
C51053 NAND2X1_LOC_35/Y NAND2X1_LOC_465/A 0.01fF
C51054 INVX1_LOC_4/Y INVX1_LOC_92/A 0.17fF
C51055 NAND2X1_LOC_9/Y VDD 2.38fF
C51056 NOR2X1_LOC_598/B INVX1_LOC_37/A 0.25fF
C51057 NOR2X1_LOC_423/Y INVX1_LOC_189/A 0.04fF
C51058 D_INPUT_1 NOR2X1_LOC_363/Y 0.10fF
C51059 INVX1_LOC_292/A INVX1_LOC_75/A 0.15fF
C51060 INVX1_LOC_233/A VDD 0.42fF
C51061 INVX1_LOC_41/A INVX1_LOC_16/A 0.03fF
C51062 NOR2X1_LOC_320/Y INVX1_LOC_161/Y 0.03fF
C51063 INVX1_LOC_174/A NAND2X1_LOC_2/a_36_24# 0.01fF
C51064 NOR2X1_LOC_226/A INVX1_LOC_168/A 0.25fF
C51065 INVX1_LOC_97/Y INVX1_LOC_37/A 0.09fF
C51066 NAND2X1_LOC_332/Y INVX1_LOC_22/A 0.03fF
C51067 NOR2X1_LOC_78/B INVX1_LOC_177/A 0.06fF
C51068 NOR2X1_LOC_457/A INVX1_LOC_69/Y 0.28fF
C51069 INVX1_LOC_35/A INVX1_LOC_12/Y 0.03fF
C51070 NOR2X1_LOC_803/A NOR2X1_LOC_148/A 0.07fF
C51071 INVX1_LOC_304/Y NAND2X1_LOC_862/A 0.01fF
C51072 INVX1_LOC_2/A NOR2X1_LOC_203/Y 0.03fF
C51073 INVX1_LOC_143/A NOR2X1_LOC_537/Y 0.07fF
C51074 NAND2X1_LOC_726/Y NAND2X1_LOC_357/B 0.01fF
C51075 NAND2X1_LOC_466/a_36_24# NOR2X1_LOC_435/A 0.00fF
C51076 NOR2X1_LOC_786/a_36_216# INVX1_LOC_286/A 0.00fF
C51077 NAND2X1_LOC_778/Y INVX1_LOC_20/A 0.01fF
C51078 NOR2X1_LOC_92/Y NAND2X1_LOC_626/a_36_24# 0.00fF
C51079 INVX1_LOC_34/A NOR2X1_LOC_521/Y 0.03fF
C51080 NOR2X1_LOC_590/A NOR2X1_LOC_188/A 0.19fF
C51081 NOR2X1_LOC_222/Y INVX1_LOC_189/A 0.18fF
C51082 NAND2X1_LOC_553/A VDD 0.34fF
C51083 INVX1_LOC_24/A INVX1_LOC_313/Y 0.07fF
C51084 INVX1_LOC_279/A INVX1_LOC_155/Y 0.01fF
C51085 NOR2X1_LOC_305/Y NOR2X1_LOC_406/A 0.01fF
C51086 NOR2X1_LOC_605/B NAND2X1_LOC_357/B 0.02fF
C51087 NOR2X1_LOC_590/A NOR2X1_LOC_548/B 0.03fF
C51088 NAND2X1_LOC_569/B NOR2X1_LOC_813/Y 0.16fF
C51089 NOR2X1_LOC_763/A NAND2X1_LOC_1/Y 0.12fF
C51090 NAND2X1_LOC_348/A INVX1_LOC_110/A 0.03fF
C51091 NOR2X1_LOC_510/Y INVX1_LOC_46/A 0.15fF
C51092 NOR2X1_LOC_798/A VDD 0.93fF
C51093 NOR2X1_LOC_191/B NAND2X1_LOC_842/B 0.04fF
C51094 INVX1_LOC_136/A NOR2X1_LOC_151/Y 0.03fF
C51095 INVX1_LOC_32/A INVX1_LOC_19/A 0.31fF
C51096 NOR2X1_LOC_742/A INVX1_LOC_18/A 0.14fF
C51097 NOR2X1_LOC_664/Y NOR2X1_LOC_719/B 0.08fF
C51098 INVX1_LOC_258/A INVX1_LOC_11/Y 0.01fF
C51099 NOR2X1_LOC_209/Y NOR2X1_LOC_687/Y 0.03fF
C51100 NOR2X1_LOC_716/B NAND2X1_LOC_862/Y 0.08fF
C51101 NAND2X1_LOC_565/B NAND2X1_LOC_338/B -0.05fF
C51102 NAND2X1_LOC_569/B INVX1_LOC_280/A 0.28fF
C51103 NAND2X1_LOC_361/Y INVX1_LOC_47/A 0.01fF
C51104 INVX1_LOC_69/Y INVX1_LOC_30/A 0.12fF
C51105 INVX1_LOC_290/Y NAND2X1_LOC_792/B 0.05fF
C51106 NAND2X1_LOC_703/Y VDD 0.00fF
C51107 NOR2X1_LOC_15/Y INVX1_LOC_20/A 7.54fF
C51108 INVX1_LOC_12/A D_INPUT_5 0.01fF
C51109 NOR2X1_LOC_722/Y INVX1_LOC_311/A 0.03fF
C51110 INVX1_LOC_82/Y D_INPUT_2 0.01fF
C51111 NAND2X1_LOC_663/a_36_24# NAND2X1_LOC_451/Y 0.00fF
C51112 INVX1_LOC_279/A NOR2X1_LOC_131/A -0.03fF
C51113 INVX1_LOC_14/A NOR2X1_LOC_558/A 0.36fF
C51114 NAND2X1_LOC_254/Y INVX1_LOC_3/Y 0.02fF
C51115 NAND2X1_LOC_853/Y NAND2X1_LOC_857/a_36_24# 0.08fF
C51116 NOR2X1_LOC_590/A NOR2X1_LOC_100/a_36_216# 0.00fF
C51117 NAND2X1_LOC_175/Y INVX1_LOC_19/A 0.07fF
C51118 NOR2X1_LOC_361/B INVX1_LOC_46/A 0.05fF
C51119 NOR2X1_LOC_647/A INVX1_LOC_63/A 0.04fF
C51120 NOR2X1_LOC_36/A NOR2X1_LOC_36/B 0.75fF
C51121 NAND2X1_LOC_552/A INVX1_LOC_54/A 0.01fF
C51122 INVX1_LOC_152/Y NOR2X1_LOC_61/A 0.45fF
C51123 NAND2X1_LOC_717/Y NOR2X1_LOC_299/Y 11.57fF
C51124 INVX1_LOC_5/A INVX1_LOC_54/A 0.13fF
C51125 INVX1_LOC_103/A NAND2X1_LOC_453/A 0.05fF
C51126 INVX1_LOC_57/A NOR2X1_LOC_430/Y 0.09fF
C51127 INVX1_LOC_13/Y INVX1_LOC_118/A 0.77fF
C51128 INVX1_LOC_241/A NAND2X1_LOC_735/B 0.01fF
C51129 NAND2X1_LOC_338/B NOR2X1_LOC_130/A 0.07fF
C51130 INVX1_LOC_163/A INVX1_LOC_166/Y 0.03fF
C51131 INVX1_LOC_182/Y INVX1_LOC_155/Y 1.15fF
C51132 INVX1_LOC_168/A INPUT_1 0.15fF
C51133 NAND2X1_LOC_784/A INVX1_LOC_285/A 0.00fF
C51134 NAND2X1_LOC_784/A INVX1_LOC_265/Y 0.01fF
C51135 NAND2X1_LOC_130/a_36_24# NOR2X1_LOC_131/Y 0.00fF
C51136 NOR2X1_LOC_25/Y INPUT_7 0.13fF
C51137 INVX1_LOC_28/A NAND2X1_LOC_477/A 0.08fF
C51138 NOR2X1_LOC_140/A INVX1_LOC_280/A 0.02fF
C51139 INVX1_LOC_178/A INVX1_LOC_54/A 0.11fF
C51140 NOR2X1_LOC_776/a_36_216# INVX1_LOC_37/A 0.00fF
C51141 NAND2X1_LOC_538/Y NOR2X1_LOC_152/A 0.06fF
C51142 INVX1_LOC_224/Y NAND2X1_LOC_773/B 0.07fF
C51143 NAND2X1_LOC_115/a_36_24# INVX1_LOC_79/A 0.00fF
C51144 NOR2X1_LOC_160/B NAND2X1_LOC_611/a_36_24# 0.00fF
C51145 NOR2X1_LOC_39/a_36_216# NAND2X1_LOC_74/B 0.00fF
C51146 INVX1_LOC_201/Y NAND2X1_LOC_126/a_36_24# -0.01fF
C51147 INVX1_LOC_93/Y INVX1_LOC_18/A 0.08fF
C51148 NOR2X1_LOC_414/Y NAND2X1_LOC_219/B 0.01fF
C51149 NOR2X1_LOC_372/A INVX1_LOC_37/A 0.32fF
C51150 INVX1_LOC_34/A INVX1_LOC_311/A 0.01fF
C51151 NAND2X1_LOC_357/B NOR2X1_LOC_323/Y 0.12fF
C51152 INVX1_LOC_253/A INVX1_LOC_15/A 0.01fF
C51153 NOR2X1_LOC_530/Y NOR2X1_LOC_813/Y 0.02fF
C51154 INVX1_LOC_16/Y INVX1_LOC_42/A 0.25fF
C51155 NAND2X1_LOC_425/Y NOR2X1_LOC_460/Y 0.03fF
C51156 NOR2X1_LOC_298/Y INPUT_5 0.03fF
C51157 NOR2X1_LOC_562/B NOR2X1_LOC_303/Y 0.08fF
C51158 INVX1_LOC_88/A INVX1_LOC_118/A 0.01fF
C51159 NOR2X1_LOC_332/A NOR2X1_LOC_195/a_36_216# 0.01fF
C51160 INVX1_LOC_31/A INVX1_LOC_33/Y 0.03fF
C51161 INVX1_LOC_250/A NOR2X1_LOC_305/Y 0.02fF
C51162 NAND2X1_LOC_833/Y NOR2X1_LOC_528/Y 0.03fF
C51163 NOR2X1_LOC_530/Y INVX1_LOC_280/A 0.10fF
C51164 NAND2X1_LOC_337/B NOR2X1_LOC_602/B 0.00fF
C51165 INVX1_LOC_78/A INVX1_LOC_21/Y 0.01fF
C51166 INVX1_LOC_77/A NAND2X1_LOC_642/Y 0.68fF
C51167 INVX1_LOC_18/A INVX1_LOC_139/A 0.00fF
C51168 INVX1_LOC_229/Y NOR2X1_LOC_576/B 2.62fF
C51169 INVX1_LOC_45/A NAND2X1_LOC_472/Y 0.07fF
C51170 INVX1_LOC_53/A NOR2X1_LOC_830/Y 0.02fF
C51171 NOR2X1_LOC_815/Y NAND2X1_LOC_655/A 0.11fF
C51172 NAND2X1_LOC_374/Y INVX1_LOC_91/Y 0.03fF
C51173 NAND2X1_LOC_205/A INVX1_LOC_42/A 0.03fF
C51174 NOR2X1_LOC_307/A NOR2X1_LOC_209/B 0.01fF
C51175 INVX1_LOC_235/A NAND2X1_LOC_659/A 0.03fF
C51176 INVX1_LOC_58/A NAND2X1_LOC_254/Y 0.10fF
C51177 NOR2X1_LOC_205/Y INVX1_LOC_92/A 0.03fF
C51178 INVX1_LOC_83/A NAND2X1_LOC_143/a_36_24# 0.01fF
C51179 NOR2X1_LOC_750/A NOR2X1_LOC_789/A 0.01fF
C51180 NAND2X1_LOC_787/A NOR2X1_LOC_89/A 0.03fF
C51181 NOR2X1_LOC_667/A INPUT_0 0.08fF
C51182 NAND2X1_LOC_323/B NOR2X1_LOC_112/B 0.19fF
C51183 INVX1_LOC_80/A INPUT_1 0.13fF
C51184 NOR2X1_LOC_816/A INVX1_LOC_54/A 0.04fF
C51185 NAND2X1_LOC_154/a_36_24# INVX1_LOC_117/Y 0.00fF
C51186 NOR2X1_LOC_382/Y NOR2X1_LOC_536/A 0.02fF
C51187 NAND2X1_LOC_363/B NOR2X1_LOC_89/A 0.03fF
C51188 NAND2X1_LOC_361/Y INVX1_LOC_95/Y 0.03fF
C51189 INVX1_LOC_166/A INVX1_LOC_32/A 0.61fF
C51190 NOR2X1_LOC_78/B INVX1_LOC_285/Y 0.00fF
C51191 NOR2X1_LOC_180/Y INVX1_LOC_91/A 0.03fF
C51192 NOR2X1_LOC_860/B NOR2X1_LOC_360/A 0.02fF
C51193 INVX1_LOC_301/Y VDD 0.41fF
C51194 NOR2X1_LOC_67/A INVX1_LOC_48/A 0.04fF
C51195 INVX1_LOC_144/A INVX1_LOC_53/Y 0.01fF
C51196 NAND2X1_LOC_866/A VDD 0.37fF
C51197 INVX1_LOC_13/Y NAND2X1_LOC_63/Y 0.03fF
C51198 NOR2X1_LOC_334/Y NOR2X1_LOC_106/a_36_216# 0.00fF
C51199 NOR2X1_LOC_172/a_36_216# INVX1_LOC_91/A 0.01fF
C51200 INVX1_LOC_41/A NOR2X1_LOC_35/Y 0.05fF
C51201 NOR2X1_LOC_791/B NOR2X1_LOC_99/a_36_216# 0.00fF
C51202 INVX1_LOC_34/A NOR2X1_LOC_670/Y 0.01fF
C51203 INVX1_LOC_35/A NOR2X1_LOC_554/A 0.04fF
C51204 INVX1_LOC_124/A NAND2X1_LOC_642/Y 0.28fF
C51205 INVX1_LOC_71/A NAND2X1_LOC_472/Y 0.07fF
C51206 NOR2X1_LOC_387/A NAND2X1_LOC_863/B 0.12fF
C51207 NAND2X1_LOC_812/A VDD -0.00fF
C51208 INVX1_LOC_172/A NAND2X1_LOC_721/A 0.16fF
C51209 NAND2X1_LOC_374/Y NOR2X1_LOC_45/B 0.09fF
C51210 INVX1_LOC_314/Y INVX1_LOC_117/A 0.00fF
C51211 NAND2X1_LOC_465/Y NAND2X1_LOC_465/A 0.00fF
C51212 INVX1_LOC_57/A INVX1_LOC_94/Y 0.07fF
C51213 NOR2X1_LOC_454/Y NOR2X1_LOC_48/Y 0.04fF
C51214 NOR2X1_LOC_858/A INVX1_LOC_271/Y 0.02fF
C51215 NOR2X1_LOC_91/A INVX1_LOC_23/Y 0.07fF
C51216 INVX1_LOC_5/A NOR2X1_LOC_48/B 0.06fF
C51217 NOR2X1_LOC_334/Y NOR2X1_LOC_493/A 0.03fF
C51218 NOR2X1_LOC_84/a_36_216# INVX1_LOC_59/Y 0.00fF
C51219 INVX1_LOC_93/Y NOR2X1_LOC_709/a_36_216# 0.01fF
C51220 NAND2X1_LOC_807/A INVX1_LOC_285/A 0.04fF
C51221 NOR2X1_LOC_78/A NOR2X1_LOC_131/a_36_216# 0.00fF
C51222 NOR2X1_LOC_78/B INVX1_LOC_65/A 0.00fF
C51223 INVX1_LOC_227/A NOR2X1_LOC_188/A 0.37fF
C51224 INVX1_LOC_53/A INVX1_LOC_4/Y 0.02fF
C51225 NOR2X1_LOC_723/Y INVX1_LOC_92/A 0.08fF
C51226 INVX1_LOC_36/A NAND2X1_LOC_798/B 0.07fF
C51227 NOR2X1_LOC_273/a_36_216# INVX1_LOC_54/A 0.00fF
C51228 NOR2X1_LOC_92/Y INVX1_LOC_109/A 0.04fF
C51229 NOR2X1_LOC_352/Y INVX1_LOC_247/A 0.01fF
C51230 NAND2X1_LOC_633/Y NOR2X1_LOC_278/A 0.16fF
C51231 NOR2X1_LOC_773/Y INVX1_LOC_95/A 0.03fF
C51232 NOR2X1_LOC_216/Y INVX1_LOC_313/Y 0.02fF
C51233 NOR2X1_LOC_598/B NAND2X1_LOC_72/B 0.01fF
C51234 NOR2X1_LOC_103/Y NAND2X1_LOC_773/B 0.15fF
C51235 INVX1_LOC_178/A NOR2X1_LOC_48/B 0.19fF
C51236 INVX1_LOC_18/A INVX1_LOC_117/Y 0.20fF
C51237 INVX1_LOC_243/Y INVX1_LOC_296/A 0.22fF
C51238 NAND2X1_LOC_731/Y INVX1_LOC_185/A 0.00fF
C51239 INVX1_LOC_23/A INVX1_LOC_23/Y 0.03fF
C51240 INVX1_LOC_26/Y NOR2X1_LOC_622/A 0.01fF
C51241 INVX1_LOC_177/A INVX1_LOC_46/A 0.03fF
C51242 NOR2X1_LOC_360/Y INVX1_LOC_307/A 0.03fF
C51243 NOR2X1_LOC_160/B NOR2X1_LOC_691/B 0.07fF
C51244 INVX1_LOC_2/Y NOR2X1_LOC_87/a_36_216# 0.00fF
C51245 INVX1_LOC_64/A INVX1_LOC_273/A 0.00fF
C51246 INVX1_LOC_286/Y INVX1_LOC_119/Y 0.00fF
C51247 INVX1_LOC_132/A INVX1_LOC_9/A 0.12fF
C51248 NOR2X1_LOC_156/B INVX1_LOC_37/A 0.01fF
C51249 INVX1_LOC_57/A INVX1_LOC_296/A 0.03fF
C51250 NOR2X1_LOC_272/Y INVX1_LOC_15/A 0.17fF
C51251 INVX1_LOC_134/A NOR2X1_LOC_777/B 0.03fF
C51252 NOR2X1_LOC_382/Y NOR2X1_LOC_649/B 0.01fF
C51253 NAND2X1_LOC_541/Y INVX1_LOC_76/A 0.01fF
C51254 NOR2X1_LOC_561/Y NOR2X1_LOC_78/A 0.01fF
C51255 INVX1_LOC_7/A NOR2X1_LOC_78/A 4.91fF
C51256 NAND2X1_LOC_840/B INVX1_LOC_20/A 0.00fF
C51257 INVX1_LOC_10/A NOR2X1_LOC_269/Y 0.07fF
C51258 NOR2X1_LOC_222/Y NAND2X1_LOC_211/Y 0.12fF
C51259 INVX1_LOC_280/Y INVX1_LOC_46/A 0.15fF
C51260 VDD NOR2X1_LOC_505/Y 0.33fF
C51261 NOR2X1_LOC_817/Y NOR2X1_LOC_847/A 0.21fF
C51262 NOR2X1_LOC_300/a_36_216# INVX1_LOC_22/A 0.00fF
C51263 INVX1_LOC_177/A NAND2X1_LOC_417/a_36_24# 0.02fF
C51264 NOR2X1_LOC_211/A NOR2X1_LOC_35/Y 0.12fF
C51265 D_INPUT_1 INVX1_LOC_29/Y 0.00fF
C51266 NAND2X1_LOC_337/B NAND2X1_LOC_807/B 0.00fF
C51267 NAND2X1_LOC_364/A INVX1_LOC_84/A 0.03fF
C51268 INVX1_LOC_45/A NAND2X1_LOC_773/B 0.46fF
C51269 NOR2X1_LOC_790/B NOR2X1_LOC_748/A 0.33fF
C51270 NOR2X1_LOC_778/B INVX1_LOC_117/A 0.03fF
C51271 NAND2X1_LOC_112/Y INVX1_LOC_76/A 0.08fF
C51272 INVX1_LOC_205/A INVX1_LOC_63/A 0.03fF
C51273 NAND2X1_LOC_555/Y NOR2X1_LOC_33/B 0.04fF
C51274 NOR2X1_LOC_318/B NAND2X1_LOC_105/a_36_24# 0.00fF
C51275 NOR2X1_LOC_15/Y INVX1_LOC_4/A 0.14fF
C51276 INVX1_LOC_234/A NOR2X1_LOC_24/a_36_216# 0.00fF
C51277 NOR2X1_LOC_816/A NOR2X1_LOC_48/B 0.11fF
C51278 NAND2X1_LOC_787/A NAND2X1_LOC_804/A 0.00fF
C51279 NOR2X1_LOC_500/B NAND2X1_LOC_63/Y 1.34fF
C51280 NOR2X1_LOC_209/Y INVX1_LOC_9/A 0.07fF
C51281 NAND2X1_LOC_474/Y INVX1_LOC_26/A 0.78fF
C51282 INVX1_LOC_161/Y INVX1_LOC_32/A 0.01fF
C51283 INVX1_LOC_5/A NAND2X1_LOC_215/A 0.00fF
C51284 INVX1_LOC_30/A NOR2X1_LOC_89/A 0.40fF
C51285 NAND2X1_LOC_573/A INVX1_LOC_46/A 0.21fF
C51286 NOR2X1_LOC_576/B INVX1_LOC_20/A 0.02fF
C51287 NOR2X1_LOC_700/Y VDD 0.12fF
C51288 INVX1_LOC_71/A NAND2X1_LOC_773/B 0.02fF
C51289 NOR2X1_LOC_652/Y INVX1_LOC_29/Y 0.20fF
C51290 NOR2X1_LOC_773/Y INVX1_LOC_54/A 0.07fF
C51291 NOR2X1_LOC_321/Y NOR2X1_LOC_65/Y 0.01fF
C51292 NAND2X1_LOC_785/A NOR2X1_LOC_88/Y 0.07fF
C51293 NAND2X1_LOC_451/Y NAND2X1_LOC_428/a_36_24# 0.00fF
C51294 INVX1_LOC_161/Y NAND2X1_LOC_175/Y 0.02fF
C51295 NOR2X1_LOC_537/Y NOR2X1_LOC_197/B 0.46fF
C51296 INVX1_LOC_303/A NAND2X1_LOC_63/Y 0.04fF
C51297 INVX1_LOC_36/A INVX1_LOC_47/Y 0.11fF
C51298 INVX1_LOC_49/A INVX1_LOC_272/A 0.07fF
C51299 NOR2X1_LOC_500/a_36_216# INVX1_LOC_91/A 0.03fF
C51300 NOR2X1_LOC_272/Y INVX1_LOC_278/A 0.10fF
C51301 NOR2X1_LOC_793/Y NOR2X1_LOC_383/B 0.14fF
C51302 NAND2X1_LOC_842/B VDD 0.31fF
C51303 NOR2X1_LOC_359/Y INVX1_LOC_290/Y 0.01fF
C51304 INVX1_LOC_299/A INVX1_LOC_57/A 0.03fF
C51305 NOR2X1_LOC_790/A INVX1_LOC_53/A 0.02fF
C51306 NOR2X1_LOC_329/B NAND2X1_LOC_211/Y 0.02fF
C51307 INPUT_0 INVX1_LOC_304/A 0.07fF
C51308 INVX1_LOC_146/A INVX1_LOC_146/Y 0.12fF
C51309 INVX1_LOC_30/A INVX1_LOC_104/Y 0.02fF
C51310 NOR2X1_LOC_87/B NOR2X1_LOC_814/A 0.02fF
C51311 NAND2X1_LOC_785/A INVX1_LOC_84/A 0.03fF
C51312 NOR2X1_LOC_690/A NAND2X1_LOC_500/B 0.01fF
C51313 NAND2X1_LOC_364/A INVX1_LOC_15/A 0.07fF
C51314 INVX1_LOC_133/Y NOR2X1_LOC_127/Y 0.01fF
C51315 INVX1_LOC_146/A VDD 0.24fF
C51316 NOR2X1_LOC_638/a_36_216# NOR2X1_LOC_584/Y -0.00fF
C51317 NOR2X1_LOC_315/Y NOR2X1_LOC_662/A 0.01fF
C51318 NOR2X1_LOC_724/Y INVX1_LOC_117/A 0.03fF
C51319 NAND2X1_LOC_652/a_36_24# INVX1_LOC_12/A 0.00fF
C51320 NOR2X1_LOC_288/A NOR2X1_LOC_691/a_36_216# 0.00fF
C51321 INVX1_LOC_53/Y NOR2X1_LOC_155/A 0.04fF
C51322 INVX1_LOC_207/A INVX1_LOC_12/A 0.03fF
C51323 NOR2X1_LOC_655/B INVX1_LOC_27/Y 0.42fF
C51324 D_GATE_741 INVX1_LOC_275/Y 0.03fF
C51325 INVX1_LOC_50/Y NOR2X1_LOC_849/A 0.59fF
C51326 INVX1_LOC_75/A NOR2X1_LOC_137/Y 0.03fF
C51327 INVX1_LOC_312/A NAND2X1_LOC_175/Y 0.03fF
C51328 INVX1_LOC_31/A INVX1_LOC_23/Y 0.08fF
C51329 NOR2X1_LOC_632/Y INVX1_LOC_179/A 0.01fF
C51330 NAND2X1_LOC_11/Y INVX1_LOC_84/A 0.00fF
C51331 NAND2X1_LOC_807/Y INVX1_LOC_33/Y 0.04fF
C51332 NAND2X1_LOC_9/Y NOR2X1_LOC_361/B 0.03fF
C51333 INVX1_LOC_35/A NOR2X1_LOC_793/A 0.02fF
C51334 INVX1_LOC_39/A INVX1_LOC_13/Y 0.01fF
C51335 NOR2X1_LOC_205/Y INVX1_LOC_53/A 0.02fF
C51336 INVX1_LOC_45/Y NOR2X1_LOC_609/Y 0.00fF
C51337 NOR2X1_LOC_665/A NOR2X1_LOC_155/A 0.03fF
C51338 INVX1_LOC_64/A NOR2X1_LOC_15/Y 0.17fF
C51339 NOR2X1_LOC_86/A NOR2X1_LOC_88/Y 0.01fF
C51340 INVX1_LOC_233/A NOR2X1_LOC_361/B 0.10fF
C51341 INVX1_LOC_31/A NOR2X1_LOC_686/a_36_216# 0.00fF
C51342 NOR2X1_LOC_312/Y INVX1_LOC_185/A 0.01fF
C51343 INVX1_LOC_224/A NAND2X1_LOC_363/B 0.08fF
C51344 INVX1_LOC_11/A NAND2X1_LOC_363/B 0.07fF
C51345 NOR2X1_LOC_91/A NAND2X1_LOC_741/B 0.04fF
C51346 INVX1_LOC_2/A INVX1_LOC_272/A 0.36fF
C51347 INVX1_LOC_285/Y INVX1_LOC_46/A 0.01fF
C51348 NOR2X1_LOC_238/a_36_216# INVX1_LOC_78/A 0.00fF
C51349 INVX1_LOC_16/A INVX1_LOC_136/Y 0.01fF
C51350 NOR2X1_LOC_152/Y INVX1_LOC_21/Y 0.05fF
C51351 NAND2X1_LOC_784/A NOR2X1_LOC_590/A 0.00fF
C51352 INVX1_LOC_150/A NOR2X1_LOC_831/B 0.03fF
C51353 NOR2X1_LOC_226/A INVX1_LOC_272/A 0.01fF
C51354 NAND2X1_LOC_722/A NOR2X1_LOC_89/A 0.08fF
C51355 NOR2X1_LOC_86/A INVX1_LOC_84/A 0.07fF
C51356 INPUT_1 NOR2X1_LOC_99/Y 0.15fF
C51357 INVX1_LOC_35/A NOR2X1_LOC_160/B 0.91fF
C51358 NOR2X1_LOC_78/B NOR2X1_LOC_830/Y 0.01fF
C51359 NOR2X1_LOC_78/A INVX1_LOC_76/A 0.09fF
C51360 NOR2X1_LOC_272/a_36_216# INVX1_LOC_88/A 0.00fF
C51361 INVX1_LOC_89/A NOR2X1_LOC_831/B 0.01fF
C51362 INVX1_LOC_140/A INVX1_LOC_54/A 1.36fF
C51363 NOR2X1_LOC_309/Y INVX1_LOC_47/Y 0.02fF
C51364 NAND2X1_LOC_564/B INVX1_LOC_19/A 0.07fF
C51365 INVX1_LOC_313/Y NOR2X1_LOC_197/B 0.10fF
C51366 NOR2X1_LOC_218/Y INVX1_LOC_272/A 0.03fF
C51367 INVX1_LOC_11/A NOR2X1_LOC_791/Y 0.04fF
C51368 NOR2X1_LOC_388/Y NOR2X1_LOC_334/Y 0.03fF
C51369 NOR2X1_LOC_237/Y NOR2X1_LOC_693/a_36_216# 0.01fF
C51370 NOR2X1_LOC_476/Y NOR2X1_LOC_476/B 0.02fF
C51371 INVX1_LOC_71/A NOR2X1_LOC_481/a_36_216# 0.00fF
C51372 NOR2X1_LOC_570/B INVX1_LOC_78/A 0.02fF
C51373 NOR2X1_LOC_557/A INVX1_LOC_117/A 0.07fF
C51374 NOR2X1_LOC_773/Y NOR2X1_LOC_48/B 0.09fF
C51375 NOR2X1_LOC_816/a_36_216# INVX1_LOC_215/Y 0.01fF
C51376 INVX1_LOC_50/A NOR2X1_LOC_238/Y 0.00fF
C51377 NAND2X1_LOC_181/Y INVX1_LOC_170/Y 0.03fF
C51378 INVX1_LOC_224/Y INVX1_LOC_24/A 1.56fF
C51379 INVX1_LOC_21/A INVX1_LOC_225/Y 0.01fF
C51380 VDD NOR2X1_LOC_545/B -0.00fF
C51381 NOR2X1_LOC_76/A NAND2X1_LOC_477/Y 0.38fF
C51382 INVX1_LOC_96/Y INVX1_LOC_4/A 0.49fF
C51383 NAND2X1_LOC_350/A INVX1_LOC_178/A 0.10fF
C51384 INVX1_LOC_35/A NAND2X1_LOC_195/Y 0.02fF
C51385 NOR2X1_LOC_567/B NOR2X1_LOC_445/B 0.07fF
C51386 NAND2X1_LOC_11/Y INVX1_LOC_15/A 0.25fF
C51387 NOR2X1_LOC_391/A NAND2X1_LOC_74/B 0.01fF
C51388 INVX1_LOC_14/Y NOR2X1_LOC_683/Y 0.02fF
C51389 NAND2X1_LOC_803/B NAND2X1_LOC_326/A 0.02fF
C51390 INVX1_LOC_31/A NOR2X1_LOC_846/A 0.01fF
C51391 INVX1_LOC_289/Y NAND2X1_LOC_799/A 4.05fF
C51392 INVX1_LOC_58/A INVX1_LOC_314/Y 0.01fF
C51393 NAND2X1_LOC_569/A NAND2X1_LOC_99/A 0.02fF
C51394 INVX1_LOC_24/A NAND2X1_LOC_793/B 0.07fF
C51395 NOR2X1_LOC_92/Y INVX1_LOC_246/A 0.01fF
C51396 NAND2X1_LOC_267/B INVX1_LOC_46/A 0.03fF
C51397 NOR2X1_LOC_78/B INVX1_LOC_4/Y 0.10fF
C51398 NOR2X1_LOC_590/A NAND2X1_LOC_326/A 0.07fF
C51399 INVX1_LOC_75/A NAND2X1_LOC_659/A 0.40fF
C51400 NAND2X1_LOC_642/Y INVX1_LOC_9/A 0.03fF
C51401 NOR2X1_LOC_201/A NAND2X1_LOC_116/A 0.00fF
C51402 INVX1_LOC_103/A NOR2X1_LOC_592/a_36_216# 0.00fF
C51403 NAND2X1_LOC_715/B NAND2X1_LOC_198/B 0.11fF
C51404 INVX1_LOC_64/A NOR2X1_LOC_860/B 0.01fF
C51405 INVX1_LOC_162/A INVX1_LOC_57/A 0.11fF
C51406 NOR2X1_LOC_290/Y INVX1_LOC_23/Y 0.01fF
C51407 INVX1_LOC_120/A NAND2X1_LOC_291/B 0.12fF
C51408 INVX1_LOC_76/A NOR2X1_LOC_60/Y 0.03fF
C51409 NOR2X1_LOC_86/A INVX1_LOC_15/A 0.03fF
C51410 NAND2X1_LOC_578/a_36_24# NAND2X1_LOC_577/A 0.01fF
C51411 NOR2X1_LOC_527/Y INVX1_LOC_285/A 0.01fF
C51412 NOR2X1_LOC_100/A NOR2X1_LOC_843/B 0.03fF
C51413 NOR2X1_LOC_527/Y INVX1_LOC_265/Y 0.06fF
C51414 NOR2X1_LOC_598/B INVX1_LOC_310/Y 0.10fF
C51415 NOR2X1_LOC_315/Y INVX1_LOC_57/A 0.07fF
C51416 NOR2X1_LOC_843/A INVX1_LOC_53/A 0.07fF
C51417 NOR2X1_LOC_160/B NOR2X1_LOC_502/Y 0.17fF
C51418 D_INPUT_1 INVX1_LOC_60/Y 0.09fF
C51419 NOR2X1_LOC_19/B NOR2X1_LOC_14/a_36_216# 0.00fF
C51420 INVX1_LOC_33/A INVX1_LOC_213/A 0.13fF
C51421 INVX1_LOC_224/A INVX1_LOC_30/A 0.00fF
C51422 INVX1_LOC_215/A INVX1_LOC_78/A 0.04fF
C51423 INVX1_LOC_226/Y INVX1_LOC_26/A 0.16fF
C51424 NAND2X1_LOC_787/A NOR2X1_LOC_52/B 0.04fF
C51425 INVX1_LOC_11/A INVX1_LOC_30/A 1.10fF
C51426 NAND2X1_LOC_722/A NAND2X1_LOC_804/A 0.01fF
C51427 NOR2X1_LOC_667/Y INVX1_LOC_236/Y 0.01fF
C51428 INVX1_LOC_5/A NOR2X1_LOC_142/Y 0.01fF
C51429 NOR2X1_LOC_83/a_36_216# NAND2X1_LOC_63/Y 0.00fF
C51430 INVX1_LOC_278/A NAND2X1_LOC_785/A 0.07fF
C51431 NAND2X1_LOC_763/B INVX1_LOC_11/A 1.73fF
C51432 NAND2X1_LOC_472/Y NOR2X1_LOC_331/B 0.09fF
C51433 INVX1_LOC_93/A NAND2X1_LOC_833/Y 0.02fF
C51434 INVX1_LOC_135/A NOR2X1_LOC_334/Y 0.02fF
C51435 NOR2X1_LOC_620/Y INVX1_LOC_27/A 0.28fF
C51436 INVX1_LOC_14/A INVX1_LOC_181/Y 0.02fF
C51437 INVX1_LOC_140/A NOR2X1_LOC_48/B 0.19fF
C51438 NOR2X1_LOC_817/Y NOR2X1_LOC_554/B 0.60fF
C51439 NOR2X1_LOC_859/a_36_216# NOR2X1_LOC_68/A 0.00fF
C51440 INVX1_LOC_58/A NAND2X1_LOC_532/a_36_24# 0.01fF
C51441 NOR2X1_LOC_373/Y INVX1_LOC_78/A 0.53fF
C51442 INVX1_LOC_64/A INVX1_LOC_96/Y 0.09fF
C51443 INVX1_LOC_64/A INVX1_LOC_15/Y 0.06fF
C51444 NOR2X1_LOC_65/B INVX1_LOC_215/A 0.18fF
C51445 NAND2X1_LOC_9/Y NOR2X1_LOC_547/a_36_216# 0.00fF
C51446 INVX1_LOC_10/A INVX1_LOC_26/A 0.12fF
C51447 NOR2X1_LOC_405/A INVX1_LOC_84/A 0.05fF
C51448 NOR2X1_LOC_427/Y INVX1_LOC_12/A 0.07fF
C51449 NOR2X1_LOC_188/A NOR2X1_LOC_67/Y 0.15fF
C51450 INVX1_LOC_24/Y NOR2X1_LOC_350/A 0.02fF
C51451 NOR2X1_LOC_754/a_36_216# INVX1_LOC_42/A 0.00fF
C51452 INVX1_LOC_24/A NOR2X1_LOC_103/Y 0.16fF
C51453 VDD NAND2X1_LOC_243/B 0.01fF
C51454 INVX1_LOC_35/A NAND2X1_LOC_350/B 0.39fF
C51455 NAND2X1_LOC_35/Y NAND2X1_LOC_717/Y 0.07fF
C51456 INVX1_LOC_37/A NOR2X1_LOC_634/A 0.18fF
C51457 INVX1_LOC_230/Y NOR2X1_LOC_68/A 0.22fF
C51458 NAND2X1_LOC_574/A NOR2X1_LOC_35/Y 0.04fF
C51459 INVX1_LOC_30/Y INVX1_LOC_129/A 0.00fF
C51460 INVX1_LOC_286/Y INVX1_LOC_72/A 0.10fF
C51461 INVX1_LOC_64/A INVX1_LOC_226/A 0.03fF
C51462 NAND2X1_LOC_373/a_36_24# NOR2X1_LOC_317/B 0.00fF
C51463 NOR2X1_LOC_655/B INVX1_LOC_5/A 0.04fF
C51464 INVX1_LOC_251/Y NOR2X1_LOC_81/Y 0.02fF
C51465 D_INPUT_3 NAND2X1_LOC_141/Y 0.06fF
C51466 NOR2X1_LOC_163/a_36_216# NAND2X1_LOC_452/Y 0.00fF
C51467 INVX1_LOC_103/A NOR2X1_LOC_577/Y 0.08fF
C51468 NOR2X1_LOC_690/A NAND2X1_LOC_725/B 0.07fF
C51469 INVX1_LOC_90/A NOR2X1_LOC_25/Y 0.03fF
C51470 NOR2X1_LOC_815/Y INVX1_LOC_88/A 0.01fF
C51471 INVX1_LOC_279/A NOR2X1_LOC_858/A 0.01fF
C51472 INVX1_LOC_226/Y NOR2X1_LOC_619/a_36_216# 0.00fF
C51473 INVX1_LOC_59/A INVX1_LOC_219/Y 0.01fF
C51474 NOR2X1_LOC_279/Y NOR2X1_LOC_653/Y 0.08fF
C51475 INVX1_LOC_286/A INVX1_LOC_42/A 0.07fF
C51476 INVX1_LOC_35/A NOR2X1_LOC_516/B 0.13fF
C51477 NAND2X1_LOC_36/A INVX1_LOC_18/A 0.12fF
C51478 NOR2X1_LOC_15/Y NOR2X1_LOC_459/B 0.00fF
C51479 INVX1_LOC_75/A NOR2X1_LOC_227/A 0.03fF
C51480 VDD INVX1_LOC_119/Y 0.67fF
C51481 INVX1_LOC_49/A INVX1_LOC_150/Y 0.23fF
C51482 INVX1_LOC_230/Y NOR2X1_LOC_204/a_36_216# 0.01fF
C51483 NAND2X1_LOC_12/a_36_24# NAND2X1_LOC_36/A 0.01fF
C51484 INVX1_LOC_14/Y NOR2X1_LOC_66/Y 0.03fF
C51485 INVX1_LOC_1/A INVX1_LOC_104/A 0.03fF
C51486 NOR2X1_LOC_366/Y INVX1_LOC_23/A 0.00fF
C51487 NAND2X1_LOC_35/Y INVX1_LOC_16/A 0.11fF
C51488 NAND2X1_LOC_563/Y INVX1_LOC_14/A 0.02fF
C51489 D_INPUT_1 NOR2X1_LOC_355/A 0.07fF
C51490 INVX1_LOC_33/A NOR2X1_LOC_745/Y 0.03fF
C51491 INVX1_LOC_292/A NOR2X1_LOC_577/Y 0.25fF
C51492 INVX1_LOC_50/A INVX1_LOC_47/A 0.03fF
C51493 INVX1_LOC_45/A INVX1_LOC_24/A 0.45fF
C51494 INVX1_LOC_27/A NAND2X1_LOC_181/Y 0.04fF
C51495 INVX1_LOC_233/A NAND2X1_LOC_573/A 0.02fF
C51496 INVX1_LOC_49/Y INVX1_LOC_20/A 0.06fF
C51497 INVX1_LOC_24/A NOR2X1_LOC_568/A 0.09fF
C51498 INVX1_LOC_140/A NOR2X1_LOC_438/Y 0.12fF
C51499 NOR2X1_LOC_233/a_36_216# INVX1_LOC_25/Y 0.01fF
C51500 NOR2X1_LOC_224/a_36_216# NOR2X1_LOC_696/Y 0.00fF
C51501 INVX1_LOC_299/A NAND2X1_LOC_164/a_36_24# 0.00fF
C51502 NOR2X1_LOC_790/B INVX1_LOC_89/A 0.03fF
C51503 NOR2X1_LOC_433/A INVX1_LOC_30/A 0.16fF
C51504 NOR2X1_LOC_15/Y NAND2X1_LOC_850/Y 0.48fF
C51505 NOR2X1_LOC_590/A NOR2X1_LOC_285/B 0.01fF
C51506 NOR2X1_LOC_74/A NOR2X1_LOC_301/A 0.07fF
C51507 NOR2X1_LOC_454/Y NOR2X1_LOC_229/a_36_216# 0.01fF
C51508 NOR2X1_LOC_349/A INVX1_LOC_15/A 0.05fF
C51509 NOR2X1_LOC_794/B INVX1_LOC_104/A 0.02fF
C51510 INVX1_LOC_11/A NAND2X1_LOC_722/A 0.57fF
C51511 NOR2X1_LOC_78/B NOR2X1_LOC_205/Y 0.10fF
C51512 NOR2X1_LOC_186/Y NOR2X1_LOC_561/Y 0.03fF
C51513 INVX1_LOC_286/A INVX1_LOC_78/A 0.10fF
C51514 NAND2X1_LOC_434/Y NOR2X1_LOC_592/B 0.01fF
C51515 NOR2X1_LOC_156/Y INVX1_LOC_92/A 0.02fF
C51516 INVX1_LOC_37/A INVX1_LOC_29/A 2.93fF
C51517 NOR2X1_LOC_636/B INVX1_LOC_191/Y 0.04fF
C51518 NAND2X1_LOC_802/A NAND2X1_LOC_354/Y 0.22fF
C51519 NAND2X1_LOC_798/B NOR2X1_LOC_435/A 0.17fF
C51520 NOR2X1_LOC_82/A INVX1_LOC_34/Y 0.46fF
C51521 NOR2X1_LOC_593/Y INVX1_LOC_30/A 0.39fF
C51522 INVX1_LOC_5/A NOR2X1_LOC_99/B 0.14fF
C51523 VDD NOR2X1_LOC_755/Y -0.00fF
C51524 NAND2X1_LOC_348/A NOR2X1_LOC_646/B 0.00fF
C51525 INVX1_LOC_30/Y NOR2X1_LOC_440/B 0.01fF
C51526 NAND2X1_LOC_116/A INVX1_LOC_31/A 0.06fF
C51527 VDD INVX1_LOC_284/A 1.01fF
C51528 NAND2X1_LOC_711/Y NAND2X1_LOC_357/B 0.01fF
C51529 INVX1_LOC_72/A NAND2X1_LOC_486/a_36_24# 0.01fF
C51530 NOR2X1_LOC_514/A NOR2X1_LOC_6/B 0.48fF
C51531 INVX1_LOC_24/A INVX1_LOC_71/A 0.03fF
C51532 INVX1_LOC_6/A INVX1_LOC_23/Y 0.00fF
C51533 INVX1_LOC_151/A INVX1_LOC_30/A 0.01fF
C51534 INVX1_LOC_5/A NOR2X1_LOC_846/B 0.02fF
C51535 INVX1_LOC_99/Y NOR2X1_LOC_180/B 0.01fF
C51536 INVX1_LOC_103/A INVX1_LOC_22/A 0.19fF
C51537 NOR2X1_LOC_52/B INVX1_LOC_30/A 0.13fF
C51538 NOR2X1_LOC_65/B INVX1_LOC_286/A 0.07fF
C51539 NAND2X1_LOC_35/Y INVX1_LOC_28/A 0.03fF
C51540 INVX1_LOC_31/A NOR2X1_LOC_511/a_36_216# 0.02fF
C51541 NAND2X1_LOC_220/a_36_24# NOR2X1_LOC_467/A 0.01fF
C51542 NOR2X1_LOC_551/Y NOR2X1_LOC_383/B 0.01fF
C51543 NOR2X1_LOC_666/A INVX1_LOC_10/A 0.17fF
C51544 NOR2X1_LOC_857/A INVX1_LOC_15/A 0.07fF
C51545 NOR2X1_LOC_789/B INVX1_LOC_89/A 0.02fF
C51546 INVX1_LOC_35/A NOR2X1_LOC_706/A 0.00fF
C51547 INVX1_LOC_9/Y INVX1_LOC_161/Y 0.01fF
C51548 NOR2X1_LOC_673/A INVX1_LOC_46/Y 0.00fF
C51549 NAND2X1_LOC_303/Y NOR2X1_LOC_298/Y 0.30fF
C51550 NOR2X1_LOC_149/a_36_216# INVX1_LOC_301/A 0.00fF
C51551 INVX1_LOC_272/A INVX1_LOC_118/A 0.10fF
C51552 INVX1_LOC_5/A INVX1_LOC_182/A 0.09fF
C51553 NOR2X1_LOC_557/Y INVX1_LOC_71/A 0.10fF
C51554 NOR2X1_LOC_441/Y NOR2X1_LOC_773/Y 0.07fF
C51555 INVX1_LOC_305/A NOR2X1_LOC_802/A 0.17fF
C51556 INVX1_LOC_45/A INVX1_LOC_143/A 0.05fF
C51557 NOR2X1_LOC_720/B INVX1_LOC_62/Y 0.01fF
C51558 NAND2X1_LOC_798/B INVX1_LOC_63/A 0.18fF
C51559 NOR2X1_LOC_91/Y NAND2X1_LOC_650/a_36_24# 0.00fF
C51560 INVX1_LOC_292/A INVX1_LOC_22/A 0.07fF
C51561 INVX1_LOC_41/A NOR2X1_LOC_350/A 0.99fF
C51562 NAND2X1_LOC_35/B INVX1_LOC_72/A 0.07fF
C51563 NAND2X1_LOC_217/a_36_24# INVX1_LOC_201/Y 0.02fF
C51564 INVX1_LOC_67/A NOR2X1_LOC_577/Y 0.03fF
C51565 NOR2X1_LOC_78/B NOR2X1_LOC_723/Y 0.01fF
C51566 NOR2X1_LOC_82/A NOR2X1_LOC_383/a_36_216# 0.00fF
C51567 INVX1_LOC_46/A INVX1_LOC_4/Y 0.21fF
C51568 INVX1_LOC_31/A INVX1_LOC_232/A 0.07fF
C51569 INVX1_LOC_207/A NAND2X1_LOC_787/B 0.05fF
C51570 NOR2X1_LOC_624/A INVX1_LOC_303/A 0.03fF
C51571 NOR2X1_LOC_685/A INVX1_LOC_23/A 0.33fF
C51572 NAND2X1_LOC_577/A INVX1_LOC_316/Y 0.03fF
C51573 INVX1_LOC_181/Y NOR2X1_LOC_612/B 0.01fF
C51574 INVX1_LOC_186/A INVX1_LOC_23/A 0.03fF
C51575 NOR2X1_LOC_743/Y INVX1_LOC_29/A 0.03fF
C51576 INVX1_LOC_118/A NOR2X1_LOC_76/B 0.06fF
C51577 NOR2X1_LOC_103/Y NOR2X1_LOC_130/A 0.03fF
C51578 NOR2X1_LOC_45/Y NOR2X1_LOC_561/Y 0.07fF
C51579 NAND2X1_LOC_340/a_36_24# NAND2X1_LOC_319/A 0.00fF
C51580 INVX1_LOC_276/A NOR2X1_LOC_512/Y 0.00fF
C51581 INVX1_LOC_54/A INVX1_LOC_42/A 0.09fF
C51582 INVX1_LOC_117/A NOR2X1_LOC_839/B 0.01fF
C51583 NOR2X1_LOC_328/Y INVX1_LOC_36/A 1.52fF
C51584 NOR2X1_LOC_577/Y INVX1_LOC_240/A 0.10fF
C51585 NOR2X1_LOC_360/Y NOR2X1_LOC_566/Y 0.03fF
C51586 NOR2X1_LOC_361/B NAND2X1_LOC_842/B 1.33fF
C51587 INVX1_LOC_89/A D_GATE_741 0.05fF
C51588 INVX1_LOC_123/A INVX1_LOC_138/Y 0.09fF
C51589 INVX1_LOC_298/Y INVX1_LOC_37/A 0.01fF
C51590 INVX1_LOC_176/A NOR2X1_LOC_843/B 0.03fF
C51591 INVX1_LOC_143/A INVX1_LOC_71/A 0.10fF
C51592 INVX1_LOC_17/A NOR2X1_LOC_356/A 0.08fF
C51593 NAND2X1_LOC_559/Y NAND2X1_LOC_560/A 0.11fF
C51594 NOR2X1_LOC_780/B INVX1_LOC_75/A 0.03fF
C51595 INVX1_LOC_17/A NOR2X1_LOC_73/a_36_216# 0.00fF
C51596 INVX1_LOC_89/A NOR2X1_LOC_785/A 0.00fF
C51597 NOR2X1_LOC_178/Y INVX1_LOC_98/A 0.01fF
C51598 NAND2X1_LOC_563/Y INVX1_LOC_217/Y 0.04fF
C51599 NAND2X1_LOC_447/Y INVX1_LOC_23/A 0.03fF
C51600 INVX1_LOC_211/Y INVX1_LOC_90/A 0.06fF
C51601 INVX1_LOC_45/A NAND2X1_LOC_783/A 0.03fF
C51602 NOR2X1_LOC_68/A GATE_479 0.02fF
C51603 NAND2X1_LOC_372/a_36_24# NOR2X1_LOC_303/Y 0.00fF
C51604 INVX1_LOC_223/A NAND2X1_LOC_656/Y 0.07fF
C51605 NOR2X1_LOC_158/Y INVX1_LOC_38/A 0.07fF
C51606 NOR2X1_LOC_536/A NOR2X1_LOC_278/Y 0.03fF
C51607 INVX1_LOC_204/A INVX1_LOC_37/A 0.02fF
C51608 INVX1_LOC_45/A NOR2X1_LOC_130/A 0.06fF
C51609 NOR2X1_LOC_434/Y NOR2X1_LOC_78/A 0.03fF
C51610 D_INPUT_5 INVX1_LOC_92/A 0.03fF
C51611 NAND2X1_LOC_21/Y NAND2X1_LOC_11/Y 0.39fF
C51612 NAND2X1_LOC_77/a_36_24# INVX1_LOC_48/A 0.01fF
C51613 NOR2X1_LOC_226/A NAND2X1_LOC_494/a_36_24# 0.01fF
C51614 INVX1_LOC_21/Y INVX1_LOC_291/A 0.04fF
C51615 NOR2X1_LOC_523/A INPUT_0 0.00fF
C51616 NOR2X1_LOC_725/A NOR2X1_LOC_460/Y 0.05fF
C51617 NAND2X1_LOC_350/A INVX1_LOC_140/A 0.34fF
C51618 INVX1_LOC_268/A INVX1_LOC_105/A 0.00fF
C51619 NOR2X1_LOC_753/Y NAND2X1_LOC_170/A 0.03fF
C51620 INVX1_LOC_78/A INVX1_LOC_54/A 0.37fF
C51621 NOR2X1_LOC_667/A NAND2X1_LOC_811/Y 0.12fF
C51622 INVX1_LOC_17/A NOR2X1_LOC_74/A 0.10fF
C51623 NOR2X1_LOC_658/Y D_GATE_366 0.02fF
C51624 NOR2X1_LOC_604/Y VDD 0.24fF
C51625 NAND2X1_LOC_659/B NOR2X1_LOC_663/A 0.04fF
C51626 INVX1_LOC_32/A NOR2X1_LOC_841/A 0.12fF
C51627 INVX1_LOC_1/A INVX1_LOC_206/Y 0.08fF
C51628 INVX1_LOC_215/A NOR2X1_LOC_152/Y 0.02fF
C51629 NOR2X1_LOC_778/B NOR2X1_LOC_344/a_36_216# 0.00fF
C51630 NOR2X1_LOC_798/A INVX1_LOC_65/A 0.03fF
C51631 INVX1_LOC_35/A NAND2X1_LOC_211/Y 0.07fF
C51632 INVX1_LOC_135/A NOR2X1_LOC_523/B 0.01fF
C51633 NAND2X1_LOC_488/a_36_24# INVX1_LOC_87/A 0.00fF
C51634 INVX1_LOC_251/Y NOR2X1_LOC_709/A 0.02fF
C51635 NOR2X1_LOC_824/A NAND2X1_LOC_623/B 0.08fF
C51636 INVX1_LOC_17/A NOR2X1_LOC_9/Y 1.12fF
C51637 INVX1_LOC_233/Y INVX1_LOC_46/A 0.10fF
C51638 NOR2X1_LOC_471/Y NOR2X1_LOC_74/A 0.09fF
C51639 NOR2X1_LOC_51/A NOR2X1_LOC_25/Y 0.07fF
C51640 INVX1_LOC_71/A NOR2X1_LOC_130/A 0.07fF
C51641 NOR2X1_LOC_273/Y NOR2X1_LOC_214/B 0.03fF
C51642 NOR2X1_LOC_65/B INVX1_LOC_54/A 0.40fF
C51643 NOR2X1_LOC_383/B NOR2X1_LOC_729/A 7.73fF
C51644 INVX1_LOC_305/A NOR2X1_LOC_174/A 0.07fF
C51645 VDD NOR2X1_LOC_663/A 0.12fF
C51646 NOR2X1_LOC_363/Y NOR2X1_LOC_678/A 0.01fF
C51647 NOR2X1_LOC_388/Y NOR2X1_LOC_569/Y 0.13fF
C51648 INVX1_LOC_229/Y NAND2X1_LOC_864/a_36_24# 0.01fF
C51649 INVX1_LOC_34/A NOR2X1_LOC_589/A 2.77fF
C51650 NOR2X1_LOC_607/Y NOR2X1_LOC_355/A 0.03fF
C51651 INVX1_LOC_45/A NOR2X1_LOC_216/Y 0.03fF
C51652 NOR2X1_LOC_214/B NOR2X1_LOC_759/Y 0.00fF
C51653 NOR2X1_LOC_186/Y INVX1_LOC_76/A 0.11fF
C51654 NOR2X1_LOC_234/Y INVX1_LOC_16/A -0.01fF
C51655 INVX1_LOC_240/A INVX1_LOC_22/A 0.30fF
C51656 INVX1_LOC_47/Y INVX1_LOC_63/A 0.52fF
C51657 NAND2X1_LOC_538/Y NOR2X1_LOC_45/B 0.07fF
C51658 INVX1_LOC_13/A NOR2X1_LOC_392/B 0.48fF
C51659 VDD NOR2X1_LOC_674/Y 0.25fF
C51660 INVX1_LOC_45/A NOR2X1_LOC_112/B 0.02fF
C51661 NAND2X1_LOC_175/Y NOR2X1_LOC_841/A 0.10fF
C51662 INVX1_LOC_33/Y NOR2X1_LOC_109/Y 0.09fF
C51663 NOR2X1_LOC_250/A NOR2X1_LOC_45/B 0.02fF
C51664 INVX1_LOC_225/A NOR2X1_LOC_561/Y 0.07fF
C51665 NOR2X1_LOC_297/a_36_216# INVX1_LOC_7/A 0.00fF
C51666 INVX1_LOC_28/A INVX1_LOC_94/A 0.04fF
C51667 NAND2X1_LOC_573/Y INVX1_LOC_76/A 0.13fF
C51668 NAND2X1_LOC_851/a_36_24# INVX1_LOC_141/Y 0.00fF
C51669 NOR2X1_LOC_557/Y NOR2X1_LOC_123/B 0.15fF
C51670 VDD NOR2X1_LOC_384/A -0.00fF
C51671 NOR2X1_LOC_843/A INVX1_LOC_83/A 0.03fF
C51672 NOR2X1_LOC_207/A INVX1_LOC_290/A 0.05fF
C51673 NOR2X1_LOC_68/Y INVX1_LOC_4/Y 0.30fF
C51674 INVX1_LOC_194/A NOR2X1_LOC_459/A 0.02fF
C51675 INVX1_LOC_93/Y NAND2X1_LOC_793/Y 0.01fF
C51676 INVX1_LOC_295/A NOR2X1_LOC_162/Y 0.03fF
C51677 NOR2X1_LOC_48/B INVX1_LOC_42/A 0.24fF
C51678 NOR2X1_LOC_533/A INVX1_LOC_22/A 0.06fF
C51679 NAND2X1_LOC_231/Y NOR2X1_LOC_589/A 0.05fF
C51680 NAND2X1_LOC_724/A INVX1_LOC_76/A 0.10fF
C51681 NOR2X1_LOC_794/B NOR2X1_LOC_600/Y 0.01fF
C51682 NOR2X1_LOC_444/a_36_216# NOR2X1_LOC_862/B 0.15fF
C51683 NOR2X1_LOC_285/Y INVX1_LOC_9/A 0.03fF
C51684 INVX1_LOC_27/A INVX1_LOC_117/A 0.25fF
C51685 NAND2X1_LOC_494/a_36_24# INPUT_1 0.00fF
C51686 NOR2X1_LOC_216/Y INVX1_LOC_71/A 3.57fF
C51687 NOR2X1_LOC_637/B NOR2X1_LOC_329/B 0.06fF
C51688 NAND2X1_LOC_724/Y NAND2X1_LOC_770/Y 0.03fF
C51689 INVX1_LOC_239/A INVX1_LOC_194/Y 0.04fF
C51690 INVX1_LOC_109/Y INVX1_LOC_15/A 0.01fF
C51691 NOR2X1_LOC_180/B NOR2X1_LOC_254/Y 0.18fF
C51692 NAND2X1_LOC_379/a_36_24# GATE_811 0.00fF
C51693 INVX1_LOC_25/Y INVX1_LOC_56/Y 0.01fF
C51694 NOR2X1_LOC_329/B INVX1_LOC_155/A 0.00fF
C51695 NOR2X1_LOC_654/A INVX1_LOC_285/A 0.00fF
C51696 INVX1_LOC_208/A NOR2X1_LOC_188/Y 0.04fF
C51697 NAND2X1_LOC_72/B INVX1_LOC_29/A 0.22fF
C51698 NOR2X1_LOC_654/A INVX1_LOC_265/Y 0.00fF
C51699 NOR2X1_LOC_655/B NOR2X1_LOC_332/A 0.12fF
C51700 INVX1_LOC_61/Y INVX1_LOC_95/Y 0.14fF
C51701 INVX1_LOC_280/Y NOR2X1_LOC_700/Y 0.00fF
C51702 INVX1_LOC_28/A NAND2X1_LOC_465/Y 0.27fF
C51703 NOR2X1_LOC_500/A NOR2X1_LOC_704/Y 0.02fF
C51704 NOR2X1_LOC_234/Y INVX1_LOC_28/A -0.01fF
C51705 NOR2X1_LOC_703/B INVX1_LOC_91/A 0.08fF
C51706 NOR2X1_LOC_45/Y INVX1_LOC_76/A 0.07fF
C51707 INVX1_LOC_161/A INVX1_LOC_20/A 0.17fF
C51708 NOR2X1_LOC_118/a_36_216# INVX1_LOC_306/Y 0.00fF
C51709 INVX1_LOC_12/A NOR2X1_LOC_316/a_36_216# 0.00fF
C51710 INVX1_LOC_239/Y NOR2X1_LOC_299/Y 0.01fF
C51711 INVX1_LOC_45/A NOR2X1_LOC_209/A 0.04fF
C51712 INVX1_LOC_19/A NAND2X1_LOC_97/a_36_24# 0.00fF
C51713 INVX1_LOC_12/A INVX1_LOC_26/A 0.03fF
C51714 INVX1_LOC_78/A NOR2X1_LOC_48/B 0.22fF
C51715 NOR2X1_LOC_607/A NOR2X1_LOC_318/B 0.02fF
C51716 INVX1_LOC_39/A NOR2X1_LOC_99/Y 0.35fF
C51717 INVX1_LOC_128/A INVX1_LOC_32/A -0.02fF
C51718 INVX1_LOC_72/A NOR2X1_LOC_56/Y 0.22fF
C51719 NAND2X1_LOC_640/Y NOR2X1_LOC_167/Y 0.00fF
C51720 INVX1_LOC_256/A INVX1_LOC_202/Y 0.01fF
C51721 NOR2X1_LOC_742/A NOR2X1_LOC_593/a_36_216# 0.01fF
C51722 INVX1_LOC_118/A NOR2X1_LOC_271/B 0.17fF
C51723 INVX1_LOC_218/A NOR2X1_LOC_560/A 0.07fF
C51724 NOR2X1_LOC_647/Y INVX1_LOC_59/Y -0.03fF
C51725 INVX1_LOC_30/A NOR2X1_LOC_40/a_36_216# 0.02fF
C51726 NOR2X1_LOC_91/A NOR2X1_LOC_46/a_36_216# 0.00fF
C51727 NAND2X1_LOC_227/Y NAND2X1_LOC_446/a_36_24# 0.01fF
C51728 NOR2X1_LOC_106/Y NOR2X1_LOC_139/Y 0.01fF
C51729 INVX1_LOC_164/A INVX1_LOC_10/A 0.01fF
C51730 INVX1_LOC_50/A NOR2X1_LOC_189/a_36_216# 0.00fF
C51731 NAND2X1_LOC_51/B INVX1_LOC_266/Y 0.05fF
C51732 INVX1_LOC_104/A NOR2X1_LOC_188/A 0.04fF
C51733 INVX1_LOC_225/A NOR2X1_LOC_167/Y 0.02fF
C51734 NOR2X1_LOC_768/a_36_216# INVX1_LOC_16/A 0.01fF
C51735 NAND2X1_LOC_866/B GATE_865 0.01fF
C51736 NAND2X1_LOC_149/Y NOR2X1_LOC_155/A 0.09fF
C51737 NOR2X1_LOC_273/Y NOR2X1_LOC_275/A 0.08fF
C51738 INVX1_LOC_21/A NAND2X1_LOC_288/A 0.40fF
C51739 NOR2X1_LOC_759/Y NOR2X1_LOC_275/A 0.01fF
C51740 INVX1_LOC_13/A INVX1_LOC_90/A 0.07fF
C51741 NOR2X1_LOC_255/Y INVX1_LOC_12/A 0.50fF
C51742 INVX1_LOC_72/A VDD 4.95fF
C51743 NAND2X1_LOC_9/Y NAND2X1_LOC_81/B 0.03fF
C51744 NOR2X1_LOC_716/B INVX1_LOC_70/Y 0.03fF
C51745 INVX1_LOC_142/Y VDD -0.00fF
C51746 INVX1_LOC_311/A INVX1_LOC_266/Y 0.10fF
C51747 INVX1_LOC_236/Y NOR2X1_LOC_536/A 0.01fF
C51748 INVX1_LOC_233/A NAND2X1_LOC_81/B 0.07fF
C51749 INVX1_LOC_64/A INVX1_LOC_49/Y 0.03fF
C51750 NOR2X1_LOC_721/Y NOR2X1_LOC_537/Y 0.03fF
C51751 INVX1_LOC_72/A NAND2X1_LOC_800/A 0.32fF
C51752 INVX1_LOC_284/Y NOR2X1_LOC_536/A 0.04fF
C51753 NAND2X1_LOC_338/B NOR2X1_LOC_721/Y 0.10fF
C51754 INVX1_LOC_36/A INVX1_LOC_33/Y 0.06fF
C51755 NOR2X1_LOC_503/Y INVX1_LOC_54/A 0.03fF
C51756 INVX1_LOC_21/A NOR2X1_LOC_653/Y 0.03fF
C51757 INVX1_LOC_198/Y VDD 1.47fF
C51758 NAND2X1_LOC_364/a_36_24# INVX1_LOC_132/Y 0.00fF
C51759 INVX1_LOC_58/A INVX1_LOC_170/Y 0.01fF
C51760 INVX1_LOC_75/A INVX1_LOC_56/Y 0.03fF
C51761 NOR2X1_LOC_332/A NOR2X1_LOC_846/B 0.02fF
C51762 NAND2X1_LOC_842/B NAND2X1_LOC_573/A 0.09fF
C51763 INVX1_LOC_64/A INVX1_LOC_99/A 0.08fF
C51764 NOR2X1_LOC_283/a_36_216# INVX1_LOC_20/A 0.01fF
C51765 NOR2X1_LOC_658/Y NOR2X1_LOC_142/a_36_216# 0.01fF
C51766 NOR2X1_LOC_764/a_36_216# D_INPUT_4 0.00fF
C51767 INVX1_LOC_78/A NOR2X1_LOC_438/Y 0.03fF
C51768 INVX1_LOC_64/A NOR2X1_LOC_672/a_36_216# 0.00fF
C51769 INVX1_LOC_17/A NOR2X1_LOC_865/Y 0.04fF
C51770 NOR2X1_LOC_246/A INVX1_LOC_90/A 0.11fF
C51771 INVX1_LOC_13/A NAND2X1_LOC_348/A 0.72fF
C51772 NOR2X1_LOC_447/Y NOR2X1_LOC_447/B 0.06fF
C51773 INVX1_LOC_21/A INVX1_LOC_19/A 0.34fF
C51774 NOR2X1_LOC_240/Y NOR2X1_LOC_240/B 0.04fF
C51775 INVX1_LOC_17/A NOR2X1_LOC_243/B 0.05fF
C51776 NOR2X1_LOC_246/A NOR2X1_LOC_389/B 0.01fF
C51777 NOR2X1_LOC_577/Y NOR2X1_LOC_137/Y 0.04fF
C51778 NOR2X1_LOC_83/Y INVX1_LOC_16/A 0.04fF
C51779 INVX1_LOC_89/A NOR2X1_LOC_702/Y 0.02fF
C51780 INVX1_LOC_53/A D_INPUT_5 0.04fF
C51781 INVX1_LOC_202/A INVX1_LOC_12/Y 0.04fF
C51782 INVX1_LOC_34/A INVX1_LOC_20/A 0.54fF
C51783 NOR2X1_LOC_381/a_36_216# NOR2X1_LOC_332/A 0.01fF
C51784 NAND2X1_LOC_860/Y INVX1_LOC_286/A 0.02fF
C51785 INVX1_LOC_50/A INVX1_LOC_271/Y 0.07fF
C51786 INVX1_LOC_232/A INVX1_LOC_6/A 0.03fF
C51787 NOR2X1_LOC_523/B INVX1_LOC_280/A 0.01fF
C51788 INVX1_LOC_90/A INVX1_LOC_55/Y 0.03fF
C51789 INVX1_LOC_225/A INVX1_LOC_76/A 0.10fF
C51790 INVX1_LOC_103/A NAND2X1_LOC_476/Y 0.02fF
C51791 NOR2X1_LOC_191/A NOR2X1_LOC_192/A 0.00fF
C51792 INVX1_LOC_24/A NOR2X1_LOC_331/B 0.16fF
C51793 NAND2X1_LOC_9/Y INVX1_LOC_4/Y 0.05fF
C51794 INVX1_LOC_10/A NOR2X1_LOC_313/Y 0.02fF
C51795 NOR2X1_LOC_68/A NOR2X1_LOC_641/Y 0.02fF
C51796 NOR2X1_LOC_383/Y INVX1_LOC_6/A 0.07fF
C51797 INVX1_LOC_103/A INVX1_LOC_186/Y 0.10fF
C51798 NOR2X1_LOC_576/B INVX1_LOC_282/A 0.03fF
C51799 INVX1_LOC_45/A NOR2X1_LOC_197/B 0.01fF
C51800 NAND2X1_LOC_214/B INVX1_LOC_3/Y 0.10fF
C51801 NAND2X1_LOC_231/Y INVX1_LOC_147/Y 0.02fF
C51802 NOR2X1_LOC_666/A INVX1_LOC_12/A 0.06fF
C51803 NOR2X1_LOC_718/B INVX1_LOC_139/Y 0.01fF
C51804 NAND2X1_LOC_741/B NAND2X1_LOC_810/B 0.45fF
C51805 NOR2X1_LOC_713/a_36_216# INVX1_LOC_174/Y 0.00fF
C51806 NOR2X1_LOC_568/A NOR2X1_LOC_197/B 0.10fF
C51807 NOR2X1_LOC_131/A NAND2X1_LOC_469/B 0.01fF
C51808 INVX1_LOC_57/A NAND2X1_LOC_99/A 0.07fF
C51809 INVX1_LOC_269/A NAND2X1_LOC_74/B 0.01fF
C51810 NOR2X1_LOC_209/Y INVX1_LOC_76/A 0.07fF
C51811 NOR2X1_LOC_366/Y INVX1_LOC_6/A 0.02fF
C51812 NOR2X1_LOC_360/Y INVX1_LOC_92/A 0.16fF
C51813 INVX1_LOC_27/A INVX1_LOC_3/Y 0.09fF
C51814 NOR2X1_LOC_152/Y INVX1_LOC_54/A 0.84fF
C51815 NOR2X1_LOC_309/Y INVX1_LOC_33/Y 0.01fF
C51816 VDD INVX1_LOC_192/Y 0.35fF
C51817 NOR2X1_LOC_361/B INVX1_LOC_284/A 0.10fF
C51818 NOR2X1_LOC_231/a_36_216# NOR2X1_LOC_814/A 0.01fF
C51819 NOR2X1_LOC_231/B INVX1_LOC_63/A 0.01fF
C51820 NOR2X1_LOC_824/A INVX1_LOC_3/Y 0.01fF
C51821 VDD NOR2X1_LOC_537/Y 0.43fF
C51822 INVX1_LOC_269/A NOR2X1_LOC_847/B -0.01fF
C51823 INVX1_LOC_113/Y INVX1_LOC_54/A 0.01fF
C51824 INVX1_LOC_286/A NAND2X1_LOC_861/Y 0.06fF
C51825 NAND2X1_LOC_338/B VDD 0.15fF
C51826 NAND2X1_LOC_852/Y INVX1_LOC_76/A 0.01fF
C51827 INVX1_LOC_24/A NOR2X1_LOC_491/Y 0.03fF
C51828 INVX1_LOC_28/A INVX1_LOC_144/A 0.08fF
C51829 NOR2X1_LOC_526/Y INVX1_LOC_46/A 0.03fF
C51830 NAND2X1_LOC_577/A NOR2X1_LOC_662/A 0.07fF
C51831 NOR2X1_LOC_203/Y INVX1_LOC_14/Y 0.04fF
C51832 NOR2X1_LOC_798/A INVX1_LOC_4/Y 0.09fF
C51833 INVX1_LOC_58/A INVX1_LOC_271/A 0.03fF
C51834 NOR2X1_LOC_561/Y NAND2X1_LOC_642/Y 0.01fF
C51835 INVX1_LOC_58/A INVX1_LOC_105/Y 0.01fF
C51836 NAND2X1_LOC_323/B VDD 0.31fF
C51837 NAND2X1_LOC_733/Y NOR2X1_LOC_36/B 0.17fF
C51838 INVX1_LOC_83/A NOR2X1_LOC_595/Y 0.01fF
C51839 NOR2X1_LOC_42/a_36_216# INVX1_LOC_316/Y 0.01fF
C51840 NOR2X1_LOC_337/Y INVX1_LOC_313/Y 0.01fF
C51841 NAND2X1_LOC_45/Y NOR2X1_LOC_78/A 0.07fF
C51842 NAND2X1_LOC_842/B NOR2X1_LOC_183/a_36_216# 0.00fF
C51843 NAND2X1_LOC_361/Y NOR2X1_LOC_624/B 0.02fF
C51844 INVX1_LOC_236/A INVX1_LOC_38/A 1.29fF
C51845 NAND2X1_LOC_200/B INVX1_LOC_117/A 0.12fF
C51846 NOR2X1_LOC_503/Y NOR2X1_LOC_48/B 0.13fF
C51847 NAND2X1_LOC_318/a_36_24# NOR2X1_LOC_536/A 0.00fF
C51848 INVX1_LOC_310/Y NOR2X1_LOC_634/A 0.02fF
C51849 INVX1_LOC_83/A INVX1_LOC_115/Y 0.01fF
C51850 INVX1_LOC_181/A INVX1_LOC_306/Y 0.01fF
C51851 INVX1_LOC_21/A INVX1_LOC_26/Y 0.10fF
C51852 NOR2X1_LOC_441/Y INVX1_LOC_42/A 0.06fF
C51853 NOR2X1_LOC_753/Y INVX1_LOC_250/Y 0.03fF
C51854 INVX1_LOC_80/A D_INPUT_3 0.01fF
C51855 INVX1_LOC_137/A INVX1_LOC_117/A 0.17fF
C51856 NOR2X1_LOC_804/B INVX1_LOC_220/A 0.28fF
C51857 INVX1_LOC_30/A NAND2X1_LOC_254/Y 0.48fF
C51858 INVX1_LOC_21/A INVX1_LOC_166/A 0.21fF
C51859 NAND2X1_LOC_198/B INVX1_LOC_29/A 0.84fF
C51860 NOR2X1_LOC_228/a_36_216# INVX1_LOC_63/A 0.01fF
C51861 INVX1_LOC_140/A INVX1_LOC_291/Y 0.01fF
C51862 NOR2X1_LOC_518/Y INVX1_LOC_102/A 0.06fF
C51863 INVX1_LOC_13/A INVX1_LOC_38/A 0.07fF
C51864 INVX1_LOC_90/A NOR2X1_LOC_357/Y 0.03fF
C51865 NOR2X1_LOC_272/Y D_INPUT_1 0.10fF
C51866 INVX1_LOC_58/A INVX1_LOC_27/A 2.33fF
C51867 NAND2X1_LOC_451/Y INVX1_LOC_92/A 1.24fF
C51868 INVX1_LOC_2/A NOR2X1_LOC_58/a_36_216# 0.00fF
C51869 NAND2X1_LOC_860/Y INVX1_LOC_54/A 0.01fF
C51870 INVX1_LOC_256/Y INVX1_LOC_70/A 0.09fF
C51871 INVX1_LOC_58/A NOR2X1_LOC_824/A 0.07fF
C51872 INVX1_LOC_64/A NOR2X1_LOC_411/Y 0.08fF
C51873 INVX1_LOC_223/Y NOR2X1_LOC_790/B 0.04fF
C51874 NOR2X1_LOC_310/a_36_216# NOR2X1_LOC_405/A 0.00fF
C51875 INVX1_LOC_313/Y VDD 2.15fF
C51876 NOR2X1_LOC_769/B NAND2X1_LOC_149/Y 0.04fF
C51877 INVX1_LOC_7/A NOR2X1_LOC_271/Y 0.00fF
C51878 INVX1_LOC_309/A INVX1_LOC_91/A 0.03fF
C51879 NAND2X1_LOC_830/a_36_24# INVX1_LOC_46/A 0.00fF
C51880 NOR2X1_LOC_525/Y NOR2X1_LOC_536/A 0.01fF
C51881 NOR2X1_LOC_598/B NAND2X1_LOC_149/Y 0.25fF
C51882 NOR2X1_LOC_815/Y INVX1_LOC_272/A 0.02fF
C51883 NOR2X1_LOC_441/Y INVX1_LOC_78/A 0.90fF
C51884 NOR2X1_LOC_312/Y NOR2X1_LOC_536/A 0.01fF
C51885 NAND2X1_LOC_553/A NAND2X1_LOC_540/a_36_24# 0.02fF
C51886 NOR2X1_LOC_130/A NOR2X1_LOC_331/B 0.10fF
C51887 NOR2X1_LOC_210/A NAND2X1_LOC_93/B 0.02fF
C51888 INVX1_LOC_215/A INVX1_LOC_291/A 0.20fF
C51889 INVX1_LOC_16/A NOR2X1_LOC_155/A 0.07fF
C51890 INVX1_LOC_232/Y NOR2X1_LOC_649/B 1.51fF
C51891 INVX1_LOC_11/Y INVX1_LOC_309/A 0.03fF
C51892 NOR2X1_LOC_132/Y INVX1_LOC_284/A 0.03fF
C51893 NOR2X1_LOC_152/Y NOR2X1_LOC_48/B 0.09fF
C51894 INVX1_LOC_77/A NOR2X1_LOC_640/B 0.01fF
C51895 INVX1_LOC_232/Y INVX1_LOC_3/A 1.24fF
C51896 NOR2X1_LOC_745/Y INVX1_LOC_275/Y 0.01fF
C51897 INPUT_0 INVX1_LOC_20/A 0.36fF
C51898 NOR2X1_LOC_528/Y NAND2X1_LOC_623/B 0.08fF
C51899 NOR2X1_LOC_667/A NOR2X1_LOC_653/Y 0.03fF
C51900 NOR2X1_LOC_272/Y NOR2X1_LOC_652/Y 0.10fF
C51901 NAND2X1_LOC_578/B INVX1_LOC_203/A 0.34fF
C51902 NAND2X1_LOC_35/Y INVX1_LOC_48/Y 0.02fF
C51903 NOR2X1_LOC_210/A NAND2X1_LOC_425/Y 0.04fF
C51904 NOR2X1_LOC_719/B NOR2X1_LOC_78/Y 0.08fF
C51905 NOR2X1_LOC_82/Y NAND2X1_LOC_572/B 0.01fF
C51906 INVX1_LOC_269/A NOR2X1_LOC_660/Y 0.03fF
C51907 NAND2X1_LOC_861/Y INVX1_LOC_54/A 0.04fF
C51908 NOR2X1_LOC_65/B NOR2X1_LOC_441/Y 0.67fF
C51909 NOR2X1_LOC_311/Y NOR2X1_LOC_595/Y 0.22fF
C51910 NAND2X1_LOC_552/A NAND2X1_LOC_579/A 0.01fF
C51911 INVX1_LOC_254/Y INVX1_LOC_15/A 0.12fF
C51912 INVX1_LOC_36/A INVX1_LOC_23/Y 0.08fF
C51913 NOR2X1_LOC_846/Y NAND2X1_LOC_473/A 0.01fF
C51914 NOR2X1_LOC_667/A INVX1_LOC_19/A 1.94fF
C51915 NOR2X1_LOC_589/a_36_216# INVX1_LOC_117/A 0.01fF
C51916 NOR2X1_LOC_78/B NOR2X1_LOC_856/B 0.03fF
C51917 NOR2X1_LOC_130/A NOR2X1_LOC_592/B 2.34fF
C51918 NOR2X1_LOC_845/A NOR2X1_LOC_35/Y 0.46fF
C51919 NOR2X1_LOC_216/Y NOR2X1_LOC_331/B 0.01fF
C51920 NOR2X1_LOC_369/Y NAND2X1_LOC_793/B 0.04fF
C51921 NOR2X1_LOC_268/a_36_216# NAND2X1_LOC_61/Y -0.00fF
C51922 INVX1_LOC_24/A NOR2X1_LOC_621/B 0.08fF
C51923 NOR2X1_LOC_664/Y INVX1_LOC_3/Y 0.03fF
C51924 NAND2X1_LOC_579/A INVX1_LOC_178/A 0.10fF
C51925 NOR2X1_LOC_590/A INVX1_LOC_58/Y 0.10fF
C51926 INVX1_LOC_34/A INVX1_LOC_4/A 0.04fF
C51927 NAND2X1_LOC_25/a_36_24# INVX1_LOC_174/A 0.01fF
C51928 NOR2X1_LOC_528/a_36_216# INVX1_LOC_119/Y 0.02fF
C51929 INVX1_LOC_64/A INVX1_LOC_161/A 0.10fF
C51930 NOR2X1_LOC_15/Y NOR2X1_LOC_440/B 0.94fF
C51931 INVX1_LOC_280/Y INVX1_LOC_284/A 0.66fF
C51932 NAND2X1_LOC_642/Y INVX1_LOC_76/A 0.01fF
C51933 NOR2X1_LOC_655/B INVX1_LOC_42/A 0.76fF
C51934 INVX1_LOC_11/A NOR2X1_LOC_460/Y 0.08fF
C51935 INVX1_LOC_316/Y NOR2X1_LOC_671/a_36_216# 0.00fF
C51936 INVX1_LOC_53/Y INVX1_LOC_29/A 0.08fF
C51937 INVX1_LOC_64/A NAND2X1_LOC_208/B 0.29fF
C51938 INVX1_LOC_28/A NOR2X1_LOC_155/A 0.16fF
C51939 INVX1_LOC_181/Y NOR2X1_LOC_383/B 0.08fF
C51940 D_INPUT_1 NAND2X1_LOC_364/A 0.03fF
C51941 INVX1_LOC_223/A NOR2X1_LOC_717/A 0.10fF
C51942 NAND2X1_LOC_563/A NOR2X1_LOC_847/B -0.00fF
C51943 INVX1_LOC_135/A NAND2X1_LOC_206/Y 0.12fF
C51944 NOR2X1_LOC_338/Y INVX1_LOC_271/A 0.00fF
C51945 NOR2X1_LOC_237/Y INVX1_LOC_23/Y 0.01fF
C51946 NOR2X1_LOC_322/Y NOR2X1_LOC_487/Y 0.02fF
C51947 NAND2X1_LOC_579/A NOR2X1_LOC_494/Y 0.02fF
C51948 INVX1_LOC_24/Y INVX1_LOC_1/A 0.10fF
C51949 INVX1_LOC_21/A INVX1_LOC_161/Y 0.09fF
C51950 NAND2X1_LOC_656/A INVX1_LOC_57/A 0.17fF
C51951 NOR2X1_LOC_312/Y NOR2X1_LOC_661/A 0.03fF
C51952 NOR2X1_LOC_360/Y INVX1_LOC_53/A 0.10fF
C51953 INVX1_LOC_135/A NAND2X1_LOC_773/B 0.27fF
C51954 NOR2X1_LOC_790/B NAND2X1_LOC_167/a_36_24# 0.01fF
C51955 NOR2X1_LOC_560/A NAND2X1_LOC_206/Y 0.06fF
C51956 INVX1_LOC_75/A NOR2X1_LOC_831/B 0.96fF
C51957 INVX1_LOC_90/A NAND2X1_LOC_489/Y 0.10fF
C51958 INVX1_LOC_58/A INVX1_LOC_249/A 0.07fF
C51959 NAND2X1_LOC_796/B INVX1_LOC_31/A 0.03fF
C51960 NOR2X1_LOC_778/a_36_216# NOR2X1_LOC_383/B 0.00fF
C51961 NOR2X1_LOC_577/Y NOR2X1_LOC_677/Y 0.04fF
C51962 NAND2X1_LOC_579/A NOR2X1_LOC_816/A 0.01fF
C51963 INVX1_LOC_120/A NOR2X1_LOC_777/B 0.00fF
C51964 INVX1_LOC_21/A INVX1_LOC_312/A 0.01fF
C51965 NOR2X1_LOC_346/a_36_216# NAND2X1_LOC_206/Y 0.01fF
C51966 INVX1_LOC_17/A NOR2X1_LOC_250/Y 1.17fF
C51967 NAND2X1_LOC_36/A D_INPUT_6 0.01fF
C51968 INVX1_LOC_36/A NOR2X1_LOC_846/A 0.07fF
C51969 INVX1_LOC_193/Y NAND2X1_LOC_425/Y 0.04fF
C51970 NAND2X1_LOC_354/B NOR2X1_LOC_654/A 0.49fF
C51971 NAND2X1_LOC_364/A NOR2X1_LOC_108/a_36_216# 0.00fF
C51972 INVX1_LOC_1/Y INVX1_LOC_47/Y 0.90fF
C51973 INVX1_LOC_50/A NOR2X1_LOC_144/Y 0.01fF
C51974 NAND2X1_LOC_656/Y INVX1_LOC_290/Y 0.08fF
C51975 NAND2X1_LOC_364/A NOR2X1_LOC_652/Y 0.11fF
C51976 NOR2X1_LOC_82/A NAND2X1_LOC_793/Y 0.41fF
C51977 INVX1_LOC_41/A INVX1_LOC_25/A 0.07fF
C51978 INVX1_LOC_85/A NOR2X1_LOC_727/B 0.05fF
C51979 NOR2X1_LOC_99/B INVX1_LOC_42/A 0.31fF
C51980 NAND2X1_LOC_842/B NAND2X1_LOC_81/B 0.03fF
C51981 INVX1_LOC_83/A NAND2X1_LOC_214/a_36_24# 0.01fF
C51982 NAND2X1_LOC_139/A INVX1_LOC_23/A 0.11fF
C51983 INVX1_LOC_25/A INVX1_LOC_201/Y 0.11fF
C51984 INVX1_LOC_226/Y NAND2X1_LOC_471/Y 0.00fF
C51985 NAND2X1_LOC_357/A NAND2X1_LOC_352/B 0.04fF
C51986 INVX1_LOC_234/A INVX1_LOC_3/Y 0.20fF
C51987 NOR2X1_LOC_335/B INVX1_LOC_84/A 0.04fF
C51988 NAND2X1_LOC_350/A NOR2X1_LOC_503/Y 0.07fF
C51989 NOR2X1_LOC_506/Y NOR2X1_LOC_56/Y 0.01fF
C51990 INVX1_LOC_245/Y NOR2X1_LOC_471/Y 0.90fF
C51991 NAND2X1_LOC_783/Y NAND2X1_LOC_803/B 0.03fF
C51992 NAND2X1_LOC_287/B NOR2X1_LOC_536/A 0.02fF
C51993 NOR2X1_LOC_92/Y NOR2X1_LOC_384/Y 0.07fF
C51994 NAND2X1_LOC_778/Y INVX1_LOC_41/Y 0.03fF
C51995 NOR2X1_LOC_357/Y INVX1_LOC_38/A 0.03fF
C51996 INPUT_0 NOR2X1_LOC_68/a_36_216# 0.00fF
C51997 NOR2X1_LOC_65/B NOR2X1_LOC_655/B 0.10fF
C51998 NOR2X1_LOC_504/Y INVX1_LOC_296/Y 0.07fF
C51999 INVX1_LOC_83/A D_INPUT_5 0.10fF
C52000 INVX1_LOC_35/A NAND2X1_LOC_569/A 0.21fF
C52001 NAND2X1_LOC_51/B INVX1_LOC_19/A 0.05fF
C52002 NOR2X1_LOC_635/A INPUT_6 0.01fF
C52003 INVX1_LOC_64/A INVX1_LOC_34/A 0.16fF
C52004 NOR2X1_LOC_272/Y NOR2X1_LOC_403/B 0.10fF
C52005 INVX1_LOC_13/A NAND2X1_LOC_223/A 0.44fF
C52006 NOR2X1_LOC_332/A NOR2X1_LOC_28/a_36_216# 0.01fF
C52007 INVX1_LOC_136/A INVX1_LOC_269/A 0.13fF
C52008 NOR2X1_LOC_536/A INVX1_LOC_129/Y 0.01fF
C52009 INVX1_LOC_10/Y NAND2X1_LOC_472/Y 0.03fF
C52010 NOR2X1_LOC_211/A INVX1_LOC_116/Y 0.00fF
C52011 INVX1_LOC_135/A NOR2X1_LOC_297/A 0.01fF
C52012 NAND2X1_LOC_783/Y NOR2X1_LOC_590/A 0.01fF
C52013 INVX1_LOC_136/A NOR2X1_LOC_232/Y 0.01fF
C52014 NOR2X1_LOC_420/Y NAND2X1_LOC_361/Y 0.11fF
C52015 NOR2X1_LOC_179/Y INVX1_LOC_91/A 0.01fF
C52016 INVX1_LOC_43/Y NAND2X1_LOC_208/B 0.19fF
C52017 INVX1_LOC_90/A INVX1_LOC_32/A 0.08fF
C52018 INVX1_LOC_103/A INVX1_LOC_18/A 0.17fF
C52019 INVX1_LOC_298/Y NOR2X1_LOC_665/A 0.02fF
C52020 VDD NOR2X1_LOC_506/Y 0.11fF
C52021 NOR2X1_LOC_15/Y INVX1_LOC_41/Y 0.10fF
C52022 INVX1_LOC_144/A INVX1_LOC_109/A 0.05fF
C52023 INVX1_LOC_53/Y NOR2X1_LOC_318/a_36_216# 0.00fF
C52024 NOR2X1_LOC_389/B INVX1_LOC_32/A 0.03fF
C52025 INVX1_LOC_84/A INVX1_LOC_264/Y 0.09fF
C52026 NAND2X1_LOC_728/Y INVX1_LOC_103/A 0.16fF
C52027 NAND2X1_LOC_451/Y INVX1_LOC_53/A 0.09fF
C52028 NAND2X1_LOC_849/A NOR2X1_LOC_490/a_36_216# 0.00fF
C52029 INVX1_LOC_213/Y INVX1_LOC_5/A 0.08fF
C52030 NOR2X1_LOC_772/Y INVX1_LOC_171/Y 0.11fF
C52031 INVX1_LOC_164/Y NAND2X1_LOC_860/A 0.04fF
C52032 NOR2X1_LOC_155/A NOR2X1_LOC_35/Y 0.03fF
C52033 NOR2X1_LOC_313/Y INVX1_LOC_12/A 0.02fF
C52034 INVX1_LOC_36/A NOR2X1_LOC_596/Y 0.01fF
C52035 NOR2X1_LOC_843/A NOR2X1_LOC_798/A 0.30fF
C52036 INVX1_LOC_38/A NOR2X1_LOC_692/Y 0.01fF
C52037 NAND2X1_LOC_35/Y NOR2X1_LOC_84/Y 0.10fF
C52038 INVX1_LOC_311/Y INVX1_LOC_15/A 0.03fF
C52039 NOR2X1_LOC_19/B INVX1_LOC_3/Y 0.76fF
C52040 INVX1_LOC_15/Y NAND2X1_LOC_624/B 0.15fF
C52041 NAND2X1_LOC_549/B NOR2X1_LOC_392/Y 0.01fF
C52042 INVX1_LOC_197/Y NOR2X1_LOC_476/B 0.32fF
C52043 INVX1_LOC_64/A NAND2X1_LOC_231/Y 0.10fF
C52044 NOR2X1_LOC_215/A NOR2X1_LOC_142/Y 0.08fF
C52045 NOR2X1_LOC_831/B NOR2X1_LOC_309/a_36_216# 0.01fF
C52046 NOR2X1_LOC_315/Y INVX1_LOC_306/Y 0.10fF
C52047 NOR2X1_LOC_254/A NOR2X1_LOC_68/A 0.07fF
C52048 NAND2X1_LOC_717/Y NAND2X1_LOC_725/A 0.03fF
C52049 NOR2X1_LOC_392/B INVX1_LOC_171/Y 0.03fF
C52050 NOR2X1_LOC_637/Y INVX1_LOC_103/A 0.05fF
C52051 INVX1_LOC_45/A INVX1_LOC_286/Y 0.00fF
C52052 INVX1_LOC_292/A INVX1_LOC_18/A 0.07fF
C52053 NAND2X1_LOC_648/A NOR2X1_LOC_409/B 0.01fF
C52054 NOR2X1_LOC_130/A NOR2X1_LOC_449/A 0.03fF
C52055 INVX1_LOC_37/A NAND2X1_LOC_244/a_36_24# 0.01fF
C52056 INVX1_LOC_129/Y NAND2X1_LOC_93/B 0.03fF
C52057 NAND2X1_LOC_563/A NOR2X1_LOC_660/Y 0.23fF
C52058 NAND2X1_LOC_112/Y INVX1_LOC_23/A 0.07fF
C52059 INVX1_LOC_177/A NOR2X1_LOC_674/Y 0.01fF
C52060 NOR2X1_LOC_321/Y NAND2X1_LOC_332/Y 0.03fF
C52061 INVX1_LOC_286/Y NAND2X1_LOC_856/A 0.04fF
C52062 INVX1_LOC_233/A NAND2X1_LOC_862/A 0.04fF
C52063 NOR2X1_LOC_91/A NAND2X1_LOC_474/a_36_24# 0.01fF
C52064 INVX1_LOC_50/A INVX1_LOC_279/A 0.14fF
C52065 NAND2X1_LOC_348/A INVX1_LOC_32/A 0.03fF
C52066 INVX1_LOC_90/A NAND2X1_LOC_175/Y 0.09fF
C52067 NOR2X1_LOC_598/B INVX1_LOC_16/A 0.03fF
C52068 NAND2X1_LOC_861/Y NOR2X1_LOC_438/Y 0.19fF
C52069 NOR2X1_LOC_273/Y NOR2X1_LOC_160/B 0.03fF
C52070 INVX1_LOC_36/A NAND2X1_LOC_741/B 3.85fF
C52071 INVX1_LOC_41/A INVX1_LOC_1/A 0.28fF
C52072 INVX1_LOC_35/A INVX1_LOC_316/Y 0.03fF
C52073 NOR2X1_LOC_626/Y INVX1_LOC_266/Y 0.06fF
C52074 NOR2X1_LOC_65/B NOR2X1_LOC_99/B 0.02fF
C52075 INVX1_LOC_224/A NAND2X1_LOC_524/a_36_24# 0.00fF
C52076 NOR2X1_LOC_160/B NOR2X1_LOC_759/Y 0.03fF
C52077 INVX1_LOC_120/A NOR2X1_LOC_843/B 0.03fF
C52078 INVX1_LOC_201/Y INVX1_LOC_1/A 0.23fF
C52079 INVX1_LOC_304/A INVX1_LOC_19/A 0.07fF
C52080 NOR2X1_LOC_825/Y INVX1_LOC_84/A 0.15fF
C52081 INVX1_LOC_182/A INVX1_LOC_78/A 0.07fF
C52082 INVX1_LOC_202/A NOR2X1_LOC_160/B 0.07fF
C52083 INVX1_LOC_5/A NAND2X1_LOC_341/a_36_24# 0.00fF
C52084 INVX1_LOC_58/A INVX1_LOC_234/A 0.55fF
C52085 INVX1_LOC_58/A NAND2X1_LOC_156/B 0.01fF
C52086 NAND2X1_LOC_579/A NAND2X1_LOC_562/B 0.01fF
C52087 NAND2X1_LOC_725/A INVX1_LOC_16/A 0.05fF
C52088 NAND2X1_LOC_149/Y NOR2X1_LOC_156/B 0.05fF
C52089 INPUT_0 INVX1_LOC_4/A 0.05fF
C52090 NOR2X1_LOC_443/Y INVX1_LOC_89/A 0.02fF
C52091 INVX1_LOC_45/A INVX1_LOC_159/A 0.03fF
C52092 NOR2X1_LOC_750/Y INVX1_LOC_7/A 0.04fF
C52093 NOR2X1_LOC_536/Y INVX1_LOC_240/A 0.06fF
C52094 NAND2X1_LOC_766/a_36_24# INVX1_LOC_174/A 0.00fF
C52095 INPUT_4 NOR2X1_LOC_18/a_36_216# 0.01fF
C52096 NOR2X1_LOC_590/A NOR2X1_LOC_419/Y 0.07fF
C52097 NOR2X1_LOC_599/Y NOR2X1_LOC_387/Y 0.07fF
C52098 NOR2X1_LOC_331/B NOR2X1_LOC_197/B 0.03fF
C52099 INVX1_LOC_291/A INVX1_LOC_54/A 0.07fF
C52100 NOR2X1_LOC_590/A NOR2X1_LOC_537/A 0.01fF
C52101 INVX1_LOC_45/A NOR2X1_LOC_191/B 0.02fF
C52102 NOR2X1_LOC_441/Y NOR2X1_LOC_152/Y 0.10fF
C52103 NAND2X1_LOC_708/Y INPUT_5 0.00fF
C52104 NOR2X1_LOC_296/Y NOR2X1_LOC_392/B 0.12fF
C52105 INVX1_LOC_50/A NOR2X1_LOC_166/a_36_216# 0.00fF
C52106 NOR2X1_LOC_813/Y NOR2X1_LOC_813/a_36_216# 0.00fF
C52107 NAND2X1_LOC_357/A NAND2X1_LOC_357/B 0.19fF
C52108 INVX1_LOC_314/Y INVX1_LOC_30/A 0.15fF
C52109 INVX1_LOC_34/A INVX1_LOC_43/Y 0.03fF
C52110 INVX1_LOC_90/A NOR2X1_LOC_622/A 0.01fF
C52111 NAND2X1_LOC_860/A NOR2X1_LOC_76/A 0.03fF
C52112 INVX1_LOC_152/Y NOR2X1_LOC_99/B 0.02fF
C52113 INVX1_LOC_200/A NOR2X1_LOC_369/a_36_216# 0.00fF
C52114 NOR2X1_LOC_138/a_36_216# NAND2X1_LOC_82/Y 0.00fF
C52115 NOR2X1_LOC_689/Y INVX1_LOC_28/A 0.72fF
C52116 NOR2X1_LOC_384/Y NAND2X1_LOC_837/Y 0.21fF
C52117 INVX1_LOC_33/Y INVX1_LOC_63/A 0.05fF
C52118 NOR2X1_LOC_859/A NOR2X1_LOC_860/B 0.01fF
C52119 INVX1_LOC_93/A NAND2X1_LOC_390/A 0.17fF
C52120 NOR2X1_LOC_361/B NAND2X1_LOC_338/B 0.10fF
C52121 NAND2X1_LOC_579/A NOR2X1_LOC_773/Y 0.03fF
C52122 NOR2X1_LOC_329/B INVX1_LOC_57/A 0.00fF
C52123 INVX1_LOC_31/A NAND2X1_LOC_139/A 0.01fF
C52124 INVX1_LOC_239/A NOR2X1_LOC_375/Y 0.01fF
C52125 INVX1_LOC_50/A INVX1_LOC_182/Y 0.15fF
C52126 NOR2X1_LOC_522/a_36_216# NAND2X1_LOC_837/Y 0.00fF
C52127 INVX1_LOC_280/A NAND2X1_LOC_206/Y 1.60fF
C52128 INVX1_LOC_93/Y INVX1_LOC_47/Y 1.41fF
C52129 NOR2X1_LOC_74/A INVX1_LOC_181/A 0.01fF
C52130 INVX1_LOC_89/A INVX1_LOC_213/A 0.01fF
C52131 INVX1_LOC_12/Y NAND2X1_LOC_74/B 0.01fF
C52132 INVX1_LOC_1/A NOR2X1_LOC_211/A 0.04fF
C52133 INVX1_LOC_214/A INVX1_LOC_161/Y 0.02fF
C52134 NOR2X1_LOC_778/B NOR2X1_LOC_457/A 0.02fF
C52135 VDD NOR2X1_LOC_226/Y 0.18fF
C52136 NOR2X1_LOC_703/A INVX1_LOC_58/Y 0.00fF
C52137 NOR2X1_LOC_220/B INVX1_LOC_171/A 0.01fF
C52138 NOR2X1_LOC_567/B INVX1_LOC_53/A 0.14fF
C52139 NOR2X1_LOC_759/A INVX1_LOC_33/A 0.73fF
C52140 INVX1_LOC_50/A NAND2X1_LOC_858/B 0.22fF
C52141 NAND2X1_LOC_860/A INVX1_LOC_73/A 0.00fF
C52142 NOR2X1_LOC_514/A NAND2X1_LOC_141/A 0.02fF
C52143 NAND2X1_LOC_725/A INVX1_LOC_28/A 0.05fF
C52144 NOR2X1_LOC_533/Y INVX1_LOC_22/A 0.03fF
C52145 NOR2X1_LOC_790/B INVX1_LOC_75/A 0.03fF
C52146 NOR2X1_LOC_208/Y NOR2X1_LOC_562/a_36_216# 0.00fF
C52147 NOR2X1_LOC_639/B INVX1_LOC_302/Y 0.15fF
C52148 INVX1_LOC_247/A NOR2X1_LOC_334/Y 0.01fF
C52149 INVX1_LOC_208/Y NAND2X1_LOC_337/B 0.00fF
C52150 NAND2X1_LOC_198/B INVX1_LOC_8/A 0.07fF
C52151 INVX1_LOC_17/A NAND2X1_LOC_660/Y 0.00fF
C52152 NOR2X1_LOC_431/Y INVX1_LOC_63/Y 0.07fF
C52153 NAND2X1_LOC_728/Y INVX1_LOC_240/A 0.00fF
C52154 NOR2X1_LOC_88/Y INVX1_LOC_84/A 0.10fF
C52155 INVX1_LOC_72/A INVX1_LOC_177/A 0.03fF
C52156 NOR2X1_LOC_389/B INVX1_LOC_171/Y 0.01fF
C52157 INVX1_LOC_73/Y NOR2X1_LOC_561/Y 0.01fF
C52158 NOR2X1_LOC_219/B INVX1_LOC_77/A 0.02fF
C52159 NOR2X1_LOC_778/B INVX1_LOC_30/A 0.06fF
C52160 INVX1_LOC_35/A INVX1_LOC_86/A 0.00fF
C52161 INVX1_LOC_64/A INPUT_0 0.92fF
C52162 NAND2X1_LOC_796/B NAND2X1_LOC_807/Y 0.04fF
C52163 NOR2X1_LOC_372/A INVX1_LOC_16/A 0.11fF
C52164 NAND2X1_LOC_711/B INVX1_LOC_240/A 0.16fF
C52165 NOR2X1_LOC_274/Y INVX1_LOC_225/A 0.02fF
C52166 INVX1_LOC_58/A NOR2X1_LOC_528/Y 0.12fF
C52167 INVX1_LOC_280/Y INVX1_LOC_72/A 0.03fF
C52168 INVX1_LOC_98/A INVX1_LOC_23/A 0.00fF
C52169 NOR2X1_LOC_33/A NAND2X1_LOC_555/Y 0.04fF
C52170 INVX1_LOC_17/A D_INPUT_0 1.75fF
C52171 NAND2X1_LOC_99/a_36_24# NAND2X1_LOC_276/Y 0.01fF
C52172 INVX1_LOC_127/Y NOR2X1_LOC_271/Y 0.03fF
C52173 NOR2X1_LOC_647/A INVX1_LOC_59/Y 0.00fF
C52174 NOR2X1_LOC_78/A INVX1_LOC_23/A 0.14fF
C52175 INVX1_LOC_36/A INVX1_LOC_232/A 0.07fF
C52176 INVX1_LOC_32/A INVX1_LOC_38/A 1.56fF
C52177 NOR2X1_LOC_436/a_36_216# INPUT_0 0.02fF
C52178 INVX1_LOC_63/Y NOR2X1_LOC_364/Y -0.01fF
C52179 NOR2X1_LOC_155/A INVX1_LOC_109/A 0.00fF
C52180 NOR2X1_LOC_269/Y INVX1_LOC_53/A 0.07fF
C52181 D_INPUT_1 NOR2X1_LOC_405/A 0.10fF
C52182 INVX1_LOC_15/Y NOR2X1_LOC_617/Y 0.53fF
C52183 NAND2X1_LOC_363/B NOR2X1_LOC_557/A 0.07fF
C52184 NAND2X1_LOC_579/A INVX1_LOC_140/A 0.10fF
C52185 NOR2X1_LOC_297/A INVX1_LOC_280/A 0.03fF
C52186 INVX1_LOC_89/A NOR2X1_LOC_745/Y 0.01fF
C52187 INVX1_LOC_225/Y INVX1_LOC_171/A 0.00fF
C52188 NOR2X1_LOC_168/B INVX1_LOC_77/A 0.07fF
C52189 INVX1_LOC_38/A NOR2X1_LOC_329/Y 0.50fF
C52190 NOR2X1_LOC_590/A NOR2X1_LOC_717/B 0.03fF
C52191 NOR2X1_LOC_48/B INVX1_LOC_291/A 0.13fF
C52192 INVX1_LOC_141/Y NAND2X1_LOC_796/Y 0.02fF
C52193 NAND2X1_LOC_555/Y D_INPUT_0 0.02fF
C52194 INVX1_LOC_300/Y NAND2X1_LOC_853/Y 0.45fF
C52195 INVX1_LOC_116/A NOR2X1_LOC_220/A 0.21fF
C52196 INVX1_LOC_12/A INVX1_LOC_260/Y 0.03fF
C52197 VDD NAND2X1_LOC_402/B 0.01fF
C52198 NOR2X1_LOC_48/B NAND2X1_LOC_802/Y 0.65fF
C52199 NOR2X1_LOC_400/B VDD -0.00fF
C52200 NOR2X1_LOC_91/A NOR2X1_LOC_176/a_36_216# 0.01fF
C52201 INVX1_LOC_208/A NOR2X1_LOC_759/Y 0.00fF
C52202 NOR2X1_LOC_553/B NOR2X1_LOC_703/B 0.00fF
C52203 NOR2X1_LOC_433/a_36_216# INVX1_LOC_266/Y 0.01fF
C52204 NOR2X1_LOC_844/Y NOR2X1_LOC_99/B 0.04fF
C52205 INVX1_LOC_224/Y VDD 1.66fF
C52206 NAND2X1_LOC_734/B NAND2X1_LOC_357/B 0.04fF
C52207 INVX1_LOC_24/A NAND2X1_LOC_479/Y 0.03fF
C52208 INVX1_LOC_299/A NOR2X1_LOC_74/A 0.07fF
C52209 NOR2X1_LOC_78/B NOR2X1_LOC_717/a_36_216# 0.01fF
C52210 INVX1_LOC_38/A NAND2X1_LOC_175/Y 0.12fF
C52211 NOR2X1_LOC_178/Y NAND2X1_LOC_642/Y 0.09fF
C52212 NOR2X1_LOC_598/B NOR2X1_LOC_35/Y 0.19fF
C52213 INVX1_LOC_304/Y NOR2X1_LOC_369/a_36_216# 0.00fF
C52214 NOR2X1_LOC_75/Y NOR2X1_LOC_741/a_36_216# 0.00fF
C52215 NOR2X1_LOC_216/B INVX1_LOC_3/Y 0.07fF
C52216 NOR2X1_LOC_13/Y NAND2X1_LOC_662/Y 0.04fF
C52217 D_GATE_741 INVX1_LOC_75/A 0.02fF
C52218 INVX1_LOC_36/Y NOR2X1_LOC_247/Y 0.07fF
C52219 NOR2X1_LOC_405/A NOR2X1_LOC_108/a_36_216# 0.00fF
C52220 INVX1_LOC_28/A NOR2X1_LOC_372/A 0.11fF
C52221 INVX1_LOC_227/A NOR2X1_LOC_609/A 0.05fF
C52222 NOR2X1_LOC_488/Y NOR2X1_LOC_716/B 0.19fF
C52223 NOR2X1_LOC_405/A NOR2X1_LOC_652/Y 0.01fF
C52224 INVX1_LOC_57/A NOR2X1_LOC_107/a_36_216# 0.00fF
C52225 NOR2X1_LOC_716/B NOR2X1_LOC_82/Y 0.05fF
C52226 VDD NAND2X1_LOC_793/B 0.71fF
C52227 NOR2X1_LOC_802/A INVX1_LOC_196/A 0.10fF
C52228 NOR2X1_LOC_538/B NOR2X1_LOC_9/Y 0.03fF
C52229 INPUT_3 NAND2X1_LOC_348/A 0.03fF
C52230 NOR2X1_LOC_554/B NOR2X1_LOC_846/B 0.02fF
C52231 NOR2X1_LOC_739/Y NOR2X1_LOC_728/B 0.01fF
C52232 INVX1_LOC_23/A NOR2X1_LOC_60/Y 0.15fF
C52233 NOR2X1_LOC_334/Y NOR2X1_LOC_862/B 0.02fF
C52234 NAND2X1_LOC_36/A NOR2X1_LOC_163/a_36_216# 0.00fF
C52235 NOR2X1_LOC_590/A NOR2X1_LOC_151/Y 0.07fF
C52236 INVX1_LOC_135/A INVX1_LOC_24/A 0.06fF
C52237 INVX1_LOC_246/A INVX1_LOC_144/A 0.02fF
C52238 INVX1_LOC_13/A INVX1_LOC_33/A 0.19fF
C52239 INVX1_LOC_225/Y INVX1_LOC_222/A 0.02fF
C52240 INVX1_LOC_43/Y INPUT_0 0.03fF
C52241 NOR2X1_LOC_619/A INVX1_LOC_8/A 0.08fF
C52242 NOR2X1_LOC_822/Y NAND2X1_LOC_839/A 0.09fF
C52243 INVX1_LOC_84/A INVX1_LOC_15/A 0.13fF
C52244 NAND2X1_LOC_81/B INVX1_LOC_284/A 0.02fF
C52245 INVX1_LOC_77/A NAND2X1_LOC_656/Y 0.18fF
C52246 NAND2X1_LOC_308/Y INVX1_LOC_16/A 0.03fF
C52247 NAND2X1_LOC_357/B INVX1_LOC_25/Y 0.08fF
C52248 NOR2X1_LOC_309/Y INVX1_LOC_232/A 0.06fF
C52249 INVX1_LOC_26/A INVX1_LOC_92/A 0.10fF
C52250 NOR2X1_LOC_770/A INVX1_LOC_83/A 0.01fF
C52251 NOR2X1_LOC_287/A NOR2X1_LOC_802/A 0.04fF
C52252 NAND2X1_LOC_231/Y NAND2X1_LOC_850/Y 0.02fF
C52253 NOR2X1_LOC_541/Y NOR2X1_LOC_337/Y 0.02fF
C52254 NAND2X1_LOC_537/Y NAND2X1_LOC_729/B 0.00fF
C52255 NOR2X1_LOC_160/B NOR2X1_LOC_334/A 6.48fF
C52256 NAND2X1_LOC_93/B NOR2X1_LOC_72/Y -0.02fF
C52257 NOR2X1_LOC_690/Y INVX1_LOC_240/A 0.03fF
C52258 NOR2X1_LOC_68/A NOR2X1_LOC_322/Y 0.15fF
C52259 NAND2X1_LOC_651/B INVX1_LOC_15/A 0.05fF
C52260 NOR2X1_LOC_589/A INVX1_LOC_266/Y 0.08fF
C52261 INVX1_LOC_223/A NOR2X1_LOC_337/A 0.27fF
C52262 NOR2X1_LOC_191/B INVX1_LOC_102/Y 0.05fF
C52263 INVX1_LOC_229/Y NOR2X1_LOC_821/Y 0.05fF
C52264 NOR2X1_LOC_178/Y NOR2X1_LOC_271/Y 0.02fF
C52265 INVX1_LOC_163/A D_GATE_662 0.01fF
C52266 NOR2X1_LOC_554/A NOR2X1_LOC_847/B 0.03fF
C52267 INVX1_LOC_55/Y INVX1_LOC_33/A 0.08fF
C52268 INVX1_LOC_124/A NAND2X1_LOC_656/Y 0.01fF
C52269 NOR2X1_LOC_392/Y NOR2X1_LOC_78/a_36_216# 0.01fF
C52270 INVX1_LOC_153/Y INVX1_LOC_313/Y 0.00fF
C52271 INVX1_LOC_31/A NOR2X1_LOC_78/A 0.30fF
C52272 NAND2X1_LOC_513/B INVX1_LOC_117/A 0.01fF
C52273 NOR2X1_LOC_91/Y NOR2X1_LOC_167/Y 0.01fF
C52274 INVX1_LOC_23/Y INVX1_LOC_63/A 0.07fF
C52275 NOR2X1_LOC_385/Y NOR2X1_LOC_577/Y 0.44fF
C52276 INVX1_LOC_13/A INVX1_LOC_40/A 0.42fF
C52277 INVX1_LOC_30/A NOR2X1_LOC_557/A 0.02fF
C52278 NOR2X1_LOC_706/A NOR2X1_LOC_550/B 0.70fF
C52279 INVX1_LOC_25/A NAND2X1_LOC_574/A 0.04fF
C52280 INVX1_LOC_83/A NAND2X1_LOC_451/Y 0.12fF
C52281 INVX1_LOC_135/A INVX1_LOC_143/A 0.29fF
C52282 NOR2X1_LOC_785/Y NAND2X1_LOC_323/B 0.02fF
C52283 NOR2X1_LOC_103/Y VDD -0.00fF
C52284 INVX1_LOC_278/A NOR2X1_LOC_88/Y 0.07fF
C52285 NAND2X1_LOC_308/Y INVX1_LOC_28/A 0.02fF
C52286 NAND2X1_LOC_74/B NOR2X1_LOC_89/Y 0.10fF
C52287 INVX1_LOC_271/A NAND2X1_LOC_475/Y 0.10fF
C52288 NOR2X1_LOC_510/Y NOR2X1_LOC_506/Y 0.05fF
C52289 INVX1_LOC_212/Y INVX1_LOC_75/A 0.07fF
C52290 INVX1_LOC_75/A NOR2X1_LOC_344/A 0.02fF
C52291 INVX1_LOC_313/Y INVX1_LOC_177/A 1.17fF
C52292 NOR2X1_LOC_541/Y VDD 0.25fF
C52293 INVX1_LOC_30/A NOR2X1_LOC_657/B 0.01fF
C52294 INVX1_LOC_17/A NOR2X1_LOC_859/Y 0.01fF
C52295 NAND2X1_LOC_778/Y INVX1_LOC_185/A 0.12fF
C52296 NOR2X1_LOC_655/B NAND2X1_LOC_492/a_36_24# 0.07fF
C52297 NOR2X1_LOC_261/Y INVX1_LOC_84/A 0.07fF
C52298 INVX1_LOC_45/A NOR2X1_LOC_56/Y 0.07fF
C52299 INVX1_LOC_34/A INVX1_LOC_282/A 0.17fF
C52300 NOR2X1_LOC_590/A NOR2X1_LOC_567/a_36_216# 0.00fF
C52301 NOR2X1_LOC_89/A NOR2X1_LOC_278/Y 0.04fF
C52302 NOR2X1_LOC_337/Y INVX1_LOC_71/A 0.00fF
C52303 INVX1_LOC_41/A NOR2X1_LOC_188/A 0.09fF
C52304 INVX1_LOC_77/A INVX1_LOC_78/Y 0.04fF
C52305 INVX1_LOC_278/A INVX1_LOC_84/A 0.10fF
C52306 INVX1_LOC_17/A NAND2X1_LOC_848/A 0.10fF
C52307 INVX1_LOC_41/A NOR2X1_LOC_548/B 0.03fF
C52308 NOR2X1_LOC_791/B INVX1_LOC_95/Y 0.12fF
C52309 NOR2X1_LOC_276/Y INVX1_LOC_12/Y 0.00fF
C52310 INVX1_LOC_24/A NOR2X1_LOC_552/A 0.07fF
C52311 INVX1_LOC_32/A NAND2X1_LOC_223/A 0.07fF
C52312 NAND2X1_LOC_717/Y NAND2X1_LOC_560/A 0.01fF
C52313 NOR2X1_LOC_15/Y INVX1_LOC_185/A 0.06fF
C52314 INVX1_LOC_45/A VDD 2.37fF
C52315 INVX1_LOC_47/Y INVX1_LOC_87/A 0.09fF
C52316 INVX1_LOC_30/Y NOR2X1_LOC_749/a_36_216# 0.00fF
C52317 INVX1_LOC_12/A NAND2X1_LOC_201/a_36_24# 0.00fF
C52318 NOR2X1_LOC_568/A VDD 0.98fF
C52319 INVX1_LOC_21/A NOR2X1_LOC_841/A 0.03fF
C52320 NAND2X1_LOC_564/B INVX1_LOC_90/A 0.00fF
C52321 NOR2X1_LOC_804/B INVX1_LOC_186/A 0.07fF
C52322 NAND2X1_LOC_856/A VDD 0.04fF
C52323 NAND2X1_LOC_785/B NAND2X1_LOC_804/Y 0.18fF
C52324 NOR2X1_LOC_250/A NAND2X1_LOC_760/a_36_24# 0.00fF
C52325 INVX1_LOC_291/Y NOR2X1_LOC_152/Y 0.03fF
C52326 NOR2X1_LOC_315/Y NOR2X1_LOC_9/Y 0.09fF
C52327 INVX1_LOC_64/A NOR2X1_LOC_84/B -0.00fF
C52328 NOR2X1_LOC_360/Y INVX1_LOC_46/A 0.10fF
C52329 INVX1_LOC_135/A NOR2X1_LOC_130/A 0.06fF
C52330 INVX1_LOC_136/A INVX1_LOC_12/Y 0.01fF
C52331 INPUT_0 NAND2X1_LOC_850/Y 0.47fF
C52332 NOR2X1_LOC_360/Y NOR2X1_LOC_98/A 0.07fF
C52333 NAND2X1_LOC_560/A INVX1_LOC_16/A 0.02fF
C52334 NOR2X1_LOC_343/B NOR2X1_LOC_814/A 0.04fF
C52335 NOR2X1_LOC_273/Y NAND2X1_LOC_211/Y 0.14fF
C52336 NOR2X1_LOC_846/A INVX1_LOC_63/A 0.01fF
C52337 INVX1_LOC_17/A INVX1_LOC_46/Y 0.00fF
C52338 NOR2X1_LOC_759/Y NAND2X1_LOC_211/Y 0.03fF
C52339 INVX1_LOC_215/A NOR2X1_LOC_135/Y 0.12fF
C52340 INVX1_LOC_202/A NAND2X1_LOC_211/Y 0.07fF
C52341 INVX1_LOC_290/Y NOR2X1_LOC_717/A 0.07fF
C52342 INVX1_LOC_233/Y INVX1_LOC_284/A 0.30fF
C52343 INVX1_LOC_1/A NAND2X1_LOC_574/A 0.01fF
C52344 INVX1_LOC_14/A NAND2X1_LOC_141/Y 0.06fF
C52345 NOR2X1_LOC_643/Y INVX1_LOC_20/A 0.00fF
C52346 INVX1_LOC_24/A INVX1_LOC_139/Y 0.01fF
C52347 INVX1_LOC_71/A VDD 4.71fF
C52348 NAND2X1_LOC_715/B INVX1_LOC_109/A 0.02fF
C52349 INVX1_LOC_57/A NOR2X1_LOC_620/a_36_216# 0.00fF
C52350 NOR2X1_LOC_188/A NOR2X1_LOC_211/A 0.03fF
C52351 NOR2X1_LOC_381/Y NOR2X1_LOC_649/B 0.02fF
C52352 NOR2X1_LOC_294/Y INVX1_LOC_9/A 0.29fF
C52353 NOR2X1_LOC_238/Y INVX1_LOC_37/Y 0.00fF
C52354 INVX1_LOC_100/A INVX1_LOC_56/Y 0.04fF
C52355 NOR2X1_LOC_381/Y INVX1_LOC_3/A 0.05fF
C52356 INVX1_LOC_24/A NOR2X1_LOC_813/Y 0.09fF
C52357 NOR2X1_LOC_548/B NOR2X1_LOC_211/A 0.05fF
C52358 NOR2X1_LOC_554/A NOR2X1_LOC_660/Y 0.00fF
C52359 NOR2X1_LOC_441/Y INVX1_LOC_291/A 0.02fF
C52360 NOR2X1_LOC_500/A INVX1_LOC_117/A 0.09fF
C52361 NOR2X1_LOC_653/B NAND2X1_LOC_74/B 0.02fF
C52362 NOR2X1_LOC_442/a_36_216# NOR2X1_LOC_814/A 0.01fF
C52363 INVX1_LOC_108/Y INVX1_LOC_15/A 0.98fF
C52364 INVX1_LOC_83/A NOR2X1_LOC_567/B 0.09fF
C52365 NAND2X1_LOC_374/Y INVX1_LOC_91/A 0.09fF
C52366 NAND2X1_LOC_811/Y INVX1_LOC_20/A 0.03fF
C52367 INVX1_LOC_278/A INVX1_LOC_15/A 0.07fF
C52368 INVX1_LOC_159/A NOR2X1_LOC_331/B 0.01fF
C52369 INVX1_LOC_207/A INVX1_LOC_46/A 0.12fF
C52370 NOR2X1_LOC_78/B NOR2X1_LOC_269/Y 0.07fF
C52371 NOR2X1_LOC_128/B INVX1_LOC_75/A 1.50fF
C52372 NAND2X1_LOC_358/Y INVX1_LOC_158/Y 0.05fF
C52373 INVX1_LOC_235/Y INVX1_LOC_29/A 0.04fF
C52374 NOR2X1_LOC_738/A INVX1_LOC_85/Y 0.02fF
C52375 NOR2X1_LOC_257/a_36_216# NOR2X1_LOC_684/Y 0.00fF
C52376 NAND2X1_LOC_149/Y INVX1_LOC_29/A 0.10fF
C52377 NAND2X1_LOC_198/B INVX1_LOC_118/Y 0.03fF
C52378 NAND2X1_LOC_568/a_36_24# NAND2X1_LOC_800/A 0.00fF
C52379 NOR2X1_LOC_380/A NOR2X1_LOC_380/Y 12.96fF
C52380 NAND2X1_LOC_842/B NAND2X1_LOC_830/a_36_24# 0.02fF
C52381 NOR2X1_LOC_557/Y NOR2X1_LOC_558/a_36_216# 0.01fF
C52382 INVX1_LOC_174/Y INVX1_LOC_86/Y 0.11fF
C52383 INVX1_LOC_33/A INVX1_LOC_66/Y 0.07fF
C52384 NOR2X1_LOC_721/Y NOR2X1_LOC_749/Y 0.18fF
C52385 NAND2X1_LOC_811/Y NOR2X1_LOC_765/Y 0.79fF
C52386 NOR2X1_LOC_816/A NAND2X1_LOC_604/a_36_24# 0.01fF
C52387 NAND2X1_LOC_579/A INVX1_LOC_42/A 0.08fF
C52388 INVX1_LOC_275/A INVX1_LOC_9/A 0.02fF
C52389 NOR2X1_LOC_717/Y NOR2X1_LOC_66/Y 0.00fF
C52390 INVX1_LOC_159/A NOR2X1_LOC_592/B 0.01fF
C52391 INVX1_LOC_174/A INVX1_LOC_19/A 0.03fF
C52392 NOR2X1_LOC_74/A NOR2X1_LOC_166/Y 0.04fF
C52393 NOR2X1_LOC_437/a_36_216# INVX1_LOC_92/A 0.00fF
C52394 NOR2X1_LOC_6/B NOR2X1_LOC_536/A 0.28fF
C52395 INVX1_LOC_313/Y INVX1_LOC_285/Y 0.02fF
C52396 INVX1_LOC_302/A INVX1_LOC_302/Y 0.09fF
C52397 NOR2X1_LOC_742/A NOR2X1_LOC_303/a_36_216# 0.01fF
C52398 NOR2X1_LOC_160/B NAND2X1_LOC_74/B 0.22fF
C52399 NOR2X1_LOC_372/Y INVX1_LOC_203/A 0.01fF
C52400 INVX1_LOC_230/Y INVX1_LOC_12/A 0.07fF
C52401 INVX1_LOC_313/A NOR2X1_LOC_78/A 0.07fF
C52402 INVX1_LOC_120/A NAND2X1_LOC_86/Y 0.01fF
C52403 INVX1_LOC_45/A INVX1_LOC_133/A 0.21fF
C52404 INVX1_LOC_35/A INVX1_LOC_57/A 0.16fF
C52405 NOR2X1_LOC_6/B NOR2X1_LOC_655/Y 0.27fF
C52406 INVX1_LOC_306/Y NAND2X1_LOC_99/A 0.17fF
C52407 INVX1_LOC_269/A NAND2X1_LOC_647/B 0.02fF
C52408 NOR2X1_LOC_400/A INVX1_LOC_166/A 0.01fF
C52409 NOR2X1_LOC_87/Y INVX1_LOC_230/A 0.01fF
C52410 NOR2X1_LOC_748/Y INVX1_LOC_37/A 0.03fF
C52411 NOR2X1_LOC_91/A NOR2X1_LOC_186/Y 0.10fF
C52412 NOR2X1_LOC_387/A NAND2X1_LOC_463/B 0.02fF
C52413 INVX1_LOC_313/Y INVX1_LOC_65/A 0.25fF
C52414 NOR2X1_LOC_6/B NAND2X1_LOC_93/B 0.00fF
C52415 NAND2X1_LOC_579/A INVX1_LOC_78/A 0.01fF
C52416 INVX1_LOC_298/Y NAND2X1_LOC_149/Y 0.02fF
C52417 NAND2X1_LOC_565/B NOR2X1_LOC_813/Y 0.01fF
C52418 NAND2X1_LOC_549/Y NOR2X1_LOC_392/Y 0.01fF
C52419 INVX1_LOC_49/A NOR2X1_LOC_450/B 0.03fF
C52420 NAND2X1_LOC_309/a_36_24# NOR2X1_LOC_188/A 0.01fF
C52421 INVX1_LOC_313/Y NOR2X1_LOC_137/B 0.09fF
C52422 INVX1_LOC_225/Y INVX1_LOC_4/A 0.20fF
C52423 NOR2X1_LOC_91/A NAND2X1_LOC_573/Y 0.10fF
C52424 INVX1_LOC_9/Y INVX1_LOC_38/A 0.02fF
C52425 INVX1_LOC_58/A INVX1_LOC_93/A 0.07fF
C52426 INVX1_LOC_269/A NOR2X1_LOC_395/Y 0.01fF
C52427 NOR2X1_LOC_250/Y INVX1_LOC_94/Y 0.48fF
C52428 NOR2X1_LOC_186/Y INVX1_LOC_23/A 0.08fF
C52429 INVX1_LOC_17/Y NOR2X1_LOC_496/Y 0.14fF
C52430 GATE_741 NAND2X1_LOC_725/Y 0.03fF
C52431 NOR2X1_LOC_32/B INVX1_LOC_5/A 0.67fF
C52432 NAND2X1_LOC_729/B NAND2X1_LOC_855/Y 0.04fF
C52433 NOR2X1_LOC_294/Y NOR2X1_LOC_861/Y 0.02fF
C52434 INVX1_LOC_30/Y NOR2X1_LOC_536/A 0.04fF
C52435 NOR2X1_LOC_67/A NAND2X1_LOC_243/Y 0.02fF
C52436 INVX1_LOC_53/Y INVX1_LOC_118/Y 0.03fF
C52437 NAND2X1_LOC_844/a_36_24# INVX1_LOC_91/A 0.00fF
C52438 INVX1_LOC_204/A NAND2X1_LOC_149/Y 0.05fF
C52439 NAND2X1_LOC_30/Y NOR2X1_LOC_30/Y 0.10fF
C52440 NOR2X1_LOC_489/B NOR2X1_LOC_772/B 0.02fF
C52441 NOR2X1_LOC_67/A INVX1_LOC_89/Y 0.02fF
C52442 NOR2X1_LOC_333/A INVX1_LOC_37/A 0.02fF
C52443 NOR2X1_LOC_91/A NAND2X1_LOC_724/A 0.50fF
C52444 NOR2X1_LOC_749/Y VDD 0.37fF
C52445 INVX1_LOC_11/A NOR2X1_LOC_278/Y 0.05fF
C52446 NOR2X1_LOC_6/B NOR2X1_LOC_649/B 0.11fF
C52447 NOR2X1_LOC_789/A INVX1_LOC_9/A 0.00fF
C52448 NOR2X1_LOC_6/B INVX1_LOC_3/A 0.19fF
C52449 NOR2X1_LOC_813/Y NOR2X1_LOC_130/A 0.07fF
C52450 INVX1_LOC_98/A INVX1_LOC_6/A 1.04fF
C52451 NAND2X1_LOC_861/Y NOR2X1_LOC_176/Y 0.01fF
C52452 INPUT_3 NAND2X1_LOC_223/A 0.07fF
C52453 INVX1_LOC_193/Y NOR2X1_LOC_725/A 0.01fF
C52454 INVX1_LOC_101/Y NOR2X1_LOC_383/B 0.00fF
C52455 D_GATE_366 INVX1_LOC_37/A 0.03fF
C52456 NOR2X1_LOC_32/B INVX1_LOC_178/A 0.10fF
C52457 NAND2X1_LOC_662/B NOR2X1_LOC_43/Y 0.05fF
C52458 NOR2X1_LOC_667/Y INVX1_LOC_273/A 0.19fF
C52459 INVX1_LOC_90/A NAND2X1_LOC_804/Y 0.03fF
C52460 INVX1_LOC_50/A NAND2X1_LOC_190/Y 0.01fF
C52461 NAND2X1_LOC_348/A NOR2X1_LOC_332/B -0.02fF
C52462 NOR2X1_LOC_78/A INVX1_LOC_6/A 0.18fF
C52463 NAND2X1_LOC_363/B INVX1_LOC_27/A 0.11fF
C52464 INVX1_LOC_72/A NAND2X1_LOC_269/a_36_24# 0.01fF
C52465 NAND2X1_LOC_794/B NAND2X1_LOC_725/A 0.10fF
C52466 INVX1_LOC_224/Y NOR2X1_LOC_361/B 0.10fF
C52467 INVX1_LOC_230/Y NOR2X1_LOC_29/a_36_216# 0.00fF
C52468 NOR2X1_LOC_419/Y NOR2X1_LOC_67/Y 0.02fF
C52469 NOR2X1_LOC_761/a_36_216# NOR2X1_LOC_409/B 0.00fF
C52470 INVX1_LOC_248/A NOR2X1_LOC_841/A 0.23fF
C52471 NAND2X1_LOC_656/Y INVX1_LOC_9/A 0.08fF
C52472 NOR2X1_LOC_130/A INVX1_LOC_280/A 0.15fF
C52473 NAND2X1_LOC_796/B NOR2X1_LOC_109/Y 0.11fF
C52474 INVX1_LOC_102/Y VDD 1.06fF
C52475 NOR2X1_LOC_798/A NOR2X1_LOC_212/a_36_216# 0.00fF
C52476 INVX1_LOC_30/Y NAND2X1_LOC_93/B 0.10fF
C52477 INVX1_LOC_22/A NOR2X1_LOC_831/B 0.41fF
C52478 INVX1_LOC_290/A NOR2X1_LOC_155/A 0.08fF
C52479 NOR2X1_LOC_606/a_36_216# INVX1_LOC_23/Y 0.01fF
C52480 NOR2X1_LOC_590/A NOR2X1_LOC_39/a_36_216# 0.00fF
C52481 NAND2X1_LOC_186/a_36_24# NOR2X1_LOC_331/B 0.04fF
C52482 NOR2X1_LOC_810/A NOR2X1_LOC_809/B 0.01fF
C52483 NAND2X1_LOC_374/Y INVX1_LOC_203/A 0.13fF
C52484 INVX1_LOC_232/A NAND2X1_LOC_609/a_36_24# 0.00fF
C52485 INVX1_LOC_90/A NOR2X1_LOC_261/A 0.02fF
C52486 NOR2X1_LOC_71/Y NAND2X1_LOC_268/a_36_24# 0.01fF
C52487 INVX1_LOC_27/A NOR2X1_LOC_791/Y 0.01fF
C52488 NAND2X1_LOC_757/a_36_24# NOR2X1_LOC_38/B 0.00fF
C52489 INVX1_LOC_50/A NOR2X1_LOC_389/A 0.01fF
C52490 NOR2X1_LOC_68/A NOR2X1_LOC_685/a_36_216# 0.00fF
C52491 INVX1_LOC_6/A NAND2X1_LOC_464/A 0.01fF
C52492 NOR2X1_LOC_91/A INVX1_LOC_170/A 0.05fF
C52493 NOR2X1_LOC_457/B NAND2X1_LOC_454/Y 0.09fF
C52494 NOR2X1_LOC_772/B INVX1_LOC_14/A 0.07fF
C52495 NOR2X1_LOC_45/Y INVX1_LOC_23/A 0.28fF
C52496 NOR2X1_LOC_192/A INVX1_LOC_95/Y 0.01fF
C52497 NAND2X1_LOC_622/B INVX1_LOC_194/Y 0.02fF
C52498 NAND2X1_LOC_21/Y INVX1_LOC_15/A 0.13fF
C52499 INVX1_LOC_33/A INVX1_LOC_32/A 2.69fF
C52500 NAND2X1_LOC_338/B NAND2X1_LOC_81/B 0.02fF
C52501 INVX1_LOC_232/A INVX1_LOC_63/A 0.35fF
C52502 INVX1_LOC_125/Y INVX1_LOC_20/A 0.01fF
C52503 INVX1_LOC_69/Y NOR2X1_LOC_168/a_36_216# 0.01fF
C52504 INVX1_LOC_196/Y NOR2X1_LOC_801/a_36_216# 0.00fF
C52505 INVX1_LOC_13/Y INVX1_LOC_14/A 0.58fF
C52506 NAND2X1_LOC_41/Y NOR2X1_LOC_814/A 0.01fF
C52507 NOR2X1_LOC_84/A INVX1_LOC_3/Y 0.08fF
C52508 INVX1_LOC_30/A INVX1_LOC_271/A 0.16fF
C52509 NOR2X1_LOC_160/B NOR2X1_LOC_660/Y 0.17fF
C52510 NOR2X1_LOC_848/Y INVX1_LOC_38/Y 0.17fF
C52511 INVX1_LOC_24/A NOR2X1_LOC_541/B 0.03fF
C52512 INVX1_LOC_170/A INVX1_LOC_23/A 0.01fF
C52513 INVX1_LOC_196/Y INVX1_LOC_307/A 0.07fF
C52514 INVX1_LOC_239/A INVX1_LOC_163/A 2.05fF
C52515 INVX1_LOC_190/Y NOR2X1_LOC_592/B 0.01fF
C52516 NOR2X1_LOC_269/Y INVX1_LOC_46/A 1.78fF
C52517 INVX1_LOC_256/A INVX1_LOC_50/Y 0.07fF
C52518 NOR2X1_LOC_589/A INVX1_LOC_19/A 0.03fF
C52519 INVX1_LOC_16/A INVX1_LOC_29/A 5.02fF
C52520 NOR2X1_LOC_516/B NAND2X1_LOC_207/Y 0.01fF
C52521 NAND2X1_LOC_341/A INVX1_LOC_12/A 0.03fF
C52522 NOR2X1_LOC_486/Y NOR2X1_LOC_357/Y 0.04fF
C52523 INVX1_LOC_28/A NOR2X1_LOC_58/Y 0.02fF
C52524 INVX1_LOC_33/A NAND2X1_LOC_175/Y 0.37fF
C52525 INVX1_LOC_50/A NOR2X1_LOC_596/A 0.03fF
C52526 NOR2X1_LOC_706/A INVX1_LOC_75/Y 0.26fF
C52527 INVX1_LOC_266/Y INVX1_LOC_4/A 0.10fF
C52528 INVX1_LOC_21/A NOR2X1_LOC_705/B 0.02fF
C52529 INVX1_LOC_77/A NOR2X1_LOC_727/B 0.00fF
C52530 NOR2X1_LOC_516/B NOR2X1_LOC_847/B 0.01fF
C52531 INVX1_LOC_233/Y INVX1_LOC_72/A 0.07fF
C52532 NAND2X1_LOC_9/Y NOR2X1_LOC_360/Y 0.03fF
C52533 NOR2X1_LOC_337/Y NOR2X1_LOC_331/B 0.04fF
C52534 INVX1_LOC_28/A NAND2X1_LOC_606/a_36_24# 0.00fF
C52535 NAND2X1_LOC_363/B NAND2X1_LOC_338/a_36_24# 0.00fF
C52536 INVX1_LOC_78/Y INVX1_LOC_9/A 0.03fF
C52537 NOR2X1_LOC_91/A NAND2X1_LOC_640/Y 0.00fF
C52538 INVX1_LOC_276/A INVX1_LOC_21/Y 0.04fF
C52539 INVX1_LOC_266/A INVX1_LOC_256/A 0.67fF
C52540 NOR2X1_LOC_92/Y NAND2X1_LOC_807/A 0.03fF
C52541 INVX1_LOC_40/A INVX1_LOC_32/A 0.12fF
C52542 INVX1_LOC_171/A INVX1_LOC_19/A 0.01fF
C52543 NOR2X1_LOC_537/Y INVX1_LOC_4/Y 0.07fF
C52544 INVX1_LOC_247/A NAND2X1_LOC_472/Y 0.05fF
C52545 NOR2X1_LOC_468/a_36_216# INVX1_LOC_12/A 0.02fF
C52546 NOR2X1_LOC_361/B NOR2X1_LOC_103/Y 0.10fF
C52547 NOR2X1_LOC_52/B NOR2X1_LOC_278/Y 0.00fF
C52548 NAND2X1_LOC_338/B INVX1_LOC_4/Y 0.49fF
C52549 NOR2X1_LOC_510/Y INVX1_LOC_45/A 0.46fF
C52550 NOR2X1_LOC_8/a_36_216# NOR2X1_LOC_392/Y 0.01fF
C52551 NOR2X1_LOC_91/A INVX1_LOC_225/A 0.03fF
C52552 NAND2X1_LOC_218/B NAND2X1_LOC_46/a_36_24# 0.00fF
C52553 NOR2X1_LOC_533/Y NAND2X1_LOC_799/A 0.01fF
C52554 INVX1_LOC_221/Y NAND2X1_LOC_538/Y 0.04fF
C52555 INVX1_LOC_17/A NAND2X1_LOC_30/Y 0.10fF
C52556 INVX1_LOC_27/A INVX1_LOC_30/A 0.03fF
C52557 NOR2X1_LOC_45/B NAND2X1_LOC_637/Y 0.09fF
C52558 NOR2X1_LOC_738/A NAND2X1_LOC_782/B 0.02fF
C52559 INVX1_LOC_216/Y NOR2X1_LOC_82/A 0.01fF
C52560 NOR2X1_LOC_481/A INVX1_LOC_23/A 0.11fF
C52561 INVX1_LOC_77/A NOR2X1_LOC_717/A 0.03fF
C52562 NOR2X1_LOC_824/A INVX1_LOC_30/A 0.07fF
C52563 INVX1_LOC_83/A NOR2X1_LOC_633/a_36_216# 0.00fF
C52564 INVX1_LOC_136/A NOR2X1_LOC_653/B 0.01fF
C52565 INVX1_LOC_2/A NOR2X1_LOC_301/A 0.00fF
C52566 NOR2X1_LOC_52/B NOR2X1_LOC_638/Y 0.02fF
C52567 INVX1_LOC_51/A NOR2X1_LOC_350/A 0.01fF
C52568 NOR2X1_LOC_56/Y NOR2X1_LOC_331/B 0.07fF
C52569 NOR2X1_LOC_388/a_36_216# NOR2X1_LOC_334/Y 0.00fF
C52570 NAND2X1_LOC_84/Y NOR2X1_LOC_772/B 0.09fF
C52571 INVX1_LOC_303/A NOR2X1_LOC_489/B 0.02fF
C52572 NOR2X1_LOC_798/A NOR2X1_LOC_360/Y 0.03fF
C52573 INVX1_LOC_313/Y NOR2X1_LOC_830/Y 0.25fF
C52574 NOR2X1_LOC_513/Y INVX1_LOC_215/Y 0.02fF
C52575 NOR2X1_LOC_226/A NOR2X1_LOC_301/A 0.08fF
C52576 NOR2X1_LOC_78/B INVX1_LOC_26/A 0.03fF
C52577 INVX1_LOC_225/A INVX1_LOC_23/A 0.07fF
C52578 NOR2X1_LOC_67/A INVX1_LOC_16/Y 0.09fF
C52579 NOR2X1_LOC_189/A NAND2X1_LOC_725/A 0.06fF
C52580 INVX1_LOC_28/A INVX1_LOC_29/A 0.14fF
C52581 NOR2X1_LOC_71/Y NAND2X1_LOC_445/a_36_24# 0.00fF
C52582 NOR2X1_LOC_160/B NOR2X1_LOC_307/A 0.03fF
C52583 NAND2X1_LOC_850/Y INVX1_LOC_183/A 0.04fF
C52584 INVX1_LOC_11/A INVX1_LOC_236/Y 0.00fF
C52585 NAND2X1_LOC_84/Y INVX1_LOC_13/Y 0.12fF
C52586 INVX1_LOC_209/Y NOR2X1_LOC_53/Y 0.02fF
C52587 NAND2X1_LOC_725/A INVX1_LOC_231/Y 0.03fF
C52588 INVX1_LOC_45/A NOR2X1_LOC_361/B 0.08fF
C52589 NOR2X1_LOC_479/B INVX1_LOC_175/A 0.29fF
C52590 INVX1_LOC_146/Y NOR2X1_LOC_331/B 0.01fF
C52591 NOR2X1_LOC_160/B NOR2X1_LOC_276/Y 0.03fF
C52592 NOR2X1_LOC_91/A NAND2X1_LOC_852/Y 0.05fF
C52593 VDD NOR2X1_LOC_331/B 0.12fF
C52594 NAND2X1_LOC_660/Y INVX1_LOC_94/Y 0.06fF
C52595 NOR2X1_LOC_734/a_36_216# NOR2X1_LOC_814/A 0.01fF
C52596 INVX1_LOC_34/A NAND2X1_LOC_624/B 0.02fF
C52597 NOR2X1_LOC_32/B NAND2X1_LOC_562/B 1.46fF
C52598 NOR2X1_LOC_552/A NOR2X1_LOC_197/B 0.10fF
C52599 INVX1_LOC_64/A NAND2X1_LOC_811/Y 0.03fF
C52600 INVX1_LOC_104/A INVX1_LOC_58/Y 0.07fF
C52601 INVX1_LOC_298/Y INVX1_LOC_16/A 0.03fF
C52602 INVX1_LOC_58/A INVX1_LOC_54/Y 0.48fF
C52603 INVX1_LOC_123/A INVX1_LOC_84/A 0.07fF
C52604 NOR2X1_LOC_209/Y INVX1_LOC_23/A 0.10fF
C52605 INVX1_LOC_38/A NAND2X1_LOC_804/Y 0.01fF
C52606 INVX1_LOC_222/A INVX1_LOC_19/A 0.70fF
C52607 INVX1_LOC_50/A NOR2X1_LOC_220/A 0.08fF
C52608 NOR2X1_LOC_67/A NAND2X1_LOC_205/A 0.10fF
C52609 INVX1_LOC_256/A NOR2X1_LOC_248/Y 0.03fF
C52610 INVX1_LOC_124/A NOR2X1_LOC_717/A 0.37fF
C52611 INVX1_LOC_5/A NOR2X1_LOC_364/Y 0.02fF
C52612 NAND2X1_LOC_39/Y INVX1_LOC_54/A 0.01fF
C52613 NAND2X1_LOC_51/B INPUT_7 0.20fF
C52614 INVX1_LOC_37/A NAND2X1_LOC_617/a_36_24# 0.01fF
C52615 NOR2X1_LOC_65/B INVX1_LOC_208/Y 0.00fF
C52616 NOR2X1_LOC_56/Y NOR2X1_LOC_592/B 0.02fF
C52617 INVX1_LOC_305/Y INVX1_LOC_57/A 0.05fF
C52618 NOR2X1_LOC_139/Y NOR2X1_LOC_127/Y 0.07fF
C52619 D_INPUT_0 INVX1_LOC_94/Y 1.10fF
C52620 NOR2X1_LOC_720/B INVX1_LOC_5/A 0.02fF
C52621 INVX1_LOC_64/A INVX1_LOC_266/Y 0.01fF
C52622 NAND2X1_LOC_392/Y INVX1_LOC_26/A 0.05fF
C52623 INVX1_LOC_136/A NAND2X1_LOC_550/A 0.07fF
C52624 NOR2X1_LOC_292/Y INVX1_LOC_12/A 0.03fF
C52625 NOR2X1_LOC_637/A INVX1_LOC_103/A 0.03fF
C52626 NOR2X1_LOC_454/Y NOR2X1_LOC_782/a_36_216# 0.01fF
C52627 INVX1_LOC_36/A NOR2X1_LOC_225/a_36_216# 0.00fF
C52628 NAND2X1_LOC_537/Y NAND2X1_LOC_306/a_36_24# 0.01fF
C52629 INVX1_LOC_203/Y INVX1_LOC_239/A 0.03fF
C52630 NAND2X1_LOC_860/A NAND2X1_LOC_181/Y 0.04fF
C52631 NOR2X1_LOC_772/B NOR2X1_LOC_612/B 0.00fF
C52632 INVX1_LOC_136/A NOR2X1_LOC_160/B 0.13fF
C52633 INVX1_LOC_21/A NOR2X1_LOC_147/B 0.02fF
C52634 NOR2X1_LOC_361/B INVX1_LOC_71/A 0.10fF
C52635 INVX1_LOC_89/A NOR2X1_LOC_158/Y 0.07fF
C52636 INVX1_LOC_237/Y INVX1_LOC_239/A -0.01fF
C52637 INVX1_LOC_201/Y NAND2X1_LOC_141/a_36_24# 0.01fF
C52638 INVX1_LOC_103/A NOR2X1_LOC_449/a_36_216# 0.01fF
C52639 NOR2X1_LOC_45/B NAND2X1_LOC_773/B 0.03fF
C52640 NOR2X1_LOC_124/A INVX1_LOC_3/A 0.03fF
C52641 INVX1_LOC_50/A NOR2X1_LOC_548/Y 0.98fF
C52642 VDD NOR2X1_LOC_491/Y 0.12fF
C52643 INVX1_LOC_230/Y INVX1_LOC_217/A 0.00fF
C52644 INVX1_LOC_21/A NOR2X1_LOC_392/B 0.01fF
C52645 NOR2X1_LOC_689/A NOR2X1_LOC_298/Y 0.09fF
C52646 NAND2X1_LOC_363/B NAND2X1_LOC_200/B 0.03fF
C52647 VDD NOR2X1_LOC_592/B 0.42fF
C52648 NOR2X1_LOC_188/Y INVX1_LOC_57/A 0.01fF
C52649 INVX1_LOC_166/A NAND2X1_LOC_377/Y 0.04fF
C52650 INVX1_LOC_315/Y NAND2X1_LOC_207/Y 0.01fF
C52651 NAND2X1_LOC_827/a_36_24# NAND2X1_LOC_859/B -0.02fF
C52652 NAND2X1_LOC_549/Y INVX1_LOC_25/Y 0.01fF
C52653 INVX1_LOC_190/Y NOR2X1_LOC_449/A 0.06fF
C52654 NOR2X1_LOC_607/A INVX1_LOC_292/A 0.00fF
C52655 INVX1_LOC_17/A INVX1_LOC_49/A 0.08fF
C52656 D_INPUT_0 INVX1_LOC_181/A 0.08fF
C52657 NOR2X1_LOC_78/A NOR2X1_LOC_633/A 0.03fF
C52658 NAND2X1_LOC_447/Y INVX1_LOC_63/A 0.00fF
C52659 NOR2X1_LOC_516/B NOR2X1_LOC_660/Y 0.03fF
C52660 NOR2X1_LOC_653/Y INVX1_LOC_20/A 0.37fF
C52661 INVX1_LOC_42/Y INVX1_LOC_4/A 0.04fF
C52662 NOR2X1_LOC_679/a_36_216# NOR2X1_LOC_433/A 0.00fF
C52663 INVX1_LOC_305/A NOR2X1_LOC_336/B 0.04fF
C52664 NAND2X1_LOC_725/Y NOR2X1_LOC_299/Y 2.90fF
C52665 NAND2X1_LOC_738/B NOR2X1_LOC_298/Y 1.03fF
C52666 D_INPUT_3 NOR2X1_LOC_673/A 0.43fF
C52667 NOR2X1_LOC_798/A NOR2X1_LOC_539/a_36_216# 0.00fF
C52668 NOR2X1_LOC_471/Y INVX1_LOC_49/A 0.05fF
C52669 INVX1_LOC_89/A NOR2X1_LOC_646/B 0.01fF
C52670 INVX1_LOC_73/A NAND2X1_LOC_454/Y 0.01fF
C52671 INVX1_LOC_25/Y NOR2X1_LOC_291/Y 0.02fF
C52672 INVX1_LOC_20/A INVX1_LOC_19/A 0.03fF
C52673 INVX1_LOC_105/A NAND2X1_LOC_199/B 0.09fF
C52674 INVX1_LOC_132/A INVX1_LOC_31/A 0.08fF
C52675 NOR2X1_LOC_360/A INVX1_LOC_19/A 0.01fF
C52676 INVX1_LOC_45/A INVX1_LOC_184/Y 0.05fF
C52677 NOR2X1_LOC_35/Y INVX1_LOC_29/A 0.06fF
C52678 NOR2X1_LOC_658/Y INVX1_LOC_77/A 0.07fF
C52679 INVX1_LOC_46/A NOR2X1_LOC_36/B 0.03fF
C52680 INVX1_LOC_256/A NOR2X1_LOC_6/B -0.01fF
C52681 INVX1_LOC_125/Y INVX1_LOC_4/A 0.15fF
C52682 NOR2X1_LOC_647/B NOR2X1_LOC_6/B 0.03fF
C52683 INVX1_LOC_17/A INVX1_LOC_2/A 0.22fF
C52684 NAND2X1_LOC_222/A INVX1_LOC_75/A 0.01fF
C52685 INVX1_LOC_206/A NOR2X1_LOC_457/A 0.20fF
C52686 INVX1_LOC_238/Y NAND2X1_LOC_736/Y 0.25fF
C52687 INVX1_LOC_277/A INVX1_LOC_41/A 0.10fF
C52688 NOR2X1_LOC_541/Y INVX1_LOC_177/A 0.00fF
C52689 INVX1_LOC_17/A NOR2X1_LOC_226/A 0.15fF
C52690 NOR2X1_LOC_89/A NAND2X1_LOC_287/B 0.07fF
C52691 NAND2X1_LOC_579/A NAND2X1_LOC_859/B 0.03fF
C52692 INPUT_0 NOR2X1_LOC_720/A 0.00fF
C52693 NOR2X1_LOC_590/A NAND2X1_LOC_114/a_36_24# 0.01fF
C52694 INVX1_LOC_135/A INVX1_LOC_38/Y 0.11fF
C52695 INVX1_LOC_255/Y NAND2X1_LOC_214/Y 0.04fF
C52696 NOR2X1_LOC_328/Y INVX1_LOC_289/Y 0.01fF
C52697 INVX1_LOC_2/A NOR2X1_LOC_471/Y 0.03fF
C52698 NAND2X1_LOC_739/B NAND2X1_LOC_730/a_36_24# 0.02fF
C52699 NOR2X1_LOC_78/A NOR2X1_LOC_80/Y 0.01fF
C52700 INVX1_LOC_102/A INVX1_LOC_37/A 0.07fF
C52701 INVX1_LOC_284/Y NAND2X1_LOC_838/Y 0.14fF
C52702 NAND2X1_LOC_785/Y NAND2X1_LOC_785/B 0.10fF
C52703 NOR2X1_LOC_89/A INVX1_LOC_129/Y 0.01fF
C52704 INVX1_LOC_186/A NOR2X1_LOC_307/Y 0.22fF
C52705 NOR2X1_LOC_296/Y INVX1_LOC_40/A 0.03fF
C52706 NOR2X1_LOC_186/Y INVX1_LOC_313/A 0.03fF
C52707 INVX1_LOC_33/Y NOR2X1_LOC_669/A 0.01fF
C52708 NOR2X1_LOC_625/Y NAND2X1_LOC_837/Y 0.06fF
C52709 NAND2X1_LOC_84/Y INVX1_LOC_303/A 0.08fF
C52710 INVX1_LOC_238/Y INVX1_LOC_282/Y 0.40fF
C52711 NAND2X1_LOC_763/B NAND2X1_LOC_26/a_36_24# 0.07fF
C52712 NOR2X1_LOC_234/Y NOR2X1_LOC_384/Y 0.01fF
C52713 NOR2X1_LOC_585/a_36_216# INVX1_LOC_266/Y 0.00fF
C52714 NAND2X1_LOC_1/Y NAND2X1_LOC_3/B 0.10fF
C52715 INVX1_LOC_25/A NOR2X1_LOC_83/Y 0.01fF
C52716 INVX1_LOC_45/A INVX1_LOC_177/A 0.03fF
C52717 INPUT_3 INVX1_LOC_40/A 0.44fF
C52718 NOR2X1_LOC_180/a_36_216# NOR2X1_LOC_678/A 0.00fF
C52719 NOR2X1_LOC_210/A INVX1_LOC_11/A 0.03fF
C52720 INVX1_LOC_21/A INVX1_LOC_90/A 2.88fF
C52721 NOR2X1_LOC_667/Y NAND2X1_LOC_840/B 0.02fF
C52722 NOR2X1_LOC_186/Y NAND2X1_LOC_807/Y 0.07fF
C52723 NOR2X1_LOC_589/A INVX1_LOC_161/Y 0.07fF
C52724 NOR2X1_LOC_609/A INVX1_LOC_104/A 0.05fF
C52725 INVX1_LOC_225/A INVX1_LOC_111/A 0.03fF
C52726 NOR2X1_LOC_405/A NOR2X1_LOC_318/A 0.07fF
C52727 INVX1_LOC_75/A INVX1_LOC_213/A 2.01fF
C52728 NAND2X1_LOC_840/Y NOR2X1_LOC_109/Y 0.03fF
C52729 INVX1_LOC_299/A D_INPUT_0 0.03fF
C52730 INVX1_LOC_34/A NOR2X1_LOC_617/Y 0.02fF
C52731 NAND2X1_LOC_579/A NAND2X1_LOC_861/Y 0.10fF
C52732 INVX1_LOC_191/Y NOR2X1_LOC_584/a_36_216# 0.00fF
C52733 INVX1_LOC_223/Y NOR2X1_LOC_564/Y 0.04fF
C52734 NOR2X1_LOC_91/A NAND2X1_LOC_642/Y 0.16fF
C52735 NOR2X1_LOC_56/Y NOR2X1_LOC_449/A 0.08fF
C52736 NOR2X1_LOC_668/Y NAND2X1_LOC_642/Y 0.01fF
C52737 NAND2X1_LOC_374/Y NOR2X1_LOC_372/Y 0.19fF
C52738 NAND2X1_LOC_200/B INVX1_LOC_30/A 0.13fF
C52739 INVX1_LOC_26/A NOR2X1_LOC_368/Y 0.04fF
C52740 NOR2X1_LOC_361/B NOR2X1_LOC_123/B 0.10fF
C52741 NOR2X1_LOC_798/A NOR2X1_LOC_567/B 0.01fF
C52742 NOR2X1_LOC_470/B INVX1_LOC_295/A 0.01fF
C52743 NOR2X1_LOC_720/a_36_216# INVX1_LOC_62/Y 0.01fF
C52744 NAND2X1_LOC_583/a_36_24# NOR2X1_LOC_763/Y 0.03fF
C52745 NOR2X1_LOC_334/Y NOR2X1_LOC_139/a_36_216# 0.00fF
C52746 INVX1_LOC_11/A NOR2X1_LOC_312/Y 0.21fF
C52747 NAND2X1_LOC_787/A NOR2X1_LOC_528/Y 0.01fF
C52748 NOR2X1_LOC_537/A INVX1_LOC_104/A 0.04fF
C52749 INVX1_LOC_177/A INVX1_LOC_71/A 0.03fF
C52750 INVX1_LOC_21/A NAND2X1_LOC_348/A 0.10fF
C52751 NOR2X1_LOC_316/a_36_216# INVX1_LOC_46/A 0.00fF
C52752 INVX1_LOC_181/Y NOR2X1_LOC_190/a_36_216# 0.01fF
C52753 VDD NOR2X1_LOC_621/B -0.00fF
C52754 INPUT_0 NOR2X1_LOC_849/A 0.94fF
C52755 INVX1_LOC_293/A D_INPUT_0 0.01fF
C52756 INVX1_LOC_130/A INVX1_LOC_279/A 0.02fF
C52757 NAND2X1_LOC_182/A NOR2X1_LOC_716/B 0.02fF
C52758 INVX1_LOC_23/A NAND2X1_LOC_642/Y 0.03fF
C52759 VDD NOR2X1_LOC_449/A 0.18fF
C52760 NAND2X1_LOC_724/A NAND2X1_LOC_807/Y 0.08fF
C52761 INVX1_LOC_17/A INPUT_1 6.65fF
C52762 INVX1_LOC_26/A INVX1_LOC_46/A 0.07fF
C52763 NAND2X1_LOC_472/Y NOR2X1_LOC_465/Y 0.14fF
C52764 INVX1_LOC_36/A NAND2X1_LOC_112/Y 0.06fF
C52765 INVX1_LOC_50/A NAND2X1_LOC_655/B 0.01fF
C52766 INVX1_LOC_33/A NOR2X1_LOC_337/a_36_216# 0.00fF
C52767 INVX1_LOC_135/A NOR2X1_LOC_369/Y 0.06fF
C52768 NAND2X1_LOC_564/A NOR2X1_LOC_368/Y 0.05fF
C52769 NAND2X1_LOC_634/Y INVX1_LOC_16/A 0.08fF
C52770 NOR2X1_LOC_351/Y INVX1_LOC_32/A 0.04fF
C52771 INVX1_LOC_83/A INVX1_LOC_141/A 0.02fF
C52772 NOR2X1_LOC_98/A INVX1_LOC_26/A 0.05fF
C52773 NOR2X1_LOC_344/A NOR2X1_LOC_348/B 0.00fF
C52774 INVX1_LOC_69/Y INVX1_LOC_50/Y 0.07fF
C52775 NOR2X1_LOC_25/Y NOR2X1_LOC_425/Y 0.01fF
C52776 NOR2X1_LOC_186/Y INVX1_LOC_6/A 0.06fF
C52777 NOR2X1_LOC_536/Y NOR2X1_LOC_385/Y 0.00fF
C52778 NOR2X1_LOC_303/Y NOR2X1_LOC_357/a_36_216# 0.00fF
C52779 NAND2X1_LOC_848/A INVX1_LOC_94/Y 0.01fF
C52780 NOR2X1_LOC_577/Y NAND2X1_LOC_655/a_36_24# 0.00fF
C52781 INVX1_LOC_45/A NOR2X1_LOC_785/Y 0.06fF
C52782 NOR2X1_LOC_536/A INVX1_LOC_273/A 0.03fF
C52783 NOR2X1_LOC_361/B INVX1_LOC_102/Y 0.18fF
C52784 INVX1_LOC_135/A INVX1_LOC_286/Y 0.10fF
C52785 NOR2X1_LOC_195/A NAND2X1_LOC_508/A 0.00fF
C52786 NOR2X1_LOC_15/Y NOR2X1_LOC_313/a_36_216# 0.00fF
C52787 INVX1_LOC_251/Y NOR2X1_LOC_557/Y 0.15fF
C52788 NOR2X1_LOC_78/Y INVX1_LOC_3/Y 0.33fF
C52789 NAND2X1_LOC_555/Y INPUT_1 0.08fF
C52790 NOR2X1_LOC_92/Y NOR2X1_LOC_815/A 0.01fF
C52791 NOR2X1_LOC_91/A NOR2X1_LOC_495/a_36_216# 0.02fF
C52792 NOR2X1_LOC_474/A INVX1_LOC_197/Y 0.05fF
C52793 NOR2X1_LOC_68/A NOR2X1_LOC_719/B 0.04fF
C52794 VDD NOR2X1_LOC_493/A 0.02fF
C52795 NOR2X1_LOC_15/Y INVX1_LOC_126/Y 0.19fF
C52796 NOR2X1_LOC_155/A NOR2X1_LOC_467/A 0.16fF
C52797 NOR2X1_LOC_267/A NAND2X1_LOC_474/a_36_24# 0.05fF
C52798 INVX1_LOC_266/A INVX1_LOC_69/Y 0.10fF
C52799 INVX1_LOC_11/A NOR2X1_LOC_97/A 0.02fF
C52800 NOR2X1_LOC_301/A INVX1_LOC_118/A 3.89fF
C52801 INVX1_LOC_9/Y INVX1_LOC_33/A 0.03fF
C52802 INVX1_LOC_279/A INVX1_LOC_81/A 0.01fF
C52803 NOR2X1_LOC_441/Y NOR2X1_LOC_135/Y 0.02fF
C52804 NOR2X1_LOC_772/A INVX1_LOC_30/A 0.11fF
C52805 INVX1_LOC_90/A NAND2X1_LOC_354/Y 0.02fF
C52806 INVX1_LOC_11/A INVX1_LOC_193/Y 0.01fF
C52807 NAND2X1_LOC_61/Y INVX1_LOC_54/A 0.03fF
C52808 INVX1_LOC_109/A INVX1_LOC_29/A 0.01fF
C52809 NAND2X1_LOC_207/B NAND2X1_LOC_74/B 0.46fF
C52810 NAND2X1_LOC_721/B INVX1_LOC_28/A 0.05fF
C52811 NAND2X1_LOC_860/A INVX1_LOC_117/A 0.00fF
C52812 INVX1_LOC_30/A NOR2X1_LOC_19/B 0.09fF
C52813 NOR2X1_LOC_68/A NOR2X1_LOC_180/B 0.17fF
C52814 NOR2X1_LOC_13/Y INVX1_LOC_190/A 0.32fF
C52815 INVX1_LOC_251/Y INVX1_LOC_143/A 0.07fF
C52816 INVX1_LOC_16/A INVX1_LOC_8/A 0.17fF
C52817 NAND2X1_LOC_207/B NAND2X1_LOC_207/Y 0.03fF
C52818 NOR2X1_LOC_168/B INVX1_LOC_179/Y 0.02fF
C52819 INVX1_LOC_28/A NAND2X1_LOC_634/Y 0.08fF
C52820 NOR2X1_LOC_632/Y NOR2X1_LOC_142/Y 0.02fF
C52821 NOR2X1_LOC_634/Y INVX1_LOC_117/A 0.03fF
C52822 INVX1_LOC_23/A NOR2X1_LOC_271/Y 0.04fF
C52823 NOR2X1_LOC_68/A NOR2X1_LOC_738/A 0.06fF
C52824 NAND2X1_LOC_538/Y INVX1_LOC_91/A 1.23fF
C52825 NAND2X1_LOC_357/B INVX1_LOC_22/A 0.01fF
C52826 NOR2X1_LOC_514/A INPUT_0 0.13fF
C52827 NAND2X1_LOC_563/Y INVX1_LOC_255/Y 0.00fF
C52828 NOR2X1_LOC_45/Y INVX1_LOC_6/A 0.01fF
C52829 INVX1_LOC_75/A NOR2X1_LOC_707/B 0.29fF
C52830 NOR2X1_LOC_177/Y NAND2X1_LOC_439/a_36_24# 0.00fF
C52831 NOR2X1_LOC_541/B NOR2X1_LOC_197/B 0.05fF
C52832 NOR2X1_LOC_250/A INVX1_LOC_91/A 0.05fF
C52833 NAND2X1_LOC_53/Y NOR2X1_LOC_562/B 0.10fF
C52834 NAND2X1_LOC_728/Y NOR2X1_LOC_385/Y 0.14fF
C52835 NOR2X1_LOC_717/A INVX1_LOC_9/A 0.36fF
C52836 INVX1_LOC_83/A INVX1_LOC_103/Y 0.03fF
C52837 INVX1_LOC_135/A NOR2X1_LOC_542/a_36_216# 0.02fF
C52838 INVX1_LOC_83/A INVX1_LOC_315/A 0.31fF
C52839 INVX1_LOC_19/A INVX1_LOC_4/A 0.09fF
C52840 INVX1_LOC_75/A NOR2X1_LOC_546/A 0.01fF
C52841 INVX1_LOC_45/A INVX1_LOC_285/Y 0.03fF
C52842 NOR2X1_LOC_859/A INPUT_0 0.00fF
C52843 INVX1_LOC_76/A NAND2X1_LOC_780/Y 0.18fF
C52844 NOR2X1_LOC_415/A NOR2X1_LOC_6/B 0.06fF
C52845 NOR2X1_LOC_717/B INVX1_LOC_104/A 0.03fF
C52846 INVX1_LOC_35/A INVX1_LOC_274/A 0.46fF
C52847 INVX1_LOC_25/A NOR2X1_LOC_155/A 0.00fF
C52848 D_INPUT_0 NOR2X1_LOC_315/Y 0.03fF
C52849 NOR2X1_LOC_67/A NOR2X1_LOC_255/a_36_216# 0.00fF
C52850 INVX1_LOC_162/A NOR2X1_LOC_389/a_36_216# 0.02fF
C52851 INVX1_LOC_38/Y INVX1_LOC_280/A 0.03fF
C52852 NOR2X1_LOC_312/Y NOR2X1_LOC_52/B 0.07fF
C52853 NAND2X1_LOC_656/A NOR2X1_LOC_74/A 0.14fF
C52854 INVX1_LOC_105/Y INVX1_LOC_113/A 0.01fF
C52855 NAND2X1_LOC_310/a_36_24# INVX1_LOC_28/A 0.00fF
C52856 INVX1_LOC_30/A NOR2X1_LOC_528/Y 0.01fF
C52857 INPUT_0 INVX1_LOC_41/Y 0.03fF
C52858 NOR2X1_LOC_510/Y NOR2X1_LOC_331/B 0.08fF
C52859 INVX1_LOC_36/A INVX1_LOC_98/A 0.01fF
C52860 NOR2X1_LOC_78/B INVX1_LOC_164/A 0.09fF
C52861 INVX1_LOC_31/A NAND2X1_LOC_642/Y 0.13fF
C52862 INVX1_LOC_310/A D_INPUT_0 0.03fF
C52863 INVX1_LOC_1/Y INVX1_LOC_232/A 0.01fF
C52864 INVX1_LOC_144/Y INVX1_LOC_10/A -0.01fF
C52865 INVX1_LOC_21/A INVX1_LOC_38/A 26.35fF
C52866 INVX1_LOC_94/A NOR2X1_LOC_188/A 0.56fF
C52867 NOR2X1_LOC_848/Y VDD 0.46fF
C52868 NOR2X1_LOC_828/A INVX1_LOC_104/A 0.10fF
C52869 NOR2X1_LOC_218/a_36_216# NOR2X1_LOC_433/A 0.01fF
C52870 INVX1_LOC_161/Y INVX1_LOC_20/A 0.04fF
C52871 INVX1_LOC_28/A INVX1_LOC_8/A 0.07fF
C52872 INVX1_LOC_85/Y NOR2X1_LOC_731/A 0.01fF
C52873 INVX1_LOC_36/A NOR2X1_LOC_78/A 14.89fF
C52874 INVX1_LOC_94/A NOR2X1_LOC_548/B 0.14fF
C52875 NOR2X1_LOC_168/Y NOR2X1_LOC_548/a_36_216# 0.00fF
C52876 INVX1_LOC_11/A NAND2X1_LOC_287/B 0.25fF
C52877 INVX1_LOC_225/A NAND2X1_LOC_807/Y 0.03fF
C52878 INVX1_LOC_21/A NOR2X1_LOC_96/Y 0.03fF
C52879 NOR2X1_LOC_742/A NOR2X1_LOC_722/a_36_216# 0.01fF
C52880 INVX1_LOC_45/A INVX1_LOC_65/A 1.17fF
C52881 INVX1_LOC_285/Y INVX1_LOC_71/A 0.30fF
C52882 INVX1_LOC_89/A INVX1_LOC_210/A 0.06fF
C52883 NAND2X1_LOC_42/a_36_24# NAND2X1_LOC_215/A 0.00fF
C52884 D_INPUT_1 INVX1_LOC_84/A 0.14fF
C52885 NOR2X1_LOC_453/Y INVX1_LOC_38/A 0.65fF
C52886 NOR2X1_LOC_15/Y NOR2X1_LOC_536/A 0.19fF
C52887 NOR2X1_LOC_276/Y NAND2X1_LOC_211/Y 0.03fF
C52888 NOR2X1_LOC_717/B INVX1_LOC_263/A 0.06fF
C52889 NOR2X1_LOC_186/Y INVX1_LOC_131/Y 0.10fF
C52890 NOR2X1_LOC_667/A INVX1_LOC_90/A 0.13fF
C52891 INVX1_LOC_7/A NOR2X1_LOC_789/A 0.01fF
C52892 INVX1_LOC_141/Y INVX1_LOC_76/A 0.02fF
C52893 INVX1_LOC_248/A INVX1_LOC_90/A 0.09fF
C52894 INVX1_LOC_222/Y NOR2X1_LOC_650/a_36_216# 0.00fF
C52895 NAND2X1_LOC_787/A NAND2X1_LOC_477/Y 0.02fF
C52896 INVX1_LOC_24/A NOR2X1_LOC_45/B 0.90fF
C52897 NOR2X1_LOC_512/Y NAND2X1_LOC_655/A 0.01fF
C52898 NOR2X1_LOC_361/B NOR2X1_LOC_331/B 0.02fF
C52899 NOR2X1_LOC_798/A NOR2X1_LOC_79/Y 0.01fF
C52900 NAND2X1_LOC_866/B NAND2X1_LOC_852/Y 0.02fF
C52901 NOR2X1_LOC_599/A INVX1_LOC_20/A 0.03fF
C52902 INVX1_LOC_2/A NOR2X1_LOC_171/Y 0.06fF
C52903 INVX1_LOC_224/Y NAND2X1_LOC_81/B 0.07fF
C52904 NAND2X1_LOC_53/Y INVX1_LOC_281/Y 0.01fF
C52905 INVX1_LOC_312/Y INVX1_LOC_76/A 0.10fF
C52906 INVX1_LOC_141/Y NAND2X1_LOC_405/a_36_24# 0.00fF
C52907 NOR2X1_LOC_561/Y NAND2X1_LOC_656/Y 0.10fF
C52908 NAND2X1_LOC_573/Y INVX1_LOC_131/Y 0.12fF
C52909 INVX1_LOC_13/A INVX1_LOC_89/A 0.79fF
C52910 INVX1_LOC_225/A INVX1_LOC_6/A 0.07fF
C52911 INVX1_LOC_17/A INVX1_LOC_118/A 9.82fF
C52912 NAND2X1_LOC_383/a_36_24# INVX1_LOC_284/A 0.00fF
C52913 INVX1_LOC_24/A INVX1_LOC_247/A 0.03fF
C52914 NOR2X1_LOC_15/Y NAND2X1_LOC_93/B 0.06fF
C52915 NOR2X1_LOC_848/Y NOR2X1_LOC_846/a_36_216# 0.00fF
C52916 INVX1_LOC_14/A NOR2X1_LOC_99/Y 0.34fF
C52917 INVX1_LOC_305/A NOR2X1_LOC_857/A 0.00fF
C52918 NOR2X1_LOC_804/B NOR2X1_LOC_78/A 0.07fF
C52919 INVX1_LOC_84/A NOR2X1_LOC_652/Y 0.03fF
C52920 INVX1_LOC_64/A INVX1_LOC_19/A 0.13fF
C52921 INVX1_LOC_11/A NAND2X1_LOC_260/a_36_24# 0.00fF
C52922 NOR2X1_LOC_359/a_36_216# INVX1_LOC_92/A 0.00fF
C52923 INVX1_LOC_286/Y NOR2X1_LOC_152/A 0.02fF
C52924 NAND2X1_LOC_374/Y NAND2X1_LOC_844/a_36_24# 0.01fF
C52925 NAND2X1_LOC_14/a_36_24# INVX1_LOC_89/A 0.00fF
C52926 INVX1_LOC_63/Y INVX1_LOC_159/Y 0.01fF
C52927 INVX1_LOC_1/A NOR2X1_LOC_155/A 0.09fF
C52928 NOR2X1_LOC_78/B NOR2X1_LOC_368/A 0.03fF
C52929 INVX1_LOC_31/A NOR2X1_LOC_271/Y 0.00fF
C52930 NOR2X1_LOC_598/B INVX1_LOC_114/Y 0.03fF
C52931 NOR2X1_LOC_13/Y NAND2X1_LOC_649/a_36_24# 0.00fF
C52932 NOR2X1_LOC_473/B INVX1_LOC_10/A 0.08fF
C52933 INVX1_LOC_263/A NOR2X1_LOC_151/Y 0.01fF
C52934 INVX1_LOC_103/A NAND2X1_LOC_798/B 0.05fF
C52935 NOR2X1_LOC_48/B NOR2X1_LOC_452/A 0.08fF
C52936 NAND2X1_LOC_849/A INVX1_LOC_22/A 0.00fF
C52937 NOR2X1_LOC_309/Y NOR2X1_LOC_78/A 0.03fF
C52938 NOR2X1_LOC_32/B INVX1_LOC_42/A 0.09fF
C52939 NOR2X1_LOC_270/Y NAND2X1_LOC_472/Y 0.02fF
C52940 NOR2X1_LOC_237/Y NAND2X1_LOC_464/A 0.02fF
C52941 INVX1_LOC_269/A INVX1_LOC_285/A 0.10fF
C52942 NOR2X1_LOC_769/B NOR2X1_LOC_467/A 0.04fF
C52943 NOR2X1_LOC_15/Y INVX1_LOC_3/A 0.13fF
C52944 INVX1_LOC_102/Y NAND2X1_LOC_573/A 0.10fF
C52945 NAND2X1_LOC_860/A INVX1_LOC_3/Y 0.04fF
C52946 NOR2X1_LOC_219/B INVX1_LOC_76/A 0.03fF
C52947 INVX1_LOC_55/Y INVX1_LOC_89/A 0.04fF
C52948 INVX1_LOC_88/A NOR2X1_LOC_127/Y 0.15fF
C52949 INVX1_LOC_224/Y INVX1_LOC_4/Y 0.03fF
C52950 INVX1_LOC_163/Y INVX1_LOC_242/A 0.01fF
C52951 INVX1_LOC_24/A INVX1_LOC_281/A 0.07fF
C52952 NOR2X1_LOC_598/B NOR2X1_LOC_467/A 0.60fF
C52953 INVX1_LOC_269/A NOR2X1_LOC_814/A 0.02fF
C52954 NOR2X1_LOC_598/B NOR2X1_LOC_801/B 0.05fF
C52955 INVX1_LOC_283/Y INVX1_LOC_139/Y 0.00fF
C52956 INVX1_LOC_220/Y NOR2X1_LOC_74/A 0.00fF
C52957 INVX1_LOC_163/A NAND2X1_LOC_82/Y 0.01fF
C52958 NOR2X1_LOC_388/Y VDD 0.59fF
C52959 NOR2X1_LOC_355/B NOR2X1_LOC_500/Y 0.52fF
C52960 INVX1_LOC_174/A NAND2X1_LOC_426/a_36_24# -0.00fF
C52961 INVX1_LOC_48/Y INVX1_LOC_29/A 0.03fF
C52962 NOR2X1_LOC_106/A INVX1_LOC_79/A 0.02fF
C52963 NAND2X1_LOC_182/A NAND2X1_LOC_633/Y 0.01fF
C52964 NOR2X1_LOC_315/Y NOR2X1_LOC_266/B 0.00fF
C52965 INVX1_LOC_8/A NOR2X1_LOC_133/a_36_216# 0.01fF
C52966 INVX1_LOC_85/A INVX1_LOC_37/A 0.04fF
C52967 INVX1_LOC_262/A NOR2X1_LOC_635/B 0.01fF
C52968 INVX1_LOC_232/Y INVX1_LOC_74/A 0.10fF
C52969 NOR2X1_LOC_486/B INVX1_LOC_117/A 0.08fF
C52970 NAND2X1_LOC_741/B NAND2X1_LOC_770/Y 0.06fF
C52971 INVX1_LOC_17/A NAND2X1_LOC_63/Y 0.04fF
C52972 INVX1_LOC_149/A INVX1_LOC_46/A 0.20fF
C52973 INVX1_LOC_93/Y INVX1_LOC_232/A 0.40fF
C52974 NAND2X1_LOC_198/B INVX1_LOC_70/A 0.08fF
C52975 NOR2X1_LOC_717/B INVX1_LOC_206/Y 0.03fF
C52976 NOR2X1_LOC_103/Y NAND2X1_LOC_81/B 0.03fF
C52977 NAND2X1_LOC_364/Y INVX1_LOC_9/A 0.03fF
C52978 INVX1_LOC_18/A NOR2X1_LOC_831/B 0.20fF
C52979 NOR2X1_LOC_635/A NAND2X1_LOC_639/A 0.05fF
C52980 NAND2X1_LOC_9/Y INVX1_LOC_26/A 2.21fF
C52981 NOR2X1_LOC_180/Y NAND2X1_LOC_472/Y 0.03fF
C52982 INVX1_LOC_90/A INVX1_LOC_311/A 0.03fF
C52983 NOR2X1_LOC_458/Y NOR2X1_LOC_331/B 0.03fF
C52984 INVX1_LOC_153/Y NOR2X1_LOC_331/B 0.19fF
C52985 NOR2X1_LOC_210/B NAND2X1_LOC_212/Y 0.01fF
C52986 NOR2X1_LOC_753/Y INVX1_LOC_54/A 0.05fF
C52987 INVX1_LOC_233/A INVX1_LOC_26/A 0.07fF
C52988 NOR2X1_LOC_210/A INVX1_LOC_199/A 0.24fF
C52989 NAND2X1_LOC_783/A NOR2X1_LOC_45/B 0.03fF
C52990 INVX1_LOC_1/Y NAND2X1_LOC_447/Y 0.08fF
C52991 INVX1_LOC_30/A NAND2X1_LOC_477/Y 0.03fF
C52992 INVX1_LOC_192/A NOR2X1_LOC_450/A 0.19fF
C52993 INVX1_LOC_77/A NOR2X1_LOC_640/Y 0.25fF
C52994 NOR2X1_LOC_667/Y INVX1_LOC_49/Y 0.00fF
C52995 INVX1_LOC_64/A INVX1_LOC_26/Y 0.03fF
C52996 NOR2X1_LOC_315/Y NAND2X1_LOC_848/A 0.03fF
C52997 INVX1_LOC_288/A NOR2X1_LOC_639/B 0.02fF
C52998 NOR2X1_LOC_366/B VDD 0.12fF
C52999 NAND2X1_LOC_785/Y INVX1_LOC_38/A 0.07fF
C53000 NOR2X1_LOC_304/Y NAND2X1_LOC_175/Y 0.04fF
C53001 NOR2X1_LOC_45/B NOR2X1_LOC_130/A 0.31fF
C53002 INVX1_LOC_174/A INPUT_7 0.33fF
C53003 NOR2X1_LOC_106/A INVX1_LOC_91/A 0.03fF
C53004 NOR2X1_LOC_392/Y NOR2X1_LOC_646/B 0.00fF
C53005 NOR2X1_LOC_717/B NOR2X1_LOC_600/Y 0.19fF
C53006 INVX1_LOC_34/A INVX1_LOC_185/A 0.05fF
C53007 INVX1_LOC_136/A NOR2X1_LOC_605/A 0.00fF
C53008 NOR2X1_LOC_789/A INVX1_LOC_76/A 0.01fF
C53009 NOR2X1_LOC_458/B NAND2X1_LOC_472/Y 0.03fF
C53010 INVX1_LOC_85/A NAND2X1_LOC_629/a_36_24# 0.00fF
C53011 NAND2X1_LOC_479/Y VDD 0.17fF
C53012 INVX1_LOC_278/A D_INPUT_1 0.07fF
C53013 INVX1_LOC_225/A NOR2X1_LOC_79/A 0.14fF
C53014 NOR2X1_LOC_772/B NOR2X1_LOC_383/B 2.00fF
C53015 NOR2X1_LOC_798/A INVX1_LOC_26/A 0.00fF
C53016 INVX1_LOC_214/A INVX1_LOC_38/A 0.03fF
C53017 NAND2X1_LOC_662/Y INVX1_LOC_37/A 0.11fF
C53018 NOR2X1_LOC_241/A INVX1_LOC_15/A 0.02fF
C53019 INVX1_LOC_135/A NAND2X1_LOC_659/B 0.16fF
C53020 NOR2X1_LOC_667/A INVX1_LOC_38/A 0.11fF
C53021 INVX1_LOC_225/A INVX1_LOC_131/Y 0.01fF
C53022 D_INPUT_2 INVX1_LOC_84/A 0.04fF
C53023 NOR2X1_LOC_730/Y INVX1_LOC_37/A 0.10fF
C53024 NOR2X1_LOC_103/Y NAND2X1_LOC_269/a_36_24# 0.00fF
C53025 INVX1_LOC_248/A INVX1_LOC_38/A 0.03fF
C53026 NOR2X1_LOC_254/A NAND2X1_LOC_253/a_36_24# 0.00fF
C53027 NOR2X1_LOC_667/A NAND2X1_LOC_264/a_36_24# 0.01fF
C53028 INVX1_LOC_200/Y NAND2X1_LOC_552/A 0.01fF
C53029 NAND2X1_LOC_656/Y INVX1_LOC_76/A 0.10fF
C53030 NAND2X1_LOC_840/B NOR2X1_LOC_536/A 0.29fF
C53031 NOR2X1_LOC_151/Y INVX1_LOC_206/Y 0.03fF
C53032 NAND2X1_LOC_9/Y NOR2X1_LOC_619/a_36_216# 0.01fF
C53033 NAND2X1_LOC_303/Y NOR2X1_LOC_409/B 0.03fF
C53034 INVX1_LOC_5/A NOR2X1_LOC_858/A 0.01fF
C53035 INVX1_LOC_13/Y NOR2X1_LOC_383/B 0.03fF
C53036 NOR2X1_LOC_562/B NOR2X1_LOC_302/Y 0.03fF
C53037 INVX1_LOC_276/A INVX1_LOC_54/A 0.08fF
C53038 NOR2X1_LOC_669/Y NAND2X1_LOC_175/Y 0.17fF
C53039 NOR2X1_LOC_186/Y INVX1_LOC_270/A 0.34fF
C53040 NOR2X1_LOC_130/a_36_216# INVX1_LOC_59/Y 0.00fF
C53041 INVX1_LOC_41/A NAND2X1_LOC_572/B 0.07fF
C53042 NAND2X1_LOC_807/Y NAND2X1_LOC_642/Y 0.03fF
C53043 INPUT_0 NOR2X1_LOC_368/a_36_216# 0.00fF
C53044 NOR2X1_LOC_103/Y INVX1_LOC_4/Y 0.11fF
C53045 INVX1_LOC_96/Y NAND2X1_LOC_93/B 0.01fF
C53046 NAND2X1_LOC_571/B INVX1_LOC_5/A 0.23fF
C53047 INVX1_LOC_90/A NOR2X1_LOC_670/Y 0.00fF
C53048 INVX1_LOC_135/A VDD 7.30fF
C53049 INVX1_LOC_17/Y INVX1_LOC_178/A 0.01fF
C53050 INVX1_LOC_279/A NOR2X1_LOC_363/Y 0.03fF
C53051 NAND2X1_LOC_383/a_36_24# NOR2X1_LOC_384/A 0.00fF
C53052 NAND2X1_LOC_725/B NOR2X1_LOC_693/Y 0.05fF
C53053 NAND2X1_LOC_117/a_36_24# INVX1_LOC_46/A 0.01fF
C53054 INVX1_LOC_295/A VDD -0.00fF
C53055 NOR2X1_LOC_151/Y NOR2X1_LOC_600/Y 0.00fF
C53056 NOR2X1_LOC_824/A NAND2X1_LOC_458/a_36_24# 0.00fF
C53057 NOR2X1_LOC_188/A NOR2X1_LOC_845/A 0.07fF
C53058 NOR2X1_LOC_828/B NOR2X1_LOC_833/Y 0.03fF
C53059 INVX1_LOC_50/A INVX1_LOC_52/Y 0.22fF
C53060 INVX1_LOC_143/A NOR2X1_LOC_862/B 0.33fF
C53061 NOR2X1_LOC_92/Y NOR2X1_LOC_654/A 0.08fF
C53062 INVX1_LOC_35/A INVX1_LOC_306/Y 0.03fF
C53063 NAND2X1_LOC_555/Y NAND2X1_LOC_618/Y 0.02fF
C53064 NAND2X1_LOC_863/A INVX1_LOC_11/Y 0.11fF
C53065 NOR2X1_LOC_87/B NAND2X1_LOC_574/A 0.02fF
C53066 NOR2X1_LOC_560/A VDD 0.14fF
C53067 NOR2X1_LOC_350/A INVX1_LOC_29/A 0.05fF
C53068 INVX1_LOC_18/A NAND2X1_LOC_430/B 0.01fF
C53069 D_INPUT_0 NAND2X1_LOC_96/A 0.54fF
C53070 INVX1_LOC_239/A INVX1_LOC_23/A 0.00fF
C53071 NOR2X1_LOC_82/A INVX1_LOC_23/Y 0.31fF
C53072 INVX1_LOC_135/A NAND2X1_LOC_463/a_36_24# 0.00fF
C53073 INVX1_LOC_72/A D_INPUT_5 0.12fF
C53074 NOR2X1_LOC_591/Y INVX1_LOC_84/A 0.03fF
C53075 INVX1_LOC_88/A NOR2X1_LOC_383/B 2.20fF
C53076 INVX1_LOC_5/A NAND2X1_LOC_746/a_36_24# 0.00fF
C53077 NOR2X1_LOC_211/Y NOR2X1_LOC_220/B 0.15fF
C53078 NAND2X1_LOC_141/A NOR2X1_LOC_649/B 0.67fF
C53079 NOR2X1_LOC_186/Y NOR2X1_LOC_109/Y 1.49fF
C53080 NOR2X1_LOC_490/Y VDD 0.20fF
C53081 VDD INVX1_LOC_169/Y 0.41fF
C53082 NOR2X1_LOC_778/A INVX1_LOC_15/A 0.26fF
C53083 INVX1_LOC_45/A INVX1_LOC_4/Y 0.10fF
C53084 NOR2X1_LOC_576/B NOR2X1_LOC_536/A 0.05fF
C53085 NOR2X1_LOC_529/Y INVX1_LOC_84/A -0.01fF
C53086 INVX1_LOC_85/Y INVX1_LOC_117/A 1.76fF
C53087 NOR2X1_LOC_15/Y NOR2X1_LOC_476/B 0.08fF
C53088 INVX1_LOC_58/A NAND2X1_LOC_537/Y 0.10fF
C53089 NOR2X1_LOC_568/A INVX1_LOC_4/Y 0.07fF
C53090 INVX1_LOC_6/A NAND2X1_LOC_642/Y 0.07fF
C53091 INVX1_LOC_54/Y NAND2X1_LOC_475/Y 0.10fF
C53092 NOR2X1_LOC_598/B INVX1_LOC_1/A 0.33fF
C53093 NAND2X1_LOC_569/A NAND2X1_LOC_74/B -0.01fF
C53094 NOR2X1_LOC_791/B NOR2X1_LOC_38/B 0.05fF
C53095 GATE_479 INVX1_LOC_92/A 0.01fF
C53096 INVX1_LOC_113/Y NOR2X1_LOC_470/a_36_216# 0.00fF
C53097 INVX1_LOC_223/A NAND2X1_LOC_72/B 0.00fF
C53098 NOR2X1_LOC_264/Y NAND2X1_LOC_74/B 0.12fF
C53099 NOR2X1_LOC_552/A NOR2X1_LOC_337/Y 0.02fF
C53100 NOR2X1_LOC_753/Y NOR2X1_LOC_48/B 0.07fF
C53101 NOR2X1_LOC_703/B NOR2X1_LOC_334/Y 0.01fF
C53102 NAND2X1_LOC_573/Y NOR2X1_LOC_109/Y 0.89fF
C53103 NOR2X1_LOC_775/a_36_216# INVX1_LOC_176/A 0.00fF
C53104 INVX1_LOC_64/A NOR2X1_LOC_122/A 0.49fF
C53105 INVX1_LOC_178/A NOR2X1_LOC_406/A 0.03fF
C53106 INVX1_LOC_182/Y NOR2X1_LOC_363/Y 0.01fF
C53107 NAND2X1_LOC_541/Y INVX1_LOC_63/A 0.06fF
C53108 NAND2X1_LOC_325/Y NOR2X1_LOC_48/B 0.03fF
C53109 NOR2X1_LOC_6/B NOR2X1_LOC_89/A 0.02fF
C53110 INVX1_LOC_12/Y INVX1_LOC_67/Y 0.03fF
C53111 INVX1_LOC_44/Y INVX1_LOC_19/A 0.01fF
C53112 NOR2X1_LOC_391/B VDD 0.16fF
C53113 INVX1_LOC_28/A INVX1_LOC_118/Y 0.09fF
C53114 NAND2X1_LOC_850/Y INVX1_LOC_19/A 0.07fF
C53115 INVX1_LOC_78/Y INVX1_LOC_76/A 0.00fF
C53116 NOR2X1_LOC_711/A VDD 0.21fF
C53117 INVX1_LOC_71/A INVX1_LOC_4/Y 0.57fF
C53118 NOR2X1_LOC_318/B NAND2X1_LOC_447/Y 0.19fF
C53119 INVX1_LOC_286/A NOR2X1_LOC_558/A 0.01fF
C53120 INVX1_LOC_216/A INVX1_LOC_29/A 0.05fF
C53121 NOR2X1_LOC_791/A NAND2X1_LOC_99/A -0.01fF
C53122 INVX1_LOC_64/A INVX1_LOC_161/Y 1.65fF
C53123 NOR2X1_LOC_706/Y NOR2X1_LOC_706/B 0.03fF
C53124 NOR2X1_LOC_171/Y INVX1_LOC_118/A 0.04fF
C53125 NOR2X1_LOC_447/Y INVX1_LOC_78/A 0.03fF
C53126 INVX1_LOC_89/A NOR2X1_LOC_259/B 0.05fF
C53127 NAND2X1_LOC_51/B INVX1_LOC_38/A 2.99fF
C53128 INVX1_LOC_144/Y INVX1_LOC_12/A 0.01fF
C53129 INVX1_LOC_97/Y NOR2X1_LOC_794/B 0.00fF
C53130 NOR2X1_LOC_91/A NOR2X1_LOC_91/Y 0.13fF
C53131 INVX1_LOC_93/Y NAND2X1_LOC_447/Y 0.15fF
C53132 INVX1_LOC_224/A INVX1_LOC_50/Y 0.10fF
C53133 INVX1_LOC_49/A INVX1_LOC_94/Y 1.21fF
C53134 NOR2X1_LOC_143/a_36_216# INVX1_LOC_3/Y 0.01fF
C53135 NAND2X1_LOC_540/a_36_24# NOR2X1_LOC_103/Y 0.00fF
C53136 INVX1_LOC_11/A INVX1_LOC_50/Y 0.03fF
C53137 INVX1_LOC_276/A NOR2X1_LOC_48/B 0.28fF
C53138 INVX1_LOC_316/Y NAND2X1_LOC_74/B 0.09fF
C53139 INVX1_LOC_79/Y INVX1_LOC_270/Y 0.01fF
C53140 INVX1_LOC_311/A INVX1_LOC_38/A 0.03fF
C53141 NOR2X1_LOC_124/B NOR2X1_LOC_38/B 0.03fF
C53142 INVX1_LOC_151/Y INVX1_LOC_109/A 0.02fF
C53143 NOR2X1_LOC_552/A VDD 0.96fF
C53144 NOR2X1_LOC_337/A INVX1_LOC_9/A 0.03fF
C53145 NAND2X1_LOC_218/B NAND2X1_LOC_222/A 0.03fF
C53146 INVX1_LOC_285/Y NOR2X1_LOC_331/B 0.10fF
C53147 NOR2X1_LOC_816/A NOR2X1_LOC_406/A 0.01fF
C53148 NOR2X1_LOC_156/B NOR2X1_LOC_467/A 0.04fF
C53149 INVX1_LOC_6/A NOR2X1_LOC_271/Y 0.03fF
C53150 INVX1_LOC_290/A INVX1_LOC_29/A 0.11fF
C53151 NOR2X1_LOC_87/a_36_216# INVX1_LOC_15/A 0.02fF
C53152 INVX1_LOC_192/Y D_INPUT_5 0.18fF
C53153 INVX1_LOC_14/A NOR2X1_LOC_271/B 0.03fF
C53154 INVX1_LOC_149/Y NAND2X1_LOC_72/B 0.02fF
C53155 NOR2X1_LOC_790/B INVX1_LOC_18/A 0.07fF
C53156 INPUT_0 INVX1_LOC_185/A 0.04fF
C53157 NOR2X1_LOC_359/Y INVX1_LOC_23/A 0.09fF
C53158 INVX1_LOC_30/Y NOR2X1_LOC_89/A 0.03fF
C53159 INVX1_LOC_266/A INVX1_LOC_11/A 0.12fF
C53160 INVX1_LOC_49/A INVX1_LOC_296/A 0.07fF
C53161 INVX1_LOC_212/Y NOR2X1_LOC_843/B 0.01fF
C53162 INVX1_LOC_256/A NOR2X1_LOC_15/Y 0.45fF
C53163 INVX1_LOC_172/Y INVX1_LOC_3/Y 0.26fF
C53164 INVX1_LOC_2/A INVX1_LOC_94/Y 0.06fF
C53165 NOR2X1_LOC_481/A INVX1_LOC_270/A 0.10fF
C53166 INVX1_LOC_93/A INVX1_LOC_30/A 0.41fF
C53167 NOR2X1_LOC_123/B NAND2X1_LOC_81/B 0.06fF
C53168 NOR2X1_LOC_294/Y NOR2X1_LOC_34/B 0.03fF
C53169 NOR2X1_LOC_186/Y INVX1_LOC_36/A 0.25fF
C53170 INVX1_LOC_57/Y INVX1_LOC_13/Y 0.00fF
C53171 NOR2X1_LOC_757/A INVX1_LOC_290/Y 0.05fF
C53172 INVX1_LOC_50/A INVX1_LOC_63/Y 0.10fF
C53173 NOR2X1_LOC_226/A INVX1_LOC_94/Y 0.10fF
C53174 INVX1_LOC_77/A NOR2X1_LOC_247/Y 0.22fF
C53175 VDD INVX1_LOC_139/Y 0.63fF
C53176 NOR2X1_LOC_111/A NOR2X1_LOC_305/Y 0.09fF
C53177 NOR2X1_LOC_679/Y INVX1_LOC_103/A 0.13fF
C53178 INVX1_LOC_166/A NOR2X1_LOC_459/B 0.04fF
C53179 NOR2X1_LOC_646/A NOR2X1_LOC_38/B 0.07fF
C53180 INVX1_LOC_64/A NOR2X1_LOC_437/Y 0.32fF
C53181 INVX1_LOC_225/A INVX1_LOC_270/A 0.06fF
C53182 NAND2X1_LOC_849/B NOR2X1_LOC_670/Y 0.02fF
C53183 INVX1_LOC_269/A NOR2X1_LOC_590/A 0.19fF
C53184 NOR2X1_LOC_209/A NOR2X1_LOC_499/B 0.12fF
C53185 INVX1_LOC_36/A NAND2X1_LOC_573/Y 0.36fF
C53186 NOR2X1_LOC_813/Y VDD 1.56fF
C53187 NOR2X1_LOC_71/a_36_216# NAND2X1_LOC_572/B 0.01fF
C53188 NOR2X1_LOC_658/Y NAND2X1_LOC_67/Y 0.07fF
C53189 INVX1_LOC_34/A NOR2X1_LOC_754/Y 0.00fF
C53190 INVX1_LOC_10/Y VDD 0.54fF
C53191 NOR2X1_LOC_390/a_36_216# INVX1_LOC_53/A 0.01fF
C53192 NOR2X1_LOC_186/Y INVX1_LOC_145/A 0.03fF
C53193 INVX1_LOC_232/A INVX1_LOC_87/A 0.03fF
C53194 INVX1_LOC_36/A NAND2X1_LOC_724/A 0.07fF
C53195 INVX1_LOC_2/A INVX1_LOC_296/A 0.03fF
C53196 INVX1_LOC_102/Y NAND2X1_LOC_81/B 0.07fF
C53197 NAND2X1_LOC_571/B NAND2X1_LOC_562/B 0.08fF
C53198 NOR2X1_LOC_226/A INVX1_LOC_181/A 0.19fF
C53199 VDD INVX1_LOC_280/A 3.68fF
C53200 VDD NOR2X1_LOC_94/Y 0.02fF
C53201 INVX1_LOC_172/A NAND2X1_LOC_169/Y 0.07fF
C53202 NOR2X1_LOC_613/Y INVX1_LOC_24/A 0.01fF
C53203 INVX1_LOC_177/A NOR2X1_LOC_493/A 0.01fF
C53204 INVX1_LOC_5/A NAND2X1_LOC_361/Y 0.07fF
C53205 NOR2X1_LOC_203/Y NOR2X1_LOC_383/B 0.01fF
C53206 NOR2X1_LOC_604/a_36_216# INVX1_LOC_266/Y 0.00fF
C53207 INVX1_LOC_89/A INVX1_LOC_32/A 0.47fF
C53208 INVX1_LOC_11/A NOR2X1_LOC_248/Y 0.01fF
C53209 NOR2X1_LOC_256/a_36_216# INVX1_LOC_48/Y 0.00fF
C53210 INPUT_5 NOR2X1_LOC_30/Y 0.02fF
C53211 INVX1_LOC_247/A NOR2X1_LOC_197/B 0.01fF
C53212 NAND2X1_LOC_848/Y NOR2X1_LOC_670/Y 0.18fF
C53213 INVX1_LOC_98/A INVX1_LOC_63/A 0.19fF
C53214 INVX1_LOC_6/A NOR2X1_LOC_48/Y 0.00fF
C53215 INVX1_LOC_5/A INVX1_LOC_219/Y 0.03fF
C53216 INVX1_LOC_21/A INVX1_LOC_33/A 0.26fF
C53217 INVX1_LOC_250/A NOR2X1_LOC_816/A 0.08fF
C53218 NOR2X1_LOC_236/a_36_216# INVX1_LOC_23/Y 0.01fF
C53219 NOR2X1_LOC_206/a_36_216# INVX1_LOC_63/Y 0.01fF
C53220 NOR2X1_LOC_78/A INVX1_LOC_63/A 0.33fF
C53221 NOR2X1_LOC_405/a_36_216# INVX1_LOC_58/Y 0.01fF
C53222 INVX1_LOC_90/A NOR2X1_LOC_248/A 0.02fF
C53223 NOR2X1_LOC_186/Y NOR2X1_LOC_309/Y 0.02fF
C53224 NOR2X1_LOC_92/Y NOR2X1_LOC_716/B 0.07fF
C53225 INVX1_LOC_306/A INVX1_LOC_23/Y 0.02fF
C53226 INVX1_LOC_175/Y INVX1_LOC_253/A 0.01fF
C53227 INVX1_LOC_299/A INVX1_LOC_49/A 0.03fF
C53228 NOR2X1_LOC_389/B NOR2X1_LOC_248/A 0.01fF
C53229 INVX1_LOC_224/A NOR2X1_LOC_559/B 0.02fF
C53230 NAND2X1_LOC_819/a_36_24# NOR2X1_LOC_649/B 0.01fF
C53231 NAND2X1_LOC_862/A NAND2X1_LOC_793/B 0.01fF
C53232 NOR2X1_LOC_770/B NOR2X1_LOC_376/A 0.04fF
C53233 INVX1_LOC_266/A NOR2X1_LOC_593/Y 0.02fF
C53234 NAND2X1_LOC_341/A INVX1_LOC_53/A 0.02fF
C53235 NOR2X1_LOC_457/A NOR2X1_LOC_303/Y 0.18fF
C53236 INVX1_LOC_48/Y INVX1_LOC_8/A 0.03fF
C53237 NOR2X1_LOC_32/B NAND2X1_LOC_859/B 0.04fF
C53238 INVX1_LOC_31/A NOR2X1_LOC_91/Y 2.23fF
C53239 INVX1_LOC_316/Y NOR2X1_LOC_660/Y 0.01fF
C53240 NAND2X1_LOC_88/a_36_24# INVX1_LOC_50/Y 0.01fF
C53241 NOR2X1_LOC_543/A INVX1_LOC_23/A 0.15fF
C53242 INVX1_LOC_14/A NAND2X1_LOC_494/a_36_24# 0.00fF
C53243 INVX1_LOC_208/A NOR2X1_LOC_665/Y 0.23fF
C53244 INVX1_LOC_279/A INVX1_LOC_29/Y 0.06fF
C53245 NOR2X1_LOC_815/Y INVX1_LOC_17/A 0.02fF
C53246 NAND2X1_LOC_350/A INVX1_LOC_180/A 0.09fF
C53247 INVX1_LOC_13/A NOR2X1_LOC_392/Y 2.63fF
C53248 INVX1_LOC_11/A NOR2X1_LOC_718/Y 0.04fF
C53249 INVX1_LOC_35/A NAND2X1_LOC_149/B 0.02fF
C53250 NOR2X1_LOC_60/a_36_216# INVX1_LOC_271/A 0.00fF
C53251 NAND2X1_LOC_842/B INVX1_LOC_26/A 0.23fF
C53252 NAND2X1_LOC_244/A NAND2X1_LOC_489/Y 0.45fF
C53253 NOR2X1_LOC_389/A INVX1_LOC_81/A 0.17fF
C53254 NOR2X1_LOC_773/Y NOR2X1_LOC_406/A 0.01fF
C53255 NOR2X1_LOC_510/Y NOR2X1_LOC_366/B 0.05fF
C53256 INVX1_LOC_79/A NOR2X1_LOC_334/Y 0.02fF
C53257 INVX1_LOC_12/Y INVX1_LOC_285/A 0.10fF
C53258 INVX1_LOC_25/Y NOR2X1_LOC_293/a_36_216# 0.00fF
C53259 NAND2X1_LOC_724/Y INVX1_LOC_173/Y 0.91fF
C53260 NAND2X1_LOC_222/B NOR2X1_LOC_6/B 0.77fF
C53261 INVX1_LOC_224/A NOR2X1_LOC_6/B 0.01fF
C53262 INVX1_LOC_233/A INVX1_LOC_164/A 0.35fF
C53263 INVX1_LOC_14/Y NOR2X1_LOC_257/Y 0.01fF
C53264 NOR2X1_LOC_176/a_36_216# INVX1_LOC_63/A 0.00fF
C53265 NOR2X1_LOC_121/A INVX1_LOC_306/Y 0.02fF
C53266 INVX1_LOC_89/A NOR2X1_LOC_622/A 0.02fF
C53267 INVX1_LOC_12/Y NOR2X1_LOC_814/A 0.01fF
C53268 INVX1_LOC_30/A NOR2X1_LOC_303/Y 0.07fF
C53269 INVX1_LOC_2/A INVX1_LOC_299/A 0.10fF
C53270 INVX1_LOC_218/Y NOR2X1_LOC_520/B 0.01fF
C53271 INVX1_LOC_279/Y NOR2X1_LOC_551/B 0.10fF
C53272 NOR2X1_LOC_524/Y INVX1_LOC_49/A 0.09fF
C53273 NOR2X1_LOC_60/Y INVX1_LOC_63/A 0.03fF
C53274 INVX1_LOC_299/A NOR2X1_LOC_226/A 0.45fF
C53275 NOR2X1_LOC_389/A INVX1_LOC_192/A 0.00fF
C53276 INVX1_LOC_117/A NAND2X1_LOC_782/B 0.01fF
C53277 INVX1_LOC_196/Y INVX1_LOC_53/A 0.17fF
C53278 INVX1_LOC_256/A INVX1_LOC_96/Y 0.15fF
C53279 INVX1_LOC_54/Y NOR2X1_LOC_457/A 0.01fF
C53280 INVX1_LOC_131/A INVX1_LOC_270/Y 0.00fF
C53281 INVX1_LOC_200/Y INVX1_LOC_140/A 0.00fF
C53282 NOR2X1_LOC_75/Y NOR2X1_LOC_207/A 0.01fF
C53283 NAND2X1_LOC_66/a_36_24# NOR2X1_LOC_232/Y 0.00fF
C53284 INVX1_LOC_118/A NOR2X1_LOC_430/Y 0.10fF
C53285 NOR2X1_LOC_361/B NOR2X1_LOC_366/B 0.46fF
C53286 NOR2X1_LOC_134/Y NOR2X1_LOC_315/Y 0.01fF
C53287 NAND2X1_LOC_347/B INVX1_LOC_22/A 0.00fF
C53288 INVX1_LOC_182/Y INVX1_LOC_29/Y 0.34fF
C53289 INVX1_LOC_45/A NOR2X1_LOC_843/A 0.03fF
C53290 INVX1_LOC_268/A NAND2X1_LOC_213/A 0.01fF
C53291 NOR2X1_LOC_334/Y INVX1_LOC_91/A 0.07fF
C53292 INVX1_LOC_207/A INVX1_LOC_72/A 8.76fF
C53293 INVX1_LOC_178/A NAND2X1_LOC_319/A 0.00fF
C53294 NAND2X1_LOC_728/Y NOR2X1_LOC_387/Y 0.02fF
C53295 INVX1_LOC_35/A NOR2X1_LOC_356/A 0.05fF
C53296 INVX1_LOC_269/A NOR2X1_LOC_82/Y 0.01fF
C53297 NOR2X1_LOC_659/a_36_216# INVX1_LOC_63/Y 0.00fF
C53298 INVX1_LOC_311/Y NOR2X1_LOC_678/A 0.14fF
C53299 NAND2X1_LOC_557/Y INVX1_LOC_282/A 0.03fF
C53300 NOR2X1_LOC_510/Y INVX1_LOC_135/A 0.11fF
C53301 INVX1_LOC_246/Y NAND2X1_LOC_593/Y 0.19fF
C53302 NOR2X1_LOC_536/A INVX1_LOC_49/Y 0.05fF
C53303 INVX1_LOC_18/A NOR2X1_LOC_344/A 0.00fF
C53304 INVX1_LOC_37/A INVX1_LOC_290/Y 0.01fF
C53305 INVX1_LOC_36/A INVX1_LOC_225/A 0.11fF
C53306 INVX1_LOC_136/A NAND2X1_LOC_569/A 0.03fF
C53307 NOR2X1_LOC_658/Y NOR2X1_LOC_367/B 0.03fF
C53308 NOR2X1_LOC_441/Y INVX1_LOC_133/Y 0.07fF
C53309 INVX1_LOC_230/Y NOR2X1_LOC_78/B 0.10fF
C53310 NOR2X1_LOC_440/Y NOR2X1_LOC_15/Y 0.72fF
C53311 NAND2X1_LOC_7/Y INVX1_LOC_314/Y 0.03fF
C53312 INVX1_LOC_12/A INVX1_LOC_281/Y 0.00fF
C53313 NOR2X1_LOC_82/A INVX1_LOC_232/A 0.08fF
C53314 INVX1_LOC_147/Y INVX1_LOC_128/A -0.00fF
C53315 NAND2X1_LOC_802/A NAND2X1_LOC_593/Y 0.01fF
C53316 INVX1_LOC_224/A INVX1_LOC_30/Y 0.01fF
C53317 INVX1_LOC_5/A NAND2X1_LOC_654/B 0.03fF
C53318 NAND2X1_LOC_471/Y NOR2X1_LOC_368/Y 0.18fF
C53319 INVX1_LOC_54/Y INVX1_LOC_30/A 0.16fF
C53320 NAND2X1_LOC_9/Y NOR2X1_LOC_368/A 0.01fF
C53321 NAND2X1_LOC_357/B INVX1_LOC_18/A 0.07fF
C53322 NOR2X1_LOC_334/A INVX1_LOC_57/A 0.07fF
C53323 NOR2X1_LOC_230/Y NAND2X1_LOC_231/Y 0.04fF
C53324 INVX1_LOC_269/A INVX1_LOC_227/A 0.01fF
C53325 NOR2X1_LOC_620/Y NOR2X1_LOC_545/A 0.00fF
C53326 NOR2X1_LOC_598/B NOR2X1_LOC_188/A 0.01fF
C53327 INVX1_LOC_118/Y INVX1_LOC_109/A 0.01fF
C53328 NOR2X1_LOC_424/a_36_216# INVX1_LOC_103/A 0.12fF
C53329 NAND2X1_LOC_447/Y INVX1_LOC_87/A 0.02fF
C53330 NOR2X1_LOC_536/A NAND2X1_LOC_288/a_36_24# 0.00fF
C53331 INVX1_LOC_35/A NOR2X1_LOC_74/A 0.10fF
C53332 INVX1_LOC_25/A INVX1_LOC_201/A 0.03fF
C53333 INVX1_LOC_2/Y NOR2X1_LOC_38/B 2.24fF
C53334 NOR2X1_LOC_644/B INVX1_LOC_263/A 0.27fF
C53335 NOR2X1_LOC_852/B NAND2X1_LOC_364/Y 0.01fF
C53336 NOR2X1_LOC_82/A NOR2X1_LOC_383/Y 0.19fF
C53337 NOR2X1_LOC_598/B NOR2X1_LOC_548/B 0.10fF
C53338 INVX1_LOC_128/Y INVX1_LOC_76/A 0.17fF
C53339 NAND2X1_LOC_149/Y D_GATE_366 0.07fF
C53340 D_INPUT_1 INVX1_LOC_123/A 0.07fF
C53341 INVX1_LOC_105/A INVX1_LOC_63/Y 0.01fF
C53342 NOR2X1_LOC_689/Y NAND2X1_LOC_688/a_36_24# 0.00fF
C53343 INVX1_LOC_125/Y INVX1_LOC_129/A 0.00fF
C53344 INVX1_LOC_242/Y NOR2X1_LOC_298/Y 0.07fF
C53345 NOR2X1_LOC_763/A INVX1_LOC_244/A 0.03fF
C53346 INVX1_LOC_49/A NAND2X1_LOC_157/a_36_24# 0.01fF
C53347 INVX1_LOC_35/A NOR2X1_LOC_9/Y 0.03fF
C53348 INVX1_LOC_41/A NOR2X1_LOC_716/B 0.10fF
C53349 NAND2X1_LOC_361/Y NAND2X1_LOC_366/A 0.03fF
C53350 NOR2X1_LOC_360/Y NOR2X1_LOC_537/Y 0.03fF
C53351 INVX1_LOC_250/A NOR2X1_LOC_773/Y 0.02fF
C53352 NAND2X1_LOC_338/B NOR2X1_LOC_360/Y 0.07fF
C53353 NAND2X1_LOC_354/Y NAND2X1_LOC_798/A 0.17fF
C53354 NOR2X1_LOC_799/a_36_216# INVX1_LOC_77/A 0.00fF
C53355 INVX1_LOC_40/Y NOR2X1_LOC_516/B 0.02fF
C53356 NOR2X1_LOC_246/A NAND2X1_LOC_357/A 0.03fF
C53357 INVX1_LOC_73/A NAND2X1_LOC_474/Y 0.41fF
C53358 INVX1_LOC_172/A NAND2X1_LOC_357/B 0.16fF
C53359 NOR2X1_LOC_92/Y NOR2X1_LOC_503/A 0.01fF
C53360 INVX1_LOC_150/Y NOR2X1_LOC_137/A 0.26fF
C53361 VDD NOR2X1_LOC_541/B 0.03fF
C53362 NOR2X1_LOC_593/Y NOR2X1_LOC_6/B 0.03fF
C53363 NOR2X1_LOC_716/B NAND2X1_LOC_477/A 0.10fF
C53364 NOR2X1_LOC_738/Y INVX1_LOC_85/Y 0.01fF
C53365 NOR2X1_LOC_727/B INVX1_LOC_76/A 0.06fF
C53366 INVX1_LOC_269/A NOR2X1_LOC_703/A 0.04fF
C53367 INVX1_LOC_310/A INVX1_LOC_49/A 0.07fF
C53368 INPUT_3 INVX1_LOC_89/A 0.15fF
C53369 NOR2X1_LOC_703/B NOR2X1_LOC_569/Y 0.02fF
C53370 INVX1_LOC_90/A INVX1_LOC_174/A 0.10fF
C53371 INVX1_LOC_225/A NOR2X1_LOC_309/Y 0.41fF
C53372 NOR2X1_LOC_382/Y INVX1_LOC_234/A 0.65fF
C53373 NOR2X1_LOC_61/Y INVX1_LOC_15/A 0.08fF
C53374 NOR2X1_LOC_127/Y INVX1_LOC_272/A 0.50fF
C53375 NAND2X1_LOC_722/a_36_24# NOR2X1_LOC_299/Y 0.01fF
C53376 D_INPUT_0 NAND2X1_LOC_577/A 0.01fF
C53377 INVX1_LOC_5/A INVX1_LOC_159/Y 0.03fF
C53378 NOR2X1_LOC_388/Y INVX1_LOC_177/A 0.01fF
C53379 NOR2X1_LOC_84/Y INVX1_LOC_8/A 0.19fF
C53380 INVX1_LOC_163/A NAND2X1_LOC_622/B 0.02fF
C53381 NAND2X1_LOC_859/Y NOR2X1_LOC_91/Y 0.00fF
C53382 NOR2X1_LOC_523/A NAND2X1_LOC_348/A 0.01fF
C53383 INVX1_LOC_41/A INVX1_LOC_98/Y 0.01fF
C53384 NAND2X1_LOC_642/Y NOR2X1_LOC_109/Y 0.07fF
C53385 INVX1_LOC_94/Y INVX1_LOC_118/A 0.02fF
C53386 INVX1_LOC_200/A NOR2X1_LOC_322/Y 0.89fF
C53387 NOR2X1_LOC_100/A NAND2X1_LOC_116/A 0.07fF
C53388 NOR2X1_LOC_720/B NOR2X1_LOC_721/A 0.00fF
C53389 NOR2X1_LOC_457/B INVX1_LOC_10/A 0.10fF
C53390 NOR2X1_LOC_537/A NOR2X1_LOC_211/A 0.02fF
C53391 NOR2X1_LOC_15/Y INVX1_LOC_69/Y 0.07fF
C53392 INVX1_LOC_2/A NOR2X1_LOC_315/Y 0.03fF
C53393 NOR2X1_LOC_730/a_36_216# NOR2X1_LOC_687/Y 0.00fF
C53394 NOR2X1_LOC_49/a_36_216# INVX1_LOC_3/Y 0.00fF
C53395 NOR2X1_LOC_13/Y NOR2X1_LOC_561/Y 0.10fF
C53396 NOR2X1_LOC_38/B NOR2X1_LOC_608/Y 0.06fF
C53397 INVX1_LOC_11/A NAND2X1_LOC_328/a_36_24# 0.00fF
C53398 NOR2X1_LOC_810/Y D_GATE_811 0.18fF
C53399 NOR2X1_LOC_226/A NOR2X1_LOC_315/Y 0.02fF
C53400 NAND2X1_LOC_862/a_36_24# INVX1_LOC_41/Y 0.00fF
C53401 INVX1_LOC_47/A NAND2X1_LOC_364/A 0.01fF
C53402 D_INPUT_0 NAND2X1_LOC_656/A 0.23fF
C53403 NOR2X1_LOC_272/Y INVX1_LOC_95/Y 0.10fF
C53404 INVX1_LOC_21/A NOR2X1_LOC_486/Y 0.03fF
C53405 NOR2X1_LOC_382/Y NOR2X1_LOC_19/B 0.01fF
C53406 INVX1_LOC_118/A INVX1_LOC_181/A 0.03fF
C53407 NOR2X1_LOC_91/Y NAND2X1_LOC_866/B 0.01fF
C53408 INVX1_LOC_223/A NAND2X1_LOC_369/a_36_24# 0.00fF
C53409 NOR2X1_LOC_620/Y NOR2X1_LOC_545/a_36_216# 0.00fF
C53410 NOR2X1_LOC_360/Y INVX1_LOC_313/Y 0.01fF
C53411 INVX1_LOC_136/A NAND2X1_LOC_850/A 0.03fF
C53412 INVX1_LOC_118/A INVX1_LOC_296/A 0.15fF
C53413 NOR2X1_LOC_67/A NOR2X1_LOC_655/B 0.10fF
C53414 NOR2X1_LOC_384/Y NAND2X1_LOC_560/A 0.02fF
C53415 INVX1_LOC_11/A INVX1_LOC_96/A 0.03fF
C53416 INVX1_LOC_2/A INVX1_LOC_52/A 0.02fF
C53417 INVX1_LOC_54/A NAND2X1_LOC_787/Y 0.00fF
C53418 INVX1_LOC_90/A NAND2X1_LOC_169/a_36_24# 0.00fF
C53419 NAND2X1_LOC_10/a_36_24# NOR2X1_LOC_536/A 0.00fF
C53420 NOR2X1_LOC_624/a_36_216# NOR2X1_LOC_78/A 0.00fF
C53421 NOR2X1_LOC_99/Y NOR2X1_LOC_383/B 0.01fF
C53422 NAND2X1_LOC_338/B NAND2X1_LOC_110/a_36_24# 0.01fF
C53423 INVX1_LOC_41/A NOR2X1_LOC_717/B 0.04fF
C53424 INVX1_LOC_18/A NAND2X1_LOC_849/A 0.09fF
C53425 INVX1_LOC_217/A NOR2X1_LOC_322/Y 0.19fF
C53426 INVX1_LOC_9/A NOR2X1_LOC_247/Y 0.07fF
C53427 NAND2X1_LOC_357/B NOR2X1_LOC_690/Y 0.05fF
C53428 NOR2X1_LOC_470/B INVX1_LOC_199/Y 0.01fF
C53429 NAND2X1_LOC_726/Y NOR2X1_LOC_667/A 0.08fF
C53430 NOR2X1_LOC_584/Y NOR2X1_LOC_48/B 0.03fF
C53431 NOR2X1_LOC_808/A NOR2X1_LOC_687/Y 0.13fF
C53432 NAND2X1_LOC_341/A NOR2X1_LOC_78/B 0.03fF
C53433 NOR2X1_LOC_456/Y INVX1_LOC_274/A 0.01fF
C53434 INVX1_LOC_271/A INVX1_LOC_180/Y 0.01fF
C53435 NAND2X1_LOC_796/B NAND2X1_LOC_721/A -0.00fF
C53436 INVX1_LOC_29/A NOR2X1_LOC_467/A 0.35fF
C53437 NOR2X1_LOC_454/Y INVX1_LOC_37/A 0.08fF
C53438 INVX1_LOC_72/A NOR2X1_LOC_427/Y 0.09fF
C53439 NOR2X1_LOC_605/B NOR2X1_LOC_667/A 0.02fF
C53440 NOR2X1_LOC_561/Y NOR2X1_LOC_504/Y 0.03fF
C53441 INVX1_LOC_41/A NOR2X1_LOC_828/A 0.01fF
C53442 NOR2X1_LOC_68/A NOR2X1_LOC_589/Y 0.05fF
C53443 NOR2X1_LOC_225/a_36_216# INVX1_LOC_93/Y 0.01fF
C53444 INVX1_LOC_286/Y NOR2X1_LOC_45/B 0.10fF
C53445 INVX1_LOC_135/A INVX1_LOC_177/A 0.06fF
C53446 INVX1_LOC_172/A NAND2X1_LOC_849/A 0.03fF
C53447 NOR2X1_LOC_688/Y NOR2X1_LOC_78/A 0.02fF
C53448 INVX1_LOC_89/A INVX1_LOC_158/A 0.05fF
C53449 NOR2X1_LOC_91/Y INVX1_LOC_6/A 0.01fF
C53450 NOR2X1_LOC_232/a_36_216# NAND2X1_LOC_721/A 0.01fF
C53451 INVX1_LOC_63/Y NAND2X1_LOC_652/Y 0.02fF
C53452 NOR2X1_LOC_315/Y INPUT_1 0.45fF
C53453 INVX1_LOC_17/A INVX1_LOC_14/Y 0.08fF
C53454 INVX1_LOC_45/A NOR2X1_LOC_595/Y 0.03fF
C53455 INVX1_LOC_181/Y INVX1_LOC_286/A 0.01fF
C53456 NOR2X1_LOC_67/A NOR2X1_LOC_99/B 0.59fF
C53457 INVX1_LOC_72/A NOR2X1_LOC_269/Y 0.07fF
C53458 NOR2X1_LOC_89/A INVX1_LOC_273/A 0.06fF
C53459 NOR2X1_LOC_831/Y NOR2X1_LOC_301/A 0.01fF
C53460 INVX1_LOC_90/A INVX1_LOC_259/A 0.01fF
C53461 INVX1_LOC_135/A NOR2X1_LOC_608/a_36_216# 0.01fF
C53462 INVX1_LOC_41/A NOR2X1_LOC_151/Y 0.24fF
C53463 NOR2X1_LOC_361/B NOR2X1_LOC_813/Y 0.10fF
C53464 INVX1_LOC_35/A NOR2X1_LOC_865/Y 0.01fF
C53465 INVX1_LOC_33/A NAND2X1_LOC_51/B 0.00fF
C53466 INVX1_LOC_36/A NAND2X1_LOC_642/Y 1.66fF
C53467 INVX1_LOC_203/A NAND2X1_LOC_464/B 0.41fF
C53468 INVX1_LOC_140/A NAND2X1_LOC_799/Y 0.44fF
C53469 INVX1_LOC_211/Y NAND2X1_LOC_453/A 0.15fF
C53470 NOR2X1_LOC_720/A INVX1_LOC_19/A 0.01fF
C53471 INVX1_LOC_35/A NOR2X1_LOC_243/B 0.07fF
C53472 INVX1_LOC_159/A NOR2X1_LOC_45/B 0.63fF
C53473 NOR2X1_LOC_471/Y INVX1_LOC_14/Y 0.03fF
C53474 NOR2X1_LOC_589/A NAND2X1_LOC_480/a_36_24# 0.00fF
C53475 NOR2X1_LOC_781/B NAND2X1_LOC_662/Y 0.00fF
C53476 NOR2X1_LOC_267/A NAND2X1_LOC_642/Y 0.03fF
C53477 NAND2X1_LOC_555/Y D_GATE_479 0.02fF
C53478 INVX1_LOC_26/A INVX1_LOC_284/A 0.01fF
C53479 NOR2X1_LOC_78/B INVX1_LOC_196/Y 0.03fF
C53480 NAND2X1_LOC_555/Y D_INPUT_3 0.14fF
C53481 INVX1_LOC_84/A NOR2X1_LOC_678/A 0.03fF
C53482 NOR2X1_LOC_361/B INVX1_LOC_280/A 0.21fF
C53483 NOR2X1_LOC_246/A INVX1_LOC_25/Y 0.12fF
C53484 NOR2X1_LOC_716/B NOR2X1_LOC_71/a_36_216# 0.01fF
C53485 INVX1_LOC_304/Y NOR2X1_LOC_322/Y 0.10fF
C53486 NOR2X1_LOC_658/Y INVX1_LOC_76/A 0.03fF
C53487 NOR2X1_LOC_205/Y NOR2X1_LOC_331/B 0.25fF
C53488 NAND2X1_LOC_63/Y NOR2X1_LOC_621/a_36_216# 0.01fF
C53489 NAND2X1_LOC_364/A INVX1_LOC_95/Y 0.07fF
C53490 INVX1_LOC_17/A INVX1_LOC_230/A 0.18fF
C53491 INVX1_LOC_11/A NOR2X1_LOC_684/Y 0.47fF
C53492 NOR2X1_LOC_644/A NOR2X1_LOC_544/A 0.03fF
C53493 INVX1_LOC_83/A GATE_479 0.07fF
C53494 NOR2X1_LOC_388/Y INVX1_LOC_285/Y 0.10fF
C53495 NOR2X1_LOC_278/Y INVX1_LOC_170/Y 0.00fF
C53496 INVX1_LOC_135/A NAND2X1_LOC_376/a_36_24# 0.01fF
C53497 INVX1_LOC_23/A NAND2X1_LOC_82/Y 0.07fF
C53498 INVX1_LOC_57/A NAND2X1_LOC_74/B 0.21fF
C53499 NOR2X1_LOC_590/A INVX1_LOC_12/Y 0.01fF
C53500 NOR2X1_LOC_180/B NOR2X1_LOC_500/Y 0.08fF
C53501 INVX1_LOC_305/Y NOR2X1_LOC_356/A 0.02fF
C53502 INVX1_LOC_181/Y INVX1_LOC_95/A 0.00fF
C53503 NAND2X1_LOC_551/A INVX1_LOC_25/Y 0.01fF
C53504 NAND2X1_LOC_7/Y NOR2X1_LOC_557/A 0.00fF
C53505 INVX1_LOC_10/A NOR2X1_LOC_335/a_36_216# 0.00fF
C53506 INVX1_LOC_14/A NOR2X1_LOC_612/Y 0.04fF
C53507 INVX1_LOC_25/A INVX1_LOC_29/A 0.07fF
C53508 NOR2X1_LOC_242/A NOR2X1_LOC_461/B 0.03fF
C53509 NOR2X1_LOC_34/Y INVX1_LOC_15/A 0.01fF
C53510 NOR2X1_LOC_478/A INVX1_LOC_117/A 0.03fF
C53511 INVX1_LOC_89/A GATE_662 0.35fF
C53512 NAND2X1_LOC_387/B VDD 0.01fF
C53513 NAND2X1_LOC_323/B NOR2X1_LOC_567/B 0.07fF
C53514 INVX1_LOC_174/A INVX1_LOC_38/A 0.23fF
C53515 INVX1_LOC_90/A NOR2X1_LOC_589/A 0.03fF
C53516 INVX1_LOC_57/A NOR2X1_LOC_847/B 0.09fF
C53517 INVX1_LOC_135/A NAND2X1_LOC_378/a_36_24# 0.00fF
C53518 NOR2X1_LOC_653/B INVX1_LOC_285/A 0.03fF
C53519 INVX1_LOC_17/Y INVX1_LOC_42/A 0.00fF
C53520 NOR2X1_LOC_255/Y INVX1_LOC_284/A 0.53fF
C53521 INVX1_LOC_200/Y INVX1_LOC_42/A 0.06fF
C53522 NOR2X1_LOC_389/B NOR2X1_LOC_589/A 0.07fF
C53523 NAND2X1_LOC_462/B NAND2X1_LOC_624/A 0.02fF
C53524 INVX1_LOC_23/A NOR2X1_LOC_461/Y 0.01fF
C53525 INVX1_LOC_24/A NOR2X1_LOC_603/Y 0.01fF
C53526 INVX1_LOC_81/A NAND2X1_LOC_469/B 0.03fF
C53527 NOR2X1_LOC_186/Y INVX1_LOC_63/A 1.38fF
C53528 NAND2X1_LOC_231/Y INVX1_LOC_126/Y 0.11fF
C53529 NOR2X1_LOC_13/Y INVX1_LOC_76/A 0.22fF
C53530 NOR2X1_LOC_329/B NAND2X1_LOC_660/Y 0.03fF
C53531 NOR2X1_LOC_794/A INVX1_LOC_177/A 0.01fF
C53532 NOR2X1_LOC_593/Y INVX1_LOC_188/Y 0.01fF
C53533 NOR2X1_LOC_68/A INVX1_LOC_117/A 4.32fF
C53534 INVX1_LOC_41/A NOR2X1_LOC_181/A 0.01fF
C53535 NOR2X1_LOC_172/Y INVX1_LOC_147/Y 0.00fF
C53536 INVX1_LOC_36/A NOR2X1_LOC_271/Y 0.03fF
C53537 NAND2X1_LOC_391/Y NAND2X1_LOC_773/B 0.01fF
C53538 NOR2X1_LOC_569/A NOR2X1_LOC_500/Y 0.01fF
C53539 INVX1_LOC_13/A INVX1_LOC_75/A 0.79fF
C53540 NOR2X1_LOC_304/a_36_216# INVX1_LOC_12/A 0.00fF
C53541 NOR2X1_LOC_309/Y NAND2X1_LOC_642/Y 0.07fF
C53542 INVX1_LOC_209/Y NOR2X1_LOC_421/Y 0.01fF
C53543 NOR2X1_LOC_388/Y NOR2X1_LOC_137/B 0.28fF
C53544 NAND2X1_LOC_573/Y INVX1_LOC_63/A 0.10fF
C53545 NAND2X1_LOC_319/A INVX1_LOC_140/A 0.23fF
C53546 NOR2X1_LOC_45/Y NOR2X1_LOC_435/A 0.03fF
C53547 NOR2X1_LOC_389/B INVX1_LOC_171/A 0.05fF
C53548 INVX1_LOC_77/A INVX1_LOC_37/A 0.16fF
C53549 NOR2X1_LOC_793/A NOR2X1_LOC_814/A 0.00fF
C53550 D_INPUT_0 NOR2X1_LOC_329/B 0.17fF
C53551 INVX1_LOC_314/Y INVX1_LOC_129/Y 0.02fF
C53552 INVX1_LOC_73/A INVX1_LOC_10/A 0.03fF
C53553 NOR2X1_LOC_570/A NOR2X1_LOC_188/A 0.01fF
C53554 NOR2X1_LOC_392/Y INVX1_LOC_32/A 0.16fF
C53555 NOR2X1_LOC_6/B INVX1_LOC_74/A 0.02fF
C53556 NOR2X1_LOC_678/A INVX1_LOC_15/A 0.11fF
C53557 NAND2X1_LOC_11/Y NOR2X1_LOC_588/A 0.00fF
C53558 NOR2X1_LOC_355/A INVX1_LOC_182/Y -0.04fF
C53559 NAND2X1_LOC_778/Y NOR2X1_LOC_89/A 0.10fF
C53560 NOR2X1_LOC_392/B INVX1_LOC_20/A 0.01fF
C53561 NOR2X1_LOC_545/A INVX1_LOC_117/A 0.04fF
C53562 NOR2X1_LOC_322/Y NAND2X1_LOC_808/A 0.04fF
C53563 INVX1_LOC_200/Y INVX1_LOC_78/A 0.02fF
C53564 INVX1_LOC_58/A NAND2X1_LOC_454/Y 0.17fF
C53565 INVX1_LOC_153/Y INVX1_LOC_139/Y 0.03fF
C53566 NAND2X1_LOC_364/A NAND2X1_LOC_289/a_36_24# 0.01fF
C53567 NAND2X1_LOC_116/A INVX1_LOC_176/A 0.03fF
C53568 INVX1_LOC_49/A NAND2X1_LOC_96/A 0.14fF
C53569 INVX1_LOC_277/A NOR2X1_LOC_155/A 0.11fF
C53570 NOR2X1_LOC_160/B INVX1_LOC_285/A 0.07fF
C53571 INVX1_LOC_292/A INVX1_LOC_220/A 0.31fF
C53572 INVX1_LOC_1/Y INVX1_LOC_98/A 0.11fF
C53573 NOR2X1_LOC_132/Y NOR2X1_LOC_813/Y 0.06fF
C53574 INVX1_LOC_1/A INVX1_LOC_29/A 0.20fF
C53575 INVX1_LOC_30/A INVX1_LOC_35/Y 0.05fF
C53576 NOR2X1_LOC_160/B NOR2X1_LOC_814/A 0.36fF
C53577 NAND2X1_LOC_633/Y NAND2X1_LOC_477/A 0.10fF
C53578 INVX1_LOC_1/Y NOR2X1_LOC_78/A 0.17fF
C53579 NOR2X1_LOC_795/Y VDD 1.06fF
C53580 NOR2X1_LOC_289/Y INVX1_LOC_28/A 0.40fF
C53581 INVX1_LOC_55/Y INVX1_LOC_75/A 0.03fF
C53582 NOR2X1_LOC_15/Y NOR2X1_LOC_89/A 1.27fF
C53583 INVX1_LOC_26/A NAND2X1_LOC_275/a_36_24# 0.00fF
C53584 NOR2X1_LOC_538/B NAND2X1_LOC_63/Y 0.00fF
C53585 NOR2X1_LOC_360/Y NOR2X1_LOC_79/a_36_216# 0.01fF
C53586 INVX1_LOC_153/Y INVX1_LOC_10/Y 0.01fF
C53587 NOR2X1_LOC_285/a_36_216# INVX1_LOC_26/Y 0.00fF
C53588 NAND2X1_LOC_839/Y VDD 0.01fF
C53589 NAND2X1_LOC_35/Y NOR2X1_LOC_394/Y 0.02fF
C53590 NOR2X1_LOC_457/B INVX1_LOC_307/A 0.03fF
C53591 NOR2X1_LOC_132/Y INVX1_LOC_280/A 0.01fF
C53592 INVX1_LOC_49/A NAND2X1_LOC_427/a_36_24# 0.01fF
C53593 INVX1_LOC_34/A NOR2X1_LOC_536/A 2.63fF
C53594 INVX1_LOC_251/Y VDD 0.44fF
C53595 INVX1_LOC_196/A NOR2X1_LOC_857/A 0.10fF
C53596 INVX1_LOC_256/Y INVX1_LOC_76/A 0.10fF
C53597 NAND2X1_LOC_342/Y NAND2X1_LOC_211/Y 0.07fF
C53598 INVX1_LOC_235/A INVX1_LOC_32/A 0.05fF
C53599 INVX1_LOC_90/A INVX1_LOC_222/A 0.05fF
C53600 INVX1_LOC_41/A NOR2X1_LOC_709/B 0.06fF
C53601 NOR2X1_LOC_550/B INVX1_LOC_274/A 0.19fF
C53602 INVX1_LOC_232/A INVX1_LOC_59/Y 0.01fF
C53603 INVX1_LOC_60/Y NOR2X1_LOC_98/B 0.20fF
C53604 NOR2X1_LOC_778/B NOR2X1_LOC_858/B 0.01fF
C53605 D_INPUT_1 NAND2X1_LOC_90/a_36_24# 0.01fF
C53606 NOR2X1_LOC_794/B INVX1_LOC_29/A 0.01fF
C53607 NAND2X1_LOC_393/a_36_24# INVX1_LOC_32/A 0.00fF
C53608 INVX1_LOC_13/Y INVX1_LOC_165/A 0.03fF
C53609 NAND2X1_LOC_729/B INVX1_LOC_10/A 0.00fF
C53610 NOR2X1_LOC_287/A NOR2X1_LOC_857/A 0.02fF
C53611 NAND2X1_LOC_276/Y NOR2X1_LOC_489/A 0.00fF
C53612 INVX1_LOC_31/A NAND2X1_LOC_82/Y 0.73fF
C53613 INVX1_LOC_162/A INVX1_LOC_118/A 0.72fF
C53614 NOR2X1_LOC_409/Y NAND2X1_LOC_463/B 0.20fF
C53615 NOR2X1_LOC_45/B NAND2X1_LOC_803/a_36_24# 0.01fF
C53616 NOR2X1_LOC_614/Y VDD 0.48fF
C53617 INVX1_LOC_230/Y NOR2X1_LOC_671/Y 0.04fF
C53618 NAND2X1_LOC_341/A INVX1_LOC_46/A 0.01fF
C53619 INVX1_LOC_136/A NOR2X1_LOC_662/A 0.07fF
C53620 NAND2X1_LOC_662/Y NOR2X1_LOC_585/Y 0.01fF
C53621 NAND2X1_LOC_811/Y INVX1_LOC_185/A 0.00fF
C53622 INVX1_LOC_57/A NOR2X1_LOC_660/Y 0.03fF
C53623 INVX1_LOC_90/A NOR2X1_LOC_311/a_36_216# 0.00fF
C53624 NAND2X1_LOC_231/Y NOR2X1_LOC_536/A 0.27fF
C53625 NOR2X1_LOC_315/Y INVX1_LOC_118/A 0.06fF
C53626 INVX1_LOC_34/A NAND2X1_LOC_93/B 0.10fF
C53627 INVX1_LOC_36/A NOR2X1_LOC_48/Y 0.03fF
C53628 NOR2X1_LOC_534/a_36_216# NOR2X1_LOC_74/A 0.01fF
C53629 INVX1_LOC_135/A INVX1_LOC_316/A 0.03fF
C53630 INVX1_LOC_142/A INVX1_LOC_19/A 0.33fF
C53631 NOR2X1_LOC_687/Y INVX1_LOC_37/A 0.07fF
C53632 NAND2X1_LOC_787/A NAND2X1_LOC_860/A 0.05fF
C53633 NAND2X1_LOC_357/A INVX1_LOC_32/A 0.14fF
C53634 INVX1_LOC_13/Y NOR2X1_LOC_693/Y 0.00fF
C53635 INVX1_LOC_26/Y NOR2X1_LOC_849/A 0.15fF
C53636 NAND2X1_LOC_725/Y NAND2X1_LOC_725/A 0.02fF
C53637 INVX1_LOC_50/A NAND2X1_LOC_552/A 0.01fF
C53638 NOR2X1_LOC_82/Y INVX1_LOC_12/Y 0.07fF
C53639 INVX1_LOC_47/A NOR2X1_LOC_405/A 0.17fF
C53640 INVX1_LOC_280/Y INVX1_LOC_280/A 0.10fF
C53641 INVX1_LOC_144/A NOR2X1_LOC_815/A 0.01fF
C53642 INVX1_LOC_50/A INVX1_LOC_5/A 0.55fF
C53643 NOR2X1_LOC_791/Y NAND2X1_LOC_286/B 0.07fF
C53644 NAND2X1_LOC_144/a_36_24# NOR2X1_LOC_706/A 0.01fF
C53645 INPUT_0 INVX1_LOC_126/Y 0.19fF
C53646 NOR2X1_LOC_612/B NOR2X1_LOC_612/Y 0.02fF
C53647 NOR2X1_LOC_608/a_36_216# INVX1_LOC_280/A 0.02fF
C53648 INVX1_LOC_26/Y NOR2X1_LOC_852/Y 0.01fF
C53649 NOR2X1_LOC_384/Y INVX1_LOC_29/A 0.22fF
C53650 INVX1_LOC_208/A NOR2X1_LOC_366/a_36_216# 0.01fF
C53651 INVX1_LOC_155/A NOR2X1_LOC_117/a_36_216# 0.00fF
C53652 INVX1_LOC_5/A NOR2X1_LOC_105/Y 0.16fF
C53653 INVX1_LOC_277/A NOR2X1_LOC_833/B 0.04fF
C53654 INVX1_LOC_21/A NOR2X1_LOC_635/B 0.53fF
C53655 NOR2X1_LOC_418/Y INVX1_LOC_38/A 0.04fF
C53656 NOR2X1_LOC_516/B NOR2X1_LOC_862/a_36_216# 0.13fF
C53657 INVX1_LOC_298/Y INVX1_LOC_1/A 0.07fF
C53658 INVX1_LOC_21/A INVX1_LOC_275/Y 0.11fF
C53659 NOR2X1_LOC_528/Y NOR2X1_LOC_527/a_36_216# 0.01fF
C53660 INVX1_LOC_21/A NOR2X1_LOC_748/A 0.03fF
C53661 INVX1_LOC_50/A INVX1_LOC_178/A 0.03fF
C53662 D_INPUT_1 NOR2X1_LOC_652/Y 0.34fF
C53663 INVX1_LOC_132/A INVX1_LOC_63/A 0.16fF
C53664 INVX1_LOC_227/A INVX1_LOC_12/Y 0.29fF
C53665 INVX1_LOC_90/A INVX1_LOC_20/A 3.60fF
C53666 INVX1_LOC_34/A INVX1_LOC_3/A 0.10fF
C53667 INVX1_LOC_179/Y NOR2X1_LOC_640/Y 0.02fF
C53668 NAND2X1_LOC_640/Y INVX1_LOC_63/A 0.00fF
C53669 NAND2X1_LOC_860/A NOR2X1_LOC_791/Y 0.02fF
C53670 NOR2X1_LOC_589/A INVX1_LOC_38/A 0.07fF
C53671 INVX1_LOC_144/Y INVX1_LOC_92/A 0.09fF
C53672 INVX1_LOC_45/A D_INPUT_5 0.01fF
C53673 NOR2X1_LOC_577/Y INVX1_LOC_264/A 0.01fF
C53674 NAND2X1_LOC_359/Y NOR2X1_LOC_240/A 0.03fF
C53675 NOR2X1_LOC_775/Y INVX1_LOC_176/A 0.01fF
C53676 NAND2X1_LOC_372/a_36_24# INVX1_LOC_307/A 0.01fF
C53677 INVX1_LOC_225/A INVX1_LOC_63/A 0.10fF
C53678 NOR2X1_LOC_68/A INVX1_LOC_3/Y 0.14fF
C53679 NOR2X1_LOC_758/Y INVX1_LOC_19/A 0.01fF
C53680 NOR2X1_LOC_468/Y INVX1_LOC_29/Y 0.11fF
C53681 NOR2X1_LOC_78/B NOR2X1_LOC_461/B 0.03fF
C53682 NOR2X1_LOC_163/A INVX1_LOC_117/A 0.00fF
C53683 NAND2X1_LOC_348/A INVX1_LOC_20/A 0.03fF
C53684 INVX1_LOC_311/A NOR2X1_LOC_486/Y 0.03fF
C53685 NAND2X1_LOC_190/Y INVX1_LOC_29/Y 0.02fF
C53686 NOR2X1_LOC_495/Y INVX1_LOC_42/A 0.02fF
C53687 NAND2X1_LOC_735/B NOR2X1_LOC_630/a_36_216# 0.00fF
C53688 NAND2X1_LOC_114/B NOR2X1_LOC_668/Y 0.11fF
C53689 INVX1_LOC_75/A NOR2X1_LOC_357/Y 0.10fF
C53690 INVX1_LOC_150/Y NOR2X1_LOC_383/B 0.05fF
C53691 NAND2X1_LOC_348/A NOR2X1_LOC_360/A 0.01fF
C53692 NOR2X1_LOC_134/Y NAND2X1_LOC_99/A 0.00fF
C53693 NOR2X1_LOC_716/B INVX1_LOC_168/Y 0.01fF
C53694 NOR2X1_LOC_318/B NOR2X1_LOC_78/A 0.07fF
C53695 INVX1_LOC_89/A NOR2X1_LOC_261/A 0.01fF
C53696 INVX1_LOC_50/A NOR2X1_LOC_816/A 1.35fF
C53697 NAND2X1_LOC_361/Y INVX1_LOC_42/A 0.07fF
C53698 INVX1_LOC_16/A INVX1_LOC_123/Y 0.75fF
C53699 NOR2X1_LOC_315/Y NAND2X1_LOC_63/Y 0.03fF
C53700 INVX1_LOC_93/Y INVX1_LOC_98/A 0.03fF
C53701 INVX1_LOC_91/Y VDD 0.41fF
C53702 NAND2X1_LOC_116/A NOR2X1_LOC_340/A 0.03fF
C53703 NOR2X1_LOC_91/A INVX1_LOC_141/Y 0.09fF
C53704 NOR2X1_LOC_329/B NAND2X1_LOC_848/A 0.10fF
C53705 INVX1_LOC_93/Y NOR2X1_LOC_78/A 0.07fF
C53706 INVX1_LOC_75/A NOR2X1_LOC_34/a_36_216# 0.00fF
C53707 INVX1_LOC_96/A NOR2X1_LOC_601/Y 0.01fF
C53708 NOR2X1_LOC_337/Y INVX1_LOC_247/A 0.02fF
C53709 INVX1_LOC_279/A NOR2X1_LOC_600/a_36_216# 0.00fF
C53710 NOR2X1_LOC_765/a_36_216# NAND2X1_LOC_175/Y 0.01fF
C53711 NOR2X1_LOC_91/A INVX1_LOC_312/Y 0.10fF
C53712 INVX1_LOC_72/A INVX1_LOC_26/A 0.01fF
C53713 INVX1_LOC_30/A NAND2X1_LOC_286/B 0.01fF
C53714 NOR2X1_LOC_552/A INVX1_LOC_65/A 0.06fF
C53715 INVX1_LOC_131/A NOR2X1_LOC_536/A 0.02fF
C53716 INVX1_LOC_35/A NOR2X1_LOC_250/Y 0.04fF
C53717 NAND2X1_LOC_799/Y INVX1_LOC_42/A 0.01fF
C53718 NOR2X1_LOC_45/B NOR2X1_LOC_56/Y 0.14fF
C53719 NOR2X1_LOC_516/B NOR2X1_LOC_814/A 0.10fF
C53720 INVX1_LOC_25/Y NAND2X1_LOC_489/Y 0.19fF
C53721 NAND2X1_LOC_858/B NOR2X1_LOC_111/A 0.04fF
C53722 INVX1_LOC_285/Y INVX1_LOC_139/Y 0.13fF
C53723 NOR2X1_LOC_744/a_36_216# NAND2X1_LOC_175/Y 0.01fF
C53724 INVX1_LOC_75/A INVX1_LOC_66/Y 0.00fF
C53725 NOR2X1_LOC_315/Y NAND2X1_LOC_455/B 0.11fF
C53726 NOR2X1_LOC_561/Y NOR2X1_LOC_697/Y 0.20fF
C53727 INVX1_LOC_96/Y NOR2X1_LOC_89/A 0.01fF
C53728 INVX1_LOC_255/Y NOR2X1_LOC_820/B 0.00fF
C53729 INPUT_3 NOR2X1_LOC_392/Y 2.94fF
C53730 INVX1_LOC_155/Y NOR2X1_LOC_609/Y 0.01fF
C53731 INPUT_0 NOR2X1_LOC_536/A 0.28fF
C53732 INVX1_LOC_77/A NAND2X1_LOC_72/B 0.05fF
C53733 NOR2X1_LOC_372/Y NAND2X1_LOC_464/B 0.06fF
C53734 NAND2X1_LOC_569/B NOR2X1_LOC_530/Y 0.31fF
C53735 NOR2X1_LOC_45/B INVX1_LOC_146/Y 0.29fF
C53736 NOR2X1_LOC_433/A INVX1_LOC_273/A 0.12fF
C53737 NOR2X1_LOC_124/A INVX1_LOC_74/A 0.06fF
C53738 INVX1_LOC_136/A INVX1_LOC_57/A 3.03fF
C53739 INVX1_LOC_161/Y NOR2X1_LOC_674/a_36_216# 0.01fF
C53740 INVX1_LOC_277/A NOR2X1_LOC_598/B 0.07fF
C53741 NOR2X1_LOC_45/B VDD 0.75fF
C53742 NAND2X1_LOC_860/A INVX1_LOC_30/A 0.10fF
C53743 NOR2X1_LOC_392/B INVX1_LOC_4/A 0.10fF
C53744 NAND2X1_LOC_361/Y INVX1_LOC_78/A 0.07fF
C53745 INVX1_LOC_34/A NAND2X1_LOC_470/B 0.03fF
C53746 INVX1_LOC_58/A NOR2X1_LOC_68/A 0.06fF
C53747 NAND2X1_LOC_472/Y INVX1_LOC_91/A 0.07fF
C53748 NOR2X1_LOC_808/A NOR2X1_LOC_812/A 0.05fF
C53749 INVX1_LOC_178/A NAND2X1_LOC_227/Y 0.20fF
C53750 NAND2X1_LOC_805/a_36_24# NOR2X1_LOC_652/Y 0.01fF
C53751 INVX1_LOC_39/A INVX1_LOC_293/A 0.00fF
C53752 NOR2X1_LOC_322/Y INVX1_LOC_92/A 0.08fF
C53753 INVX1_LOC_268/A INVX1_LOC_109/Y 0.02fF
C53754 D_INPUT_0 NOR2X1_LOC_691/B 4.64fF
C53755 INVX1_LOC_16/A INVX1_LOC_102/A 0.07fF
C53756 NAND2X1_LOC_799/Y INVX1_LOC_78/A 0.01fF
C53757 VDD INVX1_LOC_247/A -0.00fF
C53758 INVX1_LOC_13/A NAND2X1_LOC_291/B 2.10fF
C53759 INVX1_LOC_199/Y VDD 0.53fF
C53760 INVX1_LOC_224/A NOR2X1_LOC_15/Y 0.49fF
C53761 NOR2X1_LOC_546/B INVX1_LOC_23/A 0.01fF
C53762 NOR2X1_LOC_596/A INVX1_LOC_29/Y 0.02fF
C53763 NOR2X1_LOC_163/Y INVX1_LOC_107/Y 0.22fF
C53764 NOR2X1_LOC_52/B INVX1_LOC_273/A 0.00fF
C53765 INPUT_0 NAND2X1_LOC_93/B 0.10fF
C53766 INVX1_LOC_11/A NOR2X1_LOC_15/Y 0.23fF
C53767 D_INPUT_1 NOR2X1_LOC_403/B 0.01fF
C53768 D_INPUT_1 D_INPUT_2 0.03fF
C53769 NOR2X1_LOC_665/A INVX1_LOC_290/Y 0.02fF
C53770 NAND2X1_LOC_649/B NOR2X1_LOC_536/A 0.05fF
C53771 INVX1_LOC_30/Y NOR2X1_LOC_159/a_36_216# 0.00fF
C53772 INVX1_LOC_25/Y INVX1_LOC_32/A 0.03fF
C53773 NAND2X1_LOC_329/a_36_24# INVX1_LOC_9/A 0.00fF
C53774 NAND2X1_LOC_807/Y NOR2X1_LOC_661/a_36_216# 0.01fF
C53775 NOR2X1_LOC_91/Y NOR2X1_LOC_109/Y 0.09fF
C53776 INVX1_LOC_92/Y INVX1_LOC_92/A 0.09fF
C53777 NAND2X1_LOC_231/Y NAND2X1_LOC_470/B 0.10fF
C53778 INVX1_LOC_91/A NAND2X1_LOC_637/Y 0.04fF
C53779 INVX1_LOC_275/A INVX1_LOC_23/A 0.00fF
C53780 NAND2X1_LOC_158/a_36_24# NOR2X1_LOC_467/A 0.01fF
C53781 INVX1_LOC_41/Y NAND2X1_LOC_790/a_36_24# 0.00fF
C53782 NOR2X1_LOC_99/B NOR2X1_LOC_67/a_36_216# 0.01fF
C53783 NOR2X1_LOC_209/Y NOR2X1_LOC_307/Y 0.01fF
C53784 NAND2X1_LOC_349/B INVX1_LOC_32/A 0.19fF
C53785 NOR2X1_LOC_355/B INVX1_LOC_92/A 0.06fF
C53786 NOR2X1_LOC_83/Y NAND2X1_LOC_572/B 0.11fF
C53787 INVX1_LOC_27/A INVX1_LOC_122/Y 0.09fF
C53788 NOR2X1_LOC_537/Y INVX1_LOC_26/A 0.03fF
C53789 INPUT_0 NOR2X1_LOC_649/B 0.20fF
C53790 NOR2X1_LOC_367/a_36_216# INVX1_LOC_109/Y 0.01fF
C53791 NOR2X1_LOC_538/Y INVX1_LOC_26/Y 0.02fF
C53792 NAND2X1_LOC_849/B INVX1_LOC_20/A 0.13fF
C53793 INVX1_LOC_25/A INVX1_LOC_8/A 0.03fF
C53794 NOR2X1_LOC_295/Y INVX1_LOC_29/Y 0.02fF
C53795 NAND2X1_LOC_338/B INVX1_LOC_26/A 0.36fF
C53796 NOR2X1_LOC_631/B INVX1_LOC_9/A 0.07fF
C53797 INPUT_0 INVX1_LOC_3/A 0.11fF
C53798 INVX1_LOC_38/A INVX1_LOC_20/A 0.10fF
C53799 VDD INVX1_LOC_281/A 0.00fF
C53800 INVX1_LOC_304/A NOR2X1_LOC_177/a_36_216# 0.02fF
C53801 INVX1_LOC_5/A INVX1_LOC_105/A 0.14fF
C53802 NOR2X1_LOC_251/Y NOR2X1_LOC_278/Y 0.16fF
C53803 INVX1_LOC_22/A NOR2X1_LOC_158/Y 0.03fF
C53804 NOR2X1_LOC_666/A INVX1_LOC_72/A 0.08fF
C53805 VDD INVX1_LOC_299/Y 0.41fF
C53806 INVX1_LOC_314/Y INVX1_LOC_50/Y 0.05fF
C53807 NAND2X1_LOC_391/Y INVX1_LOC_24/A 0.03fF
C53808 INVX1_LOC_290/A NOR2X1_LOC_158/a_36_216# 0.01fF
C53809 NAND2X1_LOC_463/B INVX1_LOC_240/Y 0.00fF
C53810 NOR2X1_LOC_553/B NOR2X1_LOC_334/Y 0.02fF
C53811 INVX1_LOC_48/A NOR2X1_LOC_673/A 0.01fF
C53812 VDD NOR2X1_LOC_378/Y 0.23fF
C53813 INVX1_LOC_28/A INVX1_LOC_102/A 0.07fF
C53814 NAND2X1_LOC_773/Y NAND2X1_LOC_364/A 0.10fF
C53815 INVX1_LOC_22/A NOR2X1_LOC_25/Y 0.03fF
C53816 VDD NOR2X1_LOC_499/B 0.08fF
C53817 INVX1_LOC_36/A INVX1_LOC_73/Y 0.01fF
C53818 NOR2X1_LOC_168/B INVX1_LOC_23/A 0.09fF
C53819 NOR2X1_LOC_590/A NOR2X1_LOC_160/B 0.14fF
C53820 NAND2X1_LOC_374/Y NAND2X1_LOC_464/B 0.08fF
C53821 NOR2X1_LOC_598/B NOR2X1_LOC_87/B 0.09fF
C53822 NOR2X1_LOC_358/a_36_216# NAND2X1_LOC_469/B 0.00fF
C53823 NAND2X1_LOC_114/B INVX1_LOC_31/A 0.02fF
C53824 INVX1_LOC_37/A INVX1_LOC_9/A 0.38fF
C53825 INVX1_LOC_73/A INVX1_LOC_12/A 0.02fF
C53826 NOR2X1_LOC_51/A INVX1_LOC_20/A 0.00fF
C53827 NAND2X1_LOC_319/A INVX1_LOC_78/A 0.11fF
C53828 INVX1_LOC_50/A NOR2X1_LOC_773/Y 0.16fF
C53829 INVX1_LOC_135/A INVX1_LOC_4/Y 0.07fF
C53830 NOR2X1_LOC_268/a_36_216# INVX1_LOC_88/A 0.00fF
C53831 NOR2X1_LOC_188/A INVX1_LOC_29/A 1.41fF
C53832 INVX1_LOC_228/A INVX1_LOC_1/A 0.32fF
C53833 INVX1_LOC_90/A INVX1_LOC_4/A 0.21fF
C53834 INVX1_LOC_31/A INVX1_LOC_141/Y 0.03fF
C53835 INVX1_LOC_144/Y INVX1_LOC_53/A 0.03fF
C53836 INVX1_LOC_45/Y INVX1_LOC_88/A 0.05fF
C53837 NOR2X1_LOC_103/Y NOR2X1_LOC_360/Y 0.07fF
C53838 NOR2X1_LOC_389/B INVX1_LOC_4/A 0.10fF
C53839 NOR2X1_LOC_563/a_36_216# NOR2X1_LOC_383/B 0.00fF
C53840 INVX1_LOC_16/A INVX1_LOC_296/Y 0.03fF
C53841 VDD NOR2X1_LOC_676/Y 0.12fF
C53842 NOR2X1_LOC_90/a_36_216# INVX1_LOC_61/Y 0.01fF
C53843 NOR2X1_LOC_181/Y INVX1_LOC_50/Y 0.09fF
C53844 NOR2X1_LOC_68/A INVX1_LOC_215/Y 0.03fF
C53845 NOR2X1_LOC_294/Y INVX1_LOC_31/A 0.34fF
C53846 NAND2X1_LOC_386/a_36_24# INVX1_LOC_174/A 0.01fF
C53847 NOR2X1_LOC_15/Y NOR2X1_LOC_433/A 0.13fF
C53848 VDD NOR2X1_LOC_862/B 2.25fF
C53849 INVX1_LOC_91/A NAND2X1_LOC_773/B 0.06fF
C53850 NOR2X1_LOC_15/Y NOR2X1_LOC_474/A 0.03fF
C53851 NOR2X1_LOC_208/Y INVX1_LOC_73/Y 0.01fF
C53852 NAND2X1_LOC_349/a_36_24# INVX1_LOC_23/A 0.00fF
C53853 INVX1_LOC_69/Y INVX1_LOC_99/A 0.00fF
C53854 INVX1_LOC_5/A NOR2X1_LOC_720/a_36_216# 0.02fF
C53855 NAND2X1_LOC_642/Y INVX1_LOC_63/A 0.21fF
C53856 INPUT_5 INVX1_LOC_296/A 0.14fF
C53857 NOR2X1_LOC_15/Y NOR2X1_LOC_593/Y 0.07fF
C53858 INVX1_LOC_11/A NOR2X1_LOC_860/B 0.07fF
C53859 INVX1_LOC_75/A INVX1_LOC_32/A 0.10fF
C53860 NOR2X1_LOC_65/B NAND2X1_LOC_660/a_36_24# 0.00fF
C53861 NAND2X1_LOC_348/A INVX1_LOC_4/A 0.03fF
C53862 INVX1_LOC_120/A NOR2X1_LOC_342/B 0.12fF
C53863 INVX1_LOC_1/A INVX1_LOC_8/A 0.10fF
C53864 INVX1_LOC_21/A NOR2X1_LOC_493/B 0.19fF
C53865 NOR2X1_LOC_778/B INVX1_LOC_50/Y 0.03fF
C53866 INVX1_LOC_281/Y INVX1_LOC_92/A 0.01fF
C53867 NOR2X1_LOC_205/Y NOR2X1_LOC_388/Y 0.06fF
C53868 INVX1_LOC_57/Y NOR2X1_LOC_487/a_36_216# 0.13fF
C53869 INPUT_1 NAND2X1_LOC_99/A 0.08fF
C53870 INVX1_LOC_45/A NOR2X1_LOC_360/Y 0.01fF
C53871 NAND2X1_LOC_656/Y INVX1_LOC_23/A 0.17fF
C53872 NOR2X1_LOC_332/A NOR2X1_LOC_105/Y 0.05fF
C53873 INVX1_LOC_200/A NAND2X1_LOC_833/Y 0.07fF
C53874 INVX1_LOC_17/A NOR2X1_LOC_690/A 0.00fF
C53875 NOR2X1_LOC_15/Y NOR2X1_LOC_52/B 0.18fF
C53876 NOR2X1_LOC_360/Y NOR2X1_LOC_568/A 0.01fF
C53877 INPUT_3 NOR2X1_LOC_554/a_36_216# 0.00fF
C53878 NOR2X1_LOC_70/a_36_216# NOR2X1_LOC_25/Y 0.00fF
C53879 INVX1_LOC_269/A INVX1_LOC_104/A 0.09fF
C53880 INVX1_LOC_200/Y NAND2X1_LOC_861/Y 0.01fF
C53881 NAND2X1_LOC_240/a_36_24# NOR2X1_LOC_536/A 0.00fF
C53882 NOR2X1_LOC_82/A NAND2X1_LOC_139/A 0.02fF
C53883 NOR2X1_LOC_180/a_36_216# INVX1_LOC_271/Y 0.01fF
C53884 NOR2X1_LOC_276/B INVX1_LOC_72/A 0.03fF
C53885 INVX1_LOC_256/A INVX1_LOC_34/A 0.03fF
C53886 NAND2X1_LOC_326/A NAND2X1_LOC_660/A 1.24fF
C53887 INVX1_LOC_159/A NOR2X1_LOC_52/Y 0.00fF
C53888 INVX1_LOC_174/A INVX1_LOC_33/A 0.06fF
C53889 NAND2X1_LOC_346/a_36_24# NOR2X1_LOC_709/A 0.00fF
C53890 NOR2X1_LOC_657/Y NOR2X1_LOC_759/Y 0.02fF
C53891 NOR2X1_LOC_635/A INVX1_LOC_11/A 0.03fF
C53892 INVX1_LOC_136/A NOR2X1_LOC_220/a_36_216# 0.01fF
C53893 NOR2X1_LOC_186/Y INVX1_LOC_1/Y 0.04fF
C53894 INVX1_LOC_303/A NOR2X1_LOC_641/B 0.03fF
C53895 NOR2X1_LOC_124/A NAND2X1_LOC_254/Y 0.05fF
C53896 INVX1_LOC_24/A NOR2X1_LOC_703/B 0.03fF
C53897 NOR2X1_LOC_503/Y NAND2X1_LOC_799/Y 0.02fF
C53898 INVX1_LOC_35/A D_INPUT_0 6.11fF
C53899 NAND2X1_LOC_357/B NAND2X1_LOC_793/Y 0.16fF
C53900 INVX1_LOC_132/A NOR2X1_LOC_688/Y 0.12fF
C53901 NOR2X1_LOC_67/A NAND2X1_LOC_579/A 0.28fF
C53902 NOR2X1_LOC_669/Y INVX1_LOC_248/A 0.01fF
C53903 NOR2X1_LOC_392/B INVX1_LOC_43/Y 0.39fF
C53904 NOR2X1_LOC_473/B INVX1_LOC_53/A 0.10fF
C53905 INVX1_LOC_50/A INVX1_LOC_140/A 0.03fF
C53906 INVX1_LOC_298/Y NOR2X1_LOC_188/A 0.02fF
C53907 INVX1_LOC_64/A INVX1_LOC_97/A 0.08fF
C53908 NOR2X1_LOC_609/A INVX1_LOC_94/A 0.62fF
C53909 VDD NOR2X1_LOC_1/Y -0.00fF
C53910 NOR2X1_LOC_360/Y INVX1_LOC_71/A 0.01fF
C53911 NOR2X1_LOC_546/A NOR2X1_LOC_713/B 0.13fF
C53912 NAND2X1_LOC_725/Y NAND2X1_LOC_560/A 1.96fF
C53913 NAND2X1_LOC_785/B NAND2X1_LOC_833/a_36_24# 0.01fF
C53914 NAND2X1_LOC_149/Y NAND2X1_LOC_662/Y 0.14fF
C53915 INVX1_LOC_63/A NOR2X1_LOC_271/Y 0.03fF
C53916 INVX1_LOC_64/A INVX1_LOC_90/A 0.18fF
C53917 NOR2X1_LOC_272/Y INVX1_LOC_279/A 0.07fF
C53918 NAND2X1_LOC_655/A INVX1_LOC_21/Y 0.02fF
C53919 INVX1_LOC_224/A INVX1_LOC_226/A 0.47fF
C53920 NOR2X1_LOC_237/Y NOR2X1_LOC_91/Y 0.01fF
C53921 NAND2X1_LOC_96/A NAND2X1_LOC_63/Y 0.10fF
C53922 NAND2X1_LOC_198/B INVX1_LOC_77/A 0.10fF
C53923 NOR2X1_LOC_382/Y NOR2X1_LOC_84/A 0.03fF
C53924 NOR2X1_LOC_813/Y NAND2X1_LOC_81/B 0.02fF
C53925 INVX1_LOC_144/A NOR2X1_LOC_654/A 0.32fF
C53926 NOR2X1_LOC_298/a_36_216# NAND2X1_LOC_463/B 0.00fF
C53927 NOR2X1_LOC_357/Y INVX1_LOC_283/A 0.09fF
C53928 NOR2X1_LOC_552/A INVX1_LOC_4/Y 0.02fF
C53929 INVX1_LOC_13/Y NOR2X1_LOC_71/Y 0.53fF
C53930 INVX1_LOC_11/A INVX1_LOC_226/A 0.02fF
C53931 INVX1_LOC_62/A NOR2X1_LOC_849/A 0.06fF
C53932 INVX1_LOC_11/A NAND2X1_LOC_840/B 0.00fF
C53933 NOR2X1_LOC_78/A INVX1_LOC_87/A 0.03fF
C53934 NOR2X1_LOC_454/Y NOR2X1_LOC_781/B 0.02fF
C53935 INVX1_LOC_21/A NOR2X1_LOC_110/a_36_216# 0.00fF
C53936 NAND2X1_LOC_391/Y NOR2X1_LOC_130/A 0.09fF
C53937 NOR2X1_LOC_322/Y INVX1_LOC_53/A 0.24fF
C53938 NOR2X1_LOC_205/Y NAND2X1_LOC_479/Y 0.08fF
C53939 NOR2X1_LOC_824/A NOR2X1_LOC_525/Y 0.05fF
C53940 NOR2X1_LOC_230/Y INVX1_LOC_266/Y 0.01fF
C53941 NOR2X1_LOC_566/a_36_216# INVX1_LOC_4/Y 0.01fF
C53942 INVX1_LOC_21/A INVX1_LOC_89/A 7.29fF
C53943 NOR2X1_LOC_667/A NAND2X1_LOC_711/Y 0.19fF
C53944 INVX1_LOC_32/A NAND2X1_LOC_453/A 0.07fF
C53945 INVX1_LOC_119/A NAND2X1_LOC_354/Y 0.01fF
C53946 NOR2X1_LOC_309/Y NOR2X1_LOC_91/Y 0.03fF
C53947 INVX1_LOC_64/A NAND2X1_LOC_348/A 0.25fF
C53948 INVX1_LOC_91/A NOR2X1_LOC_481/a_36_216# 0.00fF
C53949 NOR2X1_LOC_160/B NOR2X1_LOC_82/Y 0.03fF
C53950 INVX1_LOC_45/A NAND2X1_LOC_451/Y 0.07fF
C53951 NOR2X1_LOC_96/a_36_216# NOR2X1_LOC_671/Y 0.00fF
C53952 INVX1_LOC_211/Y INVX1_LOC_22/A 0.01fF
C53953 INVX1_LOC_21/A NAND2X1_LOC_508/A 0.00fF
C53954 NOR2X1_LOC_346/A INVX1_LOC_230/A 0.01fF
C53955 INVX1_LOC_78/Y INVX1_LOC_23/A 0.03fF
C53956 INVX1_LOC_62/Y INVX1_LOC_60/Y 0.23fF
C53957 NOR2X1_LOC_590/A NOR2X1_LOC_516/B 0.07fF
C53958 INVX1_LOC_103/A NOR2X1_LOC_366/Y 0.02fF
C53959 NAND2X1_LOC_223/A INVX1_LOC_20/A 0.06fF
C53960 INVX1_LOC_90/A NAND2X1_LOC_704/a_36_24# 0.00fF
C53961 INVX1_LOC_22/Y NOR2X1_LOC_516/B 0.03fF
C53962 NOR2X1_LOC_503/Y NAND2X1_LOC_319/A 0.03fF
C53963 INVX1_LOC_314/Y NOR2X1_LOC_6/B 0.39fF
C53964 VDD NOR2X1_LOC_685/B -0.00fF
C53965 INVX1_LOC_37/A INVX1_LOC_274/Y 0.02fF
C53966 VDD NOR2X1_LOC_465/Y 0.31fF
C53967 NOR2X1_LOC_355/B INVX1_LOC_53/A 0.01fF
C53968 NOR2X1_LOC_808/A NOR2X1_LOC_324/Y 0.02fF
C53969 INVX1_LOC_227/A NOR2X1_LOC_160/B 0.07fF
C53970 NOR2X1_LOC_114/Y INVX1_LOC_54/A 0.02fF
C53971 INVX1_LOC_223/A INVX1_LOC_16/A 0.03fF
C53972 INVX1_LOC_112/A INVX1_LOC_112/Y 0.09fF
C53973 INVX1_LOC_59/Y INVX1_LOC_112/Y 0.01fF
C53974 NOR2X1_LOC_235/Y INVX1_LOC_284/A 0.01fF
C53975 NAND2X1_LOC_214/B NOR2X1_LOC_391/Y -0.04fF
C53976 NOR2X1_LOC_226/A NAND2X1_LOC_656/A 0.05fF
C53977 NOR2X1_LOC_798/A NOR2X1_LOC_292/Y 0.00fF
C53978 NOR2X1_LOC_793/A NOR2X1_LOC_703/A 0.03fF
C53979 NOR2X1_LOC_433/A INVX1_LOC_96/Y 0.72fF
C53980 NOR2X1_LOC_355/A NOR2X1_LOC_389/A 0.01fF
C53981 INVX1_LOC_304/Y NAND2X1_LOC_833/Y 0.22fF
C53982 INVX1_LOC_236/A NOR2X1_LOC_577/Y 0.12fF
C53983 NOR2X1_LOC_520/A NOR2X1_LOC_350/A 0.12fF
C53984 INVX1_LOC_280/A INVX1_LOC_4/Y 0.01fF
C53985 NOR2X1_LOC_593/Y INVX1_LOC_96/Y 0.03fF
C53986 NAND2X1_LOC_112/Y NAND2X1_LOC_514/Y 0.00fF
C53987 INVX1_LOC_90/A INVX1_LOC_43/Y 0.00fF
C53988 NOR2X1_LOC_205/Y NOR2X1_LOC_202/Y 0.04fF
C53989 NAND2X1_LOC_342/Y INVX1_LOC_155/A 0.14fF
C53990 NOR2X1_LOC_222/Y INVX1_LOC_49/A 0.05fF
C53991 NOR2X1_LOC_243/B NAND2X1_LOC_206/B 0.15fF
C53992 NAND2X1_LOC_72/B INVX1_LOC_9/A 0.03fF
C53993 NAND2X1_LOC_448/a_36_24# INVX1_LOC_296/Y 0.01fF
C53994 NAND2X1_LOC_227/Y INVX1_LOC_140/A 0.13fF
C53995 NOR2X1_LOC_219/Y INVX1_LOC_77/A 0.98fF
C53996 NAND2X1_LOC_30/Y D_INPUT_4 0.46fF
C53997 NOR2X1_LOC_186/Y NOR2X1_LOC_318/B 0.00fF
C53998 NOR2X1_LOC_510/Y NOR2X1_LOC_45/B 0.10fF
C53999 NAND2X1_LOC_218/B INVX1_LOC_13/A 0.09fF
C54000 INVX1_LOC_77/A INVX1_LOC_53/Y 0.63fF
C54001 NAND2X1_LOC_577/A INPUT_1 0.01fF
C54002 NOR2X1_LOC_53/Y NOR2X1_LOC_56/Y 0.09fF
C54003 NOR2X1_LOC_52/B INVX1_LOC_96/Y 0.18fF
C54004 NOR2X1_LOC_795/Y INVX1_LOC_177/A 0.00fF
C54005 INVX1_LOC_30/Y INVX1_LOC_314/Y 0.88fF
C54006 INVX1_LOC_30/A INVX1_LOC_85/Y 0.03fF
C54007 INVX1_LOC_33/A NOR2X1_LOC_131/Y 0.03fF
C54008 INVX1_LOC_132/A INVX1_LOC_1/Y 0.07fF
C54009 INVX1_LOC_11/A NAND2X1_LOC_2/a_36_24# 0.00fF
C54010 NAND2X1_LOC_121/a_36_24# INVX1_LOC_6/A 0.00fF
C54011 INVX1_LOC_2/A NOR2X1_LOC_423/Y 0.01fF
C54012 INVX1_LOC_19/A INVX1_LOC_69/A 0.04fF
C54013 INVX1_LOC_119/A INVX1_LOC_214/A 0.31fF
C54014 INPUT_3 INVX1_LOC_75/A 0.69fF
C54015 INVX1_LOC_256/A INPUT_0 0.00fF
C54016 NOR2X1_LOC_773/a_36_216# NOR2X1_LOC_773/Y 0.02fF
C54017 NOR2X1_LOC_590/A NOR2X1_LOC_706/A 0.00fF
C54018 INVX1_LOC_149/A NOR2X1_LOC_537/Y 0.02fF
C54019 INVX1_LOC_118/A NAND2X1_LOC_99/A 0.76fF
C54020 NOR2X1_LOC_89/A INVX1_LOC_49/Y 0.03fF
C54021 INVX1_LOC_223/A INVX1_LOC_28/A 0.40fF
C54022 VDD NOR2X1_LOC_53/Y 0.20fF
C54023 NOR2X1_LOC_589/A INVX1_LOC_33/A 0.13fF
C54024 INVX1_LOC_145/Y INVX1_LOC_77/A 0.03fF
C54025 INVX1_LOC_240/Y INVX1_LOC_42/A 0.22fF
C54026 NAND2X1_LOC_112/Y NAND2X1_LOC_332/Y 0.02fF
C54027 INVX1_LOC_45/A NOR2X1_LOC_567/B 0.08fF
C54028 INVX1_LOC_35/A NOR2X1_LOC_859/Y 0.00fF
C54029 INVX1_LOC_225/A INVX1_LOC_1/Y 0.23fF
C54030 INVX1_LOC_2/A NOR2X1_LOC_222/Y 0.06fF
C54031 NAND2X1_LOC_773/Y NOR2X1_LOC_405/A 0.00fF
C54032 INVX1_LOC_18/A NOR2X1_LOC_564/Y 0.03fF
C54033 INVX1_LOC_85/A INVX1_LOC_16/A 0.03fF
C54034 INVX1_LOC_41/A NOR2X1_LOC_391/A 0.77fF
C54035 INVX1_LOC_124/A INVX1_LOC_53/Y 0.02fF
C54036 NOR2X1_LOC_15/Y NOR2X1_LOC_601/Y 0.12fF
C54037 NOR2X1_LOC_350/A INVX1_LOC_65/Y 0.42fF
C54038 NOR2X1_LOC_82/A NOR2X1_LOC_78/A 0.08fF
C54039 INVX1_LOC_2/A NOR2X1_LOC_269/a_36_216# 0.00fF
C54040 NOR2X1_LOC_736/Y NOR2X1_LOC_596/A 2.75fF
C54041 INVX1_LOC_64/A INVX1_LOC_38/A 0.21fF
C54042 NAND2X1_LOC_454/Y NAND2X1_LOC_475/Y 0.01fF
C54043 NOR2X1_LOC_454/Y NOR2X1_LOC_585/Y 0.03fF
C54044 NOR2X1_LOC_613/Y VDD 0.18fF
C54045 NOR2X1_LOC_843/A INVX1_LOC_135/A 0.01fF
C54046 INVX1_LOC_292/A INVX1_LOC_186/A 0.46fF
C54047 NOR2X1_LOC_468/Y INVX1_LOC_126/A 0.21fF
C54048 INVX1_LOC_55/Y NOR2X1_LOC_577/Y 0.17fF
C54049 NOR2X1_LOC_218/Y NOR2X1_LOC_222/Y 0.02fF
C54050 NOR2X1_LOC_795/Y NOR2X1_LOC_785/Y 0.16fF
C54051 INVX1_LOC_135/A INVX1_LOC_82/A 0.04fF
C54052 NOR2X1_LOC_516/B NAND2X1_LOC_819/Y 0.05fF
C54053 INVX1_LOC_64/A NOR2X1_LOC_96/Y 0.01fF
C54054 NOR2X1_LOC_807/B NOR2X1_LOC_324/A 0.04fF
C54055 NAND2X1_LOC_483/Y NAND2X1_LOC_866/B 0.07fF
C54056 INVX1_LOC_135/A INVX1_LOC_194/A 0.35fF
C54057 INVX1_LOC_13/A NOR2X1_LOC_346/B 0.07fF
C54058 INVX1_LOC_271/A NAND2X1_LOC_792/a_36_24# 0.00fF
C54059 INVX1_LOC_49/A NOR2X1_LOC_329/B 0.21fF
C54060 INVX1_LOC_120/A NAND2X1_LOC_116/A 0.03fF
C54061 NOR2X1_LOC_454/Y INVX1_LOC_77/Y 0.85fF
C54062 INVX1_LOC_299/A INVX1_LOC_14/Y 0.05fF
C54063 INVX1_LOC_49/A D_INPUT_4 0.03fF
C54064 NAND2X1_LOC_512/a_36_24# NAND2X1_LOC_472/Y 0.00fF
C54065 NAND2X1_LOC_733/Y NAND2X1_LOC_729/B 0.46fF
C54066 NAND2X1_LOC_564/B INVX1_LOC_25/Y 0.22fF
C54067 INVX1_LOC_232/Y INVX1_LOC_234/A 0.24fF
C54068 INVX1_LOC_9/Y NAND2X1_LOC_349/B 0.02fF
C54069 NAND2X1_LOC_363/B NOR2X1_LOC_461/A -0.01fF
C54070 INVX1_LOC_292/A NAND2X1_LOC_447/Y 0.10fF
C54071 NAND2X1_LOC_181/Y INVX1_LOC_10/A 0.01fF
C54072 INVX1_LOC_303/A NOR2X1_LOC_751/A 0.06fF
C54073 INVX1_LOC_55/Y NOR2X1_LOC_348/B 0.03fF
C54074 INVX1_LOC_64/A NAND2X1_LOC_848/Y 0.00fF
C54075 NAND2X1_LOC_9/Y NOR2X1_LOC_461/B 0.09fF
C54076 INVX1_LOC_227/A INVX1_LOC_208/A 0.10fF
C54077 NOR2X1_LOC_550/B NOR2X1_LOC_74/A 0.00fF
C54078 NOR2X1_LOC_798/A NOR2X1_LOC_641/Y 0.02fF
C54079 INVX1_LOC_186/Y NAND2X1_LOC_299/a_36_24# 0.00fF
C54080 INVX1_LOC_155/A INVX1_LOC_67/Y 0.00fF
C54081 INVX1_LOC_13/Y NAND2X1_LOC_243/Y 0.01fF
C54082 NOR2X1_LOC_553/B NOR2X1_LOC_569/Y 0.11fF
C54083 NOR2X1_LOC_174/A NOR2X1_LOC_175/A 0.03fF
C54084 INVX1_LOC_64/A NOR2X1_LOC_697/a_36_216# 0.01fF
C54085 NOR2X1_LOC_716/B NOR2X1_LOC_83/Y 0.27fF
C54086 INVX1_LOC_255/Y INVX1_LOC_80/A 0.03fF
C54087 NAND2X1_LOC_53/Y INVX1_LOC_117/A 0.12fF
C54088 INVX1_LOC_24/A INVX1_LOC_91/A 0.46fF
C54089 INVX1_LOC_270/Y INVX1_LOC_19/A 0.01fF
C54090 INVX1_LOC_2/A NOR2X1_LOC_329/B 0.26fF
C54091 NOR2X1_LOC_92/Y NOR2X1_LOC_629/Y 0.04fF
C54092 NOR2X1_LOC_188/A INVX1_LOC_8/A 0.07fF
C54093 NOR2X1_LOC_757/A NOR2X1_LOC_561/Y 0.04fF
C54094 INVX1_LOC_223/A NOR2X1_LOC_35/Y 0.03fF
C54095 NOR2X1_LOC_219/B INVX1_LOC_6/A 0.01fF
C54096 NOR2X1_LOC_468/Y INVX1_LOC_127/A 0.02fF
C54097 INVX1_LOC_71/A NOR2X1_LOC_269/Y 0.07fF
C54098 NOR2X1_LOC_551/Y NOR2X1_LOC_551/B 0.01fF
C54099 NOR2X1_LOC_548/B INVX1_LOC_8/A 1.95fF
C54100 INVX1_LOC_34/A INVX1_LOC_69/Y 0.03fF
C54101 INVX1_LOC_232/Y NOR2X1_LOC_19/B 0.48fF
C54102 NOR2X1_LOC_226/A NOR2X1_LOC_329/B 0.01fF
C54103 NOR2X1_LOC_598/B NAND2X1_LOC_219/B -0.01fF
C54104 NAND2X1_LOC_467/a_36_24# D_INPUT_5 0.01fF
C54105 NOR2X1_LOC_209/Y NOR2X1_LOC_742/A 0.92fF
C54106 INVX1_LOC_24/A INVX1_LOC_11/Y 0.08fF
C54107 NOR2X1_LOC_565/A INVX1_LOC_37/A 0.01fF
C54108 NOR2X1_LOC_778/Y VDD 0.51fF
C54109 INVX1_LOC_55/Y INVX1_LOC_22/A 12.13fF
C54110 NAND2X1_LOC_358/Y INVX1_LOC_148/Y 0.06fF
C54111 NOR2X1_LOC_19/B INVX1_LOC_197/Y 0.00fF
C54112 INVX1_LOC_50/A INVX1_LOC_42/A 0.91fF
C54113 NOR2X1_LOC_723/Y INVX1_LOC_139/Y 0.01fF
C54114 NOR2X1_LOC_481/A NOR2X1_LOC_318/B 0.05fF
C54115 NAND2X1_LOC_785/A NAND2X1_LOC_858/B 0.00fF
C54116 INVX1_LOC_290/A D_GATE_366 0.07fF
C54117 NOR2X1_LOC_52/Y VDD 0.44fF
C54118 NOR2X1_LOC_343/B NAND2X1_LOC_574/A 0.06fF
C54119 NAND2X1_LOC_543/Y INVX1_LOC_28/A 0.00fF
C54120 NOR2X1_LOC_557/Y INVX1_LOC_91/A 0.04fF
C54121 INPUT_6 INPUT_7 0.04fF
C54122 NOR2X1_LOC_516/B NOR2X1_LOC_703/A 0.03fF
C54123 NOR2X1_LOC_270/Y VDD 0.60fF
C54124 INVX1_LOC_89/A NOR2X1_LOC_565/B 0.05fF
C54125 INVX1_LOC_24/A NOR2X1_LOC_421/Y 0.04fF
C54126 INVX1_LOC_174/A NAND2X1_LOC_459/a_36_24# 0.00fF
C54127 NAND2X1_LOC_656/Y INVX1_LOC_313/A 0.03fF
C54128 INVX1_LOC_48/Y INVX1_LOC_123/Y 0.03fF
C54129 NAND2X1_LOC_359/Y NAND2X1_LOC_348/a_36_24# 0.01fF
C54130 INVX1_LOC_177/Y INVX1_LOC_12/Y 0.10fF
C54131 NOR2X1_LOC_555/a_36_216# INVX1_LOC_121/Y 0.00fF
C54132 NOR2X1_LOC_238/Y NOR2X1_LOC_482/a_36_216# 0.00fF
C54133 NOR2X1_LOC_458/Y INVX1_LOC_247/A -0.01fF
C54134 INVX1_LOC_225/A INVX1_LOC_93/Y 0.01fF
C54135 NOR2X1_LOC_75/Y NOR2X1_LOC_155/A 0.03fF
C54136 NAND2X1_LOC_74/B INVX1_LOC_306/Y 1.04fF
C54137 NAND2X1_LOC_647/B INVX1_LOC_57/A 0.02fF
C54138 INVX1_LOC_33/A INVX1_LOC_20/A 0.03fF
C54139 NOR2X1_LOC_45/Y INVX1_LOC_117/Y 0.03fF
C54140 INVX1_LOC_143/A INVX1_LOC_91/A 0.07fF
C54141 NOR2X1_LOC_360/Y NOR2X1_LOC_331/B 0.09fF
C54142 INVX1_LOC_50/A INVX1_LOC_78/A 0.13fF
C54143 INVX1_LOC_280/Y NOR2X1_LOC_45/B 0.03fF
C54144 INVX1_LOC_149/Y NOR2X1_LOC_35/Y 0.06fF
C54145 INVX1_LOC_128/Y INVX1_LOC_23/A 0.22fF
C54146 INVX1_LOC_96/Y INVX1_LOC_199/A 0.05fF
C54147 NAND2X1_LOC_794/B INVX1_LOC_102/A 0.31fF
C54148 NAND2X1_LOC_198/B INVX1_LOC_9/A 0.03fF
C54149 INVX1_LOC_31/A NOR2X1_LOC_820/a_36_216# 0.01fF
C54150 INVX1_LOC_85/A NOR2X1_LOC_35/Y 0.00fF
C54151 NAND2X1_LOC_738/B NOR2X1_LOC_409/B 0.03fF
C54152 NOR2X1_LOC_817/Y NOR2X1_LOC_820/B 0.01fF
C54153 INVX1_LOC_265/A VDD 0.04fF
C54154 NAND2X1_LOC_778/Y NAND2X1_LOC_254/Y 0.01fF
C54155 NAND2X1_LOC_162/A NOR2X1_LOC_45/B 0.01fF
C54156 INVX1_LOC_2/A NOR2X1_LOC_69/A 0.01fF
C54157 INVX1_LOC_224/Y INVX1_LOC_26/A 0.23fF
C54158 INVX1_LOC_138/Y NOR2X1_LOC_38/B 0.04fF
C54159 INVX1_LOC_89/A NAND2X1_LOC_51/B 0.04fF
C54160 NOR2X1_LOC_180/Y VDD 0.12fF
C54161 NAND2X1_LOC_656/Y INVX1_LOC_6/A 0.07fF
C54162 NOR2X1_LOC_599/A NAND2X1_LOC_809/a_36_24# 0.00fF
C54163 NOR2X1_LOC_224/Y INVX1_LOC_78/A 0.01fF
C54164 NOR2X1_LOC_65/B INVX1_LOC_50/A 0.02fF
C54165 NOR2X1_LOC_717/B NOR2X1_LOC_730/B 0.01fF
C54166 INVX1_LOC_30/Y NOR2X1_LOC_557/A 0.02fF
C54167 INVX1_LOC_11/A INVX1_LOC_49/Y 0.03fF
C54168 INVX1_LOC_251/Y NAND2X1_LOC_267/B 0.06fF
C54169 NOR2X1_LOC_703/B NOR2X1_LOC_197/B 0.03fF
C54170 INVX1_LOC_104/A INVX1_LOC_12/Y 0.10fF
C54171 NAND2X1_LOC_629/Y INVX1_LOC_37/A 0.03fF
C54172 NAND2X1_LOC_652/a_36_24# NOR2X1_LOC_331/B 0.00fF
C54173 INVX1_LOC_89/A INVX1_LOC_311/A 0.07fF
C54174 INVX1_LOC_136/A NAND2X1_LOC_243/a_36_24# 0.01fF
C54175 INVX1_LOC_1/Y NAND2X1_LOC_642/Y 0.07fF
C54176 NOR2X1_LOC_15/Y NAND2X1_LOC_254/Y 0.03fF
C54177 NAND2X1_LOC_811/Y NOR2X1_LOC_536/A 0.00fF
C54178 INVX1_LOC_23/A NOR2X1_LOC_727/B 0.03fF
C54179 INVX1_LOC_64/A INVX1_LOC_18/Y 0.08fF
C54180 NOR2X1_LOC_401/Y VDD 0.24fF
C54181 NOR2X1_LOC_593/Y NAND2X1_LOC_204/a_36_24# 0.00fF
C54182 INVX1_LOC_224/Y NAND2X1_LOC_564/A 0.06fF
C54183 INVX1_LOC_310/Y INVX1_LOC_9/A 0.03fF
C54184 INVX1_LOC_210/Y NOR2X1_LOC_814/A 0.31fF
C54185 INVX1_LOC_40/A INVX1_LOC_20/A 2.16fF
C54186 NAND2X1_LOC_783/A INVX1_LOC_91/A 0.10fF
C54187 NOR2X1_LOC_272/Y NOR2X1_LOC_38/B 0.01fF
C54188 INVX1_LOC_243/A INVX1_LOC_37/A 0.00fF
C54189 NOR2X1_LOC_355/A NAND2X1_LOC_498/a_36_24# 0.00fF
C54190 NAND2X1_LOC_800/a_36_24# INVX1_LOC_16/A 0.01fF
C54191 NAND2X1_LOC_759/a_36_24# NOR2X1_LOC_536/A 0.00fF
C54192 NOR2X1_LOC_238/Y NOR2X1_LOC_88/Y 0.03fF
C54193 NOR2X1_LOC_130/A INVX1_LOC_91/A 0.10fF
C54194 INVX1_LOC_184/Y NOR2X1_LOC_862/B 0.11fF
C54195 NOR2X1_LOC_186/Y INVX1_LOC_87/A 0.03fF
C54196 NOR2X1_LOC_352/Y NAND2X1_LOC_472/Y 0.01fF
C54197 NAND2X1_LOC_860/A NAND2X1_LOC_458/a_36_24# 0.00fF
C54198 NOR2X1_LOC_357/Y INVX1_LOC_22/A 0.07fF
C54199 NOR2X1_LOC_590/A NAND2X1_LOC_207/B 0.03fF
C54200 INVX1_LOC_124/A NOR2X1_LOC_652/a_36_216# 0.03fF
C54201 INVX1_LOC_230/Y INVX1_LOC_284/A 0.34fF
C54202 INVX1_LOC_24/A NOR2X1_LOC_179/Y 0.16fF
C54203 INVX1_LOC_23/A NOR2X1_LOC_717/A 0.03fF
C54204 NOR2X1_LOC_91/Y INVX1_LOC_63/A 0.00fF
C54205 NOR2X1_LOC_78/B INVX1_LOC_281/Y 0.01fF
C54206 NOR2X1_LOC_318/A NOR2X1_LOC_652/Y 0.16fF
C54207 NOR2X1_LOC_234/a_36_216# NAND2X1_LOC_243/Y 0.00fF
C54208 NOR2X1_LOC_238/Y INVX1_LOC_84/A 0.00fF
C54209 NOR2X1_LOC_151/Y NOR2X1_LOC_730/B 0.04fF
C54210 INVX1_LOC_88/A INVX1_LOC_21/Y 0.04fF
C54211 NOR2X1_LOC_200/a_36_216# INVX1_LOC_54/A 0.00fF
C54212 NOR2X1_LOC_598/B INVX1_LOC_58/Y 0.86fF
C54213 NOR2X1_LOC_233/a_36_216# INVX1_LOC_23/Y 0.00fF
C54214 NAND2X1_LOC_491/a_36_24# INVX1_LOC_9/A 0.00fF
C54215 INVX1_LOC_61/Y INVX1_LOC_42/A 0.14fF
C54216 INVX1_LOC_24/A INVX1_LOC_203/A 0.14fF
C54217 INVX1_LOC_39/A NAND2X1_LOC_99/A 0.01fF
C54218 NAND2X1_LOC_799/Y NAND2X1_LOC_802/Y 0.29fF
C54219 INVX1_LOC_10/A NOR2X1_LOC_314/Y 0.02fF
C54220 INVX1_LOC_70/Y NAND2X1_LOC_850/A 0.14fF
C54221 INVX1_LOC_227/A NAND2X1_LOC_211/Y 0.16fF
C54222 NOR2X1_LOC_643/Y INVX1_LOC_3/A 0.03fF
C54223 NOR2X1_LOC_561/Y INVX1_LOC_37/A 0.02fF
C54224 INVX1_LOC_295/A INVX1_LOC_115/Y 0.03fF
C54225 INVX1_LOC_69/Y INPUT_0 0.26fF
C54226 INVX1_LOC_8/Y NOR2X1_LOC_814/A 0.03fF
C54227 INVX1_LOC_27/A NOR2X1_LOC_72/Y -0.02fF
C54228 INVX1_LOC_89/A NOR2X1_LOC_670/Y 0.01fF
C54229 INVX1_LOC_266/Y NAND2X1_LOC_93/B 0.07fF
C54230 INVX1_LOC_13/Y NAND2X1_LOC_205/A 0.03fF
C54231 NOR2X1_LOC_722/Y NOR2X1_LOC_89/A 0.01fF
C54232 NOR2X1_LOC_268/a_36_216# INVX1_LOC_272/A -0.01fF
C54233 NOR2X1_LOC_216/Y INVX1_LOC_91/A 0.17fF
C54234 INVX1_LOC_28/A NAND2X1_LOC_843/a_36_24# 0.01fF
C54235 NAND2X1_LOC_656/A NAND2X1_LOC_63/Y 0.02fF
C54236 INVX1_LOC_50/A NOR2X1_LOC_215/A 0.01fF
C54237 INVX1_LOC_14/A NOR2X1_LOC_301/A 0.14fF
C54238 INVX1_LOC_177/A NOR2X1_LOC_862/B 0.02fF
C54239 NOR2X1_LOC_514/a_36_216# NOR2X1_LOC_649/B 0.01fF
C54240 INVX1_LOC_49/A NOR2X1_LOC_691/B 0.06fF
C54241 INVX1_LOC_24/Y NOR2X1_LOC_621/A 0.23fF
C54242 NOR2X1_LOC_433/A INVX1_LOC_49/Y 0.03fF
C54243 NOR2X1_LOC_103/Y INVX1_LOC_26/A 0.10fF
C54244 NAND2X1_LOC_303/Y INVX1_LOC_296/A 0.27fF
C54245 INVX1_LOC_21/A NOR2X1_LOC_392/Y 0.07fF
C54246 NOR2X1_LOC_735/Y NOR2X1_LOC_357/Y 0.03fF
C54247 NOR2X1_LOC_274/B INVX1_LOC_32/A 0.15fF
C54248 NAND2X1_LOC_577/A NAND2X1_LOC_618/Y 0.13fF
C54249 NOR2X1_LOC_309/Y NOR2X1_LOC_661/a_36_216# 0.01fF
C54250 NAND2X1_LOC_783/A NAND2X1_LOC_783/a_36_24# 0.00fF
C54251 NOR2X1_LOC_283/a_36_216# NOR2X1_LOC_89/A 0.00fF
C54252 NOR2X1_LOC_152/a_36_216# INVX1_LOC_42/A 0.00fF
C54253 NAND2X1_LOC_115/a_36_24# INVX1_LOC_133/A 0.01fF
C54254 NOR2X1_LOC_561/Y INVX1_LOC_157/Y -0.04fF
C54255 NAND2X1_LOC_852/Y NAND2X1_LOC_770/Y 0.80fF
C54256 NOR2X1_LOC_189/A INVX1_LOC_102/A 0.01fF
C54257 NOR2X1_LOC_121/A INVX1_LOC_46/Y 0.05fF
C54258 INVX1_LOC_83/A INVX1_LOC_193/A 0.02fF
C54259 INVX1_LOC_30/A NAND2X1_LOC_454/Y 0.05fF
C54260 NOR2X1_LOC_433/A NAND2X1_LOC_288/a_36_24# 0.01fF
C54261 INVX1_LOC_255/Y NOR2X1_LOC_861/a_36_216# 0.02fF
C54262 NOR2X1_LOC_169/B NAND2X1_LOC_72/B 0.04fF
C54263 NOR2X1_LOC_310/Y INVX1_LOC_19/A 0.01fF
C54264 NOR2X1_LOC_322/Y INVX1_LOC_46/A 0.15fF
C54265 NAND2X1_LOC_564/A NOR2X1_LOC_103/Y 0.01fF
C54266 NOR2X1_LOC_52/B INVX1_LOC_49/Y 2.44fF
C54267 INVX1_LOC_58/A NAND2X1_LOC_53/Y 0.14fF
C54268 INVX1_LOC_34/A NOR2X1_LOC_89/A 0.52fF
C54269 NOR2X1_LOC_679/B INVX1_LOC_42/A 0.01fF
C54270 INVX1_LOC_27/A INVX1_LOC_50/Y 0.03fF
C54271 NOR2X1_LOC_109/Y NAND2X1_LOC_780/Y 0.04fF
C54272 INVX1_LOC_45/A INVX1_LOC_26/A 0.10fF
C54273 INVX1_LOC_18/A NOR2X1_LOC_158/Y 0.10fF
C54274 INVX1_LOC_31/A NOR2X1_LOC_105/a_36_216# 0.00fF
C54275 INVX1_LOC_229/Y INVX1_LOC_241/Y 0.04fF
C54276 NOR2X1_LOC_142/Y NOR2X1_LOC_114/Y 0.04fF
C54277 NOR2X1_LOC_261/a_36_216# NOR2X1_LOC_471/Y 0.00fF
C54278 NOR2X1_LOC_577/Y INVX1_LOC_32/A 0.21fF
C54279 NOR2X1_LOC_20/Y INVX1_LOC_64/A 0.01fF
C54280 NOR2X1_LOC_75/Y NOR2X1_LOC_598/B 0.01fF
C54281 INVX1_LOC_17/A NOR2X1_LOC_489/B 0.01fF
C54282 INVX1_LOC_238/A NAND2X1_LOC_725/Y 0.06fF
C54283 NOR2X1_LOC_168/B NOR2X1_LOC_633/A 0.02fF
C54284 NOR2X1_LOC_717/B NOR2X1_LOC_155/A 0.01fF
C54285 INVX1_LOC_35/A NAND2X1_LOC_30/Y 0.05fF
C54286 NOR2X1_LOC_167/Y INVX1_LOC_37/A 0.03fF
C54287 INVX1_LOC_93/Y NAND2X1_LOC_642/Y 0.01fF
C54288 INVX1_LOC_303/Y INVX1_LOC_37/A 0.01fF
C54289 NOR2X1_LOC_78/A INVX1_LOC_59/Y 0.03fF
C54290 NOR2X1_LOC_487/a_36_216# NOR2X1_LOC_693/Y 0.01fF
C54291 INVX1_LOC_22/A NAND2X1_LOC_489/Y 0.00fF
C54292 NOR2X1_LOC_329/B INVX1_LOC_118/A 0.13fF
C54293 INVX1_LOC_232/Y NAND2X1_LOC_82/a_36_24# 0.01fF
C54294 NOR2X1_LOC_91/A NOR2X1_LOC_518/Y 0.03fF
C54295 NOR2X1_LOC_93/Y NOR2X1_LOC_92/Y 0.06fF
C54296 INVX1_LOC_33/A INVX1_LOC_4/A 0.03fF
C54297 NOR2X1_LOC_272/Y NOR2X1_LOC_468/Y 0.10fF
C54298 NOR2X1_LOC_454/Y NAND2X1_LOC_149/Y 0.19fF
C54299 INVX1_LOC_282/A INVX1_LOC_38/A 0.08fF
C54300 NOR2X1_LOC_78/A INVX1_LOC_176/A 0.01fF
C54301 INVX1_LOC_35/A NOR2X1_LOC_134/Y 0.03fF
C54302 NOR2X1_LOC_658/Y INVX1_LOC_23/A 0.07fF
C54303 INVX1_LOC_105/A INVX1_LOC_78/A 0.07fF
C54304 INVX1_LOC_45/A NOR2X1_LOC_255/Y 0.09fF
C54305 NOR2X1_LOC_828/A NOR2X1_LOC_155/A 0.00fF
C54306 INVX1_LOC_285/Y INVX1_LOC_281/A 0.17fF
C54307 INVX1_LOC_132/A INVX1_LOC_87/A 0.07fF
C54308 INVX1_LOC_71/A INVX1_LOC_26/A 0.01fF
C54309 NOR2X1_LOC_348/B INVX1_LOC_32/A 0.07fF
C54310 NOR2X1_LOC_554/B NOR2X1_LOC_105/Y 0.11fF
C54311 NOR2X1_LOC_679/B INVX1_LOC_78/A 0.09fF
C54312 NOR2X1_LOC_577/Y NAND2X1_LOC_175/Y 0.00fF
C54313 INVX1_LOC_21/A NAND2X1_LOC_357/A 0.03fF
C54314 NOR2X1_LOC_91/A NOR2X1_LOC_13/Y 0.07fF
C54315 NOR2X1_LOC_657/a_36_216# INVX1_LOC_103/A 0.00fF
C54316 INVX1_LOC_141/Y NOR2X1_LOC_109/Y 0.18fF
C54317 NOR2X1_LOC_631/B INVX1_LOC_76/A 0.25fF
C54318 NOR2X1_LOC_609/a_36_216# NOR2X1_LOC_383/B 0.00fF
C54319 INVX1_LOC_269/A INVX1_LOC_24/Y 0.23fF
C54320 NOR2X1_LOC_811/B NOR2X1_LOC_812/A 0.01fF
C54321 INVX1_LOC_125/Y NOR2X1_LOC_536/A 0.35fF
C54322 INVX1_LOC_225/A INVX1_LOC_87/A 0.14fF
C54323 INVX1_LOC_31/A NOR2X1_LOC_649/Y 0.18fF
C54324 INVX1_LOC_312/Y NOR2X1_LOC_109/Y 0.03fF
C54325 INVX1_LOC_25/A NAND2X1_LOC_79/Y 0.02fF
C54326 NOR2X1_LOC_151/Y NOR2X1_LOC_155/A 2.12fF
C54327 INVX1_LOC_16/A INVX1_LOC_290/Y 0.07fF
C54328 NOR2X1_LOC_13/Y INVX1_LOC_23/A 0.01fF
C54329 NOR2X1_LOC_272/Y NOR2X1_LOC_389/A 0.39fF
C54330 NAND2X1_LOC_363/B NOR2X1_LOC_68/A 0.24fF
C54331 INVX1_LOC_17/A INVX1_LOC_14/A 0.07fF
C54332 INVX1_LOC_251/Y INVX1_LOC_4/Y 0.00fF
C54333 INVX1_LOC_266/Y NAND2X1_LOC_470/B 0.02fF
C54334 NOR2X1_LOC_711/Y INVX1_LOC_117/A 0.02fF
C54335 VDD NOR2X1_LOC_603/Y 0.12fF
C54336 NOR2X1_LOC_269/Y NOR2X1_LOC_331/B 1.32fF
C54337 NOR2X1_LOC_598/B NAND2X1_LOC_162/B 0.03fF
C54338 INVX1_LOC_39/A NAND2X1_LOC_577/A 0.01fF
C54339 INVX1_LOC_37/A INVX1_LOC_76/A 0.39fF
C54340 NAND2X1_LOC_715/a_36_24# INVX1_LOC_109/A 0.00fF
C54341 INVX1_LOC_279/A INVX1_LOC_109/Y 0.01fF
C54342 INVX1_LOC_226/Y INVX1_LOC_3/Y 0.08fF
C54343 INVX1_LOC_278/A NOR2X1_LOC_238/Y 0.07fF
C54344 NAND2X1_LOC_338/B NAND2X1_LOC_471/Y 0.02fF
C54345 INVX1_LOC_40/A INVX1_LOC_4/A 0.77fF
C54346 NAND2X1_LOC_364/Y INVX1_LOC_23/A 0.03fF
C54347 INVX1_LOC_136/A INVX1_LOC_306/Y 0.03fF
C54348 INVX1_LOC_55/Y INVX1_LOC_186/Y 0.07fF
C54349 INVX1_LOC_5/A NOR2X1_LOC_791/B 0.01fF
C54350 INVX1_LOC_22/A INVX1_LOC_32/A 0.16fF
C54351 NAND2X1_LOC_213/A NOR2X1_LOC_389/A 0.14fF
C54352 INVX1_LOC_27/A NOR2X1_LOC_248/Y 0.01fF
C54353 INVX1_LOC_40/Y INVX1_LOC_252/A 0.00fF
C54354 NOR2X1_LOC_742/A NAND2X1_LOC_252/a_36_24# 0.00fF
C54355 NOR2X1_LOC_598/B NOR2X1_LOC_537/A 0.02fF
C54356 INVX1_LOC_179/Y NAND2X1_LOC_72/B 0.72fF
C54357 NAND2X1_LOC_35/Y NAND2X1_LOC_559/a_36_24# 0.01fF
C54358 NAND2X1_LOC_363/B NOR2X1_LOC_545/A 0.01fF
C54359 INVX1_LOC_51/A NOR2X1_LOC_419/Y 0.00fF
C54360 NAND2X1_LOC_655/A INVX1_LOC_54/A 0.07fF
C54361 NAND2X1_LOC_175/B INVX1_LOC_23/A 0.07fF
C54362 NAND2X1_LOC_555/Y INVX1_LOC_14/A 0.17fF
C54363 NOR2X1_LOC_71/Y NOR2X1_LOC_76/B 0.03fF
C54364 NOR2X1_LOC_91/A NOR2X1_LOC_504/Y 0.03fF
C54365 INVX1_LOC_35/A INVX1_LOC_49/A 0.22fF
C54366 NOR2X1_LOC_356/A NAND2X1_LOC_74/B 0.00fF
C54367 INVX1_LOC_89/A NOR2X1_LOC_240/B 0.05fF
C54368 INVX1_LOC_256/A INVX1_LOC_225/Y 0.12fF
C54369 INVX1_LOC_36/A NAND2X1_LOC_780/Y 0.07fF
C54370 INVX1_LOC_147/Y NOR2X1_LOC_351/Y 0.16fF
C54371 INVX1_LOC_21/A NOR2X1_LOC_744/a_36_216# 0.00fF
C54372 NAND2X1_LOC_468/B INVX1_LOC_54/A 0.04fF
C54373 NOR2X1_LOC_91/A INVX1_LOC_256/Y 0.07fF
C54374 INVX1_LOC_64/A INVX1_LOC_33/A 0.20fF
C54375 INVX1_LOC_91/A NOR2X1_LOC_197/B 0.10fF
C54376 INVX1_LOC_48/A NAND2X1_LOC_73/a_36_24# 0.00fF
C54377 INVX1_LOC_36/A NAND2X1_LOC_121/a_36_24# 0.00fF
C54378 INVX1_LOC_22/A NAND2X1_LOC_175/Y 0.08fF
C54379 NAND2X1_LOC_800/Y INVX1_LOC_231/A 0.00fF
C54380 INVX1_LOC_22/A NOR2X1_LOC_821/a_36_216# 0.03fF
C54381 INVX1_LOC_286/Y INVX1_LOC_221/Y 0.03fF
C54382 NAND2X1_LOC_342/Y INVX1_LOC_57/A 0.00fF
C54383 INVX1_LOC_28/A INVX1_LOC_290/Y 0.07fF
C54384 INVX1_LOC_295/A D_INPUT_5 0.06fF
C54385 NOR2X1_LOC_369/a_36_216# NAND2X1_LOC_793/B 0.01fF
C54386 NOR2X1_LOC_181/A NOR2X1_LOC_155/A 0.01fF
C54387 INVX1_LOC_114/A INVX1_LOC_117/A 0.03fF
C54388 NOR2X1_LOC_256/Y INVX1_LOC_284/A 0.04fF
C54389 NOR2X1_LOC_74/A NAND2X1_LOC_74/B 0.07fF
C54390 NAND2X1_LOC_213/A NOR2X1_LOC_596/A 0.12fF
C54391 INVX1_LOC_256/Y INVX1_LOC_23/A 0.09fF
C54392 INVX1_LOC_76/A NOR2X1_LOC_743/Y 0.05fF
C54393 D_GATE_366 NOR2X1_LOC_467/A 0.07fF
C54394 NAND2X1_LOC_149/Y INVX1_LOC_77/A 0.07fF
C54395 INVX1_LOC_5/A NOR2X1_LOC_124/B 0.20fF
C54396 NOR2X1_LOC_151/Y NOR2X1_LOC_833/B 0.02fF
C54397 INVX1_LOC_27/A NOR2X1_LOC_718/Y 0.01fF
C54398 NOR2X1_LOC_106/A NOR2X1_LOC_334/Y 0.00fF
C54399 INVX1_LOC_13/A NOR2X1_LOC_843/B 0.07fF
C54400 INVX1_LOC_35/A INVX1_LOC_2/A 0.08fF
C54401 NAND2X1_LOC_214/B NOR2X1_LOC_6/B 0.02fF
C54402 INVX1_LOC_45/A INVX1_LOC_141/A 0.01fF
C54403 NOR2X1_LOC_15/Y INVX1_LOC_314/Y 0.36fF
C54404 INPUT_0 NOR2X1_LOC_89/A 0.16fF
C54405 NOR2X1_LOC_9/Y NAND2X1_LOC_74/B 0.03fF
C54406 INVX1_LOC_58/A NOR2X1_LOC_500/Y 0.10fF
C54407 INVX1_LOC_64/A NOR2X1_LOC_521/a_36_216# 0.00fF
C54408 INVX1_LOC_58/A INVX1_LOC_226/Y 0.27fF
C54409 NOR2X1_LOC_278/A INVX1_LOC_306/Y 0.51fF
C54410 INVX1_LOC_5/A NOR2X1_LOC_802/A 0.03fF
C54411 NAND2X1_LOC_162/a_36_24# NOR2X1_LOC_467/A 0.00fF
C54412 INVX1_LOC_35/A NOR2X1_LOC_226/A 0.10fF
C54413 NOR2X1_LOC_88/Y NOR2X1_LOC_305/Y 0.07fF
C54414 INVX1_LOC_17/A NAND2X1_LOC_84/Y 1.42fF
C54415 INVX1_LOC_22/A NOR2X1_LOC_622/A 0.14fF
C54416 INVX1_LOC_95/Y INVX1_LOC_84/A 0.07fF
C54417 INVX1_LOC_36/A INVX1_LOC_141/Y 0.01fF
C54418 NOR2X1_LOC_389/A NAND2X1_LOC_364/A 0.01fF
C54419 INVX1_LOC_27/A NOR2X1_LOC_6/B 0.23fF
C54420 NAND2X1_LOC_656/Y INVX1_LOC_28/Y 0.03fF
C54421 NOR2X1_LOC_123/B INVX1_LOC_26/A 0.15fF
C54422 NOR2X1_LOC_392/B NOR2X1_LOC_440/B 0.07fF
C54423 INVX1_LOC_36/A INVX1_LOC_312/Y 0.07fF
C54424 INVX1_LOC_117/A INVX1_LOC_307/A 0.07fF
C54425 NOR2X1_LOC_294/Y INVX1_LOC_36/A 0.16fF
C54426 NAND2X1_LOC_656/Y INVX1_LOC_270/A 0.10fF
C54427 INVX1_LOC_41/A INVX1_LOC_269/A 0.10fF
C54428 NOR2X1_LOC_122/a_36_216# INVX1_LOC_92/A 0.00fF
C54429 INVX1_LOC_64/A NAND2X1_LOC_726/Y 0.02fF
C54430 NOR2X1_LOC_78/A NOR2X1_LOC_340/A 0.89fF
C54431 NAND2X1_LOC_218/B INPUT_3 0.10fF
C54432 NOR2X1_LOC_275/a_36_216# NOR2X1_LOC_759/Y 0.00fF
C54433 INVX1_LOC_58/A INVX1_LOC_10/A 0.30fF
C54434 INVX1_LOC_117/A NOR2X1_LOC_445/B 0.16fF
C54435 NAND2X1_LOC_577/A INVX1_LOC_61/A 0.02fF
C54436 NOR2X1_LOC_305/Y INVX1_LOC_84/A 0.07fF
C54437 NOR2X1_LOC_68/A INVX1_LOC_30/A 0.43fF
C54438 NOR2X1_LOC_598/B NOR2X1_LOC_470/A 0.10fF
C54439 INVX1_LOC_34/A INVX1_LOC_11/A 0.07fF
C54440 NOR2X1_LOC_598/B NOR2X1_LOC_424/Y 0.09fF
C54441 NAND2X1_LOC_763/B NOR2X1_LOC_68/A 0.03fF
C54442 NAND2X1_LOC_785/B INVX1_LOC_41/Y 0.05fF
C54443 NOR2X1_LOC_536/A NAND2X1_LOC_288/A 0.09fF
C54444 NOR2X1_LOC_357/Y INVX1_LOC_186/Y 0.02fF
C54445 NOR2X1_LOC_598/B NOR2X1_LOC_717/B 0.04fF
C54446 NOR2X1_LOC_637/B NOR2X1_LOC_590/A 0.32fF
C54447 NAND2X1_LOC_775/a_36_24# NAND2X1_LOC_579/A 0.07fF
C54448 INVX1_LOC_102/Y INVX1_LOC_26/A 0.26fF
C54449 INVX1_LOC_43/Y INVX1_LOC_33/A 0.04fF
C54450 NOR2X1_LOC_246/Y INVX1_LOC_57/A 0.01fF
C54451 NAND2X1_LOC_392/A INVX1_LOC_93/A 0.05fF
C54452 NOR2X1_LOC_48/B NAND2X1_LOC_655/A 0.08fF
C54453 INVX1_LOC_24/A NOR2X1_LOC_372/Y 0.04fF
C54454 NOR2X1_LOC_197/A NOR2X1_LOC_254/Y 0.01fF
C54455 INVX1_LOC_90/A INVX1_LOC_129/A 0.00fF
C54456 NOR2X1_LOC_332/B NAND2X1_LOC_291/B 0.03fF
C54457 INVX1_LOC_21/A INVX1_LOC_25/Y 0.01fF
C54458 INVX1_LOC_87/Y INVX1_LOC_57/A 0.01fF
C54459 NOR2X1_LOC_443/Y INVX1_LOC_148/A 0.00fF
C54460 INVX1_LOC_212/A INVX1_LOC_122/Y 0.02fF
C54461 NOR2X1_LOC_288/A INVX1_LOC_134/A 0.05fF
C54462 NAND2X1_LOC_45/Y NOR2X1_LOC_247/Y 0.09fF
C54463 INVX1_LOC_97/Y NOR2X1_LOC_717/B 0.00fF
C54464 NOR2X1_LOC_614/Y NOR2X1_LOC_790/A 0.00fF
C54465 NAND2X1_LOC_656/Y NOR2X1_LOC_109/Y 0.07fF
C54466 INVX1_LOC_21/A NOR2X1_LOC_302/B 0.11fF
C54467 NOR2X1_LOC_536/A NOR2X1_LOC_653/Y 0.04fF
C54468 INVX1_LOC_25/A NOR2X1_LOC_750/A 0.03fF
C54469 NOR2X1_LOC_598/B NOR2X1_LOC_828/A 0.12fF
C54470 INVX1_LOC_17/A INVX1_LOC_111/Y 0.15fF
C54471 INVX1_LOC_12/A NOR2X1_LOC_422/Y 0.00fF
C54472 NOR2X1_LOC_180/B INVX1_LOC_53/A 0.15fF
C54473 NOR2X1_LOC_314/Y INVX1_LOC_12/A 0.03fF
C54474 NOR2X1_LOC_160/B INVX1_LOC_104/A 2.87fF
C54475 INVX1_LOC_27/A INVX1_LOC_30/Y 0.02fF
C54476 INVX1_LOC_11/A NAND2X1_LOC_231/Y 0.03fF
C54477 INVX1_LOC_35/A INPUT_1 0.51fF
C54478 NOR2X1_LOC_400/A INVX1_LOC_89/A 0.02fF
C54479 NAND2X1_LOC_562/Y NAND2X1_LOC_577/A 0.15fF
C54480 INVX1_LOC_13/Y NOR2X1_LOC_373/Y 0.01fF
C54481 INVX1_LOC_1/A NAND2X1_LOC_831/a_36_24# 0.00fF
C54482 NOR2X1_LOC_846/Y INVX1_LOC_83/A 0.01fF
C54483 INVX1_LOC_49/A NOR2X1_LOC_325/Y 0.02fF
C54484 NOR2X1_LOC_536/A INVX1_LOC_19/A 4.29fF
C54485 NOR2X1_LOC_691/A NOR2X1_LOC_729/A 0.03fF
C54486 NOR2X1_LOC_319/B NOR2X1_LOC_777/B 0.03fF
C54487 NOR2X1_LOC_147/B INVX1_LOC_142/A 0.75fF
C54488 INVX1_LOC_36/A INVX1_LOC_88/Y 0.04fF
C54489 INVX1_LOC_224/Y NOR2X1_LOC_368/A 0.06fF
C54490 NOR2X1_LOC_211/Y NOR2X1_LOC_389/B 0.02fF
C54491 INVX1_LOC_12/A INVX1_LOC_117/A 0.10fF
C54492 INVX1_LOC_230/Y NOR2X1_LOC_537/Y 0.43fF
C54493 NOR2X1_LOC_382/Y NOR2X1_LOC_143/a_36_216# 0.00fF
C54494 INVX1_LOC_33/A INVX1_LOC_130/Y 0.39fF
C54495 INVX1_LOC_73/A INVX1_LOC_53/A 0.07fF
C54496 INVX1_LOC_136/A INVX1_LOC_294/Y 0.03fF
C54497 INVX1_LOC_36/A NAND2X1_LOC_847/a_36_24# 0.00fF
C54498 NAND2X1_LOC_67/Y NOR2X1_LOC_665/A 0.08fF
C54499 NOR2X1_LOC_598/B NOR2X1_LOC_151/Y 0.17fF
C54500 NOR2X1_LOC_388/Y NOR2X1_LOC_360/Y 0.10fF
C54501 NOR2X1_LOC_295/Y NAND2X1_LOC_364/A 0.02fF
C54502 INVX1_LOC_90/A NOR2X1_LOC_849/A 0.09fF
C54503 NAND2X1_LOC_642/Y INVX1_LOC_87/A 0.03fF
C54504 INVX1_LOC_105/A NOR2X1_LOC_152/Y 0.07fF
C54505 NOR2X1_LOC_337/A INVX1_LOC_23/A 0.01fF
C54506 INVX1_LOC_233/A NOR2X1_LOC_322/Y 0.10fF
C54507 INVX1_LOC_45/A INVX1_LOC_149/A 0.01fF
C54508 INPUT_0 NAND2X1_LOC_804/A 0.01fF
C54509 NAND2X1_LOC_276/Y INVX1_LOC_24/A 0.03fF
C54510 INVX1_LOC_105/A NAND2X1_LOC_193/a_36_24# 0.02fF
C54511 NAND2X1_LOC_742/a_36_24# NOR2X1_LOC_576/B 0.04fF
C54512 NOR2X1_LOC_457/A NOR2X1_LOC_570/Y 0.03fF
C54513 INVX1_LOC_149/A NOR2X1_LOC_568/A 0.00fF
C54514 NOR2X1_LOC_208/Y NOR2X1_LOC_219/B 0.00fF
C54515 NOR2X1_LOC_569/A INVX1_LOC_53/A 0.03fF
C54516 NOR2X1_LOC_155/A NOR2X1_LOC_666/a_36_216# 0.00fF
C54517 INVX1_LOC_5/A NOR2X1_LOC_197/Y 0.04fF
C54518 NOR2X1_LOC_172/Y NAND2X1_LOC_593/Y 0.10fF
C54519 INVX1_LOC_269/A NOR2X1_LOC_299/Y 0.03fF
C54520 INVX1_LOC_90/A NOR2X1_LOC_440/B 0.01fF
C54521 INVX1_LOC_27/A NOR2X1_LOC_156/A 0.21fF
C54522 NOR2X1_LOC_71/Y NOR2X1_LOC_271/B 0.03fF
C54523 NAND2X1_LOC_57/a_36_24# NAND2X1_LOC_360/B 0.01fF
C54524 NOR2X1_LOC_208/Y INVX1_LOC_88/Y 0.07fF
C54525 NAND2X1_LOC_93/B INVX1_LOC_19/A 0.03fF
C54526 INVX1_LOC_1/A NOR2X1_LOC_333/A 0.01fF
C54527 NOR2X1_LOC_836/B NOR2X1_LOC_836/A 0.09fF
C54528 NOR2X1_LOC_68/A NAND2X1_LOC_722/A 0.16fF
C54529 INVX1_LOC_34/A NOR2X1_LOC_433/A 0.03fF
C54530 INVX1_LOC_35/A NOR2X1_LOC_706/Y 0.02fF
C54531 NOR2X1_LOC_781/Y INVX1_LOC_266/Y 0.01fF
C54532 INVX1_LOC_17/A NOR2X1_LOC_137/A 0.03fF
C54533 INVX1_LOC_1/A D_GATE_366 0.04fF
C54534 NAND2X1_LOC_425/Y INVX1_LOC_19/A 0.01fF
C54535 NOR2X1_LOC_592/A NOR2X1_LOC_130/A 0.01fF
C54536 INVX1_LOC_34/A NOR2X1_LOC_593/Y 0.02fF
C54537 INVX1_LOC_313/Y NOR2X1_LOC_359/a_36_216# 0.00fF
C54538 NOR2X1_LOC_78/B NOR2X1_LOC_457/B 0.07fF
C54539 INVX1_LOC_21/A INVX1_LOC_75/A 16.31fF
C54540 NOR2X1_LOC_662/A INVX1_LOC_285/A 0.01fF
C54541 D_GATE_662 INVX1_LOC_175/A 0.00fF
C54542 INVX1_LOC_24/A NOR2X1_LOC_352/Y 0.05fF
C54543 NOR2X1_LOC_653/Y NOR2X1_LOC_661/A 0.15fF
C54544 INVX1_LOC_208/A INVX1_LOC_177/Y 0.63fF
C54545 NOR2X1_LOC_772/B INVX1_LOC_286/A 0.10fF
C54546 NAND2X1_LOC_341/A INVX1_LOC_72/A 0.12fF
C54547 INVX1_LOC_24/A NAND2X1_LOC_374/Y 0.23fF
C54548 NOR2X1_LOC_720/B NOR2X1_LOC_520/B 0.18fF
C54549 NOR2X1_LOC_381/Y NOR2X1_LOC_19/B 0.09fF
C54550 INVX1_LOC_19/A NOR2X1_LOC_649/B -0.04fF
C54551 INVX1_LOC_174/A INVX1_LOC_89/A 0.32fF
C54552 INVX1_LOC_233/Y NOR2X1_LOC_45/B 0.16fF
C54553 NOR2X1_LOC_647/Y INVX1_LOC_13/A 0.12fF
C54554 INVX1_LOC_13/Y INVX1_LOC_286/A 0.07fF
C54555 NAND2X1_LOC_231/Y NOR2X1_LOC_433/A 0.48fF
C54556 INVX1_LOC_34/A NOR2X1_LOC_52/B 0.13fF
C54557 NOR2X1_LOC_782/a_36_216# INVX1_LOC_191/Y 0.00fF
C54558 INVX1_LOC_45/A INVX1_LOC_164/A 1.82fF
C54559 NOR2X1_LOC_447/A INVX1_LOC_37/A 0.07fF
C54560 INVX1_LOC_201/Y NAND2X1_LOC_127/a_36_24# 0.00fF
C54561 INVX1_LOC_36/A NAND2X1_LOC_656/Y 0.08fF
C54562 INVX1_LOC_278/A INVX1_LOC_95/Y 0.07fF
C54563 INVX1_LOC_64/A NOR2X1_LOC_486/Y 0.02fF
C54564 INVX1_LOC_286/Y INVX1_LOC_183/Y 0.03fF
C54565 NOR2X1_LOC_392/Y NOR2X1_LOC_670/Y 0.00fF
C54566 INVX1_LOC_90/A NOR2X1_LOC_514/A 0.03fF
C54567 NOR2X1_LOC_536/A INVX1_LOC_26/Y 0.01fF
C54568 INVX1_LOC_2/A NOR2X1_LOC_365/a_36_216# 0.00fF
C54569 NAND2X1_LOC_198/B NOR2X1_LOC_561/Y 0.03fF
C54570 INVX1_LOC_24/A NOR2X1_LOC_553/B 0.02fF
C54571 NOR2X1_LOC_598/B NOR2X1_LOC_567/a_36_216# 0.01fF
C54572 INVX1_LOC_77/A INVX1_LOC_16/A 0.14fF
C54573 NOR2X1_LOC_458/Y NOR2X1_LOC_458/B 0.03fF
C54574 INVX1_LOC_232/Y NOR2X1_LOC_84/A 0.01fF
C54575 INVX1_LOC_9/Y NOR2X1_LOC_577/Y 0.01fF
C54576 INVX1_LOC_224/A INPUT_0 0.03fF
C54577 NAND2X1_LOC_456/Y NAND2X1_LOC_254/Y 0.14fF
C54578 NAND2X1_LOC_214/B NOR2X1_LOC_124/A 0.01fF
C54579 NOR2X1_LOC_103/Y NOR2X1_LOC_368/A 0.14fF
C54580 NAND2X1_LOC_231/Y NOR2X1_LOC_52/B 0.01fF
C54581 INVX1_LOC_11/A INPUT_0 11.70fF
C54582 INVX1_LOC_135/A NOR2X1_LOC_360/Y 0.01fF
C54583 INVX1_LOC_36/A NAND2X1_LOC_638/Y 0.17fF
C54584 NOR2X1_LOC_334/Y NOR2X1_LOC_830/a_36_216# 0.01fF
C54585 NAND2X1_LOC_734/B NOR2X1_LOC_667/A 0.02fF
C54586 NAND2X1_LOC_381/Y INPUT_0 0.10fF
C54587 NAND2X1_LOC_557/Y NOR2X1_LOC_536/A 0.10fF
C54588 NOR2X1_LOC_304/Y INVX1_LOC_20/A 0.02fF
C54589 INVX1_LOC_136/A NOR2X1_LOC_356/A 0.03fF
C54590 INVX1_LOC_17/A INVX1_LOC_48/A 0.02fF
C54591 NOR2X1_LOC_222/a_36_216# INVX1_LOC_63/Y 0.01fF
C54592 INVX1_LOC_208/A INVX1_LOC_104/A 0.10fF
C54593 INVX1_LOC_55/Y INVX1_LOC_18/A 0.08fF
C54594 INVX1_LOC_166/A NAND2X1_LOC_659/a_36_24# 0.00fF
C54595 INVX1_LOC_5/A INVX1_LOC_2/Y 1.57fF
C54596 NOR2X1_LOC_470/B INVX1_LOC_91/A 0.01fF
C54597 NOR2X1_LOC_458/B INVX1_LOC_177/A 0.04fF
C54598 NAND2X1_LOC_741/B NOR2X1_LOC_385/Y 0.00fF
C54599 NOR2X1_LOC_99/Y INVX1_LOC_16/Y 0.27fF
C54600 NOR2X1_LOC_272/Y NAND2X1_LOC_469/B 0.01fF
C54601 NOR2X1_LOC_516/B INVX1_LOC_104/A 0.07fF
C54602 INVX1_LOC_225/Y INVX1_LOC_69/Y 0.10fF
C54603 NOR2X1_LOC_67/Y NAND2X1_LOC_207/B 0.07fF
C54604 D_INPUT_7 INVX1_LOC_140/A 0.19fF
C54605 INVX1_LOC_227/A INVX1_LOC_155/A 0.03fF
C54606 INVX1_LOC_90/A INVX1_LOC_41/Y 0.06fF
C54607 INVX1_LOC_177/A NOR2X1_LOC_388/a_36_216# 0.00fF
C54608 INVX1_LOC_103/A NOR2X1_LOC_78/A 0.00fF
C54609 NOR2X1_LOC_209/Y NOR2X1_LOC_731/Y 0.02fF
C54610 INVX1_LOC_147/A INVX1_LOC_30/A 0.26fF
C54611 NAND2X1_LOC_740/B INVX1_LOC_72/A 0.04fF
C54612 INVX1_LOC_32/A INVX1_LOC_186/Y 0.07fF
C54613 INVX1_LOC_124/A INVX1_LOC_16/A 0.09fF
C54614 NOR2X1_LOC_2/Y INVX1_LOC_30/A 0.19fF
C54615 INVX1_LOC_45/A NOR2X1_LOC_368/A 0.03fF
C54616 INVX1_LOC_21/A NAND2X1_LOC_453/A 0.07fF
C54617 NOR2X1_LOC_859/A NAND2X1_LOC_348/A 0.02fF
C54618 NAND2X1_LOC_372/a_36_24# NOR2X1_LOC_78/B 0.00fF
C54619 INVX1_LOC_5/A NAND2X1_LOC_230/a_36_24# 0.00fF
C54620 INVX1_LOC_90/A NAND2X1_LOC_593/Y 0.07fF
C54621 NAND2X1_LOC_391/Y VDD 0.18fF
C54622 INVX1_LOC_84/A INVX1_LOC_271/Y 0.07fF
C54623 INVX1_LOC_89/A INVX1_LOC_153/A 0.01fF
C54624 NOR2X1_LOC_99/Y NAND2X1_LOC_205/A 0.19fF
C54625 INVX1_LOC_50/A NAND2X1_LOC_802/Y 0.02fF
C54626 INVX1_LOC_136/A NOR2X1_LOC_74/A 0.30fF
C54627 INVX1_LOC_234/A NOR2X1_LOC_6/B 0.00fF
C54628 NOR2X1_LOC_667/A INVX1_LOC_25/Y 0.15fF
C54629 NOR2X1_LOC_669/Y INVX1_LOC_20/A 0.53fF
C54630 NOR2X1_LOC_82/A NAND2X1_LOC_642/Y 0.22fF
C54631 NOR2X1_LOC_292/Y INVX1_LOC_72/A 0.01fF
C54632 NOR2X1_LOC_658/Y INVX1_LOC_6/A 0.17fF
C54633 INVX1_LOC_13/A INVX1_LOC_34/Y 0.09fF
C54634 INVX1_LOC_292/A NOR2X1_LOC_78/A 0.07fF
C54635 INVX1_LOC_12/A INVX1_LOC_3/Y 0.07fF
C54636 INVX1_LOC_35/A INVX1_LOC_118/A 0.17fF
C54637 NOR2X1_LOC_778/A NAND2X1_LOC_496/a_36_24# 0.00fF
C54638 INVX1_LOC_178/A NAND2X1_LOC_687/A 0.05fF
C54639 INVX1_LOC_28/A INVX1_LOC_77/A 0.08fF
C54640 INVX1_LOC_58/A INVX1_LOC_307/A 0.10fF
C54641 NOR2X1_LOC_91/A NOR2X1_LOC_697/Y 0.00fF
C54642 INVX1_LOC_235/Y INVX1_LOC_194/Y 0.03fF
C54643 INPUT_6 NOR2X1_LOC_51/A 0.31fF
C54644 NOR2X1_LOC_79/A NOR2X1_LOC_717/A 0.01fF
C54645 INVX1_LOC_136/A NOR2X1_LOC_9/Y 0.11fF
C54646 NAND2X1_LOC_470/B INVX1_LOC_19/A 0.94fF
C54647 NOR2X1_LOC_413/Y NAND2X1_LOC_624/A 0.02fF
C54648 INVX1_LOC_286/Y INVX1_LOC_91/A 0.07fF
C54649 NAND2X1_LOC_35/Y NOR2X1_LOC_629/Y 0.11fF
C54650 INVX1_LOC_30/Y NAND2X1_LOC_200/B 0.08fF
C54651 NOR2X1_LOC_270/Y INVX1_LOC_285/Y 0.10fF
C54652 NOR2X1_LOC_389/A NOR2X1_LOC_405/A 0.30fF
C54653 NOR2X1_LOC_441/Y NOR2X1_LOC_139/Y 0.05fF
C54654 NOR2X1_LOC_390/a_36_216# INVX1_LOC_313/Y 0.00fF
C54655 NAND2X1_LOC_350/A NAND2X1_LOC_468/B 0.19fF
C54656 NOR2X1_LOC_736/Y INVX1_LOC_63/Y 0.02fF
C54657 NOR2X1_LOC_703/B NOR2X1_LOC_337/Y 0.02fF
C54658 INVX1_LOC_57/A INVX1_LOC_285/A 0.95fF
C54659 INVX1_LOC_23/A NOR2X1_LOC_697/Y 0.05fF
C54660 INVX1_LOC_57/A INVX1_LOC_265/Y 0.02fF
C54661 INVX1_LOC_89/A INVX1_LOC_259/A 0.04fF
C54662 NOR2X1_LOC_207/A NOR2X1_LOC_214/B 0.01fF
C54663 INVX1_LOC_57/A NOR2X1_LOC_814/A 0.40fF
C54664 INVX1_LOC_290/A NAND2X1_LOC_662/Y 0.07fF
C54665 NOR2X1_LOC_433/A INPUT_0 0.07fF
C54666 NOR2X1_LOC_441/Y NAND2X1_LOC_468/B 0.41fF
C54667 NOR2X1_LOC_13/Y INVX1_LOC_6/A 0.01fF
C54668 INVX1_LOC_221/Y VDD 0.26fF
C54669 NAND2X1_LOC_733/B NOR2X1_LOC_380/A 0.11fF
C54670 NOR2X1_LOC_561/Y INVX1_LOC_53/Y 0.02fF
C54671 NOR2X1_LOC_6/B NOR2X1_LOC_19/B 0.20fF
C54672 INVX1_LOC_295/A NAND2X1_LOC_451/Y 0.04fF
C54673 INVX1_LOC_217/A NAND2X1_LOC_623/B 0.01fF
C54674 INVX1_LOC_159/A INVX1_LOC_91/A 0.07fF
C54675 NOR2X1_LOC_205/Y INVX1_LOC_281/A 0.00fF
C54676 NOR2X1_LOC_790/B INVX1_LOC_220/A 0.03fF
C54677 NOR2X1_LOC_208/Y INVX1_LOC_78/Y 0.31fF
C54678 NOR2X1_LOC_711/a_36_216# INVX1_LOC_85/Y 0.00fF
C54679 INVX1_LOC_262/Y INVX1_LOC_296/A 0.04fF
C54680 NAND2X1_LOC_190/a_36_24# INVX1_LOC_307/A 0.01fF
C54681 NOR2X1_LOC_78/B NOR2X1_LOC_180/B 0.05fF
C54682 INVX1_LOC_134/A NOR2X1_LOC_863/A 0.02fF
C54683 INVX1_LOC_303/A INVX1_LOC_286/A 0.03fF
C54684 NOR2X1_LOC_191/B INVX1_LOC_91/A 0.10fF
C54685 NAND2X1_LOC_577/A D_INPUT_3 0.09fF
C54686 NOR2X1_LOC_781/A INVX1_LOC_83/A 0.10fF
C54687 INVX1_LOC_271/Y INVX1_LOC_15/A 0.11fF
C54688 NOR2X1_LOC_566/a_36_216# NOR2X1_LOC_360/Y 0.01fF
C54689 NOR2X1_LOC_82/A NOR2X1_LOC_271/Y 0.04fF
C54690 NAND2X1_LOC_577/A NAND2X1_LOC_618/a_36_24# 0.01fF
C54691 NOR2X1_LOC_52/B INPUT_0 13.27fF
C54692 INVX1_LOC_30/A NOR2X1_LOC_364/a_36_216# 0.00fF
C54693 NOR2X1_LOC_121/A INPUT_1 0.03fF
C54694 INVX1_LOC_89/A NAND2X1_LOC_666/a_36_24# 0.00fF
C54695 INVX1_LOC_88/A INVX1_LOC_54/A 2.23fF
C54696 NOR2X1_LOC_790/A NOR2X1_LOC_862/B 0.04fF
C54697 NOR2X1_LOC_29/a_36_216# INVX1_LOC_3/Y 0.01fF
C54698 NOR2X1_LOC_589/A INVX1_LOC_89/A 0.11fF
C54699 NOR2X1_LOC_544/A INVX1_LOC_182/A 0.01fF
C54700 INVX1_LOC_58/A INVX1_LOC_12/A 0.62fF
C54701 NOR2X1_LOC_565/a_36_216# INVX1_LOC_177/A 0.00fF
C54702 NOR2X1_LOC_816/A NAND2X1_LOC_846/a_36_24# 0.00fF
C54703 INVX1_LOC_164/A NOR2X1_LOC_123/B 0.04fF
C54704 INVX1_LOC_89/A NAND2X1_LOC_377/Y 0.01fF
C54705 INVX1_LOC_177/Y NAND2X1_LOC_211/Y 0.01fF
C54706 INVX1_LOC_67/A NOR2X1_LOC_78/A 0.03fF
C54707 NOR2X1_LOC_703/B VDD 0.02fF
C54708 NAND2X1_LOC_198/B INVX1_LOC_76/A 0.30fF
C54709 INVX1_LOC_58/Y INVX1_LOC_29/A 0.06fF
C54710 INVX1_LOC_35/A NAND2X1_LOC_63/Y 0.09fF
C54711 NOR2X1_LOC_457/B INVX1_LOC_46/A 0.07fF
C54712 INVX1_LOC_90/A NAND2X1_LOC_692/a_36_24# 0.00fF
C54713 NOR2X1_LOC_526/Y INVX1_LOC_91/Y 0.01fF
C54714 INVX1_LOC_286/A INVX1_LOC_168/A 0.02fF
C54715 INVX1_LOC_312/A NOR2X1_LOC_536/A 0.01fF
C54716 NAND2X1_LOC_474/Y NAND2X1_LOC_475/Y 0.01fF
C54717 INVX1_LOC_1/A INVX1_LOC_123/Y 0.03fF
C54718 NOR2X1_LOC_723/Y INVX1_LOC_281/A 0.08fF
C54719 NOR2X1_LOC_91/Y NAND2X1_LOC_721/A 0.02fF
C54720 NAND2X1_LOC_656/A D_INPUT_3 1.24fF
C54721 INVX1_LOC_77/A NOR2X1_LOC_35/Y 0.03fF
C54722 INVX1_LOC_75/A NAND2X1_LOC_6/a_36_24# 0.00fF
C54723 NAND2X1_LOC_656/A INVX1_LOC_14/Y 0.19fF
C54724 INVX1_LOC_89/A INVX1_LOC_171/A 0.03fF
C54725 NOR2X1_LOC_295/Y NOR2X1_LOC_405/A 0.02fF
C54726 NOR2X1_LOC_639/B NOR2X1_LOC_584/Y 0.11fF
C54727 NOR2X1_LOC_78/B NOR2X1_LOC_704/Y 0.02fF
C54728 INVX1_LOC_59/A INVX1_LOC_84/A 0.02fF
C54729 INVX1_LOC_256/Y INVX1_LOC_6/A 0.07fF
C54730 NOR2X1_LOC_178/Y NOR2X1_LOC_178/a_36_216# 0.00fF
C54731 INVX1_LOC_34/A INVX1_LOC_199/A 0.06fF
C54732 INVX1_LOC_18/A INVX1_LOC_66/Y 0.01fF
C54733 INVX1_LOC_83/A NOR2X1_LOC_738/A 0.05fF
C54734 INVX1_LOC_164/A INVX1_LOC_102/Y 0.05fF
C54735 INVX1_LOC_34/A INVX1_LOC_74/A 0.02fF
C54736 NAND2X1_LOC_832/Y INVX1_LOC_16/A 0.17fF
C54737 D_INPUT_4 INPUT_5 1.36fF
C54738 NOR2X1_LOC_52/B NAND2X1_LOC_649/B 0.01fF
C54739 INVX1_LOC_213/Y NOR2X1_LOC_833/Y 0.02fF
C54740 NAND2X1_LOC_837/Y NOR2X1_LOC_492/Y 0.04fF
C54741 NOR2X1_LOC_360/Y INVX1_LOC_280/A 0.04fF
C54742 INVX1_LOC_311/A NOR2X1_LOC_302/B 0.02fF
C54743 INVX1_LOC_135/A NOR2X1_LOC_567/B 0.07fF
C54744 NAND2X1_LOC_286/B NOR2X1_LOC_278/Y 0.29fF
C54745 NOR2X1_LOC_644/B NOR2X1_LOC_155/A 0.01fF
C54746 INVX1_LOC_254/A NAND2X1_LOC_96/A 0.01fF
C54747 NOR2X1_LOC_366/B NOR2X1_LOC_269/Y 0.01fF
C54748 INVX1_LOC_41/Y INVX1_LOC_38/A 0.04fF
C54749 NOR2X1_LOC_617/Y NAND2X1_LOC_849/B 0.05fF
C54750 NOR2X1_LOC_561/Y NOR2X1_LOC_113/B 0.01fF
C54751 NOR2X1_LOC_773/Y NOR2X1_LOC_192/A 0.02fF
C54752 INVX1_LOC_104/A NAND2X1_LOC_211/Y 0.01fF
C54753 INVX1_LOC_41/A INVX1_LOC_12/Y 0.01fF
C54754 NOR2X1_LOC_220/A NOR2X1_LOC_405/A 0.02fF
C54755 NOR2X1_LOC_647/A NOR2X1_LOC_646/B 0.03fF
C54756 NAND2X1_LOC_593/Y INVX1_LOC_38/A 0.07fF
C54757 INVX1_LOC_31/A NOR2X1_LOC_697/Y 0.06fF
C54758 NAND2X1_LOC_578/B NAND2X1_LOC_659/B 0.23fF
C54759 NOR2X1_LOC_717/a_36_216# INVX1_LOC_10/Y 0.00fF
C54760 NAND2X1_LOC_114/B INVX1_LOC_63/A 0.07fF
C54761 NOR2X1_LOC_222/Y NAND2X1_LOC_212/Y 0.01fF
C54762 NAND2X1_LOC_860/A NOR2X1_LOC_278/Y 0.03fF
C54763 INVX1_LOC_256/A INVX1_LOC_19/A 0.07fF
C54764 NOR2X1_LOC_401/B INVX1_LOC_20/A 0.24fF
C54765 INVX1_LOC_304/A INVX1_LOC_25/Y 0.15fF
C54766 NOR2X1_LOC_543/A NOR2X1_LOC_318/B 0.02fF
C54767 NAND2X1_LOC_181/Y NOR2X1_LOC_9/a_36_216# 0.00fF
C54768 NAND2X1_LOC_578/B VDD 0.02fF
C54769 NOR2X1_LOC_500/A NOR2X1_LOC_809/B 0.03fF
C54770 INVX1_LOC_59/A INVX1_LOC_15/A 0.03fF
C54771 INVX1_LOC_166/A NOR2X1_LOC_476/B 0.17fF
C54772 NOR2X1_LOC_219/Y INVX1_LOC_76/A 0.01fF
C54773 INPUT_5 INPUT_4 0.28fF
C54774 INVX1_LOC_312/Y INVX1_LOC_63/A 0.08fF
C54775 NOR2X1_LOC_294/Y INVX1_LOC_63/A 0.40fF
C54776 NAND2X1_LOC_187/a_36_24# NOR2X1_LOC_216/B 0.00fF
C54777 NAND2X1_LOC_347/B INVX1_LOC_47/Y 0.01fF
C54778 INVX1_LOC_53/Y INVX1_LOC_76/A 1.05fF
C54779 INVX1_LOC_30/A NAND2X1_LOC_768/Y 0.05fF
C54780 INVX1_LOC_34/A NOR2X1_LOC_675/a_36_216# 0.01fF
C54781 NAND2X1_LOC_51/B INVX1_LOC_75/A 0.12fF
C54782 INVX1_LOC_57/A NOR2X1_LOC_292/a_36_216# 0.00fF
C54783 INVX1_LOC_120/A NOR2X1_LOC_78/A 0.03fF
C54784 NAND2X1_LOC_130/a_36_24# NOR2X1_LOC_657/B 0.00fF
C54785 INVX1_LOC_306/A NAND2X1_LOC_642/Y 0.01fF
C54786 NOR2X1_LOC_679/B NAND2X1_LOC_802/Y 0.02fF
C54787 INVX1_LOC_18/A NAND2X1_LOC_489/Y 0.06fF
C54788 NOR2X1_LOC_665/A INVX1_LOC_76/A 0.03fF
C54789 NOR2X1_LOC_389/A INVX1_LOC_109/Y 0.10fF
C54790 INVX1_LOC_64/A NOR2X1_LOC_748/A 0.10fF
C54791 INVX1_LOC_311/A INVX1_LOC_75/A 0.03fF
C54792 NAND2X1_LOC_622/B NOR2X1_LOC_19/Y 0.01fF
C54793 NAND2X1_LOC_712/A VDD -0.00fF
C54794 VDD INVX1_LOC_137/Y 0.21fF
C54795 D_INPUT_6 NOR2X1_LOC_25/Y 0.45fF
C54796 NOR2X1_LOC_843/A NOR2X1_LOC_862/B 0.05fF
C54797 INVX1_LOC_225/Y NOR2X1_LOC_170/A 0.04fF
C54798 NOR2X1_LOC_507/A INVX1_LOC_122/A 0.20fF
C54799 NOR2X1_LOC_76/A NOR2X1_LOC_368/Y 0.03fF
C54800 INVX1_LOC_239/A INVX1_LOC_175/A 0.07fF
C54801 NOR2X1_LOC_92/Y NOR2X1_LOC_89/Y -0.03fF
C54802 NOR2X1_LOC_798/A NOR2X1_LOC_699/a_36_216# 0.00fF
C54803 NOR2X1_LOC_208/A INVX1_LOC_78/Y 0.01fF
C54804 NOR2X1_LOC_332/A INVX1_LOC_2/Y 0.03fF
C54805 INVX1_LOC_172/A NAND2X1_LOC_489/Y 0.03fF
C54806 NOR2X1_LOC_103/Y NAND2X1_LOC_471/Y 0.13fF
C54807 INVX1_LOC_89/A INVX1_LOC_20/A 0.07fF
C54808 GATE_811 NAND2X1_LOC_770/Y 0.07fF
C54809 NAND2X1_LOC_811/Y INVX1_LOC_297/A 0.07fF
C54810 NOR2X1_LOC_609/A INVX1_LOC_29/A 0.06fF
C54811 NOR2X1_LOC_19/B NOR2X1_LOC_124/A 0.00fF
C54812 NOR2X1_LOC_142/Y NOR2X1_LOC_66/Y 0.20fF
C54813 NAND2X1_LOC_181/a_36_24# NOR2X1_LOC_271/Y 0.00fF
C54814 INVX1_LOC_16/A INVX1_LOC_9/A 0.08fF
C54815 NOR2X1_LOC_76/A INVX1_LOC_46/A 0.46fF
C54816 NOR2X1_LOC_791/B INVX1_LOC_42/A 0.59fF
C54817 INVX1_LOC_183/Y VDD 0.21fF
C54818 NAND2X1_LOC_358/a_36_24# NAND2X1_LOC_96/A 0.00fF
C54819 NOR2X1_LOC_144/Y INVX1_LOC_84/A 0.06fF
C54820 INVX1_LOC_64/A NOR2X1_LOC_304/Y 0.02fF
C54821 INVX1_LOC_14/A INVX1_LOC_181/A 0.03fF
C54822 NOR2X1_LOC_419/Y INVX1_LOC_29/A 0.01fF
C54823 NAND2X1_LOC_387/B D_INPUT_5 0.01fF
C54824 INVX1_LOC_60/Y INVX1_LOC_27/Y 0.11fF
C54825 INVX1_LOC_35/A INVX1_LOC_39/A 0.03fF
C54826 NOR2X1_LOC_447/Y NOR2X1_LOC_584/Y 0.00fF
C54827 INVX1_LOC_256/A INVX1_LOC_26/Y 0.04fF
C54828 NOR2X1_LOC_716/B INVX1_LOC_29/A 0.07fF
C54829 INVX1_LOC_18/A INVX1_LOC_32/A 0.18fF
C54830 INVX1_LOC_215/Y NOR2X1_LOC_686/A 0.04fF
C54831 NOR2X1_LOC_6/B NOR2X1_LOC_126/a_36_216# 0.00fF
C54832 INVX1_LOC_17/A NOR2X1_LOC_383/B 0.03fF
C54833 INVX1_LOC_306/A NOR2X1_LOC_271/Y 0.26fF
C54834 NOR2X1_LOC_155/a_36_216# INVX1_LOC_117/A 0.01fF
C54835 NOR2X1_LOC_337/Y INVX1_LOC_91/A 0.02fF
C54836 INPUT_0 INVX1_LOC_74/A 0.02fF
C54837 INVX1_LOC_73/A INVX1_LOC_46/A 0.03fF
C54838 NOR2X1_LOC_168/B INVX1_LOC_63/A 0.03fF
C54839 NOR2X1_LOC_709/A NAND2X1_LOC_773/B 0.17fF
C54840 INVX1_LOC_58/A INVX1_LOC_200/A 0.07fF
C54841 NOR2X1_LOC_471/Y NOR2X1_LOC_383/B 0.07fF
C54842 INVX1_LOC_79/A VDD 0.00fF
C54843 NAND2X1_LOC_384/a_36_24# NOR2X1_LOC_99/Y 0.01fF
C54844 NAND2X1_LOC_811/Y NOR2X1_LOC_89/A 0.02fF
C54845 NOR2X1_LOC_553/B NOR2X1_LOC_197/B 0.03fF
C54846 INVX1_LOC_34/A NAND2X1_LOC_254/Y 0.07fF
C54847 NOR2X1_LOC_78/A NOR2X1_LOC_141/a_36_216# 0.00fF
C54848 INVX1_LOC_25/A INPUT_2 0.14fF
C54849 NAND2X1_LOC_778/Y NOR2X1_LOC_824/A 0.07fF
C54850 INVX1_LOC_233/Y INVX1_LOC_258/A 0.04fF
C54851 INVX1_LOC_18/A NAND2X1_LOC_175/Y 0.07fF
C54852 NAND2X1_LOC_35/Y INVX1_LOC_269/A 0.01fF
C54853 NOR2X1_LOC_590/A INVX1_LOC_57/A 0.72fF
C54854 NOR2X1_LOC_637/Y NOR2X1_LOC_329/Y 0.04fF
C54855 INVX1_LOC_291/Y NAND2X1_LOC_655/A 0.04fF
C54856 NOR2X1_LOC_124/B INVX1_LOC_42/A 0.01fF
C54857 NOR2X1_LOC_56/Y INVX1_LOC_91/A 0.07fF
C54858 INVX1_LOC_28/A INVX1_LOC_9/A 0.07fF
C54859 VDD NOR2X1_LOC_728/B -0.00fF
C54860 INVX1_LOC_143/A INVX1_LOC_125/A 0.74fF
C54861 INVX1_LOC_90/A INVX1_LOC_185/A 0.03fF
C54862 INVX1_LOC_255/Y NOR2X1_LOC_673/A 0.07fF
C54863 NOR2X1_LOC_254/a_36_216# INVX1_LOC_23/A 0.02fF
C54864 D_INPUT_1 INVX1_LOC_188/A 0.01fF
C54865 INVX1_LOC_22/Y INVX1_LOC_57/A 0.05fF
C54866 INVX1_LOC_266/Y NOR2X1_LOC_89/A 0.07fF
C54867 VDD INVX1_LOC_309/A 0.00fF
C54868 INVX1_LOC_11/A NAND2X1_LOC_25/a_36_24# 0.00fF
C54869 NOR2X1_LOC_653/B NOR2X1_LOC_92/Y 0.02fF
C54870 INVX1_LOC_201/Y NOR2X1_LOC_554/A 0.04fF
C54871 VDD NOR2X1_LOC_114/A 0.24fF
C54872 NAND2X1_LOC_721/B NOR2X1_LOC_654/A 0.19fF
C54873 NOR2X1_LOC_15/Y INVX1_LOC_27/A 0.18fF
C54874 INVX1_LOC_279/A INVX1_LOC_84/A 0.07fF
C54875 NAND2X1_LOC_59/B NAND2X1_LOC_3/B 0.35fF
C54876 NOR2X1_LOC_778/B INVX1_LOC_99/A 0.04fF
C54877 NOR2X1_LOC_15/Y NOR2X1_LOC_824/A 0.06fF
C54878 INVX1_LOC_10/A NAND2X1_LOC_475/Y 0.03fF
C54879 NOR2X1_LOC_78/A NOR2X1_LOC_137/Y 0.03fF
C54880 VDD INVX1_LOC_91/A 6.54fF
C54881 INVX1_LOC_257/Y INVX1_LOC_257/A 0.03fF
C54882 NAND2X1_LOC_468/B NAND2X1_LOC_274/a_36_24# 0.00fF
C54883 INVX1_LOC_176/A NAND2X1_LOC_642/Y 0.01fF
C54884 INVX1_LOC_64/A NAND2X1_LOC_711/Y 0.07fF
C54885 INVX1_LOC_315/Y NAND2X1_LOC_8/a_36_24# 0.00fF
C54886 NAND2X1_LOC_579/A NAND2X1_LOC_725/B 0.07fF
C54887 INVX1_LOC_58/A NAND2X1_LOC_355/Y 0.05fF
C54888 INVX1_LOC_36/A NOR2X1_LOC_717/A 0.31fF
C54889 NOR2X1_LOC_208/Y NOR2X1_LOC_727/B 0.00fF
C54890 INVX1_LOC_17/A NOR2X1_LOC_763/A 0.45fF
C54891 NOR2X1_LOC_544/A NOR2X1_LOC_850/B 0.01fF
C54892 INVX1_LOC_24/Y NOR2X1_LOC_793/A 0.31fF
C54893 VDD INVX1_LOC_11/Y 0.69fF
C54894 NOR2X1_LOC_501/a_36_216# INVX1_LOC_29/A 0.00fF
C54895 NAND2X1_LOC_244/A INVX1_LOC_20/A 0.00fF
C54896 NAND2X1_LOC_241/Y INVX1_LOC_46/A 0.01fF
C54897 INVX1_LOC_35/A INVX1_LOC_61/A 0.07fF
C54898 NOR2X1_LOC_92/Y NAND2X1_LOC_550/A 0.09fF
C54899 INVX1_LOC_25/Y INVX1_LOC_19/Y 0.09fF
C54900 NAND2X1_LOC_79/a_36_24# NAND2X1_LOC_215/A 0.00fF
C54901 INVX1_LOC_256/A NOR2X1_LOC_122/A 0.01fF
C54902 INVX1_LOC_36/A NOR2X1_LOC_649/Y 0.07fF
C54903 NOR2X1_LOC_391/Y NOR2X1_LOC_78/Y 0.01fF
C54904 D_INPUT_0 NAND2X1_LOC_74/B 0.20fF
C54905 NAND2X1_LOC_531/a_36_24# INVX1_LOC_29/A 0.00fF
C54906 NAND2X1_LOC_713/a_36_24# NAND2X1_LOC_550/A 0.00fF
C54907 INVX1_LOC_24/Y NOR2X1_LOC_160/B 0.10fF
C54908 INVX1_LOC_182/Y INVX1_LOC_84/A 0.03fF
C54909 NOR2X1_LOC_448/B INVX1_LOC_174/A 0.02fF
C54910 NAND2X1_LOC_858/B NOR2X1_LOC_88/Y 0.73fF
C54911 INVX1_LOC_30/A NAND2X1_LOC_474/Y 0.10fF
C54912 NOR2X1_LOC_322/Y INVX1_LOC_119/Y 0.21fF
C54913 NAND2X1_LOC_468/B NAND2X1_LOC_61/a_36_24# 0.00fF
C54914 NAND2X1_LOC_354/B INVX1_LOC_57/A 0.46fF
C54915 NAND2X1_LOC_662/Y NOR2X1_LOC_467/A 0.01fF
C54916 INVX1_LOC_21/A NOR2X1_LOC_274/B 0.20fF
C54917 INVX1_LOC_11/A INVX1_LOC_225/Y 0.09fF
C54918 INVX1_LOC_256/A INVX1_LOC_161/Y 0.10fF
C54919 INVX1_LOC_103/A NOR2X1_LOC_45/Y 0.07fF
C54920 INVX1_LOC_236/Y NAND2X1_LOC_537/Y 0.01fF
C54921 VDD NOR2X1_LOC_698/Y 0.27fF
C54922 NOR2X1_LOC_441/Y INVX1_LOC_88/A 0.05fF
C54923 INVX1_LOC_212/A INVX1_LOC_50/Y 0.02fF
C54924 INVX1_LOC_6/A NOR2X1_LOC_697/Y 0.01fF
C54925 INVX1_LOC_233/A NAND2X1_LOC_833/Y 0.50fF
C54926 NAND2X1_LOC_549/Y NAND2X1_LOC_549/a_36_24# 0.02fF
C54927 NOR2X1_LOC_35/Y INVX1_LOC_9/A 0.32fF
C54928 INVX1_LOC_58/A INVX1_LOC_304/Y 0.03fF
C54929 NOR2X1_LOC_352/a_36_216# NOR2X1_LOC_155/A 0.00fF
C54930 NOR2X1_LOC_569/Y NOR2X1_LOC_334/Y 0.00fF
C54931 INVX1_LOC_35/A NOR2X1_LOC_624/A 0.09fF
C54932 NOR2X1_LOC_309/Y NOR2X1_LOC_717/A 0.01fF
C54933 INVX1_LOC_79/A INVX1_LOC_133/A 0.21fF
C54934 INVX1_LOC_27/A NOR2X1_LOC_860/B 0.07fF
C54935 INVX1_LOC_17/A INVX1_LOC_57/Y 0.07fF
C54936 NAND2X1_LOC_53/Y INVX1_LOC_30/A 0.07fF
C54937 INVX1_LOC_244/A NOR2X1_LOC_48/B 0.14fF
C54938 NOR2X1_LOC_220/B NOR2X1_LOC_593/Y 0.05fF
C54939 NOR2X1_LOC_205/Y NOR2X1_LOC_270/Y 0.12fF
C54940 NAND2X1_LOC_709/a_36_24# NOR2X1_LOC_833/B 0.00fF
C54941 INVX1_LOC_21/A NOR2X1_LOC_577/Y 0.08fF
C54942 INVX1_LOC_89/A INVX1_LOC_4/A 5.45fF
C54943 NAND2X1_LOC_579/A INVX1_LOC_309/Y -0.01fF
C54944 NAND2X1_LOC_325/Y NOR2X1_LOC_406/A 0.17fF
C54945 INVX1_LOC_69/Y INVX1_LOC_19/A 0.01fF
C54946 NOR2X1_LOC_647/A INVX1_LOC_13/A 0.08fF
C54947 NOR2X1_LOC_254/Y INVX1_LOC_50/Y 0.94fF
C54948 NOR2X1_LOC_773/Y INVX1_LOC_29/Y 0.31fF
C54949 INVX1_LOC_58/A NOR2X1_LOC_566/Y 0.02fF
C54950 NOR2X1_LOC_67/A NAND2X1_LOC_571/B 0.03fF
C54951 NOR2X1_LOC_488/Y INVX1_LOC_57/A 0.03fF
C54952 NOR2X1_LOC_137/A INVX1_LOC_94/Y 0.03fF
C54953 INVX1_LOC_266/A NOR2X1_LOC_303/Y 0.10fF
C54954 INVX1_LOC_269/A INVX1_LOC_94/A 0.42fF
C54955 INVX1_LOC_2/A NOR2X1_LOC_423/a_36_216# 0.00fF
C54956 INVX1_LOC_249/A NOR2X1_LOC_15/Y 0.01fF
C54957 INVX1_LOC_299/A NAND2X1_LOC_84/Y 0.00fF
C54958 NAND2X1_LOC_773/Y NOR2X1_LOC_262/Y 0.05fF
C54959 INVX1_LOC_24/A NAND2X1_LOC_538/Y 0.07fF
C54960 INVX1_LOC_17/A NOR2X1_LOC_512/Y 0.01fF
C54961 NOR2X1_LOC_647/Y INPUT_3 0.00fF
C54962 INVX1_LOC_233/A INVX1_LOC_164/Y 0.04fF
C54963 NAND2X1_LOC_703/Y NAND2X1_LOC_833/Y 0.01fF
C54964 INVX1_LOC_256/A NOR2X1_LOC_276/a_36_216# 0.00fF
C54965 NOR2X1_LOC_632/Y INVX1_LOC_50/A 0.06fF
C54966 INVX1_LOC_24/A NOR2X1_LOC_250/A 0.00fF
C54967 INVX1_LOC_135/A INVX1_LOC_26/A 0.50fF
C54968 NOR2X1_LOC_725/A INVX1_LOC_19/A 0.16fF
C54969 NOR2X1_LOC_655/B NOR2X1_LOC_772/B 0.10fF
C54970 NAND2X1_LOC_222/B NOR2X1_LOC_643/Y 0.02fF
C54971 NAND2X1_LOC_392/A NAND2X1_LOC_860/A 0.02fF
C54972 INVX1_LOC_133/A INVX1_LOC_91/A 0.02fF
C54973 INVX1_LOC_110/Y NOR2X1_LOC_68/A 0.04fF
C54974 INVX1_LOC_311/A INVX1_LOC_283/A 0.05fF
C54975 INVX1_LOC_117/A INVX1_LOC_92/A 0.21fF
C54976 INVX1_LOC_41/A NOR2X1_LOC_793/A 0.07fF
C54977 INVX1_LOC_243/Y NOR2X1_LOC_763/Y 0.16fF
C54978 NAND2X1_LOC_550/a_36_24# NAND2X1_LOC_860/A 0.01fF
C54979 INVX1_LOC_227/A INVX1_LOC_57/A 0.07fF
C54980 NAND2X1_LOC_555/Y NOR2X1_LOC_480/A 0.00fF
C54981 NAND2X1_LOC_659/B INVX1_LOC_203/A 0.08fF
C54982 INVX1_LOC_185/A INVX1_LOC_38/A 0.03fF
C54983 INVX1_LOC_27/A NAND2X1_LOC_141/A 0.03fF
C54984 INVX1_LOC_125/Y NOR2X1_LOC_89/A 0.33fF
C54985 NOR2X1_LOC_655/B INVX1_LOC_13/Y 0.01fF
C54986 NOR2X1_LOC_111/Y INVX1_LOC_78/A 0.01fF
C54987 NOR2X1_LOC_598/B NAND2X1_LOC_41/Y 0.01fF
C54988 VDD NOR2X1_LOC_179/Y 0.25fF
C54989 INVX1_LOC_88/A NOR2X1_LOC_142/Y 0.05fF
C54990 NOR2X1_LOC_381/Y NOR2X1_LOC_84/A 0.10fF
C54991 NAND2X1_LOC_149/Y NAND2X1_LOC_629/Y 0.04fF
C54992 NAND2X1_LOC_565/B NAND2X1_LOC_569/B 0.03fF
C54993 NOR2X1_LOC_178/Y INVX1_LOC_53/Y 0.12fF
C54994 INVX1_LOC_2/A NAND2X1_LOC_714/B 0.03fF
C54995 INVX1_LOC_1/A INVX1_LOC_85/A 0.09fF
C54996 INVX1_LOC_58/A NAND2X1_LOC_808/A -0.02fF
C54997 NAND2X1_LOC_650/B NOR2X1_LOC_662/A 0.02fF
C54998 NAND2X1_LOC_787/A INVX1_LOC_10/A 0.03fF
C54999 NOR2X1_LOC_255/Y INVX1_LOC_135/A 0.10fF
C55000 NOR2X1_LOC_232/Y NOR2X1_LOC_234/Y 0.01fF
C55001 INVX1_LOC_225/Y NOR2X1_LOC_593/Y 0.04fF
C55002 INVX1_LOC_14/A NOR2X1_LOC_315/Y 0.28fF
C55003 VDD INVX1_LOC_203/A 1.36fF
C55004 NOR2X1_LOC_15/Y INVX1_LOC_206/A 0.72fF
C55005 INVX1_LOC_267/Y INVX1_LOC_163/A 0.01fF
C55006 NAND2X1_LOC_149/Y INVX1_LOC_243/A 0.02fF
C55007 INVX1_LOC_27/A INVX1_LOC_226/A 0.03fF
C55008 NOR2X1_LOC_536/A NOR2X1_LOC_841/A 0.16fF
C55009 NOR2X1_LOC_498/Y NAND2X1_LOC_550/A 0.17fF
C55010 NOR2X1_LOC_658/Y NOR2X1_LOC_208/Y 0.02fF
C55011 INVX1_LOC_226/Y NOR2X1_LOC_791/Y 0.01fF
C55012 INVX1_LOC_36/A NOR2X1_LOC_13/Y 0.00fF
C55013 INVX1_LOC_41/A NOR2X1_LOC_160/B 0.29fF
C55014 INVX1_LOC_39/A NOR2X1_LOC_121/A 0.05fF
C55015 INVX1_LOC_201/Y NOR2X1_LOC_160/B 0.07fF
C55016 D_INPUT_0 NOR2X1_LOC_660/Y 0.04fF
C55017 NAND2X1_LOC_9/Y NOR2X1_LOC_76/A 0.07fF
C55018 NOR2X1_LOC_45/B D_INPUT_5 0.03fF
C55019 INVX1_LOC_21/A INVX1_LOC_22/A 0.27fF
C55020 INVX1_LOC_235/Y NOR2X1_LOC_375/Y 0.03fF
C55021 INVX1_LOC_11/A INVX1_LOC_266/Y 0.08fF
C55022 NAND2X1_LOC_469/B INVX1_LOC_109/Y 0.12fF
C55023 NAND2X1_LOC_741/B NOR2X1_LOC_387/Y 0.01fF
C55024 INVX1_LOC_107/Y INVX1_LOC_54/A 0.04fF
C55025 NOR2X1_LOC_15/Y NAND2X1_LOC_200/B 0.01fF
C55026 NAND2X1_LOC_633/Y INVX1_LOC_29/A 0.07fF
C55027 NAND2X1_LOC_569/B NOR2X1_LOC_130/A 1.95fF
C55028 INVX1_LOC_108/Y NAND2X1_LOC_815/a_36_24# 0.00fF
C55029 NOR2X1_LOC_296/Y INVX1_LOC_34/Y 0.17fF
C55030 D_INPUT_3 NOR2X1_LOC_671/a_36_216# 0.00fF
C55031 INVX1_LOC_64/A INVX1_LOC_89/A 0.23fF
C55032 INVX1_LOC_250/A NOR2X1_LOC_753/Y 0.07fF
C55033 NOR2X1_LOC_241/A INVX1_LOC_196/A 0.09fF
C55034 NOR2X1_LOC_208/A NOR2X1_LOC_727/B 0.31fF
C55035 NOR2X1_LOC_78/A NOR2X1_LOC_227/A 0.01fF
C55036 NOR2X1_LOC_453/Y INVX1_LOC_22/A 0.00fF
C55037 NOR2X1_LOC_716/B NOR2X1_LOC_82/a_36_216# 0.01fF
C55038 INVX1_LOC_36/A NAND2X1_LOC_175/B 0.07fF
C55039 NOR2X1_LOC_454/Y INVX1_LOC_290/A 2.31fF
C55040 NOR2X1_LOC_35/Y NOR2X1_LOC_861/Y 0.10fF
C55041 NOR2X1_LOC_716/B NAND2X1_LOC_634/Y 0.01fF
C55042 INVX1_LOC_24/Y NOR2X1_LOC_516/B 0.11fF
C55043 INVX1_LOC_2/Y INVX1_LOC_42/A 0.06fF
C55044 NOR2X1_LOC_410/Y INVX1_LOC_33/A 0.03fF
C55045 NAND2X1_LOC_639/A INPUT_7 0.03fF
C55046 NOR2X1_LOC_592/B NOR2X1_LOC_832/a_36_216# 0.00fF
C55047 INVX1_LOC_246/Y NOR2X1_LOC_433/A 0.01fF
C55048 INVX1_LOC_214/Y INVX1_LOC_215/Y 0.02fF
C55049 NOR2X1_LOC_457/A NOR2X1_LOC_500/Y 0.07fF
C55050 INVX1_LOC_55/Y INVX1_LOC_298/A 0.02fF
C55051 NOR2X1_LOC_283/a_36_216# INVX1_LOC_314/Y 0.01fF
C55052 INVX1_LOC_233/A INVX1_LOC_73/A 0.04fF
C55053 NAND2X1_LOC_425/Y NAND2X1_LOC_426/a_36_24# 0.00fF
C55054 NOR2X1_LOC_336/B NOR2X1_LOC_175/A 0.06fF
C55055 NOR2X1_LOC_15/Y INVX1_LOC_234/A 0.07fF
C55056 INVX1_LOC_5/A NOR2X1_LOC_736/Y 0.08fF
C55057 NAND2X1_LOC_802/A NOR2X1_LOC_433/A 0.00fF
C55058 INVX1_LOC_135/A NOR2X1_LOC_560/a_36_216# 0.00fF
C55059 INVX1_LOC_36/A NOR2X1_LOC_504/Y 1.06fF
C55060 INVX1_LOC_289/A NAND2X1_LOC_509/a_36_24# 0.00fF
C55061 INVX1_LOC_49/A NOR2X1_LOC_550/B 0.03fF
C55062 NOR2X1_LOC_140/A NOR2X1_LOC_130/A 0.06fF
C55063 NOR2X1_LOC_598/a_36_216# INVX1_LOC_104/A 0.02fF
C55064 VDD INVX1_LOC_231/A -0.00fF
C55065 NOR2X1_LOC_400/A INVX1_LOC_75/A 0.02fF
C55066 NOR2X1_LOC_460/B INVX1_LOC_77/A 0.00fF
C55067 INVX1_LOC_54/A INVX1_LOC_272/A 0.14fF
C55068 NOR2X1_LOC_703/B INVX1_LOC_177/A 0.01fF
C55069 INVX1_LOC_293/Y INVX1_LOC_46/Y 2.15fF
C55070 NAND2X1_LOC_783/A NAND2X1_LOC_538/Y 0.10fF
C55071 INVX1_LOC_34/A INVX1_LOC_314/Y 0.03fF
C55072 NOR2X1_LOC_428/Y INVX1_LOC_22/A 0.15fF
C55073 NAND2X1_LOC_800/A INVX1_LOC_231/A 0.85fF
C55074 INVX1_LOC_36/A INVX1_LOC_256/Y 0.25fF
C55075 NOR2X1_LOC_820/a_36_216# INVX1_LOC_63/A 0.00fF
C55076 NOR2X1_LOC_74/A NOR2X1_LOC_665/Y 0.54fF
C55077 NOR2X1_LOC_408/a_36_216# INPUT_5 0.00fF
C55078 INVX1_LOC_305/A NAND2X1_LOC_690/a_36_24# 0.00fF
C55079 NOR2X1_LOC_645/a_36_216# INVX1_LOC_2/A 0.00fF
C55080 NOR2X1_LOC_419/Y INVX1_LOC_8/A 0.11fF
C55081 NOR2X1_LOC_640/Y NOR2X1_LOC_633/A 0.01fF
C55082 INVX1_LOC_13/Y NAND2X1_LOC_102/a_36_24# 0.01fF
C55083 INVX1_LOC_24/A NOR2X1_LOC_709/A 0.00fF
C55084 INVX1_LOC_30/A NOR2X1_LOC_500/Y 0.05fF
C55085 INVX1_LOC_226/Y INVX1_LOC_30/A 0.00fF
C55086 INVX1_LOC_2/A NOR2X1_LOC_273/Y 0.07fF
C55087 NOR2X1_LOC_250/A NOR2X1_LOC_130/A 0.03fF
C55088 NOR2X1_LOC_716/B INVX1_LOC_8/A 0.16fF
C55089 INVX1_LOC_125/A NOR2X1_LOC_197/B 0.09fF
C55090 INVX1_LOC_46/Y NAND2X1_LOC_74/B 0.17fF
C55091 INVX1_LOC_2/A NOR2X1_LOC_759/Y 0.05fF
C55092 NOR2X1_LOC_790/B INVX1_LOC_186/A 0.93fF
C55093 NOR2X1_LOC_15/Y NOR2X1_LOC_772/A 0.00fF
C55094 NOR2X1_LOC_246/A NAND2X1_LOC_793/Y 0.01fF
C55095 INVX1_LOC_249/A INVX1_LOC_96/Y 0.09fF
C55096 NOR2X1_LOC_15/Y NOR2X1_LOC_19/B 0.03fF
C55097 INVX1_LOC_78/A INVX1_LOC_37/Y 0.00fF
C55098 NOR2X1_LOC_433/A INVX1_LOC_266/Y 0.01fF
C55099 INVX1_LOC_104/A INVX1_LOC_155/A 0.05fF
C55100 NAND2X1_LOC_312/a_36_24# NOR2X1_LOC_703/A 0.02fF
C55101 NOR2X1_LOC_517/Y INVX1_LOC_22/A 0.17fF
C55102 INVX1_LOC_136/A NAND2X1_LOC_727/Y 0.01fF
C55103 NOR2X1_LOC_658/a_36_216# NOR2X1_LOC_357/Y 0.00fF
C55104 INVX1_LOC_202/Y NAND2X1_LOC_454/Y 0.01fF
C55105 D_INPUT_1 INVX1_LOC_95/Y 0.19fF
C55106 NAND2X1_LOC_287/B NAND2X1_LOC_286/B 0.09fF
C55107 NOR2X1_LOC_631/B INVX1_LOC_23/A 0.43fF
C55108 NAND2X1_LOC_564/B INVX1_LOC_18/A 0.07fF
C55109 INVX1_LOC_303/A NOR2X1_LOC_655/B 0.10fF
C55110 NOR2X1_LOC_91/A INVX1_LOC_37/A 0.03fF
C55111 NOR2X1_LOC_593/Y INVX1_LOC_266/Y 0.01fF
C55112 INVX1_LOC_136/A NAND2X1_LOC_660/Y 1.22fF
C55113 NOR2X1_LOC_197/A INVX1_LOC_85/Y 0.01fF
C55114 NOR2X1_LOC_89/A NAND2X1_LOC_288/A 0.01fF
C55115 INVX1_LOC_30/A INVX1_LOC_10/A 1.26fF
C55116 NOR2X1_LOC_557/Y NOR2X1_LOC_709/A 0.10fF
C55117 INVX1_LOC_214/A NOR2X1_LOC_577/Y 0.06fF
C55118 NOR2X1_LOC_273/Y NOR2X1_LOC_218/Y 0.01fF
C55119 NAND2X1_LOC_798/A NAND2X1_LOC_593/Y 0.00fF
C55120 INVX1_LOC_27/A NOR2X1_LOC_733/Y 0.03fF
C55121 NOR2X1_LOC_667/A NOR2X1_LOC_577/Y 0.00fF
C55122 NOR2X1_LOC_813/Y INVX1_LOC_26/A 0.04fF
C55123 NOR2X1_LOC_667/Y INVX1_LOC_90/A 0.02fF
C55124 NOR2X1_LOC_218/Y NOR2X1_LOC_759/Y 0.02fF
C55125 NAND2X1_LOC_850/a_36_24# NAND2X1_LOC_850/Y 0.03fF
C55126 NOR2X1_LOC_361/B INVX1_LOC_79/A 0.11fF
C55127 NAND2X1_LOC_218/B NAND2X1_LOC_6/a_36_24# 0.00fF
C55128 NOR2X1_LOC_99/B NOR2X1_LOC_500/B 0.04fF
C55129 INVX1_LOC_202/A NOR2X1_LOC_218/Y 0.06fF
C55130 NAND2X1_LOC_778/Y NOR2X1_LOC_528/Y 0.15fF
C55131 INVX1_LOC_70/Y INVX1_LOC_306/Y 0.01fF
C55132 NOR2X1_LOC_814/A NOR2X1_LOC_33/B 0.06fF
C55133 NOR2X1_LOC_510/Y INVX1_LOC_91/A 0.07fF
C55134 NOR2X1_LOC_52/B INVX1_LOC_266/Y 0.00fF
C55135 INVX1_LOC_136/A D_INPUT_0 0.39fF
C55136 NOR2X1_LOC_392/Y INVX1_LOC_20/A 0.08fF
C55137 INVX1_LOC_26/A INVX1_LOC_280/A 0.02fF
C55138 INVX1_LOC_37/A INVX1_LOC_23/A 0.80fF
C55139 NOR2X1_LOC_544/A NOR2X1_LOC_551/B 0.01fF
C55140 NOR2X1_LOC_716/B NOR2X1_LOC_315/a_36_216# 0.01fF
C55141 INVX1_LOC_64/A NOR2X1_LOC_24/Y 0.00fF
C55142 INVX1_LOC_232/Y NOR2X1_LOC_516/Y 0.01fF
C55143 NAND2X1_LOC_574/A NOR2X1_LOC_554/A 0.03fF
C55144 INVX1_LOC_290/A INVX1_LOC_77/A 0.07fF
C55145 NOR2X1_LOC_726/a_36_216# INVX1_LOC_213/A 0.01fF
C55146 INVX1_LOC_174/A INVX1_LOC_75/A 0.14fF
C55147 INVX1_LOC_35/A D_INPUT_3 0.11fF
C55148 INVX1_LOC_95/Y NOR2X1_LOC_652/Y 0.00fF
C55149 INVX1_LOC_136/A NOR2X1_LOC_389/a_36_216# 0.00fF
C55150 INVX1_LOC_41/A NOR2X1_LOC_516/B 0.04fF
C55151 NOR2X1_LOC_471/Y NOR2X1_LOC_74/Y 0.04fF
C55152 NOR2X1_LOC_89/A INVX1_LOC_19/A 0.48fF
C55153 INVX1_LOC_35/A INVX1_LOC_14/Y 0.01fF
C55154 NOR2X1_LOC_255/Y NOR2X1_LOC_813/Y 0.37fF
C55155 INVX1_LOC_143/A NOR2X1_LOC_709/A 0.17fF
C55156 NOR2X1_LOC_15/Y NOR2X1_LOC_528/Y 0.03fF
C55157 NOR2X1_LOC_603/a_36_216# INVX1_LOC_266/Y 0.01fF
C55158 NOR2X1_LOC_151/Y NOR2X1_LOC_181/a_36_216# 0.00fF
C55159 INVX1_LOC_53/A INVX1_LOC_117/A 0.21fF
C55160 NAND2X1_LOC_787/A NOR2X1_LOC_301/a_36_216# 0.00fF
C55161 NOR2X1_LOC_331/B NAND2X1_LOC_201/a_36_24# 0.01fF
C55162 NAND2X1_LOC_351/a_36_24# INVX1_LOC_37/A 0.01fF
C55163 INVX1_LOC_45/A NOR2X1_LOC_256/Y 0.01fF
C55164 NOR2X1_LOC_361/B INVX1_LOC_91/A 0.10fF
C55165 NOR2X1_LOC_255/Y INVX1_LOC_280/A 0.01fF
C55166 NAND2X1_LOC_470/B NOR2X1_LOC_841/A 0.07fF
C55167 NOR2X1_LOC_91/A NOR2X1_LOC_743/Y 0.00fF
C55168 INVX1_LOC_84/A NOR2X1_LOC_38/B 0.11fF
C55169 NAND2X1_LOC_740/B NAND2X1_LOC_856/A 0.64fF
C55170 NOR2X1_LOC_620/Y INVX1_LOC_83/A 0.03fF
C55171 NAND2X1_LOC_303/Y INPUT_4 0.16fF
C55172 INVX1_LOC_38/A NOR2X1_LOC_754/Y 0.00fF
C55173 NOR2X1_LOC_78/B NAND2X1_LOC_181/Y 0.03fF
C55174 INVX1_LOC_179/A NOR2X1_LOC_302/A 0.01fF
C55175 NAND2X1_LOC_736/Y INVX1_LOC_229/Y 0.64fF
C55176 INVX1_LOC_289/A INVX1_LOC_191/Y 0.00fF
C55177 INVX1_LOC_1/A INVX1_LOC_314/A 0.03fF
C55178 NOR2X1_LOC_409/B NAND2X1_LOC_407/a_36_24# 0.02fF
C55179 NAND2X1_LOC_149/Y INVX1_LOC_76/A 0.34fF
C55180 NOR2X1_LOC_425/a_36_216# INPUT_5 0.02fF
C55181 INVX1_LOC_223/A NOR2X1_LOC_188/A 0.77fF
C55182 NOR2X1_LOC_15/Y NOR2X1_LOC_314/a_36_216# 0.00fF
C55183 NOR2X1_LOC_1/Y D_INPUT_5 0.01fF
C55184 INVX1_LOC_23/A NOR2X1_LOC_743/Y 0.03fF
C55185 NOR2X1_LOC_329/B NOR2X1_LOC_106/Y 0.04fF
C55186 NOR2X1_LOC_667/A INVX1_LOC_22/A 0.11fF
C55187 INVX1_LOC_58/A INVX1_LOC_92/A 0.22fF
C55188 INVX1_LOC_295/A INVX1_LOC_103/Y 0.03fF
C55189 NOR2X1_LOC_111/Y NOR2X1_LOC_152/Y 0.04fF
C55190 NOR2X1_LOC_592/A NOR2X1_LOC_56/Y -0.01fF
C55191 NOR2X1_LOC_242/A INVX1_LOC_117/A 0.01fF
C55192 NOR2X1_LOC_196/A NOR2X1_LOC_196/Y 0.01fF
C55193 INVX1_LOC_83/A NOR2X1_LOC_731/A 0.52fF
C55194 NAND2X1_LOC_708/Y INVX1_LOC_54/A 0.08fF
C55195 NOR2X1_LOC_149/a_36_216# INVX1_LOC_213/A 0.01fF
C55196 NAND2X1_LOC_722/A INVX1_LOC_10/A 0.07fF
C55197 INVX1_LOC_15/Y INVX1_LOC_234/A 0.07fF
C55198 NOR2X1_LOC_67/A NOR2X1_LOC_789/a_36_216# 0.00fF
C55199 NAND2X1_LOC_327/a_36_24# NOR2X1_LOC_577/Y 0.00fF
C55200 NAND2X1_LOC_181/Y NAND2X1_LOC_392/Y 0.21fF
C55201 INVX1_LOC_16/A NOR2X1_LOC_719/A 0.15fF
C55202 NOR2X1_LOC_739/Y VDD 0.36fF
C55203 NOR2X1_LOC_292/Y INVX1_LOC_71/A 0.28fF
C55204 INVX1_LOC_314/Y INPUT_0 0.19fF
C55205 NOR2X1_LOC_468/Y NOR2X1_LOC_440/a_36_216# 0.00fF
C55206 NAND2X1_LOC_349/B NOR2X1_LOC_589/A 0.43fF
C55207 INVX1_LOC_34/A NOR2X1_LOC_597/Y 0.09fF
C55208 INVX1_LOC_89/A INVX1_LOC_44/Y 0.01fF
C55209 INVX1_LOC_18/Y INVX1_LOC_69/A 0.01fF
C55210 NOR2X1_LOC_599/Y INVX1_LOC_20/A 0.07fF
C55211 NOR2X1_LOC_560/a_36_216# INVX1_LOC_280/A 0.00fF
C55212 NOR2X1_LOC_561/Y INVX1_LOC_16/A 0.10fF
C55213 NAND2X1_LOC_714/B INVX1_LOC_118/A 0.03fF
C55214 NOR2X1_LOC_703/B INVX1_LOC_65/A 0.01fF
C55215 NAND2X1_LOC_337/B NOR2X1_LOC_111/A 0.11fF
C55216 NOR2X1_LOC_19/B NAND2X1_LOC_141/A 0.08fF
C55217 NOR2X1_LOC_795/Y NOR2X1_LOC_567/B 0.10fF
C55218 INVX1_LOC_49/A NOR2X1_LOC_334/A 0.02fF
C55219 INVX1_LOC_15/Y NOR2X1_LOC_19/B 2.84fF
C55220 INVX1_LOC_96/A NOR2X1_LOC_303/Y 0.03fF
C55221 INVX1_LOC_83/Y INVX1_LOC_85/Y 0.01fF
C55222 INVX1_LOC_31/A NOR2X1_LOC_681/Y 0.29fF
C55223 INVX1_LOC_31/A INVX1_LOC_37/A 0.07fF
C55224 NOR2X1_LOC_631/a_36_216# NOR2X1_LOC_631/Y 0.02fF
C55225 NAND2X1_LOC_561/B INVX1_LOC_118/A 0.00fF
C55226 NOR2X1_LOC_86/Y INVX1_LOC_20/A 0.01fF
C55227 INVX1_LOC_208/A NOR2X1_LOC_122/Y 0.02fF
C55228 INVX1_LOC_255/Y INVX1_LOC_20/Y 0.02fF
C55229 NOR2X1_LOC_372/Y VDD 0.12fF
C55230 NOR2X1_LOC_554/B INVX1_LOC_2/Y 0.03fF
C55231 NAND2X1_LOC_633/Y NAND2X1_LOC_634/Y 0.02fF
C55232 INVX1_LOC_207/A NOR2X1_LOC_45/B 0.09fF
C55233 NOR2X1_LOC_647/A INVX1_LOC_32/A 0.01fF
C55234 NOR2X1_LOC_667/Y INVX1_LOC_38/A 0.02fF
C55235 NOR2X1_LOC_602/A INVX1_LOC_33/Y 0.15fF
C55236 NOR2X1_LOC_614/Y NOR2X1_LOC_567/B 0.02fF
C55237 NAND2X1_LOC_787/A INVX1_LOC_12/A 0.03fF
C55238 INVX1_LOC_35/A NOR2X1_LOC_831/Y 0.30fF
C55239 NOR2X1_LOC_15/Y NOR2X1_LOC_216/B 0.03fF
C55240 INVX1_LOC_63/A NOR2X1_LOC_649/Y 0.14fF
C55241 NOR2X1_LOC_744/Y INVX1_LOC_76/A 0.03fF
C55242 INVX1_LOC_150/Y INVX1_LOC_54/A 0.09fF
C55243 NOR2X1_LOC_778/B INPUT_0 0.03fF
C55244 NOR2X1_LOC_763/A NOR2X1_LOC_430/Y 0.02fF
C55245 NAND2X1_LOC_720/a_36_24# INVX1_LOC_33/Y -0.00fF
C55246 NAND2X1_LOC_342/Y NOR2X1_LOC_9/Y 0.02fF
C55247 INVX1_LOC_244/Y VDD 0.70fF
C55248 INPUT_3 NOR2X1_LOC_860/Y 0.01fF
C55249 NOR2X1_LOC_561/Y INVX1_LOC_28/A 0.17fF
C55250 NOR2X1_LOC_457/A INVX1_LOC_307/A 0.08fF
C55251 NOR2X1_LOC_590/A INVX1_LOC_274/A 0.51fF
C55252 INVX1_LOC_280/Y INVX1_LOC_309/A 0.03fF
C55253 INVX1_LOC_21/A INVX1_LOC_186/Y 0.03fF
C55254 INVX1_LOC_136/A NAND2X1_LOC_848/A 0.07fF
C55255 NOR2X1_LOC_457/A NOR2X1_LOC_445/B 0.14fF
C55256 NOR2X1_LOC_589/A INVX1_LOC_75/A 0.03fF
C55257 INVX1_LOC_177/A INVX1_LOC_91/A 0.03fF
C55258 NOR2X1_LOC_471/Y INVX1_LOC_179/A 0.02fF
C55259 NAND2X1_LOC_53/Y INVX1_LOC_113/A 0.37fF
C55260 INVX1_LOC_211/Y NAND2X1_LOC_798/B 0.50fF
C55261 NOR2X1_LOC_15/Y NAND2X1_LOC_477/Y 0.19fF
C55262 INVX1_LOC_311/A INVX1_LOC_22/A 0.08fF
C55263 NAND2X1_LOC_190/Y INVX1_LOC_84/A 0.07fF
C55264 NOR2X1_LOC_383/B INVX1_LOC_94/Y 0.05fF
C55265 NOR2X1_LOC_705/B NAND2X1_LOC_425/Y 0.01fF
C55266 INVX1_LOC_45/A NOR2X1_LOC_641/Y 0.00fF
C55267 INVX1_LOC_18/A NOR2X1_LOC_261/A 0.03fF
C55268 NAND2X1_LOC_687/A NOR2X1_LOC_152/Y 0.03fF
C55269 NOR2X1_LOC_219/B INVX1_LOC_139/A 0.10fF
C55270 NAND2X1_LOC_736/Y INVX1_LOC_20/A 0.04fF
C55271 NOR2X1_LOC_568/A NOR2X1_LOC_641/Y 0.00fF
C55272 NOR2X1_LOC_174/B INVX1_LOC_148/A 0.00fF
C55273 NOR2X1_LOC_307/Y NOR2X1_LOC_727/B 0.21fF
C55274 INVX1_LOC_199/A INVX1_LOC_266/Y 0.07fF
C55275 INVX1_LOC_71/A INVX1_LOC_44/A 0.08fF
C55276 NAND2X1_LOC_348/A NOR2X1_LOC_349/B 0.01fF
C55277 NAND2X1_LOC_276/Y VDD 0.42fF
C55278 NAND2X1_LOC_724/Y NAND2X1_LOC_175/Y 2.53fF
C55279 NOR2X1_LOC_392/Y INVX1_LOC_4/A 0.07fF
C55280 INVX1_LOC_11/A NOR2X1_LOC_653/Y 0.03fF
C55281 INVX1_LOC_78/A INVX1_LOC_29/Y 0.03fF
C55282 NOR2X1_LOC_160/B NAND2X1_LOC_574/A 0.10fF
C55283 INVX1_LOC_23/A NAND2X1_LOC_72/B 0.03fF
C55284 INVX1_LOC_30/A INVX1_LOC_307/A 0.18fF
C55285 NOR2X1_LOC_454/Y INVX1_LOC_261/Y 0.04fF
C55286 INVX1_LOC_98/A INVX1_LOC_56/Y 0.03fF
C55287 NOR2X1_LOC_657/Y NOR2X1_LOC_364/A 0.01fF
C55288 INVX1_LOC_280/Y INVX1_LOC_11/Y 0.03fF
C55289 NAND2X1_LOC_717/Y NOR2X1_LOC_824/Y 0.01fF
C55290 NOR2X1_LOC_591/Y NOR2X1_LOC_305/Y 0.08fF
C55291 INVX1_LOC_224/A INVX1_LOC_19/A 0.03fF
C55292 NOR2X1_LOC_298/Y NOR2X1_LOC_387/A 0.03fF
C55293 INVX1_LOC_30/A NOR2X1_LOC_445/B 0.10fF
C55294 NAND2X1_LOC_349/a_36_24# NOR2X1_LOC_318/B 0.00fF
C55295 INVX1_LOC_136/A INVX1_LOC_46/Y 0.10fF
C55296 NOR2X1_LOC_553/B NOR2X1_LOC_337/Y 0.02fF
C55297 INVX1_LOC_257/Y INVX1_LOC_14/Y 0.34fF
C55298 INVX1_LOC_11/A INVX1_LOC_19/A 0.18fF
C55299 NOR2X1_LOC_172/Y NOR2X1_LOC_536/A 0.04fF
C55300 INVX1_LOC_73/A NAND2X1_LOC_842/B 0.16fF
C55301 NOR2X1_LOC_175/A NOR2X1_LOC_857/A 0.13fF
C55302 NAND2X1_LOC_717/Y INVX1_LOC_76/A 0.03fF
C55303 NOR2X1_LOC_772/Y NOR2X1_LOC_536/A 0.03fF
C55304 NOR2X1_LOC_122/A NOR2X1_LOC_89/A 0.00fF
C55305 INVX1_LOC_102/Y NOR2X1_LOC_153/a_36_216# 0.00fF
C55306 NAND2X1_LOC_505/a_36_24# NOR2X1_LOC_78/A 0.01fF
C55307 NOR2X1_LOC_82/A NAND2X1_LOC_82/Y 0.64fF
C55308 NAND2X1_LOC_151/a_36_24# INVX1_LOC_49/Y 0.00fF
C55309 NAND2X1_LOC_662/Y NOR2X1_LOC_43/Y 0.05fF
C55310 INVX1_LOC_36/A NOR2X1_LOC_697/Y 0.04fF
C55311 NOR2X1_LOC_65/B INVX1_LOC_29/Y 0.05fF
C55312 NOR2X1_LOC_773/Y INVX1_LOC_126/A 0.01fF
C55313 INVX1_LOC_87/Y NOR2X1_LOC_74/A 0.01fF
C55314 VDD NOR2X1_LOC_352/Y 0.29fF
C55315 NOR2X1_LOC_392/B NOR2X1_LOC_536/A 0.01fF
C55316 NOR2X1_LOC_13/Y NOR2X1_LOC_435/A 0.01fF
C55317 INVX1_LOC_191/Y INVX1_LOC_37/A 0.05fF
C55318 NAND2X1_LOC_55/a_36_24# NOR2X1_LOC_271/Y 0.00fF
C55319 NAND2X1_LOC_549/Y INVX1_LOC_23/Y 0.08fF
C55320 NAND2X1_LOC_374/Y VDD 0.26fF
C55321 NOR2X1_LOC_318/B NAND2X1_LOC_656/Y 0.10fF
C55322 NOR2X1_LOC_246/Y NOR2X1_LOC_9/Y 0.10fF
C55323 NOR2X1_LOC_321/Y INVX1_LOC_32/A 0.02fF
C55324 INVX1_LOC_25/Y INVX1_LOC_20/A 0.46fF
C55325 INVX1_LOC_161/Y NOR2X1_LOC_89/A 0.10fF
C55326 NOR2X1_LOC_696/a_36_216# NOR2X1_LOC_696/Y 0.00fF
C55327 NOR2X1_LOC_557/Y NOR2X1_LOC_489/A 0.01fF
C55328 NOR2X1_LOC_134/Y NAND2X1_LOC_74/B 0.03fF
C55329 INVX1_LOC_28/A NOR2X1_LOC_167/Y 0.02fF
C55330 INVX1_LOC_16/A INVX1_LOC_76/A 1.68fF
C55331 NOR2X1_LOC_468/Y INVX1_LOC_15/A 0.03fF
C55332 INVX1_LOC_178/A INVX1_LOC_253/A 0.03fF
C55333 NOR2X1_LOC_773/Y NOR2X1_LOC_111/A 0.04fF
C55334 NOR2X1_LOC_441/Y INVX1_LOC_272/A 0.45fF
C55335 NOR2X1_LOC_78/B INVX1_LOC_117/A 3.19fF
C55336 NOR2X1_LOC_355/B INVX1_LOC_313/Y 0.00fF
C55337 INVX1_LOC_58/A INVX1_LOC_53/A 0.21fF
C55338 INVX1_LOC_23/Y NOR2X1_LOC_291/Y 0.07fF
C55339 NOR2X1_LOC_794/B INVX1_LOC_290/Y 0.32fF
C55340 NAND2X1_LOC_510/A NOR2X1_LOC_509/A 0.05fF
C55341 NOR2X1_LOC_433/A NAND2X1_LOC_288/A 0.17fF
C55342 NAND2X1_LOC_390/A INVX1_LOC_46/A 0.07fF
C55343 NOR2X1_LOC_596/A INVX1_LOC_84/A 0.15fF
C55344 NOR2X1_LOC_173/Y NAND2X1_LOC_175/Y 0.02fF
C55345 NOR2X1_LOC_78/B NOR2X1_LOC_808/B 0.06fF
C55346 INVX1_LOC_141/Y NOR2X1_LOC_669/A 0.01fF
C55347 NOR2X1_LOC_392/B NAND2X1_LOC_93/B 0.10fF
C55348 NOR2X1_LOC_389/A NAND2X1_LOC_220/B 0.39fF
C55349 NOR2X1_LOC_553/B VDD 0.25fF
C55350 INVX1_LOC_30/A INVX1_LOC_12/A 0.95fF
C55351 NOR2X1_LOC_13/Y INVX1_LOC_63/A 0.07fF
C55352 NOR2X1_LOC_510/a_36_216# NOR2X1_LOC_56/Y 0.00fF
C55353 INVX1_LOC_21/A NOR2X1_LOC_843/B 0.00fF
C55354 INVX1_LOC_174/Y NOR2X1_LOC_706/a_36_216# 0.00fF
C55355 INVX1_LOC_143/A NOR2X1_LOC_489/A 0.05fF
C55356 INVX1_LOC_64/A NOR2X1_LOC_392/Y 0.29fF
C55357 INVX1_LOC_144/Y NOR2X1_LOC_506/Y 0.25fF
C55358 NOR2X1_LOC_389/A INVX1_LOC_15/A 0.10fF
C55359 NAND2X1_LOC_833/Y INVX1_LOC_119/Y 0.03fF
C55360 NOR2X1_LOC_763/A INVX1_LOC_296/A 0.77fF
C55361 INVX1_LOC_294/Y INVX1_LOC_285/A 0.02fF
C55362 NOR2X1_LOC_582/A INVX1_LOC_296/A 0.14fF
C55363 INPUT_0 NOR2X1_LOC_557/A 0.05fF
C55364 NOR2X1_LOC_433/A INVX1_LOC_19/A 0.15fF
C55365 INVX1_LOC_14/A NAND2X1_LOC_99/A 0.18fF
C55366 NOR2X1_LOC_392/B INVX1_LOC_3/A 0.01fF
C55367 INVX1_LOC_83/A INVX1_LOC_117/A 0.25fF
C55368 INVX1_LOC_224/A INVX1_LOC_26/Y 0.03fF
C55369 INVX1_LOC_5/A INVX1_LOC_138/Y 0.02fF
C55370 NAND2X1_LOC_726/Y INVX1_LOC_185/A 0.01fF
C55371 INVX1_LOC_28/A INVX1_LOC_76/A 0.32fF
C55372 NAND2X1_LOC_114/B INVX1_LOC_87/A 0.60fF
C55373 INVX1_LOC_299/A NOR2X1_LOC_383/B 0.03fF
C55374 INVX1_LOC_17/A NOR2X1_LOC_693/Y 0.07fF
C55375 INVX1_LOC_34/A NAND2X1_LOC_625/a_36_24# 0.00fF
C55376 INVX1_LOC_285/Y INVX1_LOC_91/A 0.10fF
C55377 NOR2X1_LOC_593/Y INVX1_LOC_19/A 0.61fF
C55378 INVX1_LOC_11/A INVX1_LOC_26/Y 0.06fF
C55379 NOR2X1_LOC_437/Y NOR2X1_LOC_89/A 0.15fF
C55380 NOR2X1_LOC_52/B NOR2X1_LOC_653/Y 0.05fF
C55381 INVX1_LOC_223/Y INVX1_LOC_64/A 0.03fF
C55382 NOR2X1_LOC_605/B INVX1_LOC_185/A 0.00fF
C55383 NAND2X1_LOC_10/a_36_24# INVX1_LOC_27/A 0.00fF
C55384 INPUT_0 NOR2X1_LOC_657/B 0.04fF
C55385 NAND2X1_LOC_773/Y D_INPUT_1 0.00fF
C55386 NAND2X1_LOC_807/Y INVX1_LOC_37/A 0.07fF
C55387 NOR2X1_LOC_6/B NOR2X1_LOC_721/B 0.02fF
C55388 INVX1_LOC_75/A INVX1_LOC_20/A 0.03fF
C55389 INVX1_LOC_100/A INVX1_LOC_304/A 0.42fF
C55390 NOR2X1_LOC_647/A INPUT_3 0.02fF
C55391 NOR2X1_LOC_32/B NAND2X1_LOC_725/B 0.07fF
C55392 INVX1_LOC_90/A NOR2X1_LOC_536/A 5.83fF
C55393 NOR2X1_LOC_52/B INVX1_LOC_19/A 0.06fF
C55394 NOR2X1_LOC_703/B INVX1_LOC_4/Y 0.01fF
C55395 INVX1_LOC_278/A NOR2X1_LOC_468/Y 0.29fF
C55396 NOR2X1_LOC_598/B INVX1_LOC_269/A 0.10fF
C55397 NOR2X1_LOC_68/A NAND2X1_LOC_296/a_36_24# 0.00fF
C55398 NOR2X1_LOC_596/A INVX1_LOC_15/A 0.03fF
C55399 NAND2X1_LOC_778/Y INVX1_LOC_93/A 0.10fF
C55400 NOR2X1_LOC_389/B NOR2X1_LOC_536/A 0.07fF
C55401 INVX1_LOC_233/Y NAND2X1_LOC_576/a_36_24# 0.05fF
C55402 INVX1_LOC_63/Y INVX1_LOC_109/Y 0.93fF
C55403 INVX1_LOC_60/A NAND2X1_LOC_74/B 0.02fF
C55404 INVX1_LOC_256/Y INVX1_LOC_63/A 0.10fF
C55405 D_INPUT_1 INVX1_LOC_252/Y 0.01fF
C55406 NAND2X1_LOC_787/A INVX1_LOC_200/A 0.08fF
C55407 INVX1_LOC_77/A NOR2X1_LOC_467/A 0.05fF
C55408 NOR2X1_LOC_6/B NOR2X1_LOC_610/Y 0.03fF
C55409 NOR2X1_LOC_99/B NOR2X1_LOC_99/Y 0.00fF
C55410 INVX1_LOC_269/A NAND2X1_LOC_725/A 0.30fF
C55411 NAND2X1_LOC_213/A INVX1_LOC_5/A 0.02fF
C55412 INVX1_LOC_50/Y NAND2X1_LOC_473/A 0.07fF
C55413 NAND2X1_LOC_141/A NAND2X1_LOC_82/a_36_24# 0.01fF
C55414 NOR2X1_LOC_512/Y INVX1_LOC_94/Y 0.03fF
C55415 INVX1_LOC_24/A NOR2X1_LOC_334/Y 0.07fF
C55416 INVX1_LOC_2/A NAND2X1_LOC_74/B 0.17fF
C55417 NAND2X1_LOC_722/A INVX1_LOC_12/A 0.07fF
C55418 INVX1_LOC_6/A INVX1_LOC_37/A 0.06fF
C55419 INVX1_LOC_60/Y INVX1_LOC_42/A 0.03fF
C55420 NOR2X1_LOC_15/Y INVX1_LOC_93/A 0.08fF
C55421 NOR2X1_LOC_226/A NAND2X1_LOC_74/B 0.07fF
C55422 INVX1_LOC_90/A NAND2X1_LOC_93/B 0.15fF
C55423 NOR2X1_LOC_214/B NOR2X1_LOC_155/A 0.03fF
C55424 INVX1_LOC_235/Y INVX1_LOC_163/A 0.25fF
C55425 NAND2X1_LOC_787/A NAND2X1_LOC_733/Y 0.03fF
C55426 NOR2X1_LOC_389/B NAND2X1_LOC_93/B 0.07fF
C55427 NAND2X1_LOC_35/Y NAND2X1_LOC_550/A 0.02fF
C55428 INVX1_LOC_142/A NOR2X1_LOC_748/A 0.02fF
C55429 NOR2X1_LOC_91/A NAND2X1_LOC_198/B 0.08fF
C55430 INVX1_LOC_90/A NAND2X1_LOC_425/Y 0.02fF
C55431 NOR2X1_LOC_844/A INVX1_LOC_15/A 0.02fF
C55432 NOR2X1_LOC_454/Y INVX1_LOC_1/A 0.36fF
C55433 NAND2X1_LOC_623/B INVX1_LOC_46/A 0.01fF
C55434 NOR2X1_LOC_13/Y NOR2X1_LOC_65/Y 0.06fF
C55435 NAND2X1_LOC_338/B NAND2X1_LOC_456/a_36_24# 0.00fF
C55436 NOR2X1_LOC_323/Y INVX1_LOC_185/A 0.01fF
C55437 NOR2X1_LOC_272/Y NAND2X1_LOC_337/B 0.10fF
C55438 NOR2X1_LOC_165/Y INVX1_LOC_102/A 0.05fF
C55439 INVX1_LOC_24/A NAND2X1_LOC_464/B 0.61fF
C55440 NOR2X1_LOC_567/B NOR2X1_LOC_862/B 0.10fF
C55441 NAND2X1_LOC_41/Y INVX1_LOC_29/A 0.03fF
C55442 INVX1_LOC_90/A NOR2X1_LOC_649/B 0.07fF
C55443 NAND2X1_LOC_787/A INVX1_LOC_217/A 0.06fF
C55444 NAND2X1_LOC_198/B INVX1_LOC_23/A 0.14fF
C55445 NAND2X1_LOC_214/B NAND2X1_LOC_208/B 0.00fF
C55446 NOR2X1_LOC_78/B INVX1_LOC_3/Y 0.36fF
C55447 NOR2X1_LOC_35/Y INVX1_LOC_76/A 0.01fF
C55448 NOR2X1_LOC_561/Y INVX1_LOC_109/A 0.01fF
C55449 INVX1_LOC_50/A NOR2X1_LOC_753/Y 0.03fF
C55450 NOR2X1_LOC_220/A INVX1_LOC_15/A 0.10fF
C55451 INVX1_LOC_20/A NAND2X1_LOC_453/A 0.03fF
C55452 NOR2X1_LOC_564/Y INVX1_LOC_220/A 0.01fF
C55453 NOR2X1_LOC_356/A NOR2X1_LOC_814/A 0.01fF
C55454 INPUT_1 INVX1_LOC_293/Y 0.32fF
C55455 INVX1_LOC_166/A NOR2X1_LOC_474/A 0.04fF
C55456 NOR2X1_LOC_73/a_36_216# NOR2X1_LOC_814/A 0.01fF
C55457 INVX1_LOC_8/A NOR2X1_LOC_39/a_36_216# 0.01fF
C55458 INVX1_LOC_103/A INVX1_LOC_73/Y 0.01fF
C55459 INVX1_LOC_160/A INVX1_LOC_9/A 0.10fF
C55460 NOR2X1_LOC_719/B INVX1_LOC_284/A 0.02fF
C55461 INVX1_LOC_33/A INVX1_LOC_270/Y 0.47fF
C55462 INVX1_LOC_5/A NAND2X1_LOC_364/A 0.09fF
C55463 NOR2X1_LOC_743/a_36_216# INVX1_LOC_270/Y 0.01fF
C55464 INVX1_LOC_34/A INVX1_LOC_271/A 0.09fF
C55465 NOR2X1_LOC_687/Y NOR2X1_LOC_801/B 0.00fF
C55466 NOR2X1_LOC_65/B INVX1_LOC_60/Y 0.03fF
C55467 INVX1_LOC_11/A INVX1_LOC_161/Y 0.08fF
C55468 NAND2X1_LOC_348/A INVX1_LOC_3/A 0.06fF
C55469 INVX1_LOC_310/Y INVX1_LOC_23/A 0.03fF
C55470 INPUT_1 NAND2X1_LOC_74/B 0.26fF
C55471 INVX1_LOC_251/Y INVX1_LOC_26/A 0.15fF
C55472 NAND2X1_LOC_787/A NAND2X1_LOC_787/B 0.21fF
C55473 INVX1_LOC_27/A NOR2X1_LOC_722/Y 0.03fF
C55474 NOR2X1_LOC_74/A INVX1_LOC_265/Y 0.00fF
C55475 INVX1_LOC_21/A INVX1_LOC_18/A 0.20fF
C55476 NOR2X1_LOC_315/Y NOR2X1_LOC_383/B 2.74fF
C55477 INVX1_LOC_46/A INVX1_LOC_117/A 0.03fF
C55478 INVX1_LOC_104/A INVX1_LOC_57/A 0.15fF
C55479 NOR2X1_LOC_74/A NOR2X1_LOC_814/A 0.07fF
C55480 NAND2X1_LOC_577/A INVX1_LOC_14/A 0.06fF
C55481 NOR2X1_LOC_9/Y INVX1_LOC_285/A 0.10fF
C55482 INVX1_LOC_286/Y NAND2X1_LOC_538/Y 1.06fF
C55483 INPUT_1 NOR2X1_LOC_847/B 0.34fF
C55484 INVX1_LOC_137/Y INVX1_LOC_4/Y 0.13fF
C55485 NOR2X1_LOC_331/a_36_216# NOR2X1_LOC_331/B 0.00fF
C55486 INVX1_LOC_50/A INVX1_LOC_133/Y 0.00fF
C55487 NOR2X1_LOC_337/A INVX1_LOC_63/A 0.03fF
C55488 NOR2X1_LOC_78/A NOR2X1_LOC_831/B 0.08fF
C55489 NOR2X1_LOC_538/Y NOR2X1_LOC_748/A 0.15fF
C55490 NOR2X1_LOC_537/Y NOR2X1_LOC_699/a_36_216# 0.00fF
C55491 NOR2X1_LOC_9/Y NOR2X1_LOC_814/A 0.04fF
C55492 INVX1_LOC_300/A NAND2X1_LOC_175/Y 0.04fF
C55493 NOR2X1_LOC_328/Y NOR2X1_LOC_25/Y 0.01fF
C55494 INVX1_LOC_21/A NOR2X1_LOC_713/B 0.18fF
C55495 INVX1_LOC_304/Y NAND2X1_LOC_787/A 0.28fF
C55496 NAND2X1_LOC_231/Y INVX1_LOC_271/A 0.01fF
C55497 INVX1_LOC_311/A INVX1_LOC_186/Y 0.48fF
C55498 INVX1_LOC_200/A INVX1_LOC_30/A 0.85fF
C55499 INVX1_LOC_162/Y NOR2X1_LOC_129/a_36_216# 0.00fF
C55500 NAND2X1_LOC_51/B INVX1_LOC_261/A 0.00fF
C55501 NOR2X1_LOC_721/Y INVX1_LOC_125/A 0.21fF
C55502 INVX1_LOC_64/A NAND2X1_LOC_33/Y 0.54fF
C55503 NOR2X1_LOC_486/a_36_216# NOR2X1_LOC_590/A 0.00fF
C55504 NOR2X1_LOC_155/A NOR2X1_LOC_275/A 0.01fF
C55505 NOR2X1_LOC_88/A NOR2X1_LOC_670/Y 0.16fF
C55506 NOR2X1_LOC_19/B NOR2X1_LOC_128/a_36_216# 0.00fF
C55507 INVX1_LOC_75/A NOR2X1_LOC_128/A 0.06fF
C55508 INVX1_LOC_59/A D_INPUT_2 0.01fF
C55509 NAND2X1_LOC_214/B INVX1_LOC_34/A 0.10fF
C55510 INVX1_LOC_58/A NOR2X1_LOC_78/B 0.24fF
C55511 NOR2X1_LOC_252/Y NOR2X1_LOC_693/Y 0.02fF
C55512 INVX1_LOC_45/A NOR2X1_LOC_254/A 0.07fF
C55513 NOR2X1_LOC_401/a_36_216# INVX1_LOC_23/A 0.02fF
C55514 NOR2X1_LOC_80/a_36_216# NAND2X1_LOC_572/B 0.01fF
C55515 NAND2X1_LOC_849/B NOR2X1_LOC_536/A 0.03fF
C55516 INVX1_LOC_235/Y INVX1_LOC_203/Y 0.07fF
C55517 INVX1_LOC_14/A NAND2X1_LOC_656/A 0.12fF
C55518 NOR2X1_LOC_355/A INVX1_LOC_78/A 0.50fF
C55519 NOR2X1_LOC_15/Y NOR2X1_LOC_303/Y 0.10fF
C55520 NOR2X1_LOC_536/A INVX1_LOC_38/A 0.35fF
C55521 NAND2X1_LOC_565/B NAND2X1_LOC_464/B -0.03fF
C55522 NAND2X1_LOC_364/A NAND2X1_LOC_337/B 0.31fF
C55523 INVX1_LOC_34/A INVX1_LOC_27/A 0.17fF
C55524 NOR2X1_LOC_219/Y INVX1_LOC_23/A 0.72fF
C55525 NOR2X1_LOC_637/B NOR2X1_LOC_92/Y 0.00fF
C55526 INVX1_LOC_17/A INVX1_LOC_45/Y 0.03fF
C55527 NAND2X1_LOC_785/A NAND2X1_LOC_552/A 0.09fF
C55528 NAND2X1_LOC_9/Y NAND2X1_LOC_181/Y 0.06fF
C55529 INVX1_LOC_1/A INVX1_LOC_77/A 0.70fF
C55530 INVX1_LOC_34/A NOR2X1_LOC_824/A 0.07fF
C55531 INVX1_LOC_136/A NOR2X1_LOC_134/Y 0.00fF
C55532 NAND2X1_LOC_687/A INVX1_LOC_291/A 0.01fF
C55533 INVX1_LOC_53/Y INVX1_LOC_23/A 4.40fF
C55534 INVX1_LOC_233/A NAND2X1_LOC_181/Y 0.01fF
C55535 INPUT_0 INVX1_LOC_170/Y 0.02fF
C55536 INVX1_LOC_36/A NOR2X1_LOC_426/Y 0.01fF
C55537 NAND2X1_LOC_796/B NAND2X1_LOC_357/B -0.01fF
C55538 NAND2X1_LOC_692/a_36_24# INVX1_LOC_275/Y 0.00fF
C55539 NOR2X1_LOC_447/B NOR2X1_LOC_88/Y 0.02fF
C55540 INVX1_LOC_124/Y NOR2X1_LOC_266/a_36_216# -0.00fF
C55541 NOR2X1_LOC_92/Y NAND2X1_LOC_569/A 0.00fF
C55542 NOR2X1_LOC_665/A INVX1_LOC_23/A 0.14fF
C55543 NOR2X1_LOC_813/Y NOR2X1_LOC_235/Y 0.03fF
C55544 NAND2X1_LOC_30/Y NAND2X1_LOC_17/a_36_24# 0.00fF
C55545 NOR2X1_LOC_91/A NAND2X1_LOC_728/a_36_24# 0.01fF
C55546 NOR2X1_LOC_65/B NOR2X1_LOC_355/A 0.01fF
C55547 INVX1_LOC_1/Y NOR2X1_LOC_717/A 0.01fF
C55548 NOR2X1_LOC_6/B NAND2X1_LOC_473/A 0.02fF
C55549 INVX1_LOC_75/A INVX1_LOC_4/A 0.49fF
C55550 NAND2X1_LOC_569/a_36_24# NOR2X1_LOC_384/Y 0.00fF
C55551 NAND2X1_LOC_785/A INVX1_LOC_178/A 0.10fF
C55552 INVX1_LOC_258/A INVX1_LOC_207/A 0.06fF
C55553 NAND2X1_LOC_860/A INVX1_LOC_30/Y 0.95fF
C55554 INVX1_LOC_64/A INVX1_LOC_25/Y 0.05fF
C55555 NAND2X1_LOC_190/a_36_24# NOR2X1_LOC_78/B 0.00fF
C55556 D_INPUT_1 INVX1_LOC_279/A 0.08fF
C55557 NOR2X1_LOC_286/Y NAND2X1_LOC_361/Y 0.00fF
C55558 NOR2X1_LOC_433/A INVX1_LOC_161/Y 0.13fF
C55559 INVX1_LOC_217/A INVX1_LOC_30/A 0.09fF
C55560 NAND2X1_LOC_846/a_36_24# INVX1_LOC_291/A 0.01fF
C55561 NOR2X1_LOC_216/Y NOR2X1_LOC_334/Y 0.07fF
C55562 INVX1_LOC_38/A NAND2X1_LOC_93/B 0.85fF
C55563 INVX1_LOC_145/Y INVX1_LOC_23/A 0.00fF
C55564 NOR2X1_LOC_500/A NAND2X1_LOC_321/a_36_24# 0.00fF
C55565 INVX1_LOC_59/A NOR2X1_LOC_529/Y -0.10fF
C55566 NOR2X1_LOC_178/Y INVX1_LOC_16/A 0.15fF
C55567 INVX1_LOC_58/A INVX1_LOC_83/A 0.05fF
C55568 D_INPUT_0 NOR2X1_LOC_414/Y 0.77fF
C55569 NOR2X1_LOC_226/A NAND2X1_LOC_793/a_36_24# 0.00fF
C55570 NOR2X1_LOC_272/Y NOR2X1_LOC_773/Y 0.10fF
C55571 INVX1_LOC_124/A INVX1_LOC_1/A 0.41fF
C55572 INVX1_LOC_38/A NAND2X1_LOC_425/Y 0.07fF
C55573 NOR2X1_LOC_82/Y INVX1_LOC_306/Y 0.03fF
C55574 INVX1_LOC_89/A INVX1_LOC_129/A 0.05fF
C55575 INVX1_LOC_150/Y NOR2X1_LOC_142/Y 0.30fF
C55576 NOR2X1_LOC_71/Y NAND2X1_LOC_203/a_36_24# 0.00fF
C55577 NOR2X1_LOC_15/Y INVX1_LOC_54/Y 0.05fF
C55578 NOR2X1_LOC_285/a_36_216# INVX1_LOC_89/A 0.00fF
C55579 NOR2X1_LOC_40/a_36_216# NOR2X1_LOC_11/Y 0.00fF
C55580 INVX1_LOC_123/A NOR2X1_LOC_38/B 0.07fF
C55581 NOR2X1_LOC_598/B NOR2X1_LOC_814/Y 0.02fF
C55582 INVX1_LOC_109/A INVX1_LOC_76/A 0.14fF
C55583 INVX1_LOC_131/Y NOR2X1_LOC_743/Y 0.31fF
C55584 INVX1_LOC_161/Y NOR2X1_LOC_52/B 0.17fF
C55585 NOR2X1_LOC_433/A NOR2X1_LOC_599/A 0.18fF
C55586 NOR2X1_LOC_637/Y NAND2X1_LOC_354/Y 0.15fF
C55587 NOR2X1_LOC_68/Y INVX1_LOC_117/A 0.16fF
C55588 INVX1_LOC_258/Y INVX1_LOC_22/A 0.23fF
C55589 NOR2X1_LOC_742/A NOR2X1_LOC_727/B 0.48fF
C55590 INVX1_LOC_30/A NAND2X1_LOC_787/B 0.17fF
C55591 NAND2X1_LOC_500/Y NAND2X1_LOC_483/Y 0.01fF
C55592 INVX1_LOC_9/Y NOR2X1_LOC_321/Y 0.26fF
C55593 NOR2X1_LOC_92/Y INVX1_LOC_316/Y 0.02fF
C55594 INVX1_LOC_136/A INVX1_LOC_49/A 0.05fF
C55595 INPUT_1 NOR2X1_LOC_660/Y 0.07fF
C55596 INVX1_LOC_91/A INVX1_LOC_4/Y 0.20fF
C55597 NOR2X1_LOC_68/A NAND2X1_LOC_7/Y 0.05fF
C55598 INVX1_LOC_48/Y NOR2X1_LOC_719/A 0.01fF
C55599 D_INPUT_1 INVX1_LOC_182/Y 0.04fF
C55600 INVX1_LOC_1/A NOR2X1_LOC_687/Y 0.07fF
C55601 NAND2X1_LOC_655/B INVX1_LOC_15/A 0.07fF
C55602 NOR2X1_LOC_778/B INVX1_LOC_225/Y 0.03fF
C55603 NOR2X1_LOC_78/B INVX1_LOC_215/Y 0.06fF
C55604 NAND2X1_LOC_469/B INVX1_LOC_15/A 0.01fF
C55605 INPUT_0 INVX1_LOC_271/A 0.78fF
C55606 NAND2X1_LOC_733/Y NAND2X1_LOC_722/A 0.10fF
C55607 NOR2X1_LOC_226/A INVX1_LOC_211/A 0.23fF
C55608 NOR2X1_LOC_111/A INVX1_LOC_42/A 0.12fF
C55609 INVX1_LOC_209/Y INVX1_LOC_24/A 0.03fF
C55610 INVX1_LOC_304/Y INVX1_LOC_30/A 0.07fF
C55611 NAND2X1_LOC_116/A INVX1_LOC_110/A 0.00fF
C55612 NOR2X1_LOC_322/Y NAND2X1_LOC_793/B 0.10fF
C55613 INVX1_LOC_85/Y INVX1_LOC_50/Y 0.00fF
C55614 NOR2X1_LOC_437/Y NOR2X1_LOC_433/A 0.08fF
C55615 INVX1_LOC_57/Y NOR2X1_LOC_315/Y 0.20fF
C55616 NOR2X1_LOC_67/A INVX1_LOC_61/Y 0.07fF
C55617 NOR2X1_LOC_640/Y INVX1_LOC_63/A 0.07fF
C55618 NAND2X1_LOC_475/Y INVX1_LOC_92/A 0.03fF
C55619 NAND2X1_LOC_564/B NAND2X1_LOC_793/Y 0.12fF
C55620 INVX1_LOC_64/A INVX1_LOC_75/A 0.25fF
C55621 NAND2X1_LOC_508/A NOR2X1_LOC_849/A 0.04fF
C55622 NOR2X1_LOC_82/A NOR2X1_LOC_789/A 0.00fF
C55623 INVX1_LOC_43/Y INVX1_LOC_25/Y 0.92fF
C55624 INVX1_LOC_211/Y NOR2X1_LOC_328/Y 0.04fF
C55625 INVX1_LOC_13/Y NOR2X1_LOC_756/Y 0.02fF
C55626 INVX1_LOC_118/A NAND2X1_LOC_74/B 0.15fF
C55627 INVX1_LOC_174/A INVX1_LOC_22/A 0.35fF
C55628 NAND2X1_LOC_206/B INVX1_LOC_230/A 0.75fF
C55629 NOR2X1_LOC_218/Y NOR2X1_LOC_276/Y 0.03fF
C55630 NAND2X1_LOC_736/Y NAND2X1_LOC_863/Y 0.09fF
C55631 NOR2X1_LOC_443/Y INVX1_LOC_186/A 0.01fF
C55632 INVX1_LOC_249/A INVX1_LOC_34/A 0.05fF
C55633 INVX1_LOC_2/A INVX1_LOC_136/A 0.20fF
C55634 NOR2X1_LOC_160/B NOR2X1_LOC_507/A 0.13fF
C55635 INVX1_LOC_24/A NOR2X1_LOC_718/B 1.33fF
C55636 NAND2X1_LOC_722/A INVX1_LOC_217/A 0.07fF
C55637 INVX1_LOC_41/A INVX1_LOC_8/Y 0.01fF
C55638 INVX1_LOC_73/A NOR2X1_LOC_674/Y 0.07fF
C55639 INVX1_LOC_136/A NOR2X1_LOC_226/A 0.14fF
C55640 NOR2X1_LOC_243/B NOR2X1_LOC_814/A 0.07fF
C55641 INVX1_LOC_255/Y NAND2X1_LOC_555/Y 0.02fF
C55642 NAND2X1_LOC_85/Y INVX1_LOC_63/A 0.11fF
C55643 INVX1_LOC_214/A INVX1_LOC_18/A 0.03fF
C55644 INVX1_LOC_238/Y GATE_865 0.06fF
C55645 NAND2X1_LOC_564/A NOR2X1_LOC_45/B 0.03fF
C55646 NOR2X1_LOC_859/a_36_216# INVX1_LOC_135/A 0.00fF
C55647 NOR2X1_LOC_667/A INVX1_LOC_18/A 0.07fF
C55648 INVX1_LOC_27/A INVX1_LOC_131/A 0.69fF
C55649 INVX1_LOC_246/A NOR2X1_LOC_561/Y 0.02fF
C55650 NOR2X1_LOC_738/Y INVX1_LOC_83/A 0.01fF
C55651 INVX1_LOC_17/A NOR2X1_LOC_71/Y 0.79fF
C55652 INVX1_LOC_232/Y NOR2X1_LOC_68/A 0.01fF
C55653 INVX1_LOC_289/A INVX1_LOC_36/A 0.03fF
C55654 NOR2X1_LOC_191/B NOR2X1_LOC_709/A 0.01fF
C55655 INVX1_LOC_170/A INVX1_LOC_56/Y 0.39fF
C55656 INVX1_LOC_233/Y INVX1_LOC_309/A 0.03fF
C55657 NAND2X1_LOC_214/B INPUT_0 0.07fF
C55658 INVX1_LOC_248/A INVX1_LOC_18/A 0.07fF
C55659 INVX1_LOC_119/A NAND2X1_LOC_593/Y 0.03fF
C55660 INVX1_LOC_64/A NOR2X1_LOC_7/a_36_216# 0.01fF
C55661 INVX1_LOC_111/Y NAND2X1_LOC_656/A 0.01fF
C55662 NOR2X1_LOC_92/Y NAND2X1_LOC_850/A 0.06fF
C55663 INVX1_LOC_215/Y INVX1_LOC_83/A 0.10fF
C55664 NOR2X1_LOC_111/A INVX1_LOC_78/A 0.07fF
C55665 NOR2X1_LOC_303/Y INVX1_LOC_96/Y 0.10fF
C55666 NOR2X1_LOC_287/A INVX1_LOC_305/A 0.04fF
C55667 INVX1_LOC_41/A NOR2X1_LOC_264/Y 0.21fF
C55668 NOR2X1_LOC_318/B NOR2X1_LOC_717/A 0.10fF
C55669 NOR2X1_LOC_790/B NOR2X1_LOC_78/A 0.07fF
C55670 NOR2X1_LOC_220/A NOR2X1_LOC_168/Y 0.03fF
C55671 INVX1_LOC_21/A NOR2X1_LOC_185/a_36_216# 0.02fF
C55672 INVX1_LOC_230/Y INVX1_LOC_135/A 0.29fF
C55673 INVX1_LOC_34/A NOR2X1_LOC_664/Y 0.16fF
C55674 NAND2X1_LOC_711/B NOR2X1_LOC_667/A 0.02fF
C55675 INVX1_LOC_27/A INPUT_0 0.29fF
C55676 INVX1_LOC_233/Y INVX1_LOC_91/A 0.01fF
C55677 INVX1_LOC_12/A INVX1_LOC_113/A 0.23fF
C55678 INVX1_LOC_256/A INVX1_LOC_90/A 0.13fF
C55679 INVX1_LOC_21/A NOR2X1_LOC_548/A 0.01fF
C55680 INVX1_LOC_24/A INVX1_LOC_218/A 0.04fF
C55681 NOR2X1_LOC_419/Y NOR2X1_LOC_520/A 0.00fF
C55682 NOR2X1_LOC_75/Y D_GATE_366 0.03fF
C55683 NOR2X1_LOC_781/A INVX1_LOC_72/A 0.02fF
C55684 INVX1_LOC_93/Y NOR2X1_LOC_717/A 0.10fF
C55685 NAND2X1_LOC_860/A NOR2X1_LOC_124/A 0.04fF
C55686 NOR2X1_LOC_536/A NAND2X1_LOC_223/A 0.03fF
C55687 INVX1_LOC_256/A NOR2X1_LOC_389/B 0.07fF
C55688 NOR2X1_LOC_6/B NOR2X1_LOC_516/Y 0.02fF
C55689 NAND2X1_LOC_465/A INVX1_LOC_23/A 0.02fF
C55690 INVX1_LOC_208/A INVX1_LOC_94/A 0.01fF
C55691 NOR2X1_LOC_210/A NOR2X1_LOC_68/A 0.01fF
C55692 NOR2X1_LOC_667/A INVX1_LOC_172/A 0.01fF
C55693 NOR2X1_LOC_521/Y INVX1_LOC_18/A 0.01fF
C55694 NOR2X1_LOC_808/A NOR2X1_LOC_804/B 0.03fF
C55695 NOR2X1_LOC_65/B NOR2X1_LOC_111/A 0.07fF
C55696 NAND2X1_LOC_768/Y NAND2X1_LOC_772/a_36_24# 0.00fF
C55697 NAND2X1_LOC_141/A NOR2X1_LOC_84/A 0.00fF
C55698 NOR2X1_LOC_168/Y NOR2X1_LOC_548/Y 0.34fF
C55699 INVX1_LOC_233/Y INVX1_LOC_11/Y 0.07fF
C55700 INVX1_LOC_1/A NAND2X1_LOC_832/Y 0.01fF
C55701 INVX1_LOC_32/A NAND2X1_LOC_798/B 0.07fF
C55702 INVX1_LOC_58/A INVX1_LOC_46/A 0.73fF
C55703 INVX1_LOC_24/A NOR2X1_LOC_569/Y 0.07fF
C55704 NOR2X1_LOC_590/A NOR2X1_LOC_356/A 0.10fF
C55705 INVX1_LOC_17/A NOR2X1_LOC_751/A 0.06fF
C55706 NAND2X1_LOC_514/Y NAND2X1_LOC_656/Y 0.03fF
C55707 INVX1_LOC_45/A NOR2X1_LOC_473/B 0.01fF
C55708 INVX1_LOC_171/A NOR2X1_LOC_274/B 0.01fF
C55709 INVX1_LOC_23/A INVX1_LOC_77/Y 0.07fF
C55710 NOR2X1_LOC_68/A NOR2X1_LOC_312/Y 0.17fF
C55711 INVX1_LOC_43/Y INVX1_LOC_75/A 0.03fF
C55712 INVX1_LOC_136/A NAND2X1_LOC_648/A 0.03fF
C55713 NOR2X1_LOC_226/A NOR2X1_LOC_278/A 0.03fF
C55714 INVX1_LOC_172/A NOR2X1_LOC_521/Y 0.07fF
C55715 NOR2X1_LOC_589/A NOR2X1_LOC_577/Y 0.03fF
C55716 NAND2X1_LOC_63/Y NAND2X1_LOC_74/B 0.10fF
C55717 INVX1_LOC_136/A INPUT_1 1.18fF
C55718 INVX1_LOC_64/A NAND2X1_LOC_453/A 0.07fF
C55719 NOR2X1_LOC_334/Y NOR2X1_LOC_197/B 0.10fF
C55720 NOR2X1_LOC_433/a_36_216# INVX1_LOC_22/A 0.00fF
C55721 NAND2X1_LOC_569/B VDD 0.14fF
C55722 NAND2X1_LOC_254/Y INVX1_LOC_19/A 0.08fF
C55723 INVX1_LOC_5/A NOR2X1_LOC_857/A 0.07fF
C55724 NOR2X1_LOC_34/B NOR2X1_LOC_35/Y 0.02fF
C55725 INVX1_LOC_37/A NOR2X1_LOC_109/Y 0.07fF
C55726 NOR2X1_LOC_590/A NOR2X1_LOC_74/A 0.10fF
C55727 D_INPUT_0 NOR2X1_LOC_237/a_36_216# 0.01fF
C55728 NOR2X1_LOC_167/a_36_216# INVX1_LOC_92/A 0.01fF
C55729 INVX1_LOC_230/Y NOR2X1_LOC_391/B 0.01fF
C55730 INVX1_LOC_90/A NOR2X1_LOC_781/Y 0.02fF
C55731 NAND2X1_LOC_455/B NAND2X1_LOC_74/B 0.01fF
C55732 NOR2X1_LOC_617/Y INVX1_LOC_89/A 0.21fF
C55733 NOR2X1_LOC_297/A NAND2X1_LOC_206/Y 0.06fF
C55734 INVX1_LOC_25/A INVX1_LOC_9/A 0.65fF
C55735 VDD NOR2X1_LOC_81/Y 0.12fF
C55736 NOR2X1_LOC_391/A INVX1_LOC_8/A 0.07fF
C55737 INVX1_LOC_73/A INVX1_LOC_72/A 0.03fF
C55738 NOR2X1_LOC_473/B INVX1_LOC_71/A 0.23fF
C55739 NOR2X1_LOC_440/Y NOR2X1_LOC_392/B 0.27fF
C55740 INVX1_LOC_34/A INVX1_LOC_234/A 0.14fF
C55741 NAND2X1_LOC_562/B NAND2X1_LOC_632/a_36_24# 0.01fF
C55742 NAND2X1_LOC_736/Y NOR2X1_LOC_700/a_36_216# 0.01fF
C55743 NOR2X1_LOC_393/Y NAND2X1_LOC_773/B 0.02fF
C55744 NAND2X1_LOC_361/Y INVX1_LOC_148/Y 0.01fF
C55745 INVX1_LOC_48/Y INVX1_LOC_76/A 0.08fF
C55746 NOR2X1_LOC_860/B NOR2X1_LOC_112/Y 0.04fF
C55747 NAND2X1_LOC_51/B INVX1_LOC_18/A 2.94fF
C55748 INVX1_LOC_25/Y NAND2X1_LOC_850/Y 0.07fF
C55749 NOR2X1_LOC_553/B INVX1_LOC_177/A 0.02fF
C55750 NOR2X1_LOC_785/A NOR2X1_LOC_78/A 0.00fF
C55751 INVX1_LOC_222/A NOR2X1_LOC_274/B 0.50fF
C55752 NOR2X1_LOC_671/Y INVX1_LOC_3/Y 0.04fF
C55753 NAND2X1_LOC_337/B NOR2X1_LOC_405/A 0.26fF
C55754 NOR2X1_LOC_798/A INVX1_LOC_117/A 0.03fF
C55755 NAND2X1_LOC_704/a_36_24# NAND2X1_LOC_453/A 0.00fF
C55756 INVX1_LOC_180/A NAND2X1_LOC_652/Y 0.26fF
C55757 INVX1_LOC_141/A NOR2X1_LOC_45/B 0.08fF
C55758 NOR2X1_LOC_736/Y INVX1_LOC_113/Y 0.03fF
C55759 NOR2X1_LOC_140/A VDD 0.10fF
C55760 INVX1_LOC_311/A INVX1_LOC_18/A 0.33fF
C55761 NOR2X1_LOC_218/A NAND2X1_LOC_468/B 0.03fF
C55762 NOR2X1_LOC_131/Y INVX1_LOC_22/A 0.01fF
C55763 INVX1_LOC_45/A NOR2X1_LOC_355/B 0.08fF
C55764 NOR2X1_LOC_418/Y INVX1_LOC_22/A 0.02fF
C55765 INVX1_LOC_81/Y NOR2X1_LOC_78/A 0.04fF
C55766 NOR2X1_LOC_298/Y NOR2X1_LOC_822/Y 0.11fF
C55767 NOR2X1_LOC_68/A NOR2X1_LOC_391/Y 0.02fF
C55768 NAND2X1_LOC_722/A NAND2X1_LOC_808/A 0.02fF
C55769 INVX1_LOC_41/A NAND2X1_LOC_850/A 0.04fF
C55770 NAND2X1_LOC_538/Y VDD 0.81fF
C55771 NAND2X1_LOC_198/B INVX1_LOC_6/A 0.01fF
C55772 NAND2X1_LOC_88/a_36_24# INVX1_LOC_62/A 0.00fF
C55773 NOR2X1_LOC_743/Y NOR2X1_LOC_109/Y 0.07fF
C55774 INVX1_LOC_34/A NOR2X1_LOC_19/B 0.22fF
C55775 NOR2X1_LOC_577/a_36_216# NOR2X1_LOC_500/Y 0.01fF
C55776 NOR2X1_LOC_788/B NOR2X1_LOC_802/A 0.01fF
C55777 INVX1_LOC_283/A INVX1_LOC_4/A 0.01fF
C55778 NAND2X1_LOC_152/a_36_24# NOR2X1_LOC_499/B 0.00fF
C55779 NOR2X1_LOC_589/A INVX1_LOC_22/A 0.32fF
C55780 INVX1_LOC_89/A NOR2X1_LOC_538/Y 0.01fF
C55781 INVX1_LOC_39/Y INVX1_LOC_59/Y 0.11fF
C55782 INVX1_LOC_77/A NOR2X1_LOC_188/A 0.04fF
C55783 NAND2X1_LOC_656/A INVX1_LOC_48/A 0.10fF
C55784 NAND2X1_LOC_479/Y GATE_479 0.03fF
C55785 INVX1_LOC_77/A NOR2X1_LOC_548/B 0.03fF
C55786 INVX1_LOC_215/Y INVX1_LOC_46/A 0.04fF
C55787 NOR2X1_LOC_531/a_36_216# INVX1_LOC_91/A 0.00fF
C55788 INVX1_LOC_72/A NAND2X1_LOC_729/B 0.03fF
C55789 NOR2X1_LOC_530/Y VDD 0.18fF
C55790 NOR2X1_LOC_226/A NAND2X1_LOC_862/Y 0.07fF
C55791 INVX1_LOC_229/Y INVX1_LOC_22/A 0.36fF
C55792 INVX1_LOC_290/A NOR2X1_LOC_561/Y 0.10fF
C55793 NAND2X1_LOC_736/Y INVX1_LOC_282/A 0.00fF
C55794 INVX1_LOC_53/A NAND2X1_LOC_475/Y 0.10fF
C55795 NOR2X1_LOC_409/B NOR2X1_LOC_48/B 0.02fF
C55796 NOR2X1_LOC_355/B INVX1_LOC_71/A 0.00fF
C55797 NAND2X1_LOC_785/A INVX1_LOC_140/A 0.25fF
C55798 INVX1_LOC_1/A INVX1_LOC_9/A 0.31fF
C55799 INVX1_LOC_314/Y INVX1_LOC_125/Y 0.04fF
C55800 NOR2X1_LOC_384/Y NOR2X1_LOC_670/a_36_216# 0.00fF
C55801 NOR2X1_LOC_186/Y NOR2X1_LOC_831/B 1.00fF
C55802 INVX1_LOC_171/A INVX1_LOC_22/A 0.10fF
C55803 INVX1_LOC_313/A INVX1_LOC_53/Y 0.13fF
C55804 NOR2X1_LOC_859/a_36_216# INVX1_LOC_280/A 0.01fF
C55805 NOR2X1_LOC_658/Y INVX1_LOC_139/A 0.02fF
C55806 D_INPUT_7 NAND2X1_LOC_1/Y 0.03fF
C55807 INVX1_LOC_18/A NOR2X1_LOC_670/Y 0.03fF
C55808 INVX1_LOC_256/A INVX1_LOC_38/A 0.09fF
C55809 NAND2X1_LOC_11/Y INVX1_LOC_140/A 0.13fF
C55810 NOR2X1_LOC_392/B INVX1_LOC_69/Y 0.03fF
C55811 INVX1_LOC_295/A GATE_479 0.07fF
C55812 NOR2X1_LOC_273/Y NAND2X1_LOC_212/Y 0.05fF
C55813 INVX1_LOC_136/A NOR2X1_LOC_586/Y 0.00fF
C55814 INVX1_LOC_36/A INVX1_LOC_37/A 0.10fF
C55815 NOR2X1_LOC_113/a_36_216# NOR2X1_LOC_114/Y 0.00fF
C55816 INVX1_LOC_58/A NOR2X1_LOC_671/Y 0.18fF
C55817 INVX1_LOC_124/A NOR2X1_LOC_188/A 0.08fF
C55818 INVX1_LOC_83/A NOR2X1_LOC_777/a_36_216# 0.02fF
C55819 NAND2X1_LOC_170/A NOR2X1_LOC_166/Y 0.01fF
C55820 NAND2X1_LOC_573/Y NOR2X1_LOC_831/B 0.23fF
C55821 NOR2X1_LOC_15/Y NAND2X1_LOC_656/B 0.01fF
C55822 INVX1_LOC_230/Y INVX1_LOC_280/A 4.52fF
C55823 NOR2X1_LOC_794/B INVX1_LOC_9/A 0.03fF
C55824 INVX1_LOC_230/Y NOR2X1_LOC_94/Y 0.03fF
C55825 NOR2X1_LOC_208/Y NOR2X1_LOC_631/B 0.01fF
C55826 INVX1_LOC_34/A NOR2X1_LOC_528/Y 0.34fF
C55827 INVX1_LOC_145/Y INVX1_LOC_313/A 0.02fF
C55828 INVX1_LOC_17/A NAND2X1_LOC_243/Y 0.00fF
C55829 NAND2X1_LOC_662/B NAND2X1_LOC_661/B 0.19fF
C55830 NOR2X1_LOC_15/Y INVX1_LOC_35/Y 0.38fF
C55831 NOR2X1_LOC_716/B NOR2X1_LOC_80/a_36_216# 0.01fF
C55832 INVX1_LOC_135/A NOR2X1_LOC_415/a_36_216# 0.00fF
C55833 NOR2X1_LOC_440/Y NOR2X1_LOC_389/B 0.42fF
C55834 NOR2X1_LOC_620/Y NOR2X1_LOC_545/B 0.01fF
C55835 NAND2X1_LOC_200/B INPUT_0 0.01fF
C55836 INVX1_LOC_39/A INVX1_LOC_293/Y 0.26fF
C55837 NOR2X1_LOC_112/Y NOR2X1_LOC_97/B 0.05fF
C55838 INVX1_LOC_64/A NAND2X1_LOC_291/B 0.03fF
C55839 NOR2X1_LOC_189/A INVX1_LOC_76/A 0.03fF
C55840 NOR2X1_LOC_626/Y INVX1_LOC_186/Y 0.01fF
C55841 NOR2X1_LOC_577/Y INVX1_LOC_20/A 0.08fF
C55842 NOR2X1_LOC_274/a_36_216# INVX1_LOC_14/Y 0.00fF
C55843 NAND2X1_LOC_796/a_36_24# INVX1_LOC_54/A 0.01fF
C55844 NAND2X1_LOC_711/Y INVX1_LOC_185/A 0.02fF
C55845 INVX1_LOC_24/A NAND2X1_LOC_472/Y 0.07fF
C55846 NOR2X1_LOC_532/Y NOR2X1_LOC_788/B 0.12fF
C55847 INVX1_LOC_222/A INVX1_LOC_22/A 0.03fF
C55848 INPUT_0 INVX1_LOC_137/A 0.00fF
C55849 NOR2X1_LOC_160/B NOR2X1_LOC_155/A 0.13fF
C55850 NOR2X1_LOC_237/Y INVX1_LOC_37/A 0.03fF
C55851 NOR2X1_LOC_92/Y NOR2X1_LOC_662/A 0.07fF
C55852 INVX1_LOC_5/A INVX1_LOC_109/Y 0.01fF
C55853 NOR2X1_LOC_590/A NOR2X1_LOC_650/a_36_216# 0.00fF
C55854 NAND2X1_LOC_9/Y INVX1_LOC_3/Y 0.05fF
C55855 NOR2X1_LOC_219/Y INVX1_LOC_6/A 0.16fF
C55856 INVX1_LOC_39/A NAND2X1_LOC_74/B -0.01fF
C55857 INVX1_LOC_11/A NAND2X1_LOC_426/a_36_24# -0.02fF
C55858 NOR2X1_LOC_152/Y NOR2X1_LOC_111/A 0.01fF
C55859 NOR2X1_LOC_335/B NOR2X1_LOC_188/a_36_216# 0.01fF
C55860 NOR2X1_LOC_82/Y NOR2X1_LOC_9/Y 0.14fF
C55861 D_INPUT_1 NOR2X1_LOC_38/B 0.13fF
C55862 NOR2X1_LOC_180/B INVX1_LOC_313/Y 0.07fF
C55863 NOR2X1_LOC_139/Y NOR2X1_LOC_131/A 0.05fF
C55864 INVX1_LOC_53/Y INVX1_LOC_6/A 0.11fF
C55865 INVX1_LOC_136/A INVX1_LOC_118/A 0.29fF
C55866 NOR2X1_LOC_526/Y INVX1_LOC_91/A 0.01fF
C55867 NOR2X1_LOC_589/A INVX1_LOC_100/A 0.04fF
C55868 INVX1_LOC_227/A NOR2X1_LOC_74/A 0.31fF
C55869 INVX1_LOC_234/A INPUT_0 0.07fF
C55870 INVX1_LOC_30/A INVX1_LOC_92/A 1.52fF
C55871 INVX1_LOC_57/A NOR2X1_LOC_281/a_36_216# 0.00fF
C55872 NOR2X1_LOC_548/a_36_216# NOR2X1_LOC_548/Y 0.00fF
C55873 NOR2X1_LOC_590/A NOR2X1_LOC_243/B 0.01fF
C55874 NOR2X1_LOC_272/Y INVX1_LOC_42/A 0.39fF
C55875 NOR2X1_LOC_370/a_36_216# NOR2X1_LOC_335/B 0.00fF
C55876 NOR2X1_LOC_660/Y NAND2X1_LOC_618/Y 0.09fF
C55877 NAND2X1_LOC_763/B INVX1_LOC_92/A 0.11fF
C55878 NOR2X1_LOC_131/A NAND2X1_LOC_468/B -0.00fF
C55879 NOR2X1_LOC_356/A NOR2X1_LOC_703/A 0.09fF
C55880 NOR2X1_LOC_383/B NAND2X1_LOC_99/A 0.01fF
C55881 NOR2X1_LOC_84/Y INVX1_LOC_76/A 0.19fF
C55882 INVX1_LOC_73/A INVX1_LOC_313/Y 0.23fF
C55883 NOR2X1_LOC_309/Y INVX1_LOC_37/A 0.46fF
C55884 NOR2X1_LOC_191/A INVX1_LOC_95/Y 0.00fF
C55885 INVX1_LOC_271/Y NOR2X1_LOC_678/A 0.62fF
C55886 INVX1_LOC_269/A INVX1_LOC_29/A 0.32fF
C55887 INVX1_LOC_87/A NOR2X1_LOC_717/A 0.08fF
C55888 INVX1_LOC_33/A NOR2X1_LOC_536/A 0.09fF
C55889 INVX1_LOC_135/A NOR2X1_LOC_391/a_36_216# 0.01fF
C55890 VDD NOR2X1_LOC_709/A 2.01fF
C55891 INVX1_LOC_259/Y NOR2X1_LOC_631/Y 0.01fF
C55892 INVX1_LOC_50/A NAND2X1_LOC_787/Y 0.09fF
C55893 NOR2X1_LOC_346/B NOR2X1_LOC_360/A 0.01fF
C55894 NOR2X1_LOC_13/Y INVX1_LOC_117/Y 0.00fF
C55895 INVX1_LOC_69/Y NOR2X1_LOC_355/a_36_216# 0.01fF
C55896 INVX1_LOC_90/A INVX1_LOC_69/Y 0.07fF
C55897 INVX1_LOC_147/Y INVX1_LOC_22/A 0.48fF
C55898 NAND2X1_LOC_337/B NOR2X1_LOC_841/a_36_216# 0.00fF
C55899 NOR2X1_LOC_136/Y NAND2X1_LOC_211/Y 0.03fF
C55900 NOR2X1_LOC_74/A NOR2X1_LOC_703/A 0.00fF
C55901 NOR2X1_LOC_19/B INPUT_0 0.32fF
C55902 INVX1_LOC_191/Y INVX1_LOC_77/Y 0.04fF
C55903 INVX1_LOC_22/A INVX1_LOC_20/A 3.26fF
C55904 NAND2X1_LOC_205/A NAND2X1_LOC_203/a_36_24# 0.02fF
C55905 NOR2X1_LOC_716/B INVX1_LOC_70/A 0.03fF
C55906 NOR2X1_LOC_272/Y INVX1_LOC_78/A 0.03fF
C55907 INVX1_LOC_290/A INVX1_LOC_76/A 0.19fF
C55908 INVX1_LOC_33/A NAND2X1_LOC_93/B 0.66fF
C55909 INVX1_LOC_58/A NAND2X1_LOC_9/Y 0.02fF
C55910 INVX1_LOC_64/A NOR2X1_LOC_529/a_36_216# 0.00fF
C55911 INVX1_LOC_41/A NAND2X1_LOC_487/a_36_24# 0.00fF
C55912 INVX1_LOC_24/A NOR2X1_LOC_813/a_36_216# 0.02fF
C55913 INVX1_LOC_58/A INVX1_LOC_233/A 0.07fF
C55914 INVX1_LOC_13/A NOR2X1_LOC_112/a_36_216# 0.02fF
C55915 NOR2X1_LOC_433/A NOR2X1_LOC_841/A 0.10fF
C55916 INVX1_LOC_104/A INVX1_LOC_274/A 0.08fF
C55917 NAND2X1_LOC_859/Y NAND2X1_LOC_242/a_36_24# 0.02fF
C55918 NAND2X1_LOC_474/Y NOR2X1_LOC_278/Y 0.07fF
C55919 INVX1_LOC_54/Y NAND2X1_LOC_204/a_36_24# 0.00fF
C55920 INVX1_LOC_34/A NOR2X1_LOC_216/B 2.52fF
C55921 INVX1_LOC_136/A NAND2X1_LOC_63/Y 0.03fF
C55922 NAND2X1_LOC_213/A INVX1_LOC_78/A 0.31fF
C55923 INVX1_LOC_40/A NOR2X1_LOC_536/A 0.05fF
C55924 NOR2X1_LOC_272/Y NOR2X1_LOC_65/B 0.10fF
C55925 NAND2X1_LOC_453/a_36_24# NOR2X1_LOC_435/A 0.00fF
C55926 NAND2X1_LOC_537/Y INVX1_LOC_273/A -0.02fF
C55927 INVX1_LOC_24/A NAND2X1_LOC_773/B 0.50fF
C55928 INVX1_LOC_225/A NOR2X1_LOC_831/B 0.11fF
C55929 INVX1_LOC_61/A NAND2X1_LOC_74/B 0.04fF
C55930 INVX1_LOC_56/Y NOR2X1_LOC_271/Y 0.01fF
C55931 INVX1_LOC_170/A NAND2X1_LOC_74/a_36_24# 0.01fF
C55932 INVX1_LOC_298/Y INVX1_LOC_269/A 0.02fF
C55933 INVX1_LOC_58/A NOR2X1_LOC_798/A 0.03fF
C55934 INVX1_LOC_314/Y INVX1_LOC_19/A 0.03fF
C55935 NOR2X1_LOC_52/B NOR2X1_LOC_841/A 0.01fF
C55936 INPUT_0 NOR2X1_LOC_528/Y 0.10fF
C55937 NAND2X1_LOC_364/A INVX1_LOC_42/A 0.07fF
C55938 INVX1_LOC_40/A NOR2X1_LOC_655/Y 0.02fF
C55939 NOR2X1_LOC_552/A NOR2X1_LOC_336/a_36_216# 0.01fF
C55940 NOR2X1_LOC_835/B INVX1_LOC_160/A 0.10fF
C55941 NOR2X1_LOC_701/Y INVX1_LOC_118/A 0.01fF
C55942 NOR2X1_LOC_759/a_36_216# INVX1_LOC_109/Y 0.00fF
C55943 NOR2X1_LOC_316/Y NAND2X1_LOC_572/B 0.03fF
C55944 NOR2X1_LOC_92/Y INVX1_LOC_57/A 0.18fF
C55945 INVX1_LOC_40/A NAND2X1_LOC_93/B 0.98fF
C55946 NOR2X1_LOC_246/A INVX1_LOC_33/Y 0.03fF
C55947 NOR2X1_LOC_242/A NAND2X1_LOC_363/B 0.46fF
C55948 INVX1_LOC_157/A INVX1_LOC_38/A 0.32fF
C55949 INVX1_LOC_286/Y NAND2X1_LOC_444/B 0.02fF
C55950 INVX1_LOC_24/Y INVX1_LOC_57/A 0.04fF
C55951 NAND2X1_LOC_192/B NOR2X1_LOC_383/B 0.02fF
C55952 INVX1_LOC_53/Y INVX1_LOC_131/Y 0.07fF
C55953 NOR2X1_LOC_631/B NOR2X1_LOC_208/A 0.03fF
C55954 INVX1_LOC_208/A NOR2X1_LOC_155/A 0.01fF
C55955 NOR2X1_LOC_274/B INVX1_LOC_4/A 0.39fF
C55956 D_INPUT_1 NOR2X1_LOC_468/Y 0.07fF
C55957 NOR2X1_LOC_15/Y NOR2X1_LOC_15/a_36_216# 0.03fF
C55958 NOR2X1_LOC_557/A INVX1_LOC_125/Y 0.50fF
C55959 NOR2X1_LOC_516/B NOR2X1_LOC_155/A 0.01fF
C55960 D_INPUT_1 NAND2X1_LOC_190/Y 0.01fF
C55961 NOR2X1_LOC_15/Y NAND2X1_LOC_860/A 0.20fF
C55962 INVX1_LOC_313/Y NOR2X1_LOC_122/a_36_216# 0.00fF
C55963 NAND2X1_LOC_863/A VDD -0.00fF
C55964 NOR2X1_LOC_254/Y INVX1_LOC_99/A 0.07fF
C55965 NOR2X1_LOC_473/B NOR2X1_LOC_331/B 0.01fF
C55966 INVX1_LOC_299/A NOR2X1_LOC_405/Y 0.07fF
C55967 NAND2X1_LOC_650/B NOR2X1_LOC_74/A 0.03fF
C55968 INVX1_LOC_24/A NOR2X1_LOC_393/Y 0.01fF
C55969 INVX1_LOC_100/A INVX1_LOC_20/A 0.03fF
C55970 NOR2X1_LOC_569/Y NOR2X1_LOC_197/B 0.10fF
C55971 INVX1_LOC_144/A NAND2X1_LOC_211/Y 0.02fF
C55972 INVX1_LOC_40/A NOR2X1_LOC_649/B 0.04fF
C55973 NOR2X1_LOC_595/Y INVX1_LOC_91/A -0.00fF
C55974 NAND2X1_LOC_741/B NOR2X1_LOC_25/Y 0.02fF
C55975 NOR2X1_LOC_382/Y NOR2X1_LOC_29/a_36_216# 0.00fF
C55976 INVX1_LOC_35/A INVX1_LOC_14/A 0.80fF
C55977 NOR2X1_LOC_208/A INVX1_LOC_37/A 0.05fF
C55978 INVX1_LOC_10/A INVX1_LOC_180/Y 0.04fF
C55979 INVX1_LOC_40/A INVX1_LOC_3/A 1.98fF
C55980 NAND2X1_LOC_364/A INVX1_LOC_78/A 0.10fF
C55981 NAND2X1_LOC_218/B INVX1_LOC_4/A 0.01fF
C55982 NOR2X1_LOC_457/A INVX1_LOC_53/A 0.07fF
C55983 NOR2X1_LOC_403/B NOR2X1_LOC_38/B 0.14fF
C55984 NOR2X1_LOC_256/Y NOR2X1_LOC_813/Y 0.03fF
C55985 D_INPUT_2 NOR2X1_LOC_38/B 0.03fF
C55986 INVX1_LOC_316/Y NOR2X1_LOC_23/a_36_216# 0.00fF
C55987 NOR2X1_LOC_130/A NAND2X1_LOC_434/Y 0.01fF
C55988 INVX1_LOC_21/A NOR2X1_LOC_173/Y 0.03fF
C55989 NOR2X1_LOC_778/B INVX1_LOC_19/A 0.05fF
C55990 INVX1_LOC_45/Y INVX1_LOC_94/Y 0.11fF
C55991 INVX1_LOC_115/Y INVX1_LOC_91/A 0.01fF
C55992 NOR2X1_LOC_577/Y INVX1_LOC_4/A 0.09fF
C55993 NAND2X1_LOC_848/a_36_24# INVX1_LOC_84/A 0.00fF
C55994 NOR2X1_LOC_598/B NOR2X1_LOC_160/B 0.58fF
C55995 INVX1_LOC_21/A NOR2X1_LOC_321/Y 0.01fF
C55996 NOR2X1_LOC_468/Y NOR2X1_LOC_652/Y 0.01fF
C55997 NOR2X1_LOC_188/a_36_216# INVX1_LOC_84/A 0.00fF
C55998 NOR2X1_LOC_33/A NOR2X1_LOC_814/A 0.12fF
C55999 NOR2X1_LOC_256/Y INVX1_LOC_280/A 0.03fF
C56000 NOR2X1_LOC_433/A INVX1_LOC_128/A -0.01fF
C56001 INVX1_LOC_63/Y INVX1_LOC_15/A 0.03fF
C56002 NOR2X1_LOC_65/B NAND2X1_LOC_364/A 2.21fF
C56003 NAND2X1_LOC_725/A NAND2X1_LOC_550/A 0.15fF
C56004 INVX1_LOC_6/A INVX1_LOC_77/Y 0.17fF
C56005 D_INPUT_0 INVX1_LOC_285/A 0.07fF
C56006 NOR2X1_LOC_589/A INVX1_LOC_186/Y 0.00fF
C56007 NAND2X1_LOC_276/Y INVX1_LOC_4/Y 0.08fF
C56008 INVX1_LOC_30/A INVX1_LOC_53/A 1.12fF
C56009 NOR2X1_LOC_99/B NOR2X1_LOC_673/A 0.01fF
C56010 INVX1_LOC_314/Y INVX1_LOC_26/Y 0.07fF
C56011 NAND2X1_LOC_332/Y INVX1_LOC_128/Y 0.01fF
C56012 NOR2X1_LOC_348/B INVX1_LOC_4/A 0.07fF
C56013 NOR2X1_LOC_188/A INVX1_LOC_9/A 0.18fF
C56014 INVX1_LOC_69/Y INVX1_LOC_38/A 0.07fF
C56015 NOR2X1_LOC_391/a_36_216# INVX1_LOC_280/A 0.01fF
C56016 NOR2X1_LOC_816/a_36_216# INVX1_LOC_161/Y 0.01fF
C56017 D_INPUT_0 NOR2X1_LOC_814/A 0.04fF
C56018 NAND2X1_LOC_763/B INVX1_LOC_53/A 0.35fF
C56019 NOR2X1_LOC_548/B INVX1_LOC_9/A 0.01fF
C56020 NOR2X1_LOC_389/a_36_216# INVX1_LOC_285/A 0.01fF
C56021 NOR2X1_LOC_15/Y NAND2X1_LOC_537/Y 0.07fF
C56022 NOR2X1_LOC_186/Y NAND2X1_LOC_352/B 0.01fF
C56023 D_INPUT_1 INVX1_LOC_62/Y 0.14fF
C56024 INVX1_LOC_234/A NOR2X1_LOC_84/B 0.06fF
C56025 NOR2X1_LOC_389/A NOR2X1_LOC_652/Y 0.10fF
C56026 INVX1_LOC_131/A NOR2X1_LOC_216/B 0.20fF
C56027 NAND2X1_LOC_837/Y INVX1_LOC_57/A 0.07fF
C56028 NAND2X1_LOC_466/A NAND2X1_LOC_470/B 0.02fF
C56029 INVX1_LOC_243/A NOR2X1_LOC_467/A 0.05fF
C56030 D_INPUT_1 NOR2X1_LOC_596/A 0.03fF
C56031 NOR2X1_LOC_86/A INVX1_LOC_42/A 0.07fF
C56032 NOR2X1_LOC_545/B INVX1_LOC_117/A 0.13fF
C56033 INPUT_0 NOR2X1_LOC_216/B 0.15fF
C56034 INVX1_LOC_162/A NAND2X1_LOC_288/B 0.12fF
C56035 INVX1_LOC_88/A NOR2X1_LOC_218/A 0.00fF
C56036 NOR2X1_LOC_724/Y INVX1_LOC_19/A 0.01fF
C56037 NAND2X1_LOC_198/B NOR2X1_LOC_109/Y 0.06fF
C56038 INVX1_LOC_41/A INVX1_LOC_57/A 0.31fF
C56039 NAND2X1_LOC_214/B INVX1_LOC_72/Y 0.01fF
C56040 NOR2X1_LOC_315/Y NOR2X1_LOC_693/Y 0.09fF
C56041 NAND2X1_LOC_11/Y INVX1_LOC_78/A 0.00fF
C56042 INVX1_LOC_22/A INVX1_LOC_4/A 0.21fF
C56043 NOR2X1_LOC_68/A INVX1_LOC_50/Y 0.24fF
C56044 INVX1_LOC_39/A INVX1_LOC_136/A 0.13fF
C56045 NOR2X1_LOC_328/Y NOR2X1_LOC_329/Y 0.04fF
C56046 INVX1_LOC_21/A INVX1_LOC_205/A 0.59fF
C56047 NOR2X1_LOC_32/B NOR2X1_LOC_672/Y 0.01fF
C56048 NOR2X1_LOC_598/B NOR2X1_LOC_544/a_36_216# 0.14fF
C56049 NAND2X1_LOC_53/Y NOR2X1_LOC_197/A 0.03fF
C56050 NOR2X1_LOC_705/B INVX1_LOC_11/A 0.02fF
C56051 NAND2X1_LOC_602/a_36_24# NOR2X1_LOC_331/B 0.00fF
C56052 NOR2X1_LOC_261/Y INVX1_LOC_63/Y 0.30fF
C56053 INVX1_LOC_90/A NOR2X1_LOC_89/A 0.16fF
C56054 NAND2X1_LOC_354/Y NOR2X1_LOC_173/Y 0.18fF
C56055 INVX1_LOC_64/A NOR2X1_LOC_577/Y 0.13fF
C56056 NAND2X1_LOC_833/Y NAND2X1_LOC_793/B 0.01fF
C56057 NOR2X1_LOC_91/A NAND2X1_LOC_717/Y 0.03fF
C56058 NAND2X1_LOC_477/A INVX1_LOC_57/A 0.03fF
C56059 INVX1_LOC_49/A NOR2X1_LOC_665/Y 0.02fF
C56060 NOR2X1_LOC_389/B NOR2X1_LOC_89/A 0.01fF
C56061 NOR2X1_LOC_454/Y NOR2X1_LOC_194/a_36_216# 0.01fF
C56062 INVX1_LOC_21/A NOR2X1_LOC_607/A 0.03fF
C56063 NAND2X1_LOC_214/B NOR2X1_LOC_643/Y 0.00fF
C56064 INVX1_LOC_149/Y INVX1_LOC_58/Y 0.10fF
C56065 NOR2X1_LOC_186/Y NAND2X1_LOC_573/a_36_24# 0.00fF
C56066 NOR2X1_LOC_538/B NOR2X1_LOC_641/B 0.16fF
C56067 INVX1_LOC_266/Y INVX1_LOC_105/Y 0.01fF
C56068 INVX1_LOC_1/Y NAND2X1_LOC_221/a_36_24# 0.01fF
C56069 INVX1_LOC_58/A NOR2X1_LOC_718/a_36_216# 0.00fF
C56070 NOR2X1_LOC_270/Y NOR2X1_LOC_666/A 0.26fF
C56071 NOR2X1_LOC_45/B INVX1_LOC_260/Y 0.07fF
C56072 INVX1_LOC_2/A NOR2X1_LOC_414/Y 0.14fF
C56073 NOR2X1_LOC_355/A NOR2X1_LOC_609/Y 0.02fF
C56074 NOR2X1_LOC_465/a_36_216# NOR2X1_LOC_348/B 0.01fF
C56075 NAND2X1_LOC_516/a_36_24# NOR2X1_LOC_816/A 0.00fF
C56076 INVX1_LOC_64/A NOR2X1_LOC_629/B 0.01fF
C56077 NOR2X1_LOC_538/B NOR2X1_LOC_751/Y 0.06fF
C56078 INVX1_LOC_1/A NOR2X1_LOC_324/Y 0.01fF
C56079 NOR2X1_LOC_91/A INVX1_LOC_16/A 0.19fF
C56080 INVX1_LOC_64/A NOR2X1_LOC_348/B 0.32fF
C56081 NOR2X1_LOC_524/a_36_216# INVX1_LOC_270/Y 0.02fF
C56082 NOR2X1_LOC_393/a_36_216# INVX1_LOC_42/A 0.01fF
C56083 NOR2X1_LOC_544/A NOR2X1_LOC_858/A 0.03fF
C56084 INVX1_LOC_13/A INVX1_LOC_23/Y 0.19fF
C56085 NOR2X1_LOC_598/B INVX1_LOC_189/A -0.02fF
C56086 NOR2X1_LOC_689/Y NAND2X1_LOC_853/Y 0.18fF
C56087 INVX1_LOC_45/A NAND2X1_LOC_171/a_36_24# 0.01fF
C56088 INVX1_LOC_232/A NOR2X1_LOC_646/B 0.00fF
C56089 INVX1_LOC_53/Y INVX1_LOC_270/A 0.00fF
C56090 INVX1_LOC_269/A INVX1_LOC_228/A 0.03fF
C56091 NAND2X1_LOC_30/Y NAND2X1_LOC_588/B 0.16fF
C56092 INVX1_LOC_208/A NOR2X1_LOC_125/Y 0.02fF
C56093 INVX1_LOC_35/A INVX1_LOC_111/Y 0.01fF
C56094 NOR2X1_LOC_295/Y NOR2X1_LOC_652/Y 0.00fF
C56095 NAND2X1_LOC_213/A NOR2X1_LOC_152/Y 0.09fF
C56096 NAND2X1_LOC_633/Y INVX1_LOC_70/A 0.00fF
C56097 INVX1_LOC_224/Y NOR2X1_LOC_62/a_36_216# 0.00fF
C56098 NAND2X1_LOC_182/A INVX1_LOC_306/Y 0.00fF
C56099 NOR2X1_LOC_155/A NAND2X1_LOC_211/Y 0.04fF
C56100 NAND2X1_LOC_363/B NOR2X1_LOC_78/B 0.03fF
C56101 INVX1_LOC_2/A NOR2X1_LOC_665/Y 0.12fF
C56102 NAND2X1_LOC_762/a_36_24# INVX1_LOC_174/A 0.01fF
C56103 NOR2X1_LOC_735/Y INVX1_LOC_4/A 0.01fF
C56104 NAND2X1_LOC_213/A INVX1_LOC_113/Y 0.00fF
C56105 INVX1_LOC_174/A INVX1_LOC_18/A 0.08fF
C56106 INVX1_LOC_233/Y NAND2X1_LOC_374/Y 0.10fF
C56107 INVX1_LOC_201/Y INVX1_LOC_252/A 0.03fF
C56108 NOR2X1_LOC_186/Y NAND2X1_LOC_357/B 0.15fF
C56109 NOR2X1_LOC_96/a_36_216# INVX1_LOC_280/A 0.01fF
C56110 INVX1_LOC_16/A INVX1_LOC_23/A 0.56fF
C56111 INVX1_LOC_220/Y NOR2X1_LOC_383/B 0.01fF
C56112 NOR2X1_LOC_557/A INVX1_LOC_19/A 0.04fF
C56113 INVX1_LOC_25/A NOR2X1_LOC_719/A 0.01fF
C56114 NOR2X1_LOC_576/B NOR2X1_LOC_829/A 0.33fF
C56115 NAND2X1_LOC_12/a_36_24# INVX1_LOC_174/A 0.01fF
C56116 NOR2X1_LOC_188/A NOR2X1_LOC_861/Y 0.07fF
C56117 NOR2X1_LOC_598/B NOR2X1_LOC_516/B 0.26fF
C56118 NOR2X1_LOC_156/a_36_216# INVX1_LOC_117/A 0.01fF
C56119 NOR2X1_LOC_845/A NAND2X1_LOC_207/B 0.21fF
C56120 INVX1_LOC_269/A NOR2X1_LOC_516/a_36_216# 0.01fF
C56121 INVX1_LOC_27/A INVX1_LOC_266/Y 0.17fF
C56122 NAND2X1_LOC_472/Y NOR2X1_LOC_197/B 0.10fF
C56123 INVX1_LOC_25/A NOR2X1_LOC_561/Y 0.13fF
C56124 INVX1_LOC_93/A NAND2X1_LOC_231/Y 0.02fF
C56125 INVX1_LOC_88/A INVX1_LOC_155/Y 0.11fF
C56126 INVX1_LOC_25/A INVX1_LOC_7/A 0.07fF
C56127 NOR2X1_LOC_454/Y NOR2X1_LOC_300/Y 0.04fF
C56128 INVX1_LOC_269/A INVX1_LOC_8/A 0.10fF
C56129 NAND2X1_LOC_120/a_36_24# NOR2X1_LOC_759/Y 0.01fF
C56130 INVX1_LOC_64/A INVX1_LOC_22/A 0.31fF
C56131 INVX1_LOC_11/A NOR2X1_LOC_172/Y 0.03fF
C56132 NOR2X1_LOC_78/B NOR2X1_LOC_791/Y 0.05fF
C56133 NAND2X1_LOC_787/A NAND2X1_LOC_392/Y 0.20fF
C56134 NAND2X1_LOC_475/Y INVX1_LOC_46/A 0.10fF
C56135 NOR2X1_LOC_807/B INVX1_LOC_33/A 0.15fF
C56136 INVX1_LOC_256/A INVX1_LOC_33/A 0.16fF
C56137 NAND2X1_LOC_724/A NAND2X1_LOC_357/B 0.89fF
C56138 INVX1_LOC_224/Y NOR2X1_LOC_76/A 0.87fF
C56139 INVX1_LOC_36/A NAND2X1_LOC_198/B 0.64fF
C56140 INVX1_LOC_279/A NOR2X1_LOC_678/A 0.07fF
C56141 NOR2X1_LOC_609/A INVX1_LOC_223/A 0.25fF
C56142 NOR2X1_LOC_189/A NAND2X1_LOC_188/a_36_24# 0.02fF
C56143 INVX1_LOC_1/A NAND2X1_LOC_629/Y 0.01fF
C56144 NAND2X1_LOC_725/Y NAND2X1_LOC_379/a_36_24# 0.08fF
C56145 NOR2X1_LOC_91/A INVX1_LOC_28/A 0.60fF
C56146 INVX1_LOC_136/A INVX1_LOC_61/A 0.23fF
C56147 INVX1_LOC_37/A INVX1_LOC_63/A 0.16fF
C56148 INVX1_LOC_93/A NAND2X1_LOC_858/a_36_24# 0.01fF
C56149 INVX1_LOC_36/A NAND2X1_LOC_368/a_36_24# 0.00fF
C56150 NOR2X1_LOC_405/A INVX1_LOC_42/A 0.03fF
C56151 INVX1_LOC_184/A INVX1_LOC_30/A 0.06fF
C56152 INVX1_LOC_287/Y NOR2X1_LOC_708/Y 0.01fF
C56153 NOR2X1_LOC_276/B NOR2X1_LOC_270/Y 0.06fF
C56154 NOR2X1_LOC_267/A NAND2X1_LOC_198/B 0.13fF
C56155 NAND2X1_LOC_363/B INVX1_LOC_83/A 0.07fF
C56156 INVX1_LOC_277/A INVX1_LOC_77/A 0.24fF
C56157 NAND2X1_LOC_848/A INVX1_LOC_285/A 0.10fF
C56158 INVX1_LOC_5/A NOR2X1_LOC_32/Y 0.01fF
C56159 INVX1_LOC_286/Y INVX1_LOC_209/Y 0.03fF
C56160 INVX1_LOC_243/A INVX1_LOC_1/A 0.07fF
C56161 INVX1_LOC_35/A NOR2X1_LOC_137/A 0.03fF
C56162 NOR2X1_LOC_76/A NAND2X1_LOC_793/B 0.03fF
C56163 NAND2X1_LOC_758/a_36_24# INVX1_LOC_159/A 0.01fF
C56164 INVX1_LOC_83/A NOR2X1_LOC_640/a_36_216# 0.00fF
C56165 INVX1_LOC_225/A NAND2X1_LOC_352/B 0.24fF
C56166 INVX1_LOC_28/A INVX1_LOC_23/A 1.76fF
C56167 INVX1_LOC_69/Y INVX1_LOC_18/Y 0.09fF
C56168 NOR2X1_LOC_15/Y INVX1_LOC_172/Y 0.07fF
C56169 NOR2X1_LOC_209/Y D_GATE_741 0.00fF
C56170 NAND2X1_LOC_537/Y NAND2X1_LOC_840/B 0.01fF
C56171 INVX1_LOC_12/Y INVX1_LOC_29/A 0.01fF
C56172 NOR2X1_LOC_82/A INVX1_LOC_256/Y 0.07fF
C56173 INVX1_LOC_286/A NOR2X1_LOC_301/A 0.29fF
C56174 NOR2X1_LOC_78/B NOR2X1_LOC_457/A 0.36fF
C56175 NOR2X1_LOC_45/B NAND2X1_LOC_471/Y 0.01fF
C56176 INVX1_LOC_153/A INVX1_LOC_18/A 0.06fF
C56177 INVX1_LOC_266/A NOR2X1_LOC_570/Y 0.17fF
C56178 INVX1_LOC_14/A NOR2X1_LOC_121/A 0.09fF
C56179 NAND2X1_LOC_624/A INVX1_LOC_253/Y 0.07fF
C56180 NAND2X1_LOC_53/Y INVX1_LOC_83/Y 0.04fF
C56181 NOR2X1_LOC_113/B INVX1_LOC_270/A 0.10fF
C56182 NOR2X1_LOC_598/B NOR2X1_LOC_706/A 0.00fF
C56183 NOR2X1_LOC_113/A INVX1_LOC_78/A 0.01fF
C56184 NOR2X1_LOC_405/A INVX1_LOC_78/A 0.07fF
C56185 INVX1_LOC_172/A NAND2X1_LOC_169/a_36_24# 0.01fF
C56186 INVX1_LOC_76/A NOR2X1_LOC_467/A 0.46fF
C56187 NAND2X1_LOC_851/a_36_24# NOR2X1_LOC_654/A 0.01fF
C56188 NOR2X1_LOC_174/a_36_216# NOR2X1_LOC_500/B 0.13fF
C56189 NAND2X1_LOC_383/a_36_24# INVX1_LOC_309/A 0.00fF
C56190 NOR2X1_LOC_557/A INVX1_LOC_26/Y 0.10fF
C56191 INVX1_LOC_5/A INVX1_LOC_311/Y 0.19fF
C56192 NOR2X1_LOC_743/Y INVX1_LOC_63/A 0.23fF
C56193 INVX1_LOC_40/Y NOR2X1_LOC_818/Y 0.06fF
C56194 NOR2X1_LOC_68/A NOR2X1_LOC_6/B 0.15fF
C56195 INVX1_LOC_188/Y NAND2X1_LOC_454/Y 0.00fF
C56196 NOR2X1_LOC_89/A INVX1_LOC_38/A 0.42fF
C56197 NAND2X1_LOC_198/B NOR2X1_LOC_309/Y 0.10fF
C56198 INVX1_LOC_45/A INVX1_LOC_164/Y 0.16fF
C56199 NOR2X1_LOC_78/B INVX1_LOC_30/A 0.19fF
C56200 NOR2X1_LOC_172/Y NOR2X1_LOC_433/A 0.02fF
C56201 NOR2X1_LOC_334/Y NOR2X1_LOC_136/a_36_216# 0.00fF
C56202 INVX1_LOC_13/A NAND2X1_LOC_563/a_36_24# 0.00fF
C56203 INVX1_LOC_18/A INVX1_LOC_259/A 0.08fF
C56204 NOR2X1_LOC_443/Y NOR2X1_LOC_78/A 0.02fF
C56205 NOR2X1_LOC_606/Y INVX1_LOC_40/A 0.01fF
C56206 INVX1_LOC_78/A NOR2X1_LOC_682/a_36_216# 0.00fF
C56207 NOR2X1_LOC_355/B NOR2X1_LOC_493/A 0.00fF
C56208 NOR2X1_LOC_65/B NOR2X1_LOC_405/A 0.21fF
C56209 VDD NAND2X1_LOC_444/B 0.01fF
C56210 INVX1_LOC_17/A NOR2X1_LOC_373/Y 0.01fF
C56211 INVX1_LOC_31/A INVX1_LOC_16/A 4.09fF
C56212 NOR2X1_LOC_361/B NOR2X1_LOC_106/A 0.36fF
C56213 VDD NOR2X1_LOC_334/Y 3.20fF
C56214 NOR2X1_LOC_67/A NOR2X1_LOC_791/B 0.07fF
C56215 NAND2X1_LOC_763/B NAND2X1_LOC_588/a_36_24# 0.00fF
C56216 GATE_741 NOR2X1_LOC_380/Y 0.03fF
C56217 NOR2X1_LOC_45/B NOR2X1_LOC_696/Y 0.05fF
C56218 INVX1_LOC_277/A NOR2X1_LOC_687/Y 0.07fF
C56219 NOR2X1_LOC_598/B INVX1_LOC_315/Y 0.13fF
C56220 NAND2X1_LOC_803/B D_INPUT_0 0.85fF
C56221 INVX1_LOC_249/A INVX1_LOC_266/Y 0.35fF
C56222 NOR2X1_LOC_172/Y INVX1_LOC_151/A 0.00fF
C56223 INVX1_LOC_36/A INVX1_LOC_53/Y 0.07fF
C56224 NOR2X1_LOC_668/Y NOR2X1_LOC_35/Y 0.01fF
C56225 INVX1_LOC_224/A INVX1_LOC_90/A 0.05fF
C56226 INVX1_LOC_278/Y NOR2X1_LOC_518/Y 0.02fF
C56227 NOR2X1_LOC_103/Y NOR2X1_LOC_76/A 0.04fF
C56228 INVX1_LOC_24/A INVX1_LOC_143/A 0.07fF
C56229 INVX1_LOC_292/A NAND2X1_LOC_656/Y 0.03fF
C56230 INVX1_LOC_93/A INPUT_0 0.40fF
C56231 INVX1_LOC_34/A NOR2X1_LOC_84/A 0.08fF
C56232 D_INPUT_6 NAND2X1_LOC_51/B 0.03fF
C56233 INVX1_LOC_11/A INVX1_LOC_90/A 1.73fF
C56234 NOR2X1_LOC_172/Y NOR2X1_LOC_52/B 0.06fF
C56235 NAND2X1_LOC_35/Y NOR2X1_LOC_526/a_36_216# 0.01fF
C56236 INVX1_LOC_11/A NAND2X1_LOC_769/a_36_24# 0.00fF
C56237 INVX1_LOC_2/A NAND2X1_LOC_567/Y 0.06fF
C56238 INVX1_LOC_36/A NOR2X1_LOC_665/A 0.03fF
C56239 NAND2X1_LOC_569/A NAND2X1_LOC_465/Y 0.02fF
C56240 NOR2X1_LOC_15/Y NAND2X1_LOC_855/Y 0.06fF
C56241 NOR2X1_LOC_716/B NOR2X1_LOC_316/Y 0.03fF
C56242 INVX1_LOC_30/A NAND2X1_LOC_392/Y 0.03fF
C56243 INVX1_LOC_11/A NOR2X1_LOC_389/B 0.08fF
C56244 NOR2X1_LOC_590/A D_INPUT_0 0.14fF
C56245 INVX1_LOC_33/Y NAND2X1_LOC_175/Y 0.02fF
C56246 NAND2X1_LOC_563/A INVX1_LOC_228/A 0.19fF
C56247 NOR2X1_LOC_627/Y INVX1_LOC_113/Y 0.01fF
C56248 INVX1_LOC_49/A NAND2X1_LOC_342/Y 0.00fF
C56249 INVX1_LOC_36/A NOR2X1_LOC_781/B 0.16fF
C56250 NOR2X1_LOC_589/A INVX1_LOC_18/A 0.09fF
C56251 INVX1_LOC_23/A NOR2X1_LOC_35/Y 0.01fF
C56252 INVX1_LOC_41/Y INVX1_LOC_25/Y 0.03fF
C56253 INVX1_LOC_36/A INVX1_LOC_145/Y 0.04fF
C56254 INVX1_LOC_225/A NAND2X1_LOC_357/B 0.03fF
C56255 NAND2X1_LOC_787/A NOR2X1_LOC_164/Y 0.01fF
C56256 NOR2X1_LOC_219/Y NOR2X1_LOC_208/Y 0.05fF
C56257 NOR2X1_LOC_252/a_36_216# NOR2X1_LOC_238/Y 0.00fF
C56258 NAND2X1_LOC_565/B INVX1_LOC_24/A 0.01fF
C56259 NOR2X1_LOC_67/Y NOR2X1_LOC_243/B 0.13fF
C56260 INVX1_LOC_25/A INVX1_LOC_76/A 0.15fF
C56261 INVX1_LOC_83/A INVX1_LOC_30/A 0.23fF
C56262 INVX1_LOC_145/A INVX1_LOC_53/Y 0.08fF
C56263 NOR2X1_LOC_212/a_36_216# INVX1_LOC_91/A 0.02fF
C56264 VDD NAND2X1_LOC_464/B 0.06fF
C56265 NAND2X1_LOC_141/A NOR2X1_LOC_516/Y 0.05fF
C56266 NOR2X1_LOC_331/B NOR2X1_LOC_464/Y 0.02fF
C56267 INVX1_LOC_161/Y NAND2X1_LOC_123/Y 0.07fF
C56268 NOR2X1_LOC_557/Y INVX1_LOC_143/A 0.01fF
C56269 INVX1_LOC_1/A NOR2X1_LOC_835/B 0.85fF
C56270 NOR2X1_LOC_230/Y INVX1_LOC_89/A 0.06fF
C56271 NAND2X1_LOC_763/B INVX1_LOC_83/A 0.03fF
C56272 NAND2X1_LOC_639/A NOR2X1_LOC_635/B 0.27fF
C56273 INVX1_LOC_45/A NOR2X1_LOC_76/A 0.02fF
C56274 NAND2X1_LOC_550/A NAND2X1_LOC_560/A 0.01fF
C56275 INVX1_LOC_11/A NAND2X1_LOC_348/A 0.10fF
C56276 INVX1_LOC_1/A INVX1_LOC_303/Y 0.01fF
C56277 NOR2X1_LOC_208/Y NOR2X1_LOC_665/A 0.08fF
C56278 INVX1_LOC_28/A INVX1_LOC_31/A 0.23fF
C56279 NAND2X1_LOC_787/A INVX1_LOC_46/A 0.06fF
C56280 INVX1_LOC_45/A NOR2X1_LOC_180/B 0.07fF
C56281 NOR2X1_LOC_67/A NOR2X1_LOC_124/B 0.00fF
C56282 INVX1_LOC_259/Y INVX1_LOC_14/Y 0.01fF
C56283 NAND2X1_LOC_731/Y INVX1_LOC_10/A 0.18fF
C56284 NAND2X1_LOC_89/a_36_24# INVX1_LOC_120/A 0.00fF
C56285 NAND2X1_LOC_543/Y NOR2X1_LOC_716/B 0.03fF
C56286 INVX1_LOC_77/A INVX1_LOC_174/Y 0.00fF
C56287 INVX1_LOC_171/A INVX1_LOC_18/A 0.00fF
C56288 NAND2X1_LOC_783/A INVX1_LOC_24/A 0.01fF
C56289 INVX1_LOC_145/A INVX1_LOC_145/Y 0.01fF
C56290 NOR2X1_LOC_301/A INVX1_LOC_54/A 0.09fF
C56291 NAND2X1_LOC_363/B INVX1_LOC_46/A 0.17fF
C56292 D_INPUT_3 NOR2X1_LOC_660/Y 0.15fF
C56293 INVX1_LOC_24/A NAND2X1_LOC_800/Y 0.00fF
C56294 INVX1_LOC_71/A NOR2X1_LOC_335/a_36_216# 0.00fF
C56295 NAND2X1_LOC_618/a_36_24# NOR2X1_LOC_660/Y 0.00fF
C56296 NAND2X1_LOC_347/B NOR2X1_LOC_78/A 0.55fF
C56297 INVX1_LOC_24/A NOR2X1_LOC_130/A 2.78fF
C56298 NOR2X1_LOC_168/B NAND2X1_LOC_118/a_36_24# 0.00fF
C56299 INVX1_LOC_17/A INVX1_LOC_286/A 0.09fF
C56300 INVX1_LOC_5/A NOR2X1_LOC_825/Y 0.60fF
C56301 NOR2X1_LOC_597/Y NOR2X1_LOC_599/A 0.02fF
C56302 NOR2X1_LOC_68/A NOR2X1_LOC_156/A 0.07fF
C56303 NOR2X1_LOC_309/Y INVX1_LOC_53/Y 1.94fF
C56304 INVX1_LOC_45/A INVX1_LOC_73/A 0.03fF
C56305 NAND2X1_LOC_382/a_36_24# NOR2X1_LOC_391/B 0.00fF
C56306 INVX1_LOC_71/A NOR2X1_LOC_76/A 0.02fF
C56307 INVX1_LOC_38/A NAND2X1_LOC_804/A 0.03fF
C56308 INVX1_LOC_157/A INVX1_LOC_33/A 0.06fF
C56309 NOR2X1_LOC_526/Y NAND2X1_LOC_374/Y 0.03fF
C56310 INVX1_LOC_13/A NAND2X1_LOC_116/A 0.07fF
C56311 INVX1_LOC_15/Y INVX1_LOC_172/Y 0.11fF
C56312 NOR2X1_LOC_180/B INVX1_LOC_71/A 0.07fF
C56313 NOR2X1_LOC_290/Y INVX1_LOC_16/A 0.02fF
C56314 NAND2X1_LOC_451/a_36_24# NAND2X1_LOC_451/Y 0.01fF
C56315 NOR2X1_LOC_554/A INVX1_LOC_29/A 0.01fF
C56316 INVX1_LOC_197/A INVX1_LOC_197/Y 0.15fF
C56317 INVX1_LOC_90/A NOR2X1_LOC_433/A 0.13fF
C56318 D_INPUT_0 NAND2X1_LOC_518/a_36_24# 0.00fF
C56319 NAND2X1_LOC_326/A NAND2X1_LOC_649/a_36_24# 0.01fF
C56320 NOR2X1_LOC_249/Y NOR2X1_LOC_34/a_36_216# 0.00fF
C56321 NAND2X1_LOC_72/B INVX1_LOC_63/A 0.03fF
C56322 NOR2X1_LOC_304/Y NOR2X1_LOC_536/A 0.02fF
C56323 INVX1_LOC_90/A NOR2X1_LOC_593/Y 0.07fF
C56324 INVX1_LOC_230/Y NOR2X1_LOC_45/B 0.03fF
C56325 INVX1_LOC_1/A INVX1_LOC_76/A 0.25fF
C56326 NOR2X1_LOC_437/Y NAND2X1_LOC_123/Y 0.01fF
C56327 NOR2X1_LOC_220/A NOR2X1_LOC_553/Y 0.01fF
C56328 NOR2X1_LOC_612/a_36_216# INVX1_LOC_1/Y 0.00fF
C56329 INVX1_LOC_304/A NAND2X1_LOC_793/Y 0.04fF
C56330 INVX1_LOC_284/A INVX1_LOC_3/Y 0.09fF
C56331 INVX1_LOC_18/A INVX1_LOC_222/A 0.38fF
C56332 INVX1_LOC_58/A NAND2X1_LOC_243/B 0.25fF
C56333 NOR2X1_LOC_389/B NOR2X1_LOC_593/Y 0.02fF
C56334 INVX1_LOC_73/A INVX1_LOC_71/A 0.07fF
C56335 NOR2X1_LOC_334/Y INVX1_LOC_133/A 0.00fF
C56336 NOR2X1_LOC_315/Y NOR2X1_LOC_71/Y 0.03fF
C56337 NOR2X1_LOC_431/a_36_216# INVX1_LOC_144/A 0.01fF
C56338 INVX1_LOC_23/Y NAND2X1_LOC_489/Y 1.61fF
C56339 NOR2X1_LOC_721/a_36_216# NOR2X1_LOC_346/B 0.02fF
C56340 NAND2X1_LOC_799/A INVX1_LOC_20/A 0.03fF
C56341 INVX1_LOC_249/A INVX1_LOC_42/Y 0.02fF
C56342 NOR2X1_LOC_500/A INPUT_0 0.03fF
C56343 NAND2X1_LOC_785/A NAND2X1_LOC_861/Y 0.02fF
C56344 INVX1_LOC_64/A NOR2X1_LOC_88/A 0.00fF
C56345 INVX1_LOC_90/A NOR2X1_LOC_52/B 0.28fF
C56346 VDD INVX1_LOC_308/Y 0.21fF
C56347 INVX1_LOC_13/A INVX1_LOC_232/A 0.99fF
C56348 NOR2X1_LOC_86/A NAND2X1_LOC_859/B 0.03fF
C56349 INVX1_LOC_104/A NOR2X1_LOC_356/A 0.07fF
C56350 NOR2X1_LOC_457/A INVX1_LOC_46/A 0.16fF
C56351 INVX1_LOC_29/A NOR2X1_LOC_89/Y 0.03fF
C56352 NOR2X1_LOC_389/B NOR2X1_LOC_52/B 0.07fF
C56353 INVX1_LOC_58/A INVX1_LOC_119/Y 0.02fF
C56354 NAND2X1_LOC_859/Y INVX1_LOC_16/A 0.10fF
C56355 NOR2X1_LOC_89/A NAND2X1_LOC_223/A 0.03fF
C56356 NOR2X1_LOC_637/B INVX1_LOC_144/A 0.06fF
C56357 INVX1_LOC_164/Y NOR2X1_LOC_123/B 0.02fF
C56358 NAND2X1_LOC_856/A NAND2X1_LOC_729/B 0.00fF
C56359 NOR2X1_LOC_360/Y INVX1_LOC_91/A 0.17fF
C56360 INVX1_LOC_31/A NOR2X1_LOC_35/Y 0.28fF
C56361 NAND2X1_LOC_721/a_36_24# NAND2X1_LOC_807/Y 0.00fF
C56362 NAND2X1_LOC_717/Y NAND2X1_LOC_866/B 0.00fF
C56363 NAND2X1_LOC_552/A NOR2X1_LOC_88/Y 0.03fF
C56364 NAND2X1_LOC_807/B NOR2X1_LOC_301/A 1.00fF
C56365 NOR2X1_LOC_290/Y INVX1_LOC_28/A 0.02fF
C56366 INVX1_LOC_271/A INVX1_LOC_19/A 0.03fF
C56367 NOR2X1_LOC_473/B NOR2X1_LOC_366/B 0.11fF
C56368 INVX1_LOC_224/A INVX1_LOC_38/A 0.03fF
C56369 INPUT_0 NOR2X1_LOC_84/A 0.01fF
C56370 NOR2X1_LOC_68/A NOR2X1_LOC_124/A 0.02fF
C56371 INVX1_LOC_33/A INVX1_LOC_69/Y 0.26fF
C56372 NOR2X1_LOC_836/Y VDD 0.39fF
C56373 INVX1_LOC_21/A NAND2X1_LOC_798/B 0.07fF
C56374 INVX1_LOC_207/A INVX1_LOC_309/A 0.03fF
C56375 NOR2X1_LOC_717/B NOR2X1_LOC_730/Y 0.03fF
C56376 INVX1_LOC_36/A NOR2X1_LOC_585/Y 0.01fF
C56377 INVX1_LOC_11/A INVX1_LOC_38/A 0.24fF
C56378 INVX1_LOC_104/A NOR2X1_LOC_74/A 0.24fF
C56379 NAND2X1_LOC_803/B NAND2X1_LOC_848/A 0.67fF
C56380 NOR2X1_LOC_590/A NOR2X1_LOC_859/Y 0.00fF
C56381 NOR2X1_LOC_770/A INVX1_LOC_91/A 0.01fF
C56382 NAND2X1_LOC_363/B NOR2X1_LOC_68/Y 0.02fF
C56383 INVX1_LOC_30/A INVX1_LOC_46/A 0.93fF
C56384 INVX1_LOC_178/A NOR2X1_LOC_88/Y 0.10fF
C56385 NAND2X1_LOC_866/B INVX1_LOC_16/A 0.07fF
C56386 NAND2X1_LOC_552/A INVX1_LOC_84/A 0.89fF
C56387 INVX1_LOC_18/A INVX1_LOC_20/A 2.29fF
C56388 NAND2X1_LOC_88/a_36_24# NAND2X1_LOC_348/A 0.00fF
C56389 INVX1_LOC_5/A INVX1_LOC_84/A 2.36fF
C56390 INVX1_LOC_23/A INVX1_LOC_109/A 0.40fF
C56391 NOR2X1_LOC_793/Y INVX1_LOC_307/Y 0.00fF
C56392 NOR2X1_LOC_500/A NOR2X1_LOC_324/A 0.11fF
C56393 NOR2X1_LOC_405/A NOR2X1_LOC_152/Y 0.01fF
C56394 INVX1_LOC_104/A NOR2X1_LOC_9/Y 0.16fF
C56395 INVX1_LOC_10/A NOR2X1_LOC_525/Y 0.02fF
C56396 NAND2X1_LOC_35/Y NOR2X1_LOC_662/A 0.10fF
C56397 INVX1_LOC_64/A INVX1_LOC_186/Y 0.01fF
C56398 INVX1_LOC_17/A INVX1_LOC_54/A 1.04fF
C56399 NAND2X1_LOC_728/Y INVX1_LOC_20/A 0.30fF
C56400 NOR2X1_LOC_388/Y NOR2X1_LOC_355/B 0.01fF
C56401 INVX1_LOC_280/Y NAND2X1_LOC_863/A 0.02fF
C56402 INVX1_LOC_58/A INVX1_LOC_284/A 0.28fF
C56403 INVX1_LOC_207/A INVX1_LOC_91/A 0.04fF
C56404 INVX1_LOC_32/A INVX1_LOC_23/Y 0.07fF
C56405 NOR2X1_LOC_590/A NAND2X1_LOC_848/A 0.03fF
C56406 NAND2X1_LOC_574/A INVX1_LOC_252/A 0.03fF
C56407 NOR2X1_LOC_598/B NAND2X1_LOC_207/B 0.01fF
C56408 INVX1_LOC_38/Y NAND2X1_LOC_206/Y 0.02fF
C56409 NAND2X1_LOC_729/Y INVX1_LOC_76/A 0.00fF
C56410 INVX1_LOC_36/A INVX1_LOC_77/Y 0.07fF
C56411 NOR2X1_LOC_82/a_36_216# INVX1_LOC_12/Y 0.01fF
C56412 NOR2X1_LOC_523/B VDD -0.00fF
C56413 INVX1_LOC_178/A INVX1_LOC_84/A 0.15fF
C56414 NOR2X1_LOC_632/Y NOR2X1_LOC_736/Y 0.04fF
C56415 INVX1_LOC_13/A NOR2X1_LOC_775/Y 0.01fF
C56416 INVX1_LOC_28/A NAND2X1_LOC_859/Y 0.13fF
C56417 INVX1_LOC_72/A INVX1_LOC_117/A 0.09fF
C56418 INVX1_LOC_207/A INVX1_LOC_11/Y 0.07fF
C56419 INVX1_LOC_209/Y NOR2X1_LOC_56/Y 0.04fF
C56420 NAND2X1_LOC_221/a_36_24# INVX1_LOC_87/A 0.00fF
C56421 INVX1_LOC_142/Y INVX1_LOC_117/A 0.00fF
C56422 INVX1_LOC_100/A NAND2X1_LOC_850/Y 0.07fF
C56423 INVX1_LOC_5/A NAND2X1_LOC_651/B 0.14fF
C56424 NOR2X1_LOC_152/Y NOR2X1_LOC_682/a_36_216# 0.01fF
C56425 INVX1_LOC_289/Y NOR2X1_LOC_697/Y 0.11fF
C56426 INVX1_LOC_172/A INVX1_LOC_20/A 0.03fF
C56427 NOR2X1_LOC_217/a_36_216# NOR2X1_LOC_155/A 0.00fF
C56428 INVX1_LOC_282/A INVX1_LOC_22/A 0.05fF
C56429 D_GATE_579 NAND2X1_LOC_463/B 0.01fF
C56430 INVX1_LOC_165/A NAND2X1_LOC_99/A 0.02fF
C56431 INVX1_LOC_198/Y INVX1_LOC_117/A 0.08fF
C56432 NOR2X1_LOC_151/Y NOR2X1_LOC_730/Y 0.03fF
C56433 NAND2X1_LOC_357/B NAND2X1_LOC_642/Y 0.07fF
C56434 INVX1_LOC_27/A INVX1_LOC_19/A 0.10fF
C56435 INVX1_LOC_49/A NOR2X1_LOC_562/A 0.01fF
C56436 NOR2X1_LOC_160/B NOR2X1_LOC_634/A 0.02fF
C56437 NOR2X1_LOC_68/A NOR2X1_LOC_684/Y 0.09fF
C56438 NOR2X1_LOC_828/Y INVX1_LOC_15/A 0.26fF
C56439 NOR2X1_LOC_562/a_36_216# NOR2X1_LOC_357/Y 0.00fF
C56440 NOR2X1_LOC_816/A NOR2X1_LOC_88/Y 0.07fF
C56441 INVX1_LOC_209/Y VDD 0.48fF
C56442 NOR2X1_LOC_301/A NOR2X1_LOC_438/Y 0.00fF
C56443 NAND2X1_LOC_451/Y INVX1_LOC_91/A 0.01fF
C56444 NOR2X1_LOC_590/A INVX1_LOC_46/Y 0.04fF
C56445 INVX1_LOC_28/A INVX1_LOC_313/A 0.09fF
C56446 NOR2X1_LOC_299/Y NOR2X1_LOC_380/Y 0.09fF
C56447 INVX1_LOC_16/A INVX1_LOC_6/A 6.07fF
C56448 NOR2X1_LOC_457/B NOR2X1_LOC_331/B 0.87fF
C56449 NOR2X1_LOC_516/B INVX1_LOC_201/A 0.01fF
C56450 INVX1_LOC_48/A NOR2X1_LOC_121/A 0.01fF
C56451 NOR2X1_LOC_226/A INVX1_LOC_70/Y 0.14fF
C56452 NOR2X1_LOC_162/Y VDD 0.22fF
C56453 INVX1_LOC_135/A NOR2X1_LOC_322/Y 0.10fF
C56454 NAND2X1_LOC_725/B INVX1_LOC_240/Y 0.09fF
C56455 NOR2X1_LOC_761/Y NAND2X1_LOC_802/Y 0.17fF
C56456 NOR2X1_LOC_168/B NOR2X1_LOC_542/B 0.01fF
C56457 INVX1_LOC_73/A NOR2X1_LOC_123/B 0.09fF
C56458 NAND2X1_LOC_562/B NOR2X1_LOC_825/Y 0.19fF
C56459 INVX1_LOC_221/A INVX1_LOC_76/A 0.02fF
C56460 NAND2X1_LOC_722/A NOR2X1_LOC_164/Y 0.07fF
C56461 NOR2X1_LOC_215/A INVX1_LOC_109/Y 0.07fF
C56462 NAND2X1_LOC_354/B NOR2X1_LOC_682/Y 0.01fF
C56463 NOR2X1_LOC_816/A INVX1_LOC_84/A 4.60fF
C56464 NAND2X1_LOC_537/Y INVX1_LOC_49/Y 0.17fF
C56465 NOR2X1_LOC_612/a_36_216# INVX1_LOC_93/Y 0.01fF
C56466 NOR2X1_LOC_718/B VDD 0.02fF
C56467 INVX1_LOC_28/A NAND2X1_LOC_807/Y 0.19fF
C56468 INVX1_LOC_5/A INVX1_LOC_15/A 1.41fF
C56469 NOR2X1_LOC_168/B INVX1_LOC_143/Y 0.18fF
C56470 INVX1_LOC_8/A INVX1_LOC_12/Y 0.10fF
C56471 NOR2X1_LOC_433/A INVX1_LOC_38/A 0.18fF
C56472 NAND2X1_LOC_283/a_36_24# NOR2X1_LOC_536/A 0.00fF
C56473 NOR2X1_LOC_709/A NAND2X1_LOC_267/B 0.04fF
C56474 NAND2X1_LOC_722/A INVX1_LOC_46/A 0.07fF
C56475 NOR2X1_LOC_593/Y INVX1_LOC_38/A 0.07fF
C56476 NAND2X1_LOC_198/B NOR2X1_LOC_435/A 0.02fF
C56477 INVX1_LOC_72/Y NOR2X1_LOC_216/B 0.07fF
C56478 INVX1_LOC_178/A INVX1_LOC_15/A 0.24fF
C56479 NOR2X1_LOC_218/A INVX1_LOC_272/A 0.05fF
C56480 D_INPUT_4 NOR2X1_LOC_163/Y 0.01fF
C56481 NAND2X1_LOC_51/B NOR2X1_LOC_163/a_36_216# 0.00fF
C56482 INVX1_LOC_232/Y INVX1_LOC_178/Y 0.50fF
C56483 NOR2X1_LOC_112/Y INPUT_0 0.15fF
C56484 INVX1_LOC_13/A INVX1_LOC_74/Y 0.01fF
C56485 INVX1_LOC_276/A NAND2X1_LOC_687/A 0.01fF
C56486 NOR2X1_LOC_285/B INVX1_LOC_9/A 0.05fF
C56487 INVX1_LOC_24/A NOR2X1_LOC_197/B 0.01fF
C56488 NOR2X1_LOC_52/B NAND2X1_LOC_849/B 0.07fF
C56489 NOR2X1_LOC_596/A NAND2X1_LOC_435/a_36_24# 0.00fF
C56490 NOR2X1_LOC_510/Y NOR2X1_LOC_334/Y 0.51fF
C56491 INVX1_LOC_119/A NOR2X1_LOC_536/A 0.09fF
C56492 NOR2X1_LOC_309/Y NOR2X1_LOC_652/a_36_216# 0.00fF
C56493 NOR2X1_LOC_160/B INVX1_LOC_29/A 0.21fF
C56494 INVX1_LOC_218/A VDD -0.00fF
C56495 NAND2X1_LOC_205/A NAND2X1_LOC_205/a_36_24# 0.00fF
C56496 NOR2X1_LOC_52/B INVX1_LOC_38/A 0.53fF
C56497 NOR2X1_LOC_537/Y INVX1_LOC_117/A 0.07fF
C56498 INVX1_LOC_17/A NOR2X1_LOC_48/B 0.19fF
C56499 INVX1_LOC_41/A INVX1_LOC_274/A 0.10fF
C56500 NAND2X1_LOC_338/B INVX1_LOC_117/A 0.01fF
C56501 INVX1_LOC_35/A NOR2X1_LOC_383/B 0.06fF
C56502 INVX1_LOC_28/A INVX1_LOC_6/A 0.14fF
C56503 INVX1_LOC_186/A NOR2X1_LOC_174/B 0.06fF
C56504 NOR2X1_LOC_82/Y NOR2X1_LOC_266/B 0.39fF
C56505 INVX1_LOC_58/A NOR2X1_LOC_604/Y 0.04fF
C56506 NOR2X1_LOC_87/B INVX1_LOC_9/A 0.07fF
C56507 NAND2X1_LOC_323/B INVX1_LOC_117/A 0.03fF
C56508 INVX1_LOC_36/Y NAND2X1_LOC_41/Y 0.00fF
C56509 INVX1_LOC_34/A NOR2X1_LOC_78/Y 0.01fF
C56510 INVX1_LOC_276/A NAND2X1_LOC_846/a_36_24# 0.00fF
C56511 INVX1_LOC_12/Y NOR2X1_LOC_315/a_36_216# 0.08fF
C56512 INVX1_LOC_155/A NOR2X1_LOC_155/A 0.05fF
C56513 NOR2X1_LOC_802/A NOR2X1_LOC_729/A 0.24fF
C56514 INVX1_LOC_93/A INVX1_LOC_183/A 0.03fF
C56515 NAND2X1_LOC_198/B INVX1_LOC_63/A 0.10fF
C56516 INVX1_LOC_72/A INVX1_LOC_163/Y 0.16fF
C56517 NOR2X1_LOC_844/A NOR2X1_LOC_61/Y 0.01fF
C56518 NAND2X1_LOC_35/Y INVX1_LOC_57/A 0.07fF
C56519 NOR2X1_LOC_569/Y VDD 0.08fF
C56520 NAND2X1_LOC_734/B INVX1_LOC_185/A 0.01fF
C56521 NOR2X1_LOC_91/A NAND2X1_LOC_794/B 0.39fF
C56522 NOR2X1_LOC_15/Y NAND2X1_LOC_454/Y 0.07fF
C56523 INVX1_LOC_233/A NAND2X1_LOC_787/A 0.00fF
C56524 INVX1_LOC_27/A INVX1_LOC_26/Y 0.04fF
C56525 INVX1_LOC_49/A INVX1_LOC_285/A 0.07fF
C56526 NOR2X1_LOC_349/A INVX1_LOC_156/A 0.00fF
C56527 NOR2X1_LOC_78/A NOR2X1_LOC_564/Y 0.11fF
C56528 NOR2X1_LOC_361/B NOR2X1_LOC_334/Y 0.17fF
C56529 INVX1_LOC_90/A NOR2X1_LOC_601/Y 0.05fF
C56530 INVX1_LOC_154/Y NAND2X1_LOC_359/A 0.05fF
C56531 NOR2X1_LOC_357/Y NOR2X1_LOC_366/Y 0.05fF
C56532 INVX1_LOC_206/Y NOR2X1_LOC_74/A 0.01fF
C56533 D_INPUT_0 NAND2X1_LOC_650/B 0.07fF
C56534 INVX1_LOC_49/A NOR2X1_LOC_814/A 7.17fF
C56535 INVX1_LOC_224/A NAND2X1_LOC_223/A 0.03fF
C56536 INVX1_LOC_202/A NAND2X1_LOC_479/a_36_24# 0.00fF
C56537 NOR2X1_LOC_410/Y NAND2X1_LOC_291/B 0.04fF
C56538 NOR2X1_LOC_423/Y INVX1_LOC_179/A 0.28fF
C56539 INVX1_LOC_55/Y NAND2X1_LOC_447/Y 0.03fF
C56540 NOR2X1_LOC_91/A INVX1_LOC_48/Y 0.45fF
C56541 INVX1_LOC_108/Y INVX1_LOC_5/A 0.69fF
C56542 INVX1_LOC_249/A INVX1_LOC_19/A 0.00fF
C56543 INVX1_LOC_2/A NOR2X1_LOC_364/A 0.01fF
C56544 NAND2X1_LOC_662/Y NAND2X1_LOC_423/a_36_24# 0.01fF
C56545 NOR2X1_LOC_454/Y NOR2X1_LOC_654/A 0.04fF
C56546 NAND2X1_LOC_9/Y NOR2X1_LOC_791/Y 0.01fF
C56547 NOR2X1_LOC_100/A NAND2X1_LOC_85/Y 0.00fF
C56548 INVX1_LOC_143/A NOR2X1_LOC_197/B 0.05fF
C56549 NOR2X1_LOC_222/Y INVX1_LOC_179/A 0.03fF
C56550 NAND2X1_LOC_562/B INVX1_LOC_84/A 0.07fF
C56551 INVX1_LOC_50/A NAND2X1_LOC_725/B 0.01fF
C56552 NOR2X1_LOC_296/Y INVX1_LOC_23/Y 0.03fF
C56553 INVX1_LOC_72/A INVX1_LOC_3/Y 0.01fF
C56554 INVX1_LOC_48/Y INVX1_LOC_23/A 0.03fF
C56555 INVX1_LOC_315/Y INVX1_LOC_201/A 0.60fF
C56556 INVX1_LOC_16/A NOR2X1_LOC_79/A 0.01fF
C56557 INVX1_LOC_278/A INVX1_LOC_178/A 0.01fF
C56558 NOR2X1_LOC_78/B INVX1_LOC_113/A 0.08fF
C56559 NOR2X1_LOC_122/A INVX1_LOC_271/A 0.15fF
C56560 NOR2X1_LOC_773/Y NOR2X1_LOC_88/Y 0.08fF
C56561 NAND2X1_LOC_348/A INVX1_LOC_74/A 0.03fF
C56562 INVX1_LOC_293/A INVX1_LOC_16/Y 0.03fF
C56563 INVX1_LOC_2/A INVX1_LOC_285/A 0.08fF
C56564 NOR2X1_LOC_234/Y NOR2X1_LOC_662/A 0.20fF
C56565 INVX1_LOC_1/Y NOR2X1_LOC_743/Y 0.02fF
C56566 NOR2X1_LOC_636/B INVX1_LOC_262/A 0.03fF
C56567 NOR2X1_LOC_84/A NOR2X1_LOC_84/B 0.02fF
C56568 INVX1_LOC_35/A NOR2X1_LOC_463/a_36_216# 0.00fF
C56569 INVX1_LOC_89/A NOR2X1_LOC_536/A 0.70fF
C56570 INVX1_LOC_157/A NOR2X1_LOC_351/Y 0.09fF
C56571 INVX1_LOC_18/A INVX1_LOC_4/A 0.56fF
C56572 INVX1_LOC_2/A NOR2X1_LOC_814/A 0.10fF
C56573 INVX1_LOC_228/A NOR2X1_LOC_554/A 0.15fF
C56574 NOR2X1_LOC_457/a_36_216# NOR2X1_LOC_678/A 0.00fF
C56575 NOR2X1_LOC_226/A INVX1_LOC_285/A 0.10fF
C56576 NAND2X1_LOC_30/Y NAND2X1_LOC_40/a_36_24# 0.01fF
C56577 INVX1_LOC_33/A NOR2X1_LOC_89/A 0.31fF
C56578 NAND2X1_LOC_466/Y NAND2X1_LOC_74/B 0.03fF
C56579 INVX1_LOC_256/A NOR2X1_LOC_748/A 0.10fF
C56580 NOR2X1_LOC_742/A INVX1_LOC_37/A 0.07fF
C56581 INVX1_LOC_90/A NOR2X1_LOC_376/Y 0.06fF
C56582 INVX1_LOC_50/A NOR2X1_LOC_760/a_36_216# 0.00fF
C56583 NOR2X1_LOC_354/Y NOR2X1_LOC_324/A 0.00fF
C56584 NOR2X1_LOC_226/A NOR2X1_LOC_814/A 0.01fF
C56585 INVX1_LOC_89/A NAND2X1_LOC_659/a_36_24# 0.00fF
C56586 NOR2X1_LOC_773/Y INVX1_LOC_84/A 0.08fF
C56587 NOR2X1_LOC_589/A NAND2X1_LOC_210/a_36_24# 0.00fF
C56588 INVX1_LOC_246/A INVX1_LOC_23/A 0.08fF
C56589 NOR2X1_LOC_92/Y INVX1_LOC_306/Y 0.03fF
C56590 INVX1_LOC_10/A NAND2X1_LOC_792/a_36_24# 0.01fF
C56591 NOR2X1_LOC_391/A INVX1_LOC_123/Y 0.01fF
C56592 INVX1_LOC_33/A NOR2X1_LOC_170/A 0.01fF
C56593 NOR2X1_LOC_160/B NOR2X1_LOC_843/a_36_216# 0.00fF
C56594 INVX1_LOC_64/A NAND2X1_LOC_799/A 0.03fF
C56595 INVX1_LOC_89/A NAND2X1_LOC_93/B 0.07fF
C56596 NAND2X1_LOC_200/B INVX1_LOC_19/A 0.74fF
C56597 INVX1_LOC_53/Y INVX1_LOC_63/A 0.10fF
C56598 INVX1_LOC_58/A NOR2X1_LOC_361/a_36_216# 0.00fF
C56599 INVX1_LOC_73/A NOR2X1_LOC_331/B 0.04fF
C56600 INVX1_LOC_292/A NOR2X1_LOC_717/A 0.37fF
C56601 NAND2X1_LOC_350/B INVX1_LOC_29/A 0.52fF
C56602 INVX1_LOC_232/Y INVX1_LOC_12/A 1.20fF
C56603 NOR2X1_LOC_87/B NOR2X1_LOC_861/Y 0.06fF
C56604 INVX1_LOC_196/Y NOR2X1_LOC_676/Y 0.05fF
C56605 INVX1_LOC_89/A NAND2X1_LOC_425/Y 0.13fF
C56606 NOR2X1_LOC_846/Y NOR2X1_LOC_848/Y 0.13fF
C56607 NAND2X1_LOC_562/B INVX1_LOC_15/A 0.00fF
C56608 INVX1_LOC_208/A INVX1_LOC_29/A 0.01fF
C56609 NAND2X1_LOC_53/Y INVX1_LOC_50/Y 0.01fF
C56610 INVX1_LOC_58/A INVX1_LOC_72/A 0.26fF
C56611 NOR2X1_LOC_516/B INVX1_LOC_29/A 0.06fF
C56612 NOR2X1_LOC_332/A INVX1_LOC_84/A 0.08fF
C56613 INVX1_LOC_298/A INVX1_LOC_174/A 0.01fF
C56614 NOR2X1_LOC_337/Y NAND2X1_LOC_472/Y 0.03fF
C56615 INVX1_LOC_40/A NOR2X1_LOC_89/A 0.19fF
C56616 NAND2X1_LOC_9/Y INVX1_LOC_30/A 0.16fF
C56617 NAND2X1_LOC_323/a_36_24# NOR2X1_LOC_809/B 0.01fF
C56618 NAND2X1_LOC_726/Y NOR2X1_LOC_89/A 0.07fF
C56619 INVX1_LOC_89/A NOR2X1_LOC_649/B 0.32fF
C56620 NOR2X1_LOC_473/B NOR2X1_LOC_473/a_36_216# 0.01fF
C56621 NOR2X1_LOC_757/Y INVX1_LOC_290/Y 0.06fF
C56622 INVX1_LOC_233/A INVX1_LOC_30/A 0.18fF
C56623 INVX1_LOC_27/A INVX1_LOC_161/Y 0.07fF
C56624 INVX1_LOC_89/A INVX1_LOC_3/A 0.54fF
C56625 NOR2X1_LOC_350/A NOR2X1_LOC_668/Y 0.10fF
C56626 NOR2X1_LOC_91/A NOR2X1_LOC_189/A 0.01fF
C56627 INVX1_LOC_234/A INVX1_LOC_19/A 0.42fF
C56628 NOR2X1_LOC_298/Y INVX1_LOC_240/Y 0.21fF
C56629 INVX1_LOC_94/A INVX1_LOC_57/A 0.54fF
C56630 INVX1_LOC_64/A NOR2X1_LOC_532/a_36_216# 0.01fF
C56631 NAND2X1_LOC_338/B INVX1_LOC_3/Y 0.16fF
C56632 NOR2X1_LOC_605/B NOR2X1_LOC_89/A 0.07fF
C56633 INPUT_1 INVX1_LOC_265/Y 0.01fF
C56634 INVX1_LOC_140/A NOR2X1_LOC_88/Y 0.17fF
C56635 INVX1_LOC_174/A D_INPUT_6 0.08fF
C56636 INVX1_LOC_28/A NOR2X1_LOC_117/Y 0.02fF
C56637 NOR2X1_LOC_709/A INVX1_LOC_4/Y 0.19fF
C56638 NOR2X1_LOC_75/Y NOR2X1_LOC_454/Y 0.10fF
C56639 NOR2X1_LOC_437/Y INVX1_LOC_271/A 0.61fF
C56640 D_GATE_579 INVX1_LOC_42/A 0.00fF
C56641 NOR2X1_LOC_593/Y NAND2X1_LOC_256/a_36_24# 0.01fF
C56642 INVX1_LOC_132/A NOR2X1_LOC_443/Y 0.04fF
C56643 INVX1_LOC_64/A INVX1_LOC_18/A 4.43fF
C56644 NOR2X1_LOC_773/Y INVX1_LOC_15/A 0.07fF
C56645 INVX1_LOC_311/A NOR2X1_LOC_433/Y 0.31fF
C56646 INVX1_LOC_177/A NOR2X1_LOC_334/Y 0.04fF
C56647 NAND2X1_LOC_728/Y INVX1_LOC_64/A 0.12fF
C56648 NOR2X1_LOC_602/A NOR2X1_LOC_186/Y 0.02fF
C56649 NAND2X1_LOC_477/A NAND2X1_LOC_477/a_36_24# 0.01fF
C56650 INVX1_LOC_225/A NOR2X1_LOC_282/Y 0.01fF
C56651 NOR2X1_LOC_798/A INVX1_LOC_30/A 0.06fF
C56652 NOR2X1_LOC_596/A NOR2X1_LOC_678/A 0.03fF
C56653 INVX1_LOC_286/A NOR2X1_LOC_118/a_36_216# 0.00fF
C56654 INVX1_LOC_232/A INVX1_LOC_32/A 0.00fF
C56655 NOR2X1_LOC_596/A INVX1_LOC_295/Y 0.00fF
C56656 INVX1_LOC_140/A INVX1_LOC_84/A 0.40fF
C56657 INVX1_LOC_48/Y INVX1_LOC_31/A 0.08fF
C56658 NOR2X1_LOC_601/Y INVX1_LOC_38/A 0.18fF
C56659 INVX1_LOC_5/A NOR2X1_LOC_168/Y 0.06fF
C56660 NOR2X1_LOC_744/Y NOR2X1_LOC_109/Y 0.03fF
C56661 INVX1_LOC_77/A INVX1_LOC_58/Y 0.04fF
C56662 INVX1_LOC_64/A NOR2X1_LOC_637/Y 0.15fF
C56663 NOR2X1_LOC_772/A INVX1_LOC_19/A 0.01fF
C56664 INVX1_LOC_17/A NAND2X1_LOC_350/A 0.04fF
C56665 NOR2X1_LOC_602/A NAND2X1_LOC_573/Y 0.03fF
C56666 NAND2X1_LOC_721/A INVX1_LOC_37/A 0.03fF
C56667 NOR2X1_LOC_413/a_36_216# INVX1_LOC_23/A 0.00fF
C56668 NAND2X1_LOC_149/Y INVX1_LOC_36/A 0.13fF
C56669 NAND2X1_LOC_778/Y NOR2X1_LOC_68/A 0.02fF
C56670 NOR2X1_LOC_19/B INVX1_LOC_19/A 0.06fF
C56671 VDD NAND2X1_LOC_472/Y 0.00fF
C56672 INVX1_LOC_64/A INVX1_LOC_172/A 0.00fF
C56673 INVX1_LOC_34/A NAND2X1_LOC_860/A 0.03fF
C56674 NAND2X1_LOC_231/Y NAND2X1_LOC_286/B 0.01fF
C56675 NAND2X1_LOC_650/B NAND2X1_LOC_848/A 0.10fF
C56676 INVX1_LOC_116/A INVX1_LOC_13/Y 0.01fF
C56677 NOR2X1_LOC_40/a_36_216# INVX1_LOC_38/A 0.01fF
C56678 NOR2X1_LOC_405/A INVX1_LOC_291/A 0.56fF
C56679 NOR2X1_LOC_315/Y NAND2X1_LOC_205/A 0.05fF
C56680 INVX1_LOC_90/A NAND2X1_LOC_254/Y 0.03fF
C56681 NOR2X1_LOC_629/a_36_216# INVX1_LOC_23/A 0.00fF
C56682 INVX1_LOC_17/A NOR2X1_LOC_441/Y 0.02fF
C56683 NOR2X1_LOC_533/Y INVX1_LOC_141/Y 0.02fF
C56684 NOR2X1_LOC_220/B NOR2X1_LOC_303/Y 0.02fF
C56685 NAND2X1_LOC_200/B INVX1_LOC_26/Y 0.03fF
C56686 INVX1_LOC_298/Y INVX1_LOC_208/A 0.01fF
C56687 NOR2X1_LOC_332/A INVX1_LOC_15/A 0.14fF
C56688 INVX1_LOC_139/Y INVX1_LOC_281/Y 0.01fF
C56689 NOR2X1_LOC_658/Y INVX1_LOC_103/A 0.10fF
C56690 INVX1_LOC_136/A NAND2X1_LOC_303/Y 0.10fF
C56691 NOR2X1_LOC_577/Y NOR2X1_LOC_674/a_36_216# 0.01fF
C56692 NOR2X1_LOC_312/a_36_216# INVX1_LOC_57/A 0.00fF
C56693 NOR2X1_LOC_84/Y INVX1_LOC_23/A 0.27fF
C56694 NOR2X1_LOC_56/Y NAND2X1_LOC_434/Y 0.02fF
C56695 NOR2X1_LOC_569/a_36_216# INVX1_LOC_99/A 0.02fF
C56696 NOR2X1_LOC_15/Y NOR2X1_LOC_68/A 0.02fF
C56697 INVX1_LOC_246/A INVX1_LOC_31/A 0.00fF
C56698 INVX1_LOC_216/A INVX1_LOC_23/A 0.03fF
C56699 INVX1_LOC_305/Y NOR2X1_LOC_383/B 0.14fF
C56700 VDD NAND2X1_LOC_637/Y 0.20fF
C56701 INVX1_LOC_233/A NAND2X1_LOC_722/A 0.93fF
C56702 INVX1_LOC_284/Y NAND2X1_LOC_733/Y 0.03fF
C56703 INVX1_LOC_11/A NAND2X1_LOC_386/a_36_24# 0.00fF
C56704 NAND2X1_LOC_734/a_36_24# NOR2X1_LOC_406/A 0.00fF
C56705 NAND2X1_LOC_348/A NAND2X1_LOC_254/Y 0.06fF
C56706 NAND2X1_LOC_550/A NAND2X1_LOC_634/Y 0.10fF
C56707 INVX1_LOC_16/A INVX1_LOC_270/A 0.17fF
C56708 NOR2X1_LOC_274/Y INVX1_LOC_1/A 0.02fF
C56709 NAND2X1_LOC_57/a_36_24# NOR2X1_LOC_160/B 0.00fF
C56710 INVX1_LOC_38/A NOR2X1_LOC_376/Y 0.01fF
C56711 INVX1_LOC_89/A NAND2X1_LOC_470/B 0.03fF
C56712 NOR2X1_LOC_810/A NOR2X1_LOC_798/Y 0.01fF
C56713 INVX1_LOC_103/A NOR2X1_LOC_13/Y 0.10fF
C56714 NAND2X1_LOC_349/B INVX1_LOC_270/Y 0.01fF
C56715 NOR2X1_LOC_858/B INVX1_LOC_307/A 0.04fF
C56716 NAND2X1_LOC_477/A INVX1_LOC_306/Y 0.03fF
C56717 NOR2X1_LOC_335/B INVX1_LOC_42/A 0.03fF
C56718 NOR2X1_LOC_220/A NOR2X1_LOC_678/A 0.03fF
C56719 NOR2X1_LOC_209/Y INVX1_LOC_213/A 0.07fF
C56720 INVX1_LOC_278/A NOR2X1_LOC_773/Y 0.01fF
C56721 INVX1_LOC_176/A NAND2X1_LOC_85/Y 0.09fF
C56722 INVX1_LOC_113/A INVX1_LOC_46/A 0.04fF
C56723 INVX1_LOC_290/A INVX1_LOC_23/A 1.28fF
C56724 NOR2X1_LOC_626/Y NOR2X1_LOC_593/a_36_216# 0.00fF
C56725 NOR2X1_LOC_220/B INVX1_LOC_54/Y 0.01fF
C56726 INVX1_LOC_284/Y INVX1_LOC_217/A 0.11fF
C56727 NOR2X1_LOC_71/Y NAND2X1_LOC_99/A 0.21fF
C56728 NAND2X1_LOC_724/Y INVX1_LOC_229/Y 0.04fF
C56729 INVX1_LOC_55/A NOR2X1_LOC_596/A 0.07fF
C56730 INVX1_LOC_225/Y NOR2X1_LOC_303/Y 0.10fF
C56731 NOR2X1_LOC_75/Y INVX1_LOC_77/A 0.03fF
C56732 INVX1_LOC_34/A NAND2X1_LOC_537/Y 0.19fF
C56733 NOR2X1_LOC_140/A INVX1_LOC_82/A 0.01fF
C56734 NOR2X1_LOC_577/a_36_216# INVX1_LOC_53/A 0.01fF
C56735 NAND2X1_LOC_624/B INVX1_LOC_22/A 0.00fF
C56736 NAND2X1_LOC_53/Y NOR2X1_LOC_718/Y 0.03fF
C56737 INVX1_LOC_11/A INVX1_LOC_33/A 1.82fF
C56738 INVX1_LOC_307/Y NOR2X1_LOC_729/A 0.06fF
C56739 NOR2X1_LOC_211/Y INVX1_LOC_22/A 0.03fF
C56740 INVX1_LOC_286/Y INVX1_LOC_24/A 0.10fF
C56741 INVX1_LOC_17/A NOR2X1_LOC_142/Y 0.01fF
C56742 VDD NAND2X1_LOC_206/Y 0.86fF
C56743 NOR2X1_LOC_500/Y INVX1_LOC_50/Y 0.03fF
C56744 INVX1_LOC_226/Y INVX1_LOC_50/Y 0.03fF
C56745 NOR2X1_LOC_590/A INVX1_LOC_49/A 1.56fF
C56746 INVX1_LOC_36/A NOR2X1_LOC_744/Y 0.01fF
C56747 INVX1_LOC_108/Y NOR2X1_LOC_332/A 0.01fF
C56748 VDD NAND2X1_LOC_773/B 1.28fF
C56749 INVX1_LOC_58/A INVX1_LOC_313/Y 0.10fF
C56750 INVX1_LOC_285/Y NOR2X1_LOC_334/Y 0.10fF
C56751 INVX1_LOC_28/A INVX1_LOC_270/A 0.17fF
C56752 NOR2X1_LOC_160/B INVX1_LOC_8/A 0.19fF
C56753 NOR2X1_LOC_818/a_36_216# NOR2X1_LOC_332/A 0.00fF
C56754 NOR2X1_LOC_387/A NOR2X1_LOC_409/B 0.00fF
C56755 NAND2X1_LOC_211/Y INVX1_LOC_29/A 0.07fF
C56756 NOR2X1_LOC_620/Y INVX1_LOC_45/A 0.01fF
C56757 INVX1_LOC_22/A NOR2X1_LOC_440/B 0.18fF
C56758 NOR2X1_LOC_68/A NOR2X1_LOC_860/B 0.15fF
C56759 INVX1_LOC_17/A NOR2X1_LOC_655/B 0.10fF
C56760 NAND2X1_LOC_361/Y NOR2X1_LOC_500/B 0.10fF
C56761 INVX1_LOC_256/A NOR2X1_LOC_493/B 0.12fF
C56762 INVX1_LOC_266/A NOR2X1_LOC_500/Y 0.01fF
C56763 NOR2X1_LOC_590/A INVX1_LOC_60/A 0.01fF
C56764 INVX1_LOC_232/Y INVX1_LOC_228/Y 0.10fF
C56765 INVX1_LOC_2/A NAND2X1_LOC_803/B 0.05fF
C56766 INVX1_LOC_118/A INVX1_LOC_285/A 0.09fF
C56767 INPUT_0 NAND2X1_LOC_286/B 0.06fF
C56768 INVX1_LOC_54/Y INVX1_LOC_225/Y 0.07fF
C56769 NOR2X1_LOC_201/a_36_216# NAND2X1_LOC_116/A 0.00fF
C56770 INVX1_LOC_75/A INVX1_LOC_270/Y 0.02fF
C56771 NAND2X1_LOC_181/Y NOR2X1_LOC_103/Y 0.01fF
C56772 NOR2X1_LOC_226/A NAND2X1_LOC_803/B 0.02fF
C56773 INVX1_LOC_124/Y INVX1_LOC_104/A 0.01fF
C56774 NOR2X1_LOC_482/a_36_216# INVX1_LOC_42/A 0.00fF
C56775 INVX1_LOC_136/A NOR2X1_LOC_690/A 0.15fF
C56776 INVX1_LOC_2/A NOR2X1_LOC_590/A 0.09fF
C56777 INVX1_LOC_278/A INVX1_LOC_140/A 0.07fF
C56778 INVX1_LOC_65/A NOR2X1_LOC_334/Y 0.10fF
C56779 NAND2X1_LOC_194/a_36_24# NOR2X1_LOC_103/Y 0.00fF
C56780 INVX1_LOC_28/A NOR2X1_LOC_109/Y 0.07fF
C56781 INVX1_LOC_286/A INVX1_LOC_181/A 0.23fF
C56782 INVX1_LOC_27/A INVX1_LOC_62/A 0.11fF
C56783 INVX1_LOC_24/A INVX1_LOC_283/Y -0.01fF
C56784 NAND2X1_LOC_796/B NOR2X1_LOC_246/A 0.03fF
C56785 INVX1_LOC_31/A INVX1_LOC_216/A 0.06fF
C56786 INVX1_LOC_26/A INVX1_LOC_91/A 0.04fF
C56787 NOR2X1_LOC_226/A NOR2X1_LOC_590/A 0.00fF
C56788 INVX1_LOC_24/A NAND2X1_LOC_486/a_36_24# 0.00fF
C56789 INVX1_LOC_69/Y NOR2X1_LOC_748/A 0.10fF
C56790 NAND2X1_LOC_311/a_36_24# NOR2X1_LOC_802/A 0.00fF
C56791 INVX1_LOC_11/A NOR2X1_LOC_605/B 0.04fF
C56792 NOR2X1_LOC_334/Y NOR2X1_LOC_137/B 0.01fF
C56793 NOR2X1_LOC_753/a_36_216# NOR2X1_LOC_753/Y 0.00fF
C56794 NOR2X1_LOC_537/A INVX1_LOC_77/A 0.01fF
C56795 NAND2X1_LOC_860/A INPUT_0 0.18fF
C56796 INVX1_LOC_64/A INVX1_LOC_31/Y 0.05fF
C56797 NOR2X1_LOC_635/A NOR2X1_LOC_68/A 0.00fF
C56798 NOR2X1_LOC_791/Y NAND2X1_LOC_842/B 0.16fF
C56799 NOR2X1_LOC_716/B INVX1_LOC_77/A 0.07fF
C56800 NOR2X1_LOC_598/B INVX1_LOC_86/A 0.07fF
C56801 VDD NOR2X1_LOC_393/Y 0.12fF
C56802 INVX1_LOC_36/A NAND2X1_LOC_717/Y 0.03fF
C56803 NOR2X1_LOC_589/A NAND2X1_LOC_793/Y 0.37fF
C56804 NAND2X1_LOC_794/B NAND2X1_LOC_807/Y 0.07fF
C56805 NOR2X1_LOC_168/B NAND2X1_LOC_497/a_36_24# 0.00fF
C56806 INVX1_LOC_33/A NOR2X1_LOC_433/A 0.19fF
C56807 INVX1_LOC_45/A NAND2X1_LOC_181/Y 0.03fF
C56808 NOR2X1_LOC_78/A NOR2X1_LOC_646/B 0.02fF
C56809 NOR2X1_LOC_496/Y NOR2X1_LOC_497/Y 0.17fF
C56810 NOR2X1_LOC_392/B INVX1_LOC_314/Y 0.10fF
C56811 INVX1_LOC_50/A NOR2X1_LOC_139/Y 0.01fF
C56812 NAND2X1_LOC_564/B NAND2X1_LOC_543/a_36_24# 0.01fF
C56813 INVX1_LOC_33/A NOR2X1_LOC_593/Y 6.72fF
C56814 INVX1_LOC_50/A NAND2X1_LOC_655/A 0.00fF
C56815 INVX1_LOC_17/A NOR2X1_LOC_99/B 0.06fF
C56816 INVX1_LOC_95/A INVX1_LOC_181/A 0.00fF
C56817 NOR2X1_LOC_216/B INVX1_LOC_19/A 0.01fF
C56818 NAND2X1_LOC_30/Y NOR2X1_LOC_763/Y 0.01fF
C56819 NOR2X1_LOC_338/a_36_216# INVX1_LOC_76/A 0.01fF
C56820 INVX1_LOC_18/A NAND2X1_LOC_850/Y 0.07fF
C56821 INVX1_LOC_78/A NOR2X1_LOC_482/a_36_216# 0.00fF
C56822 INVX1_LOC_255/Y NAND2X1_LOC_577/A 0.09fF
C56823 INVX1_LOC_24/Y NOR2X1_LOC_356/A 0.09fF
C56824 INVX1_LOC_188/A INVX1_LOC_279/A -0.01fF
C56825 INVX1_LOC_17/A NOR2X1_LOC_846/B 0.04fF
C56826 INVX1_LOC_36/A INVX1_LOC_16/A 0.10fF
C56827 NAND2X1_LOC_722/A NAND2X1_LOC_866/A 0.02fF
C56828 INVX1_LOC_21/A NOR2X1_LOC_196/Y 0.03fF
C56829 NOR2X1_LOC_752/a_36_216# INVX1_LOC_72/A 0.00fF
C56830 INVX1_LOC_50/A NAND2X1_LOC_468/B 0.14fF
C56831 NAND2X1_LOC_341/A NOR2X1_LOC_52/Y 0.04fF
C56832 INVX1_LOC_256/A INVX1_LOC_89/A 0.08fF
C56833 NOR2X1_LOC_15/Y NAND2X1_LOC_462/a_36_24# 0.00fF
C56834 NOR2X1_LOC_718/B INVX1_LOC_153/Y 0.07fF
C56835 INVX1_LOC_33/A NOR2X1_LOC_52/B 0.15fF
C56836 NOR2X1_LOC_67/Y INVX1_LOC_46/Y 0.20fF
C56837 NOR2X1_LOC_479/a_36_216# NOR2X1_LOC_375/Y 0.00fF
C56838 INVX1_LOC_21/A NOR2X1_LOC_775/a_36_216# 0.00fF
C56839 INVX1_LOC_5/A INVX1_LOC_123/A 0.01fF
C56840 VDD NOR2X1_LOC_639/Y 0.24fF
C56841 NAND2X1_LOC_724/Y INVX1_LOC_20/A 0.03fF
C56842 INVX1_LOC_64/A NOR2X1_LOC_43/a_36_216# 0.01fF
C56843 NOR2X1_LOC_589/A NAND2X1_LOC_16/Y 0.03fF
C56844 NAND2X1_LOC_733/Y NOR2X1_LOC_525/Y 0.01fF
C56845 NAND2X1_LOC_477/Y INVX1_LOC_19/A 0.05fF
C56846 NAND2X1_LOC_733/Y NAND2X1_LOC_809/A 0.01fF
C56847 INVX1_LOC_286/Y NAND2X1_LOC_800/Y 0.03fF
C56848 NOR2X1_LOC_248/Y INVX1_LOC_10/A 0.02fF
C56849 NOR2X1_LOC_88/Y INVX1_LOC_42/A 0.10fF
C56850 NOR2X1_LOC_92/Y NOR2X1_LOC_74/A 0.07fF
C56851 NAND2X1_LOC_574/A NOR2X1_LOC_33/B 0.06fF
C56852 NOR2X1_LOC_718/B INVX1_LOC_121/Y 0.00fF
C56853 NOR2X1_LOC_35/Y NOR2X1_LOC_416/A 0.10fF
C56854 NAND2X1_LOC_63/Y NOR2X1_LOC_814/A 0.00fF
C56855 NOR2X1_LOC_433/A NAND2X1_LOC_798/A 0.00fF
C56856 NAND2X1_LOC_363/B NOR2X1_LOC_545/B 0.06fF
C56857 NOR2X1_LOC_476/Y NOR2X1_LOC_459/A 0.01fF
C56858 INVX1_LOC_228/A NOR2X1_LOC_516/B 0.01fF
C56859 INVX1_LOC_2/A NAND2X1_LOC_354/B 0.03fF
C56860 INVX1_LOC_255/Y NAND2X1_LOC_656/A 0.11fF
C56861 NOR2X1_LOC_606/Y INVX1_LOC_89/A 0.00fF
C56862 INVX1_LOC_207/A NAND2X1_LOC_374/Y 0.05fF
C56863 INVX1_LOC_226/Y NOR2X1_LOC_559/B 0.00fF
C56864 NOR2X1_LOC_208/Y INVX1_LOC_16/A 0.58fF
C56865 D_INPUT_3 NOR2X1_LOC_414/Y 0.02fF
C56866 NOR2X1_LOC_558/A INVX1_LOC_29/Y 0.00fF
C56867 NOR2X1_LOC_617/Y INVX1_LOC_22/A 0.00fF
C56868 NOR2X1_LOC_220/A NAND2X1_LOC_536/a_36_24# 0.00fF
C56869 INVX1_LOC_94/Y INVX1_LOC_54/A 0.12fF
C56870 NOR2X1_LOC_226/A NAND2X1_LOC_354/B 0.15fF
C56871 NOR2X1_LOC_778/B NOR2X1_LOC_147/B 0.00fF
C56872 INVX1_LOC_90/A NAND2X1_LOC_185/a_36_24# 0.00fF
C56873 NAND2X1_LOC_724/Y NOR2X1_LOC_765/Y 0.08fF
C56874 INVX1_LOC_224/Y INVX1_LOC_117/A 0.02fF
C56875 NOR2X1_LOC_48/B NOR2X1_LOC_430/Y 0.37fF
C56876 INVX1_LOC_84/A INVX1_LOC_42/A 0.20fF
C56877 NOR2X1_LOC_361/Y INVX1_LOC_133/Y 0.03fF
C56878 INVX1_LOC_188/A INVX1_LOC_182/Y 0.02fF
C56879 NOR2X1_LOC_75/Y NAND2X1_LOC_832/Y 0.01fF
C56880 INVX1_LOC_36/A INVX1_LOC_28/A 0.32fF
C56881 NAND2X1_LOC_207/B INVX1_LOC_29/A 0.03fF
C56882 INVX1_LOC_72/A NOR2X1_LOC_533/a_36_216# 0.15fF
C56883 INVX1_LOC_226/Y NOR2X1_LOC_6/B 0.09fF
C56884 INVX1_LOC_54/A INVX1_LOC_181/A 0.40fF
C56885 NOR2X1_LOC_88/Y INVX1_LOC_78/A 0.06fF
C56886 NOR2X1_LOC_717/B INVX1_LOC_77/A 0.03fF
C56887 NAND2X1_LOC_56/a_36_24# INVX1_LOC_311/A 0.00fF
C56888 NOR2X1_LOC_729/A NOR2X1_LOC_809/A 0.00fF
C56889 NOR2X1_LOC_309/Y INVX1_LOC_16/A 0.03fF
C56890 NAND2X1_LOC_347/B NAND2X1_LOC_642/Y 0.24fF
C56891 NOR2X1_LOC_763/Y INVX1_LOC_49/A 0.36fF
C56892 INVX1_LOC_2/A NOR2X1_LOC_488/Y 0.06fF
C56893 INVX1_LOC_290/A NOR2X1_LOC_75/a_36_216# 0.01fF
C56894 NAND2X1_LOC_538/Y NOR2X1_LOC_595/Y 0.20fF
C56895 NAND2X1_LOC_773/Y INVX1_LOC_95/Y 0.10fF
C56896 INVX1_LOC_90/A INVX1_LOC_314/Y 1.19fF
C56897 NOR2X1_LOC_638/Y INVX1_LOC_92/A 0.02fF
C56898 INVX1_LOC_135/A NAND2X1_LOC_833/Y 0.14fF
C56899 INVX1_LOC_58/Y INVX1_LOC_9/A 0.07fF
C56900 INVX1_LOC_145/A INVX1_LOC_28/A 0.03fF
C56901 NOR2X1_LOC_538/Y INVX1_LOC_22/A 0.01fF
C56902 NOR2X1_LOC_226/A NOR2X1_LOC_488/Y 0.04fF
C56903 INVX1_LOC_78/A INVX1_LOC_84/A 0.17fF
C56904 NOR2X1_LOC_208/Y INVX1_LOC_28/A 0.08fF
C56905 NOR2X1_LOC_569/Y INVX1_LOC_177/A 0.01fF
C56906 NAND2X1_LOC_326/A INVX1_LOC_76/A 0.77fF
C56907 NOR2X1_LOC_226/A NOR2X1_LOC_82/Y 0.18fF
C56908 INVX1_LOC_290/A INVX1_LOC_191/Y 2.38fF
C56909 INVX1_LOC_7/A NOR2X1_LOC_87/B 0.13fF
C56910 NOR2X1_LOC_167/a_36_216# INVX1_LOC_119/Y 0.03fF
C56911 NOR2X1_LOC_155/A INVX1_LOC_57/A 0.00fF
C56912 INVX1_LOC_11/A NOR2X1_LOC_486/Y 0.03fF
C56913 INVX1_LOC_141/A INVX1_LOC_91/A 0.06fF
C56914 INVX1_LOC_21/A INVX1_LOC_33/Y 0.08fF
C56915 NOR2X1_LOC_373/Y NOR2X1_LOC_315/Y 0.48fF
C56916 NAND2X1_LOC_354/B NAND2X1_LOC_648/A 0.00fF
C56917 INVX1_LOC_2/A INVX1_LOC_227/A 0.07fF
C56918 INVX1_LOC_53/A INVX1_LOC_180/Y 0.01fF
C56919 INVX1_LOC_49/A NOR2X1_LOC_703/A 0.04fF
C56920 INVX1_LOC_41/A NOR2X1_LOC_356/A 0.07fF
C56921 INVX1_LOC_271/A NOR2X1_LOC_841/A 0.01fF
C56922 INVX1_LOC_24/A NOR2X1_LOC_721/Y 0.01fF
C56923 INVX1_LOC_15/A INVX1_LOC_42/A 0.07fF
C56924 INVX1_LOC_124/A NAND2X1_LOC_656/a_36_24# 0.00fF
C56925 NOR2X1_LOC_65/B INVX1_LOC_84/A 0.03fF
C56926 NOR2X1_LOC_151/Y INVX1_LOC_77/A 0.07fF
C56927 INVX1_LOC_1/Y INVX1_LOC_53/Y 0.03fF
C56928 INVX1_LOC_313/Y NOR2X1_LOC_344/a_36_216# 0.00fF
C56929 NOR2X1_LOC_756/a_36_216# INVX1_LOC_8/A 0.01fF
C56930 NAND2X1_LOC_21/Y INVX1_LOC_140/A 0.35fF
C56931 NOR2X1_LOC_334/Y NOR2X1_LOC_830/Y 0.03fF
C56932 NAND2X1_LOC_793/Y INVX1_LOC_20/A 0.01fF
C56933 INVX1_LOC_50/A NOR2X1_LOC_66/Y 0.01fF
C56934 INVX1_LOC_256/A NOR2X1_LOC_52/a_36_216# 0.00fF
C56935 D_INPUT_1 INVX1_LOC_27/Y 0.01fF
C56936 NAND2X1_LOC_402/B INVX1_LOC_163/Y 0.17fF
C56937 NOR2X1_LOC_778/B INVX1_LOC_97/A 0.02fF
C56938 NAND2X1_LOC_181/Y NOR2X1_LOC_123/B 0.00fF
C56939 NOR2X1_LOC_644/Y INVX1_LOC_55/Y 0.05fF
C56940 NAND2X1_LOC_787/A INVX1_LOC_119/Y 0.03fF
C56941 NAND2X1_LOC_198/B NOR2X1_LOC_318/B 0.03fF
C56942 NOR2X1_LOC_48/B INVX1_LOC_94/Y 0.07fF
C56943 INVX1_LOC_78/A NAND2X1_LOC_220/B 0.27fF
C56944 INVX1_LOC_41/A NOR2X1_LOC_74/A 0.05fF
C56945 NOR2X1_LOC_778/B INVX1_LOC_90/A 0.03fF
C56946 NOR2X1_LOC_103/Y INVX1_LOC_117/A 0.16fF
C56947 INVX1_LOC_50/Y INVX1_LOC_307/A 0.07fF
C56948 INVX1_LOC_208/A NAND2X1_LOC_140/A 0.03fF
C56949 NOR2X1_LOC_392/Y INVX1_LOC_3/A 0.14fF
C56950 NOR2X1_LOC_717/B NOR2X1_LOC_687/Y 0.03fF
C56951 INVX1_LOC_181/Y NOR2X1_LOC_192/A 0.03fF
C56952 INVX1_LOC_36/A NOR2X1_LOC_35/Y 0.01fF
C56953 INVX1_LOC_50/Y NOR2X1_LOC_445/B 0.07fF
C56954 INPUT_0 NOR2X1_LOC_516/Y 0.01fF
C56955 NAND2X1_LOC_198/B INVX1_LOC_93/Y 0.01fF
C56956 INVX1_LOC_41/A NOR2X1_LOC_9/Y 0.10fF
C56957 INVX1_LOC_78/A INVX1_LOC_15/A 9.84fF
C56958 INVX1_LOC_40/Y D_INPUT_3 0.00fF
C56959 NOR2X1_LOC_307/B INVX1_LOC_311/Y 0.03fF
C56960 NOR2X1_LOC_152/Y INVX1_LOC_264/Y 0.02fF
C56961 NAND2X1_LOC_477/A NOR2X1_LOC_74/A 0.10fF
C56962 NOR2X1_LOC_82/Y INPUT_1 0.99fF
C56963 NOR2X1_LOC_828/A NOR2X1_LOC_687/Y 0.03fF
C56964 INVX1_LOC_23/A INVX1_LOC_261/Y 0.07fF
C56965 INVX1_LOC_135/A NOR2X1_LOC_719/B 0.05fF
C56966 NOR2X1_LOC_448/B NAND2X1_LOC_93/B 0.03fF
C56967 NAND2X1_LOC_803/B INVX1_LOC_118/A 0.00fF
C56968 NOR2X1_LOC_48/B INVX1_LOC_296/A 0.06fF
C56969 INVX1_LOC_45/A INVX1_LOC_117/A 0.21fF
C56970 NOR2X1_LOC_615/Y INVX1_LOC_118/A 0.01fF
C56971 NOR2X1_LOC_721/Y INVX1_LOC_143/A 0.02fF
C56972 INVX1_LOC_103/Y INVX1_LOC_91/A 0.01fF
C56973 INVX1_LOC_266/A NOR2X1_LOC_445/B 0.10fF
C56974 NOR2X1_LOC_666/Y NOR2X1_LOC_155/A 0.13fF
C56975 NOR2X1_LOC_312/Y NAND2X1_LOC_808/A 0.01fF
C56976 NOR2X1_LOC_647/A INVX1_LOC_4/A 0.10fF
C56977 NOR2X1_LOC_415/A INVX1_LOC_89/A 0.02fF
C56978 NOR2X1_LOC_208/Y NOR2X1_LOC_35/Y 0.06fF
C56979 NOR2X1_LOC_448/B NAND2X1_LOC_425/Y 0.03fF
C56980 NAND2X1_LOC_576/a_36_24# INVX1_LOC_260/Y 0.00fF
C56981 NOR2X1_LOC_482/Y INVX1_LOC_6/A 0.00fF
C56982 INVX1_LOC_32/A INVX1_LOC_112/Y 0.01fF
C56983 NOR2X1_LOC_590/A INVX1_LOC_118/A 0.21fF
C56984 INVX1_LOC_224/Y INVX1_LOC_3/Y 0.17fF
C56985 INVX1_LOC_24/A VDD 1.03fF
C56986 NOR2X1_LOC_764/Y INVX1_LOC_89/A 0.01fF
C56987 NOR2X1_LOC_151/Y NOR2X1_LOC_687/Y 0.10fF
C56988 INVX1_LOC_269/A INVX1_LOC_123/Y 0.04fF
C56989 INVX1_LOC_278/A INVX1_LOC_42/A 0.10fF
C56990 INVX1_LOC_93/A INVX1_LOC_19/A 0.07fF
C56991 INVX1_LOC_77/A NOR2X1_LOC_567/a_36_216# 0.00fF
C56992 INVX1_LOC_162/A INVX1_LOC_95/A 0.02fF
C56993 NOR2X1_LOC_211/A NOR2X1_LOC_74/A 0.03fF
C56994 NOR2X1_LOC_86/Y NOR2X1_LOC_536/A 0.01fF
C56995 INVX1_LOC_149/A INVX1_LOC_91/A 0.03fF
C56996 INVX1_LOC_103/A NOR2X1_LOC_697/Y 0.02fF
C56997 NOR2X1_LOC_214/B D_GATE_366 0.03fF
C56998 NOR2X1_LOC_457/B INVX1_LOC_10/Y 0.03fF
C56999 NOR2X1_LOC_503/Y NOR2X1_LOC_88/Y 0.07fF
C57000 NOR2X1_LOC_113/B INVX1_LOC_1/Y 0.15fF
C57001 INVX1_LOC_271/A INVX1_LOC_128/A 0.01fF
C57002 NOR2X1_LOC_777/B NOR2X1_LOC_852/Y 0.03fF
C57003 NOR2X1_LOC_78/A INVX1_LOC_210/A 0.09fF
C57004 NAND2X1_LOC_516/a_36_24# INVX1_LOC_291/A 0.01fF
C57005 INVX1_LOC_71/A INVX1_LOC_117/A 0.10fF
C57006 INVX1_LOC_14/A INVX1_LOC_293/Y 0.07fF
C57007 NAND2X1_LOC_589/a_36_24# INVX1_LOC_118/A 0.00fF
C57008 INVX1_LOC_168/Y INVX1_LOC_306/Y 0.01fF
C57009 NOR2X1_LOC_557/Y VDD 1.40fF
C57010 INVX1_LOC_290/A INVX1_LOC_6/A 0.03fF
C57011 NOR2X1_LOC_609/A INVX1_LOC_9/A 0.05fF
C57012 NOR2X1_LOC_438/Y INVX1_LOC_181/A 0.07fF
C57013 NOR2X1_LOC_561/Y NOR2X1_LOC_815/A 0.01fF
C57014 NOR2X1_LOC_361/B NAND2X1_LOC_773/B 0.03fF
C57015 INVX1_LOC_314/Y INVX1_LOC_38/A 0.07fF
C57016 NOR2X1_LOC_391/B NOR2X1_LOC_719/B 0.04fF
C57017 NOR2X1_LOC_503/Y INVX1_LOC_84/A 0.70fF
C57018 NOR2X1_LOC_261/Y INVX1_LOC_78/A 0.01fF
C57019 INVX1_LOC_90/A NOR2X1_LOC_597/Y 0.01fF
C57020 NAND2X1_LOC_839/Y NAND2X1_LOC_836/Y 0.16fF
C57021 NOR2X1_LOC_458/Y NAND2X1_LOC_472/Y -0.02fF
C57022 NOR2X1_LOC_318/B INVX1_LOC_53/Y 0.01fF
C57023 INVX1_LOC_153/Y NAND2X1_LOC_472/Y 0.10fF
C57024 INVX1_LOC_14/A NAND2X1_LOC_74/B 1.76fF
C57025 INVX1_LOC_278/A INVX1_LOC_78/A 0.08fF
C57026 NOR2X1_LOC_419/Y INVX1_LOC_9/A 0.07fF
C57027 NAND2X1_LOC_205/A NAND2X1_LOC_99/A 0.02fF
C57028 INVX1_LOC_69/Y INVX1_LOC_150/A 0.20fF
C57029 NOR2X1_LOC_381/Y INVX1_LOC_12/A 0.15fF
C57030 NAND2X1_LOC_11/Y NAND2X1_LOC_1/Y 0.58fF
C57031 INVX1_LOC_308/Y NAND2X1_LOC_81/B 0.21fF
C57032 INVX1_LOC_13/A NOR2X1_LOC_78/A 0.50fF
C57033 INVX1_LOC_226/Y NOR2X1_LOC_124/A 0.02fF
C57034 INVX1_LOC_93/Y INVX1_LOC_53/Y 0.07fF
C57035 NOR2X1_LOC_433/A NOR2X1_LOC_351/Y 0.02fF
C57036 INVX1_LOC_1/Y NOR2X1_LOC_557/a_36_216# 0.00fF
C57037 NOR2X1_LOC_716/B INVX1_LOC_9/A 0.75fF
C57038 INVX1_LOC_224/A INVX1_LOC_106/Y 0.00fF
C57039 INVX1_LOC_89/A INVX1_LOC_69/Y 0.07fF
C57040 INVX1_LOC_30/A INVX1_LOC_119/Y 0.05fF
C57041 INVX1_LOC_164/A INVX1_LOC_91/A 0.06fF
C57042 INVX1_LOC_143/A VDD 0.00fF
C57043 INVX1_LOC_145/Y NOR2X1_LOC_318/B 0.01fF
C57044 INVX1_LOC_58/A INVX1_LOC_224/Y 0.01fF
C57045 NOR2X1_LOC_82/A NOR2X1_LOC_178/a_36_216# 0.00fF
C57046 INVX1_LOC_243/Y NOR2X1_LOC_598/B 0.25fF
C57047 INVX1_LOC_35/A NAND2X1_LOC_288/B 0.00fF
C57048 NAND2X1_LOC_215/A NAND2X1_LOC_205/a_36_24# 0.00fF
C57049 INVX1_LOC_72/A NAND2X1_LOC_475/Y 0.26fF
C57050 NOR2X1_LOC_590/A NAND2X1_LOC_63/Y 0.12fF
C57051 NOR2X1_LOC_219/Y INVX1_LOC_139/A 0.03fF
C57052 NOR2X1_LOC_554/B INVX1_LOC_84/A 0.03fF
C57053 NOR2X1_LOC_825/Y NAND2X1_LOC_859/B 0.30fF
C57054 NOR2X1_LOC_598/B INVX1_LOC_57/A 0.10fF
C57055 INVX1_LOC_68/Y VDD 0.49fF
C57056 INPUT_0 NAND2X1_LOC_855/Y 0.02fF
C57057 INVX1_LOC_36/Y NOR2X1_LOC_196/a_36_216# 0.00fF
C57058 INVX1_LOC_22/Y NAND2X1_LOC_63/Y 0.03fF
C57059 NOR2X1_LOC_152/Y NOR2X1_LOC_88/Y 0.07fF
C57060 NOR2X1_LOC_667/A INVX1_LOC_33/Y 0.10fF
C57061 NOR2X1_LOC_78/A NOR2X1_LOC_174/B 0.05fF
C57062 INVX1_LOC_51/A INVX1_LOC_57/A 0.03fF
C57063 INVX1_LOC_90/A NOR2X1_LOC_557/A 0.03fF
C57064 INVX1_LOC_248/A INVX1_LOC_33/Y 0.69fF
C57065 NAND2X1_LOC_565/B VDD 0.19fF
C57066 INVX1_LOC_142/A INVX1_LOC_186/Y 0.04fF
C57067 INVX1_LOC_174/Y INVX1_LOC_76/A 0.00fF
C57068 INVX1_LOC_58/A NAND2X1_LOC_793/B 0.07fF
C57069 NAND2X1_LOC_796/B NAND2X1_LOC_175/Y 0.02fF
C57070 INVX1_LOC_124/A NOR2X1_LOC_709/B 0.30fF
C57071 NAND2X1_LOC_711/Y NOR2X1_LOC_89/A 0.46fF
C57072 INVX1_LOC_210/Y INVX1_LOC_29/A 0.39fF
C57073 NOR2X1_LOC_315/Y INVX1_LOC_54/A 0.01fF
C57074 NOR2X1_LOC_52/B NOR2X1_LOC_177/a_36_216# 0.00fF
C57075 NOR2X1_LOC_130/A NOR2X1_LOC_56/Y 0.14fF
C57076 INVX1_LOC_21/A INVX1_LOC_23/Y 0.03fF
C57077 NOR2X1_LOC_843/B NOR2X1_LOC_849/A 0.03fF
C57078 INVX1_LOC_202/A NOR2X1_LOC_127/Y 0.53fF
C57079 NOR2X1_LOC_644/B INVX1_LOC_290/Y 0.02fF
C57080 NOR2X1_LOC_778/B INVX1_LOC_38/A 0.14fF
C57081 NAND2X1_LOC_123/a_36_24# NAND2X1_LOC_123/Y 0.02fF
C57082 NOR2X1_LOC_382/Y NOR2X1_LOC_671/Y 0.01fF
C57083 NAND2X1_LOC_560/A NOR2X1_LOC_526/a_36_216# 0.00fF
C57084 NOR2X1_LOC_68/A INVX1_LOC_49/Y 0.03fF
C57085 NOR2X1_LOC_152/Y INVX1_LOC_84/A 0.07fF
C57086 INVX1_LOC_300/A NOR2X1_LOC_765/Y 0.01fF
C57087 INVX1_LOC_30/A INVX1_LOC_284/A 0.00fF
C57088 NOR2X1_LOC_432/Y INVX1_LOC_54/A 0.02fF
C57089 NOR2X1_LOC_205/Y NOR2X1_LOC_334/Y 0.04fF
C57090 INVX1_LOC_50/A INVX1_LOC_13/Y 0.05fF
C57091 NOR2X1_LOC_360/Y INVX1_LOC_125/A 0.07fF
C57092 INVX1_LOC_25/Y NOR2X1_LOC_536/A 0.17fF
C57093 D_INPUT_1 INVX1_LOC_5/A 0.20fF
C57094 NAND2X1_LOC_783/A VDD 0.58fF
C57095 INVX1_LOC_35/A NOR2X1_LOC_405/Y 0.01fF
C57096 INVX1_LOC_113/Y INVX1_LOC_84/A 0.03fF
C57097 NAND2X1_LOC_800/Y VDD 0.22fF
C57098 NOR2X1_LOC_500/A INVX1_LOC_19/A 0.08fF
C57099 NOR2X1_LOC_322/Y NOR2X1_LOC_45/B 0.70fF
C57100 NOR2X1_LOC_130/A VDD 0.62fF
C57101 NOR2X1_LOC_68/A INVX1_LOC_99/A 0.01fF
C57102 INVX1_LOC_41/A NOR2X1_LOC_461/a_36_216# 0.00fF
C57103 NOR2X1_LOC_303/Y INVX1_LOC_19/A 0.06fF
C57104 NAND2X1_LOC_800/Y NAND2X1_LOC_800/A 0.01fF
C57105 NAND2X1_LOC_551/A NAND2X1_LOC_464/A 0.02fF
C57106 NOR2X1_LOC_757/a_36_216# INVX1_LOC_92/A 0.00fF
C57107 NAND2X1_LOC_652/Y NAND2X1_LOC_468/B 0.14fF
C57108 INVX1_LOC_45/A INVX1_LOC_3/Y 0.10fF
C57109 NAND2X1_LOC_650/B INPUT_1 0.00fF
C57110 NOR2X1_LOC_624/A NOR2X1_LOC_814/A -0.03fF
C57111 INVX1_LOC_64/Y NOR2X1_LOC_865/Y 0.07fF
C57112 NOR2X1_LOC_45/Y NOR2X1_LOC_158/Y 0.06fF
C57113 NOR2X1_LOC_719/B INVX1_LOC_280/A 0.03fF
C57114 INVX1_LOC_22/A INVX1_LOC_185/A 0.00fF
C57115 INVX1_LOC_134/A NOR2X1_LOC_863/B 0.35fF
C57116 INVX1_LOC_25/Y NAND2X1_LOC_93/B 0.36fF
C57117 INVX1_LOC_64/Y NOR2X1_LOC_243/B 0.55fF
C57118 INVX1_LOC_50/A INVX1_LOC_88/A 0.04fF
C57119 NOR2X1_LOC_441/Y INVX1_LOC_94/Y 0.17fF
C57120 NAND2X1_LOC_357/B NOR2X1_LOC_661/a_36_216# 0.00fF
C57121 INVX1_LOC_57/A NOR2X1_LOC_271/a_36_216# 0.01fF
C57122 NOR2X1_LOC_554/B INVX1_LOC_15/A 0.11fF
C57123 NOR2X1_LOC_254/Y INVX1_LOC_19/A 0.00fF
C57124 INVX1_LOC_11/A NOR2X1_LOC_635/B 0.03fF
C57125 INVX1_LOC_1/A INVX1_LOC_23/A 1.09fF
C57126 NAND2X1_LOC_36/a_36_24# INVX1_LOC_15/A 0.00fF
C57127 NOR2X1_LOC_717/B INVX1_LOC_9/A 0.03fF
C57128 NAND2X1_LOC_563/A INVX1_LOC_123/Y 0.02fF
C57129 NOR2X1_LOC_718/Y INVX1_LOC_12/A 0.00fF
C57130 NOR2X1_LOC_589/A NOR2X1_LOC_433/Y 0.30fF
C57131 NOR2X1_LOC_210/A INVX1_LOC_92/A 0.22fF
C57132 INVX1_LOC_150/Y NOR2X1_LOC_113/a_36_216# 0.00fF
C57133 INVX1_LOC_11/A NOR2X1_LOC_748/A 0.43fF
C57134 NOR2X1_LOC_514/Y NAND2X1_LOC_82/Y 0.02fF
C57135 NOR2X1_LOC_216/Y VDD 0.61fF
C57136 NOR2X1_LOC_784/Y INVX1_LOC_23/A 0.15fF
C57137 NOR2X1_LOC_555/a_36_216# NOR2X1_LOC_562/B 0.11fF
C57138 INVX1_LOC_113/Y NAND2X1_LOC_220/B 0.01fF
C57139 INVX1_LOC_58/A NOR2X1_LOC_103/Y 0.55fF
C57140 INVX1_LOC_66/A INVX1_LOC_54/A 0.02fF
C57141 INVX1_LOC_71/A INVX1_LOC_3/Y 0.02fF
C57142 NOR2X1_LOC_776/a_36_216# INVX1_LOC_57/A 0.02fF
C57143 NOR2X1_LOC_112/B VDD 0.07fF
C57144 INVX1_LOC_14/A NOR2X1_LOC_660/Y 0.05fF
C57145 INVX1_LOC_293/A NAND2X1_LOC_215/A 0.01fF
C57146 INVX1_LOC_162/A NAND2X1_LOC_807/B 0.38fF
C57147 INVX1_LOC_21/A NOR2X1_LOC_249/Y 1.02fF
C57148 NAND2X1_LOC_858/B NOR2X1_LOC_305/Y 0.11fF
C57149 INVX1_LOC_54/Y INVX1_LOC_19/A 0.07fF
C57150 NOR2X1_LOC_152/Y INVX1_LOC_15/A 0.30fF
C57151 NOR2X1_LOC_353/Y INVX1_LOC_19/A 0.01fF
C57152 NAND2X1_LOC_464/Y INVX1_LOC_42/A 0.02fF
C57153 INVX1_LOC_25/Y INVX1_LOC_3/A 0.03fF
C57154 NOR2X1_LOC_372/A INVX1_LOC_57/A 0.03fF
C57155 NAND2X1_LOC_656/Y NOR2X1_LOC_831/B 0.00fF
C57156 INVX1_LOC_75/A NOR2X1_LOC_536/A 0.04fF
C57157 INVX1_LOC_25/A INVX1_LOC_31/A 0.33fF
C57158 INVX1_LOC_93/Y NOR2X1_LOC_557/a_36_216# 0.01fF
C57159 INVX1_LOC_16/A INVX1_LOC_63/A 0.03fF
C57160 NOR2X1_LOC_493/B NOR2X1_LOC_89/A 0.03fF
C57161 INVX1_LOC_191/Y INVX1_LOC_261/Y 0.01fF
C57162 NAND2X1_LOC_861/Y NOR2X1_LOC_88/Y 0.07fF
C57163 NOR2X1_LOC_486/Y NOR2X1_LOC_601/Y 0.00fF
C57164 INVX1_LOC_285/Y NAND2X1_LOC_472/Y 0.10fF
C57165 NAND2X1_LOC_69/a_36_24# NAND2X1_LOC_114/B 0.00fF
C57166 INVX1_LOC_58/A INVX1_LOC_45/A 0.05fF
C57167 NOR2X1_LOC_15/Y NAND2X1_LOC_474/Y 0.01fF
C57168 NOR2X1_LOC_151/Y INVX1_LOC_9/A 0.42fF
C57169 INVX1_LOC_58/A NOR2X1_LOC_568/A 0.80fF
C57170 INVX1_LOC_174/A NAND2X1_LOC_31/a_36_24# 0.01fF
C57171 INVX1_LOC_120/A NAND2X1_LOC_85/Y 0.08fF
C57172 INVX1_LOC_58/A NAND2X1_LOC_856/A 0.03fF
C57173 NOR2X1_LOC_82/Y NAND2X1_LOC_63/Y 0.16fF
C57174 INVX1_LOC_316/Y INVX1_LOC_29/A 0.03fF
C57175 INVX1_LOC_247/A NAND2X1_LOC_602/a_36_24# 0.00fF
C57176 INVX1_LOC_21/A NOR2X1_LOC_636/B 0.13fF
C57177 INVX1_LOC_75/A NOR2X1_LOC_655/Y 0.05fF
C57178 NOR2X1_LOC_142/Y INVX1_LOC_94/Y 0.03fF
C57179 INVX1_LOC_34/A NAND2X1_LOC_454/Y 0.07fF
C57180 NAND2X1_LOC_787/A INVX1_LOC_72/A 0.03fF
C57181 INVX1_LOC_7/A NAND2X1_LOC_219/B 0.01fF
C57182 NAND2X1_LOC_861/Y INVX1_LOC_84/A 0.07fF
C57183 INVX1_LOC_18/A NOR2X1_LOC_629/A 0.02fF
C57184 NOR2X1_LOC_828/Y NOR2X1_LOC_778/A 0.20fF
C57185 NOR2X1_LOC_65/B NOR2X1_LOC_262/Y 0.09fF
C57186 INVX1_LOC_75/A NAND2X1_LOC_93/B 0.08fF
C57187 INVX1_LOC_165/Y NAND2X1_LOC_254/Y 0.01fF
C57188 NAND2X1_LOC_738/B INVX1_LOC_300/Y 0.03fF
C57189 INVX1_LOC_108/Y NOR2X1_LOC_554/B 0.06fF
C57190 INVX1_LOC_191/Y NOR2X1_LOC_467/A 0.29fF
C57191 INPUT_6 INVX1_LOC_18/A 0.62fF
C57192 INVX1_LOC_181/Y INVX1_LOC_29/Y 0.12fF
C57193 NOR2X1_LOC_209/A VDD -0.00fF
C57194 INVX1_LOC_35/A NOR2X1_LOC_751/Y 0.00fF
C57195 INVX1_LOC_30/Y INVX1_LOC_12/A -0.00fF
C57196 NOR2X1_LOC_78/A NOR2X1_LOC_319/B 0.01fF
C57197 INVX1_LOC_17/A NAND2X1_LOC_579/A 0.01fF
C57198 NOR2X1_LOC_250/Y NOR2X1_LOC_92/Y 0.07fF
C57199 INVX1_LOC_313/Y NAND2X1_LOC_475/Y 0.16fF
C57200 INVX1_LOC_303/A INVX1_LOC_50/A 0.07fF
C57201 NOR2X1_LOC_669/Y INVX1_LOC_11/A 0.01fF
C57202 INVX1_LOC_39/A NOR2X1_LOC_590/A 0.04fF
C57203 NOR2X1_LOC_557/A INVX1_LOC_38/A 0.03fF
C57204 INVX1_LOC_58/A INVX1_LOC_71/A 0.08fF
C57205 NOR2X1_LOC_818/a_36_216# NOR2X1_LOC_554/B 0.00fF
C57206 INVX1_LOC_75/A NAND2X1_LOC_425/Y 0.64fF
C57207 NOR2X1_LOC_550/B NOR2X1_LOC_383/B 0.01fF
C57208 NAND2X1_LOC_811/Y NOR2X1_LOC_829/A 0.00fF
C57209 NAND2X1_LOC_53/Y NOR2X1_LOC_15/Y 0.07fF
C57210 NOR2X1_LOC_381/Y INVX1_LOC_228/Y 0.05fF
C57211 NAND2X1_LOC_624/B INVX1_LOC_18/A 0.02fF
C57212 INVX1_LOC_176/A INVX1_LOC_37/A 0.03fF
C57213 VDD NOR2X1_LOC_280/Y 0.22fF
C57214 NOR2X1_LOC_593/Y NOR2X1_LOC_748/A 0.12fF
C57215 NAND2X1_LOC_149/a_36_24# INVX1_LOC_193/A 0.00fF
C57216 INVX1_LOC_28/A INVX1_LOC_63/A 0.04fF
C57217 NOR2X1_LOC_172/Y INVX1_LOC_271/A 0.03fF
C57218 NAND2X1_LOC_231/Y NAND2X1_LOC_454/Y 0.07fF
C57219 NOR2X1_LOC_315/Y NOR2X1_LOC_438/Y 0.02fF
C57220 INVX1_LOC_75/A NOR2X1_LOC_649/B 0.07fF
C57221 NAND2X1_LOC_112/Y INVX1_LOC_32/A 0.45fF
C57222 INVX1_LOC_75/A INVX1_LOC_3/A 2.32fF
C57223 INVX1_LOC_267/Y INVX1_LOC_175/A 0.01fF
C57224 INVX1_LOC_1/A INVX1_LOC_31/A 0.12fF
C57225 NOR2X1_LOC_513/Y INVX1_LOC_161/Y 0.05fF
C57226 NOR2X1_LOC_368/A NOR2X1_LOC_179/Y 0.07fF
C57227 INVX1_LOC_89/A NOR2X1_LOC_89/A 2.81fF
C57228 INVX1_LOC_188/A NAND2X1_LOC_190/Y 0.01fF
C57229 INVX1_LOC_309/A INVX1_LOC_260/Y 0.47fF
C57230 NOR2X1_LOC_65/B NOR2X1_LOC_63/a_36_216# -0.00fF
C57231 INVX1_LOC_36/A INVX1_LOC_48/Y 0.07fF
C57232 INVX1_LOC_136/A NOR2X1_LOC_792/a_36_216# 0.01fF
C57233 INVX1_LOC_172/A NAND2X1_LOC_624/B 0.46fF
C57234 NOR2X1_LOC_337/Y NOR2X1_LOC_197/B 0.85fF
C57235 INVX1_LOC_5/A D_INPUT_2 0.19fF
C57236 VDD NAND2X1_LOC_811/B 0.01fF
C57237 INVX1_LOC_13/Y NAND2X1_LOC_757/a_36_24# -0.01fF
C57238 NAND2X1_LOC_850/A INVX1_LOC_29/A 0.00fF
C57239 NOR2X1_LOC_510/Y INVX1_LOC_24/A 0.15fF
C57240 NOR2X1_LOC_78/A NOR2X1_LOC_259/B 0.02fF
C57241 NOR2X1_LOC_433/A NOR2X1_LOC_304/Y 0.27fF
C57242 INVX1_LOC_269/A INVX1_LOC_223/A 0.14fF
C57243 VDD NOR2X1_LOC_148/Y 0.24fF
C57244 INVX1_LOC_118/Y NAND2X1_LOC_211/Y 0.07fF
C57245 INVX1_LOC_136/A INVX1_LOC_14/A 0.21fF
C57246 NAND2X1_LOC_860/a_36_24# NAND2X1_LOC_793/Y 0.00fF
C57247 NAND2X1_LOC_650/B INVX1_LOC_118/A 0.07fF
C57248 NAND2X1_LOC_861/Y INVX1_LOC_15/A 0.07fF
C57249 NAND2X1_LOC_823/a_36_24# NOR2X1_LOC_865/Y 0.01fF
C57250 INVX1_LOC_188/Y INVX1_LOC_307/A 0.01fF
C57251 NOR2X1_LOC_166/Y NOR2X1_LOC_48/B 0.03fF
C57252 INVX1_LOC_48/A INVX1_LOC_293/Y 0.03fF
C57253 NOR2X1_LOC_717/B INVX1_LOC_274/Y 0.04fF
C57254 NAND2X1_LOC_347/B NOR2X1_LOC_81/a_36_216# 0.00fF
C57255 INVX1_LOC_45/A INVX1_LOC_215/Y 0.07fF
C57256 NAND2X1_LOC_11/Y NOR2X1_LOC_452/A 0.01fF
C57257 INVX1_LOC_1/A INVX1_LOC_111/A 0.01fF
C57258 NAND2X1_LOC_392/Y NOR2X1_LOC_278/Y 0.00fF
C57259 NOR2X1_LOC_643/Y NAND2X1_LOC_473/A 0.07fF
C57260 NAND2X1_LOC_214/B NOR2X1_LOC_392/B 0.01fF
C57261 D_INPUT_1 NOR2X1_LOC_773/Y 0.07fF
C57262 INVX1_LOC_64/Y NOR2X1_LOC_342/A 0.00fF
C57263 NOR2X1_LOC_361/B INVX1_LOC_24/A 0.13fF
C57264 NAND2X1_LOC_363/B NOR2X1_LOC_537/Y 0.07fF
C57265 INVX1_LOC_5/A NOR2X1_LOC_154/a_36_216# 0.02fF
C57266 NAND2X1_LOC_860/A NAND2X1_LOC_334/a_36_24# 0.00fF
C57267 NAND2X1_LOC_363/B NAND2X1_LOC_338/B 0.08fF
C57268 NAND2X1_LOC_303/Y NAND2X1_LOC_567/Y 0.00fF
C57269 NOR2X1_LOC_441/Y NOR2X1_LOC_524/Y 0.06fF
C57270 INVX1_LOC_48/A NAND2X1_LOC_74/B 0.59fF
C57271 INVX1_LOC_5/A NOR2X1_LOC_529/Y -0.01fF
C57272 NAND2X1_LOC_363/B NAND2X1_LOC_323/B 0.07fF
C57273 INVX1_LOC_27/A NOR2X1_LOC_392/B 0.10fF
C57274 NOR2X1_LOC_378/Y INVX1_LOC_193/A 0.10fF
C57275 NOR2X1_LOC_34/B NOR2X1_LOC_87/B 0.00fF
C57276 VDD NOR2X1_LOC_197/B 1.62fF
C57277 INVX1_LOC_31/A NOR2X1_LOC_384/Y 0.15fF
C57278 NAND2X1_LOC_561/B NAND2X1_LOC_632/B 0.02fF
C57279 NOR2X1_LOC_329/B INVX1_LOC_21/Y 0.04fF
C57280 NAND2X1_LOC_72/Y NOR2X1_LOC_203/Y 0.02fF
C57281 INVX1_LOC_129/Y INVX1_LOC_92/A 0.01fF
C57282 NAND2X1_LOC_79/Y NOR2X1_LOC_160/B 0.01fF
C57283 NAND2X1_LOC_583/a_36_24# INVX1_LOC_77/A 0.01fF
C57284 INVX1_LOC_30/A INVX1_LOC_72/A 0.46fF
C57285 NOR2X1_LOC_272/Y INVX1_LOC_133/Y 0.50fF
C57286 INVX1_LOC_123/A INVX1_LOC_42/A 0.08fF
C57287 NOR2X1_LOC_791/Y NAND2X1_LOC_338/B 0.01fF
C57288 NOR2X1_LOC_35/Y INVX1_LOC_63/A 0.12fF
C57289 INVX1_LOC_35/A INVX1_LOC_255/Y 0.07fF
C57290 NAND2X1_LOC_537/Y NAND2X1_LOC_811/Y 0.00fF
C57291 INVX1_LOC_12/Y INVX1_LOC_123/Y 0.10fF
C57292 NOR2X1_LOC_151/Y INVX1_LOC_274/Y 0.17fF
C57293 NAND2X1_LOC_464/A NAND2X1_LOC_489/Y 0.00fF
C57294 INVX1_LOC_269/A INVX1_LOC_149/Y 0.01fF
C57295 NOR2X1_LOC_773/Y NOR2X1_LOC_652/Y 0.35fF
C57296 D_INPUT_3 NOR2X1_LOC_814/A 0.10fF
C57297 NOR2X1_LOC_272/Y NOR2X1_LOC_67/A 0.35fF
C57298 INVX1_LOC_142/A INVX1_LOC_18/A 0.06fF
C57299 INVX1_LOC_75/A NAND2X1_LOC_470/B 0.16fF
C57300 D_INPUT_1 NOR2X1_LOC_332/A 0.19fF
C57301 NOR2X1_LOC_625/a_36_216# INVX1_LOC_30/A 0.00fF
C57302 INVX1_LOC_30/A INVX1_LOC_198/Y 0.01fF
C57303 INVX1_LOC_14/A NOR2X1_LOC_278/A 0.18fF
C57304 INVX1_LOC_14/Y NOR2X1_LOC_814/A 0.04fF
C57305 NOR2X1_LOC_124/A INVX1_LOC_12/A 0.02fF
C57306 INVX1_LOC_136/A NOR2X1_LOC_522/Y 0.04fF
C57307 INVX1_LOC_28/A NOR2X1_LOC_65/Y 0.03fF
C57308 NAND2X1_LOC_840/Y NAND2X1_LOC_175/Y 0.04fF
C57309 INVX1_LOC_90/A INVX1_LOC_271/A 0.03fF
C57310 INPUT_0 NAND2X1_LOC_454/Y 0.01fF
C57311 NAND2X1_LOC_739/B INVX1_LOC_136/A 0.13fF
C57312 INVX1_LOC_299/A NOR2X1_LOC_655/B 0.30fF
C57313 INVX1_LOC_136/A NAND2X1_LOC_84/Y 0.08fF
C57314 INVX1_LOC_18/A INVX1_LOC_41/Y 0.03fF
C57315 INVX1_LOC_278/A NAND2X1_LOC_861/Y 0.07fF
C57316 INVX1_LOC_35/A NOR2X1_LOC_71/Y 0.07fF
C57317 NOR2X1_LOC_15/Y INVX1_LOC_197/A 0.19fF
C57318 NOR2X1_LOC_78/A INVX1_LOC_32/A 0.05fF
C57319 NOR2X1_LOC_155/A INVX1_LOC_274/A 0.01fF
C57320 NOR2X1_LOC_189/A INVX1_LOC_36/A 0.03fF
C57321 NOR2X1_LOC_624/A NOR2X1_LOC_590/A 0.04fF
C57322 NOR2X1_LOC_478/A INVX1_LOC_34/A 0.00fF
C57323 NOR2X1_LOC_89/A NAND2X1_LOC_244/A 0.02fF
C57324 NOR2X1_LOC_591/Y NOR2X1_LOC_816/A 0.12fF
C57325 NOR2X1_LOC_78/A NOR2X1_LOC_623/B 3.88fF
C57326 INVX1_LOC_41/A INVX1_LOC_124/Y 0.07fF
C57327 NOR2X1_LOC_88/Y INVX1_LOC_291/A 0.08fF
C57328 INVX1_LOC_221/A INVX1_LOC_31/A 0.02fF
C57329 NOR2X1_LOC_188/A NOR2X1_LOC_668/Y 0.03fF
C57330 NOR2X1_LOC_168/B NOR2X1_LOC_785/A 0.12fF
C57331 NAND2X1_LOC_850/Y NAND2X1_LOC_793/Y 0.02fF
C57332 INVX1_LOC_7/Y D_INPUT_0 0.10fF
C57333 NOR2X1_LOC_92/Y NAND2X1_LOC_660/Y 0.07fF
C57334 NOR2X1_LOC_510/Y NOR2X1_LOC_130/A 0.07fF
C57335 NOR2X1_LOC_186/Y NOR2X1_LOC_246/A 0.81fF
C57336 INVX1_LOC_172/A INVX1_LOC_41/Y 0.03fF
C57337 INVX1_LOC_95/Y NOR2X1_LOC_38/B 0.09fF
C57338 INVX1_LOC_35/A NOR2X1_LOC_828/B 0.04fF
C57339 INVX1_LOC_17/A INVX1_LOC_208/Y 0.00fF
C57340 NAND2X1_LOC_198/B NAND2X1_LOC_316/a_36_24# 0.06fF
C57341 INVX1_LOC_34/A NOR2X1_LOC_68/A 0.21fF
C57342 INVX1_LOC_47/Y INVX1_LOC_20/A 0.00fF
C57343 NOR2X1_LOC_65/B INVX1_LOC_123/A -0.02fF
C57344 NOR2X1_LOC_188/A INVX1_LOC_23/A 0.28fF
C57345 NOR2X1_LOC_82/A INVX1_LOC_53/Y 0.03fF
C57346 INVX1_LOC_12/A NOR2X1_LOC_684/Y 0.00fF
C57347 INVX1_LOC_84/A NAND2X1_LOC_802/Y 0.12fF
C57348 NOR2X1_LOC_310/Y NOR2X1_LOC_274/B 0.01fF
C57349 NOR2X1_LOC_15/Y INVX1_LOC_10/A 0.66fF
C57350 INVX1_LOC_36/A NOR2X1_LOC_84/Y 0.07fF
C57351 INVX1_LOC_24/A INVX1_LOC_153/Y 0.01fF
C57352 NAND2X1_LOC_354/a_36_24# NAND2X1_LOC_798/A 0.00fF
C57353 NOR2X1_LOC_548/B INVX1_LOC_23/A 0.00fF
C57354 INVX1_LOC_256/A NAND2X1_LOC_349/B 0.10fF
C57355 NAND2X1_LOC_573/Y NOR2X1_LOC_246/A 0.01fF
C57356 INVX1_LOC_27/A INVX1_LOC_90/A 0.19fF
C57357 NOR2X1_LOC_92/Y D_INPUT_0 0.18fF
C57358 INVX1_LOC_25/A INVX1_LOC_6/A 0.07fF
C57359 INVX1_LOC_33/A INVX1_LOC_314/Y 0.04fF
C57360 INVX1_LOC_30/A NOR2X1_LOC_537/Y 0.03fF
C57361 NOR2X1_LOC_824/A INVX1_LOC_90/A 0.07fF
C57362 INVX1_LOC_247/A NOR2X1_LOC_464/Y 0.01fF
C57363 NAND2X1_LOC_722/A INVX1_LOC_72/A 0.07fF
C57364 NOR2X1_LOC_609/a_36_216# INVX1_LOC_155/Y 0.00fF
C57365 NAND2X1_LOC_338/B INVX1_LOC_30/A 0.12fF
C57366 INVX1_LOC_27/A NOR2X1_LOC_389/B 0.10fF
C57367 INVX1_LOC_305/A NOR2X1_LOC_175/A 0.32fF
C57368 INVX1_LOC_35/A NOR2X1_LOC_199/a_36_216# 0.00fF
C57369 INVX1_LOC_24/A INVX1_LOC_121/Y 0.00fF
C57370 NOR2X1_LOC_360/Y NOR2X1_LOC_709/A 0.10fF
C57371 INVX1_LOC_21/A NOR2X1_LOC_775/Y 0.04fF
C57372 INVX1_LOC_178/A NOR2X1_LOC_497/Y 0.01fF
C57373 NOR2X1_LOC_361/B NOR2X1_LOC_130/A 0.03fF
C57374 NAND2X1_LOC_656/B INVX1_LOC_19/A 0.01fF
C57375 NAND2X1_LOC_214/B NAND2X1_LOC_348/A 0.03fF
C57376 INVX1_LOC_32/A NOR2X1_LOC_60/Y 0.00fF
C57377 NAND2X1_LOC_470/B NAND2X1_LOC_453/A 0.01fF
C57378 INVX1_LOC_245/Y INVX1_LOC_121/A 0.00fF
C57379 INVX1_LOC_24/A INVX1_LOC_177/A 0.03fF
C57380 NOR2X1_LOC_78/A NOR2X1_LOC_622/A 0.01fF
C57381 INVX1_LOC_2/A NOR2X1_LOC_215/Y 0.05fF
C57382 INVX1_LOC_224/A INVX1_LOC_89/A 0.03fF
C57383 NOR2X1_LOC_230/Y INVX1_LOC_22/A 0.03fF
C57384 NOR2X1_LOC_230/a_36_216# INVX1_LOC_290/A 0.01fF
C57385 INVX1_LOC_49/A INVX1_LOC_104/A 0.12fF
C57386 NOR2X1_LOC_278/Y INVX1_LOC_46/A 2.69fF
C57387 INVX1_LOC_119/A NOR2X1_LOC_433/A 0.03fF
C57388 INVX1_LOC_27/A NAND2X1_LOC_348/A 0.07fF
C57389 INVX1_LOC_11/A INVX1_LOC_89/A 0.86fF
C57390 INVX1_LOC_293/A NOR2X1_LOC_99/B 0.01fF
C57391 NOR2X1_LOC_15/Y NOR2X1_LOC_302/Y 0.01fF
C57392 INVX1_LOC_280/Y INVX1_LOC_24/A 0.03fF
C57393 INVX1_LOC_36/A INVX1_LOC_290/A 0.10fF
C57394 NAND2X1_LOC_785/A NOR2X1_LOC_753/Y 0.23fF
C57395 NOR2X1_LOC_264/Y INVX1_LOC_8/A 0.07fF
C57396 NOR2X1_LOC_457/A INVX1_LOC_313/Y 0.07fF
C57397 INVX1_LOC_184/Y INVX1_LOC_143/A 0.04fF
C57398 NOR2X1_LOC_160/B NOR2X1_LOC_333/A 0.00fF
C57399 INVX1_LOC_71/A NOR2X1_LOC_357/a_36_216# 0.02fF
C57400 INVX1_LOC_88/A NAND2X1_LOC_652/Y 0.01fF
C57401 NOR2X1_LOC_785/A INVX1_LOC_132/Y 0.02fF
C57402 NOR2X1_LOC_654/A INVX1_LOC_76/A 0.10fF
C57403 INVX1_LOC_223/Y INVX1_LOC_69/Y 0.00fF
C57404 NAND2X1_LOC_859/Y NOR2X1_LOC_384/Y 0.15fF
C57405 NOR2X1_LOC_596/A NAND2X1_LOC_841/A 0.21fF
C57406 INVX1_LOC_314/Y INVX1_LOC_40/A 0.05fF
C57407 INVX1_LOC_291/A INVX1_LOC_15/A 0.07fF
C57408 NOR2X1_LOC_654/A NAND2X1_LOC_405/a_36_24# 0.00fF
C57409 NOR2X1_LOC_721/B INVX1_LOC_19/A 0.21fF
C57410 NOR2X1_LOC_176/Y INVX1_LOC_181/A 0.02fF
C57411 NOR2X1_LOC_778/B INVX1_LOC_33/A 0.04fF
C57412 INVX1_LOC_21/A NOR2X1_LOC_685/A 0.20fF
C57413 NOR2X1_LOC_662/A INVX1_LOC_29/A 0.03fF
C57414 VDD NOR2X1_LOC_260/Y 0.22fF
C57415 INVX1_LOC_122/Y INVX1_LOC_83/A 0.01fF
C57416 NAND2X1_LOC_81/B NAND2X1_LOC_773/B 0.03fF
C57417 NAND2X1_LOC_86/Y NOR2X1_LOC_849/A 0.01fF
C57418 INVX1_LOC_2/A INVX1_LOC_104/A 0.07fF
C57419 INVX1_LOC_136/A NOR2X1_LOC_137/A 0.39fF
C57420 INVX1_LOC_256/A INVX1_LOC_75/A 0.10fF
C57421 INVX1_LOC_1/A INVX1_LOC_6/A 0.13fF
C57422 INVX1_LOC_30/A INVX1_LOC_313/Y 0.06fF
C57423 INVX1_LOC_53/A NOR2X1_LOC_858/B 0.04fF
C57424 NOR2X1_LOC_647/B INVX1_LOC_75/A 0.01fF
C57425 NOR2X1_LOC_326/Y NOR2X1_LOC_324/Y 0.00fF
C57426 NOR2X1_LOC_142/Y INVX1_LOC_52/A 0.03fF
C57427 NAND2X1_LOC_182/A NOR2X1_LOC_226/A 0.15fF
C57428 INVX1_LOC_24/A NOR2X1_LOC_528/a_36_216# 0.01fF
C57429 INVX1_LOC_232/Y INVX1_LOC_80/Y 0.01fF
C57430 INVX1_LOC_8/A INVX1_LOC_316/Y 0.03fF
C57431 NOR2X1_LOC_332/A D_INPUT_2 0.07fF
C57432 D_INPUT_0 NAND2X1_LOC_837/Y 0.01fF
C57433 NAND2X1_LOC_53/Y NOR2X1_LOC_733/Y 0.03fF
C57434 INVX1_LOC_271/A INVX1_LOC_38/A 0.11fF
C57435 NOR2X1_LOC_778/B NOR2X1_LOC_714/Y 0.17fF
C57436 INVX1_LOC_21/A NAND2X1_LOC_447/Y 0.03fF
C57437 INVX1_LOC_17/A NOR2X1_LOC_501/B 0.01fF
C57438 INVX1_LOC_58/A NOR2X1_LOC_331/B 1.33fF
C57439 NOR2X1_LOC_392/B INVX1_LOC_137/A 0.38fF
C57440 NOR2X1_LOC_583/Y NOR2X1_LOC_584/Y 0.02fF
C57441 INVX1_LOC_31/A NOR2X1_LOC_188/A 0.07fF
C57442 VDD INVX1_LOC_38/Y 0.48fF
C57443 INVX1_LOC_2/A INVX1_LOC_263/A 0.07fF
C57444 INVX1_LOC_94/A NOR2X1_LOC_356/A -0.05fF
C57445 NOR2X1_LOC_468/Y INVX1_LOC_95/Y 0.07fF
C57446 NAND2X1_LOC_660/Y NAND2X1_LOC_477/A 0.54fF
C57447 INVX1_LOC_41/A D_INPUT_0 0.07fF
C57448 NOR2X1_LOC_142/Y INVX1_LOC_66/A 0.02fF
C57449 INVX1_LOC_89/A NOR2X1_LOC_593/Y 0.03fF
C57450 INVX1_LOC_201/Y D_INPUT_0 0.05fF
C57451 NAND2X1_LOC_286/B NAND2X1_LOC_288/A 0.04fF
C57452 INVX1_LOC_4/Y NAND2X1_LOC_773/B 0.10fF
C57453 NOR2X1_LOC_598/B INVX1_LOC_274/A 0.10fF
C57454 INVX1_LOC_230/Y INVX1_LOC_91/A -0.03fF
C57455 INVX1_LOC_57/A NOR2X1_LOC_634/A 0.08fF
C57456 INVX1_LOC_33/A NOR2X1_LOC_724/Y 0.02fF
C57457 NOR2X1_LOC_68/A INPUT_0 0.11fF
C57458 INVX1_LOC_2/A NAND2X1_LOC_854/B 0.03fF
C57459 INVX1_LOC_225/A NOR2X1_LOC_246/A 0.02fF
C57460 INVX1_LOC_310/A NAND2X1_LOC_358/Y 0.00fF
C57461 NOR2X1_LOC_67/A NOR2X1_LOC_86/A 0.42fF
C57462 INVX1_LOC_58/A NOR2X1_LOC_592/B 0.01fF
C57463 D_INPUT_0 NAND2X1_LOC_477/A 0.10fF
C57464 NOR2X1_LOC_328/Y NOR2X1_LOC_418/Y 0.15fF
C57465 INVX1_LOC_136/A INVX1_LOC_48/A 0.10fF
C57466 NOR2X1_LOC_470/B VDD 0.12fF
C57467 NOR2X1_LOC_772/Y NOR2X1_LOC_772/A 0.00fF
C57468 INVX1_LOC_94/A NOR2X1_LOC_74/A 0.07fF
C57469 NOR2X1_LOC_158/Y NOR2X1_LOC_48/Y 0.06fF
C57470 NAND2X1_LOC_286/B NOR2X1_LOC_653/Y 0.03fF
C57471 INVX1_LOC_89/A NOR2X1_LOC_52/B 0.03fF
C57472 NOR2X1_LOC_785/Y INVX1_LOC_143/A 0.02fF
C57473 INVX1_LOC_35/A NOR2X1_LOC_61/A 0.00fF
C57474 INVX1_LOC_78/A NAND2X1_LOC_449/a_36_24# 0.00fF
C57475 INVX1_LOC_27/A INVX1_LOC_38/A 0.06fF
C57476 INVX1_LOC_9/Y NAND2X1_LOC_112/Y 0.01fF
C57477 INVX1_LOC_1/Y INVX1_LOC_16/A 0.19fF
C57478 INVX1_LOC_26/Y NOR2X1_LOC_721/B 0.87fF
C57479 NOR2X1_LOC_215/a_36_216# NOR2X1_LOC_357/Y 0.01fF
C57480 NOR2X1_LOC_389/A INVX1_LOC_95/Y 0.16fF
C57481 NOR2X1_LOC_824/A INVX1_LOC_38/A 0.21fF
C57482 INVX1_LOC_5/A NOR2X1_LOC_61/Y 0.07fF
C57483 NOR2X1_LOC_831/B NOR2X1_LOC_717/A 0.10fF
C57484 INVX1_LOC_48/Y NOR2X1_LOC_102/a_36_216# 0.00fF
C57485 INVX1_LOC_103/A INVX1_LOC_37/A 0.08fF
C57486 INVX1_LOC_24/A INVX1_LOC_285/Y 0.03fF
C57487 NOR2X1_LOC_679/Y INVX1_LOC_20/A 0.16fF
C57488 NAND2X1_LOC_326/a_36_24# INVX1_LOC_28/A 0.00fF
C57489 INVX1_LOC_256/A NOR2X1_LOC_309/a_36_216# 0.01fF
C57490 INVX1_LOC_64/A NAND2X1_LOC_798/B 0.07fF
C57491 INVX1_LOC_38/Y NOR2X1_LOC_846/a_36_216# 0.01fF
C57492 INVX1_LOC_130/A NAND2X1_LOC_468/B 0.01fF
C57493 INVX1_LOC_206/A NOR2X1_LOC_355/a_36_216# 0.00fF
C57494 NOR2X1_LOC_545/A INPUT_0 0.01fF
C57495 NAND2X1_LOC_656/A INVX1_LOC_286/A 0.10fF
C57496 INVX1_LOC_26/A INVX1_LOC_125/A 0.46fF
C57497 NAND2X1_LOC_392/A NAND2X1_LOC_392/Y 0.01fF
C57498 NOR2X1_LOC_383/B INVX1_LOC_293/Y 0.01fF
C57499 NOR2X1_LOC_92/Y NAND2X1_LOC_848/A 0.18fF
C57500 NOR2X1_LOC_205/Y NAND2X1_LOC_472/Y 0.07fF
C57501 INVX1_LOC_83/A INVX1_LOC_83/Y 0.02fF
C57502 NAND2X1_LOC_286/B INVX1_LOC_19/A 0.09fF
C57503 NOR2X1_LOC_369/Y VDD 0.27fF
C57504 INVX1_LOC_284/Y NAND2X1_LOC_836/a_36_24# -0.02fF
C57505 NAND2X1_LOC_741/B NOR2X1_LOC_328/a_36_216# 0.03fF
C57506 INVX1_LOC_47/Y INVX1_LOC_4/A 0.10fF
C57507 NOR2X1_LOC_591/Y INVX1_LOC_140/A 0.05fF
C57508 INVX1_LOC_292/A INVX1_LOC_37/A 0.07fF
C57509 NOR2X1_LOC_664/Y NAND2X1_LOC_348/A 0.58fF
C57510 INVX1_LOC_34/A NOR2X1_LOC_2/Y 0.01fF
C57511 NOR2X1_LOC_551/a_36_216# INVX1_LOC_104/A 0.00fF
C57512 INVX1_LOC_243/Y INVX1_LOC_29/A 0.16fF
C57513 INVX1_LOC_109/A NOR2X1_LOC_65/Y 0.06fF
C57514 INVX1_LOC_7/Y INVX1_LOC_46/Y -0.03fF
C57515 INVX1_LOC_49/A INVX1_LOC_206/Y 0.03fF
C57516 NOR2X1_LOC_590/A INVX1_LOC_14/Y 0.49fF
C57517 NOR2X1_LOC_383/B NAND2X1_LOC_74/B 0.03fF
C57518 INVX1_LOC_284/Y INVX1_LOC_46/A 0.02fF
C57519 NOR2X1_LOC_210/A INVX1_LOC_83/A 0.01fF
C57520 INVX1_LOC_286/Y VDD 2.93fF
C57521 INVX1_LOC_287/Y INVX1_LOC_301/A -0.00fF
C57522 NOR2X1_LOC_216/Y INVX1_LOC_177/A 0.05fF
C57523 INVX1_LOC_57/A INVX1_LOC_29/A 0.85fF
C57524 INVX1_LOC_81/A NOR2X1_LOC_139/Y 0.08fF
C57525 NAND2X1_LOC_860/A INVX1_LOC_19/A 0.10fF
C57526 INVX1_LOC_286/Y NAND2X1_LOC_800/A 0.03fF
C57527 NOR2X1_LOC_457/B INVX1_LOC_247/A 0.13fF
C57528 NOR2X1_LOC_68/A NAND2X1_LOC_441/a_36_24# 0.01fF
C57529 INVX1_LOC_1/A NOR2X1_LOC_79/A 0.01fF
C57530 INVX1_LOC_218/Y NAND2X1_LOC_96/A 0.00fF
C57531 D_INPUT_1 INVX1_LOC_263/Y 0.01fF
C57532 INVX1_LOC_103/A INVX1_LOC_157/Y -0.04fF
C57533 NOR2X1_LOC_634/Y INVX1_LOC_19/A 0.04fF
C57534 NOR2X1_LOC_15/Y INVX1_LOC_307/A 0.03fF
C57535 NOR2X1_LOC_576/B INVX1_LOC_10/A 0.14fF
C57536 INVX1_LOC_223/A INVX1_LOC_12/Y 0.03fF
C57537 D_INPUT_1 NOR2X1_LOC_847/A 0.08fF
C57538 INVX1_LOC_81/A NAND2X1_LOC_468/B 0.01fF
C57539 INVX1_LOC_28/A INVX1_LOC_1/Y 0.03fF
C57540 INVX1_LOC_159/A INVX1_LOC_146/Y 0.27fF
C57541 D_INPUT_1 INVX1_LOC_42/A 0.13fF
C57542 NAND2X1_LOC_162/B INVX1_LOC_76/A 0.03fF
C57543 INVX1_LOC_90/A INVX1_LOC_234/A 0.05fF
C57544 INVX1_LOC_90/A NAND2X1_LOC_156/B 0.02fF
C57545 INVX1_LOC_215/A NOR2X1_LOC_329/B 0.03fF
C57546 NOR2X1_LOC_742/A INVX1_LOC_16/A 0.07fF
C57547 INVX1_LOC_33/A NOR2X1_LOC_657/B 0.04fF
C57548 INVX1_LOC_2/A INVX1_LOC_206/Y 0.14fF
C57549 NOR2X1_LOC_191/B VDD 0.53fF
C57550 NAND2X1_LOC_29/a_36_24# NAND2X1_LOC_207/Y 0.00fF
C57551 INVX1_LOC_279/A INVX1_LOC_182/Y 0.03fF
C57552 INVX1_LOC_48/Y INVX1_LOC_63/A 0.07fF
C57553 NOR2X1_LOC_716/B INVX1_LOC_76/A 0.12fF
C57554 NOR2X1_LOC_396/Y INVX1_LOC_240/A 0.00fF
C57555 INVX1_LOC_283/Y VDD -0.00fF
C57556 INVX1_LOC_19/A NAND2X1_LOC_473/A 0.01fF
C57557 NOR2X1_LOC_557/Y NAND2X1_LOC_267/B 0.02fF
C57558 NAND2X1_LOC_348/A INVX1_LOC_234/A 0.03fF
C57559 NOR2X1_LOC_338/Y NOR2X1_LOC_331/B 0.02fF
C57560 NAND2X1_LOC_662/B NAND2X1_LOC_660/Y 0.55fF
C57561 INVX1_LOC_41/A NOR2X1_LOC_266/B 0.20fF
C57562 NOR2X1_LOC_415/A INVX1_LOC_75/A 0.02fF
C57563 NOR2X1_LOC_160/B INVX1_LOC_123/Y 0.01fF
C57564 INVX1_LOC_30/A NAND2X1_LOC_444/a_36_24# 0.00fF
C57565 NOR2X1_LOC_545/a_36_216# INPUT_0 0.00fF
C57566 INVX1_LOC_143/A INVX1_LOC_65/A 0.04fF
C57567 INVX1_LOC_40/A NOR2X1_LOC_557/A 0.01fF
C57568 INVX1_LOC_90/A NOR2X1_LOC_19/B 0.07fF
C57569 NOR2X1_LOC_389/B NOR2X1_LOC_772/A 0.01fF
C57570 D_INPUT_1 INVX1_LOC_78/A 0.10fF
C57571 INVX1_LOC_18/A INVX1_LOC_185/A 0.03fF
C57572 NOR2X1_LOC_52/B NAND2X1_LOC_244/A 0.02fF
C57573 INVX1_LOC_278/A NOR2X1_LOC_89/a_36_216# 0.01fF
C57574 INVX1_LOC_1/A INVX1_LOC_301/A 0.61fF
C57575 INVX1_LOC_185/Y VDD -0.00fF
C57576 NOR2X1_LOC_657/Y NOR2X1_LOC_155/A 0.07fF
C57577 NOR2X1_LOC_778/B NOR2X1_LOC_486/Y 0.00fF
C57578 NOR2X1_LOC_281/Y INVX1_LOC_57/A 0.01fF
C57579 NOR2X1_LOC_276/Y NOR2X1_LOC_127/Y 0.02fF
C57580 NOR2X1_LOC_577/Y NOR2X1_LOC_536/A 0.00fF
C57581 NOR2X1_LOC_318/B INVX1_LOC_16/A 0.07fF
C57582 NOR2X1_LOC_639/B NOR2X1_LOC_158/B 0.03fF
C57583 NOR2X1_LOC_15/Y INVX1_LOC_12/A 0.35fF
C57584 INVX1_LOC_272/Y INVX1_LOC_49/Y 0.00fF
C57585 NOR2X1_LOC_340/Y NAND2X1_LOC_96/A 0.01fF
C57586 NOR2X1_LOC_447/A NOR2X1_LOC_654/A 0.02fF
C57587 INVX1_LOC_83/A INVX1_LOC_193/Y 0.03fF
C57588 NOR2X1_LOC_91/A NAND2X1_LOC_725/Y 0.03fF
C57589 NOR2X1_LOC_186/Y INVX1_LOC_32/A 0.10fF
C57590 NOR2X1_LOC_15/Y NOR2X1_LOC_519/Y 0.00fF
C57591 GATE_479 INVX1_LOC_91/A 0.03fF
C57592 NOR2X1_LOC_784/Y INVX1_LOC_301/A 0.15fF
C57593 NAND2X1_LOC_343/a_36_24# NOR2X1_LOC_318/B 0.00fF
C57594 INVX1_LOC_98/Y INVX1_LOC_76/A 0.37fF
C57595 INVX1_LOC_230/Y INVX1_LOC_203/A 0.03fF
C57596 NAND2X1_LOC_218/B NOR2X1_LOC_655/Y 0.09fF
C57597 NAND2X1_LOC_9/Y NOR2X1_LOC_278/Y 0.05fF
C57598 INVX1_LOC_93/Y INVX1_LOC_16/A 0.07fF
C57599 INVX1_LOC_72/A INVX1_LOC_113/A 0.45fF
C57600 INVX1_LOC_143/A NAND2X1_LOC_267/B -0.04fF
C57601 NOR2X1_LOC_65/B D_INPUT_1 0.37fF
C57602 NOR2X1_LOC_575/Y NAND2X1_LOC_463/B 0.01fF
C57603 INVX1_LOC_233/A NOR2X1_LOC_278/Y 0.01fF
C57604 NAND2X1_LOC_35/B VDD 0.01fF
C57605 NAND2X1_LOC_560/A NOR2X1_LOC_380/Y 0.04fF
C57606 NAND2X1_LOC_574/a_36_24# INVX1_LOC_32/A 0.00fF
C57607 NAND2X1_LOC_348/A NOR2X1_LOC_19/B 0.08fF
C57608 NAND2X1_LOC_361/a_36_24# NOR2X1_LOC_536/A 0.00fF
C57609 INVX1_LOC_13/A NAND2X1_LOC_642/Y 0.00fF
C57610 INVX1_LOC_45/A NAND2X1_LOC_475/Y 0.03fF
C57611 NAND2X1_LOC_729/Y NAND2X1_LOC_810/B 0.00fF
C57612 INVX1_LOC_172/A INVX1_LOC_185/A 0.03fF
C57613 INVX1_LOC_25/A INVX1_LOC_270/A 0.03fF
C57614 NOR2X1_LOC_78/B NOR2X1_LOC_858/B 0.19fF
C57615 NAND2X1_LOC_573/Y INVX1_LOC_32/A 0.26fF
C57616 INVX1_LOC_196/Y NOR2X1_LOC_728/B 0.38fF
C57617 INVX1_LOC_78/A NOR2X1_LOC_652/Y 0.07fF
C57618 NOR2X1_LOC_328/Y INVX1_LOC_20/A 0.03fF
C57619 NOR2X1_LOC_91/A NOR2X1_LOC_129/a_36_216# 0.00fF
C57620 NOR2X1_LOC_577/Y NAND2X1_LOC_93/B 0.07fF
C57621 INVX1_LOC_1/Y NOR2X1_LOC_35/Y 0.16fF
C57622 NOR2X1_LOC_516/B INVX1_LOC_36/Y 0.02fF
C57623 NOR2X1_LOC_590/A NOR2X1_LOC_831/Y 0.00fF
C57624 NOR2X1_LOC_186/Y NAND2X1_LOC_175/Y 0.07fF
C57625 NOR2X1_LOC_550/B INVX1_LOC_179/A 0.03fF
C57626 INVX1_LOC_16/A INVX1_LOC_139/A 0.03fF
C57627 NOR2X1_LOC_160/a_36_216# NAND2X1_LOC_425/Y 0.01fF
C57628 NOR2X1_LOC_312/Y NOR2X1_LOC_311/Y 0.01fF
C57629 INVX1_LOC_224/Y NAND2X1_LOC_363/B 0.01fF
C57630 INVX1_LOC_90/A NOR2X1_LOC_528/Y 0.01fF
C57631 INVX1_LOC_27/A NAND2X1_LOC_223/A 0.24fF
C57632 NOR2X1_LOC_718/Y INVX1_LOC_92/A 0.00fF
C57633 NOR2X1_LOC_371/a_36_216# INVX1_LOC_42/A 0.00fF
C57634 NOR2X1_LOC_246/A NAND2X1_LOC_642/Y 0.07fF
C57635 NOR2X1_LOC_428/a_36_216# NOR2X1_LOC_48/B 0.00fF
C57636 NOR2X1_LOC_379/Y NAND2X1_LOC_425/Y 0.03fF
C57637 INVX1_LOC_14/A NAND2X1_LOC_647/B 0.01fF
C57638 NOR2X1_LOC_346/B NOR2X1_LOC_536/A 0.03fF
C57639 NAND2X1_LOC_721/A INVX1_LOC_16/A 0.07fF
C57640 NAND2X1_LOC_218/B INVX1_LOC_3/A 1.24fF
C57641 NOR2X1_LOC_457/a_36_216# INVX1_LOC_271/Y 0.01fF
C57642 NOR2X1_LOC_203/a_36_216# NOR2X1_LOC_383/B 0.00fF
C57643 NOR2X1_LOC_423/Y INVX1_LOC_54/A 0.18fF
C57644 INVX1_LOC_69/Y INVX1_LOC_75/A 0.08fF
C57645 INVX1_LOC_235/Y INVX1_LOC_175/A 0.34fF
C57646 INVX1_LOC_89/A INVX1_LOC_199/A 0.02fF
C57647 NOR2X1_LOC_68/A NOR2X1_LOC_48/a_36_216# 0.00fF
C57648 INVX1_LOC_28/A NOR2X1_LOC_318/B 0.25fF
C57649 NAND2X1_LOC_573/Y NAND2X1_LOC_175/Y 0.02fF
C57650 NOR2X1_LOC_65/B NOR2X1_LOC_652/Y 0.01fF
C57651 NAND2X1_LOC_787/A NAND2X1_LOC_793/B 0.34fF
C57652 INVX1_LOC_71/A NAND2X1_LOC_475/Y 0.10fF
C57653 INVX1_LOC_219/A INVX1_LOC_20/A 0.01fF
C57654 INVX1_LOC_22/A NAND2X1_LOC_639/A 0.02fF
C57655 NOR2X1_LOC_382/Y INVX1_LOC_284/A 0.01fF
C57656 INVX1_LOC_249/Y INVX1_LOC_179/A 0.01fF
C57657 NAND2X1_LOC_479/Y INVX1_LOC_117/A 0.02fF
C57658 INVX1_LOC_89/A INVX1_LOC_74/A 0.07fF
C57659 INVX1_LOC_190/Y NOR2X1_LOC_56/Y 0.01fF
C57660 NOR2X1_LOC_251/Y INVX1_LOC_38/A 0.19fF
C57661 INVX1_LOC_227/A INVX1_LOC_14/Y 0.10fF
C57662 NAND2X1_LOC_708/Y NOR2X1_LOC_224/Y 0.12fF
C57663 NOR2X1_LOC_45/Y INVX1_LOC_32/A 0.29fF
C57664 NOR2X1_LOC_180/B INVX1_LOC_247/A 0.01fF
C57665 NAND2X1_LOC_724/A NAND2X1_LOC_175/Y 0.03fF
C57666 NOR2X1_LOC_83/Y NOR2X1_LOC_9/Y 0.08fF
C57667 INVX1_LOC_224/Y NOR2X1_LOC_791/Y 0.06fF
C57668 INVX1_LOC_22/A NOR2X1_LOC_536/A 0.12fF
C57669 NOR2X1_LOC_350/A INVX1_LOC_63/A 0.05fF
C57670 INVX1_LOC_298/Y NOR2X1_LOC_666/Y 0.07fF
C57671 NOR2X1_LOC_222/Y INVX1_LOC_54/A 0.09fF
C57672 NOR2X1_LOC_725/A INVX1_LOC_75/A 0.01fF
C57673 NOR2X1_LOC_91/A NAND2X1_LOC_326/A 0.08fF
C57674 NAND2X1_LOC_346/a_36_24# INVX1_LOC_26/A 0.00fF
C57675 NAND2X1_LOC_358/Y NAND2X1_LOC_96/A 0.06fF
C57676 INVX1_LOC_24/A NAND2X1_LOC_81/B 0.00fF
C57677 NOR2X1_LOC_336/a_36_216# INVX1_LOC_91/A 0.01fF
C57678 INVX1_LOC_5/A NOR2X1_LOC_678/A 0.49fF
C57679 INVX1_LOC_177/A NOR2X1_LOC_197/B 0.01fF
C57680 INVX1_LOC_53/A INVX1_LOC_50/Y 0.07fF
C57681 NAND2X1_LOC_740/B INVX1_LOC_11/Y 0.39fF
C57682 INVX1_LOC_13/A NOR2X1_LOC_271/Y 0.01fF
C57683 INVX1_LOC_190/Y VDD 0.32fF
C57684 INVX1_LOC_135/A INVX1_LOC_117/A 8.33fF
C57685 NOR2X1_LOC_717/B NAND2X1_LOC_418/a_36_24# 0.00fF
C57686 NAND2X1_LOC_41/Y INVX1_LOC_9/A 0.02fF
C57687 INVX1_LOC_36/A NOR2X1_LOC_467/A 0.01fF
C57688 INVX1_LOC_1/A INVX1_LOC_270/A 0.02fF
C57689 INPUT_6 D_INPUT_6 0.01fF
C57690 INVX1_LOC_314/Y INVX1_LOC_106/Y 0.01fF
C57691 INVX1_LOC_234/A INVX1_LOC_38/A 0.73fF
C57692 NAND2X1_LOC_337/B NOR2X1_LOC_318/A 0.08fF
C57693 D_INPUT_2 INVX1_LOC_42/A 0.00fF
C57694 INVX1_LOC_22/A NAND2X1_LOC_93/B 0.09fF
C57695 INVX1_LOC_6/A NOR2X1_LOC_43/Y 0.37fF
C57696 INVX1_LOC_101/Y INVX1_LOC_29/Y 0.10fF
C57697 INVX1_LOC_234/A NOR2X1_LOC_96/Y 0.03fF
C57698 D_GATE_741 NOR2X1_LOC_727/B 0.00fF
C57699 NOR2X1_LOC_690/Y INVX1_LOC_185/A 0.02fF
C57700 INVX1_LOC_28/A NAND2X1_LOC_721/A 0.17fF
C57701 INVX1_LOC_266/A INVX1_LOC_53/A 0.01fF
C57702 NOR2X1_LOC_84/Y INVX1_LOC_63/A 0.37fF
C57703 NOR2X1_LOC_143/a_36_216# INVX1_LOC_19/A 0.02fF
C57704 NOR2X1_LOC_307/A NOR2X1_LOC_383/B 0.05fF
C57705 INVX1_LOC_30/Y INVX1_LOC_92/A 0.03fF
C57706 INVX1_LOC_22/A NAND2X1_LOC_425/Y 0.01fF
C57707 NOR2X1_LOC_186/Y INVX1_LOC_171/Y 0.01fF
C57708 NOR2X1_LOC_360/Y NOR2X1_LOC_334/Y 0.10fF
C57709 NOR2X1_LOC_599/A NOR2X1_LOC_829/A 0.05fF
C57710 NOR2X1_LOC_721/Y VDD 0.26fF
C57711 INVX1_LOC_21/A NAND2X1_LOC_796/B 0.03fF
C57712 INVX1_LOC_234/A NAND2X1_LOC_848/Y -0.01fF
C57713 INVX1_LOC_24/A INVX1_LOC_4/Y 0.13fF
C57714 NOR2X1_LOC_457/B NOR2X1_LOC_465/Y 0.01fF
C57715 INVX1_LOC_17/A NOR2X1_LOC_639/B 0.17fF
C57716 INVX1_LOC_132/A INVX1_LOC_32/A 0.07fF
C57717 INVX1_LOC_11/A NOR2X1_LOC_392/Y 0.07fF
C57718 NOR2X1_LOC_33/A NAND2X1_LOC_574/A 0.06fF
C57719 INVX1_LOC_226/Y NAND2X1_LOC_456/Y 0.01fF
C57720 INVX1_LOC_83/A NOR2X1_LOC_809/B 0.45fF
C57721 NAND2X1_LOC_363/B NOR2X1_LOC_103/Y 0.63fF
C57722 INVX1_LOC_35/A NOR2X1_LOC_817/Y 0.02fF
C57723 NOR2X1_LOC_329/B NOR2X1_LOC_602/B 0.03fF
C57724 INVX1_LOC_96/Y INVX1_LOC_12/A 0.07fF
C57725 NOR2X1_LOC_596/A INVX1_LOC_271/Y 0.09fF
C57726 NOR2X1_LOC_168/A NAND2X1_LOC_74/B 0.00fF
C57727 NOR2X1_LOC_78/A NOR2X1_LOC_332/B 0.00fF
C57728 NOR2X1_LOC_689/A INVX1_LOC_136/A 0.02fF
C57729 NAND2X1_LOC_784/A INVX1_LOC_31/A 0.03fF
C57730 NOR2X1_LOC_591/Y INVX1_LOC_42/A 0.06fF
C57731 NOR2X1_LOC_804/B NOR2X1_LOC_801/B 0.01fF
C57732 NOR2X1_LOC_632/Y INVX1_LOC_84/A 0.03fF
C57733 NOR2X1_LOC_45/B NAND2X1_LOC_241/Y 0.02fF
C57734 NOR2X1_LOC_679/Y INVX1_LOC_64/A 0.02fF
C57735 NOR2X1_LOC_329/B INVX1_LOC_54/A 0.42fF
C57736 INVX1_LOC_136/A NOR2X1_LOC_383/B 0.10fF
C57737 INVX1_LOC_277/A INVX1_LOC_23/A 0.11fF
C57738 NOR2X1_LOC_337/Y VDD 0.18fF
C57739 NAND2X1_LOC_721/B INVX1_LOC_57/A 0.78fF
C57740 NOR2X1_LOC_711/A INVX1_LOC_117/A 0.01fF
C57741 INVX1_LOC_225/A INVX1_LOC_32/A 0.10fF
C57742 INVX1_LOC_90/A NOR2X1_LOC_216/B 0.03fF
C57743 D_INPUT_0 NAND2X1_LOC_574/A 0.05fF
C57744 INVX1_LOC_25/A INVX1_LOC_36/A 5.96fF
C57745 NOR2X1_LOC_156/A INVX1_LOC_92/A 0.07fF
C57746 NOR2X1_LOC_648/a_36_216# INVX1_LOC_290/Y 0.00fF
C57747 NOR2X1_LOC_557/Y INVX1_LOC_4/Y 0.03fF
C57748 INVX1_LOC_28/A INVX1_LOC_117/Y 0.00fF
C57749 NOR2X1_LOC_389/B NOR2X1_LOC_216/B 0.10fF
C57750 INVX1_LOC_223/Y INVX1_LOC_11/A 0.01fF
C57751 NOR2X1_LOC_248/Y INVX1_LOC_53/A 0.01fF
C57752 INVX1_LOC_30/A NAND2X1_LOC_793/B 0.07fF
C57753 NOR2X1_LOC_500/Y INVX1_LOC_99/A 0.03fF
C57754 D_INPUT_1 NOR2X1_LOC_554/B 0.26fF
C57755 INVX1_LOC_45/A NAND2X1_LOC_363/B 0.07fF
C57756 NAND2X1_LOC_213/A NAND2X1_LOC_209/a_36_24# 0.02fF
C57757 INVX1_LOC_25/Y NOR2X1_LOC_89/A 0.05fF
C57758 NOR2X1_LOC_244/B NOR2X1_LOC_240/B 0.14fF
C57759 NAND2X1_LOC_687/A NAND2X1_LOC_655/A 0.06fF
C57760 NAND2X1_LOC_656/A NAND2X1_LOC_215/A 0.10fF
C57761 NOR2X1_LOC_363/Y NOR2X1_LOC_139/Y 0.00fF
C57762 NAND2X1_LOC_503/a_36_24# INVX1_LOC_50/Y 0.00fF
C57763 VDD NOR2X1_LOC_56/Y 0.32fF
C57764 INVX1_LOC_62/A NOR2X1_LOC_721/B 0.01fF
C57765 VDD NAND2X1_LOC_659/B 0.02fF
C57766 NOR2X1_LOC_188/A NOR2X1_LOC_79/A 0.06fF
C57767 INVX1_LOC_8/A NOR2X1_LOC_55/a_36_216# 0.01fF
C57768 NAND2X1_LOC_348/A NOR2X1_LOC_216/B 0.03fF
C57769 NOR2X1_LOC_591/Y INVX1_LOC_78/A 0.00fF
C57770 NOR2X1_LOC_15/Y INVX1_LOC_200/A 0.01fF
C57771 INVX1_LOC_82/Y NAND2X1_LOC_141/Y 0.12fF
C57772 INVX1_LOC_37/A INVX1_LOC_143/Y 0.01fF
C57773 NOR2X1_LOC_74/A NOR2X1_LOC_155/A 0.06fF
C57774 INVX1_LOC_45/A NOR2X1_LOC_840/A 0.05fF
C57775 INVX1_LOC_143/A INVX1_LOC_4/Y 0.10fF
C57776 NOR2X1_LOC_363/Y NAND2X1_LOC_468/B 0.11fF
C57777 INVX1_LOC_45/A NOR2X1_LOC_791/Y 0.03fF
C57778 NAND2X1_LOC_187/a_36_24# INVX1_LOC_53/A 0.00fF
C57779 INVX1_LOC_146/Y VDD 0.55fF
C57780 NAND2X1_LOC_787/A INVX1_LOC_71/A 0.00fF
C57781 NAND2X1_LOC_287/B INVX1_LOC_46/A 0.07fF
C57782 NOR2X1_LOC_92/Y NOR2X1_LOC_134/Y 0.03fF
C57783 INVX1_LOC_132/A NOR2X1_LOC_622/A 0.10fF
C57784 INVX1_LOC_85/Y INVX1_LOC_19/A 0.03fF
C57785 NOR2X1_LOC_352/a_36_216# INVX1_LOC_9/A 0.02fF
C57786 NOR2X1_LOC_709/A NOR2X1_LOC_316/a_36_216# 0.01fF
C57787 INVX1_LOC_33/A INVX1_LOC_271/A 0.03fF
C57788 INVX1_LOC_11/A NAND2X1_LOC_357/A 0.07fF
C57789 INVX1_LOC_233/Y INVX1_LOC_24/A 0.22fF
C57790 NOR2X1_LOC_9/Y NOR2X1_LOC_155/A 0.01fF
C57791 NAND2X1_LOC_326/A INVX1_LOC_31/A 0.07fF
C57792 INVX1_LOC_33/Y INVX1_LOC_20/A 0.07fF
C57793 NOR2X1_LOC_709/A INVX1_LOC_26/A 0.21fF
C57794 INVX1_LOC_13/Y NOR2X1_LOC_791/B 0.01fF
C57795 INVX1_LOC_8/A INVX1_LOC_57/A 0.33fF
C57796 NAND2X1_LOC_200/B NAND2X1_LOC_223/A 0.17fF
C57797 NOR2X1_LOC_220/A INVX1_LOC_271/Y 0.10fF
C57798 INVX1_LOC_58/A NOR2X1_LOC_388/Y 0.10fF
C57799 NOR2X1_LOC_15/Y NAND2X1_LOC_733/Y 0.03fF
C57800 NAND2X1_LOC_778/Y INVX1_LOC_217/A 0.10fF
C57801 NOR2X1_LOC_285/B INVX1_LOC_23/A 0.09fF
C57802 NOR2X1_LOC_355/A NOR2X1_LOC_114/Y 0.00fF
C57803 NOR2X1_LOC_181/Y NOR2X1_LOC_748/A 0.03fF
C57804 NAND2X1_LOC_538/Y INVX1_LOC_141/A 0.07fF
C57805 NOR2X1_LOC_824/A NAND2X1_LOC_501/a_36_24# 0.00fF
C57806 INPUT_4 INVX1_LOC_54/A 0.22fF
C57807 NAND2X1_LOC_852/Y NAND2X1_LOC_175/Y 0.10fF
C57808 NOR2X1_LOC_229/a_36_216# NOR2X1_LOC_158/Y 0.01fF
C57809 INVX1_LOC_208/Y INVX1_LOC_94/Y 0.00fF
C57810 NAND2X1_LOC_852/Y NOR2X1_LOC_821/a_36_216# 0.15fF
C57811 NOR2X1_LOC_655/B NAND2X1_LOC_99/A 0.44fF
C57812 INVX1_LOC_25/A NOR2X1_LOC_309/Y 0.03fF
C57813 INVX1_LOC_22/A NAND2X1_LOC_470/B 0.07fF
C57814 NAND2X1_LOC_652/Y INVX1_LOC_272/A 0.02fF
C57815 NOR2X1_LOC_272/Y INVX1_LOC_181/Y 0.19fF
C57816 INVX1_LOC_36/A INVX1_LOC_1/A 0.51fF
C57817 INVX1_LOC_40/Y INVX1_LOC_14/A 0.02fF
C57818 INVX1_LOC_162/A INVX1_LOC_308/A 0.01fF
C57819 NOR2X1_LOC_211/A NAND2X1_LOC_71/a_36_24# 0.00fF
C57820 INVX1_LOC_16/A INVX1_LOC_87/A 0.03fF
C57821 NAND2X1_LOC_601/a_36_24# NOR2X1_LOC_109/Y 0.00fF
C57822 INVX1_LOC_135/A INVX1_LOC_3/Y 0.39fF
C57823 NOR2X1_LOC_15/Y INVX1_LOC_217/A 0.01fF
C57824 NOR2X1_LOC_575/Y INVX1_LOC_42/A 0.01fF
C57825 NOR2X1_LOC_857/A NOR2X1_LOC_729/A 0.39fF
C57826 NOR2X1_LOC_121/A INVX1_LOC_16/Y 0.39fF
C57827 NOR2X1_LOC_497/Y INVX1_LOC_42/A 0.01fF
C57828 NOR2X1_LOC_103/Y INVX1_LOC_30/A 0.05fF
C57829 NOR2X1_LOC_778/B NOR2X1_LOC_748/A 0.03fF
C57830 NAND2X1_LOC_214/B INVX1_LOC_33/A 0.01fF
C57831 NOR2X1_LOC_91/A NOR2X1_LOC_165/Y 0.01fF
C57832 NAND2X1_LOC_370/a_36_24# NOR2X1_LOC_309/Y 0.07fF
C57833 NAND2X1_LOC_587/a_36_24# INVX1_LOC_1/A 0.01fF
C57834 INVX1_LOC_75/A NOR2X1_LOC_89/A 0.10fF
C57835 INVX1_LOC_277/Y NOR2X1_LOC_307/A 0.01fF
C57836 NOR2X1_LOC_329/B NOR2X1_LOC_48/B 0.01fF
C57837 NOR2X1_LOC_173/Y NAND2X1_LOC_593/Y 0.06fF
C57838 NAND2X1_LOC_53/Y NOR2X1_LOC_722/Y 0.03fF
C57839 INVX1_LOC_122/A INVX1_LOC_9/A 0.06fF
C57840 NAND2X1_LOC_853/Y INVX1_LOC_296/Y 0.09fF
C57841 INVX1_LOC_256/A NOR2X1_LOC_274/B 0.02fF
C57842 INVX1_LOC_58/A NOR2X1_LOC_366/B 0.03fF
C57843 INVX1_LOC_223/A NOR2X1_LOC_160/B 0.68fF
C57844 NOR2X1_LOC_208/Y INVX1_LOC_1/A 0.01fF
C57845 INVX1_LOC_103/A NAND2X1_LOC_198/B 0.01fF
C57846 INVX1_LOC_27/A INVX1_LOC_33/A 0.20fF
C57847 NOR2X1_LOC_205/Y INVX1_LOC_24/A 0.00fF
C57848 NOR2X1_LOC_74/A NOR2X1_LOC_833/B 0.01fF
C57849 NOR2X1_LOC_92/Y INVX1_LOC_49/A 1.56fF
C57850 INVX1_LOC_34/A NAND2X1_LOC_474/Y 0.07fF
C57851 NOR2X1_LOC_121/A NAND2X1_LOC_205/A 0.14fF
C57852 INVX1_LOC_225/A INVX1_LOC_171/Y 0.02fF
C57853 INVX1_LOC_24/Y INVX1_LOC_49/A 0.03fF
C57854 NOR2X1_LOC_733/Y INVX1_LOC_12/A 0.21fF
C57855 INVX1_LOC_269/A INVX1_LOC_77/A 0.28fF
C57856 INVX1_LOC_58/A NAND2X1_LOC_479/Y 0.07fF
C57857 INVX1_LOC_75/A NOR2X1_LOC_170/A 0.01fF
C57858 INVX1_LOC_41/Y NAND2X1_LOC_793/Y 0.13fF
C57859 INVX1_LOC_304/Y NAND2X1_LOC_778/Y 0.10fF
C57860 INVX1_LOC_45/A INVX1_LOC_30/A 0.35fF
C57861 NAND2X1_LOC_720/a_36_24# INVX1_LOC_141/Y 0.00fF
C57862 NOR2X1_LOC_602/A INVX1_LOC_312/Y 0.12fF
C57863 NAND2X1_LOC_740/B INVX1_LOC_231/A 0.02fF
C57864 NOR2X1_LOC_457/A INVX1_LOC_71/A 0.00fF
C57865 INVX1_LOC_30/A NOR2X1_LOC_568/A 0.13fF
C57866 D_INPUT_4 NAND2X1_LOC_3/B 0.02fF
C57867 NAND2X1_LOC_218/B NOR2X1_LOC_647/B 0.03fF
C57868 NAND2X1_LOC_763/B INVX1_LOC_45/A 0.05fF
C57869 INVX1_LOC_233/A NAND2X1_LOC_392/A 0.01fF
C57870 NAND2X1_LOC_303/Y NAND2X1_LOC_354/B 0.01fF
C57871 NOR2X1_LOC_567/B NOR2X1_LOC_334/Y 0.07fF
C57872 NOR2X1_LOC_230/Y INVX1_LOC_18/A 0.01fF
C57873 NAND2X1_LOC_842/B NOR2X1_LOC_278/Y 0.05fF
C57874 NOR2X1_LOC_88/A NOR2X1_LOC_536/A 0.19fF
C57875 NOR2X1_LOC_328/Y INVX1_LOC_64/A 0.01fF
C57876 NOR2X1_LOC_78/B INVX1_LOC_50/Y 0.03fF
C57877 NAND2X1_LOC_532/a_36_24# NOR2X1_LOC_304/Y 0.01fF
C57878 INVX1_LOC_256/A NOR2X1_LOC_577/Y 0.11fF
C57879 NOR2X1_LOC_684/Y INVX1_LOC_92/A 0.02fF
C57880 NOR2X1_LOC_348/B NOR2X1_LOC_348/Y 0.19fF
C57881 NAND2X1_LOC_214/B INVX1_LOC_40/A 0.07fF
C57882 NOR2X1_LOC_561/A NOR2X1_LOC_216/B 0.01fF
C57883 INVX1_LOC_1/A NOR2X1_LOC_309/Y 0.05fF
C57884 INVX1_LOC_35/A INVX1_LOC_215/A 0.07fF
C57885 INVX1_LOC_211/Y NAND2X1_LOC_798/a_36_24# 0.00fF
C57886 NOR2X1_LOC_443/Y INVX1_LOC_132/Y 0.00fF
C57887 INVX1_LOC_58/A INVX1_LOC_135/A 0.04fF
C57888 NAND2X1_LOC_796/B NOR2X1_LOC_667/A 0.35fF
C57889 INVX1_LOC_35/A NOR2X1_LOC_195/a_36_216# 0.00fF
C57890 NOR2X1_LOC_409/Y NOR2X1_LOC_409/B 0.02fF
C57891 NAND2X1_LOC_364/Y NOR2X1_LOC_785/A 0.03fF
C57892 NAND2X1_LOC_729/Y INVX1_LOC_36/A 0.03fF
C57893 NAND2X1_LOC_53/Y INVX1_LOC_34/A 0.07fF
C57894 NAND2X1_LOC_796/B INVX1_LOC_248/A 0.01fF
C57895 INVX1_LOC_284/Y NAND2X1_LOC_866/A 0.31fF
C57896 INVX1_LOC_14/A NAND2X1_LOC_122/a_36_24# 0.06fF
C57897 INVX1_LOC_42/Y NAND2X1_LOC_454/Y 0.01fF
C57898 NOR2X1_LOC_804/B NOR2X1_LOC_794/B 0.11fF
C57899 NOR2X1_LOC_27/Y INVX1_LOC_269/A 0.01fF
C57900 INVX1_LOC_2/A NOR2X1_LOC_92/Y 0.17fF
C57901 INVX1_LOC_124/A INVX1_LOC_269/A 0.10fF
C57902 NOR2X1_LOC_455/Y NOR2X1_LOC_717/B 0.00fF
C57903 NOR2X1_LOC_615/Y NOR2X1_LOC_690/A 0.03fF
C57904 INVX1_LOC_27/A INVX1_LOC_40/A 2.05fF
C57905 NAND2X1_LOC_725/Y NAND2X1_LOC_866/B 0.10fF
C57906 INVX1_LOC_24/A NOR2X1_LOC_723/Y 0.06fF
C57907 INVX1_LOC_30/A INVX1_LOC_71/A 0.96fF
C57908 NOR2X1_LOC_270/Y NOR2X1_LOC_457/B 0.11fF
C57909 INVX1_LOC_230/Y NAND2X1_LOC_276/Y 0.07fF
C57910 NOR2X1_LOC_226/A NOR2X1_LOC_92/Y 0.15fF
C57911 INVX1_LOC_64/A INVX1_LOC_219/A 0.01fF
C57912 INVX1_LOC_228/Y NAND2X1_LOC_141/A 0.00fF
C57913 VDD INVX1_LOC_133/A 0.27fF
C57914 INVX1_LOC_172/Y NOR2X1_LOC_474/a_36_216# 0.00fF
C57915 NAND2X1_LOC_102/a_36_24# NAND2X1_LOC_99/A 0.02fF
C57916 NOR2X1_LOC_456/Y NOR2X1_LOC_644/A 0.01fF
C57917 NAND2X1_LOC_35/Y D_INPUT_0 0.07fF
C57918 NAND2X1_LOC_784/A NAND2X1_LOC_807/Y 0.59fF
C57919 INVX1_LOC_32/A NAND2X1_LOC_642/Y 0.04fF
C57920 NOR2X1_LOC_331/B NAND2X1_LOC_475/Y 0.10fF
C57921 NOR2X1_LOC_598/B NOR2X1_LOC_356/A 0.10fF
C57922 INVX1_LOC_136/A NAND2X1_LOC_632/B 0.04fF
C57923 NAND2X1_LOC_254/Y NAND2X1_LOC_244/A 0.00fF
C57924 NOR2X1_LOC_186/a_36_216# INVX1_LOC_84/A 0.01fF
C57925 INVX1_LOC_99/Y INVX1_LOC_97/A 0.02fF
C57926 NOR2X1_LOC_188/A INVX1_LOC_28/Y 0.22fF
C57927 INVX1_LOC_95/Y INVX1_LOC_251/A 0.02fF
C57928 INVX1_LOC_83/A INVX1_LOC_50/Y 0.07fF
C57929 INVX1_LOC_206/Y NOR2X1_LOC_631/Y 0.03fF
C57930 INVX1_LOC_31/A NOR2X1_LOC_87/B 0.06fF
C57931 NAND2X1_LOC_59/B D_INPUT_7 0.18fF
C57932 NOR2X1_LOC_456/a_36_216# INVX1_LOC_279/A 0.00fF
C57933 INVX1_LOC_229/A NAND2X1_LOC_579/a_36_24# 0.00fF
C57934 NOR2X1_LOC_791/Y NOR2X1_LOC_123/B 0.00fF
C57935 NAND2X1_LOC_1/Y INVX1_LOC_15/A 0.41fF
C57936 NOR2X1_LOC_150/a_36_216# NOR2X1_LOC_652/Y 0.01fF
C57937 INVX1_LOC_11/A INVX1_LOC_25/Y 0.03fF
C57938 INVX1_LOC_101/Y INVX1_LOC_101/A 0.05fF
C57939 INVX1_LOC_12/Y INVX1_LOC_290/Y 0.03fF
C57940 NOR2X1_LOC_807/B NOR2X1_LOC_325/A 0.38fF
C57941 INVX1_LOC_276/A NAND2X1_LOC_516/a_36_24# 0.00fF
C57942 NOR2X1_LOC_802/A NOR2X1_LOC_500/B 0.12fF
C57943 INVX1_LOC_93/A INVX1_LOC_90/A 0.13fF
C57944 NOR2X1_LOC_82/A INVX1_LOC_16/A 0.13fF
C57945 NOR2X1_LOC_188/A NOR2X1_LOC_416/A 0.07fF
C57946 NOR2X1_LOC_815/A INVX1_LOC_23/A 0.00fF
C57947 NAND2X1_LOC_642/Y NAND2X1_LOC_175/Y 0.39fF
C57948 NOR2X1_LOC_598/B NOR2X1_LOC_74/A 0.12fF
C57949 INVX1_LOC_103/A NOR2X1_LOC_665/A 2.55fF
C57950 INVX1_LOC_256/A INVX1_LOC_22/A 0.81fF
C57951 NAND2X1_LOC_190/Y INVX1_LOC_279/A 0.55fF
C57952 NOR2X1_LOC_312/Y NAND2X1_LOC_703/Y 0.03fF
C57953 NAND2X1_LOC_9/Y NOR2X1_LOC_97/A 0.02fF
C57954 NOR2X1_LOC_310/Y INVX1_LOC_18/A 0.01fF
C57955 NAND2X1_LOC_861/a_36_24# NAND2X1_LOC_793/Y 0.00fF
C57956 NOR2X1_LOC_454/Y NOR2X1_LOC_214/B 1.94fF
C57957 NAND2X1_LOC_93/B INVX1_LOC_186/Y 0.07fF
C57958 NAND2X1_LOC_328/a_36_24# INVX1_LOC_53/A 0.00fF
C57959 INVX1_LOC_6/Y INVX1_LOC_33/A 0.01fF
C57960 INVX1_LOC_101/Y NOR2X1_LOC_355/A 0.01fF
C57961 NOR2X1_LOC_78/B NOR2X1_LOC_248/Y 0.02fF
C57962 NOR2X1_LOC_92/Y NAND2X1_LOC_648/A 0.00fF
C57963 NOR2X1_LOC_813/Y INVX1_LOC_3/Y 0.08fF
C57964 INVX1_LOC_226/Y NAND2X1_LOC_208/B 0.53fF
C57965 INVX1_LOC_207/Y INVX1_LOC_239/A 0.01fF
C57966 INVX1_LOC_41/A INVX1_LOC_49/A 4.78fF
C57967 NOR2X1_LOC_92/Y INPUT_1 0.03fF
C57968 NOR2X1_LOC_269/a_36_216# NOR2X1_LOC_441/Y 0.00fF
C57969 INVX1_LOC_35/A INVX1_LOC_286/A 0.07fF
C57970 INVX1_LOC_223/A INVX1_LOC_208/A 0.09fF
C57971 INVX1_LOC_280/A INVX1_LOC_3/Y 0.84fF
C57972 INVX1_LOC_20/A INVX1_LOC_23/Y 0.09fF
C57973 NOR2X1_LOC_591/Y NOR2X1_LOC_152/Y 0.02fF
C57974 NOR2X1_LOC_94/Y INVX1_LOC_3/Y 0.04fF
C57975 INVX1_LOC_279/A NOR2X1_LOC_389/A 0.10fF
C57976 INVX1_LOC_265/A NAND2X1_LOC_833/Y 0.33fF
C57977 INVX1_LOC_161/A INVX1_LOC_10/A 0.07fF
C57978 INVX1_LOC_2/A NAND2X1_LOC_837/Y 0.06fF
C57979 NOR2X1_LOC_655/B NAND2X1_LOC_656/A 0.10fF
C57980 INVX1_LOC_163/A INVX1_LOC_135/Y 0.02fF
C57981 INVX1_LOC_99/A INVX1_LOC_307/A 0.04fF
C57982 NOR2X1_LOC_13/Y NAND2X1_LOC_655/a_36_24# 0.00fF
C57983 INVX1_LOC_136/A NAND2X1_LOC_170/A 0.03fF
C57984 NOR2X1_LOC_739/Y INVX1_LOC_196/Y 0.01fF
C57985 INPUT_0 NAND2X1_LOC_474/Y 0.07fF
C57986 NOR2X1_LOC_678/a_36_216# INVX1_LOC_75/A 0.13fF
C57987 INVX1_LOC_99/A NOR2X1_LOC_445/B 0.00fF
C57988 NOR2X1_LOC_401/B INVX1_LOC_314/Y 0.22fF
C57989 NAND2X1_LOC_195/Y NAND2X1_LOC_662/Y 0.00fF
C57990 NAND2X1_LOC_190/Y INVX1_LOC_182/Y 0.01fF
C57991 NAND2X1_LOC_733/Y NOR2X1_LOC_576/B 0.02fF
C57992 NOR2X1_LOC_82/A INVX1_LOC_28/A 0.07fF
C57993 NAND2X1_LOC_741/B INVX1_LOC_229/Y 0.12fF
C57994 NOR2X1_LOC_456/Y NOR2X1_LOC_540/B 0.03fF
C57995 INVX1_LOC_54/Y NOR2X1_LOC_772/Y 0.03fF
C57996 INVX1_LOC_35/A INVX1_LOC_95/A 0.03fF
C57997 INVX1_LOC_41/A INVX1_LOC_2/A 0.03fF
C57998 NOR2X1_LOC_781/Y INVX1_LOC_22/A 0.45fF
C57999 NAND2X1_LOC_222/B INVX1_LOC_75/A 0.06fF
C58000 NOR2X1_LOC_681/Y NOR2X1_LOC_677/Y 0.01fF
C58001 NAND2X1_LOC_807/Y NAND2X1_LOC_807/A 0.00fF
C58002 NOR2X1_LOC_78/B NOR2X1_LOC_718/Y 0.05fF
C58003 INVX1_LOC_76/A NOR2X1_LOC_591/A 0.05fF
C58004 NOR2X1_LOC_392/Y INVX1_LOC_74/A 0.01fF
C58005 NAND2X1_LOC_350/A NOR2X1_LOC_329/B 0.04fF
C58006 INVX1_LOC_41/A NOR2X1_LOC_226/A 0.16fF
C58007 INVX1_LOC_54/Y NOR2X1_LOC_392/B 0.29fF
C58008 INVX1_LOC_11/A INVX1_LOC_75/A 1.95fF
C58009 NOR2X1_LOC_843/A INVX1_LOC_143/A 0.02fF
C58010 INVX1_LOC_58/A INVX1_LOC_139/Y 0.02fF
C58011 INVX1_LOC_21/A NOR2X1_LOC_78/A 1.46fF
C58012 NOR2X1_LOC_222/Y NOR2X1_LOC_142/Y 0.11fF
C58013 NOR2X1_LOC_251/Y INVX1_LOC_33/A 0.04fF
C58014 NAND2X1_LOC_349/B NOR2X1_LOC_433/A 0.01fF
C58015 INVX1_LOC_2/A NAND2X1_LOC_477/A 0.07fF
C58016 INVX1_LOC_279/A NOR2X1_LOC_596/A 0.07fF
C58017 GATE_579 NAND2X1_LOC_463/B 0.03fF
C58018 NOR2X1_LOC_250/Y INVX1_LOC_144/A 0.01fF
C58019 INVX1_LOC_217/A NOR2X1_LOC_576/B 0.06fF
C58020 NAND2X1_LOC_785/A NAND2X1_LOC_775/a_36_24# 0.01fF
C58021 NAND2X1_LOC_364/A INVX1_LOC_148/Y 0.08fF
C58022 NOR2X1_LOC_441/Y NOR2X1_LOC_329/B 0.06fF
C58023 INVX1_LOC_238/A NOR2X1_LOC_380/Y 0.06fF
C58024 INVX1_LOC_58/A NOR2X1_LOC_813/Y 0.04fF
C58025 INVX1_LOC_226/Y INVX1_LOC_34/A 0.03fF
C58026 INVX1_LOC_26/A NOR2X1_LOC_489/A 0.04fF
C58027 NOR2X1_LOC_226/A NAND2X1_LOC_477/A 0.10fF
C58028 NOR2X1_LOC_664/Y INVX1_LOC_40/A 0.03fF
C58029 INVX1_LOC_273/A INVX1_LOC_92/A 0.03fF
C58030 INVX1_LOC_227/A NOR2X1_LOC_106/Y 0.02fF
C58031 NAND2X1_LOC_564/B NAND2X1_LOC_640/Y 0.01fF
C58032 NAND2X1_LOC_656/A NOR2X1_LOC_99/B 0.03fF
C58033 NOR2X1_LOC_510/Y NOR2X1_LOC_56/Y 0.01fF
C58034 INVX1_LOC_33/A INVX1_LOC_137/A 0.01fF
C58035 INVX1_LOC_268/A INVX1_LOC_63/Y 0.01fF
C58036 INVX1_LOC_27/A NOR2X1_LOC_486/Y 0.07fF
C58037 NAND2X1_LOC_551/A NOR2X1_LOC_91/Y 0.00fF
C58038 NAND2X1_LOC_35/Y NAND2X1_LOC_839/a_36_24# 0.01fF
C58039 INVX1_LOC_77/A NOR2X1_LOC_97/a_36_216# 0.01fF
C58040 INVX1_LOC_58/A INVX1_LOC_280/A 0.04fF
C58041 NOR2X1_LOC_52/B INVX1_LOC_25/Y 3.91fF
C58042 INVX1_LOC_89/A INVX1_LOC_314/Y 0.13fF
C58043 NOR2X1_LOC_351/Y INVX1_LOC_271/A 0.20fF
C58044 NAND2X1_LOC_349/B NOR2X1_LOC_52/B 0.59fF
C58045 INVX1_LOC_90/A NOR2X1_LOC_303/Y 0.03fF
C58046 NOR2X1_LOC_510/Y VDD 1.45fF
C58047 INVX1_LOC_34/A INVX1_LOC_10/A 0.46fF
C58048 NOR2X1_LOC_773/Y NOR2X1_LOC_191/A 0.04fF
C58049 INPUT_2 INVX1_LOC_315/Y 0.01fF
C58050 NOR2X1_LOC_389/B NOR2X1_LOC_303/Y 0.02fF
C58051 NOR2X1_LOC_835/A INVX1_LOC_134/Y 0.06fF
C58052 NAND2X1_LOC_35/Y NAND2X1_LOC_848/A 0.07fF
C58053 INVX1_LOC_36/A NOR2X1_LOC_188/A 0.00fF
C58054 NOR2X1_LOC_644/A NOR2X1_LOC_550/B 0.01fF
C58055 INVX1_LOC_182/Y NOR2X1_LOC_596/A 0.03fF
C58056 INVX1_LOC_63/Y NOR2X1_LOC_367/a_36_216# 0.01fF
C58057 INVX1_LOC_97/A NOR2X1_LOC_254/Y 0.06fF
C58058 INVX1_LOC_83/A NOR2X1_LOC_6/B 0.02fF
C58059 NAND2X1_LOC_390/a_36_24# NAND2X1_LOC_850/Y 0.00fF
C58060 INVX1_LOC_35/A INVX1_LOC_54/A 0.14fF
C58061 NOR2X1_LOC_234/Y D_INPUT_0 0.02fF
C58062 INVX1_LOC_41/A INPUT_1 0.05fF
C58063 INVX1_LOC_152/Y NOR2X1_LOC_61/Y 0.28fF
C58064 INVX1_LOC_278/Y INVX1_LOC_16/A 0.06fF
C58065 INVX1_LOC_2/A INVX1_LOC_121/A 0.08fF
C58066 NOR2X1_LOC_598/B NOR2X1_LOC_650/a_36_216# 0.01fF
C58067 INVX1_LOC_201/Y INPUT_1 0.09fF
C58068 INVX1_LOC_234/A NOR2X1_LOC_521/a_36_216# 0.00fF
C58069 INVX1_LOC_89/A NOR2X1_LOC_181/Y 0.03fF
C58070 NAND2X1_LOC_515/a_36_24# INVX1_LOC_79/A 0.00fF
C58071 INVX1_LOC_227/A NAND2X1_LOC_675/a_36_24# 0.00fF
C58072 INVX1_LOC_269/A NOR2X1_LOC_138/a_36_216# 0.01fF
C58073 INVX1_LOC_259/Y INVX1_LOC_179/A 0.02fF
C58074 INVX1_LOC_40/A INVX1_LOC_137/A 0.05fF
C58075 NAND2X1_LOC_231/Y INVX1_LOC_10/A 1.16fF
C58076 NOR2X1_LOC_557/Y NAND2X1_LOC_830/a_36_24# 0.01fF
C58077 NOR2X1_LOC_561/a_36_216# NAND2X1_LOC_842/B 0.00fF
C58078 NOR2X1_LOC_361/B VDD 2.71fF
C58079 NOR2X1_LOC_160/B INVX1_LOC_314/A 0.03fF
C58080 NOR2X1_LOC_286/Y NOR2X1_LOC_857/A 0.01fF
C58081 NOR2X1_LOC_433/A INVX1_LOC_75/A 0.10fF
C58082 NAND2X1_LOC_552/a_36_24# NAND2X1_LOC_862/A 0.01fF
C58083 NOR2X1_LOC_220/A INVX1_LOC_279/A 0.10fF
C58084 NAND2X1_LOC_117/a_36_24# NOR2X1_LOC_709/A 0.00fF
C58085 NOR2X1_LOC_180/B NOR2X1_LOC_180/Y 0.00fF
C58086 NAND2X1_LOC_724/A NAND2X1_LOC_804/Y 0.01fF
C58087 INVX1_LOC_11/A NAND2X1_LOC_453/A 0.07fF
C58088 NOR2X1_LOC_598/B NOR2X1_LOC_865/Y 0.07fF
C58089 NAND2X1_LOC_350/A NAND2X1_LOC_468/a_36_24# 0.01fF
C58090 NOR2X1_LOC_716/B NOR2X1_LOC_716/a_36_216# 0.00fF
C58091 NOR2X1_LOC_593/Y INVX1_LOC_75/A 0.16fF
C58092 NOR2X1_LOC_598/B NOR2X1_LOC_243/B 0.07fF
C58093 NOR2X1_LOC_47/a_36_216# NOR2X1_LOC_11/Y 0.02fF
C58094 INVX1_LOC_88/A NOR2X1_LOC_363/Y 0.03fF
C58095 NOR2X1_LOC_440/Y INVX1_LOC_22/A 0.22fF
C58096 INVX1_LOC_90/A INVX1_LOC_54/Y 0.23fF
C58097 INVX1_LOC_87/Y NOR2X1_LOC_612/B 0.01fF
C58098 NOR2X1_LOC_366/Y NOR2X1_LOC_131/Y 0.23fF
C58099 NOR2X1_LOC_778/B INVX1_LOC_89/A 0.03fF
C58100 NOR2X1_LOC_391/A NOR2X1_LOC_719/A 0.46fF
C58101 INVX1_LOC_25/A INVX1_LOC_63/A 0.23fF
C58102 NOR2X1_LOC_389/B INVX1_LOC_54/Y 0.10fF
C58103 NOR2X1_LOC_594/a_36_216# INVX1_LOC_63/Y 0.01fF
C58104 NOR2X1_LOC_33/Y NOR2X1_LOC_33/B -0.01fF
C58105 NAND2X1_LOC_778/Y INVX1_LOC_92/A 0.74fF
C58106 NOR2X1_LOC_344/A NOR2X1_LOC_337/A 0.03fF
C58107 NOR2X1_LOC_92/Y INVX1_LOC_118/A 0.24fF
C58108 NOR2X1_LOC_52/B INVX1_LOC_75/A 1.10fF
C58109 NOR2X1_LOC_521/a_36_216# NOR2X1_LOC_19/B 0.01fF
C58110 INVX1_LOC_64/A INVX1_LOC_220/A 0.47fF
C58111 NAND2X1_LOC_306/a_36_24# NOR2X1_LOC_45/B 0.01fF
C58112 NAND2X1_LOC_741/B INVX1_LOC_20/A 0.47fF
C58113 INVX1_LOC_269/A INVX1_LOC_9/A 0.10fF
C58114 NAND2X1_LOC_799/A NOR2X1_LOC_536/A 0.13fF
C58115 INVX1_LOC_171/A INVX1_LOC_232/A 0.02fF
C58116 NOR2X1_LOC_254/A NOR2X1_LOC_698/Y 0.16fF
C58117 NOR2X1_LOC_489/B NOR2X1_LOC_814/A 0.03fF
C58118 INVX1_LOC_108/A NAND2X1_LOC_473/A 0.01fF
C58119 NOR2X1_LOC_296/Y NOR2X1_LOC_271/Y 0.01fF
C58120 NOR2X1_LOC_309/Y NOR2X1_LOC_188/A 0.00fF
C58121 NOR2X1_LOC_6/B NOR2X1_LOC_193/a_36_216# 0.12fF
C58122 NOR2X1_LOC_457/A NOR2X1_LOC_331/B 0.03fF
C58123 INVX1_LOC_223/A NAND2X1_LOC_211/Y 0.30fF
C58124 NOR2X1_LOC_379/Y NOR2X1_LOC_725/A 0.14fF
C58125 NOR2X1_LOC_19/B INVX1_LOC_40/A 0.11fF
C58126 NOR2X1_LOC_15/Y INVX1_LOC_92/A 0.07fF
C58127 NOR2X1_LOC_667/A NAND2X1_LOC_840/Y 0.08fF
C58128 NAND2X1_LOC_351/A INVX1_LOC_37/A 0.09fF
C58129 NAND2X1_LOC_853/a_36_24# NAND2X1_LOC_866/A 0.01fF
C58130 INVX1_LOC_248/A NAND2X1_LOC_840/Y 0.01fF
C58131 INVX1_LOC_23/Y INVX1_LOC_4/A 0.07fF
C58132 NOR2X1_LOC_792/a_36_216# INVX1_LOC_285/A 0.00fF
C58133 NOR2X1_LOC_620/B INVX1_LOC_158/Y 0.03fF
C58134 INVX1_LOC_50/Y NOR2X1_LOC_68/Y 0.03fF
C58135 INVX1_LOC_72/A INVX1_LOC_202/Y 0.00fF
C58136 INVX1_LOC_35/A NAND2X1_LOC_807/B 0.00fF
C58137 NAND2X1_LOC_360/B INVX1_LOC_6/A 0.04fF
C58138 NOR2X1_LOC_337/Y INVX1_LOC_177/A 0.02fF
C58139 NOR2X1_LOC_678/A INVX1_LOC_42/A 0.00fF
C58140 INVX1_LOC_30/A NOR2X1_LOC_331/B 0.19fF
C58141 NAND2X1_LOC_647/B NOR2X1_LOC_383/B 0.00fF
C58142 NOR2X1_LOC_500/Y INPUT_0 0.13fF
C58143 INVX1_LOC_226/Y INPUT_0 0.03fF
C58144 INVX1_LOC_184/Y VDD -0.00fF
C58145 NAND2X1_LOC_21/Y NAND2X1_LOC_1/Y 0.52fF
C58146 INVX1_LOC_47/Y INVX1_LOC_129/A -0.03fF
C58147 INVX1_LOC_29/A INVX1_LOC_306/Y 0.03fF
C58148 INVX1_LOC_18/A NOR2X1_LOC_536/A 0.28fF
C58149 INVX1_LOC_14/A INVX1_LOC_285/A 0.09fF
C58150 INVX1_LOC_64/A NAND2X1_LOC_410/a_36_24# 0.00fF
C58151 NOR2X1_LOC_433/A NAND2X1_LOC_453/A 0.07fF
C58152 NOR2X1_LOC_142/Y NOR2X1_LOC_69/A 0.03fF
C58153 INVX1_LOC_89/A NOR2X1_LOC_724/Y 0.06fF
C58154 INVX1_LOC_14/A INVX1_LOC_265/Y 0.02fF
C58155 INVX1_LOC_131/A INVX1_LOC_10/A 0.07fF
C58156 NOR2X1_LOC_750/Y INVX1_LOC_32/A 0.04fF
C58157 NOR2X1_LOC_570/A NOR2X1_LOC_74/A 0.01fF
C58158 INVX1_LOC_62/Y NOR2X1_LOC_98/B 0.01fF
C58159 INVX1_LOC_14/A NOR2X1_LOC_814/A 0.12fF
C58160 INVX1_LOC_1/A INVX1_LOC_63/A 2.45fF
C58161 NAND2X1_LOC_660/Y INVX1_LOC_144/A 0.07fF
C58162 NOR2X1_LOC_275/a_36_216# NOR2X1_LOC_155/A 0.00fF
C58163 NOR2X1_LOC_636/A INVX1_LOC_37/A 0.01fF
C58164 NAND2X1_LOC_170/A NOR2X1_LOC_165/a_36_216# 0.00fF
C58165 NAND2X1_LOC_35/Y NOR2X1_LOC_754/A -0.01fF
C58166 INVX1_LOC_120/A NAND2X1_LOC_506/a_36_24# 0.00fF
C58167 INVX1_LOC_69/Y INVX1_LOC_22/A 0.07fF
C58168 INVX1_LOC_77/A INVX1_LOC_12/Y 0.10fF
C58169 NOR2X1_LOC_132/Y VDD 0.12fF
C58170 INVX1_LOC_50/A NOR2X1_LOC_409/B 0.03fF
C58171 INVX1_LOC_225/A NOR2X1_LOC_279/Y 0.01fF
C58172 NOR2X1_LOC_394/Y INVX1_LOC_23/A 0.02fF
C58173 NOR2X1_LOC_458/Y VDD 0.24fF
C58174 INVX1_LOC_153/Y VDD 1.06fF
C58175 NOR2X1_LOC_647/Y NOR2X1_LOC_655/Y 0.08fF
C58176 NOR2X1_LOC_65/B NOR2X1_LOC_318/A 0.03fF
C58177 INPUT_0 INVX1_LOC_10/A 3.60fF
C58178 NAND2X1_LOC_581/Y VDD 0.01fF
C58179 NOR2X1_LOC_303/Y INVX1_LOC_38/A 3.91fF
C58180 INVX1_LOC_24/Y NAND2X1_LOC_63/Y 0.07fF
C58181 INVX1_LOC_172/A NOR2X1_LOC_536/A 0.03fF
C58182 INVX1_LOC_256/A NAND2X1_LOC_476/Y 0.01fF
C58183 D_INPUT_0 INVX1_LOC_144/A 0.01fF
C58184 INVX1_LOC_53/A INVX1_LOC_273/A 0.03fF
C58185 NOR2X1_LOC_791/B NOR2X1_LOC_99/Y 0.30fF
C58186 INVX1_LOC_121/Y VDD 0.28fF
C58187 NOR2X1_LOC_78/B INVX1_LOC_188/Y 0.01fF
C58188 NOR2X1_LOC_361/B INVX1_LOC_133/A 0.42fF
C58189 INVX1_LOC_104/A INVX1_LOC_14/Y 0.10fF
C58190 NOR2X1_LOC_52/B NAND2X1_LOC_453/A 0.07fF
C58191 INVX1_LOC_18/A NAND2X1_LOC_93/B 0.14fF
C58192 NAND2X1_LOC_837/Y INVX1_LOC_118/A 0.09fF
C58193 NOR2X1_LOC_794/B INVX1_LOC_63/A 0.07fF
C58194 INVX1_LOC_78/A NOR2X1_LOC_678/A 0.03fF
C58195 NOR2X1_LOC_92/Y NAND2X1_LOC_455/B 0.11fF
C58196 INVX1_LOC_177/A VDD 1.18fF
C58197 NAND2X1_LOC_580/a_36_24# INVX1_LOC_240/Y 0.00fF
C58198 NOR2X1_LOC_807/B NOR2X1_LOC_777/B 0.06fF
C58199 NAND2X1_LOC_348/A NOR2X1_LOC_112/Y 0.01fF
C58200 NOR2X1_LOC_254/Y INVX1_LOC_38/A 0.03fF
C58201 INVX1_LOC_124/A INVX1_LOC_12/Y 0.01fF
C58202 NOR2X1_LOC_795/Y INVX1_LOC_117/A 0.10fF
C58203 INVX1_LOC_23/A NOR2X1_LOC_654/A 0.15fF
C58204 INVX1_LOC_280/Y VDD 0.73fF
C58205 INVX1_LOC_47/Y NOR2X1_LOC_440/B 0.02fF
C58206 INVX1_LOC_11/A NAND2X1_LOC_291/B 0.11fF
C58207 INVX1_LOC_31/A NAND2X1_LOC_219/B 0.13fF
C58208 INVX1_LOC_16/A INVX1_LOC_59/Y 0.09fF
C58209 INVX1_LOC_64/A INVX1_LOC_23/Y 0.02fF
C58210 NOR2X1_LOC_647/Y NOR2X1_LOC_649/B 0.13fF
C58211 NAND2X1_LOC_807/Y NOR2X1_LOC_527/Y 0.09fF
C58212 NOR2X1_LOC_498/Y INVX1_LOC_118/A 2.55fF
C58213 INVX1_LOC_251/Y INVX1_LOC_117/A 0.01fF
C58214 INVX1_LOC_232/A INVX1_LOC_20/A 0.07fF
C58215 NAND2X1_LOC_773/Y INVX1_LOC_251/A 0.08fF
C58216 NAND2X1_LOC_155/a_36_24# NOR2X1_LOC_45/B 0.00fF
C58217 NOR2X1_LOC_713/B NAND2X1_LOC_425/Y 0.03fF
C58218 INVX1_LOC_141/Y INVX1_LOC_264/A 0.01fF
C58219 INVX1_LOC_89/A NOR2X1_LOC_557/A 0.03fF
C58220 INVX1_LOC_161/A INVX1_LOC_12/A 0.07fF
C58221 GATE_579 INVX1_LOC_42/A 0.01fF
C58222 NOR2X1_LOC_639/B INVX1_LOC_296/A 0.02fF
C58223 INVX1_LOC_263/A INVX1_LOC_14/Y 0.10fF
C58224 INVX1_LOC_18/A NOR2X1_LOC_661/A 0.03fF
C58225 NOR2X1_LOC_793/Y INVX1_LOC_15/A 0.07fF
C58226 NOR2X1_LOC_352/Y INVX1_LOC_44/A 0.02fF
C58227 NOR2X1_LOC_360/Y NAND2X1_LOC_206/Y 0.04fF
C58228 NOR2X1_LOC_383/B NOR2X1_LOC_665/Y 0.07fF
C58229 NOR2X1_LOC_473/B INVX1_LOC_91/A 0.03fF
C58230 INVX1_LOC_23/A INVX1_LOC_58/Y 0.29fF
C58231 NOR2X1_LOC_700/Y NAND2X1_LOC_853/a_36_24# 0.00fF
C58232 NOR2X1_LOC_383/Y INVX1_LOC_20/A 0.00fF
C58233 NAND2X1_LOC_477/A INVX1_LOC_118/A 0.40fF
C58234 NOR2X1_LOC_160/B INVX1_LOC_290/Y 0.03fF
C58235 NOR2X1_LOC_641/B NAND2X1_LOC_74/B 0.03fF
C58236 NAND2X1_LOC_208/B INVX1_LOC_12/A 0.02fF
C58237 NOR2X1_LOC_391/A INVX1_LOC_76/A 0.07fF
C58238 NOR2X1_LOC_124/B NOR2X1_LOC_99/Y 0.05fF
C58239 INVX1_LOC_33/A NOR2X1_LOC_216/B 0.24fF
C58240 INVX1_LOC_30/Y INVX1_LOC_46/A 0.18fF
C58241 INVX1_LOC_1/A NAND2X1_LOC_452/Y 0.01fF
C58242 NAND2X1_LOC_325/Y NOR2X1_LOC_88/Y 4.07fF
C58243 NAND2X1_LOC_84/Y NOR2X1_LOC_814/A 0.05fF
C58244 NOR2X1_LOC_68/A INVX1_LOC_19/A 0.38fF
C58245 INVX1_LOC_53/A NOR2X1_LOC_434/A 0.03fF
C58246 INVX1_LOC_171/A NAND2X1_LOC_447/Y 0.01fF
C58247 NOR2X1_LOC_751/Y NAND2X1_LOC_74/B 0.11fF
C58248 NOR2X1_LOC_122/A NAND2X1_LOC_454/Y 0.02fF
C58249 NOR2X1_LOC_635/A INVX1_LOC_92/A 0.01fF
C58250 NOR2X1_LOC_591/Y INVX1_LOC_291/A 0.20fF
C58251 NAND2X1_LOC_784/A NOR2X1_LOC_109/Y 0.74fF
C58252 NOR2X1_LOC_772/B INVX1_LOC_29/Y 0.13fF
C58253 VDD NAND2X1_LOC_573/A 0.77fF
C58254 INVX1_LOC_1/A NOR2X1_LOC_307/Y 0.03fF
C58255 NOR2X1_LOC_722/Y INVX1_LOC_12/A 0.10fF
C58256 NOR2X1_LOC_446/A INVX1_LOC_4/A 0.02fF
C58257 NOR2X1_LOC_753/Y INVX1_LOC_84/A 0.36fF
C58258 INVX1_LOC_49/A INVX1_LOC_136/Y 0.01fF
C58259 NOR2X1_LOC_559/B NOR2X1_LOC_68/Y 0.05fF
C58260 INVX1_LOC_13/Y INVX1_LOC_29/Y 0.03fF
C58261 NOR2X1_LOC_322/Y INVX1_LOC_91/A 0.32fF
C58262 NOR2X1_LOC_323/Y NOR2X1_LOC_528/Y 0.09fF
C58263 INVX1_LOC_96/Y INVX1_LOC_92/A 0.07fF
C58264 NAND2X1_LOC_9/Y INVX1_LOC_50/Y 0.07fF
C58265 NAND2X1_LOC_364/A NOR2X1_LOC_114/Y 0.33fF
C58266 INVX1_LOC_276/A NOR2X1_LOC_88/Y 0.03fF
C58267 INVX1_LOC_75/A INVX1_LOC_199/A 0.14fF
C58268 INVX1_LOC_55/A INVX1_LOC_78/A 0.01fF
C58269 NAND2X1_LOC_840/B INVX1_LOC_92/A 0.01fF
C58270 NOR2X1_LOC_67/A NOR2X1_LOC_88/Y 0.42fF
C58271 INVX1_LOC_75/A INVX1_LOC_74/A 0.06fF
C58272 INVX1_LOC_41/A NAND2X1_LOC_63/Y 0.15fF
C58273 INVX1_LOC_256/A NOR2X1_LOC_843/B 0.05fF
C58274 NOR2X1_LOC_577/Y NOR2X1_LOC_89/A 0.17fF
C58275 INVX1_LOC_34/Y INVX1_LOC_3/A 0.02fF
C58276 INVX1_LOC_88/A INVX1_LOC_29/Y 0.09fF
C58277 NOR2X1_LOC_355/B INVX1_LOC_91/A 0.13fF
C58278 NAND2X1_LOC_347/B NOR2X1_LOC_717/A 0.00fF
C58279 INVX1_LOC_17/A INVX1_LOC_200/Y 0.01fF
C58280 NOR2X1_LOC_226/A NOR2X1_LOC_435/B 0.04fF
C58281 NOR2X1_LOC_15/Y INVX1_LOC_53/A 0.05fF
C58282 INVX1_LOC_24/A D_INPUT_5 0.01fF
C58283 INVX1_LOC_294/Y INVX1_LOC_29/A 0.00fF
C58284 NOR2X1_LOC_67/A INVX1_LOC_84/A 0.14fF
C58285 NOR2X1_LOC_798/A INVX1_LOC_50/Y 0.05fF
C58286 INVX1_LOC_34/A INVX1_LOC_12/A 16.26fF
C58287 NOR2X1_LOC_818/Y NAND2X1_LOC_818/a_36_24# 0.00fF
C58288 NOR2X1_LOC_814/Y INVX1_LOC_9/A 0.01fF
C58289 NOR2X1_LOC_383/a_36_216# NAND2X1_LOC_93/B 0.00fF
C58290 INVX1_LOC_62/Y NOR2X1_LOC_38/B 0.03fF
C58291 INVX1_LOC_21/A NOR2X1_LOC_186/Y 2.09fF
C58292 NOR2X1_LOC_45/B NAND2X1_LOC_623/B 0.00fF
C58293 NOR2X1_LOC_443/a_36_216# INVX1_LOC_57/A 0.00fF
C58294 INVX1_LOC_18/A NAND2X1_LOC_470/B 0.03fF
C58295 INVX1_LOC_30/A NOR2X1_LOC_449/A 0.11fF
C58296 NOR2X1_LOC_75/Y INVX1_LOC_23/A 0.00fF
C58297 NOR2X1_LOC_6/B NOR2X1_LOC_671/Y 0.06fF
C58298 INVX1_LOC_180/A INVX1_LOC_15/A 0.11fF
C58299 INVX1_LOC_31/A NOR2X1_LOC_654/A 0.35fF
C58300 NAND2X1_LOC_338/B NAND2X1_LOC_772/a_36_24# 0.00fF
C58301 NOR2X1_LOC_276/a_36_216# NAND2X1_LOC_454/Y 0.01fF
C58302 INVX1_LOC_285/Y VDD 1.61fF
C58303 INVX1_LOC_245/Y NOR2X1_LOC_598/B 0.02fF
C58304 INVX1_LOC_136/A NOR2X1_LOC_693/Y 0.07fF
C58305 INVX1_LOC_21/A NAND2X1_LOC_573/Y 0.51fF
C58306 NOR2X1_LOC_405/A NOR2X1_LOC_675/A 0.02fF
C58307 NOR2X1_LOC_520/B INVX1_LOC_15/A 0.07fF
C58308 NAND2X1_LOC_479/Y NAND2X1_LOC_475/Y 0.07fF
C58309 INVX1_LOC_136/A NAND2X1_LOC_288/B 0.05fF
C58310 INVX1_LOC_72/A NOR2X1_LOC_638/Y -0.03fF
C58311 NOR2X1_LOC_68/A INVX1_LOC_26/Y 0.18fF
C58312 NAND2X1_LOC_231/Y INVX1_LOC_12/A 0.02fF
C58313 INVX1_LOC_35/A NAND2X1_LOC_350/A 0.44fF
C58314 INVX1_LOC_64/A NOR2X1_LOC_446/A 0.01fF
C58315 NOR2X1_LOC_377/a_36_216# INVX1_LOC_37/A 0.00fF
C58316 NOR2X1_LOC_510/Y NOR2X1_LOC_361/B 0.14fF
C58317 INVX1_LOC_31/A INVX1_LOC_58/Y 0.01fF
C58318 INVX1_LOC_35/A NOR2X1_LOC_441/Y 0.11fF
C58319 NOR2X1_LOC_226/A INVX1_LOC_168/Y 0.03fF
C58320 NAND2X1_LOC_35/Y NOR2X1_LOC_134/Y 0.01fF
C58321 NAND2X1_LOC_358/Y NOR2X1_LOC_691/B 0.00fF
C58322 NAND2X1_LOC_149/Y INVX1_LOC_103/A 0.10fF
C58323 INVX1_LOC_65/A VDD 2.02fF
C58324 INPUT_1 NAND2X1_LOC_574/A 0.06fF
C58325 NOR2X1_LOC_137/A NOR2X1_LOC_814/A 0.24fF
C58326 INVX1_LOC_89/A NAND2X1_LOC_657/a_36_24# 0.00fF
C58327 INVX1_LOC_255/Y NAND2X1_LOC_207/Y 0.01fF
C58328 NOR2X1_LOC_15/Y NOR2X1_LOC_267/a_36_216# 0.00fF
C58329 NOR2X1_LOC_45/B INVX1_LOC_117/A 0.08fF
C58330 INVX1_LOC_22/A NOR2X1_LOC_89/A 0.17fF
C58331 NOR2X1_LOC_609/A INVX1_LOC_23/A 0.03fF
C58332 INVX1_LOC_316/A VDD -0.00fF
C58333 NAND2X1_LOC_348/A NOR2X1_LOC_78/Y 0.32fF
C58334 INVX1_LOC_276/A INVX1_LOC_15/A 0.50fF
C58335 INVX1_LOC_208/A INVX1_LOC_290/Y 1.14fF
C58336 INVX1_LOC_25/Y NAND2X1_LOC_254/Y 0.07fF
C58337 NOR2X1_LOC_810/A NOR2X1_LOC_777/B 0.03fF
C58338 VDD NOR2X1_LOC_137/B 0.08fF
C58339 NOR2X1_LOC_67/A INVX1_LOC_15/A 0.07fF
C58340 NOR2X1_LOC_82/A INVX1_LOC_48/Y 0.10fF
C58341 NOR2X1_LOC_763/Y INVX1_LOC_262/Y 0.02fF
C58342 NOR2X1_LOC_187/Y NAND2X1_LOC_192/B 0.00fF
C58343 NOR2X1_LOC_91/A NOR2X1_LOC_716/B 0.09fF
C58344 INVX1_LOC_255/Y NOR2X1_LOC_847/B 0.02fF
C58345 NOR2X1_LOC_443/Y NAND2X1_LOC_364/Y 0.02fF
C58346 INPUT_0 INVX1_LOC_307/A 0.08fF
C58347 NOR2X1_LOC_454/Y NOR2X1_LOC_160/B 0.28fF
C58348 INVX1_LOC_90/A NOR2X1_LOC_721/B 0.02fF
C58349 INVX1_LOC_91/A INVX1_LOC_193/A 0.01fF
C58350 INVX1_LOC_199/Y INVX1_LOC_117/A 0.08fF
C58351 VDD NAND2X1_LOC_267/B 0.01fF
C58352 INPUT_0 NOR2X1_LOC_445/B 0.07fF
C58353 NOR2X1_LOC_71/Y NAND2X1_LOC_74/B 0.10fF
C58354 NOR2X1_LOC_82/a_36_216# INVX1_LOC_306/Y 0.01fF
C58355 INVX1_LOC_230/Y NOR2X1_LOC_140/A 0.01fF
C58356 INVX1_LOC_21/A INVX1_LOC_170/A 0.00fF
C58357 NAND2X1_LOC_9/Y NOR2X1_LOC_559/B -0.01fF
C58358 NOR2X1_LOC_733/Y INVX1_LOC_92/A 0.00fF
C58359 NOR2X1_LOC_716/B INVX1_LOC_23/A 0.08fF
C58360 INVX1_LOC_232/A INVX1_LOC_4/A 0.07fF
C58361 NOR2X1_LOC_590/A INVX1_LOC_14/A 0.02fF
C58362 NOR2X1_LOC_356/A INVX1_LOC_29/A 0.16fF
C58363 NOR2X1_LOC_277/a_36_216# NOR2X1_LOC_716/B 0.01fF
C58364 NOR2X1_LOC_845/A INVX1_LOC_46/Y 0.15fF
C58365 NOR2X1_LOC_454/Y NAND2X1_LOC_195/Y -0.02fF
C58366 INVX1_LOC_36/A NAND2X1_LOC_326/A 0.13fF
C58367 INVX1_LOC_72/A NAND2X1_LOC_475/a_36_24# 0.01fF
C58368 INVX1_LOC_119/A INVX1_LOC_271/A 0.26fF
C58369 NAND2X1_LOC_39/a_36_24# INVX1_LOC_1/A 0.00fF
C58370 NAND2X1_LOC_860/A NOR2X1_LOC_392/B 0.10fF
C58371 INVX1_LOC_35/A NOR2X1_LOC_340/Y 0.09fF
C58372 NOR2X1_LOC_188/A INVX1_LOC_63/A 0.10fF
C58373 INVX1_LOC_147/A INVX1_LOC_19/A 0.01fF
C58374 INVX1_LOC_216/Y NOR2X1_LOC_514/A 0.02fF
C58375 INVX1_LOC_230/Y NOR2X1_LOC_530/Y 0.15fF
C58376 INVX1_LOC_269/A NOR2X1_LOC_169/B 0.04fF
C58377 INVX1_LOC_35/A NOR2X1_LOC_142/Y 0.17fF
C58378 INVX1_LOC_178/A NOR2X1_LOC_238/Y 0.01fF
C58379 INVX1_LOC_191/Y NOR2X1_LOC_654/A 0.00fF
C58380 NAND2X1_LOC_9/Y NOR2X1_LOC_6/B 0.16fF
C58381 NOR2X1_LOC_548/B INVX1_LOC_63/A 0.10fF
C58382 NOR2X1_LOC_92/Y INVX1_LOC_61/A 0.04fF
C58383 INVX1_LOC_98/Y INVX1_LOC_23/A 0.01fF
C58384 NOR2X1_LOC_2/Y NOR2X1_LOC_11/Y 0.77fF
C58385 INVX1_LOC_1/Y INVX1_LOC_116/Y 0.03fF
C58386 NAND2X1_LOC_733/Y INVX1_LOC_161/A 0.05fF
C58387 INVX1_LOC_75/A NOR2X1_LOC_509/a_36_216# 0.00fF
C58388 INVX1_LOC_21/A INVX1_LOC_132/A 0.07fF
C58389 INVX1_LOC_11/A NOR2X1_LOC_274/B 0.04fF
C58390 NOR2X1_LOC_74/A INVX1_LOC_29/A 0.48fF
C58391 INVX1_LOC_12/Y INVX1_LOC_9/A 0.10fF
C58392 INVX1_LOC_8/A INVX1_LOC_306/Y 0.18fF
C58393 INPUT_0 INVX1_LOC_12/A 0.24fF
C58394 INVX1_LOC_41/A INVX1_LOC_39/A 0.03fF
C58395 NAND2X1_LOC_190/Y NOR2X1_LOC_596/A 0.07fF
C58396 INVX1_LOC_256/A INVX1_LOC_18/A 0.07fF
C58397 INPUT_0 NOR2X1_LOC_519/Y 0.05fF
C58398 NOR2X1_LOC_647/Y NOR2X1_LOC_647/B -0.00fF
C58399 NOR2X1_LOC_9/Y INVX1_LOC_29/A 0.30fF
C58400 NOR2X1_LOC_68/A INVX1_LOC_161/Y 0.07fF
C58401 NAND2X1_LOC_290/a_36_24# INVX1_LOC_53/A 0.00fF
C58402 INVX1_LOC_35/A NOR2X1_LOC_655/B 0.03fF
C58403 INVX1_LOC_272/Y INVX1_LOC_246/Y 0.06fF
C58404 NOR2X1_LOC_689/Y NAND2X1_LOC_727/Y 0.01fF
C58405 INVX1_LOC_2/A NAND2X1_LOC_35/Y 0.07fF
C58406 INVX1_LOC_36/A NAND2X1_LOC_104/a_36_24# 0.00fF
C58407 NOR2X1_LOC_798/A NOR2X1_LOC_6/B 0.03fF
C58408 INVX1_LOC_21/A INVX1_LOC_225/A 0.08fF
C58409 NOR2X1_LOC_815/Y NOR2X1_LOC_92/Y 0.00fF
C58410 INVX1_LOC_25/A INVX1_LOC_1/Y 0.07fF
C58411 INVX1_LOC_284/Y INVX1_LOC_72/A 0.03fF
C58412 INVX1_LOC_272/Y NAND2X1_LOC_802/A 0.01fF
C58413 INVX1_LOC_232/Y NOR2X1_LOC_663/A 0.05fF
C58414 NOR2X1_LOC_349/A NOR2X1_LOC_509/A 0.01fF
C58415 NOR2X1_LOC_614/a_36_216# NOR2X1_LOC_614/Y 0.00fF
C58416 NOR2X1_LOC_624/A INVX1_LOC_24/Y 0.05fF
C58417 INVX1_LOC_117/A NOR2X1_LOC_862/B 0.11fF
C58418 INVX1_LOC_11/A NOR2X1_LOC_577/Y 0.07fF
C58419 NAND2X1_LOC_199/B INVX1_LOC_107/A 0.06fF
C58420 INVX1_LOC_17/A NAND2X1_LOC_361/Y 0.07fF
C58421 NOR2X1_LOC_295/Y NOR2X1_LOC_468/Y 0.02fF
C58422 NOR2X1_LOC_389/A NOR2X1_LOC_596/A 0.03fF
C58423 INVX1_LOC_255/Y NOR2X1_LOC_660/Y 0.02fF
C58424 INVX1_LOC_21/A NOR2X1_LOC_209/Y 0.06fF
C58425 NOR2X1_LOC_186/Y INVX1_LOC_248/A 0.08fF
C58426 INVX1_LOC_90/A NAND2X1_LOC_286/B 1.38fF
C58427 NOR2X1_LOC_245/a_36_216# INVX1_LOC_57/A 0.00fF
C58428 INVX1_LOC_36/A NAND2X1_LOC_481/a_36_24# 0.00fF
C58429 NOR2X1_LOC_160/B INVX1_LOC_77/A 1.70fF
C58430 NOR2X1_LOC_717/B INVX1_LOC_23/A 0.08fF
C58431 GATE_741 NAND2X1_LOC_733/B 0.01fF
C58432 NOR2X1_LOC_388/Y NOR2X1_LOC_457/A 0.03fF
C58433 NOR2X1_LOC_721/Y INVX1_LOC_4/Y 0.02fF
C58434 INVX1_LOC_55/A INVX1_LOC_113/Y 0.01fF
C58435 INVX1_LOC_268/A INVX1_LOC_5/A 0.01fF
C58436 INVX1_LOC_278/Y NAND2X1_LOC_794/B 0.09fF
C58437 NOR2X1_LOC_756/Y NAND2X1_LOC_99/A 0.00fF
C58438 INVX1_LOC_65/Y INVX1_LOC_57/A 0.04fF
C58439 NOR2X1_LOC_113/A NOR2X1_LOC_114/Y 0.00fF
C58440 NOR2X1_LOC_667/A NAND2X1_LOC_573/Y 0.03fF
C58441 NAND2X1_LOC_787/A INVX1_LOC_135/A 0.01fF
C58442 NOR2X1_LOC_91/A NOR2X1_LOC_503/A 0.01fF
C58443 NOR2X1_LOC_598/B D_INPUT_0 0.29fF
C58444 INVX1_LOC_88/A NOR2X1_LOC_361/Y 0.01fF
C58445 NOR2X1_LOC_405/A NOR2X1_LOC_114/Y 0.02fF
C58446 NAND2X1_LOC_731/Y INVX1_LOC_72/A 0.09fF
C58447 INVX1_LOC_136/A INVX1_LOC_45/Y 0.00fF
C58448 INVX1_LOC_248/A NAND2X1_LOC_573/Y 0.76fF
C58449 NOR2X1_LOC_178/Y NOR2X1_LOC_391/A 0.03fF
C58450 INVX1_LOC_11/A NOR2X1_LOC_348/B 0.01fF
C58451 NOR2X1_LOC_716/B INVX1_LOC_31/A 0.26fF
C58452 NAND2X1_LOC_363/B INVX1_LOC_135/A 0.07fF
C58453 INVX1_LOC_51/A D_INPUT_0 0.03fF
C58454 NOR2X1_LOC_45/B INVX1_LOC_3/Y 0.02fF
C58455 INVX1_LOC_35/A NOR2X1_LOC_99/B 0.08fF
C58456 NOR2X1_LOC_483/B NOR2X1_LOC_254/Y 0.07fF
C58457 INVX1_LOC_64/A NOR2X1_LOC_366/Y 0.02fF
C58458 NAND2X1_LOC_807/Y NOR2X1_LOC_654/A 0.10fF
C58459 NOR2X1_LOC_15/Y NOR2X1_LOC_78/B 0.10fF
C58460 NOR2X1_LOC_309/Y NAND2X1_LOC_807/A 0.03fF
C58461 INVX1_LOC_57/Y NOR2X1_LOC_237/a_36_216# 0.00fF
C58462 INVX1_LOC_298/Y NOR2X1_LOC_74/A 0.29fF
C58463 NOR2X1_LOC_667/A NAND2X1_LOC_724/A 0.15fF
C58464 NAND2X1_LOC_860/A INVX1_LOC_90/A 0.03fF
C58465 NOR2X1_LOC_82/A NOR2X1_LOC_84/Y 0.43fF
C58466 INVX1_LOC_24/A NOR2X1_LOC_360/Y 0.03fF
C58467 NAND2X1_LOC_53/Y INVX1_LOC_266/Y 0.11fF
C58468 NOR2X1_LOC_816/A NOR2X1_LOC_574/A 0.27fF
C58469 VDD NAND2X1_LOC_81/B 0.25fF
C58470 INVX1_LOC_34/A NAND2X1_LOC_733/Y 0.03fF
C58471 INVX1_LOC_136/A NAND2X1_LOC_740/A 0.02fF
C58472 INVX1_LOC_248/A NAND2X1_LOC_724/A 0.11fF
C58473 NOR2X1_LOC_389/B NOR2X1_LOC_15/a_36_216# 0.01fF
C58474 INVX1_LOC_269/A INVX1_LOC_179/Y 0.02fF
C58475 INVX1_LOC_166/A NAND2X1_LOC_462/a_36_24# 0.01fF
C58476 INVX1_LOC_177/Y NOR2X1_LOC_106/Y 0.20fF
C58477 NOR2X1_LOC_337/Y INVX1_LOC_4/Y 0.21fF
C58478 NOR2X1_LOC_134/Y NAND2X1_LOC_465/Y 0.03fF
C58479 NAND2X1_LOC_582/a_36_24# INVX1_LOC_174/A 0.00fF
C58480 NAND2X1_LOC_190/Y NOR2X1_LOC_220/A 0.01fF
C58481 NOR2X1_LOC_831/B NOR2X1_LOC_743/Y 0.24fF
C58482 NOR2X1_LOC_211/a_36_216# NOR2X1_LOC_389/B 0.00fF
C58483 NOR2X1_LOC_82/A INVX1_LOC_216/A 0.02fF
C58484 INVX1_LOC_223/A INVX1_LOC_155/A 0.08fF
C58485 INVX1_LOC_224/A NOR2X1_LOC_346/B 0.05fF
C58486 INVX1_LOC_124/A NOR2X1_LOC_160/B 0.05fF
C58487 NOR2X1_LOC_593/Y NOR2X1_LOC_274/B 0.19fF
C58488 INVX1_LOC_38/A NOR2X1_LOC_721/B 0.03fF
C58489 NOR2X1_LOC_363/Y INVX1_LOC_272/A 0.06fF
C58490 NOR2X1_LOC_78/A NOR2X1_LOC_248/A 0.01fF
C58491 INVX1_LOC_290/Y NAND2X1_LOC_211/Y 0.20fF
C58492 INVX1_LOC_1/A INVX1_LOC_1/Y 0.17fF
C58493 INVX1_LOC_14/A NOR2X1_LOC_82/Y 0.39fF
C58494 NAND2X1_LOC_35/Y INPUT_1 0.63fF
C58495 NOR2X1_LOC_92/Y NAND2X1_LOC_735/B 0.03fF
C58496 NAND2X1_LOC_214/B INVX1_LOC_89/A 0.14fF
C58497 NOR2X1_LOC_151/Y INVX1_LOC_23/A 0.09fF
C58498 INVX1_LOC_152/A NOR2X1_LOC_243/B 0.20fF
C58499 NOR2X1_LOC_433/A NOR2X1_LOC_351/a_36_216# 0.01fF
C58500 INVX1_LOC_269/A NOR2X1_LOC_719/A 0.10fF
C58501 NOR2X1_LOC_590/A INVX1_LOC_111/Y 0.02fF
C58502 INVX1_LOC_34/A INVX1_LOC_217/A 0.11fF
C58503 INVX1_LOC_103/A INVX1_LOC_16/A 0.10fF
C58504 INVX1_LOC_200/A NAND2X1_LOC_858/a_36_24# 0.00fF
C58505 NAND2X1_LOC_447/Y INVX1_LOC_4/A 0.13fF
C58506 INVX1_LOC_224/A INVX1_LOC_22/A 0.00fF
C58507 NOR2X1_LOC_15/Y NAND2X1_LOC_392/Y 0.00fF
C58508 NAND2X1_LOC_303/Y NAND2X1_LOC_854/B 0.02fF
C58509 NAND2X1_LOC_391/Y NOR2X1_LOC_76/A 0.12fF
C58510 INVX1_LOC_36/A NOR2X1_LOC_87/B 0.05fF
C58511 INVX1_LOC_37/A NAND2X1_LOC_430/B 0.09fF
C58512 INVX1_LOC_11/A INVX1_LOC_22/A 6.67fF
C58513 NOR2X1_LOC_15/Y NOR2X1_LOC_459/A 0.23fF
C58514 INVX1_LOC_207/A INVX1_LOC_24/A 0.02fF
C58515 INVX1_LOC_27/A INVX1_LOC_89/A 2.07fF
C58516 INVX1_LOC_225/Y NOR2X1_LOC_500/Y -0.01fF
C58517 NAND2X1_LOC_2/a_36_24# INVX1_LOC_53/A 0.00fF
C58518 INVX1_LOC_269/A NOR2X1_LOC_561/Y 0.22fF
C58519 NOR2X1_LOC_500/A INVX1_LOC_33/A 0.00fF
C58520 INVX1_LOC_33/A NOR2X1_LOC_303/Y 0.03fF
C58521 NOR2X1_LOC_361/B NAND2X1_LOC_573/A 0.51fF
C58522 NOR2X1_LOC_433/A NOR2X1_LOC_577/Y 0.09fF
C58523 INVX1_LOC_48/Y NOR2X1_LOC_132/a_36_216# 0.00fF
C58524 NOR2X1_LOC_160/B NOR2X1_LOC_687/Y 0.03fF
C58525 INVX1_LOC_292/A INVX1_LOC_16/A 0.03fF
C58526 INVX1_LOC_27/A NAND2X1_LOC_508/A 0.01fF
C58527 NOR2X1_LOC_593/Y NOR2X1_LOC_577/Y 0.07fF
C58528 NOR2X1_LOC_355/A INVX1_LOC_88/A 0.03fF
C58529 VDD INVX1_LOC_4/Y 1.31fF
C58530 INVX1_LOC_49/Y INVX1_LOC_92/A 0.03fF
C58531 NOR2X1_LOC_527/Y NOR2X1_LOC_109/Y 0.04fF
C58532 NOR2X1_LOC_383/Y INVX1_LOC_43/Y 0.26fF
C58533 NOR2X1_LOC_106/Y INVX1_LOC_104/A 0.19fF
C58534 INVX1_LOC_34/A NAND2X1_LOC_787/B 1.05fF
C58535 INVX1_LOC_58/A NOR2X1_LOC_45/B 0.19fF
C58536 INVX1_LOC_143/A NOR2X1_LOC_360/Y 0.07fF
C58537 NOR2X1_LOC_517/Y NAND2X1_LOC_852/Y 0.10fF
C58538 NOR2X1_LOC_197/a_36_216# NOR2X1_LOC_748/A 0.01fF
C58539 INVX1_LOC_90/A NAND2X1_LOC_537/Y 0.03fF
C58540 INVX1_LOC_2/A INVX1_LOC_94/A 0.07fF
C58541 INVX1_LOC_30/A NAND2X1_LOC_479/Y 0.02fF
C58542 NOR2X1_LOC_52/B NOR2X1_LOC_577/Y 0.47fF
C58543 INVX1_LOC_25/A INVX1_LOC_93/Y 0.07fF
C58544 NOR2X1_LOC_717/B NAND2X1_LOC_179/a_36_24# 0.00fF
C58545 NOR2X1_LOC_593/Y NOR2X1_LOC_348/B 0.03fF
C58546 NOR2X1_LOC_729/A INVX1_LOC_15/A 0.08fF
C58547 INVX1_LOC_226/Y INVX1_LOC_72/Y 0.03fF
C58548 INVX1_LOC_103/A INVX1_LOC_28/A 0.07fF
C58549 NOR2X1_LOC_243/B INVX1_LOC_29/A 0.07fF
C58550 INVX1_LOC_1/A NOR2X1_LOC_742/A 0.10fF
C58551 NOR2X1_LOC_590/A NOR2X1_LOC_137/A 0.12fF
C58552 NAND2X1_LOC_9/Y NOR2X1_LOC_124/A 0.02fF
C58553 NOR2X1_LOC_6/B NOR2X1_LOC_140/a_36_216# 0.01fF
C58554 INVX1_LOC_304/Y INVX1_LOC_34/A 0.08fF
C58555 NAND2X1_LOC_198/B INVX1_LOC_56/Y 0.10fF
C58556 NAND2X1_LOC_564/B NOR2X1_LOC_91/Y 0.10fF
C58557 INVX1_LOC_54/Y INVX1_LOC_33/A 0.02fF
C58558 INVX1_LOC_233/A NOR2X1_LOC_124/A 0.01fF
C58559 NOR2X1_LOC_246/A INVX1_LOC_141/Y 0.02fF
C58560 INVX1_LOC_135/A INVX1_LOC_30/A 0.01fF
C58561 INVX1_LOC_53/A NOR2X1_LOC_137/a_36_216# 0.00fF
C58562 INVX1_LOC_314/Y INVX1_LOC_25/Y 0.03fF
C58563 NOR2X1_LOC_500/A NAND2X1_LOC_754/a_36_24# 0.01fF
C58564 NOR2X1_LOC_828/B NOR2X1_LOC_307/A 0.03fF
C58565 INVX1_LOC_208/A INVX1_LOC_77/A 0.08fF
C58566 NOR2X1_LOC_735/a_36_216# NOR2X1_LOC_665/A 0.02fF
C58567 INVX1_LOC_292/A INVX1_LOC_28/A 0.03fF
C58568 NOR2X1_LOC_246/A INVX1_LOC_312/Y 0.00fF
C58569 INVX1_LOC_80/Y NAND2X1_LOC_141/A 0.20fF
C58570 INVX1_LOC_72/A NOR2X1_LOC_525/Y 0.01fF
C58571 NOR2X1_LOC_516/B INVX1_LOC_77/A 0.30fF
C58572 INVX1_LOC_295/A INVX1_LOC_30/A 0.04fF
C58573 NOR2X1_LOC_252/Y NOR2X1_LOC_495/Y 0.10fF
C58574 INVX1_LOC_136/A NOR2X1_LOC_71/Y 0.07fF
C58575 NOR2X1_LOC_433/A INVX1_LOC_22/A 0.26fF
C58576 NAND2X1_LOC_717/Y INVX1_LOC_240/A 0.03fF
C58577 INVX1_LOC_228/Y INPUT_0 0.26fF
C58578 NOR2X1_LOC_272/Y NOR2X1_LOC_139/Y 0.10fF
C58579 INVX1_LOC_225/A NOR2X1_LOC_667/A -0.04fF
C58580 NOR2X1_LOC_68/A INVX1_LOC_62/A 0.18fF
C58581 INVX1_LOC_200/A INPUT_0 0.13fF
C58582 NOR2X1_LOC_790/B INVX1_LOC_37/A 0.03fF
C58583 INVX1_LOC_102/A NOR2X1_LOC_662/A 0.02fF
C58584 NOR2X1_LOC_89/A INVX1_LOC_186/Y 0.07fF
C58585 NOR2X1_LOC_599/Y NOR2X1_LOC_597/Y 0.00fF
C58586 NOR2X1_LOC_277/a_36_216# NAND2X1_LOC_633/Y 0.00fF
C58587 NOR2X1_LOC_613/Y NAND2X1_LOC_623/B 0.06fF
C58588 NOR2X1_LOC_593/Y INVX1_LOC_22/A 0.10fF
C58589 INVX1_LOC_21/A NAND2X1_LOC_642/Y 0.10fF
C58590 INVX1_LOC_58/A INVX1_LOC_281/A 0.01fF
C58591 INVX1_LOC_126/Y NAND2X1_LOC_793/Y 0.14fF
C58592 NOR2X1_LOC_180/B NOR2X1_LOC_703/B 0.00fF
C58593 INVX1_LOC_233/Y VDD 1.55fF
C58594 NOR2X1_LOC_490/Y INVX1_LOC_30/A 0.49fF
C58595 INVX1_LOC_136/A NOR2X1_LOC_644/A 0.08fF
C58596 NOR2X1_LOC_67/A NOR2X1_LOC_63/a_36_216# 0.00fF
C58597 NAND2X1_LOC_802/A INVX1_LOC_10/A 0.00fF
C58598 NOR2X1_LOC_716/B NAND2X1_LOC_859/Y 0.01fF
C58599 INVX1_LOC_83/A NOR2X1_LOC_860/B 0.07fF
C58600 NOR2X1_LOC_78/B INVX1_LOC_96/Y 0.07fF
C58601 NOR2X1_LOC_160/B NAND2X1_LOC_832/Y 0.02fF
C58602 NOR2X1_LOC_272/Y NAND2X1_LOC_468/B 0.03fF
C58603 NAND2X1_LOC_370/a_36_24# NAND2X1_LOC_721/A 0.01fF
C58604 INVX1_LOC_151/A INVX1_LOC_22/A 0.01fF
C58605 NAND2X1_LOC_727/Y NAND2X1_LOC_308/Y 0.05fF
C58606 INVX1_LOC_240/A INVX1_LOC_16/A 0.12fF
C58607 NAND2X1_LOC_733/Y INPUT_0 0.03fF
C58608 NOR2X1_LOC_80/Y NAND2X1_LOC_572/B 0.04fF
C58609 NOR2X1_LOC_52/B INVX1_LOC_22/A 0.42fF
C58610 INVX1_LOC_2/A NOR2X1_LOC_136/Y 0.14fF
C58611 NOR2X1_LOC_500/Y INVX1_LOC_266/Y 0.08fF
C58612 NAND2X1_LOC_796/B INVX1_LOC_20/A 0.02fF
C58613 NOR2X1_LOC_401/Y NAND2X1_LOC_181/Y 0.02fF
C58614 INVX1_LOC_1/A INVX1_LOC_93/Y 0.15fF
C58615 NAND2X1_LOC_838/Y INVX1_LOC_22/A 0.03fF
C58616 NOR2X1_LOC_605/a_36_216# NAND2X1_LOC_357/B 0.00fF
C58617 NOR2X1_LOC_547/B INVX1_LOC_226/A 0.00fF
C58618 NAND2X1_LOC_778/Y INVX1_LOC_46/A 0.03fF
C58619 NOR2X1_LOC_824/A NAND2X1_LOC_244/A 0.01fF
C58620 INVX1_LOC_48/Y INVX1_LOC_59/Y 0.05fF
C58621 INVX1_LOC_10/A NAND2X1_LOC_811/Y 0.03fF
C58622 INVX1_LOC_178/A NOR2X1_LOC_305/Y 0.10fF
C58623 NOR2X1_LOC_590/A INVX1_LOC_48/A 0.01fF
C58624 INVX1_LOC_134/A INVX1_LOC_160/A 0.02fF
C58625 NOR2X1_LOC_15/Y NOR2X1_LOC_164/Y 0.00fF
C58626 NAND2X1_LOC_67/a_36_24# INVX1_LOC_76/A 0.01fF
C58627 INVX1_LOC_215/Y NOR2X1_LOC_45/B 0.07fF
C58628 NOR2X1_LOC_457/A NOR2X1_LOC_552/A 0.09fF
C58629 INVX1_LOC_247/Y NOR2X1_LOC_74/A 0.03fF
C58630 INVX1_LOC_24/A NOR2X1_LOC_567/B 0.03fF
C58631 NOR2X1_LOC_716/B NAND2X1_LOC_866/B 0.00fF
C58632 NAND2X1_LOC_660/Y NAND2X1_LOC_660/A 0.05fF
C58633 NOR2X1_LOC_552/Y NOR2X1_LOC_500/B 0.03fF
C58634 INVX1_LOC_10/A NOR2X1_LOC_821/Y 0.06fF
C58635 NAND2X1_LOC_550/a_36_24# NAND2X1_LOC_338/B 0.00fF
C58636 NOR2X1_LOC_533/A INVX1_LOC_16/A 0.05fF
C58637 NOR2X1_LOC_703/B NOR2X1_LOC_569/A 0.01fF
C58638 INVX1_LOC_69/Y NOR2X1_LOC_532/a_36_216# 0.01fF
C58639 INVX1_LOC_217/A INPUT_0 0.03fF
C58640 NOR2X1_LOC_411/A NOR2X1_LOC_629/Y 0.00fF
C58641 NAND2X1_LOC_223/A NOR2X1_LOC_721/B 0.03fF
C58642 INVX1_LOC_269/A INVX1_LOC_76/A 0.10fF
C58643 NOR2X1_LOC_647/A NOR2X1_LOC_649/B 0.02fF
C58644 INVX1_LOC_1/A INVX1_LOC_139/A 0.04fF
C58645 NOR2X1_LOC_794/A INVX1_LOC_30/A 0.08fF
C58646 NOR2X1_LOC_15/Y INVX1_LOC_46/A 0.33fF
C58647 NAND2X1_LOC_35/Y INVX1_LOC_118/A 1.54fF
C58648 NOR2X1_LOC_147/B INVX1_LOC_85/Y 0.02fF
C58649 INVX1_LOC_90/A NOR2X1_LOC_486/B 0.00fF
C58650 INVX1_LOC_14/A NAND2X1_LOC_650/B 0.03fF
C58651 INVX1_LOC_227/A INVX1_LOC_111/Y 0.01fF
C58652 INVX1_LOC_69/Y INVX1_LOC_18/A 0.02fF
C58653 INVX1_LOC_314/Y INVX1_LOC_75/A 0.03fF
C58654 NOR2X1_LOC_220/A NOR2X1_LOC_548/Y 0.10fF
C58655 INVX1_LOC_57/A INVX1_LOC_123/Y 0.06fF
C58656 NOR2X1_LOC_383/B INVX1_LOC_285/A 0.07fF
C58657 INVX1_LOC_16/Y INVX1_LOC_293/Y 0.13fF
C58658 INVX1_LOC_90/A NOR2X1_LOC_64/a_36_216# 0.02fF
C58659 NOR2X1_LOC_94/a_36_216# INVX1_LOC_316/Y 0.00fF
C58660 NOR2X1_LOC_205/Y NOR2X1_LOC_69/a_36_216# 0.00fF
C58661 NOR2X1_LOC_205/Y VDD 0.57fF
C58662 D_INPUT_0 NAND2X1_LOC_660/A 0.15fF
C58663 NOR2X1_LOC_234/Y INPUT_1 -0.00fF
C58664 INVX1_LOC_152/Y NAND2X1_LOC_60/a_36_24# 0.01fF
C58665 NOR2X1_LOC_36/A NOR2X1_LOC_11/Y 0.87fF
C58666 NOR2X1_LOC_666/A NAND2X1_LOC_472/Y 0.04fF
C58667 INVX1_LOC_26/A NAND2X1_LOC_773/B 0.05fF
C58668 NOR2X1_LOC_383/B NOR2X1_LOC_814/A 0.03fF
C58669 NOR2X1_LOC_552/A INVX1_LOC_30/A 0.10fF
C58670 NOR2X1_LOC_389/A NAND2X1_LOC_469/B 0.10fF
C58671 INVX1_LOC_292/A NOR2X1_LOC_35/Y 0.10fF
C58672 INVX1_LOC_49/A INVX1_LOC_144/A 0.08fF
C58673 INVX1_LOC_28/A INVX1_LOC_240/A 0.44fF
C58674 NAND2X1_LOC_112/Y NOR2X1_LOC_589/A 0.03fF
C58675 INVX1_LOC_83/A INVX1_LOC_226/A 0.03fF
C58676 NOR2X1_LOC_816/A NOR2X1_LOC_305/Y 0.07fF
C58677 NAND2X1_LOC_541/a_36_24# INVX1_LOC_123/Y 0.00fF
C58678 INVX1_LOC_298/A NAND2X1_LOC_93/B 0.04fF
C58679 NOR2X1_LOC_510/a_36_216# INVX1_LOC_144/Y 0.00fF
C58680 INVX1_LOC_209/Y NOR2X1_LOC_313/Y 0.01fF
C58681 D_INPUT_0 NAND2X1_LOC_528/a_36_24# 0.00fF
C58682 NOR2X1_LOC_419/Y INVX1_LOC_6/A 0.09fF
C58683 NAND2X1_LOC_714/B INVX1_LOC_54/A 0.01fF
C58684 NOR2X1_LOC_785/A INVX1_LOC_37/A 0.01fF
C58685 INVX1_LOC_298/A NAND2X1_LOC_425/Y 0.02fF
C58686 NAND2X1_LOC_537/Y INVX1_LOC_38/A 0.07fF
C58687 NOR2X1_LOC_39/Y NAND2X1_LOC_74/B 0.01fF
C58688 NOR2X1_LOC_99/B NOR2X1_LOC_121/A 0.05fF
C58689 NOR2X1_LOC_716/B INVX1_LOC_6/A 0.14fF
C58690 NOR2X1_LOC_416/A NAND2X1_LOC_219/B 0.03fF
C58691 NOR2X1_LOC_299/Y NAND2X1_LOC_735/B 0.03fF
C58692 NOR2X1_LOC_725/A NOR2X1_LOC_713/B 0.15fF
C58693 INVX1_LOC_33/A NOR2X1_LOC_354/Y 0.01fF
C58694 NAND2X1_LOC_793/Y NOR2X1_LOC_536/A 0.05fF
C58695 NAND2X1_LOC_725/A INVX1_LOC_5/Y 0.05fF
C58696 NOR2X1_LOC_309/Y NOR2X1_LOC_527/Y 0.02fF
C58697 INVX1_LOC_8/A NOR2X1_LOC_9/Y 0.00fF
C58698 NAND2X1_LOC_74/B NAND2X1_LOC_205/A 0.01fF
C58699 NOR2X1_LOC_778/B NOR2X1_LOC_439/B 0.00fF
C58700 INVX1_LOC_56/Y NOR2X1_LOC_76/a_36_216# 0.00fF
C58701 INVX1_LOC_53/A INVX1_LOC_49/Y 0.03fF
C58702 NOR2X1_LOC_716/B NOR2X1_LOC_10/a_36_216# 0.01fF
C58703 NOR2X1_LOC_723/Y VDD 0.00fF
C58704 NAND2X1_LOC_374/Y NOR2X1_LOC_322/Y 0.02fF
C58705 INVX1_LOC_102/A INVX1_LOC_57/A 0.08fF
C58706 NOR2X1_LOC_292/Y NOR2X1_LOC_709/A 0.02fF
C58707 NAND2X1_LOC_833/Y INVX1_LOC_91/A 0.07fF
C58708 INVX1_LOC_2/A INVX1_LOC_144/A 0.10fF
C58709 INVX1_LOC_227/A NOR2X1_LOC_137/A 0.03fF
C58710 NOR2X1_LOC_778/B INVX1_LOC_75/A 0.06fF
C58711 NOR2X1_LOC_486/Y NOR2X1_LOC_303/Y 0.03fF
C58712 INVX1_LOC_78/A NOR2X1_LOC_681/a_36_216# 0.00fF
C58713 INVX1_LOC_26/A NOR2X1_LOC_393/Y 0.01fF
C58714 INVX1_LOC_89/A INVX1_LOC_234/A 0.07fF
C58715 NOR2X1_LOC_160/B INVX1_LOC_9/A 10.77fF
C58716 NAND2X1_LOC_338/B NOR2X1_LOC_97/A 0.03fF
C58717 INVX1_LOC_285/Y INVX1_LOC_177/A 0.05fF
C58718 INVX1_LOC_53/A INVX1_LOC_99/A 0.47fF
C58719 NOR2X1_LOC_384/Y NAND2X1_LOC_721/A 0.04fF
C58720 NOR2X1_LOC_226/A INVX1_LOC_144/A 0.08fF
C58721 NOR2X1_LOC_209/Y INVX1_LOC_311/A 0.21fF
C58722 INVX1_LOC_235/Y NAND2X1_LOC_659/A 0.34fF
C58723 NAND2X1_LOC_323/B NOR2X1_LOC_97/A 0.05fF
C58724 NOR2X1_LOC_226/A NOR2X1_LOC_83/Y 0.01fF
C58725 INVX1_LOC_98/Y INVX1_LOC_6/A 0.36fF
C58726 NAND2X1_LOC_640/Y INVX1_LOC_304/A 0.01fF
C58727 NOR2X1_LOC_350/A INVX1_LOC_176/A 0.00fF
C58728 NOR2X1_LOC_78/B NOR2X1_LOC_733/Y 0.01fF
C58729 INVX1_LOC_116/Y INVX1_LOC_87/A 0.00fF
C58730 NOR2X1_LOC_560/a_36_216# NAND2X1_LOC_206/Y 0.01fF
C58731 NAND2X1_LOC_352/B NOR2X1_LOC_743/Y 0.57fF
C58732 NOR2X1_LOC_67/A INVX1_LOC_123/A 0.01fF
C58733 NAND2X1_LOC_326/A INVX1_LOC_63/A 0.03fF
C58734 INVX1_LOC_1/Y NOR2X1_LOC_188/A 0.10fF
C58735 INVX1_LOC_225/Y NOR2X1_LOC_445/B 0.10fF
C58736 NOR2X1_LOC_219/B NOR2X1_LOC_357/Y 0.04fF
C58737 INVX1_LOC_1/Y NOR2X1_LOC_548/B 0.05fF
C58738 INVX1_LOC_177/A INVX1_LOC_65/A 0.03fF
C58739 NOR2X1_LOC_607/A NOR2X1_LOC_536/A 0.02fF
C58740 INVX1_LOC_194/A NAND2X1_LOC_659/B 0.37fF
C58741 NOR2X1_LOC_387/A NAND2X1_LOC_857/a_36_24# 0.00fF
C58742 INVX1_LOC_89/A NOR2X1_LOC_19/B 0.12fF
C58743 NOR2X1_LOC_344/A INVX1_LOC_37/A 0.02fF
C58744 INVX1_LOC_201/Y D_GATE_479 0.01fF
C58745 INVX1_LOC_45/A INVX1_LOC_180/Y 0.09fF
C58746 INVX1_LOC_201/Y D_INPUT_3 0.07fF
C58747 NOR2X1_LOC_84/Y INVX1_LOC_59/Y 0.01fF
C58748 INVX1_LOC_177/A NOR2X1_LOC_137/B 0.01fF
C58749 NOR2X1_LOC_843/A VDD 0.22fF
C58750 INVX1_LOC_112/A NOR2X1_LOC_84/Y 0.16fF
C58751 NOR2X1_LOC_486/Y NOR2X1_LOC_353/Y 0.00fF
C58752 INVX1_LOC_68/A INVX1_LOC_15/A 0.01fF
C58753 NOR2X1_LOC_92/Y NOR2X1_LOC_831/Y 0.06fF
C58754 NOR2X1_LOC_667/A NAND2X1_LOC_642/Y 2.14fF
C58755 INVX1_LOC_136/A NAND2X1_LOC_243/Y 0.02fF
C58756 NOR2X1_LOC_78/A NOR2X1_LOC_131/Y 0.04fF
C58757 INVX1_LOC_248/A NAND2X1_LOC_642/Y 0.06fF
C58758 NOR2X1_LOC_722/Y INVX1_LOC_92/A 0.00fF
C58759 INVX1_LOC_11/A INVX1_LOC_186/Y 0.07fF
C58760 NOR2X1_LOC_273/Y INVX1_LOC_54/A 0.83fF
C58761 NOR2X1_LOC_361/B NAND2X1_LOC_81/B 0.07fF
C58762 NAND2X1_LOC_357/B INVX1_LOC_37/A 0.07fF
C58763 NOR2X1_LOC_773/Y INVX1_LOC_95/Y 0.13fF
C58764 NOR2X1_LOC_589/A INVX1_LOC_98/A 0.01fF
C58765 NOR2X1_LOC_759/Y INVX1_LOC_54/A 0.03fF
C58766 NAND2X1_LOC_714/B NOR2X1_LOC_48/B 0.07fF
C58767 INVX1_LOC_202/A INVX1_LOC_54/A 0.07fF
C58768 NOR2X1_LOC_781/A INVX1_LOC_91/A 0.07fF
C58769 INVX1_LOC_96/Y INVX1_LOC_46/A 0.02fF
C58770 NOR2X1_LOC_589/A NOR2X1_LOC_78/A 0.04fF
C58771 INVX1_LOC_134/Y NOR2X1_LOC_857/A 0.13fF
C58772 INVX1_LOC_36/A NAND2X1_LOC_572/B 0.07fF
C58773 INVX1_LOC_103/A INVX1_LOC_109/A 0.00fF
C58774 NOR2X1_LOC_720/B NAND2X1_LOC_96/A 0.02fF
C58775 NOR2X1_LOC_250/Y INVX1_LOC_29/A 0.04fF
C58776 INVX1_LOC_2/Y NOR2X1_LOC_87/Y 0.16fF
C58777 INVX1_LOC_57/A NOR2X1_LOC_280/a_36_216# 0.00fF
C58778 INVX1_LOC_199/A INVX1_LOC_22/A 0.03fF
C58779 INVX1_LOC_57/Y INVX1_LOC_285/A 0.38fF
C58780 NAND2X1_LOC_785/Y NOR2X1_LOC_495/a_36_216# 0.00fF
C58781 INVX1_LOC_5/A INVX1_LOC_271/Y 0.07fF
C58782 NAND2X1_LOC_563/A INVX1_LOC_76/A 0.00fF
C58783 NAND2X1_LOC_198/B NOR2X1_LOC_831/B 0.18fF
C58784 INVX1_LOC_57/Y INVX1_LOC_265/Y 0.03fF
C58785 NOR2X1_LOC_335/a_36_216# INVX1_LOC_91/A 0.01fF
C58786 NAND2X1_LOC_799/A NOR2X1_LOC_89/A 1.75fF
C58787 INPUT_3 NAND2X1_LOC_82/Y 0.12fF
C58788 NOR2X1_LOC_526/Y VDD 0.23fF
C58789 NOR2X1_LOC_817/Y NOR2X1_LOC_847/B 0.10fF
C58790 NOR2X1_LOC_816/A NOR2X1_LOC_189/a_36_216# 0.00fF
C58791 NOR2X1_LOC_561/Y NOR2X1_LOC_275/A 0.02fF
C58792 INVX1_LOC_49/A NOR2X1_LOC_155/A 0.06fF
C58793 INVX1_LOC_36/A NAND2X1_LOC_219/B 0.00fF
C58794 NOR2X1_LOC_516/B NOR2X1_LOC_138/a_36_216# 0.00fF
C58795 NOR2X1_LOC_234/Y INVX1_LOC_118/A -0.01fF
C58796 NAND2X1_LOC_481/a_36_24# INVX1_LOC_63/A 0.00fF
C58797 NOR2X1_LOC_180/B INVX1_LOC_91/A 0.07fF
C58798 NAND2X1_LOC_555/Y NAND2X1_LOC_20/a_36_24# 0.01fF
C58799 NOR2X1_LOC_654/A NOR2X1_LOC_109/Y 0.30fF
C58800 NAND2X1_LOC_223/A NAND2X1_LOC_473/A 0.07fF
C58801 INVX1_LOC_234/A NOR2X1_LOC_24/Y 0.07fF
C58802 INVX1_LOC_34/A INVX1_LOC_92/A 0.41fF
C58803 NOR2X1_LOC_286/Y INVX1_LOC_15/A 0.03fF
C58804 INVX1_LOC_58/A NOR2X1_LOC_53/Y 0.05fF
C58805 NOR2X1_LOC_379/a_36_216# NAND2X1_LOC_425/Y 0.01fF
C58806 NAND2X1_LOC_357/B NOR2X1_LOC_743/Y 0.01fF
C58807 INVX1_LOC_1/A INVX1_LOC_87/A 0.06fF
C58808 NOR2X1_LOC_52/B NOR2X1_LOC_88/A 0.08fF
C58809 NAND2X1_LOC_175/Y NAND2X1_LOC_780/Y 0.05fF
C58810 NOR2X1_LOC_588/A INVX1_LOC_140/A 0.10fF
C58811 INVX1_LOC_121/A INVX1_LOC_14/Y 0.02fF
C58812 INVX1_LOC_69/Y NOR2X1_LOC_548/A 0.01fF
C58813 INVX1_LOC_73/A INVX1_LOC_91/A 0.07fF
C58814 INVX1_LOC_14/A NOR2X1_LOC_415/Y 0.06fF
C58815 INVX1_LOC_1/A INVX1_LOC_175/A 0.26fF
C58816 INVX1_LOC_24/A NOR2X1_LOC_36/B 0.15fF
C58817 NOR2X1_LOC_216/Y NOR2X1_LOC_269/Y 0.00fF
C58818 INVX1_LOC_266/Y INVX1_LOC_307/A 0.10fF
C58819 INVX1_LOC_208/A INVX1_LOC_9/A 0.19fF
C58820 NOR2X1_LOC_214/B INVX1_LOC_76/A 0.08fF
C58821 INVX1_LOC_18/A NOR2X1_LOC_89/A 0.25fF
C58822 NOR2X1_LOC_576/B INVX1_LOC_46/A 3.04fF
C58823 NAND2X1_LOC_728/Y NOR2X1_LOC_89/A 0.12fF
C58824 INVX1_LOC_56/A INVX1_LOC_118/A 0.03fF
C58825 NOR2X1_LOC_516/B INVX1_LOC_9/A 0.03fF
C58826 NOR2X1_LOC_433/A INVX1_LOC_186/Y 0.08fF
C58827 NAND2X1_LOC_214/B NOR2X1_LOC_392/Y 0.08fF
C58828 INVX1_LOC_2/A NOR2X1_LOC_155/A 0.17fF
C58829 INVX1_LOC_187/Y INVX1_LOC_140/A 0.47fF
C58830 NOR2X1_LOC_318/B NOR2X1_LOC_188/A 0.05fF
C58831 NOR2X1_LOC_593/Y INVX1_LOC_186/Y 0.02fF
C58832 INVX1_LOC_75/A NOR2X1_LOC_657/B 0.19fF
C58833 INVX1_LOC_40/A NOR2X1_LOC_78/Y 0.03fF
C58834 NAND2X1_LOC_323/B NOR2X1_LOC_809/B 0.35fF
C58835 INVX1_LOC_224/A NOR2X1_LOC_843/B 0.03fF
C58836 NAND2X1_LOC_778/Y INVX1_LOC_233/A 0.10fF
C58837 NAND2X1_LOC_563/Y INVX1_LOC_84/A 0.44fF
C58838 NOR2X1_LOC_798/A NOR2X1_LOC_434/A 0.01fF
C58839 INVX1_LOC_298/Y INVX1_LOC_245/Y 0.04fF
C58840 NAND2X1_LOC_802/A INVX1_LOC_12/A 0.01fF
C58841 INVX1_LOC_188/A INVX1_LOC_78/A 0.03fF
C58842 NOR2X1_LOC_576/B NOR2X1_LOC_766/Y 0.05fF
C58843 NOR2X1_LOC_238/Y INVX1_LOC_42/A 0.08fF
C58844 INVX1_LOC_11/A NOR2X1_LOC_843/B 8.00fF
C58845 NOR2X1_LOC_363/a_36_216# INVX1_LOC_290/Y 0.01fF
C58846 INVX1_LOC_172/A NOR2X1_LOC_89/A 7.22fF
C58847 INVX1_LOC_140/A NOR2X1_LOC_305/Y 0.10fF
C58848 INVX1_LOC_17/A INVX1_LOC_50/A 0.06fF
C58849 NOR2X1_LOC_87/B INVX1_LOC_63/A 0.12fF
C58850 NOR2X1_LOC_647/A NOR2X1_LOC_647/B 0.02fF
C58851 INVX1_LOC_256/A NOR2X1_LOC_658/a_36_216# 0.02fF
C58852 NOR2X1_LOC_657/a_36_216# INVX1_LOC_64/A 0.01fF
C58853 INVX1_LOC_39/A NAND2X1_LOC_35/Y 0.02fF
C58854 NOR2X1_LOC_387/A INPUT_4 0.04fF
C58855 NAND2X1_LOC_840/Y INVX1_LOC_20/A 0.02fF
C58856 NOR2X1_LOC_218/Y NOR2X1_LOC_155/A 0.02fF
C58857 NOR2X1_LOC_826/Y NOR2X1_LOC_92/Y 0.03fF
C58858 NOR2X1_LOC_597/Y NAND2X1_LOC_453/A 0.02fF
C58859 INVX1_LOC_49/A NOR2X1_LOC_833/B 0.04fF
C58860 NOR2X1_LOC_52/B INVX1_LOC_186/Y 0.02fF
C58861 INVX1_LOC_141/Y NAND2X1_LOC_175/Y 0.09fF
C58862 INVX1_LOC_17/A NOR2X1_LOC_105/Y 0.00fF
C58863 INVX1_LOC_53/Y NOR2X1_LOC_831/B 0.07fF
C58864 INVX1_LOC_285/Y NOR2X1_LOC_137/B 0.06fF
C58865 INVX1_LOC_233/A NOR2X1_LOC_15/Y 0.09fF
C58866 NAND2X1_LOC_811/Y INVX1_LOC_12/A 3.27fF
C58867 INVX1_LOC_312/Y NAND2X1_LOC_175/Y 0.17fF
C58868 NOR2X1_LOC_272/Y INVX1_LOC_13/Y 0.10fF
C58869 NOR2X1_LOC_471/Y INVX1_LOC_50/A 0.02fF
C58870 NAND2X1_LOC_23/a_36_24# NAND2X1_LOC_555/Y 0.00fF
C58871 INVX1_LOC_45/A NOR2X1_LOC_278/Y 0.03fF
C58872 INVX1_LOC_25/A NOR2X1_LOC_82/A 0.49fF
C58873 INVX1_LOC_59/A INVX1_LOC_5/A 0.00fF
C58874 NOR2X1_LOC_411/A INVX1_LOC_269/A 0.01fF
C58875 INVX1_LOC_45/Y NAND2X1_LOC_647/B 0.04fF
C58876 NAND2X1_LOC_672/B NOR2X1_LOC_673/A 0.14fF
C58877 NAND2X1_LOC_660/Y NOR2X1_LOC_58/Y 0.06fF
C58878 NOR2X1_LOC_590/A NOR2X1_LOC_383/B 0.10fF
C58879 NOR2X1_LOC_361/Y INVX1_LOC_272/A 0.12fF
C58880 NOR2X1_LOC_178/Y INVX1_LOC_269/A 0.10fF
C58881 INVX1_LOC_235/A INVX1_LOC_27/A 0.01fF
C58882 NOR2X1_LOC_817/Y NOR2X1_LOC_660/Y 0.77fF
C58883 INVX1_LOC_266/Y INVX1_LOC_12/A 0.08fF
C58884 NOR2X1_LOC_78/B INVX1_LOC_49/Y 0.04fF
C58885 NOR2X1_LOC_357/Y INVX1_LOC_78/Y 0.00fF
C58886 NAND2X1_LOC_729/B INVX1_LOC_11/Y 0.05fF
C58887 INVX1_LOC_21/A INVX1_LOC_239/A 1.23fF
C58888 NOR2X1_LOC_449/a_36_216# NAND2X1_LOC_470/B 0.00fF
C58889 NOR2X1_LOC_238/Y INVX1_LOC_78/A 0.40fF
C58890 INVX1_LOC_98/A INVX1_LOC_20/A 0.01fF
C58891 INVX1_LOC_16/A NOR2X1_LOC_631/A 0.14fF
C58892 NOR2X1_LOC_152/Y NOR2X1_LOC_681/a_36_216# 0.01fF
C58893 NOR2X1_LOC_15/Y NOR2X1_LOC_798/A 0.03fF
C58894 INVX1_LOC_72/A NOR2X1_LOC_72/Y 0.03fF
C58895 INVX1_LOC_36/A NOR2X1_LOC_654/A 0.02fF
C58896 NOR2X1_LOC_78/A INVX1_LOC_20/A 0.07fF
C58897 INVX1_LOC_89/A NOR2X1_LOC_216/B 0.04fF
C58898 INVX1_LOC_223/A INVX1_LOC_57/A 0.05fF
C58899 INVX1_LOC_226/Y INVX1_LOC_19/A 0.08fF
C58900 INVX1_LOC_24/A INVX1_LOC_26/A 0.19fF
C58901 NOR2X1_LOC_78/B INVX1_LOC_99/A 0.04fF
C58902 INVX1_LOC_71/A NOR2X1_LOC_278/Y 0.16fF
C58903 NOR2X1_LOC_272/Y INVX1_LOC_88/A 0.03fF
C58904 NOR2X1_LOC_716/B NOR2X1_LOC_80/Y 0.42fF
C58905 NOR2X1_LOC_32/B NAND2X1_LOC_577/A 0.01fF
C58906 NAND2X1_LOC_563/Y INVX1_LOC_15/A 0.07fF
C58907 NAND2X1_LOC_783/Y NOR2X1_LOC_109/Y 0.05fF
C58908 NAND2X1_LOC_850/Y NOR2X1_LOC_46/a_36_216# 0.00fF
C58909 INVX1_LOC_58/A NOR2X1_LOC_52/Y 0.09fF
C58910 NOR2X1_LOC_92/Y NAND2X1_LOC_303/Y 0.10fF
C58911 VDD NOR2X1_LOC_595/Y 0.44fF
C58912 NAND2X1_LOC_706/Y NAND2X1_LOC_725/B 0.01fF
C58913 NOR2X1_LOC_344/A NAND2X1_LOC_72/B 0.02fF
C58914 INVX1_LOC_144/A INVX1_LOC_118/A 0.08fF
C58915 INVX1_LOC_6/A NAND2X1_LOC_423/a_36_24# 0.01fF
C58916 INVX1_LOC_269/A INVX1_LOC_163/A 0.01fF
C58917 NOR2X1_LOC_390/a_36_216# NOR2X1_LOC_334/Y 0.01fF
C58918 INVX1_LOC_215/A NAND2X1_LOC_74/B 0.07fF
C58919 INVX1_LOC_10/A INVX1_LOC_19/A 0.10fF
C58920 INVX1_LOC_79/Y INVX1_LOC_53/A 0.02fF
C58921 NOR2X1_LOC_709/B INVX1_LOC_6/A 0.00fF
C58922 NOR2X1_LOC_168/B NOR2X1_LOC_623/B 0.03fF
C58923 NOR2X1_LOC_253/a_36_216# NOR2X1_LOC_238/Y 0.00fF
C58924 NOR2X1_LOC_780/B NOR2X1_LOC_783/A 0.20fF
C58925 NOR2X1_LOC_557/Y INVX1_LOC_26/A 0.27fF
C58926 NOR2X1_LOC_252/a_36_216# INVX1_LOC_42/A 0.00fF
C58927 NAND2X1_LOC_573/A NAND2X1_LOC_81/B 0.03fF
C58928 VDD INVX1_LOC_115/Y 0.41fF
C58929 INVX1_LOC_22/A NAND2X1_LOC_254/Y 0.03fF
C58930 NAND2X1_LOC_350/A NAND2X1_LOC_714/B 0.12fF
C58931 NOR2X1_LOC_255/Y INVX1_LOC_24/A 0.00fF
C58932 NOR2X1_LOC_574/A INVX1_LOC_78/A 0.01fF
C58933 NAND2X1_LOC_303/Y NAND2X1_LOC_568/A 0.03fF
C58934 NOR2X1_LOC_516/B NOR2X1_LOC_861/Y 0.10fF
C58935 INVX1_LOC_83/A INVX1_LOC_49/Y 0.01fF
C58936 INPUT_0 INVX1_LOC_92/A 0.10fF
C58937 NOR2X1_LOC_82/A INVX1_LOC_1/A 0.14fF
C58938 NAND2X1_LOC_711/B NAND2X1_LOC_804/A 0.05fF
C58939 INVX1_LOC_315/Y INVX1_LOC_9/A 0.08fF
C58940 INVX1_LOC_134/A INVX1_LOC_1/A 0.03fF
C58941 INVX1_LOC_278/A INVX1_LOC_181/Y 0.00fF
C58942 INVX1_LOC_147/A NOR2X1_LOC_841/A 0.07fF
C58943 D_INPUT_0 INVX1_LOC_29/A 0.62fF
C58944 NOR2X1_LOC_299/Y INVX1_LOC_167/A 0.01fF
C58945 NOR2X1_LOC_772/B NAND2X1_LOC_364/A 0.35fF
C58946 NOR2X1_LOC_826/Y NAND2X1_LOC_837/Y 0.12fF
C58947 NOR2X1_LOC_619/a_36_216# INVX1_LOC_24/A 0.00fF
C58948 NAND2X1_LOC_280/a_36_24# INVX1_LOC_117/A 0.01fF
C58949 NOR2X1_LOC_113/B NOR2X1_LOC_831/B 0.14fF
C58950 INVX1_LOC_12/Y INVX1_LOC_76/A 0.06fF
C58951 NOR2X1_LOC_254/Y NOR2X1_LOC_748/A 0.65fF
C58952 INVX1_LOC_13/Y NAND2X1_LOC_364/A 0.03fF
C58953 NOR2X1_LOC_789/A INVX1_LOC_32/A 0.02fF
C58954 NOR2X1_LOC_598/B INVX1_LOC_49/A 0.50fF
C58955 NOR2X1_LOC_99/B NAND2X1_LOC_206/B 0.04fF
C58956 INVX1_LOC_46/A NOR2X1_LOC_492/a_36_216# 0.00fF
C58957 INVX1_LOC_76/A NOR2X1_LOC_492/Y 0.03fF
C58958 INVX1_LOC_103/A INVX1_LOC_246/A 0.02fF
C58959 NAND2X1_LOC_702/a_36_24# NAND2X1_LOC_198/B 0.00fF
C58960 NAND2X1_LOC_860/A INVX1_LOC_33/A 0.04fF
C58961 NOR2X1_LOC_309/Y NOR2X1_LOC_654/A 0.02fF
C58962 INVX1_LOC_162/Y INVX1_LOC_57/A 0.01fF
C58963 INVX1_LOC_51/A INVX1_LOC_49/A 0.00fF
C58964 INVX1_LOC_143/A INVX1_LOC_26/A 0.07fF
C58965 NOR2X1_LOC_848/Y INVX1_LOC_110/Y 0.04fF
C58966 INVX1_LOC_21/A NOR2X1_LOC_91/Y 0.03fF
C58967 NAND2X1_LOC_36/A INVX1_LOC_1/A 1.18fF
C58968 INVX1_LOC_34/A INVX1_LOC_53/A 0.11fF
C58969 NOR2X1_LOC_817/a_36_216# INVX1_LOC_31/A 0.01fF
C58970 INVX1_LOC_33/A NOR2X1_LOC_634/Y 0.02fF
C58971 INVX1_LOC_200/Y NOR2X1_LOC_315/Y 0.00fF
C58972 INVX1_LOC_35/A NOR2X1_LOC_551/B 0.03fF
C58973 NAND2X1_LOC_656/Y INVX1_LOC_32/A 0.23fF
C58974 NOR2X1_LOC_43/Y INVX1_LOC_117/Y 0.04fF
C58975 INVX1_LOC_268/A INVX1_LOC_78/A 0.02fF
C58976 NOR2X1_LOC_664/Y NOR2X1_LOC_392/Y 0.05fF
C58977 INVX1_LOC_64/A NAND2X1_LOC_139/A 0.02fF
C58978 NAND2X1_LOC_211/Y INVX1_LOC_9/A 0.37fF
C58979 INVX1_LOC_35/A INVX1_LOC_213/Y 0.08fF
C58980 INVX1_LOC_226/Y INVX1_LOC_26/Y 0.07fF
C58981 NOR2X1_LOC_343/a_36_216# NAND2X1_LOC_574/A 0.01fF
C58982 INVX1_LOC_166/A INVX1_LOC_197/A -0.02fF
C58983 NOR2X1_LOC_757/Y INVX1_LOC_270/A 0.10fF
C58984 INVX1_LOC_88/A NAND2X1_LOC_364/A 0.01fF
C58985 NOR2X1_LOC_33/A NOR2X1_LOC_33/Y 0.02fF
C58986 NOR2X1_LOC_67/A D_INPUT_1 0.20fF
C58987 INVX1_LOC_2/A NOR2X1_LOC_598/B 0.03fF
C58988 INVX1_LOC_5/A NOR2X1_LOC_144/Y 0.00fF
C58989 NOR2X1_LOC_2/Y INPUT_7 0.00fF
C58990 NOR2X1_LOC_83/Y NAND2X1_LOC_63/Y 0.04fF
C58991 NAND2X1_LOC_231/Y INVX1_LOC_53/A 0.03fF
C58992 NAND2X1_LOC_45/a_36_24# NOR2X1_LOC_242/A 0.00fF
C58993 NAND2X1_LOC_762/a_36_24# INVX1_LOC_11/A 0.00fF
C58994 INVX1_LOC_11/A INVX1_LOC_18/A 13.80fF
C58995 INVX1_LOC_92/Y INVX1_LOC_125/A 0.01fF
C58996 NAND2X1_LOC_560/A NOR2X1_LOC_754/A 0.00fF
C58997 INVX1_LOC_251/Y NAND2X1_LOC_363/B 0.16fF
C58998 NAND2X1_LOC_656/Y NAND2X1_LOC_175/Y 0.01fF
C58999 NOR2X1_LOC_636/A NAND2X1_LOC_149/Y 0.04fF
C59000 INVX1_LOC_64/A NOR2X1_LOC_644/Y 0.08fF
C59001 INVX1_LOC_45/A INVX1_LOC_236/Y 0.01fF
C59002 NOR2X1_LOC_252/Y INVX1_LOC_50/A 0.16fF
C59003 INVX1_LOC_286/A NAND2X1_LOC_74/B 0.07fF
C59004 INVX1_LOC_191/A INVX1_LOC_12/A 0.07fF
C59005 NAND2X1_LOC_116/A NOR2X1_LOC_849/A 0.03fF
C59006 VDD NOR2X1_LOC_156/Y 0.12fF
C59007 INVX1_LOC_232/A INVX1_LOC_129/A 0.08fF
C59008 NAND2X1_LOC_9/Y INVX1_LOC_226/A 0.03fF
C59009 NOR2X1_LOC_705/B NOR2X1_LOC_68/A 0.04fF
C59010 INVX1_LOC_196/Y NOR2X1_LOC_334/Y 0.07fF
C59011 NAND2X1_LOC_794/B INVX1_LOC_240/A 0.15fF
C59012 INVX1_LOC_33/Y INVX1_LOC_185/A 0.00fF
C59013 INVX1_LOC_233/Y INVX1_LOC_280/Y 0.07fF
C59014 INVX1_LOC_47/A INVX1_LOC_78/A 0.06fF
C59015 INVX1_LOC_2/A NAND2X1_LOC_715/B 0.64fF
C59016 NOR2X1_LOC_130/A INVX1_LOC_26/A 0.06fF
C59017 INVX1_LOC_100/A NAND2X1_LOC_254/Y -0.01fF
C59018 NOR2X1_LOC_498/Y NAND2X1_LOC_705/Y 0.09fF
C59019 NOR2X1_LOC_643/A NOR2X1_LOC_643/Y 0.06fF
C59020 INVX1_LOC_11/A NOR2X1_LOC_713/B 0.12fF
C59021 INVX1_LOC_227/A NOR2X1_LOC_383/B 0.08fF
C59022 NOR2X1_LOC_690/A NOR2X1_LOC_92/Y 0.01fF
C59023 INVX1_LOC_48/A NOR2X1_LOC_67/Y 0.13fF
C59024 NOR2X1_LOC_311/Y INVX1_LOC_49/Y 0.00fF
C59025 INVX1_LOC_269/A INVX1_LOC_237/Y 0.02fF
C59026 INVX1_LOC_35/A INVX1_LOC_208/Y 0.45fF
C59027 NOR2X1_LOC_413/Y NOR2X1_LOC_92/Y 0.02fF
C59028 D_INPUT_3 NAND2X1_LOC_574/A 0.59fF
C59029 INVX1_LOC_199/A INVX1_LOC_186/Y 0.05fF
C59030 NAND2X1_LOC_799/A NOR2X1_LOC_433/A 0.03fF
C59031 NAND2X1_LOC_338/B INVX1_LOC_50/Y 0.07fF
C59032 NOR2X1_LOC_538/B NAND2X1_LOC_361/Y 0.01fF
C59033 NOR2X1_LOC_690/Y NAND2X1_LOC_804/A 0.01fF
C59034 INVX1_LOC_2/Y NOR2X1_LOC_673/A 0.03fF
C59035 NOR2X1_LOC_205/Y INVX1_LOC_153/Y 0.18fF
C59036 NOR2X1_LOC_799/B INVX1_LOC_19/A 0.07fF
C59037 NAND2X1_LOC_543/a_36_24# INVX1_LOC_41/Y 0.00fF
C59038 NAND2X1_LOC_364/A NOR2X1_LOC_500/B 0.10fF
C59039 NOR2X1_LOC_658/Y NOR2X1_LOC_759/A 0.15fF
C59040 D_INPUT_3 NOR2X1_LOC_23/a_36_216# 0.00fF
C59041 INVX1_LOC_64/A NAND2X1_LOC_112/Y 0.02fF
C59042 INVX1_LOC_25/A INVX1_LOC_306/A 0.01fF
C59043 NAND2X1_LOC_432/a_36_24# NAND2X1_LOC_453/A 0.00fF
C59044 INVX1_LOC_95/A NAND2X1_LOC_74/B 2.23fF
C59045 INVX1_LOC_65/A NOR2X1_LOC_830/Y 0.03fF
C59046 NAND2X1_LOC_214/B INVX1_LOC_25/Y 0.01fF
C59047 NAND2X1_LOC_22/a_36_24# INVX1_LOC_174/A 0.01fF
C59048 INVX1_LOC_202/A NOR2X1_LOC_441/Y 0.40fF
C59049 NAND2X1_LOC_391/Y NAND2X1_LOC_181/Y 0.02fF
C59050 NAND2X1_LOC_35/Y NAND2X1_LOC_735/B 0.03fF
C59051 INVX1_LOC_102/Y NOR2X1_LOC_278/Y 0.07fF
C59052 NOR2X1_LOC_454/Y NAND2X1_LOC_661/B 0.02fF
C59053 INVX1_LOC_234/A NOR2X1_LOC_392/Y 0.01fF
C59054 NAND2X1_LOC_731/Y NAND2X1_LOC_856/A 0.03fF
C59055 NOR2X1_LOC_785/A INVX1_LOC_310/Y 0.04fF
C59056 INVX1_LOC_285/Y INVX1_LOC_4/Y 0.10fF
C59057 INVX1_LOC_27/A INVX1_LOC_25/Y 0.07fF
C59058 NAND2X1_LOC_654/B INVX1_LOC_296/A 0.03fF
C59059 NAND2X1_LOC_468/B INVX1_LOC_109/Y 0.00fF
C59060 NOR2X1_LOC_205/Y INVX1_LOC_177/A 0.03fF
C59061 NOR2X1_LOC_188/A INVX1_LOC_87/A 0.04fF
C59062 NOR2X1_LOC_389/A INVX1_LOC_63/Y 0.10fF
C59063 INVX1_LOC_40/A NAND2X1_LOC_473/A 0.16fF
C59064 NOR2X1_LOC_703/A NOR2X1_LOC_383/B 0.01fF
C59065 INVX1_LOC_49/Y INVX1_LOC_46/A 0.03fF
C59066 NOR2X1_LOC_824/A INVX1_LOC_25/Y 0.03fF
C59067 INVX1_LOC_95/Y INVX1_LOC_42/A 0.12fF
C59068 NOR2X1_LOC_186/Y NOR2X1_LOC_589/A 0.07fF
C59069 INVX1_LOC_5/A INVX1_LOC_279/A 0.09fF
C59070 NAND2X1_LOC_624/B NAND2X1_LOC_523/a_36_24# 0.01fF
C59071 NOR2X1_LOC_548/B INVX1_LOC_87/A 0.43fF
C59072 INVX1_LOC_27/A NOR2X1_LOC_302/B 0.05fF
C59073 NOR2X1_LOC_454/Y NOR2X1_LOC_229/Y 0.05fF
C59074 INVX1_LOC_11/A INVX1_LOC_34/Y 0.07fF
C59075 NAND2X1_LOC_733/Y NAND2X1_LOC_811/Y 0.05fF
C59076 INVX1_LOC_1/A NOR2X1_LOC_731/Y 0.01fF
C59077 NOR2X1_LOC_78/A INVX1_LOC_4/A 0.09fF
C59078 INVX1_LOC_36/A NOR2X1_LOC_716/B 0.15fF
C59079 NAND2X1_LOC_571/Y NAND2X1_LOC_735/B 0.03fF
C59080 INVX1_LOC_55/Y NOR2X1_LOC_717/A 0.03fF
C59081 INVX1_LOC_303/A NAND2X1_LOC_364/A 0.47fF
C59082 NAND2X1_LOC_67/Y INVX1_LOC_208/A 0.25fF
C59083 NAND2X1_LOC_59/a_36_24# INVX1_LOC_1/A 0.00fF
C59084 INVX1_LOC_21/A NOR2X1_LOC_543/A 0.01fF
C59085 INVX1_LOC_180/Y NOR2X1_LOC_592/B 0.01fF
C59086 NOR2X1_LOC_433/A INVX1_LOC_18/A 0.10fF
C59087 INVX1_LOC_115/A NAND2X1_LOC_220/B 0.04fF
C59088 INVX1_LOC_124/Y INVX1_LOC_8/A 0.00fF
C59089 NOR2X1_LOC_289/a_36_216# INVX1_LOC_88/A 0.00fF
C59090 NAND2X1_LOC_725/A NAND2X1_LOC_648/A 0.48fF
C59091 INVX1_LOC_99/Y INVX1_LOC_89/A 0.03fF
C59092 INVX1_LOC_75/A INVX1_LOC_271/A 0.10fF
C59093 NOR2X1_LOC_456/Y INVX1_LOC_182/A 0.10fF
C59094 NOR2X1_LOC_859/Y INVX1_LOC_29/A 0.00fF
C59095 NAND2X1_LOC_733/Y NOR2X1_LOC_821/Y 0.02fF
C59096 NAND2X1_LOC_288/a_36_24# INVX1_LOC_46/A 0.00fF
C59097 NOR2X1_LOC_593/Y INVX1_LOC_18/A 0.01fF
C59098 NOR2X1_LOC_68/A NOR2X1_LOC_172/Y 0.12fF
C59099 NOR2X1_LOC_19/B NOR2X1_LOC_392/Y 0.52fF
C59100 NOR2X1_LOC_588/A INVX1_LOC_78/A 0.08fF
C59101 NAND2X1_LOC_181/a_36_24# INVX1_LOC_1/A 0.06fF
C59102 NAND2X1_LOC_339/a_36_24# INVX1_LOC_30/A 0.01fF
C59103 NOR2X1_LOC_186/Y INVX1_LOC_171/A 0.01fF
C59104 INVX1_LOC_2/A NOR2X1_LOC_372/A 0.08fF
C59105 NOR2X1_LOC_791/A INVX1_LOC_8/A -0.00fF
C59106 NOR2X1_LOC_590/A NOR2X1_LOC_168/A 0.07fF
C59107 NOR2X1_LOC_533/Y INVX1_LOC_16/A 0.03fF
C59108 NAND2X1_LOC_848/A INVX1_LOC_29/A 0.03fF
C59109 NAND2X1_LOC_725/B NOR2X1_LOC_32/Y 0.01fF
C59110 NOR2X1_LOC_68/A NOR2X1_LOC_147/B 3.13fF
C59111 NOR2X1_LOC_763/Y NOR2X1_LOC_763/A 0.06fF
C59112 INVX1_LOC_103/A INVX1_LOC_290/A 0.10fF
C59113 INVX1_LOC_313/Y INVX1_LOC_50/Y 0.07fF
C59114 NOR2X1_LOC_859/A NAND2X1_LOC_116/A 0.00fF
C59115 INVX1_LOC_224/Y NOR2X1_LOC_391/Y -0.04fF
C59116 NOR2X1_LOC_564/a_36_216# NOR2X1_LOC_383/B 0.00fF
C59117 VDD D_INPUT_5 1.42fF
C59118 INPUT_0 INVX1_LOC_53/A 0.13fF
C59119 INVX1_LOC_227/Y INVX1_LOC_104/A 0.03fF
C59120 NOR2X1_LOC_78/B NAND2X1_LOC_208/B 0.83fF
C59121 NOR2X1_LOC_673/B INVX1_LOC_46/Y 0.02fF
C59122 NOR2X1_LOC_596/A INVX1_LOC_63/Y 0.01fF
C59123 NOR2X1_LOC_52/B INVX1_LOC_18/A 0.30fF
C59124 NOR2X1_LOC_553/a_36_216# NOR2X1_LOC_500/Y 0.01fF
C59125 NAND2X1_LOC_303/Y NOR2X1_LOC_299/Y 0.15fF
C59126 INVX1_LOC_187/Y INVX1_LOC_78/A 0.21fF
C59127 INVX1_LOC_304/Y NOR2X1_LOC_91/a_36_216# 0.00fF
C59128 NOR2X1_LOC_234/Y INVX1_LOC_61/A 0.01fF
C59129 NOR2X1_LOC_690/A NAND2X1_LOC_837/Y 0.07fF
C59130 NAND2X1_LOC_207/B INVX1_LOC_9/A 0.00fF
C59131 NOR2X1_LOC_142/Y NOR2X1_LOC_759/Y 0.05fF
C59132 NOR2X1_LOC_209/B INVX1_LOC_301/A 0.21fF
C59133 INVX1_LOC_36/A INVX1_LOC_98/Y 0.05fF
C59134 INVX1_LOC_77/A INVX1_LOC_155/A 0.10fF
C59135 NAND2X1_LOC_352/B INVX1_LOC_53/Y 0.01fF
C59136 INVX1_LOC_254/A INVX1_LOC_41/A 0.00fF
C59137 INVX1_LOC_54/A NAND2X1_LOC_74/B 0.03fF
C59138 NAND2X1_LOC_357/B NAND2X1_LOC_198/B 0.10fF
C59139 NOR2X1_LOC_160/B NOR2X1_LOC_719/A 0.07fF
C59140 NOR2X1_LOC_531/a_36_216# INVX1_LOC_177/A 0.00fF
C59141 NAND2X1_LOC_214/B INVX1_LOC_75/A 0.07fF
C59142 NAND2X1_LOC_34/a_36_24# INVX1_LOC_72/A 0.01fF
C59143 INVX1_LOC_19/A INVX1_LOC_307/A 0.07fF
C59144 NOR2X1_LOC_267/A INVX1_LOC_98/Y 0.04fF
C59145 NOR2X1_LOC_78/B NOR2X1_LOC_722/Y 0.01fF
C59146 NOR2X1_LOC_589/A NOR2X1_LOC_45/Y 0.17fF
C59147 NOR2X1_LOC_799/B INVX1_LOC_26/Y 0.03fF
C59148 INVX1_LOC_161/Y INVX1_LOC_10/A 0.07fF
C59149 NOR2X1_LOC_637/Y NOR2X1_LOC_52/B 0.17fF
C59150 NAND2X1_LOC_572/B INVX1_LOC_63/A 0.06fF
C59151 INVX1_LOC_12/A NOR2X1_LOC_508/a_36_216# 0.00fF
C59152 NOR2X1_LOC_65/B INVX1_LOC_95/Y 0.10fF
C59153 NOR2X1_LOC_160/B NOR2X1_LOC_561/Y 0.12fF
C59154 NOR2X1_LOC_574/A NOR2X1_LOC_152/Y 0.05fF
C59155 INVX1_LOC_19/A NOR2X1_LOC_445/B 3.64fF
C59156 INVX1_LOC_47/Y NOR2X1_LOC_536/A 0.19fF
C59157 NOR2X1_LOC_189/A INVX1_LOC_240/A 0.41fF
C59158 NOR2X1_LOC_15/Y NAND2X1_LOC_842/B 0.99fF
C59159 INVX1_LOC_46/Y INVX1_LOC_29/A 0.04fF
C59160 INVX1_LOC_27/A INVX1_LOC_75/A 1.77fF
C59161 INVX1_LOC_255/Y INVX1_LOC_40/Y 0.01fF
C59162 NOR2X1_LOC_498/Y NOR2X1_LOC_690/A 0.10fF
C59163 NOR2X1_LOC_716/B NOR2X1_LOC_309/Y 0.01fF
C59164 NAND2X1_LOC_787/A NOR2X1_LOC_45/B 0.04fF
C59165 INVX1_LOC_231/Y INVX1_LOC_240/A 0.03fF
C59166 NAND2X1_LOC_783/A INVX1_LOC_141/A 0.02fF
C59167 NOR2X1_LOC_769/A INVX1_LOC_268/A 0.01fF
C59168 NOR2X1_LOC_274/a_36_216# NOR2X1_LOC_655/B 0.12fF
C59169 NOR2X1_LOC_360/Y NOR2X1_LOC_568/a_36_216# 0.01fF
C59170 NAND2X1_LOC_338/B NOR2X1_LOC_559/B 0.05fF
C59171 INVX1_LOC_110/Y INVX1_LOC_135/A 0.01fF
C59172 INVX1_LOC_124/A INVX1_LOC_155/A 0.08fF
C59173 INVX1_LOC_64/A NOR2X1_LOC_78/A 2.87fF
C59174 INVX1_LOC_30/Y INVX1_LOC_72/A 0.15fF
C59175 INVX1_LOC_25/A INVX1_LOC_112/A 0.02fF
C59176 INVX1_LOC_25/A INVX1_LOC_59/Y 1.16fF
C59177 NAND2X1_LOC_219/B INVX1_LOC_63/A 0.11fF
C59178 NOR2X1_LOC_599/A INVX1_LOC_10/A 0.06fF
C59179 INVX1_LOC_310/A NAND2X1_LOC_361/Y 0.04fF
C59180 INVX1_LOC_58/A NOR2X1_LOC_603/Y 0.02fF
C59181 NAND2X1_LOC_466/Y NAND2X1_LOC_477/A 0.00fF
C59182 NAND2X1_LOC_454/Y INVX1_LOC_38/A 0.08fF
C59183 NOR2X1_LOC_483/B INVX1_LOC_85/Y 0.01fF
C59184 INVX1_LOC_93/Y NOR2X1_LOC_129/a_36_216# 0.00fF
C59185 NAND2X1_LOC_35/B INVX1_LOC_207/A 0.24fF
C59186 NOR2X1_LOC_443/Y INVX1_LOC_37/A 0.17fF
C59187 INVX1_LOC_286/A NAND2X1_LOC_793/a_36_24# 0.06fF
C59188 INVX1_LOC_47/Y NAND2X1_LOC_93/B 0.07fF
C59189 INVX1_LOC_271/A NAND2X1_LOC_453/A 0.67fF
C59190 INVX1_LOC_36/A NOR2X1_LOC_717/B 0.05fF
C59191 NAND2X1_LOC_392/A INVX1_LOC_71/A 0.01fF
C59192 INVX1_LOC_45/A NOR2X1_LOC_312/Y 0.00fF
C59193 NOR2X1_LOC_392/B NAND2X1_LOC_134/a_36_24# 0.06fF
C59194 NOR2X1_LOC_478/a_36_216# NOR2X1_LOC_68/A 0.00fF
C59195 INVX1_LOC_314/Y INVX1_LOC_22/A 0.04fF
C59196 NAND2X1_LOC_77/a_36_24# INVX1_LOC_123/A 0.01fF
C59197 NAND2X1_LOC_149/Y NOR2X1_LOC_377/a_36_216# 0.01fF
C59198 NOR2X1_LOC_476/Y INVX1_LOC_135/A 0.03fF
C59199 NOR2X1_LOC_194/Y NOR2X1_LOC_207/A 0.00fF
C59200 INVX1_LOC_34/A NOR2X1_LOC_78/B 0.19fF
C59201 INVX1_LOC_268/A NOR2X1_LOC_152/Y 0.02fF
C59202 NOR2X1_LOC_210/A INVX1_LOC_71/A 0.05fF
C59203 NOR2X1_LOC_211/Y NAND2X1_LOC_447/Y 0.06fF
C59204 INVX1_LOC_13/Y NOR2X1_LOC_405/A 0.03fF
C59205 INVX1_LOC_111/Y INVX1_LOC_104/A 0.01fF
C59206 NOR2X1_LOC_6/B NOR2X1_LOC_537/Y 0.06fF
C59207 NOR2X1_LOC_52/B INVX1_LOC_34/Y 0.00fF
C59208 NAND2X1_LOC_784/A NAND2X1_LOC_721/A 0.69fF
C59209 NAND2X1_LOC_338/B NOR2X1_LOC_6/B 0.13fF
C59210 NOR2X1_LOC_205/Y INVX1_LOC_285/Y 0.08fF
C59211 INVX1_LOC_12/A INVX1_LOC_19/A 0.10fF
C59212 NOR2X1_LOC_68/A INVX1_LOC_97/A 0.06fF
C59213 NOR2X1_LOC_778/B NOR2X1_LOC_348/B 0.02fF
C59214 INVX1_LOC_11/A NOR2X1_LOC_548/A 0.02fF
C59215 NOR2X1_LOC_498/Y NAND2X1_LOC_717/a_36_24# 0.00fF
C59216 NOR2X1_LOC_45/a_36_216# INVX1_LOC_54/A 0.00fF
C59217 INVX1_LOC_106/A INVX1_LOC_125/A 0.00fF
C59218 INVX1_LOC_12/A NOR2X1_LOC_11/Y 0.01fF
C59219 NAND2X1_LOC_470/B NAND2X1_LOC_798/B 0.01fF
C59220 NOR2X1_LOC_68/A INVX1_LOC_90/A 0.31fF
C59221 NAND2X1_LOC_714/B INVX1_LOC_291/Y 0.03fF
C59222 NOR2X1_LOC_816/A NAND2X1_LOC_858/B 0.02fF
C59223 NOR2X1_LOC_186/Y INVX1_LOC_20/A 0.11fF
C59224 NOR2X1_LOC_78/B NAND2X1_LOC_231/Y 0.10fF
C59225 NOR2X1_LOC_388/Y NOR2X1_LOC_577/a_36_216# 0.00fF
C59226 NOR2X1_LOC_576/B NAND2X1_LOC_866/A 1.01fF
C59227 NOR2X1_LOC_160/B INVX1_LOC_303/Y 0.06fF
C59228 NAND2X1_LOC_20/B INVX1_LOC_315/Y 0.01fF
C59229 NOR2X1_LOC_178/Y INVX1_LOC_12/Y 0.14fF
C59230 INVX1_LOC_225/A NOR2X1_LOC_589/A 0.07fF
C59231 INVX1_LOC_36/A NOR2X1_LOC_151/Y 0.01fF
C59232 INVX1_LOC_280/Y NOR2X1_LOC_526/Y 0.01fF
C59233 NAND2X1_LOC_708/Y NOR2X1_LOC_694/Y 0.00fF
C59234 INVX1_LOC_88/A NOR2X1_LOC_405/A 0.10fF
C59235 INVX1_LOC_45/A NOR2X1_LOC_97/A 0.19fF
C59236 INVX1_LOC_23/A NOR2X1_LOC_629/Y 0.01fF
C59237 NAND2X1_LOC_573/Y INVX1_LOC_20/A 0.17fF
C59238 NOR2X1_LOC_612/Y INVX1_LOC_29/Y 0.05fF
C59239 D_INPUT_0 NOR2X1_LOC_516/a_36_216# 0.00fF
C59240 INVX1_LOC_1/A INVX1_LOC_59/Y 0.03fF
C59241 INVX1_LOC_89/A NAND2X1_LOC_5/a_36_24# 0.00fF
C59242 INVX1_LOC_43/Y INVX1_LOC_98/A 0.00fF
C59243 NOR2X1_LOC_68/A NAND2X1_LOC_348/A 0.55fF
C59244 D_INPUT_0 INVX1_LOC_8/A 0.06fF
C59245 NOR2X1_LOC_778/B INVX1_LOC_22/A 0.04fF
C59246 INVX1_LOC_30/Y NOR2X1_LOC_537/Y 0.03fF
C59247 INVX1_LOC_89/A NOR2X1_LOC_254/Y 0.03fF
C59248 INVX1_LOC_33/A INVX1_LOC_85/Y 0.03fF
C59249 INVX1_LOC_225/A INVX1_LOC_171/A 0.01fF
C59250 NAND2X1_LOC_725/A INVX1_LOC_118/A 0.03fF
C59251 NOR2X1_LOC_457/A INVX1_LOC_247/A 0.05fF
C59252 NOR2X1_LOC_137/A INVX1_LOC_104/A 0.02fF
C59253 NAND2X1_LOC_173/a_36_24# NOR2X1_LOC_211/A 0.00fF
C59254 NAND2X1_LOC_288/B INVX1_LOC_285/A 0.01fF
C59255 NAND2X1_LOC_123/Y NOR2X1_LOC_577/Y 0.07fF
C59256 INVX1_LOC_182/A NOR2X1_LOC_550/B 0.10fF
C59257 NOR2X1_LOC_218/a_36_216# INVX1_LOC_71/A 0.02fF
C59258 INVX1_LOC_136/A INVX1_LOC_286/A 1.27fF
C59259 INVX1_LOC_24/A NOR2X1_LOC_368/A 0.12fF
C59260 NOR2X1_LOC_204/a_36_216# NAND2X1_LOC_348/A 0.00fF
C59261 INVX1_LOC_16/A INVX1_LOC_56/Y 0.09fF
C59262 INVX1_LOC_54/Y INVX1_LOC_150/A 0.00fF
C59263 NAND2X1_LOC_350/B NOR2X1_LOC_561/Y 0.01fF
C59264 INVX1_LOC_227/Y INVX1_LOC_206/Y 0.00fF
C59265 INVX1_LOC_30/A NOR2X1_LOC_45/B 3.51fF
C59266 NOR2X1_LOC_52/B NAND2X1_LOC_105/a_36_24# 0.00fF
C59267 INVX1_LOC_186/A INVX1_LOC_142/A 0.02fF
C59268 NAND2X1_LOC_363/B NOR2X1_LOC_862/B 0.10fF
C59269 NOR2X1_LOC_45/Y INVX1_LOC_147/Y 0.71fF
C59270 NOR2X1_LOC_392/Y NOR2X1_LOC_216/B 0.07fF
C59271 NOR2X1_LOC_607/A INVX1_LOC_69/Y 0.01fF
C59272 INVX1_LOC_54/Y INVX1_LOC_89/A 0.03fF
C59273 INVX1_LOC_208/A NOR2X1_LOC_561/Y 0.10fF
C59274 NAND2X1_LOC_850/Y NAND2X1_LOC_474/a_36_24# 0.00fF
C59275 NOR2X1_LOC_36/A INPUT_7 0.65fF
C59276 INVX1_LOC_147/A NOR2X1_LOC_172/Y 0.01fF
C59277 NOR2X1_LOC_160/B INVX1_LOC_76/A 0.17fF
C59278 NAND2X1_LOC_537/Y NOR2X1_LOC_816/Y 0.00fF
C59279 NOR2X1_LOC_576/B NOR2X1_LOC_505/Y 0.14fF
C59280 NOR2X1_LOC_516/B INVX1_LOC_7/A 0.25fF
C59281 INVX1_LOC_271/Y INVX1_LOC_42/A 0.01fF
C59282 INVX1_LOC_70/A INVX1_LOC_306/Y 0.03fF
C59283 NOR2X1_LOC_103/Y INVX1_LOC_129/Y 0.00fF
C59284 INVX1_LOC_136/A INVX1_LOC_95/A 0.06fF
C59285 NAND2X1_LOC_9/Y NAND2X1_LOC_456/Y 0.01fF
C59286 INVX1_LOC_18/A INVX1_LOC_199/A 0.07fF
C59287 NAND2X1_LOC_11/Y INVX1_LOC_244/A 0.16fF
C59288 INVX1_LOC_128/Y INVX1_LOC_32/A 0.00fF
C59289 INVX1_LOC_58/Y INVX1_LOC_63/A 2.34fF
C59290 NAND2X1_LOC_529/a_36_24# NAND2X1_LOC_96/A 0.00fF
C59291 NOR2X1_LOC_658/Y NOR2X1_LOC_357/Y 1.43fF
C59292 NOR2X1_LOC_758/a_36_216# NOR2X1_LOC_405/A 0.01fF
C59293 INVX1_LOC_123/Y INVX1_LOC_306/Y 0.02fF
C59294 INVX1_LOC_206/A INVX1_LOC_75/A 0.74fF
C59295 INPUT_0 INVX1_LOC_80/Y 0.01fF
C59296 INVX1_LOC_241/Y INVX1_LOC_242/A 0.17fF
C59297 NAND2X1_LOC_74/B NAND2X1_LOC_215/A 0.11fF
C59298 NOR2X1_LOC_500/B NOR2X1_LOC_857/A 0.10fF
C59299 NOR2X1_LOC_667/Y INVX1_LOC_33/Y 0.00fF
C59300 INVX1_LOC_57/Y NAND2X1_LOC_650/B 0.28fF
C59301 NOR2X1_LOC_250/Y INVX1_LOC_118/Y 0.28fF
C59302 INVX1_LOC_36/A NAND2X1_LOC_633/Y 0.06fF
C59303 NOR2X1_LOC_598/B NAND2X1_LOC_63/Y 0.34fF
C59304 INVX1_LOC_303/A NOR2X1_LOC_405/A 0.07fF
C59305 NAND2X1_LOC_778/Y INVX1_LOC_119/Y 1.06fF
C59306 NOR2X1_LOC_19/B INVX1_LOC_25/Y 0.00fF
C59307 INVX1_LOC_286/A NOR2X1_LOC_278/A 0.02fF
C59308 NOR2X1_LOC_180/B NOR2X1_LOC_553/B 0.01fF
C59309 NOR2X1_LOC_667/A NAND2X1_LOC_811/a_36_24# 0.00fF
C59310 NOR2X1_LOC_576/B NOR2X1_LOC_700/Y 0.03fF
C59311 INVX1_LOC_110/Y INVX1_LOC_280/A 0.02fF
C59312 NOR2X1_LOC_382/Y NOR2X1_LOC_813/Y 0.02fF
C59313 NOR2X1_LOC_360/Y VDD 1.50fF
C59314 INVX1_LOC_78/A INVX1_LOC_271/Y 0.08fF
C59315 NAND2X1_LOC_213/A INVX1_LOC_107/Y 0.00fF
C59316 NOR2X1_LOC_78/B INPUT_0 0.10fF
C59317 NOR2X1_LOC_276/Y INVX1_LOC_54/A 0.03fF
C59318 NOR2X1_LOC_703/B INVX1_LOC_117/A 0.12fF
C59319 NOR2X1_LOC_372/A INVX1_LOC_118/A 0.60fF
C59320 NOR2X1_LOC_843/A INVX1_LOC_65/A 0.02fF
C59321 NOR2X1_LOC_773/Y NAND2X1_LOC_858/B 0.07fF
C59322 INVX1_LOC_94/A INVX1_LOC_14/Y 0.10fF
C59323 NOR2X1_LOC_382/Y INVX1_LOC_280/A 0.00fF
C59324 INVX1_LOC_71/A NAND2X1_LOC_287/B 0.10fF
C59325 INVX1_LOC_132/A INVX1_LOC_20/A 0.07fF
C59326 NOR2X1_LOC_152/Y NOR2X1_LOC_305/Y 0.03fF
C59327 INVX1_LOC_210/Y INVX1_LOC_9/A 0.00fF
C59328 NAND2X1_LOC_634/Y NAND2X1_LOC_848/A 1.35fF
C59329 NOR2X1_LOC_486/Y NOR2X1_LOC_486/B 0.19fF
C59330 INVX1_LOC_18/A NAND2X1_LOC_699/a_36_24# 0.00fF
C59331 NOR2X1_LOC_15/Y INVX1_LOC_119/Y 0.02fF
C59332 NAND2X1_LOC_514/a_36_24# INVX1_LOC_79/A 0.00fF
C59333 INVX1_LOC_63/Y NAND2X1_LOC_469/B 0.08fF
C59334 NOR2X1_LOC_770/A VDD -0.00fF
C59335 INVX1_LOC_36/A NOR2X1_LOC_709/B 0.01fF
C59336 INVX1_LOC_82/A INVX1_LOC_316/A 0.25fF
C59337 NOR2X1_LOC_598/B INVX1_LOC_257/A 0.01fF
C59338 INVX1_LOC_298/A NOR2X1_LOC_89/A 0.09fF
C59339 INVX1_LOC_136/A NOR2X1_LOC_602/B 0.01fF
C59340 NOR2X1_LOC_68/A INVX1_LOC_38/A 0.49fF
C59341 NOR2X1_LOC_272/Y INVX1_LOC_272/A 0.27fF
C59342 NOR2X1_LOC_590/A INVX1_LOC_179/A 0.03fF
C59343 INVX1_LOC_50/A INVX1_LOC_94/Y 0.00fF
C59344 INVX1_LOC_98/A NAND2X1_LOC_850/Y 0.32fF
C59345 INPUT_3 NOR2X1_LOC_820/a_36_216# 0.00fF
C59346 INVX1_LOC_216/Y NOR2X1_LOC_649/B 0.01fF
C59347 NOR2X1_LOC_553/B NOR2X1_LOC_569/A 0.04fF
C59348 INVX1_LOC_207/A VDD 0.18fF
C59349 NAND2X1_LOC_181/Y INVX1_LOC_91/A 0.03fF
C59350 INPUT_0 NAND2X1_LOC_392/Y 0.03fF
C59351 INVX1_LOC_136/A INVX1_LOC_54/A 0.24fF
C59352 NOR2X1_LOC_602/A NOR2X1_LOC_743/Y 0.18fF
C59353 INVX1_LOC_225/A INVX1_LOC_20/A 0.03fF
C59354 NOR2X1_LOC_748/Y NOR2X1_LOC_9/Y 0.37fF
C59355 INVX1_LOC_284/Y NOR2X1_LOC_491/Y 0.00fF
C59356 INVX1_LOC_211/Y NOR2X1_LOC_697/Y 0.03fF
C59357 INVX1_LOC_34/A INVX1_LOC_46/A 2.58fF
C59358 INVX1_LOC_191/Y INVX1_LOC_187/A 0.00fF
C59359 NAND2X1_LOC_807/a_36_24# NOR2X1_LOC_652/Y 0.00fF
C59360 INVX1_LOC_8/A NOR2X1_LOC_266/B 0.00fF
C59361 NAND2X1_LOC_338/B NOR2X1_LOC_124/A 0.02fF
C59362 INVX1_LOC_27/A GATE_222 0.02fF
C59363 INVX1_LOC_83/A INPUT_0 0.06fF
C59364 NOR2X1_LOC_792/B VDD 0.00fF
C59365 NOR2X1_LOC_391/A INVX1_LOC_6/A 0.10fF
C59366 NOR2X1_LOC_300/Y INVX1_LOC_139/A 0.00fF
C59367 NOR2X1_LOC_188/Y NOR2X1_LOC_501/B 0.04fF
C59368 INVX1_LOC_27/A INVX1_LOC_283/A 0.01fF
C59369 INVX1_LOC_230/Y NAND2X1_LOC_206/Y 0.05fF
C59370 NOR2X1_LOC_184/a_36_216# NOR2X1_LOC_76/A 0.01fF
C59371 NOR2X1_LOC_15/Y INVX1_LOC_284/A 0.03fF
C59372 INVX1_LOC_5/A NOR2X1_LOC_38/B 2.01fF
C59373 INVX1_LOC_90/A NOR2X1_LOC_2/Y 0.14fF
C59374 NOR2X1_LOC_727/a_36_216# INVX1_LOC_117/A 0.00fF
C59375 NOR2X1_LOC_772/A INVX1_LOC_75/A 0.01fF
C59376 INVX1_LOC_7/A INVX1_LOC_315/Y 0.36fF
C59377 NOR2X1_LOC_657/B INVX1_LOC_22/A 0.00fF
C59378 NAND2X1_LOC_231/Y INVX1_LOC_46/A 0.03fF
C59379 NOR2X1_LOC_19/B INVX1_LOC_75/A 0.36fF
C59380 INVX1_LOC_290/A NOR2X1_LOC_141/a_36_216# 0.11fF
C59381 NAND2X1_LOC_30/Y INVX1_LOC_29/A 0.28fF
C59382 NAND2X1_LOC_852/Y INVX1_LOC_20/A 0.03fF
C59383 INVX1_LOC_155/A INVX1_LOC_9/A 0.18fF
C59384 VDD NAND2X1_LOC_451/Y 0.01fF
C59385 NOR2X1_LOC_589/A NAND2X1_LOC_642/Y 0.18fF
C59386 NOR2X1_LOC_641/B NOR2X1_LOC_814/A 0.03fF
C59387 INVX1_LOC_269/A NOR2X1_LOC_847/a_36_216# 0.01fF
C59388 NAND2X1_LOC_350/A NAND2X1_LOC_74/B 0.07fF
C59389 INVX1_LOC_208/A INVX1_LOC_76/A 0.01fF
C59390 NAND2X1_LOC_837/Y NOR2X1_LOC_88/a_36_216# 0.11fF
C59391 NOR2X1_LOC_264/Y INVX1_LOC_9/A 0.31fF
C59392 NOR2X1_LOC_594/Y NAND2X1_LOC_652/Y 0.00fF
C59393 NOR2X1_LOC_134/Y INVX1_LOC_29/A 0.03fF
C59394 NOR2X1_LOC_751/Y NOR2X1_LOC_814/A 0.07fF
C59395 NAND2X1_LOC_733/Y NOR2X1_LOC_11/Y 0.03fF
C59396 INVX1_LOC_286/Y NOR2X1_LOC_36/B 0.00fF
C59397 INVX1_LOC_49/A NOR2X1_LOC_634/A 0.03fF
C59398 NOR2X1_LOC_270/Y NAND2X1_LOC_475/Y 0.00fF
C59399 INVX1_LOC_83/A NAND2X1_LOC_649/B 0.01fF
C59400 NOR2X1_LOC_441/Y NAND2X1_LOC_74/B 0.16fF
C59401 INVX1_LOC_62/Y INVX1_LOC_27/Y 0.02fF
C59402 NAND2X1_LOC_852/Y NOR2X1_LOC_765/Y 0.03fF
C59403 NOR2X1_LOC_278/A INVX1_LOC_54/A 0.01fF
C59404 NOR2X1_LOC_67/A NOR2X1_LOC_99/a_36_216# 0.00fF
C59405 INVX1_LOC_30/A NOR2X1_LOC_1/Y 0.02fF
C59406 NOR2X1_LOC_433/A NOR2X1_LOC_127/a_36_216# 0.01fF
C59407 INVX1_LOC_8/A INVX1_LOC_46/Y 0.03fF
C59408 NOR2X1_LOC_599/A INVX1_LOC_12/A 0.03fF
C59409 NOR2X1_LOC_561/Y NAND2X1_LOC_211/Y 0.07fF
C59410 NOR2X1_LOC_574/A INVX1_LOC_291/A 0.07fF
C59411 NOR2X1_LOC_160/B INVX1_LOC_127/Y 0.00fF
C59412 INVX1_LOC_35/A NOR2X1_LOC_32/B 0.01fF
C59413 INVX1_LOC_182/Y NOR2X1_LOC_187/a_36_216# 0.00fF
C59414 INVX1_LOC_313/Y INVX1_LOC_188/Y 0.01fF
C59415 INVX1_LOC_137/Y INVX1_LOC_117/A 0.01fF
C59416 NOR2X1_LOC_419/Y INVX1_LOC_63/A 0.04fF
C59417 INVX1_LOC_266/Y INVX1_LOC_92/A 0.10fF
C59418 INVX1_LOC_136/A NAND2X1_LOC_807/B 0.18fF
C59419 NOR2X1_LOC_373/a_36_216# NAND2X1_LOC_477/Y 0.02fF
C59420 INVX1_LOC_230/Y NOR2X1_LOC_297/A 0.03fF
C59421 NAND2X1_LOC_773/a_36_24# NAND2X1_LOC_773/Y 0.00fF
C59422 NOR2X1_LOC_716/B INVX1_LOC_63/A 1.23fF
C59423 INVX1_LOC_58/A NAND2X1_LOC_391/Y 0.01fF
C59424 INVX1_LOC_18/A NAND2X1_LOC_254/Y 0.03fF
C59425 INVX1_LOC_192/A NOR2X1_LOC_450/B 0.00fF
C59426 INVX1_LOC_136/A NOR2X1_LOC_48/B 0.19fF
C59427 NOR2X1_LOC_65/B NAND2X1_LOC_773/Y 0.10fF
C59428 NOR2X1_LOC_454/Y INVX1_LOC_57/A 0.07fF
C59429 INVX1_LOC_2/A NOR2X1_LOC_58/Y 0.05fF
C59430 INVX1_LOC_33/A NAND2X1_LOC_782/B 0.01fF
C59431 INVX1_LOC_299/A INVX1_LOC_50/A 0.07fF
C59432 INVX1_LOC_161/Y NOR2X1_LOC_686/A 0.03fF
C59433 INVX1_LOC_49/A INVX1_LOC_29/A 0.18fF
C59434 NOR2X1_LOC_730/Y INVX1_LOC_274/A 0.47fF
C59435 NOR2X1_LOC_103/Y NOR2X1_LOC_72/Y 0.01fF
C59436 NAND2X1_LOC_565/B NOR2X1_LOC_235/Y 0.01fF
C59437 INPUT_0 NOR2X1_LOC_368/Y 0.00fF
C59438 INVX1_LOC_269/A INVX1_LOC_23/A 1.19fF
C59439 INPUT_0 NOR2X1_LOC_164/Y 0.03fF
C59440 INVX1_LOC_131/A INVX1_LOC_46/A 0.01fF
C59441 INVX1_LOC_25/Y NOR2X1_LOC_216/B 0.02fF
C59442 NOR2X1_LOC_567/B VDD 0.02fF
C59443 INVX1_LOC_172/A NAND2X1_LOC_254/Y 0.03fF
C59444 INVX1_LOC_249/A INVX1_LOC_283/A 0.01fF
C59445 D_INPUT_0 INVX1_LOC_118/Y 0.13fF
C59446 INVX1_LOC_16/A NOR2X1_LOC_831/B 0.03fF
C59447 INVX1_LOC_34/A NOR2X1_LOC_671/Y 0.01fF
C59448 NOR2X1_LOC_13/Y INVX1_LOC_32/A 0.03fF
C59449 NOR2X1_LOC_590/A NAND2X1_LOC_288/B 0.00fF
C59450 NAND2X1_LOC_35/Y NAND2X1_LOC_705/Y 0.03fF
C59451 NOR2X1_LOC_163/A INVX1_LOC_38/A 0.00fF
C59452 D_INPUT_7 NOR2X1_LOC_30/Y 0.03fF
C59453 INVX1_LOC_246/A NOR2X1_LOC_677/Y 0.02fF
C59454 NOR2X1_LOC_528/Y NAND2X1_LOC_620/a_36_24# 0.01fF
C59455 INVX1_LOC_264/Y NAND2X1_LOC_655/A 0.21fF
C59456 INVX1_LOC_64/A NAND2X1_LOC_724/A 0.07fF
C59457 NOR2X1_LOC_479/B NOR2X1_LOC_649/B 0.01fF
C59458 NOR2X1_LOC_311/a_36_216# NAND2X1_LOC_642/Y 0.00fF
C59459 INVX1_LOC_300/A INVX1_LOC_297/A 0.01fF
C59460 INPUT_0 INVX1_LOC_46/A 0.69fF
C59461 NOR2X1_LOC_68/A NAND2X1_LOC_223/A 0.03fF
C59462 INVX1_LOC_13/A NAND2X1_LOC_85/Y 0.01fF
C59463 NOR2X1_LOC_311/Y NAND2X1_LOC_649/B 0.17fF
C59464 NAND2X1_LOC_862/Y INVX1_LOC_54/A 0.01fF
C59465 NOR2X1_LOC_427/Y VDD 0.18fF
C59466 INVX1_LOC_24/A NAND2X1_LOC_471/Y 0.01fF
C59467 INVX1_LOC_25/Y NAND2X1_LOC_477/Y 0.08fF
C59468 NAND2X1_LOC_721/A NOR2X1_LOC_527/Y 0.06fF
C59469 INVX1_LOC_2/A INVX1_LOC_29/A 0.18fF
C59470 INVX1_LOC_225/Y INVX1_LOC_53/A -0.01fF
C59471 INVX1_LOC_132/A INVX1_LOC_4/A 0.47fF
C59472 INVX1_LOC_10/A NOR2X1_LOC_841/A 0.21fF
C59473 NOR2X1_LOC_655/B NAND2X1_LOC_74/B 0.15fF
C59474 INVX1_LOC_160/A INVX1_LOC_143/Y 0.45fF
C59475 NOR2X1_LOC_226/A INVX1_LOC_29/A 0.07fF
C59476 INVX1_LOC_21/A NAND2X1_LOC_780/Y 0.09fF
C59477 INVX1_LOC_15/Y INVX1_LOC_284/A 0.01fF
C59478 NOR2X1_LOC_130/A NOR2X1_LOC_832/a_36_216# 0.00fF
C59479 INVX1_LOC_147/A INVX1_LOC_38/A 0.00fF
C59480 NAND2X1_LOC_560/A INVX1_LOC_118/A 0.04fF
C59481 NAND2X1_LOC_581/Y D_INPUT_5 0.01fF
C59482 INVX1_LOC_11/A INVX1_LOC_298/A 0.03fF
C59483 NOR2X1_LOC_289/a_36_216# INVX1_LOC_272/A 0.01fF
C59484 NOR2X1_LOC_92/Y NOR2X1_LOC_792/a_36_216# 0.01fF
C59485 INVX1_LOC_24/A NAND2X1_LOC_616/a_36_24# 0.01fF
C59486 INVX1_LOC_64/A NOR2X1_LOC_45/Y 0.07fF
C59487 NAND2X1_LOC_9/Y NAND2X1_LOC_208/B 0.22fF
C59488 NOR2X1_LOC_2/Y INVX1_LOC_38/A 0.05fF
C59489 NOR2X1_LOC_590/A NOR2X1_LOC_405/Y 0.01fF
C59490 NOR2X1_LOC_191/B INVX1_LOC_26/A 0.00fF
C59491 NOR2X1_LOC_178/Y NOR2X1_LOC_160/B 0.20fF
C59492 INVX1_LOC_136/A NAND2X1_LOC_215/A 0.10fF
C59493 NAND2X1_LOC_642/Y INVX1_LOC_20/A 0.31fF
C59494 VDD NOR2X1_LOC_269/Y 0.15fF
C59495 NAND2X1_LOC_740/Y NAND2X1_LOC_537/a_36_24# 0.00fF
C59496 INVX1_LOC_225/A INVX1_LOC_4/A 0.14fF
C59497 INVX1_LOC_204/Y INVX1_LOC_174/A 0.03fF
C59498 INVX1_LOC_33/A NAND2X1_LOC_454/Y 0.13fF
C59499 NAND2X1_LOC_584/a_36_24# NOR2X1_LOC_467/A 0.00fF
C59500 INVX1_LOC_5/A NOR2X1_LOC_389/A 0.10fF
C59501 NOR2X1_LOC_92/Y INVX1_LOC_14/A 0.10fF
C59502 NOR2X1_LOC_717/B INVX1_LOC_63/A 0.03fF
C59503 NOR2X1_LOC_272/Y INVX1_LOC_150/Y 0.34fF
C59504 INVX1_LOC_91/A INVX1_LOC_117/A 0.14fF
C59505 INPUT_3 NOR2X1_LOC_649/Y 0.04fF
C59506 NOR2X1_LOC_741/a_36_216# INVX1_LOC_179/A 0.00fF
C59507 NAND2X1_LOC_175/B NAND2X1_LOC_175/Y 0.02fF
C59508 NOR2X1_LOC_351/a_36_216# INVX1_LOC_271/A 0.00fF
C59509 NAND2X1_LOC_579/A NAND2X1_LOC_561/B 0.41fF
C59510 NOR2X1_LOC_99/B INVX1_LOC_293/Y 0.09fF
C59511 NOR2X1_LOC_2/Y NOR2X1_LOC_51/A 0.03fF
C59512 INVX1_LOC_21/A NAND2X1_LOC_114/B 0.07fF
C59513 D_INPUT_1 INVX1_LOC_181/Y 0.04fF
C59514 INVX1_LOC_256/Y INVX1_LOC_32/A 0.10fF
C59515 INVX1_LOC_103/A INVX1_LOC_1/A 0.10fF
C59516 INVX1_LOC_279/A INVX1_LOC_263/Y 0.02fF
C59517 INVX1_LOC_75/A NOR2X1_LOC_216/B 0.16fF
C59518 NOR2X1_LOC_421/Y NOR2X1_LOC_422/Y 0.06fF
C59519 INVX1_LOC_76/A NAND2X1_LOC_211/Y 0.10fF
C59520 INVX1_LOC_77/A INVX1_LOC_57/A 8.63fF
C59521 INVX1_LOC_266/A NOR2X1_LOC_541/Y 0.01fF
C59522 INVX1_LOC_45/A INVX1_LOC_50/Y 0.03fF
C59523 INVX1_LOC_21/A INVX1_LOC_141/Y 0.03fF
C59524 INVX1_LOC_16/A NOR2X1_LOC_270/a_36_216# 0.00fF
C59525 NOR2X1_LOC_99/B NAND2X1_LOC_74/B 0.08fF
C59526 NOR2X1_LOC_286/Y NOR2X1_LOC_241/A 0.05fF
C59527 INVX1_LOC_279/A INVX1_LOC_42/A 0.07fF
C59528 INVX1_LOC_21/A INVX1_LOC_312/Y 0.04fF
C59529 INVX1_LOC_21/A NOR2X1_LOC_294/Y 0.06fF
C59530 NOR2X1_LOC_400/B NOR2X1_LOC_6/B 0.06fF
C59531 NOR2X1_LOC_613/Y INVX1_LOC_30/A 0.05fF
C59532 INVX1_LOC_298/Y INVX1_LOC_2/A 0.03fF
C59533 INVX1_LOC_36/A NAND2X1_LOC_816/a_36_24# 0.00fF
C59534 INVX1_LOC_11/A NAND2X1_LOC_793/Y 0.00fF
C59535 INVX1_LOC_5/A INVX1_LOC_62/Y 0.07fF
C59536 INVX1_LOC_238/A INVX1_LOC_229/A 1.28fF
C59537 INPUT_1 INVX1_LOC_29/A 4.42fF
C59538 NOR2X1_LOC_816/a_36_216# INVX1_LOC_18/A 0.00fF
C59539 INVX1_LOC_104/A NOR2X1_LOC_383/B 0.16fF
C59540 INVX1_LOC_125/Y INVX1_LOC_92/A 0.82fF
C59541 NAND2X1_LOC_55/a_36_24# INVX1_LOC_25/A 0.00fF
C59542 INVX1_LOC_5/A NOR2X1_LOC_596/A 0.10fF
C59543 INVX1_LOC_224/Y NOR2X1_LOC_6/B 0.05fF
C59544 INVX1_LOC_269/A INVX1_LOC_31/A 0.08fF
C59545 NOR2X1_LOC_151/Y INVX1_LOC_63/A 0.14fF
C59546 INVX1_LOC_298/Y NOR2X1_LOC_226/A 0.00fF
C59547 NOR2X1_LOC_440/Y INVX1_LOC_47/Y 0.19fF
C59548 INVX1_LOC_181/Y NOR2X1_LOC_652/Y 0.14fF
C59549 NOR2X1_LOC_751/A NOR2X1_LOC_814/A 0.02fF
C59550 NOR2X1_LOC_232/Y INVX1_LOC_31/A 0.02fF
C59551 INVX1_LOC_132/A INVX1_LOC_64/A 0.07fF
C59552 INVX1_LOC_266/A INVX1_LOC_45/A 0.03fF
C59553 INVX1_LOC_20/A NOR2X1_LOC_271/Y 0.03fF
C59554 INVX1_LOC_316/Y NOR2X1_LOC_825/a_36_216# 0.00fF
C59555 NAND2X1_LOC_9/Y INVX1_LOC_34/A 0.03fF
C59556 INVX1_LOC_266/A NOR2X1_LOC_568/A 0.56fF
C59557 NAND2X1_LOC_563/Y D_INPUT_1 0.11fF
C59558 INVX1_LOC_124/A INVX1_LOC_57/A 0.03fF
C59559 INVX1_LOC_233/A INVX1_LOC_34/A 0.07fF
C59560 INVX1_LOC_223/Y NOR2X1_LOC_500/A 0.37fF
C59561 INVX1_LOC_41/A NOR2X1_LOC_489/B 0.01fF
C59562 NOR2X1_LOC_389/A NAND2X1_LOC_337/B 0.10fF
C59563 NOR2X1_LOC_84/A NOR2X1_LOC_392/Y 0.07fF
C59564 NOR2X1_LOC_15/Y INVX1_LOC_72/A 0.04fF
C59565 INVX1_LOC_21/A NOR2X1_LOC_546/B 0.02fF
C59566 INVX1_LOC_292/A NOR2X1_LOC_794/B 0.01fF
C59567 INPUT_0 NOR2X1_LOC_68/Y 0.01fF
C59568 INVX1_LOC_256/A NOR2X1_LOC_231/B 0.08fF
C59569 NOR2X1_LOC_45/B INVX1_LOC_113/A 0.04fF
C59570 INVX1_LOC_182/Y INVX1_LOC_263/Y 0.00fF
C59571 NAND2X1_LOC_218/B INVX1_LOC_27/A 1.88fF
C59572 NOR2X1_LOC_88/Y NAND2X1_LOC_655/A 0.07fF
C59573 NOR2X1_LOC_817/Y INVX1_LOC_40/Y 0.03fF
C59574 NOR2X1_LOC_488/Y NOR2X1_LOC_693/Y 0.02fF
C59575 NAND2X1_LOC_35/Y NOR2X1_LOC_690/A 0.22fF
C59576 NOR2X1_LOC_332/A NOR2X1_LOC_38/B 0.09fF
C59577 INVX1_LOC_266/Y INVX1_LOC_53/A 0.22fF
C59578 INVX1_LOC_33/Y NOR2X1_LOC_536/A 0.03fF
C59579 INVX1_LOC_279/A INVX1_LOC_78/A 0.07fF
C59580 INVX1_LOC_17/A D_INPUT_7 0.00fF
C59581 NOR2X1_LOC_441/Y NOR2X1_LOC_276/Y 0.39fF
C59582 INVX1_LOC_27/A NOR2X1_LOC_577/Y 0.03fF
C59583 INVX1_LOC_182/Y INVX1_LOC_42/A 0.03fF
C59584 NOR2X1_LOC_502/Y NAND2X1_LOC_510/A 0.03fF
C59585 INVX1_LOC_50/A INVX1_LOC_52/A 0.02fF
C59586 INVX1_LOC_21/A INVX1_LOC_275/A 0.12fF
C59587 NOR2X1_LOC_173/Y NOR2X1_LOC_433/A 0.07fF
C59588 NOR2X1_LOC_401/B NAND2X1_LOC_860/A 0.02fF
C59589 INPUT_0 NOR2X1_LOC_671/Y 0.03fF
C59590 INVX1_LOC_266/A INVX1_LOC_71/A 0.06fF
C59591 INVX1_LOC_84/A NAND2X1_LOC_655/A 0.03fF
C59592 INVX1_LOC_5/A NOR2X1_LOC_844/A 0.03fF
C59593 INVX1_LOC_136/A NAND2X1_LOC_350/A 0.10fF
C59594 NOR2X1_LOC_772/Y NAND2X1_LOC_474/Y 0.27fF
C59595 NOR2X1_LOC_402/a_36_216# NAND2X1_LOC_860/A 0.01fF
C59596 NAND2X1_LOC_364/A INVX1_LOC_150/Y 0.09fF
C59597 NOR2X1_LOC_74/A INVX1_LOC_102/A 0.14fF
C59598 INVX1_LOC_36/A NOR2X1_LOC_644/B 0.01fF
C59599 NOR2X1_LOC_287/a_36_216# NOR2X1_LOC_798/A 0.00fF
C59600 NAND2X1_LOC_733/Y NOR2X1_LOC_599/A 0.03fF
C59601 INVX1_LOC_22/A INVX1_LOC_271/A 0.09fF
C59602 NOR2X1_LOC_473/B NOR2X1_LOC_334/Y 0.10fF
C59603 NOR2X1_LOC_479/B NOR2X1_LOC_476/B 0.26fF
C59604 VDD NOR2X1_LOC_79/Y 0.00fF
C59605 INVX1_LOC_14/Y NOR2X1_LOC_155/A 0.01fF
C59606 NOR2X1_LOC_500/Y NOR2X1_LOC_493/a_36_216# 0.03fF
C59607 NOR2X1_LOC_349/B NOR2X1_LOC_342/B 0.02fF
C59608 NAND2X1_LOC_644/a_36_24# NOR2X1_LOC_409/B 0.00fF
C59609 INVX1_LOC_52/Y INVX1_LOC_63/Y 0.01fF
C59610 INVX1_LOC_136/A NOR2X1_LOC_441/Y 0.01fF
C59611 NOR2X1_LOC_240/Y NOR2X1_LOC_78/B 0.12fF
C59612 INVX1_LOC_90/A NOR2X1_LOC_36/A 0.13fF
C59613 NOR2X1_LOC_181/A INVX1_LOC_63/A 0.01fF
C59614 NOR2X1_LOC_92/Y INVX1_LOC_217/Y -0.09fF
C59615 INVX1_LOC_233/A NAND2X1_LOC_858/a_36_24# 0.00fF
C59616 NOR2X1_LOC_173/Y NOR2X1_LOC_52/B 0.03fF
C59617 INVX1_LOC_186/A INVX1_LOC_69/A 0.03fF
C59618 NOR2X1_LOC_165/a_36_216# NOR2X1_LOC_48/B 0.00fF
C59619 INVX1_LOC_41/A INVX1_LOC_14/A 0.22fF
C59620 NOR2X1_LOC_52/Y INVX1_LOC_30/A 0.00fF
C59621 INVX1_LOC_5/A NOR2X1_LOC_220/A 0.10fF
C59622 NAND2X1_LOC_510/A NAND2X1_LOC_508/a_36_24# 0.03fF
C59623 INVX1_LOC_11/Y INVX1_LOC_163/Y 0.03fF
C59624 NAND2X1_LOC_151/a_36_24# NOR2X1_LOC_577/Y 0.00fF
C59625 INVX1_LOC_201/Y INVX1_LOC_14/A 0.20fF
C59626 NOR2X1_LOC_270/Y INVX1_LOC_30/A 0.01fF
C59627 INVX1_LOC_27/A NOR2X1_LOC_346/B 0.07fF
C59628 NAND2X1_LOC_725/A NAND2X1_LOC_735/B 0.05fF
C59629 INVX1_LOC_33/Y NAND2X1_LOC_780/a_36_24# 0.00fF
C59630 NOR2X1_LOC_434/Y NOR2X1_LOC_516/B 0.03fF
C59631 NAND2X1_LOC_53/Y NOR2X1_LOC_147/B 0.12fF
C59632 INVX1_LOC_91/A NOR2X1_LOC_460/A 0.01fF
C59633 INVX1_LOC_119/A NAND2X1_LOC_537/Y 0.30fF
C59634 INVX1_LOC_14/A NAND2X1_LOC_477/A 0.10fF
C59635 NAND2X1_LOC_358/B NAND2X1_LOC_358/Y 0.12fF
C59636 INVX1_LOC_93/A INVX1_LOC_25/Y 0.07fF
C59637 NOR2X1_LOC_331/B NAND2X1_LOC_792/a_36_24# 0.01fF
C59638 NOR2X1_LOC_34/B NOR2X1_LOC_516/B 0.01fF
C59639 NOR2X1_LOC_214/B INVX1_LOC_23/A 0.00fF
C59640 NOR2X1_LOC_739/Y NOR2X1_LOC_731/A 0.00fF
C59641 NOR2X1_LOC_103/Y NOR2X1_LOC_6/B 0.03fF
C59642 INVX1_LOC_204/Y NOR2X1_LOC_589/A 0.03fF
C59643 INVX1_LOC_50/A NOR2X1_LOC_166/Y 0.02fF
C59644 NOR2X1_LOC_15/Y NAND2X1_LOC_338/B 0.15fF
C59645 INVX1_LOC_91/A INVX1_LOC_3/Y 0.01fF
C59646 NOR2X1_LOC_276/Y NOR2X1_LOC_142/Y 0.09fF
C59647 VDD NOR2X1_LOC_36/B 0.41fF
C59648 INVX1_LOC_248/A NAND2X1_LOC_780/Y 0.02fF
C59649 INVX1_LOC_27/A INVX1_LOC_22/A 0.11fF
C59650 NOR2X1_LOC_586/Y INVX1_LOC_29/A 0.02fF
C59651 NOR2X1_LOC_824/A INVX1_LOC_22/A 0.02fF
C59652 NOR2X1_LOC_346/Y NOR2X1_LOC_861/Y 0.04fF
C59653 NOR2X1_LOC_139/Y INVX1_LOC_15/A 0.08fF
C59654 NAND2X1_LOC_655/A INVX1_LOC_15/A 0.07fF
C59655 INVX1_LOC_48/Y NOR2X1_LOC_121/a_36_216# 0.01fF
C59656 NOR2X1_LOC_514/A NAND2X1_LOC_139/A 0.01fF
C59657 NOR2X1_LOC_117/a_36_216# INVX1_LOC_54/A 0.01fF
C59658 NOR2X1_LOC_355/B NOR2X1_LOC_334/Y 0.01fF
C59659 NOR2X1_LOC_522/Y NAND2X1_LOC_837/Y 0.03fF
C59660 NOR2X1_LOC_99/B NOR2X1_LOC_845/a_36_216# 0.01fF
C59661 INVX1_LOC_237/A INVX1_LOC_22/A 0.20fF
C59662 NOR2X1_LOC_82/A NAND2X1_LOC_360/B 0.09fF
C59663 NAND2X1_LOC_642/Y INVX1_LOC_4/A 0.18fF
C59664 NAND2X1_LOC_154/Y INVX1_LOC_63/Y 0.01fF
C59665 INVX1_LOC_265/A INVX1_LOC_30/A 0.01fF
C59666 NAND2X1_LOC_468/B INVX1_LOC_15/A 0.05fF
C59667 NOR2X1_LOC_837/B NOR2X1_LOC_837/Y 0.03fF
C59668 INVX1_LOC_214/Y INVX1_LOC_161/Y 0.05fF
C59669 NOR2X1_LOC_458/B NOR2X1_LOC_457/A 0.03fF
C59670 NOR2X1_LOC_778/B NOR2X1_LOC_787/a_36_216# 0.00fF
C59671 INVX1_LOC_21/A NAND2X1_LOC_656/Y 0.12fF
C59672 INVX1_LOC_136/A NOR2X1_LOC_142/Y 0.07fF
C59673 NOR2X1_LOC_68/A INVX1_LOC_33/A 0.27fF
C59674 NOR2X1_LOC_78/B INVX1_LOC_225/Y 0.17fF
C59675 INVX1_LOC_45/A NOR2X1_LOC_6/B 0.00fF
C59676 INVX1_LOC_30/A NOR2X1_LOC_180/Y 0.10fF
C59677 NOR2X1_LOC_441/Y NOR2X1_LOC_111/a_36_216# 0.01fF
C59678 NOR2X1_LOC_6/B NOR2X1_LOC_568/A -0.00fF
C59679 NOR2X1_LOC_381/a_36_216# NOR2X1_LOC_660/Y 0.00fF
C59680 NOR2X1_LOC_514/A NAND2X1_LOC_139/a_36_24# 0.00fF
C59681 NAND2X1_LOC_361/Y NAND2X1_LOC_656/A 0.10fF
C59682 INVX1_LOC_206/Y NOR2X1_LOC_383/B 0.01fF
C59683 NOR2X1_LOC_232/Y NAND2X1_LOC_859/Y 0.00fF
C59684 INVX1_LOC_193/A NAND2X1_LOC_259/a_36_24# 0.00fF
C59685 INVX1_LOC_254/Y INVX1_LOC_303/A 0.02fF
C59686 NAND2X1_LOC_9/Y INPUT_0 0.13fF
C59687 NOR2X1_LOC_667/A INVX1_LOC_141/Y 0.03fF
C59688 NAND2X1_LOC_169/Y INVX1_LOC_28/A 0.02fF
C59689 INVX1_LOC_30/Y NOR2X1_LOC_103/Y 0.04fF
C59690 INVX1_LOC_2/A NAND2X1_LOC_721/B 0.00fF
C59691 INVX1_LOC_41/A NAND2X1_LOC_84/Y 0.03fF
C59692 INVX1_LOC_90/A NAND2X1_LOC_474/Y 0.03fF
C59693 INVX1_LOC_118/A INVX1_LOC_29/A 1.82fF
C59694 INVX1_LOC_89/A NAND2X1_LOC_473/A 0.01fF
C59695 NAND2X1_LOC_555/Y NAND2X1_LOC_672/B 0.02fF
C59696 NAND2X1_LOC_563/A INVX1_LOC_31/A 0.12fF
C59697 INVX1_LOC_21/A NAND2X1_LOC_638/Y 0.18fF
C59698 INVX1_LOC_248/A INVX1_LOC_141/Y 0.84fF
C59699 INVX1_LOC_217/Y NAND2X1_LOC_837/Y 0.01fF
C59700 NAND2X1_LOC_729/Y INVX1_LOC_240/A 0.53fF
C59701 INVX1_LOC_233/A INPUT_0 0.25fF
C59702 NOR2X1_LOC_389/B NAND2X1_LOC_474/Y 0.01fF
C59703 NOR2X1_LOC_217/a_36_216# NOR2X1_LOC_561/Y 0.01fF
C59704 INVX1_LOC_99/Y INVX1_LOC_75/A 0.02fF
C59705 NOR2X1_LOC_667/A INVX1_LOC_312/Y 0.03fF
C59706 NOR2X1_LOC_226/A NAND2X1_LOC_721/B 0.03fF
C59707 INVX1_LOC_248/A INVX1_LOC_312/Y -0.01fF
C59708 NOR2X1_LOC_360/Y INVX1_LOC_177/A 0.03fF
C59709 INVX1_LOC_136/A NOR2X1_LOC_655/B 0.10fF
C59710 INVX1_LOC_19/A INVX1_LOC_92/A 0.80fF
C59711 NAND2X1_LOC_784/a_36_24# NAND2X1_LOC_807/Y -0.01fF
C59712 NAND2X1_LOC_563/Y D_INPUT_2 0.12fF
C59713 NAND2X1_LOC_508/A NAND2X1_LOC_473/A 0.07fF
C59714 NOR2X1_LOC_458/a_36_216# INVX1_LOC_96/A -0.00fF
C59715 INVX1_LOC_58/A INVX1_LOC_91/A 0.67fF
C59716 NOR2X1_LOC_15/Y INVX1_LOC_313/Y 0.01fF
C59717 NOR2X1_LOC_778/B INVX1_LOC_18/A 0.03fF
C59718 NOR2X1_LOC_78/A INVX1_LOC_129/A 0.00fF
C59719 NAND2X1_LOC_24/a_36_24# NAND2X1_LOC_555/Y 0.00fF
C59720 NOR2X1_LOC_66/Y INVX1_LOC_84/A 0.18fF
C59721 NAND2X1_LOC_553/A INPUT_0 0.14fF
C59722 NOR2X1_LOC_78/B INVX1_LOC_72/Y 0.01fF
C59723 INVX1_LOC_224/Y NOR2X1_LOC_124/A 0.02fF
C59724 INVX1_LOC_84/A NOR2X1_LOC_820/B 0.04fF
C59725 NOR2X1_LOC_443/a_36_216# D_INPUT_0 0.02fF
C59726 NOR2X1_LOC_68/A INVX1_LOC_40/A 0.07fF
C59727 NOR2X1_LOC_798/A INPUT_0 0.08fF
C59728 INVX1_LOC_58/A INVX1_LOC_11/Y 0.03fF
C59729 D_INPUT_1 NOR2X1_LOC_675/A 0.01fF
C59730 VDD INVX1_LOC_26/A 1.23fF
C59731 INVX1_LOC_4/A NOR2X1_LOC_271/Y 0.03fF
C59732 NAND2X1_LOC_53/Y INVX1_LOC_90/A 0.07fF
C59733 INVX1_LOC_230/Y NOR2X1_LOC_130/A 0.71fF
C59734 INVX1_LOC_206/A NOR2X1_LOC_577/Y 0.01fF
C59735 NOR2X1_LOC_690/A NOR2X1_LOC_234/Y 0.14fF
C59736 NOR2X1_LOC_160/B NAND2X1_LOC_45/Y 0.10fF
C59737 INVX1_LOC_60/A INVX1_LOC_8/A 0.03fF
C59738 INVX1_LOC_12/A NOR2X1_LOC_841/A 0.10fF
C59739 INVX1_LOC_49/Y INVX1_LOC_119/Y 0.01fF
C59740 INVX1_LOC_7/Y INVX1_LOC_48/A 0.09fF
C59741 INVX1_LOC_41/A NOR2X1_LOC_612/B 0.27fF
C59742 INVX1_LOC_31/A NOR2X1_LOC_814/Y 0.23fF
C59743 NOR2X1_LOC_598/B NAND2X1_LOC_212/Y 0.03fF
C59744 NAND2X1_LOC_647/B INVX1_LOC_54/A 0.01fF
C59745 NOR2X1_LOC_720/B NAND2X1_LOC_667/a_36_24# 0.02fF
C59746 INVX1_LOC_21/A INVX1_LOC_78/Y 0.03fF
C59747 NOR2X1_LOC_34/B INVX1_LOC_315/Y 0.01fF
C59748 INVX1_LOC_38/A NOR2X1_LOC_36/A 0.13fF
C59749 INVX1_LOC_248/Y INVX1_LOC_91/A 0.10fF
C59750 NOR2X1_LOC_623/B NOR2X1_LOC_640/Y 0.01fF
C59751 INVX1_LOC_2/A INVX1_LOC_8/A 0.10fF
C59752 INVX1_LOC_207/A INVX1_LOC_280/Y 0.03fF
C59753 NOR2X1_LOC_590/A NOR2X1_LOC_644/A 0.03fF
C59754 NOR2X1_LOC_790/B NOR2X1_LOC_35/Y 0.03fF
C59755 NAND2X1_LOC_640/Y NAND2X1_LOC_850/Y -0.00fF
C59756 INVX1_LOC_249/A INVX1_LOC_22/A 0.03fF
C59757 NOR2X1_LOC_351/Y NAND2X1_LOC_454/Y 0.01fF
C59758 NOR2X1_LOC_536/A INVX1_LOC_23/Y 1.06fF
C59759 NOR2X1_LOC_445/Y NOR2X1_LOC_203/Y 0.05fF
C59760 INVX1_LOC_136/A NOR2X1_LOC_99/B 0.10fF
C59761 NOR2X1_LOC_255/Y VDD -0.00fF
C59762 NOR2X1_LOC_510/Y NOR2X1_LOC_269/Y 0.08fF
C59763 NOR2X1_LOC_75/Y NOR2X1_LOC_742/A -0.00fF
C59764 INVX1_LOC_30/Y INVX1_LOC_71/A 0.10fF
C59765 NOR2X1_LOC_226/A INVX1_LOC_8/A 0.01fF
C59766 NOR2X1_LOC_431/a_36_216# NOR2X1_LOC_561/Y 0.01fF
C59767 NOR2X1_LOC_598/B D_INPUT_3 0.08fF
C59768 INVX1_LOC_227/A INVX1_LOC_45/Y 0.08fF
C59769 INVX1_LOC_269/A INVX1_LOC_6/A 0.01fF
C59770 INVX1_LOC_12/Y INVX1_LOC_23/A 0.11fF
C59771 NOR2X1_LOC_598/B INVX1_LOC_14/Y 0.09fF
C59772 NOR2X1_LOC_675/A NOR2X1_LOC_652/Y 0.01fF
C59773 INVX1_LOC_239/A INVX1_LOC_167/Y 0.16fF
C59774 NOR2X1_LOC_51/A NOR2X1_LOC_36/A 0.40fF
C59775 NOR2X1_LOC_281/Y INVX1_LOC_118/A 0.06fF
C59776 NOR2X1_LOC_716/B INVX1_LOC_1/Y 0.07fF
C59777 NOR2X1_LOC_78/A NOR2X1_LOC_440/B 0.04fF
C59778 NOR2X1_LOC_107/Y NOR2X1_LOC_721/Y 0.06fF
C59779 NAND2X1_LOC_555/Y INVX1_LOC_82/Y 0.04fF
C59780 NAND2X1_LOC_63/Y INVX1_LOC_29/A 0.13fF
C59781 INVX1_LOC_5/A NAND2X1_LOC_469/B 0.00fF
C59782 INVX1_LOC_223/A NOR2X1_LOC_356/A 0.47fF
C59783 INVX1_LOC_314/Y NOR2X1_LOC_383/a_36_216# 0.00fF
C59784 NAND2X1_LOC_634/Y INPUT_1 0.04fF
C59785 D_INPUT_0 NAND2X1_LOC_79/Y 0.06fF
C59786 NOR2X1_LOC_78/B INVX1_LOC_266/Y 0.06fF
C59787 INVX1_LOC_226/Y NOR2X1_LOC_392/B 0.01fF
C59788 NOR2X1_LOC_637/B NOR2X1_LOC_561/Y 0.00fF
C59789 NAND2X1_LOC_190/Y NOR2X1_LOC_187/a_36_216# 0.00fF
C59790 INVX1_LOC_292/A NOR2X1_LOC_188/A 0.08fF
C59791 INVX1_LOC_203/A INVX1_LOC_3/Y 0.10fF
C59792 INVX1_LOC_57/A INVX1_LOC_9/A 0.25fF
C59793 NAND2X1_LOC_93/B INVX1_LOC_23/Y 0.02fF
C59794 NOR2X1_LOC_561/Y INVX1_LOC_155/A 0.01fF
C59795 INVX1_LOC_136/A INVX1_LOC_182/A 0.39fF
C59796 NOR2X1_LOC_643/Y INVX1_LOC_83/A 0.13fF
C59797 NAND2X1_LOC_357/B INVX1_LOC_16/A 0.07fF
C59798 NOR2X1_LOC_172/Y INVX1_LOC_10/A 0.01fF
C59799 NOR2X1_LOC_361/B NOR2X1_LOC_269/Y 0.00fF
C59800 NOR2X1_LOC_256/a_36_216# INPUT_1 0.00fF
C59801 INVX1_LOC_5/A NAND2X1_LOC_212/a_36_24# 0.00fF
C59802 INVX1_LOC_26/Y INVX1_LOC_92/A 0.08fF
C59803 INVX1_LOC_228/A INPUT_1 0.20fF
C59804 NOR2X1_LOC_84/Y INVX1_LOC_56/Y 0.06fF
C59805 NOR2X1_LOC_468/a_36_216# NOR2X1_LOC_557/Y 0.00fF
C59806 INVX1_LOC_87/A NAND2X1_LOC_572/B 0.01fF
C59807 NAND2X1_LOC_338/B INVX1_LOC_226/A 0.03fF
C59808 NOR2X1_LOC_419/Y NOR2X1_LOC_559/a_36_216# 0.00fF
C59809 INVX1_LOC_2/A INVX1_LOC_151/Y 0.03fF
C59810 NOR2X1_LOC_62/a_36_216# NOR2X1_LOC_709/A 0.01fF
C59811 NAND2X1_LOC_200/B NOR2X1_LOC_346/B 0.01fF
C59812 INVX1_LOC_179/A NOR2X1_LOC_632/a_36_216# 0.00fF
C59813 NOR2X1_LOC_772/B NOR2X1_LOC_440/a_36_216# 0.00fF
C59814 NAND2X1_LOC_736/B INVX1_LOC_229/Y 0.05fF
C59815 INVX1_LOC_223/A NOR2X1_LOC_74/A 0.03fF
C59816 NAND2X1_LOC_162/A NAND2X1_LOC_451/Y 0.02fF
C59817 INVX1_LOC_34/A NOR2X1_LOC_700/Y 0.00fF
C59818 NOR2X1_LOC_392/B INVX1_LOC_10/A 0.03fF
C59819 INVX1_LOC_229/Y GATE_811 0.02fF
C59820 INVX1_LOC_215/Y INVX1_LOC_91/A 0.05fF
C59821 NOR2X1_LOC_629/B INVX1_LOC_234/A 0.02fF
C59822 NAND2X1_LOC_218/B NOR2X1_LOC_19/B 0.12fF
C59823 INVX1_LOC_249/A NOR2X1_LOC_735/Y 0.01fF
C59824 NOR2X1_LOC_68/A NOR2X1_LOC_323/Y 0.03fF
C59825 INVX1_LOC_150/Y NOR2X1_LOC_113/A 0.36fF
C59826 INVX1_LOC_1/A INVX1_LOC_143/Y 2.76fF
C59827 NOR2X1_LOC_103/Y NOR2X1_LOC_124/A 0.02fF
C59828 INVX1_LOC_150/Y NOR2X1_LOC_405/A 0.81fF
C59829 INVX1_LOC_278/Y NOR2X1_LOC_165/Y 0.00fF
C59830 NAND2X1_LOC_564/B INVX1_LOC_256/Y 0.04fF
C59831 NOR2X1_LOC_773/Y NAND2X1_LOC_863/B 0.03fF
C59832 INVX1_LOC_89/A NOR2X1_LOC_486/B 0.24fF
C59833 INVX1_LOC_33/A NOR2X1_LOC_163/A 0.31fF
C59834 NAND2X1_LOC_265/a_36_24# INVX1_LOC_92/A 0.00fF
C59835 INVX1_LOC_212/A INVX1_LOC_75/A 0.03fF
C59836 NOR2X1_LOC_777/B NOR2X1_LOC_839/B 0.06fF
C59837 INVX1_LOC_23/Y INVX1_LOC_3/A 0.23fF
C59838 INVX1_LOC_89/A NOR2X1_LOC_516/Y 0.03fF
C59839 NOR2X1_LOC_666/A VDD 0.20fF
C59840 INVX1_LOC_255/Y NAND2X1_LOC_819/Y 0.01fF
C59841 INVX1_LOC_43/Y NAND2X1_LOC_642/Y 0.00fF
C59842 INVX1_LOC_8/A INPUT_1 0.32fF
C59843 INVX1_LOC_83/A INVX1_LOC_266/Y 0.05fF
C59844 INVX1_LOC_75/A NOR2X1_LOC_303/Y 0.03fF
C59845 NAND2X1_LOC_608/a_36_24# INVX1_LOC_9/A 0.00fF
C59846 NOR2X1_LOC_392/Y NOR2X1_LOC_78/Y 0.06fF
C59847 INVX1_LOC_34/A NAND2X1_LOC_842/B 0.03fF
C59848 NOR2X1_LOC_561/A NAND2X1_LOC_474/Y 0.05fF
C59849 NOR2X1_LOC_385/Y INVX1_LOC_231/Y 0.02fF
C59850 INVX1_LOC_17/A INVX1_LOC_2/Y 1.45fF
C59851 NOR2X1_LOC_382/Y NOR2X1_LOC_45/B 0.09fF
C59852 NOR2X1_LOC_356/A INVX1_LOC_149/Y 0.00fF
C59853 NAND2X1_LOC_323/B NOR2X1_LOC_97/B 0.00fF
C59854 D_INPUT_0 NOR2X1_LOC_520/A 0.07fF
C59855 NOR2X1_LOC_38/B INVX1_LOC_42/A 0.06fF
C59856 INVX1_LOC_53/A NAND2X1_LOC_288/A 0.08fF
C59857 NOR2X1_LOC_75/Y INVX1_LOC_139/A 0.01fF
C59858 INVX1_LOC_75/A NOR2X1_LOC_708/B 0.04fF
C59859 NOR2X1_LOC_107/Y VDD 0.25fF
C59860 NAND2X1_LOC_371/a_36_24# NOR2X1_LOC_337/Y -0.00fF
C59861 NAND2X1_LOC_357/B INVX1_LOC_28/A 0.12fF
C59862 INVX1_LOC_17/A INVX1_LOC_37/Y 0.16fF
C59863 INVX1_LOC_45/A NOR2X1_LOC_124/A 0.03fF
C59864 INVX1_LOC_36/A INVX1_LOC_187/A 0.01fF
C59865 NAND2X1_LOC_782/B INVX1_LOC_275/Y 0.20fF
C59866 INVX1_LOC_225/Y INVX1_LOC_46/A 0.09fF
C59867 INVX1_LOC_75/A NOR2X1_LOC_254/Y 0.03fF
C59868 INVX1_LOC_135/A INVX1_LOC_197/Y 0.66fF
C59869 NOR2X1_LOC_739/Y INVX1_LOC_117/A 0.00fF
C59870 INVX1_LOC_58/A INVX1_LOC_203/A 0.03fF
C59871 NOR2X1_LOC_636/B NAND2X1_LOC_639/A 0.37fF
C59872 NAND2X1_LOC_796/B INVX1_LOC_185/A -0.00fF
C59873 NOR2X1_LOC_266/a_36_216# INVX1_LOC_95/A -0.00fF
C59874 NOR2X1_LOC_89/A NOR2X1_LOC_693/a_36_216# 0.02fF
C59875 NAND2X1_LOC_465/a_36_24# INVX1_LOC_23/A 0.00fF
C59876 NOR2X1_LOC_292/Y NOR2X1_LOC_557/Y 0.02fF
C59877 NOR2X1_LOC_596/A NOR2X1_LOC_187/a_36_216# 0.02fF
C59878 INVX1_LOC_141/A VDD -0.00fF
C59879 NOR2X1_LOC_219/B INVX1_LOC_311/A 0.24fF
C59880 INVX1_LOC_96/A INVX1_LOC_71/A 1.46fF
C59881 NAND2X1_LOC_466/Y INVX1_LOC_144/A 0.03fF
C59882 NOR2X1_LOC_82/Y NOR2X1_LOC_71/Y 0.09fF
C59883 NOR2X1_LOC_477/a_36_216# INVX1_LOC_37/A 0.00fF
C59884 INVX1_LOC_162/Y NOR2X1_LOC_74/A 0.17fF
C59885 NOR2X1_LOC_68/A NOR2X1_LOC_486/Y 0.08fF
C59886 INVX1_LOC_73/A NOR2X1_LOC_709/A 0.07fF
C59887 INVX1_LOC_90/A NOR2X1_LOC_500/Y 0.07fF
C59888 INVX1_LOC_226/Y INVX1_LOC_90/A 0.03fF
C59889 NAND2X1_LOC_53/Y INVX1_LOC_38/A 0.10fF
C59890 INVX1_LOC_30/Y NOR2X1_LOC_123/B 0.02fF
C59891 NOR2X1_LOC_772/B INVX1_LOC_84/A 0.07fF
C59892 INVX1_LOC_53/A INVX1_LOC_19/A 0.19fF
C59893 INVX1_LOC_54/Y INVX1_LOC_75/A 0.01fF
C59894 NAND2X1_LOC_733/B NAND2X1_LOC_560/A 0.25fF
C59895 NOR2X1_LOC_210/A INVX1_LOC_295/A 0.02fF
C59896 INVX1_LOC_30/Y NOR2X1_LOC_749/Y 0.01fF
C59897 INVX1_LOC_48/Y NOR2X1_LOC_101/a_36_216# 0.01fF
C59898 NOR2X1_LOC_91/Y INVX1_LOC_20/A 0.34fF
C59899 NOR2X1_LOC_122/A INVX1_LOC_92/A 0.03fF
C59900 INVX1_LOC_43/Y NOR2X1_LOC_271/Y 1.41fF
C59901 INVX1_LOC_13/Y INVX1_LOC_84/A 0.07fF
C59902 NOR2X1_LOC_316/Y NOR2X1_LOC_9/Y -0.01fF
C59903 NOR2X1_LOC_820/A VDD 0.24fF
C59904 NAND2X1_LOC_463/B NOR2X1_LOC_399/Y 0.00fF
C59905 NOR2X1_LOC_245/a_36_216# D_INPUT_0 0.02fF
C59906 NOR2X1_LOC_276/B VDD -0.00fF
C59907 NOR2X1_LOC_292/Y INVX1_LOC_143/A 0.01fF
C59908 INVX1_LOC_90/A INVX1_LOC_10/A 0.13fF
C59909 NOR2X1_LOC_518/Y NAND2X1_LOC_804/Y 0.14fF
C59910 NAND2X1_LOC_849/A INVX1_LOC_16/A 0.03fF
C59911 NOR2X1_LOC_718/B NOR2X1_LOC_562/B 0.02fF
C59912 NOR2X1_LOC_389/B INVX1_LOC_10/A 0.08fF
C59913 INVX1_LOC_11/A NAND2X1_LOC_798/B 0.07fF
C59914 NAND2X1_LOC_816/a_36_24# INVX1_LOC_63/A 0.00fF
C59915 INVX1_LOC_161/Y INVX1_LOC_92/A 0.03fF
C59916 NOR2X1_LOC_68/A NOR2X1_LOC_816/Y 0.01fF
C59917 INVX1_LOC_14/A NAND2X1_LOC_574/A 0.16fF
C59918 INVX1_LOC_1/A NAND2X1_LOC_659/A 0.05fF
C59919 INVX1_LOC_27/A INVX1_LOC_186/Y 0.00fF
C59920 NOR2X1_LOC_242/A INVX1_LOC_19/A 4.34fF
C59921 NAND2X1_LOC_702/a_36_24# INVX1_LOC_109/A 0.00fF
C59922 NOR2X1_LOC_672/Y NOR2X1_LOC_825/Y 0.20fF
C59923 D_INPUT_0 NOR2X1_LOC_750/A 0.32fF
C59924 INVX1_LOC_58/A INVX1_LOC_231/A 0.03fF
C59925 INVX1_LOC_64/A NAND2X1_LOC_792/B 0.28fF
C59926 NOR2X1_LOC_344/A NOR2X1_LOC_35/Y 0.52fF
C59927 NOR2X1_LOC_712/B VDD 0.02fF
C59928 NAND2X1_LOC_175/B NOR2X1_LOC_173/a_36_216# 0.00fF
C59929 NOR2X1_LOC_773/Y INVX1_LOC_100/Y 0.01fF
C59930 NOR2X1_LOC_82/A NAND2X1_LOC_572/B 0.01fF
C59931 INVX1_LOC_39/A INVX1_LOC_29/A 0.07fF
C59932 INVX1_LOC_24/A INVX1_LOC_44/A 0.07fF
C59933 NAND2X1_LOC_634/Y INVX1_LOC_118/A 0.14fF
C59934 INVX1_LOC_305/A NOR2X1_LOC_729/A 0.26fF
C59935 NOR2X1_LOC_570/B NOR2X1_LOC_562/A 0.07fF
C59936 NAND2X1_LOC_374/Y NAND2X1_LOC_623/B 0.13fF
C59937 GATE_811 INVX1_LOC_20/A 0.00fF
C59938 NOR2X1_LOC_716/B NAND2X1_LOC_721/A 0.07fF
C59939 NAND2X1_LOC_125/a_36_24# INVX1_LOC_75/A 0.01fF
C59940 INVX1_LOC_98/Y INVX1_LOC_93/Y 0.02fF
C59941 INVX1_LOC_160/Y NOR2X1_LOC_835/B 0.28fF
C59942 VDD INVX1_LOC_103/Y -0.00fF
C59943 INVX1_LOC_290/Y NOR2X1_LOC_644/a_36_216# 0.01fF
C59944 INVX1_LOC_90/A NOR2X1_LOC_302/Y 0.01fF
C59945 NAND2X1_LOC_811/Y INVX1_LOC_46/A 0.06fF
C59946 VDD INVX1_LOC_315/A 0.00fF
C59947 NAND2X1_LOC_563/a_36_24# NOR2X1_LOC_649/B -0.02fF
C59948 NAND2X1_LOC_364/A NOR2X1_LOC_612/Y 0.00fF
C59949 NAND2X1_LOC_850/Y NAND2X1_LOC_642/Y 0.01fF
C59950 NOR2X1_LOC_710/B NAND2X1_LOC_782/B 0.04fF
C59951 INVX1_LOC_176/A NOR2X1_LOC_87/B 0.03fF
C59952 NAND2X1_LOC_276/Y INVX1_LOC_117/A 0.43fF
C59953 INVX1_LOC_24/A NOR2X1_LOC_641/Y 0.04fF
C59954 INVX1_LOC_120/A NOR2X1_LOC_188/A 0.03fF
C59955 INVX1_LOC_13/Y INVX1_LOC_15/A 0.07fF
C59956 NAND2X1_LOC_190/Y INVX1_LOC_263/Y 0.03fF
C59957 INVX1_LOC_266/Y INVX1_LOC_46/A 0.02fF
C59958 INVX1_LOC_135/A NOR2X1_LOC_391/Y 0.03fF
C59959 INVX1_LOC_49/A INVX1_LOC_118/Y 0.04fF
C59960 INVX1_LOC_33/A NOR2X1_LOC_114/a_36_216# 0.01fF
C59961 GATE_811 NOR2X1_LOC_765/Y 0.00fF
C59962 NAND2X1_LOC_811/Y NOR2X1_LOC_766/Y 0.03fF
C59963 NOR2X1_LOC_318/B NOR2X1_LOC_501/a_36_216# 0.00fF
C59964 INVX1_LOC_149/A VDD 0.00fF
C59965 NOR2X1_LOC_468/Y INVX1_LOC_42/A 0.01fF
C59966 INVX1_LOC_77/A INVX1_LOC_274/A 0.07fF
C59967 NAND2X1_LOC_842/B INPUT_0 0.03fF
C59968 NOR2X1_LOC_214/B INVX1_LOC_6/A 0.04fF
C59969 NAND2X1_LOC_190/Y INVX1_LOC_42/A 0.07fF
C59970 INVX1_LOC_233/A INVX1_LOC_183/A 0.04fF
C59971 NOR2X1_LOC_414/Y NAND2X1_LOC_215/A 0.25fF
C59972 NOR2X1_LOC_437/Y INVX1_LOC_92/A 0.02fF
C59973 NOR2X1_LOC_433/A NOR2X1_LOC_433/Y 0.21fF
C59974 NOR2X1_LOC_106/Y NOR2X1_LOC_155/A 0.42fF
C59975 INVX1_LOC_8/A INVX1_LOC_118/A 0.15fF
C59976 INVX1_LOC_286/A INVX1_LOC_87/Y 0.23fF
C59977 INVX1_LOC_35/A NOR2X1_LOC_113/a_36_216# 0.00fF
C59978 NOR2X1_LOC_433/A NAND2X1_LOC_798/B 0.07fF
C59979 NOR2X1_LOC_808/A NOR2X1_LOC_319/B 0.03fF
C59980 INVX1_LOC_50/Y NOR2X1_LOC_621/B 0.06fF
C59981 INVX1_LOC_88/A INVX1_LOC_15/A 0.03fF
C59982 NOR2X1_LOC_123/B NOR2X1_LOC_124/A 0.03fF
C59983 INVX1_LOC_2/A INVX1_LOC_118/Y 0.05fF
C59984 NAND2X1_LOC_208/B INVX1_LOC_284/A 0.01fF
C59985 NOR2X1_LOC_147/B INVX1_LOC_307/A 0.22fF
C59986 NAND2X1_LOC_394/a_36_24# INVX1_LOC_166/A 0.00fF
C59987 INVX1_LOC_232/Y INVX1_LOC_280/A 0.01fF
C59988 INVX1_LOC_13/A INVX1_LOC_37/A 0.00fF
C59989 INVX1_LOC_34/A NAND2X1_LOC_243/B 0.22fF
C59990 NOR2X1_LOC_242/A INVX1_LOC_26/Y 0.03fF
C59991 NAND2X1_LOC_690/a_36_24# NOR2X1_LOC_729/A 0.00fF
C59992 NOR2X1_LOC_468/Y INVX1_LOC_78/A 0.08fF
C59993 INVX1_LOC_164/A VDD 0.15fF
C59994 INVX1_LOC_27/A NOR2X1_LOC_843/B 0.03fF
C59995 NAND2X1_LOC_190/Y INVX1_LOC_78/A 0.03fF
C59996 NAND2X1_LOC_79/a_36_24# INVX1_LOC_84/A 0.00fF
C59997 INVX1_LOC_21/A NOR2X1_LOC_727/B 0.03fF
C59998 INVX1_LOC_232/A NOR2X1_LOC_536/A 0.03fF
C59999 NOR2X1_LOC_52/B NAND2X1_LOC_798/B 0.07fF
C60000 NOR2X1_LOC_500/Y INVX1_LOC_38/A 0.07fF
C60001 INVX1_LOC_31/A NOR2X1_LOC_554/A 0.01fF
C60002 NOR2X1_LOC_121/Y INVX1_LOC_123/Y 0.20fF
C60003 NOR2X1_LOC_209/a_36_216# INVX1_LOC_117/A 0.00fF
C60004 INVX1_LOC_143/A NOR2X1_LOC_641/Y 0.01fF
C60005 INVX1_LOC_35/A INVX1_LOC_292/Y 0.07fF
C60006 INVX1_LOC_226/Y INVX1_LOC_38/A 0.07fF
C60007 NOR2X1_LOC_391/B NOR2X1_LOC_391/Y 0.01fF
C60008 INVX1_LOC_61/A INVX1_LOC_29/A 0.04fF
C60009 NOR2X1_LOC_672/Y INVX1_LOC_84/A 0.00fF
C60010 INVX1_LOC_249/A INVX1_LOC_186/Y 0.10fF
C60011 INVX1_LOC_313/Y NOR2X1_LOC_137/a_36_216# 0.02fF
C60012 NOR2X1_LOC_68/A INVX1_LOC_106/Y 0.00fF
C60013 NOR2X1_LOC_567/B INVX1_LOC_65/A 0.10fF
C60014 NAND2X1_LOC_729/B NAND2X1_LOC_863/A 0.32fF
C60015 NOR2X1_LOC_361/B INVX1_LOC_26/A 0.13fF
C60016 NOR2X1_LOC_590/A INVX1_LOC_21/Y 0.03fF
C60017 NAND2X1_LOC_361/Y NOR2X1_LOC_691/B 0.12fF
C60018 NOR2X1_LOC_174/B INVX1_LOC_37/A 0.00fF
C60019 NOR2X1_LOC_741/A INVX1_LOC_6/A 0.01fF
C60020 INVX1_LOC_269/A INVX1_LOC_28/Y 0.03fF
C60021 INVX1_LOC_278/A INVX1_LOC_13/Y 0.00fF
C60022 INVX1_LOC_24/Y NOR2X1_LOC_383/B 0.03fF
C60023 NAND2X1_LOC_778/Y NAND2X1_LOC_793/B 0.10fF
C60024 NOR2X1_LOC_500/B INVX1_LOC_15/A 0.10fF
C60025 NAND2X1_LOC_850/A INVX1_LOC_76/A 0.30fF
C60026 INVX1_LOC_313/A INVX1_LOC_12/Y 0.07fF
C60027 INVX1_LOC_62/Y INVX1_LOC_42/A 0.01fF
C60028 INVX1_LOC_21/A NOR2X1_LOC_717/A 0.36fF
C60029 NOR2X1_LOC_689/Y NAND2X1_LOC_303/Y 0.03fF
C60030 INVX1_LOC_224/Y NOR2X1_LOC_15/Y 0.03fF
C60031 INVX1_LOC_10/A INVX1_LOC_38/A 0.21fF
C60032 INVX1_LOC_269/A INVX1_LOC_270/A 0.87fF
C60033 NOR2X1_LOC_389/A INVX1_LOC_78/A 0.04fF
C60034 INVX1_LOC_55/Y INVX1_LOC_37/A 0.04fF
C60035 NAND2X1_LOC_357/A NAND2X1_LOC_286/B 0.07fF
C60036 NAND2X1_LOC_523/a_36_24# NOR2X1_LOC_536/A 0.00fF
C60037 NOR2X1_LOC_596/A INVX1_LOC_42/A 0.14fF
C60038 INVX1_LOC_232/A NAND2X1_LOC_93/B 0.01fF
C60039 NOR2X1_LOC_15/Y NOR2X1_LOC_458/a_36_216# 0.00fF
C60040 NOR2X1_LOC_793/A INVX1_LOC_23/A 0.60fF
C60041 INPUT_0 NOR2X1_LOC_545/B 0.00fF
C60042 INVX1_LOC_70/Y INVX1_LOC_286/A 0.03fF
C60043 NOR2X1_LOC_91/A NAND2X1_LOC_550/A 0.03fF
C60044 D_INPUT_1 INVX1_LOC_101/Y 0.03fF
C60045 NOR2X1_LOC_313/Y NOR2X1_LOC_56/Y 0.01fF
C60046 NOR2X1_LOC_761/Y NOR2X1_LOC_409/B 0.06fF
C60047 NOR2X1_LOC_172/Y INVX1_LOC_12/A 0.02fF
C60048 INVX1_LOC_25/Y INVX1_LOC_35/Y 0.07fF
C60049 NOR2X1_LOC_554/B NOR2X1_LOC_38/B -0.01fF
C60050 INVX1_LOC_8/A NAND2X1_LOC_63/Y 0.03fF
C60051 NOR2X1_LOC_624/A INVX1_LOC_29/A 0.03fF
C60052 NOR2X1_LOC_255/Y NOR2X1_LOC_361/B 0.21fF
C60053 INVX1_LOC_45/A INVX1_LOC_273/A 0.03fF
C60054 NOR2X1_LOC_401/A INVX1_LOC_23/A 0.01fF
C60055 INVX1_LOC_22/A NOR2X1_LOC_216/B 0.10fF
C60056 INVX1_LOC_17/A INVX1_LOC_29/Y 0.03fF
C60057 NOR2X1_LOC_15/Y NAND2X1_LOC_793/B 0.01fF
C60058 NAND2X1_LOC_588/B NAND2X1_LOC_3/B 0.21fF
C60059 NOR2X1_LOC_798/A NOR2X1_LOC_220/B 0.01fF
C60060 NAND2X1_LOC_338/B NAND2X1_LOC_456/Y 0.01fF
C60061 NOR2X1_LOC_383/Y NAND2X1_LOC_93/B 0.55fF
C60062 NOR2X1_LOC_203/Y INVX1_LOC_84/A 0.01fF
C60063 NOR2X1_LOC_792/B NAND2X1_LOC_81/B 0.00fF
C60064 NOR2X1_LOC_65/B NOR2X1_LOC_389/A 0.10fF
C60065 INVX1_LOC_34/A INVX1_LOC_284/A 0.23fF
C60066 NOR2X1_LOC_606/Y INVX1_LOC_23/Y 0.04fF
C60067 NOR2X1_LOC_590/A NOR2X1_LOC_39/Y 0.01fF
C60068 NOR2X1_LOC_360/Y INVX1_LOC_4/Y 0.24fF
C60069 NOR2X1_LOC_392/B INVX1_LOC_12/A 3.34fF
C60070 INVX1_LOC_234/A NOR2X1_LOC_88/A 0.03fF
C60071 NOR2X1_LOC_561/Y NOR2X1_LOC_510/B 0.03fF
C60072 NOR2X1_LOC_81/a_36_216# INVX1_LOC_4/A 0.02fF
C60073 NAND2X1_LOC_725/A NAND2X1_LOC_303/Y 0.10fF
C60074 INVX1_LOC_5/A INVX1_LOC_52/Y 0.04fF
C60075 VDD NOR2X1_LOC_313/Y 0.12fF
C60076 INVX1_LOC_303/A INVX1_LOC_15/A 0.11fF
C60077 NOR2X1_LOC_278/a_36_216# INVX1_LOC_70/A 0.00fF
C60078 NOR2X1_LOC_634/B INVX1_LOC_19/A 0.59fF
C60079 NOR2X1_LOC_496/Y INVX1_LOC_178/A 0.02fF
C60080 NAND2X1_LOC_35/Y INVX1_LOC_14/A 0.07fF
C60081 INVX1_LOC_161/Y INVX1_LOC_53/A 1.49fF
C60082 NOR2X1_LOC_160/B INVX1_LOC_23/A 1.64fF
C60083 INVX1_LOC_232/A INVX1_LOC_3/A 0.10fF
C60084 NOR2X1_LOC_246/A NOR2X1_LOC_743/Y 0.18fF
C60085 NOR2X1_LOC_636/A NOR2X1_LOC_467/A 0.01fF
C60086 NOR2X1_LOC_78/B INVX1_LOC_19/A 7.92fF
C60087 INVX1_LOC_62/Y INVX1_LOC_78/A 0.02fF
C60088 INVX1_LOC_201/A D_INPUT_3 0.01fF
C60089 NOR2X1_LOC_596/A INVX1_LOC_78/A 0.09fF
C60090 NOR2X1_LOC_147/B NAND2X1_LOC_253/a_36_24# 0.01fF
C60091 NOR2X1_LOC_553/a_36_216# INVX1_LOC_53/A 0.01fF
C60092 INVX1_LOC_97/A INVX1_LOC_307/A 0.12fF
C60093 INVX1_LOC_11/A NAND2X1_LOC_31/a_36_24# 0.00fF
C60094 NAND2X1_LOC_59/B INVX1_LOC_15/A 0.00fF
C60095 NAND2X1_LOC_338/B NAND2X1_LOC_80/a_36_24# 0.00fF
C60096 INVX1_LOC_6/A INVX1_LOC_12/Y 0.64fF
C60097 INVX1_LOC_90/A INVX1_LOC_307/A 0.07fF
C60098 NAND2X1_LOC_342/Y NAND2X1_LOC_807/B 0.05fF
C60099 NOR2X1_LOC_848/Y INVX1_LOC_50/Y 0.03fF
C60100 INVX1_LOC_43/A NAND2X1_LOC_74/B 0.01fF
C60101 INVX1_LOC_125/Y INVX1_LOC_46/A 0.00fF
C60102 NOR2X1_LOC_68/A NOR2X1_LOC_635/B 0.21fF
C60103 NAND2X1_LOC_357/a_36_24# NAND2X1_LOC_288/B 0.00fF
C60104 INVX1_LOC_90/A NOR2X1_LOC_445/B 0.07fF
C60105 NOR2X1_LOC_68/A INVX1_LOC_275/Y 0.05fF
C60106 NAND2X1_LOC_757/a_36_24# NAND2X1_LOC_99/A 0.00fF
C60107 NOR2X1_LOC_68/A NOR2X1_LOC_748/A 0.07fF
C60108 INVX1_LOC_18/A INVX1_LOC_271/A 0.03fF
C60109 NOR2X1_LOC_716/B INVX1_LOC_87/A 0.08fF
C60110 NOR2X1_LOC_19/Y NOR2X1_LOC_629/Y 0.00fF
C60111 INVX1_LOC_18/A INVX1_LOC_105/Y 0.04fF
C60112 NAND2X1_LOC_18/a_36_24# INVX1_LOC_174/A 0.01fF
C60113 NOR2X1_LOC_391/Y INVX1_LOC_280/A 0.02fF
C60114 NAND2X1_LOC_392/Y INVX1_LOC_19/A 0.03fF
C60115 NOR2X1_LOC_552/A NOR2X1_LOC_168/a_36_216# 0.01fF
C60116 INVX1_LOC_136/A INVX1_LOC_308/A 0.03fF
C60117 NAND2X1_LOC_67/Y NOR2X1_LOC_666/Y 0.02fF
C60118 NOR2X1_LOC_631/B NOR2X1_LOC_357/Y 0.01fF
C60119 INVX1_LOC_136/A NAND2X1_LOC_827/a_36_24# -0.01fF
C60120 INVX1_LOC_75/A NAND2X1_LOC_656/B 0.04fF
C60121 NAND2X1_LOC_374/Y INVX1_LOC_3/Y 0.00fF
C60122 INVX1_LOC_58/A INVX1_LOC_244/Y 0.02fF
C60123 INVX1_LOC_50/A NOR2X1_LOC_484/Y 0.01fF
C60124 NAND2X1_LOC_9/Y INVX1_LOC_72/Y 0.03fF
C60125 NOR2X1_LOC_516/B NOR2X1_LOC_847/a_36_216# 0.00fF
C60126 INVX1_LOC_83/A INVX1_LOC_19/A 0.11fF
C60127 NOR2X1_LOC_9/Y NAND2X1_LOC_62/a_36_24# 0.00fF
C60128 INVX1_LOC_89/A NAND2X1_LOC_782/B 0.01fF
C60129 INVX1_LOC_96/A NOR2X1_LOC_331/B 0.52fF
C60130 NOR2X1_LOC_15/Y NOR2X1_LOC_103/Y 0.09fF
C60131 INVX1_LOC_244/A INVX1_LOC_84/A 0.09fF
C60132 NAND2X1_LOC_602/a_36_24# NAND2X1_LOC_472/Y 0.00fF
C60133 INVX1_LOC_41/A NOR2X1_LOC_383/B 0.80fF
C60134 INVX1_LOC_132/A INVX1_LOC_129/A 0.01fF
C60135 NOR2X1_LOC_295/Y NOR2X1_LOC_65/B 0.02fF
C60136 NAND2X1_LOC_391/Y INVX1_LOC_30/A 0.07fF
C60137 INVX1_LOC_64/A NOR2X1_LOC_359/Y -0.02fF
C60138 NOR2X1_LOC_455/a_36_216# NOR2X1_LOC_383/B 0.00fF
C60139 NAND2X1_LOC_447/Y NOR2X1_LOC_536/A 0.05fF
C60140 INVX1_LOC_206/Y INVX1_LOC_179/A 0.00fF
C60141 NOR2X1_LOC_52/B NAND2X1_LOC_211/a_36_24# 0.00fF
C60142 D_INPUT_0 INVX1_LOC_102/A 0.07fF
C60143 INVX1_LOC_58/A NAND2X1_LOC_276/Y 0.03fF
C60144 INVX1_LOC_93/Y NOR2X1_LOC_709/B 0.01fF
C60145 NOR2X1_LOC_797/a_36_216# INVX1_LOC_301/A 0.00fF
C60146 NOR2X1_LOC_220/A INVX1_LOC_78/A 0.08fF
C60147 INVX1_LOC_90/A INVX1_LOC_12/A 0.53fF
C60148 INPUT_0 INVX1_LOC_119/Y 0.02fF
C60149 NOR2X1_LOC_784/Y NOR2X1_LOC_803/B 0.00fF
C60150 INVX1_LOC_27/A INVX1_LOC_18/A 0.35fF
C60151 NOR2X1_LOC_405/A NOR2X1_LOC_612/Y 0.00fF
C60152 NOR2X1_LOC_262/Y NOR2X1_LOC_772/B 0.02fF
C60153 INVX1_LOC_90/A NOR2X1_LOC_519/Y 0.01fF
C60154 NOR2X1_LOC_824/A INVX1_LOC_18/A 0.07fF
C60155 INVX1_LOC_313/Y INVX1_LOC_99/A 0.08fF
C60156 INVX1_LOC_226/Y NAND2X1_LOC_223/A 0.07fF
C60157 INVX1_LOC_35/A NAND2X1_LOC_361/Y 0.07fF
C60158 NOR2X1_LOC_389/B INVX1_LOC_12/A 0.07fF
C60159 INVX1_LOC_45/A NOR2X1_LOC_15/Y 0.06fF
C60160 NAND2X1_LOC_53/Y NOR2X1_LOC_483/B 0.01fF
C60161 INVX1_LOC_163/A INVX1_LOC_195/A 0.01fF
C60162 INVX1_LOC_50/A NOR2X1_LOC_423/Y 0.04fF
C60163 NOR2X1_LOC_685/A NAND2X1_LOC_425/Y 0.03fF
C60164 NOR2X1_LOC_231/B INVX1_LOC_11/A 0.02fF
C60165 INVX1_LOC_39/A NOR2X1_LOC_256/a_36_216# 0.00fF
C60166 INVX1_LOC_233/Y INVX1_LOC_207/A 0.12fF
C60167 INVX1_LOC_286/A INVX1_LOC_285/A 0.22fF
C60168 NOR2X1_LOC_15/Y NAND2X1_LOC_856/A 0.59fF
C60169 NOR2X1_LOC_112/Y NAND2X1_LOC_291/B 0.40fF
C60170 INVX1_LOC_36/A INVX1_LOC_269/A 0.03fF
C60171 INVX1_LOC_243/Y INVX1_LOC_243/A 0.14fF
C60172 INVX1_LOC_209/Y NOR2X1_LOC_304/a_36_216# 0.00fF
C60173 INVX1_LOC_136/A NAND2X1_LOC_579/A 0.08fF
C60174 NAND2X1_LOC_550/A INVX1_LOC_31/A 0.07fF
C60175 NOR2X1_LOC_690/A NAND2X1_LOC_725/A 0.10fF
C60176 NOR2X1_LOC_167/Y NOR2X1_LOC_662/A 0.02fF
C60177 NOR2X1_LOC_143/a_36_216# NOR2X1_LOC_392/Y 0.00fF
C60178 NOR2X1_LOC_142/Y NOR2X1_LOC_665/Y 0.01fF
C60179 NOR2X1_LOC_91/A NAND2X1_LOC_853/Y 0.01fF
C60180 INVX1_LOC_286/A NOR2X1_LOC_814/A 0.10fF
C60181 NOR2X1_LOC_160/B INVX1_LOC_31/A 0.17fF
C60182 NAND2X1_LOC_1/a_36_24# INVX1_LOC_15/A 0.00fF
C60183 INVX1_LOC_50/A NOR2X1_LOC_222/Y 0.07fF
C60184 INVX1_LOC_5/A INVX1_LOC_63/Y 0.10fF
C60185 INVX1_LOC_58/A NAND2X1_LOC_374/Y 0.07fF
C60186 NAND2X1_LOC_348/A INVX1_LOC_12/A 0.03fF
C60187 NOR2X1_LOC_781/B NOR2X1_LOC_158/Y 0.01fF
C60188 INVX1_LOC_225/A NOR2X1_LOC_211/Y 0.02fF
C60189 INVX1_LOC_278/A INVX1_LOC_168/A 0.00fF
C60190 INVX1_LOC_75/A NOR2X1_LOC_610/Y 0.01fF
C60191 NOR2X1_LOC_824/A INVX1_LOC_172/A 0.07fF
C60192 INVX1_LOC_34/A NOR2X1_LOC_674/Y 0.07fF
C60193 INVX1_LOC_91/A NAND2X1_LOC_475/Y 0.10fF
C60194 INVX1_LOC_73/Y INVX1_LOC_130/Y 0.00fF
C60195 INVX1_LOC_13/Y NAND2X1_LOC_464/Y 0.05fF
C60196 NOR2X1_LOC_186/Y NOR2X1_LOC_758/Y 0.01fF
C60197 NOR2X1_LOC_15/Y INVX1_LOC_71/A 0.12fF
C60198 INVX1_LOC_33/A NAND2X1_LOC_474/Y 0.07fF
C60199 INVX1_LOC_21/A NAND2X1_LOC_175/B 0.07fF
C60200 NOR2X1_LOC_2/Y NOR2X1_LOC_12/a_36_216# 0.00fF
C60201 NAND2X1_LOC_573/A INVX1_LOC_26/A 0.02fF
C60202 NOR2X1_LOC_451/A INVX1_LOC_37/A 0.01fF
C60203 INVX1_LOC_95/A INVX1_LOC_285/A 0.06fF
C60204 INPUT_0 INVX1_LOC_284/A 0.07fF
C60205 INVX1_LOC_208/A INVX1_LOC_23/A 0.09fF
C60206 VDD NOR2X1_LOC_235/Y 0.12fF
C60207 INVX1_LOC_39/A INVX1_LOC_8/A 0.06fF
C60208 NOR2X1_LOC_92/Y NAND2X1_LOC_632/B 0.02fF
C60209 INVX1_LOC_293/A NOR2X1_LOC_791/B 0.30fF
C60210 INVX1_LOC_161/A INVX1_LOC_72/A 0.23fF
C60211 NOR2X1_LOC_74/A INVX1_LOC_290/Y 0.07fF
C60212 NOR2X1_LOC_516/B INVX1_LOC_23/A 0.05fF
C60213 INVX1_LOC_21/A NAND2X1_LOC_142/a_36_24# 0.00fF
C60214 NOR2X1_LOC_180/B NOR2X1_LOC_334/Y 0.07fF
C60215 INVX1_LOC_5/A NOR2X1_LOC_175/A 0.07fF
C60216 INVX1_LOC_235/A NOR2X1_LOC_516/Y 0.06fF
C60217 INVX1_LOC_74/Y INVX1_LOC_3/A 0.03fF
C60218 INVX1_LOC_25/Y NOR2X1_LOC_15/a_36_216# 0.00fF
C60219 NAND2X1_LOC_794/B NAND2X1_LOC_357/B 0.07fF
C60220 NAND2X1_LOC_860/A INVX1_LOC_25/Y 0.18fF
C60221 INVX1_LOC_83/A INVX1_LOC_26/Y 0.03fF
C60222 NAND2X1_LOC_573/Y NOR2X1_LOC_758/Y 0.02fF
C60223 NOR2X1_LOC_7/Y INVX1_LOC_29/A 0.03fF
C60224 INVX1_LOC_172/Y NOR2X1_LOC_392/Y 0.29fF
C60225 NAND2X1_LOC_288/A INVX1_LOC_46/A 0.13fF
C60226 VDD INVX1_LOC_260/Y 0.21fF
C60227 NOR2X1_LOC_561/Y INVX1_LOC_57/A 0.23fF
C60228 NOR2X1_LOC_459/B INVX1_LOC_239/A 0.03fF
C60229 INVX1_LOC_166/A NOR2X1_LOC_459/A 0.53fF
C60230 INVX1_LOC_202/A NOR2X1_LOC_218/A 0.05fF
C60231 INVX1_LOC_266/A NOR2X1_LOC_388/Y 0.12fF
C60232 INVX1_LOC_174/A NOR2X1_LOC_546/B 0.05fF
C60233 NAND2X1_LOC_549/Y INVX1_LOC_16/A 0.05fF
C60234 NAND2X1_LOC_785/B INVX1_LOC_217/A 0.02fF
C60235 D_INPUT_0 NAND2X1_LOC_439/a_36_24# 0.01fF
C60236 NOR2X1_LOC_703/B INVX1_LOC_30/A 0.03fF
C60237 NOR2X1_LOC_78/A INVX1_LOC_69/A 0.07fF
C60238 INVX1_LOC_73/A NOR2X1_LOC_334/Y 0.12fF
C60239 NAND2X1_LOC_423/a_36_24# INVX1_LOC_117/Y 0.00fF
C60240 NOR2X1_LOC_679/Y NOR2X1_LOC_433/A 0.03fF
C60241 NOR2X1_LOC_82/A NOR2X1_LOC_716/B 0.10fF
C60242 NOR2X1_LOC_368/Y INVX1_LOC_19/A 0.01fF
C60243 NAND2X1_LOC_53/Y INVX1_LOC_33/A 0.03fF
C60244 NAND2X1_LOC_738/B NOR2X1_LOC_299/Y 0.01fF
C60245 NAND2X1_LOC_732/a_36_24# NOR2X1_LOC_298/Y 0.09fF
C60246 NOR2X1_LOC_653/Y INVX1_LOC_46/A 0.01fF
C60247 INVX1_LOC_14/A NAND2X1_LOC_465/Y 0.03fF
C60248 INVX1_LOC_38/A INVX1_LOC_307/A 0.07fF
C60249 INVX1_LOC_44/A NOR2X1_LOC_197/B 0.25fF
C60250 INVX1_LOC_21/A INVX1_LOC_256/Y 0.07fF
C60251 INVX1_LOC_269/A NOR2X1_LOC_309/Y 0.01fF
C60252 NOR2X1_LOC_222/Y NOR2X1_LOC_206/a_36_216# 0.00fF
C60253 NAND2X1_LOC_725/A NOR2X1_LOC_32/a_36_216# 0.16fF
C60254 INVX1_LOC_299/A NOR2X1_LOC_802/A 0.03fF
C60255 INVX1_LOC_38/A NOR2X1_LOC_445/B 0.07fF
C60256 INVX1_LOC_37/A NAND2X1_LOC_489/Y 0.02fF
C60257 NOR2X1_LOC_389/A INVX1_LOC_113/Y 0.03fF
C60258 INVX1_LOC_16/A NOR2X1_LOC_291/Y 0.17fF
C60259 NAND2X1_LOC_244/a_36_24# INVX1_LOC_118/A 0.00fF
C60260 INVX1_LOC_46/A INVX1_LOC_19/A 0.45fF
C60261 NOR2X1_LOC_692/Y NOR2X1_LOC_485/a_36_216# 0.03fF
C60262 INVX1_LOC_50/A NOR2X1_LOC_329/B 0.85fF
C60263 INVX1_LOC_227/Y INVX1_LOC_94/A 0.01fF
C60264 NOR2X1_LOC_793/Y INVX1_LOC_196/A 0.40fF
C60265 NOR2X1_LOC_690/A NOR2X1_LOC_372/A 0.02fF
C60266 NOR2X1_LOC_303/Y NOR2X1_LOC_274/B 0.10fF
C60267 INVX1_LOC_46/A NOR2X1_LOC_11/Y 0.00fF
C60268 INVX1_LOC_245/Y INVX1_LOC_85/A 0.00fF
C60269 D_INPUT_3 INVX1_LOC_29/A 0.14fF
C60270 INVX1_LOC_249/A INVX1_LOC_18/A 0.16fF
C60271 INVX1_LOC_75/A NOR2X1_LOC_35/a_36_216# 0.00fF
C60272 INVX1_LOC_14/Y INVX1_LOC_29/A 0.02fF
C60273 INVX1_LOC_6/A NOR2X1_LOC_89/Y 0.27fF
C60274 NOR2X1_LOC_636/a_36_216# INVX1_LOC_30/A 0.01fF
C60275 NAND2X1_LOC_213/A NOR2X1_LOC_210/B 0.04fF
C60276 NOR2X1_LOC_468/Y NAND2X1_LOC_860/Y 0.06fF
C60277 NOR2X1_LOC_193/a_36_216# INVX1_LOC_26/Y 0.00fF
C60278 NAND2X1_LOC_550/A NOR2X1_LOC_290/Y 0.11fF
C60279 NAND2X1_LOC_347/B INVX1_LOC_16/A 0.07fF
C60280 NOR2X1_LOC_430/A NOR2X1_LOC_582/Y 0.38fF
C60281 INVX1_LOC_272/Y NAND2X1_LOC_798/A 0.02fF
C60282 INVX1_LOC_54/A INVX1_LOC_285/A 0.08fF
C60283 INVX1_LOC_1/A INVX1_LOC_56/Y 0.01fF
C60284 INVX1_LOC_2/Y NOR2X1_LOC_346/A 0.01fF
C60285 INVX1_LOC_27/A NOR2X1_LOC_383/a_36_216# 0.00fF
C60286 INVX1_LOC_135/A INVX1_LOC_50/Y 0.03fF
C60287 NOR2X1_LOC_817/Y NAND2X1_LOC_819/Y 0.01fF
C60288 NOR2X1_LOC_78/B INVX1_LOC_161/Y 0.09fF
C60289 NAND2X1_LOC_243/B NAND2X1_LOC_240/a_36_24# 0.02fF
C60290 INVX1_LOC_311/A NOR2X1_LOC_727/B 0.26fF
C60291 INVX1_LOC_34/A INVX1_LOC_72/A 13.40fF
C60292 NAND2X1_LOC_175/B NAND2X1_LOC_354/Y 0.00fF
C60293 INVX1_LOC_54/A NOR2X1_LOC_814/A 0.10fF
C60294 INVX1_LOC_284/Y NAND2X1_LOC_839/Y 0.04fF
C60295 INVX1_LOC_304/Y NAND2X1_LOC_785/B 0.02fF
C60296 NAND2X1_LOC_860/A INVX1_LOC_75/A 0.03fF
C60297 INVX1_LOC_33/Y NOR2X1_LOC_89/A 0.00fF
C60298 NOR2X1_LOC_596/A INVX1_LOC_113/Y 0.04fF
C60299 INVX1_LOC_33/Y NAND2X1_LOC_668/a_36_24# 0.00fF
C60300 NAND2X1_LOC_632/B NAND2X1_LOC_837/Y 0.03fF
C60301 NOR2X1_LOC_262/Y INVX1_LOC_303/A 0.10fF
C60302 NOR2X1_LOC_167/Y INVX1_LOC_57/A 0.06fF
C60303 NOR2X1_LOC_560/A INVX1_LOC_50/Y 0.14fF
C60304 INVX1_LOC_61/A INVX1_LOC_8/A 0.09fF
C60305 NAND2X1_LOC_640/Y INVX1_LOC_41/Y 0.19fF
C60306 NOR2X1_LOC_720/A NAND2X1_LOC_669/a_36_24# 0.02fF
C60307 NOR2X1_LOC_530/a_36_216# INVX1_LOC_25/Y 0.00fF
C60308 NAND2X1_LOC_338/B NAND2X1_LOC_208/B 0.05fF
C60309 INVX1_LOC_201/Y NOR2X1_LOC_480/A 0.39fF
C60310 NOR2X1_LOC_759/a_36_216# INVX1_LOC_63/Y 0.00fF
C60311 NOR2X1_LOC_536/A NAND2X1_LOC_263/a_36_24# 0.00fF
C60312 INVX1_LOC_12/A INVX1_LOC_38/A 0.24fF
C60313 INVX1_LOC_17/A INVX1_LOC_101/A 0.01fF
C60314 INVX1_LOC_28/A NOR2X1_LOC_291/Y 0.20fF
C60315 INVX1_LOC_37/A INVX1_LOC_32/A 0.03fF
C60316 NAND2X1_LOC_848/A INVX1_LOC_102/A 0.10fF
C60317 INVX1_LOC_78/A NAND2X1_LOC_655/B 0.02fF
C60318 INVX1_LOC_54/Y NOR2X1_LOC_274/B 0.07fF
C60319 INVX1_LOC_78/A NAND2X1_LOC_469/B 0.03fF
C60320 NAND2X1_LOC_184/a_36_24# INVX1_LOC_50/Y 0.01fF
C60321 INVX1_LOC_37/A NOR2X1_LOC_623/B -0.00fF
C60322 NOR2X1_LOC_209/Y INVX1_LOC_142/A 0.04fF
C60323 NOR2X1_LOC_653/B NAND2X1_LOC_807/Y 0.02fF
C60324 NAND2X1_LOC_550/A NAND2X1_LOC_859/Y 0.15fF
C60325 NAND2X1_LOC_231/Y INVX1_LOC_72/A 0.02fF
C60326 INVX1_LOC_45/Y INVX1_LOC_104/A 0.11fF
C60327 NOR2X1_LOC_468/Y NAND2X1_LOC_861/Y 0.21fF
C60328 INVX1_LOC_37/A NOR2X1_LOC_329/Y 0.27fF
C60329 NOR2X1_LOC_516/B INVX1_LOC_31/A 0.29fF
C60330 NOR2X1_LOC_158/Y NOR2X1_LOC_585/Y 0.03fF
C60331 NOR2X1_LOC_720/A NAND2X1_LOC_642/Y 0.01fF
C60332 INVX1_LOC_45/A NAND2X1_LOC_840/B 0.03fF
C60333 NOR2X1_LOC_78/A INVX1_LOC_270/Y 0.26fF
C60334 VDD NAND2X1_LOC_471/Y 0.04fF
C60335 INVX1_LOC_17/A NOR2X1_LOC_355/A 0.08fF
C60336 NOR2X1_LOC_606/Y INVX1_LOC_232/A 0.01fF
C60337 NOR2X1_LOC_51/A INVX1_LOC_12/A 0.46fF
C60338 NOR2X1_LOC_52/a_36_216# NAND2X1_LOC_454/Y 0.01fF
C60339 NOR2X1_LOC_303/Y NOR2X1_LOC_348/B 0.25fF
C60340 NAND2X1_LOC_21/Y NAND2X1_LOC_59/B 0.10fF
C60341 INVX1_LOC_134/A NOR2X1_LOC_326/Y 0.14fF
C60342 NOR2X1_LOC_721/A INVX1_LOC_62/Y 0.05fF
C60343 NAND2X1_LOC_812/A NAND2X1_LOC_811/Y 0.00fF
C60344 INVX1_LOC_83/A INVX1_LOC_161/Y 0.10fF
C60345 NOR2X1_LOC_447/B INVX1_LOC_78/A 0.04fF
C60346 INVX1_LOC_290/A INVX1_LOC_81/Y 0.02fF
C60347 INVX1_LOC_27/A INVX1_LOC_31/Y 0.04fF
C60348 NOR2X1_LOC_91/Y NAND2X1_LOC_850/Y 0.37fF
C60349 NOR2X1_LOC_681/Y NAND2X1_LOC_175/Y 0.51fF
C60350 INVX1_LOC_111/Y INVX1_LOC_94/A 0.05fF
C60351 NAND2X1_LOC_787/A INVX1_LOC_91/A 0.03fF
C60352 INVX1_LOC_96/Y INVX1_LOC_71/A 0.05fF
C60353 INVX1_LOC_37/A NAND2X1_LOC_175/Y 0.07fF
C60354 INVX1_LOC_26/A NAND2X1_LOC_267/B -0.00fF
C60355 NAND2X1_LOC_705/Y NAND2X1_LOC_560/A 0.01fF
C60356 NOR2X1_LOC_759/Y NOR2X1_LOC_131/A 0.01fF
C60357 INVX1_LOC_279/Y INVX1_LOC_279/A 0.03fF
C60358 INVX1_LOC_298/Y INVX1_LOC_14/Y 0.60fF
C60359 INVX1_LOC_181/Y NOR2X1_LOC_191/A 0.04fF
C60360 NAND2X1_LOC_363/B INVX1_LOC_91/A 0.46fF
C60361 INVX1_LOC_50/A NOR2X1_LOC_69/A 0.02fF
C60362 INVX1_LOC_200/A INVX1_LOC_90/A 0.11fF
C60363 NOR2X1_LOC_667/A NOR2X1_LOC_13/Y 0.00fF
C60364 NOR2X1_LOC_498/Y NAND2X1_LOC_706/a_36_24# 0.00fF
C60365 NAND2X1_LOC_472/Y NOR2X1_LOC_464/Y 0.04fF
C60366 INVX1_LOC_21/A NOR2X1_LOC_337/A 0.04fF
C60367 NOR2X1_LOC_15/Y INVX1_LOC_102/Y 0.03fF
C60368 INVX1_LOC_45/A NOR2X1_LOC_97/B 0.01fF
C60369 NOR2X1_LOC_740/Y INVX1_LOC_311/Y 0.00fF
C60370 NAND2X1_LOC_550/A NAND2X1_LOC_866/B 0.05fF
C60371 NAND2X1_LOC_341/A INVX1_LOC_159/A 0.02fF
C60372 NAND2X1_LOC_787/A INVX1_LOC_11/Y 0.03fF
C60373 NOR2X1_LOC_324/B INVX1_LOC_23/A 0.01fF
C60374 INVX1_LOC_49/A NOR2X1_LOC_520/A 0.10fF
C60375 INVX1_LOC_57/A INVX1_LOC_76/A 0.17fF
C60376 NOR2X1_LOC_84/A NOR2X1_LOC_84/a_36_216# 0.01fF
C60377 NAND2X1_LOC_43/a_36_24# NAND2X1_LOC_508/A 0.00fF
C60378 NOR2X1_LOC_478/A INVX1_LOC_89/A 0.01fF
C60379 INVX1_LOC_32/A NOR2X1_LOC_743/Y 0.01fF
C60380 INVX1_LOC_37/A INVX1_LOC_262/A 0.01fF
C60381 INVX1_LOC_269/A NOR2X1_LOC_19/Y 0.01fF
C60382 NOR2X1_LOC_500/A NOR2X1_LOC_325/A -0.02fF
C60383 NOR2X1_LOC_833/Y NOR2X1_LOC_678/A 0.02fF
C60384 NOR2X1_LOC_319/B NOR2X1_LOC_863/B 0.01fF
C60385 NAND2X1_LOC_807/B INVX1_LOC_285/A 0.36fF
C60386 NOR2X1_LOC_220/A INVX1_LOC_113/Y 0.04fF
C60387 NOR2X1_LOC_471/Y NOR2X1_LOC_736/Y 0.12fF
C60388 INVX1_LOC_90/A NAND2X1_LOC_733/Y 0.05fF
C60389 INVX1_LOC_23/A NAND2X1_LOC_211/Y 0.12fF
C60390 INVX1_LOC_234/A INVX1_LOC_18/A 0.00fF
C60391 NOR2X1_LOC_791/Y INVX1_LOC_91/A 0.01fF
C60392 INVX1_LOC_274/A INVX1_LOC_274/Y 0.01fF
C60393 NOR2X1_LOC_303/Y INVX1_LOC_22/A 0.02fF
C60394 INVX1_LOC_207/A NOR2X1_LOC_526/Y 0.01fF
C60395 INVX1_LOC_34/A NAND2X1_LOC_338/B 0.03fF
C60396 INVX1_LOC_12/Y INVX1_LOC_270/A 0.03fF
C60397 NOR2X1_LOC_666/A INVX1_LOC_285/Y 0.03fF
C60398 VDD NOR2X1_LOC_696/Y 0.02fF
C60399 NOR2X1_LOC_361/B NOR2X1_LOC_368/A 0.06fF
C60400 INVX1_LOC_36/A NOR2X1_LOC_814/Y 0.01fF
C60401 INVX1_LOC_183/Y INVX1_LOC_30/A 0.01fF
C60402 INVX1_LOC_14/A NOR2X1_LOC_83/Y 1.59fF
C60403 INVX1_LOC_37/A NOR2X1_LOC_622/A 0.15fF
C60404 NOR2X1_LOC_514/Y INVX1_LOC_216/A 0.01fF
C60405 NOR2X1_LOC_552/A INVX1_LOC_50/Y 0.07fF
C60406 NOR2X1_LOC_48/B INVX1_LOC_285/A 0.05fF
C60407 INVX1_LOC_276/A NOR2X1_LOC_574/A 0.13fF
C60408 INVX1_LOC_103/A NOR2X1_LOC_815/A 0.01fF
C60409 INVX1_LOC_33/A NOR2X1_LOC_500/Y 0.08fF
C60410 INVX1_LOC_226/Y INVX1_LOC_33/A 0.03fF
C60411 NOR2X1_LOC_718/a_36_216# INVX1_LOC_266/Y 0.00fF
C60412 INVX1_LOC_27/A NAND2X1_LOC_86/Y 0.02fF
C60413 INVX1_LOC_11/A NOR2X1_LOC_775/a_36_216# 0.00fF
C60414 NOR2X1_LOC_68/A INVX1_LOC_89/A 0.62fF
C60415 NOR2X1_LOC_246/A NAND2X1_LOC_198/B 0.10fF
C60416 NOR2X1_LOC_84/B INVX1_LOC_284/A -0.01fF
C60417 INVX1_LOC_279/A NAND2X1_LOC_140/a_36_24# 0.00fF
C60418 NAND2X1_LOC_175/Y NOR2X1_LOC_743/Y 0.18fF
C60419 INVX1_LOC_90/A INVX1_LOC_217/A 0.06fF
C60420 INVX1_LOC_286/Y NAND2X1_LOC_740/B 0.03fF
C60421 INVX1_LOC_172/A INVX1_LOC_234/A 0.01fF
C60422 NOR2X1_LOC_772/A INVX1_LOC_18/A 0.00fF
C60423 NAND2X1_LOC_550/A INVX1_LOC_6/A 0.02fF
C60424 NAND2X1_LOC_456/a_36_24# NAND2X1_LOC_773/B 0.00fF
C60425 INVX1_LOC_266/A NOR2X1_LOC_552/A 0.10fF
C60426 NOR2X1_LOC_68/A NAND2X1_LOC_508/A 0.03fF
C60427 INVX1_LOC_54/Y NOR2X1_LOC_175/B 0.13fF
C60428 NOR2X1_LOC_352/Y NOR2X1_LOC_357/a_36_216# 0.00fF
C60429 NOR2X1_LOC_632/Y NOR2X1_LOC_144/Y 0.01fF
C60430 INVX1_LOC_33/A INVX1_LOC_10/A 0.29fF
C60431 NOR2X1_LOC_160/B INVX1_LOC_6/A 0.15fF
C60432 INVX1_LOC_49/A NOR2X1_LOC_333/A 0.01fF
C60433 NOR2X1_LOC_457/A INVX1_LOC_91/A 0.03fF
C60434 NOR2X1_LOC_559/B NOR2X1_LOC_560/A 0.14fF
C60435 NOR2X1_LOC_653/Y NOR2X1_LOC_282/a_36_216# 0.00fF
C60436 INVX1_LOC_54/Y INVX1_LOC_22/A 0.15fF
C60437 NAND2X1_LOC_729/Y NOR2X1_LOC_385/Y 0.02fF
C60438 INVX1_LOC_10/A NAND2X1_LOC_466/A 0.01fF
C60439 INVX1_LOC_272/A INVX1_LOC_15/A 0.07fF
C60440 INVX1_LOC_49/A D_GATE_366 0.07fF
C60441 INVX1_LOC_72/A INPUT_0 0.12fF
C60442 INVX1_LOC_77/A NOR2X1_LOC_356/A 0.09fF
C60443 INVX1_LOC_20/A NAND2X1_LOC_780/Y 0.05fF
C60444 INVX1_LOC_31/A INVX1_LOC_315/Y 0.27fF
C60445 INVX1_LOC_30/A INVX1_LOC_309/A 0.06fF
C60446 NAND2X1_LOC_53/Y NOR2X1_LOC_486/Y 0.07fF
C60447 INVX1_LOC_135/A NOR2X1_LOC_6/B 0.26fF
C60448 NOR2X1_LOC_666/Y INVX1_LOC_76/A 0.01fF
C60449 NOR2X1_LOC_13/Y NAND2X1_LOC_327/a_36_24# 0.00fF
C60450 NOR2X1_LOC_852/Y NOR2X1_LOC_863/A 0.02fF
C60451 INVX1_LOC_24/A NOR2X1_LOC_322/Y 0.16fF
C60452 INVX1_LOC_226/Y INVX1_LOC_40/A 0.10fF
C60453 INVX1_LOC_226/Y INVX1_LOC_165/Y 0.02fF
C60454 NAND2X1_LOC_195/Y INVX1_LOC_6/A 0.00fF
C60455 INVX1_LOC_34/A INVX1_LOC_313/Y 0.04fF
C60456 INVX1_LOC_50/Y INVX1_LOC_280/A 0.07fF
C60457 INVX1_LOC_256/A NAND2X1_LOC_447/Y 0.10fF
C60458 INVX1_LOC_251/A INVX1_LOC_42/A 0.07fF
C60459 NOR2X1_LOC_75/Y NOR2X1_LOC_300/a_36_216# 0.00fF
C60460 INVX1_LOC_30/A INVX1_LOC_91/A 0.51fF
C60461 NOR2X1_LOC_430/A NAND2X1_LOC_51/B 0.04fF
C60462 INVX1_LOC_304/Y INVX1_LOC_90/A 0.51fF
C60463 NAND2X1_LOC_798/A INVX1_LOC_10/A 0.01fF
C60464 NOR2X1_LOC_644/A INVX1_LOC_104/A 0.03fF
C60465 NAND2X1_LOC_84/Y NOR2X1_LOC_83/Y 0.12fF
C60466 INVX1_LOC_77/A NOR2X1_LOC_74/A 0.10fF
C60467 INVX1_LOC_53/A NOR2X1_LOC_841/A 0.02fF
C60468 INVX1_LOC_13/A NOR2X1_LOC_619/A 0.05fF
C60469 NOR2X1_LOC_690/A NAND2X1_LOC_560/A 0.01fF
C60470 INVX1_LOC_18/A NOR2X1_LOC_528/Y 0.03fF
C60471 INVX1_LOC_17/A NOR2X1_LOC_111/A 0.14fF
C60472 INVX1_LOC_161/Y INVX1_LOC_46/A 0.16fF
C60473 INVX1_LOC_26/A NAND2X1_LOC_81/B 0.04fF
C60474 INVX1_LOC_293/A INVX1_LOC_2/Y 0.01fF
C60475 NAND2X1_LOC_726/Y INVX1_LOC_10/A 0.08fF
C60476 NOR2X1_LOC_507/B INVX1_LOC_210/A -0.06fF
C60477 NAND2X1_LOC_660/Y NAND2X1_LOC_662/Y 0.01fF
C60478 INVX1_LOC_2/A D_GATE_366 0.03fF
C60479 INVX1_LOC_77/A NOR2X1_LOC_9/Y 0.07fF
C60480 INVX1_LOC_75/A NOR2X1_LOC_486/B 0.19fF
C60481 INVX1_LOC_75/A NOR2X1_LOC_516/Y 0.08fF
C60482 INVX1_LOC_36/A NOR2X1_LOC_275/A 0.02fF
C60483 NOR2X1_LOC_15/Y NOR2X1_LOC_331/B 0.09fF
C60484 INVX1_LOC_230/Y VDD 1.57fF
C60485 INVX1_LOC_11/A INVX1_LOC_33/Y 0.10fF
C60486 INVX1_LOC_141/Y INVX1_LOC_20/A 0.03fF
C60487 NOR2X1_LOC_61/B NOR2X1_LOC_61/Y 0.11fF
C60488 NOR2X1_LOC_89/A INVX1_LOC_23/Y 0.20fF
C60489 NOR2X1_LOC_668/Y NAND2X1_LOC_207/B 0.01fF
C60490 INVX1_LOC_290/A NOR2X1_LOC_586/a_36_216# 0.01fF
C60491 INVX1_LOC_24/A NOR2X1_LOC_562/B 0.03fF
C60492 NOR2X1_LOC_705/a_36_216# INVX1_LOC_91/A 0.00fF
C60493 INVX1_LOC_208/A INVX1_LOC_313/A 0.00fF
C60494 NOR2X1_LOC_589/A NAND2X1_LOC_656/Y 0.07fF
C60495 NOR2X1_LOC_246/A INVX1_LOC_53/Y 0.19fF
C60496 INVX1_LOC_312/Y INVX1_LOC_20/A 0.09fF
C60497 NAND2X1_LOC_708/Y INVX1_LOC_84/A 0.01fF
C60498 NOR2X1_LOC_389/B NOR2X1_LOC_566/Y 0.03fF
C60499 INVX1_LOC_2/A NOR2X1_LOC_289/Y 0.02fF
C60500 NAND2X1_LOC_514/a_36_24# NOR2X1_LOC_106/A 0.00fF
C60501 INVX1_LOC_269/A NOR2X1_LOC_656/Y 0.03fF
C60502 NOR2X1_LOC_599/A INVX1_LOC_46/A 0.03fF
C60503 NOR2X1_LOC_780/A VDD -0.00fF
C60504 INVX1_LOC_263/A NOR2X1_LOC_644/A 0.01fF
C60505 NAND2X1_LOC_724/A INVX1_LOC_185/A 0.01fF
C60506 NAND2X1_LOC_9/Y INVX1_LOC_19/A 2.62fF
C60507 INVX1_LOC_124/A NOR2X1_LOC_74/A 0.09fF
C60508 INVX1_LOC_21/A NAND2X1_LOC_85/Y 0.07fF
C60509 INVX1_LOC_233/A INVX1_LOC_19/A 0.07fF
C60510 NOR2X1_LOC_791/Y NOR2X1_LOC_179/Y 0.17fF
C60511 INPUT_0 NAND2X1_LOC_633/a_36_24# 0.01fF
C60512 NOR2X1_LOC_616/Y NOR2X1_LOC_19/Y 0.15fF
C60513 NAND2X1_LOC_567/Y INVX1_LOC_291/Y 0.09fF
C60514 INVX1_LOC_21/A NOR2X1_LOC_697/Y 0.12fF
C60515 NOR2X1_LOC_180/B NOR2X1_LOC_569/Y 0.02fF
C60516 NOR2X1_LOC_32/B NAND2X1_LOC_74/B 0.04fF
C60517 INVX1_LOC_36/A INVX1_LOC_12/Y 0.01fF
C60518 NOR2X1_LOC_441/Y NOR2X1_LOC_366/a_36_216# 0.03fF
C60519 INVX1_LOC_124/A NOR2X1_LOC_9/Y 0.15fF
C60520 INPUT_0 NOR2X1_LOC_537/Y 0.07fF
C60521 D_INPUT_0 NAND2X1_LOC_364/a_36_24# 0.01fF
C60522 NAND2X1_LOC_803/B INVX1_LOC_54/A 0.02fF
C60523 NAND2X1_LOC_338/B INPUT_0 0.11fF
C60524 INVX1_LOC_24/A NAND2X1_LOC_836/Y 0.02fF
C60525 INVX1_LOC_30/A NOR2X1_LOC_698/Y 0.03fF
C60526 NOR2X1_LOC_65/B INVX1_LOC_251/A 0.01fF
C60527 NAND2X1_LOC_733/Y INVX1_LOC_38/A 0.02fF
C60528 INVX1_LOC_36/A NOR2X1_LOC_492/Y 0.08fF
C60529 NOR2X1_LOC_590/A NOR2X1_LOC_602/B 0.01fF
C60530 NOR2X1_LOC_152/Y NAND2X1_LOC_469/B 0.01fF
C60531 INVX1_LOC_26/A INVX1_LOC_4/Y 0.08fF
C60532 NAND2X1_LOC_796/B NOR2X1_LOC_661/A 0.02fF
C60533 INVX1_LOC_228/A D_INPUT_3 0.01fF
C60534 INVX1_LOC_90/A NAND2X1_LOC_808/A 0.08fF
C60535 NOR2X1_LOC_590/A INVX1_LOC_54/A 0.19fF
C60536 INVX1_LOC_278/A NOR2X1_LOC_76/B 0.00fF
C60537 NOR2X1_LOC_419/Y INVX1_LOC_176/A 0.90fF
C60538 NOR2X1_LOC_270/Y INVX1_LOC_202/Y 0.02fF
C60539 NOR2X1_LOC_457/B NAND2X1_LOC_472/Y 0.24fF
C60540 NOR2X1_LOC_798/A INVX1_LOC_19/A 1.52fF
C60541 NAND2X1_LOC_507/a_36_24# NOR2X1_LOC_387/A 0.00fF
C60542 NOR2X1_LOC_137/A NOR2X1_LOC_768/a_36_216# 0.00fF
C60543 NOR2X1_LOC_591/Y NAND2X1_LOC_655/A 0.30fF
C60544 INVX1_LOC_269/A NOR2X1_LOC_642/a_36_216# 0.00fF
C60545 NOR2X1_LOC_705/B INVX1_LOC_92/A 0.05fF
C60546 INVX1_LOC_217/A NAND2X1_LOC_849/B 0.10fF
C60547 NOR2X1_LOC_753/Y NOR2X1_LOC_305/Y 0.07fF
C60548 NAND2X1_LOC_3/B NAND2X1_LOC_40/a_36_24# 0.00fF
C60549 NAND2X1_LOC_733/Y NOR2X1_LOC_51/A 0.08fF
C60550 INVX1_LOC_89/A NOR2X1_LOC_163/A 0.02fF
C60551 INVX1_LOC_217/A INVX1_LOC_38/A 0.76fF
C60552 NAND2X1_LOC_763/a_36_24# NOR2X1_LOC_467/A 0.01fF
C60553 INVX1_LOC_208/A INVX1_LOC_6/A 0.11fF
C60554 NOR2X1_LOC_285/B INVX1_LOC_143/Y 0.01fF
C60555 NAND2X1_LOC_483/Y INVX1_LOC_20/A 0.03fF
C60556 NAND2X1_LOC_355/Y INVX1_LOC_38/A 0.00fF
C60557 NOR2X1_LOC_264/a_36_216# INVX1_LOC_63/A 0.01fF
C60558 NOR2X1_LOC_569/A NOR2X1_LOC_569/Y 0.03fF
C60559 NOR2X1_LOC_354/Y NOR2X1_LOC_325/A 0.05fF
C60560 NAND2X1_LOC_325/Y NOR2X1_LOC_305/Y 0.07fF
C60561 INVX1_LOC_269/A INVX1_LOC_63/A 0.15fF
C60562 INVX1_LOC_24/A INVX1_LOC_281/Y 0.01fF
C60563 NOR2X1_LOC_734/a_36_216# INVX1_LOC_1/Y 0.00fF
C60564 NOR2X1_LOC_718/Y INVX1_LOC_139/Y 0.01fF
C60565 NAND2X1_LOC_722/A INVX1_LOC_11/Y 0.07fF
C60566 D_INPUT_3 INVX1_LOC_8/A 0.00fF
C60567 NOR2X1_LOC_717/Y NOR2X1_LOC_155/A 0.01fF
C60568 INVX1_LOC_24/A INVX1_LOC_193/A 0.03fF
C60569 INVX1_LOC_256/Y INVX1_LOC_304/A 0.01fF
C60570 NOR2X1_LOC_496/Y INVX1_LOC_42/A 0.01fF
C60571 NOR2X1_LOC_473/B NOR2X1_LOC_216/Y 0.08fF
C60572 NOR2X1_LOC_441/Y INVX1_LOC_285/A 0.07fF
C60573 NOR2X1_LOC_447/A INVX1_LOC_57/A 0.04fF
C60574 NAND2X1_LOC_787/B INVX1_LOC_38/A 0.19fF
C60575 NOR2X1_LOC_309/Y INVX1_LOC_12/Y 0.03fF
C60576 INVX1_LOC_18/A NOR2X1_LOC_216/B 0.07fF
C60577 NAND2X1_LOC_741/B INVX1_LOC_297/A 0.01fF
C60578 NAND2X1_LOC_139/A NOR2X1_LOC_536/A 0.01fF
C60579 INVX1_LOC_295/A NAND2X1_LOC_328/a_36_24# 0.01fF
C60580 NAND2X1_LOC_335/a_36_24# INVX1_LOC_46/A 0.01fF
C60581 INVX1_LOC_313/Y INPUT_0 0.16fF
C60582 NOR2X1_LOC_52/B INVX1_LOC_33/Y 0.03fF
C60583 NAND2X1_LOC_9/Y INVX1_LOC_26/Y 0.07fF
C60584 NAND2X1_LOC_20/B NOR2X1_LOC_33/B 0.08fF
C60585 NAND2X1_LOC_354/Y NOR2X1_LOC_697/Y 0.02fF
C60586 NAND2X1_LOC_535/a_36_24# INVX1_LOC_264/A 0.00fF
C60587 NOR2X1_LOC_709/A INVX1_LOC_117/A 0.06fF
C60588 NOR2X1_LOC_6/B INVX1_LOC_280/A 0.02fF
C60589 INVX1_LOC_192/A NAND2X1_LOC_427/a_36_24# 0.00fF
C60590 INVX1_LOC_77/A NOR2X1_LOC_650/a_36_216# 0.00fF
C60591 NOR2X1_LOC_160/B NOR2X1_LOC_633/A 0.00fF
C60592 NOR2X1_LOC_219/Y NOR2X1_LOC_357/Y 0.17fF
C60593 INVX1_LOC_288/Y NOR2X1_LOC_639/B 0.04fF
C60594 INVX1_LOC_304/Y INVX1_LOC_38/A 0.07fF
C60595 NOR2X1_LOC_644/A INVX1_LOC_206/Y 0.03fF
C60596 NOR2X1_LOC_312/Y NOR2X1_LOC_45/B 0.04fF
C60597 NOR2X1_LOC_749/a_36_216# NOR2X1_LOC_78/A 0.00fF
C60598 INVX1_LOC_35/A INVX1_LOC_50/A 1.75fF
C60599 D_INPUT_2 NAND2X1_LOC_141/Y 0.13fF
C60600 NAND2X1_LOC_341/A VDD -0.00fF
C60601 INVX1_LOC_31/A NAND2X1_LOC_207/B 0.08fF
C60602 NOR2X1_LOC_811/B NOR2X1_LOC_319/B 0.01fF
C60603 INVX1_LOC_45/A INVX1_LOC_49/Y 0.06fF
C60604 INVX1_LOC_33/A INVX1_LOC_307/A 0.07fF
C60605 INVX1_LOC_77/A NOR2X1_LOC_865/Y 0.72fF
C60606 INVX1_LOC_35/A NOR2X1_LOC_105/Y 0.05fF
C60607 INVX1_LOC_135/A NOR2X1_LOC_124/A 0.02fF
C60608 INVX1_LOC_2/A NOR2X1_LOC_142/a_36_216# 0.00fF
C60609 NOR2X1_LOC_590/A NAND2X1_LOC_807/B 0.00fF
C60610 INVX1_LOC_225/A INVX1_LOC_185/A 0.00fF
C60611 NAND2X1_LOC_564/B INVX1_LOC_37/A 0.07fF
C60612 NOR2X1_LOC_357/Y NOR2X1_LOC_665/A 0.14fF
C60613 NAND2X1_LOC_149/Y NOR2X1_LOC_158/Y 0.08fF
C60614 INVX1_LOC_41/A INVX1_LOC_179/A 0.13fF
C60615 INVX1_LOC_53/A NOR2X1_LOC_493/a_36_216# 0.01fF
C60616 INVX1_LOC_77/A NOR2X1_LOC_243/B 0.08fF
C60617 NOR2X1_LOC_147/B INVX1_LOC_92/A 0.03fF
C60618 GATE_479 VDD 0.03fF
C60619 NOR2X1_LOC_798/A INVX1_LOC_26/Y 0.02fF
C60620 INVX1_LOC_33/A NOR2X1_LOC_445/B 0.15fF
C60621 INVX1_LOC_58/A NAND2X1_LOC_569/B 0.15fF
C60622 GATE_662 INVX1_LOC_37/A 0.01fF
C60623 INVX1_LOC_176/Y NOR2X1_LOC_461/A 0.01fF
C60624 INVX1_LOC_45/A INVX1_LOC_99/A 0.03fF
C60625 NOR2X1_LOC_644/A NOR2X1_LOC_600/Y 0.01fF
C60626 INVX1_LOC_196/A NOR2X1_LOC_729/A 0.21fF
C60627 NOR2X1_LOC_530/Y INVX1_LOC_3/Y 0.01fF
C60628 INVX1_LOC_13/Y NAND2X1_LOC_90/a_36_24# 0.00fF
C60629 NOR2X1_LOC_130/a_36_216# INVX1_LOC_74/A 0.00fF
C60630 NOR2X1_LOC_643/A NAND2X1_LOC_223/A 0.02fF
C60631 NOR2X1_LOC_186/Y INVX1_LOC_270/Y 1.43fF
C60632 NOR2X1_LOC_130/Y INVX1_LOC_59/Y 0.00fF
C60633 D_GATE_222 INVX1_LOC_38/A 0.00fF
C60634 INVX1_LOC_266/A NOR2X1_LOC_541/B 0.00fF
C60635 NOR2X1_LOC_303/Y INVX1_LOC_186/Y 0.01fF
C60636 NOR2X1_LOC_107/Y INVX1_LOC_4/Y 0.01fF
C60637 D_INPUT_1 INVX1_LOC_13/Y 0.15fF
C60638 NOR2X1_LOC_714/Y INVX1_LOC_307/A -0.01fF
C60639 NOR2X1_LOC_287/A NOR2X1_LOC_729/A 0.08fF
C60640 INVX1_LOC_313/A NAND2X1_LOC_211/Y 0.01fF
C60641 NAND2X1_LOC_139/A NOR2X1_LOC_649/B 0.01fF
C60642 NOR2X1_LOC_486/Y NOR2X1_LOC_302/Y 0.02fF
C60643 INVX1_LOC_25/A NOR2X1_LOC_789/B 0.01fF
C60644 NOR2X1_LOC_173/Y INVX1_LOC_271/A 0.02fF
C60645 NOR2X1_LOC_226/A INVX1_LOC_70/A -0.01fF
C60646 NOR2X1_LOC_488/Y INVX1_LOC_54/A 0.02fF
C60647 INVX1_LOC_34/Y NOR2X1_LOC_216/B 0.18fF
C60648 NOR2X1_LOC_142/Y NOR2X1_LOC_814/A 0.03fF
C60649 NOR2X1_LOC_829/Y NAND2X1_LOC_303/Y 0.01fF
C60650 INVX1_LOC_11/A INVX1_LOC_23/Y 0.07fF
C60651 NAND2X1_LOC_218/B NOR2X1_LOC_610/Y 0.02fF
C60652 INVX1_LOC_196/Y VDD 0.08fF
C60653 INVX1_LOC_177/A NOR2X1_LOC_800/a_36_216# 0.00fF
C60654 NAND2X1_LOC_555/Y INVX1_LOC_90/Y 0.02fF
C60655 INVX1_LOC_299/A NOR2X1_LOC_809/A 0.01fF
C60656 INVX1_LOC_48/A NOR2X1_LOC_845/A 0.39fF
C60657 NOR2X1_LOC_254/Y INVX1_LOC_186/Y 0.17fF
C60658 NOR2X1_LOC_781/A NAND2X1_LOC_637/Y 0.24fF
C60659 NAND2X1_LOC_564/B NOR2X1_LOC_177/Y 0.01fF
C60660 NOR2X1_LOC_99/B NOR2X1_LOC_862/a_36_216# 0.01fF
C60661 NOR2X1_LOC_772/B NOR2X1_LOC_652/Y 0.61fF
C60662 INVX1_LOC_280/Y INVX1_LOC_260/Y 0.01fF
C60663 NOR2X1_LOC_78/B NOR2X1_LOC_841/A 0.12fF
C60664 NAND2X1_LOC_808/A INVX1_LOC_38/A 0.07fF
C60665 INVX1_LOC_103/A NOR2X1_LOC_654/A 0.02fF
C60666 NOR2X1_LOC_180/B NAND2X1_LOC_472/Y 0.03fF
C60667 INVX1_LOC_214/A NOR2X1_LOC_697/Y 0.00fF
C60668 INVX1_LOC_10/A NOR2X1_LOC_351/Y 0.01fF
C60669 NAND2X1_LOC_198/B INVX1_LOC_32/A 0.16fF
C60670 NOR2X1_LOC_725/A NOR2X1_LOC_685/A 0.02fF
C60671 INVX1_LOC_33/A INVX1_LOC_12/A 0.26fF
C60672 D_INPUT_1 INVX1_LOC_88/A 0.09fF
C60673 INVX1_LOC_227/A INVX1_LOC_54/A 0.08fF
C60674 NAND2X1_LOC_740/B VDD 0.30fF
C60675 NAND2X1_LOC_549/Y INVX1_LOC_48/Y 0.00fF
C60676 INVX1_LOC_13/Y NOR2X1_LOC_652/Y 0.01fF
C60677 NOR2X1_LOC_256/Y VDD 0.18fF
C60678 INVX1_LOC_5/A INVX1_LOC_178/A 0.03fF
C60679 NOR2X1_LOC_655/B NOR2X1_LOC_814/A 0.98fF
C60680 NAND2X1_LOC_740/B NAND2X1_LOC_800/A 0.03fF
C60681 NAND2X1_LOC_9/a_36_24# INVX1_LOC_27/Y 0.00fF
C60682 INVX1_LOC_69/Y NAND2X1_LOC_447/Y 0.10fF
C60683 NOR2X1_LOC_720/B NAND2X1_LOC_74/B 0.10fF
C60684 INVX1_LOC_169/A INVX1_LOC_166/Y 0.05fF
C60685 NOR2X1_LOC_160/B INVX1_LOC_270/A 2.01fF
C60686 INVX1_LOC_314/Y INVX1_LOC_47/Y 0.00fF
C60687 INVX1_LOC_58/A NOR2X1_LOC_530/Y 0.11fF
C60688 NOR2X1_LOC_292/Y VDD 0.00fF
C60689 NOR2X1_LOC_346/B NOR2X1_LOC_721/B 0.04fF
C60690 NAND2X1_LOC_563/A INVX1_LOC_63/A 0.10fF
C60691 NOR2X1_LOC_356/A INVX1_LOC_9/A 0.09fF
C60692 NAND2X1_LOC_354/B NOR2X1_LOC_48/B 0.18fF
C60693 INVX1_LOC_6/A NAND2X1_LOC_211/Y 0.10fF
C60694 INVX1_LOC_224/Y NAND2X1_LOC_208/B 0.02fF
C60695 INVX1_LOC_286/A NAND2X1_LOC_650/B 0.10fF
C60696 INVX1_LOC_17/A INVX1_LOC_138/Y 0.33fF
C60697 NOR2X1_LOC_790/B NOR2X1_LOC_794/B 0.01fF
C60698 NOR2X1_LOC_543/a_36_216# NAND2X1_LOC_447/Y 0.14fF
C60699 INVX1_LOC_90/A INVX1_LOC_92/A 2.03fF
C60700 INVX1_LOC_88/A NOR2X1_LOC_652/Y 0.04fF
C60701 INVX1_LOC_2/A INVX1_LOC_102/A 0.07fF
C60702 NOR2X1_LOC_389/B INVX1_LOC_92/A 0.07fF
C60703 NOR2X1_LOC_739/Y NOR2X1_LOC_840/A 0.06fF
C60704 NAND2X1_LOC_798/A INVX1_LOC_12/A 0.01fF
C60705 NOR2X1_LOC_113/B INVX1_LOC_66/Y 0.04fF
C60706 NOR2X1_LOC_226/A INVX1_LOC_102/A 0.07fF
C60707 INVX1_LOC_64/A INVX1_LOC_39/Y 0.00fF
C60708 NOR2X1_LOC_237/Y NOR2X1_LOC_89/Y -0.01fF
C60709 NOR2X1_LOC_74/A INVX1_LOC_9/A 0.10fF
C60710 INVX1_LOC_17/A NOR2X1_LOC_272/Y 0.10fF
C60711 NOR2X1_LOC_516/B NOR2X1_LOC_633/A 0.21fF
C60712 NAND2X1_LOC_726/Y INVX1_LOC_12/A 0.01fF
C60713 INVX1_LOC_315/A INVX1_LOC_4/Y 0.16fF
C60714 INPUT_1 INVX1_LOC_123/Y 0.00fF
C60715 NOR2X1_LOC_99/B NOR2X1_LOC_814/A 0.07fF
C60716 INVX1_LOC_63/Y INVX1_LOC_78/A 0.03fF
C60717 NAND2X1_LOC_493/Y NAND2X1_LOC_561/B 0.04fF
C60718 NAND2X1_LOC_218/B NAND2X1_LOC_218/a_36_24# 0.00fF
C60719 INVX1_LOC_249/A NOR2X1_LOC_658/a_36_216# 0.00fF
C60720 INVX1_LOC_232/A NOR2X1_LOC_89/A 0.03fF
C60721 NOR2X1_LOC_657/a_36_216# INVX1_LOC_256/A 0.01fF
C60722 NOR2X1_LOC_9/Y INVX1_LOC_9/A 0.03fF
C60723 NOR2X1_LOC_205/Y NOR2X1_LOC_666/A 0.01fF
C60724 NOR2X1_LOC_87/Y INVX1_LOC_15/A 0.10fF
C60725 NAND2X1_LOC_451/Y D_INPUT_5 0.07fF
C60726 INVX1_LOC_178/A NOR2X1_LOC_816/A 0.10fF
C60727 NOR2X1_LOC_814/Y INVX1_LOC_63/A 0.04fF
C60728 NOR2X1_LOC_337/a_36_216# NAND2X1_LOC_72/B 0.00fF
C60729 NOR2X1_LOC_487/a_36_216# INVX1_LOC_278/A 0.01fF
C60730 NOR2X1_LOC_68/A NOR2X1_LOC_392/Y 0.08fF
C60731 NOR2X1_LOC_274/Y INVX1_LOC_57/A 0.01fF
C60732 INVX1_LOC_149/A INVX1_LOC_4/Y 0.09fF
C60733 NOR2X1_LOC_78/A NOR2X1_LOC_536/A 0.07fF
C60734 NOR2X1_LOC_498/Y NOR2X1_LOC_693/Y 0.00fF
C60735 INVX1_LOC_1/A D_GATE_741 0.00fF
C60736 NOR2X1_LOC_813/Y NOR2X1_LOC_124/A 0.16fF
C60737 NOR2X1_LOC_647/A NOR2X1_LOC_664/Y 0.03fF
C60738 NOR2X1_LOC_477/a_36_216# NAND2X1_LOC_149/Y 0.01fF
C60739 NOR2X1_LOC_667/Y NAND2X1_LOC_573/Y 0.14fF
C60740 NOR2X1_LOC_264/Y NOR2X1_LOC_668/Y 0.08fF
C60741 INVX1_LOC_287/A NOR2X1_LOC_708/B 0.14fF
C60742 NOR2X1_LOC_637/B INVX1_LOC_23/A 0.09fF
C60743 NOR2X1_LOC_188/A NOR2X1_LOC_831/B 0.07fF
C60744 INVX1_LOC_53/Y INVX1_LOC_32/A 0.07fF
C60745 NOR2X1_LOC_366/Y NOR2X1_LOC_89/A 0.00fF
C60746 NAND2X1_LOC_807/Y NOR2X1_LOC_605/A 0.15fF
C60747 NAND2X1_LOC_170/a_36_24# INVX1_LOC_30/A 0.00fF
C60748 INVX1_LOC_1/A NOR2X1_LOC_785/A 0.00fF
C60749 NOR2X1_LOC_52/B INVX1_LOC_23/Y 0.02fF
C60750 NOR2X1_LOC_294/Y NAND2X1_LOC_27/a_36_24# 0.00fF
C60751 NOR2X1_LOC_653/B INVX1_LOC_36/A 0.02fF
C60752 INVX1_LOC_123/A NOR2X1_LOC_99/Y 0.01fF
C60753 INVX1_LOC_65/Y NAND2X1_LOC_63/Y 0.02fF
C60754 NAND2X1_LOC_739/B NAND2X1_LOC_725/A 0.08fF
C60755 INVX1_LOC_34/A INVX1_LOC_224/Y 0.07fF
C60756 NOR2X1_LOC_75/Y INVX1_LOC_103/A 0.01fF
C60757 NOR2X1_LOC_204/a_36_216# NOR2X1_LOC_392/Y 0.00fF
C60758 NOR2X1_LOC_124/A INVX1_LOC_280/A 0.02fF
C60759 INVX1_LOC_155/A INVX1_LOC_23/A 0.09fF
C60760 NAND2X1_LOC_842/B INVX1_LOC_19/A 0.01fF
C60761 NOR2X1_LOC_212/a_36_216# NOR2X1_LOC_360/Y 0.01fF
C60762 INVX1_LOC_93/A INVX1_LOC_18/A 0.07fF
C60763 INVX1_LOC_230/Y NOR2X1_LOC_361/B 0.13fF
C60764 INVX1_LOC_223/Y NOR2X1_LOC_68/A 0.01fF
C60765 NOR2X1_LOC_763/Y NOR2X1_LOC_48/B 0.08fF
C60766 NOR2X1_LOC_172/Y INVX1_LOC_53/A 0.03fF
C60767 INVX1_LOC_225/A INVX1_LOC_270/Y 0.01fF
C60768 INVX1_LOC_27/A INVX1_LOC_205/A 0.01fF
C60769 INVX1_LOC_215/Y NOR2X1_LOC_250/A 0.00fF
C60770 NOR2X1_LOC_78/A NAND2X1_LOC_93/B 0.06fF
C60771 NAND2X1_LOC_803/B NAND2X1_LOC_350/A 0.02fF
C60772 NOR2X1_LOC_261/Y NOR2X1_LOC_770/B 0.00fF
C60773 INVX1_LOC_75/A NAND2X1_LOC_782/B 0.05fF
C60774 NOR2X1_LOC_147/B INVX1_LOC_53/A 0.00fF
C60775 VDD INVX1_LOC_44/A 0.26fF
C60776 NOR2X1_LOC_218/A NOR2X1_LOC_276/Y 0.09fF
C60777 INPUT_1 INVX1_LOC_102/A 0.00fF
C60778 NOR2X1_LOC_658/Y NOR2X1_LOC_202/a_36_216# 0.02fF
C60779 NOR2X1_LOC_403/B INVX1_LOC_13/Y 0.03fF
C60780 NAND2X1_LOC_363/B NAND2X1_LOC_276/Y 0.04fF
C60781 NOR2X1_LOC_392/B INVX1_LOC_53/A 0.02fF
C60782 NAND2X1_LOC_208/B NOR2X1_LOC_103/Y 0.17fF
C60783 NOR2X1_LOC_590/A NAND2X1_LOC_350/A 0.05fF
C60784 NOR2X1_LOC_226/A NAND2X1_LOC_439/a_36_24# 0.00fF
C60785 INVX1_LOC_36/A NOR2X1_LOC_401/A 0.23fF
C60786 INVX1_LOC_16/A NOR2X1_LOC_25/Y 0.53fF
C60787 NOR2X1_LOC_261/A INVX1_LOC_37/A 0.01fF
C60788 NOR2X1_LOC_486/Y INVX1_LOC_307/A 0.02fF
C60789 NOR2X1_LOC_205/a_36_216# NOR2X1_LOC_383/B 0.00fF
C60790 NAND2X1_LOC_650/B INVX1_LOC_54/A 0.07fF
C60791 NOR2X1_LOC_604/Y INVX1_LOC_266/Y 0.01fF
C60792 NOR2X1_LOC_690/A NOR2X1_LOC_291/a_36_216# 0.00fF
C60793 NOR2X1_LOC_368/A NAND2X1_LOC_81/B 0.17fF
C60794 NOR2X1_LOC_144/a_36_216# NOR2X1_LOC_66/Y 0.00fF
C60795 VDD NOR2X1_LOC_641/Y 0.20fF
C60796 NOR2X1_LOC_76/a_36_216# INVX1_LOC_32/A 0.12fF
C60797 INVX1_LOC_17/A NAND2X1_LOC_364/A 0.25fF
C60798 NOR2X1_LOC_590/A NOR2X1_LOC_441/Y 0.02fF
C60799 INVX1_LOC_208/A INVX1_LOC_270/A 0.10fF
C60800 NOR2X1_LOC_78/A INVX1_LOC_3/A 4.64fF
C60801 NOR2X1_LOC_230/Y NOR2X1_LOC_45/Y 0.04fF
C60802 NOR2X1_LOC_355/A INVX1_LOC_94/Y 0.02fF
C60803 NOR2X1_LOC_186/Y NAND2X1_LOC_300/a_36_24# 0.00fF
C60804 NAND2X1_LOC_850/a_36_24# NAND2X1_LOC_474/Y 0.00fF
C60805 NOR2X1_LOC_500/Y NOR2X1_LOC_748/A 0.05fF
C60806 NOR2X1_LOC_513/Y INVX1_LOC_18/A 0.01fF
C60807 INVX1_LOC_135/A INVX1_LOC_273/A 0.01fF
C60808 INVX1_LOC_5/A NAND2X1_LOC_562/B 0.52fF
C60809 INVX1_LOC_36/A NOR2X1_LOC_160/B 0.17fF
C60810 INVX1_LOC_64/A NOR2X1_LOC_168/B 0.03fF
C60811 NAND2X1_LOC_350/A NAND2X1_LOC_589/a_36_24# 0.01fF
C60812 INVX1_LOC_316/Y INVX1_LOC_23/A 0.03fF
C60813 NOR2X1_LOC_502/a_36_216# NOR2X1_LOC_814/A 0.01fF
C60814 NOR2X1_LOC_215/A INVX1_LOC_63/Y 0.03fF
C60815 INVX1_LOC_45/A NAND2X1_LOC_208/B 0.46fF
C60816 NOR2X1_LOC_848/Y NOR2X1_LOC_860/B 0.01fF
C60817 INVX1_LOC_90/A NAND2X1_LOC_247/a_36_24# 0.00fF
C60818 NOR2X1_LOC_653/B NOR2X1_LOC_309/Y 0.01fF
C60819 NOR2X1_LOC_858/B NOR2X1_LOC_862/B 0.03fF
C60820 NAND2X1_LOC_573/Y NAND2X1_LOC_300/a_36_24# 0.00fF
C60821 NAND2X1_LOC_537/Y NOR2X1_LOC_577/Y 0.34fF
C60822 INVX1_LOC_178/A NAND2X1_LOC_562/B 0.13fF
C60823 INVX1_LOC_224/A NAND2X1_LOC_517/a_36_24# 0.00fF
C60824 NAND2X1_LOC_714/B NAND2X1_LOC_799/Y 0.08fF
C60825 NAND2X1_LOC_860/A INVX1_LOC_22/A 0.02fF
C60826 NOR2X1_LOC_609/A INVX1_LOC_292/A 0.01fF
C60827 INVX1_LOC_222/Y NOR2X1_LOC_802/A 0.04fF
C60828 NOR2X1_LOC_841/A INVX1_LOC_46/A 0.01fF
C60829 NOR2X1_LOC_211/a_36_216# INVX1_LOC_22/A 0.00fF
C60830 NOR2X1_LOC_15/Y NOR2X1_LOC_388/Y 0.07fF
C60831 NOR2X1_LOC_250/Y INVX1_LOC_77/A 0.20fF
C60832 NAND2X1_LOC_552/A NOR2X1_LOC_773/Y 0.01fF
C60833 NOR2X1_LOC_208/Y NOR2X1_LOC_160/B 0.10fF
C60834 NOR2X1_LOC_80/a_36_216# NAND2X1_LOC_63/Y 0.00fF
C60835 NOR2X1_LOC_237/Y NAND2X1_LOC_550/A 0.01fF
C60836 INVX1_LOC_1/A NOR2X1_LOC_514/Y 0.02fF
C60837 INVX1_LOC_38/A INVX1_LOC_92/A 0.17fF
C60838 INVX1_LOC_34/A NOR2X1_LOC_103/Y 0.07fF
C60839 INVX1_LOC_75/A NAND2X1_LOC_454/Y 0.10fF
C60840 NOR2X1_LOC_231/B INVX1_LOC_314/Y 0.01fF
C60841 INVX1_LOC_72/A INVX1_LOC_72/Y 0.01fF
C60842 NOR2X1_LOC_506/a_36_216# NOR2X1_LOC_697/Y 0.00fF
C60843 NOR2X1_LOC_644/Y NOR2X1_LOC_348/Y 0.04fF
C60844 INVX1_LOC_244/Y INVX1_LOC_30/A 0.06fF
C60845 INVX1_LOC_178/A NOR2X1_LOC_773/Y 0.10fF
C60846 NOR2X1_LOC_160/B NOR2X1_LOC_804/B 0.07fF
C60847 NAND2X1_LOC_725/Y INVX1_LOC_173/Y 0.15fF
C60848 INVX1_LOC_8/Y INVX1_LOC_31/A 0.37fF
C60849 INVX1_LOC_224/A NAND2X1_LOC_116/A 0.02fF
C60850 NOR2X1_LOC_794/B NOR2X1_LOC_344/A 0.02fF
C60851 INVX1_LOC_59/A NOR2X1_LOC_67/A 0.01fF
C60852 NOR2X1_LOC_596/Y NOR2X1_LOC_593/Y 0.03fF
C60853 INVX1_LOC_119/A INVX1_LOC_272/Y 0.10fF
C60854 NOR2X1_LOC_719/A INVX1_LOC_306/Y 0.01fF
C60855 INVX1_LOC_11/A NAND2X1_LOC_116/A 0.03fF
C60856 INVX1_LOC_12/Y INVX1_LOC_63/A 0.07fF
C60857 NOR2X1_LOC_649/a_36_216# INVX1_LOC_31/A 0.00fF
C60858 INVX1_LOC_64/A NAND2X1_LOC_656/Y 0.36fF
C60859 NOR2X1_LOC_865/Y INVX1_LOC_9/A 0.07fF
C60860 INVX1_LOC_171/A NOR2X1_LOC_717/A 0.01fF
C60861 NOR2X1_LOC_557/A INVX1_LOC_47/Y 0.00fF
C60862 NOR2X1_LOC_590/A NOR2X1_LOC_340/Y 0.04fF
C60863 INVX1_LOC_288/Y INVX1_LOC_302/A 0.24fF
C60864 NOR2X1_LOC_590/A NOR2X1_LOC_142/Y 0.07fF
C60865 NOR2X1_LOC_243/B INVX1_LOC_9/A 0.07fF
C60866 NOR2X1_LOC_91/Y INVX1_LOC_41/Y 0.07fF
C60867 INVX1_LOC_22/A INVX1_LOC_242/A 0.49fF
C60868 INVX1_LOC_90/A INVX1_LOC_53/A 3.42fF
C60869 NOR2X1_LOC_160/B NOR2X1_LOC_309/Y 0.03fF
C60870 INVX1_LOC_10/A NOR2X1_LOC_304/Y 0.01fF
C60871 INVX1_LOC_18/A NOR2X1_LOC_303/Y 0.10fF
C60872 NAND2X1_LOC_769/a_36_24# INVX1_LOC_53/A 0.00fF
C60873 NAND2X1_LOC_774/a_36_24# NOR2X1_LOC_226/A 0.00fF
C60874 NAND2X1_LOC_850/A INVX1_LOC_23/A 1.20fF
C60875 NOR2X1_LOC_286/Y INVX1_LOC_196/A 1.78fF
C60876 NOR2X1_LOC_264/Y INVX1_LOC_31/A 0.23fF
C60877 NOR2X1_LOC_389/B INVX1_LOC_53/A 0.01fF
C60878 INVX1_LOC_5/A NOR2X1_LOC_332/A 0.22fF
C60879 INVX1_LOC_17/A NAND2X1_LOC_11/Y 0.06fF
C60880 INVX1_LOC_45/A INVX1_LOC_34/A 0.03fF
C60881 NOR2X1_LOC_471/Y NOR2X1_LOC_627/Y 0.02fF
C60882 INVX1_LOC_41/A NOR2X1_LOC_751/Y 0.01fF
C60883 NAND2X1_LOC_714/B NAND2X1_LOC_319/A 0.03fF
C60884 NAND2X1_LOC_729/Y NOR2X1_LOC_387/Y 0.11fF
C60885 INVX1_LOC_34/A NAND2X1_LOC_856/A 0.01fF
C60886 NAND2X1_LOC_537/Y INVX1_LOC_22/A 0.07fF
C60887 NOR2X1_LOC_83/Y NOR2X1_LOC_383/B 0.01fF
C60888 INVX1_LOC_269/A INVX1_LOC_1/Y 0.10fF
C60889 INVX1_LOC_224/Y INPUT_0 0.04fF
C60890 NOR2X1_LOC_690/A NAND2X1_LOC_634/Y 0.07fF
C60891 INVX1_LOC_72/A NAND2X1_LOC_811/Y 0.94fF
C60892 NOR2X1_LOC_773/Y NOR2X1_LOC_816/A 0.07fF
C60893 NOR2X1_LOC_655/B NOR2X1_LOC_590/A 0.07fF
C60894 INVX1_LOC_230/Y INVX1_LOC_280/Y 0.18fF
C60895 INVX1_LOC_11/A INVX1_LOC_232/A 0.07fF
C60896 INVX1_LOC_230/Y NOR2X1_LOC_608/a_36_216# 0.00fF
C60897 INVX1_LOC_24/A NAND2X1_LOC_833/Y 0.03fF
C60898 INVX1_LOC_86/A INVX1_LOC_23/A 0.01fF
C60899 NOR2X1_LOC_228/a_36_216# INVX1_LOC_314/Y 0.01fF
C60900 NOR2X1_LOC_155/A NOR2X1_LOC_127/Y 0.07fF
C60901 INVX1_LOC_147/Y INVX1_LOC_128/Y 0.04fF
C60902 INVX1_LOC_1/A NOR2X1_LOC_128/B 0.01fF
C60903 NAND2X1_LOC_432/a_36_24# NAND2X1_LOC_798/B 0.00fF
C60904 NOR2X1_LOC_405/A NOR2X1_LOC_301/A 0.05fF
C60905 NAND2X1_LOC_552/A INVX1_LOC_140/A 0.01fF
C60906 INVX1_LOC_256/A NAND2X1_LOC_112/Y 0.01fF
C60907 INVX1_LOC_2/A INVX1_LOC_223/A 0.03fF
C60908 INVX1_LOC_45/A NAND2X1_LOC_231/Y 0.01fF
C60909 INVX1_LOC_72/A INVX1_LOC_266/Y 0.04fF
C60910 NAND2X1_LOC_734/B NOR2X1_LOC_68/A 0.03fF
C60911 NAND2X1_LOC_860/A INVX1_LOC_100/A 0.07fF
C60912 NOR2X1_LOC_92/Y NOR2X1_LOC_71/Y 0.27fF
C60913 NOR2X1_LOC_15/Y INVX1_LOC_135/A 1.38fF
C60914 INVX1_LOC_34/A INVX1_LOC_71/A 0.10fF
C60915 NAND2X1_LOC_374/Y INVX1_LOC_30/A 0.07fF
C60916 INVX1_LOC_174/A NOR2X1_LOC_146/Y 0.03fF
C60917 NOR2X1_LOC_794/B NOR2X1_LOC_540/a_36_216# 0.00fF
C60918 NAND2X1_LOC_755/a_36_24# NOR2X1_LOC_68/A 0.01fF
C60919 NOR2X1_LOC_424/Y INVX1_LOC_103/A 0.73fF
C60920 INPUT_3 NOR2X1_LOC_619/A 0.17fF
C60921 INVX1_LOC_63/Y NOR2X1_LOC_152/Y 0.01fF
C60922 INVX1_LOC_31/A INVX1_LOC_316/Y 0.05fF
C60923 NOR2X1_LOC_82/A NOR2X1_LOC_391/A 0.01fF
C60924 INVX1_LOC_54/Y INVX1_LOC_18/A 0.08fF
C60925 NAND2X1_LOC_149/Y INVX1_LOC_55/Y 0.08fF
C60926 INVX1_LOC_63/Y INVX1_LOC_113/Y 0.01fF
C60927 INVX1_LOC_102/A INVX1_LOC_118/A 0.07fF
C60928 GATE_579 NOR2X1_LOC_298/Y 0.11fF
C60929 INVX1_LOC_178/A INVX1_LOC_140/A 0.14fF
C60930 NAND2X1_LOC_338/B INVX1_LOC_72/Y 0.03fF
C60931 INVX1_LOC_36/A INVX1_LOC_208/A 0.09fF
C60932 NAND2X1_LOC_361/Y NAND2X1_LOC_362/a_36_24# 0.01fF
C60933 INVX1_LOC_24/Y NOR2X1_LOC_644/A 0.19fF
C60934 NOR2X1_LOC_111/A INVX1_LOC_94/Y 0.03fF
C60935 INVX1_LOC_36/A NOR2X1_LOC_516/B 0.08fF
C60936 INVX1_LOC_49/A INVX1_LOC_85/A 0.00fF
C60937 NOR2X1_LOC_334/Y INVX1_LOC_117/A 0.07fF
C60938 NAND2X1_LOC_53/Y INVX1_LOC_89/A 0.07fF
C60939 NOR2X1_LOC_705/B INVX1_LOC_83/A 0.03fF
C60940 NOR2X1_LOC_799/B NOR2X1_LOC_748/A 0.08fF
C60941 NOR2X1_LOC_658/Y NOR2X1_LOC_589/A 0.07fF
C60942 NOR2X1_LOC_570/a_36_216# NOR2X1_LOC_500/Y 0.01fF
C60943 NOR2X1_LOC_152/A INVX1_LOC_273/A 0.15fF
C60944 NOR2X1_LOC_590/A NOR2X1_LOC_99/B 0.10fF
C60945 NOR2X1_LOC_643/Y NOR2X1_LOC_537/Y 0.03fF
C60946 INVX1_LOC_9/Y NAND2X1_LOC_198/B 0.03fF
C60947 NOR2X1_LOC_222/Y INVX1_LOC_81/A 0.15fF
C60948 NOR2X1_LOC_657/Y NOR2X1_LOC_561/Y 0.02fF
C60949 INVX1_LOC_215/A INVX1_LOC_177/Y 0.15fF
C60950 INVX1_LOC_227/Y NOR2X1_LOC_570/A 0.00fF
C60951 INVX1_LOC_11/A NOR2X1_LOC_775/Y 0.01fF
C60952 NOR2X1_LOC_208/Y INVX1_LOC_208/A 0.10fF
C60953 NOR2X1_LOC_524/Y NOR2X1_LOC_355/A 0.00fF
C60954 NAND2X1_LOC_468/B NOR2X1_LOC_678/A 0.03fF
C60955 NAND2X1_LOC_67/Y NOR2X1_LOC_74/A 0.03fF
C60956 NOR2X1_LOC_390/a_36_216# INVX1_LOC_177/A 0.00fF
C60957 NOR2X1_LOC_104/a_36_216# INVX1_LOC_3/Y 0.01fF
C60958 NOR2X1_LOC_861/Y NOR2X1_LOC_865/Y 0.21fF
C60959 NOR2X1_LOC_632/Y NOR2X1_LOC_596/A 0.68fF
C60960 NOR2X1_LOC_816/A INVX1_LOC_140/A 0.10fF
C60961 NOR2X1_LOC_861/Y NOR2X1_LOC_243/B 0.16fF
C60962 INVX1_LOC_91/A NOR2X1_LOC_460/Y 0.01fF
C60963 INVX1_LOC_27/Y INVX1_LOC_42/A 0.03fF
C60964 NOR2X1_LOC_78/B NOR2X1_LOC_147/B 0.17fF
C60965 INVX1_LOC_2/A INVX1_LOC_85/A 0.04fF
C60966 NOR2X1_LOC_78/B NOR2X1_LOC_392/B 0.07fF
C60967 NOR2X1_LOC_590/A INVX1_LOC_182/A 0.07fF
C60968 NOR2X1_LOC_103/Y INPUT_0 0.07fF
C60969 NOR2X1_LOC_516/B NOR2X1_LOC_804/B 0.08fF
C60970 INVX1_LOC_14/A INVX1_LOC_201/A 0.23fF
C60971 INVX1_LOC_49/A NAND2X1_LOC_662/Y 0.08fF
C60972 NOR2X1_LOC_593/Y INVX1_LOC_232/A 0.09fF
C60973 INVX1_LOC_50/Y INVX1_LOC_247/A 0.03fF
C60974 NOR2X1_LOC_169/B NOR2X1_LOC_356/A 0.03fF
C60975 INVX1_LOC_19/A INVX1_LOC_284/A 0.07fF
C60976 NOR2X1_LOC_226/A NOR2X1_LOC_316/Y -0.10fF
C60977 NAND2X1_LOC_211/Y NOR2X1_LOC_109/Y 0.32fF
C60978 D_INPUT_0 NAND2X1_LOC_101/a_36_24# 0.00fF
C60979 INVX1_LOC_21/A NOR2X1_LOC_631/B 0.07fF
C60980 INVX1_LOC_135/A NOR2X1_LOC_860/B 0.08fF
C60981 INVX1_LOC_76/A INVX1_LOC_306/Y 0.08fF
C60982 INVX1_LOC_20/A NOR2X1_LOC_649/Y 0.04fF
C60983 INVX1_LOC_24/A NOR2X1_LOC_76/A 0.04fF
C60984 INVX1_LOC_269/A NOR2X1_LOC_318/B 0.17fF
C60985 NOR2X1_LOC_433/A NOR2X1_LOC_366/Y 0.02fF
C60986 NOR2X1_LOC_106/Y NAND2X1_LOC_140/A 0.00fF
C60987 D_INPUT_0 INVX1_LOC_77/A 0.24fF
C60988 INVX1_LOC_24/A NOR2X1_LOC_180/B 0.07fF
C60989 INVX1_LOC_12/A NOR2X1_LOC_12/a_36_216# 0.01fF
C60990 INVX1_LOC_53/A INVX1_LOC_38/A 7.87fF
C60991 D_INPUT_7 D_INPUT_4 0.35fF
C60992 NAND2X1_LOC_338/B NAND2X1_LOC_334/a_36_24# 0.02fF
C60993 NOR2X1_LOC_493/B NOR2X1_LOC_500/Y 0.02fF
C60994 NOR2X1_LOC_384/Y NAND2X1_LOC_849/A 0.68fF
C60995 INVX1_LOC_227/A NOR2X1_LOC_142/Y 0.10fF
C60996 INVX1_LOC_269/A INVX1_LOC_93/Y 0.10fF
C60997 NOR2X1_LOC_172/Y INVX1_LOC_83/A 0.03fF
C60998 NOR2X1_LOC_68/A NOR2X1_LOC_439/B 0.01fF
C60999 INVX1_LOC_256/A INVX1_LOC_98/A 0.02fF
C61000 NOR2X1_LOC_860/B NOR2X1_LOC_560/A 0.01fF
C61001 NOR2X1_LOC_565/A NOR2X1_LOC_74/A 0.02fF
C61002 NOR2X1_LOC_36/B D_INPUT_5 0.01fF
C61003 INVX1_LOC_45/A INPUT_0 0.17fF
C61004 INVX1_LOC_17/A NOR2X1_LOC_405/A 0.15fF
C61005 INVX1_LOC_208/Y NAND2X1_LOC_342/Y 0.10fF
C61006 INVX1_LOC_256/A NOR2X1_LOC_78/A 0.04fF
C61007 NAND2X1_LOC_479/Y INVX1_LOC_96/Y 0.43fF
C61008 NOR2X1_LOC_522/a_36_216# NAND2X1_LOC_849/A 0.01fF
C61009 INVX1_LOC_21/A INVX1_LOC_37/A 0.31fF
C61010 NOR2X1_LOC_147/B INVX1_LOC_83/A 0.15fF
C61011 NOR2X1_LOC_68/A INVX1_LOC_75/A 1.26fF
C61012 INVX1_LOC_41/A NOR2X1_LOC_71/Y 0.49fF
C61013 INVX1_LOC_25/A NOR2X1_LOC_78/a_36_216# 0.00fF
C61014 NOR2X1_LOC_155/A NOR2X1_LOC_383/B 0.09fF
C61015 INVX1_LOC_313/A INVX1_LOC_155/A 0.21fF
C61016 INVX1_LOC_21/A NOR2X1_LOC_231/A 0.01fF
C61017 INVX1_LOC_34/A NOR2X1_LOC_123/B 0.07fF
C61018 INVX1_LOC_307/A NOR2X1_LOC_748/A 0.10fF
C61019 INVX1_LOC_251/Y INVX1_LOC_30/Y 0.04fF
C61020 NOR2X1_LOC_226/A NAND2X1_LOC_543/Y 0.01fF
C61021 INVX1_LOC_119/A INVX1_LOC_10/A 0.02fF
C61022 INVX1_LOC_271/A NAND2X1_LOC_798/B 0.00fF
C61023 NOR2X1_LOC_216/a_36_216# INVX1_LOC_77/A 0.01fF
C61024 NAND2X1_LOC_784/a_36_24# NAND2X1_LOC_721/A -0.00fF
C61025 NOR2X1_LOC_52/B NOR2X1_LOC_366/Y 0.02fF
C61026 NOR2X1_LOC_624/A INVX1_LOC_65/Y 0.00fF
C61027 NOR2X1_LOC_445/B NOR2X1_LOC_748/A 0.10fF
C61028 INVX1_LOC_72/A INVX1_LOC_191/A 0.04fF
C61029 NOR2X1_LOC_186/Y NOR2X1_LOC_536/A 0.26fF
C61030 INVX1_LOC_41/A NOR2X1_LOC_644/A 0.03fF
C61031 NAND2X1_LOC_477/A NOR2X1_LOC_71/Y 0.18fF
C61032 NOR2X1_LOC_65/B INVX1_LOC_27/Y 0.03fF
C61033 INVX1_LOC_135/A NAND2X1_LOC_141/A 0.01fF
C61034 NOR2X1_LOC_655/B INVX1_LOC_227/A 0.09fF
C61035 INVX1_LOC_36/A INVX1_LOC_315/Y 0.07fF
C61036 INVX1_LOC_15/Y INVX1_LOC_135/A 0.17fF
C61037 INPUT_0 INVX1_LOC_71/A 0.15fF
C61038 NOR2X1_LOC_91/A NOR2X1_LOC_662/A 0.02fF
C61039 INVX1_LOC_41/A NOR2X1_LOC_828/B 0.06fF
C61040 INVX1_LOC_13/A INVX1_LOC_16/A 0.06fF
C61041 NOR2X1_LOC_299/a_36_216# NAND2X1_LOC_463/B 0.00fF
C61042 NAND2X1_LOC_573/Y NOR2X1_LOC_536/A 0.28fF
C61043 NOR2X1_LOC_232/Y NAND2X1_LOC_721/A 0.33fF
C61044 INVX1_LOC_63/Y NAND2X1_LOC_661/A 0.01fF
C61045 NOR2X1_LOC_125/Y NOR2X1_LOC_127/Y 0.24fF
C61046 NOR2X1_LOC_557/Y INVX1_LOC_73/A 0.97fF
C61047 INVX1_LOC_45/A NAND2X1_LOC_649/B 0.02fF
C61048 INVX1_LOC_313/Y INVX1_LOC_266/Y 0.12fF
C61049 NOR2X1_LOC_15/Y INVX1_LOC_10/Y 0.03fF
C61050 INVX1_LOC_177/A INVX1_LOC_196/Y 0.40fF
C61051 NOR2X1_LOC_78/B INVX1_LOC_97/A 0.64fF
C61052 INVX1_LOC_308/A INVX1_LOC_285/A 0.04fF
C61053 INVX1_LOC_233/Y INVX1_LOC_260/Y 0.15fF
C61054 NAND2X1_LOC_785/B NOR2X1_LOC_164/Y 0.16fF
C61055 NAND2X1_LOC_483/Y INVX1_LOC_282/A 0.04fF
C61056 INVX1_LOC_124/A NOR2X1_LOC_216/a_36_216# 0.01fF
C61057 INVX1_LOC_41/A NOR2X1_LOC_751/A 0.28fF
C61058 NOR2X1_LOC_15/Y INVX1_LOC_280/A 0.03fF
C61059 INVX1_LOC_21/A NOR2X1_LOC_177/Y 0.05fF
C61060 INVX1_LOC_23/A NOR2X1_LOC_662/A 0.02fF
C61061 NOR2X1_LOC_855/A NOR2X1_LOC_812/A 0.19fF
C61062 NOR2X1_LOC_78/B INVX1_LOC_90/A 0.74fF
C61063 NOR2X1_LOC_389/A NAND2X1_LOC_39/Y 0.04fF
C61064 NAND2X1_LOC_356/a_36_24# NOR2X1_LOC_45/B 0.00fF
C61065 INVX1_LOC_236/A INVX1_LOC_28/A 0.18fF
C61066 INVX1_LOC_27/A NOR2X1_LOC_433/Y 0.04fF
C61067 NOR2X1_LOC_428/Y INVX1_LOC_37/A 0.01fF
C61068 INVX1_LOC_21/A NOR2X1_LOC_743/Y 0.72fF
C61069 NOR2X1_LOC_441/Y NAND2X1_LOC_650/B 0.08fF
C61070 NOR2X1_LOC_78/B NOR2X1_LOC_389/B 0.07fF
C61071 INVX1_LOC_89/A NOR2X1_LOC_500/Y 0.03fF
C61072 NOR2X1_LOC_605/B NAND2X1_LOC_808/A 0.04fF
C61073 INVX1_LOC_155/A INVX1_LOC_6/A 0.03fF
C61074 INVX1_LOC_226/Y INVX1_LOC_89/A 0.08fF
C61075 NAND2X1_LOC_361/Y NOR2X1_LOC_334/A 0.07fF
C61076 NAND2X1_LOC_254/Y INVX1_LOC_23/Y 1.25fF
C61077 NOR2X1_LOC_202/Y INVX1_LOC_96/Y 0.03fF
C61078 NOR2X1_LOC_657/Y INVX1_LOC_76/A 0.01fF
C61079 NOR2X1_LOC_92/Y NAND2X1_LOC_243/Y 0.04fF
C61080 NAND2X1_LOC_231/Y INVX1_LOC_102/Y 0.08fF
C61081 NAND2X1_LOC_569/A INVX1_LOC_6/A 0.00fF
C61082 INVX1_LOC_181/Y INVX1_LOC_95/Y 0.19fF
C61083 NOR2X1_LOC_570/B INVX1_LOC_206/Y 0.09fF
C61084 NAND2X1_LOC_715/B NOR2X1_LOC_127/Y 0.23fF
C61085 INVX1_LOC_36/A NAND2X1_LOC_211/Y 0.16fF
C61086 INVX1_LOC_83/A NOR2X1_LOC_512/a_36_216# 0.01fF
C61087 INVX1_LOC_269/Y NOR2X1_LOC_729/A 0.01fF
C61088 NOR2X1_LOC_186/Y NAND2X1_LOC_780/a_36_24# 0.00fF
C61089 INVX1_LOC_39/A INVX1_LOC_123/Y 0.01fF
C61090 NAND2X1_LOC_653/a_36_24# NAND2X1_LOC_661/B 0.00fF
C61091 INVX1_LOC_10/A INVX1_LOC_150/A 0.01fF
C61092 NOR2X1_LOC_836/Y INVX1_LOC_117/A 0.82fF
C61093 NOR2X1_LOC_773/Y INVX1_LOC_140/A 0.10fF
C61094 INVX1_LOC_55/Y INVX1_LOC_16/A 0.03fF
C61095 NAND2X1_LOC_207/B NOR2X1_LOC_416/A 0.03fF
C61096 NOR2X1_LOC_78/B NAND2X1_LOC_348/A 0.65fF
C61097 NAND2X1_LOC_182/A INVX1_LOC_286/A 0.03fF
C61098 NOR2X1_LOC_13/Y INVX1_LOC_147/Y 0.01fF
C61099 INVX1_LOC_286/A INVX1_LOC_104/A 0.00fF
C61100 NOR2X1_LOC_68/A NAND2X1_LOC_453/A 0.07fF
C61101 INVX1_LOC_89/A INVX1_LOC_10/A 0.17fF
C61102 NAND2X1_LOC_354/Y INVX1_LOC_37/A 0.02fF
C61103 INVX1_LOC_49/A NAND2X1_LOC_843/a_36_24# 0.00fF
C61104 INVX1_LOC_24/A NAND2X1_LOC_241/Y 0.01fF
C61105 INVX1_LOC_179/Y NOR2X1_LOC_74/A 0.03fF
C61106 NOR2X1_LOC_582/Y INVX1_LOC_37/A 0.12fF
C61107 NOR2X1_LOC_13/Y INVX1_LOC_20/A -0.01fF
C61108 NAND2X1_LOC_573/Y NAND2X1_LOC_780/a_36_24# 0.01fF
C61109 NAND2X1_LOC_656/A INVX1_LOC_2/Y 0.05fF
C61110 NOR2X1_LOC_130/A NOR2X1_LOC_76/A 0.07fF
C61111 NAND2X1_LOC_661/B INVX1_LOC_6/A 0.33fF
C61112 INVX1_LOC_289/A NAND2X1_LOC_51/B 0.03fF
C61113 NOR2X1_LOC_6/B NOR2X1_LOC_45/B 0.11fF
C61114 NOR2X1_LOC_596/A NAND2X1_LOC_39/Y 0.01fF
C61115 INVX1_LOC_90/A INVX1_LOC_83/A 0.24fF
C61116 NAND2X1_LOC_354/B INVX1_LOC_291/Y 0.01fF
C61117 NAND2X1_LOC_579/A INVX1_LOC_285/A 0.02fF
C61118 NOR2X1_LOC_593/Y NAND2X1_LOC_447/Y 0.40fF
C61119 INVX1_LOC_44/Y INVX1_LOC_78/Y 0.01fF
C61120 INVX1_LOC_41/A NOR2X1_LOC_540/B 0.06fF
C61121 NAND2X1_LOC_794/B INVX1_LOC_264/A 0.05fF
C61122 NOR2X1_LOC_304/Y INVX1_LOC_12/A 0.01fF
C61123 INVX1_LOC_209/Y NOR2X1_LOC_314/Y 0.01fF
C61124 INVX1_LOC_209/Y NOR2X1_LOC_422/Y 0.01fF
C61125 NOR2X1_LOC_390/a_36_216# NOR2X1_LOC_137/B 0.00fF
C61126 NOR2X1_LOC_192/a_36_216# INVX1_LOC_95/Y 0.01fF
C61127 NAND2X1_LOC_552/A INVX1_LOC_42/A 0.05fF
C61128 NOR2X1_LOC_229/Y INVX1_LOC_6/A 0.47fF
C61129 INVX1_LOC_5/A INVX1_LOC_42/A 0.06fF
C61130 NOR2X1_LOC_172/Y INVX1_LOC_46/A 0.05fF
C61131 INVX1_LOC_77/A NOR2X1_LOC_859/Y 0.02fF
C61132 NOR2X1_LOC_772/Y INVX1_LOC_46/A 0.04fF
C61133 NOR2X1_LOC_561/Y NOR2X1_LOC_74/A 0.00fF
C61134 INVX1_LOC_58/A NOR2X1_LOC_334/Y 0.10fF
C61135 NOR2X1_LOC_717/A INVX1_LOC_4/A -0.01fF
C61136 NAND2X1_LOC_348/A INVX1_LOC_83/A 0.07fF
C61137 NOR2X1_LOC_323/Y NAND2X1_LOC_808/A 0.01fF
C61138 NOR2X1_LOC_392/B INVX1_LOC_46/A 0.11fF
C61139 NOR2X1_LOC_860/B INVX1_LOC_280/A 0.06fF
C61140 INVX1_LOC_127/Y INVX1_LOC_306/Y 0.03fF
C61141 INVX1_LOC_178/A INVX1_LOC_42/A 0.02fF
C61142 NOR2X1_LOC_474/A INVX1_LOC_166/Y 0.15fF
C61143 NOR2X1_LOC_91/Y INVX1_LOC_185/A 0.02fF
C61144 INVX1_LOC_132/A NOR2X1_LOC_536/A 0.09fF
C61145 NOR2X1_LOC_504/Y INVX1_LOC_20/A 0.07fF
C61146 INVX1_LOC_144/Y NOR2X1_LOC_56/Y 0.62fF
C61147 NOR2X1_LOC_689/A NOR2X1_LOC_689/Y 0.32fF
C61148 NOR2X1_LOC_123/B INPUT_0 0.07fF
C61149 NOR2X1_LOC_397/a_36_216# INVX1_LOC_98/A 0.14fF
C61150 NOR2X1_LOC_723/a_36_216# INVX1_LOC_179/A 0.00fF
C61151 NOR2X1_LOC_111/Y NOR2X1_LOC_329/B 0.07fF
C61152 INVX1_LOC_18/A NAND2X1_LOC_656/B 0.03fF
C61153 INVX1_LOC_14/A INVX1_LOC_29/A 0.91fF
C61154 INVX1_LOC_30/A NOR2X1_LOC_103/a_36_216# 0.00fF
C61155 INVX1_LOC_75/A NOR2X1_LOC_163/A 0.00fF
C61156 NOR2X1_LOC_91/A INVX1_LOC_57/A 0.07fF
C61157 NOR2X1_LOC_668/Y INVX1_LOC_57/A 0.07fF
C61158 NOR2X1_LOC_122/A NOR2X1_LOC_755/Y 0.05fF
C61159 NOR2X1_LOC_160/B INVX1_LOC_63/A 1.21fF
C61160 NOR2X1_LOC_397/a_36_216# NOR2X1_LOC_78/A 0.00fF
C61161 NAND2X1_LOC_112/a_36_24# NAND2X1_LOC_211/Y 0.01fF
C61162 NOR2X1_LOC_360/Y NOR2X1_LOC_79/Y 0.03fF
C61163 INVX1_LOC_256/Y INVX1_LOC_20/A 0.22fF
C61164 NAND2X1_LOC_802/A NOR2X1_LOC_506/Y 0.00fF
C61165 NOR2X1_LOC_677/Y NOR2X1_LOC_654/A 0.59fF
C61166 NAND2X1_LOC_35/Y INVX1_LOC_165/A 0.06fF
C61167 NOR2X1_LOC_262/a_36_216# INVX1_LOC_57/A 0.00fF
C61168 INVX1_LOC_31/A NOR2X1_LOC_662/A 0.07fF
C61169 INVX1_LOC_235/Y INVX1_LOC_32/A 0.08fF
C61170 INVX1_LOC_34/A NOR2X1_LOC_331/B 0.09fF
C61171 INVX1_LOC_214/A NOR2X1_LOC_681/Y 0.09fF
C61172 INVX1_LOC_225/A NOR2X1_LOC_536/A 0.16fF
C61173 INVX1_LOC_144/Y VDD 0.13fF
C61174 NAND2X1_LOC_149/Y INVX1_LOC_32/A 0.09fF
C61175 INVX1_LOC_5/A INVX1_LOC_78/A 0.11fF
C61176 INVX1_LOC_214/A INVX1_LOC_37/A 0.06fF
C61177 NOR2X1_LOC_216/Y INVX1_LOC_73/A 1.35fF
C61178 INVX1_LOC_232/A INVX1_LOC_74/A 0.02fF
C61179 INVX1_LOC_157/A NOR2X1_LOC_78/A 0.01fF
C61180 INVX1_LOC_263/A NAND2X1_LOC_454/a_36_24# 0.00fF
C61181 NOR2X1_LOC_667/A INVX1_LOC_37/A 3.29fF
C61182 INVX1_LOC_57/A INVX1_LOC_23/A 0.47fF
C61183 NOR2X1_LOC_320/Y INVX1_LOC_28/A 0.01fF
C61184 INVX1_LOC_41/A NAND2X1_LOC_698/a_36_24# 0.00fF
C61185 INVX1_LOC_248/A INVX1_LOC_37/A 0.07fF
C61186 NOR2X1_LOC_456/Y INVX1_LOC_50/A 0.07fF
C61187 NOR2X1_LOC_624/A NAND2X1_LOC_617/a_36_24# 0.00fF
C61188 NOR2X1_LOC_598/B NOR2X1_LOC_383/B 0.22fF
C61189 INVX1_LOC_93/A NAND2X1_LOC_443/a_36_24# 0.01fF
C61190 INPUT_0 INVX1_LOC_102/Y 0.05fF
C61191 NAND2X1_LOC_866/B NOR2X1_LOC_526/a_36_216# 0.00fF
C61192 INVX1_LOC_77/A INVX1_LOC_46/Y 0.03fF
C61193 NOR2X1_LOC_272/Y INVX1_LOC_94/Y 0.01fF
C61194 NOR2X1_LOC_514/A NAND2X1_LOC_82/Y 0.04fF
C61195 INVX1_LOC_162/Y INVX1_LOC_118/A 0.02fF
C61196 NOR2X1_LOC_357/Y INVX1_LOC_16/A 0.10fF
C61197 INVX1_LOC_13/A NOR2X1_LOC_35/Y 0.10fF
C61198 INVX1_LOC_21/A NAND2X1_LOC_72/B 0.05fF
C61199 NAND2X1_LOC_850/A INVX1_LOC_6/A 0.15fF
C61200 INVX1_LOC_178/A INVX1_LOC_78/A 0.06fF
C61201 NOR2X1_LOC_816/A INVX1_LOC_42/A 0.03fF
C61202 INVX1_LOC_33/A INVX1_LOC_92/A 0.21fF
C61203 INVX1_LOC_15/Y INVX1_LOC_280/A 0.03fF
C61204 NAND2X1_LOC_711/Y INVX1_LOC_12/A 0.01fF
C61205 NAND2X1_LOC_182/A INVX1_LOC_54/A 0.03fF
C61206 INVX1_LOC_104/A INVX1_LOC_54/A 0.07fF
C61207 INVX1_LOC_30/A INVX1_LOC_125/A 0.00fF
C61208 NOR2X1_LOC_315/Y INVX1_LOC_127/A 0.03fF
C61209 NAND2X1_LOC_711/Y NOR2X1_LOC_519/Y 0.04fF
C61210 INVX1_LOC_90/A NOR2X1_LOC_311/Y 0.01fF
C61211 INVX1_LOC_72/A INVX1_LOC_19/A 0.10fF
C61212 NAND2X1_LOC_231/Y NOR2X1_LOC_331/B 0.10fF
C61213 INVX1_LOC_225/A NAND2X1_LOC_93/B 0.07fF
C61214 INVX1_LOC_166/A NOR2X1_LOC_663/A 0.01fF
C61215 NOR2X1_LOC_78/B INVX1_LOC_38/A 0.14fF
C61216 INVX1_LOC_1/Y INVX1_LOC_12/Y 0.18fF
C61217 INVX1_LOC_72/A NOR2X1_LOC_11/Y 0.26fF
C61218 INVX1_LOC_36/A NAND2X1_LOC_207/B 0.00fF
C61219 NAND2X1_LOC_738/B NAND2X1_LOC_725/A 0.43fF
C61220 INVX1_LOC_89/A NOR2X1_LOC_799/B 0.02fF
C61221 NOR2X1_LOC_74/A NOR2X1_LOC_167/Y 0.02fF
C61222 NOR2X1_LOC_742/A NOR2X1_LOC_741/A 0.17fF
C61223 INVX1_LOC_198/Y INVX1_LOC_19/A 0.05fF
C61224 INVX1_LOC_155/A NOR2X1_LOC_117/Y 0.01fF
C61225 INVX1_LOC_64/A NOR2X1_LOC_717/A 0.07fF
C61226 NAND2X1_LOC_555/Y NAND2X1_LOC_223/a_36_24# 0.01fF
C61227 INVX1_LOC_90/A NOR2X1_LOC_164/Y 0.02fF
C61228 INVX1_LOC_16/A NOR2X1_LOC_692/Y 0.01fF
C61229 NOR2X1_LOC_843/B NAND2X1_LOC_473/A 0.08fF
C61230 D_INPUT_0 NOR2X1_LOC_138/a_36_216# 0.00fF
C61231 NOR2X1_LOC_516/B NOR2X1_LOC_865/A 0.28fF
C61232 INVX1_LOC_269/A INVX1_LOC_175/A 0.00fF
C61233 NOR2X1_LOC_214/B INVX1_LOC_139/A 0.10fF
C61234 NAND2X1_LOC_149/Y INVX1_LOC_262/A 0.06fF
C61235 NOR2X1_LOC_667/A NOR2X1_LOC_743/Y 0.06fF
C61236 INVX1_LOC_89/A INVX1_LOC_178/Y 0.03fF
C61237 NOR2X1_LOC_175/A NAND2X1_LOC_255/a_36_24# 0.01fF
C61238 NAND2X1_LOC_569/B NAND2X1_LOC_565/a_36_24# 0.03fF
C61239 INVX1_LOC_230/Y INVX1_LOC_4/Y 0.01fF
C61240 NAND2X1_LOC_337/B INVX1_LOC_78/A 0.11fF
C61241 INVX1_LOC_248/A NOR2X1_LOC_743/Y 0.03fF
C61242 INVX1_LOC_48/Y NOR2X1_LOC_646/B 0.15fF
C61243 NOR2X1_LOC_516/B NOR2X1_LOC_656/Y 0.01fF
C61244 NAND2X1_LOC_350/B NOR2X1_LOC_435/A 0.00fF
C61245 NOR2X1_LOC_816/A INVX1_LOC_78/A 0.03fF
C61246 INVX1_LOC_90/A INVX1_LOC_46/A 0.15fF
C61247 NOR2X1_LOC_473/B VDD 0.58fF
C61248 NOR2X1_LOC_45/Y NAND2X1_LOC_470/B 0.07fF
C61249 INVX1_LOC_269/A NOR2X1_LOC_19/a_36_216# 0.00fF
C61250 NOR2X1_LOC_443/Y INVX1_LOC_1/A 0.01fF
C61251 NOR2X1_LOC_389/B INVX1_LOC_46/A 0.07fF
C61252 NOR2X1_LOC_658/Y INVX1_LOC_4/A 0.01fF
C61253 INVX1_LOC_225/A NOR2X1_LOC_661/A 0.67fF
C61254 NOR2X1_LOC_178/Y INVX1_LOC_306/Y 0.10fF
C61255 NOR2X1_LOC_27/Y INVX1_LOC_5/Y 0.00fF
C61256 INVX1_LOC_25/A NAND2X1_LOC_347/B 0.09fF
C61257 INVX1_LOC_23/A NOR2X1_LOC_475/A 0.01fF
C61258 INVX1_LOC_126/Y NAND2X1_LOC_642/Y 0.01fF
C61259 NAND2X1_LOC_361/Y NAND2X1_LOC_74/B 0.10fF
C61260 INVX1_LOC_83/A INVX1_LOC_38/A 0.75fF
C61261 NOR2X1_LOC_544/A NAND2X1_LOC_438/a_36_24# 0.00fF
C61262 NOR2X1_LOC_333/a_36_216# INVX1_LOC_117/A 0.00fF
C61263 INVX1_LOC_50/A NAND2X1_LOC_719/a_36_24# 0.00fF
C61264 INVX1_LOC_89/A INVX1_LOC_114/A 0.00fF
C61265 NAND2X1_LOC_11/Y NOR2X1_LOC_430/Y 0.01fF
C61266 NAND2X1_LOC_192/B INVX1_LOC_29/Y 0.01fF
C61267 D_INPUT_0 INVX1_LOC_9/A 0.09fF
C61268 NOR2X1_LOC_846/Y INVX1_LOC_38/Y 0.48fF
C61269 NOR2X1_LOC_290/Y NOR2X1_LOC_662/A 0.01fF
C61270 NAND2X1_LOC_114/B NOR2X1_LOC_720/A 0.02fF
C61271 NOR2X1_LOC_74/A INVX1_LOC_76/A 0.66fF
C61272 NOR2X1_LOC_322/Y VDD 1.52fF
C61273 INVX1_LOC_147/A NAND2X1_LOC_453/A 0.20fF
C61274 INVX1_LOC_5/A NOR2X1_LOC_215/A 0.04fF
C61275 NOR2X1_LOC_456/Y NAND2X1_LOC_178/a_36_24# 0.01fF
C61276 INVX1_LOC_88/A NOR2X1_LOC_678/A 0.01fF
C61277 NAND2X1_LOC_51/B INVX1_LOC_37/A 0.12fF
C61278 D_INPUT_1 INVX1_LOC_150/Y 0.07fF
C61279 NOR2X1_LOC_338/Y NOR2X1_LOC_334/Y 0.15fF
C61280 NOR2X1_LOC_316/Y NAND2X1_LOC_63/Y 0.01fF
C61281 INVX1_LOC_48/Y NOR2X1_LOC_293/a_36_216# 0.00fF
C61282 INVX1_LOC_1/A INVX1_LOC_213/A 0.11fF
C61283 INVX1_LOC_119/A INVX1_LOC_12/A 1.03fF
C61284 NOR2X1_LOC_537/Y INVX1_LOC_19/A 0.44fF
C61285 INVX1_LOC_96/A INVX1_LOC_247/A 0.02fF
C61286 NAND2X1_LOC_338/B INVX1_LOC_19/A 0.25fF
C61287 INVX1_LOC_311/A INVX1_LOC_37/A 0.68fF
C61288 INVX1_LOC_31/A INVX1_LOC_57/A 0.28fF
C61289 INVX1_LOC_92/Y VDD 0.51fF
C61290 INVX1_LOC_111/Y INVX1_LOC_29/A 0.02fF
C61291 NAND2X1_LOC_562/B INVX1_LOC_42/A 0.03fF
C61292 NAND2X1_LOC_323/B INVX1_LOC_19/A 0.03fF
C61293 NOR2X1_LOC_516/B INVX1_LOC_63/A 0.09fF
C61294 INVX1_LOC_16/A NAND2X1_LOC_489/Y 0.15fF
C61295 NAND2X1_LOC_728/Y NOR2X1_LOC_829/A 0.00fF
C61296 INVX1_LOC_89/A INVX1_LOC_307/A 0.07fF
C61297 NOR2X1_LOC_360/Y INVX1_LOC_26/A 0.09fF
C61298 NOR2X1_LOC_733/Y INVX1_LOC_139/Y 0.01fF
C61299 NOR2X1_LOC_744/Y NAND2X1_LOC_175/Y 0.05fF
C61300 INVX1_LOC_75/A NOR2X1_LOC_114/a_36_216# 0.00fF
C61301 NOR2X1_LOC_355/B VDD 0.08fF
C61302 INVX1_LOC_89/A NOR2X1_LOC_445/B 0.07fF
C61303 INVX1_LOC_155/Y NAND2X1_LOC_647/B 0.00fF
C61304 INVX1_LOC_2/A INVX1_LOC_290/Y 0.07fF
C61305 NOR2X1_LOC_180/B NOR2X1_LOC_197/B 0.10fF
C61306 INPUT_0 NOR2X1_LOC_331/B 0.07fF
C61307 NOR2X1_LOC_562/B VDD 0.50fF
C61308 INVX1_LOC_224/Y INVX1_LOC_72/Y 0.01fF
C61309 INVX1_LOC_161/Y NOR2X1_LOC_674/Y 0.03fF
C61310 INVX1_LOC_150/Y NOR2X1_LOC_108/a_36_216# 0.01fF
C61311 INVX1_LOC_256/A NOR2X1_LOC_186/Y 0.15fF
C61312 INVX1_LOC_150/Y NOR2X1_LOC_652/Y 0.13fF
C61313 NAND2X1_LOC_796/B INVX1_LOC_11/A 0.11fF
C61314 NOR2X1_LOC_773/Y INVX1_LOC_42/A 0.07fF
C61315 NOR2X1_LOC_318/B INVX1_LOC_12/Y 0.10fF
C61316 INVX1_LOC_136/A NAND2X1_LOC_571/B 0.04fF
C61317 INVX1_LOC_64/A NOR2X1_LOC_658/Y 0.26fF
C61318 INVX1_LOC_50/A NOR2X1_LOC_759/Y 0.04fF
C61319 NOR2X1_LOC_344/a_36_216# NOR2X1_LOC_334/Y 0.01fF
C61320 NAND2X1_LOC_860/A INVX1_LOC_18/A 0.07fF
C61321 NAND2X1_LOC_386/a_36_24# INVX1_LOC_53/A 0.00fF
C61322 NAND2X1_LOC_41/Y NOR2X1_LOC_340/A 0.01fF
C61323 INVX1_LOC_178/A NOR2X1_LOC_503/Y 0.08fF
C61324 NOR2X1_LOC_536/Y NAND2X1_LOC_537/Y 0.09fF
C61325 NAND2X1_LOC_549/Y NOR2X1_LOC_384/Y 0.01fF
C61326 INVX1_LOC_202/A INVX1_LOC_50/A 0.07fF
C61327 NAND2X1_LOC_112/Y NOR2X1_LOC_89/A 0.03fF
C61328 NOR2X1_LOC_210/B NAND2X1_LOC_220/B 0.35fF
C61329 NOR2X1_LOC_377/Y INVX1_LOC_78/A 0.03fF
C61330 NAND2X1_LOC_656/A INVX1_LOC_29/Y 0.01fF
C61331 NOR2X1_LOC_91/a_36_216# NAND2X1_LOC_793/B 0.01fF
C61332 INVX1_LOC_93/Y INVX1_LOC_12/Y 0.10fF
C61333 NOR2X1_LOC_218/Y INVX1_LOC_290/Y 0.19fF
C61334 NOR2X1_LOC_348/B NAND2X1_LOC_454/Y 0.01fF
C61335 INVX1_LOC_135/A INVX1_LOC_49/Y 0.01fF
C61336 INVX1_LOC_50/A NOR2X1_LOC_550/B 0.01fF
C61337 VDD NAND2X1_LOC_836/Y 0.03fF
C61338 NOR2X1_LOC_67/A NOR2X1_LOC_38/B 0.08fF
C61339 NAND2X1_LOC_537/Y NAND2X1_LOC_799/A 0.23fF
C61340 NOR2X1_LOC_311/Y INVX1_LOC_38/A 0.02fF
C61341 INVX1_LOC_269/A NOR2X1_LOC_82/A 0.17fF
C61342 INVX1_LOC_85/Y INVX1_LOC_186/Y 0.01fF
C61343 INVX1_LOC_85/A NOR2X1_LOC_631/Y 0.03fF
C61344 NOR2X1_LOC_536/A NAND2X1_LOC_642/Y 0.21fF
C61345 NOR2X1_LOC_285/A NAND2X1_LOC_361/Y 0.04fF
C61346 NAND2X1_LOC_182/A NOR2X1_LOC_438/Y 0.01fF
C61347 INVX1_LOC_150/A INVX1_LOC_12/A 0.03fF
C61348 INVX1_LOC_5/A NOR2X1_LOC_554/B 0.23fF
C61349 NOR2X1_LOC_137/A INVX1_LOC_29/A 0.13fF
C61350 INVX1_LOC_28/A NAND2X1_LOC_489/Y 0.01fF
C61351 INVX1_LOC_58/A INVX1_LOC_209/Y 0.03fF
C61352 INVX1_LOC_16/A INVX1_LOC_32/A 7.21fF
C61353 INVX1_LOC_313/Y INVX1_LOC_19/A 0.09fF
C61354 NAND2X1_LOC_807/Y NOR2X1_LOC_662/A 0.02fF
C61355 NOR2X1_LOC_332/A NOR2X1_LOC_847/A 0.03fF
C61356 INVX1_LOC_64/A NOR2X1_LOC_13/Y 0.13fF
C61357 NAND2X1_LOC_717/Y NAND2X1_LOC_175/Y 4.85fF
C61358 NOR2X1_LOC_99/B NOR2X1_LOC_67/Y 0.05fF
C61359 INVX1_LOC_89/A INVX1_LOC_12/A 7.12fF
C61360 NAND2X1_LOC_650/B NOR2X1_LOC_176/Y 0.04fF
C61361 NOR2X1_LOC_164/Y INVX1_LOC_38/A 0.33fF
C61362 NAND2X1_LOC_231/Y NOR2X1_LOC_449/A 0.01fF
C61363 NOR2X1_LOC_773/Y INVX1_LOC_78/A 0.15fF
C61364 INVX1_LOC_90/A NOR2X1_LOC_671/Y 0.05fF
C61365 INVX1_LOC_33/A INVX1_LOC_53/A 0.73fF
C61366 INVX1_LOC_225/Y NOR2X1_LOC_541/Y 0.04fF
C61367 NOR2X1_LOC_537/Y INVX1_LOC_26/Y 0.03fF
C61368 NAND2X1_LOC_338/B INVX1_LOC_26/Y 0.07fF
C61369 INVX1_LOC_58/A NOR2X1_LOC_718/B 0.08fF
C61370 VDD NOR2X1_LOC_863/Y 0.24fF
C61371 INVX1_LOC_21/A NAND2X1_LOC_198/B 0.22fF
C61372 INVX1_LOC_299/A NOR2X1_LOC_336/B 0.02fF
C61373 INVX1_LOC_5/A NOR2X1_LOC_152/Y 0.03fF
C61374 VDD INVX1_LOC_281/Y -0.00fF
C61375 INVX1_LOC_22/A NAND2X1_LOC_454/Y 0.08fF
C61376 INVX1_LOC_304/A NOR2X1_LOC_177/Y 0.08fF
C61377 NAND2X1_LOC_784/A NAND2X1_LOC_357/B 0.01fF
C61378 NOR2X1_LOC_263/a_36_216# INVX1_LOC_29/Y 0.00fF
C61379 NAND2X1_LOC_642/Y NAND2X1_LOC_93/B 0.69fF
C61380 NAND2X1_LOC_323/B INVX1_LOC_26/Y 0.03fF
C61381 NAND2X1_LOC_9/Y NOR2X1_LOC_392/B 0.01fF
C61382 INVX1_LOC_5/A NAND2X1_LOC_193/a_36_24# 0.00fF
C61383 NAND2X1_LOC_559/Y NOR2X1_LOC_517/Y 0.00fF
C61384 NAND2X1_LOC_472/Y INVX1_LOC_117/A 0.42fF
C61385 INVX1_LOC_16/A NAND2X1_LOC_175/Y 0.07fF
C61386 INVX1_LOC_63/Y NOR2X1_LOC_665/a_36_216# 0.01fF
C61387 NOR2X1_LOC_206/a_36_216# NOR2X1_LOC_759/Y 0.00fF
C61388 INVX1_LOC_38/A INVX1_LOC_46/A 5.54fF
C61389 NOR2X1_LOC_122/A INVX1_LOC_72/A 0.03fF
C61390 INVX1_LOC_53/A NAND2X1_LOC_466/A 0.02fF
C61391 INVX1_LOC_290/A NOR2X1_LOC_158/Y 0.04fF
C61392 NAND2X1_LOC_184/a_36_24# INVX1_LOC_99/A 0.02fF
C61393 NOR2X1_LOC_590/Y NOR2X1_LOC_550/B 0.01fF
C61394 INVX1_LOC_191/Y INVX1_LOC_57/A 0.03fF
C61395 NAND2X1_LOC_11/Y INVX1_LOC_296/A 0.01fF
C61396 NOR2X1_LOC_65/B NOR2X1_LOC_773/Y 0.01fF
C61397 INVX1_LOC_123/A NOR2X1_LOC_673/A 0.00fF
C61398 INVX1_LOC_48/A NOR2X1_LOC_673/B 0.03fF
C61399 NOR2X1_LOC_486/Y INVX1_LOC_92/A 0.01fF
C61400 INVX1_LOC_299/A NAND2X1_LOC_364/A 0.12fF
C61401 NOR2X1_LOC_250/A INVX1_LOC_30/A 0.03fF
C61402 NAND2X1_LOC_537/Y INVX1_LOC_18/A 0.07fF
C61403 INVX1_LOC_6/A NOR2X1_LOC_662/A 0.01fF
C61404 INVX1_LOC_178/A NOR2X1_LOC_152/Y 0.10fF
C61405 INVX1_LOC_140/A INVX1_LOC_42/A 0.10fF
C61406 NAND2X1_LOC_317/a_36_24# INVX1_LOC_78/A 0.01fF
C61407 INVX1_LOC_45/A INVX1_LOC_225/Y 0.04fF
C61408 INVX1_LOC_35/A NOR2X1_LOC_802/A 0.04fF
C61409 NOR2X1_LOC_538/B NAND2X1_LOC_364/A 0.04fF
C61410 INVX1_LOC_22/A NOR2X1_LOC_831/a_36_216# 0.02fF
C61411 NAND2X1_LOC_363/B NOR2X1_LOC_709/A 0.14fF
C61412 D_INPUT_7 NOR2X1_LOC_408/a_36_216# 0.00fF
C61413 INVX1_LOC_225/Y NOR2X1_LOC_568/A 0.25fF
C61414 INVX1_LOC_161/Y INVX1_LOC_72/A 0.07fF
C61415 INVX1_LOC_315/Y INVX1_LOC_63/A 0.16fF
C61416 NOR2X1_LOC_242/A INVX1_LOC_33/A 1.20fF
C61417 INVX1_LOC_83/A NAND2X1_LOC_223/A 0.07fF
C61418 INVX1_LOC_28/A INVX1_LOC_32/A 0.22fF
C61419 NOR2X1_LOC_454/Y INVX1_LOC_49/A 0.07fF
C61420 NAND2X1_LOC_463/B INVX1_LOC_42/A 0.00fF
C61421 NOR2X1_LOC_361/B NAND2X1_LOC_515/a_36_24# 0.06fF
C61422 NAND2X1_LOC_637/Y INVX1_LOC_117/A 0.04fF
C61423 NAND2X1_LOC_642/Y INVX1_LOC_3/A -0.00fF
C61424 NOR2X1_LOC_570/A NOR2X1_LOC_383/B 0.01fF
C61425 INVX1_LOC_48/A INVX1_LOC_29/A 0.06fF
C61426 NOR2X1_LOC_180/Y INVX1_LOC_50/Y 0.12fF
C61427 NOR2X1_LOC_84/Y NOR2X1_LOC_293/a_36_216# 0.02fF
C61428 NAND2X1_LOC_859/Y INVX1_LOC_57/A 0.03fF
C61429 NOR2X1_LOC_208/Y NOR2X1_LOC_217/a_36_216# 0.00fF
C61430 INVX1_LOC_5/A NOR2X1_LOC_721/A 0.06fF
C61431 NOR2X1_LOC_272/Y NOR2X1_LOC_315/Y 0.10fF
C61432 INPUT_5 INVX1_LOC_296/Y 0.01fF
C61433 NOR2X1_LOC_441/Y INVX1_LOC_177/Y 0.65fF
C61434 NAND2X1_LOC_30/Y INVX1_LOC_77/A 0.32fF
C61435 INVX1_LOC_225/Y INVX1_LOC_71/A 0.06fF
C61436 INVX1_LOC_72/A NOR2X1_LOC_599/A 0.02fF
C61437 INVX1_LOC_28/A NAND2X1_LOC_175/Y 0.15fF
C61438 NOR2X1_LOC_816/A NOR2X1_LOC_152/Y 0.08fF
C61439 INVX1_LOC_132/A INVX1_LOC_256/A 0.03fF
C61440 INVX1_LOC_14/A INVX1_LOC_8/A 0.17fF
C61441 INVX1_LOC_305/A NOR2X1_LOC_500/B 0.10fF
C61442 NOR2X1_LOC_78/A NOR2X1_LOC_89/A 0.80fF
C61443 NOR2X1_LOC_510/Y INVX1_LOC_144/Y 0.01fF
C61444 INVX1_LOC_21/A NAND2X1_LOC_491/a_36_24# 0.00fF
C61445 INVX1_LOC_140/A INVX1_LOC_78/A 1.50fF
C61446 NAND2X1_LOC_93/B NOR2X1_LOC_271/Y 0.03fF
C61447 INVX1_LOC_250/A INVX1_LOC_136/A 0.01fF
C61448 NOR2X1_LOC_242/A INVX1_LOC_120/Y 0.01fF
C61449 NOR2X1_LOC_552/A INVX1_LOC_99/A 0.01fF
C61450 INVX1_LOC_5/A NAND2X1_LOC_859/B 0.02fF
C61451 INVX1_LOC_46/Y INVX1_LOC_9/A 0.12fF
C61452 INVX1_LOC_223/Y NOR2X1_LOC_500/Y 0.02fF
C61453 NOR2X1_LOC_369/Y NAND2X1_LOC_833/Y 0.01fF
C61454 INVX1_LOC_251/Y NOR2X1_LOC_15/Y 3.27fF
C61455 INVX1_LOC_256/A INVX1_LOC_225/A 0.20fF
C61456 NAND2X1_LOC_387/a_36_24# INVX1_LOC_49/A 0.00fF
C61457 NAND2X1_LOC_582/a_36_24# INVX1_LOC_11/A 0.00fF
C61458 INVX1_LOC_136/A INVX1_LOC_116/A 0.06fF
C61459 INVX1_LOC_21/A INVX1_LOC_53/Y 0.08fF
C61460 INVX1_LOC_16/A INVX1_LOC_171/Y 0.02fF
C61461 INVX1_LOC_25/Y NAND2X1_LOC_474/Y 0.08fF
C61462 INVX1_LOC_21/A NOR2X1_LOC_619/A 0.03fF
C61463 NOR2X1_LOC_437/Y INVX1_LOC_72/A 0.07fF
C61464 NAND2X1_LOC_807/Y INVX1_LOC_57/A 1.02fF
C61465 NAND2X1_LOC_357/B NAND2X1_LOC_807/A 0.04fF
C61466 NAND2X1_LOC_9/Y INVX1_LOC_90/A 0.07fF
C61467 NOR2X1_LOC_602/A NAND2X1_LOC_601/a_36_24# 0.02fF
C61468 NOR2X1_LOC_186/Y NOR2X1_LOC_440/Y 0.01fF
C61469 NOR2X1_LOC_89/A NAND2X1_LOC_464/A 0.10fF
C61470 INVX1_LOC_3/A NOR2X1_LOC_271/Y 0.12fF
C61471 NOR2X1_LOC_454/Y NOR2X1_LOC_161/Y 0.12fF
C61472 VDD INVX1_LOC_106/A 0.12fF
C61473 NAND2X1_LOC_35/Y NOR2X1_LOC_71/Y 0.02fF
C61474 NOR2X1_LOC_488/Y NAND2X1_LOC_579/A 0.01fF
C61475 INVX1_LOC_233/A INVX1_LOC_90/A 0.07fF
C61476 INVX1_LOC_45/Y INVX1_LOC_94/A 0.05fF
C61477 NOR2X1_LOC_455/Y NOR2X1_LOC_356/A 0.01fF
C61478 INVX1_LOC_36/A INVX1_LOC_155/A 0.04fF
C61479 NOR2X1_LOC_155/A INVX1_LOC_179/A 0.38fF
C61480 NAND2X1_LOC_552/A NAND2X1_LOC_861/Y 0.01fF
C61481 INVX1_LOC_136/A NAND2X1_LOC_361/Y 0.06fF
C61482 NOR2X1_LOC_441/Y INVX1_LOC_104/A 0.02fF
C61483 NOR2X1_LOC_68/A NOR2X1_LOC_577/Y 0.07fF
C61484 NAND2X1_LOC_149/Y GATE_662 0.04fF
C61485 NOR2X1_LOC_152/A INVX1_LOC_49/Y 0.49fF
C61486 INVX1_LOC_13/A INVX1_LOC_48/Y 0.07fF
C61487 INVX1_LOC_11/A NAND2X1_LOC_541/Y 0.01fF
C61488 INVX1_LOC_35/A NOR2X1_LOC_174/A 0.03fF
C61489 INVX1_LOC_215/A NOR2X1_LOC_92/Y 0.07fF
C61490 NOR2X1_LOC_446/A NOR2X1_LOC_778/B 0.01fF
C61491 NAND2X1_LOC_856/A NAND2X1_LOC_811/Y 0.03fF
C61492 NOR2X1_LOC_82/A NAND2X1_LOC_563/A 0.57fF
C61493 INVX1_LOC_35/A NOR2X1_LOC_111/Y 0.06fF
C61494 NOR2X1_LOC_598/B NOR2X1_LOC_163/Y 0.07fF
C61495 INVX1_LOC_105/A NOR2X1_LOC_759/Y 0.04fF
C61496 NOR2X1_LOC_405/A INVX1_LOC_94/Y 0.03fF
C61497 NOR2X1_LOC_332/A NOR2X1_LOC_655/a_36_216# 0.01fF
C61498 NOR2X1_LOC_454/Y NOR2X1_LOC_781/a_36_216# 0.01fF
C61499 INVX1_LOC_315/Y NAND2X1_LOC_223/B 0.20fF
C61500 INVX1_LOC_91/A NOR2X1_LOC_278/Y 0.02fF
C61501 NAND2X1_LOC_364/A INVX1_LOC_162/A 0.05fF
C61502 NOR2X1_LOC_520/B INVX1_LOC_62/Y 0.04fF
C61503 INVX1_LOC_35/A INVX1_LOC_82/Y 0.01fF
C61504 NOR2X1_LOC_323/Y INVX1_LOC_53/A 0.00fF
C61505 NOR2X1_LOC_296/Y INVX1_LOC_16/A 0.07fF
C61506 INVX1_LOC_45/A INVX1_LOC_266/Y 0.08fF
C61507 INVX1_LOC_178/A NAND2X1_LOC_861/Y 0.23fF
C61508 NOR2X1_LOC_798/A INVX1_LOC_90/A 0.03fF
C61509 INVX1_LOC_30/A NOR2X1_LOC_709/A 0.17fF
C61510 NOR2X1_LOC_598/B NOR2X1_LOC_74/Y 0.02fF
C61511 INVX1_LOC_6/A INVX1_LOC_57/A 0.13fF
C61512 NOR2X1_LOC_92/Y NOR2X1_LOC_373/Y 0.02fF
C61513 NOR2X1_LOC_859/Y NOR2X1_LOC_861/Y 0.00fF
C61514 NOR2X1_LOC_215/Y NOR2X1_LOC_142/Y 0.02fF
C61515 NAND2X1_LOC_53/Y NOR2X1_LOC_302/B 0.03fF
C61516 INVX1_LOC_49/A INVX1_LOC_77/A 0.15fF
C61517 NOR2X1_LOC_455/Y NOR2X1_LOC_74/A 0.04fF
C61518 NOR2X1_LOC_798/A NOR2X1_LOC_389/B 0.01fF
C61519 D_GATE_741 INVX1_LOC_174/Y 0.02fF
C61520 INVX1_LOC_36/A NAND2X1_LOC_661/B 0.01fF
C61521 INVX1_LOC_280/A NOR2X1_LOC_672/a_36_216# 0.01fF
C61522 NOR2X1_LOC_96/Y NOR2X1_LOC_671/Y 0.01fF
C61523 NOR2X1_LOC_160/B INVX1_LOC_1/Y 0.15fF
C61524 INVX1_LOC_90/A NAND2X1_LOC_703/Y 0.46fF
C61525 NOR2X1_LOC_590/A INVX1_LOC_208/Y 0.68fF
C61526 INVX1_LOC_310/A NAND2X1_LOC_364/A 0.00fF
C61527 NAND2X1_LOC_656/A INVX1_LOC_60/Y 0.12fF
C61528 NAND2X1_LOC_569/A NOR2X1_LOC_237/Y -0.08fF
C61529 NOR2X1_LOC_122/A INVX1_LOC_313/Y 0.00fF
C61530 INVX1_LOC_5/A INVX1_LOC_158/Y 0.09fF
C61531 NOR2X1_LOC_68/A NOR2X1_LOC_346/B 0.03fF
C61532 VDD NOR2X1_LOC_464/Y 0.31fF
C61533 INVX1_LOC_71/A INVX1_LOC_266/Y 0.07fF
C61534 NOR2X1_LOC_275/a_36_216# NOR2X1_LOC_561/Y 0.01fF
C61535 INVX1_LOC_36/A NOR2X1_LOC_229/Y 0.05fF
C61536 INVX1_LOC_157/A NOR2X1_LOC_45/Y 0.06fF
C61537 INVX1_LOC_75/A NAND2X1_LOC_474/Y 0.07fF
C61538 NOR2X1_LOC_483/B INVX1_LOC_83/A 0.01fF
C61539 INVX1_LOC_124/A INVX1_LOC_49/A 0.47fF
C61540 INVX1_LOC_2/A INVX1_LOC_77/A 0.15fF
C61541 NOR2X1_LOC_791/B NOR2X1_LOC_121/A 0.23fF
C61542 NOR2X1_LOC_346/Y NOR2X1_LOC_416/A 0.02fF
C61543 NAND2X1_LOC_167/a_36_24# NOR2X1_LOC_500/Y 0.01fF
C61544 NOR2X1_LOC_68/A INVX1_LOC_22/A 0.22fF
C61545 NOR2X1_LOC_142/Y INVX1_LOC_104/A 0.10fF
C61546 INVX1_LOC_161/Y INVX1_LOC_313/Y 0.10fF
C61547 NAND2X1_LOC_338/B NAND2X1_LOC_119/a_36_24# 0.01fF
C61548 NOR2X1_LOC_226/A INVX1_LOC_77/A 0.00fF
C61549 INVX1_LOC_135/A NAND2X1_LOC_208/B 0.21fF
C61550 NOR2X1_LOC_861/Y INVX1_LOC_46/Y 0.02fF
C61551 INVX1_LOC_216/Y NOR2X1_LOC_19/B 0.02fF
C61552 NOR2X1_LOC_770/Y INVX1_LOC_174/A -0.03fF
C61553 NOR2X1_LOC_620/Y INVX1_LOC_143/A 0.03fF
C61554 NOR2X1_LOC_773/Y NOR2X1_LOC_152/Y 0.01fF
C61555 NOR2X1_LOC_781/A INVX1_LOC_159/A 0.40fF
C61556 INVX1_LOC_33/A NOR2X1_LOC_547/B 0.01fF
C61557 NOR2X1_LOC_78/B INVX1_LOC_33/A 0.42fF
C61558 INVX1_LOC_314/Y INVX1_LOC_232/A 0.10fF
C61559 NOR2X1_LOC_243/B NAND2X1_LOC_202/a_36_24# 0.00fF
C61560 NOR2X1_LOC_794/B NOR2X1_LOC_564/Y 0.37fF
C61561 NAND2X1_LOC_207/B INVX1_LOC_63/A 0.00fF
C61562 NOR2X1_LOC_78/B NOR2X1_LOC_743/a_36_216# 0.01fF
C61563 NOR2X1_LOC_503/Y INVX1_LOC_140/A 0.10fF
C61564 NAND2X1_LOC_778/Y NOR2X1_LOC_45/B 0.10fF
C61565 NAND2X1_LOC_53/Y INVX1_LOC_75/A 0.10fF
C61566 INVX1_LOC_11/A NAND2X1_LOC_840/Y 0.02fF
C61567 NOR2X1_LOC_332/A NOR2X1_LOC_554/B 0.02fF
C61568 INVX1_LOC_77/A NOR2X1_LOC_161/Y 0.07fF
C61569 NOR2X1_LOC_92/Y INVX1_LOC_286/A 0.07fF
C61570 NOR2X1_LOC_848/Y INPUT_0 0.00fF
C61571 NOR2X1_LOC_216/B INVX1_LOC_47/Y 0.43fF
C61572 NAND2X1_LOC_217/a_36_24# INVX1_LOC_13/A 0.00fF
C61573 NOR2X1_LOC_304/a_36_216# NOR2X1_LOC_56/Y 0.00fF
C61574 NAND2X1_LOC_364/A INVX1_LOC_66/A 0.01fF
C61575 INVX1_LOC_17/A NOR2X1_LOC_335/B 0.17fF
C61576 INVX1_LOC_49/A NOR2X1_LOC_687/Y 0.20fF
C61577 NOR2X1_LOC_655/B INVX1_LOC_104/A 0.12fF
C61578 NAND2X1_LOC_112/Y NOR2X1_LOC_433/A 0.02fF
C61579 NOR2X1_LOC_383/Y INVX1_LOC_314/Y 0.03fF
C61580 INVX1_LOC_13/A NOR2X1_LOC_350/A 0.01fF
C61581 NOR2X1_LOC_570/Y NOR2X1_LOC_577/Y 0.01fF
C61582 INVX1_LOC_58/A NAND2X1_LOC_472/Y 0.10fF
C61583 INVX1_LOC_217/A INVX1_LOC_89/A 0.04fF
C61584 INVX1_LOC_18/A INVX1_LOC_85/Y 0.71fF
C61585 NOR2X1_LOC_15/Y NOR2X1_LOC_555/a_36_216# 0.02fF
C61586 INVX1_LOC_36/A NAND2X1_LOC_850/A 0.03fF
C61587 NOR2X1_LOC_15/Y NOR2X1_LOC_45/B 0.13fF
C61588 INVX1_LOC_34/A NAND2X1_LOC_479/Y 0.14fF
C61589 NOR2X1_LOC_78/B NOR2X1_LOC_714/Y 0.01fF
C61590 NOR2X1_LOC_121/Y NOR2X1_LOC_719/A 0.01fF
C61591 NOR2X1_LOC_632/Y INVX1_LOC_63/Y 0.03fF
C61592 INVX1_LOC_136/A NAND2X1_LOC_654/B 0.00fF
C61593 INVX1_LOC_305/Y NOR2X1_LOC_802/A 0.02fF
C61594 NAND2X1_LOC_562/B NAND2X1_LOC_859/B 0.02fF
C61595 NOR2X1_LOC_267/A NAND2X1_LOC_850/A 0.02fF
C61596 NOR2X1_LOC_92/Y INVX1_LOC_95/A 0.03fF
C61597 INVX1_LOC_299/A NOR2X1_LOC_405/A 0.13fF
C61598 INVX1_LOC_11/A INVX1_LOC_98/A 0.77fF
C61599 NOR2X1_LOC_78/B INVX1_LOC_120/Y 0.11fF
C61600 NAND2X1_LOC_549/a_36_24# INVX1_LOC_234/A 0.00fF
C61601 INVX1_LOC_3/Y NAND2X1_LOC_773/B 0.20fF
C61602 NAND2X1_LOC_55/a_36_24# NOR2X1_LOC_391/A 0.01fF
C61603 NAND2X1_LOC_9/Y INVX1_LOC_38/A 0.07fF
C61604 NAND2X1_LOC_112/Y NOR2X1_LOC_52/B 0.03fF
C61605 NOR2X1_LOC_846/Y VDD 0.16fF
C61606 INVX1_LOC_225/A NOR2X1_LOC_440/Y 0.06fF
C61607 INVX1_LOC_83/A INVX1_LOC_33/A 0.18fF
C61608 INVX1_LOC_11/A NOR2X1_LOC_78/A 6.26fF
C61609 NOR2X1_LOC_635/B INVX1_LOC_92/A 0.06fF
C61610 INVX1_LOC_69/A NOR2X1_LOC_640/B 0.26fF
C61611 NOR2X1_LOC_334/Y NAND2X1_LOC_475/Y 0.10fF
C61612 NOR2X1_LOC_78/B INVX1_LOC_40/A 0.07fF
C61613 NOR2X1_LOC_15/Y INVX1_LOC_247/A 0.03fF
C61614 NOR2X1_LOC_155/A NAND2X1_LOC_288/B 0.03fF
C61615 NOR2X1_LOC_241/a_36_216# INVX1_LOC_37/A 0.00fF
C61616 INVX1_LOC_233/A INVX1_LOC_38/A 0.16fF
C61617 INVX1_LOC_274/A INVX1_LOC_23/A 0.08fF
C61618 INVX1_LOC_284/Y INVX1_LOC_309/A 0.00fF
C61619 NOR2X1_LOC_742/A NOR2X1_LOC_733/a_36_216# 0.01fF
C61620 INVX1_LOC_275/Y INVX1_LOC_92/A 0.01fF
C61621 NOR2X1_LOC_351/Y INVX1_LOC_53/A 0.00fF
C61622 INVX1_LOC_34/A INVX1_LOC_135/A 0.11fF
C61623 NOR2X1_LOC_383/B NOR2X1_LOC_634/A 0.02fF
C61624 NOR2X1_LOC_590/A NOR2X1_LOC_501/B 0.02fF
C61625 INVX1_LOC_269/A INVX1_LOC_59/Y 0.24fF
C61626 NOR2X1_LOC_598/B NOR2X1_LOC_332/Y 0.01fF
C61627 NAND2X1_LOC_454/Y NAND2X1_LOC_476/Y 0.03fF
C61628 NOR2X1_LOC_454/Y NOR2X1_LOC_586/Y 0.04fF
C61629 NOR2X1_LOC_160/B NOR2X1_LOC_318/B 0.07fF
C61630 INVX1_LOC_256/A NAND2X1_LOC_642/Y 0.02fF
C61631 INVX1_LOC_32/A INVX1_LOC_109/A 0.80fF
C61632 INVX1_LOC_289/A NOR2X1_LOC_418/Y 0.25fF
C61633 INVX1_LOC_236/Y INVX1_LOC_91/A 0.04fF
C61634 NAND2X1_LOC_477/Y NOR2X1_LOC_693/a_36_216# 0.00fF
C61635 NOR2X1_LOC_234/Y NOR2X1_LOC_71/Y -0.00fF
C61636 INVX1_LOC_140/A NOR2X1_LOC_152/Y 0.10fF
C61637 INVX1_LOC_2/A NAND2X1_LOC_796/Y 0.03fF
C61638 NOR2X1_LOC_160/B INVX1_LOC_93/Y 0.08fF
C61639 INVX1_LOC_226/Y INVX1_LOC_25/Y 0.04fF
C61640 INVX1_LOC_142/A INVX1_LOC_78/Y 0.02fF
C61641 NOR2X1_LOC_798/A INVX1_LOC_38/A 0.03fF
C61642 NAND2X1_LOC_355/a_36_24# NOR2X1_LOC_45/B 0.00fF
C61643 NOR2X1_LOC_67/a_36_216# NOR2X1_LOC_38/B 0.02fF
C61644 INVX1_LOC_64/A NOR2X1_LOC_640/Y 0.07fF
C61645 NOR2X1_LOC_538/B NOR2X1_LOC_857/A 0.01fF
C61646 NOR2X1_LOC_576/B NAND2X1_LOC_839/Y 0.28fF
C61647 NOR2X1_LOC_328/Y NOR2X1_LOC_695/Y 0.02fF
C61648 NOR2X1_LOC_551/B NOR2X1_LOC_703/A 0.01fF
C61649 NAND2X1_LOC_35/Y NAND2X1_LOC_243/Y 0.09fF
C61650 INVX1_LOC_34/A NOR2X1_LOC_490/Y 0.01fF
C61651 NOR2X1_LOC_274/Y NOR2X1_LOC_74/A 0.01fF
C61652 INVX1_LOC_284/Y INVX1_LOC_11/Y 0.03fF
C61653 NAND2X1_LOC_363/B NAND2X1_LOC_413/a_36_24# 0.00fF
C61654 NOR2X1_LOC_617/Y NAND2X1_LOC_622/B 0.04fF
C61655 NOR2X1_LOC_846/Y NOR2X1_LOC_846/a_36_216# 0.00fF
C61656 NOR2X1_LOC_612/Y NOR2X1_LOC_652/Y 0.04fF
C61657 D_INPUT_1 NOR2X1_LOC_673/A 0.03fF
C61658 INVX1_LOC_34/A NOR2X1_LOC_202/Y 0.02fF
C61659 NAND2X1_LOC_181/Y NOR2X1_LOC_130/A 0.03fF
C61660 NAND2X1_LOC_149/Y NOR2X1_LOC_261/A 0.04fF
C61661 NOR2X1_LOC_160/B INVX1_LOC_139/A 0.03fF
C61662 INVX1_LOC_287/A NAND2X1_LOC_782/B 0.10fF
C61663 INPUT_2 D_INPUT_3 0.19fF
C61664 INVX1_LOC_83/A INVX1_LOC_40/A 0.01fF
C61665 INVX1_LOC_78/A INVX1_LOC_42/A 0.53fF
C61666 NOR2X1_LOC_276/B NOR2X1_LOC_269/Y 0.09fF
C61667 NOR2X1_LOC_82/A INVX1_LOC_12/Y 0.02fF
C61668 NOR2X1_LOC_454/Y INVX1_LOC_118/A 0.07fF
C61669 INVX1_LOC_174/A INVX1_LOC_37/A 0.12fF
C61670 NAND2X1_LOC_550/A NAND2X1_LOC_721/A 0.07fF
C61671 NOR2X1_LOC_71/Y INVX1_LOC_56/A 0.02fF
C61672 NOR2X1_LOC_561/Y NAND2X1_LOC_660/Y 0.07fF
C61673 INVX1_LOC_64/A NOR2X1_LOC_697/Y 0.05fF
C61674 INVX1_LOC_224/Y INVX1_LOC_19/A 0.09fF
C61675 INVX1_LOC_58/A NAND2X1_LOC_773/B 0.02fF
C61676 INVX1_LOC_178/A INVX1_LOC_291/A 0.10fF
C61677 INVX1_LOC_124/Y INVX1_LOC_76/A 0.10fF
C61678 NOR2X1_LOC_481/A INVX1_LOC_69/Y 0.02fF
C61679 D_INPUT_0 NOR2X1_LOC_719/A 0.00fF
C61680 NOR2X1_LOC_92/Y INVX1_LOC_54/A 0.15fF
C61681 NOR2X1_LOC_383/B INVX1_LOC_29/A 4.91fF
C61682 INVX1_LOC_24/A NAND2X1_LOC_623/B 0.03fF
C61683 INVX1_LOC_50/A NAND2X1_LOC_74/B 0.03fF
C61684 INVX1_LOC_34/A NOR2X1_LOC_391/B 0.04fF
C61685 INVX1_LOC_223/Y NOR2X1_LOC_445/B 0.00fF
C61686 NOR2X1_LOC_468/Y NAND2X1_LOC_268/a_36_24# 0.00fF
C61687 NAND2X1_LOC_198/B INVX1_LOC_304/A 0.00fF
C61688 INVX1_LOC_41/A INVX1_LOC_286/A 0.05fF
C61689 NAND2X1_LOC_731/Y INVX1_LOC_11/Y 0.00fF
C61690 NAND2X1_LOC_357/B NOR2X1_LOC_527/Y 0.03fF
C61691 NOR2X1_LOC_65/B INVX1_LOC_42/A 1.77fF
C61692 NOR2X1_LOC_433/A NOR2X1_LOC_78/A 0.07fF
C61693 NOR2X1_LOC_213/a_36_216# NOR2X1_LOC_742/A 0.01fF
C61694 INVX1_LOC_219/A INVX1_LOC_234/A 0.01fF
C61695 INVX1_LOC_223/A INVX1_LOC_14/Y 0.01fF
C61696 NOR2X1_LOC_301/A INVX1_LOC_15/A 0.03fF
C61697 D_INPUT_0 INVX1_LOC_7/A 0.12fF
C61698 NOR2X1_LOC_669/Y INVX1_LOC_92/A 0.42fF
C61699 NAND2X1_LOC_208/B NOR2X1_LOC_813/Y 0.01fF
C61700 NOR2X1_LOC_479/B NOR2X1_LOC_19/B 0.01fF
C61701 NOR2X1_LOC_722/Y INVX1_LOC_139/Y 0.01fF
C61702 NOR2X1_LOC_253/a_36_216# INVX1_LOC_42/A 0.00fF
C61703 NAND2X1_LOC_564/B INVX1_LOC_28/A 0.04fF
C61704 INVX1_LOC_314/Y NAND2X1_LOC_447/Y 0.02fF
C61705 INVX1_LOC_286/A NAND2X1_LOC_477/A 0.10fF
C61706 NOR2X1_LOC_392/Y INVX1_LOC_12/A 0.07fF
C61707 NOR2X1_LOC_302/B NOR2X1_LOC_302/Y 0.00fF
C61708 INVX1_LOC_75/A NOR2X1_LOC_500/Y 0.08fF
C61709 INVX1_LOC_226/Y INVX1_LOC_75/A 0.03fF
C61710 INVX1_LOC_96/A NOR2X1_LOC_180/Y 0.10fF
C61711 NOR2X1_LOC_606/Y NOR2X1_LOC_271/Y 0.00fF
C61712 INVX1_LOC_41/A INVX1_LOC_95/A 0.06fF
C61713 INVX1_LOC_239/A NOR2X1_LOC_649/B 0.02fF
C61714 NOR2X1_LOC_562/B INVX1_LOC_121/Y 0.30fF
C61715 NOR2X1_LOC_52/B NOR2X1_LOC_78/A 0.13fF
C61716 NOR2X1_LOC_355/B INVX1_LOC_177/A 0.01fF
C61717 NOR2X1_LOC_816/A INVX1_LOC_291/A 0.17fF
C61718 NOR2X1_LOC_574/A NAND2X1_LOC_655/A 0.03fF
C61719 NOR2X1_LOC_2/Y INVX1_LOC_22/A 0.03fF
C61720 INVX1_LOC_24/A INVX1_LOC_117/A 0.14fF
C61721 NOR2X1_LOC_65/B INVX1_LOC_78/A 0.08fF
C61722 NOR2X1_LOC_355/A NOR2X1_LOC_329/B 0.01fF
C61723 NOR2X1_LOC_778/B INVX1_LOC_186/A 0.03fF
C61724 NOR2X1_LOC_186/Y NOR2X1_LOC_89/A 0.28fF
C61725 INVX1_LOC_75/A INVX1_LOC_10/A 0.12fF
C61726 INVX1_LOC_90/A NAND2X1_LOC_842/B 0.02fF
C61727 NOR2X1_LOC_458/B INVX1_LOC_96/A 0.00fF
C61728 INVX1_LOC_33/A INVX1_LOC_46/A 0.13fF
C61729 NOR2X1_LOC_121/Y INVX1_LOC_76/A 0.01fF
C61730 INVX1_LOC_153/A INVX1_LOC_37/A 0.01fF
C61731 NAND2X1_LOC_833/Y VDD 0.13fF
C61732 INVX1_LOC_286/A NOR2X1_LOC_211/A 0.00fF
C61733 INVX1_LOC_17/A INVX1_LOC_84/A 0.07fF
C61734 NOR2X1_LOC_337/a_36_216# NOR2X1_LOC_35/Y 0.12fF
C61735 NAND2X1_LOC_861/Y INVX1_LOC_140/A 0.10fF
C61736 INVX1_LOC_298/Y NOR2X1_LOC_383/B 3.27fF
C61737 NOR2X1_LOC_433/A NOR2X1_LOC_60/Y 0.07fF
C61738 INVX1_LOC_31/A NAND2X1_LOC_243/a_36_24# 0.00fF
C61739 INVX1_LOC_31/A NOR2X1_LOC_820/Y 0.32fF
C61740 INVX1_LOC_208/A NOR2X1_LOC_318/B 0.03fF
C61741 NAND2X1_LOC_724/Y NOR2X1_LOC_829/A 0.03fF
C61742 NOR2X1_LOC_817/Y NAND2X1_LOC_818/a_36_24# 0.00fF
C61743 INVX1_LOC_18/A NOR2X1_LOC_487/Y 0.03fF
C61744 NAND2X1_LOC_866/B NOR2X1_LOC_380/Y 0.04fF
C61745 NOR2X1_LOC_471/Y INVX1_LOC_84/A 0.03fF
C61746 NAND2X1_LOC_573/Y NOR2X1_LOC_89/A 0.05fF
C61747 D_INPUT_1 NAND2X1_LOC_400/a_36_24# 0.00fF
C61748 INVX1_LOC_135/A INPUT_0 0.26fF
C61749 NAND2X1_LOC_195/Y INVX1_LOC_117/Y 0.02fF
C61750 NOR2X1_LOC_78/B NOR2X1_LOC_486/Y 0.03fF
C61751 NAND2X1_LOC_9/Y NAND2X1_LOC_223/A 0.03fF
C61752 INVX1_LOC_85/A INVX1_LOC_14/Y 0.06fF
C61753 NOR2X1_LOC_92/Y NAND2X1_LOC_807/B 0.18fF
C61754 INVX1_LOC_34/A NOR2X1_LOC_813/Y 0.01fF
C61755 NOR2X1_LOC_103/Y INVX1_LOC_19/A 0.25fF
C61756 D_INPUT_0 NOR2X1_LOC_167/Y 0.03fF
C61757 NOR2X1_LOC_400/B INVX1_LOC_166/A 0.00fF
C61758 INVX1_LOC_57/A INVX1_LOC_28/Y 0.11fF
C61759 NAND2X1_LOC_563/A NOR2X1_LOC_124/a_36_216# 0.02fF
C61760 INVX1_LOC_58/A NOR2X1_LOC_639/Y 0.03fF
C61761 NAND2X1_LOC_724/A NOR2X1_LOC_89/A 0.08fF
C61762 NAND2X1_LOC_182/A NOR2X1_LOC_176/Y 0.06fF
C61763 INVX1_LOC_49/A INVX1_LOC_9/A 0.06fF
C61764 INVX1_LOC_77/A INVX1_LOC_118/A 0.16fF
C61765 NOR2X1_LOC_541/Y INVX1_LOC_19/A 0.01fF
C61766 NAND2X1_LOC_563/A INVX1_LOC_59/Y 0.06fF
C61767 INVX1_LOC_259/A INVX1_LOC_37/A 0.01fF
C61768 NOR2X1_LOC_359/Y NAND2X1_LOC_93/B 0.05fF
C61769 NOR2X1_LOC_92/Y NOR2X1_LOC_48/B 1.10fF
C61770 NOR2X1_LOC_392/Y NOR2X1_LOC_29/a_36_216# 0.01fF
C61771 INVX1_LOC_57/A INVX1_LOC_270/A 0.01fF
C61772 INVX1_LOC_34/A INVX1_LOC_280/A 0.31fF
C61773 NOR2X1_LOC_829/Y NAND2X1_LOC_738/B 0.01fF
C61774 INVX1_LOC_34/A NOR2X1_LOC_94/Y 0.39fF
C61775 INVX1_LOC_25/A NOR2X1_LOC_646/B 0.01fF
C61776 INVX1_LOC_164/Y VDD 0.21fF
C61777 INVX1_LOC_30/A INVX1_LOC_294/A 0.05fF
C61778 NAND2X1_LOC_510/A NOR2X1_LOC_814/A 0.05fF
C61779 INVX1_LOC_48/Y INVX1_LOC_32/A 0.03fF
C61780 NAND2X1_LOC_863/A NAND2X1_LOC_856/a_36_24# 0.04fF
C61781 INVX1_LOC_96/Y INVX1_LOC_281/A 0.06fF
C61782 GATE_479 INVX1_LOC_115/Y 0.11fF
C61783 INVX1_LOC_40/A INVX1_LOC_46/A 0.02fF
C61784 INVX1_LOC_53/A NOR2X1_LOC_748/A 0.10fF
C61785 NOR2X1_LOC_498/Y INVX1_LOC_54/A 2.56fF
C61786 INVX1_LOC_143/A INVX1_LOC_117/A 0.68fF
C61787 INVX1_LOC_60/A INVX1_LOC_9/A 0.03fF
C61788 INVX1_LOC_40/A NOR2X1_LOC_98/A 0.05fF
C61789 NOR2X1_LOC_405/A INVX1_LOC_66/A 0.03fF
C61790 NOR2X1_LOC_599/Y INVX1_LOC_12/A 0.04fF
C61791 INVX1_LOC_45/A INVX1_LOC_19/A 0.19fF
C61792 NAND2X1_LOC_53/Y INVX1_LOC_283/A 0.01fF
C61793 NAND2X1_LOC_794/B NAND2X1_LOC_175/Y 0.02fF
C61794 INVX1_LOC_266/Y NOR2X1_LOC_331/B 0.10fF
C61795 NOR2X1_LOC_503/Y INVX1_LOC_42/A 0.00fF
C61796 NOR2X1_LOC_657/B NOR2X1_LOC_366/Y 0.02fF
C61797 INVX1_LOC_290/A NOR2X1_LOC_357/Y 0.10fF
C61798 NOR2X1_LOC_568/A INVX1_LOC_19/A 0.08fF
C61799 NOR2X1_LOC_525/Y INVX1_LOC_11/Y 0.03fF
C61800 INVX1_LOC_182/A INVX1_LOC_206/Y 0.07fF
C61801 NOR2X1_LOC_82/A NOR2X1_LOC_554/A 0.01fF
C61802 NOR2X1_LOC_91/A INVX1_LOC_306/Y 0.03fF
C61803 INVX1_LOC_35/A INVX1_LOC_29/Y 0.03fF
C61804 INVX1_LOC_17/A INVX1_LOC_15/A 0.86fF
C61805 NAND2X1_LOC_477/A INVX1_LOC_54/A 3.08fF
C61806 NOR2X1_LOC_364/Y NOR2X1_LOC_364/A 0.16fF
C61807 NOR2X1_LOC_68/A INVX1_LOC_186/Y 0.03fF
C61808 INVX1_LOC_57/A NOR2X1_LOC_109/Y 0.03fF
C61809 INVX1_LOC_2/A INVX1_LOC_9/A 0.09fF
C61810 NOR2X1_LOC_234/Y NAND2X1_LOC_243/Y 0.01fF
C61811 INVX1_LOC_16/A NAND2X1_LOC_804/Y 0.09fF
C61812 NOR2X1_LOC_589/A INVX1_LOC_37/A 0.03fF
C61813 INVX1_LOC_27/A INVX1_LOC_23/Y 0.09fF
C61814 NOR2X1_LOC_272/Y NAND2X1_LOC_99/A 0.10fF
C61815 NOR2X1_LOC_207/A INVX1_LOC_54/A 0.02fF
C61816 NOR2X1_LOC_15/Y NOR2X1_LOC_465/Y 0.02fF
C61817 NOR2X1_LOC_598/B NOR2X1_LOC_405/Y 0.03fF
C61818 NOR2X1_LOC_561/Y NOR2X1_LOC_266/B 0.00fF
C61819 NOR2X1_LOC_824/A INVX1_LOC_23/Y 0.06fF
C61820 NAND2X1_LOC_287/a_36_24# NOR2X1_LOC_652/Y 0.01fF
C61821 INVX1_LOC_10/A NAND2X1_LOC_453/A 0.05fF
C61822 INVX1_LOC_119/A INVX1_LOC_92/A 0.03fF
C61823 NOR2X1_LOC_471/Y INVX1_LOC_15/A 0.01fF
C61824 D_INPUT_0 INVX1_LOC_76/A 0.94fF
C61825 NAND2X1_LOC_554/a_36_24# NAND2X1_LOC_211/Y 0.00fF
C61826 NOR2X1_LOC_214/B NOR2X1_LOC_300/a_36_216# 0.00fF
C61827 INVX1_LOC_273/Y VDD 0.26fF
C61828 INVX1_LOC_182/A NOR2X1_LOC_600/Y 0.02fF
C61829 INVX1_LOC_23/A INVX1_LOC_306/Y 0.05fF
C61830 NOR2X1_LOC_457/A NOR2X1_LOC_334/Y 0.07fF
C61831 NAND2X1_LOC_555/Y INVX1_LOC_15/A 0.05fF
C61832 INVX1_LOC_273/Y NAND2X1_LOC_800/A 0.01fF
C61833 NOR2X1_LOC_237/Y NOR2X1_LOC_662/A 0.47fF
C61834 NOR2X1_LOC_493/B INVX1_LOC_92/A 0.02fF
C61835 NOR2X1_LOC_554/B NOR2X1_LOC_847/A 0.03fF
C61836 INVX1_LOC_71/A INVX1_LOC_19/A 0.16fF
C61837 NOR2X1_LOC_649/a_36_216# INVX1_LOC_63/A 0.00fF
C61838 NOR2X1_LOC_131/A NOR2X1_LOC_364/A 0.01fF
C61839 VDD NOR2X1_LOC_76/A 0.86fF
C61840 NOR2X1_LOC_503/Y INVX1_LOC_78/A 0.12fF
C61841 NOR2X1_LOC_277/a_36_216# INVX1_LOC_306/Y 0.00fF
C61842 INVX1_LOC_1/A NAND2X1_LOC_299/a_36_24# 0.00fF
C61843 NAND2X1_LOC_350/B INVX1_LOC_117/Y 0.00fF
C61844 NOR2X1_LOC_180/B VDD 0.09fF
C61845 INVX1_LOC_77/A NAND2X1_LOC_63/Y 0.73fF
C61846 INVX1_LOC_193/Y INVX1_LOC_91/A 0.03fF
C61847 NOR2X1_LOC_160/B INVX1_LOC_87/A 0.07fF
C61848 NOR2X1_LOC_264/Y INVX1_LOC_63/A 0.14fF
C61849 NOR2X1_LOC_552/A INPUT_0 0.03fF
C61850 NAND2X1_LOC_303/Y INVX1_LOC_296/Y 0.02fF
C61851 INVX1_LOC_246/A NAND2X1_LOC_175/Y 0.02fF
C61852 INVX1_LOC_226/A NOR2X1_LOC_862/B 0.03fF
C61853 INVX1_LOC_239/A NOR2X1_LOC_476/B 0.10fF
C61854 NOR2X1_LOC_738/A VDD 0.35fF
C61855 NOR2X1_LOC_309/Y NOR2X1_LOC_662/A 0.02fF
C61856 NOR2X1_LOC_717/A NOR2X1_LOC_440/B 0.01fF
C61857 NAND2X1_LOC_793/Y NAND2X1_LOC_286/B 0.00fF
C61858 INVX1_LOC_30/A NAND2X1_LOC_444/B 0.01fF
C61859 INVX1_LOC_132/A NOR2X1_LOC_89/A 0.01fF
C61860 INVX1_LOC_30/A NOR2X1_LOC_334/Y 0.21fF
C61861 NOR2X1_LOC_669/Y INVX1_LOC_53/A 0.03fF
C61862 NOR2X1_LOC_152/Y INVX1_LOC_42/A 0.08fF
C61863 NOR2X1_LOC_589/A NOR2X1_LOC_743/Y 0.03fF
C61864 NOR2X1_LOC_329/B NOR2X1_LOC_111/A 1.60fF
C61865 INVX1_LOC_28/A NAND2X1_LOC_804/Y 0.00fF
C61866 NAND2X1_LOC_853/Y NAND2X1_LOC_770/Y 0.03fF
C61867 NAND2X1_LOC_852/Y INVX1_LOC_297/A 1.15fF
C61868 INVX1_LOC_24/A INVX1_LOC_3/Y 0.19fF
C61869 INVX1_LOC_73/A VDD 0.13fF
C61870 NAND2X1_LOC_842/B NOR2X1_LOC_561/A 0.04fF
C61871 NAND2X1_LOC_551/a_36_24# NOR2X1_LOC_103/Y 0.00fF
C61872 INVX1_LOC_50/A NOR2X1_LOC_276/Y 0.03fF
C61873 INVX1_LOC_17/A INVX1_LOC_108/Y 0.04fF
C61874 INVX1_LOC_27/A NOR2X1_LOC_249/Y 0.19fF
C61875 NAND2X1_LOC_33/Y INVX1_LOC_12/A 0.03fF
C61876 INVX1_LOC_225/A NOR2X1_LOC_89/A 0.05fF
C61877 INVX1_LOC_49/A NOR2X1_LOC_812/A 0.01fF
C61878 INVX1_LOC_7/A INVX1_LOC_46/Y 0.11fF
C61879 INVX1_LOC_17/A INVX1_LOC_278/A 0.07fF
C61880 NOR2X1_LOC_569/A VDD 0.24fF
C61881 NAND2X1_LOC_860/A NAND2X1_LOC_793/Y 0.00fF
C61882 INVX1_LOC_45/A INVX1_LOC_26/Y 0.08fF
C61883 NOR2X1_LOC_703/a_36_216# NOR2X1_LOC_383/B 0.00fF
C61884 NAND2X1_LOC_51/B INVX1_LOC_77/Y 0.05fF
C61885 NOR2X1_LOC_720/a_36_216# NAND2X1_LOC_74/B 0.00fF
C61886 INVX1_LOC_21/A INVX1_LOC_235/Y 0.15fF
C61887 NOR2X1_LOC_261/Y NOR2X1_LOC_471/Y 0.20fF
C61888 NOR2X1_LOC_557/A NAND2X1_LOC_447/Y 0.01fF
C61889 NOR2X1_LOC_704/Y VDD 0.24fF
C61890 INVX1_LOC_238/Y NAND2X1_LOC_725/Y 0.03fF
C61891 NOR2X1_LOC_486/a_36_216# INVX1_LOC_23/A 0.00fF
C61892 INVX1_LOC_21/A NAND2X1_LOC_149/Y 0.02fF
C61893 INVX1_LOC_17/A NOR2X1_LOC_489/a_36_216# 0.00fF
C61894 NOR2X1_LOC_168/B INVX1_LOC_69/A 0.38fF
C61895 INVX1_LOC_243/Y INVX1_LOC_36/A 0.00fF
C61896 INVX1_LOC_89/A INVX1_LOC_92/A 2.43fF
C61897 INVX1_LOC_75/A INVX1_LOC_114/A -0.01fF
C61898 INPUT_0 NOR2X1_LOC_813/Y 0.01fF
C61899 INVX1_LOC_142/A NOR2X1_LOC_727/B 0.34fF
C61900 NOR2X1_LOC_68/A NOR2X1_LOC_843/B 0.03fF
C61901 INVX1_LOC_108/Y NAND2X1_LOC_555/Y 0.03fF
C61902 INVX1_LOC_36/A INVX1_LOC_57/A 0.58fF
C61903 INVX1_LOC_42/Y NOR2X1_LOC_331/B 0.01fF
C61904 NOR2X1_LOC_152/Y INVX1_LOC_78/A 0.08fF
C61905 INVX1_LOC_136/A INVX1_LOC_50/A 0.13fF
C61906 INVX1_LOC_247/Y NOR2X1_LOC_383/B 0.02fF
C61907 NOR2X1_LOC_318/B NAND2X1_LOC_211/Y 0.06fF
C61908 NAND2X1_LOC_45/Y NOR2X1_LOC_865/Y 0.02fF
C61909 INVX1_LOC_113/Y INVX1_LOC_78/A 0.03fF
C61910 INPUT_0 INVX1_LOC_280/A 0.14fF
C61911 INVX1_LOC_287/A NOR2X1_LOC_68/A 0.04fF
C61912 NOR2X1_LOC_186/Y INVX1_LOC_11/A 0.14fF
C61913 NAND2X1_LOC_848/A NOR2X1_LOC_167/Y 0.03fF
C61914 NAND2X1_LOC_45/Y NOR2X1_LOC_243/B 0.19fF
C61915 INVX1_LOC_244/Y NOR2X1_LOC_638/Y -0.01fF
C61916 NOR2X1_LOC_168/a_36_216# INVX1_LOC_91/A 0.01fF
C61917 NAND2X1_LOC_21/Y NOR2X1_LOC_30/Y 0.05fF
C61918 NOR2X1_LOC_84/Y INVX1_LOC_32/A 0.10fF
C61919 NOR2X1_LOC_396/a_36_216# INVX1_LOC_46/A 0.02fF
C61920 INVX1_LOC_25/Y INVX1_LOC_12/A 0.16fF
C61921 NAND2X1_LOC_729/B VDD 0.28fF
C61922 NAND2X1_LOC_563/Y NOR2X1_LOC_38/B 0.10fF
C61923 NOR2X1_LOC_439/B INVX1_LOC_307/A 0.04fF
C61924 NOR2X1_LOC_828/B NOR2X1_LOC_155/A 0.15fF
C61925 NOR2X1_LOC_615/a_36_216# NOR2X1_LOC_496/Y 0.00fF
C61926 NAND2X1_LOC_99/Y INVX1_LOC_23/Y 0.04fF
C61927 INVX1_LOC_54/Y INVX1_LOC_47/Y 0.10fF
C61928 NOR2X1_LOC_65/B NOR2X1_LOC_152/Y 0.01fF
C61929 INVX1_LOC_90/A INVX1_LOC_119/Y 0.22fF
C61930 INVX1_LOC_277/A INVX1_LOC_213/A 0.06fF
C61931 NOR2X1_LOC_570/a_36_216# INVX1_LOC_53/A 0.01fF
C61932 INVX1_LOC_11/A NAND2X1_LOC_573/Y 0.62fF
C61933 INVX1_LOC_75/A INVX1_LOC_307/A 0.07fF
C61934 INVX1_LOC_31/A INVX1_LOC_306/Y 0.07fF
C61935 INVX1_LOC_58/A INVX1_LOC_24/A 0.13fF
C61936 NAND2X1_LOC_859/B INVX1_LOC_42/A 0.05fF
C61937 INVX1_LOC_136/A NAND2X1_LOC_72/Y 0.64fF
C61938 INVX1_LOC_75/A NOR2X1_LOC_445/B 0.01fF
C61939 VDD NAND2X1_LOC_241/Y 0.01fF
C61940 NOR2X1_LOC_266/B INVX1_LOC_76/A 0.03fF
C61941 INVX1_LOC_11/A NAND2X1_LOC_724/A 0.02fF
C61942 NOR2X1_LOC_681/Y INVX1_LOC_20/A 0.02fF
C61943 INVX1_LOC_139/A NAND2X1_LOC_211/Y 0.15fF
C61944 INVX1_LOC_37/A INVX1_LOC_20/A 0.03fF
C61945 INVX1_LOC_12/Y INVX1_LOC_59/Y 0.00fF
C61946 NOR2X1_LOC_209/A INVX1_LOC_117/A -0.00fF
C61947 NAND2X1_LOC_310/a_36_24# NOR2X1_LOC_383/B 0.01fF
C61948 INVX1_LOC_222/Y NOR2X1_LOC_336/B 0.01fF
C61949 INVX1_LOC_102/Y NOR2X1_LOC_653/Y 0.01fF
C61950 INVX1_LOC_8/A NOR2X1_LOC_383/B 0.02fF
C61951 NOR2X1_LOC_703/B INVX1_LOC_50/Y 0.03fF
C61952 INVX1_LOC_256/A INVX1_LOC_73/Y 0.01fF
C61953 INVX1_LOC_58/A NOR2X1_LOC_557/Y 0.15fF
C61954 NOR2X1_LOC_92/Y NOR2X1_LOC_441/Y 0.03fF
C61955 INVX1_LOC_269/A INVX1_LOC_292/A 0.01fF
C61956 NOR2X1_LOC_311/a_36_216# NOR2X1_LOC_743/Y 0.00fF
C61957 NOR2X1_LOC_78/B NOR2X1_LOC_856/a_36_216# 0.02fF
C61958 NAND2X1_LOC_725/A NAND2X1_LOC_740/A 0.07fF
C61959 NAND2X1_LOC_357/B NOR2X1_LOC_654/A 0.01fF
C61960 NOR2X1_LOC_309/Y INVX1_LOC_57/A 0.07fF
C61961 NAND2X1_LOC_9/Y INVX1_LOC_33/A 1.09fF
C61962 NAND2X1_LOC_848/A INVX1_LOC_76/A 0.10fF
C61963 NOR2X1_LOC_554/B NOR2X1_LOC_655/a_36_216# 0.00fF
C61964 INVX1_LOC_53/Y NOR2X1_LOC_248/A 0.01fF
C61965 NAND2X1_LOC_861/Y INVX1_LOC_42/A 0.29fF
C61966 NOR2X1_LOC_82/A NOR2X1_LOC_160/B 0.13fF
C61967 INVX1_LOC_90/A INVX1_LOC_284/A 0.23fF
C61968 NOR2X1_LOC_78/A NOR2X1_LOC_858/a_36_216# 0.00fF
C61969 NOR2X1_LOC_344/A INVX1_LOC_58/Y 0.01fF
C61970 INVX1_LOC_233/A INVX1_LOC_33/A 0.07fF
C61971 INVX1_LOC_205/A NAND2X1_LOC_473/A 0.00fF
C61972 NOR2X1_LOC_199/B INVX1_LOC_15/A 0.38fF
C61973 INVX1_LOC_36/A NOR2X1_LOC_666/Y 0.01fF
C61974 INVX1_LOC_21/A NOR2X1_LOC_744/Y 0.02fF
C61975 NOR2X1_LOC_130/A INVX1_LOC_3/Y 0.49fF
C61976 INVX1_LOC_22/A NOR2X1_LOC_36/A 0.16fF
C61977 INVX1_LOC_123/A NAND2X1_LOC_73/a_36_24# 0.00fF
C61978 INVX1_LOC_119/A INVX1_LOC_53/A 0.13fF
C61979 NOR2X1_LOC_15/Y NOR2X1_LOC_270/Y 0.19fF
C61980 NOR2X1_LOC_186/Y NOR2X1_LOC_433/A 0.39fF
C61981 NOR2X1_LOC_78/B NOR2X1_LOC_748/A 0.03fF
C61982 NOR2X1_LOC_351/Y INVX1_LOC_46/A 1.69fF
C61983 NOR2X1_LOC_177/Y INVX1_LOC_20/A 0.06fF
C61984 INVX1_LOC_45/A INVX1_LOC_161/Y 0.07fF
C61985 INVX1_LOC_58/A INVX1_LOC_143/A 0.07fF
C61986 INVX1_LOC_75/A INVX1_LOC_12/A 0.20fF
C61987 NOR2X1_LOC_359/Y NOR2X1_LOC_348/Y 0.11fF
C61988 INVX1_LOC_137/A INVX1_LOC_23/Y 0.01fF
C61989 NAND2X1_LOC_733/Y NOR2X1_LOC_599/Y 0.03fF
C61990 NOR2X1_LOC_540/B NOR2X1_LOC_155/A 0.01fF
C61991 NOR2X1_LOC_493/B INVX1_LOC_53/A 0.02fF
C61992 NOR2X1_LOC_468/Y INVX1_LOC_181/Y 0.02fF
C61993 INVX1_LOC_20/A NOR2X1_LOC_743/Y 0.05fF
C61994 NOR2X1_LOC_798/A INVX1_LOC_33/A 0.03fF
C61995 NAND2X1_LOC_348/A INVX1_LOC_284/A 0.01fF
C61996 NOR2X1_LOC_667/Y INVX1_LOC_141/Y 0.00fF
C61997 NAND2X1_LOC_364/Y NOR2X1_LOC_852/Y 0.02fF
C61998 NAND2X1_LOC_79/Y INVX1_LOC_14/A 0.04fF
C61999 INVX1_LOC_76/A INVX1_LOC_46/Y 0.15fF
C62000 INVX1_LOC_164/A INVX1_LOC_26/A 0.09fF
C62001 NOR2X1_LOC_208/Y NOR2X1_LOC_666/Y 0.12fF
C62002 INVX1_LOC_27/A NOR2X1_LOC_722/a_36_216# 0.01fF
C62003 NAND2X1_LOC_861/Y INVX1_LOC_78/A 0.07fF
C62004 NAND2X1_LOC_349/a_36_24# INVX1_LOC_270/Y 0.01fF
C62005 INVX1_LOC_171/A NAND2X1_LOC_72/B 0.26fF
C62006 NAND2X1_LOC_67/Y INVX1_LOC_49/A 0.01fF
C62007 NOR2X1_LOC_186/Y NOR2X1_LOC_52/B 0.11fF
C62008 NAND2X1_LOC_9/Y INVX1_LOC_40/A 0.02fF
C62009 INVX1_LOC_8/A NAND2X1_LOC_75/a_36_24# 0.00fF
C62010 INVX1_LOC_45/A INVX1_LOC_312/A 0.01fF
C62011 NAND2X1_LOC_9/Y INVX1_LOC_165/Y 0.01fF
C62012 INVX1_LOC_136/A INVX1_LOC_61/Y 0.03fF
C62013 INVX1_LOC_27/A NAND2X1_LOC_116/A 0.03fF
C62014 NOR2X1_LOC_45/B INVX1_LOC_49/Y 0.04fF
C62015 INVX1_LOC_83/A NOR2X1_LOC_798/Y 0.01fF
C62016 INVX1_LOC_25/A INVX1_LOC_13/A 0.26fF
C62017 INVX1_LOC_24/A INVX1_LOC_215/Y 0.58fF
C62018 NAND2X1_LOC_117/a_36_24# INVX1_LOC_26/A 0.00fF
C62019 INVX1_LOC_161/Y INVX1_LOC_71/A 0.07fF
C62020 NOR2X1_LOC_188/Y INVX1_LOC_29/Y 0.06fF
C62021 INVX1_LOC_83/A NOR2X1_LOC_635/B 0.03fF
C62022 INVX1_LOC_286/A INVX1_LOC_168/Y 0.02fF
C62023 INVX1_LOC_2/A NOR2X1_LOC_626/a_36_216# 0.02fF
C62024 NOR2X1_LOC_749/Y INVX1_LOC_26/Y 0.02fF
C62025 INVX1_LOC_132/A INVX1_LOC_11/A 0.07fF
C62026 INVX1_LOC_265/A NOR2X1_LOC_15/Y 0.01fF
C62027 NAND2X1_LOC_573/Y NOR2X1_LOC_52/B 0.07fF
C62028 NOR2X1_LOC_594/Y INVX1_LOC_15/A 0.30fF
C62029 INVX1_LOC_17/A NAND2X1_LOC_21/Y 0.12fF
C62030 INVX1_LOC_57/Y NAND2X1_LOC_634/Y 0.10fF
C62031 NOR2X1_LOC_366/Y INVX1_LOC_271/A 0.02fF
C62032 INVX1_LOC_249/A NOR2X1_LOC_596/Y 0.04fF
C62033 INVX1_LOC_130/A NOR2X1_LOC_759/Y 0.00fF
C62034 NAND2X1_LOC_569/a_36_24# INVX1_LOC_61/A 0.01fF
C62035 INVX1_LOC_58/A NOR2X1_LOC_130/A 0.03fF
C62036 INVX1_LOC_269/A INVX1_LOC_240/A 0.03fF
C62037 NOR2X1_LOC_45/Y NOR2X1_LOC_433/A 0.01fF
C62038 NOR2X1_LOC_89/A NAND2X1_LOC_642/Y 0.09fF
C62039 NAND2X1_LOC_214/B INVX1_LOC_232/A 0.51fF
C62040 INVX1_LOC_88/A NOR2X1_LOC_574/A 0.06fF
C62041 INVX1_LOC_108/Y NOR2X1_LOC_199/B 0.36fF
C62042 NOR2X1_LOC_68/A INVX1_LOC_18/A 0.41fF
C62043 NOR2X1_LOC_78/A NOR2X1_LOC_159/a_36_216# 0.00fF
C62044 INVX1_LOC_64/A NOR2X1_LOC_757/A 0.06fF
C62045 INVX1_LOC_11/A INVX1_LOC_225/A 0.09fF
C62046 NOR2X1_LOC_332/Y INVX1_LOC_152/A 0.08fF
C62047 NOR2X1_LOC_388/Y INVX1_LOC_225/Y 0.10fF
C62048 NAND2X1_LOC_347/B NAND2X1_LOC_360/B 0.04fF
C62049 INVX1_LOC_2/A NAND2X1_LOC_67/Y 0.14fF
C62050 NOR2X1_LOC_632/Y INVX1_LOC_5/A 0.06fF
C62051 INVX1_LOC_247/A INVX1_LOC_99/A 0.00fF
C62052 INVX1_LOC_92/Y INVX1_LOC_4/Y 0.02fF
C62053 NOR2X1_LOC_639/B NOR2X1_LOC_763/Y 0.03fF
C62054 NAND2X1_LOC_390/a_36_24# INVX1_LOC_93/A 0.00fF
C62055 INVX1_LOC_222/A NAND2X1_LOC_72/B 0.72fF
C62056 INVX1_LOC_223/A NOR2X1_LOC_106/Y 0.00fF
C62057 NOR2X1_LOC_33/A NOR2X1_LOC_34/B 0.02fF
C62058 INVX1_LOC_89/A INVX1_LOC_53/A 2.09fF
C62059 INVX1_LOC_27/A INVX1_LOC_232/A 0.11fF
C62060 INVX1_LOC_21/A INVX1_LOC_16/A 0.11fF
C62061 NAND2X1_LOC_364/A NAND2X1_LOC_656/A 0.17fF
C62062 INVX1_LOC_136/A NAND2X1_LOC_845/a_36_24# 0.01fF
C62063 INVX1_LOC_22/A NAND2X1_LOC_474/Y 0.14fF
C62064 NAND2X1_LOC_45/Y NOR2X1_LOC_342/A 0.02fF
C62065 NOR2X1_LOC_356/A INVX1_LOC_23/A 0.30fF
C62066 NOR2X1_LOC_15/Y NOR2X1_LOC_458/B 0.00fF
C62067 INVX1_LOC_38/A INVX1_LOC_119/Y 0.01fF
C62068 INVX1_LOC_313/Y NOR2X1_LOC_493/a_36_216# 0.00fF
C62069 INVX1_LOC_164/Y NOR2X1_LOC_361/B 0.10fF
C62070 NAND2X1_LOC_736/Y NAND2X1_LOC_733/Y 0.10fF
C62071 NAND2X1_LOC_350/A NAND2X1_LOC_477/A 0.03fF
C62072 NOR2X1_LOC_355/B INVX1_LOC_4/Y 0.09fF
C62073 INVX1_LOC_11/A NOR2X1_LOC_209/Y 0.15fF
C62074 NOR2X1_LOC_598/B NOR2X1_LOC_644/A 0.02fF
C62075 INVX1_LOC_12/A NAND2X1_LOC_453/A 0.14fF
C62076 NOR2X1_LOC_91/A NOR2X1_LOC_74/A 0.12fF
C62077 INVX1_LOC_27/A NOR2X1_LOC_383/Y 0.51fF
C62078 NAND2X1_LOC_254/Y NAND2X1_LOC_464/A 0.00fF
C62079 NOR2X1_LOC_813/Y NOR2X1_LOC_84/B -0.08fF
C62080 NAND2X1_LOC_30/Y INVX1_LOC_243/A 0.02fF
C62081 INVX1_LOC_172/A NOR2X1_LOC_68/A 0.22fF
C62082 NAND2X1_LOC_394/a_36_24# INVX1_LOC_89/A 0.00fF
C62083 NOR2X1_LOC_772/Y INVX1_LOC_72/A 0.01fF
C62084 NOR2X1_LOC_590/A NOR2X1_LOC_174/a_36_216# 0.00fF
C62085 INVX1_LOC_97/Y NOR2X1_LOC_644/A 0.01fF
C62086 NOR2X1_LOC_441/Y NAND2X1_LOC_477/A 0.03fF
C62087 INVX1_LOC_81/A NOR2X1_LOC_759/Y 0.30fF
C62088 INVX1_LOC_7/Y NOR2X1_LOC_99/B -0.01fF
C62089 INVX1_LOC_49/A NOR2X1_LOC_324/Y 0.01fF
C62090 INVX1_LOC_14/Y INVX1_LOC_290/Y 0.10fF
C62091 INVX1_LOC_27/A NOR2X1_LOC_366/Y 0.06fF
C62092 NOR2X1_LOC_331/B INVX1_LOC_19/A 0.07fF
C62093 INVX1_LOC_13/A INVX1_LOC_1/A 0.23fF
C62094 INVX1_LOC_280/A NOR2X1_LOC_84/B 0.08fF
C62095 NOR2X1_LOC_226/A NOR2X1_LOC_331/Y 0.00fF
C62096 NOR2X1_LOC_392/B INVX1_LOC_72/A 0.25fF
C62097 INVX1_LOC_200/A INVX1_LOC_25/Y 0.03fF
C62098 NOR2X1_LOC_74/A INVX1_LOC_23/A 0.15fF
C62099 INVX1_LOC_136/A NOR2X1_LOC_773/a_36_216# 0.00fF
C62100 INVX1_LOC_13/Y INVX1_LOC_47/A 0.00fF
C62101 INVX1_LOC_71/A NAND2X1_LOC_119/a_36_24# 0.00fF
C62102 NOR2X1_LOC_457/B INVX1_LOC_153/Y 0.10fF
C62103 INVX1_LOC_50/A NOR2X1_LOC_165/a_36_216# 0.00fF
C62104 NOR2X1_LOC_82/A NOR2X1_LOC_516/B 0.09fF
C62105 NAND2X1_LOC_53/Y INVX1_LOC_22/A 0.09fF
C62106 INVX1_LOC_101/Y INVX1_LOC_279/A 0.02fF
C62107 NAND2X1_LOC_559/Y INVX1_LOC_229/Y 0.49fF
C62108 NAND2X1_LOC_63/Y INVX1_LOC_9/A 0.05fF
C62109 NAND2X1_LOC_849/B INVX1_LOC_284/A 0.04fF
C62110 NOR2X1_LOC_295/Y INVX1_LOC_181/Y 0.02fF
C62111 NOR2X1_LOC_457/A NOR2X1_LOC_569/Y 0.01fF
C62112 INVX1_LOC_38/A INVX1_LOC_284/A 0.07fF
C62113 INVX1_LOC_180/A INVX1_LOC_63/Y 0.10fF
C62114 NAND2X1_LOC_175/B NAND2X1_LOC_593/Y 0.37fF
C62115 INVX1_LOC_24/A NOR2X1_LOC_344/a_36_216# 0.02fF
C62116 NAND2X1_LOC_134/a_36_24# INVX1_LOC_18/A 0.00fF
C62117 INVX1_LOC_21/A INVX1_LOC_28/A 0.26fF
C62118 NAND2X1_LOC_181/a_36_24# NOR2X1_LOC_160/B 0.00fF
C62119 NOR2X1_LOC_272/Y NOR2X1_LOC_329/B 0.10fF
C62120 NOR2X1_LOC_624/A INVX1_LOC_77/A 0.10fF
C62121 INVX1_LOC_1/A NOR2X1_LOC_174/B 0.02fF
C62122 NOR2X1_LOC_710/B INVX1_LOC_83/A 0.06fF
C62123 NOR2X1_LOC_592/B INVX1_LOC_19/A 0.06fF
C62124 NOR2X1_LOC_361/B NOR2X1_LOC_76/A 0.01fF
C62125 INVX1_LOC_239/A INVX1_LOC_169/A 0.03fF
C62126 NOR2X1_LOC_78/B NOR2X1_LOC_570/a_36_216# 0.02fF
C62127 INVX1_LOC_225/A NOR2X1_LOC_433/A 0.28fF
C62128 INVX1_LOC_55/Y INVX1_LOC_1/A 0.07fF
C62129 NAND2X1_LOC_783/A INVX1_LOC_215/Y 0.00fF
C62130 INVX1_LOC_158/A NOR2X1_LOC_350/A 0.08fF
C62131 NOR2X1_LOC_34/A INVX1_LOC_75/A 0.01fF
C62132 NAND2X1_LOC_741/B NOR2X1_LOC_695/Y 0.06fF
C62133 INVX1_LOC_225/A NOR2X1_LOC_593/Y 0.20fF
C62134 NOR2X1_LOC_160/B INVX1_LOC_306/A 0.03fF
C62135 NAND2X1_LOC_848/Y INVX1_LOC_284/A 0.13fF
C62136 INVX1_LOC_291/A INVX1_LOC_42/A 0.07fF
C62137 NOR2X1_LOC_661/a_36_216# NOR2X1_LOC_661/A 0.01fF
C62138 INVX1_LOC_248/A NOR2X1_LOC_744/Y 0.02fF
C62139 NOR2X1_LOC_720/B NAND2X1_LOC_518/a_36_24# 0.00fF
C62140 INVX1_LOC_104/A NOR2X1_LOC_551/B 0.12fF
C62141 NOR2X1_LOC_52/B NAND2X1_LOC_640/Y 0.00fF
C62142 INVX1_LOC_6/A INVX1_LOC_306/Y 0.15fF
C62143 NOR2X1_LOC_662/A INVX1_LOC_63/A 0.02fF
C62144 NOR2X1_LOC_601/a_36_216# INVX1_LOC_96/A 0.00fF
C62145 NAND2X1_LOC_149/Y NAND2X1_LOC_51/B 0.10fF
C62146 NAND2X1_LOC_802/Y INVX1_LOC_42/A 0.03fF
C62147 INVX1_LOC_101/Y INVX1_LOC_182/Y 0.02fF
C62148 NAND2X1_LOC_82/Y NOR2X1_LOC_649/B 0.10fF
C62149 NOR2X1_LOC_372/A NOR2X1_LOC_71/Y 0.22fF
C62150 INVX1_LOC_100/A NAND2X1_LOC_474/Y 0.05fF
C62151 NOR2X1_LOC_388/Y INVX1_LOC_266/Y 0.24fF
C62152 INVX1_LOC_225/A NOR2X1_LOC_52/B 0.10fF
C62153 INVX1_LOC_213/Y INVX1_LOC_104/A 0.21fF
C62154 INVX1_LOC_174/Y NOR2X1_LOC_546/A 0.01fF
C62155 NOR2X1_LOC_10/a_36_216# INVX1_LOC_306/Y 0.01fF
C62156 NOR2X1_LOC_643/A INVX1_LOC_75/A 0.03fF
C62157 INVX1_LOC_64/A NOR2X1_LOC_396/Y 0.00fF
C62158 NOR2X1_LOC_589/A NAND2X1_LOC_198/B 0.10fF
C62159 INVX1_LOC_50/Y INVX1_LOC_91/A 0.07fF
C62160 INVX1_LOC_41/A NOR2X1_LOC_655/B 0.03fF
C62161 NOR2X1_LOC_91/A NOR2X1_LOC_690/a_36_216# 0.00fF
C62162 NOR2X1_LOC_500/Y NOR2X1_LOC_577/Y 0.09fF
C62163 INVX1_LOC_35/A INVX1_LOC_126/A 0.03fF
C62164 NOR2X1_LOC_772/B INVX1_LOC_95/Y 0.06fF
C62165 NOR2X1_LOC_596/a_36_216# INVX1_LOC_16/A 0.00fF
C62166 NAND2X1_LOC_338/B NOR2X1_LOC_392/B 0.10fF
C62167 INVX1_LOC_2/A NOR2X1_LOC_367/B 0.01fF
C62168 INVX1_LOC_8/Y INVX1_LOC_1/Y 0.01fF
C62169 NAND2X1_LOC_99/Y INVX1_LOC_232/A 0.39fF
C62170 NOR2X1_LOC_103/Y NAND2X1_LOC_270/a_36_24# 0.00fF
C62171 INVX1_LOC_159/A NAND2X1_LOC_155/a_36_24# 0.00fF
C62172 INVX1_LOC_90/A INVX1_LOC_72/A 0.12fF
C62173 INVX1_LOC_78/A INVX1_LOC_291/A 0.06fF
C62174 INVX1_LOC_13/Y INVX1_LOC_95/Y 0.37fF
C62175 INVX1_LOC_58/A NAND2X1_LOC_811/B 0.01fF
C62176 NAND2X1_LOC_721/a_36_24# NOR2X1_LOC_667/A 0.00fF
C62177 NOR2X1_LOC_389/B INVX1_LOC_72/A 0.10fF
C62178 INVX1_LOC_78/A NAND2X1_LOC_802/Y 0.03fF
C62179 INVX1_LOC_64/A NOR2X1_LOC_681/Y 0.00fF
C62180 INVX1_LOC_266/A INVX1_LOC_91/A 0.10fF
C62181 INVX1_LOC_64/A INVX1_LOC_37/A 2.52fF
C62182 NOR2X1_LOC_561/Y INVX1_LOC_49/A 0.07fF
C62183 INVX1_LOC_27/A INVX1_LOC_74/Y 0.02fF
C62184 INVX1_LOC_35/A NOR2X1_LOC_111/A 0.02fF
C62185 INVX1_LOC_224/A NAND2X1_LOC_669/a_36_24# 0.00fF
C62186 NOR2X1_LOC_88/Y INVX1_LOC_94/Y 0.07fF
C62187 INVX1_LOC_17/A INVX1_LOC_123/A 0.03fF
C62188 NOR2X1_LOC_264/Y INVX1_LOC_1/Y 0.07fF
C62189 NOR2X1_LOC_577/Y INVX1_LOC_10/A 0.21fF
C62190 NOR2X1_LOC_274/Y D_INPUT_0 0.00fF
C62191 INVX1_LOC_208/Y INVX1_LOC_104/A 0.01fF
C62192 INVX1_LOC_90/A INVX1_LOC_198/Y 0.01fF
C62193 INVX1_LOC_298/Y INVX1_LOC_179/A 0.03fF
C62194 INVX1_LOC_31/A NOR2X1_LOC_74/A 0.07fF
C62195 NAND2X1_LOC_785/Y INVX1_LOC_16/A 0.22fF
C62196 INVX1_LOC_41/A NAND2X1_LOC_358/Y 0.03fF
C62197 INVX1_LOC_21/A NOR2X1_LOC_35/Y 0.08fF
C62198 NOR2X1_LOC_454/Y NAND2X1_LOC_212/Y 0.02fF
C62199 NOR2X1_LOC_65/B INVX1_LOC_291/A 0.04fF
C62200 INVX1_LOC_227/A INVX1_LOC_155/Y 0.02fF
C62201 NOR2X1_LOC_216/B INVX1_LOC_23/Y 0.07fF
C62202 NOR2X1_LOC_590/a_36_216# INVX1_LOC_18/A 0.00fF
C62203 INVX1_LOC_14/A NOR2X1_LOC_80/a_36_216# 0.02fF
C62204 INVX1_LOC_31/A NOR2X1_LOC_9/Y 0.05fF
C62205 NOR2X1_LOC_717/B NOR2X1_LOC_344/A 0.00fF
C62206 INVX1_LOC_84/A INVX1_LOC_94/Y 0.03fF
C62207 NAND2X1_LOC_479/Y INVX1_LOC_266/Y 0.07fF
C62208 NOR2X1_LOC_89/A NAND2X1_LOC_792/B 0.03fF
C62209 INVX1_LOC_303/A INVX1_LOC_47/A 0.06fF
C62210 INVX1_LOC_224/A NAND2X1_LOC_642/Y 0.02fF
C62211 INVX1_LOC_269/A NOR2X1_LOC_542/B 0.01fF
C62212 INVX1_LOC_147/A INVX1_LOC_18/A 0.06fF
C62213 NAND2X1_LOC_568/A INVX1_LOC_291/Y 0.00fF
C62214 NAND2X1_LOC_794/B NAND2X1_LOC_804/Y 0.02fF
C62215 INVX1_LOC_11/A NAND2X1_LOC_642/Y 0.13fF
C62216 INVX1_LOC_226/Y NOR2X1_LOC_346/B 0.07fF
C62217 NOR2X1_LOC_438/a_36_216# INVX1_LOC_304/A 0.00fF
C62218 INVX1_LOC_103/A NOR2X1_LOC_275/A 0.01fF
C62219 NOR2X1_LOC_667/A INVX1_LOC_16/A 5.16fF
C62220 NOR2X1_LOC_798/A NOR2X1_LOC_537/a_36_216# 0.00fF
C62221 INVX1_LOC_225/Y NOR2X1_LOC_552/A 0.10fF
C62222 NOR2X1_LOC_657/Y INVX1_LOC_6/A 0.04fF
C62223 NOR2X1_LOC_201/A NOR2X1_LOC_243/B -0.02fF
C62224 INVX1_LOC_1/A NOR2X1_LOC_357/Y 0.00fF
C62225 NAND2X1_LOC_734/B NAND2X1_LOC_808/A 0.02fF
C62226 INVX1_LOC_2/A NOR2X1_LOC_561/Y 0.14fF
C62227 INVX1_LOC_267/A NOR2X1_LOC_459/A 0.01fF
C62228 INVX1_LOC_33/A NAND2X1_LOC_842/B 0.03fF
C62229 INVX1_LOC_2/A INVX1_LOC_7/A 0.00fF
C62230 NAND2X1_LOC_477/Y INVX1_LOC_23/Y 0.01fF
C62231 NOR2X1_LOC_147/B INVX1_LOC_313/Y 0.02fF
C62232 NOR2X1_LOC_500/Y INVX1_LOC_22/A 0.07fF
C62233 INVX1_LOC_269/A NOR2X1_LOC_137/Y 0.01fF
C62234 NAND2X1_LOC_361/Y NAND2X1_LOC_7/a_36_24# 0.00fF
C62235 NOR2X1_LOC_226/A NOR2X1_LOC_561/Y 0.15fF
C62236 INVX1_LOC_215/A NOR2X1_LOC_136/Y 0.13fF
C62237 NOR2X1_LOC_265/a_36_216# NAND2X1_LOC_390/A 0.00fF
C62238 NOR2X1_LOC_392/B INVX1_LOC_313/Y 0.02fF
C62239 NAND2X1_LOC_30/Y INVX1_LOC_76/A 0.01fF
C62240 NOR2X1_LOC_248/Y INVX1_LOC_91/A 0.06fF
C62241 NOR2X1_LOC_160/B INVX1_LOC_59/Y 0.72fF
C62242 INVX1_LOC_84/A INVX1_LOC_296/A 0.01fF
C62243 NOR2X1_LOC_544/A INVX1_LOC_279/A 0.07fF
C62244 NOR2X1_LOC_113/a_36_216# NOR2X1_LOC_814/A 0.00fF
C62245 INVX1_LOC_39/A INVX1_LOC_9/A 0.17fF
C62246 NOR2X1_LOC_589/A INVX1_LOC_53/Y 0.03fF
C62247 NOR2X1_LOC_470/B INVX1_LOC_117/A 0.01fF
C62248 INVX1_LOC_57/A NOR2X1_LOC_654/a_36_216# 0.00fF
C62249 NOR2X1_LOC_180/B INVX1_LOC_177/A 0.03fF
C62250 NOR2X1_LOC_218/Y NOR2X1_LOC_561/Y 0.02fF
C62251 INVX1_LOC_57/A INVX1_LOC_63/A 0.28fF
C62252 INVX1_LOC_181/Y INVX1_LOC_100/Y 0.04fF
C62253 INVX1_LOC_49/A NOR2X1_LOC_835/B 0.00fF
C62254 INVX1_LOC_84/A NAND2X1_LOC_205/a_36_24# 0.00fF
C62255 NOR2X1_LOC_78/B INVX1_LOC_89/A 0.14fF
C62256 NAND2X1_LOC_723/a_36_24# NOR2X1_LOC_380/A 0.01fF
C62257 INVX1_LOC_90/A NOR2X1_LOC_537/Y 0.07fF
C62258 INVX1_LOC_101/A NOR2X1_LOC_188/Y 0.11fF
C62259 INVX1_LOC_10/A INVX1_LOC_22/A 0.94fF
C62260 INVX1_LOC_90/A NAND2X1_LOC_338/B 0.08fF
C62261 INVX1_LOC_49/A INVX1_LOC_303/Y 0.01fF
C62262 NOR2X1_LOC_122/A NOR2X1_LOC_331/B 0.01fF
C62263 NOR2X1_LOC_457/A NAND2X1_LOC_472/Y 0.14fF
C62264 NAND2X1_LOC_288/B INVX1_LOC_29/A 0.00fF
C62265 NOR2X1_LOC_389/B NOR2X1_LOC_537/Y 0.13fF
C62266 NAND2X1_LOC_651/B INVX1_LOC_296/A 0.04fF
C62267 NAND2X1_LOC_860/Y NAND2X1_LOC_861/Y 0.10fF
C62268 INVX1_LOC_145/Y NOR2X1_LOC_589/A 0.01fF
C62269 NAND2X1_LOC_733/Y NAND2X1_LOC_453/A 0.05fF
C62270 NAND2X1_LOC_190/a_36_24# NOR2X1_LOC_197/B 0.06fF
C62271 NAND2X1_LOC_711/Y INVX1_LOC_46/A 0.01fF
C62272 INVX1_LOC_314/Y INVX1_LOC_98/A 0.04fF
C62273 NOR2X1_LOC_667/A INVX1_LOC_28/A 0.26fF
C62274 INVX1_LOC_73/A INVX1_LOC_177/A 0.06fF
C62275 INVX1_LOC_94/Y INVX1_LOC_15/A 0.68fF
C62276 NAND2X1_LOC_541/a_36_24# INVX1_LOC_63/A 0.01fF
C62277 NAND2X1_LOC_656/A NOR2X1_LOC_405/A 0.00fF
C62278 INVX1_LOC_314/Y NOR2X1_LOC_78/A 1.25fF
C62279 INVX1_LOC_11/A NOR2X1_LOC_271/Y 0.03fF
C62280 INVX1_LOC_248/A INVX1_LOC_28/A 0.07fF
C62281 NAND2X1_LOC_85/Y NOR2X1_LOC_849/A 0.49fF
C62282 NOR2X1_LOC_355/A NOR2X1_LOC_188/Y 0.00fF
C62283 NAND2X1_LOC_72/B INVX1_LOC_4/A 1.97fF
C62284 NAND2X1_LOC_198/B INVX1_LOC_147/Y 0.71fF
C62285 NAND2X1_LOC_11/Y D_INPUT_4 0.03fF
C62286 NAND2X1_LOC_348/A NOR2X1_LOC_537/Y 0.03fF
C62287 NOR2X1_LOC_406/A INVX1_LOC_285/A 0.01fF
C62288 NOR2X1_LOC_569/A INVX1_LOC_177/A 0.01fF
C62289 NOR2X1_LOC_318/B INVX1_LOC_155/A 0.07fF
C62290 NAND2X1_LOC_198/B INVX1_LOC_20/A 0.03fF
C62291 INVX1_LOC_39/Y NOR2X1_LOC_536/A 0.21fF
C62292 NOR2X1_LOC_433/A NAND2X1_LOC_642/Y 0.01fF
C62293 INVX1_LOC_14/A INVX1_LOC_70/A 0.01fF
C62294 INVX1_LOC_251/Y INPUT_0 0.02fF
C62295 INVX1_LOC_89/A NOR2X1_LOC_459/A 0.62fF
C62296 NOR2X1_LOC_19/B INVX1_LOC_232/A 0.12fF
C62297 INVX1_LOC_30/A NAND2X1_LOC_472/Y 0.07fF
C62298 NAND2X1_LOC_514/Y NAND2X1_LOC_211/Y 0.03fF
C62299 INVX1_LOC_303/A INVX1_LOC_95/Y 0.10fF
C62300 INVX1_LOC_34/A NOR2X1_LOC_45/B 7.63fF
C62301 INVX1_LOC_141/Y NOR2X1_LOC_536/A 0.01fF
C62302 INVX1_LOC_2/A NOR2X1_LOC_167/Y 0.03fF
C62303 NOR2X1_LOC_704/Y INVX1_LOC_177/A 0.16fF
C62304 NOR2X1_LOC_322/Y NAND2X1_LOC_862/A 0.12fF
C62305 INVX1_LOC_181/A INVX1_LOC_15/A 0.05fF
C62306 INVX1_LOC_89/A INVX1_LOC_83/A 0.19fF
C62307 INVX1_LOC_312/Y NOR2X1_LOC_536/A 0.01fF
C62308 NOR2X1_LOC_6/B INVX1_LOC_91/A 4.11fF
C62309 INVX1_LOC_296/A INVX1_LOC_15/A 0.04fF
C62310 INVX1_LOC_262/A NOR2X1_LOC_467/A 0.01fF
C62311 NOR2X1_LOC_226/A NOR2X1_LOC_167/Y 0.03fF
C62312 INVX1_LOC_14/A INVX1_LOC_123/Y 0.02fF
C62313 NOR2X1_LOC_722/Y INVX1_LOC_281/A 0.10fF
C62314 NOR2X1_LOC_723/Y INVX1_LOC_281/Y 0.31fF
C62315 NOR2X1_LOC_791/Y NAND2X1_LOC_773/B 0.02fF
C62316 NAND2X1_LOC_98/a_36_24# INVX1_LOC_84/A 0.00fF
C62317 NOR2X1_LOC_78/B NOR2X1_LOC_703/Y 0.00fF
C62318 INVX1_LOC_159/A INVX1_LOC_117/A 0.07fF
C62319 INVX1_LOC_49/A INVX1_LOC_76/A 0.22fF
C62320 NOR2X1_LOC_503/Y NAND2X1_LOC_802/Y -0.00fF
C62321 INVX1_LOC_25/A INVX1_LOC_32/A 1.17fF
C62322 INVX1_LOC_83/A NAND2X1_LOC_508/A 0.24fF
C62323 INVX1_LOC_72/A INVX1_LOC_38/A 0.54fF
C62324 INVX1_LOC_34/A INVX1_LOC_199/Y 0.02fF
C62325 NOR2X1_LOC_372/A NAND2X1_LOC_243/Y 0.00fF
C62326 INVX1_LOC_313/Y INVX1_LOC_97/A 0.01fF
C62327 INVX1_LOC_226/Y INVX1_LOC_100/A -0.00fF
C62328 NOR2X1_LOC_52/B NAND2X1_LOC_642/Y 0.03fF
C62329 INVX1_LOC_72/A NAND2X1_LOC_264/a_36_24# 0.01fF
C62330 INVX1_LOC_77/A INVX1_LOC_14/Y 0.03fF
C62331 INVX1_LOC_30/A NAND2X1_LOC_637/Y 0.09fF
C62332 INVX1_LOC_311/A INVX1_LOC_16/A 0.11fF
C62333 NOR2X1_LOC_759/Y NOR2X1_LOC_363/Y 0.01fF
C62334 NOR2X1_LOC_52/B NAND2X1_LOC_643/a_36_24# 0.00fF
C62335 NAND2X1_LOC_860/A INVX1_LOC_47/Y 0.02fF
C62336 INVX1_LOC_26/Y NOR2X1_LOC_621/B 0.01fF
C62337 INVX1_LOC_90/A INVX1_LOC_313/Y 0.07fF
C62338 INVX1_LOC_215/A INVX1_LOC_144/A 0.73fF
C62339 NAND2X1_LOC_231/Y NOR2X1_LOC_45/B 0.34fF
C62340 NOR2X1_LOC_620/Y VDD 0.29fF
C62341 INVX1_LOC_13/A NOR2X1_LOC_188/A 0.07fF
C62342 INVX1_LOC_202/A NOR2X1_LOC_363/Y 0.15fF
C62343 NAND2X1_LOC_283/a_36_24# INVX1_LOC_46/A 0.00fF
C62344 NAND2X1_LOC_794/B NOR2X1_LOC_519/a_36_216# 0.01fF
C62345 NOR2X1_LOC_181/a_36_216# INVX1_LOC_179/A 0.01fF
C62346 NOR2X1_LOC_189/A NAND2X1_LOC_804/Y 0.17fF
C62347 NOR2X1_LOC_778/B NOR2X1_LOC_78/A 1.41fF
C62348 INVX1_LOC_13/A NOR2X1_LOC_548/B 0.03fF
C62349 NAND2X1_LOC_332/Y NAND2X1_LOC_211/Y -0.02fF
C62350 INVX1_LOC_255/Y INVX1_LOC_201/A 0.04fF
C62351 INVX1_LOC_27/A NAND2X1_LOC_263/a_36_24# 0.00fF
C62352 INVX1_LOC_72/A NOR2X1_LOC_51/A 0.13fF
C62353 NAND2X1_LOC_350/A NOR2X1_LOC_435/B 0.15fF
C62354 NOR2X1_LOC_382/Y NOR2X1_LOC_104/a_36_216# 0.00fF
C62355 NOR2X1_LOC_68/A NOR2X1_LOC_860/Y 0.01fF
C62356 NOR2X1_LOC_543/A INVX1_LOC_69/Y 0.19fF
C62357 INVX1_LOC_293/A INVX1_LOC_84/A 0.01fF
C62358 NOR2X1_LOC_437/Y NOR2X1_LOC_331/B 0.10fF
C62359 NAND2X1_LOC_181/Y NOR2X1_LOC_123/a_36_216# 0.00fF
C62360 NAND2X1_LOC_276/Y INVX1_LOC_129/Y 0.14fF
C62361 INVX1_LOC_31/A NOR2X1_LOC_243/B 0.07fF
C62362 INVX1_LOC_41/A NOR2X1_LOC_176/Y 0.05fF
C62363 NOR2X1_LOC_631/B INVX1_LOC_44/Y 0.01fF
C62364 NOR2X1_LOC_731/A VDD 0.24fF
C62365 NAND2X1_LOC_53/Y INVX1_LOC_186/Y 1.15fF
C62366 INVX1_LOC_280/Y NOR2X1_LOC_24/a_36_216# 0.00fF
C62367 INVX1_LOC_2/A INVX1_LOC_76/A 4.64fF
C62368 INVX1_LOC_45/A NOR2X1_LOC_841/A 0.01fF
C62369 INVX1_LOC_30/Y INVX1_LOC_91/A 0.03fF
C62370 INVX1_LOC_36/A NOR2X1_LOC_820/Y 0.05fF
C62371 INVX1_LOC_34/A INVX1_LOC_281/A 0.34fF
C62372 INVX1_LOC_64/A NAND2X1_LOC_72/B 0.03fF
C62373 NAND2X1_LOC_483/Y NOR2X1_LOC_536/A 0.01fF
C62374 INVX1_LOC_266/Y INVX1_LOC_139/Y 0.06fF
C62375 NOR2X1_LOC_226/A INVX1_LOC_76/A 0.20fF
C62376 INVX1_LOC_14/A INVX1_LOC_102/A 0.09fF
C62377 NOR2X1_LOC_112/Y NOR2X1_LOC_196/Y 0.07fF
C62378 NOR2X1_LOC_799/B INVX1_LOC_22/A 0.01fF
C62379 INVX1_LOC_279/A NOR2X1_LOC_139/Y 0.07fF
C62380 NAND2X1_LOC_357/B NOR2X1_LOC_322/a_36_216# 0.00fF
C62381 INPUT_1 NOR2X1_LOC_167/Y 0.00fF
C62382 NOR2X1_LOC_516/B INVX1_LOC_59/Y 0.29fF
C62383 NOR2X1_LOC_152/Y INVX1_LOC_291/A 0.09fF
C62384 INVX1_LOC_205/Y INVX1_LOC_15/A 0.01fF
C62385 NAND2X1_LOC_181/Y VDD 0.42fF
C62386 NAND2X1_LOC_850/Y INVX1_LOC_37/A 0.07fF
C62387 NOR2X1_LOC_546/B NAND2X1_LOC_425/Y 0.01fF
C62388 NOR2X1_LOC_226/A NAND2X1_LOC_84/a_36_24# 0.01fF
C62389 INVX1_LOC_53/Y INVX1_LOC_20/A 0.03fF
C62390 NOR2X1_LOC_160/B NOR2X1_LOC_340/A 0.12fF
C62391 NOR2X1_LOC_218/Y INVX1_LOC_76/A 0.01fF
C62392 NOR2X1_LOC_516/B INVX1_LOC_176/A 0.03fF
C62393 NOR2X1_LOC_52/B NOR2X1_LOC_271/Y 0.03fF
C62394 INVX1_LOC_1/A INVX1_LOC_32/A 0.29fF
C62395 NAND2X1_LOC_722/A NAND2X1_LOC_603/a_36_24# 0.01fF
C62396 INVX1_LOC_30/A NAND2X1_LOC_773/B 0.01fF
C62397 NOR2X1_LOC_384/Y NAND2X1_LOC_489/Y 0.02fF
C62398 INVX1_LOC_45/Y NAND2X1_LOC_606/a_36_24# 0.00fF
C62399 INVX1_LOC_299/A INVX1_LOC_15/A 0.03fF
C62400 INVX1_LOC_279/A NAND2X1_LOC_468/B 0.48fF
C62401 NOR2X1_LOC_301/A NOR2X1_LOC_652/Y 0.07fF
C62402 INVX1_LOC_1/A NOR2X1_LOC_623/B -0.01fF
C62403 NOR2X1_LOC_791/B INVX1_LOC_293/Y 0.00fF
C62404 INVX1_LOC_192/Y INVX1_LOC_38/A 0.39fF
C62405 INVX1_LOC_50/A NOR2X1_LOC_665/Y 0.00fF
C62406 NAND2X1_LOC_364/A NOR2X1_LOC_691/B 0.03fF
C62407 NOR2X1_LOC_724/Y NOR2X1_LOC_78/A -0.00fF
C62408 NOR2X1_LOC_537/Y INVX1_LOC_38/A 0.07fF
C62409 NAND2X1_LOC_664/a_36_24# INVX1_LOC_76/A 0.01fF
C62410 NAND2X1_LOC_338/B INVX1_LOC_38/A 0.07fF
C62411 NOR2X1_LOC_418/Y INVX1_LOC_77/Y 0.04fF
C62412 NAND2X1_LOC_593/Y NOR2X1_LOC_697/Y 0.02fF
C62413 NAND2X1_LOC_390/A VDD 0.15fF
C62414 NOR2X1_LOC_570/B NOR2X1_LOC_155/A 0.02fF
C62415 NAND2X1_LOC_621/a_36_24# NOR2X1_LOC_19/Y 0.00fF
C62416 NOR2X1_LOC_798/A NOR2X1_LOC_798/Y 0.01fF
C62417 NOR2X1_LOC_312/a_36_216# INVX1_LOC_54/A 0.02fF
C62418 INVX1_LOC_6/A NOR2X1_LOC_74/A 0.19fF
C62419 NAND2X1_LOC_505/a_36_24# INVX1_LOC_122/A 0.00fF
C62420 NOR2X1_LOC_348/B INVX1_LOC_307/A 0.12fF
C62421 INVX1_LOC_88/A INVX1_LOC_271/Y 0.02fF
C62422 INVX1_LOC_170/A NAND2X1_LOC_254/Y 0.02fF
C62423 NOR2X1_LOC_798/A NOR2X1_LOC_748/A 0.01fF
C62424 NOR2X1_LOC_419/a_36_216# NOR2X1_LOC_721/B 0.00fF
C62425 NOR2X1_LOC_329/B NOR2X1_LOC_405/A 0.02fF
C62426 INVX1_LOC_93/Y NAND2X1_LOC_850/A 0.02fF
C62427 INVX1_LOC_150/A INVX1_LOC_46/A 0.02fF
C62428 NAND2X1_LOC_361/Y NOR2X1_LOC_814/A 0.07fF
C62429 INVX1_LOC_83/A NOR2X1_LOC_319/a_36_216# 0.00fF
C62430 INVX1_LOC_6/A NOR2X1_LOC_9/Y 0.22fF
C62431 NAND2X1_LOC_648/A INVX1_LOC_76/A 0.03fF
C62432 NAND2X1_LOC_812/a_36_24# NAND2X1_LOC_770/Y 0.01fF
C62433 GATE_811 INVX1_LOC_297/A 0.26fF
C62434 INVX1_LOC_45/Y INVX1_LOC_29/A 0.03fF
C62435 NOR2X1_LOC_19/B INVX1_LOC_74/Y 0.01fF
C62436 NOR2X1_LOC_91/Y NOR2X1_LOC_89/A 0.03fF
C62437 INPUT_1 INVX1_LOC_76/A 0.11fF
C62438 NAND2X1_LOC_661/B INVX1_LOC_117/Y 0.33fF
C62439 INVX1_LOC_25/A INVX1_LOC_171/Y 0.01fF
C62440 INVX1_LOC_89/A INVX1_LOC_46/A 0.07fF
C62441 NOR2X1_LOC_144/Y NOR2X1_LOC_66/Y 0.04fF
C62442 NAND2X1_LOC_308/B NOR2X1_LOC_305/Y 0.02fF
C62443 NOR2X1_LOC_45/B INPUT_0 0.07fF
C62444 NOR2X1_LOC_359/Y NOR2X1_LOC_89/A 0.29fF
C62445 NAND2X1_LOC_7/Y INVX1_LOC_125/A 0.02fF
C62446 NAND2X1_LOC_847/a_36_24# NOR2X1_LOC_649/B 0.01fF
C62447 INVX1_LOC_182/Y NAND2X1_LOC_468/B 0.08fF
C62448 NAND2X1_LOC_656/Y NOR2X1_LOC_536/A 0.08fF
C62449 INVX1_LOC_30/A NOR2X1_LOC_393/Y 0.09fF
C62450 NOR2X1_LOC_315/Y INVX1_LOC_84/A 0.03fF
C62451 INVX1_LOC_35/A NOR2X1_LOC_272/Y 0.01fF
C62452 NOR2X1_LOC_577/Y INVX1_LOC_12/A 0.14fF
C62453 NOR2X1_LOC_561/Y INVX1_LOC_118/A 0.10fF
C62454 INVX1_LOC_230/Y INVX1_LOC_26/A 0.03fF
C62455 INVX1_LOC_22/A INVX1_LOC_307/A 0.08fF
C62456 NOR2X1_LOC_92/Y INVX1_LOC_308/A 0.03fF
C62457 INVX1_LOC_161/Y NOR2X1_LOC_106/a_36_216# 0.01fF
C62458 INVX1_LOC_232/A NOR2X1_LOC_216/B 0.09fF
C62459 INVX1_LOC_171/A NOR2X1_LOC_652/a_36_216# 0.00fF
C62460 NOR2X1_LOC_400/A INVX1_LOC_235/Y 0.01fF
C62461 NOR2X1_LOC_78/A NOR2X1_LOC_557/A 0.06fF
C62462 INVX1_LOC_17/A D_INPUT_1 0.03fF
C62463 INVX1_LOC_22/A NOR2X1_LOC_445/B 0.07fF
C62464 INVX1_LOC_268/A INVX1_LOC_107/Y 0.18fF
C62465 INVX1_LOC_25/A NOR2X1_LOC_296/Y 0.30fF
C62466 INVX1_LOC_17/Y NOR2X1_LOC_615/Y 0.24fF
C62467 INVX1_LOC_313/Y INVX1_LOC_38/A 0.07fF
C62468 NOR2X1_LOC_601/a_36_216# NOR2X1_LOC_15/Y 0.01fF
C62469 NOR2X1_LOC_590/A NOR2X1_LOC_113/a_36_216# 0.00fF
C62470 NOR2X1_LOC_383/Y NOR2X1_LOC_216/B 0.22fF
C62471 NAND2X1_LOC_656/Y NAND2X1_LOC_93/B 0.07fF
C62472 NAND2X1_LOC_773/Y NOR2X1_LOC_772/B 0.10fF
C62473 INVX1_LOC_18/A NOR2X1_LOC_36/A 0.02fF
C62474 NOR2X1_LOC_802/A NAND2X1_LOC_74/B 0.02fF
C62475 INVX1_LOC_58/A NOR2X1_LOC_369/Y 0.03fF
C62476 NOR2X1_LOC_589/Y VDD 0.24fF
C62477 NAND2X1_LOC_763/B NAND2X1_LOC_70/a_36_24# 0.01fF
C62478 INVX1_LOC_25/A INPUT_3 0.16fF
C62479 NOR2X1_LOC_78/A NOR2X1_LOC_657/B 0.08fF
C62480 INVX1_LOC_90/A NOR2X1_LOC_506/Y 0.18fF
C62481 NAND2X1_LOC_773/Y INVX1_LOC_13/Y 0.03fF
C62482 D_INPUT_1 NAND2X1_LOC_555/Y 0.08fF
C62483 NOR2X1_LOC_721/Y INVX1_LOC_117/A 0.02fF
C62484 NAND2X1_LOC_634/Y NOR2X1_LOC_693/Y 0.10fF
C62485 NOR2X1_LOC_789/A INVX1_LOC_3/A 0.01fF
C62486 INVX1_LOC_42/Y INVX1_LOC_10/Y 0.03fF
C62487 INVX1_LOC_58/A INVX1_LOC_286/Y 0.07fF
C62488 NOR2X1_LOC_647/A NOR2X1_LOC_68/A 0.01fF
C62489 INVX1_LOC_1/A INVX1_LOC_171/Y 0.03fF
C62490 INVX1_LOC_124/Y INVX1_LOC_23/A 0.09fF
C62491 NAND2X1_LOC_720/a_36_24# NOR2X1_LOC_654/A 0.04fF
C62492 NOR2X1_LOC_535/a_36_216# NOR2X1_LOC_640/Y 0.00fF
C62493 NOR2X1_LOC_669/Y NAND2X1_LOC_703/Y 0.01fF
C62494 NOR2X1_LOC_222/Y INVX1_LOC_109/Y 0.04fF
C62495 NOR2X1_LOC_315/Y INVX1_LOC_15/A 0.03fF
C62496 NAND2X1_LOC_623/B VDD 0.16fF
C62497 NOR2X1_LOC_646/A NAND2X1_LOC_74/B 0.00fF
C62498 NOR2X1_LOC_516/B NOR2X1_LOC_340/A 0.07fF
C62499 INVX1_LOC_176/A NAND2X1_LOC_109/a_36_24# 0.01fF
C62500 INVX1_LOC_35/A NOR2X1_LOC_336/B 0.00fF
C62501 INVX1_LOC_255/Y INVX1_LOC_29/A 0.07fF
C62502 INVX1_LOC_144/A INVX1_LOC_54/A 0.10fF
C62503 INVX1_LOC_22/A INVX1_LOC_12/A 0.70fF
C62504 INVX1_LOC_58/A INVX1_LOC_159/A 0.11fF
C62505 NOR2X1_LOC_314/Y NOR2X1_LOC_56/Y 0.01fF
C62506 NOR2X1_LOC_264/Y INVX1_LOC_87/A 1.24fF
C62507 NOR2X1_LOC_167/Y INVX1_LOC_118/A 0.03fF
C62508 INVX1_LOC_75/A INVX1_LOC_92/A 0.27fF
C62509 INVX1_LOC_135/A INVX1_LOC_19/A 0.09fF
C62510 INVX1_LOC_35/A NAND2X1_LOC_364/A 0.13fF
C62511 NAND2X1_LOC_149/Y INVX1_LOC_174/A 0.05fF
C62512 NAND2X1_LOC_787/A INVX1_LOC_24/A 0.07fF
C62513 NAND2X1_LOC_244/A INVX1_LOC_46/A 0.04fF
C62514 INPUT_0 NOR2X1_LOC_862/B 0.05fF
C62515 INVX1_LOC_36/A INVX1_LOC_306/Y 3.83fF
C62516 VDD NOR2X1_LOC_422/Y 0.34fF
C62517 NAND2X1_LOC_363/B INVX1_LOC_24/A 0.07fF
C62518 VDD NOR2X1_LOC_314/Y 0.34fF
C62519 NOR2X1_LOC_71/Y INVX1_LOC_29/A 0.07fF
C62520 INVX1_LOC_58/A INVX1_LOC_283/Y -0.01fF
C62521 INVX1_LOC_272/Y NAND2X1_LOC_799/A 0.47fF
C62522 NOR2X1_LOC_76/A NAND2X1_LOC_81/B 0.07fF
C62523 NAND2X1_LOC_338/B NAND2X1_LOC_223/A 0.07fF
C62524 NOR2X1_LOC_793/A INVX1_LOC_292/A 0.12fF
C62525 INPUT_2 INVX1_LOC_14/A 1.98fF
C62526 INPUT_3 INVX1_LOC_1/A 0.15fF
C62527 NOR2X1_LOC_68/A INVX1_LOC_298/A 0.01fF
C62528 INVX1_LOC_53/Y INVX1_LOC_4/A 0.50fF
C62529 INVX1_LOC_89/A NOR2X1_LOC_671/Y 0.03fF
C62530 INVX1_LOC_12/Y NOR2X1_LOC_137/Y 0.03fF
C62531 NOR2X1_LOC_302/Y INVX1_LOC_186/Y 0.02fF
C62532 INVX1_LOC_103/A NOR2X1_LOC_160/B 0.07fF
C62533 INVX1_LOC_224/Y NOR2X1_LOC_392/B 0.03fF
C62534 GATE_662 NOR2X1_LOC_467/A 0.02fF
C62535 NOR2X1_LOC_214/B NAND2X1_LOC_469/a_36_24# 0.01fF
C62536 NOR2X1_LOC_644/A INVX1_LOC_29/A 0.07fF
C62537 VDD INVX1_LOC_117/A 4.27fF
C62538 NAND2X1_LOC_573/A NAND2X1_LOC_404/a_36_24# 0.02fF
C62539 INVX1_LOC_236/Y NAND2X1_LOC_538/Y 0.04fF
C62540 INVX1_LOC_18/A NAND2X1_LOC_474/Y 0.02fF
C62541 NOR2X1_LOC_665/A INVX1_LOC_4/A 0.16fF
C62542 NOR2X1_LOC_824/Y INVX1_LOC_118/A 0.01fF
C62543 NOR2X1_LOC_791/Y INVX1_LOC_24/A 0.01fF
C62544 INVX1_LOC_245/A INVX1_LOC_78/A 0.01fF
C62545 INVX1_LOC_233/Y NAND2X1_LOC_833/Y 0.00fF
C62546 VDD NOR2X1_LOC_808/B 0.29fF
C62547 NOR2X1_LOC_226/A NOR2X1_LOC_447/A 0.03fF
C62548 INVX1_LOC_95/Y NOR2X1_LOC_99/Y 0.13fF
C62549 NOR2X1_LOC_577/a_36_216# NOR2X1_LOC_334/Y 0.00fF
C62550 INVX1_LOC_76/A INVX1_LOC_118/A 0.61fF
C62551 NOR2X1_LOC_632/Y INVX1_LOC_78/A 0.03fF
C62552 NAND2X1_LOC_734/B INVX1_LOC_53/A 0.03fF
C62553 INVX1_LOC_34/A NOR2X1_LOC_53/Y 0.12fF
C62554 NOR2X1_LOC_684/a_36_216# INVX1_LOC_117/A 0.01fF
C62555 INVX1_LOC_14/Y INVX1_LOC_9/A 0.10fF
C62556 INVX1_LOC_278/A NOR2X1_LOC_315/Y 0.28fF
C62557 INVX1_LOC_226/Y NOR2X1_LOC_843/B 0.03fF
C62558 NAND2X1_LOC_624/A INVX1_LOC_15/A 0.06fF
C62559 NOR2X1_LOC_205/Y NOR2X1_LOC_457/B 0.98fF
C62560 NAND2X1_LOC_579/A NAND2X1_LOC_837/Y 0.15fF
C62561 NAND2X1_LOC_53/Y INVX1_LOC_18/A 0.29fF
C62562 NAND2X1_LOC_510/a_36_24# INVX1_LOC_50/Y 0.00fF
C62563 INVX1_LOC_200/Y NOR2X1_LOC_488/Y 0.01fF
C62564 NOR2X1_LOC_91/A NAND2X1_LOC_660/Y 0.19fF
C62565 NAND2X1_LOC_485/a_36_24# INVX1_LOC_92/A 0.00fF
C62566 INVX1_LOC_239/A NOR2X1_LOC_474/A 0.10fF
C62567 NAND2X1_LOC_149/Y INVX1_LOC_153/A 0.06fF
C62568 NAND2X1_LOC_453/A INVX1_LOC_92/A 0.07fF
C62569 NAND2X1_LOC_773/Y INVX1_LOC_303/A 0.87fF
C62570 INVX1_LOC_233/A NOR2X1_LOC_401/B 0.05fF
C62571 NOR2X1_LOC_78/B NOR2X1_LOC_392/Y 0.01fF
C62572 INVX1_LOC_246/A NAND2X1_LOC_354/Y 0.18fF
C62573 INVX1_LOC_1/Y INVX1_LOC_57/A 0.22fF
C62574 NOR2X1_LOC_284/a_36_216# NOR2X1_LOC_598/B 0.01fF
C62575 NOR2X1_LOC_613/Y INVX1_LOC_34/A 0.03fF
C62576 NOR2X1_LOC_716/B NAND2X1_LOC_347/B 0.02fF
C62577 NAND2X1_LOC_112/Y INVX1_LOC_271/A 0.00fF
C62578 INVX1_LOC_230/A INVX1_LOC_9/A 0.07fF
C62579 INVX1_LOC_25/Y INVX1_LOC_53/A 0.00fF
C62580 INVX1_LOC_135/A INVX1_LOC_26/Y 0.03fF
C62581 NAND2X1_LOC_9/Y NOR2X1_LOC_618/a_36_216# 0.02fF
C62582 NOR2X1_LOC_426/a_36_216# INVX1_LOC_72/A 0.01fF
C62583 NOR2X1_LOC_91/A D_INPUT_0 0.12fF
C62584 NAND2X1_LOC_219/a_36_24# NOR2X1_LOC_643/Y 0.00fF
C62585 NAND2X1_LOC_660/Y INVX1_LOC_23/A 0.03fF
C62586 INVX1_LOC_24/Y NOR2X1_LOC_551/B 0.03fF
C62587 INVX1_LOC_73/Y NOR2X1_LOC_433/A 0.07fF
C62588 NOR2X1_LOC_552/A INVX1_LOC_19/A 0.05fF
C62589 NAND2X1_LOC_349/B INVX1_LOC_53/A 0.07fF
C62590 NOR2X1_LOC_446/A NOR2X1_LOC_303/Y 0.03fF
C62591 INVX1_LOC_21/A NOR2X1_LOC_84/Y 0.78fF
C62592 INVX1_LOC_64/A NOR2X1_LOC_219/Y 0.49fF
C62593 NOR2X1_LOC_454/Y NOR2X1_LOC_194/Y 0.03fF
C62594 NAND2X1_LOC_214/B NAND2X1_LOC_541/Y 0.02fF
C62595 INVX1_LOC_64/A INVX1_LOC_53/Y 0.13fF
C62596 NOR2X1_LOC_188/A INVX1_LOC_32/A 1.78fF
C62597 INVX1_LOC_166/A INVX1_LOC_135/A 1.11fF
C62598 NOR2X1_LOC_135/Y INVX1_LOC_78/A 0.10fF
C62599 NAND2X1_LOC_370/a_36_24# NAND2X1_LOC_564/B 0.00fF
C62600 NOR2X1_LOC_667/A NAND2X1_LOC_794/B 0.14fF
C62601 INVX1_LOC_276/A INVX1_LOC_178/A 0.01fF
C62602 INVX1_LOC_227/Y INVX1_LOC_223/A 0.01fF
C62603 INVX1_LOC_14/A INVX1_LOC_162/Y 0.07fF
C62604 NAND2X1_LOC_555/Y D_INPUT_2 0.19fF
C62605 NAND2X1_LOC_149/Y INVX1_LOC_259/A 0.06fF
C62606 NOR2X1_LOC_753/Y NOR2X1_LOC_816/A 0.03fF
C62607 NAND2X1_LOC_794/B INVX1_LOC_248/A 0.10fF
C62608 INVX1_LOC_143/A NAND2X1_LOC_63/a_36_24# 0.00fF
C62609 NOR2X1_LOC_67/A INVX1_LOC_178/A 0.10fF
C62610 D_INPUT_0 INVX1_LOC_23/A 1.38fF
C62611 INVX1_LOC_64/A NOR2X1_LOC_665/A 0.16fF
C62612 NOR2X1_LOC_411/A NAND2X1_LOC_462/B 0.08fF
C62613 INVX1_LOC_24/A INVX1_LOC_30/A 0.32fF
C62614 NAND2X1_LOC_468/B NAND2X1_LOC_433/a_36_24# 0.00fF
C62615 NOR2X1_LOC_540/B INVX1_LOC_29/A 0.00fF
C62616 NAND2X1_LOC_326/A INVX1_LOC_236/A 0.00fF
C62617 NOR2X1_LOC_691/B NOR2X1_LOC_857/A 0.01fF
C62618 INVX1_LOC_305/A NAND2X1_LOC_789/a_36_24# 0.02fF
C62619 NOR2X1_LOC_816/A NAND2X1_LOC_325/Y 0.07fF
C62620 NOR2X1_LOC_392/B NOR2X1_LOC_103/Y 0.10fF
C62621 INVX1_LOC_7/A INVX1_LOC_138/A 0.02fF
C62622 INVX1_LOC_256/A INVX1_LOC_88/Y 0.00fF
C62623 NAND2X1_LOC_733/Y NOR2X1_LOC_577/Y 0.23fF
C62624 NOR2X1_LOC_590/A NAND2X1_LOC_361/Y 0.08fF
C62625 NOR2X1_LOC_331/B NOR2X1_LOC_841/A 0.10fF
C62626 NAND2X1_LOC_741/Y NAND2X1_LOC_863/B 0.01fF
C62627 NOR2X1_LOC_155/A INVX1_LOC_54/A 0.06fF
C62628 NOR2X1_LOC_626/Y INVX1_LOC_16/A 0.03fF
C62629 VDD INVX1_LOC_163/Y 0.41fF
C62630 NOR2X1_LOC_9/Y NOR2X1_LOC_80/Y 0.16fF
C62631 INVX1_LOC_22/Y NAND2X1_LOC_361/Y 0.02fF
C62632 NAND2X1_LOC_9/Y INVX1_LOC_89/A 0.05fF
C62633 INVX1_LOC_39/A NOR2X1_LOC_719/A 0.01fF
C62634 INVX1_LOC_152/A NOR2X1_LOC_61/A 0.05fF
C62635 NAND2X1_LOC_557/Y NOR2X1_LOC_490/Y 0.07fF
C62636 INVX1_LOC_2/Y NAND2X1_LOC_74/B 0.00fF
C62637 INVX1_LOC_21/A INVX1_LOC_290/A 0.03fF
C62638 NOR2X1_LOC_43/Y INVX1_LOC_32/A 0.06fF
C62639 INVX1_LOC_45/A NOR2X1_LOC_172/Y 0.03fF
C62640 INVX1_LOC_13/A NAND2X1_LOC_141/a_36_24# 0.00fF
C62641 NOR2X1_LOC_292/Y INVX1_LOC_26/A 0.38fF
C62642 INVX1_LOC_90/A NAND2X1_LOC_793/B 0.08fF
C62643 NOR2X1_LOC_361/B NAND2X1_LOC_181/Y 0.03fF
C62644 INVX1_LOC_256/A NOR2X1_LOC_168/B 0.10fF
C62645 NOR2X1_LOC_813/Y INVX1_LOC_19/A 0.07fF
C62646 NOR2X1_LOC_557/Y INVX1_LOC_30/A 0.05fF
C62647 INVX1_LOC_103/A NAND2X1_LOC_350/B 0.00fF
C62648 INVX1_LOC_45/A NOR2X1_LOC_147/B 0.05fF
C62649 NAND2X1_LOC_149/Y NOR2X1_LOC_589/A 0.09fF
C62650 INVX1_LOC_39/A INVX1_LOC_7/A 0.06fF
C62651 INVX1_LOC_33/A INVX1_LOC_72/A 0.22fF
C62652 INVX1_LOC_50/A INVX1_LOC_67/Y 0.00fF
C62653 INVX1_LOC_278/A NOR2X1_LOC_166/Y 0.06fF
C62654 INVX1_LOC_235/Y NAND2X1_LOC_377/Y 0.01fF
C62655 INVX1_LOC_276/A NOR2X1_LOC_816/A 0.27fF
C62656 NOR2X1_LOC_178/Y INPUT_1 0.07fF
C62657 NAND2X1_LOC_659/B INVX1_LOC_3/Y 0.00fF
C62658 NOR2X1_LOC_74/A INVX1_LOC_270/A 0.01fF
C62659 INVX1_LOC_45/A NOR2X1_LOC_392/B 0.03fF
C62660 NAND2X1_LOC_553/A INVX1_LOC_89/A 0.00fF
C62661 NOR2X1_LOC_439/B INVX1_LOC_53/A 0.03fF
C62662 INVX1_LOC_103/A INVX1_LOC_208/A 0.01fF
C62663 INVX1_LOC_91/A INVX1_LOC_273/A 0.10fF
C62664 INVX1_LOC_36/A INVX1_LOC_294/Y 0.00fF
C62665 INVX1_LOC_34/A NOR2X1_LOC_52/Y 0.00fF
C62666 INVX1_LOC_280/A INVX1_LOC_19/A 0.14fF
C62667 VDD NOR2X1_LOC_460/A 0.00fF
C62668 NOR2X1_LOC_592/B NOR2X1_LOC_841/A 0.18fF
C62669 INVX1_LOC_163/A NAND2X1_LOC_462/B 0.01fF
C62670 INVX1_LOC_1/A GATE_662 0.03fF
C62671 NOR2X1_LOC_703/A INVX1_LOC_292/Y 0.11fF
C62672 INVX1_LOC_75/A INVX1_LOC_53/A 0.33fF
C62673 INVX1_LOC_274/A INVX1_LOC_63/A 0.08fF
C62674 NOR2X1_LOC_798/A INVX1_LOC_89/A 0.07fF
C62675 NOR2X1_LOC_82/A INVX1_LOC_316/Y 0.16fF
C62676 INVX1_LOC_33/A INVX1_LOC_198/Y 0.02fF
C62677 NAND2X1_LOC_656/Y NOR2X1_LOC_348/Y 0.00fF
C62678 INVX1_LOC_132/A INVX1_LOC_314/Y 0.09fF
C62679 NOR2X1_LOC_827/a_36_216# NOR2X1_LOC_500/B 0.05fF
C62680 VDD INVX1_LOC_3/Y 3.60fF
C62681 NOR2X1_LOC_562/a_36_216# NOR2X1_LOC_303/Y 0.00fF
C62682 NOR2X1_LOC_172/Y INVX1_LOC_71/A 0.03fF
C62683 INVX1_LOC_208/A INVX1_LOC_292/A 0.01fF
C62684 INVX1_LOC_279/A INVX1_LOC_88/A 0.07fF
C62685 NAND2X1_LOC_579/A NOR2X1_LOC_299/Y 0.02fF
C62686 INVX1_LOC_223/A INVX1_LOC_111/Y 0.02fF
C62687 INVX1_LOC_45/A NAND2X1_LOC_294/a_36_24# 0.00fF
C62688 INVX1_LOC_143/A INVX1_LOC_30/A 0.02fF
C62689 NOR2X1_LOC_52/B NOR2X1_LOC_91/Y 2.72fF
C62690 INVX1_LOC_43/Y INVX1_LOC_53/Y 0.00fF
C62691 INVX1_LOC_292/A NOR2X1_LOC_516/B 0.07fF
C62692 NOR2X1_LOC_448/B INVX1_LOC_83/A 0.03fF
C62693 INVX1_LOC_64/A NAND2X1_LOC_124/a_36_24# 0.00fF
C62694 INVX1_LOC_136/A NOR2X1_LOC_767/a_36_216# 0.01fF
C62695 INVX1_LOC_134/A INVX1_LOC_160/Y 0.11fF
C62696 NOR2X1_LOC_392/B INVX1_LOC_71/A 0.17fF
C62697 NOR2X1_LOC_74/A NOR2X1_LOC_109/Y 0.01fF
C62698 NOR2X1_LOC_820/Y INVX1_LOC_63/A 0.31fF
C62699 NOR2X1_LOC_861/Y INVX1_LOC_230/A 0.12fF
C62700 NOR2X1_LOC_318/B INVX1_LOC_57/A 0.01fF
C62701 NOR2X1_LOC_15/Y INVX1_LOC_183/Y 0.01fF
C62702 NAND2X1_LOC_96/A INVX1_LOC_15/A 0.07fF
C62703 NAND2X1_LOC_733/Y INVX1_LOC_22/A 0.03fF
C62704 NOR2X1_LOC_78/A INVX1_LOC_271/A 0.03fF
C62705 INVX1_LOC_256/A NAND2X1_LOC_656/Y 0.10fF
C62706 NOR2X1_LOC_640/Y INVX1_LOC_69/A 0.06fF
C62707 INVX1_LOC_41/A NOR2X1_LOC_551/B 0.03fF
C62708 INVX1_LOC_24/A NAND2X1_LOC_722/A 0.02fF
C62709 INVX1_LOC_76/A NOR2X1_LOC_631/Y 0.11fF
C62710 INVX1_LOC_135/A INVX1_LOC_161/Y 0.03fF
C62711 INVX1_LOC_93/Y INVX1_LOC_57/A 0.15fF
C62712 NAND2X1_LOC_726/Y INVX1_LOC_72/A 0.00fF
C62713 NAND2X1_LOC_198/B NAND2X1_LOC_850/Y 0.10fF
C62714 NOR2X1_LOC_655/B INVX1_LOC_94/A 0.10fF
C62715 INVX1_LOC_18/A NOR2X1_LOC_500/Y 0.03fF
C62716 NOR2X1_LOC_246/A NAND2X1_LOC_807/A 0.03fF
C62717 INVX1_LOC_90/A NOR2X1_LOC_103/Y 0.00fF
C62718 INVX1_LOC_41/A INVX1_LOC_213/Y 0.07fF
C62719 NOR2X1_LOC_2/Y D_INPUT_6 0.03fF
C62720 NOR2X1_LOC_155/A NAND2X1_LOC_807/B 0.03fF
C62721 INVX1_LOC_104/A INVX1_LOC_155/Y 0.03fF
C62722 INVX1_LOC_217/A INVX1_LOC_22/A 0.05fF
C62723 INVX1_LOC_58/A NOR2X1_LOC_56/Y 0.03fF
C62724 NOR2X1_LOC_160/B INVX1_LOC_120/A 0.01fF
C62725 INVX1_LOC_128/A NOR2X1_LOC_331/B -0.10fF
C62726 INVX1_LOC_35/A NOR2X1_LOC_113/A 0.01fF
C62727 INVX1_LOC_294/Y NOR2X1_LOC_309/Y 0.04fF
C62728 INVX1_LOC_224/Y NOR2X1_LOC_92/a_36_216# 0.01fF
C62729 D_INPUT_0 INVX1_LOC_31/A 0.31fF
C62730 INVX1_LOC_283/A INVX1_LOC_92/A 0.03fF
C62731 INVX1_LOC_88/A INVX1_LOC_182/Y 0.02fF
C62732 INVX1_LOC_35/A NOR2X1_LOC_405/A 0.53fF
C62733 NAND2X1_LOC_287/B NAND2X1_LOC_285/a_36_24# 0.01fF
C62734 NOR2X1_LOC_189/A NOR2X1_LOC_667/A 0.44fF
C62735 INVX1_LOC_50/A NOR2X1_LOC_562/A 0.07fF
C62736 NAND2X1_LOC_190/a_36_24# NOR2X1_LOC_337/Y 0.01fF
C62737 NOR2X1_LOC_778/B NOR2X1_LOC_374/A 0.02fF
C62738 INVX1_LOC_214/Y NOR2X1_LOC_577/Y 0.00fF
C62739 INVX1_LOC_299/A NOR2X1_LOC_310/a_36_216# 0.01fF
C62740 NOR2X1_LOC_773/Y NOR2X1_LOC_753/Y 0.07fF
C62741 NAND2X1_LOC_214/B NOR2X1_LOC_78/A 0.09fF
C62742 INVX1_LOC_27/A NOR2X1_LOC_737/a_36_216# 0.01fF
C62743 NOR2X1_LOC_320/Y NAND2X1_LOC_326/A 0.08fF
C62744 NAND2X1_LOC_338/B INVX1_LOC_33/A 0.04fF
C62745 INVX1_LOC_30/A NOR2X1_LOC_130/A 0.10fF
C62746 INVX1_LOC_58/A INVX1_LOC_146/Y 0.01fF
C62747 INVX1_LOC_18/A INVX1_LOC_10/A 0.07fF
C62748 INVX1_LOC_255/Y INVX1_LOC_228/A 0.04fF
C62749 NOR2X1_LOC_92/Y NOR2X1_LOC_387/A 0.01fF
C62750 INVX1_LOC_58/A VDD 4.62fF
C62751 INVX1_LOC_223/A NOR2X1_LOC_137/A 0.44fF
C62752 NOR2X1_LOC_266/B INVX1_LOC_23/A 0.03fF
C62753 NAND2X1_LOC_721/A INVX1_LOC_57/A 0.06fF
C62754 NAND2X1_LOC_728/Y INVX1_LOC_10/A 0.07fF
C62755 NAND2X1_LOC_323/B INVX1_LOC_33/A 1.10fF
C62756 NAND2X1_LOC_796/B NOR2X1_LOC_528/Y 0.01fF
C62757 INVX1_LOC_27/A INVX1_LOC_98/A 0.12fF
C62758 NOR2X1_LOC_814/A NAND2X1_LOC_20/a_36_24# 0.01fF
C62759 NOR2X1_LOC_91/A NAND2X1_LOC_848/A 0.03fF
C62760 INVX1_LOC_58/A NAND2X1_LOC_800/A 0.12fF
C62761 NOR2X1_LOC_773/Y NAND2X1_LOC_325/Y 0.01fF
C62762 NAND2X1_LOC_785/Y NOR2X1_LOC_482/Y 0.02fF
C62763 INVX1_LOC_45/A INVX1_LOC_90/A 1.02fF
C62764 INVX1_LOC_53/A NAND2X1_LOC_453/A 0.36fF
C62765 NAND2X1_LOC_833/Y NAND2X1_LOC_862/A 0.00fF
C62766 NAND2X1_LOC_634/Y NOR2X1_LOC_71/Y 0.03fF
C62767 INVX1_LOC_208/A INVX1_LOC_67/A 0.02fF
C62768 INVX1_LOC_235/Y INVX1_LOC_167/Y 0.16fF
C62769 INVX1_LOC_245/A INVX1_LOC_113/Y 0.01fF
C62770 INVX1_LOC_27/A NOR2X1_LOC_78/A 0.33fF
C62771 INVX1_LOC_90/A NOR2X1_LOC_568/A 1.49fF
C62772 INVX1_LOC_22/A NAND2X1_LOC_787/B 0.05fF
C62773 INVX1_LOC_12/A INVX1_LOC_186/Y 0.07fF
C62774 INVX1_LOC_286/Y NOR2X1_LOC_533/a_36_216# 0.00fF
C62775 INVX1_LOC_45/A NOR2X1_LOC_389/B 0.07fF
C62776 INPUT_6 INVX1_LOC_37/A 0.01fF
C62777 INVX1_LOC_271/A NOR2X1_LOC_60/Y 0.01fF
C62778 NOR2X1_LOC_15/Y NOR2X1_LOC_114/A 0.01fF
C62779 INVX1_LOC_35/A NOR2X1_LOC_857/A 0.30fF
C62780 NAND2X1_LOC_711/B INVX1_LOC_10/A 0.07fF
C62781 NOR2X1_LOC_323/a_36_216# INVX1_LOC_57/A 0.00fF
C62782 NOR2X1_LOC_632/Y INVX1_LOC_113/Y 0.00fF
C62783 NOR2X1_LOC_637/Y INVX1_LOC_10/A 0.00fF
C62784 NOR2X1_LOC_389/B NOR2X1_LOC_568/A 0.00fF
C62785 NAND2X1_LOC_350/A INVX1_LOC_144/A 0.13fF
C62786 NAND2X1_LOC_487/a_36_24# INVX1_LOC_87/A 0.00fF
C62787 NAND2X1_LOC_454/Y NAND2X1_LOC_798/B 0.01fF
C62788 INVX1_LOC_255/Y NOR2X1_LOC_516/a_36_216# 0.00fF
C62789 INVX1_LOC_247/Y NOR2X1_LOC_644/A 0.04fF
C62790 NOR2X1_LOC_15/Y INVX1_LOC_91/A 0.15fF
C62791 NAND2X1_LOC_276/Y INVX1_LOC_30/Y 0.02fF
C62792 NOR2X1_LOC_570/B NOR2X1_LOC_570/A 0.03fF
C62793 INVX1_LOC_245/Y INVX1_LOC_6/A 0.16fF
C62794 NOR2X1_LOC_272/a_36_216# INVX1_LOC_76/A 0.01fF
C62795 NOR2X1_LOC_441/Y INVX1_LOC_144/A 0.03fF
C62796 INVX1_LOC_248/Y VDD 0.24fF
C62797 INPUT_3 NOR2X1_LOC_548/B 0.04fF
C62798 NOR2X1_LOC_536/A NOR2X1_LOC_717/A 0.07fF
C62799 INVX1_LOC_39/A INVX1_LOC_76/A 0.02fF
C62800 INVX1_LOC_45/A NAND2X1_LOC_348/A 0.01fF
C62801 INVX1_LOC_18/A NOR2X1_LOC_302/Y 0.01fF
C62802 NOR2X1_LOC_355/a_36_216# INVX1_LOC_71/A 0.00fF
C62803 INVX1_LOC_90/A INVX1_LOC_71/A 0.07fF
C62804 INVX1_LOC_293/A INVX1_LOC_123/A 0.00fF
C62805 NAND2X1_LOC_301/a_36_24# NAND2X1_LOC_841/A 0.00fF
C62806 NAND2X1_LOC_740/B NAND2X1_LOC_854/a_36_24# 0.01fF
C62807 NOR2X1_LOC_15/Y INVX1_LOC_11/Y 0.07fF
C62808 NOR2X1_LOC_189/A NAND2X1_LOC_804/a_36_24# 0.00fF
C62809 INVX1_LOC_38/A NAND2X1_LOC_793/B 0.02fF
C62810 INVX1_LOC_35/Y INVX1_LOC_23/Y 0.01fF
C62811 NAND2X1_LOC_338/B INVX1_LOC_40/A 0.10fF
C62812 NOR2X1_LOC_793/A NOR2X1_LOC_542/B 0.00fF
C62813 INVX1_LOC_95/Y NOR2X1_LOC_271/B 0.03fF
C62814 INVX1_LOC_226/Y INVX1_LOC_34/Y 0.02fF
C62815 INVX1_LOC_234/A NAND2X1_LOC_139/A 0.06fF
C62816 NOR2X1_LOC_389/B INVX1_LOC_71/A 0.10fF
C62817 NOR2X1_LOC_780/B NAND2X1_LOC_697/a_36_24# 0.00fF
C62818 NOR2X1_LOC_828/Y NOR2X1_LOC_729/A 0.08fF
C62819 NAND2X1_LOC_166/a_36_24# INVX1_LOC_75/A 0.00fF
C62820 INVX1_LOC_54/Y INVX1_LOC_232/A 0.00fF
C62821 INVX1_LOC_36/A NOR2X1_LOC_74/A 0.25fF
C62822 NAND2X1_LOC_338/B INVX1_LOC_165/Y 0.04fF
C62823 NOR2X1_LOC_502/Y NOR2X1_LOC_349/A 0.04fF
C62824 INVX1_LOC_124/Y INVX1_LOC_6/A 0.12fF
C62825 NOR2X1_LOC_78/B INVX1_LOC_25/Y 1.01fF
C62826 INVX1_LOC_190/A NAND2X1_LOC_466/Y 0.08fF
C62827 NOR2X1_LOC_724/Y NOR2X1_LOC_374/A 0.01fF
C62828 NOR2X1_LOC_267/A NOR2X1_LOC_74/A 0.10fF
C62829 NOR2X1_LOC_71/Y INVX1_LOC_8/A 0.93fF
C62830 NAND2X1_LOC_731/Y NAND2X1_LOC_863/A 0.10fF
C62831 INVX1_LOC_36/A NOR2X1_LOC_9/Y 0.22fF
C62832 NOR2X1_LOC_78/B NAND2X1_LOC_349/B 0.02fF
C62833 INVX1_LOC_33/A INVX1_LOC_313/Y 0.07fF
C62834 NAND2X1_LOC_850/a_36_24# NAND2X1_LOC_842/B 0.00fF
C62835 NAND2X1_LOC_500/Y NOR2X1_LOC_526/a_36_216# 0.00fF
C62836 NOR2X1_LOC_479/B INVX1_LOC_172/Y 0.11fF
C62837 NOR2X1_LOC_566/Y INVX1_LOC_22/A 0.01fF
C62838 NOR2X1_LOC_389/A NOR2X1_LOC_139/Y 0.02fF
C62839 NOR2X1_LOC_135/Y NOR2X1_LOC_152/Y 0.03fF
C62840 NAND2X1_LOC_48/a_36_24# NOR2X1_LOC_196/Y 0.00fF
C62841 NOR2X1_LOC_142/Y NOR2X1_LOC_768/a_36_216# 0.01fF
C62842 NOR2X1_LOC_178/Y INVX1_LOC_118/A 0.34fF
C62843 INVX1_LOC_45/A NAND2X1_LOC_123/a_36_24# 0.00fF
C62844 NOR2X1_LOC_662/A INVX1_LOC_175/A 0.14fF
C62845 NAND2X1_LOC_725/A INVX1_LOC_54/A 0.10fF
C62846 NAND2X1_LOC_93/B NOR2X1_LOC_717/A 0.07fF
C62847 INVX1_LOC_84/A NAND2X1_LOC_99/A 0.07fF
C62848 NOR2X1_LOC_209/B INVX1_LOC_213/A 0.04fF
C62849 NOR2X1_LOC_15/Y NOR2X1_LOC_290/a_36_216# 0.00fF
C62850 NOR2X1_LOC_753/Y INVX1_LOC_140/A 0.30fF
C62851 NAND2X1_LOC_717/Y INVX1_LOC_229/Y 0.15fF
C62852 D_GATE_222 INVX1_LOC_22/A -0.00fF
C62853 NOR2X1_LOC_160/B NOR2X1_LOC_542/B 0.02fF
C62854 D_INPUT_0 NOR2X1_LOC_290/Y 0.07fF
C62855 INVX1_LOC_103/A NAND2X1_LOC_211/Y 0.07fF
C62856 INVX1_LOC_50/A INVX1_LOC_285/A 0.09fF
C62857 NOR2X1_LOC_208/Y NOR2X1_LOC_74/A 0.07fF
C62858 INVX1_LOC_50/A INVX1_LOC_265/Y 0.03fF
C62859 NAND2X1_LOC_181/Y NAND2X1_LOC_573/A 0.01fF
C62860 NOR2X1_LOC_389/A NAND2X1_LOC_468/B 0.01fF
C62861 NAND2X1_LOC_139/A NOR2X1_LOC_19/B 0.01fF
C62862 NOR2X1_LOC_541/B INVX1_LOC_19/A 0.02fF
C62863 INVX1_LOC_50/A NOR2X1_LOC_814/A 0.07fF
C62864 INVX1_LOC_16/A NAND2X1_LOC_666/a_36_24# 0.00fF
C62865 NOR2X1_LOC_160/B INVX1_LOC_143/Y 0.01fF
C62866 NAND2X1_LOC_243/Y NOR2X1_LOC_291/a_36_216# 0.00fF
C62867 NOR2X1_LOC_738/Y VDD 0.26fF
C62868 INVX1_LOC_25/Y NAND2X1_LOC_392/Y 0.00fF
C62869 NOR2X1_LOC_655/Y NOR2X1_LOC_649/Y 0.14fF
C62870 NOR2X1_LOC_619/A NOR2X1_LOC_721/a_36_216# 0.00fF
C62871 NAND2X1_LOC_508/a_36_24# NOR2X1_LOC_349/A 0.00fF
C62872 INVX1_LOC_215/Y VDD 0.49fF
C62873 NOR2X1_LOC_804/B NOR2X1_LOC_74/A 0.20fF
C62874 NOR2X1_LOC_209/Y NOR2X1_LOC_724/Y 0.05fF
C62875 NOR2X1_LOC_160/B NOR2X1_LOC_137/Y 0.03fF
C62876 NOR2X1_LOC_298/Y NAND2X1_LOC_863/B 1.96fF
C62877 NOR2X1_LOC_599/Y INVX1_LOC_46/A 0.49fF
C62878 NOR2X1_LOC_751/A INVX1_LOC_8/A 0.16fF
C62879 NOR2X1_LOC_500/A INVX1_LOC_186/A 0.07fF
C62880 INVX1_LOC_265/A INPUT_0 0.03fF
C62881 INVX1_LOC_18/A NOR2X1_LOC_799/B 0.02fF
C62882 NOR2X1_LOC_690/Y INVX1_LOC_10/A 0.03fF
C62883 NOR2X1_LOC_516/B INVX1_LOC_120/A 0.03fF
C62884 NOR2X1_LOC_309/Y NOR2X1_LOC_74/A 0.10fF
C62885 INVX1_LOC_171/A INVX1_LOC_16/A 0.02fF
C62886 NOR2X1_LOC_276/Y NOR2X1_LOC_363/Y 0.20fF
C62887 D_INPUT_0 NAND2X1_LOC_859/Y 0.00fF
C62888 INVX1_LOC_132/A NOR2X1_LOC_557/A 0.81fF
C62889 NOR2X1_LOC_78/B NOR2X1_LOC_439/B 0.02fF
C62890 NAND2X1_LOC_36/a_36_24# NAND2X1_LOC_1/Y 0.00fF
C62891 NOR2X1_LOC_309/Y NOR2X1_LOC_9/Y 0.03fF
C62892 INVX1_LOC_314/Y NAND2X1_LOC_642/Y 0.12fF
C62893 NOR2X1_LOC_649/B NOR2X1_LOC_649/Y 0.16fF
C62894 INVX1_LOC_136/A INVX1_LOC_2/Y 0.00fF
C62895 NAND2X1_LOC_739/B NAND2X1_LOC_800/a_36_24# 0.00fF
C62896 NOR2X1_LOC_78/B INVX1_LOC_75/A 0.49fF
C62897 INVX1_LOC_142/A INVX1_LOC_37/A 0.00fF
C62898 INVX1_LOC_17/A NOR2X1_LOC_61/Y 0.36fF
C62899 INVX1_LOC_31/A NAND2X1_LOC_848/A 0.08fF
C62900 NOR2X1_LOC_410/Y INVX1_LOC_37/A 0.02fF
C62901 NOR2X1_LOC_303/Y NAND2X1_LOC_447/Y 0.10fF
C62902 NOR2X1_LOC_744/Y INVX1_LOC_20/A 0.01fF
C62903 NOR2X1_LOC_620/Y INVX1_LOC_65/A 0.46fF
C62904 INVX1_LOC_306/Y INVX1_LOC_63/A 0.08fF
C62905 NOR2X1_LOC_338/Y VDD 0.00fF
C62906 NOR2X1_LOC_392/Y NOR2X1_LOC_671/Y 0.01fF
C62907 INVX1_LOC_35/A NOR2X1_LOC_841/a_36_216# 0.00fF
C62908 INVX1_LOC_36/A NOR2X1_LOC_690/a_36_216# 0.02fF
C62909 NOR2X1_LOC_589/A INVX1_LOC_28/A 0.07fF
C62910 NOR2X1_LOC_168/B INVX1_LOC_69/Y 0.08fF
C62911 INVX1_LOC_269/A NOR2X1_LOC_831/B 0.01fF
C62912 NOR2X1_LOC_664/Y NOR2X1_LOC_78/A 0.01fF
C62913 D_INPUT_0 INVX1_LOC_313/A 0.02fF
C62914 INVX1_LOC_45/A INVX1_LOC_38/A 4.05fF
C62915 INVX1_LOC_41/Y INVX1_LOC_37/A 0.03fF
C62916 INVX1_LOC_90/A NOR2X1_LOC_123/B 1.01fF
C62917 NOR2X1_LOC_568/A INVX1_LOC_38/A 0.07fF
C62918 INVX1_LOC_62/A NOR2X1_LOC_560/A 0.02fF
C62919 NOR2X1_LOC_669/Y INVX1_LOC_119/Y 0.04fF
C62920 NOR2X1_LOC_45/B INVX1_LOC_266/Y 0.09fF
C62921 INVX1_LOC_89/A NOR2X1_LOC_702/a_36_216# 0.00fF
C62922 INVX1_LOC_290/A NAND2X1_LOC_51/B 0.44fF
C62923 NOR2X1_LOC_763/Y NAND2X1_LOC_654/B 0.01fF
C62924 INVX1_LOC_90/A NOR2X1_LOC_749/Y 0.01fF
C62925 NOR2X1_LOC_496/Y NAND2X1_LOC_500/B 0.18fF
C62926 D_INPUT_0 NAND2X1_LOC_807/Y 0.07fF
C62927 NAND2X1_LOC_593/Y INVX1_LOC_37/A 0.07fF
C62928 NAND2X1_LOC_39/Y INVX1_LOC_113/Y 0.16fF
C62929 NAND2X1_LOC_53/Y NAND2X1_LOC_210/a_36_24# 0.00fF
C62930 INVX1_LOC_96/A NOR2X1_LOC_352/Y 0.01fF
C62931 NOR2X1_LOC_15/Y INVX1_LOC_203/A 0.18fF
C62932 NOR2X1_LOC_318/A NOR2X1_LOC_301/A 0.68fF
C62933 NAND2X1_LOC_725/A NOR2X1_LOC_48/B 0.20fF
C62934 INVX1_LOC_67/A NAND2X1_LOC_211/Y 0.10fF
C62935 INVX1_LOC_31/A INVX1_LOC_46/Y 0.02fF
C62936 NAND2X1_LOC_338/B NAND2X1_LOC_490/a_36_24# 0.01fF
C62937 INVX1_LOC_304/A NOR2X1_LOC_84/Y 0.12fF
C62938 NOR2X1_LOC_441/Y NOR2X1_LOC_155/A 0.03fF
C62939 NOR2X1_LOC_658/Y NAND2X1_LOC_93/B 0.07fF
C62940 NOR2X1_LOC_13/Y NOR2X1_LOC_536/A 0.17fF
C62941 INVX1_LOC_57/A INVX1_LOC_87/A 0.14fF
C62942 INVX1_LOC_21/A NOR2X1_LOC_641/a_36_216# 0.00fF
C62943 NOR2X1_LOC_242/A NAND2X1_LOC_291/B 0.03fF
C62944 INVX1_LOC_83/A INVX1_LOC_75/A 0.28fF
C62945 D_INPUT_1 INVX1_LOC_94/Y 0.03fF
C62946 NAND2X1_LOC_736/Y INVX1_LOC_46/A 0.08fF
C62947 NAND2X1_LOC_840/B INVX1_LOC_91/A 0.07fF
C62948 NAND2X1_LOC_660/Y INVX1_LOC_6/A 0.22fF
C62949 INVX1_LOC_71/A INVX1_LOC_38/A 0.07fF
C62950 NAND2X1_LOC_634/Y NAND2X1_LOC_243/Y 0.02fF
C62951 INVX1_LOC_54/Y NAND2X1_LOC_447/Y 0.03fF
C62952 NAND2X1_LOC_471/a_36_24# NAND2X1_LOC_464/A 0.01fF
C62953 NAND2X1_LOC_784/A NAND2X1_LOC_175/Y 0.03fF
C62954 INVX1_LOC_30/A NOR2X1_LOC_197/B 0.04fF
C62955 INVX1_LOC_153/Y INVX1_LOC_117/A 0.10fF
C62956 NOR2X1_LOC_106/Y INVX1_LOC_9/A 0.02fF
C62957 NOR2X1_LOC_299/Y NOR2X1_LOC_387/A 0.03fF
C62958 INVX1_LOC_18/A INVX1_LOC_307/A 0.07fF
C62959 NOR2X1_LOC_536/Y INVX1_LOC_12/A 0.01fF
C62960 NAND2X1_LOC_717/Y INVX1_LOC_20/A 0.01fF
C62961 NAND2X1_LOC_629/Y INVX1_LOC_14/Y 0.00fF
C62962 INVX1_LOC_41/Y NOR2X1_LOC_177/Y 0.01fF
C62963 NOR2X1_LOC_68/A NAND2X1_LOC_798/B 0.07fF
C62964 D_INPUT_0 INVX1_LOC_6/A 0.06fF
C62965 INVX1_LOC_110/Y NAND2X1_LOC_206/Y 0.09fF
C62966 INVX1_LOC_73/A NAND2X1_LOC_830/a_36_24# 0.01fF
C62967 NOR2X1_LOC_513/a_36_216# INVX1_LOC_54/A 0.02fF
C62968 NAND2X1_LOC_860/A INVX1_LOC_23/Y 0.03fF
C62969 NOR2X1_LOC_172/Y NOR2X1_LOC_331/B 0.04fF
C62970 INVX1_LOC_221/Y INVX1_LOC_49/Y 0.01fF
C62971 INVX1_LOC_18/A NOR2X1_LOC_445/B 0.07fF
C62972 INVX1_LOC_121/Y INVX1_LOC_117/A 0.03fF
C62973 NAND2X1_LOC_577/A INVX1_LOC_84/A 0.07fF
C62974 INVX1_LOC_21/A NOR2X1_LOC_467/A 0.08fF
C62975 INVX1_LOC_13/Y NOR2X1_LOC_38/B 0.25fF
C62976 INVX1_LOC_25/Y NOR2X1_LOC_368/Y 0.02fF
C62977 INVX1_LOC_316/Y INVX1_LOC_59/Y 0.75fF
C62978 NOR2X1_LOC_773/Y NOR2X1_LOC_558/A 0.00fF
C62979 INVX1_LOC_278/A NAND2X1_LOC_99/A 0.01fF
C62980 INVX1_LOC_177/A INVX1_LOC_117/A 0.04fF
C62981 NOR2X1_LOC_845/A NOR2X1_LOC_99/B 0.04fF
C62982 INVX1_LOC_266/Y INVX1_LOC_281/A 0.00fF
C62983 NAND2X1_LOC_338/B NAND2X1_LOC_642/a_36_24# 0.00fF
C62984 NOR2X1_LOC_446/a_36_216# INVX1_LOC_29/A 0.00fF
C62985 INVX1_LOC_303/A NOR2X1_LOC_624/B 0.04fF
C62986 INVX1_LOC_16/A INVX1_LOC_20/A 1.30fF
C62987 NOR2X1_LOC_537/a_36_216# NOR2X1_LOC_537/Y 0.02fF
C62988 NOR2X1_LOC_464/B INVX1_LOC_15/A 0.01fF
C62989 NOR2X1_LOC_577/Y INVX1_LOC_92/A 0.15fF
C62990 NOR2X1_LOC_375/Y D_GATE_479 0.01fF
C62991 NAND2X1_LOC_114/B NOR2X1_LOC_89/A 0.06fF
C62992 NOR2X1_LOC_290/Y NAND2X1_LOC_848/A 0.01fF
C62993 INVX1_LOC_25/Y INVX1_LOC_46/A 0.12fF
C62994 NOR2X1_LOC_15/Y INVX1_LOC_231/A 0.03fF
C62995 NOR2X1_LOC_361/B INVX1_LOC_3/Y 0.15fF
C62996 INVX1_LOC_163/A NAND2X1_LOC_618/Y 0.04fF
C62997 D_INPUT_6 NOR2X1_LOC_36/A 0.14fF
C62998 NOR2X1_LOC_473/B NOR2X1_LOC_269/Y 0.00fF
C62999 NAND2X1_LOC_349/B INVX1_LOC_46/A 0.07fF
C63000 NOR2X1_LOC_758/Y NOR2X1_LOC_743/Y 0.02fF
C63001 INVX1_LOC_256/Y NOR2X1_LOC_536/A 0.03fF
C63002 NOR2X1_LOC_172/Y NOR2X1_LOC_592/B 0.00fF
C63003 NAND2X1_LOC_388/a_36_24# INVX1_LOC_20/A 0.01fF
C63004 NOR2X1_LOC_576/B INVX1_LOC_11/Y 0.76fF
C63005 INVX1_LOC_12/Y INVX1_LOC_56/Y 0.03fF
C63006 INVX1_LOC_141/Y NOR2X1_LOC_89/A 0.03fF
C63007 INVX1_LOC_210/Y NOR2X1_LOC_340/A 0.01fF
C63008 NAND2X1_LOC_162/A INVX1_LOC_117/A 0.03fF
C63009 NAND2X1_LOC_675/a_36_24# INVX1_LOC_9/A 0.00fF
C63010 NOR2X1_LOC_142/Y NOR2X1_LOC_155/A 0.04fF
C63011 INVX1_LOC_141/Y NAND2X1_LOC_668/a_36_24# 0.00fF
C63012 NOR2X1_LOC_863/B NOR2X1_LOC_852/Y 0.09fF
C63013 NAND2X1_LOC_361/a_36_24# INVX1_LOC_92/A 0.01fF
C63014 NOR2X1_LOC_389/A NAND2X1_LOC_213/a_36_24# 0.06fF
C63015 NOR2X1_LOC_249/Y NOR2X1_LOC_35/a_36_216# 0.00fF
C63016 NAND2X1_LOC_326/A NAND2X1_LOC_175/Y 0.42fF
C63017 INVX1_LOC_7/A D_INPUT_3 0.10fF
C63018 NOR2X1_LOC_348/B INVX1_LOC_92/A 0.10fF
C63019 INVX1_LOC_313/Y NOR2X1_LOC_486/Y 0.00fF
C63020 INVX1_LOC_175/A NOR2X1_LOC_475/A 0.04fF
C63021 INVX1_LOC_57/Y INVX1_LOC_102/A 0.49fF
C63022 INVX1_LOC_83/A NAND2X1_LOC_453/A 0.10fF
C63023 NOR2X1_LOC_703/B INVX1_LOC_99/A 0.02fF
C63024 INVX1_LOC_18/A INVX1_LOC_12/A 3.07fF
C63025 NAND2X1_LOC_798/A NOR2X1_LOC_506/Y 0.14fF
C63026 INVX1_LOC_170/A INVX1_LOC_170/Y 0.10fF
C63027 NOR2X1_LOC_726/a_36_216# INVX1_LOC_85/Y 0.00fF
C63028 NAND2X1_LOC_728/Y INVX1_LOC_12/A 0.07fF
C63029 INVX1_LOC_58/A NOR2X1_LOC_510/Y 0.03fF
C63030 NOR2X1_LOC_103/Y NAND2X1_LOC_223/A 0.94fF
C63031 NOR2X1_LOC_160/B NOR2X1_LOC_227/A 0.01fF
C63032 NOR2X1_LOC_785/Y INVX1_LOC_117/A 0.00fF
C63033 NAND2X1_LOC_577/A INVX1_LOC_15/A 0.03fF
C63034 NOR2X1_LOC_773/a_36_216# INVX1_LOC_285/A 0.00fF
C63035 NOR2X1_LOC_75/Y NOR2X1_LOC_158/Y 0.13fF
C63036 NAND2X1_LOC_711/B INVX1_LOC_12/A 0.07fF
C63037 NOR2X1_LOC_534/a_36_216# NOR2X1_LOC_405/A 0.00fF
C63038 INVX1_LOC_28/A INVX1_LOC_20/A 0.21fF
C63039 NOR2X1_LOC_637/Y INVX1_LOC_12/A 0.05fF
C63040 INVX1_LOC_5/A INVX1_LOC_68/A 0.01fF
C63041 INVX1_LOC_17/A NOR2X1_LOC_318/A 0.14fF
C63042 INVX1_LOC_119/A INVX1_LOC_119/Y 0.04fF
C63043 INVX1_LOC_7/A INVX1_LOC_230/A 0.00fF
C63044 NOR2X1_LOC_191/a_36_216# INVX1_LOC_6/A 0.00fF
C63045 NOR2X1_LOC_184/a_36_216# NOR2X1_LOC_124/A 0.03fF
C63046 INVX1_LOC_232/A NOR2X1_LOC_78/Y 0.00fF
C63047 NOR2X1_LOC_605/a_36_216# INVX1_LOC_185/A 0.00fF
C63048 NAND2X1_LOC_555/Y NOR2X1_LOC_34/Y 0.04fF
C63049 INVX1_LOC_22/A INVX1_LOC_92/A 0.17fF
C63050 INVX1_LOC_58/A NOR2X1_LOC_361/B 0.09fF
C63051 NOR2X1_LOC_32/B NOR2X1_LOC_92/Y 0.13fF
C63052 NOR2X1_LOC_570/B INVX1_LOC_29/A 0.03fF
C63053 NAND2X1_LOC_803/B INVX1_LOC_50/A 0.02fF
C63054 NOR2X1_LOC_82/A INVX1_LOC_57/A 0.08fF
C63055 INVX1_LOC_75/A INVX1_LOC_46/A 0.06fF
C63056 NOR2X1_LOC_146/Y NAND2X1_LOC_425/Y 0.03fF
C63057 NOR2X1_LOC_790/B INVX1_LOC_269/A 0.02fF
C63058 NOR2X1_LOC_795/Y INVX1_LOC_19/A 0.03fF
C63059 INVX1_LOC_45/A INVX1_LOC_18/Y 0.05fF
C63060 INVX1_LOC_222/A NOR2X1_LOC_35/Y 0.11fF
C63061 INVX1_LOC_90/A NOR2X1_LOC_331/B 0.17fF
C63062 NAND2X1_LOC_30/Y INVX1_LOC_23/A 0.03fF
C63063 NOR2X1_LOC_186/Y INVX1_LOC_27/A 0.19fF
C63064 NAND2X1_LOC_807/Y NAND2X1_LOC_848/A 0.10fF
C63065 NOR2X1_LOC_557/A NAND2X1_LOC_642/Y 0.03fF
C63066 INVX1_LOC_88/Y NOR2X1_LOC_89/A 0.03fF
C63067 NAND2X1_LOC_325/Y INVX1_LOC_42/A 0.03fF
C63068 INVX1_LOC_60/Y NAND2X1_LOC_74/B 0.32fF
C63069 NAND2X1_LOC_35/Y NAND2X1_LOC_579/A 0.17fF
C63070 NAND2X1_LOC_741/B NOR2X1_LOC_829/A 0.02fF
C63071 NAND2X1_LOC_832/a_36_24# INVX1_LOC_186/Y 0.00fF
C63072 INVX1_LOC_50/A NOR2X1_LOC_590/A 0.10fF
C63073 NAND2X1_LOC_214/Y INVX1_LOC_5/A 0.01fF
C63074 NOR2X1_LOC_45/Y INVX1_LOC_271/A 0.06fF
C63075 NOR2X1_LOC_772/B NOR2X1_LOC_468/Y 0.02fF
C63076 NOR2X1_LOC_365/a_36_216# INVX1_LOC_109/Y 0.00fF
C63077 INVX1_LOC_155/A NOR2X1_LOC_116/a_36_216# 0.00fF
C63078 INVX1_LOC_256/A NOR2X1_LOC_717/A 0.19fF
C63079 INVX1_LOC_6/A NOR2X1_LOC_266/B 0.03fF
C63080 NOR2X1_LOC_846/A NAND2X1_LOC_473/A 0.03fF
C63081 INVX1_LOC_18/A NOR2X1_LOC_686/A 0.01fF
C63082 NOR2X1_LOC_13/Y NAND2X1_LOC_470/B 0.10fF
C63083 NAND2X1_LOC_787/A NOR2X1_LOC_369/Y 0.44fF
C63084 INVX1_LOC_41/A NOR2X1_LOC_620/A 0.05fF
C63085 NOR2X1_LOC_7/Y INVX1_LOC_76/A 0.03fF
C63086 NOR2X1_LOC_71/Y NAND2X1_LOC_244/a_36_24# 0.00fF
C63087 INVX1_LOC_34/Y INVX1_LOC_12/A 0.51fF
C63088 NOR2X1_LOC_250/Y NOR2X1_LOC_109/Y 0.03fF
C63089 NOR2X1_LOC_471/Y NOR2X1_LOC_678/A 0.02fF
C63090 INVX1_LOC_223/A NOR2X1_LOC_383/B 0.03fF
C63091 NAND2X1_LOC_655/A NAND2X1_LOC_655/B 0.01fF
C63092 NOR2X1_LOC_139/Y NAND2X1_LOC_469/B 0.05fF
C63093 NAND2X1_LOC_181/Y NAND2X1_LOC_81/B 0.03fF
C63094 NOR2X1_LOC_614/Y INVX1_LOC_19/A 0.01fF
C63095 INVX1_LOC_89/A NAND2X1_LOC_243/B 0.08fF
C63096 NAND2X1_LOC_359/Y NOR2X1_LOC_240/B 0.00fF
C63097 INVX1_LOC_21/A INVX1_LOC_1/A 0.11fF
C63098 NOR2X1_LOC_78/B NAND2X1_LOC_291/B 0.05fF
C63099 INVX1_LOC_276/A INVX1_LOC_42/A 0.03fF
C63100 INVX1_LOC_90/A NOR2X1_LOC_592/B 0.03fF
C63101 INVX1_LOC_136/A INVX1_LOC_29/Y 0.07fF
C63102 NOR2X1_LOC_67/A INVX1_LOC_42/A 0.36fF
C63103 NAND2X1_LOC_468/B NAND2X1_LOC_469/B 0.06fF
C63104 NAND2X1_LOC_848/A INVX1_LOC_6/A 0.01fF
C63105 INVX1_LOC_295/A NAND2X1_LOC_426/a_36_24# -0.02fF
C63106 INVX1_LOC_198/Y INVX1_LOC_275/Y 0.00fF
C63107 INVX1_LOC_35/A NOR2X1_LOC_726/Y 0.01fF
C63108 NOR2X1_LOC_78/B INVX1_LOC_283/A 0.00fF
C63109 INVX1_LOC_30/Y INVX1_LOC_125/A 0.02fF
C63110 INVX1_LOC_198/Y NOR2X1_LOC_748/A 0.10fF
C63111 NOR2X1_LOC_488/a_36_216# INVX1_LOC_42/A 0.00fF
C63112 NAND2X1_LOC_212/Y INVX1_LOC_76/A 0.04fF
C63113 INVX1_LOC_196/Y NOR2X1_LOC_800/a_36_216# 0.00fF
C63114 INVX1_LOC_215/A INVX1_LOC_29/A 0.07fF
C63115 NOR2X1_LOC_590/A NOR2X1_LOC_590/Y 0.02fF
C63116 NAND2X1_LOC_715/B NOR2X1_LOC_441/Y 0.29fF
C63117 INVX1_LOC_11/Y NOR2X1_LOC_27/a_36_216# 0.02fF
C63118 INVX1_LOC_21/A NOR2X1_LOC_794/B 0.05fF
C63119 NAND2X1_LOC_170/A INVX1_LOC_102/A 0.07fF
C63120 INVX1_LOC_279/A INVX1_LOC_272/A -0.02fF
C63121 NOR2X1_LOC_591/Y INVX1_LOC_94/Y 0.06fF
C63122 INVX1_LOC_11/A NAND2X1_LOC_780/Y 0.03fF
C63123 INVX1_LOC_65/A INVX1_LOC_117/A 0.19fF
C63124 INVX1_LOC_266/Y NOR2X1_LOC_465/Y 0.16fF
C63125 NAND2X1_LOC_464/Y NAND2X1_LOC_99/A 0.01fF
C63126 INVX1_LOC_14/Y INVX1_LOC_76/A 0.10fF
C63127 NOR2X1_LOC_356/A INVX1_LOC_63/A 0.07fF
C63128 NOR2X1_LOC_137/Y NAND2X1_LOC_211/Y 0.02fF
C63129 INVX1_LOC_133/Y INVX1_LOC_78/A 0.01fF
C63130 NOR2X1_LOC_32/B NAND2X1_LOC_837/Y 0.02fF
C63131 INVX1_LOC_8/A NOR2X1_LOC_39/Y 0.02fF
C63132 NAND2X1_LOC_656/Y NOR2X1_LOC_89/A 0.07fF
C63133 INVX1_LOC_103/A NOR2X1_LOC_217/a_36_216# 0.00fF
C63134 INVX1_LOC_49/A INVX1_LOC_23/A 0.38fF
C63135 INVX1_LOC_224/Y INVX1_LOC_33/A 1.76fF
C63136 NOR2X1_LOC_719/a_36_216# INVX1_LOC_284/A 0.02fF
C63137 INVX1_LOC_276/A INVX1_LOC_78/A 0.00fF
C63138 INVX1_LOC_6/A INVX1_LOC_46/Y 0.02fF
C63139 NOR2X1_LOC_313/a_36_216# NOR2X1_LOC_697/Y 0.00fF
C63140 NOR2X1_LOC_548/A NOR2X1_LOC_445/B 0.01fF
C63141 INVX1_LOC_58/A NOR2X1_LOC_132/Y 0.01fF
C63142 NOR2X1_LOC_577/Y INVX1_LOC_53/A 2.41fF
C63143 INVX1_LOC_16/A INVX1_LOC_4/A 0.25fF
C63144 INVX1_LOC_58/A INVX1_LOC_153/Y 0.10fF
C63145 INVX1_LOC_21/A NOR2X1_LOC_384/Y 0.07fF
C63146 INVX1_LOC_224/A NAND2X1_LOC_114/B 0.00fF
C63147 INVX1_LOC_8/A NAND2X1_LOC_205/A 0.10fF
C63148 NOR2X1_LOC_389/A INVX1_LOC_88/A 0.01fF
C63149 INVX1_LOC_89/A INVX1_LOC_284/A 0.24fF
C63150 NAND2X1_LOC_733/Y NOR2X1_LOC_536/Y 0.13fF
C63151 NOR2X1_LOC_489/B INVX1_LOC_77/A 0.01fF
C63152 INVX1_LOC_11/A NAND2X1_LOC_114/B 0.07fF
C63153 NOR2X1_LOC_510/Y NOR2X1_LOC_338/Y -0.03fF
C63154 NOR2X1_LOC_91/A INVX1_LOC_2/A 10.27fF
C63155 NOR2X1_LOC_388/Y NOR2X1_LOC_493/a_36_216# 0.00fF
C63156 NOR2X1_LOC_316/Y NOR2X1_LOC_383/B 0.01fF
C63157 NOR2X1_LOC_74/A INVX1_LOC_63/A 0.18fF
C63158 NOR2X1_LOC_91/A NOR2X1_LOC_226/A 0.10fF
C63159 NOR2X1_LOC_78/A NOR2X1_LOC_216/B 0.03fF
C63160 D_INPUT_1 NOR2X1_LOC_315/Y 0.07fF
C63161 NOR2X1_LOC_15/Y NOR2X1_LOC_372/Y 0.06fF
C63162 NOR2X1_LOC_67/A NOR2X1_LOC_65/B -0.02fF
C63163 INVX1_LOC_55/A NOR2X1_LOC_471/Y 0.03fF
C63164 NOR2X1_LOC_272/Y NOR2X1_LOC_759/Y 0.00fF
C63165 INVX1_LOC_11/A INVX1_LOC_141/Y 0.07fF
C63166 NAND2X1_LOC_866/B NOR2X1_LOC_754/A -0.03fF
C63167 INVX1_LOC_58/A INVX1_LOC_177/A 0.01fF
C63168 NOR2X1_LOC_272/Y INVX1_LOC_202/A 0.25fF
C63169 NOR2X1_LOC_537/Y NOR2X1_LOC_748/A 0.04fF
C63170 NOR2X1_LOC_9/Y INVX1_LOC_63/A 0.10fF
C63171 INVX1_LOC_2/A INVX1_LOC_23/A 0.14fF
C63172 INVX1_LOC_11/A INVX1_LOC_312/Y 0.07fF
C63173 INVX1_LOC_256/A NOR2X1_LOC_658/Y 0.02fF
C63174 NAND2X1_LOC_841/a_36_24# INVX1_LOC_186/Y 0.01fF
C63175 INVX1_LOC_104/A INVX1_LOC_292/Y 0.15fF
C63176 NAND2X1_LOC_51/B INVX1_LOC_261/Y 0.10fF
C63177 NOR2X1_LOC_226/A INVX1_LOC_23/A 0.14fF
C63178 INVX1_LOC_58/A INVX1_LOC_280/Y 0.02fF
C63179 INVX1_LOC_132/A INVX1_LOC_27/A 0.15fF
C63180 INVX1_LOC_224/Y INVX1_LOC_40/A 0.33fF
C63181 NAND2X1_LOC_53/Y NAND2X1_LOC_16/Y 0.11fF
C63182 NOR2X1_LOC_619/A NOR2X1_LOC_720/A 0.00fF
C63183 INVX1_LOC_200/A INVX1_LOC_18/A 0.08fF
C63184 INVX1_LOC_45/A NOR2X1_LOC_483/B 0.07fF
C63185 NOR2X1_LOC_454/Y NOR2X1_LOC_638/a_36_216# -0.01fF
C63186 INVX1_LOC_37/A INVX1_LOC_185/A 0.03fF
C63187 INVX1_LOC_162/A NOR2X1_LOC_652/Y 0.01fF
C63188 NOR2X1_LOC_489/A INVX1_LOC_129/Y 0.00fF
C63189 NOR2X1_LOC_431/a_36_216# INVX1_LOC_103/A 0.01fF
C63190 NOR2X1_LOC_329/B INVX1_LOC_15/A 0.07fF
C63191 NOR2X1_LOC_284/B NOR2X1_LOC_634/Y 0.02fF
C63192 INVX1_LOC_64/A NAND2X1_LOC_717/Y 0.06fF
C63193 NAND2X1_LOC_550/a_36_24# NAND2X1_LOC_464/B 0.00fF
C63194 NOR2X1_LOC_331/B INVX1_LOC_38/A 0.13fF
C63195 INVX1_LOC_286/A INVX1_LOC_29/A 0.12fF
C63196 NOR2X1_LOC_218/Y INVX1_LOC_23/A 0.01fF
C63197 INVX1_LOC_11/A NOR2X1_LOC_546/B 0.02fF
C63198 INVX1_LOC_14/A INVX1_LOC_77/A 0.02fF
C63199 INVX1_LOC_286/Y INVX1_LOC_30/A -0.01fF
C63200 INVX1_LOC_225/A INVX1_LOC_27/A 0.07fF
C63201 NOR2X1_LOC_817/Y INVX1_LOC_228/A 0.10fF
C63202 D_INPUT_4 INVX1_LOC_15/A 0.01fF
C63203 NAND2X1_LOC_685/a_36_24# INVX1_LOC_291/A 0.01fF
C63204 NOR2X1_LOC_45/B INVX1_LOC_19/A 0.18fF
C63205 INVX1_LOC_235/Y NOR2X1_LOC_459/B 0.05fF
C63206 INVX1_LOC_36/A INVX1_LOC_124/Y 0.17fF
C63207 INVX1_LOC_157/A NAND2X1_LOC_424/a_36_24# 0.01fF
C63208 INVX1_LOC_91/A INVX1_LOC_49/Y 0.06fF
C63209 NAND2X1_LOC_9/Y INVX1_LOC_25/Y 0.04fF
C63210 NAND2X1_LOC_563/Y INVX1_LOC_178/A 0.01fF
C63211 INVX1_LOC_22/A INVX1_LOC_53/A 0.13fF
C63212 NOR2X1_LOC_637/B INVX1_LOC_103/A 0.01fF
C63213 INVX1_LOC_50/A INVX1_LOC_227/A 0.14fF
C63214 NOR2X1_LOC_231/B NOR2X1_LOC_68/A 0.02fF
C63215 INVX1_LOC_90/A NOR2X1_LOC_621/B 0.01fF
C63216 NOR2X1_LOC_15/Y NAND2X1_LOC_276/Y 0.04fF
C63217 INVX1_LOC_233/A INVX1_LOC_25/Y 0.10fF
C63218 NAND2X1_LOC_51/B NOR2X1_LOC_467/A 0.07fF
C63219 NAND2X1_LOC_728/Y NAND2X1_LOC_733/Y 0.10fF
C63220 NOR2X1_LOC_223/B NOR2X1_LOC_222/Y 0.01fF
C63221 INVX1_LOC_17/A NOR2X1_LOC_335/A 0.04fF
C63222 INVX1_LOC_124/Y NOR2X1_LOC_267/A 0.17fF
C63223 INVX1_LOC_12/Y NOR2X1_LOC_831/B 0.05fF
C63224 NOR2X1_LOC_6/B NOR2X1_LOC_611/a_36_216# 0.01fF
C63225 NAND2X1_LOC_116/A NAND2X1_LOC_473/A 0.10fF
C63226 INVX1_LOC_6/A NOR2X1_LOC_754/A 0.02fF
C63227 NOR2X1_LOC_6/B NAND2X1_LOC_218/A 0.23fF
C63228 INVX1_LOC_91/A INVX1_LOC_99/A 0.06fF
C63229 NAND2X1_LOC_860/A NOR2X1_LOC_383/Y 0.21fF
C63230 NAND2X1_LOC_477/Y NAND2X1_LOC_464/A 0.01fF
C63231 NOR2X1_LOC_91/A NAND2X1_LOC_648/A 0.03fF
C63232 INVX1_LOC_64/A INVX1_LOC_16/A 14.30fF
C63233 NOR2X1_LOC_140/A NOR2X1_LOC_6/B 0.02fF
C63234 INVX1_LOC_11/A INVX1_LOC_275/A 0.09fF
C63235 INVX1_LOC_27/A NOR2X1_LOC_209/Y 0.26fF
C63236 NAND2X1_LOC_778/Y NAND2X1_LOC_374/Y 0.16fF
C63237 NOR2X1_LOC_52/B NAND2X1_LOC_780/Y 0.01fF
C63238 NOR2X1_LOC_91/A INPUT_1 0.39fF
C63239 INVX1_LOC_33/A NOR2X1_LOC_103/Y 0.08fF
C63240 NAND2X1_LOC_711/B NAND2X1_LOC_733/Y 0.10fF
C63241 INVX1_LOC_13/Y NOR2X1_LOC_220/A 0.05fF
C63242 NOR2X1_LOC_598/B NAND2X1_LOC_358/Y 0.02fF
C63243 NOR2X1_LOC_440/Y NOR2X1_LOC_717/A 0.09fF
C63244 INVX1_LOC_269/A NOR2X1_LOC_514/Y 0.03fF
C63245 INVX1_LOC_159/A INVX1_LOC_30/A 0.08fF
C63246 VDD NAND2X1_LOC_475/Y 0.76fF
C63247 INVX1_LOC_95/A INVX1_LOC_29/A 0.09fF
C63248 INVX1_LOC_33/A NOR2X1_LOC_541/Y 0.02fF
C63249 NAND2X1_LOC_553/A INVX1_LOC_25/Y 0.02fF
C63250 D_INPUT_0 NOR2X1_LOC_416/A 0.12fF
C63251 D_INPUT_7 NAND2X1_LOC_588/B 0.04fF
C63252 INVX1_LOC_217/A INVX1_LOC_18/A 0.10fF
C63253 INVX1_LOC_14/A NAND2X1_LOC_650/a_36_24# 0.00fF
C63254 NOR2X1_LOC_45/B NAND2X1_LOC_227/a_36_24# 0.00fF
C63255 INVX1_LOC_124/A INVX1_LOC_14/A 0.23fF
C63256 INVX1_LOC_313/Y NOR2X1_LOC_748/A 0.10fF
C63257 INVX1_LOC_49/A INVX1_LOC_31/A 0.03fF
C63258 NOR2X1_LOC_865/A NOR2X1_LOC_865/Y 0.01fF
C63259 INVX1_LOC_147/Y INVX1_LOC_109/A 0.49fF
C63260 INVX1_LOC_292/A INVX1_LOC_155/A 0.01fF
C63261 INVX1_LOC_1/Y INVX1_LOC_306/Y 0.00fF
C63262 NOR2X1_LOC_598/B NOR2X1_LOC_99/B 0.46fF
C63263 INVX1_LOC_126/A NAND2X1_LOC_74/B 0.03fF
C63264 INVX1_LOC_227/A NAND2X1_LOC_72/Y 0.01fF
C63265 NOR2X1_LOC_791/B NOR2X1_LOC_791/a_36_216# 0.00fF
C63266 NOR2X1_LOC_865/A NOR2X1_LOC_243/B 0.03fF
C63267 INPUT_1 INVX1_LOC_23/A 0.36fF
C63268 NOR2X1_LOC_15/Y NAND2X1_LOC_374/Y 0.33fF
C63269 INVX1_LOC_30/Y NOR2X1_LOC_81/Y 0.02fF
C63270 NOR2X1_LOC_598/B NOR2X1_LOC_846/B 0.03fF
C63271 NAND2X1_LOC_396/a_36_24# INVX1_LOC_168/A 0.00fF
C63272 NOR2X1_LOC_332/A INVX1_LOC_68/A 0.03fF
C63273 D_INPUT_0 NOR2X1_LOC_109/Y 0.14fF
C63274 INVX1_LOC_45/A INVX1_LOC_33/A 0.57fF
C63275 NOR2X1_LOC_384/a_36_216# NAND2X1_LOC_787/B 0.01fF
C63276 NOR2X1_LOC_866/B D_GATE_865 0.18fF
C63277 INVX1_LOC_172/A INVX1_LOC_217/A 0.07fF
C63278 NOR2X1_LOC_111/A NAND2X1_LOC_74/B 0.07fF
C63279 INPUT_3 NOR2X1_LOC_87/B 0.08fF
C63280 NOR2X1_LOC_276/Y NOR2X1_LOC_361/Y 0.00fF
C63281 NOR2X1_LOC_68/A NOR2X1_LOC_228/a_36_216# 0.02fF
C63282 INVX1_LOC_89/A NOR2X1_LOC_663/A 0.18fF
C63283 NOR2X1_LOC_598/B INVX1_LOC_182/A 0.02fF
C63284 INVX1_LOC_256/A INVX1_LOC_256/Y 0.11fF
C63285 NOR2X1_LOC_134/Y NOR2X1_LOC_290/Y 0.04fF
C63286 INVX1_LOC_141/Y NOR2X1_LOC_52/B 0.00fF
C63287 NOR2X1_LOC_830/Y INVX1_LOC_117/A 0.00fF
C63288 INVX1_LOC_185/Y INVX1_LOC_30/A 0.01fF
C63289 NOR2X1_LOC_103/Y INVX1_LOC_40/A 0.15fF
C63290 INVX1_LOC_64/A INVX1_LOC_28/A 0.38fF
C63291 INVX1_LOC_2/A INVX1_LOC_31/A 0.08fF
C63292 NOR2X1_LOC_52/B INVX1_LOC_312/Y 0.07fF
C63293 INVX1_LOC_31/A NOR2X1_LOC_818/Y 0.04fF
C63294 NAND2X1_LOC_9/Y INVX1_LOC_75/A 0.03fF
C63295 NOR2X1_LOC_226/A NAND2X1_LOC_509/a_36_24# 0.00fF
C63296 INVX1_LOC_97/Y INVX1_LOC_182/A -0.01fF
C63297 NAND2X1_LOC_303/Y NOR2X1_LOC_561/Y 0.10fF
C63298 NOR2X1_LOC_678/a_36_216# NAND2X1_LOC_656/Y 0.01fF
C63299 INVX1_LOC_225/Y NOR2X1_LOC_388/a_36_216# 0.00fF
C63300 NOR2X1_LOC_226/A INVX1_LOC_31/A 0.07fF
C63301 INVX1_LOC_136/A INVX1_LOC_60/Y 0.01fF
C63302 INVX1_LOC_233/A INVX1_LOC_75/A 0.07fF
C63303 NOR2X1_LOC_758/Y NAND2X1_LOC_198/B 0.18fF
C63304 NAND2X1_LOC_214/Y NOR2X1_LOC_332/A 0.04fF
C63305 INVX1_LOC_58/A INVX1_LOC_285/Y 0.01fF
C63306 INVX1_LOC_33/A INVX1_LOC_71/A 0.23fF
C63307 NOR2X1_LOC_160/B NOR2X1_LOC_121/a_36_216# 0.02fF
C63308 NOR2X1_LOC_186/Y NOR2X1_LOC_772/A 0.02fF
C63309 INVX1_LOC_304/Y INVX1_LOC_18/A 0.25fF
C63310 NOR2X1_LOC_160/B INVX1_LOC_56/Y 0.03fF
C63311 NAND2X1_LOC_363/B NOR2X1_LOC_721/Y 0.03fF
C63312 INVX1_LOC_269/A NOR2X1_LOC_128/B 0.01fF
C63313 NAND2X1_LOC_506/a_36_24# NOR2X1_LOC_849/A 0.00fF
C63314 INVX1_LOC_127/A NAND2X1_LOC_74/B 0.01fF
C63315 INVX1_LOC_43/Y INVX1_LOC_16/A 0.03fF
C63316 INVX1_LOC_54/A INVX1_LOC_29/A 0.17fF
C63317 INVX1_LOC_186/Y INVX1_LOC_92/A 0.08fF
C63318 NOR2X1_LOC_219/B NOR2X1_LOC_433/A 0.01fF
C63319 NAND2X1_LOC_736/Y NAND2X1_LOC_866/A 0.26fF
C63320 INVX1_LOC_69/Y NOR2X1_LOC_717/A 0.10fF
C63321 NOR2X1_LOC_265/a_36_216# INVX1_LOC_30/A 0.00fF
C63322 INVX1_LOC_19/A NOR2X1_LOC_862/B 0.02fF
C63323 NOR2X1_LOC_334/Y NOR2X1_LOC_858/B 0.03fF
C63324 NAND2X1_LOC_656/A NOR2X1_LOC_63/a_36_216# 0.08fF
C63325 INVX1_LOC_229/A NAND2X1_LOC_866/B 0.04fF
C63326 INVX1_LOC_214/Y INVX1_LOC_18/A 0.14fF
C63327 INVX1_LOC_238/A NAND2X1_LOC_866/a_36_24# 0.01fF
C63328 NAND2X1_LOC_733/Y NOR2X1_LOC_690/Y 0.03fF
C63329 INVX1_LOC_304/Y INVX1_LOC_172/A 0.07fF
C63330 INVX1_LOC_117/A INVX1_LOC_4/Y 2.00fF
C63331 NOR2X1_LOC_92/Y NAND2X1_LOC_842/a_36_24# 0.01fF
C63332 NAND2X1_LOC_717/Y NAND2X1_LOC_863/Y 0.40fF
C63333 NOR2X1_LOC_226/A INVX1_LOC_111/A 0.26fF
C63334 INVX1_LOC_41/A NOR2X1_LOC_720/B 0.00fF
C63335 NOR2X1_LOC_388/Y NOR2X1_LOC_392/B 0.01fF
C63336 NOR2X1_LOC_773/Y INVX1_LOC_181/Y 1.01fF
C63337 INVX1_LOC_59/Y INVX1_LOC_57/A 0.03fF
C63338 NAND2X1_LOC_67/Y NOR2X1_LOC_736/a_36_216# 0.01fF
C63339 NOR2X1_LOC_219/B NOR2X1_LOC_52/B 0.05fF
C63340 INVX1_LOC_276/A NOR2X1_LOC_152/Y 0.10fF
C63341 INVX1_LOC_111/Y INVX1_LOC_77/A 0.01fF
C63342 NOR2X1_LOC_751/Y NOR2X1_LOC_748/Y 0.01fF
C63343 INVX1_LOC_21/A NOR2X1_LOC_188/A 0.63fF
C63344 INVX1_LOC_21/A NOR2X1_LOC_548/B 0.12fF
C63345 NOR2X1_LOC_521/Y NOR2X1_LOC_384/Y 0.00fF
C63346 INVX1_LOC_176/A INVX1_LOC_57/A 0.02fF
C63347 INVX1_LOC_40/A INVX1_LOC_71/A 0.06fF
C63348 NOR2X1_LOC_78/B NOR2X1_LOC_577/Y 0.17fF
C63349 NOR2X1_LOC_124/B NAND2X1_LOC_122/a_36_24# 0.02fF
C63350 INVX1_LOC_1/A NAND2X1_LOC_51/B 0.03fF
C63351 NAND2X1_LOC_563/Y NAND2X1_LOC_562/B 0.09fF
C63352 NOR2X1_LOC_467/a_36_216# NOR2X1_LOC_68/A 0.00fF
C63353 NOR2X1_LOC_382/Y NOR2X1_LOC_130/A 0.07fF
C63354 INVX1_LOC_2/Y NOR2X1_LOC_414/Y 0.11fF
C63355 NOR2X1_LOC_498/Y NOR2X1_LOC_822/Y 0.04fF
C63356 NOR2X1_LOC_468/Y NOR2X1_LOC_83/a_36_216# 0.01fF
C63357 NAND2X1_LOC_773/B NAND2X1_LOC_772/a_36_24# 0.02fF
C63358 NOR2X1_LOC_848/Y NAND2X1_LOC_348/A 0.01fF
C63359 NOR2X1_LOC_424/a_36_216# NOR2X1_LOC_68/A 0.00fF
C63360 INVX1_LOC_36/A D_INPUT_0 0.09fF
C63361 INVX1_LOC_31/A INPUT_1 0.28fF
C63362 NOR2X1_LOC_373/Y NAND2X1_LOC_634/Y 0.03fF
C63363 NOR2X1_LOC_99/Y NOR2X1_LOC_38/B 0.06fF
C63364 INVX1_LOC_1/A INVX1_LOC_311/A 1.64fF
C63365 INVX1_LOC_18/A NAND2X1_LOC_808/A 0.07fF
C63366 NOR2X1_LOC_637/A INVX1_LOC_10/A 0.01fF
C63367 INVX1_LOC_89/A INVX1_LOC_72/A 0.07fF
C63368 INVX1_LOC_64/A NOR2X1_LOC_35/Y 0.03fF
C63369 NOR2X1_LOC_861/a_36_216# NOR2X1_LOC_38/B 0.00fF
C63370 NOR2X1_LOC_607/A INVX1_LOC_10/A 0.01fF
C63371 NAND2X1_LOC_787/A VDD 0.82fF
C63372 INVX1_LOC_5/A NOR2X1_LOC_833/Y 0.01fF
C63373 NOR2X1_LOC_791/Y NOR2X1_LOC_123/a_36_216# 0.00fF
C63374 INVX1_LOC_13/A NOR2X1_LOC_419/Y 0.03fF
C63375 NOR2X1_LOC_78/B NOR2X1_LOC_348/B 1.45fF
C63376 NOR2X1_LOC_334/Y NOR2X1_LOC_809/B 0.03fF
C63377 NOR2X1_LOC_773/Y NOR2X1_LOC_192/a_36_216# 0.00fF
C63378 NAND2X1_LOC_363/B VDD 0.01fF
C63379 INVX1_LOC_27/A NAND2X1_LOC_642/Y 0.84fF
C63380 NOR2X1_LOC_1/Y NOR2X1_LOC_11/Y 0.01fF
C63381 NOR2X1_LOC_91/A INVX1_LOC_118/A 0.38fF
C63382 INVX1_LOC_237/Y NAND2X1_LOC_735/B 0.01fF
C63383 D_INPUT_0 INVX1_LOC_145/A 0.02fF
C63384 INVX1_LOC_89/A INVX1_LOC_198/Y 0.01fF
C63385 NOR2X1_LOC_210/A NOR2X1_LOC_162/Y 0.06fF
C63386 INVX1_LOC_34/A NAND2X1_LOC_712/A 0.01fF
C63387 NOR2X1_LOC_433/A NAND2X1_LOC_656/Y 0.69fF
C63388 NAND2X1_LOC_807/B INVX1_LOC_29/A 0.10fF
C63389 INVX1_LOC_172/A NAND2X1_LOC_808/A 0.03fF
C63390 D_INPUT_0 NOR2X1_LOC_237/Y 0.16fF
C63391 INVX1_LOC_83/A NOR2X1_LOC_577/Y 0.10fF
C63392 NAND2X1_LOC_349/a_36_24# NOR2X1_LOC_52/B 0.00fF
C63393 INVX1_LOC_77/A NOR2X1_LOC_137/A 1.18fF
C63394 INVX1_LOC_230/Y NOR2X1_LOC_391/a_36_216# 0.01fF
C63395 NOR2X1_LOC_691/B INVX1_LOC_15/A 0.07fF
C63396 VDD NOR2X1_LOC_840/A 0.12fF
C63397 NOR2X1_LOC_134/Y INVX1_LOC_6/A 0.01fF
C63398 INVX1_LOC_26/Y NOR2X1_LOC_862/B 0.05fF
C63399 INVX1_LOC_32/A NAND2X1_LOC_219/B 0.02fF
C63400 NOR2X1_LOC_561/Y NAND2X1_LOC_466/Y 0.04fF
C63401 NOR2X1_LOC_48/B INVX1_LOC_29/A 0.09fF
C63402 NOR2X1_LOC_791/Y VDD 0.32fF
C63403 INVX1_LOC_23/A INVX1_LOC_118/A 9.64fF
C63404 D_INPUT_0 NOR2X1_LOC_804/B 0.09fF
C63405 NAND2X1_LOC_402/B INVX1_LOC_241/Y 0.60fF
C63406 INVX1_LOC_49/A INVX1_LOC_313/A 1.21fF
C63407 NOR2X1_LOC_721/Y INVX1_LOC_30/A 0.00fF
C63408 INVX1_LOC_33/A NOR2X1_LOC_123/B 0.07fF
C63409 INVX1_LOC_161/Y NOR2X1_LOC_45/B 0.15fF
C63410 NAND2X1_LOC_736/Y NOR2X1_LOC_700/Y 0.19fF
C63411 INVX1_LOC_30/Y NOR2X1_LOC_709/A 0.12fF
C63412 INVX1_LOC_270/Y NOR2X1_LOC_743/Y 0.06fF
C63413 NOR2X1_LOC_49/a_36_216# INVX1_LOC_23/Y 0.01fF
C63414 NAND2X1_LOC_848/A NOR2X1_LOC_109/Y 0.10fF
C63415 INVX1_LOC_79/A INVX1_LOC_79/Y 0.09fF
C63416 NOR2X1_LOC_67/A NAND2X1_LOC_859/B 0.03fF
C63417 NOR2X1_LOC_78/B INVX1_LOC_22/A 9.68fF
C63418 NOR2X1_LOC_703/B INPUT_0 0.06fF
C63419 INVX1_LOC_163/A D_GATE_479 0.01fF
C63420 NAND2X1_LOC_303/Y INVX1_LOC_76/A 0.32fF
C63421 NOR2X1_LOC_52/B NAND2X1_LOC_656/Y 0.10fF
C63422 D_INPUT_0 NOR2X1_LOC_309/Y 0.07fF
C63423 NAND2X1_LOC_563/Y NOR2X1_LOC_332/A -0.02fF
C63424 INVX1_LOC_222/A NAND2X1_LOC_272/a_36_24# 0.00fF
C63425 INVX1_LOC_90/A NOR2X1_LOC_388/Y 0.04fF
C63426 NOR2X1_LOC_416/A INVX1_LOC_46/Y 0.04fF
C63427 NAND2X1_LOC_3/B INVX1_LOC_29/A 0.08fF
C63428 NOR2X1_LOC_226/A NAND2X1_LOC_859/Y 0.00fF
C63429 INVX1_LOC_124/A NOR2X1_LOC_137/A 0.13fF
C63430 NOR2X1_LOC_309/Y NOR2X1_LOC_389/a_36_216# 0.00fF
C63431 NOR2X1_LOC_298/Y NAND2X1_LOC_839/A 0.04fF
C63432 NOR2X1_LOC_418/Y INVX1_LOC_290/A 0.01fF
C63433 INVX1_LOC_308/Y NAND2X1_LOC_287/B 0.03fF
C63434 INVX1_LOC_41/A NAND2X1_LOC_842/a_36_24# 0.00fF
C63435 INVX1_LOC_36/A NOR2X1_LOC_191/a_36_216# 0.00fF
C63436 INVX1_LOC_27/A NOR2X1_LOC_271/Y 0.12fF
C63437 NOR2X1_LOC_646/A NOR2X1_LOC_646/a_36_216# 0.02fF
C63438 NAND2X1_LOC_21/Y D_INPUT_4 0.25fF
C63439 INVX1_LOC_225/A NOR2X1_LOC_772/A 0.01fF
C63440 INVX1_LOC_89/A INVX1_LOC_192/Y 0.00fF
C63441 INVX1_LOC_246/A INVX1_LOC_20/A 0.02fF
C63442 NOR2X1_LOC_457/A VDD 0.48fF
C63443 NAND2X1_LOC_563/A NOR2X1_LOC_128/B 0.01fF
C63444 INVX1_LOC_89/A NOR2X1_LOC_537/Y 0.20fF
C63445 NOR2X1_LOC_290/Y INPUT_1 0.41fF
C63446 NOR2X1_LOC_589/A INVX1_LOC_290/A 0.03fF
C63447 INVX1_LOC_89/A NAND2X1_LOC_338/B 0.15fF
C63448 NAND2X1_LOC_656/A INVX1_LOC_123/A 0.10fF
C63449 NOR2X1_LOC_493/B INVX1_LOC_313/Y 0.03fF
C63450 INVX1_LOC_94/A NOR2X1_LOC_501/B 0.02fF
C63451 NOR2X1_LOC_474/A NAND2X1_LOC_622/B 0.39fF
C63452 INVX1_LOC_30/A NOR2X1_LOC_56/Y 0.07fF
C63453 INVX1_LOC_89/A NAND2X1_LOC_323/B 0.03fF
C63454 NOR2X1_LOC_488/a_36_216# NAND2X1_LOC_861/Y 0.01fF
C63455 INVX1_LOC_77/A INVX1_LOC_48/A 0.02fF
C63456 INVX1_LOC_49/A INVX1_LOC_6/A 0.37fF
C63457 INVX1_LOC_83/A NOR2X1_LOC_325/A 1.21fF
C63458 INVX1_LOC_2/A NAND2X1_LOC_807/Y 0.04fF
C63459 INVX1_LOC_83/A INVX1_LOC_22/A 0.04fF
C63460 INVX1_LOC_212/A NOR2X1_LOC_78/A 0.03fF
C63461 NOR2X1_LOC_394/Y INVX1_LOC_32/A 0.02fF
C63462 INVX1_LOC_35/A INVX1_LOC_84/A 0.10fF
C63463 NOR2X1_LOC_186/Y NOR2X1_LOC_216/B 0.13fF
C63464 NOR2X1_LOC_500/A NOR2X1_LOC_78/A 0.07fF
C63465 INVX1_LOC_14/A INVX1_LOC_9/A 0.02fF
C63466 NOR2X1_LOC_226/A NAND2X1_LOC_807/Y 0.07fF
C63467 NOR2X1_LOC_297/A NAND2X1_LOC_296/a_36_24# 0.00fF
C63468 NOR2X1_LOC_384/Y NOR2X1_LOC_670/Y 0.01fF
C63469 NOR2X1_LOC_529/a_36_216# NOR2X1_LOC_671/Y 0.00fF
C63470 INVX1_LOC_34/A INVX1_LOC_309/A 0.03fF
C63471 NOR2X1_LOC_274/a_36_216# NOR2X1_LOC_405/A 0.00fF
C63472 NOR2X1_LOC_328/Y NOR2X1_LOC_224/a_36_216# 0.00fF
C63473 INVX1_LOC_30/A VDD 8.93fF
C63474 INVX1_LOC_36/A NOR2X1_LOC_266/B 0.06fF
C63475 NAND2X1_LOC_842/B INVX1_LOC_25/Y 0.15fF
C63476 INVX1_LOC_213/Y NOR2X1_LOC_730/B 0.02fF
C63477 NOR2X1_LOC_577/Y NOR2X1_LOC_311/Y 0.00fF
C63478 INVX1_LOC_53/A NOR2X1_LOC_777/B 0.03fF
C63479 NAND2X1_LOC_763/B VDD 0.01fF
C63480 INVX1_LOC_290/Y NOR2X1_LOC_383/B 0.09fF
C63481 NOR2X1_LOC_274/B INVX1_LOC_46/A 0.15fF
C63482 NOR2X1_LOC_486/Y INVX1_LOC_71/A 1.46fF
C63483 NOR2X1_LOC_267/A NOR2X1_LOC_266/B 0.15fF
C63484 INVX1_LOC_83/A NOR2X1_LOC_784/B 0.06fF
C63485 INVX1_LOC_1/Y NOR2X1_LOC_73/a_36_216# 0.00fF
C63486 INVX1_LOC_34/A INVX1_LOC_91/A 0.23fF
C63487 NOR2X1_LOC_381/Y NOR2X1_LOC_104/a_36_216# 0.00fF
C63488 INVX1_LOC_271/A NAND2X1_LOC_792/B 0.01fF
C63489 INVX1_LOC_136/A NOR2X1_LOC_111/A 0.10fF
C63490 INVX1_LOC_230/Y NOR2X1_LOC_96/a_36_216# 0.00fF
C63491 NAND2X1_LOC_9/Y NAND2X1_LOC_291/B 0.04fF
C63492 INVX1_LOC_225/A NOR2X1_LOC_528/Y 0.01fF
C63493 NOR2X1_LOC_89/A NOR2X1_LOC_717/A 0.08fF
C63494 INVX1_LOC_2/A INVX1_LOC_6/A 0.49fF
C63495 INVX1_LOC_103/A NOR2X1_LOC_510/B 0.03fF
C63496 NAND2X1_LOC_53/Y NOR2X1_LOC_433/Y 0.02fF
C63497 NAND2X1_LOC_21/Y INPUT_4 0.14fF
C63498 INVX1_LOC_256/A NOR2X1_LOC_640/Y 0.07fF
C63499 NOR2X1_LOC_392/Y INVX1_LOC_284/A 0.01fF
C63500 INVX1_LOC_36/A NAND2X1_LOC_848/A 0.01fF
C63501 NOR2X1_LOC_219/B INVX1_LOC_199/A 0.13fF
C63502 INVX1_LOC_31/A INVX1_LOC_118/A 0.24fF
C63503 INVX1_LOC_135/A INVX1_LOC_90/A 0.57fF
C63504 NOR2X1_LOC_257/a_36_216# INVX1_LOC_37/A 0.00fF
C63505 NOR2X1_LOC_598/B NOR2X1_LOC_850/B 0.03fF
C63506 INVX1_LOC_294/Y INVX1_LOC_93/Y 0.09fF
C63507 INVX1_LOC_34/A INVX1_LOC_11/Y 0.97fF
C63508 NOR2X1_LOC_226/A INVX1_LOC_6/A 0.24fF
C63509 NOR2X1_LOC_68/A INVX1_LOC_33/Y 0.06fF
C63510 INVX1_LOC_282/A INVX1_LOC_16/A 0.19fF
C63511 NOR2X1_LOC_318/A INVX1_LOC_94/Y 0.00fF
C63512 INVX1_LOC_231/Y INVX1_LOC_20/A 0.44fF
C63513 NOR2X1_LOC_274/Y INVX1_LOC_14/Y 0.01fF
C63514 NOR2X1_LOC_690/A NOR2X1_LOC_824/Y 0.04fF
C63515 INVX1_LOC_1/Y NOR2X1_LOC_74/A 0.10fF
C63516 INVX1_LOC_89/A INVX1_LOC_313/Y 0.07fF
C63517 INVX1_LOC_295/A NAND2X1_LOC_769/a_36_24# 0.06fF
C63518 INVX1_LOC_203/Y D_GATE_479 0.26fF
C63519 INVX1_LOC_45/A NOR2X1_LOC_833/a_36_216# 0.00fF
C63520 NOR2X1_LOC_412/a_36_216# INVX1_LOC_20/A 0.00fF
C63521 NOR2X1_LOC_577/Y INVX1_LOC_46/A 0.21fF
C63522 NAND2X1_LOC_231/Y INVX1_LOC_91/A 0.10fF
C63523 NOR2X1_LOC_242/A NOR2X1_LOC_777/B 0.00fF
C63524 NAND2X1_LOC_647/B INVX1_LOC_29/Y 0.05fF
C63525 INPUT_0 INVX1_LOC_137/Y 0.01fF
C63526 NOR2X1_LOC_272/Y NAND2X1_LOC_74/B 0.01fF
C63527 NOR2X1_LOC_690/A INVX1_LOC_76/A 0.10fF
C63528 NOR2X1_LOC_160/B NOR2X1_LOC_831/B 0.01fF
C63529 NOR2X1_LOC_218/Y INVX1_LOC_6/A 0.04fF
C63530 INVX1_LOC_32/A INVX1_LOC_58/Y 0.06fF
C63531 INVX1_LOC_155/A NOR2X1_LOC_137/Y 0.00fF
C63532 NOR2X1_LOC_335/B NOR2X1_LOC_188/Y 0.16fF
C63533 INVX1_LOC_1/Y NOR2X1_LOC_9/Y 0.75fF
C63534 INVX1_LOC_23/A NAND2X1_LOC_618/Y 0.54fF
C63535 INVX1_LOC_227/Y INVX1_LOC_9/A 0.03fF
C63536 INVX1_LOC_58/A INVX1_LOC_4/Y 0.22fF
C63537 INVX1_LOC_35/A INVX1_LOC_15/A 0.24fF
C63538 INVX1_LOC_25/A NOR2X1_LOC_248/A 0.03fF
C63539 NAND2X1_LOC_634/Y INVX1_LOC_54/A 0.01fF
C63540 NAND2X1_LOC_175/Y NOR2X1_LOC_654/A 0.10fF
C63541 D_INPUT_6 INVX1_LOC_12/A 0.01fF
C63542 INVX1_LOC_135/A NAND2X1_LOC_348/A 2.67fF
C63543 NOR2X1_LOC_173/Y INVX1_LOC_12/A 0.09fF
C63544 NOR2X1_LOC_389/B NOR2X1_LOC_248/a_36_216# 0.01fF
C63545 NAND2X1_LOC_200/B NAND2X1_LOC_642/Y 0.01fF
C63546 INVX1_LOC_13/A NOR2X1_LOC_392/a_36_216# 0.01fF
C63547 NOR2X1_LOC_237/Y NAND2X1_LOC_848/A 0.10fF
C63548 INVX1_LOC_266/Y NOR2X1_LOC_603/Y 0.01fF
C63549 NOR2X1_LOC_84/Y INVX1_LOC_20/A 0.17fF
C63550 NOR2X1_LOC_348/B INVX1_LOC_46/A 0.03fF
C63551 NAND2X1_LOC_90/a_36_24# NAND2X1_LOC_99/A 0.00fF
C63552 INVX1_LOC_18/A INVX1_LOC_92/A 1.47fF
C63553 NOR2X1_LOC_843/A INVX1_LOC_117/A 0.26fF
C63554 NAND2X1_LOC_348/A NOR2X1_LOC_560/A 0.07fF
C63555 INVX1_LOC_55/Y NOR2X1_LOC_151/Y 0.03fF
C63556 NAND2X1_LOC_842/B INVX1_LOC_75/A 1.18fF
C63557 INVX1_LOC_183/Y INPUT_0 0.06fF
C63558 D_INPUT_1 NAND2X1_LOC_99/A 0.22fF
C63559 NAND2X1_LOC_722/A VDD 0.04fF
C63560 NAND2X1_LOC_510/A NAND2X1_LOC_574/A 0.02fF
C63561 INVX1_LOC_33/A NOR2X1_LOC_331/B 0.15fF
C63562 NOR2X1_LOC_468/Y NOR2X1_LOC_76/B 0.01fF
C63563 INVX1_LOC_137/A NAND2X1_LOC_642/Y 0.01fF
C63564 INPUT_3 NAND2X1_LOC_219/B 0.23fF
C63565 INVX1_LOC_50/A NOR2X1_LOC_441/a_36_216# 0.00fF
C63566 NAND2X1_LOC_474/Y INVX1_LOC_47/Y 0.34fF
C63567 NAND2X1_LOC_348/A NOR2X1_LOC_346/a_36_216# 0.00fF
C63568 INVX1_LOC_124/Y INVX1_LOC_63/A 0.07fF
C63569 NOR2X1_LOC_637/Y INVX1_LOC_92/A 2.46fF
C63570 INVX1_LOC_159/A INVX1_LOC_113/A 0.05fF
C63571 INVX1_LOC_50/Y NOR2X1_LOC_334/Y 0.07fF
C63572 NOR2X1_LOC_309/Y NAND2X1_LOC_848/A 0.10fF
C63573 INVX1_LOC_6/A INPUT_1 0.10fF
C63574 NOR2X1_LOC_389/A INVX1_LOC_272/A 0.10fF
C63575 NOR2X1_LOC_742/A NOR2X1_LOC_74/A 1.01fF
C63576 INVX1_LOC_31/A NAND2X1_LOC_63/Y 0.02fF
C63577 NOR2X1_LOC_239/a_36_216# NOR2X1_LOC_721/B 0.00fF
C63578 NOR2X1_LOC_441/Y INVX1_LOC_29/A 0.23fF
C63579 INVX1_LOC_186/A INVX1_LOC_85/Y 0.00fF
C63580 NOR2X1_LOC_620/B NAND2X1_LOC_96/A 0.04fF
C63581 INVX1_LOC_22/A INVX1_LOC_46/A 0.36fF
C63582 NAND2X1_LOC_300/a_36_24# NOR2X1_LOC_743/Y 0.00fF
C63583 NOR2X1_LOC_646/a_36_216# INVX1_LOC_2/Y 0.00fF
C63584 NAND2X1_LOC_348/A NOR2X1_LOC_391/B 0.12fF
C63585 NOR2X1_LOC_318/B NOR2X1_LOC_356/A 0.02fF
C63586 INVX1_LOC_266/A NOR2X1_LOC_334/Y 0.00fF
C63587 INVX1_LOC_90/A NOR2X1_LOC_552/A 0.07fF
C63588 INVX1_LOC_111/Y INVX1_LOC_9/A 0.05fF
C63589 INVX1_LOC_1/A NOR2X1_LOC_248/A 0.01fF
C63590 NOR2X1_LOC_290/Y INVX1_LOC_118/A 0.09fF
C63591 NOR2X1_LOC_112/Y NOR2X1_LOC_78/A 0.03fF
C63592 NOR2X1_LOC_91/A INVX1_LOC_39/A 0.03fF
C63593 INVX1_LOC_191/Y INVX1_LOC_118/A 0.03fF
C63594 INVX1_LOC_35/A INVX1_LOC_108/Y 0.18fF
C63595 NOR2X1_LOC_826/a_36_216# INVX1_LOC_64/A 0.00fF
C63596 INVX1_LOC_225/A NOR2X1_LOC_216/B 0.29fF
C63597 INVX1_LOC_35/A INVX1_LOC_278/A 0.07fF
C63598 INVX1_LOC_213/Y NOR2X1_LOC_155/A 0.03fF
C63599 INVX1_LOC_174/A NOR2X1_LOC_467/A 0.42fF
C63600 INVX1_LOC_131/A INVX1_LOC_91/A 0.10fF
C63601 NAND2X1_LOC_364/A NAND2X1_LOC_74/B 0.10fF
C63602 NAND2X1_LOC_16/Y INVX1_LOC_12/A 0.12fF
C63603 INVX1_LOC_85/A INVX1_LOC_179/A 0.00fF
C63604 NAND2X1_LOC_466/A NOR2X1_LOC_592/B 0.01fF
C63605 INVX1_LOC_69/Y NOR2X1_LOC_337/A 0.03fF
C63606 NAND2X1_LOC_538/Y INVX1_LOC_273/A 0.03fF
C63607 NOR2X1_LOC_350/A NOR2X1_LOC_68/a_36_216# 0.00fF
C63608 NOR2X1_LOC_32/B NAND2X1_LOC_35/Y 0.07fF
C63609 NOR2X1_LOC_389/B NOR2X1_LOC_566/a_36_216# 0.00fF
C63610 INVX1_LOC_73/A NOR2X1_LOC_269/Y 0.03fF
C63611 NOR2X1_LOC_86/Y INVX1_LOC_284/A 0.01fF
C63612 NOR2X1_LOC_750/Y NAND2X1_LOC_214/B 0.00fF
C63613 INVX1_LOC_276/A INVX1_LOC_291/A 1.69fF
C63614 INVX1_LOC_161/A INVX1_LOC_231/A -0.00fF
C63615 NAND2X1_LOC_721/B NOR2X1_LOC_48/B 0.03fF
C63616 INVX1_LOC_200/A NAND2X1_LOC_443/a_36_24# 0.00fF
C63617 INVX1_LOC_39/A INVX1_LOC_23/A 0.03fF
C63618 INVX1_LOC_137/A NOR2X1_LOC_271/Y 0.02fF
C63619 INVX1_LOC_21/A NAND2X1_LOC_784/A 0.01fF
C63620 INPUT_0 INVX1_LOC_91/A 3.99fF
C63621 NOR2X1_LOC_251/a_36_216# INVX1_LOC_50/A -0.00fF
C63622 NOR2X1_LOC_273/Y INVX1_LOC_109/Y 0.02fF
C63623 INVX1_LOC_34/A INVX1_LOC_203/A 0.03fF
C63624 INVX1_LOC_215/A INVX1_LOC_118/Y 0.07fF
C63625 NOR2X1_LOC_326/Y NOR2X1_LOC_319/B 0.26fF
C63626 NAND2X1_LOC_734/B INVX1_LOC_119/Y 0.04fF
C63627 NOR2X1_LOC_596/Y NAND2X1_LOC_454/Y 0.08fF
C63628 NAND2X1_LOC_821/a_36_24# INVX1_LOC_160/A 0.01fF
C63629 NOR2X1_LOC_759/Y INVX1_LOC_109/Y 0.24fF
C63630 INVX1_LOC_93/Y NOR2X1_LOC_74/A 0.00fF
C63631 NAND2X1_LOC_859/Y INVX1_LOC_118/A 0.03fF
C63632 INVX1_LOC_40/A NAND2X1_LOC_92/a_36_24# 0.00fF
C63633 INVX1_LOC_64/A NAND2X1_LOC_794/B 0.07fF
C63634 INVX1_LOC_24/Y NOR2X1_LOC_858/A 0.03fF
C63635 NOR2X1_LOC_32/B NAND2X1_LOC_571/Y 0.47fF
C63636 NAND2X1_LOC_783/Y NAND2X1_LOC_175/Y 0.05fF
C63637 INVX1_LOC_135/A NAND2X1_LOC_849/B 0.10fF
C63638 INPUT_0 INVX1_LOC_11/Y 0.06fF
C63639 INVX1_LOC_210/Y NOR2X1_LOC_227/A 0.01fF
C63640 NOR2X1_LOC_802/A NOR2X1_LOC_814/A 0.07fF
C63641 INVX1_LOC_135/A INVX1_LOC_38/A 0.03fF
C63642 NOR2X1_LOC_328/Y NOR2X1_LOC_695/a_36_216# 0.00fF
C63643 NAND2X1_LOC_571/B NOR2X1_LOC_92/Y 0.09fF
C63644 INVX1_LOC_177/A NAND2X1_LOC_475/Y 0.03fF
C63645 INVX1_LOC_90/A NOR2X1_LOC_813/Y 0.00fF
C63646 INVX1_LOC_25/Y NAND2X1_LOC_243/B 0.16fF
C63647 INVX1_LOC_93/Y NOR2X1_LOC_9/Y 0.10fF
C63648 INVX1_LOC_103/A INVX1_LOC_57/A 0.07fF
C63649 INVX1_LOC_208/Y NOR2X1_LOC_155/A 0.12fF
C63650 NOR2X1_LOC_340/Y INVX1_LOC_29/A 0.02fF
C63651 NOR2X1_LOC_142/Y INVX1_LOC_29/A 0.08fF
C63652 NOR2X1_LOC_790/B NOR2X1_LOC_793/A 0.10fF
C63653 INVX1_LOC_295/A INVX1_LOC_38/A 0.05fF
C63654 D_INPUT_1 NAND2X1_LOC_192/B 0.01fF
C63655 NAND2X1_LOC_660/Y NOR2X1_LOC_435/A 0.03fF
C63656 NOR2X1_LOC_137/A INVX1_LOC_9/A 0.02fF
C63657 INVX1_LOC_64/A INVX1_LOC_48/Y 0.02fF
C63658 NOR2X1_LOC_441/Y NOR2X1_LOC_281/Y 0.01fF
C63659 INVX1_LOC_90/A INVX1_LOC_280/A 0.25fF
C63660 INVX1_LOC_90/A NOR2X1_LOC_94/Y 0.43fF
C63661 INVX1_LOC_78/Y NOR2X1_LOC_601/Y 0.02fF
C63662 INVX1_LOC_24/Y INVX1_LOC_292/Y 0.25fF
C63663 NAND2X1_LOC_483/Y NAND2X1_LOC_254/Y 0.91fF
C63664 NAND2X1_LOC_725/A NAND2X1_LOC_579/A 0.10fF
C63665 INVX1_LOC_36/Y NOR2X1_LOC_199/a_36_216# 0.00fF
C63666 NAND2X1_LOC_649/B INVX1_LOC_91/A 0.02fF
C63667 NOR2X1_LOC_419/Y INVX1_LOC_32/A 0.07fF
C63668 INVX1_LOC_292/A INVX1_LOC_57/A 0.00fF
C63669 NAND2X1_LOC_672/B NOR2X1_LOC_814/A 0.02fF
C63670 INVX1_LOC_10/A NAND2X1_LOC_798/B 0.04fF
C63671 NAND2X1_LOC_470/a_36_24# INVX1_LOC_19/A 0.01fF
C63672 NAND2X1_LOC_866/B INVX1_LOC_118/A 0.14fF
C63673 NOR2X1_LOC_78/B INVX1_LOC_186/Y 0.07fF
C63674 NAND2X1_LOC_721/A NOR2X1_LOC_74/A 0.02fF
C63675 INVX1_LOC_5/A NAND2X1_LOC_725/B 0.05fF
C63676 INVX1_LOC_213/Y NOR2X1_LOC_833/B 0.05fF
C63677 NAND2X1_LOC_348/A NOR2X1_LOC_813/Y 0.01fF
C63678 NOR2X1_LOC_121/A INVX1_LOC_84/A 0.03fF
C63679 NOR2X1_LOC_130/A INVX1_LOC_180/Y 0.02fF
C63680 NOR2X1_LOC_716/B INVX1_LOC_32/A 0.17fF
C63681 INVX1_LOC_181/Y INVX1_LOC_78/A 0.03fF
C63682 INVX1_LOC_45/A NOR2X1_LOC_635/B 0.07fF
C63683 NOR2X1_LOC_536/a_36_216# INVX1_LOC_76/A 0.01fF
C63684 NOR2X1_LOC_334/A NOR2X1_LOC_857/A 0.02fF
C63685 NAND2X1_LOC_634/Y NOR2X1_LOC_438/Y 0.02fF
C63686 NAND2X1_LOC_807/Y INVX1_LOC_118/A 0.16fF
C63687 NOR2X1_LOC_78/B NOR2X1_LOC_777/B 0.13fF
C63688 NOR2X1_LOC_655/B INVX1_LOC_29/A 0.01fF
C63689 INVX1_LOC_45/A INVX1_LOC_275/Y 0.00fF
C63690 INVX1_LOC_21/A NAND2X1_LOC_326/A 0.07fF
C63691 INVX1_LOC_45/A NOR2X1_LOC_748/A 0.26fF
C63692 NOR2X1_LOC_188/Y INVX1_LOC_84/A 0.01fF
C63693 INVX1_LOC_22/A NOR2X1_LOC_68/Y 0.02fF
C63694 NOR2X1_LOC_626/Y INVX1_LOC_1/A 0.01fF
C63695 NAND2X1_LOC_348/A INVX1_LOC_280/A 0.13fF
C63696 NOR2X1_LOC_770/Y NAND2X1_LOC_93/B 0.03fF
C63697 NOR2X1_LOC_433/A INVX1_LOC_128/Y 1.37fF
C63698 NOR2X1_LOC_568/A NOR2X1_LOC_748/A 0.36fF
C63699 NOR2X1_LOC_361/B NOR2X1_LOC_791/Y 0.03fF
C63700 INVX1_LOC_64/A INVX1_LOC_246/A 0.07fF
C63701 NOR2X1_LOC_91/A INVX1_LOC_61/A 0.01fF
C63702 NAND2X1_LOC_660/Y INVX1_LOC_63/A 1.53fF
C63703 INVX1_LOC_5/A NAND2X1_LOC_183/a_36_24# 0.01fF
C63704 NOR2X1_LOC_335/A INVX1_LOC_94/Y 0.01fF
C63705 INVX1_LOC_256/Y NOR2X1_LOC_89/A 0.09fF
C63706 INVX1_LOC_58/A NOR2X1_LOC_723/Y 0.03fF
C63707 INVX1_LOC_50/A INVX1_LOC_177/Y 0.63fF
C63708 NOR2X1_LOC_82/A INVX1_LOC_306/Y 1.00fF
C63709 NOR2X1_LOC_770/Y NAND2X1_LOC_425/Y 0.03fF
C63710 NOR2X1_LOC_65/B INVX1_LOC_181/Y 0.00fF
C63711 NOR2X1_LOC_775/Y NOR2X1_LOC_461/A 0.31fF
C63712 NOR2X1_LOC_403/B NAND2X1_LOC_99/A 0.00fF
C63713 NOR2X1_LOC_99/B NOR2X1_LOC_673/B 0.03fF
C63714 INVX1_LOC_50/A NOR2X1_LOC_215/Y 0.06fF
C63715 INVX1_LOC_151/A INVX1_LOC_128/Y 0.03fF
C63716 NOR2X1_LOC_468/Y NOR2X1_LOC_271/B 0.01fF
C63717 INVX1_LOC_25/Y INVX1_LOC_284/A 0.84fF
C63718 INVX1_LOC_61/A INVX1_LOC_23/A 0.07fF
C63719 D_INPUT_0 INVX1_LOC_63/A 3.03fF
C63720 INVX1_LOC_18/A INVX1_LOC_53/A 0.17fF
C63721 INVX1_LOC_98/Y INVX1_LOC_32/A 0.01fF
C63722 NAND2X1_LOC_79/Y NAND2X1_LOC_205/A 0.03fF
C63723 NOR2X1_LOC_574/a_36_216# INVX1_LOC_21/Y 0.00fF
C63724 NOR2X1_LOC_186/Y NAND2X1_LOC_337/a_36_24# 0.01fF
C63725 INVX1_LOC_48/A INVX1_LOC_9/A 0.42fF
C63726 INVX1_LOC_6/A INVX1_LOC_118/A 0.43fF
C63727 INVX1_LOC_298/Y NOR2X1_LOC_142/Y 0.07fF
C63728 INVX1_LOC_77/A NOR2X1_LOC_383/B 5.24fF
C63729 NOR2X1_LOC_272/Y NOR2X1_LOC_276/Y 0.09fF
C63730 D_INPUT_1 NAND2X1_LOC_656/A 0.11fF
C63731 INVX1_LOC_39/A INVX1_LOC_31/A 0.06fF
C63732 NOR2X1_LOC_554/B INVX1_LOC_68/A 0.04fF
C63733 INVX1_LOC_83/A NOR2X1_LOC_777/B 0.06fF
C63734 INVX1_LOC_162/A NOR2X1_LOC_318/A 0.05fF
C63735 NAND2X1_LOC_466/A NOR2X1_LOC_449/A 0.03fF
C63736 NAND2X1_LOC_571/B NAND2X1_LOC_837/Y 0.04fF
C63737 NAND2X1_LOC_856/A NOR2X1_LOC_304/Y 0.03fF
C63738 INVX1_LOC_69/Y NOR2X1_LOC_640/Y 0.02fF
C63739 NOR2X1_LOC_637/Y INVX1_LOC_53/A 0.01fF
C63740 NOR2X1_LOC_99/B INVX1_LOC_29/A 0.08fF
C63741 NOR2X1_LOC_552/A INVX1_LOC_38/A 0.07fF
C63742 NOR2X1_LOC_510/Y INVX1_LOC_30/A 0.07fF
C63743 INVX1_LOC_174/A INVX1_LOC_1/A 2.21fF
C63744 NOR2X1_LOC_226/A NOR2X1_LOC_80/Y 0.23fF
C63745 INVX1_LOC_292/A NAND2X1_LOC_312/a_36_24# 0.00fF
C63746 INVX1_LOC_41/A NOR2X1_LOC_858/A 0.08fF
C63747 NOR2X1_LOC_815/Y INVX1_LOC_23/A 0.01fF
C63748 INVX1_LOC_172/A INVX1_LOC_53/A 0.04fF
C63749 NAND2X1_LOC_579/A NOR2X1_LOC_372/A 0.01fF
C63750 INVX1_LOC_272/Y NOR2X1_LOC_679/Y 0.01fF
C63751 NOR2X1_LOC_486/Y NOR2X1_LOC_331/B 0.07fF
C63752 NOR2X1_LOC_272/Y INVX1_LOC_136/A 0.01fF
C63753 INVX1_LOC_41/A NOR2X1_LOC_828/a_36_216# 0.00fF
C63754 INPUT_0 NOR2X1_LOC_179/Y 0.01fF
C63755 INVX1_LOC_50/A INVX1_LOC_104/A 0.34fF
C63756 NAND2X1_LOC_562/Y INVX1_LOC_23/A 0.37fF
C63757 NAND2X1_LOC_740/Y INVX1_LOC_300/Y 0.17fF
C63758 NOR2X1_LOC_128/B NOR2X1_LOC_554/A 0.15fF
C63759 NOR2X1_LOC_34/A INVX1_LOC_205/A 0.14fF
C63760 NOR2X1_LOC_78/A NOR2X1_LOC_78/Y 0.01fF
C63761 NOR2X1_LOC_598/B NOR2X1_LOC_551/B 0.26fF
C63762 INVX1_LOC_124/A NOR2X1_LOC_383/B 0.07fF
C63763 NAND2X1_LOC_639/A INVX1_LOC_37/A 0.01fF
C63764 NAND2X1_LOC_67/Y NOR2X1_LOC_717/Y 0.04fF
C63765 INVX1_LOC_49/A NOR2X1_LOC_109/Y 0.94fF
C63766 INVX1_LOC_64/A INVX1_LOC_231/Y 0.15fF
C63767 NOR2X1_LOC_91/A NAND2X1_LOC_733/B 0.52fF
C63768 INVX1_LOC_182/A INVX1_LOC_29/A 0.23fF
C63769 NOR2X1_LOC_717/B INVX1_LOC_32/A 0.03fF
C63770 INVX1_LOC_2/A INVX1_LOC_270/A 0.11fF
C63771 NOR2X1_LOC_536/A INVX1_LOC_37/A 0.15fF
C63772 NAND2X1_LOC_214/Y NOR2X1_LOC_554/B 0.03fF
C63773 NOR2X1_LOC_160/B NOR2X1_LOC_785/A 0.04fF
C63774 INVX1_LOC_213/Y NOR2X1_LOC_598/B 1.94fF
C63775 NOR2X1_LOC_411/A NOR2X1_LOC_413/Y 0.06fF
C63776 INVX1_LOC_64/A NOR2X1_LOC_413/a_36_216# 0.00fF
C63777 INVX1_LOC_139/Y INVX1_LOC_38/A 0.02fF
C63778 NAND2X1_LOC_13/a_36_24# NOR2X1_LOC_641/B 0.00fF
C63779 NOR2X1_LOC_45/B NOR2X1_LOC_841/A 0.10fF
C63780 INVX1_LOC_299/A INVX1_LOC_305/A 0.03fF
C63781 NOR2X1_LOC_216/B NAND2X1_LOC_642/Y 0.01fF
C63782 NOR2X1_LOC_270/Y NOR2X1_LOC_122/A 0.03fF
C63783 NOR2X1_LOC_457/B NOR2X1_LOC_666/A 0.04fF
C63784 INVX1_LOC_25/Y NOR2X1_LOC_134/a_36_216# 0.01fF
C63785 INVX1_LOC_2/A NOR2X1_LOC_416/A 0.23fF
C63786 NOR2X1_LOC_355/A NAND2X1_LOC_647/B 0.05fF
C63787 INVX1_LOC_35/A INVX1_LOC_76/Y 0.03fF
C63788 NOR2X1_LOC_813/Y NAND2X1_LOC_849/B 0.03fF
C63789 NOR2X1_LOC_130/Y INVX1_LOC_32/A 0.02fF
C63790 NOR2X1_LOC_859/Y NOR2X1_LOC_865/A 0.04fF
C63791 INVX1_LOC_64/A NOR2X1_LOC_629/a_36_216# 0.00fF
C63792 NAND2X1_LOC_72/Y INVX1_LOC_104/A 0.01fF
C63793 INVX1_LOC_93/A NAND2X1_LOC_640/Y 0.00fF
C63794 INVX1_LOC_75/A INVX1_LOC_284/A 0.07fF
C63795 NOR2X1_LOC_667/A NAND2X1_LOC_784/A 0.47fF
C63796 NAND2X1_LOC_493/Y NAND2X1_LOC_837/Y 0.09fF
C63797 NOR2X1_LOC_152/A INVX1_LOC_38/A 0.04fF
C63798 NOR2X1_LOC_636/B NOR2X1_LOC_68/A 0.09fF
C63799 NAND2X1_LOC_784/A INVX1_LOC_248/A 0.00fF
C63800 INVX1_LOC_64/A NOR2X1_LOC_84/Y 1.23fF
C63801 NOR2X1_LOC_689/a_36_216# NAND2X1_LOC_863/B 0.00fF
C63802 INVX1_LOC_135/A NAND2X1_LOC_223/A 0.03fF
C63803 NOR2X1_LOC_537/Y NOR2X1_LOC_392/Y 0.07fF
C63804 NOR2X1_LOC_685/A NAND2X1_LOC_782/B 0.16fF
C63805 NOR2X1_LOC_687/Y NOR2X1_LOC_383/B 0.03fF
C63806 NAND2X1_LOC_787/A INVX1_LOC_280/Y 0.03fF
C63807 NAND2X1_LOC_9/Y NOR2X1_LOC_346/B 0.15fF
C63808 INVX1_LOC_225/Y NOR2X1_LOC_703/B 0.10fF
C63809 NAND2X1_LOC_30/Y NAND2X1_LOC_587/a_36_24# 0.00fF
C63810 INVX1_LOC_38/A INVX1_LOC_280/A 0.02fF
C63811 INVX1_LOC_37/A NAND2X1_LOC_93/B 0.04fF
C63812 INVX1_LOC_35/Y NAND2X1_LOC_464/A 0.17fF
C63813 INVX1_LOC_2/A NOR2X1_LOC_109/Y 0.14fF
C63814 NAND2X1_LOC_35/Y NOR2X1_LOC_822/Y 0.03fF
C63815 NOR2X1_LOC_263/a_36_216# NOR2X1_LOC_652/Y 0.01fF
C63816 INVX1_LOC_11/A NOR2X1_LOC_13/Y 0.07fF
C63817 NOR2X1_LOC_653/B NAND2X1_LOC_357/B 0.02fF
C63818 NOR2X1_LOC_96/Y INVX1_LOC_280/A 0.12fF
C63819 NOR2X1_LOC_549/a_36_216# NOR2X1_LOC_383/B 0.00fF
C63820 INVX1_LOC_24/Y NAND2X1_LOC_361/Y 0.10fF
C63821 NOR2X1_LOC_151/Y INVX1_LOC_32/A 0.03fF
C63822 NOR2X1_LOC_94/Y NOR2X1_LOC_96/Y 0.17fF
C63823 NAND2X1_LOC_735/B INVX1_LOC_23/A 0.00fF
C63824 VDD INVX1_LOC_113/A 0.00fF
C63825 INVX1_LOC_37/A NAND2X1_LOC_425/Y 0.06fF
C63826 NOR2X1_LOC_351/Y NOR2X1_LOC_331/B 0.09fF
C63827 NOR2X1_LOC_137/B NAND2X1_LOC_475/Y 0.10fF
C63828 INVX1_LOC_6/A NAND2X1_LOC_455/B 0.46fF
C63829 NOR2X1_LOC_790/B NOR2X1_LOC_516/B 0.07fF
C63830 INVX1_LOC_83/A NOR2X1_LOC_843/B 0.10fF
C63831 INVX1_LOC_171/A INVX1_LOC_116/Y 0.08fF
C63832 NOR2X1_LOC_498/Y NAND2X1_LOC_493/Y 0.00fF
C63833 INVX1_LOC_21/A NOR2X1_LOC_87/B 0.03fF
C63834 NOR2X1_LOC_76/A INVX1_LOC_26/A 0.07fF
C63835 NOR2X1_LOC_186/Y INVX1_LOC_54/Y 0.06fF
C63836 NOR2X1_LOC_156/Y INVX1_LOC_117/A 0.03fF
C63837 INVX1_LOC_61/A INVX1_LOC_31/A 2.81fF
C63838 NOR2X1_LOC_536/A NOR2X1_LOC_743/Y 0.30fF
C63839 INVX1_LOC_145/Y INVX1_LOC_270/Y 0.00fF
C63840 NOR2X1_LOC_92/Y NAND2X1_LOC_799/Y 0.01fF
C63841 INVX1_LOC_233/A INVX1_LOC_22/A 0.18fF
C63842 INVX1_LOC_287/A INVX1_LOC_83/A 0.07fF
C63843 NOR2X1_LOC_400/B INVX1_LOC_89/A 0.02fF
C63844 NAND2X1_LOC_624/B INVX1_LOC_16/A 0.00fF
C63845 INVX1_LOC_284/Y INVX1_LOC_24/A 0.07fF
C63846 INVX1_LOC_64/A INVX1_LOC_290/A 0.10fF
C63847 INVX1_LOC_218/A INVX1_LOC_50/Y 0.01fF
C63848 NOR2X1_LOC_798/A NOR2X1_LOC_175/B 0.00fF
C63849 INPUT_3 NOR2X1_LOC_419/Y 0.11fF
C63850 NAND2X1_LOC_848/Y INVX1_LOC_280/A -0.01fF
C63851 INVX1_LOC_224/Y INVX1_LOC_89/A 0.03fF
C63852 INVX1_LOC_136/A NAND2X1_LOC_364/A 0.58fF
C63853 NOR2X1_LOC_266/B INVX1_LOC_63/A 0.03fF
C63854 NOR2X1_LOC_134/Y NOR2X1_LOC_237/Y 0.02fF
C63855 NOR2X1_LOC_216/B NOR2X1_LOC_271/Y 0.12fF
C63856 INVX1_LOC_37/A NOR2X1_LOC_661/A 0.05fF
C63857 NOR2X1_LOC_15/Y NOR2X1_LOC_709/A 0.03fF
C63858 NAND2X1_LOC_564/A NOR2X1_LOC_76/A 0.04fF
C63859 INVX1_LOC_214/Y NOR2X1_LOC_173/Y 0.00fF
C63860 INVX1_LOC_45/Y INVX1_LOC_223/A 0.16fF
C63861 INVX1_LOC_212/Y NOR2X1_LOC_160/B 0.07fF
C63862 INVX1_LOC_17/A NOR2X1_LOC_574/A 0.18fF
C63863 INVX1_LOC_136/A NAND2X1_LOC_100/a_36_24# 0.00fF
C63864 NOR2X1_LOC_74/A INVX1_LOC_87/A 0.08fF
C63865 INVX1_LOC_73/A INVX1_LOC_26/A 0.07fF
C63866 NOR2X1_LOC_295/Y INVX1_LOC_150/Y 0.04fF
C63867 NOR2X1_LOC_798/A INVX1_LOC_22/A 0.21fF
C63868 NOR2X1_LOC_815/Y INVX1_LOC_31/A 0.01fF
C63869 NOR2X1_LOC_667/A NAND2X1_LOC_326/A 0.10fF
C63870 INVX1_LOC_256/A NOR2X1_LOC_799/a_36_216# 0.01fF
C63871 NOR2X1_LOC_658/Y NOR2X1_LOC_433/A 0.07fF
C63872 NOR2X1_LOC_569/Y INVX1_LOC_50/Y 0.03fF
C63873 INVX1_LOC_87/Y INVX1_LOC_29/Y 0.01fF
C63874 NAND2X1_LOC_488/a_36_24# INVX1_LOC_92/A 0.01fF
C63875 NOR2X1_LOC_358/a_36_216# NOR2X1_LOC_364/A 0.03fF
C63876 NOR2X1_LOC_857/A NAND2X1_LOC_74/B 0.10fF
C63877 NOR2X1_LOC_9/Y INVX1_LOC_87/A 0.05fF
C63878 INVX1_LOC_36/A INVX1_LOC_49/A 11.62fF
C63879 NOR2X1_LOC_624/A INVX1_LOC_31/A 0.07fF
C63880 NOR2X1_LOC_457/A INVX1_LOC_177/A 0.06fF
C63881 INVX1_LOC_21/A INVX1_LOC_174/Y 0.01fF
C63882 INVX1_LOC_225/A NAND2X1_LOC_337/a_36_24# 0.01fF
C63883 NAND2X1_LOC_848/A INVX1_LOC_63/A 0.03fF
C63884 NOR2X1_LOC_808/A NOR2X1_LOC_807/B 0.03fF
C63885 NOR2X1_LOC_791/Y NAND2X1_LOC_573/A 0.09fF
C63886 INVX1_LOC_306/A INVX1_LOC_306/Y 0.01fF
C63887 INVX1_LOC_269/A NOR2X1_LOC_382/a_36_216# 0.01fF
C63888 NAND2X1_LOC_538/Y NAND2X1_LOC_840/B 0.07fF
C63889 NOR2X1_LOC_176/Y INVX1_LOC_29/A 0.11fF
C63890 NOR2X1_LOC_590/A NOR2X1_LOC_802/A 0.20fF
C63891 INPUT_1 NOR2X1_LOC_109/Y 0.03fF
C63892 NOR2X1_LOC_797/a_36_216# INVX1_LOC_213/A 0.01fF
C63893 NOR2X1_LOC_588/A NOR2X1_LOC_30/Y 0.35fF
C63894 INVX1_LOC_266/A NOR2X1_LOC_569/Y 0.01fF
C63895 INVX1_LOC_14/A NOR2X1_LOC_719/A 0.10fF
C63896 NAND2X1_LOC_622/a_36_24# INVX1_LOC_253/Y 0.00fF
C63897 NOR2X1_LOC_658/Y NOR2X1_LOC_52/B 0.55fF
C63898 INVX1_LOC_1/A NOR2X1_LOC_589/A 0.26fF
C63899 INVX1_LOC_46/Y NAND2X1_LOC_609/a_36_24# 0.01fF
C63900 NOR2X1_LOC_13/Y NOR2X1_LOC_433/A 0.10fF
C63901 INVX1_LOC_145/A INVX1_LOC_49/A 0.10fF
C63902 NOR2X1_LOC_607/a_36_216# INVX1_LOC_77/A 0.00fF
C63903 NOR2X1_LOC_500/A NOR2X1_LOC_374/A 0.03fF
C63904 INVX1_LOC_1/A NAND2X1_LOC_377/Y 0.00fF
C63905 NOR2X1_LOC_208/Y INVX1_LOC_49/A 0.01fF
C63906 INVX1_LOC_57/Y NAND2X1_LOC_650/a_36_24# 0.06fF
C63907 INVX1_LOC_11/A NOR2X1_LOC_146/Y 0.10fF
C63908 INVX1_LOC_30/A INVX1_LOC_177/A 0.06fF
C63909 INVX1_LOC_50/A INVX1_LOC_206/Y 0.03fF
C63910 NOR2X1_LOC_175/A NOR2X1_LOC_500/B 0.37fF
C63911 INVX1_LOC_14/A NOR2X1_LOC_561/Y 0.08fF
C63912 INVX1_LOC_14/A INVX1_LOC_7/A 5.88fF
C63913 NOR2X1_LOC_68/A NAND2X1_LOC_116/A 0.88fF
C63914 NOR2X1_LOC_815/a_36_216# NAND2X1_LOC_593/Y 0.01fF
C63915 NOR2X1_LOC_668/a_36_216# INPUT_0 0.00fF
C63916 NAND2X1_LOC_447/Y NAND2X1_LOC_454/Y 0.32fF
C63917 INVX1_LOC_2/A INVX1_LOC_36/A 0.19fF
C63918 INVX1_LOC_136/A NAND2X1_LOC_785/A 0.06fF
C63919 INVX1_LOC_36/A NOR2X1_LOC_818/Y 0.24fF
C63920 INVX1_LOC_83/A NAND2X1_LOC_216/a_36_24# 0.01fF
C63921 NAND2X1_LOC_9/Y INVX1_LOC_100/A 0.00fF
C63922 NOR2X1_LOC_804/B INVX1_LOC_49/A 0.29fF
C63923 NOR2X1_LOC_226/A INVX1_LOC_36/A 3.86fF
C63924 INVX1_LOC_233/A INVX1_LOC_100/A 0.07fF
C63925 INVX1_LOC_78/A INVX1_LOC_115/A 0.58fF
C63926 NAND2X1_LOC_175/B NOR2X1_LOC_433/A 1.38fF
C63927 NOR2X1_LOC_441/Y INVX1_LOC_151/Y 0.00fF
C63928 INVX1_LOC_45/A NOR2X1_LOC_524/a_36_216# 0.00fF
C63929 INVX1_LOC_1/A INVX1_LOC_171/A 2.32fF
C63930 INVX1_LOC_117/A D_INPUT_5 0.07fF
C63931 INVX1_LOC_225/A NOR2X1_LOC_303/Y 0.09fF
C63932 NOR2X1_LOC_13/Y NOR2X1_LOC_52/B 0.01fF
C63933 NOR2X1_LOC_65/B NOR2X1_LOC_675/A 0.04fF
C63934 INVX1_LOC_41/A NAND2X1_LOC_361/Y 0.14fF
C63935 INVX1_LOC_50/A NOR2X1_LOC_600/Y 0.39fF
C63936 NOR2X1_LOC_78/B INVX1_LOC_18/A 0.13fF
C63937 INVX1_LOC_37/A NAND2X1_LOC_470/B 0.02fF
C63938 INVX1_LOC_12/A NOR2X1_LOC_433/Y 0.13fF
C63939 NAND2X1_LOC_860/A INVX1_LOC_98/A 0.12fF
C63940 NOR2X1_LOC_388/Y INVX1_LOC_33/A 0.19fF
C63941 NOR2X1_LOC_309/Y INVX1_LOC_49/A 0.03fF
C63942 INVX1_LOC_239/A NOR2X1_LOC_19/B 0.00fF
C63943 NAND2X1_LOC_588/a_36_24# INVX1_LOC_18/A 0.01fF
C63944 NOR2X1_LOC_557/Y NOR2X1_LOC_561/a_36_216# 0.01fF
C63945 NOR2X1_LOC_178/a_36_216# NAND2X1_LOC_93/B 0.00fF
C63946 INVX1_LOC_34/A NAND2X1_LOC_276/Y 0.03fF
C63947 INVX1_LOC_36/A NOR2X1_LOC_218/Y 0.16fF
C63948 NAND2X1_LOC_860/A NOR2X1_LOC_78/A 0.07fF
C63949 INVX1_LOC_89/A NOR2X1_LOC_103/Y 0.07fF
C63950 NAND2X1_LOC_46/a_36_24# INVX1_LOC_315/Y 0.00fF
C63951 NAND2X1_LOC_301/a_36_24# NOR2X1_LOC_596/A 0.00fF
C63952 NAND2X1_LOC_72/Y INVX1_LOC_206/Y 0.00fF
C63953 INVX1_LOC_2/A NOR2X1_LOC_208/Y 0.08fF
C63954 INVX1_LOC_17/A INVX1_LOC_47/A 0.03fF
C63955 INVX1_LOC_72/A INVX1_LOC_25/Y 0.18fF
C63956 NOR2X1_LOC_454/Y NOR2X1_LOC_163/Y 0.05fF
C63957 INVX1_LOC_290/A NOR2X1_LOC_585/a_36_216# 0.01fF
C63958 INVX1_LOC_12/A NAND2X1_LOC_798/B 0.17fF
C63959 NAND2X1_LOC_326/A NAND2X1_LOC_327/a_36_24# 0.01fF
C63960 NAND2X1_LOC_194/a_36_24# NOR2X1_LOC_360/Y 0.01fF
C63961 NAND2X1_LOC_579/A NAND2X1_LOC_560/A 0.02fF
C63962 INVX1_LOC_2/A NOR2X1_LOC_237/Y 0.01fF
C63963 NAND2X1_LOC_175/B NOR2X1_LOC_52/B 0.07fF
C63964 NOR2X1_LOC_68/A INVX1_LOC_232/A 0.85fF
C63965 INVX1_LOC_57/A INVX1_LOC_143/Y 0.03fF
C63966 INVX1_LOC_64/A NOR2X1_LOC_41/a_36_216# 0.01fF
C63967 NOR2X1_LOC_15/Y NAND2X1_LOC_863/A 0.10fF
C63968 INVX1_LOC_136/A NOR2X1_LOC_86/A 0.34fF
C63969 NOR2X1_LOC_524/a_36_216# INVX1_LOC_71/A 0.00fF
C63970 NOR2X1_LOC_559/B INVX1_LOC_218/A 0.18fF
C63971 INVX1_LOC_25/A INVX1_LOC_20/A 0.10fF
C63972 INVX1_LOC_280/A NAND2X1_LOC_223/A 0.07fF
C63973 INVX1_LOC_45/A INVX1_LOC_150/A 0.01fF
C63974 INVX1_LOC_116/A NOR2X1_LOC_211/A 0.01fF
C63975 INVX1_LOC_41/Y INVX1_LOC_16/A 0.02fF
C63976 NOR2X1_LOC_160/B NOR2X1_LOC_702/Y 0.06fF
C63977 INVX1_LOC_45/A NOR2X1_LOC_110/a_36_216# 0.00fF
C63978 NOR2X1_LOC_220/B INVX1_LOC_91/A 0.05fF
C63979 NOR2X1_LOC_252/Y NOR2X1_LOC_238/Y 0.01fF
C63980 NOR2X1_LOC_617/Y INVX1_LOC_16/A -0.02fF
C63981 D_INPUT_3 INVX1_LOC_23/A 0.27fF
C63982 INVX1_LOC_225/A INVX1_LOC_54/Y 0.20fF
C63983 INVX1_LOC_34/A NAND2X1_LOC_374/Y 0.07fF
C63984 INVX1_LOC_45/A INVX1_LOC_89/A 0.57fF
C63985 INVX1_LOC_38/A NOR2X1_LOC_541/B 0.02fF
C63986 NOR2X1_LOC_590/A NOR2X1_LOC_174/A 0.05fF
C63987 NOR2X1_LOC_655/B INVX1_LOC_8/A 0.10fF
C63988 INVX1_LOC_14/Y INVX1_LOC_23/A 0.11fF
C63989 INVX1_LOC_1/A NAND2X1_LOC_821/a_36_24# 0.01fF
C63990 INVX1_LOC_2/A NOR2X1_LOC_309/Y 0.00fF
C63991 INVX1_LOC_89/A NOR2X1_LOC_568/A 0.03fF
C63992 INVX1_LOC_83/A INVX1_LOC_18/A 1.03fF
C63993 INVX1_LOC_245/Y NOR2X1_LOC_742/A 0.02fF
C63994 INVX1_LOC_14/A NOR2X1_LOC_167/Y 0.02fF
C63995 NOR2X1_LOC_844/A NOR2X1_LOC_87/Y 0.11fF
C63996 INVX1_LOC_93/A NAND2X1_LOC_642/Y 0.00fF
C63997 NOR2X1_LOC_351/Y NOR2X1_LOC_449/A 0.05fF
C63998 NOR2X1_LOC_82/A NOR2X1_LOC_74/A 0.01fF
C63999 INVX1_LOC_36/A INPUT_1 0.04fF
C64000 NOR2X1_LOC_226/A NOR2X1_LOC_309/Y 0.21fF
C64001 INVX1_LOC_178/A NAND2X1_LOC_655/A 0.10fF
C64002 INVX1_LOC_11/A NOR2X1_LOC_337/A 0.00fF
C64003 INVX1_LOC_295/A NAND2X1_LOC_386/a_36_24# 0.01fF
C64004 NAND2X1_LOC_564/B NOR2X1_LOC_716/B 0.05fF
C64005 NOR2X1_LOC_78/A NAND2X1_LOC_473/A 0.02fF
C64006 INVX1_LOC_33/A NAND2X1_LOC_479/Y 0.01fF
C64007 INVX1_LOC_24/A NOR2X1_LOC_525/Y 0.34fF
C64008 INVX1_LOC_59/Y INVX1_LOC_306/Y 0.02fF
C64009 INVX1_LOC_24/A NAND2X1_LOC_809/A 0.02fF
C64010 NOR2X1_LOC_82/A NOR2X1_LOC_9/Y 0.14fF
C64011 INVX1_LOC_71/A INVX1_LOC_150/A 0.10fF
C64012 NOR2X1_LOC_1/Y INPUT_7 0.03fF
C64013 INVX1_LOC_83/A NOR2X1_LOC_713/B 0.08fF
C64014 NOR2X1_LOC_383/B INVX1_LOC_9/A 0.18fF
C64015 INVX1_LOC_280/Y NAND2X1_LOC_722/A 0.07fF
C64016 NOR2X1_LOC_78/B INVX1_LOC_34/Y 0.16fF
C64017 NOR2X1_LOC_673/A NOR2X1_LOC_38/B 0.03fF
C64018 INVX1_LOC_89/A INVX1_LOC_71/A 0.03fF
C64019 INVX1_LOC_247/Y INVX1_LOC_182/A 0.02fF
C64020 NOR2X1_LOC_250/Y NOR2X1_LOC_318/B 0.03fF
C64021 INVX1_LOC_75/A INVX1_LOC_72/A 0.17fF
C64022 VDD NOR2X1_LOC_460/Y 0.12fF
C64023 INVX1_LOC_135/A INVX1_LOC_33/A 0.06fF
C64024 NOR2X1_LOC_718/a_36_216# INVX1_LOC_22/A 0.01fF
C64025 NAND2X1_LOC_741/B NOR2X1_LOC_2/Y 0.01fF
C64026 INVX1_LOC_28/A INVX1_LOC_41/Y 0.03fF
C64027 INVX1_LOC_256/A NAND2X1_LOC_329/a_36_24# 0.06fF
C64028 NAND2X1_LOC_402/a_36_24# INVX1_LOC_42/A 0.00fF
C64029 INVX1_LOC_16/Y INVX1_LOC_123/Y 0.17fF
C64030 NOR2X1_LOC_237/Y INPUT_1 0.07fF
C64031 NAND2X1_LOC_338/B INVX1_LOC_25/Y 0.04fF
C64032 INVX1_LOC_225/Y INVX1_LOC_91/A 0.10fF
C64033 NAND2X1_LOC_114/B NOR2X1_LOC_557/A 0.07fF
C64034 INVX1_LOC_50/Y NAND2X1_LOC_472/Y 0.07fF
C64035 INVX1_LOC_295/A INVX1_LOC_33/A 0.04fF
C64036 NOR2X1_LOC_617/Y INVX1_LOC_28/A 0.02fF
C64037 INVX1_LOC_17/A INVX1_LOC_95/Y 0.03fF
C64038 INVX1_LOC_1/A INVX1_LOC_20/A 0.03fF
C64039 NOR2X1_LOC_816/A NAND2X1_LOC_655/A 0.09fF
C64040 INVX1_LOC_206/A NOR2X1_LOC_543/A 0.13fF
C64041 INVX1_LOC_28/A NAND2X1_LOC_593/Y 0.32fF
C64042 NOR2X1_LOC_808/A NOR2X1_LOC_811/A 0.26fF
C64043 INVX1_LOC_47/Y INVX1_LOC_12/A 0.09fF
C64044 INVX1_LOC_14/A INVX1_LOC_76/A 0.17fF
C64045 NAND2X1_LOC_359/Y INVX1_LOC_156/Y 0.20fF
C64046 INVX1_LOC_118/A NOR2X1_LOC_109/Y 0.10fF
C64047 INVX1_LOC_191/Y INPUT_5 0.03fF
C64048 NAND2X1_LOC_206/B INVX1_LOC_15/A 0.03fF
C64049 INVX1_LOC_77/A NOR2X1_LOC_163/Y 0.03fF
C64050 NAND2X1_LOC_660/a_36_24# NAND2X1_LOC_477/A 0.06fF
C64051 NAND2X1_LOC_63/Y NOR2X1_LOC_80/Y 0.01fF
C64052 NAND2X1_LOC_205/A INVX1_LOC_123/Y 0.06fF
C64053 NOR2X1_LOC_431/Y INVX1_LOC_144/A 0.03fF
C64054 INVX1_LOC_164/Y INVX1_LOC_164/A 0.04fF
C64055 NOR2X1_LOC_309/Y INPUT_1 0.03fF
C64056 INVX1_LOC_23/Y NAND2X1_LOC_768/Y 0.01fF
C64057 INVX1_LOC_135/A NOR2X1_LOC_521/a_36_216# 0.01fF
C64058 INVX1_LOC_14/A NAND2X1_LOC_84/a_36_24# 0.01fF
C64059 NOR2X1_LOC_355/A NAND2X1_LOC_342/Y 0.00fF
C64060 NAND2X1_LOC_785/A NAND2X1_LOC_862/Y 0.03fF
C64061 NOR2X1_LOC_843/B NOR2X1_LOC_68/Y 0.03fF
C64062 INVX1_LOC_285/A INVX1_LOC_29/Y 0.17fF
C64063 INVX1_LOC_24/A NOR2X1_LOC_391/Y -0.00fF
C64064 INVX1_LOC_124/Y INVX1_LOC_93/Y 0.01fF
C64065 INVX1_LOC_49/A NOR2X1_LOC_208/A 0.01fF
C64066 INVX1_LOC_232/Y NOR2X1_LOC_130/A 0.01fF
C64067 NOR2X1_LOC_68/A NOR2X1_LOC_685/A 0.02fF
C64068 NOR2X1_LOC_401/B NOR2X1_LOC_123/B 0.01fF
C64069 NOR2X1_LOC_86/A NAND2X1_LOC_849/a_36_24# 0.00fF
C64070 INVX1_LOC_30/A INVX1_LOC_65/A 0.01fF
C64071 NOR2X1_LOC_91/Y NOR2X1_LOC_528/Y 0.01fF
C64072 INVX1_LOC_251/Y INVX1_LOC_90/A 0.03fF
C64073 INVX1_LOC_256/A INVX1_LOC_37/A 0.08fF
C64074 INVX1_LOC_29/Y NOR2X1_LOC_814/A 0.03fF
C64075 NOR2X1_LOC_658/Y INVX1_LOC_199/A 0.01fF
C64076 NOR2X1_LOC_637/a_36_216# INVX1_LOC_144/A 0.01fF
C64077 NOR2X1_LOC_766/a_36_216# INVX1_LOC_20/A 0.00fF
C64078 INVX1_LOC_135/A INVX1_LOC_40/A 0.07fF
C64079 NOR2X1_LOC_328/Y INVX1_LOC_10/A 0.02fF
C64080 INVX1_LOC_136/A NOR2X1_LOC_405/A 0.13fF
C64081 INVX1_LOC_161/Y NOR2X1_LOC_139/a_36_216# 0.00fF
C64082 INVX1_LOC_78/A NOR2X1_LOC_114/Y 0.09fF
C64083 INVX1_LOC_30/A NOR2X1_LOC_137/B 0.01fF
C64084 NOR2X1_LOC_516/B NOR2X1_LOC_128/B 0.01fF
C64085 INVX1_LOC_13/A NOR2X1_LOC_391/A 0.03fF
C64086 NAND2X1_LOC_276/Y INPUT_0 0.28fF
C64087 NOR2X1_LOC_700/Y INVX1_LOC_22/A 0.03fF
C64088 INVX1_LOC_110/Y VDD -0.00fF
C64089 NAND2X1_LOC_392/A NOR2X1_LOC_130/A 0.02fF
C64090 INVX1_LOC_31/A D_INPUT_3 0.23fF
C64091 NOR2X1_LOC_717/Y INVX1_LOC_76/A 0.07fF
C64092 INVX1_LOC_33/A NOR2X1_LOC_711/A 0.01fF
C64093 D_INPUT_0 INVX1_LOC_1/Y 0.00fF
C64094 NOR2X1_LOC_384/Y INVX1_LOC_20/A 0.25fF
C64095 INVX1_LOC_36/A NOR2X1_LOC_586/Y 0.10fF
C64096 NOR2X1_LOC_382/Y VDD 0.16fF
C64097 INVX1_LOC_5/A NOR2X1_LOC_66/Y 0.01fF
C64098 NOR2X1_LOC_65/B NOR2X1_LOC_114/Y 0.07fF
C64099 INVX1_LOC_282/A NOR2X1_LOC_482/Y 0.05fF
C64100 NAND2X1_LOC_338/B INVX1_LOC_75/A 0.03fF
C64101 INVX1_LOC_72/A NAND2X1_LOC_453/A 0.05fF
C64102 INVX1_LOC_5/A NOR2X1_LOC_820/B 0.10fF
C64103 NAND2X1_LOC_783/A NAND2X1_LOC_779/a_36_24# 0.00fF
C64104 NOR2X1_LOC_476/Y VDD 0.24fF
C64105 NOR2X1_LOC_172/Y NOR2X1_LOC_45/B 0.45fF
C64106 NAND2X1_LOC_729/Y INVX1_LOC_20/A 0.02fF
C64107 INVX1_LOC_18/A INVX1_LOC_46/A 1.31fF
C64108 INVX1_LOC_50/Y NAND2X1_LOC_206/Y 0.07fF
C64109 NAND2X1_LOC_739/B INVX1_LOC_76/A 0.01fF
C64110 INVX1_LOC_33/A NOR2X1_LOC_552/A 0.03fF
C64111 INVX1_LOC_11/A NOR2X1_LOC_640/Y 0.01fF
C64112 NOR2X1_LOC_667/A NOR2X1_LOC_527/Y 0.02fF
C64113 NAND2X1_LOC_714/B INVX1_LOC_84/A 4.51fF
C64114 NOR2X1_LOC_441/Y INVX1_LOC_118/Y 0.03fF
C64115 INVX1_LOC_256/A NOR2X1_LOC_743/Y 0.06fF
C64116 INVX1_LOC_278/Y NOR2X1_LOC_74/A 0.08fF
C64117 INVX1_LOC_111/A INVX1_LOC_14/Y 0.00fF
C64118 NAND2X1_LOC_711/B INVX1_LOC_46/A 0.03fF
C64119 INVX1_LOC_89/A NOR2X1_LOC_749/Y 0.00fF
C64120 NOR2X1_LOC_360/Y INVX1_LOC_117/A 0.07fF
C64121 INVX1_LOC_113/Y INVX1_LOC_115/A 0.01fF
C64122 NAND2X1_LOC_811/Y INVX1_LOC_11/Y 0.03fF
C64123 NOR2X1_LOC_218/A NOR2X1_LOC_155/A 0.01fF
C64124 INVX1_LOC_58/A D_INPUT_5 0.02fF
C64125 NAND2X1_LOC_387/B INVX1_LOC_38/A 0.02fF
C64126 INVX1_LOC_266/Y INVX1_LOC_91/A 0.02fF
C64127 NAND2X1_LOC_391/Y INVX1_LOC_19/A 0.03fF
C64128 NAND2X1_LOC_84/Y NAND2X1_LOC_84/a_36_24# 0.00fF
C64129 INVX1_LOC_172/A INVX1_LOC_46/A 0.03fF
C64130 NOR2X1_LOC_791/Y NAND2X1_LOC_81/B 0.05fF
C64131 NOR2X1_LOC_15/Y INVX1_LOC_294/A 0.26fF
C64132 NOR2X1_LOC_298/Y INVX1_LOC_140/A 0.05fF
C64133 NAND2X1_LOC_123/Y NAND2X1_LOC_656/Y 0.14fF
C64134 INVX1_LOC_25/A INVX1_LOC_4/A 0.27fF
C64135 INVX1_LOC_36/A INVX1_LOC_118/A 7.78fF
C64136 NAND2X1_LOC_198/B NOR2X1_LOC_536/A 0.03fF
C64137 NAND2X1_LOC_462/B NOR2X1_LOC_19/Y 0.01fF
C64138 NOR2X1_LOC_298/Y NAND2X1_LOC_463/B 0.01fF
C64139 INVX1_LOC_54/Y NAND2X1_LOC_642/Y 0.00fF
C64140 INVX1_LOC_83/A INVX1_LOC_31/Y 0.06fF
C64141 INVX1_LOC_221/A INVX1_LOC_20/A 0.03fF
C64142 INVX1_LOC_123/A NOR2X1_LOC_121/A 0.01fF
C64143 NOR2X1_LOC_576/B NAND2X1_LOC_863/A 0.33fF
C64144 NOR2X1_LOC_355/A INVX1_LOC_67/Y 0.02fF
C64145 NOR2X1_LOC_439/B INVX1_LOC_313/Y 0.00fF
C64146 NAND2X1_LOC_354/B NAND2X1_LOC_687/A 0.04fF
C64147 NAND2X1_LOC_363/B INVX1_LOC_4/Y 0.01fF
C64148 NAND2X1_LOC_538/Y INVX1_LOC_49/Y 0.04fF
C64149 INVX1_LOC_75/A INVX1_LOC_313/Y 0.10fF
C64150 INVX1_LOC_7/A INVX1_LOC_48/A 0.52fF
C64151 INVX1_LOC_33/A INVX1_LOC_10/Y 0.03fF
C64152 NOR2X1_LOC_368/A NOR2X1_LOC_76/A 0.44fF
C64153 INVX1_LOC_171/A NOR2X1_LOC_188/A 0.18fF
C64154 NOR2X1_LOC_250/A INVX1_LOC_49/Y 0.34fF
C64155 NOR2X1_LOC_237/Y INVX1_LOC_118/A 0.27fF
C64156 NAND2X1_LOC_197/a_36_24# NOR2X1_LOC_435/A 0.00fF
C64157 NOR2X1_LOC_245/a_36_216# INVX1_LOC_286/A 0.00fF
C64158 NOR2X1_LOC_677/Y INVX1_LOC_57/A 0.04fF
C64159 NAND2X1_LOC_9/Y NOR2X1_LOC_843/B 0.07fF
C64160 NAND2X1_LOC_842/B INVX1_LOC_100/A 0.00fF
C64161 INVX1_LOC_122/A INVX1_LOC_210/A 0.23fF
C64162 INVX1_LOC_276/A NAND2X1_LOC_685/a_36_24# 0.00fF
C64163 D_INPUT_0 NOR2X1_LOC_318/B 0.12fF
C64164 INVX1_LOC_49/A NOR2X1_LOC_435/A 0.03fF
C64165 NOR2X1_LOC_593/Y NOR2X1_LOC_640/Y 0.02fF
C64166 NOR2X1_LOC_645/a_36_216# INVX1_LOC_84/A 0.02fF
C64167 INVX1_LOC_224/Y NOR2X1_LOC_392/Y 0.02fF
C64168 NOR2X1_LOC_309/Y INVX1_LOC_118/A 0.09fF
C64169 NAND2X1_LOC_7/Y NOR2X1_LOC_197/B 0.10fF
C64170 NOR2X1_LOC_657/a_36_216# NAND2X1_LOC_454/Y 0.01fF
C64171 INVX1_LOC_1/A INVX1_LOC_4/A 0.06fF
C64172 D_INPUT_0 INVX1_LOC_93/Y 0.02fF
C64173 INVX1_LOC_1/Y NOR2X1_LOC_266/B 0.06fF
C64174 NOR2X1_LOC_91/Y NAND2X1_LOC_477/Y 0.03fF
C64175 NOR2X1_LOC_442/a_36_216# NOR2X1_LOC_623/B 0.02fF
C64176 INVX1_LOC_90/A NOR2X1_LOC_45/B 3.21fF
C64177 NAND2X1_LOC_564/B NAND2X1_LOC_633/Y 0.07fF
C64178 NOR2X1_LOC_521/a_36_216# INVX1_LOC_280/A 0.00fF
C64179 NOR2X1_LOC_594/a_36_216# NOR2X1_LOC_594/Y 0.00fF
C64180 INVX1_LOC_36/Y NOR2X1_LOC_195/a_36_216# 0.00fF
C64181 INVX1_LOC_35/A D_INPUT_1 0.65fF
C64182 NOR2X1_LOC_15/Y NAND2X1_LOC_444/B 0.01fF
C64183 INVX1_LOC_36/A NAND2X1_LOC_63/Y 0.03fF
C64184 INPUT_0 NOR2X1_LOC_184/a_36_216# 0.00fF
C64185 INVX1_LOC_17/Y NAND2X1_LOC_35/Y 0.03fF
C64186 NOR2X1_LOC_703/B INVX1_LOC_19/A 0.01fF
C64187 INVX1_LOC_138/A NOR2X1_LOC_416/A 0.03fF
C64188 NOR2X1_LOC_15/Y NOR2X1_LOC_334/Y 0.05fF
C64189 NOR2X1_LOC_186/Y NAND2X1_LOC_286/B 0.04fF
C64190 NOR2X1_LOC_433/A NOR2X1_LOC_697/Y 0.12fF
C64191 NOR2X1_LOC_690/Y INVX1_LOC_46/A 0.03fF
C64192 INVX1_LOC_97/A INVX1_LOC_247/A 0.02fF
C64193 NOR2X1_LOC_216/a_36_216# NOR2X1_LOC_318/B 0.00fF
C64194 INVX1_LOC_222/A NOR2X1_LOC_188/A 0.09fF
C64195 INVX1_LOC_233/Y NAND2X1_LOC_787/A 0.03fF
C64196 INVX1_LOC_40/A INVX1_LOC_280/A 0.01fF
C64197 INVX1_LOC_222/A NOR2X1_LOC_548/B 0.01fF
C64198 INVX1_LOC_90/A INVX1_LOC_247/A 0.03fF
C64199 INVX1_LOC_53/Y NOR2X1_LOC_536/A 0.56fF
C64200 NOR2X1_LOC_32/B NAND2X1_LOC_725/A 0.07fF
C64201 INVX1_LOC_140/A NAND2X1_LOC_655/A 0.03fF
C64202 NOR2X1_LOC_457/A INVX1_LOC_4/Y 0.43fF
C64203 NAND2X1_LOC_30/Y NAND2X1_LOC_452/Y 0.50fF
C64204 INVX1_LOC_298/Y NOR2X1_LOC_187/Y 0.02fF
C64205 NOR2X1_LOC_312/Y NOR2X1_LOC_280/Y 0.18fF
C64206 NAND2X1_LOC_573/Y NAND2X1_LOC_286/B 0.02fF
C64207 NOR2X1_LOC_130/A NAND2X1_LOC_287/B 0.07fF
C64208 INVX1_LOC_49/A INVX1_LOC_63/A 0.03fF
C64209 INVX1_LOC_2/A NOR2X1_LOC_435/A 0.02fF
C64210 INVX1_LOC_256/A NAND2X1_LOC_72/B 0.07fF
C64211 NOR2X1_LOC_91/A NAND2X1_LOC_303/Y 0.21fF
C64212 D_INPUT_0 NAND2X1_LOC_721/A 0.01fF
C64213 NOR2X1_LOC_52/B NOR2X1_LOC_697/Y 0.06fF
C64214 NOR2X1_LOC_131/A NOR2X1_LOC_155/A 0.01fF
C64215 INVX1_LOC_50/A NOR2X1_LOC_92/Y 0.49fF
C64216 NOR2X1_LOC_471/Y INVX1_LOC_271/Y 0.07fF
C64217 INVX1_LOC_35/A NOR2X1_LOC_108/a_36_216# 0.00fF
C64218 NOR2X1_LOC_7/Y INVX1_LOC_6/A 0.14fF
C64219 NAND2X1_LOC_67/Y NOR2X1_LOC_383/B 0.19fF
C64220 INVX1_LOC_249/Y INVX1_LOC_84/A 0.09fF
C64221 NOR2X1_LOC_100/A NOR2X1_LOC_243/B 0.01fF
C64222 NAND2X1_LOC_321/a_36_24# NOR2X1_LOC_334/Y 0.01fF
C64223 INVX1_LOC_21/A INVX1_LOC_58/Y 0.08fF
C64224 NOR2X1_LOC_15/Y NAND2X1_LOC_464/B 0.10fF
C64225 NAND2X1_LOC_571/B NAND2X1_LOC_571/Y 0.02fF
C64226 INVX1_LOC_16/A INVX1_LOC_185/A 0.03fF
C64227 NOR2X1_LOC_6/B NAND2X1_LOC_206/Y 0.05fF
C64228 INVX1_LOC_45/Y INVX1_LOC_290/Y 0.10fF
C64229 INVX1_LOC_53/Y NAND2X1_LOC_93/B 0.07fF
C64230 NOR2X1_LOC_61/B INVX1_LOC_152/Y 0.09fF
C64231 NAND2X1_LOC_357/B NOR2X1_LOC_605/A 0.01fF
C64232 INVX1_LOC_30/A INVX1_LOC_4/Y 0.07fF
C64233 NAND2X1_LOC_564/B INVX1_LOC_71/Y 0.01fF
C64234 INVX1_LOC_125/Y INVX1_LOC_91/A 0.46fF
C64235 INPUT_1 NOR2X1_LOC_102/a_36_216# 0.00fF
C64236 INVX1_LOC_157/A INVX1_LOC_157/Y 0.02fF
C64237 NAND2X1_LOC_364/A NAND2X1_LOC_647/B 0.02fF
C64238 NOR2X1_LOC_665/A NAND2X1_LOC_93/B 0.07fF
C64239 NOR2X1_LOC_464/B NOR2X1_LOC_678/A 0.01fF
C64240 NOR2X1_LOC_273/Y INVX1_LOC_15/A 0.02fF
C64241 INVX1_LOC_2/A INVX1_LOC_63/A 1.97fF
C64242 NOR2X1_LOC_92/Y NAND2X1_LOC_544/a_36_24# 0.00fF
C64243 NOR2X1_LOC_818/Y INVX1_LOC_63/A 0.03fF
C64244 NAND2X1_LOC_660/Y INVX1_LOC_117/Y 0.00fF
C64245 NOR2X1_LOC_759/Y INVX1_LOC_15/A 0.02fF
C64246 INVX1_LOC_6/A NAND2X1_LOC_212/Y 0.01fF
C64247 INVX1_LOC_90/A NOR2X1_LOC_378/Y 0.01fF
C64248 NOR2X1_LOC_443/Y NOR2X1_LOC_160/B 0.01fF
C64249 INPUT_5 NOR2X1_LOC_36/a_36_216# 0.00fF
C64250 INVX1_LOC_202/A INVX1_LOC_15/A 0.00fF
C64251 NOR2X1_LOC_226/A INVX1_LOC_63/A 0.07fF
C64252 INVX1_LOC_64/A INVX1_LOC_1/A 0.08fF
C64253 NAND2X1_LOC_35/Y NAND2X1_LOC_493/Y 0.08fF
C64254 NOR2X1_LOC_500/Y INVX1_LOC_220/A 0.01fF
C64255 NOR2X1_LOC_567/B INVX1_LOC_117/A 0.08fF
C64256 NOR2X1_LOC_191/a_36_216# INVX1_LOC_93/Y 0.01fF
C64257 NOR2X1_LOC_629/B INVX1_LOC_284/A 0.05fF
C64258 INVX1_LOC_25/A INVX1_LOC_43/Y 0.03fF
C64259 NAND2X1_LOC_198/B NAND2X1_LOC_470/B 0.03fF
C64260 NOR2X1_LOC_178/Y INVX1_LOC_14/A 0.65fF
C64261 NOR2X1_LOC_550/B INVX1_LOC_15/A 0.10fF
C64262 INVX1_LOC_48/A INVX1_LOC_76/A 0.04fF
C64263 D_GATE_366 INVX1_LOC_54/A 0.03fF
C64264 NOR2X1_LOC_590/A INVX1_LOC_29/Y 0.03fF
C64265 INVX1_LOC_6/A INVX1_LOC_14/Y 0.03fF
C64266 NOR2X1_LOC_565/A NOR2X1_LOC_383/B 0.01fF
C64267 INVX1_LOC_69/Y INVX1_LOC_37/A 0.08fF
C64268 NOR2X1_LOC_186/Y NAND2X1_LOC_537/Y 0.00fF
C64269 INVX1_LOC_89/A NOR2X1_LOC_592/B 0.01fF
C64270 INVX1_LOC_49/A NAND2X1_LOC_452/Y 0.02fF
C64271 INVX1_LOC_64/A NOR2X1_LOC_794/B 0.01fF
C64272 INVX1_LOC_28/A INVX1_LOC_185/A 0.06fF
C64273 NAND2X1_LOC_341/a_36_24# INVX1_LOC_29/A 0.01fF
C64274 INVX1_LOC_91/Y INVX1_LOC_38/A 0.09fF
C64275 NAND2X1_LOC_354/Y NOR2X1_LOC_654/A 0.02fF
C64276 NOR2X1_LOC_68/A INVX1_LOC_112/Y 0.01fF
C64277 NOR2X1_LOC_208/Y NOR2X1_LOC_631/Y 0.01fF
C64278 NOR2X1_LOC_113/B NOR2X1_LOC_536/A 0.02fF
C64279 NAND2X1_LOC_351/A INVX1_LOC_57/A 0.01fF
C64280 NOR2X1_LOC_612/a_36_216# NOR2X1_LOC_89/A 0.00fF
C64281 NOR2X1_LOC_160/B INVX1_LOC_213/A 0.07fF
C64282 NOR2X1_LOC_6/B NOR2X1_LOC_297/A 0.04fF
C64283 NOR2X1_LOC_332/A NOR2X1_LOC_820/B 0.02fF
C64284 INVX1_LOC_96/A NAND2X1_LOC_472/Y 0.03fF
C64285 NOR2X1_LOC_355/A NOR2X1_LOC_814/A 0.00fF
C64286 INVX1_LOC_93/Y NOR2X1_LOC_266/B 0.01fF
C64287 NOR2X1_LOC_328/Y INVX1_LOC_12/A 0.08fF
C64288 INVX1_LOC_58/A NOR2X1_LOC_360/Y 0.07fF
C64289 INVX1_LOC_233/Y INVX1_LOC_30/A 0.03fF
C64290 NAND2X1_LOC_79/Y NAND2X1_LOC_215/A 0.03fF
C64291 INVX1_LOC_21/A NAND2X1_LOC_783/Y 0.01fF
C64292 NOR2X1_LOC_605/a_36_216# NOR2X1_LOC_89/A 0.00fF
C64293 INVX1_LOC_233/A INVX1_LOC_18/A 0.07fF
C64294 NOR2X1_LOC_562/B INVX1_LOC_44/A 0.15fF
C64295 NOR2X1_LOC_294/Y NAND2X1_LOC_207/a_36_24# 0.00fF
C64296 NOR2X1_LOC_637/A INVX1_LOC_53/A 0.01fF
C64297 INVX1_LOC_5/A NOR2X1_LOC_500/B 0.01fF
C64298 NOR2X1_LOC_607/A INVX1_LOC_53/A 0.01fF
C64299 INPUT_1 INVX1_LOC_63/A 0.08fF
C64300 NOR2X1_LOC_45/B INVX1_LOC_38/A 0.19fF
C64301 NOR2X1_LOC_757/A NOR2X1_LOC_89/A 0.01fF
C64302 NOR2X1_LOC_91/A NOR2X1_LOC_690/A 0.07fF
C64303 NAND2X1_LOC_832/Y INVX1_LOC_179/A 0.06fF
C64304 NOR2X1_LOC_280/Y NAND2X1_LOC_287/B 0.06fF
C64305 INVX1_LOC_223/Y INVX1_LOC_45/A 0.03fF
C64306 INVX1_LOC_201/Y NAND2X1_LOC_23/a_36_24# 0.02fF
C64307 INVX1_LOC_41/A INVX1_LOC_50/A 0.06fF
C64308 INVX1_LOC_225/A NAND2X1_LOC_286/B 0.01fF
C64309 INVX1_LOC_1/A INVX1_LOC_43/Y 0.01fF
C64310 INVX1_LOC_286/A INVX1_LOC_70/A 0.09fF
C64311 INVX1_LOC_39/A INVX1_LOC_36/A 0.03fF
C64312 INVX1_LOC_136/A NAND2X1_LOC_740/Y 0.01fF
C64313 NOR2X1_LOC_639/a_36_216# NOR2X1_LOC_584/Y 0.00fF
C64314 NOR2X1_LOC_498/Y INVX1_LOC_50/A 0.05fF
C64315 INVX1_LOC_88/A NOR2X1_LOC_816/A 0.02fF
C64316 INVX1_LOC_35/A D_INPUT_2 0.26fF
C64317 NOR2X1_LOC_298/Y INVX1_LOC_42/A 0.19fF
C64318 INVX1_LOC_247/A INVX1_LOC_38/A 0.04fF
C64319 NOR2X1_LOC_45/B NOR2X1_LOC_51/A 0.19fF
C64320 INVX1_LOC_77/A NOR2X1_LOC_405/Y 0.01fF
C64321 INVX1_LOC_233/A INVX1_LOC_172/A 0.07fF
C64322 NOR2X1_LOC_690/A INVX1_LOC_23/A 0.00fF
C64323 INVX1_LOC_93/A NOR2X1_LOC_91/Y 0.16fF
C64324 NOR2X1_LOC_817/a_36_216# INPUT_3 0.00fF
C64325 NAND2X1_LOC_571/a_36_24# NOR2X1_LOC_92/Y 0.01fF
C64326 NOR2X1_LOC_391/A INVX1_LOC_32/A 0.01fF
C64327 NOR2X1_LOC_413/Y INVX1_LOC_23/A 0.01fF
C64328 NOR2X1_LOC_795/Y NAND2X1_LOC_279/a_36_24# 0.06fF
C64329 NAND2X1_LOC_796/B NOR2X1_LOC_68/A 0.23fF
C64330 INVX1_LOC_50/A NAND2X1_LOC_477/A 0.01fF
C64331 NOR2X1_LOC_19/B NAND2X1_LOC_82/Y 0.77fF
C64332 VDD INVX1_LOC_202/Y 0.26fF
C64333 NAND2X1_LOC_35/Y NOR2X1_LOC_495/Y 0.01fF
C64334 INVX1_LOC_24/A INVX1_LOC_50/Y 0.10fF
C64335 NOR2X1_LOC_770/Y NOR2X1_LOC_89/A 0.01fF
C64336 INVX1_LOC_2/A NOR2X1_LOC_65/Y 0.01fF
C64337 NOR2X1_LOC_78/A NOR2X1_LOC_461/A 0.03fF
C64338 NAND2X1_LOC_181/Y INVX1_LOC_26/A 0.03fF
C64339 NOR2X1_LOC_647/A NOR2X1_LOC_78/B 0.02fF
C64340 INVX1_LOC_21/A NOR2X1_LOC_609/A 0.04fF
C64341 NAND2X1_LOC_703/Y INVX1_LOC_18/A 0.07fF
C64342 NAND2X1_LOC_863/B NOR2X1_LOC_409/B 0.03fF
C64343 NAND2X1_LOC_852/Y NOR2X1_LOC_829/A 0.03fF
C64344 NAND2X1_LOC_794/B INVX1_LOC_41/Y 0.02fF
C64345 INVX1_LOC_303/A INVX1_LOC_5/A 0.13fF
C64346 NAND2X1_LOC_555/Y INVX1_LOC_252/Y 0.03fF
C64347 NOR2X1_LOC_644/A INVX1_LOC_290/Y 0.41fF
C64348 INVX1_LOC_5/A NOR2X1_LOC_672/Y 0.23fF
C64349 INVX1_LOC_214/A NOR2X1_LOC_654/A 0.01fF
C64350 NOR2X1_LOC_657/Y INVX1_LOC_103/A 0.01fF
C64351 INVX1_LOC_226/Y INVX1_LOC_23/Y 1.38fF
C64352 INVX1_LOC_179/Y NOR2X1_LOC_383/B 0.02fF
C64353 NOR2X1_LOC_577/Y NOR2X1_LOC_674/Y 0.04fF
C64354 NAND2X1_LOC_149/Y NOR2X1_LOC_257/a_36_216# 0.01fF
C64355 NOR2X1_LOC_56/Y INVX1_LOC_180/Y 0.01fF
C64356 NOR2X1_LOC_667/A NOR2X1_LOC_654/A 0.11fF
C64357 NOR2X1_LOC_288/A NOR2X1_LOC_634/Y 0.03fF
C64358 NOR2X1_LOC_769/a_36_216# INVX1_LOC_296/A 0.01fF
C64359 INVX1_LOC_248/A NOR2X1_LOC_654/A 0.10fF
C64360 INVX1_LOC_21/A NOR2X1_LOC_419/Y 0.03fF
C64361 NOR2X1_LOC_726/Y NOR2X1_LOC_307/A 0.01fF
C64362 NAND2X1_LOC_392/a_36_24# INVX1_LOC_71/A 0.00fF
C64363 INPUT_0 INVX1_LOC_125/A 0.02fF
C64364 INVX1_LOC_41/A NOR2X1_LOC_590/Y 0.19fF
C64365 NOR2X1_LOC_506/Y NAND2X1_LOC_453/A 0.03fF
C64366 INVX1_LOC_266/A INVX1_LOC_24/A 0.07fF
C64367 NAND2X1_LOC_9/Y INVX1_LOC_34/Y 0.02fF
C64368 INVX1_LOC_21/A NOR2X1_LOC_716/B 0.17fF
C64369 INVX1_LOC_174/A NAND2X1_LOC_3/a_36_24# 0.01fF
C64370 INVX1_LOC_236/Y INVX1_LOC_286/Y 0.00fF
C64371 INVX1_LOC_224/Y INVX1_LOC_25/Y 0.11fF
C64372 INVX1_LOC_50/A NOR2X1_LOC_211/A 0.03fF
C64373 NOR2X1_LOC_810/A NOR2X1_LOC_863/B 0.01fF
C64374 INVX1_LOC_233/Y NAND2X1_LOC_722/A 0.06fF
C64375 D_INPUT_0 INVX1_LOC_87/A 0.03fF
C64376 NAND2X1_LOC_733/A NAND2X1_LOC_733/Y 0.06fF
C64377 NOR2X1_LOC_114/A INVX1_LOC_19/A 0.00fF
C64378 INVX1_LOC_56/Y INVX1_LOC_57/A 0.03fF
C64379 NOR2X1_LOC_76/A NAND2X1_LOC_471/Y 0.01fF
C64380 VDD INVX1_LOC_180/Y 0.26fF
C64381 NOR2X1_LOC_824/A NAND2X1_LOC_483/Y 0.02fF
C64382 INVX1_LOC_38/A NOR2X1_LOC_378/Y 0.02fF
C64383 NOR2X1_LOC_124/A NOR2X1_LOC_813/a_36_216# 0.00fF
C64384 INVX1_LOC_89/A NAND2X1_LOC_467/a_36_24# 0.00fF
C64385 NOR2X1_LOC_92/Y NOR2X1_LOC_679/B 0.01fF
C64386 NAND2X1_LOC_787/A NAND2X1_LOC_862/A 0.00fF
C64387 NOR2X1_LOC_15/Y INVX1_LOC_209/Y 0.03fF
C64388 INVX1_LOC_91/A INVX1_LOC_19/A 14.03fF
C64389 NOR2X1_LOC_501/B INVX1_LOC_29/A 0.00fF
C64390 INVX1_LOC_256/A NAND2X1_LOC_368/a_36_24# 0.00fF
C64391 INVX1_LOC_89/A NOR2X1_LOC_621/B 0.01fF
C64392 NAND2X1_LOC_337/B NOR2X1_LOC_758/a_36_216# 0.00fF
C64393 INVX1_LOC_16/A NOR2X1_LOC_754/Y 0.07fF
C64394 INVX1_LOC_25/Y NAND2X1_LOC_793/B 0.01fF
C64395 INVX1_LOC_34/A NOR2X1_LOC_140/A 0.02fF
C64396 NOR2X1_LOC_220/A NAND2X1_LOC_406/a_36_24# 0.00fF
C64397 INVX1_LOC_286/A INVX1_LOC_102/A 0.18fF
C64398 NOR2X1_LOC_142/a_36_216# INVX1_LOC_54/A 0.02fF
C64399 NOR2X1_LOC_124/A NAND2X1_LOC_773/B 0.02fF
C64400 NOR2X1_LOC_127/Y INVX1_LOC_76/A 0.16fF
C64401 INVX1_LOC_122/A NOR2X1_LOC_259/B 0.21fF
C64402 INVX1_LOC_143/A INVX1_LOC_50/Y 0.10fF
C64403 NAND2X1_LOC_725/Y INVX1_LOC_229/Y 3.52fF
C64404 INVX1_LOC_10/A NOR2X1_LOC_484/a_36_216# 0.02fF
C64405 NAND2X1_LOC_76/a_36_24# NOR2X1_LOC_596/A 0.01fF
C64406 INVX1_LOC_227/A INVX1_LOC_29/Y 0.08fF
C64407 NOR2X1_LOC_15/Y NOR2X1_LOC_718/B 0.03fF
C64408 NOR2X1_LOC_272/Y NAND2X1_LOC_342/Y 0.22fF
C64409 INVX1_LOC_21/A INVX1_LOC_98/Y 0.02fF
C64410 NOR2X1_LOC_826/Y NAND2X1_LOC_859/Y 0.02fF
C64411 INVX1_LOC_246/A NAND2X1_LOC_593/Y 0.01fF
C64412 NOR2X1_LOC_188/A INVX1_LOC_4/A 0.04fF
C64413 NOR2X1_LOC_111/A INVX1_LOC_285/A 0.01fF
C64414 NOR2X1_LOC_589/A NOR2X1_LOC_129/a_36_216# 0.00fF
C64415 INVX1_LOC_254/A INVX1_LOC_31/A 0.02fF
C64416 INVX1_LOC_179/A INVX1_LOC_9/A 0.03fF
C64417 NAND2X1_LOC_655/A INVX1_LOC_42/A 0.07fF
C64418 INVX1_LOC_54/A INVX1_LOC_70/A 0.10fF
C64419 INVX1_LOC_34/A NOR2X1_LOC_530/Y 0.08fF
C64420 NAND2X1_LOC_214/B NOR2X1_LOC_789/A 0.02fF
C64421 NOR2X1_LOC_78/B NOR2X1_LOC_321/Y 0.03fF
C64422 INVX1_LOC_95/A INVX1_LOC_102/A 0.09fF
C64423 NOR2X1_LOC_629/Y INVX1_LOC_260/A 0.16fF
C64424 INVX1_LOC_299/A INVX1_LOC_196/A 0.05fF
C64425 INVX1_LOC_28/A INVX1_LOC_270/Y 0.17fF
C64426 NOR2X1_LOC_750/A NAND2X1_LOC_215/A 0.01fF
C64427 NOR2X1_LOC_703/a_36_216# NOR2X1_LOC_551/B 0.00fF
C64428 INVX1_LOC_174/A NAND2X1_LOC_163/a_36_24# 0.00fF
C64429 INVX1_LOC_69/Y NAND2X1_LOC_72/B 0.03fF
C64430 NOR2X1_LOC_690/A INVX1_LOC_31/A 0.03fF
C64431 NOR2X1_LOC_400/B INVX1_LOC_75/A 0.06fF
C64432 INVX1_LOC_27/A NOR2X1_LOC_789/A 0.02fF
C64433 INVX1_LOC_72/A NOR2X1_LOC_577/Y 0.17fF
C64434 NAND2X1_LOC_798/B INVX1_LOC_92/A 0.07fF
C64435 NOR2X1_LOC_523/B NOR2X1_LOC_860/B 0.01fF
C64436 INVX1_LOC_298/A INVX1_LOC_83/A 0.00fF
C64437 INVX1_LOC_19/A NOR2X1_LOC_698/Y 0.06fF
C64438 NOR2X1_LOC_287/A INVX1_LOC_299/A 0.02fF
C64439 INVX1_LOC_224/Y INVX1_LOC_75/A 0.07fF
C64440 NOR2X1_LOC_590/A INVX1_LOC_60/Y 0.30fF
C64441 NOR2X1_LOC_89/A INVX1_LOC_37/A 0.11fF
C64442 NOR2X1_LOC_348/B NOR2X1_LOC_348/a_36_216# 0.00fF
C64443 INVX1_LOC_223/A NOR2X1_LOC_570/B 0.00fF
C64444 NOR2X1_LOC_405/A NAND2X1_LOC_647/B 0.02fF
C64445 NOR2X1_LOC_843/A INVX1_LOC_30/A 0.07fF
C64446 INVX1_LOC_90/A NOR2X1_LOC_53/Y 0.00fF
C64447 NOR2X1_LOC_510/Y NOR2X1_LOC_60/a_36_216# 0.00fF
C64448 INVX1_LOC_298/Y NOR2X1_LOC_501/B 0.28fF
C64449 INVX1_LOC_27/A NAND2X1_LOC_656/Y 0.07fF
C64450 NOR2X1_LOC_78/A NAND2X1_LOC_454/Y 0.01fF
C64451 NOR2X1_LOC_665/A NOR2X1_LOC_348/Y 0.06fF
C64452 INVX1_LOC_45/Y INVX1_LOC_77/A 0.11fF
C64453 INVX1_LOC_21/A NOR2X1_LOC_717/B 0.03fF
C64454 INVX1_LOC_118/A INVX1_LOC_63/A 0.28fF
C64455 NAND2X1_LOC_38/a_36_24# INVX1_LOC_75/A 0.00fF
C64456 NOR2X1_LOC_570/a_36_216# NOR2X1_LOC_388/Y 0.00fF
C64457 NOR2X1_LOC_103/Y INVX1_LOC_25/Y 0.07fF
C64458 INVX1_LOC_13/A INVX1_LOC_269/A 1.65fF
C64459 NAND2X1_LOC_200/B NAND2X1_LOC_114/B 0.10fF
C64460 NAND2X1_LOC_783/Y INVX1_LOC_248/A 0.01fF
C64461 INVX1_LOC_24/A NOR2X1_LOC_718/Y 0.01fF
C64462 NOR2X1_LOC_514/A INVX1_LOC_216/A 0.02fF
C64463 INVX1_LOC_58/A NOR2X1_LOC_427/Y 0.01fF
C64464 NOR2X1_LOC_1/Y INVX1_LOC_38/A 0.01fF
C64465 INVX1_LOC_256/A INVX1_LOC_53/Y 0.24fF
C64466 NAND2X1_LOC_273/a_36_24# NAND2X1_LOC_288/A 0.00fF
C64467 INVX1_LOC_286/A NOR2X1_LOC_280/a_36_216# 0.00fF
C64468 NAND2X1_LOC_557/Y INVX1_LOC_309/A -0.00fF
C64469 NAND2X1_LOC_222/A INVX1_LOC_315/Y 0.01fF
C64470 NOR2X1_LOC_272/Y NOR2X1_LOC_246/Y 0.08fF
C64471 NAND2X1_LOC_468/B INVX1_LOC_78/A 0.03fF
C64472 NOR2X1_LOC_334/Y NOR2X1_LOC_137/a_36_216# 0.00fF
C64473 NOR2X1_LOC_691/A NOR2X1_LOC_634/A 0.09fF
C64474 NOR2X1_LOC_690/A NOR2X1_LOC_617/a_36_216# 0.02fF
C64475 INVX1_LOC_256/A NOR2X1_LOC_665/A 0.07fF
C64476 NOR2X1_LOC_389/A NOR2X1_LOC_210/B 0.10fF
C64477 INVX1_LOC_24/A NOR2X1_LOC_6/B 0.39fF
C64478 NAND2X1_LOC_705/Y NAND2X1_LOC_866/B 0.02fF
C64479 NOR2X1_LOC_588/A INVX1_LOC_296/A 0.45fF
C64480 NAND2X1_LOC_392/Y NAND2X1_LOC_793/Y 0.25fF
C64481 INVX1_LOC_249/A INVX1_LOC_88/Y 0.36fF
C64482 INVX1_LOC_225/Y NOR2X1_LOC_553/B 0.10fF
C64483 NOR2X1_LOC_590/A NOR2X1_LOC_835/A 0.10fF
C64484 NOR2X1_LOC_328/Y NAND2X1_LOC_733/Y 0.68fF
C64485 NAND2X1_LOC_364/A NAND2X1_LOC_342/Y 0.02fF
C64486 NOR2X1_LOC_78/B NAND2X1_LOC_16/Y 0.05fF
C64487 NOR2X1_LOC_51/A NOR2X1_LOC_1/Y 0.03fF
C64488 NOR2X1_LOC_305/a_36_216# NAND2X1_LOC_175/Y 0.01fF
C64489 NOR2X1_LOC_468/Y NOR2X1_LOC_72/a_36_216# 0.01fF
C64490 NAND2X1_LOC_557/Y INVX1_LOC_91/A 0.07fF
C64491 NAND2X1_LOC_67/a_36_24# INVX1_LOC_55/Y 0.01fF
C64492 INVX1_LOC_256/A INVX1_LOC_145/Y 0.01fF
C64493 INVX1_LOC_124/A INVX1_LOC_45/Y 0.10fF
C64494 INVX1_LOC_30/A NAND2X1_LOC_862/A 0.03fF
C64495 INVX1_LOC_102/A INVX1_LOC_54/A 0.07fF
C64496 NOR2X1_LOC_552/A NOR2X1_LOC_748/A 0.10fF
C64497 INVX1_LOC_45/A INVX1_LOC_25/Y 0.62fF
C64498 INVX1_LOC_58/A NOR2X1_LOC_269/Y 0.07fF
C64499 NOR2X1_LOC_82/A D_INPUT_0 5.56fF
C64500 NOR2X1_LOC_500/A NAND2X1_LOC_320/a_36_24# 0.01fF
C64501 INVX1_LOC_21/A NOR2X1_LOC_151/Y 0.46fF
C64502 INVX1_LOC_269/A INVX1_LOC_207/Y 0.01fF
C64503 NOR2X1_LOC_89/A NOR2X1_LOC_743/Y 0.01fF
C64504 INVX1_LOC_41/Y NOR2X1_LOC_482/Y 0.00fF
C64505 INVX1_LOC_230/Y NOR2X1_LOC_719/B 0.03fF
C64506 INVX1_LOC_45/A NAND2X1_LOC_349/B 0.22fF
C64507 NAND2X1_LOC_562/B NOR2X1_LOC_672/Y 0.04fF
C64508 NOR2X1_LOC_92/Y NAND2X1_LOC_652/Y 0.02fF
C64509 NOR2X1_LOC_88/A INVX1_LOC_284/A 0.04fF
C64510 VDD NOR2X1_LOC_278/Y 0.36fF
C64511 INVX1_LOC_84/A INVX1_LOC_293/Y 0.07fF
C64512 INVX1_LOC_17/A NAND2X1_LOC_815/a_36_24# 0.00fF
C64513 INVX1_LOC_234/A INVX1_LOC_39/Y 0.03fF
C64514 INVX1_LOC_72/A INVX1_LOC_22/A 0.22fF
C64515 INVX1_LOC_36/A NAND2X1_LOC_735/B 0.03fF
C64516 NOR2X1_LOC_848/Y NAND2X1_LOC_508/A 0.07fF
C64517 NAND2X1_LOC_860/A NAND2X1_LOC_642/Y 0.13fF
C64518 NOR2X1_LOC_590/A NOR2X1_LOC_355/A 0.42fF
C64519 NOR2X1_LOC_795/Y INVX1_LOC_33/A 0.03fF
C64520 NOR2X1_LOC_383/B INVX1_LOC_76/A 0.07fF
C64521 INVX1_LOC_314/Y INVX1_LOC_256/Y 0.02fF
C64522 NOR2X1_LOC_480/A NOR2X1_LOC_375/Y 0.01fF
C64523 INVX1_LOC_36/A INPUT_5 0.06fF
C64524 VDD NOR2X1_LOC_638/Y 0.26fF
C64525 NAND2X1_LOC_725/Y INVX1_LOC_20/A 0.06fF
C64526 INVX1_LOC_64/A NOR2X1_LOC_43/Y 0.03fF
C64527 NAND2X1_LOC_741/B INVX1_LOC_10/A 0.14fF
C64528 INVX1_LOC_26/A INVX1_LOC_117/A 0.07fF
C64529 INVX1_LOC_34/A NOR2X1_LOC_709/A 0.07fF
C64530 NOR2X1_LOC_405/A NOR2X1_LOC_109/a_36_216# 0.01fF
C64531 NAND2X1_LOC_738/B INVX1_LOC_76/A 0.03fF
C64532 INVX1_LOC_84/A NAND2X1_LOC_74/B 0.10fF
C64533 NAND2X1_LOC_724/Y INVX1_LOC_46/A 11.32fF
C64534 NAND2X1_LOC_784/A INVX1_LOC_20/A 0.01fF
C64535 NOR2X1_LOC_312/Y INVX1_LOC_286/Y 0.04fF
C64536 NOR2X1_LOC_140/A INPUT_0 0.03fF
C64537 NOR2X1_LOC_388/Y NOR2X1_LOC_493/B 0.01fF
C64538 INVX1_LOC_276/A NAND2X1_LOC_325/Y 0.00fF
C64539 INVX1_LOC_71/A INVX1_LOC_25/Y 0.08fF
C64540 INVX1_LOC_292/A NOR2X1_LOC_356/A 0.50fF
C64541 NAND2X1_LOC_63/Y INVX1_LOC_63/A 0.43fF
C64542 NOR2X1_LOC_253/Y NOR2X1_LOC_754/Y 0.08fF
C64543 NOR2X1_LOC_520/A NOR2X1_LOC_340/Y 0.03fF
C64544 INVX1_LOC_47/Y INVX1_LOC_92/A 0.07fF
C64545 NAND2X1_LOC_741/B NOR2X1_LOC_504/a_36_216# 0.03fF
C64546 NOR2X1_LOC_103/Y INVX1_LOC_75/A 0.07fF
C64547 D_INPUT_3 NOR2X1_LOC_416/A 0.01fF
C64548 NAND2X1_LOC_349/B INVX1_LOC_71/A 0.02fF
C64549 INVX1_LOC_83/A INVX1_LOC_205/A 0.04fF
C64550 NOR2X1_LOC_541/Y INVX1_LOC_75/A 0.16fF
C64551 INVX1_LOC_232/Y NOR2X1_LOC_4/a_36_216# 0.00fF
C64552 NOR2X1_LOC_781/B NOR2X1_LOC_781/Y 0.01fF
C64553 INVX1_LOC_157/A NAND2X1_LOC_198/B 0.02fF
C64554 NOR2X1_LOC_614/Y INVX1_LOC_33/A 0.39fF
C64555 NOR2X1_LOC_6/B INVX1_LOC_143/A 0.10fF
C64556 INVX1_LOC_161/Y INVX1_LOC_79/A 0.03fF
C64557 INVX1_LOC_49/A INVX1_LOC_1/Y 0.11fF
C64558 NAND2X1_LOC_724/Y NOR2X1_LOC_766/Y 0.03fF
C64559 INVX1_LOC_108/A NAND2X1_LOC_226/a_36_24# 0.00fF
C64560 D_INPUT_0 NAND2X1_LOC_514/Y 0.01fF
C64561 NOR2X1_LOC_710/B NOR2X1_LOC_711/A 0.01fF
C64562 NAND2X1_LOC_711/B NOR2X1_LOC_700/Y 0.10fF
C64563 NOR2X1_LOC_75/Y INVX1_LOC_311/A 0.00fF
C64564 INVX1_LOC_292/A NOR2X1_LOC_74/A 0.39fF
C64565 INVX1_LOC_45/A NOR2X1_LOC_439/B 0.02fF
C64566 NAND2X1_LOC_842/B INVX1_LOC_18/A 0.02fF
C64567 INVX1_LOC_226/Y NAND2X1_LOC_116/A 0.13fF
C64568 NOR2X1_LOC_690/A NAND2X1_LOC_859/Y 0.01fF
C64569 NAND2X1_LOC_618/Y NOR2X1_LOC_642/a_36_216# 0.00fF
C64570 NOR2X1_LOC_416/A INVX1_LOC_230/A 0.87fF
C64571 NOR2X1_LOC_590/A NOR2X1_LOC_541/a_36_216# 0.00fF
C64572 INVX1_LOC_45/A INVX1_LOC_75/A 2.86fF
C64573 NAND2X1_LOC_338/B NOR2X1_LOC_346/B 0.07fF
C64574 NOR2X1_LOC_106/Y INVX1_LOC_313/A 0.06fF
C64575 NOR2X1_LOC_175/B NOR2X1_LOC_537/Y 0.50fF
C64576 INVX1_LOC_75/A NOR2X1_LOC_568/A 0.58fF
C64577 NAND2X1_LOC_120/a_36_24# INVX1_LOC_6/A 0.00fF
C64578 INVX1_LOC_209/Y NOR2X1_LOC_576/B 0.03fF
C64579 NAND2X1_LOC_538/Y NAND2X1_LOC_649/B 0.09fF
C64580 INVX1_LOC_161/Y INVX1_LOC_91/A 0.07fF
C64581 INVX1_LOC_21/A NAND2X1_LOC_633/Y 0.30fF
C64582 INVX1_LOC_13/A NAND2X1_LOC_127/a_36_24# 0.00fF
C64583 NOR2X1_LOC_589/A NOR2X1_LOC_300/Y 0.02fF
C64584 INVX1_LOC_299/A INVX1_LOC_95/Y 0.00fF
C64585 NOR2X1_LOC_384/Y INVX1_LOC_282/A 0.04fF
C64586 INVX1_LOC_2/A INVX1_LOC_1/Y 0.03fF
C64587 NAND2X1_LOC_549/B INVX1_LOC_316/Y 0.01fF
C64588 NOR2X1_LOC_706/A NOR2X1_LOC_546/A 0.04fF
C64589 NOR2X1_LOC_644/A INVX1_LOC_77/A 0.03fF
C64590 NAND2X1_LOC_326/A INVX1_LOC_20/A 0.62fF
C64591 NOR2X1_LOC_537/Y INVX1_LOC_22/A 0.60fF
C64592 NOR2X1_LOC_620/A INVX1_LOC_29/A 0.03fF
C64593 INVX1_LOC_313/Y NOR2X1_LOC_577/Y 0.00fF
C64594 INVX1_LOC_102/A NOR2X1_LOC_48/B 0.12fF
C64595 NAND2X1_LOC_74/B INVX1_LOC_15/A 0.06fF
C64596 NOR2X1_LOC_577/a_36_216# INVX1_LOC_177/A 0.00fF
C64597 NOR2X1_LOC_226/A INVX1_LOC_1/Y 0.29fF
C64598 INVX1_LOC_57/Y NOR2X1_LOC_167/Y 0.02fF
C64599 NOR2X1_LOC_321/Y INVX1_LOC_46/A 0.07fF
C64600 NOR2X1_LOC_155/A NOR2X1_LOC_858/A 0.02fF
C64601 NAND2X1_LOC_323/B NOR2X1_LOC_325/A 0.03fF
C64602 INVX1_LOC_30/Y INVX1_LOC_143/A 0.01fF
C64603 NOR2X1_LOC_6/B NOR2X1_LOC_130/A 0.05fF
C64604 INVX1_LOC_11/A NOR2X1_LOC_631/B 0.07fF
C64605 NOR2X1_LOC_690/A NAND2X1_LOC_866/B 1.28fF
C64606 NOR2X1_LOC_828/B INVX1_LOC_77/A 0.04fF
C64607 NOR2X1_LOC_831/B INVX1_LOC_57/A 0.19fF
C64608 INVX1_LOC_35/A NOR2X1_LOC_61/Y 0.18fF
C64609 INVX1_LOC_39/A NOR2X1_LOC_102/a_36_216# 0.00fF
C64610 INVX1_LOC_206/A NAND2X1_LOC_656/Y 0.05fF
C64611 NOR2X1_LOC_516/B NOR2X1_LOC_382/a_36_216# 0.00fF
C64612 INVX1_LOC_75/A INVX1_LOC_71/A 0.40fF
C64613 INVX1_LOC_226/Y INVX1_LOC_232/A 0.10fF
C64614 INVX1_LOC_123/Y NAND2X1_LOC_215/A 0.09fF
C64615 INVX1_LOC_13/A NAND2X1_LOC_563/A 0.09fF
C64616 NAND2X1_LOC_149/Y NAND2X1_LOC_639/A 0.02fF
C64617 INVX1_LOC_53/A NAND2X1_LOC_798/B 0.57fF
C64618 INVX1_LOC_267/A INVX1_LOC_135/A 0.03fF
C64619 NOR2X1_LOC_742/A INVX1_LOC_49/A 0.10fF
C64620 NOR2X1_LOC_151/Y NOR2X1_LOC_596/a_36_216# 0.00fF
C64621 NOR2X1_LOC_299/Y INVX1_LOC_209/A 0.07fF
C64622 INVX1_LOC_268/A INVX1_LOC_268/Y 0.06fF
C64623 NOR2X1_LOC_78/B NOR2X1_LOC_686/B 0.07fF
C64624 NAND2X1_LOC_181/Y INVX1_LOC_164/A 0.14fF
C64625 NOR2X1_LOC_15/Y NAND2X1_LOC_472/Y 0.09fF
C64626 INVX1_LOC_313/Y NOR2X1_LOC_348/B 0.02fF
C64627 NOR2X1_LOC_334/Y INVX1_LOC_99/A 0.08fF
C64628 NOR2X1_LOC_756/Y INVX1_LOC_8/A 0.03fF
C64629 INVX1_LOC_50/A INVX1_LOC_136/Y 0.00fF
C64630 NOR2X1_LOC_82/A NOR2X1_LOC_266/B 0.00fF
C64631 NOR2X1_LOC_835/A NAND2X1_LOC_822/a_36_24# 0.00fF
C64632 NAND2X1_LOC_793/Y INVX1_LOC_46/A 0.03fF
C64633 INVX1_LOC_11/A INVX1_LOC_37/A 7.30fF
C64634 NOR2X1_LOC_828/B NOR2X1_LOC_732/A 0.03fF
C64635 INVX1_LOC_166/A INVX1_LOC_203/A 0.01fF
C64636 INVX1_LOC_11/A NOR2X1_LOC_231/A 0.01fF
C64637 INVX1_LOC_34/A NAND2X1_LOC_863/A 0.43fF
C64638 NOR2X1_LOC_251/Y NAND2X1_LOC_656/Y 0.08fF
C64639 NOR2X1_LOC_106/Y INVX1_LOC_6/A 0.06fF
C64640 NAND2X1_LOC_794/B INVX1_LOC_185/A 0.03fF
C64641 NOR2X1_LOC_68/A NOR2X1_LOC_78/A 0.25fF
C64642 NOR2X1_LOC_209/Y INVX1_LOC_85/Y 0.03fF
C64643 INVX1_LOC_269/A INVX1_LOC_66/Y 0.01fF
C64644 NAND2X1_LOC_803/B NOR2X1_LOC_111/A 0.04fF
C64645 NAND2X1_LOC_596/a_36_24# INVX1_LOC_90/A 0.00fF
C64646 NOR2X1_LOC_648/a_36_216# INVX1_LOC_55/Y 0.01fF
C64647 INVX1_LOC_12/A INVX1_LOC_23/Y 0.07fF
C64648 INVX1_LOC_24/A INVX1_LOC_96/A 1.48fF
C64649 INVX1_LOC_78/A NAND2X1_LOC_213/a_36_24# 0.00fF
C64650 NAND2X1_LOC_842/B NOR2X1_LOC_709/a_36_216# 0.00fF
C64651 NOR2X1_LOC_107/Y INVX1_LOC_117/A 0.01fF
C64652 NOR2X1_LOC_626/a_36_216# INVX1_LOC_179/A 0.00fF
C64653 INVX1_LOC_227/A INVX1_LOC_101/A 0.01fF
C64654 INVX1_LOC_236/Y VDD 0.54fF
C64655 NOR2X1_LOC_655/B NOR2X1_LOC_750/A 0.01fF
C64656 INVX1_LOC_284/Y VDD 0.56fF
C64657 INVX1_LOC_90/A NOR2X1_LOC_388/a_36_216# 0.01fF
C64658 NOR2X1_LOC_590/A NOR2X1_LOC_111/A 0.08fF
C64659 NOR2X1_LOC_170/A NAND2X1_LOC_72/B 0.01fF
C64660 NOR2X1_LOC_793/Y NOR2X1_LOC_729/A 1.42fF
C64661 NAND2X1_LOC_149/Y NAND2X1_LOC_93/B 0.07fF
C64662 NOR2X1_LOC_604/Y INVX1_LOC_186/Y 0.01fF
C64663 INVX1_LOC_2/A NOR2X1_LOC_742/A 0.07fF
C64664 INVX1_LOC_45/A NAND2X1_LOC_453/A 0.07fF
C64665 INVX1_LOC_89/A NAND2X1_LOC_479/Y 0.00fF
C64666 INVX1_LOC_36/A D_INPUT_3 0.03fF
C64667 INVX1_LOC_24/A NOR2X1_LOC_124/A 0.08fF
C64668 INVX1_LOC_49/A NOR2X1_LOC_318/B 1.54fF
C64669 NOR2X1_LOC_152/Y NAND2X1_LOC_655/A 0.11fF
C64670 INVX1_LOC_313/Y INVX1_LOC_22/A 0.07fF
C64671 INVX1_LOC_1/Y INPUT_1 0.05fF
C64672 INVX1_LOC_36/A INVX1_LOC_14/Y 0.01fF
C64673 INVX1_LOC_80/A NOR2X1_LOC_332/A 0.00fF
C64674 INPUT_0 NOR2X1_LOC_709/A 0.15fF
C64675 NAND2X1_LOC_149/Y NAND2X1_LOC_425/Y 0.02fF
C64676 NAND2X1_LOC_276/Y INVX1_LOC_125/Y 0.00fF
C64677 INVX1_LOC_26/A INVX1_LOC_3/Y 0.14fF
C64678 NAND2X1_LOC_16/Y INVX1_LOC_46/A 0.23fF
C64679 NOR2X1_LOC_858/A NOR2X1_LOC_833/B 0.00fF
C64680 INVX1_LOC_33/A NOR2X1_LOC_45/B 3.28fF
C64681 INVX1_LOC_122/Y VDD 0.21fF
C64682 INVX1_LOC_135/A NOR2X1_LOC_719/a_36_216# 0.00fF
C64683 NOR2X1_LOC_272/Y INVX1_LOC_285/A 0.10fF
C64684 NOR2X1_LOC_32/B INVX1_LOC_29/A 0.37fF
C64685 NOR2X1_LOC_448/a_36_216# NAND2X1_LOC_93/B 0.00fF
C64686 NOR2X1_LOC_516/B NOR2X1_LOC_564/Y 0.04fF
C64687 INVX1_LOC_49/A INVX1_LOC_93/Y 0.08fF
C64688 NOR2X1_LOC_512/Y INVX1_LOC_76/A 0.03fF
C64689 INVX1_LOC_266/A NOR2X1_LOC_197/B 0.10fF
C64690 INVX1_LOC_108/Y NAND2X1_LOC_207/Y 0.05fF
C64691 INVX1_LOC_278/A NAND2X1_LOC_74/B 0.14fF
C64692 NOR2X1_LOC_152/Y NAND2X1_LOC_468/B 0.03fF
C64693 NAND2X1_LOC_303/Y NAND2X1_LOC_810/B 0.74fF
C64694 NOR2X1_LOC_778/B NOR2X1_LOC_337/A -0.00fF
C64695 INVX1_LOC_11/A NOR2X1_LOC_743/Y 0.04fF
C64696 NOR2X1_LOC_716/B INVX1_LOC_304/A 1.44fF
C64697 NAND2X1_LOC_338/B INVX1_LOC_100/A 0.04fF
C64698 INVX1_LOC_39/A INVX1_LOC_63/A 0.03fF
C64699 NOR2X1_LOC_448/a_36_216# NAND2X1_LOC_425/Y 0.01fF
C64700 NOR2X1_LOC_831/Y NOR2X1_LOC_109/Y 1.68fF
C64701 INVX1_LOC_135/A INVX1_LOC_89/A 0.43fF
C64702 NAND2X1_LOC_116/A NOR2X1_LOC_340/a_36_216# 0.00fF
C64703 NOR2X1_LOC_82/A INVX1_LOC_46/Y 1.51fF
C64704 INVX1_LOC_295/A INVX1_LOC_89/A 0.14fF
C64705 NOR2X1_LOC_446/A INVX1_LOC_307/A 0.01fF
C64706 NOR2X1_LOC_641/B INVX1_LOC_9/A 0.07fF
C64707 NOR2X1_LOC_208/Y INVX1_LOC_14/Y 0.10fF
C64708 INVX1_LOC_162/Y INVX1_LOC_95/A 0.12fF
C64709 INVX1_LOC_135/A NAND2X1_LOC_508/A 0.03fF
C64710 NOR2X1_LOC_52/Y INVX1_LOC_38/A 0.04fF
C64711 NAND2X1_LOC_7/Y VDD -0.00fF
C64712 INVX1_LOC_89/A NOR2X1_LOC_560/A 0.00fF
C64713 INVX1_LOC_2/A NOR2X1_LOC_318/B 0.07fF
C64714 NOR2X1_LOC_433/A INVX1_LOC_37/A 0.07fF
C64715 NOR2X1_LOC_772/B INVX1_LOC_42/A 1.49fF
C64716 NAND2X1_LOC_170/A NOR2X1_LOC_167/Y 0.11fF
C64717 NOR2X1_LOC_751/Y INVX1_LOC_9/A 0.03fF
C64718 INVX1_LOC_53/A INVX1_LOC_47/Y 0.14fF
C64719 INVX1_LOC_223/A INVX1_LOC_54/A 0.72fF
C64720 NOR2X1_LOC_315/Y INVX1_LOC_95/Y 0.27fF
C64721 INVX1_LOC_271/A INVX1_LOC_128/Y 0.13fF
C64722 NOR2X1_LOC_593/Y INVX1_LOC_37/A 0.07fF
C64723 INVX1_LOC_2/A INVX1_LOC_93/Y 0.19fF
C64724 NOR2X1_LOC_660/Y INVX1_LOC_15/A 0.04fF
C64725 INVX1_LOC_13/Y INVX1_LOC_42/A 0.06fF
C64726 NOR2X1_LOC_591/a_36_216# INVX1_LOC_76/A 0.00fF
C64727 INVX1_LOC_75/A NOR2X1_LOC_123/B 0.07fF
C64728 NOR2X1_LOC_226/A INVX1_LOC_93/Y 0.09fF
C64729 INVX1_LOC_45/Y INVX1_LOC_9/A 0.08fF
C64730 NOR2X1_LOC_541/B NOR2X1_LOC_748/A 0.03fF
C64731 INVX1_LOC_211/A INVX1_LOC_84/A 0.03fF
C64732 NOR2X1_LOC_309/Y INVX1_LOC_14/Y 0.01fF
C64733 INVX1_LOC_58/A INVX1_LOC_26/A 0.31fF
C64734 INVX1_LOC_232/Y NAND2X1_LOC_659/B 0.00fF
C64735 NOR2X1_LOC_52/B INVX1_LOC_37/A 0.07fF
C64736 INVX1_LOC_233/A NAND2X1_LOC_443/a_36_24# 0.00fF
C64737 NAND2X1_LOC_360/B INVX1_LOC_20/A 0.39fF
C64738 INVX1_LOC_14/A NOR2X1_LOC_664/a_36_216# 0.02fF
C64739 INVX1_LOC_2/A INVX1_LOC_139/A 0.03fF
C64740 INVX1_LOC_136/A NOR2X1_LOC_88/Y 0.02fF
C64741 NOR2X1_LOC_621/A NOR2X1_LOC_622/A 0.29fF
C64742 NOR2X1_LOC_624/a_36_216# NAND2X1_LOC_63/Y 0.01fF
C64743 INVX1_LOC_135/A NOR2X1_LOC_703/Y 0.03fF
C64744 INVX1_LOC_89/A NOR2X1_LOC_711/A 0.01fF
C64745 NOR2X1_LOC_500/Y NAND2X1_LOC_447/Y 0.10fF
C64746 NOR2X1_LOC_142/Y NOR2X1_LOC_142/a_36_216# 0.12fF
C64747 INVX1_LOC_2/A NAND2X1_LOC_721/A 8.73fF
C64748 INVX1_LOC_232/Y VDD 0.62fF
C64749 NOR2X1_LOC_816/A INVX1_LOC_272/A 0.09fF
C64750 INVX1_LOC_88/A INVX1_LOC_42/A 0.00fF
C64751 INVX1_LOC_35/A NOR2X1_LOC_318/A 2.82fF
C64752 INVX1_LOC_77/A NOR2X1_LOC_61/A 0.02fF
C64753 INVX1_LOC_83/Y VDD 0.41fF
C64754 NAND2X1_LOC_364/A INVX1_LOC_285/A 0.13fF
C64755 NOR2X1_LOC_433/A NOR2X1_LOC_743/Y 0.05fF
C64756 INVX1_LOC_136/A INVX1_LOC_84/A 0.17fF
C64757 NOR2X1_LOC_455/Y NOR2X1_LOC_383/B 0.00fF
C64758 INVX1_LOC_13/Y INVX1_LOC_78/A 0.03fF
C64759 NOR2X1_LOC_226/A NAND2X1_LOC_721/A 0.10fF
C64760 INVX1_LOC_197/Y VDD 0.23fF
C64761 INVX1_LOC_49/A INVX1_LOC_117/Y 0.03fF
C64762 INVX1_LOC_72/A NAND2X1_LOC_476/Y 0.03fF
C64763 NOR2X1_LOC_218/Y INVX1_LOC_139/A 0.03fF
C64764 NOR2X1_LOC_598/B NOR2X1_LOC_858/A 0.01fF
C64765 NOR2X1_LOC_554/B NOR2X1_LOC_820/B 0.01fF
C64766 NAND2X1_LOC_364/A NOR2X1_LOC_814/A 0.21fF
C64767 INPUT_0 NAND2X1_LOC_863/A 0.07fF
C64768 INVX1_LOC_269/A INVX1_LOC_32/A 0.24fF
C64769 NOR2X1_LOC_456/Y D_INPUT_1 0.05fF
C64770 NOR2X1_LOC_552/Y NOR2X1_LOC_703/A 0.02fF
C64771 NOR2X1_LOC_65/B NOR2X1_LOC_772/B 0.09fF
C64772 NAND2X1_LOC_717/Y NOR2X1_LOC_536/A 0.03fF
C64773 NOR2X1_LOC_172/a_36_216# INVX1_LOC_38/A 0.00fF
C64774 INVX1_LOC_300/A INVX1_LOC_46/A 0.02fF
C64775 INVX1_LOC_255/Y NOR2X1_LOC_138/a_36_216# 0.01fF
C64776 INVX1_LOC_305/A NOR2X1_LOC_691/B 0.02fF
C64777 INVX1_LOC_33/A NOR2X1_LOC_862/B 0.07fF
C64778 INVX1_LOC_89/A NOR2X1_LOC_552/A 0.07fF
C64779 NOR2X1_LOC_130/A NOR2X1_LOC_124/A 0.13fF
C64780 NOR2X1_LOC_446/a_36_216# INVX1_LOC_290/Y 0.01fF
C64781 NOR2X1_LOC_210/A VDD 0.00fF
C64782 D_INPUT_0 INVX1_LOC_59/Y 0.06fF
C64783 NOR2X1_LOC_65/B INVX1_LOC_13/Y 0.03fF
C64784 NOR2X1_LOC_441/Y INVX1_LOC_102/A 0.08fF
C64785 NOR2X1_LOC_52/B NOR2X1_LOC_177/Y 0.08fF
C64786 D_INPUT_0 INVX1_LOC_112/A 0.01fF
C64787 INVX1_LOC_93/Y INPUT_1 0.02fF
C64788 NAND2X1_LOC_741/B INVX1_LOC_12/A 0.02fF
C64789 NOR2X1_LOC_458/B INVX1_LOC_38/A 0.03fF
C64790 INVX1_LOC_45/A NAND2X1_LOC_291/B 0.04fF
C64791 NOR2X1_LOC_860/B NAND2X1_LOC_206/Y 0.04fF
C64792 INVX1_LOC_72/A INVX1_LOC_261/A 0.04fF
C64793 NOR2X1_LOC_598/B INVX1_LOC_292/Y 0.08fF
C64794 INVX1_LOC_161/Y INVX1_LOC_231/A 0.01fF
C64795 D_INPUT_0 INVX1_LOC_176/A 0.01fF
C64796 INVX1_LOC_88/A INVX1_LOC_78/A 0.05fF
C64797 INVX1_LOC_27/A NOR2X1_LOC_727/B 0.00fF
C64798 NOR2X1_LOC_276/Y INVX1_LOC_15/A 0.02fF
C64799 NOR2X1_LOC_6/B NOR2X1_LOC_197/B 0.13fF
C64800 INVX1_LOC_16/A NOR2X1_LOC_536/A 0.64fF
C64801 NOR2X1_LOC_356/A NOR2X1_LOC_542/B 0.02fF
C64802 NOR2X1_LOC_121/A NOR2X1_LOC_99/a_36_216# 0.00fF
C64803 NAND2X1_LOC_629/Y INVX1_LOC_179/A 0.02fF
C64804 NOR2X1_LOC_168/Y NAND2X1_LOC_74/B 0.09fF
C64805 INVX1_LOC_18/A INVX1_LOC_284/A 0.07fF
C64806 NOR2X1_LOC_361/B NOR2X1_LOC_278/Y 0.07fF
C64807 INVX1_LOC_11/A NAND2X1_LOC_72/B 1.06fF
C64808 INVX1_LOC_2/A INVX1_LOC_117/Y 0.00fF
C64809 NAND2X1_LOC_809/A VDD -0.00fF
C64810 NOR2X1_LOC_214/B NOR2X1_LOC_357/Y 0.02fF
C64811 NOR2X1_LOC_312/Y VDD 0.16fF
C64812 NOR2X1_LOC_78/B NOR2X1_LOC_433/Y 0.01fF
C64813 NAND2X1_LOC_198/B NOR2X1_LOC_89/A 1.35fF
C64814 NAND2X1_LOC_551/A NAND2X1_LOC_457/a_36_24# 0.01fF
C64815 NOR2X1_LOC_91/A INVX1_LOC_14/A 0.04fF
C64816 INVX1_LOC_30/A D_INPUT_5 0.07fF
C64817 INVX1_LOC_33/Y NAND2X1_LOC_808/A 0.06fF
C64818 NAND2X1_LOC_543/Y INVX1_LOC_54/A 0.03fF
C64819 NOR2X1_LOC_45/Y NAND2X1_LOC_454/Y 0.07fF
C64820 INVX1_LOC_235/Y NOR2X1_LOC_476/B 0.15fF
C64821 NOR2X1_LOC_65/B INVX1_LOC_88/A 0.07fF
C64822 NAND2X1_LOC_763/B D_INPUT_5 0.03fF
C64823 NOR2X1_LOC_284/B NOR2X1_LOC_445/B 0.09fF
C64824 NAND2X1_LOC_662/Y INVX1_LOC_54/A 0.10fF
C64825 NAND2X1_LOC_721/A INPUT_1 0.02fF
C64826 INVX1_LOC_136/A INVX1_LOC_15/A 0.23fF
C64827 NOR2X1_LOC_719/a_36_216# INVX1_LOC_280/A 0.00fF
C64828 INVX1_LOC_89/A NOR2X1_LOC_813/Y 0.38fF
C64829 INVX1_LOC_16/A NAND2X1_LOC_93/B 0.13fF
C64830 NOR2X1_LOC_163/Y INVX1_LOC_76/A 0.13fF
C64831 NOR2X1_LOC_328/Y INVX1_LOC_92/A 0.03fF
C64832 NAND2X1_LOC_357/B NOR2X1_LOC_662/A 0.03fF
C64833 INVX1_LOC_172/A INVX1_LOC_284/A 0.03fF
C64834 INVX1_LOC_14/A INVX1_LOC_23/A 0.05fF
C64835 NOR2X1_LOC_468/Y NAND2X1_LOC_203/a_36_24# 0.00fF
C64836 NOR2X1_LOC_84/A NAND2X1_LOC_82/Y 0.23fF
C64837 INVX1_LOC_303/A INVX1_LOC_42/A 0.07fF
C64838 INVX1_LOC_50/Y INVX1_LOC_38/Y 0.04fF
C64839 NAND2X1_LOC_464/Y NAND2X1_LOC_74/B 0.00fF
C64840 INVX1_LOC_89/A INVX1_LOC_280/A 0.36fF
C64841 NAND2X1_LOC_553/a_36_24# INVX1_LOC_123/Y 0.00fF
C64842 NOR2X1_LOC_197/a_36_216# INVX1_LOC_78/Y 0.00fF
C64843 NOR2X1_LOC_722/a_36_216# INVX1_LOC_12/A 0.00fF
C64844 INPUT_6 INVX1_LOC_1/A 0.03fF
C64845 INVX1_LOC_89/A NOR2X1_LOC_94/Y 0.03fF
C64846 NOR2X1_LOC_91/A NOR2X1_LOC_595/a_36_216# 0.14fF
C64847 INVX1_LOC_79/Y NOR2X1_LOC_334/Y 0.02fF
C64848 NAND2X1_LOC_725/A NAND2X1_LOC_493/Y 0.01fF
C64849 NAND2X1_LOC_195/Y NOR2X1_LOC_158/Y -0.00fF
C64850 INVX1_LOC_28/A NOR2X1_LOC_536/A 0.25fF
C64851 NOR2X1_LOC_785/A INVX1_LOC_57/A 0.05fF
C64852 NOR2X1_LOC_97/A VDD 0.33fF
C64853 NOR2X1_LOC_211/Y INVX1_LOC_1/A 0.01fF
C64854 NAND2X1_LOC_508/A INVX1_LOC_280/A 0.07fF
C64855 NOR2X1_LOC_570/B INVX1_LOC_290/Y 0.07fF
C64856 NAND2X1_LOC_767/a_36_24# NAND2X1_LOC_215/A 0.01fF
C64857 NAND2X1_LOC_17/a_36_24# INVX1_LOC_15/A 0.00fF
C64858 INVX1_LOC_162/Y NAND2X1_LOC_807/B 0.09fF
C64859 NAND2X1_LOC_352/B INVX1_LOC_57/A 0.15fF
C64860 INVX1_LOC_21/A NOR2X1_LOC_343/B 0.02fF
C64861 NOR2X1_LOC_34/A NOR2X1_LOC_249/Y 0.08fF
C64862 NOR2X1_LOC_644/A INVX1_LOC_9/A 0.03fF
C64863 INVX1_LOC_17/Y NOR2X1_LOC_372/A 0.16fF
C64864 NOR2X1_LOC_352/Y INVX1_LOC_19/A 0.00fF
C64865 NOR2X1_LOC_234/a_36_216# INVX1_LOC_42/A 0.01fF
C64866 INVX1_LOC_193/Y VDD 0.22fF
C64867 INVX1_LOC_16/A INVX1_LOC_3/A 0.13fF
C64868 INVX1_LOC_306/A INVX1_LOC_46/Y 0.04fF
C64869 INVX1_LOC_83/A NAND2X1_LOC_798/B 0.10fF
C64870 INVX1_LOC_147/A NOR2X1_LOC_60/Y 0.19fF
C64871 NOR2X1_LOC_391/Y VDD 0.12fF
C64872 INVX1_LOC_233/A NAND2X1_LOC_793/Y 0.02fF
C64873 INVX1_LOC_24/A INVX1_LOC_273/A 0.49fF
C64874 NAND2X1_LOC_733/Y NOR2X1_LOC_484/a_36_216# 0.00fF
C64875 INVX1_LOC_2/A NOR2X1_LOC_669/A 0.01fF
C64876 INVX1_LOC_239/A INVX1_LOC_242/A 0.10fF
C64877 NAND2X1_LOC_364/Y NOR2X1_LOC_839/B 0.18fF
C64878 INVX1_LOC_75/A NOR2X1_LOC_331/B 0.13fF
C64879 INVX1_LOC_303/A INVX1_LOC_78/A 0.07fF
C64880 NOR2X1_LOC_486/Y INVX1_LOC_247/A 0.06fF
C64881 INVX1_LOC_120/A NOR2X1_LOC_865/Y 0.03fF
C64882 NAND2X1_LOC_519/a_36_24# NAND2X1_LOC_96/A 0.00fF
C64883 INVX1_LOC_28/A NAND2X1_LOC_93/B 0.05fF
C64884 INVX1_LOC_120/A NOR2X1_LOC_243/B 0.30fF
C64885 INVX1_LOC_33/A NOR2X1_LOC_685/B 0.03fF
C64886 NOR2X1_LOC_751/A INVX1_LOC_9/A 0.01fF
C64887 NOR2X1_LOC_593/Y NAND2X1_LOC_72/B 0.07fF
C64888 INVX1_LOC_1/Y NAND2X1_LOC_63/Y 0.04fF
C64889 INVX1_LOC_34/A NOR2X1_LOC_334/Y 0.07fF
C64890 NAND2X1_LOC_35/Y INVX1_LOC_61/Y 0.02fF
C64891 INVX1_LOC_232/A INVX1_LOC_12/A 0.18fF
C64892 INVX1_LOC_256/Y INVX1_LOC_170/Y 0.04fF
C64893 NAND2X1_LOC_773/Y INVX1_LOC_299/A 1.88fF
C64894 INVX1_LOC_53/Y NOR2X1_LOC_89/A 0.42fF
C64895 NAND2X1_LOC_633/Y INVX1_LOC_304/A 0.24fF
C64896 NOR2X1_LOC_604/Y INVX1_LOC_18/A 0.02fF
C64897 NAND2X1_LOC_862/Y INVX1_LOC_84/A 0.01fF
C64898 INVX1_LOC_278/A INVX1_LOC_136/A 1.49fF
C64899 NOR2X1_LOC_45/B NOR2X1_LOC_816/Y 0.02fF
C64900 NOR2X1_LOC_65/B INVX1_LOC_303/A 0.26fF
C64901 INVX1_LOC_199/A INVX1_LOC_37/A 0.02fF
C64902 NAND2X1_LOC_860/A NOR2X1_LOC_91/Y 0.04fF
C64903 NOR2X1_LOC_13/Y INVX1_LOC_271/A 0.01fF
C64904 INVX1_LOC_22/A NOR2X1_LOC_226/Y 0.01fF
C64905 NOR2X1_LOC_569/Y INVX1_LOC_99/A 0.07fF
C64906 NAND2X1_LOC_725/Y NAND2X1_LOC_863/Y 0.71fF
C64907 INVX1_LOC_35/A INVX1_LOC_305/A 0.04fF
C64908 INVX1_LOC_126/A NAND2X1_LOC_650/B 0.27fF
C64909 NOR2X1_LOC_225/a_36_216# NAND2X1_LOC_474/Y 0.00fF
C64910 NOR2X1_LOC_383/Y INVX1_LOC_12/A 0.06fF
C64911 NAND2X1_LOC_624/B NOR2X1_LOC_384/Y 0.02fF
C64912 D_INPUT_1 NOR2X1_LOC_759/Y 0.03fF
C64913 NAND2X1_LOC_360/B INVX1_LOC_4/A 1.27fF
C64914 NOR2X1_LOC_665/A NOR2X1_LOC_89/A 0.02fF
C64915 NOR2X1_LOC_272/Y NOR2X1_LOC_590/A 0.01fF
C64916 NAND2X1_LOC_363/B NOR2X1_LOC_360/Y 0.07fF
C64917 INVX1_LOC_202/A D_INPUT_1 0.75fF
C64918 NAND2X1_LOC_563/A INVX1_LOC_32/A 0.02fF
C64919 GATE_811 NOR2X1_LOC_829/A 0.25fF
C64920 NAND2X1_LOC_860/A NOR2X1_LOC_81/a_36_216# 0.01fF
C64921 INVX1_LOC_28/A INVX1_LOC_3/A 0.25fF
C64922 NAND2X1_LOC_218/B NAND2X1_LOC_38/a_36_24# 0.00fF
C64923 INVX1_LOC_255/Y NOR2X1_LOC_861/Y 0.03fF
C64924 INVX1_LOC_239/A NOR2X1_LOC_573/Y 0.03fF
C64925 INVX1_LOC_2/A INVX1_LOC_87/A 0.01fF
C64926 NOR2X1_LOC_318/B INVX1_LOC_118/A 0.04fF
C64927 VDD NAND2X1_LOC_287/B 0.01fF
C64928 NAND2X1_LOC_370/a_36_24# INVX1_LOC_41/Y 0.00fF
C64929 NOR2X1_LOC_658/Y INVX1_LOC_27/A 0.07fF
C64930 INVX1_LOC_13/A NOR2X1_LOC_554/A 0.03fF
C64931 VDD NOR2X1_LOC_858/B 0.31fF
C64932 NAND2X1_LOC_175/B INVX1_LOC_271/A 0.03fF
C64933 NAND2X1_LOC_571/a_36_24# NAND2X1_LOC_571/Y 0.01fF
C64934 NAND2X1_LOC_72/Y INVX1_LOC_94/A 0.27fF
C64935 NOR2X1_LOC_226/A INVX1_LOC_87/A 0.03fF
C64936 INVX1_LOC_269/A INPUT_3 0.01fF
C64937 NOR2X1_LOC_186/Y NOR2X1_LOC_68/A 0.07fF
C64938 NAND2X1_LOC_126/a_36_24# INVX1_LOC_3/A 0.00fF
C64939 VDD INVX1_LOC_129/Y 0.46fF
C64940 NOR2X1_LOC_536/A NOR2X1_LOC_35/Y 0.01fF
C64941 NOR2X1_LOC_598/B NAND2X1_LOC_361/Y 0.10fF
C64942 INVX1_LOC_217/Y INVX1_LOC_23/A 0.04fF
C64943 INVX1_LOC_14/A INVX1_LOC_31/A 0.17fF
C64944 INVX1_LOC_1/A NOR2X1_LOC_514/A 0.68fF
C64945 NOR2X1_LOC_161/a_36_216# NAND2X1_LOC_425/Y 0.01fF
C64946 NOR2X1_LOC_275/a_36_216# INVX1_LOC_103/A 0.00fF
C64947 INVX1_LOC_186/A INVX1_LOC_307/A 0.07fF
C64948 NAND2X1_LOC_337/B INVX1_LOC_150/Y 0.01fF
C64949 INVX1_LOC_17/A NOR2X1_LOC_389/A 0.10fF
C64950 NAND2X1_LOC_655/A INVX1_LOC_291/A 0.23fF
C64951 NAND2X1_LOC_357/B INVX1_LOC_57/A 0.21fF
C64952 INVX1_LOC_35/A NAND2X1_LOC_536/a_36_24# 0.00fF
C64953 INVX1_LOC_96/A NOR2X1_LOC_197/B 0.01fF
C64954 INVX1_LOC_104/A INVX1_LOC_29/Y 0.09fF
C64955 INVX1_LOC_36/A NAND2X1_LOC_303/Y 3.09fF
C64956 NAND2X1_LOC_338/B NOR2X1_LOC_843/B 0.07fF
C64957 NAND2X1_LOC_778/Y INVX1_LOC_24/A 0.28fF
C64958 INVX1_LOC_186/A NOR2X1_LOC_445/B 0.07fF
C64959 NAND2X1_LOC_573/Y NOR2X1_LOC_68/A 0.07fF
C64960 INVX1_LOC_1/A INVX1_LOC_142/A 0.09fF
C64961 NOR2X1_LOC_331/B NAND2X1_LOC_453/A 0.12fF
C64962 INVX1_LOC_304/A INVX1_LOC_71/Y 0.32fF
C64963 INVX1_LOC_91/A NOR2X1_LOC_841/A 2.15fF
C64964 INVX1_LOC_58/A INVX1_LOC_149/A 0.01fF
C64965 NOR2X1_LOC_480/A INVX1_LOC_163/A 0.04fF
C64966 NAND2X1_LOC_149/Y NOR2X1_LOC_781/Y 0.00fF
C64967 NAND2X1_LOC_30/Y NAND2X1_LOC_36/A 1.73fF
C64968 NOR2X1_LOC_68/A NAND2X1_LOC_724/A 0.37fF
C64969 INVX1_LOC_111/Y INVX1_LOC_23/A 0.02fF
C64970 NOR2X1_LOC_490/Y NOR2X1_LOC_490/a_36_216# 0.01fF
C64971 NAND2X1_LOC_724/Y NOR2X1_LOC_505/Y 0.03fF
C64972 NAND2X1_LOC_447/Y INVX1_LOC_307/A 0.00fF
C64973 INVX1_LOC_206/A NOR2X1_LOC_717/A 0.10fF
C64974 INVX1_LOC_50/A NOR2X1_LOC_136/Y 0.28fF
C64975 INVX1_LOC_123/A INVX1_LOC_293/Y -0.04fF
C64976 NOR2X1_LOC_482/Y NOR2X1_LOC_754/Y 0.04fF
C64977 NOR2X1_LOC_15/Y INVX1_LOC_24/A 0.16fF
C64978 NAND2X1_LOC_721/A INVX1_LOC_118/A 0.07fF
C64979 NOR2X1_LOC_541/Y NOR2X1_LOC_274/B 0.04fF
C64980 NOR2X1_LOC_405/A INVX1_LOC_285/A 0.01fF
C64981 NAND2X1_LOC_573/A NOR2X1_LOC_278/Y 1.04fF
C64982 INVX1_LOC_179/A INVX1_LOC_76/A 0.03fF
C64983 NOR2X1_LOC_349/A NOR2X1_LOC_814/A 0.12fF
C64984 INVX1_LOC_17/A INVX1_LOC_62/Y 0.02fF
C64985 NOR2X1_LOC_643/Y NAND2X1_LOC_218/A 0.05fF
C64986 NOR2X1_LOC_590/A NOR2X1_LOC_336/B 0.16fF
C64987 NOR2X1_LOC_113/A NOR2X1_LOC_814/A 0.00fF
C64988 INVX1_LOC_11/A NAND2X1_LOC_198/B 0.01fF
C64989 INVX1_LOC_36/A NAND2X1_LOC_120/a_36_24# 0.00fF
C64990 NOR2X1_LOC_405/A NOR2X1_LOC_814/A 0.34fF
C64991 VDD NOR2X1_LOC_809/B 0.06fF
C64992 NAND2X1_LOC_733/Y NAND2X1_LOC_741/B 2.53fF
C64993 NOR2X1_LOC_792/B NOR2X1_LOC_791/Y 0.17fF
C64994 NOR2X1_LOC_441/Y INVX1_LOC_223/A 0.10fF
C64995 INVX1_LOC_88/A NOR2X1_LOC_152/Y 0.03fF
C64996 NOR2X1_LOC_592/B NAND2X1_LOC_453/A 0.06fF
C64997 INVX1_LOC_125/Y INVX1_LOC_125/A 0.10fF
C64998 INVX1_LOC_123/A NAND2X1_LOC_74/B 0.74fF
C64999 INVX1_LOC_20/A NAND2X1_LOC_572/B 0.71fF
C65000 NOR2X1_LOC_844/Y NOR2X1_LOC_500/B 0.15fF
C65001 NOR2X1_LOC_590/A NAND2X1_LOC_364/A 3.50fF
C65002 NOR2X1_LOC_328/Y INVX1_LOC_53/A 0.03fF
C65003 NOR2X1_LOC_15/Y NOR2X1_LOC_557/Y 0.36fF
C65004 NOR2X1_LOC_329/B NOR2X1_LOC_681/a_36_216# 0.01fF
C65005 INVX1_LOC_89/A NOR2X1_LOC_541/B 0.01fF
C65006 NAND2X1_LOC_551/A NOR2X1_LOC_89/Y 0.00fF
C65007 NAND2X1_LOC_549/Y INVX1_LOC_316/Y 0.01fF
C65008 INVX1_LOC_33/Y INVX1_LOC_92/A 0.03fF
C65009 NOR2X1_LOC_471/Y NOR2X1_LOC_596/A 0.07fF
C65010 NOR2X1_LOC_656/a_36_216# INVX1_LOC_31/A 0.01fF
C65011 INVX1_LOC_244/A INVX1_LOC_78/A 0.03fF
C65012 INVX1_LOC_45/A NOR2X1_LOC_274/B 0.02fF
C65013 NAND2X1_LOC_714/B NOR2X1_LOC_591/Y 2.48fF
C65014 INVX1_LOC_89/A NAND2X1_LOC_416/a_36_24# 0.00fF
C65015 NOR2X1_LOC_568/A NOR2X1_LOC_274/B 0.03fF
C65016 NAND2X1_LOC_725/Y NOR2X1_LOC_700/a_36_216# 0.16fF
C65017 INVX1_LOC_93/Y NAND2X1_LOC_63/Y 0.01fF
C65018 INVX1_LOC_134/A INVX1_LOC_49/A 0.06fF
C65019 NOR2X1_LOC_857/A NOR2X1_LOC_814/A 0.07fF
C65020 INVX1_LOC_30/A NOR2X1_LOC_360/Y 0.23fF
C65021 NOR2X1_LOC_335/B NAND2X1_LOC_647/B 0.11fF
C65022 INVX1_LOC_72/A INVX1_LOC_18/A 1.27fF
C65023 INVX1_LOC_20/A NAND2X1_LOC_219/B 0.00fF
C65024 D_INPUT_3 INVX1_LOC_63/A 0.03fF
C65025 INVX1_LOC_17/A NOR2X1_LOC_295/Y 0.01fF
C65026 NOR2X1_LOC_121/a_36_216# INVX1_LOC_306/Y 0.01fF
C65027 NOR2X1_LOC_137/A INVX1_LOC_23/A 0.07fF
C65028 NAND2X1_LOC_728/Y INVX1_LOC_72/A 0.10fF
C65029 INVX1_LOC_24/Y NOR2X1_LOC_802/A 0.05fF
C65030 INPUT_0 NAND2X1_LOC_444/B 0.03fF
C65031 INVX1_LOC_56/Y INVX1_LOC_306/Y 0.13fF
C65032 INPUT_0 NOR2X1_LOC_334/Y 0.14fF
C65033 NAND2X1_LOC_16/a_36_24# NOR2X1_LOC_596/A 0.00fF
C65034 NOR2X1_LOC_75/Y NOR2X1_LOC_433/a_36_216# 0.00fF
C65035 INVX1_LOC_17/A NOR2X1_LOC_844/A 0.01fF
C65036 NOR2X1_LOC_742/A NOR2X1_LOC_631/Y 0.01fF
C65037 INVX1_LOC_249/A NOR2X1_LOC_658/Y 0.04fF
C65038 INVX1_LOC_135/A NOR2X1_LOC_392/Y 2.01fF
C65039 NAND2X1_LOC_711/B INVX1_LOC_72/A 0.15fF
C65040 NOR2X1_LOC_15/Y INVX1_LOC_143/A 0.07fF
C65041 INVX1_LOC_36/A NOR2X1_LOC_106/Y 0.19fF
C65042 NOR2X1_LOC_637/Y INVX1_LOC_72/A 0.01fF
C65043 NAND2X1_LOC_36/A INVX1_LOC_49/A 0.02fF
C65044 INVX1_LOC_171/A INVX1_LOC_58/Y 0.01fF
C65045 INVX1_LOC_289/Y NOR2X1_LOC_226/A 0.14fF
C65046 NAND2X1_LOC_236/a_36_24# INVX1_LOC_3/A 0.00fF
C65047 NOR2X1_LOC_617/Y NOR2X1_LOC_384/Y 0.02fF
C65048 INVX1_LOC_45/A NOR2X1_LOC_577/Y 0.09fF
C65049 INVX1_LOC_278/A NAND2X1_LOC_862/Y 0.01fF
C65050 INVX1_LOC_30/A NAND2X1_LOC_652/a_36_24# 0.00fF
C65051 INVX1_LOC_21/A NAND2X1_LOC_41/Y 0.00fF
C65052 INVX1_LOC_17/Y NAND2X1_LOC_560/A 0.00fF
C65053 INVX1_LOC_2/A NOR2X1_LOC_82/A 0.18fF
C65054 NOR2X1_LOC_778/Y INVX1_LOC_33/A 0.07fF
C65055 INVX1_LOC_230/A INVX1_LOC_63/A 0.46fF
C65056 NAND2X1_LOC_84/Y INVX1_LOC_111/A 0.03fF
C65057 INVX1_LOC_132/A NOR2X1_LOC_68/A 0.07fF
C65058 NOR2X1_LOC_690/A INVX1_LOC_36/A 2.32fF
C65059 NOR2X1_LOC_226/A NOR2X1_LOC_82/A 0.09fF
C65060 INVX1_LOC_223/A NOR2X1_LOC_142/Y 0.01fF
C65061 NOR2X1_LOC_52/Y INVX1_LOC_33/A 0.19fF
C65062 NOR2X1_LOC_188/A NOR2X1_LOC_720/A 0.03fF
C65063 NAND2X1_LOC_198/B NOR2X1_LOC_433/A 0.10fF
C65064 INVX1_LOC_50/A INVX1_LOC_144/A 0.01fF
C65065 NAND2X1_LOC_725/Y INVX1_LOC_282/A 0.05fF
C65066 INVX1_LOC_75/A NOR2X1_LOC_493/A 0.02fF
C65067 NOR2X1_LOC_160/B INVX1_LOC_210/A 0.05fF
C65068 INVX1_LOC_203/Y NOR2X1_LOC_480/A 0.01fF
C65069 INVX1_LOC_37/A NAND2X1_LOC_254/Y 0.00fF
C65070 NOR2X1_LOC_270/Y INVX1_LOC_33/A 0.01fF
C65071 INVX1_LOC_41/A NOR2X1_LOC_791/B 0.01fF
C65072 NAND2X1_LOC_474/a_36_24# NAND2X1_LOC_474/Y 0.02fF
C65073 INVX1_LOC_235/A INVX1_LOC_135/A 0.06fF
C65074 NAND2X1_LOC_30/Y NAND2X1_LOC_59/a_36_24# 0.00fF
C65075 NOR2X1_LOC_653/B NOR2X1_LOC_246/A 0.03fF
C65076 NOR2X1_LOC_176/Y INVX1_LOC_102/A 0.03fF
C65077 INVX1_LOC_224/Y INVX1_LOC_100/A 0.09fF
C65078 INVX1_LOC_58/A NOR2X1_LOC_368/A 0.08fF
C65079 NOR2X1_LOC_324/A NOR2X1_LOC_334/Y 0.13fF
C65080 INVX1_LOC_11/A INVX1_LOC_53/Y 0.04fF
C65081 NOR2X1_LOC_577/Y INVX1_LOC_71/A 0.07fF
C65082 NOR2X1_LOC_195/A NOR2X1_LOC_516/B 0.00fF
C65083 INPUT_3 NAND2X1_LOC_563/A 0.07fF
C65084 INVX1_LOC_225/A NOR2X1_LOC_68/A 0.02fF
C65085 INVX1_LOC_103/A NAND2X1_LOC_660/Y 0.07fF
C65086 INVX1_LOC_256/A INVX1_LOC_16/A 0.10fF
C65087 NOR2X1_LOC_541/Y INVX1_LOC_22/A 0.03fF
C65088 NAND2X1_LOC_393/a_36_24# INVX1_LOC_135/A 0.01fF
C65089 INVX1_LOC_34/A NAND2X1_LOC_758/a_36_24# 0.00fF
C65090 INVX1_LOC_284/Y INVX1_LOC_280/Y 0.14fF
C65091 INVX1_LOC_47/Y INVX1_LOC_46/A 0.29fF
C65092 INVX1_LOC_279/Y NOR2X1_LOC_544/A 0.19fF
C65093 INVX1_LOC_30/A NAND2X1_LOC_451/Y 0.19fF
C65094 NOR2X1_LOC_15/Y NOR2X1_LOC_130/A 0.03fF
C65095 INVX1_LOC_222/A INVX1_LOC_58/Y 0.38fF
C65096 NOR2X1_LOC_655/B INVX1_LOC_223/A 0.10fF
C65097 NOR2X1_LOC_75/Y NOR2X1_LOC_589/A 0.07fF
C65098 INVX1_LOC_72/A INVX1_LOC_34/Y 0.01fF
C65099 NAND2X1_LOC_198/B NOR2X1_LOC_52/B 0.03fF
C65100 INVX1_LOC_12/Y INVX1_LOC_32/A 0.01fF
C65101 INVX1_LOC_11/A NOR2X1_LOC_781/B 0.07fF
C65102 NOR2X1_LOC_391/B NOR2X1_LOC_392/Y 0.09fF
C65103 INVX1_LOC_223/Y NAND2X1_LOC_184/a_36_24# 0.00fF
C65104 NAND2X1_LOC_763/B NAND2X1_LOC_451/Y 0.14fF
C65105 INVX1_LOC_283/Y NOR2X1_LOC_718/Y 0.21fF
C65106 NAND2X1_LOC_789/a_36_24# NOR2X1_LOC_175/A 0.00fF
C65107 INVX1_LOC_13/A NOR2X1_LOC_160/B 0.37fF
C65108 INVX1_LOC_235/Y INVX1_LOC_169/A 0.01fF
C65109 NOR2X1_LOC_68/A NOR2X1_LOC_209/Y 0.07fF
C65110 INVX1_LOC_95/Y NAND2X1_LOC_99/A 0.19fF
C65111 NOR2X1_LOC_348/B INVX1_LOC_71/A 0.01fF
C65112 INVX1_LOC_34/A INVX1_LOC_209/Y 0.03fF
C65113 INVX1_LOC_45/A INVX1_LOC_22/A 0.10fF
C65114 INVX1_LOC_290/Y INVX1_LOC_54/A 0.03fF
C65115 NOR2X1_LOC_230/Y INVX1_LOC_290/A 0.06fF
C65116 NOR2X1_LOC_568/A INVX1_LOC_22/A 1.50fF
C65117 NOR2X1_LOC_449/A NAND2X1_LOC_453/A 0.03fF
C65118 NOR2X1_LOC_188/A NOR2X1_LOC_849/A 0.03fF
C65119 NAND2X1_LOC_856/A INVX1_LOC_22/A 0.03fF
C65120 NAND2X1_LOC_288/B INVX1_LOC_76/A 0.10fF
C65121 INVX1_LOC_247/A NOR2X1_LOC_748/A 0.03fF
C65122 NOR2X1_LOC_99/Y INVX1_LOC_42/A 0.19fF
C65123 NOR2X1_LOC_364/A INVX1_LOC_109/Y 0.01fF
C65124 NAND2X1_LOC_493/Y NAND2X1_LOC_560/A 0.03fF
C65125 NOR2X1_LOC_82/A INPUT_1 0.32fF
C65126 NAND2X1_LOC_456/Y NAND2X1_LOC_773/B 0.01fF
C65127 INVX1_LOC_20/A NOR2X1_LOC_654/A 0.01fF
C65128 NOR2X1_LOC_638/a_36_216# INVX1_LOC_191/Y -0.00fF
C65129 NAND2X1_LOC_551/A NAND2X1_LOC_550/A 0.02fF
C65130 NOR2X1_LOC_142/Y INVX1_LOC_85/A 0.02fF
C65131 NOR2X1_LOC_787/a_36_216# INVX1_LOC_313/Y 0.00fF
C65132 INVX1_LOC_24/A NAND2X1_LOC_840/B 0.01fF
C65133 NOR2X1_LOC_160/B NOR2X1_LOC_174/B 0.05fF
C65134 INVX1_LOC_41/A NOR2X1_LOC_802/A 0.07fF
C65135 NOR2X1_LOC_4/a_36_216# NOR2X1_LOC_6/B 0.03fF
C65136 NOR2X1_LOC_690/Y INVX1_LOC_72/A 0.03fF
C65137 VDD NOR2X1_LOC_72/Y 0.12fF
C65138 INVX1_LOC_33/A NOR2X1_LOC_172/a_36_216# 0.00fF
C65139 INVX1_LOC_256/A INVX1_LOC_28/A 1.37fF
C65140 NOR2X1_LOC_8/a_36_216# INVX1_LOC_316/Y 0.01fF
C65141 NOR2X1_LOC_284/a_36_216# INVX1_LOC_77/A 0.00fF
C65142 NOR2X1_LOC_308/a_36_216# INVX1_LOC_117/A 0.00fF
C65143 INVX1_LOC_2/A NAND2X1_LOC_332/Y 0.06fF
C65144 NOR2X1_LOC_831/Y INVX1_LOC_63/A 0.08fF
C65145 INVX1_LOC_71/A INVX1_LOC_22/A 0.26fF
C65146 NAND2X1_LOC_425/Y NOR2X1_LOC_460/a_36_216# 0.01fF
C65147 NOR2X1_LOC_219/Y NOR2X1_LOC_433/A 0.04fF
C65148 INVX1_LOC_98/A NAND2X1_LOC_474/Y -0.04fF
C65149 NOR2X1_LOC_433/A INVX1_LOC_53/Y 0.07fF
C65150 INVX1_LOC_45/Y NOR2X1_LOC_561/Y 0.01fF
C65151 NAND2X1_LOC_387/B INVX1_LOC_89/A 0.01fF
C65152 NOR2X1_LOC_355/A INVX1_LOC_177/Y 0.15fF
C65153 NAND2X1_LOC_80/a_36_24# NAND2X1_LOC_773/B 0.00fF
C65154 INVX1_LOC_34/A NOR2X1_LOC_44/a_36_216# 0.00fF
C65155 NOR2X1_LOC_100/a_36_216# NOR2X1_LOC_849/A 0.00fF
C65156 NOR2X1_LOC_78/A NAND2X1_LOC_474/Y 0.07fF
C65157 INVX1_LOC_223/Y NOR2X1_LOC_552/A 0.00fF
C65158 INVX1_LOC_14/A INVX1_LOC_6/A 1.28fF
C65159 NAND2X1_LOC_180/a_36_24# NOR2X1_LOC_226/A 0.00fF
C65160 NOR2X1_LOC_103/Y INVX1_LOC_100/A 0.03fF
C65161 INVX1_LOC_90/A NOR2X1_LOC_703/B 0.05fF
C65162 NAND2X1_LOC_447/a_36_24# INVX1_LOC_92/A 0.00fF
C65163 NOR2X1_LOC_39/Y INVX1_LOC_9/A 0.07fF
C65164 NAND2X1_LOC_223/a_36_24# NOR2X1_LOC_814/A 0.01fF
C65165 NAND2X1_LOC_572/B INVX1_LOC_4/A 0.18fF
C65166 INVX1_LOC_18/A INVX1_LOC_313/Y 0.03fF
C65167 INVX1_LOC_33/Y INVX1_LOC_53/A 0.05fF
C65168 NOR2X1_LOC_241/A NOR2X1_LOC_334/A 0.28fF
C65169 NAND2X1_LOC_338/B INVX1_LOC_34/Y 0.27fF
C65170 INVX1_LOC_145/Y NOR2X1_LOC_433/A 0.03fF
C65171 INVX1_LOC_30/A NOR2X1_LOC_567/B 0.19fF
C65172 NOR2X1_LOC_219/Y NOR2X1_LOC_52/B 0.19fF
C65173 NOR2X1_LOC_778/B NOR2X1_LOC_724/a_36_216# 0.00fF
C65174 INVX1_LOC_217/Y NAND2X1_LOC_859/Y 0.01fF
C65175 INVX1_LOC_78/A INVX1_LOC_107/Y 0.02fF
C65176 INVX1_LOC_17/A NAND2X1_LOC_498/a_36_24# 0.00fF
C65177 NOR2X1_LOC_52/B INVX1_LOC_53/Y 0.04fF
C65178 NOR2X1_LOC_488/Y NAND2X1_LOC_785/A 0.01fF
C65179 NAND2X1_LOC_647/B INVX1_LOC_84/A 0.02fF
C65180 NAND2X1_LOC_727/Y INVX1_LOC_240/A 0.12fF
C65181 VDD INVX1_LOC_50/Y 1.92fF
C65182 NOR2X1_LOC_392/Y INVX1_LOC_280/A 0.16fF
C65183 INVX1_LOC_104/A INVX1_LOC_101/A 0.02fF
C65184 NOR2X1_LOC_94/Y NOR2X1_LOC_392/Y 0.02fF
C65185 NAND2X1_LOC_308/B NOR2X1_LOC_152/Y 0.01fF
C65186 INVX1_LOC_158/Y NOR2X1_LOC_500/B 0.10fF
C65187 NOR2X1_LOC_705/B INVX1_LOC_91/A 0.00fF
C65188 NOR2X1_LOC_717/Y INVX1_LOC_6/A 0.31fF
C65189 INVX1_LOC_50/A NOR2X1_LOC_155/A 0.10fF
C65190 INVX1_LOC_145/Y NOR2X1_LOC_52/B 0.01fF
C65191 INVX1_LOC_58/A NOR2X1_LOC_235/Y 0.01fF
C65192 NOR2X1_LOC_208/Y NOR2X1_LOC_736/a_36_216# 0.01fF
C65193 NOR2X1_LOC_589/A INVX1_LOC_98/Y 0.01fF
C65194 NOR2X1_LOC_566/Y INVX1_LOC_232/A 0.04fF
C65195 NOR2X1_LOC_355/A INVX1_LOC_104/A 0.01fF
C65196 INVX1_LOC_17/A NAND2X1_LOC_655/B 0.01fF
C65197 NOR2X1_LOC_523/B INPUT_0 0.01fF
C65198 INVX1_LOC_266/A VDD 1.18fF
C65199 NOR2X1_LOC_495/Y NAND2X1_LOC_560/A 0.00fF
C65200 NOR2X1_LOC_590/A NOR2X1_LOC_113/A 0.01fF
C65201 NOR2X1_LOC_381/Y VDD 0.63fF
C65202 NOR2X1_LOC_590/A NOR2X1_LOC_405/A 0.08fF
C65203 INVX1_LOC_136/A INVX1_LOC_123/A 0.10fF
C65204 INVX1_LOC_271/A NOR2X1_LOC_697/Y 0.02fF
C65205 INVX1_LOC_256/A NOR2X1_LOC_35/Y 0.10fF
C65206 INVX1_LOC_78/A INVX1_LOC_272/A 0.07fF
C65207 INVX1_LOC_11/A NOR2X1_LOC_585/Y 0.03fF
C65208 NAND2X1_LOC_63/Y INVX1_LOC_87/A 0.03fF
C65209 INVX1_LOC_30/A NOR2X1_LOC_269/Y 0.01fF
C65210 NAND2X1_LOC_660/a_36_24# NAND2X1_LOC_660/A 0.00fF
C65211 INVX1_LOC_282/A NOR2X1_LOC_625/Y 0.01fF
C65212 INVX1_LOC_13/A NOR2X1_LOC_516/B 0.36fF
C65213 NAND2X1_LOC_11/Y NOR2X1_LOC_763/Y 0.64fF
C65214 NAND2X1_LOC_81/B NOR2X1_LOC_278/Y 0.03fF
C65215 NOR2X1_LOC_15/Y NAND2X1_LOC_811/B 0.06fF
C65216 INVX1_LOC_48/Y NOR2X1_LOC_536/A 0.03fF
C65217 NOR2X1_LOC_322/Y NAND2X1_LOC_833/Y 0.01fF
C65218 INVX1_LOC_24/A NOR2X1_LOC_733/Y 0.01fF
C65219 NOR2X1_LOC_479/B NOR2X1_LOC_459/A 0.03fF
C65220 INVX1_LOC_23/A NOR2X1_LOC_127/Y 0.17fF
C65221 NAND2X1_LOC_545/a_36_24# NOR2X1_LOC_78/A 0.01fF
C65222 NAND2X1_LOC_783/Y INVX1_LOC_20/A 0.01fF
C65223 NOR2X1_LOC_440/Y INVX1_LOC_16/A 0.16fF
C65224 INVX1_LOC_26/Y INVX1_LOC_125/A 0.07fF
C65225 INVX1_LOC_201/Y INVX1_LOC_82/Y 0.05fF
C65226 INVX1_LOC_35/A NAND2X1_LOC_438/a_36_24# 0.01fF
C65227 NOR2X1_LOC_160/B NOR2X1_LOC_357/Y 0.07fF
C65228 NOR2X1_LOC_388/Y INVX1_LOC_75/A 0.15fF
C65229 NOR2X1_LOC_537/A INVX1_LOC_222/A 0.03fF
C65230 NAND2X1_LOC_555/Y NAND2X1_LOC_414/a_36_24# 0.00fF
C65231 INVX1_LOC_255/Y INVX1_LOC_7/A 0.14fF
C65232 NOR2X1_LOC_303/Y INVX1_LOC_78/Y 0.00fF
C65233 NOR2X1_LOC_590/A NOR2X1_LOC_857/A 0.08fF
C65234 NOR2X1_LOC_101/a_36_216# INVX1_LOC_306/Y 0.01fF
C65235 D_INPUT_1 INVX1_LOC_293/Y 0.02fF
C65236 INVX1_LOC_77/A INVX1_LOC_286/A 0.07fF
C65237 INVX1_LOC_135/A INVX1_LOC_25/Y 0.01fF
C65238 NOR2X1_LOC_413/Y NOR2X1_LOC_19/Y 0.04fF
C65239 NOR2X1_LOC_68/A NAND2X1_LOC_642/Y 0.19fF
C65240 NOR2X1_LOC_454/Y INVX1_LOC_54/A 0.16fF
C65241 NOR2X1_LOC_424/Y NOR2X1_LOC_589/A 0.11fF
C65242 NOR2X1_LOC_644/A INVX1_LOC_179/Y 0.03fF
C65243 INVX1_LOC_33/A NOR2X1_LOC_500/a_36_216# 0.00fF
C65244 NOR2X1_LOC_123/B INVX1_LOC_22/A 0.11fF
C65245 INVX1_LOC_289/Y INVX1_LOC_118/A 0.05fF
C65246 NOR2X1_LOC_516/B NOR2X1_LOC_174/B 0.03fF
C65247 NOR2X1_LOC_209/Y NOR2X1_LOC_590/a_36_216# 0.00fF
C65248 NOR2X1_LOC_627/a_36_216# NOR2X1_LOC_742/A 0.01fF
C65249 NAND2X1_LOC_265/a_36_24# INVX1_LOC_125/A 0.02fF
C65250 INVX1_LOC_221/Y INVX1_LOC_38/A 0.05fF
C65251 NAND2X1_LOC_550/A NOR2X1_LOC_692/Y 0.00fF
C65252 NOR2X1_LOC_248/Y VDD 0.26fF
C65253 INVX1_LOC_5/A NOR2X1_LOC_673/A 0.03fF
C65254 NOR2X1_LOC_286/Y NOR2X1_LOC_729/A 0.01fF
C65255 D_INPUT_1 NAND2X1_LOC_74/B 0.08fF
C65256 NOR2X1_LOC_113/B NOR2X1_LOC_52/B 0.02fF
C65257 NOR2X1_LOC_254/Y INVX1_LOC_78/Y 0.04fF
C65258 INVX1_LOC_27/A NAND2X1_LOC_85/Y 0.03fF
C65259 NOR2X1_LOC_592/a_36_216# NOR2X1_LOC_331/B 0.02fF
C65260 INVX1_LOC_50/A NOR2X1_LOC_833/B 0.01fF
C65261 NOR2X1_LOC_552/Y INVX1_LOC_104/A 0.02fF
C65262 INVX1_LOC_14/A NOR2X1_LOC_79/A 0.01fF
C65263 NOR2X1_LOC_82/A INVX1_LOC_118/A 0.46fF
C65264 NOR2X1_LOC_172/Y INVX1_LOC_91/A 0.05fF
C65265 NOR2X1_LOC_268/a_36_216# INVX1_LOC_76/A -0.01fF
C65266 NAND2X1_LOC_725/A INVX1_LOC_240/Y 0.03fF
C65267 D_INPUT_1 NOR2X1_LOC_847/B 0.70fF
C65268 NOR2X1_LOC_795/Y NOR2X1_LOC_703/Y 0.02fF
C65269 INVX1_LOC_41/A NOR2X1_LOC_192/A 0.02fF
C65270 NOR2X1_LOC_662/A NOR2X1_LOC_291/Y 0.01fF
C65271 NAND2X1_LOC_140/a_36_24# NAND2X1_LOC_468/B 0.00fF
C65272 INVX1_LOC_124/A INVX1_LOC_286/A 0.03fF
C65273 NAND2X1_LOC_618/Y INVX1_LOC_175/A 0.00fF
C65274 NAND2X1_LOC_356/a_36_24# INVX1_LOC_146/Y 0.01fF
C65275 INVX1_LOC_181/Y NOR2X1_LOC_558/A 0.00fF
C65276 NOR2X1_LOC_392/B INVX1_LOC_91/A 0.07fF
C65277 INVX1_LOC_90/Y NOR2X1_LOC_415/Y 0.01fF
C65278 NOR2X1_LOC_636/B INVX1_LOC_92/A 0.08fF
C65279 NOR2X1_LOC_86/Y NOR2X1_LOC_813/Y 0.03fF
C65280 NOR2X1_LOC_353/Y INVX1_LOC_78/Y 0.01fF
C65281 INVX1_LOC_125/Y NOR2X1_LOC_709/A 0.02fF
C65282 INVX1_LOC_48/Y INVX1_LOC_3/A 0.03fF
C65283 NAND2X1_LOC_500/Y INVX1_LOC_118/A 0.01fF
C65284 INVX1_LOC_49/A INVX1_LOC_176/A 0.03fF
C65285 INVX1_LOC_314/Y INVX1_LOC_37/A 1.79fF
C65286 NOR2X1_LOC_716/B INVX1_LOC_20/A 0.17fF
C65287 NOR2X1_LOC_742/A NOR2X1_LOC_302/a_36_216# 0.01fF
C65288 NOR2X1_LOC_703/B INVX1_LOC_38/A 0.03fF
C65289 NOR2X1_LOC_592/a_36_216# NOR2X1_LOC_592/B 0.00fF
C65290 INVX1_LOC_314/Y NOR2X1_LOC_231/A 0.01fF
C65291 INVX1_LOC_30/Y NOR2X1_LOC_721/Y 0.02fF
C65292 NOR2X1_LOC_160/B NOR2X1_LOC_259/B 0.05fF
C65293 INVX1_LOC_69/Y INVX1_LOC_16/A 0.03fF
C65294 NOR2X1_LOC_112/B NOR2X1_LOC_97/B 0.00fF
C65295 NOR2X1_LOC_52/Y NOR2X1_LOC_351/Y 0.00fF
C65296 INVX1_LOC_58/Y INVX1_LOC_4/A 0.85fF
C65297 NOR2X1_LOC_374/a_36_216# NOR2X1_LOC_78/A 0.00fF
C65298 INVX1_LOC_135/A INVX1_LOC_75/A 0.90fF
C65299 NOR2X1_LOC_91/A NOR2X1_LOC_689/A 0.06fF
C65300 INVX1_LOC_143/A NAND2X1_LOC_108/a_36_24# 0.00fF
C65301 INVX1_LOC_30/A NOR2X1_LOC_79/Y 0.09fF
C65302 NAND2X1_LOC_149/Y NOR2X1_LOC_89/A 0.08fF
C65303 INVX1_LOC_226/Y NOR2X1_LOC_78/A 0.07fF
C65304 INVX1_LOC_232/Y INVX1_LOC_316/A 0.01fF
C65305 INVX1_LOC_295/A INVX1_LOC_75/A 0.17fF
C65306 NOR2X1_LOC_818/Y INVX1_LOC_59/Y 0.00fF
C65307 NOR2X1_LOC_6/B VDD 3.49fF
C65308 NOR2X1_LOC_181/Y INVX1_LOC_37/A 0.26fF
C65309 NAND2X1_LOC_550/A NAND2X1_LOC_489/Y 0.01fF
C65310 NOR2X1_LOC_282/Y INVX1_LOC_57/A 0.01fF
C65311 INVX1_LOC_13/A INVX1_LOC_315/Y 0.00fF
C65312 NOR2X1_LOC_250/A INVX1_LOC_19/A 0.03fF
C65313 NOR2X1_LOC_147/B NOR2X1_LOC_698/Y 0.05fF
C65314 NOR2X1_LOC_91/A NAND2X1_LOC_738/B 0.03fF
C65315 NAND2X1_LOC_579/A INVX1_LOC_102/A 0.07fF
C65316 NOR2X1_LOC_454/Y NOR2X1_LOC_48/B 0.10fF
C65317 NOR2X1_LOC_219/Y INVX1_LOC_199/A 0.02fF
C65318 NOR2X1_LOC_798/A INVX1_LOC_47/Y 0.02fF
C65319 NOR2X1_LOC_689/Y INVX1_LOC_50/A 0.03fF
C65320 NOR2X1_LOC_82/A NAND2X1_LOC_63/Y 0.02fF
C65321 NOR2X1_LOC_443/Y INVX1_LOC_57/A 0.01fF
C65322 INVX1_LOC_72/A NAND2X1_LOC_210/a_36_24# 0.01fF
C65323 NOR2X1_LOC_52/B INVX1_LOC_77/Y 0.04fF
C65324 NOR2X1_LOC_512/a_36_216# INVX1_LOC_91/A 0.00fF
C65325 INVX1_LOC_77/A INVX1_LOC_54/A 0.12fF
C65326 INVX1_LOC_98/A INVX1_LOC_10/A 0.00fF
C65327 NAND2X1_LOC_184/a_36_24# INVX1_LOC_75/A 0.00fF
C65328 NOR2X1_LOC_579/a_36_216# NAND2X1_LOC_463/B 0.00fF
C65329 INVX1_LOC_143/A NAND2X1_LOC_266/a_36_24# 0.00fF
C65330 NAND2X1_LOC_363/B INVX1_LOC_26/A 0.07fF
C65331 NOR2X1_LOC_383/B INVX1_LOC_23/A 0.90fF
C65332 NOR2X1_LOC_78/A INVX1_LOC_10/A 12.02fF
C65333 NOR2X1_LOC_570/B INVX1_LOC_9/A 0.01fF
C65334 NOR2X1_LOC_778/B INVX1_LOC_37/A 0.24fF
C65335 NAND2X1_LOC_739/B NAND2X1_LOC_810/B 0.01fF
C65336 NAND2X1_LOC_208/B NAND2X1_LOC_773/B 0.10fF
C65337 INVX1_LOC_144/A NAND2X1_LOC_652/Y 0.02fF
C65338 INVX1_LOC_226/Y NAND2X1_LOC_464/A 0.00fF
C65339 INVX1_LOC_208/A NOR2X1_LOC_357/Y 0.12fF
C65340 INVX1_LOC_196/Y NAND2X1_LOC_679/a_36_24# 0.00fF
C65341 INVX1_LOC_227/A NOR2X1_LOC_405/A 0.03fF
C65342 NOR2X1_LOC_598/B INVX1_LOC_50/A 0.10fF
C65343 INVX1_LOC_58/A NOR2X1_LOC_696/Y 0.03fF
C65344 NOR2X1_LOC_82/A NAND2X1_LOC_455/B 0.76fF
C65345 NOR2X1_LOC_6/a_36_216# NAND2X1_LOC_93/B 0.00fF
C65346 INVX1_LOC_45/A INVX1_LOC_186/Y 0.51fF
C65347 INVX1_LOC_97/A INVX1_LOC_91/A 0.03fF
C65348 INVX1_LOC_69/Y INVX1_LOC_28/A 0.01fF
C65349 NOR2X1_LOC_598/B NOR2X1_LOC_105/Y 0.02fF
C65350 NAND2X1_LOC_755/a_36_24# INVX1_LOC_280/A 0.01fF
C65351 INVX1_LOC_36/A NAND2X1_LOC_479/a_36_24# 0.00fF
C65352 NOR2X1_LOC_590/A NOR2X1_LOC_841/a_36_216# 0.00fF
C65353 INVX1_LOC_89/A NOR2X1_LOC_45/B 1.72fF
C65354 NOR2X1_LOC_78/B INVX1_LOC_33/Y 0.00fF
C65355 INVX1_LOC_100/A INVX1_LOC_102/Y 0.01fF
C65356 NOR2X1_LOC_152/Y INVX1_LOC_107/Y 0.19fF
C65357 NOR2X1_LOC_355/a_36_216# INVX1_LOC_91/A 0.01fF
C65358 INVX1_LOC_64/A NOR2X1_LOC_654/A 0.02fF
C65359 INVX1_LOC_90/A INVX1_LOC_91/A 0.26fF
C65360 NOR2X1_LOC_401/A INVX1_LOC_32/A 0.44fF
C65361 NAND2X1_LOC_361/Y NOR2X1_LOC_634/A 0.01fF
C65362 INVX1_LOC_50/A NAND2X1_LOC_725/A 0.10fF
C65363 NOR2X1_LOC_791/Y INVX1_LOC_26/A 0.02fF
C65364 D_INPUT_0 NOR2X1_LOC_542/B 0.01fF
C65365 NOR2X1_LOC_389/B INVX1_LOC_91/A 0.13fF
C65366 D_INPUT_1 NOR2X1_LOC_660/Y 0.59fF
C65367 NOR2X1_LOC_460/B NAND2X1_LOC_425/Y 0.03fF
C65368 INVX1_LOC_24/A NAND2X1_LOC_456/Y 0.03fF
C65369 NAND2X1_LOC_694/a_36_24# INVX1_LOC_19/A 0.00fF
C65370 NAND2X1_LOC_466/Y NOR2X1_LOC_435/A 0.01fF
C65371 INVX1_LOC_30/Y VDD 1.30fF
C65372 INVX1_LOC_124/A INVX1_LOC_54/A 0.11fF
C65373 NOR2X1_LOC_813/Y INVX1_LOC_25/Y 0.40fF
C65374 NAND2X1_LOC_217/a_36_24# INVX1_LOC_3/A 0.01fF
C65375 NOR2X1_LOC_464/B INVX1_LOC_271/Y 0.03fF
C65376 INPUT_3 NOR2X1_LOC_554/A 0.00fF
C65377 NOR2X1_LOC_242/A NOR2X1_LOC_342/B 0.01fF
C65378 NOR2X1_LOC_68/A NOR2X1_LOC_48/Y 0.01fF
C65379 INVX1_LOC_89/A INVX1_LOC_247/A 0.03fF
C65380 INVX1_LOC_14/A NOR2X1_LOC_80/Y 0.01fF
C65381 INVX1_LOC_89/A INVX1_LOC_199/Y 0.04fF
C65382 NAND2X1_LOC_573/A NAND2X1_LOC_287/B 0.10fF
C65383 INVX1_LOC_230/Y INVX1_LOC_3/Y 0.99fF
C65384 NOR2X1_LOC_160/B INVX1_LOC_32/A 0.14fF
C65385 INVX1_LOC_254/A INVX1_LOC_63/A 0.05fF
C65386 NOR2X1_LOC_71/Y INVX1_LOC_76/A 0.07fF
C65387 GATE_479 INVX1_LOC_117/A 0.02fF
C65388 NOR2X1_LOC_82/A NAND2X1_LOC_618/Y 0.04fF
C65389 INPUT_1 INVX1_LOC_59/Y 0.35fF
C65390 INVX1_LOC_71/A INVX1_LOC_186/Y 0.08fF
C65391 INVX1_LOC_293/A NOR2X1_LOC_38/B 0.01fF
C65392 INVX1_LOC_73/Y NAND2X1_LOC_454/Y 0.01fF
C65393 INVX1_LOC_24/A INVX1_LOC_49/Y 0.08fF
C65394 NOR2X1_LOC_160/B NOR2X1_LOC_623/B -0.01fF
C65395 INVX1_LOC_177/A NOR2X1_LOC_809/B -0.00fF
C65396 NAND2X1_LOC_348/A INVX1_LOC_91/A -0.00fF
C65397 NOR2X1_LOC_644/Y INVX1_LOC_307/A 0.03fF
C65398 INVX1_LOC_22/A NOR2X1_LOC_331/B 0.20fF
C65399 NAND2X1_LOC_773/Y NAND2X1_LOC_99/A 0.10fF
C65400 INVX1_LOC_90/A NOR2X1_LOC_421/Y 0.08fF
C65401 NOR2X1_LOC_498/Y NOR2X1_LOC_485/Y 0.01fF
C65402 NOR2X1_LOC_552/A INVX1_LOC_75/A 0.01fF
C65403 INVX1_LOC_150/Y INVX1_LOC_78/A 0.07fF
C65404 NOR2X1_LOC_468/Y INVX1_LOC_181/A 0.02fF
C65405 INVX1_LOC_34/A NAND2X1_LOC_206/Y 0.02fF
C65406 NOR2X1_LOC_152/Y INVX1_LOC_272/A 0.10fF
C65407 INVX1_LOC_53/Y NOR2X1_LOC_675/a_36_216# 0.00fF
C65408 NOR2X1_LOC_763/A INVX1_LOC_23/A 0.52fF
C65409 INVX1_LOC_215/A INVX1_LOC_9/A 0.02fF
C65410 INVX1_LOC_240/A INVX1_LOC_5/Y 0.05fF
C65411 NOR2X1_LOC_53/Y NOR2X1_LOC_304/Y 0.01fF
C65412 NOR2X1_LOC_389/A INVX1_LOC_94/Y 0.01fF
C65413 NOR2X1_LOC_724/Y INVX1_LOC_37/A 0.03fF
C65414 INVX1_LOC_120/A NOR2X1_LOC_859/Y 0.02fF
C65415 INVX1_LOC_314/Y NOR2X1_LOC_178/a_36_216# 0.00fF
C65416 VDD NOR2X1_LOC_156/A 0.12fF
C65417 INVX1_LOC_34/A NAND2X1_LOC_773/B 0.08fF
C65418 NOR2X1_LOC_329/B NOR2X1_LOC_305/Y 0.20fF
C65419 NAND2X1_LOC_361/Y INVX1_LOC_29/A 0.07fF
C65420 NOR2X1_LOC_322/Y NAND2X1_LOC_241/Y 0.01fF
C65421 NOR2X1_LOC_337/Y INVX1_LOC_96/A 0.00fF
C65422 INVX1_LOC_232/A INVX1_LOC_92/A 0.10fF
C65423 INVX1_LOC_286/Y INVX1_LOC_273/A 0.01fF
C65424 INVX1_LOC_216/A NOR2X1_LOC_649/B 0.00fF
C65425 NOR2X1_LOC_65/B INVX1_LOC_150/Y 0.10fF
C65426 NAND2X1_LOC_154/Y NOR2X1_LOC_158/B 0.00fF
C65427 NOR2X1_LOC_516/Y NAND2X1_LOC_82/Y 0.01fF
C65428 NAND2X1_LOC_796/Y INVX1_LOC_54/A 0.08fF
C65429 INVX1_LOC_22/A NOR2X1_LOC_491/Y 0.31fF
C65430 NOR2X1_LOC_122/Y NOR2X1_LOC_363/Y 0.25fF
C65431 INVX1_LOC_22/A NOR2X1_LOC_592/B 0.05fF
C65432 INVX1_LOC_77/A NOR2X1_LOC_48/B 0.07fF
C65433 NOR2X1_LOC_742/A INVX1_LOC_14/Y 0.09fF
C65434 NAND2X1_LOC_672/B NAND2X1_LOC_574/A 0.02fF
C65435 INVX1_LOC_190/A INVX1_LOC_54/A 0.04fF
C65436 INVX1_LOC_219/Y INVX1_LOC_29/A 0.01fF
C65437 NOR2X1_LOC_709/A INVX1_LOC_19/A 0.00fF
C65438 NOR2X1_LOC_186/Y NAND2X1_LOC_474/Y 0.00fF
C65439 NOR2X1_LOC_487/a_36_216# INVX1_LOC_78/A 0.00fF
C65440 INVX1_LOC_69/Y NOR2X1_LOC_35/Y 0.10fF
C65441 INVX1_LOC_163/A INVX1_LOC_253/Y 0.13fF
C65442 INVX1_LOC_30/A INVX1_LOC_26/A 0.24fF
C65443 NOR2X1_LOC_142/Y INVX1_LOC_290/Y 0.10fF
C65444 NAND2X1_LOC_656/Y NAND2X1_LOC_656/B 0.09fF
C65445 INVX1_LOC_14/A NOR2X1_LOC_109/Y 0.52fF
C65446 INVX1_LOC_58/A INVX1_LOC_230/Y 0.01fF
C65447 NAND2X1_LOC_49/a_36_24# INVX1_LOC_84/A 0.00fF
C65448 NOR2X1_LOC_457/B NOR2X1_LOC_464/Y 0.28fF
C65449 NOR2X1_LOC_91/A INVX1_LOC_57/Y 0.20fF
C65450 INVX1_LOC_77/A NAND2X1_LOC_3/B 0.17fF
C65451 NAND2X1_LOC_363/B NOR2X1_LOC_107/Y 0.06fF
C65452 INPUT_0 NAND2X1_LOC_472/Y 0.03fF
C65453 NOR2X1_LOC_632/Y NOR2X1_LOC_66/Y 0.01fF
C65454 INVX1_LOC_287/A INVX1_LOC_45/A 0.00fF
C65455 NOR2X1_LOC_716/B INVX1_LOC_4/A 1.29fF
C65456 NOR2X1_LOC_123/a_36_216# NOR2X1_LOC_124/A 0.02fF
C65457 INVX1_LOC_120/A INVX1_LOC_46/Y -0.00fF
C65458 NOR2X1_LOC_45/B NOR2X1_LOC_24/Y 0.02fF
C65459 INVX1_LOC_75/A INVX1_LOC_280/A 0.07fF
C65460 INVX1_LOC_89/A NOR2X1_LOC_862/B 0.05fF
C65461 INVX1_LOC_79/A INVX1_LOC_38/A 0.07fF
C65462 NAND2X1_LOC_156/B NOR2X1_LOC_697/Y 0.01fF
C65463 NOR2X1_LOC_45/B NAND2X1_LOC_244/A 0.01fF
C65464 INVX1_LOC_96/A VDD 0.46fF
C65465 NOR2X1_LOC_78/A NOR2X1_LOC_850/a_36_216# 0.02fF
C65466 INVX1_LOC_34/A NOR2X1_LOC_297/A 0.01fF
C65467 NAND2X1_LOC_541/Y INVX1_LOC_12/A 0.01fF
C65468 INVX1_LOC_21/A INVX1_LOC_269/A 0.23fF
C65469 INVX1_LOC_132/Y NAND2X1_LOC_412/a_36_24# 0.00fF
C65470 INVX1_LOC_21/A NOR2X1_LOC_232/Y 0.01fF
C65471 NOR2X1_LOC_655/B INVX1_LOC_290/Y 0.05fF
C65472 NOR2X1_LOC_332/A NOR2X1_LOC_673/A 0.07fF
C65473 INVX1_LOC_63/Y NOR2X1_LOC_158/B 0.01fF
C65474 NOR2X1_LOC_703/a_36_216# INVX1_LOC_292/Y 0.01fF
C65475 INVX1_LOC_136/A D_INPUT_1 3.38fF
C65476 NAND2X1_LOC_849/B INVX1_LOC_309/A -0.03fF
C65477 INVX1_LOC_39/A NOR2X1_LOC_82/A 0.13fF
C65478 NAND2X1_LOC_659/B NAND2X1_LOC_658/a_36_24# 0.02fF
C65479 INVX1_LOC_309/A INVX1_LOC_38/A 0.03fF
C65480 NOR2X1_LOC_1/a_36_216# D_INPUT_5 0.00fF
C65481 INVX1_LOC_65/A NOR2X1_LOC_858/B 0.25fF
C65482 NOR2X1_LOC_770/B INVX1_LOC_78/A 0.03fF
C65483 NOR2X1_LOC_295/Y INVX1_LOC_94/Y 0.01fF
C65484 INVX1_LOC_16/A NOR2X1_LOC_89/A 0.36fF
C65485 NAND2X1_LOC_832/Y INVX1_LOC_54/A 0.32fF
C65486 VDD NOR2X1_LOC_124/A 0.35fF
C65487 INVX1_LOC_13/A NAND2X1_LOC_207/B 0.07fF
C65488 NOR2X1_LOC_750/Y NOR2X1_LOC_68/A -0.01fF
C65489 INVX1_LOC_139/A NAND2X1_LOC_212/Y 0.32fF
C65490 NAND2X1_LOC_149/Y INVX1_LOC_11/A 2.09fF
C65491 VDD INVX1_LOC_188/Y 0.21fF
C65492 NOR2X1_LOC_311/Y INVX1_LOC_33/Y 0.01fF
C65493 NOR2X1_LOC_542/Y NOR2X1_LOC_814/A 0.05fF
C65494 INVX1_LOC_18/A NAND2X1_LOC_793/B 0.07fF
C65495 NAND2X1_LOC_783/A INVX1_LOC_49/Y 0.01fF
C65496 NOR2X1_LOC_577/Y NOR2X1_LOC_106/a_36_216# 0.00fF
C65497 INVX1_LOC_266/Y NOR2X1_LOC_334/Y 0.08fF
C65498 INVX1_LOC_90/A INVX1_LOC_203/A 0.03fF
C65499 INVX1_LOC_91/A INVX1_LOC_38/A 5.07fF
C65500 NOR2X1_LOC_130/A INVX1_LOC_49/Y 0.06fF
C65501 NAND2X1_LOC_633/Y INVX1_LOC_20/A 0.28fF
C65502 NOR2X1_LOC_357/Y NAND2X1_LOC_211/Y 0.05fF
C65503 INVX1_LOC_82/Y NAND2X1_LOC_574/A 0.03fF
C65504 NAND2X1_LOC_721/B NOR2X1_LOC_406/A 0.02fF
C65505 INVX1_LOC_219/A NOR2X1_LOC_671/Y 0.01fF
C65506 NOR2X1_LOC_759/Y NOR2X1_LOC_678/A 0.02fF
C65507 INVX1_LOC_125/Y NOR2X1_LOC_489/A 0.11fF
C65508 NOR2X1_LOC_577/Y NOR2X1_LOC_493/A 0.01fF
C65509 NOR2X1_LOC_516/B INVX1_LOC_32/A 0.03fF
C65510 NAND2X1_LOC_661/B NOR2X1_LOC_158/Y 0.00fF
C65511 NAND2X1_LOC_96/A NAND2X1_LOC_411/a_36_24# 0.00fF
C65512 INVX1_LOC_202/A NOR2X1_LOC_678/A 0.01fF
C65513 INVX1_LOC_204/Y NOR2X1_LOC_68/A 0.03fF
C65514 INVX1_LOC_136/A NOR2X1_LOC_652/Y 0.09fF
C65515 D_INPUT_2 NOR2X1_LOC_660/Y 0.04fF
C65516 INVX1_LOC_11/Y INVX1_LOC_38/A 0.03fF
C65517 INVX1_LOC_59/A NAND2X1_LOC_577/A 0.16fF
C65518 NOR2X1_LOC_778/B NAND2X1_LOC_72/B 0.04fF
C65519 NOR2X1_LOC_852/A NOR2X1_LOC_852/Y 0.17fF
C65520 INVX1_LOC_278/A NOR2X1_LOC_237/a_36_216# 0.01fF
C65521 NOR2X1_LOC_606/Y INVX1_LOC_48/Y 0.32fF
C65522 INVX1_LOC_172/A NAND2X1_LOC_793/B 0.07fF
C65523 INVX1_LOC_41/A INVX1_LOC_29/Y 0.03fF
C65524 NOR2X1_LOC_250/A INVX1_LOC_161/Y 0.02fF
C65525 INVX1_LOC_50/A NAND2X1_LOC_308/Y 0.01fF
C65526 NOR2X1_LOC_550/B NOR2X1_LOC_678/A 0.03fF
C65527 NOR2X1_LOC_7/Y INVX1_LOC_117/Y 0.01fF
C65528 NOR2X1_LOC_272/Y INVX1_LOC_177/Y 0.09fF
C65529 NOR2X1_LOC_294/Y NAND2X1_LOC_473/A 0.44fF
C65530 NOR2X1_LOC_15/Y INVX1_LOC_286/Y 0.07fF
C65531 INVX1_LOC_33/Y INVX1_LOC_46/A 0.03fF
C65532 NOR2X1_LOC_180/Y NOR2X1_LOC_748/A 0.05fF
C65533 NAND2X1_LOC_537/Y INVX1_LOC_141/Y 0.02fF
C65534 NOR2X1_LOC_78/B INVX1_LOC_23/Y 0.08fF
C65535 NAND2X1_LOC_654/B INVX1_LOC_29/A 0.48fF
C65536 NOR2X1_LOC_78/A INVX1_LOC_307/A 0.00fF
C65537 NOR2X1_LOC_335/B NOR2X1_LOC_814/A 0.24fF
C65538 NAND2X1_LOC_853/Y NAND2X1_LOC_175/Y 0.86fF
C65539 NOR2X1_LOC_229/Y NOR2X1_LOC_158/Y 0.05fF
C65540 NOR2X1_LOC_353/Y NOR2X1_LOC_727/B 0.00fF
C65541 NOR2X1_LOC_71/Y INVX1_LOC_127/Y 0.00fF
C65542 NOR2X1_LOC_860/B INVX1_LOC_38/Y 0.00fF
C65543 INVX1_LOC_6/A NOR2X1_LOC_127/Y 0.07fF
C65544 VDD NOR2X1_LOC_684/Y 0.35fF
C65545 INVX1_LOC_50/A NAND2X1_LOC_660/A 0.13fF
C65546 NAND2X1_LOC_537/Y INVX1_LOC_312/Y 0.02fF
C65547 INVX1_LOC_36/A INVX1_LOC_14/A 0.31fF
C65548 INVX1_LOC_28/A NOR2X1_LOC_89/A 0.16fF
C65549 NOR2X1_LOC_78/A NOR2X1_LOC_445/B 0.08fF
C65550 INVX1_LOC_224/Y INVX1_LOC_34/Y 0.34fF
C65551 INPUT_3 NOR2X1_LOC_160/B 0.03fF
C65552 INPUT_0 NAND2X1_LOC_773/B 0.07fF
C65553 NOR2X1_LOC_717/B INVX1_LOC_4/A 0.03fF
C65554 INVX1_LOC_45/A NAND2X1_LOC_154/a_36_24# 0.01fF
C65555 NAND2X1_LOC_787/A NOR2X1_LOC_369/a_36_216# 0.00fF
C65556 INVX1_LOC_22/A NOR2X1_LOC_449/A 2.49fF
C65557 NOR2X1_LOC_168/A INVX1_LOC_23/A 0.01fF
C65558 NOR2X1_LOC_719/A INVX1_LOC_16/Y 0.32fF
C65559 NAND2X1_LOC_447/Y INVX1_LOC_92/A 0.04fF
C65560 NOR2X1_LOC_91/A NAND2X1_LOC_170/A 0.36fF
C65561 INVX1_LOC_182/A INVX1_LOC_290/Y 0.09fF
C65562 NAND2X1_LOC_334/a_36_24# NAND2X1_LOC_464/B 0.00fF
C65563 NAND2X1_LOC_773/Y NAND2X1_LOC_656/A 0.08fF
C65564 INVX1_LOC_89/Y INVX1_LOC_76/A 0.04fF
C65565 NOR2X1_LOC_98/B NAND2X1_LOC_93/a_36_24# 0.02fF
C65566 NOR2X1_LOC_15/Y NOR2X1_LOC_191/B 0.01fF
C65567 INVX1_LOC_54/Y NOR2X1_LOC_717/A 0.21fF
C65568 NOR2X1_LOC_684/a_36_216# NOR2X1_LOC_684/Y 0.00fF
C65569 NAND2X1_LOC_842/B INVX1_LOC_47/Y 0.11fF
C65570 INVX1_LOC_235/Y NOR2X1_LOC_474/A 0.76fF
C65571 NOR2X1_LOC_168/B NOR2X1_LOC_634/Y 0.36fF
C65572 NOR2X1_LOC_541/Y INVX1_LOC_18/A 0.02fF
C65573 NOR2X1_LOC_82/A INVX1_LOC_61/A 0.07fF
C65574 INVX1_LOC_89/A NOR2X1_LOC_685/B 0.02fF
C65575 INVX1_LOC_58/A NAND2X1_LOC_341/A 0.05fF
C65576 INVX1_LOC_11/A NOR2X1_LOC_744/Y 0.01fF
C65577 INVX1_LOC_57/Y INVX1_LOC_31/A 0.09fF
C65578 NOR2X1_LOC_719/A NAND2X1_LOC_205/A 0.15fF
C65579 NOR2X1_LOC_237/Y INVX1_LOC_14/A 1.75fF
C65580 NOR2X1_LOC_256/Y INVX1_LOC_3/Y 0.05fF
C65581 INVX1_LOC_225/A NAND2X1_LOC_474/Y 0.01fF
C65582 NOR2X1_LOC_737/a_36_216# INVX1_LOC_12/A 0.00fF
C65583 NOR2X1_LOC_272/Y INVX1_LOC_104/A 0.60fF
C65584 INVX1_LOC_177/A INVX1_LOC_50/Y 0.03fF
C65585 INVX1_LOC_64/A NOR2X1_LOC_757/Y 0.01fF
C65586 INVX1_LOC_36/A NOR2X1_LOC_717/Y 0.01fF
C65587 INVX1_LOC_35/A NOR2X1_LOC_287/A 0.03fF
C65588 INVX1_LOC_277/A INVX1_LOC_142/A 0.18fF
C65589 INVX1_LOC_103/A INVX1_LOC_49/A 0.07fF
C65590 NOR2X1_LOC_792/a_36_216# NOR2X1_LOC_309/Y 0.01fF
C65591 NOR2X1_LOC_757/A INVX1_LOC_271/A 0.07fF
C65592 NOR2X1_LOC_151/Y INVX1_LOC_4/A 0.03fF
C65593 INVX1_LOC_31/A NOR2X1_LOC_512/Y 0.01fF
C65594 INVX1_LOC_54/A INVX1_LOC_9/A 0.11fF
C65595 INVX1_LOC_45/A INVX1_LOC_18/A 13.49fF
C65596 NOR2X1_LOC_78/A INVX1_LOC_12/A 0.06fF
C65597 NAND2X1_LOC_355/a_36_24# INVX1_LOC_159/A 0.00fF
C65598 INVX1_LOC_302/Y NOR2X1_LOC_158/B 0.00fF
C65599 NOR2X1_LOC_137/A INVX1_LOC_270/A 0.10fF
C65600 NOR2X1_LOC_15/Y INVX1_LOC_185/Y 0.01fF
C65601 INVX1_LOC_72/A NAND2X1_LOC_16/Y -0.02fF
C65602 INVX1_LOC_18/A NOR2X1_LOC_568/A 0.08fF
C65603 NOR2X1_LOC_276/B INVX1_LOC_30/A 0.02fF
C65604 INVX1_LOC_24/A NAND2X1_LOC_208/B 0.01fF
C65605 INVX1_LOC_14/A NOR2X1_LOC_309/Y 0.37fF
C65606 NOR2X1_LOC_468/Y NOR2X1_LOC_315/Y 1.29fF
C65607 INVX1_LOC_292/A INVX1_LOC_49/A 0.01fF
C65608 NAND2X1_LOC_784/a_36_24# NOR2X1_LOC_667/A -0.02fF
C65609 INVX1_LOC_266/A INVX1_LOC_177/A 0.00fF
C65610 NAND2X1_LOC_739/B INVX1_LOC_36/A 0.03fF
C65611 NOR2X1_LOC_208/Y NOR2X1_LOC_717/Y 0.14fF
C65612 NOR2X1_LOC_151/a_36_216# NAND2X1_LOC_454/Y 0.01fF
C65613 NOR2X1_LOC_441/Y INVX1_LOC_77/A 0.01fF
C65614 NOR2X1_LOC_242/A NOR2X1_LOC_244/B 0.01fF
C65615 NOR2X1_LOC_471/Y INVX1_LOC_63/Y 0.10fF
C65616 NOR2X1_LOC_607/A INVX1_LOC_72/A 0.03fF
C65617 NOR2X1_LOC_438/a_36_216# NOR2X1_LOC_52/B 0.00fF
C65618 INVX1_LOC_176/A NAND2X1_LOC_63/Y 0.05fF
C65619 INVX1_LOC_24/A NOR2X1_LOC_722/Y 0.01fF
C65620 INVX1_LOC_72/A NOR2X1_LOC_95/a_36_216# 0.00fF
C65621 INVX1_LOC_64/A NOR2X1_LOC_717/B 1.92fF
C65622 INVX1_LOC_136/A NOR2X1_LOC_403/B 0.03fF
C65623 INVX1_LOC_2/A INVX1_LOC_103/A 0.15fF
C65624 NOR2X1_LOC_389/A INVX1_LOC_162/A 0.17fF
C65625 INVX1_LOC_18/A INVX1_LOC_71/A 0.19fF
C65626 NAND2X1_LOC_465/A NAND2X1_LOC_254/Y 0.01fF
C65627 INVX1_LOC_299/A NOR2X1_LOC_220/A 0.10fF
C65628 NOR2X1_LOC_265/a_36_216# NOR2X1_LOC_15/Y 0.00fF
C65629 NAND2X1_LOC_633/a_36_24# NAND2X1_LOC_793/Y 0.00fF
C65630 NOR2X1_LOC_178/Y NOR2X1_LOC_71/Y 0.28fF
C65631 NOR2X1_LOC_226/A INVX1_LOC_103/A 0.16fF
C65632 NAND2X1_LOC_53/Y NOR2X1_LOC_209/Y 0.04fF
C65633 NOR2X1_LOC_455/Y NOR2X1_LOC_644/A 0.02fF
C65634 NOR2X1_LOC_186/Y INVX1_LOC_10/A 0.12fF
C65635 NOR2X1_LOC_858/B NOR2X1_LOC_830/Y 0.25fF
C65636 NOR2X1_LOC_790/B NOR2X1_LOC_356/A 0.09fF
C65637 NOR2X1_LOC_740/Y NOR2X1_LOC_307/B 0.08fF
C65638 INVX1_LOC_58/A NAND2X1_LOC_740/B 0.03fF
C65639 INVX1_LOC_255/Y INVX1_LOC_163/A 0.01fF
C65640 NAND2X1_LOC_543/Y NAND2X1_LOC_579/A 0.03fF
C65641 NAND2X1_LOC_751/a_36_24# NOR2X1_LOC_750/A 0.00fF
C65642 INVX1_LOC_92/A NAND2X1_LOC_750/a_36_24# 0.00fF
C65643 INVX1_LOC_33/A NOR2X1_LOC_703/B 0.00fF
C65644 INVX1_LOC_2/A INVX1_LOC_292/A 0.07fF
C65645 NOR2X1_LOC_446/A NOR2X1_LOC_78/B 0.17fF
C65646 INVX1_LOC_83/A NOR2X1_LOC_846/A 0.03fF
C65647 NAND2X1_LOC_21/Y NAND2X1_LOC_588/B 0.13fF
C65648 INVX1_LOC_5/A INVX1_LOC_20/Y 0.00fF
C65649 NAND2X1_LOC_796/B NAND2X1_LOC_808/A 0.06fF
C65650 NOR2X1_LOC_218/Y INVX1_LOC_103/A 0.02fF
C65651 INVX1_LOC_12/A NOR2X1_LOC_60/Y 0.00fF
C65652 INVX1_LOC_139/Y INVX1_LOC_283/A 0.00fF
C65653 INVX1_LOC_39/A NOR2X1_LOC_132/a_36_216# 0.00fF
C65654 INVX1_LOC_6/A NOR2X1_LOC_383/B 0.21fF
C65655 INVX1_LOC_11/A INVX1_LOC_16/A 0.06fF
C65656 NOR2X1_LOC_387/A INVX1_LOC_296/Y 0.05fF
C65657 NAND2X1_LOC_637/Y NOR2X1_LOC_48/a_36_216# 0.00fF
C65658 INVX1_LOC_32/A NAND2X1_LOC_211/Y 0.01fF
C65659 NOR2X1_LOC_807/B NOR2X1_LOC_374/B 0.16fF
C65660 INVX1_LOC_149/A INVX1_LOC_30/A 0.32fF
C65661 INVX1_LOC_36/A NOR2X1_LOC_612/B 0.14fF
C65662 NAND2X1_LOC_170/a_36_24# INVX1_LOC_90/A 0.01fF
C65663 NOR2X1_LOC_88/Y INVX1_LOC_285/A 0.07fF
C65664 NOR2X1_LOC_790/B NOR2X1_LOC_74/A 0.80fF
C65665 NAND2X1_LOC_724/A INVX1_LOC_10/A 0.08fF
C65666 NAND2X1_LOC_364/A INVX1_LOC_104/A 0.09fF
C65667 INVX1_LOC_210/Y INVX1_LOC_210/A 0.05fF
C65668 INVX1_LOC_34/A INVX1_LOC_24/A 0.35fF
C65669 INVX1_LOC_280/A NAND2X1_LOC_291/B 0.01fF
C65670 NAND2X1_LOC_192/a_36_24# NOR2X1_LOC_665/A 0.01fF
C65671 NAND2X1_LOC_655/B INVX1_LOC_94/Y 0.02fF
C65672 INVX1_LOC_256/A INVX1_LOC_290/A 0.04fF
C65673 NOR2X1_LOC_546/B NOR2X1_LOC_486/B 0.04fF
C65674 NAND2X1_LOC_192/B INVX1_LOC_279/A 0.03fF
C65675 NAND2X1_LOC_9/Y NOR2X1_LOC_775/a_36_216# 0.00fF
C65676 INVX1_LOC_181/Y NOR2X1_LOC_192/a_36_216# 0.00fF
C65677 NAND2X1_LOC_499/a_36_24# INVX1_LOC_118/A 0.00fF
C65678 NAND2X1_LOC_848/Y INVX1_LOC_203/A 0.05fF
C65679 INPUT_3 NOR2X1_LOC_516/B 3.08fF
C65680 INVX1_LOC_286/Y NAND2X1_LOC_840/B 0.07fF
C65681 INVX1_LOC_225/Y NOR2X1_LOC_569/Y 0.06fF
C65682 INVX1_LOC_77/A NOR2X1_LOC_142/Y 1.58fF
C65683 NAND2X1_LOC_84/Y NOR2X1_LOC_309/Y 0.03fF
C65684 NAND2X1_LOC_639/A NOR2X1_LOC_467/A 0.20fF
C65685 NAND2X1_LOC_468/B NAND2X1_LOC_61/Y 0.01fF
C65686 NOR2X1_LOC_388/Y NOR2X1_LOC_577/Y 1.20fF
C65687 INVX1_LOC_84/A INVX1_LOC_285/A 0.65fF
C65688 INVX1_LOC_226/Y INVX1_LOC_170/A 0.02fF
C65689 NOR2X1_LOC_718/Y INVX1_LOC_153/Y 0.06fF
C65690 VDD INVX1_LOC_273/A 0.13fF
C65691 INVX1_LOC_275/A NOR2X1_LOC_486/B 0.04fF
C65692 NAND2X1_LOC_169/Y NOR2X1_LOC_74/A 0.05fF
C65693 NAND2X1_LOC_361/Y INVX1_LOC_8/A 0.03fF
C65694 INVX1_LOC_129/Y INVX1_LOC_4/Y 0.01fF
C65695 NAND2X1_LOC_96/A NOR2X1_LOC_38/B 0.04fF
C65696 INVX1_LOC_186/A INVX1_LOC_53/A 0.06fF
C65697 INVX1_LOC_34/A NOR2X1_LOC_557/Y 1.25fF
C65698 INVX1_LOC_16/Y INVX1_LOC_76/A 0.09fF
C65699 INVX1_LOC_84/A NOR2X1_LOC_814/A 0.07fF
C65700 INVX1_LOC_103/A NAND2X1_LOC_648/A 0.03fF
C65701 NOR2X1_LOC_45/Y INVX1_LOC_10/A 0.07fF
C65702 NAND2X1_LOC_800/A INVX1_LOC_273/A 0.01fF
C65703 NOR2X1_LOC_432/Y NOR2X1_LOC_596/A 0.01fF
C65704 D_GATE_479 INVX1_LOC_175/A 0.00fF
C65705 NOR2X1_LOC_96/a_36_216# INVX1_LOC_3/Y 0.01fF
C65706 INVX1_LOC_161/Y NOR2X1_LOC_106/A 0.01fF
C65707 NOR2X1_LOC_791/Y NOR2X1_LOC_368/A 0.01fF
C65708 NAND2X1_LOC_350/A INVX1_LOC_190/A 0.02fF
C65709 INVX1_LOC_71/A INVX1_LOC_34/Y 0.32fF
C65710 NOR2X1_LOC_45/B NOR2X1_LOC_392/Y 0.01fF
C65711 INVX1_LOC_90/A NOR2X1_LOC_592/A 0.02fF
C65712 INVX1_LOC_161/A NAND2X1_LOC_800/Y 0.10fF
C65713 INVX1_LOC_46/A INVX1_LOC_23/Y 0.01fF
C65714 NOR2X1_LOC_461/A NOR2X1_LOC_461/Y 0.16fF
C65715 NOR2X1_LOC_655/B INVX1_LOC_77/A 0.01fF
C65716 NOR2X1_LOC_135/Y INVX1_LOC_88/A 0.02fF
C65717 INVX1_LOC_11/A INVX1_LOC_28/A 0.09fF
C65718 INVX1_LOC_124/A NOR2X1_LOC_142/Y 0.10fF
C65719 NAND2X1_LOC_192/B INVX1_LOC_182/Y 0.01fF
C65720 INVX1_LOC_76/A NAND2X1_LOC_205/A 0.10fF
C65721 INVX1_LOC_53/A NAND2X1_LOC_447/Y 0.10fF
C65722 INVX1_LOC_58/A NOR2X1_LOC_331/a_36_216# 0.00fF
C65723 NOR2X1_LOC_366/B NOR2X1_LOC_577/Y 0.00fF
C65724 INVX1_LOC_20/A NOR2X1_LOC_591/A 0.02fF
C65725 NOR2X1_LOC_781/Y INVX1_LOC_290/A 0.04fF
C65726 INVX1_LOC_314/Y INVX1_LOC_53/Y 0.03fF
C65727 INVX1_LOC_271/A INVX1_LOC_37/A 0.12fF
C65728 NOR2X1_LOC_718/B INVX1_LOC_266/Y 0.03fF
C65729 NOR2X1_LOC_364/A INVX1_LOC_15/A 0.61fF
C65730 NOR2X1_LOC_78/B NOR2X1_LOC_722/a_36_216# 0.00fF
C65731 INVX1_LOC_111/Y NOR2X1_LOC_309/Y 0.26fF
C65732 NOR2X1_LOC_673/A INVX1_LOC_42/A 0.00fF
C65733 D_GATE_741 NOR2X1_LOC_74/A 0.02fF
C65734 NAND2X1_LOC_559/a_36_24# INVX1_LOC_229/Y 0.07fF
C65735 NAND2X1_LOC_717/Y NAND2X1_LOC_838/Y 0.00fF
C65736 NOR2X1_LOC_593/Y INVX1_LOC_16/A 0.04fF
C65737 NOR2X1_LOC_419/Y NOR2X1_LOC_721/a_36_216# 0.00fF
C65738 NAND2X1_LOC_474/Y NAND2X1_LOC_642/Y 0.05fF
C65739 INVX1_LOC_238/Y NOR2X1_LOC_380/Y 0.91fF
C65740 INVX1_LOC_285/A INVX1_LOC_15/A 0.07fF
C65741 NOR2X1_LOC_826/Y NAND2X1_LOC_721/A 0.01fF
C65742 NOR2X1_LOC_541/Y NOR2X1_LOC_548/A 0.36fF
C65743 INVX1_LOC_57/Y NAND2X1_LOC_807/Y 0.01fF
C65744 INVX1_LOC_25/A NOR2X1_LOC_536/A 0.10fF
C65745 INVX1_LOC_194/A INVX1_LOC_197/Y 0.41fF
C65746 INVX1_LOC_39/A INVX1_LOC_59/Y 0.15fF
C65747 INVX1_LOC_136/A NOR2X1_LOC_497/Y 0.39fF
C65748 INVX1_LOC_15/A NOR2X1_LOC_814/A 1.07fF
C65749 NOR2X1_LOC_401/B NOR2X1_LOC_401/Y 0.02fF
C65750 NOR2X1_LOC_65/B NOR2X1_LOC_612/Y 0.02fF
C65751 NOR2X1_LOC_590/A NOR2X1_LOC_335/B 0.07fF
C65752 NAND2X1_LOC_149/Y INVX1_LOC_199/A 0.05fF
C65753 INVX1_LOC_98/Y NAND2X1_LOC_850/Y 0.01fF
C65754 INVX1_LOC_77/A NOR2X1_LOC_99/B 0.11fF
C65755 NOR2X1_LOC_607/A INVX1_LOC_313/Y 0.00fF
C65756 NOR2X1_LOC_481/A INVX1_LOC_10/A 0.01fF
C65757 NOR2X1_LOC_52/B INVX1_LOC_16/A 0.10fF
C65758 NAND2X1_LOC_352/B NOR2X1_LOC_9/Y 0.01fF
C65759 INVX1_LOC_135/A NOR2X1_LOC_577/Y 0.10fF
C65760 INVX1_LOC_245/Y NOR2X1_LOC_377/a_36_216# 0.00fF
C65761 NAND2X1_LOC_35/Y INVX1_LOC_37/Y 0.02fF
C65762 NOR2X1_LOC_445/Y INVX1_LOC_227/A 0.02fF
C65763 INVX1_LOC_213/Y NOR2X1_LOC_730/Y 0.01fF
C65764 NAND2X1_LOC_343/a_36_24# NOR2X1_LOC_52/B 0.00fF
C65765 NAND2X1_LOC_778/Y VDD 1.10fF
C65766 INVX1_LOC_269/A INVX1_LOC_255/A 0.02fF
C65767 NOR2X1_LOC_15/Y NOR2X1_LOC_56/Y 0.03fF
C65768 NOR2X1_LOC_381/Y INVX1_LOC_316/A 0.01fF
C65769 NOR2X1_LOC_15/Y NAND2X1_LOC_659/B 0.07fF
C65770 NOR2X1_LOC_361/B NOR2X1_LOC_124/A 0.01fF
C65771 INVX1_LOC_25/A NOR2X1_LOC_655/Y 0.01fF
C65772 NOR2X1_LOC_244/B NOR2X1_LOC_78/B 0.11fF
C65773 INVX1_LOC_225/A INVX1_LOC_10/A 0.07fF
C65774 INVX1_LOC_34/A NAND2X1_LOC_800/Y 0.03fF
C65775 NOR2X1_LOC_594/Y NAND2X1_LOC_154/Y 0.04fF
C65776 INPUT_3 INVX1_LOC_315/Y 0.02fF
C65777 INVX1_LOC_34/A NOR2X1_LOC_130/A 0.01fF
C65778 INVX1_LOC_27/A INVX1_LOC_37/A 0.14fF
C65779 NAND2X1_LOC_784/A INVX1_LOC_185/A 0.00fF
C65780 NOR2X1_LOC_568/A NOR2X1_LOC_548/A 0.00fF
C65781 NOR2X1_LOC_824/A INVX1_LOC_37/A 0.08fF
C65782 NOR2X1_LOC_78/B INVX1_LOC_232/A 0.35fF
C65783 INVX1_LOC_21/A INVX1_LOC_12/Y 0.01fF
C65784 INVX1_LOC_25/A NAND2X1_LOC_93/B 0.07fF
C65785 NOR2X1_LOC_629/B INVX1_LOC_135/A 0.03fF
C65786 NOR2X1_LOC_232/Y NOR2X1_LOC_670/Y 0.01fF
C65787 INVX1_LOC_83/A NAND2X1_LOC_116/A 0.03fF
C65788 NOR2X1_LOC_433/A INVX1_LOC_28/A 0.18fF
C65789 INVX1_LOC_57/Y INVX1_LOC_6/A 0.22fF
C65790 NAND2X1_LOC_276/Y INVX1_LOC_90/A 0.00fF
C65791 INVX1_LOC_23/A INVX1_LOC_179/A 0.03fF
C65792 NOR2X1_LOC_334/Y INVX1_LOC_19/A 0.08fF
C65793 NAND2X1_LOC_569/A NAND2X1_LOC_551/A 0.01fF
C65794 INVX1_LOC_224/A NOR2X1_LOC_35/Y 0.03fF
C65795 NOR2X1_LOC_91/A INVX1_LOC_250/Y 0.04fF
C65796 NOR2X1_LOC_15/Y VDD 3.27fF
C65797 NOR2X1_LOC_364/Y D_GATE_366 0.01fF
C65798 INVX1_LOC_223/A NOR2X1_LOC_501/B 0.01fF
C65799 INVX1_LOC_13/Y NAND2X1_LOC_297/a_36_24# 0.01fF
C65800 NOR2X1_LOC_92/Y NOR2X1_LOC_111/A 0.07fF
C65801 NOR2X1_LOC_15/Y NAND2X1_LOC_800/A 0.03fF
C65802 INVX1_LOC_11/A NOR2X1_LOC_35/Y 0.01fF
C65803 INVX1_LOC_89/A NOR2X1_LOC_180/Y 0.03fF
C65804 INVX1_LOC_24/A INPUT_0 0.14fF
C65805 NAND2X1_LOC_703/Y INVX1_LOC_33/Y 0.12fF
C65806 INVX1_LOC_13/A INVX1_LOC_316/Y 0.01fF
C65807 INVX1_LOC_129/A NAND2X1_LOC_572/B 0.08fF
C65808 NAND2X1_LOC_479/Y INVX1_LOC_22/A 1.20fF
C65809 NAND2X1_LOC_231/Y NOR2X1_LOC_130/A 0.04fF
C65810 INVX1_LOC_71/A NOR2X1_LOC_548/A 0.03fF
C65811 NOR2X1_LOC_284/B INVX1_LOC_83/A 0.01fF
C65812 INVX1_LOC_10/A NAND2X1_LOC_852/Y 0.10fF
C65813 NOR2X1_LOC_82/A D_INPUT_3 0.24fF
C65814 INVX1_LOC_25/A NOR2X1_LOC_649/B 0.29fF
C65815 NOR2X1_LOC_15/Y NAND2X1_LOC_463/a_36_24# 0.00fF
C65816 INVX1_LOC_135/A NOR2X1_LOC_346/B 0.00fF
C65817 NOR2X1_LOC_716/B INVX1_LOC_282/A 0.04fF
C65818 NAND2X1_LOC_593/Y NOR2X1_LOC_815/A 0.02fF
C65819 INVX1_LOC_25/A INVX1_LOC_3/A 0.64fF
C65820 INVX1_LOC_33/A INVX1_LOC_79/A 0.46fF
C65821 INVX1_LOC_28/A NOR2X1_LOC_52/B 1.14fF
C65822 NAND2X1_LOC_276/Y NAND2X1_LOC_348/A 0.03fF
C65823 INVX1_LOC_1/A NOR2X1_LOC_536/A 0.07fF
C65824 NOR2X1_LOC_25/Y NOR2X1_LOC_18/a_36_216# 0.00fF
C65825 NOR2X1_LOC_409/B INVX1_LOC_42/A 0.31fF
C65826 INVX1_LOC_90/A NAND2X1_LOC_374/Y 0.07fF
C65827 NOR2X1_LOC_344/A NOR2X1_LOC_74/A 0.02fF
C65828 NOR2X1_LOC_596/Y INVX1_LOC_46/A 0.00fF
C65829 NOR2X1_LOC_391/A NAND2X1_LOC_666/a_36_24# 0.01fF
C65830 NOR2X1_LOC_594/Y INVX1_LOC_63/Y 0.01fF
C65831 INVX1_LOC_108/Y NOR2X1_LOC_814/A 0.32fF
C65832 NOR2X1_LOC_383/B INVX1_LOC_301/A 0.10fF
C65833 NOR2X1_LOC_209/Y NOR2X1_LOC_302/Y 0.02fF
C65834 INVX1_LOC_50/A INVX1_LOC_29/A 0.06fF
C65835 NAND2X1_LOC_355/a_36_24# INVX1_LOC_146/Y 0.00fF
C65836 NAND2X1_LOC_470/B NOR2X1_LOC_467/A 0.05fF
C65837 INVX1_LOC_295/A INVX1_LOC_22/A 0.03fF
C65838 INVX1_LOC_14/A NOR2X1_LOC_656/Y 0.07fF
C65839 NOR2X1_LOC_489/a_36_216# NOR2X1_LOC_814/A 0.01fF
C65840 NAND2X1_LOC_35/Y NOR2X1_LOC_485/Y 0.01fF
C65841 NAND2X1_LOC_741/B INVX1_LOC_46/A 0.03fF
C65842 INVX1_LOC_103/A INVX1_LOC_118/A 0.12fF
C65843 INVX1_LOC_61/A INVX1_LOC_59/Y 0.13fF
C65844 NOR2X1_LOC_553/B INVX1_LOC_97/A 0.01fF
C65845 INVX1_LOC_1/A NAND2X1_LOC_93/B 0.18fF
C65846 NOR2X1_LOC_458/Y INVX1_LOC_96/A 0.01fF
C65847 NOR2X1_LOC_460/B NOR2X1_LOC_725/A 0.03fF
C65848 INVX1_LOC_33/A INVX1_LOC_91/A 0.19fF
C65849 NOR2X1_LOC_328/Y INVX1_LOC_146/A 0.01fF
C65850 INVX1_LOC_143/A INPUT_0 0.07fF
C65851 INVX1_LOC_1/A NAND2X1_LOC_425/Y 0.02fF
C65852 NAND2X1_LOC_354/B INVX1_LOC_264/Y 0.01fF
C65853 NAND2X1_LOC_72/Y INVX1_LOC_29/A 0.01fF
C65854 NOR2X1_LOC_38/B NAND2X1_LOC_99/A 0.00fF
C65855 NOR2X1_LOC_441/Y INVX1_LOC_9/A 0.02fF
C65856 NOR2X1_LOC_332/A INVX1_LOC_20/Y 0.02fF
C65857 INVX1_LOC_49/A INVX1_LOC_143/Y 0.04fF
C65858 NOR2X1_LOC_384/Y NOR2X1_LOC_536/A 0.48fF
C65859 NOR2X1_LOC_860/B VDD 0.12fF
C65860 INVX1_LOC_1/A NOR2X1_LOC_649/B 0.16fF
C65861 INVX1_LOC_104/A NOR2X1_LOC_405/A 0.12fF
C65862 INVX1_LOC_211/Y NOR2X1_LOC_510/B 0.43fF
C65863 NOR2X1_LOC_593/Y NOR2X1_LOC_35/Y 0.10fF
C65864 INVX1_LOC_1/A INVX1_LOC_3/A 0.15fF
C65865 NAND2X1_LOC_565/B INPUT_0 0.00fF
C65866 INVX1_LOC_62/Y NAND2X1_LOC_96/A 0.03fF
C65867 INVX1_LOC_41/A INVX1_LOC_126/A 0.03fF
C65868 INVX1_LOC_133/Y NOR2X1_LOC_139/Y 0.79fF
C65869 NOR2X1_LOC_250/A NOR2X1_LOC_841/A 0.03fF
C65870 INVX1_LOC_18/A NOR2X1_LOC_331/B 0.08fF
C65871 NOR2X1_LOC_186/Y INVX1_LOC_12/A 0.03fF
C65872 NOR2X1_LOC_78/B INVX1_LOC_186/A 0.03fF
C65873 NOR2X1_LOC_570/B INVX1_LOC_76/A 0.00fF
C65874 INVX1_LOC_276/A NAND2X1_LOC_655/A 0.95fF
C65875 NOR2X1_LOC_354/B NOR2X1_LOC_729/A 0.03fF
C65876 INVX1_LOC_14/A INVX1_LOC_63/A 3.09fF
C65877 NAND2X1_LOC_794/B NOR2X1_LOC_89/A 0.03fF
C65878 INVX1_LOC_130/A NOR2X1_LOC_155/A 0.01fF
C65879 INVX1_LOC_244/Y INVX1_LOC_38/A 0.00fF
C65880 INVX1_LOC_27/A NOR2X1_LOC_178/a_36_216# 0.01fF
C65881 NOR2X1_LOC_542/Y NOR2X1_LOC_703/A 0.00fF
C65882 NOR2X1_LOC_91/A NOR2X1_LOC_693/Y 0.03fF
C65883 INVX1_LOC_165/A INVX1_LOC_23/A 0.02fF
C65884 INVX1_LOC_40/A INVX1_LOC_91/A 1.17fF
C65885 INVX1_LOC_298/Y INVX1_LOC_50/A 0.03fF
C65886 NAND2X1_LOC_477/A INVX1_LOC_126/A 0.07fF
C65887 NOR2X1_LOC_577/Y NOR2X1_LOC_152/A 0.01fF
C65888 NOR2X1_LOC_690/A NAND2X1_LOC_721/A 0.02fF
C65889 NOR2X1_LOC_45/B INVX1_LOC_25/Y 0.14fF
C65890 NOR2X1_LOC_619/A NOR2X1_LOC_557/A 0.01fF
C65891 INPUT_0 NOR2X1_LOC_130/A 0.07fF
C65892 NOR2X1_LOC_561/Y INVX1_LOC_286/A 0.00fF
C65893 NOR2X1_LOC_78/B NAND2X1_LOC_447/Y 0.00fF
C65894 NAND2X1_LOC_601/a_36_24# NOR2X1_LOC_536/A 0.00fF
C65895 INVX1_LOC_155/A INVX1_LOC_66/Y 0.09fF
C65896 NOR2X1_LOC_590/A INVX1_LOC_84/A 0.06fF
C65897 NAND2X1_LOC_724/A INVX1_LOC_12/A 0.07fF
C65898 INVX1_LOC_50/A NOR2X1_LOC_318/a_36_216# 0.00fF
C65899 INVX1_LOC_226/Y NAND2X1_LOC_642/Y 0.01fF
C65900 NOR2X1_LOC_418/Y INVX1_LOC_187/A 0.42fF
C65901 NOR2X1_LOC_355/A NAND2X1_LOC_309/a_36_24# 0.00fF
C65902 NOR2X1_LOC_552/A INVX1_LOC_22/A 0.07fF
C65903 NAND2X1_LOC_141/A VDD -0.00fF
C65904 NOR2X1_LOC_829/Y INVX1_LOC_50/A 0.08fF
C65905 INVX1_LOC_18/A NOR2X1_LOC_592/B 0.03fF
C65906 INVX1_LOC_96/Y NOR2X1_LOC_69/a_36_216# 0.00fF
C65907 INVX1_LOC_23/A NAND2X1_LOC_288/B 0.21fF
C65908 NAND2X1_LOC_477/A NOR2X1_LOC_111/A 0.10fF
C65909 INVX1_LOC_96/Y VDD 0.69fF
C65910 NOR2X1_LOC_602/a_36_216# NOR2X1_LOC_841/A 0.12fF
C65911 INVX1_LOC_15/Y VDD 0.12fF
C65912 NOR2X1_LOC_810/A INVX1_LOC_160/A 0.02fF
C65913 NAND2X1_LOC_707/a_36_24# NOR2X1_LOC_45/B 0.00fF
C65914 INVX1_LOC_171/A NOR2X1_LOC_734/a_36_216# 0.02fF
C65915 NAND2X1_LOC_9/Y INVX1_LOC_23/Y 0.35fF
C65916 NOR2X1_LOC_187/Y INVX1_LOC_290/Y 0.03fF
C65917 NOR2X1_LOC_566/a_36_216# INVX1_LOC_22/A 0.00fF
C65918 INVX1_LOC_36/A NOR2X1_LOC_127/Y 0.01fF
C65919 INVX1_LOC_50/Y INVX1_LOC_4/Y 0.67fF
C65920 INVX1_LOC_266/Y NAND2X1_LOC_472/Y 0.10fF
C65921 INVX1_LOC_221/A NOR2X1_LOC_536/A 0.01fF
C65922 NOR2X1_LOC_142/Y INVX1_LOC_9/A 0.10fF
C65923 INVX1_LOC_83/A INVX1_LOC_186/A 0.37fF
C65924 INVX1_LOC_121/Y NOR2X1_LOC_684/Y 0.02fF
C65925 NOR2X1_LOC_111/Y INVX1_LOC_144/A 0.01fF
C65926 NOR2X1_LOC_629/B INVX1_LOC_280/A 0.01fF
C65927 INVX1_LOC_226/A VDD 0.12fF
C65928 D_INPUT_1 NOR2X1_LOC_414/Y 0.46fF
C65929 INVX1_LOC_81/A NOR2X1_LOC_155/A 0.09fF
C65930 NOR2X1_LOC_554/B NOR2X1_LOC_673/A 0.07fF
C65931 INVX1_LOC_10/A NAND2X1_LOC_642/Y 0.03fF
C65932 NOR2X1_LOC_329/B NAND2X1_LOC_858/B 0.02fF
C65933 NAND2X1_LOC_840/B VDD 0.17fF
C65934 NOR2X1_LOC_45/Y INVX1_LOC_12/A 0.05fF
C65935 INVX1_LOC_9/Y NAND2X1_LOC_211/Y 0.01fF
C65936 NOR2X1_LOC_216/Y INPUT_0 0.11fF
C65937 INVX1_LOC_286/Y INVX1_LOC_49/Y 0.01fF
C65938 NOR2X1_LOC_374/A INVX1_LOC_307/A 0.01fF
C65939 INVX1_LOC_240/A INVX1_LOC_118/A 0.03fF
C65940 INVX1_LOC_215/A INVX1_LOC_76/A 0.10fF
C65941 NAND2X1_LOC_580/a_36_24# INVX1_LOC_42/A 0.00fF
C65942 NOR2X1_LOC_100/A INVX1_LOC_230/A 0.03fF
C65943 NOR2X1_LOC_447/a_36_216# NOR2X1_LOC_447/B 0.00fF
C65944 NOR2X1_LOC_656/a_36_216# INVX1_LOC_63/A 0.00fF
C65945 INVX1_LOC_30/Y NAND2X1_LOC_267/B 0.02fF
C65946 NOR2X1_LOC_690/A NOR2X1_LOC_823/a_36_216# 0.01fF
C65947 INVX1_LOC_22/A INVX1_LOC_139/Y 0.03fF
C65948 INVX1_LOC_266/A INVX1_LOC_4/Y 0.10fF
C65949 NAND2X1_LOC_364/Y NAND2X1_LOC_412/a_36_24# 0.00fF
C65950 NOR2X1_LOC_352/Y INVX1_LOC_38/A 0.04fF
C65951 NAND2X1_LOC_374/Y INVX1_LOC_38/A 0.07fF
C65952 INVX1_LOC_266/Y NAND2X1_LOC_637/Y 0.04fF
C65953 INVX1_LOC_72/Y NAND2X1_LOC_773/B 0.02fF
C65954 NOR2X1_LOC_178/Y NAND2X1_LOC_205/A 0.02fF
C65955 NOR2X1_LOC_346/B INVX1_LOC_280/A 0.02fF
C65956 NOR2X1_LOC_558/a_36_216# INVX1_LOC_22/A 0.00fF
C65957 NOR2X1_LOC_655/B INVX1_LOC_9/A 0.13fF
C65958 INVX1_LOC_1/A NAND2X1_LOC_470/B 0.06fF
C65959 NAND2X1_LOC_354/B NOR2X1_LOC_88/Y 0.46fF
C65960 NAND2X1_LOC_84/Y INVX1_LOC_63/A 1.66fF
C65961 INVX1_LOC_53/A NAND2X1_LOC_431/a_36_24# 0.00fF
C65962 NAND2X1_LOC_777/a_36_24# NOR2X1_LOC_109/Y 0.01fF
C65963 INVX1_LOC_10/Y INVX1_LOC_22/A 0.03fF
C65964 NAND2X1_LOC_1/a_36_24# NAND2X1_LOC_1/Y 0.01fF
C65965 NOR2X1_LOC_288/A NOR2X1_LOC_445/B 0.03fF
C65966 INVX1_LOC_49/A NOR2X1_LOC_631/A 0.30fF
C65967 NOR2X1_LOC_590/A INVX1_LOC_15/A 0.31fF
C65968 INVX1_LOC_75/A NOR2X1_LOC_45/B 0.16fF
C65969 INVX1_LOC_161/Y NOR2X1_LOC_334/Y 1.54fF
C65970 INVX1_LOC_286/A NOR2X1_LOC_167/Y 0.02fF
C65971 NOR2X1_LOC_576/B VDD 1.68fF
C65972 INVX1_LOC_311/A NOR2X1_LOC_741/A 0.03fF
C65973 NAND2X1_LOC_354/B INVX1_LOC_84/A 0.03fF
C65974 INVX1_LOC_88/A NAND2X1_LOC_61/Y 0.02fF
C65975 NAND2X1_LOC_794/B NAND2X1_LOC_804/A 0.03fF
C65976 NOR2X1_LOC_553/B INVX1_LOC_38/A 0.03fF
C65977 NAND2X1_LOC_569/A NAND2X1_LOC_489/Y 0.02fF
C65978 INVX1_LOC_105/A INVX1_LOC_29/A 0.07fF
C65979 NOR2X1_LOC_848/Y NOR2X1_LOC_843/B 0.04fF
C65980 INVX1_LOC_75/A INVX1_LOC_247/A 0.03fF
C65981 NAND2X1_LOC_337/B NOR2X1_LOC_301/A 0.01fF
C65982 NAND2X1_LOC_76/a_36_24# INVX1_LOC_78/A 0.00fF
C65983 INVX1_LOC_72/A INVX1_LOC_47/Y 0.10fF
C65984 NOR2X1_LOC_433/A INVX1_LOC_109/A 0.00fF
C65985 NAND2X1_LOC_834/a_36_24# INVX1_LOC_92/A 0.00fF
C65986 NOR2X1_LOC_148/B NOR2X1_LOC_148/Y 0.00fF
C65987 NOR2X1_LOC_561/Y INVX1_LOC_54/A 0.32fF
C65988 INVX1_LOC_30/A NAND2X1_LOC_471/Y 0.02fF
C65989 NOR2X1_LOC_481/A INVX1_LOC_12/A 0.03fF
C65990 INVX1_LOC_35/A INVX1_LOC_59/A 0.04fF
C65991 NOR2X1_LOC_488/Y NOR2X1_LOC_88/Y 0.03fF
C65992 NOR2X1_LOC_99/B INVX1_LOC_9/A 0.09fF
C65993 INVX1_LOC_77/A NOR2X1_LOC_850/B 0.05fF
C65994 INVX1_LOC_35/A NAND2X1_LOC_773/Y 0.03fF
C65995 INVX1_LOC_31/A NOR2X1_LOC_693/Y 0.07fF
C65996 INVX1_LOC_174/A NAND2X1_LOC_64/a_36_24# -0.02fF
C65997 INVX1_LOC_151/A INVX1_LOC_109/A 0.06fF
C65998 INVX1_LOC_225/A INVX1_LOC_12/A 0.07fF
C65999 INVX1_LOC_25/A INVX1_LOC_256/A 0.39fF
C66000 NOR2X1_LOC_846/B INVX1_LOC_9/A 0.01fF
C66001 NAND2X1_LOC_656/A NOR2X1_LOC_38/B 0.03fF
C66002 NOR2X1_LOC_589/a_36_216# INVX1_LOC_37/A 0.00fF
C66003 NOR2X1_LOC_382/Y INVX1_LOC_26/A 0.09fF
C66004 NOR2X1_LOC_75/Y NOR2X1_LOC_604/a_36_216# 0.00fF
C66005 NOR2X1_LOC_488/Y INVX1_LOC_84/A 0.01fF
C66006 NOR2X1_LOC_649/Y NAND2X1_LOC_473/A 0.07fF
C66007 NOR2X1_LOC_340/Y NOR2X1_LOC_861/Y 0.11fF
C66008 INVX1_LOC_135/A NOR2X1_LOC_88/A 0.02fF
C66009 INVX1_LOC_286/A INVX1_LOC_76/A 0.07fF
C66010 INVX1_LOC_42/Y NAND2X1_LOC_472/Y 0.03fF
C66011 NAND2X1_LOC_347/B INVX1_LOC_306/Y 0.02fF
C66012 NAND2X1_LOC_793/Y NAND2X1_LOC_793/B 0.02fF
C66013 INVX1_LOC_75/A INVX1_LOC_281/A 0.10fF
C66014 INVX1_LOC_136/A NOR2X1_LOC_318/A 0.00fF
C66015 NOR2X1_LOC_733/Y VDD 0.16fF
C66016 INVX1_LOC_182/A INVX1_LOC_9/A 0.07fF
C66017 INVX1_LOC_218/A INVX1_LOC_19/A 0.03fF
C66018 INVX1_LOC_36/A NOR2X1_LOC_383/B 5.93fF
C66019 INVX1_LOC_17/A NAND2X1_LOC_552/A 0.03fF
C66020 NOR2X1_LOC_456/Y INVX1_LOC_188/A 0.18fF
C66021 NAND2X1_LOC_479/Y NAND2X1_LOC_476/Y 0.00fF
C66022 INVX1_LOC_25/A NOR2X1_LOC_606/Y 0.05fF
C66023 INVX1_LOC_17/A INVX1_LOC_5/A 7.03fF
C66024 NOR2X1_LOC_276/Y NOR2X1_LOC_678/A 0.10fF
C66025 INVX1_LOC_72/A NOR2X1_LOC_651/a_36_216# 0.00fF
C66026 INVX1_LOC_30/A NAND2X1_LOC_201/a_36_24# 0.00fF
C66027 NOR2X1_LOC_264/Y INVX1_LOC_32/A 0.06fF
C66028 INVX1_LOC_92/Y INVX1_LOC_117/A 0.03fF
C66029 D_INPUT_1 INVX1_LOC_40/Y 0.00fF
C66030 INVX1_LOC_51/Y NAND2X1_LOC_96/A 0.01fF
C66031 NAND2X1_LOC_479/Y INVX1_LOC_186/Y 0.07fF
C66032 NAND2X1_LOC_738/B INVX1_LOC_36/A 0.03fF
C66033 INVX1_LOC_227/A INVX1_LOC_84/A 0.07fF
C66034 NOR2X1_LOC_45/B NAND2X1_LOC_453/A 0.07fF
C66035 NOR2X1_LOC_528/Y INVX1_LOC_37/A 0.03fF
C66036 NOR2X1_LOC_703/B NOR2X1_LOC_748/A 0.01fF
C66037 INVX1_LOC_64/A NOR2X1_LOC_644/B 0.02fF
C66038 NOR2X1_LOC_471/Y INVX1_LOC_5/A 0.02fF
C66039 NOR2X1_LOC_637/B NAND2X1_LOC_175/Y 0.00fF
C66040 INVX1_LOC_11/A NAND2X1_LOC_794/B 0.01fF
C66041 INVX1_LOC_95/A INVX1_LOC_76/A 0.03fF
C66042 INVX1_LOC_243/A NOR2X1_LOC_48/B 0.01fF
C66043 NOR2X1_LOC_300/a_36_216# NAND2X1_LOC_212/Y 0.03fF
C66044 INPUT_0 NOR2X1_LOC_16/a_36_216# 0.00fF
C66045 INVX1_LOC_6/A NAND2X1_LOC_476/a_36_24# 0.00fF
C66046 NAND2X1_LOC_555/Y INVX1_LOC_5/A 0.06fF
C66047 NAND2X1_LOC_198/B INVX1_LOC_271/A 0.07fF
C66048 INVX1_LOC_201/Y INVX1_LOC_90/Y 0.07fF
C66049 NOR2X1_LOC_6/B INVX1_LOC_4/Y 0.23fF
C66050 NOR2X1_LOC_208/Y NOR2X1_LOC_383/B 0.07fF
C66051 INVX1_LOC_21/A NAND2X1_LOC_550/A 0.07fF
C66052 INVX1_LOC_88/Y NAND2X1_LOC_454/Y 0.01fF
C66053 NOR2X1_LOC_15/Y NOR2X1_LOC_361/B 0.07fF
C66054 INVX1_LOC_136/A NOR2X1_LOC_678/A 0.03fF
C66055 NOR2X1_LOC_419/Y NOR2X1_LOC_720/A 0.00fF
C66056 NOR2X1_LOC_527/Y INVX1_LOC_185/A 0.01fF
C66057 NOR2X1_LOC_167/Y INVX1_LOC_54/A 0.03fF
C66058 INVX1_LOC_11/A INVX1_LOC_48/Y 0.07fF
C66059 INVX1_LOC_290/A NOR2X1_LOC_89/A 0.00fF
C66060 NAND2X1_LOC_447/Y INVX1_LOC_46/A 0.54fF
C66061 INVX1_LOC_45/Y INVX1_LOC_23/A 0.01fF
C66062 NOR2X1_LOC_246/A NOR2X1_LOC_662/A 0.01fF
C66063 INVX1_LOC_21/A NOR2X1_LOC_160/B 1.99fF
C66064 INVX1_LOC_94/A INVX1_LOC_29/Y 0.07fF
C66065 D_INPUT_3 INVX1_LOC_59/Y 1.33fF
C66066 INVX1_LOC_16/A NAND2X1_LOC_254/Y 0.17fF
C66067 INVX1_LOC_57/Y NOR2X1_LOC_109/Y 0.09fF
C66068 INVX1_LOC_13/Y NAND2X1_LOC_768/a_36_24# 0.01fF
C66069 NAND2X1_LOC_593/Y NOR2X1_LOC_654/A 0.03fF
C66070 INVX1_LOC_36/A NAND2X1_LOC_29/a_36_24# 0.00fF
C66071 NOR2X1_LOC_763/Y NAND2X1_LOC_651/B 0.05fF
C66072 NAND2X1_LOC_190/Y NAND2X1_LOC_192/B 0.18fF
C66073 NOR2X1_LOC_188/A NAND2X1_LOC_93/B 1.18fF
C66074 NOR2X1_LOC_130/A NOR2X1_LOC_84/B 0.05fF
C66075 NOR2X1_LOC_807/B INVX1_LOC_1/A 0.15fF
C66076 INVX1_LOC_255/Y NOR2X1_LOC_847/a_36_216# 0.01fF
C66077 INVX1_LOC_243/A NAND2X1_LOC_3/B 0.06fF
C66078 INVX1_LOC_256/A INVX1_LOC_1/A 0.07fF
C66079 NOR2X1_LOC_804/B NOR2X1_LOC_383/B 0.01fF
C66080 INVX1_LOC_316/Y INVX1_LOC_32/A 1.39fF
C66081 INVX1_LOC_120/A NAND2X1_LOC_63/Y 0.00fF
C66082 NOR2X1_LOC_413/Y NOR2X1_LOC_19/a_36_216# 0.01fF
C66083 NOR2X1_LOC_667/Y NAND2X1_LOC_326/A 0.00fF
C66084 NOR2X1_LOC_189/A NAND2X1_LOC_804/A 0.02fF
C66085 NOR2X1_LOC_716/B INVX1_LOC_129/A 0.01fF
C66086 INVX1_LOC_6/A INVX1_LOC_179/A 0.00fF
C66087 NOR2X1_LOC_561/Y NOR2X1_LOC_48/B 0.10fF
C66088 INVX1_LOC_90/A INVX1_LOC_125/A 0.34fF
C66089 INVX1_LOC_50/A INVX1_LOC_8/A 0.06fF
C66090 INVX1_LOC_10/A NAND2X1_LOC_792/B 0.04fF
C66091 NOR2X1_LOC_309/Y NOR2X1_LOC_383/B 0.03fF
C66092 INVX1_LOC_17/A NOR2X1_LOC_816/A 0.12fF
C66093 NAND2X1_LOC_724/A NAND2X1_LOC_733/Y 0.10fF
C66094 NOR2X1_LOC_92/Y NOR2X1_LOC_761/Y 0.08fF
C66095 NOR2X1_LOC_264/Y NOR2X1_LOC_622/A 0.00fF
C66096 NOR2X1_LOC_99/B NOR2X1_LOC_861/Y 0.02fF
C66097 NOR2X1_LOC_78/A INVX1_LOC_92/A 0.02fF
C66098 NOR2X1_LOC_773/Y NOR2X1_LOC_301/A 0.18fF
C66099 NOR2X1_LOC_210/B INVX1_LOC_78/A 0.10fF
C66100 INVX1_LOC_176/A INVX1_LOC_230/A 0.03fF
C66101 NOR2X1_LOC_135/Y INVX1_LOC_272/A 0.01fF
C66102 INVX1_LOC_30/Y INVX1_LOC_4/Y 0.06fF
C66103 NOR2X1_LOC_763/Y INVX1_LOC_15/A 0.17fF
C66104 NOR2X1_LOC_420/a_36_216# INVX1_LOC_77/A 0.02fF
C66105 NAND2X1_LOC_9/Y NAND2X1_LOC_116/A 0.07fF
C66106 NOR2X1_LOC_419/Y NOR2X1_LOC_849/A 0.04fF
C66107 NOR2X1_LOC_68/A NAND2X1_LOC_780/Y 0.02fF
C66108 INVX1_LOC_24/Y NAND2X1_LOC_364/A 0.10fF
C66109 INVX1_LOC_28/A NAND2X1_LOC_254/Y 0.02fF
C66110 INVX1_LOC_76/A INVX1_LOC_54/A 0.41fF
C66111 NOR2X1_LOC_226/A NOR2X1_LOC_677/Y 0.04fF
C66112 INVX1_LOC_22/A NOR2X1_LOC_541/B 0.01fF
C66113 NOR2X1_LOC_598/B NOR2X1_LOC_802/A 0.12fF
C66114 INVX1_LOC_48/A INVX1_LOC_63/A 0.03fF
C66115 INVX1_LOC_13/A NOR2X1_LOC_55/a_36_216# 0.00fF
C66116 INVX1_LOC_286/Y INVX1_LOC_161/A 0.07fF
C66117 NAND2X1_LOC_860/A INVX1_LOC_256/Y 0.04fF
C66118 NAND2X1_LOC_859/Y NOR2X1_LOC_693/Y 0.07fF
C66119 NOR2X1_LOC_272/Y INVX1_LOC_41/A 0.03fF
C66120 NAND2X1_LOC_850/A INVX1_LOC_32/A 0.03fF
C66121 NOR2X1_LOC_716/B NOR2X1_LOC_440/B 0.02fF
C66122 NOR2X1_LOC_719/A NAND2X1_LOC_215/A 0.21fF
C66123 NOR2X1_LOC_68/A NAND2X1_LOC_114/B 0.23fF
C66124 INVX1_LOC_13/A INVX1_LOC_57/A 0.03fF
C66125 INVX1_LOC_255/Y INVX1_LOC_23/A 0.22fF
C66126 INVX1_LOC_224/A NOR2X1_LOC_350/A 0.02fF
C66127 NOR2X1_LOC_665/A INVX1_LOC_271/A 0.16fF
C66128 NAND2X1_LOC_35/B NOR2X1_LOC_411/Y 0.32fF
C66129 INVX1_LOC_278/A NOR2X1_LOC_488/Y 0.04fF
C66130 INVX1_LOC_24/A INVX1_LOC_225/Y 0.05fF
C66131 NAND2X1_LOC_9/Y INVX1_LOC_232/A 0.07fF
C66132 INVX1_LOC_71/A NAND2X1_LOC_793/Y 0.75fF
C66133 INVX1_LOC_135/A NOR2X1_LOC_843/B 0.03fF
C66134 NOR2X1_LOC_458/Y NOR2X1_LOC_15/Y 0.04fF
C66135 NOR2X1_LOC_167/Y NOR2X1_LOC_48/B 0.12fF
C66136 NOR2X1_LOC_15/Y INVX1_LOC_153/Y 0.10fF
C66137 NOR2X1_LOC_91/A NOR2X1_LOC_71/Y 0.07fF
C66138 INVX1_LOC_278/A NOR2X1_LOC_82/Y 0.05fF
C66139 NOR2X1_LOC_590/A NOR2X1_LOC_168/Y 0.06fF
C66140 INVX1_LOC_294/Y NAND2X1_LOC_347/B 0.01fF
C66141 INVX1_LOC_11/A NOR2X1_LOC_350/A 0.03fF
C66142 NAND2X1_LOC_112/Y INVX1_LOC_53/A 0.01fF
C66143 INVX1_LOC_7/A NAND2X1_LOC_215/A 1.10fF
C66144 NAND2X1_LOC_67/Y NOR2X1_LOC_142/Y 0.22fF
C66145 NAND2X1_LOC_342/Y NOR2X1_LOC_652/Y 0.03fF
C66146 NOR2X1_LOC_272/Y NOR2X1_LOC_398/Y 0.05fF
C66147 NAND2X1_LOC_866/B NOR2X1_LOC_693/Y 0.02fF
C66148 NAND2X1_LOC_199/B NAND2X1_LOC_199/a_36_24# 0.00fF
C66149 NOR2X1_LOC_489/B INVX1_LOC_1/Y 0.01fF
C66150 NOR2X1_LOC_99/Y NAND2X1_LOC_297/a_36_24# 0.01fF
C66151 NOR2X1_LOC_256/a_36_216# INVX1_LOC_61/Y 0.00fF
C66152 NOR2X1_LOC_88/A INVX1_LOC_280/A 0.01fF
C66153 NOR2X1_LOC_68/A INVX1_LOC_312/Y 0.07fF
C66154 NOR2X1_LOC_15/Y INVX1_LOC_121/Y 0.48fF
C66155 INVX1_LOC_140/A NOR2X1_LOC_30/Y 0.05fF
C66156 INVX1_LOC_50/A NAND2X1_LOC_140/A 0.03fF
C66157 INVX1_LOC_200/A NAND2X1_LOC_640/Y 0.01fF
C66158 NOR2X1_LOC_294/Y NOR2X1_LOC_68/A 0.00fF
C66159 NOR2X1_LOC_124/A NAND2X1_LOC_81/B 0.06fF
C66160 NOR2X1_LOC_560/A NOR2X1_LOC_843/B 0.05fF
C66161 INVX1_LOC_246/A NOR2X1_LOC_433/A 0.00fF
C66162 VDD NAND2X1_LOC_456/Y 0.02fF
C66163 NOR2X1_LOC_246/A INVX1_LOC_57/A 0.15fF
C66164 INVX1_LOC_233/A NOR2X1_LOC_383/Y 0.22fF
C66165 INVX1_LOC_12/A NAND2X1_LOC_642/Y 0.10fF
C66166 INVX1_LOC_85/Y NOR2X1_LOC_727/B 0.02fF
C66167 INVX1_LOC_45/A NOR2X1_LOC_607/A 0.09fF
C66168 NAND2X1_LOC_553/A INVX1_LOC_232/A 0.01fF
C66169 INVX1_LOC_36/A NOR2X1_LOC_512/Y 0.01fF
C66170 INVX1_LOC_140/A NOR2X1_LOC_301/A 0.03fF
C66171 NOR2X1_LOC_71/Y INVX1_LOC_23/A 0.08fF
C66172 INVX1_LOC_35/A INVX1_LOC_279/A 0.07fF
C66173 NOR2X1_LOC_453/Y INVX1_LOC_189/A 0.00fF
C66174 NOR2X1_LOC_15/Y INVX1_LOC_177/A 0.03fF
C66175 NOR2X1_LOC_649/a_36_216# INPUT_3 0.01fF
C66176 INVX1_LOC_299/A NOR2X1_LOC_175/A 0.70fF
C66177 INVX1_LOC_33/Y INVX1_LOC_119/Y 0.02fF
C66178 INVX1_LOC_21/A INVX1_LOC_208/A 0.37fF
C66179 INVX1_LOC_239/A INVX1_LOC_197/A 0.12fF
C66180 NOR2X1_LOC_798/A INVX1_LOC_232/A 0.02fF
C66181 INVX1_LOC_27/A NOR2X1_LOC_219/Y 0.70fF
C66182 INVX1_LOC_139/Y INVX1_LOC_186/Y 0.01fF
C66183 NOR2X1_LOC_506/Y NAND2X1_LOC_798/B 0.21fF
C66184 INVX1_LOC_88/A INVX1_LOC_133/Y 0.12fF
C66185 INVX1_LOC_21/A NOR2X1_LOC_516/B 0.03fF
C66186 VDD INVX1_LOC_49/Y 0.08fF
C66187 NOR2X1_LOC_538/B NOR2X1_LOC_175/A 0.02fF
C66188 INVX1_LOC_27/A INVX1_LOC_53/Y 0.08fF
C66189 NOR2X1_LOC_644/A INVX1_LOC_23/A 0.03fF
C66190 INVX1_LOC_284/Y INVX1_LOC_207/A 0.03fF
C66191 INVX1_LOC_276/A INVX1_LOC_88/A 0.07fF
C66192 INVX1_LOC_11/A NOR2X1_LOC_84/Y 0.07fF
C66193 INVX1_LOC_24/A INVX1_LOC_72/Y 0.29fF
C66194 NOR2X1_LOC_254/a_36_216# NOR2X1_LOC_254/Y 0.01fF
C66195 INVX1_LOC_52/Y INVX1_LOC_52/A -0.01fF
C66196 NOR2X1_LOC_471/Y NOR2X1_LOC_377/Y 0.00fF
C66197 INVX1_LOC_2/A NOR2X1_LOC_533/Y 0.05fF
C66198 INVX1_LOC_57/Y NOR2X1_LOC_237/Y 0.73fF
C66199 NAND2X1_LOC_800/A INVX1_LOC_49/Y 0.03fF
C66200 INVX1_LOC_5/A NOR2X1_LOC_199/B 0.04fF
C66201 NOR2X1_LOC_358/a_36_216# NOR2X1_LOC_155/A 0.00fF
C66202 INVX1_LOC_61/Y INVX1_LOC_8/A 0.08fF
C66203 NAND2X1_LOC_807/B INVX1_LOC_76/A 0.36fF
C66204 NAND2X1_LOC_741/B NAND2X1_LOC_812/A 0.01fF
C66205 NAND2X1_LOC_254/Y NOR2X1_LOC_253/Y 0.03fF
C66206 INVX1_LOC_62/Y NAND2X1_LOC_656/A 0.09fF
C66207 INVX1_LOC_34/A INVX1_LOC_286/Y 0.18fF
C66208 NOR2X1_LOC_690/A NAND2X1_LOC_500/Y 0.03fF
C66209 INVX1_LOC_13/A INVX1_LOC_252/A 0.01fF
C66210 NAND2X1_LOC_472/Y INVX1_LOC_19/A 0.07fF
C66211 NOR2X1_LOC_828/B INVX1_LOC_23/A 0.40fF
C66212 INVX1_LOC_246/Y INVX1_LOC_24/A 0.01fF
C66213 NOR2X1_LOC_722/Y INVX1_LOC_283/Y 0.31fF
C66214 VDD INVX1_LOC_99/A 0.04fF
C66215 NOR2X1_LOC_607/A INVX1_LOC_71/A 0.01fF
C66216 INVX1_LOC_224/A NAND2X1_LOC_292/a_36_24# 0.00fF
C66217 NOR2X1_LOC_48/B INVX1_LOC_76/A 0.14fF
C66218 INVX1_LOC_17/A NOR2X1_LOC_773/Y 0.07fF
C66219 NAND2X1_LOC_9/Y NOR2X1_LOC_775/Y 0.01fF
C66220 NOR2X1_LOC_186/Y NAND2X1_LOC_808/A 0.09fF
C66221 NOR2X1_LOC_593/Y NAND2X1_LOC_272/a_36_24# 0.01fF
C66222 INVX1_LOC_58/A NOR2X1_LOC_322/Y 0.51fF
C66223 NOR2X1_LOC_68/A INVX1_LOC_275/A 0.02fF
C66224 INVX1_LOC_6/A NOR2X1_LOC_693/Y 0.25fF
C66225 NOR2X1_LOC_92/Y NOR2X1_LOC_86/A 0.06fF
C66226 NAND2X1_LOC_124/a_36_24# INVX1_LOC_271/A 0.00fF
C66227 NAND2X1_LOC_802/A INVX1_LOC_24/A 0.49fF
C66228 INVX1_LOC_14/A INVX1_LOC_1/Y 0.30fF
C66229 NOR2X1_LOC_92/Y NAND2X1_LOC_632/a_36_24# 0.01fF
C66230 INVX1_LOC_41/A NAND2X1_LOC_364/A 0.07fF
C66231 NOR2X1_LOC_48/B NAND2X1_LOC_405/a_36_24# 0.01fF
C66232 INVX1_LOC_57/Y NOR2X1_LOC_309/Y 0.10fF
C66233 INVX1_LOC_38/A INVX1_LOC_125/A 0.03fF
C66234 INVX1_LOC_287/A NOR2X1_LOC_711/A 0.05fF
C66235 NOR2X1_LOC_440/Y INVX1_LOC_1/A 0.27fF
C66236 INVX1_LOC_90/A NOR2X1_LOC_81/Y 0.07fF
C66237 NOR2X1_LOC_716/B INVX1_LOC_41/Y 0.00fF
C66238 NOR2X1_LOC_810/A INVX1_LOC_1/A 0.03fF
C66239 INVX1_LOC_34/A INVX1_LOC_159/A 0.11fF
C66240 NOR2X1_LOC_246/Y NOR2X1_LOC_652/Y 0.03fF
C66241 NAND2X1_LOC_573/Y NAND2X1_LOC_808/A 0.00fF
C66242 NOR2X1_LOC_15/Y NAND2X1_LOC_573/A 0.10fF
C66243 NAND2X1_LOC_650/B INVX1_LOC_15/A 0.07fF
C66244 NAND2X1_LOC_637/Y INVX1_LOC_19/A 0.03fF
C66245 INVX1_LOC_87/Y NOR2X1_LOC_652/Y 0.01fF
C66246 INVX1_LOC_11/A INVX1_LOC_290/A 0.07fF
C66247 INVX1_LOC_12/A NOR2X1_LOC_271/Y 0.01fF
C66248 NAND2X1_LOC_538/Y NOR2X1_LOC_512/a_36_216# 0.01fF
C66249 NAND2X1_LOC_733/Y NAND2X1_LOC_852/Y 0.10fF
C66250 INPUT_3 INVX1_LOC_316/Y 0.04fF
C66251 NOR2X1_LOC_42/a_36_216# NOR2X1_LOC_38/B 0.00fF
C66252 NAND2X1_LOC_724/A NAND2X1_LOC_808/A 0.14fF
C66253 NOR2X1_LOC_816/a_36_216# INVX1_LOC_28/A 0.02fF
C66254 NOR2X1_LOC_764/Y INVX1_LOC_1/A 0.01fF
C66255 NOR2X1_LOC_68/A NOR2X1_LOC_168/B 0.03fF
C66256 INVX1_LOC_27/A NAND2X1_LOC_506/a_36_24# 0.00fF
C66257 NOR2X1_LOC_295/a_36_216# INVX1_LOC_77/A 0.01fF
C66258 INVX1_LOC_91/A NOR2X1_LOC_748/A 0.17fF
C66259 INVX1_LOC_126/Y NOR2X1_LOC_129/a_36_216# 0.00fF
C66260 INVX1_LOC_17/A NOR2X1_LOC_332/A 0.15fF
C66261 NAND2X1_LOC_501/a_36_24# NAND2X1_LOC_374/Y 0.00fF
C66262 INVX1_LOC_255/Y INVX1_LOC_31/A 0.12fF
C66263 NAND2X1_LOC_350/A NOR2X1_LOC_561/Y 0.03fF
C66264 INVX1_LOC_136/A NOR2X1_LOC_191/A 0.04fF
C66265 NOR2X1_LOC_596/A NOR2X1_LOC_423/Y 0.02fF
C66266 INVX1_LOC_24/A INVX1_LOC_266/Y 0.03fF
C66267 NOR2X1_LOC_721/B NAND2X1_LOC_85/Y 0.15fF
C66268 INVX1_LOC_2/A NOR2X1_LOC_735/a_36_216# 0.00fF
C66269 NAND2X1_LOC_231/Y INVX1_LOC_159/A 0.02fF
C66270 NOR2X1_LOC_391/A INVX1_LOC_43/Y 0.12fF
C66271 INVX1_LOC_21/A NOR2X1_LOC_706/A 1.68fF
C66272 NAND2X1_LOC_341/A INVX1_LOC_30/A 0.22fF
C66273 INVX1_LOC_217/A NAND2X1_LOC_852/Y 0.10fF
C66274 INVX1_LOC_90/A NAND2X1_LOC_538/Y 0.07fF
C66275 NOR2X1_LOC_259/a_36_216# INVX1_LOC_89/A 0.00fF
C66276 NOR2X1_LOC_78/A INVX1_LOC_53/A 1.12fF
C66277 NOR2X1_LOC_808/A NOR2X1_LOC_500/A 0.03fF
C66278 NOR2X1_LOC_328/Y INVX1_LOC_72/A 0.05fF
C66279 NOR2X1_LOC_222/Y NOR2X1_LOC_596/A 0.03fF
C66280 NAND2X1_LOC_195/a_36_24# INVX1_LOC_159/A 0.00fF
C66281 NOR2X1_LOC_445/Y INVX1_LOC_104/A 0.02fF
C66282 NOR2X1_LOC_251/Y NAND2X1_LOC_198/B 0.14fF
C66283 NOR2X1_LOC_662/A NAND2X1_LOC_489/Y 0.10fF
C66284 NOR2X1_LOC_273/Y NAND2X1_LOC_841/A 0.06fF
C66285 NAND2X1_LOC_792/B INVX1_LOC_307/A 0.05fF
C66286 INVX1_LOC_18/A NAND2X1_LOC_479/Y 0.07fF
C66287 NAND2X1_LOC_139/A INVX1_LOC_80/Y 0.03fF
C66288 NAND2X1_LOC_348/A NOR2X1_LOC_140/A 0.11fF
C66289 INVX1_LOC_90/A NOR2X1_LOC_530/Y 0.24fF
C66290 INVX1_LOC_31/A NOR2X1_LOC_71/Y 0.03fF
C66291 INVX1_LOC_19/A NAND2X1_LOC_206/Y 0.07fF
C66292 NAND2X1_LOC_581/Y NOR2X1_LOC_635/A 0.11fF
C66293 NOR2X1_LOC_68/A NOR2X1_LOC_789/A 0.03fF
C66294 INVX1_LOC_45/A NOR2X1_LOC_686/B 0.02fF
C66295 NOR2X1_LOC_6/B INVX1_LOC_82/A 0.06fF
C66296 NOR2X1_LOC_295/a_36_216# INVX1_LOC_124/A 0.01fF
C66297 NAND2X1_LOC_352/B NOR2X1_LOC_389/a_36_216# 0.00fF
C66298 NAND2X1_LOC_347/B NOR2X1_LOC_74/A 0.00fF
C66299 INVX1_LOC_17/A INVX1_LOC_140/A 0.07fF
C66300 NOR2X1_LOC_489/B INVX1_LOC_93/Y 0.02fF
C66301 INVX1_LOC_153/Y INVX1_LOC_96/Y 0.10fF
C66302 INVX1_LOC_19/A NAND2X1_LOC_773/B 0.03fF
C66303 NOR2X1_LOC_392/B NOR2X1_LOC_709/A 0.10fF
C66304 NOR2X1_LOC_798/A INVX1_LOC_186/A 0.06fF
C66305 INVX1_LOC_102/Y NAND2X1_LOC_793/Y 0.07fF
C66306 NOR2X1_LOC_717/B INVX1_LOC_142/A 0.00fF
C66307 NAND2X1_LOC_84/Y INVX1_LOC_1/Y 0.03fF
C66308 INVX1_LOC_314/Y INVX1_LOC_16/A 0.07fF
C66309 INVX1_LOC_21/A INVX1_LOC_315/Y 0.02fF
C66310 INVX1_LOC_1/A NOR2X1_LOC_710/a_36_216# 0.00fF
C66311 INVX1_LOC_208/Y INVX1_LOC_77/A 0.01fF
C66312 INVX1_LOC_94/A INVX1_LOC_101/A 0.01fF
C66313 NAND2X1_LOC_866/A GATE_865 0.10fF
C66314 NOR2X1_LOC_86/A NAND2X1_LOC_837/Y 0.10fF
C66315 NOR2X1_LOC_210/B INVX1_LOC_113/Y 0.00fF
C66316 NOR2X1_LOC_389/A NOR2X1_LOC_329/B 0.10fF
C66317 NOR2X1_LOC_598/B INVX1_LOC_2/Y 0.03fF
C66318 INVX1_LOC_11/Y NOR2X1_LOC_304/Y 0.02fF
C66319 INVX1_LOC_135/A INVX1_LOC_18/A 0.16fF
C66320 NOR2X1_LOC_698/Y NOR2X1_LOC_748/A 0.03fF
C66321 INVX1_LOC_249/A NOR2X1_LOC_665/A 0.04fF
C66322 NAND2X1_LOC_276/Y INVX1_LOC_40/A 0.05fF
C66323 INVX1_LOC_63/Y INVX1_LOC_52/A 0.04fF
C66324 NOR2X1_LOC_843/B INVX1_LOC_280/A 0.07fF
C66325 INVX1_LOC_89/A NOR2X1_LOC_703/B 0.03fF
C66326 NOR2X1_LOC_363/Y NOR2X1_LOC_125/Y 0.10fF
C66327 INVX1_LOC_290/A NOR2X1_LOC_433/A 0.02fF
C66328 NOR2X1_LOC_15/Y NOR2X1_LOC_183/a_36_216# 0.00fF
C66329 NOR2X1_LOC_602/a_36_216# INVX1_LOC_90/A 0.00fF
C66330 INVX1_LOC_225/A NOR2X1_LOC_566/Y 0.02fF
C66331 INVX1_LOC_12/A NOR2X1_LOC_48/Y 0.01fF
C66332 INVX1_LOC_256/A NOR2X1_LOC_188/A 0.19fF
C66333 INVX1_LOC_24/A NAND2X1_LOC_862/a_36_24# 0.01fF
C66334 INVX1_LOC_45/A INVX1_LOC_148/A 0.01fF
C66335 NOR2X1_LOC_551/B NOR2X1_LOC_687/Y 0.12fF
C66336 NOR2X1_LOC_554/B INVX1_LOC_20/Y 0.02fF
C66337 NOR2X1_LOC_355/A INVX1_LOC_94/A 0.10fF
C66338 NOR2X1_LOC_409/B NAND2X1_LOC_802/Y 0.01fF
C66339 NOR2X1_LOC_798/A NAND2X1_LOC_447/Y 0.03fF
C66340 NOR2X1_LOC_53/Y NAND2X1_LOC_453/A 0.01fF
C66341 INVX1_LOC_58/A INVX1_LOC_281/Y 0.00fF
C66342 INVX1_LOC_256/A NOR2X1_LOC_548/B 0.10fF
C66343 NOR2X1_LOC_590/A NOR2X1_LOC_310/a_36_216# 0.00fF
C66344 NOR2X1_LOC_644/Y NOR2X1_LOC_78/B 0.01fF
C66345 NAND2X1_LOC_564/B NAND2X1_LOC_569/A 0.03fF
C66346 NOR2X1_LOC_68/A NAND2X1_LOC_638/Y 0.01fF
C66347 INVX1_LOC_50/A INVX1_LOC_118/Y 0.03fF
C66348 NOR2X1_LOC_751/A INVX1_LOC_31/A 0.08fF
C66349 NOR2X1_LOC_92/Y NOR2X1_LOC_405/A 3.83fF
C66350 NOR2X1_LOC_160/B INVX1_LOC_311/A 0.06fF
C66351 NOR2X1_LOC_742/A NOR2X1_LOC_717/Y 0.01fF
C66352 INVX1_LOC_99/Y INVX1_LOC_37/A 0.10fF
C66353 INVX1_LOC_213/Y NOR2X1_LOC_687/Y 2.09fF
C66354 NOR2X1_LOC_411/Y VDD 0.02fF
C66355 NOR2X1_LOC_490/Y INVX1_LOC_18/A 0.04fF
C66356 INVX1_LOC_172/A INVX1_LOC_135/A 0.01fF
C66357 INVX1_LOC_131/Y NAND2X1_LOC_288/B 0.03fF
C66358 NAND2X1_LOC_727/Y NAND2X1_LOC_357/B 0.01fF
C66359 NOR2X1_LOC_561/Y NOR2X1_LOC_142/Y 0.19fF
C66360 NAND2X1_LOC_28/a_36_24# D_INPUT_2 0.00fF
C66361 INVX1_LOC_286/Y INPUT_0 -0.01fF
C66362 INVX1_LOC_240/A NAND2X1_LOC_735/B 0.03fF
C66363 INVX1_LOC_164/Y NAND2X1_LOC_181/Y 0.01fF
C66364 INVX1_LOC_290/A NOR2X1_LOC_52/B 0.02fF
C66365 NOR2X1_LOC_151/Y INVX1_LOC_142/A 0.05fF
C66366 INVX1_LOC_185/A NOR2X1_LOC_654/A 0.00fF
C66367 INVX1_LOC_14/A INVX1_LOC_93/Y 0.10fF
C66368 INVX1_LOC_21/A NAND2X1_LOC_211/Y 0.10fF
C66369 INVX1_LOC_93/A INVX1_LOC_37/A 0.07fF
C66370 INVX1_LOC_12/A NAND2X1_LOC_792/B 0.06fF
C66371 INVX1_LOC_1/Y NOR2X1_LOC_612/B 0.00fF
C66372 NOR2X1_LOC_441/Y NOR2X1_LOC_167/Y 0.03fF
C66373 NAND2X1_LOC_839/Y INVX1_LOC_22/A 0.02fF
C66374 NAND2X1_LOC_315/a_36_24# INVX1_LOC_28/A 0.01fF
C66375 INVX1_LOC_207/A NOR2X1_LOC_525/Y 0.03fF
C66376 INVX1_LOC_251/Y INVX1_LOC_22/A 0.00fF
C66377 NAND2X1_LOC_579/A NOR2X1_LOC_670/a_36_216# 0.03fF
C66378 NAND2X1_LOC_714/B NOR2X1_LOC_305/Y 0.01fF
C66379 NOR2X1_LOC_590/A INVX1_LOC_123/A 0.02fF
C66380 NAND2X1_LOC_361/Y INVX1_LOC_65/Y 0.00fF
C66381 INVX1_LOC_225/A NAND2X1_LOC_808/A -0.03fF
C66382 INVX1_LOC_78/A NOR2X1_LOC_257/Y 0.07fF
C66383 NAND2X1_LOC_513/B INVX1_LOC_37/A 0.02fF
C66384 INVX1_LOC_239/A INVX1_LOC_178/Y 0.01fF
C66385 NOR2X1_LOC_596/A D_INPUT_4 0.01fF
C66386 INVX1_LOC_172/A NOR2X1_LOC_490/Y 0.03fF
C66387 NOR2X1_LOC_647/Y NOR2X1_LOC_391/B 0.39fF
C66388 NOR2X1_LOC_78/B NAND2X1_LOC_112/Y 0.08fF
C66389 INVX1_LOC_269/A INVX1_LOC_20/A 0.05fF
C66390 INVX1_LOC_24/Y NOR2X1_LOC_857/A 0.10fF
C66391 D_INPUT_0 NAND2X1_LOC_357/B 0.07fF
C66392 INVX1_LOC_64/A NOR2X1_LOC_629/Y 0.37fF
C66393 NOR2X1_LOC_232/Y INVX1_LOC_20/A 0.00fF
C66394 NOR2X1_LOC_666/Y NOR2X1_LOC_357/Y 0.14fF
C66395 NOR2X1_LOC_251/Y INVX1_LOC_53/Y 0.00fF
C66396 NOR2X1_LOC_67/Y INVX1_LOC_15/A 0.10fF
C66397 NOR2X1_LOC_631/A NOR2X1_LOC_631/Y 0.41fF
C66398 INVX1_LOC_90/A NAND2X1_LOC_484/a_36_24# 0.00fF
C66399 NOR2X1_LOC_703/B NOR2X1_LOC_703/Y 0.01fF
C66400 INVX1_LOC_14/A NAND2X1_LOC_641/a_36_24# 0.00fF
C66401 NOR2X1_LOC_655/B INVX1_LOC_7/A 0.06fF
C66402 NAND2X1_LOC_223/A INVX1_LOC_125/A 0.02fF
C66403 NOR2X1_LOC_290/Y NOR2X1_LOC_71/Y 0.01fF
C66404 NOR2X1_LOC_68/A INVX1_LOC_78/Y 0.03fF
C66405 INVX1_LOC_14/A NAND2X1_LOC_721/A 0.07fF
C66406 NOR2X1_LOC_122/A NAND2X1_LOC_472/Y 0.20fF
C66407 NOR2X1_LOC_383/B INVX1_LOC_63/A 0.03fF
C66408 NOR2X1_LOC_173/Y NOR2X1_LOC_331/B 0.03fF
C66409 D_INPUT_1 INVX1_LOC_285/A 0.07fF
C66410 INVX1_LOC_90/A NOR2X1_LOC_709/A 0.13fF
C66411 NOR2X1_LOC_552/A NOR2X1_LOC_532/a_36_216# 0.01fF
C66412 NOR2X1_LOC_738/A NOR2X1_LOC_731/A 0.04fF
C66413 NAND2X1_LOC_326/A NOR2X1_LOC_536/A 0.11fF
C66414 INVX1_LOC_57/A NAND2X1_LOC_489/Y 0.03fF
C66415 INVX1_LOC_163/A NAND2X1_LOC_403/a_36_24# 0.00fF
C66416 NAND2X1_LOC_61/Y INVX1_LOC_272/A 0.03fF
C66417 NAND2X1_LOC_363/B NOR2X1_LOC_461/B 0.05fF
C66418 NOR2X1_LOC_389/B NOR2X1_LOC_709/A 0.18fF
C66419 D_INPUT_1 NOR2X1_LOC_814/A 0.06fF
C66420 INVX1_LOC_41/A NOR2X1_LOC_180/a_36_216# 0.00fF
C66421 NAND2X1_LOC_784/A NOR2X1_LOC_661/A 0.01fF
C66422 NOR2X1_LOC_552/A INVX1_LOC_18/A 0.02fF
C66423 NOR2X1_LOC_439/B NOR2X1_LOC_180/Y 0.09fF
C66424 NOR2X1_LOC_441/Y INVX1_LOC_76/A 0.01fF
C66425 INVX1_LOC_292/A INVX1_LOC_14/Y 0.10fF
C66426 INVX1_LOC_161/A VDD 0.00fF
C66427 INVX1_LOC_23/Y INVX1_LOC_284/A 0.02fF
C66428 NAND2X1_LOC_538/Y INVX1_LOC_38/A 0.08fF
C66429 INVX1_LOC_161/A NAND2X1_LOC_800/A 0.04fF
C66430 NOR2X1_LOC_137/A INVX1_LOC_1/Y 0.17fF
C66431 NOR2X1_LOC_380/A NAND2X1_LOC_863/B 0.05fF
C66432 NAND2X1_LOC_208/B VDD 0.30fF
C66433 NOR2X1_LOC_416/A NAND2X1_LOC_215/a_36_24# 0.01fF
C66434 NOR2X1_LOC_789/B INVX1_LOC_46/Y 0.03fF
C66435 INVX1_LOC_185/Y INPUT_0 0.04fF
C66436 NAND2X1_LOC_725/A NOR2X1_LOC_485/Y 0.02fF
C66437 NOR2X1_LOC_250/A INVX1_LOC_38/A 0.01fF
C66438 NOR2X1_LOC_372/A INVX1_LOC_37/Y 0.17fF
C66439 NOR2X1_LOC_121/a_36_216# INPUT_1 0.00fF
C66440 NOR2X1_LOC_445/Y INVX1_LOC_206/Y 0.00fF
C66441 NAND2X1_LOC_859/Y NOR2X1_LOC_71/Y 0.01fF
C66442 INVX1_LOC_182/A INVX1_LOC_179/Y 0.25fF
C66443 NAND2X1_LOC_84/Y INVX1_LOC_93/Y 0.09fF
C66444 NOR2X1_LOC_45/B NOR2X1_LOC_577/Y 0.07fF
C66445 NOR2X1_LOC_447/A NOR2X1_LOC_48/B 0.05fF
C66446 NOR2X1_LOC_589/A NOR2X1_LOC_214/B 0.04fF
C66447 NOR2X1_LOC_332/A NOR2X1_LOC_199/B 0.03fF
C66448 NOR2X1_LOC_652/Y INVX1_LOC_285/A 0.83fF
C66449 INVX1_LOC_7/A NOR2X1_LOC_99/B 0.09fF
C66450 NOR2X1_LOC_722/Y VDD 0.11fF
C66451 NOR2X1_LOC_108/a_36_216# NOR2X1_LOC_814/A 0.00fF
C66452 NOR2X1_LOC_645/a_36_216# NOR2X1_LOC_305/Y 0.00fF
C66453 VDD INVX1_LOC_79/Y 0.41fF
C66454 INVX1_LOC_251/A NAND2X1_LOC_99/A 0.01fF
C66455 NOR2X1_LOC_631/B NOR2X1_LOC_303/Y 0.03fF
C66456 INVX1_LOC_285/Y INVX1_LOC_96/Y 0.65fF
C66457 NOR2X1_LOC_483/a_36_216# NOR2X1_LOC_748/A 0.00fF
C66458 INVX1_LOC_41/A NOR2X1_LOC_405/A 0.03fF
C66459 INVX1_LOC_314/Y NOR2X1_LOC_35/Y 0.10fF
C66460 INVX1_LOC_58/A NAND2X1_LOC_456/a_36_24# 0.01fF
C66461 NAND2X1_LOC_633/Y INVX1_LOC_41/Y 0.00fF
C66462 INVX1_LOC_254/A INVX1_LOC_176/A 0.01fF
C66463 INVX1_LOC_32/A INVX1_LOC_57/A 0.17fF
C66464 INVX1_LOC_119/A INVX1_LOC_91/A 0.02fF
C66465 INVX1_LOC_78/A NOR2X1_LOC_301/A 3.79fF
C66466 NOR2X1_LOC_190/a_36_216# INVX1_LOC_6/A 0.00fF
C66467 INVX1_LOC_18/A NOR2X1_LOC_152/A 0.01fF
C66468 INVX1_LOC_217/A NOR2X1_LOC_495/a_36_216# 0.00fF
C66469 NOR2X1_LOC_91/Y NOR2X1_LOC_301/a_36_216# 0.00fF
C66470 INVX1_LOC_36/A NAND2X1_LOC_476/a_36_24# 0.00fF
C66471 NOR2X1_LOC_500/A INVX1_LOC_37/A 0.01fF
C66472 INVX1_LOC_91/Y INVX1_LOC_22/A 0.01fF
C66473 NOR2X1_LOC_78/B NOR2X1_LOC_737/a_36_216# 0.00fF
C66474 NOR2X1_LOC_631/B NOR2X1_LOC_254/Y 0.33fF
C66475 INVX1_LOC_143/A INVX1_LOC_125/Y 0.41fF
C66476 INVX1_LOC_31/A NAND2X1_LOC_243/Y 0.03fF
C66477 INVX1_LOC_26/A NOR2X1_LOC_278/Y 0.03fF
C66478 INVX1_LOC_57/A NOR2X1_LOC_329/Y 0.10fF
C66479 INVX1_LOC_111/Y NOR2X1_LOC_318/B 0.02fF
C66480 INVX1_LOC_18/A INVX1_LOC_280/A 0.02fF
C66481 NAND2X1_LOC_672/B INVX1_LOC_201/A 0.01fF
C66482 NOR2X1_LOC_78/B INVX1_LOC_98/A 0.07fF
C66483 INVX1_LOC_93/Y NOR2X1_LOC_612/B 0.03fF
C66484 INVX1_LOC_30/A NOR2X1_LOC_641/Y 0.01fF
C66485 NOR2X1_LOC_142/Y INVX1_LOC_76/A 0.02fF
C66486 INVX1_LOC_41/A NOR2X1_LOC_857/A 0.07fF
C66487 NOR2X1_LOC_78/B NOR2X1_LOC_78/A 0.11fF
C66488 NAND2X1_LOC_141/A INVX1_LOC_316/A 0.50fF
C66489 NOR2X1_LOC_440/Y NOR2X1_LOC_188/A 0.01fF
C66490 NOR2X1_LOC_524/a_36_216# INVX1_LOC_91/A 0.09fF
C66491 INVX1_LOC_34/A VDD 1.46fF
C66492 INVX1_LOC_57/A NAND2X1_LOC_175/Y 0.07fF
C66493 NOR2X1_LOC_254/Y INVX1_LOC_37/A 0.32fF
C66494 NOR2X1_LOC_84/Y INVX1_LOC_74/A 0.01fF
C66495 INVX1_LOC_45/A NAND2X1_LOC_798/B 0.10fF
C66496 NOR2X1_LOC_334/Y NOR2X1_LOC_493/a_36_216# 0.00fF
C66497 INVX1_LOC_177/A NOR2X1_LOC_137/a_36_216# 0.00fF
C66498 INVX1_LOC_34/A NAND2X1_LOC_800/A 0.07fF
C66499 NOR2X1_LOC_625/Y NOR2X1_LOC_536/A 0.01fF
C66500 NAND2X1_LOC_231/Y NOR2X1_LOC_56/Y 0.10fF
C66501 NOR2X1_LOC_15/Y NAND2X1_LOC_81/B 0.03fF
C66502 NOR2X1_LOC_631/B NOR2X1_LOC_353/Y 0.01fF
C66503 NOR2X1_LOC_486/Y NOR2X1_LOC_352/Y 0.00fF
C66504 NOR2X1_LOC_792/B NAND2X1_LOC_287/B 0.02fF
C66505 INVX1_LOC_172/A INVX1_LOC_280/A 0.00fF
C66506 NAND2X1_LOC_454/Y NOR2X1_LOC_717/A 0.01fF
C66507 NOR2X1_LOC_45/B INVX1_LOC_22/A 0.75fF
C66508 INVX1_LOC_28/A NAND2X1_LOC_123/Y 0.04fF
C66509 NOR2X1_LOC_304/Y INVX1_LOC_231/A 0.02fF
C66510 NAND2X1_LOC_104/a_36_24# NOR2X1_LOC_649/B 0.01fF
C66511 NOR2X1_LOC_405/A NOR2X1_LOC_211/A 0.03fF
C66512 INVX1_LOC_48/Y NAND2X1_LOC_254/Y 0.03fF
C66513 INVX1_LOC_1/A NOR2X1_LOC_89/A 0.12fF
C66514 NAND2X1_LOC_811/Y NAND2X1_LOC_811/B 0.05fF
C66515 NOR2X1_LOC_655/B INVX1_LOC_76/A 0.10fF
C66516 NOR2X1_LOC_778/B NOR2X1_LOC_35/Y 1.47fF
C66517 NOR2X1_LOC_222/Y NAND2X1_LOC_469/B 0.12fF
C66518 NOR2X1_LOC_489/B INVX1_LOC_87/A 0.01fF
C66519 NOR2X1_LOC_71/Y INVX1_LOC_6/A 0.13fF
C66520 NAND2X1_LOC_470/a_36_24# NAND2X1_LOC_453/A 0.00fF
C66521 INVX1_LOC_41/Y INVX1_LOC_71/Y 0.01fF
C66522 NAND2X1_LOC_231/Y VDD 2.35fF
C66523 NOR2X1_LOC_359/Y INVX1_LOC_307/A 0.01fF
C66524 NAND2X1_LOC_596/a_36_24# NAND2X1_LOC_453/A 0.00fF
C66525 NAND2X1_LOC_361/Y NAND2X1_LOC_617/a_36_24# 0.00fF
C66526 INVX1_LOC_89/A INVX1_LOC_309/A -0.00fF
C66527 NOR2X1_LOC_361/B NAND2X1_LOC_288/a_36_24# 0.06fF
C66528 INVX1_LOC_304/Y NOR2X1_LOC_495/a_36_216# 0.01fF
C66529 NOR2X1_LOC_564/Y NOR2X1_LOC_74/A 0.05fF
C66530 NAND2X1_LOC_357/B NAND2X1_LOC_848/A 0.10fF
C66531 NOR2X1_LOC_113/B NOR2X1_LOC_772/A 0.00fF
C66532 INVX1_LOC_150/A INVX1_LOC_91/A 0.02fF
C66533 NOR2X1_LOC_449/a_36_216# NOR2X1_LOC_592/B 0.00fF
C66534 INVX1_LOC_17/A INVX1_LOC_42/A 9.88fF
C66535 INVX1_LOC_83/A NOR2X1_LOC_78/A 0.30fF
C66536 NOR2X1_LOC_561/A NOR2X1_LOC_709/A 0.01fF
C66537 NOR2X1_LOC_137/A NOR2X1_LOC_318/B 0.07fF
C66538 NOR2X1_LOC_817/Y NOR2X1_LOC_847/a_36_216# 0.00fF
C66539 INVX1_LOC_132/A INVX1_LOC_92/A 0.10fF
C66540 NOR2X1_LOC_211/A NOR2X1_LOC_857/A 0.08fF
C66541 INVX1_LOC_89/A INVX1_LOC_91/A 0.25fF
C66542 INVX1_LOC_178/A INVX1_LOC_94/Y 0.10fF
C66543 NOR2X1_LOC_218/A INVX1_LOC_290/Y 0.11fF
C66544 INVX1_LOC_45/Y NOR2X1_LOC_117/Y 0.24fF
C66545 NAND2X1_LOC_30/Y NAND2X1_LOC_430/B 0.03fF
C66546 INVX1_LOC_49/A NOR2X1_LOC_831/B 0.08fF
C66547 D_GATE_366 INVX1_LOC_159/Y 0.01fF
C66548 NAND2X1_LOC_112/Y INVX1_LOC_46/A 0.04fF
C66549 INVX1_LOC_269/A INVX1_LOC_4/A 0.55fF
C66550 NOR2X1_LOC_15/Y INVX1_LOC_4/Y 0.15fF
C66551 NOR2X1_LOC_721/Y INPUT_0 0.06fF
C66552 INVX1_LOC_11/A NOR2X1_LOC_467/A 0.03fF
C66553 INVX1_LOC_5/A INVX1_LOC_296/A 0.00fF
C66554 NOR2X1_LOC_288/a_36_216# INVX1_LOC_15/A 0.02fF
C66555 NAND2X1_LOC_550/A INVX1_LOC_19/Y 0.00fF
C66556 INVX1_LOC_225/A INVX1_LOC_92/A 0.07fF
C66557 NOR2X1_LOC_99/B INVX1_LOC_76/A 0.11fF
C66558 INVX1_LOC_14/A INVX1_LOC_87/A 0.03fF
C66559 NOR2X1_LOC_290/Y NAND2X1_LOC_243/Y 0.00fF
C66560 INVX1_LOC_69/Y NOR2X1_LOC_188/A 0.17fF
C66561 NOR2X1_LOC_781/A INVX1_LOC_117/A 0.12fF
C66562 NAND2X1_LOC_163/a_36_24# NAND2X1_LOC_425/Y 0.00fF
C66563 INVX1_LOC_24/A INVX1_LOC_19/A 2.24fF
C66564 INVX1_LOC_17/A INVX1_LOC_78/A 0.68fF
C66565 INVX1_LOC_69/Y NOR2X1_LOC_548/B 0.15fF
C66566 INVX1_LOC_171/Y INVX1_LOC_57/A 0.13fF
C66567 INVX1_LOC_24/A NOR2X1_LOC_11/Y 0.03fF
C66568 INVX1_LOC_14/A INVX1_LOC_175/A 0.03fF
C66569 NOR2X1_LOC_148/B VDD 0.25fF
C66570 NAND2X1_LOC_360/B NAND2X1_LOC_93/B 0.32fF
C66571 NOR2X1_LOC_67/A NOR2X1_LOC_99/Y 0.22fF
C66572 NOR2X1_LOC_652/Y NOR2X1_LOC_292/a_36_216# 0.00fF
C66573 NOR2X1_LOC_186/Y INVX1_LOC_53/A 0.51fF
C66574 INVX1_LOC_56/Y INVX1_LOC_118/A 0.31fF
C66575 NOR2X1_LOC_816/A INVX1_LOC_94/Y 0.46fF
C66576 INVX1_LOC_31/A INVX1_LOC_21/Y 0.04fF
C66577 NOR2X1_LOC_471/Y INVX1_LOC_78/A 0.09fF
C66578 NOR2X1_LOC_193/a_36_216# NOR2X1_LOC_78/A 0.00fF
C66579 INVX1_LOC_104/A INVX1_LOC_84/A 0.07fF
C66580 NOR2X1_LOC_112/Y NOR2X1_LOC_332/a_36_216# 0.02fF
C66581 NOR2X1_LOC_226/A NOR2X1_LOC_831/B 0.18fF
C66582 NOR2X1_LOC_552/A NOR2X1_LOC_548/A 0.02fF
C66583 INVX1_LOC_17/A NOR2X1_LOC_65/B 1.27fF
C66584 NOR2X1_LOC_93/Y INVX1_LOC_64/A 0.01fF
C66585 NOR2X1_LOC_805/a_36_216# NOR2X1_LOC_383/B 0.00fF
C66586 NOR2X1_LOC_106/A INVX1_LOC_38/A 0.12fF
C66587 NOR2X1_LOC_639/B NOR2X1_LOC_454/Y 0.08fF
C66588 INVX1_LOC_131/A VDD 0.18fF
C66589 INVX1_LOC_53/Y NOR2X1_LOC_216/B 0.01fF
C66590 NAND2X1_LOC_360/B INVX1_LOC_3/A -0.01fF
C66591 NAND2X1_LOC_724/A INVX1_LOC_53/A 0.05fF
C66592 INVX1_LOC_31/A INVX1_LOC_16/Y 0.10fF
C66593 NOR2X1_LOC_738/A INVX1_LOC_117/A 0.02fF
C66594 NAND2X1_LOC_656/A INVX1_LOC_251/A 0.15fF
C66595 NAND2X1_LOC_139/A NOR2X1_LOC_671/Y 0.02fF
C66596 INVX1_LOC_35/A NOR2X1_LOC_468/Y 0.03fF
C66597 INVX1_LOC_25/A INVX1_LOC_11/A 0.11fF
C66598 NOR2X1_LOC_735/Y INVX1_LOC_281/A -0.02fF
C66599 INVX1_LOC_135/A NOR2X1_LOC_860/Y 0.01fF
C66600 INVX1_LOC_286/Y INVX1_LOC_183/A 0.02fF
C66601 INVX1_LOC_71/A INVX1_LOC_47/Y 0.10fF
C66602 INVX1_LOC_174/Y NAND2X1_LOC_425/Y 0.05fF
C66603 NOR2X1_LOC_667/A NOR2X1_LOC_605/A 0.04fF
C66604 INPUT_0 VDD 2.80fF
C66605 INVX1_LOC_155/Y INVX1_LOC_290/Y 0.14fF
C66606 INPUT_3 INVX1_LOC_57/A 0.03fF
C66607 INVX1_LOC_64/A INVX1_LOC_269/A 0.13fF
C66608 NOR2X1_LOC_667/Y NOR2X1_LOC_654/A 0.00fF
C66609 NOR2X1_LOC_802/A INVX1_LOC_29/A 0.01fF
C66610 NOR2X1_LOC_52/B INVX1_LOC_261/Y 0.02fF
C66611 INVX1_LOC_263/A INVX1_LOC_84/A 1.24fF
C66612 INVX1_LOC_143/A INVX1_LOC_19/A 0.07fF
C66613 INVX1_LOC_133/Y INVX1_LOC_272/A 0.28fF
C66614 INVX1_LOC_144/A NOR2X1_LOC_111/A 0.06fF
C66615 INVX1_LOC_72/A INVX1_LOC_23/Y 0.01fF
C66616 INVX1_LOC_299/A INVX1_LOC_5/A 0.07fF
C66617 INVX1_LOC_235/Y INVX1_LOC_27/A 0.09fF
C66618 INVX1_LOC_18/A NOR2X1_LOC_541/B 0.03fF
C66619 NAND2X1_LOC_149/Y INVX1_LOC_27/A 0.09fF
C66620 NAND2X1_LOC_796/B NAND2X1_LOC_703/Y 0.03fF
C66621 D_INPUT_1 NOR2X1_LOC_590/A 1.05fF
C66622 NOR2X1_LOC_355/A NOR2X1_LOC_155/A 0.03fF
C66623 INVX1_LOC_177/A INVX1_LOC_99/A 0.03fF
C66624 NOR2X1_LOC_45/Y INVX1_LOC_53/A 0.03fF
C66625 NOR2X1_LOC_557/A NOR2X1_LOC_35/Y 1.19fF
C66626 INVX1_LOC_21/A NAND2X1_LOC_578/a_36_24# 0.01fF
C66627 NOR2X1_LOC_538/B INVX1_LOC_5/A 0.03fF
C66628 NAND2X1_LOC_84/Y INVX1_LOC_87/A 0.04fF
C66629 NOR2X1_LOC_84/Y NAND2X1_LOC_254/Y 0.10fF
C66630 INVX1_LOC_16/A NAND2X1_LOC_625/a_36_24# 0.01fF
C66631 NOR2X1_LOC_303/Y NAND2X1_LOC_72/B 0.08fF
C66632 NAND2X1_LOC_564/B NOR2X1_LOC_662/A 0.02fF
C66633 INVX1_LOC_40/A INVX1_LOC_125/A 0.01fF
C66634 NAND2X1_LOC_854/B INVX1_LOC_84/A 0.19fF
C66635 NOR2X1_LOC_482/Y NAND2X1_LOC_254/Y 0.06fF
C66636 INPUT_1 NOR2X1_LOC_101/a_36_216# 0.00fF
C66637 INVX1_LOC_35/A NOR2X1_LOC_389/A 0.03fF
C66638 NOR2X1_LOC_68/A NOR2X1_LOC_727/B 0.03fF
C66639 NOR2X1_LOC_550/B INVX1_LOC_271/Y 0.10fF
C66640 INVX1_LOC_24/A INVX1_LOC_26/Y 2.30fF
C66641 NAND2X1_LOC_182/A INVX1_LOC_15/A 0.01fF
C66642 NOR2X1_LOC_78/A INVX1_LOC_46/A 1.58fF
C66643 INVX1_LOC_104/A INVX1_LOC_15/A 0.16fF
C66644 INVX1_LOC_293/A INVX1_LOC_5/A 0.01fF
C66645 INVX1_LOC_291/Y INVX1_LOC_76/A 0.03fF
C66646 INVX1_LOC_35/A NAND2X1_LOC_199/B 0.02fF
C66647 NOR2X1_LOC_137/B NOR2X1_LOC_137/a_36_216# 0.00fF
C66648 NOR2X1_LOC_147/B NOR2X1_LOC_334/Y 0.01fF
C66649 NOR2X1_LOC_130/A NOR2X1_LOC_653/Y 0.02fF
C66650 INVX1_LOC_22/A NOR2X1_LOC_1/Y 0.00fF
C66651 VDD NAND2X1_LOC_649/B 0.01fF
C66652 INVX1_LOC_45/Y INVX1_LOC_270/A 1.05fF
C66653 NOR2X1_LOC_567/B NOR2X1_LOC_809/B 0.06fF
C66654 INVX1_LOC_58/A NOR2X1_LOC_457/B 0.10fF
C66655 INVX1_LOC_213/Y INVX1_LOC_274/Y 0.11fF
C66656 NOR2X1_LOC_392/B NOR2X1_LOC_334/Y 0.01fF
C66657 NOR2X1_LOC_237/Y NOR2X1_LOC_693/Y 0.42fF
C66658 INVX1_LOC_232/A INVX1_LOC_284/A 0.45fF
C66659 NOR2X1_LOC_590/A NOR2X1_LOC_108/a_36_216# 0.00fF
C66660 NOR2X1_LOC_15/Y NOR2X1_LOC_205/Y 0.07fF
C66661 NOR2X1_LOC_328/Y NOR2X1_LOC_226/Y 0.01fF
C66662 INVX1_LOC_89/A INVX1_LOC_203/A 0.03fF
C66663 NOR2X1_LOC_348/B NOR2X1_LOC_465/Y 0.29fF
C66664 NOR2X1_LOC_252/Y INVX1_LOC_42/A 0.12fF
C66665 NOR2X1_LOC_130/A INVX1_LOC_19/A 0.17fF
C66666 INVX1_LOC_11/A INVX1_LOC_1/A 1.16fF
C66667 NOR2X1_LOC_389/B INVX1_LOC_294/A 0.01fF
C66668 NOR2X1_LOC_612/B INVX1_LOC_87/A 0.08fF
C66669 NAND2X1_LOC_711/B NAND2X1_LOC_794/a_36_24# 0.00fF
C66670 NOR2X1_LOC_82/A INVX1_LOC_14/A 3.88fF
C66671 NAND2X1_LOC_267/B NAND2X1_LOC_266/a_36_24# 0.02fF
C66672 INVX1_LOC_54/Y NAND2X1_LOC_72/B 0.06fF
C66673 INVX1_LOC_263/A INVX1_LOC_15/A 0.01fF
C66674 INVX1_LOC_21/A INVX1_LOC_210/Y 0.13fF
C66675 INVX1_LOC_12/Y INVX1_LOC_20/A 0.10fF
C66676 NAND2X1_LOC_560/A NOR2X1_LOC_485/Y 0.00fF
C66677 NOR2X1_LOC_309/Y NAND2X1_LOC_288/B 0.01fF
C66678 INVX1_LOC_269/A INVX1_LOC_43/Y 0.03fF
C66679 INVX1_LOC_58/A NAND2X1_LOC_833/Y 0.03fF
C66680 INVX1_LOC_20/A NOR2X1_LOC_492/Y 0.04fF
C66681 NOR2X1_LOC_790/B INVX1_LOC_49/A 0.02fF
C66682 INVX1_LOC_223/Y NOR2X1_LOC_703/B 0.00fF
C66683 NOR2X1_LOC_639/B INVX1_LOC_77/A 0.09fF
C66684 INVX1_LOC_11/A NOR2X1_LOC_794/B 0.03fF
C66685 INVX1_LOC_46/A NOR2X1_LOC_60/Y 0.14fF
C66686 NAND2X1_LOC_338/B INVX1_LOC_23/Y 0.04fF
C66687 INVX1_LOC_143/A INVX1_LOC_26/Y 0.08fF
C66688 NOR2X1_LOC_590/A NOR2X1_LOC_241/A 0.01fF
C66689 INVX1_LOC_22/A NOR2X1_LOC_465/Y 0.02fF
C66690 NOR2X1_LOC_527/Y NOR2X1_LOC_661/A 0.09fF
C66691 INVX1_LOC_25/A NOR2X1_LOC_52/B 0.07fF
C66692 NOR2X1_LOC_817/Y INVX1_LOC_31/A 0.49fF
C66693 INVX1_LOC_35/A NOR2X1_LOC_712/Y 0.43fF
C66694 INVX1_LOC_225/A INVX1_LOC_53/A 0.08fF
C66695 INVX1_LOC_174/A NOR2X1_LOC_160/B 0.12fF
C66696 INVX1_LOC_133/Y NOR2X1_LOC_125/a_36_216# 0.02fF
C66697 NOR2X1_LOC_288/A INVX1_LOC_53/A 0.37fF
C66698 NOR2X1_LOC_843/A NOR2X1_LOC_434/A 0.05fF
C66699 INVX1_LOC_82/Y INVX1_LOC_29/A 0.02fF
C66700 INVX1_LOC_35/A NOR2X1_LOC_295/Y 0.02fF
C66701 NOR2X1_LOC_773/Y INVX1_LOC_181/A 0.01fF
C66702 NOR2X1_LOC_123/B INVX1_LOC_47/Y 0.12fF
C66703 NAND2X1_LOC_354/a_36_24# INVX1_LOC_246/A 0.00fF
C66704 INVX1_LOC_35/A NOR2X1_LOC_844/A 0.03fF
C66705 NOR2X1_LOC_349/A NAND2X1_LOC_574/A 0.05fF
C66706 INVX1_LOC_17/A NOR2X1_LOC_554/B 0.29fF
C66707 NOR2X1_LOC_447/Y NOR2X1_LOC_454/Y 0.00fF
C66708 NOR2X1_LOC_254/A INVX1_LOC_30/A 0.07fF
C66709 INVX1_LOC_21/A INVX1_LOC_155/A 0.39fF
C66710 INVX1_LOC_230/Y NOR2X1_LOC_382/Y 0.80fF
C66711 INVX1_LOC_1/Y NOR2X1_LOC_383/B 0.07fF
C66712 INVX1_LOC_97/A NOR2X1_LOC_334/Y 0.03fF
C66713 INVX1_LOC_200/A NOR2X1_LOC_91/Y 0.16fF
C66714 NAND2X1_LOC_552/A NOR2X1_LOC_315/Y 0.00fF
C66715 NOR2X1_LOC_188/A NOR2X1_LOC_89/A 0.22fF
C66716 INVX1_LOC_64/A NOR2X1_LOC_648/a_36_216# 0.01fF
C66717 INVX1_LOC_200/Y NAND2X1_LOC_543/Y 0.13fF
C66718 INVX1_LOC_16/A INVX1_LOC_271/A 0.07fF
C66719 INVX1_LOC_21/A NOR2X1_LOC_264/Y 0.07fF
C66720 INVX1_LOC_90/A NOR2X1_LOC_334/Y 0.07fF
C66721 INVX1_LOC_1/A NOR2X1_LOC_433/A 0.16fF
C66722 NOR2X1_LOC_548/B NOR2X1_LOC_89/A 0.05fF
C66723 INVX1_LOC_136/A INVX1_LOC_188/A 0.01fF
C66724 INVX1_LOC_35/A NOR2X1_LOC_220/A 0.07fF
C66725 INVX1_LOC_24/A INVX1_LOC_161/Y 0.11fF
C66726 NOR2X1_LOC_322/a_36_216# INVX1_LOC_185/A 0.00fF
C66727 NAND2X1_LOC_861/Y NOR2X1_LOC_301/A 0.01fF
C66728 NOR2X1_LOC_647/A INVX1_LOC_135/A 0.04fF
C66729 INVX1_LOC_255/Y NOR2X1_LOC_416/A 0.01fF
C66730 INVX1_LOC_1/A NOR2X1_LOC_593/Y 0.20fF
C66731 INVX1_LOC_17/A NOR2X1_LOC_152/Y 0.08fF
C66732 INVX1_LOC_215/A INVX1_LOC_23/A 0.07fF
C66733 INVX1_LOC_58/A NOR2X1_LOC_781/A 0.01fF
C66734 NOR2X1_LOC_498/Y NAND2X1_LOC_706/Y 0.06fF
C66735 NAND2X1_LOC_551/A NAND2X1_LOC_477/a_36_24# 0.01fF
C66736 INVX1_LOC_37/A NAND2X1_LOC_412/a_36_24# 0.01fF
C66737 NOR2X1_LOC_860/Y INVX1_LOC_280/A 0.04fF
C66738 INVX1_LOC_123/A NOR2X1_LOC_67/Y 0.08fF
C66739 INVX1_LOC_24/A NOR2X1_LOC_553/a_36_216# 0.02fF
C66740 NOR2X1_LOC_510/Y NAND2X1_LOC_231/Y 0.10fF
C66741 NOR2X1_LOC_226/A NAND2X1_LOC_169/Y 0.02fF
C66742 NOR2X1_LOC_443/Y D_INPUT_0 0.13fF
C66743 INVX1_LOC_140/A INVX1_LOC_94/Y 0.03fF
C66744 NOR2X1_LOC_163/Y NAND2X1_LOC_452/Y 0.03fF
C66745 D_INPUT_1 INVX1_LOC_227/A 0.07fF
C66746 INVX1_LOC_34/A NOR2X1_LOC_361/B 0.01fF
C66747 NOR2X1_LOC_186/Y NOR2X1_LOC_78/B 0.07fF
C66748 NOR2X1_LOC_280/Y NOR2X1_LOC_653/Y 0.40fF
C66749 INVX1_LOC_5/A INVX1_LOC_52/A 0.01fF
C66750 NOR2X1_LOC_690/Y NAND2X1_LOC_794/a_36_24# 0.00fF
C66751 NOR2X1_LOC_456/Y INVX1_LOC_279/A 0.22fF
C66752 NAND2X1_LOC_303/Y INVX1_LOC_240/A 0.03fF
C66753 INVX1_LOC_22/A NOR2X1_LOC_53/Y 0.02fF
C66754 NOR2X1_LOC_15/Y INVX1_LOC_194/A 0.06fF
C66755 NOR2X1_LOC_824/A NAND2X1_LOC_717/Y 0.11fF
C66756 INVX1_LOC_103/A NAND2X1_LOC_466/Y 0.03fF
C66757 INVX1_LOC_1/A NOR2X1_LOC_52/B 0.10fF
C66758 NOR2X1_LOC_471/Y INVX1_LOC_113/Y 1.37fF
C66759 NOR2X1_LOC_785/A INVX1_LOC_49/A 0.01fF
C66760 NOR2X1_LOC_331/B NAND2X1_LOC_798/B 0.07fF
C66761 INVX1_LOC_95/Y NAND2X1_LOC_74/B 0.23fF
C66762 NAND2X1_LOC_214/B INVX1_LOC_16/A 0.58fF
C66763 INVX1_LOC_24/A NOR2X1_LOC_599/A 0.97fF
C66764 INVX1_LOC_206/Y INVX1_LOC_15/A 0.07fF
C66765 NAND2X1_LOC_746/a_36_24# NAND2X1_LOC_662/Y 0.00fF
C66766 INVX1_LOC_58/A NOR2X1_LOC_76/A 0.02fF
C66767 NAND2X1_LOC_573/Y NOR2X1_LOC_78/B 0.01fF
C66768 NOR2X1_LOC_536/A NAND2X1_LOC_572/B 0.01fF
C66769 INVX1_LOC_39/A NOR2X1_LOC_121/a_36_216# 0.00fF
C66770 INVX1_LOC_21/A INVX1_LOC_316/Y 0.03fF
C66771 NAND2X1_LOC_391/Y INVX1_LOC_25/Y 0.06fF
C66772 INVX1_LOC_13/A INVX1_LOC_306/Y 0.10fF
C66773 INVX1_LOC_136/A NOR2X1_LOC_238/Y 0.03fF
C66774 NOR2X1_LOC_222/Y INVX1_LOC_52/Y 0.02fF
C66775 NAND2X1_LOC_549/Y D_INPUT_0 0.00fF
C66776 NOR2X1_LOC_831/B INVX1_LOC_118/A 0.07fF
C66777 NOR2X1_LOC_205/Y INVX1_LOC_96/Y 0.03fF
C66778 INVX1_LOC_140/A INVX1_LOC_181/A 0.02fF
C66779 NOR2X1_LOC_668/a_36_216# INVX1_LOC_89/A 0.01fF
C66780 INVX1_LOC_178/Y NAND2X1_LOC_82/Y 0.03fF
C66781 INVX1_LOC_27/A INVX1_LOC_16/A 0.14fF
C66782 NAND2X1_LOC_651/a_36_24# INVX1_LOC_296/A 0.03fF
C66783 INVX1_LOC_28/A INVX1_LOC_271/A 0.42fF
C66784 NOR2X1_LOC_533/A NAND2X1_LOC_303/Y 0.04fF
C66785 INVX1_LOC_140/A INVX1_LOC_296/A 0.10fF
C66786 NOR2X1_LOC_824/A INVX1_LOC_16/A 0.11fF
C66787 INVX1_LOC_17/A NOR2X1_LOC_721/A 0.03fF
C66788 INVX1_LOC_233/Y NOR2X1_LOC_576/B 0.07fF
C66789 NOR2X1_LOC_742/A NOR2X1_LOC_383/B 0.07fF
C66790 NOR2X1_LOC_600/Y INVX1_LOC_15/A 0.01fF
C66791 NOR2X1_LOC_15/Y NAND2X1_LOC_862/A 0.01fF
C66792 INVX1_LOC_64/A NOR2X1_LOC_214/B 0.02fF
C66793 INVX1_LOC_286/Y NAND2X1_LOC_811/Y 0.15fF
C66794 INVX1_LOC_281/A INVX1_LOC_186/Y 1.12fF
C66795 NOR2X1_LOC_637/B NAND2X1_LOC_354/Y 0.32fF
C66796 INVX1_LOC_234/Y NAND2X1_LOC_735/B 0.16fF
C66797 NAND2X1_LOC_571/Y NAND2X1_LOC_632/a_36_24# 0.00fF
C66798 NOR2X1_LOC_647/A NOR2X1_LOC_391/B 0.07fF
C66799 NAND2X1_LOC_741/Y NOR2X1_LOC_298/Y 0.04fF
C66800 D_INPUT_0 NOR2X1_LOC_291/Y 0.16fF
C66801 NAND2X1_LOC_798/B NOR2X1_LOC_592/B 0.06fF
C66802 NAND2X1_LOC_220/a_36_24# NAND2X1_LOC_220/B 0.00fF
C66803 NAND2X1_LOC_725/A NAND2X1_LOC_644/a_36_24# 0.06fF
C66804 INVX1_LOC_174/A INVX1_LOC_189/A 0.02fF
C66805 NAND2X1_LOC_93/B NAND2X1_LOC_572/B 0.07fF
C66806 NOR2X1_LOC_456/Y INVX1_LOC_182/Y 0.10fF
C66807 INVX1_LOC_258/A INVX1_LOC_22/A 0.01fF
C66808 NOR2X1_LOC_92/Y NOR2X1_LOC_32/Y 0.01fF
C66809 NOR2X1_LOC_61/Y NOR2X1_LOC_814/A 0.07fF
C66810 NOR2X1_LOC_91/A INVX1_LOC_286/A 0.12fF
C66811 NAND2X1_LOC_181/a_36_24# INVX1_LOC_14/A 0.01fF
C66812 NAND2X1_LOC_787/A NOR2X1_LOC_322/Y 0.01fF
C66813 NOR2X1_LOC_791/B INVX1_LOC_8/A 0.08fF
C66814 INVX1_LOC_135/A NOR2X1_LOC_173/Y 0.00fF
C66815 NOR2X1_LOC_750/A NAND2X1_LOC_749/a_36_24# 0.00fF
C66816 NOR2X1_LOC_52/B NOR2X1_LOC_384/Y 0.03fF
C66817 NAND2X1_LOC_725/B NOR2X1_LOC_298/Y 0.08fF
C66818 NAND2X1_LOC_35/Y NOR2X1_LOC_393/a_36_216# 0.01fF
C66819 INVX1_LOC_178/A NAND2X1_LOC_624/A 0.02fF
C66820 INVX1_LOC_6/A NAND2X1_LOC_205/A 0.02fF
C66821 NOR2X1_LOC_598/B NOR2X1_LOC_541/a_36_216# 0.01fF
C66822 NOR2X1_LOC_6/B NOR2X1_LOC_360/Y 0.03fF
C66823 NOR2X1_LOC_106/Y INVX1_LOC_67/A 0.74fF
C66824 NAND2X1_LOC_748/a_36_24# INVX1_LOC_89/A 0.00fF
C66825 INVX1_LOC_179/A INVX1_LOC_63/A 0.00fF
C66826 NOR2X1_LOC_673/a_36_216# INVX1_LOC_46/Y 0.01fF
C66827 INVX1_LOC_304/Y NOR2X1_LOC_91/Y 0.08fF
C66828 INVX1_LOC_286/A INVX1_LOC_23/A 0.07fF
C66829 INVX1_LOC_14/A INVX1_LOC_306/A 0.00fF
C66830 NOR2X1_LOC_318/B NOR2X1_LOC_383/B 0.07fF
C66831 INVX1_LOC_77/A INVX1_LOC_155/Y 0.03fF
C66832 INVX1_LOC_254/Y INVX1_LOC_41/A 0.00fF
C66833 INVX1_LOC_21/A NAND2X1_LOC_850/A 0.03fF
C66834 INVX1_LOC_27/A INVX1_LOC_28/A 0.07fF
C66835 NOR2X1_LOC_567/B INVX1_LOC_50/Y 0.08fF
C66836 NOR2X1_LOC_160/B NOR2X1_LOC_589/A 0.03fF
C66837 NOR2X1_LOC_91/A INVX1_LOC_95/A 1.06fF
C66838 NOR2X1_LOC_824/A INVX1_LOC_28/A 0.10fF
C66839 NAND2X1_LOC_363/B INVX1_LOC_92/Y 0.02fF
C66840 NOR2X1_LOC_48/Y INVX1_LOC_92/A 0.03fF
C66841 NOR2X1_LOC_218/Y INVX1_LOC_81/Y 0.32fF
C66842 INVX1_LOC_24/Y NOR2X1_LOC_542/Y 0.01fF
C66843 NOR2X1_LOC_266/a_36_216# NOR2X1_LOC_191/A -0.00fF
C66844 NAND2X1_LOC_54/a_36_24# INVX1_LOC_136/A 0.01fF
C66845 INVX1_LOC_93/Y NOR2X1_LOC_383/B 0.07fF
C66846 INVX1_LOC_19/A NOR2X1_LOC_197/B 0.01fF
C66847 NAND2X1_LOC_783/A INVX1_LOC_161/Y 0.01fF
C66848 NOR2X1_LOC_277/a_36_216# INVX1_LOC_286/A 0.00fF
C66849 INVX1_LOC_17/A NAND2X1_LOC_861/Y 0.07fF
C66850 INVX1_LOC_314/Y NOR2X1_LOC_84/Y 0.04fF
C66851 INVX1_LOC_161/Y NOR2X1_LOC_130/A 0.07fF
C66852 INVX1_LOC_34/A INVX1_LOC_153/Y 0.01fF
C66853 INVX1_LOC_90/A INVX1_LOC_308/Y 0.01fF
C66854 INVX1_LOC_233/A INVX1_LOC_98/A 0.10fF
C66855 NOR2X1_LOC_454/Y INVX1_LOC_302/A 0.06fF
C66856 NAND2X1_LOC_9/Y NOR2X1_LOC_78/A 0.05fF
C66857 NOR2X1_LOC_392/Y INVX1_LOC_91/A -0.03fF
C66858 INVX1_LOC_255/Y INVX1_LOC_36/A 0.03fF
C66859 INVX1_LOC_95/A INVX1_LOC_23/A 0.03fF
C66860 NOR2X1_LOC_52/Y INVX1_LOC_22/A 0.30fF
C66861 NAND2X1_LOC_703/Y NAND2X1_LOC_840/Y 0.02fF
C66862 INVX1_LOC_233/A NOR2X1_LOC_78/A 0.12fF
C66863 INVX1_LOC_3/A NAND2X1_LOC_219/B 0.40fF
C66864 INVX1_LOC_283/Y INVX1_LOC_266/Y -0.04fF
C66865 NOR2X1_LOC_274/Y NOR2X1_LOC_655/B 0.34fF
C66866 NOR2X1_LOC_690/A INVX1_LOC_240/A 0.10fF
C66867 NAND2X1_LOC_149/Y NOR2X1_LOC_589/a_36_216# 0.01fF
C66868 INVX1_LOC_21/A INVX1_LOC_86/A 0.01fF
C66869 NAND2X1_LOC_792/B INVX1_LOC_92/A 0.01fF
C66870 NOR2X1_LOC_160/B INVX1_LOC_171/A 0.01fF
C66871 NOR2X1_LOC_589/A NAND2X1_LOC_195/Y 0.01fF
C66872 NOR2X1_LOC_446/A INVX1_LOC_313/Y 0.03fF
C66873 NOR2X1_LOC_279/Y INVX1_LOC_57/A 0.01fF
C66874 INVX1_LOC_33/A NOR2X1_LOC_709/A 0.10fF
C66875 NOR2X1_LOC_334/Y INVX1_LOC_38/A 0.14fF
C66876 INVX1_LOC_25/A INVX1_LOC_74/A 0.13fF
C66877 NOR2X1_LOC_591/Y NAND2X1_LOC_354/B 0.06fF
C66878 NOR2X1_LOC_738/Y NOR2X1_LOC_738/A 0.04fF
C66879 NOR2X1_LOC_383/Y INVX1_LOC_72/A 0.03fF
C66880 NOR2X1_LOC_423/Y INVX1_LOC_63/Y 0.02fF
C66881 INVX1_LOC_58/A NAND2X1_LOC_241/Y 0.07fF
C66882 NAND2X1_LOC_151/a_36_24# INVX1_LOC_28/A 0.00fF
C66883 NAND2X1_LOC_553/A INVX1_LOC_98/A 0.08fF
C66884 INVX1_LOC_34/A INVX1_LOC_177/A 0.03fF
C66885 INVX1_LOC_30/Y NOR2X1_LOC_360/Y 0.03fF
C66886 NOR2X1_LOC_78/B NOR2X1_LOC_374/A 0.41fF
C66887 INVX1_LOC_36/Y NOR2X1_LOC_105/Y 0.13fF
C66888 NOR2X1_LOC_599/A NAND2X1_LOC_800/Y 0.00fF
C66889 INVX1_LOC_312/A NOR2X1_LOC_130/A 0.01fF
C66890 NOR2X1_LOC_615/Y NOR2X1_LOC_497/Y 0.07fF
C66891 NOR2X1_LOC_554/B NOR2X1_LOC_199/B 0.41fF
C66892 INVX1_LOC_36/A NOR2X1_LOC_71/Y 0.07fF
C66893 INVX1_LOC_249/A INVX1_LOC_16/A 0.03fF
C66894 NOR2X1_LOC_238/a_36_216# NAND2X1_LOC_859/Y 0.00fF
C66895 NAND2X1_LOC_579/A NOR2X1_LOC_167/Y 0.03fF
C66896 INVX1_LOC_35/A NAND2X1_LOC_469/B 0.03fF
C66897 INVX1_LOC_223/Y INVX1_LOC_91/A 0.04fF
C66898 NOR2X1_LOC_216/Y INVX1_LOC_161/Y 0.07fF
C66899 NOR2X1_LOC_361/B INPUT_0 0.03fF
C66900 NOR2X1_LOC_798/A NOR2X1_LOC_78/A 0.03fF
C66901 NOR2X1_LOC_186/Y NOR2X1_LOC_311/Y 0.01fF
C66902 INVX1_LOC_34/A INVX1_LOC_280/Y 6.70fF
C66903 NOR2X1_LOC_222/Y INVX1_LOC_63/Y 0.22fF
C66904 INVX1_LOC_6/Y INVX1_LOC_16/A 0.01fF
C66905 INVX1_LOC_2/A NAND2X1_LOC_357/B 0.07fF
C66906 NOR2X1_LOC_647/A INVX1_LOC_280/A 0.05fF
C66907 NOR2X1_LOC_273/Y INVX1_LOC_279/A 0.00fF
C66908 NOR2X1_LOC_288/A NOR2X1_LOC_634/B 0.00fF
C66909 INVX1_LOC_224/A NOR2X1_LOC_188/A 0.15fF
C66910 INVX1_LOC_225/A NOR2X1_LOC_78/B 0.07fF
C66911 NAND2X1_LOC_338/B NAND2X1_LOC_116/A 0.15fF
C66912 INVX1_LOC_174/A NOR2X1_LOC_706/A 0.18fF
C66913 NOR2X1_LOC_416/a_36_216# INVX1_LOC_2/Y 0.00fF
C66914 INVX1_LOC_279/A NOR2X1_LOC_759/Y 0.01fF
C66915 NAND2X1_LOC_860/A INVX1_LOC_37/A 0.01fF
C66916 INVX1_LOC_224/A NOR2X1_LOC_548/B 0.02fF
C66917 NOR2X1_LOC_91/A NOR2X1_LOC_602/B 0.03fF
C66918 INVX1_LOC_202/A INVX1_LOC_279/A 0.48fF
C66919 NOR2X1_LOC_226/A NAND2X1_LOC_357/B 0.07fF
C66920 NOR2X1_LOC_536/A NOR2X1_LOC_654/A 0.03fF
C66921 INVX1_LOC_58/A NAND2X1_LOC_837/a_36_24# 0.00fF
C66922 NOR2X1_LOC_458/B NOR2X1_LOC_348/B 0.02fF
C66923 INVX1_LOC_11/A NOR2X1_LOC_548/B 0.03fF
C66924 NAND2X1_LOC_573/Y NOR2X1_LOC_311/Y 0.01fF
C66925 NOR2X1_LOC_607/Y INVX1_LOC_227/A 0.01fF
C66926 NAND2X1_LOC_364/A NOR2X1_LOC_768/a_36_216# 0.00fF
C66927 INVX1_LOC_106/Y INVX1_LOC_125/A 0.00fF
C66928 NOR2X1_LOC_91/A INVX1_LOC_54/A 0.13fF
C66929 INVX1_LOC_279/A NOR2X1_LOC_550/B 0.10fF
C66930 NOR2X1_LOC_240/Y VDD 0.12fF
C66931 NAND2X1_LOC_9/Y NOR2X1_LOC_98/a_36_216# 0.00fF
C66932 NOR2X1_LOC_448/B INVX1_LOC_91/A 0.01fF
C66933 NOR2X1_LOC_82/A INVX1_LOC_48/A 0.02fF
C66934 INVX1_LOC_81/A NAND2X1_LOC_140/A 0.01fF
C66935 INVX1_LOC_40/A NOR2X1_LOC_709/A 0.08fF
C66936 NOR2X1_LOC_449/A NAND2X1_LOC_798/B 0.09fF
C66937 NOR2X1_LOC_322/Y INVX1_LOC_30/A 0.01fF
C66938 INVX1_LOC_132/A INVX1_LOC_83/A 0.07fF
C66939 INVX1_LOC_305/A NAND2X1_LOC_172/a_36_24# 0.01fF
C66940 NAND2X1_LOC_286/B NOR2X1_LOC_743/Y 0.11fF
C66941 INVX1_LOC_27/A NOR2X1_LOC_35/Y 0.11fF
C66942 INVX1_LOC_83/A NOR2X1_LOC_374/A 0.08fF
C66943 NOR2X1_LOC_220/B VDD 0.24fF
C66944 INVX1_LOC_303/A INVX1_LOC_148/Y 0.01fF
C66945 NOR2X1_LOC_237/Y NOR2X1_LOC_71/Y 0.14fF
C66946 NAND2X1_LOC_578/B NAND2X1_LOC_577/a_36_24# 0.04fF
C66947 NOR2X1_LOC_186/Y INVX1_LOC_46/A 0.66fF
C66948 NAND2X1_LOC_19/a_36_24# INVX1_LOC_315/Y 0.00fF
C66949 NOR2X1_LOC_234/Y NOR2X1_LOC_86/A 0.01fF
C66950 NAND2X1_LOC_361/Y NAND2X1_LOC_364/a_36_24# 0.00fF
C66951 INVX1_LOC_225/Y NOR2X1_LOC_337/Y 0.04fF
C66952 INVX1_LOC_1/A INVX1_LOC_199/A 0.07fF
C66953 NOR2X1_LOC_394/Y INVX1_LOC_3/A 0.01fF
C66954 INVX1_LOC_23/A INVX1_LOC_54/A 0.50fF
C66955 NAND2X1_LOC_725/A NOR2X1_LOC_694/Y 0.06fF
C66956 INVX1_LOC_25/A NOR2X1_LOC_675/a_36_216# 0.00fF
C66957 INVX1_LOC_26/Y NOR2X1_LOC_197/B 0.08fF
C66958 NOR2X1_LOC_703/B INVX1_LOC_75/A 0.05fF
C66959 NOR2X1_LOC_716/B NOR2X1_LOC_749/a_36_216# 0.00fF
C66960 INVX1_LOC_10/A INVX1_LOC_88/Y 0.01fF
C66961 NOR2X1_LOC_629/A NOR2X1_LOC_629/Y 0.00fF
C66962 INVX1_LOC_33/A NOR2X1_LOC_106/A 0.01fF
C66963 INVX1_LOC_5/A NAND2X1_LOC_96/A 0.08fF
C66964 NAND2X1_LOC_338/B INVX1_LOC_232/A 0.10fF
C66965 INVX1_LOC_1/A INVX1_LOC_74/A 0.07fF
C66966 INVX1_LOC_14/A INVX1_LOC_59/Y 0.03fF
C66967 NOR2X1_LOC_128/A NOR2X1_LOC_554/A 0.00fF
C66968 NAND2X1_LOC_563/Y INVX1_LOC_80/A 0.02fF
C66969 INVX1_LOC_90/A INVX1_LOC_209/Y 0.09fF
C66970 INVX1_LOC_14/A INVX1_LOC_112/A 0.08fF
C66971 NOR2X1_LOC_92/Y NOR2X1_LOC_825/Y 0.03fF
C66972 NOR2X1_LOC_523/B NAND2X1_LOC_348/A 0.03fF
C66973 NAND2X1_LOC_276/Y INVX1_LOC_89/A 0.11fF
C66974 NOR2X1_LOC_589/A INVX1_LOC_189/A 0.04fF
C66975 INVX1_LOC_182/Y NOR2X1_LOC_759/Y 0.00fF
C66976 NAND2X1_LOC_573/Y INVX1_LOC_46/A 0.35fF
C66977 NAND2X1_LOC_579/A INVX1_LOC_76/A 0.08fF
C66978 INVX1_LOC_41/A NOR2X1_LOC_542/Y 0.03fF
C66979 NOR2X1_LOC_34/Y NOR2X1_LOC_814/A 0.05fF
C66980 NOR2X1_LOC_318/A INVX1_LOC_285/A 0.01fF
C66981 NAND2X1_LOC_848/A NOR2X1_LOC_291/Y 1.22fF
C66982 NOR2X1_LOC_458/B INVX1_LOC_22/A 0.00fF
C66983 INVX1_LOC_202/A INVX1_LOC_182/Y 0.04fF
C66984 NOR2X1_LOC_644/A NOR2X1_LOC_804/B 0.01fF
C66985 NOR2X1_LOC_723/Y NOR2X1_LOC_733/Y 0.03fF
C66986 NOR2X1_LOC_383/Y NAND2X1_LOC_338/B 0.00fF
C66987 NOR2X1_LOC_401/A INVX1_LOC_20/A 0.15fF
C66988 INVX1_LOC_27/Y NAND2X1_LOC_99/A 0.25fF
C66989 INVX1_LOC_77/A INVX1_LOC_302/A 0.02fF
C66990 INVX1_LOC_90/A NOR2X1_LOC_718/B 0.42fF
C66991 INVX1_LOC_41/A INVX1_LOC_311/Y 0.09fF
C66992 NAND2X1_LOC_738/B NAND2X1_LOC_770/Y 0.10fF
C66993 NAND2X1_LOC_537/Y INVX1_LOC_37/A 0.08fF
C66994 INVX1_LOC_24/A NAND2X1_LOC_270/a_36_24# 0.01fF
C66995 NOR2X1_LOC_209/Y INVX1_LOC_83/A 0.10fF
C66996 NOR2X1_LOC_695/Y INVX1_LOC_16/A 0.02fF
C66997 NAND2X1_LOC_288/B INVX1_LOC_63/A 0.05fF
C66998 NAND2X1_LOC_550/A INVX1_LOC_20/A 0.37fF
C66999 NOR2X1_LOC_238/a_36_216# INVX1_LOC_6/A -0.00fF
C67000 INVX1_LOC_186/A INVX1_LOC_142/Y 0.00fF
C67001 NOR2X1_LOC_654/A NOR2X1_LOC_661/A 0.01fF
C67002 NOR2X1_LOC_160/B INVX1_LOC_20/A 0.12fF
C67003 INVX1_LOC_286/A INVX1_LOC_111/A 0.01fF
C67004 INVX1_LOC_229/Y NAND2X1_LOC_853/Y 0.00fF
C67005 INVX1_LOC_18/A NOR2X1_LOC_45/B 0.21fF
C67006 INVX1_LOC_204/Y INVX1_LOC_92/A 0.04fF
C67007 INVX1_LOC_94/Y INVX1_LOC_42/A 0.42fF
C67008 INVX1_LOC_225/Y VDD 1.26fF
C67009 INVX1_LOC_241/A NOR2X1_LOC_298/Y 0.66fF
C67010 INVX1_LOC_234/A INVX1_LOC_16/A 0.20fF
C67011 INVX1_LOC_186/A INVX1_LOC_198/Y 0.81fF
C67012 D_INPUT_0 NOR2X1_LOC_382/a_36_216# 0.00fF
C67013 INVX1_LOC_206/A INVX1_LOC_28/A 0.01fF
C67014 NOR2X1_LOC_593/Y NOR2X1_LOC_188/A 0.06fF
C67015 NOR2X1_LOC_315/Y INVX1_LOC_140/A 0.01fF
C67016 INVX1_LOC_45/A NOR2X1_LOC_726/a_36_216# 0.02fF
C67017 INVX1_LOC_136/A INVX1_LOC_95/Y 0.23fF
C67018 NOR2X1_LOC_593/Y NOR2X1_LOC_548/B 0.10fF
C67019 INVX1_LOC_90/A INVX1_LOC_218/A 0.05fF
C67020 INVX1_LOC_43/Y INVX1_LOC_12/Y 0.01fF
C67021 INVX1_LOC_39/A NOR2X1_LOC_101/a_36_216# 0.00fF
C67022 NOR2X1_LOC_637/Y NOR2X1_LOC_45/B 0.03fF
C67023 NOR2X1_LOC_272/Y NOR2X1_LOC_155/A 1.73fF
C67024 INVX1_LOC_34/A INVX1_LOC_285/Y 0.03fF
C67025 NOR2X1_LOC_392/Y INVX1_LOC_203/A 0.10fF
C67026 INVX1_LOC_1/A NOR2X1_LOC_675/a_36_216# 0.01fF
C67027 INVX1_LOC_45/A NOR2X1_LOC_112/a_36_216# 0.00fF
C67028 NOR2X1_LOC_658/Y NOR2X1_LOC_364/a_36_216# 0.01fF
C67029 INVX1_LOC_271/A INVX1_LOC_109/A 0.03fF
C67030 INVX1_LOC_172/A NOR2X1_LOC_45/B 0.07fF
C67031 NOR2X1_LOC_775/Y NAND2X1_LOC_323/B 0.07fF
C67032 NAND2X1_LOC_656/Y INVX1_LOC_10/A 0.14fF
C67033 INVX1_LOC_29/A INVX1_LOC_29/Y 0.13fF
C67034 NOR2X1_LOC_251/Y INVX1_LOC_28/A -0.10fF
C67035 NOR2X1_LOC_91/A NOR2X1_LOC_48/B 0.27fF
C67036 INVX1_LOC_50/A INVX1_LOC_102/A 0.11fF
C67037 INVX1_LOC_89/A NOR2X1_LOC_553/B 0.03fF
C67038 NOR2X1_LOC_751/a_36_216# NOR2X1_LOC_197/B 0.03fF
C67039 INPUT_0 INVX1_LOC_177/A 0.03fF
C67040 INVX1_LOC_90/A NOR2X1_LOC_569/Y 0.07fF
C67041 NOR2X1_LOC_772/A INVX1_LOC_16/A 0.09fF
C67042 NAND2X1_LOC_807/B INVX1_LOC_23/A 0.98fF
C67043 NAND2X1_LOC_213/A NOR2X1_LOC_155/A 0.02fF
C67044 INVX1_LOC_57/Y NAND2X1_LOC_721/A 0.15fF
C67045 NOR2X1_LOC_92/Y NOR2X1_LOC_88/Y 0.07fF
C67046 INVX1_LOC_173/Y INPUT_5 0.08fF
C67047 INVX1_LOC_45/A INVX1_LOC_33/Y 0.01fF
C67048 INVX1_LOC_54/Y NOR2X1_LOC_113/B 0.02fF
C67049 NOR2X1_LOC_19/B INVX1_LOC_16/A 0.80fF
C67050 INVX1_LOC_72/Y VDD 0.46fF
C67051 NAND2X1_LOC_802/A NOR2X1_LOC_56/Y 0.01fF
C67052 INVX1_LOC_17/A INVX1_LOC_291/A 0.09fF
C67053 INVX1_LOC_78/A INVX1_LOC_94/Y 0.06fF
C67054 INVX1_LOC_280/Y INPUT_0 0.22fF
C67055 NOR2X1_LOC_48/B INVX1_LOC_23/A 0.07fF
C67056 INVX1_LOC_197/A NAND2X1_LOC_622/B 0.30fF
C67057 INVX1_LOC_246/Y VDD 0.26fF
C67058 NOR2X1_LOC_75/Y NAND2X1_LOC_93/B 0.03fF
C67059 INVX1_LOC_21/A NOR2X1_LOC_662/A 1.73fF
C67060 INVX1_LOC_31/A INVX1_LOC_54/A 0.15fF
C67061 NOR2X1_LOC_106/Y NOR2X1_LOC_137/Y 0.01fF
C67062 NOR2X1_LOC_92/Y INVX1_LOC_84/A 0.69fF
C67063 NAND2X1_LOC_349/B INVX1_LOC_79/A 0.01fF
C67064 INVX1_LOC_63/Y NOR2X1_LOC_69/A 0.03fF
C67065 NOR2X1_LOC_764/a_36_216# NAND2X1_LOC_51/B 0.00fF
C67066 NOR2X1_LOC_486/Y NAND2X1_LOC_484/a_36_24# 0.00fF
C67067 NOR2X1_LOC_65/B INVX1_LOC_94/Y 1.02fF
C67068 NOR2X1_LOC_643/Y VDD 0.12fF
C67069 INVX1_LOC_135/A INVX1_LOC_148/A 0.05fF
C67070 INVX1_LOC_78/A INVX1_LOC_181/A 0.03fF
C67071 NAND2X1_LOC_773/Y INVX1_LOC_293/Y 0.00fF
C67072 NOR2X1_LOC_240/Y NAND2X1_LOC_232/a_36_24# 0.00fF
C67073 INVX1_LOC_78/A INVX1_LOC_296/A 0.01fF
C67074 NOR2X1_LOC_577/Y NOR2X1_LOC_139/a_36_216# 0.02fF
C67075 INPUT_3 NOR2X1_LOC_820/Y 0.10fF
C67076 INVX1_LOC_55/Y NOR2X1_LOC_356/A -0.00fF
C67077 INVX1_LOC_59/A NAND2X1_LOC_74/B 0.03fF
C67078 NOR2X1_LOC_78/B NAND2X1_LOC_642/Y 0.03fF
C67079 NAND2X1_LOC_811/Y VDD 0.25fF
C67080 NOR2X1_LOC_620/Y INVX1_LOC_117/A 0.00fF
C67081 NOR2X1_LOC_486/B INVX1_LOC_37/A 0.04fF
C67082 INVX1_LOC_61/Y INVX1_LOC_123/Y 0.01fF
C67083 NOR2X1_LOC_419/Y NOR2X1_LOC_536/A 0.01fF
C67084 INVX1_LOC_225/A INVX1_LOC_46/A 0.21fF
C67085 INVX1_LOC_25/Y INVX1_LOC_91/A 0.01fF
C67086 INVX1_LOC_224/Y INVX1_LOC_23/Y 0.07fF
C67087 NAND2X1_LOC_773/Y NAND2X1_LOC_74/B 0.03fF
C67088 NAND2X1_LOC_811/Y NAND2X1_LOC_800/A 0.00fF
C67089 NOR2X1_LOC_68/A NOR2X1_LOC_640/Y 0.10fF
C67090 INVX1_LOC_298/Y INVX1_LOC_29/Y 0.07fF
C67091 INVX1_LOC_140/A NOR2X1_LOC_166/Y 0.11fF
C67092 VDD NOR2X1_LOC_821/Y 0.12fF
C67093 INVX1_LOC_32/A INVX1_LOC_306/Y 0.03fF
C67094 NOR2X1_LOC_147/B NAND2X1_LOC_472/Y 0.10fF
C67095 NAND2X1_LOC_349/B INVX1_LOC_91/A 0.02fF
C67096 NOR2X1_LOC_716/B NOR2X1_LOC_536/A 0.20fF
C67097 NOR2X1_LOC_507/A NOR2X1_LOC_349/A 0.11fF
C67098 NOR2X1_LOC_373/Y INVX1_LOC_6/A 0.02fF
C67099 VDD INVX1_LOC_266/Y 4.20fF
C67100 NOR2X1_LOC_609/A NAND2X1_LOC_93/B 0.03fF
C67101 NOR2X1_LOC_617/Y NOR2X1_LOC_629/Y 0.00fF
C67102 NOR2X1_LOC_593/a_36_216# INVX1_LOC_139/Y 0.00fF
C67103 NOR2X1_LOC_725/A INVX1_LOC_174/Y 0.02fF
C67104 NAND2X1_LOC_364/A NOR2X1_LOC_155/A 0.15fF
C67105 INVX1_LOC_48/A INVX1_LOC_306/A 0.01fF
C67106 NAND2X1_LOC_374/Y NAND2X1_LOC_244/A 0.00fF
C67107 NOR2X1_LOC_289/Y NAND2X1_LOC_652/Y 0.01fF
C67108 INVX1_LOC_45/A INVX1_LOC_220/A 0.23fF
C67109 NOR2X1_LOC_162/Y INVX1_LOC_38/A 0.01fF
C67110 INVX1_LOC_55/Y NOR2X1_LOC_74/A 0.22fF
C67111 INVX1_LOC_286/Y NOR2X1_LOC_653/Y 0.00fF
C67112 NAND2X1_LOC_200/B NOR2X1_LOC_35/Y 0.13fF
C67113 NOR2X1_LOC_731/A INVX1_LOC_117/A 0.02fF
C67114 NOR2X1_LOC_359/Y INVX1_LOC_92/A 0.26fF
C67115 INVX1_LOC_299/A INVX1_LOC_42/A 0.07fF
C67116 NOR2X1_LOC_68/A NAND2X1_LOC_85/Y 0.05fF
C67117 INVX1_LOC_290/A NOR2X1_LOC_657/B 0.12fF
C67118 NAND2X1_LOC_853/Y INVX1_LOC_20/A 0.03fF
C67119 INVX1_LOC_155/Y INVX1_LOC_9/A 0.03fF
C67120 INVX1_LOC_88/A NOR2X1_LOC_114/Y 0.07fF
C67121 NOR2X1_LOC_641/B INVX1_LOC_63/A 0.05fF
C67122 NAND2X1_LOC_392/Y NAND2X1_LOC_642/Y 0.03fF
C67123 NOR2X1_LOC_419/Y NAND2X1_LOC_93/B 0.16fF
C67124 NOR2X1_LOC_718/B INVX1_LOC_38/A 0.03fF
C67125 NAND2X1_LOC_852/Y INVX1_LOC_46/A 0.49fF
C67126 INVX1_LOC_208/Y INVX1_LOC_76/A 0.01fF
C67127 NOR2X1_LOC_516/B INVX1_LOC_20/A 0.03fF
C67128 NOR2X1_LOC_92/Y INVX1_LOC_15/A 6.31fF
C67129 NAND2X1_LOC_837/Y NOR2X1_LOC_88/Y 0.36fF
C67130 INVX1_LOC_24/A NOR2X1_LOC_841/A 0.01fF
C67131 NOR2X1_LOC_594/Y NAND2X1_LOC_661/A 0.18fF
C67132 INVX1_LOC_24/Y INVX1_LOC_15/A 0.10fF
C67133 INVX1_LOC_305/A NOR2X1_LOC_814/A 0.07fF
C67134 NOR2X1_LOC_716/B NAND2X1_LOC_93/B 0.07fF
C67135 NOR2X1_LOC_172/Y NAND2X1_LOC_434/Y 0.17fF
C67136 NOR2X1_LOC_751/Y INVX1_LOC_63/A 0.01fF
C67137 NOR2X1_LOC_78/B NOR2X1_LOC_863/A 0.05fF
C67138 INVX1_LOC_286/Y NOR2X1_LOC_11/Y 0.03fF
C67139 INVX1_LOC_83/A NAND2X1_LOC_642/Y 0.08fF
C67140 INVX1_LOC_293/A INVX1_LOC_42/A 0.00fF
C67141 NOR2X1_LOC_270/Y NAND2X1_LOC_476/Y 0.01fF
C67142 NAND2X1_LOC_357/B INVX1_LOC_118/A 1.20fF
C67143 NAND2X1_LOC_656/A INVX1_LOC_27/Y 0.02fF
C67144 NOR2X1_LOC_75/a_36_216# INVX1_LOC_54/A 0.00fF
C67145 NAND2X1_LOC_842/B INVX1_LOC_98/A 0.06fF
C67146 NOR2X1_LOC_589/A NAND2X1_LOC_211/Y 0.42fF
C67147 NAND2X1_LOC_852/Y NOR2X1_LOC_766/Y 0.03fF
C67148 NAND2X1_LOC_853/Y NOR2X1_LOC_765/Y 0.36fF
C67149 INVX1_LOC_28/A NOR2X1_LOC_528/Y 0.07fF
C67150 NAND2X1_LOC_842/B NOR2X1_LOC_78/A 0.03fF
C67151 NOR2X1_LOC_778/Y NOR2X1_LOC_777/B 0.02fF
C67152 NOR2X1_LOC_768/a_36_216# NOR2X1_LOC_405/A 0.00fF
C67153 INVX1_LOC_310/Y NAND2X1_LOC_412/a_36_24# 0.00fF
C67154 INVX1_LOC_159/A INVX1_LOC_19/A 0.07fF
C67155 INVX1_LOC_31/A NOR2X1_LOC_48/B 0.15fF
C67156 NOR2X1_LOC_459/A D_GATE_662 0.01fF
C67157 NOR2X1_LOC_586/a_36_216# NOR2X1_LOC_586/Y 0.00fF
C67158 INVX1_LOC_75/A NOR2X1_LOC_114/A 0.15fF
C67159 INVX1_LOC_299/A INVX1_LOC_78/A 0.07fF
C67160 INVX1_LOC_243/Y INVX1_LOC_21/A 0.01fF
C67161 INVX1_LOC_18/A NOR2X1_LOC_1/Y 0.12fF
C67162 INVX1_LOC_313/Y NAND2X1_LOC_447/Y 0.10fF
C67163 INVX1_LOC_75/A INVX1_LOC_91/A 3.33fF
C67164 NOR2X1_LOC_160/B INVX1_LOC_4/A 1.36fF
C67165 INVX1_LOC_21/A INVX1_LOC_57/A 0.17fF
C67166 NOR2X1_LOC_272/Y NOR2X1_LOC_125/Y 0.34fF
C67167 INVX1_LOC_41/A INVX1_LOC_84/A 0.03fF
C67168 NOR2X1_LOC_381/Y INVX1_LOC_26/A 0.01fF
C67169 INVX1_LOC_286/A INVX1_LOC_6/A 0.15fF
C67170 NOR2X1_LOC_569/Y INVX1_LOC_38/A 0.07fF
C67171 NOR2X1_LOC_457/A NOR2X1_LOC_464/Y 0.00fF
C67172 NOR2X1_LOC_168/B NOR2X1_LOC_445/B 0.12fF
C67173 INVX1_LOC_68/Y INVX1_LOC_108/A 0.09fF
C67174 NAND2X1_LOC_354/Y NAND2X1_LOC_419/a_36_24# 0.00fF
C67175 NOR2X1_LOC_103/Y INVX1_LOC_23/Y 0.09fF
C67176 NAND2X1_LOC_140/A NOR2X1_LOC_363/Y 0.19fF
C67177 INVX1_LOC_255/Y NOR2X1_LOC_656/Y 0.01fF
C67178 INPUT_0 INVX1_LOC_65/A 0.07fF
C67179 NOR2X1_LOC_456/Y NOR2X1_LOC_456/a_36_216# 0.00fF
C67180 NAND2X1_LOC_474/Y NOR2X1_LOC_717/A 0.42fF
C67181 INPUT_0 INVX1_LOC_316/A 0.01fF
C67182 NAND2X1_LOC_859/Y INVX1_LOC_54/A 0.01fF
C67183 INVX1_LOC_90/A NAND2X1_LOC_472/Y 0.07fF
C67184 NOR2X1_LOC_392/B NAND2X1_LOC_773/B 0.10fF
C67185 NAND2X1_LOC_479/Y NOR2X1_LOC_433/Y 0.01fF
C67186 NAND2X1_LOC_53/Y NOR2X1_LOC_727/B 0.01fF
C67187 NOR2X1_LOC_598/B NAND2X1_LOC_213/A 0.03fF
C67188 NOR2X1_LOC_82/A NOR2X1_LOC_383/B 0.03fF
C67189 INVX1_LOC_222/Y INVX1_LOC_5/A 0.03fF
C67190 NOR2X1_LOC_524/Y INVX1_LOC_78/A 0.01fF
C67191 INVX1_LOC_278/A NOR2X1_LOC_92/Y 0.09fF
C67192 INVX1_LOC_16/A NOR2X1_LOC_216/B 0.06fF
C67193 NAND2X1_LOC_483/Y INVX1_LOC_12/A 0.43fF
C67194 NOR2X1_LOC_590/A NOR2X1_LOC_318/A 0.03fF
C67195 NOR2X1_LOC_67/A NOR2X1_LOC_673/A 0.02fF
C67196 NOR2X1_LOC_456/Y NAND2X1_LOC_190/Y 0.20fF
C67197 INVX1_LOC_21/A NAND2X1_LOC_608/a_36_24# 0.00fF
C67198 NOR2X1_LOC_186/Y NOR2X1_LOC_798/A 0.01fF
C67199 INVX1_LOC_136/A INVX1_LOC_271/Y 0.07fF
C67200 INVX1_LOC_42/Y VDD 0.76fF
C67201 NOR2X1_LOC_357/Y NOR2X1_LOC_74/A 0.56fF
C67202 INVX1_LOC_11/A NAND2X1_LOC_784/A 0.01fF
C67203 NAND2X1_LOC_139/A INVX1_LOC_284/A 0.02fF
C67204 NOR2X1_LOC_91/A NOR2X1_LOC_441/Y 0.05fF
C67205 INVX1_LOC_13/A NOR2X1_LOC_865/Y 0.07fF
C67206 INVX1_LOC_45/A INVX1_LOC_23/Y 0.07fF
C67207 INVX1_LOC_246/A INVX1_LOC_271/A 0.39fF
C67208 NOR2X1_LOC_667/A NOR2X1_LOC_662/A 0.01fF
C67209 INVX1_LOC_269/A NAND2X1_LOC_624/B 0.05fF
C67210 NAND2X1_LOC_214/B INVX1_LOC_48/Y 0.02fF
C67211 NAND2X1_LOC_350/A INVX1_LOC_23/A 0.04fF
C67212 INVX1_LOC_36/A INVX1_LOC_16/Y 0.01fF
C67213 NAND2X1_LOC_577/a_36_24# INVX1_LOC_203/A 0.00fF
C67214 INVX1_LOC_24/A INVX1_LOC_128/A 0.05fF
C67215 NAND2X1_LOC_656/Y INVX1_LOC_307/A 0.00fF
C67216 NOR2X1_LOC_311/Y NAND2X1_LOC_642/Y 0.05fF
C67217 INVX1_LOC_13/A NOR2X1_LOC_243/B 0.07fF
C67218 NOR2X1_LOC_186/Y NAND2X1_LOC_703/Y 0.79fF
C67219 INVX1_LOC_269/A NOR2X1_LOC_662/a_36_216# 0.01fF
C67220 INVX1_LOC_255/Y NOR2X1_LOC_642/a_36_216# 0.01fF
C67221 NAND2X1_LOC_866/B INVX1_LOC_54/A 0.00fF
C67222 INVX1_LOC_176/A INVX1_LOC_48/A 0.02fF
C67223 NOR2X1_LOC_65/B NOR2X1_LOC_524/Y 0.02fF
C67224 INVX1_LOC_256/A INVX1_LOC_58/Y 1.48fF
C67225 NOR2X1_LOC_844/A NAND2X1_LOC_206/B 0.17fF
C67226 INVX1_LOC_31/A NAND2X1_LOC_215/A 0.56fF
C67227 INVX1_LOC_191/A VDD 0.00fF
C67228 INVX1_LOC_282/A NOR2X1_LOC_492/Y 0.03fF
C67229 NOR2X1_LOC_139/Y NAND2X1_LOC_468/B 0.03fF
C67230 INVX1_LOC_315/Y INVX1_LOC_20/A 0.03fF
C67231 NOR2X1_LOC_315/Y INVX1_LOC_42/A 0.02fF
C67232 NOR2X1_LOC_480/A INVX1_LOC_175/A 0.01fF
C67233 INVX1_LOC_41/A INVX1_LOC_15/A 0.24fF
C67234 NOR2X1_LOC_441/Y INVX1_LOC_23/A 0.29fF
C67235 NAND2X1_LOC_807/Y INVX1_LOC_54/A 0.07fF
C67236 NOR2X1_LOC_589/Y INVX1_LOC_117/A 0.11fF
C67237 INVX1_LOC_50/A INVX1_LOC_223/A 0.03fF
C67238 INVX1_LOC_64/A NAND2X1_LOC_550/A 0.10fF
C67239 INVX1_LOC_255/Y INVX1_LOC_63/A 0.04fF
C67240 NOR2X1_LOC_619/A NOR2X1_LOC_721/B 0.02fF
C67241 NOR2X1_LOC_152/Y INVX1_LOC_94/Y 0.00fF
C67242 NAND2X1_LOC_573/Y NAND2X1_LOC_703/Y 0.23fF
C67243 NAND2X1_LOC_813/a_36_24# NOR2X1_LOC_35/Y 0.06fF
C67244 NAND2X1_LOC_638/Y NAND2X1_LOC_428/a_36_24# 0.00fF
C67245 NOR2X1_LOC_130/A NOR2X1_LOC_841/A 0.17fF
C67246 NOR2X1_LOC_590/A NOR2X1_LOC_678/A 0.03fF
C67247 INVX1_LOC_64/A NOR2X1_LOC_160/B 0.25fF
C67248 VDD INVX1_LOC_125/Y 0.21fF
C67249 NAND2X1_LOC_849/A INVX1_LOC_118/A 0.01fF
C67250 NOR2X1_LOC_296/Y INVX1_LOC_306/Y 0.07fF
C67251 NAND2X1_LOC_198/B NAND2X1_LOC_286/B 0.01fF
C67252 NOR2X1_LOC_635/A D_INPUT_5 0.01fF
C67253 INVX1_LOC_91/A NAND2X1_LOC_453/A 0.07fF
C67254 INVX1_LOC_33/A NOR2X1_LOC_334/Y 0.17fF
C67255 NAND2X1_LOC_541/Y INVX1_LOC_284/A 0.02fF
C67256 NAND2X1_LOC_354/Y INVX1_LOC_57/A 0.18fF
C67257 INVX1_LOC_71/A INVX1_LOC_23/Y 0.03fF
C67258 INVX1_LOC_34/A INVX1_LOC_4/Y 0.03fF
C67259 INVX1_LOC_83/A NAND2X1_LOC_252/a_36_24# 0.00fF
C67260 INVX1_LOC_191/Y NOR2X1_LOC_48/B 0.06fF
C67261 NOR2X1_LOC_433/A NOR2X1_LOC_338/a_36_216# 0.01fF
C67262 NOR2X1_LOC_598/B NOR2X1_LOC_336/B 0.00fF
C67263 NAND2X1_LOC_9/Y INVX1_LOC_170/A 0.01fF
C67264 NAND2X1_LOC_477/A INVX1_LOC_15/A 0.01fF
C67265 NOR2X1_LOC_582/Y INVX1_LOC_57/A 0.32fF
C67266 INVX1_LOC_28/A NOR2X1_LOC_216/B 0.02fF
C67267 NAND2X1_LOC_642/Y INVX1_LOC_46/A 7.10fF
C67268 NOR2X1_LOC_134/Y NOR2X1_LOC_291/Y 0.27fF
C67269 INVX1_LOC_225/A NOR2X1_LOC_282/a_36_216# 0.00fF
C67270 NOR2X1_LOC_71/Y INVX1_LOC_63/A 0.07fF
C67271 INVX1_LOC_101/A INVX1_LOC_29/A 0.01fF
C67272 NOR2X1_LOC_742/A INVX1_LOC_179/A 0.26fF
C67273 INVX1_LOC_5/A NAND2X1_LOC_577/A 0.07fF
C67274 INVX1_LOC_101/Y INVX1_LOC_88/A 0.02fF
C67275 NAND2X1_LOC_72/Y INVX1_LOC_223/A 0.12fF
C67276 NAND2X1_LOC_860/A NAND2X1_LOC_198/B 0.24fF
C67277 INVX1_LOC_11/A NAND2X1_LOC_326/A 0.03fF
C67278 INVX1_LOC_90/A NAND2X1_LOC_206/Y 0.01fF
C67279 INVX1_LOC_64/A NAND2X1_LOC_195/Y 0.03fF
C67280 NAND2X1_LOC_303/Y NOR2X1_LOC_533/Y 0.03fF
C67281 INVX1_LOC_6/A INVX1_LOC_54/A 0.87fF
C67282 NOR2X1_LOC_443/Y INVX1_LOC_49/A 0.03fF
C67283 NOR2X1_LOC_180/a_36_216# NOR2X1_LOC_155/A 0.00fF
C67284 NOR2X1_LOC_315/Y INVX1_LOC_78/A 0.03fF
C67285 INVX1_LOC_25/A INVX1_LOC_314/Y 0.07fF
C67286 NOR2X1_LOC_714/Y NOR2X1_LOC_334/Y 0.02fF
C67287 NOR2X1_LOC_421/Y NAND2X1_LOC_453/A 0.01fF
C67288 NOR2X1_LOC_201/A NOR2X1_LOC_340/Y 0.59fF
C67289 NOR2X1_LOC_644/A INVX1_LOC_63/A 0.03fF
C67290 NAND2X1_LOC_656/Y INVX1_LOC_12/A 0.07fF
C67291 NOR2X1_LOC_355/A INVX1_LOC_29/A 0.08fF
C67292 INVX1_LOC_286/A NOR2X1_LOC_79/A 0.04fF
C67293 NOR2X1_LOC_6/B INVX1_LOC_26/A 0.04fF
C67294 INVX1_LOC_178/A NAND2X1_LOC_577/A 0.80fF
C67295 INVX1_LOC_89/A INVX1_LOC_125/A 0.13fF
C67296 INVX1_LOC_75/A NOR2X1_LOC_179/Y 0.03fF
C67297 INVX1_LOC_208/A INVX1_LOC_4/A 0.03fF
C67298 NOR2X1_LOC_516/B INVX1_LOC_4/A 0.11fF
C67299 INVX1_LOC_50/A INVX1_LOC_149/Y 0.12fF
C67300 INVX1_LOC_11/A NAND2X1_LOC_807/A 0.02fF
C67301 INVX1_LOC_5/A NAND2X1_LOC_656/A 0.08fF
C67302 NOR2X1_LOC_142/Y INVX1_LOC_23/A 0.10fF
C67303 NAND2X1_LOC_348/A NAND2X1_LOC_206/Y 0.11fF
C67304 INVX1_LOC_238/Y INVX1_LOC_229/A 0.14fF
C67305 INVX1_LOC_50/A INVX1_LOC_85/A 0.32fF
C67306 NAND2X1_LOC_357/a_36_24# NOR2X1_LOC_652/Y 0.00fF
C67307 NAND2X1_LOC_787/A NAND2X1_LOC_833/Y 0.07fF
C67308 INVX1_LOC_269/A NOR2X1_LOC_514/A 0.06fF
C67309 NAND2X1_LOC_111/a_36_24# NOR2X1_LOC_243/B 0.01fF
C67310 INVX1_LOC_59/A INVX1_LOC_136/A 0.00fF
C67311 NOR2X1_LOC_589/A NAND2X1_LOC_53/a_36_24# 0.00fF
C67312 NOR2X1_LOC_321/a_36_216# INVX1_LOC_78/A 0.00fF
C67313 INVX1_LOC_233/A NAND2X1_LOC_640/Y 0.06fF
C67314 NOR2X1_LOC_751/A INVX1_LOC_63/A 0.00fF
C67315 NAND2X1_LOC_276/Y NOR2X1_LOC_392/Y 0.07fF
C67316 INVX1_LOC_41/A INVX1_LOC_278/A 0.01fF
C67317 D_INPUT_1 INVX1_LOC_104/A 0.07fF
C67318 NAND2X1_LOC_633/Y NOR2X1_LOC_536/A 0.07fF
C67319 INVX1_LOC_35/A INVX1_LOC_63/Y 0.03fF
C67320 NAND2X1_LOC_773/Y INVX1_LOC_136/A 0.10fF
C67321 NAND2X1_LOC_807/Y NAND2X1_LOC_807/B 0.17fF
C67322 NOR2X1_LOC_160/B INVX1_LOC_43/Y 0.19fF
C67323 INVX1_LOC_233/Y INVX1_LOC_34/A 0.14fF
C67324 INVX1_LOC_46/A NOR2X1_LOC_271/Y 0.05fF
C67325 NOR2X1_LOC_508/a_36_216# NOR2X1_LOC_56/Y 0.00fF
C67326 NOR2X1_LOC_405/A NOR2X1_LOC_155/A 0.09fF
C67327 INVX1_LOC_45/A NOR2X1_LOC_636/B 0.07fF
C67328 NOR2X1_LOC_721/Y INVX1_LOC_19/A 0.07fF
C67329 INVX1_LOC_214/A INVX1_LOC_57/A 0.03fF
C67330 INVX1_LOC_11/A NAND2X1_LOC_3/a_36_24# 0.00fF
C67331 NOR2X1_LOC_15/Y NOR2X1_LOC_360/Y 3.28fF
C67332 NOR2X1_LOC_817/Y INVX1_LOC_36/A 0.44fF
C67333 NOR2X1_LOC_667/A INVX1_LOC_57/A 0.10fF
C67334 INVX1_LOC_30/Y NOR2X1_LOC_316/a_36_216# 0.00fF
C67335 NAND2X1_LOC_807/Y NOR2X1_LOC_48/B 0.11fF
C67336 NAND2X1_LOC_860/Y INVX1_LOC_181/A 0.03fF
C67337 INVX1_LOC_278/A NAND2X1_LOC_477/A 0.10fF
C67338 NOR2X1_LOC_655/B INVX1_LOC_23/A 0.01fF
C67339 INVX1_LOC_248/A INVX1_LOC_57/A 0.07fF
C67340 INPUT_0 NAND2X1_LOC_81/B 0.03fF
C67341 INVX1_LOC_298/Y INVX1_LOC_101/A 0.13fF
C67342 NAND2X1_LOC_472/Y INVX1_LOC_38/A 0.09fF
C67343 INVX1_LOC_30/Y INVX1_LOC_26/A 0.03fF
C67344 NOR2X1_LOC_356/A INVX1_LOC_32/A 0.03fF
C67345 INVX1_LOC_35/A NOR2X1_LOC_175/A 0.01fF
C67346 NOR2X1_LOC_401/a_36_216# NAND2X1_LOC_860/A 0.01fF
C67347 INVX1_LOC_37/A NOR2X1_LOC_487/Y 0.01fF
C67348 INVX1_LOC_224/Y INVX1_LOC_232/A 0.03fF
C67349 INVX1_LOC_1/A INVX1_LOC_314/Y 0.04fF
C67350 NOR2X1_LOC_456/Y NOR2X1_LOC_220/A 0.10fF
C67351 NOR2X1_LOC_590/Y INVX1_LOC_85/A 0.00fF
C67352 INVX1_LOC_139/A INVX1_LOC_179/A 0.00fF
C67353 INVX1_LOC_269/A NOR2X1_LOC_617/Y 0.02fF
C67354 D_INPUT_1 INVX1_LOC_263/A 0.05fF
C67355 NOR2X1_LOC_328/Y NOR2X1_LOC_696/a_36_216# 0.00fF
C67356 INVX1_LOC_294/Y INVX1_LOC_171/Y 0.01fF
C67357 INVX1_LOC_104/A NOR2X1_LOC_652/Y 0.10fF
C67358 INVX1_LOC_5/A NOR2X1_LOC_423/Y 0.00fF
C67359 INVX1_LOC_298/Y NOR2X1_LOC_355/A 0.05fF
C67360 INVX1_LOC_36/A NAND2X1_LOC_597/a_36_24# 0.00fF
C67361 NOR2X1_LOC_288/A NOR2X1_LOC_798/A 0.00fF
C67362 INVX1_LOC_286/Y NOR2X1_LOC_599/A 0.03fF
C67363 NAND2X1_LOC_214/B NOR2X1_LOC_84/Y 0.38fF
C67364 INVX1_LOC_290/A INVX1_LOC_271/A 0.02fF
C67365 INVX1_LOC_227/Y INVX1_LOC_292/A 0.02fF
C67366 NOR2X1_LOC_160/B INVX1_LOC_130/Y 0.03fF
C67367 INVX1_LOC_51/Y NAND2X1_LOC_206/B 0.09fF
C67368 INVX1_LOC_53/Y NOR2X1_LOC_15/a_36_216# 0.00fF
C67369 INVX1_LOC_64/A NAND2X1_LOC_350/B 0.01fF
C67370 INVX1_LOC_290/A INVX1_LOC_105/Y 0.03fF
C67371 NOR2X1_LOC_590/A INVX1_LOC_305/A 0.09fF
C67372 NOR2X1_LOC_521/Y INVX1_LOC_57/A 0.01fF
C67373 NAND2X1_LOC_860/A INVX1_LOC_53/Y 0.19fF
C67374 NOR2X1_LOC_15/Y NOR2X1_LOC_717/a_36_216# 0.00fF
C67375 NOR2X1_LOC_500/Y NOR2X1_LOC_717/A 0.18fF
C67376 INVX1_LOC_14/Y NOR2X1_LOC_831/B 0.04fF
C67377 INVX1_LOC_304/A NOR2X1_LOC_662/A 0.01fF
C67378 INVX1_LOC_225/A NAND2X1_LOC_703/Y 0.01fF
C67379 NOR2X1_LOC_595/Y INVX1_LOC_49/Y 0.01fF
C67380 NOR2X1_LOC_201/A NOR2X1_LOC_99/B 0.03fF
C67381 INVX1_LOC_64/A INVX1_LOC_208/A 0.06fF
C67382 NOR2X1_LOC_74/A INVX1_LOC_32/A 0.14fF
C67383 INVX1_LOC_5/A NOR2X1_LOC_222/Y 0.08fF
C67384 NAND2X1_LOC_348/A NOR2X1_LOC_297/A 0.01fF
C67385 NAND2X1_LOC_861/Y INVX1_LOC_181/A 0.03fF
C67386 INVX1_LOC_64/A NOR2X1_LOC_516/B 0.32fF
C67387 D_INPUT_0 NOR2X1_LOC_646/B 0.02fF
C67388 INVX1_LOC_256/A NOR2X1_LOC_537/A 0.03fF
C67389 NOR2X1_LOC_389/A NOR2X1_LOC_759/Y 0.01fF
C67390 NOR2X1_LOC_723/Y NOR2X1_LOC_722/Y 0.05fF
C67391 NOR2X1_LOC_687/Y INVX1_LOC_292/Y 0.75fF
C67392 INVX1_LOC_34/A NOR2X1_LOC_205/Y 0.00fF
C67393 NOR2X1_LOC_56/Y INVX1_LOC_19/A 0.07fF
C67394 NAND2X1_LOC_326/A NOR2X1_LOC_52/B 0.09fF
C67395 INVX1_LOC_202/A NOR2X1_LOC_389/A 0.10fF
C67396 INVX1_LOC_256/A NOR2X1_LOC_716/B 0.01fF
C67397 NOR2X1_LOC_9/Y INVX1_LOC_32/A 0.03fF
C67398 VDD NOR2X1_LOC_653/Y 0.28fF
C67399 NOR2X1_LOC_826/a_36_216# INVX1_LOC_234/A 0.00fF
C67400 NOR2X1_LOC_603/Y INVX1_LOC_186/Y 0.01fF
C67401 NAND2X1_LOC_213/A NOR2X1_LOC_156/B 0.04fF
C67402 INPUT_0 INVX1_LOC_4/Y 0.03fF
C67403 INVX1_LOC_215/A NOR2X1_LOC_109/Y 0.05fF
C67404 INVX1_LOC_266/A INVX1_LOC_149/A 0.00fF
C67405 INVX1_LOC_119/A NAND2X1_LOC_538/Y 0.02fF
C67406 INVX1_LOC_11/A NAND2X1_LOC_163/a_36_24# 0.00fF
C67407 NAND2X1_LOC_564/B INVX1_LOC_306/Y 0.05fF
C67408 INVX1_LOC_126/A INVX1_LOC_29/A 0.04fF
C67409 NAND2X1_LOC_708/Y NOR2X1_LOC_53/a_36_216# 0.00fF
C67410 NOR2X1_LOC_738/Y NOR2X1_LOC_731/A 0.05fF
C67411 INVX1_LOC_5/A INVX1_LOC_220/Y 0.01fF
C67412 VDD INVX1_LOC_19/A 1.44fF
C67413 NAND2X1_LOC_787/A NOR2X1_LOC_76/A 0.03fF
C67414 NOR2X1_LOC_778/B INVX1_LOC_1/A 0.03fF
C67415 VDD NOR2X1_LOC_11/Y 0.38fF
C67416 NOR2X1_LOC_340/Y INVX1_LOC_31/A 0.03fF
C67417 INVX1_LOC_27/A INVX1_LOC_290/A 0.17fF
C67418 INVX1_LOC_93/A NAND2X1_LOC_388/a_36_24# 0.01fF
C67419 INVX1_LOC_38/A NAND2X1_LOC_206/Y 0.01fF
C67420 NOR2X1_LOC_721/Y INVX1_LOC_26/Y 0.05fF
C67421 NAND2X1_LOC_833/Y INVX1_LOC_30/A 1.36fF
C67422 NOR2X1_LOC_860/B NOR2X1_LOC_360/Y 0.05fF
C67423 NAND2X1_LOC_549/Y INPUT_1 0.00fF
C67424 INVX1_LOC_182/A INVX1_LOC_23/A 0.07fF
C67425 NOR2X1_LOC_273/Y NOR2X1_LOC_596/A 0.12fF
C67426 NOR2X1_LOC_117/Y INVX1_LOC_54/A 0.10fF
C67427 INVX1_LOC_225/Y INVX1_LOC_177/A 0.00fF
C67428 INVX1_LOC_36/A NOR2X1_LOC_570/B 0.02fF
C67429 INVX1_LOC_6/A NOR2X1_LOC_438/Y 0.03fF
C67430 NAND2X1_LOC_562/B NAND2X1_LOC_577/A 0.22fF
C67431 INVX1_LOC_62/A INVX1_LOC_38/Y 0.01fF
C67432 NAND2X1_LOC_51/B INVX1_LOC_57/A 0.10fF
C67433 INVX1_LOC_292/A INVX1_LOC_111/Y 0.08fF
C67434 NOR2X1_LOC_837/a_36_216# NOR2X1_LOC_837/Y 0.02fF
C67435 NOR2X1_LOC_778/B NOR2X1_LOC_794/B 0.04fF
C67436 NAND2X1_LOC_483/Y INVX1_LOC_217/A 0.02fF
C67437 INVX1_LOC_239/A NOR2X1_LOC_459/A 0.18fF
C67438 INVX1_LOC_232/Y INVX1_LOC_230/Y 0.01fF
C67439 NOR2X1_LOC_791/Y NOR2X1_LOC_76/A 0.01fF
C67440 INPUT_1 NOR2X1_LOC_291/Y 0.14fF
C67441 INVX1_LOC_265/A INVX1_LOC_18/A 0.03fF
C67442 NOR2X1_LOC_103/Y INVX1_LOC_232/A 0.10fF
C67443 NOR2X1_LOC_655/B INVX1_LOC_31/A 0.13fF
C67444 INVX1_LOC_24/A NOR2X1_LOC_172/Y 0.03fF
C67445 INVX1_LOC_174/A NAND2X1_LOC_452/a_36_24# 0.01fF
C67446 NOR2X1_LOC_837/Y NOR2X1_LOC_852/B 0.03fF
C67447 NOR2X1_LOC_186/Y NAND2X1_LOC_842/B 0.02fF
C67448 NOR2X1_LOC_445/Y INVX1_LOC_94/A 0.00fF
C67449 INVX1_LOC_18/A NOR2X1_LOC_180/Y 0.03fF
C67450 INVX1_LOC_11/A INVX1_LOC_174/Y 0.01fF
C67451 INVX1_LOC_245/A NOR2X1_LOC_471/Y 0.04fF
C67452 NAND2X1_LOC_361/Y INVX1_LOC_77/A 0.12fF
C67453 NOR2X1_LOC_208/Y NOR2X1_LOC_570/B 0.28fF
C67454 INVX1_LOC_93/A INVX1_LOC_28/A 0.38fF
C67455 NOR2X1_LOC_383/Y NOR2X1_LOC_103/Y 0.02fF
C67456 INVX1_LOC_41/A NOR2X1_LOC_262/Y 0.02fF
C67457 NAND2X1_LOC_555/Y NAND2X1_LOC_671/a_36_24# 0.00fF
C67458 NAND2X1_LOC_79/Y NOR2X1_LOC_124/B 0.16fF
C67459 INVX1_LOC_24/A NOR2X1_LOC_392/B 0.06fF
C67460 D_INPUT_1 INVX1_LOC_206/Y 0.06fF
C67461 NOR2X1_LOC_124/A INVX1_LOC_26/A 0.02fF
C67462 INVX1_LOC_174/A NOR2X1_LOC_764/a_36_216# 0.00fF
C67463 NAND2X1_LOC_739/B INVX1_LOC_240/A 0.03fF
C67464 NOR2X1_LOC_632/Y NOR2X1_LOC_471/Y 0.02fF
C67465 NOR2X1_LOC_91/A INVX1_LOC_291/Y 0.03fF
C67466 NOR2X1_LOC_218/A NOR2X1_LOC_561/Y 0.02fF
C67467 INVX1_LOC_69/Y INVX1_LOC_58/Y 0.09fF
C67468 NOR2X1_LOC_558/a_36_216# INVX1_LOC_47/Y 0.02fF
C67469 NAND2X1_LOC_303/Y INVX1_LOC_173/Y 0.04fF
C67470 NAND2X1_LOC_483/Y NAND2X1_LOC_787/B 0.12fF
C67471 NOR2X1_LOC_807/B NOR2X1_LOC_326/Y 0.02fF
C67472 INVX1_LOC_1/A NOR2X1_LOC_724/Y 0.07fF
C67473 NOR2X1_LOC_772/Y NOR2X1_LOC_557/Y 0.23fF
C67474 NOR2X1_LOC_454/Y NAND2X1_LOC_654/B 0.15fF
C67475 NOR2X1_LOC_607/Y INVX1_LOC_104/A 0.10fF
C67476 INVX1_LOC_279/A NOR2X1_LOC_276/Y 0.01fF
C67477 INVX1_LOC_48/Y NOR2X1_LOC_19/B 0.00fF
C67478 NAND2X1_LOC_540/a_36_24# INPUT_0 0.01fF
C67479 INVX1_LOC_29/A NOR2X1_LOC_600/a_36_216# 0.00fF
C67480 NOR2X1_LOC_831/B NOR2X1_LOC_831/Y 0.05fF
C67481 INVX1_LOC_133/A NAND2X1_LOC_288/A 0.21fF
C67482 NAND2X1_LOC_807/B INVX1_LOC_131/Y 0.03fF
C67483 NOR2X1_LOC_568/A INVX1_LOC_232/A 0.06fF
C67484 NOR2X1_LOC_655/B INVX1_LOC_111/A 0.45fF
C67485 NOR2X1_LOC_392/B NOR2X1_LOC_557/Y 0.10fF
C67486 NOR2X1_LOC_319/B NOR2X1_LOC_855/A 0.02fF
C67487 NOR2X1_LOC_299/Y NOR2X1_LOC_380/a_36_216# 0.02fF
C67488 NAND2X1_LOC_802/A NAND2X1_LOC_799/a_36_24# 0.00fF
C67489 INVX1_LOC_166/A NAND2X1_LOC_659/B 0.07fF
C67490 NOR2X1_LOC_769/A INVX1_LOC_268/Y 0.01fF
C67491 NOR2X1_LOC_751/Y INVX1_LOC_1/Y 0.02fF
C67492 NOR2X1_LOC_703/B INVX1_LOC_22/A 0.03fF
C67493 INVX1_LOC_63/Y NOR2X1_LOC_365/a_36_216# 0.00fF
C67494 NOR2X1_LOC_155/A INVX1_LOC_109/Y 0.08fF
C67495 NOR2X1_LOC_255/Y NOR2X1_LOC_124/A 0.01fF
C67496 INVX1_LOC_292/A NOR2X1_LOC_137/A 0.00fF
C67497 NAND2X1_LOC_303/Y NOR2X1_LOC_385/Y 0.22fF
C67498 D_INPUT_1 NAND2X1_LOC_674/a_36_24# 0.00fF
C67499 VDD INVX1_LOC_26/Y 1.41fF
C67500 NAND2X1_LOC_96/A INVX1_LOC_78/A 0.19fF
C67501 NOR2X1_LOC_616/Y NOR2X1_LOC_617/Y 0.04fF
C67502 NAND2X1_LOC_9/Y NAND2X1_LOC_642/Y 0.02fF
C67503 INVX1_LOC_31/A NOR2X1_LOC_99/B 0.07fF
C67504 NOR2X1_LOC_364/Y NOR2X1_LOC_367/B 0.09fF
C67505 INVX1_LOC_141/Y NAND2X1_LOC_808/A 0.03fF
C67506 INVX1_LOC_60/Y INVX1_LOC_8/A 0.16fF
C67507 NAND2X1_LOC_721/A NOR2X1_LOC_693/Y 0.07fF
C67508 NAND2X1_LOC_722/A NAND2X1_LOC_833/Y 0.25fF
C67509 INVX1_LOC_153/Y INVX1_LOC_266/Y 0.10fF
C67510 INVX1_LOC_300/Y NAND2X1_LOC_863/B 0.15fF
C67511 INVX1_LOC_245/Y INVX1_LOC_55/Y 0.04fF
C67512 NOR2X1_LOC_89/A NAND2X1_LOC_572/B 0.28fF
C67513 INVX1_LOC_7/Y INVX1_LOC_123/A 0.02fF
C67514 INVX1_LOC_136/A INVX1_LOC_279/A 0.07fF
C67515 NOR2X1_LOC_441/Y INVX1_LOC_313/A 0.03fF
C67516 INVX1_LOC_166/A VDD 0.12fF
C67517 NOR2X1_LOC_91/A NOR2X1_LOC_176/Y 0.01fF
C67518 INVX1_LOC_31/A NOR2X1_LOC_846/B 0.01fF
C67519 NOR2X1_LOC_351/Y NOR2X1_LOC_334/Y 0.01fF
C67520 NAND2X1_LOC_337/B NOR2X1_LOC_329/B 0.21fF
C67521 NAND2X1_LOC_557/Y VDD 0.00fF
C67522 NOR2X1_LOC_816/A NOR2X1_LOC_329/B 0.07fF
C67523 NOR2X1_LOC_849/a_36_216# NOR2X1_LOC_99/B 0.01fF
C67524 INVX1_LOC_30/A NOR2X1_LOC_76/A 0.10fF
C67525 INVX1_LOC_133/A INVX1_LOC_19/A 0.01fF
C67526 INVX1_LOC_157/Y NAND2X1_LOC_454/Y -0.06fF
C67527 NOR2X1_LOC_598/B NOR2X1_LOC_857/A 0.10fF
C67528 NOR2X1_LOC_392/B INVX1_LOC_143/A 0.01fF
C67529 INVX1_LOC_38/A NOR2X1_LOC_639/Y 0.02fF
C67530 NAND2X1_LOC_81/B NOR2X1_LOC_84/B 0.03fF
C67531 NOR2X1_LOC_441/Y NAND2X1_LOC_807/Y 0.07fF
C67532 NOR2X1_LOC_180/B INVX1_LOC_30/A 0.19fF
C67533 NOR2X1_LOC_635/A NAND2X1_LOC_451/Y 0.13fF
C67534 INVX1_LOC_182/Y NOR2X1_LOC_276/Y 0.00fF
C67535 NOR2X1_LOC_431/Y NOR2X1_LOC_561/Y 0.04fF
C67536 INVX1_LOC_177/A INVX1_LOC_266/Y 0.04fF
C67537 NAND2X1_LOC_550/A INVX1_LOC_282/A 0.07fF
C67538 INVX1_LOC_166/A NAND2X1_LOC_463/a_36_24# 0.01fF
C67539 INVX1_LOC_58/A INVX1_LOC_117/A 0.00fF
C67540 INVX1_LOC_5/A NOR2X1_LOC_69/A 0.03fF
C67541 NOR2X1_LOC_381/a_36_216# INVX1_LOC_31/A 0.01fF
C67542 NOR2X1_LOC_13/Y INVX1_LOC_10/A 0.97fF
C67543 NAND2X1_LOC_574/A INVX1_LOC_15/A 0.02fF
C67544 INVX1_LOC_64/A NAND2X1_LOC_211/Y 0.01fF
C67545 NOR2X1_LOC_282/Y INVX1_LOC_118/A 0.02fF
C67546 NAND2X1_LOC_656/A NOR2X1_LOC_332/A 0.12fF
C67547 NOR2X1_LOC_321/Y NOR2X1_LOC_45/B 0.45fF
C67548 NOR2X1_LOC_716/B NOR2X1_LOC_397/a_36_216# 0.01fF
C67549 NOR2X1_LOC_435/B INVX1_LOC_15/A 0.06fF
C67550 NOR2X1_LOC_263/a_36_216# NOR2X1_LOC_773/Y 0.00fF
C67551 INVX1_LOC_1/A NOR2X1_LOC_557/A 0.01fF
C67552 NAND2X1_LOC_36/A NOR2X1_LOC_163/Y 0.12fF
C67553 NOR2X1_LOC_637/a_36_216# NOR2X1_LOC_561/Y 0.01fF
C67554 NOR2X1_LOC_662/A INVX1_LOC_19/Y 0.01fF
C67555 NOR2X1_LOC_536/A NOR2X1_LOC_591/A 0.04fF
C67556 NOR2X1_LOC_373/Y NOR2X1_LOC_237/Y 0.43fF
C67557 INVX1_LOC_73/A INVX1_LOC_30/A 0.01fF
C67558 NOR2X1_LOC_553/Y INVX1_LOC_104/A 0.07fF
C67559 INVX1_LOC_90/A INVX1_LOC_24/A 0.30fF
C67560 INVX1_LOC_270/A INVX1_LOC_54/A 0.14fF
C67561 INVX1_LOC_88/A NOR2X1_LOC_139/Y 0.45fF
C67562 INVX1_LOC_136/A INVX1_LOC_182/Y 0.03fF
C67563 INVX1_LOC_230/Y NOR2X1_LOC_391/Y 0.02fF
C67564 NOR2X1_LOC_413/a_36_216# INVX1_LOC_234/A 0.00fF
C67565 NOR2X1_LOC_172/Y NOR2X1_LOC_130/A 0.03fF
C67566 NAND2X1_LOC_852/Y NOR2X1_LOC_505/Y 0.00fF
C67567 NOR2X1_LOC_441/Y INVX1_LOC_6/A 0.05fF
C67568 INVX1_LOC_54/Y INVX1_LOC_16/A 0.07fF
C67569 INVX1_LOC_207/A NOR2X1_LOC_576/B 0.19fF
C67570 NAND2X1_LOC_854/B NOR2X1_LOC_591/Y 0.06fF
C67571 NAND2X1_LOC_223/A NAND2X1_LOC_206/Y 0.07fF
C67572 INVX1_LOC_88/A NAND2X1_LOC_468/B 0.01fF
C67573 NOR2X1_LOC_646/B INVX1_LOC_46/Y 0.39fF
C67574 NOR2X1_LOC_629/a_36_216# INVX1_LOC_234/A 0.00fF
C67575 INVX1_LOC_215/A NAND2X1_LOC_112/a_36_24# 0.00fF
C67576 NOR2X1_LOC_602/B NOR2X1_LOC_109/Y 0.03fF
C67577 INVX1_LOC_150/Y NAND2X1_LOC_107/a_36_24# 0.01fF
C67578 INVX1_LOC_90/A NOR2X1_LOC_557/Y 0.05fF
C67579 INVX1_LOC_234/A NOR2X1_LOC_84/Y 0.19fF
C67580 INVX1_LOC_278/Y NAND2X1_LOC_170/A 0.03fF
C67581 INVX1_LOC_36/A INVX1_LOC_286/A 0.17fF
C67582 NAND2X1_LOC_553/A NOR2X1_LOC_271/Y 0.08fF
C67583 NOR2X1_LOC_38/B NAND2X1_LOC_74/B 0.08fF
C67584 NOR2X1_LOC_504/Y INVX1_LOC_10/A 0.16fF
C67585 INVX1_LOC_49/A NOR2X1_LOC_564/Y 0.04fF
C67586 NOR2X1_LOC_389/B NOR2X1_LOC_557/Y 0.19fF
C67587 INVX1_LOC_17/A NAND2X1_LOC_1/Y 1.24fF
C67588 NOR2X1_LOC_561/Y NOR2X1_LOC_131/A 0.03fF
C67589 INVX1_LOC_54/A NOR2X1_LOC_109/Y 0.07fF
C67590 NOR2X1_LOC_315/Y NAND2X1_LOC_861/Y 0.01fF
C67591 INVX1_LOC_45/A INVX1_LOC_186/A 0.07fF
C67592 NOR2X1_LOC_717/A INVX1_LOC_307/A 0.02fF
C67593 INVX1_LOC_94/A NOR2X1_LOC_335/B 0.12fF
C67594 NOR2X1_LOC_504/Y NOR2X1_LOC_504/a_36_216# 0.01fF
C67595 INVX1_LOC_118/A NOR2X1_LOC_291/Y 0.31fF
C67596 INVX1_LOC_161/Y NOR2X1_LOC_136/a_36_216# 0.01fF
C67597 INVX1_LOC_89/A NOR2X1_LOC_709/A 0.92fF
C67598 NOR2X1_LOC_589/A NOR2X1_LOC_229/Y 0.43fF
C67599 INVX1_LOC_256/A NOR2X1_LOC_567/a_36_216# 0.01fF
C67600 INVX1_LOC_314/Y NOR2X1_LOC_188/A 0.10fF
C67601 NOR2X1_LOC_259/B NOR2X1_LOC_342/A 0.06fF
C67602 NOR2X1_LOC_592/A NAND2X1_LOC_453/A -0.00fF
C67603 INVX1_LOC_79/A NOR2X1_LOC_577/Y 0.01fF
C67604 NOR2X1_LOC_274/B INVX1_LOC_91/A 0.03fF
C67605 INVX1_LOC_72/A NOR2X1_LOC_78/A 0.13fF
C67606 INVX1_LOC_314/Y NOR2X1_LOC_548/B 0.10fF
C67607 NOR2X1_LOC_700/Y NAND2X1_LOC_852/Y 0.10fF
C67608 INVX1_LOC_161/Y VDD 1.97fF
C67609 NOR2X1_LOC_644/Y INVX1_LOC_313/Y 0.01fF
C67610 NOR2X1_LOC_433/A NOR2X1_LOC_815/A 0.02fF
C67611 INVX1_LOC_36/A INVX1_LOC_95/A 0.03fF
C67612 INVX1_LOC_153/Y INVX1_LOC_42/Y 0.34fF
C67613 INVX1_LOC_161/Y NAND2X1_LOC_800/A 0.02fF
C67614 NAND2X1_LOC_35/Y NOR2X1_LOC_88/Y 0.07fF
C67615 INVX1_LOC_21/A INVX1_LOC_274/A 0.04fF
C67616 INVX1_LOC_90/A INVX1_LOC_143/A 0.08fF
C67617 NOR2X1_LOC_479/B INVX1_LOC_135/A 0.08fF
C67618 NAND2X1_LOC_781/a_36_24# INVX1_LOC_275/Y 0.00fF
C67619 INVX1_LOC_45/A NAND2X1_LOC_447/Y 0.01fF
C67620 NOR2X1_LOC_738/Y INVX1_LOC_117/A 0.01fF
C67621 NAND2X1_LOC_583/a_36_24# NAND2X1_LOC_639/A 0.00fF
C67622 INVX1_LOC_41/A NOR2X1_LOC_728/a_36_216# 0.00fF
C67623 INVX1_LOC_45/Y NOR2X1_LOC_318/B 0.01fF
C67624 NOR2X1_LOC_267/A INVX1_LOC_95/A 0.09fF
C67625 NOR2X1_LOC_568/A NAND2X1_LOC_447/Y 0.50fF
C67626 NOR2X1_LOC_843/A INPUT_0 0.03fF
C67627 NOR2X1_LOC_19/B INVX1_LOC_216/A 0.04fF
C67628 NOR2X1_LOC_478/A INVX1_LOC_37/A 0.02fF
C67629 INVX1_LOC_13/A D_INPUT_0 1.74fF
C67630 NAND2X1_LOC_99/A INVX1_LOC_42/A 0.01fF
C67631 NOR2X1_LOC_142/Y INVX1_LOC_6/A 0.20fF
C67632 INVX1_LOC_312/A VDD 0.00fF
C67633 NAND2X1_LOC_35/Y INVX1_LOC_84/A 0.07fF
C67634 NAND2X1_LOC_16/a_36_24# NAND2X1_LOC_39/Y 0.00fF
C67635 NOR2X1_LOC_810/A NOR2X1_LOC_326/Y 0.00fF
C67636 NOR2X1_LOC_599/A VDD 0.16fF
C67637 NOR2X1_LOC_577/Y INVX1_LOC_91/A 0.07fF
C67638 INVX1_LOC_18/A NOR2X1_LOC_603/Y 0.06fF
C67639 NOR2X1_LOC_383/Y NOR2X1_LOC_123/B 0.00fF
C67640 NOR2X1_LOC_379/Y INVX1_LOC_91/A 0.01fF
C67641 INVX1_LOC_50/A INVX1_LOC_290/Y 0.75fF
C67642 NOR2X1_LOC_817/Y NOR2X1_LOC_656/Y 0.01fF
C67643 NOR2X1_LOC_273/Y NAND2X1_LOC_469/B 0.24fF
C67644 INVX1_LOC_48/Y NOR2X1_LOC_216/B 0.09fF
C67645 NOR2X1_LOC_309/Y INVX1_LOC_286/A 0.01fF
C67646 NOR2X1_LOC_596/Y NOR2X1_LOC_331/B 0.00fF
C67647 NOR2X1_LOC_759/Y NAND2X1_LOC_469/B 0.94fF
C67648 INVX1_LOC_71/A NAND2X1_LOC_447/Y 0.01fF
C67649 INVX1_LOC_285/Y INVX1_LOC_266/Y 0.00fF
C67650 NAND2X1_LOC_776/a_36_24# NAND2X1_LOC_804/Y 0.01fF
C67651 NOR2X1_LOC_91/Y INVX1_LOC_46/A 0.00fF
C67652 INVX1_LOC_12/A NOR2X1_LOC_717/A 0.07fF
C67653 NOR2X1_LOC_68/A INVX1_LOC_37/A 4.37fF
C67654 NOR2X1_LOC_246/A D_INPUT_0 0.47fF
C67655 INVX1_LOC_64/A NAND2X1_LOC_81/a_36_24# -0.00fF
C67656 NOR2X1_LOC_68/A NOR2X1_LOC_231/A 0.02fF
C67657 NOR2X1_LOC_303/Y NOR2X1_LOC_35/Y 0.11fF
C67658 NOR2X1_LOC_589/A NAND2X1_LOC_850/A 0.10fF
C67659 NOR2X1_LOC_629/B INVX1_LOC_91/A 0.06fF
C67660 NAND2X1_LOC_783/A INVX1_LOC_90/A 0.01fF
C67661 INVX1_LOC_135/A NOR2X1_LOC_130/a_36_216# 0.01fF
C67662 NOR2X1_LOC_655/B INVX1_LOC_6/A 0.05fF
C67663 NOR2X1_LOC_81/a_36_216# INVX1_LOC_46/A 0.00fF
C67664 NOR2X1_LOC_361/B NAND2X1_LOC_288/A 0.29fF
C67665 NOR2X1_LOC_273/Y NAND2X1_LOC_212/a_36_24# 0.01fF
C67666 INVX1_LOC_53/A NOR2X1_LOC_640/B 0.21fF
C67667 INPUT_0 NAND2X1_LOC_862/A 0.01fF
C67668 INVX1_LOC_90/A NOR2X1_LOC_130/A 0.06fF
C67669 NOR2X1_LOC_510/Y INVX1_LOC_19/A 0.07fF
C67670 NAND2X1_LOC_214/Y NOR2X1_LOC_673/A 0.02fF
C67671 INVX1_LOC_58/A INVX1_LOC_3/Y 0.02fF
C67672 NOR2X1_LOC_437/Y VDD -0.00fF
C67673 NOR2X1_LOC_751/A INVX1_LOC_1/Y 0.00fF
C67674 NOR2X1_LOC_553/B INVX1_LOC_75/A 0.03fF
C67675 INVX1_LOC_14/A NAND2X1_LOC_659/A 0.13fF
C67676 NOR2X1_LOC_230/a_36_216# INVX1_LOC_54/A 0.00fF
C67677 NOR2X1_LOC_309/Y INVX1_LOC_95/A 0.05fF
C67678 NOR2X1_LOC_718/B NOR2X1_LOC_486/Y 0.07fF
C67679 INVX1_LOC_64/A NAND2X1_LOC_791/a_36_24# 0.00fF
C67680 NOR2X1_LOC_78/A NOR2X1_LOC_537/Y 0.04fF
C67681 NOR2X1_LOC_272/Y INVX1_LOC_29/A 0.03fF
C67682 NAND2X1_LOC_338/B NOR2X1_LOC_78/A 0.07fF
C67683 NOR2X1_LOC_334/Y NOR2X1_LOC_748/A 0.10fF
C67684 INVX1_LOC_36/A INVX1_LOC_54/A 3.23fF
C67685 NOR2X1_LOC_48/B NOR2X1_LOC_109/Y 1.60fF
C67686 INVX1_LOC_57/A NOR2X1_LOC_248/A 0.01fF
C67687 NOR2X1_LOC_364/Y INVX1_LOC_76/A 0.02fF
C67688 NOR2X1_LOC_320/Y NAND2X1_LOC_660/Y 0.18fF
C67689 INVX1_LOC_141/Y INVX1_LOC_92/A 0.03fF
C67690 D_INPUT_6 NOR2X1_LOC_1/Y 0.02fF
C67691 INVX1_LOC_24/A INVX1_LOC_38/A 0.73fF
C67692 NAND2X1_LOC_323/B NOR2X1_LOC_78/A 0.03fF
C67693 NAND2X1_LOC_347/B NAND2X1_LOC_63/Y 1.09fF
C67694 INVX1_LOC_27/A INVX1_LOC_114/Y 0.00fF
C67695 NAND2X1_LOC_348/A NOR2X1_LOC_130/A 0.02fF
C67696 INVX1_LOC_69/Y NOR2X1_LOC_501/a_36_216# 0.01fF
C67697 NOR2X1_LOC_190/a_36_216# INVX1_LOC_93/Y 0.01fF
C67698 NAND2X1_LOC_35/Y INVX1_LOC_15/A 0.07fF
C67699 NOR2X1_LOC_817/Y INVX1_LOC_63/A 0.20fF
C67700 NOR2X1_LOC_660/Y NOR2X1_LOC_38/B 0.02fF
C67701 NAND2X1_LOC_222/B NAND2X1_LOC_219/B 0.06fF
C67702 GATE_811 INVX1_LOC_46/A 0.04fF
C67703 NOR2X1_LOC_361/B INVX1_LOC_19/A 0.03fF
C67704 NOR2X1_LOC_514/Y D_INPUT_3 0.03fF
C67705 INVX1_LOC_33/A NAND2X1_LOC_472/Y 0.09fF
C67706 NAND2X1_LOC_700/a_36_24# NAND2X1_LOC_782/B 0.01fF
C67707 NOR2X1_LOC_468/Y NAND2X1_LOC_74/B 0.18fF
C67708 INVX1_LOC_22/A INVX1_LOC_91/A 0.29fF
C67709 NOR2X1_LOC_353/Y NOR2X1_LOC_35/Y 0.01fF
C67710 NOR2X1_LOC_557/Y NOR2X1_LOC_561/A 0.15fF
C67711 NOR2X1_LOC_208/Y INVX1_LOC_54/A 0.03fF
C67712 INVX1_LOC_24/A NOR2X1_LOC_51/A 0.03fF
C67713 NAND2X1_LOC_338/B NAND2X1_LOC_464/A 0.10fF
C67714 INVX1_LOC_161/Y INVX1_LOC_133/A 0.01fF
C67715 GATE_811 NOR2X1_LOC_766/Y 0.00fF
C67716 INVX1_LOC_11/Y INVX1_LOC_22/A 0.13fF
C67717 INVX1_LOC_27/A NOR2X1_LOC_467/A 0.10fF
C67718 NAND2X1_LOC_361/Y INVX1_LOC_9/A 0.33fF
C67719 D_INPUT_4 INVX1_LOC_140/A 0.02fF
C67720 NOR2X1_LOC_546/B INVX1_LOC_92/A 0.04fF
C67721 INVX1_LOC_120/A INVX1_LOC_48/A 0.53fF
C67722 NOR2X1_LOC_220/B INVX1_LOC_4/Y 0.09fF
C67723 NOR2X1_LOC_45/B NOR2X1_LOC_686/B 0.03fF
C67724 INVX1_LOC_316/Y INVX1_LOC_20/A 0.01fF
C67725 NOR2X1_LOC_416/A NAND2X1_LOC_215/A 0.54fF
C67726 NOR2X1_LOC_75/Y NOR2X1_LOC_89/A 0.00fF
C67727 NOR2X1_LOC_721/A NAND2X1_LOC_96/A 0.03fF
C67728 INVX1_LOC_218/A NAND2X1_LOC_642/a_36_24# 0.00fF
C67729 INVX1_LOC_275/A INVX1_LOC_92/A 0.58fF
C67730 INVX1_LOC_150/Y NOR2X1_LOC_114/Y 0.01fF
C67731 NOR2X1_LOC_309/Y INVX1_LOC_54/A 0.28fF
C67732 INVX1_LOC_94/A INVX1_LOC_84/A 0.16fF
C67733 INVX1_LOC_143/A INVX1_LOC_38/A 0.07fF
C67734 NOR2X1_LOC_658/Y INVX1_LOC_12/A 0.10fF
C67735 NOR2X1_LOC_543/A INVX1_LOC_46/A 0.01fF
C67736 NOR2X1_LOC_464/B INVX1_LOC_78/A 0.04fF
C67737 NAND2X1_LOC_842/B NAND2X1_LOC_642/Y 0.05fF
C67738 INVX1_LOC_36/A NAND2X1_LOC_807/B 0.05fF
C67739 NAND2X1_LOC_364/A INVX1_LOC_29/A 0.12fF
C67740 INVX1_LOC_25/A NAND2X1_LOC_214/B 0.10fF
C67741 NOR2X1_LOC_128/B D_INPUT_3 0.00fF
C67742 NOR2X1_LOC_124/B INVX1_LOC_123/Y 0.26fF
C67743 NOR2X1_LOC_15/Y INVX1_LOC_26/A 0.07fF
C67744 INVX1_LOC_62/Y NAND2X1_LOC_74/B 0.03fF
C67745 INVX1_LOC_62/A VDD 0.12fF
C67746 INVX1_LOC_36/A NOR2X1_LOC_48/B 0.03fF
C67747 INVX1_LOC_225/Y INVX1_LOC_4/Y 0.10fF
C67748 NOR2X1_LOC_84/Y NOR2X1_LOC_216/B 0.00fF
C67749 INVX1_LOC_140/A INPUT_4 0.07fF
C67750 NOR2X1_LOC_91/A NAND2X1_LOC_579/A 0.09fF
C67751 INVX1_LOC_31/A NOR2X1_LOC_28/a_36_216# 0.01fF
C67752 INVX1_LOC_35/A INVX1_LOC_5/A 1.40fF
C67753 NOR2X1_LOC_250/Y NAND2X1_LOC_175/Y 0.03fF
C67754 INVX1_LOC_25/A INVX1_LOC_27/A 0.66fF
C67755 INVX1_LOC_124/Y INVX1_LOC_32/A 0.32fF
C67756 NOR2X1_LOC_557/A NOR2X1_LOC_188/A 0.17fF
C67757 NOR2X1_LOC_71/Y NAND2X1_LOC_721/A 0.03fF
C67758 NAND2X1_LOC_729/B NAND2X1_LOC_856/a_36_24# 0.00fF
C67759 NOR2X1_LOC_13/Y INVX1_LOC_12/A 0.16fF
C67760 INVX1_LOC_135/A INVX1_LOC_33/Y 0.01fF
C67761 NOR2X1_LOC_557/A NOR2X1_LOC_548/B 0.10fF
C67762 INVX1_LOC_33/A NAND2X1_LOC_773/B 0.07fF
C67763 NOR2X1_LOC_163/A INVX1_LOC_37/A 0.01fF
C67764 INVX1_LOC_39/A NAND2X1_LOC_549/Y 0.00fF
C67765 NOR2X1_LOC_750/A INVX1_LOC_2/Y 0.02fF
C67766 NOR2X1_LOC_789/a_36_216# INVX1_LOC_9/A 0.00fF
C67767 NAND2X1_LOC_656/A INVX1_LOC_42/A 0.98fF
C67768 NAND2X1_LOC_740/Y NAND2X1_LOC_725/A 0.03fF
C67769 D_INPUT_1 NOR2X1_LOC_92/Y 0.02fF
C67770 NAND2X1_LOC_783/A INVX1_LOC_38/A 0.01fF
C67771 NOR2X1_LOC_368/A NOR2X1_LOC_124/A 0.01fF
C67772 NOR2X1_LOC_772/B INVX1_LOC_13/Y 0.07fF
C67773 NOR2X1_LOC_419/Y NOR2X1_LOC_89/A 0.03fF
C67774 INVX1_LOC_219/A INVX1_LOC_280/A 0.03fF
C67775 NOR2X1_LOC_366/Y NOR2X1_LOC_331/B 0.02fF
C67776 NOR2X1_LOC_246/A NAND2X1_LOC_848/A 0.01fF
C67777 NOR2X1_LOC_750/a_36_216# INVX1_LOC_2/Y 0.00fF
C67778 NOR2X1_LOC_130/A INVX1_LOC_38/A 0.06fF
C67779 INVX1_LOC_136/A NOR2X1_LOC_38/B 0.00fF
C67780 INVX1_LOC_11/A NOR2X1_LOC_654/A 0.03fF
C67781 NOR2X1_LOC_716/B NOR2X1_LOC_89/A 0.17fF
C67782 NOR2X1_LOC_140/A NOR2X1_LOC_392/Y 0.02fF
C67783 NAND2X1_LOC_175/B INVX1_LOC_12/A 0.15fF
C67784 NOR2X1_LOC_130/a_36_216# INVX1_LOC_280/A 0.01fF
C67785 INVX1_LOC_16/A INVX1_LOC_35/Y 0.08fF
C67786 INVX1_LOC_13/A INVX1_LOC_46/Y 0.04fF
C67787 INVX1_LOC_226/Y NAND2X1_LOC_85/Y 0.01fF
C67788 INVX1_LOC_80/Y NAND2X1_LOC_82/Y 0.07fF
C67789 INVX1_LOC_21/A INVX1_LOC_306/Y 0.03fF
C67790 NOR2X1_LOC_391/A NAND2X1_LOC_93/B 0.02fF
C67791 NOR2X1_LOC_570/a_36_216# NOR2X1_LOC_334/Y 0.00fF
C67792 INVX1_LOC_292/A NOR2X1_LOC_383/B 1.59fF
C67793 INVX1_LOC_177/A INVX1_LOC_19/A 0.06fF
C67794 NOR2X1_LOC_68/A NAND2X1_LOC_72/B 0.03fF
C67795 INVX1_LOC_2/A INVX1_LOC_264/A 0.01fF
C67796 NAND2X1_LOC_656/Y INVX1_LOC_92/A 0.25fF
C67797 INVX1_LOC_11/A INVX1_LOC_58/Y 0.11fF
C67798 NOR2X1_LOC_309/Y NAND2X1_LOC_807/B 0.40fF
C67799 NOR2X1_LOC_595/Y NAND2X1_LOC_649/B 0.06fF
C67800 NAND2X1_LOC_198/B NAND2X1_LOC_454/Y 0.01fF
C67801 NOR2X1_LOC_285/a_36_216# NOR2X1_LOC_160/B 0.02fF
C67802 NAND2X1_LOC_214/B INVX1_LOC_1/A 0.10fF
C67803 INVX1_LOC_298/Y NAND2X1_LOC_364/A 0.04fF
C67804 NOR2X1_LOC_92/Y NOR2X1_LOC_652/Y 0.01fF
C67805 NOR2X1_LOC_577/Y INVX1_LOC_231/A 0.00fF
C67806 NAND2X1_LOC_573/A NAND2X1_LOC_288/A 0.23fF
C67807 NOR2X1_LOC_526/a_36_216# INVX1_LOC_20/A 0.00fF
C67808 INVX1_LOC_24/A NAND2X1_LOC_223/A 0.03fF
C67809 NOR2X1_LOC_504/Y INVX1_LOC_12/A 0.14fF
C67810 INVX1_LOC_40/A NAND2X1_LOC_773/B 0.03fF
C67811 NOR2X1_LOC_530/Y NOR2X1_LOC_392/Y 0.00fF
C67812 INVX1_LOC_35/A NAND2X1_LOC_337/B 0.38fF
C67813 INVX1_LOC_165/Y NAND2X1_LOC_773/B 0.01fF
C67814 INVX1_LOC_158/Y NAND2X1_LOC_96/A 0.06fF
C67815 INVX1_LOC_36/A NAND2X1_LOC_215/A 0.07fF
C67816 NOR2X1_LOC_391/A INVX1_LOC_3/A 0.03fF
C67817 INVX1_LOC_27/A INVX1_LOC_1/A 0.24fF
C67818 NAND2X1_LOC_638/Y INVX1_LOC_92/A 0.07fF
C67819 INVX1_LOC_196/Y NOR2X1_LOC_809/B 0.24fF
C67820 INVX1_LOC_141/Y INVX1_LOC_53/A 0.03fF
C67821 INVX1_LOC_49/A NOR2X1_LOC_158/Y 0.07fF
C67822 INVX1_LOC_90/A NOR2X1_LOC_197/B 0.02fF
C67823 NOR2X1_LOC_848/Y NOR2X1_LOC_846/A 0.19fF
C67824 NOR2X1_LOC_757/Y NOR2X1_LOC_89/A 0.34fF
C67825 INVX1_LOC_24/A NAND2X1_LOC_256/a_36_24# 0.00fF
C67826 NOR2X1_LOC_65/B NAND2X1_LOC_656/A 0.69fF
C67827 NOR2X1_LOC_780/B NOR2X1_LOC_779/Y 0.01fF
C67828 NOR2X1_LOC_15/Y NOR2X1_LOC_666/A 0.02fF
C67829 NOR2X1_LOC_510/Y INVX1_LOC_161/Y 0.02fF
C67830 NOR2X1_LOC_441/Y NOR2X1_LOC_109/Y 0.02fF
C67831 NOR2X1_LOC_237/Y NOR2X1_LOC_438/Y 0.01fF
C67832 INVX1_LOC_28/A INVX1_LOC_35/Y 0.11fF
C67833 NOR2X1_LOC_447/Y NOR2X1_LOC_447/A 0.14fF
C67834 D_INPUT_0 NAND2X1_LOC_489/Y 0.07fF
C67835 NOR2X1_LOC_5/a_36_216# NAND2X1_LOC_574/A 0.01fF
C67836 NOR2X1_LOC_346/Y NOR2X1_LOC_360/A 0.00fF
C67837 NAND2X1_LOC_364/A NOR2X1_LOC_843/a_36_216# 0.00fF
C67838 NAND2X1_LOC_573/A INVX1_LOC_19/A 0.03fF
C67839 INVX1_LOC_251/Y INVX1_LOC_47/Y 0.01fF
C67840 NOR2X1_LOC_315/Y NOR2X1_LOC_89/a_36_216# 0.00fF
C67841 INVX1_LOC_47/A NOR2X1_LOC_814/A 0.17fF
C67842 INVX1_LOC_50/A INVX1_LOC_77/A 0.08fF
C67843 NOR2X1_LOC_433/A NOR2X1_LOC_654/A 0.03fF
C67844 INVX1_LOC_233/A NOR2X1_LOC_91/Y 0.15fF
C67845 NAND2X1_LOC_549/Y INVX1_LOC_61/A 0.09fF
C67846 NOR2X1_LOC_486/Y NAND2X1_LOC_472/Y 0.12fF
C67847 NOR2X1_LOC_576/B NOR2X1_LOC_36/B 0.11fF
C67848 NOR2X1_LOC_423/Y INVX1_LOC_78/A 0.04fF
C67849 NOR2X1_LOC_493/B NOR2X1_LOC_334/Y 0.02fF
C67850 NOR2X1_LOC_424/Y NOR2X1_LOC_89/A 0.06fF
C67851 INVX1_LOC_144/A NOR2X1_LOC_88/Y 0.04fF
C67852 NOR2X1_LOC_361/B INVX1_LOC_161/Y 0.17fF
C67853 NOR2X1_LOC_337/A NOR2X1_LOC_445/B 0.03fF
C67854 NOR2X1_LOC_186/Y INVX1_LOC_72/A 0.12fF
C67855 NOR2X1_LOC_142/Y INVX1_LOC_270/A 0.75fF
C67856 INVX1_LOC_143/A NAND2X1_LOC_223/A 0.01fF
C67857 NOR2X1_LOC_507/A INVX1_LOC_15/A 0.20fF
C67858 INVX1_LOC_64/A NOR2X1_LOC_363/a_36_216# 0.01fF
C67859 INVX1_LOC_22/A INVX1_LOC_231/A 0.03fF
C67860 NAND2X1_LOC_535/a_36_24# NAND2X1_LOC_537/Y 0.01fF
C67861 NAND2X1_LOC_579/A INVX1_LOC_31/A 2.18fF
C67862 INVX1_LOC_41/A D_INPUT_1 0.03fF
C67863 NOR2X1_LOC_222/Y INVX1_LOC_78/A 0.03fF
C67864 NAND2X1_LOC_660/Y INVX1_LOC_32/A 3.05fF
C67865 INVX1_LOC_35/A NOR2X1_LOC_546/a_36_216# 0.00fF
C67866 NOR2X1_LOC_803/A INVX1_LOC_301/A 0.01fF
C67867 INVX1_LOC_83/A NOR2X1_LOC_640/B 0.01fF
C67868 INVX1_LOC_201/Y D_INPUT_1 0.09fF
C67869 NOR2X1_LOC_620/Y NAND2X1_LOC_363/B 0.01fF
C67870 NOR2X1_LOC_52/B NOR2X1_LOC_654/A 0.20fF
C67871 NOR2X1_LOC_593/Y INVX1_LOC_58/Y 0.03fF
C67872 INVX1_LOC_25/A NOR2X1_LOC_664/Y 0.07fF
C67873 NAND2X1_LOC_783/Y INVX1_LOC_11/A 0.02fF
C67874 INVX1_LOC_213/Y INVX1_LOC_23/A 0.01fF
C67875 INVX1_LOC_303/A NOR2X1_LOC_772/B 0.02fF
C67876 NOR2X1_LOC_83/Y INVX1_LOC_84/A 0.01fF
C67877 NAND2X1_LOC_738/B INVX1_LOC_240/A 0.02fF
C67878 NOR2X1_LOC_45/B NAND2X1_LOC_798/B 0.12fF
C67879 INVX1_LOC_163/A INVX1_LOC_195/Y 0.03fF
C67880 NOR2X1_LOC_423/a_36_216# INVX1_LOC_63/Y 0.01fF
C67881 INVX1_LOC_136/A NOR2X1_LOC_468/Y 0.07fF
C67882 D_INPUT_0 INVX1_LOC_32/A 0.76fF
C67883 NAND2X1_LOC_724/A INVX1_LOC_72/A 0.07fF
C67884 NOR2X1_LOC_799/B NOR2X1_LOC_640/Y 0.04fF
C67885 INVX1_LOC_209/Y NOR2X1_LOC_304/Y 0.00fF
C67886 NOR2X1_LOC_665/A NAND2X1_LOC_454/Y 0.07fF
C67887 INVX1_LOC_311/Y NOR2X1_LOC_833/B 0.03fF
C67888 INVX1_LOC_136/A NAND2X1_LOC_190/Y 0.03fF
C67889 NOR2X1_LOC_389/A NOR2X1_LOC_276/Y 0.01fF
C67890 NAND2X1_LOC_35/Y NAND2X1_LOC_464/Y 0.03fF
C67891 INVX1_LOC_255/Y INVX1_LOC_175/A 0.02fF
C67892 NOR2X1_LOC_329/B INVX1_LOC_42/A 0.10fF
C67893 INVX1_LOC_286/A INVX1_LOC_63/A 0.07fF
C67894 INVX1_LOC_52/Y NOR2X1_LOC_759/Y -0.00fF
C67895 NOR2X1_LOC_168/B INVX1_LOC_53/A 0.18fF
C67896 INVX1_LOC_285/Y INVX1_LOC_19/A 0.01fF
C67897 NOR2X1_LOC_781/a_36_216# NOR2X1_LOC_158/Y 0.01fF
C67898 NOR2X1_LOC_296/a_36_216# NOR2X1_LOC_791/B 0.00fF
C67899 INVX1_LOC_36/A NAND2X1_LOC_350/A 0.07fF
C67900 NOR2X1_LOC_454/Y INVX1_LOC_105/A 0.02fF
C67901 NOR2X1_LOC_332/B NOR2X1_LOC_865/Y 0.03fF
C67902 NOR2X1_LOC_56/Y NOR2X1_LOC_841/A 0.10fF
C67903 VDD INVX1_LOC_108/A 0.12fF
C67904 NOR2X1_LOC_217/a_36_216# INVX1_LOC_130/Y 0.00fF
C67905 INVX1_LOC_89/A NOR2X1_LOC_334/Y 0.07fF
C67906 INVX1_LOC_249/A INVX1_LOC_1/A 0.12fF
C67907 INVX1_LOC_215/A NOR2X1_LOC_65/Y 0.01fF
C67908 NOR2X1_LOC_332/B NOR2X1_LOC_243/B 0.01fF
C67909 NAND2X1_LOC_44/a_36_24# INVX1_LOC_174/A 0.00fF
C67910 D_INPUT_0 NAND2X1_LOC_175/Y 0.10fF
C67911 NOR2X1_LOC_634/A NOR2X1_LOC_857/A 0.07fF
C67912 NOR2X1_LOC_272/Y INVX1_LOC_8/A 1.52fF
C67913 NOR2X1_LOC_140/A NOR2X1_LOC_554/a_36_216# 0.00fF
C67914 INVX1_LOC_64/A NAND2X1_LOC_661/B 0.01fF
C67915 NOR2X1_LOC_45/Y INVX1_LOC_72/A 0.03fF
C67916 INVX1_LOC_95/Y INVX1_LOC_285/A 0.00fF
C67917 INVX1_LOC_208/Y INVX1_LOC_23/A 0.04fF
C67918 NOR2X1_LOC_785/Y INVX1_LOC_26/Y 0.01fF
C67919 INVX1_LOC_91/A INVX1_LOC_186/Y 2.23fF
C67920 NAND2X1_LOC_303/Y NOR2X1_LOC_387/Y 0.03fF
C67921 INVX1_LOC_36/A NOR2X1_LOC_441/Y 0.06fF
C67922 INVX1_LOC_136/A NOR2X1_LOC_389/A 0.00fF
C67923 NOR2X1_LOC_569/Y NOR2X1_LOC_748/A 0.03fF
C67924 INVX1_LOC_35/A NOR2X1_LOC_773/Y 0.07fF
C67925 NOR2X1_LOC_589/A INVX1_LOC_57/A 0.03fF
C67926 INVX1_LOC_135/A INVX1_LOC_23/Y 0.08fF
C67927 INVX1_LOC_95/Y NOR2X1_LOC_814/A 0.12fF
C67928 INVX1_LOC_235/Y NOR2X1_LOC_516/Y 0.26fF
C67929 INVX1_LOC_25/A INVX1_LOC_137/A 0.04fF
C67930 NAND2X1_LOC_860/A INVX1_LOC_16/A 0.15fF
C67931 INVX1_LOC_263/A NOR2X1_LOC_678/A 0.00fF
C67932 NAND2X1_LOC_363/B NAND2X1_LOC_194/a_36_24# 0.01fF
C67933 VDD NOR2X1_LOC_841/A 1.12fF
C67934 NOR2X1_LOC_139/Y INVX1_LOC_272/A 0.07fF
C67935 INVX1_LOC_65/A INVX1_LOC_19/A 2.40fF
C67936 INVX1_LOC_166/A NAND2X1_LOC_378/a_36_24# 0.01fF
C67937 INVX1_LOC_11/A NOR2X1_LOC_537/A 0.03fF
C67938 NOR2X1_LOC_349/A INVX1_LOC_29/A 0.09fF
C67939 INVX1_LOC_64/A INVX1_LOC_316/Y 0.38fF
C67940 INVX1_LOC_144/A INVX1_LOC_15/A 0.04fF
C67941 NOR2X1_LOC_329/B INVX1_LOC_78/A 0.33fF
C67942 VDD NOR2X1_LOC_801/A 0.24fF
C67943 NAND2X1_LOC_569/B INVX1_LOC_25/Y 0.10fF
C67944 INVX1_LOC_11/A NOR2X1_LOC_716/B 0.07fF
C67945 NOR2X1_LOC_75/Y NOR2X1_LOC_433/A 0.01fF
C67946 NOR2X1_LOC_607/a_36_216# INVX1_LOC_292/A 0.00fF
C67947 NOR2X1_LOC_584/a_36_216# INVX1_LOC_72/A 0.00fF
C67948 NOR2X1_LOC_405/A INVX1_LOC_29/A 0.16fF
C67949 NAND2X1_LOC_26/a_36_24# INVX1_LOC_1/A 0.01fF
C67950 NOR2X1_LOC_92/Y NOR2X1_LOC_591/Y 0.03fF
C67951 NOR2X1_LOC_35/Y NOR2X1_LOC_721/B 0.03fF
C67952 NOR2X1_LOC_468/Y NOR2X1_LOC_278/A 0.04fF
C67953 NOR2X1_LOC_662/A INVX1_LOC_20/A 0.13fF
C67954 NAND2X1_LOC_303/Y NAND2X1_LOC_357/B 0.02fF
C67955 NAND2X1_LOC_181/Y NOR2X1_LOC_791/Y 0.31fF
C67956 NOR2X1_LOC_730/B INVX1_LOC_15/A 0.03fF
C67957 NOR2X1_LOC_703/B INVX1_LOC_18/A 0.03fF
C67958 NAND2X1_LOC_468/B INVX1_LOC_272/A 0.01fF
C67959 NAND2X1_LOC_656/Y INVX1_LOC_53/A 0.21fF
C67960 INVX1_LOC_38/A NOR2X1_LOC_197/B 0.14fF
C67961 NOR2X1_LOC_848/Y NAND2X1_LOC_116/A 0.05fF
C67962 INVX1_LOC_89/A NAND2X1_LOC_607/a_36_24# 0.00fF
C67963 NOR2X1_LOC_222/Y NOR2X1_LOC_215/A 0.01fF
C67964 NAND2X1_LOC_725/A NOR2X1_LOC_32/Y 0.78fF
C67965 NOR2X1_LOC_516/B NOR2X1_LOC_849/A 0.01fF
C67966 INVX1_LOC_136/A INVX1_LOC_62/Y 0.11fF
C67967 NOR2X1_LOC_435/A INVX1_LOC_54/A 0.03fF
C67968 INVX1_LOC_108/A NAND2X1_LOC_41/a_36_24# 0.00fF
C67969 NOR2X1_LOC_65/B NOR2X1_LOC_329/B 0.01fF
C67970 INVX1_LOC_35/A NOR2X1_LOC_332/A 0.09fF
C67971 NAND2X1_LOC_656/A NOR2X1_LOC_554/B 0.19fF
C67972 INVX1_LOC_303/A NOR2X1_LOC_500/B 0.10fF
C67973 NOR2X1_LOC_703/Y NOR2X1_LOC_334/Y 2.01fF
C67974 NOR2X1_LOC_75/Y NOR2X1_LOC_52/B 0.00fF
C67975 NOR2X1_LOC_857/A INVX1_LOC_29/A 0.08fF
C67976 NOR2X1_LOC_620/Y INVX1_LOC_30/A 0.00fF
C67977 INVX1_LOC_17/A INVX1_LOC_276/A 0.22fF
C67978 NOR2X1_LOC_168/Y INVX1_LOC_94/A 0.12fF
C67979 INVX1_LOC_230/Y NOR2X1_LOC_6/B 0.11fF
C67980 INVX1_LOC_186/Y NOR2X1_LOC_698/Y 0.21fF
C67981 NAND2X1_LOC_848/A NAND2X1_LOC_489/Y 0.07fF
C67982 INVX1_LOC_125/Y INVX1_LOC_4/Y 0.10fF
C67983 D_INPUT_3 NOR2X1_LOC_610/a_36_216# 0.00fF
C67984 VDD INPUT_7 0.18fF
C67985 INVX1_LOC_161/Y INVX1_LOC_177/A 0.16fF
C67986 INVX1_LOC_25/A NOR2X1_LOC_19/B 0.71fF
C67987 NOR2X1_LOC_590/A NOR2X1_LOC_574/A 0.06fF
C67988 NAND2X1_LOC_860/A INVX1_LOC_28/A 0.02fF
C67989 NOR2X1_LOC_690/A NOR2X1_LOC_372/a_36_216# 0.00fF
C67990 NOR2X1_LOC_441/Y NOR2X1_LOC_309/Y 0.07fF
C67991 NOR2X1_LOC_598/B INVX1_LOC_311/Y 0.03fF
C67992 NAND2X1_LOC_213/A NAND2X1_LOC_158/a_36_24# 0.01fF
C67993 NOR2X1_LOC_553/a_36_216# INVX1_LOC_177/A 0.00fF
C67994 NOR2X1_LOC_602/B INVX1_LOC_63/A 0.10fF
C67995 INVX1_LOC_36/A NOR2X1_LOC_142/Y 0.04fF
C67996 INVX1_LOC_14/A INVX1_LOC_56/Y 0.03fF
C67997 NOR2X1_LOC_75/Y NOR2X1_LOC_603/a_36_216# 0.00fF
C67998 NAND2X1_LOC_537/Y INVX1_LOC_16/A 0.07fF
C67999 NAND2X1_LOC_611/a_36_24# INVX1_LOC_42/A 0.01fF
C68000 NAND2X1_LOC_725/A NOR2X1_LOC_597/A 0.04fF
C68001 INVX1_LOC_211/Y NOR2X1_LOC_226/A 0.02fF
C68002 INVX1_LOC_41/A NOR2X1_LOC_778/A 0.00fF
C68003 NAND2X1_LOC_579/A NAND2X1_LOC_859/Y 0.09fF
C68004 INVX1_LOC_54/A INVX1_LOC_63/A 0.10fF
C68005 NAND2X1_LOC_733/Y NOR2X1_LOC_504/Y 0.70fF
C68006 INPUT_1 NOR2X1_LOC_293/a_36_216# 0.00fF
C68007 NOR2X1_LOC_590/A INVX1_LOC_196/A 0.01fF
C68008 INVX1_LOC_225/A INVX1_LOC_72/A 0.10fF
C68009 NOR2X1_LOC_272/Y NAND2X1_LOC_140/A 0.03fF
C68010 INVX1_LOC_90/A INVX1_LOC_38/Y 0.13fF
C68011 NAND2X1_LOC_364/A INVX1_LOC_8/A 0.00fF
C68012 NOR2X1_LOC_322/a_36_216# NOR2X1_LOC_89/A 0.00fF
C68013 INPUT_2 NAND2X1_LOC_672/B 0.00fF
C68014 INVX1_LOC_24/A INVX1_LOC_33/A 0.15fF
C68015 INVX1_LOC_238/Y NAND2X1_LOC_733/B 0.04fF
C68016 NOR2X1_LOC_266/B INVX1_LOC_32/A 0.03fF
C68017 NOR2X1_LOC_155/A INVX1_LOC_84/A 0.03fF
C68018 INVX1_LOC_255/Y NOR2X1_LOC_82/A 0.09fF
C68019 NOR2X1_LOC_723/Y INVX1_LOC_266/Y 0.01fF
C68020 NOR2X1_LOC_530/Y INVX1_LOC_25/Y 0.03fF
C68021 INVX1_LOC_298/Y NOR2X1_LOC_405/A 0.02fF
C68022 NOR2X1_LOC_759/Y INVX1_LOC_63/Y 0.10fF
C68023 NAND2X1_LOC_338/B INVX1_LOC_170/A 0.00fF
C68024 NOR2X1_LOC_208/Y NOR2X1_LOC_142/Y 0.16fF
C68025 INVX1_LOC_21/A NOR2X1_LOC_356/A 0.08fF
C68026 NOR2X1_LOC_655/B INVX1_LOC_36/A 0.00fF
C68027 NOR2X1_LOC_78/B INVX1_LOC_312/Y 0.19fF
C68028 INVX1_LOC_201/Y D_INPUT_2 0.06fF
C68029 NOR2X1_LOC_537/A NOR2X1_LOC_593/Y 0.04fF
C68030 INVX1_LOC_65/A INVX1_LOC_26/Y 0.00fF
C68031 NOR2X1_LOC_852/B NAND2X1_LOC_361/Y 0.02fF
C68032 NOR2X1_LOC_209/Y INVX1_LOC_142/Y 0.03fF
C68033 NOR2X1_LOC_501/B INVX1_LOC_23/A 0.01fF
C68034 NAND2X1_LOC_594/a_36_24# NAND2X1_LOC_807/Y 0.00fF
C68035 VDD INVX1_LOC_128/A 0.12fF
C68036 INVX1_LOC_224/Y NOR2X1_LOC_78/A 0.04fF
C68037 INVX1_LOC_2/A NOR2X1_LOC_759/A 0.16fF
C68038 NOR2X1_LOC_516/B NOR2X1_LOC_514/A 0.04fF
C68039 INVX1_LOC_11/A NOR2X1_LOC_717/B 0.03fF
C68040 NAND2X1_LOC_348/A INVX1_LOC_38/Y 0.01fF
C68041 NOR2X1_LOC_158/Y NOR2X1_LOC_586/Y 0.21fF
C68042 INVX1_LOC_206/Y NOR2X1_LOC_678/A 0.03fF
C68043 NOR2X1_LOC_557/Y INVX1_LOC_33/A 0.11fF
C68044 INVX1_LOC_299/A NOR2X1_LOC_788/B 0.00fF
C68045 INVX1_LOC_136/A NOR2X1_LOC_220/A 0.02fF
C68046 NOR2X1_LOC_209/Y INVX1_LOC_198/Y 0.10fF
C68047 NOR2X1_LOC_82/A NOR2X1_LOC_71/Y 0.16fF
C68048 NOR2X1_LOC_403/B NOR2X1_LOC_398/Y 0.10fF
C68049 NAND2X1_LOC_812/A GATE_811 0.14fF
C68050 NAND2X1_LOC_579/A NAND2X1_LOC_807/Y 0.04fF
C68051 INVX1_LOC_1/A NOR2X1_LOC_772/A 0.01fF
C68052 INVX1_LOC_26/A NAND2X1_LOC_266/a_36_24# 0.00fF
C68053 INVX1_LOC_1/A NOR2X1_LOC_19/B 0.09fF
C68054 INVX1_LOC_21/A NOR2X1_LOC_74/A 0.63fF
C68055 NAND2X1_LOC_537/Y INVX1_LOC_28/A 0.48fF
C68056 NAND2X1_LOC_390/A INVX1_LOC_30/A 0.50fF
C68057 NOR2X1_LOC_716/B NOR2X1_LOC_52/B 0.80fF
C68058 NOR2X1_LOC_423/Y INVX1_LOC_113/Y 0.06fF
C68059 INPUT_3 D_INPUT_0 0.08fF
C68060 NOR2X1_LOC_383/B INVX1_LOC_143/Y 0.03fF
C68061 INVX1_LOC_24/A NAND2X1_LOC_798/A 0.03fF
C68062 NAND2X1_LOC_360/B INVX1_LOC_314/Y 0.01fF
C68063 INVX1_LOC_27/A NOR2X1_LOC_188/A 0.07fF
C68064 INVX1_LOC_75/A NAND2X1_LOC_218/A 0.02fF
C68065 INVX1_LOC_24/A INVX1_LOC_40/A 0.03fF
C68066 NAND2X1_LOC_222/A D_INPUT_3 0.02fF
C68067 NOR2X1_LOC_140/A INVX1_LOC_75/A 0.02fF
C68068 NOR2X1_LOC_600/Y NOR2X1_LOC_678/A 0.00fF
C68069 NOR2X1_LOC_433/A INVX1_LOC_98/Y 0.33fF
C68070 INVX1_LOC_57/A INVX1_LOC_20/A 0.55fF
C68071 INVX1_LOC_132/A NOR2X1_LOC_537/Y 0.07fF
C68072 NOR2X1_LOC_742/a_36_216# INVX1_LOC_311/Y 0.00fF
C68073 INVX1_LOC_83/A INVX1_LOC_141/Y 0.23fF
C68074 INVX1_LOC_21/A NOR2X1_LOC_9/Y 0.03fF
C68075 INVX1_LOC_24/A INVX1_LOC_165/Y 0.01fF
C68076 NOR2X1_LOC_836/Y NAND2X1_LOC_363/Y 0.03fF
C68077 INVX1_LOC_12/A NOR2X1_LOC_697/Y 0.08fF
C68078 NAND2X1_LOC_228/a_36_24# INVX1_LOC_159/A 0.00fF
C68079 NOR2X1_LOC_369/Y INVX1_LOC_90/A 0.40fF
C68080 INVX1_LOC_244/Y INVX1_LOC_22/A 0.00fF
C68081 NAND2X1_LOC_848/A NAND2X1_LOC_175/Y 0.10fF
C68082 NOR2X1_LOC_813/Y INVX1_LOC_23/Y 0.02fF
C68083 NOR2X1_LOC_84/A NOR2X1_LOC_84/Y 0.05fF
C68084 INVX1_LOC_33/A INVX1_LOC_143/A 0.06fF
C68085 NOR2X1_LOC_222/Y INVX1_LOC_113/Y 0.17fF
C68086 INVX1_LOC_234/A NOR2X1_LOC_384/Y 0.00fF
C68087 NOR2X1_LOC_41/Y INVX1_LOC_63/Y 0.01fF
C68088 INVX1_LOC_83/A INVX1_LOC_312/Y 0.02fF
C68089 NOR2X1_LOC_294/Y INVX1_LOC_83/A 0.25fF
C68090 INVX1_LOC_36/A NOR2X1_LOC_99/B 0.01fF
C68091 NOR2X1_LOC_15/Y NOR2X1_LOC_313/Y 0.02fF
C68092 NAND2X1_LOC_223/A NOR2X1_LOC_16/a_36_216# 0.00fF
C68093 INVX1_LOC_32/A INVX1_LOC_46/Y 0.09fF
C68094 INVX1_LOC_90/A INVX1_LOC_286/Y 0.04fF
C68095 INVX1_LOC_11/A NOR2X1_LOC_151/Y 0.03fF
C68096 INVX1_LOC_41/A NOR2X1_LOC_620/B 0.00fF
C68097 NOR2X1_LOC_89/A NOR2X1_LOC_666/a_36_216# 0.02fF
C68098 NOR2X1_LOC_155/A INVX1_LOC_15/A 0.11fF
C68099 NAND2X1_LOC_487/a_36_24# INVX1_LOC_4/A 0.01fF
C68100 NOR2X1_LOC_159/a_36_216# NAND2X1_LOC_572/B 0.00fF
C68101 NAND2X1_LOC_579/A INVX1_LOC_6/A 0.03fF
C68102 NAND2X1_LOC_472/Y NOR2X1_LOC_748/A 0.10fF
C68103 NAND2X1_LOC_807/B INVX1_LOC_63/A 0.04fF
C68104 INVX1_LOC_277/A NOR2X1_LOC_724/Y 0.07fF
C68105 INVX1_LOC_36/A NOR2X1_LOC_846/B 0.02fF
C68106 INVX1_LOC_224/Y NOR2X1_LOC_98/a_36_216# 0.03fF
C68107 NOR2X1_LOC_655/B NOR2X1_LOC_309/Y 0.03fF
C68108 INVX1_LOC_304/A INVX1_LOC_306/Y 0.44fF
C68109 NOR2X1_LOC_830/Y INVX1_LOC_19/A 0.07fF
C68110 INVX1_LOC_13/A INVX1_LOC_49/A 0.02fF
C68111 NOR2X1_LOC_288/A NAND2X1_LOC_323/B 0.05fF
C68112 INVX1_LOC_5/A NOR2X1_LOC_347/a_36_216# 0.02fF
C68113 INVX1_LOC_83/A NOR2X1_LOC_546/B 0.03fF
C68114 NOR2X1_LOC_168/B NOR2X1_LOC_634/B 0.03fF
C68115 NOR2X1_LOC_220/a_36_216# INVX1_LOC_171/A 0.00fF
C68116 NOR2X1_LOC_663/A D_GATE_662 0.01fF
C68117 INVX1_LOC_90/A INVX1_LOC_159/A 0.02fF
C68118 INVX1_LOC_50/A INVX1_LOC_9/A 0.16fF
C68119 INVX1_LOC_186/Y NOR2X1_LOC_483/a_36_216# 0.00fF
C68120 NAND2X1_LOC_363/B INVX1_LOC_117/A 0.02fF
C68121 NOR2X1_LOC_384/Y NOR2X1_LOC_19/B 0.00fF
C68122 NOR2X1_LOC_105/Y INVX1_LOC_9/A 0.01fF
C68123 INVX1_LOC_90/A NOR2X1_LOC_191/B 0.01fF
C68124 NOR2X1_LOC_103/Y INVX1_LOC_98/A 0.00fF
C68125 INVX1_LOC_25/Y NOR2X1_LOC_709/A 0.02fF
C68126 INVX1_LOC_13/A INVX1_LOC_60/A 0.01fF
C68127 INVX1_LOC_83/A INVX1_LOC_275/A 0.05fF
C68128 NOR2X1_LOC_717/B NOR2X1_LOC_593/Y 0.03fF
C68129 NOR2X1_LOC_389/B NOR2X1_LOC_191/B 0.08fF
C68130 NOR2X1_LOC_103/Y NOR2X1_LOC_78/A 0.07fF
C68131 NOR2X1_LOC_35/Y NAND2X1_LOC_473/A 0.10fF
C68132 NOR2X1_LOC_755/Y NAND2X1_LOC_792/B 0.00fF
C68133 NAND2X1_LOC_256/a_36_24# NOR2X1_LOC_197/B 0.00fF
C68134 NAND2X1_LOC_739/B NOR2X1_LOC_385/Y 0.04fF
C68135 INVX1_LOC_251/A NAND2X1_LOC_74/B 0.01fF
C68136 INVX1_LOC_2/A INVX1_LOC_13/A 0.01fF
C68137 NAND2X1_LOC_374/Y INVX1_LOC_22/A 0.03fF
C68138 INVX1_LOC_55/Y INVX1_LOC_49/A 0.06fF
C68139 NAND2X1_LOC_72/Y INVX1_LOC_9/A 0.08fF
C68140 INVX1_LOC_19/A INVX1_LOC_4/Y 0.37fF
C68141 NOR2X1_LOC_329/B NOR2X1_LOC_152/Y 0.67fF
C68142 INVX1_LOC_135/A NAND2X1_LOC_116/A 0.02fF
C68143 NOR2X1_LOC_360/Y INPUT_0 0.03fF
C68144 NOR2X1_LOC_75/Y INVX1_LOC_199/A 0.06fF
C68145 NOR2X1_LOC_415/a_36_216# NOR2X1_LOC_6/B 0.01fF
C68146 NOR2X1_LOC_503/A NOR2X1_LOC_433/A 0.01fF
C68147 INVX1_LOC_24/A NOR2X1_LOC_323/Y 0.01fF
C68148 D_INPUT_0 INVX1_LOC_158/A 0.01fF
C68149 NAND2X1_LOC_456/Y INVX1_LOC_26/A 0.02fF
C68150 INVX1_LOC_25/A NOR2X1_LOC_216/B 0.30fF
C68151 INVX1_LOC_89/A NOR2X1_LOC_718/B 0.19fF
C68152 NOR2X1_LOC_833/B INVX1_LOC_15/A 0.03fF
C68153 INVX1_LOC_161/Y NOR2X1_LOC_137/B 0.04fF
C68154 INVX1_LOC_135/Y NOR2X1_LOC_474/A 0.15fF
C68155 INVX1_LOC_45/A INVX1_LOC_98/A 0.14fF
C68156 NOR2X1_LOC_717/A INVX1_LOC_92/A 0.15fF
C68157 INVX1_LOC_18/A INVX1_LOC_309/A 0.01fF
C68158 INVX1_LOC_230/Y NOR2X1_LOC_124/A 0.03fF
C68159 NAND2X1_LOC_609/a_36_24# NAND2X1_LOC_215/A 0.01fF
C68160 NOR2X1_LOC_168/B INVX1_LOC_83/A 0.03fF
C68161 NAND2X1_LOC_572/a_36_24# NOR2X1_LOC_123/B 0.00fF
C68162 NOR2X1_LOC_392/Y NOR2X1_LOC_104/a_36_216# 0.00fF
C68163 INVX1_LOC_45/A NOR2X1_LOC_78/A 0.19fF
C68164 NOR2X1_LOC_532/a_36_216# INVX1_LOC_91/A 0.01fF
C68165 INVX1_LOC_18/A NOR2X1_LOC_114/A 0.02fF
C68166 NOR2X1_LOC_78/B NAND2X1_LOC_656/Y 0.29fF
C68167 INVX1_LOC_30/A NAND2X1_LOC_623/B 2.21fF
C68168 D_INPUT_1 NAND2X1_LOC_574/A 0.04fF
C68169 INVX1_LOC_312/Y NOR2X1_LOC_311/Y 0.00fF
C68170 INVX1_LOC_2/A NOR2X1_LOC_246/A 0.09fF
C68171 INVX1_LOC_2/A NOR2X1_LOC_503/a_36_216# 0.02fF
C68172 NOR2X1_LOC_216/Y INVX1_LOC_33/A 0.26fF
C68173 NOR2X1_LOC_151/Y NOR2X1_LOC_593/Y 0.03fF
C68174 NOR2X1_LOC_366/B NOR2X1_LOC_366/Y 0.01fF
C68175 NAND2X1_LOC_53/Y INVX1_LOC_37/A 0.07fF
C68176 NOR2X1_LOC_394/Y NAND2X1_LOC_254/Y 0.08fF
C68177 INVX1_LOC_18/A INVX1_LOC_91/A 0.45fF
C68178 NOR2X1_LOC_690/A NAND2X1_LOC_849/A 0.02fF
C68179 NOR2X1_LOC_68/a_36_216# INVX1_LOC_57/A 0.00fF
C68180 NOR2X1_LOC_112/B INVX1_LOC_33/A 0.01fF
C68181 INVX1_LOC_13/Y NOR2X1_LOC_99/Y 0.07fF
C68182 NAND2X1_LOC_7/Y INVX1_LOC_92/Y 0.04fF
C68183 INVX1_LOC_72/A NAND2X1_LOC_642/Y 0.55fF
C68184 INVX1_LOC_2/A INVX1_LOC_55/Y 0.06fF
C68185 INVX1_LOC_269/A NOR2X1_LOC_536/A 0.04fF
C68186 INVX1_LOC_284/Y NAND2X1_LOC_836/Y -0.04fF
C68187 INVX1_LOC_172/A INVX1_LOC_309/A 0.03fF
C68188 NOR2X1_LOC_598/B INVX1_LOC_84/A 0.07fF
C68189 NOR2X1_LOC_470/B INVX1_LOC_38/A 0.01fF
C68190 NOR2X1_LOC_590/A NOR2X1_LOC_305/Y 0.00fF
C68191 INVX1_LOC_89/A INVX1_LOC_218/A 0.04fF
C68192 NOR2X1_LOC_232/Y NOR2X1_LOC_536/A 0.05fF
C68193 INVX1_LOC_78/A NOR2X1_LOC_477/B 0.01fF
C68194 INVX1_LOC_36/A NAND2X1_LOC_274/a_36_24# 0.00fF
C68195 INVX1_LOC_135/A INVX1_LOC_232/A 0.16fF
C68196 NOR2X1_LOC_720/A NAND2X1_LOC_207/B 0.02fF
C68197 NAND2X1_LOC_564/B D_INPUT_0 0.07fF
C68198 NOR2X1_LOC_561/Y NAND2X1_LOC_319/A 0.02fF
C68199 NOR2X1_LOC_713/B INVX1_LOC_91/A 0.08fF
C68200 INVX1_LOC_208/Y INVX1_LOC_313/A 0.03fF
C68201 NOR2X1_LOC_78/A INVX1_LOC_71/A 0.08fF
C68202 INVX1_LOC_266/A NOR2X1_LOC_641/Y 0.08fF
C68203 NAND2X1_LOC_349/B NOR2X1_LOC_106/A 0.17fF
C68204 NAND2X1_LOC_181/a_36_24# NOR2X1_LOC_71/Y 0.01fF
C68205 INVX1_LOC_75/A NOR2X1_LOC_709/A 0.03fF
C68206 NAND2X1_LOC_850/A NAND2X1_LOC_850/Y 0.18fF
C68207 NOR2X1_LOC_389/B NOR2X1_LOC_568/a_36_216# 0.00fF
C68208 NAND2X1_LOC_785/B VDD 0.02fF
C68209 NOR2X1_LOC_510/Y NOR2X1_LOC_841/A 0.10fF
C68210 INVX1_LOC_172/A INVX1_LOC_91/A 0.12fF
C68211 INVX1_LOC_312/Y INVX1_LOC_46/A 0.07fF
C68212 INVX1_LOC_24/A NOR2X1_LOC_486/Y 5.13fF
C68213 INVX1_LOC_89/A NOR2X1_LOC_569/Y 0.68fF
C68214 NAND2X1_LOC_711/B INVX1_LOC_11/Y 0.19fF
C68215 INVX1_LOC_64/A NOR2X1_LOC_662/A 0.03fF
C68216 INVX1_LOC_269/A NOR2X1_LOC_655/Y 0.00fF
C68217 INVX1_LOC_21/A NOR2X1_LOC_865/Y 0.02fF
C68218 NOR2X1_LOC_828/B NOR2X1_LOC_731/Y 0.04fF
C68219 INVX1_LOC_21/A NOR2X1_LOC_243/B 0.09fF
C68220 INVX1_LOC_245/Y NOR2X1_LOC_261/A 0.01fF
C68221 INVX1_LOC_206/A NOR2X1_LOC_188/A 0.78fF
C68222 INVX1_LOC_13/A INPUT_1 0.06fF
C68223 INVX1_LOC_269/A NAND2X1_LOC_93/B 0.17fF
C68224 INVX1_LOC_30/A INVX1_LOC_117/A 0.27fF
C68225 INVX1_LOC_1/A NOR2X1_LOC_216/B 0.10fF
C68226 INVX1_LOC_211/Y INVX1_LOC_118/A 0.22fF
C68227 INVX1_LOC_34/A NOR2X1_LOC_269/Y 0.01fF
C68228 NOR2X1_LOC_667/A NOR2X1_LOC_74/A 0.01fF
C68229 INVX1_LOC_103/A INVX1_LOC_179/A 0.03fF
C68230 INVX1_LOC_286/Y INVX1_LOC_38/A 0.07fF
C68231 NAND2X1_LOC_763/B INVX1_LOC_117/A 0.01fF
C68232 INVX1_LOC_14/A NOR2X1_LOC_831/B 0.01fF
C68233 NAND2X1_LOC_200/B NOR2X1_LOC_188/A 0.03fF
C68234 INVX1_LOC_35/A NOR2X1_LOC_847/A 0.05fF
C68235 NOR2X1_LOC_367/B INVX1_LOC_159/Y 0.24fF
C68236 NOR2X1_LOC_598/B NAND2X1_LOC_220/B 0.08fF
C68237 NOR2X1_LOC_172/Y NOR2X1_LOC_56/Y 0.03fF
C68238 INVX1_LOC_26/Y INVX1_LOC_4/Y 0.07fF
C68239 NAND2X1_LOC_200/B NOR2X1_LOC_548/B 0.12fF
C68240 NAND2X1_LOC_350/A NOR2X1_LOC_435/A 0.20fF
C68241 NOR2X1_LOC_503/a_36_216# NAND2X1_LOC_648/A 0.00fF
C68242 INVX1_LOC_35/A INVX1_LOC_42/A 0.11fF
C68243 INVX1_LOC_43/A INVX1_LOC_6/A 0.01fF
C68244 NOR2X1_LOC_388/Y NAND2X1_LOC_447/Y 0.10fF
C68245 INVX1_LOC_49/A NOR2X1_LOC_357/Y 0.05fF
C68246 INVX1_LOC_57/A INVX1_LOC_4/A 1.79fF
C68247 INVX1_LOC_72/A NOR2X1_LOC_271/Y 0.01fF
C68248 INVX1_LOC_269/A NOR2X1_LOC_649/B 1.42fF
C68249 NAND2X1_LOC_773/Y NOR2X1_LOC_814/A 1.60fF
C68250 INVX1_LOC_34/Y INVX1_LOC_91/A 0.21fF
C68251 INVX1_LOC_269/A INVX1_LOC_3/A 0.07fF
C68252 INPUT_3 INVX1_LOC_46/Y 0.07fF
C68253 INVX1_LOC_286/Y NOR2X1_LOC_51/A 0.03fF
C68254 NOR2X1_LOC_414/Y NOR2X1_LOC_38/B 0.01fF
C68255 NOR2X1_LOC_391/B INVX1_LOC_232/A 0.02fF
C68256 INVX1_LOC_24/A NOR2X1_LOC_816/Y 0.02fF
C68257 NOR2X1_LOC_598/B INVX1_LOC_15/A 0.43fF
C68258 NOR2X1_LOC_790/A INVX1_LOC_19/A 0.01fF
C68259 INVX1_LOC_159/A INVX1_LOC_38/A 0.15fF
C68260 NOR2X1_LOC_172/Y VDD 0.57fF
C68261 NOR2X1_LOC_772/Y VDD 0.09fF
C68262 NOR2X1_LOC_372/A NOR2X1_LOC_88/Y 0.03fF
C68263 NAND2X1_LOC_483/Y INVX1_LOC_46/A 0.01fF
C68264 INVX1_LOC_286/A INVX1_LOC_1/Y 0.16fF
C68265 NOR2X1_LOC_537/Y NAND2X1_LOC_642/Y 0.03fF
C68266 NOR2X1_LOC_565/B NOR2X1_LOC_74/A 0.00fF
C68267 NOR2X1_LOC_658/Y INVX1_LOC_92/A 0.42fF
C68268 NOR2X1_LOC_147/B VDD 0.78fF
C68269 NOR2X1_LOC_722/a_36_216# INVX1_LOC_139/Y 0.00fF
C68270 NAND2X1_LOC_338/B NAND2X1_LOC_642/Y 0.03fF
C68271 INVX1_LOC_271/A NOR2X1_LOC_338/a_36_216# 0.00fF
C68272 INVX1_LOC_49/A NOR2X1_LOC_319/B 0.03fF
C68273 NOR2X1_LOC_392/B VDD 2.09fF
C68274 INVX1_LOC_1/A NAND2X1_LOC_82/a_36_24# 0.00fF
C68275 NOR2X1_LOC_328/Y NOR2X1_LOC_45/B 0.12fF
C68276 NOR2X1_LOC_52/B NAND2X1_LOC_633/Y 0.14fF
C68277 NAND2X1_LOC_350/A INVX1_LOC_63/A 0.08fF
C68278 INVX1_LOC_88/A INVX1_LOC_272/A 0.76fF
C68279 NOR2X1_LOC_791/Y INVX1_LOC_3/Y 0.03fF
C68280 INVX1_LOC_35/A INVX1_LOC_78/A 0.10fF
C68281 INVX1_LOC_2/A NOR2X1_LOC_357/Y 1.17fF
C68282 NAND2X1_LOC_114/B NOR2X1_LOC_68/Y 0.04fF
C68283 NOR2X1_LOC_134/Y NAND2X1_LOC_489/Y 0.26fF
C68284 INVX1_LOC_90/A NOR2X1_LOC_721/Y 0.02fF
C68285 INVX1_LOC_218/Y INVX1_LOC_63/A 0.03fF
C68286 NAND2X1_LOC_137/a_36_24# NOR2X1_LOC_536/A 0.00fF
C68287 NOR2X1_LOC_441/Y INVX1_LOC_63/A 0.09fF
C68288 INVX1_LOC_24/A INVX1_LOC_241/Y 0.08fF
C68289 INVX1_LOC_296/A NOR2X1_LOC_452/A 0.03fF
C68290 INVX1_LOC_17/A NOR2X1_LOC_584/Y 0.03fF
C68291 NOR2X1_LOC_510/Y INVX1_LOC_128/A 0.01fF
C68292 NAND2X1_LOC_20/B NAND2X1_LOC_20/a_36_24# 0.00fF
C68293 NOR2X1_LOC_210/B INVX1_LOC_115/A 0.01fF
C68294 INVX1_LOC_141/A INVX1_LOC_49/Y 0.01fF
C68295 NOR2X1_LOC_123/B INVX1_LOC_98/A 0.14fF
C68296 NOR2X1_LOC_690/Y INVX1_LOC_11/Y 0.03fF
C68297 INVX1_LOC_255/Y INVX1_LOC_59/Y 0.13fF
C68298 NAND2X1_LOC_116/A INVX1_LOC_280/A 0.23fF
C68299 INVX1_LOC_35/A NOR2X1_LOC_65/B 0.10fF
C68300 NOR2X1_LOC_470/A INVX1_LOC_199/A 0.07fF
C68301 NOR2X1_LOC_123/B NOR2X1_LOC_78/A 0.07fF
C68302 INPUT_0 NOR2X1_LOC_567/B 0.07fF
C68303 NOR2X1_LOC_218/Y NOR2X1_LOC_357/Y 0.10fF
C68304 NOR2X1_LOC_91/Y INVX1_LOC_119/Y 0.03fF
C68305 NOR2X1_LOC_500/Y INVX1_LOC_37/A 0.46fF
C68306 INVX1_LOC_58/A NAND2X1_LOC_787/A 0.03fF
C68307 NOR2X1_LOC_749/Y NOR2X1_LOC_78/A 0.09fF
C68308 NOR2X1_LOC_32/B INVX1_LOC_23/A 0.70fF
C68309 D_INPUT_2 NAND2X1_LOC_574/A 0.06fF
C68310 NOR2X1_LOC_666/Y INVX1_LOC_4/A -0.01fF
C68311 NOR2X1_LOC_6/B NOR2X1_LOC_641/Y 0.85fF
C68312 INVX1_LOC_314/Y NAND2X1_LOC_572/B 0.28fF
C68313 INVX1_LOC_64/A INVX1_LOC_57/A 0.16fF
C68314 NOR2X1_LOC_261/Y NOR2X1_LOC_598/B 0.54fF
C68315 NAND2X1_LOC_338/B NOR2X1_LOC_271/Y 0.06fF
C68316 INVX1_LOC_33/A NOR2X1_LOC_197/B 0.01fF
C68317 INVX1_LOC_72/A NOR2X1_LOC_48/Y 0.01fF
C68318 INVX1_LOC_108/Y NOR2X1_LOC_598/B 0.08fF
C68319 INVX1_LOC_53/A NOR2X1_LOC_717/A 0.16fF
C68320 INVX1_LOC_63/Y NOR2X1_LOC_13/a_36_216# 0.00fF
C68321 NAND2X1_LOC_142/a_36_24# INVX1_LOC_92/A 0.01fF
C68322 INVX1_LOC_311/A NOR2X1_LOC_74/A 0.07fF
C68323 INVX1_LOC_232/A NOR2X1_LOC_813/Y 0.04fF
C68324 NAND2X1_LOC_35/Y D_INPUT_1 0.03fF
C68325 NAND2X1_LOC_740/Y NOR2X1_LOC_829/Y 0.01fF
C68326 INVX1_LOC_58/A NAND2X1_LOC_565/a_36_24# 0.00fF
C68327 NOR2X1_LOC_776/a_36_216# INVX1_LOC_15/A 0.01fF
C68328 INVX1_LOC_98/A INVX1_LOC_102/Y 0.00fF
C68329 NOR2X1_LOC_52/B INVX1_LOC_71/Y 0.01fF
C68330 INVX1_LOC_35/A INVX1_LOC_152/Y 0.02fF
C68331 INVX1_LOC_90/A NOR2X1_LOC_56/Y 0.07fF
C68332 INVX1_LOC_10/A INVX1_LOC_37/A 0.02fF
C68333 NAND2X1_LOC_656/Y INVX1_LOC_46/A 0.09fF
C68334 INVX1_LOC_39/A NOR2X1_LOC_646/B 0.01fF
C68335 NOR2X1_LOC_130/Y INVX1_LOC_74/A 0.04fF
C68336 NAND2X1_LOC_595/a_36_24# NAND2X1_LOC_223/A 0.01fF
C68337 NOR2X1_LOC_456/Y INVX1_LOC_5/A 0.04fF
C68338 NOR2X1_LOC_92/Y NOR2X1_LOC_318/A 0.01fF
C68339 NAND2X1_LOC_564/B NAND2X1_LOC_848/A 0.10fF
C68340 INVX1_LOC_232/A INVX1_LOC_280/A 0.16fF
C68341 INVX1_LOC_97/A VDD 0.00fF
C68342 NAND2X1_LOC_112/Y NOR2X1_LOC_331/B 0.01fF
C68343 NAND2X1_LOC_470/a_36_24# NAND2X1_LOC_798/B 0.00fF
C68344 INPUT_0 NOR2X1_LOC_269/Y 0.12fF
C68345 INVX1_LOC_90/A VDD 2.46fF
C68346 INVX1_LOC_111/Y NOR2X1_LOC_831/B 0.00fF
C68347 NOR2X1_LOC_256/Y NOR2X1_LOC_124/A 0.01fF
C68348 NOR2X1_LOC_548/A INVX1_LOC_91/A 0.02fF
C68349 NOR2X1_LOC_151/Y NOR2X1_LOC_601/Y 0.15fF
C68350 INVX1_LOC_1/Y INVX1_LOC_54/A 1.29fF
C68351 INVX1_LOC_50/A NAND2X1_LOC_67/Y 0.01fF
C68352 NOR2X1_LOC_389/B VDD 0.57fF
C68353 NOR2X1_LOC_590/A INVX1_LOC_271/Y 0.07fF
C68354 INVX1_LOC_89/A NAND2X1_LOC_472/Y 0.09fF
C68355 NAND2X1_LOC_7/Y INVX1_LOC_106/A 0.02fF
C68356 INVX1_LOC_136/A INVX1_LOC_251/A 0.03fF
C68357 NAND2X1_LOC_127/a_36_24# INVX1_LOC_3/A 0.01fF
C68358 INVX1_LOC_177/A NOR2X1_LOC_801/A 0.01fF
C68359 NOR2X1_LOC_354/Y INVX1_LOC_160/A 0.11fF
C68360 INVX1_LOC_208/Y INVX1_LOC_131/Y 0.04fF
C68361 INVX1_LOC_123/A NOR2X1_LOC_845/A 0.03fF
C68362 INVX1_LOC_34/A NOR2X1_LOC_36/B 0.00fF
C68363 INVX1_LOC_88/A NOR2X1_LOC_125/a_36_216# 0.00fF
C68364 INVX1_LOC_256/A NOR2X1_LOC_621/A 0.01fF
C68365 NOR2X1_LOC_852/A NOR2X1_LOC_839/B 0.02fF
C68366 NOR2X1_LOC_99/B NOR2X1_LOC_865/A 0.05fF
C68367 INVX1_LOC_214/Y NOR2X1_LOC_697/Y 0.02fF
C68368 NAND2X1_LOC_176/a_36_24# NAND2X1_LOC_472/Y 0.00fF
C68369 NOR2X1_LOC_445/Y INVX1_LOC_29/A 0.01fF
C68370 INVX1_LOC_63/Y NAND2X1_LOC_74/B 0.02fF
C68371 INVX1_LOC_10/A INVX1_LOC_157/Y 0.03fF
C68372 NAND2X1_LOC_728/Y INVX1_LOC_231/A 0.01fF
C68373 NOR2X1_LOC_68/A NAND2X1_LOC_278/a_36_24# 0.06fF
C68374 INVX1_LOC_286/A INVX1_LOC_93/Y 0.18fF
C68375 INVX1_LOC_2/A NAND2X1_LOC_489/Y 0.03fF
C68376 NOR2X1_LOC_643/Y NAND2X1_LOC_214/a_36_24# 0.00fF
C68377 INVX1_LOC_39/A NOR2X1_LOC_293/a_36_216# 0.00fF
C68378 NOR2X1_LOC_82/A NAND2X1_LOC_205/A 0.01fF
C68379 NAND2X1_LOC_348/A VDD 0.83fF
C68380 NOR2X1_LOC_655/B INVX1_LOC_63/A 0.11fF
C68381 NAND2X1_LOC_563/A NOR2X1_LOC_649/B 0.02fF
C68382 INVX1_LOC_58/A NOR2X1_LOC_457/A 0.07fF
C68383 NOR2X1_LOC_246/A INVX1_LOC_118/A 0.48fF
C68384 INVX1_LOC_113/Y NOR2X1_LOC_477/B 0.01fF
C68385 NAND2X1_LOC_563/A INVX1_LOC_3/A 0.16fF
C68386 NOR2X1_LOC_716/B NOR2X1_LOC_159/a_36_216# 0.00fF
C68387 INVX1_LOC_43/Y INVX1_LOC_57/A 0.03fF
C68388 NOR2X1_LOC_441/Y NOR2X1_LOC_65/Y 0.65fF
C68389 NAND2X1_LOC_579/A NOR2X1_LOC_109/Y 0.03fF
C68390 NAND2X1_LOC_850/Y NOR2X1_LOC_662/A 0.02fF
C68391 NAND2X1_LOC_551/A INVX1_LOC_118/A 0.01fF
C68392 INVX1_LOC_49/A INVX1_LOC_32/A 0.10fF
C68393 NOR2X1_LOC_175/A NAND2X1_LOC_74/B 0.10fF
C68394 NAND2X1_LOC_550/A NOR2X1_LOC_754/Y 0.02fF
C68395 INVX1_LOC_93/Y INVX1_LOC_95/A 0.13fF
C68396 INVX1_LOC_224/Y INVX1_LOC_170/A 0.01fF
C68397 NOR2X1_LOC_255/Y NAND2X1_LOC_208/B 0.01fF
C68398 NOR2X1_LOC_552/A NAND2X1_LOC_447/Y 0.46fF
C68399 NOR2X1_LOC_137/A NOR2X1_LOC_831/B 0.77fF
C68400 INVX1_LOC_159/Y INVX1_LOC_76/A 0.03fF
C68401 INVX1_LOC_32/Y NOR2X1_LOC_257/Y 0.08fF
C68402 INVX1_LOC_5/A NAND2X1_LOC_719/a_36_24# 0.00fF
C68403 NOR2X1_LOC_32/B INVX1_LOC_31/A 0.01fF
C68404 INVX1_LOC_58/A INVX1_LOC_30/A 0.39fF
C68405 NOR2X1_LOC_753/Y INVX1_LOC_94/Y 0.01fF
C68406 INVX1_LOC_223/A INVX1_LOC_29/Y 0.07fF
C68407 NAND2X1_LOC_35/Y NOR2X1_LOC_371/a_36_216# 0.01fF
C68408 INVX1_LOC_89/A NAND2X1_LOC_257/a_36_24# 0.00fF
C68409 INVX1_LOC_99/Y NOR2X1_LOC_794/B 0.01fF
C68410 NOR2X1_LOC_329/B INVX1_LOC_291/A 0.12fF
C68411 INVX1_LOC_49/A NAND2X1_LOC_175/Y 0.00fF
C68412 NOR2X1_LOC_303/Y INVX1_LOC_116/Y 0.01fF
C68413 NAND2X1_LOC_325/Y INVX1_LOC_94/Y 0.01fF
C68414 INVX1_LOC_35/A NOR2X1_LOC_844/Y 0.01fF
C68415 INVX1_LOC_266/Y D_INPUT_5 0.09fF
C68416 INVX1_LOC_21/A NOR2X1_LOC_250/Y 0.18fF
C68417 NOR2X1_LOC_516/B INVX1_LOC_69/A 0.01fF
C68418 INVX1_LOC_13/A NAND2X1_LOC_63/Y 0.10fF
C68419 NAND2X1_LOC_391/Y NAND2X1_LOC_793/Y 0.00fF
C68420 NOR2X1_LOC_151/Y NOR2X1_LOC_676/a_36_216# 0.00fF
C68421 NOR2X1_LOC_99/B INVX1_LOC_63/A 0.07fF
C68422 INVX1_LOC_2/A INVX1_LOC_32/A 0.04fF
C68423 INVX1_LOC_24/A NOR2X1_LOC_748/A 0.41fF
C68424 NOR2X1_LOC_494/Y NAND2X1_LOC_561/B 0.08fF
C68425 NOR2X1_LOC_45/B INVX1_LOC_33/Y 0.03fF
C68426 INVX1_LOC_96/A INVX1_LOC_44/A 0.02fF
C68427 INVX1_LOC_35/A NOR2X1_LOC_769/A 0.06fF
C68428 NOR2X1_LOC_337/Y INVX1_LOC_38/A 0.03fF
C68429 NOR2X1_LOC_226/A INVX1_LOC_32/A 0.10fF
C68430 NOR2X1_LOC_121/A INVX1_LOC_42/A 0.06fF
C68431 INVX1_LOC_35/A NOR2X1_LOC_554/B 0.08fF
C68432 NAND2X1_LOC_714/B NOR2X1_LOC_816/A 0.09fF
C68433 NOR2X1_LOC_846/B INVX1_LOC_63/A 0.03fF
C68434 INVX1_LOC_34/A INVX1_LOC_26/A 0.18fF
C68435 INVX1_LOC_48/Y NOR2X1_LOC_530/a_36_216# 0.00fF
C68436 INPUT_1 NAND2X1_LOC_489/Y 0.03fF
C68437 NAND2X1_LOC_335/a_36_24# INVX1_LOC_4/Y 0.01fF
C68438 NOR2X1_LOC_843/A INVX1_LOC_26/Y 0.02fF
C68439 NOR2X1_LOC_78/A NOR2X1_LOC_331/B 0.07fF
C68440 NOR2X1_LOC_13/Y INVX1_LOC_53/A 0.03fF
C68441 NOR2X1_LOC_226/A NOR2X1_LOC_329/Y 0.21fF
C68442 INVX1_LOC_45/A NOR2X1_LOC_186/Y 0.14fF
C68443 NOR2X1_LOC_728/a_36_216# NOR2X1_LOC_155/A 0.00fF
C68444 INVX1_LOC_256/A INVX1_LOC_269/A 0.10fF
C68445 NAND2X1_LOC_510/a_36_24# NOR2X1_LOC_843/B 0.00fF
C68446 NOR2X1_LOC_478/A NAND2X1_LOC_149/Y 0.06fF
C68447 NOR2X1_LOC_720/B NOR2X1_LOC_668/Y 0.02fF
C68448 INVX1_LOC_88/A INVX1_LOC_150/Y 0.10fF
C68449 INVX1_LOC_287/Y NOR2X1_LOC_708/B 0.01fF
C68450 INVX1_LOC_230/Y NOR2X1_LOC_15/Y 0.03fF
C68451 NOR2X1_LOC_647/B INVX1_LOC_269/A 0.02fF
C68452 INVX1_LOC_2/A NAND2X1_LOC_175/Y 0.16fF
C68453 INVX1_LOC_182/A INVX1_LOC_63/A 0.07fF
C68454 NOR2X1_LOC_405/A INVX1_LOC_118/Y 0.02fF
C68455 NOR2X1_LOC_318/B INVX1_LOC_54/A 0.08fF
C68456 NAND2X1_LOC_807/Y NAND2X1_LOC_604/a_36_24# 0.01fF
C68457 NAND2X1_LOC_703/Y INVX1_LOC_141/Y 0.13fF
C68458 NOR2X1_LOC_817/Y NOR2X1_LOC_82/A 0.47fF
C68459 NAND2X1_LOC_773/Y NOR2X1_LOC_590/A 0.00fF
C68460 NOR2X1_LOC_596/A NOR2X1_LOC_665/Y 0.03fF
C68461 NOR2X1_LOC_56/Y INVX1_LOC_38/A 0.07fF
C68462 INVX1_LOC_35/A NOR2X1_LOC_152/Y 0.07fF
C68463 NOR2X1_LOC_220/B NOR2X1_LOC_360/Y 0.02fF
C68464 INVX1_LOC_136/A NOR2X1_LOC_496/Y 0.01fF
C68465 NOR2X1_LOC_273/Y INVX1_LOC_5/A 0.07fF
C68466 NOR2X1_LOC_226/A NAND2X1_LOC_175/Y 0.10fF
C68467 INVX1_LOC_45/A NAND2X1_LOC_573/Y 0.01fF
C68468 INVX1_LOC_54/Y INVX1_LOC_116/Y 0.00fF
C68469 NAND2X1_LOC_35/Y NOR2X1_LOC_403/B 0.01fF
C68470 INVX1_LOC_24/A NOR2X1_LOC_304/Y 0.16fF
C68471 NAND2X1_LOC_858/B INVX1_LOC_285/A 0.07fF
C68472 INVX1_LOC_5/A NOR2X1_LOC_759/Y 0.01fF
C68473 INVX1_LOC_166/A INVX1_LOC_194/A 0.38fF
C68474 NOR2X1_LOC_646/a_36_216# NOR2X1_LOC_38/B 0.00fF
C68475 NAND2X1_LOC_858/B INVX1_LOC_265/Y 0.00fF
C68476 NAND2X1_LOC_640/Y NAND2X1_LOC_793/B 0.02fF
C68477 INVX1_LOC_239/A INVX1_LOC_72/A 0.01fF
C68478 INVX1_LOC_166/A NOR2X1_LOC_399/A 0.16fF
C68479 INVX1_LOC_36/A NAND2X1_LOC_579/A 0.07fF
C68480 INVX1_LOC_41/A NOR2X1_LOC_678/A 0.03fF
C68481 INVX1_LOC_16/A NAND2X1_LOC_454/Y 0.10fF
C68482 NAND2X1_LOC_149/Y NOR2X1_LOC_68/A 0.09fF
C68483 NAND2X1_LOC_849/B VDD 0.46fF
C68484 NOR2X1_LOC_186/Y INVX1_LOC_71/A 0.17fF
C68485 INVX1_LOC_146/Y INVX1_LOC_38/A 0.05fF
C68486 INVX1_LOC_5/A NOR2X1_LOC_550/B 0.10fF
C68487 INVX1_LOC_114/A INVX1_LOC_37/A 0.01fF
C68488 VDD INVX1_LOC_38/A 2.24fF
C68489 NOR2X1_LOC_309/Y INVX1_LOC_308/A 0.03fF
C68490 NAND2X1_LOC_198/a_36_24# NOR2X1_LOC_103/Y 0.00fF
C68491 INVX1_LOC_305/A INVX1_LOC_24/Y 0.10fF
C68492 INVX1_LOC_58/A NAND2X1_LOC_722/A 0.02fF
C68493 INVX1_LOC_12/Y NOR2X1_LOC_536/A 0.01fF
C68494 INVX1_LOC_170/A NOR2X1_LOC_103/Y 0.02fF
C68495 INVX1_LOC_25/A INVX1_LOC_54/Y 0.10fF
C68496 NAND2X1_LOC_860/A NOR2X1_LOC_84/Y 0.20fF
C68497 VDD NOR2X1_LOC_96/Y 0.43fF
C68498 INVX1_LOC_139/A INVX1_LOC_54/A 0.04fF
C68499 NOR2X1_LOC_536/A NOR2X1_LOC_492/Y 0.01fF
C68500 INVX1_LOC_73/Y INVX1_LOC_72/A 0.01fF
C68501 INVX1_LOC_177/A NOR2X1_LOC_493/a_36_216# 0.00fF
C68502 NAND2X1_LOC_573/Y INVX1_LOC_71/A 0.10fF
C68503 INPUT_1 INVX1_LOC_32/A 0.11fF
C68504 NOR2X1_LOC_669/Y INVX1_LOC_24/A 0.42fF
C68505 NOR2X1_LOC_298/Y NOR2X1_LOC_409/B 0.03fF
C68506 NOR2X1_LOC_242/A NAND2X1_LOC_364/Y 0.03fF
C68507 NAND2X1_LOC_218/B NAND2X1_LOC_218/A 0.11fF
C68508 NOR2X1_LOC_510/Y NOR2X1_LOC_172/Y 0.45fF
C68509 NOR2X1_LOC_690/A NOR2X1_LOC_291/Y 0.02fF
C68510 NOR2X1_LOC_335/B INVX1_LOC_29/A 0.77fF
C68511 NOR2X1_LOC_331/B NOR2X1_LOC_60/Y 0.01fF
C68512 INPUT_5 NOR2X1_LOC_25/Y 0.03fF
C68513 INVX1_LOC_208/A INVX1_LOC_270/Y 0.02fF
C68514 VDD NOR2X1_LOC_51/A 0.42fF
C68515 NAND2X1_LOC_721/A INVX1_LOC_54/A 0.07fF
C68516 INVX1_LOC_25/Y NAND2X1_LOC_464/B 0.07fF
C68517 NAND2X1_LOC_112/Y NOR2X1_LOC_106/a_36_216# 0.00fF
C68518 NAND2X1_LOC_331/a_36_24# INVX1_LOC_94/Y 0.00fF
C68519 INVX1_LOC_1/A NOR2X1_LOC_303/Y 0.01fF
C68520 NOR2X1_LOC_639/B INVX1_LOC_191/Y 0.00fF
C68521 D_INPUT_1 INVX1_LOC_56/A 0.08fF
C68522 VDD NAND2X1_LOC_848/Y -0.00fF
C68523 INVX1_LOC_37/A INVX1_LOC_307/A 0.07fF
C68524 NOR2X1_LOC_645/a_36_216# NOR2X1_LOC_816/A 0.00fF
C68525 INVX1_LOC_12/Y NAND2X1_LOC_93/B 0.10fF
C68526 INVX1_LOC_5/A NOR2X1_LOC_41/Y 0.01fF
C68527 INVX1_LOC_50/A NOR2X1_LOC_561/Y 0.11fF
C68528 NAND2X1_LOC_538/Y NOR2X1_LOC_577/Y 0.01fF
C68529 INVX1_LOC_37/A NOR2X1_LOC_445/B 0.10fF
C68530 INVX1_LOC_27/A NOR2X1_LOC_300/Y 0.08fF
C68531 INVX1_LOC_27/A NOR2X1_LOC_87/B 0.04fF
C68532 NOR2X1_LOC_798/A NOR2X1_LOC_168/B 0.02fF
C68533 INVX1_LOC_28/A NAND2X1_LOC_454/Y 0.01fF
C68534 INVX1_LOC_83/A NOR2X1_LOC_727/B 0.01fF
C68535 INVX1_LOC_45/Y INVX1_LOC_292/A 0.03fF
C68536 INVX1_LOC_135/A INVX1_LOC_112/Y 0.03fF
C68537 NOR2X1_LOC_439/B NOR2X1_LOC_334/Y 0.00fF
C68538 NOR2X1_LOC_689/Y NAND2X1_LOC_691/a_36_24# 0.00fF
C68539 INVX1_LOC_1/A NOR2X1_LOC_84/A 0.03fF
C68540 NOR2X1_LOC_250/A NOR2X1_LOC_577/Y 0.01fF
C68541 NOR2X1_LOC_32/B NAND2X1_LOC_859/Y 0.18fF
C68542 NOR2X1_LOC_328/Y NOR2X1_LOC_53/Y 0.01fF
C68543 INVX1_LOC_75/A NOR2X1_LOC_334/Y 0.18fF
C68544 INVX1_LOC_27/A NAND2X1_LOC_360/B 0.14fF
C68545 INVX1_LOC_191/A D_INPUT_5 0.01fF
C68546 NAND2X1_LOC_562/B NAND2X1_LOC_561/B 0.02fF
C68547 NAND2X1_LOC_357/B INVX1_LOC_14/A 0.07fF
C68548 INVX1_LOC_95/Y NOR2X1_LOC_77/a_36_216# 0.01fF
C68549 INVX1_LOC_54/A INVX1_LOC_117/Y 0.03fF
C68550 NAND2X1_LOC_738/B INVX1_LOC_173/Y 1.23fF
C68551 INVX1_LOC_54/Y INVX1_LOC_1/A 0.10fF
C68552 NOR2X1_LOC_721/Y NAND2X1_LOC_223/A 0.44fF
C68553 INVX1_LOC_224/A NAND2X1_LOC_114/a_36_24# 0.00fF
C68554 NOR2X1_LOC_794/B NOR2X1_LOC_254/Y 0.00fF
C68555 NOR2X1_LOC_176/Y INVX1_LOC_63/A 0.08fF
C68556 NOR2X1_LOC_9/Y NOR2X1_LOC_248/A 0.03fF
C68557 INVX1_LOC_239/Y INVX1_LOC_242/A 0.03fF
C68558 INVX1_LOC_53/Y NAND2X1_LOC_474/Y 1.56fF
C68559 INVX1_LOC_298/Y NOR2X1_LOC_335/B 0.02fF
C68560 INVX1_LOC_14/A NAND2X1_LOC_549/B 0.01fF
C68561 INVX1_LOC_39/A INVX1_LOC_13/A 0.12fF
C68562 INPUT_0 INVX1_LOC_26/A 0.13fF
C68563 D_INPUT_7 INVX1_LOC_77/A 0.03fF
C68564 INVX1_LOC_126/A INVX1_LOC_102/A 0.06fF
C68565 NOR2X1_LOC_481/A INVX1_LOC_45/A 0.37fF
C68566 INVX1_LOC_286/A INVX1_LOC_87/A 0.71fF
C68567 NOR2X1_LOC_720/B INVX1_LOC_31/A 0.01fF
C68568 NAND2X1_LOC_563/Y NAND2X1_LOC_555/Y 0.01fF
C68569 INVX1_LOC_160/Y NOR2X1_LOC_852/Y 0.02fF
C68570 INVX1_LOC_12/A INVX1_LOC_37/A 0.11fF
C68571 NAND2X1_LOC_738/B NOR2X1_LOC_385/Y 0.00fF
C68572 INVX1_LOC_83/A NOR2X1_LOC_649/Y 0.09fF
C68573 INVX1_LOC_230/Y INVX1_LOC_15/Y 0.03fF
C68574 INVX1_LOC_45/A INVX1_LOC_225/A 0.80fF
C68575 INVX1_LOC_136/A INVX1_LOC_63/Y 0.01fF
C68576 INPUT_3 NOR2X1_LOC_818/Y 0.52fF
C68577 INVX1_LOC_41/A INVX1_LOC_305/A 0.07fF
C68578 NOR2X1_LOC_67/A INVX1_LOC_293/A 0.01fF
C68579 NAND2X1_LOC_739/B NOR2X1_LOC_387/Y 0.01fF
C68580 INVX1_LOC_225/A NOR2X1_LOC_568/A 0.01fF
C68581 NOR2X1_LOC_697/Y INVX1_LOC_92/A 0.03fF
C68582 NAND2X1_LOC_796/B INVX1_LOC_135/A 0.01fF
C68583 INVX1_LOC_21/A D_INPUT_0 15.90fF
C68584 NOR2X1_LOC_827/a_36_216# INVX1_LOC_22/Y 0.00fF
C68585 INVX1_LOC_159/A INVX1_LOC_33/A 0.07fF
C68586 INVX1_LOC_50/A NOR2X1_LOC_167/Y 0.81fF
C68587 NOR2X1_LOC_815/A INVX1_LOC_271/A 0.05fF
C68588 NOR2X1_LOC_419/Y INVX1_LOC_314/Y 0.04fF
C68589 NOR2X1_LOC_78/A NOR2X1_LOC_621/B 0.01fF
C68590 NAND2X1_LOC_35/Y NOR2X1_LOC_497/Y 0.05fF
C68591 INVX1_LOC_34/A NOR2X1_LOC_276/B 0.00fF
C68592 NAND2X1_LOC_721/A NOR2X1_LOC_48/B 0.15fF
C68593 NOR2X1_LOC_78/A NOR2X1_LOC_449/A 0.01fF
C68594 INVX1_LOC_185/A NOR2X1_LOC_605/A 0.01fF
C68595 NOR2X1_LOC_510/Y INVX1_LOC_90/A 0.04fF
C68596 NOR2X1_LOC_441/Y NOR2X1_LOC_362/a_36_216# 0.00fF
C68597 NOR2X1_LOC_363/Y INVX1_LOC_290/Y 0.05fF
C68598 NOR2X1_LOC_45/B INVX1_LOC_23/Y 0.04fF
C68599 NOR2X1_LOC_637/B NAND2X1_LOC_593/Y 0.02fF
C68600 NOR2X1_LOC_481/A INVX1_LOC_71/A 0.05fF
C68601 NOR2X1_LOC_716/B INVX1_LOC_314/Y 0.23fF
C68602 INVX1_LOC_45/A NOR2X1_LOC_209/Y 0.08fF
C68603 NAND2X1_LOC_640/Y INVX1_LOC_71/A 0.06fF
C68604 INVX1_LOC_14/A NOR2X1_LOC_128/B 0.02fF
C68605 INVX1_LOC_1/A NAND2X1_LOC_125/a_36_24# 0.00fF
C68606 NAND2X1_LOC_30/Y GATE_662 0.01fF
C68607 NOR2X1_LOC_658/Y NOR2X1_LOC_78/B 0.07fF
C68608 INVX1_LOC_188/A INVX1_LOC_263/A -0.00fF
C68609 NAND2X1_LOC_149/Y NOR2X1_LOC_163/A 0.02fF
C68610 INVX1_LOC_174/A NAND2X1_LOC_149/B 0.03fF
C68611 INVX1_LOC_225/A INVX1_LOC_71/A 0.11fF
C68612 NOR2X1_LOC_561/Y NAND2X1_LOC_227/Y 0.01fF
C68613 INVX1_LOC_119/A INVX1_LOC_24/A 0.25fF
C68614 INVX1_LOC_128/Y INVX1_LOC_46/A 0.01fF
C68615 INVX1_LOC_192/A INVX1_LOC_77/A 0.03fF
C68616 INVX1_LOC_59/Y INVX1_LOC_16/Y 0.10fF
C68617 NAND2X1_LOC_374/Y INVX1_LOC_18/A 0.07fF
C68618 NAND2X1_LOC_213/A D_GATE_366 0.07fF
C68619 NOR2X1_LOC_639/B INVX1_LOC_6/A 0.15fF
C68620 NOR2X1_LOC_804/B NOR2X1_LOC_551/B 0.10fF
C68621 NAND2X1_LOC_784/A NOR2X1_LOC_528/Y 0.01fF
C68622 VDD NAND2X1_LOC_223/A 0.34fF
C68623 NAND2X1_LOC_580/a_36_24# NOR2X1_LOC_298/Y 0.07fF
C68624 INVX1_LOC_224/Y NAND2X1_LOC_642/Y 0.01fF
C68625 NAND2X1_LOC_714/B INVX1_LOC_140/A 1.70fF
C68626 INVX1_LOC_235/Y NAND2X1_LOC_462/a_36_24# 0.01fF
C68627 INVX1_LOC_33/A NOR2X1_LOC_542/a_36_216# 0.00fF
C68628 NOR2X1_LOC_361/B INVX1_LOC_90/A 0.05fF
C68629 INVX1_LOC_36/A INVX1_LOC_208/Y 0.01fF
C68630 NAND2X1_LOC_724/Y INVX1_LOC_11/Y 0.03fF
C68631 NOR2X1_LOC_357/Y NOR2X1_LOC_631/Y 0.15fF
C68632 NOR2X1_LOC_229/a_36_216# INVX1_LOC_72/A 0.00fF
C68633 VDD INVX1_LOC_18/Y 0.21fF
C68634 NOR2X1_LOC_590/A INVX1_LOC_279/A 0.07fF
C68635 NOR2X1_LOC_802/A INVX1_LOC_77/A 0.08fF
C68636 NOR2X1_LOC_15/Y NOR2X1_LOC_153/a_36_216# 0.00fF
C68637 NOR2X1_LOC_336/B NOR2X1_LOC_748/Y 0.00fF
C68638 INVX1_LOC_49/A INVX1_LOC_158/A 0.01fF
C68639 NAND2X1_LOC_213/A NAND2X1_LOC_162/a_36_24# 0.00fF
C68640 NOR2X1_LOC_246/A NAND2X1_LOC_352/a_36_24# 0.01fF
C68641 NOR2X1_LOC_361/B NOR2X1_LOC_389/B 0.43fF
C68642 NOR2X1_LOC_209/Y INVX1_LOC_71/A 0.03fF
C68643 NOR2X1_LOC_773/Y INVX1_LOC_300/Y 0.00fF
C68644 NOR2X1_LOC_296/Y INPUT_1 0.16fF
C68645 NOR2X1_LOC_78/B NOR2X1_LOC_13/Y 0.17fF
C68646 INVX1_LOC_32/A INVX1_LOC_118/A 0.10fF
C68647 NOR2X1_LOC_447/Y INVX1_LOC_191/Y 0.00fF
C68648 INVX1_LOC_223/A INVX1_LOC_101/A 0.04fF
C68649 NOR2X1_LOC_15/Y NAND2X1_LOC_740/B 0.05fF
C68650 NOR2X1_LOC_68/A INVX1_LOC_16/A 0.02fF
C68651 INVX1_LOC_59/Y NAND2X1_LOC_205/A 0.00fF
C68652 NOR2X1_LOC_321/Y INVX1_LOC_79/A 0.03fF
C68653 INVX1_LOC_112/A NAND2X1_LOC_205/A 0.10fF
C68654 INVX1_LOC_50/A INVX1_LOC_76/A 5.48fF
C68655 NAND2X1_LOC_424/a_36_24# INVX1_LOC_46/A 0.01fF
C68656 NOR2X1_LOC_740/a_36_216# INVX1_LOC_85/Y 0.00fF
C68657 INVX1_LOC_172/A NAND2X1_LOC_374/Y 0.07fF
C68658 NOR2X1_LOC_329/Y INVX1_LOC_118/A 0.07fF
C68659 INVX1_LOC_27/Y NAND2X1_LOC_74/B 0.04fF
C68660 INPUT_3 INPUT_1 0.04fF
C68661 NOR2X1_LOC_78/B NAND2X1_LOC_364/Y 0.07fF
C68662 INVX1_LOC_298/A INVX1_LOC_91/A 0.01fF
C68663 INVX1_LOC_215/A NAND2X1_LOC_514/Y 0.04fF
C68664 INVX1_LOC_145/A INVX1_LOC_208/Y 0.00fF
C68665 INVX1_LOC_270/Y NAND2X1_LOC_211/Y 0.02fF
C68666 NOR2X1_LOC_789/B INVX1_LOC_48/A 0.04fF
C68667 NOR2X1_LOC_553/Y INVX1_LOC_94/A 0.00fF
C68668 INVX1_LOC_84/A INVX1_LOC_29/A 0.28fF
C68669 NOR2X1_LOC_361/B NAND2X1_LOC_348/A 0.00fF
C68670 INVX1_LOC_223/A NOR2X1_LOC_355/A 1.40fF
C68671 NOR2X1_LOC_392/B INVX1_LOC_177/A 0.01fF
C68672 NOR2X1_LOC_634/A INVX1_LOC_15/A 0.03fF
C68673 NOR2X1_LOC_865/a_36_216# NOR2X1_LOC_865/Y 0.02fF
C68674 INVX1_LOC_41/A NOR2X1_LOC_191/A 0.03fF
C68675 NOR2X1_LOC_224/Y INVX1_LOC_76/A 0.07fF
C68676 NAND2X1_LOC_175/Y INVX1_LOC_118/A 0.10fF
C68677 NAND2X1_LOC_198/B INVX1_LOC_10/A 0.02fF
C68678 NAND2X1_LOC_297/a_36_24# NAND2X1_LOC_99/A 0.00fF
C68679 INVX1_LOC_1/A NOR2X1_LOC_354/Y 0.01fF
C68680 NOR2X1_LOC_380/a_36_216# NAND2X1_LOC_560/A 0.00fF
C68681 INVX1_LOC_269/A INVX1_LOC_69/Y 0.18fF
C68682 INVX1_LOC_46/A NOR2X1_LOC_717/A 0.17fF
C68683 NOR2X1_LOC_19/B NAND2X1_LOC_104/a_36_24# 0.00fF
C68684 NAND2X1_LOC_368/a_36_24# INVX1_LOC_10/A 0.00fF
C68685 NAND2X1_LOC_364/A NOR2X1_LOC_333/A 0.11fF
C68686 NOR2X1_LOC_554/A NOR2X1_LOC_649/B 0.03fF
C68687 NAND2X1_LOC_651/B INVX1_LOC_29/A 0.27fF
C68688 NOR2X1_LOC_107/Y INPUT_0 0.01fF
C68689 NOR2X1_LOC_820/Y INVX1_LOC_4/A 0.08fF
C68690 NOR2X1_LOC_554/A INVX1_LOC_3/A 0.03fF
C68691 INVX1_LOC_280/A INVX1_LOC_112/Y 0.05fF
C68692 NOR2X1_LOC_321/Y INVX1_LOC_91/A 0.01fF
C68693 INVX1_LOC_49/A GATE_662 0.46fF
C68694 NOR2X1_LOC_795/Y NOR2X1_LOC_284/B 0.45fF
C68695 NOR2X1_LOC_13/Y INVX1_LOC_83/A 0.10fF
C68696 NOR2X1_LOC_142/Y INVX1_LOC_1/Y 0.01fF
C68697 INVX1_LOC_245/Y INVX1_LOC_311/A 0.01fF
C68698 INVX1_LOC_20/A INVX1_LOC_306/Y 0.05fF
C68699 NOR2X1_LOC_82/A INVX1_LOC_286/A 0.07fF
C68700 INVX1_LOC_24/A INVX1_LOC_89/A 0.33fF
C68701 NAND2X1_LOC_72/B NOR2X1_LOC_445/B 0.04fF
C68702 INVX1_LOC_215/A NAND2X1_LOC_332/Y 0.03fF
C68703 NAND2X1_LOC_527/a_36_24# INVX1_LOC_158/Y 0.00fF
C68704 NOR2X1_LOC_590/A NAND2X1_LOC_858/B 0.00fF
C68705 NOR2X1_LOC_68/A INVX1_LOC_28/A 0.26fF
C68706 NOR2X1_LOC_718/B NOR2X1_LOC_302/B 0.05fF
C68707 NOR2X1_LOC_359/Y INVX1_LOC_313/Y 0.00fF
C68708 NAND2X1_LOC_208/B NOR2X1_LOC_368/A 0.06fF
C68709 NOR2X1_LOC_78/B INVX1_LOC_256/Y 0.15fF
C68710 NOR2X1_LOC_848/Y NOR2X1_LOC_78/A 0.00fF
C68711 INVX1_LOC_245/A NOR2X1_LOC_423/Y 0.00fF
C68712 NOR2X1_LOC_106/A NOR2X1_LOC_577/Y 0.00fF
C68713 NOR2X1_LOC_709/A INVX1_LOC_22/A 0.12fF
C68714 INVX1_LOC_19/A D_INPUT_5 0.00fF
C68715 INVX1_LOC_2/A INVX1_LOC_9/Y 0.06fF
C68716 INVX1_LOC_132/A NOR2X1_LOC_749/Y 0.01fF
C68717 NAND2X1_LOC_574/A NOR2X1_LOC_34/Y 0.06fF
C68718 NOR2X1_LOC_669/A NOR2X1_LOC_48/B 0.03fF
C68719 NOR2X1_LOC_11/Y D_INPUT_5 0.03fF
C68720 NAND2X1_LOC_63/Y INVX1_LOC_32/A 0.03fF
C68721 INVX1_LOC_2/A NAND2X1_LOC_564/B 0.07fF
C68722 NOR2X1_LOC_103/Y NAND2X1_LOC_642/Y 0.00fF
C68723 NOR2X1_LOC_522/Y NAND2X1_LOC_849/A 0.01fF
C68724 NOR2X1_LOC_655/B INVX1_LOC_1/Y 0.01fF
C68725 NAND2X1_LOC_308/Y NAND2X1_LOC_691/a_36_24# 0.00fF
C68726 INVX1_LOC_89/A NOR2X1_LOC_557/Y 0.03fF
C68727 INVX1_LOC_29/A INVX1_LOC_15/A 4.07fF
C68728 NAND2X1_LOC_360/B INVX1_LOC_137/A 0.24fF
C68729 NOR2X1_LOC_831/B NOR2X1_LOC_383/B 0.03fF
C68730 INVX1_LOC_25/A NOR2X1_LOC_78/Y 0.10fF
C68731 NOR2X1_LOC_82/A INVX1_LOC_95/A 0.00fF
C68732 INVX1_LOC_298/Y INVX1_LOC_84/A 0.02fF
C68733 NOR2X1_LOC_226/A NAND2X1_LOC_564/B 1.34fF
C68734 NOR2X1_LOC_197/B NOR2X1_LOC_748/A 0.04fF
C68735 INVX1_LOC_271/A NAND2X1_LOC_436/a_36_24# 0.00fF
C68736 INVX1_LOC_53/A NOR2X1_LOC_640/Y 0.18fF
C68737 INVX1_LOC_256/A NOR2X1_LOC_275/A 0.01fF
C68738 D_INPUT_1 NOR2X1_LOC_155/A 0.08fF
C68739 INVX1_LOC_119/A NOR2X1_LOC_130/A 0.02fF
C68740 NOR2X1_LOC_441/Y NOR2X1_LOC_318/B 0.01fF
C68741 INVX1_LOC_58/A INVX1_LOC_113/A 0.06fF
C68742 NOR2X1_LOC_510/Y INVX1_LOC_38/A 0.34fF
C68743 INVX1_LOC_256/Y NAND2X1_LOC_392/Y 0.02fF
C68744 INVX1_LOC_226/Y NOR2X1_LOC_619/A 0.20fF
C68745 INVX1_LOC_21/A NAND2X1_LOC_848/A 0.01fF
C68746 INVX1_LOC_190/Y NAND2X1_LOC_466/A 0.08fF
C68747 INVX1_LOC_90/A INVX1_LOC_121/Y 0.01fF
C68748 NOR2X1_LOC_772/B NOR2X1_LOC_612/Y 0.03fF
C68749 INVX1_LOC_47/A INVX1_LOC_104/A 0.03fF
C68750 NAND2X1_LOC_741/B NOR2X1_LOC_45/B 0.02fF
C68751 NOR2X1_LOC_20/Y VDD 0.24fF
C68752 NAND2X1_LOC_454/Y INVX1_LOC_109/A 0.01fF
C68753 NOR2X1_LOC_303/Y NOR2X1_LOC_188/A 0.11fF
C68754 NOR2X1_LOC_717/B NOR2X1_LOC_778/B 0.61fF
C68755 INVX1_LOC_26/A NOR2X1_LOC_84/B 0.05fF
C68756 NOR2X1_LOC_471/Y INVX1_LOC_115/A 0.01fF
C68757 INVX1_LOC_200/A INVX1_LOC_37/A 0.07fF
C68758 INVX1_LOC_45/A NAND2X1_LOC_642/Y 0.06fF
C68759 NOR2X1_LOC_667/A D_INPUT_0 0.08fF
C68760 INVX1_LOC_90/A INVX1_LOC_177/A 0.03fF
C68761 INVX1_LOC_248/A D_INPUT_0 0.07fF
C68762 NOR2X1_LOC_15/Y INVX1_LOC_44/A 0.07fF
C68763 INVX1_LOC_53/A NOR2X1_LOC_697/Y 0.06fF
C68764 NOR2X1_LOC_162/Y INVX1_LOC_75/A 0.00fF
C68765 INVX1_LOC_89/A INVX1_LOC_143/A 0.09fF
C68766 INVX1_LOC_53/Y INVX1_LOC_10/A 0.03fF
C68767 INVX1_LOC_90/A NAND2X1_LOC_630/a_36_24# 0.01fF
C68768 INVX1_LOC_61/Y INVX1_LOC_76/A 0.12fF
C68769 NOR2X1_LOC_483/B VDD 0.02fF
C68770 NOR2X1_LOC_778/B NOR2X1_LOC_828/A 0.05fF
C68771 NOR2X1_LOC_607/A INVX1_LOC_91/A 0.02fF
C68772 NOR2X1_LOC_718/B INVX1_LOC_75/A 0.07fF
C68773 NOR2X1_LOC_151/Y NOR2X1_LOC_181/Y 0.07fF
C68774 INVX1_LOC_83/A NOR2X1_LOC_146/Y 0.12fF
C68775 NOR2X1_LOC_361/B INVX1_LOC_38/A 3.22fF
C68776 NOR2X1_LOC_155/A NOR2X1_LOC_652/Y 0.03fF
C68777 INVX1_LOC_10/A NOR2X1_LOC_665/A 0.10fF
C68778 NOR2X1_LOC_392/Y NAND2X1_LOC_206/Y 0.10fF
C68779 NOR2X1_LOC_541/a_36_216# INVX1_LOC_149/Y 0.00fF
C68780 INVX1_LOC_299/A NOR2X1_LOC_729/A 0.03fF
C68781 INVX1_LOC_21/A INVX1_LOC_46/Y 2.53fF
C68782 NOR2X1_LOC_125/a_36_216# INVX1_LOC_272/A 0.01fF
C68783 NOR2X1_LOC_13/Y NOR2X1_LOC_311/Y 0.00fF
C68784 NAND2X1_LOC_731/Y NAND2X1_LOC_729/B 0.30fF
C68785 NOR2X1_LOC_518/Y NOR2X1_LOC_164/Y 0.18fF
C68786 INVX1_LOC_289/Y INVX1_LOC_54/A 0.03fF
C68787 NOR2X1_LOC_103/Y NOR2X1_LOC_271/Y 0.01fF
C68788 NOR2X1_LOC_419/Y NOR2X1_LOC_557/A 0.00fF
C68789 NOR2X1_LOC_364/Y INVX1_LOC_6/A 0.01fF
C68790 NAND2X1_LOC_550/A NOR2X1_LOC_536/A 0.07fF
C68791 INVX1_LOC_191/Y INVX1_LOC_302/A 0.01fF
C68792 NAND2X1_LOC_63/Y NOR2X1_LOC_622/A 0.06fF
C68793 INVX1_LOC_71/A NAND2X1_LOC_642/Y 0.11fF
C68794 INVX1_LOC_33/A NOR2X1_LOC_337/Y 0.01fF
C68795 NOR2X1_LOC_68/A NOR2X1_LOC_35/Y 0.03fF
C68796 NOR2X1_LOC_160/B NOR2X1_LOC_536/A 4.38fF
C68797 NOR2X1_LOC_272/Y INVX1_LOC_123/Y 0.02fF
C68798 NAND2X1_LOC_564/B INPUT_1 0.07fF
C68799 NOR2X1_LOC_716/B NOR2X1_LOC_557/A 0.59fF
C68800 INVX1_LOC_298/Y INVX1_LOC_15/A 0.03fF
C68801 NOR2X1_LOC_590/A NOR2X1_LOC_98/B 0.00fF
C68802 INVX1_LOC_54/Y NOR2X1_LOC_188/A 0.04fF
C68803 NOR2X1_LOC_33/Y INVX1_LOC_15/A 0.01fF
C68804 INVX1_LOC_108/Y INVX1_LOC_29/A 0.13fF
C68805 NOR2X1_LOC_45/Y NOR2X1_LOC_331/B 0.08fF
C68806 NOR2X1_LOC_788/B INVX1_LOC_220/Y 0.16fF
C68807 NOR2X1_LOC_82/A INVX1_LOC_54/A 0.06fF
C68808 NOR2X1_LOC_420/a_36_216# INVX1_LOC_63/A 0.01fF
C68809 NOR2X1_LOC_379/a_36_216# INVX1_LOC_91/A 0.00fF
C68810 INVX1_LOC_278/A INVX1_LOC_29/A 0.07fF
C68811 NOR2X1_LOC_608/a_36_216# NAND2X1_LOC_348/A 0.00fF
C68812 NOR2X1_LOC_142/Y NOR2X1_LOC_318/B 0.10fF
C68813 NAND2X1_LOC_355/Y INVX1_LOC_37/A 0.02fF
C68814 INVX1_LOC_24/A NAND2X1_LOC_244/A 0.28fF
C68815 INVX1_LOC_90/A NAND2X1_LOC_573/A 0.01fF
C68816 INVX1_LOC_290/Y INVX1_LOC_29/Y 0.14fF
C68817 NAND2X1_LOC_214/B NAND2X1_LOC_219/B 0.15fF
C68818 INVX1_LOC_88/A NOR2X1_LOC_58/a_36_216# 0.00fF
C68819 NOR2X1_LOC_660/Y NAND2X1_LOC_83/a_36_24# 0.01fF
C68820 NOR2X1_LOC_663/A NAND2X1_LOC_82/Y 0.04fF
C68821 INVX1_LOC_89/A NOR2X1_LOC_130/A 0.03fF
C68822 NOR2X1_LOC_152/a_36_216# INVX1_LOC_76/A 0.00fF
C68823 NAND2X1_LOC_863/A INVX1_LOC_22/A 0.07fF
C68824 NOR2X1_LOC_160/B NOR2X1_LOC_655/Y 1.19fF
C68825 NOR2X1_LOC_147/B INVX1_LOC_65/A 0.02fF
C68826 NOR2X1_LOC_717/B NOR2X1_LOC_724/Y 0.05fF
C68827 NOR2X1_LOC_13/Y INVX1_LOC_46/A 0.08fF
C68828 INVX1_LOC_105/A INVX1_LOC_76/A 0.49fF
C68829 NOR2X1_LOC_561/Y NAND2X1_LOC_652/Y 0.03fF
C68830 INVX1_LOC_5/A NAND2X1_LOC_74/B 0.20fF
C68831 INVX1_LOC_5/A NAND2X1_LOC_207/Y 0.16fF
C68832 NOR2X1_LOC_523/A NOR2X1_LOC_243/B 0.04fF
C68833 NOR2X1_LOC_160/B NAND2X1_LOC_93/B 0.13fF
C68834 INVX1_LOC_75/A NOR2X1_LOC_569/Y 0.07fF
C68835 NOR2X1_LOC_679/B INVX1_LOC_76/A 0.01fF
C68836 INVX1_LOC_227/A INVX1_LOC_182/Y -0.04fF
C68837 NOR2X1_LOC_843/a_36_216# INVX1_LOC_15/A 0.01fF
C68838 INVX1_LOC_209/Y NAND2X1_LOC_453/A 0.14fF
C68839 NOR2X1_LOC_392/B NOR2X1_LOC_137/B 0.01fF
C68840 INVX1_LOC_104/A INVX1_LOC_95/Y 0.20fF
C68841 NOR2X1_LOC_589/A NOR2X1_LOC_74/A 1.03fF
C68842 NOR2X1_LOC_655/B NOR2X1_LOC_318/B 0.10fF
C68843 NAND2X1_LOC_466/A NOR2X1_LOC_56/Y 0.03fF
C68844 NOR2X1_LOC_828/A NOR2X1_LOC_724/Y 0.02fF
C68845 NOR2X1_LOC_160/B NAND2X1_LOC_425/Y 0.01fF
C68846 INVX1_LOC_33/A VDD 2.20fF
C68847 INVX1_LOC_162/Y INVX1_LOC_126/A 0.17fF
C68848 INVX1_LOC_77/A NOR2X1_LOC_363/Y 0.01fF
C68849 NOR2X1_LOC_142/Y INVX1_LOC_139/A 0.00fF
C68850 INVX1_LOC_138/A INVX1_LOC_32/A 0.04fF
C68851 NOR2X1_LOC_392/Y NOR2X1_LOC_297/A 0.02fF
C68852 INVX1_LOC_164/A INPUT_0 0.06fF
C68853 NOR2X1_LOC_614/Y INVX1_LOC_186/A 0.03fF
C68854 INVX1_LOC_135/A NAND2X1_LOC_840/Y 0.01fF
C68855 NOR2X1_LOC_655/B INVX1_LOC_93/Y 0.10fF
C68856 INVX1_LOC_71/A NOR2X1_LOC_271/Y 0.03fF
C68857 NOR2X1_LOC_160/B NOR2X1_LOC_649/B 0.12fF
C68858 NOR2X1_LOC_456/Y INVX1_LOC_78/A 0.08fF
C68859 NOR2X1_LOC_391/Y NOR2X1_LOC_719/B 0.18fF
C68860 NOR2X1_LOC_389/A INVX1_LOC_285/A 0.00fF
C68861 NOR2X1_LOC_160/B INVX1_LOC_3/A 0.04fF
C68862 NOR2X1_LOC_520/B NAND2X1_LOC_96/A 0.47fF
C68863 NAND2X1_LOC_714/B INVX1_LOC_42/A 0.03fF
C68864 NOR2X1_LOC_91/Y NAND2X1_LOC_444/a_36_24# 0.00fF
C68865 INVX1_LOC_171/A NOR2X1_LOC_74/A 0.03fF
C68866 NOR2X1_LOC_151/Y NOR2X1_LOC_724/Y 1.97fF
C68867 NAND2X1_LOC_798/A NOR2X1_LOC_56/Y 0.01fF
C68868 NAND2X1_LOC_139/A NOR2X1_LOC_813/Y 0.04fF
C68869 INVX1_LOC_304/Y INVX1_LOC_37/A 0.04fF
C68870 NOR2X1_LOC_135/Y NOR2X1_LOC_329/B 0.09fF
C68871 INVX1_LOC_14/A NOR2X1_LOC_610/a_36_216# 0.01fF
C68872 INVX1_LOC_18/A NAND2X1_LOC_647/a_36_24# 0.00fF
C68873 INVX1_LOC_49/A NOR2X1_LOC_261/A 0.01fF
C68874 NOR2X1_LOC_720/A INVX1_LOC_57/A 0.02fF
C68875 NOR2X1_LOC_504/Y INVX1_LOC_46/A 0.19fF
C68876 INVX1_LOC_141/Y INVX1_LOC_119/Y 0.02fF
C68877 INVX1_LOC_306/Y INVX1_LOC_4/A 0.03fF
C68878 INVX1_LOC_39/A INVX1_LOC_32/A 0.03fF
C68879 INVX1_LOC_269/A NOR2X1_LOC_89/A 0.07fF
C68880 NOR2X1_LOC_458/Y INVX1_LOC_38/A -0.00fF
C68881 INVX1_LOC_171/A NOR2X1_LOC_9/Y 0.03fF
C68882 INVX1_LOC_147/A INVX1_LOC_28/A 0.32fF
C68883 INVX1_LOC_300/A INVX1_LOC_11/Y 0.01fF
C68884 INVX1_LOC_271/A NOR2X1_LOC_654/A 0.26fF
C68885 NAND2X1_LOC_561/B INVX1_LOC_42/A 0.03fF
C68886 NAND2X1_LOC_139/A INVX1_LOC_280/A 0.03fF
C68887 INVX1_LOC_289/Y NOR2X1_LOC_48/B 0.10fF
C68888 INVX1_LOC_226/Y NAND2X1_LOC_465/A 0.00fF
C68889 NAND2X1_LOC_337/B NAND2X1_LOC_74/B 0.07fF
C68890 INVX1_LOC_30/A NAND2X1_LOC_475/Y 0.62fF
C68891 INVX1_LOC_120/Y VDD -0.00fF
C68892 INVX1_LOC_57/A INVX1_LOC_129/A 0.00fF
C68893 NOR2X1_LOC_220/A NOR2X1_LOC_562/A 0.01fF
C68894 INVX1_LOC_136/A INVX1_LOC_27/Y 0.03fF
C68895 INVX1_LOC_121/Y INVX1_LOC_38/A 0.39fF
C68896 NOR2X1_LOC_790/B NOR2X1_LOC_383/B 0.01fF
C68897 INVX1_LOC_17/A NOR2X1_LOC_114/Y 0.01fF
C68898 INVX1_LOC_135/A NOR2X1_LOC_78/A 0.09fF
C68899 INVX1_LOC_40/A VDD 1.10fF
C68900 INVX1_LOC_96/Y INVX1_LOC_44/A 0.09fF
C68901 INVX1_LOC_269/A NOR2X1_LOC_170/A 0.04fF
C68902 INVX1_LOC_25/A NOR2X1_LOC_15/a_36_216# 0.00fF
C68903 INVX1_LOC_13/Y NAND2X1_LOC_400/a_36_24# 0.01fF
C68904 INVX1_LOC_165/Y VDD 0.41fF
C68905 NOR2X1_LOC_711/a_36_216# INVX1_LOC_117/A 0.02fF
C68906 INVX1_LOC_25/A NAND2X1_LOC_860/A 0.07fF
C68907 NAND2X1_LOC_361/a_36_24# NOR2X1_LOC_489/A 0.00fF
C68908 INVX1_LOC_177/A INVX1_LOC_38/A 0.03fF
C68909 D_INPUT_1 NOR2X1_LOC_598/B 1.29fF
C68910 NOR2X1_LOC_802/A INVX1_LOC_9/A 0.07fF
C68911 NOR2X1_LOC_748/Y NOR2X1_LOC_857/A 0.06fF
C68912 NOR2X1_LOC_123/B NAND2X1_LOC_642/Y 0.09fF
C68913 NOR2X1_LOC_278/a_36_216# INVX1_LOC_304/A 0.01fF
C68914 NAND2X1_LOC_714/B INVX1_LOC_78/A 0.03fF
C68915 INVX1_LOC_230/Y NOR2X1_LOC_672/a_36_216# 0.00fF
C68916 D_INPUT_0 INVX1_LOC_304/A 0.07fF
C68917 NOR2X1_LOC_605/B VDD -0.00fF
C68918 INVX1_LOC_39/Y INVX1_LOC_284/A 0.02fF
C68919 NOR2X1_LOC_667/A NAND2X1_LOC_848/A 0.10fF
C68920 INVX1_LOC_13/A D_INPUT_3 2.97fF
C68921 NAND2X1_LOC_624/B INVX1_LOC_57/A 0.06fF
C68922 INPUT_0 NOR2X1_LOC_368/A 0.01fF
C68923 INVX1_LOC_248/A NAND2X1_LOC_848/A 0.10fF
C68924 INVX1_LOC_222/A NOR2X1_LOC_74/A 0.03fF
C68925 INVX1_LOC_280/Y INVX1_LOC_38/A 0.05fF
C68926 INVX1_LOC_90/A INVX1_LOC_65/A 0.02fF
C68927 NOR2X1_LOC_730/A INVX1_LOC_37/A 0.01fF
C68928 D_INPUT_0 NOR2X1_LOC_670/Y 0.03fF
C68929 INVX1_LOC_41/Y NOR2X1_LOC_662/A 0.02fF
C68930 NOR2X1_LOC_360/Y INVX1_LOC_19/A 0.07fF
C68931 NAND2X1_LOC_14/a_36_24# D_INPUT_3 0.01fF
C68932 NOR2X1_LOC_22/a_36_216# D_INPUT_5 0.00fF
C68933 INVX1_LOC_174/A NAND2X1_LOC_421/a_36_24# 0.01fF
C68934 NOR2X1_LOC_427/Y INVX1_LOC_191/A 0.09fF
C68935 NAND2X1_LOC_303/Y NOR2X1_LOC_25/Y 0.03fF
C68936 INVX1_LOC_239/A NAND2X1_LOC_402/B 0.25fF
C68937 NAND2X1_LOC_808/A INVX1_LOC_37/A 0.07fF
C68938 INVX1_LOC_189/A NAND2X1_LOC_93/B 0.01fF
C68939 INVX1_LOC_102/Y NAND2X1_LOC_642/Y 0.06fF
C68940 NOR2X1_LOC_295/Y INVX1_LOC_285/A 0.02fF
C68941 INVX1_LOC_30/A NOR2X1_LOC_452/a_36_216# 0.01fF
C68942 NOR2X1_LOC_590/A NOR2X1_LOC_38/B 0.03fF
C68943 NOR2X1_LOC_528/Y NOR2X1_LOC_527/Y 0.04fF
C68944 INVX1_LOC_90/A NAND2X1_LOC_267/B 0.02fF
C68945 INVX1_LOC_57/A NOR2X1_LOC_440/B 0.18fF
C68946 INVX1_LOC_8/A INVX1_LOC_84/A 0.15fF
C68947 NOR2X1_LOC_382/Y INVX1_LOC_3/Y 0.03fF
C68948 INVX1_LOC_189/A NAND2X1_LOC_425/Y 0.01fF
C68949 NOR2X1_LOC_295/Y NOR2X1_LOC_814/A 0.02fF
C68950 NAND2X1_LOC_336/a_36_24# INVX1_LOC_78/A 0.01fF
C68951 NOR2X1_LOC_798/A NOR2X1_LOC_717/A 0.03fF
C68952 NAND2X1_LOC_564/B INVX1_LOC_118/A 0.08fF
C68953 NOR2X1_LOC_155/a_36_216# INVX1_LOC_37/A 0.00fF
C68954 NOR2X1_LOC_516/B NOR2X1_LOC_655/Y 0.01fF
C68955 INVX1_LOC_208/A NAND2X1_LOC_93/B 0.07fF
C68956 NAND2X1_LOC_36/A NAND2X1_LOC_3/B 0.28fF
C68957 INVX1_LOC_64/A NOR2X1_LOC_644/a_36_216# 0.02fF
C68958 INVX1_LOC_55/Y INVX1_LOC_14/Y 0.01fF
C68959 NAND2X1_LOC_652/Y INVX1_LOC_76/A 0.03fF
C68960 INVX1_LOC_11/A NOR2X1_LOC_621/A 0.03fF
C68961 INVX1_LOC_33/A INVX1_LOC_133/A 0.02fF
C68962 D_INPUT_4 NAND2X1_LOC_1/Y 0.02fF
C68963 NOR2X1_LOC_45/Y NOR2X1_LOC_449/A 0.03fF
C68964 NAND2X1_LOC_21/Y INVX1_LOC_29/A 0.00fF
C68965 INVX1_LOC_11/A NAND2X1_LOC_64/a_36_24# -0.02fF
C68966 INVX1_LOC_174/A NAND2X1_LOC_425/a_36_24# 0.01fF
C68967 INVX1_LOC_1/A NOR2X1_LOC_15/a_36_216# 0.01fF
C68968 NAND2X1_LOC_860/A INVX1_LOC_1/A 0.05fF
C68969 NOR2X1_LOC_792/B INVX1_LOC_19/A 0.01fF
C68970 NOR2X1_LOC_211/a_36_216# INVX1_LOC_1/A 0.00fF
C68971 NOR2X1_LOC_74/A INVX1_LOC_20/A 0.10fF
C68972 NOR2X1_LOC_82/A NAND2X1_LOC_215/A 0.07fF
C68973 NOR2X1_LOC_147/B NOR2X1_LOC_830/Y 0.04fF
C68974 NAND2X1_LOC_735/B INVX1_LOC_260/A 0.01fF
C68975 NOR2X1_LOC_665/A INVX1_LOC_307/A 0.04fF
C68976 NOR2X1_LOC_323/Y VDD 0.16fF
C68977 NOR2X1_LOC_785/A NOR2X1_LOC_383/B 0.09fF
C68978 NAND2X1_LOC_483/Y INVX1_LOC_284/A 0.01fF
C68979 INVX1_LOC_158/A NAND2X1_LOC_63/Y 0.13fF
C68980 NAND2X1_LOC_549/Y INVX1_LOC_14/A 0.00fF
C68981 NOR2X1_LOC_757/A INVX1_LOC_92/A 0.00fF
C68982 NOR2X1_LOC_439/B NAND2X1_LOC_472/Y 0.01fF
C68983 NAND2X1_LOC_768/a_36_24# NAND2X1_LOC_99/A 0.00fF
C68984 NOR2X1_LOC_75/Y INVX1_LOC_105/Y 0.00fF
C68985 NOR2X1_LOC_6/B INVX1_LOC_106/A 0.27fF
C68986 NOR2X1_LOC_716/B INVX1_LOC_170/Y 0.01fF
C68987 NAND2X1_LOC_858/B NAND2X1_LOC_650/B 0.08fF
C68988 NOR2X1_LOC_9/Y INVX1_LOC_20/A 0.28fF
C68989 INVX1_LOC_83/A NOR2X1_LOC_640/Y 0.08fF
C68990 INVX1_LOC_75/A NAND2X1_LOC_472/Y 0.07fF
C68991 NOR2X1_LOC_516/B NOR2X1_LOC_649/B 0.01fF
C68992 NOR2X1_LOC_779/Y INVX1_LOC_213/A 0.05fF
C68993 NAND2X1_LOC_451/Y INVX1_LOC_19/A 0.12fF
C68994 INVX1_LOC_17/Y INVX1_LOC_31/A 0.08fF
C68995 NOR2X1_LOC_516/B INVX1_LOC_3/A 0.06fF
C68996 NOR2X1_LOC_539/a_36_216# INVX1_LOC_19/A 0.02fF
C68997 INVX1_LOC_200/Y INVX1_LOC_31/A 0.16fF
C68998 INVX1_LOC_120/A NOR2X1_LOC_61/A 0.03fF
C68999 INVX1_LOC_208/Y INVX1_LOC_63/A 0.01fF
C69000 NOR2X1_LOC_91/A INVX1_LOC_250/A 0.06fF
C69001 NAND2X1_LOC_785/A INVX1_LOC_102/A 0.01fF
C69002 NOR2X1_LOC_516/B NOR2X1_LOC_814/a_36_216# 0.00fF
C69003 NAND2X1_LOC_729/Y NOR2X1_LOC_829/A 0.10fF
C69004 INVX1_LOC_25/Y NAND2X1_LOC_773/B 0.08fF
C69005 NOR2X1_LOC_737/a_36_216# INVX1_LOC_139/Y 0.00fF
C69006 NOR2X1_LOC_773/Y NAND2X1_LOC_74/B 0.07fF
C69007 NOR2X1_LOC_577/Y NOR2X1_LOC_334/Y 0.12fF
C69008 INVX1_LOC_89/A NOR2X1_LOC_197/B 0.28fF
C69009 INVX1_LOC_58/A NOR2X1_LOC_382/Y 0.02fF
C69010 NOR2X1_LOC_624/A NOR2X1_LOC_623/B 0.02fF
C69011 NOR2X1_LOC_448/Y NOR2X1_LOC_453/Y 0.00fF
C69012 INVX1_LOC_181/Y INVX1_LOC_181/A 0.01fF
C69013 NAND2X1_LOC_787/A INVX1_LOC_30/A 0.06fF
C69014 INVX1_LOC_132/A NOR2X1_LOC_621/B 0.04fF
C69015 INVX1_LOC_17/A NOR2X1_LOC_61/B 0.07fF
C69016 INVX1_LOC_21/A NAND2X1_LOC_30/Y 0.02fF
C69017 NOR2X1_LOC_499/a_36_216# NOR2X1_LOC_383/B 0.00fF
C69018 INVX1_LOC_53/Y INVX1_LOC_12/A 0.07fF
C69019 NOR2X1_LOC_392/B INVX1_LOC_4/Y 0.46fF
C69020 INVX1_LOC_43/Y INVX1_LOC_306/Y 0.16fF
C69021 INVX1_LOC_14/A NAND2X1_LOC_347/B 0.13fF
C69022 NAND2X1_LOC_363/B INVX1_LOC_30/A 0.01fF
C69023 NOR2X1_LOC_91/A NOR2X1_LOC_495/Y 0.09fF
C69024 INVX1_LOC_245/Y NOR2X1_LOC_626/Y 0.02fF
C69025 NOR2X1_LOC_639/B INVX1_LOC_36/A 0.24fF
C69026 NOR2X1_LOC_75/Y INVX1_LOC_27/A 0.04fF
C69027 INVX1_LOC_136/A NAND2X1_LOC_561/a_36_24# 0.01fF
C69028 INVX1_LOC_41/Y INVX1_LOC_57/A 0.03fF
C69029 NOR2X1_LOC_357/Y NAND2X1_LOC_212/Y 0.01fF
C69030 NOR2X1_LOC_486/Y VDD 0.25fF
C69031 INVX1_LOC_64/A NOR2X1_LOC_657/Y 0.07fF
C69032 INVX1_LOC_278/Y NOR2X1_LOC_48/B 0.25fF
C69033 INVX1_LOC_17/Y NOR2X1_LOC_617/a_36_216# -0.00fF
C69034 INVX1_LOC_278/A NAND2X1_LOC_634/Y 0.10fF
C69035 D_GATE_741 NOR2X1_LOC_463/a_36_216# 0.03fF
C69036 NOR2X1_LOC_348/B NOR2X1_LOC_334/Y 0.02fF
C69037 INVX1_LOC_286/Y NOR2X1_LOC_304/Y 0.02fF
C69038 NOR2X1_LOC_665/A INVX1_LOC_12/A 0.07fF
C69039 INVX1_LOC_31/A NOR2X1_LOC_406/A 0.03fF
C69040 NAND2X1_LOC_714/B NOR2X1_LOC_503/Y 0.07fF
C69041 INVX1_LOC_178/A INVX1_LOC_211/A 0.03fF
C69042 NOR2X1_LOC_617/Y INVX1_LOC_57/A 0.06fF
C69043 NOR2X1_LOC_210/B NAND2X1_LOC_213/a_36_24# 0.00fF
C69044 NOR2X1_LOC_706/A NAND2X1_LOC_425/Y 0.01fF
C69045 NOR2X1_LOC_91/Y NAND2X1_LOC_793/B 1.22fF
C69046 NAND2X1_LOC_593/Y INVX1_LOC_57/A 0.03fF
C69047 NAND2X1_LOC_802/a_36_24# INVX1_LOC_78/A 0.00fF
C69048 INVX1_LOC_13/A NAND2X1_LOC_233/a_36_24# 0.01fF
C69049 NOR2X1_LOC_78/A INVX1_LOC_280/A 0.12fF
C69050 NOR2X1_LOC_188/A NAND2X1_LOC_656/B 0.02fF
C69051 INVX1_LOC_11/A INVX1_LOC_269/A 0.15fF
C69052 INVX1_LOC_77/A INVX1_LOC_29/Y 0.03fF
C69053 INVX1_LOC_24/A NOR2X1_LOC_392/Y 0.00fF
C69054 INVX1_LOC_136/A INVX1_LOC_5/A 0.44fF
C69055 NAND2X1_LOC_538/Y NAND2X1_LOC_799/A 0.08fF
C69056 NAND2X1_LOC_537/Y NAND2X1_LOC_539/a_36_24# 0.01fF
C69057 NOR2X1_LOC_344/A NOR2X1_LOC_383/B 0.02fF
C69058 NOR2X1_LOC_357/Y INVX1_LOC_14/Y 0.10fF
C69059 NOR2X1_LOC_332/A NAND2X1_LOC_207/Y 0.02fF
C69060 NAND2X1_LOC_656/Y NOR2X1_LOC_755/Y 0.03fF
C69061 INVX1_LOC_269/A NAND2X1_LOC_381/Y 0.03fF
C69062 INVX1_LOC_155/Y INVX1_LOC_270/A 0.01fF
C69063 INVX1_LOC_155/A INVX1_LOC_270/Y 0.08fF
C69064 NOR2X1_LOC_756/Y INVX1_LOC_63/A 0.10fF
C69065 INVX1_LOC_304/A NAND2X1_LOC_848/A 0.21fF
C69066 INVX1_LOC_315/Y NOR2X1_LOC_655/Y 0.02fF
C69067 INVX1_LOC_28/A NAND2X1_LOC_768/Y 0.04fF
C69068 NOR2X1_LOC_655/B INVX1_LOC_87/A 0.03fF
C69069 NAND2X1_LOC_361/Y INVX1_LOC_23/A 0.07fF
C69070 NAND2X1_LOC_350/B NAND2X1_LOC_470/B 0.26fF
C69071 NOR2X1_LOC_758/Y INVX1_LOC_57/A 0.00fF
C69072 INVX1_LOC_90/A NAND2X1_LOC_81/B 0.00fF
C69073 NOR2X1_LOC_332/A NOR2X1_LOC_847/B -0.07fF
C69074 INVX1_LOC_95/Y NOR2X1_LOC_119/a_36_216# 0.01fF
C69075 NAND2X1_LOC_794/B NOR2X1_LOC_68/A 0.03fF
C69076 INVX1_LOC_136/A INVX1_LOC_178/A 0.10fF
C69077 NOR2X1_LOC_325/A NOR2X1_LOC_334/Y 0.03fF
C69078 VDD NOR2X1_LOC_816/Y 0.24fF
C69079 INVX1_LOC_263/A INVX1_LOC_271/Y 0.04fF
C69080 NAND2X1_LOC_181/Y NOR2X1_LOC_278/Y 0.01fF
C69081 INVX1_LOC_22/A NOR2X1_LOC_334/Y 0.11fF
C69082 INVX1_LOC_186/A NOR2X1_LOC_862/B 0.78fF
C69083 NOR2X1_LOC_567/B INVX1_LOC_19/A 0.64fF
C69084 INVX1_LOC_256/A NOR2X1_LOC_160/B 1.15fF
C69085 INVX1_LOC_91/A NAND2X1_LOC_798/B 0.07fF
C69086 INVX1_LOC_75/A NAND2X1_LOC_773/B 0.07fF
C69087 D_GATE_366 INVX1_LOC_109/Y 0.02fF
C69088 NOR2X1_LOC_536/A NAND2X1_LOC_211/Y 0.01fF
C69089 D_INPUT_0 INVX1_LOC_19/Y 0.02fF
C69090 INVX1_LOC_299/A NAND2X1_LOC_311/a_36_24# 0.00fF
C69091 INVX1_LOC_16/A NOR2X1_LOC_36/A 0.95fF
C69092 NOR2X1_LOC_279/Y INVX1_LOC_118/A 0.03fF
C69093 INVX1_LOC_278/A INVX1_LOC_8/A 0.02fF
C69094 INVX1_LOC_290/A NAND2X1_LOC_454/Y 0.24fF
C69095 INVX1_LOC_124/A INVX1_LOC_29/Y 0.28fF
C69096 NOR2X1_LOC_188/A NOR2X1_LOC_721/B 0.01fF
C69097 NOR2X1_LOC_300/a_36_216# INVX1_LOC_54/A 0.00fF
C69098 NAND2X1_LOC_559/Y INVX1_LOC_217/A 0.04fF
C69099 INVX1_LOC_2/Y INVX1_LOC_9/A 0.09fF
C69100 INVX1_LOC_63/Y NOR2X1_LOC_665/Y 0.05fF
C69101 NOR2X1_LOC_215/A NOR2X1_LOC_759/Y 0.01fF
C69102 NAND2X1_LOC_140/A INVX1_LOC_15/A 0.03fF
C69103 NAND2X1_LOC_121/a_36_24# INVX1_LOC_72/A 0.01fF
C69104 INVX1_LOC_315/Y NOR2X1_LOC_649/B 0.13fF
C69105 INVX1_LOC_123/A NOR2X1_LOC_673/B 0.01fF
C69106 NOR2X1_LOC_590/A NOR2X1_LOC_389/A 0.09fF
C69107 INVX1_LOC_27/A NOR2X1_LOC_419/Y 0.01fF
C69108 VDD NOR2X1_LOC_351/Y 0.02fF
C69109 NAND2X1_LOC_538/Y INVX1_LOC_18/A 0.07fF
C69110 INVX1_LOC_315/Y INVX1_LOC_3/A 0.03fF
C69111 INVX1_LOC_21/A INVX1_LOC_49/A 0.19fF
C69112 INVX1_LOC_36/A NOR2X1_LOC_218/A 0.03fF
C69113 NAND2X1_LOC_787/A NAND2X1_LOC_722/A 0.01fF
C69114 NAND2X1_LOC_714/B NOR2X1_LOC_152/Y 0.07fF
C69115 NOR2X1_LOC_364/A NAND2X1_LOC_469/B 0.11fF
C69116 NOR2X1_LOC_510/Y INVX1_LOC_33/A 0.07fF
C69117 NOR2X1_LOC_757/Y INVX1_LOC_271/A 0.02fF
C69118 NAND2X1_LOC_729/Y NAND2X1_LOC_537/Y 0.06fF
C69119 NAND2X1_LOC_84/Y NAND2X1_LOC_347/B 0.00fF
C69120 INVX1_LOC_27/A NOR2X1_LOC_716/B 0.10fF
C69121 INVX1_LOC_136/A NOR2X1_LOC_786/a_36_216# 0.02fF
C69122 INVX1_LOC_136/A NAND2X1_LOC_337/B 0.10fF
C69123 NAND2X1_LOC_434/Y NAND2X1_LOC_453/A 0.02fF
C69124 INVX1_LOC_136/A NOR2X1_LOC_816/A 0.03fF
C69125 NAND2X1_LOC_9/Y INVX1_LOC_256/Y 0.12fF
C69126 NOR2X1_LOC_598/B NOR2X1_LOC_620/B 0.03fF
C69127 NOR2X1_LOC_356/A INVX1_LOC_4/A 0.46fF
C69128 INVX1_LOC_90/A INVX1_LOC_4/Y 0.15fF
C69129 NOR2X1_LOC_453/Y INVX1_LOC_49/A 0.01fF
C69130 NOR2X1_LOC_681/Y INVX1_LOC_92/A 0.28fF
C69131 NOR2X1_LOC_91/A NAND2X1_LOC_319/A 0.02fF
C69132 INVX1_LOC_233/A INVX1_LOC_256/Y 1.28fF
C69133 VDD INVX1_LOC_241/Y 0.60fF
C69134 INVX1_LOC_37/A INVX1_LOC_92/A 0.27fF
C69135 NOR2X1_LOC_389/B INVX1_LOC_4/Y 0.03fF
C69136 INVX1_LOC_123/A INVX1_LOC_29/A 0.01fF
C69137 INVX1_LOC_17/Y NAND2X1_LOC_859/Y 0.34fF
C69138 INVX1_LOC_200/Y NAND2X1_LOC_859/Y 0.05fF
C69139 INVX1_LOC_269/A NOR2X1_LOC_474/A 0.00fF
C69140 NOR2X1_LOC_220/B INVX1_LOC_149/A 0.00fF
C69141 NOR2X1_LOC_208/Y NOR2X1_LOC_218/A 0.01fF
C69142 INVX1_LOC_269/A NOR2X1_LOC_593/Y 0.01fF
C69143 INVX1_LOC_249/A NOR2X1_LOC_75/Y 0.00fF
C69144 NOR2X1_LOC_361/B INVX1_LOC_33/A 2.51fF
C69145 NAND2X1_LOC_763/B INVX1_LOC_30/A 0.02fF
C69146 NOR2X1_LOC_590/A INVX1_LOC_62/Y 0.02fF
C69147 INVX1_LOC_24/A NOR2X1_LOC_599/Y 0.03fF
C69148 INVX1_LOC_1/A NOR2X1_LOC_516/Y 0.01fF
C69149 INVX1_LOC_21/A INVX1_LOC_2/A 0.14fF
C69150 NOR2X1_LOC_74/A INVX1_LOC_4/A 0.36fF
C69151 NAND2X1_LOC_348/A INVX1_LOC_4/Y 0.06fF
C69152 INVX1_LOC_120/A NAND2X1_LOC_246/a_36_24# 0.00fF
C69153 NAND2X1_LOC_347/B NOR2X1_LOC_612/B 0.09fF
C69154 NAND2X1_LOC_92/a_36_24# NOR2X1_LOC_271/Y 0.00fF
C69155 INVX1_LOC_21/A NOR2X1_LOC_226/A 0.21fF
C69156 INVX1_LOC_245/Y INVX1_LOC_153/A 0.01fF
C69157 INVX1_LOC_221/A NAND2X1_LOC_537/Y 0.10fF
C69158 NOR2X1_LOC_9/Y INVX1_LOC_4/A 1.28fF
C69159 INVX1_LOC_17/Y NAND2X1_LOC_866/B 0.01fF
C69160 INVX1_LOC_235/Y INVX1_LOC_197/A 0.03fF
C69161 NAND2X1_LOC_169/Y NAND2X1_LOC_170/A 0.19fF
C69162 INVX1_LOC_89/A NOR2X1_LOC_260/Y 0.02fF
C69163 NOR2X1_LOC_332/A NOR2X1_LOC_660/Y 0.04fF
C69164 NOR2X1_LOC_130/A NOR2X1_LOC_392/Y 0.01fF
C69165 INVX1_LOC_292/A NOR2X1_LOC_570/B 0.01fF
C69166 NAND2X1_LOC_361/Y INVX1_LOC_31/A 0.09fF
C69167 INVX1_LOC_230/Y INVX1_LOC_34/A 0.28fF
C69168 NOR2X1_LOC_447/Y INVX1_LOC_36/A 0.01fF
C69169 INVX1_LOC_47/Y INVX1_LOC_91/A 0.03fF
C69170 NOR2X1_LOC_295/Y NOR2X1_LOC_590/A 0.44fF
C69171 NOR2X1_LOC_503/Y NAND2X1_LOC_802/a_36_24# 0.00fF
C69172 INVX1_LOC_208/A NOR2X1_LOC_348/Y 0.10fF
C69173 INVX1_LOC_206/Y INVX1_LOC_271/Y 0.07fF
C69174 NOR2X1_LOC_441/Y NAND2X1_LOC_332/Y 0.22fF
C69175 NOR2X1_LOC_91/Y INVX1_LOC_71/A 0.07fF
C69176 NOR2X1_LOC_590/A NOR2X1_LOC_844/A 0.00fF
C69177 INVX1_LOC_149/A INVX1_LOC_225/Y 0.00fF
C69178 NOR2X1_LOC_68/A NOR2X1_LOC_350/A 0.00fF
C69179 NOR2X1_LOC_685/A NOR2X1_LOC_685/B 0.00fF
C69180 NAND2X1_LOC_842/B NOR2X1_LOC_717/A 0.00fF
C69181 VDD INVX1_LOC_106/Y 0.23fF
C69182 NOR2X1_LOC_655/B NOR2X1_LOC_82/A 0.03fF
C69183 NAND2X1_LOC_787/a_36_24# NOR2X1_LOC_667/A 0.00fF
C69184 INVX1_LOC_64/A NOR2X1_LOC_356/A 0.07fF
C69185 INVX1_LOC_96/A NOR2X1_LOC_464/Y 0.00fF
C69186 NAND2X1_LOC_114/B NOR2X1_LOC_537/Y 0.39fF
C69187 INVX1_LOC_119/A INVX1_LOC_286/Y 0.00fF
C69188 INVX1_LOC_11/A NAND2X1_LOC_563/A 1.49fF
C69189 INVX1_LOC_12/A INVX1_LOC_77/Y 0.07fF
C69190 INVX1_LOC_2/Y NOR2X1_LOC_861/Y 0.10fF
C69191 INVX1_LOC_12/Y NOR2X1_LOC_89/A 0.12fF
C69192 INVX1_LOC_58/A NOR2X1_LOC_527/a_36_216# 0.02fF
C69193 NOR2X1_LOC_446/A NOR2X1_LOC_458/B 0.14fF
C69194 NAND2X1_LOC_381/Y NAND2X1_LOC_563/A 0.03fF
C69195 NOR2X1_LOC_600/Y INVX1_LOC_271/Y 0.01fF
C69196 NOR2X1_LOC_335/A INVX1_LOC_94/A 0.19fF
C69197 INVX1_LOC_256/A INVX1_LOC_208/A 0.28fF
C69198 NAND2X1_LOC_574/a_36_24# INVX1_LOC_135/A 0.01fF
C69199 INVX1_LOC_57/Y NAND2X1_LOC_357/B 0.00fF
C69200 NOR2X1_LOC_536/A NAND2X1_LOC_207/B 0.03fF
C69201 INVX1_LOC_185/A NOR2X1_LOC_662/A 0.02fF
C69202 NOR2X1_LOC_180/B INVX1_LOC_50/Y 0.07fF
C69203 NAND2X1_LOC_53/Y INVX1_LOC_16/A 0.15fF
C69204 NAND2X1_LOC_392/a_36_24# NOR2X1_LOC_130/A 0.01fF
C69205 NAND2X1_LOC_573/Y INVX1_LOC_135/A 0.01fF
C69206 INVX1_LOC_178/A NAND2X1_LOC_862/Y 0.06fF
C69207 INVX1_LOC_65/A INVX1_LOC_18/Y 0.01fF
C69208 D_INPUT_3 INVX1_LOC_32/A 0.10fF
C69209 INVX1_LOC_200/Y INVX1_LOC_6/A 0.02fF
C69210 NOR2X1_LOC_590/A NOR2X1_LOC_220/A 0.02fF
C69211 INVX1_LOC_21/A INPUT_1 0.03fF
C69212 INVX1_LOC_14/Y INVX1_LOC_32/A 0.16fF
C69213 NOR2X1_LOC_647/B NOR2X1_LOC_516/B 0.00fF
C69214 NOR2X1_LOC_67/A NAND2X1_LOC_577/A 0.00fF
C69215 NAND2X1_LOC_807/Y NOR2X1_LOC_406/A 0.27fF
C69216 D_INPUT_1 INVX1_LOC_201/A 0.09fF
C69217 NOR2X1_LOC_142/a_36_216# INVX1_LOC_109/Y 0.00fF
C69218 INVX1_LOC_18/A NOR2X1_LOC_709/A 0.02fF
C69219 INVX1_LOC_64/A NOR2X1_LOC_74/A 0.10fF
C69220 NOR2X1_LOC_68/A NOR2X1_LOC_84/Y 0.28fF
C69221 NOR2X1_LOC_162/Y NOR2X1_LOC_160/a_36_216# 0.00fF
C69222 NOR2X1_LOC_528/Y NOR2X1_LOC_654/A 0.01fF
C69223 NOR2X1_LOC_331/B NAND2X1_LOC_792/B 0.02fF
C69224 NAND2X1_LOC_493/Y NAND2X1_LOC_866/B 0.01fF
C69225 NOR2X1_LOC_470/B INVX1_LOC_89/A 0.03fF
C69226 NAND2X1_LOC_848/A INVX1_LOC_19/Y 0.10fF
C69227 NOR2X1_LOC_226/A NAND2X1_LOC_354/Y 0.05fF
C69228 INVX1_LOC_1/A INVX1_LOC_85/Y 0.10fF
C69229 NOR2X1_LOC_590/A NOR2X1_LOC_548/Y 1.73fF
C69230 NOR2X1_LOC_230/Y NOR2X1_LOC_229/Y 0.15fF
C69231 INVX1_LOC_136/A NOR2X1_LOC_773/Y 0.15fF
C69232 NAND2X1_LOC_778/Y NOR2X1_LOC_322/Y 0.10fF
C69233 INVX1_LOC_33/A INVX1_LOC_153/Y 0.03fF
C69234 NOR2X1_LOC_82/A NOR2X1_LOC_99/B 0.11fF
C69235 INVX1_LOC_77/A INVX1_LOC_60/Y 0.72fF
C69236 NOR2X1_LOC_58/a_36_216# INVX1_LOC_272/A 0.01fF
C69237 INVX1_LOC_249/Y INVX1_LOC_113/Y 0.01fF
C69238 INVX1_LOC_17/A NAND2X1_LOC_189/a_36_24# 0.00fF
C69239 INVX1_LOC_130/A NOR2X1_LOC_561/Y 0.03fF
C69240 INVX1_LOC_124/Y NOR2X1_LOC_589/A 0.15fF
C69241 NOR2X1_LOC_67/A NAND2X1_LOC_656/A 0.12fF
C69242 NOR2X1_LOC_219/a_36_216# INVX1_LOC_96/Y 0.00fF
C69243 NOR2X1_LOC_599/Y NAND2X1_LOC_800/Y 0.02fF
C69244 INVX1_LOC_59/Y NAND2X1_LOC_215/A 0.07fF
C69245 INVX1_LOC_112/A NAND2X1_LOC_215/A 0.02fF
C69246 VDD NOR2X1_LOC_798/Y 0.26fF
C69247 INVX1_LOC_38/A INVX1_LOC_4/Y 0.12fF
C69248 NOR2X1_LOC_361/a_36_216# NAND2X1_LOC_656/Y 0.00fF
C69249 NOR2X1_LOC_15/Y NOR2X1_LOC_322/Y 0.05fF
C69250 INVX1_LOC_290/Y NOR2X1_LOC_600/a_36_216# 0.00fF
C69251 INVX1_LOC_33/A INVX1_LOC_177/A 0.04fF
C69252 NOR2X1_LOC_68/A INVX1_LOC_290/A 0.07fF
C69253 INVX1_LOC_24/A INVX1_LOC_25/Y 0.06fF
C69254 NOR2X1_LOC_188/A NAND2X1_LOC_473/A 0.01fF
C69255 VDD INVX1_LOC_275/Y 0.41fF
C69256 VDD NOR2X1_LOC_748/A 2.15fF
C69257 INVX1_LOC_41/A INVX1_LOC_196/A 0.01fF
C69258 NAND2X1_LOC_656/Y INVX1_LOC_72/A 0.07fF
C69259 INVX1_LOC_24/A NOR2X1_LOC_302/B 0.03fF
C69260 INVX1_LOC_33/A NOR2X1_LOC_547/a_36_216# 0.00fF
C69261 NOR2X1_LOC_372/A NOR2X1_LOC_497/Y 0.04fF
C69262 NAND2X1_LOC_796/B NOR2X1_LOC_45/B 1.75fF
C69263 NOR2X1_LOC_36/B NOR2X1_LOC_11/Y 0.03fF
C69264 NAND2X1_LOC_30/Y NAND2X1_LOC_51/B 0.44fF
C69265 INVX1_LOC_77/A NOR2X1_LOC_160/Y 0.01fF
C69266 NOR2X1_LOC_681/Y INVX1_LOC_53/A 0.46fF
C69267 NOR2X1_LOC_627/Y INVX1_LOC_85/A 0.01fF
C69268 INVX1_LOC_209/Y INVX1_LOC_22/A 0.03fF
C69269 NOR2X1_LOC_543/A INVX1_LOC_71/A 0.01fF
C69270 NOR2X1_LOC_304/Y NOR2X1_LOC_56/Y 0.01fF
C69271 INVX1_LOC_53/A INVX1_LOC_37/A 1.68fF
C69272 INVX1_LOC_227/A NOR2X1_LOC_596/A 0.01fF
C69273 NOR2X1_LOC_557/Y INVX1_LOC_25/Y 0.04fF
C69274 INVX1_LOC_81/A NOR2X1_LOC_561/Y 0.07fF
C69275 NOR2X1_LOC_804/a_36_216# INVX1_LOC_177/A 0.00fF
C69276 INVX1_LOC_293/Y INVX1_LOC_42/A -0.00fF
C69277 NOR2X1_LOC_569/Y NOR2X1_LOC_577/Y 0.04fF
C69278 INVX1_LOC_35/A NOR2X1_LOC_145/Y 0.18fF
C69279 NAND2X1_LOC_341/A INVX1_LOC_34/A 0.06fF
C69280 INVX1_LOC_89/A INVX1_LOC_159/A 0.07fF
C69281 NOR2X1_LOC_802/A INVX1_LOC_179/Y 0.18fF
C69282 NAND2X1_LOC_37/a_36_24# INVX1_LOC_75/A 0.00fF
C69283 INVX1_LOC_230/Y INPUT_0 0.14fF
C69284 NOR2X1_LOC_15/Y NOR2X1_LOC_562/B 1.39fF
C69285 INVX1_LOC_250/A NAND2X1_LOC_807/Y 0.03fF
C69286 NOR2X1_LOC_809/A INVX1_LOC_9/A 0.02fF
C69287 NOR2X1_LOC_504/Y NOR2X1_LOC_505/Y 0.00fF
C69288 INVX1_LOC_2/A NOR2X1_LOC_667/A 0.28fF
C69289 INVX1_LOC_34/A GATE_479 0.05fF
C69290 NAND2X1_LOC_545/a_36_24# INVX1_LOC_28/A 0.01fF
C69291 NOR2X1_LOC_808/A NOR2X1_LOC_78/B 0.03fF
C69292 NOR2X1_LOC_124/B NOR2X1_LOC_719/A 0.36fF
C69293 NOR2X1_LOC_718/B INVX1_LOC_22/A 0.02fF
C69294 INVX1_LOC_2/A INVX1_LOC_248/A 0.98fF
C69295 NOR2X1_LOC_816/A NOR2X1_LOC_165/a_36_216# 0.00fF
C69296 VDD NOR2X1_LOC_304/Y 0.77fF
C69297 INVX1_LOC_36/A INVX1_LOC_302/A 0.01fF
C69298 NOR2X1_LOC_355/A INVX1_LOC_77/A 0.09fF
C69299 NOR2X1_LOC_168/B NAND2X1_LOC_323/B 0.07fF
C69300 NOR2X1_LOC_785/Y INVX1_LOC_33/A 0.03fF
C69301 NOR2X1_LOC_267/A NAND2X1_LOC_842/a_36_24# 0.01fF
C69302 NOR2X1_LOC_226/A NOR2X1_LOC_667/A 0.07fF
C69303 INVX1_LOC_9/A INVX1_LOC_29/Y 0.14fF
C69304 INVX1_LOC_132/A INVX1_LOC_135/A 0.28fF
C69305 NAND2X1_LOC_74/B INVX1_LOC_42/A 0.18fF
C69306 INVX1_LOC_289/Y INVX1_LOC_291/Y 0.03fF
C69307 NOR2X1_LOC_590/A INVX1_LOC_51/Y 0.01fF
C69308 NAND2X1_LOC_800/A NOR2X1_LOC_304/Y 0.02fF
C69309 NOR2X1_LOC_226/A INVX1_LOC_248/A 0.10fF
C69310 NAND2X1_LOC_785/A NAND2X1_LOC_543/Y -0.02fF
C69311 INVX1_LOC_185/A INVX1_LOC_57/A 0.03fF
C69312 INVX1_LOC_17/A NAND2X1_LOC_655/A 0.10fF
C69313 NOR2X1_LOC_847/A NOR2X1_LOC_847/B 0.55fF
C69314 NAND2X1_LOC_866/B NOR2X1_LOC_495/Y 0.01fF
C69315 NOR2X1_LOC_620/B NAND2X1_LOC_528/a_36_24# 0.02fF
C69316 NOR2X1_LOC_242/A INVX1_LOC_37/A 0.05fF
C69317 INVX1_LOC_233/Y INVX1_LOC_38/A 0.04fF
C69318 INVX1_LOC_279/A INVX1_LOC_104/A 0.07fF
C69319 NOR2X1_LOC_831/B NAND2X1_LOC_288/B 0.02fF
C69320 INVX1_LOC_206/A NOR2X1_LOC_501/a_36_216# 0.01fF
C69321 INVX1_LOC_157/Y INVX1_LOC_53/A 0.01fF
C69322 INVX1_LOC_269/A INVX1_LOC_74/A 0.02fF
C69323 NOR2X1_LOC_297/a_36_216# INVX1_LOC_135/A 0.00fF
C69324 D_INPUT_5 INPUT_7 0.06fF
C69325 NAND2X1_LOC_392/A NAND2X1_LOC_181/Y 0.00fF
C69326 NOR2X1_LOC_186/Y NOR2X1_LOC_152/A 0.01fF
C69327 NOR2X1_LOC_264/Y NOR2X1_LOC_749/a_36_216# 0.00fF
C69328 NOR2X1_LOC_288/A INVX1_LOC_135/A 0.04fF
C69329 INVX1_LOC_41/A INVX1_LOC_47/A 0.02fF
C69330 INVX1_LOC_24/A INVX1_LOC_75/A 0.06fF
C69331 NOR2X1_LOC_468/Y NAND2X1_LOC_650/B 0.01fF
C69332 NOR2X1_LOC_384/Y NOR2X1_LOC_86/a_36_216# 0.01fF
C69333 INVX1_LOC_53/A NOR2X1_LOC_743/Y 0.19fF
C69334 NOR2X1_LOC_669/Y VDD 0.38fF
C69335 NOR2X1_LOC_807/B NOR2X1_LOC_324/B 0.06fF
C69336 INVX1_LOC_249/A NOR2X1_LOC_151/Y 0.02fF
C69337 INVX1_LOC_226/Y INVX1_LOC_16/A 0.10fF
C69338 NAND2X1_LOC_565/B INVX1_LOC_25/Y 0.01fF
C69339 NAND2X1_LOC_579/A NAND2X1_LOC_721/A 0.04fF
C69340 NOR2X1_LOC_214/B NOR2X1_LOC_52/B 0.00fF
C69341 NOR2X1_LOC_100/A NOR2X1_LOC_99/B 0.02fF
C69342 NOR2X1_LOC_67/Y NOR2X1_LOC_38/B 0.05fF
C69343 NAND2X1_LOC_564/B NAND2X1_LOC_182/a_36_24# 0.00fF
C69344 NOR2X1_LOC_808/A INVX1_LOC_83/A 0.03fF
C69345 NOR2X1_LOC_155/A NOR2X1_LOC_678/A 0.03fF
C69346 NOR2X1_LOC_710/B VDD -0.00fF
C69347 INVX1_LOC_310/A INVX1_LOC_148/Y 0.01fF
C69348 NOR2X1_LOC_655/B INVX1_LOC_306/A 0.13fF
C69349 INVX1_LOC_78/A NAND2X1_LOC_74/B 0.08fF
C69350 NOR2X1_LOC_328/Y NAND2X1_LOC_712/A 0.02fF
C69351 INVX1_LOC_157/A NAND2X1_LOC_350/B 0.05fF
C69352 NOR2X1_LOC_831/Y NAND2X1_LOC_175/Y 0.00fF
C69353 INVX1_LOC_26/A INVX1_LOC_19/A 0.10fF
C69354 NAND2X1_LOC_149/Y INVX1_LOC_114/A 0.06fF
C69355 INVX1_LOC_49/A NAND2X1_LOC_51/B 0.11fF
C69356 NOR2X1_LOC_510/Y NOR2X1_LOC_351/Y 0.01fF
C69357 NOR2X1_LOC_553/Y NOR2X1_LOC_570/A 0.02fF
C69358 INVX1_LOC_256/A NAND2X1_LOC_211/Y 0.13fF
C69359 NOR2X1_LOC_569/Y INVX1_LOC_22/A 0.07fF
C69360 NAND2X1_LOC_9/Y NAND2X1_LOC_85/Y 0.01fF
C69361 NOR2X1_LOC_541/a_36_216# INVX1_LOC_77/A 0.00fF
C69362 NAND2X1_LOC_579/A NOR2X1_LOC_323/a_36_216# 0.03fF
C69363 INVX1_LOC_27/A NOR2X1_LOC_709/B 0.41fF
C69364 INVX1_LOC_198/Y INVX1_LOC_78/Y 0.05fF
C69365 INVX1_LOC_263/A INVX1_LOC_279/A 0.08fF
C69366 INVX1_LOC_21/A INVX1_LOC_118/A 0.29fF
C69367 NOR2X1_LOC_646/A INVX1_LOC_7/A 0.01fF
C69368 INVX1_LOC_11/A INVX1_LOC_12/Y 0.07fF
C69369 INVX1_LOC_49/A INVX1_LOC_311/A 0.07fF
C69370 INVX1_LOC_77/A NOR2X1_LOC_552/Y 0.09fF
C69371 NOR2X1_LOC_114/Y INVX1_LOC_94/Y 0.00fF
C69372 NOR2X1_LOC_89/A NOR2X1_LOC_89/Y 0.10fF
C69373 INVX1_LOC_218/Y INVX1_LOC_176/A 0.00fF
C69374 INVX1_LOC_10/A INVX1_LOC_16/A 0.11fF
C69375 INPUT_3 D_INPUT_3 0.55fF
C69376 INVX1_LOC_36/A NAND2X1_LOC_271/a_36_24# 0.00fF
C69377 INVX1_LOC_182/Y INVX1_LOC_104/A 0.03fF
C69378 NOR2X1_LOC_532/Y INVX1_LOC_179/Y 0.20fF
C69379 NAND2X1_LOC_323/B INVX1_LOC_132/Y 0.03fF
C69380 INVX1_LOC_64/A NOR2X1_LOC_243/B 0.07fF
C69381 NOR2X1_LOC_233/a_36_216# NAND2X1_LOC_243/Y 0.01fF
C69382 NOR2X1_LOC_130/A INVX1_LOC_25/Y 0.14fF
C69383 NOR2X1_LOC_65/B NAND2X1_LOC_74/B 0.14fF
C69384 NOR2X1_LOC_329/B INVX1_LOC_133/Y 0.01fF
C69385 NAND2X1_LOC_564/A INVX1_LOC_19/A 0.02fF
C69386 NOR2X1_LOC_71/Y INVX1_LOC_56/Y 0.08fF
C69387 INVX1_LOC_33/A INVX1_LOC_285/Y 0.05fF
C69388 NAND2X1_LOC_711/Y VDD 0.17fF
C69389 INVX1_LOC_276/A NOR2X1_LOC_329/B 0.07fF
C69390 NAND2X1_LOC_364/A INVX1_LOC_314/A 0.04fF
C69391 INVX1_LOC_90/A NAND2X1_LOC_862/A 0.00fF
C69392 NOR2X1_LOC_437/Y NOR2X1_LOC_269/Y 0.00fF
C69393 INVX1_LOC_24/A NAND2X1_LOC_620/a_36_24# 0.00fF
C69394 NAND2X1_LOC_714/B NAND2X1_LOC_802/Y 0.00fF
C69395 NOR2X1_LOC_716/B NOR2X1_LOC_528/Y 0.10fF
C69396 INVX1_LOC_286/Y NOR2X1_LOC_425/Y 0.04fF
C69397 D_INPUT_1 INVX1_LOC_29/A 0.63fF
C69398 NOR2X1_LOC_791/B INVX1_LOC_76/A 0.07fF
C69399 INVX1_LOC_103/A INVX1_LOC_54/A 1.76fF
C69400 NAND2X1_LOC_470/B NAND2X1_LOC_53/a_36_24# 0.01fF
C69401 INVX1_LOC_226/Y INVX1_LOC_28/A 0.01fF
C69402 NAND2X1_LOC_531/a_36_24# INVX1_LOC_234/A 0.01fF
C69403 NAND2X1_LOC_223/A INVX1_LOC_4/Y 0.07fF
C69404 INPUT_3 INVX1_LOC_230/A 0.72fF
C69405 INVX1_LOC_306/A NOR2X1_LOC_99/B 0.02fF
C69406 INVX1_LOC_2/A INVX1_LOC_311/A 0.07fF
C69407 INVX1_LOC_263/A INVX1_LOC_182/Y 0.00fF
C69408 NOR2X1_LOC_295/a_36_216# NOR2X1_LOC_318/B 0.00fF
C69409 NAND2X1_LOC_139/A NOR2X1_LOC_45/B 0.14fF
C69410 NAND2X1_LOC_850/Y NOR2X1_LOC_74/A 1.08fF
C69411 INVX1_LOC_33/A INVX1_LOC_65/A 0.03fF
C69412 NOR2X1_LOC_428/Y INVX1_LOC_118/A 0.16fF
C69413 INVX1_LOC_24/A NAND2X1_LOC_453/A 0.03fF
C69414 NAND2X1_LOC_656/Y INVX1_LOC_313/Y 0.01fF
C69415 NOR2X1_LOC_592/A NAND2X1_LOC_798/B 0.01fF
C69416 NOR2X1_LOC_660/Y NOR2X1_LOC_847/A 0.20fF
C69417 NOR2X1_LOC_678/A NOR2X1_LOC_833/B 0.43fF
C69418 NOR2X1_LOC_770/Y INVX1_LOC_83/A 0.04fF
C69419 INVX1_LOC_41/A INVX1_LOC_95/Y 0.07fF
C69420 NOR2X1_LOC_106/A NAND2X1_LOC_105/a_36_24# 0.02fF
C69421 INVX1_LOC_28/A INVX1_LOC_10/A 0.71fF
C69422 INVX1_LOC_184/A INVX1_LOC_37/A 0.02fF
C69423 NOR2X1_LOC_652/Y INVX1_LOC_29/A 0.15fF
C69424 INVX1_LOC_251/Y NOR2X1_LOC_78/A 0.32fF
C69425 INVX1_LOC_208/A INVX1_LOC_69/Y 0.02fF
C69426 INVX1_LOC_21/A NAND2X1_LOC_63/Y 0.03fF
C69427 NOR2X1_LOC_340/Y INVX1_LOC_176/A 0.02fF
C69428 INVX1_LOC_26/A INVX1_LOC_26/Y 0.04fF
C69429 INVX1_LOC_119/A NOR2X1_LOC_56/Y 0.01fF
C69430 NAND2X1_LOC_354/Y INVX1_LOC_118/A 0.02fF
C69431 INVX1_LOC_1/A NAND2X1_LOC_782/B 0.02fF
C69432 NOR2X1_LOC_433/A INVX1_LOC_12/Y 0.10fF
C69433 NOR2X1_LOC_124/B INVX1_LOC_76/A 0.00fF
C69434 INVX1_LOC_142/A INVX1_LOC_274/A 0.01fF
C69435 INVX1_LOC_75/A NOR2X1_LOC_130/A 0.10fF
C69436 NOR2X1_LOC_359/Y NOR2X1_LOC_331/B 0.06fF
C69437 NAND2X1_LOC_862/Y INVX1_LOC_140/A 0.03fF
C69438 NAND2X1_LOC_555/Y NAND2X1_LOC_141/Y 0.14fF
C69439 INVX1_LOC_267/A NAND2X1_LOC_659/B 0.01fF
C69440 NAND2X1_LOC_149/Y INVX1_LOC_12/A 0.11fF
C69441 NOR2X1_LOC_614/Y NOR2X1_LOC_78/A 0.04fF
C69442 NOR2X1_LOC_454/Y NOR2X1_LOC_583/Y 0.06fF
C69443 INVX1_LOC_208/Y NOR2X1_LOC_318/B 0.00fF
C69444 NOR2X1_LOC_226/A INVX1_LOC_304/A 0.02fF
C69445 NAND2X1_LOC_159/a_36_24# INVX1_LOC_48/A 0.00fF
C69446 INVX1_LOC_2/A NOR2X1_LOC_670/Y 0.02fF
C69447 INVX1_LOC_298/Y D_INPUT_1 0.03fF
C69448 NOR2X1_LOC_91/A INVX1_LOC_50/A 0.22fF
C69449 INVX1_LOC_279/A INVX1_LOC_206/Y 0.07fF
C69450 INVX1_LOC_119/A VDD 0.45fF
C69451 INVX1_LOC_89/A NOR2X1_LOC_721/Y 0.33fF
C69452 NAND2X1_LOC_112/Y NOR2X1_LOC_45/B 0.12fF
C69453 NOR2X1_LOC_497/Y NAND2X1_LOC_560/A 0.01fF
C69454 NOR2X1_LOC_107/Y INVX1_LOC_19/A 0.02fF
C69455 INVX1_LOC_34/A INVX1_LOC_44/A 0.02fF
C69456 INVX1_LOC_267/A VDD -0.00fF
C69457 NOR2X1_LOC_52/B INVX1_LOC_12/Y 2.11fF
C69458 NAND2X1_LOC_563/A INVX1_LOC_74/A 0.28fF
C69459 INVX1_LOC_58/A NOR2X1_LOC_638/Y -0.02fF
C69460 NOR2X1_LOC_493/B VDD -0.00fF
C69461 NAND2X1_LOC_569/A NOR2X1_LOC_536/A 0.00fF
C69462 NOR2X1_LOC_401/B VDD 0.02fF
C69463 INVX1_LOC_50/A INVX1_LOC_23/A 0.10fF
C69464 NOR2X1_LOC_297/a_36_216# INVX1_LOC_280/A 0.01fF
C69465 INVX1_LOC_230/Y NOR2X1_LOC_84/B 0.02fF
C69466 NOR2X1_LOC_500/Y NOR2X1_LOC_35/Y 0.10fF
C69467 INVX1_LOC_226/Y NOR2X1_LOC_35/Y 0.10fF
C69468 NOR2X1_LOC_78/B INVX1_LOC_37/A 0.24fF
C69469 INVX1_LOC_279/A NOR2X1_LOC_600/Y 0.01fF
C69470 NOR2X1_LOC_703/B INVX1_LOC_220/A 0.01fF
C69471 NOR2X1_LOC_216/Y INVX1_LOC_75/A 0.21fF
C69472 INVX1_LOC_21/A NAND2X1_LOC_618/Y 0.03fF
C69473 INVX1_LOC_103/A NOR2X1_LOC_48/B 0.17fF
C69474 NOR2X1_LOC_328/Y NOR2X1_LOC_421/Y 0.04fF
C69475 NAND2X1_LOC_550/A NOR2X1_LOC_89/A 0.02fF
C69476 NAND2X1_LOC_462/B INVX1_LOC_255/A 0.01fF
C69477 INVX1_LOC_25/Y NOR2X1_LOC_280/Y 0.11fF
C69478 NOR2X1_LOC_160/B NOR2X1_LOC_89/A 0.12fF
C69479 INVX1_LOC_240/A INVX1_LOC_54/A 0.12fF
C69480 NOR2X1_LOC_716/B NOR2X1_LOC_216/B 0.10fF
C69481 NOR2X1_LOC_383/B INVX1_LOC_213/A 0.05fF
C69482 NAND2X1_LOC_79/Y INVX1_LOC_84/A 0.03fF
C69483 INVX1_LOC_63/Y NOR2X1_LOC_364/A 0.04fF
C69484 NOR2X1_LOC_589/A NOR2X1_LOC_266/B 0.02fF
C69485 INVX1_LOC_182/Y INVX1_LOC_206/Y 0.53fF
C69486 NAND2X1_LOC_358/Y INVX1_LOC_176/A 0.01fF
C69487 NAND2X1_LOC_391/Y INVX1_LOC_23/Y 0.03fF
C69488 NOR2X1_LOC_76/A NOR2X1_LOC_124/A 0.03fF
C69489 NOR2X1_LOC_598/B NOR2X1_LOC_678/A 0.03fF
C69490 NOR2X1_LOC_526/Y INVX1_LOC_38/A 0.03fF
C69491 NAND2X1_LOC_72/Y INVX1_LOC_23/A 0.01fF
C69492 INVX1_LOC_22/A NAND2X1_LOC_472/Y 0.07fF
C69493 NOR2X1_LOC_214/B INVX1_LOC_199/A 0.10fF
C69494 NOR2X1_LOC_82/A NOR2X1_LOC_28/a_36_216# 0.00fF
C69495 INVX1_LOC_7/A INVX1_LOC_2/Y 0.08fF
C69496 INVX1_LOC_304/A INPUT_1 0.05fF
C69497 INVX1_LOC_89/A NAND2X1_LOC_659/B 0.10fF
C69498 NOR2X1_LOC_15/Y NOR2X1_LOC_464/Y 0.15fF
C69499 D_INPUT_0 INVX1_LOC_20/A 1.18fF
C69500 NOR2X1_LOC_134/Y INVX1_LOC_19/Y 0.08fF
C69501 INVX1_LOC_176/A NOR2X1_LOC_99/B 0.07fF
C69502 NAND2X1_LOC_303/Y NAND2X1_LOC_175/Y 0.07fF
C69503 NOR2X1_LOC_210/A INVX1_LOC_117/A 0.01fF
C69504 NOR2X1_LOC_679/Y INVX1_LOC_231/A 0.24fF
C69505 NAND2X1_LOC_740/Y INVX1_LOC_296/Y 0.15fF
C69506 NOR2X1_LOC_667/A INVX1_LOC_118/A 0.69fF
C69507 NOR2X1_LOC_576/B NAND2X1_LOC_836/Y 0.06fF
C69508 INVX1_LOC_229/Y NAND2X1_LOC_839/a_36_24# 0.07fF
C69509 INVX1_LOC_24/A NAND2X1_LOC_478/a_36_24# 0.01fF
C69510 NOR2X1_LOC_554/B NAND2X1_LOC_207/Y 0.01fF
C69511 INVX1_LOC_248/A INVX1_LOC_118/A 0.10fF
C69512 NOR2X1_LOC_524/Y NOR2X1_LOC_114/Y 0.04fF
C69513 INVX1_LOC_152/Y NAND2X1_LOC_358/B 0.21fF
C69514 INVX1_LOC_135/A D_GATE_662 0.02fF
C69515 NOR2X1_LOC_111/A NAND2X1_LOC_796/Y 0.04fF
C69516 VDD INVX1_LOC_150/A 0.35fF
C69517 NOR2X1_LOC_130/A NAND2X1_LOC_453/A 0.04fF
C69518 INVX1_LOC_83/A INVX1_LOC_37/A 0.38fF
C69519 NOR2X1_LOC_68/A NOR2X1_LOC_641/a_36_216# 0.01fF
C69520 NOR2X1_LOC_561/Y NOR2X1_LOC_363/Y 0.01fF
C69521 NAND2X1_LOC_363/Y VDD 0.13fF
C69522 INVX1_LOC_136/A INVX1_LOC_42/A 0.27fF
C69523 NOR2X1_LOC_68/A INVX1_LOC_114/Y 0.08fF
C69524 NOR2X1_LOC_160/B INVX1_LOC_104/Y 0.02fF
C69525 NOR2X1_LOC_554/B NOR2X1_LOC_847/B 0.05fF
C69526 INVX1_LOC_89/A VDD 1.80fF
C69527 NOR2X1_LOC_78/B NOR2X1_LOC_743/Y 0.19fF
C69528 NAND2X1_LOC_347/B NOR2X1_LOC_383/B 0.09fF
C69529 D_INPUT_2 INVX1_LOC_29/A 0.22fF
C69530 NOR2X1_LOC_712/B INVX1_LOC_19/A 0.01fF
C69531 INVX1_LOC_62/Y NOR2X1_LOC_67/Y 0.02fF
C69532 NOR2X1_LOC_690/A NAND2X1_LOC_489/Y 1.14fF
C69533 INVX1_LOC_22/A NAND2X1_LOC_637/Y 0.04fF
C69534 INVX1_LOC_5/A NOR2X1_LOC_665/Y 0.02fF
C69535 NOR2X1_LOC_152/Y NAND2X1_LOC_74/B 0.07fF
C69536 INVX1_LOC_101/A INVX1_LOC_9/A 0.02fF
C69537 NAND2X1_LOC_341/a_36_24# INVX1_LOC_117/Y 0.00fF
C69538 INVX1_LOC_6/A INVX1_LOC_159/Y 0.02fF
C69539 NAND2X1_LOC_508/A VDD 0.06fF
C69540 NOR2X1_LOC_406/A NOR2X1_LOC_109/Y 0.05fF
C69541 NOR2X1_LOC_197/Y INVX1_LOC_76/A 0.01fF
C69542 NOR2X1_LOC_736/a_36_216# NOR2X1_LOC_357/Y 0.00fF
C69543 INVX1_LOC_24/A INVX1_LOC_283/A 0.02fF
C69544 NOR2X1_LOC_718/B INVX1_LOC_186/Y 0.47fF
C69545 NOR2X1_LOC_68/A NOR2X1_LOC_467/A 0.42fF
C69546 NOR2X1_LOC_318/B NOR2X1_LOC_501/B 0.00fF
C69547 NAND2X1_LOC_807/A NAND2X1_LOC_286/B 0.01fF
C69548 NOR2X1_LOC_355/A INVX1_LOC_9/A 0.94fF
C69549 NOR2X1_LOC_340/Y NOR2X1_LOC_340/A 0.12fF
C69550 NAND2X1_LOC_352/B NAND2X1_LOC_288/B 0.19fF
C69551 NOR2X1_LOC_561/Y NOR2X1_LOC_358/a_36_216# 0.00fF
C69552 NOR2X1_LOC_665/A INVX1_LOC_92/A 0.00fF
C69553 INVX1_LOC_18/A NOR2X1_LOC_334/Y 0.07fF
C69554 NOR2X1_LOC_91/A INVX1_LOC_61/Y 0.38fF
C69555 INVX1_LOC_136/A INVX1_LOC_78/A 0.04fF
C69556 NOR2X1_LOC_346/B NAND2X1_LOC_206/Y 0.01fF
C69557 INVX1_LOC_149/A INVX1_LOC_19/A 0.01fF
C69558 INVX1_LOC_316/Y NOR2X1_LOC_649/B 0.00fF
C69559 NOR2X1_LOC_6/B NOR2X1_LOC_14/a_36_216# 0.01fF
C69560 INVX1_LOC_27/A NOR2X1_LOC_343/B 0.04fF
C69561 INVX1_LOC_50/A INVX1_LOC_31/A 0.39fF
C69562 INVX1_LOC_7/A NOR2X1_LOC_608/Y 0.02fF
C69563 NOR2X1_LOC_529/Y INVX1_LOC_29/A 0.00fF
C69564 INVX1_LOC_31/A NOR2X1_LOC_105/Y 0.19fF
C69565 NOR2X1_LOC_721/A NAND2X1_LOC_74/B 0.06fF
C69566 INVX1_LOC_45/A NOR2X1_LOC_840/Y 0.01fF
C69567 INVX1_LOC_55/A NOR2X1_LOC_598/B 0.01fF
C69568 NOR2X1_LOC_703/Y VDD 0.24fF
C69569 INVX1_LOC_17/A NOR2X1_LOC_772/B 0.16fF
C69570 NOR2X1_LOC_65/B INVX1_LOC_136/A 0.10fF
C69571 NAND2X1_LOC_717/Y INVX1_LOC_12/A 0.03fF
C69572 INVX1_LOC_35/A NAND2X1_LOC_47/a_36_24# 0.02fF
C69573 INVX1_LOC_75/A NOR2X1_LOC_148/Y 0.03fF
C69574 INVX1_LOC_189/A NOR2X1_LOC_89/A 0.00fF
C69575 NAND2X1_LOC_337/B NOR2X1_LOC_109/a_36_216# 0.00fF
C69576 NOR2X1_LOC_620/B INVX1_LOC_29/A 0.03fF
C69577 INVX1_LOC_142/Y NOR2X1_LOC_727/B 0.24fF
C69578 NOR2X1_LOC_45/B NAND2X1_LOC_464/A 0.02fF
C69579 INVX1_LOC_17/A INVX1_LOC_13/Y 0.03fF
C69580 INVX1_LOC_59/A NOR2X1_LOC_92/Y 0.38fF
C69581 INVX1_LOC_33/A INVX1_LOC_4/Y 0.07fF
C69582 INVX1_LOC_198/Y NOR2X1_LOC_727/B 0.05fF
C69583 NOR2X1_LOC_653/B INVX1_LOC_11/A 0.01fF
C69584 INVX1_LOC_195/A NOR2X1_LOC_476/B 0.01fF
C69585 INVX1_LOC_41/A INVX1_LOC_271/Y 0.10fF
C69586 INVX1_LOC_208/A NOR2X1_LOC_89/A 0.85fF
C69587 NOR2X1_LOC_666/A NOR2X1_LOC_122/A 0.06fF
C69588 INVX1_LOC_25/A NOR2X1_LOC_68/A 0.11fF
C69589 INVX1_LOC_16/A INVX1_LOC_12/A 0.46fF
C69590 NAND2X1_LOC_326/A NAND2X1_LOC_537/Y 0.01fF
C69591 NOR2X1_LOC_396/Y INVX1_LOC_46/A 0.07fF
C69592 INVX1_LOC_72/A NOR2X1_LOC_717/A 0.10fF
C69593 INVX1_LOC_33/Y INVX1_LOC_91/A 0.03fF
C69594 NOR2X1_LOC_598/B INVX1_LOC_305/A 0.11fF
C69595 NOR2X1_LOC_615/Y NOR2X1_LOC_496/Y 0.05fF
C69596 NOR2X1_LOC_321/Y NOR2X1_LOC_250/A 0.02fF
C69597 INVX1_LOC_277/Y INVX1_LOC_213/A 0.04fF
C69598 NOR2X1_LOC_554/B NOR2X1_LOC_660/Y 0.07fF
C69599 D_INPUT_1 INVX1_LOC_228/A 0.33fF
C69600 NAND2X1_LOC_198/B INVX1_LOC_53/A 0.01fF
C69601 INVX1_LOC_75/A NOR2X1_LOC_197/B 0.10fF
C69602 VDD NOR2X1_LOC_24/Y 0.32fF
C69603 NOR2X1_LOC_266/B INVX1_LOC_20/A 0.01fF
C69604 INVX1_LOC_197/Y INVX1_LOC_3/Y 0.00fF
C69605 INVX1_LOC_10/A INVX1_LOC_109/A 0.01fF
C69606 INVX1_LOC_25/A NOR2X1_LOC_204/a_36_216# 0.00fF
C69607 INVX1_LOC_17/A INVX1_LOC_88/A 0.05fF
C69608 NAND2X1_LOC_567/a_36_24# INVX1_LOC_49/Y 0.00fF
C69609 INVX1_LOC_200/Y NOR2X1_LOC_237/Y 0.01fF
C69610 NOR2X1_LOC_448/Y INVX1_LOC_174/A 0.01fF
C69611 INVX1_LOC_12/Y INVX1_LOC_74/A 0.00fF
C69612 NOR2X1_LOC_111/a_36_216# INVX1_LOC_78/A 0.00fF
C69613 NOR2X1_LOC_682/Y INVX1_LOC_20/A 0.03fF
C69614 NOR2X1_LOC_595/Y INVX1_LOC_38/A 0.04fF
C69615 NOR2X1_LOC_303/Y INVX1_LOC_58/Y 0.10fF
C69616 INVX1_LOC_86/A NAND2X1_LOC_425/Y 0.01fF
C69617 INVX1_LOC_37/A INVX1_LOC_46/A 0.03fF
C69618 NOR2X1_LOC_78/B NAND2X1_LOC_72/B 0.00fF
C69619 NAND2X1_LOC_357/B NAND2X1_LOC_288/B 0.01fF
C69620 INVX1_LOC_259/Y INVX1_LOC_113/Y 0.02fF
C69621 INVX1_LOC_40/A INVX1_LOC_4/Y 0.25fF
C69622 INVX1_LOC_256/A NOR2X1_LOC_217/a_36_216# 0.00fF
C69623 NAND2X1_LOC_350/A INVX1_LOC_103/A 0.02fF
C69624 VDD NOR2X1_LOC_425/Y 0.24fF
C69625 INVX1_LOC_272/Y INVX1_LOC_246/A 0.04fF
C69626 INVX1_LOC_115/Y INVX1_LOC_38/A 0.01fF
C69627 INVX1_LOC_304/A INVX1_LOC_118/A 0.07fF
C69628 NAND2X1_LOC_848/A INVX1_LOC_20/A 0.04fF
C69629 D_INPUT_1 INVX1_LOC_8/A 0.20fF
C69630 NAND2X1_LOC_30/Y INVX1_LOC_174/A 0.04fF
C69631 INVX1_LOC_11/A NOR2X1_LOC_160/B 0.69fF
C69632 INVX1_LOC_45/A NAND2X1_LOC_780/Y 0.01fF
C69633 NAND2X1_LOC_363/B NAND2X1_LOC_524/a_36_24# 0.00fF
C69634 NOR2X1_LOC_858/B INVX1_LOC_117/A 0.01fF
C69635 NOR2X1_LOC_311/Y NOR2X1_LOC_743/Y 0.13fF
C69636 INVX1_LOC_21/A INVX1_LOC_61/A 0.04fF
C69637 NOR2X1_LOC_78/B NOR2X1_LOC_863/B 0.13fF
C69638 NAND2X1_LOC_862/Y INVX1_LOC_42/A 0.01fF
C69639 NOR2X1_LOC_71/Y NAND2X1_LOC_74/a_36_24# 0.01fF
C69640 NOR2X1_LOC_804/B INVX1_LOC_292/Y 0.02fF
C69641 NOR2X1_LOC_503/Y INVX1_LOC_211/A 0.06fF
C69642 NOR2X1_LOC_78/A NOR2X1_LOC_862/B 0.11fF
C69643 INVX1_LOC_28/A INVX1_LOC_12/A 8.31fF
C69644 INVX1_LOC_129/Y INVX1_LOC_117/A 0.00fF
C69645 INVX1_LOC_177/A NOR2X1_LOC_748/A 0.05fF
C69646 INVX1_LOC_299/A NOR2X1_LOC_354/B 0.01fF
C69647 NOR2X1_LOC_333/A INVX1_LOC_15/A 0.04fF
C69648 NOR2X1_LOC_368/A INVX1_LOC_19/A 0.24fF
C69649 D_INPUT_0 INVX1_LOC_4/A 0.03fF
C69650 NOR2X1_LOC_91/A NOR2X1_LOC_701/a_36_216# 0.00fF
C69651 NOR2X1_LOC_68/A INVX1_LOC_1/A 0.26fF
C69652 INVX1_LOC_100/A NAND2X1_LOC_773/B 0.03fF
C69653 NOR2X1_LOC_272/Y INVX1_LOC_77/A 0.10fF
C69654 NOR2X1_LOC_15/Y NOR2X1_LOC_457/B 1.00fF
C69655 NOR2X1_LOC_241/a_36_216# INVX1_LOC_49/A 0.02fF
C69656 NOR2X1_LOC_137/Y INVX1_LOC_54/A 0.03fF
C69657 INVX1_LOC_91/A INVX1_LOC_220/A 0.05fF
C69658 INVX1_LOC_22/A NOR2X1_LOC_639/Y 0.04fF
C69659 NOR2X1_LOC_68/A NAND2X1_LOC_131/a_36_24# 0.00fF
C69660 NOR2X1_LOC_163/A NOR2X1_LOC_467/A 0.04fF
C69661 INVX1_LOC_33/Y NAND2X1_LOC_783/a_36_24# 0.00fF
C69662 NAND2X1_LOC_778/Y NAND2X1_LOC_833/Y 0.01fF
C69663 NOR2X1_LOC_35/Y INVX1_LOC_307/A 0.10fF
C69664 INVX1_LOC_286/Y NOR2X1_LOC_599/Y 0.06fF
C69665 INVX1_LOC_54/Y INVX1_LOC_58/Y 1.03fF
C69666 NAND2X1_LOC_860/A NAND2X1_LOC_360/B 0.01fF
C69667 NOR2X1_LOC_112/B NAND2X1_LOC_291/B 0.05fF
C69668 NOR2X1_LOC_822/a_36_216# INVX1_LOC_54/A 0.02fF
C69669 INVX1_LOC_20/A INVX1_LOC_46/Y 0.09fF
C69670 NOR2X1_LOC_242/A INVX1_LOC_310/Y 0.01fF
C69671 INVX1_LOC_46/A NOR2X1_LOC_743/Y 0.56fF
C69672 NOR2X1_LOC_264/a_36_216# INVX1_LOC_314/Y 0.01fF
C69673 NOR2X1_LOC_35/Y NOR2X1_LOC_445/B 0.10fF
C69674 INVX1_LOC_56/Y NAND2X1_LOC_205/A 0.03fF
C69675 INVX1_LOC_269/A INVX1_LOC_314/Y 0.03fF
C69676 NOR2X1_LOC_790/A INVX1_LOC_33/A 0.01fF
C69677 INVX1_LOC_35/A NOR2X1_LOC_67/A 0.07fF
C69678 INVX1_LOC_45/A INVX1_LOC_141/Y 0.01fF
C69679 INVX1_LOC_224/Y NOR2X1_LOC_789/A 0.00fF
C69680 NOR2X1_LOC_289/Y INVX1_LOC_15/A 0.07fF
C69681 INVX1_LOC_119/A NOR2X1_LOC_510/Y 0.03fF
C69682 NOR2X1_LOC_33/a_36_216# NAND2X1_LOC_574/A -0.00fF
C69683 NOR2X1_LOC_389/A INVX1_LOC_177/Y 0.01fF
C69684 INVX1_LOC_294/Y NOR2X1_LOC_440/B 0.01fF
C69685 INPUT_5 INVX1_LOC_173/A 0.34fF
C69686 NOR2X1_LOC_15/Y NAND2X1_LOC_833/Y 0.02fF
C69687 INVX1_LOC_45/A INVX1_LOC_312/Y 0.08fF
C69688 INVX1_LOC_53/Y INVX1_LOC_53/A 0.23fF
C69689 INVX1_LOC_41/A NAND2X1_LOC_773/Y 0.03fF
C69690 INVX1_LOC_17/A INVX1_LOC_303/A 0.07fF
C69691 INVX1_LOC_77/Y INVX1_LOC_92/A 0.07fF
C69692 INVX1_LOC_83/A NOR2X1_LOC_802/a_36_216# 0.00fF
C69693 NOR2X1_LOC_658/Y INVX1_LOC_72/A 0.07fF
C69694 NOR2X1_LOC_205/Y INVX1_LOC_33/A 0.03fF
C69695 NOR2X1_LOC_561/Y INVX1_LOC_29/Y 0.01fF
C69696 INVX1_LOC_2/A NOR2X1_LOC_626/Y 0.09fF
C69697 NOR2X1_LOC_87/B NAND2X1_LOC_473/A 0.10fF
C69698 NAND2X1_LOC_182/A NOR2X1_LOC_468/Y 0.02fF
C69699 INVX1_LOC_103/A NOR2X1_LOC_142/Y 0.29fF
C69700 NOR2X1_LOC_394/a_36_216# NOR2X1_LOC_38/B 0.00fF
C69701 NAND2X1_LOC_218/B NAND2X1_LOC_37/a_36_24# 0.00fF
C69702 NOR2X1_LOC_769/A NAND2X1_LOC_764/a_36_24# 0.02fF
C69703 INVX1_LOC_31/A NAND2X1_LOC_845/a_36_24# 0.00fF
C69704 NOR2X1_LOC_160/B NOR2X1_LOC_433/A 0.07fF
C69705 INVX1_LOC_174/A INVX1_LOC_49/A 1.43fF
C69706 INVX1_LOC_50/A INVX1_LOC_313/A 0.01fF
C69707 INVX1_LOC_100/A NOR2X1_LOC_393/Y 0.06fF
C69708 INVX1_LOC_64/A NAND2X1_LOC_660/Y 0.06fF
C69709 NAND2X1_LOC_803/B INVX1_LOC_63/Y 0.02fF
C69710 NOR2X1_LOC_750/Y INVX1_LOC_135/A 0.06fF
C69711 INVX1_LOC_204/Y NAND2X1_LOC_479/Y 0.09fF
C69712 NAND2X1_LOC_776/a_36_24# INVX1_LOC_41/Y 0.00fF
C69713 INVX1_LOC_201/Y INVX1_LOC_252/Y 0.02fF
C69714 NOR2X1_LOC_20/Y NOR2X1_LOC_399/A 0.12fF
C69715 NOR2X1_LOC_61/Y INVX1_LOC_152/A 0.03fF
C69716 NOR2X1_LOC_536/A NAND2X1_LOC_286/a_36_24# 0.00fF
C69717 INVX1_LOC_2/A NOR2X1_LOC_202/a_36_216# 0.00fF
C69718 INVX1_LOC_292/A NOR2X1_LOC_142/Y 0.03fF
C69719 NOR2X1_LOC_564/Y NOR2X1_LOC_383/B 0.93fF
C69720 INVX1_LOC_50/A NAND2X1_LOC_807/Y 0.03fF
C69721 NOR2X1_LOC_336/B INVX1_LOC_77/A 0.01fF
C69722 NOR2X1_LOC_441/Y INVX1_LOC_67/A 0.02fF
C69723 NAND2X1_LOC_214/B NOR2X1_LOC_391/A 0.07fF
C69724 INVX1_LOC_64/A D_INPUT_0 0.50fF
C69725 NAND2X1_LOC_550/A NOR2X1_LOC_52/B 0.07fF
C69726 NOR2X1_LOC_401/B NOR2X1_LOC_361/B 0.03fF
C69727 NOR2X1_LOC_678/a_36_216# INVX1_LOC_208/A 0.01fF
C69728 INVX1_LOC_269/A NOR2X1_LOC_778/B -0.01fF
C69729 INVX1_LOC_45/A INVX1_LOC_275/A 0.20fF
C69730 INVX1_LOC_136/A NOR2X1_LOC_152/Y 0.10fF
C69731 INVX1_LOC_99/Y NOR2X1_LOC_717/B 0.01fF
C69732 NOR2X1_LOC_614/Y NOR2X1_LOC_790/a_36_216# 0.00fF
C69733 NOR2X1_LOC_160/B NOR2X1_LOC_52/B 0.15fF
C69734 INVX1_LOC_311/A NOR2X1_LOC_631/Y 0.05fF
C69735 NOR2X1_LOC_782/a_36_216# INVX1_LOC_72/A 0.00fF
C69736 INVX1_LOC_11/A INVX1_LOC_189/A 0.03fF
C69737 INVX1_LOC_313/Y NOR2X1_LOC_717/A 0.08fF
C69738 NOR2X1_LOC_402/a_36_216# NOR2X1_LOC_361/B 0.12fF
C69739 NOR2X1_LOC_536/A NOR2X1_LOC_662/A 0.03fF
C69740 NOR2X1_LOC_89/A NAND2X1_LOC_211/Y 0.03fF
C69741 NOR2X1_LOC_389/A INVX1_LOC_104/A 0.19fF
C69742 NAND2X1_LOC_652/Y INVX1_LOC_23/A 0.01fF
C69743 NAND2X1_LOC_364/A INVX1_LOC_77/A 0.21fF
C69744 NAND2X1_LOC_724/Y NAND2X1_LOC_863/A 0.02fF
C69745 NOR2X1_LOC_793/Y INVX1_LOC_305/Y 0.18fF
C69746 NAND2X1_LOC_794/B INVX1_LOC_10/A 0.01fF
C69747 NOR2X1_LOC_445/Y INVX1_LOC_223/A 0.28fF
C69748 INVX1_LOC_27/A NOR2X1_LOC_391/A 0.02fF
C69749 NOR2X1_LOC_754/A INVX1_LOC_20/A -0.00fF
C69750 INVX1_LOC_263/A NAND2X1_LOC_190/Y 0.14fF
C69751 NAND2X1_LOC_563/Y NAND2X1_LOC_577/A 0.20fF
C69752 NOR2X1_LOC_590/A NOR2X1_LOC_175/A 0.05fF
C69753 NOR2X1_LOC_82/A INVX1_LOC_43/A 0.01fF
C69754 NAND2X1_LOC_222/B NOR2X1_LOC_516/B 0.00fF
C69755 NAND2X1_LOC_655/A INVX1_LOC_94/Y 0.02fF
C69756 NOR2X1_LOC_655/B INVX1_LOC_292/A 0.08fF
C69757 INVX1_LOC_224/A NOR2X1_LOC_516/B 0.39fF
C69758 INVX1_LOC_24/A NOR2X1_LOC_577/Y 0.11fF
C69759 NOR2X1_LOC_691/B NOR2X1_LOC_729/A 0.05fF
C69760 NOR2X1_LOC_74/A INVX1_LOC_129/A -0.02fF
C69761 INVX1_LOC_13/A INVX1_LOC_14/A 0.12fF
C69762 NAND2X1_LOC_717/Y NAND2X1_LOC_733/Y 0.03fF
C69763 INVX1_LOC_11/A NOR2X1_LOC_516/B 0.06fF
C69764 NOR2X1_LOC_717/B NAND2X1_LOC_513/B 0.01fF
C69765 NOR2X1_LOC_212/a_36_216# NOR2X1_LOC_389/B 0.00fF
C69766 INVX1_LOC_36/Y INVX1_LOC_15/A 0.10fF
C69767 INVX1_LOC_50/A INVX1_LOC_6/A 0.13fF
C69768 INVX1_LOC_24/Y INVX1_LOC_279/A 0.01fF
C69769 NOR2X1_LOC_434/Y NOR2X1_LOC_174/A 0.05fF
C69770 NOR2X1_LOC_718/B INVX1_LOC_18/A 0.01fF
C69771 INVX1_LOC_91/A INVX1_LOC_23/Y 0.91fF
C69772 INVX1_LOC_45/A NOR2X1_LOC_168/B 0.06fF
C69773 INVX1_LOC_135/A INVX1_LOC_239/A 0.09fF
C69774 NAND2X1_LOC_381/Y NOR2X1_LOC_516/B 0.01fF
C69775 NOR2X1_LOC_9/Y INVX1_LOC_129/A 0.03fF
C69776 NOR2X1_LOC_632/Y NAND2X1_LOC_719/a_36_24# 0.00fF
C69777 NAND2X1_LOC_53/Y INVX1_LOC_290/A 0.05fF
C69778 INVX1_LOC_229/A INVX1_LOC_229/Y 0.12fF
C69779 NOR2X1_LOC_321/Y NOR2X1_LOC_106/A 0.02fF
C69780 NOR2X1_LOC_168/B NOR2X1_LOC_568/A 0.03fF
C69781 NOR2X1_LOC_266/B INVX1_LOC_4/A 0.04fF
C69782 INVX1_LOC_174/A NOR2X1_LOC_161/Y 0.01fF
C69783 INVX1_LOC_124/Y NAND2X1_LOC_850/Y 0.10fF
C69784 INVX1_LOC_124/A NAND2X1_LOC_364/A 0.27fF
C69785 NAND2X1_LOC_149/Y NOR2X1_LOC_155/a_36_216# 0.01fF
C69786 NOR2X1_LOC_403/B INVX1_LOC_8/A 0.08fF
C69787 D_INPUT_2 INVX1_LOC_8/A 0.13fF
C69788 NOR2X1_LOC_570/a_36_216# INVX1_LOC_177/A 0.00fF
C69789 NOR2X1_LOC_61/Y INVX1_LOC_29/A 0.07fF
C69790 NOR2X1_LOC_263/a_36_216# INVX1_LOC_181/Y 0.00fF
C69791 NOR2X1_LOC_15/Y NOR2X1_LOC_76/A 0.03fF
C69792 INVX1_LOC_24/A NOR2X1_LOC_348/B 0.05fF
C69793 NOR2X1_LOC_596/A INVX1_LOC_104/A 0.02fF
C69794 NOR2X1_LOC_246/A INVX1_LOC_14/A 0.07fF
C69795 INVX1_LOC_34/A NOR2X1_LOC_219/a_36_216# 0.01fF
C69796 NAND2X1_LOC_733/Y INVX1_LOC_16/A 0.03fF
C69797 INVX1_LOC_291/A NAND2X1_LOC_74/B 0.07fF
C69798 NOR2X1_LOC_266/a_36_216# NOR2X1_LOC_773/Y -0.01fF
C69799 INVX1_LOC_1/A NOR2X1_LOC_163/A 0.04fF
C69800 INVX1_LOC_35/A NAND2X1_LOC_103/a_36_24# 0.00fF
C69801 INVX1_LOC_239/A INVX1_LOC_169/Y 0.03fF
C69802 INVX1_LOC_246/A INVX1_LOC_10/A 0.00fF
C69803 NOR2X1_LOC_781/Y NAND2X1_LOC_661/B 0.10fF
C69804 INVX1_LOC_38/A D_INPUT_5 0.03fF
C69805 NOR2X1_LOC_78/B NAND2X1_LOC_198/B 0.10fF
C69806 NOR2X1_LOC_662/A NOR2X1_LOC_649/B 0.08fF
C69807 NOR2X1_LOC_592/a_36_216# NOR2X1_LOC_130/A 0.00fF
C69808 NAND2X1_LOC_67/Y NOR2X1_LOC_736/Y 0.02fF
C69809 INVX1_LOC_19/Y INVX1_LOC_118/A 0.05fF
C69810 INVX1_LOC_136/A NAND2X1_LOC_859/B 0.17fF
C69811 NAND2X1_LOC_741/B NAND2X1_LOC_712/A 0.05fF
C69812 NAND2X1_LOC_513/B NOR2X1_LOC_151/Y 0.07fF
C69813 NOR2X1_LOC_152/Y NOR2X1_LOC_111/a_36_216# 0.00fF
C69814 INVX1_LOC_24/A NOR2X1_LOC_346/B 0.03fF
C69815 NOR2X1_LOC_662/A NOR2X1_LOC_661/A 0.18fF
C69816 INVX1_LOC_23/Y NOR2X1_LOC_290/a_36_216# 0.00fF
C69817 INVX1_LOC_217/A INVX1_LOC_16/A 0.51fF
C69818 INVX1_LOC_269/A NAND2X1_LOC_123/Y 0.02fF
C69819 INVX1_LOC_54/Y NOR2X1_LOC_537/A 0.48fF
C69820 NOR2X1_LOC_74/A NOR2X1_LOC_440/B 0.14fF
C69821 NOR2X1_LOC_15/Y INVX1_LOC_73/A 0.03fF
C69822 INVX1_LOC_88/A NOR2X1_LOC_171/Y 0.01fF
C69823 NOR2X1_LOC_88/Y INVX1_LOC_102/A 0.07fF
C69824 INVX1_LOC_200/A INVX1_LOC_28/A 0.14fF
C69825 INVX1_LOC_2/A INVX1_LOC_153/A 0.04fF
C69826 NAND2X1_LOC_11/Y INVX1_LOC_77/A 0.06fF
C69827 NAND2X1_LOC_717/Y NAND2X1_LOC_787/B 0.05fF
C69828 NOR2X1_LOC_51/A D_INPUT_5 0.08fF
C69829 INVX1_LOC_45/A NAND2X1_LOC_656/Y 0.04fF
C69830 INVX1_LOC_40/Y NOR2X1_LOC_332/A 0.01fF
C69831 INVX1_LOC_24/A INVX1_LOC_22/A 0.15fF
C69832 NOR2X1_LOC_815/a_36_216# INVX1_LOC_214/Y 0.00fF
C69833 NOR2X1_LOC_9/Y NOR2X1_LOC_440/B 0.02fF
C69834 NOR2X1_LOC_795/Y NOR2X1_LOC_288/A 0.46fF
C69835 NOR2X1_LOC_392/Y NAND2X1_LOC_659/B 0.02fF
C69836 NAND2X1_LOC_364/Y NAND2X1_LOC_323/B 0.03fF
C69837 NOR2X1_LOC_186/Y NOR2X1_LOC_45/B 0.07fF
C69838 INVX1_LOC_208/A NOR2X1_LOC_433/A 0.50fF
C69839 INVX1_LOC_11/A NOR2X1_LOC_706/A 0.09fF
C69840 NAND2X1_LOC_198/B NAND2X1_LOC_392/Y 0.03fF
C69841 INVX1_LOC_45/A INVX1_LOC_132/Y 0.03fF
C69842 INVX1_LOC_102/A INVX1_LOC_84/A 0.07fF
C69843 INVX1_LOC_108/Y INVX1_LOC_36/Y 0.12fF
C69844 INVX1_LOC_277/A INVX1_LOC_85/Y 0.00fF
C69845 NAND2X1_LOC_803/B INVX1_LOC_302/Y 0.06fF
C69846 NAND2X1_LOC_35/B NAND2X1_LOC_33/Y 0.21fF
C69847 INVX1_LOC_46/Y INVX1_LOC_4/A 0.06fF
C69848 NAND2X1_LOC_733/Y INVX1_LOC_28/A 0.03fF
C69849 NOR2X1_LOC_89/A NOR2X1_LOC_605/A 0.04fF
C69850 INVX1_LOC_55/Y NOR2X1_LOC_717/Y 0.15fF
C69851 INVX1_LOC_135/A NOR2X1_LOC_91/Y 0.01fF
C69852 INVX1_LOC_136/A NOR2X1_LOC_150/a_36_216# 0.00fF
C69853 INVX1_LOC_16/A NAND2X1_LOC_787/B 0.02fF
C69854 NAND2X1_LOC_99/a_36_24# INVX1_LOC_232/A 0.06fF
C69855 NAND2X1_LOC_9/Y INVX1_LOC_37/A 0.01fF
C69856 VDD NOR2X1_LOC_392/Y 3.88fF
C69857 NOR2X1_LOC_493/B INVX1_LOC_177/A 0.01fF
C69858 NAND2X1_LOC_190/Y INVX1_LOC_206/Y 0.03fF
C69859 NAND2X1_LOC_573/Y NOR2X1_LOC_45/B 0.07fF
C69860 NOR2X1_LOC_589/A INVX1_LOC_49/A 0.10fF
C69861 INVX1_LOC_233/A INVX1_LOC_37/A 0.07fF
C69862 NOR2X1_LOC_557/Y INVX1_LOC_22/A 0.63fF
C69863 NOR2X1_LOC_220/A INVX1_LOC_104/A 0.17fF
C69864 NOR2X1_LOC_32/B NAND2X1_LOC_721/A 0.02fF
C69865 NOR2X1_LOC_536/A INVX1_LOC_57/A 7.02fF
C69866 NAND2X1_LOC_656/Y INVX1_LOC_71/A 0.65fF
C69867 NOR2X1_LOC_500/A NOR2X1_LOC_717/B 0.11fF
C69868 NOR2X1_LOC_171/a_36_216# NAND2X1_LOC_593/Y 0.00fF
C69869 INVX1_LOC_232/Y NOR2X1_LOC_515/a_36_216# 0.00fF
C69870 INVX1_LOC_36/A NAND2X1_LOC_654/B 0.00fF
C69871 INVX1_LOC_90/A NOR2X1_LOC_360/Y 0.03fF
C69872 NOR2X1_LOC_717/B NOR2X1_LOC_303/Y 0.03fF
C69873 NOR2X1_LOC_189/A INVX1_LOC_10/A 0.03fF
C69874 INVX1_LOC_64/A NOR2X1_LOC_682/Y 0.02fF
C69875 INVX1_LOC_185/Y INVX1_LOC_25/Y 0.09fF
C69876 NAND2X1_LOC_222/B INVX1_LOC_315/Y 0.02fF
C69877 INVX1_LOC_5/A NOR2X1_LOC_562/A 0.03fF
C69878 INVX1_LOC_12/A INVX1_LOC_109/A 0.02fF
C69879 INVX1_LOC_208/A NOR2X1_LOC_52/B 0.00fF
C69880 NAND2X1_LOC_839/Y NAND2X1_LOC_852/Y 0.11fF
C69881 NAND2X1_LOC_363/B NAND2X1_LOC_613/a_36_24# 0.01fF
C69882 NAND2X1_LOC_783/A NOR2X1_LOC_577/Y 0.10fF
C69883 NOR2X1_LOC_389/B NOR2X1_LOC_360/Y 0.10fF
C69884 INVX1_LOC_217/A INVX1_LOC_28/A 1.05fF
C69885 INVX1_LOC_64/A NOR2X1_LOC_859/Y 0.03fF
C69886 INVX1_LOC_231/Y INVX1_LOC_10/A 0.14fF
C69887 INVX1_LOC_255/Y NOR2X1_LOC_514/Y 0.04fF
C69888 NOR2X1_LOC_15/Y NAND2X1_LOC_729/B 0.02fF
C69889 INVX1_LOC_41/A INVX1_LOC_279/A 0.07fF
C69890 NOR2X1_LOC_811/B NOR2X1_LOC_78/B 0.00fF
C69891 NOR2X1_LOC_577/Y NAND2X1_LOC_800/Y 0.02fF
C69892 NOR2X1_LOC_750/Y INVX1_LOC_280/A 0.05fF
C69893 INVX1_LOC_226/Y NOR2X1_LOC_84/Y 0.33fF
C69894 INVX1_LOC_304/Y INVX1_LOC_16/A 0.08fF
C69895 NOR2X1_LOC_577/Y NOR2X1_LOC_130/A 0.07fF
C69896 NOR2X1_LOC_34/A NOR2X1_LOC_35/Y 0.13fF
C69897 NAND2X1_LOC_190/Y NOR2X1_LOC_600/Y 0.14fF
C69898 INVX1_LOC_104/A NOR2X1_LOC_548/Y 0.01fF
C69899 INVX1_LOC_223/Y VDD 0.21fF
C69900 NOR2X1_LOC_798/A INVX1_LOC_37/A 0.03fF
C69901 INVX1_LOC_64/A NAND2X1_LOC_848/A 0.00fF
C69902 NOR2X1_LOC_770/A INVX1_LOC_90/A 0.02fF
C69903 INVX1_LOC_21/A INVX1_LOC_14/Y 0.03fF
C69904 INVX1_LOC_235/A VDD -0.00fF
C69905 NOR2X1_LOC_717/B NOR2X1_LOC_254/Y 0.29fF
C69906 INVX1_LOC_103/A INVX1_LOC_291/Y 0.03fF
C69907 INVX1_LOC_223/A NOR2X1_LOC_335/B 0.01fF
C69908 INVX1_LOC_142/A NOR2X1_LOC_74/A 0.03fF
C69909 NOR2X1_LOC_226/A NOR2X1_LOC_418/Y 0.02fF
C69910 INVX1_LOC_57/A NAND2X1_LOC_93/B 2.65fF
C69911 INVX1_LOC_143/A INVX1_LOC_22/A 0.02fF
C69912 INVX1_LOC_120/A NOR2X1_LOC_340/Y 0.25fF
C69913 NOR2X1_LOC_78/B INVX1_LOC_53/Y 0.03fF
C69914 NAND2X1_LOC_348/A NOR2X1_LOC_360/Y 0.00fF
C69915 NOR2X1_LOC_67/A NOR2X1_LOC_121/A 0.24fF
C69916 INVX1_LOC_50/Y INVX1_LOC_117/A 0.10fF
C69917 INVX1_LOC_2/A NOR2X1_LOC_589/A 0.07fF
C69918 NOR2X1_LOC_45/Y NOR2X1_LOC_45/B 0.33fF
C69919 INVX1_LOC_89/A INVX1_LOC_153/Y 0.04fF
C69920 NAND2X1_LOC_703/Y INVX1_LOC_37/A 0.07fF
C69921 INVX1_LOC_138/Y INVX1_LOC_9/A 0.03fF
C69922 INVX1_LOC_50/A NAND2X1_LOC_810/B 0.05fF
C69923 INVX1_LOC_45/A INVX1_LOC_78/Y 0.03fF
C69924 NOR2X1_LOC_191/B INVX1_LOC_75/A 0.08fF
C69925 NAND2X1_LOC_471/Y INVX1_LOC_19/A 0.02fF
C69926 NOR2X1_LOC_68/A NOR2X1_LOC_188/A 0.17fF
C69927 NAND2X1_LOC_65/a_36_24# NOR2X1_LOC_243/B 0.00fF
C69928 NOR2X1_LOC_644/A NOR2X1_LOC_344/A 0.02fF
C69929 NAND2X1_LOC_721/a_36_24# NAND2X1_LOC_808/A 0.00fF
C69930 INVX1_LOC_233/A NOR2X1_LOC_177/Y 0.09fF
C69931 INVX1_LOC_267/Y NOR2X1_LOC_459/A 0.01fF
C69932 INVX1_LOC_102/A INVX1_LOC_15/A 0.07fF
C69933 NOR2X1_LOC_151/Y NOR2X1_LOC_303/Y 0.03fF
C69934 INVX1_LOC_89/A INVX1_LOC_121/Y 0.01fF
C69935 NOR2X1_LOC_448/B VDD -0.00fF
C69936 NOR2X1_LOC_89/a_36_216# NAND2X1_LOC_74/B 0.01fF
C69937 INVX1_LOC_41/Y NOR2X1_LOC_74/A 0.05fF
C69938 INVX1_LOC_203/A INVX1_LOC_23/Y 2.46fF
C69939 NOR2X1_LOC_160/B INVX1_LOC_199/A 2.46fF
C69940 INVX1_LOC_90/A NOR2X1_LOC_792/B 0.02fF
C69941 NOR2X1_LOC_843/B NAND2X1_LOC_206/Y 0.07fF
C69942 NOR2X1_LOC_216/Y NOR2X1_LOC_577/Y 0.07fF
C69943 INVX1_LOC_21/A INVX1_LOC_230/A 0.03fF
C69944 INVX1_LOC_106/Y INVX1_LOC_4/Y 0.03fF
C69945 INVX1_LOC_24/A INVX1_LOC_100/A 0.25fF
C69946 INVX1_LOC_57/A NOR2X1_LOC_649/B 0.02fF
C69947 INVX1_LOC_89/A INVX1_LOC_177/A 0.03fF
C69948 NAND2X1_LOC_357/A VDD 0.08fF
C69949 INVX1_LOC_2/A INVX1_LOC_171/A 0.01fF
C69950 NOR2X1_LOC_703/B INVX1_LOC_186/A 0.03fF
C69951 NOR2X1_LOC_272/Y INVX1_LOC_9/A 0.01fF
C69952 INVX1_LOC_233/Y INVX1_LOC_241/Y 0.02fF
C69953 NAND2X1_LOC_860/A NAND2X1_LOC_572/B 0.00fF
C69954 D_INPUT_0 NAND2X1_LOC_850/Y 0.07fF
C69955 NOR2X1_LOC_52/Y NOR2X1_LOC_78/A 0.41fF
C69956 NAND2X1_LOC_740/B NAND2X1_LOC_811/Y 0.02fF
C69957 INVX1_LOC_57/A NOR2X1_LOC_661/A 0.04fF
C69958 NOR2X1_LOC_134/Y INVX1_LOC_20/A 0.03fF
C69959 INVX1_LOC_304/Y INVX1_LOC_28/A 0.07fF
C69960 NOR2X1_LOC_226/A INVX1_LOC_171/A 0.03fF
C69961 NOR2X1_LOC_151/Y NOR2X1_LOC_254/Y 0.07fF
C69962 NOR2X1_LOC_521/Y NAND2X1_LOC_735/B 0.01fF
C69963 INVX1_LOC_5/A NOR2X1_LOC_364/A 0.06fF
C69964 INVX1_LOC_105/A INVX1_LOC_6/A 0.08fF
C69965 INVX1_LOC_71/A INVX1_LOC_78/Y 0.06fF
C69966 INVX1_LOC_55/Y INVX1_LOC_111/Y 0.00fF
C69967 NOR2X1_LOC_655/Y INVX1_LOC_252/A 0.01fF
C69968 NAND2X1_LOC_778/a_36_24# INVX1_LOC_118/A 0.00fF
C69969 INVX1_LOC_290/A INVX1_LOC_10/A 0.12fF
C69970 NOR2X1_LOC_599/Y VDD 0.17fF
C69971 INVX1_LOC_255/Y NOR2X1_LOC_128/B 0.00fF
C69972 NAND2X1_LOC_634/a_36_24# INVX1_LOC_118/A 0.00fF
C69973 INVX1_LOC_237/A NOR2X1_LOC_629/Y 0.00fF
C69974 INVX1_LOC_286/Y NAND2X1_LOC_453/A 0.03fF
C69975 NOR2X1_LOC_717/Y NOR2X1_LOC_357/Y 0.46fF
C69976 INVX1_LOC_64/A INVX1_LOC_5/Y 0.09fF
C69977 NOR2X1_LOC_242/A NAND2X1_LOC_238/a_36_24# 0.00fF
C69978 NAND2X1_LOC_552/A INVX1_LOC_285/A 0.01fF
C69979 NAND2X1_LOC_149/Y INVX1_LOC_92/A 0.34fF
C69980 INVX1_LOC_217/A NOR2X1_LOC_253/Y 0.05fF
C69981 NOR2X1_LOC_243/B NOR2X1_LOC_849/A 0.19fF
C69982 NOR2X1_LOC_781/B INVX1_LOC_83/A 0.10fF
C69983 NOR2X1_LOC_355/A NOR2X1_LOC_561/Y 0.10fF
C69984 INVX1_LOC_77/A NOR2X1_LOC_405/A 2.68fF
C69985 INVX1_LOC_5/A NOR2X1_LOC_814/A 0.11fF
C69986 NOR2X1_LOC_644/A NOR2X1_LOC_540/a_36_216# 0.00fF
C69987 NOR2X1_LOC_45/B NAND2X1_LOC_640/Y 0.12fF
C69988 NOR2X1_LOC_589/A INPUT_1 0.01fF
C69989 NOR2X1_LOC_86/Y VDD 0.24fF
C69990 NOR2X1_LOC_677/Y NOR2X1_LOC_48/B 0.04fF
C69991 NOR2X1_LOC_785/Y INVX1_LOC_89/A 0.01fF
C69992 NOR2X1_LOC_414/Y INVX1_LOC_42/A 0.18fF
C69993 INVX1_LOC_89/A NAND2X1_LOC_378/a_36_24# 0.00fF
C69994 NAND2X1_LOC_198/B INVX1_LOC_46/A 0.14fF
C69995 INVX1_LOC_3/A INVX1_LOC_252/A 0.01fF
C69996 NOR2X1_LOC_703/Y INVX1_LOC_177/A 0.07fF
C69997 INVX1_LOC_120/A NOR2X1_LOC_99/B 0.01fF
C69998 INVX1_LOC_225/A NOR2X1_LOC_45/B 0.03fF
C69999 INVX1_LOC_49/A INVX1_LOC_147/Y 0.01fF
C70000 INVX1_LOC_279/A NOR2X1_LOC_122/Y 0.02fF
C70001 INVX1_LOC_18/A NAND2X1_LOC_472/Y 0.07fF
C70002 INVX1_LOC_278/A INVX1_LOC_102/A -0.00fF
C70003 NOR2X1_LOC_753/a_36_216# INVX1_LOC_76/A 0.00fF
C70004 NAND2X1_LOC_475/a_36_24# NAND2X1_LOC_475/Y 0.02fF
C70005 NAND2X1_LOC_861/Y NAND2X1_LOC_862/Y 0.17fF
C70006 NOR2X1_LOC_722/Y INVX1_LOC_281/Y 0.02fF
C70007 NOR2X1_LOC_181/A NOR2X1_LOC_254/Y 0.00fF
C70008 INVX1_LOC_77/A NOR2X1_LOC_857/A 0.07fF
C70009 NOR2X1_LOC_433/A NAND2X1_LOC_211/Y 0.10fF
C70010 INVX1_LOC_28/A NAND2X1_LOC_808/A 0.19fF
C70011 INVX1_LOC_124/A NOR2X1_LOC_113/A 0.35fF
C70012 NOR2X1_LOC_401/Y INVX1_LOC_98/A 0.02fF
C70013 NOR2X1_LOC_835/B NOR2X1_LOC_835/A 0.04fF
C70014 INVX1_LOC_124/A NOR2X1_LOC_405/A 0.04fF
C70015 NAND2X1_LOC_219/B NAND2X1_LOC_473/A 0.01fF
C70016 NOR2X1_LOC_570/Y NOR2X1_LOC_188/A 0.04fF
C70017 INVX1_LOC_21/A NOR2X1_LOC_831/Y 0.43fF
C70018 INVX1_LOC_314/Y INVX1_LOC_12/Y 0.11fF
C70019 INVX1_LOC_138/Y NOR2X1_LOC_861/Y 0.04fF
C70020 NAND2X1_LOC_794/B INVX1_LOC_12/A 0.07fF
C70021 NAND2X1_LOC_364/A INVX1_LOC_9/A 0.09fF
C70022 NOR2X1_LOC_559/B INVX1_LOC_117/A 0.02fF
C70023 NOR2X1_LOC_372/a_36_216# NAND2X1_LOC_243/Y 0.00fF
C70024 NAND2X1_LOC_794/B NOR2X1_LOC_519/Y 0.03fF
C70025 INVX1_LOC_251/Y NAND2X1_LOC_642/Y 0.01fF
C70026 INVX1_LOC_252/Y NAND2X1_LOC_574/A 0.03fF
C70027 INVX1_LOC_18/A NAND2X1_LOC_637/Y 0.38fF
C70028 NAND2X1_LOC_736/Y VDD 0.70fF
C70029 INVX1_LOC_13/A INVX1_LOC_48/A 0.00fF
C70030 INVX1_LOC_176/Y VDD -0.00fF
C70031 INVX1_LOC_136/A INVX1_LOC_291/A 0.10fF
C70032 NOR2X1_LOC_220/A NOR2X1_LOC_600/Y 0.10fF
C70033 INVX1_LOC_11/A NOR2X1_LOC_605/A 0.02fF
C70034 INVX1_LOC_2/A INVX1_LOC_147/Y 0.36fF
C70035 INVX1_LOC_48/Y INVX1_LOC_12/A 0.08fF
C70036 NAND2X1_LOC_33/Y VDD -0.00fF
C70037 NOR2X1_LOC_52/B NAND2X1_LOC_211/Y 0.12fF
C70038 NAND2X1_LOC_767/a_36_24# INVX1_LOC_84/A 0.00fF
C70039 NOR2X1_LOC_770/A INVX1_LOC_38/A 0.01fF
C70040 INVX1_LOC_136/A NAND2X1_LOC_802/Y 0.12fF
C70041 NAND2X1_LOC_181/Y NOR2X1_LOC_124/A 0.01fF
C70042 NAND2X1_LOC_734/B VDD 0.01fF
C70043 INVX1_LOC_2/A INVX1_LOC_20/A 1.21fF
C70044 NOR2X1_LOC_590/A INVX1_LOC_27/Y 0.01fF
C70045 INVX1_LOC_182/Y NOR2X1_LOC_122/Y 0.00fF
C70046 INVX1_LOC_285/Y INVX1_LOC_150/A 0.10fF
C70047 NAND2X1_LOC_577/a_36_24# NAND2X1_LOC_659/B 0.00fF
C70048 INVX1_LOC_280/Y NOR2X1_LOC_24/Y 0.03fF
C70049 INVX1_LOC_17/A INVX1_LOC_272/A 0.09fF
C70050 NOR2X1_LOC_326/Y NOR2X1_LOC_354/Y 0.01fF
C70051 NAND2X1_LOC_523/a_36_24# INVX1_LOC_309/A 0.00fF
C70052 NOR2X1_LOC_473/B INPUT_0 0.39fF
C70053 INVX1_LOC_50/A INVX1_LOC_270/A 0.00fF
C70054 INVX1_LOC_282/Y VDD 0.68fF
C70055 NOR2X1_LOC_226/A INVX1_LOC_20/A 1.94fF
C70056 INVX1_LOC_224/A NAND2X1_LOC_207/B 0.02fF
C70057 INVX1_LOC_167/Y NAND2X1_LOC_462/B 0.06fF
C70058 NOR2X1_LOC_6/B INVX1_LOC_117/A 0.11fF
C70059 INVX1_LOC_298/Y NOR2X1_LOC_678/A 0.03fF
C70060 INVX1_LOC_16/A NOR2X1_LOC_56/a_36_216# 0.02fF
C70061 INVX1_LOC_178/Y INVX1_LOC_216/A 0.04fF
C70062 NOR2X1_LOC_859/A NOR2X1_LOC_243/B 0.04fF
C70063 INVX1_LOC_230/Y INVX1_LOC_19/A 0.07fF
C70064 NAND2X1_LOC_735/B INVX1_LOC_255/A 0.05fF
C70065 NAND2X1_LOC_850/Y NOR2X1_LOC_266/B 0.11fF
C70066 NOR2X1_LOC_516/B INVX1_LOC_74/A 0.02fF
C70067 INVX1_LOC_223/A INVX1_LOC_84/A 0.42fF
C70068 INVX1_LOC_88/Y NOR2X1_LOC_331/B 0.01fF
C70069 INVX1_LOC_246/A INVX1_LOC_12/A 0.37fF
C70070 NOR2X1_LOC_798/A NAND2X1_LOC_72/B 0.00fF
C70071 NOR2X1_LOC_160/B NOR2X1_LOC_509/a_36_216# 0.00fF
C70072 INVX1_LOC_132/A NOR2X1_LOC_862/B 0.23fF
C70073 INVX1_LOC_14/A INVX1_LOC_32/A 0.29fF
C70074 VDD INVX1_LOC_25/Y 1.88fF
C70075 NAND2X1_LOC_550/A NAND2X1_LOC_254/Y 0.04fF
C70076 NOR2X1_LOC_322/Y INPUT_0 0.10fF
C70077 INVX1_LOC_53/Y INVX1_LOC_46/A 0.10fF
C70078 NAND2X1_LOC_652/Y INVX1_LOC_6/A 0.00fF
C70079 NOR2X1_LOC_791/Y NOR2X1_LOC_278/Y 0.03fF
C70080 NOR2X1_LOC_321/Y NOR2X1_LOC_334/Y 0.01fF
C70081 NAND2X1_LOC_349/B VDD 0.08fF
C70082 NOR2X1_LOC_626/Y NOR2X1_LOC_631/Y 0.29fF
C70083 NOR2X1_LOC_589/A NOR2X1_LOC_586/Y 0.01fF
C70084 INVX1_LOC_50/A NOR2X1_LOC_109/Y 2.93fF
C70085 INVX1_LOC_89/A INVX1_LOC_65/A 0.00fF
C70086 NAND2X1_LOC_451/Y INVX1_LOC_38/A 0.09fF
C70087 NOR2X1_LOC_522/Y NAND2X1_LOC_489/Y 0.30fF
C70088 NAND2X1_LOC_848/A NAND2X1_LOC_850/Y 0.10fF
C70089 NOR2X1_LOC_368/A NAND2X1_LOC_270/a_36_24# 0.00fF
C70090 INVX1_LOC_89/A INVX1_LOC_316/A 0.03fF
C70091 INVX1_LOC_174/A INVX1_LOC_257/A 0.06fF
C70092 INVX1_LOC_92/Y INPUT_0 0.02fF
C70093 INVX1_LOC_22/A NAND2X1_LOC_811/B 0.05fF
C70094 INVX1_LOC_83/A NOR2X1_LOC_585/Y 0.05fF
C70095 INVX1_LOC_24/A INVX1_LOC_186/Y 0.10fF
C70096 INVX1_LOC_88/A INVX1_LOC_94/Y 0.10fF
C70097 INVX1_LOC_75/A NOR2X1_LOC_337/Y 0.03fF
C70098 INVX1_LOC_305/A INVX1_LOC_29/A 0.15fF
C70099 INVX1_LOC_30/Y INVX1_LOC_117/A 0.04fF
C70100 NOR2X1_LOC_419/Y NOR2X1_LOC_721/B 0.12fF
C70101 INVX1_LOC_35/A INVX1_LOC_68/A 0.02fF
C70102 NAND2X1_LOC_648/A INVX1_LOC_20/A 0.02fF
C70103 INPUT_1 INVX1_LOC_20/A 0.05fF
C70104 NAND2X1_LOC_361/Y INVX1_LOC_63/A 0.08fF
C70105 INVX1_LOC_25/A NAND2X1_LOC_474/Y 0.01fF
C70106 INVX1_LOC_190/Y NAND2X1_LOC_453/A 0.12fF
C70107 NOR2X1_LOC_736/Y INVX1_LOC_76/A 0.09fF
C70108 NAND2X1_LOC_303/Y INVX1_LOC_173/A 0.09fF
C70109 INVX1_LOC_85/A INVX1_LOC_84/A 0.12fF
C70110 NAND2X1_LOC_338/B NAND2X1_LOC_94/a_36_24# 0.00fF
C70111 NOR2X1_LOC_175/B NOR2X1_LOC_197/B 0.39fF
C70112 NAND2X1_LOC_537/Y NOR2X1_LOC_654/A 0.10fF
C70113 NOR2X1_LOC_335/A INVX1_LOC_29/A 0.03fF
C70114 NAND2X1_LOC_338/B NAND2X1_LOC_85/Y 0.00fF
C70115 NAND2X1_LOC_149/Y INVX1_LOC_53/A 0.07fF
C70116 INVX1_LOC_16/A INVX1_LOC_92/A 0.07fF
C70117 INVX1_LOC_231/Y INVX1_LOC_12/A 0.03fF
C70118 INVX1_LOC_146/A INVX1_LOC_37/A 0.01fF
C70119 NOR2X1_LOC_439/B VDD -0.00fF
C70120 NOR2X1_LOC_447/Y NAND2X1_LOC_636/a_36_24# 0.00fF
C70121 INVX1_LOC_234/A NOR2X1_LOC_629/Y -0.02fF
C70122 NOR2X1_LOC_685/A INVX1_LOC_91/A 0.03fF
C70123 NOR2X1_LOC_156/A INVX1_LOC_117/A 0.03fF
C70124 INVX1_LOC_22/A NOR2X1_LOC_197/B 0.03fF
C70125 NAND2X1_LOC_543/Y NOR2X1_LOC_88/Y 0.06fF
C70126 NOR2X1_LOC_773/Y INVX1_LOC_285/A 2.25fF
C70127 INVX1_LOC_256/A INVX1_LOC_57/A 0.03fF
C70128 NAND2X1_LOC_394/a_36_24# INVX1_LOC_235/Y 0.00fF
C70129 INVX1_LOC_75/A VDD 4.95fF
C70130 NOR2X1_LOC_636/A NOR2X1_LOC_48/B 0.01fF
C70131 NAND2X1_LOC_569/A NOR2X1_LOC_89/A -0.00fF
C70132 INVX1_LOC_283/Y INVX1_LOC_283/A -0.01fF
C70133 NOR2X1_LOC_361/B NOR2X1_LOC_392/Y 0.00fF
C70134 INVX1_LOC_34/Y NAND2X1_LOC_773/B 0.36fF
C70135 NOR2X1_LOC_360/Y NAND2X1_LOC_223/A 0.03fF
C70136 NOR2X1_LOC_113/B INVX1_LOC_46/A 0.09fF
C70137 NOR2X1_LOC_32/B NOR2X1_LOC_82/A 0.14fF
C70138 NOR2X1_LOC_607/A NOR2X1_LOC_334/Y 0.00fF
C70139 INVX1_LOC_311/A INVX1_LOC_14/Y 0.10fF
C70140 NAND2X1_LOC_543/Y INVX1_LOC_84/A 0.01fF
C70141 NOR2X1_LOC_84/Y INVX1_LOC_12/A 0.46fF
C70142 INVX1_LOC_45/A NOR2X1_LOC_727/B 0.03fF
C70143 NAND2X1_LOC_447/Y INVX1_LOC_91/A 1.32fF
C70144 INVX1_LOC_49/A INVX1_LOC_4/A 0.39fF
C70145 INVX1_LOC_33/A D_INPUT_5 0.00fF
C70146 NAND2X1_LOC_214/B INVX1_LOC_269/A 0.10fF
C70147 NOR2X1_LOC_151/a_36_216# INVX1_LOC_10/Y 0.00fF
C70148 INVX1_LOC_50/A INVX1_LOC_36/A 11.59fF
C70149 NOR2X1_LOC_237/a_36_216# INVX1_LOC_78/A 0.00fF
C70150 NOR2X1_LOC_657/B NOR2X1_LOC_275/A 0.06fF
C70151 INVX1_LOC_36/A NOR2X1_LOC_105/Y 0.01fF
C70152 INVX1_LOC_1/A NAND2X1_LOC_474/Y 0.12fF
C70153 NOR2X1_LOC_6/B INVX1_LOC_3/Y 0.04fF
C70154 NOR2X1_LOC_181/a_36_216# NOR2X1_LOC_678/A 0.00fF
C70155 INVX1_LOC_269/A INVX1_LOC_27/A 0.10fF
C70156 NOR2X1_LOC_389/B NOR2X1_LOC_79/Y 0.01fF
C70157 INVX1_LOC_28/A INVX1_LOC_92/A 4.11fF
C70158 NAND2X1_LOC_349/B INVX1_LOC_133/A 0.26fF
C70159 D_INPUT_7 INVX1_LOC_23/A 0.00fF
C70160 NOR2X1_LOC_778/B NOR2X1_LOC_842/a_36_216# 0.00fF
C70161 NOR2X1_LOC_427/Y INVX1_LOC_38/A 0.01fF
C70162 INVX1_LOC_45/A NOR2X1_LOC_717/A 0.03fF
C70163 NOR2X1_LOC_92/Y NOR2X1_LOC_468/Y 0.08fF
C70164 NOR2X1_LOC_332/A NOR2X1_LOC_814/A 0.08fF
C70165 NOR2X1_LOC_646/A NOR2X1_LOC_664/a_36_216# 0.01fF
C70166 NOR2X1_LOC_709/A INVX1_LOC_47/Y 0.19fF
C70167 NOR2X1_LOC_590/A INVX1_LOC_5/A 0.17fF
C70168 INVX1_LOC_36/A NOR2X1_LOC_224/Y 0.01fF
C70169 NAND2X1_LOC_784/A NOR2X1_LOC_68/A 0.02fF
C70170 INVX1_LOC_186/A NOR2X1_LOC_698/Y 0.07fF
C70171 NOR2X1_LOC_74/A INVX1_LOC_185/A 0.01fF
C70172 NOR2X1_LOC_56/Y NAND2X1_LOC_453/A 0.02fF
C70173 INVX1_LOC_50/A NOR2X1_LOC_208/Y 0.32fF
C70174 INVX1_LOC_290/A INVX1_LOC_12/A 0.12fF
C70175 NOR2X1_LOC_615/Y INVX1_LOC_178/A 0.05fF
C70176 INVX1_LOC_78/Y NOR2X1_LOC_331/B 0.04fF
C70177 NOR2X1_LOC_398/Y NOR2X1_LOC_38/B 0.01fF
C70178 INVX1_LOC_2/A INVX1_LOC_4/A 2.80fF
C70179 NOR2X1_LOC_818/Y INVX1_LOC_4/A 0.14fF
C70180 INVX1_LOC_148/Y NOR2X1_LOC_691/B 0.01fF
C70181 NAND2X1_LOC_276/Y INVX1_LOC_23/Y 0.07fF
C70182 NOR2X1_LOC_427/Y NOR2X1_LOC_51/A 0.04fF
C70183 NAND2X1_LOC_794/B NAND2X1_LOC_733/Y 0.20fF
C70184 INVX1_LOC_81/A INVX1_LOC_23/A 0.03fF
C70185 NAND2X1_LOC_53/Y INVX1_LOC_1/A 3.80fF
C70186 NOR2X1_LOC_226/A INVX1_LOC_4/A 0.34fF
C70187 NOR2X1_LOC_269/Y INVX1_LOC_38/A 0.07fF
C70188 NAND2X1_LOC_724/Y INVX1_LOC_209/Y 0.03fF
C70189 INVX1_LOC_233/A NAND2X1_LOC_198/B 0.10fF
C70190 NOR2X1_LOC_392/B INVX1_LOC_26/A 0.10fF
C70191 NOR2X1_LOC_361/B NAND2X1_LOC_357/A 0.02fF
C70192 INVX1_LOC_256/A NOR2X1_LOC_666/Y 0.00fF
C70193 INVX1_LOC_71/A NOR2X1_LOC_717/A 0.12fF
C70194 NOR2X1_LOC_349/A INVX1_LOC_9/A 0.11fF
C70195 NOR2X1_LOC_111/A INVX1_LOC_76/A 0.12fF
C70196 INVX1_LOC_90/A NOR2X1_LOC_36/B 0.11fF
C70197 INVX1_LOC_196/Y INVX1_LOC_19/A 0.03fF
C70198 INVX1_LOC_58/A NOR2X1_LOC_718/Y 0.03fF
C70199 NOR2X1_LOC_405/A INVX1_LOC_9/A 0.01fF
C70200 INPUT_3 INVX1_LOC_14/A 3.93fF
C70201 NAND2X1_LOC_794/B INVX1_LOC_217/A 0.02fF
C70202 NAND2X1_LOC_860/A NOR2X1_LOC_716/B 0.40fF
C70203 NOR2X1_LOC_730/Y INVX1_LOC_15/A 0.15fF
C70204 INVX1_LOC_30/A NAND2X1_LOC_475/a_36_24# 0.01fF
C70205 INVX1_LOC_50/A NOR2X1_LOC_309/Y 0.01fF
C70206 NAND2X1_LOC_663/a_36_24# NOR2X1_LOC_467/A 0.00fF
C70207 INVX1_LOC_64/A INVX1_LOC_49/A 0.13fF
C70208 NOR2X1_LOC_180/B INVX1_LOC_99/A 0.20fF
C70209 NAND2X1_LOC_803/B NOR2X1_LOC_816/A 0.15fF
C70210 NAND2X1_LOC_374/Y INVX1_LOC_23/Y 0.20fF
C70211 NOR2X1_LOC_65/B NAND2X1_LOC_342/Y 0.01fF
C70212 NOR2X1_LOC_171/Y INVX1_LOC_272/A 0.04fF
C70213 INVX1_LOC_143/A NOR2X1_LOC_843/B 0.09fF
C70214 INVX1_LOC_299/A NOR2X1_LOC_500/B 0.03fF
C70215 NAND2X1_LOC_592/a_36_24# INVX1_LOC_78/A 0.00fF
C70216 NOR2X1_LOC_802/A INVX1_LOC_23/A 0.12fF
C70217 NOR2X1_LOC_590/A NAND2X1_LOC_337/B 0.24fF
C70218 INVX1_LOC_20/A INVX1_LOC_118/A 0.36fF
C70219 NOR2X1_LOC_226/A NAND2X1_LOC_420/a_36_24# 0.00fF
C70220 NOR2X1_LOC_590/A NOR2X1_LOC_816/A 0.15fF
C70221 NOR2X1_LOC_68/A NAND2X1_LOC_326/A 0.98fF
C70222 NOR2X1_LOC_857/A INVX1_LOC_9/A 0.22fF
C70223 INVX1_LOC_21/A NOR2X1_LOC_106/Y 0.60fF
C70224 INVX1_LOC_35/A NAND2X1_LOC_563/Y 0.04fF
C70225 NOR2X1_LOC_684/Y INVX1_LOC_117/A 0.18fF
C70226 INVX1_LOC_150/A INVX1_LOC_4/Y 0.01fF
C70227 INVX1_LOC_36/A NAND2X1_LOC_227/Y 0.03fF
C70228 INPUT_1 INVX1_LOC_4/A 5.61fF
C70229 INVX1_LOC_89/A INVX1_LOC_4/Y 0.24fF
C70230 NAND2X1_LOC_559/Y NAND2X1_LOC_866/A 0.18fF
C70231 INVX1_LOC_2/A INVX1_LOC_64/A 2.27fF
C70232 NOR2X1_LOC_156/a_36_216# INVX1_LOC_37/A 0.00fF
C70233 INVX1_LOC_25/A INVX1_LOC_226/Y 0.02fF
C70234 INVX1_LOC_13/A NOR2X1_LOC_383/B 0.01fF
C70235 INVX1_LOC_282/A NOR2X1_LOC_754/A 0.03fF
C70236 INVX1_LOC_178/A NAND2X1_LOC_354/B 0.14fF
C70237 NOR2X1_LOC_608/a_36_216# NOR2X1_LOC_392/Y 0.01fF
C70238 NAND2X1_LOC_773/Y NAND2X1_LOC_786/a_36_24# 0.06fF
C70239 INVX1_LOC_24/A NAND2X1_LOC_799/A 0.12fF
C70240 INVX1_LOC_13/Y NOR2X1_LOC_315/Y 0.00fF
C70241 INVX1_LOC_64/A NOR2X1_LOC_226/A 0.08fF
C70242 NOR2X1_LOC_287/A NOR2X1_LOC_598/B 0.02fF
C70243 NOR2X1_LOC_656/a_36_216# INPUT_3 0.00fF
C70244 NOR2X1_LOC_45/B NOR2X1_LOC_48/Y 0.00fF
C70245 INVX1_LOC_303/A NOR2X1_LOC_538/B 0.03fF
C70246 INVX1_LOC_58/A INVX1_LOC_30/Y 0.00fF
C70247 NOR2X1_LOC_440/Y INVX1_LOC_57/A 0.03fF
C70248 INVX1_LOC_16/A INVX1_LOC_53/A 0.07fF
C70249 NOR2X1_LOC_791/B INVX1_LOC_31/A 0.05fF
C70250 INVX1_LOC_268/A NOR2X1_LOC_598/B 0.00fF
C70251 INVX1_LOC_41/A NOR2X1_LOC_468/Y 0.12fF
C70252 NAND2X1_LOC_9/Y NOR2X1_LOC_619/A 0.11fF
C70253 NOR2X1_LOC_426/Y INVX1_LOC_72/A 0.36fF
C70254 INVX1_LOC_223/Y INVX1_LOC_177/A 0.00fF
C70255 D_INPUT_0 NOR2X1_LOC_720/A 0.03fF
C70256 INVX1_LOC_233/A INVX1_LOC_53/Y 0.12fF
C70257 INVX1_LOC_90/A INVX1_LOC_26/A 0.10fF
C70258 NOR2X1_LOC_626/Y NOR2X1_LOC_627/a_36_216# 0.00fF
C70259 NOR2X1_LOC_632/Y INVX1_LOC_259/Y 0.11fF
C70260 INVX1_LOC_40/Y NOR2X1_LOC_554/B 0.03fF
C70261 INVX1_LOC_64/A NOR2X1_LOC_218/Y 0.01fF
C70262 INVX1_LOC_21/A NAND2X1_LOC_675/a_36_24# 0.00fF
C70263 INVX1_LOC_25/A INVX1_LOC_10/A 0.35fF
C70264 NOR2X1_LOC_160/B INVX1_LOC_314/Y 0.26fF
C70265 NAND2X1_LOC_214/B NAND2X1_LOC_563/A 0.02fF
C70266 NOR2X1_LOC_488/Y NAND2X1_LOC_552/A 0.00fF
C70267 NAND2X1_LOC_579/A INVX1_LOC_240/A 0.10fF
C70268 INVX1_LOC_224/A NOR2X1_LOC_264/Y 0.00fF
C70269 D_INPUT_0 INVX1_LOC_129/A 0.03fF
C70270 NOR2X1_LOC_468/Y NAND2X1_LOC_477/A 0.03fF
C70271 INVX1_LOC_223/A NOR2X1_LOC_168/Y 0.00fF
C70272 NOR2X1_LOC_567/B INVX1_LOC_18/Y 0.11fF
C70273 NAND2X1_LOC_788/a_36_24# INVX1_LOC_248/A 0.00fF
C70274 INVX1_LOC_48/A INVX1_LOC_32/A 0.08fF
C70275 NOR2X1_LOC_536/A NAND2X1_LOC_243/a_36_24# 0.00fF
C70276 NAND2X1_LOC_549/a_36_24# NOR2X1_LOC_530/Y 0.01fF
C70277 INVX1_LOC_67/Y INVX1_LOC_78/A 0.01fF
C70278 NOR2X1_LOC_189/A NAND2X1_LOC_733/Y 0.01fF
C70279 NAND2X1_LOC_149/Y NOR2X1_LOC_78/B 0.09fF
C70280 NOR2X1_LOC_214/B INVX1_LOC_105/Y 0.28fF
C70281 INVX1_LOC_55/Y NOR2X1_LOC_383/B 0.59fF
C70282 INVX1_LOC_45/A NOR2X1_LOC_13/Y 0.15fF
C70283 NOR2X1_LOC_658/Y INVX1_LOC_71/A 0.07fF
C70284 INVX1_LOC_64/A NAND2X1_LOC_462/B 0.78fF
C70285 INVX1_LOC_269/A INVX1_LOC_206/A 0.02fF
C70286 NOR2X1_LOC_532/Y INVX1_LOC_23/A 0.01fF
C70287 INVX1_LOC_292/A NOR2X1_LOC_551/B 0.01fF
C70288 NAND2X1_LOC_63/Y INVX1_LOC_20/A 0.06fF
C70289 INVX1_LOC_244/A INVX1_LOC_296/A 0.04fF
C70290 INVX1_LOC_7/A INVX1_LOC_138/Y 0.01fF
C70291 NOR2X1_LOC_471/Y NOR2X1_LOC_770/B 0.00fF
C70292 INVX1_LOC_286/Y NOR2X1_LOC_577/Y 0.07fF
C70293 NOR2X1_LOC_123/B NOR2X1_LOC_717/A 0.00fF
C70294 NAND2X1_LOC_348/A INVX1_LOC_26/A 0.04fF
C70295 INVX1_LOC_269/A NAND2X1_LOC_570/Y 0.01fF
C70296 INVX1_LOC_24/A INVX1_LOC_18/A 0.38fF
C70297 GATE_741 NAND2X1_LOC_863/B 0.07fF
C70298 NOR2X1_LOC_831/B INVX1_LOC_54/A 0.10fF
C70299 INVX1_LOC_45/A NAND2X1_LOC_364/Y 0.03fF
C70300 NOR2X1_LOC_67/A NAND2X1_LOC_561/B 0.88fF
C70301 INVX1_LOC_2/Y NOR2X1_LOC_664/a_36_216# 0.00fF
C70302 INVX1_LOC_5/A NOR2X1_LOC_763/Y -0.04fF
C70303 NOR2X1_LOC_474/A INVX1_LOC_195/A 0.01fF
C70304 INVX1_LOC_258/Y NAND2X1_LOC_735/B 0.01fF
C70305 NOR2X1_LOC_65/B INVX1_LOC_67/Y 0.02fF
C70306 NOR2X1_LOC_189/A INVX1_LOC_217/A 0.02fF
C70307 NOR2X1_LOC_15/Y NAND2X1_LOC_194/a_36_24# 0.00fF
C70308 NOR2X1_LOC_506/Y NOR2X1_LOC_697/Y 0.01fF
C70309 INVX1_LOC_64/A NAND2X1_LOC_648/A 0.02fF
C70310 NOR2X1_LOC_124/A INVX1_LOC_3/Y 0.03fF
C70311 VDD NAND2X1_LOC_291/B 0.63fF
C70312 INVX1_LOC_226/Y INVX1_LOC_1/A 0.01fF
C70313 NOR2X1_LOC_272/Y NOR2X1_LOC_561/Y 0.01fF
C70314 INVX1_LOC_28/A INVX1_LOC_53/A 0.75fF
C70315 INVX1_LOC_64/A INPUT_1 0.05fF
C70316 INVX1_LOC_44/A INVX1_LOC_19/A 0.03fF
C70317 INVX1_LOC_50/A NOR2X1_LOC_208/A 0.05fF
C70318 INVX1_LOC_115/A NOR2X1_LOC_477/B 0.03fF
C70319 NOR2X1_LOC_550/a_36_216# INVX1_LOC_104/A 0.00fF
C70320 INVX1_LOC_314/A INVX1_LOC_15/A 0.06fF
C70321 NOR2X1_LOC_71/Y NOR2X1_LOC_291/Y 0.00fF
C70322 NOR2X1_LOC_93/Y INVX1_LOC_234/A 0.03fF
C70323 NOR2X1_LOC_361/B INVX1_LOC_25/Y 0.01fF
C70324 NAND2X1_LOC_794/B NAND2X1_LOC_808/A 0.07fF
C70325 VDD GATE_222 0.18fF
C70326 INVX1_LOC_235/Y NOR2X1_LOC_459/A 0.24fF
C70327 INVX1_LOC_11/A NAND2X1_LOC_452/a_36_24# 0.00fF
C70328 INVX1_LOC_172/A INVX1_LOC_24/A 0.03fF
C70329 NOR2X1_LOC_15/Y NAND2X1_LOC_390/A 0.58fF
C70330 NOR2X1_LOC_860/Y NAND2X1_LOC_206/Y 0.05fF
C70331 VDD INVX1_LOC_283/A 0.00fF
C70332 NOR2X1_LOC_361/B NAND2X1_LOC_349/B 0.10fF
C70333 NOR2X1_LOC_778/B NOR2X1_LOC_160/B 0.09fF
C70334 INVX1_LOC_284/Y NAND2X1_LOC_722/A 0.00fF
C70335 NOR2X1_LOC_832/a_36_216# NOR2X1_LOC_841/A 0.00fF
C70336 NAND2X1_LOC_149/Y INVX1_LOC_83/A 0.11fF
C70337 NAND2X1_LOC_567/Y NOR2X1_LOC_152/Y 0.01fF
C70338 NOR2X1_LOC_828/B INVX1_LOC_213/A 0.07fF
C70339 INVX1_LOC_27/A NOR2X1_LOC_214/B 0.11fF
C70340 INVX1_LOC_69/Y INVX1_LOC_57/A 0.03fF
C70341 NOR2X1_LOC_215/Y INVX1_LOC_63/Y 0.03fF
C70342 NOR2X1_LOC_794/B NOR2X1_LOC_500/Y 0.50fF
C70343 INVX1_LOC_1/A INVX1_LOC_10/A 0.01fF
C70344 NOR2X1_LOC_168/Y INVX1_LOC_149/Y 0.02fF
C70345 NOR2X1_LOC_641/Y INVX1_LOC_19/A 0.00fF
C70346 NOR2X1_LOC_637/B NOR2X1_LOC_433/A 0.00fF
C70347 NOR2X1_LOC_226/A NAND2X1_LOC_860/a_36_24# 0.01fF
C70348 NOR2X1_LOC_189/A NAND2X1_LOC_787/B 0.00fF
C70349 NAND2X1_LOC_363/B NOR2X1_LOC_97/A 0.07fF
C70350 NOR2X1_LOC_820/Y NOR2X1_LOC_649/B 0.04fF
C70351 NOR2X1_LOC_68/A NOR2X1_LOC_87/B 0.00fF
C70352 NOR2X1_LOC_51/A NOR2X1_LOC_36/B 0.52fF
C70353 INVX1_LOC_45/A INVX1_LOC_256/Y 0.33fF
C70354 INVX1_LOC_217/A NOR2X1_LOC_482/Y 0.09fF
C70355 NOR2X1_LOC_646/A INVX1_LOC_31/A 0.16fF
C70356 NOR2X1_LOC_335/A NAND2X1_LOC_310/a_36_24# 0.02fF
C70357 NOR2X1_LOC_817/Y NOR2X1_LOC_128/B 0.02fF
C70358 INVX1_LOC_286/Y INVX1_LOC_22/A 0.07fF
C70359 INVX1_LOC_174/A INPUT_5 0.51fF
C70360 NOR2X1_LOC_207/A NOR2X1_LOC_596/A 0.02fF
C70361 INVX1_LOC_24/A INVX1_LOC_34/Y 0.51fF
C70362 INVX1_LOC_114/A NOR2X1_LOC_467/A 0.04fF
C70363 INVX1_LOC_289/A INVX1_LOC_72/A 0.03fF
C70364 INVX1_LOC_19/A NOR2X1_LOC_461/B 0.03fF
C70365 INVX1_LOC_202/A INVX1_LOC_133/Y 0.01fF
C70366 INVX1_LOC_41/A NOR2X1_LOC_295/Y 0.00fF
C70367 INVX1_LOC_58/A NOR2X1_LOC_124/A 0.16fF
C70368 NOR2X1_LOC_360/Y INVX1_LOC_40/A 0.03fF
C70369 INVX1_LOC_1/A NOR2X1_LOC_302/Y 0.05fF
C70370 NOR2X1_LOC_52/B INVX1_LOC_155/A 0.04fF
C70371 INVX1_LOC_310/A INVX1_LOC_303/A 0.01fF
C70372 INVX1_LOC_269/A NOR2X1_LOC_19/B 0.42fF
C70373 NOR2X1_LOC_831/B NAND2X1_LOC_807/B 0.00fF
C70374 INVX1_LOC_256/Y INVX1_LOC_71/A 0.16fF
C70375 NOR2X1_LOC_632/Y INVX1_LOC_136/A 0.00fF
C70376 NOR2X1_LOC_357/Y NOR2X1_LOC_383/B 0.01fF
C70377 NAND2X1_LOC_802/A INVX1_LOC_144/Y 0.01fF
C70378 INVX1_LOC_271/A NAND2X1_LOC_434/a_36_24# 0.00fF
C70379 INVX1_LOC_47/Y NOR2X1_LOC_489/A 0.01fF
C70380 INVX1_LOC_159/A INVX1_LOC_22/A 0.07fF
C70381 INVX1_LOC_49/A INVX1_LOC_44/Y 0.02fF
C70382 INVX1_LOC_128/Y NOR2X1_LOC_331/B 0.03fF
C70383 INVX1_LOC_135/A INVX1_LOC_141/Y 0.01fF
C70384 INPUT_2 NOR2X1_LOC_5/a_36_216# 0.00fF
C70385 D_INPUT_0 NOR2X1_LOC_514/A 0.00fF
C70386 NOR2X1_LOC_773/a_36_216# NOR2X1_LOC_309/Y 0.00fF
C70387 INVX1_LOC_43/Y INPUT_1 0.03fF
C70388 NOR2X1_LOC_757/A INVX1_LOC_72/A 0.07fF
C70389 NOR2X1_LOC_160/B NOR2X1_LOC_724/Y 0.01fF
C70390 INVX1_LOC_90/A INVX1_LOC_141/A 0.01fF
C70391 INVX1_LOC_229/A INVX1_LOC_282/A 0.00fF
C70392 INVX1_LOC_33/A NAND2X1_LOC_451/Y 0.07fF
C70393 NAND2X1_LOC_9/Y NAND2X1_LOC_465/A 0.05fF
C70394 NOR2X1_LOC_561/Y NAND2X1_LOC_364/A 0.03fF
C70395 NOR2X1_LOC_778/B NOR2X1_LOC_544/a_36_216# 0.00fF
C70396 NAND2X1_LOC_727/a_36_24# INVX1_LOC_28/A 0.00fF
C70397 NOR2X1_LOC_561/A INVX1_LOC_26/A 0.03fF
C70398 NOR2X1_LOC_294/Y INVX1_LOC_135/A 0.16fF
C70399 NAND2X1_LOC_428/a_36_24# NOR2X1_LOC_467/A 0.01fF
C70400 INVX1_LOC_53/A NOR2X1_LOC_35/Y 0.10fF
C70401 INVX1_LOC_35/A NOR2X1_LOC_833/Y 0.16fF
C70402 INVX1_LOC_27/A NOR2X1_LOC_741/A 0.03fF
C70403 NAND2X1_LOC_740/B INVX1_LOC_161/Y 0.13fF
C70404 NAND2X1_LOC_783/A INVX1_LOC_18/A 0.01fF
C70405 INVX1_LOC_285/A INVX1_LOC_42/A 0.08fF
C70406 NOR2X1_LOC_690/A NOR2X1_LOC_667/A 0.03fF
C70407 INVX1_LOC_200/Y NAND2X1_LOC_721/A 0.03fF
C70408 INVX1_LOC_233/Y NOR2X1_LOC_24/Y 0.02fF
C70409 INVX1_LOC_12/Y INVX1_LOC_271/A 0.02fF
C70410 NAND2X1_LOC_860/A NAND2X1_LOC_633/Y 0.10fF
C70411 NAND2X1_LOC_778/Y NAND2X1_LOC_623/B 0.12fF
C70412 INVX1_LOC_18/A NOR2X1_LOC_130/A 0.03fF
C70413 NOR2X1_LOC_89/A NOR2X1_LOC_662/A 0.03fF
C70414 INVX1_LOC_84/A INVX1_LOC_290/Y 0.07fF
C70415 NAND2X1_LOC_728/Y NAND2X1_LOC_800/Y 0.00fF
C70416 INVX1_LOC_304/Y NOR2X1_LOC_482/Y 0.02fF
C70417 NOR2X1_LOC_814/A INVX1_LOC_42/A 0.19fF
C70418 NOR2X1_LOC_132/Y INVX1_LOC_25/Y 0.03fF
C70419 INVX1_LOC_223/Y INVX1_LOC_65/A 0.01fF
C70420 INVX1_LOC_136/A NOR2X1_LOC_246/a_36_216# 0.00fF
C70421 NAND2X1_LOC_361/Y INVX1_LOC_1/Y 0.07fF
C70422 NOR2X1_LOC_627/Y NAND2X1_LOC_629/Y 0.09fF
C70423 INVX1_LOC_11/A INVX1_LOC_86/A 0.00fF
C70424 NOR2X1_LOC_363/Y INVX1_LOC_23/A 0.02fF
C70425 NOR2X1_LOC_434/a_36_216# NOR2X1_LOC_174/B 0.00fF
C70426 NAND2X1_LOC_276/Y INVX1_LOC_232/A 2.51fF
C70427 NOR2X1_LOC_541/Y NOR2X1_LOC_337/A 0.10fF
C70428 D_INPUT_0 INVX1_LOC_41/Y 0.03fF
C70429 NOR2X1_LOC_364/A INVX1_LOC_78/A 1.94fF
C70430 INVX1_LOC_26/Y NOR2X1_LOC_641/Y 0.02fF
C70431 NOR2X1_LOC_155/A INVX1_LOC_271/Y 1.04fF
C70432 INVX1_LOC_32/A NOR2X1_LOC_127/Y 0.06fF
C70433 NAND2X1_LOC_363/B INVX1_LOC_129/Y 0.00fF
C70434 NOR2X1_LOC_828/B NOR2X1_LOC_707/B 0.04fF
C70435 NOR2X1_LOC_637/Y NOR2X1_LOC_130/A 0.32fF
C70436 NOR2X1_LOC_617/Y D_INPUT_0 0.03fF
C70437 INVX1_LOC_2/A NAND2X1_LOC_850/Y 0.07fF
C70438 NOR2X1_LOC_434/A INVX1_LOC_117/A 0.01fF
C70439 INVX1_LOC_39/A INVX1_LOC_20/A 0.00fF
C70440 NOR2X1_LOC_272/Y INVX1_LOC_76/A 0.04fF
C70441 NOR2X1_LOC_510/Y NAND2X1_LOC_453/A 0.02fF
C70442 NOR2X1_LOC_791/Y NAND2X1_LOC_287/B 0.01fF
C70443 INPUT_3 INVX1_LOC_48/A 0.07fF
C70444 INVX1_LOC_34/A NOR2X1_LOC_719/B 0.06fF
C70445 INVX1_LOC_1/A NOR2X1_LOC_711/Y 0.08fF
C70446 NOR2X1_LOC_388/Y NAND2X1_LOC_656/Y 0.07fF
C70447 NAND2X1_LOC_214/B INVX1_LOC_12/Y 0.44fF
C70448 NOR2X1_LOC_331/B NOR2X1_LOC_717/A 0.01fF
C70449 NOR2X1_LOC_542/Y INVX1_LOC_77/A 0.27fF
C70450 INVX1_LOC_78/A INVX1_LOC_285/A 0.16fF
C70451 NOR2X1_LOC_103/a_36_216# INVX1_LOC_23/Y 0.00fF
C70452 INVX1_LOC_234/A NAND2X1_LOC_137/a_36_24# 0.00fF
C70453 NAND2X1_LOC_721/A NOR2X1_LOC_406/A 0.64fF
C70454 INVX1_LOC_95/Y NOR2X1_LOC_271/a_36_216# 0.01fF
C70455 INVX1_LOC_78/A NOR2X1_LOC_814/A 0.10fF
C70456 NOR2X1_LOC_859/Y NOR2X1_LOC_849/A 0.37fF
C70457 NOR2X1_LOC_68/A NOR2X1_LOC_74/a_36_216# 0.00fF
C70458 NOR2X1_LOC_160/B NOR2X1_LOC_557/A 0.02fF
C70459 NOR2X1_LOC_778/B NOR2X1_LOC_516/B 0.03fF
C70460 NAND2X1_LOC_213/A INVX1_LOC_76/A 0.02fF
C70461 NOR2X1_LOC_78/B INVX1_LOC_16/A 0.07fF
C70462 INVX1_LOC_27/A INVX1_LOC_12/Y 0.10fF
C70463 INVX1_LOC_77/A INVX1_LOC_311/Y 0.08fF
C70464 NOR2X1_LOC_220/A NOR2X1_LOC_211/A 0.12fF
C70465 NAND2X1_LOC_63/Y INVX1_LOC_4/A 0.29fF
C70466 NOR2X1_LOC_536/A INVX1_LOC_306/Y 0.03fF
C70467 INVX1_LOC_64/A INVX1_LOC_118/A 0.14fF
C70468 NOR2X1_LOC_15/Y NOR2X1_LOC_314/Y 0.02fF
C70469 NOR2X1_LOC_68/A NOR2X1_LOC_527/Y 0.02fF
C70470 NOR2X1_LOC_433/A NAND2X1_LOC_850/A 0.00fF
C70471 INVX1_LOC_174/A NOR2X1_LOC_448/A -0.03fF
C70472 NOR2X1_LOC_92/Y NOR2X1_LOC_447/B 0.02fF
C70473 NOR2X1_LOC_568/a_36_216# INVX1_LOC_22/A 0.00fF
C70474 NOR2X1_LOC_65/B INVX1_LOC_285/A 0.10fF
C70475 NOR2X1_LOC_48/B NAND2X1_LOC_430/B 0.17fF
C70476 NOR2X1_LOC_178/Y INVX1_LOC_127/A 0.01fF
C70477 INVX1_LOC_89/A INVX1_LOC_82/A 0.06fF
C70478 INVX1_LOC_1/A INVX1_LOC_178/Y 0.00fF
C70479 NOR2X1_LOC_160/B NOR2X1_LOC_657/B 0.05fF
C70480 NAND2X1_LOC_352/B INVX1_LOC_95/A 0.05fF
C70481 INVX1_LOC_255/Y NOR2X1_LOC_382/a_36_216# 0.01fF
C70482 NOR2X1_LOC_798/A NOR2X1_LOC_652/a_36_216# 0.00fF
C70483 INVX1_LOC_135/A NOR2X1_LOC_168/B 0.03fF
C70484 NOR2X1_LOC_65/B NOR2X1_LOC_814/A 0.01fF
C70485 INVX1_LOC_33/A NOR2X1_LOC_567/B 0.02fF
C70486 NOR2X1_LOC_15/Y INVX1_LOC_117/A 0.93fF
C70487 INVX1_LOC_193/Y NOR2X1_LOC_705/a_36_216# 0.00fF
C70488 NOR2X1_LOC_219/B NOR2X1_LOC_202/Y 0.28fF
C70489 NAND2X1_LOC_354/B INVX1_LOC_140/A 0.03fF
C70490 NOR2X1_LOC_366/B NAND2X1_LOC_656/Y 0.08fF
C70491 INVX1_LOC_50/A INVX1_LOC_63/A 0.10fF
C70492 NAND2X1_LOC_243/Y NOR2X1_LOC_291/Y 0.14fF
C70493 NOR2X1_LOC_703/B NOR2X1_LOC_78/A 0.03fF
C70494 NOR2X1_LOC_332/A NAND2X1_LOC_819/Y 0.03fF
C70495 INVX1_LOC_256/Y NOR2X1_LOC_123/B 0.16fF
C70496 INVX1_LOC_34/A INVX1_LOC_73/A 0.07fF
C70497 NAND2X1_LOC_746/a_36_24# INVX1_LOC_117/Y 0.00fF
C70498 NOR2X1_LOC_389/B INVX1_LOC_149/A 0.02fF
C70499 NAND2X1_LOC_61/Y NAND2X1_LOC_74/B 0.03fF
C70500 NOR2X1_LOC_105/Y INVX1_LOC_63/A 0.01fF
C70501 NOR2X1_LOC_91/Y NOR2X1_LOC_45/B 0.04fF
C70502 NAND2X1_LOC_93/B INVX1_LOC_306/Y 0.25fF
C70503 NOR2X1_LOC_299/Y NAND2X1_LOC_863/B 6.64fF
C70504 NAND2X1_LOC_850/Y INPUT_1 0.15fF
C70505 NAND2X1_LOC_704/a_36_24# INVX1_LOC_118/A 0.00fF
C70506 INVX1_LOC_229/Y NAND2X1_LOC_735/B 0.01fF
C70507 INVX1_LOC_31/A INVX1_LOC_2/Y 0.09fF
C70508 NOR2X1_LOC_609/Y NAND2X1_LOC_647/B 0.10fF
C70509 INVX1_LOC_135/A NOR2X1_LOC_789/A 0.00fF
C70510 NOR2X1_LOC_78/B INVX1_LOC_28/A 0.15fF
C70511 NOR2X1_LOC_585/a_36_216# NOR2X1_LOC_586/Y 0.01fF
C70512 INVX1_LOC_75/A INVX1_LOC_177/A 0.03fF
C70513 INVX1_LOC_31/A INVX1_LOC_37/Y 0.03fF
C70514 INVX1_LOC_30/A NAND2X1_LOC_287/B 0.10fF
C70515 INVX1_LOC_190/Y INVX1_LOC_22/A 0.04fF
C70516 INVX1_LOC_39/Y NOR2X1_LOC_813/Y 0.06fF
C70517 NAND2X1_LOC_563/A NOR2X1_LOC_19/B 0.02fF
C70518 NOR2X1_LOC_89/A INVX1_LOC_57/A 0.18fF
C70519 INVX1_LOC_41/A INVX1_LOC_100/Y 0.02fF
C70520 NAND2X1_LOC_364/A INVX1_LOC_76/A 0.10fF
C70521 INVX1_LOC_25/A INVX1_LOC_12/A 0.07fF
C70522 NAND2X1_LOC_842/B INVX1_LOC_53/Y 0.02fF
C70523 VDD NOR2X1_LOC_274/B 0.02fF
C70524 INVX1_LOC_61/Y NOR2X1_LOC_102/a_36_216# 0.01fF
C70525 INVX1_LOC_61/A INVX1_LOC_20/A 0.04fF
C70526 INVX1_LOC_3/A INVX1_LOC_306/Y 0.03fF
C70527 INVX1_LOC_208/A NAND2X1_LOC_123/Y 0.07fF
C70528 INVX1_LOC_72/A INVX1_LOC_37/A 0.07fF
C70529 INVX1_LOC_33/A NOR2X1_LOC_269/Y 0.07fF
C70530 INVX1_LOC_53/A INVX1_LOC_109/A 0.00fF
C70531 NAND2X1_LOC_785/A NOR2X1_LOC_167/Y 0.01fF
C70532 INVX1_LOC_141/A INVX1_LOC_38/A 0.01fF
C70533 NOR2X1_LOC_488/Y INVX1_LOC_140/A 0.01fF
C70534 INVX1_LOC_39/Y INVX1_LOC_280/A 0.15fF
C70535 INVX1_LOC_64/A NAND2X1_LOC_63/Y 0.39fF
C70536 INVX1_LOC_1/A NOR2X1_LOC_445/B 0.03fF
C70537 INVX1_LOC_43/Y INVX1_LOC_118/A -0.01fF
C70538 NOR2X1_LOC_859/A NOR2X1_LOC_859/Y 0.04fF
C70539 INVX1_LOC_269/A NOR2X1_LOC_216/B 0.07fF
C70540 NOR2X1_LOC_721/Y NOR2X1_LOC_346/B 0.18fF
C70541 NAND2X1_LOC_162/A INVX1_LOC_75/A 0.03fF
C70542 INVX1_LOC_32/A NOR2X1_LOC_383/B 0.03fF
C70543 NAND2X1_LOC_17/a_36_24# NAND2X1_LOC_1/Y 0.00fF
C70544 INVX1_LOC_34/A NAND2X1_LOC_729/B 0.04fF
C70545 INVX1_LOC_135/A INVX1_LOC_132/Y 0.04fF
C70546 INVX1_LOC_198/Y INVX1_LOC_37/A 0.09fF
C70547 NOR2X1_LOC_454/Y INVX1_LOC_84/A 0.46fF
C70548 NAND2X1_LOC_218/B VDD 0.01fF
C70549 INVX1_LOC_26/A NAND2X1_LOC_223/A 0.03fF
C70550 NOR2X1_LOC_294/Y INVX1_LOC_280/A 0.06fF
C70551 NOR2X1_LOC_577/Y NOR2X1_LOC_136/a_36_216# 0.00fF
C70552 NOR2X1_LOC_413/Y INVX1_LOC_255/A 0.02fF
C70553 NOR2X1_LOC_500/Y NOR2X1_LOC_188/A 0.03fF
C70554 INVX1_LOC_35/A NOR2X1_LOC_114/Y 0.32fF
C70555 INVX1_LOC_226/Y NOR2X1_LOC_188/A 0.03fF
C70556 NAND2X1_LOC_112/Y INVX1_LOC_79/A 0.01fF
C70557 INVX1_LOC_246/A INVX1_LOC_92/A 0.07fF
C70558 NOR2X1_LOC_794/B INVX1_LOC_307/A 0.01fF
C70559 INVX1_LOC_21/A INVX1_LOC_262/Y 0.01fF
C70560 INVX1_LOC_83/A INVX1_LOC_28/A 0.03fF
C70561 NOR2X1_LOC_763/Y NAND2X1_LOC_651/a_36_24# 0.01fF
C70562 NAND2X1_LOC_357/B INVX1_LOC_95/A 0.01fF
C70563 INVX1_LOC_226/Y NOR2X1_LOC_548/B 0.03fF
C70564 NOR2X1_LOC_577/Y VDD 2.33fF
C70565 INVX1_LOC_5/A NOR2X1_LOC_67/Y 0.07fF
C70566 NOR2X1_LOC_689/A NAND2X1_LOC_175/Y 0.03fF
C70567 NOR2X1_LOC_379/Y VDD 0.01fF
C70568 INVX1_LOC_136/A NOR2X1_LOC_186/a_36_216# 0.01fF
C70569 NOR2X1_LOC_168/B NOR2X1_LOC_552/A 0.07fF
C70570 INVX1_LOC_153/A INVX1_LOC_14/Y 0.02fF
C70571 NOR2X1_LOC_577/Y NAND2X1_LOC_800/A 0.05fF
C70572 NAND2X1_LOC_371/a_36_24# INVX1_LOC_38/A 0.01fF
C70573 INVX1_LOC_41/Y NAND2X1_LOC_848/A 0.01fF
C70574 INVX1_LOC_45/A NOR2X1_LOC_640/Y 0.07fF
C70575 INVX1_LOC_201/Y NAND2X1_LOC_414/a_36_24# 0.01fF
C70576 NOR2X1_LOC_568/A NOR2X1_LOC_640/Y 0.36fF
C70577 NAND2X1_LOC_169/Y NOR2X1_LOC_48/B 0.02fF
C70578 NOR2X1_LOC_13/Y NOR2X1_LOC_331/B 0.10fF
C70579 NAND2X1_LOC_308/Y NOR2X1_LOC_305/Y 0.00fF
C70580 NOR2X1_LOC_392/Y INVX1_LOC_4/Y 0.07fF
C70581 NOR2X1_LOC_629/B VDD -0.00fF
C70582 NAND2X1_LOC_738/B NAND2X1_LOC_175/Y 0.02fF
C70583 NOR2X1_LOC_598/B INVX1_LOC_271/Y 0.10fF
C70584 NOR2X1_LOC_249/a_36_216# NAND2X1_LOC_574/A 0.01fF
C70585 NOR2X1_LOC_348/B VDD 0.51fF
C70586 INVX1_LOC_135/A NAND2X1_LOC_622/B 0.03fF
C70587 NAND2X1_LOC_35/Y NOR2X1_LOC_38/B 0.00fF
C70588 NAND2X1_LOC_555/Y NOR2X1_LOC_673/A 0.08fF
C70589 INVX1_LOC_1/A INVX1_LOC_12/A 1.96fF
C70590 NAND2X1_LOC_717/Y NAND2X1_LOC_836/a_36_24# -0.00fF
C70591 INVX1_LOC_27/A NOR2X1_LOC_554/A 0.05fF
C70592 INPUT_0 NOR2X1_LOC_76/A 0.01fF
C70593 INVX1_LOC_34/A NOR2X1_LOC_122/a_36_216# 0.00fF
C70594 NOR2X1_LOC_78/B NOR2X1_LOC_35/Y 0.05fF
C70595 NOR2X1_LOC_666/Y NOR2X1_LOC_89/A 0.81fF
C70596 NAND2X1_LOC_357/A NAND2X1_LOC_81/B 0.10fF
C70597 INVX1_LOC_18/A NOR2X1_LOC_197/B 0.10fF
C70598 INVX1_LOC_259/A INVX1_LOC_14/Y 0.03fF
C70599 NOR2X1_LOC_180/B INPUT_0 0.39fF
C70600 INVX1_LOC_61/Y INVX1_LOC_63/A 0.07fF
C70601 INVX1_LOC_90/A NOR2X1_LOC_313/Y 0.01fF
C70602 INVX1_LOC_10/Y INVX1_LOC_88/Y 0.15fF
C70603 NAND2X1_LOC_717/Y INVX1_LOC_46/A 0.03fF
C70604 NOR2X1_LOC_502/Y NOR2X1_LOC_509/A 0.11fF
C70605 NOR2X1_LOC_254/A INVX1_LOC_19/A 0.67fF
C70606 NAND2X1_LOC_175/B NOR2X1_LOC_331/B 0.31fF
C70607 INVX1_LOC_294/Y NOR2X1_LOC_536/A 0.02fF
C70608 INVX1_LOC_103/Y INVX1_LOC_38/A 0.02fF
C70609 INVX1_LOC_39/A INVX1_LOC_4/A 0.03fF
C70610 INVX1_LOC_22/A NOR2X1_LOC_56/Y 0.10fF
C70611 NOR2X1_LOC_537/Y INVX1_LOC_37/A 0.07fF
C70612 INVX1_LOC_179/Y NOR2X1_LOC_857/A 0.01fF
C70613 INVX1_LOC_16/A NOR2X1_LOC_164/Y 0.07fF
C70614 NAND2X1_LOC_338/B INVX1_LOC_37/A 0.10fF
C70615 NOR2X1_LOC_289/a_36_216# INVX1_LOC_76/A 0.00fF
C70616 NOR2X1_LOC_445/Y INVX1_LOC_9/A 0.07fF
C70617 INVX1_LOC_23/A NOR2X1_LOC_809/A 0.04fF
C70618 NOR2X1_LOC_113/B NAND2X1_LOC_842/B 0.01fF
C70619 INVX1_LOC_24/A NAND2X1_LOC_489/a_36_24# 0.00fF
C70620 VDD NOR2X1_LOC_346/B 0.11fF
C70621 NOR2X1_LOC_454/Y INVX1_LOC_15/A 0.07fF
C70622 NOR2X1_LOC_561/Y NOR2X1_LOC_405/A 0.08fF
C70623 NOR2X1_LOC_175/B VDD 0.30fF
C70624 INVX1_LOC_10/A NOR2X1_LOC_43/Y 0.03fF
C70625 NOR2X1_LOC_13/Y NOR2X1_LOC_592/B 0.14fF
C70626 NOR2X1_LOC_445/a_36_216# INVX1_LOC_29/A 0.00fF
C70627 NAND2X1_LOC_569/B INVX1_LOC_23/Y 0.05fF
C70628 NAND2X1_LOC_325/a_36_24# NAND2X1_LOC_807/Y 0.01fF
C70629 INVX1_LOC_23/A INVX1_LOC_29/Y 0.06fF
C70630 NOR2X1_LOC_589/A NAND2X1_LOC_212/Y 0.06fF
C70631 NAND2X1_LOC_323/B INVX1_LOC_37/A 0.06fF
C70632 NOR2X1_LOC_15/Y INVX1_LOC_3/Y 2.34fF
C70633 INVX1_LOC_266/Y INVX1_LOC_281/Y 0.01fF
C70634 NOR2X1_LOC_298/Y INPUT_4 0.55fF
C70635 INVX1_LOC_188/A INVX1_LOC_29/A 0.01fF
C70636 NOR2X1_LOC_554/B NOR2X1_LOC_814/A 0.05fF
C70637 NOR2X1_LOC_85/a_36_216# INVX1_LOC_20/A 0.00fF
C70638 NAND2X1_LOC_803/B INVX1_LOC_42/A 0.02fF
C70639 NAND2X1_LOC_735/B INVX1_LOC_20/A 0.03fF
C70640 NAND2X1_LOC_352/B NAND2X1_LOC_807/B 0.16fF
C70641 NOR2X1_LOC_615/Y INVX1_LOC_42/A 0.01fF
C70642 INVX1_LOC_16/A INVX1_LOC_46/A 0.31fF
C70643 NAND2X1_LOC_20/B NAND2X1_LOC_223/a_36_24# 0.00fF
C70644 VDD INVX1_LOC_22/A 3.29fF
C70645 NOR2X1_LOC_493/A NOR2X1_LOC_717/A 0.13fF
C70646 NAND2X1_LOC_357/B INVX1_LOC_54/A 0.07fF
C70647 INVX1_LOC_163/A INVX1_LOC_253/A 0.03fF
C70648 INVX1_LOC_207/A INVX1_LOC_241/Y 0.03fF
C70649 INPUT_5 INVX1_LOC_20/A 0.15fF
C70650 NAND2X1_LOC_800/A INVX1_LOC_22/A 0.03fF
C70651 INVX1_LOC_13/Y NAND2X1_LOC_99/A 1.64fF
C70652 NAND2X1_LOC_343/a_36_24# INVX1_LOC_46/A 0.01fF
C70653 INVX1_LOC_75/A INVX1_LOC_285/Y 0.00fF
C70654 INVX1_LOC_38/Y NOR2X1_LOC_843/B 0.39fF
C70655 NOR2X1_LOC_68/A NAND2X1_LOC_219/B 0.01fF
C70656 NOR2X1_LOC_590/A INVX1_LOC_42/A 0.57fF
C70657 NAND2X1_LOC_510/A NOR2X1_LOC_340/A 0.95fF
C70658 NOR2X1_LOC_74/A INVX1_LOC_126/Y 0.03fF
C70659 INVX1_LOC_83/A NOR2X1_LOC_35/Y 0.12fF
C70660 NOR2X1_LOC_142/Y NOR2X1_LOC_831/B 0.00fF
C70661 INVX1_LOC_77/A INVX1_LOC_84/A 0.03fF
C70662 NOR2X1_LOC_329/B NOR2X1_LOC_139/Y 0.01fF
C70663 NOR2X1_LOC_329/B NAND2X1_LOC_655/A 0.07fF
C70664 NAND2X1_LOC_859/Y INVX1_LOC_37/Y 0.01fF
C70665 NOR2X1_LOC_384/Y INVX1_LOC_12/A 0.01fF
C70666 NAND2X1_LOC_850/Y INVX1_LOC_118/A 0.07fF
C70667 INVX1_LOC_171/Y NOR2X1_LOC_383/B 0.03fF
C70668 NOR2X1_LOC_583/a_36_216# INVX1_LOC_77/Y 0.01fF
C70669 NOR2X1_LOC_784/B VDD 0.14fF
C70670 NAND2X1_LOC_306/a_36_24# INVX1_LOC_49/Y 0.00fF
C70671 INVX1_LOC_143/A NAND2X1_LOC_488/a_36_24# 0.00fF
C70672 INVX1_LOC_58/A NAND2X1_LOC_778/Y 0.11fF
C70673 NOR2X1_LOC_665/a_36_216# NOR2X1_LOC_665/Y 0.00fF
C70674 NOR2X1_LOC_789/A INVX1_LOC_280/A 0.02fF
C70675 NAND2X1_LOC_803/B INVX1_LOC_78/A 0.02fF
C70676 INVX1_LOC_283/Y INVX1_LOC_186/Y -0.02fF
C70677 NOR2X1_LOC_795/a_36_216# INVX1_LOC_117/A 0.00fF
C70678 NAND2X1_LOC_794/B INVX1_LOC_53/A 0.03fF
C70679 NAND2X1_LOC_363/B INVX1_LOC_50/Y 0.09fF
C70680 NOR2X1_LOC_577/Y INVX1_LOC_133/A 0.00fF
C70681 NOR2X1_LOC_655/B NOR2X1_LOC_831/B 0.00fF
C70682 INVX1_LOC_313/Y INVX1_LOC_37/A 0.09fF
C70683 NOR2X1_LOC_590/A INVX1_LOC_78/A 0.13fF
C70684 NAND2X1_LOC_727/Y INVX1_LOC_185/A 0.15fF
C70685 INVX1_LOC_28/A INVX1_LOC_46/A 0.22fF
C70686 INVX1_LOC_124/A INVX1_LOC_84/A 2.25fF
C70687 NOR2X1_LOC_848/Y NOR2X1_LOC_105/a_36_216# 0.00fF
C70688 INVX1_LOC_39/A INVX1_LOC_64/A 0.02fF
C70689 NOR2X1_LOC_735/Y VDD -0.00fF
C70690 INVX1_LOC_58/A NOR2X1_LOC_15/Y 0.31fF
C70691 NOR2X1_LOC_192/A INVX1_LOC_6/A 0.02fF
C70692 NOR2X1_LOC_530/Y INVX1_LOC_23/Y 0.00fF
C70693 NOR2X1_LOC_52/B NOR2X1_LOC_662/A 0.05fF
C70694 NOR2X1_LOC_520/B NAND2X1_LOC_74/B 0.11fF
C70695 INVX1_LOC_224/A INVX1_LOC_57/A 0.04fF
C70696 INVX1_LOC_98/A INVX1_LOC_91/A 0.10fF
C70697 INVX1_LOC_290/A INVX1_LOC_92/A 0.03fF
C70698 NAND2X1_LOC_537/Y NOR2X1_LOC_591/A 0.03fF
C70699 INVX1_LOC_11/A INVX1_LOC_57/A 0.31fF
C70700 NOR2X1_LOC_78/A INVX1_LOC_91/A 0.10fF
C70701 NOR2X1_LOC_391/A NOR2X1_LOC_78/Y 0.00fF
C70702 NAND2X1_LOC_149/B NAND2X1_LOC_425/Y 0.03fF
C70703 NOR2X1_LOC_65/B NOR2X1_LOC_590/A 0.04fF
C70704 NOR2X1_LOC_453/Y NOR2X1_LOC_221/a_36_216# 0.00fF
C70705 NOR2X1_LOC_67/A INVX1_LOC_293/Y -0.02fF
C70706 D_INPUT_0 INVX1_LOC_185/A 0.08fF
C70707 NOR2X1_LOC_835/B NOR2X1_LOC_857/A 0.01fF
C70708 NAND2X1_LOC_569/A NAND2X1_LOC_254/Y 0.02fF
C70709 INVX1_LOC_279/A NOR2X1_LOC_155/A 0.07fF
C70710 NOR2X1_LOC_160/B INVX1_LOC_271/A 0.07fF
C70711 INVX1_LOC_77/A INVX1_LOC_15/A 0.79fF
C70712 NAND2X1_LOC_354/B INVX1_LOC_42/A 0.04fF
C70713 NOR2X1_LOC_802/A NOR2X1_LOC_633/A 0.01fF
C70714 D_INPUT_1 INPUT_2 0.17fF
C70715 INPUT_6 NAND2X1_LOC_30/Y 0.08fF
C70716 INVX1_LOC_85/Y NOR2X1_LOC_209/B 0.21fF
C70717 NAND2X1_LOC_357/B NAND2X1_LOC_807/B 0.16fF
C70718 INVX1_LOC_100/A VDD 0.08fF
C70719 NOR2X1_LOC_367/B INVX1_LOC_109/Y 0.04fF
C70720 INVX1_LOC_246/A INVX1_LOC_53/A 0.08fF
C70721 NOR2X1_LOC_315/Y NOR2X1_LOC_76/B 0.02fF
C70722 NAND2X1_LOC_357/B NOR2X1_LOC_48/B 0.07fF
C70723 NOR2X1_LOC_67/A NAND2X1_LOC_74/B 0.15fF
C70724 INVX1_LOC_58/A NAND2X1_LOC_355/a_36_24# 0.01fF
C70725 NOR2X1_LOC_74/A NOR2X1_LOC_536/A 0.14fF
C70726 NAND2X1_LOC_656/Y NOR2X1_LOC_473/a_36_216# 0.01fF
C70727 INVX1_LOC_6/A INVX1_LOC_37/Y 0.00fF
C70728 INVX1_LOC_21/A INVX1_LOC_14/A 0.07fF
C70729 D_INPUT_1 INVX1_LOC_223/A 0.72fF
C70730 INVX1_LOC_55/Y INVX1_LOC_179/A 0.03fF
C70731 NOR2X1_LOC_405/A INVX1_LOC_76/A 0.10fF
C70732 INVX1_LOC_25/Y NAND2X1_LOC_81/B 0.03fF
C70733 INVX1_LOC_276/Y INVX1_LOC_42/A 0.02fF
C70734 NOR2X1_LOC_68/A NOR2X1_LOC_654/A 0.01fF
C70735 INVX1_LOC_256/A INVX1_LOC_306/Y 0.01fF
C70736 INVX1_LOC_282/A INVX1_LOC_118/A 0.03fF
C70737 NAND2X1_LOC_819/Y NOR2X1_LOC_847/A 0.12fF
C70738 NOR2X1_LOC_9/Y NOR2X1_LOC_536/A 0.17fF
C70739 NAND2X1_LOC_361/Y INVX1_LOC_87/A 0.07fF
C70740 NAND2X1_LOC_214/B NOR2X1_LOC_160/B 0.07fF
C70741 INVX1_LOC_268/A INVX1_LOC_29/A 0.05fF
C70742 NOR2X1_LOC_150/a_36_216# INVX1_LOC_285/A 0.00fF
C70743 INVX1_LOC_15/Y INVX1_LOC_3/Y 0.01fF
C70744 NOR2X1_LOC_657/B NAND2X1_LOC_211/Y 0.07fF
C70745 NAND2X1_LOC_354/B INVX1_LOC_78/A 0.00fF
C70746 NOR2X1_LOC_488/Y INVX1_LOC_42/A 0.33fF
C70747 INVX1_LOC_91/A NOR2X1_LOC_60/Y 0.04fF
C70748 INVX1_LOC_196/Y NOR2X1_LOC_801/A 0.01fF
C70749 INVX1_LOC_33/A INVX1_LOC_26/A 0.07fF
C70750 NOR2X1_LOC_785/a_36_216# NOR2X1_LOC_634/A 0.00fF
C70751 NOR2X1_LOC_824/A NAND2X1_LOC_550/A 0.05fF
C70752 NAND2X1_LOC_866/B NOR2X1_LOC_485/Y 0.01fF
C70753 NOR2X1_LOC_68/A INVX1_LOC_58/Y 0.05fF
C70754 INVX1_LOC_27/A NOR2X1_LOC_160/B 0.32fF
C70755 NOR2X1_LOC_74/A NAND2X1_LOC_93/B 0.07fF
C70756 NOR2X1_LOC_665/A NOR2X1_LOC_755/Y 0.06fF
C70757 NOR2X1_LOC_334/A NOR2X1_LOC_729/A 0.03fF
C70758 INVX1_LOC_228/Y INVX1_LOC_1/A 0.01fF
C70759 NOR2X1_LOC_253/Y INVX1_LOC_46/A 0.01fF
C70760 INVX1_LOC_266/A NOR2X1_LOC_457/A 0.10fF
C70761 NAND2X1_LOC_192/B INVX1_LOC_88/A 0.02fF
C70762 D_INPUT_3 INVX1_LOC_20/A 0.03fF
C70763 NOR2X1_LOC_433/A INVX1_LOC_57/A 0.06fF
C70764 NOR2X1_LOC_708/A INVX1_LOC_117/A 0.01fF
C70765 INVX1_LOC_30/A INVX1_LOC_50/Y 0.03fF
C70766 NOR2X1_LOC_561/Y INVX1_LOC_109/Y 0.03fF
C70767 NOR2X1_LOC_9/Y NAND2X1_LOC_93/B 0.07fF
C70768 NOR2X1_LOC_188/A NOR2X1_LOC_445/B 0.55fF
C70769 INVX1_LOC_227/A INVX1_LOC_42/A 0.07fF
C70770 INVX1_LOC_103/A NOR2X1_LOC_218/A 0.01fF
C70771 NOR2X1_LOC_687/Y INVX1_LOC_15/A 0.08fF
C70772 NAND2X1_LOC_363/B NOR2X1_LOC_559/B 0.03fF
C70773 NOR2X1_LOC_709/A INVX1_LOC_23/Y 0.17fF
C70774 NOR2X1_LOC_548/B NOR2X1_LOC_445/B 0.01fF
C70775 NOR2X1_LOC_772/B NAND2X1_LOC_656/A 0.14fF
C70776 INVX1_LOC_5/A NOR2X1_LOC_215/Y 0.05fF
C70777 INVX1_LOC_286/Y NOR2X1_LOC_536/Y 0.07fF
C70778 NOR2X1_LOC_174/A NOR2X1_LOC_633/A 0.00fF
C70779 NOR2X1_LOC_488/Y INVX1_LOC_78/A 0.03fF
C70780 INVX1_LOC_13/Y NAND2X1_LOC_656/A 0.01fF
C70781 INVX1_LOC_27/A NOR2X1_LOC_733/a_36_216# 0.01fF
C70782 NOR2X1_LOC_510/Y NOR2X1_LOC_351/a_36_216# 0.01fF
C70783 NOR2X1_LOC_52/B INVX1_LOC_57/A 0.35fF
C70784 INVX1_LOC_158/Y NOR2X1_LOC_814/A 0.03fF
C70785 NOR2X1_LOC_572/a_36_216# NOR2X1_LOC_38/B 0.00fF
C70786 NOR2X1_LOC_388/Y NOR2X1_LOC_717/A 0.10fF
C70787 NOR2X1_LOC_82/Y INVX1_LOC_78/A 0.02fF
C70788 NOR2X1_LOC_360/A INVX1_LOC_230/A 0.02fF
C70789 NAND2X1_LOC_451/Y NOR2X1_LOC_635/B 0.12fF
C70790 INVX1_LOC_40/A INVX1_LOC_26/A 0.04fF
C70791 NAND2X1_LOC_338/B NAND2X1_LOC_96/a_36_24# 0.01fF
C70792 INVX1_LOC_24/A D_INPUT_6 0.01fF
C70793 INVX1_LOC_190/A INVX1_LOC_15/A 0.01fF
C70794 NOR2X1_LOC_361/Y INVX1_LOC_23/A 0.15fF
C70795 INVX1_LOC_286/Y NAND2X1_LOC_799/A 0.04fF
C70796 INVX1_LOC_165/Y INVX1_LOC_26/A 0.01fF
C70797 NOR2X1_LOC_624/A INVX1_LOC_64/A 0.10fF
C70798 INVX1_LOC_58/A INVX1_LOC_96/Y 0.10fF
C70799 INVX1_LOC_89/A D_INPUT_5 0.09fF
C70800 NAND2X1_LOC_363/B NOR2X1_LOC_6/B 0.13fF
C70801 NOR2X1_LOC_510/Y NOR2X1_LOC_577/Y 0.00fF
C70802 INVX1_LOC_24/A NOR2X1_LOC_321/Y 0.07fF
C70803 INVX1_LOC_256/A NOR2X1_LOC_657/Y 0.04fF
C70804 INVX1_LOC_278/A INVX1_LOC_124/A 0.16fF
C70805 INVX1_LOC_92/Y INVX1_LOC_19/A 0.02fF
C70806 NAND2X1_LOC_44/a_36_24# INVX1_LOC_11/A 0.00fF
C70807 NOR2X1_LOC_717/B NAND2X1_LOC_454/Y 0.06fF
C70808 NOR2X1_LOC_88/Y NOR2X1_LOC_670/a_36_216# 0.00fF
C70809 NOR2X1_LOC_19/B NOR2X1_LOC_554/A 0.01fF
C70810 INVX1_LOC_64/A NOR2X1_LOC_93/a_36_216# 0.00fF
C70811 NOR2X1_LOC_844/Y NOR2X1_LOC_590/A 0.01fF
C70812 INVX1_LOC_5/A INVX1_LOC_104/A 0.07fF
C70813 INVX1_LOC_159/A NAND2X1_LOC_154/a_36_24# 0.00fF
C70814 NOR2X1_LOC_500/A INVX1_LOC_269/A 0.85fF
C70815 INVX1_LOC_50/A INVX1_LOC_1/Y 0.03fF
C70816 INVX1_LOC_162/Y NOR2X1_LOC_652/Y 0.00fF
C70817 NOR2X1_LOC_75/Y NOR2X1_LOC_68/A 0.03fF
C70818 INVX1_LOC_269/A NOR2X1_LOC_303/Y 0.10fF
C70819 NOR2X1_LOC_431/Y INVX1_LOC_103/A 0.04fF
C70820 INVX1_LOC_130/A INVX1_LOC_36/A 0.02fF
C70821 NOR2X1_LOC_474/A NOR2X1_LOC_475/A 0.00fF
C70822 NOR2X1_LOC_369/Y INVX1_LOC_18/A 0.06fF
C70823 INVX1_LOC_35/A NOR2X1_LOC_544/A 0.49fF
C70824 NAND2X1_LOC_783/Y NOR2X1_LOC_68/A 0.07fF
C70825 NOR2X1_LOC_666/A INVX1_LOC_33/A 0.13fF
C70826 NOR2X1_LOC_562/B INVX1_LOC_19/A 0.03fF
C70827 NOR2X1_LOC_361/B NOR2X1_LOC_577/Y 0.04fF
C70828 NAND2X1_LOC_9/Y INVX1_LOC_16/A 0.06fF
C70829 NAND2X1_LOC_848/A INVX1_LOC_185/A 0.01fF
C70830 INVX1_LOC_101/A INVX1_LOC_23/A 0.01fF
C70831 INVX1_LOC_12/Y NOR2X1_LOC_216/B 0.11fF
C70832 INVX1_LOC_286/Y INVX1_LOC_18/A 0.07fF
C70833 NOR2X1_LOC_557/A NAND2X1_LOC_207/B 0.06fF
C70834 INVX1_LOC_290/A INVX1_LOC_53/A 0.07fF
C70835 NOR2X1_LOC_637/a_36_216# INVX1_LOC_103/A 0.00fF
C70836 NOR2X1_LOC_246/A NAND2X1_LOC_288/B 0.87fF
C70837 NOR2X1_LOC_231/a_36_216# NOR2X1_LOC_68/A 0.01fF
C70838 INVX1_LOC_90/A NAND2X1_LOC_616/a_36_24# 0.00fF
C70839 NAND2X1_LOC_803/B NOR2X1_LOC_152/Y 0.02fF
C70840 INVX1_LOC_233/A INVX1_LOC_16/A 0.01fF
C70841 NAND2X1_LOC_729/Y NAND2X1_LOC_733/Y 0.05fF
C70842 NAND2X1_LOC_728/Y INVX1_LOC_286/Y 0.07fF
C70843 INVX1_LOC_21/A INVX1_LOC_111/Y 0.02fF
C70844 INVX1_LOC_269/A NOR2X1_LOC_84/A 0.23fF
C70845 INVX1_LOC_289/Y NAND2X1_LOC_799/Y 0.11fF
C70846 INVX1_LOC_75/A INVX1_LOC_4/Y 0.27fF
C70847 INVX1_LOC_36/A NOR2X1_LOC_791/B 1.72fF
C70848 NAND2X1_LOC_363/B INVX1_LOC_30/Y 0.03fF
C70849 NOR2X1_LOC_43/Y INVX1_LOC_12/A 0.01fF
C70850 NOR2X1_LOC_598/B INVX1_LOC_279/A 0.20fF
C70851 INVX1_LOC_64/A NAND2X1_LOC_735/B 0.80fF
C70852 INVX1_LOC_217/A NOR2X1_LOC_384/Y 0.03fF
C70853 NOR2X1_LOC_315/Y NOR2X1_LOC_271/B 0.02fF
C70854 NOR2X1_LOC_151/Y NAND2X1_LOC_454/Y 0.05fF
C70855 NOR2X1_LOC_355/A INVX1_LOC_23/A 0.09fF
C70856 NOR2X1_LOC_590/A NOR2X1_LOC_152/Y 0.07fF
C70857 VDD NAND2X1_LOC_476/Y 0.04fF
C70858 INVX1_LOC_95/Y INVX1_LOC_29/A 0.01fF
C70859 NAND2X1_LOC_214/B NOR2X1_LOC_516/B 0.33fF
C70860 NOR2X1_LOC_632/Y NOR2X1_LOC_665/Y 0.01fF
C70861 NOR2X1_LOC_824/A NAND2X1_LOC_500/a_36_24# 0.01fF
C70862 NAND2X1_LOC_553/A INVX1_LOC_16/A 0.00fF
C70863 NOR2X1_LOC_226/A NOR2X1_LOC_440/B 0.03fF
C70864 INVX1_LOC_24/Y NOR2X1_LOC_175/A 0.03fF
C70865 INVX1_LOC_97/Y INVX1_LOC_279/A -0.01fF
C70866 INVX1_LOC_38/A INVX1_LOC_260/Y 0.03fF
C70867 NOR2X1_LOC_349/B NOR2X1_LOC_342/A 0.00fF
C70868 NAND2X1_LOC_624/B NAND2X1_LOC_462/B 0.00fF
C70869 VDD INVX1_LOC_186/Y 0.28fF
C70870 INVX1_LOC_159/A INVX1_LOC_18/A 0.17fF
C70871 NAND2X1_LOC_500/Y NOR2X1_LOC_495/Y 0.01fF
C70872 NOR2X1_LOC_78/B INVX1_LOC_48/Y 0.07fF
C70873 INVX1_LOC_27/A INVX1_LOC_208/A 0.48fF
C70874 NOR2X1_LOC_510/Y INVX1_LOC_22/A 0.07fF
C70875 INVX1_LOC_292/A INVX1_LOC_155/Y 0.01fF
C70876 NOR2X1_LOC_567/B NOR2X1_LOC_798/Y 0.06fF
C70877 NOR2X1_LOC_798/A INVX1_LOC_16/A 0.00fF
C70878 NOR2X1_LOC_397/a_36_216# INVX1_LOC_306/Y 0.01fF
C70879 INVX1_LOC_36/A INVX1_LOC_81/A 0.03fF
C70880 INVX1_LOC_269/A INVX1_LOC_54/Y 0.01fF
C70881 INVX1_LOC_1/A NAND2X1_LOC_832/a_36_24# 0.00fF
C70882 NOR2X1_LOC_331/B NOR2X1_LOC_697/Y 0.05fF
C70883 INVX1_LOC_27/A NOR2X1_LOC_516/B 0.09fF
C70884 NAND2X1_LOC_53/Y NOR2X1_LOC_300/Y 0.00fF
C70885 NAND2X1_LOC_715/B INVX1_LOC_279/A 0.03fF
C70886 NOR2X1_LOC_607/Y INVX1_LOC_223/A 0.01fF
C70887 NOR2X1_LOC_824/A NAND2X1_LOC_705/a_36_24# 0.01fF
C70888 NAND2X1_LOC_337/B INVX1_LOC_104/A 0.10fF
C70889 NOR2X1_LOC_191/B INVX1_LOC_18/A 1.01fF
C70890 VDD NOR2X1_LOC_777/B 0.61fF
C70891 NOR2X1_LOC_68/A NAND2X1_LOC_162/B 0.02fF
C70892 NAND2X1_LOC_434/Y NAND2X1_LOC_798/B 0.15fF
C70893 NOR2X1_LOC_667/A INVX1_LOC_14/A 0.01fF
C70894 INVX1_LOC_103/A NOR2X1_LOC_131/A 0.02fF
C70895 VDD INVX1_LOC_261/A 0.00fF
C70896 INVX1_LOC_1/A NOR2X1_LOC_566/Y 0.03fF
C70897 INVX1_LOC_109/A INVX1_LOC_46/A 0.01fF
C70898 INVX1_LOC_49/A INVX1_LOC_142/A 0.03fF
C70899 INVX1_LOC_109/Y INVX1_LOC_76/A 0.01fF
C70900 NOR2X1_LOC_567/B NOR2X1_LOC_748/A 0.10fF
C70901 INVX1_LOC_136/A NOR2X1_LOC_753/Y 4.38fF
C70902 D_INPUT_3 NOR2X1_LOC_128/A 0.01fF
C70903 NOR2X1_LOC_468/Y INVX1_LOC_56/A 0.02fF
C70904 INVX1_LOC_84/A INVX1_LOC_9/A 0.07fF
C70905 NOR2X1_LOC_68/A NOR2X1_LOC_419/Y 0.03fF
C70906 NOR2X1_LOC_384/Y NAND2X1_LOC_787/B 0.16fF
C70907 NOR2X1_LOC_140/A INVX1_LOC_232/A 0.00fF
C70908 NAND2X1_LOC_9/Y INVX1_LOC_28/A 0.11fF
C70909 NOR2X1_LOC_92/Y NAND2X1_LOC_848/a_36_24# 0.01fF
C70910 NAND2X1_LOC_650/B INVX1_LOC_42/A 0.07fF
C70911 NAND2X1_LOC_41/Y NAND2X1_LOC_473/A 0.02fF
C70912 NOR2X1_LOC_441/Y NAND2X1_LOC_357/B 0.07fF
C70913 INVX1_LOC_92/Y INVX1_LOC_26/Y 0.03fF
C70914 NOR2X1_LOC_276/Y INVX1_LOC_133/Y 0.01fF
C70915 INVX1_LOC_233/A INVX1_LOC_28/A 0.07fF
C70916 NOR2X1_LOC_68/A NOR2X1_LOC_716/B 0.08fF
C70917 NAND2X1_LOC_374/a_36_24# INVX1_LOC_24/A 0.00fF
C70918 NOR2X1_LOC_269/a_36_216# INVX1_LOC_88/A 0.00fF
C70919 INVX1_LOC_45/A NOR2X1_LOC_799/a_36_216# 0.00fF
C70920 NOR2X1_LOC_6/B INVX1_LOC_30/A 0.03fF
C70921 NOR2X1_LOC_361/B INVX1_LOC_22/A 0.00fF
C70922 NOR2X1_LOC_276/B INVX1_LOC_33/A 0.02fF
C70923 NOR2X1_LOC_799/a_36_216# NOR2X1_LOC_568/A 0.00fF
C70924 NOR2X1_LOC_789/B NOR2X1_LOC_99/B 0.03fF
C70925 INVX1_LOC_27/A NAND2X1_LOC_133/a_36_24# 0.00fF
C70926 INVX1_LOC_21/A NOR2X1_LOC_137/A 0.03fF
C70927 NAND2X1_LOC_649/a_36_24# INVX1_LOC_15/A 0.01fF
C70928 NOR2X1_LOC_592/B NOR2X1_LOC_697/Y 0.66fF
C70929 INVX1_LOC_289/Y NAND2X1_LOC_319/A 0.27fF
C70930 INVX1_LOC_265/A NOR2X1_LOC_91/Y 0.22fF
C70931 NOR2X1_LOC_321/Y NOR2X1_LOC_130/A 0.07fF
C70932 NOR2X1_LOC_552/Y INVX1_LOC_23/A 0.01fF
C70933 NOR2X1_LOC_487/a_36_216# NOR2X1_LOC_315/Y 0.00fF
C70934 INVX1_LOC_6/A INVX1_LOC_29/Y 0.05fF
C70935 INVX1_LOC_58/A NOR2X1_LOC_733/Y 0.03fF
C70936 D_INPUT_3 INVX1_LOC_4/A 0.28fF
C70937 NAND2X1_LOC_21/Y INVX1_LOC_77/A 0.56fF
C70938 INVX1_LOC_232/Y NOR2X1_LOC_382/Y 0.02fF
C70939 INVX1_LOC_14/Y INVX1_LOC_4/A 0.10fF
C70940 NOR2X1_LOC_82/A NOR2X1_LOC_789/a_36_216# 0.00fF
C70941 NOR2X1_LOC_160/B INVX1_LOC_137/A 0.03fF
C70942 NOR2X1_LOC_590/Y NOR2X1_LOC_742/A 0.04fF
C70943 INVX1_LOC_50/A NOR2X1_LOC_318/B 0.03fF
C70944 NOR2X1_LOC_264/Y INVX1_LOC_314/Y 0.11fF
C70945 NOR2X1_LOC_457/B INVX1_LOC_266/Y 0.10fF
C70946 NAND2X1_LOC_354/B NOR2X1_LOC_152/Y 0.07fF
C70947 NOR2X1_LOC_396/Y NAND2X1_LOC_402/B 0.06fF
C70948 NOR2X1_LOC_67/A INVX1_LOC_136/A 0.15fF
C70949 NAND2X1_LOC_650/B INVX1_LOC_78/A 0.07fF
C70950 NAND2X1_LOC_854/B NOR2X1_LOC_816/A 0.15fF
C70951 NAND2X1_LOC_703/Y INVX1_LOC_28/A 0.39fF
C70952 NAND2X1_LOC_819/Y NOR2X1_LOC_554/B 0.03fF
C70953 NOR2X1_LOC_130/A NAND2X1_LOC_793/Y 0.03fF
C70954 INVX1_LOC_2/A INVX1_LOC_41/Y 0.03fF
C70955 NOR2X1_LOC_778/B NOR2X1_LOC_598/a_36_216# 0.00fF
C70956 INVX1_LOC_261/Y INVX1_LOC_92/A 0.03fF
C70957 INVX1_LOC_150/Y INVX1_LOC_66/A -0.02fF
C70958 NOR2X1_LOC_658/Y NAND2X1_LOC_479/Y 0.07fF
C70959 NOR2X1_LOC_219/Y INVX1_LOC_72/A 0.07fF
C70960 INVX1_LOC_223/A NOR2X1_LOC_553/Y 0.01fF
C70961 INVX1_LOC_160/A INVX1_LOC_53/A 0.43fF
C70962 NOR2X1_LOC_91/A INVX1_LOC_126/A 0.01fF
C70963 INVX1_LOC_125/A NAND2X1_LOC_750/a_36_24# 0.00fF
C70964 NOR2X1_LOC_191/B NOR2X1_LOC_709/a_36_216# 0.01fF
C70965 NOR2X1_LOC_820/A INVX1_LOC_40/A 0.01fF
C70966 INVX1_LOC_114/Y INVX1_LOC_92/A 0.01fF
C70967 INVX1_LOC_57/Y NAND2X1_LOC_564/B 0.10fF
C70968 INVX1_LOC_72/A INVX1_LOC_53/Y -0.01fF
C70969 INVX1_LOC_30/Y INVX1_LOC_30/A 0.02fF
C70970 INVX1_LOC_64/A NOR2X1_LOC_7/Y 0.04fF
C70971 NOR2X1_LOC_226/A INVX1_LOC_41/Y 0.03fF
C70972 INVX1_LOC_9/A INVX1_LOC_15/A 1.54fF
C70973 INVX1_LOC_5/A INVX1_LOC_206/Y 0.07fF
C70974 INVX1_LOC_2/A NAND2X1_LOC_593/Y 0.38fF
C70975 NAND2X1_LOC_717/Y NAND2X1_LOC_866/A 2.08fF
C70976 NAND2X1_LOC_733/B NAND2X1_LOC_863/Y 0.28fF
C70977 INVX1_LOC_74/A INVX1_LOC_57/A 0.03fF
C70978 NOR2X1_LOC_577/Y INVX1_LOC_177/A 0.03fF
C70979 NOR2X1_LOC_473/B INVX1_LOC_161/Y 0.10fF
C70980 INVX1_LOC_88/A NOR2X1_LOC_329/B 0.01fF
C70981 INVX1_LOC_153/Y NOR2X1_LOC_348/B 0.00fF
C70982 INVX1_LOC_276/Y NOR2X1_LOC_152/Y 0.03fF
C70983 NAND2X1_LOC_72/Y NOR2X1_LOC_318/B -0.03fF
C70984 INVX1_LOC_305/A NOR2X1_LOC_748/Y 0.01fF
C70985 VDD NOR2X1_LOC_843/B 0.17fF
C70986 NOR2X1_LOC_226/A NAND2X1_LOC_593/Y 0.03fF
C70987 NOR2X1_LOC_180/B INVX1_LOC_225/Y 0.13fF
C70988 NOR2X1_LOC_862/B NOR2X1_LOC_640/B 0.05fF
C70989 NOR2X1_LOC_186/Y NOR2X1_LOC_114/A 0.04fF
C70990 NOR2X1_LOC_91/A NOR2X1_LOC_111/A 0.10fF
C70991 NAND2X1_LOC_214/B INVX1_LOC_315/Y 0.11fF
C70992 INVX1_LOC_50/A INVX1_LOC_139/A 0.00fF
C70993 NOR2X1_LOC_74/A NOR2X1_LOC_348/Y 0.73fF
C70994 NOR2X1_LOC_419/Y NOR2X1_LOC_520/a_36_216# 0.00fF
C70995 INVX1_LOC_230/Y INVX1_LOC_90/A 0.60fF
C70996 INVX1_LOC_21/A INVX1_LOC_48/A 0.03fF
C70997 NOR2X1_LOC_781/B INVX1_LOC_72/A 0.15fF
C70998 INVX1_LOC_249/A INVX1_LOC_208/A 0.04fF
C70999 INVX1_LOC_271/A NAND2X1_LOC_211/Y 0.03fF
C71000 NOR2X1_LOC_205/Y INVX1_LOC_75/A 0.15fF
C71001 NAND2X1_LOC_555/Y INVX1_LOC_20/Y 0.05fF
C71002 NOR2X1_LOC_470/A NOR2X1_LOC_68/A 0.10fF
C71003 INVX1_LOC_35/A NAND2X1_LOC_468/B 0.03fF
C71004 NOR2X1_LOC_467/A INVX1_LOC_92/A 0.28fF
C71005 INVX1_LOC_32/A INVX1_LOC_179/A 0.03fF
C71006 NAND2X1_LOC_9/Y NOR2X1_LOC_35/Y 0.10fF
C71007 NOR2X1_LOC_769/A NOR2X1_LOC_763/Y 0.18fF
C71008 NOR2X1_LOC_186/Y INVX1_LOC_91/A 0.22fF
C71009 INVX1_LOC_2/Y NOR2X1_LOC_416/A 0.58fF
C71010 INVX1_LOC_50/A NAND2X1_LOC_721/A 0.05fF
C71011 NOR2X1_LOC_468/Y NOR2X1_LOC_83/Y 0.05fF
C71012 NOR2X1_LOC_514/A INPUT_1 0.17fF
C71013 NOR2X1_LOC_424/Y NOR2X1_LOC_68/A 0.11fF
C71014 NOR2X1_LOC_160/B NOR2X1_LOC_19/B 0.04fF
C71015 INVX1_LOC_64/A NAND2X1_LOC_212/Y 0.00fF
C71016 INVX1_LOC_177/A NOR2X1_LOC_348/B 0.00fF
C71017 INVX1_LOC_225/A NOR2X1_LOC_279/a_36_216# 0.00fF
C71018 NOR2X1_LOC_363/Y INVX1_LOC_270/A 0.10fF
C71019 NAND2X1_LOC_323/B INVX1_LOC_310/Y 0.19fF
C71020 INVX1_LOC_1/A NAND2X1_LOC_841/a_36_24# 0.00fF
C71021 NOR2X1_LOC_309/Y NOR2X1_LOC_767/a_36_216# 0.00fF
C71022 NAND2X1_LOC_347/B INVX1_LOC_286/A 0.02fF
C71023 NOR2X1_LOC_717/B NOR2X1_LOC_68/A 0.01fF
C71024 NOR2X1_LOC_589/A NOR2X1_LOC_106/Y 0.28fF
C71025 NOR2X1_LOC_361/B INVX1_LOC_100/A 0.05fF
C71026 INVX1_LOC_80/Y INVX1_LOC_216/A 0.01fF
C71027 NOR2X1_LOC_795/Y NOR2X1_LOC_168/B 0.05fF
C71028 NOR2X1_LOC_328/Y INVX1_LOC_209/Y 0.06fF
C71029 INVX1_LOC_256/A NOR2X1_LOC_74/A 0.10fF
C71030 INVX1_LOC_24/A NOR2X1_LOC_686/B 0.02fF
C71031 INVX1_LOC_269/A NOR2X1_LOC_354/Y 0.03fF
C71032 INVX1_LOC_40/A INVX1_LOC_315/A 0.23fF
C71033 NAND2X1_LOC_795/a_36_24# NAND2X1_LOC_722/A 0.00fF
C71034 INVX1_LOC_37/A NAND2X1_LOC_793/B 0.07fF
C71035 NAND2X1_LOC_254/Y NOR2X1_LOC_662/A 0.01fF
C71036 NOR2X1_LOC_791/Y NOR2X1_LOC_124/A 0.02fF
C71037 NOR2X1_LOC_617/Y NAND2X1_LOC_462/B 0.00fF
C71038 NOR2X1_LOC_637/A NOR2X1_LOC_130/A 0.00fF
C71039 INVX1_LOC_230/Y NAND2X1_LOC_348/A 0.02fF
C71040 INVX1_LOC_89/A NOR2X1_LOC_360/Y 0.10fF
C71041 INVX1_LOC_64/A D_INPUT_3 0.11fF
C71042 NOR2X1_LOC_773/Y INVX1_LOC_104/A 0.14fF
C71043 NAND2X1_LOC_9/Y NOR2X1_LOC_133/a_36_216# 0.00fF
C71044 INVX1_LOC_153/Y INVX1_LOC_22/A 0.47fF
C71045 INVX1_LOC_64/A INVX1_LOC_14/Y 0.10fF
C71046 NOR2X1_LOC_68/A NOR2X1_LOC_130/Y 0.01fF
C71047 NAND2X1_LOC_794/B NOR2X1_LOC_164/Y 0.01fF
C71048 NOR2X1_LOC_449/a_36_216# NOR2X1_LOC_130/A 0.00fF
C71049 INVX1_LOC_256/A NOR2X1_LOC_9/Y 0.16fF
C71050 NOR2X1_LOC_664/Y NOR2X1_LOC_516/B 0.12fF
C71051 NAND2X1_LOC_724/A INVX1_LOC_91/A 0.44fF
C71052 NOR2X1_LOC_658/Y NOR2X1_LOC_202/Y 0.02fF
C71053 NAND2X1_LOC_740/Y INVX1_LOC_76/A 0.07fF
C71054 NOR2X1_LOC_798/A NOR2X1_LOC_35/Y 0.05fF
C71055 NOR2X1_LOC_434/Y NOR2X1_LOC_857/A 0.03fF
C71056 NOR2X1_LOC_99/Y NAND2X1_LOC_99/A 0.07fF
C71057 INVX1_LOC_10/Y NOR2X1_LOC_717/A 0.00fF
C71058 NAND2X1_LOC_456/a_36_24# INVX1_LOC_19/A 0.01fF
C71059 INVX1_LOC_41/Y INPUT_1 0.03fF
C71060 INVX1_LOC_206/A INVX1_LOC_208/A 0.01fF
C71061 NOR2X1_LOC_614/Y NOR2X1_LOC_168/B 0.00fF
C71062 INVX1_LOC_57/A NOR2X1_LOC_675/a_36_216# 0.00fF
C71063 NOR2X1_LOC_440/Y INVX1_LOC_294/Y 0.00fF
C71064 NAND2X1_LOC_162/B NOR2X1_LOC_163/A 0.11fF
C71065 NOR2X1_LOC_194/Y NOR2X1_LOC_589/A 0.04fF
C71066 NOR2X1_LOC_175/A NOR2X1_LOC_211/A 0.04fF
C71067 NAND2X1_LOC_724/A INVX1_LOC_11/Y 0.07fF
C71068 NAND2X1_LOC_794/B INVX1_LOC_46/A 0.00fF
C71069 INVX1_LOC_23/A INVX1_LOC_127/A 0.01fF
C71070 INVX1_LOC_27/A NAND2X1_LOC_211/Y 0.01fF
C71071 NAND2X1_LOC_425/a_36_24# NAND2X1_LOC_425/Y 0.00fF
C71072 INVX1_LOC_177/A INVX1_LOC_22/A 0.07fF
C71073 INVX1_LOC_14/A INVX1_LOC_304/A 0.07fF
C71074 NAND2X1_LOC_550/A NOR2X1_LOC_528/Y 0.04fF
C71075 INVX1_LOC_135/A NAND2X1_LOC_175/B 0.06fF
C71076 INVX1_LOC_108/Y INVX1_LOC_9/A 0.08fF
C71077 NAND2X1_LOC_401/a_36_24# INVX1_LOC_241/Y 0.01fF
C71078 NOR2X1_LOC_717/Y INVX1_LOC_311/A 1.09fF
C71079 NAND2X1_LOC_705/Y INVX1_LOC_20/A 0.00fF
C71080 NOR2X1_LOC_67/Y INVX1_LOC_42/A 0.09fF
C71081 NOR2X1_LOC_68/A NOR2X1_LOC_151/Y 0.09fF
C71082 NAND2X1_LOC_454/Y NOR2X1_LOC_666/a_36_216# 0.01fF
C71083 NAND2X1_LOC_175/Y INVX1_LOC_250/Y 0.09fF
C71084 NOR2X1_LOC_79/A INVX1_LOC_29/Y 0.02fF
C71085 NOR2X1_LOC_781/A INVX1_LOC_266/Y 0.00fF
C71086 NOR2X1_LOC_619/A NAND2X1_LOC_338/B 0.02fF
C71087 NAND2X1_LOC_303/Y INVX1_LOC_20/A 0.06fF
C71088 NOR2X1_LOC_113/B INVX1_LOC_72/A 0.03fF
C71089 NOR2X1_LOC_457/B INVX1_LOC_42/Y 0.01fF
C71090 NOR2X1_LOC_78/B NOR2X1_LOC_374/B 0.02fF
C71091 INVX1_LOC_280/Y INVX1_LOC_22/A 0.08fF
C71092 INVX1_LOC_16/A NOR2X1_LOC_505/Y 0.05fF
C71093 NAND2X1_LOC_231/Y NAND2X1_LOC_390/A 0.19fF
C71094 NAND2X1_LOC_477/Y NOR2X1_LOC_89/Y 0.01fF
C71095 NOR2X1_LOC_78/B INVX1_LOC_290/A 0.02fF
C71096 NOR2X1_LOC_226/A NAND2X1_LOC_861/a_36_24# 0.01fF
C71097 NAND2X1_LOC_624/B INVX1_LOC_118/A 0.01fF
C71098 NOR2X1_LOC_177/Y NAND2X1_LOC_793/B 0.27fF
C71099 NOR2X1_LOC_672/a_36_216# INVX1_LOC_3/Y 0.01fF
C71100 INVX1_LOC_47/A INVX1_LOC_8/A 0.01fF
C71101 INVX1_LOC_141/Y NOR2X1_LOC_45/B 0.03fF
C71102 NOR2X1_LOC_536/Y VDD 0.25fF
C71103 INVX1_LOC_136/A NAND2X1_LOC_103/a_36_24# 0.01fF
C71104 NOR2X1_LOC_186/Y NAND2X1_LOC_783/a_36_24# 0.00fF
C71105 NAND2X1_LOC_123/Y INVX1_LOC_155/A 0.02fF
C71106 NOR2X1_LOC_536/Y NAND2X1_LOC_800/A 0.01fF
C71107 NOR2X1_LOC_693/Y NAND2X1_LOC_489/Y 0.00fF
C71108 NAND2X1_LOC_717/Y NOR2X1_LOC_700/Y 0.03fF
C71109 INVX1_LOC_312/Y NOR2X1_LOC_45/B 0.72fF
C71110 NOR2X1_LOC_861/Y INVX1_LOC_15/A 0.29fF
C71111 INVX1_LOC_182/A NOR2X1_LOC_344/A 0.02fF
C71112 INVX1_LOC_77/A NOR2X1_LOC_310/a_36_216# 0.00fF
C71113 INVX1_LOC_36/A NOR2X1_LOC_192/A 0.01fF
C71114 NAND2X1_LOC_799/A VDD 0.21fF
C71115 NAND2X1_LOC_303/Y NOR2X1_LOC_765/Y 0.09fF
C71116 NAND2X1_LOC_59/B D_INPUT_4 0.51fF
C71117 INVX1_LOC_255/Y INVX1_LOC_13/A 0.30fF
C71118 INVX1_LOC_277/A NOR2X1_LOC_711/Y 0.16fF
C71119 NAND2X1_LOC_799/A NAND2X1_LOC_800/A 0.17fF
C71120 INVX1_LOC_89/A NAND2X1_LOC_451/Y 0.12fF
C71121 NOR2X1_LOC_620/Y INPUT_0 0.35fF
C71122 INVX1_LOC_58/A NAND2X1_LOC_456/Y 0.26fF
C71123 INVX1_LOC_35/A NAND2X1_LOC_141/Y 0.52fF
C71124 INVX1_LOC_62/Y NOR2X1_LOC_845/A 0.00fF
C71125 INVX1_LOC_45/A NOR2X1_LOC_631/B 0.05fF
C71126 INVX1_LOC_285/Y NOR2X1_LOC_577/Y 0.10fF
C71127 INVX1_LOC_94/A NAND2X1_LOC_498/a_36_24# 0.00fF
C71128 INVX1_LOC_106/A INVX1_LOC_26/Y 0.01fF
C71129 INVX1_LOC_75/A INVX1_LOC_82/A 0.04fF
C71130 NOR2X1_LOC_488/a_36_216# NAND2X1_LOC_862/Y 0.01fF
C71131 NOR2X1_LOC_488/Y NAND2X1_LOC_861/Y 0.09fF
C71132 INVX1_LOC_77/A INVX1_LOC_123/A 0.02fF
C71133 NAND2X1_LOC_662/B INVX1_LOC_63/Y 0.01fF
C71134 INVX1_LOC_83/A NOR2X1_LOC_374/B 0.04fF
C71135 INVX1_LOC_274/Y INVX1_LOC_15/A 0.22fF
C71136 NOR2X1_LOC_250/Y NOR2X1_LOC_536/A 0.21fF
C71137 INVX1_LOC_143/A INVX1_LOC_148/A 0.02fF
C71138 INVX1_LOC_290/A INVX1_LOC_83/A 0.10fF
C71139 INVX1_LOC_18/A NOR2X1_LOC_56/Y 0.07fF
C71140 NOR2X1_LOC_68/A NOR2X1_LOC_181/A 0.02fF
C71141 NOR2X1_LOC_292/Y NOR2X1_LOC_392/B 0.01fF
C71142 NAND2X1_LOC_149/Y NOR2X1_LOC_156/a_36_216# 0.01fF
C71143 NAND2X1_LOC_63/Y INVX1_LOC_129/A 0.00fF
C71144 INVX1_LOC_36/A INVX1_LOC_2/Y 0.04fF
C71145 NAND2X1_LOC_721/B NOR2X1_LOC_305/Y -0.02fF
C71146 NOR2X1_LOC_186/Y NAND2X1_LOC_273/a_36_24# 0.00fF
C71147 INVX1_LOC_72/A NOR2X1_LOC_585/Y 0.04fF
C71148 INVX1_LOC_132/A INVX1_LOC_91/A 0.07fF
C71149 INVX1_LOC_45/A INVX1_LOC_37/A 6.86fF
C71150 NOR2X1_LOC_274/Y NOR2X1_LOC_405/A 0.01fF
C71151 NAND2X1_LOC_785/a_36_24# INVX1_LOC_84/A 0.00fF
C71152 NOR2X1_LOC_568/A INVX1_LOC_37/A 0.15fF
C71153 NOR2X1_LOC_457/a_36_216# NOR2X1_LOC_155/A 0.00fF
C71154 NOR2X1_LOC_481/A INVX1_LOC_91/A 0.06fF
C71155 NOR2X1_LOC_647/Y VDD 0.12fF
C71156 INVX1_LOC_1/A INVX1_LOC_92/A 0.54fF
C71157 INVX1_LOC_269/A NOR2X1_LOC_78/Y 0.01fF
C71158 INVX1_LOC_57/A NAND2X1_LOC_254/Y 0.03fF
C71159 NOR2X1_LOC_637/Y NOR2X1_LOC_56/Y 0.10fF
C71160 NOR2X1_LOC_631/B INVX1_LOC_71/A 0.07fF
C71161 NOR2X1_LOC_112/Y NOR2X1_LOC_196/a_36_216# 0.02fF
C71162 INVX1_LOC_18/A VDD 1.82fF
C71163 NOR2X1_LOC_516/B NOR2X1_LOC_19/B 0.10fF
C71164 NAND2X1_LOC_276/Y NOR2X1_LOC_78/A 0.02fF
C71165 INVX1_LOC_32/A NAND2X1_LOC_288/B 0.10fF
C71166 INVX1_LOC_36/A NOR2X1_LOC_363/Y 0.02fF
C71167 NOR2X1_LOC_264/Y NOR2X1_LOC_557/A 0.10fF
C71168 INVX1_LOC_230/Y NOR2X1_LOC_96/Y 0.35fF
C71169 NOR2X1_LOC_208/Y NOR2X1_LOC_556/a_36_216# 0.00fF
C71170 INVX1_LOC_271/A NAND2X1_LOC_791/a_36_24# 0.00fF
C71171 D_INPUT_1 INVX1_LOC_290/Y 0.09fF
C71172 INVX1_LOC_182/A NOR2X1_LOC_540/a_36_216# 0.01fF
C71173 INVX1_LOC_34/A NAND2X1_LOC_623/B 0.02fF
C71174 INVX1_LOC_72/A INVX1_LOC_77/Y 1.76fF
C71175 INVX1_LOC_225/A INVX1_LOC_91/A 0.28fF
C71176 NOR2X1_LOC_561/Y NOR2X1_LOC_597/A 0.06fF
C71177 NAND2X1_LOC_728/Y NAND2X1_LOC_800/A 0.03fF
C71178 NOR2X1_LOC_355/A INVX1_LOC_313/A 0.04fF
C71179 NOR2X1_LOC_577/Y NOR2X1_LOC_137/B 0.01fF
C71180 NAND2X1_LOC_181/Y INPUT_0 0.07fF
C71181 NAND2X1_LOC_803/B INVX1_LOC_291/A 0.07fF
C71182 NAND2X1_LOC_661/a_36_24# NAND2X1_LOC_661/B 0.00fF
C71183 NAND2X1_LOC_729/B NAND2X1_LOC_811/Y 0.02fF
C71184 INVX1_LOC_298/Y INVX1_LOC_271/Y 0.07fF
C71185 INVX1_LOC_256/A NOR2X1_LOC_650/a_36_216# 0.00fF
C71186 NOR2X1_LOC_637/Y INVX1_LOC_146/Y 0.01fF
C71187 NAND2X1_LOC_711/B VDD 0.01fF
C71188 NOR2X1_LOC_754/A NOR2X1_LOC_754/Y 0.00fF
C71189 NOR2X1_LOC_637/Y VDD 0.23fF
C71190 NAND2X1_LOC_551/A NOR2X1_LOC_71/Y 0.38fF
C71191 NAND2X1_LOC_854/B INVX1_LOC_140/A 0.19fF
C71192 INVX1_LOC_71/A INVX1_LOC_37/A 3.22fF
C71193 INVX1_LOC_95/Y INVX1_LOC_8/A 1.43fF
C71194 INVX1_LOC_64/A NAND2X1_LOC_233/a_36_24# 0.00fF
C71195 NAND2X1_LOC_63/Y NOR2X1_LOC_849/A 0.00fF
C71196 NOR2X1_LOC_590/A INVX1_LOC_291/A 0.07fF
C71197 INVX1_LOC_172/A VDD 0.28fF
C71198 NOR2X1_LOC_15/Y NAND2X1_LOC_475/Y 0.01fF
C71199 NOR2X1_LOC_189/A INVX1_LOC_46/A 0.01fF
C71200 INVX1_LOC_64/A NOR2X1_LOC_38/a_36_216# 0.00fF
C71201 NOR2X1_LOC_728/a_36_216# NOR2X1_LOC_687/Y 0.00fF
C71202 NOR2X1_LOC_209/Y INVX1_LOC_91/A 0.07fF
C71203 INVX1_LOC_230/Y NAND2X1_LOC_848/Y 0.01fF
C71204 NOR2X1_LOC_160/B NOR2X1_LOC_216/B 0.19fF
C71205 NOR2X1_LOC_690/A INVX1_LOC_20/A 0.12fF
C71206 INVX1_LOC_53/A NOR2X1_LOC_467/A 0.05fF
C71207 NAND2X1_LOC_390/A INPUT_0 0.09fF
C71208 NOR2X1_LOC_89/A INVX1_LOC_306/Y 0.03fF
C71209 NOR2X1_LOC_389/A NOR2X1_LOC_155/A 0.76fF
C71210 NOR2X1_LOC_78/B INVX1_LOC_160/A 0.00fF
C71211 NOR2X1_LOC_440/Y NOR2X1_LOC_74/A 0.01fF
C71212 INVX1_LOC_27/A NAND2X1_LOC_207/B 0.07fF
C71213 NAND2X1_LOC_63/Y NOR2X1_LOC_440/B 0.01fF
C71214 INVX1_LOC_50/A INVX1_LOC_87/A 0.06fF
C71215 INVX1_LOC_155/Y NOR2X1_LOC_137/Y 0.27fF
C71216 NOR2X1_LOC_598/B NOR2X1_LOC_38/B 0.01fF
C71217 INVX1_LOC_23/A INVX1_LOC_253/A 0.01fF
C71218 INVX1_LOC_45/A NOR2X1_LOC_743/Y 0.68fF
C71219 NOR2X1_LOC_168/Y INVX1_LOC_9/A 0.03fF
C71220 NOR2X1_LOC_183/a_36_216# INVX1_LOC_22/A -0.01fF
C71221 INVX1_LOC_59/A INVX1_LOC_29/A 0.03fF
C71222 INVX1_LOC_10/A NOR2X1_LOC_815/A 0.00fF
C71223 INVX1_LOC_100/A NAND2X1_LOC_573/A 0.54fF
C71224 NOR2X1_LOC_227/B NOR2X1_LOC_340/A 0.00fF
C71225 NAND2X1_LOC_550/A NAND2X1_LOC_477/Y 0.01fF
C71226 NAND2X1_LOC_464/B INVX1_LOC_23/Y 0.45fF
C71227 INVX1_LOC_41/Y INVX1_LOC_118/A 0.03fF
C71228 NAND2X1_LOC_852/Y INVX1_LOC_11/Y 0.03fF
C71229 NOR2X1_LOC_219/B INVX1_LOC_281/A 0.02fF
C71230 INVX1_LOC_34/A INVX1_LOC_117/A 0.16fF
C71231 INVX1_LOC_225/A NOR2X1_LOC_653/a_36_216# 0.00fF
C71232 NAND2X1_LOC_338/B NAND2X1_LOC_465/A 0.01fF
C71233 NOR2X1_LOC_471/Y NOR2X1_LOC_257/Y 0.00fF
C71234 NOR2X1_LOC_617/Y INVX1_LOC_118/A 0.00fF
C71235 NOR2X1_LOC_287/a_36_216# INVX1_LOC_117/A 0.01fF
C71236 NOR2X1_LOC_355/A INVX1_LOC_6/A 0.03fF
C71237 NAND2X1_LOC_593/Y INVX1_LOC_118/A 0.10fF
C71238 INVX1_LOC_24/A NOR2X1_LOC_433/Y 0.17fF
C71239 INVX1_LOC_71/A NOR2X1_LOC_177/Y 0.07fF
C71240 NOR2X1_LOC_482/Y INVX1_LOC_46/A 0.37fF
C71241 VDD INVX1_LOC_34/Y 0.24fF
C71242 INVX1_LOC_173/Y NOR2X1_LOC_387/A 0.02fF
C71243 INVX1_LOC_71/A NOR2X1_LOC_743/Y 0.31fF
C71244 NAND2X1_LOC_852/Y NOR2X1_LOC_421/Y 0.18fF
C71245 INVX1_LOC_137/Y NAND2X1_LOC_642/Y 0.01fF
C71246 NOR2X1_LOC_822/Y NOR2X1_LOC_822/a_36_216# 0.01fF
C71247 NOR2X1_LOC_596/A NOR2X1_LOC_155/A 4.60fF
C71248 INVX1_LOC_83/A INVX1_LOC_160/A 0.02fF
C71249 NOR2X1_LOC_256/Y NAND2X1_LOC_348/A 0.06fF
C71250 INVX1_LOC_105/A INVX1_LOC_117/Y 0.15fF
C71251 NAND2X1_LOC_184/a_36_24# NOR2X1_LOC_337/A 0.00fF
C71252 INVX1_LOC_69/Y NOR2X1_LOC_356/A 0.02fF
C71253 NOR2X1_LOC_736/Y INVX1_LOC_6/A 0.03fF
C71254 INVX1_LOC_22/A NAND2X1_LOC_267/B 0.01fF
C71255 INVX1_LOC_25/A INVX1_LOC_53/A 0.02fF
C71256 NOR2X1_LOC_791/B INVX1_LOC_63/A 1.85fF
C71257 NAND2X1_LOC_354/B INVX1_LOC_291/A 0.19fF
C71258 NOR2X1_LOC_63/a_36_216# INVX1_LOC_9/A 0.00fF
C71259 NAND2X1_LOC_778/Y NOR2X1_LOC_167/a_36_216# 0.12fF
C71260 INVX1_LOC_290/A INVX1_LOC_46/A 0.05fF
C71261 NOR2X1_LOC_16/Y INVX1_LOC_9/A 0.01fF
C71262 NAND2X1_LOC_170/A NAND2X1_LOC_804/Y 0.14fF
C71263 NAND2X1_LOC_20/B INVX1_LOC_15/A 0.17fF
C71264 NAND2X1_LOC_348/A NOR2X1_LOC_391/a_36_216# 0.00fF
C71265 NOR2X1_LOC_19/B INVX1_LOC_315/Y 0.06fF
C71266 NOR2X1_LOC_690/Y VDD 0.47fF
C71267 INVX1_LOC_221/A INVX1_LOC_92/A 0.03fF
C71268 INVX1_LOC_69/Y NOR2X1_LOC_74/A 0.07fF
C71269 INVX1_LOC_2/A INVX1_LOC_185/A 0.03fF
C71270 NOR2X1_LOC_826/Y INVX1_LOC_64/A 0.01fF
C71271 INVX1_LOC_21/A NOR2X1_LOC_383/B 0.07fF
C71272 NAND2X1_LOC_341/A INVX1_LOC_38/A 0.08fF
C71273 NOR2X1_LOC_15/Y NOR2X1_LOC_167/a_36_216# 0.00fF
C71274 INVX1_LOC_63/Y NOR2X1_LOC_435/B 0.14fF
C71275 NOR2X1_LOC_350/A NOR2X1_LOC_68/Y 0.01fF
C71276 NOR2X1_LOC_226/A INVX1_LOC_185/A 0.03fF
C71277 INVX1_LOC_303/A NOR2X1_LOC_691/B 0.02fF
C71278 NAND2X1_LOC_208/B INVX1_LOC_3/Y 0.10fF
C71279 INVX1_LOC_276/Y INVX1_LOC_291/A 0.01fF
C71280 NOR2X1_LOC_168/B NOR2X1_LOC_862/B 0.05fF
C71281 NAND2X1_LOC_660/Y NOR2X1_LOC_536/A 0.00fF
C71282 NAND2X1_LOC_99/A NOR2X1_LOC_271/B 0.01fF
C71283 NOR2X1_LOC_272/Y INVX1_LOC_23/A 0.37fF
C71284 NAND2X1_LOC_720/a_36_24# NOR2X1_LOC_48/B -0.00fF
C71285 NOR2X1_LOC_541/Y NAND2X1_LOC_72/B 0.02fF
C71286 GATE_479 INVX1_LOC_38/A 0.03fF
C71287 NAND2X1_LOC_778/Y NAND2X1_LOC_787/A 0.01fF
C71288 INVX1_LOC_232/A NOR2X1_LOC_489/A 0.17fF
C71289 NOR2X1_LOC_246/A NAND2X1_LOC_284/a_36_24# 0.00fF
C71290 INVX1_LOC_35/A INVX1_LOC_13/Y 0.14fF
C71291 INVX1_LOC_311/Y INVX1_LOC_76/A 0.03fF
C71292 INVX1_LOC_230/Y NAND2X1_LOC_223/A 0.07fF
C71293 NOR2X1_LOC_757/A NOR2X1_LOC_331/B 0.04fF
C71294 INVX1_LOC_153/Y INVX1_LOC_186/Y 0.10fF
C71295 NOR2X1_LOC_220/A NOR2X1_LOC_155/A 0.03fF
C71296 NOR2X1_LOC_644/B NAND2X1_LOC_454/Y 0.02fF
C71297 NOR2X1_LOC_552/A NOR2X1_LOC_337/A 0.03fF
C71298 NOR2X1_LOC_181/a_36_216# INVX1_LOC_271/Y 0.00fF
C71299 D_INPUT_0 NOR2X1_LOC_536/A 0.25fF
C71300 NOR2X1_LOC_32/B INVX1_LOC_234/Y 0.04fF
C71301 NOR2X1_LOC_148/B NOR2X1_LOC_808/B 0.16fF
C71302 INVX1_LOC_272/Y NOR2X1_LOC_654/A 0.35fF
C71303 NOR2X1_LOC_802/A INVX1_LOC_63/A 0.01fF
C71304 INVX1_LOC_121/Y INVX1_LOC_186/Y 0.00fF
C71305 NAND2X1_LOC_807/Y NOR2X1_LOC_111/A 0.14fF
C71306 NAND2X1_LOC_35/Y NOR2X1_LOC_496/Y 0.05fF
C71307 INVX1_LOC_16/A NAND2X1_LOC_243/B 0.20fF
C71308 NAND2X1_LOC_787/A NOR2X1_LOC_15/Y 0.03fF
C71309 NOR2X1_LOC_274/B INVX1_LOC_4/Y 0.03fF
C71310 INVX1_LOC_90/A INVX1_LOC_44/A 0.07fF
C71311 NOR2X1_LOC_516/B NOR2X1_LOC_216/B 0.03fF
C71312 INVX1_LOC_1/A INVX1_LOC_53/A 2.27fF
C71313 INVX1_LOC_208/Y NOR2X1_LOC_831/B 0.01fF
C71314 INVX1_LOC_45/A NAND2X1_LOC_72/B 0.12fF
C71315 INVX1_LOC_31/Y VDD 0.45fF
C71316 INVX1_LOC_269/A NAND2X1_LOC_860/A 0.19fF
C71317 INVX1_LOC_64/A NAND2X1_LOC_705/Y 0.04fF
C71318 NOR2X1_LOC_568/A NAND2X1_LOC_72/B 0.07fF
C71319 INVX1_LOC_235/Y NOR2X1_LOC_663/A 0.01fF
C71320 NOR2X1_LOC_15/Y NAND2X1_LOC_363/B 1.01fF
C71321 NOR2X1_LOC_345/A NOR2X1_LOC_260/Y 0.05fF
C71322 NOR2X1_LOC_441/Y NOR2X1_LOC_282/Y 0.01fF
C71323 INVX1_LOC_64/A NAND2X1_LOC_303/Y 0.07fF
C71324 INVX1_LOC_90/A NOR2X1_LOC_96/a_36_216# 0.00fF
C71325 INVX1_LOC_78/Y INVX1_LOC_247/A 0.01fF
C71326 INVX1_LOC_35/A INVX1_LOC_88/A 0.06fF
C71327 INVX1_LOC_177/Y INVX1_LOC_78/A 0.61fF
C71328 INVX1_LOC_91/A NAND2X1_LOC_642/Y 0.12fF
C71329 INVX1_LOC_97/Y NAND2X1_LOC_190/Y 0.17fF
C71330 NAND2X1_LOC_553/A INVX1_LOC_48/Y 0.01fF
C71331 NOR2X1_LOC_92/Y INVX1_LOC_5/A 0.03fF
C71332 D_INPUT_0 NAND2X1_LOC_93/B 0.03fF
C71333 NOR2X1_LOC_400/A INVX1_LOC_14/A 0.10fF
C71334 NOR2X1_LOC_375/Y INVX1_LOC_84/A 0.00fF
C71335 NOR2X1_LOC_561/Y NOR2X1_LOC_88/Y 0.01fF
C71336 NOR2X1_LOC_300/Y INVX1_LOC_12/A 0.02fF
C71337 NAND2X1_LOC_671/a_36_24# NOR2X1_LOC_814/A 0.01fF
C71338 NOR2X1_LOC_389/A NOR2X1_LOC_125/Y 0.10fF
C71339 INVX1_LOC_58/A INVX1_LOC_161/A 0.01fF
C71340 INVX1_LOC_41/A NOR2X1_LOC_462/a_36_216# 0.00fF
C71341 INVX1_LOC_243/A NAND2X1_LOC_651/B 0.08fF
C71342 NOR2X1_LOC_794/B INVX1_LOC_53/A 0.00fF
C71343 NAND2X1_LOC_725/Y NAND2X1_LOC_733/Y 0.56fF
C71344 INVX1_LOC_104/A INVX1_LOC_42/A 0.07fF
C71345 NOR2X1_LOC_719/A INVX1_LOC_84/A 0.03fF
C71346 NOR2X1_LOC_130/A NAND2X1_LOC_798/B 0.08fF
C71347 INPUT_0 INVX1_LOC_117/A 0.11fF
C71348 NOR2X1_LOC_15/Y NOR2X1_LOC_791/Y 0.02fF
C71349 NOR2X1_LOC_557/Y INVX1_LOC_47/Y 0.18fF
C71350 INVX1_LOC_34/A INVX1_LOC_3/Y 0.26fF
C71351 INVX1_LOC_71/A NAND2X1_LOC_72/B 0.05fF
C71352 NOR2X1_LOC_92/Y INVX1_LOC_178/A 0.19fF
C71353 NOR2X1_LOC_598/B NOR2X1_LOC_389/A 0.10fF
C71354 INVX1_LOC_191/Y NOR2X1_LOC_583/Y 0.01fF
C71355 NOR2X1_LOC_242/A INVX1_LOC_1/A 0.00fF
C71356 NOR2X1_LOC_561/Y INVX1_LOC_84/A 0.07fF
C71357 NOR2X1_LOC_336/B INVX1_LOC_23/A 0.00fF
C71358 INVX1_LOC_11/A INVX1_LOC_306/Y 0.07fF
C71359 NAND2X1_LOC_740/A NAND2X1_LOC_175/Y 0.03fF
C71360 INVX1_LOC_36/A INVX1_LOC_29/Y 1.20fF
C71361 INVX1_LOC_58/A NOR2X1_LOC_722/Y 0.03fF
C71362 INVX1_LOC_50/A NAND2X1_LOC_514/Y 0.06fF
C71363 D_INPUT_0 NOR2X1_LOC_649/B 0.14fF
C71364 VDD NAND2X1_LOC_86/Y -0.00fF
C71365 NOR2X1_LOC_781/A INVX1_LOC_19/A 0.07fF
C71366 D_INPUT_0 INVX1_LOC_3/A 0.61fF
C71367 NOR2X1_LOC_560/A NAND2X1_LOC_85/Y 0.26fF
C71368 NAND2X1_LOC_652/Y INVX1_LOC_117/Y 0.00fF
C71369 NAND2X1_LOC_364/A INVX1_LOC_23/A 0.08fF
C71370 INVX1_LOC_224/Y NAND2X1_LOC_198/B 0.33fF
C71371 NOR2X1_LOC_775/Y NAND2X1_LOC_413/a_36_24# 0.00fF
C71372 NOR2X1_LOC_246/a_36_216# INVX1_LOC_285/A 0.00fF
C71373 INVX1_LOC_35/A NOR2X1_LOC_500/B 0.04fF
C71374 NOR2X1_LOC_99/B NOR2X1_LOC_673/a_36_216# 0.01fF
C71375 NAND2X1_LOC_725/B NAND2X1_LOC_561/B 0.03fF
C71376 NAND2X1_LOC_850/a_36_24# INVX1_LOC_26/A 0.00fF
C71377 NOR2X1_LOC_468/Y NOR2X1_LOC_271/a_36_216# 0.00fF
C71378 NOR2X1_LOC_71/Y NAND2X1_LOC_489/Y 0.02fF
C71379 INVX1_LOC_16/A INVX1_LOC_284/A 0.12fF
C71380 INVX1_LOC_75/A NOR2X1_LOC_156/Y 0.03fF
C71381 INVX1_LOC_143/A INVX1_LOC_47/Y 0.00fF
C71382 INVX1_LOC_113/Y NOR2X1_LOC_632/a_36_216# 0.00fF
C71383 INVX1_LOC_6/A INVX1_LOC_127/A 0.00fF
C71384 INVX1_LOC_104/A INVX1_LOC_78/A 0.14fF
C71385 INVX1_LOC_314/Y INVX1_LOC_57/A 0.10fF
C71386 INVX1_LOC_279/A INVX1_LOC_29/A 0.06fF
C71387 INVX1_LOC_236/A INVX1_LOC_21/Y 0.02fF
C71388 NOR2X1_LOC_553/Y INVX1_LOC_290/Y 0.01fF
C71389 INVX1_LOC_123/A INVX1_LOC_9/A 0.21fF
C71390 INVX1_LOC_234/A NAND2X1_LOC_81/a_36_24# -0.00fF
C71391 NOR2X1_LOC_92/Y NAND2X1_LOC_337/B 0.07fF
C71392 NOR2X1_LOC_376/A INVX1_LOC_174/A 0.04fF
C71393 NOR2X1_LOC_15/Y NOR2X1_LOC_457/A 0.01fF
C71394 INVX1_LOC_28/A INVX1_LOC_119/Y 0.01fF
C71395 INVX1_LOC_91/A NOR2X1_LOC_271/Y 0.07fF
C71396 NOR2X1_LOC_188/A INVX1_LOC_92/A 0.17fF
C71397 NOR2X1_LOC_598/B NOR2X1_LOC_596/A 0.14fF
C71398 INVX1_LOC_49/A INVX1_LOC_270/Y 0.73fF
C71399 INVX1_LOC_289/Y NAND2X1_LOC_227/Y 0.02fF
C71400 NOR2X1_LOC_428/Y NOR2X1_LOC_763/A 0.08fF
C71401 NOR2X1_LOC_92/Y NOR2X1_LOC_816/A 0.01fF
C71402 NOR2X1_LOC_637/B INVX1_LOC_271/A 0.13fF
C71403 NOR2X1_LOC_76/A INVX1_LOC_19/A 0.07fF
C71404 INVX1_LOC_162/Y NOR2X1_LOC_318/A 0.01fF
C71405 D_INPUT_1 INVX1_LOC_77/A 0.76fF
C71406 NOR2X1_LOC_548/B INVX1_LOC_92/A 0.10fF
C71407 NAND2X1_LOC_453/a_36_24# NOR2X1_LOC_449/A 0.00fF
C71408 NAND2X1_LOC_778/Y INVX1_LOC_30/A 0.03fF
C71409 INVX1_LOC_35/A NOR2X1_LOC_758/a_36_216# 0.00fF
C71410 NOR2X1_LOC_346/B INVX1_LOC_4/Y 0.00fF
C71411 NAND2X1_LOC_9/Y NOR2X1_LOC_350/A 0.02fF
C71412 INVX1_LOC_21/A INVX1_LOC_57/Y 0.07fF
C71413 NOR2X1_LOC_88/Y NOR2X1_LOC_167/Y 0.03fF
C71414 INVX1_LOC_255/Y INVX1_LOC_32/A 0.04fF
C71415 INVX1_LOC_78/Y NOR2X1_LOC_676/Y 0.11fF
C71416 NOR2X1_LOC_65/B INVX1_LOC_104/A 0.10fF
C71417 NOR2X1_LOC_510/Y INVX1_LOC_18/A 0.07fF
C71418 INVX1_LOC_35/A INVX1_LOC_303/A 0.07fF
C71419 INVX1_LOC_58/A INVX1_LOC_34/A 0.31fF
C71420 NOR2X1_LOC_75/Y NAND2X1_LOC_53/Y 0.01fF
C71421 NOR2X1_LOC_91/A NAND2X1_LOC_785/A 0.15fF
C71422 INVX1_LOC_41/A NOR2X1_LOC_828/Y 0.11fF
C71423 INVX1_LOC_226/Y NOR2X1_LOC_394/Y 0.01fF
C71424 INVX1_LOC_5/A NAND2X1_LOC_837/Y 0.01fF
C71425 INVX1_LOC_22/A INVX1_LOC_4/Y 0.15fF
C71426 NOR2X1_LOC_561/Y INVX1_LOC_15/A 0.08fF
C71427 NAND2X1_LOC_149/Y INVX1_LOC_72/A 0.14fF
C71428 NOR2X1_LOC_790/B NOR2X1_LOC_551/B 0.02fF
C71429 NOR2X1_LOC_773/Y NOR2X1_LOC_281/a_36_216# 0.01fF
C71430 INVX1_LOC_17/A NAND2X1_LOC_555/Y 0.09fF
C71431 NOR2X1_LOC_455/Y NOR2X1_LOC_445/Y 0.01fF
C71432 NOR2X1_LOC_309/Y INVX1_LOC_29/Y 0.40fF
C71433 NAND2X1_LOC_32/a_36_24# INVX1_LOC_205/A 0.02fF
C71434 NOR2X1_LOC_329/B INVX1_LOC_272/A 0.97fF
C71435 NOR2X1_LOC_15/Y INVX1_LOC_30/A 0.36fF
C71436 INVX1_LOC_21/A NOR2X1_LOC_480/A 0.10fF
C71437 NOR2X1_LOC_266/B NOR2X1_LOC_536/A 0.07fF
C71438 INVX1_LOC_73/A INVX1_LOC_19/A 0.03fF
C71439 NOR2X1_LOC_381/Y NOR2X1_LOC_382/Y 0.02fF
C71440 INVX1_LOC_256/A NOR2X1_LOC_275/a_36_216# 0.00fF
C71441 INVX1_LOC_227/A NOR2X1_LOC_609/Y 0.00fF
C71442 NOR2X1_LOC_811/A NOR2X1_LOC_855/A 0.05fF
C71443 NOR2X1_LOC_82/A INVX1_LOC_61/Y 0.91fF
C71444 NOR2X1_LOC_763/A NOR2X1_LOC_582/Y 0.02fF
C71445 NAND2X1_LOC_833/Y NAND2X1_LOC_790/a_36_24# 0.01fF
C71446 INVX1_LOC_160/Y NOR2X1_LOC_839/B 0.01fF
C71447 INVX1_LOC_83/A NOR2X1_LOC_467/A 0.03fF
C71448 NOR2X1_LOC_215/A NOR2X1_LOC_215/Y 0.30fF
C71449 NOR2X1_LOC_582/A NOR2X1_LOC_582/Y 0.10fF
C71450 INVX1_LOC_124/A D_INPUT_1 0.07fF
C71451 INVX1_LOC_64/A NOR2X1_LOC_690/A 0.07fF
C71452 INVX1_LOC_221/A INVX1_LOC_53/A 0.14fF
C71453 NOR2X1_LOC_71/Y INVX1_LOC_32/A 0.10fF
C71454 INVX1_LOC_178/A NAND2X1_LOC_837/Y 0.10fF
C71455 NAND2X1_LOC_357/B INVX1_LOC_308/A 0.01fF
C71456 NOR2X1_LOC_618/a_36_216# INVX1_LOC_26/A 0.00fF
C71457 INVX1_LOC_37/A NOR2X1_LOC_331/B 0.15fF
C71458 INVX1_LOC_64/A NOR2X1_LOC_413/Y 0.08fF
C71459 INVX1_LOC_256/A INVX1_LOC_124/Y 0.03fF
C71460 INVX1_LOC_41/A INVX1_LOC_5/A 3.44fF
C71461 NAND2X1_LOC_563/Y NOR2X1_LOC_660/Y 0.11fF
C71462 INVX1_LOC_58/A NAND2X1_LOC_231/Y 0.10fF
C71463 NAND2X1_LOC_9/Y NOR2X1_LOC_84/Y 0.07fF
C71464 INVX1_LOC_285/Y INVX1_LOC_186/Y 0.07fF
C71465 NOR2X1_LOC_355/A NAND2X1_LOC_646/a_36_24# 0.00fF
C71466 NAND2X1_LOC_11/Y INVX1_LOC_23/A 0.06fF
C71467 INVX1_LOC_201/Y INVX1_LOC_5/A 0.16fF
C71468 INVX1_LOC_13/A INVX1_LOC_16/Y 0.98fF
C71469 INVX1_LOC_50/A INVX1_LOC_278/Y 0.14fF
C71470 INVX1_LOC_25/A NOR2X1_LOC_78/B 0.08fF
C71471 NOR2X1_LOC_704/Y INVX1_LOC_19/A 0.02fF
C71472 NOR2X1_LOC_356/A NOR2X1_LOC_170/A 0.03fF
C71473 NAND2X1_LOC_840/a_36_24# NOR2X1_LOC_109/Y 0.01fF
C71474 INVX1_LOC_233/A NOR2X1_LOC_84/Y 0.40fF
C71475 NOR2X1_LOC_644/A INVX1_LOC_32/A 0.03fF
C71476 INVX1_LOC_251/Y NOR2X1_LOC_717/A 0.01fF
C71477 NAND2X1_LOC_848/A NOR2X1_LOC_536/A 0.04fF
C71478 NOR2X1_LOC_155/A NAND2X1_LOC_469/B 2.12fF
C71479 NOR2X1_LOC_145/a_36_216# NAND2X1_LOC_93/B 0.00fF
C71480 INVX1_LOC_298/Y INVX1_LOC_279/A 0.07fF
C71481 NOR2X1_LOC_500/A NOR2X1_LOC_793/A 0.15fF
C71482 INVX1_LOC_44/A INVX1_LOC_38/A 0.07fF
C71483 NOR2X1_LOC_494/Y NAND2X1_LOC_837/Y 0.04fF
C71484 INVX1_LOC_27/A INVX1_LOC_155/A 0.03fF
C71485 NOR2X1_LOC_74/A NOR2X1_LOC_89/A 0.23fF
C71486 INVX1_LOC_1/A INVX1_LOC_184/A 0.02fF
C71487 INVX1_LOC_13/A NOR2X1_LOC_39/Y 0.01fF
C71488 NOR2X1_LOC_815/A INVX1_LOC_12/A 0.04fF
C71489 NOR2X1_LOC_689/Y NAND2X1_LOC_863/B 0.08fF
C71490 NAND2X1_LOC_198/B NOR2X1_LOC_103/Y 0.13fF
C71491 NOR2X1_LOC_88/Y INVX1_LOC_76/A 0.07fF
C71492 NOR2X1_LOC_145/a_36_216# NAND2X1_LOC_425/Y 0.01fF
C71493 NOR2X1_LOC_598/B NOR2X1_LOC_220/A 0.11fF
C71494 NOR2X1_LOC_9/Y NOR2X1_LOC_89/A 0.02fF
C71495 INVX1_LOC_124/A NOR2X1_LOC_652/Y 0.55fF
C71496 NOR2X1_LOC_443/Y NAND2X1_LOC_358/Y 0.04fF
C71497 INVX1_LOC_75/A D_INPUT_5 0.19fF
C71498 INVX1_LOC_37/A NOR2X1_LOC_592/B 0.33fF
C71499 INVX1_LOC_59/A INVX1_LOC_8/A 0.10fF
C71500 NOR2X1_LOC_679/Y INVX1_LOC_24/A 0.01fF
C71501 NAND2X1_LOC_364/A INVX1_LOC_31/A 0.10fF
C71502 NOR2X1_LOC_565/B NOR2X1_LOC_383/B 0.01fF
C71503 NOR2X1_LOC_205/Y NOR2X1_LOC_577/Y 0.02fF
C71504 NOR2X1_LOC_78/A INVX1_LOC_125/A 0.03fF
C71505 NOR2X1_LOC_137/a_36_216# NAND2X1_LOC_475/Y 0.12fF
C71506 INVX1_LOC_89/A INVX1_LOC_26/A 0.05fF
C71507 NAND2X1_LOC_735/B NOR2X1_LOC_629/A 0.01fF
C71508 INVX1_LOC_212/A NOR2X1_LOC_160/B 0.02fF
C71509 NOR2X1_LOC_576/B NAND2X1_LOC_828/a_36_24# 0.04fF
C71510 NOR2X1_LOC_34/A NOR2X1_LOC_87/B 0.06fF
C71511 NAND2X1_LOC_773/Y INVX1_LOC_8/A 0.02fF
C71512 INPUT_0 INVX1_LOC_3/Y 0.14fF
C71513 NOR2X1_LOC_500/A NOR2X1_LOC_160/B 0.07fF
C71514 INVX1_LOC_84/A INVX1_LOC_76/A 0.32fF
C71515 NAND2X1_LOC_100/a_36_24# INVX1_LOC_31/A 0.00fF
C71516 NOR2X1_LOC_355/A INVX1_LOC_270/A 0.10fF
C71517 NOR2X1_LOC_92/Y NAND2X1_LOC_562/B 0.02fF
C71518 NAND2X1_LOC_813/a_36_24# NAND2X1_LOC_207/B 0.01fF
C71519 NAND2X1_LOC_493/Y INVX1_LOC_240/A 0.08fF
C71520 INVX1_LOC_233/Y INVX1_LOC_22/A 0.05fF
C71521 NOR2X1_LOC_536/A INVX1_LOC_46/Y 0.08fF
C71522 INVX1_LOC_269/A NOR2X1_LOC_516/Y 0.04fF
C71523 NAND2X1_LOC_579/A NAND2X1_LOC_357/B 0.03fF
C71524 INVX1_LOC_98/Y NAND2X1_LOC_474/Y 0.01fF
C71525 INVX1_LOC_1/A INVX1_LOC_80/Y 0.00fF
C71526 INPUT_6 INPUT_5 0.02fF
C71527 INVX1_LOC_303/Y INVX1_LOC_15/A 0.04fF
C71528 NOR2X1_LOC_167/Y INVX1_LOC_15/A 0.07fF
C71529 INVX1_LOC_25/A INVX1_LOC_83/A 0.25fF
C71530 INVX1_LOC_45/A NAND2X1_LOC_198/B 1.85fF
C71531 NAND2X1_LOC_624/B NAND2X1_LOC_735/B 0.03fF
C71532 INVX1_LOC_2/Y INVX1_LOC_63/A 0.18fF
C71533 NAND2X1_LOC_784/A NAND2X1_LOC_808/A 0.44fF
C71534 INVX1_LOC_298/Y INVX1_LOC_182/Y 0.03fF
C71535 NOR2X1_LOC_594/Y NOR2X1_LOC_158/B 0.02fF
C71536 NOR2X1_LOC_205/Y NOR2X1_LOC_348/B 0.02fF
C71537 NAND2X1_LOC_626/a_36_24# INVX1_LOC_284/A 0.00fF
C71538 NOR2X1_LOC_15/Y NAND2X1_LOC_722/A 0.02fF
C71539 NAND2X1_LOC_578/B INVX1_LOC_239/A 0.00fF
C71540 NOR2X1_LOC_9/Y INVX1_LOC_104/Y 0.01fF
C71541 INVX1_LOC_224/Y NOR2X1_LOC_76/a_36_216# 0.01fF
C71542 NOR2X1_LOC_255/Y INVX1_LOC_89/A 0.01fF
C71543 INVX1_LOC_136/A INVX1_LOC_181/Y 0.09fF
C71544 NOR2X1_LOC_254/A NOR2X1_LOC_147/B 0.80fF
C71545 NOR2X1_LOC_736/Y INVX1_LOC_270/A 0.16fF
C71546 NAND2X1_LOC_725/A NAND2X1_LOC_795/Y 0.03fF
C71547 NAND2X1_LOC_364/A INVX1_LOC_111/A 0.01fF
C71548 NOR2X1_LOC_92/Y NOR2X1_LOC_773/Y 0.07fF
C71549 NOR2X1_LOC_78/B INVX1_LOC_1/A 0.19fF
C71550 NOR2X1_LOC_179/Y NOR2X1_LOC_271/Y 0.11fF
C71551 NAND2X1_LOC_337/B NAND2X1_LOC_477/A 0.10fF
C71552 NAND2X1_LOC_741/B INVX1_LOC_209/Y 0.02fF
C71553 NOR2X1_LOC_209/Y NOR2X1_LOC_739/Y 0.00fF
C71554 NAND2X1_LOC_588/a_36_24# INVX1_LOC_1/A 0.01fF
C71555 NAND2X1_LOC_513/B NOR2X1_LOC_516/B 0.11fF
C71556 NAND2X1_LOC_93/B INVX1_LOC_46/Y 0.02fF
C71557 NOR2X1_LOC_425/Y NOR2X1_LOC_36/B 0.00fF
C71558 NAND2X1_LOC_848/A NOR2X1_LOC_661/A 0.14fF
C71559 INVX1_LOC_206/Y INVX1_LOC_78/A 2.53fF
C71560 NOR2X1_LOC_48/a_36_216# INVX1_LOC_117/A 0.01fF
C71561 INVX1_LOC_45/A INVX1_LOC_310/Y 0.72fF
C71562 NAND2X1_LOC_198/B INVX1_LOC_71/A 0.10fF
C71563 INVX1_LOC_186/A NOR2X1_LOC_334/Y 0.07fF
C71564 NOR2X1_LOC_45/B INVX1_LOC_128/Y 0.07fF
C71565 INVX1_LOC_269/A INVX1_LOC_172/Y 0.02fF
C71566 NOR2X1_LOC_340/Y INVX1_LOC_110/A 0.20fF
C71567 NAND2X1_LOC_785/A INVX1_LOC_31/A 0.07fF
C71568 INVX1_LOC_230/Y NOR2X1_LOC_521/a_36_216# 0.00fF
C71569 NOR2X1_LOC_667/Y INVX1_LOC_2/A 0.04fF
C71570 INVX1_LOC_311/A NOR2X1_LOC_383/B 0.07fF
C71571 NOR2X1_LOC_635/A INVX1_LOC_30/A 0.02fF
C71572 NOR2X1_LOC_78/B NOR2X1_LOC_794/B 0.01fF
C71573 NOR2X1_LOC_382/Y NOR2X1_LOC_6/B 0.08fF
C71574 INVX1_LOC_153/Y INVX1_LOC_18/A 0.25fF
C71575 NOR2X1_LOC_205/Y INVX1_LOC_22/A 0.05fF
C71576 NOR2X1_LOC_803/A INVX1_LOC_213/A 0.04fF
C71577 INVX1_LOC_266/A NOR2X1_LOC_577/a_36_216# 0.01fF
C71578 INVX1_LOC_78/A NOR2X1_LOC_600/Y 0.03fF
C71579 NOR2X1_LOC_657/Y NOR2X1_LOC_52/B 0.02fF
C71580 INVX1_LOC_14/A NOR2X1_LOC_589/A 0.72fF
C71581 INVX1_LOC_58/A INPUT_0 0.13fF
C71582 INVX1_LOC_76/A INVX1_LOC_15/A 0.13fF
C71583 NOR2X1_LOC_103/Y INVX1_LOC_53/Y -0.04fF
C71584 NOR2X1_LOC_272/Y INVX1_LOC_313/A 0.03fF
C71585 NOR2X1_LOC_454/Y NOR2X1_LOC_747/a_36_216# 0.01fF
C71586 NAND2X1_LOC_581/Y INVX1_LOC_18/A 0.02fF
C71587 NOR2X1_LOC_607/Y INVX1_LOC_77/A 0.04fF
C71588 NOR2X1_LOC_231/B INVX1_LOC_143/A 0.04fF
C71589 NAND2X1_LOC_243/Y NAND2X1_LOC_489/Y 0.23fF
C71590 INVX1_LOC_14/A NAND2X1_LOC_377/Y 0.30fF
C71591 INVX1_LOC_18/A INVX1_LOC_121/Y 0.47fF
C71592 INVX1_LOC_46/Y INVX1_LOC_3/A 0.23fF
C71593 INVX1_LOC_230/Y INVX1_LOC_40/A 0.03fF
C71594 NAND2X1_LOC_447/Y NOR2X1_LOC_334/Y 0.10fF
C71595 INVX1_LOC_11/A NAND2X1_LOC_149/B 0.02fF
C71596 NOR2X1_LOC_817/Y INVX1_LOC_13/A 0.02fF
C71597 NOR2X1_LOC_188/A INVX1_LOC_53/A 0.03fF
C71598 NOR2X1_LOC_814/Y NAND2X1_LOC_473/A 0.03fF
C71599 NOR2X1_LOC_500/A NOR2X1_LOC_317/B 0.10fF
C71600 NOR2X1_LOC_523/B NAND2X1_LOC_116/A 0.01fF
C71601 INVX1_LOC_103/A NAND2X1_LOC_319/A 0.03fF
C71602 INVX1_LOC_1/A INVX1_LOC_83/A 8.35fF
C71603 NOR2X1_LOC_815/Y NAND2X1_LOC_593/Y 0.03fF
C71604 INVX1_LOC_18/A INVX1_LOC_177/A 0.03fF
C71605 NAND2X1_LOC_717/Y INVX1_LOC_72/A 0.03fF
C71606 INVX1_LOC_255/Y INPUT_3 2.31fF
C71607 INVX1_LOC_57/Y NOR2X1_LOC_667/A 0.01fF
C71608 INVX1_LOC_278/A NOR2X1_LOC_167/Y 0.00fF
C71609 NOR2X1_LOC_557/A INVX1_LOC_57/A 0.07fF
C71610 INVX1_LOC_108/Y NAND2X1_LOC_251/a_36_24# 0.00fF
C71611 INVX1_LOC_78/A NAND2X1_LOC_220/a_36_24# 0.00fF
C71612 INVX1_LOC_132/A NAND2X1_LOC_276/Y 0.01fF
C71613 NAND2X1_LOC_562/B NAND2X1_LOC_837/Y 0.06fF
C71614 INVX1_LOC_14/A INVX1_LOC_171/A 0.03fF
C71615 INVX1_LOC_18/A NAND2X1_LOC_630/a_36_24# 0.00fF
C71616 INVX1_LOC_280/Y INVX1_LOC_18/A 0.01fF
C71617 INVX1_LOC_273/Y INVX1_LOC_161/Y 0.01fF
C71618 NOR2X1_LOC_65/B NAND2X1_LOC_674/a_36_24# 0.01fF
C71619 INVX1_LOC_31/A NOR2X1_LOC_86/A 1.18fF
C71620 INVX1_LOC_5/A NAND2X1_LOC_662/B 0.09fF
C71621 INVX1_LOC_45/A INVX1_LOC_53/Y 0.18fF
C71622 INVX1_LOC_256/A D_INPUT_0 0.10fF
C71623 NOR2X1_LOC_750/Y INVX1_LOC_91/A -0.01fF
C71624 NAND2X1_LOC_287/B NOR2X1_LOC_278/Y 0.08fF
C71625 GATE_741 NAND2X1_LOC_463/B 0.03fF
C71626 NOR2X1_LOC_405/A INVX1_LOC_23/A 0.12fF
C71627 NOR2X1_LOC_92/Y INVX1_LOC_140/A 0.10fF
C71628 INVX1_LOC_37/A NOR2X1_LOC_621/B 0.02fF
C71629 INVX1_LOC_72/A INVX1_LOC_16/A 0.34fF
C71630 NAND2X1_LOC_711/B INVX1_LOC_280/Y 0.04fF
C71631 NOR2X1_LOC_647/A VDD 0.20fF
C71632 NOR2X1_LOC_205/Y NOR2X1_LOC_735/Y 0.00fF
C71633 NOR2X1_LOC_763/A NAND2X1_LOC_51/B 0.02fF
C71634 INVX1_LOC_224/Y NAND2X1_LOC_465/A 0.02fF
C71635 NOR2X1_LOC_668/a_36_216# NAND2X1_LOC_642/Y 0.00fF
C71636 INVX1_LOC_11/A NOR2X1_LOC_356/A 0.07fF
C71637 NAND2X1_LOC_579/A NAND2X1_LOC_849/A 0.09fF
C71638 INVX1_LOC_272/Y NOR2X1_LOC_503/A 0.01fF
C71639 INVX1_LOC_45/A INVX1_LOC_145/Y 0.01fF
C71640 INVX1_LOC_12/A NAND2X1_LOC_572/B 0.65fF
C71641 NOR2X1_LOC_272/Y INVX1_LOC_6/A 1.81fF
C71642 NOR2X1_LOC_15/Y NAND2X1_LOC_856/a_36_24# 0.00fF
C71643 NOR2X1_LOC_799/B INVX1_LOC_58/Y 0.01fF
C71644 NOR2X1_LOC_328/Y INVX1_LOC_24/A 0.07fF
C71645 NOR2X1_LOC_219/Y INVX1_LOC_71/A 0.07fF
C71646 NAND2X1_LOC_724/Y VDD 0.27fF
C71647 NOR2X1_LOC_500/A NOR2X1_LOC_516/B 0.14fF
C71648 NAND2X1_LOC_21/Y INVX1_LOC_243/A 0.02fF
C71649 INVX1_LOC_247/Y INVX1_LOC_279/A 0.01fF
C71650 NOR2X1_LOC_590/A NOR2X1_LOC_788/B 0.02fF
C71651 NOR2X1_LOC_68/A NOR2X1_LOC_391/A 0.08fF
C71652 INVX1_LOC_36/A NOR2X1_LOC_355/A 0.07fF
C71653 INVX1_LOC_53/Y INVX1_LOC_71/A 0.15fF
C71654 INVX1_LOC_23/A NOR2X1_LOC_857/A 0.07fF
C71655 NOR2X1_LOC_78/A NOR2X1_LOC_81/Y 0.01fF
C71656 NAND2X1_LOC_35/Y NOR2X1_LOC_823/Y 0.03fF
C71657 INVX1_LOC_226/Y NOR2X1_LOC_419/Y 0.10fF
C71658 INVX1_LOC_25/A INVX1_LOC_46/A 0.11fF
C71659 INVX1_LOC_161/Y INVX1_LOC_73/A 0.07fF
C71660 INVX1_LOC_278/A INVX1_LOC_76/A 0.03fF
C71661 NOR2X1_LOC_158/Y INVX1_LOC_54/A 0.06fF
C71662 NOR2X1_LOC_617/Y NAND2X1_LOC_735/B 0.04fF
C71663 NOR2X1_LOC_609/A INVX1_LOC_10/A 0.06fF
C71664 INVX1_LOC_2/A NOR2X1_LOC_310/Y 0.06fF
C71665 INVX1_LOC_11/A NOR2X1_LOC_74/A 0.14fF
C71666 NAND2X1_LOC_341/A INVX1_LOC_33/A 0.03fF
C71667 NOR2X1_LOC_25/Y INVX1_LOC_54/A 0.01fF
C71668 INVX1_LOC_12/Y NOR2X1_LOC_15/a_36_216# 0.12fF
C71669 NOR2X1_LOC_50/a_36_216# INPUT_5 0.00fF
C71670 NAND2X1_LOC_714/B NAND2X1_LOC_655/A 0.15fF
C71671 INVX1_LOC_145/Y INVX1_LOC_71/A 0.01fF
C71672 NAND2X1_LOC_198/B NOR2X1_LOC_123/B 0.20fF
C71673 NAND2X1_LOC_860/A INVX1_LOC_12/Y 0.04fF
C71674 INVX1_LOC_11/A NOR2X1_LOC_9/Y 0.61fF
C71675 INVX1_LOC_183/Y NOR2X1_LOC_91/Y 0.01fF
C71676 INVX1_LOC_145/A NOR2X1_LOC_355/A 0.11fF
C71677 NAND2X1_LOC_360/a_36_24# INVX1_LOC_46/A 0.01fF
C71678 NOR2X1_LOC_773/Y NAND2X1_LOC_477/A 0.10fF
C71679 NOR2X1_LOC_516/B NOR2X1_LOC_84/A 0.16fF
C71680 NOR2X1_LOC_843/A INVX1_LOC_22/A 0.17fF
C71681 NAND2X1_LOC_182/A NAND2X1_LOC_860/Y 0.01fF
C71682 INVX1_LOC_28/A INVX1_LOC_72/A 3.08fF
C71683 INVX1_LOC_237/Y NOR2X1_LOC_32/Y 0.00fF
C71684 NAND2X1_LOC_11/Y INVX1_LOC_191/Y 0.00fF
C71685 NAND2X1_LOC_84/Y INVX1_LOC_171/A 0.03fF
C71686 INVX1_LOC_239/A INVX1_LOC_11/Y 0.08fF
C71687 INVX1_LOC_298/A VDD 0.12fF
C71688 NOR2X1_LOC_716/B INVX1_LOC_10/A 0.02fF
C71689 NOR2X1_LOC_111/A NOR2X1_LOC_109/Y 3.82fF
C71690 D_INPUT_1 INVX1_LOC_9/A 0.10fF
C71691 NAND2X1_LOC_569/A INVX1_LOC_234/A 0.00fF
C71692 NOR2X1_LOC_84/B INVX1_LOC_3/Y 0.00fF
C71693 INVX1_LOC_256/A NOR2X1_LOC_191/a_36_216# 0.00fF
C71694 NOR2X1_LOC_321/Y NOR2X1_LOC_136/a_36_216# 0.00fF
C71695 NAND2X1_LOC_198/B INVX1_LOC_102/Y 0.10fF
C71696 D_INPUT_6 VDD 0.07fF
C71697 INVX1_LOC_121/A NOR2X1_LOC_377/Y 0.30fF
C71698 NOR2X1_LOC_208/Y NOR2X1_LOC_736/Y 0.01fF
C71699 NAND2X1_LOC_763/B NAND2X1_LOC_2/a_36_24# 0.01fF
C71700 NAND2X1_LOC_785/A NAND2X1_LOC_859/Y 0.00fF
C71701 INVX1_LOC_75/A NOR2X1_LOC_360/Y 0.10fF
C71702 NAND2X1_LOC_338/B INVX1_LOC_16/A 0.14fF
C71703 NOR2X1_LOC_173/Y VDD 0.24fF
C71704 NOR2X1_LOC_609/A NAND2X1_LOC_132/a_36_24# 0.00fF
C71705 NOR2X1_LOC_321/Y VDD 0.80fF
C71706 NOR2X1_LOC_526/Y INVX1_LOC_22/A 0.05fF
C71707 INVX1_LOC_14/A INVX1_LOC_20/A 1.47fF
C71708 NOR2X1_LOC_38/B INVX1_LOC_29/A 0.03fF
C71709 NOR2X1_LOC_593/Y NOR2X1_LOC_356/A 0.39fF
C71710 NOR2X1_LOC_437/Y INVX1_LOC_73/A 0.02fF
C71711 NAND2X1_LOC_182/A NAND2X1_LOC_861/Y 0.02fF
C71712 INVX1_LOC_1/A INVX1_LOC_46/A 0.35fF
C71713 INVX1_LOC_18/A INVX1_LOC_285/Y 0.00fF
C71714 NOR2X1_LOC_103/Y NAND2X1_LOC_465/A 0.02fF
C71715 INVX1_LOC_280/Y NOR2X1_LOC_690/Y 0.02fF
C71716 NAND2X1_LOC_364/A INVX1_LOC_6/A 0.03fF
C71717 NAND2X1_LOC_656/Y NOR2X1_LOC_172/a_36_216# 0.01fF
C71718 INVX1_LOC_58/A NAND2X1_LOC_240/a_36_24# 0.00fF
C71719 NOR2X1_LOC_401/B INVX1_LOC_164/A 0.05fF
C71720 NOR2X1_LOC_315/Y NOR2X1_LOC_72/a_36_216# 0.00fF
C71721 NAND2X1_LOC_722/A NOR2X1_LOC_576/B 0.07fF
C71722 INVX1_LOC_23/Y NAND2X1_LOC_773/B 1.45fF
C71723 INVX1_LOC_58/Y NOR2X1_LOC_445/B 0.02fF
C71724 NAND2X1_LOC_785/A NAND2X1_LOC_866/B 0.03fF
C71725 NOR2X1_LOC_433/A NOR2X1_LOC_74/A 0.01fF
C71726 VDD NAND2X1_LOC_793/Y 0.14fF
C71727 INVX1_LOC_256/A NOR2X1_LOC_266/B 0.02fF
C71728 NOR2X1_LOC_709/B NAND2X1_LOC_474/Y 0.03fF
C71729 INVX1_LOC_61/Y INVX1_LOC_59/Y 0.27fF
C71730 INVX1_LOC_33/A NOR2X1_LOC_336/a_36_216# 0.00fF
C71731 INVX1_LOC_234/A INVX1_LOC_316/Y 0.02fF
C71732 INVX1_LOC_290/A NOR2X1_LOC_583/a_36_216# 0.00fF
C71733 NOR2X1_LOC_593/Y NOR2X1_LOC_74/A 0.18fF
C71734 NAND2X1_LOC_859/Y NOR2X1_LOC_86/A 0.10fF
C71735 INVX1_LOC_229/A NOR2X1_LOC_536/A 0.09fF
C71736 NOR2X1_LOC_690/A INVX1_LOC_282/A 0.07fF
C71737 NOR2X1_LOC_387/A NOR2X1_LOC_387/Y 0.00fF
C71738 INVX1_LOC_90/A INVX1_LOC_144/Y -0.00fF
C71739 INVX1_LOC_136/A NOR2X1_LOC_675/A 0.01fF
C71740 INVX1_LOC_63/Y INVX1_LOC_144/A 0.10fF
C71741 NOR2X1_LOC_272/Y INVX1_LOC_131/Y 0.69fF
C71742 NOR2X1_LOC_804/B NOR2X1_LOC_552/Y 0.01fF
C71743 NOR2X1_LOC_123/B INVX1_LOC_53/Y 0.07fF
C71744 INVX1_LOC_206/Y INVX1_LOC_113/Y 0.00fF
C71745 NOR2X1_LOC_13/Y NOR2X1_LOC_45/B 0.51fF
C71746 NAND2X1_LOC_338/B INVX1_LOC_28/A 0.21fF
C71747 NOR2X1_LOC_514/A D_INPUT_3 0.20fF
C71748 NOR2X1_LOC_759/Y NOR2X1_LOC_139/Y 0.00fF
C71749 INVX1_LOC_21/A INVX1_LOC_179/A 0.03fF
C71750 INVX1_LOC_5/A NAND2X1_LOC_574/A 0.02fF
C71751 NOR2X1_LOC_596/Y NAND2X1_LOC_472/Y 0.01fF
C71752 INVX1_LOC_111/A NOR2X1_LOC_405/A 0.00fF
C71753 NAND2X1_LOC_112/Y NOR2X1_LOC_106/A 0.00fF
C71754 INVX1_LOC_202/A NOR2X1_LOC_139/Y 0.01fF
C71755 NOR2X1_LOC_52/B NOR2X1_LOC_74/A 0.14fF
C71756 INVX1_LOC_12/A NOR2X1_LOC_654/A 0.08fF
C71757 NOR2X1_LOC_340/A NOR2X1_LOC_105/Y 0.05fF
C71758 NOR2X1_LOC_448/Y NAND2X1_LOC_93/B 0.16fF
C71759 NOR2X1_LOC_637/A NOR2X1_LOC_56/Y 0.05fF
C71760 NOR2X1_LOC_241/A INVX1_LOC_9/A 0.03fF
C71761 INVX1_LOC_313/Y INVX1_LOC_16/A 0.03fF
C71762 NOR2X1_LOC_273/Y NAND2X1_LOC_468/B 0.00fF
C71763 NOR2X1_LOC_510/Y NOR2X1_LOC_127/a_36_216# 0.00fF
C71764 NOR2X1_LOC_766/a_36_216# NOR2X1_LOC_766/Y 0.01fF
C71765 INVX1_LOC_5/A INVX1_LOC_136/Y 0.00fF
C71766 NOR2X1_LOC_134/Y NOR2X1_LOC_536/A 0.02fF
C71767 INVX1_LOC_279/A NAND2X1_LOC_140/A 0.02fF
C71768 NOR2X1_LOC_577/Y NOR2X1_LOC_595/Y 0.01fF
C71769 NOR2X1_LOC_52/B NOR2X1_LOC_9/Y 0.08fF
C71770 INVX1_LOC_36/A NOR2X1_LOC_111/A 0.07fF
C71771 INVX1_LOC_32/A INVX1_LOC_16/Y 0.01fF
C71772 NOR2X1_LOC_415/A D_INPUT_0 0.01fF
C71773 NOR2X1_LOC_19/B INVX1_LOC_316/Y 1.30fF
C71774 INVX1_LOC_23/A INVX1_LOC_109/Y 0.07fF
C71775 INVX1_LOC_21/Y NAND2X1_LOC_175/Y 0.11fF
C71776 NOR2X1_LOC_448/Y NAND2X1_LOC_425/Y 0.03fF
C71777 NAND2X1_LOC_175/B NOR2X1_LOC_45/B 0.24fF
C71778 INVX1_LOC_202/A NAND2X1_LOC_468/B 0.02fF
C71779 NOR2X1_LOC_805/a_36_216# INVX1_LOC_307/Y 0.00fF
C71780 NOR2X1_LOC_500/A NOR2X1_LOC_324/B 0.19fF
C71781 INVX1_LOC_35/A INVX1_LOC_272/A 0.08fF
C71782 NAND2X1_LOC_739/B INVX1_LOC_20/A 0.03fF
C71783 NOR2X1_LOC_393/Y INVX1_LOC_23/Y 0.03fF
C71784 NOR2X1_LOC_826/a_36_216# INVX1_LOC_284/A 0.00fF
C71785 NOR2X1_LOC_658/Y INVX1_LOC_281/A 0.06fF
C71786 INVX1_LOC_211/Y INVX1_LOC_54/A 0.03fF
C71787 NAND2X1_LOC_84/Y INVX1_LOC_20/A 0.01fF
C71788 NOR2X1_LOC_78/B NOR2X1_LOC_188/A 0.03fF
C71789 NOR2X1_LOC_637/A VDD -0.00fF
C71790 INVX1_LOC_36/A NOR2X1_LOC_694/Y 0.22fF
C71791 INVX1_LOC_214/Y NOR2X1_LOC_815/A 0.00fF
C71792 NAND2X1_LOC_276/Y NAND2X1_LOC_642/Y 0.12fF
C71793 INVX1_LOC_68/Y NOR2X1_LOC_196/Y 0.09fF
C71794 INVX1_LOC_98/A NOR2X1_LOC_709/A 0.08fF
C71795 NOR2X1_LOC_824/A NOR2X1_LOC_662/A 0.03fF
C71796 INVX1_LOC_163/A INVX1_LOC_84/A 0.15fF
C71797 INVX1_LOC_32/A NAND2X1_LOC_205/A 0.01fF
C71798 INVX1_LOC_290/Y NOR2X1_LOC_678/A 0.00fF
C71799 GATE_811 INVX1_LOC_11/Y 0.00fF
C71800 INVX1_LOC_30/A NAND2X1_LOC_204/a_36_24# 0.00fF
C71801 NOR2X1_LOC_78/A NOR2X1_LOC_709/A 0.37fF
C71802 INVX1_LOC_11/A NOR2X1_LOC_865/Y 0.07fF
C71803 INVX1_LOC_239/A INVX1_LOC_203/A 0.01fF
C71804 NOR2X1_LOC_755/a_36_216# NAND2X1_LOC_656/Y -0.01fF
C71805 NAND2X1_LOC_550/A INVX1_LOC_35/Y 0.01fF
C71806 INVX1_LOC_24/A INVX1_LOC_33/Y 0.03fF
C71807 NOR2X1_LOC_299/Y INVX1_LOC_140/A 0.07fF
C71808 INVX1_LOC_11/A NOR2X1_LOC_243/B 0.07fF
C71809 NAND2X1_LOC_400/a_36_24# NAND2X1_LOC_99/A 0.00fF
C71810 INVX1_LOC_17/A NOR2X1_LOC_430/Y 0.03fF
C71811 NOR2X1_LOC_570/B NOR2X1_LOC_357/Y 0.01fF
C71812 NOR2X1_LOC_30/Y INVX1_LOC_296/A 0.18fF
C71813 NAND2X1_LOC_198/B NOR2X1_LOC_331/B 0.30fF
C71814 NOR2X1_LOC_301/A INVX1_LOC_181/A 0.16fF
C71815 NOR2X1_LOC_456/a_36_216# INVX1_LOC_29/A 0.00fF
C71816 NOR2X1_LOC_606/Y INVX1_LOC_46/Y 0.04fF
C71817 INVX1_LOC_28/A INVX1_LOC_313/Y 0.01fF
C71818 NOR2X1_LOC_299/Y NAND2X1_LOC_463/B 0.01fF
C71819 INVX1_LOC_7/Y INVX1_LOC_42/A 0.02fF
C71820 NOR2X1_LOC_788/B NOR2X1_LOC_703/A 0.02fF
C71821 NOR2X1_LOC_489/B INVX1_LOC_4/A 0.07fF
C71822 NAND2X1_LOC_660/A NAND2X1_LOC_655/B 0.08fF
C71823 NOR2X1_LOC_716/B NOR2X1_LOC_301/a_36_216# 0.01fF
C71824 NOR2X1_LOC_761/Y NAND2X1_LOC_810/B 0.05fF
C71825 NOR2X1_LOC_168/B NAND2X1_LOC_280/a_36_24# 0.00fF
C71826 INVX1_LOC_49/A NOR2X1_LOC_536/A 0.43fF
C71827 NOR2X1_LOC_527/Y NAND2X1_LOC_808/A 0.01fF
C71828 NOR2X1_LOC_468/Y INVX1_LOC_29/A 0.04fF
C71829 INVX1_LOC_83/A NOR2X1_LOC_188/A 0.01fF
C71830 INVX1_LOC_90/A NOR2X1_LOC_322/Y 0.83fF
C71831 NAND2X1_LOC_364/A INVX1_LOC_131/Y 0.19fF
C71832 INVX1_LOC_48/Y INVX1_LOC_284/A 0.76fF
C71833 NAND2X1_LOC_354/B NAND2X1_LOC_685/a_36_24# 0.00fF
C71834 NAND2X1_LOC_190/Y INVX1_LOC_29/A 0.26fF
C71835 NOR2X1_LOC_607/Y INVX1_LOC_9/A 0.02fF
C71836 NAND2X1_LOC_860/A NOR2X1_LOC_89/Y 0.06fF
C71837 NOR2X1_LOC_537/Y NOR2X1_LOC_35/Y 0.16fF
C71838 NAND2X1_LOC_338/B NOR2X1_LOC_35/Y 0.10fF
C71839 NOR2X1_LOC_34/B INVX1_LOC_15/A 0.02fF
C71840 INVX1_LOC_7/A INVX1_LOC_123/A 0.34fF
C71841 NAND2X1_LOC_270/a_36_24# NOR2X1_LOC_76/A 0.00fF
C71842 INVX1_LOC_14/A NOR2X1_LOC_128/A 0.04fF
C71843 NOR2X1_LOC_92/Y INVX1_LOC_42/A 0.22fF
C71844 INVX1_LOC_8/A NOR2X1_LOC_98/B 0.00fF
C71845 NOR2X1_LOC_543/A INVX1_LOC_91/A 0.04fF
C71846 NOR2X1_LOC_646/B NAND2X1_LOC_215/A 0.00fF
C71847 NOR2X1_LOC_392/Y INVX1_LOC_26/A 0.01fF
C71848 NOR2X1_LOC_246/A INVX1_LOC_286/A 0.01fF
C71849 INVX1_LOC_90/A INVX1_LOC_92/Y 0.01fF
C71850 INVX1_LOC_30/A NAND2X1_LOC_456/Y 0.04fF
C71851 NAND2X1_LOC_112/a_36_24# NOR2X1_LOC_111/A 0.00fF
C71852 INVX1_LOC_266/Y INVX1_LOC_117/A 0.03fF
C71853 NOR2X1_LOC_75/Y INVX1_LOC_12/A 0.02fF
C71854 INVX1_LOC_163/A INVX1_LOC_15/A 0.08fF
C71855 INVX1_LOC_154/A NOR2X1_LOC_349/B 0.35fF
C71856 NAND2X1_LOC_51/B NOR2X1_LOC_163/Y 0.02fF
C71857 INVX1_LOC_49/A NAND2X1_LOC_93/B 0.06fF
C71858 INVX1_LOC_245/Y NOR2X1_LOC_89/A 0.04fF
C71859 NOR2X1_LOC_389/A INVX1_LOC_29/A 0.12fF
C71860 NOR2X1_LOC_355/B NOR2X1_LOC_355/a_36_216# 0.00fF
C71861 INVX1_LOC_2/A NOR2X1_LOC_536/A 2.38fF
C71862 NOR2X1_LOC_723/Y INVX1_LOC_186/Y 0.02fF
C71863 NAND2X1_LOC_9/Y INVX1_LOC_25/A 0.05fF
C71864 NAND2X1_LOC_199/B INVX1_LOC_29/A 0.07fF
C71865 INVX1_LOC_49/A NAND2X1_LOC_425/Y 0.89fF
C71866 INVX1_LOC_30/A INVX1_LOC_49/Y 0.03fF
C71867 INVX1_LOC_300/A VDD 0.00fF
C71868 INVX1_LOC_90/A NOR2X1_LOC_562/B 0.66fF
C71869 NOR2X1_LOC_181/Y INVX1_LOC_274/A 0.22fF
C71870 INVX1_LOC_14/A INVX1_LOC_4/A 1.37fF
C71871 NOR2X1_LOC_82/Y NAND2X1_LOC_262/a_36_24# 0.00fF
C71872 INVX1_LOC_211/Y NOR2X1_LOC_48/B 0.17fF
C71873 NOR2X1_LOC_226/A NOR2X1_LOC_536/A 0.47fF
C71874 NOR2X1_LOC_798/A INVX1_LOC_116/Y 0.02fF
C71875 NAND2X1_LOC_479/Y INVX1_LOC_37/A 0.03fF
C71876 INVX1_LOC_155/A NOR2X1_LOC_216/B 0.03fF
C71877 NOR2X1_LOC_246/A INVX1_LOC_95/A 0.02fF
C71878 NOR2X1_LOC_91/A NAND2X1_LOC_740/Y 0.03fF
C71879 INVX1_LOC_136/A NAND2X1_LOC_500/B 0.01fF
C71880 INVX1_LOC_63/Y NOR2X1_LOC_155/A 0.03fF
C71881 NOR2X1_LOC_92/Y INVX1_LOC_78/A 0.30fF
C71882 NOR2X1_LOC_497/a_36_216# NAND2X1_LOC_35/Y 0.01fF
C71883 INVX1_LOC_138/Y NOR2X1_LOC_416/A 0.03fF
C71884 NOR2X1_LOC_653/B NAND2X1_LOC_286/B 0.01fF
C71885 INVX1_LOC_93/A NAND2X1_LOC_442/a_36_24# 0.01fF
C71886 NOR2X1_LOC_65/B INVX1_LOC_7/Y -0.00fF
C71887 INVX1_LOC_30/A INVX1_LOC_99/A 0.04fF
C71888 INVX1_LOC_33/A NOR2X1_LOC_461/B 0.01fF
C71889 NAND2X1_LOC_214/B INVX1_LOC_57/A 0.07fF
C71890 NOR2X1_LOC_686/B VDD -0.00fF
C71891 INVX1_LOC_107/A INVX1_LOC_29/A 0.01fF
C71892 NOR2X1_LOC_400/B INVX1_LOC_235/Y 0.01fF
C71893 INVX1_LOC_17/A INVX1_LOC_94/Y 1.78fF
C71894 NAND2X1_LOC_325/Y INVX1_LOC_285/A 0.01fF
C71895 INVX1_LOC_2/A NAND2X1_LOC_93/B 0.06fF
C71896 NOR2X1_LOC_2/Y NOR2X1_LOC_587/a_36_216# 0.00fF
C71897 INVX1_LOC_75/A NOR2X1_LOC_269/Y 0.10fF
C71898 INVX1_LOC_62/Y INVX1_LOC_29/A 0.01fF
C71899 INVX1_LOC_298/Y NAND2X1_LOC_190/Y 0.07fF
C71900 NOR2X1_LOC_312/Y NAND2X1_LOC_287/B 0.23fF
C71901 INVX1_LOC_27/A INVX1_LOC_57/A 0.15fF
C71902 NAND2X1_LOC_30/Y NAND2X1_LOC_470/B 0.10fF
C71903 INVX1_LOC_135/A INVX1_LOC_37/A 4.60fF
C71904 NOR2X1_LOC_91/A NAND2X1_LOC_706/Y 0.07fF
C71905 INVX1_LOC_313/Y NOR2X1_LOC_35/Y 0.10fF
C71906 NOR2X1_LOC_65/B NOR2X1_LOC_92/Y 0.15fF
C71907 NOR2X1_LOC_824/A INVX1_LOC_57/A 0.07fF
C71908 NAND2X1_LOC_68/a_36_24# INVX1_LOC_50/A 0.00fF
C71909 NOR2X1_LOC_553/Y INVX1_LOC_9/A 0.05fF
C71910 NOR2X1_LOC_226/A NAND2X1_LOC_93/B 0.07fF
C71911 NAND2X1_LOC_214/B NAND2X1_LOC_541/a_36_24# 0.01fF
C71912 INVX1_LOC_34/A NAND2X1_LOC_475/Y 0.13fF
C71913 NAND2X1_LOC_783/A INVX1_LOC_33/Y 0.14fF
C71914 INVX1_LOC_295/A INVX1_LOC_37/A 0.08fF
C71915 INVX1_LOC_57/Y INVX1_LOC_19/Y 0.41fF
C71916 NOR2X1_LOC_665/A NOR2X1_LOC_331/B 0.51fF
C71917 NAND2X1_LOC_35/Y INVX1_LOC_5/A 0.03fF
C71918 INVX1_LOC_33/Y NOR2X1_LOC_130/A 0.03fF
C71919 NOR2X1_LOC_614/Y NOR2X1_LOC_640/Y 0.03fF
C71920 INVX1_LOC_132/A INVX1_LOC_125/A 0.01fF
C71921 NOR2X1_LOC_717/Y INVX1_LOC_4/A 0.07fF
C71922 INVX1_LOC_11/A NAND2X1_LOC_425/a_36_24# 0.00fF
C71923 NAND2X1_LOC_116/A NAND2X1_LOC_206/Y 0.18fF
C71924 INVX1_LOC_143/A NAND2X1_LOC_52/a_36_24# 0.00fF
C71925 NOR2X1_LOC_121/A NOR2X1_LOC_99/Y 0.04fF
C71926 NAND2X1_LOC_837/Y INVX1_LOC_42/A 0.14fF
C71927 INVX1_LOC_148/A VDD 0.24fF
C71928 NOR2X1_LOC_113/A INVX1_LOC_6/A 0.01fF
C71929 NOR2X1_LOC_161/Y NAND2X1_LOC_93/B 0.02fF
C71930 INVX1_LOC_10/A NOR2X1_LOC_709/B 0.00fF
C71931 INVX1_LOC_72/Y INVX1_LOC_3/Y 0.02fF
C71932 INVX1_LOC_17/A INVX1_LOC_296/A 0.07fF
C71933 INVX1_LOC_50/A INVX1_LOC_103/A 0.12fF
C71934 NOR2X1_LOC_818/Y NOR2X1_LOC_649/B 0.02fF
C71935 INVX1_LOC_16/A NOR2X1_LOC_79/a_36_216# 0.00fF
C71936 INVX1_LOC_2/A INVX1_LOC_3/A 0.48fF
C71937 NOR2X1_LOC_405/A INVX1_LOC_6/A 0.07fF
C71938 NOR2X1_LOC_716/B INVX1_LOC_12/A 0.46fF
C71939 NAND2X1_LOC_35/Y INVX1_LOC_178/A 0.10fF
C71940 INVX1_LOC_240/A INVX1_LOC_240/Y 0.01fF
C71941 NAND2X1_LOC_9/Y INVX1_LOC_1/A 0.01fF
C71942 NOR2X1_LOC_161/Y NAND2X1_LOC_425/Y 0.06fF
C71943 INPUT_1 NOR2X1_LOC_536/A 0.06fF
C71944 INVX1_LOC_35/A INVX1_LOC_198/A 0.01fF
C71945 NOR2X1_LOC_295/Y INVX1_LOC_29/A 0.12fF
C71946 NOR2X1_LOC_412/a_36_216# INVX1_LOC_284/A 0.00fF
C71947 INVX1_LOC_18/A INVX1_LOC_4/Y 0.07fF
C71948 INVX1_LOC_233/A INVX1_LOC_1/A 0.10fF
C71949 INVX1_LOC_5/A NAND2X1_LOC_571/Y 0.10fF
C71950 INVX1_LOC_174/A NOR2X1_LOC_383/B 0.08fF
C71951 NAND2X1_LOC_860/A NOR2X1_LOC_401/A 0.05fF
C71952 NOR2X1_LOC_844/A INVX1_LOC_29/A 0.03fF
C71953 NOR2X1_LOC_246/A INVX1_LOC_54/A 0.03fF
C71954 INVX1_LOC_41/A INVX1_LOC_42/A 0.03fF
C71955 INVX1_LOC_90/A INVX1_LOC_193/A 0.57fF
C71956 INVX1_LOC_50/A INVX1_LOC_292/A 0.16fF
C71957 INVX1_LOC_64/A INVX1_LOC_14/A 0.02fF
C71958 INVX1_LOC_58/A INVX1_LOC_225/Y 0.25fF
C71959 NOR2X1_LOC_438/a_36_216# NAND2X1_LOC_793/B 0.01fF
C71960 NAND2X1_LOC_84/Y INVX1_LOC_4/A 0.04fF
C71961 NOR2X1_LOC_188/A INVX1_LOC_46/A 0.14fF
C71962 NOR2X1_LOC_510/Y NOR2X1_LOC_173/Y 0.01fF
C71963 NOR2X1_LOC_192/A INVX1_LOC_93/Y 0.03fF
C71964 INVX1_LOC_48/A INVX1_LOC_20/A 0.07fF
C71965 NOR2X1_LOC_717/B INVX1_LOC_307/A 0.15fF
C71966 INVX1_LOC_27/A INVX1_LOC_252/A 0.05fF
C71967 INVX1_LOC_11/A NOR2X1_LOC_342/A 0.00fF
C71968 NAND2X1_LOC_860/A NAND2X1_LOC_550/A 0.10fF
C71969 INVX1_LOC_123/A INVX1_LOC_76/A 0.03fF
C71970 NAND2X1_LOC_860/A NOR2X1_LOC_160/B 0.18fF
C71971 NOR2X1_LOC_690/A NOR2X1_LOC_496/a_36_216# 0.01fF
C71972 NOR2X1_LOC_84/Y INVX1_LOC_284/A 0.17fF
C71973 NAND2X1_LOC_325/a_36_24# NAND2X1_LOC_721/A 0.00fF
C71974 NOR2X1_LOC_589/A NOR2X1_LOC_127/Y 0.07fF
C71975 INVX1_LOC_35/A INVX1_LOC_150/Y 0.02fF
C71976 NOR2X1_LOC_322/Y INVX1_LOC_38/A 0.15fF
C71977 NAND2X1_LOC_198/B NOR2X1_LOC_449/A 0.00fF
C71978 NOR2X1_LOC_798/A INVX1_LOC_1/A 0.03fF
C71979 INPUT_1 NAND2X1_LOC_93/B 0.14fF
C71980 NOR2X1_LOC_160/B NOR2X1_LOC_634/Y 0.03fF
C71981 INVX1_LOC_298/Y NOR2X1_LOC_596/A 8.99fF
C71982 NOR2X1_LOC_186/Y NAND2X1_LOC_538/Y 0.07fF
C71983 NOR2X1_LOC_220/A INVX1_LOC_29/A 0.01fF
C71984 INVX1_LOC_190/Y NAND2X1_LOC_798/B 0.01fF
C71985 NOR2X1_LOC_828/A INVX1_LOC_307/A 0.19fF
C71986 INVX1_LOC_49/A NAND2X1_LOC_470/B 0.11fF
C71987 NAND2X1_LOC_124/a_36_24# NOR2X1_LOC_331/B 0.00fF
C71988 INVX1_LOC_24/A INVX1_LOC_23/Y 0.11fF
C71989 NOR2X1_LOC_757/Y INVX1_LOC_12/A 0.05fF
C71990 NAND2X1_LOC_72/Y INVX1_LOC_292/A 0.13fF
C71991 NAND2X1_LOC_364/A INVX1_LOC_270/A 0.03fF
C71992 INVX1_LOC_8/A NOR2X1_LOC_38/B 0.19fF
C71993 NAND2X1_LOC_399/a_36_24# NOR2X1_LOC_38/B 0.00fF
C71994 NAND2X1_LOC_390/A INVX1_LOC_19/A 1.20fF
C71995 INVX1_LOC_104/A NOR2X1_LOC_609/Y 0.04fF
C71996 INVX1_LOC_234/A NOR2X1_LOC_662/A 0.07fF
C71997 INVX1_LOC_41/A INVX1_LOC_78/A 0.06fF
C71998 NOR2X1_LOC_197/A INVX1_LOC_50/Y 0.48fF
C71999 INVX1_LOC_186/A NAND2X1_LOC_472/Y 0.07fF
C72000 NOR2X1_LOC_361/B NOR2X1_LOC_321/Y 0.06fF
C72001 NOR2X1_LOC_552/A INVX1_LOC_37/A 0.08fF
C72002 NOR2X1_LOC_320/Y INVX1_LOC_54/A 0.04fF
C72003 NOR2X1_LOC_620/Y INVX1_LOC_26/Y 0.02fF
C72004 INPUT_1 NOR2X1_LOC_649/B 1.55fF
C72005 INVX1_LOC_16/A NOR2X1_LOC_226/Y 0.00fF
C72006 INPUT_1 INVX1_LOC_3/A 1.05fF
C72007 NOR2X1_LOC_583/a_36_216# INVX1_LOC_261/Y 0.00fF
C72008 INVX1_LOC_111/Y INVX1_LOC_4/A 0.02fF
C72009 INVX1_LOC_17/A INVX1_LOC_299/A 0.07fF
C72010 NOR2X1_LOC_791/Y NAND2X1_LOC_208/B 0.01fF
C72011 INVX1_LOC_233/Y INVX1_LOC_18/A 0.01fF
C72012 NAND2X1_LOC_477/A INVX1_LOC_78/A 0.03fF
C72013 NOR2X1_LOC_92/Y NOR2X1_LOC_503/Y 0.30fF
C72014 INVX1_LOC_41/A NOR2X1_LOC_65/B 0.11fF
C72015 INVX1_LOC_2/A NAND2X1_LOC_470/B 2.40fF
C72016 NOR2X1_LOC_843/A NOR2X1_LOC_843/B 0.03fF
C72017 INVX1_LOC_311/A INVX1_LOC_179/A 0.95fF
C72018 INVX1_LOC_50/A INVX1_LOC_67/A 0.70fF
C72019 NOR2X1_LOC_749/a_36_216# NAND2X1_LOC_63/Y 0.00fF
C72020 INVX1_LOC_205/Y NAND2X1_LOC_555/Y 0.21fF
C72021 INVX1_LOC_21/A NOR2X1_LOC_641/B 0.00fF
C72022 NOR2X1_LOC_486/Y INVX1_LOC_44/A 0.08fF
C72023 NAND2X1_LOC_739/B INVX1_LOC_64/A 0.08fF
C72024 INVX1_LOC_22/A D_INPUT_5 0.01fF
C72025 INVX1_LOC_103/A NAND2X1_LOC_227/Y 0.00fF
C72026 INVX1_LOC_122/Y INVX1_LOC_50/Y 0.22fF
C72027 NOR2X1_LOC_272/Y INVX1_LOC_36/A 0.17fF
C72028 D_INPUT_0 NOR2X1_LOC_89/A 0.09fF
C72029 NAND2X1_LOC_794/B INVX1_LOC_72/A 0.68fF
C72030 INVX1_LOC_14/A INVX1_LOC_43/Y 0.03fF
C72031 NOR2X1_LOC_19/B NOR2X1_LOC_662/A 0.01fF
C72032 NOR2X1_LOC_405/a_36_216# INVX1_LOC_78/A 0.02fF
C72033 NOR2X1_LOC_299/Y INVX1_LOC_42/A 0.50fF
C72034 INVX1_LOC_77/A NOR2X1_LOC_678/A 0.10fF
C72035 NOR2X1_LOC_706/Y NAND2X1_LOC_425/Y 0.03fF
C72036 INVX1_LOC_45/A NAND2X1_LOC_149/Y 2.01fF
C72037 INVX1_LOC_215/A INVX1_LOC_32/A 0.01fF
C72038 NOR2X1_LOC_445/Y INVX1_LOC_23/A 0.03fF
C72039 NOR2X1_LOC_246/A NAND2X1_LOC_807/B 0.07fF
C72040 INVX1_LOC_21/A NOR2X1_LOC_751/Y 0.35fF
C72041 NOR2X1_LOC_65/B NAND2X1_LOC_477/A 0.01fF
C72042 INVX1_LOC_245/Y INVX1_LOC_11/A 0.04fF
C72043 INVX1_LOC_90/A INVX1_LOC_106/A 0.01fF
C72044 INVX1_LOC_50/A INVX1_LOC_240/A 0.05fF
C72045 INVX1_LOC_58/A NAND2X1_LOC_811/Y 0.04fF
C72046 NAND2X1_LOC_633/Y NOR2X1_LOC_301/a_36_216# 0.00fF
C72047 NOR2X1_LOC_750/Y NAND2X1_LOC_276/Y 0.01fF
C72048 NOR2X1_LOC_711/Y NOR2X1_LOC_209/B 0.05fF
C72049 NOR2X1_LOC_817/Y INPUT_3 0.17fF
C72050 NOR2X1_LOC_598/B INVX1_LOC_63/Y 0.18fF
C72051 NOR2X1_LOC_78/A NOR2X1_LOC_830/a_36_216# 0.00fF
C72052 INVX1_LOC_34/A NAND2X1_LOC_787/A 0.03fF
C72053 NOR2X1_LOC_211/A INVX1_LOC_78/A 0.03fF
C72054 NOR2X1_LOC_152/A INVX1_LOC_37/A 0.09fF
C72055 INVX1_LOC_211/Y NAND2X1_LOC_350/A 0.11fF
C72056 NAND2X1_LOC_112/Y NOR2X1_LOC_334/Y 0.15fF
C72057 INVX1_LOC_314/Y INVX1_LOC_306/Y 0.16fF
C72058 NOR2X1_LOC_332/a_36_216# INVX1_LOC_280/A 0.00fF
C72059 NOR2X1_LOC_405/A INVX1_LOC_131/Y 0.03fF
C72060 INVX1_LOC_21/A INVX1_LOC_45/Y 0.45fF
C72061 INVX1_LOC_206/A INVX1_LOC_57/A 0.01fF
C72062 NAND2X1_LOC_853/Y NOR2X1_LOC_829/A 0.03fF
C72063 NOR2X1_LOC_254/A NOR2X1_LOC_483/B 0.26fF
C72064 INVX1_LOC_58/A INVX1_LOC_266/Y 0.00fF
C72065 INVX1_LOC_64/A INVX1_LOC_217/Y 0.77fF
C72066 INVX1_LOC_17/A NOR2X1_LOC_524/Y 0.01fF
C72067 NOR2X1_LOC_690/A NAND2X1_LOC_624/B 0.02fF
C72068 INVX1_LOC_25/Y INVX1_LOC_26/A 0.03fF
C72069 NAND2X1_LOC_45/Y INVX1_LOC_15/A 0.00fF
C72070 NOR2X1_LOC_413/Y NAND2X1_LOC_624/B 0.04fF
C72071 NAND2X1_LOC_724/Y INVX1_LOC_280/Y 0.06fF
C72072 NAND2X1_LOC_565/B INVX1_LOC_23/Y 0.03fF
C72073 NOR2X1_LOC_357/Y INVX1_LOC_54/A 0.07fF
C72074 NOR2X1_LOC_45/B NOR2X1_LOC_697/Y 0.03fF
C72075 INVX1_LOC_269/A NOR2X1_LOC_68/A 0.19fF
C72076 NOR2X1_LOC_56/Y NAND2X1_LOC_798/B 1.57fF
C72077 NAND2X1_LOC_149/Y INVX1_LOC_71/A 0.07fF
C72078 INVX1_LOC_121/A INVX1_LOC_78/A 0.02fF
C72079 NAND2X1_LOC_200/B INVX1_LOC_57/A 0.09fF
C72080 INVX1_LOC_213/Y INVX1_LOC_213/A 0.04fF
C72081 INVX1_LOC_11/A NOR2X1_LOC_791/A 0.01fF
C72082 NOR2X1_LOC_82/A NOR2X1_LOC_791/B 0.03fF
C72083 NOR2X1_LOC_92/Y NOR2X1_LOC_152/Y 0.07fF
C72084 INVX1_LOC_51/Y INVX1_LOC_29/A 0.00fF
C72085 VDD NOR2X1_LOC_433/Y 0.13fF
C72086 NOR2X1_LOC_32/B NAND2X1_LOC_549/B 0.05fF
C72087 NAND2X1_LOC_639/A INVX1_LOC_118/A 0.02fF
C72088 NAND2X1_LOC_78/a_36_24# INVX1_LOC_54/Y 0.00fF
C72089 NAND2X1_LOC_785/A NOR2X1_LOC_109/Y 0.01fF
C72090 INVX1_LOC_88/A NOR2X1_LOC_759/Y 0.00fF
C72091 NOR2X1_LOC_242/A NOR2X1_LOC_285/B 0.02fF
C72092 INVX1_LOC_224/Y INVX1_LOC_16/A 0.10fF
C72093 INVX1_LOC_249/A NOR2X1_LOC_666/Y 0.11fF
C72094 INVX1_LOC_202/A INVX1_LOC_88/A 0.01fF
C72095 NOR2X1_LOC_255/Y INVX1_LOC_25/Y 0.20fF
C72096 VDD NAND2X1_LOC_798/B 0.01fF
C72097 NOR2X1_LOC_689/A INVX1_LOC_229/Y 0.06fF
C72098 INVX1_LOC_38/A INVX1_LOC_193/A 0.04fF
C72099 NOR2X1_LOC_536/A INVX1_LOC_118/A 0.21fF
C72100 INVX1_LOC_1/Y INVX1_LOC_29/Y 0.04fF
C72101 NOR2X1_LOC_272/Y NOR2X1_LOC_309/Y 0.03fF
C72102 INVX1_LOC_13/A NAND2X1_LOC_215/A 0.03fF
C72103 INVX1_LOC_66/Y INVX1_LOC_54/A 0.08fF
C72104 NOR2X1_LOC_130/A INVX1_LOC_23/Y 0.03fF
C72105 INVX1_LOC_6/A INVX1_LOC_109/Y 0.15fF
C72106 INVX1_LOC_100/Y INVX1_LOC_29/A 0.01fF
C72107 INVX1_LOC_36/A NOR2X1_LOC_761/Y 0.03fF
C72108 NOR2X1_LOC_692/Y INVX1_LOC_54/A 0.02fF
C72109 NAND2X1_LOC_568/A NOR2X1_LOC_152/Y 0.01fF
C72110 NAND2X1_LOC_571/Y NAND2X1_LOC_562/B 0.02fF
C72111 D_INPUT_7 NAND2X1_LOC_36/A 0.06fF
C72112 INVX1_LOC_234/A INVX1_LOC_57/A 0.01fF
C72113 INVX1_LOC_103/A NOR2X1_LOC_679/B 0.01fF
C72114 INVX1_LOC_291/Y INVX1_LOC_264/A 0.09fF
C72115 NOR2X1_LOC_468/Y INVX1_LOC_8/A 0.07fF
C72116 D_INPUT_1 NOR2X1_LOC_561/Y 0.07fF
C72117 NOR2X1_LOC_807/B INVX1_LOC_49/A 0.48fF
C72118 NOR2X1_LOC_99/B NOR2X1_LOC_646/B 0.15fF
C72119 NAND2X1_LOC_808/A NOR2X1_LOC_654/A 0.50fF
C72120 NOR2X1_LOC_71/Y NAND2X1_LOC_97/a_36_24# 0.01fF
C72121 INVX1_LOC_256/A INVX1_LOC_49/A 0.01fF
C72122 NAND2X1_LOC_738/B INVX1_LOC_229/Y 0.27fF
C72123 INVX1_LOC_200/A NOR2X1_LOC_716/B 0.15fF
C72124 D_INPUT_1 INVX1_LOC_7/A 0.47fF
C72125 NAND2X1_LOC_462/B NOR2X1_LOC_476/B 0.03fF
C72126 INVX1_LOC_36/A NAND2X1_LOC_364/A 0.03fF
C72127 INVX1_LOC_110/Y NOR2X1_LOC_860/B 0.37fF
C72128 NOR2X1_LOC_763/Y NOR2X1_LOC_452/A 0.03fF
C72129 INVX1_LOC_21/A NOR2X1_LOC_190/a_36_216# 0.02fF
C72130 NOR2X1_LOC_91/A NOR2X1_LOC_597/A 0.05fF
C72131 INVX1_LOC_45/A NOR2X1_LOC_744/Y 0.00fF
C72132 INVX1_LOC_286/A INVX1_LOC_32/A 0.18fF
C72133 NAND2X1_LOC_468/B NAND2X1_LOC_74/B 0.03fF
C72134 NOR2X1_LOC_212/a_36_216# INVX1_LOC_22/A 0.00fF
C72135 NAND2X1_LOC_741/B INVX1_LOC_24/A 0.03fF
C72136 INVX1_LOC_254/Y INVX1_LOC_31/A 0.09fF
C72137 NOR2X1_LOC_548/A INVX1_LOC_4/Y 0.01fF
C72138 NOR2X1_LOC_82/A NOR2X1_LOC_124/B 0.04fF
C72139 NOR2X1_LOC_266/a_36_216# INVX1_LOC_181/Y -0.01fF
C72140 NAND2X1_LOC_469/B INVX1_LOC_29/A 0.03fF
C72141 INVX1_LOC_48/A INVX1_LOC_4/A 0.42fF
C72142 NOR2X1_LOC_111/A INVX1_LOC_63/A 0.09fF
C72143 INVX1_LOC_17/A NOR2X1_LOC_315/Y 0.03fF
C72144 NOR2X1_LOC_542/Y INVX1_LOC_23/A 0.05fF
C72145 NOR2X1_LOC_78/B NAND2X1_LOC_326/A 0.00fF
C72146 NOR2X1_LOC_250/Y NOR2X1_LOC_52/B -0.00fF
C72147 INVX1_LOC_124/Y NOR2X1_LOC_433/A 0.01fF
C72148 INVX1_LOC_75/A INVX1_LOC_26/A 0.03fF
C72149 NOR2X1_LOC_772/A INVX1_LOC_57/A 0.00fF
C72150 INVX1_LOC_25/A NAND2X1_LOC_842/B 0.02fF
C72151 INVX1_LOC_21/A INVX1_LOC_255/Y 0.07fF
C72152 INVX1_LOC_232/Y NOR2X1_LOC_381/Y 0.04fF
C72153 NOR2X1_LOC_857/A NOR2X1_LOC_633/A 0.03fF
C72154 NOR2X1_LOC_640/Y NOR2X1_LOC_862/B 0.19fF
C72155 NOR2X1_LOC_19/B INVX1_LOC_57/A 0.03fF
C72156 INVX1_LOC_14/A NAND2X1_LOC_850/Y 0.19fF
C72157 NOR2X1_LOC_516/B NAND2X1_LOC_473/A 0.13fF
C72158 INVX1_LOC_311/Y INVX1_LOC_23/A 0.13fF
C72159 NOR2X1_LOC_189/A INVX1_LOC_72/A 0.12fF
C72160 NOR2X1_LOC_561/Y NOR2X1_LOC_652/Y 0.10fF
C72161 NAND2X1_LOC_785/B NAND2X1_LOC_833/Y 0.44fF
C72162 INVX1_LOC_305/A INVX1_LOC_77/A 0.07fF
C72163 INVX1_LOC_19/A INVX1_LOC_117/A 9.34fF
C72164 INVX1_LOC_2/A INVX1_LOC_256/A 0.13fF
C72165 NOR2X1_LOC_92/Y NAND2X1_LOC_859/B 0.11fF
C72166 INVX1_LOC_95/A INVX1_LOC_32/A 0.01fF
C72167 INVX1_LOC_212/Y NAND2X1_LOC_510/A 0.11fF
C72168 INVX1_LOC_276/A NAND2X1_LOC_803/B 0.39fF
C72169 INVX1_LOC_34/A INVX1_LOC_30/A 0.29fF
C72170 INVX1_LOC_118/A INVX1_LOC_3/A 0.03fF
C72171 NOR2X1_LOC_78/A NOR2X1_LOC_334/Y 0.14fF
C72172 INVX1_LOC_28/A NAND2X1_LOC_793/B 0.07fF
C72173 NOR2X1_LOC_360/Y NOR2X1_LOC_577/Y 0.10fF
C72174 INVX1_LOC_256/A NOR2X1_LOC_226/A 0.02fF
C72175 INVX1_LOC_118/A NOR2X1_LOC_661/A 0.01fF
C72176 NOR2X1_LOC_255/Y INVX1_LOC_75/A 0.01fF
C72177 NOR2X1_LOC_186/Y NOR2X1_LOC_106/A 0.00fF
C72178 NAND2X1_LOC_572/B INVX1_LOC_92/A 0.02fF
C72179 INVX1_LOC_298/Y NAND2X1_LOC_498/a_36_24# 0.01fF
C72180 NAND2X1_LOC_63/Y NOR2X1_LOC_536/A 0.04fF
C72181 INVX1_LOC_276/A NOR2X1_LOC_590/A 0.07fF
C72182 NOR2X1_LOC_552/A NAND2X1_LOC_72/B 0.33fF
C72183 INVX1_LOC_21/A NOR2X1_LOC_71/Y 0.05fF
C72184 NOR2X1_LOC_335/B INVX1_LOC_23/A 0.02fF
C72185 NOR2X1_LOC_67/A NOR2X1_LOC_590/A 0.05fF
C72186 NOR2X1_LOC_103/Y INVX1_LOC_16/A 0.11fF
C72187 NOR2X1_LOC_382/Y NAND2X1_LOC_141/A 0.05fF
C72188 INVX1_LOC_256/A NOR2X1_LOC_218/Y 0.02fF
C72189 NAND2X1_LOC_364/A NOR2X1_LOC_309/Y 0.18fF
C72190 NAND2X1_LOC_848/A NOR2X1_LOC_89/A 0.12fF
C72191 NAND2X1_LOC_454/Y NOR2X1_LOC_275/A 0.02fF
C72192 INVX1_LOC_62/Y INVX1_LOC_8/A 0.02fF
C72193 INVX1_LOC_58/A INVX1_LOC_191/A 0.40fF
C72194 NAND2X1_LOC_326/A INVX1_LOC_83/A 0.04fF
C72195 NOR2X1_LOC_335/A INVX1_LOC_77/A 0.01fF
C72196 VDD INVX1_LOC_47/Y 1.15fF
C72197 NAND2X1_LOC_9/Y NOR2X1_LOC_188/A 0.07fF
C72198 NAND2X1_LOC_218/a_36_24# INVX1_LOC_315/Y 0.00fF
C72199 NAND2X1_LOC_231/Y INVX1_LOC_30/A 0.19fF
C72200 INVX1_LOC_11/A NAND2X1_LOC_660/Y 0.10fF
C72201 NOR2X1_LOC_815/A INVX1_LOC_53/A 0.01fF
C72202 INVX1_LOC_21/A NOR2X1_LOC_644/A 0.03fF
C72203 NAND2X1_LOC_363/B INPUT_0 0.09fF
C72204 NAND2X1_LOC_740/B NOR2X1_LOC_304/Y 0.02fF
C72205 NOR2X1_LOC_690/A NOR2X1_LOC_617/Y 0.33fF
C72206 NOR2X1_LOC_435/a_36_216# INVX1_LOC_144/A 0.01fF
C72207 NAND2X1_LOC_9/Y NOR2X1_LOC_548/B 0.04fF
C72208 NOR2X1_LOC_48/B NOR2X1_LOC_692/Y 0.03fF
C72209 NOR2X1_LOC_528/Y INVX1_LOC_57/A 0.58fF
C72210 NOR2X1_LOC_413/Y NOR2X1_LOC_617/Y 0.10fF
C72211 NOR2X1_LOC_669/a_36_216# INVX1_LOC_90/A 0.00fF
C72212 INVX1_LOC_58/A INVX1_LOC_125/Y 0.09fF
C72213 NAND2X1_LOC_63/Y NAND2X1_LOC_93/B 0.03fF
C72214 NOR2X1_LOC_19/B INVX1_LOC_252/A 0.02fF
C72215 NOR2X1_LOC_113/A INVX1_LOC_270/A 0.26fF
C72216 NOR2X1_LOC_328/Y INVX1_LOC_286/Y 0.09fF
C72217 INVX1_LOC_13/A INVX1_LOC_218/Y 0.01fF
C72218 NOR2X1_LOC_318/B INVX1_LOC_29/Y 0.07fF
C72219 NOR2X1_LOC_607/A INVX1_LOC_177/A 0.00fF
C72220 NOR2X1_LOC_405/A INVX1_LOC_270/A 2.87fF
C72221 NOR2X1_LOC_496/Y NAND2X1_LOC_560/A 0.08fF
C72222 INVX1_LOC_30/A NAND2X1_LOC_858/a_36_24# 0.00fF
C72223 INVX1_LOC_11/A D_INPUT_0 0.53fF
C72224 NAND2X1_LOC_7/Y NOR2X1_LOC_6/B 0.07fF
C72225 NOR2X1_LOC_520/B NAND2X1_LOC_518/a_36_24# 0.02fF
C72226 INVX1_LOC_1/A NAND2X1_LOC_842/B 0.03fF
C72227 INVX1_LOC_45/A INVX1_LOC_16/A 0.09fF
C72228 NOR2X1_LOC_794/a_36_216# INVX1_LOC_104/A -0.02fF
C72229 NAND2X1_LOC_477/A NOR2X1_LOC_152/Y 0.07fF
C72230 NAND2X1_LOC_30/Y NOR2X1_LOC_764/Y 0.06fF
C72231 NAND2X1_LOC_325/Y NAND2X1_LOC_354/B 0.02fF
C72232 NAND2X1_LOC_563/A NOR2X1_LOC_68/A 0.02fF
C72233 NOR2X1_LOC_791/Y INPUT_0 1.63fF
C72234 NOR2X1_LOC_19/B NOR2X1_LOC_475/A 0.01fF
C72235 INVX1_LOC_230/Y NOR2X1_LOC_719/a_36_216# 0.01fF
C72236 INVX1_LOC_93/Y INVX1_LOC_29/Y 0.16fF
C72237 NAND2X1_LOC_856/A INVX1_LOC_16/A 0.03fF
C72238 NOR2X1_LOC_798/A NOR2X1_LOC_188/A 0.03fF
C72239 NOR2X1_LOC_61/Y NOR2X1_LOC_861/Y 0.17fF
C72240 INVX1_LOC_124/A NOR2X1_LOC_335/A 0.01fF
C72241 INVX1_LOC_304/Y NOR2X1_LOC_716/B 0.98fF
C72242 NAND2X1_LOC_477/Y NOR2X1_LOC_662/A 0.10fF
C72243 NOR2X1_LOC_451/A NOR2X1_LOC_48/B 0.04fF
C72244 INVX1_LOC_132/A NOR2X1_LOC_709/A 0.11fF
C72245 NOR2X1_LOC_383/B INVX1_LOC_20/A 0.03fF
C72246 NOR2X1_LOC_798/A NOR2X1_LOC_548/B 0.05fF
C72247 INVX1_LOC_290/A INVX1_LOC_72/A 0.21fF
C72248 INVX1_LOC_50/A NAND2X1_LOC_440/a_36_24# 0.01fF
C72249 INVX1_LOC_256/A INPUT_1 0.02fF
C72250 INVX1_LOC_32/A INVX1_LOC_54/A 0.03fF
C72251 INVX1_LOC_83/A NAND2X1_LOC_104/a_36_24# 0.01fF
C72252 NOR2X1_LOC_389/A NAND2X1_LOC_140/A 0.04fF
C72253 NAND2X1_LOC_338/B NOR2X1_LOC_350/A 0.04fF
C72254 NOR2X1_LOC_360/Y INVX1_LOC_22/A 0.72fF
C72255 INVX1_LOC_230/Y INVX1_LOC_89/A 0.17fF
C72256 INVX1_LOC_103/A NAND2X1_LOC_652/Y 0.03fF
C72257 NAND2X1_LOC_724/A NAND2X1_LOC_863/A 0.46fF
C72258 INVX1_LOC_28/A NOR2X1_LOC_103/Y 0.02fF
C72259 NOR2X1_LOC_160/B INVX1_LOC_85/Y 0.03fF
C72260 INVX1_LOC_5/A NOR2X1_LOC_845/A 0.02fF
C72261 INVX1_LOC_277/A INVX1_LOC_83/A 0.03fF
C72262 NOR2X1_LOC_246/A NOR2X1_LOC_441/Y 0.64fF
C72263 NAND2X1_LOC_738/B INVX1_LOC_20/A 0.03fF
C72264 INVX1_LOC_257/A NAND2X1_LOC_93/B 0.03fF
C72265 INVX1_LOC_50/A NOR2X1_LOC_137/Y 0.05fF
C72266 INVX1_LOC_24/A INVX1_LOC_232/A 0.10fF
C72267 INVX1_LOC_34/A NAND2X1_LOC_722/A 0.07fF
C72268 D_INPUT_1 INVX1_LOC_76/A 0.14fF
C72269 INVX1_LOC_26/Y INVX1_LOC_117/A 0.10fF
C72270 NOR2X1_LOC_405/A NOR2X1_LOC_109/Y 0.10fF
C72271 NAND2X1_LOC_837/Y NAND2X1_LOC_859/B 0.25fF
C72272 NAND2X1_LOC_725/Y INVX1_LOC_46/A 0.06fF
C72273 INVX1_LOC_225/A NOR2X1_LOC_709/A 0.76fF
C72274 INVX1_LOC_71/A INVX1_LOC_16/A 0.15fF
C72275 INVX1_LOC_276/A NAND2X1_LOC_354/B 0.13fF
C72276 NOR2X1_LOC_602/B NAND2X1_LOC_175/Y 0.01fF
C72277 NAND2X1_LOC_363/B NAND2X1_LOC_441/a_36_24# 0.00fF
C72278 NOR2X1_LOC_606/Y INPUT_1 0.06fF
C72279 INVX1_LOC_257/A NAND2X1_LOC_425/Y 0.02fF
C72280 NAND2X1_LOC_207/B NOR2X1_LOC_721/B 0.03fF
C72281 NOR2X1_LOC_770/A INVX1_LOC_22/A 0.01fF
C72282 INVX1_LOC_83/A NAND2X1_LOC_481/a_36_24# 0.01fF
C72283 INVX1_LOC_174/A NOR2X1_LOC_163/Y 0.17fF
C72284 NAND2X1_LOC_175/Y INVX1_LOC_54/A 0.07fF
C72285 NOR2X1_LOC_856/B NOR2X1_LOC_777/B 0.04fF
C72286 INVX1_LOC_315/Y NAND2X1_LOC_473/A 0.08fF
C72287 INVX1_LOC_232/Y NOR2X1_LOC_6/B 0.08fF
C72288 INVX1_LOC_157/A NAND2X1_LOC_197/a_36_24# 0.00fF
C72289 NOR2X1_LOC_795/Y NOR2X1_LOC_808/A 0.04fF
C72290 NOR2X1_LOC_433/A NAND2X1_LOC_660/Y 0.07fF
C72291 NOR2X1_LOC_557/Y INVX1_LOC_232/A 0.10fF
C72292 NAND2X1_LOC_738/B NOR2X1_LOC_765/Y 0.02fF
C72293 INVX1_LOC_207/A INVX1_LOC_22/A 0.78fF
C72294 NOR2X1_LOC_78/B NOR2X1_LOC_300/Y 0.07fF
C72295 INVX1_LOC_45/A INVX1_LOC_28/A 5.64fF
C72296 NOR2X1_LOC_811/A INVX1_LOC_49/A 0.09fF
C72297 NAND2X1_LOC_338/B NOR2X1_LOC_84/Y 0.14fF
C72298 NOR2X1_LOC_84/A INVX1_LOC_316/Y 0.08fF
C72299 NOR2X1_LOC_810/A INVX1_LOC_49/A 0.04fF
C72300 NOR2X1_LOC_516/B NOR2X1_LOC_516/Y 0.00fF
C72301 NAND2X1_LOC_326/A NOR2X1_LOC_311/Y 0.00fF
C72302 INVX1_LOC_13/A NOR2X1_LOC_340/Y 0.01fF
C72303 INVX1_LOC_276/A INVX1_LOC_276/Y 0.09fF
C72304 INVX1_LOC_76/A NOR2X1_LOC_652/Y 0.10fF
C72305 INVX1_LOC_19/A NOR2X1_LOC_460/A 0.01fF
C72306 NAND2X1_LOC_830/a_36_24# INVX1_LOC_18/A 0.00fF
C72307 NOR2X1_LOC_401/Y INVX1_LOC_256/Y 0.03fF
C72308 NOR2X1_LOC_773/Y NOR2X1_LOC_312/a_36_216# 0.01fF
C72309 NAND2X1_LOC_736/Y NAND2X1_LOC_863/a_36_24# 0.01fF
C72310 NAND2X1_LOC_618/Y NOR2X1_LOC_649/B 0.06fF
C72311 NOR2X1_LOC_189/a_36_216# INVX1_LOC_102/A 0.02fF
C72312 NOR2X1_LOC_641/Y NOR2X1_LOC_748/A 0.02fF
C72313 INVX1_LOC_144/Y NAND2X1_LOC_798/A 0.08fF
C72314 NOR2X1_LOC_764/Y INVX1_LOC_49/A 0.01fF
C72315 INVX1_LOC_19/A INVX1_LOC_3/Y 0.07fF
C72316 INVX1_LOC_30/A INPUT_0 0.21fF
C72317 NOR2X1_LOC_52/B NAND2X1_LOC_660/Y 0.02fF
C72318 NOR2X1_LOC_91/A NOR2X1_LOC_88/Y 0.03fF
C72319 NOR2X1_LOC_678/A INVX1_LOC_9/A 0.03fF
C72320 NOR2X1_LOC_654/A INVX1_LOC_92/A 1.06fF
C72321 INVX1_LOC_143/A INVX1_LOC_232/A 0.10fF
C72322 INVX1_LOC_28/A INVX1_LOC_71/A 0.07fF
C72323 NAND2X1_LOC_330/a_36_24# INVX1_LOC_28/A 0.01fF
C72324 NAND2X1_LOC_371/a_36_24# INVX1_LOC_75/A 0.00fF
C72325 NOR2X1_LOC_539/a_36_216# INVX1_LOC_22/A 0.00fF
C72326 NOR2X1_LOC_296/a_36_216# INVX1_LOC_95/Y 0.00fF
C72327 NOR2X1_LOC_488/a_36_216# NOR2X1_LOC_488/Y 0.00fF
C72328 NOR2X1_LOC_473/B INVX1_LOC_33/A 0.01fF
C72329 INVX1_LOC_90/A NAND2X1_LOC_833/Y 0.45fF
C72330 INVX1_LOC_13/A NOR2X1_LOC_655/B 0.05fF
C72331 NOR2X1_LOC_276/Y NOR2X1_LOC_139/Y 0.03fF
C72332 NOR2X1_LOC_216/B INVX1_LOC_57/A 0.01fF
C72333 NAND2X1_LOC_326/A INVX1_LOC_46/A 0.06fF
C72334 NAND2X1_LOC_807/B INVX1_LOC_32/A 0.10fF
C72335 INVX1_LOC_35/A NOR2X1_LOC_612/Y 0.02fF
C72336 D_INPUT_0 NOR2X1_LOC_52/B 0.24fF
C72337 INVX1_LOC_83/A NOR2X1_LOC_87/B 0.11fF
C72338 INVX1_LOC_141/Y INVX1_LOC_91/A 0.04fF
C72339 INVX1_LOC_2/A INVX1_LOC_157/A 0.03fF
C72340 INVX1_LOC_55/Y NOR2X1_LOC_142/Y 0.07fF
C72341 NOR2X1_LOC_88/Y INVX1_LOC_23/A 0.03fF
C72342 NOR2X1_LOC_91/A INVX1_LOC_84/A 2.44fF
C72343 INVX1_LOC_39/A NOR2X1_LOC_536/A 0.06fF
C72344 INVX1_LOC_296/A NOR2X1_LOC_430/Y 0.03fF
C72345 INVX1_LOC_267/Y INVX1_LOC_135/A 0.03fF
C72346 INVX1_LOC_75/A NOR2X1_LOC_712/B 0.08fF
C72347 NOR2X1_LOC_276/Y NAND2X1_LOC_468/B 0.22fF
C72348 NOR2X1_LOC_541/Y NOR2X1_LOC_35/Y 0.16fF
C72349 NOR2X1_LOC_533/a_36_216# NAND2X1_LOC_811/Y 0.00fF
C72350 INVX1_LOC_314/Y NOR2X1_LOC_74/A 0.01fF
C72351 INVX1_LOC_11/A NOR2X1_LOC_266/B 0.03fF
C72352 INVX1_LOC_9/Y INVX1_LOC_215/A 0.02fF
C72353 INVX1_LOC_216/Y VDD 0.41fF
C72354 INVX1_LOC_200/A NAND2X1_LOC_633/Y 0.09fF
C72355 INVX1_LOC_141/Y INVX1_LOC_11/Y 0.32fF
C72356 INVX1_LOC_36/A NOR2X1_LOC_113/A 0.06fF
C72357 INVX1_LOC_226/Y NOR2X1_LOC_391/A 0.03fF
C72358 INVX1_LOC_50/A NOR2X1_LOC_631/A 0.04fF
C72359 INVX1_LOC_36/A NOR2X1_LOC_405/A 0.07fF
C72360 INVX1_LOC_314/Y NOR2X1_LOC_9/Y -0.00fF
C72361 INVX1_LOC_84/A INVX1_LOC_23/A 0.13fF
C72362 NOR2X1_LOC_679/Y VDD 0.35fF
C72363 INVX1_LOC_5/A NOR2X1_LOC_155/A 0.10fF
C72364 INVX1_LOC_17/A NAND2X1_LOC_96/A 0.07fF
C72365 NOR2X1_LOC_679/Y NAND2X1_LOC_800/A 0.00fF
C72366 INVX1_LOC_13/A NAND2X1_LOC_358/Y 0.06fF
C72367 INVX1_LOC_21/A NAND2X1_LOC_243/Y 0.03fF
C72368 NOR2X1_LOC_655/B INVX1_LOC_55/Y 0.12fF
C72369 NOR2X1_LOC_667/A NAND2X1_LOC_703/a_36_24# 0.00fF
C72370 INVX1_LOC_232/A NOR2X1_LOC_130/A 0.03fF
C72371 NOR2X1_LOC_546/B INVX1_LOC_91/A 0.00fF
C72372 INVX1_LOC_45/A NOR2X1_LOC_35/Y 0.03fF
C72373 INVX1_LOC_136/A NAND2X1_LOC_468/B 0.03fF
C72374 INVX1_LOC_21/A NOR2X1_LOC_61/A 0.01fF
C72375 NOR2X1_LOC_510/Y NAND2X1_LOC_798/B 0.05fF
C72376 NOR2X1_LOC_778/B NOR2X1_LOC_356/A 0.03fF
C72377 NOR2X1_LOC_48/B NAND2X1_LOC_175/Y 0.09fF
C72378 NOR2X1_LOC_103/Y NAND2X1_LOC_236/a_36_24# 0.00fF
C72379 NOR2X1_LOC_626/Y INVX1_LOC_179/A 0.01fF
C72380 INVX1_LOC_64/A NOR2X1_LOC_127/Y 0.06fF
C72381 INVX1_LOC_58/A INVX1_LOC_19/A 0.21fF
C72382 INVX1_LOC_11/A NAND2X1_LOC_848/A 0.01fF
C72383 NOR2X1_LOC_568/A NOR2X1_LOC_35/Y 0.10fF
C72384 NAND2X1_LOC_538/a_36_24# NOR2X1_LOC_52/B 0.00fF
C72385 INVX1_LOC_13/A NOR2X1_LOC_99/B 0.01fF
C72386 INVX1_LOC_83/A INVX1_LOC_174/Y 0.02fF
C72387 NOR2X1_LOC_717/B NOR2X1_LOC_730/A 0.01fF
C72388 NAND2X1_LOC_733/A VDD 0.15fF
C72389 INVX1_LOC_57/Y INVX1_LOC_20/A 0.04fF
C72390 NOR2X1_LOC_791/B INVX1_LOC_59/Y 0.18fF
C72391 INVX1_LOC_58/A NOR2X1_LOC_11/Y 0.01fF
C72392 NAND2X1_LOC_483/Y INVX1_LOC_309/A 0.01fF
C72393 NAND2X1_LOC_560/A NAND2X1_LOC_839/A 0.00fF
C72394 NOR2X1_LOC_68/A NAND2X1_LOC_434/a_36_24# 0.01fF
C72395 INVX1_LOC_89/A GATE_479 0.01fF
C72396 NOR2X1_LOC_92/Y NAND2X1_LOC_802/Y 0.01fF
C72397 NOR2X1_LOC_607/A NOR2X1_LOC_137/B 0.00fF
C72398 INVX1_LOC_275/A INVX1_LOC_91/A 0.03fF
C72399 NAND2X1_LOC_722/A INPUT_0 0.02fF
C72400 INVX1_LOC_286/Y INVX1_LOC_33/Y 0.01fF
C72401 NOR2X1_LOC_248/a_36_216# INVX1_LOC_53/Y 0.00fF
C72402 INVX1_LOC_25/A INVX1_LOC_284/A 0.77fF
C72403 NOR2X1_LOC_48/B INVX1_LOC_262/A 0.03fF
C72404 NAND2X1_LOC_863/A NAND2X1_LOC_852/Y 0.10fF
C72405 NAND2X1_LOC_483/Y INVX1_LOC_91/A 0.02fF
C72406 NOR2X1_LOC_186/Y INVX1_LOC_294/A 0.12fF
C72407 NOR2X1_LOC_91/A INVX1_LOC_15/A 0.03fF
C72408 INVX1_LOC_39/A INVX1_LOC_3/A 0.03fF
C72409 NOR2X1_LOC_778/B NOR2X1_LOC_74/A 0.06fF
C72410 NOR2X1_LOC_201/A INVX1_LOC_15/A 0.17fF
C72411 NOR2X1_LOC_219/Y NOR2X1_LOC_202/Y 0.09fF
C72412 INVX1_LOC_71/A NOR2X1_LOC_35/Y 0.39fF
C72413 INVX1_LOC_2/A INVX1_LOC_69/Y 0.07fF
C72414 INVX1_LOC_93/A NOR2X1_LOC_662/A 0.02fF
C72415 NAND2X1_LOC_303/Y NAND2X1_LOC_809/a_36_24# 0.06fF
C72416 NOR2X1_LOC_403/B INVX1_LOC_76/A 0.01fF
C72417 INVX1_LOC_200/A INVX1_LOC_71/Y 0.16fF
C72418 NOR2X1_LOC_272/Y INVX1_LOC_63/A 0.49fF
C72419 NAND2X1_LOC_550/A NOR2X1_LOC_487/Y 0.04fF
C72420 NOR2X1_LOC_68/A INVX1_LOC_12/Y 0.02fF
C72421 NOR2X1_LOC_383/B INVX1_LOC_4/A 0.52fF
C72422 INVX1_LOC_32/A NAND2X1_LOC_215/A -0.00fF
C72423 NOR2X1_LOC_75/Y INVX1_LOC_92/A 0.02fF
C72424 NOR2X1_LOC_589/A NOR2X1_LOC_163/Y 0.00fF
C72425 NOR2X1_LOC_309/Y NOR2X1_LOC_405/A 0.01fF
C72426 NOR2X1_LOC_557/Y NAND2X1_LOC_447/Y 0.04fF
C72427 INVX1_LOC_23/A INVX1_LOC_15/A 2.00fF
C72428 NAND2X1_LOC_337/B NOR2X1_LOC_155/A 0.13fF
C72429 NOR2X1_LOC_180/B INVX1_LOC_97/A 0.03fF
C72430 NOR2X1_LOC_716/B NOR2X1_LOC_9/a_36_216# 0.00fF
C72431 NOR2X1_LOC_160/B NOR2X1_LOC_461/A 0.03fF
C72432 INVX1_LOC_13/Y NAND2X1_LOC_74/B 0.10fF
C72433 NOR2X1_LOC_168/B INVX1_LOC_91/A 0.08fF
C72434 NAND2X1_LOC_743/a_36_24# INVX1_LOC_301/A 0.01fF
C72435 NAND2X1_LOC_35/Y INVX1_LOC_42/A 2.13fF
C72436 INVX1_LOC_61/A NOR2X1_LOC_536/A 1.11fF
C72437 INVX1_LOC_143/A INVX1_LOC_186/A 0.02fF
C72438 INVX1_LOC_90/A NOR2X1_LOC_180/B 2.98fF
C72439 INVX1_LOC_5/A NOR2X1_LOC_833/B 0.06fF
C72440 NOR2X1_LOC_644/B INVX1_LOC_307/A 0.01fF
C72441 INVX1_LOC_75/A INVX1_LOC_164/A 0.05fF
C72442 NOR2X1_LOC_124/B INVX1_LOC_112/A 0.01fF
C72443 NOR2X1_LOC_709/A NAND2X1_LOC_642/Y 0.55fF
C72444 NAND2X1_LOC_348/A NOR2X1_LOC_719/B 0.01fF
C72445 NOR2X1_LOC_142/Y NOR2X1_LOC_357/Y 0.46fF
C72446 NAND2X1_LOC_656/Y INVX1_LOC_79/A 0.10fF
C72447 INVX1_LOC_27/A NOR2X1_LOC_33/B 0.03fF
C72448 NAND2X1_LOC_564/B INVX1_LOC_286/A 0.17fF
C72449 INVX1_LOC_31/A NOR2X1_LOC_88/Y 23.15fF
C72450 NAND2X1_LOC_207/B NAND2X1_LOC_473/A 0.01fF
C72451 INVX1_LOC_87/A INVX1_LOC_29/Y 0.04fF
C72452 INVX1_LOC_170/Y INVX1_LOC_306/Y 0.02fF
C72453 INVX1_LOC_289/A NOR2X1_LOC_45/B 0.33fF
C72454 NOR2X1_LOC_591/Y INVX1_LOC_76/A 0.12fF
C72455 INVX1_LOC_173/Y NOR2X1_LOC_409/Y 0.70fF
C72456 INVX1_LOC_90/A INVX1_LOC_73/A 0.03fF
C72457 NOR2X1_LOC_52/B NOR2X1_LOC_266/B 0.05fF
C72458 NAND2X1_LOC_571/Y INVX1_LOC_42/A 0.46fF
C72459 NOR2X1_LOC_300/Y INVX1_LOC_46/A 0.00fF
C72460 NOR2X1_LOC_269/Y INVX1_LOC_22/A 0.06fF
C72461 NOR2X1_LOC_384/Y NAND2X1_LOC_243/B 0.01fF
C72462 NOR2X1_LOC_310/Y INVX1_LOC_14/Y 0.00fF
C72463 NOR2X1_LOC_389/B INVX1_LOC_73/A 0.07fF
C72464 INVX1_LOC_88/A NAND2X1_LOC_74/B 0.03fF
C72465 NOR2X1_LOC_795/Y INVX1_LOC_37/A 0.01fF
C72466 INVX1_LOC_1/A INVX1_LOC_284/A 0.10fF
C72467 INVX1_LOC_31/A INVX1_LOC_84/A 0.81fF
C72468 NOR2X1_LOC_318/B INVX1_LOC_101/A 0.00fF
C72469 NOR2X1_LOC_160/B NAND2X1_LOC_782/B 0.07fF
C72470 NOR2X1_LOC_736/Y NOR2X1_LOC_742/A 0.20fF
C72471 NOR2X1_LOC_142/Y INVX1_LOC_66/Y 0.24fF
C72472 NAND2X1_LOC_833/Y INVX1_LOC_38/A 0.18fF
C72473 NOR2X1_LOC_342/B NOR2X1_LOC_260/Y 0.19fF
C72474 INVX1_LOC_215/Y INVX1_LOC_19/A 0.01fF
C72475 NOR2X1_LOC_479/B NAND2X1_LOC_659/B 0.16fF
C72476 INVX1_LOC_256/A NAND2X1_LOC_63/Y 0.03fF
C72477 NAND2X1_LOC_564/B INVX1_LOC_95/A 0.06fF
C72478 NAND2X1_LOC_360/B INVX1_LOC_46/A 0.47fF
C72479 INVX1_LOC_255/Y INVX1_LOC_255/A 0.13fF
C72480 NAND2X1_LOC_162/B INVX1_LOC_92/A 0.17fF
C72481 NAND2X1_LOC_656/Y INVX1_LOC_91/A 1.14fF
C72482 NOR2X1_LOC_91/A INVX1_LOC_278/A 0.12fF
C72483 NOR2X1_LOC_336/B INVX1_LOC_63/A 0.09fF
C72484 NOR2X1_LOC_52/B NAND2X1_LOC_848/A 0.28fF
C72485 NOR2X1_LOC_355/A NOR2X1_LOC_318/B 0.35fF
C72486 NOR2X1_LOC_419/Y INVX1_LOC_92/A 0.01fF
C72487 INVX1_LOC_53/A NOR2X1_LOC_654/A 0.16fF
C72488 NOR2X1_LOC_703/Y INVX1_LOC_196/Y 0.02fF
C72489 NOR2X1_LOC_322/Y NOR2X1_LOC_323/Y 0.01fF
C72490 NOR2X1_LOC_479/B VDD 0.03fF
C72491 NOR2X1_LOC_667/A NAND2X1_LOC_284/a_36_24# 0.00fF
C72492 NAND2X1_LOC_662/B NAND2X1_LOC_661/A 0.09fF
C72493 NOR2X1_LOC_82/Y NOR2X1_LOC_558/A 0.03fF
C72494 NOR2X1_LOC_328/Y INVX1_LOC_146/Y 0.15fF
C72495 INVX1_LOC_30/A NOR2X1_LOC_48/a_36_216# 0.01fF
C72496 INVX1_LOC_181/Y INVX1_LOC_285/A 0.01fF
C72497 NOR2X1_LOC_716/B INVX1_LOC_92/A 0.05fF
C72498 INVX1_LOC_64/A NOR2X1_LOC_383/B 1.27fF
C72499 NOR2X1_LOC_709/A NOR2X1_LOC_271/Y 0.08fF
C72500 NOR2X1_LOC_134/Y NOR2X1_LOC_89/A 0.03fF
C72501 NOR2X1_LOC_328/Y VDD 1.08fF
C72502 NOR2X1_LOC_551/Y NOR2X1_LOC_703/A 0.01fF
C72503 NAND2X1_LOC_364/A INVX1_LOC_63/A 0.17fF
C72504 NOR2X1_LOC_590/A NOR2X1_LOC_67/a_36_216# 0.00fF
C72505 NOR2X1_LOC_455/Y D_INPUT_1 0.00fF
C72506 NAND2X1_LOC_859/Y NOR2X1_LOC_825/Y 0.00fF
C72507 INVX1_LOC_278/A INVX1_LOC_23/A 0.03fF
C72508 INVX1_LOC_188/A INVX1_LOC_290/Y -0.01fF
C72509 D_INPUT_0 INVX1_LOC_74/A 0.41fF
C72510 NOR2X1_LOC_32/B NAND2X1_LOC_549/Y 0.02fF
C72511 NAND2X1_LOC_477/A INVX1_LOC_291/A 0.10fF
C72512 NAND2X1_LOC_140/A NAND2X1_LOC_469/B 0.01fF
C72513 NAND2X1_LOC_350/A INVX1_LOC_32/A 0.07fF
C72514 INVX1_LOC_30/Y INVX1_LOC_129/Y 0.02fF
C72515 INVX1_LOC_304/Y INVX1_LOC_71/Y 0.13fF
C72516 INVX1_LOC_72/A INVX1_LOC_261/Y 0.04fF
C72517 NAND2X1_LOC_182/a_36_24# NOR2X1_LOC_536/A 0.01fF
C72518 NOR2X1_LOC_15/Y NOR2X1_LOC_278/Y 0.03fF
C72519 NAND2X1_LOC_725/B NOR2X1_LOC_395/Y 0.01fF
C72520 INVX1_LOC_93/A INVX1_LOC_57/A 0.08fF
C72521 INVX1_LOC_219/A VDD -0.00fF
C72522 NOR2X1_LOC_92/a_36_216# NOR2X1_LOC_76/A 0.01fF
C72523 NOR2X1_LOC_384/Y INVX1_LOC_284/A 0.18fF
C72524 NOR2X1_LOC_341/a_36_216# INVX1_LOC_19/A 0.02fF
C72525 INVX1_LOC_40/A NOR2X1_LOC_54/a_36_216# 0.01fF
C72526 NOR2X1_LOC_598/B INVX1_LOC_5/A 0.72fF
C72527 INVX1_LOC_35/A NAND2X1_LOC_406/a_36_24# 0.00fF
C72528 INVX1_LOC_31/A INVX1_LOC_15/A 0.39fF
C72529 INVX1_LOC_16/A NOR2X1_LOC_331/B 0.07fF
C72530 NOR2X1_LOC_441/Y INVX1_LOC_32/A 0.02fF
C72531 NOR2X1_LOC_557/A NOR2X1_LOC_74/A 0.02fF
C72532 NAND2X1_LOC_560/A NOR2X1_LOC_823/Y 0.01fF
C72533 NAND2X1_LOC_562/Y NOR2X1_LOC_649/B 0.03fF
C72534 INVX1_LOC_202/A INVX1_LOC_272/A 0.03fF
C72535 NOR2X1_LOC_45/Y NOR2X1_LOC_334/Y 0.11fF
C72536 INVX1_LOC_224/Y INVX1_LOC_48/Y 0.50fF
C72537 NOR2X1_LOC_160/B NAND2X1_LOC_454/Y 0.07fF
C72538 NAND2X1_LOC_725/A INVX1_LOC_5/A 0.10fF
C72539 INVX1_LOC_221/A INVX1_LOC_119/Y 0.00fF
C72540 INVX1_LOC_225/A INVX1_LOC_294/A 0.12fF
C72541 NOR2X1_LOC_757/Y INVX1_LOC_92/A 0.53fF
C72542 INVX1_LOC_33/Y NAND2X1_LOC_803/a_36_24# 0.00fF
C72543 NOR2X1_LOC_557/A NOR2X1_LOC_9/Y 0.06fF
C72544 INVX1_LOC_303/A NAND2X1_LOC_74/B 0.10fF
C72545 NOR2X1_LOC_658/a_36_216# NOR2X1_LOC_205/Y 0.00fF
C72546 NAND2X1_LOC_784/A NAND2X1_LOC_703/Y 0.31fF
C72547 NAND2X1_LOC_564/B INVX1_LOC_54/A 0.09fF
C72548 NOR2X1_LOC_414/a_36_216# NOR2X1_LOC_38/B 0.00fF
C72549 NOR2X1_LOC_208/Y INVX1_LOC_109/Y 0.03fF
C72550 INVX1_LOC_94/A INVX1_LOC_42/A 0.07fF
C72551 NOR2X1_LOC_706/Y NOR2X1_LOC_725/A 0.00fF
C72552 INVX1_LOC_18/A D_INPUT_5 0.08fF
C72553 INVX1_LOC_25/Y NOR2X1_LOC_235/Y 0.03fF
C72554 INVX1_LOC_78/Y INVX1_LOC_91/A 0.03fF
C72555 INVX1_LOC_49/A NOR2X1_LOC_89/A 0.05fF
C72556 NOR2X1_LOC_441/Y NAND2X1_LOC_175/Y 0.02fF
C72557 NOR2X1_LOC_524/Y INVX1_LOC_94/Y 0.01fF
C72558 INVX1_LOC_63/Y INVX1_LOC_29/A 0.03fF
C72559 INVX1_LOC_22/A NOR2X1_LOC_79/Y 0.02fF
C72560 INVX1_LOC_191/Y INVX1_LOC_84/A 0.03fF
C72561 NOR2X1_LOC_211/A NAND2X1_LOC_255/a_36_24# 0.01fF
C72562 INVX1_LOC_38/Y NOR2X1_LOC_846/A 0.04fF
C72563 NOR2X1_LOC_180/B INVX1_LOC_38/A 0.07fF
C72564 NOR2X1_LOC_470/A INVX1_LOC_92/A 0.19fF
C72565 INVX1_LOC_27/A INVX1_LOC_306/Y 0.48fF
C72566 INVX1_LOC_43/Y NOR2X1_LOC_383/B 0.09fF
C72567 VDD NOR2X1_LOC_196/Y -0.00fF
C72568 NOR2X1_LOC_254/A NOR2X1_LOC_748/A 0.02fF
C72569 NAND2X1_LOC_859/Y NOR2X1_LOC_88/Y 0.10fF
C72570 NAND2X1_LOC_79/Y NOR2X1_LOC_38/B 0.01fF
C72571 NOR2X1_LOC_424/Y INVX1_LOC_92/A 0.19fF
C72572 NAND2X1_LOC_725/A NOR2X1_LOC_494/Y 0.10fF
C72573 NOR2X1_LOC_313/Y NAND2X1_LOC_453/A 0.01fF
C72574 INVX1_LOC_89/A NOR2X1_LOC_641/Y 0.02fF
C72575 INVX1_LOC_286/A NOR2X1_LOC_279/Y 0.00fF
C72576 INVX1_LOC_30/A INVX1_LOC_183/A 0.01fF
C72577 INVX1_LOC_28/A NOR2X1_LOC_331/B 0.15fF
C72578 NAND2X1_LOC_32/a_36_24# NOR2X1_LOC_249/Y 0.00fF
C72579 NOR2X1_LOC_175/A INVX1_LOC_29/A 0.03fF
C72580 NOR2X1_LOC_562/B NOR2X1_LOC_486/Y 0.04fF
C72581 INVX1_LOC_73/A NOR2X1_LOC_561/A 0.02fF
C72582 INVX1_LOC_47/A NAND2X1_LOC_62/a_36_24# 0.02fF
C72583 NAND2X1_LOC_465/Y INVX1_LOC_42/A 0.02fF
C72584 NOR2X1_LOC_234/Y INVX1_LOC_42/A 0.04fF
C72585 NOR2X1_LOC_668/a_36_216# NAND2X1_LOC_114/B 0.01fF
C72586 INVX1_LOC_94/A INVX1_LOC_78/A 0.07fF
C72587 INVX1_LOC_2/A NOR2X1_LOC_89/A 0.15fF
C72588 NAND2X1_LOC_859/Y INVX1_LOC_84/A 0.00fF
C72589 INVX1_LOC_230/Y NOR2X1_LOC_392/Y 0.08fF
C72590 INVX1_LOC_58/A NOR2X1_LOC_599/A 0.03fF
C72591 NAND2X1_LOC_725/A NOR2X1_LOC_816/A 0.03fF
C72592 INVX1_LOC_108/Y INVX1_LOC_31/A 0.02fF
C72593 NOR2X1_LOC_374/A NOR2X1_LOC_334/Y 0.01fF
C72594 NOR2X1_LOC_226/A NOR2X1_LOC_89/A 0.24fF
C72595 INVX1_LOC_278/A INVX1_LOC_31/A 0.07fF
C72596 INVX1_LOC_269/A NAND2X1_LOC_474/Y 0.10fF
C72597 NOR2X1_LOC_67/A NOR2X1_LOC_67/Y 0.11fF
C72598 INVX1_LOC_89/A NOR2X1_LOC_461/B 0.03fF
C72599 INVX1_LOC_25/A INVX1_LOC_72/A 0.07fF
C72600 INVX1_LOC_14/A NOR2X1_LOC_440/B 0.98fF
C72601 NOR2X1_LOC_818/a_36_216# INVX1_LOC_31/A 0.01fF
C72602 NOR2X1_LOC_45/B INVX1_LOC_37/A 0.10fF
C72603 NOR2X1_LOC_341/a_36_216# INVX1_LOC_26/Y 0.00fF
C72604 INVX1_LOC_78/Y NOR2X1_LOC_698/Y 0.01fF
C72605 INVX1_LOC_120/A NAND2X1_LOC_235/a_36_24# 0.01fF
C72606 NOR2X1_LOC_272/a_36_216# INVX1_LOC_256/A 0.12fF
C72607 INVX1_LOC_28/A NOR2X1_LOC_592/B 0.03fF
C72608 NAND2X1_LOC_807/Y NOR2X1_LOC_88/Y 0.07fF
C72609 NOR2X1_LOC_290/Y INVX1_LOC_15/A 0.05fF
C72610 NOR2X1_LOC_218/Y NOR2X1_LOC_89/A 0.00fF
C72611 NOR2X1_LOC_188/a_36_216# INVX1_LOC_29/A 0.00fF
C72612 NOR2X1_LOC_168/Y INVX1_LOC_23/A 0.30fF
C72613 NAND2X1_LOC_773/Y NAND2X1_LOC_774/a_36_24# 0.01fF
C72614 NAND2X1_LOC_787/A NOR2X1_LOC_91/a_36_216# 0.00fF
C72615 NOR2X1_LOC_655/B INVX1_LOC_32/A 0.10fF
C72616 NOR2X1_LOC_500/A INVX1_LOC_57/A 0.02fF
C72617 INVX1_LOC_298/Y INVX1_LOC_63/Y 0.10fF
C72618 INVX1_LOC_2/Y INVX1_LOC_59/Y 0.11fF
C72619 NAND2X1_LOC_866/B INVX1_LOC_84/A 0.01fF
C72620 NOR2X1_LOC_448/Y INVX1_LOC_11/A 0.04fF
C72621 NOR2X1_LOC_65/B NAND2X1_LOC_786/a_36_24# 0.01fF
C72622 INVX1_LOC_247/A INVX1_LOC_37/A 0.03fF
C72623 INVX1_LOC_199/Y INVX1_LOC_37/A 0.39fF
C72624 NAND2X1_LOC_763/B NAND2X1_LOC_25/a_36_24# 0.00fF
C72625 NOR2X1_LOC_609/A INVX1_LOC_53/A 0.02fF
C72626 NAND2X1_LOC_725/Y NAND2X1_LOC_866/A 0.03fF
C72627 INVX1_LOC_108/Y NAND2X1_LOC_106/a_36_24# 0.01fF
C72628 INVX1_LOC_2/Y INVX1_LOC_176/A 0.01fF
C72629 INVX1_LOC_136/A NOR2X1_LOC_772/B 0.57fF
C72630 INVX1_LOC_214/A INVX1_LOC_21/Y 0.06fF
C72631 NOR2X1_LOC_220/B INVX1_LOC_30/A 0.01fF
C72632 NOR2X1_LOC_370/a_36_216# INVX1_LOC_29/A 0.00fF
C72633 NAND2X1_LOC_807/Y INVX1_LOC_84/A 0.16fF
C72634 INVX1_LOC_39/A NOR2X1_LOC_606/Y 0.20fF
C72635 NAND2X1_LOC_740/Y INVX1_LOC_36/A 0.03fF
C72636 NOR2X1_LOC_471/Y NOR2X1_LOC_464/B 0.02fF
C72637 NAND2X1_LOC_624/B NOR2X1_LOC_522/Y 0.16fF
C72638 INVX1_LOC_136/A INVX1_LOC_13/Y 0.17fF
C72639 NAND2X1_LOC_21/Y INVX1_LOC_23/A 0.05fF
C72640 INVX1_LOC_11/A NAND2X1_LOC_30/Y 0.23fF
C72641 NAND2X1_LOC_350/B NAND2X1_LOC_454/Y 0.25fF
C72642 INVX1_LOC_6/A NOR2X1_LOC_88/Y 0.03fF
C72643 INVX1_LOC_88/A NOR2X1_LOC_276/Y 0.01fF
C72644 D_INPUT_0 NAND2X1_LOC_254/Y 0.06fF
C72645 INVX1_LOC_45/A INVX1_LOC_48/Y 0.03fF
C72646 NOR2X1_LOC_136/Y INVX1_LOC_78/A 0.01fF
C72647 INVX1_LOC_225/Y NOR2X1_LOC_457/A 0.50fF
C72648 INVX1_LOC_75/A NAND2X1_LOC_225/a_36_24# 0.00fF
C72649 NAND2X1_LOC_648/A NOR2X1_LOC_89/A 0.03fF
C72650 INVX1_LOC_25/Y NAND2X1_LOC_471/Y 0.00fF
C72651 INVX1_LOC_208/A NAND2X1_LOC_454/Y 0.10fF
C72652 NAND2X1_LOC_721/A NOR2X1_LOC_111/A 0.15fF
C72653 INVX1_LOC_1/A NAND2X1_LOC_136/a_36_24# 0.00fF
C72654 INVX1_LOC_215/Y INVX1_LOC_161/Y 0.40fF
C72655 INPUT_1 NOR2X1_LOC_89/A 0.07fF
C72656 NOR2X1_LOC_70/a_36_216# NOR2X1_LOC_36/B 0.00fF
C72657 NOR2X1_LOC_590/A NOR2X1_LOC_286/Y 0.03fF
C72658 NOR2X1_LOC_331/B NOR2X1_LOC_35/Y 0.19fF
C72659 INVX1_LOC_130/A INVX1_LOC_103/A 0.04fF
C72660 GATE_662 NAND2X1_LOC_3/B 0.18fF
C72661 INVX1_LOC_224/Y NOR2X1_LOC_84/Y 0.19fF
C72662 NOR2X1_LOC_448/A NAND2X1_LOC_93/B 0.01fF
C72663 NOR2X1_LOC_166/a_36_216# INVX1_LOC_102/A 0.01fF
C72664 NOR2X1_LOC_71/Y INVX1_LOC_19/Y 0.03fF
C72665 NOR2X1_LOC_559/B INVX1_LOC_50/Y 0.02fF
C72666 INVX1_LOC_6/A INVX1_LOC_84/A 0.10fF
C72667 INVX1_LOC_1/A INVX1_LOC_72/A 0.35fF
C72668 NOR2X1_LOC_598/B NOR2X1_LOC_377/Y 0.01fF
C72669 NOR2X1_LOC_99/B INVX1_LOC_32/A 0.09fF
C72670 INVX1_LOC_54/Y INVX1_LOC_57/A 0.14fF
C72671 INVX1_LOC_1/A INVX1_LOC_142/Y 0.01fF
C72672 INVX1_LOC_58/A NAND2X1_LOC_335/a_36_24# 0.00fF
C72673 INVX1_LOC_136/A INVX1_LOC_88/A 0.02fF
C72674 NOR2X1_LOC_448/A NAND2X1_LOC_425/Y 0.01fF
C72675 INVX1_LOC_37/A NOR2X1_LOC_499/B 0.03fF
C72676 INVX1_LOC_22/A INVX1_LOC_26/A 0.01fF
C72677 INVX1_LOC_239/Y NAND2X1_LOC_402/B 0.01fF
C72678 NAND2X1_LOC_84/Y NOR2X1_LOC_440/B 0.01fF
C72679 INVX1_LOC_64/A NAND2X1_LOC_706/a_36_24# 0.01fF
C72680 NOR2X1_LOC_689/Y NOR2X1_LOC_773/Y 0.04fF
C72681 NAND2X1_LOC_564/B NOR2X1_LOC_438/Y 0.01fF
C72682 INVX1_LOC_25/A NAND2X1_LOC_338/B 0.11fF
C72683 INVX1_LOC_1/A INVX1_LOC_198/Y 0.10fF
C72684 NAND2X1_LOC_725/Y NOR2X1_LOC_505/Y 0.11fF
C72685 NOR2X1_LOC_15/Y NAND2X1_LOC_731/Y 0.02fF
C72686 D_INPUT_3 NOR2X1_LOC_655/Y 2.20fF
C72687 NAND2X1_LOC_555/Y NAND2X1_LOC_577/A 0.05fF
C72688 NOR2X1_LOC_2/Y NOR2X1_LOC_25/a_36_216# 0.00fF
C72689 INVX1_LOC_14/A INVX1_LOC_41/Y 0.02fF
C72690 NAND2X1_LOC_804/Y INVX1_LOC_54/A 0.00fF
C72691 NAND2X1_LOC_807/Y INVX1_LOC_15/A 0.07fF
C72692 NOR2X1_LOC_675/A INVX1_LOC_285/A -0.03fF
C72693 INVX1_LOC_67/Y NOR2X1_LOC_114/Y 0.00fF
C72694 INVX1_LOC_17/A NAND2X1_LOC_656/A 0.09fF
C72695 INVX1_LOC_37/A NOR2X1_LOC_676/Y 0.01fF
C72696 NOR2X1_LOC_6/B INVX1_LOC_50/Y 0.44fF
C72697 NOR2X1_LOC_750/A NOR2X1_LOC_38/B 0.01fF
C72698 NAND2X1_LOC_357/B NOR2X1_LOC_406/A 0.02fF
C72699 NAND2X1_LOC_858/B INVX1_LOC_102/A 0.15fF
C72700 NOR2X1_LOC_78/A NAND2X1_LOC_773/B 0.07fF
C72701 INVX1_LOC_5/A NOR2X1_LOC_156/B 0.03fF
C72702 NOR2X1_LOC_405/A INVX1_LOC_63/A 0.02fF
C72703 INVX1_LOC_103/A INVX1_LOC_81/A 0.03fF
C72704 NOR2X1_LOC_68/A NOR2X1_LOC_160/B 0.40fF
C72705 INVX1_LOC_286/Y NAND2X1_LOC_741/B 0.61fF
C72706 INVX1_LOC_37/A NOR2X1_LOC_862/B 0.03fF
C72707 NOR2X1_LOC_750/a_36_216# NOR2X1_LOC_38/B 0.00fF
C72708 NAND2X1_LOC_725/A NOR2X1_LOC_773/Y 0.10fF
C72709 NOR2X1_LOC_203/a_36_216# NOR2X1_LOC_203/Y 0.00fF
C72710 INVX1_LOC_46/A NAND2X1_LOC_572/B 0.15fF
C72711 INVX1_LOC_11/A INVX1_LOC_49/A 3.45fF
C72712 D_INPUT_3 NOR2X1_LOC_649/B 0.17fF
C72713 VDD INVX1_LOC_220/A 0.12fF
C72714 NOR2X1_LOC_612/B NOR2X1_LOC_440/B 0.51fF
C72715 INVX1_LOC_266/A NOR2X1_LOC_6/B -0.04fF
C72716 NAND2X1_LOC_725/Y NOR2X1_LOC_700/Y 0.47fF
C72717 D_INPUT_3 INVX1_LOC_3/A 0.11fF
C72718 INVX1_LOC_278/A NAND2X1_LOC_859/Y 0.16fF
C72719 INVX1_LOC_78/Y NOR2X1_LOC_483/a_36_216# 0.00fF
C72720 NOR2X1_LOC_381/Y NOR2X1_LOC_6/B 0.00fF
C72721 D_INPUT_4 NOR2X1_LOC_30/Y 0.03fF
C72722 NAND2X1_LOC_391/Y INVX1_LOC_256/Y 0.00fF
C72723 NOR2X1_LOC_857/A INVX1_LOC_63/A 0.07fF
C72724 INVX1_LOC_6/A INVX1_LOC_15/A 0.31fF
C72725 NOR2X1_LOC_561/Y NOR2X1_LOC_678/A 0.07fF
C72726 INVX1_LOC_225/A INVX1_LOC_308/Y 0.01fF
C72727 NAND2X1_LOC_361/Y NOR2X1_LOC_785/A 0.01fF
C72728 INVX1_LOC_141/A NOR2X1_LOC_577/Y 0.02fF
C72729 NOR2X1_LOC_717/B INVX1_LOC_53/A 0.06fF
C72730 INVX1_LOC_80/A NOR2X1_LOC_660/Y 0.08fF
C72731 NOR2X1_LOC_598/B NOR2X1_LOC_332/A 2.80fF
C72732 INVX1_LOC_124/Y INVX1_LOC_314/Y 0.01fF
C72733 NOR2X1_LOC_625/a_36_216# NOR2X1_LOC_384/Y 0.00fF
C72734 INVX1_LOC_18/A NOR2X1_LOC_360/Y 0.10fF
C72735 INVX1_LOC_144/A INVX1_LOC_78/A 0.03fF
C72736 INVX1_LOC_1/A INVX1_LOC_192/Y 0.04fF
C72737 INVX1_LOC_137/A INVX1_LOC_306/Y 0.00fF
C72738 NOR2X1_LOC_246/A INVX1_LOC_308/A 0.03fF
C72739 INVX1_LOC_1/A NOR2X1_LOC_537/Y 0.52fF
C72740 INVX1_LOC_1/A NAND2X1_LOC_338/B 0.01fF
C72741 NOR2X1_LOC_272/Y INVX1_LOC_1/Y 0.19fF
C72742 NOR2X1_LOC_454/Y NAND2X1_LOC_841/A 0.09fF
C72743 NOR2X1_LOC_103/Y NOR2X1_LOC_84/Y 0.14fF
C72744 INVX1_LOC_171/A NOR2X1_LOC_405/Y 0.12fF
C72745 NOR2X1_LOC_828/A INVX1_LOC_53/A 0.06fF
C72746 INVX1_LOC_1/A NAND2X1_LOC_323/B 0.07fF
C72747 INVX1_LOC_50/A NOR2X1_LOC_385/Y 0.05fF
C72748 INVX1_LOC_136/A INVX1_LOC_303/A 0.10fF
C72749 INVX1_LOC_21/A INVX1_LOC_215/A 0.04fF
C72750 INVX1_LOC_2/A INVX1_LOC_11/A 2.11fF
C72751 NOR2X1_LOC_15/Y INVX1_LOC_197/Y 0.03fF
C72752 NOR2X1_LOC_454/Y INVX1_LOC_268/A 0.04fF
C72753 NAND2X1_LOC_149/Y NAND2X1_LOC_479/Y 0.15fF
C72754 NOR2X1_LOC_471/Y NOR2X1_LOC_423/Y 0.14fF
C72755 INVX1_LOC_100/A INVX1_LOC_26/A 0.04fF
C72756 NOR2X1_LOC_723/a_36_216# INVX1_LOC_113/Y 0.00fF
C72757 NOR2X1_LOC_65/B INVX1_LOC_144/A 0.00fF
C72758 NOR2X1_LOC_7/Y NAND2X1_LOC_470/B 0.04fF
C72759 NOR2X1_LOC_335/B INVX1_LOC_28/Y 0.03fF
C72760 NOR2X1_LOC_78/A NAND2X1_LOC_615/a_36_24# 0.01fF
C72761 NOR2X1_LOC_382/Y INVX1_LOC_34/A 0.07fF
C72762 NOR2X1_LOC_226/A INVX1_LOC_11/A 0.10fF
C72763 INVX1_LOC_230/Y NAND2X1_LOC_755/a_36_24# 0.00fF
C72764 NAND2X1_LOC_392/A NOR2X1_LOC_15/Y 0.01fF
C72765 INVX1_LOC_269/A NOR2X1_LOC_500/Y 0.02fF
C72766 INVX1_LOC_226/Y INVX1_LOC_269/A 0.01fF
C72767 NOR2X1_LOC_75/Y NOR2X1_LOC_78/B 0.02fF
C72768 NAND2X1_LOC_796/B NAND2X1_LOC_783/A 0.21fF
C72769 INVX1_LOC_21/A NOR2X1_LOC_373/Y 0.01fF
C72770 NOR2X1_LOC_655/B INPUT_3 0.15fF
C72771 NOR2X1_LOC_536/A NOR2X1_LOC_831/Y 0.27fF
C72772 NOR2X1_LOC_457/B INVX1_LOC_33/A 0.08fF
C72773 NOR2X1_LOC_471/Y NOR2X1_LOC_222/Y 0.07fF
C72774 NOR2X1_LOC_151/Y INVX1_LOC_53/A 0.14fF
C72775 INVX1_LOC_235/Y INVX1_LOC_135/A 0.43fF
C72776 NAND2X1_LOC_594/a_36_24# NOR2X1_LOC_246/A 0.00fF
C72777 NOR2X1_LOC_68/A NOR2X1_LOC_523/a_36_216# 0.00fF
C72778 INVX1_LOC_11/A NOR2X1_LOC_161/Y 0.02fF
C72779 INVX1_LOC_45/A NOR2X1_LOC_84/Y 0.11fF
C72780 INVX1_LOC_30/A INVX1_LOC_266/Y 0.03fF
C72781 INVX1_LOC_250/A NAND2X1_LOC_357/B 0.03fF
C72782 INVX1_LOC_47/Y NAND2X1_LOC_267/B 0.01fF
C72783 NOR2X1_LOC_48/B NAND2X1_LOC_804/Y 0.45fF
C72784 NOR2X1_LOC_99/Y INVX1_LOC_293/Y 0.20fF
C72785 NOR2X1_LOC_331/B INVX1_LOC_109/A 0.03fF
C72786 INVX1_LOC_136/A INVX1_LOC_168/A 0.05fF
C72787 NOR2X1_LOC_433/A INVX1_LOC_49/A 0.08fF
C72788 INVX1_LOC_269/A INVX1_LOC_10/A 0.13fF
C72789 INVX1_LOC_149/A NOR2X1_LOC_274/B 0.21fF
C72790 NAND2X1_LOC_848/A NAND2X1_LOC_254/Y 0.04fF
C72791 INVX1_LOC_236/Y NAND2X1_LOC_840/B 0.09fF
C72792 NAND2X1_LOC_634/a_36_24# NOR2X1_LOC_71/Y 0.00fF
C72793 INVX1_LOC_91/A NOR2X1_LOC_727/B 0.03fF
C72794 NOR2X1_LOC_617/Y INVX1_LOC_217/Y 0.12fF
C72795 INVX1_LOC_49/A NOR2X1_LOC_593/Y 0.02fF
C72796 INVX1_LOC_177/Y INVX1_LOC_133/Y 0.06fF
C72797 INVX1_LOC_222/A NOR2X1_LOC_405/Y 0.01fF
C72798 INVX1_LOC_12/A NOR2X1_LOC_629/Y 0.03fF
C72799 NOR2X1_LOC_89/A INVX1_LOC_118/A 0.52fF
C72800 INVX1_LOC_57/Y NAND2X1_LOC_850/Y 0.11fF
C72801 INVX1_LOC_35/Y NOR2X1_LOC_662/A 0.20fF
C72802 NOR2X1_LOC_405/A NOR2X1_LOC_65/Y 0.14fF
C72803 NOR2X1_LOC_391/a_36_216# NOR2X1_LOC_392/Y 0.01fF
C72804 NOR2X1_LOC_68/A INVX1_LOC_189/A -0.02fF
C72805 INVX1_LOC_278/A INVX1_LOC_6/A 0.18fF
C72806 INVX1_LOC_18/A NAND2X1_LOC_451/Y 0.07fF
C72807 NAND2X1_LOC_454/Y NAND2X1_LOC_211/Y 0.07fF
C72808 INVX1_LOC_235/Y INVX1_LOC_169/Y 0.01fF
C72809 INVX1_LOC_24/Y NOR2X1_LOC_788/B 0.12fF
C72810 INVX1_LOC_178/A NAND2X1_LOC_560/A 0.23fF
C72811 INVX1_LOC_163/A NOR2X1_LOC_575/Y 0.11fF
C72812 INVX1_LOC_305/A INVX1_LOC_179/Y 0.01fF
C72813 INVX1_LOC_32/A NAND2X1_LOC_61/a_36_24# 0.00fF
C72814 INVX1_LOC_49/A NOR2X1_LOC_52/B 0.06fF
C72815 INVX1_LOC_45/A INVX1_LOC_290/A 0.07fF
C72816 NAND2X1_LOC_53/Y NOR2X1_LOC_214/B 0.04fF
C72817 INVX1_LOC_91/A NOR2X1_LOC_717/A 0.10fF
C72818 INPUT_3 NOR2X1_LOC_99/B 0.07fF
C72819 INVX1_LOC_27/A NOR2X1_LOC_74/A 0.17fF
C72820 INVX1_LOC_11/A INPUT_1 0.06fF
C72821 INVX1_LOC_5/A INVX1_LOC_201/A 0.01fF
C72822 VDD INVX1_LOC_23/Y 1.82fF
C72823 NAND2X1_LOC_541/Y INVX1_LOC_24/A 0.02fF
C72824 NOR2X1_LOC_68/A NOR2X1_LOC_516/B 0.03fF
C72825 INVX1_LOC_2/A NOR2X1_LOC_433/A 1.43fF
C72826 INVX1_LOC_269/A NAND2X1_LOC_323/a_36_24# 0.00fF
C72827 VDD NOR2X1_LOC_342/B 0.21fF
C72828 NAND2X1_LOC_364/A INVX1_LOC_1/Y 0.04fF
C72829 NOR2X1_LOC_340/Y INVX1_LOC_158/A 0.12fF
C72830 NAND2X1_LOC_475/Y INVX1_LOC_19/A 0.01fF
C72831 NOR2X1_LOC_155/A INVX1_LOC_42/A 0.00fF
C72832 INVX1_LOC_48/A NOR2X1_LOC_849/A 0.01fF
C72833 INVX1_LOC_17/A NOR2X1_LOC_329/B 0.15fF
C72834 INVX1_LOC_27/A NOR2X1_LOC_9/Y 0.10fF
C72835 NOR2X1_LOC_144/Y INVX1_LOC_85/A 0.12fF
C72836 NOR2X1_LOC_794/B INVX1_LOC_313/Y 0.07fF
C72837 INVX1_LOC_284/Y NOR2X1_LOC_576/B 0.02fF
C72838 INVX1_LOC_2/A NOR2X1_LOC_593/Y 0.01fF
C72839 NOR2X1_LOC_509/A NOR2X1_LOC_814/A 0.04fF
C72840 NOR2X1_LOC_226/A NOR2X1_LOC_433/A 0.08fF
C72841 NOR2X1_LOC_380/a_36_216# NAND2X1_LOC_866/B 0.00fF
C72842 INVX1_LOC_21/A INVX1_LOC_286/A 0.16fF
C72843 NOR2X1_LOC_596/A NAND2X1_LOC_831/a_36_24# 0.00fF
C72844 NOR2X1_LOC_78/B NOR2X1_LOC_716/B 0.07fF
C72845 INVX1_LOC_17/A D_INPUT_4 0.01fF
C72846 NOR2X1_LOC_226/A NOR2X1_LOC_593/Y 0.03fF
C72847 NOR2X1_LOC_287/A INVX1_LOC_77/A 0.05fF
C72848 INVX1_LOC_209/Y NAND2X1_LOC_852/Y 0.00fF
C72849 NAND2X1_LOC_483/Y NAND2X1_LOC_374/Y 0.03fF
C72850 INVX1_LOC_2/A INVX1_LOC_151/A 0.04fF
C72851 INVX1_LOC_133/Y INVX1_LOC_104/A 0.01fF
C72852 NOR2X1_LOC_272/Y NOR2X1_LOC_318/B 0.39fF
C72853 NOR2X1_LOC_209/Y NOR2X1_LOC_718/B 0.02fF
C72854 NOR2X1_LOC_218/Y NOR2X1_LOC_433/A 0.02fF
C72855 INPUT_3 NOR2X1_LOC_381/a_36_216# 0.00fF
C72856 INVX1_LOC_2/A NOR2X1_LOC_52/B 0.63fF
C72857 NOR2X1_LOC_114/Y NOR2X1_LOC_814/A 0.01fF
C72858 NOR2X1_LOC_802/A NAND2X1_LOC_118/a_36_24# 0.00fF
C72859 INVX1_LOC_230/Y INVX1_LOC_75/A 0.07fF
C72860 NOR2X1_LOC_272/Y INVX1_LOC_93/Y 0.10fF
C72861 NOR2X1_LOC_226/A NOR2X1_LOC_52/B 0.43fF
C72862 INVX1_LOC_119/A INVX1_LOC_144/Y 0.11fF
C72863 NAND2X1_LOC_308/Y NOR2X1_LOC_773/Y 0.02fF
C72864 INVX1_LOC_272/A NAND2X1_LOC_74/B 0.07fF
C72865 NOR2X1_LOC_808/A NOR2X1_LOC_806/Y 0.00fF
C72866 INVX1_LOC_21/A INVX1_LOC_95/A 0.03fF
C72867 NOR2X1_LOC_38/B INVX1_LOC_123/Y 0.03fF
C72868 INVX1_LOC_232/Y NAND2X1_LOC_141/A 0.01fF
C72869 INVX1_LOC_103/Y INVX1_LOC_22/A 0.01fF
C72870 INVX1_LOC_11/A NOR2X1_LOC_706/Y 0.01fF
C72871 NAND2X1_LOC_854/B NOR2X1_LOC_753/Y 0.05fF
C72872 NOR2X1_LOC_89/A NAND2X1_LOC_63/Y 0.77fF
C72873 INVX1_LOC_78/A NOR2X1_LOC_155/A 0.19fF
C72874 NOR2X1_LOC_474/A NAND2X1_LOC_462/B 0.02fF
C72875 NOR2X1_LOC_716/B NAND2X1_LOC_392/Y 0.01fF
C72876 D_INPUT_0 INVX1_LOC_314/Y 0.07fF
C72877 NOR2X1_LOC_143/a_36_216# INVX1_LOC_316/Y 0.00fF
C72878 NOR2X1_LOC_175/B INVX1_LOC_149/A 0.02fF
C72879 INVX1_LOC_110/Y INPUT_0 0.07fF
C72880 INVX1_LOC_94/A NAND2X1_LOC_492/a_36_24# 0.01fF
C72881 NOR2X1_LOC_218/Y NOR2X1_LOC_52/B 0.16fF
C72882 NAND2X1_LOC_53/Y NOR2X1_LOC_741/A 0.03fF
C72883 NOR2X1_LOC_780/A INVX1_LOC_75/A 0.01fF
C72884 NAND2X1_LOC_74/B NOR2X1_LOC_76/B 0.05fF
C72885 INVX1_LOC_15/Y INVX1_LOC_197/Y 0.01fF
C72886 NOR2X1_LOC_454/Y INVX1_LOC_187/Y 0.02fF
C72887 NOR2X1_LOC_596/A D_GATE_366 0.51fF
C72888 INVX1_LOC_18/A NOR2X1_LOC_567/B 0.42fF
C72889 NAND2X1_LOC_796/B NOR2X1_LOC_280/Y 0.06fF
C72890 NOR2X1_LOC_89/A NAND2X1_LOC_455/B 0.09fF
C72891 VDD NOR2X1_LOC_249/Y 0.34fF
C72892 NOR2X1_LOC_80/Y INVX1_LOC_84/A 0.19fF
C72893 VDD NOR2X1_LOC_846/A 0.00fF
C72894 NOR2X1_LOC_382/Y INPUT_0 0.01fF
C72895 INVX1_LOC_258/A NOR2X1_LOC_396/Y 0.02fF
C72896 NOR2X1_LOC_519/a_36_216# NOR2X1_LOC_48/B 0.00fF
C72897 NOR2X1_LOC_433/A NAND2X1_LOC_648/A 0.75fF
C72898 NOR2X1_LOC_65/B NOR2X1_LOC_155/A 0.07fF
C72899 NOR2X1_LOC_96/a_36_216# NOR2X1_LOC_392/Y 0.01fF
C72900 NOR2X1_LOC_68/A NOR2X1_LOC_706/A 0.00fF
C72901 NOR2X1_LOC_433/A INPUT_1 0.01fF
C72902 NAND2X1_LOC_555/Y NAND2X1_LOC_4/a_36_24# 0.01fF
C72903 INVX1_LOC_31/A INVX1_LOC_123/A 0.15fF
C72904 NOR2X1_LOC_620/Y INVX1_LOC_90/A 0.05fF
C72905 NOR2X1_LOC_754/A NAND2X1_LOC_254/Y 0.00fF
C72906 NOR2X1_LOC_89/A INVX1_LOC_257/A 0.04fF
C72907 INVX1_LOC_12/Y NAND2X1_LOC_474/Y 0.10fF
C72908 NOR2X1_LOC_591/A INVX1_LOC_92/A 0.01fF
C72909 INVX1_LOC_237/Y NOR2X1_LOC_575/Y 0.00fF
C72910 INVX1_LOC_64/A NOR2X1_LOC_332/Y 0.01fF
C72911 INVX1_LOC_33/A NOR2X1_LOC_738/A 0.02fF
C72912 INVX1_LOC_269/A INVX1_LOC_178/Y 0.24fF
C72913 INVX1_LOC_84/A INVX1_LOC_28/Y 0.01fF
C72914 NOR2X1_LOC_123/B NOR2X1_LOC_84/Y 0.16fF
C72915 NOR2X1_LOC_388/Y INVX1_LOC_28/A 0.42fF
C72916 NOR2X1_LOC_15/Y INVX1_LOC_129/Y 0.00fF
C72917 INVX1_LOC_249/A NOR2X1_LOC_74/A 0.03fF
C72918 NOR2X1_LOC_52/B INPUT_1 0.10fF
C72919 NAND2X1_LOC_479/Y INVX1_LOC_16/A 0.03fF
C72920 INVX1_LOC_11/A NOR2X1_LOC_586/Y 0.02fF
C72921 INVX1_LOC_21/A NOR2X1_LOC_602/B 0.06fF
C72922 INVX1_LOC_144/A NOR2X1_LOC_152/Y 0.07fF
C72923 NOR2X1_LOC_717/B NOR2X1_LOC_78/B 0.03fF
C72924 INVX1_LOC_64/A INVX1_LOC_179/A 0.01fF
C72925 INVX1_LOC_282/A NAND2X1_LOC_632/B 0.03fF
C72926 INVX1_LOC_33/A INVX1_LOC_73/A 0.00fF
C72927 NOR2X1_LOC_75/Y INVX1_LOC_46/A 0.01fF
C72928 INVX1_LOC_256/A INVX1_LOC_14/Y 0.07fF
C72929 NOR2X1_LOC_446/A VDD 0.00fF
C72930 NOR2X1_LOC_516/B NOR2X1_LOC_545/a_36_216# 0.13fF
C72931 INVX1_LOC_21/A INVX1_LOC_54/A 0.15fF
C72932 NAND2X1_LOC_303/Y NOR2X1_LOC_536/A 0.12fF
C72933 NOR2X1_LOC_647/B D_INPUT_3 0.01fF
C72934 INVX1_LOC_209/A INVX1_LOC_173/Y 0.28fF
C72935 INVX1_LOC_206/A NOR2X1_LOC_356/A 0.03fF
C72936 INVX1_LOC_164/A INVX1_LOC_22/A 0.01fF
C72937 NOR2X1_LOC_441/Y NOR2X1_LOC_279/Y 0.01fF
C72938 INVX1_LOC_233/A NAND2X1_LOC_572/B 0.28fF
C72939 NOR2X1_LOC_716/B NOR2X1_LOC_193/a_36_216# 0.00fF
C72940 NAND2X1_LOC_519/a_36_24# INVX1_LOC_77/A 0.01fF
C72941 NOR2X1_LOC_596/Y VDD 0.23fF
C72942 NOR2X1_LOC_78/B NOR2X1_LOC_828/A 0.01fF
C72943 NAND2X1_LOC_364/A INVX1_LOC_93/Y 0.26fF
C72944 NOR2X1_LOC_353/a_36_216# INVX1_LOC_78/Y 0.00fF
C72945 NAND2X1_LOC_513/B INVX1_LOC_274/A 0.02fF
C72946 NOR2X1_LOC_216/B INVX1_LOC_306/Y 0.09fF
C72947 INVX1_LOC_135/A INVX1_LOC_16/A 0.14fF
C72948 INVX1_LOC_24/A NOR2X1_LOC_78/A 0.07fF
C72949 NAND2X1_LOC_860/A NOR2X1_LOC_662/A 0.03fF
C72950 NOR2X1_LOC_13/Y INVX1_LOC_91/A 0.08fF
C72951 INVX1_LOC_47/Y INVX1_LOC_4/Y 0.01fF
C72952 NOR2X1_LOC_705/B INVX1_LOC_117/A 0.03fF
C72953 INVX1_LOC_284/Y NOR2X1_LOC_492/a_36_216# 0.01fF
C72954 NOR2X1_LOC_782/a_36_216# INVX1_LOC_91/A 0.00fF
C72955 NOR2X1_LOC_627/Y NOR2X1_LOC_742/A 0.03fF
C72956 INVX1_LOC_279/A NAND2X1_LOC_715/a_36_24# 0.02fF
C72957 NAND2X1_LOC_787/A INVX1_LOC_19/A 0.08fF
C72958 NAND2X1_LOC_741/B VDD 0.39fF
C72959 NAND2X1_LOC_223/B NAND2X1_LOC_223/a_36_24# 0.00fF
C72960 INVX1_LOC_27/A NOR2X1_LOC_865/Y 0.03fF
C72961 INVX1_LOC_206/A NOR2X1_LOC_74/A 0.00fF
C72962 INVX1_LOC_14/A INVX1_LOC_185/A 0.08fF
C72963 NOR2X1_LOC_778/Y INVX1_LOC_37/A 0.03fF
C72964 INVX1_LOC_11/A INVX1_LOC_118/A 0.15fF
C72965 NAND2X1_LOC_363/B INVX1_LOC_19/A 0.10fF
C72966 NOR2X1_LOC_78/B NOR2X1_LOC_151/Y 0.03fF
C72967 INVX1_LOC_27/A NOR2X1_LOC_243/B 0.03fF
C72968 INVX1_LOC_246/A NOR2X1_LOC_331/B 0.79fF
C72969 INVX1_LOC_1/A NOR2X1_LOC_79/a_36_216# 0.00fF
C72970 NOR2X1_LOC_82/A INVX1_LOC_127/A 0.01fF
C72971 NOR2X1_LOC_551/Y INVX1_LOC_104/A 0.05fF
C72972 INVX1_LOC_83/A NOR2X1_LOC_326/Y 0.10fF
C72973 NOR2X1_LOC_717/B INVX1_LOC_83/A 0.16fF
C72974 INVX1_LOC_103/A NOR2X1_LOC_358/a_36_216# 0.00fF
C72975 INVX1_LOC_77/A INVX1_LOC_95/Y 0.07fF
C72976 NOR2X1_LOC_188/A NOR2X1_LOC_537/Y 0.07fF
C72977 NAND2X1_LOC_338/B NOR2X1_LOC_188/A 0.07fF
C72978 NOR2X1_LOC_714/Y NOR2X1_LOC_704/Y 0.08fF
C72979 INVX1_LOC_24/A NAND2X1_LOC_464/A 0.00fF
C72980 INVX1_LOC_36/A NOR2X1_LOC_440/a_36_216# 0.01fF
C72981 NOR2X1_LOC_256/Y INVX1_LOC_25/Y 0.02fF
C72982 NOR2X1_LOC_520/A INVX1_LOC_51/Y 0.14fF
C72983 NOR2X1_LOC_548/B NOR2X1_LOC_537/Y 0.03fF
C72984 NOR2X1_LOC_202/Y INVX1_LOC_16/A 0.01fF
C72985 INVX1_LOC_269/A NOR2X1_LOC_445/B 2.12fF
C72986 NAND2X1_LOC_338/B NOR2X1_LOC_548/B 0.04fF
C72987 INVX1_LOC_270/A INVX1_LOC_15/A 0.14fF
C72988 INVX1_LOC_90/Y INVX1_LOC_175/A 0.00fF
C72989 NAND2X1_LOC_552/A INVX1_LOC_29/A 0.02fF
C72990 INVX1_LOC_5/A INVX1_LOC_29/A 0.26fF
C72991 INVX1_LOC_88/A NOR2X1_LOC_117/a_36_216# 0.12fF
C72992 INVX1_LOC_314/Y NOR2X1_LOC_266/B 0.03fF
C72993 NOR2X1_LOC_355/B NOR2X1_LOC_493/B 0.20fF
C72994 NOR2X1_LOC_352/Y INVX1_LOC_78/Y 0.42fF
C72995 NOR2X1_LOC_122/A NAND2X1_LOC_475/Y 0.01fF
C72996 INVX1_LOC_135/A INVX1_LOC_28/A 0.19fF
C72997 NOR2X1_LOC_419/Y NOR2X1_LOC_98/A -0.01fF
C72998 INVX1_LOC_246/A NOR2X1_LOC_592/B 0.09fF
C72999 INVX1_LOC_174/A NAND2X1_LOC_50/a_36_24# 0.01fF
C73000 NAND2X1_LOC_579/A NAND2X1_LOC_489/Y 0.05fF
C73001 NOR2X1_LOC_716/B INVX1_LOC_46/A 0.27fF
C73002 INVX1_LOC_143/A NOR2X1_LOC_78/A 0.08fF
C73003 INVX1_LOC_215/Y NOR2X1_LOC_841/A 0.09fF
C73004 NOR2X1_LOC_802/A NOR2X1_LOC_542/B 0.06fF
C73005 NOR2X1_LOC_52/Y INVX1_LOC_157/Y -0.01fF
C73006 NOR2X1_LOC_97/A NOR2X1_LOC_97/B 0.00fF
C73007 NAND2X1_LOC_354/Y INVX1_LOC_54/A 0.02fF
C73008 INVX1_LOC_21/A NAND2X1_LOC_807/B 0.07fF
C73009 INVX1_LOC_2/A INVX1_LOC_199/A 0.02fF
C73010 NOR2X1_LOC_109/Y INVX1_LOC_15/A 0.07fF
C73011 INVX1_LOC_161/Y NAND2X1_LOC_475/Y 0.10fF
C73012 INVX1_LOC_265/A INVX1_LOC_37/A 0.05fF
C73013 NAND2X1_LOC_9/Y NOR2X1_LOC_394/Y 0.30fF
C73014 NOR2X1_LOC_360/Y NOR2X1_LOC_860/Y 0.04fF
C73015 NAND2X1_LOC_74/B NOR2X1_LOC_271/B 0.01fF
C73016 INVX1_LOC_218/A NAND2X1_LOC_642/Y 0.03fF
C73017 NOR2X1_LOC_598/B INVX1_LOC_78/A 0.76fF
C73018 INVX1_LOC_21/A NOR2X1_LOC_48/B 0.18fF
C73019 NAND2X1_LOC_116/A VDD 0.35fF
C73020 NOR2X1_LOC_504/Y NOR2X1_LOC_421/Y 0.13fF
C73021 NOR2X1_LOC_146/Y INVX1_LOC_91/A 0.01fF
C73022 NAND2X1_LOC_726/Y NAND2X1_LOC_729/B 0.11fF
C73023 NOR2X1_LOC_147/B INVX1_LOC_117/A 0.06fF
C73024 NOR2X1_LOC_180/Y INVX1_LOC_37/A 0.03fF
C73025 INVX1_LOC_224/A NAND2X1_LOC_63/Y 0.01fF
C73026 NAND2X1_LOC_286/B INVX1_LOC_57/A 0.17fF
C73027 INVX1_LOC_269/A INVX1_LOC_12/A 0.28fF
C73028 NOR2X1_LOC_639/B NOR2X1_LOC_158/Y 0.46fF
C73029 INVX1_LOC_1/Y NOR2X1_LOC_113/A 0.03fF
C73030 NOR2X1_LOC_392/B INVX1_LOC_117/A 0.01fF
C73031 NOR2X1_LOC_332/A INVX1_LOC_201/A 0.02fF
C73032 INVX1_LOC_1/Y NOR2X1_LOC_405/A 0.14fF
C73033 INVX1_LOC_11/A NAND2X1_LOC_63/Y 0.12fF
C73034 NOR2X1_LOC_468/Y INVX1_LOC_102/A 0.01fF
C73035 NOR2X1_LOC_690/A NOR2X1_LOC_536/A 0.14fF
C73036 NOR2X1_LOC_433/A INVX1_LOC_118/A 0.13fF
C73037 INVX1_LOC_89/A INVX1_LOC_92/Y 0.01fF
C73038 NOR2X1_LOC_191/A INVX1_LOC_76/A 0.02fF
C73039 D_INPUT_6 D_INPUT_5 0.11fF
C73040 INVX1_LOC_35/A NOR2X1_LOC_301/A 0.04fF
C73041 NAND2X1_LOC_715/B INVX1_LOC_78/A 0.07fF
C73042 INVX1_LOC_30/A NOR2X1_LOC_653/Y 0.02fF
C73043 NAND2X1_LOC_337/B INVX1_LOC_29/A 0.07fF
C73044 NOR2X1_LOC_284/B VDD -0.00fF
C73045 INVX1_LOC_25/A INVX1_LOC_224/Y 1.44fF
C73046 INVX1_LOC_36/A INVX1_LOC_84/A 0.32fF
C73047 NAND2X1_LOC_363/B INVX1_LOC_26/Y 0.07fF
C73048 NOR2X1_LOC_276/Y INVX1_LOC_272/A 0.03fF
C73049 INVX1_LOC_314/Y INVX1_LOC_46/Y -0.04fF
C73050 D_INPUT_0 NOR2X1_LOC_557/A 0.01fF
C73051 INVX1_LOC_236/Y INVX1_LOC_49/Y 0.01fF
C73052 INVX1_LOC_64/A NOR2X1_LOC_693/Y 0.05fF
C73053 INVX1_LOC_57/A NOR2X1_LOC_15/a_36_216# 0.00fF
C73054 D_INPUT_1 INVX1_LOC_23/A 0.29fF
C73055 INVX1_LOC_298/Y INVX1_LOC_5/A 0.07fF
C73056 NAND2X1_LOC_860/A INVX1_LOC_57/A 0.03fF
C73057 NOR2X1_LOC_152/Y NOR2X1_LOC_155/A 0.01fF
C73058 INVX1_LOC_170/A NAND2X1_LOC_773/B 0.03fF
C73059 INVX1_LOC_255/Y INVX1_LOC_20/A 0.04fF
C73060 NOR2X1_LOC_254/Y INVX1_LOC_274/A 0.07fF
C73061 NOR2X1_LOC_34/B NOR2X1_LOC_34/Y 0.03fF
C73062 INVX1_LOC_30/A INVX1_LOC_19/A 1.40fF
C73063 INVX1_LOC_232/A VDD 1.83fF
C73064 INVX1_LOC_57/A NOR2X1_LOC_634/Y 0.04fF
C73065 NOR2X1_LOC_52/B INVX1_LOC_118/A 0.37fF
C73066 NOR2X1_LOC_68/A NOR2X1_LOC_605/A 0.01fF
C73067 NAND2X1_LOC_785/Y INVX1_LOC_54/A 0.01fF
C73068 INVX1_LOC_16/A INVX1_LOC_139/Y 0.03fF
C73069 INVX1_LOC_30/A NOR2X1_LOC_11/Y 0.16fF
C73070 NAND2X1_LOC_763/B INVX1_LOC_19/A 0.14fF
C73071 NOR2X1_LOC_134/Y NAND2X1_LOC_254/Y 1.38fF
C73072 INVX1_LOC_226/Y INVX1_LOC_12/Y 0.03fF
C73073 NOR2X1_LOC_471/Y NOR2X1_LOC_477/B 0.03fF
C73074 NOR2X1_LOC_576/B NAND2X1_LOC_853/a_36_24# 0.01fF
C73075 NOR2X1_LOC_372/A INVX1_LOC_42/A 0.00fF
C73076 INVX1_LOC_21/A NOR2X1_LOC_438/Y 0.03fF
C73077 NOR2X1_LOC_208/Y INVX1_LOC_84/A 0.09fF
C73078 NOR2X1_LOC_428/Y NOR2X1_LOC_48/B 0.08fF
C73079 NOR2X1_LOC_590/A NOR2X1_LOC_114/Y 0.22fF
C73080 NOR2X1_LOC_383/Y VDD 0.56fF
C73081 INVX1_LOC_196/A INVX1_LOC_9/A 0.10fF
C73082 INVX1_LOC_136/A INVX1_LOC_272/A 0.10fF
C73083 NOR2X1_LOC_437/Y NAND2X1_LOC_475/Y 0.10fF
C73084 NOR2X1_LOC_219/Y INVX1_LOC_281/A 0.02fF
C73085 NAND2X1_LOC_633/Y NAND2X1_LOC_392/Y 0.11fF
C73086 INVX1_LOC_100/A NOR2X1_LOC_368/A 0.08fF
C73087 NOR2X1_LOC_598/B INVX1_LOC_152/Y 0.01fF
C73088 NOR2X1_LOC_667/A NOR2X1_LOC_602/B 0.14fF
C73089 NAND2X1_LOC_564/B NOR2X1_LOC_176/Y 0.00fF
C73090 NOR2X1_LOC_813/Y INVX1_LOC_16/A 0.15fF
C73091 NAND2X1_LOC_721/A NOR2X1_LOC_86/A 0.05fF
C73092 INVX1_LOC_135/A NOR2X1_LOC_35/Y 0.05fF
C73093 NAND2X1_LOC_218/B NAND2X1_LOC_225/a_36_24# 0.00fF
C73094 INVX1_LOC_248/A NOR2X1_LOC_602/B 0.01fF
C73095 INVX1_LOC_50/A NAND2X1_LOC_169/Y 0.18fF
C73096 NOR2X1_LOC_237/Y INVX1_LOC_84/A 0.07fF
C73097 INVX1_LOC_121/A NOR2X1_LOC_145/Y 0.02fF
C73098 NAND2X1_LOC_579/A NAND2X1_LOC_175/Y 0.04fF
C73099 NOR2X1_LOC_71/Y INVX1_LOC_20/A 0.25fF
C73100 INVX1_LOC_10/Y INVX1_LOC_16/A 0.03fF
C73101 NOR2X1_LOC_366/Y VDD 0.44fF
C73102 NOR2X1_LOC_717/B INVX1_LOC_46/A 0.03fF
C73103 NOR2X1_LOC_92/Y NAND2X1_LOC_61/Y 0.07fF
C73104 NOR2X1_LOC_667/A INVX1_LOC_54/A 0.07fF
C73105 NOR2X1_LOC_68/A NAND2X1_LOC_207/B 0.19fF
C73106 INVX1_LOC_248/A INVX1_LOC_54/A 0.07fF
C73107 INVX1_LOC_23/A NOR2X1_LOC_652/Y 0.07fF
C73108 INVX1_LOC_10/A INVX1_LOC_12/Y 0.01fF
C73109 INVX1_LOC_16/A INVX1_LOC_280/A 0.45fF
C73110 NOR2X1_LOC_217/a_36_216# NAND2X1_LOC_454/Y 0.01fF
C73111 NAND2X1_LOC_656/a_36_24# INVX1_LOC_46/A 0.01fF
C73112 INVX1_LOC_136/A NOR2X1_LOC_76/B 0.07fF
C73113 NOR2X1_LOC_528/Y NOR2X1_LOC_74/A 0.10fF
C73114 NOR2X1_LOC_478/a_36_216# INVX1_LOC_117/A 0.00fF
C73115 NOR2X1_LOC_112/B NOR2X1_LOC_78/A 0.26fF
C73116 INVX1_LOC_8/A INVX1_LOC_27/Y 0.04fF
C73117 NAND2X1_LOC_703/Y NOR2X1_LOC_654/A 0.10fF
C73118 NOR2X1_LOC_361/B INVX1_LOC_23/Y 0.10fF
C73119 INVX1_LOC_90/A NOR2X1_LOC_314/Y 0.01fF
C73120 INVX1_LOC_90/A NOR2X1_LOC_422/Y 0.04fF
C73121 INVX1_LOC_290/A NOR2X1_LOC_331/B 0.01fF
C73122 INVX1_LOC_266/Y INVX1_LOC_113/A 0.01fF
C73123 NAND2X1_LOC_354/Y NOR2X1_LOC_48/B 0.12fF
C73124 NOR2X1_LOC_337/A INVX1_LOC_91/A 0.04fF
C73125 INVX1_LOC_45/A NOR2X1_LOC_467/A 0.14fF
C73126 NOR2X1_LOC_297/a_36_216# NAND2X1_LOC_206/Y 0.01fF
C73127 INVX1_LOC_11/A NOR2X1_LOC_631/Y 0.08fF
C73128 NAND2X1_LOC_795/Y NOR2X1_LOC_692/a_36_216# 0.00fF
C73129 NOR2X1_LOC_582/Y NOR2X1_LOC_48/B 0.16fF
C73130 INVX1_LOC_36/A INVX1_LOC_15/A 3.13fF
C73131 NOR2X1_LOC_309/Y INVX1_LOC_84/A 0.07fF
C73132 INVX1_LOC_240/A NOR2X1_LOC_485/Y 0.03fF
C73133 INVX1_LOC_224/Y INVX1_LOC_1/A 0.10fF
C73134 INVX1_LOC_177/A INVX1_LOC_220/A 0.01fF
C73135 NAND2X1_LOC_537/Y INVX1_LOC_57/A 0.07fF
C73136 NOR2X1_LOC_775/Y VDD 0.19fF
C73137 NOR2X1_LOC_625/Y INVX1_LOC_284/A 0.01fF
C73138 INVX1_LOC_90/A INVX1_LOC_117/A 0.17fF
C73139 INVX1_LOC_161/Y NOR2X1_LOC_135/a_36_216# 0.01fF
C73140 NOR2X1_LOC_322/Y NAND2X1_LOC_244/A 0.00fF
C73141 INVX1_LOC_103/A INVX1_LOC_29/Y 0.02fF
C73142 NOR2X1_LOC_151/Y INVX1_LOC_46/A 0.03fF
C73143 INVX1_LOC_83/A NOR2X1_LOC_209/B 0.07fF
C73144 INVX1_LOC_286/A INVX1_LOC_304/A 0.11fF
C73145 INVX1_LOC_25/A NOR2X1_LOC_103/Y 0.07fF
C73146 INVX1_LOC_28/A NOR2X1_LOC_152/A 0.09fF
C73147 INVX1_LOC_94/A NOR2X1_LOC_609/Y 0.04fF
C73148 NOR2X1_LOC_91/Y NAND2X1_LOC_444/B 0.01fF
C73149 INVX1_LOC_71/A NOR2X1_LOC_467/A 1.22fF
C73150 NOR2X1_LOC_318/B NOR2X1_LOC_405/A 0.02fF
C73151 INVX1_LOC_230/Y NOR2X1_LOC_529/a_36_216# 0.01fF
C73152 NAND2X1_LOC_364/A INVX1_LOC_87/A -0.02fF
C73153 NOR2X1_LOC_237/Y INVX1_LOC_15/A 0.07fF
C73154 INVX1_LOC_30/A INVX1_LOC_26/Y 0.71fF
C73155 INVX1_LOC_35/A INVX1_LOC_17/A 0.14fF
C73156 INVX1_LOC_292/A INVX1_LOC_29/Y 0.04fF
C73157 INVX1_LOC_75/A INVX1_LOC_44/A 0.07fF
C73158 INVX1_LOC_89/A NOR2X1_LOC_259/A 0.00fF
C73159 INVX1_LOC_18/A INVX1_LOC_26/A 0.01fF
C73160 D_INPUT_1 INVX1_LOC_31/A 0.20fF
C73161 NAND2X1_LOC_360/a_36_24# NOR2X1_LOC_103/Y 0.00fF
C73162 NAND2X1_LOC_785/Y NOR2X1_LOC_48/B -0.00fF
C73163 INVX1_LOC_95/A INVX1_LOC_304/A 0.01fF
C73164 NOR2X1_LOC_632/Y INVX1_LOC_136/Y 0.00fF
C73165 NOR2X1_LOC_474/A NAND2X1_LOC_618/Y 0.02fF
C73166 NOR2X1_LOC_513/a_36_216# INVX1_LOC_78/A 0.00fF
C73167 NAND2X1_LOC_557/Y INVX1_LOC_30/A 0.01fF
C73168 INVX1_LOC_222/Y INVX1_LOC_299/A 0.02fF
C73169 NOR2X1_LOC_392/B INVX1_LOC_3/Y 0.10fF
C73170 INVX1_LOC_77/A INVX1_LOC_271/Y 0.03fF
C73171 NOR2X1_LOC_773/Y INVX1_LOC_29/A 0.08fF
C73172 INVX1_LOC_2/A NAND2X1_LOC_254/Y 0.03fF
C73173 NOR2X1_LOC_552/A NOR2X1_LOC_35/Y 0.10fF
C73174 INVX1_LOC_35/A NAND2X1_LOC_555/Y 0.09fF
C73175 INVX1_LOC_186/A VDD 0.21fF
C73176 NOR2X1_LOC_309/Y INVX1_LOC_15/A 0.07fF
C73177 NAND2X1_LOC_563/A INVX1_LOC_12/A 0.26fF
C73178 NOR2X1_LOC_669/a_36_216# NOR2X1_LOC_669/Y 0.02fF
C73179 INVX1_LOC_39/A INVX1_LOC_11/A 0.03fF
C73180 INVX1_LOC_25/A NOR2X1_LOC_819/a_36_216# 0.02fF
C73181 INVX1_LOC_214/A NOR2X1_LOC_48/B 0.01fF
C73182 NAND2X1_LOC_51/B INVX1_LOC_54/A 0.03fF
C73183 INVX1_LOC_108/Y INVX1_LOC_36/A 0.04fF
C73184 NOR2X1_LOC_667/A NOR2X1_LOC_48/B 0.56fF
C73185 NOR2X1_LOC_769/A NOR2X1_LOC_598/B 0.01fF
C73186 INVX1_LOC_248/A NOR2X1_LOC_48/B 0.08fF
C73187 INVX1_LOC_278/A INVX1_LOC_36/A 0.05fF
C73188 NAND2X1_LOC_466/Y NAND2X1_LOC_470/B 0.02fF
C73189 NOR2X1_LOC_598/B NOR2X1_LOC_554/B 1.72fF
C73190 INVX1_LOC_21/A NAND2X1_LOC_350/A 0.07fF
C73191 INVX1_LOC_74/Y VDD 0.21fF
C73192 INVX1_LOC_245/Y INVX1_LOC_27/A 0.02fF
C73193 INVX1_LOC_311/A INVX1_LOC_54/A 0.11fF
C73194 NOR2X1_LOC_244/B NAND2X1_LOC_232/a_36_24# 0.01fF
C73195 VDD NAND2X1_LOC_447/Y 1.24fF
C73196 NOR2X1_LOC_160/B NAND2X1_LOC_474/Y 0.07fF
C73197 NOR2X1_LOC_635/a_36_216# NOR2X1_LOC_68/A 0.00fF
C73198 NOR2X1_LOC_366/a_36_216# NOR2X1_LOC_139/Y 0.00fF
C73199 NOR2X1_LOC_403/B INVX1_LOC_23/A 0.04fF
C73200 INVX1_LOC_1/A NOR2X1_LOC_103/Y 0.10fF
C73201 INVX1_LOC_50/A NOR2X1_LOC_387/Y 0.06fF
C73202 INVX1_LOC_25/A INVX1_LOC_71/A 0.17fF
C73203 D_INPUT_2 INVX1_LOC_23/A 0.70fF
C73204 INVX1_LOC_269/A INVX1_LOC_228/Y 0.03fF
C73205 NOR2X1_LOC_443/Y NAND2X1_LOC_361/Y 0.03fF
C73206 INVX1_LOC_21/A NOR2X1_LOC_441/Y 0.07fF
C73207 NOR2X1_LOC_74/A NOR2X1_LOC_216/B 0.10fF
C73208 NOR2X1_LOC_332/A INVX1_LOC_29/A 0.07fF
C73209 NOR2X1_LOC_156/B INVX1_LOC_78/A 0.01fF
C73210 NAND2X1_LOC_552/A NAND2X1_LOC_634/Y 0.02fF
C73211 NAND2X1_LOC_796/B INVX1_LOC_286/Y 0.10fF
C73212 NAND2X1_LOC_660/A INVX1_LOC_78/A 2.03fF
C73213 INVX1_LOC_27/A INVX1_LOC_124/Y 0.01fF
C73214 INVX1_LOC_247/Y INVX1_LOC_5/A 0.01fF
C73215 INVX1_LOC_208/Y INVX1_LOC_32/A 0.08fF
C73216 NAND2X1_LOC_633/Y INVX1_LOC_46/A 0.07fF
C73217 INVX1_LOC_64/A INVX1_LOC_45/Y 0.01fF
C73218 NOR2X1_LOC_434/Y INVX1_LOC_305/A 0.04fF
C73219 NAND2X1_LOC_284/a_36_24# INVX1_LOC_20/A 0.01fF
C73220 NAND2X1_LOC_477/A NAND2X1_LOC_61/Y 0.05fF
C73221 NOR2X1_LOC_598/B NOR2X1_LOC_152/Y 0.01fF
C73222 NAND2X1_LOC_9/Y NOR2X1_LOC_419/Y 0.04fF
C73223 NOR2X1_LOC_740/Y NOR2X1_LOC_307/A 0.02fF
C73224 NOR2X1_LOC_9/Y NOR2X1_LOC_216/B 0.10fF
C73225 NOR2X1_LOC_315/Y NAND2X1_LOC_99/A 0.01fF
C73226 NAND2X1_LOC_721/B INVX1_LOC_178/A 0.01fF
C73227 INVX1_LOC_89/A INVX1_LOC_106/A 0.02fF
C73228 NOR2X1_LOC_214/B INVX1_LOC_12/A 0.08fF
C73229 INVX1_LOC_278/A NOR2X1_LOC_237/Y 1.39fF
C73230 INVX1_LOC_255/Y INVX1_LOC_4/A 0.04fF
C73231 NAND2X1_LOC_9/Y NOR2X1_LOC_716/B 0.08fF
C73232 INVX1_LOC_50/A NAND2X1_LOC_357/B 0.18fF
C73233 NAND2X1_LOC_53/Y NOR2X1_LOC_160/B 0.42fF
C73234 INVX1_LOC_233/A NOR2X1_LOC_716/B 0.17fF
C73235 INVX1_LOC_280/A NOR2X1_LOC_35/Y 0.10fF
C73236 NOR2X1_LOC_794/B NOR2X1_LOC_541/Y 0.00fF
C73237 NOR2X1_LOC_65/B NAND2X1_LOC_660/A 0.20fF
C73238 INVX1_LOC_304/A INVX1_LOC_54/A 0.02fF
C73239 INVX1_LOC_45/A INVX1_LOC_1/A 1.06fF
C73240 NOR2X1_LOC_373/Y INVX1_LOC_19/Y 0.05fF
C73241 NOR2X1_LOC_139/Y NOR2X1_LOC_364/A 1.23fF
C73242 NAND2X1_LOC_715/B NOR2X1_LOC_152/Y 0.10fF
C73243 NOR2X1_LOC_122/A INVX1_LOC_30/A 0.03fF
C73244 VDD INVX1_LOC_166/Y 0.25fF
C73245 NAND2X1_LOC_538/Y INVX1_LOC_141/Y 0.14fF
C73246 NOR2X1_LOC_773/Y NOR2X1_LOC_281/Y 0.03fF
C73247 INVX1_LOC_1/A NOR2X1_LOC_568/A 0.00fF
C73248 INPUT_1 NAND2X1_LOC_254/Y 0.07fF
C73249 NOR2X1_LOC_860/B INVX1_LOC_50/Y 0.07fF
C73250 INVX1_LOC_256/A NAND2X1_LOC_120/a_36_24# 0.00fF
C73251 NOR2X1_LOC_78/A NOR2X1_LOC_197/B 0.00fF
C73252 NAND2X1_LOC_538/Y INVX1_LOC_312/Y 0.29fF
C73253 NAND2X1_LOC_549/Y INVX1_LOC_219/Y 0.00fF
C73254 NOR2X1_LOC_272/a_36_216# NOR2X1_LOC_433/A 0.00fF
C73255 NOR2X1_LOC_798/A NOR2X1_LOC_537/A 0.00fF
C73256 NOR2X1_LOC_250/A INVX1_LOC_312/Y 0.02fF
C73257 NOR2X1_LOC_71/Y INVX1_LOC_4/A 0.01fF
C73258 INVX1_LOC_90/A INVX1_LOC_3/Y 0.39fF
C73259 NAND2X1_LOC_468/B NOR2X1_LOC_364/A 0.00fF
C73260 NAND2X1_LOC_243/Y INVX1_LOC_20/A 0.01fF
C73261 INVX1_LOC_161/Y INVX1_LOC_30/A 0.70fF
C73262 INVX1_LOC_38/A INVX1_LOC_117/A 0.21fF
C73263 INVX1_LOC_5/A INVX1_LOC_8/A 0.08fF
C73264 NAND2X1_LOC_666/a_36_24# INVX1_LOC_16/Y 0.00fF
C73265 NAND2X1_LOC_560/A INVX1_LOC_42/A 0.04fF
C73266 NOR2X1_LOC_186/Y NOR2X1_LOC_557/Y 0.04fF
C73267 NAND2X1_LOC_276/Y NOR2X1_LOC_649/Y 0.01fF
C73268 NAND2X1_LOC_214/B NOR2X1_LOC_121/Y 0.01fF
C73269 INVX1_LOC_182/Y INVX1_LOC_290/Y 0.14fF
C73270 NAND2X1_LOC_721/B NOR2X1_LOC_816/A -0.03fF
C73271 INVX1_LOC_299/A NAND2X1_LOC_656/A 0.17fF
C73272 INVX1_LOC_136/A INVX1_LOC_150/Y 0.08fF
C73273 INVX1_LOC_172/Y INVX1_LOC_57/A 0.01fF
C73274 INVX1_LOC_1/A INVX1_LOC_71/A 0.17fF
C73275 NOR2X1_LOC_644/A INVX1_LOC_4/A 0.03fF
C73276 NOR2X1_LOC_163/a_36_216# D_INPUT_5 0.00fF
C73277 INVX1_LOC_21/A NOR2X1_LOC_142/Y 0.01fF
C73278 NAND2X1_LOC_350/A NAND2X1_LOC_354/Y 0.01fF
C73279 NAND2X1_LOC_773/Y INVX1_LOC_77/A 0.09fF
C73280 INVX1_LOC_22/A NOR2X1_LOC_696/Y 0.22fF
C73281 NOR2X1_LOC_272/a_36_216# NOR2X1_LOC_52/B 0.01fF
C73282 NAND2X1_LOC_348/A INVX1_LOC_3/Y 0.05fF
C73283 NAND2X1_LOC_660/Y INVX1_LOC_271/A 0.16fF
C73284 NOR2X1_LOC_741/A INVX1_LOC_12/A 0.02fF
C73285 NOR2X1_LOC_329/B INVX1_LOC_94/Y 0.12fF
C73286 NOR2X1_LOC_794/B INVX1_LOC_71/A 0.03fF
C73287 INVX1_LOC_211/Y NOR2X1_LOC_447/Y 0.24fF
C73288 NAND2X1_LOC_51/B NAND2X1_LOC_3/B 0.23fF
C73289 NOR2X1_LOC_67/A INVX1_LOC_7/Y -0.03fF
C73290 NOR2X1_LOC_15/Y NOR2X1_LOC_6/B 0.02fF
C73291 INVX1_LOC_21/A NOR2X1_LOC_655/B 0.01fF
C73292 INVX1_LOC_302/Y NOR2X1_LOC_158/a_36_216# 0.00fF
C73293 INVX1_LOC_31/A D_INPUT_2 0.07fF
C73294 INVX1_LOC_24/A INVX1_LOC_170/A 0.01fF
C73295 NOR2X1_LOC_826/a_36_216# INVX1_LOC_135/A 0.01fF
C73296 INVX1_LOC_57/Y INVX1_LOC_41/Y 0.03fF
C73297 NOR2X1_LOC_180/B NOR2X1_LOC_748/A 0.10fF
C73298 INVX1_LOC_35/A NOR2X1_LOC_199/B 0.01fF
C73299 NOR2X1_LOC_381/Y NAND2X1_LOC_141/A 0.00fF
C73300 NOR2X1_LOC_437/Y INVX1_LOC_30/A 0.10fF
C73301 NOR2X1_LOC_67/A NOR2X1_LOC_92/Y 0.07fF
C73302 INVX1_LOC_58/A INVX1_LOC_90/A 0.56fF
C73303 INVX1_LOC_58/A NOR2X1_LOC_389/B 0.03fF
C73304 INVX1_LOC_146/A NOR2X1_LOC_654/A 0.05fF
C73305 INVX1_LOC_136/A NOR2X1_LOC_403/a_36_216# 0.02fF
C73306 INVX1_LOC_64/A NOR2X1_LOC_71/Y 0.02fF
C73307 INVX1_LOC_282/A NOR2X1_LOC_693/Y 0.07fF
C73308 NOR2X1_LOC_33/A INVX1_LOC_27/A 0.03fF
C73309 INVX1_LOC_230/Y NOR2X1_LOC_629/B 0.01fF
C73310 INVX1_LOC_172/Y NOR2X1_LOC_475/A 0.01fF
C73311 NOR2X1_LOC_446/A INVX1_LOC_177/A 0.01fF
C73312 INVX1_LOC_139/A INVX1_LOC_109/Y 0.02fF
C73313 NAND2X1_LOC_214/B D_INPUT_0 0.03fF
C73314 NOR2X1_LOC_465/a_36_216# NOR2X1_LOC_644/A 0.00fF
C73315 NOR2X1_LOC_186/Y NAND2X1_LOC_783/A 0.00fF
C73316 INVX1_LOC_14/Y NOR2X1_LOC_89/A 0.00fF
C73317 NAND2X1_LOC_564/B NAND2X1_LOC_579/A 0.01fF
C73318 INVX1_LOC_228/Y NAND2X1_LOC_563/A 0.07fF
C73319 INVX1_LOC_64/A NOR2X1_LOC_644/A 0.14fF
C73320 NOR2X1_LOC_186/Y NOR2X1_LOC_130/A 0.08fF
C73321 INVX1_LOC_12/Y INVX1_LOC_12/A 0.72fF
C73322 INVX1_LOC_244/Y NOR2X1_LOC_430/A 0.09fF
C73323 NOR2X1_LOC_271/Y NAND2X1_LOC_773/B 0.00fF
C73324 INVX1_LOC_45/A INVX1_LOC_221/A 0.03fF
C73325 NOR2X1_LOC_15/Y INVX1_LOC_30/Y 0.08fF
C73326 INVX1_LOC_21/A NOR2X1_LOC_99/B 0.12fF
C73327 INVX1_LOC_49/A NAND2X1_LOC_315/a_36_24# 0.00fF
C73328 NOR2X1_LOC_569/A NOR2X1_LOC_748/A 0.04fF
C73329 NOR2X1_LOC_772/B INVX1_LOC_87/Y 0.03fF
C73330 INVX1_LOC_132/A INVX1_LOC_24/A 0.07fF
C73331 INVX1_LOC_27/A D_INPUT_0 0.13fF
C73332 INVX1_LOC_83/A NAND2X1_LOC_816/a_36_24# 0.01fF
C73333 NAND2X1_LOC_21/Y NAND2X1_LOC_587/a_36_24# 0.00fF
C73334 NAND2X1_LOC_59/B NAND2X1_LOC_588/B 0.04fF
C73335 NAND2X1_LOC_784/a_36_24# NAND2X1_LOC_808/A -0.02fF
C73336 NOR2X1_LOC_513/a_36_216# NOR2X1_LOC_152/Y 0.01fF
C73337 NAND2X1_LOC_573/Y NAND2X1_LOC_783/A 0.10fF
C73338 NOR2X1_LOC_824/A D_INPUT_0 0.06fF
C73339 NOR2X1_LOC_405/A INVX1_LOC_87/A 0.03fF
C73340 NOR2X1_LOC_264/Y NOR2X1_LOC_68/A 0.07fF
C73341 NOR2X1_LOC_644/B NOR2X1_LOC_78/B 0.02fF
C73342 NAND2X1_LOC_573/Y NOR2X1_LOC_130/A 0.07fF
C73343 NOR2X1_LOC_667/A NOR2X1_LOC_441/Y 0.09fF
C73344 INVX1_LOC_135/A INVX1_LOC_48/Y 0.01fF
C73345 NAND2X1_LOC_637/Y NOR2X1_LOC_48/Y 0.08fF
C73346 INVX1_LOC_227/A INVX1_LOC_101/Y 0.00fF
C73347 INVX1_LOC_34/A NAND2X1_LOC_731/Y 0.01fF
C73348 INVX1_LOC_17/A NOR2X1_LOC_188/Y 0.01fF
C73349 NAND2X1_LOC_335/a_36_24# INVX1_LOC_30/A 0.00fF
C73350 NOR2X1_LOC_598/B INVX1_LOC_158/Y 0.03fF
C73351 INVX1_LOC_226/Y NOR2X1_LOC_160/B 0.03fF
C73352 NOR2X1_LOC_802/A NAND2X1_LOC_497/a_36_24# 0.01fF
C73353 INVX1_LOC_18/A NOR2X1_LOC_369/a_36_216# 0.02fF
C73354 NAND2X1_LOC_753/a_36_24# NOR2X1_LOC_74/A 0.00fF
C73355 D_INPUT_1 INVX1_LOC_6/A 0.18fF
C73356 NAND2X1_LOC_807/Y NOR2X1_LOC_652/Y 0.07fF
C73357 NAND2X1_LOC_11/Y NAND2X1_LOC_36/A 0.86fF
C73358 NOR2X1_LOC_815/Y NOR2X1_LOC_433/A 0.00fF
C73359 INVX1_LOC_1/A NOR2X1_LOC_123/B 0.10fF
C73360 INVX1_LOC_149/A INVX1_LOC_18/A 0.01fF
C73361 INVX1_LOC_181/Y INVX1_LOC_104/A 0.23fF
C73362 INVX1_LOC_304/A NOR2X1_LOC_438/Y 0.10fF
C73363 INVX1_LOC_21/A INVX1_LOC_182/A 0.07fF
C73364 NOR2X1_LOC_220/A INVX1_LOC_223/A 0.05fF
C73365 NAND2X1_LOC_721/B NOR2X1_LOC_773/Y 0.01fF
C73366 INVX1_LOC_292/A INVX1_LOC_101/A 0.00fF
C73367 NOR2X1_LOC_250/A NAND2X1_LOC_656/Y 0.02fF
C73368 D_INPUT_1 NOR2X1_LOC_10/a_36_216# 0.02fF
C73369 NAND2X1_LOC_254/Y INVX1_LOC_118/A 0.03fF
C73370 NAND2X1_LOC_849/B INVX1_LOC_3/Y 0.28fF
C73371 NOR2X1_LOC_390/a_36_216# NOR2X1_LOC_577/Y 0.01fF
C73372 NAND2X1_LOC_308/Y NOR2X1_LOC_152/Y 0.03fF
C73373 INPUT_4 INVX1_LOC_296/A 0.16fF
C73374 NOR2X1_LOC_35/Y NOR2X1_LOC_541/B 0.50fF
C73375 NOR2X1_LOC_160/B INVX1_LOC_10/A 0.03fF
C73376 NOR2X1_LOC_209/Y INVX1_LOC_24/A 0.07fF
C73377 INVX1_LOC_275/A NAND2X1_LOC_484/a_36_24# 0.00fF
C73378 INVX1_LOC_93/A NOR2X1_LOC_74/A 0.19fF
C73379 INVX1_LOC_84/A INVX1_LOC_63/A 0.13fF
C73380 INVX1_LOC_2/A INVX1_LOC_314/Y 0.10fF
C73381 INVX1_LOC_225/A NOR2X1_LOC_557/Y 0.19fF
C73382 INVX1_LOC_109/Y INVX1_LOC_117/Y 0.00fF
C73383 NOR2X1_LOC_96/Y INVX1_LOC_3/Y 0.03fF
C73384 NOR2X1_LOC_355/A INVX1_LOC_292/A 0.00fF
C73385 NAND2X1_LOC_223/A INVX1_LOC_117/A 0.07fF
C73386 INVX1_LOC_223/A NOR2X1_LOC_548/Y 0.02fF
C73387 INVX1_LOC_43/Y NOR2X1_LOC_71/Y 0.05fF
C73388 NOR2X1_LOC_67/A NAND2X1_LOC_837/Y 0.12fF
C73389 INVX1_LOC_24/A NAND2X1_LOC_852/Y 0.20fF
C73390 INVX1_LOC_6/A NOR2X1_LOC_652/Y 0.09fF
C73391 NOR2X1_LOC_226/A INVX1_LOC_314/Y 0.02fF
C73392 INVX1_LOC_90/A INVX1_LOC_215/Y 0.03fF
C73393 INVX1_LOC_132/A INVX1_LOC_143/A 0.18fF
C73394 VDD INVX1_LOC_112/Y 0.26fF
C73395 NOR2X1_LOC_778/B INVX1_LOC_49/A 0.03fF
C73396 NOR2X1_LOC_270/Y NOR2X1_LOC_665/A 0.04fF
C73397 NAND2X1_LOC_170/A INVX1_LOC_41/Y 0.00fF
C73398 INVX1_LOC_271/Y INVX1_LOC_9/A 0.07fF
C73399 NOR2X1_LOC_435/A INVX1_LOC_15/A 0.01fF
C73400 NAND2X1_LOC_848/Y INVX1_LOC_3/Y -0.02fF
C73401 NAND2X1_LOC_349/B NAND2X1_LOC_515/a_36_24# 0.01fF
C73402 INVX1_LOC_54/Y INVX1_LOC_294/Y 0.05fF
C73403 NOR2X1_LOC_6/B NAND2X1_LOC_141/A 0.06fF
C73404 INVX1_LOC_232/Y INVX1_LOC_34/A 0.00fF
C73405 INVX1_LOC_14/A INVX1_LOC_126/Y 0.08fF
C73406 NOR2X1_LOC_673/B INVX1_LOC_42/A 0.01fF
C73407 NOR2X1_LOC_220/A INVX1_LOC_149/Y 0.02fF
C73408 NOR2X1_LOC_103/Y NOR2X1_LOC_188/A 0.08fF
C73409 NAND2X1_LOC_149/Y NOR2X1_LOC_45/B 0.09fF
C73410 INVX1_LOC_233/A NAND2X1_LOC_633/Y 0.59fF
C73411 NAND2X1_LOC_717/Y NAND2X1_LOC_839/Y 0.01fF
C73412 INVX1_LOC_279/A INVX1_LOC_77/A 0.14fF
C73413 INVX1_LOC_228/A NOR2X1_LOC_332/A 0.03fF
C73414 NOR2X1_LOC_15/Y INVX1_LOC_96/A 0.03fF
C73415 NOR2X1_LOC_220/A INVX1_LOC_85/A 0.03fF
C73416 NOR2X1_LOC_806/Y NOR2X1_LOC_811/B 0.01fF
C73417 INVX1_LOC_58/A NAND2X1_LOC_849/B 0.07fF
C73418 INVX1_LOC_35/A NOR2X1_LOC_706/B 0.00fF
C73419 INVX1_LOC_26/A NAND2X1_LOC_488/a_36_24# 0.00fF
C73420 NAND2X1_LOC_338/B NAND2X1_LOC_360/B 0.10fF
C73421 INVX1_LOC_58/A INVX1_LOC_38/A 2.46fF
C73422 NOR2X1_LOC_201/A NOR2X1_LOC_61/Y 0.00fF
C73423 INVX1_LOC_15/A INVX1_LOC_63/A 0.31fF
C73424 NOR2X1_LOC_401/B INVX1_LOC_164/Y 0.14fF
C73425 NOR2X1_LOC_548/Y INVX1_LOC_149/Y 0.02fF
C73426 NAND2X1_LOC_149/Y INVX1_LOC_199/Y 0.03fF
C73427 INVX1_LOC_292/A NOR2X1_LOC_552/Y 0.00fF
C73428 NAND2X1_LOC_634/Y INVX1_LOC_140/A 0.02fF
C73429 NAND2X1_LOC_99/Y D_INPUT_0 0.00fF
C73430 INVX1_LOC_29/A INVX1_LOC_42/A 0.14fF
C73431 INVX1_LOC_13/A NOR2X1_LOC_720/B 0.03fF
C73432 NOR2X1_LOC_826/a_36_216# INVX1_LOC_280/A 0.00fF
C73433 NOR2X1_LOC_250/a_36_216# INVX1_LOC_91/A 0.01fF
C73434 NAND2X1_LOC_63/Y NOR2X1_LOC_159/a_36_216# 0.00fF
C73435 INVX1_LOC_58/A NOR2X1_LOC_96/Y 0.00fF
C73436 NOR2X1_LOC_52/B NAND2X1_LOC_735/B 0.00fF
C73437 INVX1_LOC_314/Y INPUT_1 0.06fF
C73438 NOR2X1_LOC_500/A NOR2X1_LOC_356/A 1.11fF
C73439 INVX1_LOC_27/A NOR2X1_LOC_266/B 0.01fF
C73440 NOR2X1_LOC_172/a_36_216# INVX1_LOC_53/Y 0.00fF
C73441 INVX1_LOC_45/A NOR2X1_LOC_188/A 0.23fF
C73442 NAND2X1_LOC_796/B VDD 0.01fF
C73443 NOR2X1_LOC_303/Y NOR2X1_LOC_356/A 0.10fF
C73444 NOR2X1_LOC_748/Y NOR2X1_LOC_175/A 0.01fF
C73445 NAND2X1_LOC_392/A NAND2X1_LOC_231/Y 0.01fF
C73446 INVX1_LOC_58/A NOR2X1_LOC_51/A 0.02fF
C73447 NAND2X1_LOC_803/B NAND2X1_LOC_655/A 0.12fF
C73448 NOR2X1_LOC_568/A NOR2X1_LOC_188/A 0.10fF
C73449 NOR2X1_LOC_413/a_36_216# INVX1_LOC_135/A 0.01fF
C73450 INVX1_LOC_11/A NOR2X1_LOC_448/A 0.01fF
C73451 INVX1_LOC_45/A NOR2X1_LOC_548/B 0.03fF
C73452 INVX1_LOC_57/A NOR2X1_LOC_461/A 0.04fF
C73453 NOR2X1_LOC_664/Y D_INPUT_0 0.01fF
C73454 NOR2X1_LOC_568/A NOR2X1_LOC_548/B 0.10fF
C73455 INVX1_LOC_225/A NOR2X1_LOC_130/A 0.03fF
C73456 INVX1_LOC_27/A NOR2X1_LOC_859/Y 0.03fF
C73457 INVX1_LOC_208/A NOR2X1_LOC_500/Y 0.05fF
C73458 INVX1_LOC_58/A NAND2X1_LOC_848/Y 0.01fF
C73459 NOR2X1_LOC_629/a_36_216# INVX1_LOC_135/A 0.01fF
C73460 NOR2X1_LOC_68/A INVX1_LOC_86/A 0.04fF
C73461 INVX1_LOC_248/Y INVX1_LOC_38/A 0.01fF
C73462 NOR2X1_LOC_590/A NAND2X1_LOC_655/A 0.07fF
C73463 INVX1_LOC_63/Y D_GATE_366 0.03fF
C73464 NOR2X1_LOC_604/a_36_216# INVX1_LOC_179/A 0.00fF
C73465 INVX1_LOC_36/A INVX1_LOC_123/A 0.07fF
C73466 INVX1_LOC_182/Y INVX1_LOC_77/A 0.07fF
C73467 NAND2X1_LOC_564/a_36_24# NAND2X1_LOC_551/A 0.00fF
C73468 INVX1_LOC_135/A NOR2X1_LOC_84/Y 0.10fF
C73469 NOR2X1_LOC_391/A NOR2X1_LOC_78/B 0.03fF
C73470 NOR2X1_LOC_554/B INVX1_LOC_201/A 0.02fF
C73471 INVX1_LOC_152/Y INVX1_LOC_152/A 0.28fF
C73472 INVX1_LOC_223/A NAND2X1_LOC_498/a_36_24# 0.00fF
C73473 NAND2X1_LOC_341/A INVX1_LOC_22/A 0.02fF
C73474 NAND2X1_LOC_740/B NOR2X1_LOC_577/Y 0.00fF
C73475 NOR2X1_LOC_32/B INVX1_LOC_260/A 0.05fF
C73476 INVX1_LOC_58/A NOR2X1_LOC_697/a_36_216# 0.00fF
C73477 NOR2X1_LOC_824/A NAND2X1_LOC_848/A 0.03fF
C73478 INVX1_LOC_191/Y NOR2X1_LOC_747/a_36_216# 0.00fF
C73479 INVX1_LOC_48/Y NOR2X1_LOC_813/Y 0.26fF
C73480 NOR2X1_LOC_303/Y NOR2X1_LOC_74/A 0.10fF
C73481 NOR2X1_LOC_174/B NOR2X1_LOC_174/a_36_216# 0.00fF
C73482 INVX1_LOC_64/A NOR2X1_LOC_61/A 0.02fF
C73483 INVX1_LOC_78/A INVX1_LOC_29/A 0.17fF
C73484 NAND2X1_LOC_350/B INVX1_LOC_10/A 0.01fF
C73485 INVX1_LOC_71/A NOR2X1_LOC_188/A 0.44fF
C73486 INVX1_LOC_11/A INVX1_LOC_14/Y 0.07fF
C73487 NAND2X1_LOC_725/A NAND2X1_LOC_802/Y 0.10fF
C73488 INVX1_LOC_134/A NOR2X1_LOC_857/A 0.03fF
C73489 INVX1_LOC_71/A NOR2X1_LOC_548/B 0.03fF
C73490 NAND2X1_LOC_724/A NAND2X1_LOC_811/B 0.12fF
C73491 INVX1_LOC_208/A INVX1_LOC_10/A 0.17fF
C73492 NOR2X1_LOC_79/A NOR2X1_LOC_652/Y 0.00fF
C73493 NAND2X1_LOC_81/B INVX1_LOC_23/Y 0.01fF
C73494 NOR2X1_LOC_15/Y NOR2X1_LOC_684/Y 0.01fF
C73495 NOR2X1_LOC_221/a_36_216# NAND2X1_LOC_425/Y 0.01fF
C73496 INVX1_LOC_279/A NOR2X1_LOC_687/Y 0.11fF
C73497 NAND2X1_LOC_214/B INVX1_LOC_46/Y 0.63fF
C73498 D_INPUT_0 NOR2X1_LOC_251/Y 0.11fF
C73499 INVX1_LOC_14/A NOR2X1_LOC_536/A 0.25fF
C73500 INVX1_LOC_88/A NOR2X1_LOC_366/a_36_216# 0.00fF
C73501 INVX1_LOC_54/Y NOR2X1_LOC_356/A 0.00fF
C73502 NOR2X1_LOC_468/a_36_216# INVX1_LOC_22/A 0.00fF
C73503 INVX1_LOC_98/Y NAND2X1_LOC_842/B 0.04fF
C73504 NOR2X1_LOC_65/B INVX1_LOC_29/A 0.49fF
C73505 NAND2X1_LOC_734/B NOR2X1_LOC_322/Y 0.21fF
C73506 NOR2X1_LOC_191/B NOR2X1_LOC_78/A 0.07fF
C73507 INVX1_LOC_108/Y INVX1_LOC_63/A 1.02fF
C73508 INVX1_LOC_14/A NAND2X1_LOC_659/a_36_24# 0.01fF
C73509 NOR2X1_LOC_68/A NOR2X1_LOC_346/Y 0.01fF
C73510 INVX1_LOC_184/Y INVX1_LOC_186/A 0.25fF
C73511 NOR2X1_LOC_772/B INVX1_LOC_285/A 0.11fF
C73512 INVX1_LOC_278/A INVX1_LOC_63/A 0.01fF
C73513 INVX1_LOC_27/A INVX1_LOC_46/Y 0.21fF
C73514 INVX1_LOC_34/A NOR2X1_LOC_391/Y 0.01fF
C73515 NOR2X1_LOC_376/A NAND2X1_LOC_93/B 0.05fF
C73516 NAND2X1_LOC_740/Y NAND2X1_LOC_770/Y 0.27fF
C73517 INVX1_LOC_24/A NAND2X1_LOC_642/Y 0.05fF
C73518 NOR2X1_LOC_818/a_36_216# INVX1_LOC_63/A 0.00fF
C73519 INVX1_LOC_49/A NOR2X1_LOC_557/A 0.01fF
C73520 INVX1_LOC_14/A NOR2X1_LOC_655/Y 0.15fF
C73521 NOR2X1_LOC_772/B NOR2X1_LOC_814/A 0.20fF
C73522 NOR2X1_LOC_781/A INVX1_LOC_89/A 0.03fF
C73523 NOR2X1_LOC_815/a_36_216# NOR2X1_LOC_45/B 0.00fF
C73524 INVX1_LOC_215/Y INVX1_LOC_38/A 0.04fF
C73525 INVX1_LOC_19/Y NOR2X1_LOC_438/Y 0.24fF
C73526 INVX1_LOC_226/Y NOR2X1_LOC_756/a_36_216# 0.00fF
C73527 D_INPUT_0 INVX1_LOC_234/A 0.14fF
C73528 NOR2X1_LOC_335/a_36_216# INVX1_LOC_150/A 0.02fF
C73529 NOR2X1_LOC_376/A NAND2X1_LOC_425/Y 0.03fF
C73530 NAND2X1_LOC_545/a_36_24# NAND2X1_LOC_211/Y 0.00fF
C73531 NAND2X1_LOC_337/B INVX1_LOC_118/Y 0.02fF
C73532 INVX1_LOC_54/Y NOR2X1_LOC_74/A 0.12fF
C73533 INVX1_LOC_14/A NAND2X1_LOC_93/B 5.41fF
C73534 NOR2X1_LOC_329/B NOR2X1_LOC_321/a_36_216# 0.01fF
C73535 NOR2X1_LOC_445/Y NOR2X1_LOC_318/B 0.34fF
C73536 NOR2X1_LOC_703/B INVX1_LOC_37/A 0.03fF
C73537 INVX1_LOC_269/A INVX1_LOC_92/A 0.07fF
C73538 INVX1_LOC_13/Y NOR2X1_LOC_814/A 0.03fF
C73539 INVX1_LOC_232/Y INPUT_0 0.09fF
C73540 NOR2X1_LOC_793/A NOR2X1_LOC_445/B 0.34fF
C73541 NAND2X1_LOC_354/B NAND2X1_LOC_655/A 0.59fF
C73542 NOR2X1_LOC_557/Y NAND2X1_LOC_642/Y 0.03fF
C73543 NAND2X1_LOC_740/B INVX1_LOC_22/A 0.03fF
C73544 INVX1_LOC_23/Y INVX1_LOC_4/Y 0.10fF
C73545 NOR2X1_LOC_500/B NOR2X1_LOC_862/a_36_216# 0.00fF
C73546 NAND2X1_LOC_528/a_36_24# INVX1_LOC_158/Y 0.00fF
C73547 INVX1_LOC_298/Y INVX1_LOC_78/A 0.01fF
C73548 NOR2X1_LOC_785/Y NOR2X1_LOC_775/Y 0.11fF
C73549 INVX1_LOC_186/A INVX1_LOC_177/A 0.03fF
C73550 INVX1_LOC_96/A INVX1_LOC_96/Y 0.04fF
C73551 INVX1_LOC_19/A NOR2X1_LOC_460/Y 0.37fF
C73552 NAND2X1_LOC_392/A INPUT_0 0.00fF
C73553 INVX1_LOC_230/Y NOR2X1_LOC_88/A 0.01fF
C73554 INVX1_LOC_70/Y INVX1_LOC_168/A 0.53fF
C73555 INVX1_LOC_14/A NOR2X1_LOC_649/B 0.29fF
C73556 INVX1_LOC_89/A NOR2X1_LOC_180/B 0.07fF
C73557 NOR2X1_LOC_160/B INVX1_LOC_307/A 0.39fF
C73558 INVX1_LOC_88/A INVX1_LOC_285/A 0.01fF
C73559 NOR2X1_LOC_335/B INVX1_LOC_1/Y 0.41fF
C73560 NOR2X1_LOC_292/Y INVX1_LOC_22/A 0.21fF
C73561 D_INPUT_6 NOR2X1_LOC_36/B 0.29fF
C73562 INVX1_LOC_14/A INVX1_LOC_3/A 0.28fF
C73563 D_INPUT_0 NOR2X1_LOC_19/B 0.39fF
C73564 NOR2X1_LOC_592/A NOR2X1_LOC_697/Y 0.08fF
C73565 NOR2X1_LOC_522/Y NOR2X1_LOC_536/A 0.01fF
C73566 INVX1_LOC_89/A NOR2X1_LOC_738/A 0.03fF
C73567 INVX1_LOC_50/Y INVX1_LOC_99/A 3.18fF
C73568 INVX1_LOC_88/A NOR2X1_LOC_814/A 0.01fF
C73569 NOR2X1_LOC_160/B NOR2X1_LOC_445/B 0.08fF
C73570 NOR2X1_LOC_291/a_36_216# INVX1_LOC_42/A 0.01fF
C73571 INVX1_LOC_204/A INVX1_LOC_78/A 0.01fF
C73572 NOR2X1_LOC_52/B NAND2X1_LOC_212/Y 0.01fF
C73573 NOR2X1_LOC_180/B NAND2X1_LOC_176/a_36_24# 0.02fF
C73574 INVX1_LOC_41/A NOR2X1_LOC_558/A 0.03fF
C73575 NOR2X1_LOC_357/Y NOR2X1_LOC_364/Y 0.02fF
C73576 INVX1_LOC_276/Y NAND2X1_LOC_655/A 0.05fF
C73577 INVX1_LOC_57/Y INVX1_LOC_185/A 0.16fF
C73578 NAND2X1_LOC_866/B NOR2X1_LOC_497/Y 0.27fF
C73579 NOR2X1_LOC_636/a_36_216# INVX1_LOC_37/A 0.00fF
C73580 NAND2X1_LOC_84/Y NOR2X1_LOC_536/A 0.50fF
C73581 NAND2X1_LOC_139/A VDD 0.21fF
C73582 INVX1_LOC_225/A NOR2X1_LOC_280/Y 0.01fF
C73583 INVX1_LOC_177/A NAND2X1_LOC_447/Y 0.03fF
C73584 NAND2X1_LOC_344/a_36_24# INVX1_LOC_42/A 0.01fF
C73585 NOR2X1_LOC_589/A INVX1_LOC_286/A 0.03fF
C73586 NOR2X1_LOC_209/Y NOR2X1_LOC_209/A 0.08fF
C73587 INVX1_LOC_39/A NAND2X1_LOC_254/Y 0.03fF
C73588 INVX1_LOC_33/A INVX1_LOC_117/A 0.55fF
C73589 NOR2X1_LOC_412/a_36_216# NOR2X1_LOC_813/Y 0.01fF
C73590 NOR2X1_LOC_45/B INVX1_LOC_16/A 0.19fF
C73591 INVX1_LOC_77/A NOR2X1_LOC_450/A 0.04fF
C73592 INVX1_LOC_35/A INVX1_LOC_94/Y 0.03fF
C73593 NOR2X1_LOC_824/A NOR2X1_LOC_754/A -0.02fF
C73594 INVX1_LOC_30/A NOR2X1_LOC_841/A 0.11fF
C73595 INVX1_LOC_89/A NOR2X1_LOC_569/A 0.01fF
C73596 NOR2X1_LOC_742/A INVX1_LOC_311/Y 0.01fF
C73597 NOR2X1_LOC_644/Y VDD 0.23fF
C73598 NOR2X1_LOC_218/Y NOR2X1_LOC_657/B 0.06fF
C73599 INVX1_LOC_52/A NOR2X1_LOC_69/A 0.00fF
C73600 NOR2X1_LOC_749/Y NOR2X1_LOC_548/B 0.07fF
C73601 NAND2X1_LOC_231/Y NAND2X1_LOC_287/B 0.10fF
C73602 INVX1_LOC_72/A NAND2X1_LOC_572/B 0.12fF
C73603 NOR2X1_LOC_413/a_36_216# INVX1_LOC_280/A 0.00fF
C73604 INVX1_LOC_63/Y NOR2X1_LOC_142/a_36_216# 0.01fF
C73605 NAND2X1_LOC_9/Y NOR2X1_LOC_39/a_36_216# 0.00fF
C73606 INVX1_LOC_171/A INVX1_LOC_286/A 0.50fF
C73607 INVX1_LOC_144/Y NAND2X1_LOC_453/A -0.02fF
C73608 INVX1_LOC_16/A INVX1_LOC_247/A 0.00fF
C73609 NAND2X1_LOC_190/Y INVX1_LOC_290/Y 0.01fF
C73610 D_INPUT_1 INVX1_LOC_270/A 0.11fF
C73611 NOR2X1_LOC_589/A INVX1_LOC_95/A 0.00fF
C73612 NOR2X1_LOC_500/B NOR2X1_LOC_814/A 0.10fF
C73613 NOR2X1_LOC_813/Y NOR2X1_LOC_84/Y 0.17fF
C73614 INVX1_LOC_41/A NOR2X1_LOC_729/A 0.00fF
C73615 NAND2X1_LOC_541/Y VDD 0.01fF
C73616 NAND2X1_LOC_550/A INVX1_LOC_12/A 0.03fF
C73617 INVX1_LOC_53/A NAND2X1_LOC_64/a_36_24# -0.00fF
C73618 NOR2X1_LOC_835/A INVX1_LOC_143/Y 0.02fF
C73619 INVX1_LOC_35/A INVX1_LOC_181/A 0.07fF
C73620 NOR2X1_LOC_629/a_36_216# INVX1_LOC_280/A 0.00fF
C73621 D_INPUT_1 NOR2X1_LOC_416/A 0.01fF
C73622 NOR2X1_LOC_160/B INVX1_LOC_12/A 0.17fF
C73623 NOR2X1_LOC_433/a_36_216# INVX1_LOC_54/A 0.00fF
C73624 INVX1_LOC_268/A INVX1_LOC_76/A 0.05fF
C73625 NAND2X1_LOC_140/a_36_24# NOR2X1_LOC_155/A 0.01fF
C73626 NAND2X1_LOC_112/Y NOR2X1_LOC_136/a_36_216# 0.00fF
C73627 NOR2X1_LOC_84/Y INVX1_LOC_280/A 0.09fF
C73628 NOR2X1_LOC_382/Y INVX1_LOC_19/A 0.03fF
C73629 NOR2X1_LOC_130/A NAND2X1_LOC_642/Y 0.03fF
C73630 INVX1_LOC_132/A NOR2X1_LOC_197/B 0.01fF
C73631 NOR2X1_LOC_844/Y INVX1_LOC_29/A 0.02fF
C73632 NAND2X1_LOC_88/a_36_24# INVX1_LOC_230/A 0.00fF
C73633 INVX1_LOC_23/A NOR2X1_LOC_678/A 0.04fF
C73634 NOR2X1_LOC_770/Y INVX1_LOC_91/A 0.01fF
C73635 NOR2X1_LOC_68/A NOR2X1_LOC_662/A 0.03fF
C73636 NAND2X1_LOC_112/Y VDD 0.54fF
C73637 INVX1_LOC_40/A INVX1_LOC_117/A 0.12fF
C73638 NOR2X1_LOC_97/A INPUT_0 0.05fF
C73639 INVX1_LOC_180/A NOR2X1_LOC_435/B 0.27fF
C73640 INVX1_LOC_30/A INPUT_7 0.02fF
C73641 INVX1_LOC_28/A NOR2X1_LOC_45/B 0.40fF
C73642 NOR2X1_LOC_817/Y INVX1_LOC_4/A 0.19fF
C73643 NOR2X1_LOC_664/Y INVX1_LOC_46/Y 0.00fF
C73644 NOR2X1_LOC_121/Y NOR2X1_LOC_216/B 0.13fF
C73645 NOR2X1_LOC_769/A INVX1_LOC_29/A 0.01fF
C73646 INVX1_LOC_270/A NOR2X1_LOC_108/a_36_216# 0.01fF
C73647 NOR2X1_LOC_373/Y INVX1_LOC_20/A 0.07fF
C73648 INVX1_LOC_10/A NAND2X1_LOC_211/Y 3.80fF
C73649 NOR2X1_LOC_666/Y NAND2X1_LOC_454/Y 0.09fF
C73650 INVX1_LOC_1/A NAND2X1_LOC_467/a_36_24# 0.00fF
C73651 INVX1_LOC_16/A INVX1_LOC_281/A 0.07fF
C73652 NOR2X1_LOC_554/B INVX1_LOC_29/A 0.03fF
C73653 INVX1_LOC_303/A NOR2X1_LOC_814/A 0.07fF
C73654 NAND2X1_LOC_195/Y INVX1_LOC_12/A 0.01fF
C73655 NAND2X1_LOC_326/a_36_24# NOR2X1_LOC_88/Y 0.01fF
C73656 NOR2X1_LOC_612/B NAND2X1_LOC_93/B 0.07fF
C73657 NOR2X1_LOC_355/B INVX1_LOC_75/A 0.06fF
C73658 NOR2X1_LOC_716/B INVX1_LOC_119/Y 0.07fF
C73659 NOR2X1_LOC_772/B NOR2X1_LOC_292/a_36_216# 0.00fF
C73660 NOR2X1_LOC_355/A NOR2X1_LOC_137/Y 0.01fF
C73661 NOR2X1_LOC_733/a_36_216# INVX1_LOC_12/A 0.00fF
C73662 INVX1_LOC_174/A NAND2X1_LOC_3/B 0.35fF
C73663 INVX1_LOC_217/Y NOR2X1_LOC_649/B 0.05fF
C73664 NOR2X1_LOC_772/Y NAND2X1_LOC_475/Y 0.10fF
C73665 NAND2X1_LOC_860/A INVX1_LOC_306/Y 0.59fF
C73666 NAND2X1_LOC_634/Y INVX1_LOC_42/A 0.17fF
C73667 INVX1_LOC_314/Y NAND2X1_LOC_63/Y 0.56fF
C73668 NOR2X1_LOC_318/B NOR2X1_LOC_335/B 0.49fF
C73669 NOR2X1_LOC_721/Y NOR2X1_LOC_78/A 0.44fF
C73670 D_INPUT_7 NAND2X1_LOC_430/B 0.00fF
C73671 INVX1_LOC_22/A NOR2X1_LOC_641/Y 0.02fF
C73672 NOR2X1_LOC_152/Y INVX1_LOC_29/A 0.07fF
C73673 INVX1_LOC_234/A NAND2X1_LOC_848/A 0.09fF
C73674 NAND2X1_LOC_569/A NAND2X1_LOC_768/Y 0.29fF
C73675 NAND2X1_LOC_170/A INVX1_LOC_185/A 1.03fF
C73676 INVX1_LOC_228/A NOR2X1_LOC_847/A 0.09fF
C73677 NAND2X1_LOC_793/Y INVX1_LOC_26/A 0.15fF
C73678 INVX1_LOC_279/A INVX1_LOC_9/A 0.07fF
C73679 NOR2X1_LOC_596/A INVX1_LOC_290/Y 0.07fF
C73680 NOR2X1_LOC_589/A INVX1_LOC_54/A 0.66fF
C73681 INVX1_LOC_208/A INVX1_LOC_307/A 0.04fF
C73682 INVX1_LOC_30/A INVX1_LOC_128/A 0.01fF
C73683 NOR2X1_LOC_516/B INVX1_LOC_307/A 0.12fF
C73684 NOR2X1_LOC_516/B NOR2X1_LOC_445/B 0.10fF
C73685 INVX1_LOC_269/A INVX1_LOC_53/A 0.11fF
C73686 NAND2X1_LOC_840/Y VDD 0.00fF
C73687 INVX1_LOC_310/A NOR2X1_LOC_691/B 0.28fF
C73688 INVX1_LOC_136/A NOR2X1_LOC_409/B 0.00fF
C73689 INVX1_LOC_35/A INVX1_LOC_299/A 0.22fF
C73690 NAND2X1_LOC_634/Y INVX1_LOC_78/A 0.03fF
C73691 NAND2X1_LOC_339/a_36_24# INVX1_LOC_109/A 0.00fF
C73692 NOR2X1_LOC_703/B NAND2X1_LOC_72/B 0.00fF
C73693 INVX1_LOC_186/A INVX1_LOC_65/A 0.12fF
C73694 INPUT_0 NAND2X1_LOC_287/B 0.07fF
C73695 INVX1_LOC_43/Y NAND2X1_LOC_205/A 0.02fF
C73696 INVX1_LOC_35/A NOR2X1_LOC_538/B 0.00fF
C73697 INVX1_LOC_8/A INVX1_LOC_42/A 0.27fF
C73698 INVX1_LOC_286/A INVX1_LOC_20/A 0.49fF
C73699 NOR2X1_LOC_75/Y NOR2X1_LOC_604/Y 0.01fF
C73700 NAND2X1_LOC_842/B NOR2X1_LOC_709/B 0.44fF
C73701 INVX1_LOC_33/A INVX1_LOC_3/Y 0.07fF
C73702 NOR2X1_LOC_631/B INVX1_LOC_91/A 0.46fF
C73703 INVX1_LOC_1/Y INVX1_LOC_84/A 0.25fF
C73704 INPUT_0 INVX1_LOC_129/Y 0.02fF
C73705 NOR2X1_LOC_6/B NOR2X1_LOC_128/a_36_216# 0.01fF
C73706 NOR2X1_LOC_728/B INVX1_LOC_37/A 0.03fF
C73707 D_INPUT_0 NOR2X1_LOC_216/B 0.03fF
C73708 NOR2X1_LOC_45/B NOR2X1_LOC_253/Y 0.05fF
C73709 NAND2X1_LOC_778/Y NOR2X1_LOC_15/Y 0.03fF
C73710 NOR2X1_LOC_647/A NOR2X1_LOC_820/A 0.01fF
C73711 INVX1_LOC_182/Y INVX1_LOC_9/A -0.01fF
C73712 NOR2X1_LOC_455/Y INVX1_LOC_188/A 0.01fF
C73713 NAND2X1_LOC_35/Y NOR2X1_LOC_615/a_36_216# 0.01fF
C73714 INVX1_LOC_279/Y NOR2X1_LOC_598/B 0.01fF
C73715 INVX1_LOC_72/A NOR2X1_LOC_654/A 0.03fF
C73716 INVX1_LOC_166/A NOR2X1_LOC_476/Y 0.04fF
C73717 INVX1_LOC_243/Y NOR2X1_LOC_68/A 0.01fF
C73718 INVX1_LOC_98/A VDD 0.62fF
C73719 D_INPUT_1 INVX1_LOC_36/A 1.00fF
C73720 NOR2X1_LOC_757/Y NOR2X1_LOC_755/Y 0.02fF
C73721 NOR2X1_LOC_272/Y INVX1_LOC_103/A 0.00fF
C73722 NOR2X1_LOC_78/A VDD 1.81fF
C73723 NAND2X1_LOC_785/B NAND2X1_LOC_787/A 0.01fF
C73724 INVX1_LOC_37/A INVX1_LOC_91/A 0.22fF
C73725 INVX1_LOC_95/A INVX1_LOC_20/A 0.01fF
C73726 INVX1_LOC_226/Y NAND2X1_LOC_207/B 0.12fF
C73727 INVX1_LOC_208/A INVX1_LOC_12/A 0.07fF
C73728 NOR2X1_LOC_833/Y NOR2X1_LOC_840/a_36_216# -0.02fF
C73729 NAND2X1_LOC_112/Y INVX1_LOC_133/A 0.00fF
C73730 NOR2X1_LOC_68/A INVX1_LOC_57/A 0.33fF
C73731 NOR2X1_LOC_510/a_36_216# NOR2X1_LOC_697/Y 0.00fF
C73732 INVX1_LOC_247/A NOR2X1_LOC_35/Y 0.03fF
C73733 INVX1_LOC_298/Y INVX1_LOC_113/Y 0.06fF
C73734 NOR2X1_LOC_24/a_36_216# NOR2X1_LOC_24/Y 0.03fF
C73735 INVX1_LOC_48/A NOR2X1_LOC_536/A 0.49fF
C73736 NOR2X1_LOC_19/B INVX1_LOC_46/Y 0.27fF
C73737 D_INPUT_0 NAND2X1_LOC_477/Y 0.07fF
C73738 NOR2X1_LOC_220/A INVX1_LOC_290/Y 0.01fF
C73739 NOR2X1_LOC_516/B INVX1_LOC_12/A 0.03fF
C73740 NOR2X1_LOC_112/Y NOR2X1_LOC_865/Y 0.01fF
C73741 INVX1_LOC_8/A INVX1_LOC_78/A 0.06fF
C73742 NAND2X1_LOC_241/Y NAND2X1_LOC_244/A 0.28fF
C73743 NOR2X1_LOC_590/A INVX1_LOC_13/Y 0.08fF
C73744 NOR2X1_LOC_112/Y NOR2X1_LOC_243/B 0.01fF
C73745 NOR2X1_LOC_326/Y NOR2X1_LOC_854/a_36_216# 0.00fF
C73746 NOR2X1_LOC_607/Y INVX1_LOC_270/A 0.06fF
C73747 D_INPUT_3 INVX1_LOC_74/A 0.00fF
C73748 NOR2X1_LOC_34/A NOR2X1_LOC_160/B 0.02fF
C73749 NOR2X1_LOC_589/A NAND2X1_LOC_807/B 0.06fF
C73750 NOR2X1_LOC_186/Y INVX1_LOC_286/Y 0.13fF
C73751 NOR2X1_LOC_389/B NAND2X1_LOC_475/Y 0.00fF
C73752 INVX1_LOC_304/A NOR2X1_LOC_176/Y 0.02fF
C73753 NOR2X1_LOC_545/A INVX1_LOC_57/A 0.03fF
C73754 INVX1_LOC_40/A INVX1_LOC_3/Y 2.61fF
C73755 INVX1_LOC_204/A INVX1_LOC_113/Y 0.01fF
C73756 INVX1_LOC_93/Y NOR2X1_LOC_440/a_36_216# 0.00fF
C73757 NOR2X1_LOC_763/Y NAND2X1_LOC_639/a_36_24# 0.01fF
C73758 NOR2X1_LOC_486/Y INVX1_LOC_117/A 0.09fF
C73759 INVX1_LOC_49/A INVX1_LOC_271/A 0.03fF
C73760 NOR2X1_LOC_454/Y NOR2X1_LOC_389/A 0.10fF
C73761 INVX1_LOC_36/A NOR2X1_LOC_652/Y 0.19fF
C73762 NOR2X1_LOC_65/B INVX1_LOC_8/A 0.07fF
C73763 NAND2X1_LOC_803/B INVX1_LOC_88/A 0.02fF
C73764 NOR2X1_LOC_335/A INVX1_LOC_23/A 0.03fF
C73765 NAND2X1_LOC_861/Y INVX1_LOC_29/A 0.03fF
C73766 NOR2X1_LOC_647/B INVX1_LOC_14/A 0.02fF
C73767 NAND2X1_LOC_721/A NOR2X1_LOC_825/Y 0.04fF
C73768 NAND2X1_LOC_573/Y INVX1_LOC_286/Y 0.10fF
C73769 INVX1_LOC_58/A INVX1_LOC_33/A 8.31fF
C73770 NOR2X1_LOC_454/Y NAND2X1_LOC_199/B 0.06fF
C73771 NOR2X1_LOC_742/A INVX1_LOC_84/A 0.07fF
C73772 INVX1_LOC_71/A NOR2X1_LOC_129/a_36_216# 0.12fF
C73773 NOR2X1_LOC_72/a_36_216# NAND2X1_LOC_74/B 0.00fF
C73774 NOR2X1_LOC_822/Y NOR2X1_LOC_821/a_36_216# 0.00fF
C73775 NOR2X1_LOC_741/A INVX1_LOC_92/A 0.02fF
C73776 NAND2X1_LOC_642/Y NOR2X1_LOC_16/a_36_216# 0.00fF
C73777 INVX1_LOC_20/Y NAND2X1_LOC_207/Y 0.11fF
C73778 NOR2X1_LOC_590/A INVX1_LOC_88/A 0.01fF
C73779 INVX1_LOC_5/A NAND2X1_LOC_79/Y 0.01fF
C73780 INVX1_LOC_232/A INVX1_LOC_4/Y 0.19fF
C73781 NAND2X1_LOC_840/B INVX1_LOC_273/A 0.01fF
C73782 INVX1_LOC_45/A NAND2X1_LOC_326/A 0.48fF
C73783 VDD NOR2X1_LOC_60/Y 0.03fF
C73784 NOR2X1_LOC_99/B NOR2X1_LOC_865/a_36_216# 0.01fF
C73785 NOR2X1_LOC_186/Y NOR2X1_LOC_191/B 0.10fF
C73786 D_INPUT_1 NOR2X1_LOC_309/Y 0.03fF
C73787 NOR2X1_LOC_614/a_36_216# INVX1_LOC_33/A 0.00fF
C73788 NAND2X1_LOC_158/a_36_24# INVX1_LOC_78/A 0.00fF
C73789 INVX1_LOC_147/Y INVX1_LOC_54/A 0.13fF
C73790 NOR2X1_LOC_454/Y INVX1_LOC_107/A 0.04fF
C73791 NAND2X1_LOC_134/a_36_24# INVX1_LOC_57/A 0.00fF
C73792 INVX1_LOC_64/A NOR2X1_LOC_570/B 0.02fF
C73793 NOR2X1_LOC_420/Y INVX1_LOC_77/A 0.05fF
C73794 INVX1_LOC_48/A INVX1_LOC_3/A 0.52fF
C73795 NOR2X1_LOC_43/Y NOR2X1_LOC_592/B 0.01fF
C73796 INVX1_LOC_2/A INVX1_LOC_271/A 0.28fF
C73797 INVX1_LOC_20/A INVX1_LOC_54/A 1.40fF
C73798 NOR2X1_LOC_826/Y NOR2X1_LOC_52/B 0.05fF
C73799 INVX1_LOC_269/A NAND2X1_LOC_166/a_36_24# 0.00fF
C73800 NOR2X1_LOC_92/Y INVX1_LOC_181/Y 0.07fF
C73801 INVX1_LOC_295/A NOR2X1_LOC_467/A 0.38fF
C73802 NOR2X1_LOC_454/Y NOR2X1_LOC_596/A 0.07fF
C73803 NOR2X1_LOC_226/A INVX1_LOC_271/A 0.65fF
C73804 NAND2X1_LOC_656/Y NOR2X1_LOC_334/Y 0.34fF
C73805 INVX1_LOC_35/A NOR2X1_LOC_315/Y 0.03fF
C73806 NOR2X1_LOC_709/A NOR2X1_LOC_717/A 0.46fF
C73807 INVX1_LOC_27/A INVX1_LOC_49/A 0.15fF
C73808 INVX1_LOC_158/Y INVX1_LOC_29/A 0.03fF
C73809 NOR2X1_LOC_191/A INVX1_LOC_23/A 0.01fF
C73810 NOR2X1_LOC_318/B INVX1_LOC_84/A 0.07fF
C73811 NOR2X1_LOC_389/A NAND2X1_LOC_387/a_36_24# 0.02fF
C73812 NOR2X1_LOC_272/Y INVX1_LOC_67/A 0.01fF
C73813 NOR2X1_LOC_75/Y INVX1_LOC_72/A 0.01fF
C73814 NAND2X1_LOC_740/a_36_24# INVX1_LOC_72/A 0.07fF
C73815 NAND2X1_LOC_550/A INVX1_LOC_217/A 0.10fF
C73816 NOR2X1_LOC_218/Y INVX1_LOC_271/A 0.02fF
C73817 NOR2X1_LOC_590/A NOR2X1_LOC_500/B 0.48fF
C73818 INVX1_LOC_58/A NAND2X1_LOC_726/Y 0.07fF
C73819 NOR2X1_LOC_98/B INVX1_LOC_9/A 0.03fF
C73820 INVX1_LOC_93/Y INVX1_LOC_84/A 0.07fF
C73821 NOR2X1_LOC_13/Y NAND2X1_LOC_538/Y 0.02fF
C73822 NOR2X1_LOC_309/Y NOR2X1_LOC_652/Y 0.14fF
C73823 INVX1_LOC_22/Y NOR2X1_LOC_500/B 0.03fF
C73824 NOR2X1_LOC_216/B NOR2X1_LOC_266/B 0.01fF
C73825 INVX1_LOC_230/Y INVX1_LOC_18/A 0.03fF
C73826 NAND2X1_LOC_199/B NAND2X1_LOC_196/a_36_24# 0.02fF
C73827 INVX1_LOC_277/A INVX1_LOC_45/A 0.20fF
C73828 NOR2X1_LOC_689/Y NAND2X1_LOC_731/a_36_24# 0.00fF
C73829 INVX1_LOC_58/A NOR2X1_LOC_605/B 0.01fF
C73830 INVX1_LOC_254/A INVX1_LOC_224/A 0.02fF
C73831 NOR2X1_LOC_742/A INVX1_LOC_15/A 0.03fF
C73832 NOR2X1_LOC_13/Y NOR2X1_LOC_250/A 0.04fF
C73833 INVX1_LOC_2/A NAND2X1_LOC_214/B 0.03fF
C73834 NOR2X1_LOC_67/A NAND2X1_LOC_35/Y 0.02fF
C73835 NOR2X1_LOC_45/Y INVX1_LOC_159/A 0.07fF
C73836 NOR2X1_LOC_533/Y NOR2X1_LOC_753/a_36_216# 0.00fF
C73837 NOR2X1_LOC_557/A NAND2X1_LOC_63/Y 0.08fF
C73838 INVX1_LOC_245/A NOR2X1_LOC_598/B 0.03fF
C73839 NOR2X1_LOC_545/a_36_216# INVX1_LOC_57/A 0.00fF
C73840 INVX1_LOC_71/A NAND2X1_LOC_807/A 0.07fF
C73841 NAND2X1_LOC_721/A NOR2X1_LOC_88/Y 0.21fF
C73842 NOR2X1_LOC_45/B INVX1_LOC_109/A 0.04fF
C73843 NAND2X1_LOC_654/B NOR2X1_LOC_158/Y 0.02fF
C73844 NOR2X1_LOC_349/A NOR2X1_LOC_340/A 0.07fF
C73845 NOR2X1_LOC_590/A NOR2X1_LOC_758/a_36_216# 0.00fF
C73846 INVX1_LOC_2/A INVX1_LOC_27/A 0.24fF
C73847 INVX1_LOC_2/A NOR2X1_LOC_824/A 0.07fF
C73848 INVX1_LOC_16/A NOR2X1_LOC_53/Y 0.06fF
C73849 NOR2X1_LOC_489/a_36_216# INVX1_LOC_1/Y 0.00fF
C73850 NAND2X1_LOC_9/Y NOR2X1_LOC_391/A 0.03fF
C73851 NAND2X1_LOC_550/A NAND2X1_LOC_787/B 0.05fF
C73852 INVX1_LOC_101/Y INVX1_LOC_104/A 0.02fF
C73853 INVX1_LOC_64/A INVX1_LOC_215/A 0.02fF
C73854 NOR2X1_LOC_226/A INVX1_LOC_27/A 0.10fF
C73855 INVX1_LOC_25/A INVX1_LOC_135/A 0.30fF
C73856 INVX1_LOC_230/Y INVX1_LOC_172/A 0.00fF
C73857 INVX1_LOC_255/Y NOR2X1_LOC_662/a_36_216# 0.01fF
C73858 INVX1_LOC_269/A INVX1_LOC_80/Y 0.02fF
C73859 NOR2X1_LOC_389/A INVX1_LOC_77/A 0.10fF
C73860 INVX1_LOC_303/A NOR2X1_LOC_590/A 0.07fF
C73861 NOR2X1_LOC_719/B NOR2X1_LOC_392/Y 0.05fF
C73862 INVX1_LOC_81/A INVX1_LOC_81/Y 0.16fF
C73863 NAND2X1_LOC_721/A INVX1_LOC_84/A 0.09fF
C73864 INVX1_LOC_5/A NOR2X1_LOC_748/Y 0.03fF
C73865 INVX1_LOC_303/A INVX1_LOC_22/Y 0.02fF
C73866 NOR2X1_LOC_388/Y NOR2X1_LOC_794/B 0.00fF
C73867 INVX1_LOC_286/A INVX1_LOC_4/A 0.14fF
C73868 INVX1_LOC_36/A NOR2X1_LOC_403/B 0.26fF
C73869 NOR2X1_LOC_429/a_36_216# INVX1_LOC_30/A 0.01fF
C73870 INVX1_LOC_35/A INVX1_LOC_66/A 0.01fF
C73871 NOR2X1_LOC_510/Y NAND2X1_LOC_112/Y 0.02fF
C73872 INVX1_LOC_228/A NOR2X1_LOC_554/B 0.17fF
C73873 NOR2X1_LOC_760/a_36_216# INVX1_LOC_104/A 0.00fF
C73874 INVX1_LOC_248/A NAND2X1_LOC_579/A 0.02fF
C73875 INVX1_LOC_24/A NOR2X1_LOC_91/Y 0.03fF
C73876 INVX1_LOC_269/A NOR2X1_LOC_78/B 0.18fF
C73877 NOR2X1_LOC_598/B NOR2X1_LOC_788/B 0.01fF
C73878 INVX1_LOC_25/A NOR2X1_LOC_248/a_36_216# 0.00fF
C73879 NAND2X1_LOC_787/A INVX1_LOC_90/A 0.04fF
C73880 NAND2X1_LOC_848/A NAND2X1_LOC_477/Y 0.62fF
C73881 NOR2X1_LOC_172/Y INVX1_LOC_30/A 0.08fF
C73882 NAND2X1_LOC_363/B INVX1_LOC_90/A 0.07fF
C73883 INVX1_LOC_299/A INVX1_LOC_305/Y 0.00fF
C73884 NOR2X1_LOC_772/Y INVX1_LOC_30/A 0.09fF
C73885 NAND2X1_LOC_360/B NOR2X1_LOC_103/Y 0.16fF
C73886 INVX1_LOC_256/A INVX1_LOC_111/Y 0.02fF
C73887 NOR2X1_LOC_716/B INVX1_LOC_72/A 0.10fF
C73888 INVX1_LOC_225/A INVX1_LOC_286/Y 0.01fF
C73889 NOR2X1_LOC_48/B INVX1_LOC_20/A 8.41fF
C73890 NOR2X1_LOC_147/B INVX1_LOC_30/A 0.01fF
C73891 INPUT_0 NOR2X1_LOC_72/Y -0.00fF
C73892 INVX1_LOC_62/Y INVX1_LOC_77/A 0.46fF
C73893 NAND2X1_LOC_273/a_36_24# NOR2X1_LOC_743/Y 0.00fF
C73894 D_INPUT_0 INVX1_LOC_93/A 0.07fF
C73895 INVX1_LOC_91/A NAND2X1_LOC_72/B 0.14fF
C73896 NOR2X1_LOC_392/B INVX1_LOC_30/A 0.10fF
C73897 INVX1_LOC_1/A NAND2X1_LOC_479/Y 0.07fF
C73898 NOR2X1_LOC_186/Y NAND2X1_LOC_803/a_36_24# 0.00fF
C73899 NOR2X1_LOC_643/A NOR2X1_LOC_516/B 0.00fF
C73900 INVX1_LOC_58/A NOR2X1_LOC_323/Y 0.01fF
C73901 NOR2X1_LOC_596/A INVX1_LOC_77/A 0.05fF
C73902 NOR2X1_LOC_366/a_36_216# INVX1_LOC_272/A 0.01fF
C73903 NAND2X1_LOC_579/A NOR2X1_LOC_521/Y 0.02fF
C73904 NOR2X1_LOC_628/a_36_216# NAND2X1_LOC_735/B 0.00fF
C73905 INVX1_LOC_5/A D_GATE_366 4.39fF
C73906 INVX1_LOC_106/Y INVX1_LOC_117/A 0.03fF
C73907 NAND2X1_LOC_214/B INPUT_1 0.03fF
C73908 NOR2X1_LOC_361/B NAND2X1_LOC_112/Y 0.04fF
C73909 INVX1_LOC_228/Y NOR2X1_LOC_516/B 0.01fF
C73910 NOR2X1_LOC_433/A NOR2X1_LOC_106/Y 0.15fF
C73911 INVX1_LOC_102/Y NOR2X1_LOC_129/a_36_216# 0.00fF
C73912 INVX1_LOC_249/A INVX1_LOC_49/A 0.03fF
C73913 NAND2X1_LOC_447/Y INVX1_LOC_4/Y 0.12fF
C73914 NOR2X1_LOC_440/Y INVX1_LOC_14/A 0.07fF
C73915 INVX1_LOC_90/A NOR2X1_LOC_791/Y 0.01fF
C73916 NAND2X1_LOC_785/B NAND2X1_LOC_722/A 0.28fF
C73917 INVX1_LOC_41/A INVX1_LOC_181/Y 0.01fF
C73918 INVX1_LOC_25/A NOR2X1_LOC_391/B 0.03fF
C73919 NAND2X1_LOC_715/B NOR2X1_LOC_135/Y 0.05fF
C73920 INVX1_LOC_27/A INPUT_1 0.19fF
C73921 INVX1_LOC_293/A NOR2X1_LOC_121/A 0.00fF
C73922 INVX1_LOC_227/A INVX1_LOC_88/A 0.10fF
C73923 NOR2X1_LOC_824/A INPUT_1 0.69fF
C73924 NOR2X1_LOC_415/A INVX1_LOC_14/A 0.04fF
C73925 INVX1_LOC_135/A INVX1_LOC_1/A 0.29fF
C73926 NAND2X1_LOC_860/A NOR2X1_LOC_9/Y 0.01fF
C73927 NOR2X1_LOC_126/a_36_216# INVX1_LOC_46/Y 0.01fF
C73928 INVX1_LOC_269/A INVX1_LOC_83/A 0.46fF
C73929 INVX1_LOC_225/A NOR2X1_LOC_191/B 0.03fF
C73930 NOR2X1_LOC_441/Y NOR2X1_LOC_131/Y 0.03fF
C73931 NOR2X1_LOC_361/B NAND2X1_LOC_474/a_36_24# 0.00fF
C73932 NOR2X1_LOC_598/B NOR2X1_LOC_147/A 0.03fF
C73933 NOR2X1_LOC_726/Y NOR2X1_LOC_731/Y 0.01fF
C73934 NOR2X1_LOC_523/A NOR2X1_LOC_99/B -0.02fF
C73935 INVX1_LOC_295/A INVX1_LOC_1/A 0.14fF
C73936 NAND2X1_LOC_850/A NAND2X1_LOC_474/Y 0.10fF
C73937 INVX1_LOC_163/A INVX1_LOC_175/Y 0.01fF
C73938 INVX1_LOC_6/A NOR2X1_LOC_678/A 0.03fF
C73939 NOR2X1_LOC_295/Y INVX1_LOC_77/A 0.04fF
C73940 NOR2X1_LOC_300/Y INVX1_LOC_71/A 0.01fF
C73941 INVX1_LOC_255/Y NOR2X1_LOC_514/A 0.05fF
C73942 INVX1_LOC_77/A NOR2X1_LOC_844/A 0.02fF
C73943 NOR2X1_LOC_441/Y NOR2X1_LOC_589/A 3.02fF
C73944 NAND2X1_LOC_384/a_36_24# INVX1_LOC_43/Y 0.01fF
C73945 INVX1_LOC_20/A NOR2X1_LOC_438/Y 0.04fF
C73946 INVX1_LOC_170/Y INVX1_LOC_118/A 0.01fF
C73947 NOR2X1_LOC_134/Y INVX1_LOC_234/A 0.00fF
C73948 INPUT_0 INVX1_LOC_50/Y 0.08fF
C73949 INVX1_LOC_249/A INVX1_LOC_2/A 0.09fF
C73950 NOR2X1_LOC_712/Y NOR2X1_LOC_732/A 0.05fF
C73951 NAND2X1_LOC_360/B INVX1_LOC_71/A 0.12fF
C73952 INVX1_LOC_90/A NOR2X1_LOC_457/A 0.17fF
C73953 INVX1_LOC_34/A NOR2X1_LOC_6/B 0.16fF
C73954 NOR2X1_LOC_419/Y NOR2X1_LOC_537/Y 0.07fF
C73955 NOR2X1_LOC_270/Y INVX1_LOC_16/A 0.41fF
C73956 NOR2X1_LOC_38/B INVX1_LOC_9/A 0.03fF
C73957 NOR2X1_LOC_419/Y NAND2X1_LOC_338/B 0.10fF
C73958 NOR2X1_LOC_690/A NOR2X1_LOC_52/B 0.14fF
C73959 NOR2X1_LOC_537/A NOR2X1_LOC_537/Y 0.00fF
C73960 INVX1_LOC_278/A INVX1_LOC_93/Y 0.02fF
C73961 INVX1_LOC_20/A NAND2X1_LOC_215/A 0.07fF
C73962 NAND2X1_LOC_73/a_36_24# NAND2X1_LOC_74/B 0.03fF
C73963 NOR2X1_LOC_413/Y NOR2X1_LOC_52/B 0.01fF
C73964 NOR2X1_LOC_716/B NOR2X1_LOC_537/Y 0.07fF
C73965 NOR2X1_LOC_220/A INVX1_LOC_77/A 0.01fF
C73966 NOR2X1_LOC_644/Y INVX1_LOC_153/Y 0.01fF
C73967 NOR2X1_LOC_295/Y INVX1_LOC_124/A 0.04fF
C73968 NAND2X1_LOC_795/a_36_24# INVX1_LOC_34/A 0.01fF
C73969 NAND2X1_LOC_647/B NOR2X1_LOC_612/Y 0.00fF
C73970 INVX1_LOC_299/A NOR2X1_LOC_534/a_36_216# 0.00fF
C73971 NOR2X1_LOC_489/a_36_216# INVX1_LOC_93/Y 0.01fF
C73972 INVX1_LOC_78/A INVX1_LOC_118/Y 0.03fF
C73973 INVX1_LOC_117/Y INVX1_LOC_15/A 0.03fF
C73974 NOR2X1_LOC_381/Y INPUT_0 0.03fF
C73975 NAND2X1_LOC_303/Y INVX1_LOC_140/Y 0.08fF
C73976 NOR2X1_LOC_251/Y INVX1_LOC_49/A 0.00fF
C73977 INVX1_LOC_117/A NOR2X1_LOC_635/B 0.02fF
C73978 INVX1_LOC_135/A NOR2X1_LOC_384/Y 0.31fF
C73979 NOR2X1_LOC_664/Y NOR2X1_LOC_818/Y 0.00fF
C73980 INVX1_LOC_232/Y NOR2X1_LOC_514/a_36_216# 0.00fF
C73981 NOR2X1_LOC_510/Y NOR2X1_LOC_78/A 0.00fF
C73982 NOR2X1_LOC_262/Y INVX1_LOC_1/Y 0.01fF
C73983 NOR2X1_LOC_178/Y INVX1_LOC_95/Y 0.18fF
C73984 INVX1_LOC_255/Y NOR2X1_LOC_617/Y 0.04fF
C73985 INVX1_LOC_1/A NOR2X1_LOC_711/A 1.01fF
C73986 NAND2X1_LOC_705/a_36_24# NAND2X1_LOC_787/B 0.06fF
C73987 NOR2X1_LOC_848/Y NOR2X1_LOC_188/A 0.36fF
C73988 INVX1_LOC_117/A NOR2X1_LOC_748/A 0.47fF
C73989 INVX1_LOC_90/A INVX1_LOC_30/A 1.76fF
C73990 INVX1_LOC_64/A NAND2X1_LOC_454/a_36_24# 0.00fF
C73991 NAND2X1_LOC_861/Y NAND2X1_LOC_634/Y 0.13fF
C73992 NOR2X1_LOC_283/a_36_216# INVX1_LOC_30/Y 0.00fF
C73993 NOR2X1_LOC_67/A NOR2X1_LOC_234/Y 0.01fF
C73994 NOR2X1_LOC_536/A NOR2X1_LOC_383/B 0.03fF
C73995 NOR2X1_LOC_717/B INVX1_LOC_198/Y 0.00fF
C73996 NOR2X1_LOC_389/B INVX1_LOC_30/A 0.12fF
C73997 INVX1_LOC_226/Y NAND2X1_LOC_569/A 0.02fF
C73998 NOR2X1_LOC_544/A INVX1_LOC_104/A 0.07fF
C73999 INVX1_LOC_12/Y INVX1_LOC_53/A 0.12fF
C74000 INVX1_LOC_48/Y NOR2X1_LOC_45/B 0.03fF
C74001 NOR2X1_LOC_65/B INVX1_LOC_118/Y 0.07fF
C74002 INVX1_LOC_278/A NAND2X1_LOC_721/A 0.07fF
C74003 NOR2X1_LOC_500/A D_INPUT_0 0.07fF
C74004 INVX1_LOC_5/A INVX1_LOC_36/Y 0.06fF
C74005 NOR2X1_LOC_222/Y NOR2X1_LOC_423/Y 1.23fF
C74006 INVX1_LOC_63/Y NAND2X1_LOC_662/Y 0.01fF
C74007 INVX1_LOC_289/Y INVX1_LOC_264/Y 0.01fF
C74008 NOR2X1_LOC_361/B INVX1_LOC_98/A 0.10fF
C74009 NOR2X1_LOC_643/A INVX1_LOC_315/Y 0.00fF
C74010 NOR2X1_LOC_637/B INVX1_LOC_10/A 0.02fF
C74011 NOR2X1_LOC_490/Y NOR2X1_LOC_384/Y 0.43fF
C74012 INVX1_LOC_25/A INVX1_LOC_280/A 0.34fF
C74013 NOR2X1_LOC_609/A INVX1_LOC_313/Y 0.09fF
C74014 NOR2X1_LOC_617/Y NOR2X1_LOC_71/Y 0.05fF
C74015 INVX1_LOC_35/A NAND2X1_LOC_96/A 0.07fF
C74016 NOR2X1_LOC_270/Y INVX1_LOC_28/A 0.16fF
C74017 INVX1_LOC_155/A INVX1_LOC_10/A 0.70fF
C74018 NOR2X1_LOC_506/Y NOR2X1_LOC_654/A 0.11fF
C74019 INVX1_LOC_271/A INVX1_LOC_118/A 0.32fF
C74020 NOR2X1_LOC_401/B NAND2X1_LOC_181/Y 0.01fF
C74021 NOR2X1_LOC_186/Y VDD 0.31fF
C74022 NAND2X1_LOC_787/A INVX1_LOC_38/A 0.49fF
C74023 NAND2X1_LOC_141/Y NOR2X1_LOC_415/Y 0.18fF
C74024 NAND2X1_LOC_659/A INVX1_LOC_90/Y 0.03fF
C74025 NAND2X1_LOC_731/a_36_24# NAND2X1_LOC_308/Y 0.00fF
C74026 NAND2X1_LOC_288/A NOR2X1_LOC_278/Y 0.10fF
C74027 NAND2X1_LOC_363/B INVX1_LOC_38/A 0.07fF
C74028 NOR2X1_LOC_402/a_36_216# NAND2X1_LOC_181/Y 0.00fF
C74029 NOR2X1_LOC_383/B NAND2X1_LOC_93/B 0.50fF
C74030 INVX1_LOC_1/A NOR2X1_LOC_566/a_36_216# 0.00fF
C74031 NOR2X1_LOC_16/Y INVX1_LOC_1/Y 0.14fF
C74032 NOR2X1_LOC_620/Y INVX1_LOC_89/A 0.02fF
C74033 NAND2X1_LOC_728/Y NAND2X1_LOC_740/B 0.02fF
C74034 INVX1_LOC_84/A INVX1_LOC_87/A 4.35fF
C74035 NAND2X1_LOC_579/A NOR2X1_LOC_670/Y 0.03fF
C74036 NOR2X1_LOC_473/B NOR2X1_LOC_577/Y 0.10fF
C74037 INVX1_LOC_41/A INVX1_LOC_148/Y 0.22fF
C74038 D_INPUT_0 NOR2X1_LOC_84/A 3.29fF
C74039 NOR2X1_LOC_606/Y INVX1_LOC_48/A 0.01fF
C74040 NOR2X1_LOC_440/Y NOR2X1_LOC_612/B 0.02fF
C74041 NOR2X1_LOC_383/B NAND2X1_LOC_425/Y 0.02fF
C74042 NOR2X1_LOC_151/Y INVX1_LOC_198/Y 0.18fF
C74043 NAND2X1_LOC_573/Y VDD 0.29fF
C74044 INVX1_LOC_84/A INVX1_LOC_175/A 0.06fF
C74045 NOR2X1_LOC_510/Y NOR2X1_LOC_60/Y 0.01fF
C74046 NAND2X1_LOC_198/B INVX1_LOC_79/A 0.39fF
C74047 INVX1_LOC_64/A INVX1_LOC_54/A 0.21fF
C74048 INVX1_LOC_93/A NAND2X1_LOC_848/A 0.10fF
C74049 INVX1_LOC_292/A NOR2X1_LOC_405/A 0.00fF
C74050 NOR2X1_LOC_831/B INVX1_LOC_29/Y 0.27fF
C74051 INVX1_LOC_269/A INVX1_LOC_46/A 0.12fF
C74052 INVX1_LOC_1/A INVX1_LOC_139/Y 0.01fF
C74053 NOR2X1_LOC_763/A NAND2X1_LOC_639/A 0.32fF
C74054 INVX1_LOC_49/Y INVX1_LOC_273/A 0.15fF
C74055 NOR2X1_LOC_664/Y INPUT_1 0.00fF
C74056 NOR2X1_LOC_596/A NAND2X1_LOC_832/Y 0.01fF
C74057 INVX1_LOC_279/A INVX1_LOC_179/Y 0.00fF
C74058 NOR2X1_LOC_278/Y INVX1_LOC_19/A 0.03fF
C74059 NOR2X1_LOC_45/Y NOR2X1_LOC_56/Y 0.72fF
C74060 INVX1_LOC_227/A NOR2X1_LOC_203/Y 0.03fF
C74061 NOR2X1_LOC_383/B INVX1_LOC_3/A 0.01fF
C74062 INVX1_LOC_180/A INVX1_LOC_144/A 0.03fF
C74063 NOR2X1_LOC_559/B INPUT_0 0.00fF
C74064 NOR2X1_LOC_739/Y INVX1_LOC_37/A 0.01fF
C74065 NAND2X1_LOC_208/B NOR2X1_LOC_124/A 0.02fF
C74066 NAND2X1_LOC_121/a_36_24# NAND2X1_LOC_472/Y 0.00fF
C74067 NOR2X1_LOC_861/Y NOR2X1_LOC_38/B 0.02fF
C74068 NOR2X1_LOC_36/A NOR2X1_LOC_18/a_36_216# 0.03fF
C74069 INVX1_LOC_90/A NAND2X1_LOC_722/A 0.02fF
C74070 NOR2X1_LOC_655/B INVX1_LOC_171/A 0.01fF
C74071 NOR2X1_LOC_301/A NAND2X1_LOC_74/B 0.03fF
C74072 INVX1_LOC_269/A NAND2X1_LOC_417/a_36_24# 0.00fF
C74073 INVX1_LOC_27/A INVX1_LOC_118/A 0.01fF
C74074 INVX1_LOC_17/Y NAND2X1_LOC_489/Y 0.01fF
C74075 NOR2X1_LOC_441/Y INVX1_LOC_147/Y 0.00fF
C74076 INVX1_LOC_119/Y NOR2X1_LOC_591/A 0.12fF
C74077 NOR2X1_LOC_245/a_36_216# NOR2X1_LOC_773/Y 0.01fF
C74078 NOR2X1_LOC_824/A INVX1_LOC_118/A 0.62fF
C74079 INVX1_LOC_200/Y NAND2X1_LOC_489/Y 0.01fF
C74080 INVX1_LOC_177/Y NOR2X1_LOC_139/Y 0.04fF
C74081 NOR2X1_LOC_78/B NOR2X1_LOC_214/B 0.95fF
C74082 NOR2X1_LOC_710/B INVX1_LOC_117/A 0.00fF
C74083 NAND2X1_LOC_198/B INVX1_LOC_91/A 0.10fF
C74084 INVX1_LOC_1/A INVX1_LOC_280/A 0.09fF
C74085 D_INPUT_1 INVX1_LOC_63/A 0.08fF
C74086 NOR2X1_LOC_441/Y INVX1_LOC_20/A 0.03fF
C74087 NOR2X1_LOC_45/Y VDD 0.17fF
C74088 INVX1_LOC_121/A INVX1_LOC_32/Y 0.00fF
C74089 NOR2X1_LOC_208/Y NOR2X1_LOC_144/a_36_216# 0.00fF
C74090 NOR2X1_LOC_388/Y NOR2X1_LOC_188/A 0.05fF
C74091 NOR2X1_LOC_757/Y INVX1_LOC_313/Y 0.00fF
C74092 INVX1_LOC_279/A NOR2X1_LOC_561/Y 0.10fF
C74093 INVX1_LOC_25/Y NOR2X1_LOC_76/A 0.02fF
C74094 NAND2X1_LOC_190/Y INVX1_LOC_9/A 0.01fF
C74095 INVX1_LOC_215/Y NOR2X1_LOC_816/Y 0.03fF
C74096 NOR2X1_LOC_355/B NOR2X1_LOC_577/Y 0.00fF
C74097 NOR2X1_LOC_6/B INPUT_0 0.13fF
C74098 NOR2X1_LOC_191/B NAND2X1_LOC_642/Y 0.15fF
C74099 INVX1_LOC_170/A VDD 0.12fF
C74100 INVX1_LOC_33/A NOR2X1_LOC_356/a_36_216# 0.00fF
C74101 NAND2X1_LOC_619/a_36_24# INVX1_LOC_15/A 0.00fF
C74102 NAND2X1_LOC_527/a_36_24# NAND2X1_LOC_96/A 0.00fF
C74103 NOR2X1_LOC_262/Y INVX1_LOC_93/Y 0.07fF
C74104 INPUT_1 INVX1_LOC_137/A 0.01fF
C74105 INVX1_LOC_175/A INVX1_LOC_15/A 0.02fF
C74106 NAND2X1_LOC_425/Y NOR2X1_LOC_463/a_36_216# 0.01fF
C74107 NAND2X1_LOC_303/B INPUT_5 0.06fF
C74108 INVX1_LOC_128/Y NOR2X1_LOC_334/Y 0.13fF
C74109 INVX1_LOC_47/Y INVX1_LOC_26/A 0.10fF
C74110 NOR2X1_LOC_843/A INVX1_LOC_186/A 0.03fF
C74111 NOR2X1_LOC_652/Y INVX1_LOC_63/A 0.07fF
C74112 NOR2X1_LOC_389/A INVX1_LOC_9/A 0.03fF
C74113 INVX1_LOC_83/A NOR2X1_LOC_814/Y 0.03fF
C74114 INVX1_LOC_234/A INPUT_1 0.03fF
C74115 INVX1_LOC_111/Y INVX1_LOC_69/Y 0.10fF
C74116 INVX1_LOC_30/A NAND2X1_LOC_849/B 0.08fF
C74117 NOR2X1_LOC_384/Y NOR2X1_LOC_813/Y 0.79fF
C74118 INVX1_LOC_53/A NOR2X1_LOC_842/a_36_216# 0.00fF
C74119 NOR2X1_LOC_817/Y NAND2X1_LOC_817/a_36_24# -0.02fF
C74120 INVX1_LOC_244/Y INVX1_LOC_37/A 0.01fF
C74121 NAND2X1_LOC_656/A NAND2X1_LOC_611/a_36_24# 0.01fF
C74122 INVX1_LOC_30/A INVX1_LOC_38/A 0.35fF
C74123 INVX1_LOC_104/A NOR2X1_LOC_139/Y 0.03fF
C74124 INVX1_LOC_34/A NOR2X1_LOC_124/A 0.01fF
C74125 NOR2X1_LOC_19/B NAND2X1_LOC_462/B 0.00fF
C74126 NOR2X1_LOC_191/A INVX1_LOC_6/A 0.26fF
C74127 NOR2X1_LOC_186/Y INVX1_LOC_133/A 0.04fF
C74128 INVX1_LOC_286/A NAND2X1_LOC_850/Y 0.10fF
C74129 INVX1_LOC_2/A NOR2X1_LOC_528/Y 0.42fF
C74130 NOR2X1_LOC_561/Y INVX1_LOC_182/Y 0.01fF
C74131 INVX1_LOC_4/A NAND2X1_LOC_215/A 0.07fF
C74132 NOR2X1_LOC_160/B INVX1_LOC_92/A 0.10fF
C74133 NOR2X1_LOC_384/Y INVX1_LOC_280/A 0.03fF
C74134 INVX1_LOC_177/A NOR2X1_LOC_78/A 0.05fF
C74135 INVX1_LOC_289/Y INVX1_LOC_84/A 0.11fF
C74136 INVX1_LOC_249/A NAND2X1_LOC_605/a_36_24# 0.01fF
C74137 NOR2X1_LOC_78/B NOR2X1_LOC_741/A 0.01fF
C74138 INVX1_LOC_64/A NOR2X1_LOC_48/B 0.17fF
C74139 NOR2X1_LOC_45/B NOR2X1_LOC_482/Y 0.14fF
C74140 INVX1_LOC_132/A VDD 0.16fF
C74141 NOR2X1_LOC_374/A VDD 0.09fF
C74142 NOR2X1_LOC_226/A NOR2X1_LOC_528/Y 0.10fF
C74143 INVX1_LOC_30/Y INPUT_0 2.31fF
C74144 INVX1_LOC_27/A NAND2X1_LOC_63/Y 0.02fF
C74145 NOR2X1_LOC_837/B NAND2X1_LOC_96/A 0.10fF
C74146 NOR2X1_LOC_512/Y NOR2X1_LOC_536/A 0.03fF
C74147 NAND2X1_LOC_671/a_36_24# INVX1_LOC_201/A 0.00fF
C74148 NOR2X1_LOC_710/A NOR2X1_LOC_155/A 0.01fF
C74149 NOR2X1_LOC_144/Y INVX1_LOC_76/A 0.01fF
C74150 NOR2X1_LOC_93/Y NOR2X1_LOC_671/Y 0.01fF
C74151 INVX1_LOC_256/A NOR2X1_LOC_127/Y 0.10fF
C74152 NOR2X1_LOC_82/A INVX1_LOC_84/A 0.55fF
C74153 INVX1_LOC_62/Y INVX1_LOC_9/A 0.07fF
C74154 NOR2X1_LOC_338/Y NOR2X1_LOC_351/Y 0.11fF
C74155 INVX1_LOC_18/A NOR2X1_LOC_641/Y 0.01fF
C74156 NOR2X1_LOC_19/B INPUT_1 2.89fF
C74157 INVX1_LOC_130/Y INVX1_LOC_54/A 0.03fF
C74158 INVX1_LOC_178/A INVX1_LOC_102/A 0.10fF
C74159 NOR2X1_LOC_381/Y NOR2X1_LOC_84/B 0.00fF
C74160 NOR2X1_LOC_68/A INVX1_LOC_274/A 0.08fF
C74161 NOR2X1_LOC_180/B NOR2X1_LOC_439/B 0.01fF
C74162 NOR2X1_LOC_596/A INVX1_LOC_9/A 0.01fF
C74163 INVX1_LOC_150/Y NOR2X1_LOC_814/A 0.21fF
C74164 INVX1_LOC_225/A VDD 0.59fF
C74165 INVX1_LOC_95/A NAND2X1_LOC_850/Y 0.05fF
C74166 NOR2X1_LOC_376/A NOR2X1_LOC_89/A 0.01fF
C74167 NOR2X1_LOC_334/Y NOR2X1_LOC_717/A 0.08fF
C74168 NOR2X1_LOC_288/A VDD 0.16fF
C74169 INVX1_LOC_53/Y INVX1_LOC_91/A 0.09fF
C74170 NAND2X1_LOC_632/B NOR2X1_LOC_536/A 0.03fF
C74171 NOR2X1_LOC_631/B NOR2X1_LOC_352/Y 0.01fF
C74172 NOR2X1_LOC_265/a_36_216# NAND2X1_LOC_642/Y 0.01fF
C74173 INVX1_LOC_135/A NOR2X1_LOC_188/A 0.03fF
C74174 NOR2X1_LOC_180/B INVX1_LOC_75/A 0.07fF
C74175 NOR2X1_LOC_243/Y VDD 0.05fF
C74176 NOR2X1_LOC_152/Y INVX1_LOC_118/Y 0.55fF
C74177 NAND2X1_LOC_363/B NAND2X1_LOC_223/A 0.07fF
C74178 NOR2X1_LOC_134/Y NAND2X1_LOC_477/Y 0.02fF
C74179 INVX1_LOC_290/A NOR2X1_LOC_45/B 0.13fF
C74180 INVX1_LOC_88/Y NAND2X1_LOC_472/Y 0.03fF
C74181 NOR2X1_LOC_655/B INVX1_LOC_20/A 0.00fF
C74182 INVX1_LOC_89/A NOR2X1_LOC_589/Y 0.01fF
C74183 INVX1_LOC_85/Y NOR2X1_LOC_74/A 0.03fF
C74184 INVX1_LOC_17/A NAND2X1_LOC_74/B 0.09fF
C74185 NOR2X1_LOC_254/A INVX1_LOC_186/Y 0.15fF
C74186 INVX1_LOC_14/A NOR2X1_LOC_89/A 0.23fF
C74187 INVX1_LOC_54/Y NOR2X1_LOC_266/B 0.00fF
C74188 INVX1_LOC_69/Y NOR2X1_LOC_137/A 0.03fF
C74189 NOR2X1_LOC_197/A INVX1_LOC_19/A 0.00fF
C74190 NOR2X1_LOC_209/Y VDD 0.66fF
C74191 NAND2X1_LOC_803/B INVX1_LOC_272/A 0.02fF
C74192 NOR2X1_LOC_781/B INVX1_LOC_91/A 0.57fF
C74193 NOR2X1_LOC_693/Y NOR2X1_LOC_754/Y 0.02fF
C74194 INVX1_LOC_103/A INVX1_LOC_109/Y 1.03fF
C74195 INVX1_LOC_145/Y INVX1_LOC_91/A 0.02fF
C74196 NOR2X1_LOC_785/Y NOR2X1_LOC_78/A 0.01fF
C74197 NAND2X1_LOC_374/Y INVX1_LOC_37/A 0.07fF
C74198 NOR2X1_LOC_294/Y NAND2X1_LOC_206/Y 0.01fF
C74199 INVX1_LOC_35/A NAND2X1_LOC_99/A 0.06fF
C74200 INVX1_LOC_73/A INVX1_LOC_75/A 0.07fF
C74201 VDD NAND2X1_LOC_852/Y 2.08fF
C74202 INVX1_LOC_22/A NAND2X1_LOC_836/Y 0.21fF
C74203 NOR2X1_LOC_590/A INVX1_LOC_272/A 0.07fF
C74204 NOR2X1_LOC_78/B INVX1_LOC_12/Y 0.03fF
C74205 NOR2X1_LOC_318/A NOR2X1_LOC_109/Y 0.17fF
C74206 INVX1_LOC_270/A NOR2X1_LOC_678/A 0.03fF
C74207 NAND2X1_LOC_175/Y NOR2X1_LOC_406/A 0.03fF
C74208 NAND2X1_LOC_555/Y NAND2X1_LOC_207/Y 0.05fF
C74209 NOR2X1_LOC_816/A INVX1_LOC_102/A 0.11fF
C74210 NAND2X1_LOC_714/B INVX1_LOC_94/Y 0.03fF
C74211 NAND2X1_LOC_722/A INVX1_LOC_38/A 0.10fF
C74212 INVX1_LOC_71/A NAND2X1_LOC_572/B 0.10fF
C74213 INVX1_LOC_27/A NOR2X1_LOC_631/Y 0.08fF
C74214 INVX1_LOC_279/A INVX1_LOC_76/A -0.01fF
C74215 NOR2X1_LOC_553/B INVX1_LOC_37/A 0.03fF
C74216 NOR2X1_LOC_31/a_36_216# INPUT_5 0.00fF
C74217 INVX1_LOC_134/A INVX1_LOC_15/A 0.10fF
C74218 NOR2X1_LOC_99/B INVX1_LOC_20/A 0.07fF
C74219 NOR2X1_LOC_52/Y INVX1_LOC_109/A 0.02fF
C74220 INVX1_LOC_305/A NOR2X1_LOC_633/A 0.13fF
C74221 NAND2X1_LOC_858/B NOR2X1_LOC_167/Y 0.14fF
C74222 NOR2X1_LOC_332/A INVX1_LOC_36/Y 0.15fF
C74223 INVX1_LOC_58/A NOR2X1_LOC_304/Y 0.20fF
C74224 NOR2X1_LOC_220/A INVX1_LOC_9/A 0.10fF
C74225 NAND2X1_LOC_511/a_36_24# NAND2X1_LOC_782/B 0.01fF
C74226 NAND2X1_LOC_850/Y INVX1_LOC_54/A 0.07fF
C74227 INVX1_LOC_33/A NAND2X1_LOC_475/Y 0.00fF
C74228 NOR2X1_LOC_113/B NOR2X1_LOC_114/A 0.00fF
C74229 NAND2X1_LOC_474/Y INVX1_LOC_57/A 0.09fF
C74230 NOR2X1_LOC_214/B INVX1_LOC_46/A 0.00fF
C74231 NOR2X1_LOC_348/Y NOR2X1_LOC_383/B 0.07fF
C74232 INVX1_LOC_56/Y INVX1_LOC_127/A 0.07fF
C74233 NAND2X1_LOC_36/A INVX1_LOC_15/A 0.42fF
C74234 NOR2X1_LOC_548/Y INVX1_LOC_9/A 0.07fF
C74235 INVX1_LOC_31/A NOR2X1_LOC_681/a_36_216# 0.00fF
C74236 INVX1_LOC_21/A NOR2X1_LOC_32/B 0.07fF
C74237 NAND2X1_LOC_84/Y NOR2X1_LOC_89/A 0.02fF
C74238 NOR2X1_LOC_226/A NOR2X1_LOC_216/B 0.10fF
C74239 NOR2X1_LOC_721/Y NAND2X1_LOC_642/Y 0.02fF
C74240 NOR2X1_LOC_552/A NOR2X1_LOC_188/A 0.12fF
C74241 INVX1_LOC_89/A INVX1_LOC_117/A 0.77fF
C74242 INVX1_LOC_208/A INVX1_LOC_92/A 0.15fF
C74243 INVX1_LOC_21/A NOR2X1_LOC_639/B 0.08fF
C74244 INPUT_0 NOR2X1_LOC_124/A 0.02fF
C74245 NOR2X1_LOC_637/B INVX1_LOC_12/A 0.01fF
C74246 NOR2X1_LOC_552/A NOR2X1_LOC_548/B 0.10fF
C74247 NOR2X1_LOC_576/B NAND2X1_LOC_770/a_36_24# 0.03fF
C74248 INVX1_LOC_272/Y INVX1_LOC_57/A 0.07fF
C74249 NOR2X1_LOC_807/B NOR2X1_LOC_383/B 0.09fF
C74250 INVX1_LOC_256/A NOR2X1_LOC_383/B 0.08fF
C74251 NOR2X1_LOC_793/A INVX1_LOC_53/A 0.98fF
C74252 NOR2X1_LOC_647/A INVX1_LOC_230/Y 0.00fF
C74253 INVX1_LOC_30/A NAND2X1_LOC_223/A 0.01fF
C74254 NOR2X1_LOC_657/Y NAND2X1_LOC_454/Y 0.02fF
C74255 INVX1_LOC_39/A NAND2X1_LOC_214/B 0.01fF
C74256 NAND2X1_LOC_9/Y INVX1_LOC_269/A 0.01fF
C74257 NOR2X1_LOC_793/Y NOR2X1_LOC_598/B 0.46fF
C74258 INVX1_LOC_116/A INVX1_LOC_32/A 0.01fF
C74259 INVX1_LOC_233/A INVX1_LOC_269/A 0.19fF
C74260 INVX1_LOC_278/Y INVX1_LOC_84/A 0.07fF
C74261 NAND2X1_LOC_741/Y GATE_741 0.00fF
C74262 INVX1_LOC_250/A NAND2X1_LOC_175/Y 0.03fF
C74263 NOR2X1_LOC_690/A NAND2X1_LOC_254/Y 0.25fF
C74264 INVX1_LOC_10/A NOR2X1_LOC_510/B 0.09fF
C74265 NOR2X1_LOC_78/A INVX1_LOC_65/A 0.01fF
C74266 NOR2X1_LOC_667/A NAND2X1_LOC_604/a_36_24# 0.00fF
C74267 INVX1_LOC_39/A INVX1_LOC_27/A 0.06fF
C74268 INVX1_LOC_136/A NOR2X1_LOC_301/A 0.07fF
C74269 D_INPUT_0 NOR2X1_LOC_78/Y 0.01fF
C74270 INVX1_LOC_278/A NOR2X1_LOC_82/A 0.36fF
C74271 INVX1_LOC_232/Y INVX1_LOC_19/A 0.14fF
C74272 NAND2X1_LOC_638/Y NAND2X1_LOC_637/Y 0.01fF
C74273 NOR2X1_LOC_541/Y INVX1_LOC_58/Y 0.02fF
C74274 NAND2X1_LOC_361/Y INVX1_LOC_32/A 0.03fF
C74275 NOR2X1_LOC_612/B NOR2X1_LOC_89/A 0.00fF
C74276 NOR2X1_LOC_160/B INVX1_LOC_53/A 0.49fF
C74277 INVX1_LOC_58/A NAND2X1_LOC_711/Y 0.03fF
C74278 INVX1_LOC_45/A NOR2X1_LOC_654/A 0.03fF
C74279 NOR2X1_LOC_61/B NAND2X1_LOC_58/a_36_24# 0.00fF
C74280 D_INPUT_0 INVX1_LOC_35/Y 0.38fF
C74281 NOR2X1_LOC_844/A NOR2X1_LOC_861/Y 0.17fF
C74282 NAND2X1_LOC_840/B INVX1_LOC_49/Y 0.27fF
C74283 INVX1_LOC_64/A NAND2X1_LOC_350/A 0.07fF
C74284 NOR2X1_LOC_186/Y NOR2X1_LOC_361/B 0.10fF
C74285 NOR2X1_LOC_262/Y INVX1_LOC_87/A 0.01fF
C74286 NAND2X1_LOC_13/a_36_24# INVX1_LOC_5/A 0.00fF
C74287 INVX1_LOC_91/A NOR2X1_LOC_585/Y 0.01fF
C74288 NOR2X1_LOC_303/Y NAND2X1_LOC_71/a_36_24# 0.00fF
C74289 NOR2X1_LOC_142/Y INVX1_LOC_4/A 0.70fF
C74290 NOR2X1_LOC_78/A NAND2X1_LOC_267/B 0.00fF
C74291 NOR2X1_LOC_328/Y NOR2X1_LOC_36/B 0.03fF
C74292 NOR2X1_LOC_703/Y INVX1_LOC_117/A -0.00fF
C74293 NOR2X1_LOC_123/B NAND2X1_LOC_572/B 0.01fF
C74294 INPUT_1 NOR2X1_LOC_216/B 0.05fF
C74295 NOR2X1_LOC_188/A INVX1_LOC_280/A 0.07fF
C74296 INVX1_LOC_78/Y NAND2X1_LOC_472/Y 0.02fF
C74297 INVX1_LOC_291/Y INVX1_LOC_20/A 0.01fF
C74298 NOR2X1_LOC_815/A NOR2X1_LOC_331/B 0.05fF
C74299 INVX1_LOC_125/Y INVX1_LOC_129/Y 0.00fF
C74300 NOR2X1_LOC_92/Y NAND2X1_LOC_725/B 0.07fF
C74301 INVX1_LOC_64/A NOR2X1_LOC_441/Y 0.05fF
C74302 INVX1_LOC_45/A INVX1_LOC_58/Y 0.04fF
C74303 NOR2X1_LOC_773/Y INVX1_LOC_102/A 0.11fF
C74304 INVX1_LOC_282/A INVX1_LOC_54/A 0.02fF
C74305 NAND2X1_LOC_570/a_36_24# INVX1_LOC_15/A 0.00fF
C74306 NOR2X1_LOC_229/Y INVX1_LOC_12/A 0.12fF
C74307 NOR2X1_LOC_795/Y NOR2X1_LOC_801/B 0.08fF
C74308 NAND2X1_LOC_573/Y NOR2X1_LOC_361/B 0.35fF
C74309 VDD NAND2X1_LOC_642/Y 1.44fF
C74310 NOR2X1_LOC_568/A INVX1_LOC_58/Y 0.09fF
C74311 NAND2X1_LOC_850/Y NOR2X1_LOC_48/B 0.06fF
C74312 NOR2X1_LOC_100/A INVX1_LOC_15/A 0.33fF
C74313 INVX1_LOC_36/A NOR2X1_LOC_678/A 0.03fF
C74314 NOR2X1_LOC_312/Y NOR2X1_LOC_653/Y 0.13fF
C74315 NAND2X1_LOC_7/Y INVX1_LOC_26/Y 0.02fF
C74316 NAND2X1_LOC_808/A NOR2X1_LOC_605/A 0.07fF
C74317 NOR2X1_LOC_706/A INVX1_LOC_92/A 0.39fF
C74318 INVX1_LOC_61/Y NOR2X1_LOC_293/a_36_216# 0.01fF
C74319 NOR2X1_LOC_510/Y NOR2X1_LOC_45/Y 0.00fF
C74320 D_INPUT_0 NOR2X1_LOC_721/B 0.00fF
C74321 NOR2X1_LOC_480/A NOR2X1_LOC_476/B 0.10fF
C74322 NOR2X1_LOC_242/A NOR2X1_LOC_160/B 0.05fF
C74323 INVX1_LOC_143/Y NOR2X1_LOC_857/A 0.07fF
C74324 INVX1_LOC_224/Y NOR2X1_LOC_419/Y 0.03fF
C74325 NOR2X1_LOC_168/B NAND2X1_LOC_615/a_36_24# 0.00fF
C74326 NOR2X1_LOC_655/B INVX1_LOC_4/A 0.39fF
C74327 NAND2X1_LOC_570/Y NAND2X1_LOC_618/Y 0.05fF
C74328 NOR2X1_LOC_335/A INVX1_LOC_270/A 0.05fF
C74329 INVX1_LOC_11/A INVX1_LOC_14/A 0.13fF
C74330 NOR2X1_LOC_574/a_36_216# INVX1_LOC_78/A 0.00fF
C74331 INVX1_LOC_266/A INVX1_LOC_225/Y 0.10fF
C74332 NAND2X1_LOC_59/a_36_24# INVX1_LOC_15/A 0.00fF
C74333 INVX1_LOC_35/A NAND2X1_LOC_656/A 0.18fF
C74334 NOR2X1_LOC_309/Y NOR2X1_LOC_318/A 0.01fF
C74335 VDD D_GATE_662 0.23fF
C74336 NOR2X1_LOC_815/A NOR2X1_LOC_592/B 0.01fF
C74337 NOR2X1_LOC_208/Y NOR2X1_LOC_678/A 0.03fF
C74338 NOR2X1_LOC_176/Y INVX1_LOC_20/A 0.05fF
C74339 INVX1_LOC_21/A NAND2X1_LOC_510/A 0.10fF
C74340 NOR2X1_LOC_299/Y NAND2X1_LOC_402/a_36_24# 0.00fF
C74341 NAND2X1_LOC_361/Y NOR2X1_LOC_622/A 0.02fF
C74342 NOR2X1_LOC_718/B NOR2X1_LOC_727/B 0.09fF
C74343 NOR2X1_LOC_788/B INVX1_LOC_29/A 0.07fF
C74344 INVX1_LOC_12/Y INVX1_LOC_46/A 0.03fF
C74345 NOR2X1_LOC_719/A NOR2X1_LOC_38/B 0.00fF
C74346 VDD NOR2X1_LOC_863/A 0.24fF
C74347 NOR2X1_LOC_716/B NAND2X1_LOC_793/B 1.55fF
C74348 INVX1_LOC_46/A NOR2X1_LOC_492/Y 0.38fF
C74349 NAND2X1_LOC_363/B INVX1_LOC_33/A 0.07fF
C74350 NOR2X1_LOC_317/B INVX1_LOC_53/A 0.01fF
C74351 NOR2X1_LOC_135/Y INVX1_LOC_29/A 0.00fF
C74352 NAND2X1_LOC_387/B INVX1_LOC_1/A 0.01fF
C74353 INVX1_LOC_7/A NOR2X1_LOC_38/B 2.07fF
C74354 INVX1_LOC_35/A NOR2X1_LOC_725/a_36_216# 0.00fF
C74355 NOR2X1_LOC_590/A INVX1_LOC_150/Y 0.14fF
C74356 INVX1_LOC_316/Y NOR2X1_LOC_29/a_36_216# 0.00fF
C74357 VDD NOR2X1_LOC_271/Y 0.12fF
C74358 INVX1_LOC_226/Y NOR2X1_LOC_55/a_36_216# 0.00fF
C74359 INVX1_LOC_64/A NOR2X1_LOC_142/Y 0.01fF
C74360 INVX1_LOC_133/Y NOR2X1_LOC_125/Y 0.02fF
C74361 INVX1_LOC_11/A NOR2X1_LOC_717/Y 0.05fF
C74362 INVX1_LOC_89/A INVX1_LOC_3/Y 0.09fF
C74363 NOR2X1_LOC_99/B INVX1_LOC_4/A 0.07fF
C74364 NOR2X1_LOC_15/Y NOR2X1_LOC_518/a_36_216# 0.00fF
C74365 INVX1_LOC_140/A INVX1_LOC_102/A 0.10fF
C74366 INVX1_LOC_196/A INVX1_LOC_23/A 0.01fF
C74367 NOR2X1_LOC_773/Y NOR2X1_LOC_280/a_36_216# 0.00fF
C74368 INVX1_LOC_17/A INVX1_LOC_136/A 0.18fF
C74369 INVX1_LOC_298/Y NOR2X1_LOC_632/Y 0.10fF
C74370 INVX1_LOC_166/A INVX1_LOC_197/Y 0.05fF
C74371 NAND2X1_LOC_67/Y NOR2X1_LOC_596/A 0.03fF
C74372 INVX1_LOC_2/Y NOR2X1_LOC_78/a_36_216# 0.00fF
C74373 NAND2X1_LOC_725/B NAND2X1_LOC_837/Y 0.07fF
C74374 INVX1_LOC_13/A NAND2X1_LOC_23/a_36_24# 0.00fF
C74375 INVX1_LOC_22/A NOR2X1_LOC_699/a_36_216# 0.00fF
C74376 NAND2X1_LOC_778/Y INVX1_LOC_34/A 0.35fF
C74377 INVX1_LOC_226/Y INVX1_LOC_57/A 0.11fF
C74378 INVX1_LOC_5/A INVX1_LOC_85/A 0.01fF
C74379 INVX1_LOC_21/A INVX1_LOC_155/Y 0.01fF
C74380 NAND2X1_LOC_350/B INVX1_LOC_53/A 0.43fF
C74381 INVX1_LOC_136/A NOR2X1_LOC_471/Y 0.48fF
C74382 NOR2X1_LOC_624/A INVX1_LOC_27/A 0.00fF
C74383 INVX1_LOC_13/Y INVX1_LOC_104/A 0.03fF
C74384 NOR2X1_LOC_254/A INVX1_LOC_18/A 0.07fF
C74385 NAND2X1_LOC_740/Y INVX1_LOC_240/A 0.02fF
C74386 NOR2X1_LOC_636/a_36_216# NAND2X1_LOC_149/Y 0.01fF
C74387 INVX1_LOC_64/A NOR2X1_LOC_655/B 0.02fF
C74388 INVX1_LOC_200/Y NAND2X1_LOC_564/B 0.14fF
C74389 NOR2X1_LOC_562/B INVX1_LOC_186/Y 0.10fF
C74390 INVX1_LOC_21/A NOR2X1_LOC_720/B 0.01fF
C74391 INVX1_LOC_208/A INVX1_LOC_53/A 0.10fF
C74392 D_INPUT_1 INVX1_LOC_1/Y 0.14fF
C74393 INVX1_LOC_182/A INVX1_LOC_4/A 0.50fF
C74394 D_GATE_366 INVX1_LOC_78/A 0.03fF
C74395 NAND2X1_LOC_363/B INVX1_LOC_40/A 0.12fF
C74396 INVX1_LOC_59/Y INVX1_LOC_84/A 0.10fF
C74397 NOR2X1_LOC_486/a_36_216# NOR2X1_LOC_68/A 0.00fF
C74398 NOR2X1_LOC_516/B INVX1_LOC_53/A 0.16fF
C74399 NOR2X1_LOC_19/B NAND2X1_LOC_618/Y 0.61fF
C74400 INVX1_LOC_112/A INVX1_LOC_84/A 0.01fF
C74401 NOR2X1_LOC_419/Y NOR2X1_LOC_103/Y 0.10fF
C74402 NOR2X1_LOC_75/Y INVX1_LOC_71/A 0.03fF
C74403 INVX1_LOC_24/A NAND2X1_LOC_114/B 0.46fF
C74404 INVX1_LOC_2/A INVX1_LOC_93/A 0.07fF
C74405 NOR2X1_LOC_498/Y NAND2X1_LOC_725/B 0.22fF
C74406 INVX1_LOC_34/A NOR2X1_LOC_15/Y 0.10fF
C74407 INVX1_LOC_10/A INVX1_LOC_57/A 2.98fF
C74408 NOR2X1_LOC_78/A NOR2X1_LOC_830/Y 0.01fF
C74409 INVX1_LOC_286/Y NOR2X1_LOC_91/Y 0.11fF
C74410 NOR2X1_LOC_160/B INVX1_LOC_184/A 0.03fF
C74411 NAND2X1_LOC_162/a_36_24# INVX1_LOC_78/A 0.00fF
C74412 NOR2X1_LOC_124/A NOR2X1_LOC_84/B -0.01fF
C74413 NOR2X1_LOC_32/B NOR2X1_LOC_521/Y 0.02fF
C74414 NOR2X1_LOC_226/A INVX1_LOC_93/A 0.44fF
C74415 NAND2X1_LOC_553/A NAND2X1_LOC_563/A 0.01fF
C74416 NOR2X1_LOC_238/Y INVX1_LOC_31/A 0.03fF
C74417 INVX1_LOC_50/A NOR2X1_LOC_246/A 0.03fF
C74418 INVX1_LOC_24/A INVX1_LOC_141/Y 0.03fF
C74419 INVX1_LOC_33/A NOR2X1_LOC_457/A 0.36fF
C74420 NAND2X1_LOC_287/B NOR2X1_LOC_653/Y 0.17fF
C74421 INVX1_LOC_225/A NOR2X1_LOC_361/B 0.81fF
C74422 NOR2X1_LOC_455/Y INVX1_LOC_279/A 0.03fF
C74423 NAND2X1_LOC_543/Y NAND2X1_LOC_552/A 0.01fF
C74424 NAND2X1_LOC_848/A INVX1_LOC_35/Y 0.10fF
C74425 INVX1_LOC_22/A NOR2X1_LOC_304/a_36_216# 0.02fF
C74426 NAND2X1_LOC_784/A INVX1_LOC_135/A 0.10fF
C74427 NOR2X1_LOC_795/Y INVX1_LOC_1/A 0.01fF
C74428 INVX1_LOC_88/A INVX1_LOC_104/A 0.10fF
C74429 INVX1_LOC_14/A NOR2X1_LOC_52/B 0.21fF
C74430 NAND2X1_LOC_860/A NOR2X1_LOC_278/a_36_216# 0.01fF
C74431 INVX1_LOC_178/Y NOR2X1_LOC_662/A 0.03fF
C74432 INVX1_LOC_58/A INVX1_LOC_89/A 0.79fF
C74433 NAND2X1_LOC_860/A D_INPUT_0 0.03fF
C74434 NOR2X1_LOC_74/A NAND2X1_LOC_454/Y 0.07fF
C74435 NAND2X1_LOC_208/a_36_24# INVX1_LOC_16/A 0.00fF
C74436 INVX1_LOC_5/A NAND2X1_LOC_662/Y 0.05fF
C74437 INVX1_LOC_50/A INVX1_LOC_55/Y 0.03fF
C74438 NOR2X1_LOC_155/A NOR2X1_LOC_729/A 0.00fF
C74439 INVX1_LOC_1/Y NOR2X1_LOC_652/Y 0.64fF
C74440 NOR2X1_LOC_848/Y NOR2X1_LOC_87/B 0.00fF
C74441 NAND2X1_LOC_287/B INVX1_LOC_19/A 0.07fF
C74442 NOR2X1_LOC_445/Y INVX1_LOC_292/A 0.01fF
C74443 NOR2X1_LOC_15/Y NAND2X1_LOC_231/Y 0.01fF
C74444 NOR2X1_LOC_536/A NAND2X1_LOC_267/a_36_24# 0.00fF
C74445 NOR2X1_LOC_836/Y NAND2X1_LOC_364/Y 0.02fF
C74446 NOR2X1_LOC_272/Y INVX1_LOC_56/Y 0.01fF
C74447 D_INPUT_0 NOR2X1_LOC_634/Y 0.03fF
C74448 NOR2X1_LOC_644/Y NOR2X1_LOC_205/Y 0.02fF
C74449 NAND2X1_LOC_391/Y INVX1_LOC_16/A 0.00fF
C74450 NAND2X1_LOC_433/a_36_24# INVX1_LOC_76/A 0.01fF
C74451 NOR2X1_LOC_858/B INVX1_LOC_19/A 0.06fF
C74452 INVX1_LOC_224/Y NOR2X1_LOC_120/a_36_216# 0.00fF
C74453 VDD NOR2X1_LOC_48/Y 0.58fF
C74454 INVX1_LOC_45/A NOR2X1_LOC_537/A 0.01fF
C74455 INVX1_LOC_64/A NOR2X1_LOC_99/B 0.07fF
C74456 NOR2X1_LOC_45/B NOR2X1_LOC_467/A 0.02fF
C74457 INVX1_LOC_39/A INVX1_LOC_137/A 0.00fF
C74458 INVX1_LOC_37/A INVX1_LOC_125/A 0.00fF
C74459 NOR2X1_LOC_82/A NOR2X1_LOC_63/a_36_216# 0.00fF
C74460 INVX1_LOC_179/A NAND2X1_LOC_93/B 0.03fF
C74461 NAND2X1_LOC_21/Y NAND2X1_LOC_36/A 1.27fF
C74462 INVX1_LOC_24/Y NOR2X1_LOC_544/A 0.01fF
C74463 INVX1_LOC_45/A NOR2X1_LOC_716/B 0.08fF
C74464 INVX1_LOC_2/A NOR2X1_LOC_513/Y 0.01fF
C74465 INVX1_LOC_33/A INVX1_LOC_30/A 0.20fF
C74466 NOR2X1_LOC_636/B NAND2X1_LOC_451/Y 0.35fF
C74467 NOR2X1_LOC_186/Y NAND2X1_LOC_573/A 0.22fF
C74468 INVX1_LOC_281/Y INVX1_LOC_186/Y 0.01fF
C74469 NOR2X1_LOC_759/A INVX1_LOC_105/A 0.78fF
C74470 NOR2X1_LOC_828/A NAND2X1_LOC_599/a_36_24# 0.00fF
C74471 NOR2X1_LOC_78/A INVX1_LOC_4/Y 0.09fF
C74472 NOR2X1_LOC_349/A NOR2X1_LOC_227/A 0.13fF
C74473 NOR2X1_LOC_574/A INVX1_LOC_31/A 0.04fF
C74474 INVX1_LOC_309/Y NAND2X1_LOC_837/Y 0.01fF
C74475 INVX1_LOC_39/A INVX1_LOC_234/A 0.02fF
C74476 INVX1_LOC_237/A NAND2X1_LOC_735/B 0.01fF
C74477 GATE_741 NOR2X1_LOC_298/Y 0.56fF
C74478 NAND2X1_LOC_741/Y NOR2X1_LOC_299/Y 0.01fF
C74479 NAND2X1_LOC_477/Y INVX1_LOC_118/A 0.10fF
C74480 NOR2X1_LOC_458/a_36_216# NOR2X1_LOC_151/Y -0.00fF
C74481 INVX1_LOC_55/Y NAND2X1_LOC_72/Y 0.18fF
C74482 VDD NAND2X1_LOC_792/B 0.01fF
C74483 INVX1_LOC_35/A NOR2X1_LOC_329/B 0.07fF
C74484 NOR2X1_LOC_455/Y INVX1_LOC_182/Y 0.02fF
C74485 NOR2X1_LOC_612/Y NOR2X1_LOC_814/A 0.00fF
C74486 INVX1_LOC_228/Y INVX1_LOC_316/Y 0.05fF
C74487 NAND2X1_LOC_573/Y NAND2X1_LOC_573/A 0.69fF
C74488 NOR2X1_LOC_78/B NOR2X1_LOC_160/B 0.37fF
C74489 NAND2X1_LOC_726/a_36_24# NAND2X1_LOC_308/Y 0.00fF
C74490 NAND2X1_LOC_244/A INVX1_LOC_3/Y 0.06fF
C74491 NOR2X1_LOC_500/A INVX1_LOC_49/A 0.10fF
C74492 INVX1_LOC_64/A INVX1_LOC_182/A 0.09fF
C74493 INVX1_LOC_69/Y NOR2X1_LOC_383/B 0.03fF
C74494 INVX1_LOC_176/A INVX1_LOC_15/A 0.03fF
C74495 INVX1_LOC_24/A INVX1_LOC_275/A 0.07fF
C74496 NOR2X1_LOC_142/Y INVX1_LOC_130/Y 0.05fF
C74497 INVX1_LOC_35/A D_INPUT_4 0.01fF
C74498 NOR2X1_LOC_788/a_36_216# NOR2X1_LOC_383/B 0.00fF
C74499 INVX1_LOC_49/A NOR2X1_LOC_303/Y 0.60fF
C74500 INVX1_LOC_93/A INPUT_1 0.08fF
C74501 NAND2X1_LOC_579/A INVX1_LOC_229/Y 0.14fF
C74502 D_INPUT_0 NAND2X1_LOC_473/A 0.03fF
C74503 NOR2X1_LOC_590/A NAND2X1_LOC_165/a_36_24# 0.01fF
C74504 NAND2X1_LOC_783/A NAND2X1_LOC_780/Y 0.01fF
C74505 NOR2X1_LOC_716/B INVX1_LOC_71/A 0.12fF
C74506 NAND2X1_LOC_483/Y INVX1_LOC_24/A 0.03fF
C74507 INVX1_LOC_76/A NOR2X1_LOC_38/B 0.10fF
C74508 NAND2X1_LOC_54/a_36_24# INVX1_LOC_31/A 0.00fF
C74509 NOR2X1_LOC_666/Y INVX1_LOC_10/A 0.02fF
C74510 NOR2X1_LOC_441/Y NAND2X1_LOC_850/Y 0.10fF
C74511 NAND2X1_LOC_725/B NOR2X1_LOC_299/Y 0.03fF
C74512 INVX1_LOC_135/A NAND2X1_LOC_326/A 0.10fF
C74513 INVX1_LOC_224/Y NOR2X1_LOC_392/a_36_216# 0.00fF
C74514 NOR2X1_LOC_721/B INVX1_LOC_46/Y 0.04fF
C74515 NAND2X1_LOC_391/Y INVX1_LOC_28/A 0.07fF
C74516 D_INPUT_0 NAND2X1_LOC_537/Y 0.06fF
C74517 NAND2X1_LOC_303/Y NAND2X1_LOC_303/B 0.19fF
C74518 NOR2X1_LOC_790/B NOR2X1_LOC_552/Y 0.04fF
C74519 INVX1_LOC_77/A INVX1_LOC_63/Y 0.07fF
C74520 INVX1_LOC_36/A NOR2X1_LOC_191/A 0.06fF
C74521 INVX1_LOC_39/A NOR2X1_LOC_19/B 0.00fF
C74522 INVX1_LOC_49/A NOR2X1_LOC_254/Y 0.11fF
C74523 NOR2X1_LOC_629/Y INVX1_LOC_284/A 0.03fF
C74524 NOR2X1_LOC_746/a_36_216# INVX1_LOC_23/A 0.00fF
C74525 D_INPUT_1 NOR2X1_LOC_318/B 0.07fF
C74526 NOR2X1_LOC_267/A NOR2X1_LOC_191/A 0.08fF
C74527 NOR2X1_LOC_643/Y NOR2X1_LOC_6/B 0.02fF
C74528 NOR2X1_LOC_78/B NOR2X1_LOC_733/a_36_216# 0.00fF
C74529 INVX1_LOC_24/A NOR2X1_LOC_168/B 0.89fF
C74530 INVX1_LOC_303/A INVX1_LOC_104/A 0.18fF
C74531 NOR2X1_LOC_673/A NOR2X1_LOC_814/A 0.42fF
C74532 NOR2X1_LOC_498/a_36_216# NOR2X1_LOC_498/Y 0.01fF
C74533 NOR2X1_LOC_389/A NOR2X1_LOC_561/Y 0.10fF
C74534 D_INPUT_0 NOR2X1_LOC_530/a_36_216# 0.00fF
C74535 INVX1_LOC_46/A NOR2X1_LOC_89/Y 0.37fF
C74536 INVX1_LOC_12/A NOR2X1_LOC_510/B 0.05fF
C74537 NOR2X1_LOC_211/Y INVX1_LOC_286/A 0.03fF
C74538 NOR2X1_LOC_574/a_36_216# NOR2X1_LOC_152/Y 0.00fF
C74539 D_INPUT_1 INVX1_LOC_93/Y 0.07fF
C74540 NAND2X1_LOC_778/Y INPUT_0 0.10fF
C74541 NOR2X1_LOC_160/B INVX1_LOC_83/A 0.16fF
C74542 INVX1_LOC_2/A NOR2X1_LOC_303/Y 0.09fF
C74543 INVX1_LOC_77/A NOR2X1_LOC_175/A 0.07fF
C74544 NOR2X1_LOC_454/Y INVX1_LOC_302/Y 0.07fF
C74545 NOR2X1_LOC_91/A NOR2X1_LOC_305/Y 0.08fF
C74546 INVX1_LOC_95/Y INVX1_LOC_23/A 0.01fF
C74547 NOR2X1_LOC_374/A INVX1_LOC_177/A 0.02fF
C74548 INVX1_LOC_209/Y NOR2X1_LOC_504/Y 0.01fF
C74549 NAND2X1_LOC_783/A INVX1_LOC_141/Y 1.08fF
C74550 INVX1_LOC_49/A NOR2X1_LOC_353/Y 0.01fF
C74551 NOR2X1_LOC_718/Y INVX1_LOC_266/Y 0.01fF
C74552 NOR2X1_LOC_360/Y INVX1_LOC_232/A 0.12fF
C74553 INVX1_LOC_217/Y NOR2X1_LOC_52/B -0.01fF
C74554 NOR2X1_LOC_457/B INVX1_LOC_22/A 0.07fF
C74555 NOR2X1_LOC_759/Y INVX1_LOC_52/A 0.01fF
C74556 INVX1_LOC_50/A NOR2X1_LOC_357/Y 0.15fF
C74557 NAND2X1_LOC_783/A INVX1_LOC_312/Y 0.10fF
C74558 NOR2X1_LOC_391/A INVX1_LOC_72/A 0.02fF
C74559 INVX1_LOC_58/A NAND2X1_LOC_244/A 0.03fF
C74560 INVX1_LOC_45/A NOR2X1_LOC_717/B 0.03fF
C74561 INVX1_LOC_34/A INVX1_LOC_96/Y 0.29fF
C74562 INVX1_LOC_64/A INVX1_LOC_291/Y 0.07fF
C74563 INVX1_LOC_123/Y INVX1_LOC_42/A 0.11fF
C74564 INVX1_LOC_47/A INVX1_LOC_31/A 0.03fF
C74565 NOR2X1_LOC_644/B INVX1_LOC_313/Y 0.00fF
C74566 NOR2X1_LOC_15/Y INPUT_0 0.22fF
C74567 NOR2X1_LOC_516/B INVX1_LOC_184/A 0.08fF
C74568 NOR2X1_LOC_599/A NAND2X1_LOC_809/A 0.02fF
C74569 NOR2X1_LOC_32/B NOR2X1_LOC_670/Y 0.01fF
C74570 NOR2X1_LOC_89/A NOR2X1_LOC_127/Y 0.27fF
C74571 INVX1_LOC_24/A NOR2X1_LOC_789/A 0.00fF
C74572 NOR2X1_LOC_68/A NOR2X1_LOC_171/a_36_216# 0.01fF
C74573 INVX1_LOC_286/A NOR2X1_LOC_440/B 0.22fF
C74574 NOR2X1_LOC_615/a_36_216# NAND2X1_LOC_560/A 0.00fF
C74575 NAND2X1_LOC_562/Y NAND2X1_LOC_570/Y 0.02fF
C74576 NOR2X1_LOC_408/a_36_216# D_INPUT_4 0.00fF
C74577 INVX1_LOC_234/A INVX1_LOC_61/A 0.05fF
C74578 NOR2X1_LOC_78/B NOR2X1_LOC_317/B 0.05fF
C74579 NOR2X1_LOC_468/Y NOR2X1_LOC_167/Y 0.35fF
C74580 NOR2X1_LOC_238/Y NAND2X1_LOC_859/Y 0.53fF
C74581 INVX1_LOC_53/A NAND2X1_LOC_211/Y 0.07fF
C74582 INVX1_LOC_41/A NOR2X1_LOC_544/A 0.07fF
C74583 NOR2X1_LOC_536/A NAND2X1_LOC_288/B 0.02fF
C74584 NAND2X1_LOC_860/A NOR2X1_LOC_266/B 0.05fF
C74585 NOR2X1_LOC_750/Y VDD 0.43fF
C74586 NOR2X1_LOC_501/a_36_216# INVX1_LOC_71/A 0.00fF
C74587 INVX1_LOC_93/Y NOR2X1_LOC_652/Y 0.75fF
C74588 NAND2X1_LOC_633/Y NAND2X1_LOC_793/B 0.51fF
C74589 NAND2X1_LOC_149/Y INVX1_LOC_91/A 0.07fF
C74590 NOR2X1_LOC_773/Y INVX1_LOC_162/Y 0.07fF
C74591 NOR2X1_LOC_203/Y INVX1_LOC_104/A 0.09fF
C74592 NOR2X1_LOC_82/Y NAND2X1_LOC_494/a_36_24# 0.00fF
C74593 INVX1_LOC_50/A NOR2X1_LOC_692/Y 0.02fF
C74594 NOR2X1_LOC_299/Y INVX1_LOC_309/Y 0.01fF
C74595 NOR2X1_LOC_401/Y NOR2X1_LOC_84/Y 0.03fF
C74596 INVX1_LOC_2/A INVX1_LOC_54/Y 0.01fF
C74597 NAND2X1_LOC_9/Y INVX1_LOC_12/Y 0.03fF
C74598 INVX1_LOC_110/Y NAND2X1_LOC_348/A 0.41fF
C74599 NOR2X1_LOC_717/B INVX1_LOC_71/A 0.03fF
C74600 NOR2X1_LOC_285/Y VDD 0.24fF
C74601 NAND2X1_LOC_472/Y NOR2X1_LOC_717/A 0.03fF
C74602 INVX1_LOC_233/A INVX1_LOC_12/Y 0.18fF
C74603 NOR2X1_LOC_226/A INVX1_LOC_54/Y 0.17fF
C74604 NOR2X1_LOC_68/A NOR2X1_LOC_356/A 0.10fF
C74605 INVX1_LOC_27/A NAND2X1_LOC_212/Y 0.02fF
C74606 NOR2X1_LOC_448/a_36_216# INVX1_LOC_91/A 0.00fF
C74607 NAND2X1_LOC_860/A NAND2X1_LOC_848/A 0.03fF
C74608 NAND2X1_LOC_214/B D_INPUT_3 0.03fF
C74609 NOR2X1_LOC_82/A INVX1_LOC_123/A 0.01fF
C74610 INVX1_LOC_204/Y VDD 0.21fF
C74611 INVX1_LOC_273/Y NOR2X1_LOC_577/Y 0.03fF
C74612 INVX1_LOC_45/A NOR2X1_LOC_151/Y 0.24fF
C74613 NOR2X1_LOC_238/Y NAND2X1_LOC_866/B 0.02fF
C74614 INVX1_LOC_239/A NAND2X1_LOC_659/B 0.14fF
C74615 NOR2X1_LOC_206/a_36_216# NOR2X1_LOC_357/Y 0.01fF
C74616 NOR2X1_LOC_92/Y NAND2X1_LOC_468/B 0.03fF
C74617 NOR2X1_LOC_172/Y NOR2X1_LOC_60/a_36_216# 0.00fF
C74618 INVX1_LOC_243/Y NAND2X1_LOC_428/a_36_24# 0.01fF
C74619 INVX1_LOC_280/Y NAND2X1_LOC_852/Y 0.08fF
C74620 NOR2X1_LOC_361/B NAND2X1_LOC_642/Y 0.07fF
C74621 NOR2X1_LOC_716/B NOR2X1_LOC_123/B 0.01fF
C74622 NAND2X1_LOC_553/A INVX1_LOC_12/Y 0.16fF
C74623 INVX1_LOC_240/A NOR2X1_LOC_32/Y 0.01fF
C74624 NOR2X1_LOC_322/Y INVX1_LOC_18/A 0.07fF
C74625 INVX1_LOC_225/A NAND2X1_LOC_573/A 0.01fF
C74626 INVX1_LOC_27/A D_INPUT_3 0.19fF
C74627 NOR2X1_LOC_605/B NAND2X1_LOC_722/A 0.28fF
C74628 INVX1_LOC_27/A INVX1_LOC_14/Y 0.10fF
C74629 INVX1_LOC_102/A INVX1_LOC_42/A 0.07fF
C74630 NOR2X1_LOC_598/B NOR2X1_LOC_729/A 0.10fF
C74631 INVX1_LOC_83/A NOR2X1_LOC_317/B 0.03fF
C74632 NOR2X1_LOC_716/B NOR2X1_LOC_749/Y 0.07fF
C74633 NOR2X1_LOC_78/B NOR2X1_LOC_516/B 0.03fF
C74634 INVX1_LOC_14/A INVX1_LOC_74/A 0.02fF
C74635 NAND2X1_LOC_579/A INVX1_LOC_20/A 0.10fF
C74636 D_INPUT_0 NOR2X1_LOC_516/Y 0.01fF
C74637 NAND2X1_LOC_787/A NOR2X1_LOC_177/a_36_216# 0.00fF
C74638 NAND2X1_LOC_181/Y INVX1_LOC_25/Y 0.06fF
C74639 NOR2X1_LOC_468/Y INVX1_LOC_76/A 0.07fF
C74640 NOR2X1_LOC_340/A INVX1_LOC_15/A 0.05fF
C74641 INVX1_LOC_223/Y INVX1_LOC_117/A 0.01fF
C74642 NOR2X1_LOC_68/A NOR2X1_LOC_74/A 2.63fF
C74643 NAND2X1_LOC_521/a_36_24# NAND2X1_LOC_348/A 0.01fF
C74644 INVX1_LOC_57/A NOR2X1_LOC_445/B 0.03fF
C74645 NOR2X1_LOC_151/Y INVX1_LOC_71/A 0.03fF
C74646 INVX1_LOC_135/A NOR2X1_LOC_87/B 0.08fF
C74647 NOR2X1_LOC_722/Y NOR2X1_LOC_733/Y 0.01fF
C74648 NOR2X1_LOC_391/A NAND2X1_LOC_338/B 0.07fF
C74649 NOR2X1_LOC_84/A INPUT_1 0.01fF
C74650 INVX1_LOC_295/A NAND2X1_LOC_163/a_36_24# 0.01fF
C74651 NOR2X1_LOC_68/A NOR2X1_LOC_9/Y 0.12fF
C74652 INVX1_LOC_71/Y NAND2X1_LOC_793/B 0.01fF
C74653 NAND2X1_LOC_860/A INVX1_LOC_46/Y 0.44fF
C74654 NOR2X1_LOC_318/A INVX1_LOC_63/A 0.07fF
C74655 INVX1_LOC_77/A INVX1_LOC_302/Y 0.04fF
C74656 NOR2X1_LOC_447/Y NAND2X1_LOC_51/B 0.00fF
C74657 INVX1_LOC_172/A NOR2X1_LOC_322/Y 0.30fF
C74658 INVX1_LOC_241/A NAND2X1_LOC_579/a_36_24# 0.02fF
C74659 INVX1_LOC_73/A NOR2X1_LOC_577/Y 0.07fF
C74660 INVX1_LOC_94/Y NAND2X1_LOC_74/B 0.05fF
C74661 INVX1_LOC_83/A INVX1_LOC_189/A 0.01fF
C74662 NAND2X1_LOC_738/B INVX1_LOC_297/A 0.03fF
C74663 INVX1_LOC_27/A INVX1_LOC_230/A 0.07fF
C74664 NAND2X1_LOC_538/Y INVX1_LOC_37/A 0.09fF
C74665 NOR2X1_LOC_860/B INPUT_0 0.21fF
C74666 INVX1_LOC_73/Y VDD -0.00fF
C74667 NOR2X1_LOC_180/B NOR2X1_LOC_348/B 0.09fF
C74668 NAND2X1_LOC_321/a_36_24# NOR2X1_LOC_324/A 0.02fF
C74669 INVX1_LOC_208/Y NOR2X1_LOC_589/A 0.03fF
C74670 INVX1_LOC_93/A INVX1_LOC_118/A 0.07fF
C74671 NAND2X1_LOC_712/A INVX1_LOC_16/A 0.02fF
C74672 NAND2X1_LOC_326/A NOR2X1_LOC_152/A 0.01fF
C74673 INVX1_LOC_31/A INVX1_LOC_95/Y 0.07fF
C74674 NAND2X1_LOC_562/Y NOR2X1_LOC_19/B 0.44fF
C74675 NAND2X1_LOC_349/B NAND2X1_LOC_514/a_36_24# 0.00fF
C74676 NOR2X1_LOC_384/Y NOR2X1_LOC_45/B 1.46fF
C74677 NOR2X1_LOC_781/A INVX1_LOC_22/A 0.03fF
C74678 NOR2X1_LOC_376/A NOR2X1_LOC_376/Y 0.05fF
C74679 NOR2X1_LOC_793/A NAND2X1_LOC_417/a_36_24# 0.00fF
C74680 NOR2X1_LOC_238/Y INVX1_LOC_6/A 0.01fF
C74681 INVX1_LOC_1/A INVX1_LOC_281/A 0.08fF
C74682 INVX1_LOC_286/A INVX1_LOC_41/Y 0.48fF
C74683 INVX1_LOC_24/A INVX1_LOC_78/Y 0.03fF
C74684 NOR2X1_LOC_562/B INVX1_LOC_18/A 0.39fF
C74685 INVX1_LOC_143/A INVX1_LOC_132/Y 0.63fF
C74686 NAND2X1_LOC_550/A INVX1_LOC_46/A 0.04fF
C74687 INVX1_LOC_102/A INVX1_LOC_78/A 0.07fF
C74688 NOR2X1_LOC_389/A INVX1_LOC_76/A 0.43fF
C74689 INVX1_LOC_14/A NAND2X1_LOC_699/a_36_24# 0.00fF
C74690 NOR2X1_LOC_160/B INVX1_LOC_46/A 0.10fF
C74691 INVX1_LOC_72/A INVX1_LOC_187/A 0.02fF
C74692 NAND2X1_LOC_537/Y NAND2X1_LOC_848/A 0.07fF
C74693 NAND2X1_LOC_579/a_36_24# NOR2X1_LOC_298/Y 0.06fF
C74694 INVX1_LOC_241/A NOR2X1_LOC_299/Y 0.08fF
C74695 INVX1_LOC_31/A NOR2X1_LOC_305/Y 0.07fF
C74696 NAND2X1_LOC_74/B INVX1_LOC_181/A 0.07fF
C74697 NOR2X1_LOC_516/B INVX1_LOC_83/A 5.76fF
C74698 NOR2X1_LOC_91/A NOR2X1_LOC_189/a_36_216# 0.00fF
C74699 NOR2X1_LOC_371/a_36_216# NAND2X1_LOC_721/A 0.03fF
C74700 INVX1_LOC_234/A NAND2X1_LOC_735/B 0.14fF
C74701 NOR2X1_LOC_78/B NOR2X1_LOC_756/a_36_216# 0.00fF
C74702 INVX1_LOC_45/A NOR2X1_LOC_567/a_36_216# 0.00fF
C74703 NOR2X1_LOC_678/A INVX1_LOC_63/A 0.00fF
C74704 INVX1_LOC_39/A NOR2X1_LOC_216/B 0.04fF
C74705 NOR2X1_LOC_272/Y NOR2X1_LOC_831/B 0.10fF
C74706 NOR2X1_LOC_89/A NOR2X1_LOC_383/B 0.17fF
C74707 NOR2X1_LOC_567/a_36_216# NOR2X1_LOC_568/A 0.00fF
C74708 INVX1_LOC_98/Y INVX1_LOC_102/Y 0.01fF
C74709 NOR2X1_LOC_360/Y NAND2X1_LOC_447/Y 0.10fF
C74710 NOR2X1_LOC_703/B NOR2X1_LOC_35/Y 0.01fF
C74711 INVX1_LOC_12/A INVX1_LOC_57/A 4.26fF
C74712 NOR2X1_LOC_284/B NOR2X1_LOC_567/B 0.03fF
C74713 NOR2X1_LOC_67/A NAND2X1_LOC_560/A 0.01fF
C74714 NOR2X1_LOC_180/B INVX1_LOC_22/A 3.21fF
C74715 NOR2X1_LOC_272/Y NOR2X1_LOC_179/a_36_216# 0.12fF
C74716 NOR2X1_LOC_298/Y NOR2X1_LOC_299/Y 0.48fF
C74717 INPUT_0 NAND2X1_LOC_141/A 0.03fF
C74718 INVX1_LOC_36/Y NOR2X1_LOC_554/B 0.14fF
C74719 NAND2X1_LOC_656/Y NOR2X1_LOC_130/A 0.07fF
C74720 NAND2X1_LOC_181/Y INVX1_LOC_75/A 0.03fF
C74721 INVX1_LOC_1/A NOR2X1_LOC_862/B 0.10fF
C74722 INVX1_LOC_132/A INVX1_LOC_65/A 0.02fF
C74723 INVX1_LOC_108/Y NOR2X1_LOC_340/A 0.07fF
C74724 NOR2X1_LOC_91/Y VDD 0.59fF
C74725 NAND2X1_LOC_35/Y NAND2X1_LOC_500/B 0.02fF
C74726 NOR2X1_LOC_843/A NOR2X1_LOC_78/A 0.03fF
C74727 NOR2X1_LOC_596/A INVX1_LOC_76/A 0.07fF
C74728 NAND2X1_LOC_543/Y INVX1_LOC_140/A 0.09fF
C74729 NOR2X1_LOC_19/B NAND2X1_LOC_735/B 0.03fF
C74730 NAND2X1_LOC_363/B INVX1_LOC_106/Y 0.01fF
C74731 NOR2X1_LOC_168/A INVX1_LOC_69/Y 0.01fF
C74732 INVX1_LOC_73/A INVX1_LOC_22/A 0.42fF
C74733 INVX1_LOC_50/A INVX1_LOC_32/A 0.06fF
C74734 NOR2X1_LOC_359/Y VDD 0.15fF
C74735 INPUT_0 INVX1_LOC_226/A 0.06fF
C74736 INVX1_LOC_50/Y INVX1_LOC_19/A 0.22fF
C74737 INVX1_LOC_103/A NOR2X1_LOC_88/Y 0.00fF
C74738 INVX1_LOC_235/Y INVX1_LOC_203/A 0.02fF
C74739 NOR2X1_LOC_590/A NOR2X1_LOC_612/Y 0.00fF
C74740 NAND2X1_LOC_633/Y INVX1_LOC_71/A 0.16fF
C74741 INVX1_LOC_249/A INVX1_LOC_14/Y 0.34fF
C74742 NOR2X1_LOC_203/Y INVX1_LOC_206/Y 0.05fF
C74743 INVX1_LOC_244/Y INVX1_LOC_77/Y 0.02fF
C74744 NAND2X1_LOC_349/B NAND2X1_LOC_138/a_36_24# 0.00fF
C74745 NOR2X1_LOC_570/Y NOR2X1_LOC_74/A 0.38fF
C74746 INVX1_LOC_45/A NOR2X1_LOC_209/B 0.15fF
C74747 NOR2X1_LOC_392/Y INVX1_LOC_3/Y 0.17fF
C74748 NOR2X1_LOC_216/Y NAND2X1_LOC_656/Y 0.07fF
C74749 INVX1_LOC_26/A INVX1_LOC_23/Y 0.34fF
C74750 NOR2X1_LOC_495/Y NAND2X1_LOC_804/Y 0.01fF
C74751 INVX1_LOC_103/A INVX1_LOC_84/A 0.07fF
C74752 INVX1_LOC_45/Y NOR2X1_LOC_536/A 0.00fF
C74753 NOR2X1_LOC_134/Y INVX1_LOC_35/Y 0.04fF
C74754 INVX1_LOC_268/A INVX1_LOC_6/A 0.01fF
C74755 NAND2X1_LOC_477/A NAND2X1_LOC_468/B 0.12fF
C74756 INVX1_LOC_83/A NOR2X1_LOC_706/A 0.08fF
C74757 INVX1_LOC_266/Y INVX1_LOC_188/Y 0.32fF
C74758 INPUT_6 NAND2X1_LOC_3/B 0.32fF
C74759 INVX1_LOC_50/A NAND2X1_LOC_175/Y 0.16fF
C74760 INVX1_LOC_266/A INVX1_LOC_19/A 0.01fF
C74761 NAND2X1_LOC_72/Y INVX1_LOC_32/A 0.19fF
C74762 INVX1_LOC_23/A INVX1_LOC_271/Y 0.10fF
C74763 NAND2X1_LOC_717/Y INVX1_LOC_11/Y 0.15fF
C74764 NAND2X1_LOC_736/B VDD 0.17fF
C74765 NOR2X1_LOC_602/a_36_216# NOR2X1_LOC_743/Y 0.00fF
C74766 INVX1_LOC_200/A NOR2X1_LOC_662/A 0.02fF
C74767 INVX1_LOC_191/Y INVX1_LOC_187/Y 0.01fF
C74768 INVX1_LOC_135/A NOR2X1_LOC_527/Y 0.06fF
C74769 INVX1_LOC_229/Y NOR2X1_LOC_387/A 0.06fF
C74770 INVX1_LOC_16/A INVX1_LOC_91/A 5.16fF
C74771 INVX1_LOC_292/A INVX1_LOC_84/A 0.07fF
C74772 INVX1_LOC_299/A NAND2X1_LOC_74/B 0.10fF
C74773 INVX1_LOC_30/Y INVX1_LOC_125/Y 0.01fF
C74774 INVX1_LOC_41/Y INVX1_LOC_54/A 0.05fF
C74775 NAND2X1_LOC_357/B NOR2X1_LOC_111/A 0.03fF
C74776 D_INPUT_0 NOR2X1_LOC_86/a_36_216# 0.00fF
C74777 NOR2X1_LOC_51/a_36_216# INPUT_5 0.00fF
C74778 NAND2X1_LOC_729/B INVX1_LOC_22/A 0.00fF
C74779 NOR2X1_LOC_538/B NAND2X1_LOC_74/B 0.43fF
C74780 INVX1_LOC_206/A INVX1_LOC_14/Y 0.34fF
C74781 NAND2X1_LOC_505/a_36_24# NOR2X1_LOC_349/A 0.02fF
C74782 NAND2X1_LOC_364/A NOR2X1_LOC_831/B 0.36fF
C74783 INVX1_LOC_100/A NOR2X1_LOC_76/A 0.10fF
C74784 INVX1_LOC_16/A INVX1_LOC_11/Y 0.03fF
C74785 INVX1_LOC_123/A INVX1_LOC_306/A 0.02fF
C74786 NOR2X1_LOC_131/a_36_216# NAND2X1_LOC_469/B 0.00fF
C74787 NAND2X1_LOC_593/Y INVX1_LOC_54/A 0.08fF
C74788 NOR2X1_LOC_232/Y INVX1_LOC_284/A 0.03fF
C74789 INVX1_LOC_14/A NAND2X1_LOC_254/Y 0.03fF
C74790 NOR2X1_LOC_220/A INVX1_LOC_76/A 0.10fF
C74791 NOR2X1_LOC_78/B NAND2X1_LOC_211/Y 0.01fF
C74792 INVX1_LOC_286/Y NOR2X1_LOC_661/a_36_216# 0.00fF
C74793 NOR2X1_LOC_363/a_36_216# INVX1_LOC_92/A 0.00fF
C74794 INVX1_LOC_83/A INVX1_LOC_315/Y 0.10fF
C74795 NOR2X1_LOC_468/Y INVX1_LOC_127/Y 0.01fF
C74796 NOR2X1_LOC_68/A NOR2X1_LOC_243/B 0.53fF
C74797 NOR2X1_LOC_366/Y NOR2X1_LOC_269/Y 0.01fF
C74798 NAND2X1_LOC_573/A NAND2X1_LOC_642/Y 0.02fF
C74799 INVX1_LOC_87/A NOR2X1_LOC_652/Y 0.03fF
C74800 NAND2X1_LOC_853/Y INVX1_LOC_46/A 1.04fF
C74801 NOR2X1_LOC_87/B INVX1_LOC_280/A 0.02fF
C74802 NAND2X1_LOC_850/Y NOR2X1_LOC_176/Y 0.29fF
C74803 INVX1_LOC_305/A INVX1_LOC_63/A 0.12fF
C74804 NOR2X1_LOC_561/Y NAND2X1_LOC_469/B 0.32fF
C74805 NAND2X1_LOC_741/B NOR2X1_LOC_36/B 0.08fF
C74806 INVX1_LOC_58/A NOR2X1_LOC_392/Y 0.00fF
C74807 INVX1_LOC_170/A NAND2X1_LOC_81/B 0.18fF
C74808 INVX1_LOC_103/A INVX1_LOC_15/A 0.11fF
C74809 NOR2X1_LOC_175/A INVX1_LOC_9/A 0.07fF
C74810 INVX1_LOC_50/Y INVX1_LOC_26/Y 0.09fF
C74811 NAND2X1_LOC_101/a_36_24# INVX1_LOC_27/Y 0.00fF
C74812 NOR2X1_LOC_264/Y INVX1_LOC_92/A 0.05fF
C74813 NAND2X1_LOC_853/Y NOR2X1_LOC_766/Y 0.03fF
C74814 NOR2X1_LOC_278/A NOR2X1_LOC_118/a_36_216# 0.00fF
C74815 INVX1_LOC_33/A INVX1_LOC_113/A 0.08fF
C74816 INVX1_LOC_28/A INVX1_LOC_91/A 0.18fF
C74817 NOR2X1_LOC_543/A VDD -0.00fF
C74818 INVX1_LOC_17/A NAND2X1_LOC_647/B 0.02fF
C74819 INVX1_LOC_77/A INVX1_LOC_27/Y 0.03fF
C74820 INVX1_LOC_209/Y NOR2X1_LOC_697/Y 0.75fF
C74821 NOR2X1_LOC_542/Y NOR2X1_LOC_542/B 0.15fF
C74822 INVX1_LOC_30/A NOR2X1_LOC_12/a_36_216# 0.00fF
C74823 NOR2X1_LOC_757/Y NOR2X1_LOC_331/B 0.02fF
C74824 NOR2X1_LOC_433/A NOR2X1_LOC_127/Y 0.05fF
C74825 INVX1_LOC_186/A NOR2X1_LOC_567/B 0.07fF
C74826 NOR2X1_LOC_561/Y NOR2X1_LOC_447/B 0.01fF
C74827 INVX1_LOC_57/Y NOR2X1_LOC_89/A 0.15fF
C74828 INVX1_LOC_181/A NAND2X1_LOC_793/a_36_24# 0.00fF
C74829 NOR2X1_LOC_598/B INVX1_LOC_68/A 0.01fF
C74830 NOR2X1_LOC_476/B INVX1_LOC_253/Y 0.01fF
C74831 INVX1_LOC_201/Y NAND2X1_LOC_141/Y 0.36fF
C74832 NOR2X1_LOC_91/A INVX1_LOC_59/A 0.00fF
C74833 INVX1_LOC_223/A INVX1_LOC_42/A 0.07fF
C74834 INVX1_LOC_28/A INVX1_LOC_11/Y 3.01fF
C74835 INVX1_LOC_61/Y INVX1_LOC_32/A 0.07fF
C74836 NOR2X1_LOC_15/Y INVX1_LOC_183/A 0.01fF
C74837 NAND2X1_LOC_164/a_36_24# NOR2X1_LOC_445/B 0.00fF
C74838 INVX1_LOC_59/A INVX1_LOC_23/A 0.04fF
C74839 NOR2X1_LOC_52/B NOR2X1_LOC_127/Y 0.07fF
C74840 NOR2X1_LOC_275/a_36_216# NAND2X1_LOC_454/Y 0.01fF
C74841 NAND2X1_LOC_347/B INVX1_LOC_29/Y 0.01fF
C74842 INVX1_LOC_255/Y NOR2X1_LOC_655/Y 0.04fF
C74843 NOR2X1_LOC_32/B INVX1_LOC_258/Y 0.30fF
C74844 NOR2X1_LOC_71/Y NOR2X1_LOC_536/A 0.07fF
C74845 INVX1_LOC_41/Y NOR2X1_LOC_48/B 0.01fF
C74846 NOR2X1_LOC_19/B D_INPUT_3 4.23fF
C74847 NOR2X1_LOC_717/B NOR2X1_LOC_331/B 0.05fF
C74848 NAND2X1_LOC_842/B INVX1_LOC_12/Y 0.01fF
C74849 INVX1_LOC_11/A NOR2X1_LOC_383/B 0.06fF
C74850 NAND2X1_LOC_214/Y NOR2X1_LOC_598/B 0.03fF
C74851 NOR2X1_LOC_456/Y NOR2X1_LOC_464/B 0.01fF
C74852 NOR2X1_LOC_4/a_36_216# NAND2X1_LOC_82/Y 0.00fF
C74853 NOR2X1_LOC_6/B INVX1_LOC_19/A 0.14fF
C74854 INVX1_LOC_186/A NAND2X1_LOC_677/a_36_24# 0.01fF
C74855 INVX1_LOC_200/A INVX1_LOC_57/A 3.76fF
C74856 NAND2X1_LOC_593/Y NOR2X1_LOC_48/B 0.06fF
C74857 INVX1_LOC_95/Y INVX1_LOC_6/A 0.10fF
C74858 INVX1_LOC_223/A INVX1_LOC_78/A 0.06fF
C74859 INVX1_LOC_225/A NAND2X1_LOC_81/B 0.03fF
C74860 NOR2X1_LOC_67/A NOR2X1_LOC_673/B 0.05fF
C74861 NOR2X1_LOC_455/Y NAND2X1_LOC_190/Y 0.02fF
C74862 INVX1_LOC_136/A INVX1_LOC_94/Y 0.11fF
C74863 INVX1_LOC_64/A NAND2X1_LOC_579/A 0.07fF
C74864 D_INPUT_1 NOR2X1_LOC_82/A 0.82fF
C74865 NOR2X1_LOC_454/Y INVX1_LOC_5/A 0.14fF
C74866 NOR2X1_LOC_45/B NOR2X1_LOC_43/Y 0.46fF
C74867 NAND2X1_LOC_584/a_36_24# NAND2X1_LOC_651/B 0.00fF
C74868 INVX1_LOC_64/A NOR2X1_LOC_187/Y 0.05fF
C74869 NOR2X1_LOC_191/A INVX1_LOC_63/A 0.03fF
C74870 NOR2X1_LOC_387/A INVX1_LOC_20/A 0.06fF
C74871 NOR2X1_LOC_315/Y NAND2X1_LOC_74/B 2.79fF
C74872 NAND2X1_LOC_35/Y NAND2X1_LOC_725/B 0.08fF
C74873 INVX1_LOC_233/A NOR2X1_LOC_401/A 0.03fF
C74874 NOR2X1_LOC_178/Y NOR2X1_LOC_468/Y 0.15fF
C74875 INVX1_LOC_123/A INVX1_LOC_59/Y 0.17fF
C74876 INVX1_LOC_246/A NAND2X1_LOC_678/a_36_24# 0.00fF
C74877 INVX1_LOC_75/A INVX1_LOC_117/A 0.23fF
C74878 INVX1_LOC_54/Y NAND2X1_LOC_63/Y 0.00fF
C74879 NOR2X1_LOC_71/Y NAND2X1_LOC_93/B 0.01fF
C74880 NOR2X1_LOC_92/Y INVX1_LOC_13/Y 0.72fF
C74881 INVX1_LOC_269/A NOR2X1_LOC_663/A 0.02fF
C74882 INVX1_LOC_255/Y NOR2X1_LOC_649/B 0.04fF
C74883 INVX1_LOC_30/A NOR2X1_LOC_635/B 0.06fF
C74884 INVX1_LOC_255/Y INVX1_LOC_3/A 0.19fF
C74885 NOR2X1_LOC_65/B INVX1_LOC_223/A 0.02fF
C74886 INVX1_LOC_256/A NOR2X1_LOC_405/Y 0.03fF
C74887 NAND2X1_LOC_9/Y NOR2X1_LOC_160/B 0.06fF
C74888 NAND2X1_LOC_860/A NOR2X1_LOC_134/Y 0.02fF
C74889 INVX1_LOC_21/A NOR2X1_LOC_227/B 0.02fF
C74890 NAND2X1_LOC_391/Y INVX1_LOC_48/Y 0.01fF
C74891 NOR2X1_LOC_223/B INVX1_LOC_103/A 0.03fF
C74892 NOR2X1_LOC_135/Y INVX1_LOC_118/Y 0.17fF
C74893 INVX1_LOC_91/A NOR2X1_LOC_253/Y 0.05fF
C74894 INVX1_LOC_16/A INVX1_LOC_203/A 0.07fF
C74895 INVX1_LOC_30/A INVX1_LOC_275/Y 0.00fF
C74896 NOR2X1_LOC_67/A INVX1_LOC_29/A 0.12fF
C74897 INVX1_LOC_269/A NOR2X1_LOC_674/Y 0.04fF
C74898 NOR2X1_LOC_824/A NAND2X1_LOC_705/Y 0.06fF
C74899 INVX1_LOC_30/A NOR2X1_LOC_748/A 0.07fF
C74900 INVX1_LOC_91/A NOR2X1_LOC_35/Y 0.10fF
C74901 INVX1_LOC_132/A INVX1_LOC_4/Y 0.10fF
C74902 NOR2X1_LOC_151/Y NOR2X1_LOC_331/B 0.03fF
C74903 INVX1_LOC_233/A NOR2X1_LOC_160/B 0.10fF
C74904 NOR2X1_LOC_481/A INVX1_LOC_4/Y 0.03fF
C74905 INVX1_LOC_41/Y NOR2X1_LOC_438/Y 0.00fF
C74906 NOR2X1_LOC_303/Y NOR2X1_LOC_631/Y 0.14fF
C74907 INPUT_1 INVX1_LOC_35/Y 0.07fF
C74908 INVX1_LOC_217/A INVX1_LOC_57/A 0.07fF
C74909 NOR2X1_LOC_334/A NAND2X1_LOC_96/A 0.27fF
C74910 INVX1_LOC_52/Y NAND2X1_LOC_67/Y 0.13fF
C74911 NAND2X1_LOC_563/A INVX1_LOC_284/A 0.01fF
C74912 INVX1_LOC_30/Y INVX1_LOC_19/A 0.03fF
C74913 NAND2X1_LOC_553/A NOR2X1_LOC_160/B 0.01fF
C74914 INVX1_LOC_225/A INVX1_LOC_4/Y 0.07fF
C74915 NAND2X1_LOC_170/A NOR2X1_LOC_89/A 0.03fF
C74916 NAND2X1_LOC_11/Y NAND2X1_LOC_430/B 0.06fF
C74917 NOR2X1_LOC_92/Y INVX1_LOC_88/A 0.14fF
C74918 NOR2X1_LOC_828/B NAND2X1_LOC_425/Y 0.01fF
C74919 D_INPUT_1 NAND2X1_LOC_153/a_36_24# 0.01fF
C74920 NOR2X1_LOC_798/A NOR2X1_LOC_160/B 0.05fF
C74921 NAND2X1_LOC_469/B INVX1_LOC_76/A 0.03fF
C74922 NOR2X1_LOC_272/Y NAND2X1_LOC_352/B 0.02fF
C74923 INVX1_LOC_135/A NAND2X1_LOC_219/B 0.03fF
C74924 NOR2X1_LOC_598/a_36_216# INVX1_LOC_53/A 0.00fF
C74925 NAND2X1_LOC_543/Y INVX1_LOC_42/A 0.03fF
C74926 INVX1_LOC_20/Y NOR2X1_LOC_814/A 0.05fF
C74927 INVX1_LOC_85/A INVX1_LOC_78/A 0.03fF
C74928 INVX1_LOC_86/A INVX1_LOC_92/A 0.03fF
C74929 NOR2X1_LOC_593/Y NOR2X1_LOC_383/B 0.03fF
C74930 NOR2X1_LOC_422/Y NAND2X1_LOC_453/A 0.08fF
C74931 NOR2X1_LOC_272/Y INVX1_LOC_81/Y 0.10fF
C74932 NOR2X1_LOC_724/a_36_216# NOR2X1_LOC_334/Y 0.01fF
C74933 INVX1_LOC_286/A INVX1_LOC_185/A 0.92fF
C74934 NOR2X1_LOC_808/A NOR2X1_LOC_334/Y 0.03fF
C74935 NOR2X1_LOC_314/Y NAND2X1_LOC_453/A 0.01fF
C74936 INVX1_LOC_25/Y INVX1_LOC_3/Y 0.11fF
C74937 INVX1_LOC_83/A NAND2X1_LOC_207/B 0.01fF
C74938 INVX1_LOC_76/A NAND2X1_LOC_212/a_36_24# 0.01fF
C74939 INVX1_LOC_46/A NAND2X1_LOC_211/Y 0.12fF
C74940 INVX1_LOC_28/A INVX1_LOC_203/A 0.07fF
C74941 INVX1_LOC_59/A INVX1_LOC_31/A 0.03fF
C74942 NOR2X1_LOC_6/B INVX1_LOC_26/Y 0.14fF
C74943 INVX1_LOC_16/A INVX1_LOC_231/A 0.03fF
C74944 NOR2X1_LOC_637/B INVX1_LOC_53/A 0.02fF
C74945 NOR2X1_LOC_278/A INVX1_LOC_181/A 0.01fF
C74946 INVX1_LOC_166/A NOR2X1_LOC_6/B 0.04fF
C74947 NOR2X1_LOC_240/Y NOR2X1_LOC_860/B 0.10fF
C74948 INVX1_LOC_155/A INVX1_LOC_53/A 0.01fF
C74949 NAND2X1_LOC_153/a_36_24# NOR2X1_LOC_652/Y 0.00fF
C74950 INVX1_LOC_78/Y NOR2X1_LOC_197/B 0.03fF
C74951 INVX1_LOC_50/A NAND2X1_LOC_147/a_36_24# 0.00fF
C74952 NOR2X1_LOC_557/Y NOR2X1_LOC_717/A 0.56fF
C74953 INVX1_LOC_304/Y INVX1_LOC_57/A 0.07fF
C74954 INVX1_LOC_24/Y NOR2X1_LOC_500/B 0.33fF
C74955 INVX1_LOC_58/A NAND2X1_LOC_734/B 0.01fF
C74956 NOR2X1_LOC_468/a_36_216# INVX1_LOC_47/Y 0.01fF
C74957 INVX1_LOC_5/A INVX1_LOC_77/A 0.21fF
C74958 INVX1_LOC_299/A INVX1_LOC_136/A 0.10fF
C74959 INVX1_LOC_269/A INVX1_LOC_72/A 1.49fF
C74960 NOR2X1_LOC_113/A NOR2X1_LOC_831/B 0.01fF
C74961 INVX1_LOC_41/A NOR2X1_LOC_772/B 0.01fF
C74962 INVX1_LOC_232/A INVX1_LOC_26/A 0.03fF
C74963 INVX1_LOC_27/A NOR2X1_LOC_106/Y 0.03fF
C74964 INVX1_LOC_120/A INVX1_LOC_15/A 0.08fF
C74965 NOR2X1_LOC_778/Y NOR2X1_LOC_784/Y 0.08fF
C74966 NOR2X1_LOC_405/A NOR2X1_LOC_831/B 0.07fF
C74967 NAND2X1_LOC_316/a_36_24# NOR2X1_LOC_652/Y 0.00fF
C74968 NOR2X1_LOC_155/A NOR2X1_LOC_833/Y 0.07fF
C74969 NAND2X1_LOC_773/Y INVX1_LOC_111/A 0.06fF
C74970 INVX1_LOC_41/A INVX1_LOC_13/Y 0.06fF
C74971 NOR2X1_LOC_340/Y NOR2X1_LOC_849/A 0.02fF
C74972 INVX1_LOC_21/A NAND2X1_LOC_361/Y 0.07fF
C74973 INVX1_LOC_30/Y INVX1_LOC_26/Y 0.14fF
C74974 NOR2X1_LOC_74/Y NOR2X1_LOC_89/A 0.02fF
C74975 NOR2X1_LOC_226/A NAND2X1_LOC_860/A 0.01fF
C74976 NOR2X1_LOC_646/A NOR2X1_LOC_646/B 0.02fF
C74977 INPUT_0 INVX1_LOC_99/A 0.02fF
C74978 NAND2X1_LOC_555/Y INVX1_LOC_40/Y 0.02fF
C74979 INVX1_LOC_286/Y INVX1_LOC_141/Y 0.01fF
C74980 INVX1_LOC_75/A NOR2X1_LOC_460/A 0.01fF
C74981 NOR2X1_LOC_27/Y INVX1_LOC_5/A 0.00fF
C74982 INVX1_LOC_14/A INVX1_LOC_314/Y 0.11fF
C74983 INVX1_LOC_58/A INVX1_LOC_25/Y 0.01fF
C74984 INVX1_LOC_303/A INVX1_LOC_24/Y 0.10fF
C74985 INVX1_LOC_245/Y NOR2X1_LOC_68/A 0.02fF
C74986 NOR2X1_LOC_690/A NOR2X1_LOC_824/A 0.02fF
C74987 INVX1_LOC_96/A INVX1_LOC_19/A 0.02fF
C74988 NAND2X1_LOC_452/a_36_24# INVX1_LOC_53/A 0.00fF
C74989 NOR2X1_LOC_92/Y NOR2X1_LOC_672/Y 0.02fF
C74990 NOR2X1_LOC_328/Y NOR2X1_LOC_696/Y 0.01fF
C74991 INVX1_LOC_294/Y NAND2X1_LOC_474/Y 0.44fF
C74992 INVX1_LOC_286/Y INVX1_LOC_312/Y 0.04fF
C74993 NOR2X1_LOC_255/Y INVX1_LOC_232/A 0.02fF
C74994 NAND2X1_LOC_364/A NAND2X1_LOC_352/B 0.25fF
C74995 NOR2X1_LOC_423/a_36_216# NOR2X1_LOC_222/Y 0.00fF
C74996 INVX1_LOC_75/A INVX1_LOC_3/Y 0.10fF
C74997 NAND2X1_LOC_208/a_36_24# NOR2X1_LOC_84/Y 0.06fF
C74998 NOR2X1_LOC_82/A D_INPUT_2 2.75fF
C74999 INVX1_LOC_13/Y NOR2X1_LOC_398/Y 0.02fF
C75000 INVX1_LOC_224/Y NOR2X1_LOC_391/A 0.07fF
C75001 NAND2X1_LOC_9/Y NOR2X1_LOC_516/B 0.03fF
C75002 INVX1_LOC_285/Y NAND2X1_LOC_792/B 0.19fF
C75003 INVX1_LOC_90/A NOR2X1_LOC_278/Y 0.05fF
C75004 NOR2X1_LOC_536/A NAND2X1_LOC_243/Y 0.01fF
C75005 NAND2X1_LOC_67/Y INVX1_LOC_63/Y 0.60fF
C75006 NOR2X1_LOC_15/Y NAND2X1_LOC_811/Y 0.09fF
C75007 NAND2X1_LOC_649/B INVX1_LOC_49/Y 0.06fF
C75008 INVX1_LOC_279/A INVX1_LOC_23/A 0.21fF
C75009 INVX1_LOC_135/A NOR2X1_LOC_654/A 0.12fF
C75010 NOR2X1_LOC_667/A NOR2X1_LOC_406/A 0.03fF
C75011 NOR2X1_LOC_292/Y INVX1_LOC_47/Y 0.03fF
C75012 NAND2X1_LOC_808/A INVX1_LOC_57/A 0.07fF
C75013 NAND2X1_LOC_81/B NAND2X1_LOC_642/Y 0.04fF
C75014 NOR2X1_LOC_815/Y NOR2X1_LOC_513/Y 0.07fF
C75015 INVX1_LOC_248/A NOR2X1_LOC_406/A 0.02fF
C75016 D_INPUT_1 INVX1_LOC_306/A 0.02fF
C75017 NOR2X1_LOC_187/a_36_216# INVX1_LOC_290/Y 0.01fF
C75018 NOR2X1_LOC_91/A NOR2X1_LOC_166/a_36_216# 0.01fF
C75019 NAND2X1_LOC_659/B NAND2X1_LOC_82/Y 0.01fF
C75020 INVX1_LOC_185/A INVX1_LOC_54/A 0.05fF
C75021 INVX1_LOC_226/Y INVX1_LOC_306/Y 0.06fF
C75022 NOR2X1_LOC_826/Y INVX1_LOC_234/A 0.03fF
C75023 NOR2X1_LOC_658/Y INVX1_LOC_24/A 0.00fF
C75024 NOR2X1_LOC_15/Y INVX1_LOC_266/Y 0.10fF
C75025 INVX1_LOC_5/A NOR2X1_LOC_687/Y 0.05fF
C75026 INVX1_LOC_88/A NAND2X1_LOC_477/A 0.03fF
C75027 INVX1_LOC_13/Y NOR2X1_LOC_211/A 0.10fF
C75028 NOR2X1_LOC_634/A NOR2X1_LOC_729/A 0.01fF
C75029 NOR2X1_LOC_798/A NOR2X1_LOC_516/B 0.03fF
C75030 INVX1_LOC_91/A NOR2X1_LOC_460/a_36_216# 0.00fF
C75031 INVX1_LOC_2/A NAND2X1_LOC_537/Y 0.79fF
C75032 INVX1_LOC_35/Y INVX1_LOC_118/A 0.01fF
C75033 INVX1_LOC_163/A NOR2X1_LOC_399/Y 0.05fF
C75034 INVX1_LOC_34/A INVX1_LOC_161/A 0.19fF
C75035 NOR2X1_LOC_824/A NAND2X1_LOC_717/a_36_24# 0.00fF
C75036 NAND2X1_LOC_363/B NAND2X1_LOC_363/Y 0.27fF
C75037 NAND2X1_LOC_579/A NAND2X1_LOC_850/Y 0.03fF
C75038 VDD NAND2X1_LOC_82/Y 0.46fF
C75039 NOR2X1_LOC_833/Y NOR2X1_LOC_833/B 0.19fF
C75040 INVX1_LOC_215/Y NOR2X1_LOC_320/a_36_216# 0.00fF
C75041 INVX1_LOC_269/A NAND2X1_LOC_338/B 0.33fF
C75042 INVX1_LOC_6/A INVX1_LOC_271/Y 0.11fF
C75043 NAND2X1_LOC_860/A INPUT_1 0.25fF
C75044 NOR2X1_LOC_226/A NAND2X1_LOC_537/Y 0.10fF
C75045 NAND2X1_LOC_363/B INVX1_LOC_89/A 0.18fF
C75046 INVX1_LOC_17/A NAND2X1_LOC_342/Y 0.01fF
C75047 INVX1_LOC_10/A INVX1_LOC_306/Y 0.02fF
C75048 NAND2X1_LOC_9/Y NOR2X1_LOC_756/a_36_216# 0.00fF
C75049 INVX1_LOC_41/A NOR2X1_LOC_500/B 0.03fF
C75050 NOR2X1_LOC_13/Y INVX1_LOC_24/A 0.01fF
C75051 NAND2X1_LOC_721/B NAND2X1_LOC_325/Y 0.22fF
C75052 NOR2X1_LOC_91/A NAND2X1_LOC_858/B 0.03fF
C75053 INVX1_LOC_182/Y INVX1_LOC_23/A 0.03fF
C75054 VDD NOR2X1_LOC_461/Y 0.12fF
C75055 NOR2X1_LOC_99/B NOR2X1_LOC_849/A 0.04fF
C75056 INVX1_LOC_58/A INVX1_LOC_75/A 0.11fF
C75057 INVX1_LOC_62/A INVX1_LOC_50/Y 0.08fF
C75058 NAND2X1_LOC_303/Y NOR2X1_LOC_695/Y 0.32fF
C75059 INVX1_LOC_280/A NAND2X1_LOC_219/B 0.02fF
C75060 INVX1_LOC_299/Y NOR2X1_LOC_810/Y 0.01fF
C75061 NAND2X1_LOC_833/Y INVX1_LOC_18/A 0.08fF
C75062 NAND2X1_LOC_96/A NAND2X1_LOC_74/B 0.10fF
C75063 NAND2X1_LOC_642/Y INVX1_LOC_4/Y 0.04fF
C75064 INVX1_LOC_12/Y INVX1_LOC_284/A 0.06fF
C75065 VDD NOR2X1_LOC_640/B 0.12fF
C75066 INVX1_LOC_136/A INVX1_LOC_162/A 0.02fF
C75067 INVX1_LOC_143/Y INVX1_LOC_15/A 0.05fF
C75068 INVX1_LOC_36/A NOR2X1_LOC_574/A 0.04fF
C75069 NAND2X1_LOC_306/a_36_24# NOR2X1_LOC_577/Y 0.00fF
C75070 INVX1_LOC_57/Y NOR2X1_LOC_52/B 0.10fF
C75071 INVX1_LOC_43/Y INVX1_LOC_43/A 0.19fF
C75072 NOR2X1_LOC_609/A NOR2X1_LOC_388/Y 0.04fF
C75073 NOR2X1_LOC_794/B NOR2X1_LOC_388/a_36_216# 0.00fF
C75074 INVX1_LOC_136/A NOR2X1_LOC_315/Y 0.07fF
C75075 NOR2X1_LOC_754/a_36_216# NOR2X1_LOC_754/Y 0.00fF
C75076 NAND2X1_LOC_357/B NAND2X1_LOC_364/A 0.11fF
C75077 NAND2X1_LOC_141/Y NAND2X1_LOC_574/A 0.74fF
C75078 NOR2X1_LOC_75/Y NAND2X1_LOC_479/Y 0.03fF
C75079 INVX1_LOC_58/A NOR2X1_LOC_7/a_36_216# 0.00fF
C75080 INVX1_LOC_255/Y NOR2X1_LOC_647/B 0.00fF
C75081 INVX1_LOC_172/A NAND2X1_LOC_833/Y 1.24fF
C75082 NAND2X1_LOC_170/a_36_24# INVX1_LOC_28/A 0.00fF
C75083 NOR2X1_LOC_391/A NOR2X1_LOC_103/Y 0.09fF
C75084 NOR2X1_LOC_52/B NOR2X1_LOC_512/Y 0.02fF
C75085 INVX1_LOC_41/A INVX1_LOC_303/A 0.18fF
C75086 INVX1_LOC_21/A NAND2X1_LOC_654/B 0.01fF
C75087 NAND2X1_LOC_740/Y NOR2X1_LOC_385/Y 0.02fF
C75088 NAND2X1_LOC_447/Y INVX1_LOC_26/A 0.11fF
C75089 INVX1_LOC_250/A NOR2X1_LOC_667/A 0.01fF
C75090 NOR2X1_LOC_334/Y INVX1_LOC_37/A 0.07fF
C75091 NOR2X1_LOC_759/Y NOR2X1_LOC_423/Y 0.01fF
C75092 INVX1_LOC_24/A NOR2X1_LOC_504/Y 0.07fF
C75093 NAND2X1_LOC_785/Y NOR2X1_LOC_495/Y 0.34fF
C75094 INVX1_LOC_269/A INVX1_LOC_313/Y 0.00fF
C75095 NOR2X1_LOC_226/A NAND2X1_LOC_640/a_36_24# 0.00fF
C75096 INVX1_LOC_85/A INVX1_LOC_113/Y 0.00fF
C75097 INVX1_LOC_230/Y INVX1_LOC_219/A 0.05fF
C75098 NOR2X1_LOC_67/A NOR2X1_LOC_256/a_36_216# 0.00fF
C75099 NAND2X1_LOC_269/a_36_24# NOR2X1_LOC_271/Y 0.01fF
C75100 NOR2X1_LOC_372/Y INVX1_LOC_16/A 0.04fF
C75101 NOR2X1_LOC_89/A INVX1_LOC_179/A 0.03fF
C75102 INVX1_LOC_185/A NOR2X1_LOC_48/B 0.05fF
C75103 INVX1_LOC_88/A NOR2X1_LOC_122/Y 0.02fF
C75104 NOR2X1_LOC_273/Y NOR2X1_LOC_222/Y 0.02fF
C75105 NOR2X1_LOC_74/A NAND2X1_LOC_474/Y 0.24fF
C75106 NOR2X1_LOC_222/Y NOR2X1_LOC_759/Y 1.20fF
C75107 NOR2X1_LOC_552/A INVX1_LOC_58/Y 0.09fF
C75108 INVX1_LOC_63/Y NOR2X1_LOC_367/B 0.03fF
C75109 NOR2X1_LOC_843/A NOR2X1_LOC_288/A -0.00fF
C75110 INVX1_LOC_4/Y NOR2X1_LOC_271/Y 0.02fF
C75111 D_INPUT_1 INVX1_LOC_59/Y 0.03fF
C75112 NOR2X1_LOC_447/B NOR2X1_LOC_447/A 0.00fF
C75113 INVX1_LOC_17/A NAND2X1_LOC_7/a_36_24# 0.01fF
C75114 INVX1_LOC_13/A NOR2X1_LOC_791/B 0.03fF
C75115 NOR2X1_LOC_9/Y NAND2X1_LOC_474/Y 0.10fF
C75116 INVX1_LOC_2/Y NOR2X1_LOC_646/B 0.00fF
C75117 VDD NOR2X1_LOC_840/Y -0.00fF
C75118 NOR2X1_LOC_781/A INVX1_LOC_18/A 0.02fF
C75119 NOR2X1_LOC_657/Y INVX1_LOC_10/A 0.02fF
C75120 NOR2X1_LOC_15/Y INVX1_LOC_42/Y 0.00fF
C75121 NAND2X1_LOC_364/Y INVX1_LOC_143/A 0.32fF
C75122 NAND2X1_LOC_579/A INVX1_LOC_282/A 0.16fF
C75123 NOR2X1_LOC_598/B NOR2X1_LOC_833/Y 0.19fF
C75124 INVX1_LOC_141/Y NAND2X1_LOC_803/a_36_24# 0.00fF
C75125 INVX1_LOC_77/A NAND2X1_LOC_9/a_36_24# 0.01fF
C75126 NAND2X1_LOC_555/Y NAND2X1_LOC_28/a_36_24# 0.00fF
C75127 NAND2X1_LOC_866/A NAND2X1_LOC_853/Y 1.03fF
C75128 NOR2X1_LOC_160/B NAND2X1_LOC_842/B 0.03fF
C75129 INVX1_LOC_24/A NOR2X1_LOC_146/Y 0.05fF
C75130 INVX1_LOC_41/A NAND2X1_LOC_610/a_36_24# 0.00fF
C75131 NOR2X1_LOC_89/A NAND2X1_LOC_267/a_36_24# 0.01fF
C75132 NOR2X1_LOC_89/A INVX1_LOC_250/Y 0.01fF
C75133 INVX1_LOC_236/Y INVX1_LOC_90/A 0.03fF
C75134 INVX1_LOC_11/A NOR2X1_LOC_163/Y 0.02fF
C75135 NOR2X1_LOC_78/B INVX1_LOC_155/A 0.02fF
C75136 INVX1_LOC_34/A NAND2X1_LOC_231/Y 0.00fF
C75137 INVX1_LOC_58/A NAND2X1_LOC_453/A 0.03fF
C75138 NOR2X1_LOC_598/B INVX1_LOC_115/A 0.00fF
C75139 INVX1_LOC_38/A NOR2X1_LOC_278/Y 0.02fF
C75140 INVX1_LOC_50/A NAND2X1_LOC_804/Y 0.11fF
C75141 NAND2X1_LOC_794/B INVX1_LOC_91/A 0.10fF
C75142 NOR2X1_LOC_32/B INVX1_LOC_20/A 0.33fF
C75143 INVX1_LOC_89/A INVX1_LOC_30/A 1.14fF
C75144 INVX1_LOC_17/A INVX1_LOC_67/Y 0.05fF
C75145 NOR2X1_LOC_859/A NOR2X1_LOC_99/B 0.03fF
C75146 NAND2X1_LOC_773/Y INVX1_LOC_6/A 0.03fF
C75147 NOR2X1_LOC_67/A INVX1_LOC_8/A 0.13fF
C75148 NAND2X1_LOC_728/Y INVX1_LOC_273/Y 0.24fF
C75149 NOR2X1_LOC_536/A NOR2X1_LOC_39/Y 0.46fF
C75150 INVX1_LOC_11/A NOR2X1_LOC_74/Y 0.01fF
C75151 NAND2X1_LOC_763/B INVX1_LOC_89/A 0.45fF
C75152 NOR2X1_LOC_68/A D_INPUT_0 0.12fF
C75153 NAND2X1_LOC_53/Y NOR2X1_LOC_74/A 0.17fF
C75154 NOR2X1_LOC_214/B INVX1_LOC_72/A 0.01fF
C75155 INVX1_LOC_96/Y INVX1_LOC_266/Y 0.10fF
C75156 NOR2X1_LOC_391/A INVX1_LOC_71/A 0.07fF
C75157 INVX1_LOC_38/A NOR2X1_LOC_638/Y 0.00fF
C75158 NAND2X1_LOC_500/Y NOR2X1_LOC_497/Y 0.05fF
C75159 INVX1_LOC_34/A NAND2X1_LOC_195/a_36_24# 0.01fF
C75160 NAND2X1_LOC_794/B INVX1_LOC_11/Y 0.06fF
C75161 NOR2X1_LOC_305/Y NOR2X1_LOC_109/Y 0.01fF
C75162 NAND2X1_LOC_286/B INVX1_LOC_118/A 0.04fF
C75163 NOR2X1_LOC_180/B INVX1_LOC_18/A 0.07fF
C75164 NAND2X1_LOC_326/A NOR2X1_LOC_45/B 0.08fF
C75165 NAND2X1_LOC_114/B NOR2X1_LOC_721/Y 0.19fF
C75166 INVX1_LOC_251/Y NAND2X1_LOC_360/B 0.09fF
C75167 NOR2X1_LOC_13/Y NOR2X1_LOC_130/A 0.05fF
C75168 INVX1_LOC_28/A NOR2X1_LOC_372/Y 0.13fF
C75169 NOR2X1_LOC_175/A INVX1_LOC_179/Y 0.02fF
C75170 INVX1_LOC_124/A NOR2X1_LOC_773/Y 0.01fF
C75171 NOR2X1_LOC_68/A NAND2X1_LOC_665/a_36_24# 0.01fF
C75172 INVX1_LOC_161/A INPUT_0 0.11fF
C75173 NOR2X1_LOC_705/B INVX1_LOC_193/Y 0.00fF
C75174 INVX1_LOC_77/A NOR2X1_LOC_332/A 0.03fF
C75175 NOR2X1_LOC_589/A NOR2X1_LOC_364/Y 0.05fF
C75176 NAND2X1_LOC_189/a_36_24# INVX1_LOC_94/A 0.00fF
C75177 NAND2X1_LOC_858/B INVX1_LOC_31/A 0.07fF
C75178 NOR2X1_LOC_561/Y INVX1_LOC_63/Y 0.14fF
C75179 NOR2X1_LOC_563/a_36_216# INVX1_LOC_104/A 0.00fF
C75180 NOR2X1_LOC_536/Y NAND2X1_LOC_729/B 0.19fF
C75181 NAND2X1_LOC_208/B INPUT_0 0.00fF
C75182 NAND2X1_LOC_358/B NAND2X1_LOC_96/A 0.03fF
C75183 NAND2X1_LOC_839/A NAND2X1_LOC_835/a_36_24# 0.02fF
C75184 INVX1_LOC_290/Y INVX1_LOC_263/Y 0.04fF
C75185 INVX1_LOC_135/A NOR2X1_LOC_716/B 0.10fF
C75186 INVX1_LOC_53/Y NOR2X1_LOC_709/A 0.07fF
C75187 NOR2X1_LOC_690/A INVX1_LOC_234/A 0.01fF
C75188 INVX1_LOC_243/Y INVX1_LOC_92/A 0.03fF
C75189 NOR2X1_LOC_131/A NOR2X1_LOC_131/Y 0.19fF
C75190 INVX1_LOC_73/A INVX1_LOC_18/A 0.07fF
C75191 NOR2X1_LOC_413/Y INVX1_LOC_234/A 0.03fF
C75192 INVX1_LOC_90/A NAND2X1_LOC_7/Y 0.01fF
C75193 NAND2X1_LOC_860/A INVX1_LOC_118/A 0.15fF
C75194 NOR2X1_LOC_419/Y NOR2X1_LOC_560/A 0.02fF
C75195 NAND2X1_LOC_853/Y NOR2X1_LOC_505/Y 0.09fF
C75196 INVX1_LOC_52/Y INVX1_LOC_76/A -0.07fF
C75197 INVX1_LOC_49/A INVX1_LOC_85/Y 0.03fF
C75198 INVX1_LOC_290/Y INVX1_LOC_42/A 0.07fF
C75199 NOR2X1_LOC_301/A INVX1_LOC_285/A 0.07fF
C75200 INVX1_LOC_57/A INVX1_LOC_92/A 14.57fF
C75201 NOR2X1_LOC_754/Y INVX1_LOC_54/A 0.01fF
C75202 NAND2X1_LOC_374/Y INVX1_LOC_16/A 0.21fF
C75203 NAND2X1_LOC_93/B NAND2X1_LOC_205/A 0.02fF
C75204 INVX1_LOC_1/A NOR2X1_LOC_603/Y 0.01fF
C75205 NOR2X1_LOC_589/A NOR2X1_LOC_131/A 0.06fF
C75206 INVX1_LOC_249/A NOR2X1_LOC_736/a_36_216# 0.00fF
C75207 NOR2X1_LOC_677/Y NOR2X1_LOC_88/Y 0.01fF
C75208 VDD NAND2X1_LOC_780/Y 0.02fF
C75209 NAND2X1_LOC_600/a_36_24# NOR2X1_LOC_109/Y 0.01fF
C75210 NOR2X1_LOC_6/B INVX1_LOC_62/A 0.00fF
C75211 NAND2X1_LOC_352/B NOR2X1_LOC_405/A 0.03fF
C75212 NOR2X1_LOC_273/a_36_216# NAND2X1_LOC_832/Y 0.00fF
C75213 INVX1_LOC_229/Y NOR2X1_LOC_822/Y 0.03fF
C75214 NOR2X1_LOC_38/B NOR2X1_LOC_664/a_36_216# 0.00fF
C75215 INVX1_LOC_5/A INVX1_LOC_9/A 2.90fF
C75216 NOR2X1_LOC_576/B NOR2X1_LOC_821/Y 0.04fF
C75217 NAND2X1_LOC_540/a_36_24# NOR2X1_LOC_271/Y 0.00fF
C75218 NOR2X1_LOC_516/Y INPUT_1 0.01fF
C75219 NOR2X1_LOC_78/B INVX1_LOC_160/Y 0.06fF
C75220 INVX1_LOC_13/A NAND2X1_LOC_672/B 0.01fF
C75221 INVX1_LOC_24/A NOR2X1_LOC_337/A 0.06fF
C75222 INVX1_LOC_83/A NAND2X1_LOC_661/B 0.28fF
C75223 INVX1_LOC_36/A NOR2X1_LOC_588/A 0.01fF
C75224 INVX1_LOC_45/Y INVX1_LOC_69/Y 0.00fF
C75225 NOR2X1_LOC_413/Y NOR2X1_LOC_19/B 0.19fF
C75226 INVX1_LOC_256/Y NOR2X1_LOC_130/A 0.03fF
C75227 NAND2X1_LOC_323/B NOR2X1_LOC_97/a_36_216# 0.00fF
C75228 NOR2X1_LOC_75/Y INVX1_LOC_139/Y 0.48fF
C75229 NOR2X1_LOC_700/Y NAND2X1_LOC_853/Y 0.01fF
C75230 NOR2X1_LOC_648/a_36_216# INVX1_LOC_313/Y 0.00fF
C75231 NOR2X1_LOC_360/Y NOR2X1_LOC_78/A 0.03fF
C75232 NAND2X1_LOC_114/B VDD 0.38fF
C75233 INVX1_LOC_78/A INVX1_LOC_290/Y 0.07fF
C75234 INVX1_LOC_36/A INVX1_LOC_95/Y 0.10fF
C75235 NAND2X1_LOC_74/B NAND2X1_LOC_99/A 1.26fF
C75236 INVX1_LOC_232/Y INVX1_LOC_90/A 0.03fF
C75237 INVX1_LOC_34/A INPUT_0 0.28fF
C75238 INVX1_LOC_15/A NOR2X1_LOC_227/A 0.20fF
C75239 INVX1_LOC_72/A NOR2X1_LOC_275/A 0.00fF
C75240 NOR2X1_LOC_89/A NOR2X1_LOC_693/Y 1.11fF
C75241 INVX1_LOC_39/Y VDD 0.41fF
C75242 NOR2X1_LOC_106/A INVX1_LOC_53/Y 0.01fF
C75243 NAND2X1_LOC_543/Y NAND2X1_LOC_861/Y 0.02fF
C75244 NOR2X1_LOC_264/Y NOR2X1_LOC_193/a_36_216# 0.00fF
C75245 NAND2X1_LOC_374/Y INVX1_LOC_28/A 0.19fF
C75246 INVX1_LOC_141/Y VDD 0.41fF
C75247 NOR2X1_LOC_836/Y INVX1_LOC_37/A 0.00fF
C75248 NAND2X1_LOC_537/Y INVX1_LOC_118/A 0.01fF
C75249 INVX1_LOC_50/A NOR2X1_LOC_519/a_36_216# 0.00fF
C75250 NOR2X1_LOC_45/B NOR2X1_LOC_625/Y 0.01fF
C75251 INVX1_LOC_96/Y INVX1_LOC_42/Y 0.01fF
C75252 NOR2X1_LOC_500/Y NOR2X1_LOC_356/A 0.01fF
C75253 INVX1_LOC_312/Y VDD 1.04fF
C75254 NOR2X1_LOC_294/Y VDD 0.69fF
C75255 NOR2X1_LOC_392/B NOR2X1_LOC_391/Y -0.00fF
C75256 NOR2X1_LOC_335/A NOR2X1_LOC_318/B 0.01fF
C75257 NOR2X1_LOC_602/A NOR2X1_LOC_111/A 0.02fF
C75258 NAND2X1_LOC_807/B INVX1_LOC_270/Y 0.20fF
C75259 NAND2X1_LOC_860/A NAND2X1_LOC_63/Y 0.20fF
C75260 NOR2X1_LOC_460/B INVX1_LOC_91/A 0.01fF
C75261 INVX1_LOC_232/Y NAND2X1_LOC_348/A 0.16fF
C75262 INVX1_LOC_145/Y NOR2X1_LOC_106/A 0.00fF
C75263 NOR2X1_LOC_759/Y NOR2X1_LOC_69/A 0.00fF
C75264 NAND2X1_LOC_9/Y NAND2X1_LOC_207/B 0.07fF
C75265 NOR2X1_LOC_817/Y NOR2X1_LOC_655/Y 0.03fF
C75266 NOR2X1_LOC_189/A INVX1_LOC_11/Y 0.03fF
C75267 INVX1_LOC_212/Y NOR2X1_LOC_349/A 0.01fF
C75268 D_INPUT_2 INVX1_LOC_59/Y 0.05fF
C75269 NAND2X1_LOC_231/Y INPUT_0 1.13fF
C75270 NOR2X1_LOC_644/B NOR2X1_LOC_331/B 0.03fF
C75271 INVX1_LOC_236/Y INVX1_LOC_38/A 0.03fF
C75272 NOR2X1_LOC_733/Y INVX1_LOC_266/Y 0.02fF
C75273 INVX1_LOC_284/Y INVX1_LOC_38/A 0.03fF
C75274 INVX1_LOC_58/A INVX1_LOC_283/A 0.02fF
C75275 NOR2X1_LOC_529/a_36_216# INVX1_LOC_3/Y 0.01fF
C75276 NOR2X1_LOC_286/Y NOR2X1_LOC_634/A 0.01fF
C75277 NOR2X1_LOC_353/a_36_216# NOR2X1_LOC_35/Y 0.00fF
C75278 NOR2X1_LOC_68/A NOR2X1_LOC_859/Y 0.01fF
C75279 INVX1_LOC_36/A NAND2X1_LOC_446/a_36_24# 0.00fF
C75280 INVX1_LOC_11/A INVX1_LOC_179/A 0.05fF
C75281 NAND2X1_LOC_471/Y INVX1_LOC_23/Y 0.05fF
C75282 NAND2X1_LOC_181/Y INVX1_LOC_100/A 0.03fF
C75283 INVX1_LOC_135/A NOR2X1_LOC_130/Y -0.02fF
C75284 INVX1_LOC_13/A INVX1_LOC_82/Y 0.01fF
C75285 INVX1_LOC_135/A NOR2X1_LOC_828/A 0.04fF
C75286 NOR2X1_LOC_500/Y NOR2X1_LOC_74/A 1.50fF
C75287 INVX1_LOC_277/A NOR2X1_LOC_499/B 0.07fF
C75288 INVX1_LOC_90/A NOR2X1_LOC_312/Y 0.00fF
C75289 NAND2X1_LOC_849/A NOR2X1_LOC_86/A 0.06fF
C75290 NAND2X1_LOC_569/A NOR2X1_LOC_368/Y 0.01fF
C75291 INVX1_LOC_53/A NAND2X1_LOC_419/a_36_24# 0.01fF
C75292 INVX1_LOC_41/Y NOR2X1_LOC_176/Y 0.18fF
C75293 INVX1_LOC_147/A NAND2X1_LOC_660/Y 0.07fF
C75294 NOR2X1_LOC_68/A NAND2X1_LOC_848/A 2.42fF
C75295 NOR2X1_LOC_441/Y INVX1_LOC_185/A 0.15fF
C75296 NOR2X1_LOC_482/Y INVX1_LOC_91/A 0.03fF
C75297 INVX1_LOC_12/A INVX1_LOC_306/Y 0.07fF
C75298 NOR2X1_LOC_230/Y INVX1_LOC_54/A 0.04fF
C75299 NOR2X1_LOC_309/Y INVX1_LOC_95/Y 0.03fF
C75300 INVX1_LOC_222/Y NAND2X1_LOC_74/B 0.03fF
C75301 INVX1_LOC_17/A INVX1_LOC_285/A 0.07fF
C75302 NOR2X1_LOC_174/A NOR2X1_LOC_174/B 0.02fF
C75303 INVX1_LOC_23/A NOR2X1_LOC_38/B 0.00fF
C75304 INVX1_LOC_63/Y INVX1_LOC_76/A 0.12fF
C75305 INVX1_LOC_275/A VDD -0.00fF
C75306 INVX1_LOC_270/A INVX1_LOC_271/Y 0.09fF
C75307 NOR2X1_LOC_533/Y INVX1_LOC_84/A 0.03fF
C75308 NOR2X1_LOC_817/Y NOR2X1_LOC_649/B 0.03fF
C75309 INVX1_LOC_11/A INVX1_LOC_250/Y 0.01fF
C75310 NOR2X1_LOC_219/B VDD 0.12fF
C75311 INVX1_LOC_5/A NOR2X1_LOC_861/Y 0.14fF
C75312 INVX1_LOC_17/A NOR2X1_LOC_814/A 0.15fF
C75313 NAND2X1_LOC_483/Y VDD 0.08fF
C75314 INVX1_LOC_10/A NOR2X1_LOC_74/A 0.07fF
C75315 NOR2X1_LOC_15/Y INVX1_LOC_19/A 0.10fF
C75316 NOR2X1_LOC_84/A D_INPUT_3 0.07fF
C75317 INVX1_LOC_149/A NAND2X1_LOC_447/Y 0.03fF
C75318 NOR2X1_LOC_147/B NOR2X1_LOC_858/B 0.26fF
C75319 NOR2X1_LOC_92/Y INVX1_LOC_272/A 0.10fF
C75320 NAND2X1_LOC_550/A INVX1_LOC_119/Y 0.00fF
C75321 VDD INVX1_LOC_88/Y 0.31fF
C75322 NOR2X1_LOC_191/A INVX1_LOC_93/Y 0.03fF
C75323 INVX1_LOC_279/A INVX1_LOC_6/A 0.07fF
C75324 NAND2X1_LOC_323/a_36_24# NOR2X1_LOC_356/A 0.00fF
C75325 NAND2X1_LOC_7/Y INVX1_LOC_38/A 0.03fF
C75326 NOR2X1_LOC_718/B INVX1_LOC_37/A 0.07fF
C75327 INVX1_LOC_33/A INVX1_LOC_202/Y 0.00fF
C75328 INVX1_LOC_10/A NOR2X1_LOC_9/Y 0.04fF
C75329 NAND2X1_LOC_623/B INVX1_LOC_22/A 0.03fF
C75330 INVX1_LOC_290/A INVX1_LOC_91/A 0.04fF
C75331 NOR2X1_LOC_352/Y NOR2X1_LOC_35/Y 0.29fF
C75332 NAND2X1_LOC_112/Y NOR2X1_LOC_269/Y 0.00fF
C75333 NAND2X1_LOC_555/Y NOR2X1_LOC_814/A 1.33fF
C75334 NOR2X1_LOC_68/A INVX1_LOC_46/Y 0.38fF
C75335 NAND2X1_LOC_839/A INVX1_LOC_76/A 0.08fF
C75336 NOR2X1_LOC_168/B VDD 0.32fF
C75337 INVX1_LOC_24/A NOR2X1_LOC_640/Y 0.02fF
C75338 NOR2X1_LOC_541/B INVX1_LOC_58/Y 0.02fF
C75339 NOR2X1_LOC_516/B NOR2X1_LOC_545/B 0.06fF
C75340 NOR2X1_LOC_620/B INVX1_LOC_176/A 0.01fF
C75341 NOR2X1_LOC_690/Y NAND2X1_LOC_729/B 0.06fF
C75342 NAND2X1_LOC_858/B NAND2X1_LOC_807/Y 0.07fF
C75343 NAND2X1_LOC_338/B INVX1_LOC_12/Y 0.03fF
C75344 INVX1_LOC_233/A NAND2X1_LOC_442/a_36_24# 0.00fF
C75345 INVX1_LOC_24/A NAND2X1_LOC_85/Y 0.03fF
C75346 INVX1_LOC_53/A INVX1_LOC_57/A 15.85fF
C75347 NOR2X1_LOC_552/Y NOR2X1_LOC_564/Y 0.00fF
C75348 NOR2X1_LOC_160/B INVX1_LOC_284/A 0.04fF
C75349 NOR2X1_LOC_718/B NAND2X1_LOC_629/a_36_24# 0.00fF
C75350 INVX1_LOC_24/A NOR2X1_LOC_697/Y 0.00fF
C75351 INVX1_LOC_41/A NOR2X1_LOC_99/Y 0.02fF
C75352 NOR2X1_LOC_346/B INVX1_LOC_117/A 0.00fF
C75353 NAND2X1_LOC_686/a_36_24# INVX1_LOC_92/A 0.01fF
C75354 NOR2X1_LOC_593/Y INVX1_LOC_179/A 0.01fF
C75355 NOR2X1_LOC_454/Y INVX1_LOC_78/A 0.12fF
C75356 NAND2X1_LOC_348/A NOR2X1_LOC_391/Y 0.00fF
C75357 NOR2X1_LOC_569/Y INVX1_LOC_37/A 0.07fF
C75358 NOR2X1_LOC_667/Y NOR2X1_LOC_48/B 0.01fF
C75359 INVX1_LOC_22/A INVX1_LOC_117/A 0.19fF
C75360 NOR2X1_LOC_828/B NOR2X1_LOC_725/A 0.30fF
C75361 NOR2X1_LOC_32/B INVX1_LOC_64/A 0.08fF
C75362 NOR2X1_LOC_52/B INVX1_LOC_179/A 0.00fF
C75363 NAND2X1_LOC_656/Y VDD 2.17fF
C75364 NOR2X1_LOC_567/B NOR2X1_LOC_78/A 0.08fF
C75365 INVX1_LOC_30/A NOR2X1_LOC_490/a_36_216# 0.00fF
C75366 INVX1_LOC_288/A NOR2X1_LOC_454/Y 0.06fF
C75367 INVX1_LOC_21/A INVX1_LOC_50/A 0.16fF
C75368 NOR2X1_LOC_242/A INVX1_LOC_57/A 0.19fF
C75369 NAND2X1_LOC_803/B NOR2X1_LOC_158/B 0.61fF
C75370 NOR2X1_LOC_860/B INVX1_LOC_19/A 0.07fF
C75371 INVX1_LOC_181/Y INVX1_LOC_29/A 0.08fF
C75372 NAND2X1_LOC_656/A NAND2X1_LOC_74/B 0.00fF
C75373 NAND2X1_LOC_673/a_36_24# INVX1_LOC_84/A 0.00fF
C75374 NOR2X1_LOC_210/A INVX1_LOC_38/A 0.01fF
C75375 NOR2X1_LOC_91/A NOR2X1_LOC_468/Y 0.73fF
C75376 INVX1_LOC_161/Y INVX1_LOC_273/A 0.00fF
C75377 INVX1_LOC_132/Y VDD 0.27fF
C75378 INVX1_LOC_31/A NOR2X1_LOC_38/B 0.15fF
C75379 INVX1_LOC_269/A NAND2X1_LOC_402/B 0.01fF
C75380 NOR2X1_LOC_603/a_36_216# INVX1_LOC_179/A 0.00fF
C75381 INVX1_LOC_45/Y NOR2X1_LOC_89/A 0.13fF
C75382 INVX1_LOC_90/A NAND2X1_LOC_287/B 0.21fF
C75383 NOR2X1_LOC_395/a_36_216# INVX1_LOC_46/A 0.02fF
C75384 INVX1_LOC_144/Y NAND2X1_LOC_798/B -0.02fF
C75385 NOR2X1_LOC_45/B NOR2X1_LOC_815/A 0.07fF
C75386 INVX1_LOC_166/A NOR2X1_LOC_15/Y 0.05fF
C75387 NAND2X1_LOC_638/Y VDD 0.00fF
C75388 NOR2X1_LOC_636/A NAND2X1_LOC_651/B 0.02fF
C75389 NOR2X1_LOC_717/B INVX1_LOC_10/Y 0.14fF
C75390 INVX1_LOC_223/A NOR2X1_LOC_609/Y 0.01fF
C75391 INVX1_LOC_251/Y NAND2X1_LOC_572/B 0.12fF
C75392 NOR2X1_LOC_264/Y NOR2X1_LOC_68/Y 0.08fF
C75393 NOR2X1_LOC_330/a_36_216# NOR2X1_LOC_447/B 0.00fF
C75394 INVX1_LOC_224/Y INVX1_LOC_269/A 0.10fF
C75395 INVX1_LOC_11/A NAND2X1_LOC_288/B 0.24fF
C75396 INVX1_LOC_90/A INVX1_LOC_129/Y 0.00fF
C75397 NAND2X1_LOC_35/Y INVX1_LOC_13/Y 0.01fF
C75398 NAND2X1_LOC_101/a_36_24# INVX1_LOC_42/A 0.01fF
C75399 NOR2X1_LOC_791/B INVX1_LOC_32/A 0.01fF
C75400 INVX1_LOC_34/A NOR2X1_LOC_84/B 0.01fF
C75401 NOR2X1_LOC_468/Y INVX1_LOC_23/A 0.11fF
C75402 INVX1_LOC_144/A NAND2X1_LOC_468/B 0.03fF
C75403 INVX1_LOC_95/A INVX1_LOC_126/Y 0.01fF
C75404 NOR2X1_LOC_525/Y INVX1_LOC_38/A 0.03fF
C75405 INVX1_LOC_21/A NAND2X1_LOC_72/Y 0.01fF
C75406 NAND2X1_LOC_352/a_36_24# NAND2X1_LOC_286/B 0.01fF
C75407 NOR2X1_LOC_590/A NOR2X1_LOC_301/A 0.01fF
C75408 NOR2X1_LOC_332/A INVX1_LOC_9/A 0.11fF
C75409 INVX1_LOC_77/A INVX1_LOC_42/A 0.04fF
C75410 INVX1_LOC_36/A INVX1_LOC_271/Y 0.02fF
C75411 D_INPUT_1 INVX1_LOC_103/A 0.01fF
C75412 NAND2X1_LOC_218/B INVX1_LOC_3/Y 0.04fF
C75413 NOR2X1_LOC_468/Y NOR2X1_LOC_277/a_36_216# 0.00fF
C75414 NOR2X1_LOC_78/A NOR2X1_LOC_269/Y 0.07fF
C75415 NOR2X1_LOC_130/Y INVX1_LOC_280/A -0.02fF
C75416 NAND2X1_LOC_141/A INVX1_LOC_19/A -0.00fF
C75417 NAND2X1_LOC_563/Y INVX1_LOC_29/A 0.04fF
C75418 NAND2X1_LOC_579/A NAND2X1_LOC_624/B 0.03fF
C75419 NAND2X1_LOC_338/B NAND2X1_LOC_465/a_36_24# 0.00fF
C75420 NAND2X1_LOC_477/A INVX1_LOC_272/A 0.07fF
C75421 INVX1_LOC_96/Y INVX1_LOC_19/A 0.14fF
C75422 NAND2X1_LOC_725/A NAND2X1_LOC_725/B 0.07fF
C75423 NAND2X1_LOC_198/B NOR2X1_LOC_334/Y 0.11fF
C75424 VDD NAND2X1_LOC_622/B 0.08fF
C75425 NOR2X1_LOC_595/Y NAND2X1_LOC_642/Y 0.03fF
C75426 D_INPUT_1 INVX1_LOC_292/A 0.03fF
C75427 INVX1_LOC_5/A NAND2X1_LOC_67/Y 0.02fF
C75428 INVX1_LOC_90/A NAND2X1_LOC_260/a_36_24# 0.01fF
C75429 NOR2X1_LOC_389/A INVX1_LOC_23/A 0.22fF
C75430 NOR2X1_LOC_441/Y INVX1_LOC_270/Y 0.01fF
C75431 NOR2X1_LOC_151/Y INVX1_LOC_10/Y 0.03fF
C75432 NAND2X1_LOC_214/B INVX1_LOC_14/A 0.13fF
C75433 INVX1_LOC_136/A NAND2X1_LOC_99/A 0.07fF
C75434 NAND2X1_LOC_11/a_36_24# INPUT_7 0.00fF
C75435 INVX1_LOC_64/A NOR2X1_LOC_218/A 0.01fF
C75436 NOR2X1_LOC_208/Y INVX1_LOC_271/Y 0.11fF
C75437 VDD INVX1_LOC_78/Y 0.51fF
C75438 NAND2X1_LOC_567/Y INVX1_LOC_94/Y 0.02fF
C75439 NAND2X1_LOC_783/A NOR2X1_LOC_697/Y 0.00fF
C75440 NAND2X1_LOC_622/B NAND2X1_LOC_463/a_36_24# 0.01fF
C75441 NOR2X1_LOC_823/Y NOR2X1_LOC_824/Y 0.02fF
C75442 NOR2X1_LOC_124/B INVX1_LOC_32/A 0.07fF
C75443 INVX1_LOC_77/A INVX1_LOC_78/A 0.14fF
C75444 NOR2X1_LOC_443/Y NAND2X1_LOC_364/A 0.02fF
C75445 INVX1_LOC_27/A INVX1_LOC_14/A 2.34fF
C75446 NOR2X1_LOC_130/A NOR2X1_LOC_697/Y 0.17fF
C75447 NOR2X1_LOC_199/B NOR2X1_LOC_814/A 0.06fF
C75448 NOR2X1_LOC_84/a_36_216# INVX1_LOC_3/Y 0.01fF
C75449 INVX1_LOC_58/A NOR2X1_LOC_274/B 0.12fF
C75450 NOR2X1_LOC_823/Y INVX1_LOC_76/A 0.06fF
C75451 NAND2X1_LOC_577/A NOR2X1_LOC_660/Y 0.30fF
C75452 INVX1_LOC_208/A NOR2X1_LOC_755/Y 0.02fF
C75453 INVX1_LOC_316/Y NOR2X1_LOC_671/Y 1.94fF
C75454 NOR2X1_LOC_356/A NOR2X1_LOC_445/B 0.02fF
C75455 INVX1_LOC_286/A NOR2X1_LOC_536/A 0.14fF
C75456 NOR2X1_LOC_160/B NOR2X1_LOC_674/Y 0.39fF
C75457 NOR2X1_LOC_802/A NOR2X1_LOC_623/B 0.02fF
C75458 INVX1_LOC_39/A NOR2X1_LOC_530/a_36_216# 0.00fF
C75459 NAND2X1_LOC_44/a_36_24# INVX1_LOC_53/A 0.00fF
C75460 INVX1_LOC_288/A INVX1_LOC_77/A 0.02fF
C75461 INVX1_LOC_33/A NOR2X1_LOC_278/Y 0.11fF
C75462 NOR2X1_LOC_65/B INVX1_LOC_77/A 0.22fF
C75463 NOR2X1_LOC_433/A NAND2X1_LOC_288/B 0.10fF
C75464 INVX1_LOC_314/Y NOR2X1_LOC_383/B 0.07fF
C75465 NOR2X1_LOC_711/A NOR2X1_LOC_209/B 0.01fF
C75466 NOR2X1_LOC_596/A INVX1_LOC_23/A 0.03fF
C75467 NOR2X1_LOC_556/a_36_216# NOR2X1_LOC_357/Y 0.00fF
C75468 NOR2X1_LOC_516/B NOR2X1_LOC_643/a_36_216# 0.00fF
C75469 INVX1_LOC_47/A INVX1_LOC_63/A 0.00fF
C75470 NOR2X1_LOC_74/A INVX1_LOC_307/A 0.13fF
C75471 INVX1_LOC_124/A INVX1_LOC_78/A 0.05fF
C75472 INVX1_LOC_269/A NOR2X1_LOC_103/Y 0.10fF
C75473 NOR2X1_LOC_15/Y INVX1_LOC_161/Y 0.03fF
C75474 INVX1_LOC_2/A NAND2X1_LOC_454/Y 0.14fF
C75475 NOR2X1_LOC_74/A NOR2X1_LOC_445/B 1.18fF
C75476 INVX1_LOC_269/A NOR2X1_LOC_541/Y 0.02fF
C75477 INVX1_LOC_223/Y INVX1_LOC_30/A 0.03fF
C75478 INVX1_LOC_58/A NOR2X1_LOC_577/Y 0.17fF
C75479 NAND2X1_LOC_342/Y INVX1_LOC_94/Y 0.03fF
C75480 INVX1_LOC_95/A NOR2X1_LOC_536/A 2.28fF
C75481 NOR2X1_LOC_337/A NOR2X1_LOC_197/B 0.01fF
C75482 NOR2X1_LOC_646/A INVX1_LOC_32/A 0.03fF
C75483 INVX1_LOC_124/Y NAND2X1_LOC_474/Y 0.28fF
C75484 INVX1_LOC_286/A NAND2X1_LOC_93/B 0.07fF
C75485 INVX1_LOC_27/A NOR2X1_LOC_717/Y 0.01fF
C75486 NOR2X1_LOC_617/Y NAND2X1_LOC_827/a_36_24# 0.01fF
C75487 NOR2X1_LOC_52/B NOR2X1_LOC_693/Y 0.07fF
C75488 NOR2X1_LOC_668/a_36_216# NOR2X1_LOC_350/A 0.00fF
C75489 INVX1_LOC_17/A NAND2X1_LOC_803/B 0.03fF
C75490 NOR2X1_LOC_201/A NOR2X1_LOC_844/A 0.16fF
C75491 INVX1_LOC_143/A NAND2X1_LOC_221/a_36_24# 0.00fF
C75492 NOR2X1_LOC_71/Y NOR2X1_LOC_89/A 0.12fF
C75493 INVX1_LOC_152/Y INVX1_LOC_77/A 0.03fF
C75494 NAND2X1_LOC_391/Y NOR2X1_LOC_384/Y 0.16fF
C75495 INVX1_LOC_75/A NAND2X1_LOC_475/Y 0.10fF
C75496 INVX1_LOC_172/Y NAND2X1_LOC_618/Y 0.02fF
C75497 NOR2X1_LOC_817/Y NOR2X1_LOC_647/B 0.02fF
C75498 INVX1_LOC_245/Y NAND2X1_LOC_53/Y 0.02fF
C75499 NOR2X1_LOC_65/B INVX1_LOC_124/A 0.27fF
C75500 INVX1_LOC_35/A NOR2X1_LOC_550/B 0.01fF
C75501 NOR2X1_LOC_592/A INVX1_LOC_246/A 0.00fF
C75502 NAND2X1_LOC_472/Y INVX1_LOC_37/A 0.08fF
C75503 NOR2X1_LOC_295/Y INVX1_LOC_23/A 0.00fF
C75504 INVX1_LOC_17/A NOR2X1_LOC_590/A 0.18fF
C75505 NOR2X1_LOC_15/Y NOR2X1_LOC_599/A 0.02fF
C75506 NOR2X1_LOC_593/Y NOR2X1_LOC_405/Y 0.01fF
C75507 NAND2X1_LOC_560/A NAND2X1_LOC_500/B 0.01fF
C75508 NOR2X1_LOC_218/Y NAND2X1_LOC_454/Y 0.02fF
C75509 NOR2X1_LOC_329/B NAND2X1_LOC_74/B 0.07fF
C75510 INVX1_LOC_58/A NOR2X1_LOC_348/B 0.03fF
C75511 INVX1_LOC_45/A INVX1_LOC_269/A 0.17fF
C75512 NOR2X1_LOC_139/Y NOR2X1_LOC_155/A 0.38fF
C75513 INVX1_LOC_313/Y NOR2X1_LOC_842/a_36_216# 0.00fF
C75514 INVX1_LOC_64/A INVX1_LOC_155/Y 0.01fF
C75515 NOR2X1_LOC_474/A INVX1_LOC_253/Y 0.32fF
C75516 NOR2X1_LOC_543/A INVX1_LOC_4/Y 0.02fF
C75517 INVX1_LOC_64/A NOR2X1_LOC_364/Y 0.01fF
C75518 NAND2X1_LOC_363/B INVX1_LOC_176/Y 0.03fF
C75519 NOR2X1_LOC_778/B NOR2X1_LOC_383/B 0.10fF
C75520 NOR2X1_LOC_641/B INVX1_LOC_11/A 0.05fF
C75521 INVX1_LOC_233/Y NAND2X1_LOC_736/B 0.01fF
C75522 NOR2X1_LOC_634/B INVX1_LOC_57/A 0.05fF
C75523 INVX1_LOC_50/A NOR2X1_LOC_667/A 0.19fF
C75524 NOR2X1_LOC_78/B INVX1_LOC_57/A 0.06fF
C75525 INVX1_LOC_50/A INVX1_LOC_248/A 0.07fF
C75526 NAND2X1_LOC_35/Y NOR2X1_LOC_234/a_36_216# 0.01fF
C75527 NOR2X1_LOC_215/A INVX1_LOC_77/A 0.01fF
C75528 NAND2X1_LOC_468/B NOR2X1_LOC_155/A 0.03fF
C75529 INVX1_LOC_37/A NAND2X1_LOC_637/Y 0.22fF
C75530 INVX1_LOC_11/A NOR2X1_LOC_751/Y 0.50fF
C75531 NAND2X1_LOC_579/A INVX1_LOC_41/Y 0.03fF
C75532 NOR2X1_LOC_454/Y NOR2X1_LOC_152/Y 0.07fF
C75533 NOR2X1_LOC_74/A INVX1_LOC_12/A 0.10fF
C75534 NOR2X1_LOC_439/a_36_216# NOR2X1_LOC_383/B 0.01fF
C75535 NOR2X1_LOC_220/A INVX1_LOC_23/A 0.11fF
C75536 NOR2X1_LOC_296/Y NOR2X1_LOC_791/B 0.00fF
C75537 NAND2X1_LOC_198/B INVX1_LOC_308/Y 0.01fF
C75538 INVX1_LOC_256/A NAND2X1_LOC_342/a_36_24# 0.01fF
C75539 INVX1_LOC_5/A NOR2X1_LOC_367/B 0.45fF
C75540 NOR2X1_LOC_454/Y INVX1_LOC_113/Y 0.05fF
C75541 NOR2X1_LOC_174/A NOR2X1_LOC_623/B 0.03fF
C75542 NOR2X1_LOC_218/A INVX1_LOC_130/Y 0.18fF
C75543 NOR2X1_LOC_794/B NOR2X1_LOC_703/B 0.01fF
C75544 INVX1_LOC_269/A INVX1_LOC_71/A 0.67fF
C75545 NOR2X1_LOC_602/B NOR2X1_LOC_536/A 0.02fF
C75546 INVX1_LOC_13/Y NAND2X1_LOC_465/Y 0.03fF
C75547 NOR2X1_LOC_160/B INVX1_LOC_72/A 0.70fF
C75548 NOR2X1_LOC_598/B NOR2X1_LOC_544/A 1.12fF
C75549 NOR2X1_LOC_186/Y NOR2X1_LOC_792/B 0.05fF
C75550 NOR2X1_LOC_9/Y INVX1_LOC_12/A 0.10fF
C75551 INVX1_LOC_58/A INVX1_LOC_22/A 17.65fF
C75552 NAND2X1_LOC_474/a_36_24# INVX1_LOC_26/A 0.00fF
C75553 NOR2X1_LOC_434/Y NOR2X1_LOC_175/A 0.01fF
C75554 NOR2X1_LOC_536/A INVX1_LOC_54/A 0.37fF
C75555 NAND2X1_LOC_787/A INVX1_LOC_25/Y 0.07fF
C75556 INVX1_LOC_279/A INVX1_LOC_270/A 0.10fF
C75557 NOR2X1_LOC_548/Y INVX1_LOC_23/A 0.16fF
C75558 INVX1_LOC_95/Y INVX1_LOC_63/A 0.34fF
C75559 INVX1_LOC_5/A INVX1_LOC_243/A 0.06fF
C75560 NOR2X1_LOC_815/Y NAND2X1_LOC_537/Y 0.00fF
C75561 INVX1_LOC_136/A NAND2X1_LOC_577/A 0.01fF
C75562 INVX1_LOC_278/A INVX1_LOC_56/Y 0.13fF
C75563 NAND2X1_LOC_573/Y NOR2X1_LOC_792/B 0.07fF
C75564 NAND2X1_LOC_286/a_36_24# INVX1_LOC_46/A 0.00fF
C75565 INVX1_LOC_194/A INVX1_LOC_239/A 0.01fF
C75566 NAND2X1_LOC_773/Y NOR2X1_LOC_309/Y 0.01fF
C75567 INVX1_LOC_83/A INVX1_LOC_57/A 0.14fF
C75568 INVX1_LOC_239/A NOR2X1_LOC_399/A 0.03fF
C75569 NAND2X1_LOC_195/Y INVX1_LOC_72/A -0.01fF
C75570 NAND2X1_LOC_569/B INVX1_LOC_16/A 0.09fF
C75571 NOR2X1_LOC_664/Y INVX1_LOC_14/A 0.10fF
C75572 NOR2X1_LOC_658/Y INVX1_LOC_159/A 0.03fF
C75573 NOR2X1_LOC_607/Y INVX1_LOC_292/A 0.01fF
C75574 NOR2X1_LOC_78/A NOR2X1_LOC_633/a_36_216# 0.00fF
C75575 NOR2X1_LOC_675/A INVX1_LOC_29/A 0.00fF
C75576 INVX1_LOC_315/Y NOR2X1_LOC_643/a_36_216# 0.00fF
C75577 INVX1_LOC_67/Y INVX1_LOC_94/Y 0.04fF
C75578 NAND2X1_LOC_585/a_36_24# INVX1_LOC_246/A 0.00fF
C75579 NOR2X1_LOC_662/A INVX1_LOC_46/A 0.01fF
C75580 INVX1_LOC_5/A NOR2X1_LOC_719/A 0.00fF
C75581 NOR2X1_LOC_435/a_36_216# NOR2X1_LOC_561/Y 0.01fF
C75582 NOR2X1_LOC_35/Y INVX1_LOC_125/A 0.19fF
C75583 NOR2X1_LOC_791/Y INVX1_LOC_25/Y 0.02fF
C75584 INVX1_LOC_249/A NOR2X1_LOC_717/Y 0.23fF
C75585 NOR2X1_LOC_859/a_36_216# NAND2X1_LOC_116/A 0.00fF
C75586 NOR2X1_LOC_844/Y INVX1_LOC_77/A 0.04fF
C75587 INVX1_LOC_136/A NAND2X1_LOC_656/A 0.32fF
C75588 INVX1_LOC_37/Y NAND2X1_LOC_489/Y 0.01fF
C75589 NAND2X1_LOC_725/A NOR2X1_LOC_298/Y 0.17fF
C75590 INVX1_LOC_5/A INVX1_LOC_7/A 0.05fF
C75591 NOR2X1_LOC_790/B NOR2X1_LOC_542/Y 0.00fF
C75592 NOR2X1_LOC_692/Y NOR2X1_LOC_485/Y 0.14fF
C75593 INVX1_LOC_182/Y INVX1_LOC_270/A 0.01fF
C75594 NOR2X1_LOC_13/Y INVX1_LOC_159/A 0.01fF
C75595 INPUT_0 INVX1_LOC_183/A 0.03fF
C75596 D_INPUT_3 NOR2X1_LOC_610/Y 0.01fF
C75597 INVX1_LOC_31/A NOR2X1_LOC_844/A 0.03fF
C75598 NOR2X1_LOC_510/Y NAND2X1_LOC_656/Y 0.16fF
C75599 INVX1_LOC_178/A NOR2X1_LOC_561/Y 0.10fF
C75600 NOR2X1_LOC_68/A INVX1_LOC_49/A 7.91fF
C75601 NOR2X1_LOC_777/B INVX1_LOC_117/A 0.03fF
C75602 INVX1_LOC_132/A NOR2X1_LOC_360/Y 0.07fF
C75603 NAND2X1_LOC_550/A NAND2X1_LOC_338/B 0.24fF
C75604 NAND2X1_LOC_600/a_36_24# INVX1_LOC_63/A 0.01fF
C75605 NOR2X1_LOC_160/B NOR2X1_LOC_537/Y 0.07fF
C75606 NOR2X1_LOC_160/B NAND2X1_LOC_338/B 0.56fF
C75607 INVX1_LOC_97/A INVX1_LOC_50/Y 0.03fF
C75608 INVX1_LOC_54/A NOR2X1_LOC_661/A 0.03fF
C75609 INVX1_LOC_255/Y NAND2X1_LOC_222/B 0.03fF
C75610 INVX1_LOC_161/Y NAND2X1_LOC_840/B 0.01fF
C75611 INVX1_LOC_34/A INVX1_LOC_72/Y 0.01fF
C75612 INVX1_LOC_98/A INVX1_LOC_26/A 0.25fF
C75613 NOR2X1_LOC_78/A NOR2X1_LOC_316/a_36_216# 0.00fF
C75614 INVX1_LOC_90/A INVX1_LOC_50/Y 0.50fF
C75615 NOR2X1_LOC_160/B NAND2X1_LOC_323/B 0.07fF
C75616 INVX1_LOC_284/Y NAND2X1_LOC_852/a_36_24# 0.00fF
C75617 NOR2X1_LOC_78/A INVX1_LOC_26/A 0.06fF
C75618 INVX1_LOC_2/Y INVX1_LOC_32/A 0.18fF
C75619 INVX1_LOC_58/A INVX1_LOC_100/A 0.13fF
C75620 INVX1_LOC_255/Y INVX1_LOC_11/A 0.03fF
C75621 NAND2X1_LOC_807/B NOR2X1_LOC_536/A 0.03fF
C75622 INVX1_LOC_225/A NOR2X1_LOC_360/Y 0.10fF
C75623 INVX1_LOC_77/A INVX1_LOC_113/Y 0.03fF
C75624 NAND2X1_LOC_639/A NOR2X1_LOC_48/B 0.06fF
C75625 INVX1_LOC_303/A NAND2X1_LOC_786/a_36_24# 0.01fF
C75626 NOR2X1_LOC_220/A INVX1_LOC_31/A 0.10fF
C75627 INVX1_LOC_14/A INVX1_LOC_234/A 0.68fF
C75628 INVX1_LOC_255/Y NAND2X1_LOC_381/Y 0.01fF
C75629 NOR2X1_LOC_722/Y INVX1_LOC_266/Y 0.02fF
C75630 NOR2X1_LOC_530/Y INVX1_LOC_16/A 0.02fF
C75631 NOR2X1_LOC_831/B INVX1_LOC_84/A 0.07fF
C75632 INVX1_LOC_256/A INVX1_LOC_215/A 0.10fF
C75633 NOR2X1_LOC_361/B NAND2X1_LOC_656/Y 0.61fF
C75634 INVX1_LOC_230/Y INVX1_LOC_232/A 0.48fF
C75635 INVX1_LOC_292/A NOR2X1_LOC_553/Y 0.01fF
C75636 NOR2X1_LOC_536/A NOR2X1_LOC_48/B 0.03fF
C75637 NOR2X1_LOC_208/Y NOR2X1_LOC_144/Y 0.04fF
C75638 INVX1_LOC_269/A NOR2X1_LOC_123/B 0.10fF
C75639 NOR2X1_LOC_45/B NOR2X1_LOC_654/A 0.02fF
C75640 INVX1_LOC_17/A NOR2X1_LOC_763/Y 0.39fF
C75641 INVX1_LOC_2/A NOR2X1_LOC_68/A 0.40fF
C75642 VDD INVX1_LOC_128/Y 0.28fF
C75643 INVX1_LOC_266/A INVX1_LOC_90/A 0.07fF
C75644 INVX1_LOC_9/A INVX1_LOC_42/A 0.20fF
C75645 NAND2X1_LOC_858/B NOR2X1_LOC_109/Y 0.06fF
C75646 NAND2X1_LOC_348/A INVX1_LOC_50/Y 0.07fF
C75647 INVX1_LOC_25/A INVX1_LOC_91/A 0.10fF
C75648 NOR2X1_LOC_791/Y INVX1_LOC_75/A 0.03fF
C75649 NOR2X1_LOC_139/Y NOR2X1_LOC_125/Y 0.46fF
C75650 INVX1_LOC_30/A INVX1_LOC_25/Y 0.13fF
C75651 NOR2X1_LOC_226/A NOR2X1_LOC_68/A 0.10fF
C75652 INVX1_LOC_11/A NOR2X1_LOC_71/Y 0.07fF
C75653 NOR2X1_LOC_237/a_36_216# NOR2X1_LOC_315/Y 0.00fF
C75654 NAND2X1_LOC_552/A NOR2X1_LOC_167/Y 0.02fF
C75655 INVX1_LOC_208/A INVX1_LOC_72/A 0.07fF
C75656 NAND2X1_LOC_650/B NOR2X1_LOC_301/A 0.07fF
C75657 NOR2X1_LOC_590/Y INVX1_LOC_311/A 0.14fF
C75658 INVX1_LOC_226/Y NOR2X1_LOC_791/A -0.00fF
C75659 INVX1_LOC_34/A NAND2X1_LOC_811/Y 0.03fF
C75660 NOR2X1_LOC_91/Y NAND2X1_LOC_862/A 0.03fF
C75661 NOR2X1_LOC_203/Y INVX1_LOC_94/A 0.01fF
C75662 NAND2X1_LOC_725/B NAND2X1_LOC_560/A 0.03fF
C75663 INVX1_LOC_14/A NOR2X1_LOC_19/B 0.20fF
C75664 NAND2X1_LOC_214/B INVX1_LOC_48/A 0.21fF
C75665 NAND2X1_LOC_30/Y NOR2X1_LOC_163/A 0.01fF
C75666 NAND2X1_LOC_538/Y INVX1_LOC_28/A 0.09fF
C75667 INVX1_LOC_11/A NOR2X1_LOC_644/A 0.03fF
C75668 INVX1_LOC_204/A INVX1_LOC_115/A 0.01fF
C75669 NAND2X1_LOC_537/Y NAND2X1_LOC_680/a_36_24# 0.01fF
C75670 INVX1_LOC_124/Y INVX1_LOC_10/A 0.14fF
C75671 NAND2X1_LOC_456/Y INVX1_LOC_19/A 0.06fF
C75672 INVX1_LOC_17/Y INVX1_LOC_20/A 0.06fF
C75673 INVX1_LOC_178/A NOR2X1_LOC_167/Y 0.11fF
C75674 INVX1_LOC_23/A NAND2X1_LOC_469/B 0.07fF
C75675 INVX1_LOC_36/A INVX1_LOC_279/A 0.07fF
C75676 INVX1_LOC_251/Y NOR2X1_LOC_716/B 0.07fF
C75677 NOR2X1_LOC_338/Y INVX1_LOC_22/A 0.03fF
C75678 NAND2X1_LOC_726/Y NAND2X1_LOC_731/Y 0.08fF
C75679 INVX1_LOC_225/A NOR2X1_LOC_792/B 0.00fF
C75680 NOR2X1_LOC_389/A INVX1_LOC_313/A 0.01fF
C75681 NOR2X1_LOC_516/B INVX1_LOC_198/Y 0.01fF
C75682 VDD NOR2X1_LOC_727/B 0.02fF
C75683 NOR2X1_LOC_250/A INVX1_LOC_28/A 0.07fF
C75684 NOR2X1_LOC_160/B INVX1_LOC_313/Y 0.03fF
C75685 NOR2X1_LOC_307/B INVX1_LOC_77/A 0.03fF
C75686 INVX1_LOC_45/A NOR2X1_LOC_97/a_36_216# 0.00fF
C75687 D_GATE_741 INVX1_LOC_311/Y 0.00fF
C75688 INVX1_LOC_34/A INVX1_LOC_266/Y 0.10fF
C75689 NOR2X1_LOC_98/a_36_216# INVX1_LOC_26/A 0.01fF
C75690 NOR2X1_LOC_381/Y NAND2X1_LOC_348/A 0.12fF
C75691 NAND2X1_LOC_288/A NAND2X1_LOC_288/a_36_24# 0.01fF
C75692 INVX1_LOC_27/A INVX1_LOC_48/A 1.94fF
C75693 NOR2X1_LOC_598/B NOR2X1_LOC_683/Y 0.01fF
C75694 NAND2X1_LOC_736/Y NAND2X1_LOC_722/A 0.16fF
C75695 INVX1_LOC_57/A INVX1_LOC_46/A 0.17fF
C75696 INVX1_LOC_217/Y NAND2X1_LOC_570/Y 0.04fF
C75697 INVX1_LOC_244/Y INVX1_LOC_290/A 0.02fF
C75698 NAND2X1_LOC_803/B NOR2X1_LOC_171/Y 0.04fF
C75699 NOR2X1_LOC_843/B INVX1_LOC_117/A 0.07fF
C75700 INVX1_LOC_78/A INVX1_LOC_9/A 0.15fF
C75701 NOR2X1_LOC_576/B NOR2X1_LOC_599/A 0.03fF
C75702 NOR2X1_LOC_98/A INVX1_LOC_57/A 0.00fF
C75703 D_INPUT_1 NOR2X1_LOC_137/Y 0.07fF
C75704 INVX1_LOC_88/A INVX1_LOC_144/A 0.09fF
C75705 INVX1_LOC_110/Y NAND2X1_LOC_508/A 0.07fF
C75706 NOR2X1_LOC_612/a_36_216# NOR2X1_LOC_557/Y 0.00fF
C75707 INVX1_LOC_224/Y INVX1_LOC_12/Y 0.03fF
C75708 INVX1_LOC_49/Y INVX1_LOC_19/A 0.03fF
C75709 NAND2X1_LOC_470/B INVX1_LOC_54/A 0.99fF
C75710 INVX1_LOC_32/A NOR2X1_LOC_608/Y -0.01fF
C75711 NOR2X1_LOC_457/A INVX1_LOC_75/A 0.12fF
C75712 NOR2X1_LOC_662/A NOR2X1_LOC_671/Y 0.03fF
C75713 INVX1_LOC_287/A INVX1_LOC_117/A 0.00fF
C75714 NOR2X1_LOC_468/Y INVX1_LOC_6/A 0.21fF
C75715 INVX1_LOC_90/A NOR2X1_LOC_248/Y 0.01fF
C75716 INVX1_LOC_200/A NOR2X1_LOC_74/A 0.00fF
C75717 INPUT_3 INVX1_LOC_82/Y 0.12fF
C75718 INVX1_LOC_36/A NAND2X1_LOC_815/a_36_24# 0.00fF
C75719 VDD NOR2X1_LOC_717/A 1.43fF
C75720 INVX1_LOC_255/Y NOR2X1_LOC_474/A 0.00fF
C75721 NOR2X1_LOC_389/B NOR2X1_LOC_248/Y 0.03fF
C75722 NAND2X1_LOC_803/B NOR2X1_LOC_594/Y 0.03fF
C75723 INVX1_LOC_206/A INVX1_LOC_111/Y 0.04fF
C75724 NAND2X1_LOC_231/Y INVX1_LOC_266/Y 0.00fF
C75725 NOR2X1_LOC_65/B INVX1_LOC_9/A 0.00fF
C75726 NOR2X1_LOC_68/A INPUT_1 0.08fF
C75727 INVX1_LOC_5/A INVX1_LOC_76/A 3.95fF
C75728 INVX1_LOC_1/A INVX1_LOC_91/A 0.10fF
C75729 NOR2X1_LOC_439/B INVX1_LOC_30/A 0.04fF
C75730 NOR2X1_LOC_9/a_36_216# INVX1_LOC_306/Y 0.01fF
C75731 INVX1_LOC_116/A INVX1_LOC_171/A 0.01fF
C75732 INVX1_LOC_20/A NOR2X1_LOC_406/A 0.00fF
C75733 INVX1_LOC_136/A NOR2X1_LOC_329/B 0.12fF
C75734 INVX1_LOC_30/A INVX1_LOC_75/A 0.24fF
C75735 NOR2X1_LOC_214/B INVX1_LOC_71/A 2.75fF
C75736 INVX1_LOC_30/Y NOR2X1_LOC_392/B 0.10fF
C75737 VDD NOR2X1_LOC_649/Y 0.15fF
C75738 INVX1_LOC_178/A INVX1_LOC_76/A 0.10fF
C75739 INVX1_LOC_90/A NAND2X1_LOC_187/a_36_24# 0.00fF
C75740 NOR2X1_LOC_389/A INVX1_LOC_6/A 0.03fF
C75741 INVX1_LOC_16/A NOR2X1_LOC_709/A 0.10fF
C75742 INVX1_LOC_217/Y INVX1_LOC_234/A -0.01fF
C75743 NOR2X1_LOC_632/Y INVX1_LOC_85/A 0.91fF
C75744 INVX1_LOC_13/A INVX1_LOC_60/Y 0.02fF
C75745 NAND2X1_LOC_474/Y NOR2X1_LOC_266/B 0.02fF
C75746 NOR2X1_LOC_75/Y NOR2X1_LOC_45/B 0.04fF
C75747 NOR2X1_LOC_516/B NOR2X1_LOC_537/Y 0.03fF
C75748 NAND2X1_LOC_199/B INVX1_LOC_6/A 0.03fF
C75749 NOR2X1_LOC_516/B NAND2X1_LOC_338/B 0.10fF
C75750 NOR2X1_LOC_794/B INVX1_LOC_91/A 0.02fF
C75751 NAND2X1_LOC_493/Y INVX1_LOC_20/A 0.46fF
C75752 INVX1_LOC_49/A NOR2X1_LOC_163/A 0.02fF
C75753 INVX1_LOC_271/Y INVX1_LOC_63/A 0.01fF
C75754 D_INPUT_3 NAND2X1_LOC_473/A 1.03fF
C75755 INVX1_LOC_58/A NOR2X1_LOC_88/A 0.05fF
C75756 INVX1_LOC_53/A INVX1_LOC_274/A 0.53fF
C75757 NOR2X1_LOC_703/B NOR2X1_LOC_188/A 0.02fF
C75758 INVX1_LOC_256/A INVX1_LOC_95/A 0.10fF
C75759 INVX1_LOC_18/A NOR2X1_LOC_589/Y 0.06fF
C75760 NOR2X1_LOC_644/A NOR2X1_LOC_593/Y 0.03fF
C75761 NOR2X1_LOC_809/a_36_216# INVX1_LOC_196/A 0.17fF
C75762 NOR2X1_LOC_619/A INVX1_LOC_218/A 0.17fF
C75763 NOR2X1_LOC_785/Y NOR2X1_LOC_168/B 0.00fF
C75764 NOR2X1_LOC_384/Y INVX1_LOC_309/A -0.00fF
C75765 NAND2X1_LOC_656/Y INVX1_LOC_177/A 0.03fF
C75766 NOR2X1_LOC_52/B NOR2X1_LOC_71/Y 0.15fF
C75767 NOR2X1_LOC_241/A INVX1_LOC_143/Y 0.01fF
C75768 INVX1_LOC_161/Y NOR2X1_LOC_137/a_36_216# 0.01fF
C75769 INVX1_LOC_107/A INVX1_LOC_6/A 0.01fF
C75770 INVX1_LOC_35/A INVX1_LOC_75/Y 0.01fF
C75771 INVX1_LOC_17/A NAND2X1_LOC_650/B 0.07fF
C75772 INVX1_LOC_90/A NOR2X1_LOC_6/B 0.03fF
C75773 INVX1_LOC_172/Y NAND2X1_LOC_735/B 0.05fF
C75774 NOR2X1_LOC_773/Y NOR2X1_LOC_561/Y 0.01fF
C75775 NOR2X1_LOC_620/Y INVX1_LOC_31/Y 0.07fF
C75776 NAND2X1_LOC_337/B INVX1_LOC_76/A 0.10fF
C75777 INVX1_LOC_217/Y NOR2X1_LOC_19/B 0.05fF
C75778 NAND2X1_LOC_430/B INVX1_LOC_15/A 0.01fF
C75779 INVX1_LOC_271/A NOR2X1_LOC_127/Y 0.01fF
C75780 INVX1_LOC_3/A NAND2X1_LOC_215/A 0.07fF
C75781 NOR2X1_LOC_384/Y INVX1_LOC_91/A 0.03fF
C75782 NOR2X1_LOC_596/A INVX1_LOC_6/A 0.06fF
C75783 NOR2X1_LOC_816/A INVX1_LOC_76/A 0.19fF
C75784 INVX1_LOC_165/A NAND2X1_LOC_254/Y 0.03fF
C75785 NOR2X1_LOC_103/Y INVX1_LOC_12/Y 0.10fF
C75786 INVX1_LOC_266/A INVX1_LOC_38/A 0.07fF
C75787 NOR2X1_LOC_68/Y INVX1_LOC_57/A 0.13fF
C75788 INPUT_3 INVX1_LOC_2/Y 0.03fF
C75789 INVX1_LOC_34/A INVX1_LOC_42/Y 0.00fF
C75790 NOR2X1_LOC_97/A INVX1_LOC_33/A 0.20fF
C75791 NAND2X1_LOC_341/A NOR2X1_LOC_366/Y 0.02fF
C75792 NAND2X1_LOC_727/Y INVX1_LOC_10/A 0.07fF
C75793 INVX1_LOC_226/Y D_INPUT_0 0.04fF
C75794 NAND2X1_LOC_504/a_36_24# INVX1_LOC_210/A 0.00fF
C75795 INVX1_LOC_58/A INVX1_LOC_186/Y 0.10fF
C75796 NOR2X1_LOC_329/B NOR2X1_LOC_111/a_36_216# 0.01fF
C75797 NAND2X1_LOC_348/A NOR2X1_LOC_6/B 0.02fF
C75798 NAND2X1_LOC_338/B NOR2X1_LOC_756/a_36_216# 0.00fF
C75799 INPUT_0 NAND2X1_LOC_811/Y 0.03fF
C75800 NOR2X1_LOC_360/Y NAND2X1_LOC_642/Y 0.03fF
C75801 NAND2X1_LOC_660/Y INVX1_LOC_10/A 0.07fF
C75802 NAND2X1_LOC_162/B NOR2X1_LOC_45/B 0.02fF
C75803 NOR2X1_LOC_61/B INVX1_LOC_152/A 0.03fF
C75804 INVX1_LOC_31/A NOR2X1_LOC_447/B 0.01fF
C75805 NOR2X1_LOC_89/A NOR2X1_LOC_39/Y 0.03fF
C75806 INVX1_LOC_208/A INVX1_LOC_313/Y 0.04fF
C75807 NAND2X1_LOC_254/Y NOR2X1_LOC_693/Y 0.02fF
C75808 NAND2X1_LOC_579/A INVX1_LOC_185/A 0.05fF
C75809 INVX1_LOC_233/A NOR2X1_LOC_662/A 0.02fF
C75810 NOR2X1_LOC_658/Y NOR2X1_LOC_69/a_36_216# 0.00fF
C75811 NOR2X1_LOC_309/Y NAND2X1_LOC_858/B 0.17fF
C75812 NOR2X1_LOC_658/Y VDD 0.69fF
C75813 NAND2X1_LOC_842/a_36_24# NAND2X1_LOC_850/Y 0.00fF
C75814 NAND2X1_LOC_717/Y NAND2X1_LOC_863/A 0.03fF
C75815 INVX1_LOC_58/A INVX1_LOC_261/A 0.02fF
C75816 INVX1_LOC_47/A INVX1_LOC_1/Y 0.78fF
C75817 INVX1_LOC_135/A NOR2X1_LOC_391/A 0.02fF
C75818 INVX1_LOC_2/A INVX1_LOC_147/A 0.03fF
C75819 INVX1_LOC_72/A NAND2X1_LOC_211/Y 0.07fF
C75820 INVX1_LOC_7/A NOR2X1_LOC_332/A 0.04fF
C75821 INVX1_LOC_172/A NAND2X1_LOC_623/B 0.02fF
C75822 INVX1_LOC_24/A NOR2X1_LOC_631/B 0.07fF
C75823 NOR2X1_LOC_716/B NOR2X1_LOC_45/B 0.08fF
C75824 INVX1_LOC_2/A NOR2X1_LOC_2/Y 0.01fF
C75825 NOR2X1_LOC_599/a_36_216# INVX1_LOC_46/A 0.02fF
C75826 INVX1_LOC_30/Y INVX1_LOC_90/A 1.38fF
C75827 INVX1_LOC_45/A INVX1_LOC_12/Y 0.01fF
C75828 NOR2X1_LOC_13/Y NOR2X1_LOC_56/Y 0.10fF
C75829 INVX1_LOC_71/A NOR2X1_LOC_275/A 0.01fF
C75830 NOR2X1_LOC_226/A INVX1_LOC_147/A 0.07fF
C75831 NOR2X1_LOC_518/Y VDD 0.12fF
C75832 INVX1_LOC_256/A INVX1_LOC_54/A 0.03fF
C75833 NOR2X1_LOC_441/Y NOR2X1_LOC_536/A 0.04fF
C75834 NOR2X1_LOC_785/Y INVX1_LOC_132/Y 0.33fF
C75835 INVX1_LOC_27/A NOR2X1_LOC_127/Y 0.07fF
C75836 INVX1_LOC_35/A NAND2X1_LOC_74/B 0.09fF
C75837 INVX1_LOC_88/A NOR2X1_LOC_155/A 0.03fF
C75838 INVX1_LOC_14/A NOR2X1_LOC_216/B 1.98fF
C75839 NAND2X1_LOC_363/B NAND2X1_LOC_291/B 0.15fF
C75840 INVX1_LOC_221/A INVX1_LOC_91/A 0.02fF
C75841 INVX1_LOC_24/A NOR2X1_LOC_681/Y 0.40fF
C75842 INVX1_LOC_18/A INVX1_LOC_117/A 0.30fF
C75843 NOR2X1_LOC_495/Y INVX1_LOC_20/A 0.00fF
C75844 INVX1_LOC_24/A INVX1_LOC_37/A 0.19fF
C75845 NOR2X1_LOC_13/Y VDD 1.04fF
C75846 INVX1_LOC_205/Y NOR2X1_LOC_814/A 0.03fF
C75847 NOR2X1_LOC_773/Y NOR2X1_LOC_167/Y 0.02fF
C75848 INVX1_LOC_24/A NOR2X1_LOC_231/A 0.02fF
C75849 INVX1_LOC_1/A NOR2X1_LOC_179/Y 0.03fF
C75850 NOR2X1_LOC_216/a_36_216# INVX1_LOC_10/A 0.00fF
C75851 NOR2X1_LOC_561/Y INVX1_LOC_140/A 0.10fF
C75852 INVX1_LOC_315/Y NOR2X1_LOC_537/Y 0.03fF
C75853 NAND2X1_LOC_368/a_36_24# NAND2X1_LOC_472/Y 0.00fF
C75854 NOR2X1_LOC_389/A INVX1_LOC_131/Y 0.11fF
C75855 NOR2X1_LOC_298/Y NAND2X1_LOC_560/A 0.05fF
C75856 NOR2X1_LOC_137/A NOR2X1_LOC_772/A 0.01fF
C75857 INVX1_LOC_71/A INVX1_LOC_12/Y 0.48fF
C75858 INVX1_LOC_299/A NOR2X1_LOC_814/A 0.23fF
C75859 INVX1_LOC_28/A NOR2X1_LOC_106/A 0.05fF
C75860 NAND2X1_LOC_660/A NAND2X1_LOC_655/A 0.01fF
C75861 NAND2X1_LOC_364/Y VDD 0.01fF
C75862 NOR2X1_LOC_416/A NOR2X1_LOC_38/B 0.08fF
C75863 INVX1_LOC_229/Y NOR2X1_LOC_409/Y 2.59fF
C75864 NOR2X1_LOC_554/B INVX1_LOC_9/A 0.89fF
C75865 NOR2X1_LOC_168/B INVX1_LOC_65/A 0.05fF
C75866 INVX1_LOC_57/A NOR2X1_LOC_282/a_36_216# 0.00fF
C75867 NAND2X1_LOC_356/a_36_24# INVX1_LOC_38/A 0.01fF
C75868 NOR2X1_LOC_538/B NOR2X1_LOC_814/A 0.02fF
C75869 NAND2X1_LOC_175/B VDD 0.31fF
C75870 NOR2X1_LOC_68/A INVX1_LOC_118/A 0.07fF
C75871 INVX1_LOC_167/A INVX1_LOC_242/A 0.03fF
C75872 INVX1_LOC_219/Y INVX1_LOC_20/A 0.02fF
C75873 INVX1_LOC_33/A NOR2X1_LOC_168/a_36_216# 0.00fF
C75874 INVX1_LOC_256/Y NOR2X1_LOC_123/a_36_216# 0.01fF
C75875 NAND2X1_LOC_842/B NAND2X1_LOC_850/A 0.08fF
C75876 D_INPUT_3 NOR2X1_LOC_143/a_36_216# 0.00fF
C75877 INVX1_LOC_24/A NAND2X1_LOC_629/a_36_24# 0.00fF
C75878 NOR2X1_LOC_440/Y INVX1_LOC_286/A 0.01fF
C75879 NAND2X1_LOC_656/Y INVX1_LOC_285/Y 0.10fF
C75880 NOR2X1_LOC_562/a_36_216# INVX1_LOC_44/A 0.00fF
C75881 NOR2X1_LOC_152/Y INVX1_LOC_9/A 0.01fF
C75882 NOR2X1_LOC_504/Y VDD 0.02fF
C75883 INVX1_LOC_28/A NAND2X1_LOC_863/A 0.17fF
C75884 NAND2X1_LOC_9/Y NOR2X1_LOC_55/a_36_216# 0.00fF
C75885 INVX1_LOC_2/A NOR2X1_LOC_364/a_36_216# 0.00fF
C75886 INVX1_LOC_161/Y INVX1_LOC_49/Y 0.04fF
C75887 NOR2X1_LOC_142/Y NOR2X1_LOC_536/A 0.01fF
C75888 NOR2X1_LOC_134/Y NAND2X1_LOC_768/Y 0.05fF
C75889 INVX1_LOC_164/A INVX1_LOC_98/A 0.32fF
C75890 NOR2X1_LOC_441/Y NOR2X1_LOC_661/A 0.03fF
C75891 NOR2X1_LOC_773/Y INVX1_LOC_76/A 0.19fF
C75892 INVX1_LOC_95/Y INVX1_LOC_1/Y 0.03fF
C75893 INVX1_LOC_164/A NOR2X1_LOC_78/A 0.01fF
C75894 INVX1_LOC_143/A INVX1_LOC_37/A 0.21fF
C75895 INVX1_LOC_256/Y VDD 0.60fF
C75896 INVX1_LOC_17/A NOR2X1_LOC_67/Y 0.04fF
C75897 INVX1_LOC_143/A NOR2X1_LOC_231/A 0.01fF
C75898 NOR2X1_LOC_510/Y INVX1_LOC_128/Y 0.02fF
C75899 NAND2X1_LOC_841/A INVX1_LOC_139/A 0.12fF
C75900 NOR2X1_LOC_6/B INVX1_LOC_38/A 0.03fF
C75901 INVX1_LOC_255/Y INVX1_LOC_74/A 0.02fF
C75902 INVX1_LOC_245/Y INVX1_LOC_12/A 0.03fF
C75903 INVX1_LOC_159/A NOR2X1_LOC_697/Y 0.00fF
C75904 NOR2X1_LOC_210/B NAND2X1_LOC_220/a_36_24# 0.00fF
C75905 INVX1_LOC_41/A NOR2X1_LOC_612/Y 0.01fF
C75906 NOR2X1_LOC_470/A INVX1_LOC_199/Y 0.09fF
C75907 NAND2X1_LOC_9/Y INVX1_LOC_57/A 0.58fF
C75908 NOR2X1_LOC_384/Y INVX1_LOC_203/A 0.10fF
C75909 INVX1_LOC_90/A INVX1_LOC_96/A 0.03fF
C75910 NOR2X1_LOC_222/a_36_216# NOR2X1_LOC_357/Y 0.01fF
C75911 INVX1_LOC_233/A INVX1_LOC_57/A 0.16fF
C75912 INVX1_LOC_33/A NOR2X1_LOC_809/B 0.02fF
C75913 NOR2X1_LOC_19/B INVX1_LOC_48/A 0.21fF
C75914 NOR2X1_LOC_146/Y VDD 0.15fF
C75915 INVX1_LOC_40/A INVX1_LOC_129/Y 0.01fF
C75916 NOR2X1_LOC_655/B NOR2X1_LOC_536/A 0.05fF
C75917 NOR2X1_LOC_142/Y NAND2X1_LOC_93/B 0.07fF
C75918 NOR2X1_LOC_32/B NOR2X1_LOC_629/A 0.04fF
C75919 NOR2X1_LOC_717/B INVX1_LOC_247/A 0.16fF
C75920 NOR2X1_LOC_92/Y NOR2X1_LOC_409/B 1.59fF
C75921 NOR2X1_LOC_613/a_36_216# NOR2X1_LOC_693/Y 0.01fF
C75922 INVX1_LOC_225/A NOR2X1_LOC_79/Y 0.02fF
C75923 NOR2X1_LOC_181/Y INVX1_LOC_179/A 0.00fF
C75924 INVX1_LOC_10/A NOR2X1_LOC_266/B 0.11fF
C75925 NOR2X1_LOC_68/A NAND2X1_LOC_63/Y 0.03fF
C75926 NOR2X1_LOC_785/A INVX1_LOC_15/A 0.03fF
C75927 NOR2X1_LOC_32/B NAND2X1_LOC_624/B 0.07fF
C75928 INVX1_LOC_35/A NOR2X1_LOC_660/Y 0.43fF
C75929 NOR2X1_LOC_577/Y NAND2X1_LOC_475/Y 0.10fF
C75930 NOR2X1_LOC_665/A NAND2X1_LOC_472/Y 0.07fF
C75931 NOR2X1_LOC_655/B NOR2X1_LOC_655/Y 0.00fF
C75932 NOR2X1_LOC_798/A INVX1_LOC_57/A 0.05fF
C75933 INVX1_LOC_27/A NOR2X1_LOC_383/B 0.15fF
C75934 NAND2X1_LOC_357/B NOR2X1_LOC_88/Y 0.07fF
C75935 NAND2X1_LOC_303/Y NOR2X1_LOC_829/A 0.01fF
C75936 NOR2X1_LOC_130/A INVX1_LOC_37/A 0.02fF
C75937 INVX1_LOC_162/A INVX1_LOC_285/A 0.03fF
C75938 NOR2X1_LOC_337/Y NOR2X1_LOC_337/A 0.03fF
C75939 NAND2X1_LOC_803/B INVX1_LOC_94/Y 0.24fF
C75940 NOR2X1_LOC_655/B NAND2X1_LOC_93/B 0.03fF
C75941 INVX1_LOC_171/Y INVX1_LOC_29/Y 0.00fF
C75942 INVX1_LOC_81/Y INVX1_LOC_15/A 0.01fF
C75943 NAND2X1_LOC_114/B INVX1_LOC_4/Y 0.13fF
C75944 INVX1_LOC_244/Y INVX1_LOC_261/Y 0.02fF
C75945 NAND2X1_LOC_30/Y NOR2X1_LOC_36/A 0.60fF
C75946 NAND2X1_LOC_350/A NAND2X1_LOC_470/B 0.02fF
C75947 NAND2X1_LOC_703/Y INVX1_LOC_57/A 0.08fF
C75948 INVX1_LOC_278/A NAND2X1_LOC_169/Y 0.01fF
C75949 NOR2X1_LOC_238/a_36_216# NOR2X1_LOC_89/A -0.02fF
C75950 NOR2X1_LOC_246/A NOR2X1_LOC_111/A 0.02fF
C75951 NOR2X1_LOC_188/A INVX1_LOC_91/A 0.19fF
C75952 INVX1_LOC_100/Y INVX1_LOC_6/A 0.01fF
C75953 NOR2X1_LOC_123/B INVX1_LOC_12/Y 0.10fF
C75954 NOR2X1_LOC_778/B INVX1_LOC_179/A 0.00fF
C75955 NOR2X1_LOC_545/A NAND2X1_LOC_63/Y 0.05fF
C75956 NOR2X1_LOC_391/A INVX1_LOC_280/A 0.01fF
C75957 NAND2X1_LOC_348/A NOR2X1_LOC_124/A 0.01fF
C75958 NOR2X1_LOC_548/B INVX1_LOC_91/A 0.10fF
C75959 NOR2X1_LOC_590/A INVX1_LOC_94/Y 0.07fF
C75960 NOR2X1_LOC_736/Y NOR2X1_LOC_357/Y 0.10fF
C75961 NOR2X1_LOC_151/Y INVX1_LOC_247/A 0.01fF
C75962 NAND2X1_LOC_357/B INVX1_LOC_84/A 0.08fF
C75963 INVX1_LOC_224/A NOR2X1_LOC_39/Y 0.06fF
C75964 INVX1_LOC_18/A INVX1_LOC_3/Y 0.10fF
C75965 INVX1_LOC_140/A INVX1_LOC_76/A 0.19fF
C75966 NOR2X1_LOC_99/B NOR2X1_LOC_536/A 0.09fF
C75967 INVX1_LOC_36/A NOR2X1_LOC_38/B 0.03fF
C75968 NOR2X1_LOC_67/A INVX1_LOC_123/Y 0.04fF
C75969 INVX1_LOC_34/A INVX1_LOC_19/A 0.11fF
C75970 NOR2X1_LOC_68/A INVX1_LOC_257/A 0.01fF
C75971 NAND2X1_LOC_7/Y INVX1_LOC_106/Y 0.13fF
C75972 NAND2X1_LOC_555/Y NOR2X1_LOC_415/Y 0.02fF
C75973 INVX1_LOC_226/Y INVX1_LOC_46/Y 0.02fF
C75974 INVX1_LOC_34/A NOR2X1_LOC_11/Y 0.03fF
C75975 INVX1_LOC_5/A NOR2X1_LOC_34/B 0.01fF
C75976 INVX1_LOC_48/A NAND2X1_LOC_813/a_36_24# 0.00fF
C75977 NOR2X1_LOC_781/B NAND2X1_LOC_637/Y 0.02fF
C75978 NOR2X1_LOC_717/B NOR2X1_LOC_499/B 0.00fF
C75979 INVX1_LOC_88/A NOR2X1_LOC_125/Y 0.01fF
C75980 NOR2X1_LOC_753/Y INVX1_LOC_102/A 0.07fF
C75981 INVX1_LOC_310/A NOR2X1_LOC_814/A 0.19fF
C75982 NOR2X1_LOC_655/B NOR2X1_LOC_649/B 0.02fF
C75983 NOR2X1_LOC_655/B INVX1_LOC_3/A 0.10fF
C75984 INVX1_LOC_90/A NOR2X1_LOC_684/Y 0.10fF
C75985 NOR2X1_LOC_169/B INVX1_LOC_78/A 0.01fF
C75986 NOR2X1_LOC_690/A NOR2X1_LOC_824/a_36_216# 0.01fF
C75987 NAND2X1_LOC_549/B INVX1_LOC_84/A 0.02fF
C75988 INVX1_LOC_135/A NOR2X1_LOC_629/Y 0.01fF
C75989 INVX1_LOC_64/A NAND2X1_LOC_493/Y 0.05fF
C75990 NAND2X1_LOC_569/B INVX1_LOC_48/Y 0.09fF
C75991 INVX1_LOC_230/Y INVX1_LOC_112/Y 0.05fF
C75992 NOR2X1_LOC_197/A NOR2X1_LOC_748/A 0.02fF
C75993 NAND2X1_LOC_569/A INVX1_LOC_284/A 0.01fF
C75994 NOR2X1_LOC_43/Y INVX1_LOC_91/A 0.03fF
C75995 INVX1_LOC_6/A NAND2X1_LOC_469/B 0.96fF
C75996 NAND2X1_LOC_492/a_36_24# INVX1_LOC_9/A 0.01fF
C75997 INVX1_LOC_224/Y NOR2X1_LOC_160/B 0.13fF
C75998 NOR2X1_LOC_112/B INVX1_LOC_37/A 0.15fF
C75999 INVX1_LOC_170/A INVX1_LOC_26/A 0.01fF
C76000 INVX1_LOC_103/A NOR2X1_LOC_678/A 0.28fF
C76001 VDD NOR2X1_LOC_337/A 0.12fF
C76002 NAND2X1_LOC_231/Y INVX1_LOC_19/A 0.14fF
C76003 NAND2X1_LOC_21/Y NAND2X1_LOC_430/B 0.09fF
C76004 NOR2X1_LOC_717/B NOR2X1_LOC_676/Y 0.00fF
C76005 NOR2X1_LOC_130/A NOR2X1_LOC_743/Y 0.03fF
C76006 NOR2X1_LOC_322/Y INVX1_LOC_33/Y 0.01fF
C76007 NAND2X1_LOC_451/Y NOR2X1_LOC_48/Y 0.01fF
C76008 INVX1_LOC_16/A INVX1_LOC_294/A 0.02fF
C76009 INVX1_LOC_24/A NAND2X1_LOC_72/B 0.03fF
C76010 NAND2X1_LOC_715/B INVX1_LOC_88/A 0.48fF
C76011 INVX1_LOC_35/A NOR2X1_LOC_307/A 0.03fF
C76012 NOR2X1_LOC_433/A INVX1_LOC_21/Y 0.03fF
C76013 NOR2X1_LOC_121/A INVX1_LOC_293/Y 0.02fF
C76014 NAND2X1_LOC_338/B NAND2X1_LOC_207/B 0.03fF
C76015 D_INPUT_0 NOR2X1_LOC_445/B 0.07fF
C76016 NAND2X1_LOC_361/Y INVX1_LOC_4/A 0.07fF
C76017 INVX1_LOC_93/Y INVX1_LOC_95/Y 0.15fF
C76018 NOR2X1_LOC_828/A NOR2X1_LOC_676/Y 0.04fF
C76019 INVX1_LOC_93/A INVX1_LOC_14/A 1.40fF
C76020 NOR2X1_LOC_151/Y NOR2X1_LOC_499/B 0.01fF
C76021 NOR2X1_LOC_181/A INVX1_LOC_247/A 0.04fF
C76022 NOR2X1_LOC_644/A NOR2X1_LOC_858/a_36_216# 0.00fF
C76023 NOR2X1_LOC_763/Y NOR2X1_LOC_430/Y 0.06fF
C76024 NOR2X1_LOC_45/B NAND2X1_LOC_633/Y 0.20fF
C76025 INVX1_LOC_279/A INVX1_LOC_63/A 0.07fF
C76026 NAND2X1_LOC_357/B INVX1_LOC_15/A 0.07fF
C76027 NOR2X1_LOC_121/A NAND2X1_LOC_74/B 0.01fF
C76028 NOR2X1_LOC_598/B NOR2X1_LOC_500/B 0.25fF
C76029 NOR2X1_LOC_99/B INVX1_LOC_3/A 0.16fF
C76030 INVX1_LOC_58/A INVX1_LOC_18/A 2.39fF
C76031 NOR2X1_LOC_382/Y NOR2X1_LOC_392/Y 0.02fF
C76032 INVX1_LOC_66/A NOR2X1_LOC_814/A 0.02fF
C76033 NAND2X1_LOC_354/B INVX1_LOC_94/Y 0.00fF
C76034 INVX1_LOC_58/A NAND2X1_LOC_728/Y 0.07fF
C76035 INVX1_LOC_132/A INVX1_LOC_26/A 0.07fF
C76036 INVX1_LOC_34/Y INVX1_LOC_3/Y 1.19fF
C76037 INVX1_LOC_56/A NOR2X1_LOC_76/B 0.00fF
C76038 NOR2X1_LOC_151/Y NOR2X1_LOC_676/Y 0.03fF
C76039 NAND2X1_LOC_303/Y NAND2X1_LOC_537/Y 0.46fF
C76040 INVX1_LOC_249/A NOR2X1_LOC_383/B 0.03fF
C76041 NOR2X1_LOC_726/Y INVX1_LOC_213/A 0.04fF
C76042 INVX1_LOC_35/A INVX1_LOC_136/A 0.16fF
C76043 NOR2X1_LOC_6/B NAND2X1_LOC_223/A 0.03fF
C76044 NAND2X1_LOC_660/Y INVX1_LOC_12/A 0.08fF
C76045 NOR2X1_LOC_577/Y NOR2X1_LOC_135/a_36_216# 0.00fF
C76046 INVX1_LOC_215/A NOR2X1_LOC_89/A 0.07fF
C76047 INVX1_LOC_58/A NAND2X1_LOC_711/B 0.14fF
C76048 INVX1_LOC_1/A NOR2X1_LOC_739/Y 0.03fF
C76049 INVX1_LOC_96/A INVX1_LOC_38/A 0.33fF
C76050 INVX1_LOC_58/A NOR2X1_LOC_637/Y 0.14fF
C76051 NOR2X1_LOC_74/A INVX1_LOC_92/A 3.34fF
C76052 NOR2X1_LOC_719/A INVX1_LOC_42/A 0.01fF
C76053 NAND2X1_LOC_815/a_36_24# INVX1_LOC_63/A 0.00fF
C76054 NOR2X1_LOC_68/A INVX1_LOC_138/A 0.01fF
C76055 NAND2X1_LOC_629/Y INVX1_LOC_78/A 0.05fF
C76056 INVX1_LOC_33/A NOR2X1_LOC_72/Y 0.01fF
C76057 INVX1_LOC_48/Y NOR2X1_LOC_530/Y 0.01fF
C76058 INVX1_LOC_58/A INVX1_LOC_172/A 0.09fF
C76059 NOR2X1_LOC_9/Y INVX1_LOC_92/A 0.64fF
C76060 NOR2X1_LOC_381/a_36_216# INVX1_LOC_3/A 0.02fF
C76061 NOR2X1_LOC_561/Y INVX1_LOC_42/A 0.02fF
C76062 D_INPUT_0 INVX1_LOC_12/A 0.03fF
C76063 NOR2X1_LOC_32/B NOR2X1_LOC_617/Y 0.04fF
C76064 NOR2X1_LOC_373/Y NOR2X1_LOC_89/A 0.07fF
C76065 NOR2X1_LOC_423/a_36_216# NOR2X1_LOC_759/Y 0.00fF
C76066 INVX1_LOC_7/A INVX1_LOC_42/A 0.09fF
C76067 NOR2X1_LOC_817/Y INVX1_LOC_11/A 0.01fF
C76068 NOR2X1_LOC_667/Y NAND2X1_LOC_579/A 0.07fF
C76069 NOR2X1_LOC_456/Y NOR2X1_LOC_550/B 0.10fF
C76070 NOR2X1_LOC_647/a_36_216# INVX1_LOC_269/A 0.05fF
C76071 NAND2X1_LOC_557/Y INVX1_LOC_34/A 0.06fF
C76072 NAND2X1_LOC_102/a_36_24# INVX1_LOC_3/A 0.00fF
C76073 NOR2X1_LOC_817/Y NAND2X1_LOC_381/Y 0.03fF
C76074 INVX1_LOC_21/A D_INPUT_7 0.00fF
C76075 INVX1_LOC_299/A NOR2X1_LOC_590/A 0.09fF
C76076 INVX1_LOC_63/Y INVX1_LOC_23/A 0.07fF
C76077 NOR2X1_LOC_71/Y NAND2X1_LOC_254/Y 0.00fF
C76078 NAND2X1_LOC_35/Y NOR2X1_LOC_403/a_36_216# 0.01fF
C76079 NOR2X1_LOC_160/B NOR2X1_LOC_103/Y 0.09fF
C76080 NOR2X1_LOC_690/A NAND2X1_LOC_860/A 0.01fF
C76081 INVX1_LOC_16/A NOR2X1_LOC_334/Y 0.07fF
C76082 INVX1_LOC_131/A INVX1_LOC_19/A 0.13fF
C76083 INVX1_LOC_206/A NOR2X1_LOC_383/B 0.00fF
C76084 NOR2X1_LOC_220/a_36_216# NOR2X1_LOC_798/A 0.00fF
C76085 INVX1_LOC_36/A NOR2X1_LOC_468/Y 0.30fF
C76086 INVX1_LOC_64/A NAND2X1_LOC_361/Y 0.07fF
C76087 INVX1_LOC_161/A INVX1_LOC_161/Y 0.09fF
C76088 NOR2X1_LOC_510/Y NOR2X1_LOC_13/Y 0.10fF
C76089 INVX1_LOC_256/A NOR2X1_LOC_441/Y 0.01fF
C76090 INVX1_LOC_30/Y NAND2X1_LOC_223/A 0.02fF
C76091 INVX1_LOC_259/Y INVX1_LOC_257/Y 0.01fF
C76092 INVX1_LOC_237/Y INVX1_LOC_5/A 0.01fF
C76093 NOR2X1_LOC_585/Y NAND2X1_LOC_637/Y 0.02fF
C76094 NOR2X1_LOC_210/a_36_216# NOR2X1_LOC_68/A -0.02fF
C76095 INPUT_0 INVX1_LOC_19/A 10.89fF
C76096 NOR2X1_LOC_409/a_36_216# NOR2X1_LOC_409/B 0.00fF
C76097 NOR2X1_LOC_626/a_36_216# INVX1_LOC_113/Y 0.00fF
C76098 NAND2X1_LOC_656/Y INVX1_LOC_4/Y 0.07fF
C76099 NOR2X1_LOC_561/Y INVX1_LOC_78/A 0.14fF
C76100 INVX1_LOC_64/A INVX1_LOC_219/Y 0.01fF
C76101 INVX1_LOC_36/A NAND2X1_LOC_396/a_36_24# 0.00fF
C76102 INVX1_LOC_144/A INVX1_LOC_272/A 0.13fF
C76103 INVX1_LOC_12/Y NOR2X1_LOC_331/B 0.01fF
C76104 INVX1_LOC_33/A INVX1_LOC_50/Y 0.03fF
C76105 INVX1_LOC_177/A NOR2X1_LOC_717/A 0.04fF
C76106 INVX1_LOC_49/A NAND2X1_LOC_474/Y 0.01fF
C76107 NOR2X1_LOC_631/B NOR2X1_LOC_197/B 0.01fF
C76108 NAND2X1_LOC_468/B NOR2X1_LOC_58/Y 0.26fF
C76109 NOR2X1_LOC_717/B NOR2X1_LOC_465/Y 0.12fF
C76110 NOR2X1_LOC_299/Y NOR2X1_LOC_409/B 0.07fF
C76111 NOR2X1_LOC_510/Y NAND2X1_LOC_175/B 0.01fF
C76112 INVX1_LOC_45/A NOR2X1_LOC_160/B 5.80fF
C76113 INVX1_LOC_35/A NOR2X1_LOC_111/a_36_216# 0.02fF
C76114 VDD NOR2X1_LOC_640/Y 0.57fF
C76115 INVX1_LOC_38/A NOR2X1_LOC_684/Y 0.07fF
C76116 INVX1_LOC_208/Y INVX1_LOC_270/Y 0.08fF
C76117 INVX1_LOC_161/Y INVX1_LOC_79/Y 0.02fF
C76118 INVX1_LOC_137/A NOR2X1_LOC_383/B 0.13fF
C76119 INVX1_LOC_16/A NAND2X1_LOC_464/B 0.01fF
C76120 INVX1_LOC_36/A NOR2X1_LOC_389/A 0.01fF
C76121 INVX1_LOC_215/Y INVX1_LOC_18/A 0.00fF
C76122 NOR2X1_LOC_468/Y NOR2X1_LOC_237/Y 0.00fF
C76123 D_INPUT_1 INVX1_LOC_56/Y 0.12fF
C76124 NAND2X1_LOC_363/B NOR2X1_LOC_346/B 0.07fF
C76125 INVX1_LOC_50/A NOR2X1_LOC_589/A 0.03fF
C76126 NOR2X1_LOC_65/B NOR2X1_LOC_561/Y 0.07fF
C76127 INVX1_LOC_47/A INVX1_LOC_87/A 0.25fF
C76128 INVX1_LOC_266/A INVX1_LOC_33/A 0.01fF
C76129 INVX1_LOC_73/A INVX1_LOC_47/Y 0.19fF
C76130 INVX1_LOC_286/A NOR2X1_LOC_89/A 0.08fF
C76131 INVX1_LOC_37/A NOR2X1_LOC_197/B 0.08fF
C76132 NOR2X1_LOC_167/Y INVX1_LOC_42/A 0.03fF
C76133 INVX1_LOC_28/A NOR2X1_LOC_334/Y 0.07fF
C76134 NOR2X1_LOC_15/Y NOR2X1_LOC_772/Y 0.34fF
C76135 INVX1_LOC_280/A NOR2X1_LOC_629/Y 0.00fF
C76136 VDD NAND2X1_LOC_85/Y 0.41fF
C76137 INVX1_LOC_36/A NAND2X1_LOC_708/a_36_24# 0.00fF
C76138 NOR2X1_LOC_763/Y INVX1_LOC_296/A 0.44fF
C76139 INVX1_LOC_34/A NOR2X1_LOC_122/A 0.00fF
C76140 INVX1_LOC_30/A NOR2X1_LOC_274/B 0.01fF
C76141 NAND2X1_LOC_714/B NAND2X1_LOC_802/a_36_24# 0.00fF
C76142 NAND2X1_LOC_363/B INVX1_LOC_22/A 0.00fF
C76143 NOR2X1_LOC_491/Y NOR2X1_LOC_492/Y 0.01fF
C76144 VDD NOR2X1_LOC_697/Y 1.04fF
C76145 NAND2X1_LOC_53/Y INVX1_LOC_49/A 0.14fF
C76146 NOR2X1_LOC_78/B INVX1_LOC_306/Y 0.17fF
C76147 NOR2X1_LOC_160/B INVX1_LOC_71/A 0.17fF
C76148 NOR2X1_LOC_15/Y NOR2X1_LOC_392/B 0.01fF
C76149 NAND2X1_LOC_87/a_36_24# NAND2X1_LOC_859/B 0.01fF
C76150 NAND2X1_LOC_465/A NAND2X1_LOC_773/B 0.02fF
C76151 INVX1_LOC_6/A INVX1_LOC_251/A 0.05fF
C76152 INVX1_LOC_48/Y NOR2X1_LOC_709/A 0.18fF
C76153 NOR2X1_LOC_151/Y NOR2X1_LOC_465/Y 0.00fF
C76154 NOR2X1_LOC_140/A NOR2X1_LOC_84/Y 0.02fF
C76155 NOR2X1_LOC_226/A NAND2X1_LOC_474/Y 0.04fF
C76156 NAND2X1_LOC_468/B INVX1_LOC_29/A 0.03fF
C76157 INVX1_LOC_95/A NOR2X1_LOC_89/A 0.03fF
C76158 INVX1_LOC_34/A INVX1_LOC_161/Y 0.07fF
C76159 INVX1_LOC_256/A NOR2X1_LOC_142/Y 0.14fF
C76160 INVX1_LOC_36/A NOR2X1_LOC_596/A 0.31fF
C76161 INVX1_LOC_17/A INVX1_LOC_104/A 0.13fF
C76162 NOR2X1_LOC_641/B INVX1_LOC_314/Y 0.48fF
C76163 NOR2X1_LOC_533/Y NOR2X1_LOC_591/Y 0.02fF
C76164 INVX1_LOC_54/Y INVX1_LOC_14/A 0.03fF
C76165 NAND2X1_LOC_732/a_36_24# INVX1_LOC_173/Y 0.01fF
C76166 NAND2X1_LOC_842/B INVX1_LOC_57/A 0.14fF
C76167 NAND2X1_LOC_96/A NOR2X1_LOC_814/A 0.07fF
C76168 NOR2X1_LOC_457/A NOR2X1_LOC_348/B 0.35fF
C76169 INVX1_LOC_230/Y NAND2X1_LOC_139/A 0.03fF
C76170 INVX1_LOC_28/A NAND2X1_LOC_464/B 0.03fF
C76171 NOR2X1_LOC_167/Y INVX1_LOC_78/A 0.03fF
C76172 NOR2X1_LOC_360/Y NOR2X1_LOC_359/Y 0.03fF
C76173 INVX1_LOC_30/A NOR2X1_LOC_577/Y 0.17fF
C76174 INVX1_LOC_2/A INVX1_LOC_272/Y 0.03fF
C76175 NAND2X1_LOC_392/Y INVX1_LOC_306/Y 0.01fF
C76176 INVX1_LOC_146/A INVX1_LOC_57/A 0.01fF
C76177 NOR2X1_LOC_361/B INVX1_LOC_256/Y 0.10fF
C76178 INVX1_LOC_227/Y NOR2X1_LOC_303/Y 0.05fF
C76179 INVX1_LOC_24/A NAND2X1_LOC_198/B 0.06fF
C76180 NOR2X1_LOC_590/A NOR2X1_LOC_350/a_36_216# 0.02fF
C76181 INVX1_LOC_2/A NAND2X1_LOC_53/Y 0.07fF
C76182 NOR2X1_LOC_34/A NOR2X1_LOC_33/A 0.21fF
C76183 NOR2X1_LOC_669/A NOR2X1_LOC_305/Y 0.01fF
C76184 INVX1_LOC_12/A NOR2X1_LOC_266/B 0.02fF
C76185 INPUT_0 INVX1_LOC_26/Y 0.06fF
C76186 NOR2X1_LOC_356/A INVX1_LOC_53/A 0.07fF
C76187 NOR2X1_LOC_389/A NOR2X1_LOC_309/Y 0.00fF
C76188 INVX1_LOC_272/Y NOR2X1_LOC_226/A 0.07fF
C76189 NOR2X1_LOC_273/Y NOR2X1_LOC_759/Y 0.02fF
C76190 INVX1_LOC_76/A INVX1_LOC_42/A 0.79fF
C76191 INVX1_LOC_34/A NOR2X1_LOC_599/A 0.03fF
C76192 INVX1_LOC_134/A INVX1_LOC_196/A 0.05fF
C76193 NAND2X1_LOC_231/Y INVX1_LOC_161/Y 0.10fF
C76194 INVX1_LOC_72/A INVX1_LOC_155/A 0.03fF
C76195 INVX1_LOC_256/A NOR2X1_LOC_655/B 0.10fF
C76196 NAND2X1_LOC_773/Y INVX1_LOC_1/Y 0.03fF
C76197 NOR2X1_LOC_208/Y NOR2X1_LOC_596/A 0.07fF
C76198 INVX1_LOC_5/A NAND2X1_LOC_45/Y 0.27fF
C76199 NOR2X1_LOC_34/B NOR2X1_LOC_332/A 0.02fF
C76200 INVX1_LOC_246/Y NAND2X1_LOC_802/A 0.01fF
C76201 NOR2X1_LOC_295/Y INVX1_LOC_36/A 0.03fF
C76202 NAND2X1_LOC_181/Y NAND2X1_LOC_793/Y 0.01fF
C76203 INVX1_LOC_50/A INVX1_LOC_222/A 0.05fF
C76204 NAND2X1_LOC_704/a_36_24# NAND2X1_LOC_319/A 0.01fF
C76205 NAND2X1_LOC_725/A NOR2X1_LOC_385/a_36_216# 0.15fF
C76206 NOR2X1_LOC_168/Y NOR2X1_LOC_344/A 0.02fF
C76207 INVX1_LOC_310/A INVX1_LOC_22/Y 0.12fF
C76208 NOR2X1_LOC_418/Y NAND2X1_LOC_227/Y 0.16fF
C76209 NAND2X1_LOC_571/B INVX1_LOC_282/A 0.06fF
C76210 NOR2X1_LOC_454/Y NOR2X1_LOC_639/a_36_216# 0.01fF
C76211 NAND2X1_LOC_778/Y INVX1_LOC_90/A 0.01fF
C76212 NOR2X1_LOC_457/A INVX1_LOC_22/A 0.15fF
C76213 NOR2X1_LOC_74/A INVX1_LOC_53/A 0.14fF
C76214 INVX1_LOC_95/Y INVX1_LOC_87/A 0.01fF
C76215 NOR2X1_LOC_496/Y NAND2X1_LOC_866/B 0.07fF
C76216 INPUT_1 NAND2X1_LOC_474/Y 0.01fF
C76217 INVX1_LOC_226/Y NOR2X1_LOC_134/Y 0.03fF
C76218 NOR2X1_LOC_334/Y NOR2X1_LOC_35/Y 0.10fF
C76219 INVX1_LOC_26/A NAND2X1_LOC_642/Y 0.40fF
C76220 INVX1_LOC_34/A NOR2X1_LOC_437/Y 0.09fF
C76221 NAND2X1_LOC_471/Y NAND2X1_LOC_464/A 0.20fF
C76222 NOR2X1_LOC_9/Y INVX1_LOC_53/A 0.01fF
C76223 INVX1_LOC_269/A INVX1_LOC_135/A 0.29fF
C76224 INVX1_LOC_72/A NAND2X1_LOC_661/B 0.02fF
C76225 NOR2X1_LOC_232/Y INVX1_LOC_135/A 0.01fF
C76226 NAND2X1_LOC_574/A NOR2X1_LOC_673/A 0.02fF
C76227 INVX1_LOC_78/A INVX1_LOC_76/A 0.31fF
C76228 NOR2X1_LOC_794/B NOR2X1_LOC_553/B 0.03fF
C76229 INVX1_LOC_36/A NOR2X1_LOC_220/A 0.06fF
C76230 NOR2X1_LOC_89/A INVX1_LOC_54/A 0.12fF
C76231 NOR2X1_LOC_561/Y NOR2X1_LOC_503/Y 0.07fF
C76232 INVX1_LOC_279/Y NOR2X1_LOC_687/Y 0.09fF
C76233 NOR2X1_LOC_401/A NOR2X1_LOC_123/B 0.01fF
C76234 INVX1_LOC_228/Y D_INPUT_0 0.05fF
C76235 NOR2X1_LOC_15/Y INVX1_LOC_90/A 1.45fF
C76236 INVX1_LOC_45/A INVX1_LOC_208/A 0.03fF
C76237 NAND2X1_LOC_727/Y NAND2X1_LOC_733/Y 0.04fF
C76238 INVX1_LOC_200/A D_INPUT_0 0.03fF
C76239 NAND2X1_LOC_433/a_36_24# NOR2X1_LOC_435/A 0.02fF
C76240 INVX1_LOC_14/Y NAND2X1_LOC_454/Y 0.10fF
C76241 NOR2X1_LOC_848/Y NOR2X1_LOC_814/Y 0.01fF
C76242 NOR2X1_LOC_382/Y INVX1_LOC_25/Y 0.02fF
C76243 INVX1_LOC_58/A NOR2X1_LOC_43/a_36_216# 0.00fF
C76244 INVX1_LOC_75/A NOR2X1_LOC_460/Y 0.01fF
C76245 INVX1_LOC_45/A NOR2X1_LOC_516/B 0.10fF
C76246 NOR2X1_LOC_15/Y NOR2X1_LOC_389/B 0.24fF
C76247 NOR2X1_LOC_155/A INVX1_LOC_272/A 0.07fF
C76248 INVX1_LOC_207/A NAND2X1_LOC_736/B 0.02fF
C76249 INVX1_LOC_30/A INVX1_LOC_22/A 0.63fF
C76250 INVX1_LOC_272/Y NAND2X1_LOC_648/A 0.00fF
C76251 INVX1_LOC_49/Y NOR2X1_LOC_841/A 0.01fF
C76252 NAND2X1_LOC_475/Y NAND2X1_LOC_476/Y 0.05fF
C76253 NAND2X1_LOC_84/Y INVX1_LOC_54/Y 0.00fF
C76254 NAND2X1_LOC_254/Y NAND2X1_LOC_243/Y 0.33fF
C76255 NOR2X1_LOC_229/Y INVX1_LOC_72/A 0.03fF
C76256 NOR2X1_LOC_545/B INVX1_LOC_57/A -0.01fF
C76257 NOR2X1_LOC_443/a_36_216# INVX1_LOC_148/Y 0.00fF
C76258 NOR2X1_LOC_111/A NAND2X1_LOC_175/Y 1.53fF
C76259 NOR2X1_LOC_819/a_36_216# NOR2X1_LOC_516/B 0.01fF
C76260 NOR2X1_LOC_65/B INVX1_LOC_76/A -0.00fF
C76261 NAND2X1_LOC_629/Y INVX1_LOC_113/Y 0.02fF
C76262 NOR2X1_LOC_791/Y INVX1_LOC_100/A 0.57fF
C76263 NOR2X1_LOC_160/B NOR2X1_LOC_123/B 0.07fF
C76264 INVX1_LOC_269/A NAND2X1_LOC_184/a_36_24# 0.00fF
C76265 NAND2X1_LOC_141/Y INVX1_LOC_29/A 0.35fF
C76266 INVX1_LOC_64/A INVX1_LOC_159/Y 0.10fF
C76267 NOR2X1_LOC_609/Y INVX1_LOC_9/A 0.01fF
C76268 INVX1_LOC_297/Y INVX1_LOC_300/Y 0.01fF
C76269 NOR2X1_LOC_590/A INVX1_LOC_66/A 0.00fF
C76270 INVX1_LOC_50/A INVX1_LOC_20/A 0.15fF
C76271 INVX1_LOC_163/A NAND2X1_LOC_463/B 0.00fF
C76272 INVX1_LOC_150/Y NOR2X1_LOC_768/a_36_216# 0.00fF
C76273 NOR2X1_LOC_220/A NOR2X1_LOC_208/Y 0.03fF
C76274 NOR2X1_LOC_295/Y NOR2X1_LOC_309/Y 0.02fF
C76275 NAND2X1_LOC_493/Y INVX1_LOC_282/A 0.05fF
C76276 NOR2X1_LOC_606/Y NOR2X1_LOC_99/B 0.04fF
C76277 INVX1_LOC_38/A INVX1_LOC_273/A 0.39fF
C76278 NOR2X1_LOC_401/Y NOR2X1_LOC_716/B 0.04fF
C76279 INVX1_LOC_208/A INVX1_LOC_71/A 0.08fF
C76280 NOR2X1_LOC_619/A INVX1_LOC_24/A 0.41fF
C76281 INVX1_LOC_77/Y NOR2X1_LOC_639/Y 0.04fF
C76282 INVX1_LOC_7/A NOR2X1_LOC_554/B 0.08fF
C76283 NOR2X1_LOC_789/B INVX1_LOC_123/A 0.04fF
C76284 INVX1_LOC_310/Y INVX1_LOC_143/A 0.09fF
C76285 INVX1_LOC_225/A INVX1_LOC_149/A 0.02fF
C76286 NAND2X1_LOC_562/B NAND2X1_LOC_556/a_36_24# 0.02fF
C76287 NAND2X1_LOC_569/A NAND2X1_LOC_338/B 0.02fF
C76288 NOR2X1_LOC_264/Y NOR2X1_LOC_537/Y 1.20fF
C76289 INVX1_LOC_49/A NOR2X1_LOC_500/Y 0.09fF
C76290 NAND2X1_LOC_483/Y NOR2X1_LOC_526/Y 0.08fF
C76291 INVX1_LOC_226/Y INVX1_LOC_49/A 0.11fF
C76292 INVX1_LOC_269/A NOR2X1_LOC_391/B 0.25fF
C76293 D_INPUT_0 INVX1_LOC_217/A 0.00fF
C76294 NAND2X1_LOC_267/B NOR2X1_LOC_717/A 0.21fF
C76295 NAND2X1_LOC_544/a_36_24# INVX1_LOC_20/A 0.01fF
C76296 NOR2X1_LOC_662/A INVX1_LOC_284/A 0.03fF
C76297 INVX1_LOC_209/Y INVX1_LOC_16/A 0.03fF
C76298 VDD NOR2X1_LOC_247/Y 0.03fF
C76299 INVX1_LOC_105/A NOR2X1_LOC_589/A 0.15fF
C76300 NOR2X1_LOC_246/A NAND2X1_LOC_364/A 0.11fF
C76301 INVX1_LOC_54/Y NOR2X1_LOC_612/B 0.03fF
C76302 INVX1_LOC_161/Y INPUT_0 0.07fF
C76303 NOR2X1_LOC_557/Y INVX1_LOC_53/Y 0.19fF
C76304 NAND2X1_LOC_364/A NOR2X1_LOC_174/B 0.03fF
C76305 INVX1_LOC_36/Y INVX1_LOC_68/A 0.01fF
C76306 NOR2X1_LOC_561/Y NOR2X1_LOC_152/Y 0.10fF
C76307 NOR2X1_LOC_585/a_36_216# NAND2X1_LOC_654/B 0.00fF
C76308 NOR2X1_LOC_413/Y INVX1_LOC_172/Y 0.02fF
C76309 NAND2X1_LOC_326/A INVX1_LOC_91/A 0.09fF
C76310 NOR2X1_LOC_6/B INVX1_LOC_40/A 0.91fF
C76311 INVX1_LOC_30/Y INVX1_LOC_33/A 0.02fF
C76312 NAND2X1_LOC_166/a_36_24# NOR2X1_LOC_356/A 0.01fF
C76313 INVX1_LOC_11/A INVX1_LOC_286/A 0.07fF
C76314 INVX1_LOC_122/Y NAND2X1_LOC_508/A 0.05fF
C76315 INVX1_LOC_226/Y INVX1_LOC_60/A 0.01fF
C76316 NAND2X1_LOC_72/B NOR2X1_LOC_197/B 0.01fF
C76317 INVX1_LOC_234/A NAND2X1_LOC_632/B 0.06fF
C76318 INVX1_LOC_49/A INVX1_LOC_10/A 0.49fF
C76319 NAND2X1_LOC_364/Y NOR2X1_LOC_785/Y 0.01fF
C76320 NOR2X1_LOC_488/Y NOR2X1_LOC_315/Y 0.28fF
C76321 NOR2X1_LOC_718/B INVX1_LOC_16/A 0.03fF
C76322 INVX1_LOC_314/Y NOR2X1_LOC_71/Y 0.02fF
C76323 INVX1_LOC_45/A NOR2X1_LOC_706/A 0.00fF
C76324 NOR2X1_LOC_315/Y NOR2X1_LOC_82/Y 0.00fF
C76325 INVX1_LOC_46/A INVX1_LOC_306/Y 0.06fF
C76326 NAND2X1_LOC_773/Y INVX1_LOC_93/Y 0.10fF
C76327 INVX1_LOC_135/A NOR2X1_LOC_360/a_36_216# 0.00fF
C76328 NOR2X1_LOC_89/A NAND2X1_LOC_807/B 0.03fF
C76329 NAND2X1_LOC_827/a_36_24# NOR2X1_LOC_536/A -0.00fF
C76330 INVX1_LOC_269/A NOR2X1_LOC_552/A 0.15fF
C76331 NOR2X1_LOC_363/a_36_216# INVX1_LOC_313/Y 0.00fF
C76332 NAND2X1_LOC_198/a_36_24# NOR2X1_LOC_368/A 0.00fF
C76333 INVX1_LOC_2/A NOR2X1_LOC_500/Y 0.07fF
C76334 INVX1_LOC_90/A NOR2X1_LOC_860/B 0.08fF
C76335 NAND2X1_LOC_7/Y INVX1_LOC_89/A 0.27fF
C76336 NOR2X1_LOC_215/A INVX1_LOC_76/A 0.03fF
C76337 NOR2X1_LOC_38/B INVX1_LOC_63/A 0.08fF
C76338 INVX1_LOC_2/A INVX1_LOC_226/Y 0.10fF
C76339 INVX1_LOC_170/A NOR2X1_LOC_368/A 0.08fF
C76340 INVX1_LOC_215/A NOR2X1_LOC_52/B 0.07fF
C76341 INVX1_LOC_21/A INVX1_LOC_2/Y 0.03fF
C76342 NOR2X1_LOC_599/A INPUT_0 0.00fF
C76343 NAND2X1_LOC_722/A INVX1_LOC_22/A 0.05fF
C76344 D_INPUT_7 NAND2X1_LOC_51/B 0.10fF
C76345 NAND2X1_LOC_588/B D_INPUT_4 0.01fF
C76346 NAND2X1_LOC_530/a_36_24# INVX1_LOC_75/A 0.00fF
C76347 NOR2X1_LOC_788/B INVX1_LOC_77/A 0.02fF
C76348 INVX1_LOC_298/A INVX1_LOC_117/A 0.02fF
C76349 NOR2X1_LOC_89/A NOR2X1_LOC_48/B 0.21fF
C76350 INVX1_LOC_45/Y NAND2X1_LOC_123/Y 0.02fF
C76351 INVX1_LOC_54/A NAND2X1_LOC_804/A 0.01fF
C76352 INVX1_LOC_30/A INVX1_LOC_100/A 0.02fF
C76353 NOR2X1_LOC_658/Y INVX1_LOC_285/Y 0.03fF
C76354 NAND2X1_LOC_668/a_36_24# NOR2X1_LOC_48/B 0.00fF
C76355 NOR2X1_LOC_454/Y NAND2X1_LOC_39/Y 0.03fF
C76356 INVX1_LOC_11/A INVX1_LOC_95/A 0.04fF
C76357 NOR2X1_LOC_107/Y NAND2X1_LOC_642/Y 0.01fF
C76358 INVX1_LOC_230/Y NOR2X1_LOC_78/A 0.84fF
C76359 NAND2X1_LOC_154/Y INVX1_LOC_6/A 0.02fF
C76360 NAND2X1_LOC_360/B INVX1_LOC_137/Y 0.06fF
C76361 NOR2X1_LOC_717/B NOR2X1_LOC_180/Y 0.00fF
C76362 NOR2X1_LOC_82/A INVX1_LOC_95/Y 0.09fF
C76363 NAND2X1_LOC_670/a_36_24# INVX1_LOC_48/A 0.01fF
C76364 NAND2X1_LOC_866/A NOR2X1_LOC_380/Y 0.16fF
C76365 INVX1_LOC_2/A INVX1_LOC_10/A 0.14fF
C76366 NOR2X1_LOC_817/Y INVX1_LOC_74/A 0.04fF
C76367 D_INPUT_1 NOR2X1_LOC_831/B 0.03fF
C76368 NAND2X1_LOC_348/A NOR2X1_LOC_860/B 0.12fF
C76369 NOR2X1_LOC_470/B INVX1_LOC_37/A 0.00fF
C76370 INVX1_LOC_229/Y INVX1_LOC_209/A 0.03fF
C76371 NAND2X1_LOC_308/Y NAND2X1_LOC_308/B 0.00fF
C76372 INVX1_LOC_30/Y INVX1_LOC_40/A 0.02fF
C76373 INVX1_LOC_256/Y NAND2X1_LOC_573/A 0.03fF
C76374 NOR2X1_LOC_226/A INVX1_LOC_10/A 0.16fF
C76375 NOR2X1_LOC_334/Y INVX1_LOC_109/A 0.01fF
C76376 INVX1_LOC_57/Y NOR2X1_LOC_528/Y 0.10fF
C76377 NOR2X1_LOC_751/A INVX1_LOC_314/Y 0.01fF
C76378 D_INPUT_1 NOR2X1_LOC_179/a_36_216# 0.00fF
C76379 NOR2X1_LOC_93/Y INVX1_LOC_280/A 0.03fF
C76380 NOR2X1_LOC_75/Y NOR2X1_LOC_603/Y 0.01fF
C76381 NOR2X1_LOC_437/Y INPUT_0 0.12fF
C76382 INVX1_LOC_54/Y NOR2X1_LOC_137/A 0.02fF
C76383 NOR2X1_LOC_267/A INVX1_LOC_100/Y 0.07fF
C76384 NOR2X1_LOC_93/Y NOR2X1_LOC_94/Y 0.14fF
C76385 INVX1_LOC_57/A INVX1_LOC_119/Y 0.01fF
C76386 NOR2X1_LOC_616/Y INVX1_LOC_135/A 0.04fF
C76387 INVX1_LOC_312/Y NOR2X1_LOC_595/Y 0.09fF
C76388 NOR2X1_LOC_717/B NOR2X1_LOC_458/B 0.02fF
C76389 INVX1_LOC_237/Y NAND2X1_LOC_463/B 0.00fF
C76390 NAND2X1_LOC_53/Y NAND2X1_LOC_605/a_36_24# 0.01fF
C76391 NAND2X1_LOC_579/A NOR2X1_LOC_536/A 0.15fF
C76392 NOR2X1_LOC_15/Y NAND2X1_LOC_849/B 0.08fF
C76393 NOR2X1_LOC_232/Y NOR2X1_LOC_813/Y 0.04fF
C76394 NAND2X1_LOC_563/A INVX1_LOC_135/A 0.17fF
C76395 INVX1_LOC_232/Y INVX1_LOC_89/A 0.15fF
C76396 NOR2X1_LOC_218/Y INVX1_LOC_10/A 0.03fF
C76397 NAND2X1_LOC_866/B NAND2X1_LOC_839/A 0.02fF
C76398 NOR2X1_LOC_15/Y INVX1_LOC_38/A 0.29fF
C76399 NOR2X1_LOC_625/Y INVX1_LOC_309/A 0.01fF
C76400 NAND2X1_LOC_149/Y NAND2X1_LOC_637/Y 0.15fF
C76401 NOR2X1_LOC_831/Y NOR2X1_LOC_831/a_36_216# 0.02fF
C76402 NOR2X1_LOC_369/Y INVX1_LOC_37/A 0.04fF
C76403 INVX1_LOC_269/A INVX1_LOC_280/A 0.10fF
C76404 NOR2X1_LOC_763/Y INVX1_LOC_268/Y 0.00fF
C76405 NAND2X1_LOC_776/a_36_24# NOR2X1_LOC_164/Y 0.00fF
C76406 NOR2X1_LOC_89/A NOR2X1_LOC_438/Y 0.00fF
C76407 NOR2X1_LOC_778/B NOR2X1_LOC_644/A 2.79fF
C76408 NAND2X1_LOC_549/Y INVX1_LOC_84/A 0.01fF
C76409 NOR2X1_LOC_151/Y NOR2X1_LOC_180/Y 0.03fF
C76410 NOR2X1_LOC_78/B NOR2X1_LOC_356/A 0.08fF
C76411 INVX1_LOC_200/A NAND2X1_LOC_848/A 0.01fF
C76412 INVX1_LOC_83/A NAND2X1_LOC_149/B 0.04fF
C76413 INVX1_LOC_90/A NAND2X1_LOC_840/B 0.02fF
C76414 INVX1_LOC_32/A INVX1_LOC_90/Y 0.03fF
C76415 INVX1_LOC_27/A INVX1_LOC_179/A 0.02fF
C76416 NOR2X1_LOC_593/Y INVX1_LOC_286/A 0.01fF
C76417 NOR2X1_LOC_690/A NOR2X1_LOC_86/a_36_216# 0.00fF
C76418 INVX1_LOC_63/Y INVX1_LOC_6/A 0.17fF
C76419 NOR2X1_LOC_68/A NAND2X1_LOC_212/Y 0.05fF
C76420 NOR2X1_LOC_125/Y INVX1_LOC_272/A 0.02fF
C76421 INVX1_LOC_286/Y INVX1_LOC_37/A 0.07fF
C76422 INVX1_LOC_69/Y NOR2X1_LOC_142/Y 0.01fF
C76423 NAND2X1_LOC_555/Y NAND2X1_LOC_8/a_36_24# 0.01fF
C76424 NOR2X1_LOC_426/Y VDD 0.03fF
C76425 INVX1_LOC_226/Y INPUT_1 0.74fF
C76426 NOR2X1_LOC_778/B NOR2X1_LOC_828/B 0.00fF
C76427 NOR2X1_LOC_769/A INVX1_LOC_76/A 0.15fF
C76428 NOR2X1_LOC_242/A NOR2X1_LOC_865/Y 0.07fF
C76429 NOR2X1_LOC_210/A INVX1_LOC_89/A 0.03fF
C76430 INVX1_LOC_194/A NAND2X1_LOC_622/B 0.00fF
C76431 INVX1_LOC_191/Y INVX1_LOC_302/Y 0.08fF
C76432 NOR2X1_LOC_755/a_36_216# NOR2X1_LOC_757/Y -0.00fF
C76433 NOR2X1_LOC_590/A NAND2X1_LOC_96/A 0.08fF
C76434 NOR2X1_LOC_644/A NOR2X1_LOC_439/a_36_216# 0.00fF
C76435 NOR2X1_LOC_510/Y NOR2X1_LOC_697/Y 0.03fF
C76436 INVX1_LOC_36/A NOR2X1_LOC_447/B 0.00fF
C76437 INVX1_LOC_57/A INVX1_LOC_284/A 0.24fF
C76438 NOR2X1_LOC_647/A INVX1_LOC_3/Y 0.03fF
C76439 NOR2X1_LOC_160/B NOR2X1_LOC_331/B 0.07fF
C76440 INVX1_LOC_11/A INVX1_LOC_54/A 0.12fF
C76441 INVX1_LOC_24/A NAND2X1_LOC_465/A 0.00fF
C76442 NOR2X1_LOC_662/A NOR2X1_LOC_663/A 0.14fF
C76443 NOR2X1_LOC_561/Y NOR2X1_LOC_150/a_36_216# 0.03fF
C76444 NOR2X1_LOC_458/B NOR2X1_LOC_151/Y 0.00fF
C76445 INVX1_LOC_277/A NOR2X1_LOC_698/Y 0.00fF
C76446 INVX1_LOC_14/A NAND2X1_LOC_656/B 0.01fF
C76447 NAND2X1_LOC_363/B NOR2X1_LOC_777/B 0.06fF
C76448 INVX1_LOC_286/A NOR2X1_LOC_52/B 0.07fF
C76449 NOR2X1_LOC_68/A D_INPUT_3 0.00fF
C76450 NOR2X1_LOC_433/A INVX1_LOC_95/A 0.12fF
C76451 NOR2X1_LOC_420/Y INVX1_LOC_63/A 0.03fF
C76452 NOR2X1_LOC_78/B NOR2X1_LOC_74/A 0.15fF
C76453 NOR2X1_LOC_68/A INVX1_LOC_14/Y 0.09fF
C76454 INVX1_LOC_10/A NAND2X1_LOC_648/A 0.03fF
C76455 INVX1_LOC_159/A INVX1_LOC_37/A 0.01fF
C76456 INVX1_LOC_10/A INPUT_1 0.03fF
C76457 INVX1_LOC_24/A NAND2X1_LOC_242/a_36_24# 0.00fF
C76458 NOR2X1_LOC_667/A NAND2X1_LOC_325/a_36_24# 0.00fF
C76459 NAND2X1_LOC_214/B NAND2X1_LOC_215/a_36_24# 0.00fF
C76460 NAND2X1_LOC_541/a_36_24# INVX1_LOC_284/A 0.00fF
C76461 INVX1_LOC_88/A NOR2X1_LOC_58/Y 0.01fF
C76462 NOR2X1_LOC_473/B NOR2X1_LOC_366/Y 0.01fF
C76463 NOR2X1_LOC_443/Y INVX1_LOC_15/A 0.02fF
C76464 NOR2X1_LOC_772/B INVX1_LOC_29/A 0.05fF
C76465 NOR2X1_LOC_655/B INVX1_LOC_69/Y 0.10fF
C76466 INVX1_LOC_33/A INVX1_LOC_188/Y 0.09fF
C76467 NAND2X1_LOC_715/B INVX1_LOC_272/A 0.01fF
C76468 NOR2X1_LOC_78/B NOR2X1_LOC_9/Y 0.50fF
C76469 NOR2X1_LOC_152/Y INVX1_LOC_76/A 0.57fF
C76470 NAND2X1_LOC_347/B INVX1_LOC_84/A 0.03fF
C76471 NOR2X1_LOC_411/A INVX1_LOC_42/A 0.19fF
C76472 INVX1_LOC_245/Y INVX1_LOC_92/A 0.03fF
C76473 INVX1_LOC_50/A INVX1_LOC_4/A 0.00fF
C76474 NAND2X1_LOC_364/A INVX1_LOC_66/Y 0.05fF
C76475 INVX1_LOC_150/Y NOR2X1_LOC_155/A 0.90fF
C76476 NOR2X1_LOC_301/A NOR2X1_LOC_281/a_36_216# 0.00fF
C76477 INVX1_LOC_13/Y INVX1_LOC_29/A 0.07fF
C76478 NAND2X1_LOC_522/a_36_24# NOR2X1_LOC_243/B -0.02fF
C76479 NOR2X1_LOC_178/Y INVX1_LOC_42/A 0.05fF
C76480 NOR2X1_LOC_68/A INVX1_LOC_230/A 0.30fF
C76481 NOR2X1_LOC_181/A NOR2X1_LOC_180/Y 0.02fF
C76482 NOR2X1_LOC_540/B NOR2X1_LOC_181/Y 0.09fF
C76483 NOR2X1_LOC_468/Y INVX1_LOC_63/A 0.12fF
C76484 NOR2X1_LOC_349/A INVX1_LOC_210/A 0.41fF
C76485 NOR2X1_LOC_74/A NAND2X1_LOC_392/Y 0.01fF
C76486 NOR2X1_LOC_2/Y INPUT_5 0.04fF
C76487 INVX1_LOC_35/A NAND2X1_LOC_647/B 0.00fF
C76488 NOR2X1_LOC_717/A INVX1_LOC_4/Y 0.10fF
C76489 NOR2X1_LOC_860/B INVX1_LOC_38/A 0.01fF
C76490 NOR2X1_LOC_828/B NOR2X1_LOC_724/Y 4.60fF
C76491 INVX1_LOC_1/A INVX1_LOC_125/A 0.11fF
C76492 INVX1_LOC_83/A NOR2X1_LOC_74/A 0.07fF
C76493 NAND2X1_LOC_72/Y INVX1_LOC_4/A 0.12fF
C76494 NAND2X1_LOC_833/Y INVX1_LOC_33/Y 0.02fF
C76495 NOR2X1_LOC_360/a_36_216# INVX1_LOC_280/A 0.01fF
C76496 NOR2X1_LOC_778/B NOR2X1_LOC_540/B 0.00fF
C76497 NAND2X1_LOC_518/a_36_24# NAND2X1_LOC_96/A 0.00fF
C76498 INVX1_LOC_88/A INVX1_LOC_29/A 0.04fF
C76499 INVX1_LOC_163/A INVX1_LOC_42/A 0.08fF
C76500 INVX1_LOC_174/Y INVX1_LOC_91/A 0.04fF
C76501 INVX1_LOC_165/Y NOR2X1_LOC_124/A 0.20fF
C76502 NOR2X1_LOC_389/A INVX1_LOC_63/A 0.76fF
C76503 INVX1_LOC_14/A NOR2X1_LOC_610/Y 0.04fF
C76504 NOR2X1_LOC_272/Y INVX1_LOC_32/A 0.06fF
C76505 INVX1_LOC_225/Y INVX1_LOC_19/A 0.10fF
C76506 INVX1_LOC_53/A NAND2X1_LOC_425/a_36_24# 0.00fF
C76507 INVX1_LOC_151/Y NAND2X1_LOC_468/B 0.01fF
C76508 INVX1_LOC_89/A NOR2X1_LOC_391/Y 0.03fF
C76509 NOR2X1_LOC_808/A VDD 0.12fF
C76510 NOR2X1_LOC_433/A INVX1_LOC_54/A 8.64fF
C76511 NOR2X1_LOC_329/B INVX1_LOC_67/Y 0.01fF
C76512 NAND2X1_LOC_137/a_36_24# INVX1_LOC_280/A 0.00fF
C76513 INVX1_LOC_11/A NAND2X1_LOC_807/B 0.27fF
C76514 INVX1_LOC_30/A NAND2X1_LOC_476/Y 0.02fF
C76515 NAND2X1_LOC_363/B NOR2X1_LOC_843/B 0.07fF
C76516 INVX1_LOC_249/A INVX1_LOC_179/A 0.01fF
C76517 INVX1_LOC_57/Y NAND2X1_LOC_477/Y 0.37fF
C76518 NOR2X1_LOC_844/A NOR2X1_LOC_865/A 0.07fF
C76519 INVX1_LOC_30/A INVX1_LOC_186/Y 0.03fF
C76520 INVX1_LOC_49/A INVX1_LOC_307/A 0.07fF
C76521 INVX1_LOC_18/A NAND2X1_LOC_475/Y 0.10fF
C76522 INVX1_LOC_289/A VDD -0.00fF
C76523 NAND2X1_LOC_140/A NOR2X1_LOC_139/Y 0.10fF
C76524 INVX1_LOC_11/A NOR2X1_LOC_48/B 0.77fF
C76525 NOR2X1_LOC_569/Y NOR2X1_LOC_35/Y 0.10fF
C76526 NOR2X1_LOC_91/A NAND2X1_LOC_552/A 0.02fF
C76527 INVX1_LOC_64/A INVX1_LOC_50/A 0.15fF
C76528 INVX1_LOC_5/A NOR2X1_LOC_668/Y 0.12fF
C76529 INVX1_LOC_49/A NOR2X1_LOC_445/B 0.13fF
C76530 INVX1_LOC_95/Y INVX1_LOC_306/A 0.01fF
C76531 INVX1_LOC_17/Y NAND2X1_LOC_624/B 0.06fF
C76532 NOR2X1_LOC_78/A INVX1_LOC_196/Y 0.03fF
C76533 NOR2X1_LOC_52/B INVX1_LOC_54/A 0.34fF
C76534 NAND2X1_LOC_117/a_36_24# NAND2X1_LOC_642/Y 0.01fF
C76535 NOR2X1_LOC_441/Y NOR2X1_LOC_89/A 0.08fF
C76536 NAND2X1_LOC_656/A NOR2X1_LOC_814/A 0.47fF
C76537 NOR2X1_LOC_500/B INVX1_LOC_29/A 0.04fF
C76538 NAND2X1_LOC_140/A NAND2X1_LOC_468/B 0.16fF
C76539 INVX1_LOC_16/A NAND2X1_LOC_472/Y 0.02fF
C76540 NAND2X1_LOC_773/Y INVX1_LOC_87/A 0.03fF
C76541 NOR2X1_LOC_15/Y NAND2X1_LOC_223/A 0.03fF
C76542 NAND2X1_LOC_866/B NOR2X1_LOC_823/Y 0.02fF
C76543 NOR2X1_LOC_91/A INVX1_LOC_178/A 0.03fF
C76544 NAND2X1_LOC_563/A INVX1_LOC_280/A 0.12fF
C76545 INVX1_LOC_11/A NAND2X1_LOC_3/B 0.16fF
C76546 NAND2X1_LOC_840/B INVX1_LOC_38/A 0.03fF
C76547 NOR2X1_LOC_92/Y NOR2X1_LOC_301/A 0.16fF
C76548 INVX1_LOC_5/A INVX1_LOC_23/A 7.04fF
C76549 INVX1_LOC_50/Y NOR2X1_LOC_748/A 0.02fF
C76550 INVX1_LOC_208/Y NOR2X1_LOC_536/A 0.00fF
C76551 INVX1_LOC_208/A NOR2X1_LOC_331/B 0.10fF
C76552 INVX1_LOC_35/A NOR2X1_LOC_109/a_36_216# 0.00fF
C76553 INVX1_LOC_2/A INVX1_LOC_307/A 0.07fF
C76554 NAND2X1_LOC_11/Y NOR2X1_LOC_451/A 0.01fF
C76555 NOR2X1_LOC_174/B NOR2X1_LOC_857/A 0.01fF
C76556 NOR2X1_LOC_751/A NOR2X1_LOC_557/A 0.00fF
C76557 NOR2X1_LOC_759/A INVX1_LOC_109/Y 0.00fF
C76558 INVX1_LOC_21/A INVX1_LOC_29/Y 0.29fF
C76559 NAND2X1_LOC_9/Y INVX1_LOC_306/Y 0.09fF
C76560 INVX1_LOC_226/Y INVX1_LOC_118/A 0.01fF
C76561 INVX1_LOC_178/A INVX1_LOC_23/A 0.12fF
C76562 INVX1_LOC_135/A INVX1_LOC_12/Y 0.01fF
C76563 NAND2X1_LOC_357/A NOR2X1_LOC_278/Y 0.00fF
C76564 INVX1_LOC_14/A NAND2X1_LOC_286/B 0.03fF
C76565 INVX1_LOC_217/A NOR2X1_LOC_754/A 0.06fF
C76566 INVX1_LOC_233/A INVX1_LOC_306/Y 0.01fF
C76567 INVX1_LOC_43/A NAND2X1_LOC_93/B 0.04fF
C76568 NAND2X1_LOC_53/Y NOR2X1_LOC_631/Y 0.08fF
C76569 NOR2X1_LOC_770/Y VDD 0.12fF
C76570 INVX1_LOC_303/A INVX1_LOC_29/A 0.07fF
C76571 INVX1_LOC_89/A INVX1_LOC_129/Y 0.00fF
C76572 NOR2X1_LOC_356/A INVX1_LOC_46/A 0.03fF
C76573 INVX1_LOC_110/A INVX1_LOC_15/A 0.03fF
C76574 NOR2X1_LOC_78/B NOR2X1_LOC_865/Y 0.07fF
C76575 INVX1_LOC_49/A INVX1_LOC_12/A 4.10fF
C76576 NAND2X1_LOC_364/A INVX1_LOC_32/A 0.50fF
C76577 NOR2X1_LOC_91/A NAND2X1_LOC_337/B 0.34fF
C76578 NOR2X1_LOC_433/A NAND2X1_LOC_807/B 0.13fF
C76579 INVX1_LOC_25/A NAND2X1_LOC_346/a_36_24# 0.01fF
C76580 NOR2X1_LOC_274/Y INVX1_LOC_42/A 0.06fF
C76581 INVX1_LOC_10/A INVX1_LOC_118/A 0.13fF
C76582 NAND2X1_LOC_59/B INVX1_LOC_29/A 0.05fF
C76583 NOR2X1_LOC_91/A NOR2X1_LOC_816/A 0.64fF
C76584 NAND2X1_LOC_364/A NOR2X1_LOC_623/B 0.08fF
C76585 NOR2X1_LOC_196/A INVX1_LOC_15/A 0.01fF
C76586 NOR2X1_LOC_356/A NAND2X1_LOC_417/a_36_24# 0.00fF
C76587 INVX1_LOC_28/A NAND2X1_LOC_472/Y 0.08fF
C76588 NAND2X1_LOC_860/A INVX1_LOC_14/A 0.45fF
C76589 INVX1_LOC_148/A INVX1_LOC_117/A 0.01fF
C76590 NOR2X1_LOC_433/A NOR2X1_LOC_48/B 0.05fF
C76591 NOR2X1_LOC_590/A NAND2X1_LOC_99/A 0.03fF
C76592 INVX1_LOC_22/A INVX1_LOC_113/A 0.02fF
C76593 INVX1_LOC_237/Y INVX1_LOC_42/A 0.02fF
C76594 NOR2X1_LOC_142/Y NOR2X1_LOC_89/A 0.09fF
C76595 NOR2X1_LOC_846/Y NOR2X1_LOC_846/A 0.02fF
C76596 INVX1_LOC_266/Y INVX1_LOC_19/A 0.17fF
C76597 NOR2X1_LOC_205/Y NOR2X1_LOC_717/A 0.51fF
C76598 NAND2X1_LOC_67/Y NOR2X1_LOC_665/a_36_216# 0.02fF
C76599 INVX1_LOC_28/A NAND2X1_LOC_603/a_36_24# 0.00fF
C76600 NOR2X1_LOC_74/A INVX1_LOC_46/A 0.29fF
C76601 NAND2X1_LOC_337/B INVX1_LOC_23/A 0.08fF
C76602 NOR2X1_LOC_816/A INVX1_LOC_23/A 0.00fF
C76603 INVX1_LOC_96/A NOR2X1_LOC_486/Y 0.03fF
C76604 NOR2X1_LOC_45/B INVX1_LOC_187/A 0.03fF
C76605 NOR2X1_LOC_175/A NOR2X1_LOC_633/A 0.51fF
C76606 D_INPUT_0 INVX1_LOC_92/A 0.07fF
C76607 INVX1_LOC_30/A NOR2X1_LOC_843/B 0.00fF
C76608 NOR2X1_LOC_9/Y INVX1_LOC_46/A 0.08fF
C76609 NAND2X1_LOC_858/B NAND2X1_LOC_721/A 0.02fF
C76610 INVX1_LOC_2/A INVX1_LOC_12/A 0.29fF
C76611 INVX1_LOC_256/Y NAND2X1_LOC_81/B 0.07fF
C76612 INVX1_LOC_120/A NAND2X1_LOC_60/a_36_24# 0.00fF
C76613 NOR2X1_LOC_135/Y INVX1_LOC_9/A 0.01fF
C76614 INVX1_LOC_16/A NAND2X1_LOC_773/B 0.27fF
C76615 NOR2X1_LOC_655/B NOR2X1_LOC_89/A 0.03fF
C76616 NOR2X1_LOC_226/A INVX1_LOC_12/A 0.14fF
C76617 NAND2X1_LOC_739/B NOR2X1_LOC_829/A 0.06fF
C76618 INVX1_LOC_83/A NOR2X1_LOC_243/B 0.07fF
C76619 NOR2X1_LOC_337/Y INVX1_LOC_37/A 0.02fF
C76620 NOR2X1_LOC_741/A INVX1_LOC_139/Y 0.01fF
C76621 INVX1_LOC_72/A INVX1_LOC_57/A 1.07fF
C76622 INPUT_3 INVX1_LOC_138/Y 0.03fF
C76623 NOR2X1_LOC_368/A NOR2X1_LOC_271/Y 0.10fF
C76624 INVX1_LOC_50/A INVX1_LOC_130/Y 0.03fF
C76625 INVX1_LOC_64/A INVX1_LOC_61/Y 0.02fF
C76626 INVX1_LOC_58/A NAND2X1_LOC_16/Y 0.00fF
C76627 NOR2X1_LOC_453/a_36_216# NOR2X1_LOC_453/Y 0.00fF
C76628 INVX1_LOC_121/A NOR2X1_LOC_257/Y 0.02fF
C76629 NOR2X1_LOC_187/Y NOR2X1_LOC_348/Y 0.02fF
C76630 INVX1_LOC_1/A NOR2X1_LOC_140/A 0.07fF
C76631 NOR2X1_LOC_456/Y INVX1_LOC_136/A 0.13fF
C76632 NOR2X1_LOC_268/a_36_216# INVX1_LOC_271/A 0.00fF
C76633 NAND2X1_LOC_552/A INVX1_LOC_31/A 0.03fF
C76634 INVX1_LOC_20/Y NAND2X1_LOC_574/A 0.02fF
C76635 NOR2X1_LOC_396/Y VDD 0.25fF
C76636 NOR2X1_LOC_500/A NOR2X1_LOC_383/B 5.15fF
C76637 NOR2X1_LOC_65/B NOR2X1_LOC_274/Y -0.00fF
C76638 INVX1_LOC_5/A INVX1_LOC_31/A 0.42fF
C76639 NAND2X1_LOC_352/B NOR2X1_LOC_652/Y 0.13fF
C76640 NOR2X1_LOC_627/Y INVX1_LOC_32/A 0.00fF
C76641 INVX1_LOC_45/Y INVX1_LOC_271/A 0.02fF
C76642 NOR2X1_LOC_303/Y NOR2X1_LOC_383/B 0.03fF
C76643 INVX1_LOC_200/Y INVX1_LOC_41/Y 0.00fF
C76644 NAND2X1_LOC_787/A INVX1_LOC_18/A 0.03fF
C76645 INVX1_LOC_59/A NOR2X1_LOC_82/A 0.63fF
C76646 INVX1_LOC_17/A NOR2X1_LOC_92/Y 0.15fF
C76647 INVX1_LOC_104/A INVX1_LOC_94/Y 0.01fF
C76648 NOR2X1_LOC_631/B VDD 0.24fF
C76649 INVX1_LOC_64/A NOR2X1_LOC_659/a_36_216# 0.01fF
C76650 INVX1_LOC_17/Y NOR2X1_LOC_617/Y 0.06fF
C76651 NOR2X1_LOC_56/Y INVX1_LOC_37/A 0.03fF
C76652 INVX1_LOC_222/Y NOR2X1_LOC_590/A 0.03fF
C76653 INVX1_LOC_80/A INVX1_LOC_29/A 0.01fF
C76654 NAND2X1_LOC_569/B NOR2X1_LOC_384/Y 0.09fF
C76655 INVX1_LOC_215/Y NOR2X1_LOC_321/Y 0.28fF
C76656 NAND2X1_LOC_462/B INVX1_LOC_12/A 0.00fF
C76657 NOR2X1_LOC_405/A INVX1_LOC_66/Y 0.06fF
C76658 INVX1_LOC_256/A NOR2X1_LOC_187/Y 0.27fF
C76659 NAND2X1_LOC_84/Y NAND2X1_LOC_860/A 0.01fF
C76660 NOR2X1_LOC_78/B NOR2X1_LOC_855/A 0.03fF
C76661 NAND2X1_LOC_477/A NOR2X1_LOC_301/A 0.03fF
C76662 INVX1_LOC_57/Y INVX1_LOC_93/A 0.10fF
C76663 INVX1_LOC_63/Y INVX1_LOC_270/A 0.08fF
C76664 INVX1_LOC_146/Y INVX1_LOC_37/A 0.00fF
C76665 NOR2X1_LOC_52/B NOR2X1_LOC_438/Y 0.03fF
C76666 NOR2X1_LOC_681/Y VDD 0.03fF
C76667 INVX1_LOC_90/A INVX1_LOC_49/Y 0.03fF
C76668 NAND2X1_LOC_472/Y NOR2X1_LOC_35/Y 0.10fF
C76669 NOR2X1_LOC_486/Y NOR2X1_LOC_684/Y 0.45fF
C76670 VDD INVX1_LOC_37/A 2.21fF
C76671 NOR2X1_LOC_703/Y NOR2X1_LOC_809/B 0.01fF
C76672 NOR2X1_LOC_45/B NOR2X1_LOC_629/Y 0.03fF
C76673 NAND2X1_LOC_787/A INVX1_LOC_172/A 0.03fF
C76674 NAND2X1_LOC_182/A INVX1_LOC_181/A 0.29fF
C76675 NOR2X1_LOC_34/B NOR2X1_LOC_554/B 0.03fF
C76676 VDD NOR2X1_LOC_231/A -0.00fF
C76677 INVX1_LOC_28/A NAND2X1_LOC_773/B 0.14fF
C76678 INVX1_LOC_97/A INVX1_LOC_99/A 0.01fF
C76679 NOR2X1_LOC_332/A NOR2X1_LOC_847/a_36_216# 0.01fF
C76680 NAND2X1_LOC_648/A INVX1_LOC_12/A 0.12fF
C76681 INVX1_LOC_11/A NAND2X1_LOC_350/A 0.07fF
C76682 INVX1_LOC_64/A INVX1_LOC_105/A 0.01fF
C76683 NOR2X1_LOC_6/B NOR2X1_LOC_748/A 0.02fF
C76684 NOR2X1_LOC_241/A NOR2X1_LOC_785/A 0.00fF
C76685 INPUT_1 INVX1_LOC_12/A 0.11fF
C76686 INVX1_LOC_224/A INVX1_LOC_218/Y 0.25fF
C76687 NAND2X1_LOC_350/B NOR2X1_LOC_449/A 0.02fF
C76688 INVX1_LOC_199/A INVX1_LOC_54/A 0.03fF
C76689 NOR2X1_LOC_71/Y INVX1_LOC_170/Y 0.01fF
C76690 NOR2X1_LOC_598/B NOR2X1_LOC_770/B 0.00fF
C76691 INVX1_LOC_90/A NOR2X1_LOC_672/a_36_216# 0.00fF
C76692 NAND2X1_LOC_562/B INVX1_LOC_23/A 0.01fF
C76693 INVX1_LOC_65/A NOR2X1_LOC_640/Y 0.10fF
C76694 INVX1_LOC_54/Y NOR2X1_LOC_383/B 0.07fF
C76695 INVX1_LOC_37/A NOR2X1_LOC_684/a_36_216# 0.00fF
C76696 INVX1_LOC_11/A NOR2X1_LOC_441/Y 0.03fF
C76697 NOR2X1_LOC_658/Y NOR2X1_LOC_205/Y 0.01fF
C76698 NOR2X1_LOC_813/Y INVX1_LOC_12/Y 0.75fF
C76699 NOR2X1_LOC_331/B NAND2X1_LOC_211/Y 0.07fF
C76700 NOR2X1_LOC_349/A NOR2X1_LOC_259/B 0.04fF
C76701 INVX1_LOC_277/A NOR2X1_LOC_739/Y 0.19fF
C76702 NOR2X1_LOC_91/A NOR2X1_LOC_773/Y 0.42fF
C76703 INVX1_LOC_25/A NOR2X1_LOC_709/A 0.24fF
C76704 INVX1_LOC_50/A INVX1_LOC_44/Y 0.01fF
C76705 INVX1_LOC_136/A NAND2X1_LOC_561/B 0.09fF
C76706 NOR2X1_LOC_537/Y INVX1_LOC_57/A 0.07fF
C76707 NOR2X1_LOC_816/A INVX1_LOC_31/A 0.16fF
C76708 NAND2X1_LOC_854/B INVX1_LOC_94/Y 0.02fF
C76709 NAND2X1_LOC_338/B INVX1_LOC_57/A 0.25fF
C76710 INVX1_LOC_50/A NAND2X1_LOC_850/Y 0.00fF
C76711 INVX1_LOC_12/Y INVX1_LOC_280/A 0.01fF
C76712 NOR2X1_LOC_379/Y NOR2X1_LOC_460/Y 0.05fF
C76713 NAND2X1_LOC_469/B NOR2X1_LOC_435/A 0.02fF
C76714 NOR2X1_LOC_188/A INVX1_LOC_125/A 0.10fF
C76715 VDD INVX1_LOC_157/Y 0.27fF
C76716 INPUT_5 NOR2X1_LOC_36/A 0.25fF
C76717 INVX1_LOC_48/A NOR2X1_LOC_721/B 0.03fF
C76718 NAND2X1_LOC_323/B INVX1_LOC_57/A 12.39fF
C76719 INVX1_LOC_291/A INVX1_LOC_76/A 0.10fF
C76720 NAND2X1_LOC_391/Y NOR2X1_LOC_716/B 0.01fF
C76721 NOR2X1_LOC_548/B INVX1_LOC_125/A 0.10fF
C76722 NOR2X1_LOC_567/B NOR2X1_LOC_640/B 0.08fF
C76723 VDD NOR2X1_LOC_177/Y 0.13fF
C76724 NOR2X1_LOC_773/Y INVX1_LOC_23/A 0.07fF
C76725 NAND2X1_LOC_802/Y INVX1_LOC_76/A 0.07fF
C76726 NAND2X1_LOC_361/Y NOR2X1_LOC_852/Y 0.15fF
C76727 INVX1_LOC_13/Y INVX1_LOC_8/A 0.16fF
C76728 INVX1_LOC_13/Y NAND2X1_LOC_399/a_36_24# 0.01fF
C76729 VDD NOR2X1_LOC_743/Y 0.32fF
C76730 NOR2X1_LOC_530/Y NOR2X1_LOC_384/Y 0.02fF
C76731 INVX1_LOC_35/A NAND2X1_LOC_342/Y 0.02fF
C76732 D_INPUT_7 INVX1_LOC_174/A 0.03fF
C76733 INVX1_LOC_180/Y NAND2X1_LOC_453/A 0.01fF
C76734 INVX1_LOC_232/Y NOR2X1_LOC_392/Y 0.00fF
C76735 INVX1_LOC_28/A NOR2X1_LOC_393/Y 0.02fF
C76736 NAND2X1_LOC_357/B NOR2X1_LOC_652/Y 0.01fF
C76737 NOR2X1_LOC_682/Y INVX1_LOC_92/A 0.01fF
C76738 NOR2X1_LOC_91/A NAND2X1_LOC_317/a_36_24# 0.01fF
C76739 NOR2X1_LOC_15/Y INVX1_LOC_33/A 0.06fF
C76740 NOR2X1_LOC_596/Y NOR2X1_LOC_457/B 0.01fF
C76741 NOR2X1_LOC_790/B NOR2X1_LOC_553/Y 0.05fF
C76742 NOR2X1_LOC_791/Y INVX1_LOC_34/Y 0.01fF
C76743 NOR2X1_LOC_35/Y NAND2X1_LOC_206/Y 0.10fF
C76744 NAND2X1_LOC_660/Y INVX1_LOC_53/A 0.03fF
C76745 NOR2X1_LOC_590/A NAND2X1_LOC_656/A 0.01fF
C76746 INVX1_LOC_30/A INVX1_LOC_18/A 9.36fF
C76747 INVX1_LOC_202/A NOR2X1_LOC_276/Y 0.04fF
C76748 INVX1_LOC_17/A INVX1_LOC_41/A 0.03fF
C76749 INVX1_LOC_14/A NOR2X1_LOC_516/Y 0.02fF
C76750 NAND2X1_LOC_350/A NOR2X1_LOC_433/A 0.69fF
C76751 D_INPUT_1 NOR2X1_LOC_128/B 0.03fF
C76752 INVX1_LOC_299/A INVX1_LOC_104/A 0.07fF
C76753 NAND2X1_LOC_763/B INVX1_LOC_18/A 0.04fF
C76754 INVX1_LOC_11/A NOR2X1_LOC_340/Y 0.02fF
C76755 NAND2X1_LOC_569/A NOR2X1_LOC_103/Y 0.02fF
C76756 INVX1_LOC_221/A NAND2X1_LOC_538/Y 0.03fF
C76757 INVX1_LOC_291/Y NOR2X1_LOC_89/A 0.03fF
C76758 NOR2X1_LOC_795/Y INVX1_LOC_269/A 0.10fF
C76759 INVX1_LOC_1/A NOR2X1_LOC_709/A 0.20fF
C76760 NOR2X1_LOC_337/A INVX1_LOC_4/Y 0.08fF
C76761 NAND2X1_LOC_39/a_36_24# NOR2X1_LOC_596/A 0.00fF
C76762 INVX1_LOC_255/Y NAND2X1_LOC_214/B 0.24fF
C76763 D_INPUT_0 INVX1_LOC_53/A 0.31fF
C76764 NOR2X1_LOC_441/Y NOR2X1_LOC_433/A 0.09fF
C76765 INVX1_LOC_313/Y INVX1_LOC_57/A 0.01fF
C76766 INVX1_LOC_39/A INVX1_LOC_226/Y 0.08fF
C76767 NOR2X1_LOC_506/Y NOR2X1_LOC_510/B 0.06fF
C76768 INVX1_LOC_17/A NAND2X1_LOC_477/A 0.10fF
C76769 INVX1_LOC_5/A NAND2X1_LOC_859/Y 0.00fF
C76770 NOR2X1_LOC_91/A INVX1_LOC_140/A 0.16fF
C76771 INVX1_LOC_174/A INVX1_LOC_192/A 0.01fF
C76772 INVX1_LOC_172/A INVX1_LOC_30/A 0.06fF
C76773 NOR2X1_LOC_20/Y INVX1_LOC_15/Y 0.05fF
C76774 INVX1_LOC_230/Y NOR2X1_LOC_297/a_36_216# 0.00fF
C76775 INVX1_LOC_201/Y NAND2X1_LOC_555/Y 1.07fF
C76776 NAND2X1_LOC_350/A NOR2X1_LOC_52/B 0.07fF
C76777 INVX1_LOC_2/A INVX1_LOC_200/A 0.07fF
C76778 NAND2X1_LOC_736/Y INVX1_LOC_284/Y 0.07fF
C76779 INVX1_LOC_21/A INVX1_LOC_101/A 0.03fF
C76780 INVX1_LOC_45/A INVX1_LOC_155/A 0.04fF
C76781 NOR2X1_LOC_405/A INVX1_LOC_32/A 1.11fF
C76782 NOR2X1_LOC_15/Y INVX1_LOC_40/A 0.08fF
C76783 INVX1_LOC_254/A NOR2X1_LOC_68/A 0.03fF
C76784 NOR2X1_LOC_357/Y INVX1_LOC_109/Y 0.15fF
C76785 NOR2X1_LOC_337/Y NAND2X1_LOC_72/B 0.01fF
C76786 NOR2X1_LOC_614/Y INVX1_LOC_269/A 0.01fF
C76787 NOR2X1_LOC_226/A INVX1_LOC_200/A 0.11fF
C76788 INVX1_LOC_88/A INVX1_LOC_151/Y 0.01fF
C76789 NOR2X1_LOC_441/Y NOR2X1_LOC_52/B 0.24fF
C76790 INVX1_LOC_245/Y NOR2X1_LOC_78/B 0.03fF
C76791 INVX1_LOC_41/Y NOR2X1_LOC_495/Y 0.01fF
C76792 NOR2X1_LOC_848/Y NOR2X1_LOC_516/B 1.16fF
C76793 INVX1_LOC_11/A NAND2X1_LOC_553/a_36_24# 0.01fF
C76794 NOR2X1_LOC_632/Y NAND2X1_LOC_67/Y 0.02fF
C76795 INVX1_LOC_38/A INVX1_LOC_49/Y 0.11fF
C76796 INVX1_LOC_21/A NOR2X1_LOC_355/A 0.03fF
C76797 INVX1_LOC_89/A INVX1_LOC_50/Y 0.20fF
C76798 NOR2X1_LOC_446/A NAND2X1_LOC_372/a_36_24# 0.00fF
C76799 INVX1_LOC_64/A NAND2X1_LOC_652/Y 0.02fF
C76800 INVX1_LOC_27/A NOR2X1_LOC_71/Y 0.01fF
C76801 NAND2X1_LOC_552/A NAND2X1_LOC_807/Y 0.00fF
C76802 NOR2X1_LOC_824/A NOR2X1_LOC_71/Y 0.02fF
C76803 INVX1_LOC_256/A INVX1_LOC_208/Y 0.07fF
C76804 NOR2X1_LOC_405/A NAND2X1_LOC_175/Y 0.24fF
C76805 NOR2X1_LOC_528/Y NOR2X1_LOC_693/Y 0.20fF
C76806 INVX1_LOC_315/Y NAND2X1_LOC_222/a_36_24# 0.00fF
C76807 NAND2X1_LOC_357/a_36_24# INVX1_LOC_162/A 0.00fF
C76808 NOR2X1_LOC_285/A NOR2X1_LOC_334/A 0.01fF
C76809 NOR2X1_LOC_623/B NOR2X1_LOC_857/A 0.07fF
C76810 NAND2X1_LOC_508/A INVX1_LOC_50/Y 0.05fF
C76811 INVX1_LOC_155/A INVX1_LOC_71/A 0.04fF
C76812 NOR2X1_LOC_773/Y INVX1_LOC_31/A 0.07fF
C76813 NAND2X1_LOC_773/Y INVX1_LOC_306/A 0.32fF
C76814 INVX1_LOC_124/Y NOR2X1_LOC_78/B 0.46fF
C76815 NOR2X1_LOC_601/a_36_216# NOR2X1_LOC_151/Y 0.00fF
C76816 INVX1_LOC_181/Y INVX1_LOC_162/Y 0.69fF
C76817 NOR2X1_LOC_208/Y INVX1_LOC_63/Y 0.33fF
C76818 INVX1_LOC_233/A NOR2X1_LOC_74/A 0.02fF
C76819 INVX1_LOC_135/A NOR2X1_LOC_793/A 0.68fF
C76820 NOR2X1_LOC_647/a_36_216# NOR2X1_LOC_516/B 0.00fF
C76821 INVX1_LOC_11/A NAND2X1_LOC_358/Y 0.01fF
C76822 D_INPUT_1 NAND2X1_LOC_473/a_36_24# 0.00fF
C76823 INVX1_LOC_12/A INVX1_LOC_118/A 0.68fF
C76824 INVX1_LOC_91/A NOR2X1_LOC_654/A 0.10fF
C76825 INVX1_LOC_133/A NOR2X1_LOC_743/Y 0.00fF
C76826 INVX1_LOC_178/A NAND2X1_LOC_807/Y 0.10fF
C76827 INVX1_LOC_178/Y NAND2X1_LOC_618/Y 0.14fF
C76828 NOR2X1_LOC_389/A INVX1_LOC_1/Y 0.00fF
C76829 NOR2X1_LOC_391/Y NOR2X1_LOC_392/Y 0.08fF
C76830 NOR2X1_LOC_433/A NOR2X1_LOC_142/Y 0.37fF
C76831 INVX1_LOC_88/A NAND2X1_LOC_140/A 0.03fF
C76832 INVX1_LOC_303/A INVX1_LOC_8/A 0.06fF
C76833 INVX1_LOC_233/A NOR2X1_LOC_9/Y 0.38fF
C76834 NOR2X1_LOC_78/B NOR2X1_LOC_791/A 0.00fF
C76835 NOR2X1_LOC_331/B NAND2X1_LOC_791/a_36_24# 0.01fF
C76836 VDD NAND2X1_LOC_72/B 0.51fF
C76837 NOR2X1_LOC_226/A NAND2X1_LOC_355/Y 0.02fF
C76838 NOR2X1_LOC_471/Y INVX1_LOC_121/A 0.00fF
C76839 INVX1_LOC_215/Y NOR2X1_LOC_686/B 0.05fF
C76840 INVX1_LOC_34/A NOR2X1_LOC_772/Y 0.06fF
C76841 NAND2X1_LOC_288/A INVX1_LOC_19/A 0.16fF
C76842 NAND2X1_LOC_778/Y NOR2X1_LOC_323/Y 0.19fF
C76843 INVX1_LOC_135/A NAND2X1_LOC_550/A 0.10fF
C76844 NAND2X1_LOC_717/Y INVX1_LOC_24/A 0.03fF
C76845 NOR2X1_LOC_58/Y INVX1_LOC_272/A 0.03fF
C76846 NOR2X1_LOC_798/A NOR2X1_LOC_74/A 0.06fF
C76847 NOR2X1_LOC_92/Y NOR2X1_LOC_171/Y 0.03fF
C76848 INVX1_LOC_91/A INVX1_LOC_58/Y 0.11fF
C76849 INVX1_LOC_5/A INVX1_LOC_6/A 0.92fF
C76850 INVX1_LOC_135/A NOR2X1_LOC_160/B 0.14fF
C76851 INVX1_LOC_200/A INPUT_1 0.05fF
C76852 NOR2X1_LOC_691/B NOR2X1_LOC_814/A 0.03fF
C76853 NAND2X1_LOC_530/a_36_24# INVX1_LOC_22/A 0.01fF
C76854 INVX1_LOC_31/A NOR2X1_LOC_332/A 3.67fF
C76855 NOR2X1_LOC_599/Y NAND2X1_LOC_809/A 0.01fF
C76856 NOR2X1_LOC_798/A NOR2X1_LOC_9/Y 0.02fF
C76857 INVX1_LOC_295/A NOR2X1_LOC_160/B 0.06fF
C76858 NOR2X1_LOC_653/Y INVX1_LOC_19/A 0.01fF
C76859 NOR2X1_LOC_142/Y NOR2X1_LOC_52/B 0.27fF
C76860 INVX1_LOC_84/A INVX1_LOC_264/A 0.06fF
C76861 NOR2X1_LOC_67/A INVX1_LOC_77/A 0.00fF
C76862 INVX1_LOC_178/A INVX1_LOC_6/A 0.10fF
C76863 INVX1_LOC_11/A INVX1_LOC_182/A 0.07fF
C76864 NAND2X1_LOC_231/Y NOR2X1_LOC_172/Y 0.03fF
C76865 INVX1_LOC_24/A INVX1_LOC_16/A 1.34fF
C76866 INVX1_LOC_81/A NOR2X1_LOC_131/Y 0.01fF
C76867 NOR2X1_LOC_191/B INVX1_LOC_53/Y 0.02fF
C76868 NOR2X1_LOC_655/B NOR2X1_LOC_593/Y 0.01fF
C76869 NAND2X1_LOC_303/Y NOR2X1_LOC_2/Y 0.05fF
C76870 NAND2X1_LOC_803/B NOR2X1_LOC_329/B 0.02fF
C76871 NOR2X1_LOC_816/A NAND2X1_LOC_807/Y 0.07fF
C76872 NOR2X1_LOC_778/B NOR2X1_LOC_570/B 0.06fF
C76873 INVX1_LOC_33/A INVX1_LOC_226/A 0.01fF
C76874 D_GATE_222 INVX1_LOC_49/A 0.00fF
C76875 NAND2X1_LOC_656/Y NOR2X1_LOC_360/Y 0.63fF
C76876 NOR2X1_LOC_590/A NOR2X1_LOC_329/B 0.19fF
C76877 INVX1_LOC_304/Y INVX1_LOC_2/A 0.03fF
C76878 INVX1_LOC_77/A NOR2X1_LOC_162/a_36_216# 0.00fF
C76879 INVX1_LOC_208/A NOR2X1_LOC_388/Y 0.10fF
C76880 NOR2X1_LOC_667/A NAND2X1_LOC_840/a_36_24# 0.01fF
C76881 NOR2X1_LOC_772/a_36_216# NOR2X1_LOC_772/Y 0.02fF
C76882 INVX1_LOC_31/A INVX1_LOC_140/A 0.07fF
C76883 INVX1_LOC_17/A NAND2X1_LOC_309/a_36_24# 0.00fF
C76884 NOR2X1_LOC_557/Y INVX1_LOC_16/A 0.72fF
C76885 NOR2X1_LOC_553/Y NOR2X1_LOC_344/A 0.06fF
C76886 INVX1_LOC_272/A INVX1_LOC_29/A 0.07fF
C76887 INVX1_LOC_304/Y NOR2X1_LOC_226/A 0.03fF
C76888 NOR2X1_LOC_808/A INVX1_LOC_177/A 0.00fF
C76889 NOR2X1_LOC_577/a_36_216# NOR2X1_LOC_577/Y 0.02fF
C76890 NOR2X1_LOC_529/Y NAND2X1_LOC_549/B 0.00fF
C76891 INVX1_LOC_12/A NAND2X1_LOC_63/Y 0.02fF
C76892 NAND2X1_LOC_228/a_36_24# INVX1_LOC_34/A 0.00fF
C76893 NOR2X1_LOC_295/Y INVX1_LOC_1/Y 0.03fF
C76894 INVX1_LOC_2/A INVX1_LOC_214/Y 0.03fF
C76895 NOR2X1_LOC_160/B NOR2X1_LOC_391/B 0.03fF
C76896 INVX1_LOC_255/Y NOR2X1_LOC_664/Y 0.57fF
C76897 NOR2X1_LOC_639/B NAND2X1_LOC_639/A 0.02fF
C76898 INVX1_LOC_36/A INVX1_LOC_302/Y 0.01fF
C76899 NAND2X1_LOC_164/a_36_24# NAND2X1_LOC_323/B 0.01fF
C76900 NOR2X1_LOC_468/Y INVX1_LOC_93/Y 0.02fF
C76901 INVX1_LOC_89/A NOR2X1_LOC_559/B 0.01fF
C76902 NOR2X1_LOC_506/Y INVX1_LOC_57/A 0.01fF
C76903 INVX1_LOC_59/A INVX1_LOC_59/Y 0.00fF
C76904 NOR2X1_LOC_478/a_36_216# INVX1_LOC_34/A 0.02fF
C76905 NOR2X1_LOC_15/Y NOR2X1_LOC_486/Y 0.19fF
C76906 NAND2X1_LOC_562/B NAND2X1_LOC_859/Y 0.00fF
C76907 NAND2X1_LOC_785/A NAND2X1_LOC_564/B 0.35fF
C76908 NOR2X1_LOC_510/Y INVX1_LOC_37/A 0.03fF
C76909 NOR2X1_LOC_831/B NOR2X1_LOC_318/A 0.46fF
C76910 INVX1_LOC_122/Y INVX1_LOC_75/A 0.43fF
C76911 INVX1_LOC_24/A INVX1_LOC_28/A 1.37fF
C76912 NAND2X1_LOC_391/Y NAND2X1_LOC_633/Y 0.04fF
C76913 INVX1_LOC_45/A INVX1_LOC_86/A 0.04fF
C76914 INVX1_LOC_255/Y NAND2X1_LOC_570/Y 0.04fF
C76915 INVX1_LOC_58/A NOR2X1_LOC_433/Y 0.05fF
C76916 INVX1_LOC_135/A NOR2X1_LOC_523/a_36_216# 0.00fF
C76917 INVX1_LOC_208/A NOR2X1_LOC_366/B 0.00fF
C76918 INVX1_LOC_21/A NOR2X1_LOC_111/A 0.09fF
C76919 NOR2X1_LOC_389/A NOR2X1_LOC_318/B 0.10fF
C76920 NOR2X1_LOC_742/A NOR2X1_LOC_596/A 0.08fF
C76921 NOR2X1_LOC_264/Y NOR2X1_LOC_749/Y 0.05fF
C76922 INVX1_LOC_34/A INVX1_LOC_90/A 0.08fF
C76923 NAND2X1_LOC_53/Y NAND2X1_LOC_212/Y 0.02fF
C76924 NOR2X1_LOC_78/B NAND2X1_LOC_660/Y 0.14fF
C76925 NAND2X1_LOC_559/Y VDD 0.01fF
C76926 NOR2X1_LOC_445/Y INVX1_LOC_55/Y 0.00fF
C76927 INVX1_LOC_89/A NOR2X1_LOC_6/B 0.30fF
C76928 INVX1_LOC_34/A NOR2X1_LOC_389/B 0.07fF
C76929 NAND2X1_LOC_477/Y NOR2X1_LOC_693/Y 0.06fF
C76930 INVX1_LOC_2/A NAND2X1_LOC_808/A 0.08fF
C76931 NAND2X1_LOC_565/B INVX1_LOC_16/A 0.02fF
C76932 INVX1_LOC_84/A NOR2X1_LOC_646/B 0.05fF
C76933 NAND2X1_LOC_357/A NAND2X1_LOC_287/B 0.02fF
C76934 NAND2X1_LOC_9/Y NOR2X1_LOC_865/Y 0.04fF
C76935 NOR2X1_LOC_226/A NAND2X1_LOC_808/A 0.07fF
C76936 INVX1_LOC_171/A NOR2X1_LOC_767/a_36_216# 0.00fF
C76937 D_INPUT_0 NOR2X1_LOC_547/B 0.02fF
C76938 D_INPUT_0 NOR2X1_LOC_78/B 0.41fF
C76939 NAND2X1_LOC_53/Y INVX1_LOC_14/Y 0.10fF
C76940 NOR2X1_LOC_200/a_36_216# D_GATE_366 0.02fF
C76941 INVX1_LOC_295/A INVX1_LOC_189/A 0.03fF
C76942 NOR2X1_LOC_841/a_36_216# NAND2X1_LOC_175/Y 0.00fF
C76943 INVX1_LOC_26/Y INVX1_LOC_19/A 0.21fF
C76944 NOR2X1_LOC_816/a_36_216# INVX1_LOC_54/A 0.00fF
C76945 INVX1_LOC_185/A NOR2X1_LOC_406/A 0.00fF
C76946 NAND2X1_LOC_214/B INVX1_LOC_89/Y 0.01fF
C76947 INVX1_LOC_27/A NAND2X1_LOC_698/a_36_24# 0.06fF
C76948 INVX1_LOC_36/A NOR2X1_LOC_823/Y 0.00fF
C76949 INVX1_LOC_90/A NAND2X1_LOC_231/Y 0.01fF
C76950 INVX1_LOC_34/A NAND2X1_LOC_348/A 0.00fF
C76951 INVX1_LOC_232/A NOR2X1_LOC_719/B 0.01fF
C76952 INVX1_LOC_314/Y INVX1_LOC_286/A 0.01fF
C76953 NOR2X1_LOC_598/B NOR2X1_LOC_673/A 0.10fF
C76954 NAND2X1_LOC_638/Y NAND2X1_LOC_451/Y 0.14fF
C76955 INVX1_LOC_35/A INVX1_LOC_285/A 0.10fF
C76956 INVX1_LOC_135/A NOR2X1_LOC_516/B 0.08fF
C76957 NAND2X1_LOC_800/Y INVX1_LOC_16/A 0.13fF
C76958 NOR2X1_LOC_824/A NAND2X1_LOC_243/Y 0.02fF
C76959 NOR2X1_LOC_147/B INPUT_0 0.12fF
C76960 NOR2X1_LOC_312/Y INVX1_LOC_25/Y 0.14fF
C76961 NOR2X1_LOC_130/A INVX1_LOC_16/A 0.07fF
C76962 INVX1_LOC_88/A INVX1_LOC_118/Y 0.06fF
C76963 NOR2X1_LOC_793/Y INVX1_LOC_9/A 0.12fF
C76964 INVX1_LOC_35/A NOR2X1_LOC_814/A 1.20fF
C76965 NAND2X1_LOC_551/a_36_24# INVX1_LOC_19/A 0.00fF
C76966 NOR2X1_LOC_392/B INPUT_0 0.01fF
C76967 NOR2X1_LOC_168/B NOR2X1_LOC_567/B 0.07fF
C76968 INVX1_LOC_191/Y INVX1_LOC_140/A 0.03fF
C76969 NOR2X1_LOC_662/A NAND2X1_LOC_793/B 0.07fF
C76970 NOR2X1_LOC_13/Y NOR2X1_LOC_595/Y 0.00fF
C76971 NOR2X1_LOC_158/Y INVX1_LOC_15/A 0.07fF
C76972 NOR2X1_LOC_91/A INVX1_LOC_42/A 0.12fF
C76973 NOR2X1_LOC_295/a_36_216# INVX1_LOC_69/Y 0.00fF
C76974 NOR2X1_LOC_419/Y INVX1_LOC_91/A 1.59fF
C76975 NOR2X1_LOC_773/Y NAND2X1_LOC_807/Y 0.01fF
C76976 NAND2X1_LOC_198/B NOR2X1_LOC_56/Y 0.03fF
C76977 INVX1_LOC_30/Y INVX1_LOC_89/A 0.03fF
C76978 NOR2X1_LOC_716/B INVX1_LOC_91/A 0.17fF
C76979 INVX1_LOC_286/Y INVX1_LOC_77/Y 0.06fF
C76980 INVX1_LOC_200/A INVX1_LOC_118/A 0.06fF
C76981 NOR2X1_LOC_160/B INVX1_LOC_280/A 0.07fF
C76982 NAND2X1_LOC_303/Y NOR2X1_LOC_695/a_36_216# 0.15fF
C76983 NOR2X1_LOC_361/B NOR2X1_LOC_743/Y 0.27fF
C76984 NOR2X1_LOC_220/A NOR2X1_LOC_742/A 0.14fF
C76985 INVX1_LOC_24/A NOR2X1_LOC_253/Y 0.04fF
C76986 NAND2X1_LOC_565/B INVX1_LOC_28/A 0.00fF
C76987 D_INPUT_0 INVX1_LOC_83/A 0.25fF
C76988 INVX1_LOC_24/A NOR2X1_LOC_35/Y 0.43fF
C76989 INVX1_LOC_207/Y NOR2X1_LOC_32/Y 0.04fF
C76990 INVX1_LOC_269/A NOR2X1_LOC_862/B 0.10fF
C76991 INVX1_LOC_23/A INVX1_LOC_42/A 0.11fF
C76992 INVX1_LOC_308/A NOR2X1_LOC_89/A 0.00fF
C76993 INVX1_LOC_255/Y NOR2X1_LOC_19/B 0.14fF
C76994 NOR2X1_LOC_733/a_36_216# INVX1_LOC_139/Y 0.00fF
C76995 NOR2X1_LOC_295/Y NOR2X1_LOC_318/B 0.07fF
C76996 NAND2X1_LOC_198/B VDD 2.84fF
C76997 NAND2X1_LOC_552/a_36_24# INVX1_LOC_28/A 0.01fF
C76998 NOR2X1_LOC_596/A INVX1_LOC_139/A 1.83fF
C76999 INVX1_LOC_33/A NOR2X1_LOC_708/A 0.63fF
C77000 INVX1_LOC_220/Y NOR2X1_LOC_703/A 0.00fF
C77001 NAND2X1_LOC_733/Y INVX1_LOC_118/A 0.07fF
C77002 NAND2X1_LOC_337/B INVX1_LOC_131/Y 0.61fF
C77003 NAND2X1_LOC_859/Y INVX1_LOC_140/A 0.01fF
C77004 INVX1_LOC_48/Y NOR2X1_LOC_813/a_36_216# 0.01fF
C77005 NOR2X1_LOC_660/Y NOR2X1_LOC_847/B 0.10fF
C77006 NOR2X1_LOC_295/Y INVX1_LOC_93/Y 0.01fF
C77007 NAND2X1_LOC_783/A INVX1_LOC_28/A 0.10fF
C77008 NOR2X1_LOC_210/A INVX1_LOC_75/A 0.46fF
C77009 INVX1_LOC_227/A NOR2X1_LOC_329/B 0.05fF
C77010 NOR2X1_LOC_773/Y INVX1_LOC_6/A 0.10fF
C77011 INVX1_LOC_58/A INVX1_LOC_47/Y 0.03fF
C77012 NOR2X1_LOC_619/A NOR2X1_LOC_721/Y 0.06fF
C77013 INVX1_LOC_184/Y INVX1_LOC_37/A 0.01fF
C77014 NOR2X1_LOC_91/A INVX1_LOC_78/A 0.14fF
C77015 INVX1_LOC_1/A INVX1_LOC_294/A 0.03fF
C77016 INVX1_LOC_28/A NOR2X1_LOC_130/A 0.13fF
C77017 INVX1_LOC_17/A NAND2X1_LOC_574/A 0.02fF
C77018 NOR2X1_LOC_516/B NOR2X1_LOC_391/B 0.04fF
C77019 NOR2X1_LOC_678/A NOR2X1_LOC_270/a_36_216# 0.00fF
C77020 INVX1_LOC_211/Y NOR2X1_LOC_88/Y 0.08fF
C77021 NOR2X1_LOC_763/Y D_INPUT_4 0.00fF
C77022 INVX1_LOC_39/A INVX1_LOC_12/A 0.03fF
C77023 INVX1_LOC_217/A INVX1_LOC_118/A 0.10fF
C77024 INVX1_LOC_310/Y VDD 0.21fF
C77025 INVX1_LOC_250/A INVX1_LOC_185/A 0.00fF
C77026 INVX1_LOC_153/Y INVX1_LOC_37/A 0.04fF
C77027 INVX1_LOC_78/A INVX1_LOC_23/A 0.20fF
C77028 NAND2X1_LOC_562/Y INVX1_LOC_178/Y 0.13fF
C77029 NAND2X1_LOC_866/B INVX1_LOC_140/A 0.01fF
C77030 NOR2X1_LOC_502/Y NOR2X1_LOC_814/A 0.15fF
C77031 NAND2X1_LOC_555/Y NAND2X1_LOC_574/A 0.07fF
C77032 NOR2X1_LOC_471/Y INVX1_LOC_136/Y 0.34fF
C77033 NOR2X1_LOC_454/Y NOR2X1_LOC_584/Y 0.06fF
C77034 NAND2X1_LOC_159/a_36_24# INVX1_LOC_123/A 0.01fF
C77035 INVX1_LOC_121/Y INVX1_LOC_37/A 0.01fF
C77036 INVX1_LOC_198/Y INVX1_LOC_274/A 0.00fF
C77037 NAND2X1_LOC_738/B NOR2X1_LOC_829/A 0.06fF
C77038 NOR2X1_LOC_67/A NOR2X1_LOC_670/a_36_216# 0.01fF
C77039 INVX1_LOC_196/A INVX1_LOC_143/Y 0.03fF
C77040 NAND2X1_LOC_579/A NOR2X1_LOC_89/A 0.10fF
C77041 INVX1_LOC_140/A NAND2X1_LOC_807/Y 0.10fF
C77042 NOR2X1_LOC_717/B NOR2X1_LOC_728/B 0.37fF
C77043 NOR2X1_LOC_65/B NOR2X1_LOC_262/a_36_216# 0.02fF
C77044 INVX1_LOC_143/A NOR2X1_LOC_35/Y 0.10fF
C77045 NAND2X1_LOC_850/A INVX1_LOC_102/Y 0.01fF
C77046 INVX1_LOC_34/A NOR2X1_LOC_561/A 0.00fF
C77047 NOR2X1_LOC_187/Y NOR2X1_LOC_89/A 0.01fF
C77048 NOR2X1_LOC_216/Y INVX1_LOC_28/A 0.12fF
C77049 NOR2X1_LOC_287/A NOR2X1_LOC_542/B 0.08fF
C77050 NOR2X1_LOC_667/A INVX1_LOC_126/A 0.07fF
C77051 INVX1_LOC_161/Y INVX1_LOC_19/A 0.07fF
C77052 NOR2X1_LOC_501/a_36_216# INVX1_LOC_91/A 0.01fF
C77053 NAND2X1_LOC_527/a_36_24# NOR2X1_LOC_814/A 0.01fF
C77054 NOR2X1_LOC_497/Y NAND2X1_LOC_849/A 0.02fF
C77055 INVX1_LOC_177/A INVX1_LOC_37/A 0.03fF
C77056 INVX1_LOC_89/A NAND2X1_LOC_328/a_36_24# 0.00fF
C77057 INVX1_LOC_90/A INPUT_0 0.31fF
C77058 INVX1_LOC_34/A NAND2X1_LOC_849/B 0.01fF
C77059 NAND2X1_LOC_725/A NOR2X1_LOC_409/B 0.03fF
C77060 INVX1_LOC_267/Y VDD -0.00fF
C77061 NOR2X1_LOC_65/B INVX1_LOC_23/A 0.04fF
C77062 INVX1_LOC_18/A INVX1_LOC_113/A 0.01fF
C77063 NAND2X1_LOC_842/B NOR2X1_LOC_74/A 0.08fF
C77064 NOR2X1_LOC_590/A NOR2X1_LOC_691/B 0.03fF
C77065 INVX1_LOC_34/A INVX1_LOC_38/A 0.13fF
C77066 INVX1_LOC_224/Y INVX1_LOC_57/A 0.11fF
C77067 NAND2X1_LOC_787/B INVX1_LOC_118/A 0.19fF
C77068 NOR2X1_LOC_389/B INPUT_0 0.07fF
C77069 NOR2X1_LOC_78/B NOR2X1_LOC_266/B 0.03fF
C77070 NOR2X1_LOC_811/B VDD 0.02fF
C77071 INVX1_LOC_150/Y INVX1_LOC_29/A 0.03fF
C77072 NOR2X1_LOC_523/a_36_216# INVX1_LOC_280/A 0.00fF
C77073 NOR2X1_LOC_431/a_36_216# NOR2X1_LOC_592/B 0.00fF
C77074 INVX1_LOC_135/A INVX1_LOC_315/Y 0.02fF
C77075 NOR2X1_LOC_717/B INVX1_LOC_91/A 0.05fF
C77076 NAND2X1_LOC_860/A NOR2X1_LOC_383/B 0.07fF
C77077 NOR2X1_LOC_303/Y INVX1_LOC_179/A 0.01fF
C77078 INVX1_LOC_34/A NOR2X1_LOC_96/Y 0.20fF
C77079 NAND2X1_LOC_842/B NOR2X1_LOC_9/Y 0.06fF
C77080 NOR2X1_LOC_736/Y INVX1_LOC_311/A 0.06fF
C77081 NOR2X1_LOC_667/A NOR2X1_LOC_111/A 2.98fF
C77082 INVX1_LOC_49/A INVX1_LOC_92/A 0.23fF
C77083 D_INPUT_0 NOR2X1_LOC_311/Y 0.01fF
C77084 INVX1_LOC_248/A NOR2X1_LOC_111/A 0.09fF
C77085 NOR2X1_LOC_219/Y VDD 0.28fF
C77086 NAND2X1_LOC_740/Y NAND2X1_LOC_175/Y 0.16fF
C77087 NOR2X1_LOC_383/B NOR2X1_LOC_634/Y 0.12fF
C77088 NOR2X1_LOC_500/Y INVX1_LOC_14/Y 0.10fF
C77089 INVX1_LOC_312/A INVX1_LOC_19/A 0.02fF
C77090 INVX1_LOC_57/A NAND2X1_LOC_793/B 0.07fF
C77091 NAND2X1_LOC_214/B INVX1_LOC_16/Y 0.38fF
C77092 NAND2X1_LOC_162/A INVX1_LOC_37/A 0.01fF
C77093 INVX1_LOC_34/A NOR2X1_LOC_51/A 0.03fF
C77094 NOR2X1_LOC_822/Y NOR2X1_LOC_536/A 0.01fF
C77095 NOR2X1_LOC_632/Y INVX1_LOC_76/A 0.05fF
C77096 INVX1_LOC_53/Y VDD 1.31fF
C77097 NAND2X1_LOC_348/A INPUT_0 0.07fF
C77098 NOR2X1_LOC_619/A VDD 0.21fF
C77099 INVX1_LOC_155/Y NAND2X1_LOC_93/B 0.15fF
C77100 NOR2X1_LOC_473/B NOR2X1_LOC_78/A 0.07fF
C77101 INVX1_LOC_8/A NOR2X1_LOC_99/Y 0.07fF
C77102 NAND2X1_LOC_231/Y INVX1_LOC_38/A 0.03fF
C77103 NOR2X1_LOC_607/A NAND2X1_LOC_475/Y 0.02fF
C77104 INVX1_LOC_31/A NOR2X1_LOC_847/A 0.03fF
C77105 INVX1_LOC_193/Y INVX1_LOC_75/A 0.03fF
C77106 INVX1_LOC_133/Y INVX1_LOC_9/A 0.01fF
C77107 NOR2X1_LOC_92/Y INVX1_LOC_94/Y 0.03fF
C77108 NOR2X1_LOC_151/Y NOR2X1_LOC_728/B -0.01fF
C77109 NOR2X1_LOC_254/Y INVX1_LOC_179/A 2.01fF
C77110 NAND2X1_LOC_660/Y INVX1_LOC_46/A 0.50fF
C77111 NOR2X1_LOC_665/A VDD 0.04fF
C77112 INVX1_LOC_5/A INVX1_LOC_270/A 0.01fF
C77113 INVX1_LOC_89/A NOR2X1_LOC_124/A 0.02fF
C77114 INVX1_LOC_31/A INVX1_LOC_42/A 0.17fF
C77115 NOR2X1_LOC_68/A INVX1_LOC_262/Y 0.02fF
C77116 INVX1_LOC_50/A NOR2X1_LOC_674/a_36_216# 0.02fF
C77117 NOR2X1_LOC_67/A INVX1_LOC_9/A 0.22fF
C77118 INVX1_LOC_136/A NAND2X1_LOC_74/B 0.92fF
C77119 NOR2X1_LOC_781/B VDD 0.03fF
C77120 NAND2X1_LOC_303/Y NOR2X1_LOC_36/A 0.07fF
C77121 NAND2X1_LOC_214/B NAND2X1_LOC_205/A 0.10fF
C77122 NOR2X1_LOC_82/A NOR2X1_LOC_38/B 6.77fF
C77123 INVX1_LOC_145/Y VDD 0.30fF
C77124 INVX1_LOC_71/A NOR2X1_LOC_662/A 0.02fF
C77125 INVX1_LOC_5/A NOR2X1_LOC_416/A 0.07fF
C77126 NOR2X1_LOC_15/Y NOR2X1_LOC_471/a_36_216# 0.00fF
C77127 NOR2X1_LOC_785/Y INVX1_LOC_37/A 0.03fF
C77128 INVX1_LOC_166/A NAND2X1_LOC_398/a_36_24# 0.01fF
C77129 INVX1_LOC_103/A INVX1_LOC_271/Y 0.31fF
C77130 NOR2X1_LOC_467/a_36_216# INVX1_LOC_117/A 0.00fF
C77131 NOR2X1_LOC_151/Y INVX1_LOC_91/A 0.07fF
C77132 NOR2X1_LOC_516/B INVX1_LOC_280/A 0.10fF
C77133 D_INPUT_0 INVX1_LOC_46/A 0.17fF
C77134 NOR2X1_LOC_424/a_36_216# INVX1_LOC_117/A 0.01fF
C77135 INVX1_LOC_2/A INVX1_LOC_92/A 3.28fF
C77136 NOR2X1_LOC_321/Y NOR2X1_LOC_135/a_36_216# 0.00fF
C77137 D_INPUT_0 NOR2X1_LOC_98/A 0.02fF
C77138 INVX1_LOC_27/A NAND2X1_LOC_205/A 0.00fF
C77139 NAND2X1_LOC_367/B VDD 0.01fF
C77140 NOR2X1_LOC_794/B NOR2X1_LOC_334/Y 0.07fF
C77141 INVX1_LOC_24/A INVX1_LOC_109/A 0.01fF
C77142 NAND2X1_LOC_728/a_36_24# NAND2X1_LOC_800/A 0.00fF
C77143 INVX1_LOC_83/A NOR2X1_LOC_859/Y 0.03fF
C77144 NOR2X1_LOC_226/A INVX1_LOC_92/A 0.26fF
C77145 INVX1_LOC_69/Y NOR2X1_LOC_501/B 0.02fF
C77146 NOR2X1_LOC_507/B VDD -0.00fF
C77147 NOR2X1_LOC_78/B INVX1_LOC_46/Y 0.20fF
C77148 NOR2X1_LOC_289/Y NAND2X1_LOC_468/B 0.01fF
C77149 D_INPUT_0 NAND2X1_LOC_417/a_36_24# 0.01fF
C77150 INVX1_LOC_290/A NAND2X1_LOC_637/Y 0.11fF
C77151 INVX1_LOC_92/Y NOR2X1_LOC_78/A 0.03fF
C77152 NOR2X1_LOC_135/Y INVX1_LOC_76/A 0.02fF
C77153 INVX1_LOC_83/A NAND2X1_LOC_848/A 0.10fF
C77154 INVX1_LOC_31/A INVX1_LOC_78/A 0.12fF
C77155 NOR2X1_LOC_214/B INVX1_LOC_281/A 0.07fF
C77156 NOR2X1_LOC_91/A NOR2X1_LOC_503/Y 0.03fF
C77157 NAND2X1_LOC_738/B NAND2X1_LOC_537/Y 0.01fF
C77158 NOR2X1_LOC_815/Y INVX1_LOC_12/A 0.01fF
C77159 NOR2X1_LOC_717/Y NAND2X1_LOC_454/Y 0.02fF
C77160 INVX1_LOC_89/A NOR2X1_LOC_684/Y 0.09fF
C77161 INVX1_LOC_280/Y NOR2X1_LOC_485/a_36_216# 0.01fF
C77162 NOR2X1_LOC_175/A INVX1_LOC_63/A 0.03fF
C77163 INVX1_LOC_39/Y INVX1_LOC_26/A 0.16fF
C77164 INVX1_LOC_33/A INVX1_LOC_99/A 0.01fF
C77165 INVX1_LOC_30/A NAND2X1_LOC_443/a_36_24# 0.00fF
C77166 NOR2X1_LOC_103/Y INVX1_LOC_57/A 0.16fF
C77167 NOR2X1_LOC_92/a_36_216# INPUT_0 0.00fF
C77168 NOR2X1_LOC_84/Y NAND2X1_LOC_773/B 0.07fF
C77169 INVX1_LOC_223/Y INVX1_LOC_50/Y 0.03fF
C77170 INVX1_LOC_255/Y NOR2X1_LOC_216/B 0.03fF
C77171 INVX1_LOC_28/A NAND2X1_LOC_811/B 0.01fF
C77172 NAND2X1_LOC_573/A NOR2X1_LOC_743/Y 0.14fF
C77173 NOR2X1_LOC_381/Y NOR2X1_LOC_392/Y 0.11fF
C77174 NAND2X1_LOC_863/B NAND2X1_LOC_770/Y 0.23fF
C77175 INVX1_LOC_93/Y INVX1_LOC_100/Y 0.01fF
C77176 INVX1_LOC_21/A NOR2X1_LOC_272/Y 0.05fF
C77177 NAND2X1_LOC_30/Y INVX1_LOC_53/A 0.02fF
C77178 INVX1_LOC_11/A INVX1_LOC_308/A 0.01fF
C77179 INVX1_LOC_8/A NOR2X1_LOC_76/B 0.04fF
C77180 NOR2X1_LOC_113/B VDD -0.00fF
C77181 NAND2X1_LOC_787/A NAND2X1_LOC_793/Y 0.01fF
C77182 NOR2X1_LOC_181/A INVX1_LOC_91/A 0.01fF
C77183 NOR2X1_LOC_195/A INVX1_LOC_108/Y 0.03fF
C77184 NOR2X1_LOC_15/Y NOR2X1_LOC_304/Y 0.06fF
C77185 NAND2X1_LOC_347/B NOR2X1_LOC_652/Y 0.01fF
C77186 NOR2X1_LOC_750/Y INVX1_LOC_230/Y 0.01fF
C77187 INVX1_LOC_17/A NAND2X1_LOC_35/Y 0.01fF
C77188 INVX1_LOC_13/A INVX1_LOC_84/A 0.11fF
C77189 INVX1_LOC_45/A NOR2X1_LOC_851/a_36_216# 0.00fF
C77190 INVX1_LOC_266/A INVX1_LOC_223/Y 0.01fF
C77191 NOR2X1_LOC_71/Y NOR2X1_LOC_216/B 0.10fF
C77192 NOR2X1_LOC_112/Y NOR2X1_LOC_332/Y 0.03fF
C77193 NAND2X1_LOC_33/a_36_24# INVX1_LOC_64/A 0.00fF
C77194 INVX1_LOC_45/A INVX1_LOC_57/A 0.20fF
C77195 NOR2X1_LOC_387/a_36_216# NOR2X1_LOC_409/B 0.00fF
C77196 NAND2X1_LOC_337/B NOR2X1_LOC_109/Y 0.10fF
C77197 NOR2X1_LOC_290/Y INVX1_LOC_42/A 0.06fF
C77198 INVX1_LOC_35/A NOR2X1_LOC_590/A 0.87fF
C77199 INVX1_LOC_151/Y INVX1_LOC_272/A 0.01fF
C77200 INPUT_0 INVX1_LOC_38/A 0.11fF
C77201 NAND2X1_LOC_98/a_36_24# NOR2X1_LOC_92/Y 0.01fF
C77202 INVX1_LOC_35/A INVX1_LOC_22/Y 0.03fF
C77203 INVX1_LOC_64/A INVX1_LOC_130/A 0.04fF
C77204 NOR2X1_LOC_470/B NAND2X1_LOC_149/Y 0.02fF
C77205 NOR2X1_LOC_655/B NOR2X1_LOC_159/a_36_216# 0.12fF
C77206 INVX1_LOC_195/Y NOR2X1_LOC_476/B 0.26fF
C77207 NOR2X1_LOC_261/a_36_216# NOR2X1_LOC_68/A 0.00fF
C77208 INVX1_LOC_244/Y NOR2X1_LOC_654/A 0.07fF
C77209 NAND2X1_LOC_36/a_36_24# INVX1_LOC_23/A 0.02fF
C77210 INVX1_LOC_208/Y NOR2X1_LOC_89/A 0.26fF
C77211 NOR2X1_LOC_91/A NOR2X1_LOC_152/Y 0.09fF
C77212 NAND2X1_LOC_533/a_36_24# INVX1_LOC_30/A 0.06fF
C77213 INVX1_LOC_50/A INVX1_LOC_41/Y 0.00fF
C77214 INVX1_LOC_65/A INVX1_LOC_37/A 0.01fF
C77215 NOR2X1_LOC_71/Y NAND2X1_LOC_477/Y 0.04fF
C77216 INVX1_LOC_299/A INVX1_LOC_24/Y 0.03fF
C77217 NAND2X1_LOC_9/Y NOR2X1_LOC_791/A 0.01fF
C77218 NAND2X1_LOC_326/A NAND2X1_LOC_538/Y 0.04fF
C77219 NOR2X1_LOC_667/Y NOR2X1_LOC_406/A 0.16fF
C77220 NOR2X1_LOC_322/a_36_216# INVX1_LOC_91/A 0.00fF
C77221 NAND2X1_LOC_735/B INVX1_LOC_12/A 0.15fF
C77222 INVX1_LOC_145/Y INVX1_LOC_133/A 0.02fF
C77223 INVX1_LOC_139/A NAND2X1_LOC_469/B 0.00fF
C77224 INVX1_LOC_226/Y NOR2X1_LOC_38/a_36_216# 0.01fF
C77225 INVX1_LOC_71/A INVX1_LOC_57/A 0.03fF
C77226 NOR2X1_LOC_264/Y NOR2X1_LOC_621/B 0.01fF
C77227 NAND2X1_LOC_477/A INVX1_LOC_94/Y 0.06fF
C77228 NOR2X1_LOC_360/Y NOR2X1_LOC_717/A 0.10fF
C77229 NOR2X1_LOC_75/a_36_216# INVX1_LOC_78/A 0.01fF
C77230 NAND2X1_LOC_326/A NOR2X1_LOC_250/A 0.03fF
C77231 INVX1_LOC_11/A NAND2X1_LOC_579/A 0.01fF
C77232 INVX1_LOC_119/A INVX1_LOC_273/A 0.01fF
C77233 INVX1_LOC_55/Y INVX1_LOC_84/A 0.03fF
C77234 INVX1_LOC_2/Y INVX1_LOC_20/A 0.03fF
C77235 NOR2X1_LOC_82/A NOR2X1_LOC_468/Y 0.15fF
C77236 INVX1_LOC_36/A INVX1_LOC_5/A 0.09fF
C77237 NOR2X1_LOC_479/B INVX1_LOC_3/Y 0.07fF
C77238 INVX1_LOC_41/A INVX1_LOC_181/A 0.03fF
C77239 NOR2X1_LOC_152/Y INVX1_LOC_23/A 0.01fF
C77240 INVX1_LOC_31/A NOR2X1_LOC_655/a_36_216# 0.00fF
C77241 INVX1_LOC_2/Y NOR2X1_LOC_360/A 0.02fF
C77242 VDD NOR2X1_LOC_585/Y 0.12fF
C77243 NAND2X1_LOC_859/Y INVX1_LOC_42/A 0.04fF
C77244 INVX1_LOC_254/Y NOR2X1_LOC_622/A 0.12fF
C77245 NOR2X1_LOC_709/B INVX1_LOC_91/A 0.01fF
C77246 NAND2X1_LOC_140/A INVX1_LOC_272/A 0.03fF
C77247 INVX1_LOC_135/A NAND2X1_LOC_207/B 0.02fF
C77248 NOR2X1_LOC_639/B NOR2X1_LOC_781/Y 0.01fF
C77249 NAND2X1_LOC_553/A NOR2X1_LOC_791/A 0.07fF
C77250 NOR2X1_LOC_266/B INVX1_LOC_46/A 0.05fF
C77251 INVX1_LOC_178/Y D_INPUT_3 0.07fF
C77252 NOR2X1_LOC_130/A INVX1_LOC_109/A 0.01fF
C77253 NAND2X1_LOC_687/A INVX1_LOC_20/A 0.01fF
C77254 NAND2X1_LOC_649/B INVX1_LOC_38/A 0.01fF
C77255 INVX1_LOC_72/A INVX1_LOC_306/Y 0.35fF
C77256 D_INPUT_0 NOR2X1_LOC_671/Y 0.03fF
C77257 INVX1_LOC_139/A NAND2X1_LOC_212/a_36_24# 0.00fF
C77258 INVX1_LOC_191/Y INVX1_LOC_78/A 0.03fF
C77259 NAND2X1_LOC_357/B NOR2X1_LOC_318/A 0.00fF
C77260 INVX1_LOC_37/Y INVX1_LOC_20/A 0.01fF
C77261 NOR2X1_LOC_726/a_36_216# INVX1_LOC_117/A 0.00fF
C77262 D_INPUT_6 INVX1_LOC_30/A 0.05fF
C77263 NOR2X1_LOC_303/Y NOR2X1_LOC_405/Y 0.09fF
C77264 INVX1_LOC_36/A INVX1_LOC_178/A 0.11fF
C77265 NOR2X1_LOC_646/A INVX1_LOC_4/A 0.07fF
C77266 NOR2X1_LOC_635/A NOR2X1_LOC_635/B 0.00fF
C77267 INVX1_LOC_49/A INVX1_LOC_53/A 0.26fF
C77268 INVX1_LOC_114/A NAND2X1_LOC_212/Y 0.03fF
C77269 INVX1_LOC_13/A INVX1_LOC_15/A 0.07fF
C77270 NAND2X1_LOC_477/A INVX1_LOC_181/A 0.10fF
C77271 INVX1_LOC_256/A NOR2X1_LOC_218/A 0.01fF
C77272 NOR2X1_LOC_321/Y INVX1_LOC_30/A 0.46fF
C77273 NOR2X1_LOC_74/A INVX1_LOC_119/Y 0.02fF
C77274 VDD INVX1_LOC_77/Y 0.75fF
C77275 INVX1_LOC_21/A NAND2X1_LOC_364/A 0.09fF
C77276 NOR2X1_LOC_78/A NOR2X1_LOC_259/A 0.01fF
C77277 NOR2X1_LOC_510/Y NAND2X1_LOC_198/B 0.10fF
C77278 INVX1_LOC_5/A NOR2X1_LOC_208/Y 0.06fF
C77279 NOR2X1_LOC_107/Y NAND2X1_LOC_114/B 0.13fF
C77280 INVX1_LOC_288/A INVX1_LOC_191/Y 0.01fF
C77281 NOR2X1_LOC_188/A INVX1_LOC_294/A 0.17fF
C77282 NAND2X1_LOC_555/Y NAND2X1_LOC_377/a_36_24# 0.01fF
C77283 INVX1_LOC_219/A INVX1_LOC_3/Y 0.03fF
C77284 NAND2X1_LOC_848/A INVX1_LOC_46/A 0.01fF
C77285 NAND2X1_LOC_866/B INVX1_LOC_42/A 1.44fF
C77286 NOR2X1_LOC_236/a_36_216# NOR2X1_LOC_38/B 0.00fF
C77287 NAND2X1_LOC_785/a_36_24# NOR2X1_LOC_753/Y 0.02fF
C77288 INVX1_LOC_201/A NOR2X1_LOC_673/A 0.13fF
C77289 NAND2X1_LOC_200/B NOR2X1_LOC_39/Y 0.00fF
C77290 NOR2X1_LOC_246/A INVX1_LOC_15/A 0.07fF
C77291 NAND2X1_LOC_859/Y INVX1_LOC_78/A 0.03fF
C77292 NOR2X1_LOC_6/B NOR2X1_LOC_392/Y 0.03fF
C77293 NAND2X1_LOC_807/Y INVX1_LOC_42/A 0.07fF
C77294 NOR2X1_LOC_174/B INVX1_LOC_15/A 0.04fF
C77295 NOR2X1_LOC_68/A INVX1_LOC_14/A 0.08fF
C77296 INVX1_LOC_30/A NAND2X1_LOC_793/Y 0.03fF
C77297 INVX1_LOC_48/Y INVX1_LOC_24/A 0.10fF
C77298 NOR2X1_LOC_242/A INVX1_LOC_49/A 0.03fF
C77299 INVX1_LOC_2/A INVX1_LOC_53/A 0.13fF
C77300 INVX1_LOC_22/A NOR2X1_LOC_638/Y 0.01fF
C77301 NAND2X1_LOC_537/Y NOR2X1_LOC_512/Y 0.02fF
C77302 INVX1_LOC_141/A INVX1_LOC_141/Y 0.16fF
C77303 INVX1_LOC_64/A NOR2X1_LOC_802/A 0.05fF
C77304 INVX1_LOC_36/A NOR2X1_LOC_816/A 0.06fF
C77305 INVX1_LOC_55/Y INVX1_LOC_15/A 0.03fF
C77306 NOR2X1_LOC_361/B NAND2X1_LOC_198/B 0.19fF
C77307 INVX1_LOC_290/A NOR2X1_LOC_639/Y 0.01fF
C77308 NOR2X1_LOC_359/Y NOR2X1_LOC_359/a_36_216# 0.00fF
C77309 NAND2X1_LOC_552/A NOR2X1_LOC_309/Y 0.34fF
C77310 NAND2X1_LOC_796/B NAND2X1_LOC_833/Y 0.02fF
C77311 NAND2X1_LOC_36/A NOR2X1_LOC_389/A 0.01fF
C77312 INVX1_LOC_54/Y NOR2X1_LOC_405/Y 0.01fF
C77313 NOR2X1_LOC_226/A INVX1_LOC_53/A 0.10fF
C77314 NOR2X1_LOC_35/Y NOR2X1_LOC_197/B 0.45fF
C77315 NOR2X1_LOC_437/Y NOR2X1_LOC_122/A 0.06fF
C77316 INVX1_LOC_141/A INVX1_LOC_312/Y 0.05fF
C77317 INVX1_LOC_17/A INVX1_LOC_94/A 0.19fF
C77318 INVX1_LOC_313/A INVX1_LOC_78/A 1.20fF
C77319 INVX1_LOC_46/A INVX1_LOC_46/Y 0.16fF
C77320 INVX1_LOC_58/A NOR2X1_LOC_328/Y 0.03fF
C77321 INVX1_LOC_14/Y INVX1_LOC_307/A 0.10fF
C77322 NAND2X1_LOC_605/a_36_24# INVX1_LOC_92/A 0.00fF
C77323 NAND2X1_LOC_866/B INVX1_LOC_78/A 0.02fF
C77324 INVX1_LOC_235/A NOR2X1_LOC_6/B 0.06fF
C77325 NOR2X1_LOC_598/B NOR2X1_LOC_210/B 0.42fF
C77326 INVX1_LOC_31/A NOR2X1_LOC_554/B 1.78fF
C77327 INVX1_LOC_62/A INVX1_LOC_26/Y 0.00fF
C77328 NOR2X1_LOC_89/A NOR2X1_LOC_501/B 0.02fF
C77329 INVX1_LOC_6/A INVX1_LOC_42/A 0.28fF
C77330 NOR2X1_LOC_773/Y NOR2X1_LOC_109/Y 0.07fF
C77331 NOR2X1_LOC_729/A INVX1_LOC_9/A 4.93fF
C77332 INVX1_LOC_24/A INVX1_LOC_246/A 0.00fF
C77333 NOR2X1_LOC_92/Y INVX1_LOC_162/A 0.01fF
C77334 INVX1_LOC_41/A INVX1_LOC_299/A 0.03fF
C77335 NAND2X1_LOC_338/B INVX1_LOC_306/Y 0.23fF
C77336 NAND2X1_LOC_807/Y INVX1_LOC_78/A 0.07fF
C77337 NOR2X1_LOC_666/A INVX1_LOC_88/Y 0.02fF
C77338 INVX1_LOC_20/A NOR2X1_LOC_485/Y 0.00fF
C77339 NOR2X1_LOC_78/A INVX1_LOC_106/A 0.01fF
C77340 NOR2X1_LOC_357/Y INVX1_LOC_84/A 0.09fF
C77341 NOR2X1_LOC_65/B INVX1_LOC_313/A 0.08fF
C77342 INVX1_LOC_286/A INVX1_LOC_170/Y 0.03fF
C77343 INVX1_LOC_1/A NOR2X1_LOC_718/B 0.71fF
C77344 NOR2X1_LOC_92/Y NOR2X1_LOC_315/Y 0.72fF
C77345 NOR2X1_LOC_20/Y INVX1_LOC_34/A 0.09fF
C77346 NAND2X1_LOC_579/A NOR2X1_LOC_52/B 2.78fF
C77347 NOR2X1_LOC_123/B INVX1_LOC_57/A 0.07fF
C77348 INVX1_LOC_21/A NAND2X1_LOC_11/Y 0.44fF
C77349 NAND2X1_LOC_579/A NAND2X1_LOC_838/Y 0.02fF
C77350 NOR2X1_LOC_795/Y NOR2X1_LOC_793/A 0.03fF
C77351 INVX1_LOC_85/Y NOR2X1_LOC_383/B 0.87fF
C77352 NAND2X1_LOC_36/A NOR2X1_LOC_596/A 0.01fF
C77353 NOR2X1_LOC_607/A INVX1_LOC_30/A 0.14fF
C77354 INVX1_LOC_31/A NOR2X1_LOC_152/Y 0.17fF
C77355 INVX1_LOC_171/A INVX1_LOC_29/Y 0.03fF
C77356 INVX1_LOC_118/A INVX1_LOC_92/A 0.16fF
C77357 NOR2X1_LOC_188/A NOR2X1_LOC_334/Y 0.00fF
C77358 NOR2X1_LOC_554/B NAND2X1_LOC_106/a_36_24# 0.02fF
C77359 NAND2X1_LOC_9/Y D_INPUT_0 0.18fF
C77360 INPUT_0 NAND2X1_LOC_223/A 0.63fF
C77361 INVX1_LOC_204/Y GATE_479 0.33fF
C77362 INVX1_LOC_35/A NOR2X1_LOC_763/Y 0.49fF
C77363 NAND2X1_LOC_53/Y NOR2X1_LOC_194/Y 0.01fF
C77364 INVX1_LOC_233/A D_INPUT_0 0.07fF
C77365 INVX1_LOC_64/A NAND2X1_LOC_756/a_36_24# 0.00fF
C77366 INPUT_0 INVX1_LOC_18/Y 0.03fF
C77367 INVX1_LOC_202/Y NAND2X1_LOC_476/Y 0.32fF
C77368 NOR2X1_LOC_569/a_36_216# NOR2X1_LOC_383/B 0.00fF
C77369 INVX1_LOC_299/A NOR2X1_LOC_405/a_36_216# 0.00fF
C77370 NOR2X1_LOC_598/B INVX1_LOC_20/Y 0.02fF
C77371 INVX1_LOC_6/A INVX1_LOC_78/A 2.53fF
C77372 NOR2X1_LOC_261/Y INVX1_LOC_55/Y 0.08fF
C77373 INVX1_LOC_21/A NOR2X1_LOC_86/A 0.07fF
C77374 INVX1_LOC_100/A NOR2X1_LOC_278/Y 0.68fF
C77375 INVX1_LOC_278/A NAND2X1_LOC_551/A 0.02fF
C77376 INVX1_LOC_64/A NOR2X1_LOC_532/Y 0.03fF
C77377 NOR2X1_LOC_614/Y NOR2X1_LOC_793/A 0.02fF
C77378 NOR2X1_LOC_795/Y NOR2X1_LOC_160/B 0.01fF
C77379 NAND2X1_LOC_565/B INVX1_LOC_48/Y 0.02fF
C77380 INVX1_LOC_14/Y INVX1_LOC_12/A 0.44fF
C77381 INVX1_LOC_256/A NOR2X1_LOC_131/A 0.03fF
C77382 NOR2X1_LOC_269/Y INVX1_LOC_128/Y 0.04fF
C77383 D_INPUT_2 NOR2X1_LOC_8/a_36_216# 0.00fF
C77384 INVX1_LOC_251/Y NOR2X1_LOC_160/B 0.00fF
C77385 NOR2X1_LOC_798/A D_INPUT_0 0.03fF
C77386 INVX1_LOC_24/A NOR2X1_LOC_350/A 0.03fF
C77387 NOR2X1_LOC_361/B INVX1_LOC_53/Y 0.03fF
C77388 INVX1_LOC_5/A NAND2X1_LOC_482/a_36_24# 0.00fF
C77389 NOR2X1_LOC_65/B INVX1_LOC_6/A 0.08fF
C77390 INVX1_LOC_294/Y INVX1_LOC_72/A 0.02fF
C77391 NOR2X1_LOC_754/A INVX1_LOC_46/A 0.04fF
C77392 INVX1_LOC_99/Y NOR2X1_LOC_644/A 0.01fF
C77393 NOR2X1_LOC_124/a_36_216# NOR2X1_LOC_38/B 0.00fF
C77394 NOR2X1_LOC_45/B NOR2X1_LOC_89/Y 0.01fF
C77395 INVX1_LOC_59/Y NOR2X1_LOC_38/B 1.59fF
C77396 NAND2X1_LOC_11/Y NOR2X1_LOC_428/Y 0.02fF
C77397 INVX1_LOC_112/A NOR2X1_LOC_38/B 0.01fF
C77398 INVX1_LOC_280/A NAND2X1_LOC_81/a_36_24# -0.01fF
C77399 INVX1_LOC_313/Y NOR2X1_LOC_644/a_36_216# 0.01fF
C77400 NAND2X1_LOC_848/A NOR2X1_LOC_671/Y 0.00fF
C77401 INVX1_LOC_280/A NAND2X1_LOC_207/B 0.02fF
C77402 NOR2X1_LOC_717/B NAND2X1_LOC_512/a_36_24# 0.00fF
C77403 INVX1_LOC_118/Y INVX1_LOC_272/A 0.01fF
C77404 NOR2X1_LOC_220/B NOR2X1_LOC_389/B 0.01fF
C77405 NAND2X1_LOC_733/B NAND2X1_LOC_733/Y 0.00fF
C77406 NAND2X1_LOC_303/Y INVX1_LOC_10/A 0.07fF
C77407 NOR2X1_LOC_448/Y INVX1_LOC_83/A 0.03fF
C77408 INVX1_LOC_48/Y NOR2X1_LOC_130/A 0.03fF
C77409 INVX1_LOC_123/A NOR2X1_LOC_646/B 0.02fF
C77410 INVX1_LOC_2/Y INVX1_LOC_4/A 0.03fF
C77411 INVX1_LOC_103/A INVX1_LOC_279/A 0.02fF
C77412 NOR2X1_LOC_240/Y NAND2X1_LOC_348/A 0.05fF
C77413 INVX1_LOC_174/A NOR2X1_LOC_160/Y 0.01fF
C77414 NOR2X1_LOC_88/Y NAND2X1_LOC_489/Y 0.03fF
C77415 NOR2X1_LOC_15/Y INVX1_LOC_89/A 0.16fF
C77416 INVX1_LOC_31/A NAND2X1_LOC_859/B 0.02fF
C77417 INVX1_LOC_36/A NOR2X1_LOC_773/Y 0.37fF
C77418 NOR2X1_LOC_717/B NOR2X1_LOC_739/Y 0.00fF
C77419 INVX1_LOC_124/A INVX1_LOC_181/Y 0.02fF
C77420 INVX1_LOC_284/Y INVX1_LOC_22/A 0.10fF
C77421 INVX1_LOC_5/A NOR2X1_LOC_208/A 0.03fF
C77422 INVX1_LOC_75/A INVX1_LOC_50/Y 0.03fF
C77423 NAND2X1_LOC_276/Y NOR2X1_LOC_716/B 0.06fF
C77424 INVX1_LOC_286/Y INVX1_LOC_16/A 0.10fF
C77425 INVX1_LOC_24/A NOR2X1_LOC_84/Y 0.06fF
C77426 NAND2X1_LOC_63/Y INVX1_LOC_92/A 0.31fF
C77427 NAND2X1_LOC_30/Y INVX1_LOC_83/A 0.07fF
C77428 NOR2X1_LOC_590/A NOR2X1_LOC_188/Y 0.05fF
C77429 INVX1_LOC_34/A INVX1_LOC_33/A 13.26fF
C77430 NAND2X1_LOC_11/Y NOR2X1_LOC_582/Y 0.78fF
C77431 INVX1_LOC_91/A NOR2X1_LOC_591/A 0.06fF
C77432 NOR2X1_LOC_267/A NOR2X1_LOC_773/Y 0.12fF
C77433 INVX1_LOC_24/A NOR2X1_LOC_482/Y 0.02fF
C77434 INVX1_LOC_76/A NAND2X1_LOC_61/Y 0.02fF
C77435 NOR2X1_LOC_841/A INVX1_LOC_19/A 0.16fF
C77436 INVX1_LOC_84/A NAND2X1_LOC_489/Y 0.03fF
C77437 INVX1_LOC_35/A NOR2X1_LOC_713/a_36_216# 0.00fF
C77438 D_INPUT_3 NOR2X1_LOC_29/a_36_216# 0.00fF
C77439 NOR2X1_LOC_781/Y NAND2X1_LOC_654/a_36_24# 0.00fF
C77440 NAND2X1_LOC_733/Y INPUT_5 0.12fF
C77441 INVX1_LOC_246/A NOR2X1_LOC_130/A 0.01fF
C77442 NOR2X1_LOC_812/A NOR2X1_LOC_729/A 0.07fF
C77443 NOR2X1_LOC_222/Y NOR2X1_LOC_215/Y 0.01fF
C77444 INVX1_LOC_136/A NAND2X1_LOC_849/a_36_24# 0.01fF
C77445 NOR2X1_LOC_655/B INVX1_LOC_314/Y 0.10fF
C77446 INVX1_LOC_41/A NOR2X1_LOC_315/Y 0.03fF
C77447 NAND2X1_LOC_637/Y NOR2X1_LOC_467/A 0.01fF
C77448 INVX1_LOC_266/A INVX1_LOC_75/A 0.01fF
C77449 INVX1_LOC_90/A INVX1_LOC_225/Y 1.97fF
C77450 INVX1_LOC_315/A NAND2X1_LOC_847/a_36_24# 0.01fF
C77451 INVX1_LOC_227/Y NOR2X1_LOC_570/Y 0.05fF
C77452 INVX1_LOC_49/A NOR2X1_LOC_634/B 0.03fF
C77453 NAND2X1_LOC_213/A NAND2X1_LOC_51/B 0.03fF
C77454 INVX1_LOC_11/A NOR2X1_LOC_756/Y 0.03fF
C77455 INVX1_LOC_88/A NOR2X1_LOC_289/Y 0.01fF
C77456 NAND2X1_LOC_724/A NOR2X1_LOC_322/Y 0.01fF
C77457 INVX1_LOC_31/A NAND2X1_LOC_861/Y 0.07fF
C77458 INVX1_LOC_49/A NOR2X1_LOC_547/B 0.04fF
C77459 NOR2X1_LOC_392/Y NOR2X1_LOC_124/A 0.00fF
C77460 INVX1_LOC_103/A INVX1_LOC_182/Y 0.00fF
C77461 NOR2X1_LOC_78/B INVX1_LOC_49/A 0.26fF
C77462 INVX1_LOC_310/A INVX1_LOC_41/A 0.07fF
C77463 NOR2X1_LOC_215/A INVX1_LOC_6/A 0.08fF
C77464 NAND2X1_LOC_731/Y INVX1_LOC_22/A 0.01fF
C77465 NAND2X1_LOC_231/Y INVX1_LOC_33/A 0.01fF
C77466 INVX1_LOC_27/A INVX1_LOC_286/A 0.10fF
C77467 INVX1_LOC_233/Y NOR2X1_LOC_396/Y -0.03fF
C77468 INVX1_LOC_257/A INVX1_LOC_92/A 0.02fF
C77469 INVX1_LOC_36/A NOR2X1_LOC_332/A 0.09fF
C77470 NOR2X1_LOC_815/Y INVX1_LOC_214/Y 0.63fF
C77471 INVX1_LOC_254/A INVX1_LOC_226/Y 0.01fF
C77472 NOR2X1_LOC_151/Y NOR2X1_LOC_739/Y 0.03fF
C77473 NOR2X1_LOC_315/Y NAND2X1_LOC_477/A 0.03fF
C77474 INVX1_LOC_135/A INVX1_LOC_195/A 0.01fF
C77475 INVX1_LOC_208/Y NOR2X1_LOC_433/A 0.03fF
C77476 NOR2X1_LOC_259/B INVX1_LOC_15/A 0.01fF
C77477 NOR2X1_LOC_100/A NOR2X1_LOC_844/A 0.48fF
C77478 NAND2X1_LOC_198/B NAND2X1_LOC_573/A 0.03fF
C77479 INVX1_LOC_17/A INVX1_LOC_144/A 0.10fF
C77480 INVX1_LOC_223/A NAND2X1_LOC_189/a_36_24# 0.00fF
C77481 INVX1_LOC_21/A NOR2X1_LOC_349/A 0.10fF
C77482 INVX1_LOC_277/Y INVX1_LOC_85/Y 0.01fF
C77483 INVX1_LOC_99/Y NOR2X1_LOC_540/B 0.08fF
C77484 INVX1_LOC_292/A INVX1_LOC_182/Y 0.06fF
C77485 INVX1_LOC_124/Y NAND2X1_LOC_842/B 0.34fF
C77486 INVX1_LOC_34/A INVX1_LOC_40/A 0.03fF
C77487 INVX1_LOC_286/Y INVX1_LOC_28/A 0.07fF
C77488 INVX1_LOC_21/A NOR2X1_LOC_405/A 0.39fF
C77489 INVX1_LOC_58/A INVX1_LOC_33/Y 0.16fF
C77490 INVX1_LOC_233/A NOR2X1_LOC_266/B 0.01fF
C77491 NAND2X1_LOC_726/Y INVX1_LOC_34/A 0.01fF
C77492 INVX1_LOC_180/A NOR2X1_LOC_561/Y 0.06fF
C77493 NOR2X1_LOC_437/a_36_216# NAND2X1_LOC_656/Y 0.01fF
C77494 NOR2X1_LOC_773/Y NOR2X1_LOC_309/Y 1.35fF
C77495 NOR2X1_LOC_106/Y INVX1_LOC_10/A 0.03fF
C77496 NOR2X1_LOC_11/Y INPUT_7 0.00fF
C77497 NAND2X1_LOC_360/B NOR2X1_LOC_709/A 0.33fF
C77498 NOR2X1_LOC_561/a_36_216# INVX1_LOC_22/A 0.00fF
C77499 INVX1_LOC_32/A INVX1_LOC_84/A 0.23fF
C77500 NOR2X1_LOC_590/A NOR2X1_LOC_534/a_36_216# 0.00fF
C77501 INVX1_LOC_2/A NOR2X1_LOC_78/B 0.14fF
C77502 INVX1_LOC_36/A INVX1_LOC_140/A 0.03fF
C77503 INVX1_LOC_255/Y NOR2X1_LOC_84/A 0.05fF
C77504 INVX1_LOC_64/A NAND2X1_LOC_687/A 0.01fF
C77505 NAND2X1_LOC_571/B NOR2X1_LOC_536/A 0.03fF
C77506 INVX1_LOC_208/Y NOR2X1_LOC_52/B 0.00fF
C77507 INVX1_LOC_15/A NAND2X1_LOC_489/Y 0.03fF
C77508 NOR2X1_LOC_88/Y NAND2X1_LOC_175/Y 0.07fF
C77509 INVX1_LOC_235/Y NAND2X1_LOC_659/B 0.34fF
C77510 INVX1_LOC_89/A NOR2X1_LOC_860/B 0.08fF
C77511 INVX1_LOC_83/A INVX1_LOC_49/A 0.48fF
C77512 INVX1_LOC_64/A NOR2X1_LOC_363/Y 1.00fF
C77513 NOR2X1_LOC_91/A INVX1_LOC_291/A 0.14fF
C77514 INVX1_LOC_177/Y NOR2X1_LOC_329/B 0.27fF
C77515 NOR2X1_LOC_65/B NOR2X1_LOC_79/A 0.01fF
C77516 NOR2X1_LOC_248/Y INVX1_LOC_75/A 0.03fF
C77517 NOR2X1_LOC_226/A NOR2X1_LOC_78/B 0.07fF
C77518 NOR2X1_LOC_637/B INVX1_LOC_135/A 0.03fF
C77519 INVX1_LOC_159/A INVX1_LOC_28/A 0.00fF
C77520 NOR2X1_LOC_785/Y INVX1_LOC_310/Y 0.04fF
C77521 NOR2X1_LOC_91/A NAND2X1_LOC_802/Y 0.07fF
C77522 INVX1_LOC_233/A NAND2X1_LOC_848/A 0.10fF
C77523 INVX1_LOC_271/A INVX1_LOC_54/A 0.58fF
C77524 NOR2X1_LOC_829/a_36_216# NAND2X1_LOC_811/Y 0.00fF
C77525 INVX1_LOC_50/A INVX1_LOC_185/A 0.03fF
C77526 NOR2X1_LOC_690/A INVX1_LOC_10/A 0.08fF
C77527 INVX1_LOC_21/A NOR2X1_LOC_857/A 0.94fF
C77528 INVX1_LOC_105/Y INVX1_LOC_54/A 0.00fF
C77529 INVX1_LOC_303/A INVX1_LOC_65/Y 0.01fF
C77530 NOR2X1_LOC_454/Y INVX1_LOC_115/A 0.10fF
C77531 NAND2X1_LOC_466/Y INVX1_LOC_10/A 0.09fF
C77532 NAND2X1_LOC_802/A INVX1_LOC_90/A 0.01fF
C77533 INVX1_LOC_104/A INVX1_LOC_220/Y 0.00fF
C77534 NOR2X1_LOC_644/A NOR2X1_LOC_303/Y 0.03fF
C77535 INVX1_LOC_53/A INVX1_LOC_118/A 0.07fF
C77536 NAND2X1_LOC_508/A NOR2X1_LOC_860/B 0.07fF
C77537 INVX1_LOC_248/Y INVX1_LOC_33/Y 0.01fF
C77538 NAND2X1_LOC_550/A NOR2X1_LOC_45/B 0.11fF
C77539 INVX1_LOC_72/A NOR2X1_LOC_74/A 0.10fF
C77540 INVX1_LOC_235/Y VDD 0.21fF
C77541 INVX1_LOC_84/A NAND2X1_LOC_175/Y 0.07fF
C77542 INVX1_LOC_52/Y INVX1_LOC_139/A -0.00fF
C77543 NOR2X1_LOC_781/Y INVX1_LOC_302/A 0.15fF
C77544 NAND2X1_LOC_149/Y VDD 3.25fF
C77545 NAND2X1_LOC_807/Y NOR2X1_LOC_152/Y 0.18fF
C77546 NOR2X1_LOC_15/Y NAND2X1_LOC_244/A 0.01fF
C77547 NOR2X1_LOC_67/A NOR2X1_LOC_719/A 0.00fF
C77548 INVX1_LOC_5/A NOR2X1_LOC_865/A 0.00fF
C77549 INVX1_LOC_68/A INVX1_LOC_9/A 0.02fF
C77550 NAND2X1_LOC_530/a_36_24# NOR2X1_LOC_548/A 0.00fF
C77551 INVX1_LOC_72/A NOR2X1_LOC_9/Y 0.10fF
C77552 NAND2X1_LOC_593/Y NAND2X1_LOC_652/Y 0.03fF
C77553 NOR2X1_LOC_216/B NAND2X1_LOC_205/A 0.05fF
C77554 INVX1_LOC_198/Y NOR2X1_LOC_74/A 0.09fF
C77555 NOR2X1_LOC_614/Y NOR2X1_LOC_516/B 0.33fF
C77556 NOR2X1_LOC_644/A NOR2X1_LOC_254/Y 0.01fF
C77557 NOR2X1_LOC_226/A NAND2X1_LOC_392/Y 0.03fF
C77558 NOR2X1_LOC_84/Y NOR2X1_LOC_130/A 0.09fF
C77559 NAND2X1_LOC_9/Y INVX1_LOC_46/Y 0.31fF
C77560 NOR2X1_LOC_67/A INVX1_LOC_7/A 0.09fF
C77561 INVX1_LOC_2/A INVX1_LOC_83/A 0.54fF
C77562 INVX1_LOC_83/A NOR2X1_LOC_818/Y 0.04fF
C77563 NOR2X1_LOC_160/B INVX1_LOC_199/Y 0.13fF
C77564 NOR2X1_LOC_533/Y NOR2X1_LOC_305/Y 0.02fF
C77565 NAND2X1_LOC_149/Y NOR2X1_LOC_684/a_36_216# 0.01fF
C77566 INVX1_LOC_89/A NAND2X1_LOC_141/A 0.02fF
C77567 INVX1_LOC_228/Y D_INPUT_3 0.02fF
C77568 NOR2X1_LOC_441/Y NOR2X1_LOC_657/B 0.36fF
C77569 NAND2X1_LOC_859/Y NAND2X1_LOC_859/B 0.39fF
C77570 NAND2X1_LOC_195/Y NOR2X1_LOC_45/B 0.03fF
C77571 NAND2X1_LOC_493/Y NOR2X1_LOC_536/A 1.73fF
C77572 NOR2X1_LOC_742/A INVX1_LOC_63/Y 0.10fF
C77573 NAND2X1_LOC_833/Y NAND2X1_LOC_840/Y 0.14fF
C77574 INVX1_LOC_32/A INVX1_LOC_15/A 0.06fF
C77575 NOR2X1_LOC_383/B NAND2X1_LOC_782/B 0.01fF
C77576 NOR2X1_LOC_329/B INVX1_LOC_104/A 0.22fF
C77577 INVX1_LOC_27/A INVX1_LOC_54/A 0.08fF
C77578 NOR2X1_LOC_521/Y NOR2X1_LOC_86/A 0.14fF
C77579 NOR2X1_LOC_309/Y INVX1_LOC_140/A 0.01fF
C77580 NOR2X1_LOC_152/Y INVX1_LOC_6/A 2.56fF
C77581 INVX1_LOC_33/A INPUT_0 0.39fF
C77582 NOR2X1_LOC_623/B INVX1_LOC_15/A 0.08fF
C77583 INVX1_LOC_132/A INVX1_LOC_92/Y 0.01fF
C77584 NOR2X1_LOC_134/Y INVX1_LOC_46/A 0.00fF
C77585 INVX1_LOC_89/A INVX1_LOC_226/A 0.01fF
C77586 NOR2X1_LOC_78/B INPUT_1 0.08fF
C77587 INVX1_LOC_113/Y INVX1_LOC_6/A 0.00fF
C77588 NOR2X1_LOC_6/B INVX1_LOC_75/A 0.13fF
C77589 NOR2X1_LOC_639/Y INVX1_LOC_261/Y 0.17fF
C77590 NAND2X1_LOC_651/B INVX1_LOC_262/A 0.02fF
C77591 INVX1_LOC_295/A NAND2X1_LOC_452/a_36_24# 0.01fF
C77592 INVX1_LOC_83/A NOR2X1_LOC_161/Y 0.03fF
C77593 NOR2X1_LOC_525/Y INVX1_LOC_22/A 0.00fF
C77594 INVX1_LOC_25/A NAND2X1_LOC_773/B 0.03fF
C77595 NOR2X1_LOC_598/B NOR2X1_LOC_257/Y 0.01fF
C77596 NAND2X1_LOC_572/a_36_24# INVX1_LOC_73/A 0.01fF
C77597 INVX1_LOC_278/A NAND2X1_LOC_489/Y 0.01fF
C77598 NAND2X1_LOC_323/B NOR2X1_LOC_356/A 0.01fF
C77599 NOR2X1_LOC_717/B NOR2X1_LOC_553/B 0.00fF
C77600 NOR2X1_LOC_355/A NOR2X1_LOC_589/A 0.06fF
C77601 NOR2X1_LOC_778/B INVX1_LOC_182/A 0.20fF
C77602 NOR2X1_LOC_160/B INVX1_LOC_281/A 0.07fF
C77603 NOR2X1_LOC_286/Y INVX1_LOC_9/A 3.76fF
C77604 NAND2X1_LOC_572/B NOR2X1_LOC_81/Y 0.03fF
C77605 NAND2X1_LOC_175/Y INVX1_LOC_15/A 0.07fF
C77606 INVX1_LOC_99/A NOR2X1_LOC_748/A 0.04fF
C77607 NAND2X1_LOC_859/Y NAND2X1_LOC_861/Y 0.01fF
C77608 NOR2X1_LOC_151/Y NOR2X1_LOC_352/Y 0.01fF
C77609 INVX1_LOC_225/Y INVX1_LOC_38/A 0.02fF
C77610 NAND2X1_LOC_552/A INVX1_LOC_63/A 0.02fF
C77611 INVX1_LOC_23/Y INVX1_LOC_3/Y 0.17fF
C77612 INVX1_LOC_13/A NOR2X1_LOC_5/a_36_216# 0.00fF
C77613 INVX1_LOC_5/A INVX1_LOC_63/A 3.03fF
C77614 NAND2X1_LOC_72/B INVX1_LOC_4/Y 0.01fF
C77615 NAND2X1_LOC_11/Y NAND2X1_LOC_51/B 0.26fF
C77616 NOR2X1_LOC_160/B NOR2X1_LOC_499/B 0.03fF
C77617 NOR2X1_LOC_793/A NOR2X1_LOC_862/B 0.34fF
C77618 NOR2X1_LOC_100/A INVX1_LOC_51/Y 0.01fF
C77619 NOR2X1_LOC_439/a_36_216# INVX1_LOC_182/A 0.02fF
C77620 NOR2X1_LOC_627/Y INVX1_LOC_311/A 0.01fF
C77621 NOR2X1_LOC_416/A INVX1_LOC_42/A 0.07fF
C77622 INVX1_LOC_205/Y NAND2X1_LOC_574/A 0.05fF
C77623 NOR2X1_LOC_537/Y NOR2X1_LOC_9/Y 0.03fF
C77624 INVX1_LOC_186/A NOR2X1_LOC_731/A 0.05fF
C77625 NOR2X1_LOC_744/Y VDD 0.23fF
C77626 INVX1_LOC_33/A NOR2X1_LOC_324/A 0.01fF
C77627 INVX1_LOC_17/A NOR2X1_LOC_155/A 0.07fF
C77628 INVX1_LOC_77/A INVX1_LOC_115/A 0.07fF
C77629 INVX1_LOC_40/A INPUT_0 0.02fF
C77630 NOR2X1_LOC_817/Y NOR2X1_LOC_216/B 0.00fF
C77631 NOR2X1_LOC_753/Y INVX1_LOC_76/A 0.01fF
C77632 NAND2X1_LOC_861/Y NAND2X1_LOC_866/B 0.07fF
C77633 NOR2X1_LOC_540/B NOR2X1_LOC_254/Y 0.04fF
C77634 NOR2X1_LOC_471/Y NOR2X1_LOC_155/A 0.01fF
C77635 NOR2X1_LOC_109/Y INVX1_LOC_42/A 0.07fF
C77636 NOR2X1_LOC_160/B NOR2X1_LOC_862/B 0.10fF
C77637 INVX1_LOC_49/A INVX1_LOC_46/A 0.18fF
C77638 INVX1_LOC_31/A INVX1_LOC_291/A 0.08fF
C77639 INVX1_LOC_29/Y INVX1_LOC_4/A 0.05fF
C77640 INVX1_LOC_161/Y NOR2X1_LOC_841/A 0.10fF
C77641 NAND2X1_LOC_325/Y INVX1_LOC_76/A 0.14fF
C77642 INVX1_LOC_2/A NOR2X1_LOC_311/Y 0.03fF
C77643 INVX1_LOC_124/A NAND2X1_LOC_107/a_36_24# 0.01fF
C77644 INVX1_LOC_164/Y INVX1_LOC_98/A 0.05fF
C77645 NAND2X1_LOC_454/Y NOR2X1_LOC_383/B 0.07fF
C77646 INVX1_LOC_45/A INVX1_LOC_274/A 0.07fF
C77647 NAND2X1_LOC_219/B NAND2X1_LOC_218/A 0.04fF
C77648 INVX1_LOC_278/A INVX1_LOC_32/A 0.03fF
C77649 INVX1_LOC_78/A INVX1_LOC_270/A 0.01fF
C77650 NOR2X1_LOC_569/Y NOR2X1_LOC_188/A 0.24fF
C77651 INVX1_LOC_21/A NOR2X1_LOC_841/a_36_216# 0.00fF
C77652 INVX1_LOC_63/Y INVX1_LOC_139/A 0.01fF
C77653 INVX1_LOC_1/A NAND2X1_LOC_773/B 0.10fF
C77654 INVX1_LOC_110/A NOR2X1_LOC_61/Y 0.10fF
C77655 INVX1_LOC_14/A NAND2X1_LOC_768/Y 0.06fF
C77656 INVX1_LOC_57/Y NOR2X1_LOC_487/Y 0.16fF
C77657 INVX1_LOC_202/A NOR2X1_LOC_366/a_36_216# 0.00fF
C77658 INVX1_LOC_285/Y NOR2X1_LOC_665/A 0.10fF
C77659 INPUT_7 VSS -0.29fF
C77660 INVX1_LOC_5/Y VSS 0.18fF
C77661 NAND2X1_LOC_780/Y VSS 0.22fF
C77662 NAND2X1_LOC_804/A VSS 0.37fF
C77663 NAND2X1_LOC_787/Y VSS 0.37fF
C77664 NOR2X1_LOC_801/B VSS 0.38fF
C77665 NAND2X1_LOC_773/B VSS 0.38fF
C77666 NAND2X1_LOC_768/Y VSS 0.18fF
C77667 NAND2X1_LOC_489/Y VSS 0.45fF
C77668 INVX1_LOC_92/A VSS -5.78fF
C77669 NOR2X1_LOC_271/Y VSS 0.72fF
C77670 NOR2X1_LOC_271/B VSS 0.12fF
C77671 NOR2X1_LOC_260/Y VSS 0.12fF
C77672 NOR2X1_LOC_226/Y VSS 0.06fF
C77673 NAND2X1_LOC_218/A VSS 0.34fF
C77674 NAND2X1_LOC_473/A VSS 0.33fF
C77675 NAND2X1_LOC_215/A VSS 0.61fF
C77676 INVX1_LOC_112/Y VSS 0.06fF
C77677 INVX1_LOC_42/A VSS 1.53fF
C77678 NOR2X1_LOC_485/Y VSS 0.34fF
C77679 NOR2X1_LOC_475/A VSS 0.17fF
C77680 NOR2X1_LOC_467/A VSS 0.63fF
C77681 NOR2X1_LOC_430/Y VSS 0.14fF
C77682 INVX1_LOC_198/A VSS -0.00fF
C77683 NOR2X1_LOC_460/Y VSS -0.10fF
C77684 INVX1_LOC_173/A VSS 0.35fF
C77685 NOR2X1_LOC_649/Y VSS 0.16fF
C77686 NOR2X1_LOC_748/A VSS 0.73fF
C77687 NOR2X1_LOC_624/B VSS 0.07fF
C77688 D_INPUT_5 VSS 0.10fF
C77689 NOR2X1_LOC_33/B VSS -0.05fF
C77690 NAND2X1_LOC_99/A VSS 1.04fF
C77691 NOR2X1_LOC_89/Y VSS 0.10fF
C77692 NOR2X1_LOC_640/B VSS 0.15fF
C77693 INVX1_LOC_69/A VSS 0.26fF
C77694 NOR2X1_LOC_633/A VSS 0.55fF
C77695 INVX1_LOC_275/Y VSS 0.33fF
C77696 INVX1_LOC_231/A VSS 0.44fF
C77697 INVX1_LOC_264/A VSS 0.13fF
C77698 INVX1_LOC_220/A VSS 0.25fF
C77699 INVX1_LOC_242/A VSS -0.73fF
C77700 INVX1_LOC_253/Y VSS 0.34fF
C77701 NOR2X1_LOC_836/A VSS 0.26fF
C77702 NOR2X1_LOC_847/B VSS 0.01fF
C77703 NOR2X1_LOC_847/A VSS 0.20fF
C77704 INVX1_LOC_63/A VSS 1.00fF
C77705 NOR2X1_LOC_814/A VSS 0.81fF
C77706 NOR2X1_LOC_862/B VSS 0.47fF
C77707 NOR2X1_LOC_808/B VSS 0.36fF
C77708 NOR2X1_LOC_591/A VSS 0.22fF
C77709 INVX1_LOC_4/Y VSS -6.48fF
C77710 INVX1_LOC_4/A VSS 0.73fF
C77711 INVX1_LOC_301/A VSS 0.48fF
C77712 INVX1_LOC_297/A VSS -0.06fF
C77713 NAND2X1_LOC_770/Y VSS 0.29fF
C77714 INVX1_LOC_306/Y VSS -3.06fF
C77715 INVX1_LOC_29/Y VSS 0.42fF
C77716 NOR2X1_LOC_258/Y VSS 0.11fF
C77717 NOR2X1_LOC_257/Y VSS 0.24fF
C77718 NOR2X1_LOC_445/B VSS -2.18fF
C77719 NOR2X1_LOC_342/A VSS 0.17fF
C77720 NOR2X1_LOC_247/Y VSS 0.12fF
C77721 NOR2X1_LOC_227/A VSS 0.38fF
C77722 INVX1_LOC_15/A VSS -7.74fF
C77723 NAND2X1_LOC_219/B VSS -0.16fF
C77724 NAND2X1_LOC_206/Y VSS 0.13fF
C77725 NOR2X1_LOC_461/Y VSS 0.11fF
C77726 NOR2X1_LOC_440/B VSS -0.15fF
C77727 NOR2X1_LOC_452/A VSS 0.09fF
C77728 NOR2X1_LOC_635/B VSS 0.25fF
C77729 NAND2X1_LOC_430/B VSS -0.09fF
C77730 NOR2X1_LOC_622/A VSS 0.03fF
C77731 NOR2X1_LOC_621/A VSS 0.08fF
C77732 NOR2X1_LOC_661/A VSS 0.05fF
C77733 INVX1_LOC_265/Y VSS 0.14fF
C77734 NOR2X1_LOC_676/Y VSS -0.20fF
C77735 NOR2X1_LOC_698/Y VSS 0.19fF
C77736 NOR2X1_LOC_665/Y VSS 0.14fF
C77737 NOR2X1_LOC_631/Y VSS -0.53fF
C77738 NOR2X1_LOC_685/Y VSS 0.04fF
C77739 NOR2X1_LOC_610/Y VSS 0.07fF
C77740 INVX1_LOC_29/A VSS -4.29fF
C77741 INVX1_LOC_9/A VSS 1.79fF
C77742 NOR2X1_LOC_76/B VSS 0.10fF
C77743 NOR2X1_LOC_197/B VSS 0.73fF
C77744 INVX1_LOC_296/Y VSS 0.24fF
C77745 INVX1_LOC_296/A VSS 0.32fF
C77746 INVX1_LOC_274/Y VSS 0.74fF
C77747 INVX1_LOC_263/Y VSS 0.15fF
C77748 INVX1_LOC_285/A VSS 0.58fF
C77749 INVX1_LOC_241/Y VSS 0.24fF
C77750 INVX1_LOC_230/A VSS 0.11fF
C77751 INVX1_LOC_252/A VSS 0.09fF
C77752 NOR2X1_LOC_109/Y VSS 0.56fF
C77753 NOR2X1_LOC_839/B VSS 0.31fF
C77754 INVX1_LOC_123/Y VSS 0.60fF
C77755 NOR2X1_LOC_863/A VSS 0.09fF
C77756 NOR2X1_LOC_852/Y VSS 0.25fF
C77757 NOR2X1_LOC_809/A VSS 0.11fF
C77758 NOR2X1_LOC_798/Y VSS 0.07fF
C77759 INVX1_LOC_3/Y VSS 0.56fF
C77760 NAND2X1_LOC_782/B VSS 0.55fF
C77761 INVX1_LOC_307/A VSS -1.65fF
C77762 NOR2X1_LOC_766/Y VSS -0.12fF
C77763 NOR2X1_LOC_291/Y VSS 0.33fF
C77764 NOR2X1_LOC_248/A VSS 0.12fF
C77765 NAND2X1_LOC_207/Y VSS 0.60fF
C77766 INVX1_LOC_3/A VSS 0.79fF
C77767 NOR2X1_LOC_259/A VSS 0.12fF
C77768 INVX1_LOC_117/A VSS 0.52fF
C77769 NAND2X1_LOC_205/A VSS 0.44fF
C77770 NOR2X1_LOC_72/Y VSS 0.07fF
C77771 INVX1_LOC_127/Y VSS 0.06fF
C77772 NOR2X1_LOC_461/B VSS 0.23fF
C77773 NOR2X1_LOC_384/A VSS 0.27fF
C77774 NOR2X1_LOC_476/B VSS 0.21fF
C77775 NOR2X1_LOC_833/B VSS 0.43fF
C77776 NOR2X1_LOC_450/B VSS 0.09fF
C77777 NOR2X1_LOC_405/Y VSS 0.11fF
C77778 INVX1_LOC_58/Y VSS 0.46fF
C77779 INVX1_LOC_181/A VSS 0.54fF
C77780 NOR2X1_LOC_438/Y VSS 0.19fF
C77781 NOR2X1_LOC_620/A VSS 0.12fF
C77782 NAND2X1_LOC_74/B VSS 0.96fF
C77783 NOR2X1_LOC_649/B VSS 1.40fF
C77784 NOR2X1_LOC_652/Y VSS -2.94fF
C77785 NOR2X1_LOC_686/A VSS 0.12fF
C77786 NOR2X1_LOC_697/Y VSS 0.16fF
C77787 INVX1_LOC_117/Y VSS -0.14fF
C77788 NOR2X1_LOC_81/Y VSS 0.13fF
C77789 INVX1_LOC_295/Y VSS 0.39fF
C77790 INVX1_LOC_262/A VSS 0.09fF
C77791 INVX1_LOC_273/A VSS -0.23fF
C77792 INVX1_LOC_251/A VSS 0.17fF
C77793 INVX1_LOC_284/A VSS 0.72fF
C77794 INVX1_LOC_240/Y VSS 0.19fF
C77795 NOR2X1_LOC_608/Y VSS 0.11fF
C77796 INVX1_LOC_46/Y VSS 0.67fF
C77797 NOR2X1_LOC_11/Y VSS -0.37fF
C77798 NOR2X1_LOC_36/B VSS 0.68fF
C77799 INVX1_LOC_118/A VSS 1.66fF
C77800 NOR2X1_LOC_849/A VSS 0.39fF
C77801 NOR2X1_LOC_863/B VSS 0.23fF
C77802 D_GATE_811 VSS 0.02fF
C77803 NOR2X1_LOC_810/Y VSS 0.14fF
C77804 NOR2X1_LOC_809/B VSS 0.31fF
C77805 NOR2X1_LOC_840/A VSS 0.11fF
C77806 INVX1_LOC_213/A VSS 0.26fF
C77807 NOR2X1_LOC_678/A VSS 0.41fF
C77808 NAND2X1_LOC_792/B VSS 0.27fF
C77809 NOR2X1_LOC_755/Y VSS 0.07fF
C77810 NOR2X1_LOC_743/Y VSS 0.47fF
C77811 NAND2X1_LOC_220/B VSS 0.14fF
C77812 INVX1_LOC_114/Y VSS 0.06fF
C77813 NOR2X1_LOC_259/B VSS 0.19fF
C77814 NOR2X1_LOC_342/B VSS 0.46fF
C77815 NAND2X1_LOC_206/B VSS 0.29fF
C77816 NOR2X1_LOC_243/B VSS -0.88fF
C77817 NAND2X1_LOC_85/Y VSS 0.20fF
C77818 INVX1_LOC_127/A VSS 0.12fF
C77819 NOR2X1_LOC_717/A VSS 0.77fF
C77820 NOR2X1_LOC_493/A VSS 0.25fF
C77821 NOR2X1_LOC_464/Y VSS 0.12fF
C77822 NOR2X1_LOC_465/Y VSS 0.58fF
C77823 NOR2X1_LOC_460/A VSS 0.08fF
C77824 NOR2X1_LOC_450/A VSS 0.12fF
C77825 NOR2X1_LOC_406/A VSS 0.30fF
C77826 INVX1_LOC_175/A VSS 0.49fF
C77827 NOR2X1_LOC_415/Y VSS 0.08fF
C77828 INVX1_LOC_90/Y VSS 0.25fF
C77829 INVX1_LOC_125/A VSS -0.22fF
C77830 INVX1_LOC_260/A VSS 0.11fF
C77831 NOR2X1_LOC_629/Y VSS -0.27fF
C77832 D_GATE_662 VSS 0.14fF
C77833 NAND2X1_LOC_82/Y VSS 0.46fF
C77834 INVX1_LOC_19/A VSS 1.30fF
C77835 NOR2X1_LOC_674/Y VSS 0.21fF
C77836 NOR2X1_LOC_696/Y VSS 0.26fF
C77837 NOR2X1_LOC_685/B VSS 0.19fF
C77838 INVX1_LOC_283/A VSS -0.02fF
C77839 INVX1_LOC_272/A VSS 0.15fF
C77840 INVX1_LOC_294/A VSS -0.06fF
C77841 NOR2X1_LOC_60/Y VSS 0.14fF
C77842 INVX1_LOC_253/A VSS 0.26fF
C77843 NAND2X1_LOC_618/Y VSS 0.30fF
C77844 INVX1_LOC_261/Y VSS 0.19fF
C77845 INVX1_LOC_261/A VSS 0.11fF
C77846 INVX1_LOC_250/Y VSS 0.28fF
C77847 INVX1_LOC_70/A VSS -0.13fF
C77848 INVX1_LOC_54/A VSS 0.84fF
C77849 NOR2X1_LOC_39/Y VSS 0.27fF
C77850 INVX1_LOC_23/Y VSS 0.45fF
C77851 NOR2X1_LOC_38/B VSS -1.30fF
C77852 D_GATE_865 VSS 0.02fF
C77853 NOR2X1_LOC_865/Y VSS 0.58fF
C77854 NOR2X1_LOC_856/A VSS 0.17fF
C77855 NOR2X1_LOC_729/A VSS 0.30fF
C77856 NOR2X1_LOC_812/A VSS 0.30fF
C77857 NOR2X1_LOC_801/A VSS 0.09fF
C77858 NOR2X1_LOC_499/B VSS 0.14fF
C77859 NAND2X1_LOC_793/B VSS 0.31fF
C77860 NOR2X1_LOC_754/Y VSS 0.16fF
C77861 NOR2X1_LOC_541/B VSS 0.35fF
C77862 NOR2X1_LOC_777/B VSS 0.55fF
C77863 NAND2X1_LOC_572/B VSS -0.90fF
C77864 NAND2X1_LOC_211/Y VSS 0.77fF
C77865 NOR2X1_LOC_65/Y VSS 0.15fF
C77866 NAND2X1_LOC_61/Y VSS 0.30fF
C77867 GATE_222 VSS 0.22fF
C77868 NOR2X1_LOC_240/A VSS 0.29fF
C77869 NOR2X1_LOC_492/Y VSS 0.10fF
C77870 INVX1_LOC_46/A VSS -4.50fF
C77871 INVX1_LOC_76/A VSS -20.09fF
C77872 NOR2X1_LOC_477/B VSS 0.11fF
C77873 NAND2X1_LOC_425/Y VSS 0.37fF
C77874 INVX1_LOC_193/A VSS 0.19fF
C77875 NOR2X1_LOC_378/Y VSS -0.04fF
C77876 NOR2X1_LOC_376/Y VSS 0.07fF
C77877 NAND2X1_LOC_453/A VSS -1.03fF
C77878 NOR2X1_LOC_422/Y VSS 0.08fF
C77879 NOR2X1_LOC_421/Y VSS 0.15fF
C77880 NOR2X1_LOC_416/A VSS -0.48fF
C77881 NOR2X1_LOC_414/Y VSS 0.30fF
C77882 INVX1_LOC_87/A VSS 0.51fF
C77883 INVX1_LOC_170/Y VSS 0.33fF
C77884 INVX1_LOC_168/Y VSS 0.25fF
C77885 NOR2X1_LOC_721/B VSS 0.32fF
C77886 NOR2X1_LOC_673/B VSS 0.13fF
C77887 NOR2X1_LOC_673/A VSS 0.58fF
C77888 NOR2X1_LOC_684/Y VSS 0.35fF
C77889 NOR2X1_LOC_663/A VSS 0.18fF
C77890 NOR2X1_LOC_660/Y VSS 0.94fF
C77891 NAND2X1_LOC_72/B VSS 0.32fF
C77892 NOR2X1_LOC_61/A VSS 0.26fF
C77893 NOR2X1_LOC_98/B VSS 0.34fF
C77894 NOR2X1_LOC_634/Y VSS 0.14fF
C77895 NOR2X1_LOC_654/A VSS -2.18fF
C77896 NOR2X1_LOC_638/Y VSS 0.07fF
C77897 NOR2X1_LOC_639/Y VSS 0.11fF
C77898 INVX1_LOC_271/Y VSS 0.29fF
C77899 INVX1_LOC_19/Y VSS -0.03fF
C77900 INVX1_LOC_293/Y VSS 0.54fF
C77901 INVX1_LOC_260/Y VSS 0.07fF
C77902 NOR2X1_LOC_646/B VSS 0.21fF
C77903 INVX1_LOC_16/Y VSS 0.50fF
C77904 NOR2X1_LOC_554/A VSS 0.34fF
C77905 NOR2X1_LOC_128/A VSS 0.12fF
C77906 NOR2X1_LOC_117/Y VSS 0.07fF
C77907 NOR2X1_LOC_137/Y VSS -0.12fF
C77908 INVX1_LOC_20/A VSS 0.86fF
C77909 NOR2X1_LOC_861/Y VSS 0.64fF
C77910 NOR2X1_LOC_856/B VSS 0.11fF
C77911 NOR2X1_LOC_841/A VSS -2.47fF
C77912 NOR2X1_LOC_592/B VSS 0.13fF
C77913 NOR2X1_LOC_435/A VSS 0.26fF
C77914 INVX1_LOC_299/Y VSS 0.45fF
C77915 NOR2X1_LOC_302/A VSS 0.12fF
C77916 NAND2X1_LOC_223/B VSS 0.30fF
C77917 NAND2X1_LOC_291/B VSS 0.35fF
C77918 NAND2X1_LOC_243/Y VSS 0.06fF
C77919 NAND2X1_LOC_267/B VSS 0.38fF
C77920 NAND2X1_LOC_175/Y VSS 0.34fF
C77921 INVX1_LOC_94/Y VSS -1.52fF
C77922 NAND2X1_LOC_207/B VSS 0.29fF
C77923 NOR2X1_LOC_491/Y VSS 0.19fF
C77924 D_GATE_479 VSS -0.05fF
C77925 INVX1_LOC_186/Y VSS -2.28fF
C77926 NAND2X1_LOC_798/B VSS 0.29fF
C77927 INVX1_LOC_180/Y VSS 0.06fF
C77928 NAND2X1_LOC_434/Y VSS 0.17fF
C77929 INVX1_LOC_166/Y VSS 0.31fF
C77930 NAND2X1_LOC_464/B VSS 0.41fF
C77931 NOR2X1_LOC_671/Y VSS 0.08fF
C77932 NOR2X1_LOC_662/A VSS 0.73fF
C77933 NOR2X1_LOC_653/Y VSS -0.27fF
C77934 NOR2X1_LOC_640/Y VSS 0.12fF
C77935 NOR2X1_LOC_641/Y VSS 0.11fF
C77936 NOR2X1_LOC_694/Y VSS 0.14fF
C77937 INVX1_LOC_77/Y VSS 0.24fF
C77938 NOR2X1_LOC_425/Y VSS 0.22fF
C77939 NOR2X1_LOC_683/Y VSS 0.07fF
C77940 NAND2X1_LOC_3/B VSS 0.69fF
C77941 NOR2X1_LOC_84/B VSS 0.07fF
C77942 NAND2X1_LOC_93/B VSS -4.78fF
C77943 INVX1_LOC_281/Y VSS 0.15fF
C77944 INVX1_LOC_281/A VSS 0.89fF
C77945 INVX1_LOC_292/Y VSS 0.44fF
C77946 INVX1_LOC_270/Y VSS 0.26fF
C77947 INVX1_LOC_270/A VSS 0.47fF
C77948 INVX1_LOC_18/Y VSS 0.09fF
C77949 INVX1_LOC_257/A VSS 0.28fF
C77950 NAND2X1_LOC_651/B VSS 0.17fF
C77951 INVX1_LOC_262/Y VSS 0.06fF
C77952 NOR2X1_LOC_105/Y VSS 0.22fF
C77953 NOR2X1_LOC_114/Y VSS -0.30fF
C77954 NOR2X1_LOC_127/Y VSS 0.27fF
C77955 NOR2X1_LOC_209/B VSS 0.44fF
C77956 NOR2X1_LOC_148/Y VSS 0.25fF
C77957 NOR2X1_LOC_36/A VSS 1.01fF
C77958 NOR2X1_LOC_48/Y VSS 0.19fF
C77959 NOR2X1_LOC_820/Y VSS 0.35fF
C77960 NOR2X1_LOC_866/B VSS 0.14fF
C77961 NOR2X1_LOC_863/Y VSS 0.09fF
C77962 NOR2X1_LOC_857/A VSS -1.36fF
C77963 NOR2X1_LOC_35/Y VSS -7.98fF
C77964 NOR2X1_LOC_301/A VSS 0.68fF
C77965 NOR2X1_LOC_850/B VSS 0.13fF
C77966 INVX1_LOC_99/A VSS 0.43fF
C77967 NOR2X1_LOC_830/Y VSS 0.04fF
C77968 NAND2X1_LOC_810/B VSS 0.11fF
C77969 NAND2X1_LOC_802/Y VSS 0.24fF
C77970 INVX1_LOC_143/Y VSS 0.47fF
C77971 NOR2X1_LOC_727/B VSS 0.58fF
C77972 NOR2X1_LOC_307/Y VSS 0.22fF
C77973 INVX1_LOC_109/Y VSS 0.29fF
C77974 INVX1_LOC_109/A VSS 0.84fF
C77975 INVX1_LOC_113/A VSS 0.65fF
C77976 NAND2X1_LOC_288/B VSS 0.51fF
C77977 NOR2X1_LOC_278/Y VSS 0.40fF
C77978 NOR2X1_LOC_240/B VSS 0.13fF
C77979 NOR2X1_LOC_235/Y VSS 0.07fF
C77980 NOR2X1_LOC_253/Y VSS 0.11fF
C77981 NAND2X1_LOC_223/A VSS 0.38fF
C77982 INVX1_LOC_104/Y VSS 0.25fF
C77983 NAND2X1_LOC_476/Y VSS 0.14fF
C77984 NAND2X1_LOC_475/Y VSS -2.38fF
C77985 INVX1_LOC_179/A VSS -0.39fF
C77986 NOR2X1_LOC_433/Y VSS 0.22fF
C77987 NAND2X1_LOC_469/B VSS 0.30fF
C77988 NOR2X1_LOC_449/A VSS 0.07fF
C77989 INVX1_LOC_167/A VSS 0.12fF
C77990 INVX1_LOC_163/Y VSS 0.19fF
C77991 NOR2X1_LOC_461/A VSS 0.17fF
C77992 NAND2X1_LOC_464/A VSS 0.25fF
C77993 NOR2X1_LOC_368/Y VSS 0.21fF
C77994 NOR2X1_LOC_693/Y VSS -0.05fF
C77995 NOR2X1_LOC_655/Y VSS 0.18fF
C77996 NOR2X1_LOC_656/Y VSS 0.11fF
C77997 INVX1_LOC_28/Y VSS -0.10fF
C77998 NAND2X1_LOC_637/Y VSS -0.09fF
C77999 NAND2X1_LOC_655/B VSS 0.13fF
C78000 NAND2X1_LOC_642/Y VSS 0.36fF
C78001 NAND2X1_LOC_81/B VSS -0.13fF
C78002 INVX1_LOC_291/A VSS -0.93fF
C78003 INVX1_LOC_280/A VSS 1.18fF
C78004 NOR2X1_LOC_603/Y VSS 0.07fF
C78005 NOR2X1_LOC_629/A VSS 0.12fF
C78006 INVX1_LOC_23/A VSS 1.40fF
C78007 NOR2X1_LOC_621/B VSS 0.13fF
C78008 NOR2X1_LOC_137/B VSS 0.17fF
C78009 NOR2X1_LOC_58/Y VSS 0.21fF
C78010 NOR2X1_LOC_69/A VSS 0.12fF
C78011 NOR2X1_LOC_25/Y VSS 0.41fF
C78012 NOR2X1_LOC_30/Y VSS 0.50fF
C78013 NOR2X1_LOC_831/Y VSS -0.99fF
C78014 NAND2X1_LOC_811/B VSS 0.26fF
C78015 NAND2X1_LOC_804/Y VSS 0.34fF
C78016 NOR2X1_LOC_318/A VSS 0.20fF
C78017 NOR2X1_LOC_329/Y VSS 0.34fF
C78018 INVX1_LOC_119/Y VSS 0.43fF
C78019 INVX1_LOC_108/A VSS 0.34fF
C78020 INVX1_LOC_115/A VSS 0.66fF
C78021 NAND2X1_LOC_212/Y VSS -0.16fF
C78022 NAND2X1_LOC_288/A VSS 0.51fF
C78023 INVX1_LOC_131/Y VSS -0.28fF
C78024 NAND2X1_LOC_244/A VSS 0.36fF
C78025 NAND2X1_LOC_241/Y VSS 0.11fF
C78026 INVX1_LOC_129/A VSS 0.26fF
C78027 NAND2X1_LOC_470/B VSS 0.29fF
C78028 NAND2X1_LOC_452/Y VSS -0.07fF
C78029 NAND2X1_LOC_254/Y VSS 0.40fF
C78030 INVX1_LOC_203/A VSS -1.57fF
C78031 NAND2X1_LOC_477/Y VSS 0.23fF
C78032 NOR2X1_LOC_487/Y VSS -0.11fF
C78033 NAND2X1_LOC_402/B VSS 0.34fF
C78034 NOR2X1_LOC_395/Y VSS 0.05fF
C78035 NAND2X1_LOC_455/B VSS 0.32fF
C78036 NOR2X1_LOC_634/A VSS 0.55fF
C78037 NOR2X1_LOC_692/Y VSS -0.32fF
C78038 NOR2X1_LOC_670/Y VSS 0.46fF
C78039 NOR2X1_LOC_383/B VSS 0.75fF
C78040 INVX1_LOC_21/Y VSS -0.06fF
C78041 INVX1_LOC_290/Y VSS 0.33fF
C78042 INVX1_LOC_49/Y VSS 0.61fF
C78043 INVX1_LOC_27/Y VSS 0.35fF
C78044 INVX1_LOC_38/A VSS -4.43fF
C78045 NOR2X1_LOC_586/Y VSS -0.23fF
C78046 NOR2X1_LOC_585/Y VSS 0.12fF
C78047 NAND2X1_LOC_655/A VSS 0.40fF
C78048 INVX1_LOC_264/Y VSS 0.06fF
C78049 NOR2X1_LOC_623/B VSS 0.27fF
C78050 NOR2X1_LOC_605/A VSS 0.22fF
C78051 INVX1_LOC_91/A VSS 1.24fF
C78052 INVX1_LOC_57/A VSS -5.70fF
C78053 NOR2X1_LOC_170/A VSS -0.05fF
C78054 INVX1_LOC_35/Y VSS 0.48fF
C78055 INVX1_LOC_66/Y VSS -0.09fF
C78056 NOR2X1_LOC_125/Y VSS 0.34fF
C78057 NOR2X1_LOC_158/Y VSS 0.28fF
C78058 NOR2X1_LOC_158/B VSS 0.07fF
C78059 NOR2X1_LOC_68/Y VSS 0.15fF
C78060 NOR2X1_LOC_79/Y VSS 0.11fF
C78061 NOR2X1_LOC_79/A VSS 0.22fF
C78062 INVX1_LOC_44/A VSS -0.32fF
C78063 NOR2X1_LOC_24/Y VSS 0.09fF
C78064 NOR2X1_LOC_33/Y VSS 0.07fF
C78065 NOR2X1_LOC_34/Y VSS 0.09fF
C78066 NOR2X1_LOC_48/B VSS 0.82fF
C78067 NOR2X1_LOC_865/A VSS 0.31fF
C78068 NOR2X1_LOC_859/Y VSS 0.19fF
C78069 NOR2X1_LOC_833/Y VSS -0.04fF
C78070 NOR2X1_LOC_858/A VSS 0.27fF
C78071 NOR2X1_LOC_840/Y VSS -0.01fF
C78072 NOR2X1_LOC_855/A VSS 0.25fF
C78073 NOR2X1_LOC_820/B VSS 0.13fF
C78074 INVX1_LOC_84/A VSS -5.55fF
C78075 INVX1_LOC_152/A VSS 0.56fF
C78076 NOR2X1_LOC_61/Y VSS 0.40fF
C78077 NOR2X1_LOC_332/Y VSS -0.02fF
C78078 NOR2X1_LOC_319/B VSS 0.11fF
C78079 INPUT_4 VSS -0.45fF
C78080 NOR2X1_LOC_340/A VSS -0.59fF
C78081 NOR2X1_LOC_509/A VSS -0.11fF
C78082 INVX1_LOC_107/Y VSS 0.44fF
C78083 INVX1_LOC_118/Y VSS 0.49fF
C78084 INVX1_LOC_129/Y VSS 0.21fF
C78085 NOR2X1_LOC_275/A VSS 0.12fF
C78086 NAND2X1_LOC_286/B VSS 0.53fF
C78087 NOR2X1_LOC_282/Y VSS 0.06fF
C78088 NOR2X1_LOC_281/Y VSS 0.07fF
C78089 NOR2X1_LOC_297/A VSS 0.23fF
C78090 INVX1_LOC_32/A VSS -8.05fF
C78091 NOR2X1_LOC_231/A VSS 0.12fF
C78092 NOR2X1_LOC_448/A VSS 0.12fF
C78093 NAND2X1_LOC_454/Y VSS 0.35fF
C78094 INVX1_LOC_185/A VSS 0.34fF
C78095 NAND2X1_LOC_465/A VSS 0.25fF
C78096 NAND2X1_LOC_471/Y VSS 0.38fF
C78097 NAND2X1_LOC_500/B VSS 0.11fF
C78098 NOR2X1_LOC_489/A VSS 0.41fF
C78099 INVX1_LOC_165/A VSS 0.12fF
C78100 NOR2X1_LOC_394/Y VSS 0.07fF
C78101 NOR2X1_LOC_393/Y VSS 0.07fF
C78102 NOR2X1_LOC_691/B VSS 0.28fF
C78103 NOR2X1_LOC_691/A VSS 0.23fF
C78104 INVX1_LOC_274/A VSS 0.55fF
C78105 NOR2X1_LOC_331/B VSS 1.11fF
C78106 INVX1_LOC_37/Y VSS 0.54fF
C78107 INVX1_LOC_37/A VSS 1.22fF
C78108 INVX1_LOC_59/Y VSS 0.54fF
C78109 INVX1_LOC_26/Y VSS 0.35fF
C78110 INVX1_LOC_26/A VSS 0.89fF
C78111 NOR2X1_LOC_584/Y VSS 0.12fF
C78112 NOR2X1_LOC_583/Y VSS 0.07fF
C78113 NOR2X1_LOC_631/A VSS 0.12fF
C78114 INVX1_LOC_136/Y VSS 0.19fF
C78115 NOR2X1_LOC_66/Y VSS -0.19fF
C78116 NAND2X1_LOC_656/B VSS 0.11fF
C78117 NOR2X1_LOC_612/Y VSS 0.20fF
C78118 NAND2X1_LOC_659/B VSS 0.72fF
C78119 INVX1_LOC_255/A VSS 0.34fF
C78120 NOR2X1_LOC_720/A VSS 0.23fF
C78121 NOR2X1_LOC_668/Y VSS 0.12fF
C78122 NOR2X1_LOC_754/A VSS 0.11fF
C78123 NOR2X1_LOC_179/Y VSS 0.16fF
C78124 INVX1_LOC_75/Y VSS 0.22fF
C78125 NOR2X1_LOC_536/A VSS 1.47fF
C78126 INVX1_LOC_74/A VSS 0.48fF
C78127 NOR2X1_LOC_114/A VSS 0.29fF
C78128 NOR2X1_LOC_67/Y VSS -0.39fF
C78129 NOR2X1_LOC_78/Y VSS -0.17fF
C78130 NOR2X1_LOC_56/Y VSS -1.50fF
C78131 NOR2X1_LOC_1/Y VSS 0.03fF
C78132 NOR2X1_LOC_860/Y VSS 0.06fF
C78133 NOR2X1_LOC_858/B VSS 0.22fF
C78134 NOR2X1_LOC_829/A VSS 0.16fF
C78135 NOR2X1_LOC_409/B VSS 0.12fF
C78136 NAND2X1_LOC_807/B VSS 0.39fF
C78137 INVX1_LOC_133/A VSS 0.69fF
C78138 NAND2X1_LOC_836/Y VSS 0.18fF
C78139 NOR2X1_LOC_80/Y VSS 0.17fF
C78140 NAND2X1_LOC_63/Y VSS 0.72fF
C78141 NOR2X1_LOC_305/Y VSS 0.25fF
C78142 NOR2X1_LOC_334/Y VSS 0.24fF
C78143 NOR2X1_LOC_519/Y VSS 0.11fF
C78144 NOR2X1_LOC_510/B VSS 0.37fF
C78145 NOR2X1_LOC_506/Y VSS -0.05fF
C78146 INVX1_LOC_139/Y VSS 0.39fF
C78147 INVX1_LOC_139/A VSS 0.68fF
C78148 INVX1_LOC_128/Y VSS 0.06fF
C78149 INVX1_LOC_128/A VSS 0.11fF
C78150 INVX1_LOC_106/Y VSS 0.08fF
C78151 INVX1_LOC_106/A VSS 0.09fF
C78152 NOR2X1_LOC_831/B VSS 0.63fF
C78153 NOR2X1_LOC_155/A VSS 0.51fF
C78154 NAND2X1_LOC_287/B VSS -0.81fF
C78155 NOR2X1_LOC_280/Y VSS 0.26fF
C78156 NOR2X1_LOC_279/Y VSS 0.07fF
C78157 NOR2X1_LOC_843/B VSS 0.60fF
C78158 NOR2X1_LOC_346/A VSS -0.09fF
C78159 NAND2X1_LOC_243/B VSS 0.31fF
C78160 NOR2X1_LOC_266/B VSS 0.46fF
C78161 INVX1_LOC_309/A VSS -0.03fF
C78162 NOR2X1_LOC_435/B VSS 0.15fF
C78163 INVX1_LOC_202/Y VSS 0.06fF
C78164 NAND2X1_LOC_472/Y VSS 1.24fF
C78165 NAND2X1_LOC_447/Y VSS 0.59fF
C78166 INVX1_LOC_188/Y VSS 0.15fF
C78167 NOR2X1_LOC_501/B VSS 0.13fF
C78168 NAND2X1_LOC_444/B VSS 0.11fF
C78169 INVX1_LOC_12/A VSS -7.10fF
C78170 NAND2X1_LOC_456/Y VSS 0.07fF
C78171 INVX1_LOC_47/Y VSS 0.38fF
C78172 NAND2X1_LOC_639/A VSS 0.73fF
C78173 INVX1_LOC_247/A VSS -0.65fF
C78174 NOR2X1_LOC_601/Y VSS 0.14fF
C78175 NOR2X1_LOC_600/Y VSS 0.25fF
C78176 NOR2X1_LOC_728/B VSS 0.26fF
C78177 NAND2X1_LOC_647/B VSS 0.40fF
C78178 NOR2X1_LOC_609/Y VSS 0.06fF
C78179 NOR2X1_LOC_669/A VSS 0.12fF
C78180 NAND2X1_LOC_659/A VSS -0.73fF
C78181 NAND2X1_LOC_574/A VSS 0.13fF
C78182 NAND2X1_LOC_141/Y VSS 0.34fF
C78183 NOR2X1_LOC_124/A VSS -0.23fF
C78184 INVX1_LOC_78/A VSS 1.52fF
C78185 NOR2X1_LOC_216/B VSS 0.66fF
C78186 NOR2X1_LOC_99/Y VSS -0.46fF
C78187 NOR2X1_LOC_332/B VSS 0.35fF
C78188 NOR2X1_LOC_167/Y VSS 0.26fF
C78189 INVX1_LOC_102/A VSS -2.33fF
C78190 NOR2X1_LOC_156/Y VSS -0.26fF
C78191 NOR2X1_LOC_145/Y VSS 0.13fF
C78192 NOR2X1_LOC_89/A VSS -4.65fF
C78193 NOR2X1_LOC_88/Y VSS 0.35fF
C78194 NOR2X1_LOC_88/A VSS 0.27fF
C78195 NOR2X1_LOC_392/Y VSS -5.03fF
C78196 NAND2X1_LOC_859/B VSS 0.43fF
C78197 NAND2X1_LOC_837/Y VSS 0.41fF
C78198 INVX1_LOC_309/Y VSS 0.30fF
C78199 NAND2X1_LOC_807/A VSS 0.19fF
C78200 NAND2X1_LOC_793/Y VSS 0.52fF
C78201 INVX1_LOC_308/Y VSS 0.30fF
C78202 NOR2X1_LOC_846/A VSS 0.23fF
C78203 INVX1_LOC_38/Y VSS 0.43fF
C78204 INVX1_LOC_149/Y VSS 0.18fF
C78205 NOR2X1_LOC_324/Y VSS 0.07fF
C78206 NOR2X1_LOC_325/Y VSS 0.07fF
C78207 NOR2X1_LOC_348/Y VSS 0.37fF
C78208 NOR2X1_LOC_304/Y VSS 0.44fF
C78209 NOR2X1_LOC_53/Y VSS 0.21fF
C78210 INVX1_LOC_210/A VSS 0.14fF
C78211 INVX1_LOC_138/Y VSS 0.32fF
C78212 INVX1_LOC_138/A VSS 0.09fF
C78213 INVX1_LOC_105/Y VSS 0.22fF
C78214 INVX1_LOC_116/Y VSS 0.39fF
C78215 NOR2X1_LOC_274/B VSS 0.68fF
C78216 NOR2X1_LOC_345/A VSS 0.26fF
C78217 NOR2X1_LOC_343/B VSS 0.09fF
C78218 NOR2X1_LOC_249/Y VSS 0.24fF
C78219 INVX1_LOC_50/Y VSS -3.55fF
C78220 INVX1_LOC_308/A VSS 0.09fF
C78221 NOR2X1_LOC_447/A VSS 0.24fF
C78222 NAND2X1_LOC_466/A VSS 0.19fF
C78223 NOR2X1_LOC_500/B VSS 0.55fF
C78224 NAND2X1_LOC_474/Y VSS 0.56fF
C78225 INVX1_LOC_171/Y VSS 0.14fF
C78226 NOR2X1_LOC_434/A VSS 0.12fF
C78227 INVX1_LOC_53/A VSS 1.32fF
C78228 INVX1_LOC_183/A VSS 0.12fF
C78229 NAND2X1_LOC_787/B VSS 0.34fF
C78230 NOR2X1_LOC_484/Y VSS 0.07fF
C78231 INVX1_LOC_79/Y VSS 0.15fF
C78232 INVX1_LOC_68/A VSS 0.09fF
C78233 INVX1_LOC_271/A VSS 1.08fF
C78234 NOR2X1_LOC_677/Y VSS -0.23fF
C78235 NOR2X1_LOC_720/B VSS 0.36fF
C78236 NOR2X1_LOC_264/Y VSS 0.32fF
C78237 NOR2X1_LOC_688/Y VSS 0.06fF
C78238 INVX1_LOC_22/Y VSS 0.31fF
C78239 INVX1_LOC_24/Y VSS 0.60fF
C78240 INVX1_LOC_263/A VSS -0.01fF
C78241 INVX1_LOC_252/Y VSS 0.06fF
C78242 NAND2X1_LOC_624/B VSS 0.31fF
C78243 NOR2X1_LOC_177/Y VSS 0.24fF
C78244 NAND2X1_LOC_86/Y VSS 0.13fF
C78245 NOR2X1_LOC_196/Y VSS 0.06fF
C78246 NOR2X1_LOC_166/Y VSS 0.14fF
C78247 NOR2X1_LOC_188/Y VSS 0.17fF
C78248 NOR2X1_LOC_156/A VSS 0.11fF
C78249 NOR2X1_LOC_98/A VSS 0.12fF
C78250 NOR2X1_LOC_9/Y VSS 0.57fF
C78251 NOR2X1_LOC_76/A VSS 0.49fF
C78252 NOR2X1_LOC_32/Y VSS 0.19fF
C78253 INVX1_LOC_22/A VSS 1.73fF
C78254 NOR2X1_LOC_87/Y VSS 0.10fF
C78255 NOR2X1_LOC_87/B VSS 0.33fF
C78256 NOR2X1_LOC_43/Y VSS 0.30fF
C78257 NOR2X1_LOC_846/B VSS 0.13fF
C78258 NOR2X1_LOC_814/Y VSS 0.05fF
C78259 INVX1_LOC_316/Y VSS 0.21fF
C78260 NAND2X1_LOC_848/Y VSS 0.15fF
C78261 NOR2X1_LOC_825/Y VSS 0.12fF
C78262 NOR2X1_LOC_837/A VSS 0.12fF
C78263 NAND2X1_LOC_795/Y VSS 0.00fF
C78264 INVX1_LOC_71/Y VSS 0.10fF
C78265 NOR2X1_LOC_360/A VSS 0.09fF
C78266 NOR2X1_LOC_346/Y VSS 0.09fF
C78267 NOR2X1_LOC_337/A VSS 0.23fF
C78268 NOR2X1_LOC_703/A VSS -0.40fF
C78269 NOR2X1_LOC_374/B VSS 0.30fF
C78270 NOR2X1_LOC_325/A VSS 0.09fF
C78271 NOR2X1_LOC_364/A VSS -0.41fF
C78272 INVX1_LOC_157/Y VSS 0.21fF
C78273 NOR2X1_LOC_351/Y VSS 0.55fF
C78274 NOR2X1_LOC_314/Y VSS 0.11fF
C78275 NOR2X1_LOC_302/Y VSS 0.26fF
C78276 NOR2X1_LOC_537/Y VSS 0.37fF
C78277 NOR2X1_LOC_538/Y VSS 0.09fF
C78278 NOR2X1_LOC_447/B VSS 0.47fF
C78279 INVX1_LOC_115/Y VSS 0.15fF
C78280 INVX1_LOC_159/Y VSS 0.15fF
C78281 INVX1_LOC_126/Y VSS 0.41fF
C78282 INVX1_LOC_148/Y VSS 0.44fF
C78283 INVX1_LOC_137/Y VSS 0.25fF
C78284 INVX1_LOC_137/A VSS 0.52fF
C78285 NOR2X1_LOC_709/A VSS 0.79fF
C78286 NOR2X1_LOC_261/A VSS 0.12fF
C78287 NOR2X1_LOC_269/Y VSS 0.56fF
C78288 INPUT_1 VSS 0.87fF
C78289 INVX1_LOC_307/Y VSS 0.28fF
C78290 NAND2X1_LOC_573/A VSS 0.67fF
C78291 NAND2X1_LOC_392/Y VSS 0.03fF
C78292 NAND2X1_LOC_451/Y VSS 0.57fF
C78293 INVX1_LOC_192/Y VSS 0.35fF
C78294 NOR2X1_LOC_451/A VSS 0.29fF
C78295 INVX1_LOC_194/Y VSS 0.25fF
C78296 NOR2X1_LOC_545/B VSS 0.27fF
C78297 INVX1_LOC_78/Y VSS 0.39fF
C78298 INVX1_LOC_67/Y VSS 0.34fF
C78299 INVX1_LOC_56/Y VSS 0.44fF
C78300 INVX1_LOC_56/A VSS 0.11fF
C78301 INVX1_LOC_34/Y VSS 0.61fF
C78302 INVX1_LOC_89/Y VSS 0.23fF
C78303 INVX1_LOC_12/Y VSS 1.26fF
C78304 NAND2X1_LOC_648/A VSS 0.26fF
C78305 NAND2X1_LOC_660/A VSS 0.33fF
C78306 INVX1_LOC_14/Y VSS 1.05fF
C78307 NAND2X1_LOC_624/A VSS 0.24fF
C78308 NOR2X1_LOC_719/A VSS 0.48fF
C78309 NOR2X1_LOC_121/A VSS 0.12fF
C78310 NOR2X1_LOC_278/A VSS 0.34fF
C78311 NOR2X1_LOC_602/B VSS 0.07fF
C78312 NOR2X1_LOC_208/A VSS 0.19fF
C78313 NOR2X1_LOC_197/Y VSS 0.09fF
C78314 INVX1_LOC_8/A VSS 0.91fF
C78315 NOR2X1_LOC_176/Y VSS 0.15fF
C78316 NOR2X1_LOC_74/A VSS 0.64fF
C78317 NOR2X1_LOC_156/B VSS -0.20fF
C78318 D_INPUT_3 VSS -2.51fF
C78319 NOR2X1_LOC_99/B VSS 0.01fF
C78320 NOR2X1_LOC_97/B VSS 0.25fF
C78321 NOR2X1_LOC_19/Y VSS 0.12fF
C78322 INPUT_5 VSS 0.11fF
C78323 NOR2X1_LOC_51/A VSS 0.49fF
C78324 NOR2X1_LOC_815/A VSS 0.32fF
C78325 NAND2X1_LOC_808/A VSS 0.73fF
C78326 NAND2X1_LOC_796/Y VSS 0.19fF
C78327 NAND2X1_LOC_862/A VSS -0.06fF
C78328 NAND2X1_LOC_850/Y VSS 0.83fF
C78329 INVX1_LOC_315/A VSS 0.44fF
C78330 NAND2X1_LOC_96/A VSS 0.69fF
C78331 NOR2X1_LOC_824/Y VSS -0.08fF
C78332 NOR2X1_LOC_823/Y VSS 0.07fF
C78333 INVX1_LOC_6/A VSS -3.43fF
C78334 INVX1_LOC_150/A VSS 0.08fF
C78335 NOR2X1_LOC_352/Y VSS 0.21fF
C78336 NOR2X1_LOC_353/Y VSS 0.09fF
C78337 NOR2X1_LOC_324/B VSS 0.28fF
C78338 NOR2X1_LOC_324/A VSS 0.40fF
C78339 NOR2X1_LOC_313/Y VSS 0.13fF
C78340 NOR2X1_LOC_302/B VSS 0.13fF
C78341 NOR2X1_LOC_516/Y VSS 0.20fF
C78342 NOR2X1_LOC_527/Y VSS 0.15fF
C78343 NOR2X1_LOC_565/B VSS 0.07fF
C78344 INVX1_LOC_220/Y VSS 0.24fF
C78345 NOR2X1_LOC_548/Y VSS 0.43fF
C78346 NOR2X1_LOC_505/Y VSS 0.03fF
C78347 INVX1_LOC_103/Y VSS 0.15fF
C78348 INVX1_LOC_114/A VSS 0.09fF
C78349 INVX1_LOC_147/Y VSS 0.25fF
C78350 INVX1_LOC_125/Y VSS 0.59fF
C78351 INVX1_LOC_158/Y VSS 0.47fF
C78352 INVX1_LOC_169/Y VSS 0.15fF
C78353 INVX1_LOC_169/A VSS -0.07fF
C78354 NOR2X1_LOC_719/B VSS 0.20fF
C78355 NOR2X1_LOC_346/B VSS 0.41fF
C78356 NOR2X1_LOC_285/B VSS 0.32fF
C78357 NOR2X1_LOC_368/A VSS 0.41fF
C78358 INVX1_LOC_306/A VSS 0.56fF
C78359 NOR2X1_LOC_486/B VSS 0.30fF
C78360 NAND2X1_LOC_468/B VSS 0.63fF
C78361 INVX1_LOC_201/A VSS 0.08fF
C78362 INVX1_LOC_175/Y VSS 0.42fF
C78363 INVX1_LOC_44/Y VSS 0.15fF
C78364 INVX1_LOC_88/Y VSS 0.33fF
C78365 INVX1_LOC_11/Y VSS -0.82fF
C78366 INVX1_LOC_66/A VSS 0.25fF
C78367 NAND2X1_LOC_661/B VSS 0.31fF
C78368 INVX1_LOC_266/Y VSS 0.42fF
C78369 NOR2X1_LOC_679/B VSS 0.07fF
C78370 NAND2X1_LOC_800/A VSS 0.42fF
C78371 NAND2X1_LOC_649/B VSS 0.31fF
C78372 NOR2X1_LOC_595/Y VSS 0.01fF
C78373 NAND2X1_LOC_622/B VSS 0.33fF
C78374 NAND2X1_LOC_735/B VSS 0.25fF
C78375 NOR2X1_LOC_612/B VSS 0.67fF
C78376 NOR2X1_LOC_709/B VSS 0.14fF
C78377 NOR2X1_LOC_164/Y VSS 0.48fF
C78378 NOR2X1_LOC_211/A VSS -0.68fF
C78379 NOR2X1_LOC_131/Y VSS 0.21fF
C78380 NOR2X1_LOC_131/A VSS 0.12fF
C78381 NOR2X1_LOC_86/A VSS 0.84fF
C78382 INVX1_LOC_16/A VSS 0.92fF
C78383 INVX1_LOC_25/Y VSS 0.45fF
C78384 NOR2X1_LOC_96/Y VSS 0.12fF
C78385 NOR2X1_LOC_94/Y VSS 0.09fF
C78386 NOR2X1_LOC_74/Y VSS -0.26fF
C78387 NAND2X1_LOC_863/B VSS 0.38fF
C78388 NAND2X1_LOC_853/Y VSS 0.61fF
C78389 NAND2X1_LOC_852/Y VSS 1.11fF
C78390 NAND2X1_LOC_799/Y VSS 0.25fF
C78391 NAND2X1_LOC_848/A VSS -3.46fF
C78392 NOR2X1_LOC_816/Y VSS 0.02fF
C78393 NOR2X1_LOC_845/A VSS 0.64fF
C78394 INVX1_LOC_123/A VSS 0.97fF
C78395 INVX1_LOC_48/A VSS 0.72fF
C78396 NAND2X1_LOC_839/A VSS 0.40fF
C78397 NOR2X1_LOC_822/Y VSS -0.16fF
C78398 NOR2X1_LOC_821/Y VSS 0.07fF
C78399 INVX1_LOC_122/A VSS 0.34fF
C78400 VDD VSS 2.56fF
C78401 NOR2X1_LOC_334/A VSS -0.19fF
C78402 NOR2X1_LOC_111/A VSS 0.39fF
C78403 INVX1_LOC_160/A VSS -0.61fF
C78404 NOR2X1_LOC_354/Y VSS -0.09fF
C78405 D_GATE_366 VSS 0.16fF
C78406 NOR2X1_LOC_366/Y VSS 0.01fF
C78407 NOR2X1_LOC_377/Y VSS 0.16fF
C78408 NOR2X1_LOC_560/A VSS 0.11fF
C78409 INVX1_LOC_216/A VSS 0.25fF
C78410 NOR2X1_LOC_514/Y VSS 0.09fF
C78411 NOR2X1_LOC_548/B VSS 0.48fF
C78412 NOR2X1_LOC_548/A VSS 0.22fF
C78413 INVX1_LOC_179/Y VSS -0.01fF
C78414 INVX1_LOC_113/Y VSS 0.34fF
C78415 INVX1_LOC_146/Y VSS 0.33fF
C78416 INVX1_LOC_102/Y VSS 0.53fF
C78417 INVX1_LOC_168/A VSS -0.09fF
C78418 NOR2X1_LOC_542/B VSS 0.26fF
C78419 NOR2X1_LOC_730/A VSS -0.12fF
C78420 NOR2X1_LOC_687/Y VSS -0.67fF
C78421 INVX1_LOC_249/Y VSS 0.23fF
C78422 NOR2X1_LOC_712/B VSS 0.15fF
C78423 NOR2X1_LOC_707/A VSS 0.22fF
C78424 INVX1_LOC_316/A VSS 0.22fF
C78425 INVX1_LOC_191/A VSS 0.42fF
C78426 NOR2X1_LOC_427/Y VSS 0.06fF
C78427 INVX1_LOC_196/Y VSS 0.13fF
C78428 NAND2X1_LOC_462/B VSS -0.15fF
C78429 NOR2X1_LOC_482/Y VSS 0.14fF
C78430 INVX1_LOC_87/Y VSS 0.15fF
C78431 INVX1_LOC_32/Y VSS 0.28fF
C78432 INVX1_LOC_76/Y VSS 0.25fF
C78433 INVX1_LOC_10/Y VSS 0.28fF
C78434 INVX1_LOC_65/Y VSS 0.26fF
C78435 INVX1_LOC_43/A VSS 0.14fF
C78436 INVX1_LOC_275/A VSS -0.14fF
C78437 NOR2X1_LOC_708/A VSS 0.34fF
C78438 NAND2X1_LOC_661/A VSS 0.23fF
C78439 NAND2X1_LOC_652/Y VSS 0.34fF
C78440 NOR2X1_LOC_665/A VSS 0.01fF
C78441 NAND2X1_LOC_632/B VSS 0.27fF
C78442 NOR2X1_LOC_625/Y VSS 0.11fF
C78443 INVX1_LOC_176/A VSS 0.49fF
C78444 NAND2X1_LOC_623/B VSS 0.26fF
C78445 NOR2X1_LOC_528/Y VSS -1.99fF
C78446 NOR2X1_LOC_188/A VSS 0.63fF
C78447 NOR2X1_LOC_130/Y VSS 0.11fF
C78448 NOR2X1_LOC_130/A VSS -1.29fF
C78449 NOR2X1_LOC_175/A VSS 0.35fF
C78450 NOR2X1_LOC_152/Y VSS 0.80fF
C78451 NOR2X1_LOC_152/A VSS 0.18fF
C78452 NOR2X1_LOC_657/B VSS 0.55fF
C78453 NOR2X1_LOC_139/Y VSS 0.03fF
C78454 NOR2X1_LOC_163/Y VSS -0.08fF
C78455 NOR2X1_LOC_163/A VSS 0.31fF
C78456 INVX1_LOC_71/A VSS 1.13fF
C78457 INVX1_LOC_65/A VSS 1.00fF
C78458 NOR2X1_LOC_84/Y VSS -4.17fF
C78459 NOR2X1_LOC_84/A VSS -0.15fF
C78460 NAND2X1_LOC_863/A VSS 0.32fF
C78461 NAND2X1_LOC_855/Y VSS 0.13fF
C78462 NAND2X1_LOC_809/A VSS 0.23fF
C78463 NAND2X1_LOC_800/Y VSS 0.06fF
C78464 NAND2X1_LOC_840/B VSS 0.33fF
C78465 GATE_811 VSS 0.22fF
C78466 NAND2X1_LOC_811/Y VSS 0.22fF
C78467 NAND2X1_LOC_849/B VSS 0.11fF
C78468 NOR2X1_LOC_813/Y VSS 0.26fF
C78469 NAND2X1_LOC_721/A VSS 0.60fF
C78470 NOR2X1_LOC_836/B VSS 0.22fF
C78471 INVX1_LOC_148/A VSS -0.19fF
C78472 NOR2X1_LOC_174/B VSS 0.20fF
C78473 NOR2X1_LOC_333/A VSS 0.12fF
C78474 NOR2X1_LOC_399/Y VSS 0.36fF
C78475 NOR2X1_LOC_399/A VSS 0.31fF
C78476 INVX1_LOC_33/Y VSS 0.68fF
C78477 NOR2X1_LOC_311/Y VSS 0.24fF
C78478 NOR2X1_LOC_356/A VSS -1.11fF
C78479 NOR2X1_LOC_348/B VSS 0.18fF
C78480 NOR2X1_LOC_254/Y VSS 0.26fF
C78481 NOR2X1_LOC_344/A VSS -0.37fF
C78482 NOR2X1_LOC_363/Y VSS -0.53fF
C78483 NOR2X1_LOC_564/Y VSS 0.12fF
C78484 NOR2X1_LOC_525/Y VSS 0.31fF
C78485 INVX1_LOC_10/A VSS 0.90fF
C78486 INVX1_LOC_226/A VSS 0.18fF
C78487 NOR2X1_LOC_547/B VSS -0.05fF
C78488 NOR2X1_LOC_561/A VSS 0.14fF
C78489 NOR2X1_LOC_558/A VSS 0.19fF
C78490 INVX1_LOC_189/Y VSS 0.15fF
C78491 INVX1_LOC_189/A VSS 0.29fF
C78492 INVX1_LOC_178/Y VSS 0.05fF
C78493 INVX1_LOC_167/Y VSS 0.42fF
C78494 INVX1_LOC_156/A VSS 0.09fF
C78495 INVX1_LOC_101/A VSS 0.30fF
C78496 INVX1_LOC_134/Y VSS 0.28fF
C78497 INVX1_LOC_112/A VSS 0.11fF
C78498 NOR2X1_LOC_730/B VSS 0.07fF
C78499 NOR2X1_LOC_730/Y VSS 0.43fF
C78500 NOR2X1_LOC_634/B VSS 0.28fF
C78501 NOR2X1_LOC_706/B VSS 0.28fF
C78502 INVX1_LOC_304/A VSS 0.08fF
C78503 INVX1_LOC_315/Y VSS -0.31fF
C78504 NAND2X1_LOC_463/B VSS -1.43fF
C78505 NOR2X1_LOC_409/Y VSS 0.20fF
C78506 NOR2X1_LOC_380/Y VSS 0.18fF
C78507 NAND2X1_LOC_465/Y VSS -0.19fF
C78508 NAND2X1_LOC_464/Y VSS 0.11fF
C78509 INVX1_LOC_86/A VSS 0.22fF
C78510 INVX1_LOC_97/A VSS 0.09fF
C78511 INVX1_LOC_53/Y VSS 0.06fF
C78512 INVX1_LOC_64/Y VSS 0.62fF
C78513 NOR2X1_LOC_708/B VSS 0.19fF
C78514 NAND2X1_LOC_687/A VSS 0.19fF
C78515 NOR2X1_LOC_682/Y VSS 0.11fF
C78516 NOR2X1_LOC_681/Y VSS 0.20fF
C78517 NOR2X1_LOC_675/A VSS 0.09fF
C78518 NOR2X1_LOC_405/A VSS 0.54fF
C78519 INVX1_LOC_31/Y VSS 0.22fF
C78520 INVX1_LOC_20/Y VSS 0.44fF
C78521 GATE_662 VSS -0.03fF
C78522 NAND2X1_LOC_662/Y VSS 0.47fF
C78523 INVX1_LOC_268/Y VSS 0.28fF
C78524 INVX1_LOC_259/A VSS 0.26fF
C78525 NAND2X1_LOC_629/Y VSS 0.17fF
C78526 INVX1_LOC_257/Y VSS -0.08fF
C78527 NAND2X1_LOC_593/Y VSS 0.11fF
C78528 NAND2X1_LOC_650/B VSS 0.03fF
C78529 INVX1_LOC_126/A VSS 0.28fF
C78530 INVX1_LOC_100/A VSS 0.45fF
C78531 NOR2X1_LOC_199/B VSS 0.16fF
C78532 NAND2X1_LOC_41/Y VSS 0.23fF
C78533 INVX1_LOC_82/A VSS 0.19fF
C78534 INVX1_LOC_42/Y VSS 0.21fF
C78535 NOR2X1_LOC_160/Y VSS 0.11fF
C78536 NOR2X1_LOC_161/Y VSS -0.09fF
C78537 D_INPUT_2 VSS -0.91fF
C78538 NOR2X1_LOC_113/A VSS 0.25fF
C78539 NOR2X1_LOC_83/Y VSS 0.24fF
C78540 NOR2X1_LOC_71/Y VSS 0.85fF
C78541 NAND2X1_LOC_729/B VSS 0.54fF
C78542 NAND2X1_LOC_849/A VSS 0.48fF
C78543 NAND2X1_LOC_560/A VSS 0.25fF
C78544 NOR2X1_LOC_497/Y VSS 0.10fF
C78545 GATE_865 VSS 0.06fF
C78546 NOR2X1_LOC_495/Y VSS -0.23fF
C78547 INVX1_LOC_291/Y VSS 0.24fF
C78548 NAND2X1_LOC_807/Y VSS 0.31fF
C78549 NOR2X1_LOC_835/A VSS 0.28fF
C78550 NOR2X1_LOC_398/Y VSS 0.06fF
C78551 NOR2X1_LOC_387/Y VSS 0.17fF
C78552 NOR2X1_LOC_349/A VSS -0.80fF
C78553 NOR2X1_LOC_326/Y VSS 0.37fF
C78554 NOR2X1_LOC_367/B VSS 0.23fF
C78555 NOR2X1_LOC_364/Y VSS -0.02fF
C78556 NOR2X1_LOC_557/A VSS -0.60fF
C78557 NOR2X1_LOC_575/Y VSS 0.10fF
C78558 INVX1_LOC_232/A VSS -5.22fF
C78559 NOR2X1_LOC_566/Y VSS 0.09fF
C78560 NOR2X1_LOC_550/B VSS 0.36fF
C78561 NOR2X1_LOC_546/B VSS 0.28fF
C78562 NOR2X1_LOC_78/A VSS 0.92fF
C78563 NOR2X1_LOC_567/B VSS 0.38fF
C78564 NOR2X1_LOC_512/Y VSS 0.32fF
C78565 INVX1_LOC_199/Y VSS 0.02fF
C78566 INVX1_LOC_199/A VSS 0.32fF
C78567 INVX1_LOC_144/A VSS 0.44fF
C78568 INVX1_LOC_177/A VSS -0.91fF
C78569 INVX1_LOC_155/Y VSS 0.10fF
C78570 INVX1_LOC_155/A VSS 0.38fF
C78571 INVX1_LOC_111/A VSS 0.26fF
C78572 INVX1_LOC_100/Y VSS 0.15fF
C78573 INVX1_LOC_282/A VSS 0.16fF
C78574 INVX1_LOC_140/A VSS 1.15fF
C78575 NOR2X1_LOC_749/Y VSS 0.11fF
C78576 NOR2X1_LOC_731/Y VSS 0.07fF
C78577 NOR2X1_LOC_731/A VSS 0.23fF
C78578 NOR2X1_LOC_713/B VSS 0.47fF
C78579 NOR2X1_LOC_546/A VSS 0.13fF
C78580 INVX1_LOC_314/A VSS 0.09fF
C78581 INVX1_LOC_303/Y VSS 0.15fF
C78582 NAND2X1_LOC_477/A VSS 1.10fF
C78583 NAND2X1_LOC_466/Y VSS 0.29fF
C78584 INVX1_LOC_205/A VSS 0.18fF
C78585 INVX1_LOC_2/Y VSS -0.37fF
C78586 NOR2X1_LOC_7/Y VSS 0.15fF
C78587 INVX1_LOC_85/Y VSS 0.29fF
C78588 INVX1_LOC_52/A VSS 0.09fF
C78589 INVX1_LOC_96/Y VSS 0.28fF
C78590 INVX1_LOC_63/Y VSS 0.50fF
C78591 INVX1_LOC_41/Y VSS 0.69fF
C78592 INVX1_LOC_74/Y VSS 0.01fF
C78593 NAND2X1_LOC_654/B VSS 0.07fF
C78594 NAND2X1_LOC_638/Y VSS -0.20fF
C78595 NAND2X1_LOC_660/Y VSS 0.23fF
C78596 NOR2X1_LOC_672/Y VSS 0.12fF
C78597 NAND2X1_LOC_634/Y VSS -1.04fF
C78598 NAND2X1_LOC_633/Y VSS 0.13fF
C78599 INVX1_LOC_98/A VSS -0.79fF
C78600 NAND2X1_LOC_16/Y VSS 0.13fF
C78601 NAND2X1_LOC_39/Y VSS 0.19fF
C78602 NAND2X1_LOC_140/A VSS 0.52fF
C78603 NAND2X1_LOC_141/A VSS 0.54fF
C78604 INVX1_LOC_80/Y VSS -0.17fF
C78605 NOR2X1_LOC_554/B VSS 0.58fF
C78606 INVX1_LOC_36/Y VSS 0.27fF
C78607 INPUT_0 VSS -6.44fF
C78608 NOR2X1_LOC_123/B VSS 0.50fF
C78609 NOR2X1_LOC_423/Y VSS 0.55fF
C78610 NAND2X1_LOC_812/A VSS 0.24fF
C78611 NAND2X1_LOC_856/A VSS 0.07fF
C78612 NOR2X1_LOC_835/B VSS -0.04fF
C78613 NAND2X1_LOC_866/B VSS 0.16fF
C78614 NAND2X1_LOC_862/Y VSS 0.29fF
C78615 NAND2X1_LOC_861/Y VSS 0.07fF
C78616 INVX1_LOC_1/Y VSS 0.47fF
C78617 NOR2X1_LOC_82/Y VSS 0.21fF
C78618 NOR2X1_LOC_303/Y VSS 0.50fF
C78619 NOR2X1_LOC_357/Y VSS 0.08fF
C78620 NOR2X1_LOC_387/A VSS -1.17fF
C78621 NOR2X1_LOC_349/B VSS 0.32fF
C78622 NOR2X1_LOC_335/B VSS 0.28fF
C78623 NOR2X1_LOC_844/A VSS 0.51fF
C78624 NOR2X1_LOC_568/A VSS 0.31fF
C78625 NOR2X1_LOC_799/B VSS 0.27fF
C78626 INVX1_LOC_222/A VSS 0.36fF
C78627 INVX1_LOC_240/A VSS 0.85fF
C78628 INVX1_LOC_231/Y VSS 0.04fF
C78629 NOR2X1_LOC_577/Y VSS 0.48fF
C78630 NOR2X1_LOC_562/A VSS 0.12fF
C78631 NOR2X1_LOC_631/B VSS 0.22fF
C78632 NOR2X1_LOC_486/Y VSS -0.18fF
C78633 NOR2X1_LOC_589/Y VSS 0.10fF
C78634 NOR2X1_LOC_500/Y VSS -1.27fF
C78635 INVX1_LOC_121/Y VSS 0.25fF
C78636 INVX1_LOC_198/Y VSS 0.55fF
C78637 INVX1_LOC_187/Y VSS 0.11fF
C78638 INVX1_LOC_187/A VSS 0.35fF
C78639 INVX1_LOC_132/Y VSS 0.02fF
C78640 INVX1_LOC_165/Y VSS 0.15fF
C78641 INVX1_LOC_176/Y VSS 0.15fF
C78642 INVX1_LOC_110/A VSS 0.11fF
C78643 INVX1_LOC_154/A VSS 0.28fF
C78644 NOR2X1_LOC_112/Y VSS 0.34fF
C78645 NOR2X1_LOC_702/Y VSS 0.11fF
C78646 NOR2X1_LOC_748/Y VSS -0.09fF
C78647 NOR2X1_LOC_317/B VSS 0.48fF
C78648 NOR2X1_LOC_759/Y VSS 0.35fF
C78649 NOR2X1_LOC_209/A VSS 0.33fF
C78650 NOR2X1_LOC_711/Y VSS 0.12fF
C78651 NOR2X1_LOC_741/A VSS 0.09fF
C78652 NOR2X1_LOC_733/Y VSS 0.13fF
C78653 INVX1_LOC_285/Y VSS 0.62fF
C78654 INVX1_LOC_302/Y VSS 0.23fF
C78655 INVX1_LOC_302/A VSS 0.11fF
C78656 INVX1_LOC_313/Y VSS -6.71fF
C78657 INVX1_LOC_313/A VSS 0.35fF
C78658 GATE_479 VSS 0.08fF
C78659 NAND2X1_LOC_479/Y VSS 0.09fF
C78660 NOR2X1_LOC_493/B VSS 0.27fF
C78661 INVX1_LOC_95/Y VSS 0.68fF
C78662 INVX1_LOC_95/A VSS -0.08fF
C78663 INVX1_LOC_51/Y VSS 0.19fF
C78664 INVX1_LOC_62/A VSS 0.44fF
C78665 INVX1_LOC_40/A VSS 0.48fF
C78666 NOR2X1_LOC_707/B VSS 0.19fF
C78667 NAND2X1_LOC_662/B VSS 0.32fF
C78668 NOR2X1_LOC_686/B VSS 0.13fF
C78669 NAND2X1_LOC_640/Y VSS 0.39fF
C78670 NOR2X1_LOC_180/Y VSS 0.16fF
C78671 NOR2X1_LOC_181/Y VSS 0.13fF
C78672 NAND2X1_LOC_1/Y VSS 0.43fF
C78673 INVX1_LOC_86/Y VSS -0.39fF
C78674 INVX1_LOC_79/A VSS 0.51fF
C78675 NOR2X1_LOC_106/A VSS 0.66fF
C78676 INVX1_LOC_68/Y VSS 0.18fF
C78677 NAND2X1_LOC_841/A VSS 0.20fF
C78678 NAND2X1_LOC_866/A VSS 0.35fF
C78679 NAND2X1_LOC_863/Y VSS 0.23fF
C78680 INVX1_LOC_300/Y VSS 0.31fF
C78681 NAND2X1_LOC_850/A VSS 0.34fF
C78682 NAND2X1_LOC_819/Y VSS 0.11fF
C78683 NOR2X1_LOC_818/Y VSS -0.35fF
C78684 NOR2X1_LOC_350/A VSS -0.02fF
C78685 NOR2X1_LOC_396/Y VSS 0.04fF
C78686 NOR2X1_LOC_45/B VSS 0.84fF
C78687 NOR2X1_LOC_385/Y VSS 0.46fF
C78688 NOR2X1_LOC_359/Y VSS -0.03fF
C78689 NOR2X1_LOC_360/Y VSS -3.47fF
C78690 INVX1_LOC_96/A VSS 0.19fF
C78691 NOR2X1_LOC_337/Y VSS -0.31fF
C78692 INVX1_LOC_146/A VSS -0.11fF
C78693 NAND2X1_LOC_798/A VSS 0.49fF
C78694 INVX1_LOC_144/Y VSS -0.07fF
C78695 NOR2X1_LOC_522/Y VSS 0.17fF
C78696 INVX1_LOC_18/A VSS 1.07fF
C78697 INVX1_LOC_93/Y VSS 0.72fF
C78698 NOR2X1_LOC_569/Y VSS 0.23fF
C78699 NOR2X1_LOC_570/Y VSS 0.16fF
C78700 NOR2X1_LOC_551/B VSS 0.11fF
C78701 NOR2X1_LOC_374/A VSS 0.23fF
C78702 NOR2X1_LOC_599/A VSS -0.34fF
C78703 NOR2X1_LOC_562/B VSS 0.50fF
C78704 INVX1_LOC_206/Y VSS -0.14fF
C78705 INVX1_LOC_244/A VSS 0.21fF
C78706 INVX1_LOC_197/Y VSS 0.32fF
C78707 INVX1_LOC_197/A VSS -0.07fF
C78708 INVX1_LOC_153/Y VSS -2.41fF
C78709 INVX1_LOC_153/A VSS 0.12fF
C78710 INVX1_LOC_142/Y VSS 0.15fF
C78711 INVX1_LOC_142/A VSS 0.44fF
C78712 INVX1_LOC_186/A VSS -0.05fF
C78713 INVX1_LOC_131/A VSS -0.27fF
C78714 INVX1_LOC_164/A VSS 0.31fF
C78715 INVX1_LOC_120/Y VSS 0.15fF
C78716 NOR2X1_LOC_703/Y VSS 0.20fF
C78717 NOR2X1_LOC_704/Y VSS 0.11fF
C78718 NOR2X1_LOC_735/Y VSS 0.11fF
C78719 NOR2X1_LOC_732/A VSS 0.26fF
C78720 NOR2X1_LOC_712/Y VSS 0.12fF
C78721 INVX1_LOC_301/Y VSS 0.15fF
C78722 INVX1_LOC_312/A VSS 0.08fF
C78723 INVX1_LOC_83/Y VSS 0.15fF
C78724 INVX1_LOC_72/Y VSS 0.46fF
C78725 INVX1_LOC_72/A VSS 1.85fF
C78726 INVX1_LOC_61/Y VSS 0.45fF
C78727 NOR2X1_LOC_685/A VSS 0.39fF
C78728 NOR2X1_LOC_706/A VSS 0.64fF
C78729 NAND2X1_LOC_656/Y VSS 0.16fF
C78730 NAND2X1_LOC_672/B VSS -0.03fF
C78731 INVX1_LOC_104/A VSS 0.45fF
C78732 INVX1_LOC_94/A VSS -1.02fF
C78733 NOR2X1_LOC_168/Y VSS 0.16fF
C78734 NOR2X1_LOC_540/B VSS 0.36fF
C78735 NOR2X1_LOC_181/A VSS 0.12fF
C78736 NAND2X1_LOC_149/B VSS 0.11fF
C78737 NOR2X1_LOC_146/Y VSS 0.14fF
C78738 INVX1_LOC_67/A VSS 0.17fF
C78739 NOR2X1_LOC_106/Y VSS -0.05fF
C78740 INVX1_LOC_75/A VSS 1.41fF
C78741 NOR2X1_LOC_19/B VSS -3.77fF
C78742 NAND2X1_LOC_139/A VSS 0.36fF
C78743 NOR2X1_LOC_132/Y VSS 0.07fF
C78744 NOR2X1_LOC_91/Y VSS 0.28fF
C78745 INVX1_LOC_311/A VSS 0.76fF
C78746 NAND2X1_LOC_832/Y VSS 0.16fF
C78747 NAND2X1_LOC_842/B VSS 0.29fF
C78748 NAND2X1_LOC_839/Y VSS 0.11fF
C78749 NAND2X1_LOC_838/Y VSS 0.26fF
C78750 NOR2X1_LOC_384/Y VSS -1.66fF
C78751 INVX1_LOC_30/A VSS 2.44fF
C78752 NOR2X1_LOC_366/B VSS 0.22fF
C78753 INVX1_LOC_133/Y VSS 0.20fF
C78754 NOR2X1_LOC_361/Y VSS 0.18fF
C78755 NOR2X1_LOC_338/Y VSS 0.09fF
C78756 NOR2X1_LOC_355/B VSS 0.30fF
C78757 NAND2X1_LOC_308/B VSS 0.07fF
C78758 INVX1_LOC_143/A VSS 1.23fF
C78759 NOR2X1_LOC_316/Y VSS 0.05fF
C78760 NOR2X1_LOC_315/Y VSS 0.24fF
C78761 NOR2X1_LOC_588/A VSS -0.09fF
C78762 NOR2X1_LOC_52/B VSS 1.35fF
C78763 NOR2X1_LOC_552/A VSS -4.09fF
C78764 NOR2X1_LOC_318/B VSS -1.70fF
C78765 NOR2X1_LOC_569/A VSS 0.19fF
C78766 INVX1_LOC_174/Y VSS -0.18fF
C78767 INVX1_LOC_196/A VSS 0.30fF
C78768 INVX1_LOC_185/Y VSS 0.15fF
C78769 INVX1_LOC_130/Y VSS 0.24fF
C78770 INVX1_LOC_141/Y VSS 0.17fF
C78771 INVX1_LOC_141/A VSS 0.11fF
C78772 NOR2X1_LOC_772/A VSS 0.26fF
C78773 NOR2X1_LOC_137/A VSS 0.21fF
C78774 NOR2X1_LOC_757/Y VSS 0.18fF
C78775 NOR2X1_LOC_746/Y VSS 0.19fF
C78776 NAND2X1_LOC_45/Y VSS -0.40fF
C78777 NOR2X1_LOC_332/A VSS -4.70fF
C78778 NOR2X1_LOC_714/Y VSS 0.14fF
C78779 NOR2X1_LOC_725/A VSS 0.53fF
C78780 NOR2X1_LOC_706/Y VSS 0.09fF
C78781 INVX1_LOC_311/Y VSS 0.20fF
C78782 INVX1_LOC_300/A VSS 0.11fF
C78783 NOR2X1_LOC_6/B VSS 1.10fF
C78784 INVX1_LOC_60/Y VSS 0.42fF
C78785 INVX1_LOC_60/A VSS -0.22fF
C78786 NOR2X1_LOC_192/A VSS -0.12fF
C78787 NOR2X1_LOC_439/B VSS 0.39fF
C78788 NOR2X1_LOC_210/B VSS 0.01fF
C78789 INVX1_LOC_85/A VSS 0.89fF
C78790 NOR2X1_LOC_144/Y VSS 0.11fF
C78791 NOR2X1_LOC_142/Y VSS 0.84fF
C78792 NOR2X1_LOC_514/A VSS 0.68fF
C78793 INVX1_LOC_31/A VSS 0.77fF
C78794 NOR2X1_LOC_113/B VSS 0.25fF
C78795 NOR2X1_LOC_128/B VSS 0.34fF
C78796 NAND2X1_LOC_116/A VSS 0.54fF
C78797 INVX1_LOC_39/Y VSS 0.28fF
C78798 NAND2X1_LOC_858/B VSS -0.47fF
C78799 NAND2X1_LOC_840/Y VSS 0.11fF
C78800 NAND2X1_LOC_859/Y VSS 0.79fF
C78801 NAND2X1_LOC_833/Y VSS 0.78fF
C78802 NOR2X1_LOC_372/Y VSS 0.10fF
C78803 INVX1_LOC_158/A VSS 0.25fF
C78804 NOR2X1_LOC_340/Y VSS 0.17fF
C78805 NOR2X1_LOC_276/Y VSS -0.03fF
C78806 NAND2X1_LOC_51/B VSS 0.48fF
C78807 D_INPUT_4 VSS -1.16fF
C78808 NAND2X1_LOC_319/A VSS -0.36fF
C78809 INVX1_LOC_151/A VSS 0.12fF
C78810 NAND2X1_LOC_332/Y VSS 0.01fF
C78811 NOR2X1_LOC_573/Y VSS 0.11fF
C78812 NOR2X1_LOC_551/Y VSS 0.07fF
C78813 NOR2X1_LOC_552/Y VSS -0.17fF
C78814 NOR2X1_LOC_597/Y VSS 0.24fF
C78815 NOR2X1_LOC_597/A VSS -0.04fF
C78816 INVX1_LOC_218/A VSS 0.02fF
C78817 NOR2X1_LOC_520/A VSS -0.10fF
C78818 NOR2X1_LOC_541/Y VSS 0.38fF
C78819 INVX1_LOC_140/Y VSS 0.24fF
C78820 INVX1_LOC_173/Y VSS 0.40fF
C78821 INVX1_LOC_151/Y VSS 0.15fF
C78822 INVX1_LOC_162/Y VSS 0.29fF
C78823 INVX1_LOC_162/A VSS 0.09fF
C78824 INVX1_LOC_184/Y VSS 0.15fF
C78825 INVX1_LOC_184/A VSS 0.09fF
C78826 INVX1_LOC_195/Y VSS 0.15fF
C78827 INVX1_LOC_195/A VSS -0.07fF
C78828 INVX1_LOC_211/A VSS 0.24fF
C78829 NOR2X1_LOC_503/Y VSS -0.69fF
C78830 NAND2X1_LOC_227/Y VSS 0.35fF
C78831 INVX1_LOC_286/A VSS 0.17fF
C78832 NOR2X1_LOC_721/Y VSS 0.05fF
C78833 NOR2X1_LOC_756/Y VSS -0.18fF
C78834 NOR2X1_LOC_789/A VSS 0.28fF
C78835 NOR2X1_LOC_717/Y VSS 0.02fF
C78836 NOR2X1_LOC_745/Y VSS 0.07fF
C78837 NOR2X1_LOC_708/Y VSS 0.24fF
C78838 NOR2X1_LOC_701/Y VSS 0.06fF
C78839 INVX1_LOC_310/Y VSS 0.57fF
C78840 INVX1_LOC_81/Y VSS 0.31fF
C78841 INVX1_LOC_70/Y VSS 0.16fF
C78842 INVX1_LOC_92/Y VSS 0.41fF
C78843 NOR2X1_LOC_690/Y VSS 0.17fF
C78844 NOR2X1_LOC_191/A VSS 0.26fF
C78845 INVX1_LOC_98/Y VSS 0.23fF
C78846 NOR2X1_LOC_148/A VSS 0.12fF
C78847 INVX1_LOC_73/A VSS 0.63fF
C78848 NAND2X1_LOC_123/Y VSS 0.20fF
C78849 NOR2X1_LOC_122/Y VSS 0.14fF
C78850 NAND2X1_LOC_170/A VSS 0.34fF
C78851 NOR2X1_LOC_165/Y VSS 0.08fF
C78852 INVX1_LOC_77/A VSS 0.71fF
C78853 NAND2X1_LOC_114/B VSS 0.37fF
C78854 NOR2X1_LOC_107/Y VSS 0.07fF
C78855 NOR2X1_LOC_103/Y VSS 0.96fF
C78856 NAND2X1_LOC_860/Y VSS 0.11fF
C78857 INVX1_LOC_256/Y VSS 0.22fF
C78858 INVX1_LOC_314/Y VSS 0.46fF
C78859 NOR2X1_LOC_372/A VSS -0.36fF
C78860 INVX1_LOC_28/A VSS -6.51fF
C78861 NOR2X1_LOC_860/B VSS 0.16fF
C78862 NOR2X1_LOC_307/A VSS 0.05fF
C78863 NOR2X1_LOC_329/B VSS 0.81fF
C78864 NAND2X1_LOC_342/Y VSS 0.38fF
C78865 NAND2X1_LOC_351/A VSS 0.33fF
C78866 NOR2X1_LOC_530/Y VSS 0.18fF
C78867 NOR2X1_LOC_542/Y VSS 0.06fF
C78868 NOR2X1_LOC_570/A VSS 0.09fF
C78869 NOR2X1_LOC_553/Y VSS 0.08fF
C78870 INVX1_LOC_236/A VSS 0.16fF
C78871 NOR2X1_LOC_574/A VSS 0.42fF
C78872 NOR2X1_LOC_596/A VSS 0.98fF
C78873 INVX1_LOC_161/Y VSS 0.43fF
C78874 INVX1_LOC_183/Y VSS 0.25fF
C78875 INVX1_LOC_172/Y VSS 0.34fF
C78876 NAND2X1_LOC_510/A VSS 0.19fF
C78877 INVX1_LOC_210/Y VSS 0.29fF
C78878 NOR2X1_LOC_700/Y VSS -0.09fF
C78879 NOR2X1_LOC_802/A VSS 0.50fF
C78880 NOR2X1_LOC_593/Y VSS 0.94fF
C78881 NOR2X1_LOC_744/Y VSS 0.11fF
C78882 NOR2X1_LOC_794/A VSS 0.11fF
C78883 NOR2X1_LOC_784/B VSS 0.04fF
C78884 NOR2X1_LOC_718/Y VSS 0.13fF
C78885 INVX1_LOC_283/Y VSS 0.22fF
C78886 NOR2X1_LOC_722/Y VSS 0.17fF
C78887 NOR2X1_LOC_723/Y VSS 0.24fF
C78888 INVX1_LOC_91/Y VSS 0.15fF
C78889 INVX1_LOC_80/A VSS 0.18fF
C78890 NAND2X1_LOC_154/Y VSS 0.19fF
C78891 NOR2X1_LOC_148/B VSS 0.30fF
C78892 NOR2X1_LOC_703/B VSS 0.67fF
C78893 INVX1_LOC_69/Y VSS 0.21fF
C78894 NAND2X1_LOC_656/A VSS 0.90fF
C78895 INVX1_LOC_62/Y VSS 0.10fF
C78896 NOR2X1_LOC_391/Y VSS 0.27fF
C78897 NOR2X1_LOC_543/A VSS 0.22fF
C78898 NOR2X1_LOC_307/B VSS 0.18fF
C78899 NAND2X1_LOC_354/B VSS -0.17fF
C78900 NAND2X1_LOC_325/Y VSS -0.16fF
C78901 NAND2X1_LOC_352/B VSS 0.11fF
C78902 INVX1_LOC_150/Y VSS -1.43fF
C78903 NAND2X1_LOC_359/A VSS 0.24fF
C78904 INVX1_LOC_154/Y VSS 0.31fF
C78905 INVX1_LOC_156/Y VSS 0.06fF
C78906 NOR2X1_LOC_474/A VSS 0.44fF
C78907 NOR2X1_LOC_250/A VSS 0.34fF
C78908 NOR2X1_LOC_553/B VSS 0.08fF
C78909 NOR2X1_LOC_570/B VSS 0.09fF
C78910 INVX1_LOC_193/Y VSS 0.28fF
C78911 INVX1_LOC_182/Y VSS 0.19fF
C78912 INVX1_LOC_182/A VSS 0.08fF
C78913 INVX1_LOC_171/A VSS 0.34fF
C78914 INVX1_LOC_160/Y VSS 0.40fF
C78915 INVX1_LOC_209/A VSS 0.12fF
C78916 NOR2X1_LOC_504/Y VSS 0.21fF
C78917 NOR2X1_LOC_520/B VSS 0.36fF
C78918 INVX1_LOC_49/A VSS 1.00fF
C78919 NOR2X1_LOC_354/B VSS -0.14fF
C78920 NOR2X1_LOC_785/A VSS 0.30fF
C78921 NOR2X1_LOC_241/A VSS 0.22fF
C78922 NOR2X1_LOC_433/A VSS 0.98fF
C78923 NOR2X1_LOC_794/B VSS -0.19fF
C78924 NOR2X1_LOC_457/A VSS 0.37fF
C78925 NOR2X1_LOC_711/A VSS -0.07fF
C78926 NOR2X1_LOC_738/A VSS 0.17fF
C78927 NOR2X1_LOC_724/Y VSS -0.23fF
C78928 INVX1_LOC_107/A VSS 0.12fF
C78929 NAND2X1_LOC_195/Y VSS 0.19fF
C78930 NOR2X1_LOC_816/A VSS 0.48fF
C78931 NOR2X1_LOC_147/A VSS 0.03fF
C78932 NAND2X1_LOC_156/B VSS 0.03fF
C78933 NOR2X1_LOC_169/B VSS 0.07fF
C78934 NOR2X1_LOC_124/B VSS 0.31fF
C78935 NOR2X1_LOC_121/Y VSS 0.11fF
C78936 INVX1_LOC_33/A VSS 0.90fF
C78937 INVX1_LOC_61/A VSS 0.81fF
C78938 NOR2X1_LOC_86/Y VSS 0.07fF
C78939 NOR2X1_LOC_391/B VSS -0.14fF
C78940 NAND2X1_LOC_360/B VSS 0.38fF
C78941 NOR2X1_LOC_317/A VSS 0.12fF
C78942 NAND2X1_LOC_337/B VSS 0.19fF
C78943 NOR2X1_LOC_323/Y VSS 0.08fF
C78944 NOR2X1_LOC_322/Y VSS 0.59fF
C78945 INVX1_LOC_234/A VSS 0.69fF
C78946 NOR2X1_LOC_557/Y VSS 0.38fF
C78947 NOR2X1_LOC_565/A VSS 0.09fF
C78948 INVX1_LOC_225/Y VSS -0.82fF
C78949 NOR2X1_LOC_594/Y VSS 0.39fF
C78950 INVX1_LOC_192/A VSS 0.29fF
C78951 INVX1_LOC_181/Y VSS 0.52fF
C78952 NAND2X1_LOC_799/A VSS 0.41fF
C78953 NAND2X1_LOC_538/Y VSS 0.07fF
C78954 NAND2X1_LOC_537/Y VSS -1.53fF
C78955 NAND2X1_LOC_508/A VSS 0.62fF
C78956 INVX1_LOC_120/A VSS 0.58fF
C78957 NOR2X1_LOC_620/B VSS 0.37fF
C78958 NOR2X1_LOC_559/B VSS 0.36fF
C78959 INVX1_LOC_170/A VSS 0.25fF
C78960 NOR2X1_LOC_97/A VSS 0.46fF
C78961 NOR2X1_LOC_112/B VSS 0.03fF
C78962 NOR2X1_LOC_803/A VSS 0.19fF
C78963 NOR2X1_LOC_721/A VSS 0.11fF
C78964 NOR2X1_LOC_753/Y VSS 0.34fF
C78965 NOR2X1_LOC_726/Y VSS 0.17fF
C78966 D_GATE_741 VSS 0.07fF
C78967 NOR2X1_LOC_740/Y VSS -0.45fF
C78968 NOR2X1_LOC_215/Y VSS 0.07fF
C78969 NOR2X1_LOC_180/B VSS 0.77fF
C78970 NOR2X1_LOC_168/A VSS 0.12fF
C78971 NOR2X1_LOC_191/B VSS 0.15fF
C78972 NAND2X1_LOC_208/B VSS -0.62fF
C78973 INVX1_LOC_43/Y VSS 0.02fF
C78974 NOR2X1_LOC_122/A VSS 0.21fF
C78975 NOR2X1_LOC_666/A VSS 0.58fF
C78976 INVX1_LOC_83/A VSS -13.69fF
C78977 INVX1_LOC_7/A VSS 0.65fF
C78978 NAND2X1_LOC_323/B VSS -0.45fF
C78979 NOR2X1_LOC_392/B VSS -4.35fF
C78980 NOR2X1_LOC_388/Y VSS 0.12fF
C78981 NOR2X1_LOC_457/B VSS 0.94fF
C78982 NOR2X1_LOC_270/Y VSS -0.21fF
C78983 NAND2X1_LOC_326/A VSS 0.28fF
C78984 NOR2X1_LOC_321/Y VSS 0.12fF
C78985 NOR2X1_LOC_320/Y VSS 0.07fF
C78986 NOR2X1_LOC_380/A VSS -0.07fF
C78987 INVX1_LOC_149/A VSS 0.67fF
C78988 NOR2X1_LOC_310/Y VSS 0.06fF
C78989 NOR2X1_LOC_309/Y VSS 0.44fF
C78990 NAND2X1_LOC_364/A VSS 0.53fF
C78991 NAND2X1_LOC_347/B VSS 0.40fF
C78992 NOR2X1_LOC_292/Y VSS 0.14fF
C78993 NAND2X1_LOC_303/B VSS 0.21fF
C78994 NOR2X1_LOC_299/Y VSS 0.37fF
C78995 NOR2X1_LOC_298/Y VSS 1.27fF
C78996 NOR2X1_LOC_718/B VSS 0.34fF
C78997 NOR2X1_LOC_582/Y VSS 0.18fF
C78998 NOR2X1_LOC_576/B VSS 0.65fF
C78999 INVX1_LOC_229/Y VSS -3.37fF
C79000 NOR2X1_LOC_561/Y VSS 0.30fF
C79001 INVX1_LOC_191/Y VSS 0.32fF
C79002 INVX1_LOC_180/A VSS -0.04fF
C79003 INVX1_LOC_215/Y VSS 0.18fF
C79004 NOR2X1_LOC_513/Y VSS 0.07fF
C79005 NOR2X1_LOC_507/A VSS 0.29fF
C79006 NOR2X1_LOC_775/Y VSS -0.20fF
C79007 INVX1_LOC_297/Y VSS -0.06fF
C79008 NOR2X1_LOC_773/Y VSS 0.16fF
C79009 NOR2X1_LOC_803/B VSS 0.32fF
C79010 NOR2X1_LOC_784/Y VSS 0.33fF
C79011 NOR2X1_LOC_742/A VSS 0.42fF
C79012 NOR2X1_LOC_736/Y VSS 0.03fF
C79013 INVX1_LOC_290/A VSS -3.47fF
C79014 NOR2X1_LOC_666/Y VSS -0.34fF
C79015 NOR2X1_LOC_216/Y VSS 0.36fF
C79016 NOR2X1_LOC_214/B VSS 0.26fF
C79017 NOR2X1_LOC_229/Y VSS 0.19fF
C79018 NOR2X1_LOC_147/B VSS -0.45fF
C79019 NAND2X1_LOC_198/B VSS 0.65fF
C79020 NOR2X1_LOC_52/Y VSS 0.12fF
C79021 NOR2X1_LOC_173/Y VSS 0.12fF
C79022 NOR2X1_LOC_168/B VSS 0.32fF
C79023 NOR2X1_LOC_140/A VSS 0.16fF
C79024 INVX1_LOC_121/A VSS 0.40fF
C79025 NOR2X1_LOC_300/Y VSS 0.09fF
C79026 INVX1_LOC_159/A VSS -0.58fF
C79027 NAND2X1_LOC_355/Y VSS 0.13fF
C79028 NAND2X1_LOC_354/Y VSS 0.50fF
C79029 INVX1_LOC_161/A VSS 0.33fF
C79030 NOR2X1_LOC_459/A VSS -0.00fF
C79031 NAND2X1_LOC_377/Y VSS 0.20fF
C79032 NAND2X1_LOC_338/B VSS 1.00fF
C79033 NOR2X1_LOC_290/Y VSS 0.24fF
C79034 GATE_366 VSS 0.02fF
C79035 INVX1_LOC_246/A VSS -0.34fF
C79036 NOR2X1_LOC_592/A VSS 0.12fF
C79037 NOR2X1_LOC_582/A VSS 0.01fF
C79038 D_INPUT_6 VSS 0.28fF
C79039 NOR2X1_LOC_2/Y VSS -0.03fF
C79040 INVX1_LOC_190/Y VSS 0.31fF
C79041 INVX1_LOC_190/A VSS 0.11fF
C79042 NAND2X1_LOC_514/Y VSS 0.13fF
C79043 INVX1_LOC_177/Y VSS 0.24fF
C79044 NOR2X1_LOC_536/Y VSS 0.11fF
C79045 NOR2X1_LOC_507/B VSS 0.13fF
C79046 INVX1_LOC_89/A VSS 1.30fF
C79047 NAND2X1_LOC_549/B VSS 0.11fF
C79048 NOR2X1_LOC_529/Y VSS 0.05fF
C79049 INVX1_LOC_217/A VSS -3.42fF
C79050 NOR2X1_LOC_517/Y VSS 0.07fF
C79051 NOR2X1_LOC_751/A VSS 0.37fF
C79052 NOR2X1_LOC_785/Y VSS 0.24fF
C79053 INVX1_LOC_294/Y VSS -0.10fF
C79054 NOR2X1_LOC_772/Y VSS 0.23fF
C79055 NOR2X1_LOC_778/Y VSS 0.23fF
C79056 NOR2X1_LOC_738/Y VSS 0.07fF
C79057 NOR2X1_LOC_739/Y VSS 0.30fF
C79058 NOR2X1_LOC_763/A VSS -0.36fF
C79059 NAND2X1_LOC_712/A VSS 0.17fF
C79060 NOR2X1_LOC_695/Y VSS 0.11fF
C79061 NAND2X1_LOC_722/A VSS 0.29fF
C79062 NOR2X1_LOC_716/B VSS 0.28fF
C79063 NAND2X1_LOC_7/Y VSS 0.28fF
C79064 NOR2X1_LOC_218/A VSS 0.39fF
C79065 INVX1_LOC_73/Y VSS 0.15fF
C79066 NOR2X1_LOC_215/A VSS 0.20fF
C79067 NOR2X1_LOC_202/Y VSS 0.10fF
C79068 NOR2X1_LOC_162/Y VSS 0.10fF
C79069 NAND2X1_LOC_199/B VSS 0.25fF
C79070 NOR2X1_LOC_45/Y VSS 0.31fF
C79071 NOR2X1_LOC_151/Y VSS -1.99fF
C79072 NOR2X1_LOC_589/A VSS -2.42fF
C79073 NAND2X1_LOC_175/B VSS 0.30fF
C79074 NOR2X1_LOC_172/Y VSS -0.25fF
C79075 INVX1_LOC_82/Y VSS 0.12fF
C79076 NAND2X1_LOC_390/A VSS 0.43fF
C79077 NOR2X1_LOC_331/Y VSS -0.28fF
C79078 INVX1_LOC_147/A VSS -0.03fF
C79079 NOR2X1_LOC_289/Y VSS 0.11fF
C79080 NOR2X1_LOC_171/Y VSS 0.13fF
C79081 NOR2X1_LOC_336/B VSS 0.23fF
C79082 INVX1_LOC_14/A VSS 0.86fF
C79083 INVX1_LOC_1/A VSS -13.72fF
C79084 NAND2X1_LOC_348/A VSS 0.70fF
C79085 NOR2X1_LOC_256/Y VSS 0.06fF
C79086 NAND2X1_LOC_367/B VSS 0.23fF
C79087 NAND2X1_LOC_363/Y VSS 0.14fF
C79088 D_GATE_579 VSS -0.00fF
C79089 INVX1_LOC_239/Y VSS -0.07fF
C79090 NOR2X1_LOC_591/Y VSS 0.11fF
C79091 NAND2X1_LOC_577/A VSS 0.58fF
C79092 NAND2X1_LOC_561/B VSS 0.31fF
C79093 NOR2X1_LOC_494/Y VSS 0.11fF
C79094 NAND2X1_LOC_493/Y VSS 0.35fF
C79095 NOR2X1_LOC_136/Y VSS 0.16fF
C79096 NOR2X1_LOC_537/A VSS 0.16fF
C79097 NOR2X1_LOC_502/Y VSS 0.08fF
C79098 NOR2X1_LOC_804/B VSS 0.39fF
C79099 NOR2X1_LOC_761/Y VSS 0.16fF
C79100 NOR2X1_LOC_599/Y VSS 0.29fF
C79101 NOR2X1_LOC_796/B VSS 0.17fF
C79102 NOR2X1_LOC_779/Y VSS 0.07fF
C79103 NAND2X1_LOC_740/B VSS 0.19fF
C79104 INVX1_LOC_273/Y VSS 0.06fF
C79105 NAND2X1_LOC_374/Y VSS 0.79fF
C79106 NOR2X1_LOC_238/Y VSS 0.25fF
C79107 NOR2X1_LOC_160/B VSS 1.64fF
C79108 NOR2X1_LOC_227/B VSS 0.13fF
C79109 NOR2X1_LOC_473/B VSS -0.99fF
C79110 NOR2X1_LOC_203/Y VSS 0.12fF
C79111 INVX1_LOC_111/Y VSS 0.49fF
C79112 NOR2X1_LOC_419/Y VSS 0.35fF
C79113 INVX1_LOC_24/A VSS 1.79fF
C79114 INVX1_LOC_174/A VSS 2.15fF
C79115 NOR2X1_LOC_41/Y VSS 0.07fF
C79116 INVX1_LOC_81/A VSS 0.38fF
C79117 INVX1_LOC_88/A VSS 0.76fF
C79118 NOR2X1_LOC_175/B VSS 0.56fF
C79119 INVX1_LOC_54/Y VSS -1.36fF
C79120 INVX1_LOC_209/Y VSS 0.41fF
C79121 NOR2X1_LOC_389/A VSS 0.93fF
C79122 INVX1_LOC_135/Y VSS 0.31fF
C79123 NOR2X1_LOC_375/Y VSS 0.08fF
C79124 INVX1_LOC_84/Y VSS -0.07fF
C79125 NAND2X1_LOC_367/A VSS 0.23fF
C79126 NAND2X1_LOC_364/Y VSS 0.42fF
C79127 NOR2X1_LOC_135/Y VSS 0.37fF
C79128 NOR2X1_LOC_111/Y VSS 0.18fF
C79129 NAND2X1_LOC_349/B VSS -0.85fF
C79130 NOR2X1_LOC_251/Y VSS -0.01fF
C79131 NOR2X1_LOC_335/A VSS 0.27fF
C79132 NOR2X1_LOC_590/Y VSS 0.14fF
C79133 NOR2X1_LOC_516/B VSS 0.76fF
C79134 NAND2X1_LOC_567/Y VSS 0.22fF
C79135 INVX1_LOC_221/Y VSS -0.06fF
C79136 NOR2X1_LOC_533/Y VSS 0.26fF
C79137 NOR2X1_LOC_490/Y VSS 0.12fF
C79138 INVX1_LOC_241/A VSS 0.31fF
C79139 NOR2X1_LOC_545/A VSS 0.12fF
C79140 NAND2X1_LOC_550/A VSS 1.00fF
C79141 NOR2X1_LOC_503/A VSS 0.12fF
C79142 INVX1_LOC_305/Y VSS 0.14fF
C79143 NOR2X1_LOC_781/Y VSS 0.25fF
C79144 INVX1_LOC_292/A VSS 0.73fF
C79145 INVX1_LOC_298/A VSS 0.18fF
C79146 NOR2X1_LOC_770/Y VSS 0.17fF
C79147 NAND2X1_LOC_740/A VSS -0.12fF
C79148 NAND2X1_LOC_731/Y VSS -0.23fF
C79149 NOR2X1_LOC_750/A VSS -0.07fF
C79150 NOR2X1_LOC_526/Y VSS -0.09fF
C79151 NOR2X1_LOC_237/Y VSS 0.38fF
C79152 NAND2X1_LOC_79/Y VSS 0.22fF
C79153 NOR2X1_LOC_205/Y VSS 0.23fF
C79154 NOR2X1_LOC_828/B VSS -0.22fF
C79155 NOR2X1_LOC_418/Y VSS 0.35fF
C79156 NOR2X1_LOC_430/A VSS 0.12fF
C79157 NOR2X1_LOC_174/A VSS 0.32fF
C79158 NAND2X1_LOC_200/B VSS 0.30fF
C79159 NOR2X1_LOC_16/Y VSS 0.17fF
C79160 NAND2X1_LOC_162/B VSS 0.11fF
C79161 NAND2X1_LOC_20/B VSS 0.32fF
C79162 INVX1_LOC_47/A VSS 0.20fF
C79163 INVX1_LOC_208/Y VSS 0.29fF
C79164 INVX1_LOC_208/A VSS -3.24fF
C79165 INVX1_LOC_219/Y VSS 0.25fF
C79166 NAND2X1_LOC_387/B VSS 0.11fF
C79167 NAND2X1_LOC_36/A VSS -1.59fF
C79168 NOR2X1_LOC_376/A VSS 0.27fF
C79169 NOR2X1_LOC_355/A VSS -2.39fF
C79170 INVX1_LOC_145/Y VSS -0.06fF
C79171 NAND2X1_LOC_357/B VSS 0.35fF
C79172 NAND2X1_LOC_308/Y VSS 0.46fF
C79173 NOR2X1_LOC_248/Y VSS 0.14fF
C79174 INVX1_LOC_163/A VSS 0.40fF
C79175 NAND2X1_LOC_358/Y VSS 0.22fF
C79176 NAND2X1_LOC_513/B VSS 0.11fF
C79177 NAND2X1_LOC_854/B VSS 0.39fF
C79178 INVX1_LOC_221/A VSS 0.30fF
C79179 INVX1_LOC_223/A VSS -0.53fF
C79180 NOR2X1_LOC_524/Y VSS 0.10fF
C79181 NOR2X1_LOC_441/Y VSS 0.77fF
C79182 INVX1_LOC_239/A VSS -2.19fF
C79183 NOR2X1_LOC_521/Y VSS 0.30fF
C79184 NAND2X1_LOC_562/B VSS 0.32fF
C79185 NAND2X1_LOC_483/Y VSS 0.24fF
C79186 NAND2X1_LOC_500/Y VSS 0.07fF
C79187 NOR2X1_LOC_791/Y VSS -0.46fF
C79188 NOR2X1_LOC_781/B VSS 0.29fF
C79189 NOR2X1_LOC_781/A VSS 0.39fF
C79190 NOR2X1_LOC_770/B VSS 0.31fF
C79191 NAND2X1_LOC_741/B VSS 0.25fF
C79192 INVX1_LOC_286/Y VSS -3.08fF
C79193 NAND2X1_LOC_733/Y VSS 0.96fF
C79194 NAND2X1_LOC_714/B VSS 0.42fF
C79195 INVX1_LOC_178/A VSS 1.75fF
C79196 INVX1_LOC_279/A VSS -3.79fF
C79197 NAND2X1_LOC_112/Y VSS -0.22fF
C79198 NOR2X1_LOC_792/B VSS 0.28fF
C79199 NOR2X1_LOC_758/Y VSS -0.02fF
C79200 NAND2X1_LOC_711/Y VSS 0.21fF
C79201 NOR2X1_LOC_789/B VSS 0.13fF
C79202 NAND2X1_LOC_72/Y VSS 0.23fF
C79203 INVX1_LOC_55/Y VSS 0.03fF
C79204 NOR2X1_LOC_219/B VSS -0.04fF
C79205 NOR2X1_LOC_208/Y VSS -2.31fF
C79206 NOR2X1_LOC_544/A VSS -0.13fF
C79207 NOR2X1_LOC_428/Y VSS -0.37fF
C79208 NAND2X1_LOC_162/A VSS 0.12fF
C79209 INVX1_LOC_105/A VSS 0.52fF
C79210 NOR2X1_LOC_13/Y VSS 0.50fF
C79211 NAND2X1_LOC_181/Y VSS 0.06fF
C79212 INVX1_LOC_45/Y VSS 0.55fF
C79213 NOR2X1_LOC_609/A VSS 0.25fF
C79214 INVX1_LOC_218/Y VSS 0.42fF
C79215 INVX1_LOC_207/Y VSS 0.24fF
C79216 NAND2X1_LOC_350/B VSS 0.18fF
C79217 NAND2X1_LOC_231/Y VSS -4.85fF
C79218 INVX1_LOC_145/A VSS 0.21fF
C79219 NAND2X1_LOC_357/A VSS 0.06fF
C79220 NOR2X1_LOC_389/B VSS 0.19fF
C79221 NAND2X1_LOC_359/Y VSS 0.38fF
C79222 NOR2X1_LOC_401/A VSS 0.22fF
C79223 NOR2X1_LOC_644/A VSS 0.25fF
C79224 NOR2X1_LOC_828/A VSS 0.64fF
C79225 INVX1_LOC_243/A VSS 0.39fF
C79226 NAND2X1_LOC_568/A VSS 0.21fF
C79227 NAND2X1_LOC_303/Y VSS 0.79fF
C79228 NOR2X1_LOC_788/B VSS 0.39fF
C79229 NOR2X1_LOC_532/Y VSS 0.11fF
C79230 NAND2X1_LOC_578/B VSS 0.11fF
C79231 NAND2X1_LOC_570/Y VSS 0.13fF
C79232 INVX1_LOC_122/Y VSS -1.25fF
C79233 NOR2X1_LOC_523/A VSS -0.00fF
C79234 NAND2X1_LOC_551/A VSS 0.49fF
C79235 NOR2X1_LOC_373/Y VSS -0.11fF
C79236 NOR2X1_LOC_791/B VSS -0.33fF
C79237 NOR2X1_LOC_791/A VSS 0.03fF
C79238 NOR2X1_LOC_783/A VSS 0.24fF
C79239 NOR2X1_LOC_780/B VSS 0.48fF
C79240 INVX1_LOC_295/A VSS 0.77fF
C79241 NOR2X1_LOC_764/Y VSS 0.06fF
C79242 NOR2X1_LOC_763/Y VSS 0.63fF
C79243 NOR2X1_LOC_759/A VSS 0.10fF
C79244 NAND2X1_LOC_724/A VSS 0.26fF
C79245 NAND2X1_LOC_703/Y VSS 0.24fF
C79246 NOR2X1_LOC_312/Y VSS -1.08fF
C79247 NOR2X1_LOC_246/Y VSS 0.13fF
C79248 NAND2X1_LOC_67/Y VSS 0.07fF
C79249 INVX1_LOC_52/Y VSS 0.12fF
C79250 NOR2X1_LOC_224/Y VSS -0.20fF
C79251 NOR2X1_LOC_220/A VSS 0.79fF
C79252 NOR2X1_LOC_209/Y VSS -1.19fF
C79253 INVX1_LOC_90/A VSS -4.38fF
C79254 NOR2X1_LOC_78/B VSS 0.74fF
C79255 INVX1_LOC_103/A VSS 0.39fF
C79256 INVX1_LOC_101/Y VSS 0.17fF
C79257 INVX1_LOC_93/A VSS 0.80fF
C79258 NAND2X1_LOC_169/Y VSS 0.28fF
C79259 D_INPUT_0 VSS 0.86fF
C79260 INVX1_LOC_206/A VSS 0.41fF
C79261 INVX1_LOC_217/Y VSS 0.20fF
C79262 INVX1_LOC_228/A VSS 0.30fF
C79263 NAND2X1_LOC_350/A VSS 0.65fF
C79264 NAND2X1_LOC_358/B VSS 0.11fF
C79265 INVX1_LOC_152/Y VSS 0.32fF
C79266 NOR2X1_LOC_391/A VSS 0.23fF
C79267 NOR2X1_LOC_383/Y VSS 0.34fF
C79268 INVX1_LOC_30/Y VSS 0.36fF
C79269 NAND2X1_LOC_366/A VSS 0.23fF
C79270 NAND2X1_LOC_361/Y VSS 0.45fF
C79271 NAND2X1_LOC_588/B VSS 0.34fF
C79272 D_INPUT_7 VSS 0.05fF
C79273 INVX1_LOC_237/A VSS 0.09fF
C79274 INVX1_LOC_234/Y VSS 0.31fF
C79275 NAND2X1_LOC_571/Y VSS -0.04fF
C79276 NAND2X1_LOC_569/B VSS 0.53fF
C79277 NAND2X1_LOC_549/Y VSS 0.27fF
C79278 INVX1_LOC_227/A VSS 0.54fF
C79279 NOR2X1_LOC_533/A VSS 0.17fF
C79280 INVX1_LOC_212/Y VSS 0.31fF
C79281 NOR2X1_LOC_523/B VSS 0.13fF
C79282 NOR2X1_LOC_68/A VSS 1.45fF
C79283 NOR2X1_LOC_369/Y VSS 0.17fF
C79284 NOR2X1_LOC_793/A VSS 0.01fF
C79285 NOR2X1_LOC_790/A VSS 0.12fF
C79286 NAND2X1_LOC_783/A VSS -1.06fF
C79287 INVX1_LOC_280/Y VSS 0.34fF
C79288 NAND2X1_LOC_736/B VSS 0.10fF
C79289 INVX1_LOC_207/A VSS 0.19fF
C79290 NOR2X1_LOC_134/Y VSS 0.22fF
C79291 NAND2X1_LOC_725/B VSS 0.27fF
C79292 NAND2X1_LOC_706/Y VSS 0.23fF
C79293 NAND2X1_LOC_705/Y VSS 0.19fF
C79294 NAND2X1_LOC_715/B VSS 0.22fF
C79295 NOR2X1_LOC_234/Y VSS 0.14fF
C79296 NOR2X1_LOC_361/B VSS 0.87fF
C79297 NOR2X1_LOC_220/B VSS 0.17fF
C79298 NOR2X1_LOC_211/Y VSS 0.09fF
C79299 NOR2X1_LOC_246/A VSS -0.94fF
C79300 D_GATE_222 VSS -0.07fF
C79301 NOR2X1_LOC_222/Y VSS 0.38fF
C79302 INVX1_LOC_194/A VSS 0.42fF
C79303 NOR2X1_LOC_459/B VSS 0.19fF
C79304 NOR2X1_LOC_437/Y VSS 0.01fF
C79305 NOR2X1_LOC_426/Y VSS 0.25fF
C79306 NOR2X1_LOC_448/B VSS 0.13fF
C79307 INVX1_LOC_135/A VSS -45.56fF
C79308 NOR2X1_LOC_415/A VSS 0.12fF
C79309 NOR2X1_LOC_619/A VSS 0.18fF
C79310 NOR2X1_LOC_629/B VSS 0.13fF
C79311 NOR2X1_LOC_607/Y VSS 0.16fF
C79312 NOR2X1_LOC_607/A VSS 0.40fF
C79313 NAND2X1_LOC_192/B VSS 0.11fF
C79314 NAND2X1_LOC_190/Y VSS -0.75fF
C79315 NOR2X1_LOC_187/Y VSS 0.07fF
C79316 NOR2X1_LOC_34/B VSS 0.24fF
C79317 INVX1_LOC_5/A VSS 0.64fF
C79318 INVX1_LOC_25/A VSS 0.60fF
C79319 NAND2X1_LOC_182/A VSS 0.33fF
C79320 INVX1_LOC_249/A VSS -0.32fF
C79321 INVX1_LOC_227/Y VSS 0.15fF
C79322 INVX1_LOC_238/Y VSS 0.21fF
C79323 INVX1_LOC_238/A VSS -0.19fF
C79324 INVX1_LOC_216/Y VSS 0.15fF
C79325 INVX1_LOC_205/Y VSS 0.06fF
C79326 NOR2X1_LOC_400/A VSS -0.01fF
C79327 INVX1_LOC_35/A VSS 1.42fF
C79328 NOR2X1_LOC_91/A VSS -4.42fF
C79329 INVX1_LOC_157/A VSS -0.19fF
C79330 NOR2X1_LOC_458/B VSS -0.14fF
C79331 NOR2X1_LOC_778/B VSS -0.41fF
C79332 NAND2X1_LOC_276/Y VSS 0.34fF
C79333 NOR2X1_LOC_637/A VSS 0.12fF
C79334 NOR2X1_LOC_644/B VSS 0.32fF
C79335 NOR2X1_LOC_596/Y VSS 0.11fF
C79336 NAND2X1_LOC_579/A VSS 0.37fF
C79337 NAND2X1_LOC_573/Y VSS -1.67fF
C79338 NAND2X1_LOC_552/A VSS 0.18fF
C79339 INVX1_LOC_219/A VSS 0.12fF
C79340 NAND2X1_LOC_563/A VSS 0.20fF
C79341 NAND2X1_LOC_541/Y VSS 0.11fF
C79342 NAND2X1_LOC_569/A VSS 0.01fF
C79343 NOR2X1_LOC_518/Y VSS 0.12fF
C79344 NOR2X1_LOC_710/A VSS 0.12fF
C79345 NAND2X1_LOC_725/A VSS 0.65fF
C79346 NAND2X1_LOC_708/Y VSS 0.19fF
C79347 NOR2X1_LOC_757/A VSS 0.25fF
C79348 NAND2X1_LOC_733/B VSS 0.26fF
C79349 NAND2X1_LOC_717/Y VSS 0.17fF
C79350 INVX1_LOC_282/Y VSS 0.36fF
C79351 INVX1_LOC_172/A VSS 0.49fF
C79352 INVX1_LOC_305/A VSS 0.74fF
C79353 NOR2X1_LOC_751/Y VSS 0.16fF
C79354 INVX1_LOC_293/A VSS -0.20fF
C79355 NOR2X1_LOC_496/Y VSS 0.30fF
C79356 NOR2X1_LOC_243/Y VSS 0.13fF
C79357 NOR2X1_LOC_267/A VSS -0.84fF
C79358 INVX1_LOC_124/Y VSS 0.68fF
C79359 INVX1_LOC_134/A VSS 0.39fF
C79360 NOR2X1_LOC_286/Y VSS 0.10fF
C79361 NOR2X1_LOC_824/A VSS -1.31fF
C79362 INVX1_LOC_13/Y VSS 1.06fF
C79363 NOR2X1_LOC_218/Y VSS 0.12fF
C79364 NOR2X1_LOC_219/Y VSS -0.95fF
C79365 NOR2X1_LOC_207/A VSS 0.09fF
C79366 NOR2X1_LOC_194/Y VSS 0.09fF
C79367 NOR2X1_LOC_403/B VSS 0.17fF
C79368 INVX1_LOC_200/A VSS 0.53fF
C79369 NOR2X1_LOC_468/Y VSS 0.35fF
C79370 NOR2X1_LOC_798/A VSS 0.38fF
C79371 NOR2X1_LOC_434/Y VSS -0.10fF
C79372 NOR2X1_LOC_717/B VSS 0.61fF
C79373 NOR2X1_LOC_617/Y VSS -0.53fF
C79374 NOR2X1_LOC_606/Y VSS 0.05fF
C79375 NOR2X1_LOC_590/A VSS 0.65fF
C79376 INVX1_LOC_258/A VSS 0.11fF
C79377 NOR2X1_LOC_92/Y VSS 0.90fF
C79378 INVX1_LOC_99/Y VSS 0.21fF
C79379 INVX1_LOC_97/Y VSS 0.10fF
C79380 NAND2X1_LOC_11/Y VSS 1.12fF
C79381 NAND2X1_LOC_59/B VSS 0.52fF
C79382 NAND2X1_LOC_21/Y VSS 0.29fF
C79383 NOR2X1_LOC_196/A VSS 0.23fF
C79384 INPUT_3 VSS 0.34fF
C79385 INPUT_2 VSS 0.27fF
C79386 INVX1_LOC_204/Y VSS 0.24fF
C79387 INVX1_LOC_259/Y VSS 0.19fF
C79388 INVX1_LOC_215/A VSS 0.44fF
C79389 INVX1_LOC_248/A VSS 0.22fF
C79390 INVX1_LOC_237/Y VSS -0.64fF
C79391 NAND2X1_LOC_381/Y VSS -0.01fF
C79392 NOR2X1_LOC_82/A VSS 0.67fF
C79393 INVX1_LOC_27/A VSS 0.90fF
C79394 NAND2X1_LOC_363/B VSS 0.90fF
C79395 NAND2X1_LOC_860/A VSS 0.48fF
C79396 NOR2X1_LOC_810/A VSS 0.18fF
C79397 INVX1_LOC_228/Y VSS 0.07fF
C79398 NOR2X1_LOC_255/Y VSS 0.50fF
C79399 NAND2X1_LOC_564/B VSS -1.15fF
C79400 NAND2X1_LOC_543/Y VSS 0.20fF
C79401 NOR2X1_LOC_770/A VSS -0.11fF
C79402 NOR2X1_LOC_780/A VSS 0.12fF
C79403 NOR2X1_LOC_710/B VSS 0.08fF
C79404 NAND2X1_LOC_794/B VSS 0.19fF
C79405 INVX1_LOC_248/Y VSS -0.20fF
C79406 NAND2X1_LOC_784/A VSS 0.33fF
C79407 INVX1_LOC_278/Y VSS -0.30fF
C79408 NOR2X1_LOC_664/Y VSS 0.27fF
C79409 NAND2X1_LOC_733/A VSS 0.16fF
C79410 INVX1_LOC_284/Y VSS 0.11fF
C79411 NOR2X1_LOC_232/Y VSS 0.29fF
C79412 NOR2X1_LOC_15/Y VSS 0.77fF
C79413 NOR2X1_LOC_240/Y VSS 0.16fF
C79414 NOR2X1_LOC_667/A VSS 0.81fF
C79415 NOR2X1_LOC_288/A VSS -0.23fF
C79416 NOR2X1_LOC_843/A VSS -0.12fF
C79417 NOR2X1_LOC_276/B VSS 0.19fF
C79418 NOR2X1_LOC_483/B VSS 0.31fF
C79419 NOR2X1_LOC_254/A VSS 0.24fF
C79420 NOR2X1_LOC_223/B VSS -0.15fF
C79421 NOR2X1_LOC_440/Y VSS -0.48fF
C79422 INVX1_LOC_164/Y VSS 0.15fF
C79423 NOR2X1_LOC_401/Y VSS 0.09fF
C79424 NOR2X1_LOC_413/Y VSS 0.02fF
C79425 NOR2X1_LOC_480/A VSS -0.34fF
C79426 NOR2X1_LOC_476/Y VSS 0.09fF
C79427 INVX1_LOC_188/A VSS 0.26fF
C79428 NOR2X1_LOC_446/A VSS 0.09fF
C79429 NOR2X1_LOC_464/B VSS 0.07fF
C79430 NOR2X1_LOC_424/Y VSS 0.22fF
C79431 NOR2X1_LOC_616/Y VSS 0.13fF
C79432 INVX1_LOC_15/Y VSS 0.27fF
C79433 NOR2X1_LOC_643/Y VSS 0.26fF
C79434 NAND2X1_LOC_30/Y VSS -3.04fF
C79435 NOR2X1_LOC_61/B VSS 0.17fF
C79436 INVX1_LOC_51/A VSS 0.18fF
C79437 NOR2X1_LOC_605/B VSS 0.07fF
C79438 NOR2X1_LOC_627/Y VSS 0.11fF
C79439 NOR2X1_LOC_637/Y VSS 0.19fF
C79440 INVX1_LOC_247/Y VSS 0.18fF
C79441 INVX1_LOC_236/Y VSS 0.28fF
C79442 INVX1_LOC_269/Y VSS 0.15fF
C79443 INVX1_LOC_269/A VSS -11.00fF
C79444 INVX1_LOC_258/Y VSS 0.22fF
C79445 INPUT_6 VSS 0.05fF
C79446 INVX1_LOC_214/Y VSS 0.22fF
C79447 INVX1_LOC_214/A VSS 0.25fF
C79448 INVX1_LOC_225/A VSS 0.96fF
C79449 INVX1_LOC_203/Y VSS 0.15fF
C79450 NOR2X1_LOC_820/A VSS 0.09fF
C79451 INVX1_LOC_36/A VSS 1.09fF
C79452 INVX1_LOC_40/Y VSS 0.33fF
C79453 INVX1_LOC_11/A VSS 1.34fF
C79454 NAND2X1_LOC_391/Y VSS 0.13fF
C79455 NAND2X1_LOC_787/A VSS 0.31fF
C79456 NOR2X1_LOC_811/A VSS 0.08fF
C79457 NAND2X1_LOC_555/Y VSS 1.68fF
C79458 NOR2X1_LOC_643/A VSS 0.32fF
C79459 NAND2X1_LOC_553/A VSS 0.08fF
C79460 NOR2X1_LOC_178/Y VSS 0.17fF
C79461 NAND2X1_LOC_564/A VSS 0.23fF
C79462 INVX1_LOC_224/Y VSS -2.05fF
C79463 INVX1_LOC_9/Y VSS 0.26fF
C79464 NAND2X1_LOC_802/A VSS 0.32fF
C79465 NAND2X1_LOC_785/B VSS 0.24fF
C79466 NAND2X1_LOC_738/B VSS 0.34fF
C79467 NAND2X1_LOC_725/Y VSS 0.69fF
C79468 NAND2X1_LOC_724/Y VSS 0.24fF
C79469 NOR2X1_LOC_614/Y VSS 0.23fF
C79470 NAND2X1_LOC_734/B VSS 0.33fF
C79471 NAND2X1_LOC_711/B VSS -0.33fF
C79472 NOR2X1_LOC_641/B VSS 0.42fF
C79473 NOR2X1_LOC_231/B VSS 0.13fF
C79474 NOR2X1_LOC_285/Y VSS 0.09fF
C79475 INVX1_LOC_50/A VSS 0.48fF
C79476 NOR2X1_LOC_244/B VSS 0.16fF
C79477 INVX1_LOC_34/A VSS -6.36fF
C79478 INVX1_LOC_116/A VSS 0.09fF
C79479 INVX1_LOC_130/A VSS 0.09fF
C79480 NAND2X1_LOC_213/A VSS 0.64fF
C79481 NAND2X1_LOC_149/Y VSS 0.22fF
C79482 NOR2X1_LOC_772/B VSS 0.44fF
C79483 NOR2X1_LOC_489/B VSS 0.13fF
C79484 INVX1_LOC_204/A VSS 0.11fF
C79485 NOR2X1_LOC_401/B VSS 0.07fF
C79486 NOR2X1_LOC_690/A VSS -3.40fF
C79487 NOR2X1_LOC_470/A VSS 0.13fF
C79488 NOR2X1_LOC_210/A VSS 0.33fF
C79489 NOR2X1_LOC_655/B VSS 0.52fF
C79490 NOR2X1_LOC_644/Y VSS 0.15fF
C79491 NOR2X1_LOC_637/B VSS 0.43fF
C79492 NOR2X1_LOC_657/Y VSS 0.15fF
C79493 NOR2X1_LOC_658/Y VSS 0.08fF
C79494 NOR2X1_LOC_615/Y VSS 0.13fF
C79495 NOR2X1_LOC_598/B VSS 1.45fF
C79496 D_INPUT_1 VSS 0.92fF
C79497 NOR2X1_LOC_33/A VSS 0.27fF
C79498 NAND2X1_LOC_33/Y VSS 0.17fF
C79499 NOR2X1_LOC_538/B VSS 0.41fF
C79500 NOR2X1_LOC_626/Y VSS 0.15fF
C79501 NOR2X1_LOC_604/Y VSS 0.02fF
C79502 INVX1_LOC_268/A VSS 0.15fF
C79503 INVX1_LOC_213/Y VSS 0.29fF
C79504 INVX1_LOC_202/A VSS 0.44fF
C79505 INVX1_LOC_279/Y VSS 0.32fF
C79506 INVX1_LOC_224/A VSS 0.41fF
C79507 INVX1_LOC_235/Y VSS 0.49fF
C79508 INVX1_LOC_235/A VSS 0.12fF
C79509 NOR2X1_LOC_829/Y VSS 0.13fF
C79510 NOR2X1_LOC_811/B VSS 0.07fF
C79511 NOR2X1_LOC_806/Y VSS 0.24fF
C79512 NOR2X1_LOC_460/B VSS 0.13fF
C79513 NOR2X1_LOC_379/Y VSS 0.13fF
C79514 NOR2X1_LOC_382/Y VSS 0.06fF
C79515 NOR2X1_LOC_636/B VSS 0.30fF
C79516 NOR2X1_LOC_653/B VSS 0.09fF
C79517 NOR2X1_LOC_186/Y VSS 0.68fF
C79518 NAND2X1_LOC_571/B VSS 0.25fF
C79519 NAND2X1_LOC_557/Y VSS 0.16fF
C79520 NAND2X1_LOC_565/B VSS 0.17fF
C79521 INVX1_LOC_226/Y VSS 0.19fF
C79522 INVX1_LOC_8/Y VSS 0.25fF
C79523 NOR2X1_LOC_769/A VSS 0.12fF
C79524 NAND2X1_LOC_803/B VSS 0.51fF
C79525 GATE_741 VSS 0.27fF
C79526 NAND2X1_LOC_741/Y VSS 0.07fF
C79527 NAND2X1_LOC_740/Y VSS 0.15fF
C79528 NOR2X1_LOC_790/B VSS 0.49fF
C79529 NAND2X1_LOC_727/Y VSS 0.11fF
C79530 NAND2X1_LOC_726/Y VSS 0.14fF
C79531 NAND2X1_LOC_785/A VSS 0.34fF
C79532 INVX1_LOC_303/A VSS 1.05fF
C79533 NOR2X1_LOC_262/Y VSS 0.18fF
C79534 NAND2X1_LOC_84/Y VSS 0.37fF
C79535 NAND2X1_LOC_721/B VSS 0.01fF
C79536 NOR2X1_LOC_296/Y VSS -0.10fF
C79537 NOR2X1_LOC_242/A VSS 0.44fF
C79538 NOR2X1_LOC_285/A VSS 0.12fF
C79539 NOR2X1_LOC_252/Y VSS 0.15fF
C79540 INVX1_LOC_124/A VSS -1.49fF
C79541 NOR2X1_LOC_274/Y VSS 0.15fF
C79542 NOR2X1_LOC_230/Y VSS 0.13fF
C79543 NAND2X1_LOC_222/B VSS 0.07fF
C79544 NAND2X1_LOC_214/Y VSS 0.19fF
C79545 NAND2X1_LOC_214/B VSS 0.61fF
C79546 NAND2X1_LOC_35/Y VSS 0.47fF
C79547 NOR2X1_LOC_443/Y VSS 0.10fF
C79548 NOR2X1_LOC_488/Y VSS 0.19fF
C79549 NOR2X1_LOC_226/A VSS -7.10fF
C79550 NOR2X1_LOC_445/Y VSS 0.40fF
C79551 NOR2X1_LOC_500/A VSS 0.61fF
C79552 NOR2X1_LOC_778/A VSS 0.38fF
C79553 NOR2X1_LOC_478/A VSS 0.14fF
C79554 NOR2X1_LOC_471/Y VSS 0.03fF
C79555 NOR2X1_LOC_470/B VSS 0.18fF
C79556 NOR2X1_LOC_453/Y VSS 0.12fF
C79557 NOR2X1_LOC_454/Y VSS 0.56fF
C79558 NOR2X1_LOC_411/Y VSS 0.15fF
C79559 INVX1_LOC_64/A VSS -7.98fF
C79560 NOR2X1_LOC_411/A VSS 0.47fF
C79561 INVX1_LOC_166/A VSS 0.29fF
C79562 NOR2X1_LOC_400/B VSS 0.13fF
C79563 INVX1_LOC_136/A VSS -11.39fF
C79564 NOR2X1_LOC_647/B VSS 0.34fF
C79565 NOR2X1_LOC_669/Y VSS -0.29fF
C79566 NOR2X1_LOC_632/Y VSS 0.44fF
C79567 NOR2X1_LOC_636/A VSS -0.11fF
C79568 NOR2X1_LOC_197/A VSS 0.32fF
C79569 NAND2X1_LOC_53/Y VSS 0.66fF
C79570 INVX1_LOC_13/A VSS 0.69fF
C79571 NAND2X1_LOC_35/B VSS 0.21fF
C79572 NOR2X1_LOC_27/Y VSS 0.07fF
C79573 INVX1_LOC_45/A VSS 1.22fF
C79574 INVX1_LOC_245/Y VSS -0.23fF
C79575 INVX1_LOC_289/Y VSS 0.33fF
C79576 INVX1_LOC_223/Y VSS 0.82fF
C79577 INVX1_LOC_278/A VSS 0.34fF
C79578 INVX1_LOC_267/Y VSS 0.15fF
C79579 INVX1_LOC_267/A VSS 0.12fF
C79580 INVX1_LOC_201/Y VSS 0.62fF
C79581 INVX1_LOC_212/A VSS 0.09fF
C79582 NOR2X1_LOC_852/A VSS 0.09fF
C79583 NOR2X1_LOC_836/Y VSS 0.07fF
C79584 NOR2X1_LOC_817/Y VSS 0.44fF
C79585 NOR2X1_LOC_381/Y VSS 0.44fF
C79586 NOR2X1_LOC_828/Y VSS 0.30fF
C79587 NAND2X1_LOC_392/A VSS 0.31fF
C79588 NOR2X1_LOC_635/A VSS 0.03fF
C79589 NAND2X1_LOC_581/Y VSS 0.11fF
C79590 INVX1_LOC_246/Y VSS 0.06fF
C79591 INVX1_LOC_230/Y VSS 0.43fF
C79592 INVX1_LOC_229/A VSS -0.19fF
C79593 NAND2X1_LOC_559/Y VSS 0.15fF
C79594 INVX1_LOC_7/Y VSS 0.28fF
C79595 NOR2X1_LOC_769/B VSS 0.13fF
C79596 INVX1_LOC_289/A VSS 0.42fF
C79597 NAND2X1_LOC_736/Y VSS 0.54fF
C79598 NAND2X1_LOC_739/B VSS 0.33fF
C79599 NAND2X1_LOC_729/Y VSS 0.24fF
C79600 NAND2X1_LOC_728/Y VSS 0.20fF
C79601 NAND2X1_LOC_783/Y VSS -0.01fF
C79602 INVX1_LOC_299/A VSS 0.66fF
C79603 NAND2X1_LOC_773/Y VSS 0.67fF
C79604 NOR2X1_LOC_65/B VSS 0.69fF
C79605 NOR2X1_LOC_287/A VSS 0.33fF
C79606 NOR2X1_LOC_284/B VSS 0.13fF
C79607 NOR2X1_LOC_295/Y VSS 0.36fF
C79608 NOR2X1_LOC_481/A VSS 0.09fF
C79609 NOR2X1_LOC_273/Y VSS 0.24fF
C79610 INVX1_LOC_108/Y VSS 0.69fF
C79611 NAND2X1_LOC_222/A VSS 0.19fF
C79612 NOR2X1_LOC_498/Y VSS 0.38fF
C79613 NOR2X1_LOC_189/A VSS 0.49fF
C79614 INVX1_LOC_57/Y VSS 0.39fF
C79615 NOR2X1_LOC_455/Y VSS 0.17fF
C79616 NOR2X1_LOC_456/Y VSS 0.29fF
C79617 NOR2X1_LOC_328/Y VSS -0.38fF
C79618 NOR2X1_LOC_432/Y VSS 0.07fF
C79619 NOR2X1_LOC_447/Y VSS 0.24fF
C79620 NOR2X1_LOC_410/Y VSS -0.02fF
C79621 INVX1_LOC_256/A VSS 0.55fF
C79622 NOR2X1_LOC_613/Y VSS 0.06fF
C79623 NOR2X1_LOC_647/A VSS 0.08fF
C79624 NOR2X1_LOC_646/A VSS -0.24fF
C79625 NOR2X1_LOC_100/A VSS 0.49fF
C79626 NAND2X1_LOC_99/Y VSS 0.12fF
C79627 NOR2X1_LOC_602/A VSS 0.23fF
C79628 NOR2X1_LOC_679/Y VSS -0.14fF
C79629 INVX1_LOC_272/Y VSS 0.36fF
C79630 NOR2X1_LOC_510/Y VSS 0.41fF
C79631 NOR2X1_LOC_639/B VSS 0.08fF
C79632 INVX1_LOC_288/Y VSS 0.15fF
C79633 INVX1_LOC_288/A VSS 0.09fF
C79634 NOR2X1_LOC_20/Y VSS 0.15fF
C79635 INVX1_LOC_39/A VSS -0.58fF
C79636 NOR2X1_LOC_67/A VSS -5.02fF
C79637 INVX1_LOC_2/A VSS 0.71fF
C79638 INVX1_LOC_41/A VSS 0.93fF
C79639 INVX1_LOC_244/Y VSS -0.05fF
C79640 INVX1_LOC_277/Y VSS 0.15fF
C79641 INVX1_LOC_277/A VSS 0.58fF
C79642 INVX1_LOC_211/Y VSS 0.40fF
C79643 INVX1_LOC_266/A VSS 0.03fF
C79644 INVX1_LOC_222/Y VSS 0.32fF
C79645 INVX1_LOC_233/Y VSS 0.86fF
C79646 INVX1_LOC_233/A VSS 0.69fF
C79647 INVX1_LOC_200/Y VSS 0.36fF
C79648 INVX1_LOC_255/Y VSS 0.39fF
C79649 INVX1_LOC_310/A VSS -0.03fF
C79650 NOR2X1_LOC_852/B VSS 0.04fF
C79651 NOR2X1_LOC_837/Y VSS -0.05fF
C79652 NOR2X1_LOC_859/A VSS 0.29fF
C79653 NOR2X1_LOC_844/Y VSS 0.11fF
C79654 NOR2X1_LOC_807/B VSS 0.30fF
C79655 NOR2X1_LOC_793/Y VSS 0.36fF
C79656 INVX1_LOC_245/A VSS 0.12fF
C79657 NAND2X1_LOC_563/Y VSS -2.09fF
C79658 NAND2X1_LOC_562/Y VSS 0.28fF
C79659 INVX1_LOC_6/Y VSS 0.25fF
C79660 NAND2X1_LOC_763/B VSS 0.51fF
C79661 NAND2X1_LOC_796/B VSS 0.38fF
C79662 NAND2X1_LOC_778/Y VSS -1.91fF
C79663 NOR2X1_LOC_750/Y VSS -0.00fF
C79664 INVX1_LOC_304/Y VSS -1.45fF
C79665 NAND2X1_LOC_785/Y VSS 0.19fF
C79666 INVX1_LOC_132/A VSS -1.61fF
C79667 NOR2X1_LOC_294/Y VSS -0.74fF
C79668 NOR2X1_LOC_250/Y VSS 0.41fF
C79669 NOR2X1_LOC_272/Y VSS 0.83fF
C79670 NOR2X1_LOC_261/Y VSS 0.27fF
C79671 NAND2X1_LOC_341/A VSS 0.46fF
C79672 INVX1_LOC_119/A VSS 0.89fF
C79673 NAND2X1_LOC_218/B VSS 0.63fF
C79674 INVX1_LOC_110/Y VSS -0.08fF
C79675 NOR2X1_LOC_420/Y VSS 0.11fF
C79676 INVX1_LOC_17/Y VSS 0.22fF
C79677 NOR2X1_LOC_479/B VSS 0.24fF
C79678 NOR2X1_LOC_458/Y VSS 0.07fF
C79679 NOR2X1_LOC_431/Y VSS 0.11fF
C79680 NOR2X1_LOC_705/B VSS 0.37fF
C79681 NOR2X1_LOC_448/Y VSS 0.12fF
C79682 NOR2X1_LOC_689/Y VSS -0.27fF
C79683 NOR2X1_LOC_689/A VSS 0.32fF
C79684 INVX1_LOC_251/Y VSS 0.02fF
C79685 NOR2X1_LOC_624/A VSS 0.12fF
C79686 NOR2X1_LOC_620/Y VSS 0.11fF
C79687 NOR2X1_LOC_647/Y VSS -0.04fF
C79688 INVX1_LOC_55/A VSS 0.12fF
C79689 NOR2X1_LOC_75/Y VSS 0.16fF
C79690 INVX1_LOC_59/A VSS 1.21fF
C79691 NOR2X1_LOC_93/Y VSS 0.13fF
C79692 NOR2X1_LOC_32/B VSS 0.20fF
C79693 NOR2X1_LOC_201/A VSS 0.35fF
C79694 INVX1_LOC_250/A VSS 0.37fF
C79695 NOR2X1_LOC_667/Y VSS 0.08fF
C79696 INVX1_LOC_287/Y VSS 0.31fF
C79697 INVX1_LOC_287/A VSS 0.41fF
C79698 INVX1_LOC_298/Y VSS 0.35fF
C79699 INVX1_LOC_276/Y VSS 0.06fF
C79700 INVX1_LOC_276/A VSS 0.80fF
C79701 INVX1_LOC_265/A VSS -0.10fF
C79702 INVX1_LOC_254/Y VSS 0.30fF
C79703 INVX1_LOC_254/A VSS 0.33fF
C79704 NOR2X1_LOC_195/A VSS 0.12fF
C79705 INVX1_LOC_17/A VSS 1.55fF
C79706 NOR2X1_LOC_34/A VSS 0.15fF
C79707 INVX1_LOC_21/A VSS -5.22fF
C79708 NAND2X1_LOC_9/Y VSS 0.32fF
C79709 INVX1_LOC_243/Y VSS 0.28fF
C79710 INVX1_LOC_232/Y VSS 0.21fF
C79711 NOR2X1_LOC_837/B VSS 0.42fF
C79712 NOR2X1_LOC_848/Y VSS 0.22fF
C79713 NOR2X1_LOC_846/Y VSS 0.13fF
C79714 NOR2X1_LOC_826/Y VSS 0.11fF
C79715 INVX1_LOC_58/A VSS 1.79fF
C79716 NOR2X1_LOC_808/A VSS 0.35fF
C79717 NOR2X1_LOC_795/Y VSS 0.32fF
C79718 NOR2X1_LOC_815/Y VSS 0.20fF
C79719 GATE_579 VSS 0.14fF
C79720 INVX1_LOC_242/Y VSS 0.06fF
.ends

