*** static inverter ***
*
* ngSPICE compensed 3-inverter inverter with feedback inverter
*
*
* Author: Jan Belohoubek, 01/2020
* jan.belohoubek@fit.cvut.cz
*
* https://users.fit.cvut.cz/~belohja4/
*
*
* **************************************

.subckt INV A O VSS VDD

*** Compensation Inverter Chain ***
Xinv0 O2 VSS A  VDD INVX1
Xinv1 O1 VSS O2 VDD INVX1
Xinv2 O  VSS O1 VDD INVX1


*** Compensation feedback inverter ***
Xpmos O1 O VDD VDD VSS LaserTrig SUBCKT_PMOS beamDistance = beamDistanceTop ch_w=1u ch_l=0.2u mos_ad=1p mos_pd=5u mos_as=1.2p mos_ps=6.6u

Xnmos O1 O VSS VSS psubIn LaserTrig SUBCKT_NMOS beamDistance = beamDistanceBot ch_w=0.5u ch_l=0.2u mos_ad=0.5p mos_pd=3u mos_as=0.66p mos_ps=4.6u

* common NMOS substarte virtual node
XpsubIn psubIn VSS PSUB_IN

.ends
