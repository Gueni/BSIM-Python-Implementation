* SPICE3 file created from POR2X1.ext - technology: scmos

.subckt POR2X1 VDD GND B A Y
X0 O CTRL2 GND GND NMOS_MAGIC ad=1.04p pd=5.2u as=3.39p ps=17u w=2u l=0.2u
**devattr s=S d=D
X1 O CTRL VDD VDD PMOS_MAGIC ad=1.72p pd=7.8u as=5.94p ps=27.8u w=3.3u l=0.2u
**devattr s=S d=D
X2 CTRL2 CTRL VDD VDD PMOS_MAGIC ad=1.95p pd=8.8u as=0p ps=0u w=3.9u l=0.2u
**devattr s=S d=D
X3 a_112_344# A a_92_344# VDD PMOS_MAGIC ad=0.42p pd=2.6u as=0.21p ps=2u w=0.7u l=0.2u
**devattr s=S d=D
X4 CTRL GND GND GND NMOS_MAGIC ad=1.75p pd=8u as=0p ps=0u w=3.5u l=0.2u
**devattr s=S d=D
X5 Y O VDD VDD PMOS_MAGIC ad=1.95p pd=8.8u as=0p ps=0u w=3.9u l=0.2u
**devattr s=S d=D
X6 a_52_28# B GND GND NMOS_MAGIC ad=0.44p pd=3.8u as=0p ps=0u w=0.4u l=0.2u
**devattr s=S d=D
X7 a_52_28# A GND GND NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=0.4u l=0.2u
**devattr s=S d=D
X8 O CTRL2 a_112_344# VDD PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=0.7u l=0.2u
**devattr s=S d=D
X9 CTRL GND VDD VDD PMOS_MAGIC ad=0.2p pd=1.8u as=0p ps=0u w=0.4u l=0.2u
**devattr s=S d=D
X10 CTRL2 CTRL GND GND NMOS_MAGIC ad=0.2p pd=1.8u as=0p ps=0u w=0.4u l=0.2u
**devattr s=S d=D
X11 a_92_344# B VDD VDD PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=0.7u l=0.2u
**devattr s=S d=D
X12 O CTRL a_52_28# GND NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=0.4u l=0.2u
**devattr s=S d=D
X13 Y O GND GND NMOS_MAGIC ad=1p pd=5u as=0p ps=0u w=2u l=0.2u
**devattr s=S d=D
C0 Y O 0.05fF
C1 B a_52_28# 0.02fF
C2 CTRL2 CTRL 0.32fF
C3 VDD a_112_344# 0.05fF
C4 A a_52_28# 0.06fF
C5 CTRL2 O 0.27fF
C6 CTRL O 0.15fF
C7 B A 0.51fF
C8 B VDD 0.38fF
C9 A VDD 0.28fF
C10 Y VDD 0.54fF
C11 O a_112_344# 0.07fF
C12 O a_52_28# 0.21fF
C13 A CTRL2 0.13fF
C14 VDD CTRL2 1.37fF
C15 B O 0.04fF
C16 A CTRL 0.16fF
C17 VDD CTRL 1.32fF
C18 A O 0.11fF
C19 VDD O 0.59fF
.ends

