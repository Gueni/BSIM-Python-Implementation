* SPICE3 file created from SECLIBAND.ext - technology: scmos

.subckt NOR3X1_LOC a_8_256# a_100_256# Y gnd vdd A B C
X0 a_8_256# B a_100_256# vdd PMOS_MAGIC ad=4.78p pd=21.2u as=4.8p ps=21.2u w=3u l=0.2u
X1 a_8_256# A vdd vdd PMOS_MAGIC ad=0p pd=0u as=1.8p ps=7.2u w=3u l=0.2u
X2 vdd A a_8_256# vdd PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=3u l=0.2u
X3 a_100_256# C Y vdd PMOS_MAGIC ad=0p pd=0u as=1.8p ps=7.2u w=3u l=0.2u
X4 Y A gnd gnd NMOS_MAGIC ad=1.1p pd=6.2u as=1.1p ps=6.2u w=1u l=0.2u
X5 Y C a_100_256# vdd PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=3u l=0.2u
X6 a_100_256# B a_8_256# vdd PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=3u l=0.2u
X7 gnd B Y gnd NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=1u l=0.2u
X8 Y C gnd gnd NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=1u l=0.2u
C0 a_100_256# vdd 0.45fF
C1 a_8_256# A 0.03fF
C2 C a_100_256# 0.02fF
C3 a_8_256# vdd 1.16fF
C4 B A 0.23fF
C5 Y a_100_256# 0.76fF
C6 B vdd 0.22fF
C7 C B 0.16fF
C8 A vdd 0.22fF
C9 Y B 0.02fF
C10 Y A 0.01fF
C11 C vdd 0.30fF
C12 Y vdd 0.07fF
C13 C Y 0.12fF
C14 a_100_256# a_8_256# 0.94fF
C15 a_100_256# B 0.02fF
C16 a_8_256# B 0.03fF
C17 Y gnd 0.20fF
C18 C gnd 0.29fF
C19 a_100_256# gnd 0.00fF
C20 a_8_256# gnd 0.00fF
C21 B gnd 0.29fF
C22 A gnd 0.31fF
C23 vdd gnd 3.25fF
.ends

.subckt CELM2X1 a_36_24# Y a_8_24# gnd vdd A B
X0 Y a_8_24# vdd vdd PMOS_MAGIC ad=1p pd=5u as=1.2p ps=5.2u w=2u l=0.2u
**devattr s=S d=D
X1 a_36_296# B vdd vdd PMOS_MAGIC ad=0.6p pd=4.6u as=0p ps=0u w=2u l=0.2u
**devattr s=S d=D
X2 a_8_24# A a_36_24# gnd NMOS_MAGIC ad=1p pd=5u as=0.6p ps=4.6u w=2u l=0.2u
**devattr s=S d=D
X3 Y a_8_24# gnd gnd NMOS_MAGIC ad=0.5p pd=3u as=1.1p ps=5.2u w=1u l=0.2u
**devattr s=S d=D
X4 a_36_24# B gnd gnd NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=2u l=0.2u
**devattr s=S d=D
X5 a_8_24# A a_36_296# vdd PMOS_MAGIC ad=1p pd=5u as=0p ps=0u w=2u l=0.2u
**devattr s=S d=D
C0 a_8_24# A 0.12fF
C1 B A 0.41fF
C2 a_8_24# vdd 0.41fF
C3 Y a_8_24# 0.51fF
C4 B vdd 0.25fF
C5 a_36_24# a_8_24# 0.00fF
C6 A vdd 0.20fF
C7 Y vdd 0.39fF
C8 a_36_296# a_8_24# 0.00fF
C9 a_8_24# B 0.38fF
C10 Y gnd 0.17fF
C11 a_8_24# gnd 0.45fF
C12 B gnd 0.17fF
C13 A gnd 0.25fF
C14 vdd gnd 1.95fF
.ends

.subckt INVX1_LOC Y gnd vdd A
X0 Y A gnd gnd NMOS_MAGIC ad=0.5p pd=3u as=0.5p ps=3u w=1u l=0.2u
X1 Y A vdd vdd PMOS_MAGIC ad=1p pd=5u as=1p ps=5u w=2u l=0.2u
C0 Y A 0.08fF
C1 Y vdd 0.39fF
C2 A vdd 0.20fF
C3 Y gnd 0.07fF
C4 A gnd 0.37fF
C5 vdd gnd 1.52fF
.ends


* Top level circuit SECLIBAND

.subckt SECLIBAND INVX1_LOC_1/vdd INVX1_LOC_1/gnd CELM2X1_4/A A1 CELM2X1_0/B B1 INVX1_LOC_0/Y INVX1_LOC_1/Y

XNOR3X1_LOC_0 NOR3X1_LOC_0/a_8_256# NOR3X1_LOC_0/a_100_256# INVX1_LOC_0/A INVX1_LOC_1/gnd INVX1_LOC_1/vdd
+ NOR3X1_LOC_0/A NOR3X1_LOC_0/B NOR3X1_LOC_0/C NOR3X1_LOC
XNOR3X1_LOC_1 NOR3X1_LOC_1/a_8_256# NOR3X1_LOC_1/a_100_256# INVX1_LOC_1/A INVX1_LOC_1/gnd INVX1_LOC_1/vdd
+ NOR3X1_LOC_1/A NOR3X1_LOC_1/B NOR3X1_LOC_1/A NOR3X1_LOC
XCELM2X1_0 CELM2X1_0/a_36_24# NOR3X1_LOC_0/C CELM2X1_0/a_8_24# INVX1_LOC_1/gnd INVX1_LOC_1/vdd
+ CELM2X1_4/A CELM2X1_0/B CELM2X1
XCELM2X1_1 CELM2X1_1/a_36_24# NOR3X1_LOC_0/A CELM2X1_1/a_8_24# INVX1_LOC_1/gnd INVX1_LOC_1/vdd
+ CELM2X1_4/A B1 CELM2X1
XCELM2X1_2 CELM2X1_2/a_36_24# NOR3X1_LOC_0/B CELM2X1_2/a_8_24# INVX1_LOC_1/gnd INVX1_LOC_1/vdd
+ A1 CELM2X1_0/B CELM2X1
XCELM2X1_3 CELM2X1_3/a_36_24# NOR3X1_LOC_1/B CELM2X1_3/a_8_24# INVX1_LOC_1/gnd INVX1_LOC_1/vdd
+ A1 B1 CELM2X1
XCELM2X1_4 CELM2X1_4/a_36_24# NOR3X1_LOC_1/A CELM2X1_4/a_8_24# INVX1_LOC_1/gnd INVX1_LOC_1/vdd
+ CELM2X1_4/A A1 CELM2X1
XINVX1_LOC_0 INVX1_LOC_0/Y INVX1_LOC_1/gnd INVX1_LOC_1/vdd INVX1_LOC_0/A INVX1_LOC
XINVX1_LOC_1 INVX1_LOC_1/Y INVX1_LOC_1/gnd INVX1_LOC_1/vdd INVX1_LOC_1/A INVX1_LOC
C0 INVX1_LOC_1/A NOR3X1_LOC_1/A 0.00fF
C1 INVX1_LOC_1/vdd CELM2X1_2/a_8_24# -0.00fF
C2 INVX1_LOC_1/vdd NOR3X1_LOC_0/C 0.11fF
C3 CELM2X1_2/a_8_24# NOR3X1_LOC_1/A 0.02fF
C4 NOR3X1_LOC_0/A CELM2X1_2/a_36_24# 0.00fF
C5 NOR3X1_LOC_0/C CELM2X1_3/a_8_24# 0.05fF
C6 NOR3X1_LOC_1/B NOR3X1_LOC_1/A 0.25fF
C7 NOR3X1_LOC_0/C NOR3X1_LOC_1/A 0.03fF
C8 INVX1_LOC_1/A INVX1_LOC_0/A 0.06fF
C9 NOR3X1_LOC_0/A CELM2X1_3/a_8_24# 0.05fF
C10 NOR3X1_LOC_0/A NOR3X1_LOC_1/A 1.27fF
C11 CELM2X1_4/A A1 0.65fF
C12 NOR3X1_LOC_0/B INVX1_LOC_1/vdd 0.07fF
C13 CELM2X1_3/a_36_24# NOR3X1_LOC_1/A 0.00fF
C14 CELM2X1_0/a_36_24# NOR3X1_LOC_1/A 0.00fF
C15 CELM2X1_4/A B1 0.01fF
C16 CELM2X1_0/a_8_24# CELM2X1_4/A 0.06fF
C17 NOR3X1_LOC_0/B CELM2X1_3/a_8_24# 0.54fF
C18 INVX1_LOC_0/A NOR3X1_LOC_1/B 0.03fF
C19 NOR3X1_LOC_0/B NOR3X1_LOC_1/A 0.03fF
C20 CELM2X1_1/a_36_24# NOR3X1_LOC_1/A 0.00fF
C21 CELM2X1_4/A CELM2X1_0/B 0.01fF
C22 B1 A1 0.02fF
C23 CELM2X1_0/a_8_24# A1 0.02fF
C24 CELM2X1_2/a_36_24# NOR3X1_LOC_1/A 0.00fF
C25 A1 CELM2X1_0/B 0.75fF
C26 CELM2X1_1/a_8_24# A1 0.02fF
C27 B1 CELM2X1_0/B 0.51fF
C28 CELM2X1_4/A CELM2X1_4/a_8_24# 0.06fF
C29 B1 CELM2X1_1/a_8_24# 0.04fF
C30 CELM2X1_0/a_8_24# CELM2X1_0/B 0.02fF
C31 INVX1_LOC_1/A INVX1_LOC_0/Y 0.43fF
C32 NOR3X1_LOC_0/C CELM2X1_4/A 0.14fF
C33 INVX1_LOC_1/vdd CELM2X1_3/a_8_24# 0.00fF
C34 INVX1_LOC_1/vdd NOR3X1_LOC_1/A 0.00fF
C35 CELM2X1_3/a_8_24# NOR3X1_LOC_1/A 0.03fF
C36 A1 CELM2X1_2/a_8_24# 0.02fF
C37 A1 CELM2X1_4/a_8_24# 0.02fF
C38 CELM2X1_1/a_8_24# CELM2X1_0/B 0.02fF
C39 B1 CELM2X1_2/a_8_24# 0.02fF
C40 INVX1_LOC_1/A INVX1_LOC_1/Y 0.31fF
C41 NOR3X1_LOC_0/C A1 0.03fF
C42 NOR3X1_LOC_0/C B1 0.98fF
C43 INVX1_LOC_0/A INVX1_LOC_1/vdd 0.00fF
C44 NOR3X1_LOC_0/A A1 0.24fF
C45 NOR3X1_LOC_0/C CELM2X1_0/B 0.03fF
C46 B1 NOR3X1_LOC_0/A 0.03fF
C47 INVX1_LOC_0/A NOR3X1_LOC_1/A 0.46fF
C48 NOR3X1_LOC_0/C CELM2X1_1/a_8_24# 0.57fF
C49 NOR3X1_LOC_0/B A1 0.31fF
C50 NOR3X1_LOC_0/B B1 0.24fF
C51 NOR3X1_LOC_0/a_100_256# NOR3X1_LOC_0/C 0.04fF
C52 NOR3X1_LOC_0/A CELM2X1_0/B 0.03fF
C53 NOR3X1_LOC_0/C CELM2X1_2/a_8_24# 0.05fF
C54 NOR3X1_LOC_1/a_8_256# NOR3X1_LOC_0/a_100_256# 0.33fF
C55 NOR3X1_LOC_0/C NOR3X1_LOC_1/B 0.04fF
C56 INVX1_LOC_1/vdd CELM2X1_4/A 0.00fF
C57 NOR3X1_LOC_0/a_8_256# NOR3X1_LOC_1/B 0.29fF
C58 NOR3X1_LOC_0/a_8_256# NOR3X1_LOC_0/C 0.05fF
C59 NOR3X1_LOC_0/A CELM2X1_2/a_8_24# 0.69fF
C60 NOR3X1_LOC_1/a_100_256# INVX1_LOC_1/vdd 0.20fF
C61 CELM2X1_4/A NOR3X1_LOC_1/A 0.14fF
C62 NOR3X1_LOC_0/A NOR3X1_LOC_1/B 0.26fF
C63 NOR3X1_LOC_0/C NOR3X1_LOC_0/A 0.04fF
C64 INVX1_LOC_1/vdd INVX1_LOC_0/Y 0.21fF
C65 NOR3X1_LOC_0/B CELM2X1_2/a_8_24# 0.00fF
C66 INVX1_LOC_1/vdd A1 0.00fF
C67 INVX1_LOC_1/vdd B1 0.07fF
C68 NOR3X1_LOC_0/B NOR3X1_LOC_1/B 0.06fF
C69 INVX1_LOC_1/vdd CELM2X1_0/a_8_24# 0.00fF
C70 NOR3X1_LOC_0/B NOR3X1_LOC_0/C 0.16fF
C71 B1 CELM2X1_3/a_8_24# 0.02fF
C72 A1 NOR3X1_LOC_1/A 0.03fF
C73 B1 NOR3X1_LOC_1/A 0.01fF
C74 CELM2X1_0/a_8_24# NOR3X1_LOC_1/A 0.55fF
C75 NOR3X1_LOC_0/A CELM2X1_3/a_36_24# 0.00fF
C76 INVX1_LOC_1/vdd CELM2X1_0/B 0.05fF
C77 INVX1_LOC_1/vdd CELM2X1_1/a_8_24# 0.00fF
C78 NOR3X1_LOC_0/B NOR3X1_LOC_0/A 0.03fF
C79 CELM2X1_0/B NOR3X1_LOC_1/A 0.01fF
C80 INVX1_LOC_1/A INVX1_LOC_1/vdd 0.08fF
C81 CELM2X1_1/a_8_24# NOR3X1_LOC_1/A 0.03fF
C82 INVX1_LOC_0/Y INVX1_LOC_1/gnd 0.10fF
C83 NOR3X1_LOC_1/A INVX1_LOC_1/gnd 0.30fF
C84 NOR3X1_LOC_1/B INVX1_LOC_1/gnd 0.17fF
C85 CELM2X1_0/B INVX1_LOC_1/gnd -0.22fF
C86 A1 INVX1_LOC_1/gnd 0.21fF
C87 NOR3X1_LOC_0/A INVX1_LOC_1/gnd 0.20fF
C88 B1 INVX1_LOC_1/gnd 0.14fF
C89 CELM2X1_4/A INVX1_LOC_1/gnd 0.16fF
C90 NOR3X1_LOC_0/C INVX1_LOC_1/gnd 0.13fF
C91 INVX1_LOC_1/A INVX1_LOC_1/gnd -0.22fF
C92 INVX1_LOC_0/A INVX1_LOC_1/gnd 0.34fF
C93 NOR3X1_LOC_0/B INVX1_LOC_1/gnd 0.17fF
C94 INVX1_LOC_1/vdd INVX1_LOC_1/gnd 0.02fF

.ends

