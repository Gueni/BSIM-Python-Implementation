* SPICE3 file created from POR2X1.ext - technology: scmos

*.subckt POR2X1 VDD GND B A Y a_24_28# O m4_240_n4# a_8_268# a_36_268# CTRL2 a_88_268# CTRL
.subckt POR2X1 VDD GND B A Y
X0 O B a_88_268# VDD PMOS_MAGIC ad=1.76p pd=8.2u as=0.78p ps=5.8u w=2.6u l=0.2u
**devattr s=S d=D
X1 CTRL GND VDD VDD PMOS_MAGIC ad=0.2p pd=1.8u as=5.28p ps=24.2u w=0.4u l=0.2u
**devattr s=S d=D
X2 O A a_36_268# VDD PMOS_MAGIC ad=0p pd=0u as=0.78p ps=5.8u w=2.6u l=0.2u
**devattr s=S d=D
X3 CTRL2 CTRL VDD VDD PMOS_MAGIC ad=1.95p pd=8.8u as=0p ps=0u w=3.9u l=0.2u
**devattr s=S d=D
X4 Y O GND GND NMOS_MAGIC ad=0.8p pd=4.2u as=2.83p ps=13.6u w=1.6u l=0.2u
**devattr s=S d=D
X5 O CTRL2 GND GND NMOS_MAGIC ad=0.84p pd=5.4u as=0p ps=0u w=1.2u l=0.2u
**devattr s=S d=D
X6 CTRL2 CTRL GND GND NMOS_MAGIC ad=0.2p pd=1.8u as=0p ps=0u w=0.4u l=0.2u
**devattr s=S d=D
X7 CTRL GND GND GND NMOS_MAGIC ad=1.75p pd=8u as=0p ps=0u w=3.5u l=0.2u
**devattr s=S d=D
X8 a_88_268# A a_8_268# VDD PMOS_MAGIC ad=0p pd=0u as=2.86p ps=12.6u w=2.6u l=0.2u
**devattr s=S d=D
X9 a_36_268# B a_8_268# VDD PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=2.6u l=0.2u
**devattr s=S d=D
X10 O B a_24_28# GND NMOS_MAGIC ad=0p pd=0u as=1.4p ps=6.6u w=0.4u l=0.2u
**devattr s=S d=D
X11 O A a_24_28# GND NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=0.4u l=0.2u
**devattr s=S d=D
X12 Y O VDD VDD PMOS_MAGIC ad=1.95p pd=8.8u as=0p ps=0u w=3.9u l=0.2u
**devattr s=S d=D
X13 a_8_268# CTRL2 VDD VDD PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=2.6u l=0.2u
**devattr s=S d=D
X14 a_24_28# CTRL3 GND GND NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=1.2u l=0.2u
**devattr s=S d=D
X15 O CTRL3 VDD VDD PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=0.4u l=0.2u
**devattr s=S d=D

*X33 CTRL3 CTRL2 VDD VDD PMOS_MAGIC ad=1.95p pd=8.8u as=0p ps=0u w=3.9u l=0.2u
*X66 CTRL3 CTRL2 GND GND NMOS_MAGIC ad=0.2p pd=1.8u as=0p ps=0u w=0.4u l=0.2u

X11 CTRL3 CTRL2 VDD VDD PMOS_MAGIC ad=0.2p pd=1.8u as=5.28p ps=24.2u w=0.4u l=0.2u
X77 CTRL3 CTRL2 GND GND NMOS_MAGIC ad=1.75p pd=8u as=0p ps=0u w=3.5u l=0.2u

C0 a_24_28# A 0.01fF
C1 CTRL2 VDD 0.73fF
C2 CTRL2 CTRL 0.37fF
C3 CTRL VDD 1.51fF
C4 CTRL2 O 1.08fF
C5 VDD B 0.41fF
C6 CTRL2 A 0.06fF
C7 O VDD 0.77fF
C8 CTRL O 0.21fF
C9 VDD A 0.31fF
C10 a_8_268# VDD 0.41fF
C11 CTRL A 0.06fF
C12 O B 0.12fF
C13 VDD Y 0.54fF
C14 B A 0.68fF
C15 O A 0.15fF
C16 a_8_268# B 0.01fF
C17 O a_8_268# 0.08fF
C18 O Y 0.05fF
C19 a_8_268# A 0.01fF
C20 a_8_268# a_36_268# 0.00fF
C21 a_24_28# B 0.01fF
C22 a_8_268# a_88_268# 0.00fF
C23 O a_24_28# 0.28fF
C24 Y GND 0.50fF
C25 A GND 0.45fF
C26 B GND 0.27fF
C27 VDD GND 4.94fF
C28 GND GND -0.17fF

*C29 m4_240_n4# GND 0.01fF
Rcorr m4_240_n4# GND 0.001

C30 a_24_28# GND 0.32fF
C31 a_8_268# GND -0.00fF
C32 O GND 0.50fF
C33 CTRL GND 0.65fF
C34 CTRL2 GND 0.44fF
.ends
