* SPICE3 file created from SECLIBAND.ext - technology: scmos

.subckt NOR3X1_LOC a_8_256# a_100_256# Y gnd vdd A B C
X0 a_8_256# B a_100_256# vdd PMOS_MAGIC ad=4.78p pd=21.2u as=4.8p ps=21.2u w=3u l=0.2u
X1 a_8_256# A vdd vdd PMOS_MAGIC ad=0p pd=0u as=1.8p ps=7.2u w=3u l=0.2u
X2 vdd A a_8_256# vdd PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=3u l=0.2u
X3 a_100_256# C Y vdd PMOS_MAGIC ad=0p pd=0u as=1.8p ps=7.2u w=3u l=0.2u
X4 Y A gnd gnd NMOS_MAGIC ad=1.1p pd=6.2u as=1.1p ps=6.2u w=1u l=0.2u
X5 Y C a_100_256# vdd PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=3u l=0.2u
X6 a_100_256# B a_8_256# vdd PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=3u l=0.2u
X7 gnd B Y gnd NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=1u l=0.2u
X8 Y C gnd gnd NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=1u l=0.2u
C0 vdd a_100_256# 0.45fF
C1 vdd Y 0.07fF
C2 B vdd 0.22fF
C3 A vdd 0.22fF
C4 a_8_256# a_100_256# 0.94fF
C5 C a_100_256# 0.02fF
C6 B a_8_256# 0.03fF
C7 C Y 0.12fF
C8 B C 0.16fF
C9 Y a_100_256# 0.76fF
C10 A a_8_256# 0.03fF
C11 B a_100_256# 0.02fF
C12 B Y 0.02fF
C13 vdd a_8_256# 1.16fF
C14 A Y 0.01fF
C15 vdd C 0.30fF
C16 B A 0.23fF
C17 Y gnd 0.20fF
C18 C gnd 0.29fF
C19 a_100_256# gnd 0.00fF
C20 a_8_256# gnd 0.00fF
C21 B gnd 0.29fF
C22 A gnd 0.31fF
C23 vdd gnd 3.25fF
.ends

.subckt CELM2X1 a_36_24# Y a_8_24# gnd vdd A B
X0 Y a_8_24# vdd vdd PMOS_MAGIC ad=1p pd=5u as=1.2p ps=5.2u w=2u l=0.2u
**devattr s=S d=D
X1 a_36_296# B vdd vdd PMOS_MAGIC ad=0.6p pd=4.6u as=0p ps=0u w=2u l=0.2u
**devattr s=S d=D
X2 a_8_24# A a_36_24# gnd NMOS_MAGIC ad=1p pd=5u as=0.6p ps=4.6u w=2u l=0.2u
**devattr s=S d=D
X3 Y a_8_24# gnd gnd NMOS_MAGIC ad=0.5p pd=3u as=1.1p ps=5.2u w=1u l=0.2u
**devattr s=S d=D
X4 a_36_24# B gnd gnd NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=2u l=0.2u
**devattr s=S d=D
X5 a_8_24# A a_36_296# vdd PMOS_MAGIC ad=1p pd=5u as=0p ps=0u w=2u l=0.2u
**devattr s=S d=D
C0 B vdd 0.25fF
C1 A vdd 0.20fF
C2 Y a_8_24# 0.51fF
C3 a_8_24# a_36_296# 0.00fF
C4 a_36_24# a_8_24# 0.00fF
C5 B a_8_24# 0.38fF
C6 A a_8_24# 0.12fF
C7 vdd a_8_24# 0.41fF
C8 vdd Y 0.39fF
C9 B A 0.41fF
C10 Y gnd 0.17fF
C11 a_8_24# gnd 0.45fF
C12 B gnd 0.17fF
C13 A gnd 0.25fF
C14 vdd gnd 1.95fF
.ends

.subckt INVX1_LOC Y gnd vdd A
X0 Y A gnd gnd NMOS_MAGIC ad=0.5p pd=3u as=0.5p ps=3u w=1u l=0.2u
X1 Y A vdd vdd PMOS_MAGIC ad=1p pd=5u as=1p ps=5u w=2u l=0.2u
C0 Y vdd 0.39fF
C1 A vdd 0.20fF
C2 Y A 0.08fF
C3 Y gnd 0.07fF
C4 A gnd 0.37fF
C5 vdd gnd 1.52fF
.ends


* Top level circuit SECLIBAND

.subckt SECLIBAND INVX1_LOC_0/vdd NOR3X1_LOC_1/A CELM2X1_0/A A1 CELM2X1_0/B B1 INVX1_LOC_0/Y INVX1_LOC_1/Y

XNOR3X1_LOC_0 NOR3X1_LOC_0/a_8_256# NOR3X1_LOC_0/a_100_256# INVX1_LOC_0/A NOR3X1_LOC_1/A INVX1_LOC_0/vdd NOR3X1_LOC_0/A
+ NOR3X1_LOC_0/B NOR3X1_LOC_0/C NOR3X1_LOC
XNOR3X1_LOC_1 NOR3X1_LOC_1/a_8_256# NOR3X1_LOC_1/a_100_256# INVX1_LOC_1/A NOR3X1_LOC_1/A INVX1_LOC_0/vdd NOR3X1_LOC_1/A
+ NOR3X1_LOC_1/B NOR3X1_LOC_1/A NOR3X1_LOC
XCELM2X1_0 CELM2X1_0/a_36_24# NOR3X1_LOC_0/C CELM2X1_0/a_8_24# NOR3X1_LOC_1/A INVX1_LOC_0/vdd
+ CELM2X1_0/A CELM2X1_0/B CELM2X1
XCELM2X1_1 CELM2X1_1/a_36_24# NOR3X1_LOC_0/A CELM2X1_1/a_8_24# NOR3X1_LOC_1/A INVX1_LOC_0/vdd
+ CELM2X1_0/A B1 CELM2X1
XCELM2X1_2 CELM2X1_2/a_36_24# NOR3X1_LOC_0/B CELM2X1_2/a_8_24# NOR3X1_LOC_1/A INVX1_LOC_0/vdd
+ A1 CELM2X1_0/B CELM2X1
XCELM2X1_3 CELM2X1_3/a_36_24# NOR3X1_LOC_1/B CELM2X1_3/a_8_24# NOR3X1_LOC_1/A INVX1_LOC_0/vdd
+ A1 B1 CELM2X1
XINVX1_LOC_0 INVX1_LOC_0/Y NOR3X1_LOC_1/A INVX1_LOC_0/vdd INVX1_LOC_0/A INVX1_LOC
XINVX1_LOC_1 INVX1_LOC_1/Y NOR3X1_LOC_1/A INVX1_LOC_0/vdd INVX1_LOC_1/A INVX1_LOC
C0 NOR3X1_LOC_0/B CELM2X1_2/a_8_24# 0.00fF
C1 INVX1_LOC_0/vdd A1 0.00fF
C2 INVX1_LOC_0/vdd CELM2X1_3/a_8_24# 0.00fF
C3 NOR3X1_LOC_0/a_8_256# NOR3X1_LOC_1/B 0.29fF
C4 INVX1_LOC_0/vdd NOR3X1_LOC_1/a_100_256# 0.20fF
C5 INVX1_LOC_0/vdd INVX1_LOC_0/A 0.00fF
C6 NOR3X1_LOC_0/A CELM2X1_3/a_36_24# 0.00fF
C7 NOR3X1_LOC_0/B INVX1_LOC_0/vdd 0.07fF
C8 INVX1_LOC_0/A INVX1_LOC_1/A 0.06fF
C9 INVX1_LOC_0/vdd CELM2X1_0/B 0.05fF
C10 NOR3X1_LOC_0/C NOR3X1_LOC_1/B 0.04fF
C11 B1 NOR3X1_LOC_0/A 0.03fF
C12 NOR3X1_LOC_0/C CELM2X1_0/A 0.14fF
C13 INVX1_LOC_0/A NOR3X1_LOC_1/B 0.03fF
C14 INVX1_LOC_0/vdd CELM2X1_2/a_8_24# -0.00fF
C15 NOR3X1_LOC_0/B NOR3X1_LOC_1/B 0.06fF
C16 NOR3X1_LOC_0/C B1 0.98fF
C17 CELM2X1_2/a_36_24# NOR3X1_LOC_0/A 0.00fF
C18 CELM2X1_0/B CELM2X1_0/A 0.01fF
C19 A1 B1 0.02fF
C20 B1 CELM2X1_3/a_8_24# 0.02fF
C21 INVX1_LOC_0/vdd INVX1_LOC_1/A 0.08fF
C22 NOR3X1_LOC_0/C CELM2X1_1/a_8_24# 0.57fF
C23 NOR3X1_LOC_0/B B1 0.24fF
C24 CELM2X1_0/B B1 0.51fF
C25 INVX1_LOC_0/vdd CELM2X1_0/A 0.00fF
C26 CELM2X1_0/B CELM2X1_1/a_8_24# 0.02fF
C27 CELM2X1_2/a_8_24# B1 0.02fF
C28 NOR3X1_LOC_0/C NOR3X1_LOC_0/A 0.04fF
C29 INVX1_LOC_0/vdd B1 0.07fF
C30 A1 NOR3X1_LOC_0/A 0.21fF
C31 NOR3X1_LOC_0/A CELM2X1_3/a_8_24# 0.05fF
C32 CELM2X1_0/B CELM2X1_0/a_8_24# 0.02fF
C33 NOR3X1_LOC_0/a_8_256# NOR3X1_LOC_0/C 0.05fF
C34 INVX1_LOC_0/vdd CELM2X1_1/a_8_24# 0.00fF
C35 NOR3X1_LOC_0/B NOR3X1_LOC_0/A 0.03fF
C36 CELM2X1_0/B NOR3X1_LOC_0/A 0.03fF
C37 NOR3X1_LOC_1/a_8_256# NOR3X1_LOC_0/a_100_256# 0.33fF
C38 A1 NOR3X1_LOC_0/C 0.01fF
C39 NOR3X1_LOC_0/a_100_256# NOR3X1_LOC_0/C 0.04fF
C40 NOR3X1_LOC_0/C CELM2X1_3/a_8_24# 0.05fF
C41 CELM2X1_0/A B1 0.01fF
C42 CELM2X1_2/a_8_24# NOR3X1_LOC_0/A 0.69fF
C43 NOR3X1_LOC_0/B NOR3X1_LOC_0/C 0.16fF
C44 INVX1_LOC_0/vdd INVX1_LOC_0/Y 0.21fF
C45 CELM2X1_0/B NOR3X1_LOC_0/C 0.03fF
C46 NOR3X1_LOC_0/B A1 0.31fF
C47 INVX1_LOC_1/A INVX1_LOC_0/Y 0.43fF
C48 NOR3X1_LOC_0/B CELM2X1_3/a_8_24# 0.54fF
C49 A1 CELM2X1_0/B 0.18fF
C50 INVX1_LOC_1/A INVX1_LOC_1/Y 0.31fF
C51 CELM2X1_2/a_8_24# NOR3X1_LOC_0/C 0.05fF
C52 A1 CELM2X1_2/a_8_24# 0.02fF
C53 B1 CELM2X1_1/a_8_24# 0.04fF
C54 CELM2X1_0/a_8_24# CELM2X1_0/A 0.06fF
C55 INVX1_LOC_0/vdd NOR3X1_LOC_0/C 0.11fF
C56 NOR3X1_LOC_0/A NOR3X1_LOC_1/B 0.26fF
C57 INVX1_LOC_0/Y NOR3X1_LOC_1/A 0.10fF
C58 NOR3X1_LOC_1/B NOR3X1_LOC_1/A 0.34fF
C59 CELM2X1_0/B NOR3X1_LOC_1/A -0.22fF
C60 A1 NOR3X1_LOC_1/A -0.03fF
C61 NOR3X1_LOC_0/A NOR3X1_LOC_1/A 0.20fF
C62 B1 NOR3X1_LOC_1/A 0.14fF
C63 CELM2X1_0/A NOR3X1_LOC_1/A 0.09fF
C64 NOR3X1_LOC_0/C NOR3X1_LOC_1/A 0.13fF
C65 INVX1_LOC_1/A NOR3X1_LOC_1/A -0.19fF
C66 INVX1_LOC_0/A NOR3X1_LOC_1/A 0.35fF
C67 NOR3X1_LOC_0/B NOR3X1_LOC_1/A 0.17fF
C68 INVX1_LOC_0/vdd NOR3X1_LOC_1/A 0.02fF

.ends

