VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO INVX1
  CLASS BLOCK ;
  FOREIGN INVX1 ;
  ORIGIN 0.900 0.300 ;
  SIZE 3.500 BY 10.800 ;
  OBS
      LAYER metal1 ;
        RECT -0.200 9.700 1.800 10.300 ;
        RECT 0.200 7.400 0.600 9.700 ;
        RECT 0.200 1.900 0.600 2.700 ;
        RECT 0.200 0.300 0.600 1.600 ;
        RECT 1.000 0.600 1.400 9.400 ;
        RECT -0.200 -0.300 1.800 0.300 ;
  END
END INVX1
END LIBRARY

