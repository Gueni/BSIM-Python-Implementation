*** TEST 005 - partitioning ***
*
* ngSPICE test for PLS experiments
*
* AES SBOX PLS test init file generator - protected dualRail SBOX area illuminated
*
* Author: Jan Belohoubek, 08/2020
* jan.belohoubek@fit.cvut.cz
*
* https://users.fit.cvut.cz/~belohja4/
*
*
* **************************************

.include ../../models.lib
.include ../../tsmc180nmcmos.lib
.include secLibDualRail.spice

* **************************************
* --- Test ---
* **************************************

* --- Settings
.param showPlots = 0
.param writeFile = 1
.param run_inputSet = 0

* redefine defaults ...
.include test00X_settings.inc

.csparam showPlots = {showPlots}
.csparam writeFile = {writeFile}
.csparam run_inputSet = {run_inputSet}

.global showPlots writeFile run_inputSet

* --- End of Settins

Vtrig LaserTrig 0 0 PWL(0ns 0V 40ns 0V 41ns SUPP)

.param beamDistanceTop = 0
.param beamDistanceBot = 0

.global LaserTrig beamDistanceTop beamDistanceBot

* --- inputs
Vvin0 INPUT_0 0 0 PWL(0ns 0V 5ns  0V 7ns  0V)
Vvin1 INPUT_1 0 0 PWL(0ns 0V 6ns  0V 8ns  0V)
Vvin2 INPUT_2 0 0 PWL(0ns 0V 7ns  0V 9ns  0V)
Vvin3 INPUT_3 0 0 PWL(0ns 0V 8ns  0V 10ns 0V)
Vvin4 INPUT_4 0 0 PWL(0ns 0V 9ns  0V 11ns 0V)
Vvin5 INPUT_5 0 0 PWL(0ns 0V 10ns 0V 12ns 0V)
Vvin6 INPUT_6 0 0 PWL(0ns 0V 11ns 0V 13ns 0V)
Vvin7 INPUT_7 0 0 PWL(0ns 0V 12ns 0V 14ns 0V)

Vvin0D D_INPUT_0 0 0 PWL(0ns 0V 5ns  0V 7ns  0V)
Vvin1D D_INPUT_1 0 0 PWL(0ns 0V 6ns  0V 8ns  0V)
Vvin2D D_INPUT_2 0 0 PWL(0ns 0V 7ns  0V 9ns  0V)
Vvin3D D_INPUT_3 0 0 PWL(0ns 0V 8ns  0V 10ns 0V)
Vvin4D D_INPUT_4 0 0 PWL(0ns 0V 9ns  0V 11ns 0V)
Vvin5D D_INPUT_5 0 0 PWL(0ns 0V 10ns 0V 12ns 0V)
Vvin6D D_INPUT_6 0 0 PWL(0ns 0V 11ns 0V 13ns 0V)
Vvin7D D_INPUT_7 0 0 PWL(0ns 0V 12ns 0V 14ns 0V)


* --- circuit layout model

Xsbox1 
+ INVX1_1164/A INVX1_1506/A INVX1_1096/A INVX1_1095/A INVX1_1386/A INVX1_1385/A INVX1_526/A INVX1_300/A INVX1_114/A INVX1_136/A INVX1_620/A INVX1_142/A INVX1_135/A INVX1_1344/A INVX1_755/A INVX1_592/A INVX1_591/A INVX1_1654/A INVX1_86/A INVX1_838/A INVX1_1068/A INVX1_756/A INVX1_1170/A INVX1_588/A INVX1_829/A INVX1_1250/A INVX1_796/A INVX1_795/A INVX1_587/A INVX1_186/A INVX1_1256/A INVX1_844/A INVX1_600/A INVX1_242/A INVX1_598/A INVX1_241/A INVX1_1212/A INVX1_1211/A INVX1_738/A INVX1_1026/A INVX1_492/A INVX1_556/A INVX1_491/A INVX1_922/A INVX1_921/A INVX1_511/A INVX1_252/A INVX1_12/A INVX1_1496/A INVX1_979/A INVX1_46/A 
+ INVX1_512/A INVX1_38/A INVX1_980/A INVX1_199/A INVX1_200/A INVX1_187/A INVX1_1222/A INVX1_764/A INVX1_258/A INVX1_160/A INVX1_163/A INVX1_582/A INVX1_1648/A INVX1_468/A INVX1_860/A INVX1_859/A INVX1_1175/A INVX1_818/A INVX1_817/A INVX1_1163/A INVX1_1525/A INVX1_1505/A INVX1_112/A INVX1_111/A INVX1_607/A INVX1_608/A INVX1_852/A INVX1_1387/A INVX1_1388/A INVX1_851/A INVX1_774/A INVX1_773/A INVX1_658/A INVX1_1192/A INVX1_1191/A INVX1_842/A INVX1_657/A INVX1_841/A INVX1_525/A INVX1_257/A INVX1_251/A INVX1_299/A INVX1_37/A INVX1_11/A INVX1_619/A INVX1_141/A INVX1_159/A INVX1_113/A INVX1_1221/A INVX1_188/A INVX1_164/A 
+ INVX1_45/A INVX1_1238/A INVX1_830/A INVX1_1237/A INVX1_763/A INVX1_1343/A INVX1_916/A INVX1_915/A INVX1_752/A INVX1_1176/A INVX1_1003/A INVX1_328/A INVX1_1004/A INVX1_1392/A INVX1_288/A INVX1_578/A INVX1_1627/A INVX1_566/A INVX1_618/A INVX1_976/A INVX1_1628/A INVX1_452/A INVX1_751/A INVX1_327/A INVX1_287/A INVX1_1391/A INVX1_809/A INVX1_1038/A INVX1_810/A INVX1_96/A INVX1_1384/A INVX1_1526/A INVX1_1653/A INVX1_1067/A INVX1_837/A INVX1_85/A INVX1_1694/A INVX1_1693/A INVX1_1037/A INVX1_95/A INVX1_1383/A INVX1_1495/A INVX1_310/A INVX1_309/A INVX1_1486/A INVX1_866/A INVX1_185/A INVX1_1255/A INVX1_843/A INVX1_555/A INVX1_737/A 
+ INVX1_597/A INVX1_599/A INVX1_1485/A INVX1_865/A INVX1_451/A INVX1_577/A INVX1_617/A INVX1_565/A INVX1_975/A INVX1_1169/A INVX1_1249/A INVX1_1602/A INVX1_581/A INVX1_1647/A INVX1_467/A INVX1_1382/A INVX1_646/A INVX1_1053/A INVX1_645/A INVX1_1054/A INVX1_222/A INVX1_221/A INVX1_1025/A INVX1_1381/A INVX1_1030/A INVX1_1029/A INVX1_552/A INVX1_1500/A INVX1_551/A INVX1_1499/A INVX1_1601/A INVX1_51/Y INVX1_24/Y INVX1_23/Y INVX1_52/Y INVX1_741/Y INVX1_742/Y INVX1_1198/Y INVX1_272/Y INVX1_612/Y INVX1_271/Y INVX1_823/Y INVX1_824/Y INVX1_611/Y INVX1_548/Y INVX1_547/Y INVX1_170/Y INVX1_169/Y INVX1_1197/Y INVX1_176/Y INVX1_175/Y 
+ INVX1_822/Y INVX1_821/Y INVX1_317/Y INVX1_318/Y INVX1_541/Y INVX1_542/Y INVX1_833/Y INVX1_834/Y INVX1_61/Y INVX1_62/Y INVX1_127/Y INVX1_128/Y INVX1_189/Y INVX1_190/Y INVX1_1377/Y INVX1_1378/Y INVX1_1021/Y INVX1_1022/Y INVX1_94/Y INVX1_93/Y INVX1_72/Y INVX1_71/Y INVX1_76/Y INVX1_75/Y INVX1_30/Y INVX1_29/Y INVX1_131/Y INVX1_132/Y INVX1_20/Y INVX1_44/Y INVX1_19/Y INVX1_43/Y INVX1_35/Y INVX1_102/Y INVX1_314/Y INVX1_208/Y INVX1_207/Y INVX1_313/Y INVX1_101/Y INVX1_36/Y INVX1_747/Y INVX1_748/Y INVX1_1640/Y INVX1_1639/Y INVX1_140/Y INVX1_139/Y INVX1_6/Y INVX1_97/Y INVX1_5/Y 
+ INVX1_110/Y INVX1_98/Y INVX1_109/Y INVX1_204/Y INVX1_203/Y INVX1_239/Y INVX1_240/Y INVX1_118/Y INVX1_117/Y INVX1_554/Y INVX1_489/Y INVX1_490/Y INVX1_553/Y INVX1_509/Y INVX1_510/Y INVX1_1398/Y INVX1_1397/Y INVX1_653/Y INVX1_654/Y INVX1_754/Y INVX1_753/Y INVX1_750/Y INVX1_154/Y INVX1_153/Y INVX1_87/Y INVX1_749/Y INVX1_88/Y INVX1_1060/Y INVX1_1059/Y INVX1_124/Y INVX1_123/Y INVX1_79/Y INVX1_80/Y INVX1_180/Y INVX1_179/Y INVX1_471/Y INVX1_472/Y INVX1_265/Y INVX1_266/Y INVX1_369/Y INVX1_370/Y INVX1_814/Y INVX1_813/Y INVX1_1198/A INVX1_548/A INVX1_547/A INVX1_1197/A INVX1_176/A INVX1_175/A INVX1_822/A INVX1_821/A 
+ INVX1_541/A INVX1_1377/A INVX1_1378/A INVX1_131/A INVX1_132/A INVX1_747/A INVX1_748/A INVX1_1640/A INVX1_1639/A INVX1_239/A INVX1_240/A INVX1_653/A INVX1_654/A INVX1_750/A INVX1_749/A INVX1_1060/A INVX1_1059/A INVX1_369/A INVX1_370/A NOR3X1_175/B NOR3X1_821/B NOR3X1_1599/C NOR3X1_747/B NOR3X1_653/B INVX1_1196/Y INVX1_1195/Y INVX1_546/Y INVX1_544/Y INVX1_545/Y INVX1_543/Y INVX1_174/Y INVX1_173/Y INVX1_820/Y INVX1_819/Y INVX1_1520/Y INVX1_1373/Y INVX1_1519/Y INVX1_1374/Y INVX1_537/Y INVX1_539/Y INVX1_540/Y INVX1_538/Y INVX1_1375/Y INVX1_1376/Y INVX1_643/Y INVX1_745/Y INVX1_746/Y INVX1_644/Y 
+ INVX1_1637/Y INVX1_1636/Y INVX1_1638/Y INVX1_1635/Y INVX1_125/Y INVX1_528/Y INVX1_527/Y INVX1_126/Y INVX1_145/Y INVX1_146/Y INVX1_174/A INVX1_173/A INVX1_820/A INVX1_819/A INVX1_1520/A INVX1_1373/A INVX1_1519/A INVX1_1374/A INVX1_537/A INVX1_539/A INVX1_540/A INVX1_538/A INVX1_745/A INVX1_746/A INVX1_528/A INVX1_527/A NOR3X1_1519/B INVX1_58/Y INVX1_57/Y INVX1_1370/Y INVX1_1372/Y INVX1_1371/Y INVX1_1369/Y INVX1_535/Y INVX1_536/Y INVX1_1370/A INVX1_1372/A INVX1_1371/A INVX1_1369/A NOR3X1_1371/C NOR3X1_1369/B INVX1_1364/Y INVX1_1362/Y INVX1_1363/Y INVX1_1361/Y INVX1_1368/Y INVX1_1366/Y INVX1_1367/Y INVX1_1365/Y INVX1_1364/A INVX1_1363/A 
+ INVX1_1366/A INVX1_1365/A 
+ VSS VDD 
+ NOR3X1_1270/C NOR3X1_1269/B NOR3X1_1270/A NOR3X1_1579/C NOR3X1_1580/A NOR3X1_1580/B NOR3X1_377/C NOR3X1_367/B NOR3X1_267/C NOR3X1_378/C NOR3X1_368/B NOR3X1_268/C NOR3X1_377/A NOR3X1_264/B NOR3X1_1187/C NOR3X1_250/C NOR3X1_1188/C NOR3X1_263/A NOR3X1_263/B NOR3X1_267/A NOR3X1_367/A NOR3X1_249/A NOR3X1_1187/A NOR3X1_249/C NOR3X1_811/A NOR3X1_811/C NOR3X1_812/C NOR3X1_120/B NOR3X1_873/C NOR3X1_1217/C NOR3X1_984/C NOR3X1_1399/A NOR3X1_1509/A NOR3X1_1218/C NOR3X1_1399/C NOR3X1_161/A NOR3X1_1509/C NOR3X1_161/C NOR3X1_790/C NOR3X1_983/A NOR3X1_1217/A NOR3X1_162/C NOR3X1_983/C NOR3X1_789/A NOR3X1_789/C NOR3X1_1400/C NOR3X1_590/C NOR3X1_874/C NOR3X1_589/A NOR3X1_119/A NOR3X1_119/B 
+ NOR3X1_1510/C NOR3X1_589/C NOR3X1_873/A NOR3X1_1529/C NOR3X1_458/C NOR3X1_987/C NOR3X1_988/C NOR3X1_457/A NOR3X1_1205/A NOR3X1_1205/C NOR3X1_987/A NOR3X1_1206/C NOR3X1_261/A NOR3X1_261/C NOR3X1_262/C NOR3X1_1355/C NOR3X1_1356/A NOR3X1_1356/B NOR3X1_1530/C NOR3X1_457/C NOR3X1_1529/A NOR3X1_1214/C NOR3X1_39/A NOR3X1_513/A NOR3X1_39/C NOR3X1_513/C NOR3X1_157/C NOR3X1_1213/A NOR3X1_158/C NOR3X1_1331/A NOR3X1_1213/C NOR3X1_1010/C NOR3X1_1331/C NOR3X1_1332/C NOR3X1_157/A NOR3X1_1009/A NOR3X1_1009/C NOR3X1_1041/A NOR3X1_1041/C NOR3X1_40/C NOR3X1_514/C NOR3X1_1042/C NOR3X1_1533/C NOR3X1_1330/C NOR3X1_794/C NOR3X1_31/A NOR3X1_1329/A NOR3X1_793/A NOR3X1_31/C NOR3X1_1329/C NOR3X1_793/C 
+ NOR3X1_961/A NOR3X1_1534/C NOR3X1_32/C NOR3X1_14/C NOR3X1_961/C NOR3X1_254/C NOR3X1_962/C NOR3X1_13/A NOR3X1_253/A NOR3X1_13/C NOR3X1_253/C NOR3X1_1533/A NOR3X1_515/B NOR3X1_516/B NOR3X1_1007/B NOR3X1_1491/A NOR3X1_1491/B NOR3X1_1008/B NOR3X1_1492/B NOR3X1_315/A NOR3X1_1007/A NOR3X1_315/B NOR3X1_355/A NOR3X1_355/B NOR3X1_316/B NOR3X1_356/B NOR3X1_515/A NOR3X1_995/C NOR3X1_1207/C NOR3X1_996/A NOR3X1_1208/A NOR3X1_996/B NOR3X1_1208/B NOR3X1_233/B NOR3X1_144/A NOR3X1_144/B NOR3X1_143/C NOR3X1_354/A NOR3X1_354/C NOR3X1_1347/C NOR3X1_1348/A NOR3X1_234/A NOR3X1_1348/B NOR3X1_234/C NOR3X1_345/C NOR3X1_346/A NOR3X1_353/B NOR3X1_346/B NOR3X1_1641/B NOR3X1_875/B NOR3X1_1642/A 
+ NOR3X1_876/A NOR3X1_1642/C NOR3X1_876/C NOR3X1_583/A NOR3X1_1225/A NOR3X1_583/C NOR3X1_1225/C NOR3X1_1226/C NOR3X1_374/C NOR3X1_373/A NOR3X1_1490/C NOR3X1_785/A NOR3X1_373/C NOR3X1_785/B NOR3X1_331/A NOR3X1_331/B NOR3X1_786/B NOR3X1_332/B NOR3X1_1489/A NOR3X1_365/A NOR3X1_365/B NOR3X1_1489/C NOR3X1_366/B NOR3X1_881/A NOR3X1_884/C NOR3X1_881/C NOR3X1_584/C NOR3X1_882/C NOR3X1_883/A NOR3X1_883/C NOR3X1_53/A NOR3X1_53/B NOR3X1_165/A NOR3X1_165/C NOR3X1_166/C NOR3X1_1190/C NOR3X1_474/C NOR3X1_351/A NOR3X1_1189/A NOR3X1_351/C NOR3X1_1189/C NOR3X1_473/A NOR3X1_352/C NOR3X1_473/C NOR3X1_54/B NOR3X1_1043/A NOR3X1_994/C NOR3X1_116/C NOR3X1_1043/C NOR3X1_1229/A NOR3X1_1229/C 
+ NOR3X1_47/A NOR3X1_993/A NOR3X1_993/C NOR3X1_1044/C NOR3X1_115/A NOR3X1_1230/C NOR3X1_47/C NOR3X1_115/C NOR3X1_48/C NOR3X1_500/C NOR3X1_1643/C NOR3X1_624/B NOR3X1_623/A NOR3X1_623/B NOR3X1_499/A NOR3X1_1333/A NOR3X1_1005/A NOR3X1_499/C NOR3X1_1333/C NOR3X1_1005/C NOR3X1_333/A NOR3X1_1006/C NOR3X1_333/C NOR3X1_334/C NOR3X1_1334/C NOR3X1_641/A NOR3X1_1531/A NOR3X1_129/A NOR3X1_1644/C NOR3X1_641/B NOR3X1_129/B NOR3X1_1531/C NOR3X1_642/B NOR3X1_130/B NOR3X1_1532/C NOR3X1_1643/A NOR3X1_639/C NOR3X1_291/A NOR3X1_291/C NOR3X1_989/A NOR3X1_292/C NOR3X1_967/B NOR3X1_989/C NOR3X1_968/B NOR3X1_791/A NOR3X1_791/B NOR3X1_137/C NOR3X1_792/B NOR3X1_77/C NOR3X1_138/C NOR3X1_78/C 
+ NOR3X1_357/C NOR3X1_137/A NOR3X1_77/A NOR3X1_358/C NOR3X1_967/A NOR3X1_640/C NOR3X1_357/A NOR3X1_639/A NOR3X1_990/C NOR3X1_459/A NOR3X1_1165/A NOR3X1_459/B NOR3X1_981/A NOR3X1_1165/C NOR3X1_1200/C NOR3X1_981/C NOR3X1_460/B NOR3X1_1166/C NOR3X1_982/C NOR3X1_147/C NOR3X1_148/C NOR3X1_1033/A NOR3X1_1033/C NOR3X1_147/A NOR3X1_1199/A NOR3X1_1199/C NOR3X1_1051/A NOR3X1_64/B NOR3X1_1051/C NOR3X1_1052/C NOR3X1_1034/C NOR3X1_63/A NOR3X1_63/B NOR3X1_1513/A NOR3X1_970/C NOR3X1_1513/C NOR3X1_797/C NOR3X1_847/C NOR3X1_798/C NOR3X1_969/A NOR3X1_848/C NOR3X1_969/C NOR3X1_797/A NOR3X1_847/A NOR3X1_1401/A NOR3X1_244/C NOR3X1_1401/C NOR3X1_594/C NOR3X1_1402/C NOR3X1_243/A NOR3X1_243/C 
+ NOR3X1_593/A NOR3X1_1514/C NOR3X1_593/C NOR3X1_1047/A NOR3X1_1201/A NOR3X1_1201/B NOR3X1_1202/B NOR3X1_787/C NOR3X1_788/C NOR3X1_1494/C NOR3X1_787/A NOR3X1_1493/A NOR3X1_1493/C NOR3X1_304/C NOR3X1_1047/C NOR3X1_303/A NOR3X1_1048/C NOR3X1_303/C NOR3X1_1050/B NOR3X1_289/A NOR3X1_289/C NOR3X1_1167/A NOR3X1_325/A NOR3X1_1360/C NOR3X1_325/C NOR3X1_326/C NOR3X1_1167/B NOR3X1_1359/A NOR3X1_1359/C NOR3X1_1168/B NOR3X1_1049/A NOR3X1_1049/B NOR3X1_290/C NOR3X1_1097/B NOR3X1_1098/B NOR3X1_1097/A NOR3X1_1098/A NOR3X1_1098/C NOR3X1_1411/B NOR3X1_1412/A NOR3X1_1412/C NOR3X1_1417/B NOR3X1_1418/B NOR3X1_1417/A NOR3X1_1411/A NOR3X1_1412/B NOR3X1_1418/A NOR3X1_1418/C NOR3X1_233/A NOR3X1_233/C NOR3X1_130/C 
+ NOR3X1_129/C NOR3X1_1625/A NOR3X1_1625/B NOR3X1_1626/B NOR3X1_469/A NOR3X1_469/B NOR3X1_470/B NOR3X1_1267/B NOR3X1_1268/A NOR3X1_1268/C NOR3X1_1554/A NOR3X1_1554/B NOR3X1_1553/C NOR3X1_1265/B NOR3X1_1266/A NOR3X1_1266/C NOR3X1_1081/C NOR3X1_1082/A NOR3X1_1082/B NOR3X1_873/B NOR3X1_583/B NOR3X1_345/A NOR3X1_345/B NOR3X1_874/B NOR3X1_584/B NOR3X1_395/C NOR3X1_396/A NOR3X1_396/B NOR3X1_137/B NOR3X1_138/A NOR3X1_670/C NOR3X1_669/B NOR3X1_670/A NOR3X1_993/B NOR3X1_367/C NOR3X1_368/C NOR3X1_143/A NOR3X1_143/B NOR3X1_994/B NOR3X1_138/B NOR3X1_1555/C NOR3X1_1556/A NOR3X1_1556/B NOR3X1_1345/B NOR3X1_1346/A NOR3X1_1346/C NOR3X1_917/B NOR3X1_918/B NOR3X1_917/A NOR3X1_594/A NOR3X1_593/B 
+ NOR3X1_594/B NOR3X1_1675/C NOR3X1_1676/A NOR3X1_1676/B NOR3X1_389/B NOR3X1_390/A NOR3X1_390/C NOR3X1_1081/B NOR3X1_1082/C NOR3X1_1011/B NOR3X1_1012/A NOR3X1_1012/C NOR3X1_894/A NOR3X1_894/B NOR3X1_893/C NOR3X1_1070/C NOR3X1_1069/B NOR3X1_1070/A NOR3X1_275/B NOR3X1_276/A NOR3X1_276/C NOR3X1_918/A NOR3X1_918/C NOR3X1_961/B NOR3X1_962/A NOR3X1_589/B NOR3X1_590/A NOR3X1_1261/B NOR3X1_1262/A NOR3X1_1262/C NOR3X1_797/B NOR3X1_798/A NOR3X1_798/B NOR3X1_590/B NOR3X1_962/B NOR3X1_1259/C NOR3X1_1260/A NOR3X1_1260/B NOR3X1_895/B NOR3X1_896/A NOR3X1_896/C NOR3X1_601/B NOR3X1_602/A NOR3X1_602/C NOR3X1_1661/B NOR3X1_1662/A NOR3X1_1662/C NOR3X1_244/A NOR3X1_243/B NOR3X1_604/A NOR3X1_604/C 
+ NOR3X1_603/B NOR3X1_244/B NOR3X1_1214/A NOR3X1_1213/B NOR3X1_1214/B NOR3X1_1085/B NOR3X1_1086/A NOR3X1_1086/C NOR3X1_1031/C NOR3X1_1032/A NOR3X1_1032/B NOR3X1_967/C NOR3X1_968/C NOR3X1_1007/C NOR3X1_1008/C NOR3X1_1194/C NOR3X1_1193/A NOR3X1_1050/C NOR3X1_1193/C NOR3X1_1641/A NOR3X1_641/C NOR3X1_1641/C NOR3X1_642/C NOR3X1_1049/C NOR3X1_1337/A NOR3X1_1207/B NOR3X1_1207/A NOR3X1_1489/B NOR3X1_333/B NOR3X1_1490/B NOR3X1_1337/C NOR3X1_334/B NOR3X1_1051/B NOR3X1_1338/C NOR3X1_1052/B NOR3X1_1530/A NOR3X1_1201/C NOR3X1_1202/A NOR3X1_31/B NOR3X1_331/C NOR3X1_32/A NOR3X1_332/A NOR3X1_1529/B NOR3X1_683/C NOR3X1_684/A NOR3X1_684/B NOR3X1_1685/B NOR3X1_1686/A NOR3X1_573/C NOR3X1_1686/C NOR3X1_574/A 
+ NOR3X1_574/B NOR3X1_147/B NOR3X1_148/B NOR3X1_1491/C NOR3X1_1492/C NOR3X1_683/A NOR3X1_684/C NOR3X1_924/B NOR3X1_923/A NOR3X1_923/B NOR3X1_924/A NOR3X1_924/C NOR3X1_687/A NOR3X1_687/B NOR3X1_688/B NOR3X1_291/B NOR3X1_984/B NOR3X1_292/B NOR3X1_787/B NOR3X1_983/B NOR3X1_788/B NOR3X1_254/B NOR3X1_253/B NOR3X1_53/C NOR3X1_459/C NOR3X1_14/B NOR3X1_365/C NOR3X1_366/C NOR3X1_1167/C NOR3X1_13/B NOR3X1_1168/C NOR3X1_54/C NOR3X1_460/C NOR3X1_1577/C NOR3X1_1578/A NOR3X1_1578/B NOR3X1_522/C NOR3X1_789/B NOR3X1_790/B NOR3X1_357/B NOR3X1_1199/B NOR3X1_358/B NOR3X1_1200/B NOR3X1_884/B NOR3X1_249/B NOR3X1_250/B NOR3X1_521/A NOR3X1_883/B NOR3X1_521/C NOR3X1_1114/B NOR3X1_1113/A 
+ NOR3X1_1113/B NOR3X1_791/C NOR3X1_792/C NOR3X1_1009/B NOR3X1_1010/B NOR3X1_875/A NOR3X1_47/B NOR3X1_875/C NOR3X1_457/B NOR3X1_48/B NOR3X1_458/B NOR3X1_688/C NOR3X1_688/A NOR3X1_39/B NOR3X1_40/B NOR3X1_1114/A NOR3X1_1114/C NOR3X1_201/B NOR3X1_202/A NOR3X1_202/C NOR3X1_201/A NOR3X1_202/B NOR3X1_640/B NOR3X1_1399/B NOR3X1_1400/B NOR3X1_264/C NOR3X1_351/B NOR3X1_352/B NOR3X1_263/C NOR3X1_1531/B NOR3X1_1532/B NOR3X1_639/B NOR3X1_1625/C NOR3X1_1626/A NOR3X1_469/C NOR3X1_470/A NOR3X1_515/C NOR3X1_516/C NOR3X1_289/B NOR3X1_847/B NOR3X1_290/B NOR3X1_848/B NOR3X1_1643/B NOR3X1_1043/B NOR3X1_981/B NOR3X1_982/B NOR3X1_969/B NOR3X1_970/B NOR3X1_1644/B NOR3X1_1044/B NOR3X1_1223/A 
+ NOR3X1_1223/B NOR3X1_1224/B NOR3X1_1225/B NOR3X1_1226/B NOR3X1_989/B NOR3X1_624/C NOR3X1_990/B NOR3X1_134/C NOR3X1_623/C NOR3X1_355/C NOR3X1_356/C NOR3X1_133/A NOR3X1_133/C NOR3X1_63/C NOR3X1_64/C NOR3X1_781/C NOR3X1_782/A NOR3X1_782/B NOR3X1_513/B NOR3X1_267/B NOR3X1_268/B NOR3X1_1351/C NOR3X1_1352/A NOR3X1_1352/B NOR3X1_1047/B NOR3X1_1048/B NOR3X1_514/B NOR3X1_1518/C NOR3X1_1517/A NOR3X1_474/B NOR3X1_1401/B NOR3X1_473/B NOR3X1_1402/B NOR3X1_1517/C NOR3X1_77/B NOR3X1_785/C NOR3X1_78/B NOR3X1_786/C NOR3X1_120/C NOR3X1_119/C NOR3X1_161/B NOR3X1_162/B NOR3X1_165/B NOR3X1_794/A NOR3X1_166/A NOR3X1_793/B NOR3X1_1165/B NOR3X1_1166/B NOR3X1_1205/B NOR3X1_1206/B NOR3X1_1494/B 
+ NOR3X1_1493/B NOR3X1_881/B NOR3X1_353/A NOR3X1_882/B NOR3X1_353/C NOR3X1_1041/B NOR3X1_115/B NOR3X1_1042/B NOR3X1_116/B NOR3X1_667/B NOR3X1_668/A NOR3X1_668/C NOR3X1_1671/B NOR3X1_1672/A NOR3X1_1672/C NOR3X1_480/C NOR3X1_479/B NOR3X1_480/A NOR3X1_166/B NOR3X1_474/A NOR3X1_352/A NOR3X1_1190/A NOR3X1_1190/B NOR3X1_54/A NOR3X1_984/A NOR3X1_1218/A NOR3X1_1218/B NOR3X1_1400/A NOR3X1_1510/A NOR3X1_1510/B NOR3X1_162/A NOR3X1_790/A NOR3X1_874/A NOR3X1_120/A NOR3X1_1226/A NOR3X1_374/A NOR3X1_374/B NOR3X1_786/A NOR3X1_332/C NOR3X1_1490/A NOR3X1_366/A NOR3X1_884/A NOR3X1_584/A NOR3X1_882/A NOR3X1_1202/C NOR3X1_788/A NOR3X1_1494/A NOR3X1_304/A NOR3X1_304/B NOR3X1_1048/A NOR3X1_901/B 
+ NOR3X1_902/A NOR3X1_902/C NOR3X1_901/A NOR3X1_902/B NOR3X1_290/A NOR3X1_326/A NOR3X1_326/B NOR3X1_1168/A NOR3X1_1360/A NOR3X1_1360/B NOR3X1_1050/A NOR3X1_378/A NOR3X1_378/B NOR3X1_268/A NOR3X1_368/A NOR3X1_264/A NOR3X1_1188/A NOR3X1_1188/B NOR3X1_250/A NOR3X1_812/A NOR3X1_812/B NOR3X1_624/A NOR3X1_500/A NOR3X1_1006/A NOR3X1_500/B NOR3X1_1006/B NOR3X1_334/A NOR3X1_1334/A NOR3X1_1644/A NOR3X1_1334/B NOR3X1_642/A NOR3X1_1532/A NOR3X1_130/A NOR3X1_995/A NOR3X1_996/C NOR3X1_1208/C NOR3X1_144/C NOR3X1_354/B NOR3X1_234/B NOR3X1_1348/C NOR3X1_346/C NOR3X1_1347/A NOR3X1_1642/B NOR3X1_876/B NOR3X1_460/A NOR3X1_1166/A NOR3X1_982/A NOR3X1_148/A NOR3X1_1200/A NOR3X1_64/A NOR3X1_1052/A 
+ NOR3X1_1034/A NOR3X1_1034/B NOR3X1_794/B NOR3X1_1534/A NOR3X1_1534/B NOR3X1_1330/A NOR3X1_14/A NOR3X1_32/B NOR3X1_1330/B NOR3X1_254/A NOR3X1_1530/B NOR3X1_988/A NOR3X1_988/B NOR3X1_1206/A NOR3X1_262/A NOR3X1_262/B NOR3X1_1355/A NOR3X1_1356/C NOR3X1_458/A NOR3X1_1230/A NOR3X1_1230/B NOR3X1_1044/A NOR3X1_48/A NOR3X1_994/A NOR3X1_116/A NOR3X1_1275/A NOR3X1_1275/C NOR3X1_1276/C NOR3X1_516/A NOR3X1_1008/A NOR3X1_1492/A NOR3X1_316/A NOR3X1_356/A NOR3X1_316/C NOR3X1_640/A NOR3X1_292/A NOR3X1_968/A NOR3X1_990/A NOR3X1_792/A NOR3X1_78/A NOR3X1_358/A NOR3X1_848/A NOR3X1_970/A NOR3X1_1402/A NOR3X1_1514/A NOR3X1_1514/B NOR3X1_40/A NOR3X1_158/A NOR3X1_158/B NOR3X1_1332/A NOR3X1_1332/B 
+ NOR3X1_1010/A NOR3X1_514/A NOR3X1_1042/A NOR3X1_920/C NOR3X1_919/B NOR3X1_920/A NOR3X1_919/A NOR3X1_920/B NOR3X1_1269/A NOR3X1_1270/B NOR3X1_1537/C NOR3X1_1538/C NOR3X1_1537/A NOR3X1_1579/A NOR3X1_1580/C NOR3X1_899/C NOR3X1_900/A NOR3X1_900/B NOR3X1_1414/C NOR3X1_1413/A NOR3X1_1413/C NOR3X1_1414/A NOR3X1_1414/B NOR3X1_900/C NOR3X1_899/A NOR3X1_777/B NOR3X1_778/A NOR3X1_778/C NOR3X1_778/B NOR3X1_777/A NOR3X1_709/C NOR3X1_710/A NOR3X1_710/B NOR3X1_1194/A NOR3X1_1193/B NOR3X1_1194/B NOR3X1_895/C NOR3X1_896/B NOR3X1_710/C NOR3X1_709/A NOR3X1_895/A NOR3X1_1268/B NOR3X1_1267/A NOR3X1_470/C NOR3X1_1626/C NOR3X1_1265/A NOR3X1_1266/B NOR3X1_1554/C NOR3X1_1553/A NOR3X1_1081/A NOR3X1_1555/A 
+ NOR3X1_1556/C NOR3X1_1338/A NOR3X1_1338/B NOR3X1_1518/A NOR3X1_1518/B NOR3X1_669/A NOR3X1_670/B NOR3X1_395/A NOR3X1_396/C NOR3X1_1224/C NOR3X1_1224/A NOR3X1_134/A NOR3X1_134/B NOR3X1_1244/A NOR3X1_1244/B NOR3X1_1243/C NOR3X1_1351/A NOR3X1_1352/C NOR3X1_522/A NOR3X1_522/B NOR3X1_1244/C NOR3X1_1243/A NOR3X1_781/A NOR3X1_782/C NOR3X1_1345/A NOR3X1_1346/B NOR3X1_927/B NOR3X1_928/B NOR3X1_927/A NOR3X1_928/A NOR3X1_928/C NOR3X1_917/C NOR3X1_1276/A NOR3X1_1276/B NOR3X1_649/C NOR3X1_650/A NOR3X1_650/B NOR3X1_1005/B NOR3X1_1551/C NOR3X1_1552/A NOR3X1_1552/B NOR3X1_335/C NOR3X1_336/A NOR3X1_336/B NOR3X1_615/C NOR3X1_616/A NOR3X1_616/B NOR3X1_1415/C NOR3X1_1416/A NOR3X1_1416/B NOR3X1_294/C 
+ NOR3X1_293/B NOR3X1_294/A NOR3X1_665/B NOR3X1_666/A NOR3X1_666/C NOR3X1_572/A NOR3X1_572/B NOR3X1_571/C NOR3X1_1407/B NOR3X1_1408/A NOR3X1_891/C NOR3X1_1408/C NOR3X1_892/A NOR3X1_892/B NOR3X1_669/C NOR3X1_453/B NOR3X1_454/A NOR3X1_454/C NOR3X1_650/C NOR3X1_649/A NOR3X1_1551/A NOR3X1_1552/C NOR3X1_335/A NOR3X1_336/C NOR3X1_615/A NOR3X1_616/C NOR3X1_293/A NOR3X1_294/B NOR3X1_1415/A NOR3X1_1416/C NOR3X1_811/B NOR3X1_1039/B NOR3X1_1040/A NOR3X1_1040/C NOR3X1_1351/B NOR3X1_391/B NOR3X1_392/A NOR3X1_392/C NOR3X1_1667/C NOR3X1_1668/A NOR3X1_1668/B NOR3X1_1557/C NOR3X1_1558/A NOR3X1_1558/B NOR3X1_1411/C NOR3X1_1538/A NOR3X1_1538/B NOR3X1_1675/A NOR3X1_1676/C NOR3X1_1069/A NOR3X1_1070/B 
+ NOR3X1_1011/A NOR3X1_1012/B NOR3X1_894/C NOR3X1_893/A NOR3X1_389/A NOR3X1_390/B NOR3X1_275/A NOR3X1_276/B NOR3X1_1696/B NOR3X1_1695/A NOR3X1_1695/B NOR3X1_1696/A NOR3X1_1696/C NOR3X1_1040/B NOR3X1_1039/A NOR3X1_391/A NOR3X1_392/B NOR3X1_1668/C NOR3X1_1558/C NOR3X1_1557/A NOR3X1_1667/A NOR3X1_1577/A NOR3X1_1578/C NOR3X1_1559/C NOR3X1_1560/A NOR3X1_1560/B NOR3X1_1661/C NOR3X1_1662/B NOR3X1_1664/A NOR3X1_1664/C NOR3X1_1663/B NOR3X1_1260/C NOR3X1_1259/A NOR3X1_1685/A NOR3X1_573/A NOR3X1_1686/B NOR3X1_574/C NOR3X1_1085/A NOR3X1_1086/B NOR3X1_604/B NOR3X1_603/A NOR3X1_601/A NOR3X1_602/B NOR3X1_1661/A NOR3X1_1560/C NOR3X1_1559/A NOR3X1_1664/B NOR3X1_1663/A NOR3X1_453/A NOR3X1_454/B NOR3X1_891/A 
+ NOR3X1_1408/B NOR3X1_892/C NOR3X1_1407/A NOR3X1_665/A NOR3X1_666/B NOR3X1_572/C NOR3X1_571/A NOR3X1_1261/A NOR3X1_1262/B NOR3X1_1617/C NOR3X1_1618/C NOR3X1_1617/A NOR3X1_668/B NOR3X1_667/A NOR3X1_1671/A NOR3X1_1672/B NOR3X1_479/A NOR3X1_480/B NOR3X1_1458/B NOR3X1_1457/A NOR3X1_1710/C NOR3X1_1709/A NOR3X1_1709/C NOR3X1_1457/B NOR3X1_649/B NOR3X1_1094/C NOR3X1_1093/A NOR3X1_1093/C NOR3X1_1094/A NOR3X1_1094/B NOR3X1_664/A NOR3X1_664/B NOR3X1_663/C NOR3X1_664/C NOR3X1_663/A NOR3X1_1031/A NOR3X1_1032/C NOR3X1_1458/C NOR3X1_1710/A NOR3X1_1710/B NOR3X1_1458/A NOR3X1_1031/B NOR3X1_721/A NOR3X1_721/B NOR3X1_722/B NOR3X1_945/A NOR3X1_945/B NOR3X1_946/B NOR3X1_722/A NOR3X1_722/C NOR3X1_946/A 
+ NOR3X1_946/C NOR3X1_1618/A NOR3X1_1618/B INVX1_1198/Y INVX1_1197/Y INVX1_176/Y INVX1_175/Y INVX1_131/Y INVX1_132/Y INVX1_747/Y INVX1_748/Y INVX1_239/Y INVX1_240/Y INVX1_653/Y INVX1_654/Y INVX1_1198/A INVX1_548/A INVX1_547/A INVX1_1197/A INVX1_176/A INVX1_175/A INVX1_822/A INVX1_821/A INVX1_1377/A INVX1_1378/A INVX1_131/A INVX1_132/A INVX1_747/A INVX1_748/A INVX1_1640/A INVX1_1639/A INVX1_239/A INVX1_240/A INVX1_653/A INVX1_654/A INVX1_750/A INVX1_749/A INVX1_1060/A INVX1_1059/A INVX1_369/A INVX1_370/A NOR3X1_175/B NOR3X1_821/B NOR3X1_747/B NOR3X1_653/B INVX1_174/Y INVX1_173/Y INVX1_820/Y INVX1_819/Y INVX1_1520/Y INVX1_1519/Y 
+ INVX1_537/Y INVX1_538/Y INVX1_745/Y INVX1_746/Y INVX1_528/Y INVX1_527/Y INVX1_174/A INVX1_173/A INVX1_820/A INVX1_819/A INVX1_1520/A INVX1_1519/A INVX1_537/A INVX1_539/A INVX1_540/A INVX1_538/A INVX1_745/A INVX1_746/A INVX1_528/A INVX1_527/A NOR3X1_1519/B INVX1_1370/Y INVX1_1372/Y INVX1_1371/Y INVX1_1369/Y INVX1_1370/A INVX1_1372/A INVX1_1371/A INVX1_1369/A NOR3X1_1371/C NOR3X1_1369/B INVX1_1364/Y INVX1_1363/Y INVX1_1366/Y INVX1_1365/Y INVX1_1364/A INVX1_1363/A INVX1_1366/A INVX1_1365/A INVX1_855/Y INVX1_856/Y INVX1_1508/Y INVX1_1507/Y INVX1_376/Y INVX1_375/Y INVX1_372/Y INVX1_1063/Y INVX1_371/Y INVX1_1064/Y INVX1_1327/Y INVX1_1216/Y 
+ INVX1_1215/Y INVX1_1328/Y INVX1_766/Y INVX1_765/Y INVX1_259/Y INVX1_260/Y INVX1_1354/Y INVX1_1353/Y INVX1_156/Y INVX1_155/Y INVX1_311/Y INVX1_312/Y INVX1_498/Y INVX1_497/Y INVX1_1227/Y INVX1_1228/Y INVX1_1179/Y INVX1_1180/Y INVX1_1656/Y INVX1_1655/Y INVX1_1511/Y INVX1_1512/Y INVX1_209/Y INVX1_210/Y INVX1_493/Y INVX1_494/Y INVX1_302/Y INVX1_301/Y INVX1_323/Y INVX1_324/Y INVX1_1062/Y INVX1_1061/Y INVX1_1396/Y INVX1_1395/Y INVX1_524/Y INVX1_523/Y INVX1_580/Y INVX1_579/Y INVX1_610/Y INVX1_609/Y INVX1_236/Y INVX1_235/Y INVX1_393/Y INVX1_394/Y INVX1_992/Y INVX1_991/Y INVX1_1340/Y INVX1_1339/Y INVX1_1673/Y INVX1_1674/Y INVX1_82/Y 
+ INVX1_81/Y INVX1_478/Y INVX1_477/Y INVX1_840/Y INVX1_839/Y INVX1_1065/Y INVX1_1066/Y INVX1_270/Y INVX1_269/Y INVX1_1172/Y INVX1_1171/Y INVX1_965/Y INVX1_966/Y INVX1_192/Y INVX1_191/Y INVX1_1257/Y INVX1_1258/Y INVX1_150/Y INVX1_149/Y INVX1_596/Y INVX1_595/Y INVX1_630/Y INVX1_629/Y INVX1_1335/Y INVX1_1336/Y INVX1_496/Y INVX1_495/Y INVX1_502/Y INVX1_501/Y INVX1_567/Y INVX1_568/Y INVX1_832/Y INVX1_831/Y INVX1_508/Y INVX1_507/Y INVX1_758/Y INVX1_757/Y INVX1_1502/Y INVX1_1501/Y INVX1_520/Y INVX1_519/Y INVX1_977/Y INVX1_978/Y INVX1_197/Y INVX1_198/Y INVX1_1219/Y INVX1_1220/Y INVX1_768/Y INVX1_767/Y INVX1_1516/Y INVX1_1515/Y 
+ INVX1_1646/Y INVX1_1645/Y INVX1_463/Y INVX1_464/Y INVX1_1274/Y INVX1_1273/Y INVX1_759/Y INVX1_760/Y INVX1_1528/Y INVX1_1527/Y INVX1_103/Y INVX1_104/Y INVX1_854/Y INVX1_853/Y INVX1_1390/Y INVX1_1389/Y INVX1_770/Y INVX1_769/Y INVX1_662/Y INVX1_661/Y INVX1_1241/Y INVX1_1242/Y INVX1_913/Y INVX1_914/Y INVX1_476/Y INVX1_475/Y INVX1_330/Y INVX1_329/Y INVX1_613/Y INVX1_614/Y INVX1_1394/Y INVX1_1393/Y INVX1_283/Y INVX1_284/Y INVX1_342/Y INVX1_341/Y INVX1_569/Y INVX1_570/Y INVX1_626/Y INVX1_625/Y INVX1_836/Y INVX1_835/Y INVX1_974/Y INVX1_973/Y INVX1_448/Y INVX1_447/Y INVX1_1036/Y INVX1_1035/Y INVX1_90/Y INVX1_89/Y INVX1_1691/Y 
+ INVX1_1692/Y INVX1_308/Y INVX1_307/Y INVX1_1488/Y INVX1_1487/Y INVX1_864/Y INVX1_846/Y INVX1_845/Y INVX1_863/Y INVX1_1603/Y INVX1_1604/Y INVX1_1658/Y INVX1_1657/Y INVX1_1056/Y INVX1_1055/Y INVX1_218/Y INVX1_217/Y INVX1_534/Y INVX1_533/Y INVX1_232/Y INVX1_231/Y INVX1_855/A INVX1_856/A INVX1_1508/A INVX1_1507/A INVX1_376/A INVX1_375/A INVX1_372/A INVX1_1063/A INVX1_371/A INVX1_1064/A INVX1_1327/A INVX1_1216/A INVX1_1215/A INVX1_1328/A INVX1_766/A INVX1_765/A INVX1_259/A INVX1_260/A INVX1_1354/A INVX1_1353/A INVX1_156/A INVX1_155/A INVX1_311/A INVX1_312/A INVX1_498/A INVX1_497/A INVX1_1227/A INVX1_1228/A INVX1_1179/A INVX1_1180/A 
+ INVX1_1656/A INVX1_1655/A INVX1_1511/A INVX1_1512/A INVX1_209/A INVX1_210/A INVX1_493/A INVX1_494/A INVX1_302/A INVX1_301/A INVX1_323/A INVX1_324/A INVX1_1062/A INVX1_1061/A INVX1_1396/A INVX1_1395/A INVX1_524/A INVX1_523/A INVX1_580/A INVX1_579/A INVX1_610/A INVX1_609/A INVX1_236/A INVX1_235/A INVX1_393/A INVX1_394/A INVX1_992/A INVX1_991/A INVX1_1340/A INVX1_1339/A INVX1_1673/A INVX1_1674/A INVX1_82/A INVX1_81/A INVX1_478/A INVX1_477/A INVX1_840/A INVX1_839/A INVX1_1065/A INVX1_1066/A INVX1_270/A INVX1_269/A INVX1_1172/A INVX1_1171/A INVX1_965/A INVX1_966/A INVX1_192/A INVX1_191/A INVX1_1257/A INVX1_1258/A INVX1_150/A 
+ INVX1_149/A INVX1_596/A INVX1_595/A INVX1_630/A INVX1_629/A INVX1_1335/A INVX1_1336/A INVX1_496/A INVX1_495/A INVX1_502/A INVX1_501/A INVX1_567/A INVX1_568/A INVX1_832/A INVX1_831/A INVX1_508/A INVX1_507/A INVX1_758/A INVX1_757/A INVX1_1502/A INVX1_1501/A INVX1_520/A INVX1_519/A INVX1_977/A INVX1_978/A INVX1_197/A INVX1_198/A INVX1_1219/A INVX1_1220/A INVX1_768/A INVX1_767/A INVX1_1516/A INVX1_1515/A INVX1_1646/A INVX1_1645/A INVX1_463/A INVX1_464/A INVX1_1274/A INVX1_1273/A INVX1_759/A INVX1_760/A INVX1_1528/A INVX1_1527/A INVX1_103/A INVX1_104/A INVX1_854/A INVX1_853/A INVX1_1390/A INVX1_1389/A INVX1_770/A INVX1_769/A 
+ INVX1_662/A INVX1_661/A INVX1_1241/A INVX1_1242/A INVX1_913/A INVX1_914/A INVX1_476/A INVX1_475/A INVX1_330/A INVX1_329/A INVX1_613/A INVX1_614/A INVX1_1394/A INVX1_1393/A INVX1_283/A INVX1_284/A INVX1_342/A INVX1_341/A INVX1_569/A INVX1_570/A INVX1_626/A INVX1_625/A INVX1_836/A INVX1_835/A INVX1_974/A INVX1_973/A INVX1_448/A INVX1_447/A INVX1_1036/A INVX1_1035/A INVX1_90/A INVX1_89/A INVX1_1691/A INVX1_1692/A INVX1_308/A INVX1_307/A INVX1_1488/A INVX1_1487/A INVX1_864/A INVX1_846/A INVX1_845/A INVX1_863/A INVX1_1603/A INVX1_1604/A INVX1_1658/A INVX1_1657/A INVX1_1056/A INVX1_1055/A INVX1_218/A INVX1_217/A INVX1_534/A 
+ INVX1_533/A NOR3X1_1507/B NOR3X1_375/B NOR3X1_371/B NOR3X1_311/C NOR3X1_393/C NOR3X1_1065/B NOR3X1_495/B NOR3X1_501/B NOR3X1_977/C NOR3X1_197/C NOR3X1_767/B NOR3X1_1273/B NOR3X1_759/B NOR3X1_613/B NOR3X1_1603/A NOR3X1_1603/B NOR3X1_1603/C NOR3X1_1604/A NOR3X1_1604/B NOR3X1_1604/C NOR3X1_1657/B NOR3X1_232/A NOR3X1_232/B NOR3X1_232/C NOR3X1_231/A NOR3X1_231/B NOR3X1_231/C INVX1_320/Y INVX1_322/Y INVX1_321/Y INVX1_319/Y INVX1_1649/Y INVX1_1651/Y INVX1_1652/Y INVX1_1650/Y INVX1_503/Y INVX1_963/Y INVX1_964/Y INVX1_504/Y INVX1_1251/Y INVX1_1253/Y INVX1_1254/Y INVX1_1252/Y INVX1_557/Y INVX1_559/Y INVX1_560/Y INVX1_558/Y INVX1_506/Y INVX1_505/Y INVX1_194/Y 
+ INVX1_196/Y INVX1_195/Y INVX1_193/Y INVX1_660/Y INVX1_659/Y INVX1_1231/Y INVX1_1233/Y INVX1_1234/Y INVX1_1232/Y INVX1_735/Y INVX1_740/Y INVX1_739/Y INVX1_736/Y INVX1_561/Y INVX1_563/Y INVX1_564/Y INVX1_562/Y INVX1_1629/Y INVX1_1631/Y INVX1_1632/Y INVX1_1630/Y INVX1_1596/Y INVX1_1598/Y INVX1_1597/Y INVX1_1595/Y INVX1_531/Y INVX1_530/Y INVX1_532/Y INVX1_529/Y INVX1_229/Y INVX1_227/Y INVX1_230/Y INVX1_228/Y INVX1_320/A INVX1_322/A INVX1_321/A INVX1_319/A INVX1_1649/A INVX1_1651/A INVX1_1652/A INVX1_1650/A INVX1_503/A INVX1_963/A INVX1_964/A INVX1_504/A INVX1_1251/A INVX1_1253/A INVX1_1254/A INVX1_1252/A INVX1_557/A INVX1_559/A 
+ INVX1_560/A INVX1_558/A INVX1_506/A INVX1_505/A INVX1_194/A INVX1_196/A INVX1_195/A INVX1_193/A INVX1_660/A INVX1_659/A INVX1_1231/A INVX1_1233/A INVX1_1234/A INVX1_1232/A INVX1_735/A INVX1_740/A INVX1_739/A INVX1_736/A INVX1_561/A INVX1_563/A INVX1_564/A INVX1_562/A INVX1_1629/A INVX1_1631/A INVX1_1632/A INVX1_1630/A INVX1_531/A INVX1_530/A INVX1_532/A INVX1_529/A INVX1_229/A INVX1_227/A INVX1_230/A INVX1_228/A NOR3X1_195/B NOR3X1_735/B NOR3X1_1631/B NOR3X1_1596/A NOR3X1_1596/B NOR3X1_1596/C NOR3X1_1598/A NOR3X1_1598/B NOR3X1_1598/C NOR3X1_1597/A NOR3X1_1597/B NOR3X1_1595/A NOR3X1_1595/B NOR3X1_531/C NOR3X1_529/B NOR3X1_227/B INVX1_182/Y 
+ INVX1_178/Y INVX1_181/Y INVX1_177/Y INVX1_871/Y INVX1_637/Y INVX1_872/Y INVX1_638/Y INVX1_1185/Y INVX1_1077/Y INVX1_1186/Y INVX1_1078/Y INVX1_211/Y INVX1_224/Y INVX1_223/Y INVX1_212/Y INVX1_215/Y INVX1_226/Y INVX1_225/Y INVX1_216/Y INVX1_182/A INVX1_178/A INVX1_181/A INVX1_177/A INVX1_871/A INVX1_872/A INVX1_1185/A INVX1_1186/A INVX1_211/A INVX1_224/A INVX1_223/A INVX1_212/A INVX1_215/A INVX1_226/A INVX1_225/A INVX1_216/A NOR3X1_871/C NOR3X1_637/A NOR3X1_637/B NOR3X1_637/C NOR3X1_638/A NOR3X1_638/B NOR3X1_638/C NOR3X1_1185/B NOR3X1_1077/A NOR3X1_1077/B NOR3X1_1077/C NOR3X1_1078/A NOR3X1_1078/B NOR3X1_1078/C NOR3X1_211/B NOR3X1_223/C 
+ INVX1_868/Y INVX1_870/Y INVX1_869/Y INVX1_867/Y INVX1_634/Y INVX1_636/Y INVX1_635/Y INVX1_633/Y INVX1_1181/Y INVX1_1184/Y INVX1_1183/Y INVX1_1182/Y INVX1_1074/Y INVX1_1076/Y INVX1_1075/Y INVX1_1073/Y INVX1_214/Y INVX1_206/Y INVX1_213/Y INVX1_205/Y INVX1_868/A INVX1_870/A INVX1_869/A INVX1_867/A INVX1_634/A INVX1_636/A INVX1_635/A INVX1_633/A INVX1_1181/A INVX1_1184/A INVX1_1183/A INVX1_1182/A INVX1_1074/A INVX1_1076/A INVX1_1075/A INVX1_1073/A INVX1_214/A INVX1_206/A INVX1_213/A INVX1_205/A NOR3X1_869/C NOR3X1_1181/B INVX1_862/Y INVX1_344/Y INVX1_861/Y INVX1_343/Y INVX1_628/Y INVX1_627/Y INVX1_632/Y INVX1_631/Y INVX1_1178/Y 
+ INVX1_1177/Y INVX1_1072/Y INVX1_1071/Y INVX1_622/Y INVX1_26/Y INVX1_621/Y INVX1_25/Y INVX1_862/A INVX1_344/A INVX1_861/A INVX1_343/A INVX1_628/A INVX1_627/A INVX1_632/A INVX1_631/A INVX1_1178/A INVX1_1177/A INVX1_1072/A INVX1_1071/A INVX1_622/A INVX1_26/A INVX1_621/A INVX1_25/A INVX1_370/Y INVX1_369/Y INVX1_540/Y INVX1_539/Y INVX1_1374/Y INVX1_1373/Y 
+ AES_SBOX_1

.include outputs_0.plw

* **************************************
* --- Simulation Settings ---
* **************************************

.param SIM_LEN = 50ns
.csparam SIM_LEN = {SIM_LEN}

.tran 0.1ns 'SIM_LEN'
.param SIMSTEP = 'SIM_LEN/0.1ns'
.csparam SIMSTEP = {SIMSTEP}

* **************************************
* --- Simulation Control ---
* **************************************

.control
    .include ../inputsD.inc

    run
    
    if ('writeFile' > 0)   
      wrdata ivdd_1.out i(vvdd)
      wrdata ivss_1.out i(vvss)
      *snsave sim_1.snap
    end
    
    set wr_vecnames
    set wr_singlescale
    wrdata outputs_1.out V("NOR3X1_1270/C") V("NOR3X1_1269/B") V("NOR3X1_1270/A") V("NOR3X1_1579/C") V("NOR3X1_1580/A") V("NOR3X1_1580/B") V("NOR3X1_377/C") V("NOR3X1_367/B") V("NOR3X1_267/C") V("NOR3X1_378/C") V("NOR3X1_368/B") V("NOR3X1_268/C") V("NOR3X1_377/A") V("NOR3X1_264/B") V("NOR3X1_1187/C") V("NOR3X1_250/C") V("NOR3X1_1188/C") V("NOR3X1_263/A") V("NOR3X1_263/B") V("NOR3X1_267/A") V("NOR3X1_367/A") V("NOR3X1_249/A") V("NOR3X1_1187/A") V("NOR3X1_249/C") V("NOR3X1_811/A") V("NOR3X1_811/C") V("NOR3X1_812/C") V("NOR3X1_120/B") V("NOR3X1_873/C") V("NOR3X1_1217/C") V("NOR3X1_984/C") V("NOR3X1_1399/A") V("NOR3X1_1509/A") V("NOR3X1_1218/C") V("NOR3X1_1399/C") V("NOR3X1_161/A") V("NOR3X1_1509/C") V("NOR3X1_161/C") V("NOR3X1_790/C") V("NOR3X1_983/A") V("NOR3X1_1217/A") V("NOR3X1_162/C") V("NOR3X1_983/C") V("NOR3X1_789/A") V("NOR3X1_789/C") V("NOR3X1_1400/C") V("NOR3X1_590/C") V("NOR3X1_874/C") V("NOR3X1_589/A") V("NOR3X1_119/A") V("NOR3X1_119/B") V("NOR3X1_1510/C") V("NOR3X1_589/C") V("NOR3X1_873/A") V("NOR3X1_1529/C") V("NOR3X1_458/C") V("NOR3X1_987/C") V("NOR3X1_988/C") V("NOR3X1_457/A") V("NOR3X1_1205/A") V("NOR3X1_1205/C") V("NOR3X1_987/A") V("NOR3X1_1206/C") V("NOR3X1_261/A") V("NOR3X1_261/C") V("NOR3X1_262/C") V("NOR3X1_1355/C") V("NOR3X1_1356/A") V("NOR3X1_1356/B") V("NOR3X1_1530/C") V("NOR3X1_457/C") V("NOR3X1_1529/A") V("NOR3X1_1214/C") V("NOR3X1_39/A") V("NOR3X1_513/A") V("NOR3X1_39/C") V("NOR3X1_513/C") V("NOR3X1_157/C") V("NOR3X1_1213/A") V("NOR3X1_158/C") V("NOR3X1_1331/A") V("NOR3X1_1213/C") V("NOR3X1_1010/C") V("NOR3X1_1331/C") V("NOR3X1_1332/C") V("NOR3X1_157/A") V("NOR3X1_1009/A") V("NOR3X1_1009/C") V("NOR3X1_1041/A") V("NOR3X1_1041/C") V("NOR3X1_40/C") V("NOR3X1_514/C") V("NOR3X1_1042/C") V("NOR3X1_1533/C") V("NOR3X1_1330/C") V("NOR3X1_794/C") V("NOR3X1_31/A") V("NOR3X1_1329/A") V("NOR3X1_793/A") V("NOR3X1_31/C") V("NOR3X1_1329/C") V("NOR3X1_793/C") V("NOR3X1_961/A") V("NOR3X1_1534/C") V("NOR3X1_32/C") V("NOR3X1_14/C") V("NOR3X1_961/C") V("NOR3X1_254/C") V("NOR3X1_962/C") V("NOR3X1_13/A") V("NOR3X1_253/A") V("NOR3X1_13/C") V("NOR3X1_253/C") V("NOR3X1_1533/A") V("NOR3X1_515/B") V("NOR3X1_516/B") V("NOR3X1_1007/B") V("NOR3X1_1491/A") V("NOR3X1_1491/B") V("NOR3X1_1008/B") V("NOR3X1_1492/B") V("NOR3X1_315/A") V("NOR3X1_1007/A") V("NOR3X1_315/B") V("NOR3X1_355/A") V("NOR3X1_355/B") V("NOR3X1_316/B") V("NOR3X1_356/B") V("NOR3X1_515/A") V("NOR3X1_995/C") V("NOR3X1_1207/C") V("NOR3X1_996/A") V("NOR3X1_1208/A") V("NOR3X1_996/B") V("NOR3X1_1208/B") V("NOR3X1_233/B") V("NOR3X1_144/A") V("NOR3X1_144/B") V("NOR3X1_143/C") V("NOR3X1_354/A") V("NOR3X1_354/C") V("NOR3X1_1347/C") V("NOR3X1_1348/A") V("NOR3X1_234/A") V("NOR3X1_1348/B") V("NOR3X1_234/C") V("NOR3X1_345/C") V("NOR3X1_346/A") V("NOR3X1_353/B") V("NOR3X1_346/B") V("NOR3X1_1641/B") V("NOR3X1_875/B") V("NOR3X1_1642/A") V("NOR3X1_876/A") V("NOR3X1_1642/C") V("NOR3X1_876/C") V("NOR3X1_583/A") V("NOR3X1_1225/A") V("NOR3X1_583/C") V("NOR3X1_1225/C") V("NOR3X1_1226/C") V("NOR3X1_374/C") V("NOR3X1_373/A") V("NOR3X1_1490/C") V("NOR3X1_785/A") V("NOR3X1_373/C") V("NOR3X1_785/B") V("NOR3X1_331/A") V("NOR3X1_331/B") V("NOR3X1_786/B") V("NOR3X1_332/B") V("NOR3X1_1489/A") V("NOR3X1_365/A") V("NOR3X1_365/B") V("NOR3X1_1489/C") V("NOR3X1_366/B") V("NOR3X1_881/A") V("NOR3X1_884/C") V("NOR3X1_881/C") V("NOR3X1_584/C") V("NOR3X1_882/C") V("NOR3X1_883/A") V("NOR3X1_883/C") V("NOR3X1_53/A") V("NOR3X1_53/B") V("NOR3X1_165/A") V("NOR3X1_165/C") V("NOR3X1_166/C") V("NOR3X1_1190/C") V("NOR3X1_474/C") V("NOR3X1_351/A") V("NOR3X1_1189/A") V("NOR3X1_351/C") V("NOR3X1_1189/C") V("NOR3X1_473/A") V("NOR3X1_352/C") V("NOR3X1_473/C") V("NOR3X1_54/B") V("NOR3X1_1043/A") V("NOR3X1_994/C") V("NOR3X1_116/C") V("NOR3X1_1043/C") V("NOR3X1_1229/A") V("NOR3X1_1229/C") V("NOR3X1_47/A") V("NOR3X1_993/A") V("NOR3X1_993/C") V("NOR3X1_1044/C") V("NOR3X1_115/A") V("NOR3X1_1230/C") V("NOR3X1_47/C") V("NOR3X1_115/C") V("NOR3X1_48/C") V("NOR3X1_500/C") V("NOR3X1_1643/C") V("NOR3X1_624/B") V("NOR3X1_623/A") V("NOR3X1_623/B") V("NOR3X1_499/A") V("NOR3X1_1333/A") V("NOR3X1_1005/A") V("NOR3X1_499/C") V("NOR3X1_1333/C") V("NOR3X1_1005/C") V("NOR3X1_333/A") V("NOR3X1_1006/C") V("NOR3X1_333/C") V("NOR3X1_334/C") V("NOR3X1_1334/C") V("NOR3X1_641/A") V("NOR3X1_1531/A") V("NOR3X1_129/A") V("NOR3X1_1644/C") V("NOR3X1_641/B") V("NOR3X1_129/B") V("NOR3X1_1531/C") V("NOR3X1_642/B") V("NOR3X1_130/B") V("NOR3X1_1532/C") V("NOR3X1_1643/A") V("NOR3X1_639/C") V("NOR3X1_291/A") V("NOR3X1_291/C") V("NOR3X1_989/A") V("NOR3X1_292/C") V("NOR3X1_967/B") V("NOR3X1_989/C") V("NOR3X1_968/B") V("NOR3X1_791/A") V("NOR3X1_791/B") V("NOR3X1_137/C") V("NOR3X1_792/B") V("NOR3X1_77/C") V("NOR3X1_138/C") V("NOR3X1_78/C") V("NOR3X1_357/C") V("NOR3X1_137/A") V("NOR3X1_77/A") V("NOR3X1_358/C") V("NOR3X1_967/A") V("NOR3X1_640/C") V("NOR3X1_357/A") V("NOR3X1_639/A") V("NOR3X1_990/C") V("NOR3X1_459/A") V("NOR3X1_1165/A") V("NOR3X1_459/B") V("NOR3X1_981/A") V("NOR3X1_1165/C") V("NOR3X1_1200/C") V("NOR3X1_981/C") V("NOR3X1_460/B") V("NOR3X1_1166/C") V("NOR3X1_982/C") V("NOR3X1_147/C") V("NOR3X1_148/C") V("NOR3X1_1033/A") V("NOR3X1_1033/C") V("NOR3X1_147/A") V("NOR3X1_1199/A") V("NOR3X1_1199/C") V("NOR3X1_1051/A") V("NOR3X1_64/B") V("NOR3X1_1051/C") V("NOR3X1_1052/C") V("NOR3X1_1034/C") V("NOR3X1_63/A") V("NOR3X1_63/B") V("NOR3X1_1513/A") V("NOR3X1_970/C") V("NOR3X1_1513/C") V("NOR3X1_797/C") V("NOR3X1_847/C") V("NOR3X1_798/C") V("NOR3X1_969/A") V("NOR3X1_848/C") V("NOR3X1_969/C") V("NOR3X1_797/A") V("NOR3X1_847/A") V("NOR3X1_1401/A") V("NOR3X1_244/C") V("NOR3X1_1401/C") V("NOR3X1_594/C") V("NOR3X1_1402/C") V("NOR3X1_243/A") V("NOR3X1_243/C") V("NOR3X1_593/A") V("NOR3X1_1514/C") V("NOR3X1_593/C") V("NOR3X1_1047/A") V("NOR3X1_1201/A") V("NOR3X1_1201/B") V("NOR3X1_1202/B") V("NOR3X1_787/C") V("NOR3X1_788/C") V("NOR3X1_1494/C") V("NOR3X1_787/A") V("NOR3X1_1493/A") V("NOR3X1_1493/C") V("NOR3X1_304/C") V("NOR3X1_1047/C") V("NOR3X1_303/A") V("NOR3X1_1048/C") V("NOR3X1_303/C") V("NOR3X1_1050/B") V("NOR3X1_289/A") V("NOR3X1_289/C") V("NOR3X1_1167/A") V("NOR3X1_325/A") V("NOR3X1_1360/C") V("NOR3X1_325/C") V("NOR3X1_326/C") V("NOR3X1_1167/B") V("NOR3X1_1359/A") V("NOR3X1_1359/C") V("NOR3X1_1168/B") V("NOR3X1_1049/A") V("NOR3X1_1049/B") V("NOR3X1_290/C") V("NOR3X1_1097/B") V("NOR3X1_1098/B") V("NOR3X1_1097/A") V("NOR3X1_1098/A") V("NOR3X1_1098/C") V("NOR3X1_1411/B") V("NOR3X1_1412/A") V("NOR3X1_1412/C") V("NOR3X1_1417/B") V("NOR3X1_1418/B") V("NOR3X1_1417/A") V("NOR3X1_1411/A") V("NOR3X1_1412/B") V("NOR3X1_1418/A") V("NOR3X1_1418/C") V("NOR3X1_233/A") V("NOR3X1_233/C") V("NOR3X1_130/C") V("NOR3X1_129/C") V("NOR3X1_1625/A") V("NOR3X1_1625/B") V("NOR3X1_1626/B") V("NOR3X1_469/A") V("NOR3X1_469/B") V("NOR3X1_470/B") V("NOR3X1_1267/B") V("NOR3X1_1268/A") V("NOR3X1_1268/C") V("NOR3X1_1554/A") V("NOR3X1_1554/B") V("NOR3X1_1553/C") V("NOR3X1_1265/B") V("NOR3X1_1266/A") V("NOR3X1_1266/C") V("NOR3X1_1081/C") V("NOR3X1_1082/A") V("NOR3X1_1082/B") V("NOR3X1_873/B") V("NOR3X1_583/B") V("NOR3X1_345/A") V("NOR3X1_345/B") V("NOR3X1_874/B") V("NOR3X1_584/B") V("NOR3X1_395/C") V("NOR3X1_396/A") V("NOR3X1_396/B") V("NOR3X1_137/B") V("NOR3X1_138/A") V("NOR3X1_670/C") V("NOR3X1_669/B") V("NOR3X1_670/A") V("NOR3X1_993/B") V("NOR3X1_367/C") V("NOR3X1_368/C") V("NOR3X1_143/A") V("NOR3X1_143/B") V("NOR3X1_994/B") V("NOR3X1_138/B") V("NOR3X1_1555/C") V("NOR3X1_1556/A") V("NOR3X1_1556/B") V("NOR3X1_1345/B") V("NOR3X1_1346/A") V("NOR3X1_1346/C") V("NOR3X1_917/B") V("NOR3X1_918/B") V("NOR3X1_917/A") V("NOR3X1_594/A") V("NOR3X1_593/B") V("NOR3X1_594/B") V("NOR3X1_1675/C") V("NOR3X1_1676/A") V("NOR3X1_1676/B") V("NOR3X1_389/B") V("NOR3X1_390/A") V("NOR3X1_390/C") V("NOR3X1_1081/B") V("NOR3X1_1082/C") V("NOR3X1_1011/B") V("NOR3X1_1012/A") V("NOR3X1_1012/C") V("NOR3X1_894/A") V("NOR3X1_894/B") V("NOR3X1_893/C") V("NOR3X1_1070/C") V("NOR3X1_1069/B") V("NOR3X1_1070/A") V("NOR3X1_275/B") V("NOR3X1_276/A") V("NOR3X1_276/C") V("NOR3X1_918/A") V("NOR3X1_918/C") V("NOR3X1_961/B") V("NOR3X1_962/A") V("NOR3X1_589/B") V("NOR3X1_590/A") V("NOR3X1_1261/B") V("NOR3X1_1262/A") V("NOR3X1_1262/C") V("NOR3X1_797/B") V("NOR3X1_798/A") V("NOR3X1_798/B") V("NOR3X1_590/B") V("NOR3X1_962/B") V("NOR3X1_1259/C") V("NOR3X1_1260/A") V("NOR3X1_1260/B") V("NOR3X1_895/B") V("NOR3X1_896/A") V("NOR3X1_896/C") V("NOR3X1_601/B") V("NOR3X1_602/A") V("NOR3X1_602/C") V("NOR3X1_1661/B") V("NOR3X1_1662/A") V("NOR3X1_1662/C") V("NOR3X1_244/A") V("NOR3X1_243/B") V("NOR3X1_604/A") V("NOR3X1_604/C") V("NOR3X1_603/B") V("NOR3X1_244/B") V("NOR3X1_1214/A") V("NOR3X1_1213/B") V("NOR3X1_1214/B") V("NOR3X1_1085/B") V("NOR3X1_1086/A") V("NOR3X1_1086/C") V("NOR3X1_1031/C") V("NOR3X1_1032/A") V("NOR3X1_1032/B") V("NOR3X1_967/C") V("NOR3X1_968/C") V("NOR3X1_1007/C") V("NOR3X1_1008/C") V("NOR3X1_1194/C") V("NOR3X1_1193/A") V("NOR3X1_1050/C") V("NOR3X1_1193/C") V("NOR3X1_1641/A") V("NOR3X1_641/C") V("NOR3X1_1641/C") V("NOR3X1_642/C") V("NOR3X1_1049/C") V("NOR3X1_1337/A") V("NOR3X1_1207/B") V("NOR3X1_1207/A") V("NOR3X1_1489/B") V("NOR3X1_333/B") V("NOR3X1_1490/B") V("NOR3X1_1337/C") V("NOR3X1_334/B") V("NOR3X1_1051/B") V("NOR3X1_1338/C") V("NOR3X1_1052/B") V("NOR3X1_1530/A") V("NOR3X1_1201/C") V("NOR3X1_1202/A") V("NOR3X1_31/B") V("NOR3X1_331/C") V("NOR3X1_32/A") V("NOR3X1_332/A") V("NOR3X1_1529/B") V("NOR3X1_683/C") V("NOR3X1_684/A") V("NOR3X1_684/B") V("NOR3X1_1685/B") V("NOR3X1_1686/A") V("NOR3X1_573/C") V("NOR3X1_1686/C") V("NOR3X1_574/A") V("NOR3X1_574/B") V("NOR3X1_147/B") V("NOR3X1_148/B") V("NOR3X1_1491/C") V("NOR3X1_1492/C") V("NOR3X1_683/A") V("NOR3X1_684/C") V("NOR3X1_924/B") V("NOR3X1_923/A") V("NOR3X1_923/B") V("NOR3X1_924/A") V("NOR3X1_924/C") V("NOR3X1_687/A") V("NOR3X1_687/B") V("NOR3X1_688/B") V("NOR3X1_291/B") V("NOR3X1_984/B") V("NOR3X1_292/B") V("NOR3X1_787/B") V("NOR3X1_983/B") V("NOR3X1_788/B") V("NOR3X1_254/B") V("NOR3X1_253/B") V("NOR3X1_53/C") V("NOR3X1_459/C") V("NOR3X1_14/B") V("NOR3X1_365/C") V("NOR3X1_366/C") V("NOR3X1_1167/C") V("NOR3X1_13/B") V("NOR3X1_1168/C") V("NOR3X1_54/C") V("NOR3X1_460/C") V("NOR3X1_1577/C") V("NOR3X1_1578/A") V("NOR3X1_1578/B") V("NOR3X1_522/C") V("NOR3X1_789/B") V("NOR3X1_790/B") V("NOR3X1_357/B") V("NOR3X1_1199/B") V("NOR3X1_358/B") V("NOR3X1_1200/B") V("NOR3X1_884/B") V("NOR3X1_249/B") V("NOR3X1_250/B") V("NOR3X1_521/A") V("NOR3X1_883/B") V("NOR3X1_521/C") V("NOR3X1_1114/B") V("NOR3X1_1113/A") V("NOR3X1_1113/B") V("NOR3X1_791/C") V("NOR3X1_792/C") V("NOR3X1_1009/B") V("NOR3X1_1010/B") V("NOR3X1_875/A") V("NOR3X1_47/B") V("NOR3X1_875/C") V("NOR3X1_457/B") V("NOR3X1_48/B") V("NOR3X1_458/B") V("NOR3X1_688/C") V("NOR3X1_688/A") V("NOR3X1_39/B") V("NOR3X1_40/B") V("NOR3X1_1114/A") V("NOR3X1_1114/C") V("NOR3X1_201/B") V("NOR3X1_202/A") V("NOR3X1_202/C") V("NOR3X1_201/A") V("NOR3X1_202/B") V("NOR3X1_640/B") V("NOR3X1_1399/B") V("NOR3X1_1400/B") V("NOR3X1_264/C") V("NOR3X1_351/B") V("NOR3X1_352/B") V("NOR3X1_263/C") V("NOR3X1_1531/B") V("NOR3X1_1532/B") V("NOR3X1_639/B") V("NOR3X1_1625/C") V("NOR3X1_1626/A") V("NOR3X1_469/C") V("NOR3X1_470/A") V("NOR3X1_515/C") V("NOR3X1_516/C") V("NOR3X1_289/B") V("NOR3X1_847/B") V("NOR3X1_290/B") V("NOR3X1_848/B") V("NOR3X1_1643/B") V("NOR3X1_1043/B") V("NOR3X1_981/B") V("NOR3X1_982/B") V("NOR3X1_969/B") V("NOR3X1_970/B") V("NOR3X1_1644/B") V("NOR3X1_1044/B") V("NOR3X1_1223/A") V("NOR3X1_1223/B") V("NOR3X1_1224/B") V("NOR3X1_1225/B") V("NOR3X1_1226/B") V("NOR3X1_989/B") V("NOR3X1_624/C") V("NOR3X1_990/B") V("NOR3X1_134/C") V("NOR3X1_623/C") V("NOR3X1_355/C") V("NOR3X1_356/C") V("NOR3X1_133/A") V("NOR3X1_133/C") V("NOR3X1_63/C") V("NOR3X1_64/C") V("NOR3X1_781/C") V("NOR3X1_782/A") V("NOR3X1_782/B") V("NOR3X1_513/B") V("NOR3X1_267/B") V("NOR3X1_268/B") V("NOR3X1_1351/C") V("NOR3X1_1352/A") V("NOR3X1_1352/B") V("NOR3X1_1047/B") V("NOR3X1_1048/B") V("NOR3X1_514/B") V("NOR3X1_1518/C") V("NOR3X1_1517/A") V("NOR3X1_474/B") V("NOR3X1_1401/B") V("NOR3X1_473/B") V("NOR3X1_1402/B") V("NOR3X1_1517/C") V("NOR3X1_77/B") V("NOR3X1_785/C") V("NOR3X1_78/B") V("NOR3X1_786/C") V("NOR3X1_120/C") V("NOR3X1_119/C") V("NOR3X1_161/B") V("NOR3X1_162/B") V("NOR3X1_165/B") V("NOR3X1_794/A") V("NOR3X1_166/A") V("NOR3X1_793/B") V("NOR3X1_1165/B") V("NOR3X1_1166/B") V("NOR3X1_1205/B") V("NOR3X1_1206/B") V("NOR3X1_1494/B") V("NOR3X1_1493/B") V("NOR3X1_881/B") V("NOR3X1_353/A") V("NOR3X1_882/B") V("NOR3X1_353/C") V("NOR3X1_1041/B") V("NOR3X1_115/B") V("NOR3X1_1042/B") V("NOR3X1_116/B") V("NOR3X1_667/B") V("NOR3X1_668/A") V("NOR3X1_668/C") V("NOR3X1_1671/B") V("NOR3X1_1672/A") V("NOR3X1_1672/C") V("NOR3X1_480/C") V("NOR3X1_479/B") V("NOR3X1_480/A") V("NOR3X1_166/B") V("NOR3X1_474/A") V("NOR3X1_352/A") V("NOR3X1_1190/A") V("NOR3X1_1190/B") V("NOR3X1_54/A") V("NOR3X1_984/A") V("NOR3X1_1218/A") V("NOR3X1_1218/B") V("NOR3X1_1400/A") V("NOR3X1_1510/A") V("NOR3X1_1510/B") V("NOR3X1_162/A") V("NOR3X1_790/A") V("NOR3X1_874/A") V("NOR3X1_120/A") V("NOR3X1_1226/A") V("NOR3X1_374/A") V("NOR3X1_374/B") V("NOR3X1_786/A") V("NOR3X1_332/C") V("NOR3X1_1490/A") V("NOR3X1_366/A") V("NOR3X1_884/A") V("NOR3X1_584/A") V("NOR3X1_882/A") V("NOR3X1_1202/C") V("NOR3X1_788/A") V("NOR3X1_1494/A") V("NOR3X1_304/A") V("NOR3X1_304/B") V("NOR3X1_1048/A") V("NOR3X1_901/B") V("NOR3X1_902/A") V("NOR3X1_902/C") V("NOR3X1_901/A") V("NOR3X1_902/B") V("NOR3X1_290/A") V("NOR3X1_326/A") V("NOR3X1_326/B") V("NOR3X1_1168/A") V("NOR3X1_1360/A") V("NOR3X1_1360/B") V("NOR3X1_1050/A") V("NOR3X1_378/A") V("NOR3X1_378/B") V("NOR3X1_268/A") V("NOR3X1_368/A") V("NOR3X1_264/A") V("NOR3X1_1188/A") V("NOR3X1_1188/B") V("NOR3X1_250/A") V("NOR3X1_812/A") V("NOR3X1_812/B") V("NOR3X1_624/A") V("NOR3X1_500/A") V("NOR3X1_1006/A") V("NOR3X1_500/B") V("NOR3X1_1006/B") V("NOR3X1_334/A") V("NOR3X1_1334/A") V("NOR3X1_1644/A") V("NOR3X1_1334/B") V("NOR3X1_642/A") V("NOR3X1_1532/A") V("NOR3X1_130/A") V("NOR3X1_995/A") V("NOR3X1_996/C") V("NOR3X1_1208/C") V("NOR3X1_144/C") V("NOR3X1_354/B") V("NOR3X1_234/B") V("NOR3X1_1348/C") V("NOR3X1_346/C") V("NOR3X1_1347/A") V("NOR3X1_1642/B") V("NOR3X1_876/B") V("NOR3X1_460/A") V("NOR3X1_1166/A") V("NOR3X1_982/A") V("NOR3X1_148/A") V("NOR3X1_1200/A") V("NOR3X1_64/A") V("NOR3X1_1052/A") V("NOR3X1_1034/A") V("NOR3X1_1034/B") V("NOR3X1_794/B") V("NOR3X1_1534/A") V("NOR3X1_1534/B") V("NOR3X1_1330/A") V("NOR3X1_14/A") V("NOR3X1_32/B") V("NOR3X1_1330/B") V("NOR3X1_254/A") V("NOR3X1_1530/B") V("NOR3X1_988/A") V("NOR3X1_988/B") V("NOR3X1_1206/A") V("NOR3X1_262/A") V("NOR3X1_262/B") V("NOR3X1_1355/A") V("NOR3X1_1356/C") V("NOR3X1_458/A") V("NOR3X1_1230/A") V("NOR3X1_1230/B") V("NOR3X1_1044/A") V("NOR3X1_48/A") V("NOR3X1_994/A") V("NOR3X1_116/A") V("NOR3X1_1275/A") V("NOR3X1_1275/C") V("NOR3X1_1276/C") V("NOR3X1_516/A") V("NOR3X1_1008/A") V("NOR3X1_1492/A") V("NOR3X1_316/A") V("NOR3X1_356/A") V("NOR3X1_316/C") V("NOR3X1_640/A") V("NOR3X1_292/A") V("NOR3X1_968/A") V("NOR3X1_990/A") V("NOR3X1_792/A") V("NOR3X1_78/A") V("NOR3X1_358/A") V("NOR3X1_848/A") V("NOR3X1_970/A") V("NOR3X1_1402/A") V("NOR3X1_1514/A") V("NOR3X1_1514/B") V("NOR3X1_40/A") V("NOR3X1_158/A") V("NOR3X1_158/B") V("NOR3X1_1332/A") V("NOR3X1_1332/B") V("NOR3X1_1010/A") V("NOR3X1_514/A") V("NOR3X1_1042/A") V("NOR3X1_920/C") V("NOR3X1_919/B") V("NOR3X1_920/A") V("NOR3X1_919/A") V("NOR3X1_920/B") V("NOR3X1_1269/A") V("NOR3X1_1270/B") V("NOR3X1_1537/C") V("NOR3X1_1538/C") V("NOR3X1_1537/A") V("NOR3X1_1579/A") V("NOR3X1_1580/C") V("NOR3X1_899/C") V("NOR3X1_900/A") V("NOR3X1_900/B") V("NOR3X1_1414/C") V("NOR3X1_1413/A") V("NOR3X1_1413/C") V("NOR3X1_1414/A") V("NOR3X1_1414/B") V("NOR3X1_900/C") V("NOR3X1_899/A") V("NOR3X1_777/B") V("NOR3X1_778/A") V("NOR3X1_778/C") V("NOR3X1_778/B") V("NOR3X1_777/A") V("NOR3X1_709/C") V("NOR3X1_710/A") V("NOR3X1_710/B") V("NOR3X1_1194/A") V("NOR3X1_1193/B") V("NOR3X1_1194/B") V("NOR3X1_895/C") V("NOR3X1_896/B") V("NOR3X1_710/C") V("NOR3X1_709/A") V("NOR3X1_895/A") V("NOR3X1_1268/B") V("NOR3X1_1267/A") V("NOR3X1_470/C") V("NOR3X1_1626/C") V("NOR3X1_1265/A") V("NOR3X1_1266/B") V("NOR3X1_1554/C") V("NOR3X1_1553/A") V("NOR3X1_1081/A") V("NOR3X1_1555/A") V("NOR3X1_1556/C") V("NOR3X1_1338/A") V("NOR3X1_1338/B") V("NOR3X1_1518/A") V("NOR3X1_1518/B") V("NOR3X1_669/A") V("NOR3X1_670/B") V("NOR3X1_395/A") V("NOR3X1_396/C") V("NOR3X1_1224/C") V("NOR3X1_1224/A") V("NOR3X1_134/A") V("NOR3X1_134/B") V("NOR3X1_1244/A") V("NOR3X1_1244/B") V("NOR3X1_1243/C") V("NOR3X1_1351/A") V("NOR3X1_1352/C") V("NOR3X1_522/A") V("NOR3X1_522/B") V("NOR3X1_1244/C") V("NOR3X1_1243/A") V("NOR3X1_781/A") V("NOR3X1_782/C") V("NOR3X1_1345/A") V("NOR3X1_1346/B") V("NOR3X1_927/B") V("NOR3X1_928/B") V("NOR3X1_927/A") V("NOR3X1_928/A") V("NOR3X1_928/C") V("NOR3X1_917/C") V("NOR3X1_1276/A") V("NOR3X1_1276/B") V("NOR3X1_649/C") V("NOR3X1_650/A") V("NOR3X1_650/B") V("NOR3X1_1005/B") V("NOR3X1_1551/C") V("NOR3X1_1552/A") V("NOR3X1_1552/B") V("NOR3X1_335/C") V("NOR3X1_336/A") V("NOR3X1_336/B") V("NOR3X1_615/C") V("NOR3X1_616/A") V("NOR3X1_616/B") V("NOR3X1_1415/C") V("NOR3X1_1416/A") V("NOR3X1_1416/B") V("NOR3X1_294/C") V("NOR3X1_293/B") V("NOR3X1_294/A") V("NOR3X1_665/B") V("NOR3X1_666/A") V("NOR3X1_666/C") V("NOR3X1_572/A") V("NOR3X1_572/B") V("NOR3X1_571/C") V("NOR3X1_1407/B") V("NOR3X1_1408/A") V("NOR3X1_891/C") V("NOR3X1_1408/C") V("NOR3X1_892/A") V("NOR3X1_892/B") V("NOR3X1_669/C") V("NOR3X1_453/B") V("NOR3X1_454/A") V("NOR3X1_454/C") V("NOR3X1_650/C") V("NOR3X1_649/A") V("NOR3X1_1551/A") V("NOR3X1_1552/C") V("NOR3X1_335/A") V("NOR3X1_336/C") V("NOR3X1_615/A") V("NOR3X1_616/C") V("NOR3X1_293/A") V("NOR3X1_294/B") V("NOR3X1_1415/A") V("NOR3X1_1416/C") V("NOR3X1_811/B") V("NOR3X1_1039/B") V("NOR3X1_1040/A") V("NOR3X1_1040/C") V("NOR3X1_1351/B") V("NOR3X1_391/B") V("NOR3X1_392/A") V("NOR3X1_392/C") V("NOR3X1_1667/C") V("NOR3X1_1668/A") V("NOR3X1_1668/B") V("NOR3X1_1557/C") V("NOR3X1_1558/A") V("NOR3X1_1558/B") V("NOR3X1_1411/C") V("NOR3X1_1538/A") V("NOR3X1_1538/B") V("NOR3X1_1675/A") V("NOR3X1_1676/C") V("NOR3X1_1069/A") V("NOR3X1_1070/B") V("NOR3X1_1011/A") V("NOR3X1_1012/B") V("NOR3X1_894/C") V("NOR3X1_893/A") V("NOR3X1_389/A") V("NOR3X1_390/B") V("NOR3X1_275/A") V("NOR3X1_276/B") V("NOR3X1_1696/B") V("NOR3X1_1695/A") V("NOR3X1_1695/B") V("NOR3X1_1696/A") V("NOR3X1_1696/C") V("NOR3X1_1040/B") V("NOR3X1_1039/A") V("NOR3X1_391/A") V("NOR3X1_392/B") V("NOR3X1_1668/C") V("NOR3X1_1558/C") V("NOR3X1_1557/A") V("NOR3X1_1667/A") V("NOR3X1_1577/A") V("NOR3X1_1578/C") V("NOR3X1_1559/C") V("NOR3X1_1560/A") V("NOR3X1_1560/B") V("NOR3X1_1661/C") V("NOR3X1_1662/B") V("NOR3X1_1664/A") V("NOR3X1_1664/C") V("NOR3X1_1663/B") V("NOR3X1_1260/C") V("NOR3X1_1259/A") V("NOR3X1_1685/A") V("NOR3X1_573/A") V("NOR3X1_1686/B") V("NOR3X1_574/C") V("NOR3X1_1085/A") V("NOR3X1_1086/B") V("NOR3X1_604/B") V("NOR3X1_603/A") V("NOR3X1_601/A") V("NOR3X1_602/B") V("NOR3X1_1661/A") V("NOR3X1_1560/C") V("NOR3X1_1559/A") V("NOR3X1_1664/B") V("NOR3X1_1663/A") V("NOR3X1_453/A") V("NOR3X1_454/B") V("NOR3X1_891/A") V("NOR3X1_1408/B") V("NOR3X1_892/C") V("NOR3X1_1407/A") V("NOR3X1_665/A") V("NOR3X1_666/B") V("NOR3X1_572/C") V("NOR3X1_571/A") V("NOR3X1_1261/A") V("NOR3X1_1262/B") V("NOR3X1_1617/C") V("NOR3X1_1618/C") V("NOR3X1_1617/A") V("NOR3X1_668/B") V("NOR3X1_667/A") V("NOR3X1_1671/A") V("NOR3X1_1672/B") V("NOR3X1_479/A") V("NOR3X1_480/B") V("NOR3X1_1458/B") V("NOR3X1_1457/A") V("NOR3X1_1710/C") V("NOR3X1_1709/A") V("NOR3X1_1709/C") V("NOR3X1_1457/B") V("NOR3X1_649/B") V("NOR3X1_1094/C") V("NOR3X1_1093/A") V("NOR3X1_1093/C") V("NOR3X1_1094/A") V("NOR3X1_1094/B") V("NOR3X1_664/A") V("NOR3X1_664/B") V("NOR3X1_663/C") V("NOR3X1_664/C") V("NOR3X1_663/A") V("NOR3X1_1031/A") V("NOR3X1_1032/C") V("NOR3X1_1458/C") V("NOR3X1_1710/A") V("NOR3X1_1710/B") V("NOR3X1_1458/A") V("NOR3X1_1031/B") V("NOR3X1_721/A") V("NOR3X1_721/B") V("NOR3X1_722/B") V("NOR3X1_945/A") V("NOR3X1_945/B") V("NOR3X1_946/B") V("NOR3X1_722/A") V("NOR3X1_722/C") V("NOR3X1_946/A") V("NOR3X1_946/C") V("NOR3X1_1618/A") V("NOR3X1_1618/B") V("INVX1_1198/Y") V("INVX1_1197/Y") V("INVX1_176/Y") V("INVX1_175/Y") V("INVX1_131/Y") V("INVX1_132/Y") V("INVX1_747/Y") V("INVX1_748/Y") V("INVX1_239/Y") V("INVX1_240/Y") V("INVX1_653/Y") V("INVX1_654/Y") V("INVX1_1198/A") V("INVX1_548/A") V("INVX1_547/A") V("INVX1_1197/A") V("INVX1_176/A") V("INVX1_175/A") V("INVX1_822/A") V("INVX1_821/A") V("INVX1_1377/A") V("INVX1_1378/A") V("INVX1_131/A") V("INVX1_132/A") V("INVX1_747/A") V("INVX1_748/A") V("INVX1_1640/A") V("INVX1_1639/A") V("INVX1_239/A") V("INVX1_240/A") V("INVX1_653/A") V("INVX1_654/A") V("INVX1_750/A") V("INVX1_749/A") V("INVX1_1060/A") V("INVX1_1059/A") V("INVX1_369/A") V("INVX1_370/A") V("NOR3X1_175/B") V("NOR3X1_821/B") V("NOR3X1_747/B") V("NOR3X1_653/B") V("INVX1_174/Y") V("INVX1_173/Y") V("INVX1_820/Y") V("INVX1_819/Y") V("INVX1_1520/Y") V("INVX1_1519/Y") V("INVX1_537/Y") V("INVX1_538/Y") V("INVX1_745/Y") V("INVX1_746/Y") V("INVX1_528/Y") V("INVX1_527/Y") V("INVX1_174/A") V("INVX1_173/A") V("INVX1_820/A") V("INVX1_819/A") V("INVX1_1520/A") V("INVX1_1519/A") V("INVX1_537/A") V("INVX1_539/A") V("INVX1_540/A") V("INVX1_538/A") V("INVX1_745/A") V("INVX1_746/A") V("INVX1_528/A") V("INVX1_527/A") V("NOR3X1_1519/B") V("INVX1_1370/Y") V("INVX1_1372/Y") V("INVX1_1371/Y") V("INVX1_1369/Y") V("INVX1_1370/A") V("INVX1_1372/A") V("INVX1_1371/A") V("INVX1_1369/A") V("NOR3X1_1371/C") V("NOR3X1_1369/B") V("INVX1_1364/Y") V("INVX1_1363/Y") V("INVX1_1366/Y") V("INVX1_1365/Y") V("INVX1_1364/A") V("INVX1_1363/A") V("INVX1_1366/A") V("INVX1_1365/A") V("INVX1_855/Y") V("INVX1_856/Y") V("INVX1_1508/Y") V("INVX1_1507/Y") V("INVX1_376/Y") V("INVX1_375/Y") V("INVX1_372/Y") V("INVX1_1063/Y") V("INVX1_371/Y") V("INVX1_1064/Y") V("INVX1_1327/Y") V("INVX1_1216/Y") V("INVX1_1215/Y") V("INVX1_1328/Y") V("INVX1_766/Y") V("INVX1_765/Y") V("INVX1_259/Y") V("INVX1_260/Y") V("INVX1_1354/Y") V("INVX1_1353/Y") V("INVX1_156/Y") V("INVX1_155/Y") V("INVX1_311/Y") V("INVX1_312/Y") V("INVX1_498/Y") V("INVX1_497/Y") V("INVX1_1227/Y") V("INVX1_1228/Y") V("INVX1_1179/Y") V("INVX1_1180/Y") V("INVX1_1656/Y") V("INVX1_1655/Y") V("INVX1_1511/Y") V("INVX1_1512/Y") V("INVX1_209/Y") V("INVX1_210/Y") V("INVX1_493/Y") V("INVX1_494/Y") V("INVX1_302/Y") V("INVX1_301/Y") V("INVX1_323/Y") V("INVX1_324/Y") V("INVX1_1062/Y") V("INVX1_1061/Y") V("INVX1_1396/Y") V("INVX1_1395/Y") V("INVX1_524/Y") V("INVX1_523/Y") V("INVX1_580/Y") V("INVX1_579/Y") V("INVX1_610/Y") V("INVX1_609/Y") V("INVX1_236/Y") V("INVX1_235/Y") V("INVX1_393/Y") V("INVX1_394/Y") V("INVX1_992/Y") V("INVX1_991/Y") V("INVX1_1340/Y") V("INVX1_1339/Y") V("INVX1_1673/Y") V("INVX1_1674/Y") V("INVX1_82/Y") V("INVX1_81/Y") V("INVX1_478/Y") V("INVX1_477/Y") V("INVX1_840/Y") V("INVX1_839/Y") V("INVX1_1065/Y") V("INVX1_1066/Y") V("INVX1_270/Y") V("INVX1_269/Y") V("INVX1_1172/Y") V("INVX1_1171/Y") V("INVX1_965/Y") V("INVX1_966/Y") V("INVX1_192/Y") V("INVX1_191/Y") V("INVX1_1257/Y") V("INVX1_1258/Y") V("INVX1_150/Y") V("INVX1_149/Y") V("INVX1_596/Y") V("INVX1_595/Y") V("INVX1_630/Y") V("INVX1_629/Y") V("INVX1_1335/Y") V("INVX1_1336/Y") V("INVX1_496/Y") V("INVX1_495/Y") V("INVX1_502/Y") V("INVX1_501/Y") V("INVX1_567/Y") V("INVX1_568/Y") V("INVX1_832/Y") V("INVX1_831/Y") V("INVX1_508/Y") V("INVX1_507/Y") V("INVX1_758/Y") V("INVX1_757/Y") V("INVX1_1502/Y") V("INVX1_1501/Y") V("INVX1_520/Y") V("INVX1_519/Y") V("INVX1_977/Y") V("INVX1_978/Y") V("INVX1_197/Y") V("INVX1_198/Y") V("INVX1_1219/Y") V("INVX1_1220/Y") V("INVX1_768/Y") V("INVX1_767/Y") V("INVX1_1516/Y") V("INVX1_1515/Y") V("INVX1_1646/Y") V("INVX1_1645/Y") V("INVX1_463/Y") V("INVX1_464/Y") V("INVX1_1274/Y") V("INVX1_1273/Y") V("INVX1_759/Y") V("INVX1_760/Y") V("INVX1_1528/Y") V("INVX1_1527/Y") V("INVX1_103/Y") V("INVX1_104/Y") V("INVX1_854/Y") V("INVX1_853/Y") V("INVX1_1390/Y") V("INVX1_1389/Y") V("INVX1_770/Y") V("INVX1_769/Y") V("INVX1_662/Y") V("INVX1_661/Y") V("INVX1_1241/Y") V("INVX1_1242/Y") V("INVX1_913/Y") V("INVX1_914/Y") V("INVX1_476/Y") V("INVX1_475/Y") V("INVX1_330/Y") V("INVX1_329/Y") V("INVX1_613/Y") V("INVX1_614/Y") V("INVX1_1394/Y") V("INVX1_1393/Y") V("INVX1_283/Y") V("INVX1_284/Y") V("INVX1_342/Y") V("INVX1_341/Y") V("INVX1_569/Y") V("INVX1_570/Y") V("INVX1_626/Y") V("INVX1_625/Y") V("INVX1_836/Y") V("INVX1_835/Y") V("INVX1_974/Y") V("INVX1_973/Y") V("INVX1_448/Y") V("INVX1_447/Y") V("INVX1_1036/Y") V("INVX1_1035/Y") V("INVX1_90/Y") V("INVX1_89/Y") V("INVX1_1691/Y") V("INVX1_1692/Y") V("INVX1_308/Y") V("INVX1_307/Y") V("INVX1_1488/Y") V("INVX1_1487/Y") V("INVX1_864/Y") V("INVX1_846/Y") V("INVX1_845/Y") V("INVX1_863/Y") V("INVX1_1603/Y") V("INVX1_1604/Y") V("INVX1_1658/Y") V("INVX1_1657/Y") V("INVX1_1056/Y") V("INVX1_1055/Y") V("INVX1_218/Y") V("INVX1_217/Y") V("INVX1_534/Y") V("INVX1_533/Y") V("INVX1_232/Y") V("INVX1_231/Y") V("INVX1_855/A") V("INVX1_856/A") V("INVX1_1508/A") V("INVX1_1507/A") V("INVX1_376/A") V("INVX1_375/A") V("INVX1_372/A") V("INVX1_1063/A") V("INVX1_371/A") V("INVX1_1064/A") V("INVX1_1327/A") V("INVX1_1216/A") V("INVX1_1215/A") V("INVX1_1328/A") V("INVX1_766/A") V("INVX1_765/A") V("INVX1_259/A") V("INVX1_260/A") V("INVX1_1354/A") V("INVX1_1353/A") V("INVX1_156/A") V("INVX1_155/A") V("INVX1_311/A") V("INVX1_312/A") V("INVX1_498/A") V("INVX1_497/A") V("INVX1_1227/A") V("INVX1_1228/A") V("INVX1_1179/A") V("INVX1_1180/A") V("INVX1_1656/A") V("INVX1_1655/A") V("INVX1_1511/A") V("INVX1_1512/A") V("INVX1_209/A") V("INVX1_210/A") V("INVX1_493/A") V("INVX1_494/A") V("INVX1_302/A") V("INVX1_301/A") V("INVX1_323/A") V("INVX1_324/A") V("INVX1_1062/A") V("INVX1_1061/A") V("INVX1_1396/A") V("INVX1_1395/A") V("INVX1_524/A") V("INVX1_523/A") V("INVX1_580/A") V("INVX1_579/A") V("INVX1_610/A") V("INVX1_609/A") V("INVX1_236/A") V("INVX1_235/A") V("INVX1_393/A") V("INVX1_394/A") V("INVX1_992/A") V("INVX1_991/A") V("INVX1_1340/A") V("INVX1_1339/A") V("INVX1_1673/A") V("INVX1_1674/A") V("INVX1_82/A") V("INVX1_81/A") V("INVX1_478/A") V("INVX1_477/A") V("INVX1_840/A") V("INVX1_839/A") V("INVX1_1065/A") V("INVX1_1066/A") V("INVX1_270/A") V("INVX1_269/A") V("INVX1_1172/A") V("INVX1_1171/A") V("INVX1_965/A") V("INVX1_966/A") V("INVX1_192/A") V("INVX1_191/A") V("INVX1_1257/A") V("INVX1_1258/A") V("INVX1_150/A") V("INVX1_149/A") V("INVX1_596/A") V("INVX1_595/A") V("INVX1_630/A") V("INVX1_629/A") V("INVX1_1335/A") V("INVX1_1336/A") V("INVX1_496/A") V("INVX1_495/A") V("INVX1_502/A") V("INVX1_501/A") V("INVX1_567/A") V("INVX1_568/A") V("INVX1_832/A") V("INVX1_831/A") V("INVX1_508/A") V("INVX1_507/A") V("INVX1_758/A") V("INVX1_757/A") V("INVX1_1502/A") V("INVX1_1501/A") V("INVX1_520/A") V("INVX1_519/A") V("INVX1_977/A") V("INVX1_978/A") V("INVX1_197/A") V("INVX1_198/A") V("INVX1_1219/A") V("INVX1_1220/A") V("INVX1_768/A") V("INVX1_767/A") V("INVX1_1516/A") V("INVX1_1515/A") V("INVX1_1646/A") V("INVX1_1645/A") V("INVX1_463/A") V("INVX1_464/A") V("INVX1_1274/A") V("INVX1_1273/A") V("INVX1_759/A") V("INVX1_760/A") V("INVX1_1528/A") V("INVX1_1527/A") V("INVX1_103/A") V("INVX1_104/A") V("INVX1_854/A") V("INVX1_853/A") V("INVX1_1390/A") V("INVX1_1389/A") V("INVX1_770/A") V("INVX1_769/A") V("INVX1_662/A") V("INVX1_661/A") V("INVX1_1241/A") V("INVX1_1242/A") V("INVX1_913/A") V("INVX1_914/A") V("INVX1_476/A") V("INVX1_475/A") V("INVX1_330/A") V("INVX1_329/A") V("INVX1_613/A") V("INVX1_614/A") V("INVX1_1394/A") V("INVX1_1393/A") V("INVX1_283/A") V("INVX1_284/A") V("INVX1_342/A") V("INVX1_341/A") V("INVX1_569/A") V("INVX1_570/A") V("INVX1_626/A") V("INVX1_625/A") V("INVX1_836/A") V("INVX1_835/A") V("INVX1_974/A") V("INVX1_973/A") V("INVX1_448/A") V("INVX1_447/A") V("INVX1_1036/A") V("INVX1_1035/A") V("INVX1_90/A") V("INVX1_89/A") V("INVX1_1691/A") V("INVX1_1692/A") V("INVX1_308/A") V("INVX1_307/A") V("INVX1_1488/A") V("INVX1_1487/A") V("INVX1_864/A") V("INVX1_846/A") V("INVX1_845/A") V("INVX1_863/A") V("INVX1_1603/A") V("INVX1_1604/A") V("INVX1_1658/A") V("INVX1_1657/A") V("INVX1_1056/A") V("INVX1_1055/A") V("INVX1_218/A") V("INVX1_217/A") V("INVX1_534/A") V("INVX1_533/A") V("NOR3X1_1507/B") V("NOR3X1_375/B") V("NOR3X1_371/B") V("NOR3X1_311/C") V("NOR3X1_393/C") V("NOR3X1_1065/B") V("NOR3X1_495/B") V("NOR3X1_501/B") V("NOR3X1_977/C") V("NOR3X1_197/C") V("NOR3X1_767/B") V("NOR3X1_1273/B") V("NOR3X1_759/B") V("NOR3X1_613/B") V("NOR3X1_1603/A") V("NOR3X1_1603/B") V("NOR3X1_1603/C") V("NOR3X1_1604/A") V("NOR3X1_1604/B") V("NOR3X1_1604/C") V("NOR3X1_1657/B") V("NOR3X1_232/A") V("NOR3X1_232/B") V("NOR3X1_232/C") V("NOR3X1_231/A") V("NOR3X1_231/B") V("NOR3X1_231/C") V("INVX1_320/Y") V("INVX1_322/Y") V("INVX1_321/Y") V("INVX1_319/Y") V("INVX1_1649/Y") V("INVX1_1651/Y") V("INVX1_1652/Y") V("INVX1_1650/Y") V("INVX1_503/Y") V("INVX1_963/Y") V("INVX1_964/Y") V("INVX1_504/Y") V("INVX1_1251/Y") V("INVX1_1253/Y") V("INVX1_1254/Y") V("INVX1_1252/Y") V("INVX1_557/Y") V("INVX1_559/Y") V("INVX1_560/Y") V("INVX1_558/Y") V("INVX1_506/Y") V("INVX1_505/Y") V("INVX1_194/Y") V("INVX1_196/Y") V("INVX1_195/Y") V("INVX1_193/Y") V("INVX1_660/Y") V("INVX1_659/Y") V("INVX1_1231/Y") V("INVX1_1233/Y") V("INVX1_1234/Y") V("INVX1_1232/Y") V("INVX1_735/Y") V("INVX1_740/Y") V("INVX1_739/Y") V("INVX1_736/Y") V("INVX1_561/Y") V("INVX1_563/Y") V("INVX1_564/Y") V("INVX1_562/Y") V("INVX1_1629/Y") V("INVX1_1631/Y") V("INVX1_1632/Y") V("INVX1_1630/Y") V("INVX1_1596/Y") V("INVX1_1598/Y") V("INVX1_1597/Y") V("INVX1_1595/Y") V("INVX1_531/Y") V("INVX1_530/Y") V("INVX1_532/Y") V("INVX1_529/Y") V("INVX1_229/Y") V("INVX1_227/Y") V("INVX1_230/Y") V("INVX1_228/Y") V("INVX1_320/A") V("INVX1_322/A") V("INVX1_321/A") V("INVX1_319/A") V("INVX1_1649/A") V("INVX1_1651/A") V("INVX1_1652/A") V("INVX1_1650/A") V("INVX1_503/A") V("INVX1_963/A") V("INVX1_964/A") V("INVX1_504/A") V("INVX1_1251/A") V("INVX1_1253/A") V("INVX1_1254/A") V("INVX1_1252/A") V("INVX1_557/A") V("INVX1_559/A") V("INVX1_560/A") V("INVX1_558/A") V("INVX1_506/A") V("INVX1_505/A") V("INVX1_194/A") V("INVX1_196/A") V("INVX1_195/A") V("INVX1_193/A") V("INVX1_660/A") V("INVX1_659/A") V("INVX1_1231/A") V("INVX1_1233/A") V("INVX1_1234/A") V("INVX1_1232/A") V("INVX1_735/A") V("INVX1_740/A") V("INVX1_739/A") V("INVX1_736/A") V("INVX1_561/A") V("INVX1_563/A") V("INVX1_564/A") V("INVX1_562/A") V("INVX1_1629/A") V("INVX1_1631/A") V("INVX1_1632/A") V("INVX1_1630/A") V("INVX1_531/A") V("INVX1_530/A") V("INVX1_532/A") V("INVX1_529/A") V("INVX1_229/A") V("INVX1_227/A") V("INVX1_230/A") V("INVX1_228/A") V("NOR3X1_195/B") V("NOR3X1_735/B") V("NOR3X1_1631/B") V("NOR3X1_1596/A") V("NOR3X1_1596/B") V("NOR3X1_1596/C") V("NOR3X1_1598/A") V("NOR3X1_1598/B") V("NOR3X1_1598/C") V("NOR3X1_1597/A") V("NOR3X1_1597/B") V("NOR3X1_1595/A") V("NOR3X1_1595/B") V("NOR3X1_531/C") V("NOR3X1_529/B") V("NOR3X1_227/B") V("INVX1_182/Y") V("INVX1_178/Y") V("INVX1_181/Y") V("INVX1_177/Y") V("INVX1_871/Y") V("INVX1_637/Y") V("INVX1_872/Y") V("INVX1_638/Y") V("INVX1_1185/Y") V("INVX1_1077/Y") V("INVX1_1186/Y") V("INVX1_1078/Y") V("INVX1_211/Y") V("INVX1_224/Y") V("INVX1_223/Y") V("INVX1_212/Y") V("INVX1_215/Y") V("INVX1_226/Y") V("INVX1_225/Y") V("INVX1_216/Y") V("INVX1_182/A") V("INVX1_178/A") V("INVX1_181/A") V("INVX1_177/A") V("INVX1_871/A") V("INVX1_872/A") V("INVX1_1185/A") V("INVX1_1186/A") V("INVX1_211/A") V("INVX1_224/A") V("INVX1_223/A") V("INVX1_212/A") V("INVX1_215/A") V("INVX1_226/A") V("INVX1_225/A") V("INVX1_216/A") V("NOR3X1_871/C") V("NOR3X1_637/A") V("NOR3X1_637/B") V("NOR3X1_637/C") V("NOR3X1_638/A") V("NOR3X1_638/B") V("NOR3X1_638/C") V("NOR3X1_1185/B") V("NOR3X1_1077/A") V("NOR3X1_1077/B") V("NOR3X1_1077/C") V("NOR3X1_1078/A") V("NOR3X1_1078/B") V("NOR3X1_1078/C") V("NOR3X1_211/B") V("NOR3X1_223/C") V("INVX1_868/Y") V("INVX1_870/Y") V("INVX1_869/Y") V("INVX1_867/Y") V("INVX1_634/Y") V("INVX1_636/Y") V("INVX1_635/Y") V("INVX1_633/Y") V("INVX1_1181/Y") V("INVX1_1184/Y") V("INVX1_1183/Y") V("INVX1_1182/Y") V("INVX1_1074/Y") V("INVX1_1076/Y") V("INVX1_1075/Y") V("INVX1_1073/Y") V("INVX1_214/Y") V("INVX1_206/Y") V("INVX1_213/Y") V("INVX1_205/Y") V("INVX1_868/A") V("INVX1_870/A") V("INVX1_869/A") V("INVX1_867/A") V("INVX1_634/A") V("INVX1_636/A") V("INVX1_635/A") V("INVX1_633/A") V("INVX1_1181/A") V("INVX1_1184/A") V("INVX1_1183/A") V("INVX1_1182/A") V("INVX1_1074/A") V("INVX1_1076/A") V("INVX1_1075/A") V("INVX1_1073/A") V("INVX1_214/A") V("INVX1_206/A") V("INVX1_213/A") V("INVX1_205/A") V("NOR3X1_869/C") V("NOR3X1_1181/B") V("INVX1_862/Y") V("INVX1_344/Y") V("INVX1_861/Y") V("INVX1_343/Y") V("INVX1_628/Y") V("INVX1_627/Y") V("INVX1_632/Y") V("INVX1_631/Y") V("INVX1_1178/Y") V("INVX1_1177/Y") V("INVX1_1072/Y") V("INVX1_1071/Y") V("INVX1_622/Y") V("INVX1_26/Y") V("INVX1_621/Y") V("INVX1_25/Y") V("INVX1_862/A") V("INVX1_344/A") V("INVX1_861/A") V("INVX1_343/A") V("INVX1_628/A") V("INVX1_627/A") V("INVX1_632/A") V("INVX1_631/A") V("INVX1_1178/A") V("INVX1_1177/A") V("INVX1_1072/A") V("INVX1_1071/A") V("INVX1_622/A") V("INVX1_26/A") V("INVX1_621/A") V("INVX1_25/A") V("INVX1_370/Y") V("INVX1_369/Y") V("INVX1_540/Y") V("INVX1_539/Y") V("INVX1_1374/Y") V("INVX1_1373/Y") 
    
    if ('showPlots' < 1)
        quit
    end
       
.endc

.end
