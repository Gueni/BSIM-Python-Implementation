*** TEST 004 partitioning ***
*
* ngSPICE test for PLS experiments
*
* AES SBOX PLS test init file generator - protected dualRail SBOX area illuminated
*
* Author: Jan Belohoubek, 08/2020
* jan.belohoubek@fit.cvut.cz
*
* https://users.fit.cvut.cz/~belohja4/
*
*
* **************************************

.include ../../models.lib
.include ../../tsmc180nmcmos.lib
.include pDualRail.spice

* **************************************
* --- Test ---
* **************************************

* --- Settings
.param showPlots = 0
.param writeFile = 1
.param run_inputSet = 0

* redefine defaults ...
.include test00X_settings.inc

.csparam showPlots = {showPlots}
.csparam writeFile = {writeFile}
.csparam run_inputSet = {run_inputSet}

.global showPlots writeFile run_inputSet

* --- End of Settins

Vtrig LaserTrig 0 0 PWL(0ns 0V 20ns 0V 21ns SUPP)

.param beamDistanceTop = 0
.param beamDistanceBot = 0

.global LaserTrig beamDistanceTop beamDistanceBot

* --- inputs
Vvin0 INPUT_0 0 0 PWL(0ns 0V 5ns  0V 7ns  0V)
Vvin1 INPUT_1 0 0 PWL(0ns 0V 6ns  0V 8ns  0V)
Vvin2 INPUT_2 0 0 PWL(0ns 0V 7ns  0V 9ns  0V)
Vvin3 INPUT_3 0 0 PWL(0ns 0V 8ns  0V 10ns 0V)
Vvin4 INPUT_4 0 0 PWL(0ns 0V 9ns  0V 11ns 0V)
Vvin5 INPUT_5 0 0 PWL(0ns 0V 10ns 0V 12ns 0V)
Vvin6 INPUT_6 0 0 PWL(0ns 0V 11ns 0V 13ns 0V)
Vvin7 INPUT_7 0 0 PWL(0ns 0V 12ns 0V 14ns 0V)

Vvin0D D_INPUT_0 0 0 PWL(0ns 0V 5ns  0V 7ns  0V)
Vvin1D D_INPUT_1 0 0 PWL(0ns 0V 6ns  0V 8ns  0V)
Vvin2D D_INPUT_2 0 0 PWL(0ns 0V 7ns  0V 9ns  0V)
Vvin3D D_INPUT_3 0 0 PWL(0ns 0V 8ns  0V 10ns 0V)
Vvin4D D_INPUT_4 0 0 PWL(0ns 0V 9ns  0V 11ns 0V)
Vvin5D D_INPUT_5 0 0 PWL(0ns 0V 10ns 0V 12ns 0V)
Vvin6D D_INPUT_6 0 0 PWL(0ns 0V 11ns 0V 13ns 0V)
Vvin7D D_INPUT_7 0 0 PWL(0ns 0V 12ns 0V 14ns 0V)


* --- circuit layout model

Xsbox1 
+ INPUT_0 INPUT_1 INPUT_2 INPUT_3 INPUT_4 INPUT_5 INPUT_6 INPUT_7 D_INPUT_0 D_INPUT_1 D_INPUT_2 D_INPUT_3 D_INPUT_4 D_INPUT_5 D_INPUT_6 D_INPUT_7 
+ VSS VDD 
+ POR2X1_751/A POR2X1_516/B PAND2X1_809/A PAND2X1_473/B POR2X1_101/A POR2X1_334/A POR2X1_836/A POR2X1_240/A POR2X1_461/Y PAND2X1_691/Y POR2X1_323/Y POR2X1_527/Y POR2X1_111/Y POR2X1_515/Y POR2X1_73/Y POR2X1_41/B POR2X1_669/B PAND2X1_63/B POR2X1_16/A POR2X1_287/B POR2X1_246/Y PAND2X1_464/B POR2X1_815/A POR2X1_309/Y POR2X1_283/Y POR2X1_488/Y POR2X1_289/Y POR2X1_417/Y POR2X1_226/Y PAND2X1_848/B POR2X1_96/B POR2X1_62/Y PAND2X1_90/Y POR2X1_612/A POR2X1_78/A PAND2X1_55/Y POR2X1_590/A POR2X1_378/Y POR2X1_274/B POR2X1_838/B POR2X1_195/A POR2X1_296/Y POR2X1_447/B POR2X1_535/A POR2X1_138/A POR2X1_519/Y POR2X1_692/Y POR2X1_48/Y POR2X1_406/A POR2X1_599/A POR2X1_763/Y 
+ POR2X1_511/Y POR2X1_98/B POR2X1_448/A POR2X1_630/B POR2X1_389/A POR2X1_631/A POR2X1_294/Y POR2X1_415/Y POR2X1_637/B POR2X1_828/A POR2X1_398/Y POR2X1_121/Y POR2X1_302/A POR2X1_450/B POR2X1_606/Y POR2X1_301/A POR2X1_543/A POR2X1_322/Y POR2X1_164/Y POR2X1_144/Y POR2X1_306/Y POR2X1_696/Y POR2X1_503/A POR2X1_588/Y POR2X1_376/Y POR2X1_273/Y POR2X1_433/Y POR2X1_409/B POR2X1_743/Y PAND2X1_156/B POR2X1_673/A POR2X1_549/A POR2X1_391/B POR2X1_619/Y POR2X1_532/A POR2X1_130/A POR2X1_266/A POR2X1_634/A PAND2X1_73/Y PAND2X1_85/Y POR2X1_541/B POR2X1_633/A POR2X1_777/B PAND2X1_39/B POR2X1_186/B POR2X1_83/A POR2X1_77/Y POR2X1_693/Y POR2X1_23/Y POR2X1_49/Y POR2X1_748/A 
+ PAND2X1_377/Y POR2X1_387/Y POR2X1_329/Y POR2X1_421/Y POR2X1_597/A POR2X1_72/B POR2X1_40/Y POR2X1_416/B POR2X1_7/B POR2X1_790/B POR2X1_694/Y POR2X1_426/Y PAND2X1_52/B PAND2X1_32/B PAND2X1_57/B PAND2X1_48/B POR2X1_304/Y POR2X1_56/Y POR2X1_409/Y POR2X1_635/A POR2X1_769/B POR2X1_430/Y PAND2X1_69/A PAND2X1_20/A POR2X1_260/A POR2X1_52/A POR2X1_96/A POR2X1_65/A POR2X1_513/Y POR2X1_855/B POR2X1_325/A POR2X1_547/B POR2X1_332/B POR2X1_557/A POR2X1_411/B POR2X1_394/A POR2X1_344/A PAND2X1_19/Y POR2X1_7/A POR2X1_748/Y POR2X1_516/A POR2X1_750/Y POR2X1_129/Y POR2X1_29/Y POR2X1_383/A POR2X1_68/A POR2X1_614/A POR2X1_81/A POR2X1_291/Y POR2X1_824/Y POR2X1_234/Y 
+ PAND2X1_462/B POR2X1_809/B POR2X1_276/Y PAND2X1_101/B POR2X1_708/B POR2X1_638/B POR2X1_459/B POR2X1_325/B POR2X1_776/B POR2X1_147/A POR2X1_502/Y POR2X1_308/B POR2X1_155/Y POR2X1_274/A POR2X1_832/A POR2X1_780/B POR2X1_407/Y POR2X1_458/Y PAND2X1_48/Y POR2X1_405/Y POR2X1_513/B POR2X1_520/A POR2X1_706/B POR2X1_335/B POR2X1_286/B POR2X1_489/A POR2X1_814/Y POR2X1_333/A POR2X1_446/B POR2X1_227/A POR2X1_481/A POR2X1_416/A POR2X1_625/Y POR2X1_399/A POR2X1_585/Y POR2X1_257/A PAND2X1_81/B PAND2X1_82/Y POR2X1_38/Y POR2X1_87/B POR2X1_236/Y POR2X1_382/Y POR2X1_300/Y POR2X1_369/Y POR2X1_607/A POR2X1_299/Y POR2X1_122/A POR2X1_848/A POR2X1_750/B POR2X1_294/B POR2X1_342/B 
+ POR2X1_78/B POR2X1_278/Y POR2X1_102/Y PAND2X1_612/B POR2X1_55/Y PAND2X1_94/Y POR2X1_90/Y POR2X1_136/Y POR2X1_43/Y POR2X1_297/A POR2X1_272/Y POR2X1_827/Y POR2X1_419/Y POR2X1_459/A POR2X1_534/Y POR2X1_814/B PAND2X1_6/Y POR2X1_490/Y POR2X1_20/A PAND2X1_23/Y POR2X1_256/Y POR2X1_789/B POR2X1_93/Y POR2X1_422/Y POR2X1_628/Y POR2X1_63/Y POR2X1_672/Y PAND2X1_71/Y POR2X1_68/Y POR2X1_198/B POR2X1_778/B POR2X1_335/A POR2X1_71/Y POR2X1_57/Y POR2X1_69/A POR2X1_372/A POR2X1_310/Y POR2X1_378/A POR2X1_706/A POR2X1_709/A POR2X1_622/B POR2X1_85/Y POR2X1_263/Y POR2X1_413/A POR2X1_278/A POR2X1_255/Y POR2X1_245/Y POR2X1_150/Y PAND2X1_63/Y PAND2X1_549/B POR2X1_355/B 
+ POR2X1_448/B POR2X1_596/Y PAND2X1_96/B POR2X1_260/B PAND2X1_60/B POR2X1_43/B POR2X1_39/B POR2X1_83/B POR2X1_66/B PAND2X1_72/A PAND2X1_41/B POR2X1_753/Y PAND2X1_65/B PAND2X1_58/A POR2X1_66/A PAND2X1_56/Y POR2X1_307/B POR2X1_707/B POR2X1_13/A POR2X1_60/A POR2X1_20/B POR2X1_32/A POR2X1_57/A POR2X1_48/A POR2X1_582/Y POR2X1_460/A POR2X1_451/A POR2X1_760/A POR2X1_66/Y POR2X1_121/A POR2X1_188/A POR2X1_327/Y POR2X1_67/A POR2X1_666/A POR2X1_816/A PAND2X1_687/Y POR2X1_271/A POR2X1_87/Y POR2X1_410/Y POR2X1_373/Y POR2X1_667/A POR2X1_411/A POR2X1_687/Y POR2X1_270/Y POR2X1_88/A POR2X1_544/B POR2X1_264/Y POR2X1_683/Y POR2X1_682/Y POR2X1_685/A POR2X1_686/B 
+ POR2X1_88/Y PAND2X1_717/A POR2X1_761/A POR2X1_644/A POR2X1_717/B PAND2X1_88/Y
+ AES_SBOX_0


* **************************************
* --- Simulation Settings ---
* **************************************

.param SIM_LEN = 35ns
.csparam SIM_LEN = {SIM_LEN}

.tran 0.1ns 'SIM_LEN'
.param SIMSTEP = 'SIM_LEN/0.1ns'
.csparam SIMSTEP = {SIMSTEP}

* **************************************
* --- Simulation Control ---
* **************************************

.control
    .include ../inputsD.inc

    run
    
    if ('writeFile' > 0)   
      wrdata ivdd_0.out i(vvdd)
      wrdata ivss_0.out i(vvss)
      *snsave sim_0.snap
    end
    
    set wr_vecnames
    set wr_singlescale
    wrdata outputs_0.out V("POR2X1_751/A") V("POR2X1_516/B") V("PAND2X1_809/A") V("PAND2X1_473/B") V("POR2X1_101/A") V("POR2X1_334/A") V("POR2X1_836/A") V("POR2X1_240/A") V("POR2X1_461/Y") V("PAND2X1_691/Y") V("POR2X1_323/Y") V("POR2X1_527/Y") V("POR2X1_111/Y") V("POR2X1_515/Y") V("POR2X1_73/Y") V("POR2X1_41/B") V("POR2X1_669/B") V("PAND2X1_63/B") V("POR2X1_16/A") V("POR2X1_287/B") V("POR2X1_246/Y") V("PAND2X1_464/B") V("POR2X1_815/A") V("POR2X1_309/Y") V("POR2X1_283/Y") V("POR2X1_488/Y") V("POR2X1_289/Y") V("POR2X1_417/Y") V("POR2X1_226/Y") V("PAND2X1_848/B") V("POR2X1_96/B") V("POR2X1_62/Y") V("PAND2X1_90/Y") V("POR2X1_612/A") V("POR2X1_78/A") V("PAND2X1_55/Y") V("POR2X1_590/A") V("POR2X1_378/Y") V("POR2X1_274/B") V("POR2X1_838/B") V("POR2X1_195/A") V("POR2X1_296/Y") V("POR2X1_447/B") V("POR2X1_535/A") V("POR2X1_138/A") V("POR2X1_519/Y") V("POR2X1_692/Y") V("POR2X1_48/Y") V("POR2X1_406/A") V("POR2X1_599/A") V("POR2X1_763/Y") V("POR2X1_511/Y") V("POR2X1_98/B") V("POR2X1_448/A") V("POR2X1_630/B") V("POR2X1_389/A") V("POR2X1_631/A") V("POR2X1_294/Y") V("POR2X1_415/Y") V("POR2X1_637/B") V("POR2X1_828/A") V("POR2X1_398/Y") V("POR2X1_121/Y") V("POR2X1_302/A") V("POR2X1_450/B") V("POR2X1_606/Y") V("POR2X1_301/A") V("POR2X1_543/A") V("POR2X1_322/Y") V("POR2X1_164/Y") V("POR2X1_144/Y") V("POR2X1_306/Y") V("POR2X1_696/Y") V("POR2X1_503/A") V("POR2X1_588/Y") V("POR2X1_376/Y") V("POR2X1_273/Y") V("POR2X1_433/Y") V("POR2X1_409/B") V("POR2X1_743/Y") V("PAND2X1_156/B") V("POR2X1_673/A") V("POR2X1_549/A") V("POR2X1_391/B") V("POR2X1_619/Y") V("POR2X1_532/A") V("POR2X1_130/A") V("POR2X1_266/A") V("POR2X1_634/A") V("PAND2X1_73/Y") V("PAND2X1_85/Y") V("POR2X1_541/B") V("POR2X1_633/A") V("POR2X1_777/B") V("PAND2X1_39/B") V("POR2X1_186/B") V("POR2X1_83/A") V("POR2X1_77/Y") V("POR2X1_693/Y") V("POR2X1_23/Y") V("POR2X1_49/Y") V("POR2X1_748/A") V("PAND2X1_377/Y") V("POR2X1_387/Y") V("POR2X1_329/Y") V("POR2X1_421/Y") V("POR2X1_597/A") V("POR2X1_72/B") V("POR2X1_40/Y") V("POR2X1_416/B") V("POR2X1_7/B") V("POR2X1_790/B") V("POR2X1_694/Y") V("POR2X1_426/Y") V("PAND2X1_52/B") V("PAND2X1_32/B") V("PAND2X1_57/B") V("PAND2X1_48/B") V("POR2X1_304/Y") V("POR2X1_56/Y") V("POR2X1_409/Y") V("POR2X1_635/A") V("POR2X1_769/B") V("POR2X1_430/Y") V("PAND2X1_69/A") V("PAND2X1_20/A") V("POR2X1_260/A") V("POR2X1_52/A") V("POR2X1_96/A") V("POR2X1_65/A") V("POR2X1_513/Y") V("POR2X1_855/B") V("POR2X1_325/A") V("POR2X1_547/B") V("POR2X1_332/B") V("POR2X1_557/A") V("POR2X1_411/B") V("POR2X1_394/A") V("POR2X1_344/A") V("PAND2X1_19/Y") V("POR2X1_7/A") V("POR2X1_748/Y") V("POR2X1_516/A") V("POR2X1_750/Y") V("POR2X1_129/Y") V("POR2X1_29/Y") V("POR2X1_383/A") V("POR2X1_68/A") V("POR2X1_614/A") V("POR2X1_81/A") V("POR2X1_291/Y") V("POR2X1_824/Y") V("POR2X1_234/Y") V("PAND2X1_462/B") V("POR2X1_809/B") V("POR2X1_276/Y") V("PAND2X1_101/B") V("POR2X1_708/B") V("POR2X1_638/B") V("POR2X1_459/B") V("POR2X1_325/B") V("POR2X1_776/B") V("POR2X1_147/A") V("POR2X1_502/Y") V("POR2X1_308/B") V("POR2X1_155/Y") V("POR2X1_274/A") V("POR2X1_832/A") V("POR2X1_780/B") V("POR2X1_407/Y") V("POR2X1_458/Y") V("PAND2X1_48/Y") V("POR2X1_405/Y") V("POR2X1_513/B") V("POR2X1_520/A") V("POR2X1_706/B") V("POR2X1_335/B") V("POR2X1_286/B") V("POR2X1_489/A") V("POR2X1_814/Y") V("POR2X1_333/A") V("POR2X1_446/B") V("POR2X1_227/A") V("POR2X1_481/A") V("POR2X1_416/A") V("POR2X1_625/Y") V("POR2X1_399/A") V("POR2X1_585/Y") V("POR2X1_257/A") V("PAND2X1_81/B") V("PAND2X1_82/Y") V("POR2X1_38/Y") V("POR2X1_87/B") V("POR2X1_236/Y") V("POR2X1_382/Y") V("POR2X1_300/Y") V("POR2X1_369/Y") V("POR2X1_607/A") V("POR2X1_299/Y") V("POR2X1_122/A") V("POR2X1_848/A") V("POR2X1_750/B") V("POR2X1_294/B") V("POR2X1_342/B") V("POR2X1_78/B") V("POR2X1_278/Y") V("POR2X1_102/Y") V("PAND2X1_612/B") V("POR2X1_55/Y") V("PAND2X1_94/Y") V("POR2X1_90/Y") V("POR2X1_136/Y") V("POR2X1_43/Y") V("POR2X1_297/A") V("POR2X1_272/Y") V("POR2X1_827/Y") V("POR2X1_419/Y") V("POR2X1_459/A") V("POR2X1_534/Y") V("POR2X1_814/B") V("PAND2X1_6/Y") V("POR2X1_490/Y") V("POR2X1_20/A") V("PAND2X1_23/Y") V("POR2X1_256/Y") V("POR2X1_789/B") V("POR2X1_93/Y") V("POR2X1_422/Y") V("POR2X1_628/Y") V("POR2X1_63/Y") V("POR2X1_672/Y") V("PAND2X1_71/Y") V("POR2X1_68/Y") V("POR2X1_198/B") V("POR2X1_778/B") V("POR2X1_335/A") V("POR2X1_71/Y") V("POR2X1_57/Y") V("POR2X1_69/A") V("POR2X1_372/A") V("POR2X1_310/Y") V("POR2X1_378/A") V("POR2X1_706/A") V("POR2X1_709/A") V("POR2X1_622/B") V("POR2X1_85/Y") V("POR2X1_263/Y") V("POR2X1_413/A") V("POR2X1_278/A") V("POR2X1_255/Y") V("POR2X1_245/Y") V("POR2X1_150/Y") V("PAND2X1_63/Y") V("PAND2X1_549/B") V("POR2X1_355/B") V("POR2X1_448/B") V("POR2X1_596/Y") V("PAND2X1_96/B") V("POR2X1_260/B") V("PAND2X1_60/B") V("POR2X1_43/B") V("POR2X1_39/B") V("POR2X1_83/B") V("POR2X1_66/B") V("PAND2X1_72/A") V("PAND2X1_41/B") V("POR2X1_753/Y") V("PAND2X1_65/B") V("PAND2X1_58/A") V("POR2X1_66/A") V("PAND2X1_56/Y") V("POR2X1_307/B") V("POR2X1_707/B") V("POR2X1_13/A") V("POR2X1_60/A") V("POR2X1_20/B") V("POR2X1_32/A") V("POR2X1_57/A") V("POR2X1_48/A") V("POR2X1_582/Y") V("POR2X1_460/A") V("POR2X1_451/A") V("POR2X1_760/A") V("POR2X1_66/Y") V("POR2X1_121/A") V("POR2X1_188/A") V("POR2X1_327/Y") V("POR2X1_67/A") V("POR2X1_666/A") V("POR2X1_816/A") V("PAND2X1_687/Y") V("POR2X1_271/A") V("POR2X1_87/Y") V("POR2X1_410/Y") V("POR2X1_373/Y") V("POR2X1_667/A") V("POR2X1_411/A") V("POR2X1_687/Y") V("POR2X1_270/Y") V("POR2X1_88/A") V("POR2X1_544/B") V("POR2X1_264/Y") V("POR2X1_683/Y") V("POR2X1_682/Y") V("POR2X1_685/A") V("POR2X1_686/B") V("POR2X1_88/Y") V("PAND2X1_717/A") V("POR2X1_761/A") V("POR2X1_644/A") V("POR2X1_717/B") V("PAND2X1_88/Y") 
    
    if ('showPlots' < 1)
        quit
    end
       
.endc

.end
