magic
tech scmos
magscale 1 2
timestamp 1598351945
<< error_s >>
rect 2524 2996 2532 3004
rect 220 2976 228 2984
rect 524 2976 532 2984
rect 860 2976 868 2984
rect 1692 2976 1700 2984
rect 2972 2976 2980 2984
rect 3996 2976 4004 2984
rect 12 2956 20 2964
rect 156 2956 164 2964
rect 700 2956 708 2964
rect 972 2956 980 2964
rect 1100 2956 1108 2964
rect 1164 2956 1172 2964
rect 1436 2956 1444 2964
rect 1516 2956 1524 2964
rect 1532 2956 1540 2964
rect 1596 2956 1604 2964
rect 1740 2956 1748 2964
rect 1772 2956 1780 2964
rect 2012 2956 2020 2964
rect 2124 2956 2132 2964
rect 2156 2956 2164 2964
rect 2220 2956 2228 2964
rect 2364 2956 2372 2964
rect 2572 2956 2580 2964
rect 2668 2956 2676 2964
rect 2764 2956 2772 2964
rect 3564 2956 3572 2964
rect 3708 2956 3716 2964
rect 764 2936 772 2944
rect 844 2936 852 2944
rect 1148 2936 1156 2944
rect 1692 2936 1700 2944
rect 2956 2936 2964 2944
rect 3084 2936 3092 2944
rect 3228 2936 3236 2944
rect 3244 2936 3252 2944
rect 3292 2936 3300 2944
rect 3372 2936 3380 2944
rect 3628 2936 3636 2944
rect 460 2916 468 2924
rect 764 2916 772 2924
rect 2396 2916 2404 2924
rect 2412 2916 2420 2924
rect 3148 2916 3156 2924
rect 3276 2916 3284 2924
rect 3532 2916 3540 2924
rect 92 2896 100 2904
rect 124 2896 132 2904
rect 252 2896 260 2904
rect 332 2896 340 2904
rect 476 2896 484 2904
rect 572 2896 580 2904
rect 652 2896 660 2904
rect 908 2896 916 2904
rect 972 2896 980 2904
rect 1116 2896 1124 2904
rect 2476 2896 2484 2904
rect 2604 2896 2612 2904
rect 3644 2896 3652 2904
rect 3836 2896 3844 2904
rect 3884 2896 3892 2904
rect 4156 2896 4164 2904
rect 684 2876 692 2884
rect 1564 2876 1572 2884
rect 3724 2876 3732 2884
rect 3756 2876 3764 2884
rect 1276 2856 1284 2864
rect 2444 2856 2452 2864
rect 1388 2836 1396 2844
rect 3420 2816 3428 2824
rect 4204 2796 4212 2804
rect 652 2776 660 2784
rect 2092 2776 2100 2784
rect 4060 2776 4068 2784
rect 4092 2776 4100 2784
rect 1452 2756 1460 2764
rect 2412 2756 2420 2764
rect 3836 2756 3844 2764
rect 4156 2756 4164 2764
rect 1020 2736 1028 2744
rect 1708 2736 1716 2744
rect 2444 2736 2452 2744
rect 124 2716 132 2724
rect 412 2716 420 2724
rect 716 2716 724 2724
rect 956 2716 964 2724
rect 1356 2716 1364 2724
rect 1484 2716 1492 2724
rect 1532 2716 1540 2724
rect 2636 2716 2644 2724
rect 2780 2716 2788 2724
rect 2876 2716 2884 2724
rect 3004 2716 3012 2724
rect 3228 2716 3236 2724
rect 3468 2716 3476 2724
rect 3596 2716 3604 2724
rect 3660 2716 3668 2724
rect 3724 2716 3732 2724
rect 3756 2716 3764 2724
rect 3852 2716 3860 2724
rect 3900 2716 3908 2724
rect 1004 2696 1012 2704
rect 380 2676 388 2684
rect 828 2676 836 2684
rect 1244 2676 1252 2684
rect 1436 2676 1444 2684
rect 2092 2676 2100 2684
rect 2108 2676 2116 2684
rect 2204 2676 2212 2684
rect 3548 2676 3556 2684
rect 3644 2676 3652 2684
rect 3932 2676 3940 2684
rect 524 2656 532 2664
rect 636 2656 644 2664
rect 876 2656 884 2664
rect 972 2656 980 2664
rect 1164 2656 1172 2664
rect 1292 2656 1300 2664
rect 1548 2656 1556 2664
rect 1820 2656 1828 2664
rect 2348 2656 2356 2664
rect 2540 2656 2548 2664
rect 2572 2656 2580 2664
rect 2732 2656 2740 2664
rect 3404 2656 3412 2664
rect 3724 2656 3732 2664
rect 3820 2656 3828 2664
rect 4108 2656 4116 2664
rect 4140 2656 4148 2664
rect 44 2636 52 2644
rect 524 2636 532 2644
rect 1196 2636 1204 2644
rect 1660 2636 1668 2644
rect 1756 2636 1764 2644
rect 1772 2636 1780 2644
rect 1932 2636 1940 2644
rect 2044 2636 2052 2644
rect 284 2616 292 2624
rect 812 2616 820 2624
rect 908 2616 916 2624
rect 2236 2616 2244 2624
rect 2444 2616 2452 2624
rect 2556 2616 2564 2624
rect 2972 2616 2980 2624
rect 652 2596 660 2604
rect 1564 2596 1572 2604
rect 1868 2596 1876 2604
rect 3100 2596 3108 2604
rect 3164 2596 3172 2604
rect 3180 2596 3188 2604
rect 3500 2596 3508 2604
rect 3516 2596 3524 2604
rect 3916 2596 3924 2604
rect 76 2576 84 2584
rect 396 2576 404 2584
rect 1388 2576 1396 2584
rect 3708 2576 3716 2584
rect 3804 2576 3812 2584
rect 4092 2576 4100 2584
rect 172 2556 180 2564
rect 444 2556 452 2564
rect 508 2556 516 2564
rect 556 2556 564 2564
rect 668 2556 676 2564
rect 844 2556 852 2564
rect 1276 2556 1284 2564
rect 1324 2556 1332 2564
rect 1420 2556 1428 2564
rect 1692 2556 1700 2564
rect 1724 2556 1732 2564
rect 348 2536 356 2544
rect 732 2536 740 2544
rect 892 2536 900 2544
rect 1020 2536 1028 2544
rect 1116 2536 1124 2544
rect 1916 2536 1924 2544
rect 2876 2536 2884 2544
rect 3036 2536 3044 2544
rect 3052 2536 3060 2544
rect 3468 2536 3476 2544
rect 3756 2536 3764 2544
rect 3772 2536 3780 2544
rect 1836 2516 1844 2524
rect 1964 2516 1972 2524
rect 2108 2516 2116 2524
rect 2348 2516 2356 2524
rect 2540 2516 2548 2524
rect 2764 2516 2772 2524
rect 44 2496 52 2504
rect 396 2496 404 2504
rect 492 2496 500 2504
rect 540 2496 548 2504
rect 1132 2496 1140 2504
rect 1404 2496 1412 2504
rect 1516 2496 1524 2504
rect 1580 2496 1588 2504
rect 1676 2496 1684 2504
rect 2236 2496 2244 2504
rect 2316 2496 2324 2504
rect 2364 2496 2372 2504
rect 2700 2496 2708 2504
rect 2716 2496 2724 2504
rect 3084 2496 3092 2504
rect 3196 2496 3204 2504
rect 3500 2496 3508 2504
rect 3612 2496 3620 2504
rect 3788 2496 3796 2504
rect 3820 2496 3828 2504
rect 4140 2496 4148 2504
rect 4220 2496 4228 2504
rect 1804 2476 1812 2484
rect 1820 2456 1828 2464
rect 3308 2456 3316 2464
rect 3324 2456 3332 2464
rect 3852 2436 3860 2444
rect 764 2396 772 2404
rect 1148 2376 1156 2384
rect 2012 2376 2020 2384
rect 3996 2376 4004 2384
rect 268 2356 276 2364
rect 620 2356 628 2364
rect 1020 2356 1028 2364
rect 1436 2356 1444 2364
rect 1612 2356 1620 2364
rect 1884 2356 1892 2364
rect 2268 2356 2276 2364
rect 2892 2356 2900 2364
rect 3100 2356 3108 2364
rect 3676 2356 3684 2364
rect 220 2336 228 2344
rect 1324 2336 1332 2344
rect 2092 2336 2100 2344
rect 2860 2336 2868 2344
rect 2940 2336 2948 2344
rect 76 2316 84 2324
rect 156 2316 164 2324
rect 364 2316 372 2324
rect 588 2316 596 2324
rect 1004 2316 1012 2324
rect 1084 2316 1092 2324
rect 1196 2316 1204 2324
rect 1548 2316 1556 2324
rect 2588 2316 2596 2324
rect 3868 2316 3876 2324
rect 3948 2316 3956 2324
rect 4108 2316 4116 2324
rect 220 2296 228 2304
rect 380 2296 388 2304
rect 332 2276 340 2284
rect 460 2276 468 2284
rect 588 2276 596 2284
rect 2092 2276 2100 2284
rect 2124 2276 2132 2284
rect 2140 2276 2148 2284
rect 2316 2276 2324 2284
rect 2348 2276 2356 2284
rect 2412 2276 2420 2284
rect 188 2256 196 2264
rect 428 2256 436 2264
rect 492 2256 500 2264
rect 556 2256 564 2264
rect 1020 2256 1028 2264
rect 1452 2256 1460 2264
rect 1484 2256 1492 2264
rect 1676 2256 1684 2264
rect 1836 2256 1844 2264
rect 1900 2256 1908 2264
rect 1996 2256 2004 2264
rect 3068 2256 3076 2264
rect 3948 2256 3956 2264
rect 4028 2256 4036 2264
rect 4188 2256 4196 2264
rect 1292 2236 1300 2244
rect 1356 2236 1364 2244
rect 1516 2236 1524 2244
rect 1740 2236 1748 2244
rect 1756 2236 1764 2244
rect 2556 2236 2564 2244
rect 2588 2236 2596 2244
rect 2684 2236 2692 2244
rect 2796 2236 2804 2244
rect 3228 2236 3236 2244
rect 3548 2236 3556 2244
rect 3564 2236 3572 2244
rect 3580 2236 3588 2244
rect 1340 2216 1348 2224
rect 1708 2216 1716 2224
rect 2300 2216 2308 2224
rect 252 2196 260 2204
rect 2364 2196 2372 2204
rect 2844 2196 2852 2204
rect 3820 2196 3828 2204
rect 4012 2196 4020 2204
rect 844 2176 852 2184
rect 988 2176 996 2184
rect 1020 2176 1028 2184
rect 1084 2176 1092 2184
rect 1212 2176 1220 2184
rect 1308 2176 1316 2184
rect 1324 2176 1332 2184
rect 1436 2176 1444 2184
rect 1756 2176 1764 2184
rect 1772 2176 1780 2184
rect 1852 2176 1860 2184
rect 1932 2176 1940 2184
rect 1964 2176 1972 2184
rect 3564 2176 3572 2184
rect 4028 2176 4036 2184
rect 4092 2176 4100 2184
rect 28 2156 36 2164
rect 60 2156 68 2164
rect 252 2156 260 2164
rect 540 2156 548 2164
rect 1676 2156 1684 2164
rect 1708 2156 1716 2164
rect 1788 2156 1796 2164
rect 1804 2156 1812 2164
rect 1836 2156 1844 2164
rect 1916 2156 1924 2164
rect 2028 2156 2036 2164
rect 2556 2156 2564 2164
rect 3692 2156 3700 2164
rect 3916 2156 3924 2164
rect 60 2136 68 2144
rect 92 2136 100 2144
rect 428 2136 436 2144
rect 1068 2136 1076 2144
rect 1180 2136 1188 2144
rect 1292 2136 1300 2144
rect 1388 2136 1396 2144
rect 1500 2136 1508 2144
rect 3580 2136 3588 2144
rect 3596 2136 3604 2144
rect 3660 2136 3668 2144
rect 3804 2136 3812 2144
rect 3916 2136 3924 2144
rect 3964 2136 3972 2144
rect 4060 2136 4068 2144
rect 284 2116 292 2124
rect 348 2116 356 2124
rect 476 2116 484 2124
rect 780 2116 788 2124
rect 828 2116 836 2124
rect 876 2116 884 2124
rect 1052 2116 1060 2124
rect 1196 2116 1204 2124
rect 1308 2116 1316 2124
rect 1580 2116 1588 2124
rect 2380 2116 2388 2124
rect 3580 2116 3588 2124
rect 3804 2116 3812 2124
rect 284 2096 292 2104
rect 316 2096 324 2104
rect 556 2096 564 2104
rect 812 2096 820 2104
rect 860 2096 868 2104
rect 2796 2096 2804 2104
rect 2908 2096 2916 2104
rect 2956 2096 2964 2104
rect 3100 2096 3108 2104
rect 3500 2096 3508 2104
rect 3964 2096 3972 2104
rect 3996 2096 4004 2104
rect 4044 2096 4052 2104
rect 4172 2096 4180 2104
rect 4204 2096 4212 2104
rect 1020 2076 1028 2084
rect 1740 2076 1748 2084
rect 2092 2076 2100 2084
rect 2236 2076 2244 2084
rect 2588 2076 2596 2084
rect 2652 2076 2660 2084
rect 764 2056 772 2064
rect 1708 2056 1716 2064
rect 2940 2056 2948 2064
rect 3580 2056 3588 2064
rect 876 2036 884 2044
rect 1484 2036 1492 2044
rect 1628 2036 1636 2044
rect 3020 2036 3028 2044
rect 1692 2016 1700 2024
rect 2124 2016 2132 2024
rect 236 1996 244 2004
rect 2412 1996 2420 2004
rect 348 1976 356 1984
rect 732 1976 740 1984
rect 316 1956 324 1964
rect 1740 1956 1748 1964
rect 2124 1956 2132 1964
rect 2364 1956 2372 1964
rect 3452 1956 3460 1964
rect 3596 1956 3604 1964
rect 908 1936 916 1944
rect 1484 1936 1492 1944
rect 1564 1936 1572 1944
rect 2588 1936 2596 1944
rect 3724 1936 3732 1944
rect 540 1916 548 1924
rect 716 1916 724 1924
rect 828 1916 836 1924
rect 876 1916 884 1924
rect 1884 1916 1892 1924
rect 2412 1916 2420 1924
rect 2428 1916 2436 1924
rect 2460 1916 2468 1924
rect 2476 1916 2484 1924
rect 3308 1916 3316 1924
rect 3340 1916 3348 1924
rect 3548 1916 3556 1924
rect 3868 1916 3876 1924
rect 124 1896 132 1904
rect 140 1896 148 1904
rect 3260 1896 3268 1904
rect 12 1876 20 1884
rect 44 1876 52 1884
rect 508 1876 516 1884
rect 940 1876 948 1884
rect 1036 1876 1044 1884
rect 1164 1876 1172 1884
rect 1180 1876 1188 1884
rect 1196 1876 1204 1884
rect 1228 1876 1236 1884
rect 1308 1876 1316 1884
rect 1356 1876 1364 1884
rect 1388 1876 1396 1884
rect 1660 1876 1668 1884
rect 1820 1876 1828 1884
rect 1836 1876 1844 1884
rect 1900 1876 1908 1884
rect 2012 1876 2020 1884
rect 2492 1876 2500 1884
rect 2620 1876 2628 1884
rect 2636 1876 2644 1884
rect 3004 1876 3012 1884
rect 3052 1876 3060 1884
rect 3516 1876 3524 1884
rect 3580 1876 3588 1884
rect 4156 1876 4164 1884
rect 4220 1876 4228 1884
rect 28 1856 36 1864
rect 1116 1856 1124 1864
rect 2924 1856 2932 1864
rect 3292 1856 3300 1864
rect 3308 1856 3316 1864
rect 3980 1856 3988 1864
rect 4044 1856 4052 1864
rect 380 1836 388 1844
rect 716 1836 724 1844
rect 1244 1836 1252 1844
rect 1404 1836 1412 1844
rect 1452 1836 1460 1844
rect 2140 1836 2148 1844
rect 2156 1836 2164 1844
rect 2220 1836 2228 1844
rect 2300 1836 2308 1844
rect 2732 1836 2740 1844
rect 3660 1836 3668 1844
rect 780 1816 788 1824
rect 1692 1816 1700 1824
rect 2460 1816 2468 1824
rect 284 1796 292 1804
rect 1676 1796 1684 1804
rect 2380 1796 2388 1804
rect 3388 1796 3396 1804
rect 12 1776 20 1784
rect 1356 1776 1364 1784
rect 1740 1776 1748 1784
rect 1916 1776 1924 1784
rect 3100 1776 3108 1784
rect 316 1756 324 1764
rect 332 1756 340 1764
rect 508 1756 516 1764
rect 780 1756 788 1764
rect 828 1756 836 1764
rect 860 1756 868 1764
rect 972 1756 980 1764
rect 1052 1756 1060 1764
rect 1100 1756 1108 1764
rect 1180 1756 1188 1764
rect 1196 1756 1204 1764
rect 1292 1756 1300 1764
rect 1948 1756 1956 1764
rect 2300 1756 2308 1764
rect 2316 1756 2324 1764
rect 2460 1756 2468 1764
rect 2524 1756 2532 1764
rect 2556 1756 2564 1764
rect 2716 1756 2724 1764
rect 2796 1756 2804 1764
rect 2860 1756 2868 1764
rect 3500 1756 3508 1764
rect 3628 1756 3636 1764
rect 3772 1756 3780 1764
rect 3868 1756 3876 1764
rect 3884 1756 3892 1764
rect 4012 1756 4020 1764
rect 4044 1756 4052 1764
rect 236 1736 244 1744
rect 492 1736 500 1744
rect 1596 1736 1604 1744
rect 1612 1736 1620 1744
rect 1852 1736 1860 1744
rect 1900 1736 1908 1744
rect 2204 1736 2212 1744
rect 2588 1736 2596 1744
rect 2748 1736 2756 1744
rect 3164 1736 3172 1744
rect 3980 1736 3988 1744
rect 4028 1736 4036 1744
rect 924 1716 932 1724
rect 1660 1716 1668 1724
rect 2156 1716 2164 1724
rect 3244 1716 3252 1724
rect 3852 1716 3860 1724
rect 1212 1696 1220 1704
rect 1772 1696 1780 1704
rect 2172 1696 2180 1704
rect 2252 1696 2260 1704
rect 2620 1696 2628 1704
rect 3036 1696 3044 1704
rect 3116 1696 3124 1704
rect 3676 1696 3684 1704
rect 3708 1696 3716 1704
rect 4076 1696 4084 1704
rect 764 1676 772 1684
rect 1932 1676 1940 1684
rect 1948 1676 1956 1684
rect 3340 1676 3348 1684
rect 2284 1656 2292 1664
rect 3388 1656 3396 1664
rect 3788 1656 3796 1664
rect 812 1636 820 1644
rect 4092 1636 4100 1644
rect 780 1616 788 1624
rect 1196 1616 1204 1624
rect 2364 1616 2372 1624
rect 3516 1616 3524 1624
rect 4172 1616 4180 1624
rect 2428 1596 2436 1604
rect 172 1576 180 1584
rect 1324 1576 1332 1584
rect 1484 1576 1492 1584
rect 4124 1576 4132 1584
rect 236 1556 244 1564
rect 508 1556 516 1564
rect 860 1556 868 1564
rect 1340 1556 1348 1564
rect 1692 1556 1700 1564
rect 3068 1556 3076 1564
rect 3596 1556 3604 1564
rect 3628 1556 3636 1564
rect 2396 1536 2404 1544
rect 2572 1536 2580 1544
rect 3724 1536 3732 1544
rect 3964 1536 3972 1544
rect 524 1516 532 1524
rect 588 1516 596 1524
rect 620 1516 628 1524
rect 732 1516 740 1524
rect 892 1516 900 1524
rect 924 1516 932 1524
rect 1196 1516 1204 1524
rect 1244 1516 1252 1524
rect 2332 1516 2340 1524
rect 2348 1516 2356 1524
rect 2396 1516 2404 1524
rect 2652 1516 2660 1524
rect 2892 1516 2900 1524
rect 2940 1516 2948 1524
rect 3164 1516 3172 1524
rect 3436 1516 3444 1524
rect 4060 1516 4068 1524
rect 4092 1516 4100 1524
rect 4172 1516 4180 1524
rect 4220 1516 4228 1524
rect 4252 1516 4260 1524
rect 1404 1496 1412 1504
rect 156 1476 164 1484
rect 188 1476 196 1484
rect 300 1476 308 1484
rect 588 1476 596 1484
rect 684 1476 692 1484
rect 924 1476 932 1484
rect 956 1476 964 1484
rect 1132 1476 1140 1484
rect 1580 1476 1588 1484
rect 1692 1476 1700 1484
rect 2012 1476 2020 1484
rect 2076 1476 2084 1484
rect 2268 1476 2276 1484
rect 2460 1476 2468 1484
rect 2508 1476 2516 1484
rect 2588 1476 2596 1484
rect 2604 1476 2612 1484
rect 2716 1476 2724 1484
rect 3516 1476 3524 1484
rect 3580 1476 3588 1484
rect 3756 1476 3764 1484
rect 3996 1476 4004 1484
rect 76 1456 84 1464
rect 108 1456 116 1464
rect 412 1456 420 1464
rect 620 1456 628 1464
rect 1532 1456 1540 1464
rect 1628 1456 1636 1464
rect 1788 1456 1796 1464
rect 2492 1456 2500 1464
rect 2540 1456 2548 1464
rect 2684 1456 2692 1464
rect 3020 1456 3028 1464
rect 3964 1456 3972 1464
rect 4092 1456 4100 1464
rect 4188 1456 4196 1464
rect 332 1436 340 1444
rect 652 1436 660 1444
rect 828 1436 836 1444
rect 1116 1436 1124 1444
rect 1212 1436 1220 1444
rect 1372 1436 1380 1444
rect 2092 1436 2100 1444
rect 2220 1436 2228 1444
rect 2396 1436 2404 1444
rect 2780 1436 2788 1444
rect 2828 1436 2836 1444
rect 3628 1436 3636 1444
rect 3708 1436 3716 1444
rect 4156 1436 4164 1444
rect 1356 1416 1364 1424
rect 1724 1416 1732 1424
rect 1756 1416 1764 1424
rect 2572 1416 2580 1424
rect 2892 1416 2900 1424
rect 3580 1416 3588 1424
rect 2028 1396 2036 1404
rect 2076 1396 2084 1404
rect 3532 1396 3540 1404
rect 3548 1396 3556 1404
rect 844 1376 852 1384
rect 1068 1376 1076 1384
rect 1308 1376 1316 1384
rect 1324 1376 1332 1384
rect 1452 1376 1460 1384
rect 2140 1376 2148 1384
rect 2172 1376 2180 1384
rect 2316 1376 2324 1384
rect 2348 1376 2356 1384
rect 2412 1376 2420 1384
rect 2508 1376 2516 1384
rect 2812 1376 2820 1384
rect 2956 1376 2964 1384
rect 3004 1376 3012 1384
rect 3052 1376 3060 1384
rect 3100 1376 3108 1384
rect 3212 1376 3220 1384
rect 3228 1376 3236 1384
rect 3244 1376 3252 1384
rect 3340 1376 3348 1384
rect 3692 1376 3700 1384
rect 3852 1376 3860 1384
rect 3980 1376 3988 1384
rect 4044 1376 4052 1384
rect 108 1356 116 1364
rect 140 1356 148 1364
rect 380 1356 388 1364
rect 396 1356 404 1364
rect 460 1356 468 1364
rect 492 1356 500 1364
rect 732 1356 740 1364
rect 764 1356 772 1364
rect 1020 1356 1028 1364
rect 1516 1356 1524 1364
rect 1564 1356 1572 1364
rect 1580 1356 1588 1364
rect 1820 1356 1828 1364
rect 2316 1356 2324 1364
rect 2588 1356 2596 1364
rect 2956 1356 2964 1364
rect 3132 1356 3140 1364
rect 3772 1356 3780 1364
rect 3884 1356 3892 1364
rect 4124 1356 4132 1364
rect 4156 1356 4164 1364
rect 4204 1356 4212 1364
rect 44 1336 52 1344
rect 364 1336 372 1344
rect 540 1336 548 1344
rect 588 1336 596 1344
rect 748 1336 756 1344
rect 1020 1336 1028 1344
rect 1404 1336 1412 1344
rect 1692 1336 1700 1344
rect 1804 1336 1812 1344
rect 2188 1336 2196 1344
rect 2284 1336 2292 1344
rect 2876 1336 2884 1344
rect 3820 1336 3828 1344
rect 956 1296 964 1304
rect 1004 1296 1012 1304
rect 1068 1296 1076 1304
rect 1388 1296 1396 1304
rect 1932 1296 1940 1304
rect 2012 1296 2020 1304
rect 2028 1296 2036 1304
rect 2540 1296 2548 1304
rect 2668 1296 2676 1304
rect 2796 1296 2804 1304
rect 3260 1296 3268 1304
rect 3468 1296 3476 1304
rect 3772 1296 3780 1304
rect 3788 1296 3796 1304
rect 3900 1296 3908 1304
rect 3948 1296 3956 1304
rect 3996 1296 4004 1304
rect 2252 1256 2260 1264
rect 3164 1256 3172 1264
rect 988 1236 996 1244
rect 1740 1236 1748 1244
rect 2060 1236 2068 1244
rect 3644 1216 3652 1224
rect 1180 1176 1188 1184
rect 2316 1176 2324 1184
rect 2892 1176 2900 1184
rect 3724 1176 3732 1184
rect 1596 1156 1604 1164
rect 2092 1156 2100 1164
rect 3452 1156 3460 1164
rect 3852 1156 3860 1164
rect 4188 1156 4196 1164
rect 652 1136 660 1144
rect 716 1136 724 1144
rect 1004 1136 1012 1144
rect 1660 1136 1668 1144
rect 1804 1136 1812 1144
rect 2012 1136 2020 1144
rect 2140 1136 2148 1144
rect 2396 1136 2404 1144
rect 4044 1136 4052 1144
rect 236 1116 244 1124
rect 332 1116 340 1124
rect 1100 1116 1108 1124
rect 1276 1116 1284 1124
rect 1324 1116 1332 1124
rect 1820 1116 1828 1124
rect 2636 1116 2644 1124
rect 2764 1116 2772 1124
rect 2796 1116 2804 1124
rect 2876 1116 2884 1124
rect 2940 1116 2948 1124
rect 2988 1116 2996 1124
rect 3084 1116 3092 1124
rect 3132 1116 3140 1124
rect 3404 1116 3412 1124
rect 3436 1116 3444 1124
rect 3996 1116 4004 1124
rect 4220 1116 4228 1124
rect 604 1096 612 1104
rect 652 1096 660 1104
rect 2956 1096 2964 1104
rect 76 1076 84 1084
rect 284 1076 292 1084
rect 316 1076 324 1084
rect 364 1076 372 1084
rect 732 1076 740 1084
rect 812 1076 820 1084
rect 1132 1076 1140 1084
rect 1660 1076 1668 1084
rect 1852 1076 1860 1084
rect 1964 1076 1972 1084
rect 2620 1076 2628 1084
rect 2668 1076 2676 1084
rect 2828 1076 2836 1084
rect 3084 1076 3092 1084
rect 3676 1076 3684 1084
rect 3820 1076 3828 1084
rect 3836 1076 3844 1084
rect 4012 1076 4020 1084
rect 4108 1076 4116 1084
rect 92 1056 100 1064
rect 140 1056 148 1064
rect 380 1056 388 1064
rect 524 1056 532 1064
rect 1212 1056 1220 1064
rect 1244 1056 1252 1064
rect 1468 1056 1476 1064
rect 1516 1056 1524 1064
rect 1596 1056 1604 1064
rect 1724 1056 1732 1064
rect 1772 1056 1780 1064
rect 1868 1056 1876 1064
rect 2476 1056 2484 1064
rect 2572 1056 2580 1064
rect 2684 1056 2692 1064
rect 2924 1056 2932 1064
rect 3068 1056 3076 1064
rect 3100 1056 3108 1064
rect 92 1036 100 1044
rect 428 1036 436 1044
rect 716 1036 724 1044
rect 780 1036 788 1044
rect 796 1036 804 1044
rect 844 1036 852 1044
rect 956 1036 964 1044
rect 972 1036 980 1044
rect 2076 1036 2084 1044
rect 2716 1036 2724 1044
rect 3148 1036 3156 1044
rect 3484 1036 3492 1044
rect 3580 1036 3588 1044
rect 3996 1036 4004 1044
rect 1644 1016 1652 1024
rect 588 996 596 1004
rect 2860 996 2868 1004
rect 3532 996 3540 1004
rect 4172 996 4180 1004
rect 124 976 132 984
rect 444 976 452 984
rect 780 976 788 984
rect 828 976 836 984
rect 988 976 996 984
rect 1244 976 1252 984
rect 1356 976 1364 984
rect 2972 976 2980 984
rect 3036 976 3044 984
rect 3084 976 3092 984
rect 3308 976 3316 984
rect 3324 976 3332 984
rect 3644 976 3652 984
rect 3948 976 3956 984
rect 4044 976 4052 984
rect 4204 976 4212 984
rect 124 956 132 964
rect 156 956 164 964
rect 300 956 308 964
rect 364 956 372 964
rect 428 956 436 964
rect 460 956 468 964
rect 492 956 500 964
rect 1276 956 1284 964
rect 1356 956 1364 964
rect 2412 956 2420 964
rect 2444 956 2452 964
rect 3660 956 3668 964
rect 3980 956 3988 964
rect 4108 956 4116 964
rect 236 936 244 944
rect 1740 936 1748 944
rect 1948 936 1956 944
rect 2092 936 2100 944
rect 2124 936 2132 944
rect 2188 936 2196 944
rect 2220 936 2228 944
rect 2300 936 2308 944
rect 2364 936 2372 944
rect 2460 936 2468 944
rect 2620 936 2628 944
rect 2860 936 2868 944
rect 3772 936 3780 944
rect 3804 936 3812 944
rect 3884 936 3892 944
rect 4028 936 4036 944
rect 4060 936 4068 944
rect 4092 936 4100 944
rect 60 916 68 924
rect 1292 916 1300 924
rect 2044 916 2052 924
rect 2252 916 2260 924
rect 2428 916 2436 924
rect 2988 916 2996 924
rect 3356 916 3364 924
rect 92 896 100 904
rect 396 896 404 904
rect 668 896 676 904
rect 764 896 772 904
rect 972 896 980 904
rect 1244 896 1252 904
rect 1260 896 1268 904
rect 1276 896 1284 904
rect 1484 896 1492 904
rect 1612 896 1620 904
rect 1980 896 1988 904
rect 2028 896 2036 904
rect 2572 896 2580 904
rect 2652 896 2660 904
rect 2684 896 2692 904
rect 2940 896 2948 904
rect 3020 896 3028 904
rect 3196 896 3204 904
rect 3420 896 3428 904
rect 3596 896 3604 904
rect 3612 896 3620 904
rect 3644 896 3652 904
rect 4028 896 4036 904
rect 1692 876 1700 884
rect 2828 876 2836 884
rect 3452 876 3460 884
rect 3628 876 3636 884
rect 1516 856 1524 864
rect 1100 816 1108 824
rect 2524 816 2532 824
rect 428 776 436 784
rect 892 776 900 784
rect 1676 776 1684 784
rect 668 756 676 764
rect 1068 756 1076 764
rect 1692 756 1700 764
rect 2572 756 2580 764
rect 1292 736 1300 744
rect 1772 736 1780 744
rect 1852 736 1860 744
rect 1932 736 1940 744
rect 2188 736 2196 744
rect 2236 736 2244 744
rect 2300 736 2308 744
rect 3500 736 3508 744
rect 508 716 516 724
rect 1068 716 1076 724
rect 1116 716 1124 724
rect 2156 716 2164 724
rect 2412 716 2420 724
rect 2460 716 2468 724
rect 2764 716 2772 724
rect 2956 716 2964 724
rect 2988 716 2996 724
rect 3020 716 3028 724
rect 3052 716 3060 724
rect 3868 716 3876 724
rect 3948 716 3956 724
rect 4188 716 4196 724
rect 364 696 372 704
rect 732 696 740 704
rect 1084 696 1092 704
rect 1260 696 1268 704
rect 2924 696 2932 704
rect 156 676 164 684
rect 236 676 244 684
rect 604 676 612 684
rect 1452 676 1460 684
rect 1612 676 1620 684
rect 1836 676 1844 684
rect 1964 676 1972 684
rect 2188 676 2196 684
rect 2716 676 2724 684
rect 3132 676 3140 684
rect 3308 676 3316 684
rect 3628 676 3636 684
rect 3676 676 3684 684
rect 4108 676 4116 684
rect 4156 676 4164 684
rect 108 656 116 664
rect 220 656 228 664
rect 412 656 420 664
rect 652 656 660 664
rect 860 656 868 664
rect 2012 656 2020 664
rect 2060 656 2068 664
rect 2236 656 2244 664
rect 3516 656 3524 664
rect 3532 656 3540 664
rect 3548 656 3556 664
rect 3676 656 3684 664
rect 3740 656 3748 664
rect 3852 656 3860 664
rect 4076 656 4084 664
rect 4108 656 4116 664
rect 1532 636 1540 644
rect 1916 636 1924 644
rect 2300 636 2308 644
rect 2460 636 2468 644
rect 2684 636 2692 644
rect 2732 636 2740 644
rect 2876 636 2884 644
rect 3356 636 3364 644
rect 3404 636 3412 644
rect 684 616 692 624
rect 1916 616 1924 624
rect 1340 596 1348 604
rect 1404 596 1412 604
rect 2732 596 2740 604
rect 4028 596 4036 604
rect 284 576 292 584
rect 2012 576 2020 584
rect 2220 576 2228 584
rect 3036 576 3044 584
rect 3260 576 3268 584
rect 3324 576 3332 584
rect 3356 576 3364 584
rect 3372 576 3380 584
rect 364 556 372 564
rect 604 556 612 564
rect 620 556 628 564
rect 716 556 724 564
rect 812 556 820 564
rect 1020 556 1028 564
rect 1388 556 1396 564
rect 1548 556 1556 564
rect 1644 556 1652 564
rect 1916 556 1924 564
rect 1980 556 1988 564
rect 1996 556 2004 564
rect 2428 556 2436 564
rect 2508 556 2516 564
rect 2748 556 2756 564
rect 3516 556 3524 564
rect 3852 556 3860 564
rect 92 536 100 544
rect 124 536 132 544
rect 268 536 276 544
rect 428 536 436 544
rect 460 536 468 544
rect 796 536 804 544
rect 844 536 852 544
rect 1212 536 1220 544
rect 1324 536 1332 544
rect 1420 536 1428 544
rect 1532 536 1540 544
rect 2524 536 2532 544
rect 2668 536 2676 544
rect 2780 536 2788 544
rect 3580 536 3588 544
rect 3676 536 3684 544
rect 3868 536 3876 544
rect 4028 536 4036 544
rect 4060 536 4068 544
rect 4076 536 4084 544
rect 1932 516 1940 524
rect 2844 516 2852 524
rect 3420 516 3428 524
rect 3468 516 3476 524
rect 3532 516 3540 524
rect 3756 516 3764 524
rect 188 496 196 504
rect 220 496 228 504
rect 284 496 292 504
rect 940 496 948 504
rect 972 496 980 504
rect 1596 496 1604 504
rect 2476 496 2484 504
rect 4076 496 4084 504
rect 364 476 372 484
rect 668 476 676 484
rect 1404 476 1412 484
rect 2284 476 2292 484
rect 2348 476 2356 484
rect 3324 476 3332 484
rect 2092 456 2100 464
rect 3244 456 3252 464
rect 252 416 260 424
rect 300 376 308 384
rect 1036 376 1044 384
rect 1740 376 1748 384
rect 2732 376 2740 384
rect 3148 376 3156 384
rect 3420 376 3428 384
rect 3452 376 3460 384
rect 3868 376 3876 384
rect 156 356 164 364
rect 364 356 372 364
rect 2044 356 2052 364
rect 3068 356 3076 364
rect 3388 356 3396 364
rect 3500 356 3508 364
rect 3612 356 3620 364
rect 812 336 820 344
rect 1004 336 1012 344
rect 1804 336 1812 344
rect 2092 336 2100 344
rect 2572 336 2580 344
rect 2956 336 2964 344
rect 3772 336 3780 344
rect 60 316 68 324
rect 652 316 660 324
rect 956 316 964 324
rect 1244 316 1252 324
rect 1260 316 1268 324
rect 1996 316 2004 324
rect 2764 316 2772 324
rect 2988 316 2996 324
rect 3212 316 3220 324
rect 3292 316 3300 324
rect 3436 316 3444 324
rect 3644 316 3652 324
rect 3708 316 3716 324
rect 1596 296 1604 304
rect 2204 296 2212 304
rect 2252 296 2260 304
rect 3916 296 3924 304
rect 284 276 292 284
rect 332 276 340 284
rect 700 276 708 284
rect 844 276 852 284
rect 1180 276 1188 284
rect 2764 276 2772 284
rect 2812 276 2820 284
rect 2940 276 2948 284
rect 2972 276 2980 284
rect 4124 276 4132 284
rect 396 256 404 264
rect 620 256 628 264
rect 780 256 788 264
rect 1308 256 1316 264
rect 1324 256 1332 264
rect 1500 256 1508 264
rect 2044 256 2052 264
rect 2444 256 2452 264
rect 2524 256 2532 264
rect 3164 256 3172 264
rect 3468 256 3476 264
rect 3596 256 3604 264
rect 3948 256 3956 264
rect 4140 256 4148 264
rect 1628 236 1636 244
rect 2092 236 2100 244
rect 2380 236 2388 244
rect 3324 236 3332 244
rect 3644 236 3652 244
rect 1004 216 1012 224
rect 2428 216 2436 224
rect 3004 216 3012 224
rect 3740 216 3748 224
rect 3804 216 3812 224
rect 1548 196 1556 204
rect 1580 196 1588 204
rect 1900 196 1908 204
rect 2684 196 2692 204
rect 4012 196 4020 204
rect 1612 176 1620 184
rect 1660 176 1668 184
rect 1772 176 1780 184
rect 1820 176 1828 184
rect 1836 176 1844 184
rect 1932 176 1940 184
rect 2044 176 2052 184
rect 2092 176 2100 184
rect 2636 176 2644 184
rect 2748 176 2756 184
rect 3580 176 3588 184
rect 4188 176 4196 184
rect 4204 176 4212 184
rect 92 156 100 164
rect 428 156 436 164
rect 2460 156 2468 164
rect 2524 156 2532 164
rect 2588 156 2596 164
rect 2844 156 2852 164
rect 2908 156 2916 164
rect 2956 156 2964 164
rect 3452 156 3460 164
rect 3516 156 3524 164
rect 3788 156 3796 164
rect 3948 156 3956 164
rect 92 136 100 144
rect 140 136 148 144
rect 780 136 788 144
rect 1132 136 1140 144
rect 1148 136 1156 144
rect 1196 136 1204 144
rect 1804 136 1812 144
rect 1836 136 1844 144
rect 2108 136 2116 144
rect 2300 136 2308 144
rect 2556 136 2564 144
rect 3036 136 3044 144
rect 3148 136 3156 144
rect 3180 136 3188 144
rect 3468 136 3476 144
rect 3692 136 3700 144
rect 540 116 548 124
rect 2556 116 2564 124
rect 3452 116 3460 124
rect 3676 116 3684 124
rect 4188 116 4196 124
rect 44 96 52 104
rect 124 96 132 104
rect 396 96 404 104
rect 1052 96 1060 104
rect 1100 96 1108 104
rect 1116 96 1124 104
rect 1564 96 1572 104
rect 1756 96 1764 104
rect 1996 96 2004 104
rect 2204 96 2212 104
rect 2252 96 2260 104
rect 2796 96 2804 104
rect 2956 96 2964 104
rect 3036 96 3044 104
rect 3084 96 3092 104
rect 3164 96 3172 104
rect 3820 96 3828 104
rect 3852 96 3860 104
rect 4140 96 4148 104
rect 892 76 900 84
rect 1164 76 1172 84
rect 1212 76 1220 84
rect 1532 76 1540 84
rect 1804 76 1812 84
rect 2012 76 2020 84
rect 2156 76 2164 84
rect 3052 56 3060 64
rect 2876 16 2884 24
<< metal1 >>
rect -412 3004 8 3016
rect -412 2616 -312 3004
rect 586 2976 588 2984
rect 858 2976 860 2984
rect 2868 2976 2870 2984
rect 68 2957 99 2963
rect 324 2957 355 2963
rect 644 2957 675 2963
rect 788 2957 819 2963
rect 980 2956 988 2964
rect 1092 2956 1100 2964
rect 1220 2957 1251 2963
rect 1293 2957 1324 2963
rect 1604 2956 1612 2964
rect 1876 2957 1907 2963
rect 1949 2957 1980 2963
rect 2020 2956 2028 2964
rect 2212 2956 2220 2964
rect 2404 2956 2412 2964
rect 2461 2957 2492 2963
rect 2589 2957 2620 2963
rect 29 2937 51 2943
rect 173 2937 195 2943
rect 285 2937 307 2943
rect 397 2937 428 2943
rect 612 2937 627 2943
rect 829 2937 844 2943
rect 1037 2937 1075 2943
rect 1181 2937 1203 2943
rect 1341 2937 1363 2943
rect 1453 2937 1491 2943
rect 1629 2937 1667 2943
rect 445 2917 460 2923
rect 749 2917 764 2923
rect 1853 2923 1859 2943
rect 2173 2937 2195 2943
rect 2260 2937 2275 2943
rect 2349 2937 2364 2943
rect 2749 2943 2755 2963
rect 2772 2956 2780 2964
rect 2932 2956 2940 2964
rect 2653 2937 2691 2943
rect 2749 2937 2764 2943
rect 3053 2943 3059 2963
rect 3092 2957 3123 2963
rect 3325 2957 3356 2963
rect 3405 2957 3436 2963
rect 3757 2957 3788 2963
rect 3869 2957 3900 2963
rect 3053 2937 3068 2943
rect 1101 2917 1139 2923
rect 1821 2917 1859 2923
rect 2285 2917 2323 2923
rect 77 2897 92 2903
rect 1101 2897 1107 2917
rect 1636 2897 1651 2903
rect 1716 2897 1731 2903
rect 2221 2897 2243 2903
rect 2317 2897 2323 2917
rect 2381 2917 2396 2923
rect 3229 2923 3235 2943
rect 3197 2917 3235 2923
rect 3453 2923 3459 2943
rect 3597 2937 3619 2943
rect 3805 2937 3827 2943
rect 3917 2937 3939 2943
rect 4029 2937 4051 2943
rect 4109 2937 4131 2943
rect 4221 2937 4268 2943
rect 3453 2917 3491 2923
rect 3540 2917 3555 2923
rect 2756 2897 2771 2903
rect 2877 2897 2892 2903
rect 2909 2897 2931 2903
rect 3101 2897 3116 2903
rect 3693 2897 3708 2903
rect 3844 2897 3859 2903
rect 100 2877 115 2883
rect 548 2877 563 2883
rect 924 2883 932 2888
rect 708 2877 723 2883
rect 924 2877 947 2883
rect 1780 2877 1795 2883
rect 3037 2877 3052 2883
rect 3309 2877 3324 2883
rect 3772 2883 3780 2888
rect 3996 2883 4004 2888
rect 4188 2883 4196 2888
rect 3764 2877 3780 2883
rect 3981 2877 4004 2883
rect 4173 2877 4196 2883
rect 4582 2816 4682 3016
rect 4242 2804 4682 2816
rect 44 2737 67 2743
rect 44 2732 52 2737
rect 1581 2737 1604 2743
rect 1613 2737 1628 2743
rect 1596 2732 1604 2737
rect 1884 2737 1907 2743
rect 2364 2737 2387 2743
rect 1884 2732 1892 2737
rect 2364 2732 2372 2737
rect 2588 2737 2611 2743
rect 3100 2737 3123 2743
rect 3341 2737 3364 2743
rect 2588 2732 2596 2737
rect 3100 2732 3108 2737
rect 3356 2732 3364 2737
rect 109 2717 124 2723
rect 420 2717 435 2723
rect 1108 2717 1123 2723
rect 1277 2717 1292 2723
rect 1364 2717 1379 2723
rect 2029 2717 2051 2723
rect 2797 2717 2835 2723
rect 3021 2717 3043 2723
rect 3140 2717 3155 2723
rect 3309 2717 3324 2723
rect 3741 2717 3756 2723
rect 3940 2717 3955 2723
rect 4029 2717 4044 2723
rect 365 2697 380 2703
rect 109 2677 131 2683
rect 189 2677 211 2683
rect 317 2677 332 2683
rect 365 2677 371 2697
rect 3076 2697 3091 2703
rect 3261 2697 3299 2703
rect 3965 2697 4003 2703
rect 461 2677 483 2683
rect 1069 2677 1091 2683
rect 1476 2677 1507 2683
rect 1629 2677 1651 2683
rect 1732 2677 1747 2683
rect 1837 2677 1859 2683
rect 1965 2677 1987 2683
rect 2116 2677 2147 2683
rect 2269 2677 2291 2683
rect 2669 2677 2691 2683
rect 2861 2677 2876 2683
rect 2909 2677 2931 2683
rect 2973 2677 2995 2683
rect 3060 2677 3075 2683
rect 3181 2677 3203 2683
rect 3261 2677 3267 2697
rect 3389 2677 3427 2683
rect 3508 2677 3523 2683
rect 3556 2677 3571 2683
rect 3997 2677 4003 2697
rect 228 2657 259 2663
rect 573 2657 604 2663
rect 788 2657 819 2663
rect 868 2656 876 2664
rect 1101 2657 1132 2663
rect 1389 2657 1420 2663
rect 2180 2656 2188 2664
rect 2836 2656 2844 2664
rect 3213 2657 3244 2663
rect 3364 2656 3372 2664
rect 3453 2657 3484 2663
rect 3581 2657 3612 2663
rect 3716 2656 3724 2664
rect 3757 2657 3788 2663
rect 4020 2657 4051 2663
rect 4100 2656 4108 2664
rect 4173 2657 4204 2663
rect 298 2636 300 2644
rect 346 2636 348 2644
rect 442 2636 444 2644
rect 682 2636 684 2644
rect 730 2636 732 2644
rect 1876 2636 1878 2644
rect 1946 2636 1948 2644
rect 2890 2636 2892 2644
rect 3162 2636 3164 2644
rect 3866 2636 3868 2644
rect -412 2604 34 2616
rect -412 2216 -312 2604
rect 532 2576 534 2584
rect 1156 2576 1158 2584
rect 1396 2576 1398 2584
rect 1466 2576 1468 2584
rect 2132 2576 2134 2584
rect 3108 2576 3110 2584
rect 3498 2576 3500 2584
rect 3924 2576 3926 2584
rect 4154 2576 4156 2584
rect 36 2557 67 2563
rect 116 2557 147 2563
rect 580 2557 611 2563
rect 685 2557 716 2563
rect 836 2557 867 2563
rect 1332 2556 1340 2564
rect 1572 2557 1603 2563
rect 2365 2557 2396 2563
rect 3380 2556 3388 2564
rect 3725 2557 3756 2563
rect 77 2537 99 2543
rect 189 2537 211 2543
rect 301 2537 323 2543
rect 356 2537 371 2543
rect 548 2537 563 2543
rect 877 2537 892 2543
rect 925 2537 963 2543
rect 973 2537 988 2543
rect 909 2517 940 2523
rect 1037 2523 1043 2543
rect 1213 2537 1235 2543
rect 1645 2537 1676 2543
rect 2045 2537 2083 2543
rect 2452 2537 2483 2543
rect 2637 2537 2659 2543
rect 2733 2537 2755 2543
rect 2813 2537 2851 2543
rect 2861 2537 2876 2543
rect 2996 2537 3011 2543
rect 3348 2537 3363 2543
rect 3428 2537 3459 2543
rect 3581 2537 3612 2543
rect 4013 2537 4035 2543
rect 1005 2517 1043 2523
rect 1069 2517 1107 2523
rect 1165 2517 1203 2523
rect 1949 2517 1964 2523
rect 237 2497 252 2503
rect 349 2497 364 2503
rect 1069 2497 1075 2517
rect 1165 2497 1171 2517
rect 2221 2517 2259 2523
rect 1309 2497 1331 2503
rect 1876 2497 1891 2503
rect 2004 2497 2019 2503
rect 2253 2497 2259 2517
rect 3229 2517 3267 2523
rect 2372 2497 2387 2503
rect 2772 2497 2787 2503
rect 3069 2497 3084 2503
rect 3261 2497 3267 2517
rect 3597 2517 3635 2523
rect 3597 2497 3603 2517
rect 3732 2497 3747 2503
rect 4077 2497 4099 2503
rect 1180 2484 1188 2488
rect 1773 2477 1804 2483
rect 2420 2477 2435 2483
rect 2572 2483 2580 2488
rect 2500 2477 2515 2483
rect 2572 2477 2595 2483
rect 3116 2483 3124 2488
rect 3932 2484 3940 2488
rect 2660 2477 2675 2483
rect 3116 2477 3139 2483
rect 3405 2477 3420 2483
rect 4582 2416 4682 2804
rect 4242 2404 4682 2416
rect 653 2337 676 2343
rect 668 2332 676 2337
rect 1309 2337 1324 2343
rect 1741 2337 1764 2343
rect 2061 2337 2092 2343
rect 1756 2332 1764 2337
rect 2396 2337 2412 2343
rect 2396 2332 2404 2337
rect 4173 2337 4196 2343
rect 573 2317 588 2323
rect 788 2317 803 2323
rect 813 2317 844 2323
rect 909 2317 924 2323
rect 349 2297 380 2303
rect 445 2297 460 2303
rect 685 2297 700 2303
rect 1213 2303 1219 2323
rect 1332 2317 1347 2323
rect 1709 2317 1724 2323
rect 1181 2297 1219 2303
rect 2013 2297 2044 2303
rect 2445 2303 2451 2323
rect 2637 2317 2652 2323
rect 2685 2317 2700 2323
rect 2733 2317 2748 2323
rect 3021 2323 3027 2336
rect 4188 2332 4196 2337
rect 3021 2317 3043 2323
rect 3124 2317 3139 2323
rect 3341 2317 3356 2323
rect 3549 2317 3564 2323
rect 3757 2317 3795 2323
rect 2173 2297 2211 2303
rect 2445 2297 2460 2303
rect 29 2277 51 2283
rect 109 2277 131 2283
rect 173 2277 204 2283
rect 701 2277 723 2283
rect 1085 2277 1107 2283
rect 1533 2277 1571 2283
rect 1844 2277 1859 2283
rect 1933 2277 1955 2283
rect 2173 2277 2179 2297
rect 2493 2297 2556 2303
rect 2333 2277 2371 2283
rect 2493 2277 2499 2297
rect 2605 2277 2611 2316
rect 3053 2297 3084 2303
rect 3213 2297 3228 2303
rect 2692 2277 2707 2283
rect 2973 2277 3011 2283
rect 3165 2277 3203 2283
rect 3213 2277 3219 2297
rect 3837 2297 3868 2303
rect 3885 2297 3923 2303
rect 3325 2277 3363 2283
rect 3469 2277 3491 2283
rect 3917 2277 3923 2297
rect 4221 2277 4243 2283
rect 484 2256 492 2264
rect 868 2257 899 2263
rect 1828 2256 1836 2264
rect 2148 2256 2156 2264
rect 2253 2257 2284 2263
rect 2788 2256 2796 2264
rect 2852 2257 2883 2263
rect 2925 2257 2956 2263
rect 3421 2257 3452 2263
rect 3661 2257 3692 2263
rect 3940 2256 3948 2264
rect 4196 2256 4204 2264
rect 68 2236 70 2244
rect 148 2236 150 2244
rect 260 2236 262 2244
rect 612 2236 614 2244
rect 762 2236 764 2244
rect 1306 2236 1308 2244
rect 1354 2236 1356 2244
rect 1514 2236 1516 2244
rect 1652 2236 1654 2244
rect 1972 2236 1974 2244
rect 2474 2236 2476 2244
rect 2628 2236 2630 2244
rect 3146 2236 3148 2244
rect 3380 2236 3382 2244
rect 3588 2236 3590 2244
rect 4074 2236 4076 2244
rect 4122 2236 4124 2244
rect -412 2204 12 2216
rect -412 1816 -312 2204
rect 852 2176 854 2184
rect 922 2176 924 2184
rect 1092 2176 1094 2184
rect 1236 2176 1238 2184
rect 1274 2176 1276 2184
rect 1444 2176 1446 2184
rect 1562 2176 1564 2184
rect 1684 2176 1686 2184
rect 2362 2176 2364 2184
rect 3098 2176 3100 2184
rect 452 2156 460 2164
rect 685 2157 716 2163
rect 1005 2157 1036 2163
rect 1492 2157 1523 2163
rect 1716 2156 1724 2164
rect 1828 2156 1836 2164
rect 2100 2157 2131 2163
rect 2669 2157 2700 2163
rect 3188 2157 3219 2163
rect 45 2137 60 2143
rect 477 2137 515 2143
rect 605 2137 643 2143
rect 1149 2137 1164 2143
rect 2045 2137 2083 2143
rect 2221 2137 2259 2143
rect 2717 2137 2732 2143
rect 2781 2137 2819 2143
rect 2957 2137 2979 2143
rect 3124 2137 3139 2143
rect 3277 2137 3299 2143
rect 3325 2143 3331 2163
rect 3380 2157 3411 2163
rect 3485 2157 3516 2163
rect 3748 2156 3756 2164
rect 3828 2157 3859 2163
rect 3908 2156 3916 2164
rect 3988 2157 4019 2163
rect 4196 2157 4227 2163
rect 3316 2137 3331 2143
rect 3533 2137 3555 2143
rect 292 2117 307 2123
rect 356 2117 371 2123
rect 797 2117 828 2123
rect 1588 2117 1603 2123
rect 2772 2117 2787 2123
rect 3789 2117 3804 2123
rect 4077 2123 4083 2143
rect 4077 2117 4115 2123
rect 324 2097 339 2103
rect 413 2097 451 2103
rect 484 2097 499 2103
rect 692 2097 707 2103
rect 1453 2097 1468 2103
rect 1533 2097 1555 2103
rect 2285 2097 2307 2103
rect 2340 2097 2355 2103
rect 2877 2097 2908 2103
rect 2980 2097 2995 2103
rect 3229 2097 3251 2103
rect 3949 2097 3964 2103
rect 4157 2097 4172 2103
rect 1100 2084 1108 2088
rect 260 2077 275 2083
rect 1756 2084 1764 2088
rect 2188 2083 2196 2088
rect 2173 2077 2196 2083
rect 2205 2077 2236 2083
rect 3004 2083 3012 2088
rect 2916 2077 2931 2083
rect 3004 2077 3027 2083
rect 3060 2077 3075 2083
rect 3860 2077 3875 2083
rect 4237 2037 4252 2043
rect 4582 2016 4682 2404
rect 4242 2004 4682 2016
rect 1260 1937 1283 1943
rect 1260 1932 1268 1937
rect 1492 1937 1507 1943
rect 1572 1937 1587 1943
rect 2020 1937 2035 1943
rect 205 1917 227 1923
rect 413 1917 435 1923
rect 621 1917 636 1923
rect 909 1917 931 1923
rect 1172 1917 1187 1923
rect 1421 1917 1443 1923
rect 1901 1917 1939 1923
rect 2093 1917 2108 1923
rect 132 1897 147 1903
rect 52 1877 67 1883
rect 141 1877 147 1897
rect 493 1897 531 1903
rect 861 1897 892 1903
rect 493 1877 499 1897
rect 2573 1903 2579 1923
rect 2733 1917 2755 1923
rect 2852 1917 2867 1923
rect 3165 1917 3180 1923
rect 3213 1917 3228 1923
rect 3453 1917 3468 1923
rect 3485 1917 3500 1923
rect 3629 1917 3667 1923
rect 4173 1917 4195 1923
rect 2573 1897 2611 1903
rect 2797 1897 2812 1903
rect 3245 1897 3260 1903
rect 573 1877 595 1883
rect 653 1877 691 1883
rect 1165 1877 1180 1883
rect 1965 1877 2003 1883
rect 2052 1877 2067 1883
rect 2356 1877 2371 1883
rect 2509 1877 2547 1883
rect 2557 1877 2588 1883
rect 2692 1877 2707 1883
rect 2973 1877 2995 1883
rect 3124 1877 3139 1883
rect 3412 1877 3427 1883
rect 3693 1877 3731 1883
rect 3757 1877 3795 1883
rect 3901 1877 3916 1883
rect 4029 1877 4067 1883
rect 4141 1877 4156 1883
rect 77 1857 108 1863
rect 1517 1857 1548 1863
rect 1940 1856 1948 1864
rect 2340 1856 2348 1864
rect 3204 1857 3235 1863
rect 3284 1856 3292 1864
rect 3444 1857 3475 1863
rect 3853 1857 3884 1863
rect 3940 1857 3971 1863
rect 4084 1856 4092 1864
rect 164 1836 166 1844
rect 234 1836 236 1844
rect 282 1836 284 1844
rect 474 1836 476 1844
rect 612 1836 614 1844
rect 660 1836 662 1844
rect 868 1836 870 1844
rect 1076 1836 1078 1844
rect 1146 1836 1148 1844
rect 1252 1836 1254 1844
rect 1322 1836 1324 1844
rect 1412 1836 1414 1844
rect 1994 1836 1996 1844
rect 2196 1836 2198 1844
rect 2388 1836 2390 1844
rect 2836 1836 2838 1844
rect 2874 1836 2876 1844
rect 3156 1836 3158 1844
rect 3322 1836 3324 1844
rect 4010 1836 4012 1844
rect 4202 1836 4204 1844
rect -412 1804 10 1816
rect -412 1416 -312 1804
rect 186 1776 188 1784
rect 554 1776 556 1784
rect 1924 1776 1926 1784
rect 2394 1776 2396 1784
rect 2692 1776 2694 1784
rect 2948 1776 2950 1784
rect 3108 1776 3110 1784
rect 3930 1776 3932 1784
rect 77 1757 108 1763
rect 356 1756 364 1764
rect 644 1757 675 1763
rect 1108 1756 1116 1764
rect 1300 1756 1308 1764
rect 1380 1756 1388 1764
rect 1437 1757 1468 1763
rect 1524 1757 1555 1763
rect 1677 1757 1708 1763
rect 1956 1756 1964 1764
rect 2013 1757 2044 1763
rect 2244 1757 2275 1763
rect 2468 1756 2476 1764
rect 2612 1757 2643 1763
rect 2804 1756 2812 1764
rect 4205 1757 4236 1763
rect 45 1737 67 1743
rect 244 1737 259 1743
rect 381 1737 403 1743
rect 573 1737 588 1743
rect 605 1737 627 1743
rect 765 1737 787 1743
rect 1053 1737 1075 1743
rect 1245 1737 1267 1743
rect 1773 1737 1811 1743
rect 1860 1737 1875 1743
rect 1981 1737 2003 1743
rect 2333 1737 2348 1743
rect 2653 1737 2675 1743
rect 2733 1737 2748 1743
rect 2868 1737 2899 1743
rect 3076 1737 3091 1743
rect 3453 1737 3475 1743
rect 3517 1737 3532 1743
rect 3741 1737 3763 1743
rect 3949 1737 3971 1743
rect 3988 1737 4003 1743
rect 1005 1717 1043 1723
rect 157 1697 179 1703
rect 525 1697 547 1703
rect 653 1697 668 1703
rect 877 1697 899 1703
rect 1005 1697 1011 1717
rect 2164 1717 2195 1723
rect 3181 1717 3219 1723
rect 2477 1697 2515 1703
rect 2701 1697 2716 1703
rect 3213 1697 3219 1717
rect 3661 1697 3676 1703
rect 3901 1697 3923 1703
rect 460 1683 468 1688
rect 732 1683 740 1688
rect 276 1677 291 1683
rect 445 1677 468 1683
rect 717 1677 740 1683
rect 1149 1677 1164 1683
rect 2564 1677 2579 1683
rect 2845 1677 2860 1683
rect 3420 1683 3428 1688
rect 3405 1677 3428 1683
rect 3549 1677 3564 1683
rect 4582 1616 4682 2004
rect 4242 1604 4682 1616
rect 3964 1532 3972 1536
rect 349 1517 371 1523
rect 477 1517 492 1523
rect 532 1517 547 1523
rect 557 1517 588 1523
rect 932 1517 947 1523
rect 1252 1517 1267 1523
rect 1533 1517 1571 1523
rect 1741 1517 1763 1523
rect 1981 1517 2003 1523
rect 2205 1517 2227 1523
rect 2301 1517 2316 1523
rect 2589 1517 2604 1523
rect 2637 1517 2652 1523
rect 3085 1517 3123 1523
rect 3252 1517 3267 1523
rect 3421 1517 3436 1523
rect 3476 1517 3491 1523
rect 1021 1497 1059 1503
rect 29 1477 51 1483
rect 196 1477 211 1483
rect 669 1477 684 1483
rect 964 1477 979 1483
rect 1053 1477 1059 1497
rect 2036 1497 2067 1503
rect 3293 1497 3308 1503
rect 1140 1477 1155 1483
rect 1172 1477 1187 1483
rect 68 1456 76 1464
rect 612 1456 620 1464
rect 740 1456 748 1464
rect 1181 1457 1187 1477
rect 1405 1477 1443 1483
rect 1805 1477 1827 1483
rect 2132 1477 2147 1483
rect 2596 1477 2611 1483
rect 2973 1477 3011 1483
rect 3037 1477 3059 1483
rect 3293 1477 3299 1497
rect 3709 1503 3715 1523
rect 4013 1517 4060 1523
rect 4205 1517 4220 1523
rect 3677 1497 3715 1503
rect 3741 1497 3779 1503
rect 3741 1477 3747 1497
rect 3869 1477 3907 1483
rect 1268 1456 1276 1464
rect 1524 1456 1532 1464
rect 1940 1457 1971 1463
rect 2164 1456 2172 1464
rect 2292 1457 2323 1463
rect 2628 1457 2659 1463
rect 2692 1456 2700 1464
rect 3156 1457 3187 1463
rect 3492 1456 3500 1464
rect 3821 1457 3852 1463
rect 3956 1456 3964 1464
rect 4084 1456 4092 1464
rect 340 1436 342 1444
rect 452 1436 454 1444
rect 650 1436 652 1444
rect 826 1436 828 1444
rect 1124 1436 1126 1444
rect 1732 1436 1734 1444
rect 1844 1436 1846 1444
rect 2372 1436 2374 1444
rect 2580 1436 2582 1444
rect 2788 1436 2790 1444
rect 2826 1436 2828 1444
rect 2884 1436 2886 1444
rect 3226 1436 3228 1444
rect 3412 1436 3414 1444
rect 3636 1436 3638 1444
rect 4164 1436 4166 1444
rect 4244 1436 4246 1444
rect -412 1404 8 1416
rect -412 1016 -312 1404
rect 186 1376 188 1384
rect 634 1376 636 1384
rect 986 1376 988 1384
rect 1786 1376 1788 1384
rect 1866 1376 1868 1384
rect 2410 1376 2412 1384
rect 2458 1376 2460 1384
rect 2506 1376 2508 1384
rect 3108 1376 3110 1384
rect 3732 1376 3734 1384
rect 3860 1376 3862 1384
rect 3988 1376 3990 1384
rect 228 1356 236 1364
rect 285 1357 316 1363
rect 804 1356 812 1364
rect 916 1357 947 1363
rect 1028 1356 1036 1364
rect 269 1337 300 1343
rect 333 1337 355 1343
rect 884 1337 899 1343
rect 1005 1337 1020 1343
rect 1213 1343 1219 1363
rect 1629 1357 1660 1363
rect 1917 1357 1948 1363
rect 2020 1356 2028 1364
rect 2308 1356 2316 1364
rect 3149 1357 3180 1363
rect 3453 1357 3484 1363
rect 3533 1357 3548 1363
rect 1133 1337 1155 1343
rect 1213 1337 1228 1343
rect 1245 1337 1267 1343
rect 1444 1337 1459 1343
rect 1492 1337 1507 1343
rect 1677 1323 1683 1343
rect 2077 1337 2099 1343
rect 2525 1337 2540 1343
rect 2884 1337 2899 1343
rect 3501 1337 3523 1343
rect 3565 1337 3580 1343
rect 3693 1337 3715 1343
rect 3837 1323 3843 1343
rect 1677 1317 1715 1323
rect 3805 1317 3843 1323
rect 157 1297 179 1303
rect 685 1297 723 1303
rect 1012 1297 1027 1303
rect 1636 1297 1651 1303
rect 2157 1297 2172 1303
rect 2708 1297 2723 1303
rect 3268 1297 3283 1303
rect 4045 1297 4067 1303
rect 4189 1297 4227 1303
rect 52 1277 67 1283
rect 413 1277 428 1283
rect 508 1283 516 1288
rect 493 1277 516 1283
rect 948 1277 963 1283
rect 1197 1277 1228 1283
rect 3044 1277 3059 1283
rect 3293 1277 3308 1283
rect 3437 1277 3452 1283
rect 3740 1283 3748 1288
rect 3740 1277 3779 1283
rect 4582 1216 4682 1604
rect 4242 1204 4682 1216
rect 109 1137 132 1143
rect 44 1132 52 1136
rect 124 1132 132 1137
rect 1012 1137 1027 1143
rect 1629 1137 1660 1143
rect 716 1132 724 1136
rect 1837 1117 1875 1123
rect 1940 1117 1955 1123
rect 1988 1117 2003 1123
rect 2180 1117 2195 1123
rect 2253 1117 2275 1123
rect 2996 1117 3011 1123
rect 3053 1117 3084 1123
rect 3229 1117 3251 1123
rect 3357 1117 3372 1123
rect 3693 1117 3708 1123
rect 4093 1117 4115 1123
rect 653 1097 691 1103
rect 157 1077 179 1083
rect 269 1077 284 1083
rect 324 1077 355 1083
rect 445 1077 483 1083
rect 685 1077 691 1097
rect 2989 1097 3004 1103
rect 804 1077 819 1083
rect 925 1077 947 1083
rect 1085 1077 1123 1083
rect 1357 1077 1379 1083
rect 1437 1077 1452 1083
rect 2333 1077 2348 1083
rect 1037 1057 1068 1063
rect 1236 1056 1244 1064
rect 1309 1057 1340 1063
rect 1389 1057 1420 1063
rect 1556 1057 1587 1063
rect 1876 1056 1884 1064
rect 2173 1057 2204 1063
rect 2333 1057 2339 1077
rect 2509 1077 2547 1083
rect 2836 1077 2851 1083
rect 2909 1077 2924 1083
rect 2484 1056 2492 1064
rect 2756 1057 2787 1063
rect 2909 1057 2915 1077
rect 2989 1077 2995 1097
rect 3629 1097 3667 1103
rect 3661 1084 3667 1097
rect 3597 1077 3612 1083
rect 4061 1077 4099 1083
rect 3012 1056 3020 1064
rect 3348 1057 3379 1063
rect 3844 1056 3852 1064
rect 4061 1057 4067 1077
rect 250 1036 252 1044
rect 426 1036 428 1044
rect 2442 1036 2444 1044
rect 3146 1036 3148 1044
rect 3578 1036 3580 1044
rect 4212 1036 4214 1044
rect -412 1004 12 1016
rect -412 616 -312 1004
rect 36 976 38 984
rect 410 976 412 984
rect 954 976 956 984
rect 1156 976 1158 984
rect 1252 976 1254 984
rect 1460 976 1462 984
rect 1764 976 1766 984
rect 1924 976 1926 984
rect 2116 976 2118 984
rect 2202 976 2204 984
rect 2954 976 2956 984
rect 3012 976 3014 984
rect 3082 976 3084 984
rect 3812 976 3814 984
rect 4042 976 4044 984
rect 4202 976 4204 984
rect 1284 956 1292 964
rect 2020 956 2028 964
rect 2500 957 2531 963
rect 2868 956 2876 964
rect 3268 957 3299 963
rect 317 937 339 943
rect 525 937 547 943
rect 701 917 739 923
rect 269 897 291 903
rect 733 897 739 917
rect 1005 917 1043 923
rect 1101 917 1116 923
rect 772 897 787 903
rect 1037 897 1043 917
rect 1229 923 1235 943
rect 1325 923 1331 943
rect 1837 937 1859 943
rect 1988 937 2003 943
rect 2157 937 2188 943
rect 2388 937 2403 943
rect 3101 937 3123 943
rect 3405 937 3443 943
rect 4013 937 4028 943
rect 1197 917 1235 923
rect 1293 917 1331 923
rect 1501 917 1516 923
rect 2237 917 2252 923
rect 2612 917 2643 923
rect 3364 917 3395 923
rect 3581 917 3596 923
rect 3613 917 3644 923
rect 3725 917 3763 923
rect 1117 897 1132 903
rect 1469 897 1484 903
rect 2509 897 2524 903
rect 2580 897 2595 903
rect 2781 897 2803 903
rect 3204 897 3219 903
rect 3309 897 3331 903
rect 3725 897 3731 917
rect 3901 897 3916 903
rect 3949 897 3971 903
rect 4173 897 4195 903
rect 204 883 212 888
rect 132 877 147 883
rect 173 877 212 883
rect 572 883 580 888
rect 2652 883 2660 888
rect 372 877 387 883
rect 572 877 611 883
rect 2652 877 2668 883
rect 2700 883 2708 888
rect 2700 877 2723 883
rect 2836 877 2851 883
rect 3068 883 3076 888
rect 3724 884 3732 888
rect 2916 877 2931 883
rect 3053 877 3076 883
rect 3437 877 3452 883
rect 4582 816 4682 1204
rect 4242 804 4682 816
rect 269 737 292 743
rect 284 732 292 737
rect 732 737 755 743
rect 732 732 740 737
rect 1532 737 1555 743
rect 1821 737 1852 743
rect 924 732 932 736
rect 1532 732 1540 737
rect 2173 737 2188 743
rect 2244 737 2259 743
rect 525 703 531 723
rect 564 717 579 723
rect 1037 717 1052 723
rect 1357 717 1372 723
rect 2045 717 2067 723
rect 2125 717 2140 723
rect 2676 717 2691 723
rect 3060 717 3075 723
rect 3613 717 3628 723
rect 493 697 531 703
rect 1021 697 1036 703
rect 3293 697 3331 703
rect 77 677 99 683
rect 317 677 339 683
rect 461 677 483 683
rect 557 677 595 683
rect 989 677 1011 683
rect 1197 677 1219 683
rect 1492 677 1507 683
rect 1844 677 1859 683
rect 2397 677 2435 683
rect 2797 677 2819 683
rect 3325 677 3331 697
rect 3597 677 3628 683
rect 3684 677 3699 683
rect 3965 677 4003 683
rect 4093 677 4108 683
rect 29 657 60 663
rect 372 656 380 664
rect 644 656 652 664
rect 1636 656 1644 664
rect 1709 657 1740 663
rect 1876 656 1884 664
rect 2068 656 2076 664
rect 2749 657 2780 663
rect 2980 657 3011 663
rect 3053 657 3084 663
rect 3748 656 3756 664
rect 4116 656 4124 664
rect 4180 657 4211 663
rect 180 636 182 644
rect 298 636 300 644
rect 724 636 726 644
rect 1130 636 1132 644
rect 1428 636 1430 644
rect 1476 636 1478 644
rect 1786 636 1788 644
rect 1924 636 1926 644
rect 2490 636 2492 644
rect 3812 636 3814 644
rect 3940 636 3942 644
rect -412 604 24 616
rect -412 216 -312 604
rect 570 576 572 584
rect 916 576 918 584
rect 1306 576 1308 584
rect 1882 576 1884 584
rect 2218 576 2220 584
rect 2378 576 2380 584
rect 3044 576 3046 584
rect 3082 576 3084 584
rect 3188 576 3190 584
rect 3604 576 3606 584
rect 4042 576 4044 584
rect 36 557 67 563
rect 221 557 252 563
rect 644 556 652 564
rect 724 556 732 564
rect 1156 557 1187 563
rect 1236 557 1267 563
rect 1437 557 1468 563
rect 1556 556 1564 564
rect 1693 557 1724 563
rect 1773 557 1804 563
rect 2029 557 2060 563
rect 2109 557 2140 563
rect 2461 557 2492 563
rect 2596 557 2627 563
rect 2996 556 3004 564
rect 3828 556 3836 564
rect 3860 556 3868 564
rect 4180 557 4211 563
rect 132 537 147 543
rect 468 537 483 543
rect 541 537 556 543
rect 877 537 899 543
rect 2397 537 2419 543
rect 2541 537 2579 543
rect 2676 537 2707 543
rect 2717 537 2739 543
rect 2925 537 2947 543
rect 4013 537 4028 543
rect 4068 537 4099 543
rect 4141 537 4163 543
rect 2829 517 2844 523
rect 3316 517 3347 523
rect 3908 517 3923 523
rect 228 497 243 503
rect 436 497 451 503
rect 500 497 515 503
rect 525 497 563 503
rect 925 497 940 503
rect 1101 497 1132 503
rect 1277 497 1299 503
rect 1444 497 1459 503
rect 1748 497 1763 503
rect 2301 497 2323 503
rect 3060 497 3075 503
rect 3197 497 3219 503
rect 3437 497 3459 503
rect 3693 497 3724 503
rect 3869 497 3907 503
rect 3972 497 3987 503
rect 4020 497 4035 503
rect 349 477 364 483
rect 676 477 691 483
rect 1053 477 1068 483
rect 1372 483 1380 488
rect 1372 477 1388 483
rect 2253 477 2284 483
rect 2364 483 2372 488
rect 2356 477 2372 483
rect 3517 477 3532 483
rect 4582 416 4682 804
rect 4242 404 4682 416
rect 1404 337 1427 343
rect 1404 332 1412 337
rect 1869 337 1892 343
rect 1804 332 1812 336
rect 1884 332 1892 337
rect 2092 332 2100 336
rect 2508 337 2531 343
rect 2508 332 2516 337
rect 2684 332 2692 336
rect 3757 337 3772 343
rect 3548 332 3556 336
rect 468 317 483 323
rect 717 317 739 323
rect 900 317 915 323
rect 1085 317 1107 323
rect 1213 317 1228 323
rect 2029 317 2051 323
rect 2685 317 2707 323
rect 2772 317 2787 323
rect 3300 317 3315 323
rect 4045 317 4067 323
rect 4205 317 4220 323
rect 2189 297 2204 303
rect 2589 297 2604 303
rect 340 277 355 283
rect 381 277 396 283
rect 260 256 268 264
rect 381 257 387 277
rect 461 277 499 283
rect 541 277 563 283
rect 637 277 675 283
rect 685 277 700 283
rect 893 277 931 283
rect 1565 277 1587 283
rect 1837 277 1852 283
rect 1949 277 1971 283
rect 2077 277 2092 283
rect 2125 277 2147 283
rect 2237 277 2259 283
rect 2317 277 2339 283
rect 2397 277 2419 283
rect 2461 277 2483 283
rect 2589 277 2595 297
rect 2925 277 2940 283
rect 3997 277 4019 283
rect 4157 277 4179 283
rect 740 256 748 264
rect 1268 256 1276 264
rect 1684 257 1715 263
rect 1988 257 2019 263
rect 2052 256 2060 264
rect 2269 257 2300 263
rect 2788 256 2796 264
rect 3156 256 3164 264
rect 3588 256 3596 264
rect 3956 257 3987 263
rect 74 236 76 244
rect 122 236 124 244
rect 826 236 828 244
rect 1146 236 1148 244
rect 1204 236 1206 244
rect 1626 236 1628 244
rect 1818 236 1820 244
rect 2378 236 2380 244
rect 2570 236 2572 244
rect 2628 236 2630 244
rect 2884 236 2886 244
rect 3108 236 3110 244
rect 3274 236 3276 244
rect 3322 236 3324 244
rect 3380 236 3382 244
rect 3428 236 3430 244
rect 3540 236 3542 244
rect 4196 236 4198 244
rect -412 204 26 216
rect -412 -2 -312 204
rect 218 176 220 184
rect 330 176 332 184
rect 410 176 412 184
rect 490 176 492 184
rect 682 176 684 184
rect 1338 176 1340 184
rect 1508 176 1510 184
rect 1578 176 1580 184
rect 1658 176 1660 184
rect 1940 176 1942 184
rect 2090 176 2092 184
rect 3204 176 3206 184
rect 3316 176 3318 184
rect 3396 176 3398 184
rect 3578 176 3580 184
rect 3882 176 3884 184
rect 4212 176 4214 184
rect 29 157 60 163
rect 980 157 1011 163
rect 2340 157 2371 163
rect 2532 156 2540 164
rect 2788 157 2819 163
rect 2852 156 2860 164
rect 2964 156 2972 164
rect 3508 156 3516 164
rect 77 137 92 143
rect 237 137 259 143
rect 349 137 371 143
rect 509 137 531 143
rect 589 137 611 143
rect 701 137 723 143
rect 797 123 803 143
rect 957 123 963 143
rect 1069 137 1091 143
rect 1396 137 1411 143
rect 548 117 579 123
rect 765 117 803 123
rect 925 117 963 123
rect 1229 117 1244 123
rect 109 97 124 103
rect 189 97 211 103
rect 461 97 483 103
rect 740 97 755 103
rect 829 97 851 103
rect 989 97 1004 103
rect 1021 97 1043 103
rect 1309 97 1331 103
rect 1437 103 1443 143
rect 1476 137 1491 143
rect 1677 137 1699 143
rect 1844 137 1859 143
rect 2173 137 2195 143
rect 2317 123 2323 143
rect 2381 137 2403 143
rect 2669 137 2691 143
rect 2877 137 2899 143
rect 2989 137 3004 143
rect 3277 137 3299 143
rect 3901 137 3923 143
rect 3965 137 3987 143
rect 4045 137 4067 143
rect 1956 117 1987 123
rect 2285 117 2323 123
rect 2564 117 2579 123
rect 2916 117 2931 123
rect 3437 117 3452 123
rect 4157 117 4188 123
rect 1428 97 1443 103
rect 2260 97 2275 103
rect 2429 97 2451 103
rect 2493 97 2531 103
rect 2605 97 2643 103
rect 2829 97 2851 103
rect 3021 97 3036 103
rect 3213 97 3235 103
rect 3517 97 3539 103
rect 3629 97 3651 103
rect 3860 97 3875 103
rect 316 83 324 88
rect 668 83 676 88
rect 285 77 324 83
rect 653 77 676 83
rect 1812 77 1827 83
rect 2076 83 2084 88
rect 2061 77 2084 83
rect 2141 77 2156 83
rect 2220 83 2228 88
rect 3324 83 3332 88
rect 3724 83 3732 88
rect 2220 77 2243 83
rect 3324 77 3347 83
rect 3724 77 3747 83
rect 4582 16 4682 404
rect 4242 4 4682 16
rect 4582 0 4682 4
<< m2contact >>
rect 220 2976 228 2984
rect 524 2976 532 2984
rect 588 2976 596 2984
rect 860 2976 868 2984
rect 1580 2976 1588 2984
rect 2524 2976 2532 2984
rect 2732 2976 2740 2984
rect 2860 2976 2868 2984
rect 2972 2976 2980 2984
rect 3388 2976 3396 2984
rect 3996 2976 4004 2984
rect 12 2956 20 2964
rect 140 2956 148 2964
rect 156 2956 164 2964
rect 236 2956 244 2964
rect 268 2956 276 2964
rect 428 2956 436 2964
rect 460 2956 468 2964
rect 540 2956 548 2964
rect 700 2956 708 2964
rect 732 2956 740 2964
rect 956 2956 964 2964
rect 972 2956 980 2964
rect 1100 2956 1108 2964
rect 1164 2956 1172 2964
rect 1372 2956 1380 2964
rect 1404 2956 1412 2964
rect 1436 2956 1444 2964
rect 1516 2956 1524 2964
rect 1596 2956 1604 2964
rect 1708 2956 1716 2964
rect 1740 2956 1748 2964
rect 1772 2956 1780 2964
rect 2012 2956 2020 2964
rect 2124 2956 2132 2964
rect 2156 2956 2164 2964
rect 2220 2956 2228 2964
rect 2252 2956 2260 2964
rect 2364 2956 2372 2964
rect 2396 2956 2404 2964
rect 2572 2956 2580 2964
rect 2668 2956 2676 2964
rect 380 2936 388 2944
rect 428 2936 436 2944
rect 492 2936 500 2944
rect 604 2936 612 2944
rect 764 2936 772 2944
rect 844 2936 852 2944
rect 876 2936 884 2944
rect 892 2936 900 2944
rect 1004 2936 1012 2944
rect 1020 2936 1028 2944
rect 1148 2936 1156 2944
rect 1500 2936 1508 2944
rect 1548 2936 1556 2944
rect 1676 2936 1684 2944
rect 1692 2936 1700 2944
rect 1756 2936 1764 2944
rect 1836 2936 1844 2944
rect 460 2916 468 2924
rect 764 2916 772 2924
rect 1996 2936 2004 2944
rect 2044 2936 2052 2944
rect 2060 2936 2068 2944
rect 2140 2936 2148 2944
rect 2252 2936 2260 2944
rect 2364 2936 2372 2944
rect 2428 2936 2436 2944
rect 2508 2936 2516 2944
rect 2556 2936 2564 2944
rect 2636 2936 2644 2944
rect 2764 2956 2772 2964
rect 2828 2956 2836 2964
rect 2892 2956 2900 2964
rect 2924 2956 2932 2964
rect 2988 2956 2996 2964
rect 3004 2956 3012 2964
rect 2764 2936 2772 2944
rect 2796 2936 2804 2944
rect 2844 2936 2852 2944
rect 2956 2936 2964 2944
rect 3164 2956 3172 2964
rect 3292 2956 3300 2964
rect 3532 2956 3540 2964
rect 3564 2956 3572 2964
rect 3580 2956 3588 2964
rect 3708 2956 3716 2964
rect 3836 2956 3844 2964
rect 3948 2956 3956 2964
rect 3964 2956 3972 2964
rect 4060 2956 4068 2964
rect 4140 2956 4148 2964
rect 4156 2956 4164 2964
rect 3068 2936 3076 2944
rect 3212 2936 3220 2944
rect 92 2896 100 2904
rect 124 2896 132 2904
rect 220 2896 228 2904
rect 252 2896 260 2904
rect 332 2896 340 2904
rect 412 2896 420 2904
rect 476 2896 484 2904
rect 524 2896 532 2904
rect 572 2896 580 2904
rect 652 2896 660 2904
rect 796 2896 804 2904
rect 844 2896 852 2904
rect 908 2896 916 2904
rect 972 2896 980 2904
rect 1052 2896 1060 2904
rect 1116 2896 1124 2904
rect 1228 2896 1236 2904
rect 1308 2896 1316 2904
rect 1420 2896 1428 2904
rect 1468 2896 1476 2904
rect 1580 2896 1588 2904
rect 1596 2896 1604 2904
rect 1628 2896 1636 2904
rect 1708 2896 1716 2904
rect 1804 2896 1812 2904
rect 1884 2896 1892 2904
rect 1964 2896 1972 2904
rect 2012 2896 2020 2904
rect 2092 2896 2100 2904
rect 2108 2896 2116 2904
rect 2300 2896 2308 2904
rect 2332 2916 2340 2924
rect 2396 2916 2404 2924
rect 3148 2916 3156 2924
rect 3244 2936 3252 2944
rect 3372 2936 3380 2944
rect 3276 2916 3284 2924
rect 3468 2936 3476 2944
rect 3628 2936 3636 2944
rect 3660 2936 3668 2944
rect 3676 2936 3684 2944
rect 4268 2936 4276 2944
rect 3532 2916 3540 2924
rect 3740 2916 3748 2924
rect 2396 2896 2404 2904
rect 2476 2896 2484 2904
rect 2524 2896 2532 2904
rect 2604 2896 2612 2904
rect 2700 2896 2708 2904
rect 2716 2896 2724 2904
rect 2748 2896 2756 2904
rect 2892 2896 2900 2904
rect 3116 2896 3124 2904
rect 3180 2896 3188 2904
rect 3260 2896 3268 2904
rect 3340 2896 3348 2904
rect 3420 2896 3428 2904
rect 3500 2896 3508 2904
rect 3644 2896 3652 2904
rect 3708 2896 3716 2904
rect 3836 2896 3844 2904
rect 3884 2896 3892 2904
rect 4076 2896 4084 2904
rect 92 2876 100 2884
rect 540 2876 548 2884
rect 684 2876 692 2884
rect 700 2876 708 2884
rect 1772 2876 1780 2884
rect 3052 2876 3060 2884
rect 3132 2876 3140 2884
rect 3324 2876 3332 2884
rect 3724 2876 3732 2884
rect 3756 2876 3764 2884
rect 1276 2856 1284 2864
rect 1532 2856 1540 2864
rect 1916 2856 1924 2864
rect 2444 2856 2452 2864
rect 364 2836 372 2844
rect 1260 2836 1268 2844
rect 1388 2836 1396 2844
rect 1932 2836 1940 2844
rect 2076 2836 2084 2844
rect 2652 2836 2660 2844
rect 2812 2836 2820 2844
rect 3020 2836 3028 2844
rect 3516 2836 3524 2844
rect 3820 2836 3828 2844
rect 4092 2836 4100 2844
rect 4204 2836 4212 2844
rect 652 2776 660 2784
rect 892 2776 900 2784
rect 1180 2776 1188 2784
rect 1308 2776 1316 2784
rect 1340 2776 1348 2784
rect 1788 2776 1796 2784
rect 2092 2776 2100 2784
rect 2220 2776 2228 2784
rect 2300 2776 2308 2784
rect 2716 2776 2724 2784
rect 2748 2776 2756 2784
rect 4060 2776 4068 2784
rect 4124 2776 4132 2784
rect 1452 2756 1460 2764
rect 2412 2756 2420 2764
rect 3836 2756 3844 2764
rect 4156 2756 4164 2764
rect 1020 2736 1028 2744
rect 1628 2736 1636 2744
rect 1708 2736 1716 2744
rect 2444 2736 2452 2744
rect 124 2716 132 2724
rect 156 2716 164 2724
rect 236 2716 244 2724
rect 284 2716 292 2724
rect 332 2716 340 2724
rect 412 2716 420 2724
rect 540 2716 548 2724
rect 588 2716 596 2724
rect 668 2716 676 2724
rect 716 2716 724 2724
rect 796 2716 804 2724
rect 876 2716 884 2724
rect 956 2716 964 2724
rect 1036 2716 1044 2724
rect 1100 2716 1108 2724
rect 1196 2716 1204 2724
rect 1292 2716 1300 2724
rect 1356 2716 1364 2724
rect 1404 2716 1412 2724
rect 1484 2716 1492 2724
rect 1532 2716 1540 2724
rect 1772 2716 1780 2724
rect 1932 2716 1940 2724
rect 2124 2716 2132 2724
rect 2172 2716 2180 2724
rect 2316 2716 2324 2724
rect 2476 2716 2484 2724
rect 2524 2716 2532 2724
rect 2636 2716 2644 2724
rect 2780 2716 2788 2724
rect 2876 2716 2884 2724
rect 3004 2716 3012 2724
rect 3132 2716 3140 2724
rect 3228 2716 3236 2724
rect 3324 2716 3332 2724
rect 3468 2716 3476 2724
rect 3548 2716 3556 2724
rect 3596 2716 3604 2724
rect 3660 2716 3668 2724
rect 3676 2716 3684 2724
rect 3724 2716 3732 2724
rect 3756 2716 3764 2724
rect 3772 2716 3780 2724
rect 3852 2716 3860 2724
rect 3900 2716 3908 2724
rect 3932 2716 3940 2724
rect 4044 2716 4052 2724
rect 4108 2716 4116 2724
rect 4188 2716 4196 2724
rect 12 2676 20 2684
rect 332 2676 340 2684
rect 380 2696 388 2704
rect 3068 2696 3076 2704
rect 380 2676 388 2684
rect 508 2676 516 2684
rect 620 2676 628 2684
rect 700 2676 708 2684
rect 748 2676 756 2684
rect 764 2676 772 2684
rect 828 2676 836 2684
rect 844 2676 852 2684
rect 924 2676 932 2684
rect 1148 2676 1156 2684
rect 1228 2676 1236 2684
rect 1244 2676 1252 2684
rect 1324 2676 1332 2684
rect 1436 2676 1444 2684
rect 1468 2676 1476 2684
rect 1516 2676 1524 2684
rect 1692 2676 1700 2684
rect 1724 2676 1732 2684
rect 2076 2676 2084 2684
rect 2108 2676 2116 2684
rect 2156 2676 2164 2684
rect 2204 2676 2212 2684
rect 2332 2676 2340 2684
rect 2508 2676 2516 2684
rect 2556 2676 2564 2684
rect 2812 2676 2820 2684
rect 2876 2676 2884 2684
rect 3052 2676 3060 2684
rect 3276 2676 3284 2684
rect 3500 2676 3508 2684
rect 3548 2676 3556 2684
rect 3628 2676 3636 2684
rect 3644 2676 3652 2684
rect 3692 2676 3700 2684
rect 3804 2676 3812 2684
rect 3884 2676 3892 2684
rect 3932 2676 3940 2684
rect 3980 2676 3988 2684
rect 4076 2676 4084 2684
rect 4220 2676 4228 2684
rect 76 2656 84 2664
rect 92 2656 100 2664
rect 172 2656 180 2664
rect 492 2656 500 2664
rect 524 2656 532 2664
rect 636 2656 644 2664
rect 876 2656 884 2664
rect 908 2656 916 2664
rect 972 2656 980 2664
rect 1004 2656 1012 2664
rect 1164 2656 1172 2664
rect 1292 2656 1300 2664
rect 1468 2656 1476 2664
rect 1548 2656 1556 2664
rect 1564 2656 1572 2664
rect 1660 2656 1668 2664
rect 1676 2656 1684 2664
rect 1724 2656 1732 2664
rect 1804 2656 1812 2664
rect 1820 2656 1828 2664
rect 1916 2656 1924 2664
rect 1996 2656 2004 2664
rect 2012 2656 2020 2664
rect 2108 2656 2116 2664
rect 2172 2656 2180 2664
rect 2236 2656 2244 2664
rect 2252 2656 2260 2664
rect 2348 2656 2356 2664
rect 2396 2656 2404 2664
rect 2428 2656 2436 2664
rect 2460 2656 2468 2664
rect 2540 2656 2548 2664
rect 2572 2656 2580 2664
rect 2620 2656 2628 2664
rect 2700 2656 2708 2664
rect 2732 2656 2740 2664
rect 2764 2656 2772 2664
rect 2828 2656 2836 2664
rect 2940 2656 2948 2664
rect 2956 2656 2964 2664
rect 3052 2656 3060 2664
rect 3132 2656 3140 2664
rect 3324 2656 3332 2664
rect 3356 2656 3364 2664
rect 3404 2656 3412 2664
rect 3724 2656 3732 2664
rect 3820 2656 3828 2664
rect 4108 2656 4116 2664
rect 4140 2656 4148 2664
rect 44 2636 52 2644
rect 156 2636 164 2644
rect 268 2636 276 2644
rect 300 2636 308 2644
rect 348 2636 356 2644
rect 412 2636 420 2644
rect 444 2636 452 2644
rect 556 2636 564 2644
rect 652 2636 660 2644
rect 684 2636 692 2644
rect 732 2636 740 2644
rect 956 2636 964 2644
rect 988 2636 996 2644
rect 1036 2636 1044 2644
rect 1196 2636 1204 2644
rect 1276 2636 1284 2644
rect 1772 2636 1780 2644
rect 1868 2636 1876 2644
rect 1948 2636 1956 2644
rect 2028 2636 2036 2644
rect 2044 2636 2052 2644
rect 2476 2636 2484 2644
rect 2636 2636 2644 2644
rect 2892 2636 2900 2644
rect 3164 2636 3172 2644
rect 3436 2636 3444 2644
rect 3548 2636 3556 2644
rect 3868 2636 3876 2644
rect 3900 2636 3908 2644
rect 76 2576 84 2584
rect 396 2576 404 2584
rect 524 2576 532 2584
rect 796 2576 804 2584
rect 1068 2576 1076 2584
rect 1148 2576 1156 2584
rect 1260 2576 1268 2584
rect 1388 2576 1396 2584
rect 1468 2576 1476 2584
rect 1740 2576 1748 2584
rect 1836 2576 1844 2584
rect 2012 2576 2020 2584
rect 2124 2576 2132 2584
rect 2156 2576 2164 2584
rect 2252 2576 2260 2584
rect 2780 2576 2788 2584
rect 2876 2576 2884 2584
rect 2924 2576 2932 2584
rect 2988 2576 2996 2584
rect 3100 2576 3108 2584
rect 3260 2576 3268 2584
rect 3500 2576 3508 2584
rect 3532 2576 3540 2584
rect 3692 2576 3700 2584
rect 3708 2576 3716 2584
rect 3804 2576 3812 2584
rect 3820 2576 3828 2584
rect 3884 2576 3892 2584
rect 3916 2576 3924 2584
rect 3980 2576 3988 2584
rect 4092 2576 4100 2584
rect 4156 2576 4164 2584
rect 4220 2576 4228 2584
rect 172 2556 180 2564
rect 252 2556 260 2564
rect 284 2556 292 2564
rect 412 2556 420 2564
rect 444 2556 452 2564
rect 476 2556 484 2564
rect 636 2556 644 2564
rect 668 2556 676 2564
rect 748 2556 756 2564
rect 780 2556 788 2564
rect 1244 2556 1252 2564
rect 1276 2556 1284 2564
rect 1292 2556 1300 2564
rect 1324 2556 1332 2564
rect 1420 2556 1428 2564
rect 1436 2556 1444 2564
rect 1692 2556 1700 2564
rect 1724 2556 1732 2564
rect 1868 2556 1876 2564
rect 1996 2556 2004 2564
rect 2444 2556 2452 2564
rect 2524 2556 2532 2564
rect 2556 2556 2564 2564
rect 2604 2556 2612 2564
rect 2620 2556 2628 2564
rect 2764 2556 2772 2564
rect 2940 2556 2948 2564
rect 3020 2556 3028 2564
rect 3052 2556 3060 2564
rect 3148 2556 3156 2564
rect 3388 2556 3396 2564
rect 3420 2556 3428 2564
rect 3548 2556 3556 2564
rect 3788 2556 3796 2564
rect 3868 2556 3876 2564
rect 3964 2556 3972 2564
rect 4044 2556 4052 2564
rect 4060 2556 4068 2564
rect 12 2536 20 2544
rect 348 2536 356 2544
rect 508 2536 516 2544
rect 540 2536 548 2544
rect 732 2536 740 2544
rect 812 2536 820 2544
rect 892 2536 900 2544
rect 988 2536 996 2544
rect 1020 2536 1028 2544
rect 940 2516 948 2524
rect 1116 2536 1124 2544
rect 1132 2536 1140 2544
rect 1356 2536 1364 2544
rect 1372 2536 1380 2544
rect 1484 2536 1492 2544
rect 1500 2536 1508 2544
rect 1548 2536 1556 2544
rect 1628 2536 1636 2544
rect 1676 2536 1684 2544
rect 1708 2536 1716 2544
rect 1788 2536 1796 2544
rect 1804 2536 1812 2544
rect 1900 2536 1908 2544
rect 1916 2536 1924 2544
rect 1932 2536 1940 2544
rect 2092 2536 2100 2544
rect 2108 2536 2116 2544
rect 2188 2536 2196 2544
rect 2204 2536 2212 2544
rect 2284 2536 2292 2544
rect 2332 2536 2340 2544
rect 2412 2536 2420 2544
rect 2444 2536 2452 2544
rect 2492 2536 2500 2544
rect 2540 2536 2548 2544
rect 2876 2536 2884 2544
rect 2908 2536 2916 2544
rect 2956 2536 2964 2544
rect 2988 2536 2996 2544
rect 3084 2536 3092 2544
rect 3164 2536 3172 2544
rect 3212 2536 3220 2544
rect 3292 2536 3300 2544
rect 3308 2536 3316 2544
rect 3340 2536 3348 2544
rect 3420 2536 3428 2544
rect 3468 2536 3476 2544
rect 3516 2536 3524 2544
rect 3564 2536 3572 2544
rect 3612 2536 3620 2544
rect 3644 2536 3652 2544
rect 3660 2536 3668 2544
rect 3772 2536 3780 2544
rect 3852 2536 3860 2544
rect 3900 2536 3908 2544
rect 4124 2536 4132 2544
rect 4172 2536 4180 2544
rect 4188 2536 4196 2544
rect 44 2496 52 2504
rect 124 2496 132 2504
rect 252 2496 260 2504
rect 364 2496 372 2504
rect 396 2496 404 2504
rect 492 2496 500 2504
rect 540 2496 548 2504
rect 588 2496 596 2504
rect 700 2496 708 2504
rect 844 2496 852 2504
rect 892 2496 900 2504
rect 940 2496 948 2504
rect 988 2496 996 2504
rect 1084 2496 1092 2504
rect 1964 2516 1972 2524
rect 1404 2496 1412 2504
rect 1452 2496 1460 2504
rect 1516 2496 1524 2504
rect 1532 2496 1540 2504
rect 1580 2496 1588 2504
rect 1660 2496 1668 2504
rect 1676 2496 1684 2504
rect 1756 2496 1764 2504
rect 1836 2496 1844 2504
rect 1868 2496 1876 2504
rect 1964 2496 1972 2504
rect 1996 2496 2004 2504
rect 2060 2496 2068 2504
rect 2140 2496 2148 2504
rect 2156 2496 2164 2504
rect 2236 2496 2244 2504
rect 2348 2516 2356 2524
rect 2300 2496 2308 2504
rect 2316 2496 2324 2504
rect 2364 2496 2372 2504
rect 2460 2496 2468 2504
rect 2684 2496 2692 2504
rect 2700 2496 2708 2504
rect 2764 2496 2772 2504
rect 2828 2496 2836 2504
rect 2876 2496 2884 2504
rect 2988 2496 2996 2504
rect 3036 2496 3044 2504
rect 3084 2496 3092 2504
rect 3196 2496 3204 2504
rect 3244 2496 3252 2504
rect 3340 2496 3348 2504
rect 3388 2496 3396 2504
rect 3436 2496 3444 2504
rect 3484 2496 3492 2504
rect 3612 2496 3620 2504
rect 3692 2496 3700 2504
rect 3724 2496 3732 2504
rect 3820 2496 3828 2504
rect 3980 2496 3988 2504
rect 4140 2496 4148 2504
rect 4220 2496 4228 2504
rect 1180 2476 1188 2484
rect 1804 2476 1812 2484
rect 2412 2476 2420 2484
rect 2492 2476 2500 2484
rect 2652 2476 2660 2484
rect 3420 2476 3428 2484
rect 3932 2476 3940 2484
rect 1612 2456 1620 2464
rect 2716 2456 2724 2464
rect 3324 2456 3332 2464
rect 156 2436 164 2444
rect 220 2436 228 2444
rect 268 2436 276 2444
rect 332 2436 340 2444
rect 428 2436 436 2444
rect 460 2436 468 2444
rect 620 2436 628 2444
rect 652 2436 660 2444
rect 668 2436 676 2444
rect 764 2436 772 2444
rect 1852 2436 1860 2444
rect 1980 2436 1988 2444
rect 3180 2436 3188 2444
rect 3948 2436 3956 2444
rect 940 2376 948 2384
rect 1148 2376 1156 2384
rect 1564 2376 1572 2384
rect 2012 2376 2020 2384
rect 2236 2376 2244 2384
rect 2764 2376 2772 2384
rect 2908 2376 2916 2384
rect 3244 2376 3252 2384
rect 3404 2376 3412 2384
rect 3612 2376 3620 2384
rect 3644 2376 3652 2384
rect 3980 2376 3988 2384
rect 3996 2376 4004 2384
rect 4044 2376 4052 2384
rect 1436 2356 1444 2364
rect 1612 2356 1620 2364
rect 1884 2356 1892 2364
rect 2892 2356 2900 2364
rect 1276 2336 1284 2344
rect 1324 2336 1332 2344
rect 2092 2336 2100 2344
rect 2412 2336 2420 2344
rect 3020 2336 3028 2344
rect 76 2316 84 2324
rect 156 2316 164 2324
rect 268 2316 276 2324
rect 316 2316 324 2324
rect 364 2316 372 2324
rect 380 2316 388 2324
rect 492 2316 500 2324
rect 508 2316 516 2324
rect 588 2316 596 2324
rect 620 2316 628 2324
rect 748 2316 756 2324
rect 780 2316 788 2324
rect 844 2316 852 2324
rect 876 2316 884 2324
rect 924 2316 932 2324
rect 956 2316 964 2324
rect 1004 2316 1012 2324
rect 1020 2316 1028 2324
rect 1052 2316 1060 2324
rect 1196 2316 1204 2324
rect 220 2296 228 2304
rect 380 2296 388 2304
rect 460 2296 468 2304
rect 700 2296 708 2304
rect 1292 2316 1300 2324
rect 1324 2316 1332 2324
rect 1420 2316 1428 2324
rect 1500 2316 1508 2324
rect 1548 2316 1556 2324
rect 1660 2316 1668 2324
rect 1724 2316 1732 2324
rect 1836 2316 1844 2324
rect 1980 2316 1988 2324
rect 1996 2316 2004 2324
rect 2044 2316 2052 2324
rect 2124 2316 2132 2324
rect 2140 2316 2148 2324
rect 2220 2316 2228 2324
rect 2268 2316 2276 2324
rect 2348 2316 2356 2324
rect 2044 2296 2052 2304
rect 2460 2316 2468 2324
rect 2540 2316 2548 2324
rect 2588 2316 2596 2324
rect 2604 2316 2612 2324
rect 2652 2316 2660 2324
rect 2700 2316 2708 2324
rect 2748 2316 2756 2324
rect 2780 2316 2788 2324
rect 2860 2316 2868 2324
rect 2940 2316 2948 2324
rect 2988 2316 2996 2324
rect 3084 2316 3092 2324
rect 3116 2316 3124 2324
rect 3180 2316 3188 2324
rect 3260 2316 3268 2324
rect 3356 2316 3364 2324
rect 3388 2316 3396 2324
rect 3436 2316 3444 2324
rect 3564 2316 3572 2324
rect 3596 2316 3604 2324
rect 3676 2316 3684 2324
rect 3804 2316 3812 2324
rect 3820 2316 3828 2324
rect 3868 2316 3876 2324
rect 3948 2316 3956 2324
rect 4060 2316 4068 2324
rect 4108 2316 4116 2324
rect 204 2276 212 2284
rect 236 2276 244 2284
rect 284 2276 292 2284
rect 332 2276 340 2284
rect 412 2276 420 2284
rect 460 2276 468 2284
rect 540 2276 548 2284
rect 588 2276 596 2284
rect 780 2276 788 2284
rect 828 2276 836 2284
rect 844 2276 852 2284
rect 988 2276 996 2284
rect 1036 2276 1044 2284
rect 1164 2276 1172 2284
rect 1244 2276 1252 2284
rect 1324 2276 1332 2284
rect 1372 2276 1380 2284
rect 1388 2276 1396 2284
rect 1580 2276 1588 2284
rect 1628 2276 1636 2284
rect 1676 2276 1684 2284
rect 1788 2276 1796 2284
rect 1804 2276 1812 2284
rect 1836 2276 1844 2284
rect 2028 2276 2036 2284
rect 2076 2276 2084 2284
rect 2092 2276 2100 2284
rect 2460 2296 2468 2304
rect 2188 2276 2196 2284
rect 2300 2276 2308 2284
rect 2316 2276 2324 2284
rect 2412 2276 2420 2284
rect 2556 2296 2564 2304
rect 2508 2276 2516 2284
rect 2556 2276 2564 2284
rect 3084 2296 3092 2304
rect 2652 2276 2660 2284
rect 2684 2276 2692 2284
rect 2812 2276 2820 2284
rect 2828 2276 2836 2284
rect 3020 2276 3028 2284
rect 3068 2276 3076 2284
rect 3116 2276 3124 2284
rect 3228 2296 3236 2304
rect 3868 2296 3876 2304
rect 3228 2276 3236 2284
rect 3308 2276 3316 2284
rect 3516 2276 3524 2284
rect 3564 2276 3572 2284
rect 3708 2276 3716 2284
rect 3724 2276 3732 2284
rect 3772 2276 3780 2284
rect 3852 2276 3860 2284
rect 3900 2276 3908 2284
rect 4092 2276 4100 2284
rect 4140 2276 4148 2284
rect 12 2256 20 2264
rect 92 2256 100 2264
rect 188 2256 196 2264
rect 204 2256 212 2264
rect 428 2256 436 2264
rect 492 2256 500 2264
rect 556 2256 564 2264
rect 636 2256 644 2264
rect 732 2256 740 2264
rect 924 2256 932 2264
rect 1116 2256 1124 2264
rect 1132 2256 1140 2264
rect 1260 2256 1268 2264
rect 1452 2256 1460 2264
rect 1468 2256 1476 2264
rect 1484 2256 1492 2264
rect 1596 2256 1604 2264
rect 1724 2256 1732 2264
rect 1836 2256 1844 2264
rect 1868 2256 1876 2264
rect 1900 2256 1908 2264
rect 1916 2256 1924 2264
rect 2140 2256 2148 2264
rect 2748 2256 2756 2264
rect 2780 2256 2788 2264
rect 3276 2256 3284 2264
rect 3500 2256 3508 2264
rect 3628 2256 3636 2264
rect 3948 2256 3956 2264
rect 3964 2256 3972 2264
rect 4012 2256 4020 2264
rect 4028 2256 4036 2264
rect 4156 2256 4164 2264
rect 4188 2256 4196 2264
rect 4252 2256 4260 2264
rect 60 2236 68 2244
rect 140 2236 148 2244
rect 252 2236 260 2244
rect 316 2236 324 2244
rect 380 2236 388 2244
rect 508 2236 516 2244
rect 604 2236 612 2244
rect 764 2236 772 2244
rect 956 2236 964 2244
rect 1052 2236 1060 2244
rect 1212 2236 1220 2244
rect 1308 2236 1316 2244
rect 1356 2236 1364 2244
rect 1420 2236 1428 2244
rect 1516 2236 1524 2244
rect 1644 2236 1652 2244
rect 1708 2236 1716 2244
rect 1756 2236 1764 2244
rect 1964 2236 1972 2244
rect 2124 2236 2132 2244
rect 2236 2236 2244 2244
rect 2396 2236 2404 2244
rect 2444 2236 2452 2244
rect 2476 2236 2484 2244
rect 2588 2236 2596 2244
rect 2620 2236 2628 2244
rect 2684 2236 2692 2244
rect 2732 2236 2740 2244
rect 3084 2236 3092 2244
rect 3148 2236 3156 2244
rect 3292 2236 3300 2244
rect 3372 2236 3380 2244
rect 3548 2236 3556 2244
rect 3580 2236 3588 2244
rect 3756 2236 3764 2244
rect 4076 2236 4084 2244
rect 4124 2236 4132 2244
rect 156 2176 164 2184
rect 668 2176 676 2184
rect 844 2176 852 2184
rect 924 2176 932 2184
rect 988 2176 996 2184
rect 1084 2176 1092 2184
rect 1116 2176 1124 2184
rect 1228 2176 1236 2184
rect 1276 2176 1284 2184
rect 1308 2176 1316 2184
rect 1356 2176 1364 2184
rect 1436 2176 1444 2184
rect 1564 2176 1572 2184
rect 1676 2176 1684 2184
rect 1756 2176 1764 2184
rect 1852 2176 1860 2184
rect 1932 2176 1940 2184
rect 2364 2176 2372 2184
rect 2604 2176 2612 2184
rect 2844 2176 2852 2184
rect 3100 2176 3108 2184
rect 3468 2176 3476 2184
rect 3628 2176 3636 2184
rect 4028 2176 4036 2184
rect 28 2156 36 2164
rect 60 2156 68 2164
rect 108 2156 116 2164
rect 124 2156 132 2164
rect 172 2156 180 2164
rect 204 2156 212 2164
rect 220 2156 228 2164
rect 252 2156 260 2164
rect 348 2156 356 2164
rect 380 2156 388 2164
rect 444 2156 452 2164
rect 540 2156 548 2164
rect 748 2156 756 2164
rect 892 2156 900 2164
rect 956 2156 964 2164
rect 1372 2156 1380 2164
rect 1404 2156 1412 2164
rect 1612 2156 1620 2164
rect 1644 2156 1652 2164
rect 1708 2156 1716 2164
rect 1836 2156 1844 2164
rect 1900 2156 1908 2164
rect 1916 2156 1924 2164
rect 2156 2156 2164 2164
rect 2236 2156 2244 2164
rect 2268 2156 2276 2164
rect 2396 2156 2404 2164
rect 2444 2156 2452 2164
rect 2476 2156 2484 2164
rect 2508 2156 2516 2164
rect 2540 2156 2548 2164
rect 2556 2156 2564 2164
rect 2620 2156 2628 2164
rect 2732 2156 2740 2164
rect 2908 2156 2916 2164
rect 2940 2156 2948 2164
rect 3036 2156 3044 2164
rect 3052 2156 3060 2164
rect 3148 2156 3156 2164
rect 3308 2156 3316 2164
rect 60 2136 68 2144
rect 92 2136 100 2144
rect 316 2136 324 2144
rect 428 2136 436 2144
rect 524 2136 532 2144
rect 652 2136 660 2144
rect 732 2136 740 2144
rect 780 2136 788 2144
rect 828 2136 836 2144
rect 940 2136 948 2144
rect 1052 2136 1060 2144
rect 1068 2136 1076 2144
rect 1164 2136 1172 2144
rect 1180 2136 1188 2144
rect 1196 2136 1204 2144
rect 1212 2136 1220 2144
rect 1292 2136 1300 2144
rect 1340 2136 1348 2144
rect 1388 2136 1396 2144
rect 1420 2136 1428 2144
rect 1468 2136 1476 2144
rect 1580 2136 1588 2144
rect 1660 2136 1668 2144
rect 1740 2136 1748 2144
rect 1788 2136 1796 2144
rect 1804 2136 1812 2144
rect 1884 2136 1892 2144
rect 1964 2136 1972 2144
rect 1980 2136 1988 2144
rect 2028 2136 2036 2144
rect 2332 2136 2340 2144
rect 2380 2136 2388 2144
rect 2492 2136 2500 2144
rect 2572 2136 2580 2144
rect 2732 2136 2740 2144
rect 2764 2136 2772 2144
rect 2892 2136 2900 2144
rect 3116 2136 3124 2144
rect 3164 2136 3172 2144
rect 3260 2136 3268 2144
rect 3308 2136 3316 2144
rect 3436 2156 3444 2164
rect 3564 2156 3572 2164
rect 3692 2156 3700 2164
rect 3756 2156 3764 2164
rect 3772 2156 3780 2164
rect 3916 2156 3924 2164
rect 3932 2156 3940 2164
rect 4140 2156 4148 2164
rect 3356 2136 3364 2144
rect 3596 2136 3604 2144
rect 3612 2136 3620 2144
rect 3660 2136 3668 2144
rect 3708 2136 3716 2144
rect 3724 2136 3732 2144
rect 3804 2136 3812 2144
rect 3884 2136 3892 2144
rect 3964 2136 3972 2144
rect 4060 2136 4068 2144
rect 284 2116 292 2124
rect 348 2116 356 2124
rect 828 2116 836 2124
rect 1580 2116 1588 2124
rect 2140 2116 2148 2124
rect 2764 2116 2772 2124
rect 3804 2116 3812 2124
rect 4092 2136 4100 2144
rect 4172 2136 4180 2144
rect 12 2096 20 2104
rect 284 2096 292 2104
rect 316 2096 324 2104
rect 396 2096 404 2104
rect 476 2096 484 2104
rect 556 2096 564 2104
rect 572 2096 580 2104
rect 620 2096 628 2104
rect 684 2096 692 2104
rect 812 2096 820 2104
rect 860 2096 868 2104
rect 908 2096 916 2104
rect 1020 2096 1028 2104
rect 1116 2096 1124 2104
rect 1164 2096 1172 2104
rect 1244 2096 1252 2104
rect 1260 2096 1268 2104
rect 1308 2096 1316 2104
rect 1468 2096 1476 2104
rect 1500 2096 1508 2104
rect 1692 2096 1700 2104
rect 1708 2096 1716 2104
rect 1836 2096 1844 2104
rect 1852 2096 1860 2104
rect 1932 2096 1940 2104
rect 2012 2096 2020 2104
rect 2060 2096 2068 2104
rect 2108 2096 2116 2104
rect 2332 2096 2340 2104
rect 2524 2096 2532 2104
rect 2604 2096 2612 2104
rect 2684 2096 2692 2104
rect 2796 2096 2804 2104
rect 2844 2096 2852 2104
rect 2860 2096 2868 2104
rect 2908 2096 2916 2104
rect 2972 2096 2980 2104
rect 3084 2096 3092 2104
rect 3196 2096 3204 2104
rect 3388 2096 3396 2104
rect 3500 2096 3508 2104
rect 3580 2096 3588 2104
rect 3628 2096 3636 2104
rect 3676 2096 3684 2104
rect 3756 2096 3764 2104
rect 3836 2096 3844 2104
rect 3916 2096 3924 2104
rect 3964 2096 3972 2104
rect 3996 2096 4004 2104
rect 4044 2096 4052 2104
rect 4124 2096 4132 2104
rect 4172 2096 4180 2104
rect 4204 2096 4212 2104
rect 252 2076 260 2084
rect 1100 2076 1108 2084
rect 1756 2076 1764 2084
rect 2236 2076 2244 2084
rect 2908 2076 2916 2084
rect 3052 2076 3060 2084
rect 3852 2076 3860 2084
rect 588 2056 596 2064
rect 764 2056 772 2064
rect 1996 2056 2004 2064
rect 76 2036 84 2044
rect 140 2036 148 2044
rect 188 2036 196 2044
rect 236 2036 244 2044
rect 876 2036 884 2044
rect 972 2036 980 2044
rect 1532 2036 1540 2044
rect 1628 2036 1636 2044
rect 2316 2036 2324 2044
rect 2412 2036 2420 2044
rect 2428 2036 2436 2044
rect 2460 2036 2468 2044
rect 2636 2036 2644 2044
rect 2652 2036 2660 2044
rect 2748 2036 2756 2044
rect 3340 2036 3348 2044
rect 3420 2036 3428 2044
rect 3452 2036 3460 2044
rect 4028 2036 4036 2044
rect 4252 2036 4260 2044
rect 348 1976 356 1984
rect 732 1976 740 1984
rect 780 1976 788 1984
rect 1100 1976 1108 1984
rect 1356 1976 1364 1984
rect 1468 1976 1476 1984
rect 1772 1976 1780 1984
rect 1804 1976 1812 1984
rect 1852 1976 1860 1984
rect 2076 1976 2084 1984
rect 2668 1976 2676 1984
rect 3068 1976 3076 1984
rect 3100 1976 3108 1984
rect 3356 1976 3364 1984
rect 3836 1976 3844 1984
rect 316 1956 324 1964
rect 1740 1956 1748 1964
rect 2124 1956 2132 1964
rect 2156 1956 2164 1964
rect 3596 1956 3604 1964
rect 908 1936 916 1944
rect 1484 1936 1492 1944
rect 1564 1936 1572 1944
rect 2012 1936 2020 1944
rect 44 1916 52 1924
rect 92 1916 100 1924
rect 172 1916 180 1924
rect 268 1916 276 1924
rect 460 1916 468 1924
rect 540 1916 548 1924
rect 636 1916 644 1924
rect 668 1916 676 1924
rect 716 1916 724 1924
rect 796 1916 804 1924
rect 876 1916 884 1924
rect 972 1916 980 1924
rect 1084 1916 1092 1924
rect 1132 1916 1140 1924
rect 1164 1916 1172 1924
rect 1308 1916 1316 1924
rect 1532 1916 1540 1924
rect 1612 1916 1620 1924
rect 1724 1916 1732 1924
rect 1868 1916 1876 1924
rect 1884 1916 1892 1924
rect 1980 1916 1988 1924
rect 2108 1916 2116 1924
rect 2204 1916 2212 1924
rect 2252 1916 2260 1924
rect 2300 1916 2308 1924
rect 2348 1916 2356 1924
rect 2396 1916 2404 1924
rect 2412 1916 2420 1924
rect 2476 1916 2484 1924
rect 2524 1916 2532 1924
rect 124 1896 132 1904
rect 12 1876 20 1884
rect 44 1876 52 1884
rect 124 1876 132 1884
rect 252 1876 260 1884
rect 300 1876 308 1884
rect 380 1876 388 1884
rect 892 1896 900 1904
rect 2588 1916 2596 1924
rect 2844 1916 2852 1924
rect 2908 1916 2916 1924
rect 3020 1916 3028 1924
rect 3180 1916 3188 1924
rect 3228 1916 3236 1924
rect 3292 1916 3300 1924
rect 3308 1916 3316 1924
rect 3468 1916 3476 1924
rect 3500 1916 3508 1924
rect 3532 1916 3540 1924
rect 3548 1916 3556 1924
rect 3708 1916 3716 1924
rect 3820 1916 3828 1924
rect 3868 1916 3876 1924
rect 3948 1916 3956 1924
rect 3996 1916 4004 1924
rect 4076 1916 4084 1924
rect 2812 1896 2820 1904
rect 3260 1896 3268 1904
rect 508 1876 516 1884
rect 636 1876 644 1884
rect 828 1876 836 1884
rect 844 1876 852 1884
rect 940 1876 948 1884
rect 956 1876 964 1884
rect 1004 1876 1012 1884
rect 1036 1876 1044 1884
rect 1052 1876 1060 1884
rect 1180 1876 1188 1884
rect 1212 1876 1220 1884
rect 1228 1876 1236 1884
rect 1340 1876 1348 1884
rect 1388 1876 1396 1884
rect 1564 1876 1572 1884
rect 1644 1876 1652 1884
rect 1660 1876 1668 1884
rect 1692 1876 1700 1884
rect 1836 1876 1844 1884
rect 1916 1876 1924 1884
rect 2012 1876 2020 1884
rect 2044 1876 2052 1884
rect 2172 1876 2180 1884
rect 2220 1876 2228 1884
rect 2268 1876 2276 1884
rect 2316 1876 2324 1884
rect 2348 1876 2356 1884
rect 2444 1876 2452 1884
rect 2492 1876 2500 1884
rect 2588 1876 2596 1884
rect 2620 1876 2628 1884
rect 2652 1876 2660 1884
rect 2684 1876 2692 1884
rect 2812 1876 2820 1884
rect 2892 1876 2900 1884
rect 2940 1876 2948 1884
rect 3004 1876 3012 1884
rect 3052 1876 3060 1884
rect 3116 1876 3124 1884
rect 3180 1876 3188 1884
rect 3260 1876 3268 1884
rect 3340 1876 3348 1884
rect 3404 1876 3412 1884
rect 3500 1876 3508 1884
rect 3516 1876 3524 1884
rect 3580 1876 3588 1884
rect 3740 1876 3748 1884
rect 3916 1876 3924 1884
rect 4108 1876 4116 1884
rect 4156 1876 4164 1884
rect 4220 1876 4228 1884
rect 28 1856 36 1864
rect 188 1856 196 1864
rect 332 1856 340 1864
rect 364 1856 372 1864
rect 444 1856 452 1864
rect 556 1856 564 1864
rect 748 1856 756 1864
rect 764 1856 772 1864
rect 892 1856 900 1864
rect 1020 1856 1028 1864
rect 1116 1856 1124 1864
rect 1292 1856 1300 1864
rect 1372 1856 1380 1864
rect 1452 1856 1460 1864
rect 1484 1856 1492 1864
rect 1596 1856 1604 1864
rect 1676 1856 1684 1864
rect 1756 1856 1764 1864
rect 1788 1856 1796 1864
rect 1820 1856 1828 1864
rect 1932 1856 1940 1864
rect 2044 1856 2052 1864
rect 2108 1856 2116 1864
rect 2140 1856 2148 1864
rect 2348 1856 2356 1864
rect 2428 1856 2436 1864
rect 2460 1856 2468 1864
rect 2636 1856 2644 1864
rect 2684 1856 2692 1864
rect 2764 1856 2772 1864
rect 2780 1856 2788 1864
rect 2924 1856 2932 1864
rect 2956 1856 2964 1864
rect 3036 1856 3044 1864
rect 3084 1856 3092 1864
rect 3116 1856 3124 1864
rect 3292 1856 3300 1864
rect 3372 1856 3380 1864
rect 3404 1856 3412 1864
rect 3612 1856 3620 1864
rect 3644 1856 3652 1864
rect 3772 1856 3780 1864
rect 3980 1856 3988 1864
rect 4044 1856 4052 1864
rect 4076 1856 4084 1864
rect 4124 1856 4132 1864
rect 4156 1856 4164 1864
rect 156 1836 164 1844
rect 236 1836 244 1844
rect 284 1836 292 1844
rect 412 1836 420 1844
rect 476 1836 484 1844
rect 604 1836 612 1844
rect 652 1836 660 1844
rect 716 1836 724 1844
rect 796 1836 804 1844
rect 860 1836 868 1844
rect 972 1836 980 1844
rect 1068 1836 1076 1844
rect 1148 1836 1156 1844
rect 1180 1836 1188 1844
rect 1244 1836 1252 1844
rect 1324 1836 1332 1844
rect 1404 1836 1412 1844
rect 1500 1836 1508 1844
rect 1612 1836 1620 1844
rect 1724 1836 1732 1844
rect 1868 1836 1876 1844
rect 1996 1836 2004 1844
rect 2188 1836 2196 1844
rect 2252 1836 2260 1844
rect 2300 1836 2308 1844
rect 2380 1836 2388 1844
rect 2732 1836 2740 1844
rect 2828 1836 2836 1844
rect 2876 1836 2884 1844
rect 3148 1836 3156 1844
rect 3324 1836 3332 1844
rect 3388 1836 3396 1844
rect 3548 1836 3556 1844
rect 3660 1836 3668 1844
rect 3820 1836 3828 1844
rect 3836 1836 3844 1844
rect 4012 1836 4020 1844
rect 4204 1836 4212 1844
rect 12 1776 20 1784
rect 188 1776 196 1784
rect 460 1776 468 1784
rect 556 1776 564 1784
rect 892 1776 900 1784
rect 940 1776 948 1784
rect 1004 1776 1012 1784
rect 1212 1776 1220 1784
rect 1356 1776 1364 1784
rect 1420 1776 1428 1784
rect 1740 1776 1748 1784
rect 1916 1776 1924 1784
rect 2108 1776 2116 1784
rect 2396 1776 2404 1784
rect 2444 1776 2452 1784
rect 2684 1776 2692 1784
rect 2780 1776 2788 1784
rect 2940 1776 2948 1784
rect 3052 1776 3060 1784
rect 3100 1776 3108 1784
rect 3212 1776 3220 1784
rect 3308 1776 3316 1784
rect 3420 1776 3428 1784
rect 3612 1776 3620 1784
rect 3708 1776 3716 1784
rect 3788 1776 3796 1784
rect 3932 1776 3940 1784
rect 140 1756 148 1764
rect 236 1756 244 1764
rect 268 1756 276 1764
rect 300 1756 308 1764
rect 316 1756 324 1764
rect 332 1756 340 1764
rect 348 1756 356 1764
rect 412 1756 420 1764
rect 428 1756 436 1764
rect 508 1756 516 1764
rect 588 1756 596 1764
rect 700 1756 708 1764
rect 796 1756 804 1764
rect 828 1756 836 1764
rect 860 1756 868 1764
rect 956 1756 964 1764
rect 1084 1756 1092 1764
rect 1100 1756 1108 1764
rect 1164 1756 1172 1764
rect 1180 1756 1188 1764
rect 1276 1756 1284 1764
rect 1292 1756 1300 1764
rect 1340 1756 1348 1764
rect 1372 1756 1380 1764
rect 1628 1756 1636 1764
rect 1852 1756 1860 1764
rect 1884 1756 1892 1764
rect 1948 1756 1956 1764
rect 2316 1756 2324 1764
rect 2348 1756 2356 1764
rect 2428 1756 2436 1764
rect 2460 1756 2468 1764
rect 2524 1756 2532 1764
rect 2556 1756 2564 1764
rect 2716 1756 2724 1764
rect 2796 1756 2804 1764
rect 2860 1756 2868 1764
rect 3020 1756 3028 1764
rect 3068 1756 3076 1764
rect 3132 1756 3140 1764
rect 3324 1756 3332 1764
rect 3388 1756 3396 1764
rect 3484 1756 3492 1764
rect 3500 1756 3508 1764
rect 3580 1756 3588 1764
rect 3628 1756 3636 1764
rect 3644 1756 3652 1764
rect 3676 1756 3684 1764
rect 3772 1756 3780 1764
rect 3884 1756 3892 1764
rect 3980 1756 3988 1764
rect 4012 1756 4020 1764
rect 4044 1756 4052 1764
rect 4124 1756 4132 1764
rect 4172 1756 4180 1764
rect 124 1736 132 1744
rect 204 1736 212 1744
rect 236 1736 244 1744
rect 492 1736 500 1744
rect 588 1736 596 1744
rect 844 1736 852 1744
rect 924 1736 932 1744
rect 972 1736 980 1744
rect 1132 1736 1140 1744
rect 1324 1736 1332 1744
rect 1404 1736 1412 1744
rect 1484 1736 1492 1744
rect 1500 1736 1508 1744
rect 1580 1736 1588 1744
rect 1596 1736 1604 1744
rect 1724 1736 1732 1744
rect 1820 1736 1828 1744
rect 1852 1736 1860 1744
rect 1900 1736 1908 1744
rect 2060 1736 2068 1744
rect 2076 1736 2084 1744
rect 2124 1736 2132 1744
rect 2204 1736 2212 1744
rect 2220 1736 2228 1744
rect 2348 1736 2356 1744
rect 2412 1736 2420 1744
rect 2492 1736 2500 1744
rect 2540 1736 2548 1744
rect 2588 1736 2596 1744
rect 2748 1736 2756 1744
rect 2828 1736 2836 1744
rect 2860 1736 2868 1744
rect 2908 1736 2916 1744
rect 2924 1736 2932 1744
rect 2972 1736 2980 1744
rect 3068 1736 3076 1744
rect 3164 1736 3172 1744
rect 3244 1736 3252 1744
rect 3260 1736 3268 1744
rect 3340 1736 3348 1744
rect 3532 1736 3540 1744
rect 3564 1736 3572 1744
rect 3820 1736 3828 1744
rect 3836 1736 3844 1744
rect 3980 1736 3988 1744
rect 4028 1736 4036 1744
rect 4108 1736 4116 1744
rect 4252 1736 4260 1744
rect 12 1696 20 1704
rect 92 1696 100 1704
rect 348 1696 356 1704
rect 668 1696 676 1704
rect 812 1696 820 1704
rect 1660 1716 1668 1724
rect 2156 1716 2164 1724
rect 1020 1696 1028 1704
rect 1100 1696 1108 1704
rect 1212 1696 1220 1704
rect 1292 1696 1300 1704
rect 1372 1696 1380 1704
rect 1452 1696 1460 1704
rect 1532 1696 1540 1704
rect 1612 1696 1620 1704
rect 1692 1696 1700 1704
rect 1740 1696 1748 1704
rect 1788 1696 1796 1704
rect 1932 1696 1940 1704
rect 1948 1696 1956 1704
rect 2028 1696 2036 1704
rect 2108 1696 2116 1704
rect 2156 1696 2164 1704
rect 2172 1696 2180 1704
rect 2252 1696 2260 1704
rect 2300 1696 2308 1704
rect 2380 1696 2388 1704
rect 2460 1696 2468 1704
rect 2620 1696 2628 1704
rect 2716 1696 2724 1704
rect 2780 1696 2788 1704
rect 2796 1696 2804 1704
rect 2876 1696 2884 1704
rect 2956 1696 2964 1704
rect 3004 1696 3012 1704
rect 3036 1696 3044 1704
rect 3116 1696 3124 1704
rect 3196 1696 3204 1704
rect 3276 1716 3284 1724
rect 3852 1716 3860 1724
rect 3292 1696 3300 1704
rect 3372 1696 3380 1704
rect 3532 1696 3540 1704
rect 3676 1696 3684 1704
rect 3708 1696 3716 1704
rect 3788 1696 3796 1704
rect 3868 1696 3876 1704
rect 4060 1696 4068 1704
rect 4076 1696 4084 1704
rect 4220 1696 4228 1704
rect 268 1676 276 1684
rect 1164 1676 1172 1684
rect 2556 1676 2564 1684
rect 2860 1676 2868 1684
rect 3564 1676 3572 1684
rect 2284 1656 2292 1664
rect 3356 1656 3364 1664
rect 220 1636 228 1644
rect 684 1636 692 1644
rect 748 1636 756 1644
rect 1196 1636 1204 1644
rect 1564 1636 1572 1644
rect 1644 1636 1652 1644
rect 1836 1636 1844 1644
rect 2140 1636 2148 1644
rect 2364 1636 2372 1644
rect 2988 1636 2996 1644
rect 3148 1636 3156 1644
rect 3596 1636 3604 1644
rect 3692 1636 3700 1644
rect 4092 1636 4100 1644
rect 4140 1636 4148 1644
rect 4156 1636 4164 1644
rect 4188 1636 4196 1644
rect 92 1576 100 1584
rect 172 1576 180 1584
rect 396 1576 404 1584
rect 780 1576 788 1584
rect 1324 1576 1332 1584
rect 1484 1576 1492 1584
rect 1884 1576 1892 1584
rect 2204 1576 2212 1584
rect 2524 1576 2532 1584
rect 2668 1576 2676 1584
rect 2732 1576 2740 1584
rect 2924 1576 2932 1584
rect 3196 1576 3204 1584
rect 3356 1576 3364 1584
rect 3804 1576 3812 1584
rect 4124 1576 4132 1584
rect 236 1556 244 1564
rect 508 1556 516 1564
rect 860 1556 868 1564
rect 1340 1556 1348 1564
rect 3068 1556 3076 1564
rect 3596 1556 3604 1564
rect 3964 1536 3972 1544
rect 76 1516 84 1524
rect 124 1516 132 1524
rect 268 1516 276 1524
rect 460 1516 468 1524
rect 492 1516 500 1524
rect 524 1516 532 1524
rect 588 1516 596 1524
rect 620 1516 628 1524
rect 636 1516 644 1524
rect 684 1516 692 1524
rect 732 1516 740 1524
rect 812 1516 820 1524
rect 892 1516 900 1524
rect 924 1516 932 1524
rect 1004 1516 1012 1524
rect 1084 1516 1092 1524
rect 1132 1516 1140 1524
rect 1196 1516 1204 1524
rect 1212 1516 1220 1524
rect 1244 1516 1252 1524
rect 1372 1516 1380 1524
rect 1420 1516 1428 1524
rect 1612 1516 1620 1524
rect 1660 1516 1668 1524
rect 1852 1516 1860 1524
rect 1868 1516 1876 1524
rect 1948 1516 1956 1524
rect 2044 1516 2052 1524
rect 2092 1516 2100 1524
rect 2172 1516 2180 1524
rect 2316 1516 2324 1524
rect 2332 1516 2340 1524
rect 2380 1516 2388 1524
rect 2396 1516 2404 1524
rect 2476 1516 2484 1524
rect 2604 1516 2612 1524
rect 2652 1516 2660 1524
rect 2684 1516 2692 1524
rect 2796 1516 2804 1524
rect 2812 1516 2820 1524
rect 2892 1516 2900 1524
rect 2940 1516 2948 1524
rect 3164 1516 3172 1524
rect 3212 1516 3220 1524
rect 3244 1516 3252 1524
rect 3340 1516 3348 1524
rect 3436 1516 3444 1524
rect 3468 1516 3476 1524
rect 3532 1516 3540 1524
rect 3644 1516 3652 1524
rect 3692 1516 3700 1524
rect 156 1476 164 1484
rect 188 1476 196 1484
rect 300 1476 308 1484
rect 316 1476 324 1484
rect 428 1476 436 1484
rect 572 1476 580 1484
rect 588 1476 596 1484
rect 684 1476 692 1484
rect 716 1476 724 1484
rect 764 1476 772 1484
rect 844 1476 852 1484
rect 924 1476 932 1484
rect 956 1476 964 1484
rect 1036 1476 1044 1484
rect 2028 1496 2036 1504
rect 2956 1496 2964 1504
rect 1100 1476 1108 1484
rect 1132 1476 1140 1484
rect 1164 1476 1172 1484
rect 12 1456 20 1464
rect 76 1456 84 1464
rect 108 1456 116 1464
rect 188 1456 196 1464
rect 220 1456 228 1464
rect 252 1456 260 1464
rect 380 1456 388 1464
rect 412 1456 420 1464
rect 492 1456 500 1464
rect 524 1456 532 1464
rect 620 1456 628 1464
rect 732 1456 740 1464
rect 796 1456 804 1464
rect 876 1456 884 1464
rect 956 1456 964 1464
rect 988 1456 996 1464
rect 1164 1456 1172 1464
rect 1244 1476 1252 1484
rect 1292 1476 1300 1484
rect 1452 1476 1460 1484
rect 1500 1476 1508 1484
rect 1580 1476 1588 1484
rect 1692 1476 1700 1484
rect 1708 1476 1716 1484
rect 1900 1476 1908 1484
rect 1916 1476 1924 1484
rect 2028 1476 2036 1484
rect 2076 1476 2084 1484
rect 2124 1476 2132 1484
rect 2252 1476 2260 1484
rect 2268 1476 2276 1484
rect 2348 1476 2356 1484
rect 2428 1476 2436 1484
rect 2444 1476 2452 1484
rect 2460 1476 2468 1484
rect 2508 1476 2516 1484
rect 2556 1476 2564 1484
rect 2588 1476 2596 1484
rect 2716 1476 2724 1484
rect 2764 1476 2772 1484
rect 2844 1476 2852 1484
rect 2860 1476 2868 1484
rect 3132 1476 3140 1484
rect 3244 1476 3252 1484
rect 3308 1496 3316 1504
rect 3452 1496 3460 1504
rect 3788 1516 3796 1524
rect 3836 1516 3844 1524
rect 3884 1516 3892 1524
rect 4060 1516 4068 1524
rect 4092 1516 4100 1524
rect 4172 1516 4180 1524
rect 4220 1516 4228 1524
rect 4252 1516 4260 1524
rect 3308 1476 3316 1484
rect 3388 1476 3396 1484
rect 3468 1476 3476 1484
rect 3516 1476 3524 1484
rect 3564 1476 3572 1484
rect 3612 1476 3620 1484
rect 3660 1476 3668 1484
rect 3756 1476 3764 1484
rect 3916 1476 3924 1484
rect 3932 1476 3940 1484
rect 3980 1476 3988 1484
rect 3996 1476 4004 1484
rect 4060 1476 4068 1484
rect 4140 1476 4148 1484
rect 4220 1476 4228 1484
rect 1260 1456 1268 1464
rect 1308 1456 1316 1464
rect 1356 1456 1364 1464
rect 1468 1456 1476 1464
rect 1532 1456 1540 1464
rect 1548 1456 1556 1464
rect 1628 1456 1636 1464
rect 1772 1456 1780 1464
rect 1788 1456 1796 1464
rect 2172 1456 2180 1464
rect 2188 1456 2196 1464
rect 2492 1456 2500 1464
rect 2540 1456 2548 1464
rect 2684 1456 2692 1464
rect 2748 1456 2756 1464
rect 2908 1456 2916 1464
rect 2988 1456 2996 1464
rect 3020 1456 3028 1464
rect 3100 1456 3108 1464
rect 3372 1456 3380 1464
rect 3484 1456 3492 1464
rect 3580 1456 3588 1464
rect 3964 1456 3972 1464
rect 4028 1456 4036 1464
rect 4092 1456 4100 1464
rect 4108 1456 4116 1464
rect 4188 1456 4196 1464
rect 124 1436 132 1444
rect 268 1436 276 1444
rect 332 1436 340 1444
rect 444 1436 452 1444
rect 652 1436 660 1444
rect 684 1436 692 1444
rect 828 1436 836 1444
rect 892 1436 900 1444
rect 1084 1436 1092 1444
rect 1116 1436 1124 1444
rect 1212 1436 1220 1444
rect 1372 1436 1380 1444
rect 1612 1436 1620 1444
rect 1644 1436 1652 1444
rect 1660 1436 1668 1444
rect 1724 1436 1732 1444
rect 1836 1436 1844 1444
rect 1996 1436 2004 1444
rect 2044 1436 2052 1444
rect 2092 1436 2100 1444
rect 2220 1436 2228 1444
rect 2364 1436 2372 1444
rect 2396 1436 2404 1444
rect 2572 1436 2580 1444
rect 2780 1436 2788 1444
rect 2828 1436 2836 1444
rect 2876 1436 2884 1444
rect 3228 1436 3236 1444
rect 3260 1436 3268 1444
rect 3340 1436 3348 1444
rect 3404 1436 3412 1444
rect 3532 1436 3540 1444
rect 3628 1436 3636 1444
rect 3708 1436 3716 1444
rect 4156 1436 4164 1444
rect 4236 1436 4244 1444
rect 12 1376 20 1384
rect 188 1376 196 1384
rect 444 1376 452 1384
rect 508 1376 516 1384
rect 572 1376 580 1384
rect 636 1376 644 1384
rect 844 1376 852 1384
rect 988 1376 996 1384
rect 1068 1376 1076 1384
rect 1180 1376 1188 1384
rect 1308 1376 1316 1384
rect 1436 1376 1444 1384
rect 1548 1376 1556 1384
rect 1788 1376 1796 1384
rect 1868 1376 1876 1384
rect 2124 1376 2132 1384
rect 2332 1376 2340 1384
rect 2412 1376 2420 1384
rect 2460 1376 2468 1384
rect 2508 1376 2516 1384
rect 2556 1376 2564 1384
rect 2652 1376 2660 1384
rect 2668 1376 2676 1384
rect 2812 1376 2820 1384
rect 3004 1376 3012 1384
rect 3100 1376 3108 1384
rect 3212 1376 3220 1384
rect 3244 1376 3252 1384
rect 3388 1376 3396 1384
rect 3580 1376 3588 1384
rect 3660 1376 3668 1384
rect 3724 1376 3732 1384
rect 3852 1376 3860 1384
rect 3948 1376 3956 1384
rect 3980 1376 3988 1384
rect 4044 1376 4052 1384
rect 76 1356 84 1364
rect 108 1356 116 1364
rect 140 1356 148 1364
rect 220 1356 228 1364
rect 364 1356 372 1364
rect 380 1356 388 1364
rect 396 1356 404 1364
rect 428 1356 436 1364
rect 460 1356 468 1364
rect 476 1356 484 1364
rect 556 1356 564 1364
rect 604 1356 612 1364
rect 732 1356 740 1364
rect 764 1356 772 1364
rect 796 1356 804 1364
rect 1020 1356 1028 1364
rect 1116 1356 1124 1364
rect 44 1336 52 1344
rect 124 1336 132 1344
rect 204 1336 212 1344
rect 252 1336 260 1344
rect 300 1336 308 1344
rect 540 1336 548 1344
rect 588 1336 596 1344
rect 652 1336 660 1344
rect 700 1336 708 1344
rect 748 1336 756 1344
rect 828 1336 836 1344
rect 876 1336 884 1344
rect 1020 1336 1028 1344
rect 1052 1336 1060 1344
rect 1100 1336 1108 1344
rect 1228 1356 1236 1364
rect 1468 1356 1476 1364
rect 1516 1356 1524 1364
rect 1564 1356 1572 1364
rect 1596 1356 1604 1364
rect 1756 1356 1764 1364
rect 1820 1356 1828 1364
rect 1836 1356 1844 1364
rect 1996 1356 2004 1364
rect 2012 1356 2020 1364
rect 2060 1356 2068 1364
rect 2204 1356 2212 1364
rect 2220 1356 2228 1364
rect 2268 1356 2276 1364
rect 2316 1356 2324 1364
rect 2348 1356 2356 1364
rect 2364 1356 2372 1364
rect 2540 1356 2548 1364
rect 2588 1356 2596 1364
rect 2780 1356 2788 1364
rect 2876 1356 2884 1364
rect 2908 1356 2916 1364
rect 2940 1356 2948 1364
rect 2956 1356 2964 1364
rect 2972 1356 2980 1364
rect 3068 1356 3076 1364
rect 3132 1356 3140 1364
rect 3228 1356 3236 1364
rect 3260 1356 3268 1364
rect 3340 1356 3348 1364
rect 3372 1356 3380 1364
rect 3548 1356 3556 1364
rect 3676 1356 3684 1364
rect 3756 1356 3764 1364
rect 3884 1356 3892 1364
rect 4076 1356 4084 1364
rect 4092 1356 4100 1364
rect 4124 1356 4132 1364
rect 4204 1356 4212 1364
rect 1228 1336 1236 1344
rect 1276 1336 1284 1344
rect 1340 1336 1348 1344
rect 1356 1336 1364 1344
rect 1404 1336 1412 1344
rect 1436 1336 1444 1344
rect 1484 1336 1492 1344
rect 1692 1336 1700 1344
rect 1804 1336 1812 1344
rect 1884 1336 1892 1344
rect 1900 1336 1908 1344
rect 1964 1336 1972 1344
rect 2044 1336 2052 1344
rect 2172 1336 2180 1344
rect 2188 1336 2196 1344
rect 2284 1336 2292 1344
rect 2428 1336 2436 1344
rect 2476 1336 2484 1344
rect 2540 1336 2548 1344
rect 2572 1336 2580 1344
rect 2620 1336 2628 1344
rect 2700 1336 2708 1344
rect 2748 1336 2756 1344
rect 2764 1336 2772 1344
rect 2844 1336 2852 1344
rect 2876 1336 2884 1344
rect 3036 1336 3044 1344
rect 3084 1336 3092 1344
rect 3196 1336 3204 1344
rect 3308 1336 3316 1344
rect 3420 1336 3428 1344
rect 3580 1336 3588 1344
rect 3612 1336 3620 1344
rect 3628 1336 3636 1344
rect 3820 1336 3828 1344
rect 3916 1336 3924 1344
rect 3964 1336 3972 1344
rect 4012 1336 4020 1344
rect 4156 1336 4164 1344
rect 12 1296 20 1304
rect 92 1296 100 1304
rect 220 1296 228 1304
rect 300 1296 308 1304
rect 620 1296 628 1304
rect 668 1296 676 1304
rect 796 1296 804 1304
rect 844 1296 852 1304
rect 924 1296 932 1304
rect 956 1296 964 1304
rect 972 1296 980 1304
rect 1004 1296 1012 1304
rect 1068 1296 1076 1304
rect 1180 1296 1188 1304
rect 1292 1296 1300 1304
rect 1308 1296 1316 1304
rect 1372 1296 1380 1304
rect 1388 1296 1396 1304
rect 1436 1296 1444 1304
rect 1484 1296 1492 1304
rect 1532 1296 1540 1304
rect 1628 1296 1636 1304
rect 1724 1296 1732 1304
rect 1772 1296 1780 1304
rect 1852 1296 1860 1304
rect 1932 1296 1940 1304
rect 2012 1296 2020 1304
rect 2124 1296 2132 1304
rect 2140 1296 2148 1304
rect 2172 1296 2180 1304
rect 2316 1296 2324 1304
rect 2396 1296 2404 1304
rect 2444 1296 2452 1304
rect 2492 1296 2500 1304
rect 2604 1296 2612 1304
rect 2652 1296 2660 1304
rect 2668 1296 2676 1304
rect 2700 1296 2708 1304
rect 2796 1296 2804 1304
rect 2812 1296 2820 1304
rect 2924 1296 2932 1304
rect 3004 1296 3012 1304
rect 3116 1296 3124 1304
rect 3164 1296 3172 1304
rect 3260 1296 3268 1304
rect 3388 1296 3396 1304
rect 3468 1296 3476 1304
rect 3580 1296 3588 1304
rect 3660 1296 3668 1304
rect 3788 1296 3796 1304
rect 3868 1296 3876 1304
rect 3900 1296 3908 1304
rect 3948 1296 3956 1304
rect 3996 1296 4004 1304
rect 44 1276 52 1284
rect 428 1276 436 1284
rect 940 1276 948 1284
rect 1228 1276 1236 1284
rect 1580 1276 1588 1284
rect 3036 1276 3044 1284
rect 3308 1276 3316 1284
rect 3452 1276 3460 1284
rect 2252 1256 2260 1264
rect 2988 1256 2996 1264
rect 780 1236 788 1244
rect 1612 1236 1620 1244
rect 1740 1236 1748 1244
rect 1980 1236 1988 1244
rect 2236 1236 2244 1244
rect 2380 1236 2388 1244
rect 2732 1236 2740 1244
rect 2860 1236 2868 1244
rect 3324 1236 3332 1244
rect 3356 1236 3364 1244
rect 4108 1236 4116 1244
rect 4140 1236 4148 1244
rect 4172 1236 4180 1244
rect 12 1176 20 1184
rect 220 1176 228 1184
rect 780 1176 788 1184
rect 924 1176 932 1184
rect 988 1176 996 1184
rect 1164 1176 1172 1184
rect 1180 1176 1188 1184
rect 1292 1176 1300 1184
rect 1756 1176 1764 1184
rect 2156 1176 2164 1184
rect 2316 1176 2324 1184
rect 2364 1176 2372 1184
rect 2572 1176 2580 1184
rect 2812 1176 2820 1184
rect 2892 1176 2900 1184
rect 3388 1176 3396 1184
rect 3420 1176 3428 1184
rect 3532 1176 3540 1184
rect 3724 1176 3732 1184
rect 3756 1176 3764 1184
rect 3788 1176 3796 1184
rect 4028 1176 4036 1184
rect 4252 1176 4260 1184
rect 1596 1156 1604 1164
rect 1916 1156 1924 1164
rect 2092 1156 2100 1164
rect 3452 1156 3460 1164
rect 44 1136 52 1144
rect 396 1136 404 1144
rect 716 1136 724 1144
rect 1004 1136 1012 1144
rect 1660 1136 1668 1144
rect 1804 1136 1812 1144
rect 2012 1136 2020 1144
rect 2140 1136 2148 1144
rect 2284 1136 2292 1144
rect 2396 1136 2404 1144
rect 4044 1136 4052 1144
rect 236 1116 244 1124
rect 284 1116 292 1124
rect 332 1116 340 1124
rect 412 1116 420 1124
rect 460 1116 468 1124
rect 508 1116 516 1124
rect 588 1116 596 1124
rect 636 1116 644 1124
rect 764 1116 772 1124
rect 844 1116 852 1124
rect 860 1116 868 1124
rect 972 1116 980 1124
rect 1052 1116 1060 1124
rect 1100 1116 1108 1124
rect 1244 1116 1252 1124
rect 1276 1116 1284 1124
rect 1324 1116 1332 1124
rect 1404 1116 1412 1124
rect 1452 1116 1460 1124
rect 1564 1116 1572 1124
rect 1612 1116 1620 1124
rect 1692 1116 1700 1124
rect 1708 1116 1716 1124
rect 1820 1116 1828 1124
rect 1932 1116 1940 1124
rect 1980 1116 1988 1124
rect 2076 1116 2084 1124
rect 2172 1116 2180 1124
rect 2412 1116 2420 1124
rect 2428 1116 2436 1124
rect 2476 1116 2484 1124
rect 2524 1116 2532 1124
rect 2636 1116 2644 1124
rect 2716 1116 2724 1124
rect 2764 1116 2772 1124
rect 2796 1116 2804 1124
rect 2876 1116 2884 1124
rect 2940 1116 2948 1124
rect 2956 1116 2964 1124
rect 2988 1116 2996 1124
rect 3084 1116 3092 1124
rect 3116 1116 3124 1124
rect 3132 1116 3140 1124
rect 3180 1116 3188 1124
rect 3372 1116 3380 1124
rect 3436 1116 3444 1124
rect 3484 1116 3492 1124
rect 3564 1116 3572 1124
rect 3612 1116 3620 1124
rect 3708 1116 3716 1124
rect 3740 1116 3748 1124
rect 3852 1116 3860 1124
rect 3900 1116 3908 1124
rect 3916 1116 3924 1124
rect 3996 1116 4004 1124
rect 4220 1116 4228 1124
rect 604 1096 612 1104
rect 76 1076 84 1084
rect 284 1076 292 1084
rect 316 1076 324 1084
rect 364 1076 372 1084
rect 492 1076 500 1084
rect 540 1076 548 1084
rect 556 1076 564 1084
rect 668 1076 676 1084
rect 732 1076 740 1084
rect 796 1076 804 1084
rect 892 1076 900 1084
rect 1132 1076 1140 1084
rect 1212 1076 1220 1084
rect 1452 1076 1460 1084
rect 1484 1076 1492 1084
rect 1532 1076 1540 1084
rect 1644 1076 1652 1084
rect 1660 1076 1668 1084
rect 1740 1076 1748 1084
rect 1852 1076 1860 1084
rect 1900 1076 1908 1084
rect 1964 1076 1972 1084
rect 1980 1076 1988 1084
rect 2028 1076 2036 1084
rect 2044 1076 2052 1084
rect 2220 1076 2228 1084
rect 2300 1076 2308 1084
rect 28 1056 36 1064
rect 92 1056 100 1064
rect 188 1056 196 1064
rect 204 1056 212 1064
rect 380 1056 388 1064
rect 524 1056 532 1064
rect 620 1056 628 1064
rect 796 1056 804 1064
rect 908 1056 916 1064
rect 1004 1056 1012 1064
rect 1148 1056 1156 1064
rect 1196 1056 1204 1064
rect 1244 1056 1252 1064
rect 1260 1056 1268 1064
rect 1468 1056 1476 1064
rect 1500 1056 1508 1064
rect 1516 1056 1524 1064
rect 1724 1056 1732 1064
rect 1772 1056 1780 1064
rect 1788 1056 1796 1064
rect 1868 1056 1876 1064
rect 1932 1056 1940 1064
rect 2108 1056 2116 1064
rect 2124 1056 2132 1064
rect 2236 1056 2244 1064
rect 2348 1076 2356 1084
rect 2380 1076 2388 1084
rect 2460 1076 2468 1084
rect 2556 1076 2564 1084
rect 2604 1076 2612 1084
rect 2620 1076 2628 1084
rect 2668 1076 2676 1084
rect 2684 1076 2692 1084
rect 2732 1076 2740 1084
rect 2828 1076 2836 1084
rect 2348 1056 2356 1064
rect 2476 1056 2484 1064
rect 2588 1056 2596 1064
rect 2652 1056 2660 1064
rect 2828 1056 2836 1064
rect 2860 1056 2868 1064
rect 2924 1076 2932 1084
rect 3004 1096 3012 1104
rect 3036 1076 3044 1084
rect 3084 1076 3092 1084
rect 3164 1076 3172 1084
rect 3276 1076 3284 1084
rect 3324 1076 3332 1084
rect 3404 1076 3412 1084
rect 3516 1076 3524 1084
rect 3612 1076 3620 1084
rect 3644 1076 3652 1084
rect 3660 1076 3668 1084
rect 3676 1076 3684 1084
rect 3708 1076 3716 1084
rect 3820 1076 3828 1084
rect 3868 1076 3876 1084
rect 3948 1076 3956 1084
rect 3964 1076 3972 1084
rect 2924 1056 2932 1064
rect 3004 1056 3012 1064
rect 3068 1056 3076 1064
rect 3100 1056 3108 1064
rect 3196 1056 3204 1064
rect 3212 1056 3220 1064
rect 3260 1056 3268 1064
rect 3292 1056 3300 1064
rect 3468 1056 3476 1064
rect 3548 1056 3556 1064
rect 3772 1056 3780 1064
rect 3804 1056 3812 1064
rect 3852 1056 3860 1064
rect 4012 1056 4020 1064
rect 4140 1076 4148 1084
rect 4188 1076 4196 1084
rect 4076 1056 4084 1064
rect 4156 1056 4164 1064
rect 4236 1056 4244 1064
rect 44 1036 52 1044
rect 124 1036 132 1044
rect 252 1036 260 1044
rect 284 1036 292 1044
rect 428 1036 436 1044
rect 588 1036 596 1044
rect 716 1036 724 1044
rect 764 1036 772 1044
rect 844 1036 852 1044
rect 860 1036 868 1044
rect 972 1036 980 1044
rect 1692 1036 1700 1044
rect 2076 1036 2084 1044
rect 2444 1036 2452 1044
rect 2716 1036 2724 1044
rect 2956 1036 2964 1044
rect 3148 1036 3156 1044
rect 3308 1036 3316 1044
rect 3436 1036 3444 1044
rect 3484 1036 3492 1044
rect 3580 1036 3588 1044
rect 3900 1036 3908 1044
rect 3916 1036 3924 1044
rect 3996 1036 4004 1044
rect 4108 1036 4116 1044
rect 4172 1036 4180 1044
rect 4204 1036 4212 1044
rect 28 976 36 984
rect 92 976 100 984
rect 204 976 212 984
rect 412 976 420 984
rect 444 976 452 984
rect 780 976 788 984
rect 876 976 884 984
rect 956 976 964 984
rect 1036 976 1044 984
rect 1148 976 1156 984
rect 1244 976 1252 984
rect 1356 976 1364 984
rect 1452 976 1460 984
rect 1644 976 1652 984
rect 1660 976 1668 984
rect 1756 976 1764 984
rect 1916 976 1924 984
rect 2044 976 2052 984
rect 2108 976 2116 984
rect 2204 976 2212 984
rect 2332 976 2340 984
rect 2780 976 2788 984
rect 2956 976 2964 984
rect 3004 976 3012 984
rect 3084 976 3092 984
rect 3180 976 3188 984
rect 3324 976 3332 984
rect 3500 976 3508 984
rect 3644 976 3652 984
rect 3724 976 3732 984
rect 3804 976 3812 984
rect 3836 976 3844 984
rect 3948 976 3956 984
rect 4044 976 4052 984
rect 4204 976 4212 984
rect 124 956 132 964
rect 156 956 164 964
rect 188 956 196 964
rect 252 956 260 964
rect 300 956 308 964
rect 348 956 356 964
rect 364 956 372 964
rect 460 956 468 964
rect 492 956 500 964
rect 508 956 516 964
rect 588 956 596 964
rect 620 956 628 964
rect 652 956 660 964
rect 892 956 900 964
rect 908 956 916 964
rect 1276 956 1284 964
rect 1388 956 1396 964
rect 1404 956 1412 964
rect 1484 956 1492 964
rect 1676 956 1684 964
rect 1708 956 1716 964
rect 1788 956 1796 964
rect 1820 956 1828 964
rect 2028 956 2036 964
rect 2252 956 2260 964
rect 2284 956 2292 964
rect 2412 956 2420 964
rect 2444 956 2452 964
rect 2572 956 2580 964
rect 2604 956 2612 964
rect 2732 956 2740 964
rect 2812 956 2820 964
rect 2828 956 2836 964
rect 2860 956 2868 964
rect 2908 956 2916 964
rect 3036 956 3044 964
rect 3132 956 3140 964
rect 3564 956 3572 964
rect 3852 956 3860 964
rect 3980 956 3988 964
rect 3996 956 4004 964
rect 4124 956 4132 964
rect 4156 956 4164 964
rect 12 936 20 944
rect 60 936 68 944
rect 236 936 244 944
rect 428 936 436 944
rect 684 936 692 944
rect 764 936 772 944
rect 812 936 820 944
rect 828 936 836 944
rect 972 936 980 944
rect 988 936 996 944
rect 1068 936 1076 944
rect 1084 936 1092 944
rect 1132 936 1140 944
rect 1212 936 1220 944
rect 44 896 52 904
rect 92 896 100 904
rect 396 896 404 904
rect 668 896 676 904
rect 716 896 724 904
rect 748 916 756 924
rect 764 896 772 904
rect 860 896 868 904
rect 940 896 948 904
rect 1020 896 1028 904
rect 1116 916 1124 924
rect 1308 936 1316 944
rect 1436 936 1444 944
rect 1548 936 1556 944
rect 1564 936 1572 944
rect 1612 936 1620 944
rect 1692 936 1700 944
rect 1740 936 1748 944
rect 1900 936 1908 944
rect 1948 936 1956 944
rect 1980 936 1988 944
rect 2076 936 2084 944
rect 2092 936 2100 944
rect 2140 936 2148 944
rect 2188 936 2196 944
rect 2220 936 2228 944
rect 2300 936 2308 944
rect 2348 936 2356 944
rect 2364 936 2372 944
rect 2380 936 2388 944
rect 2460 936 2468 944
rect 2476 936 2484 944
rect 2620 936 2628 944
rect 2668 936 2676 944
rect 2748 936 2756 944
rect 2892 936 2900 944
rect 2972 936 2980 944
rect 2988 936 2996 944
rect 3148 936 3156 944
rect 3196 936 3204 944
rect 3244 936 3252 944
rect 3356 936 3364 944
rect 3452 936 3460 944
rect 3468 936 3476 944
rect 3516 936 3524 944
rect 3628 936 3636 944
rect 3676 936 3684 944
rect 3692 936 3700 944
rect 3772 936 3780 944
rect 3788 936 3796 944
rect 3868 936 3876 944
rect 3884 936 3892 944
rect 3916 936 3924 944
rect 4028 936 4036 944
rect 4060 936 4068 944
rect 4092 936 4100 944
rect 4108 936 4116 944
rect 4220 936 4228 944
rect 1516 916 1524 924
rect 1964 916 1972 924
rect 2252 916 2260 924
rect 2604 916 2612 924
rect 3356 916 3364 924
rect 3596 916 3604 924
rect 3644 916 3652 924
rect 1132 896 1140 904
rect 1164 896 1172 904
rect 1180 896 1188 904
rect 1260 896 1268 904
rect 1276 896 1284 904
rect 1356 896 1364 904
rect 1484 896 1492 904
rect 1516 896 1524 904
rect 1596 896 1604 904
rect 1644 896 1652 904
rect 1724 896 1732 904
rect 1772 896 1780 904
rect 1884 896 1892 904
rect 1932 896 1940 904
rect 1980 896 1988 904
rect 2028 896 2036 904
rect 2044 896 2052 904
rect 2124 896 2132 904
rect 2172 896 2180 904
rect 2188 896 2196 904
rect 2332 896 2340 904
rect 2380 896 2388 904
rect 2428 896 2436 904
rect 2524 896 2532 904
rect 2572 896 2580 904
rect 2652 896 2660 904
rect 2684 896 2692 904
rect 2860 896 2868 904
rect 2940 896 2948 904
rect 3020 896 3028 904
rect 3180 896 3188 904
rect 3196 896 3204 904
rect 3228 896 3236 904
rect 3276 896 3284 904
rect 3372 896 3380 904
rect 3420 896 3428 904
rect 3500 896 3508 904
rect 3532 896 3540 904
rect 3548 896 3556 904
rect 3596 896 3604 904
rect 3644 896 3652 904
rect 3740 896 3748 904
rect 3820 896 3828 904
rect 3916 896 3924 904
rect 4028 896 4036 904
rect 4076 896 4084 904
rect 124 876 132 884
rect 364 876 372 884
rect 2668 876 2676 884
rect 2828 876 2836 884
rect 2908 876 2916 884
rect 3452 876 3460 884
rect 3724 876 3732 884
rect 1532 856 1540 864
rect 1580 856 1588 864
rect 108 836 116 844
rect 476 836 484 844
rect 556 836 564 844
rect 636 836 644 844
rect 844 836 852 844
rect 924 836 932 844
rect 1372 836 1380 844
rect 1420 836 1428 844
rect 1804 836 1812 844
rect 1868 836 1876 844
rect 2268 836 2276 844
rect 2540 836 2548 844
rect 2556 836 2564 844
rect 3308 836 3316 844
rect 4140 836 4148 844
rect 12 776 20 784
rect 140 776 148 784
rect 428 776 436 784
rect 876 776 884 784
rect 892 776 900 784
rect 1580 776 1588 784
rect 1676 776 1684 784
rect 1996 776 2004 784
rect 2348 776 2356 784
rect 2844 776 2852 784
rect 3036 776 3044 784
rect 3164 776 3172 784
rect 3244 776 3252 784
rect 3564 776 3572 784
rect 3644 776 3652 784
rect 3660 776 3668 784
rect 3900 776 3908 784
rect 3964 776 3972 784
rect 4060 776 4068 784
rect 4220 776 4228 784
rect 668 756 676 764
rect 1068 756 1076 764
rect 1692 756 1700 764
rect 2572 756 2580 764
rect 924 736 932 744
rect 1292 736 1300 744
rect 1852 736 1860 744
rect 2188 736 2196 744
rect 2236 736 2244 744
rect 2300 736 2308 744
rect 3436 736 3444 744
rect 44 716 52 724
rect 188 716 196 724
rect 204 716 212 724
rect 364 716 372 724
rect 508 716 516 724
rect 556 716 564 724
rect 652 716 660 724
rect 844 716 852 724
rect 1052 716 1060 724
rect 1116 716 1124 724
rect 1164 716 1172 724
rect 1244 716 1252 724
rect 1372 716 1380 724
rect 1436 716 1444 724
rect 1484 716 1492 724
rect 1644 716 1652 724
rect 1724 716 1732 724
rect 1772 716 1780 724
rect 1884 716 1892 724
rect 1932 716 1940 724
rect 1948 716 1956 724
rect 2108 716 2116 724
rect 2140 716 2148 724
rect 2156 716 2164 724
rect 2204 716 2212 724
rect 2316 716 2324 724
rect 2364 716 2372 724
rect 2412 716 2420 724
rect 2460 716 2468 724
rect 2476 716 2484 724
rect 2524 716 2532 724
rect 2636 716 2644 724
rect 2668 716 2676 724
rect 2764 716 2772 724
rect 2876 716 2884 724
rect 2988 716 2996 724
rect 3020 716 3028 724
rect 3052 716 3060 724
rect 3116 716 3124 724
rect 3228 716 3236 724
rect 3276 716 3284 724
rect 3356 716 3364 724
rect 3404 716 3412 724
rect 3452 716 3460 724
rect 3500 716 3508 724
rect 3628 716 3636 724
rect 3724 716 3732 724
rect 3740 716 3748 724
rect 3820 716 3828 724
rect 3868 716 3876 724
rect 3948 716 3956 724
rect 4028 716 4036 724
rect 4108 716 4116 724
rect 4188 716 4196 724
rect 828 696 836 704
rect 1036 696 1044 704
rect 1084 696 1092 704
rect 1260 696 1268 704
rect 2924 696 2932 704
rect 156 676 164 684
rect 236 676 244 684
rect 396 676 404 684
rect 604 676 612 684
rect 620 676 628 684
rect 700 676 708 684
rect 812 676 820 684
rect 956 676 964 684
rect 1148 676 1156 684
rect 1276 676 1284 684
rect 1324 676 1332 684
rect 1404 676 1412 684
rect 1452 676 1460 684
rect 1484 676 1492 684
rect 1612 676 1620 684
rect 1756 676 1764 684
rect 1804 676 1812 684
rect 1836 676 1844 684
rect 1900 676 1908 684
rect 1964 676 1972 684
rect 1980 676 1988 684
rect 2092 676 2100 684
rect 2140 676 2148 684
rect 2188 676 2196 684
rect 2236 676 2244 684
rect 2284 676 2292 684
rect 2332 676 2340 684
rect 2380 676 2388 684
rect 2508 676 2516 684
rect 2556 676 2564 684
rect 2604 676 2612 684
rect 2716 676 2724 684
rect 2908 676 2916 684
rect 2956 676 2964 684
rect 3100 676 3108 684
rect 3132 676 3140 684
rect 3148 676 3156 684
rect 3196 676 3204 684
rect 3308 676 3316 684
rect 3372 676 3380 684
rect 3420 676 3428 684
rect 3468 676 3476 684
rect 3580 676 3588 684
rect 3628 676 3636 684
rect 3676 676 3684 684
rect 3772 676 3780 684
rect 3788 676 3796 684
rect 3836 676 3844 684
rect 3916 676 3924 684
rect 4108 676 4116 684
rect 4140 676 4148 684
rect 4156 676 4164 684
rect 108 656 116 664
rect 124 656 132 664
rect 220 656 228 664
rect 252 656 260 664
rect 348 656 356 664
rect 364 656 372 664
rect 412 656 420 664
rect 444 656 452 664
rect 652 656 660 664
rect 684 656 692 664
rect 764 656 772 664
rect 796 656 804 664
rect 860 656 868 664
rect 908 656 916 664
rect 972 656 980 664
rect 1052 656 1060 664
rect 1100 656 1108 664
rect 1228 656 1236 664
rect 1308 656 1316 664
rect 1372 656 1380 664
rect 1388 656 1396 664
rect 1564 656 1572 664
rect 1596 656 1604 664
rect 1644 656 1652 664
rect 1660 656 1668 664
rect 1836 656 1844 664
rect 1884 656 1892 664
rect 2012 656 2020 664
rect 2028 656 2036 664
rect 2060 656 2068 664
rect 2268 656 2276 664
rect 2588 656 2596 664
rect 2652 656 2660 664
rect 2668 656 2676 664
rect 2828 656 2836 664
rect 2860 656 2868 664
rect 2940 656 2948 664
rect 3180 656 3188 664
rect 3260 656 3268 664
rect 3340 656 3348 664
rect 3516 656 3524 664
rect 3548 656 3556 664
rect 3628 656 3636 664
rect 3676 656 3684 664
rect 3740 656 3748 664
rect 3852 656 3860 664
rect 3884 656 3892 664
rect 3980 656 3988 664
rect 4044 656 4052 664
rect 4076 656 4084 664
rect 4108 656 4116 664
rect 12 636 20 644
rect 172 636 180 644
rect 300 636 308 644
rect 524 636 532 644
rect 716 636 724 644
rect 780 636 788 644
rect 924 636 932 644
rect 1132 636 1140 644
rect 1164 636 1172 644
rect 1356 636 1364 644
rect 1420 636 1428 644
rect 1468 636 1476 644
rect 1532 636 1540 644
rect 1788 636 1796 644
rect 1916 636 1924 644
rect 2044 636 2052 644
rect 2204 636 2212 644
rect 2460 636 2468 644
rect 2492 636 2500 644
rect 2524 636 2532 644
rect 2636 636 2644 644
rect 2684 636 2692 644
rect 2732 636 2740 644
rect 2876 636 2884 644
rect 3228 636 3236 644
rect 3404 636 3412 644
rect 3500 636 3508 644
rect 3532 636 3540 644
rect 3724 636 3732 644
rect 3804 636 3812 644
rect 3932 636 3940 644
rect 4028 636 4036 644
rect 124 576 132 584
rect 284 576 292 584
rect 572 576 580 584
rect 828 576 836 584
rect 908 576 916 584
rect 1308 576 1316 584
rect 1372 576 1380 584
rect 1500 576 1508 584
rect 1596 576 1604 584
rect 1836 576 1844 584
rect 1884 576 1892 584
rect 2012 576 2020 584
rect 2220 576 2228 584
rect 2300 576 2308 584
rect 2380 576 2388 584
rect 2444 576 2452 584
rect 2876 576 2884 584
rect 2892 576 2900 584
rect 3036 576 3044 584
rect 3084 576 3092 584
rect 3116 576 3124 584
rect 3180 576 3188 584
rect 3276 576 3284 584
rect 3372 576 3380 584
rect 3596 576 3604 584
rect 3628 576 3636 584
rect 3948 576 3956 584
rect 3980 576 3988 584
rect 4044 576 4052 584
rect 4140 576 4148 584
rect 156 556 164 564
rect 172 556 180 564
rect 332 556 340 564
rect 364 556 372 564
rect 460 556 468 564
rect 492 556 500 564
rect 604 556 612 564
rect 620 556 628 564
rect 636 556 644 564
rect 700 556 708 564
rect 716 556 724 564
rect 780 556 788 564
rect 812 556 820 564
rect 844 556 852 564
rect 860 556 868 564
rect 940 556 948 564
rect 988 556 996 564
rect 1004 556 1012 564
rect 1020 556 1028 564
rect 1388 556 1396 564
rect 1548 556 1556 564
rect 1644 556 1652 564
rect 1852 556 1860 564
rect 1916 556 1924 564
rect 1948 556 1956 564
rect 1980 556 1988 564
rect 1996 556 2004 564
rect 2188 556 2196 564
rect 2268 556 2276 564
rect 2284 556 2292 564
rect 2428 556 2436 564
rect 2668 556 2676 564
rect 2748 556 2756 564
rect 2812 556 2820 564
rect 2956 556 2964 564
rect 3004 556 3012 564
rect 3228 556 3236 564
rect 3260 556 3268 564
rect 3420 556 3428 564
rect 3564 556 3572 564
rect 3788 556 3796 564
rect 3836 556 3844 564
rect 3852 556 3860 564
rect 3964 556 3972 564
rect 4124 556 4132 564
rect 12 536 20 544
rect 92 536 100 544
rect 124 536 132 544
rect 268 536 276 544
rect 316 536 324 544
rect 380 536 388 544
rect 428 536 436 544
rect 460 536 468 544
rect 556 536 564 544
rect 588 536 596 544
rect 668 536 676 544
rect 748 536 756 544
rect 796 536 804 544
rect 1068 536 1076 544
rect 1116 536 1124 544
rect 1132 536 1140 544
rect 1212 536 1220 544
rect 1324 536 1332 544
rect 1340 536 1348 544
rect 1420 536 1428 544
rect 1484 536 1492 544
rect 1532 536 1540 544
rect 1580 536 1588 544
rect 1628 536 1636 544
rect 1740 536 1748 544
rect 1820 536 1828 544
rect 1900 536 1908 544
rect 2076 536 2084 544
rect 2156 536 2164 544
rect 2236 536 2244 544
rect 2348 536 2356 544
rect 2508 536 2516 544
rect 2524 536 2532 544
rect 2668 536 2676 544
rect 2780 536 2788 544
rect 2796 536 2804 544
rect 2844 536 2852 544
rect 2972 536 2980 544
rect 3020 536 3028 544
rect 3100 536 3108 544
rect 3148 536 3156 544
rect 3164 536 3172 544
rect 3308 536 3316 544
rect 3356 536 3364 544
rect 3404 536 3412 544
rect 3484 536 3492 544
rect 3532 536 3540 544
rect 3580 536 3588 544
rect 3660 536 3668 544
rect 3708 536 3716 544
rect 3724 536 3732 544
rect 3804 536 3812 544
rect 3884 536 3892 544
rect 3932 536 3940 544
rect 4028 536 4036 544
rect 4060 536 4068 544
rect 4108 536 4116 544
rect 1932 516 1940 524
rect 2844 516 2852 524
rect 3308 516 3316 524
rect 3468 516 3476 524
rect 3900 516 3908 524
rect 44 496 52 504
rect 124 496 132 504
rect 188 496 196 504
rect 220 496 228 504
rect 284 496 292 504
rect 396 496 404 504
rect 428 496 436 504
rect 492 496 500 504
rect 636 496 644 504
rect 716 496 724 504
rect 940 496 948 504
rect 972 496 980 504
rect 1036 496 1044 504
rect 1084 496 1092 504
rect 1132 496 1140 504
rect 1164 496 1172 504
rect 1244 496 1252 504
rect 1436 496 1444 504
rect 1500 496 1508 504
rect 1548 496 1556 504
rect 1596 496 1604 504
rect 1708 496 1716 504
rect 1740 496 1748 504
rect 1788 496 1796 504
rect 1868 496 1876 504
rect 2044 496 2052 504
rect 2124 496 2132 504
rect 2204 496 2212 504
rect 2476 496 2484 504
rect 2556 496 2564 504
rect 2604 496 2612 504
rect 2684 496 2692 504
rect 2764 496 2772 504
rect 2876 496 2884 504
rect 2892 496 2900 504
rect 3004 496 3012 504
rect 3052 496 3060 504
rect 3116 496 3124 504
rect 3276 496 3284 504
rect 3324 496 3332 504
rect 3372 496 3380 504
rect 3500 496 3508 504
rect 3612 496 3620 504
rect 3628 496 3636 504
rect 3676 496 3684 504
rect 3724 496 3732 504
rect 3756 496 3764 504
rect 3836 496 3844 504
rect 3852 496 3860 504
rect 3964 496 3972 504
rect 4012 496 4020 504
rect 4076 496 4084 504
rect 4188 496 4196 504
rect 364 476 372 484
rect 668 476 676 484
rect 1068 476 1076 484
rect 1388 476 1396 484
rect 1404 476 1412 484
rect 2284 476 2292 484
rect 2348 476 2356 484
rect 3532 476 3540 484
rect 2092 456 2100 464
rect 3244 456 3252 464
rect 3740 456 3748 464
rect 3772 456 3780 464
rect 76 436 84 444
rect 204 436 212 444
rect 412 436 420 444
rect 572 436 580 444
rect 764 436 772 444
rect 956 436 964 444
rect 1196 436 1204 444
rect 1660 436 1668 444
rect 1676 436 1684 444
rect 1964 436 1972 444
rect 2172 436 2180 444
rect 2332 436 2340 444
rect 2636 436 2644 444
rect 2652 436 2660 444
rect 3548 436 3556 444
rect 4220 436 4228 444
rect 172 376 180 384
rect 300 376 308 384
rect 1244 376 1252 384
rect 1356 376 1364 384
rect 1452 376 1460 384
rect 1740 376 1748 384
rect 1788 376 1796 384
rect 2844 376 2852 384
rect 3148 376 3156 384
rect 3180 376 3188 384
rect 3452 376 3460 384
rect 3868 376 3876 384
rect 4108 376 4116 384
rect 4236 376 4244 384
rect 364 356 372 364
rect 1724 356 1732 364
rect 3500 356 3508 364
rect 3612 356 3620 364
rect 412 336 420 344
rect 796 336 804 344
rect 1804 336 1812 344
rect 2092 336 2100 344
rect 2684 336 2692 344
rect 3548 336 3556 344
rect 3772 336 3780 344
rect 44 316 52 324
rect 60 316 68 324
rect 108 316 116 324
rect 188 316 196 324
rect 204 316 212 324
rect 252 316 260 324
rect 428 316 436 324
rect 460 316 468 324
rect 588 316 596 324
rect 604 316 612 324
rect 652 316 660 324
rect 812 316 820 324
rect 860 316 868 324
rect 892 316 900 324
rect 956 316 964 324
rect 1004 316 1012 324
rect 1132 316 1140 324
rect 1228 316 1236 324
rect 1260 316 1268 324
rect 1484 316 1492 324
rect 1532 316 1540 324
rect 1612 316 1620 324
rect 1692 316 1700 324
rect 1996 316 2004 324
rect 2204 316 2212 324
rect 2220 316 2228 324
rect 2284 316 2292 324
rect 2364 316 2372 324
rect 2556 316 2564 324
rect 2636 316 2644 324
rect 2732 316 2740 324
rect 2764 316 2772 324
rect 2892 316 2900 324
rect 2940 316 2948 324
rect 2988 316 2996 324
rect 3036 316 3044 324
rect 3116 316 3124 324
rect 3164 316 3172 324
rect 3212 316 3220 324
rect 3260 316 3268 324
rect 3292 316 3300 324
rect 3388 316 3396 324
rect 3436 316 3444 324
rect 3596 316 3604 324
rect 3644 316 3652 324
rect 3692 316 3700 324
rect 3708 316 3716 324
rect 3804 316 3812 324
rect 3820 316 3828 324
rect 3964 316 3972 324
rect 4092 316 4100 324
rect 4220 316 4228 324
rect 2204 296 2212 304
rect 12 276 20 284
rect 92 276 100 284
rect 140 276 148 284
rect 156 276 164 284
rect 236 276 244 284
rect 284 276 292 284
rect 332 276 340 284
rect 252 256 260 264
rect 316 256 324 264
rect 332 256 340 264
rect 396 276 404 284
rect 508 276 516 284
rect 700 276 708 284
rect 764 276 772 284
rect 844 276 852 284
rect 940 276 948 284
rect 988 276 996 284
rect 1036 276 1044 284
rect 1052 276 1060 284
rect 1164 276 1172 284
rect 1180 276 1188 284
rect 1292 276 1300 284
rect 1372 276 1380 284
rect 1516 276 1524 284
rect 1644 276 1652 284
rect 1660 276 1668 284
rect 1852 276 1860 284
rect 1916 276 1924 284
rect 2092 276 2100 284
rect 2604 296 2612 304
rect 3916 296 3924 304
rect 2604 276 2612 284
rect 2652 276 2660 284
rect 2764 276 2772 284
rect 2812 276 2820 284
rect 2860 276 2868 284
rect 2940 276 2948 284
rect 2972 276 2980 284
rect 3020 276 3028 284
rect 3068 276 3076 284
rect 3084 276 3092 284
rect 3132 276 3140 284
rect 3244 276 3252 284
rect 3292 276 3300 284
rect 3340 276 3348 284
rect 3356 276 3364 284
rect 3404 276 3412 284
rect 3516 276 3524 284
rect 3564 276 3572 284
rect 3676 276 3684 284
rect 3724 276 3732 284
rect 3772 276 3780 284
rect 3852 276 3860 284
rect 3932 276 3940 284
rect 4124 276 4132 284
rect 396 256 404 264
rect 524 256 532 264
rect 620 256 628 264
rect 700 256 708 264
rect 732 256 740 264
rect 780 256 788 264
rect 1116 256 1124 264
rect 1228 256 1236 264
rect 1260 256 1268 264
rect 1308 256 1316 264
rect 1324 256 1332 264
rect 1340 256 1348 264
rect 1436 256 1444 264
rect 1468 256 1476 264
rect 1500 256 1508 264
rect 1596 256 1604 264
rect 1756 256 1764 264
rect 1772 256 1780 264
rect 1852 256 1860 264
rect 1932 256 1940 264
rect 2044 256 2052 264
rect 2156 256 2164 264
rect 2172 256 2180 264
rect 2348 256 2356 264
rect 2428 256 2436 264
rect 2444 256 2452 264
rect 2540 256 2548 264
rect 2716 256 2724 264
rect 2780 256 2788 264
rect 2828 256 2836 264
rect 2908 256 2916 264
rect 3164 256 3172 264
rect 3196 256 3204 264
rect 3468 256 3476 264
rect 3484 256 3492 264
rect 3596 256 3604 264
rect 3628 256 3636 264
rect 3740 256 3748 264
rect 3884 256 3892 264
rect 3900 256 3908 264
rect 4076 256 4084 264
rect 4140 256 4148 264
rect 4220 256 4228 264
rect 44 236 52 244
rect 76 236 84 244
rect 124 236 132 244
rect 204 236 212 244
rect 428 236 436 244
rect 588 236 596 244
rect 828 236 836 244
rect 860 236 868 244
rect 956 236 964 244
rect 1004 236 1012 244
rect 1084 236 1092 244
rect 1148 236 1156 244
rect 1196 236 1204 244
rect 1404 236 1412 244
rect 1532 236 1540 244
rect 1628 236 1636 244
rect 1820 236 1828 244
rect 1884 236 1892 244
rect 2092 236 2100 244
rect 2380 236 2388 244
rect 2508 236 2516 244
rect 2572 236 2580 244
rect 2620 236 2628 244
rect 2684 236 2692 244
rect 2732 236 2740 244
rect 2876 236 2884 244
rect 2940 236 2948 244
rect 2988 236 2996 244
rect 3036 236 3044 244
rect 3100 236 3108 244
rect 3212 236 3220 244
rect 3276 236 3284 244
rect 3324 236 3332 244
rect 3372 236 3380 244
rect 3420 236 3428 244
rect 3532 236 3540 244
rect 3644 236 3652 244
rect 3804 236 3812 244
rect 3820 236 3828 244
rect 4044 236 4052 244
rect 4188 236 4196 244
rect 12 176 20 184
rect 220 176 228 184
rect 332 176 340 184
rect 412 176 420 184
rect 492 176 500 184
rect 684 176 692 184
rect 1116 176 1124 184
rect 1340 176 1348 184
rect 1372 176 1380 184
rect 1500 176 1508 184
rect 1580 176 1588 184
rect 1612 176 1620 184
rect 1660 176 1668 184
rect 1756 176 1764 184
rect 1772 176 1780 184
rect 1884 176 1892 184
rect 1932 176 1940 184
rect 2092 176 2100 184
rect 2428 176 2436 184
rect 2636 176 2644 184
rect 2748 176 2756 184
rect 3196 176 3204 184
rect 3308 176 3316 184
rect 3388 176 3396 184
rect 3580 176 3588 184
rect 3644 176 3652 184
rect 3724 176 3732 184
rect 3772 176 3780 184
rect 3884 176 3892 184
rect 4012 176 4020 184
rect 4108 176 4116 184
rect 4204 176 4212 184
rect 92 156 100 164
rect 172 156 180 164
rect 268 156 276 164
rect 300 156 308 164
rect 380 156 388 164
rect 444 156 452 164
rect 540 156 548 164
rect 620 156 628 164
rect 636 156 644 164
rect 732 156 740 164
rect 860 156 868 164
rect 876 156 884 164
rect 1100 156 1108 164
rect 1212 156 1220 164
rect 1260 156 1268 164
rect 1292 156 1300 164
rect 1388 156 1396 164
rect 1420 156 1428 164
rect 1452 156 1460 164
rect 1548 156 1556 164
rect 1628 156 1636 164
rect 1708 156 1716 164
rect 1836 156 1844 164
rect 1868 156 1876 164
rect 1900 156 1908 164
rect 2028 156 2036 164
rect 2044 156 2052 164
rect 2124 156 2132 164
rect 2156 156 2164 164
rect 2252 156 2260 164
rect 2460 156 2468 164
rect 2524 156 2532 164
rect 2588 156 2596 164
rect 2620 156 2628 164
rect 2700 156 2708 164
rect 2844 156 2852 164
rect 2908 156 2916 164
rect 2940 156 2948 164
rect 2956 156 2964 164
rect 3004 156 3012 164
rect 3244 156 3252 164
rect 3260 156 3268 164
rect 3356 156 3364 164
rect 3420 156 3428 164
rect 3452 156 3460 164
rect 3516 156 3524 164
rect 3548 156 3556 164
rect 3612 156 3620 164
rect 3756 156 3764 164
rect 3788 156 3796 164
rect 3804 156 3812 164
rect 3836 156 3844 164
rect 3852 156 3860 164
rect 3932 156 3940 164
rect 3948 156 3956 164
rect 4028 156 4036 164
rect 4124 156 4132 164
rect 92 136 100 144
rect 124 136 132 144
rect 140 136 148 144
rect 428 136 436 144
rect 780 136 788 144
rect 540 116 548 124
rect 940 136 948 144
rect 1148 136 1156 144
rect 1196 136 1204 144
rect 1276 136 1284 144
rect 1356 136 1364 144
rect 1388 136 1396 144
rect 1244 116 1252 124
rect 44 96 52 104
rect 124 96 132 104
rect 156 96 164 104
rect 396 96 404 104
rect 556 96 564 104
rect 732 96 740 104
rect 812 96 820 104
rect 908 96 916 104
rect 1004 96 1012 104
rect 1052 96 1060 104
rect 1116 96 1124 104
rect 1164 96 1172 104
rect 1180 96 1188 104
rect 1244 96 1252 104
rect 1420 96 1428 104
rect 1468 136 1476 144
rect 1596 136 1604 144
rect 1724 136 1732 144
rect 1804 136 1812 144
rect 1836 136 1844 144
rect 1916 136 1924 144
rect 1964 136 1972 144
rect 2108 136 2116 144
rect 2300 136 2308 144
rect 1948 116 1956 124
rect 2508 136 2516 144
rect 2556 136 2564 144
rect 2716 136 2724 144
rect 2764 136 2772 144
rect 3004 136 3012 144
rect 3036 136 3044 144
rect 3116 136 3124 144
rect 3132 136 3140 144
rect 3148 136 3156 144
rect 3180 136 3188 144
rect 3372 136 3380 144
rect 3468 136 3476 144
rect 3484 136 3492 144
rect 3596 136 3604 144
rect 3676 136 3684 144
rect 3692 136 3700 144
rect 4076 136 4084 144
rect 4172 136 4180 144
rect 4188 136 4196 144
rect 2556 116 2564 124
rect 2908 116 2916 124
rect 3452 116 3460 124
rect 4188 116 4196 124
rect 1468 96 1476 104
rect 1516 96 1524 104
rect 1564 96 1572 104
rect 1644 96 1652 104
rect 1756 96 1764 104
rect 1772 96 1780 104
rect 1948 96 1956 104
rect 1996 96 2004 104
rect 2204 96 2212 104
rect 2252 96 2260 104
rect 2348 96 2356 104
rect 2476 96 2484 104
rect 2748 96 2756 104
rect 2796 96 2804 104
rect 2956 96 2964 104
rect 3036 96 3044 104
rect 3068 96 3076 104
rect 3084 96 3092 104
rect 3100 96 3108 104
rect 3164 96 3172 104
rect 3404 96 3412 104
rect 3564 96 3572 104
rect 3820 96 3828 104
rect 3852 96 3860 104
rect 4012 96 4020 104
rect 4092 96 4100 104
rect 4140 96 4148 104
rect 4220 96 4228 104
rect 892 76 900 84
rect 1532 76 1540 84
rect 1804 76 1812 84
rect 2012 76 2020 84
rect 2156 76 2164 84
rect 3052 56 3060 64
<< metal2 >>
rect 141 2964 147 3083
rect 1581 2984 1587 3083
rect 596 2977 627 2983
rect 429 2964 435 2976
rect 141 2944 147 2956
rect 221 2904 227 2936
rect 93 2744 99 2876
rect 157 2724 163 2736
rect 237 2724 243 2956
rect 269 2803 275 2956
rect 381 2944 387 2956
rect 445 2943 451 2976
rect 509 2963 515 2976
rect 621 2964 627 2977
rect 733 2964 739 2976
rect 1709 2964 1715 2976
rect 509 2957 540 2963
rect 1380 2957 1388 2963
rect 1412 2957 1420 2963
rect 461 2944 467 2956
rect 605 2944 611 2956
rect 877 2944 883 2956
rect 436 2937 451 2943
rect 365 2804 371 2836
rect 253 2797 275 2803
rect 237 2704 243 2716
rect 253 2684 259 2797
rect 285 2724 291 2736
rect 333 2724 339 2796
rect 333 2684 339 2716
rect 381 2704 387 2936
rect 413 2904 419 2936
rect 493 2924 499 2936
rect 493 2744 499 2916
rect 525 2904 531 2936
rect 525 2804 531 2896
rect 13 2664 19 2676
rect 77 2664 83 2676
rect 173 2664 179 2676
rect 493 2664 499 2696
rect 509 2684 515 2796
rect 541 2724 547 2876
rect 541 2684 547 2716
rect 589 2704 595 2716
rect 621 2684 627 2736
rect 669 2704 675 2716
rect 701 2704 707 2876
rect 701 2684 707 2696
rect 749 2684 755 2736
rect 797 2724 803 2896
rect 845 2764 851 2896
rect 893 2784 899 2936
rect 957 2804 963 2956
rect 1757 2944 1763 2976
rect 1837 2944 1843 2956
rect 1997 2944 2003 2976
rect 2061 2944 2067 3083
rect 2525 2984 2531 2996
rect 2260 2957 2275 2963
rect 1508 2937 1516 2943
rect 1005 2904 1011 2936
rect 765 2684 771 2716
rect 797 2704 803 2716
rect 877 2704 883 2716
rect 925 2684 931 2796
rect 1005 2704 1011 2896
rect 1021 2804 1027 2936
rect 1053 2884 1059 2896
rect 1037 2724 1043 2856
rect 1181 2784 1187 2796
rect 1101 2724 1107 2736
rect 1197 2724 1203 2836
rect 1229 2804 1235 2896
rect 1261 2704 1267 2836
rect 1309 2784 1315 2896
rect 1421 2824 1427 2896
rect 1341 2784 1347 2816
rect 1469 2784 1475 2896
rect 1549 2884 1555 2936
rect 1581 2904 1587 2936
rect 1677 2924 1683 2936
rect 1613 2917 1651 2923
rect 1533 2844 1539 2856
rect 1597 2804 1603 2896
rect 1613 2884 1619 2917
rect 1645 2903 1651 2917
rect 1645 2897 1708 2903
rect 1629 2884 1635 2896
rect 1805 2884 1811 2896
rect 1885 2884 1891 2896
rect 1293 2724 1299 2756
rect 1629 2744 1635 2876
rect 1405 2704 1411 2716
rect 1229 2684 1235 2696
rect 1517 2684 1523 2736
rect 1773 2724 1779 2876
rect 1917 2844 1923 2856
rect 1789 2784 1795 2796
rect 1933 2724 1939 2836
rect 1965 2724 1971 2896
rect 1997 2884 2003 2936
rect 2013 2864 2019 2896
rect 2045 2784 2051 2936
rect 2061 2884 2067 2936
rect 2093 2884 2099 2896
rect 2093 2864 2099 2876
rect 2109 2864 2115 2896
rect 2077 2744 2083 2836
rect 2141 2804 2147 2936
rect 2253 2924 2259 2936
rect 2221 2784 2227 2796
rect 2180 2717 2195 2723
rect 2125 2684 2131 2716
rect 2157 2684 2163 2716
rect 1453 2677 1468 2683
rect 13 2544 19 2656
rect 93 2644 99 2656
rect 157 2544 163 2636
rect 253 2544 259 2556
rect 269 2544 275 2636
rect 285 2564 291 2616
rect 301 2564 307 2636
rect 349 2604 355 2636
rect 13 2264 19 2536
rect 125 2504 131 2516
rect 269 2503 275 2536
rect 365 2504 371 2576
rect 413 2564 419 2636
rect 445 2583 451 2636
rect 525 2584 531 2636
rect 445 2577 467 2583
rect 461 2563 467 2577
rect 461 2557 476 2563
rect 509 2544 515 2556
rect 541 2544 547 2676
rect 557 2564 563 2636
rect 653 2604 659 2636
rect 685 2584 691 2636
rect 637 2564 643 2576
rect 733 2563 739 2636
rect 733 2557 748 2563
rect 541 2524 547 2536
rect 260 2497 275 2503
rect 93 2264 99 2496
rect 157 2364 163 2436
rect 221 2344 227 2436
rect 269 2364 275 2436
rect 269 2324 275 2336
rect 317 2324 323 2496
rect 365 2484 371 2496
rect 333 2324 339 2436
rect 381 2324 387 2356
rect 429 2304 435 2436
rect 461 2324 467 2436
rect 509 2363 515 2516
rect 701 2504 707 2516
rect 589 2484 595 2496
rect 765 2463 771 2636
rect 797 2584 803 2596
rect 781 2564 787 2576
rect 813 2544 819 2616
rect 845 2544 851 2676
rect 909 2624 915 2656
rect 964 2637 972 2643
rect 845 2504 851 2536
rect 941 2524 947 2616
rect 989 2544 995 2636
rect 1005 2624 1011 2656
rect 989 2524 995 2536
rect 893 2504 899 2516
rect 749 2457 771 2463
rect 621 2364 627 2436
rect 493 2357 515 2363
rect 493 2344 499 2357
rect 493 2324 499 2336
rect 621 2324 627 2336
rect 509 2303 515 2316
rect 468 2297 515 2303
rect 413 2284 419 2296
rect 212 2277 236 2283
rect 548 2277 556 2283
rect 285 2264 291 2276
rect 637 2264 643 2456
rect 653 2404 659 2436
rect 669 2364 675 2436
rect 749 2324 755 2457
rect 765 2404 771 2436
rect 941 2424 947 2496
rect 989 2484 995 2496
rect 1037 2424 1043 2636
rect 1069 2584 1075 2656
rect 1149 2584 1155 2676
rect 1261 2584 1267 2616
rect 1277 2583 1283 2636
rect 1325 2604 1331 2676
rect 1277 2577 1299 2583
rect 1245 2564 1251 2576
rect 1293 2564 1299 2577
rect 1453 2563 1459 2677
rect 1700 2677 1724 2683
rect 2077 2664 2083 2676
rect 2173 2664 2179 2676
rect 2189 2664 2195 2717
rect 2253 2684 2259 2916
rect 2269 2804 2275 2957
rect 2397 2943 2403 2956
rect 2372 2937 2403 2943
rect 2429 2924 2435 2936
rect 2340 2917 2348 2923
rect 2301 2864 2307 2896
rect 2397 2864 2403 2896
rect 2301 2784 2307 2796
rect 2317 2724 2323 2756
rect 2333 2684 2339 2736
rect 2477 2724 2483 2836
rect 2461 2664 2467 2716
rect 2509 2704 2515 2936
rect 2525 2904 2531 2956
rect 2637 2944 2643 2996
rect 2733 2984 2739 2996
rect 2781 2943 2787 2956
rect 2797 2944 2803 2996
rect 3389 2984 3395 2996
rect 2829 2977 2860 2983
rect 2829 2964 2835 2977
rect 3005 2964 3011 2976
rect 3165 2964 3171 2976
rect 3837 2964 3843 2976
rect 3965 2964 3971 3083
rect 4061 2964 4067 3083
rect 3540 2957 3548 2963
rect 2845 2944 2851 2956
rect 2893 2944 2899 2956
rect 2925 2944 2931 2956
rect 2989 2944 2995 2956
rect 3293 2944 3299 2956
rect 3469 2944 3475 2956
rect 3581 2944 3587 2956
rect 2772 2937 2787 2943
rect 2557 2864 2563 2936
rect 3069 2904 3075 2936
rect 3213 2924 3219 2936
rect 3117 2904 3123 2916
rect 3261 2904 3267 2936
rect 3501 2904 3507 2916
rect 2692 2897 2700 2903
rect 2653 2804 2659 2836
rect 2717 2784 2723 2896
rect 2749 2784 2755 2896
rect 2813 2844 2819 2876
rect 2525 2724 2531 2736
rect 2797 2703 2803 2736
rect 2813 2724 2819 2836
rect 2893 2804 2899 2896
rect 3181 2884 3187 2896
rect 3021 2744 3027 2836
rect 2797 2697 2819 2703
rect 2813 2684 2819 2697
rect 3053 2684 3059 2876
rect 3133 2844 3139 2876
rect 3325 2744 3331 2876
rect 3341 2804 3347 2896
rect 3421 2824 3427 2896
rect 3133 2724 3139 2736
rect 2509 2664 2515 2676
rect 2436 2657 2444 2663
rect 1469 2644 1475 2656
rect 1565 2604 1571 2656
rect 1661 2644 1667 2656
rect 1476 2577 1507 2583
rect 1501 2564 1507 2577
rect 1444 2557 1459 2563
rect 1357 2544 1363 2556
rect 1485 2544 1491 2556
rect 1549 2544 1555 2556
rect 1629 2544 1635 2556
rect 1133 2504 1139 2536
rect 1373 2504 1379 2536
rect 1444 2497 1452 2503
rect 941 2384 947 2396
rect 765 2317 780 2323
rect 765 2303 771 2317
rect 852 2317 876 2323
rect 932 2317 956 2323
rect 708 2297 771 2303
rect 781 2284 787 2296
rect 733 2264 739 2276
rect 829 2264 835 2276
rect 13 2244 19 2256
rect 205 2244 211 2256
rect 13 2104 19 2196
rect 61 2184 67 2236
rect 141 2184 147 2236
rect 157 2184 163 2196
rect 125 2164 131 2176
rect 205 2164 211 2216
rect 253 2204 259 2236
rect 317 2164 323 2236
rect 381 2183 387 2236
rect 509 2204 515 2236
rect 589 2203 595 2236
rect 573 2197 595 2203
rect 365 2177 387 2183
rect 365 2163 371 2177
rect 356 2157 371 2163
rect 388 2157 444 2163
rect 109 2144 115 2156
rect 173 2124 179 2156
rect 221 2144 227 2156
rect 317 2124 323 2136
rect 525 2124 531 2136
rect 477 2104 483 2116
rect 573 2104 579 2197
rect 605 2164 611 2236
rect 637 2203 643 2256
rect 845 2244 851 2276
rect 621 2197 643 2203
rect 621 2104 627 2197
rect 669 2184 675 2236
rect 749 2164 755 2176
rect 653 2124 659 2136
rect 733 2124 739 2136
rect 637 2103 643 2116
rect 637 2097 684 2103
rect 397 2084 403 2096
rect 45 1924 51 1956
rect 77 1904 83 2036
rect 93 1924 99 1936
rect 141 1904 147 2036
rect 173 1924 179 1976
rect 189 1944 195 2036
rect 237 2004 243 2036
rect 253 1884 259 2076
rect 596 2057 604 2063
rect 269 1924 275 1936
rect 301 1884 307 1896
rect 381 1884 387 2056
rect 621 1964 627 2096
rect 765 2083 771 2236
rect 893 2164 899 2236
rect 925 2184 931 2256
rect 973 2244 979 2416
rect 989 2284 995 2356
rect 1053 2324 1059 2356
rect 1085 2324 1091 2496
rect 1181 2384 1187 2476
rect 1501 2364 1507 2536
rect 1661 2504 1667 2596
rect 1677 2544 1683 2656
rect 1725 2644 1731 2656
rect 1805 2604 1811 2656
rect 1741 2584 1747 2596
rect 1837 2584 1843 2656
rect 1917 2644 1923 2656
rect 1869 2624 1875 2636
rect 1533 2444 1539 2496
rect 1613 2444 1619 2456
rect 1565 2384 1571 2416
rect 1284 2337 1315 2343
rect 1028 2317 1036 2323
rect 1037 2244 1043 2276
rect 1133 2264 1139 2336
rect 1165 2284 1171 2336
rect 1309 2323 1315 2337
rect 1309 2317 1324 2323
rect 1117 2244 1123 2256
rect 829 2144 835 2156
rect 941 2144 947 2176
rect 957 2164 963 2236
rect 1053 2224 1059 2236
rect 1117 2184 1123 2196
rect 1165 2144 1171 2196
rect 1197 2144 1203 2276
rect 1245 2244 1251 2276
rect 1213 2184 1219 2236
rect 1261 2223 1267 2256
rect 1293 2244 1299 2316
rect 1325 2284 1331 2296
rect 1373 2284 1379 2356
rect 1405 2303 1411 2336
rect 1421 2324 1427 2336
rect 1453 2317 1500 2323
rect 1453 2303 1459 2317
rect 1405 2297 1459 2303
rect 1389 2264 1395 2276
rect 1469 2244 1475 2256
rect 1309 2224 1315 2236
rect 1261 2217 1283 2223
rect 1277 2184 1283 2217
rect 1236 2177 1244 2183
rect 1037 2137 1052 2143
rect 781 2124 787 2136
rect 1037 2124 1043 2137
rect 749 2077 771 2083
rect 637 1924 643 1976
rect 669 1924 675 1936
rect 749 1924 755 2077
rect 781 1984 787 2076
rect 797 1924 803 1936
rect 125 1864 131 1876
rect 253 1864 259 1876
rect 333 1864 339 1876
rect 157 1803 163 1836
rect 141 1797 163 1803
rect 141 1764 147 1797
rect 189 1784 195 1856
rect 365 1844 371 1856
rect 445 1844 451 1856
rect 237 1764 243 1836
rect 285 1804 291 1836
rect 301 1764 307 1776
rect 413 1764 419 1836
rect 461 1784 467 1916
rect 829 1884 835 1916
rect 893 1904 899 2116
rect 909 2084 915 2096
rect 1021 2084 1027 2096
rect 845 1884 851 1896
rect 957 1884 963 1936
rect 973 1924 979 2036
rect 1053 1884 1059 2116
rect 1117 2104 1123 2136
rect 1213 2124 1219 2136
rect 1261 2104 1267 2176
rect 1325 2144 1331 2196
rect 1357 2184 1363 2216
rect 1421 2164 1427 2236
rect 1565 2184 1571 2356
rect 1581 2284 1587 2436
rect 1709 2384 1715 2536
rect 1789 2504 1795 2536
rect 1748 2497 1756 2503
rect 1805 2503 1811 2536
rect 1837 2504 1843 2516
rect 1805 2497 1827 2503
rect 1821 2464 1827 2497
rect 1853 2464 1859 2596
rect 1869 2564 1875 2596
rect 1933 2544 1939 2576
rect 1901 2524 1907 2536
rect 1869 2484 1875 2496
rect 1853 2404 1859 2436
rect 1725 2324 1731 2396
rect 1837 2324 1843 2356
rect 1581 2164 1587 2276
rect 1629 2264 1635 2276
rect 1597 2244 1603 2256
rect 1661 2243 1667 2316
rect 1821 2277 1836 2283
rect 1677 2264 1683 2276
rect 1725 2244 1731 2256
rect 1789 2244 1795 2276
rect 1805 2264 1811 2276
rect 1821 2244 1827 2277
rect 1869 2244 1875 2256
rect 1661 2237 1683 2243
rect 1613 2164 1619 2176
rect 1645 2164 1651 2236
rect 1677 2184 1683 2237
rect 1885 2243 1891 2256
rect 1917 2243 1923 2256
rect 1885 2237 1923 2243
rect 1709 2224 1715 2236
rect 1901 2164 1907 2176
rect 1341 2124 1347 2136
rect 1309 2104 1315 2116
rect 1341 2104 1347 2116
rect 1373 2104 1379 2156
rect 1085 1924 1091 2036
rect 1101 1984 1107 2076
rect 1165 2044 1171 2096
rect 1245 2084 1251 2096
rect 1405 2084 1411 2156
rect 1469 2144 1475 2156
rect 1661 2144 1667 2156
rect 1789 2144 1795 2156
rect 1805 2144 1811 2156
rect 1885 2144 1891 2156
rect 1588 2137 1596 2143
rect 1421 2024 1427 2136
rect 1501 2104 1507 2136
rect 1709 2104 1715 2116
rect 1133 1884 1139 1916
rect 1165 1884 1171 1916
rect 1213 1884 1219 1996
rect 1357 1984 1363 2016
rect 1469 1984 1475 2096
rect 1693 2084 1699 2096
rect 1709 2064 1715 2096
rect 1741 2084 1747 2136
rect 1533 2004 1539 2036
rect 1725 2024 1731 2076
rect 1533 1924 1539 1936
rect 1613 1924 1619 1996
rect 1309 1884 1315 1916
rect 1645 1884 1651 1956
rect 1693 1904 1699 2016
rect 1757 1983 1763 2076
rect 1757 1977 1772 1983
rect 1789 1964 1795 2136
rect 1837 2084 1843 2096
rect 1805 1984 1811 2076
rect 1853 1984 1859 2096
rect 1933 2064 1939 2096
rect 1725 1924 1731 1936
rect 1693 1884 1699 1896
rect 1869 1884 1875 1916
rect 1924 1877 1932 1883
rect 637 1864 643 1876
rect 477 1764 483 1836
rect 557 1784 563 1856
rect 605 1803 611 1836
rect 589 1797 611 1803
rect 589 1764 595 1797
rect 653 1764 659 1836
rect 125 1744 131 1756
rect 269 1744 275 1756
rect 349 1744 355 1756
rect 13 1704 19 1736
rect 93 1584 99 1696
rect 77 1524 83 1556
rect 125 1524 131 1596
rect 125 1504 131 1516
rect 13 1384 19 1456
rect 77 1364 83 1376
rect 125 1344 131 1436
rect 189 1384 195 1456
rect 205 1424 211 1736
rect 221 1604 227 1636
rect 221 1464 227 1576
rect 269 1524 275 1676
rect 349 1604 355 1696
rect 429 1604 435 1756
rect 685 1743 691 1796
rect 701 1764 707 1776
rect 749 1764 755 1856
rect 765 1844 771 1856
rect 804 1837 812 1843
rect 669 1737 691 1743
rect 589 1604 595 1736
rect 669 1704 675 1737
rect 397 1584 403 1596
rect 461 1524 467 1556
rect 493 1524 499 1596
rect 685 1524 691 1636
rect 429 1484 435 1496
rect 317 1464 323 1476
rect 260 1457 268 1463
rect 205 1344 211 1396
rect 221 1384 227 1456
rect 381 1444 387 1456
rect 221 1344 227 1356
rect 253 1344 259 1356
rect 269 1343 275 1436
rect 445 1424 451 1436
rect 493 1423 499 1456
rect 525 1444 531 1456
rect 493 1417 515 1423
rect 301 1344 307 1416
rect 445 1384 451 1396
rect 509 1384 515 1417
rect 573 1384 579 1476
rect 637 1384 643 1516
rect 717 1484 723 1556
rect 749 1504 755 1636
rect 765 1484 771 1676
rect 781 1624 787 1816
rect 861 1783 867 1836
rect 893 1784 899 1856
rect 941 1784 947 1796
rect 845 1777 867 1783
rect 797 1644 803 1756
rect 845 1744 851 1777
rect 973 1783 979 1836
rect 1005 1824 1011 1876
rect 1021 1864 1027 1876
rect 1005 1784 1011 1816
rect 957 1777 979 1783
rect 957 1764 963 1777
rect 1053 1764 1059 1876
rect 1341 1864 1347 1876
rect 1293 1844 1299 1856
rect 973 1744 979 1756
rect 925 1724 931 1736
rect 813 1644 819 1696
rect 973 1604 979 1736
rect 781 1584 787 1596
rect 1021 1584 1027 1696
rect 1069 1603 1075 1836
rect 1149 1764 1155 1836
rect 1181 1804 1187 1836
rect 1165 1777 1212 1783
rect 1165 1764 1171 1777
rect 1277 1764 1283 1776
rect 1325 1764 1331 1836
rect 1341 1784 1347 1856
rect 1373 1844 1379 1856
rect 1453 1844 1459 1856
rect 1485 1844 1491 1856
rect 1565 1844 1571 1876
rect 1421 1784 1427 1796
rect 1085 1664 1091 1756
rect 1341 1744 1347 1756
rect 1373 1744 1379 1756
rect 1485 1744 1491 1756
rect 1501 1744 1507 1836
rect 1597 1784 1603 1856
rect 1620 1837 1628 1843
rect 1677 1804 1683 1856
rect 1725 1844 1731 1876
rect 1901 1863 1907 1876
rect 1901 1857 1932 1863
rect 1757 1844 1763 1856
rect 1789 1844 1795 1856
rect 1620 1757 1628 1763
rect 1069 1597 1091 1603
rect 1005 1524 1011 1536
rect 1085 1524 1091 1597
rect 813 1504 819 1516
rect 845 1484 851 1496
rect 1037 1484 1043 1496
rect 1101 1484 1107 1696
rect 1133 1684 1139 1736
rect 1325 1724 1331 1736
rect 1405 1724 1411 1736
rect 1293 1704 1299 1716
rect 1453 1704 1459 1716
rect 1533 1704 1539 1756
rect 1581 1744 1587 1756
rect 1725 1744 1731 1836
rect 1821 1784 1827 1856
rect 1853 1764 1859 1816
rect 1869 1804 1875 1836
rect 1949 1824 1955 2636
rect 1997 2623 2003 2656
rect 1988 2617 2003 2623
rect 2013 2584 2019 2656
rect 2109 2644 2115 2656
rect 2029 2624 2035 2636
rect 2237 2624 2243 2656
rect 2125 2584 2131 2616
rect 2157 2584 2163 2596
rect 2253 2584 2259 2656
rect 2397 2644 2403 2656
rect 2445 2564 2451 2616
rect 2004 2557 2019 2563
rect 2013 2544 2019 2557
rect 2093 2524 2099 2536
rect 2109 2524 2115 2536
rect 2189 2524 2195 2536
rect 1997 2504 2003 2516
rect 1965 2464 1971 2496
rect 2061 2484 2067 2496
rect 1981 2324 1987 2436
rect 2141 2404 2147 2496
rect 2157 2484 2163 2496
rect 2205 2404 2211 2536
rect 2285 2524 2291 2536
rect 2301 2504 2307 2556
rect 2420 2537 2444 2543
rect 2237 2384 2243 2396
rect 2045 2324 2051 2336
rect 1965 2184 1971 2236
rect 1981 2144 1987 2296
rect 1997 2184 2003 2316
rect 2045 2284 2051 2296
rect 2077 2284 2083 2376
rect 2333 2364 2339 2536
rect 2461 2504 2467 2636
rect 2141 2324 2147 2336
rect 2221 2324 2227 2336
rect 2269 2324 2275 2356
rect 2413 2344 2419 2476
rect 2461 2384 2467 2496
rect 2445 2317 2460 2323
rect 2125 2284 2131 2316
rect 2349 2284 2355 2316
rect 2445 2284 2451 2317
rect 2477 2303 2483 2636
rect 2557 2624 2563 2676
rect 2628 2657 2636 2663
rect 2692 2657 2700 2663
rect 2772 2657 2828 2663
rect 2637 2604 2643 2636
rect 2877 2584 2883 2676
rect 2893 2584 2899 2636
rect 2941 2624 2947 2656
rect 2957 2643 2963 2656
rect 2957 2637 2979 2643
rect 2973 2624 2979 2637
rect 3053 2624 3059 2656
rect 2925 2584 2931 2596
rect 2788 2577 2796 2583
rect 2765 2564 2771 2576
rect 2532 2557 2556 2563
rect 2493 2524 2499 2536
rect 2541 2524 2547 2536
rect 2605 2523 2611 2556
rect 2621 2524 2627 2556
rect 2765 2524 2771 2556
rect 2941 2544 2947 2556
rect 2957 2544 2963 2616
rect 2980 2577 2988 2583
rect 2973 2557 3020 2563
rect 2973 2544 2979 2557
rect 3053 2544 3059 2556
rect 2996 2537 3004 2543
rect 2596 2517 2611 2523
rect 2685 2504 2691 2516
rect 2829 2504 2835 2516
rect 2468 2297 2483 2303
rect 2196 2277 2204 2283
rect 2029 2264 2035 2276
rect 2141 2264 2147 2276
rect 2125 2183 2131 2236
rect 2237 2204 2243 2236
rect 2301 2224 2307 2276
rect 2365 2184 2371 2196
rect 2125 2177 2275 2183
rect 2269 2164 2275 2177
rect 2397 2164 2403 2236
rect 2445 2164 2451 2236
rect 2477 2164 2483 2236
rect 2493 2224 2499 2476
rect 2605 2384 2611 2416
rect 2605 2324 2611 2376
rect 2653 2324 2659 2476
rect 2717 2444 2723 2456
rect 2765 2384 2771 2496
rect 2781 2324 2787 2336
rect 2548 2317 2556 2323
rect 2564 2297 2691 2303
rect 2685 2284 2691 2297
rect 2509 2264 2515 2276
rect 2557 2244 2563 2276
rect 2653 2244 2659 2276
rect 2541 2164 2547 2196
rect 2605 2184 2611 2216
rect 2621 2164 2627 2236
rect 2701 2224 2707 2316
rect 2749 2283 2755 2316
rect 2829 2284 2835 2376
rect 2861 2344 2867 2496
rect 2861 2324 2867 2336
rect 2877 2284 2883 2496
rect 2909 2464 2915 2536
rect 3037 2504 3043 2536
rect 2989 2464 2995 2496
rect 3069 2464 3075 2696
rect 3133 2664 3139 2676
rect 3133 2644 3139 2656
rect 3085 2544 3091 2596
rect 3101 2584 3107 2596
rect 3149 2564 3155 2696
rect 3325 2683 3331 2716
rect 3501 2684 3507 2856
rect 3517 2724 3523 2836
rect 3581 2724 3587 2936
rect 3661 2924 3667 2936
rect 3677 2924 3683 2936
rect 3709 2904 3715 2916
rect 3741 2824 3747 2916
rect 3949 2864 3955 2956
rect 3965 2904 3971 2956
rect 3677 2724 3683 2736
rect 3773 2724 3779 2756
rect 3556 2717 3564 2723
rect 3821 2704 3827 2836
rect 3629 2684 3635 2696
rect 3885 2684 3891 2776
rect 3933 2724 3939 2816
rect 4061 2803 4067 2956
rect 4141 2944 4147 2956
rect 4157 2904 4163 2956
rect 4077 2884 4083 2896
rect 4061 2797 4083 2803
rect 4045 2724 4051 2756
rect 4077 2684 4083 2797
rect 4093 2784 4099 2836
rect 4205 2804 4211 2836
rect 4125 2784 4131 2796
rect 4109 2724 4115 2736
rect 3325 2677 3363 2683
rect 3277 2644 3283 2676
rect 3357 2664 3363 2677
rect 3165 2624 3171 2636
rect 3325 2623 3331 2656
rect 3309 2617 3331 2623
rect 3165 2544 3171 2596
rect 3261 2584 3267 2596
rect 3309 2544 3315 2617
rect 3437 2604 3443 2636
rect 3396 2557 3420 2563
rect 3469 2563 3475 2616
rect 3501 2584 3507 2596
rect 3533 2584 3539 2596
rect 3549 2564 3555 2636
rect 3693 2584 3699 2676
rect 3805 2643 3811 2676
rect 3981 2664 3987 2676
rect 3805 2637 3827 2643
rect 3821 2584 3827 2637
rect 3869 2564 3875 2636
rect 3885 2584 3891 2596
rect 3901 2584 3907 2636
rect 3917 2584 3923 2596
rect 3981 2584 3987 2616
rect 4189 2604 4195 2716
rect 4157 2584 4163 2596
rect 4221 2584 4227 2676
rect 3965 2564 3971 2576
rect 4045 2564 4051 2576
rect 3453 2557 3475 2563
rect 3348 2537 3356 2543
rect 3389 2537 3420 2543
rect 3188 2437 3196 2443
rect 2909 2384 2915 2416
rect 3005 2337 3020 2343
rect 2941 2324 2947 2336
rect 2973 2303 2979 2336
rect 2989 2324 2995 2336
rect 3005 2303 3011 2337
rect 3085 2324 3091 2356
rect 2973 2297 3011 2303
rect 3021 2284 3027 2316
rect 3117 2303 3123 2316
rect 3092 2297 3123 2303
rect 2749 2277 2787 2283
rect 2781 2264 2787 2277
rect 2813 2264 2819 2276
rect 3021 2264 3027 2276
rect 3069 2264 3075 2276
rect 2749 2244 2755 2256
rect 2733 2164 2739 2236
rect 2845 2184 2851 2216
rect 2909 2164 2915 2196
rect 3085 2184 3091 2236
rect 3101 2184 3107 2236
rect 3037 2164 3043 2176
rect 3053 2164 3059 2176
rect 2516 2157 2524 2163
rect 1965 1904 1971 2136
rect 2029 2124 2035 2136
rect 2132 2117 2140 2123
rect 1997 2064 2003 2076
rect 2013 2064 2019 2096
rect 2029 2003 2035 2116
rect 2061 2024 2067 2096
rect 2029 1997 2051 2003
rect 2013 1944 2019 1996
rect 1981 1904 1987 1916
rect 1997 1883 2003 1896
rect 2045 1884 2051 1997
rect 2077 1984 2083 2056
rect 2109 2024 2115 2096
rect 2157 2004 2163 2156
rect 2237 2104 2243 2156
rect 2493 2144 2499 2156
rect 2765 2144 2771 2156
rect 2333 2124 2339 2136
rect 2381 2124 2387 2136
rect 1988 1877 2003 1883
rect 1997 1824 2003 1836
rect 1885 1744 1891 1756
rect 1901 1744 1907 1796
rect 2045 1764 2051 1856
rect 2077 1804 2083 1956
rect 2109 1924 2115 1996
rect 2148 1957 2156 1963
rect 2093 1883 2099 1896
rect 2173 1884 2179 2036
rect 2253 1924 2259 1956
rect 2093 1877 2163 1883
rect 2109 1784 2115 1856
rect 2141 1844 2147 1856
rect 2157 1844 2163 1877
rect 2125 1744 2131 1816
rect 1789 1704 1795 1716
rect 1165 1584 1171 1676
rect 1197 1624 1203 1636
rect 1373 1584 1379 1696
rect 1613 1684 1619 1696
rect 1133 1524 1139 1556
rect 1165 1484 1171 1576
rect 1565 1564 1571 1636
rect 1613 1524 1619 1576
rect 1364 1517 1372 1523
rect 1645 1523 1651 1636
rect 1693 1564 1699 1696
rect 1741 1624 1747 1696
rect 1821 1644 1827 1736
rect 1645 1517 1660 1523
rect 1213 1484 1219 1516
rect 1421 1504 1427 1516
rect 1453 1484 1459 1516
rect 1837 1484 1843 1636
rect 1853 1524 1859 1596
rect 1885 1584 1891 1616
rect 1869 1524 1875 1576
rect 1885 1503 1891 1556
rect 1901 1523 1907 1736
rect 2061 1724 2067 1736
rect 1933 1684 1939 1696
rect 1949 1684 1955 1696
rect 1901 1517 1923 1523
rect 1869 1497 1891 1503
rect 733 1464 739 1476
rect 877 1464 883 1476
rect 429 1364 435 1376
rect 365 1344 371 1356
rect 477 1344 483 1356
rect 269 1337 291 1343
rect 13 1184 19 1296
rect 93 1284 99 1296
rect 45 1144 51 1276
rect 221 1184 227 1296
rect 221 1164 227 1176
rect 285 1124 291 1337
rect 29 984 35 1056
rect 189 1044 195 1056
rect 13 784 19 936
rect 45 904 51 1036
rect 93 984 99 1036
rect 125 984 131 1036
rect 205 984 211 1056
rect 189 964 195 976
rect 253 964 259 1036
rect 285 1024 291 1036
rect 301 1003 307 1296
rect 404 1137 412 1143
rect 285 997 307 1003
rect 61 924 67 936
rect 45 724 51 736
rect 109 684 115 836
rect 125 744 131 876
rect 285 824 291 997
rect 349 964 355 1036
rect 413 984 419 1116
rect 429 1104 435 1276
rect 557 1204 563 1356
rect 605 1264 611 1356
rect 653 1324 659 1336
rect 660 1297 668 1303
rect 461 1124 467 1136
rect 493 1084 499 1196
rect 621 1164 627 1296
rect 589 1124 595 1136
rect 509 1104 515 1116
rect 637 1104 643 1116
rect 541 1084 547 1096
rect 669 1084 675 1256
rect 557 1064 563 1076
rect 621 1064 627 1076
rect 493 964 499 1036
rect 589 1004 595 1036
rect 685 1004 691 1436
rect 797 1384 803 1456
rect 797 1344 803 1356
rect 877 1344 883 1436
rect 893 1424 899 1436
rect 957 1364 963 1456
rect 989 1384 995 1456
rect 1165 1444 1171 1456
rect 1085 1363 1091 1436
rect 1245 1404 1251 1476
rect 1261 1464 1267 1476
rect 1188 1377 1235 1383
rect 1229 1364 1235 1377
rect 1085 1357 1116 1363
rect 1053 1344 1059 1356
rect 1236 1337 1276 1343
rect 701 1324 707 1336
rect 829 1324 835 1336
rect 1101 1324 1107 1336
rect 1293 1324 1299 1476
rect 1309 1444 1315 1456
rect 1357 1423 1363 1456
rect 1357 1417 1372 1423
rect 1437 1384 1443 1416
rect 1453 1384 1459 1476
rect 1501 1464 1507 1476
rect 1709 1464 1715 1476
rect 1469 1444 1475 1456
rect 1549 1424 1555 1456
rect 1773 1443 1779 1456
rect 1773 1437 1795 1443
rect 1549 1384 1555 1396
rect 1421 1363 1427 1376
rect 1597 1364 1603 1416
rect 1421 1357 1468 1363
rect 1421 1337 1436 1343
rect 932 1297 940 1303
rect 797 1284 803 1296
rect 781 1203 787 1236
rect 845 1224 851 1296
rect 781 1197 803 1203
rect 772 1177 780 1183
rect 765 1124 771 1136
rect 797 1084 803 1197
rect 925 1184 931 1236
rect 845 1124 851 1176
rect 861 1104 867 1116
rect 893 1084 899 1136
rect 941 1104 947 1276
rect 973 1244 979 1296
rect 989 1184 995 1236
rect 973 1124 979 1136
rect 1053 1124 1059 1276
rect 1181 1223 1187 1296
rect 1165 1217 1187 1223
rect 1165 1184 1171 1217
rect 1213 1084 1219 1316
rect 1293 1284 1299 1296
rect 797 1044 803 1056
rect 909 1044 915 1056
rect 509 964 515 976
rect 589 964 595 976
rect 621 964 627 996
rect 653 964 659 976
rect 429 944 435 956
rect 685 944 691 956
rect 765 944 771 1036
rect 861 1024 867 1036
rect 813 944 819 996
rect 877 984 883 996
rect 829 944 835 976
rect 893 964 899 996
rect 957 984 963 1036
rect 909 964 915 976
rect 973 944 979 1016
rect 1005 1004 1011 1056
rect 1037 984 1043 996
rect 989 944 995 976
rect 1069 944 1075 956
rect 1085 944 1091 1056
rect 1149 984 1155 1056
rect 1197 984 1203 1056
rect 1133 944 1139 956
rect 1213 944 1219 1056
rect 1229 1024 1235 1276
rect 1309 1263 1315 1296
rect 1293 1257 1315 1263
rect 1293 1184 1299 1257
rect 1341 1244 1347 1336
rect 1357 1304 1363 1336
rect 1373 1304 1379 1316
rect 1245 1104 1251 1116
rect 1405 1064 1411 1116
rect 1261 1024 1267 1056
rect 1421 1024 1427 1337
rect 1492 1337 1500 1343
rect 1613 1303 1619 1436
rect 1645 1404 1651 1436
rect 1661 1424 1667 1436
rect 1725 1424 1731 1436
rect 1757 1364 1763 1416
rect 1789 1384 1795 1437
rect 1757 1304 1763 1336
rect 1773 1304 1779 1376
rect 1837 1364 1843 1436
rect 1869 1384 1875 1497
rect 1901 1484 1907 1496
rect 1917 1484 1923 1517
rect 1949 1484 1955 1516
rect 2029 1504 2035 1696
rect 2077 1624 2083 1736
rect 2109 1704 2115 1716
rect 2045 1484 2051 1516
rect 2077 1484 2083 1596
rect 2093 1524 2099 1556
rect 2125 1484 2131 1696
rect 2157 1664 2163 1696
rect 2029 1444 2035 1476
rect 1997 1364 2003 1436
rect 2020 1357 2028 1363
rect 1885 1344 1891 1356
rect 2045 1344 2051 1436
rect 2077 1404 2083 1476
rect 2125 1384 2131 1436
rect 2141 1384 2147 1636
rect 2173 1524 2179 1596
rect 2189 1564 2195 1836
rect 2205 1784 2211 1916
rect 2269 1884 2275 2116
rect 2333 2104 2339 2116
rect 2317 1964 2323 2036
rect 2413 2004 2419 2036
rect 2285 1937 2323 1943
rect 2221 1844 2227 1876
rect 2285 1844 2291 1937
rect 2301 1864 2307 1916
rect 2317 1903 2323 1937
rect 2349 1924 2355 1956
rect 2397 1924 2403 1956
rect 2429 1924 2435 2036
rect 2317 1897 2355 1903
rect 2349 1884 2355 1897
rect 2445 1884 2451 2036
rect 2461 2004 2467 2036
rect 2525 1964 2531 2096
rect 2573 2064 2579 2136
rect 2685 2104 2691 2136
rect 2733 2123 2739 2136
rect 2893 2124 2899 2136
rect 2733 2117 2764 2123
rect 2605 2084 2611 2096
rect 2637 1944 2643 2036
rect 2653 2024 2659 2036
rect 2749 2004 2755 2036
rect 2669 1984 2675 1996
rect 2845 1964 2851 2096
rect 2861 2084 2867 2096
rect 2909 1964 2915 2076
rect 2941 2064 2947 2156
rect 3117 2144 3123 2276
rect 3181 2264 3187 2316
rect 3213 2304 3219 2536
rect 3245 2464 3251 2496
rect 3293 2423 3299 2536
rect 3389 2504 3395 2537
rect 3453 2543 3459 2557
rect 3613 2557 3683 2563
rect 3613 2544 3619 2557
rect 3677 2544 3683 2557
rect 3444 2537 3459 2543
rect 3508 2537 3516 2543
rect 3556 2537 3564 2543
rect 3645 2504 3651 2536
rect 3341 2464 3347 2496
rect 3437 2484 3443 2496
rect 3277 2417 3299 2423
rect 3277 2403 3283 2417
rect 3245 2397 3283 2403
rect 3357 2397 3411 2403
rect 3229 2304 3235 2396
rect 3245 2384 3251 2397
rect 3261 2324 3267 2356
rect 3357 2324 3363 2397
rect 3405 2384 3411 2397
rect 3421 2323 3427 2476
rect 3485 2404 3491 2496
rect 3437 2324 3443 2376
rect 3396 2317 3427 2323
rect 3309 2284 3315 2296
rect 3229 2244 3235 2276
rect 3149 2164 3155 2236
rect 3277 2224 3283 2256
rect 3437 2244 3443 2316
rect 3517 2303 3523 2496
rect 3565 2397 3619 2403
rect 3565 2324 3571 2397
rect 3613 2384 3619 2397
rect 3645 2384 3651 2396
rect 3501 2297 3523 2303
rect 3501 2264 3507 2297
rect 3517 2244 3523 2276
rect 3565 2264 3571 2276
rect 3300 2237 3308 2243
rect 3373 2224 3379 2236
rect 3309 2164 3315 2216
rect 3469 2184 3475 2236
rect 3565 2184 3571 2256
rect 3597 2223 3603 2316
rect 3661 2283 3667 2536
rect 3789 2504 3795 2556
rect 4061 2544 4067 2556
rect 4189 2544 4195 2556
rect 3908 2537 3916 2543
rect 3853 2524 3859 2536
rect 3693 2484 3699 2496
rect 3725 2384 3731 2496
rect 3853 2444 3859 2516
rect 3933 2384 3939 2476
rect 3949 2364 3955 2436
rect 3981 2384 3987 2496
rect 4125 2424 4131 2536
rect 4173 2524 4179 2536
rect 4045 2384 4051 2416
rect 3677 2324 3683 2356
rect 4061 2324 4067 2336
rect 3805 2304 3811 2316
rect 3661 2277 3683 2283
rect 3581 2217 3603 2223
rect 3437 2164 3443 2176
rect 3565 2144 3571 2156
rect 3268 2137 3308 2143
rect 3165 2104 3171 2136
rect 3357 2104 3363 2136
rect 3581 2123 3587 2217
rect 3613 2164 3619 2236
rect 3629 2184 3635 2256
rect 3613 2144 3619 2156
rect 3572 2117 3587 2123
rect 3389 2104 3395 2116
rect 3629 2104 3635 2156
rect 3677 2104 3683 2277
rect 3709 2184 3715 2276
rect 3725 2224 3731 2276
rect 3773 2264 3779 2276
rect 3757 2183 3763 2236
rect 3821 2204 3827 2316
rect 3901 2303 3907 2316
rect 3876 2297 3907 2303
rect 3853 2224 3859 2276
rect 3901 2224 3907 2276
rect 4013 2264 4019 2316
rect 4141 2304 4147 2496
rect 4093 2284 4099 2296
rect 4141 2264 4147 2276
rect 4157 2264 4163 2276
rect 3965 2224 3971 2256
rect 4013 2204 4019 2256
rect 4253 2244 4259 2256
rect 3757 2177 3779 2183
rect 3773 2164 3779 2177
rect 3709 2144 3715 2156
rect 3757 2144 3763 2156
rect 3885 2144 3891 2156
rect 3725 2124 3731 2136
rect 3837 2104 3843 2116
rect 3933 2104 3939 2156
rect 4077 2104 4083 2236
rect 4125 2184 4131 2236
rect 4093 2144 4099 2176
rect 4141 2144 4147 2156
rect 4173 2144 4179 2156
rect 2980 2097 2988 2103
rect 3069 2097 3084 2103
rect 2589 1924 2595 1936
rect 2845 1924 2851 1936
rect 2532 1917 2540 1923
rect 2861 1903 2867 1936
rect 2909 1924 2915 1936
rect 2820 1897 2867 1903
rect 2893 1884 2899 1896
rect 2941 1884 2947 1936
rect 3021 1924 3027 1996
rect 3053 1944 3059 2076
rect 3069 1984 3075 2097
rect 3197 2024 3203 2096
rect 3581 2084 3587 2096
rect 3581 2064 3587 2076
rect 3757 2044 3763 2096
rect 3101 1984 3107 2016
rect 3117 1884 3123 1956
rect 3229 1924 3235 1936
rect 3341 1924 3347 2036
rect 3357 1984 3363 1996
rect 3181 1884 3187 1916
rect 3293 1904 3299 1916
rect 3341 1884 3347 1896
rect 3405 1884 3411 1956
rect 3421 1924 3427 2036
rect 3453 1964 3459 2036
rect 3837 1984 3843 2056
rect 3469 1924 3475 1956
rect 3821 1924 3827 1936
rect 3508 1917 3532 1923
rect 2660 1877 2684 1883
rect 2253 1784 2259 1836
rect 2317 1804 2323 1876
rect 2356 1857 2403 1863
rect 2397 1843 2403 1857
rect 2436 1857 2460 1863
rect 2477 1857 2563 1863
rect 2477 1843 2483 1857
rect 2397 1837 2483 1843
rect 2557 1843 2563 1857
rect 2557 1837 2572 1843
rect 2381 1804 2387 1836
rect 2397 1784 2403 1816
rect 2445 1784 2451 1796
rect 2429 1764 2435 1776
rect 2333 1757 2348 1763
rect 2221 1744 2227 1756
rect 2301 1743 2307 1756
rect 2333 1743 2339 1757
rect 2301 1737 2339 1743
rect 2349 1724 2355 1736
rect 2301 1704 2307 1716
rect 2205 1584 2211 1656
rect 2253 1484 2259 1556
rect 2349 1544 2355 1716
rect 2381 1704 2387 1756
rect 2413 1744 2419 1756
rect 2493 1744 2499 1756
rect 2541 1744 2547 1836
rect 2589 1764 2595 1876
rect 2813 1864 2819 1876
rect 2941 1857 2956 1863
rect 2637 1844 2643 1856
rect 2685 1784 2691 1856
rect 2765 1784 2771 1856
rect 2781 1784 2787 1856
rect 2829 1763 2835 1836
rect 2813 1757 2835 1763
rect 2797 1704 2803 1736
rect 2365 1624 2371 1636
rect 2381 1624 2387 1696
rect 2381 1524 2387 1616
rect 2461 1604 2467 1696
rect 2404 1537 2419 1543
rect 2317 1484 2323 1516
rect 2349 1484 2355 1516
rect 2413 1503 2419 1537
rect 2429 1524 2435 1596
rect 2525 1584 2531 1596
rect 2477 1524 2483 1536
rect 2557 1524 2563 1676
rect 2669 1604 2675 1656
rect 2717 1603 2723 1696
rect 2781 1683 2787 1696
rect 2813 1683 2819 1757
rect 2845 1743 2851 1776
rect 2845 1737 2860 1743
rect 2781 1677 2819 1683
rect 2829 1624 2835 1736
rect 2877 1704 2883 1836
rect 2941 1784 2947 1857
rect 3037 1844 3043 1856
rect 2717 1597 2739 1603
rect 2669 1584 2675 1596
rect 2733 1584 2739 1597
rect 2637 1537 2675 1543
rect 2637 1524 2643 1537
rect 2669 1523 2675 1537
rect 2797 1524 2803 1536
rect 2813 1524 2819 1616
rect 2669 1517 2684 1523
rect 2413 1497 2444 1503
rect 2605 1483 2611 1516
rect 2605 1477 2620 1483
rect 2173 1464 2179 1476
rect 2189 1444 2195 1456
rect 1908 1337 1916 1343
rect 1613 1297 1628 1303
rect 1437 1284 1443 1296
rect 1485 1284 1491 1296
rect 1453 1124 1459 1276
rect 1485 1084 1491 1256
rect 1533 1204 1539 1296
rect 1725 1284 1731 1296
rect 1588 1277 1596 1283
rect 1613 1224 1619 1236
rect 1533 1084 1539 1176
rect 1565 1124 1571 1216
rect 1613 1124 1619 1196
rect 1757 1184 1763 1296
rect 1853 1204 1859 1296
rect 1965 1204 1971 1336
rect 2061 1244 2067 1356
rect 2173 1344 2179 1376
rect 2221 1364 2227 1436
rect 2333 1384 2339 1396
rect 2269 1364 2275 1376
rect 2349 1364 2355 1376
rect 2365 1364 2371 1436
rect 2397 1363 2403 1416
rect 2413 1404 2419 1436
rect 2429 1424 2435 1476
rect 2445 1404 2451 1476
rect 2461 1384 2467 1416
rect 2477 1364 2483 1376
rect 2397 1357 2419 1363
rect 2125 1304 2131 1336
rect 2164 1297 2172 1303
rect 2141 1284 2147 1296
rect 1908 1157 1916 1163
rect 1693 1124 1699 1156
rect 1709 1124 1715 1136
rect 1933 1124 1939 1136
rect 1981 1124 1987 1236
rect 2205 1204 2211 1356
rect 2317 1304 2323 1316
rect 2397 1304 2403 1316
rect 2397 1284 2403 1296
rect 2157 1184 2163 1196
rect 1389 964 1395 996
rect 1453 984 1459 1076
rect 1613 1064 1619 1116
rect 1645 1084 1651 1116
rect 1981 1084 1987 1116
rect 2029 1084 2035 1156
rect 2077 1124 2083 1176
rect 2173 1124 2179 1136
rect 2221 1084 2227 1156
rect 2237 1144 2243 1236
rect 2365 1184 2371 1216
rect 2381 1164 2387 1236
rect 2413 1224 2419 1357
rect 2429 1344 2435 1356
rect 2477 1344 2483 1356
rect 2493 1304 2499 1436
rect 2541 1364 2547 1416
rect 2557 1384 2563 1476
rect 2573 1424 2579 1436
rect 2653 1384 2659 1496
rect 2765 1484 2771 1516
rect 2861 1484 2867 1676
rect 2909 1564 2915 1736
rect 2925 1684 2931 1736
rect 2957 1704 2963 1796
rect 3053 1784 3059 1796
rect 2973 1744 2979 1776
rect 3021 1764 3027 1776
rect 3069 1764 3075 1776
rect 3069 1704 3075 1736
rect 3005 1684 3011 1696
rect 2925 1584 2931 1616
rect 2989 1564 2995 1636
rect 2957 1504 2963 1516
rect 2845 1464 2851 1476
rect 2909 1464 2915 1496
rect 2756 1457 2771 1463
rect 2669 1384 2675 1396
rect 2445 1264 2451 1296
rect 2509 1264 2515 1356
rect 2525 1304 2531 1356
rect 2573 1344 2579 1376
rect 2621 1344 2627 1376
rect 2701 1344 2707 1356
rect 2541 1304 2547 1336
rect 2701 1304 2707 1336
rect 2612 1297 2620 1303
rect 2285 1144 2291 1156
rect 2301 1084 2307 1156
rect 2477 1124 2483 1136
rect 2525 1124 2531 1296
rect 2573 1184 2579 1296
rect 2653 1264 2659 1296
rect 2717 1244 2723 1456
rect 2765 1384 2771 1457
rect 2989 1444 2995 1456
rect 2749 1344 2755 1376
rect 2788 1357 2796 1363
rect 2765 1344 2771 1356
rect 2845 1344 2851 1396
rect 2877 1364 2883 1436
rect 3085 1424 3091 1856
rect 3117 1784 3123 1856
rect 3149 1803 3155 1836
rect 3261 1824 3267 1876
rect 3373 1864 3379 1876
rect 3412 1857 3427 1863
rect 3133 1797 3155 1803
rect 3133 1764 3139 1797
rect 3309 1784 3315 1796
rect 3204 1777 3212 1783
rect 3325 1764 3331 1836
rect 3389 1804 3395 1836
rect 3421 1784 3427 1857
rect 3501 1823 3507 1876
rect 3613 1844 3619 1856
rect 3501 1817 3523 1823
rect 3341 1744 3347 1756
rect 3197 1724 3203 1736
rect 3197 1704 3203 1716
rect 3245 1684 3251 1736
rect 3261 1724 3267 1736
rect 3284 1717 3292 1723
rect 3293 1684 3299 1696
rect 3149 1504 3155 1636
rect 3197 1584 3203 1676
rect 3213 1524 3219 1616
rect 3309 1564 3315 1716
rect 3341 1604 3347 1736
rect 3373 1684 3379 1696
rect 3357 1664 3363 1676
rect 3389 1664 3395 1756
rect 3469 1743 3475 1796
rect 3485 1764 3491 1776
rect 3469 1737 3491 1743
rect 3325 1583 3331 1596
rect 3325 1577 3356 1583
rect 3245 1504 3251 1516
rect 3309 1504 3315 1556
rect 3341 1504 3347 1516
rect 3133 1484 3139 1496
rect 3389 1484 3395 1556
rect 3485 1524 3491 1737
rect 3517 1624 3523 1817
rect 3533 1744 3539 1756
rect 3549 1723 3555 1836
rect 3581 1764 3587 1816
rect 3613 1784 3619 1796
rect 3645 1784 3651 1856
rect 3709 1784 3715 1916
rect 3741 1864 3747 1876
rect 3780 1857 3795 1863
rect 3789 1784 3795 1857
rect 3821 1784 3827 1836
rect 3837 1764 3843 1836
rect 3565 1744 3571 1756
rect 3645 1744 3651 1756
rect 3677 1724 3683 1756
rect 3853 1743 3859 2076
rect 3917 2024 3923 2096
rect 3933 2003 3939 2096
rect 3917 1997 3939 2003
rect 3917 1884 3923 1997
rect 4029 1944 4035 2036
rect 4093 2003 4099 2136
rect 4125 2104 4131 2116
rect 4093 1997 4115 2003
rect 3949 1924 3955 1936
rect 4077 1924 4083 1936
rect 3997 1884 4003 1916
rect 4109 1904 4115 1997
rect 4109 1884 4115 1896
rect 4077 1864 4083 1876
rect 4116 1857 4124 1863
rect 4157 1844 4163 1856
rect 3933 1784 3939 1836
rect 4013 1784 4019 1836
rect 4205 1784 4211 1836
rect 3981 1764 3987 1776
rect 4173 1764 4179 1776
rect 4116 1757 4124 1763
rect 4253 1744 4259 2036
rect 3844 1737 3859 1743
rect 3533 1717 3555 1723
rect 3533 1704 3539 1717
rect 3789 1684 3795 1696
rect 3533 1524 3539 1656
rect 3444 1497 3452 1503
rect 3469 1484 3475 1516
rect 3565 1504 3571 1676
rect 3700 1637 3708 1643
rect 3597 1624 3603 1636
rect 3645 1504 3651 1516
rect 3613 1484 3619 1496
rect 3661 1484 3667 1616
rect 3693 1544 3699 1596
rect 3693 1524 3699 1536
rect 3789 1524 3795 1656
rect 3821 1644 3827 1736
rect 3869 1704 3875 1736
rect 4061 1704 4067 1736
rect 3805 1584 3811 1616
rect 3837 1524 3843 1556
rect 3885 1504 3891 1516
rect 3252 1477 3260 1483
rect 3101 1444 3107 1456
rect 2941 1364 2947 1416
rect 2973 1364 2979 1376
rect 2916 1357 2924 1363
rect 3037 1344 3043 1376
rect 3069 1364 3075 1376
rect 3085 1344 3091 1356
rect 2781 1317 2867 1323
rect 2781 1304 2787 1317
rect 2365 1097 2403 1103
rect 2365 1083 2371 1097
rect 2356 1077 2371 1083
rect 1492 1057 1500 1063
rect 1405 964 1411 976
rect 1485 964 1491 976
rect 1549 964 1555 1016
rect 1645 984 1651 1016
rect 1661 984 1667 1056
rect 1693 983 1699 1036
rect 1741 1023 1747 1076
rect 1757 1043 1763 1056
rect 1789 1044 1795 1056
rect 1901 1044 1907 1076
rect 1757 1037 1779 1043
rect 1741 1017 1756 1023
rect 1757 984 1763 1016
rect 1693 977 1731 983
rect 1684 957 1708 963
rect 1725 963 1731 977
rect 1773 963 1779 1037
rect 1901 1023 1907 1036
rect 1933 1023 1939 1056
rect 2045 1044 2051 1076
rect 2381 1064 2387 1076
rect 2397 1064 2403 1097
rect 2413 1084 2419 1116
rect 2429 1104 2435 1116
rect 2461 1084 2467 1116
rect 2557 1084 2563 1096
rect 2605 1084 2611 1176
rect 2717 1124 2723 1196
rect 2685 1084 2691 1116
rect 2733 1104 2739 1236
rect 2813 1184 2819 1296
rect 2861 1283 2867 1317
rect 2925 1304 2931 1336
rect 3117 1304 3123 1376
rect 3197 1344 3203 1436
rect 3229 1364 3235 1436
rect 3261 1364 3267 1436
rect 3309 1404 3315 1476
rect 3341 1424 3347 1436
rect 3357 1403 3363 1476
rect 3380 1457 3395 1463
rect 3341 1397 3363 1403
rect 3341 1364 3347 1397
rect 3389 1384 3395 1457
rect 3373 1364 3379 1376
rect 3309 1344 3315 1356
rect 3373 1304 3379 1336
rect 2861 1277 2915 1283
rect 2909 1264 2915 1277
rect 2989 1244 2995 1256
rect 2733 1064 2739 1076
rect 2221 1057 2236 1063
rect 1901 1017 1923 1023
rect 1933 1017 1955 1023
rect 1917 984 1923 1017
rect 1949 983 1955 1017
rect 2109 984 2115 1056
rect 2125 1044 2131 1056
rect 2221 1003 2227 1057
rect 2596 1057 2604 1063
rect 2349 1043 2355 1056
rect 2205 997 2227 1003
rect 2333 1037 2355 1043
rect 2205 984 2211 997
rect 2333 984 2339 1037
rect 1949 977 2044 983
rect 2253 977 2307 983
rect 2253 964 2259 977
rect 1725 957 1763 963
rect 1773 957 1788 963
rect 756 917 764 923
rect 141 784 147 816
rect 189 724 195 756
rect 13 544 19 636
rect 125 584 131 656
rect 157 564 163 616
rect 173 564 179 636
rect 205 584 211 716
rect 253 664 259 716
rect 349 664 355 896
rect 717 884 723 896
rect 365 744 371 876
rect 365 704 371 716
rect 397 684 403 696
rect 365 664 371 676
rect 301 584 307 636
rect 349 604 355 656
rect 445 644 451 656
rect 333 564 339 576
rect 461 564 467 836
rect 477 704 483 836
rect 557 724 563 836
rect 525 624 531 636
rect 621 624 627 676
rect 573 584 579 616
rect 637 583 643 836
rect 829 804 835 936
rect 1309 924 1315 936
rect 861 904 867 916
rect 1021 904 1027 916
rect 653 724 659 736
rect 701 684 707 696
rect 765 664 771 716
rect 797 664 803 796
rect 845 724 851 836
rect 877 784 883 816
rect 925 744 931 836
rect 941 824 947 896
rect 836 697 844 703
rect 813 684 819 696
rect 957 684 963 736
rect 973 664 979 896
rect 1117 883 1123 916
rect 1133 904 1139 916
rect 1181 904 1187 916
rect 1165 883 1171 896
rect 1117 877 1171 883
rect 1037 737 1091 743
rect 1037 704 1043 737
rect 1085 724 1091 737
rect 1053 704 1059 716
rect 1101 664 1107 816
rect 1172 717 1180 723
rect 1149 684 1155 696
rect 1229 664 1235 756
rect 1245 704 1251 716
rect 1277 684 1283 836
rect 1309 664 1315 916
rect 1357 904 1363 956
rect 1437 944 1443 956
rect 1549 944 1555 956
rect 1613 944 1619 956
rect 1757 944 1763 957
rect 2301 963 2307 977
rect 2301 957 2323 963
rect 1821 943 1827 956
rect 2029 944 2035 956
rect 2141 944 2147 956
rect 1812 937 1827 943
rect 1988 937 1996 943
rect 1565 923 1571 936
rect 1524 917 1571 923
rect 1517 864 1523 896
rect 1540 857 1548 863
rect 1373 724 1379 836
rect 1325 684 1331 696
rect 1373 664 1379 696
rect 1405 684 1411 856
rect 1581 844 1587 856
rect 1421 804 1427 836
rect 1437 724 1443 836
rect 1581 784 1587 796
rect 1597 784 1603 896
rect 1645 864 1651 896
rect 1693 884 1699 936
rect 1901 924 1907 936
rect 2077 924 2083 936
rect 1972 917 1980 923
rect 2036 917 2051 923
rect 1725 884 1731 896
rect 1485 724 1491 736
rect 1645 724 1651 776
rect 1725 724 1731 876
rect 1773 824 1779 896
rect 1885 864 1891 896
rect 1437 697 1491 703
rect 1437 663 1443 697
rect 1485 684 1491 697
rect 1565 664 1571 716
rect 1757 684 1763 776
rect 1773 724 1779 736
rect 1805 684 1811 836
rect 1645 664 1651 676
rect 1396 657 1443 663
rect 685 624 691 656
rect 765 637 780 643
rect 637 577 659 583
rect 317 544 323 556
rect 493 544 499 556
rect 557 544 563 556
rect 637 544 643 556
rect 388 537 396 543
rect 45 504 51 536
rect 589 524 595 536
rect 77 344 83 436
rect 45 324 51 336
rect 93 284 99 516
rect 404 497 428 503
rect 125 404 131 496
rect 493 484 499 496
rect 637 484 643 496
rect 173 384 179 396
rect 109 324 115 336
rect 141 284 147 376
rect 157 284 163 356
rect 205 324 211 436
rect 189 284 195 316
rect 237 284 243 356
rect 253 344 259 416
rect 253 324 259 336
rect 13 184 19 276
rect 253 264 259 276
rect 317 264 323 456
rect 413 403 419 436
rect 397 397 419 403
rect 397 284 403 397
rect 413 344 419 356
rect 429 324 435 336
rect 461 324 467 456
rect 573 404 579 436
rect 589 324 595 336
rect 605 324 611 396
rect 653 344 659 577
rect 669 544 675 596
rect 717 583 723 636
rect 701 577 723 583
rect 701 564 707 577
rect 765 563 771 637
rect 781 564 787 616
rect 829 584 835 596
rect 909 584 915 656
rect 925 624 931 636
rect 861 564 867 576
rect 1005 564 1011 596
rect 749 557 771 563
rect 749 544 755 557
rect 845 544 851 556
rect 941 544 947 556
rect 717 504 723 536
rect 509 284 515 296
rect 765 284 771 436
rect 797 344 803 356
rect 813 324 819 336
rect 893 324 899 496
rect 989 444 995 556
rect 1037 484 1043 496
rect 1053 444 1059 656
rect 1373 644 1379 656
rect 1069 544 1075 556
rect 1117 544 1123 556
rect 1133 544 1139 636
rect 1165 624 1171 636
rect 1309 584 1315 616
rect 1341 544 1347 596
rect 1357 564 1363 636
rect 1373 584 1379 596
rect 1421 564 1427 636
rect 1469 544 1475 636
rect 1501 584 1507 596
rect 1597 584 1603 656
rect 1645 604 1651 656
rect 1661 644 1667 656
rect 1837 644 1843 656
rect 1485 544 1491 556
rect 1501 504 1507 556
rect 1581 544 1587 556
rect 1741 544 1747 596
rect 1789 544 1795 636
rect 1837 584 1843 596
rect 1869 563 1875 836
rect 1933 764 1939 896
rect 1997 784 2003 916
rect 2045 904 2051 917
rect 2125 904 2131 936
rect 2285 924 2291 956
rect 2317 944 2323 957
rect 2349 944 2355 956
rect 2381 944 2387 1056
rect 2445 983 2451 1036
rect 2445 977 2467 983
rect 2461 963 2467 977
rect 2573 964 2579 1056
rect 2653 1044 2659 1056
rect 2829 1004 2835 1056
rect 2605 964 2611 996
rect 2781 984 2787 996
rect 2845 983 2851 1216
rect 2861 1204 2867 1236
rect 3005 1223 3011 1296
rect 3005 1217 3027 1223
rect 2957 1104 2963 1116
rect 3005 1104 3011 1196
rect 2932 1077 3011 1083
rect 3005 1064 3011 1077
rect 2868 1057 2876 1063
rect 2957 1023 2963 1036
rect 2941 1017 2963 1023
rect 2941 1004 2947 1017
rect 2973 1004 2979 1056
rect 2957 984 2963 996
rect 2829 977 2851 983
rect 2733 964 2739 976
rect 2829 964 2835 977
rect 2909 964 2915 976
rect 2461 957 2483 963
rect 2477 944 2483 957
rect 2845 957 2860 963
rect 2669 944 2675 956
rect 2813 944 2819 956
rect 2845 944 2851 957
rect 2973 944 2979 976
rect 2989 944 2995 1036
rect 3005 984 3011 996
rect 3021 963 3027 1217
rect 3037 1084 3043 1276
rect 3165 1264 3171 1296
rect 3389 1283 3395 1296
rect 3316 1277 3395 1283
rect 3037 964 3043 976
rect 3005 957 3027 963
rect 2525 917 2604 923
rect 2189 904 2195 916
rect 2333 904 2339 916
rect 2429 904 2435 916
rect 2525 904 2531 917
rect 2173 884 2179 896
rect 1885 724 1891 736
rect 1933 724 1939 736
rect 1949 724 1955 736
rect 1901 684 1907 696
rect 1981 684 1987 696
rect 2093 684 2099 876
rect 2189 744 2195 896
rect 2109 724 2115 736
rect 2205 724 2211 736
rect 2132 717 2140 723
rect 2141 684 2147 696
rect 2269 683 2275 836
rect 2349 784 2355 836
rect 2381 804 2387 896
rect 2317 724 2323 756
rect 2365 724 2371 736
rect 2381 684 2387 716
rect 2244 677 2275 683
rect 1885 664 1891 676
rect 2029 664 2035 676
rect 2285 664 2291 676
rect 2333 664 2339 676
rect 1917 583 1923 616
rect 1892 577 1923 583
rect 1949 564 1955 596
rect 1981 564 1987 656
rect 1860 557 1875 563
rect 1821 544 1827 556
rect 1901 544 1907 556
rect 1549 504 1555 516
rect 1140 497 1164 503
rect 1069 464 1075 476
rect 1085 464 1091 496
rect 957 343 963 436
rect 957 337 979 343
rect 733 264 739 276
rect 861 264 867 316
rect 941 264 947 276
rect 685 257 700 263
rect 45 164 51 236
rect 77 104 83 236
rect 125 144 131 236
rect 205 184 211 236
rect 221 184 227 256
rect 173 164 179 176
rect 269 164 275 216
rect 333 184 339 256
rect 429 224 435 236
rect 525 204 531 256
rect 493 184 499 196
rect 420 177 451 183
rect 381 164 387 176
rect 445 164 451 177
rect 548 157 556 163
rect 157 104 163 156
rect 301 144 307 156
rect 429 144 435 156
rect 557 104 563 116
rect 589 -43 595 236
rect 685 184 691 257
rect 973 263 979 337
rect 989 284 995 436
rect 1197 404 1203 436
rect 1245 384 1251 496
rect 1437 484 1443 496
rect 1629 484 1635 536
rect 1853 524 1859 536
rect 1716 497 1740 503
rect 1357 384 1363 416
rect 1389 404 1395 476
rect 1453 384 1459 396
rect 1005 324 1011 336
rect 1037 284 1043 376
rect 1133 324 1139 336
rect 1229 324 1235 336
rect 1165 284 1171 316
rect 1293 284 1299 376
rect 1053 263 1059 276
rect 1373 264 1379 276
rect 1437 264 1443 316
rect 1469 264 1475 356
rect 1533 344 1539 476
rect 1661 404 1667 436
rect 1533 324 1539 336
rect 1485 304 1491 316
rect 1613 304 1619 316
rect 973 257 1059 263
rect 1236 257 1260 263
rect 925 243 931 256
rect 925 237 956 243
rect 621 164 627 176
rect 733 164 739 176
rect 637 144 643 156
rect 733 104 739 156
rect 829 124 835 236
rect 861 164 867 236
rect 1005 224 1011 236
rect 1085 224 1091 236
rect 1117 184 1123 256
rect 1149 163 1155 236
rect 1197 224 1203 236
rect 1341 184 1347 256
rect 1437 244 1443 256
rect 1373 184 1379 196
rect 1389 164 1395 216
rect 1149 157 1171 163
rect 877 144 883 156
rect 909 104 915 156
rect 941 144 947 156
rect 1101 144 1107 156
rect 1165 104 1171 157
rect 1268 157 1292 163
rect 1213 104 1219 156
rect 1364 137 1388 143
rect 1405 143 1411 236
rect 1517 223 1523 276
rect 1597 264 1603 296
rect 1645 284 1651 296
rect 1661 284 1667 336
rect 1677 304 1683 436
rect 1725 364 1731 396
rect 1789 384 1795 496
rect 1693 264 1699 316
rect 1853 284 1859 516
rect 1869 504 1875 516
rect 2045 504 2051 636
rect 2205 563 2211 636
rect 2196 557 2211 563
rect 2077 544 2083 556
rect 2157 544 2163 556
rect 2237 544 2243 656
rect 2269 644 2275 656
rect 2301 584 2307 616
rect 2285 564 2291 576
rect 2269 544 2275 556
rect 2349 544 2355 656
rect 2413 604 2419 716
rect 2429 703 2435 736
rect 2477 724 2483 736
rect 2525 724 2531 816
rect 2541 744 2547 836
rect 2557 744 2563 836
rect 2621 703 2627 736
rect 2637 724 2643 756
rect 2669 744 2675 876
rect 2749 804 2755 936
rect 2861 904 2867 936
rect 2893 844 2899 936
rect 2973 924 2979 936
rect 3005 883 3011 957
rect 3117 904 3123 1116
rect 3165 1084 3171 1176
rect 3181 1104 3187 1116
rect 3133 964 3139 1076
rect 3277 1064 3283 1076
rect 3293 1064 3299 1156
rect 3325 1123 3331 1236
rect 3357 1184 3363 1236
rect 3389 1184 3395 1236
rect 3405 1224 3411 1436
rect 3469 1424 3475 1476
rect 3485 1464 3491 1476
rect 3565 1443 3571 1476
rect 3661 1464 3667 1476
rect 3588 1457 3603 1463
rect 3565 1437 3587 1443
rect 3421 1184 3427 1336
rect 3437 1244 3443 1416
rect 3533 1404 3539 1436
rect 3549 1364 3555 1396
rect 3581 1384 3587 1437
rect 3597 1424 3603 1457
rect 3661 1384 3667 1416
rect 3725 1384 3731 1496
rect 3917 1484 3923 1496
rect 3981 1484 3987 1636
rect 4109 1604 4115 1736
rect 4141 1504 4147 1636
rect 4157 1604 4163 1636
rect 4189 1624 4195 1636
rect 4221 1584 4227 1696
rect 3933 1464 3939 1476
rect 4061 1464 4067 1476
rect 3677 1364 3683 1376
rect 3757 1364 3763 1456
rect 4029 1444 4035 1456
rect 3949 1384 3955 1416
rect 3581 1357 3635 1363
rect 3581 1344 3587 1357
rect 3629 1344 3635 1357
rect 3613 1324 3619 1336
rect 3869 1304 3875 1376
rect 4077 1364 4083 1436
rect 4109 1424 4115 1456
rect 4093 1364 4099 1376
rect 3965 1344 3971 1356
rect 4141 1343 4147 1476
rect 4221 1464 4227 1476
rect 4237 1344 4243 1436
rect 4125 1337 4147 1343
rect 3453 1284 3459 1296
rect 3581 1284 3587 1296
rect 3373 1124 3379 1156
rect 3485 1124 3491 1136
rect 3309 1117 3331 1123
rect 3309 1064 3315 1117
rect 3325 1084 3331 1096
rect 3405 1084 3411 1116
rect 3517 1084 3523 1216
rect 3533 1184 3539 1196
rect 3613 1124 3619 1156
rect 3565 1104 3571 1116
rect 3613 1084 3619 1116
rect 3645 1104 3651 1216
rect 3661 1184 3667 1296
rect 3917 1264 3923 1336
rect 3709 1124 3715 1236
rect 3757 1184 3763 1256
rect 3789 1184 3795 1236
rect 4013 1223 4019 1336
rect 4013 1217 4035 1223
rect 4029 1184 4035 1217
rect 3853 1124 3859 1156
rect 3901 1124 3907 1136
rect 3645 1084 3651 1096
rect 3700 1077 3708 1083
rect 3549 1064 3555 1076
rect 3252 1057 3260 1063
rect 3197 1023 3203 1056
rect 3213 1044 3219 1056
rect 3181 1017 3203 1023
rect 3149 944 3155 996
rect 3181 984 3187 1017
rect 3197 944 3203 956
rect 3229 904 3235 976
rect 3309 964 3315 1036
rect 3437 1004 3443 1036
rect 3469 1023 3475 1056
rect 3453 1017 3475 1023
rect 3453 984 3459 1017
rect 3661 1003 3667 1076
rect 3661 997 3683 1003
rect 3245 944 3251 956
rect 3357 944 3363 956
rect 3453 944 3459 956
rect 3469 944 3475 996
rect 3508 977 3571 983
rect 3565 964 3571 977
rect 3517 944 3523 956
rect 3629 944 3635 956
rect 3277 904 3283 936
rect 3645 924 3651 956
rect 3677 944 3683 997
rect 3725 984 3731 1036
rect 3741 1024 3747 1116
rect 3869 1084 3875 1096
rect 3917 1084 3923 1116
rect 3949 1084 3955 1136
rect 3965 1084 3971 1096
rect 4109 1084 4115 1236
rect 3853 1064 3859 1076
rect 4013 1064 4019 1076
rect 3773 1044 3779 1056
rect 3805 984 3811 1056
rect 4077 1044 4083 1056
rect 3837 984 3843 996
rect 3853 944 3859 956
rect 3869 944 3875 956
rect 3796 937 3804 943
rect 3604 917 3635 923
rect 3373 904 3379 916
rect 3005 877 3027 883
rect 2845 784 2851 796
rect 2909 764 2915 876
rect 3021 803 3027 877
rect 3181 864 3187 896
rect 3245 804 3251 836
rect 3309 824 3315 836
rect 3021 797 3043 803
rect 3037 784 3043 797
rect 3165 784 3171 796
rect 3245 784 3251 796
rect 2669 724 2675 736
rect 2877 704 2883 716
rect 2429 697 2515 703
rect 2621 697 2643 703
rect 2509 684 2515 697
rect 2637 683 2643 697
rect 2909 684 2915 756
rect 3229 724 3235 756
rect 3277 724 3283 736
rect 3405 724 3411 796
rect 2637 677 2675 683
rect 2557 664 2563 676
rect 2605 663 2611 676
rect 2669 664 2675 677
rect 2829 664 2835 676
rect 2941 664 2947 676
rect 2605 657 2652 663
rect 2381 584 2387 596
rect 2445 584 2451 616
rect 1965 344 1971 436
rect 1917 284 1923 296
rect 1533 224 1539 236
rect 1501 217 1523 223
rect 1501 184 1507 217
rect 1428 157 1452 163
rect 1405 137 1427 143
rect 1277 124 1283 136
rect 1252 117 1267 123
rect 1012 97 1020 103
rect 1261 103 1267 117
rect 1421 123 1427 137
rect 1469 123 1475 136
rect 1293 117 1363 123
rect 1421 117 1475 123
rect 1293 103 1299 117
rect 1261 97 1299 103
rect 1357 103 1363 117
rect 1517 104 1523 176
rect 1549 164 1555 196
rect 1581 184 1587 196
rect 1597 144 1603 236
rect 1629 164 1635 216
rect 1645 104 1651 196
rect 1757 184 1763 256
rect 1773 244 1779 256
rect 1853 244 1859 256
rect 1821 184 1827 236
rect 1885 224 1891 236
rect 1933 224 1939 256
rect 1885 184 1891 196
rect 1709 164 1715 176
rect 1837 164 1843 176
rect 1869 164 1875 176
rect 1901 164 1907 196
rect 1965 144 1971 256
rect 2029 164 2035 436
rect 2045 364 2051 496
rect 2077 304 2083 536
rect 2237 504 2243 536
rect 2125 484 2131 496
rect 2205 484 2211 496
rect 2093 284 2099 296
rect 2157 264 2163 376
rect 2173 304 2179 436
rect 2205 324 2211 336
rect 2221 324 2227 336
rect 2237 324 2243 496
rect 2269 304 2275 536
rect 2349 524 2355 536
rect 2333 424 2339 436
rect 2285 324 2291 416
rect 2349 264 2355 356
rect 2365 324 2371 396
rect 2429 264 2435 496
rect 2493 444 2499 636
rect 2525 564 2531 636
rect 2509 544 2515 556
rect 2589 544 2595 656
rect 2557 504 2563 516
rect 2605 504 2611 636
rect 2637 563 2643 636
rect 2733 604 2739 636
rect 2861 604 2867 656
rect 2957 643 2963 676
rect 3101 644 3107 676
rect 2941 637 2963 643
rect 2877 584 2883 616
rect 2893 584 2899 596
rect 2637 557 2668 563
rect 2685 524 2691 556
rect 2797 544 2803 556
rect 2813 544 2819 556
rect 2845 544 2851 576
rect 2685 504 2691 516
rect 2765 504 2771 516
rect 2877 504 2883 536
rect 2893 504 2899 516
rect 2557 337 2572 343
rect 2541 264 2547 336
rect 2557 324 2563 337
rect 2621 303 2627 396
rect 2637 324 2643 436
rect 2653 404 2659 436
rect 2941 404 2947 637
rect 2957 564 2963 576
rect 3005 544 3011 556
rect 3021 544 3027 616
rect 3085 584 3091 616
rect 3117 584 3123 716
rect 3149 684 3155 696
rect 3181 584 3187 656
rect 3197 624 3203 676
rect 3325 657 3340 663
rect 3117 564 3123 576
rect 3229 564 3235 636
rect 3261 623 3267 656
rect 3261 617 3283 623
rect 3277 584 3283 617
rect 3325 604 3331 657
rect 3357 643 3363 716
rect 3421 684 3427 876
rect 3437 744 3443 756
rect 3453 724 3459 736
rect 3469 684 3475 916
rect 3629 904 3635 917
rect 3693 904 3699 936
rect 3901 924 3907 1036
rect 3917 964 3923 1036
rect 3997 964 4003 976
rect 4109 964 4115 1036
rect 4125 1024 4131 1337
rect 4157 1324 4163 1336
rect 4141 1084 4147 1236
rect 4173 1084 4179 1236
rect 4253 1184 4259 1196
rect 4189 1084 4195 1156
rect 4189 1064 4195 1076
rect 4157 1044 4163 1056
rect 4173 1004 4179 1036
rect 4205 1004 4211 1036
rect 4237 984 4243 1056
rect 4157 964 4163 976
rect 4125 944 4131 956
rect 3917 924 3923 936
rect 4109 924 4115 936
rect 3501 884 3507 896
rect 3533 884 3539 896
rect 3549 884 3555 896
rect 3565 784 3571 816
rect 3501 724 3507 736
rect 3629 724 3635 876
rect 3645 784 3651 896
rect 3741 884 3747 896
rect 3661 784 3667 836
rect 3725 724 3731 876
rect 3629 704 3635 716
rect 3741 684 3747 716
rect 3789 684 3795 916
rect 3821 904 3827 916
rect 3901 784 3907 896
rect 3917 824 3923 896
rect 3965 784 3971 816
rect 4061 784 4067 916
rect 4077 844 4083 896
rect 4029 724 4035 776
rect 4109 724 4115 756
rect 4141 724 4147 836
rect 4221 784 4227 936
rect 3821 704 3827 716
rect 3828 677 3836 683
rect 3348 637 3363 643
rect 3373 624 3379 676
rect 3581 664 3587 676
rect 3773 664 3779 676
rect 3261 564 3267 576
rect 3309 544 3315 576
rect 2973 524 2979 536
rect 3053 504 3059 536
rect 3005 484 3011 496
rect 2845 384 2851 396
rect 2685 344 2691 356
rect 2733 324 2739 376
rect 2893 324 2899 336
rect 2941 324 2947 336
rect 2612 297 2627 303
rect 2861 284 2867 296
rect 3021 284 3027 496
rect 3101 384 3107 536
rect 3149 504 3155 536
rect 3117 484 3123 496
rect 3165 423 3171 536
rect 3277 464 3283 496
rect 3309 464 3315 516
rect 3325 504 3331 576
rect 3412 557 3420 563
rect 3357 544 3363 556
rect 3485 544 3491 556
rect 3405 524 3411 536
rect 3501 524 3507 636
rect 3533 544 3539 636
rect 3597 584 3603 616
rect 3629 584 3635 656
rect 3885 644 3891 656
rect 3572 557 3580 563
rect 3661 544 3667 556
rect 3709 544 3715 616
rect 3725 563 3731 636
rect 3725 557 3747 563
rect 3741 543 3747 557
rect 3789 544 3795 556
rect 3805 544 3811 636
rect 3917 584 3923 676
rect 3837 544 3843 556
rect 3885 544 3891 556
rect 3933 544 3939 636
rect 3949 584 3955 596
rect 3981 584 3987 656
rect 4029 604 4035 636
rect 4045 584 4051 656
rect 4141 584 4147 676
rect 3965 564 3971 576
rect 4125 544 4131 556
rect 3741 537 3756 543
rect 3501 504 3507 516
rect 3165 417 3187 423
rect 3181 384 3187 417
rect 3037 324 3043 336
rect 3069 284 3075 356
rect 3117 324 3123 336
rect 3172 317 3180 323
rect 3252 317 3260 323
rect 3085 284 3091 316
rect 3252 277 3260 283
rect 2173 244 2179 256
rect 2605 244 2611 276
rect 2653 264 2659 276
rect 2909 264 2915 276
rect 3133 264 3139 276
rect 3293 264 3299 276
rect 2724 257 2780 263
rect 2045 164 2051 176
rect 2125 164 2131 176
rect 2157 164 2163 176
rect 2253 164 2259 196
rect 2429 184 2435 216
rect 2509 144 2515 236
rect 1725 124 1731 136
rect 1917 104 1923 136
rect 1949 124 1955 136
rect 1357 97 1420 103
rect 2356 97 2364 103
rect 813 84 819 96
rect 1181 84 1187 96
rect 1245 84 1251 96
rect 1469 84 1475 96
rect 1773 84 1779 96
rect 1949 84 1955 96
rect 2477 84 2483 96
rect 2573 -37 2579 236
rect 2621 164 2627 236
rect 2685 204 2691 236
rect 2701 164 2707 176
rect 2733 163 2739 236
rect 2717 157 2739 163
rect 2717 144 2723 157
rect 2765 144 2771 216
rect 2829 204 2835 256
rect 2877 224 2883 236
rect 2941 224 2947 236
rect 2941 124 2947 156
rect 2916 117 2924 123
rect 2989 104 2995 236
rect 3005 164 3011 216
rect 3037 204 3043 236
rect 3101 203 3107 236
rect 3085 197 3107 203
rect 3005 124 3011 136
rect 3069 104 3075 136
rect 3085 104 3091 197
rect 3117 144 3123 196
rect 3133 144 3139 256
rect 3197 184 3203 256
rect 3213 204 3219 236
rect 3261 164 3267 176
rect 3245 143 3251 156
rect 3277 143 3283 236
rect 3309 184 3315 396
rect 3341 284 3347 316
rect 3357 284 3363 496
rect 3373 484 3379 496
rect 3389 324 3395 356
rect 3405 284 3411 356
rect 3517 284 3523 416
rect 3533 264 3539 476
rect 3549 344 3555 436
rect 3565 324 3571 516
rect 3629 504 3635 536
rect 3677 504 3683 536
rect 3709 524 3715 536
rect 3725 524 3731 536
rect 4109 524 4115 536
rect 3741 503 3747 516
rect 3757 504 3763 516
rect 3837 504 3843 516
rect 3853 504 3859 516
rect 3732 497 3747 503
rect 3613 404 3619 496
rect 3853 484 3859 496
rect 3741 444 3747 456
rect 3773 444 3779 456
rect 3693 324 3699 396
rect 3821 324 3827 336
rect 3588 317 3596 323
rect 3565 284 3571 316
rect 3725 284 3731 296
rect 3773 284 3779 316
rect 3805 304 3811 316
rect 3853 284 3859 296
rect 3677 264 3683 276
rect 3901 264 3907 516
rect 3965 484 3971 496
rect 4013 484 4019 496
rect 4189 424 4195 496
rect 4109 384 4115 416
rect 4221 324 4227 436
rect 4237 384 4243 396
rect 3972 317 3980 323
rect 4013 277 4083 283
rect 3933 264 3939 276
rect 4013 264 4019 277
rect 4077 264 4083 277
rect 3485 244 3491 256
rect 3357 164 3363 176
rect 3373 144 3379 236
rect 3389 184 3395 236
rect 3421 183 3427 236
rect 3533 224 3539 236
rect 3405 177 3427 183
rect 3245 137 3283 143
rect 3405 124 3411 177
rect 3549 164 3555 236
rect 3629 223 3635 256
rect 3629 217 3651 223
rect 3405 104 3411 116
rect 2756 97 2764 103
rect 3101 84 3107 96
rect 3421 64 3427 156
rect 3597 144 3603 196
rect 3645 184 3651 217
rect 3725 184 3731 236
rect 3741 224 3747 256
rect 3805 224 3811 236
rect 3773 184 3779 196
rect 3613 164 3619 176
rect 3757 164 3763 176
rect 3821 164 3827 236
rect 3885 184 3891 256
rect 4093 244 4099 316
rect 4221 264 4227 296
rect 3933 164 3939 216
rect 4013 184 4019 196
rect 4029 164 4035 196
rect 3860 157 3868 163
rect 3805 144 3811 156
rect 3837 144 3843 156
rect 4045 144 4051 236
rect 4189 224 4195 236
rect 4269 204 4275 2936
rect 4109 184 4115 196
rect 4125 164 4131 176
rect 4173 144 4179 156
rect 4189 144 4195 156
rect 3485 124 3491 136
rect 3677 124 3683 136
rect 4077 124 4083 136
rect 4013 104 4019 116
rect 4093 104 4099 116
rect 3556 97 3564 103
rect 4228 97 4236 103
rect 2557 -43 2579 -37
rect 2877 -43 2883 16
<< m3contact >>
rect 220 2976 228 2984
rect 428 2976 436 2984
rect 444 2976 452 2984
rect 508 2976 516 2984
rect 524 2976 532 2984
rect 12 2956 20 2964
rect 156 2956 164 2964
rect 380 2956 388 2964
rect 140 2936 148 2944
rect 220 2936 228 2944
rect 92 2896 100 2904
rect 124 2896 132 2904
rect 92 2736 100 2744
rect 156 2736 164 2744
rect 252 2896 260 2904
rect 412 2936 420 2944
rect 732 2976 740 2984
rect 860 2976 868 2984
rect 1708 2976 1716 2984
rect 1756 2976 1764 2984
rect 1996 2976 2004 2984
rect 604 2956 612 2964
rect 620 2956 628 2964
rect 700 2956 708 2964
rect 876 2956 884 2964
rect 972 2956 980 2964
rect 1100 2956 1108 2964
rect 1164 2956 1172 2964
rect 1388 2956 1396 2964
rect 1420 2956 1428 2964
rect 1436 2956 1444 2964
rect 1516 2956 1524 2964
rect 1596 2956 1604 2964
rect 1740 2956 1748 2964
rect 460 2936 468 2944
rect 524 2936 532 2944
rect 764 2936 772 2944
rect 844 2936 852 2944
rect 332 2896 340 2904
rect 124 2716 132 2724
rect 236 2696 244 2704
rect 332 2796 340 2804
rect 364 2796 372 2804
rect 284 2736 292 2744
rect 460 2916 468 2924
rect 492 2916 500 2924
rect 476 2896 484 2904
rect 764 2916 772 2924
rect 572 2896 580 2904
rect 652 2896 660 2904
rect 684 2876 692 2884
rect 508 2796 516 2804
rect 524 2796 532 2804
rect 492 2736 500 2744
rect 412 2716 420 2724
rect 380 2696 388 2704
rect 492 2696 500 2704
rect 76 2676 84 2684
rect 172 2676 180 2684
rect 252 2676 260 2684
rect 380 2676 388 2684
rect 652 2776 660 2784
rect 620 2736 628 2744
rect 588 2696 596 2704
rect 748 2736 756 2744
rect 716 2716 724 2724
rect 668 2696 676 2704
rect 700 2696 708 2704
rect 908 2896 916 2904
rect 1772 2956 1780 2964
rect 1836 2956 1844 2964
rect 2012 2956 2020 2964
rect 2524 2996 2532 3004
rect 2636 2996 2644 3004
rect 2732 2996 2740 3004
rect 2796 2996 2804 3004
rect 3388 2996 3396 3004
rect 2124 2956 2132 2964
rect 2156 2956 2164 2964
rect 2220 2956 2228 2964
rect 1148 2936 1156 2944
rect 1516 2936 1524 2944
rect 1580 2936 1588 2944
rect 1692 2936 1700 2944
rect 972 2896 980 2904
rect 1004 2896 1012 2904
rect 924 2796 932 2804
rect 956 2796 964 2804
rect 844 2756 852 2764
rect 764 2716 772 2724
rect 796 2696 804 2704
rect 876 2696 884 2704
rect 956 2716 964 2724
rect 1116 2896 1124 2904
rect 1468 2896 1476 2904
rect 1052 2876 1060 2884
rect 1036 2856 1044 2864
rect 1020 2796 1028 2804
rect 1020 2736 1028 2744
rect 1196 2836 1204 2844
rect 1180 2796 1188 2804
rect 1100 2736 1108 2744
rect 1276 2856 1284 2864
rect 1228 2796 1236 2804
rect 1388 2836 1396 2844
rect 1340 2816 1348 2824
rect 1420 2816 1428 2824
rect 1548 2876 1556 2884
rect 1532 2836 1540 2844
rect 1676 2916 1684 2924
rect 1612 2876 1620 2884
rect 1628 2876 1636 2884
rect 1804 2876 1812 2884
rect 1884 2876 1892 2884
rect 1596 2796 1604 2804
rect 1468 2776 1476 2784
rect 1292 2756 1300 2764
rect 1452 2756 1460 2764
rect 1516 2736 1524 2744
rect 1708 2736 1716 2744
rect 1356 2716 1364 2724
rect 1484 2716 1492 2724
rect 1004 2696 1012 2704
rect 1228 2696 1236 2704
rect 1260 2696 1268 2704
rect 1404 2696 1412 2704
rect 1916 2836 1924 2844
rect 1788 2796 1796 2804
rect 1996 2876 2004 2884
rect 2012 2856 2020 2864
rect 2060 2876 2068 2884
rect 2092 2876 2100 2884
rect 2092 2856 2100 2864
rect 2108 2856 2116 2864
rect 2044 2776 2052 2784
rect 2252 2916 2260 2924
rect 2140 2796 2148 2804
rect 2220 2796 2228 2804
rect 2092 2776 2100 2784
rect 2076 2736 2084 2744
rect 1532 2716 1540 2724
rect 1964 2716 1972 2724
rect 2156 2716 2164 2724
rect 540 2676 548 2684
rect 828 2676 836 2684
rect 924 2676 932 2684
rect 1244 2676 1252 2684
rect 1436 2676 1444 2684
rect 12 2656 20 2664
rect 172 2656 180 2664
rect 524 2656 532 2664
rect 44 2636 52 2644
rect 92 2636 100 2644
rect 524 2636 532 2644
rect 76 2576 84 2584
rect 172 2556 180 2564
rect 284 2616 292 2624
rect 348 2596 356 2604
rect 364 2576 372 2584
rect 396 2576 404 2584
rect 284 2556 292 2564
rect 300 2556 308 2564
rect 156 2536 164 2544
rect 252 2536 260 2544
rect 268 2536 276 2544
rect 348 2536 356 2544
rect 124 2516 132 2524
rect 44 2496 52 2504
rect 92 2496 100 2504
rect 444 2556 452 2564
rect 508 2556 516 2564
rect 636 2656 644 2664
rect 764 2636 772 2644
rect 652 2596 660 2604
rect 636 2576 644 2584
rect 684 2576 692 2584
rect 556 2556 564 2564
rect 668 2556 676 2564
rect 732 2536 740 2544
rect 508 2516 516 2524
rect 540 2516 548 2524
rect 700 2516 708 2524
rect 316 2496 324 2504
rect 396 2496 404 2504
rect 492 2496 500 2504
rect 76 2316 84 2324
rect 156 2356 164 2364
rect 268 2356 276 2364
rect 220 2336 228 2344
rect 268 2336 276 2344
rect 364 2476 372 2484
rect 380 2356 388 2364
rect 156 2316 164 2324
rect 316 2316 324 2324
rect 332 2316 340 2324
rect 364 2316 372 2324
rect 540 2496 548 2504
rect 588 2476 596 2484
rect 636 2456 644 2464
rect 812 2616 820 2624
rect 796 2596 804 2604
rect 780 2576 788 2584
rect 876 2656 884 2664
rect 972 2656 980 2664
rect 1068 2656 1076 2664
rect 972 2636 980 2644
rect 908 2616 916 2624
rect 940 2616 948 2624
rect 844 2536 852 2544
rect 892 2536 900 2544
rect 1004 2616 1012 2624
rect 1020 2536 1028 2544
rect 892 2516 900 2524
rect 988 2516 996 2524
rect 620 2356 628 2364
rect 492 2336 500 2344
rect 620 2336 628 2344
rect 460 2316 468 2324
rect 588 2316 596 2324
rect 220 2296 228 2304
rect 380 2296 388 2304
rect 412 2296 420 2304
rect 428 2296 436 2304
rect 332 2276 340 2284
rect 460 2276 468 2284
rect 556 2276 564 2284
rect 588 2276 596 2284
rect 652 2396 660 2404
rect 668 2356 676 2364
rect 988 2476 996 2484
rect 1164 2656 1172 2664
rect 1292 2656 1300 2664
rect 1196 2636 1204 2644
rect 1260 2616 1268 2624
rect 1244 2576 1252 2584
rect 1324 2596 1332 2604
rect 1388 2576 1396 2584
rect 1276 2556 1284 2564
rect 1324 2556 1332 2564
rect 1356 2556 1364 2564
rect 1420 2556 1428 2564
rect 2108 2676 2116 2684
rect 2124 2676 2132 2684
rect 2172 2676 2180 2684
rect 2364 2956 2372 2964
rect 2524 2956 2532 2964
rect 2572 2956 2580 2964
rect 2348 2916 2356 2924
rect 2396 2916 2404 2924
rect 2428 2916 2436 2924
rect 2476 2896 2484 2904
rect 2300 2856 2308 2864
rect 2396 2856 2404 2864
rect 2444 2856 2452 2864
rect 2476 2836 2484 2844
rect 2268 2796 2276 2804
rect 2300 2796 2308 2804
rect 2316 2756 2324 2764
rect 2412 2756 2420 2764
rect 2332 2736 2340 2744
rect 2444 2736 2452 2744
rect 2460 2716 2468 2724
rect 2204 2676 2212 2684
rect 2252 2676 2260 2684
rect 2668 2956 2676 2964
rect 2764 2956 2772 2964
rect 2780 2956 2788 2964
rect 2972 2976 2980 2984
rect 3004 2976 3012 2984
rect 3164 2976 3172 2984
rect 3836 2976 3844 2984
rect 3996 2976 4004 2984
rect 2844 2956 2852 2964
rect 3468 2956 3476 2964
rect 3548 2956 3556 2964
rect 3564 2956 3572 2964
rect 3708 2956 3716 2964
rect 3948 2956 3956 2964
rect 4060 2956 4068 2964
rect 2844 2936 2852 2944
rect 2892 2936 2900 2944
rect 2924 2936 2932 2944
rect 2956 2936 2964 2944
rect 2988 2936 2996 2944
rect 3244 2936 3252 2944
rect 3260 2936 3268 2944
rect 3292 2936 3300 2944
rect 3372 2936 3380 2944
rect 3580 2936 3588 2944
rect 3628 2936 3636 2944
rect 3116 2916 3124 2924
rect 3148 2916 3156 2924
rect 3212 2916 3220 2924
rect 3276 2916 3284 2924
rect 3500 2916 3508 2924
rect 3532 2916 3540 2924
rect 2604 2896 2612 2904
rect 2684 2896 2692 2904
rect 3068 2896 3076 2904
rect 2556 2856 2564 2864
rect 2652 2796 2660 2804
rect 2812 2876 2820 2884
rect 2524 2736 2532 2744
rect 2796 2736 2804 2744
rect 2524 2716 2532 2724
rect 2636 2716 2644 2724
rect 2780 2716 2788 2724
rect 2508 2696 2516 2704
rect 3132 2876 3140 2884
rect 3180 2876 3188 2884
rect 2892 2796 2900 2804
rect 3020 2736 3028 2744
rect 2812 2716 2820 2724
rect 2876 2716 2884 2724
rect 3004 2716 3012 2724
rect 3132 2836 3140 2844
rect 3500 2856 3508 2864
rect 3420 2816 3428 2824
rect 3340 2796 3348 2804
rect 3132 2736 3140 2744
rect 3324 2736 3332 2744
rect 3228 2716 3236 2724
rect 3468 2716 3476 2724
rect 3148 2696 3156 2704
rect 1548 2656 1556 2664
rect 1564 2656 1572 2664
rect 1820 2656 1828 2664
rect 1836 2656 1844 2664
rect 2076 2656 2084 2664
rect 2172 2656 2180 2664
rect 2188 2656 2196 2664
rect 2348 2656 2356 2664
rect 2444 2656 2452 2664
rect 2508 2656 2516 2664
rect 2540 2656 2548 2664
rect 1468 2636 1476 2644
rect 1660 2636 1668 2644
rect 1564 2596 1572 2604
rect 1660 2596 1668 2604
rect 1484 2556 1492 2564
rect 1500 2556 1508 2564
rect 1548 2556 1556 2564
rect 1628 2556 1636 2564
rect 1116 2536 1124 2544
rect 1132 2496 1140 2504
rect 1372 2496 1380 2504
rect 1404 2496 1412 2504
rect 1436 2496 1444 2504
rect 940 2416 948 2424
rect 972 2416 980 2424
rect 1036 2416 1044 2424
rect 764 2396 772 2404
rect 940 2396 948 2404
rect 780 2296 788 2304
rect 732 2276 740 2284
rect 12 2256 20 2264
rect 92 2256 100 2264
rect 188 2256 196 2264
rect 284 2256 292 2264
rect 428 2256 436 2264
rect 492 2256 500 2264
rect 556 2256 564 2264
rect 828 2256 836 2264
rect 12 2236 20 2244
rect 204 2236 212 2244
rect 588 2236 596 2244
rect 12 2196 20 2204
rect 204 2216 212 2224
rect 156 2196 164 2204
rect 60 2176 68 2184
rect 124 2176 132 2184
rect 140 2176 148 2184
rect 252 2196 260 2204
rect 508 2196 516 2204
rect 28 2156 36 2164
rect 60 2156 68 2164
rect 252 2156 260 2164
rect 316 2156 324 2164
rect 540 2156 548 2164
rect 60 2136 68 2144
rect 92 2136 100 2144
rect 108 2136 116 2144
rect 220 2136 228 2144
rect 428 2136 436 2144
rect 172 2116 180 2124
rect 284 2116 292 2124
rect 316 2116 324 2124
rect 348 2116 356 2124
rect 476 2116 484 2124
rect 524 2116 532 2124
rect 668 2236 676 2244
rect 844 2236 852 2244
rect 892 2236 900 2244
rect 604 2156 612 2164
rect 748 2176 756 2184
rect 636 2116 644 2124
rect 652 2116 660 2124
rect 732 2116 740 2124
rect 284 2096 292 2104
rect 316 2096 324 2104
rect 556 2096 564 2104
rect 396 2076 404 2084
rect 44 1956 52 1964
rect 92 1936 100 1944
rect 172 1976 180 1984
rect 236 1996 244 2004
rect 188 1936 196 1944
rect 76 1896 84 1904
rect 124 1896 132 1904
rect 140 1896 148 1904
rect 380 2056 388 2064
rect 604 2056 612 2064
rect 348 1976 356 1984
rect 316 1956 324 1964
rect 268 1936 276 1944
rect 300 1896 308 1904
rect 844 2176 852 2184
rect 988 2356 996 2364
rect 1052 2356 1060 2364
rect 1148 2376 1156 2384
rect 1180 2376 1188 2384
rect 1724 2636 1732 2644
rect 1772 2636 1780 2644
rect 1740 2596 1748 2604
rect 1804 2596 1812 2604
rect 1916 2636 1924 2644
rect 1868 2616 1876 2624
rect 1852 2596 1860 2604
rect 1868 2596 1876 2604
rect 1692 2556 1700 2564
rect 1724 2556 1732 2564
rect 1788 2536 1796 2544
rect 1516 2496 1524 2504
rect 1580 2496 1588 2504
rect 1676 2496 1684 2504
rect 1532 2436 1540 2444
rect 1580 2436 1588 2444
rect 1612 2436 1620 2444
rect 1564 2416 1572 2424
rect 1372 2356 1380 2364
rect 1436 2356 1444 2364
rect 1500 2356 1508 2364
rect 1564 2356 1572 2364
rect 1132 2336 1140 2344
rect 1164 2336 1172 2344
rect 1004 2316 1012 2324
rect 1036 2316 1044 2324
rect 1084 2316 1092 2324
rect 1196 2316 1204 2324
rect 1324 2336 1332 2344
rect 1196 2276 1204 2284
rect 972 2236 980 2244
rect 1036 2236 1044 2244
rect 1116 2236 1124 2244
rect 940 2176 948 2184
rect 828 2156 836 2164
rect 1052 2216 1060 2224
rect 1116 2196 1124 2204
rect 1164 2196 1172 2204
rect 988 2176 996 2184
rect 1084 2176 1092 2184
rect 1244 2236 1252 2244
rect 1324 2296 1332 2304
rect 1404 2336 1412 2344
rect 1420 2336 1428 2344
rect 1548 2316 1556 2324
rect 1388 2256 1396 2264
rect 1452 2256 1460 2264
rect 1484 2256 1492 2264
rect 1292 2236 1300 2244
rect 1356 2236 1364 2244
rect 1468 2236 1476 2244
rect 1516 2236 1524 2244
rect 1308 2216 1316 2224
rect 1356 2216 1364 2224
rect 1324 2196 1332 2204
rect 1212 2176 1220 2184
rect 1244 2176 1252 2184
rect 1260 2176 1268 2184
rect 1308 2176 1316 2184
rect 1068 2136 1076 2144
rect 1116 2136 1124 2144
rect 1180 2136 1188 2144
rect 780 2116 788 2124
rect 828 2116 836 2124
rect 892 2116 900 2124
rect 1036 2116 1044 2124
rect 1052 2116 1060 2124
rect 812 2096 820 2104
rect 860 2096 868 2104
rect 636 1976 644 1984
rect 732 1976 740 1984
rect 620 1956 628 1964
rect 668 1936 676 1944
rect 780 2076 788 2084
rect 764 2056 772 2064
rect 876 2036 884 2044
rect 796 1936 804 1944
rect 540 1916 548 1924
rect 716 1916 724 1924
rect 748 1916 756 1924
rect 828 1916 836 1924
rect 876 1916 884 1924
rect 12 1876 20 1884
rect 44 1876 52 1884
rect 332 1876 340 1884
rect 28 1856 36 1864
rect 124 1856 132 1864
rect 252 1856 260 1864
rect 12 1776 20 1784
rect 364 1836 372 1844
rect 444 1836 452 1844
rect 284 1796 292 1804
rect 300 1776 308 1784
rect 908 2076 916 2084
rect 1020 2076 1028 2084
rect 908 1936 916 1944
rect 956 1936 964 1944
rect 844 1896 852 1904
rect 1212 2116 1220 2124
rect 1740 2496 1748 2504
rect 1788 2496 1796 2504
rect 1836 2516 1844 2524
rect 1804 2476 1812 2484
rect 1932 2576 1940 2584
rect 1916 2536 1924 2544
rect 1900 2516 1908 2524
rect 1868 2476 1876 2484
rect 1820 2456 1828 2464
rect 1852 2456 1860 2464
rect 1724 2396 1732 2404
rect 1852 2396 1860 2404
rect 1708 2376 1716 2384
rect 1612 2356 1620 2364
rect 1836 2356 1844 2364
rect 1884 2356 1892 2364
rect 1436 2176 1444 2184
rect 1628 2256 1636 2264
rect 1596 2236 1604 2244
rect 1676 2256 1684 2264
rect 1804 2256 1812 2264
rect 1836 2256 1844 2264
rect 1884 2256 1892 2264
rect 1900 2256 1908 2264
rect 1612 2176 1620 2184
rect 1724 2236 1732 2244
rect 1756 2236 1764 2244
rect 1788 2236 1796 2244
rect 1820 2236 1828 2244
rect 1868 2236 1876 2244
rect 1708 2216 1716 2224
rect 1756 2176 1764 2184
rect 1852 2176 1860 2184
rect 1900 2176 1908 2184
rect 1932 2176 1940 2184
rect 1420 2156 1428 2164
rect 1468 2156 1476 2164
rect 1580 2156 1588 2164
rect 1660 2156 1668 2164
rect 1708 2156 1716 2164
rect 1788 2156 1796 2164
rect 1804 2156 1812 2164
rect 1836 2156 1844 2164
rect 1884 2156 1892 2164
rect 1916 2156 1924 2164
rect 1292 2136 1300 2144
rect 1324 2136 1332 2144
rect 1308 2116 1316 2124
rect 1340 2116 1348 2124
rect 1388 2136 1396 2144
rect 1340 2096 1348 2104
rect 1372 2096 1380 2104
rect 1084 2036 1092 2044
rect 1500 2136 1508 2144
rect 1596 2136 1604 2144
rect 1660 2136 1668 2144
rect 1244 2076 1252 2084
rect 1404 2076 1412 2084
rect 1164 2036 1172 2044
rect 1580 2116 1588 2124
rect 1708 2116 1716 2124
rect 1356 2016 1364 2024
rect 1420 2016 1428 2024
rect 1212 1996 1220 2004
rect 1692 2076 1700 2084
rect 1724 2076 1732 2084
rect 1740 2076 1748 2084
rect 1708 2056 1716 2064
rect 1628 2036 1636 2044
rect 1692 2016 1700 2024
rect 1724 2016 1732 2024
rect 1532 1996 1540 2004
rect 1612 1996 1620 2004
rect 1484 1936 1492 1944
rect 1532 1936 1540 1944
rect 1564 1936 1572 1944
rect 1644 1956 1652 1964
rect 1804 2076 1812 2084
rect 1836 2076 1844 2084
rect 1932 2056 1940 2064
rect 1740 1956 1748 1964
rect 1788 1956 1796 1964
rect 1724 1936 1732 1944
rect 1884 1916 1892 1924
rect 1692 1896 1700 1904
rect 508 1876 516 1884
rect 940 1876 948 1884
rect 1020 1876 1028 1884
rect 1036 1876 1044 1884
rect 1132 1876 1140 1884
rect 1164 1876 1172 1884
rect 1180 1876 1188 1884
rect 1228 1876 1236 1884
rect 1308 1876 1316 1884
rect 1388 1876 1396 1884
rect 1660 1876 1668 1884
rect 1724 1876 1732 1884
rect 1836 1876 1844 1884
rect 1868 1876 1876 1884
rect 1900 1876 1908 1884
rect 1932 1876 1940 1884
rect 636 1856 644 1864
rect 716 1836 724 1844
rect 684 1796 692 1804
rect 124 1756 132 1764
rect 316 1756 324 1764
rect 332 1756 340 1764
rect 476 1756 484 1764
rect 508 1756 516 1764
rect 652 1756 660 1764
rect 12 1736 20 1744
rect 236 1736 244 1744
rect 268 1736 276 1744
rect 348 1736 356 1744
rect 124 1596 132 1604
rect 76 1556 84 1564
rect 172 1576 180 1584
rect 124 1496 132 1504
rect 156 1476 164 1484
rect 188 1476 196 1484
rect 76 1456 84 1464
rect 108 1456 116 1464
rect 76 1376 84 1384
rect 108 1356 116 1364
rect 220 1596 228 1604
rect 220 1576 228 1584
rect 236 1556 244 1564
rect 492 1736 500 1744
rect 700 1776 708 1784
rect 764 1836 772 1844
rect 812 1836 820 1844
rect 780 1816 788 1824
rect 748 1756 756 1764
rect 764 1676 772 1684
rect 348 1596 356 1604
rect 396 1596 404 1604
rect 428 1596 436 1604
rect 492 1596 500 1604
rect 588 1596 596 1604
rect 460 1556 468 1564
rect 508 1556 516 1564
rect 716 1556 724 1564
rect 492 1516 500 1524
rect 524 1516 532 1524
rect 588 1516 596 1524
rect 620 1516 628 1524
rect 428 1496 436 1504
rect 300 1476 308 1484
rect 588 1476 596 1484
rect 268 1456 276 1464
rect 316 1456 324 1464
rect 412 1456 420 1464
rect 204 1416 212 1424
rect 204 1396 212 1404
rect 140 1356 148 1364
rect 332 1436 340 1444
rect 380 1436 388 1444
rect 220 1376 228 1384
rect 252 1356 260 1364
rect 44 1336 52 1344
rect 220 1336 228 1344
rect 300 1416 308 1424
rect 444 1416 452 1424
rect 524 1436 532 1444
rect 444 1396 452 1404
rect 620 1456 628 1464
rect 732 1516 740 1524
rect 748 1496 756 1504
rect 940 1796 948 1804
rect 828 1756 836 1764
rect 1004 1816 1012 1824
rect 1116 1856 1124 1864
rect 1340 1856 1348 1864
rect 1244 1836 1252 1844
rect 1292 1836 1300 1844
rect 860 1756 868 1764
rect 972 1756 980 1764
rect 1052 1756 1060 1764
rect 924 1716 932 1724
rect 796 1636 804 1644
rect 812 1636 820 1644
rect 780 1616 788 1624
rect 780 1596 788 1604
rect 972 1596 980 1604
rect 1180 1796 1188 1804
rect 1276 1776 1284 1784
rect 1372 1836 1380 1844
rect 1404 1836 1412 1844
rect 1452 1836 1460 1844
rect 1484 1836 1492 1844
rect 1564 1836 1572 1844
rect 1420 1796 1428 1804
rect 1340 1776 1348 1784
rect 1356 1776 1364 1784
rect 1100 1756 1108 1764
rect 1148 1756 1156 1764
rect 1180 1756 1188 1764
rect 1292 1756 1300 1764
rect 1324 1756 1332 1764
rect 1484 1756 1492 1764
rect 1628 1836 1636 1844
rect 1756 1836 1764 1844
rect 1788 1836 1796 1844
rect 1676 1796 1684 1804
rect 1596 1776 1604 1784
rect 1532 1756 1540 1764
rect 1580 1756 1588 1764
rect 1612 1756 1620 1764
rect 1340 1736 1348 1744
rect 1372 1736 1380 1744
rect 1084 1656 1092 1664
rect 1020 1576 1028 1584
rect 860 1556 868 1564
rect 1004 1536 1012 1544
rect 892 1516 900 1524
rect 924 1516 932 1524
rect 812 1496 820 1504
rect 844 1496 852 1504
rect 1036 1496 1044 1504
rect 1292 1716 1300 1724
rect 1324 1716 1332 1724
rect 1404 1716 1412 1724
rect 1452 1716 1460 1724
rect 1852 1816 1860 1824
rect 1740 1776 1748 1784
rect 1820 1776 1828 1784
rect 1980 2616 1988 2624
rect 2044 2636 2052 2644
rect 2108 2636 2116 2644
rect 2028 2616 2036 2624
rect 2124 2616 2132 2624
rect 2236 2616 2244 2624
rect 2156 2596 2164 2604
rect 2396 2636 2404 2644
rect 2460 2636 2468 2644
rect 2444 2616 2452 2624
rect 2300 2556 2308 2564
rect 2012 2536 2020 2544
rect 1964 2516 1972 2524
rect 1996 2516 2004 2524
rect 2092 2516 2100 2524
rect 2108 2516 2116 2524
rect 2188 2516 2196 2524
rect 2060 2476 2068 2484
rect 1964 2456 1972 2464
rect 2156 2476 2164 2484
rect 2284 2516 2292 2524
rect 2236 2496 2244 2504
rect 2316 2496 2324 2504
rect 2140 2396 2148 2404
rect 2204 2396 2212 2404
rect 2236 2396 2244 2404
rect 2012 2376 2020 2384
rect 2076 2376 2084 2384
rect 2044 2336 2052 2344
rect 1980 2296 1988 2304
rect 1964 2176 1972 2184
rect 2348 2516 2356 2524
rect 2364 2496 2372 2504
rect 2268 2356 2276 2364
rect 2332 2356 2340 2364
rect 2092 2336 2100 2344
rect 2140 2336 2148 2344
rect 2220 2336 2228 2344
rect 2460 2376 2468 2384
rect 2572 2656 2580 2664
rect 2636 2656 2644 2664
rect 2684 2656 2692 2664
rect 2732 2656 2740 2664
rect 2556 2616 2564 2624
rect 2636 2596 2644 2604
rect 2940 2616 2948 2624
rect 2956 2616 2964 2624
rect 2972 2616 2980 2624
rect 3052 2616 3060 2624
rect 2924 2596 2932 2604
rect 2764 2576 2772 2584
rect 2796 2576 2804 2584
rect 2892 2576 2900 2584
rect 2492 2516 2500 2524
rect 2540 2516 2548 2524
rect 2588 2516 2596 2524
rect 2972 2576 2980 2584
rect 2876 2536 2884 2544
rect 2940 2536 2948 2544
rect 2972 2536 2980 2544
rect 3004 2536 3012 2544
rect 3036 2536 3044 2544
rect 3052 2536 3060 2544
rect 2620 2516 2628 2524
rect 2684 2516 2692 2524
rect 2764 2516 2772 2524
rect 2828 2516 2836 2524
rect 2700 2496 2708 2504
rect 2860 2496 2868 2504
rect 2028 2276 2036 2284
rect 2044 2276 2052 2284
rect 2092 2276 2100 2284
rect 2124 2276 2132 2284
rect 2140 2276 2148 2284
rect 2204 2276 2212 2284
rect 2316 2276 2324 2284
rect 2348 2276 2356 2284
rect 2412 2276 2420 2284
rect 2444 2276 2452 2284
rect 2028 2256 2036 2264
rect 1996 2176 2004 2184
rect 2300 2216 2308 2224
rect 2236 2196 2244 2204
rect 2364 2196 2372 2204
rect 2604 2416 2612 2424
rect 2604 2376 2612 2384
rect 2716 2436 2724 2444
rect 2828 2376 2836 2384
rect 2780 2336 2788 2344
rect 2556 2316 2564 2324
rect 2588 2316 2596 2324
rect 2508 2276 2516 2284
rect 2508 2256 2516 2264
rect 2556 2236 2564 2244
rect 2588 2236 2596 2244
rect 2652 2236 2660 2244
rect 2684 2236 2692 2244
rect 2492 2216 2500 2224
rect 2604 2216 2612 2224
rect 2540 2196 2548 2204
rect 2860 2336 2868 2344
rect 3036 2496 3044 2504
rect 3132 2676 3140 2684
rect 3132 2636 3140 2644
rect 3084 2596 3092 2604
rect 3100 2596 3108 2604
rect 3660 2916 3668 2924
rect 3676 2916 3684 2924
rect 3708 2916 3716 2924
rect 3740 2916 3748 2924
rect 3644 2896 3652 2904
rect 3724 2876 3732 2884
rect 3836 2896 3844 2904
rect 3884 2896 3892 2904
rect 3756 2876 3764 2884
rect 3964 2896 3972 2904
rect 3948 2856 3956 2864
rect 3740 2816 3748 2824
rect 3772 2756 3780 2764
rect 3676 2736 3684 2744
rect 3516 2716 3524 2724
rect 3564 2716 3572 2724
rect 3580 2716 3588 2724
rect 3596 2716 3604 2724
rect 3660 2716 3668 2724
rect 3724 2716 3732 2724
rect 3756 2716 3764 2724
rect 3932 2816 3940 2824
rect 3884 2776 3892 2784
rect 3836 2756 3844 2764
rect 3852 2716 3860 2724
rect 3628 2696 3636 2704
rect 3820 2696 3828 2704
rect 4140 2936 4148 2944
rect 4156 2896 4164 2904
rect 4076 2876 4084 2884
rect 4060 2776 4068 2784
rect 4044 2756 4052 2764
rect 3900 2716 3908 2724
rect 4124 2796 4132 2804
rect 4204 2796 4212 2804
rect 4092 2776 4100 2784
rect 4156 2756 4164 2764
rect 4108 2736 4116 2744
rect 3548 2676 3556 2684
rect 3644 2676 3652 2684
rect 3932 2676 3940 2684
rect 3404 2656 3412 2664
rect 3276 2636 3284 2644
rect 3164 2616 3172 2624
rect 3164 2596 3172 2604
rect 3260 2596 3268 2604
rect 3468 2616 3476 2624
rect 3436 2596 3444 2604
rect 3500 2596 3508 2604
rect 3532 2596 3540 2604
rect 3724 2656 3732 2664
rect 3820 2656 3828 2664
rect 3980 2656 3988 2664
rect 4108 2656 4116 2664
rect 4140 2656 4148 2664
rect 3708 2576 3716 2584
rect 3804 2576 3812 2584
rect 3884 2596 3892 2604
rect 3980 2616 3988 2624
rect 3916 2596 3924 2604
rect 4156 2596 4164 2604
rect 4188 2596 4196 2604
rect 3900 2576 3908 2584
rect 3964 2576 3972 2584
rect 4044 2576 4052 2584
rect 4092 2576 4100 2584
rect 3308 2536 3316 2544
rect 3356 2536 3364 2544
rect 3084 2496 3092 2504
rect 3196 2496 3204 2504
rect 2908 2456 2916 2464
rect 2988 2456 2996 2464
rect 3068 2456 3076 2464
rect 3196 2436 3204 2444
rect 2908 2416 2916 2424
rect 2892 2356 2900 2364
rect 3084 2356 3092 2364
rect 2940 2336 2948 2344
rect 2972 2336 2980 2344
rect 2988 2336 2996 2344
rect 2988 2316 2996 2324
rect 3020 2316 3028 2324
rect 2876 2276 2884 2284
rect 2812 2256 2820 2264
rect 3020 2256 3028 2264
rect 3068 2256 3076 2264
rect 2748 2236 2756 2244
rect 3100 2236 3108 2244
rect 2700 2216 2708 2224
rect 2844 2216 2852 2224
rect 2908 2196 2916 2204
rect 3036 2176 3044 2184
rect 3052 2176 3060 2184
rect 3084 2176 3092 2184
rect 2492 2156 2500 2164
rect 2524 2156 2532 2164
rect 2556 2156 2564 2164
rect 2764 2156 2772 2164
rect 1964 2136 1972 2144
rect 2028 2116 2036 2124
rect 2124 2116 2132 2124
rect 1996 2076 2004 2084
rect 2012 2056 2020 2064
rect 2012 1996 2020 2004
rect 2076 2056 2084 2064
rect 2060 2016 2068 2024
rect 1964 1896 1972 1904
rect 1980 1896 1988 1904
rect 1996 1896 2004 1904
rect 1980 1876 1988 1884
rect 2108 2016 2116 2024
rect 2684 2136 2692 2144
rect 2268 2116 2276 2124
rect 2332 2116 2340 2124
rect 2380 2116 2388 2124
rect 2236 2096 2244 2104
rect 2236 2076 2244 2084
rect 2172 2036 2180 2044
rect 2108 1996 2116 2004
rect 2156 1996 2164 2004
rect 2076 1956 2084 1964
rect 2012 1876 2020 1884
rect 2044 1876 2052 1884
rect 1948 1816 1956 1824
rect 1996 1816 2004 1824
rect 1868 1796 1876 1804
rect 1900 1796 1908 1804
rect 1916 1776 1924 1784
rect 2124 1956 2132 1964
rect 2140 1956 2148 1964
rect 2108 1916 2116 1924
rect 2092 1896 2100 1904
rect 2252 1956 2260 1964
rect 2076 1796 2084 1804
rect 2140 1836 2148 1844
rect 2156 1836 2164 1844
rect 2124 1816 2132 1824
rect 1948 1756 1956 1764
rect 2044 1756 2052 1764
rect 1596 1736 1604 1744
rect 1852 1736 1860 1744
rect 1884 1736 1892 1744
rect 1660 1716 1668 1724
rect 1788 1716 1796 1724
rect 1212 1696 1220 1704
rect 1132 1676 1140 1684
rect 1196 1616 1204 1624
rect 1612 1676 1620 1684
rect 1164 1576 1172 1584
rect 1324 1576 1332 1584
rect 1372 1576 1380 1584
rect 1484 1576 1492 1584
rect 1132 1556 1140 1564
rect 1612 1576 1620 1584
rect 1340 1556 1348 1564
rect 1564 1556 1572 1564
rect 1196 1516 1204 1524
rect 1244 1516 1252 1524
rect 1356 1516 1364 1524
rect 1452 1516 1460 1524
rect 1820 1636 1828 1644
rect 1740 1616 1748 1624
rect 1692 1556 1700 1564
rect 1420 1496 1428 1504
rect 1884 1616 1892 1624
rect 1852 1596 1860 1604
rect 1868 1576 1876 1584
rect 1884 1556 1892 1564
rect 2060 1716 2068 1724
rect 1932 1676 1940 1684
rect 1948 1676 1956 1684
rect 684 1476 692 1484
rect 732 1476 740 1484
rect 876 1476 884 1484
rect 924 1476 932 1484
rect 956 1476 964 1484
rect 1100 1476 1108 1484
rect 1132 1476 1140 1484
rect 1212 1476 1220 1484
rect 1260 1476 1268 1484
rect 1292 1476 1300 1484
rect 1580 1476 1588 1484
rect 1692 1476 1700 1484
rect 1836 1476 1844 1484
rect 652 1436 660 1444
rect 428 1376 436 1384
rect 380 1356 388 1364
rect 396 1356 404 1364
rect 460 1356 468 1364
rect 92 1276 100 1284
rect 220 1156 228 1164
rect 364 1336 372 1344
rect 476 1336 484 1344
rect 540 1336 548 1344
rect 236 1116 244 1124
rect 76 1076 84 1084
rect 284 1076 292 1084
rect 92 1056 100 1064
rect 92 1036 100 1044
rect 188 1036 196 1044
rect 124 976 132 984
rect 188 976 196 984
rect 284 1016 292 1024
rect 412 1136 420 1144
rect 332 1116 340 1124
rect 316 1076 324 1084
rect 364 1076 372 1084
rect 380 1056 388 1064
rect 348 1036 356 1044
rect 124 956 132 964
rect 156 956 164 964
rect 236 936 244 944
rect 60 916 68 924
rect 92 896 100 904
rect 44 736 52 744
rect 588 1336 596 1344
rect 652 1316 660 1324
rect 652 1296 660 1304
rect 604 1256 612 1264
rect 492 1196 500 1204
rect 556 1196 564 1204
rect 460 1136 468 1144
rect 428 1096 436 1104
rect 668 1256 676 1264
rect 620 1156 628 1164
rect 588 1136 596 1144
rect 508 1096 516 1104
rect 540 1096 548 1104
rect 604 1096 612 1104
rect 636 1096 644 1104
rect 620 1076 628 1084
rect 524 1056 532 1064
rect 556 1056 564 1064
rect 428 1036 436 1044
rect 492 1036 500 1044
rect 444 976 452 984
rect 828 1436 836 1444
rect 876 1436 884 1444
rect 796 1376 804 1384
rect 844 1376 852 1384
rect 732 1356 740 1364
rect 764 1356 772 1364
rect 892 1416 900 1424
rect 1116 1436 1124 1444
rect 1164 1436 1172 1444
rect 1212 1436 1220 1444
rect 1068 1376 1076 1384
rect 956 1356 964 1364
rect 1020 1356 1028 1364
rect 1052 1356 1060 1364
rect 1244 1396 1252 1404
rect 748 1336 756 1344
rect 796 1336 804 1344
rect 1020 1336 1028 1344
rect 1308 1436 1316 1444
rect 1372 1436 1380 1444
rect 1372 1416 1380 1424
rect 1436 1416 1444 1424
rect 1500 1456 1508 1464
rect 1532 1456 1540 1464
rect 1628 1456 1636 1464
rect 1708 1456 1716 1464
rect 1788 1456 1796 1464
rect 1468 1436 1476 1444
rect 1548 1416 1556 1424
rect 1596 1416 1604 1424
rect 1548 1396 1556 1404
rect 1308 1376 1316 1384
rect 1420 1376 1428 1384
rect 1452 1376 1460 1384
rect 1516 1356 1524 1364
rect 1564 1356 1572 1364
rect 1340 1336 1348 1344
rect 1404 1336 1412 1344
rect 700 1316 708 1324
rect 828 1316 836 1324
rect 1100 1316 1108 1324
rect 1212 1316 1220 1324
rect 1292 1316 1300 1324
rect 940 1296 948 1304
rect 956 1296 964 1304
rect 1004 1296 1012 1304
rect 1068 1296 1076 1304
rect 796 1276 804 1284
rect 924 1236 932 1244
rect 844 1216 852 1224
rect 764 1176 772 1184
rect 716 1136 724 1144
rect 764 1136 772 1144
rect 844 1176 852 1184
rect 892 1136 900 1144
rect 860 1096 868 1104
rect 1052 1276 1060 1284
rect 972 1236 980 1244
rect 988 1236 996 1244
rect 972 1136 980 1144
rect 1004 1136 1012 1144
rect 1180 1176 1188 1184
rect 1100 1116 1108 1124
rect 940 1096 948 1104
rect 1308 1296 1316 1304
rect 1292 1276 1300 1284
rect 732 1076 740 1084
rect 1132 1076 1140 1084
rect 1084 1056 1092 1064
rect 1212 1056 1220 1064
rect 716 1036 724 1044
rect 796 1036 804 1044
rect 844 1036 852 1044
rect 908 1036 916 1044
rect 956 1036 964 1044
rect 972 1036 980 1044
rect 588 996 596 1004
rect 620 996 628 1004
rect 684 996 692 1004
rect 508 976 516 984
rect 588 976 596 984
rect 652 976 660 984
rect 300 956 308 964
rect 364 956 372 964
rect 428 956 436 964
rect 460 956 468 964
rect 684 956 692 964
rect 860 1016 868 1024
rect 812 996 820 1004
rect 876 996 884 1004
rect 892 996 900 1004
rect 780 976 788 984
rect 828 976 836 984
rect 972 1016 980 1024
rect 908 976 916 984
rect 1004 996 1012 1004
rect 1036 996 1044 1004
rect 988 976 996 984
rect 1068 956 1076 964
rect 1196 976 1204 984
rect 1132 956 1140 964
rect 1372 1316 1380 1324
rect 1356 1296 1364 1304
rect 1388 1296 1396 1304
rect 1340 1236 1348 1244
rect 1276 1116 1284 1124
rect 1324 1116 1332 1124
rect 1244 1096 1252 1104
rect 1244 1056 1252 1064
rect 1404 1056 1412 1064
rect 1500 1336 1508 1344
rect 1660 1416 1668 1424
rect 1724 1416 1732 1424
rect 1756 1416 1764 1424
rect 1644 1396 1652 1404
rect 1772 1376 1780 1384
rect 1692 1336 1700 1344
rect 1756 1336 1764 1344
rect 1900 1496 1908 1504
rect 2108 1716 2116 1724
rect 2156 1716 2164 1724
rect 2124 1696 2132 1704
rect 2172 1696 2180 1704
rect 2076 1616 2084 1624
rect 2076 1596 2084 1604
rect 2092 1556 2100 1564
rect 2156 1656 2164 1664
rect 1948 1476 1956 1484
rect 2044 1476 2052 1484
rect 2028 1436 2036 1444
rect 1820 1356 1828 1364
rect 1884 1356 1892 1364
rect 2028 1356 2036 1364
rect 2092 1436 2100 1444
rect 2124 1436 2132 1444
rect 2076 1396 2084 1404
rect 2172 1596 2180 1604
rect 2444 2036 2452 2044
rect 2412 1996 2420 2004
rect 2316 1956 2324 1964
rect 2348 1956 2356 1964
rect 2396 1956 2404 1964
rect 2412 1916 2420 1924
rect 2428 1916 2436 1924
rect 2460 1996 2468 2004
rect 2892 2116 2900 2124
rect 2796 2096 2804 2104
rect 2908 2096 2916 2104
rect 2604 2076 2612 2084
rect 2572 2056 2580 2064
rect 2524 1956 2532 1964
rect 2652 2016 2660 2024
rect 2668 1996 2676 2004
rect 2748 1996 2756 2004
rect 2860 2076 2868 2084
rect 3244 2456 3252 2464
rect 3436 2536 3444 2544
rect 4188 2556 4196 2564
rect 3468 2536 3476 2544
rect 3500 2536 3508 2544
rect 3548 2536 3556 2544
rect 3660 2536 3668 2544
rect 3676 2536 3684 2544
rect 3772 2536 3780 2544
rect 3516 2496 3524 2504
rect 3612 2496 3620 2504
rect 3644 2496 3652 2504
rect 3436 2476 3444 2484
rect 3324 2456 3332 2464
rect 3340 2456 3348 2464
rect 3228 2396 3236 2404
rect 3260 2356 3268 2364
rect 3484 2396 3492 2404
rect 3436 2376 3444 2384
rect 3212 2296 3220 2304
rect 3308 2296 3316 2304
rect 3180 2256 3188 2264
rect 3228 2236 3236 2244
rect 3644 2396 3652 2404
rect 3564 2256 3572 2264
rect 3308 2236 3316 2244
rect 3436 2236 3444 2244
rect 3468 2236 3476 2244
rect 3516 2236 3524 2244
rect 3548 2236 3556 2244
rect 3276 2216 3284 2224
rect 3308 2216 3316 2224
rect 3372 2216 3380 2224
rect 3580 2236 3588 2244
rect 3916 2536 3924 2544
rect 4060 2536 4068 2544
rect 3852 2516 3860 2524
rect 3788 2496 3796 2504
rect 3820 2496 3828 2504
rect 3692 2476 3700 2484
rect 3852 2436 3860 2444
rect 3724 2376 3732 2384
rect 3932 2376 3940 2384
rect 4172 2516 4180 2524
rect 4220 2496 4228 2504
rect 4044 2416 4052 2424
rect 4124 2416 4132 2424
rect 3996 2376 4004 2384
rect 3676 2356 3684 2364
rect 3948 2356 3956 2364
rect 4060 2336 4068 2344
rect 3868 2316 3876 2324
rect 3900 2316 3908 2324
rect 3948 2316 3956 2324
rect 4012 2316 4020 2324
rect 4108 2316 4116 2324
rect 3804 2296 3812 2304
rect 3612 2236 3620 2244
rect 3436 2176 3444 2184
rect 3564 2176 3572 2184
rect 3564 2136 3572 2144
rect 3388 2116 3396 2124
rect 3564 2116 3572 2124
rect 3612 2156 3620 2164
rect 3628 2156 3636 2164
rect 3596 2136 3604 2144
rect 3660 2136 3668 2144
rect 3772 2256 3780 2264
rect 3724 2216 3732 2224
rect 3708 2176 3716 2184
rect 4092 2296 4100 2304
rect 4140 2296 4148 2304
rect 4156 2276 4164 2284
rect 3948 2256 3956 2264
rect 4028 2256 4036 2264
rect 4140 2256 4148 2264
rect 4188 2256 4196 2264
rect 3852 2216 3860 2224
rect 3900 2216 3908 2224
rect 3964 2216 3972 2224
rect 4252 2236 4260 2244
rect 3820 2196 3828 2204
rect 4012 2196 4020 2204
rect 4028 2176 4036 2184
rect 3692 2156 3700 2164
rect 3708 2156 3716 2164
rect 3884 2156 3892 2164
rect 3916 2156 3924 2164
rect 3756 2136 3764 2144
rect 3804 2136 3812 2144
rect 3724 2116 3732 2124
rect 3804 2116 3812 2124
rect 3836 2116 3844 2124
rect 3964 2136 3972 2144
rect 4060 2136 4068 2144
rect 4092 2176 4100 2184
rect 4124 2176 4132 2184
rect 4172 2156 4180 2164
rect 4140 2136 4148 2144
rect 2988 2096 2996 2104
rect 2940 2056 2948 2064
rect 3020 1996 3028 2004
rect 2844 1956 2852 1964
rect 2908 1956 2916 1964
rect 2588 1936 2596 1944
rect 2636 1936 2644 1944
rect 2844 1936 2852 1944
rect 2860 1936 2868 1944
rect 2908 1936 2916 1944
rect 2940 1936 2948 1944
rect 2476 1916 2484 1924
rect 2540 1916 2548 1924
rect 2892 1896 2900 1904
rect 3164 2096 3172 2104
rect 3356 2096 3364 2104
rect 3500 2096 3508 2104
rect 3932 2096 3940 2104
rect 3964 2096 3972 2104
rect 3996 2096 4004 2104
rect 4044 2096 4052 2104
rect 4076 2096 4084 2104
rect 3580 2076 3588 2084
rect 3580 2056 3588 2064
rect 3836 2056 3844 2064
rect 3420 2036 3428 2044
rect 3756 2036 3764 2044
rect 3100 2016 3108 2024
rect 3196 2016 3204 2024
rect 3116 1956 3124 1964
rect 3052 1936 3060 1944
rect 3228 1936 3236 1944
rect 3356 1996 3364 2004
rect 3404 1956 3412 1964
rect 3308 1916 3316 1924
rect 3340 1916 3348 1924
rect 3260 1896 3268 1904
rect 3292 1896 3300 1904
rect 3340 1896 3348 1904
rect 3452 1956 3460 1964
rect 3468 1956 3476 1964
rect 3596 1956 3604 1964
rect 3820 1936 3828 1944
rect 3420 1916 3428 1924
rect 3548 1916 3556 1924
rect 2492 1876 2500 1884
rect 2620 1876 2628 1884
rect 3004 1876 3012 1884
rect 3052 1876 3060 1884
rect 3180 1876 3188 1884
rect 3372 1876 3380 1884
rect 3516 1876 3524 1884
rect 3580 1876 3588 1884
rect 2300 1856 2308 1864
rect 2220 1836 2228 1844
rect 2284 1836 2292 1844
rect 2300 1836 2308 1844
rect 2540 1836 2548 1844
rect 2572 1836 2580 1844
rect 2396 1816 2404 1824
rect 2316 1796 2324 1804
rect 2380 1796 2388 1804
rect 2444 1796 2452 1804
rect 2204 1776 2212 1784
rect 2252 1776 2260 1784
rect 2428 1776 2436 1784
rect 2220 1756 2228 1764
rect 2300 1756 2308 1764
rect 2316 1756 2324 1764
rect 2204 1736 2212 1744
rect 2380 1756 2388 1764
rect 2412 1756 2420 1764
rect 2460 1756 2468 1764
rect 2492 1756 2500 1764
rect 2524 1756 2532 1764
rect 2300 1716 2308 1724
rect 2348 1716 2356 1724
rect 2252 1696 2260 1704
rect 2204 1656 2212 1664
rect 2284 1656 2292 1664
rect 2188 1556 2196 1564
rect 2252 1556 2260 1564
rect 2812 1856 2820 1864
rect 2924 1856 2932 1864
rect 2636 1836 2644 1844
rect 2732 1836 2740 1844
rect 2764 1776 2772 1784
rect 2556 1756 2564 1764
rect 2588 1756 2596 1764
rect 2716 1756 2724 1764
rect 2796 1756 2804 1764
rect 2844 1776 2852 1784
rect 2588 1736 2596 1744
rect 2748 1736 2756 1744
rect 2796 1736 2804 1744
rect 2620 1696 2628 1704
rect 2364 1616 2372 1624
rect 2380 1616 2388 1624
rect 2348 1536 2356 1544
rect 2428 1596 2436 1604
rect 2460 1596 2468 1604
rect 2524 1596 2532 1604
rect 2396 1536 2404 1544
rect 2332 1516 2340 1524
rect 2348 1516 2356 1524
rect 2396 1516 2404 1524
rect 2476 1536 2484 1544
rect 2668 1656 2676 1664
rect 2668 1596 2676 1604
rect 2860 1756 2868 1764
rect 3036 1836 3044 1844
rect 2956 1796 2964 1804
rect 3052 1796 3060 1804
rect 2812 1616 2820 1624
rect 2828 1616 2836 1624
rect 2428 1516 2436 1524
rect 2556 1516 2564 1524
rect 2636 1516 2644 1524
rect 2652 1516 2660 1524
rect 2796 1536 2804 1544
rect 2764 1516 2772 1524
rect 2444 1496 2452 1504
rect 2172 1476 2180 1484
rect 2268 1476 2276 1484
rect 2316 1476 2324 1484
rect 2460 1476 2468 1484
rect 2508 1476 2516 1484
rect 2588 1476 2596 1484
rect 2652 1496 2660 1504
rect 2620 1476 2628 1484
rect 2188 1436 2196 1444
rect 2396 1436 2404 1444
rect 2412 1436 2420 1444
rect 2140 1376 2148 1384
rect 2172 1376 2180 1384
rect 1804 1336 1812 1344
rect 1916 1336 1924 1344
rect 1756 1296 1764 1304
rect 1932 1296 1940 1304
rect 1436 1276 1444 1284
rect 1452 1276 1460 1284
rect 1484 1276 1492 1284
rect 1484 1256 1492 1264
rect 1596 1276 1604 1284
rect 1724 1276 1732 1284
rect 1740 1236 1748 1244
rect 1564 1216 1572 1224
rect 1612 1216 1620 1224
rect 1532 1196 1540 1204
rect 1532 1176 1540 1184
rect 1612 1196 1620 1204
rect 1596 1156 1604 1164
rect 2012 1296 2020 1304
rect 2332 1396 2340 1404
rect 2268 1376 2276 1384
rect 2348 1376 2356 1384
rect 2396 1416 2404 1424
rect 2204 1356 2212 1364
rect 2316 1356 2324 1364
rect 2428 1416 2436 1424
rect 2492 1456 2500 1464
rect 2540 1456 2548 1464
rect 2492 1436 2500 1444
rect 2460 1416 2468 1424
rect 2412 1396 2420 1404
rect 2444 1396 2452 1404
rect 2412 1376 2420 1384
rect 2476 1376 2484 1384
rect 2124 1336 2132 1344
rect 2188 1336 2196 1344
rect 2156 1296 2164 1304
rect 2140 1276 2148 1284
rect 2060 1236 2068 1244
rect 1852 1196 1860 1204
rect 1964 1196 1972 1204
rect 1692 1156 1700 1164
rect 1900 1156 1908 1164
rect 1660 1136 1668 1144
rect 1708 1136 1716 1144
rect 1804 1136 1812 1144
rect 1932 1136 1940 1144
rect 2284 1336 2292 1344
rect 2316 1316 2324 1324
rect 2396 1316 2404 1324
rect 2396 1276 2404 1284
rect 2252 1256 2260 1264
rect 2156 1196 2164 1204
rect 2204 1196 2212 1204
rect 2076 1176 2084 1184
rect 2028 1156 2036 1164
rect 2012 1136 2020 1144
rect 1644 1116 1652 1124
rect 1820 1116 1828 1124
rect 1228 1016 1236 1024
rect 1260 1016 1268 1024
rect 1420 1016 1428 1024
rect 1388 996 1396 1004
rect 1244 976 1252 984
rect 1356 976 1364 984
rect 2092 1156 2100 1164
rect 2220 1156 2228 1164
rect 2140 1136 2148 1144
rect 2172 1136 2180 1144
rect 2364 1216 2372 1224
rect 2316 1176 2324 1184
rect 2428 1356 2436 1364
rect 2476 1356 2484 1364
rect 2540 1416 2548 1424
rect 2508 1376 2516 1384
rect 2572 1416 2580 1424
rect 2972 1776 2980 1784
rect 3020 1776 3028 1784
rect 3068 1776 3076 1784
rect 3036 1696 3044 1704
rect 3068 1696 3076 1704
rect 2924 1676 2932 1684
rect 3004 1676 3012 1684
rect 2924 1616 2932 1624
rect 2908 1556 2916 1564
rect 2988 1556 2996 1564
rect 3068 1556 3076 1564
rect 2892 1516 2900 1524
rect 2940 1516 2948 1524
rect 2956 1516 2964 1524
rect 2908 1496 2916 1504
rect 2716 1476 2724 1484
rect 2764 1476 2772 1484
rect 2684 1456 2692 1464
rect 2716 1456 2724 1464
rect 2668 1396 2676 1404
rect 2572 1376 2580 1384
rect 2620 1376 2628 1384
rect 2508 1356 2516 1364
rect 2524 1356 2532 1364
rect 2588 1356 2596 1364
rect 2700 1356 2708 1364
rect 2524 1296 2532 1304
rect 2540 1296 2548 1304
rect 2572 1296 2580 1304
rect 2620 1296 2628 1304
rect 2668 1296 2676 1304
rect 2444 1256 2452 1264
rect 2508 1256 2516 1264
rect 2412 1216 2420 1224
rect 2284 1156 2292 1164
rect 2300 1156 2308 1164
rect 2380 1156 2388 1164
rect 2236 1136 2244 1144
rect 2396 1136 2404 1144
rect 2476 1136 2484 1144
rect 2652 1256 2660 1264
rect 2844 1456 2852 1464
rect 3020 1456 3028 1464
rect 2780 1436 2788 1444
rect 2828 1436 2836 1444
rect 2988 1436 2996 1444
rect 2844 1396 2852 1404
rect 2748 1376 2756 1384
rect 2764 1376 2772 1384
rect 2812 1376 2820 1384
rect 2764 1356 2772 1364
rect 2796 1356 2804 1364
rect 3292 1856 3300 1864
rect 3260 1816 3268 1824
rect 3100 1776 3108 1784
rect 3116 1776 3124 1784
rect 3308 1796 3316 1804
rect 3196 1776 3204 1784
rect 3388 1796 3396 1804
rect 3612 1836 3620 1844
rect 3468 1796 3476 1804
rect 3340 1756 3348 1764
rect 3164 1736 3172 1744
rect 3196 1736 3204 1744
rect 3196 1716 3204 1724
rect 3116 1696 3124 1704
rect 3260 1716 3268 1724
rect 3292 1716 3300 1724
rect 3308 1716 3316 1724
rect 3196 1676 3204 1684
rect 3244 1676 3252 1684
rect 3292 1676 3300 1684
rect 3212 1616 3220 1624
rect 3356 1676 3364 1684
rect 3372 1676 3380 1684
rect 3484 1776 3492 1784
rect 3500 1756 3508 1764
rect 3356 1656 3364 1664
rect 3388 1656 3396 1664
rect 3324 1596 3332 1604
rect 3340 1596 3348 1604
rect 3308 1556 3316 1564
rect 3388 1556 3396 1564
rect 3164 1516 3172 1524
rect 3132 1496 3140 1504
rect 3148 1496 3156 1504
rect 3244 1496 3252 1504
rect 3340 1496 3348 1504
rect 3532 1756 3540 1764
rect 3580 1816 3588 1824
rect 3612 1796 3620 1804
rect 3660 1836 3668 1844
rect 3740 1856 3748 1864
rect 3644 1776 3652 1784
rect 3820 1776 3828 1784
rect 3564 1756 3572 1764
rect 3628 1756 3636 1764
rect 3772 1756 3780 1764
rect 3836 1756 3844 1764
rect 3644 1736 3652 1744
rect 3916 2016 3924 2024
rect 3868 1916 3876 1924
rect 4124 2116 4132 2124
rect 4172 2096 4180 2104
rect 4204 2096 4212 2104
rect 3948 1936 3956 1944
rect 4028 1936 4036 1944
rect 4076 1936 4084 1944
rect 4108 1896 4116 1904
rect 3996 1876 4004 1884
rect 4076 1876 4084 1884
rect 4156 1876 4164 1884
rect 4220 1876 4228 1884
rect 3980 1856 3988 1864
rect 4044 1856 4052 1864
rect 4108 1856 4116 1864
rect 3932 1836 3940 1844
rect 4156 1836 4164 1844
rect 3980 1776 3988 1784
rect 4012 1776 4020 1784
rect 4172 1776 4180 1784
rect 4204 1776 4212 1784
rect 3884 1756 3892 1764
rect 4012 1756 4020 1764
rect 4044 1756 4052 1764
rect 4108 1756 4116 1764
rect 3868 1736 3876 1744
rect 3980 1736 3988 1744
rect 4028 1736 4036 1744
rect 4060 1736 4068 1744
rect 3676 1716 3684 1724
rect 3676 1696 3684 1704
rect 3708 1696 3716 1704
rect 3788 1676 3796 1684
rect 3532 1656 3540 1664
rect 3516 1616 3524 1624
rect 3436 1516 3444 1524
rect 3484 1516 3492 1524
rect 3436 1496 3444 1504
rect 3788 1656 3796 1664
rect 3708 1636 3716 1644
rect 3596 1616 3604 1624
rect 3660 1616 3668 1624
rect 3596 1556 3604 1564
rect 3564 1496 3572 1504
rect 3612 1496 3620 1504
rect 3644 1496 3652 1504
rect 3692 1596 3700 1604
rect 3692 1536 3700 1544
rect 3852 1716 3860 1724
rect 4076 1696 4084 1704
rect 3820 1636 3828 1644
rect 3980 1636 3988 1644
rect 4092 1636 4100 1644
rect 3804 1616 3812 1624
rect 3836 1556 3844 1564
rect 3964 1536 3972 1544
rect 3724 1496 3732 1504
rect 3884 1496 3892 1504
rect 3916 1496 3924 1504
rect 3260 1476 3268 1484
rect 3356 1476 3364 1484
rect 3484 1476 3492 1484
rect 3516 1476 3524 1484
rect 3100 1436 3108 1444
rect 3196 1436 3204 1444
rect 2940 1416 2948 1424
rect 3084 1416 3092 1424
rect 2972 1376 2980 1384
rect 3004 1376 3012 1384
rect 3036 1376 3044 1384
rect 3068 1376 3076 1384
rect 3100 1376 3108 1384
rect 3116 1376 3124 1384
rect 2924 1356 2932 1364
rect 2956 1356 2964 1364
rect 3084 1356 3092 1364
rect 2876 1336 2884 1344
rect 2924 1336 2932 1344
rect 2780 1296 2788 1304
rect 2796 1296 2804 1304
rect 2716 1236 2724 1244
rect 2716 1196 2724 1204
rect 2604 1176 2612 1184
rect 2460 1116 2468 1124
rect 1644 1076 1652 1084
rect 1660 1076 1668 1084
rect 1852 1076 1860 1084
rect 1964 1076 1972 1084
rect 1468 1056 1476 1064
rect 1484 1056 1492 1064
rect 1516 1056 1524 1064
rect 1612 1056 1620 1064
rect 1660 1056 1668 1064
rect 1724 1056 1732 1064
rect 1548 1016 1556 1024
rect 1644 1016 1652 1024
rect 1404 976 1412 984
rect 1484 976 1492 984
rect 1756 1056 1764 1064
rect 1772 1056 1780 1064
rect 1868 1056 1876 1064
rect 1756 1016 1764 1024
rect 1276 956 1284 964
rect 1356 956 1364 964
rect 1436 956 1444 964
rect 1548 956 1556 964
rect 1612 956 1620 964
rect 1788 1036 1796 1044
rect 1900 1036 1908 1044
rect 2428 1096 2436 1104
rect 2556 1096 2564 1104
rect 2636 1116 2644 1124
rect 2684 1116 2692 1124
rect 3132 1356 3140 1364
rect 3212 1376 3220 1384
rect 3244 1376 3252 1384
rect 3340 1416 3348 1424
rect 3308 1396 3316 1404
rect 3372 1376 3380 1384
rect 3308 1356 3316 1364
rect 3372 1336 3380 1344
rect 3260 1296 3268 1304
rect 3372 1296 3380 1304
rect 2908 1256 2916 1264
rect 2988 1236 2996 1244
rect 2844 1216 2852 1224
rect 2812 1176 2820 1184
rect 2764 1116 2772 1124
rect 2796 1116 2804 1124
rect 2732 1096 2740 1104
rect 2412 1076 2420 1084
rect 2620 1076 2628 1084
rect 2668 1076 2676 1084
rect 2828 1076 2836 1084
rect 2044 1036 2052 1044
rect 2076 1036 2084 1044
rect 2124 1036 2132 1044
rect 2380 1056 2388 1064
rect 2396 1056 2404 1064
rect 2476 1056 2484 1064
rect 2572 1056 2580 1064
rect 2604 1056 2612 1064
rect 2732 1056 2740 1064
rect 764 916 772 924
rect 348 896 356 904
rect 396 896 404 904
rect 668 896 676 904
rect 764 896 772 904
rect 140 816 148 824
rect 284 816 292 824
rect 188 756 196 764
rect 124 736 132 744
rect 252 716 260 724
rect 108 676 116 684
rect 156 676 164 684
rect 108 656 116 664
rect 156 616 164 624
rect 236 676 244 684
rect 716 876 724 884
rect 460 836 468 844
rect 428 776 436 784
rect 364 736 372 744
rect 364 696 372 704
rect 396 696 404 704
rect 364 676 372 684
rect 220 656 228 664
rect 412 656 420 664
rect 444 636 452 644
rect 348 596 356 604
rect 204 576 212 584
rect 284 576 292 584
rect 300 576 308 584
rect 332 576 340 584
rect 508 716 516 724
rect 476 696 484 704
rect 604 676 612 684
rect 524 616 532 624
rect 572 616 580 624
rect 620 616 628 624
rect 860 916 868 924
rect 1020 916 1028 924
rect 1132 916 1140 924
rect 1180 916 1188 924
rect 1308 916 1316 924
rect 972 896 980 904
rect 796 796 804 804
rect 828 796 836 804
rect 668 756 676 764
rect 652 736 660 744
rect 764 716 772 724
rect 700 696 708 704
rect 876 816 884 824
rect 892 776 900 784
rect 940 816 948 824
rect 956 736 964 744
rect 812 696 820 704
rect 844 696 852 704
rect 1260 896 1268 904
rect 1276 896 1284 904
rect 1276 836 1284 844
rect 1100 816 1108 824
rect 1068 756 1076 764
rect 1084 716 1092 724
rect 1052 696 1060 704
rect 1084 696 1092 704
rect 1228 756 1236 764
rect 1116 716 1124 724
rect 1180 716 1188 724
rect 1148 696 1156 704
rect 1244 696 1252 704
rect 1260 696 1268 704
rect 1292 736 1300 744
rect 2140 956 2148 964
rect 1740 936 1748 944
rect 1756 936 1764 944
rect 1804 936 1812 944
rect 1948 936 1956 944
rect 1996 936 2004 944
rect 2028 936 2036 944
rect 2092 936 2100 944
rect 2124 936 2132 944
rect 2188 936 2196 944
rect 2220 936 2228 944
rect 1484 896 1492 904
rect 1404 856 1412 864
rect 1516 856 1524 864
rect 1548 856 1556 864
rect 1580 856 1588 864
rect 1324 696 1332 704
rect 1372 696 1380 704
rect 1436 836 1444 844
rect 1580 836 1588 844
rect 1420 796 1428 804
rect 1580 796 1588 804
rect 1900 916 1908 924
rect 1980 916 1988 924
rect 1996 916 2004 924
rect 2028 916 2036 924
rect 1980 896 1988 904
rect 1692 876 1700 884
rect 1724 876 1732 884
rect 1644 856 1652 864
rect 1596 776 1604 784
rect 1644 776 1652 784
rect 1676 776 1684 784
rect 1484 736 1492 744
rect 1692 756 1700 764
rect 1884 856 1892 864
rect 1772 816 1780 824
rect 1756 776 1764 784
rect 1564 716 1572 724
rect 652 656 660 664
rect 860 656 868 664
rect 972 656 980 664
rect 1452 676 1460 684
rect 1772 736 1780 744
rect 1852 736 1860 744
rect 1612 676 1620 684
rect 1644 676 1652 684
rect 1836 676 1844 684
rect 684 616 692 624
rect 668 596 676 604
rect 316 556 324 564
rect 364 556 372 564
rect 556 556 564 564
rect 604 556 612 564
rect 620 556 628 564
rect 44 536 52 544
rect 92 536 100 544
rect 124 536 132 544
rect 268 536 276 544
rect 396 536 404 544
rect 428 536 436 544
rect 460 536 468 544
rect 492 536 500 544
rect 636 536 644 544
rect 92 516 100 524
rect 588 516 596 524
rect 44 336 52 344
rect 76 336 84 344
rect 60 316 68 324
rect 188 496 196 504
rect 220 496 228 504
rect 284 496 292 504
rect 364 476 372 484
rect 492 476 500 484
rect 636 476 644 484
rect 316 456 324 464
rect 460 456 468 464
rect 124 396 132 404
rect 172 396 180 404
rect 140 376 148 384
rect 108 336 116 344
rect 156 356 164 364
rect 252 416 260 424
rect 236 356 244 364
rect 300 376 308 384
rect 252 336 260 344
rect 188 276 196 284
rect 252 276 260 284
rect 284 276 292 284
rect 364 356 372 364
rect 412 356 420 364
rect 428 336 436 344
rect 572 396 580 404
rect 604 396 612 404
rect 588 336 596 344
rect 716 556 724 564
rect 780 616 788 624
rect 828 596 836 604
rect 924 616 932 624
rect 1004 596 1012 604
rect 860 576 868 584
rect 812 556 820 564
rect 1020 556 1028 564
rect 716 536 724 544
rect 796 536 804 544
rect 844 536 852 544
rect 940 536 948 544
rect 892 496 900 504
rect 940 496 948 504
rect 972 496 980 504
rect 668 476 676 484
rect 652 336 660 344
rect 460 316 468 324
rect 652 316 660 324
rect 508 296 516 304
rect 796 356 804 364
rect 812 336 820 344
rect 1036 476 1044 484
rect 1372 636 1380 644
rect 1532 636 1540 644
rect 1068 556 1076 564
rect 1116 556 1124 564
rect 1164 616 1172 624
rect 1308 616 1316 624
rect 1340 596 1348 604
rect 1372 596 1380 604
rect 1356 556 1364 564
rect 1388 556 1396 564
rect 1420 556 1428 564
rect 1500 596 1508 604
rect 1660 636 1668 644
rect 1836 636 1844 644
rect 1644 596 1652 604
rect 1740 596 1748 604
rect 1484 556 1492 564
rect 1500 556 1508 564
rect 1548 556 1556 564
rect 1580 556 1588 564
rect 1644 556 1652 564
rect 1212 536 1220 544
rect 1324 536 1332 544
rect 1420 536 1428 544
rect 1468 536 1476 544
rect 1836 596 1844 604
rect 1820 556 1828 564
rect 2076 916 2084 924
rect 2348 956 2356 964
rect 2412 956 2420 964
rect 2444 956 2452 964
rect 2652 1036 2660 1044
rect 2716 1036 2724 1044
rect 2604 996 2612 1004
rect 2780 996 2788 1004
rect 2828 996 2836 1004
rect 2732 976 2740 984
rect 2860 1196 2868 1204
rect 3004 1196 3012 1204
rect 2892 1176 2900 1184
rect 2876 1116 2884 1124
rect 2940 1116 2948 1124
rect 2988 1116 2996 1124
rect 2956 1096 2964 1104
rect 2876 1056 2884 1064
rect 2924 1056 2932 1064
rect 2972 1056 2980 1064
rect 2988 1036 2996 1044
rect 2940 996 2948 1004
rect 2956 996 2964 1004
rect 2972 996 2980 1004
rect 2908 976 2916 984
rect 2972 976 2980 984
rect 2668 956 2676 964
rect 3004 996 3012 1004
rect 3164 1256 3172 1264
rect 3388 1236 3396 1244
rect 3164 1176 3172 1184
rect 3084 1116 3092 1124
rect 3132 1116 3140 1124
rect 3084 1076 3092 1084
rect 3068 1056 3076 1064
rect 3100 1056 3108 1064
rect 3036 976 3044 984
rect 3084 976 3092 984
rect 2300 936 2308 944
rect 2316 936 2324 944
rect 2364 936 2372 944
rect 2460 936 2468 944
rect 2620 936 2628 944
rect 2812 936 2820 944
rect 2844 936 2852 944
rect 2860 936 2868 944
rect 2188 916 2196 924
rect 2252 916 2260 924
rect 2284 916 2292 924
rect 2332 916 2340 924
rect 2428 916 2436 924
rect 2028 896 2036 904
rect 2572 896 2580 904
rect 2652 896 2660 904
rect 2684 896 2692 904
rect 2092 876 2100 884
rect 2172 876 2180 884
rect 1932 756 1940 764
rect 1884 736 1892 744
rect 1932 736 1940 744
rect 1948 736 1956 744
rect 1900 696 1908 704
rect 1980 696 1988 704
rect 2348 836 2356 844
rect 2108 736 2116 744
rect 2188 736 2196 744
rect 2204 736 2212 744
rect 2236 736 2244 744
rect 2124 716 2132 724
rect 2156 716 2164 724
rect 2140 696 2148 704
rect 1884 676 1892 684
rect 1964 676 1972 684
rect 2028 676 2036 684
rect 2188 676 2196 684
rect 2524 816 2532 824
rect 2380 796 2388 804
rect 2316 756 2324 764
rect 2300 736 2308 744
rect 2364 736 2372 744
rect 2428 736 2436 744
rect 2476 736 2484 744
rect 2380 716 2388 724
rect 1980 656 1988 664
rect 2012 656 2020 664
rect 2060 656 2068 664
rect 2236 656 2244 664
rect 2284 656 2292 664
rect 2332 656 2340 664
rect 2348 656 2356 664
rect 1916 636 1924 644
rect 1916 616 1924 624
rect 1948 596 1956 604
rect 2012 576 2020 584
rect 1900 556 1908 564
rect 1916 556 1924 564
rect 1996 556 2004 564
rect 1532 536 1540 544
rect 1788 536 1796 544
rect 1852 536 1860 544
rect 1548 516 1556 524
rect 1596 496 1604 504
rect 1068 476 1076 484
rect 1068 456 1076 464
rect 1084 456 1092 464
rect 988 436 996 444
rect 1052 436 1060 444
rect 956 316 964 324
rect 332 276 340 284
rect 700 276 708 284
rect 732 276 740 284
rect 844 276 852 284
rect 220 256 228 264
rect 396 256 404 264
rect 620 256 628 264
rect 44 156 52 164
rect 92 156 100 164
rect 268 216 276 224
rect 172 176 180 184
rect 204 176 212 184
rect 428 216 436 224
rect 492 196 500 204
rect 524 196 532 204
rect 380 176 388 184
rect 156 156 164 164
rect 428 156 436 164
rect 556 156 564 164
rect 92 136 100 144
rect 140 136 148 144
rect 300 136 308 144
rect 540 116 548 124
rect 556 116 564 124
rect 44 96 52 104
rect 76 96 84 104
rect 124 96 132 104
rect 396 96 404 104
rect 780 256 788 264
rect 860 256 868 264
rect 924 256 932 264
rect 940 256 948 264
rect 1196 396 1204 404
rect 1852 516 1860 524
rect 1868 516 1876 524
rect 1932 516 1940 524
rect 1404 476 1412 484
rect 1436 476 1444 484
rect 1532 476 1540 484
rect 1628 476 1636 484
rect 1356 416 1364 424
rect 1388 396 1396 404
rect 1452 396 1460 404
rect 1036 376 1044 384
rect 1292 376 1300 384
rect 1004 336 1012 344
rect 1132 336 1140 344
rect 1228 336 1236 344
rect 1164 316 1172 324
rect 1260 316 1268 324
rect 1468 356 1476 364
rect 1436 316 1444 324
rect 1180 276 1188 284
rect 1660 396 1668 404
rect 1532 336 1540 344
rect 1660 336 1668 344
rect 1484 296 1492 304
rect 1596 296 1604 304
rect 1612 296 1620 304
rect 1644 296 1652 304
rect 1308 256 1316 264
rect 1324 256 1332 264
rect 1372 256 1380 264
rect 1500 256 1508 264
rect 620 176 628 184
rect 732 176 740 184
rect 636 156 644 164
rect 636 136 644 144
rect 780 136 788 144
rect 1004 216 1012 224
rect 1084 216 1092 224
rect 908 156 916 164
rect 940 156 948 164
rect 1196 216 1204 224
rect 1436 236 1444 244
rect 1388 216 1396 224
rect 1372 196 1380 204
rect 876 136 884 144
rect 828 116 836 124
rect 1100 136 1108 144
rect 1148 136 1156 144
rect 1196 136 1204 144
rect 1724 396 1732 404
rect 1740 376 1748 384
rect 1724 356 1732 364
rect 1804 336 1812 344
rect 1692 316 1700 324
rect 1676 296 1684 304
rect 2076 556 2084 564
rect 2156 556 2164 564
rect 2220 576 2228 584
rect 2268 636 2276 644
rect 2300 616 2308 624
rect 2284 576 2292 584
rect 2300 576 2308 584
rect 2572 756 2580 764
rect 2636 756 2644 764
rect 2540 736 2548 744
rect 2556 736 2564 744
rect 2620 736 2628 744
rect 2460 716 2468 724
rect 2828 876 2836 884
rect 2972 916 2980 924
rect 2940 896 2948 904
rect 3292 1156 3300 1164
rect 3180 1096 3188 1104
rect 3132 1076 3140 1084
rect 3436 1416 3444 1424
rect 3468 1416 3476 1424
rect 3404 1216 3412 1224
rect 3532 1396 3540 1404
rect 3548 1396 3556 1404
rect 3660 1456 3668 1464
rect 3628 1436 3636 1444
rect 3708 1436 3716 1444
rect 3596 1416 3604 1424
rect 3660 1416 3668 1424
rect 4108 1596 4116 1604
rect 4124 1576 4132 1584
rect 4060 1516 4068 1524
rect 4092 1516 4100 1524
rect 4188 1616 4196 1624
rect 4156 1596 4164 1604
rect 4220 1576 4228 1584
rect 4172 1516 4180 1524
rect 4220 1516 4228 1524
rect 4252 1516 4260 1524
rect 4140 1496 4148 1504
rect 3756 1476 3764 1484
rect 3996 1476 4004 1484
rect 3756 1456 3764 1464
rect 3932 1456 3940 1464
rect 3964 1456 3972 1464
rect 4060 1456 4068 1464
rect 4092 1456 4100 1464
rect 3676 1376 3684 1384
rect 4028 1436 4036 1444
rect 4076 1436 4084 1444
rect 3948 1416 3956 1424
rect 3852 1376 3860 1384
rect 3868 1376 3876 1384
rect 3980 1376 3988 1384
rect 4044 1376 4052 1384
rect 3756 1356 3764 1364
rect 3820 1336 3828 1344
rect 3612 1316 3620 1324
rect 4108 1416 4116 1424
rect 4092 1376 4100 1384
rect 3884 1356 3892 1364
rect 3964 1356 3972 1364
rect 4124 1356 4132 1364
rect 4188 1456 4196 1464
rect 4220 1456 4228 1464
rect 4156 1436 4164 1444
rect 4204 1356 4212 1364
rect 3452 1296 3460 1304
rect 3468 1296 3476 1304
rect 3788 1296 3796 1304
rect 3900 1296 3908 1304
rect 3452 1276 3460 1284
rect 3580 1276 3588 1284
rect 3436 1236 3444 1244
rect 3516 1216 3524 1224
rect 3644 1216 3652 1224
rect 3356 1176 3364 1184
rect 3372 1156 3380 1164
rect 3452 1156 3460 1164
rect 3484 1136 3492 1144
rect 3404 1116 3412 1124
rect 3436 1116 3444 1124
rect 3324 1096 3332 1104
rect 3532 1196 3540 1204
rect 3612 1156 3620 1164
rect 3564 1096 3572 1104
rect 3948 1296 3956 1304
rect 3996 1296 4004 1304
rect 3756 1256 3764 1264
rect 3916 1256 3924 1264
rect 3708 1236 3716 1244
rect 3660 1176 3668 1184
rect 3788 1236 3796 1244
rect 3724 1176 3732 1184
rect 3852 1156 3860 1164
rect 3900 1136 3908 1144
rect 3948 1136 3956 1144
rect 4044 1136 4052 1144
rect 3644 1096 3652 1104
rect 3516 1076 3524 1084
rect 3548 1076 3556 1084
rect 3676 1076 3684 1084
rect 3692 1076 3700 1084
rect 3244 1056 3252 1064
rect 3276 1056 3284 1064
rect 3308 1056 3316 1064
rect 3148 1036 3156 1044
rect 3212 1036 3220 1044
rect 3148 996 3156 1004
rect 3228 976 3236 984
rect 3196 956 3204 964
rect 3484 1036 3492 1044
rect 3580 1036 3588 1044
rect 3436 996 3444 1004
rect 3468 996 3476 1004
rect 3724 1036 3732 1044
rect 3324 976 3332 984
rect 3452 976 3460 984
rect 3244 956 3252 964
rect 3308 956 3316 964
rect 3356 956 3364 964
rect 3452 956 3460 964
rect 3644 976 3652 984
rect 3516 956 3524 964
rect 3628 956 3636 964
rect 3644 956 3652 964
rect 3276 936 3284 944
rect 3868 1096 3876 1104
rect 3996 1116 4004 1124
rect 3964 1096 3972 1104
rect 3820 1076 3828 1084
rect 3852 1076 3860 1084
rect 3916 1076 3924 1084
rect 4012 1076 4020 1084
rect 4108 1076 4116 1084
rect 3772 1036 3780 1044
rect 3740 1016 3748 1024
rect 3996 1036 4004 1044
rect 4076 1036 4084 1044
rect 3836 996 3844 1004
rect 3868 956 3876 964
rect 3772 936 3780 944
rect 3804 936 3812 944
rect 3852 936 3860 944
rect 3884 936 3892 944
rect 3356 916 3364 924
rect 3372 916 3380 924
rect 3468 916 3476 924
rect 3020 896 3028 904
rect 3116 896 3124 904
rect 3196 896 3204 904
rect 3420 896 3428 904
rect 2892 836 2900 844
rect 2748 796 2756 804
rect 2844 796 2852 804
rect 3420 876 3428 884
rect 3452 876 3460 884
rect 3180 856 3188 864
rect 3244 836 3252 844
rect 3308 816 3316 824
rect 3164 796 3172 804
rect 3244 796 3252 804
rect 3404 796 3412 804
rect 2908 756 2916 764
rect 3228 756 3236 764
rect 2668 736 2676 744
rect 2764 716 2772 724
rect 2876 696 2884 704
rect 3276 736 3284 744
rect 2988 716 2996 724
rect 3020 716 3028 724
rect 3052 716 3060 724
rect 2924 696 2932 704
rect 2556 656 2564 664
rect 2716 676 2724 684
rect 2828 676 2836 684
rect 2940 676 2948 684
rect 2460 636 2468 644
rect 2444 616 2452 624
rect 2380 596 2388 604
rect 2412 596 2420 604
rect 2428 556 2436 564
rect 2268 536 2276 544
rect 2028 436 2036 444
rect 1964 336 1972 344
rect 1996 316 2004 324
rect 1916 296 1924 304
rect 1692 256 1700 264
rect 1964 256 1972 264
rect 1596 236 1604 244
rect 1628 236 1636 244
rect 1532 216 1540 224
rect 1548 196 1556 204
rect 1580 196 1588 204
rect 1516 176 1524 184
rect 908 96 916 104
rect 1020 96 1028 104
rect 1052 96 1060 104
rect 1116 96 1124 104
rect 1164 96 1172 104
rect 1212 96 1220 104
rect 1276 116 1284 124
rect 1628 216 1636 224
rect 1612 176 1620 184
rect 1644 196 1652 204
rect 1596 136 1604 144
rect 1772 236 1780 244
rect 1852 236 1860 244
rect 1884 216 1892 224
rect 1932 216 1940 224
rect 1884 196 1892 204
rect 1900 196 1908 204
rect 1660 176 1668 184
rect 1708 176 1716 184
rect 1772 176 1780 184
rect 1820 176 1828 184
rect 1836 176 1844 184
rect 1868 176 1876 184
rect 1932 176 1940 184
rect 2044 356 2052 364
rect 2124 496 2132 504
rect 2236 496 2244 504
rect 2124 476 2132 484
rect 2204 476 2212 484
rect 2092 456 2100 464
rect 2156 376 2164 384
rect 2092 336 2100 344
rect 2076 296 2084 304
rect 2092 296 2100 304
rect 2204 336 2212 344
rect 2220 336 2228 344
rect 2236 316 2244 324
rect 2348 516 2356 524
rect 2428 496 2436 504
rect 2476 496 2484 504
rect 2284 476 2292 484
rect 2348 476 2356 484
rect 2284 416 2292 424
rect 2332 416 2340 424
rect 2364 396 2372 404
rect 2348 356 2356 364
rect 2172 296 2180 304
rect 2204 296 2212 304
rect 2268 296 2276 304
rect 2508 556 2516 564
rect 2524 556 2532 564
rect 2604 636 2612 644
rect 2684 636 2692 644
rect 2524 536 2532 544
rect 2588 536 2596 544
rect 2556 516 2564 524
rect 2876 636 2884 644
rect 2876 616 2884 624
rect 2732 596 2740 604
rect 2860 596 2868 604
rect 2892 596 2900 604
rect 2844 576 2852 584
rect 2684 556 2692 564
rect 2748 556 2756 564
rect 2796 556 2804 564
rect 2668 536 2676 544
rect 2780 536 2788 544
rect 2812 536 2820 544
rect 2876 536 2884 544
rect 2684 516 2692 524
rect 2764 516 2772 524
rect 2844 516 2852 524
rect 2892 516 2900 524
rect 2876 496 2884 504
rect 2492 436 2500 444
rect 2620 396 2628 404
rect 2540 336 2548 344
rect 2572 336 2580 344
rect 3100 636 3108 644
rect 3020 616 3028 624
rect 3084 616 3092 624
rect 2956 576 2964 584
rect 3148 696 3156 704
rect 3132 676 3140 684
rect 3308 676 3316 684
rect 3196 616 3204 624
rect 3036 576 3044 584
rect 3340 636 3348 644
rect 3436 756 3444 764
rect 3452 736 3460 744
rect 3948 976 3956 984
rect 3996 976 4004 984
rect 4044 976 4052 984
rect 4236 1336 4244 1344
rect 4156 1316 4164 1324
rect 4252 1196 4260 1204
rect 4188 1156 4196 1164
rect 4220 1116 4228 1124
rect 4172 1076 4180 1084
rect 4188 1056 4196 1064
rect 4156 1036 4164 1044
rect 4124 1016 4132 1024
rect 4172 996 4180 1004
rect 4204 996 4212 1004
rect 4156 976 4164 984
rect 4204 976 4212 984
rect 4236 976 4244 984
rect 3916 956 3924 964
rect 3980 956 3988 964
rect 4108 956 4116 964
rect 4028 936 4036 944
rect 4060 936 4068 944
rect 4092 936 4100 944
rect 4124 936 4132 944
rect 3788 916 3796 924
rect 3820 916 3828 924
rect 3900 916 3908 924
rect 3916 916 3924 924
rect 4060 916 4068 924
rect 4108 916 4116 924
rect 3596 896 3604 904
rect 3628 896 3636 904
rect 3692 896 3700 904
rect 3500 876 3508 884
rect 3532 876 3540 884
rect 3548 876 3556 884
rect 3628 876 3636 884
rect 3564 816 3572 824
rect 3500 736 3508 744
rect 3740 876 3748 884
rect 3660 836 3668 844
rect 3628 696 3636 704
rect 3900 896 3908 904
rect 4028 896 4036 904
rect 3916 816 3924 824
rect 3964 816 3972 824
rect 4076 836 4084 844
rect 4028 776 4036 784
rect 4108 756 4116 764
rect 3868 716 3876 724
rect 3948 716 3956 724
rect 4140 716 4148 724
rect 4188 716 4196 724
rect 3820 696 3828 704
rect 3468 676 3476 684
rect 3628 676 3636 684
rect 3676 676 3684 684
rect 3740 676 3748 684
rect 3820 676 3828 684
rect 4108 676 4116 684
rect 4156 676 4164 684
rect 3516 656 3524 664
rect 3548 656 3556 664
rect 3580 656 3588 664
rect 3676 656 3684 664
rect 3740 656 3748 664
rect 3772 656 3780 664
rect 3852 656 3860 664
rect 3404 636 3412 644
rect 3372 616 3380 624
rect 3324 596 3332 604
rect 3260 576 3268 584
rect 3308 576 3316 584
rect 3324 576 3332 584
rect 3372 576 3380 584
rect 3116 556 3124 564
rect 2972 536 2980 544
rect 3004 536 3012 544
rect 3052 536 3060 544
rect 2972 516 2980 524
rect 3020 496 3028 504
rect 3004 476 3012 484
rect 2652 396 2660 404
rect 2844 396 2852 404
rect 2940 396 2948 404
rect 2732 376 2740 384
rect 2684 356 2692 364
rect 2892 336 2900 344
rect 2940 336 2948 344
rect 2764 316 2772 324
rect 2988 316 2996 324
rect 2860 296 2868 304
rect 3148 496 3156 504
rect 3116 476 3124 484
rect 3356 556 3364 564
rect 3404 556 3412 564
rect 3484 556 3492 564
rect 3596 616 3604 624
rect 3884 636 3892 644
rect 3708 616 3716 624
rect 3580 556 3588 564
rect 3660 556 3668 564
rect 3580 536 3588 544
rect 3628 536 3636 544
rect 3676 536 3684 544
rect 4076 656 4084 664
rect 4108 656 4116 664
rect 3916 576 3924 584
rect 3852 556 3860 564
rect 3884 556 3892 564
rect 3948 596 3956 604
rect 4028 596 4036 604
rect 3964 576 3972 584
rect 3756 536 3764 544
rect 3788 536 3796 544
rect 3836 536 3844 544
rect 3932 536 3940 544
rect 4028 536 4036 544
rect 4060 536 4068 544
rect 4124 536 4132 544
rect 3404 516 3412 524
rect 3468 516 3476 524
rect 3500 516 3508 524
rect 3564 516 3572 524
rect 3356 496 3364 504
rect 3244 456 3252 464
rect 3276 456 3284 464
rect 3308 456 3316 464
rect 3308 396 3316 404
rect 3100 376 3108 384
rect 3148 376 3156 384
rect 3068 356 3076 364
rect 3036 336 3044 344
rect 3116 336 3124 344
rect 3084 316 3092 324
rect 3180 316 3188 324
rect 3212 316 3220 324
rect 3244 316 3252 324
rect 3292 316 3300 324
rect 2764 276 2772 284
rect 2812 276 2820 284
rect 2908 276 2916 284
rect 2940 276 2948 284
rect 2972 276 2980 284
rect 3260 276 3268 284
rect 2044 256 2052 264
rect 2428 256 2436 264
rect 2444 256 2452 264
rect 2652 256 2660 264
rect 3132 256 3140 264
rect 3164 256 3172 264
rect 3292 256 3300 264
rect 2092 236 2100 244
rect 2172 236 2180 244
rect 2380 236 2388 244
rect 2604 236 2612 244
rect 2428 216 2436 224
rect 2252 196 2260 204
rect 2044 176 2052 184
rect 2092 176 2100 184
rect 2124 176 2132 184
rect 2156 176 2164 184
rect 2460 156 2468 164
rect 2524 156 2532 164
rect 1804 136 1812 144
rect 1836 136 1844 144
rect 1916 136 1924 144
rect 1948 136 1956 144
rect 1964 136 1972 144
rect 2108 136 2116 144
rect 2300 136 2308 144
rect 2556 136 2564 144
rect 1724 116 1732 124
rect 2556 116 2564 124
rect 1564 96 1572 104
rect 1756 96 1764 104
rect 1916 96 1924 104
rect 1996 96 2004 104
rect 2204 96 2212 104
rect 2252 96 2260 104
rect 2364 96 2372 104
rect 812 76 820 84
rect 892 76 900 84
rect 1180 76 1188 84
rect 1244 76 1252 84
rect 1468 76 1476 84
rect 1532 76 1540 84
rect 1772 76 1780 84
rect 1804 76 1812 84
rect 1948 76 1956 84
rect 2012 76 2020 84
rect 2156 76 2164 84
rect 2476 76 2484 84
rect 2684 196 2692 204
rect 2636 176 2644 184
rect 2700 176 2708 184
rect 2588 156 2596 164
rect 2764 216 2772 224
rect 2748 176 2756 184
rect 2876 216 2884 224
rect 2940 216 2948 224
rect 2828 196 2836 204
rect 2844 156 2852 164
rect 2908 156 2916 164
rect 2956 156 2964 164
rect 2924 116 2932 124
rect 2940 116 2948 124
rect 3004 216 3012 224
rect 3036 196 3044 204
rect 3036 136 3044 144
rect 3068 136 3076 144
rect 3004 116 3012 124
rect 3116 196 3124 204
rect 3212 196 3220 204
rect 3260 176 3268 184
rect 3148 136 3156 144
rect 3180 136 3188 144
rect 3340 316 3348 324
rect 3372 476 3380 484
rect 3516 416 3524 424
rect 3452 376 3460 384
rect 3388 356 3396 364
rect 3404 356 3412 364
rect 3500 356 3508 364
rect 3436 316 3444 324
rect 3708 516 3716 524
rect 3724 516 3732 524
rect 3740 516 3748 524
rect 3756 516 3764 524
rect 3836 516 3844 524
rect 3852 516 3860 524
rect 4108 516 4116 524
rect 3852 476 3860 484
rect 3740 436 3748 444
rect 3772 436 3780 444
rect 3612 396 3620 404
rect 3692 396 3700 404
rect 3612 356 3620 364
rect 3868 376 3876 384
rect 3772 336 3780 344
rect 3820 336 3828 344
rect 3564 316 3572 324
rect 3580 316 3588 324
rect 3644 316 3652 324
rect 3708 316 3716 324
rect 3772 316 3780 324
rect 3724 296 3732 304
rect 3804 296 3812 304
rect 3852 296 3860 304
rect 4076 496 4084 504
rect 3964 476 3972 484
rect 4012 476 4020 484
rect 4108 416 4116 424
rect 4188 416 4196 424
rect 4236 396 4244 404
rect 3980 316 3988 324
rect 3916 296 3924 304
rect 3468 256 3476 264
rect 3532 256 3540 264
rect 3596 256 3604 264
rect 3676 256 3684 264
rect 3932 256 3940 264
rect 4012 256 4020 264
rect 3324 236 3332 244
rect 3388 236 3396 244
rect 3484 236 3492 244
rect 3548 236 3556 244
rect 3356 176 3364 184
rect 3532 216 3540 224
rect 3372 136 3380 144
rect 3644 236 3652 244
rect 3724 236 3732 244
rect 3596 196 3604 204
rect 3580 176 3588 184
rect 3452 156 3460 164
rect 3516 156 3524 164
rect 3404 116 3412 124
rect 2764 96 2772 104
rect 2796 96 2804 104
rect 2956 96 2964 104
rect 2988 96 2996 104
rect 3036 96 3044 104
rect 3164 96 3172 104
rect 3100 76 3108 84
rect 3740 216 3748 224
rect 3804 216 3812 224
rect 3772 196 3780 204
rect 3612 176 3620 184
rect 3756 176 3764 184
rect 4220 296 4228 304
rect 4124 276 4132 284
rect 4140 256 4148 264
rect 4092 236 4100 244
rect 3932 216 3940 224
rect 4012 196 4020 204
rect 4028 196 4036 204
rect 3788 156 3796 164
rect 3820 156 3828 164
rect 3868 156 3876 164
rect 3948 156 3956 164
rect 4188 216 4196 224
rect 4108 196 4116 204
rect 4268 196 4276 204
rect 4124 176 4132 184
rect 4204 176 4212 184
rect 4172 156 4180 164
rect 4188 156 4196 164
rect 3468 136 3476 144
rect 3692 136 3700 144
rect 3804 136 3812 144
rect 3836 136 3844 144
rect 4044 136 4052 144
rect 3452 116 3460 124
rect 3484 116 3492 124
rect 3676 116 3684 124
rect 4012 116 4020 124
rect 4076 116 4084 124
rect 4092 116 4100 124
rect 4188 116 4196 124
rect 3548 96 3556 104
rect 3820 96 3828 104
rect 3852 96 3860 104
rect 4140 96 4148 104
rect 4236 96 4244 104
rect 3052 56 3060 64
rect 3420 56 3428 64
rect 2876 16 2884 24
<< metal3 >>
rect 2644 2997 2732 3003
rect 2804 2997 3388 3003
rect 228 2977 428 2983
rect 452 2977 508 2983
rect 532 2977 732 2983
rect 868 2977 1692 2983
rect 1764 2977 1859 2983
rect -51 2957 12 2963
rect 20 2957 156 2963
rect 164 2957 380 2963
rect 388 2957 604 2963
rect 628 2957 700 2963
rect 884 2957 972 2963
rect 1108 2957 1164 2963
rect 1380 2957 1388 2963
rect 1405 2957 1420 2963
rect 1444 2957 1516 2963
rect 1540 2957 1596 2963
rect 1709 2963 1715 2976
rect 1709 2957 1724 2963
rect 1748 2957 1772 2963
rect 1853 2963 1859 2977
rect 2004 2977 2972 2983
rect 2996 2977 3004 2983
rect 3172 2977 3612 2983
rect 3844 2977 3996 2983
rect 1853 2957 2012 2963
rect 2132 2957 2156 2963
rect 2228 2957 2364 2963
rect 2532 2957 2572 2963
rect 2676 2957 2764 2963
rect 2788 2957 2796 2963
rect 2852 2957 3164 2963
rect 3172 2957 3468 2963
rect 3533 2957 3548 2963
rect 3572 2957 3603 2963
rect 1837 2944 1843 2956
rect 148 2937 220 2943
rect 228 2937 284 2943
rect 292 2937 412 2943
rect 420 2937 460 2943
rect 532 2937 764 2943
rect 852 2937 1148 2943
rect 1156 2937 1244 2943
rect 1508 2937 1516 2943
rect 1588 2937 1692 2943
rect 1844 2937 2844 2943
rect 2884 2937 2892 2943
rect 2916 2937 2924 2943
rect 2964 2937 2972 2943
rect 2996 2937 3084 2943
rect 3236 2937 3244 2943
rect 3268 2937 3276 2943
rect 3380 2937 3580 2943
rect 3597 2943 3603 2957
rect 3620 2957 3708 2963
rect 3956 2957 4060 2963
rect 4141 2957 4156 2963
rect 4141 2944 4147 2957
rect 3597 2937 3628 2943
rect 3213 2924 3219 2936
rect 3661 2924 3667 2936
rect 3677 2924 3683 2943
rect 468 2917 492 2923
rect 740 2917 764 2923
rect 772 2917 1676 2923
rect 1684 2917 2252 2923
rect 2340 2917 2348 2923
rect 2404 2917 2412 2923
rect 2436 2917 2940 2923
rect 3124 2917 3148 2923
rect 3252 2917 3276 2923
rect 3508 2917 3532 2923
rect 3716 2917 3740 2923
rect 100 2897 124 2903
rect 260 2897 332 2903
rect 484 2897 572 2903
rect 660 2897 668 2903
rect 916 2897 972 2903
rect 1012 2897 1116 2903
rect 1476 2897 2460 2903
rect 2468 2897 2476 2903
rect 2532 2897 2604 2903
rect 2692 2897 2700 2903
rect 2932 2897 3068 2903
rect 3076 2897 3644 2903
rect 3652 2897 3836 2903
rect 3844 2897 3868 2903
rect 3892 2897 3964 2903
rect 3972 2897 3980 2903
rect 4077 2884 4083 2896
rect 692 2877 1052 2883
rect 1524 2877 1548 2883
rect 1572 2877 1612 2883
rect 1636 2877 1804 2883
rect 1892 2877 1996 2883
rect 2068 2877 2076 2883
rect 2100 2877 2812 2883
rect 3140 2877 3180 2883
rect 3732 2877 3756 2883
rect 1044 2857 1276 2863
rect 1533 2844 1539 2856
rect 1917 2844 1923 2863
rect 2020 2857 2092 2863
rect 2116 2857 2124 2863
rect 2308 2857 2316 2863
rect 2404 2857 2444 2863
rect 2564 2857 2572 2863
rect 3508 2857 3948 2863
rect 1204 2837 1388 2843
rect 2484 2837 3132 2843
rect 1348 2817 1420 2823
rect 3748 2817 3932 2823
rect 340 2797 364 2803
rect 372 2797 508 2803
rect 516 2797 524 2803
rect 932 2797 956 2803
rect 1028 2797 1036 2803
rect 1188 2797 1228 2803
rect 1604 2797 1788 2803
rect 2148 2797 2220 2803
rect 2276 2797 2300 2803
rect 2644 2797 2652 2803
rect 2900 2797 3036 2803
rect 3044 2797 3340 2803
rect 3348 2797 4108 2803
rect 4116 2797 4124 2803
rect 660 2777 1468 2783
rect 2052 2777 2092 2783
rect 3892 2777 4060 2783
rect 532 2757 844 2763
rect 1300 2757 1452 2763
rect 2324 2757 2412 2763
rect 3780 2757 3836 2763
rect 4052 2757 4156 2763
rect 100 2737 124 2743
rect 132 2737 156 2743
rect 164 2737 284 2743
rect 500 2737 620 2743
rect 628 2737 748 2743
rect 756 2737 812 2743
rect 1028 2737 1100 2743
rect 1524 2737 1708 2743
rect 2084 2737 2092 2743
rect 2340 2737 2444 2743
rect 2532 2737 2796 2743
rect 3028 2737 3132 2743
rect 3332 2737 3676 2743
rect 3988 2737 4092 2743
rect 4100 2737 4108 2743
rect 132 2717 412 2723
rect 420 2717 716 2723
rect 724 2717 764 2723
rect 948 2717 956 2723
rect 964 2717 1356 2723
rect 1492 2717 1532 2723
rect 1972 2717 2108 2723
rect 2148 2717 2156 2723
rect 2468 2717 2524 2723
rect 2644 2717 2652 2723
rect 2772 2717 2780 2723
rect 2820 2717 2876 2723
rect 3012 2717 3228 2723
rect 3476 2717 3516 2723
rect 3556 2717 3564 2723
rect 3572 2717 3580 2723
rect 3604 2717 3612 2723
rect 3668 2717 3724 2723
rect 3764 2717 3852 2723
rect 3876 2717 3900 2723
rect 109 2697 236 2703
rect 68 2677 76 2683
rect 109 2683 115 2697
rect 388 2697 492 2703
rect 596 2697 668 2703
rect 708 2697 796 2703
rect 804 2697 876 2703
rect 1236 2697 1260 2703
rect 1412 2697 1788 2703
rect 1796 2697 2508 2703
rect 2516 2697 3148 2703
rect 3156 2697 3628 2703
rect 3636 2697 3676 2703
rect 3684 2697 3820 2703
rect 84 2677 115 2683
rect 180 2677 252 2683
rect 388 2677 540 2683
rect 836 2677 924 2683
rect 1028 2677 1244 2683
rect 1444 2677 2076 2683
rect 2100 2677 2108 2683
rect 2132 2677 2172 2683
rect 2212 2677 2252 2683
rect 2260 2677 3068 2683
rect 3140 2677 3548 2683
rect 3556 2677 3580 2683
rect 3604 2677 3644 2683
rect 3940 2677 3948 2683
rect 3981 2664 3987 2676
rect 20 2657 172 2663
rect 532 2657 636 2663
rect 884 2657 972 2663
rect 1076 2657 1164 2663
rect 1284 2657 1292 2663
rect 1540 2657 1548 2663
rect 1572 2657 1820 2663
rect 1844 2657 1900 2663
rect 1917 2657 1932 2663
rect 1469 2644 1475 2656
rect 1917 2644 1923 2657
rect 2084 2657 2172 2663
rect 2196 2657 2348 2663
rect 2436 2657 2444 2663
rect 2516 2657 2524 2663
rect 2548 2657 2572 2663
rect 2628 2657 2636 2663
rect 2692 2657 2700 2663
rect 2740 2657 2748 2663
rect 2772 2657 3404 2663
rect 3732 2657 3820 2663
rect 4116 2657 4140 2663
rect 52 2637 92 2643
rect 772 2637 940 2643
rect 957 2637 972 2643
rect 996 2637 1196 2643
rect 1732 2637 1756 2643
rect 1780 2637 1852 2643
rect 1940 2637 2044 2643
rect 2116 2637 2268 2643
rect 2404 2637 2460 2643
rect 2468 2637 3132 2643
rect 3268 2637 3276 2643
rect 948 2617 1004 2623
rect 1124 2617 1260 2623
rect 1828 2617 1868 2623
rect 1908 2617 1980 2623
rect 2004 2617 2028 2623
rect 2116 2617 2124 2623
rect 2948 2617 2956 2623
rect 3156 2617 3164 2623
rect 3476 2617 3980 2623
rect 3053 2604 3059 2616
rect 356 2597 364 2603
rect 804 2597 860 2603
rect 868 2597 1324 2603
rect 1668 2597 1740 2603
rect 1812 2597 1852 2603
rect 1892 2597 2156 2603
rect 2324 2597 2636 2603
rect 2724 2597 2924 2603
rect 3076 2597 3084 2603
rect 3188 2597 3260 2603
rect 3396 2597 3436 2603
rect 3524 2597 3532 2603
rect 3556 2597 3884 2603
rect 4164 2597 4188 2603
rect 84 2577 364 2583
rect 404 2577 636 2583
rect 692 2577 780 2583
rect 1268 2577 1388 2583
rect 1492 2577 1836 2583
rect 1844 2577 1932 2583
rect 1940 2577 2060 2583
rect 2084 2577 2764 2583
rect 2781 2577 2796 2583
rect 2900 2577 2908 2583
rect 2980 2577 3004 2583
rect 3028 2577 3484 2583
rect 3492 2577 3708 2583
rect 3812 2577 3820 2583
rect 3908 2577 3964 2583
rect 4052 2577 4092 2583
rect 1245 2564 1251 2576
rect 180 2557 284 2563
rect 308 2557 444 2563
rect 676 2557 844 2563
rect 1284 2557 1324 2563
rect 1364 2557 1420 2563
rect 1476 2557 1484 2563
rect 1508 2557 1548 2563
rect 1588 2557 1628 2563
rect 1700 2557 1724 2563
rect 1812 2557 2300 2563
rect 2308 2557 3212 2563
rect 3220 2557 3964 2563
rect 3972 2557 4188 2563
rect 164 2537 252 2543
rect 276 2537 348 2543
rect 356 2537 668 2543
rect 676 2537 732 2543
rect 740 2537 844 2543
rect 900 2537 908 2543
rect 916 2537 1020 2543
rect 1028 2537 1052 2543
rect 1076 2537 1116 2543
rect 1124 2537 1788 2543
rect 1901 2524 1907 2543
rect 1924 2537 1996 2543
rect 2020 2537 2028 2543
rect 2100 2537 2764 2543
rect 2884 2537 2924 2543
rect 2948 2537 2972 2543
rect 2996 2537 3004 2543
rect 3076 2537 3308 2543
rect 3348 2537 3356 2543
rect 3412 2537 3436 2543
rect 3460 2537 3468 2543
rect 3508 2537 3523 2543
rect 3556 2537 3564 2543
rect 3636 2537 3660 2543
rect 3684 2537 3756 2543
rect 3780 2537 3868 2543
rect 3908 2537 3916 2543
rect 4052 2537 4060 2543
rect 2093 2524 2099 2536
rect 4173 2524 4179 2536
rect 516 2517 540 2523
rect 548 2517 700 2523
rect 996 2517 1804 2523
rect 1972 2517 1996 2523
rect 2196 2517 2284 2523
rect 2292 2517 2348 2523
rect 2484 2517 2492 2523
rect 2580 2517 2588 2523
rect 2612 2517 2620 2523
rect 2692 2517 2716 2523
rect 2836 2517 3852 2523
rect 125 2504 131 2516
rect 893 2504 899 2516
rect -51 2497 44 2503
rect 52 2497 60 2503
rect 68 2497 92 2503
rect 132 2497 316 2503
rect 324 2497 396 2503
rect 500 2497 540 2503
rect 1364 2497 1372 2503
rect 1412 2497 1420 2503
rect 1444 2497 1468 2503
rect 1524 2497 1580 2503
rect 1588 2497 1676 2503
rect 1748 2497 1756 2503
rect 1796 2497 2236 2503
rect 2244 2497 2252 2503
rect 2324 2497 2364 2503
rect 2564 2497 2700 2503
rect 2708 2497 2716 2503
rect 2868 2497 3036 2503
rect 3060 2497 3084 2503
rect 3092 2497 3196 2503
rect 3204 2497 3500 2503
rect 3524 2497 3532 2503
rect 3604 2497 3612 2503
rect 3636 2497 3644 2503
rect 3828 2497 3836 2503
rect 4148 2497 4220 2503
rect 989 2484 995 2496
rect 3693 2484 3699 2496
rect 372 2477 588 2483
rect 996 2477 1500 2483
rect 1508 2477 1660 2483
rect 1812 2477 1868 2483
rect 2068 2477 2076 2483
rect 2164 2477 2172 2483
rect 2580 2477 3436 2483
rect 644 2457 652 2463
rect 1860 2457 1916 2463
rect 1972 2457 1980 2463
rect 2900 2457 2908 2463
rect 2996 2457 3004 2463
rect 3076 2457 3244 2463
rect 3316 2457 3324 2463
rect 3348 2457 3356 2463
rect 1613 2444 1619 2456
rect 2717 2444 2723 2456
rect 1540 2437 1580 2443
rect 3188 2437 3196 2443
rect 948 2417 956 2423
rect 980 2417 1036 2423
rect 1572 2417 1580 2423
rect 2612 2417 2908 2423
rect 4052 2417 4124 2423
rect 644 2397 652 2403
rect 948 2397 1020 2403
rect 1732 2397 1852 2403
rect 2148 2397 2204 2403
rect 2212 2397 2236 2403
rect 2340 2397 3228 2403
rect 3236 2397 3484 2403
rect 3492 2397 3500 2403
rect 3508 2397 3644 2403
rect 1156 2377 1180 2383
rect 1716 2377 2012 2383
rect 2068 2377 2076 2383
rect 2452 2377 2460 2383
rect 2500 2377 2604 2383
rect 2628 2377 2828 2383
rect 2836 2377 2876 2383
rect 2884 2377 3436 2383
rect 3444 2377 3612 2383
rect 3620 2377 3724 2383
rect 3940 2377 3996 2383
rect 164 2357 188 2363
rect 388 2357 476 2363
rect 660 2357 668 2363
rect 996 2357 1020 2363
rect 1060 2357 1116 2363
rect 1380 2357 1436 2363
rect 1540 2357 1564 2363
rect 1620 2357 1628 2363
rect 1844 2357 1884 2363
rect 2340 2357 2892 2363
rect 2900 2357 2908 2363
rect 3092 2357 3100 2363
rect 3268 2357 3644 2363
rect 3940 2357 3948 2363
rect 276 2337 492 2343
rect 628 2337 636 2343
rect 644 2337 972 2343
rect 980 2337 1132 2343
rect 1140 2337 1164 2343
rect 1172 2337 1308 2343
rect 1332 2337 1404 2343
rect 1501 2343 1507 2356
rect 1428 2337 1692 2343
rect 1700 2337 2044 2343
rect 2052 2337 2060 2343
rect 2100 2337 2140 2343
rect 2228 2337 2460 2343
rect 2477 2337 2780 2343
rect 84 2317 156 2323
rect 164 2317 316 2323
rect 340 2317 348 2323
rect 372 2317 428 2323
rect 468 2317 476 2323
rect 596 2317 1004 2323
rect 1028 2317 1036 2323
rect 1188 2317 1196 2323
rect 1204 2317 1548 2323
rect 2477 2323 2483 2337
rect 2964 2337 2972 2343
rect 2996 2337 3900 2343
rect 3908 2337 4060 2343
rect 2781 2324 2787 2336
rect 1556 2317 2483 2323
rect 2548 2317 2556 2323
rect 2580 2317 2588 2323
rect 2788 2317 2988 2323
rect 3028 2317 3692 2323
rect 3700 2317 3868 2323
rect 3876 2317 3884 2323
rect 3908 2317 3948 2323
rect 4020 2317 4108 2323
rect 4116 2317 4156 2323
rect 228 2297 355 2303
rect 196 2277 332 2283
rect 349 2283 355 2297
rect 388 2297 412 2303
rect 436 2297 780 2303
rect 788 2297 1324 2303
rect 1332 2297 1436 2303
rect 1444 2297 1980 2303
rect 1988 2297 3212 2303
rect 3220 2297 3308 2303
rect 3316 2297 3708 2303
rect 3716 2297 3804 2303
rect 3812 2297 4092 2303
rect 4100 2297 4140 2303
rect 349 2277 460 2283
rect 532 2277 556 2283
rect 596 2277 604 2283
rect 724 2277 732 2283
rect 740 2277 828 2283
rect 836 2277 1196 2283
rect 1204 2277 2028 2283
rect 2052 2277 2092 2283
rect 2196 2277 2204 2283
rect 2260 2277 2316 2283
rect 2372 2277 2412 2283
rect 2436 2277 2444 2283
rect 2516 2277 2876 2283
rect 2884 2277 3196 2283
rect 3204 2277 3660 2283
rect 3668 2277 4124 2283
rect 4132 2277 4156 2283
rect -51 2257 12 2263
rect 100 2257 188 2263
rect 196 2257 284 2263
rect 356 2257 428 2263
rect 500 2257 556 2263
rect 820 2257 828 2263
rect 836 2257 1020 2263
rect 1060 2257 1388 2263
rect 1396 2257 1404 2263
rect 1460 2257 1468 2263
rect 1492 2257 1532 2263
rect 1556 2257 1628 2263
rect 1780 2257 1804 2263
rect 1844 2257 1884 2263
rect 1908 2257 1996 2263
rect 2036 2257 2492 2263
rect 2500 2257 2508 2263
rect 2532 2257 2812 2263
rect 2916 2257 3020 2263
rect 3188 2257 3564 2263
rect 3620 2257 3772 2263
rect 3780 2257 3932 2263
rect 3956 2257 4028 2263
rect 4084 2257 4140 2263
rect 4148 2257 4188 2263
rect 1725 2244 1731 2256
rect 20 2237 204 2243
rect 221 2237 387 2243
rect 221 2223 227 2237
rect 212 2217 227 2223
rect 381 2223 387 2237
rect 596 2237 668 2243
rect 836 2237 844 2243
rect 900 2237 972 2243
rect 1044 2237 1100 2243
rect 1124 2237 1132 2243
rect 1252 2237 1283 2243
rect 381 2217 1052 2223
rect 1277 2223 1283 2237
rect 1364 2237 1468 2243
rect 1524 2237 1596 2243
rect 1748 2237 1756 2243
rect 1796 2237 1820 2243
rect 1876 2237 2076 2243
rect 2084 2237 2540 2243
rect 2596 2237 2652 2243
rect 2660 2237 2668 2243
rect 2692 2237 2748 2243
rect 2804 2237 3100 2243
rect 3293 2237 3308 2243
rect 3444 2237 3468 2243
rect 3556 2237 3564 2243
rect 3588 2237 3603 2243
rect 3517 2224 3523 2236
rect 1277 2217 1308 2223
rect 1348 2217 1356 2223
rect 2468 2217 2492 2223
rect 2612 2217 2700 2223
rect 2852 2217 3276 2223
rect 3316 2217 3372 2223
rect 3597 2223 3603 2237
rect 3620 2237 3980 2243
rect 3988 2237 4188 2243
rect 4196 2237 4252 2243
rect 3597 2217 3724 2223
rect 3844 2217 3852 2223
rect 3908 2217 3916 2223
rect 3940 2217 3964 2223
rect 20 2197 156 2203
rect 500 2197 508 2203
rect 532 2197 956 2203
rect 964 2197 1116 2203
rect 1172 2197 1324 2203
rect 1348 2197 2236 2203
rect 2452 2197 2540 2203
rect 2852 2197 2908 2203
rect 68 2177 124 2183
rect 148 2177 748 2183
rect 804 2177 844 2183
rect 948 2177 988 2183
rect 1028 2177 1084 2183
rect 1236 2177 1244 2183
rect 1268 2177 1308 2183
rect 1332 2177 1436 2183
rect 1620 2177 1756 2183
rect 1780 2177 1852 2183
rect 1924 2177 1932 2183
rect 2004 2177 2012 2183
rect 2020 2177 3020 2183
rect 3028 2177 3036 2183
rect 3060 2177 3084 2183
rect 3156 2177 3436 2183
rect 3716 2177 3948 2183
rect 3956 2177 4028 2183
rect 4132 2177 4140 2183
rect 36 2157 60 2163
rect 260 2157 284 2163
rect 324 2157 540 2163
rect 596 2157 604 2163
rect 628 2157 828 2163
rect 836 2157 1356 2163
rect 1428 2157 1468 2163
rect 1588 2157 1660 2163
rect 1684 2157 1708 2163
rect 1844 2157 1884 2163
rect 1901 2157 1907 2176
rect 1924 2157 2028 2163
rect 2068 2157 2492 2163
rect 2509 2157 2524 2163
rect 2564 2157 2620 2163
rect 2772 2157 3084 2163
rect 3092 2157 3612 2163
rect 3636 2157 3692 2163
rect 3924 2157 4172 2163
rect 109 2144 115 2156
rect 221 2144 227 2156
rect 3709 2144 3715 2156
rect 3885 2144 3891 2156
rect 68 2137 92 2143
rect 276 2137 428 2143
rect 436 2137 844 2143
rect 852 2137 1068 2143
rect 1124 2137 1164 2143
rect 1188 2137 1292 2143
rect 1332 2137 1388 2143
rect 1588 2137 1596 2143
rect 1668 2137 1964 2143
rect 1972 2137 2572 2143
rect 2676 2137 2684 2143
rect 2772 2137 3548 2143
rect 3556 2137 3564 2143
rect 3572 2137 3580 2143
rect 3604 2137 3660 2143
rect 3764 2137 3804 2143
rect 3844 2137 3884 2143
rect 3924 2137 3964 2143
rect 4068 2137 4140 2143
rect 180 2117 284 2123
rect 324 2117 348 2123
rect 532 2117 540 2123
rect 596 2117 636 2123
rect 660 2117 700 2123
rect 740 2117 748 2123
rect 836 2117 876 2123
rect 900 2117 1036 2123
rect 1204 2117 1212 2123
rect 1348 2117 1580 2123
rect 1716 2117 2028 2123
rect 2036 2117 2092 2123
rect 2132 2117 2156 2123
rect 2196 2117 2268 2123
rect 2324 2117 2332 2123
rect 2484 2117 2892 2123
rect 2900 2117 2988 2123
rect 3012 2117 3132 2123
rect 3140 2117 3388 2123
rect 3572 2117 3580 2123
rect 3604 2117 3724 2123
rect 3812 2117 3836 2123
rect 4125 2104 4131 2116
rect 292 2097 316 2103
rect 564 2097 812 2103
rect 868 2097 1340 2103
rect 1380 2097 1564 2103
rect 1572 2097 1836 2103
rect 1844 2097 2236 2103
rect 2804 2097 2892 2103
rect 2916 2097 2956 2103
rect 2980 2097 2988 2103
rect 3108 2097 3164 2103
rect 3364 2097 3500 2103
rect 3508 2097 3932 2103
rect 3972 2097 3996 2103
rect 4052 2097 4076 2103
rect 4180 2097 4204 2103
rect 1837 2084 1843 2096
rect 2605 2084 2611 2096
rect 404 2077 684 2083
rect 788 2077 908 2083
rect 1252 2077 1260 2083
rect 1412 2077 1548 2083
rect 1556 2077 1692 2083
rect 1700 2077 1724 2083
rect 1812 2077 1820 2083
rect 2100 2077 2236 2083
rect 2244 2077 2588 2083
rect 2660 2077 2860 2083
rect 3588 2077 3788 2083
rect 388 2057 563 2063
rect 557 2043 563 2057
rect 596 2057 604 2063
rect 772 2057 1699 2063
rect 557 2037 876 2043
rect 1092 2037 1100 2043
rect 1108 2037 1164 2043
rect 1172 2037 1484 2043
rect 1604 2037 1628 2043
rect 1693 2043 1699 2057
rect 1940 2057 1980 2063
rect 1997 2057 2003 2076
rect 2020 2057 2028 2063
rect 2084 2057 2124 2063
rect 2285 2057 2572 2063
rect 1693 2037 2172 2043
rect 2285 2043 2291 2057
rect 3828 2057 3836 2063
rect 2180 2037 2291 2043
rect 2308 2037 2444 2043
rect 2452 2037 3004 2043
rect 3028 2037 3420 2043
rect 3428 2037 3756 2043
rect 1364 2017 1420 2023
rect 1732 2017 2028 2023
rect 2036 2017 2060 2023
rect 2100 2017 2108 2023
rect 2132 2017 2652 2023
rect 3108 2017 3196 2023
rect 3348 2017 3788 2023
rect 3796 2017 3916 2023
rect 1220 1997 1532 2003
rect 1620 1997 2012 2003
rect 2116 1997 2156 2003
rect 2452 1997 2460 2003
rect 2564 1997 2668 2003
rect 2740 1997 2748 2003
rect 3028 1997 3356 2003
rect 180 1977 348 1983
rect 644 1977 732 1983
rect 756 1977 4012 1983
rect 52 1957 316 1963
rect 628 1957 636 1963
rect 1652 1957 1740 1963
rect 1796 1957 1868 1963
rect 2084 1957 2124 1963
rect 2148 1957 2156 1963
rect 2244 1957 2252 1963
rect 2260 1957 2268 1963
rect 2308 1957 2316 1963
rect 2356 1957 2364 1963
rect 2404 1957 2460 1963
rect 2516 1957 2524 1963
rect 2564 1957 2844 1963
rect 2916 1957 3116 1963
rect 3124 1957 3404 1963
rect 3476 1957 3596 1963
rect 100 1937 188 1943
rect 244 1937 268 1943
rect 676 1937 716 1943
rect 804 1937 908 1943
rect 964 1937 1484 1943
rect 1540 1937 1564 1943
rect 1732 1937 1804 1943
rect 1812 1937 2508 1943
rect 2644 1937 2668 1943
rect 2836 1937 2844 1943
rect 2868 1937 2908 1943
rect 2948 1937 3052 1943
rect 3236 1937 3532 1943
rect 3732 1937 3820 1943
rect 3876 1937 3948 1943
rect 4036 1937 4076 1943
rect 4084 1937 4092 1943
rect -51 1863 -45 1923
rect 532 1917 540 1923
rect 724 1917 748 1923
rect 884 1917 1244 1923
rect 1252 1917 1788 1923
rect 1796 1917 1884 1923
rect 2116 1917 2412 1923
rect 2468 1917 2476 1923
rect 2532 1917 2540 1923
rect 2548 1917 2780 1923
rect 2820 1917 2972 1923
rect 2980 1917 3308 1923
rect 3428 1917 3548 1923
rect 3876 1917 3884 1923
rect 3892 1917 4108 1923
rect 1981 1904 1987 1916
rect 84 1897 124 1903
rect 308 1897 812 1903
rect 836 1897 844 1903
rect 852 1897 1692 1903
rect 1860 1897 1964 1903
rect 2004 1897 2092 1903
rect 2116 1897 2892 1903
rect 2900 1897 2908 1903
rect 3268 1897 3292 1903
rect 3348 1897 4108 1903
rect 20 1877 44 1883
rect 516 1877 732 1883
rect 948 1877 1020 1883
rect 1044 1877 1132 1883
rect 1188 1877 1196 1883
rect 1236 1877 1244 1883
rect 1252 1877 1260 1883
rect 1364 1877 1388 1883
rect 1396 1877 1660 1883
rect 1732 1877 1820 1883
rect 1844 1877 1852 1883
rect 1876 1877 1884 1883
rect 1924 1877 1932 1883
rect 1956 1877 1980 1883
rect 2004 1877 2012 1883
rect 2052 1877 2492 1883
rect 2516 1877 2620 1883
rect 2644 1877 3004 1883
rect 3060 1877 3180 1883
rect 3380 1877 3516 1883
rect 3588 1877 3708 1883
rect 4004 1877 4076 1883
rect 4164 1877 4220 1883
rect 125 1864 131 1876
rect -51 1857 28 1863
rect 212 1857 252 1863
rect 333 1863 339 1876
rect 1341 1864 1347 1876
rect 333 1857 348 1863
rect 644 1857 716 1863
rect 724 1857 988 1863
rect 1124 1857 1292 1863
rect 1412 1857 2300 1863
rect 2308 1857 2812 1863
rect 2932 1857 2956 1863
rect 3300 1857 3308 1863
rect 3380 1857 3740 1863
rect 3748 1857 3852 1863
rect 3988 1857 4012 1863
rect 4020 1857 4044 1863
rect 4116 1857 4131 1863
rect 445 1844 451 1856
rect 1293 1844 1299 1856
rect 372 1837 380 1843
rect 724 1837 764 1843
rect 797 1837 812 1843
rect 1236 1837 1244 1843
rect 1380 1837 1404 1843
rect 1492 1837 1500 1843
rect 1572 1837 1596 1843
rect 1620 1837 1628 1843
rect 1764 1837 1772 1843
rect 1796 1837 2124 1843
rect 2276 1837 2284 1843
rect 2308 1837 2540 1843
rect 2548 1837 2556 1843
rect 2580 1837 2636 1843
rect 2740 1837 3036 1843
rect 3620 1837 3660 1843
rect 3940 1837 4156 1843
rect 1012 1817 1692 1823
rect 1860 1817 1948 1823
rect 2004 1817 2124 1823
rect 2276 1817 2396 1823
rect 2468 1817 3260 1823
rect 3460 1817 3580 1823
rect 692 1797 940 1803
rect 1172 1797 1180 1803
rect 1332 1797 1420 1803
rect 1876 1797 1900 1803
rect 2084 1797 2316 1803
rect 2452 1797 2508 1803
rect 2964 1797 3052 1803
rect 3092 1797 3308 1803
rect 3476 1797 3612 1803
rect -51 1777 12 1783
rect 308 1777 364 1783
rect 692 1777 700 1783
rect 708 1777 796 1783
rect 804 1777 1180 1783
rect 1284 1777 1340 1783
rect 1364 1777 1507 1783
rect 132 1757 204 1763
rect 260 1757 316 1763
rect 340 1757 460 1763
rect 484 1757 508 1763
rect 660 1757 684 1763
rect 756 1757 780 1763
rect 836 1757 860 1763
rect 1076 1757 1100 1763
rect 1156 1757 1180 1763
rect 1204 1757 1292 1763
rect 1332 1757 1340 1763
rect 1501 1763 1507 1777
rect 1604 1777 1740 1783
rect 1828 1777 1916 1783
rect 2020 1777 2204 1783
rect 2212 1777 2220 1783
rect 2260 1777 2428 1783
rect 2772 1777 2844 1783
rect 2884 1777 2972 1783
rect 3012 1777 3020 1783
rect 3076 1777 3100 1783
rect 3124 1777 3196 1783
rect 3220 1777 3484 1783
rect 3652 1777 3660 1783
rect 3828 1777 3980 1783
rect 4020 1777 4028 1783
rect 4180 1777 4204 1783
rect 1501 1757 1532 1763
rect 1540 1757 1580 1763
rect 1620 1757 1628 1763
rect 1684 1757 1948 1763
rect 2052 1757 2156 1763
rect 2212 1757 2220 1763
rect 2324 1757 2380 1763
rect 2420 1757 2460 1763
rect 2532 1757 2556 1763
rect 2596 1757 2716 1763
rect 2756 1757 2796 1763
rect 2868 1757 2876 1763
rect 2900 1757 3340 1763
rect 3508 1757 3516 1763
rect 3540 1757 3564 1763
rect 3636 1757 3683 1763
rect 1485 1744 1491 1756
rect 2493 1744 2499 1756
rect 20 1737 236 1743
rect 276 1737 348 1743
rect 500 1737 652 1743
rect 660 1737 1212 1743
rect 1348 1737 1372 1743
rect 1508 1737 1596 1743
rect 1620 1737 1852 1743
rect 1892 1737 1900 1743
rect 2212 1737 2444 1743
rect 2452 1737 2492 1743
rect 2580 1737 2588 1743
rect 2756 1737 2796 1743
rect 2916 1737 3164 1743
rect 3204 1737 3228 1743
rect 3236 1737 3404 1743
rect 3412 1737 3644 1743
rect 3677 1743 3683 1757
rect 3780 1757 3836 1763
rect 3844 1757 3852 1763
rect 3876 1757 3884 1763
rect 4020 1757 4044 1763
rect 4116 1757 4124 1763
rect 3677 1737 3859 1743
rect 1325 1724 1331 1736
rect 3853 1724 3859 1737
rect 3876 1737 3980 1743
rect 4036 1737 4044 1743
rect 4068 1737 4140 1743
rect 1284 1717 1292 1723
rect 1412 1717 1452 1723
rect 1460 1717 1660 1723
rect 2068 1717 2108 1723
rect 2116 1717 2156 1723
rect 2260 1717 2300 1723
rect 2356 1717 2604 1723
rect 2612 1717 3196 1723
rect 3252 1717 3260 1723
rect 3284 1717 3292 1723
rect 3316 1717 3340 1723
rect 3396 1717 3676 1723
rect 1789 1704 1795 1716
rect 1220 1697 1292 1703
rect 1300 1697 1772 1703
rect 1796 1697 2108 1703
rect 2116 1697 2124 1703
rect 2164 1697 2172 1703
rect 2212 1697 2252 1703
rect 2628 1697 3020 1703
rect 3044 1697 3068 1703
rect 3076 1697 3100 1703
rect 3124 1697 3292 1703
rect 3684 1697 3708 1703
rect 4036 1697 4076 1703
rect 3293 1684 3299 1696
rect 3373 1684 3379 1696
rect 1140 1677 1356 1683
rect 1412 1677 1484 1683
rect 1620 1677 1916 1683
rect 2004 1677 2476 1683
rect 2653 1677 2924 1683
rect 916 1657 1036 1663
rect 1044 1657 1084 1663
rect 1092 1657 1660 1663
rect 2148 1657 2156 1663
rect 2212 1657 2236 1663
rect 2292 1657 2300 1663
rect 2653 1663 2659 1677
rect 3012 1677 3084 1683
rect 3204 1677 3212 1683
rect 3252 1677 3283 1683
rect 2596 1657 2659 1663
rect 2676 1657 3260 1663
rect 3277 1663 3283 1677
rect 3348 1677 3356 1683
rect 3684 1677 3788 1683
rect 3277 1657 3356 1663
rect 3524 1657 3532 1663
rect 516 1637 796 1643
rect 1828 1637 1964 1643
rect 1972 1637 3580 1643
rect 3700 1637 3708 1643
rect 3828 1637 3980 1643
rect 3988 1637 4092 1643
rect 1748 1617 1884 1623
rect 1892 1617 2076 1623
rect 2084 1617 2348 1623
rect 2388 1617 2812 1623
rect 2836 1617 2924 1623
rect 2932 1617 3212 1623
rect 3588 1617 3596 1623
rect 3636 1617 3660 1623
rect 3796 1617 3804 1623
rect 4180 1617 4188 1623
rect 132 1597 140 1603
rect 228 1597 236 1603
rect 356 1597 396 1603
rect 436 1597 492 1603
rect 596 1597 780 1603
rect 980 1597 1388 1603
rect 1860 1597 1868 1603
rect 2084 1597 2172 1603
rect 2180 1597 2396 1603
rect 2468 1597 2524 1603
rect 2564 1597 2668 1603
rect 2692 1597 3324 1603
rect 3348 1597 3436 1603
rect 3444 1597 3612 1603
rect 3700 1597 4108 1603
rect 4164 1597 4172 1603
rect 132 1577 172 1583
rect 228 1577 1020 1583
rect 1028 1577 1164 1583
rect 1332 1577 1372 1583
rect 1492 1577 1516 1583
rect 1620 1577 1724 1583
rect 1732 1577 1868 1583
rect 1876 1577 2428 1583
rect 2436 1577 2700 1583
rect 2708 1577 3628 1583
rect 3636 1577 3740 1583
rect 4132 1577 4220 1583
rect 84 1557 236 1563
rect 468 1557 508 1563
rect 724 1557 860 1563
rect 1140 1557 1340 1563
rect 1572 1557 1580 1563
rect 1892 1557 2028 1563
rect 2084 1557 2092 1563
rect 2196 1557 2204 1563
rect 2244 1557 2252 1563
rect 2260 1557 2860 1563
rect 2916 1557 2988 1563
rect 3076 1557 3116 1563
rect 3316 1557 3388 1563
rect 3604 1557 3628 1563
rect 3700 1557 3836 1563
rect 420 1537 1004 1543
rect 1428 1537 2348 1543
rect 2420 1537 2476 1543
rect 2580 1537 2796 1543
rect 3076 1537 3420 1543
rect 3428 1537 3692 1543
rect 3732 1537 3964 1543
rect -51 1517 -29 1523
rect -35 1483 -29 1517
rect 500 1517 524 1523
rect 596 1517 620 1523
rect 740 1517 748 1523
rect 900 1517 924 1523
rect 1204 1517 1244 1523
rect 1364 1517 1372 1523
rect 1460 1517 1708 1523
rect 1716 1517 2268 1523
rect 2324 1517 2332 1523
rect 2404 1517 2428 1523
rect 2564 1517 2636 1523
rect 2660 1517 2764 1523
rect 2868 1517 2892 1523
rect 2916 1517 2940 1523
rect 3156 1517 3164 1523
rect 3444 1517 3484 1523
rect 4068 1517 4092 1523
rect 4164 1517 4172 1523
rect 4228 1517 4252 1523
rect 1421 1504 1427 1516
rect 2957 1504 2963 1516
rect 3341 1504 3347 1516
rect 132 1497 412 1503
rect 436 1497 492 1503
rect 756 1497 812 1503
rect 1044 1497 1084 1503
rect 1092 1497 1404 1503
rect 1476 1497 1900 1503
rect 1908 1497 2252 1503
rect 2260 1497 2428 1503
rect 2452 1497 2604 1503
rect 2660 1497 2908 1503
rect 3156 1497 3244 1503
rect 3444 1497 3452 1503
rect 3572 1497 3587 1503
rect 845 1484 851 1496
rect 3133 1484 3139 1496
rect 3581 1484 3587 1497
rect 3652 1497 3724 1503
rect 3732 1497 3884 1503
rect 4132 1497 4140 1503
rect 3613 1484 3619 1496
rect -35 1477 12 1483
rect 164 1477 188 1483
rect 244 1477 291 1483
rect 84 1457 108 1463
rect 260 1457 268 1463
rect 285 1463 291 1477
rect 308 1477 332 1483
rect 596 1477 620 1483
rect 692 1477 732 1483
rect 884 1477 892 1483
rect 932 1477 956 1483
rect 1108 1477 1132 1483
rect 1220 1477 1260 1483
rect 1300 1477 1308 1483
rect 1316 1477 1564 1483
rect 1572 1477 1580 1483
rect 1700 1477 1708 1483
rect 1828 1477 1836 1483
rect 1956 1477 2012 1483
rect 2052 1477 2060 1483
rect 2084 1477 2172 1483
rect 2180 1477 2268 1483
rect 2324 1477 2460 1483
rect 2516 1477 2588 1483
rect 2612 1477 2620 1483
rect 2724 1477 2732 1483
rect 2772 1477 3132 1483
rect 3252 1477 3260 1483
rect 3364 1477 3484 1483
rect 3524 1477 3532 1483
rect 3732 1477 3756 1483
rect 3917 1483 3923 1496
rect 3917 1477 3932 1483
rect 3956 1477 3996 1483
rect 4221 1464 4227 1476
rect 285 1457 316 1463
rect 404 1457 412 1463
rect 628 1457 1500 1463
rect 1540 1457 1628 1463
rect 1684 1457 1708 1463
rect 1796 1457 1948 1463
rect 1956 1457 2492 1463
rect 2500 1457 2508 1463
rect 2548 1457 2579 1463
rect 381 1444 387 1456
rect 20 1437 332 1443
rect 532 1437 652 1443
rect 836 1437 876 1443
rect 900 1437 1116 1443
rect 1172 1437 1212 1443
rect 1316 1437 1372 1443
rect 1412 1437 1468 1443
rect 2036 1437 2092 1443
rect 2132 1437 2188 1443
rect 2228 1437 2396 1443
rect 2420 1437 2476 1443
rect 2500 1437 2556 1443
rect 2573 1443 2579 1457
rect 2612 1457 2684 1463
rect 2724 1457 2844 1463
rect 2900 1457 3020 1463
rect 3284 1457 3660 1463
rect 3716 1457 3756 1463
rect 3796 1457 3932 1463
rect 3972 1457 4060 1463
rect 4100 1457 4188 1463
rect 3101 1444 3107 1456
rect 2573 1437 2780 1443
rect 2836 1437 2988 1443
rect 3204 1437 3628 1443
rect 3716 1437 4028 1443
rect 4084 1437 4156 1443
rect 212 1417 300 1423
rect 436 1417 444 1423
rect 1364 1417 1372 1423
rect 1444 1417 1548 1423
rect 1604 1417 1660 1423
rect 2308 1417 2387 1423
rect 893 1404 899 1416
rect 212 1397 444 1403
rect 1236 1397 1244 1403
rect 1252 1397 1548 1403
rect 1652 1397 2028 1403
rect 2093 1397 2332 1403
rect 84 1377 220 1383
rect 420 1377 428 1383
rect 804 1377 844 1383
rect 932 1377 1068 1383
rect 1092 1377 1308 1383
rect 1332 1377 1420 1383
rect 1469 1377 1772 1383
rect 116 1357 140 1363
rect 260 1357 380 1363
rect 404 1357 444 1363
rect 468 1357 492 1363
rect 740 1357 764 1363
rect 964 1357 1020 1363
rect 1469 1363 1475 1377
rect 2093 1383 2099 1397
rect 2381 1403 2387 1417
rect 2404 1417 2428 1423
rect 2468 1417 2540 1423
rect 2660 1417 2876 1423
rect 2900 1417 2940 1423
rect 3092 1417 3100 1423
rect 3444 1417 3468 1423
rect 3588 1417 3596 1423
rect 3668 1417 3692 1423
rect 3956 1417 4108 1423
rect 3341 1404 3347 1416
rect 2381 1397 2412 1403
rect 2452 1397 2460 1403
rect 2484 1397 2668 1403
rect 2692 1397 2812 1403
rect 2836 1397 2844 1403
rect 2852 1397 3308 1403
rect 1780 1377 2099 1383
rect 2276 1377 2316 1383
rect 2420 1377 2476 1383
rect 2516 1377 2572 1383
rect 2580 1377 2620 1383
rect 2740 1377 2748 1383
rect 2772 1377 2812 1383
rect 2964 1377 2972 1383
rect 2996 1377 3004 1383
rect 3044 1377 3052 1383
rect 3076 1377 3100 1383
rect 3124 1377 3212 1383
rect 3236 1377 3244 1383
rect 3348 1377 3372 1383
rect 3476 1377 3612 1383
rect 3620 1377 3676 1383
rect 3700 1377 3852 1383
rect 3876 1377 3980 1383
rect 4052 1377 4092 1383
rect 1060 1357 1475 1363
rect 1508 1357 1516 1363
rect 1572 1357 1580 1363
rect 1668 1357 1820 1363
rect 1892 1357 1996 1363
rect 2013 1357 2028 1363
rect 2132 1357 2204 1363
rect 2292 1357 2316 1363
rect 2324 1357 2396 1363
rect 2436 1357 2444 1363
rect 2484 1357 2508 1363
rect 2532 1357 2540 1363
rect 2580 1357 2588 1363
rect 2708 1357 2716 1363
rect 2756 1357 2764 1363
rect 2788 1357 2796 1363
rect 2909 1363 2915 1376
rect 2909 1357 2924 1363
rect 2964 1357 3068 1363
rect 3092 1357 3132 1363
rect 3316 1357 3452 1363
rect 3460 1357 3756 1363
rect 3780 1357 3884 1363
rect 4100 1357 4124 1363
rect 4164 1357 4204 1363
rect 1885 1344 1891 1356
rect 3965 1344 3971 1356
rect 52 1337 220 1343
rect 484 1337 508 1343
rect 548 1337 588 1343
rect 756 1337 796 1343
rect 804 1337 812 1343
rect 1028 1337 1340 1343
rect 1364 1337 1404 1343
rect 1492 1337 1500 1343
rect 1508 1337 1692 1343
rect 1764 1337 1804 1343
rect 1908 1337 1916 1343
rect 2132 1337 2188 1343
rect 2276 1337 2284 1343
rect 2292 1337 2556 1343
rect 2564 1337 2876 1343
rect 2900 1337 2924 1343
rect 2932 1337 3372 1343
rect 3444 1337 3820 1343
rect 3828 1337 3836 1343
rect 4100 1337 4236 1343
rect 436 1317 476 1323
rect 484 1317 652 1323
rect 660 1317 700 1323
rect 708 1317 828 1323
rect 836 1317 1100 1323
rect 1108 1317 1212 1323
rect 1220 1317 1292 1323
rect 1844 1317 2012 1323
rect 2020 1317 2316 1323
rect 2324 1317 2396 1323
rect 2436 1317 3612 1323
rect 3620 1317 3724 1323
rect 4148 1317 4156 1323
rect 660 1297 668 1303
rect 932 1297 940 1303
rect 964 1297 1004 1303
rect 1076 1297 1084 1303
rect 1316 1297 1356 1303
rect 1373 1297 1379 1316
rect 1396 1297 1756 1303
rect 1828 1297 1932 1303
rect 2020 1297 2028 1303
rect 2068 1297 2140 1303
rect 2164 1297 2179 1303
rect 93 1284 99 1296
rect 797 1284 803 1296
rect 1293 1284 1299 1296
rect 2141 1284 2147 1296
rect 2173 1284 2179 1297
rect 2404 1297 2524 1303
rect 2580 1297 2588 1303
rect 2612 1297 2620 1303
rect 2676 1297 2780 1303
rect 2804 1297 2892 1303
rect 2916 1297 3260 1303
rect 3268 1297 3340 1303
rect 3380 1297 3452 1303
rect 3476 1297 3484 1303
rect 3780 1297 3788 1303
rect 3908 1297 3948 1303
rect 4004 1297 4204 1303
rect 804 1277 972 1283
rect 1060 1277 1228 1283
rect 1348 1277 1436 1283
rect 1460 1277 1468 1283
rect 1492 1277 1516 1283
rect 1588 1277 1596 1283
rect 1732 1277 2076 1283
rect 2180 1277 2387 1283
rect 548 1257 604 1263
rect 612 1257 668 1263
rect 676 1257 1484 1263
rect 1492 1257 2188 1263
rect 2228 1257 2252 1263
rect 2381 1263 2387 1277
rect 2404 1277 2892 1283
rect 2900 1277 3388 1283
rect 3460 1277 3580 1283
rect 2381 1257 2444 1263
rect 2516 1257 2652 1263
rect 2916 1257 2940 1263
rect 3220 1257 3484 1263
rect 3764 1257 3916 1263
rect 2989 1244 2995 1256
rect 932 1237 972 1243
rect 1348 1237 1740 1243
rect 2708 1237 2716 1243
rect 3396 1237 3436 1243
rect 3716 1237 3788 1243
rect 3796 1237 4220 1243
rect 852 1217 1564 1223
rect 1572 1217 1612 1223
rect 2372 1217 2412 1223
rect 2852 1217 3404 1223
rect 3508 1217 3516 1223
rect 500 1197 556 1203
rect 564 1197 1100 1203
rect 1108 1197 1532 1203
rect 1540 1197 1612 1203
rect 1620 1197 1852 1203
rect 1972 1197 2156 1203
rect 2212 1197 2220 1203
rect 2484 1197 2716 1203
rect 2740 1197 2860 1203
rect 3012 1197 3532 1203
rect 4068 1197 4252 1203
rect 772 1177 780 1183
rect 852 1177 1180 1183
rect 1540 1177 2076 1183
rect 2084 1177 2316 1183
rect 2612 1177 2812 1183
rect 2852 1177 2892 1183
rect 3172 1177 3356 1183
rect 3668 1177 3724 1183
rect 228 1157 252 1163
rect 628 1157 1020 1163
rect 1604 1157 1692 1163
rect 1716 1157 1900 1163
rect 1924 1157 2028 1163
rect 2036 1157 2092 1163
rect 2228 1157 2268 1163
rect 2308 1157 2380 1163
rect 2516 1157 2908 1163
rect 2916 1157 3292 1163
rect 3300 1157 3356 1163
rect 3380 1157 3452 1163
rect 3620 1157 3628 1163
rect 2285 1144 2291 1156
rect 388 1137 412 1143
rect 468 1137 588 1143
rect 660 1137 716 1143
rect 900 1137 972 1143
rect 980 1137 1004 1143
rect 1668 1137 1692 1143
rect 1700 1137 1708 1143
rect 1812 1137 1932 1143
rect 2004 1137 2012 1143
rect 2148 1137 2172 1143
rect 2244 1137 2252 1143
rect 2404 1137 2476 1143
rect 2548 1137 3372 1143
rect 3380 1137 3484 1143
rect 3492 1137 3580 1143
rect 3636 1137 3900 1143
rect 3956 1137 4044 1143
rect 765 1124 771 1136
rect 244 1117 284 1123
rect 340 1117 668 1123
rect 772 1117 988 1123
rect 1092 1117 1100 1123
rect 1284 1117 1292 1123
rect 1332 1117 1372 1123
rect 1652 1117 1804 1123
rect 1812 1117 1820 1123
rect 1828 1117 2460 1123
rect 2628 1117 2636 1123
rect 2644 1117 2684 1123
rect 2772 1117 2780 1123
rect 2804 1117 2876 1123
rect 2948 1117 2988 1123
rect 3092 1117 3132 1123
rect 3428 1117 3436 1123
rect 3444 1117 3756 1123
rect 3764 1117 3996 1123
rect 4212 1117 4220 1123
rect 3181 1104 3187 1116
rect 436 1097 508 1103
rect 548 1097 604 1103
rect 644 1097 652 1103
rect 868 1097 940 1103
rect 1140 1097 1244 1103
rect 1252 1097 2012 1103
rect 2164 1097 2284 1103
rect 2292 1097 2428 1103
rect 2436 1097 2444 1103
rect 2724 1097 2732 1103
rect 3316 1097 3324 1103
rect 3412 1097 3564 1103
rect 3652 1097 3868 1103
rect 3892 1097 3964 1103
rect 2557 1084 2563 1096
rect 84 1077 156 1083
rect 164 1077 268 1083
rect 292 1077 316 1083
rect 372 1077 396 1083
rect 404 1077 556 1083
rect 724 1077 732 1083
rect 740 1077 812 1083
rect 1124 1077 1132 1083
rect 1140 1077 1644 1083
rect 1668 1077 1676 1083
rect 1844 1077 1852 1083
rect 1860 1077 1900 1083
rect 1972 1077 2172 1083
rect 2212 1077 2412 1083
rect 2420 1077 2460 1083
rect 2612 1077 2620 1083
rect 2676 1077 2828 1083
rect 2868 1077 3084 1083
rect 3140 1077 3516 1083
rect 3556 1077 3676 1083
rect 3700 1077 3715 1083
rect 3796 1077 3820 1083
rect 3844 1077 3852 1083
rect 3860 1077 3916 1083
rect 4180 1077 4204 1083
rect 621 1064 627 1076
rect 100 1057 140 1063
rect 260 1057 380 1063
rect 532 1057 540 1063
rect 564 1057 572 1063
rect 628 1057 1036 1063
rect 1044 1057 1084 1063
rect 1252 1057 1340 1063
rect 1412 1057 1468 1063
rect 1492 1057 1507 1063
rect 1524 1057 1596 1063
rect 1620 1057 1660 1063
rect 1732 1057 1756 1063
rect 1780 1057 1868 1063
rect 1972 1057 2380 1063
rect 2404 1057 2476 1063
rect 2596 1057 2604 1063
rect 2692 1057 2732 1063
rect 2868 1057 2876 1063
rect 2932 1057 2972 1063
rect 3076 1057 3100 1063
rect 3213 1057 3228 1063
rect 189 1044 195 1056
rect 3213 1044 3219 1057
rect 3252 1057 3267 1063
rect 3261 1044 3267 1057
rect 3284 1057 3308 1063
rect 3380 1057 4188 1063
rect 356 1037 428 1043
rect 500 1037 675 1043
rect 148 1017 284 1023
rect 669 1023 675 1037
rect 724 1037 780 1043
rect 852 1037 908 1043
rect 980 1037 1788 1043
rect 1908 1037 2044 1043
rect 2084 1037 2124 1043
rect 2180 1037 2652 1043
rect 2724 1037 2828 1043
rect 2852 1037 2988 1043
rect 3012 1037 3148 1043
rect 3396 1037 3484 1043
rect 3588 1037 3692 1043
rect 3732 1037 3772 1043
rect 4004 1037 4076 1043
rect 4148 1037 4156 1043
rect 669 1017 860 1023
rect 980 1017 1228 1023
rect 1252 1017 1260 1023
rect 1428 1017 1500 1023
rect 1556 1017 1564 1023
rect 1764 1017 3740 1023
rect 4132 1017 4140 1023
rect 628 997 684 1003
rect 820 997 876 1003
rect 900 997 908 1003
rect 1012 997 1036 1003
rect 1396 997 2572 1003
rect 2612 997 2620 1003
rect 2724 997 2755 1003
rect 196 977 252 983
rect 260 977 444 983
rect 596 977 652 983
rect 660 977 748 983
rect 772 977 780 983
rect 916 977 924 983
rect 1204 977 1244 983
rect 1364 977 1404 983
rect 1684 977 2732 983
rect 2749 983 2755 997
rect 2788 997 2828 1003
rect 2868 997 2940 1003
rect 2980 997 3004 1003
rect 3156 997 3164 1003
rect 3444 997 3468 1003
rect 3540 997 3836 1003
rect 4196 997 4204 1003
rect 2957 984 2963 996
rect 2749 977 2908 983
rect 3092 977 3228 983
rect 3236 977 3292 983
rect 3316 977 3324 983
rect 3460 977 3644 983
rect 3956 977 3996 983
rect 4052 977 4156 983
rect 4212 977 4236 983
rect 509 964 515 976
rect 1485 964 1491 976
rect 2733 964 2739 976
rect 132 957 140 963
rect 164 957 172 963
rect 308 957 364 963
rect 468 957 492 963
rect 628 957 684 963
rect 692 957 1052 963
rect 1076 957 1132 963
rect 1140 957 1276 963
rect 1556 957 1612 963
rect 1620 957 2140 963
rect 2196 957 2348 963
rect 2372 957 2412 963
rect 2452 957 2492 963
rect 2509 957 2668 963
rect 1437 944 1443 956
rect 244 937 316 943
rect 324 937 1436 943
rect 1444 937 1740 943
rect 1764 937 1804 943
rect 1828 937 1948 943
rect 1956 937 1964 943
rect 1988 937 1996 943
rect 2036 937 2092 943
rect 2196 937 2220 943
rect 2228 937 2300 943
rect 2324 937 2364 943
rect 2509 943 2515 957
rect 2836 957 3196 963
rect 3236 957 3244 963
rect 3316 957 3356 963
rect 3460 957 3468 963
rect 3492 957 3516 963
rect 3524 957 3564 963
rect 3620 957 3628 963
rect 3652 957 3660 963
rect 3700 957 3868 963
rect 3924 957 3980 963
rect 2468 937 2515 943
rect 2548 937 2620 943
rect 2820 937 2844 943
rect 2884 937 3276 943
rect 3284 937 3772 943
rect 3780 937 3788 943
rect 3860 937 3884 943
rect 4036 937 4060 943
rect 4100 937 4124 943
rect 3917 924 3923 936
rect 756 917 764 923
rect 1188 917 1292 923
rect 1316 917 1372 923
rect 1396 917 1900 923
rect 1965 917 1980 923
rect 2004 917 2012 923
rect 2036 917 2044 923
rect 2084 917 2188 923
rect 2260 917 2268 923
rect 2292 917 2316 923
rect 2340 917 2348 923
rect 2452 917 2972 923
rect 2996 917 3356 923
rect 3380 917 3459 923
rect 861 904 867 916
rect 1021 904 1027 916
rect 1133 904 1139 916
rect 100 897 124 903
rect 340 897 348 903
rect 356 897 396 903
rect 404 897 572 903
rect 676 897 764 903
rect 1252 897 1260 903
rect 1284 897 1468 903
rect 1492 897 1612 903
rect 1661 897 1836 903
rect 708 877 716 883
rect 1661 883 1667 897
rect 1860 897 1980 903
rect 2036 897 2300 903
rect 2564 897 2572 903
rect 2644 897 2652 903
rect 2692 897 2940 903
rect 3028 897 3052 903
rect 3124 897 3196 903
rect 3428 897 3436 903
rect 3453 903 3459 917
rect 3476 917 3612 923
rect 3620 917 3788 923
rect 3828 917 3900 923
rect 4052 917 4060 923
rect 4068 917 4108 923
rect 3453 897 3516 903
rect 3604 897 3612 903
rect 3636 897 3644 903
rect 3668 897 3692 903
rect 3908 897 4028 903
rect 3533 884 3539 896
rect 3549 884 3555 896
rect 3741 884 3747 896
rect 724 877 1667 883
rect 1732 877 1868 883
rect 1876 877 2092 883
rect 2116 877 2172 883
rect 2180 877 2284 883
rect 2420 877 2556 883
rect 2692 877 2828 883
rect 3428 877 3436 883
rect 3460 877 3500 883
rect 1396 857 1404 863
rect 1540 857 1548 863
rect 1588 857 1644 863
rect 1892 857 1900 863
rect 3188 857 3267 863
rect 468 837 1164 843
rect 1268 837 1276 843
rect 1444 837 1580 843
rect 2356 837 2476 843
rect 2900 837 3244 843
rect 3261 843 3267 857
rect 3261 837 3660 843
rect 3668 837 4076 843
rect 148 817 284 823
rect 884 817 940 823
rect 1764 817 1772 823
rect 3316 817 3356 823
rect 3572 817 3676 823
rect 3924 817 3964 823
rect 804 797 828 803
rect 1428 797 1436 803
rect 1572 797 1580 803
rect 2356 797 2380 803
rect 2756 797 2844 803
rect 3028 797 3164 803
rect 3252 797 3404 803
rect 436 777 524 783
rect 804 777 892 783
rect 900 777 1052 783
rect 1060 777 1596 783
rect 1604 777 1628 783
rect 1652 777 1660 783
rect 1684 777 1756 783
rect 1764 777 2060 783
rect 2068 777 2156 783
rect 2164 777 3148 783
rect 4036 777 4108 783
rect 196 757 668 763
rect 1076 757 1084 763
rect 1236 757 1692 763
rect 1700 757 1708 763
rect 1924 757 1932 763
rect 2324 757 2572 763
rect 2644 757 2684 763
rect 2916 757 3228 763
rect 4116 757 4188 763
rect 3437 744 3443 756
rect 52 737 124 743
rect 372 737 652 743
rect 964 737 1292 743
rect 1476 737 1484 743
rect 1492 737 1724 743
rect 1860 737 1884 743
rect 2212 737 2236 743
rect 2308 737 2364 743
rect 2420 737 2428 743
rect 2484 737 2540 743
rect 2564 737 2572 743
rect 2612 737 2620 743
rect 2676 737 3196 743
rect 3268 737 3276 743
rect 1949 724 1955 736
rect 260 717 300 723
rect 516 717 764 723
rect 772 717 1068 723
rect 1092 717 1116 723
rect 1172 717 1180 723
rect 1572 717 1596 723
rect 1604 717 1692 723
rect 1700 717 1948 723
rect 2109 723 2115 736
rect 3453 724 3459 736
rect 2100 717 2115 723
rect 2132 717 2147 723
rect 2164 717 2268 723
rect 2276 717 2332 723
rect 2388 717 2396 723
rect 2420 717 2460 723
rect 2516 717 2764 723
rect 2772 717 2924 723
rect 2964 717 2988 723
rect 3028 717 3052 723
rect 3076 717 3452 723
rect 3460 717 3868 723
rect 3876 717 3884 723
rect 3956 717 3964 723
rect 4148 717 4188 723
rect 468 697 476 703
rect 692 697 700 703
rect 740 697 812 703
rect 836 697 844 703
rect 1060 697 1084 703
rect 1156 697 1212 703
rect 1236 697 1244 703
rect 1268 697 1324 703
rect 1380 697 1900 703
rect 1908 697 1980 703
rect 1988 697 2140 703
rect 2148 697 2764 703
rect 2884 697 2924 703
rect 3396 697 3628 703
rect 3684 697 3820 703
rect 397 684 403 696
rect 3149 684 3155 696
rect 116 677 156 683
rect 244 677 364 683
rect 404 677 604 683
rect 612 677 1452 683
rect 1460 677 1612 683
rect 1652 677 1836 683
rect 1892 677 1948 683
rect 1972 677 2028 683
rect 2116 677 2188 683
rect 2196 677 2204 683
rect 2212 677 2716 683
rect 2836 677 2908 683
rect 2948 677 3132 683
rect 3316 677 3468 683
rect 3636 677 3676 683
rect 3684 677 3740 683
rect 3828 677 3843 683
rect 4116 677 4156 683
rect 3581 664 3587 676
rect 116 657 220 663
rect 356 657 412 663
rect 660 657 860 663
rect 980 657 1980 663
rect 2020 657 2060 663
rect 2260 657 2284 663
rect 2324 657 2332 663
rect 2356 657 2556 663
rect 2564 657 3244 663
rect 3364 657 3516 663
rect 3540 657 3548 663
rect 3684 657 3740 663
rect 3780 657 3852 663
rect 4084 657 4108 663
rect 452 637 1372 643
rect 1540 637 1660 643
rect 1844 637 1916 643
rect 2276 637 2300 643
rect 2468 637 2572 643
rect 2612 637 2684 643
rect 2692 637 2700 643
rect 2740 637 2876 643
rect 3108 637 3116 643
rect 3348 637 3356 643
rect 3412 637 3884 643
rect 164 617 524 623
rect 580 617 620 623
rect 788 617 924 623
rect 1140 617 1164 623
rect 1316 617 1404 623
rect 2292 617 2300 623
rect 2436 617 2444 623
rect 2884 617 3020 623
rect 3092 617 3100 623
rect 3204 617 3372 623
rect 3380 617 3596 623
rect 3716 617 3724 623
rect 340 597 348 603
rect 676 597 828 603
rect 1012 597 1020 603
rect 1364 597 1372 603
rect 1412 597 1500 603
rect 1620 597 1644 603
rect 1748 597 1836 603
rect 1956 597 1964 603
rect 2388 597 2412 603
rect 2868 597 2892 603
rect 3332 597 3356 603
rect 3588 597 3948 603
rect 3309 584 3315 596
rect 212 577 284 583
rect 308 577 332 583
rect 612 577 860 583
rect 868 577 1420 583
rect 1428 577 2012 583
rect 2020 577 2140 583
rect 2228 577 2284 583
rect 2308 577 2844 583
rect 2964 577 3036 583
rect 3364 577 3372 583
rect 3476 577 3916 583
rect 3924 577 3964 583
rect 372 557 412 563
rect 564 557 604 563
rect 628 557 716 563
rect 820 557 1004 563
rect 1028 557 1068 563
rect 1364 557 1388 563
rect 1428 557 1484 563
rect 1508 557 1548 563
rect 1636 557 1644 563
rect 1892 557 1900 563
rect 1924 557 1964 563
rect 1988 557 1996 563
rect 2084 557 2092 563
rect 2164 557 2300 563
rect 2436 557 2444 563
rect 2532 557 2684 563
rect 2756 557 2764 563
rect 2804 557 2940 563
rect 2948 557 3116 563
rect 3252 557 3356 563
rect 3364 557 3372 563
rect 3412 557 3436 563
rect 3492 557 3516 563
rect 3572 557 3580 563
rect 3668 557 3852 563
rect 317 544 323 556
rect 1117 544 1123 556
rect 1581 544 1587 556
rect 1821 544 1827 556
rect 3885 544 3891 556
rect 52 537 92 543
rect 100 537 124 543
rect 276 537 284 543
rect 388 537 396 543
rect 436 537 460 543
rect 500 537 636 543
rect 724 537 796 543
rect 932 537 940 543
rect 1204 537 1212 543
rect 1316 537 1324 543
rect 1332 537 1420 543
rect 1476 537 1532 543
rect 1796 537 1804 543
rect 1860 537 2268 543
rect 2301 537 2524 543
rect 100 517 188 523
rect 196 517 588 523
rect 596 517 1548 523
rect 1556 517 1852 523
rect 1876 517 1932 523
rect 2301 523 2307 537
rect 2532 537 2540 543
rect 2596 537 2668 543
rect 2788 537 2812 543
rect 2884 537 2972 543
rect 3012 537 3052 543
rect 3156 537 3580 543
rect 3588 537 3596 543
rect 3620 537 3628 543
rect 3716 537 3731 543
rect 3725 524 3731 537
rect 3764 537 3788 543
rect 3844 537 3868 543
rect 3940 537 3980 543
rect 4036 537 4060 543
rect 4084 537 4124 543
rect 3741 524 3747 536
rect 1997 517 2307 523
rect 196 497 220 503
rect 292 497 300 503
rect 308 497 892 503
rect 948 497 972 503
rect 1044 497 1596 503
rect 1997 503 2003 517
rect 2324 517 2348 523
rect 2692 517 2764 523
rect 2852 517 2892 523
rect 2980 517 3404 523
rect 3428 517 3468 523
rect 3508 517 3532 523
rect 3572 517 3708 523
rect 3780 517 3836 523
rect 3860 517 4108 523
rect 2557 504 2563 516
rect 1604 497 2003 503
rect 2132 497 2236 503
rect 2308 497 2428 503
rect 2436 497 2476 503
rect 2756 497 2876 503
rect 3028 497 3148 503
rect 3156 497 3356 503
rect 3364 497 3964 503
rect 3972 497 4076 503
rect 372 477 492 483
rect 644 477 668 483
rect 1044 477 1052 483
rect 1076 477 1228 483
rect 1412 477 1436 483
rect 1540 477 1628 483
rect 1636 477 2124 483
rect 2196 477 2204 483
rect 2292 477 2348 483
rect 2564 477 3004 483
rect 3012 477 3116 483
rect 3124 477 3324 483
rect 3348 477 3372 483
rect 3508 477 3852 483
rect 3956 477 3964 483
rect 3988 477 4012 483
rect 324 457 332 463
rect 468 457 1068 463
rect 1092 457 1132 463
rect 1421 457 1548 463
rect 996 437 1052 443
rect 1421 443 1427 457
rect 1556 457 2092 463
rect 2180 457 3244 463
rect 3284 457 3308 463
rect 3741 444 3747 456
rect 3773 444 3779 456
rect 1060 437 1427 443
rect 2036 437 2492 443
rect 1364 417 1500 423
rect 2292 417 2332 423
rect 2340 417 2348 423
rect 3524 417 3580 423
rect 4116 417 4188 423
rect 132 397 172 403
rect 580 397 604 403
rect 1204 397 1212 403
rect 1396 397 1452 403
rect 1668 397 1676 403
rect 1732 397 2364 403
rect 2628 397 2652 403
rect 2852 397 2940 403
rect 3316 397 3612 403
rect 3620 397 3692 403
rect 4148 397 4236 403
rect 148 377 300 383
rect 1300 377 1740 383
rect 2148 377 2156 383
rect 3108 377 3148 383
rect 3428 377 3452 383
rect 3492 377 3868 383
rect 3405 364 3411 376
rect 244 357 364 363
rect 1476 357 1724 363
rect 2356 357 2684 363
rect 3508 357 3516 363
rect 3540 357 3612 363
rect 52 337 76 343
rect 116 337 252 343
rect 413 337 419 356
rect 797 344 803 356
rect 436 337 460 343
rect 596 337 652 343
rect 1140 337 1148 343
rect 1540 337 1660 343
rect 1684 337 1804 343
rect 1972 337 2092 343
rect 2548 337 2556 343
rect 2948 337 2956 343
rect 3124 337 3756 343
rect 3780 337 3820 343
rect 1229 324 1235 336
rect 2205 324 2211 336
rect 2221 324 2227 336
rect 2893 324 2899 336
rect 3037 324 3043 336
rect 68 317 460 323
rect 644 317 652 323
rect 660 317 956 323
rect 964 317 1164 323
rect 1252 317 1260 323
rect 1444 317 1692 323
rect 2004 317 2028 323
rect 2244 317 2764 323
rect 2948 317 2988 323
rect 3092 317 3180 323
rect 3204 317 3212 323
rect 3252 317 3260 323
rect 3284 317 3292 323
rect 3348 317 3436 323
rect 3444 317 3564 323
rect 3588 317 3596 323
rect 3652 317 3708 323
rect 3716 317 3772 323
rect 3956 317 3980 323
rect 3805 304 3811 316
rect 516 297 1388 303
rect 1492 297 1500 303
rect 1620 297 1628 303
rect 1652 297 1676 303
rect 1924 297 2076 303
rect 2100 297 2172 303
rect 2212 297 2252 303
rect 2276 297 2860 303
rect 2868 297 3548 303
rect 3556 297 3724 303
rect 3860 297 3916 303
rect 4020 297 4220 303
rect 196 277 252 283
rect 292 277 332 283
rect 340 277 348 283
rect 708 277 732 283
rect 852 277 1180 283
rect 1188 277 2764 283
rect 2772 277 2812 283
rect 2820 277 2828 283
rect 2884 277 2908 283
rect 2948 277 2972 283
rect 3252 277 3260 283
rect 3348 277 4124 283
rect 228 257 396 263
rect 628 257 780 263
rect 868 257 924 263
rect 948 257 1260 263
rect 1268 257 1308 263
rect 1332 257 1372 263
rect 1508 257 1683 263
rect 868 237 1436 243
rect 1604 237 1612 243
rect 1636 237 1660 243
rect 1677 243 1683 257
rect 1700 257 1964 263
rect 1988 257 2044 263
rect 2164 257 2179 263
rect 2173 244 2179 257
rect 2420 257 2428 263
rect 2452 257 2508 263
rect 2532 257 2652 263
rect 2724 257 3132 263
rect 3140 257 3148 263
rect 3172 257 3292 263
rect 3476 257 3532 263
rect 3604 257 3676 263
rect 3700 257 3932 263
rect 3956 257 4012 263
rect 4036 257 4140 263
rect 1677 237 1772 243
rect 1860 237 2044 243
rect 2068 237 2092 243
rect 2388 237 2604 243
rect 2612 237 2940 243
rect 3268 237 3324 243
rect 3396 237 3484 243
rect 3556 237 3644 243
rect 3732 237 4092 243
rect 276 217 428 223
rect 1076 217 1084 223
rect 1188 217 1196 223
rect 1396 217 1532 223
rect 1636 217 1884 223
rect 1924 217 1932 223
rect 2772 217 2876 223
rect 2948 217 2956 223
rect 3188 217 3532 223
rect 3940 217 4188 223
rect 500 197 524 203
rect 964 197 1372 203
rect 1652 197 1884 203
rect 2260 197 2268 203
rect 2804 197 2828 203
rect 2868 197 3036 203
rect 3124 197 3212 203
rect 3604 197 3772 203
rect 4036 197 4044 203
rect 4116 197 4268 203
rect 180 177 204 183
rect 388 177 604 183
rect 740 177 1468 183
rect 1524 177 1612 183
rect 1636 177 1660 183
rect 1716 177 1772 183
rect 1876 177 1932 183
rect 2100 177 2124 183
rect 2164 177 2396 183
rect 2596 177 2636 183
rect 2708 177 2748 183
rect 2900 177 3260 183
rect 3268 177 3276 183
rect 3348 177 3356 183
rect 3588 177 3612 183
rect 3844 177 4124 183
rect 4196 177 4204 183
rect 4228 177 4323 183
rect 621 164 627 176
rect 3757 164 3763 176
rect 52 157 92 163
rect 164 157 332 163
rect 541 157 556 163
rect 644 157 908 163
rect 948 157 2316 163
rect 2468 157 2524 163
rect 2596 157 2844 163
rect 2916 157 2956 163
rect 2980 157 3452 163
rect 3524 157 3747 163
rect 100 137 140 143
rect 308 137 364 143
rect 372 137 636 143
rect 788 137 860 143
rect 884 137 892 143
rect 1108 137 1132 143
rect 1156 137 1180 143
rect 1204 137 1596 143
rect 1812 137 1836 143
rect 1924 137 1948 143
rect 1972 137 2108 143
rect 2308 137 2316 143
rect 2564 137 2604 143
rect 2692 137 3036 143
rect 3076 137 3148 143
rect 3188 137 3372 143
rect 3476 137 3692 143
rect 3741 143 3747 157
rect 3796 157 3820 163
rect 3837 144 3843 163
rect 3860 157 3868 163
rect 3956 157 4092 163
rect 4173 144 4179 156
rect 3741 137 3804 143
rect 4052 137 4060 143
rect 4189 137 4195 156
rect 4077 124 4083 136
rect 340 117 540 123
rect 564 117 828 123
rect 836 117 1251 123
rect 52 97 76 103
rect 132 97 396 103
rect 916 97 956 103
rect 1012 97 1020 103
rect 1060 97 1100 103
rect 1124 97 1164 103
rect 1204 97 1212 103
rect 1245 103 1251 117
rect 1284 117 1724 123
rect 1732 117 2556 123
rect 2916 117 2924 123
rect 2948 117 2956 123
rect 3012 117 3404 123
rect 3460 117 3484 123
rect 4196 117 4323 123
rect 1245 97 1564 103
rect 1764 97 1916 103
rect 2004 97 2044 103
rect 2212 97 2252 103
rect 2340 97 2364 103
rect 2756 97 2764 103
rect 2804 97 2860 103
rect 2964 97 2988 103
rect 3044 97 3084 103
rect 3172 97 3180 103
rect 3556 97 3571 103
rect 3828 97 3852 103
rect 4013 103 4019 116
rect 4004 97 4019 103
rect 4093 97 4099 116
rect 4148 97 4156 103
rect 4212 97 4236 103
rect 813 84 819 96
rect 1181 84 1187 96
rect 3101 84 3107 96
rect 900 77 1164 83
rect 1220 77 1244 83
rect 1476 77 1532 83
rect 1780 77 1804 83
rect 1956 77 2012 83
rect 2164 77 2476 83
rect 3060 57 3420 63
<< m4contact >>
rect 2524 2996 2532 3004
rect 1692 2976 1700 2984
rect 1372 2956 1380 2964
rect 1420 2956 1428 2964
rect 1532 2956 1540 2964
rect 1724 2956 1732 2964
rect 2988 2976 2996 2984
rect 3612 2976 3620 2984
rect 2796 2956 2804 2964
rect 3164 2956 3172 2964
rect 3468 2956 3476 2964
rect 3548 2956 3556 2964
rect 284 2936 292 2944
rect 1244 2936 1252 2944
rect 1500 2936 1508 2944
rect 1836 2936 1844 2944
rect 2876 2936 2884 2944
rect 2908 2936 2916 2944
rect 2972 2936 2980 2944
rect 3084 2936 3092 2944
rect 3212 2936 3220 2944
rect 3228 2936 3236 2944
rect 3276 2936 3284 2944
rect 3292 2936 3300 2944
rect 3612 2956 3620 2964
rect 4156 2956 4164 2964
rect 3660 2936 3668 2944
rect 732 2916 740 2924
rect 2332 2916 2340 2924
rect 2412 2916 2420 2924
rect 2940 2916 2948 2924
rect 3244 2916 3252 2924
rect 3676 2916 3684 2924
rect 668 2896 676 2904
rect 2460 2896 2468 2904
rect 2524 2896 2532 2904
rect 2700 2896 2708 2904
rect 2924 2896 2932 2904
rect 3868 2896 3876 2904
rect 3884 2896 3892 2904
rect 3980 2896 3988 2904
rect 4076 2896 4084 2904
rect 4156 2896 4164 2904
rect 1516 2876 1524 2884
rect 1564 2876 1572 2884
rect 2076 2876 2084 2884
rect 1532 2856 1540 2864
rect 2124 2856 2132 2864
rect 2316 2856 2324 2864
rect 2444 2856 2452 2864
rect 2572 2856 2580 2864
rect 1916 2836 1924 2844
rect 3420 2816 3428 2824
rect 1036 2796 1044 2804
rect 2636 2796 2644 2804
rect 3036 2796 3044 2804
rect 4108 2796 4116 2804
rect 4204 2796 4212 2804
rect 4092 2776 4100 2784
rect 524 2756 532 2764
rect 124 2736 132 2744
rect 812 2736 820 2744
rect 2092 2736 2100 2744
rect 3324 2736 3332 2744
rect 3980 2736 3988 2744
rect 4092 2736 4100 2744
rect 940 2716 948 2724
rect 2108 2716 2116 2724
rect 2140 2716 2148 2724
rect 2652 2716 2660 2724
rect 2764 2716 2772 2724
rect 3548 2716 3556 2724
rect 3612 2716 3620 2724
rect 3868 2716 3876 2724
rect 60 2676 68 2684
rect 588 2696 596 2704
rect 1004 2696 1012 2704
rect 1788 2696 1796 2704
rect 3676 2696 3684 2704
rect 828 2676 836 2684
rect 1020 2676 1028 2684
rect 2076 2676 2084 2684
rect 2092 2676 2100 2684
rect 3068 2676 3076 2684
rect 3580 2676 3588 2684
rect 3596 2676 3604 2684
rect 3948 2676 3956 2684
rect 3980 2676 3988 2684
rect 1276 2656 1284 2664
rect 1468 2656 1476 2664
rect 1532 2656 1540 2664
rect 1900 2656 1908 2664
rect 1932 2656 1940 2664
rect 2428 2656 2436 2664
rect 2524 2656 2532 2664
rect 2620 2656 2628 2664
rect 2700 2656 2708 2664
rect 2748 2656 2756 2664
rect 2764 2656 2772 2664
rect 524 2636 532 2644
rect 940 2636 948 2644
rect 972 2636 980 2644
rect 988 2636 996 2644
rect 1660 2636 1668 2644
rect 1756 2636 1764 2644
rect 1852 2636 1860 2644
rect 1932 2636 1940 2644
rect 2268 2636 2276 2644
rect 3260 2636 3268 2644
rect 284 2616 292 2624
rect 812 2616 820 2624
rect 908 2616 916 2624
rect 1116 2616 1124 2624
rect 1820 2616 1828 2624
rect 1900 2616 1908 2624
rect 1996 2616 2004 2624
rect 2108 2616 2116 2624
rect 2236 2616 2244 2624
rect 2444 2616 2452 2624
rect 2556 2616 2564 2624
rect 2940 2616 2948 2624
rect 2972 2616 2980 2624
rect 3148 2616 3156 2624
rect 364 2596 372 2604
rect 652 2596 660 2604
rect 860 2596 868 2604
rect 1564 2596 1572 2604
rect 1868 2596 1876 2604
rect 1884 2596 1892 2604
rect 2316 2596 2324 2604
rect 2716 2596 2724 2604
rect 3052 2596 3060 2604
rect 3068 2596 3076 2604
rect 3084 2596 3092 2604
rect 3100 2596 3108 2604
rect 3164 2596 3172 2604
rect 3180 2596 3188 2604
rect 3388 2596 3396 2604
rect 3500 2596 3508 2604
rect 3516 2596 3524 2604
rect 3548 2596 3556 2604
rect 3916 2596 3924 2604
rect 1260 2576 1268 2584
rect 1484 2576 1492 2584
rect 1836 2576 1844 2584
rect 2060 2576 2068 2584
rect 2076 2576 2084 2584
rect 2796 2576 2804 2584
rect 2908 2576 2916 2584
rect 3004 2576 3012 2584
rect 3020 2576 3028 2584
rect 3484 2576 3492 2584
rect 3820 2576 3828 2584
rect 508 2556 516 2564
rect 556 2556 564 2564
rect 844 2556 852 2564
rect 1244 2556 1252 2564
rect 1468 2556 1476 2564
rect 1548 2556 1556 2564
rect 1580 2556 1588 2564
rect 1804 2556 1812 2564
rect 3212 2556 3220 2564
rect 3964 2556 3972 2564
rect 668 2536 676 2544
rect 908 2536 916 2544
rect 1052 2536 1060 2544
rect 1068 2536 1076 2544
rect 1996 2536 2004 2544
rect 2028 2536 2036 2544
rect 2092 2536 2100 2544
rect 2764 2536 2772 2544
rect 2924 2536 2932 2544
rect 2988 2536 2996 2544
rect 3036 2536 3044 2544
rect 3052 2536 3060 2544
rect 3068 2536 3076 2544
rect 3340 2536 3348 2544
rect 3404 2536 3412 2544
rect 3452 2536 3460 2544
rect 3500 2536 3508 2544
rect 3564 2536 3572 2544
rect 3628 2536 3636 2544
rect 3756 2536 3764 2544
rect 3868 2536 3876 2544
rect 3900 2536 3908 2544
rect 4044 2536 4052 2544
rect 4172 2536 4180 2544
rect 1804 2516 1812 2524
rect 1836 2516 1844 2524
rect 1900 2516 1908 2524
rect 2108 2516 2116 2524
rect 2476 2516 2484 2524
rect 2540 2516 2548 2524
rect 2572 2516 2580 2524
rect 2604 2516 2612 2524
rect 2716 2516 2724 2524
rect 2764 2516 2772 2524
rect 60 2496 68 2504
rect 124 2496 132 2504
rect 892 2496 900 2504
rect 988 2496 996 2504
rect 1132 2496 1140 2504
rect 1356 2496 1364 2504
rect 1420 2496 1428 2504
rect 1468 2496 1476 2504
rect 1756 2496 1764 2504
rect 2252 2496 2260 2504
rect 2556 2496 2564 2504
rect 2716 2496 2724 2504
rect 3052 2496 3060 2504
rect 3500 2496 3508 2504
rect 3532 2496 3540 2504
rect 3596 2496 3604 2504
rect 3628 2496 3636 2504
rect 3692 2496 3700 2504
rect 3788 2496 3796 2504
rect 3836 2496 3844 2504
rect 4140 2496 4148 2504
rect 588 2476 596 2484
rect 1500 2476 1508 2484
rect 1660 2476 1668 2484
rect 2076 2476 2084 2484
rect 2172 2476 2180 2484
rect 2572 2476 2580 2484
rect 652 2456 660 2464
rect 1612 2456 1620 2464
rect 1820 2456 1828 2464
rect 1916 2456 1924 2464
rect 1980 2456 1988 2464
rect 2716 2456 2724 2464
rect 2892 2456 2900 2464
rect 3004 2456 3012 2464
rect 3308 2456 3316 2464
rect 3356 2456 3364 2464
rect 3180 2436 3188 2444
rect 3852 2436 3860 2444
rect 956 2416 964 2424
rect 1580 2416 1588 2424
rect 636 2396 644 2404
rect 764 2396 772 2404
rect 1020 2396 1028 2404
rect 2332 2396 2340 2404
rect 3500 2396 3508 2404
rect 3644 2396 3652 2404
rect 2060 2376 2068 2384
rect 2444 2376 2452 2384
rect 2492 2376 2500 2384
rect 2620 2376 2628 2384
rect 2876 2376 2884 2384
rect 3612 2376 3620 2384
rect 188 2356 196 2364
rect 268 2356 276 2364
rect 476 2356 484 2364
rect 620 2356 628 2364
rect 652 2356 660 2364
rect 1020 2356 1028 2364
rect 1116 2356 1124 2364
rect 1532 2356 1540 2364
rect 1628 2356 1636 2364
rect 2268 2356 2276 2364
rect 2908 2356 2916 2364
rect 3100 2356 3108 2364
rect 3644 2356 3652 2364
rect 3676 2356 3684 2364
rect 3932 2356 3940 2364
rect 220 2336 228 2344
rect 636 2336 644 2344
rect 972 2336 980 2344
rect 1308 2336 1316 2344
rect 1692 2336 1700 2344
rect 2060 2336 2068 2344
rect 2460 2336 2468 2344
rect 348 2316 356 2324
rect 428 2316 436 2324
rect 476 2316 484 2324
rect 1020 2316 1028 2324
rect 1084 2316 1092 2324
rect 1180 2316 1188 2324
rect 2860 2336 2868 2344
rect 2940 2336 2948 2344
rect 2956 2336 2964 2344
rect 3900 2336 3908 2344
rect 2540 2316 2548 2324
rect 2572 2316 2580 2324
rect 2780 2316 2788 2324
rect 3692 2316 3700 2324
rect 3884 2316 3892 2324
rect 4156 2316 4164 2324
rect 188 2276 196 2284
rect 1436 2296 1444 2304
rect 3708 2296 3716 2304
rect 524 2276 532 2284
rect 604 2276 612 2284
rect 716 2276 724 2284
rect 828 2276 836 2284
rect 2124 2276 2132 2284
rect 2140 2276 2148 2284
rect 2188 2276 2196 2284
rect 2252 2276 2260 2284
rect 2348 2276 2356 2284
rect 2364 2276 2372 2284
rect 2428 2276 2436 2284
rect 3196 2276 3204 2284
rect 3660 2276 3668 2284
rect 4124 2276 4132 2284
rect 348 2256 356 2264
rect 812 2256 820 2264
rect 1020 2256 1028 2264
rect 1052 2256 1060 2264
rect 1404 2256 1412 2264
rect 1468 2256 1476 2264
rect 1532 2256 1540 2264
rect 1548 2256 1556 2264
rect 1676 2256 1684 2264
rect 1724 2256 1732 2264
rect 1772 2256 1780 2264
rect 1996 2256 2004 2264
rect 2492 2256 2500 2264
rect 2524 2256 2532 2264
rect 2812 2256 2820 2264
rect 2908 2256 2916 2264
rect 3068 2256 3076 2264
rect 3612 2256 3620 2264
rect 3932 2256 3940 2264
rect 4076 2256 4084 2264
rect 828 2236 836 2244
rect 1100 2236 1108 2244
rect 1132 2236 1140 2244
rect 1292 2236 1300 2244
rect 1740 2236 1748 2244
rect 2076 2236 2084 2244
rect 2540 2236 2548 2244
rect 2556 2236 2564 2244
rect 2668 2236 2676 2244
rect 2796 2236 2804 2244
rect 3228 2236 3236 2244
rect 3308 2236 3316 2244
rect 3564 2236 3572 2244
rect 1340 2216 1348 2224
rect 1708 2216 1716 2224
rect 2300 2216 2308 2224
rect 2460 2216 2468 2224
rect 3516 2216 3524 2224
rect 3980 2236 3988 2244
rect 4188 2236 4196 2244
rect 3836 2216 3844 2224
rect 3916 2216 3924 2224
rect 3932 2216 3940 2224
rect 252 2196 260 2204
rect 492 2196 500 2204
rect 524 2196 532 2204
rect 956 2196 964 2204
rect 1340 2196 1348 2204
rect 2364 2196 2372 2204
rect 2444 2196 2452 2204
rect 2844 2196 2852 2204
rect 3820 2196 3828 2204
rect 4012 2196 4020 2204
rect 796 2176 804 2184
rect 1020 2176 1028 2184
rect 1212 2176 1220 2184
rect 1228 2176 1236 2184
rect 1324 2176 1332 2184
rect 1772 2176 1780 2184
rect 1900 2176 1908 2184
rect 1916 2176 1924 2184
rect 1964 2176 1972 2184
rect 2012 2176 2020 2184
rect 3020 2176 3028 2184
rect 3148 2176 3156 2184
rect 3564 2176 3572 2184
rect 3948 2176 3956 2184
rect 4092 2176 4100 2184
rect 4140 2176 4148 2184
rect 108 2156 116 2164
rect 220 2156 228 2164
rect 284 2156 292 2164
rect 588 2156 596 2164
rect 620 2156 628 2164
rect 1356 2156 1364 2164
rect 1676 2156 1684 2164
rect 1788 2156 1796 2164
rect 1804 2156 1812 2164
rect 2028 2156 2036 2164
rect 2060 2156 2068 2164
rect 2524 2156 2532 2164
rect 2620 2156 2628 2164
rect 3084 2156 3092 2164
rect 268 2136 276 2144
rect 844 2136 852 2144
rect 1068 2136 1076 2144
rect 1164 2136 1172 2144
rect 1500 2136 1508 2144
rect 1580 2136 1588 2144
rect 2572 2136 2580 2144
rect 2668 2136 2676 2144
rect 2764 2136 2772 2144
rect 3548 2136 3556 2144
rect 3580 2136 3588 2144
rect 3708 2136 3716 2144
rect 3836 2136 3844 2144
rect 3884 2136 3892 2144
rect 3916 2136 3924 2144
rect 476 2116 484 2124
rect 540 2116 548 2124
rect 588 2116 596 2124
rect 700 2116 708 2124
rect 748 2116 756 2124
rect 780 2116 788 2124
rect 876 2116 884 2124
rect 1052 2116 1060 2124
rect 1196 2116 1204 2124
rect 1308 2116 1316 2124
rect 2092 2116 2100 2124
rect 2156 2116 2164 2124
rect 2188 2116 2196 2124
rect 2316 2116 2324 2124
rect 2380 2116 2388 2124
rect 2476 2116 2484 2124
rect 2988 2116 2996 2124
rect 3004 2116 3012 2124
rect 3132 2116 3140 2124
rect 3388 2116 3396 2124
rect 3580 2116 3588 2124
rect 3596 2116 3604 2124
rect 1564 2096 1572 2104
rect 1836 2096 1844 2104
rect 2604 2096 2612 2104
rect 2892 2096 2900 2104
rect 2956 2096 2964 2104
rect 2972 2096 2980 2104
rect 3100 2096 3108 2104
rect 3356 2096 3364 2104
rect 4124 2096 4132 2104
rect 684 2076 692 2084
rect 1020 2076 1028 2084
rect 1260 2076 1268 2084
rect 1548 2076 1556 2084
rect 1740 2076 1748 2084
rect 1820 2076 1828 2084
rect 1996 2076 2004 2084
rect 2092 2076 2100 2084
rect 2588 2076 2596 2084
rect 2652 2076 2660 2084
rect 3788 2076 3796 2084
rect 588 2056 596 2064
rect 1100 2036 1108 2044
rect 1484 2036 1492 2044
rect 1596 2036 1604 2044
rect 1708 2056 1716 2064
rect 1980 2056 1988 2064
rect 2028 2056 2036 2064
rect 2124 2056 2132 2064
rect 2940 2056 2948 2064
rect 3580 2056 3588 2064
rect 3820 2056 3828 2064
rect 2300 2036 2308 2044
rect 3004 2036 3012 2044
rect 3020 2036 3028 2044
rect 1692 2016 1700 2024
rect 2028 2016 2036 2024
rect 2092 2016 2100 2024
rect 2124 2016 2132 2024
rect 3340 2016 3348 2024
rect 3788 2016 3796 2024
rect 236 1996 244 2004
rect 2412 1996 2420 2004
rect 2444 1996 2452 2004
rect 2556 1996 2564 2004
rect 2732 1996 2740 2004
rect 748 1976 756 1984
rect 4012 1976 4020 1984
rect 636 1956 644 1964
rect 1868 1956 1876 1964
rect 2156 1956 2164 1964
rect 2236 1956 2244 1964
rect 2268 1956 2276 1964
rect 2300 1956 2308 1964
rect 2364 1956 2372 1964
rect 2460 1956 2468 1964
rect 2508 1956 2516 1964
rect 2556 1956 2564 1964
rect 3452 1956 3460 1964
rect 236 1936 244 1944
rect 716 1936 724 1944
rect 1804 1936 1812 1944
rect 2508 1936 2516 1944
rect 2588 1936 2596 1944
rect 2668 1936 2676 1944
rect 2828 1936 2836 1944
rect 3532 1936 3540 1944
rect 3724 1936 3732 1944
rect 3868 1936 3876 1944
rect 4092 1936 4100 1944
rect 524 1916 532 1924
rect 828 1916 836 1924
rect 1244 1916 1252 1924
rect 1788 1916 1796 1924
rect 1980 1916 1988 1924
rect 2412 1916 2420 1924
rect 2428 1916 2436 1924
rect 2460 1916 2468 1924
rect 2524 1916 2532 1924
rect 2780 1916 2788 1924
rect 2812 1916 2820 1924
rect 2972 1916 2980 1924
rect 3340 1916 3348 1924
rect 3884 1916 3892 1924
rect 4108 1916 4116 1924
rect 140 1896 148 1904
rect 300 1896 308 1904
rect 812 1896 820 1904
rect 828 1896 836 1904
rect 1852 1896 1860 1904
rect 2108 1896 2116 1904
rect 2908 1896 2916 1904
rect 124 1876 132 1884
rect 732 1876 740 1884
rect 1164 1876 1172 1884
rect 1196 1876 1204 1884
rect 1244 1876 1252 1884
rect 1260 1876 1268 1884
rect 1308 1876 1316 1884
rect 1340 1876 1348 1884
rect 1356 1876 1364 1884
rect 1820 1876 1828 1884
rect 1852 1876 1860 1884
rect 1884 1876 1892 1884
rect 1900 1876 1908 1884
rect 1916 1876 1924 1884
rect 1948 1876 1956 1884
rect 1996 1876 2004 1884
rect 2508 1876 2516 1884
rect 2636 1876 2644 1884
rect 3708 1876 3716 1884
rect 204 1856 212 1864
rect 348 1856 356 1864
rect 444 1856 452 1864
rect 716 1856 724 1864
rect 988 1856 996 1864
rect 1292 1856 1300 1864
rect 1404 1856 1412 1864
rect 2812 1856 2820 1864
rect 2956 1856 2964 1864
rect 3308 1856 3316 1864
rect 3372 1856 3380 1864
rect 3852 1856 3860 1864
rect 4012 1856 4020 1864
rect 4108 1856 4116 1864
rect 380 1836 388 1844
rect 812 1836 820 1844
rect 1228 1836 1236 1844
rect 1452 1836 1460 1844
rect 1500 1836 1508 1844
rect 1596 1836 1604 1844
rect 1612 1836 1620 1844
rect 1772 1836 1780 1844
rect 2124 1836 2132 1844
rect 2140 1836 2148 1844
rect 2156 1836 2164 1844
rect 2220 1836 2228 1844
rect 2268 1836 2276 1844
rect 2556 1836 2564 1844
rect 780 1816 788 1824
rect 1692 1816 1700 1824
rect 2268 1816 2276 1824
rect 2460 1816 2468 1824
rect 3452 1816 3460 1824
rect 284 1796 292 1804
rect 1164 1796 1172 1804
rect 1324 1796 1332 1804
rect 1676 1796 1684 1804
rect 2380 1796 2388 1804
rect 2508 1796 2516 1804
rect 3084 1796 3092 1804
rect 3388 1796 3396 1804
rect 364 1776 372 1784
rect 684 1776 692 1784
rect 796 1776 804 1784
rect 1180 1776 1188 1784
rect 204 1756 212 1764
rect 252 1756 260 1764
rect 460 1756 468 1764
rect 684 1756 692 1764
rect 780 1756 788 1764
rect 972 1756 980 1764
rect 1052 1756 1060 1764
rect 1068 1756 1076 1764
rect 1196 1756 1204 1764
rect 1340 1756 1348 1764
rect 2012 1776 2020 1784
rect 2220 1776 2228 1784
rect 2876 1776 2884 1784
rect 3004 1776 3012 1784
rect 3212 1776 3220 1784
rect 3660 1776 3668 1784
rect 4028 1776 4036 1784
rect 1628 1756 1636 1764
rect 1676 1756 1684 1764
rect 2156 1756 2164 1764
rect 2204 1756 2212 1764
rect 2300 1756 2308 1764
rect 2748 1756 2756 1764
rect 2876 1756 2884 1764
rect 2892 1756 2900 1764
rect 3516 1756 3524 1764
rect 652 1736 660 1744
rect 1212 1736 1220 1744
rect 1324 1736 1332 1744
rect 1484 1736 1492 1744
rect 1500 1736 1508 1744
rect 1612 1736 1620 1744
rect 1900 1736 1908 1744
rect 2444 1736 2452 1744
rect 2492 1736 2500 1744
rect 2572 1736 2580 1744
rect 2908 1736 2916 1744
rect 3228 1736 3236 1744
rect 3404 1736 3412 1744
rect 3852 1756 3860 1764
rect 3868 1756 3876 1764
rect 4124 1756 4132 1764
rect 4044 1736 4052 1744
rect 4140 1736 4148 1744
rect 924 1716 932 1724
rect 1276 1716 1284 1724
rect 2252 1716 2260 1724
rect 2604 1716 2612 1724
rect 3244 1716 3252 1724
rect 3276 1716 3284 1724
rect 3340 1716 3348 1724
rect 3388 1716 3396 1724
rect 1292 1696 1300 1704
rect 1772 1696 1780 1704
rect 1788 1696 1796 1704
rect 2108 1696 2116 1704
rect 2156 1696 2164 1704
rect 2204 1696 2212 1704
rect 3020 1696 3028 1704
rect 3100 1696 3108 1704
rect 3292 1696 3300 1704
rect 3372 1696 3380 1704
rect 4028 1696 4036 1704
rect 764 1676 772 1684
rect 1356 1676 1364 1684
rect 1404 1676 1412 1684
rect 1484 1676 1492 1684
rect 1916 1676 1924 1684
rect 1932 1676 1940 1684
rect 1948 1676 1956 1684
rect 1996 1676 2004 1684
rect 2476 1676 2484 1684
rect 908 1656 916 1664
rect 1036 1656 1044 1664
rect 1660 1656 1668 1664
rect 2140 1656 2148 1664
rect 2236 1656 2244 1664
rect 2300 1656 2308 1664
rect 2588 1656 2596 1664
rect 3084 1676 3092 1684
rect 3212 1676 3220 1684
rect 3260 1656 3268 1664
rect 3340 1676 3348 1684
rect 3676 1676 3684 1684
rect 3388 1656 3396 1664
rect 3516 1656 3524 1664
rect 3788 1656 3796 1664
rect 508 1636 516 1644
rect 812 1636 820 1644
rect 1964 1636 1972 1644
rect 3580 1636 3588 1644
rect 3692 1636 3700 1644
rect 780 1616 788 1624
rect 1196 1616 1204 1624
rect 2348 1616 2356 1624
rect 2364 1616 2372 1624
rect 3516 1616 3524 1624
rect 3580 1616 3588 1624
rect 3628 1616 3636 1624
rect 3788 1616 3796 1624
rect 4172 1616 4180 1624
rect 140 1596 148 1604
rect 236 1596 244 1604
rect 1388 1596 1396 1604
rect 1868 1596 1876 1604
rect 2396 1596 2404 1604
rect 2428 1596 2436 1604
rect 2524 1596 2532 1604
rect 2556 1596 2564 1604
rect 2684 1596 2692 1604
rect 3436 1596 3444 1604
rect 3612 1596 3620 1604
rect 4172 1596 4180 1604
rect 124 1576 132 1584
rect 1516 1576 1524 1584
rect 1724 1576 1732 1584
rect 2428 1576 2436 1584
rect 2700 1576 2708 1584
rect 3628 1576 3636 1584
rect 3740 1576 3748 1584
rect 1580 1556 1588 1564
rect 1692 1556 1700 1564
rect 2028 1556 2036 1564
rect 2076 1556 2084 1564
rect 2204 1556 2212 1564
rect 2236 1556 2244 1564
rect 2860 1556 2868 1564
rect 3116 1556 3124 1564
rect 3628 1556 3636 1564
rect 3692 1556 3700 1564
rect 412 1536 420 1544
rect 1420 1536 1428 1544
rect 2396 1536 2404 1544
rect 2412 1536 2420 1544
rect 2572 1536 2580 1544
rect 3068 1536 3076 1544
rect 3420 1536 3428 1544
rect 3724 1536 3732 1544
rect 748 1516 756 1524
rect 1372 1516 1380 1524
rect 1420 1516 1428 1524
rect 1708 1516 1716 1524
rect 2268 1516 2276 1524
rect 2316 1516 2324 1524
rect 2348 1516 2356 1524
rect 2860 1516 2868 1524
rect 2908 1516 2916 1524
rect 3148 1516 3156 1524
rect 3340 1516 3348 1524
rect 4156 1516 4164 1524
rect 412 1496 420 1504
rect 492 1496 500 1504
rect 1084 1496 1092 1504
rect 1404 1496 1412 1504
rect 1468 1496 1476 1504
rect 2252 1496 2260 1504
rect 2428 1496 2436 1504
rect 2604 1496 2612 1504
rect 2956 1496 2964 1504
rect 3452 1496 3460 1504
rect 4124 1496 4132 1504
rect 12 1476 20 1484
rect 236 1476 244 1484
rect 252 1456 260 1464
rect 332 1476 340 1484
rect 620 1476 628 1484
rect 844 1476 852 1484
rect 892 1476 900 1484
rect 1308 1476 1316 1484
rect 1564 1476 1572 1484
rect 1708 1476 1716 1484
rect 1820 1476 1828 1484
rect 2012 1476 2020 1484
rect 2060 1476 2068 1484
rect 2076 1476 2084 1484
rect 2604 1476 2612 1484
rect 2732 1476 2740 1484
rect 3132 1476 3140 1484
rect 3244 1476 3252 1484
rect 3532 1476 3540 1484
rect 3580 1476 3588 1484
rect 3612 1476 3620 1484
rect 3724 1476 3732 1484
rect 3932 1476 3940 1484
rect 3948 1476 3956 1484
rect 4220 1476 4228 1484
rect 380 1456 388 1464
rect 396 1456 404 1464
rect 1676 1456 1684 1464
rect 1948 1456 1956 1464
rect 2508 1456 2516 1464
rect 12 1436 20 1444
rect 892 1436 900 1444
rect 1404 1436 1412 1444
rect 2220 1436 2228 1444
rect 2476 1436 2484 1444
rect 2556 1436 2564 1444
rect 2604 1456 2612 1464
rect 2892 1456 2900 1464
rect 3100 1456 3108 1464
rect 3276 1456 3284 1464
rect 3708 1456 3716 1464
rect 3788 1456 3796 1464
rect 428 1416 436 1424
rect 1356 1416 1364 1424
rect 1724 1416 1732 1424
rect 1756 1416 1764 1424
rect 2300 1416 2308 1424
rect 892 1396 900 1404
rect 1228 1396 1236 1404
rect 2028 1396 2036 1404
rect 2076 1396 2084 1404
rect 412 1376 420 1384
rect 924 1376 932 1384
rect 1084 1376 1092 1384
rect 1324 1376 1332 1384
rect 1452 1376 1460 1384
rect 444 1356 452 1364
rect 492 1356 500 1364
rect 2572 1416 2580 1424
rect 2652 1416 2660 1424
rect 2876 1416 2884 1424
rect 2892 1416 2900 1424
rect 3100 1416 3108 1424
rect 3580 1416 3588 1424
rect 3692 1416 3700 1424
rect 2460 1396 2468 1404
rect 2476 1396 2484 1404
rect 2684 1396 2692 1404
rect 2812 1396 2820 1404
rect 2828 1396 2836 1404
rect 3340 1396 3348 1404
rect 3532 1396 3540 1404
rect 3548 1396 3556 1404
rect 2140 1376 2148 1384
rect 2172 1376 2180 1384
rect 2316 1376 2324 1384
rect 2348 1376 2356 1384
rect 2732 1376 2740 1384
rect 2908 1376 2916 1384
rect 2956 1376 2964 1384
rect 2988 1376 2996 1384
rect 3052 1376 3060 1384
rect 3228 1376 3236 1384
rect 3340 1376 3348 1384
rect 3468 1376 3476 1384
rect 3612 1376 3620 1384
rect 3692 1376 3700 1384
rect 1500 1356 1508 1364
rect 1580 1356 1588 1364
rect 1660 1356 1668 1364
rect 1996 1356 2004 1364
rect 2028 1356 2036 1364
rect 2124 1356 2132 1364
rect 2284 1356 2292 1364
rect 2396 1356 2404 1364
rect 2444 1356 2452 1364
rect 2540 1356 2548 1364
rect 2572 1356 2580 1364
rect 2716 1356 2724 1364
rect 2748 1356 2756 1364
rect 2780 1356 2788 1364
rect 3068 1356 3076 1364
rect 3452 1356 3460 1364
rect 3772 1356 3780 1364
rect 4092 1356 4100 1364
rect 4156 1356 4164 1364
rect 364 1336 372 1344
rect 508 1336 516 1344
rect 812 1336 820 1344
rect 1356 1336 1364 1344
rect 1484 1336 1492 1344
rect 1884 1336 1892 1344
rect 1900 1336 1908 1344
rect 2268 1336 2276 1344
rect 2556 1336 2564 1344
rect 2876 1336 2884 1344
rect 2892 1336 2900 1344
rect 3436 1336 3444 1344
rect 3836 1336 3844 1344
rect 3964 1336 3972 1344
rect 4092 1336 4100 1344
rect 428 1316 436 1324
rect 476 1316 484 1324
rect 1372 1316 1380 1324
rect 1836 1316 1844 1324
rect 2012 1316 2020 1324
rect 2428 1316 2436 1324
rect 3724 1316 3732 1324
rect 4140 1316 4148 1324
rect 92 1296 100 1304
rect 668 1296 676 1304
rect 796 1296 804 1304
rect 924 1296 932 1304
rect 1084 1296 1092 1304
rect 1292 1296 1300 1304
rect 1820 1296 1828 1304
rect 2028 1296 2036 1304
rect 2060 1296 2068 1304
rect 2140 1296 2148 1304
rect 2396 1296 2404 1304
rect 2540 1296 2548 1304
rect 2588 1296 2596 1304
rect 2604 1296 2612 1304
rect 2892 1296 2900 1304
rect 2908 1296 2916 1304
rect 3340 1296 3348 1304
rect 3484 1296 3492 1304
rect 3772 1296 3780 1304
rect 4204 1296 4212 1304
rect 972 1276 980 1284
rect 1228 1276 1236 1284
rect 1340 1276 1348 1284
rect 1468 1276 1476 1284
rect 1516 1276 1524 1284
rect 1580 1276 1588 1284
rect 1724 1276 1732 1284
rect 2076 1276 2084 1284
rect 2172 1276 2180 1284
rect 540 1256 548 1264
rect 2188 1256 2196 1264
rect 2220 1256 2228 1264
rect 2892 1276 2900 1284
rect 3388 1276 3396 1284
rect 2940 1256 2948 1264
rect 2988 1256 2996 1264
rect 3164 1256 3172 1264
rect 3212 1256 3220 1264
rect 3484 1256 3492 1264
rect 988 1236 996 1244
rect 2060 1236 2068 1244
rect 2700 1236 2708 1244
rect 4220 1236 4228 1244
rect 3500 1216 3508 1224
rect 3644 1216 3652 1224
rect 1100 1196 1108 1204
rect 2220 1196 2228 1204
rect 2476 1196 2484 1204
rect 2732 1196 2740 1204
rect 4060 1196 4068 1204
rect 780 1176 788 1184
rect 2844 1176 2852 1184
rect 252 1156 260 1164
rect 1020 1156 1028 1164
rect 1708 1156 1716 1164
rect 1916 1156 1924 1164
rect 2268 1156 2276 1164
rect 2508 1156 2516 1164
rect 2908 1156 2916 1164
rect 3356 1156 3364 1164
rect 3628 1156 3636 1164
rect 3852 1156 3860 1164
rect 4188 1156 4196 1164
rect 380 1136 388 1144
rect 460 1136 468 1144
rect 652 1136 660 1144
rect 1692 1136 1700 1144
rect 1996 1136 2004 1144
rect 2252 1136 2260 1144
rect 2284 1136 2292 1144
rect 2540 1136 2548 1144
rect 3372 1136 3380 1144
rect 3580 1136 3588 1144
rect 3628 1136 3636 1144
rect 3900 1136 3908 1144
rect 284 1116 292 1124
rect 668 1116 676 1124
rect 764 1116 772 1124
rect 988 1116 996 1124
rect 1084 1116 1092 1124
rect 1292 1116 1300 1124
rect 1372 1116 1380 1124
rect 1804 1116 1812 1124
rect 2620 1116 2628 1124
rect 2780 1116 2788 1124
rect 3180 1116 3188 1124
rect 3404 1116 3412 1124
rect 3420 1116 3428 1124
rect 3756 1116 3764 1124
rect 4204 1116 4212 1124
rect 652 1096 660 1104
rect 1132 1096 1140 1104
rect 2012 1096 2020 1104
rect 2156 1096 2164 1104
rect 2284 1096 2292 1104
rect 2444 1096 2452 1104
rect 2716 1096 2724 1104
rect 2956 1096 2964 1104
rect 3308 1096 3316 1104
rect 3404 1096 3412 1104
rect 3564 1096 3572 1104
rect 3884 1096 3892 1104
rect 156 1076 164 1084
rect 268 1076 276 1084
rect 396 1076 404 1084
rect 556 1076 564 1084
rect 716 1076 724 1084
rect 812 1076 820 1084
rect 1116 1076 1124 1084
rect 1676 1076 1684 1084
rect 1836 1076 1844 1084
rect 1900 1076 1908 1084
rect 2172 1076 2180 1084
rect 2204 1076 2212 1084
rect 2460 1076 2468 1084
rect 2556 1076 2564 1084
rect 2604 1076 2612 1084
rect 2860 1076 2868 1084
rect 3692 1076 3700 1084
rect 3788 1076 3796 1084
rect 3836 1076 3844 1084
rect 4012 1076 4020 1084
rect 4108 1076 4116 1084
rect 4204 1076 4212 1084
rect 140 1056 148 1064
rect 188 1056 196 1064
rect 252 1056 260 1064
rect 540 1056 548 1064
rect 572 1056 580 1064
rect 620 1056 628 1064
rect 1036 1056 1044 1064
rect 1212 1056 1220 1064
rect 1340 1056 1348 1064
rect 1484 1056 1492 1064
rect 1596 1056 1604 1064
rect 1964 1056 1972 1064
rect 2572 1056 2580 1064
rect 2588 1056 2596 1064
rect 2684 1056 2692 1064
rect 2860 1056 2868 1064
rect 3228 1056 3236 1064
rect 3372 1056 3380 1064
rect 92 1036 100 1044
rect 140 1016 148 1024
rect 780 1036 788 1044
rect 796 1036 804 1044
rect 956 1036 964 1044
rect 2172 1036 2180 1044
rect 2828 1036 2836 1044
rect 2844 1036 2852 1044
rect 3004 1036 3012 1044
rect 3260 1036 3268 1044
rect 3388 1036 3396 1044
rect 3692 1036 3700 1044
rect 4140 1036 4148 1044
rect 1244 1016 1252 1024
rect 1500 1016 1508 1024
rect 1564 1016 1572 1024
rect 1644 1016 1652 1024
rect 4140 1016 4148 1024
rect 588 996 596 1004
rect 908 996 916 1004
rect 2572 996 2580 1004
rect 2620 996 2628 1004
rect 2716 996 2724 1004
rect 124 976 132 984
rect 252 976 260 984
rect 748 976 756 984
rect 764 976 772 984
rect 828 976 836 984
rect 924 976 932 984
rect 988 976 996 984
rect 1676 976 1684 984
rect 2860 996 2868 1004
rect 3164 996 3172 1004
rect 3532 996 3540 1004
rect 4172 996 4180 1004
rect 4188 996 4196 1004
rect 2956 976 2964 984
rect 2972 976 2980 984
rect 3036 976 3044 984
rect 3292 976 3300 984
rect 3308 976 3316 984
rect 140 956 148 964
rect 172 956 180 964
rect 428 956 436 964
rect 492 956 500 964
rect 508 956 516 964
rect 620 956 628 964
rect 1052 956 1060 964
rect 1356 956 1364 964
rect 1484 956 1492 964
rect 2140 956 2148 964
rect 2188 956 2196 964
rect 2364 956 2372 964
rect 2492 956 2500 964
rect 316 936 324 944
rect 1436 936 1444 944
rect 1820 936 1828 944
rect 1964 936 1972 944
rect 1980 936 1988 944
rect 2028 936 2036 944
rect 2124 936 2132 944
rect 2732 956 2740 964
rect 2828 956 2836 964
rect 3196 956 3204 964
rect 3228 956 3236 964
rect 3468 956 3476 964
rect 3484 956 3492 964
rect 3564 956 3572 964
rect 3612 956 3620 964
rect 3660 956 3668 964
rect 3692 956 3700 964
rect 4108 956 4116 964
rect 2540 936 2548 944
rect 2860 936 2868 944
rect 2876 936 2884 944
rect 3788 936 3796 944
rect 3804 936 3812 944
rect 3916 936 3924 944
rect 60 916 68 924
rect 748 916 756 924
rect 1292 916 1300 924
rect 1372 916 1380 924
rect 1388 916 1396 924
rect 1980 916 1988 924
rect 2012 916 2020 924
rect 2044 916 2052 924
rect 2268 916 2276 924
rect 2316 916 2324 924
rect 2348 916 2356 924
rect 2428 916 2436 924
rect 2444 916 2452 924
rect 2988 916 2996 924
rect 124 896 132 904
rect 332 896 340 904
rect 572 896 580 904
rect 860 896 868 904
rect 972 896 980 904
rect 1020 896 1028 904
rect 1132 896 1140 904
rect 1244 896 1252 904
rect 1468 896 1476 904
rect 1612 896 1620 904
rect 700 876 708 884
rect 1836 896 1844 904
rect 1852 896 1860 904
rect 2300 896 2308 904
rect 2556 896 2564 904
rect 2636 896 2644 904
rect 3052 896 3060 904
rect 3436 896 3444 904
rect 3612 916 3620 924
rect 4044 916 4052 924
rect 3516 896 3524 904
rect 3532 896 3540 904
rect 3548 896 3556 904
rect 3612 896 3620 904
rect 3644 896 3652 904
rect 3660 896 3668 904
rect 3740 896 3748 904
rect 1692 876 1700 884
rect 1868 876 1876 884
rect 2108 876 2116 884
rect 2284 876 2292 884
rect 2412 876 2420 884
rect 2556 876 2564 884
rect 2684 876 2692 884
rect 3436 876 3444 884
rect 3628 876 3636 884
rect 1388 856 1396 864
rect 1516 856 1524 864
rect 1532 856 1540 864
rect 1900 856 1908 864
rect 1164 836 1172 844
rect 1260 836 1268 844
rect 2476 836 2484 844
rect 1100 816 1108 824
rect 1756 816 1764 824
rect 2524 816 2532 824
rect 3356 816 3364 824
rect 3676 816 3684 824
rect 1436 796 1444 804
rect 1564 796 1572 804
rect 2348 796 2356 804
rect 3020 796 3028 804
rect 524 776 532 784
rect 796 776 804 784
rect 1052 776 1060 784
rect 1628 776 1636 784
rect 1660 776 1668 784
rect 2060 776 2068 784
rect 2156 776 2164 784
rect 3148 776 3156 784
rect 4108 776 4116 784
rect 1084 756 1092 764
rect 1228 756 1236 764
rect 1708 756 1716 764
rect 1916 756 1924 764
rect 2684 756 2692 764
rect 4188 756 4196 764
rect 1468 736 1476 744
rect 1724 736 1732 744
rect 1772 736 1780 744
rect 1932 736 1940 744
rect 2188 736 2196 744
rect 2412 736 2420 744
rect 2572 736 2580 744
rect 2604 736 2612 744
rect 3196 736 3204 744
rect 3260 736 3268 744
rect 3436 736 3444 744
rect 3500 736 3508 744
rect 300 716 308 724
rect 1068 716 1076 724
rect 1164 716 1172 724
rect 1596 716 1604 724
rect 1692 716 1700 724
rect 1948 716 1956 724
rect 2092 716 2100 724
rect 2124 716 2132 724
rect 2268 716 2276 724
rect 2332 716 2340 724
rect 2396 716 2404 724
rect 2412 716 2420 724
rect 2508 716 2516 724
rect 2924 716 2932 724
rect 2956 716 2964 724
rect 3068 716 3076 724
rect 3452 716 3460 724
rect 3884 716 3892 724
rect 3964 716 3972 724
rect 364 696 372 704
rect 460 696 468 704
rect 684 696 692 704
rect 732 696 740 704
rect 828 696 836 704
rect 1212 696 1220 704
rect 1228 696 1236 704
rect 2764 696 2772 704
rect 3388 696 3396 704
rect 3676 696 3684 704
rect 396 676 404 684
rect 1452 676 1460 684
rect 1948 676 1956 684
rect 2108 676 2116 684
rect 2204 676 2212 684
rect 2716 676 2724 684
rect 2908 676 2916 684
rect 3148 676 3156 684
rect 3580 676 3588 684
rect 3820 676 3828 684
rect 348 656 356 664
rect 2236 656 2244 664
rect 2252 656 2260 664
rect 2316 656 2324 664
rect 3244 656 3252 664
rect 3356 656 3364 664
rect 3532 656 3540 664
rect 444 636 452 644
rect 2300 636 2308 644
rect 2572 636 2580 644
rect 2700 636 2708 644
rect 2732 636 2740 644
rect 3116 636 3124 644
rect 3356 636 3364 644
rect 684 616 692 624
rect 1132 616 1140 624
rect 1404 616 1412 624
rect 1916 616 1924 624
rect 2284 616 2292 624
rect 2428 616 2436 624
rect 3100 616 3108 624
rect 3724 616 3732 624
rect 332 596 340 604
rect 1020 596 1028 604
rect 1340 596 1348 604
rect 1356 596 1364 604
rect 1404 596 1412 604
rect 1612 596 1620 604
rect 1964 596 1972 604
rect 2732 596 2740 604
rect 3308 596 3316 604
rect 3356 596 3364 604
rect 3580 596 3588 604
rect 4028 596 4036 604
rect 604 576 612 584
rect 1420 576 1428 584
rect 2140 576 2148 584
rect 3260 576 3268 584
rect 3324 576 3332 584
rect 3356 576 3364 584
rect 3468 576 3476 584
rect 412 556 420 564
rect 1004 556 1012 564
rect 1628 556 1636 564
rect 1884 556 1892 564
rect 1964 556 1972 564
rect 1980 556 1988 564
rect 2092 556 2100 564
rect 2156 556 2164 564
rect 2300 556 2308 564
rect 2444 556 2452 564
rect 2508 556 2516 564
rect 2764 556 2772 564
rect 2940 556 2948 564
rect 3244 556 3252 564
rect 3372 556 3380 564
rect 3436 556 3444 564
rect 3516 556 3524 564
rect 3564 556 3572 564
rect 284 536 292 544
rect 316 536 324 544
rect 380 536 388 544
rect 844 536 852 544
rect 924 536 932 544
rect 1116 536 1124 544
rect 1196 536 1204 544
rect 1308 536 1316 544
rect 1580 536 1588 544
rect 1804 536 1812 544
rect 1820 536 1828 544
rect 1852 536 1860 544
rect 188 516 196 524
rect 2540 536 2548 544
rect 3148 536 3156 544
rect 3596 536 3604 544
rect 3612 536 3620 544
rect 3676 536 3684 544
rect 3708 536 3716 544
rect 3740 536 3748 544
rect 3868 536 3876 544
rect 3884 536 3892 544
rect 3980 536 3988 544
rect 4076 536 4084 544
rect 300 496 308 504
rect 1036 496 1044 504
rect 2316 516 2324 524
rect 3404 516 3412 524
rect 3420 516 3428 524
rect 3532 516 3540 524
rect 3756 516 3764 524
rect 3772 516 3780 524
rect 2300 496 2308 504
rect 2556 496 2564 504
rect 2748 496 2756 504
rect 3964 496 3972 504
rect 1052 476 1060 484
rect 1228 476 1236 484
rect 2188 476 2196 484
rect 2556 476 2564 484
rect 3324 476 3332 484
rect 3340 476 3348 484
rect 3500 476 3508 484
rect 3948 476 3956 484
rect 3980 476 3988 484
rect 332 456 340 464
rect 1132 456 1140 464
rect 1548 456 1556 464
rect 2172 456 2180 464
rect 3740 456 3748 464
rect 3772 456 3780 464
rect 252 416 260 424
rect 1500 416 1508 424
rect 2348 416 2356 424
rect 3580 416 3588 424
rect 1212 396 1220 404
rect 1676 396 1684 404
rect 4140 396 4148 404
rect 1036 376 1044 384
rect 2140 376 2148 384
rect 2732 376 2740 384
rect 3404 376 3412 384
rect 3420 376 3428 384
rect 3484 376 3492 384
rect 156 356 164 364
rect 412 356 420 364
rect 2044 356 2052 364
rect 3068 356 3076 364
rect 3388 356 3396 364
rect 3516 356 3524 364
rect 3532 356 3540 364
rect 460 336 468 344
rect 796 336 804 344
rect 812 336 820 344
rect 1004 336 1012 344
rect 1148 336 1156 344
rect 1676 336 1684 344
rect 2556 336 2564 344
rect 2572 336 2580 344
rect 2956 336 2964 344
rect 3756 336 3764 344
rect 60 316 68 324
rect 636 316 644 324
rect 1228 316 1236 324
rect 1244 316 1252 324
rect 2028 316 2036 324
rect 2204 316 2212 324
rect 2220 316 2228 324
rect 2892 316 2900 324
rect 2940 316 2948 324
rect 3036 316 3044 324
rect 3180 316 3188 324
rect 3196 316 3204 324
rect 3260 316 3268 324
rect 3276 316 3284 324
rect 3596 316 3604 324
rect 3804 316 3812 324
rect 3948 316 3956 324
rect 1388 296 1396 304
rect 1500 296 1508 304
rect 1596 296 1604 304
rect 1628 296 1636 304
rect 2252 296 2260 304
rect 3548 296 3556 304
rect 4012 296 4020 304
rect 348 276 356 284
rect 2828 276 2836 284
rect 2876 276 2884 284
rect 2908 276 2916 284
rect 3244 276 3252 284
rect 3340 276 3348 284
rect 1260 256 1268 264
rect 860 236 868 244
rect 1612 236 1620 244
rect 1660 236 1668 244
rect 1980 256 1988 264
rect 2156 256 2164 264
rect 2412 256 2420 264
rect 2508 256 2516 264
rect 2524 256 2532 264
rect 2716 256 2724 264
rect 3148 256 3156 264
rect 3692 256 3700 264
rect 3948 256 3956 264
rect 4028 256 4036 264
rect 2044 236 2052 244
rect 2060 236 2068 244
rect 2940 236 2948 244
rect 3260 236 3268 244
rect 1004 216 1012 224
rect 1068 216 1076 224
rect 1180 216 1188 224
rect 1916 216 1924 224
rect 2428 216 2436 224
rect 2956 216 2964 224
rect 3004 216 3012 224
rect 3180 216 3188 224
rect 3740 216 3748 224
rect 3804 216 3812 224
rect 956 196 964 204
rect 1372 196 1380 204
rect 1548 196 1556 204
rect 1580 196 1588 204
rect 1900 196 1908 204
rect 2268 196 2276 204
rect 2684 196 2692 204
rect 2796 196 2804 204
rect 2860 196 2868 204
rect 4012 196 4020 204
rect 4044 196 4052 204
rect 604 176 612 184
rect 1468 176 1476 184
rect 1628 176 1636 184
rect 1820 176 1828 184
rect 1836 176 1844 184
rect 2044 176 2052 184
rect 2396 176 2404 184
rect 2588 176 2596 184
rect 2892 176 2900 184
rect 3276 176 3284 184
rect 3340 176 3348 184
rect 3836 176 3844 184
rect 4188 176 4196 184
rect 4220 176 4228 184
rect 332 156 340 164
rect 428 156 436 164
rect 556 156 564 164
rect 620 156 628 164
rect 2316 156 2324 164
rect 2972 156 2980 164
rect 364 136 372 144
rect 860 136 868 144
rect 892 136 900 144
rect 1132 136 1140 144
rect 1180 136 1188 144
rect 2108 136 2116 144
rect 2316 136 2324 144
rect 2604 136 2612 144
rect 2684 136 2692 144
rect 3756 156 3764 164
rect 3852 156 3860 164
rect 4092 156 4100 164
rect 4188 156 4196 164
rect 3836 136 3844 144
rect 4060 136 4068 144
rect 4076 136 4084 144
rect 4172 136 4180 144
rect 332 116 340 124
rect 812 96 820 104
rect 956 96 964 104
rect 1004 96 1012 104
rect 1100 96 1108 104
rect 1180 96 1188 104
rect 1196 96 1204 104
rect 2908 116 2916 124
rect 2956 116 2964 124
rect 3676 116 3684 124
rect 4092 116 4100 124
rect 2044 96 2052 104
rect 2332 96 2340 104
rect 2748 96 2756 104
rect 2860 96 2868 104
rect 3084 96 3092 104
rect 3100 96 3108 104
rect 3180 96 3188 104
rect 3548 96 3556 104
rect 3996 96 4004 104
rect 4156 96 4164 104
rect 4204 96 4212 104
rect 1164 76 1172 84
rect 1212 76 1220 84
rect 2876 16 2884 24
<< metal4 >>
rect 2525 2964 2531 2996
rect 2996 2977 3004 2983
rect 3613 2964 3619 2976
rect 1412 2957 1420 2963
rect 1716 2957 1724 2963
rect 2788 2957 2796 2963
rect 3540 2957 3548 2963
rect 4148 2957 4156 2963
rect 1373 2944 1379 2956
rect 2909 2944 2915 2956
rect 2973 2944 2979 2956
rect 2884 2937 2892 2943
rect 61 2504 67 2676
rect 125 2504 131 2736
rect 285 2624 291 2936
rect 525 2644 531 2756
rect 189 2284 195 2356
rect 109 2144 115 2156
rect 125 1584 131 1876
rect 141 1604 147 1896
rect 13 1444 19 1476
rect 93 1044 99 1296
rect 61 324 67 916
rect 125 904 131 976
rect 141 964 147 1016
rect 157 364 163 1076
rect 189 1064 195 2276
rect 221 2164 227 2336
rect 237 1944 243 1996
rect 205 1764 211 1856
rect 253 1764 259 2196
rect 269 2144 275 2356
rect 285 2164 291 2516
rect 349 2264 355 2316
rect 237 1484 243 1596
rect 253 1444 259 1456
rect 253 1064 259 1156
rect 269 1084 275 2136
rect 285 1124 291 1796
rect 173 944 179 956
rect 189 524 195 1056
rect 253 424 259 976
rect 301 724 307 1896
rect 340 1857 348 1863
rect 365 1784 371 2596
rect 477 2364 483 2636
rect 429 2324 435 2336
rect 477 2124 483 2316
rect 445 1784 451 1856
rect 413 1504 419 1536
rect 285 544 291 556
rect 301 504 307 716
rect 317 544 323 936
rect 333 904 339 1476
rect 365 1304 371 1336
rect 381 1324 387 1456
rect 397 1384 403 1456
rect 413 1384 419 1496
rect 429 1343 435 1416
rect 413 1337 435 1343
rect 388 1137 396 1143
rect 333 464 339 596
rect 349 284 355 656
rect 333 124 339 156
rect 365 144 371 696
rect 397 684 403 1076
rect 413 564 419 1337
rect 429 1064 435 1316
rect 429 964 435 1056
rect 445 644 451 1356
rect 461 1144 467 1756
rect 477 1324 483 2116
rect 493 1504 499 2196
rect 509 1663 515 2556
rect 532 2277 540 2283
rect 525 1924 531 2196
rect 509 1657 531 1663
rect 509 1344 515 1636
rect 509 984 515 1336
rect 509 964 515 976
rect 525 784 531 1657
rect 541 1264 547 2116
rect 541 1064 547 1096
rect 557 1084 563 2556
rect 589 2484 595 2696
rect 653 2464 659 2596
rect 669 2544 675 2896
rect 589 2124 595 2156
rect 589 2064 595 2096
rect 573 904 579 1056
rect 573 884 579 896
rect 589 704 595 996
rect 381 544 387 556
rect 413 344 419 356
rect 429 164 435 396
rect 461 344 467 696
rect 605 584 611 2276
rect 621 2164 627 2356
rect 637 2344 643 2396
rect 621 1484 627 2156
rect 621 1064 627 1476
rect 605 184 611 576
rect 621 164 627 956
rect 637 324 643 1956
rect 653 1744 659 2356
rect 669 1304 675 2336
rect 701 2124 707 2136
rect 685 1784 691 2076
rect 669 1124 675 1296
rect 669 1104 675 1116
rect 685 704 691 1756
rect 701 884 707 2116
rect 717 1944 723 2276
rect 733 1884 739 2916
rect 813 2624 819 2736
rect 749 2124 755 2156
rect 717 1084 723 1856
rect 749 1524 755 1976
rect 765 1684 771 2396
rect 829 2284 835 2676
rect 941 2644 947 2716
rect 964 2637 972 2643
rect 797 2164 803 2176
rect 781 1824 787 2116
rect 813 1904 819 2256
rect 829 2184 835 2236
rect 845 2163 851 2436
rect 829 2157 851 2163
rect 829 1924 835 2157
rect 804 1837 812 1843
rect 749 984 755 1516
rect 765 1124 771 1676
rect 781 1184 787 1616
rect 797 1304 803 1776
rect 813 1344 819 1636
rect 765 964 771 976
rect 749 924 755 936
rect 797 784 803 1036
rect 829 984 835 1896
rect 845 1484 851 2136
rect 861 904 867 2596
rect 909 2544 915 2616
rect 893 2504 899 2536
rect 989 2524 995 2636
rect 957 2204 963 2416
rect 973 1764 979 2336
rect 989 1864 995 2496
rect 893 1444 899 1476
rect 893 1404 899 1416
rect 909 1004 915 1656
rect 925 1384 931 1716
rect 925 1244 931 1296
rect 957 1044 963 1056
rect 916 977 924 983
rect 973 904 979 1276
rect 989 1224 995 1236
rect 989 984 995 1116
rect 989 964 995 976
rect 685 584 691 616
rect 813 344 819 876
rect 829 544 835 696
rect 845 544 851 556
rect 797 324 803 336
rect 861 244 867 896
rect 1005 564 1011 2696
rect 1021 2404 1027 2676
rect 1021 2304 1027 2316
rect 1021 2084 1027 2156
rect 1037 1664 1043 2796
rect 1053 2264 1059 2536
rect 1053 2124 1059 2256
rect 1069 2144 1075 2536
rect 1117 2364 1123 2616
rect 1245 2564 1251 2936
rect 1133 2344 1139 2496
rect 1069 1764 1075 1776
rect 1021 924 1027 1156
rect 1021 904 1027 916
rect 1021 604 1027 836
rect 1005 544 1011 556
rect 932 537 940 543
rect 1005 344 1011 536
rect 1037 504 1043 1056
rect 1053 964 1059 1756
rect 1085 1504 1091 2316
rect 1101 2044 1107 2236
rect 1133 2184 1139 2236
rect 1165 2144 1171 2216
rect 1165 1884 1171 1896
rect 1085 1364 1091 1376
rect 1085 1124 1091 1296
rect 1085 844 1091 1116
rect 1101 824 1107 1196
rect 1037 384 1043 496
rect 1053 484 1059 776
rect 1085 744 1091 756
rect 1117 544 1123 1076
rect 1133 904 1139 1096
rect 1133 464 1139 616
rect 1149 344 1155 1096
rect 1165 844 1171 1796
rect 1181 1784 1187 2316
rect 1229 2184 1235 2196
rect 1213 1784 1219 2176
rect 1245 1924 1251 2556
rect 1261 2544 1267 2576
rect 1277 2204 1283 2656
rect 1469 2584 1475 2656
rect 1485 2564 1491 2576
rect 1476 2557 1484 2563
rect 1460 2497 1468 2503
rect 1293 2144 1299 2236
rect 1309 2124 1315 2336
rect 1261 2064 1267 2076
rect 1229 1844 1235 1896
rect 1245 1884 1251 1916
rect 1341 1884 1347 2196
rect 1357 2164 1363 2496
rect 1165 724 1171 736
rect 1197 544 1203 1616
rect 1213 1064 1219 1736
rect 1229 1284 1235 1396
rect 1213 704 1219 1056
rect 1229 764 1235 1076
rect 1245 1024 1251 1036
rect 1261 844 1267 1876
rect 1277 1724 1283 1736
rect 1293 1704 1299 1856
rect 1309 1484 1315 1876
rect 1405 1864 1411 2256
rect 1421 2244 1427 2496
rect 1325 1744 1331 1796
rect 1341 1343 1347 1756
rect 1405 1684 1411 1856
rect 1357 1664 1363 1676
rect 1389 1564 1395 1596
rect 1373 1384 1379 1516
rect 1341 1337 1356 1343
rect 1293 1304 1299 1336
rect 1373 1304 1379 1316
rect 1293 1104 1299 1116
rect 1341 1064 1347 1276
rect 1373 1124 1379 1276
rect 1229 484 1235 696
rect 1213 304 1219 396
rect 1229 324 1235 336
rect 1261 264 1267 836
rect 1341 604 1347 1056
rect 1357 904 1363 956
rect 1373 924 1379 936
rect 1389 924 1395 1556
rect 1421 1524 1427 1536
rect 1389 864 1395 916
rect 1357 564 1363 596
rect 1309 404 1315 536
rect 548 157 556 163
rect 861 144 867 236
rect 1076 217 1084 223
rect 884 137 892 143
rect 813 104 819 136
rect 957 104 963 196
rect 1005 104 1011 216
rect 1181 144 1187 216
rect 1373 204 1379 476
rect 1389 304 1395 856
rect 1405 624 1411 1436
rect 1421 584 1427 1516
rect 1437 944 1443 2296
rect 1453 2284 1459 2496
rect 1501 2484 1507 2936
rect 1469 2184 1475 2256
rect 1501 2144 1507 2156
rect 1453 1844 1459 1856
rect 1485 1744 1491 2016
rect 1501 1744 1507 1836
rect 1437 764 1443 796
rect 1453 684 1459 1376
rect 1469 1284 1475 1496
rect 1485 1344 1491 1676
rect 1517 1584 1523 2876
rect 1533 2864 1539 2876
rect 1533 2364 1539 2656
rect 1533 2264 1539 2276
rect 1549 2264 1555 2556
rect 1565 2104 1571 2596
rect 1581 2424 1587 2556
rect 1661 2484 1667 2636
rect 1757 2504 1763 2516
rect 1613 2464 1619 2476
rect 1629 2324 1635 2356
rect 1677 2264 1683 2276
rect 1501 1364 1507 1376
rect 1517 1284 1523 1396
rect 1469 904 1475 1276
rect 1492 1057 1500 1063
rect 1485 964 1491 976
rect 1469 184 1475 736
rect 1501 424 1507 1016
rect 1533 864 1539 896
rect 1517 484 1523 856
rect 1549 464 1555 2076
rect 1581 2024 1587 2136
rect 1597 1844 1603 2036
rect 1693 2024 1699 2336
rect 1773 2264 1779 2276
rect 1709 2164 1715 2216
rect 1613 1844 1619 1856
rect 1629 1764 1635 1776
rect 1677 1764 1683 1796
rect 1581 1484 1587 1556
rect 1565 1024 1571 1476
rect 1661 1364 1667 1656
rect 1677 1464 1683 1476
rect 1581 1284 1587 1336
rect 1645 1024 1651 1076
rect 1565 724 1571 796
rect 1581 544 1587 936
rect 1661 784 1667 1356
rect 1693 1144 1699 1556
rect 1709 1524 1715 2056
rect 1725 1584 1731 2256
rect 1789 2164 1795 2696
rect 1805 2524 1811 2556
rect 1821 2524 1827 2616
rect 1837 2584 1843 2936
rect 2333 2924 2339 2936
rect 2525 2904 2531 2916
rect 2701 2904 2707 2936
rect 1917 2844 1923 2856
rect 2077 2684 2083 2876
rect 2116 2857 2124 2863
rect 2093 2724 2099 2736
rect 2148 2717 2156 2723
rect 1805 2164 1811 2516
rect 1837 2484 1843 2516
rect 1709 1164 1715 1476
rect 1725 1384 1731 1416
rect 1677 1084 1683 1096
rect 1677 924 1683 976
rect 1597 304 1603 716
rect 1492 297 1500 303
rect 1549 204 1555 296
rect 1613 244 1619 596
rect 1629 564 1635 776
rect 1661 744 1667 776
rect 1693 724 1699 876
rect 1709 764 1715 916
rect 1725 744 1731 1276
rect 1741 944 1747 2076
rect 1805 1944 1811 2156
rect 1821 2084 1827 2456
rect 1853 2204 1859 2636
rect 1869 2604 1875 2676
rect 1924 2657 1932 2663
rect 1901 2624 1907 2656
rect 1885 2584 1891 2596
rect 1901 2524 1907 2536
rect 1917 2504 1923 2656
rect 1997 2544 2003 2616
rect 2077 2584 2083 2676
rect 2109 2624 2115 2716
rect 2020 2537 2028 2543
rect 1917 2244 1923 2456
rect 1901 2164 1907 2176
rect 1917 2144 1923 2176
rect 1965 2144 1971 2176
rect 1773 1844 1779 1856
rect 1789 1704 1795 1916
rect 1757 1424 1763 1436
rect 1805 1124 1811 1936
rect 1821 1304 1827 1476
rect 1837 1324 1843 2096
rect 1981 2064 1987 2456
rect 2061 2384 2067 2576
rect 2109 2564 2115 2616
rect 2052 2337 2060 2343
rect 2013 2184 2019 2336
rect 1997 2064 2003 2076
rect 1853 1884 1859 1896
rect 1821 924 1827 936
rect 1837 904 1843 1076
rect 1853 904 1859 1876
rect 1869 1604 1875 1956
rect 1981 1924 1987 2056
rect 1981 1904 1987 1916
rect 1949 1884 1955 1896
rect 1885 1724 1891 1876
rect 1901 1864 1907 1876
rect 1917 1864 1923 1876
rect 1757 484 1763 816
rect 1773 744 1779 756
rect 1853 544 1859 896
rect 1869 884 1875 1596
rect 1885 1504 1891 1716
rect 1997 1684 2003 1876
rect 2013 1784 2019 2176
rect 2029 2064 2035 2076
rect 2029 2004 2035 2016
rect 2045 1964 2051 2336
rect 2077 2324 2083 2476
rect 1901 1344 1907 1396
rect 1885 964 1891 1336
rect 1917 1164 1923 1676
rect 1933 1464 1939 1676
rect 1949 1604 1955 1676
rect 1901 1084 1907 1096
rect 1901 864 1907 996
rect 1917 624 1923 756
rect 1933 704 1939 736
rect 1949 724 1955 1456
rect 1965 1064 1971 1636
rect 1997 1364 2003 1676
rect 2029 1564 2035 1576
rect 2061 1484 2067 2156
rect 2077 1564 2083 2236
rect 2093 2124 2099 2536
rect 2093 1884 2099 2016
rect 2109 1904 2115 2516
rect 2125 2284 2131 2296
rect 2125 2064 2131 2276
rect 2141 2264 2147 2276
rect 2148 2117 2156 2123
rect 2173 2103 2179 2476
rect 2189 2264 2195 2276
rect 2189 2124 2195 2256
rect 2157 2097 2179 2103
rect 2157 1964 2163 2097
rect 2109 1704 2115 1896
rect 2157 1844 2163 1876
rect 2125 1544 2131 1836
rect 2141 1804 2147 1836
rect 2157 1764 2163 1776
rect 2157 1704 2163 1716
rect 2141 1664 2147 1676
rect 2141 1584 2147 1656
rect 2020 1357 2028 1363
rect 1965 944 1971 1056
rect 1981 944 1987 956
rect 1972 917 1980 923
rect 1949 664 1955 676
rect 1965 604 1971 836
rect 1892 557 1900 563
rect 1965 544 1971 556
rect 1677 344 1683 396
rect 1629 304 1635 316
rect 1661 244 1667 256
rect 1581 204 1587 236
rect 1805 184 1811 536
rect 1821 524 1827 536
rect 1997 284 2003 1136
rect 2013 1104 2019 1316
rect 2061 1304 2067 1476
rect 2077 1284 2083 1396
rect 2125 1364 2131 1536
rect 2141 1344 2147 1376
rect 2013 924 2019 1096
rect 2029 704 2035 936
rect 2061 784 2067 1236
rect 2141 964 2147 1296
rect 2157 1104 2163 1696
rect 2173 1384 2179 1956
rect 2173 1284 2179 1296
rect 2189 1264 2195 2116
rect 2205 1764 2211 2296
rect 2237 2184 2243 2616
rect 2269 2544 2275 2636
rect 2317 2604 2323 2856
rect 2429 2584 2435 2656
rect 2445 2624 2451 2856
rect 2253 2284 2259 2496
rect 2269 2364 2275 2536
rect 2221 1844 2227 1856
rect 2205 1684 2211 1696
rect 2221 1604 2227 1776
rect 2237 1664 2243 1956
rect 2253 1724 2259 2276
rect 2269 1964 2275 2356
rect 2333 2344 2339 2396
rect 2349 2284 2355 2316
rect 2365 2284 2371 2296
rect 2429 2284 2435 2296
rect 2445 2284 2451 2376
rect 2461 2344 2467 2896
rect 2557 2857 2572 2863
rect 2557 2844 2563 2857
rect 2461 2304 2467 2336
rect 2301 2044 2307 2216
rect 2324 2117 2332 2123
rect 2276 1837 2284 1843
rect 2269 1784 2275 1816
rect 2301 1764 2307 1956
rect 2349 1944 2355 2276
rect 2365 2184 2371 2196
rect 2381 2124 2387 2156
rect 2205 1103 2211 1556
rect 2221 1264 2227 1276
rect 2189 1097 2211 1103
rect 2173 1044 2179 1076
rect 2189 964 2195 1097
rect 2125 944 2131 956
rect 2109 884 2115 896
rect 2100 717 2108 723
rect 2132 717 2140 723
rect 2084 557 2092 563
rect 2029 324 2035 496
rect 2045 364 2051 476
rect 1837 184 1843 276
rect 1981 244 1987 256
rect 2045 244 2051 356
rect 1901 204 1907 236
rect 1924 217 1932 223
rect 2045 184 2051 236
rect 1629 164 1635 176
rect 1181 104 1187 116
rect 1821 104 1827 176
rect 2061 123 2067 236
rect 2109 144 2115 676
rect 2141 384 2147 576
rect 2157 564 2163 776
rect 2189 704 2195 736
rect 2205 684 2211 1076
rect 2189 504 2195 536
rect 2173 464 2179 496
rect 2221 484 2227 1196
rect 2237 664 2243 1556
rect 2253 1504 2259 1716
rect 2301 1524 2307 1656
rect 2269 1344 2275 1516
rect 2317 1484 2323 1516
rect 2285 1364 2291 1456
rect 2301 1384 2307 1416
rect 2253 1144 2259 1276
rect 2269 1144 2275 1156
rect 2253 844 2259 1136
rect 2285 1124 2291 1136
rect 2269 924 2275 956
rect 2285 884 2291 1096
rect 2317 924 2323 1116
rect 2301 904 2307 916
rect 2253 664 2259 696
rect 2196 477 2204 483
rect 2205 324 2211 376
rect 2269 324 2275 716
rect 2285 624 2291 876
rect 2333 724 2339 1896
rect 2381 1784 2387 1796
rect 2349 1524 2355 1616
rect 2349 1384 2355 1436
rect 2365 983 2371 1616
rect 2397 1604 2403 2276
rect 2445 2144 2451 2196
rect 2413 1984 2419 1996
rect 2445 1964 2451 1996
rect 2461 1964 2467 2216
rect 2477 2124 2483 2516
rect 2493 2364 2499 2376
rect 2525 2264 2531 2656
rect 2541 2524 2547 2556
rect 2557 2504 2563 2616
rect 2605 2524 2611 2536
rect 2580 2517 2588 2523
rect 2541 2324 2547 2336
rect 2573 2324 2579 2476
rect 2621 2384 2627 2656
rect 2637 2444 2643 2796
rect 2653 2544 2659 2716
rect 2765 2664 2771 2716
rect 2413 1544 2419 1916
rect 2429 1604 2435 1916
rect 2397 1524 2403 1536
rect 2381 1344 2387 1416
rect 2397 1344 2403 1356
rect 2365 977 2387 983
rect 2381 964 2387 977
rect 2365 943 2371 956
rect 2349 937 2371 943
rect 2349 924 2355 937
rect 2324 657 2332 663
rect 2301 504 2307 556
rect 2221 304 2227 316
rect 2164 257 2172 263
rect 2269 204 2275 316
rect 2317 164 2323 516
rect 2349 424 2355 796
rect 2397 724 2403 1296
rect 2413 884 2419 1536
rect 2429 1524 2435 1576
rect 2429 1324 2435 1496
rect 2445 1364 2451 1736
rect 2477 1684 2483 2116
rect 2493 1744 2499 2256
rect 2541 2244 2547 2316
rect 2557 2244 2563 2276
rect 2516 2157 2524 2163
rect 2516 1957 2531 1963
rect 2509 1884 2515 1936
rect 2509 1804 2515 1836
rect 2509 1524 2515 1796
rect 2525 1604 2531 1916
rect 2477 1423 2483 1436
rect 2477 1417 2499 1423
rect 2429 924 2435 1316
rect 2445 1104 2451 1296
rect 2461 1084 2467 1396
rect 2477 1364 2483 1396
rect 2493 1364 2499 1417
rect 2413 744 2419 756
rect 2397 184 2403 716
rect 2429 624 2435 896
rect 2445 564 2451 916
rect 2477 844 2483 1196
rect 2509 1164 2515 1456
rect 2541 1364 2547 2236
rect 2557 2004 2563 2216
rect 2573 2144 2579 2316
rect 2557 1844 2563 1956
rect 2573 1744 2579 1756
rect 2589 1684 2595 1936
rect 2605 1724 2611 2096
rect 2557 1444 2563 1596
rect 2557 1364 2563 1436
rect 2573 1424 2579 1456
rect 2573 1364 2579 1376
rect 2541 1324 2547 1356
rect 2541 1144 2547 1296
rect 2493 944 2499 956
rect 2525 824 2531 1096
rect 2541 944 2547 1136
rect 2557 1084 2563 1336
rect 2589 1304 2595 1656
rect 2605 1504 2611 1536
rect 2605 1444 2611 1456
rect 2605 1304 2611 1376
rect 2621 1124 2627 2156
rect 2669 2144 2675 2236
rect 2573 1044 2579 1056
rect 2509 564 2515 716
rect 2509 264 2515 556
rect 2541 544 2547 936
rect 2557 904 2563 996
rect 2573 924 2579 996
rect 2557 504 2563 876
rect 2573 724 2579 736
rect 2573 644 2579 656
rect 2557 484 2563 496
rect 2548 337 2556 343
rect 2573 304 2579 336
rect 2420 257 2428 263
rect 2429 224 2435 236
rect 2589 184 2595 1056
rect 2605 744 2611 1076
rect 2621 1004 2627 1036
rect 2637 904 2643 1596
rect 2653 1424 2659 1436
rect 2669 1124 2675 1936
rect 2685 1584 2691 1596
rect 2701 1584 2707 2656
rect 2717 2524 2723 2596
rect 2749 2584 2755 2656
rect 2765 2544 2771 2656
rect 2788 2577 2796 2583
rect 2909 2544 2915 2576
rect 2925 2544 2931 2896
rect 2941 2684 2947 2916
rect 2941 2624 2947 2676
rect 2717 2464 2723 2476
rect 2765 2144 2771 2516
rect 2733 1484 2739 1996
rect 2749 1744 2755 1756
rect 2733 1464 2739 1476
rect 2685 1364 2691 1396
rect 2708 1357 2716 1363
rect 2733 1344 2739 1376
rect 2749 1364 2755 1556
rect 2685 764 2691 876
rect 2701 644 2707 1236
rect 2717 1004 2723 1096
rect 2733 964 2739 1196
rect 2717 264 2723 676
rect 2733 384 2739 596
rect 2749 504 2755 1356
rect 2765 704 2771 2136
rect 2781 1924 2787 2316
rect 2813 1924 2819 2256
rect 2836 1937 2844 1943
rect 2813 1864 2819 1916
rect 2861 1564 2867 2336
rect 2877 1924 2883 2376
rect 2893 2104 2899 2456
rect 2909 2364 2915 2516
rect 2909 2284 2915 2356
rect 2877 1784 2883 1916
rect 2877 1764 2883 1776
rect 2893 1764 2899 2096
rect 2909 1904 2915 2256
rect 2909 1744 2915 1896
rect 2925 1864 2931 2536
rect 2941 2344 2947 2456
rect 2957 2324 2963 2336
rect 2973 2324 2979 2616
rect 2996 2577 3004 2583
rect 2973 2104 2979 2136
rect 2989 2124 2995 2536
rect 3005 2464 3011 2496
rect 3005 2124 3011 2456
rect 3021 2184 3027 2576
rect 3037 2544 3043 2796
rect 3053 2604 3059 2616
rect 3069 2604 3075 2676
rect 3053 2544 3059 2576
rect 3053 2344 3059 2496
rect 3069 2304 3075 2536
rect 3069 2264 3075 2296
rect 2861 1524 2867 1556
rect 2909 1524 2915 1536
rect 2836 1397 2844 1403
rect 2813 1384 2819 1396
rect 2781 1364 2787 1376
rect 2845 1164 2851 1176
rect 2781 1124 2787 1156
rect 2861 1084 2867 1456
rect 2893 1444 2899 1456
rect 2877 1404 2883 1416
rect 2909 1364 2915 1376
rect 2829 1044 2835 1056
rect 2861 1044 2867 1056
rect 2845 964 2851 1036
rect 2765 564 2771 696
rect 2733 324 2739 376
rect 2829 284 2835 956
rect 2861 944 2867 956
rect 2877 944 2883 1336
rect 2893 1304 2899 1336
rect 2909 1304 2915 1316
rect 2893 324 2899 1276
rect 2909 684 2915 1156
rect 2925 964 2931 1856
rect 2941 1304 2947 2056
rect 3005 2044 3011 2116
rect 2957 1804 2963 1856
rect 2957 1484 2963 1496
rect 2925 724 2931 956
rect 2317 144 2323 156
rect 2605 144 2611 216
rect 2797 204 2803 236
rect 2685 144 2691 196
rect 2045 117 2067 123
rect 2045 104 2051 117
rect 2749 104 2755 136
rect 2861 104 2867 196
rect 1204 97 1212 103
rect 2340 97 2348 103
rect 2877 24 2883 276
rect 2893 184 2899 316
rect 2909 284 2915 676
rect 2941 564 2947 1256
rect 2957 1104 2963 1116
rect 2957 984 2963 996
rect 2973 984 2979 1916
rect 3012 1777 3020 1783
rect 3021 1704 3027 1716
rect 2989 1384 2995 1396
rect 2989 1264 2995 1316
rect 3005 1024 3011 1036
rect 2941 324 2947 336
rect 2941 244 2947 296
rect 2948 217 2956 223
rect 2973 164 2979 976
rect 3021 804 3027 1696
rect 3037 984 3043 1636
rect 3069 1544 3075 2256
rect 3085 2164 3091 2596
rect 3101 2584 3107 2596
rect 3149 2184 3155 2616
rect 3165 2604 3171 2956
rect 3213 2564 3219 2936
rect 3245 2924 3251 2956
rect 3268 2937 3276 2943
rect 3261 2644 3267 2656
rect 3181 2444 3187 2556
rect 3085 1684 3091 1796
rect 3069 1304 3075 1356
rect 3053 904 3059 996
rect 3037 324 3043 496
rect 3069 364 3075 716
rect 3085 344 3091 1676
rect 3101 1664 3107 1696
rect 3117 1564 3123 1736
rect 3133 1484 3139 2116
rect 3101 1464 3107 1476
rect 3101 624 3107 1416
rect 3149 784 3155 1516
rect 3165 1264 3171 1296
rect 3165 1004 3171 1256
rect 3181 1124 3187 1136
rect 3197 964 3203 2276
rect 3213 1784 3219 2256
rect 3213 1684 3219 1776
rect 3229 1744 3235 2236
rect 3213 1264 3219 1676
rect 3261 1664 3267 2636
rect 3293 2584 3299 2936
rect 3300 2237 3308 2243
rect 3277 1724 3283 1756
rect 3293 1644 3299 1696
rect 3325 1684 3331 2736
rect 3341 2544 3347 2556
rect 3357 2464 3363 2596
rect 3389 2124 3395 2596
rect 3421 2584 3427 2816
rect 3405 2544 3411 2576
rect 3453 2524 3459 2536
rect 3341 2004 3347 2016
rect 3341 1724 3347 1916
rect 3220 1057 3228 1063
rect 3245 984 3251 1476
rect 3261 1044 3267 1056
rect 3236 957 3244 963
rect 3277 744 3283 1456
rect 3309 1084 3315 1096
rect 3268 737 3276 743
rect 3149 684 3155 696
rect 3117 404 3123 636
rect 3149 264 3155 536
rect 3197 324 3203 736
rect 3245 564 3251 656
rect 3172 317 3180 323
rect 3245 284 3251 556
rect 3261 524 3267 576
rect 3277 324 3283 536
rect 3293 344 3299 976
rect 3309 584 3315 596
rect 3325 584 3331 1676
rect 3341 1524 3347 1656
rect 3341 1404 3347 1416
rect 3325 504 3331 576
rect 3341 484 3347 1296
rect 3357 1164 3363 2096
rect 3453 1944 3459 1956
rect 3373 1704 3379 1856
rect 3453 1804 3459 1816
rect 3389 1724 3395 1796
rect 3389 1704 3395 1716
rect 3373 1144 3379 1696
rect 3389 1284 3395 1656
rect 3357 664 3363 816
rect 3357 604 3363 616
rect 3373 564 3379 1056
rect 3389 1044 3395 1256
rect 3405 1164 3411 1736
rect 3405 1124 3411 1156
rect 3421 1124 3427 1536
rect 3437 1364 3443 1596
rect 3453 1464 3459 1496
rect 3469 1384 3475 2956
rect 3501 2584 3507 2596
rect 3485 1984 3491 2576
rect 3508 2537 3516 2543
rect 3389 724 3395 1036
rect 3261 244 3267 316
rect 3005 184 3011 216
rect 2909 124 2915 136
rect 2948 117 2956 123
rect 3101 104 3107 116
rect 3181 104 3187 216
rect 3277 184 3283 316
rect 3341 284 3347 476
rect 3389 364 3395 696
rect 3405 524 3411 1096
rect 3437 904 3443 1336
rect 3421 883 3427 896
rect 3421 877 3436 883
rect 3437 644 3443 736
rect 3453 724 3459 1356
rect 3469 964 3475 1356
rect 3485 1304 3491 1956
rect 3485 1284 3491 1296
rect 3485 964 3491 1256
rect 3501 1224 3507 2396
rect 3517 2304 3523 2536
rect 3533 2504 3539 2956
rect 3613 2724 3619 2956
rect 3549 2684 3555 2716
rect 3549 2243 3555 2596
rect 3565 2544 3571 2556
rect 3533 2237 3555 2243
rect 3517 2224 3523 2236
rect 3517 1764 3523 1976
rect 3533 1944 3539 2237
rect 3517 1664 3523 1676
rect 3469 944 3475 956
rect 3469 584 3475 936
rect 3428 557 3436 563
rect 3485 384 3491 936
rect 3501 744 3507 1156
rect 3517 944 3523 1616
rect 3533 1484 3539 1936
rect 3549 1404 3555 2136
rect 3533 1364 3539 1396
rect 3565 1104 3571 2176
rect 3581 2164 3587 2676
rect 3597 2504 3603 2676
rect 3597 2124 3603 2496
rect 3613 2384 3619 2716
rect 3629 2524 3635 2536
rect 3581 1644 3587 2056
rect 3581 1544 3587 1616
rect 3533 904 3539 936
rect 3517 884 3523 896
rect 3501 484 3507 736
rect 3405 364 3411 376
rect 3533 364 3539 396
rect 3389 324 3395 356
rect 3517 324 3523 356
rect 3549 304 3555 896
rect 3565 684 3571 956
rect 3581 684 3587 1136
rect 3565 564 3571 676
rect 3581 424 3587 596
rect 3597 544 3603 2116
rect 3613 1604 3619 2256
rect 3629 1624 3635 2496
rect 3645 2404 3651 2516
rect 3645 2344 3651 2356
rect 3613 1484 3619 1596
rect 3629 1584 3635 1596
rect 3613 964 3619 1376
rect 3629 1164 3635 1516
rect 3645 1224 3651 2296
rect 3661 2284 3667 2936
rect 3677 2924 3683 2936
rect 3885 2904 3891 2956
rect 3869 2724 3875 2896
rect 3981 2744 3987 2896
rect 3677 2364 3683 2696
rect 3821 2564 3827 2576
rect 3837 2504 3843 2576
rect 3869 2544 3875 2716
rect 3917 2584 3923 2596
rect 3901 2544 3907 2556
rect 3677 1964 3683 2356
rect 3693 2324 3699 2496
rect 3709 2144 3715 2296
rect 3709 1884 3715 2136
rect 3789 2084 3795 2496
rect 3821 2204 3827 2316
rect 3837 2224 3843 2296
rect 3821 2064 3827 2196
rect 3661 1384 3667 1776
rect 3613 924 3619 956
rect 3629 884 3635 1136
rect 3661 904 3667 936
rect 3677 824 3683 1676
rect 3693 1624 3699 1636
rect 3693 1424 3699 1556
rect 3709 1464 3715 1876
rect 3789 1664 3795 2016
rect 3789 1624 3795 1636
rect 3725 1324 3731 1476
rect 3700 1077 3708 1083
rect 3693 964 3699 1036
rect 3693 884 3699 956
rect 3677 544 3683 696
rect 3613 524 3619 536
rect 3677 484 3683 536
rect 3597 324 3603 336
rect 3341 184 3347 276
rect 3693 264 3699 876
rect 3725 624 3731 1316
rect 3741 904 3747 1576
rect 3716 537 3724 543
rect 3741 524 3747 536
rect 3757 524 3763 1116
rect 3789 1084 3795 1456
rect 3837 1344 3843 2136
rect 3853 1864 3859 2436
rect 3869 1944 3875 2536
rect 3885 2144 3891 2316
rect 3853 1164 3859 1756
rect 3853 1104 3859 1156
rect 3885 1104 3891 1916
rect 3901 1144 3907 2336
rect 3933 2264 3939 2356
rect 3917 2224 3923 2256
rect 3933 2224 3939 2236
rect 3949 2184 3955 2676
rect 3924 1477 3932 1483
rect 3949 1444 3955 1476
rect 3965 1344 3971 2556
rect 3981 2244 3987 2676
rect 4052 2537 4060 2543
rect 4077 2523 4083 2896
rect 4093 2764 4099 2776
rect 4061 2517 4083 2523
rect 4013 1984 4019 2196
rect 4013 1864 4019 1976
rect 4029 1704 4035 1776
rect 3789 944 3795 1076
rect 3805 944 3811 956
rect 3917 904 3923 936
rect 3965 724 3971 1336
rect 4013 1064 4019 1076
rect 4045 924 4051 1736
rect 4061 1204 4067 2517
rect 4077 2264 4083 2336
rect 4093 2184 4099 2736
rect 4093 1364 4099 1936
rect 4109 1924 4115 2796
rect 4157 2324 4163 2896
rect 4173 2524 4179 2536
rect 4125 2104 4131 2276
rect 4116 1857 4124 1863
rect 4125 1744 4131 1756
rect 4141 1744 4147 2176
rect 4157 1524 4163 1556
rect 3828 677 3836 683
rect 3741 464 3747 496
rect 3757 344 3763 516
rect 3773 504 3779 516
rect 3773 464 3779 476
rect 3741 204 3747 216
rect 3757 164 3763 336
rect 3805 304 3811 316
rect 3805 224 3811 256
rect 3837 184 3843 676
rect 3885 544 3891 716
rect 3949 484 3955 516
rect 3965 504 3971 716
rect 3981 484 3987 536
rect 3956 317 3964 323
rect 3853 164 3859 216
rect 4013 204 4019 296
rect 4029 264 4035 596
rect 4036 197 4044 203
rect 3677 124 3683 156
rect 3837 144 3843 156
rect 4061 144 4067 216
rect 4093 164 4099 1336
rect 4109 984 4115 1076
rect 4109 784 4115 956
rect 4077 144 4083 156
rect 4125 144 4131 1496
rect 4148 1317 4156 1323
rect 4148 1037 4156 1043
rect 4173 1023 4179 1596
rect 4189 1164 4195 2236
rect 4205 1304 4211 2796
rect 4205 1124 4211 1296
rect 4221 1244 4227 1476
rect 4157 1017 4179 1023
rect 4141 404 4147 1016
rect 3556 97 3564 103
rect 4004 97 4012 103
rect 4093 97 4099 116
rect 4157 104 4163 1017
rect 4173 144 4179 996
rect 4189 764 4195 996
rect 4205 204 4211 1076
rect 4221 164 4227 176
rect 4189 144 4195 156
rect 4212 97 4220 103
<< m5contact >>
rect 1692 2976 1700 2984
rect 3004 2976 3012 2984
rect 1404 2956 1412 2964
rect 1532 2956 1540 2964
rect 1708 2956 1716 2964
rect 2524 2956 2532 2964
rect 2780 2956 2788 2964
rect 2908 2956 2916 2964
rect 2972 2956 2980 2964
rect 3244 2956 3252 2964
rect 3532 2956 3540 2964
rect 3884 2956 3892 2964
rect 4140 2956 4148 2964
rect 1372 2936 1380 2944
rect 2332 2936 2340 2944
rect 2700 2936 2708 2944
rect 2892 2936 2900 2944
rect 3084 2936 3092 2944
rect 476 2636 484 2644
rect 284 2516 292 2524
rect 108 2136 116 2144
rect 140 1056 148 1064
rect 252 1436 260 1444
rect 172 936 180 944
rect 332 1856 340 1864
rect 428 2336 436 2344
rect 380 1836 388 1844
rect 444 1776 452 1784
rect 284 556 292 564
rect 396 1376 404 1384
rect 380 1316 388 1324
rect 364 1296 372 1304
rect 396 1136 404 1144
rect 428 1056 436 1064
rect 540 2276 548 2284
rect 492 1356 500 1364
rect 508 976 516 984
rect 492 956 500 964
rect 540 1096 548 1104
rect 588 2096 596 2104
rect 572 876 580 884
rect 588 696 596 704
rect 380 556 388 564
rect 428 396 436 404
rect 412 336 420 344
rect 668 2336 676 2344
rect 700 2136 708 2144
rect 652 1136 660 1144
rect 652 1096 660 1104
rect 668 1096 676 1104
rect 748 2156 756 2164
rect 956 2636 964 2644
rect 844 2556 852 2564
rect 844 2436 852 2444
rect 796 2156 804 2164
rect 828 2176 836 2184
rect 796 1836 804 1844
rect 780 1756 788 1764
rect 812 1076 820 1084
rect 780 1036 788 1044
rect 764 956 772 964
rect 748 936 756 944
rect 892 2536 900 2544
rect 988 2516 996 2524
rect 876 2116 884 2124
rect 892 1416 900 1424
rect 924 1236 932 1244
rect 956 1056 964 1064
rect 908 976 916 984
rect 988 1216 996 1224
rect 988 956 996 964
rect 812 876 820 884
rect 732 696 740 704
rect 684 576 692 584
rect 844 556 852 564
rect 828 536 836 544
rect 796 316 804 324
rect 1020 2356 1028 2364
rect 1020 2296 1028 2304
rect 1020 2256 1028 2264
rect 1020 2176 1028 2184
rect 1020 2156 1028 2164
rect 1132 2336 1140 2344
rect 1068 1776 1076 1784
rect 1020 916 1028 924
rect 1020 836 1028 844
rect 940 536 948 544
rect 1004 536 1012 544
rect 1164 2216 1172 2224
rect 1132 2176 1140 2184
rect 1164 1896 1172 1904
rect 1084 1356 1092 1364
rect 1084 836 1092 844
rect 1148 1096 1156 1104
rect 1084 736 1092 744
rect 1068 716 1076 724
rect 1228 2196 1236 2204
rect 1196 2116 1204 2124
rect 1196 1876 1204 1884
rect 1260 2536 1268 2544
rect 1468 2576 1476 2584
rect 1484 2556 1492 2564
rect 1452 2496 1460 2504
rect 1276 2196 1284 2204
rect 1292 2136 1300 2144
rect 1340 2216 1348 2224
rect 1324 2176 1332 2184
rect 1260 2056 1268 2064
rect 1228 1896 1236 1904
rect 1356 1876 1364 1884
rect 1228 1836 1236 1844
rect 1212 1776 1220 1784
rect 1196 1756 1204 1764
rect 1164 736 1172 744
rect 1228 1076 1236 1084
rect 1244 1036 1252 1044
rect 1244 896 1252 904
rect 1276 1736 1284 1744
rect 1420 2236 1428 2244
rect 1324 1376 1332 1384
rect 1292 1336 1300 1344
rect 1356 1656 1364 1664
rect 1388 1556 1396 1564
rect 1356 1416 1364 1424
rect 1372 1376 1380 1384
rect 1372 1296 1380 1304
rect 1372 1276 1380 1284
rect 1292 1096 1300 1104
rect 1292 916 1300 924
rect 1228 336 1236 344
rect 1244 316 1252 324
rect 1212 296 1220 304
rect 1372 936 1380 944
rect 1404 1496 1412 1504
rect 1356 896 1364 904
rect 1356 556 1364 564
rect 1372 476 1380 484
rect 1308 396 1316 404
rect 540 156 548 164
rect 1084 216 1092 224
rect 812 136 820 144
rect 876 136 884 144
rect 1404 596 1412 604
rect 1532 2876 1540 2884
rect 1564 2876 1572 2884
rect 1452 2276 1460 2284
rect 1468 2176 1476 2184
rect 1500 2156 1508 2164
rect 1484 2036 1492 2044
rect 1484 2016 1492 2024
rect 1452 1856 1460 1864
rect 1436 756 1444 764
rect 1756 2636 1764 2644
rect 1532 2276 1540 2284
rect 1756 2516 1764 2524
rect 1612 2476 1620 2484
rect 1628 2316 1636 2324
rect 1676 2276 1684 2284
rect 1676 2156 1684 2164
rect 1516 1396 1524 1404
rect 1500 1376 1508 1384
rect 1500 1056 1508 1064
rect 1484 976 1492 984
rect 1532 896 1540 904
rect 1516 476 1524 484
rect 1580 2016 1588 2024
rect 1772 2276 1780 2284
rect 1724 2256 1732 2264
rect 1708 2156 1716 2164
rect 1612 1856 1620 1864
rect 1692 1816 1700 1824
rect 1628 1776 1636 1784
rect 1612 1736 1620 1744
rect 1580 1476 1588 1484
rect 1676 1476 1684 1484
rect 1580 1356 1588 1364
rect 1580 1336 1588 1344
rect 1644 1076 1652 1084
rect 1596 1056 1604 1064
rect 1580 936 1588 944
rect 1564 716 1572 724
rect 1612 896 1620 904
rect 1740 2236 1748 2244
rect 1772 2176 1780 2184
rect 2412 2916 2420 2924
rect 2524 2916 2532 2924
rect 1916 2856 1924 2864
rect 2108 2856 2116 2864
rect 2092 2716 2100 2724
rect 2156 2716 2164 2724
rect 1868 2676 1876 2684
rect 2092 2676 2100 2684
rect 1820 2516 1828 2524
rect 1836 2476 1844 2484
rect 1724 1376 1732 1384
rect 1676 1096 1684 1104
rect 1676 916 1684 924
rect 1708 916 1716 924
rect 1484 296 1492 304
rect 1548 296 1556 304
rect 1660 736 1668 744
rect 1916 2656 1924 2664
rect 1884 2576 1892 2584
rect 1900 2536 1908 2544
rect 1932 2636 1940 2644
rect 2012 2536 2020 2544
rect 1916 2496 1924 2504
rect 1916 2236 1924 2244
rect 1852 2196 1860 2204
rect 1900 2156 1908 2164
rect 1916 2136 1924 2144
rect 1964 2136 1972 2144
rect 1772 1856 1780 1864
rect 1772 1696 1780 1704
rect 1756 1436 1764 1444
rect 1820 1876 1828 1884
rect 2108 2556 2116 2564
rect 2012 2336 2020 2344
rect 2044 2336 2052 2344
rect 1996 2256 2004 2264
rect 1996 2056 2004 2064
rect 1740 936 1748 944
rect 1820 916 1828 924
rect 1948 1896 1956 1904
rect 1980 1896 1988 1904
rect 1900 1856 1908 1864
rect 1916 1856 1924 1864
rect 1900 1736 1908 1744
rect 1884 1716 1892 1724
rect 1772 756 1780 764
rect 2028 2156 2036 2164
rect 2028 2076 2036 2084
rect 2028 1996 2036 2004
rect 2076 2316 2084 2324
rect 2044 1956 2052 1964
rect 1884 1496 1892 1504
rect 1900 1396 1908 1404
rect 1948 1596 1956 1604
rect 1932 1456 1940 1464
rect 1900 1096 1908 1104
rect 1900 996 1908 1004
rect 1884 956 1892 964
rect 2028 1576 2036 1584
rect 2092 2076 2100 2084
rect 2124 2296 2132 2304
rect 2140 2256 2148 2264
rect 2140 2116 2148 2124
rect 2204 2296 2212 2304
rect 2188 2256 2196 2264
rect 2124 2016 2132 2024
rect 2172 1956 2180 1964
rect 2092 1876 2100 1884
rect 2156 1876 2164 1884
rect 2140 1796 2148 1804
rect 2156 1776 2164 1784
rect 2156 1716 2164 1724
rect 2140 1676 2148 1684
rect 2140 1576 2148 1584
rect 2124 1536 2132 1544
rect 2012 1476 2020 1484
rect 2076 1476 2084 1484
rect 2028 1396 2036 1404
rect 2012 1356 2020 1364
rect 1980 956 1988 964
rect 1964 916 1972 924
rect 1964 836 1972 844
rect 1932 696 1940 704
rect 1948 656 1956 664
rect 1900 556 1908 564
rect 1980 556 1988 564
rect 1964 536 1972 544
rect 1756 476 1764 484
rect 1628 316 1636 324
rect 1660 256 1668 264
rect 1580 236 1588 244
rect 1820 516 1828 524
rect 2028 1296 2036 1304
rect 2140 1336 2148 1344
rect 2044 916 2052 924
rect 2172 1296 2180 1304
rect 2428 2576 2436 2584
rect 2268 2536 2276 2544
rect 2236 2176 2244 2184
rect 2220 1856 2228 1864
rect 2204 1676 2212 1684
rect 2332 2336 2340 2344
rect 2348 2316 2356 2324
rect 2364 2296 2372 2304
rect 2428 2296 2436 2304
rect 2556 2836 2564 2844
rect 2460 2296 2468 2304
rect 2396 2276 2404 2284
rect 2444 2276 2452 2284
rect 2332 2116 2340 2124
rect 2284 1836 2292 1844
rect 2268 1776 2276 1784
rect 2364 2176 2372 2184
rect 2380 2156 2388 2164
rect 2364 1956 2372 1964
rect 2348 1936 2356 1944
rect 2332 1896 2340 1904
rect 2220 1596 2228 1604
rect 2220 1436 2228 1444
rect 2220 1276 2228 1284
rect 2124 956 2132 964
rect 2108 896 2116 904
rect 2108 716 2116 724
rect 2140 716 2148 724
rect 2028 696 2036 704
rect 2076 556 2084 564
rect 2028 496 2036 504
rect 2044 476 2052 484
rect 1836 276 1844 284
rect 1996 276 2004 284
rect 1900 236 1908 244
rect 1980 236 1988 244
rect 1932 216 1940 224
rect 1804 176 1812 184
rect 1628 156 1636 164
rect 1132 136 1140 144
rect 1180 116 1188 124
rect 2188 696 2196 704
rect 2188 536 2196 544
rect 2172 496 2180 504
rect 2188 496 2196 504
rect 2300 1516 2308 1524
rect 2316 1476 2324 1484
rect 2284 1456 2292 1464
rect 2300 1376 2308 1384
rect 2316 1376 2324 1384
rect 2252 1276 2260 1284
rect 2268 1136 2276 1144
rect 2284 1116 2292 1124
rect 2316 1116 2324 1124
rect 2268 956 2276 964
rect 2300 916 2308 924
rect 2252 836 2260 844
rect 2252 696 2260 704
rect 2204 476 2212 484
rect 2220 476 2228 484
rect 2204 376 2212 384
rect 2380 1776 2388 1784
rect 2348 1436 2356 1444
rect 2444 2136 2452 2144
rect 2412 1976 2420 1984
rect 2492 2356 2500 2364
rect 2540 2556 2548 2564
rect 2604 2536 2612 2544
rect 2588 2516 2596 2524
rect 2540 2336 2548 2344
rect 2652 2536 2660 2544
rect 2636 2436 2644 2444
rect 2444 1956 2452 1964
rect 2460 1916 2468 1924
rect 2460 1816 2468 1824
rect 2396 1516 2404 1524
rect 2380 1416 2388 1424
rect 2380 1336 2388 1344
rect 2396 1336 2404 1344
rect 2380 956 2388 964
rect 2332 656 2340 664
rect 2300 636 2308 644
rect 2268 316 2276 324
rect 2220 296 2228 304
rect 2252 296 2260 304
rect 2172 256 2180 264
rect 2428 1516 2436 1524
rect 2556 2276 2564 2284
rect 2508 2156 2516 2164
rect 2508 1956 2516 1964
rect 2508 1836 2516 1844
rect 2508 1516 2516 1524
rect 2444 1296 2452 1304
rect 2476 1356 2484 1364
rect 2492 1356 2500 1364
rect 2428 896 2436 904
rect 2412 876 2420 884
rect 2412 756 2420 764
rect 2412 716 2420 724
rect 2556 2216 2564 2224
rect 2588 2076 2596 2084
rect 2588 1936 2596 1944
rect 2572 1756 2580 1764
rect 2588 1676 2596 1684
rect 2588 1656 2596 1664
rect 2572 1536 2580 1544
rect 2572 1456 2580 1464
rect 2572 1376 2580 1384
rect 2556 1356 2564 1364
rect 2540 1316 2548 1324
rect 2524 1096 2532 1104
rect 2492 936 2500 944
rect 2604 1536 2612 1544
rect 2604 1476 2612 1484
rect 2604 1436 2612 1444
rect 2604 1376 2612 1384
rect 2652 2076 2660 2084
rect 2636 1876 2644 1884
rect 2636 1596 2644 1604
rect 2572 1036 2580 1044
rect 2556 996 2564 1004
rect 2508 556 2516 564
rect 2572 916 2580 924
rect 2572 716 2580 724
rect 2572 656 2580 664
rect 2540 336 2548 344
rect 2572 296 2580 304
rect 2428 256 2436 264
rect 2524 256 2532 264
rect 2428 236 2436 244
rect 2620 1036 2628 1044
rect 2652 1436 2660 1444
rect 2748 2576 2756 2584
rect 2780 2576 2788 2584
rect 2940 2676 2948 2684
rect 2908 2536 2916 2544
rect 2716 2516 2724 2524
rect 2908 2516 2916 2524
rect 2716 2496 2724 2504
rect 2716 2476 2724 2484
rect 2684 1576 2692 1584
rect 2748 1736 2756 1744
rect 2748 1556 2756 1564
rect 2732 1456 2740 1464
rect 2684 1356 2692 1364
rect 2700 1356 2708 1364
rect 2732 1336 2740 1344
rect 2668 1116 2676 1124
rect 2684 1056 2692 1064
rect 2732 636 2740 644
rect 2796 2236 2804 2244
rect 2844 2196 2852 2204
rect 2844 1936 2852 1944
rect 2908 2276 2916 2284
rect 2876 1916 2884 1924
rect 2940 2456 2948 2464
rect 2988 2576 2996 2584
rect 2988 2536 2996 2544
rect 2956 2316 2964 2324
rect 2972 2316 2980 2324
rect 2972 2136 2980 2144
rect 3004 2496 3012 2504
rect 3052 2616 3060 2624
rect 3052 2576 3060 2584
rect 3052 2336 3060 2344
rect 3068 2296 3076 2304
rect 2956 2096 2964 2104
rect 2924 1856 2932 1864
rect 2908 1536 2916 1544
rect 2860 1456 2868 1464
rect 2844 1396 2852 1404
rect 2780 1376 2788 1384
rect 2812 1376 2820 1384
rect 2780 1156 2788 1164
rect 2844 1156 2852 1164
rect 2892 1436 2900 1444
rect 2892 1416 2900 1424
rect 2876 1396 2884 1404
rect 2908 1356 2916 1364
rect 2828 1056 2836 1064
rect 2860 1036 2868 1044
rect 2860 996 2868 1004
rect 2844 956 2852 964
rect 2860 956 2868 964
rect 2732 316 2740 324
rect 2908 1316 2916 1324
rect 3020 2036 3028 2044
rect 2956 1796 2964 1804
rect 2956 1476 2964 1484
rect 2956 1376 2964 1384
rect 2940 1296 2948 1304
rect 2924 956 2932 964
rect 2796 236 2804 244
rect 2604 216 2612 224
rect 2748 136 2756 144
rect 1100 96 1108 104
rect 1212 96 1220 104
rect 1820 96 1828 104
rect 2348 96 2356 104
rect 1164 76 1172 84
rect 1212 76 1220 84
rect 2956 1116 2964 1124
rect 2956 996 2964 1004
rect 3020 1776 3028 1784
rect 3020 1716 3028 1724
rect 2988 1396 2996 1404
rect 2988 1316 2996 1324
rect 3004 1016 3012 1024
rect 2956 716 2964 724
rect 2940 336 2948 344
rect 2956 336 2964 344
rect 2940 296 2948 304
rect 2940 216 2948 224
rect 2988 916 2996 924
rect 3036 1636 3044 1644
rect 3100 2576 3108 2584
rect 3100 2356 3108 2364
rect 3228 2936 3236 2944
rect 3180 2596 3188 2604
rect 3260 2936 3268 2944
rect 3260 2656 3268 2664
rect 3180 2556 3188 2564
rect 3100 2096 3108 2104
rect 3116 1736 3124 1744
rect 3052 1376 3060 1384
rect 3068 1296 3076 1304
rect 3052 996 3060 1004
rect 3036 976 3044 984
rect 3036 496 3044 504
rect 3100 1656 3108 1664
rect 3100 1476 3108 1484
rect 3164 1296 3172 1304
rect 3180 1136 3188 1144
rect 3212 2256 3220 2264
rect 3244 1716 3252 1724
rect 3292 2576 3300 2584
rect 3308 2456 3316 2464
rect 3292 2236 3300 2244
rect 3308 1856 3316 1864
rect 3276 1756 3284 1764
rect 3356 2596 3364 2604
rect 3340 2556 3348 2564
rect 3404 2576 3412 2584
rect 3420 2576 3428 2584
rect 3452 2516 3460 2524
rect 3340 1996 3348 2004
rect 3324 1676 3332 1684
rect 3340 1676 3348 1684
rect 3292 1636 3300 1644
rect 3228 1376 3236 1384
rect 3212 1056 3220 1064
rect 3260 1056 3268 1064
rect 3244 976 3252 984
rect 3244 956 3252 964
rect 3308 1076 3316 1084
rect 3308 976 3316 984
rect 3276 736 3284 744
rect 3148 696 3156 704
rect 3116 396 3124 404
rect 3084 336 3092 344
rect 3164 316 3172 324
rect 3276 536 3284 544
rect 3260 516 3268 524
rect 3340 1656 3348 1664
rect 3340 1416 3348 1424
rect 3340 1376 3348 1384
rect 3308 576 3316 584
rect 3324 496 3332 504
rect 3452 1936 3460 1944
rect 3452 1796 3460 1804
rect 3388 1696 3396 1704
rect 3388 1256 3396 1264
rect 3356 636 3364 644
rect 3356 616 3364 624
rect 3356 576 3364 584
rect 3404 1156 3412 1164
rect 3452 1456 3460 1464
rect 3516 2596 3524 2604
rect 3500 2576 3508 2584
rect 3516 2536 3524 2544
rect 3500 2496 3508 2504
rect 3484 1976 3492 1984
rect 3484 1956 3492 1964
rect 3436 1356 3444 1364
rect 3468 1356 3476 1364
rect 3388 716 3396 724
rect 3324 476 3332 484
rect 3292 336 3300 344
rect 3004 176 3012 184
rect 2908 136 2916 144
rect 2940 116 2948 124
rect 3100 116 3108 124
rect 3420 896 3428 904
rect 3484 1276 3492 1284
rect 3676 2936 3684 2944
rect 3548 2676 3556 2684
rect 3516 2296 3524 2304
rect 3516 2236 3524 2244
rect 3564 2556 3572 2564
rect 3516 1976 3524 1984
rect 3564 2236 3572 2244
rect 3516 1676 3524 1684
rect 3500 1156 3508 1164
rect 3468 936 3476 944
rect 3484 936 3492 944
rect 3436 636 3444 644
rect 3420 556 3428 564
rect 3420 516 3428 524
rect 3532 1356 3540 1364
rect 3580 2156 3588 2164
rect 3580 2136 3588 2144
rect 3628 2516 3636 2524
rect 3644 2516 3652 2524
rect 3580 2116 3588 2124
rect 3580 1536 3588 1544
rect 3580 1476 3588 1484
rect 3580 1416 3588 1424
rect 3532 996 3540 1004
rect 3516 936 3524 944
rect 3532 936 3540 944
rect 3516 876 3524 884
rect 3532 656 3540 664
rect 3516 556 3524 564
rect 3532 516 3540 524
rect 3532 396 3540 404
rect 3420 376 3428 384
rect 3404 356 3412 364
rect 3388 316 3396 324
rect 3516 316 3524 324
rect 3564 676 3572 684
rect 3644 2336 3652 2344
rect 3644 2296 3652 2304
rect 3628 1596 3636 1604
rect 3628 1556 3636 1564
rect 3628 1516 3636 1524
rect 3836 2576 3844 2584
rect 3820 2556 3828 2564
rect 3756 2536 3764 2544
rect 3948 2676 3956 2684
rect 3916 2576 3924 2584
rect 3900 2556 3908 2564
rect 3676 1956 3684 1964
rect 3820 2316 3828 2324
rect 3836 2296 3844 2304
rect 3724 1936 3732 1944
rect 3660 1376 3668 1384
rect 3612 896 3620 904
rect 3660 956 3668 964
rect 3660 936 3668 944
rect 3644 896 3652 904
rect 3692 1616 3700 1624
rect 3788 1636 3796 1644
rect 3724 1536 3732 1544
rect 3692 1376 3700 1384
rect 3708 1076 3716 1084
rect 3692 876 3700 884
rect 3612 516 3620 524
rect 3676 476 3684 484
rect 3596 336 3604 344
rect 3772 1356 3780 1364
rect 3772 1296 3780 1304
rect 3724 536 3732 544
rect 3868 1756 3876 1764
rect 3916 2256 3924 2264
rect 3932 2236 3940 2244
rect 3916 2136 3924 2144
rect 3916 1476 3924 1484
rect 3948 1436 3956 1444
rect 4060 2536 4068 2544
rect 4092 2756 4100 2764
rect 3852 1096 3860 1104
rect 3836 1076 3844 1084
rect 3804 956 3812 964
rect 3916 896 3924 904
rect 4012 1056 4020 1064
rect 4076 2336 4084 2344
rect 4140 2496 4148 2504
rect 4172 2516 4180 2524
rect 4124 1856 4132 1864
rect 4124 1736 4132 1744
rect 4172 1616 4180 1624
rect 4156 1556 4164 1564
rect 3836 676 3844 684
rect 3740 516 3748 524
rect 3740 496 3748 504
rect 3772 496 3780 504
rect 3772 476 3780 484
rect 3740 196 3748 204
rect 3804 296 3812 304
rect 3804 256 3812 264
rect 3868 536 3876 544
rect 3948 516 3956 524
rect 3964 316 3972 324
rect 3948 256 3956 264
rect 3852 216 3860 224
rect 4076 536 4084 544
rect 4060 216 4068 224
rect 4028 196 4036 204
rect 3676 156 3684 164
rect 3836 156 3844 164
rect 4108 976 4116 984
rect 4076 156 4084 164
rect 4156 1356 4164 1364
rect 4156 1316 4164 1324
rect 4156 1036 4164 1044
rect 4124 136 4132 144
rect 4092 116 4100 124
rect 3084 96 3092 104
rect 3564 96 3572 104
rect 4012 96 4020 104
rect 4204 196 4212 204
rect 4188 176 4196 184
rect 4220 156 4228 164
rect 4188 136 4196 144
rect 4220 96 4228 104
<< metal5 >>
rect 1700 2977 3004 2983
rect 1412 2957 1532 2963
rect 1716 2957 2524 2963
rect 2788 2957 2908 2963
rect 2980 2957 3244 2963
rect 3540 2957 3884 2963
rect 4148 2957 4155 2963
rect 1380 2937 2332 2943
rect 2708 2937 2892 2943
rect 3092 2937 3228 2943
rect 3268 2937 3676 2943
rect 2420 2917 2524 2923
rect 1540 2877 1564 2883
rect 1924 2857 2108 2863
rect 2557 2844 2563 2855
rect 2100 2717 2156 2723
rect 1876 2677 2092 2683
rect 2948 2677 3548 2683
rect 3556 2677 3948 2683
rect 1924 2657 3260 2663
rect 484 2637 956 2643
rect 1764 2637 1932 2643
rect 3060 2617 3067 2623
rect 2605 2597 3180 2603
rect 1476 2577 1884 2583
rect 2605 2583 2611 2597
rect 3364 2597 3516 2603
rect 2436 2577 2611 2583
rect 2756 2577 2780 2583
rect 2996 2577 3052 2583
rect 3077 2577 3100 2583
rect 3300 2577 3404 2583
rect 3428 2577 3500 2583
rect 3844 2577 3916 2583
rect 852 2557 1484 2563
rect 2116 2557 2540 2563
rect 3188 2557 3340 2563
rect 3397 2557 3564 2563
rect 3828 2557 3900 2563
rect 900 2537 1260 2543
rect 1908 2537 2012 2543
rect 2276 2537 2604 2543
rect 2660 2537 2715 2543
rect 2996 2537 3516 2543
rect 3764 2537 4060 2543
rect 292 2517 988 2523
rect 1764 2517 1820 2523
rect 2596 2517 2716 2523
rect 2916 2517 3452 2523
rect 3460 2517 3628 2523
rect 3652 2517 4172 2523
rect 1460 2497 1916 2503
rect 2724 2497 3004 2503
rect 3508 2497 4140 2503
rect 1620 2477 1836 2483
rect 2948 2457 3308 2463
rect 852 2437 2636 2443
rect 1028 2357 2492 2363
rect 3077 2357 3100 2363
rect 436 2337 668 2343
rect 676 2337 1132 2343
rect 1140 2337 2012 2343
rect 2052 2337 2332 2343
rect 2548 2337 3052 2343
rect 3652 2337 4076 2343
rect 2084 2317 2348 2323
rect 2373 2317 2956 2323
rect 2980 2317 3820 2323
rect 1028 2297 2115 2303
rect 548 2277 1452 2283
rect 1540 2277 1676 2283
rect 1701 2277 1772 2283
rect 2109 2283 2115 2297
rect 2132 2297 2204 2303
rect 2212 2297 2364 2303
rect 2381 2297 2428 2303
rect 2381 2283 2387 2297
rect 2468 2297 3068 2303
rect 3524 2297 3644 2303
rect 3652 2297 3836 2303
rect 2109 2277 2387 2283
rect 2404 2277 2444 2283
rect 2452 2277 2556 2283
rect 1028 2257 1724 2263
rect 2004 2257 2140 2263
rect 2196 2257 3212 2263
rect 3220 2257 3916 2263
rect 1428 2237 1740 2243
rect 1924 2237 2796 2243
rect 3300 2237 3516 2243
rect 3572 2237 3932 2243
rect 1172 2217 1340 2223
rect 1236 2197 1276 2203
rect 1860 2197 2844 2203
rect 836 2177 1020 2183
rect 1140 2177 1324 2183
rect 1476 2177 1772 2183
rect 2244 2177 2364 2183
rect 756 2157 796 2163
rect 1028 2157 1315 2163
rect 116 2137 595 2143
rect 589 2104 595 2137
rect 708 2137 1292 2143
rect 1309 2143 1315 2157
rect 1508 2157 1676 2163
rect 1716 2157 1900 2163
rect 2036 2157 2107 2163
rect 2388 2157 2508 2163
rect 1309 2137 1916 2143
rect 1972 2137 2444 2143
rect 2885 2137 2972 2143
rect 3588 2137 3916 2143
rect 884 2117 1196 2123
rect 2148 2117 2332 2123
rect 3588 2117 3611 2123
rect 2964 2097 3100 2103
rect 2036 2077 2092 2083
rect 2596 2077 2652 2083
rect 1268 2057 1996 2063
rect 1492 2037 3020 2043
rect 1492 2017 1580 2023
rect 1588 2017 2124 2023
rect 2036 1997 3340 2003
rect 2405 1977 2412 1983
rect 3492 1977 3516 1983
rect 2052 1957 2172 1963
rect 2372 1957 2444 1963
rect 2516 1957 2523 1963
rect 3492 1957 3676 1963
rect 2356 1937 2588 1943
rect 2852 1937 2875 1943
rect 3460 1937 3724 1943
rect 2468 1917 2876 1923
rect 1172 1897 1228 1903
rect 1253 1897 1948 1903
rect 1988 1897 2332 1903
rect 2340 1897 2363 1903
rect 1204 1877 1356 1883
rect 1828 1877 2092 1883
rect 2164 1877 2636 1883
rect 340 1857 1243 1863
rect 1460 1857 1612 1863
rect 1780 1857 1900 1863
rect 1924 1857 2220 1863
rect 2228 1857 2924 1863
rect 3316 1857 4124 1863
rect 388 1837 796 1843
rect 1236 1837 2284 1843
rect 2516 1837 2523 1843
rect 1700 1817 2460 1823
rect 2964 1797 3452 1803
rect 452 1777 1068 1783
rect 1220 1777 1628 1783
rect 2164 1777 2268 1783
rect 2388 1777 3020 1783
rect 788 1757 1196 1763
rect 2117 1757 2572 1763
rect 3284 1757 3868 1763
rect 1284 1737 1612 1743
rect 1908 1737 2748 1743
rect 3124 1737 4124 1743
rect 1892 1717 2156 1723
rect 3028 1717 3244 1723
rect 1780 1697 3388 1703
rect 2148 1677 2204 1683
rect 2596 1677 3324 1683
rect 3348 1677 3516 1683
rect 1364 1657 2588 1663
rect 3108 1657 3340 1663
rect 2917 1637 3036 1643
rect 3300 1637 3788 1643
rect 3700 1617 3707 1623
rect 4180 1617 4187 1623
rect 1956 1597 2163 1603
rect 2036 1577 2140 1583
rect 2157 1583 2163 1597
rect 2228 1597 2636 1603
rect 3621 1597 3628 1603
rect 2157 1577 2684 1583
rect 1396 1557 2748 1563
rect 3636 1557 4156 1563
rect 2132 1537 2572 1543
rect 2612 1537 2908 1543
rect 3588 1537 3611 1543
rect 3717 1537 3724 1543
rect 2308 1517 2396 1523
rect 2516 1517 3628 1523
rect 1412 1497 1884 1503
rect 1588 1477 1676 1483
rect 2020 1477 2076 1483
rect 2324 1477 2604 1483
rect 2629 1477 2883 1483
rect 1940 1457 2284 1463
rect 2309 1457 2555 1463
rect 2580 1457 2723 1463
rect 260 1437 899 1443
rect 893 1424 899 1437
rect 1764 1437 2220 1443
rect 2356 1437 2604 1443
rect 2629 1437 2652 1443
rect 2717 1443 2723 1457
rect 2740 1457 2860 1463
rect 2877 1463 2883 1477
rect 2964 1477 3100 1483
rect 3588 1477 3916 1483
rect 2877 1457 3452 1463
rect 2717 1437 2892 1443
rect 3365 1437 3948 1443
rect 1364 1417 2299 1423
rect 2388 1417 2892 1423
rect 3348 1417 3580 1423
rect 1524 1397 1900 1403
rect 2036 1397 2844 1403
rect 2884 1397 2988 1403
rect 404 1377 1324 1383
rect 1380 1377 1500 1383
rect 1732 1377 2300 1383
rect 2324 1377 2572 1383
rect 2612 1377 2780 1383
rect 2820 1377 2956 1383
rect 3060 1377 3228 1383
rect 3348 1377 3355 1383
rect 3668 1377 3692 1383
rect 500 1357 1084 1363
rect 1588 1357 2012 1363
rect 2149 1357 2476 1363
rect 2500 1357 2523 1363
rect 2597 1357 2684 1363
rect 2708 1357 2908 1363
rect 3444 1357 3468 1363
rect 3540 1357 3772 1363
rect 4101 1357 4156 1363
rect 1300 1337 1580 1343
rect 2148 1337 2380 1343
rect 2404 1337 2732 1343
rect 388 1317 2491 1323
rect 2548 1317 2908 1323
rect 2996 1317 4156 1323
rect 372 1297 1372 1303
rect 2036 1297 2172 1303
rect 2452 1297 2940 1303
rect 3076 1297 3164 1303
rect 3405 1297 3772 1303
rect 1380 1277 2220 1283
rect 3405 1283 3411 1297
rect 2260 1277 3411 1283
rect 3429 1277 3484 1283
rect 932 1237 995 1243
rect 989 1224 995 1237
rect 2788 1157 2844 1163
rect 3412 1157 3500 1163
rect 404 1137 652 1143
rect 2276 1137 3180 1143
rect 2292 1117 2316 1123
rect 2676 1117 2956 1123
rect 548 1097 652 1103
rect 676 1097 1148 1103
rect 1300 1097 1676 1103
rect 1908 1097 2524 1103
rect 2532 1097 3852 1103
rect 820 1077 1228 1083
rect 1652 1077 3308 1083
rect 3716 1077 3836 1083
rect 148 1057 428 1063
rect 964 1057 1500 1063
rect 1604 1057 2684 1063
rect 2709 1057 2747 1063
rect 2836 1057 3212 1063
rect 3268 1057 4012 1063
rect 788 1037 1244 1043
rect 2580 1037 2587 1043
rect 2628 1037 2787 1043
rect 2781 1023 2787 1037
rect 2868 1037 4156 1043
rect 2781 1017 3004 1023
rect 1908 997 2556 1003
rect 2757 997 2860 1003
rect 2949 997 2956 1003
rect 3060 997 3532 1003
rect 516 977 908 983
rect 916 977 1484 983
rect 1492 977 3036 983
rect 3252 977 3308 983
rect 4101 977 4108 983
rect 500 957 764 963
rect 996 957 1884 963
rect 1892 957 1980 963
rect 2132 957 2268 963
rect 2388 957 2844 963
rect 2868 957 2907 963
rect 2932 957 3244 963
rect 3668 957 3804 963
rect 180 937 748 943
rect 1380 937 1580 943
rect 1588 937 1740 943
rect 1748 937 2492 943
rect 2500 937 3468 943
rect 3492 937 3516 943
rect 3540 937 3660 943
rect 1028 917 1292 923
rect 1300 917 1676 923
rect 1716 917 1820 923
rect 1972 917 2044 923
rect 2308 917 2555 923
rect 2580 917 2988 923
rect 3397 917 3579 923
rect 1252 897 1356 903
rect 1364 897 1532 903
rect 1620 897 2108 903
rect 3421 885 3427 896
rect 3589 897 3612 903
rect 3652 897 3916 903
rect 580 877 812 883
rect 820 877 2412 883
rect 3524 877 3692 883
rect 1028 837 1084 843
rect 1092 837 1964 843
rect 1972 837 2252 843
rect 1444 757 1772 763
rect 2405 757 2412 763
rect 1092 737 1164 743
rect 1668 737 3276 743
rect 1076 717 1564 723
rect 1572 717 2108 723
rect 2148 717 2412 723
rect 2580 717 2956 723
rect 596 697 732 703
rect 1940 697 2028 703
rect 2196 697 2252 703
rect 3389 703 3395 716
rect 3156 697 3395 703
rect 3572 677 3836 683
rect 1956 657 2332 663
rect 2580 657 3532 663
rect 2308 637 2732 643
rect 3364 637 3436 643
rect 3357 605 3363 616
rect 861 597 1404 603
rect 861 583 867 597
rect 692 577 867 583
rect 3316 577 3356 583
rect 292 557 380 563
rect 852 557 1356 563
rect 1908 557 1980 563
rect 2084 557 2508 563
rect 3365 557 3420 563
rect 3524 557 3771 563
rect 836 537 940 543
rect 1012 537 1964 543
rect 1972 537 2188 543
rect 3284 537 3724 543
rect 3876 537 4076 543
rect 1828 517 2107 523
rect 3268 517 3420 523
rect 3540 517 3612 523
rect 3748 517 3948 523
rect 2036 497 2172 503
rect 2196 497 3036 503
rect 3044 497 3324 503
rect 3748 497 3772 503
rect 1380 477 1516 483
rect 1524 477 1756 483
rect 2052 477 2204 483
rect 2212 477 2220 483
rect 3332 477 3676 483
rect 436 397 1308 403
rect 3124 397 3532 403
rect 2212 377 3420 383
rect 3397 357 3404 363
rect 420 337 1211 343
rect 1236 337 2540 343
rect 2548 337 2555 343
rect 2565 337 2940 343
rect 2964 337 3084 343
rect 3300 337 3596 343
rect 804 317 1244 323
rect 1285 317 1628 323
rect 2276 317 2732 323
rect 3172 317 3388 323
rect 3524 317 3964 323
rect 1220 297 1484 303
rect 1556 297 2220 303
rect 2260 297 2572 303
rect 2948 297 3804 303
rect 1844 277 1996 283
rect 1668 257 2172 263
rect 2436 257 2524 263
rect 3812 257 3948 263
rect 1588 237 1883 243
rect 1908 237 1980 243
rect 2436 237 2796 243
rect 1092 217 1932 223
rect 2612 217 2940 223
rect 3860 217 4060 223
rect 1893 197 3740 203
rect 4036 197 4204 203
rect 1812 177 3004 183
rect 4165 177 4188 183
rect 548 157 1628 163
rect 3684 157 3836 163
rect 4084 157 4220 163
rect 820 137 876 143
rect 1140 137 1187 143
rect 1181 124 1187 137
rect 2756 137 2908 143
rect 4132 137 4188 143
rect 2948 117 3100 123
rect 4093 105 4099 116
rect 1108 97 1212 103
rect 1828 97 2348 103
rect 3092 97 3564 103
rect 3621 97 4012 103
rect 4197 97 4220 103
rect 1172 77 1212 83
<< m6contact >>
rect 4155 2955 4165 2965
rect 2555 2855 2565 2865
rect 4091 2764 4101 2765
rect 4091 2756 4092 2764
rect 4092 2756 4100 2764
rect 4100 2756 4101 2764
rect 4091 2755 4101 2756
rect 3067 2615 3077 2625
rect 3067 2575 3077 2585
rect 3387 2555 3397 2565
rect 2715 2535 2725 2545
rect 2907 2544 2917 2545
rect 2907 2536 2908 2544
rect 2908 2536 2916 2544
rect 2916 2536 2917 2544
rect 2907 2535 2917 2536
rect 2715 2484 2725 2485
rect 2715 2476 2716 2484
rect 2716 2476 2724 2484
rect 2724 2476 2725 2484
rect 2715 2475 2725 2476
rect 3067 2355 3077 2365
rect 1627 2324 1637 2325
rect 1627 2316 1628 2324
rect 1628 2316 1636 2324
rect 1636 2316 1637 2324
rect 1627 2315 1637 2316
rect 2363 2315 2373 2325
rect 1691 2275 1701 2285
rect 2907 2284 2917 2285
rect 2907 2276 2908 2284
rect 2908 2276 2916 2284
rect 2916 2276 2917 2284
rect 2907 2275 2917 2276
rect 2555 2224 2565 2225
rect 2555 2216 2556 2224
rect 2556 2216 2564 2224
rect 2564 2216 2565 2224
rect 2555 2215 2565 2216
rect 2107 2155 2117 2165
rect 3579 2164 3589 2165
rect 3579 2156 3580 2164
rect 3580 2156 3588 2164
rect 3588 2156 3589 2164
rect 3579 2155 3589 2156
rect 2875 2135 2885 2145
rect 3611 2115 3621 2125
rect 2395 1975 2405 1985
rect 2523 1955 2533 1965
rect 2875 1935 2885 1945
rect 1243 1895 1253 1905
rect 2363 1895 2373 1905
rect 1243 1855 1253 1865
rect 2523 1835 2533 1845
rect 2139 1804 2149 1805
rect 2139 1796 2140 1804
rect 2140 1796 2148 1804
rect 2148 1796 2149 1804
rect 2139 1795 2149 1796
rect 2107 1755 2117 1765
rect 2907 1635 2917 1645
rect 3707 1615 3717 1625
rect 4187 1615 4197 1625
rect 3611 1595 3621 1605
rect 3611 1535 3621 1545
rect 3707 1535 3717 1545
rect 2427 1524 2437 1525
rect 2427 1516 2428 1524
rect 2428 1516 2436 1524
rect 2436 1516 2437 1524
rect 2427 1515 2437 1516
rect 2619 1475 2629 1485
rect 2299 1455 2309 1465
rect 2555 1455 2565 1465
rect 2619 1435 2629 1445
rect 3355 1435 3365 1445
rect 2299 1415 2309 1425
rect 3355 1375 3365 1385
rect 2139 1355 2149 1365
rect 2523 1355 2533 1365
rect 2555 1364 2565 1365
rect 2555 1356 2556 1364
rect 2556 1356 2564 1364
rect 2564 1356 2565 1364
rect 2555 1355 2565 1356
rect 2587 1355 2597 1365
rect 4091 1355 4101 1365
rect 2491 1315 2501 1325
rect 3419 1275 3429 1285
rect 3387 1264 3397 1265
rect 3387 1256 3388 1264
rect 3388 1256 3396 1264
rect 3396 1256 3397 1264
rect 3387 1255 3397 1256
rect 2699 1055 2709 1065
rect 2747 1055 2757 1065
rect 2587 1035 2597 1045
rect 2747 995 2757 1005
rect 2939 995 2949 1005
rect 4091 975 4101 985
rect 2907 955 2917 965
rect 2555 915 2565 925
rect 3387 915 3397 925
rect 3579 915 3589 925
rect 2427 904 2437 905
rect 2427 896 2428 904
rect 2428 896 2436 904
rect 2436 896 2437 904
rect 2427 895 2437 896
rect 3579 895 3589 905
rect 3419 875 3429 885
rect 2395 755 2405 765
rect 3355 595 3365 605
rect 3355 555 3365 565
rect 3771 555 3781 565
rect 2107 515 2117 525
rect 3771 484 3781 485
rect 3771 476 3772 484
rect 3772 476 3780 484
rect 3780 476 3781 484
rect 3771 475 3781 476
rect 3387 355 3397 365
rect 1211 335 1221 345
rect 2555 335 2565 345
rect 1275 315 1285 325
rect 1883 235 1893 245
rect 1883 195 1893 205
rect 4155 175 4165 185
rect 3611 95 3621 105
rect 4091 95 4101 105
rect 4187 95 4197 105
<< metal6 >>
rect 1627 2305 1637 2315
rect 1627 2295 1701 2305
rect 1691 2285 1701 2295
rect 1243 1865 1253 1895
rect 2107 1765 2117 2155
rect 2363 1905 2373 2315
rect 2555 2225 2565 2855
rect 3067 2585 3077 2615
rect 2715 2485 2725 2535
rect 2907 2345 2917 2535
rect 3067 2345 3077 2355
rect 2907 2335 3077 2345
rect 2107 525 2117 1755
rect 2139 1365 2149 1795
rect 2299 1425 2309 1455
rect 2395 765 2405 1975
rect 2523 1845 2533 1955
rect 2875 1945 2885 2135
rect 2907 1645 2917 2275
rect 2427 905 2437 1515
rect 2619 1465 2629 1475
rect 2565 1455 2629 1465
rect 2619 1425 2629 1435
rect 2491 1415 2629 1425
rect 2491 1325 2501 1415
rect 3355 1385 3365 1435
rect 2523 1375 2597 1385
rect 2523 1365 2533 1375
rect 2587 1365 2597 1375
rect 2555 925 2565 1355
rect 3387 1265 3397 2555
rect 2587 1055 2699 1065
rect 2587 1045 2597 1055
rect 2747 1005 2757 1055
rect 2939 985 2949 995
rect 2907 975 2949 985
rect 2907 965 2917 975
rect 2555 345 2565 915
rect 3355 565 3365 595
rect 3387 365 3397 915
rect 3419 885 3429 1275
rect 3579 925 3589 2155
rect 3611 1605 3621 2115
rect 3707 1545 3717 1615
rect 3579 905 3589 915
rect 1221 335 1285 345
rect 1275 325 1285 335
rect 1883 205 1893 235
rect 3611 105 3621 1535
rect 4091 1365 4101 2755
rect 3771 485 3781 555
rect 4091 105 4101 975
rect 4155 185 4165 2955
rect 4187 105 4197 1615
use NAND2X1  NAND2X1_294
timestamp 1598351757
transform -1 0 4232 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_245
timestamp 1598351757
transform 1 0 4152 0 -1 3010
box -18 -6 52 210
use FILL  FILL_15_2
timestamp 1598351757
transform -1 0 4264 0 -1 3010
box -16 -6 32 210
use FILL  FILL_15_1
timestamp 1598351757
transform -1 0 4248 0 -1 3010
box -16 -6 32 210
use NAND2X1  NAND2X1_577
timestamp 1598351757
transform -1 0 4120 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_14
timestamp 1598351757
transform -1 0 4040 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_443
timestamp 1598351757
transform -1 0 4152 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_22
timestamp 1598351757
transform -1 0 4072 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_5
timestamp 1598351757
transform -1 0 3928 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_23
timestamp 1598351757
transform 1 0 3960 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_10
timestamp 1598351757
transform -1 0 3960 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_9
timestamp 1598351757
transform -1 0 3880 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_82
timestamp 1598351757
transform -1 0 3816 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_21
timestamp 1598351757
transform -1 0 3848 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_83
timestamp 1598351757
transform -1 0 3768 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_84
timestamp 1598351757
transform 1 0 3704 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_83
timestamp 1598351757
transform 1 0 3656 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_19
timestamp 1598351757
transform 1 0 3608 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_28
timestamp 1598351757
transform 1 0 3576 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_27
timestamp 1598351757
transform -1 0 3576 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_20
timestamp 1598351757
transform 1 0 3464 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_33
timestamp 1598351757
transform -1 0 3464 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_13
timestamp 1598351757
transform -1 0 3544 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_42
timestamp 1598351757
transform -1 0 3416 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_126
timestamp 1598351757
transform -1 0 3384 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_84
timestamp 1598351757
transform 1 0 3224 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_117
timestamp 1598351757
transform -1 0 3336 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_183
timestamp 1598351757
transform -1 0 3304 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_81
timestamp 1598351757
transform -1 0 3224 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_80
timestamp 1598351757
transform 1 0 3064 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_82
timestamp 1598351757
transform -1 0 3176 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_81
timestamp 1598351757
transform 1 0 3112 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_214
timestamp 1598351757
transform -1 0 2968 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_72
timestamp 1598351757
transform -1 0 3064 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_366
timestamp 1598351757
transform 1 0 3000 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_85
timestamp 1598351757
transform -1 0 3000 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_85
timestamp 1598351757
transform 1 0 2840 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_35
timestamp 1598351757
transform -1 0 2808 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_184
timestamp 1598351757
transform 1 0 2888 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_86
timestamp 1598351757
transform -1 0 2840 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_208
timestamp 1598351757
transform 1 0 2680 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_219
timestamp 1598351757
transform -1 0 2648 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_190
timestamp 1598351757
transform -1 0 2760 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_44
timestamp 1598351757
transform -1 0 2680 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_222
timestamp 1598351757
transform -1 0 2568 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_699
timestamp 1598351757
transform -1 0 2520 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_195
timestamp 1598351757
transform -1 0 2600 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_748
timestamp 1598351757
transform -1 0 2440 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_789
timestamp 1598351757
transform -1 0 2360 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_543
timestamp 1598351757
transform -1 0 2472 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_191
timestamp 1598351757
transform 1 0 2360 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_751
timestamp 1598351757
transform 1 0 2264 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_215
timestamp 1598351757
transform 1 0 2184 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_182
timestamp 1598351757
transform -1 0 2264 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_181
timestamp 1598351757
transform 1 0 2152 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_205
timestamp 1598351757
transform -1 0 2152 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_86
timestamp 1598351757
transform 1 0 2056 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_235
timestamp 1598351757
transform -1 0 2056 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_786
timestamp 1598351757
transform -1 0 2008 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_204
timestamp 1598351757
transform 1 0 1848 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_616
timestamp 1598351757
transform -1 0 1960 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_180
timestamp 1598351757
transform 1 0 1896 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_79
timestamp 1598351757
transform -1 0 1848 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_243
timestamp 1598351757
transform -1 0 1768 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_210
timestamp 1598351757
transform 1 0 1768 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_198
timestamp 1598351757
transform -1 0 1720 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_767
timestamp 1598351757
transform -1 0 1688 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_773
timestamp 1598351757
transform -1 0 1640 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_223
timestamp 1598351757
transform 1 0 1544 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_232
timestamp 1598351757
transform -1 0 1512 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_240
timestamp 1598351757
transform -1 0 1464 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_207
timestamp 1598351757
transform 1 0 1512 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_601
timestamp 1598351757
transform -1 0 1416 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_793
timestamp 1598351757
transform -1 0 1352 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_619
timestamp 1598351757
transform -1 0 1384 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_623
timestamp 1598351757
transform -1 0 1304 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_599
timestamp 1598351757
transform 1 0 1240 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_771
timestamp 1598351757
transform 1 0 1192 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_764
timestamp 1598351757
transform -1 0 1160 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_597
timestamp 1598351757
transform 1 0 1160 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_769
timestamp 1598351757
transform 1 0 1064 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_763
timestamp 1598351757
transform 1 0 1016 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_380
timestamp 1598351757
transform -1 0 1016 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_311
timestamp 1598351757
transform -1 0 968 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_379
timestamp 1598351757
transform 1 0 888 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_460
timestamp 1598351757
transform -1 0 888 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_48
timestamp 1598351757
transform 1 0 808 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_40
timestamp 1598351757
transform 1 0 760 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_762
timestamp 1598351757
transform 1 0 616 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_6
timestamp 1598351757
transform 1 0 728 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_33
timestamp 1598351757
transform 1 0 696 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_595
timestamp 1598351757
transform 1 0 664 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_25
timestamp 1598351757
transform -1 0 616 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_3
timestamp 1598351757
transform 1 0 488 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_25
timestamp 1598351757
transform 1 0 536 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_17
timestamp 1598351757
transform 1 0 376 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_34
timestamp 1598351757
transform 1 0 456 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_1
timestamp 1598351757
transform 1 0 424 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_3
timestamp 1598351757
transform 1 0 344 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_2
timestamp 1598351757
transform 1 0 296 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_1
timestamp 1598351757
transform 1 0 184 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_4
timestamp 1598351757
transform 1 0 264 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_5
timestamp 1598351757
transform 1 0 232 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_56
timestamp 1598351757
transform 1 0 8 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_50
timestamp 1598351757
transform 1 0 40 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_2
timestamp 1598351757
transform 1 0 152 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_57
timestamp 1598351757
transform -1 0 152 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_55
timestamp 1598351757
transform 1 0 88 0 -1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_401
timestamp 1598351757
transform -1 0 4232 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_395
timestamp 1598351757
transform 1 0 4184 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_396
timestamp 1598351757
transform -1 0 4184 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_325
timestamp 1598351757
transform -1 0 4184 0 1 2610
box -18 -6 52 210
use FILL  FILL_14_2
timestamp 1598351757
transform 1 0 4248 0 1 2610
box -16 -6 32 210
use FILL  FILL_14_1
timestamp 1598351757
transform 1 0 4232 0 1 2610
box -16 -6 32 210
use FILL  FILL_13_2
timestamp 1598351757
transform -1 0 4264 0 -1 2610
box -16 -6 32 210
use FILL  FILL_13_1
timestamp 1598351757
transform -1 0 4248 0 -1 2610
box -16 -6 32 210
use NAND2X1  NAND2X1_37
timestamp 1598351757
transform 1 0 4072 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_402
timestamp 1598351757
transform 1 0 3992 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_199
timestamp 1598351757
transform -1 0 4136 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_207
timestamp 1598351757
transform -1 0 4024 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_46
timestamp 1598351757
transform -1 0 4152 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_326
timestamp 1598351757
transform 1 0 4040 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_172
timestamp 1598351757
transform 1 0 4056 0 -1 2610
box -18 -6 52 210
use INVX1  INVX1_175
timestamp 1598351757
transform -1 0 4056 0 -1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_397
timestamp 1598351757
transform -1 0 3992 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_6
timestamp 1598351757
transform -1 0 3944 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_404
timestamp 1598351757
transform -1 0 3896 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_398
timestamp 1598351757
transform 1 0 3896 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_11
timestamp 1598351757
transform -1 0 3976 0 -1 2610
box -18 -6 52 210
use INVX1  INVX1_328
timestamp 1598351757
transform 1 0 3864 0 -1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_403
timestamp 1598351757
transform -1 0 3816 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_400
timestamp 1598351757
transform 1 0 3688 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_399
timestamp 1598351757
transform -1 0 3864 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_236
timestamp 1598351757
transform -1 0 3784 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_324
timestamp 1598351757
transform 1 0 3816 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_327
timestamp 1598351757
transform -1 0 3768 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_322
timestamp 1598351757
transform 1 0 3784 0 -1 2610
box -18 -6 52 210
use INVX1  INVX1_206
timestamp 1598351757
transform -1 0 3736 0 -1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_394
timestamp 1598351757
transform 1 0 3640 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_49
timestamp 1598351757
transform -1 0 3640 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_393
timestamp 1598351757
transform 1 0 3656 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_48
timestamp 1598351757
transform -1 0 3656 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_196
timestamp 1598351757
transform 1 0 3560 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_54
timestamp 1598351757
transform -1 0 3592 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_530
timestamp 1598351757
transform -1 0 3560 0 -1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_671
timestamp 1598351757
transform 1 0 3512 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_8
timestamp 1598351757
transform -1 0 3512 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_24
timestamp 1598351757
transform -1 0 3528 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_617
timestamp 1598351757
transform -1 0 3480 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_12
timestamp 1598351757
transform -1 0 3464 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_305
timestamp 1598351757
transform 1 0 3400 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_483
timestamp 1598351757
transform -1 0 3432 0 -1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_375
timestamp 1598351757
transform -1 0 3400 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_376
timestamp 1598351757
transform 1 0 3272 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_459
timestamp 1598351757
transform -1 0 3272 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_621
timestamp 1598351757
transform 1 0 3352 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_672
timestamp 1598351757
transform 1 0 3304 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_202
timestamp 1598351757
transform -1 0 3304 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_306
timestamp 1598351757
transform 1 0 3320 0 1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_463
timestamp 1598351757
transform -1 0 3192 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_68
timestamp 1598351757
transform 1 0 3064 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_69
timestamp 1598351757
transform 1 0 3208 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_616
timestamp 1598351757
transform 1 0 3160 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_377
timestamp 1598351757
transform 1 0 3080 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_365
timestamp 1598351757
transform -1 0 3224 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_73
timestamp 1598351757
transform -1 0 3144 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_308
timestamp 1598351757
transform -1 0 3160 0 -1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_378
timestamp 1598351757
transform 1 0 2984 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_263
timestamp 1598351757
transform 1 0 3000 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_104
timestamp 1598351757
transform 1 0 2952 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_307
timestamp 1598351757
transform -1 0 3064 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_309
timestamp 1598351757
transform 1 0 2952 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_389
timestamp 1598351757
transform -1 0 2952 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_100
timestamp 1598351757
transform 1 0 3048 0 -1 2610
box -18 -6 52 210
use INVX1  INVX1_223
timestamp 1598351757
transform -1 0 2952 0 -1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_490
timestamp 1598351757
transform -1 0 2920 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_34
timestamp 1598351757
transform -1 0 2872 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_32
timestamp 1598351757
transform -1 0 2824 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_27
timestamp 1598351757
transform -1 0 2920 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_57
timestamp 1598351757
transform -1 0 2872 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_198
timestamp 1598351757
transform -1 0 2824 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_750
timestamp 1598351757
transform -1 0 2680 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_749
timestamp 1598351757
transform -1 0 2744 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_813
timestamp 1598351757
transform 1 0 2648 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_43
timestamp 1598351757
transform -1 0 2776 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_174
timestamp 1598351757
transform -1 0 2744 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_586
timestamp 1598351757
transform -1 0 2712 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_585
timestamp 1598351757
transform -1 0 2776 0 -1 2610
box -18 -6 52 210
use INVX1  INVX1_642
timestamp 1598351757
transform 1 0 2616 0 -1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_29
timestamp 1598351757
transform 1 0 2552 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_316
timestamp 1598351757
transform -1 0 2520 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_266
timestamp 1598351757
transform 1 0 2536 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_58
timestamp 1598351757
transform -1 0 2504 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_39
timestamp 1598351757
transform -1 0 2632 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_38
timestamp 1598351757
transform -1 0 2552 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_229
timestamp 1598351757
transform -1 0 2616 0 -1 2610
box -18 -6 52 210
use INVX1  INVX1_228
timestamp 1598351757
transform -1 0 2536 0 -1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_87
timestamp 1598351757
transform 1 0 2328 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_61
timestamp 1598351757
transform -1 0 2424 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_60
timestamp 1598351757
transform -1 0 2344 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_87
timestamp 1598351757
transform -1 0 2472 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_178
timestamp 1598351757
transform -1 0 2440 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_88
timestamp 1598351757
transform -1 0 2408 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_552
timestamp 1598351757
transform -1 0 2456 0 -1 2610
box -18 -6 52 210
use INVX1  INVX1_64
timestamp 1598351757
transform -1 0 2376 0 -1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_206
timestamp 1598351757
transform 1 0 2280 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_88
timestamp 1598351757
transform -1 0 2216 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_201
timestamp 1598351757
transform -1 0 2296 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_65
timestamp 1598351757
transform 1 0 2200 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_339
timestamp 1598351757
transform -1 0 2200 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_177
timestamp 1598351757
transform 1 0 2248 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_179
timestamp 1598351757
transform -1 0 2248 0 1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_100
timestamp 1598351757
transform -1 0 2168 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_340
timestamp 1598351757
transform -1 0 2088 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_262
timestamp 1598351757
transform 1 0 2104 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_224
timestamp 1598351757
transform -1 0 2104 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_227
timestamp 1598351757
transform -1 0 2056 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_205
timestamp 1598351757
transform -1 0 2120 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_201
timestamp 1598351757
transform 1 0 2008 0 1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_795
timestamp 1598351757
transform -1 0 1976 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_502
timestamp 1598351757
transform 1 0 1848 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_226
timestamp 1598351757
transform 1 0 1928 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_509
timestamp 1598351757
transform -1 0 1928 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_615
timestamp 1598351757
transform -1 0 2008 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_395
timestamp 1598351757
transform -1 0 1928 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_399
timestamp 1598351757
transform -1 0 2008 0 -1 2610
box -18 -6 52 210
use INVX1  INVX1_97
timestamp 1598351757
transform -1 0 1880 0 -1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_244
timestamp 1598351757
transform 1 0 1736 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_785
timestamp 1598351757
transform 1 0 1800 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_503
timestamp 1598351757
transform -1 0 1800 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_394
timestamp 1598351757
transform 1 0 1816 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_600
timestamp 1598351757
transform -1 0 1816 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_274
timestamp 1598351757
transform -1 0 1736 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_208
timestamp 1598351757
transform 1 0 1720 0 -1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_78
timestamp 1598351757
transform -1 0 1640 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_241
timestamp 1598351757
transform -1 0 1720 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_242
timestamp 1598351757
transform 1 0 1624 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_776
timestamp 1598351757
transform 1 0 1544 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_209
timestamp 1598351757
transform 1 0 1672 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_79
timestamp 1598351757
transform -1 0 1672 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_80
timestamp 1598351757
transform 1 0 1560 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_604
timestamp 1598351757
transform 1 0 1592 0 -1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_350
timestamp 1598351757
transform -1 0 1528 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_233
timestamp 1598351757
transform -1 0 1448 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_238
timestamp 1598351757
transform 1 0 1496 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_164
timestamp 1598351757
transform -1 0 1496 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_275
timestamp 1598351757
transform -1 0 1560 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_273
timestamp 1598351757
transform -1 0 1480 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_284
timestamp 1598351757
transform -1 0 1448 0 -1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_234
timestamp 1598351757
transform 1 0 1320 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_351
timestamp 1598351757
transform 1 0 1240 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_757
timestamp 1598351757
transform 1 0 1368 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_358
timestamp 1598351757
transform -1 0 1368 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_204
timestamp 1598351757
transform -1 0 1400 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_620
timestamp 1598351757
transform 1 0 1288 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_285
timestamp 1598351757
transform 1 0 1288 0 -1 2610
box -18 -6 52 210
use INVX1  INVX1_292
timestamp 1598351757
transform -1 0 1288 0 -1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_774
timestamp 1598351757
transform -1 0 1240 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_792
timestamp 1598351757
transform -1 0 1160 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_758
timestamp 1598351757
transform -1 0 1224 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_759
timestamp 1598351757
transform 1 0 1128 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_766
timestamp 1598351757
transform -1 0 1128 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_598
timestamp 1598351757
transform 1 0 1160 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_622
timestamp 1598351757
transform -1 0 1112 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_591
timestamp 1598351757
transform -1 0 1256 0 -1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_805
timestamp 1598351757
transform -1 0 1080 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_824
timestamp 1598351757
transform 1 0 920 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_770
timestamp 1598351757
transform 1 0 1032 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_765
timestamp 1598351757
transform -1 0 1032 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_755
timestamp 1598351757
transform -1 0 984 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_621
timestamp 1598351757
transform 1 0 1000 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_63
timestamp 1598351757
transform 1 0 968 0 1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_59
timestamp 1598351757
transform 1 0 840 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_791
timestamp 1598351757
transform -1 0 936 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_12
timestamp 1598351757
transform 1 0 808 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_310
timestamp 1598351757
transform -1 0 920 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_35
timestamp 1598351757
transform 1 0 808 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_20
timestamp 1598351757
transform 1 0 856 0 -1 2610
box -18 -6 52 210
use INVX1  INVX1_53
timestamp 1598351757
transform 1 0 776 0 -1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_26
timestamp 1598351757
transform 1 0 760 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_22
timestamp 1598351757
transform -1 0 760 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_47
timestamp 1598351757
transform -1 0 712 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_18
timestamp 1598351757
transform -1 0 744 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_145
timestamp 1598351757
transform 1 0 632 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_31
timestamp 1598351757
transform 1 0 744 0 -1 2610
box -18 -6 52 210
use INVX1  INVX1_26
timestamp 1598351757
transform -1 0 696 0 -1 2610
box -18 -6 52 210
use INVX1  INVX1_93
timestamp 1598351757
transform 1 0 632 0 -1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_31
timestamp 1598351757
transform -1 0 632 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_157
timestamp 1598351757
transform 1 0 504 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_44
timestamp 1598351757
transform 1 0 552 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_409
timestamp 1598351757
transform 1 0 504 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_41
timestamp 1598351757
transform -1 0 584 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_334
timestamp 1598351757
transform -1 0 504 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_50
timestamp 1598351757
transform 1 0 600 0 -1 2610
box -18 -6 52 210
use INVX1  INVX1_333
timestamp 1598351757
transform 1 0 472 0 -1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_408
timestamp 1598351757
transform -1 0 472 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_36
timestamp 1598351757
transform 1 0 376 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_581
timestamp 1598351757
transform -1 0 376 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_95
timestamp 1598351757
transform 1 0 360 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_587
timestamp 1598351757
transform 1 0 312 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_74
timestamp 1598351757
transform 1 0 440 0 -1 2610
box -18 -6 52 210
use INVX1  INVX1_45
timestamp 1598351757
transform 1 0 408 0 -1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_70
timestamp 1598351757
transform -1 0 328 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_11
timestamp 1598351757
transform 1 0 200 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_429
timestamp 1598351757
transform 1 0 200 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_18
timestamp 1598351757
transform 1 0 248 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_19
timestamp 1598351757
transform 1 0 168 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_456
timestamp 1598351757
transform 1 0 280 0 -1 2610
box -18 -6 52 210
use INVX1  INVX1_69
timestamp 1598351757
transform 1 0 248 0 -1 2610
box -18 -6 52 210
use INVX1  INVX1_343
timestamp 1598351757
transform 1 0 168 0 -1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_21
timestamp 1598351757
transform 1 0 8 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_30
timestamp 1598351757
transform 1 0 8 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_64
timestamp 1598351757
transform 1 0 120 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_51
timestamp 1598351757
transform 1 0 88 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_29
timestamp 1598351757
transform 1 0 88 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_30
timestamp 1598351757
transform -1 0 88 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_58
timestamp 1598351757
transform 1 0 136 0 -1 2610
box -18 -6 52 210
use INVX1  INVX1_40
timestamp 1598351757
transform 1 0 56 0 -1 2610
box -18 -6 52 210
use INVX1  INVX1_70
timestamp 1598351757
transform -1 0 4264 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_66
timestamp 1598351757
transform -1 0 4232 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_71
timestamp 1598351757
transform 1 0 4152 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_625
timestamp 1598351757
transform -1 0 4152 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_530
timestamp 1598351757
transform -1 0 4104 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_171
timestamp 1598351757
transform 1 0 4024 0 1 2210
box -18 -6 52 210
use INVX1  INVX1_323
timestamp 1598351757
transform -1 0 4024 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_195
timestamp 1598351757
transform 1 0 3912 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_41
timestamp 1598351757
transform -1 0 3912 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_176
timestamp 1598351757
transform 1 0 3960 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_43
timestamp 1598351757
transform -1 0 3864 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_627
timestamp 1598351757
transform 1 0 3768 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_629
timestamp 1598351757
transform 1 0 3720 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_23
timestamp 1598351757
transform -1 0 3720 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_626
timestamp 1598351757
transform 1 0 3560 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_32
timestamp 1598351757
transform -1 0 3672 0 1 2210
box -18 -6 52 210
use INVX1  INVX1_170
timestamp 1598351757
transform -1 0 3640 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_200
timestamp 1598351757
transform 1 0 3512 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_618
timestamp 1598351757
transform -1 0 3480 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_481
timestamp 1598351757
transform -1 0 3512 0 1 2210
box -18 -6 52 210
use INVX1  INVX1_480
timestamp 1598351757
transform -1 0 3432 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_622
timestamp 1598351757
transform 1 0 3352 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_619
timestamp 1598351757
transform 1 0 3304 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_67
timestamp 1598351757
transform 1 0 3224 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_169
timestamp 1598351757
transform 1 0 3272 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_487
timestamp 1598351757
transform -1 0 3224 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_489
timestamp 1598351757
transform -1 0 3176 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_557
timestamp 1598351757
transform -1 0 3128 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_488
timestamp 1598351757
transform -1 0 3080 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_670
timestamp 1598351757
transform -1 0 3032 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_673
timestamp 1598351757
transform -1 0 2984 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_38
timestamp 1598351757
transform 1 0 2824 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_536
timestamp 1598351757
transform -1 0 2824 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_531
timestamp 1598351757
transform -1 0 2936 0 1 2210
box -18 -6 52 210
use INVX1  INVX1_47
timestamp 1598351757
transform 1 0 2872 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_537
timestamp 1598351757
transform 1 0 2696 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_197
timestamp 1598351757
transform 1 0 2648 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_845
timestamp 1598351757
transform 1 0 2600 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_173
timestamp 1598351757
transform 1 0 2744 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_52
timestamp 1598351757
transform 1 0 2552 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_385
timestamp 1598351757
transform 1 0 2504 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_389
timestamp 1598351757
transform -1 0 2504 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_318
timestamp 1598351757
transform 1 0 2408 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_709
timestamp 1598351757
transform 1 0 2360 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_698
timestamp 1598351757
transform 1 0 2312 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_63
timestamp 1598351757
transform -1 0 2312 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_504
timestamp 1598351757
transform 1 0 2184 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_68
timestamp 1598351757
transform -1 0 2264 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_507
timestamp 1598351757
transform -1 0 2184 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_445
timestamp 1598351757
transform 1 0 2088 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_505
timestamp 1598351757
transform -1 0 2088 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_237
timestamp 1598351757
transform -1 0 2040 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_510
timestamp 1598351757
transform 1 0 1944 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_398
timestamp 1598351757
transform 1 0 1912 0 1 2210
box -18 -6 52 210
use INVX1  INVX1_397
timestamp 1598351757
transform -1 0 1912 0 1 2210
box -18 -6 52 210
use INVX1  INVX1_589
timestamp 1598351757
transform -1 0 1880 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_508
timestamp 1598351757
transform 1 0 1800 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_756
timestamp 1598351757
transform -1 0 1800 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_590
timestamp 1598351757
transform 1 0 1720 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_101
timestamp 1598351757
transform 1 0 1672 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_168
timestamp 1598351757
transform 1 0 1624 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_239
timestamp 1598351757
transform -1 0 1592 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_396
timestamp 1598351757
transform 1 0 1592 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_506
timestamp 1598351757
transform -1 0 1544 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_229
timestamp 1598351757
transform 1 0 1384 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_96
timestamp 1598351757
transform 1 0 1464 0 1 2210
box -18 -6 52 210
use INVX1  INVX1_94
timestamp 1598351757
transform -1 0 1464 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_99
timestamp 1598351757
transform -1 0 1384 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_419
timestamp 1598351757
transform -1 0 1336 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_95
timestamp 1598351757
transform 1 0 1256 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_447
timestamp 1598351757
transform -1 0 1256 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_420
timestamp 1598351757
transform 1 0 1160 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_592
timestamp 1598351757
transform 1 0 1128 0 1 2210
box -18 -6 52 210
use INVX1  INVX1_291
timestamp 1598351757
transform -1 0 1128 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_364
timestamp 1598351757
transform -1 0 1096 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_387
timestamp 1598351757
transform -1 0 1048 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_721
timestamp 1598351757
transform -1 0 1000 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_272
timestamp 1598351757
transform 1 0 920 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_720
timestamp 1598351757
transform 1 0 840 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_669
timestamp 1598351757
transform -1 0 840 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_563
timestamp 1598351757
transform 1 0 888 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_291
timestamp 1598351757
transform -1 0 792 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_668
timestamp 1598351757
transform -1 0 712 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_528
timestamp 1598351757
transform -1 0 744 0 1 2210
box -18 -6 52 210
use INVX1  INVX1_529
timestamp 1598351757
transform 1 0 632 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_826
timestamp 1598351757
transform 1 0 584 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_588
timestamp 1598351757
transform -1 0 552 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_315
timestamp 1598351757
transform 1 0 552 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_386
timestamp 1598351757
transform 1 0 456 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_836
timestamp 1598351757
transform -1 0 424 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_823
timestamp 1598351757
transform 1 0 328 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_455
timestamp 1598351757
transform 1 0 424 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_752
timestamp 1598351757
transform 1 0 280 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_425
timestamp 1598351757
transform 1 0 232 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_316
timestamp 1598351757
transform 1 0 200 0 1 2210
box -18 -6 52 210
use INVX1  INVX1_341
timestamp 1598351757
transform -1 0 200 0 1 2210
box -18 -6 52 210
use INVX1  INVX1_262
timestamp 1598351757
transform 1 0 8 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_53
timestamp 1598351757
transform 1 0 120 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_328
timestamp 1598351757
transform 1 0 40 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_60
timestamp 1598351757
transform 1 0 88 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_549
timestamp 1598351757
transform 1 0 4168 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_423
timestamp 1598351757
transform 1 0 4216 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_422
timestamp 1598351757
transform 1 0 4136 0 -1 2210
box -18 -6 52 210
use FILL  FILL_11_1
timestamp 1598351757
transform -1 0 4264 0 -1 2210
box -16 -6 32 210
use NAND2X1  NAND2X1_529
timestamp 1598351757
transform 1 0 4088 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_548
timestamp 1598351757
transform -1 0 4088 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_7
timestamp 1598351757
transform 1 0 4008 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_4
timestamp 1598351757
transform 1 0 3960 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_531
timestamp 1598351757
transform 1 0 3880 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_8
timestamp 1598351757
transform 1 0 3928 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_488
timestamp 1598351757
transform 1 0 3848 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_630
timestamp 1598351757
transform 1 0 3800 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_628
timestamp 1598351757
transform 1 0 3720 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_39
timestamp 1598351757
transform -1 0 3720 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_487
timestamp 1598351757
transform 1 0 3768 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_194
timestamp 1598351757
transform -1 0 3672 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_16
timestamp 1598351757
transform -1 0 3624 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_37
timestamp 1598351757
transform -1 0 3576 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_28
timestamp 1598351757
transform -1 0 3544 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_36
timestamp 1598351757
transform -1 0 3496 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_369
timestamp 1598351757
transform 1 0 3432 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_90
timestamp 1598351757
transform 1 0 3400 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_92
timestamp 1598351757
transform 1 0 3352 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_624
timestamp 1598351757
transform -1 0 3288 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_486
timestamp 1598351757
transform 1 0 3320 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_484
timestamp 1598351757
transform -1 0 3320 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_623
timestamp 1598351757
transform 1 0 3160 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_772
timestamp 1598351757
transform -1 0 3128 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_485
timestamp 1598351757
transform 1 0 3208 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_388
timestamp 1598351757
transform -1 0 3160 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_383
timestamp 1598351757
transform 1 0 2968 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_431
timestamp 1598351757
transform 1 0 3048 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_314
timestamp 1598351757
transform -1 0 3048 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_313
timestamp 1598351757
transform 1 0 2936 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_615
timestamp 1598351757
transform -1 0 2904 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_193
timestamp 1598351757
transform 1 0 2808 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_7
timestamp 1598351757
transform 1 0 2760 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_211
timestamp 1598351757
transform 1 0 2904 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_228
timestamp 1598351757
transform -1 0 2728 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_410
timestamp 1598351757
transform 1 0 2728 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_202
timestamp 1598351757
transform -1 0 2680 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_666
timestamp 1598351757
transform 1 0 2616 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_56
timestamp 1598351757
transform 1 0 2568 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_72
timestamp 1598351757
transform 1 0 2488 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_400
timestamp 1598351757
transform 1 0 2536 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_318
timestamp 1598351757
transform -1 0 2488 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_203
timestamp 1598351757
transform -1 0 2392 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_455
timestamp 1598351757
transform -1 0 2344 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_254
timestamp 1598351757
transform -1 0 2456 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_551
timestamp 1598351757
transform 1 0 2392 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_614
timestamp 1598351757
transform -1 0 2232 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_351
timestamp 1598351757
transform 1 0 2264 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_478
timestamp 1598351757
transform 1 0 2232 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_479
timestamp 1598351757
transform 1 0 2152 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_76
timestamp 1598351757
transform 1 0 2072 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_74
timestamp 1598351757
transform 1 0 2024 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_77
timestamp 1598351757
transform 1 0 2120 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_754
timestamp 1598351757
transform 1 0 1976 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_289
timestamp 1598351757
transform -1 0 1976 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_97
timestamp 1598351757
transform -1 0 1896 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_98
timestamp 1598351757
transform 1 0 1896 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_89
timestamp 1598351757
transform 1 0 1800 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_94
timestamp 1598351757
transform -1 0 1800 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_230
timestamp 1598351757
transform -1 0 1752 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_165
timestamp 1598351757
transform 1 0 1656 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_341
timestamp 1598351757
transform -1 0 1592 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_153
timestamp 1598351757
transform -1 0 1656 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_91
timestamp 1598351757
transform -1 0 1624 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_231
timestamp 1598351757
transform 1 0 1464 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_357
timestamp 1598351757
transform 1 0 1416 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_203
timestamp 1598351757
transform 1 0 1512 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_524
timestamp 1598351757
transform -1 0 1416 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_96
timestamp 1598351757
transform -1 0 1352 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_98
timestamp 1598351757
transform -1 0 1304 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_525
timestamp 1598351757
transform -1 0 1384 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_790
timestamp 1598351757
transform 1 0 1208 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_93
timestamp 1598351757
transform -1 0 1208 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_664
timestamp 1598351757
transform -1 0 1160 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_667
timestamp 1598351757
transform 1 0 1064 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_333
timestamp 1598351757
transform -1 0 1064 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_267
timestamp 1598351757
transform -1 0 1016 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_564
timestamp 1598351757
transform 1 0 952 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_338
timestamp 1598351757
transform -1 0 952 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_825
timestamp 1598351757
transform 1 0 824 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_753
timestamp 1598351757
transform 1 0 776 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_635
timestamp 1598351757
transform -1 0 904 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_837
timestamp 1598351757
transform -1 0 744 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_827
timestamp 1598351757
transform -1 0 664 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_59
timestamp 1598351757
transform 1 0 744 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_658
timestamp 1598351757
transform -1 0 696 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_838
timestamp 1598351757
transform -1 0 616 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_821
timestamp 1598351757
transform -1 0 536 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_587
timestamp 1598351757
transform 1 0 536 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_835
timestamp 1598351757
transform -1 0 488 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_822
timestamp 1598351757
transform -1 0 440 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_656
timestamp 1598351757
transform -1 0 392 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_657
timestamp 1598351757
transform -1 0 360 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_839
timestamp 1598351757
transform -1 0 328 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_602
timestamp 1598351757
transform 1 0 248 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_342
timestamp 1598351757
transform 1 0 216 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_298
timestamp 1598351757
transform -1 0 216 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_852
timestamp 1598351757
transform -1 0 56 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_660
timestamp 1598351757
transform -1 0 184 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_261
timestamp 1598351757
transform 1 0 120 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_659
timestamp 1598351757
transform -1 0 120 0 -1 2210
box -18 -6 52 210
use INVX1  INVX1_673
timestamp 1598351757
transform 1 0 56 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_479
timestamp 1598351757
transform -1 0 4232 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_382
timestamp 1598351757
transform 1 0 4152 0 1 1810
box -18 -6 52 210
use FILL  FILL_10_2
timestamp 1598351757
transform 1 0 4248 0 1 1810
box -16 -6 32 210
use FILL  FILL_10_1
timestamp 1598351757
transform 1 0 4232 0 1 1810
box -16 -6 32 210
use NAND2X1  NAND2X1_414
timestamp 1598351757
transform -1 0 4120 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_415
timestamp 1598351757
transform -1 0 4040 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_381
timestamp 1598351757
transform 1 0 4120 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_339
timestamp 1598351757
transform 1 0 4040 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_293
timestamp 1598351757
transform 1 0 3912 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_42
timestamp 1598351757
transform -1 0 3912 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_243
timestamp 1598351757
transform 1 0 3960 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_49
timestamp 1598351757
transform -1 0 3864 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_472
timestamp 1598351757
transform 1 0 3784 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_297
timestamp 1598351757
transform -1 0 3752 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_368
timestamp 1598351757
transform -1 0 3784 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_347
timestamp 1598351757
transform -1 0 3704 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_268
timestamp 1598351757
transform -1 0 3592 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_280
timestamp 1598351757
transform -1 0 3656 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_281
timestamp 1598351757
transform -1 0 3624 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_363
timestamp 1598351757
transform 1 0 3496 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_360
timestamp 1598351757
transform 1 0 3416 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_294
timestamp 1598351757
transform 1 0 3464 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_224
timestamp 1598351757
transform -1 0 3416 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_381
timestamp 1598351757
transform -1 0 3352 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_475
timestamp 1598351757
transform 1 0 3256 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_297
timestamp 1598351757
transform -1 0 3384 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_380
timestamp 1598351757
transform 1 0 3224 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_474
timestamp 1598351757
transform 1 0 3176 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_860
timestamp 1598351757
transform 1 0 3128 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_482
timestamp 1598351757
transform -1 0 3128 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_596
timestamp 1598351757
transform -1 0 3096 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_366
timestamp 1598351757
transform 1 0 2984 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_321
timestamp 1598351757
transform 1 0 3032 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_296
timestamp 1598351757
transform 1 0 2952 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_561
timestamp 1598351757
transform -1 0 2952 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_384
timestamp 1598351757
transform -1 0 2904 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_494
timestamp 1598351757
transform 1 0 2808 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_432
timestamp 1598351757
transform 1 0 2776 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_392
timestamp 1598351757
transform 1 0 2696 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_320
timestamp 1598351757
transform -1 0 2776 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_194
timestamp 1598351757
transform -1 0 2696 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_319
timestamp 1598351757
transform 1 0 2632 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_492
timestamp 1598351757
transform -1 0 2632 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_493
timestamp 1598351757
transform 1 0 2536 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_491
timestamp 1598351757
transform 1 0 2488 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_133
timestamp 1598351757
transform 1 0 2440 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_267
timestamp 1598351757
transform 1 0 2360 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_390
timestamp 1598351757
transform 1 0 2312 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_123
timestamp 1598351757
transform -1 0 2440 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_13
timestamp 1598351757
transform 1 0 2264 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_71
timestamp 1598351757
transform 1 0 2216 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_304
timestamp 1598351757
transform 1 0 2168 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_315
timestamp 1598351757
transform 1 0 2056 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_266
timestamp 1598351757
transform 1 0 2136 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_317
timestamp 1598351757
transform 1 0 2104 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_270
timestamp 1598351757
transform -1 0 2056 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_309
timestamp 1598351757
transform -1 0 2024 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_335
timestamp 1598351757
transform -1 0 1976 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_310
timestamp 1598351757
transform -1 0 1928 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_91
timestamp 1598351757
transform 1 0 1832 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_75
timestamp 1598351757
transform 1 0 1688 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_603
timestamp 1598351757
transform -1 0 1832 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_92
timestamp 1598351757
transform -1 0 1800 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_269
timestamp 1598351757
transform -1 0 1768 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_337
timestamp 1598351757
transform -1 0 1656 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_170
timestamp 1598351757
transform -1 0 1576 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_160
timestamp 1598351757
transform -1 0 1688 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_154
timestamp 1598351757
transform -1 0 1608 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_352
timestamp 1598351757
transform 1 0 1384 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_155
timestamp 1598351757
transform -1 0 1528 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_287
timestamp 1598351757
transform -1 0 1496 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_271
timestamp 1598351757
transform -1 0 1464 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_117
timestamp 1598351757
transform -1 0 1352 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_265
timestamp 1598351757
transform 1 0 1224 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_286
timestamp 1598351757
transform -1 0 1384 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_227
timestamp 1598351757
transform -1 0 1304 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_641
timestamp 1598351757
transform -1 0 1224 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_212
timestamp 1598351757
transform -1 0 1176 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_527
timestamp 1598351757
transform -1 0 1128 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_422
timestamp 1598351757
transform 1 0 1048 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_734
timestamp 1598351757
transform -1 0 1016 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_211
timestamp 1598351757
transform -1 0 968 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_187
timestamp 1598351757
transform 1 0 1016 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_171
timestamp 1598351757
transform 1 0 840 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_853
timestamp 1598351757
transform -1 0 840 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_157
timestamp 1598351757
transform 1 0 888 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_334
timestamp 1598351757
transform 1 0 680 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_290
timestamp 1598351757
transform 1 0 632 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_268
timestamp 1598351757
transform 1 0 760 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_566
timestamp 1598351757
transform -1 0 760 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_733
timestamp 1598351757
transform 1 0 584 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_665
timestamp 1598351757
transform 1 0 504 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_565
timestamp 1598351757
transform 1 0 552 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_719
timestamp 1598351757
transform -1 0 504 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_807
timestamp 1598351757
transform 1 0 376 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_636
timestamp 1598351757
transform -1 0 456 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_674
timestamp 1598351757
transform -1 0 376 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_300
timestamp 1598351757
transform -1 0 344 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_430
timestamp 1598351757
transform -1 0 312 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_864
timestamp 1598351757
transform -1 0 264 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_684
timestamp 1598351757
transform 1 0 184 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_367
timestamp 1598351757
transform 1 0 8 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_857
timestamp 1598351757
transform 1 0 136 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_365
timestamp 1598351757
transform -1 0 136 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_299
timestamp 1598351757
transform -1 0 88 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_565
timestamp 1598351757
transform -1 0 4264 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_439
timestamp 1598351757
transform -1 0 4216 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_385
timestamp 1598351757
transform -1 0 4184 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_416
timestamp 1598351757
transform -1 0 4120 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_631
timestamp 1598351757
transform 1 0 4024 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_438
timestamp 1598351757
transform 1 0 4120 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_489
timestamp 1598351757
transform -1 0 4024 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_476
timestamp 1598351757
transform -1 0 3960 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_632
timestamp 1598351757
transform 1 0 3832 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_378
timestamp 1598351757
transform -1 0 3992 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_379
timestamp 1598351757
transform 1 0 3880 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_462
timestamp 1598351757
transform -1 0 3832 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_296
timestamp 1598351757
transform -1 0 3752 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_246
timestamp 1598351757
transform -1 0 3784 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_404
timestamp 1598351757
transform 1 0 3672 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_269
timestamp 1598351757
transform -1 0 3576 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_247
timestamp 1598351757
transform 1 0 3640 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_490
timestamp 1598351757
transform -1 0 3640 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_435
timestamp 1598351757
transform 1 0 3576 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_264
timestamp 1598351757
transform -1 0 3464 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_231
timestamp 1598351757
transform 1 0 3496 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_225
timestamp 1598351757
transform -1 0 3496 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_226
timestamp 1598351757
transform 1 0 3384 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_528
timestamp 1598351757
transform 1 0 3336 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_473
timestamp 1598351757
transform 1 0 3256 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_312
timestamp 1598351757
transform -1 0 3336 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_620
timestamp 1598351757
transform -1 0 3256 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_613
timestamp 1598351757
transform 1 0 3160 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_361
timestamp 1598351757
transform 1 0 3080 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_681
timestamp 1598351757
transform 1 0 3128 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_382
timestamp 1598351757
transform 1 0 2968 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_362
timestamp 1598351757
transform 1 0 2920 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_295
timestamp 1598351757
transform -1 0 3080 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_230
timestamp 1598351757
transform 1 0 3016 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_391
timestamp 1598351757
transform -1 0 2920 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_717
timestamp 1598351757
transform -1 0 2840 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_120
timestamp 1598351757
transform -1 0 2872 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_558
timestamp 1598351757
transform 1 0 2744 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_218
timestamp 1598351757
transform 1 0 2664 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_390
timestamp 1598351757
transform 1 0 2712 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_192
timestamp 1598351757
transform 1 0 2632 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_216
timestamp 1598351757
transform 1 0 2584 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_538
timestamp 1598351757
transform -1 0 2552 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_311
timestamp 1598351757
transform -1 0 2504 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_411
timestamp 1598351757
transform 1 0 2552 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_336
timestamp 1598351757
transform -1 0 2424 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_312
timestamp 1598351757
transform -1 0 2344 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_75
timestamp 1598351757
transform 1 0 2424 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_361
timestamp 1598351757
transform 1 0 2344 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_543
timestamp 1598351757
transform 1 0 2216 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_176
timestamp 1598351757
transform -1 0 2216 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_417
timestamp 1598351757
transform 1 0 2264 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_370
timestamp 1598351757
transform 1 0 2120 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_388
timestamp 1598351757
transform 1 0 2072 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_180
timestamp 1598351757
transform -1 0 2072 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_158
timestamp 1598351757
transform -1 0 2024 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_182
timestamp 1598351757
transform -1 0 1992 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_775
timestamp 1598351757
transform 1 0 1896 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_560
timestamp 1598351757
transform -1 0 1896 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_166
timestamp 1598351757
transform -1 0 1832 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_169
timestamp 1598351757
transform -1 0 1784 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_301
timestamp 1598351757
transform -1 0 1736 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_625
timestamp 1598351757
transform -1 0 1864 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_353
timestamp 1598351757
transform 1 0 1576 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_248
timestamp 1598351757
transform -1 0 1688 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_353
timestamp 1598351757
transform 1 0 1624 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_440
timestamp 1598351757
transform 1 0 1544 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_566
timestamp 1598351757
transform 1 0 1496 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_716
timestamp 1598351757
transform -1 0 1496 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_559
timestamp 1598351757
transform -1 0 1448 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_303
timestamp 1598351757
transform -1 0 1416 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_723
timestamp 1598351757
transform -1 0 1336 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_250
timestamp 1598351757
transform 1 0 1336 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_260
timestamp 1598351757
transform -1 0 1288 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_327
timestamp 1598351757
transform -1 0 1256 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_806
timestamp 1598351757
transform -1 0 1144 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_188
timestamp 1598351757
transform 1 0 1176 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_259
timestamp 1598351757
transform -1 0 1176 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_405
timestamp 1598351757
transform -1 0 1064 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_406
timestamp 1598351757
transform 1 0 968 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_329
timestamp 1598351757
transform -1 0 1096 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_577
timestamp 1598351757
transform -1 0 968 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_175
timestamp 1598351757
transform -1 0 936 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_174
timestamp 1598351757
transform -1 0 856 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_156
timestamp 1598351757
transform 1 0 856 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_457
timestamp 1598351757
transform -1 0 808 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_590
timestamp 1598351757
transform -1 0 776 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_737
timestamp 1598351757
transform 1 0 616 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_458
timestamp 1598351757
transform 1 0 696 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_580
timestamp 1598351757
transform 1 0 664 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_722
timestamp 1598351757
transform -1 0 584 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_576
timestamp 1598351757
transform 1 0 584 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_562
timestamp 1598351757
transform 1 0 504 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_666
timestamp 1598351757
transform -1 0 504 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_811
timestamp 1598351757
transform -1 0 392 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_526
timestamp 1598351757
transform 1 0 424 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_637
timestamp 1598351757
transform -1 0 424 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_340
timestamp 1598351757
transform 1 0 312 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_863
timestamp 1598351757
transform -1 0 216 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_454
timestamp 1598351757
transform -1 0 312 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_641
timestamp 1598351757
transform -1 0 280 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_685
timestamp 1598351757
transform -1 0 248 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_812
timestamp 1598351757
transform -1 0 56 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_810
timestamp 1598351757
transform -1 0 136 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_678
timestamp 1598351757
transform 1 0 136 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_640
timestamp 1598351757
transform -1 0 88 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_560
timestamp 1598351757
transform 1 0 4216 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_576
timestamp 1598351757
transform 1 0 4136 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_433
timestamp 1598351757
transform 1 0 4184 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_559
timestamp 1598351757
transform 1 0 4056 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_642
timestamp 1598351757
transform 1 0 3976 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_424
timestamp 1598351757
transform 1 0 4104 0 1 1410
box -18 -6 52 210
use INVX1  INVX1_405
timestamp 1598351757
transform 1 0 4024 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_517
timestamp 1598351757
transform 1 0 3928 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_271
timestamp 1598351757
transform -1 0 3928 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_276
timestamp 1598351757
transform -1 0 3880 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_518
timestamp 1598351757
transform 1 0 3752 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_520
timestamp 1598351757
transform -1 0 3752 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_235
timestamp 1598351757
transform -1 0 3832 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_519
timestamp 1598351757
transform 1 0 3656 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_368
timestamp 1598351757
transform 1 0 3608 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_547
timestamp 1598351757
transform -1 0 3576 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_446
timestamp 1598351757
transform 1 0 3576 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_573
timestamp 1598351757
transform -1 0 3528 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_735
timestamp 1598351757
transform -1 0 3480 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_658
timestamp 1598351757
transform 1 0 3384 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_572
timestamp 1598351757
transform 1 0 3304 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_861
timestamp 1598351757
transform -1 0 3304 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_159
timestamp 1598351757
transform -1 0 3384 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_458
timestamp 1598351757
transform -1 0 3256 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_10
timestamp 1598351757
transform 1 0 3128 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_17
timestamp 1598351757
transform 1 0 3176 0 1 1410
box -18 -6 52 210
use INVX1  INVX1_426
timestamp 1598351757
transform 1 0 3096 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_564
timestamp 1598351757
transform 1 0 3048 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_552
timestamp 1598351757
transform -1 0 2984 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_425
timestamp 1598351757
transform 1 0 3016 0 1 1410
box -18 -6 52 210
use INVX1  INVX1_416
timestamp 1598351757
transform 1 0 2984 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_129
timestamp 1598351757
transform 1 0 2856 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_542
timestamp 1598351757
transform -1 0 2856 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_102
timestamp 1598351757
transform 1 0 2760 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_304
timestamp 1598351757
transform 1 0 2904 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_539
timestamp 1598351757
transform -1 0 2728 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_143
timestamp 1598351757
transform 1 0 2600 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_193
timestamp 1598351757
transform -1 0 2760 0 1 1410
box -18 -6 52 210
use INVX1  INVX1_129
timestamp 1598351757
transform 1 0 2648 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_551
timestamp 1598351757
transform 1 0 2552 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_99
timestamp 1598351757
transform -1 0 2552 0 1 1410
box -18 -6 52 210
use INVX1  INVX1_130
timestamp 1598351757
transform 1 0 2488 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_524
timestamp 1598351757
transform 1 0 2440 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_319
timestamp 1598351757
transform -1 0 2440 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_703
timestamp 1598351757
transform 1 0 2344 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_419
timestamp 1598351757
transform 1 0 2312 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_545
timestamp 1598351757
transform 1 0 2264 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_150
timestamp 1598351757
transform -1 0 2264 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_65
timestamp 1598351757
transform 1 0 2184 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_441
timestamp 1598351757
transform 1 0 2136 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_442
timestamp 1598351757
transform -1 0 2136 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_177
timestamp 1598351757
transform -1 0 2088 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_444
timestamp 1598351757
transform -1 0 2040 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_443
timestamp 1598351757
transform 1 0 1912 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_167
timestamp 1598351757
transform -1 0 1912 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_349
timestamp 1598351757
transform 1 0 1960 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_46
timestamp 1598351757
transform 1 0 1816 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_568
timestamp 1598351757
transform 1 0 1704 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_52
timestamp 1598351757
transform 1 0 1784 0 1 1410
box -18 -6 52 210
use INVX1  INVX1_441
timestamp 1598351757
transform -1 0 1784 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_454
timestamp 1598351757
transform -1 0 1704 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_604
timestamp 1598351757
transform 1 0 1576 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_116
timestamp 1598351757
transform 1 0 1624 0 1 1410
box -18 -6 52 210
use INVX1  INVX1_115
timestamp 1598351757
transform 1 0 1544 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_124
timestamp 1598351757
transform 1 0 1496 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_298
timestamp 1598351757
transform -1 0 1464 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_197
timestamp 1598351757
transform 1 0 1464 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_302
timestamp 1598351757
transform -1 0 1416 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_674
timestamp 1598351757
transform -1 0 1304 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_578
timestamp 1598351757
transform -1 0 1368 0 1 1410
box -18 -6 52 210
use INVX1  INVX1_249
timestamp 1598351757
transform 1 0 1304 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_675
timestamp 1598351757
transform -1 0 1256 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_736
timestamp 1598351757
transform 1 0 1096 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_532
timestamp 1598351757
transform 1 0 1176 0 1 1410
box -18 -6 52 210
use INVX1  INVX1_533
timestamp 1598351757
transform -1 0 1176 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_448
timestamp 1598351757
transform 1 0 1048 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_421
timestamp 1598351757
transform -1 0 1048 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_628
timestamp 1598351757
transform -1 0 1000 0 1 1410
box -18 -6 52 210
use INVX1  INVX1_629
timestamp 1598351757
transform -1 0 968 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_802
timestamp 1598351757
transform -1 0 936 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_591
timestamp 1598351757
transform -1 0 856 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_579
timestamp 1598351757
transform -1 0 888 0 1 1410
box -18 -6 52 210
use INVX1  INVX1_561
timestamp 1598351757
transform -1 0 808 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_585
timestamp 1598351757
transform -1 0 776 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_741
timestamp 1598351757
transform -1 0 728 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_637
timestamp 1598351757
transform -1 0 680 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_122
timestamp 1598351757
transform 1 0 584 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_121
timestamp 1598351757
transform -1 0 584 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_497
timestamp 1598351757
transform -1 0 536 0 1 1410
box -18 -6 52 210
use INVX1  INVX1_111
timestamp 1598351757
transform -1 0 504 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_638
timestamp 1598351757
transform 1 0 424 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_866
timestamp 1598351757
transform 1 0 312 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_638
timestamp 1598351757
transform -1 0 424 0 1 1410
box -18 -6 52 210
use INVX1  INVX1_686
timestamp 1598351757
transform -1 0 392 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_582
timestamp 1598351757
transform -1 0 312 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_632
timestamp 1598351757
transform -1 0 264 0 1 1410
box -18 -6 52 210
use INVX1  INVX1_263
timestamp 1598351757
transform -1 0 232 0 1 1410
box -18 -6 52 210
use INVX1  INVX1_290
timestamp 1598351757
transform -1 0 200 0 1 1410
box -18 -6 52 210
use INVX1  INVX1_631
timestamp 1598351757
transform 1 0 8 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_329
timestamp 1598351757
transform -1 0 168 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_809
timestamp 1598351757
transform 1 0 40 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_639
timestamp 1598351757
transform -1 0 120 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_578
timestamp 1598351757
transform 1 0 4152 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_451
timestamp 1598351757
transform 1 0 4200 0 -1 1410
box -18 -6 52 210
use FILL  FILL_7_2
timestamp 1598351757
transform -1 0 4264 0 -1 1410
box -16 -6 32 210
use FILL  FILL_7_1
timestamp 1598351757
transform -1 0 4248 0 -1 1410
box -16 -6 32 210
use NAND2X1  NAND2X1_579
timestamp 1598351757
transform 1 0 4008 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_219
timestamp 1598351757
transform 1 0 4120 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_453
timestamp 1598351757
transform 1 0 4088 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_450
timestamp 1598351757
transform -1 0 4088 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_295
timestamp 1598351757
transform 1 0 3960 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_550
timestamp 1598351757
transform 1 0 3912 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_346
timestamp 1598351757
transform 1 0 3832 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_421
timestamp 1598351757
transform 1 0 3880 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_292
timestamp 1598351757
transform -1 0 3832 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_270
timestamp 1598351757
transform 1 0 3704 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_233
timestamp 1598351757
transform 1 0 3752 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_232
timestamp 1598351757
transform 1 0 3672 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_275
timestamp 1598351757
transform 1 0 3624 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_527
timestamp 1598351757
transform -1 0 3624 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_234
timestamp 1598351757
transform 1 0 3544 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_110
timestamp 1598351757
transform -1 0 3512 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_181
timestamp 1598351757
transform -1 0 3432 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_104
timestamp 1598351757
transform -1 0 3544 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_103
timestamp 1598351757
transform -1 0 3464 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_179
timestamp 1598351757
transform -1 0 3320 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_502
timestamp 1598351757
transform -1 0 3384 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_447
timestamp 1598351757
transform -1 0 3352 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_682
timestamp 1598351757
transform -1 0 3272 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_457
timestamp 1598351757
transform -1 0 3208 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_464
timestamp 1598351757
transform 1 0 3080 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_364
timestamp 1598351757
transform -1 0 3240 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_363
timestamp 1598351757
transform -1 0 3160 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_865
timestamp 1598351757
transform -1 0 3048 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_370
timestamp 1598351757
transform -1 0 3080 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_442
timestamp 1598351757
transform 1 0 2968 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_301
timestamp 1598351757
transform 1 0 2936 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_111
timestamp 1598351757
transform 1 0 2888 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_217
timestamp 1598351757
transform -1 0 2856 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_323
timestamp 1598351757
transform 1 0 2760 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_119
timestamp 1598351757
transform -1 0 2888 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_112
timestamp 1598351757
transform -1 0 2760 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_332
timestamp 1598351757
transform -1 0 2712 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_374
timestamp 1598351757
transform 1 0 2616 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_325
timestamp 1598351757
transform 1 0 2568 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_322
timestamp 1598351757
transform -1 0 2536 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_418
timestamp 1598351757
transform 1 0 2536 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_544
timestamp 1598351757
transform -1 0 2488 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_373
timestamp 1598351757
transform -1 0 2440 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_545
timestamp 1598351757
transform 1 0 2360 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_412
timestamp 1598351757
transform -1 0 2360 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_109
timestamp 1598351757
transform 1 0 2280 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_257
timestamp 1598351757
transform -1 0 2280 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_134
timestamp 1598351757
transform 1 0 2216 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_67
timestamp 1598351757
transform -1 0 2216 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_438
timestamp 1598351757
transform -1 0 2184 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_62
timestamp 1598351757
transform 1 0 2088 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_439
timestamp 1598351757
transform -1 0 2056 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_66
timestamp 1598351757
transform 1 0 2056 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_804
timestamp 1598351757
transform -1 0 1976 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_369
timestamp 1598351757
transform -1 0 1896 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_350
timestamp 1598351757
transform -1 0 2008 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_634
timestamp 1598351757
transform -1 0 1928 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_567
timestamp 1598351757
transform -1 0 1816 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_603
timestamp 1598351757
transform 1 0 1688 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_51
timestamp 1598351757
transform -1 0 1848 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_255
timestamp 1598351757
transform -1 0 1768 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_605
timestamp 1598351757
transform -1 0 1688 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_469
timestamp 1598351757
transform -1 0 1640 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_360
timestamp 1598351757
transform -1 0 1608 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_347
timestamp 1598351757
transform -1 0 1576 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_299
timestamp 1598351757
transform 1 0 1496 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_808
timestamp 1598351757
transform 1 0 1448 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_123
timestamp 1598351757
transform 1 0 1400 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_854
timestamp 1598351757
transform 1 0 1352 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_354
timestamp 1598351757
transform -1 0 1352 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_466
timestamp 1598351757
transform 1 0 1256 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_359
timestamp 1598351757
transform 1 0 1224 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_453
timestamp 1598351757
transform 1 0 1144 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_372
timestamp 1598351757
transform -1 0 1224 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_354
timestamp 1598351757
transform 1 0 1112 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_173
timestamp 1598351757
transform -1 0 1112 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_799
timestamp 1598351757
transform -1 0 1064 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_798
timestamp 1598351757
transform -1 0 1016 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_460
timestamp 1598351757
transform 1 0 936 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_593
timestamp 1598351757
transform 1 0 888 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_718
timestamp 1598351757
transform -1 0 888 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_172
timestamp 1598351757
transform -1 0 840 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_434
timestamp 1598351757
transform -1 0 760 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_431
timestamp 1598351757
transform -1 0 712 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_586
timestamp 1598351757
transform -1 0 664 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_344
timestamp 1598351757
transform 1 0 760 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_120
timestamp 1598351757
transform -1 0 552 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_112
timestamp 1598351757
transform -1 0 616 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_114
timestamp 1598351757
transform 1 0 552 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_113
timestamp 1598351757
transform 1 0 472 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_288
timestamp 1598351757
transform -1 0 472 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_462
timestamp 1598351757
transform -1 0 440 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_594
timestamp 1598351757
transform -1 0 408 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_675
timestamp 1598351757
transform -1 0 376 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_856
timestamp 1598351757
transform -1 0 344 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_761
timestamp 1598351757
transform -1 0 264 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_356
timestamp 1598351757
transform -1 0 216 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_677
timestamp 1598351757
transform -1 0 296 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_801
timestamp 1598351757
transform -1 0 56 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_355
timestamp 1598351757
transform -1 0 136 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_289
timestamp 1598351757
transform 1 0 136 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_593
timestamp 1598351757
transform -1 0 88 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_444
timestamp 1598351757
transform 1 0 4232 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_481
timestamp 1598351757
transform 1 0 4184 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_384
timestamp 1598351757
transform 1 0 4152 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_256
timestamp 1598351757
transform -1 0 4152 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_218
timestamp 1598351757
transform 1 0 4072 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_415
timestamp 1598351757
transform -1 0 4072 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_449
timestamp 1598351757
transform 1 0 4008 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_255
timestamp 1598351757
transform 1 0 3960 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_541
timestamp 1598351757
transform -1 0 3960 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_522
timestamp 1598351757
transform 1 0 3864 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_272
timestamp 1598351757
transform 1 0 3816 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_274
timestamp 1598351757
transform 1 0 3704 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_406
timestamp 1598351757
transform -1 0 3816 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_420
timestamp 1598351757
transform -1 0 3784 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_844
timestamp 1598351757
transform 1 0 3656 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_497
timestamp 1598351757
transform -1 0 3656 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_184
timestamp 1598351757
transform -1 0 3608 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_665
timestamp 1598351757
transform -1 0 3560 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_45
timestamp 1598351757
transform -1 0 3528 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_178
timestamp 1598351757
transform 1 0 3400 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_392
timestamp 1598351757
transform -1 0 3480 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_393
timestamp 1598351757
transform 1 0 3368 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_501
timestamp 1598351757
transform 1 0 3320 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_575
timestamp 1598351757
transform -1 0 3288 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_303
timestamp 1598351757
transform 1 0 3288 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_649
timestamp 1598351757
transform -1 0 3176 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_643
timestamp 1598351757
transform 1 0 3080 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_448
timestamp 1598351757
transform 1 0 3208 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_617
timestamp 1598351757
transform -1 0 3208 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_471
timestamp 1598351757
transform -1 0 3048 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_849
timestamp 1598351757
transform -1 0 3000 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_503
timestamp 1598351757
transform -1 0 3080 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_371
timestamp 1598351757
transform 1 0 2920 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_478
timestamp 1598351757
transform 1 0 2840 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_377
timestamp 1598351757
transform -1 0 2920 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_128
timestamp 1598351757
transform -1 0 2840 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_383
timestamp 1598351757
transform 1 0 2776 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_477
timestamp 1598351757
transform 1 0 2728 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_574
timestamp 1598351757
transform 1 0 2680 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_657
timestamp 1598351757
transform 1 0 2600 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_375
timestamp 1598351757
transform 1 0 2648 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_600
timestamp 1598351757
transform -1 0 2568 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_602
timestamp 1598351757
transform -1 0 2520 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_242
timestamp 1598351757
transform -1 0 2600 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_700
timestamp 1598351757
transform -1 0 2472 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_601
timestamp 1598351757
transform 1 0 2376 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_253
timestamp 1598351757
transform 1 0 2344 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_468
timestamp 1598351757
transform -1 0 2344 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_714
timestamp 1598351757
transform -1 0 2312 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_794
timestamp 1598351757
transform -1 0 2232 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_546
timestamp 1598351757
transform 1 0 2232 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_624
timestamp 1598351757
transform -1 0 2184 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_788
timestamp 1598351757
transform 1 0 2040 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_727
timestamp 1598351757
transform -1 0 2040 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_618
timestamp 1598351757
transform 1 0 2120 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_252
timestamp 1598351757
transform -1 0 2120 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_469
timestamp 1598351757
transform -1 0 1992 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_535
timestamp 1598351757
transform -1 0 1912 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_352
timestamp 1598351757
transform -1 0 1944 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_534
timestamp 1598351757
transform -1 0 1864 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_831
timestamp 1598351757
transform -1 0 1752 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_374
timestamp 1598351757
transform 1 0 1784 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_409
timestamp 1598351757
transform -1 0 1784 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_648
timestamp 1598351757
transform 1 0 1656 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_300
timestamp 1598351757
transform -1 0 1656 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_645
timestamp 1598351757
transform 1 0 1528 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_506
timestamp 1598351757
transform 1 0 1576 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_321
timestamp 1598351757
transform -1 0 1496 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_324
timestamp 1598351757
transform -1 0 1448 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_376
timestamp 1598351757
transform 1 0 1496 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_326
timestamp 1598351757
transform -1 0 1368 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_256
timestamp 1598351757
transform -1 0 1400 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_258
timestamp 1598351757
transform -1 0 1320 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_504
timestamp 1598351757
transform 1 0 1256 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_118
timestamp 1598351757
transform 1 0 1208 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_437
timestamp 1598351757
transform -1 0 1144 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_345
timestamp 1598351757
transform -1 0 1208 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_355
timestamp 1598351757
transform 1 0 1144 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_440
timestamp 1598351757
transform -1 0 1096 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_468
timestamp 1598351757
transform 1 0 936 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_348
timestamp 1598351757
transform -1 0 1048 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_459
timestamp 1598351757
transform -1 0 1016 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_652
timestamp 1598351757
transform -1 0 904 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_436
timestamp 1598351757
transform 1 0 808 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_346
timestamp 1598351757
transform 1 0 904 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_588
timestamp 1598351757
transform -1 0 808 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_683
timestamp 1598351757
transform 1 0 728 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_644
timestamp 1598351757
transform 1 0 680 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_597
timestamp 1598351757
transform -1 0 680 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_694
timestamp 1598351757
transform 1 0 552 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_596
timestamp 1598351757
transform -1 0 552 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_461
timestamp 1598351757
transform -1 0 632 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_426
timestamp 1598351757
transform -1 0 504 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_450
timestamp 1598351757
transform -1 0 456 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_428
timestamp 1598351757
transform -1 0 376 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_505
timestamp 1598351757
transform 1 0 376 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_635
timestamp 1598351757
transform -1 0 328 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_451
timestamp 1598351757
transform -1 0 280 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_466
timestamp 1598351757
transform 1 0 200 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_264
timestamp 1598351757
transform -1 0 200 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_630
timestamp 1598351757
transform -1 0 40 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_330
timestamp 1598351757
transform -1 0 168 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_760
timestamp 1598351757
transform -1 0 88 0 1 1010
box -16 -6 64 210
use INVX1  INVX1_265
timestamp 1598351757
transform 1 0 88 0 1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_570
timestamp 1598351757
transform -1 0 4232 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_437
timestamp 1598351757
transform 1 0 4152 0 -1 1010
box -18 -6 52 210
use FILL  FILL_5_2
timestamp 1598351757
transform -1 0 4264 0 -1 1010
box -16 -6 32 210
use FILL  FILL_5_1
timestamp 1598351757
transform -1 0 4248 0 -1 1010
box -16 -6 32 210
use NAND2X1  NAND2X1_556
timestamp 1598351757
transform -1 0 4120 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_563
timestamp 1598351757
transform -1 0 4072 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_430
timestamp 1598351757
transform 1 0 4120 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_427
timestamp 1598351757
transform 1 0 3992 0 -1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_553
timestamp 1598351757
transform 1 0 3912 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_456
timestamp 1598351757
transform 1 0 3864 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_414
timestamp 1598351757
transform -1 0 3992 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_362
timestamp 1598351757
transform -1 0 3864 0 -1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_523
timestamp 1598351757
transform 1 0 3784 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_526
timestamp 1598351757
transform -1 0 3784 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_546
timestamp 1598351757
transform 1 0 3688 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_500
timestamp 1598351757
transform -1 0 3688 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_521
timestamp 1598351757
transform -1 0 3640 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_413
timestamp 1598351757
transform 1 0 3560 0 -1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_525
timestamp 1598351757
transform 1 0 3512 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_540
timestamp 1598351757
transform 1 0 3464 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_183
timestamp 1598351757
transform -1 0 3464 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_190
timestamp 1598351757
transform -1 0 3416 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_372
timestamp 1598351757
transform -1 0 3368 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_371
timestamp 1598351757
transform 1 0 3240 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_302
timestamp 1598351757
transform 1 0 3288 0 -1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_595
timestamp 1598351757
transform 1 0 3192 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_787
timestamp 1598351757
transform 1 0 3144 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_249
timestamp 1598351757
transform -1 0 3112 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_215
timestamp 1598351757
transform -1 0 3144 0 -1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_465
timestamp 1598351757
transform 1 0 2984 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_131
timestamp 1598351757
transform -1 0 2984 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_216
timestamp 1598351757
transform 1 0 3032 0 -1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_140
timestamp 1598351757
transform -1 0 2904 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_105
timestamp 1598351757
transform 1 0 2904 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_519
timestamp 1598351757
transform 1 0 2824 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_127
timestamp 1598351757
transform -1 0 2824 0 -1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_141
timestamp 1598351757
transform 1 0 2744 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_130
timestamp 1598351757
transform 1 0 2664 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_701
timestamp 1598351757
transform 1 0 2616 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_122
timestamp 1598351757
transform -1 0 2744 0 -1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_710
timestamp 1598351757
transform 1 0 2472 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_510
timestamp 1598351757
transform -1 0 2616 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_670
timestamp 1598351757
transform -1 0 2584 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_553
timestamp 1598351757
transform 1 0 2520 0 -1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_314
timestamp 1598351757
transform 1 0 2392 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_307
timestamp 1598351757
transform 1 0 2344 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_317
timestamp 1598351757
transform 1 0 2296 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_121
timestamp 1598351757
transform 1 0 2440 0 -1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_704
timestamp 1598351757
transform -1 0 2232 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_557
timestamp 1598351757
transform -1 0 2296 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_251
timestamp 1598351757
transform -1 0 2264 0 -1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_313
timestamp 1598351757
transform 1 0 2136 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_308
timestamp 1598351757
transform 1 0 2088 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_446
timestamp 1598351757
transform -1 0 2088 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_306
timestamp 1598351757
transform 1 0 1992 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_418
timestamp 1598351757
transform 1 0 1944 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_533
timestamp 1598351757
transform 1 0 1896 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_655
timestamp 1598351757
transform 1 0 1848 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_273
timestamp 1598351757
transform 1 0 1736 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_119
timestamp 1598351757
transform 1 0 1688 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_509
timestamp 1598351757
transform 1 0 1816 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_652
timestamp 1598351757
transform 1 0 1784 0 -1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_498
timestamp 1598351757
transform 1 0 1608 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_188
timestamp 1598351757
transform 1 0 1560 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_110
timestamp 1598351757
transform -1 0 1688 0 -1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_433
timestamp 1598351757
transform -1 0 1560 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_320
timestamp 1598351757
transform 1 0 1432 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_165
timestamp 1598351757
transform 1 0 1480 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_653
timestamp 1598351757
transform 1 0 1400 0 -1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_832
timestamp 1598351757
transform 1 0 1320 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_423
timestamp 1598351757
transform -1 0 1320 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_435
timestamp 1598351757
transform 1 0 1224 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_166
timestamp 1598351757
transform -1 0 1400 0 -1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_432
timestamp 1598351757
transform -1 0 1224 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_449
timestamp 1598351757
transform 1 0 1128 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_424
timestamp 1598351757
transform 1 0 1080 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_592
timestamp 1598351757
transform -1 0 1080 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_589
timestamp 1598351757
transform 1 0 984 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_470
timestamp 1598351757
transform -1 0 984 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_695
timestamp 1598351757
transform 1 0 824 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_598
timestamp 1598351757
transform -1 0 824 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_141
timestamp 1598351757
transform 1 0 904 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_464
timestamp 1598351757
transform -1 0 904 0 -1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_686
timestamp 1598351757
transform -1 0 776 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_684
timestamp 1598351757
transform 1 0 680 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_465
timestamp 1598351757
transform 1 0 648 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_584
timestamp 1598351757
transform 1 0 616 0 -1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_688
timestamp 1598351757
transform 1 0 536 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_540
timestamp 1598351757
transform 1 0 584 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_539
timestamp 1598351757
transform 1 0 504 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_513
timestamp 1598351757
transform -1 0 504 0 -1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_427
timestamp 1598351757
transform -1 0 440 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_463
timestamp 1598351757
transform -1 0 472 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_358
timestamp 1598351757
transform 1 0 360 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_356
timestamp 1598351757
transform -1 0 360 0 -1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_452
timestamp 1598351757
transform -1 0 328 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_599
timestamp 1598351757
transform -1 0 248 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_357
timestamp 1598351757
transform 1 0 248 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_467
timestamp 1598351757
transform -1 0 200 0 -1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_800
timestamp 1598351757
transform 1 0 8 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_331
timestamp 1598351757
transform 1 0 56 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_537
timestamp 1598351757
transform -1 0 168 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_495
timestamp 1598351757
transform -1 0 136 0 -1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_562
timestamp 1598351757
transform 1 0 4152 0 1 610
box -16 -6 64 210
use INVX1  INVX1_436
timestamp 1598351757
transform 1 0 4200 0 1 610
box -18 -6 52 210
use FILL  FILL_4_2
timestamp 1598351757
transform 1 0 4248 0 1 610
box -16 -6 32 210
use FILL  FILL_4_1
timestamp 1598351757
transform 1 0 4232 0 1 610
box -16 -6 32 210
use NAND2X1  NAND2X1_555
timestamp 1598351757
transform -1 0 4152 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_344
timestamp 1598351757
transform 1 0 3992 0 1 610
box -16 -6 64 210
use INVX1  INVX1_429
timestamp 1598351757
transform 1 0 4072 0 1 610
box -18 -6 52 210
use INVX1  INVX1_386
timestamp 1598351757
transform 1 0 4040 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_482
timestamp 1598351757
transform 1 0 3912 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_484
timestamp 1598351757
transform 1 0 3832 0 1 610
box -16 -6 64 210
use INVX1  INVX1_217
timestamp 1598351757
transform -1 0 3992 0 1 610
box -18 -6 52 210
use INVX1  INVX1_428
timestamp 1598351757
transform 1 0 3880 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_257
timestamp 1598351757
transform 1 0 3784 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_486
timestamp 1598351757
transform -1 0 3784 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_705
timestamp 1598351757
transform 1 0 3688 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_485
timestamp 1598351757
transform 1 0 3576 0 1 610
box -16 -6 64 210
use INVX1  INVX1_387
timestamp 1598351757
transform -1 0 3688 0 1 610
box -18 -6 52 210
use INVX1  INVX1_391
timestamp 1598351757
transform 1 0 3624 0 1 610
box -18 -6 52 210
use INVX1  INVX1_367
timestamp 1598351757
transform 1 0 3544 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_496
timestamp 1598351757
transform 1 0 3464 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_693
timestamp 1598351757
transform 1 0 3416 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_554
timestamp 1598351757
transform 1 0 3368 0 1 610
box -16 -6 64 210
use INVX1  INVX1_608
timestamp 1598351757
transform 1 0 3512 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_706
timestamp 1598351757
transform 1 0 3320 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_692
timestamp 1598351757
transform -1 0 3320 0 1 610
box -16 -6 64 210
use INVX1  INVX1_118
timestamp 1598351757
transform -1 0 3272 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_115
timestamp 1598351757
transform 1 0 3192 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_702
timestamp 1598351757
transform -1 0 3160 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_862
timestamp 1598351757
transform -1 0 3112 0 1 610
box -16 -6 64 210
use INVX1  INVX1_109
timestamp 1598351757
transform -1 0 3192 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_859
timestamp 1598351757
transform 1 0 2952 0 1 610
box -16 -6 64 210
use INVX1  INVX1_683
timestamp 1598351757
transform -1 0 3064 0 1 610
box -18 -6 52 210
use INVX1  INVX1_680
timestamp 1598351757
transform 1 0 3000 0 1 610
box -18 -6 52 210
use INVX1  INVX1_544
timestamp 1598351757
transform -1 0 2952 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_715
timestamp 1598351757
transform -1 0 2920 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_225
timestamp 1598351757
transform -1 0 2808 0 1 610
box -16 -6 64 210
use INVX1  INVX1_126
timestamp 1598351757
transform -1 0 2872 0 1 610
box -18 -6 52 210
use INVX1  INVX1_200
timestamp 1598351757
transform -1 0 2840 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_280
timestamp 1598351757
transform -1 0 2728 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_659
timestamp 1598351757
transform 1 0 2600 0 1 610
box -16 -6 64 210
use INVX1  INVX1_199
timestamp 1598351757
transform -1 0 2760 0 1 610
box -18 -6 52 210
use INVX1  INVX1_518
timestamp 1598351757
transform -1 0 2680 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_136
timestamp 1598351757
transform -1 0 2568 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_711
timestamp 1598351757
transform -1 0 2520 0 1 610
box -16 -6 64 210
use INVX1  INVX1_402
timestamp 1598351757
transform -1 0 2600 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_461
timestamp 1598351757
transform 1 0 2424 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_411
timestamp 1598351757
transform 1 0 2376 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_516
timestamp 1598351757
transform 1 0 2328 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_515
timestamp 1598351757
transform 1 0 2280 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_724
timestamp 1598351757
transform -1 0 2248 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_417
timestamp 1598351757
transform -1 0 2200 0 1 610
box -16 -6 64 210
use INVX1  INVX1_558
timestamp 1598351757
transform -1 0 2280 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_413
timestamp 1598351757
transform -1 0 2152 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_77
timestamp 1598351757
transform -1 0 2104 0 1 610
box -16 -6 64 210
use INVX1  INVX1_61
timestamp 1598351757
transform 1 0 2024 0 1 610
box -18 -6 52 210
use INVX1  INVX1_78
timestamp 1598351757
transform -1 0 2024 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_54
timestamp 1598351757
transform -1 0 1992 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_512
timestamp 1598351757
transform 1 0 1896 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_513
timestamp 1598351757
transform 1 0 1848 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_841
timestamp 1598351757
transform -1 0 1816 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_15
timestamp 1598351757
transform -1 0 1768 0 1 610
box -16 -6 64 210
use INVX1  INVX1_401
timestamp 1598351757
transform -1 0 1848 0 1 610
box -18 -6 52 210
use INVX1  INVX1_24
timestamp 1598351757
transform -1 0 1720 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_511
timestamp 1598351757
transform 1 0 1608 0 1 610
box -16 -6 64 210
use INVX1  INVX1_14
timestamp 1598351757
transform 1 0 1656 0 1 610
box -18 -6 52 210
use INVX1  INVX1_338
timestamp 1598351757
transform -1 0 1608 0 1 610
box -18 -6 52 210
use INVX1  INVX1_16
timestamp 1598351757
transform -1 0 1576 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_9
timestamp 1598351757
transform 1 0 1496 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_583
timestamp 1598351757
transform 1 0 1448 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_189
timestamp 1598351757
transform 1 0 1400 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_191
timestamp 1598351757
transform 1 0 1320 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_187
timestamp 1598351757
transform -1 0 1288 0 1 610
box -16 -6 64 210
use INVX1  INVX1_15
timestamp 1598351757
transform 1 0 1368 0 1 610
box -18 -6 52 210
use INVX1  INVX1_140
timestamp 1598351757
transform -1 0 1320 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_608
timestamp 1598351757
transform -1 0 1208 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_607
timestamp 1598351757
transform -1 0 1160 0 1 610
box -16 -6 64 210
use INVX1  INVX1_472
timestamp 1598351757
transform -1 0 1240 0 1 610
box -18 -6 52 210
use INVX1  INVX1_471
timestamp 1598351757
transform -1 0 1112 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_606
timestamp 1598351757
transform 1 0 1000 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_154
timestamp 1598351757
transform -1 0 968 0 1 610
box -16 -6 64 210
use INVX1  INVX1_473
timestamp 1598351757
transform 1 0 1048 0 1 610
box -18 -6 52 210
use INVX1  INVX1_470
timestamp 1598351757
transform 1 0 968 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_707
timestamp 1598351757
transform 1 0 808 0 1 610
box -16 -6 64 210
use INVX1  INVX1_161
timestamp 1598351757
transform -1 0 920 0 1 610
box -18 -6 52 210
use INVX1  INVX1_373
timestamp 1598351757
transform 1 0 856 0 1 610
box -18 -6 52 210
use INVX1  INVX1_148
timestamp 1598351757
transform -1 0 808 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_634
timestamp 1598351757
transform 1 0 696 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_467
timestamp 1598351757
transform 1 0 616 0 1 610
box -16 -6 64 210
use INVX1  INVX1_494
timestamp 1598351757
transform -1 0 776 0 1 610
box -18 -6 52 210
use INVX1  INVX1_496
timestamp 1598351757
transform -1 0 696 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_689
timestamp 1598351757
transform -1 0 616 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_691
timestamp 1598351757
transform -1 0 568 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_690
timestamp 1598351757
transform 1 0 472 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_681
timestamp 1598351757
transform -1 0 408 0 1 610
box -16 -6 64 210
use INVX1  INVX1_541
timestamp 1598351757
transform 1 0 440 0 1 610
box -18 -6 52 210
use INVX1  INVX1_335
timestamp 1598351757
transform 1 0 408 0 1 610
box -18 -6 52 210
use INVX1  INVX1_151
timestamp 1598351757
transform -1 0 360 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_161
timestamp 1598351757
transform -1 0 328 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_685
timestamp 1598351757
transform -1 0 248 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_639
timestamp 1598351757
transform 1 0 152 0 1 610
box -16 -6 64 210
use INVX1  INVX1_152
timestamp 1598351757
transform 1 0 248 0 1 610
box -18 -6 52 210
use INVX1  INVX1_538
timestamp 1598351757
transform -1 0 40 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_687
timestamp 1598351757
transform -1 0 88 0 1 610
box -16 -6 64 210
use INVX1  INVX1_676
timestamp 1598351757
transform 1 0 120 0 1 610
box -18 -6 52 210
use INVX1  INVX1_536
timestamp 1598351757
transform -1 0 120 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_345
timestamp 1598351757
transform 1 0 4152 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_279
timestamp 1598351757
transform 1 0 4200 0 -1 610
box -18 -6 52 210
use FILL  FILL_3_2
timestamp 1598351757
transform -1 0 4264 0 -1 610
box -16 -6 32 210
use FILL  FILL_3_1
timestamp 1598351757
transform -1 0 4248 0 -1 610
box -16 -6 32 210
use NAND2X1  NAND2X1_252
timestamp 1598351757
transform -1 0 4120 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_483
timestamp 1598351757
transform -1 0 4072 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_254
timestamp 1598351757
transform -1 0 4024 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_220
timestamp 1598351757
transform 1 0 4120 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_833
timestamp 1598351757
transform -1 0 3944 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_495
timestamp 1598351757
transform -1 0 3896 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_213
timestamp 1598351757
transform -1 0 3976 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_259
timestamp 1598351757
transform 1 0 3800 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_258
timestamp 1598351757
transform 1 0 3720 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_253
timestamp 1598351757
transform -1 0 3720 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_547
timestamp 1598351757
transform -1 0 3800 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_499
timestamp 1598351757
transform -1 0 3672 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_106
timestamp 1598351757
transform 1 0 3576 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_214
timestamp 1598351757
transform -1 0 3576 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_778
timestamp 1598351757
transform -1 0 3544 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_713
timestamp 1598351757
transform -1 0 3496 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_125
timestamp 1598351757
transform -1 0 3416 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_548
timestamp 1598351757
transform 1 0 3416 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_127
timestamp 1598351757
transform -1 0 3368 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_128
timestamp 1598351757
transform -1 0 3320 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_556
timestamp 1598351757
transform -1 0 3272 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_116
timestamp 1598351757
transform 1 0 3160 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_135
timestamp 1598351757
transform -1 0 3160 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_768
timestamp 1598351757
transform -1 0 3112 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_108
timestamp 1598351757
transform -1 0 3240 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_137
timestamp 1598351757
transform 1 0 3016 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_134
timestamp 1598351757
transform 1 0 2968 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_124
timestamp 1598351757
transform -1 0 2968 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_139
timestamp 1598351757
transform -1 0 2936 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_132
timestamp 1598351757
transform 1 0 2840 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_138
timestamp 1598351757
transform -1 0 2808 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_125
timestamp 1598351757
transform 1 0 2808 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_514
timestamp 1598351757
transform -1 0 2728 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_403
timestamp 1598351757
transform -1 0 2760 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_520
timestamp 1598351757
transform -1 0 2680 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_238
timestamp 1598351757
transform 1 0 2616 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_284
timestamp 1598351757
transform 1 0 2568 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_279
timestamp 1598351757
transform 1 0 2520 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_159
timestamp 1598351757
transform -1 0 2520 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_410
timestamp 1598351757
transform -1 0 2408 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_305
timestamp 1598351757
transform -1 0 2360 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_146
timestamp 1598351757
transform -1 0 2472 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_336
timestamp 1598351757
transform -1 0 2440 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_90
timestamp 1598351757
transform -1 0 2248 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_89
timestamp 1598351757
transform 1 0 2280 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_337
timestamp 1598351757
transform -1 0 2280 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_567
timestamp 1598351757
transform -1 0 2200 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_73
timestamp 1598351757
transform -1 0 2168 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_55
timestamp 1598351757
transform -1 0 2088 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_76
timestamp 1598351757
transform -1 0 2120 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_62
timestamp 1598351757
transform -1 0 2040 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_532
timestamp 1598351757
transform -1 0 1912 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_407
timestamp 1598351757
transform 1 0 1976 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_136
timestamp 1598351757
transform 1 0 1944 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_408
timestamp 1598351757
transform 1 0 1912 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_656
timestamp 1598351757
transform -1 0 1832 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_660
timestamp 1598351757
transform -1 0 1752 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_516
timestamp 1598351757
transform -1 0 1864 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_517
timestamp 1598351757
transform -1 0 1784 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_412
timestamp 1598351757
transform -1 0 1640 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_584
timestamp 1598351757
transform -1 0 1592 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_521
timestamp 1598351757
transform -1 0 1704 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_645
timestamp 1598351757
transform 1 0 1640 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_636
timestamp 1598351757
transform -1 0 1544 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_192
timestamp 1598351757
transform -1 0 1496 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_168
timestamp 1598351757
transform -1 0 1448 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_167
timestamp 1598351757
transform 1 0 1384 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_633
timestamp 1598351757
transform 1 0 1336 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_221
timestamp 1598351757
transform -1 0 1336 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_196
timestamp 1598351757
transform 1 0 1256 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_220
timestamp 1598351757
transform 1 0 1208 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_646
timestamp 1598351757
transform 1 0 1128 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_609
timestamp 1598351757
transform -1 0 1128 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_507
timestamp 1598351757
transform 1 0 1176 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_186
timestamp 1598351757
transform -1 0 1080 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_164
timestamp 1598351757
transform 1 0 1000 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_163
timestamp 1598351757
transform -1 0 1000 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_549
timestamp 1598351757
transform 1 0 936 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_185
timestamp 1598351757
transform 1 0 888 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_162
timestamp 1598351757
transform 1 0 856 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_491
timestamp 1598351757
transform -1 0 856 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_149
timestamp 1598351757
transform -1 0 824 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_160
timestamp 1598351757
transform -1 0 760 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_640
timestamp 1598351757
transform -1 0 680 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_139
timestamp 1598351757
transform -1 0 792 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_493
timestamp 1598351757
transform -1 0 712 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_163
timestamp 1598351757
transform -1 0 600 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_162
timestamp 1598351757
transform -1 0 552 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_147
timestamp 1598351757
transform -1 0 632 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_500
timestamp 1598351757
transform -1 0 504 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_650
timestamp 1598351757
transform -1 0 440 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_501
timestamp 1598351757
transform -1 0 472 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_498
timestamp 1598351757
transform 1 0 360 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_150
timestamp 1598351757
transform 1 0 328 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_682
timestamp 1598351757
transform -1 0 328 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_651
timestamp 1598351757
transform -1 0 280 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_512
timestamp 1598351757
transform -1 0 232 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_499
timestamp 1598351757
transform 1 0 168 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_729
timestamp 1598351757
transform 1 0 8 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_855
timestamp 1598351757
transform 1 0 88 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_542
timestamp 1598351757
transform -1 0 168 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_572
timestamp 1598351757
transform 1 0 56 0 -1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_348
timestamp 1598351757
transform 1 0 4168 0 1 210
box -16 -6 64 210
use INVX1  INVX1_445
timestamp 1598351757
transform 1 0 4216 0 1 210
box -18 -6 52 210
use INVX1  INVX1_278
timestamp 1598351757
transform 1 0 4136 0 1 210
box -18 -6 52 210
use FILL  FILL_2_1
timestamp 1598351757
transform 1 0 4248 0 1 210
box -16 -6 32 210
use NAND2X1  NAND2X1_261
timestamp 1598351757
transform -1 0 4136 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_850
timestamp 1598351757
transform 1 0 4008 0 1 210
box -16 -6 64 210
use INVX1  INVX1_664
timestamp 1598351757
transform -1 0 4088 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_842
timestamp 1598351757
transform 1 0 3928 0 1 210
box -16 -6 64 210
use INVX1  INVX1_663
timestamp 1598351757
transform 1 0 3976 0 1 210
box -18 -6 52 210
use INVX1  INVX1_654
timestamp 1598351757
transform 1 0 3896 0 1 210
box -18 -6 52 210
use INVX1  INVX1_293
timestamp 1598351757
transform -1 0 3896 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_840
timestamp 1598351757
transform -1 0 3864 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_843
timestamp 1598351757
transform 1 0 3768 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_251
timestamp 1598351757
transform -1 0 3736 0 1 210
box -16 -6 64 210
use INVX1  INVX1_655
timestamp 1598351757
transform 1 0 3736 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_343
timestamp 1598351757
transform -1 0 3688 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_250
timestamp 1598351757
transform 1 0 3560 0 1 210
box -16 -6 64 210
use INVX1  INVX1_679
timestamp 1598351757
transform -1 0 3640 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_247
timestamp 1598351757
transform 1 0 3512 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_142
timestamp 1598351757
transform 1 0 3400 0 1 210
box -16 -6 64 210
use INVX1  INVX1_651
timestamp 1598351757
transform 1 0 3480 0 1 210
box -18 -6 52 210
use INVX1  INVX1_607
timestamp 1598351757
transform -1 0 3480 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_108
timestamp 1598351757
transform 1 0 3352 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_107
timestamp 1598351757
transform -1 0 3352 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_113
timestamp 1598351757
transform -1 0 3304 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_281
timestamp 1598351757
transform -1 0 3256 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_103
timestamp 1598351757
transform 1 0 3128 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_282
timestamp 1598351757
transform 1 0 3080 0 1 210
box -16 -6 64 210
use INVX1  INVX1_107
timestamp 1598351757
transform -1 0 3208 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_146
timestamp 1598351757
transform -1 0 3080 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_144
timestamp 1598351757
transform -1 0 3032 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_817
timestamp 1598351757
transform -1 0 2984 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_145
timestamp 1598351757
transform 1 0 2856 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_245
timestamp 1598351757
transform -1 0 2824 0 1 210
box -16 -6 64 210
use INVX1  INVX1_646
timestamp 1598351757
transform 1 0 2904 0 1 210
box -18 -6 52 210
use INVX1  INVX1_669
timestamp 1598351757
transform 1 0 2824 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_283
timestamp 1598351757
transform -1 0 2776 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_246
timestamp 1598351757
transform 1 0 2648 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_287
timestamp 1598351757
transform 1 0 2600 0 1 210
box -16 -6 64 210
use INVX1  INVX1_212
timestamp 1598351757
transform -1 0 2728 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_663
timestamp 1598351757
transform -1 0 2600 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_818
timestamp 1598351757
transform 1 0 2472 0 1 210
box -16 -6 64 210
use INVX1  INVX1_648
timestamp 1598351757
transform -1 0 2552 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_278
timestamp 1598351757
transform -1 0 2408 0 1 210
box -16 -6 64 210
use INVX1  INVX1_647
timestamp 1598351757
transform 1 0 2440 0 1 210
box -18 -6 52 210
use INVX1  INVX1_237
timestamp 1598351757
transform -1 0 2440 0 1 210
box -18 -6 52 210
use INVX1  INVX1_606
timestamp 1598351757
transform -1 0 2360 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_777
timestamp 1598351757
transform -1 0 2328 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_784
timestamp 1598351757
transform -1 0 2248 0 1 210
box -16 -6 64 210
use INVX1  INVX1_605
timestamp 1598351757
transform -1 0 2280 0 1 210
box -18 -6 52 210
use INVX1  INVX1_523
timestamp 1598351757
transform 1 0 2168 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_151
timestamp 1598351757
transform -1 0 2136 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_732
timestamp 1598351757
transform -1 0 2088 0 1 210
box -16 -6 64 210
use INVX1  INVX1_135
timestamp 1598351757
transform -1 0 2168 0 1 210
box -18 -6 52 210
use INVX1  INVX1_568
timestamp 1598351757
transform 1 0 2008 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_725
timestamp 1598351757
transform 1 0 1960 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_611
timestamp 1598351757
transform -1 0 1928 0 1 210
box -16 -6 64 210
use INVX1  INVX1_555
timestamp 1598351757
transform 1 0 1928 0 1 210
box -18 -6 52 210
use INVX1  INVX1_477
timestamp 1598351757
transform 1 0 1848 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_816
timestamp 1598351757
transform -1 0 1848 0 1 210
box -16 -6 64 210
use INVX1  INVX1_508
timestamp 1598351757
transform 1 0 1768 0 1 210
box -18 -6 52 210
use INVX1  INVX1_185
timestamp 1598351757
transform -1 0 1768 0 1 210
box -18 -6 52 210
use INVX1  INVX1_236
timestamp 1598351757
transform 1 0 1704 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_277
timestamp 1598351757
transform 1 0 1656 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_662
timestamp 1598351757
transform -1 0 1656 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_153
timestamp 1598351757
transform -1 0 1576 0 1 210
box -16 -6 64 210
use INVX1  INVX1_138
timestamp 1598351757
transform -1 0 1608 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_647
timestamp 1598351757
transform -1 0 1528 0 1 210
box -16 -6 64 210
use INVX1  INVX1_492
timestamp 1598351757
transform -1 0 1480 0 1 210
box -18 -6 52 210
use INVX1  INVX1_475
timestamp 1598351757
transform -1 0 1448 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_610
timestamp 1598351757
transform 1 0 1368 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_213
timestamp 1598351757
transform -1 0 1304 0 1 210
box -16 -6 64 210
use INVX1  INVX1_633
timestamp 1598351757
transform 1 0 1336 0 1 210
box -18 -6 52 210
use INVX1  INVX1_474
timestamp 1598351757
transform 1 0 1304 0 1 210
box -18 -6 52 210
use INVX1  INVX1_189
timestamp 1598351757
transform 1 0 1224 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_696
timestamp 1598351757
transform 1 0 1176 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_697
timestamp 1598351757
transform -1 0 1176 0 1 210
box -16 -6 64 210
use INVX1  INVX1_550
timestamp 1598351757
transform -1 0 1128 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_712
timestamp 1598351757
transform 1 0 1048 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_744
timestamp 1598351757
transform -1 0 1048 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_746
timestamp 1598351757
transform -1 0 1000 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_745
timestamp 1598351757
transform -1 0 952 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_781
timestamp 1598351757
transform -1 0 904 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_677
timestamp 1598351757
transform -1 0 856 0 1 210
box -16 -6 64 210
use INVX1  INVX1_186
timestamp 1598351757
transform 1 0 776 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_156
timestamp 1598351757
transform -1 0 776 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_158
timestamp 1598351757
transform -1 0 696 0 1 210
box -16 -6 64 210
use INVX1  INVX1_142
timestamp 1598351757
transform 1 0 696 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_210
timestamp 1598351757
transform -1 0 648 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_742
timestamp 1598351757
transform 1 0 552 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_594
timestamp 1598351757
transform -1 0 520 0 1 210
box -16 -6 64 210
use INVX1  INVX1_583
timestamp 1598351757
transform 1 0 520 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_653
timestamp 1598351757
transform -1 0 472 0 1 210
box -16 -6 64 210
use INVX1  INVX1_522
timestamp 1598351757
transform 1 0 392 0 1 210
box -18 -6 52 210
use INVX1  INVX1_511
timestamp 1598351757
transform -1 0 392 0 1 210
box -18 -6 52 210
use INVX1  INVX1_330
timestamp 1598351757
transform 1 0 328 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_828
timestamp 1598351757
transform -1 0 296 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_654
timestamp 1598351757
transform -1 0 248 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_829
timestamp 1598351757
transform 1 0 152 0 1 210
box -16 -6 64 210
use INVX1  INVX1_534
timestamp 1598351757
transform -1 0 328 0 1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_730
timestamp 1598351757
transform 1 0 8 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_676
timestamp 1598351757
transform -1 0 152 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_680
timestamp 1598351757
transform -1 0 104 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_569
timestamp 1598351757
transform 1 0 4184 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_480
timestamp 1598351757
transform -1 0 4184 0 -1 210
box -16 -6 64 210
use FILL  FILL_1_2
timestamp 1598351757
transform -1 0 4264 0 -1 210
box -16 -6 32 210
use FILL  FILL_1_1
timestamp 1598351757
transform -1 0 4248 0 -1 210
box -16 -6 32 210
use NAND2X1  NAND2X1_580
timestamp 1598351757
transform 1 0 4056 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_571
timestamp 1598351757
transform 1 0 3976 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_244
timestamp 1598351757
transform -1 0 4136 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_452
timestamp 1598351757
transform 1 0 4024 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_359
timestamp 1598351757
transform -1 0 3912 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_434
timestamp 1598351757
transform 1 0 3944 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_282
timestamp 1598351757
transform -1 0 3944 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_671
timestamp 1598351757
transform -1 0 3864 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_260
timestamp 1598351757
transform 1 0 3688 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_283
timestamp 1598351757
transform 1 0 3800 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_661
timestamp 1598351757
transform -1 0 3800 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_222
timestamp 1598351757
transform -1 0 3768 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_858
timestamp 1598351757
transform -1 0 3688 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_851
timestamp 1598351757
transform -1 0 3608 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_672
timestamp 1598351757
transform 1 0 3608 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_277
timestamp 1598351757
transform -1 0 3560 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_349
timestamp 1598351757
transform 1 0 3480 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_830
timestamp 1598351757
transform 1 0 3368 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_221
timestamp 1598351757
transform 1 0 3448 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_276
timestamp 1598351757
transform 1 0 3416 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_105
timestamp 1598351757
transform 1 0 3288 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_102
timestamp 1598351757
transform -1 0 3368 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_101
timestamp 1598351757
transform 1 0 3256 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_106
timestamp 1598351757
transform -1 0 3256 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_114
timestamp 1598351757
transform 1 0 3176 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_248
timestamp 1598351757
transform 1 0 3128 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_285
timestamp 1598351757
transform -1 0 3128 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_342
timestamp 1598351757
transform 1 0 3032 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_147
timestamp 1598351757
transform -1 0 3000 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_662
timestamp 1598351757
transform 1 0 3000 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_239
timestamp 1598351757
transform -1 0 2952 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_149
timestamp 1598351757
transform -1 0 2888 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_148
timestamp 1598351757
transform 1 0 2760 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_131
timestamp 1598351757
transform -1 0 2920 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_132
timestamp 1598351757
transform 1 0 2808 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_286
timestamp 1598351757
transform 1 0 2712 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_288
timestamp 1598351757
transform -1 0 2680 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_240
timestamp 1598351757
transform -1 0 2712 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_847
timestamp 1598351757
transform -1 0 2568 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_820
timestamp 1598351757
transform -1 0 2520 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_241
timestamp 1598351757
transform -1 0 2632 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_133
timestamp 1598351757
transform -1 0 2600 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_848
timestamp 1598351757
transform 1 0 2392 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_846
timestamp 1598351757
transform 1 0 2312 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_668
timestamp 1598351757
transform -1 0 2472 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_667
timestamp 1598351757
transform 1 0 2360 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_815
timestamp 1598351757
transform -1 0 2312 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_814
timestamp 1598351757
transform 1 0 2184 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_644
timestamp 1598351757
transform -1 0 2264 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_643
timestamp 1598351757
transform 1 0 2152 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_819
timestamp 1598351757
transform -1 0 2120 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_649
timestamp 1598351757
transform 1 0 2120 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_650
timestamp 1598351757
transform 1 0 2040 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_554
timestamp 1598351757
transform -1 0 2040 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_152
timestamp 1598351757
transform 1 0 1960 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_726
timestamp 1598351757
transform 1 0 1912 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_575
timestamp 1598351757
transform -1 0 1912 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_569
timestamp 1598351757
transform -1 0 1880 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_731
timestamp 1598351757
transform -1 0 1816 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_209
timestamp 1598351757
transform 1 0 1720 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_570
timestamp 1598351757
transform -1 0 1848 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_574
timestamp 1598351757
transform -1 0 1720 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_738
timestamp 1598351757
transform -1 0 1688 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_834
timestamp 1598351757
transform -1 0 1608 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_476
timestamp 1598351757
transform -1 0 1640 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_612
timestamp 1598351757
transform 1 0 1480 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_796
timestamp 1598351757
transform 1 0 1432 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_614
timestamp 1598351757
transform -1 0 1560 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_626
timestamp 1598351757
transform -1 0 1432 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_803
timestamp 1598351757
transform -1 0 1368 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_797
timestamp 1598351757
transform -1 0 1288 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_137
timestamp 1598351757
transform -1 0 1400 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_627
timestamp 1598351757
transform 1 0 1288 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_779
timestamp 1598351757
transform -1 0 1208 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_708
timestamp 1598351757
transform -1 0 1160 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_613
timestamp 1598351757
transform 1 0 1208 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_609
timestamp 1598351757
transform -1 0 1112 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_783
timestamp 1598351757
transform -1 0 1080 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_780
timestamp 1598351757
transform 1 0 952 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_610
timestamp 1598351757
transform 1 0 1000 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_743
timestamp 1598351757
transform -1 0 952 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_782
timestamp 1598351757
transform 1 0 792 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_612
timestamp 1598351757
transform 1 0 872 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_611
timestamp 1598351757
transform -1 0 872 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_747
timestamp 1598351757
transform -1 0 792 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_155
timestamp 1598351757
transform -1 0 712 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_143
timestamp 1598351757
transform -1 0 744 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_144
timestamp 1598351757
transform 1 0 632 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_678
timestamp 1598351757
transform -1 0 600 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_740
timestamp 1598351757
transform -1 0 520 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_535
timestamp 1598351757
transform -1 0 632 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_581
timestamp 1598351757
transform -1 0 552 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_739
timestamp 1598351757
transform -1 0 440 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_407
timestamp 1598351757
transform -1 0 360 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_582
timestamp 1598351757
transform 1 0 440 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_331
timestamp 1598351757
transform -1 0 392 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_661
timestamp 1598351757
transform -1 0 248 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_332
timestamp 1598351757
transform -1 0 312 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_514
timestamp 1598351757
transform -1 0 280 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_515
timestamp 1598351757
transform 1 0 168 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_679
timestamp 1598351757
transform 1 0 120 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_728
timestamp 1598351757
transform -1 0 88 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_573
timestamp 1598351757
transform 1 0 88 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_571
timestamp 1598351757
transform -1 0 40 0 -1 210
box -18 -6 52 210
<< labels >>
rlabel metal2 s 2064 3080 2064 3080 6 INPUT_0
port 0 nsew
rlabel metal2 s 2880 -40 2880 -40 8 INPUT_1
port 1 nsew
rlabel metal2 s 4064 3080 4064 3080 6 INPUT_2
port 2 nsew
rlabel metal2 s 3968 3080 3968 3080 6 INPUT_3
port 3 nsew
rlabel metal3 s -48 2260 -48 2260 4 INPUT_4
port 4 nsew
rlabel metal3 s -48 2500 -48 2500 4 INPUT_5
port 5 nsew
rlabel metal3 s -48 2960 -48 2960 4 INPUT_6
port 6 nsew
rlabel metal2 s 144 3080 144 3080 6 INPUT_7
port 7 nsew
rlabel metal2 s 1584 3080 1584 3080 6 GATE_222
port 8 nsew
rlabel metal3 s -48 1920 -48 1920 4 GATE_366
port 9 nsew
rlabel metal3 s 4320 120 4320 120 6 GATE_479
port 10 nsew
rlabel metal3 s 4320 180 4320 180 6 GATE_579
port 11 nsew
rlabel metal2 s 2560 -40 2560 -40 8 GATE_662
port 12 nsew
rlabel metal2 s 592 -40 592 -40 8 GATE_741
port 13 nsew
rlabel metal3 s -48 1780 -48 1780 4 GATE_811
port 14 nsew
rlabel metal3 s -48 1520 -48 1520 4 GATE_865
port 15 nsew
rlabel metal3 s -48 2760 -48 2760 4 gate
port 16 nsew
rlabel metal3 s -48 1160 -48 1160 4 type:
port 17 nsew
rlabel metal2 s 3584 -40 3584 -40 8 NAND;
port 18 nsew
rlabel metal3 s -48 1280 -48 1280 4 name:
port 19 nsew
rlabel metal3 s -48 360 -48 360 4 GATE_0_I0
port 20 nsew
rlabel space -412 -43 4682 3083 1 vdd
rlabel space -412 -43 4682 3083 1 gnd
<< end >>
