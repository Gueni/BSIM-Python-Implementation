magic
tech scmos
magscale 1 2
timestamp 1611069007
<< nwell >>
rect -16 96 64 210
<< ntransistor >>
rect 14 12 18 32
rect 30 12 34 32
<< ptransistor >>
rect 14 108 18 188
rect 24 108 28 188
<< ndiffusion >>
rect 4 31 14 32
rect 12 13 14 31
rect 4 12 14 13
rect 18 31 30 32
rect 18 13 20 31
rect 28 13 30 31
rect 18 12 30 13
rect 34 31 44 32
rect 34 13 36 31
rect 34 12 44 13
<< pdiffusion >>
rect 4 186 14 188
rect 12 108 14 186
rect 18 108 24 188
rect 28 186 38 188
rect 28 108 30 186
<< ndcontact >>
rect 4 13 12 31
rect 20 13 28 31
rect 36 13 44 31
<< pdcontact >>
rect 4 108 12 186
rect 30 108 38 186
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
<< polysilicon >>
rect 14 188 18 192
rect 24 188 28 192
rect 14 46 18 108
rect 24 106 28 108
rect 24 102 34 106
rect 12 38 18 46
rect 14 32 18 38
rect 30 94 36 102
rect 30 32 34 94
rect 14 8 18 12
rect 30 8 34 12
<< polycontact >>
rect 4 38 12 46
rect 36 94 44 102
<< metal1 >>
rect -4 204 52 206
rect 4 196 28 204
rect 36 196 52 204
rect -4 194 52 196
rect 4 186 12 194
rect 30 186 38 188
rect 20 108 30 116
rect 22 74 28 108
rect 36 86 44 94
rect 20 66 28 74
rect 4 46 12 54
rect 22 32 28 66
rect 4 31 12 32
rect 4 6 12 13
rect 20 31 28 32
rect 20 12 28 13
rect 36 31 44 32
rect 36 6 44 13
rect -4 4 52 6
rect 4 -4 28 4
rect 36 -4 52 4
rect -4 -6 52 -4
<< m1p >>
rect 36 86 44 94
rect 20 66 28 74
rect 4 46 12 54
<< labels >>
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 40 90 40 90 4 B
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 24 70 24 70 4 Y
rlabel metal1 8 50 8 50 4 A
rlabel ptransistor 24 164 24 164 1 S$
rlabel ptransistor 14 164 14 164 1 S$
rlabel ptransistor 18 164 18 164 1 D$
rlabel ptransistor 28 164 28 164 1 D$
rlabel ntransistor 18 22 18 22 1 D$
rlabel ntransistor 14 24 14 24 1 S$
rlabel ntransistor 34 22 34 22 1 S$
rlabel ntransistor 30 24 30 24 1 D$
rlabel space -16 -6 64 210 1 vdd
rlabel space -16 -6 64 210 1 gnd
<< end >>
