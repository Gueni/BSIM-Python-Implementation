*** TEST 004 - partitioning ***
*
* ngSPICE test for PLS experiments
*
* AES SBOX PLS test init file generator - protected dualRail SBOX area illuminated
*
* Author: Jan Belohoubek, 08/2020
* jan.belohoubek@fit.cvut.cz
*
* https://users.fit.cvut.cz/~belohja4/
*
*
* **************************************

.include ../../models.lib
.include ../../tsmc180nmcmos.lib
.include pDualRail.spice

* **************************************
* --- Test ---
* **************************************

* --- Settings
.param showPlots = 0
.param writeFile = 1
.param run_inputSet = 0

* redefine defaults ...
.include test00X_settings.inc

.csparam showPlots = {showPlots}
.csparam writeFile = {writeFile}
.csparam run_inputSet = {run_inputSet}

.global showPlots writeFile run_inputSet

* --- End of Settins

Vtrig LaserTrig 0 0 PWL(0ns 0V 20ns 0V 21ns SUPP)

.param beamDistanceTop = 0
.param beamDistanceBot = 0

.global LaserTrig beamDistanceTop beamDistanceBot

* --- inputs
Vvin0 INPUT_0 0 0 PWL(0ns 0V 5ns  0V 7ns  0V)
Vvin1 INPUT_1 0 0 PWL(0ns 0V 6ns  0V 8ns  0V)
Vvin2 INPUT_2 0 0 PWL(0ns 0V 7ns  0V 9ns  0V)
Vvin3 INPUT_3 0 0 PWL(0ns 0V 8ns  0V 10ns 0V)
Vvin4 INPUT_4 0 0 PWL(0ns 0V 9ns  0V 11ns 0V)
Vvin5 INPUT_5 0 0 PWL(0ns 0V 10ns 0V 12ns 0V)
Vvin6 INPUT_6 0 0 PWL(0ns 0V 11ns 0V 13ns 0V)
Vvin7 INPUT_7 0 0 PWL(0ns 0V 12ns 0V 14ns 0V)

Vvin0D D_INPUT_0 0 0 PWL(0ns 0V 5ns  0V 7ns  0V)
Vvin1D D_INPUT_1 0 0 PWL(0ns 0V 6ns  0V 8ns  0V)
Vvin2D D_INPUT_2 0 0 PWL(0ns 0V 7ns  0V 9ns  0V)
Vvin3D D_INPUT_3 0 0 PWL(0ns 0V 8ns  0V 10ns 0V)
Vvin4D D_INPUT_4 0 0 PWL(0ns 0V 9ns  0V 11ns 0V)
Vvin5D D_INPUT_5 0 0 PWL(0ns 0V 10ns 0V 12ns 0V)
Vvin6D D_INPUT_6 0 0 PWL(0ns 0V 11ns 0V 13ns 0V)
Vvin7D D_INPUT_7 0 0 PWL(0ns 0V 12ns 0V 14ns 0V)


* --- circuit layout model

Xsbox1 
+ POR2X1_751/A POR2X1_516/B PAND2X1_809/A PAND2X1_473/B POR2X1_101/A POR2X1_334/A POR2X1_836/A POR2X1_240/A POR2X1_461/Y PAND2X1_691/Y POR2X1_323/Y POR2X1_527/Y POR2X1_111/Y POR2X1_515/Y POR2X1_73/Y POR2X1_41/B POR2X1_669/B PAND2X1_63/B POR2X1_16/A POR2X1_287/B POR2X1_246/Y PAND2X1_464/B POR2X1_815/A POR2X1_309/Y POR2X1_283/Y POR2X1_488/Y POR2X1_289/Y POR2X1_417/Y POR2X1_226/Y PAND2X1_848/B POR2X1_96/B POR2X1_62/Y PAND2X1_90/Y POR2X1_612/A POR2X1_78/A PAND2X1_55/Y POR2X1_590/A POR2X1_378/Y POR2X1_274/B POR2X1_838/B POR2X1_195/A POR2X1_296/Y POR2X1_447/B POR2X1_535/A POR2X1_138/A POR2X1_519/Y POR2X1_692/Y POR2X1_48/Y POR2X1_406/A POR2X1_599/A POR2X1_763/Y 
+ POR2X1_511/Y POR2X1_98/B POR2X1_448/A POR2X1_630/B POR2X1_389/A POR2X1_631/A POR2X1_294/Y POR2X1_415/Y POR2X1_637/B POR2X1_828/A POR2X1_398/Y POR2X1_121/Y POR2X1_302/A POR2X1_450/B POR2X1_606/Y POR2X1_301/A POR2X1_543/A POR2X1_322/Y POR2X1_164/Y POR2X1_144/Y POR2X1_306/Y POR2X1_696/Y POR2X1_503/A POR2X1_588/Y POR2X1_376/Y POR2X1_273/Y POR2X1_433/Y POR2X1_409/B POR2X1_743/Y PAND2X1_156/B POR2X1_673/A POR2X1_549/A POR2X1_391/B POR2X1_619/Y POR2X1_532/A POR2X1_130/A POR2X1_266/A POR2X1_634/A PAND2X1_73/Y PAND2X1_85/Y POR2X1_541/B POR2X1_633/A POR2X1_777/B PAND2X1_39/B POR2X1_186/B POR2X1_83/A POR2X1_77/Y POR2X1_693/Y POR2X1_23/Y POR2X1_49/Y POR2X1_748/A 
+ PAND2X1_377/Y POR2X1_387/Y POR2X1_329/Y POR2X1_421/Y POR2X1_597/A POR2X1_72/B POR2X1_40/Y POR2X1_416/B POR2X1_7/B POR2X1_790/B POR2X1_694/Y POR2X1_426/Y PAND2X1_52/B PAND2X1_32/B PAND2X1_57/B PAND2X1_48/B POR2X1_304/Y POR2X1_56/Y POR2X1_409/Y POR2X1_635/A POR2X1_769/B POR2X1_430/Y PAND2X1_69/A PAND2X1_20/A POR2X1_260/A POR2X1_52/A POR2X1_96/A POR2X1_65/A POR2X1_513/Y POR2X1_855/B POR2X1_325/A POR2X1_547/B POR2X1_332/B POR2X1_557/A POR2X1_411/B POR2X1_394/A POR2X1_344/A PAND2X1_19/Y POR2X1_7/A POR2X1_748/Y POR2X1_516/A POR2X1_750/Y POR2X1_129/Y POR2X1_29/Y POR2X1_383/A POR2X1_68/A POR2X1_614/A POR2X1_81/A POR2X1_291/Y POR2X1_824/Y POR2X1_234/Y 
+ PAND2X1_462/B POR2X1_809/B POR2X1_276/Y PAND2X1_101/B POR2X1_708/B POR2X1_638/B POR2X1_459/B POR2X1_325/B POR2X1_776/B POR2X1_147/A POR2X1_502/Y POR2X1_308/B POR2X1_155/Y POR2X1_274/A POR2X1_832/A POR2X1_780/B POR2X1_407/Y POR2X1_458/Y PAND2X1_48/Y POR2X1_405/Y POR2X1_513/B POR2X1_520/A POR2X1_706/B POR2X1_335/B POR2X1_286/B POR2X1_489/A POR2X1_814/Y POR2X1_333/A POR2X1_446/B POR2X1_227/A POR2X1_481/A POR2X1_416/A POR2X1_625/Y POR2X1_399/A POR2X1_585/Y POR2X1_257/A PAND2X1_81/B PAND2X1_82/Y POR2X1_38/Y POR2X1_87/B POR2X1_236/Y POR2X1_382/Y POR2X1_300/Y POR2X1_369/Y POR2X1_607/A POR2X1_299/Y POR2X1_122/A POR2X1_848/A POR2X1_750/B POR2X1_294/B POR2X1_342/B 
+ POR2X1_78/B POR2X1_278/Y POR2X1_102/Y PAND2X1_612/B POR2X1_55/Y PAND2X1_94/Y POR2X1_90/Y POR2X1_136/Y POR2X1_43/Y POR2X1_297/A POR2X1_272/Y POR2X1_827/Y POR2X1_419/Y POR2X1_459/A POR2X1_534/Y POR2X1_814/B PAND2X1_6/Y POR2X1_490/Y POR2X1_20/A PAND2X1_23/Y POR2X1_256/Y POR2X1_789/B POR2X1_93/Y POR2X1_422/Y POR2X1_628/Y POR2X1_63/Y POR2X1_672/Y PAND2X1_71/Y POR2X1_68/Y POR2X1_198/B POR2X1_778/B POR2X1_335/A POR2X1_71/Y POR2X1_57/Y POR2X1_69/A POR2X1_372/A POR2X1_310/Y POR2X1_378/A POR2X1_706/A POR2X1_709/A POR2X1_622/B POR2X1_85/Y POR2X1_263/Y POR2X1_413/A POR2X1_278/A POR2X1_255/Y POR2X1_245/Y POR2X1_150/Y PAND2X1_63/Y PAND2X1_549/B POR2X1_355/B 
+ POR2X1_448/B POR2X1_596/Y PAND2X1_96/B POR2X1_260/B PAND2X1_60/B POR2X1_43/B POR2X1_39/B POR2X1_83/B POR2X1_66/B PAND2X1_72/A PAND2X1_41/B POR2X1_753/Y PAND2X1_65/B PAND2X1_58/A POR2X1_66/A PAND2X1_56/Y POR2X1_307/B POR2X1_707/B POR2X1_13/A POR2X1_60/A POR2X1_20/B POR2X1_32/A POR2X1_57/A POR2X1_48/A POR2X1_582/Y POR2X1_460/A POR2X1_451/A POR2X1_760/A POR2X1_66/Y POR2X1_121/A POR2X1_188/A POR2X1_327/Y POR2X1_67/A POR2X1_666/A POR2X1_816/A PAND2X1_687/Y POR2X1_271/A POR2X1_87/Y POR2X1_410/Y POR2X1_373/Y POR2X1_667/A POR2X1_411/A POR2X1_687/Y POR2X1_270/Y POR2X1_88/A POR2X1_544/B POR2X1_264/Y POR2X1_683/Y POR2X1_682/Y POR2X1_685/A POR2X1_686/B 
+ POR2X1_88/Y PAND2X1_717/A POR2X1_761/A POR2X1_644/A POR2X1_717/B PAND2X1_88/Y 
+ VSS VDD 
+ POR2X1_452/A POR2X1_460/Y PAND2X1_635/Y POR2X1_152/Y POR2X1_612/B POR2X1_103/Y POR2X1_106/Y POR2X1_695/Y POR2X1_280/Y POR2X1_601/Y POR2X1_248/Y POR2X1_394/Y POR2X1_747/Y POR2X1_524/Y POR2X1_399/Y POR2X1_528/Y POR2X1_122/Y POR2X1_45/Y POR2X1_485/Y POR2X1_297/Y POR2X1_424/Y POR2X1_744/Y POR2X1_701/Y POR2X1_757/Y POR2X1_526/Y POR2X1_517/Y POR2X1_315/Y POR2X1_74/Y POR2X1_32/Y POR2X1_491/Y POR2X1_109/Y POR2X1_600/Y POR2X1_230/Y POR2X1_298/Y POR2X1_224/Y POR2X1_428/Y POR2X1_583/Y POR2X1_505/Y POR2X1_20/Y POR2X1_79/Y POR2X1_666/Y POR2X1_496/Y POR2X1_432/Y POR2X1_607/Y POR2X1_257/Y POR2X1_521/Y POR2X1_81/Y POR2X1_60/Y POR2X1_135/Y POR2X1_75/Y POR2X1_492/Y 
+ POR2X1_482/Y POR2X1_108/Y POR2X1_295/Y POR2X1_437/Y POR2X1_609/Y POR2X1_700/Y POR2X1_755/Y POR2X1_395/Y POR2X1_131/Y POR2X1_261/A POR2X1_679/A POR2X1_13/Y POR2X1_494/Y POR2X1_603/Y POR2X1_229/Y POR2X1_765/Y POR2X1_380/A POR2X1_707/Y POR2X1_307/Y POR2X1_197/Y POR2X1_379/Y POR2X1_334/B POR2X1_678/A POR2X1_84/A POR2X1_668/Y POR2X1_241/B POR2X1_34/B POR2X1_643/A POR2X1_538/A POR2X1_180/B POR2X1_844/B POR2X1_623/B POR2X1_33/A POR2X1_61/B POR2X1_523/A POR2X1_835/A POR2X1_709/B POR2X1_720/B POR2X1_343/B POR2X1_855/A POR2X1_832/B PAND2X1_65/Y POR2X1_593/B POR2X1_770/A POR2X1_324/A POR2X1_509/A POR2X1_703/A POR2X1_830/A POR2X1_520/B POR2X1_169/A PAND2X1_790/Y 
+ POR2X1_346/B POR2X1_443/A POR2X1_444/B POR2X1_620/A POR2X1_786/A POR2X1_267/B PAND2X1_41/Y POR2X1_610/Y POR2X1_769/A POR2X1_400/B POR2X1_781/B POR2X1_549/B POR2X1_391/A POR2X1_174/B POR2X1_540/A POR2X1_191/B POR2X1_169/B POR2X1_758/Y POR2X1_673/B POR2X1_835/B POR2X1_123/B POR2X1_123/A POR2X1_675/A POR2X1_501/B PAND2X1_72/Y POR2X1_605/A POR2X1_450/A POR2X1_544/A POR2X1_637/A POR2X1_174/A POR2X1_175/B POR2X1_180/A POR2X1_128/A POR2X1_555/A PAND2X1_7/Y POR2X1_719/B POR2X1_789/A POR2X1_194/B POR2X1_773/B POR2X1_402/B POR2X1_307/A POR2X1_311/Y POR2X1_176/Y POR2X1_83/Y POR2X1_669/A POR2X1_290/Y POR2X1_27/Y POR2X1_677/Y POR2X1_237/Y POR2X1_595/Y POR2X1_146/Y 
+ POR2X1_179/Y POR2X1_69/Y POR2X1_484/Y POR2X1_495/Y POR2X1_39/Y POR2X1_754/Y POR2X1_396/Y POR2X1_320/Y POR2X1_24/Y POR2X1_58/Y POR2X1_497/Y POR2X1_615/Y POR2X1_522/Y POR2X1_493/A POR2X1_483/A POR2X1_114/B POR2X1_84/B POR2X1_346/A POR2X1_61/A POR2X1_76/A POR2X1_440/B POR2X1_646/A POR2X1_710/B POR2X1_791/B POR2X1_401/B POR2X1_702/A POR2X1_558/A POR2X1_605/B POR2X1_260/Y POR2X1_678/Y POR2X1_193/A POR2X1_231/B POR2X1_770/B POR2X1_140/A POR2X1_447/A POR2X1_489/B POR2X1_98/A POR2X1_734/B POR2X1_653/B POR2X1_788/B POR2X1_456/B POR2X1_137/B POR2X1_768/A POR2X1_192/B POR2X1_128/B POR2X1_644/B POR2X1_448/Y POR2X1_356/A PAND2X1_565/A POR2X1_292/Y POR2X1_152/A 
+ POR2X1_173/Y PAND2X1_784/A PAND2X1_553/B PAND2X1_633/Y PAND2X1_640/B POR2X1_813/Y POR2X1_235/Y POR2X1_624/B POR2X1_711/B POR2X1_713/A PAND2X1_337/A PAND2X1_778/Y PAND2X1_198/Y POR2X1_72/Y POR2X1_184/Y POR2X1_335/Y POR2X1_784/A POR2X1_208/A POR2X1_202/A PAND2X1_673/Y POR2X1_65/Y POR2X1_117/Y POR2X1_262/Y PAND2X1_632/A PAND2X1_453/A POR2X1_789/Y PAND2X1_348/A POR2X1_707/A POR2X1_702/B POR2X1_776/A POR2X1_249/Y POR2X1_401/A POR2X1_507/A PAND2X1_561/A POR2X1_130/Y POR2X1_156/B POR2X1_231/A POR2X1_636/A POR2X1_247/Y POR2X1_620/B POR2X1_602/B POR2X1_345/A POR2X1_105/Y POR2X1_756/Y POR2X1_181/A PAND2X1_535/Y POR2X1_459/Y PAND2X1_454/B PAND2X1_506/Y PAND2X1_852/A PAND2X1_199/A 
+ PAND2X1_139/B POR2X1_132/Y POR2X1_305/Y POR2X1_384/A POR2X1_766/Y POR2X1_91/Y POR2X1_312/Y POR2X1_178/Y POR2X1_67/Y POR2X1_613/Y POR2X1_647/B POR2X1_670/Y POR2X1_822/Y POR2X1_420/Y POR2X1_591/A POR2X1_533/A POR2X1_239/Y POR2X1_172/Y PAND2X1_843/Y PAND2X1_287/Y POR2X1_602/A POR2X1_78/Y POR2X1_240/B POR2X1_446/A POR2X1_608/Y POR2X1_342/Y POR2X1_486/B POR2X1_546/B POR2X1_507/B POR2X1_720/A POR2X1_546/A POR2X1_848/Y PAND2X1_303/B PAND2X1_787/A PAND2X1_552/B PAND2X1_831/Y PAND2X1_716/B PAND2X1_392/B POR2X1_823/Y POR2X1_697/Y POR2X1_759/Y POR2X1_34/A POR2X1_250/A POR2X1_393/Y PAND2X1_156/A POR2X1_498/A POR2X1_134/Y POR2X1_679/B POR2X1_754/A POR2X1_427/Y PAND2X1_638/B 
+ PAND2X1_632/B POR2X1_416/Y POR2X1_481/Y POR2X1_509/B POR2X1_454/B POR2X1_704/Y POR2X1_333/Y POR2X1_557/B POR2X1_286/Y POR2X1_370/Y POR2X1_559/A POR2X1_834/Y POR2X1_783/B POR2X1_196/Y POR2X1_464/Y POR2X1_828/Y POR2X1_783/A POR2X1_832/Y POR2X1_841/B POR2X1_156/Y POR2X1_353/A POR2X1_149/B POR2X1_170/B POR2X1_785/A POR2X1_326/A POR2X1_638/Y POR2X1_712/A PAND2X1_656/A POR2X1_476/A POR2X1_362/A POR2X1_809/Y PAND2X1_472/A PAND2X1_243/B PAND2X1_839/B PAND2X1_338/B POR2X1_676/Y POR2X1_259/B POR2X1_614/Y POR2X1_545/A POR2X1_445/A PAND2X1_52/Y POR2X1_636/B POR2X1_523/B POR2X1_782/B POR2X1_836/B POR2X1_779/A POR2X1_542/B POR2X1_635/B POR2X1_710/A POR2X1_792/B POR2X1_383/Y 
+ POR2X1_131/A POR2X1_586/Y POR2X1_516/Y PAND2X1_793/A POR2X1_248/A POR2X1_423/Y POR2X1_584/Y POR2X1_7/Y POR2X1_183/Y POR2X1_33/B POR2X1_344/Y POR2X1_127/Y POR2X1_698/Y POR2X1_764/Y POR2X1_380/Y POR2X1_251/A POR2X1_125/Y POR2X1_442/Y POR2X1_261/Y POR2X1_757/A POR2X1_561/B POR2X1_112/Y POR2X1_332/Y POR2X1_550/A POR2X1_729/Y POR2X1_855/Y POR2X1_574/A POR2X1_503/Y POR2X1_142/Y POR2X1_518/Y POR2X1_167/Y POR2X1_667/Y POR2X1_250/Y POR2X1_829/Y POR2X1_591/Y POR2X1_321/Y POR2X1_189/Y POR2X1_96/Y POR2X1_487/Y POR2X1_406/Y POR2X1_759/A POR2X1_594/Y POR2X1_533/Y POR2X1_525/Y POR2X1_163/Y POR2X1_165/Y POR2X1_145/Y POR2X1_52/Y POR2X1_680/Y POR2X1_251/Y POR2X1_418/Y 
+ POR2X1_238/Y POR2X1_462/B POR2X1_259/A POR2X1_781/A POR2X1_181/B POR2X1_210/B POR2X1_719/A POR2X1_499/A POR2X1_435/B POR2X1_646/B PAND2X1_79/Y POR2X1_833/A POR2X1_194/A POR2X1_790/A POR2X1_324/B POR2X1_148/A PAND2X1_452/B POR2X1_769/Y POR2X1_635/Y PAND2X1_460/Y PAND2X1_197/Y PAND2X1_308/B POR2X1_554/B POR2X1_342/A POR2X1_400/A POR2X1_209/A POR2X1_113/B POR2X1_705/B POR2X1_347/B POR2X1_449/A POR2X1_780/A POR2X1_791/A POR2X1_403/B POR2X1_124/B POR2X1_493/B POR2X1_775/A POR2X1_302/B POR2X1_76/B POR2X1_227/B POR2X1_559/B POR2X1_97/A POR2X1_343/A POR2X1_506/B POR2X1_210/A POR2X1_168/A POR2X1_148/B POR2X1_728/A PAND2X1_452/A PAND2X1_707/Y POR2X1_793/A POR2X1_16/Y 
+ POR2X1_665/Y POR2X1_751/Y POR2X1_767/Y POR2X1_397/Y POR2X1_504/Y POR2X1_158/Y POR2X1_232/Y POR2X1_258/Y POR2X1_746/Y POR2X1_187/Y POR2X1_166/Y POR2X1_41/Y POR2X1_441/Y POR2X1_265/Y POR2X1_745/Y POR2X1_531/Y POR2X1_384/Y POR2X1_171/Y POR2X1_177/Y POR2X1_821/Y POR2X1_118/Y POR2X1_674/Y POR2X1_498/Y POR2X1_604/Y POR2X1_438/Y POR2X1_597/Y PAND2X1_356/B PAND2X1_389/Y PAND2X1_711/A PAND2X1_713/B POR2X1_665/A POR2X1_79/A POR2X1_151/Y POR2X1_188/Y POR2X1_590/Y POR2X1_777/Y POR2X1_633/Y POR2X1_553/A POR2X1_243/B POR2X1_664/Y POR2X1_640/A POR2X1_845/A POR2X1_460/B POR2X1_532/Y PAND2X1_624/A POR2X1_391/Y POR2X1_565/B POR2X1_673/Y POR2X1_158/B PAND2X1_783/B POR2X1_829/A 
+ PAND2X1_841/B PAND2X1_459/Y PAND2X1_651/A PAND2X1_712/B PAND2X1_308/Y PAND2X1_149/A PAND2X1_776/Y PAND2X1_168/Y PAND2X1_326/B POR2X1_552/A POR2X1_303/B POR2X1_450/Y POR2X1_302/Y POR2X1_638/A POR2X1_632/A POR2X1_389/Y POR2X1_632/B PAND2X1_840/B PAND2X1_779/Y PAND2X1_769/Y PAND2X1_199/B PAND2X1_642/B POR2X1_139/A POR2X1_567/B POR2X1_508/B POR2X1_454/A POR2X1_199/B POR2X1_852/B POR2X1_202/B POR2X1_612/Y PAND2X1_859/A PAND2X1_340/B PAND2X1_446/Y PAND2X1_714/B PAND2X1_333/Y PAND2X1_557/A PAND2X1_288/A PAND2X1_464/Y PAND2X1_349/A POR2X1_850/A POR2X1_288/A POR2X1_609/A POR2X1_669/Y PAND2X1_332/Y PAND2X1_115/B PAND2X1_550/B PAND2X1_856/B PAND2X1_730/B POR2X1_472/B POR2X1_243/A POR2X1_836/Y 
+ POR2X1_334/Y POR2X1_101/Y PAND2X1_473/Y PAND2X1_362/B PAND2X1_810/B PAND2X1_687/Y POR2X1_687/Y PAND2X1_254/Y POR2X1_254/Y PAND2X1_97/Y POR2X1_802/B POR2X1_802/A POR2X1_99/B PAND2X1_802/B PAND2X1_798/Y POR2X1_113/Y POR2X1_319/Y POR2X1_567/A PAND2X1_114/B PAND2X1_539/Y PAND2X1_354/A POR2X1_436/B POR2X1_537/Y POR2X1_592/Y PAND2X1_592/Y PAND2X1_643/A PAND2X1_436/A PAND2X1_593/Y POR2X1_652/A POR2X1_116/Y POR2X1_88/Y PAND2X1_717/A POR2X1_761/A POR2X1_373/Y POR2X1_644/A PAND2X1_216/B POR2X1_717/B PAND2X1_88/Y POR2X1_483/B POR2X1_544/B POR2X1_252/Y PAND2X1_267/Y PAND2X1_631/A PAND2X1_798/B POR2X1_631/B POR2X1_468/B POR2X1_267/Y 
+ AES_SBOX_1

.include outputs_0.plw

* **************************************
* --- Simulation Settings ---
* **************************************

.param SIM_LEN = 35ns
.csparam SIM_LEN = {SIM_LEN}

.tran 0.1ns 'SIM_LEN'
.param SIMSTEP = 'SIM_LEN/0.1ns'
.csparam SIMSTEP = {SIMSTEP}

* **************************************
* --- Simulation Control ---
* **************************************

.control
    .include ../inputsD.inc

    run
    
    if ('writeFile' > 0)   
      wrdata ivdd_1.out i(vvdd)
      wrdata ivss_1.out i(vvss)
      *snsave sim_1.snap
    end
    
    set wr_vecnames
    set wr_singlescale
    wrdata outputs_1.out V("POR2X1_452/A") V("POR2X1_460/Y") V("PAND2X1_635/Y") V("POR2X1_152/Y") V("POR2X1_612/B") V("POR2X1_103/Y") V("POR2X1_106/Y") V("POR2X1_695/Y") V("POR2X1_280/Y") V("POR2X1_601/Y") V("POR2X1_248/Y") V("POR2X1_394/Y") V("POR2X1_747/Y") V("POR2X1_524/Y") V("POR2X1_399/Y") V("POR2X1_528/Y") V("POR2X1_122/Y") V("POR2X1_45/Y") V("POR2X1_485/Y") V("POR2X1_297/Y") V("POR2X1_424/Y") V("POR2X1_744/Y") V("POR2X1_701/Y") V("POR2X1_757/Y") V("POR2X1_526/Y") V("POR2X1_517/Y") V("POR2X1_315/Y") V("POR2X1_74/Y") V("POR2X1_32/Y") V("POR2X1_491/Y") V("POR2X1_109/Y") V("POR2X1_600/Y") V("POR2X1_230/Y") V("POR2X1_298/Y") V("POR2X1_224/Y") V("POR2X1_428/Y") V("POR2X1_583/Y") V("POR2X1_505/Y") V("POR2X1_20/Y") V("POR2X1_79/Y") V("POR2X1_666/Y") V("POR2X1_496/Y") V("POR2X1_432/Y") V("POR2X1_607/Y") V("POR2X1_257/Y") V("POR2X1_521/Y") V("POR2X1_81/Y") V("POR2X1_60/Y") V("POR2X1_135/Y") V("POR2X1_75/Y") V("POR2X1_492/Y") V("POR2X1_482/Y") V("POR2X1_108/Y") V("POR2X1_295/Y") V("POR2X1_437/Y") V("POR2X1_609/Y") V("POR2X1_700/Y") V("POR2X1_755/Y") V("POR2X1_395/Y") V("POR2X1_131/Y") V("POR2X1_261/A") V("POR2X1_679/A") V("POR2X1_13/Y") V("POR2X1_494/Y") V("POR2X1_603/Y") V("POR2X1_229/Y") V("POR2X1_765/Y") V("POR2X1_380/A") V("POR2X1_707/Y") V("POR2X1_307/Y") V("POR2X1_197/Y") V("POR2X1_379/Y") V("POR2X1_334/B") V("POR2X1_678/A") V("POR2X1_84/A") V("POR2X1_668/Y") V("POR2X1_241/B") V("POR2X1_34/B") V("POR2X1_643/A") V("POR2X1_538/A") V("POR2X1_180/B") V("POR2X1_844/B") V("POR2X1_623/B") V("POR2X1_33/A") V("POR2X1_61/B") V("POR2X1_523/A") V("POR2X1_835/A") V("POR2X1_709/B") V("POR2X1_720/B") V("POR2X1_343/B") V("POR2X1_855/A") V("POR2X1_832/B") V("PAND2X1_65/Y") V("POR2X1_593/B") V("POR2X1_770/A") V("POR2X1_324/A") V("POR2X1_509/A") V("POR2X1_703/A") V("POR2X1_830/A") V("POR2X1_520/B") V("POR2X1_169/A") V("PAND2X1_790/Y") V("POR2X1_346/B") V("POR2X1_443/A") V("POR2X1_444/B") V("POR2X1_620/A") V("POR2X1_786/A") V("POR2X1_267/B") V("PAND2X1_41/Y") V("POR2X1_610/Y") V("POR2X1_769/A") V("POR2X1_400/B") V("POR2X1_781/B") V("POR2X1_549/B") V("POR2X1_391/A") V("POR2X1_174/B") V("POR2X1_540/A") V("POR2X1_191/B") V("POR2X1_169/B") V("POR2X1_758/Y") V("POR2X1_673/B") V("POR2X1_835/B") V("POR2X1_123/B") V("POR2X1_123/A") V("POR2X1_675/A") V("POR2X1_501/B") V("PAND2X1_72/Y") V("POR2X1_605/A") V("POR2X1_450/A") V("POR2X1_544/A") V("POR2X1_637/A") V("POR2X1_174/A") V("POR2X1_175/B") V("POR2X1_180/A") V("POR2X1_128/A") V("POR2X1_555/A") V("PAND2X1_7/Y") V("POR2X1_719/B") V("POR2X1_789/A") V("POR2X1_194/B") V("POR2X1_773/B") V("POR2X1_402/B") V("POR2X1_307/A") V("POR2X1_311/Y") V("POR2X1_176/Y") V("POR2X1_83/Y") V("POR2X1_669/A") V("POR2X1_290/Y") V("POR2X1_27/Y") V("POR2X1_677/Y") V("POR2X1_237/Y") V("POR2X1_595/Y") V("POR2X1_146/Y") V("POR2X1_179/Y") V("POR2X1_69/Y") V("POR2X1_484/Y") V("POR2X1_495/Y") V("POR2X1_39/Y") V("POR2X1_754/Y") V("POR2X1_396/Y") V("POR2X1_320/Y") V("POR2X1_24/Y") V("POR2X1_58/Y") V("POR2X1_497/Y") V("POR2X1_615/Y") V("POR2X1_522/Y") V("POR2X1_493/A") V("POR2X1_483/A") V("POR2X1_114/B") V("POR2X1_84/B") V("POR2X1_346/A") V("POR2X1_61/A") V("POR2X1_76/A") V("POR2X1_440/B") V("POR2X1_646/A") V("POR2X1_710/B") V("POR2X1_791/B") V("POR2X1_401/B") V("POR2X1_702/A") V("POR2X1_558/A") V("POR2X1_605/B") V("POR2X1_260/Y") V("POR2X1_678/Y") V("POR2X1_193/A") V("POR2X1_231/B") V("POR2X1_770/B") V("POR2X1_140/A") V("POR2X1_447/A") V("POR2X1_489/B") V("POR2X1_98/A") V("POR2X1_734/B") V("POR2X1_653/B") V("POR2X1_788/B") V("POR2X1_456/B") V("POR2X1_137/B") V("POR2X1_768/A") V("POR2X1_192/B") V("POR2X1_128/B") V("POR2X1_644/B") V("POR2X1_448/Y") V("POR2X1_356/A") V("PAND2X1_565/A") V("POR2X1_292/Y") V("POR2X1_152/A") V("POR2X1_173/Y") V("PAND2X1_784/A") V("PAND2X1_553/B") V("PAND2X1_633/Y") V("PAND2X1_640/B") V("POR2X1_813/Y") V("POR2X1_235/Y") V("POR2X1_624/B") V("POR2X1_711/B") V("POR2X1_713/A") V("PAND2X1_337/A") V("PAND2X1_778/Y") V("PAND2X1_198/Y") V("POR2X1_72/Y") V("POR2X1_184/Y") V("POR2X1_335/Y") V("POR2X1_784/A") V("POR2X1_208/A") V("POR2X1_202/A") V("PAND2X1_673/Y") V("POR2X1_65/Y") V("POR2X1_117/Y") V("POR2X1_262/Y") V("PAND2X1_632/A") V("PAND2X1_453/A") V("POR2X1_789/Y") V("PAND2X1_348/A") V("POR2X1_707/A") V("POR2X1_702/B") V("POR2X1_776/A") V("POR2X1_249/Y") V("POR2X1_401/A") V("POR2X1_507/A") V("PAND2X1_561/A") V("POR2X1_130/Y") V("POR2X1_156/B") V("POR2X1_231/A") V("POR2X1_636/A") V("POR2X1_247/Y") V("POR2X1_620/B") V("POR2X1_602/B") V("POR2X1_345/A") V("POR2X1_105/Y") V("POR2X1_756/Y") V("POR2X1_181/A") V("PAND2X1_535/Y") V("POR2X1_459/Y") V("PAND2X1_454/B") V("PAND2X1_506/Y") V("PAND2X1_852/A") V("PAND2X1_199/A") V("PAND2X1_139/B") V("POR2X1_132/Y") V("POR2X1_305/Y") V("POR2X1_384/A") V("POR2X1_766/Y") V("POR2X1_91/Y") V("POR2X1_312/Y") V("POR2X1_178/Y") V("POR2X1_67/Y") V("POR2X1_613/Y") V("POR2X1_647/B") V("POR2X1_670/Y") V("POR2X1_822/Y") V("POR2X1_420/Y") V("POR2X1_591/A") V("POR2X1_533/A") V("POR2X1_239/Y") V("POR2X1_172/Y") V("PAND2X1_843/Y") V("PAND2X1_287/Y") V("POR2X1_602/A") V("POR2X1_78/Y") V("POR2X1_240/B") V("POR2X1_446/A") V("POR2X1_608/Y") V("POR2X1_342/Y") V("POR2X1_486/B") V("POR2X1_546/B") V("POR2X1_507/B") V("POR2X1_720/A") V("POR2X1_546/A") V("POR2X1_848/Y") V("PAND2X1_303/B") V("PAND2X1_787/A") V("PAND2X1_552/B") V("PAND2X1_831/Y") V("PAND2X1_716/B") V("PAND2X1_392/B") V("POR2X1_823/Y") V("POR2X1_697/Y") V("POR2X1_759/Y") V("POR2X1_34/A") V("POR2X1_250/A") V("POR2X1_393/Y") V("PAND2X1_156/A") V("POR2X1_498/A") V("POR2X1_134/Y") V("POR2X1_679/B") V("POR2X1_754/A") V("POR2X1_427/Y") V("PAND2X1_638/B") V("PAND2X1_632/B") V("POR2X1_416/Y") V("POR2X1_481/Y") V("POR2X1_509/B") V("POR2X1_454/B") V("POR2X1_704/Y") V("POR2X1_333/Y") V("POR2X1_557/B") V("POR2X1_286/Y") V("POR2X1_370/Y") V("POR2X1_559/A") V("POR2X1_834/Y") V("POR2X1_783/B") V("POR2X1_196/Y") V("POR2X1_464/Y") V("POR2X1_828/Y") V("POR2X1_783/A") V("POR2X1_832/Y") V("POR2X1_841/B") V("POR2X1_156/Y") V("POR2X1_353/A") V("POR2X1_149/B") V("POR2X1_170/B") V("POR2X1_785/A") V("POR2X1_326/A") V("POR2X1_638/Y") V("POR2X1_712/A") V("PAND2X1_656/A") V("POR2X1_476/A") V("POR2X1_362/A") V("POR2X1_809/Y") V("PAND2X1_472/A") V("PAND2X1_243/B") V("PAND2X1_839/B") V("PAND2X1_338/B") V("POR2X1_676/Y") V("POR2X1_259/B") V("POR2X1_614/Y") V("POR2X1_545/A") V("POR2X1_445/A") V("PAND2X1_52/Y") V("POR2X1_636/B") V("POR2X1_523/B") V("POR2X1_782/B") V("POR2X1_836/B") V("POR2X1_779/A") V("POR2X1_542/B") V("POR2X1_635/B") V("POR2X1_710/A") V("POR2X1_792/B") V("POR2X1_383/Y") V("POR2X1_131/A") V("POR2X1_586/Y") V("POR2X1_516/Y") V("PAND2X1_793/A") V("POR2X1_248/A") V("POR2X1_423/Y") V("POR2X1_584/Y") V("POR2X1_7/Y") V("POR2X1_183/Y") V("POR2X1_33/B") V("POR2X1_344/Y") V("POR2X1_127/Y") V("POR2X1_698/Y") V("POR2X1_764/Y") V("POR2X1_380/Y") V("POR2X1_251/A") V("POR2X1_125/Y") V("POR2X1_442/Y") V("POR2X1_261/Y") V("POR2X1_757/A") V("POR2X1_561/B") V("POR2X1_112/Y") V("POR2X1_332/Y") V("POR2X1_550/A") V("POR2X1_729/Y") V("POR2X1_855/Y") V("POR2X1_574/A") V("POR2X1_503/Y") V("POR2X1_142/Y") V("POR2X1_518/Y") V("POR2X1_167/Y") V("POR2X1_667/Y") V("POR2X1_250/Y") V("POR2X1_829/Y") V("POR2X1_591/Y") V("POR2X1_321/Y") V("POR2X1_189/Y") V("POR2X1_96/Y") V("POR2X1_487/Y") V("POR2X1_406/Y") V("POR2X1_759/A") V("POR2X1_594/Y") V("POR2X1_533/Y") V("POR2X1_525/Y") V("POR2X1_163/Y") V("POR2X1_165/Y") V("POR2X1_145/Y") V("POR2X1_52/Y") V("POR2X1_680/Y") V("POR2X1_251/Y") V("POR2X1_418/Y") V("POR2X1_238/Y") V("POR2X1_462/B") V("POR2X1_259/A") V("POR2X1_781/A") V("POR2X1_181/B") V("POR2X1_210/B") V("POR2X1_719/A") V("POR2X1_499/A") V("POR2X1_435/B") V("POR2X1_646/B") V("PAND2X1_79/Y") V("POR2X1_833/A") V("POR2X1_194/A") V("POR2X1_790/A") V("POR2X1_324/B") V("POR2X1_148/A") V("PAND2X1_452/B") V("POR2X1_769/Y") V("POR2X1_635/Y") V("PAND2X1_460/Y") V("PAND2X1_197/Y") V("PAND2X1_308/B") V("POR2X1_554/B") V("POR2X1_342/A") V("POR2X1_400/A") V("POR2X1_209/A") V("POR2X1_113/B") V("POR2X1_705/B") V("POR2X1_347/B") V("POR2X1_449/A") V("POR2X1_780/A") V("POR2X1_791/A") V("POR2X1_403/B") V("POR2X1_124/B") V("POR2X1_493/B") V("POR2X1_775/A") V("POR2X1_302/B") V("POR2X1_76/B") V("POR2X1_227/B") V("POR2X1_559/B") V("POR2X1_97/A") V("POR2X1_343/A") V("POR2X1_506/B") V("POR2X1_210/A") V("POR2X1_168/A") V("POR2X1_148/B") V("POR2X1_728/A") V("PAND2X1_452/A") V("PAND2X1_707/Y") V("POR2X1_793/A") V("POR2X1_16/Y") V("POR2X1_665/Y") V("POR2X1_751/Y") V("POR2X1_767/Y") V("POR2X1_397/Y") V("POR2X1_504/Y") V("POR2X1_158/Y") V("POR2X1_232/Y") V("POR2X1_258/Y") V("POR2X1_746/Y") V("POR2X1_187/Y") V("POR2X1_166/Y") V("POR2X1_41/Y") V("POR2X1_441/Y") V("POR2X1_265/Y") V("POR2X1_745/Y") V("POR2X1_531/Y") V("POR2X1_384/Y") V("POR2X1_171/Y") V("POR2X1_177/Y") V("POR2X1_821/Y") V("POR2X1_118/Y") V("POR2X1_674/Y") V("POR2X1_498/Y") V("POR2X1_604/Y") V("POR2X1_438/Y") V("POR2X1_597/Y") V("PAND2X1_356/B") V("PAND2X1_389/Y") V("PAND2X1_711/A") V("PAND2X1_713/B") V("POR2X1_665/A") V("POR2X1_79/A") V("POR2X1_151/Y") V("POR2X1_188/Y") V("POR2X1_590/Y") V("POR2X1_777/Y") V("POR2X1_633/Y") V("POR2X1_553/A") V("POR2X1_243/B") V("POR2X1_664/Y") V("POR2X1_640/A") V("POR2X1_845/A") V("POR2X1_460/B") V("POR2X1_532/Y") V("PAND2X1_624/A") V("POR2X1_391/Y") V("POR2X1_565/B") V("POR2X1_673/Y") V("POR2X1_158/B") V("PAND2X1_783/B") V("POR2X1_829/A") V("PAND2X1_841/B") V("PAND2X1_459/Y") V("PAND2X1_651/A") V("PAND2X1_712/B") V("PAND2X1_308/Y") V("PAND2X1_149/A") V("PAND2X1_776/Y") V("PAND2X1_168/Y") V("PAND2X1_326/B") V("POR2X1_552/A") V("POR2X1_303/B") V("POR2X1_450/Y") V("POR2X1_302/Y") V("POR2X1_638/A") V("POR2X1_632/A") V("POR2X1_389/Y") V("POR2X1_632/B") V("PAND2X1_840/B") V("PAND2X1_779/Y") V("PAND2X1_769/Y") V("PAND2X1_199/B") V("PAND2X1_642/B") V("POR2X1_139/A") V("POR2X1_567/B") V("POR2X1_508/B") V("POR2X1_454/A") V("POR2X1_199/B") V("POR2X1_852/B") V("POR2X1_202/B") V("POR2X1_612/Y") V("PAND2X1_859/A") V("PAND2X1_340/B") V("PAND2X1_446/Y") V("PAND2X1_714/B") V("PAND2X1_333/Y") V("PAND2X1_557/A") V("PAND2X1_288/A") V("PAND2X1_464/Y") V("PAND2X1_349/A") V("POR2X1_850/A") V("POR2X1_288/A") V("POR2X1_609/A") V("POR2X1_669/Y") V("PAND2X1_332/Y") V("PAND2X1_115/B") V("PAND2X1_550/B") V("PAND2X1_856/B") V("PAND2X1_730/B") V("POR2X1_472/B") V("POR2X1_243/A") V("POR2X1_836/Y") V("POR2X1_334/Y") V("POR2X1_101/Y") V("PAND2X1_473/Y") V("PAND2X1_362/B") V("PAND2X1_810/B") V("PAND2X1_687/Y") V("POR2X1_687/Y") V("PAND2X1_254/Y") V("POR2X1_254/Y") V("PAND2X1_97/Y") V("POR2X1_802/B") V("POR2X1_802/A") V("POR2X1_99/B") V("PAND2X1_802/B") V("PAND2X1_798/Y") V("POR2X1_113/Y") V("POR2X1_319/Y") V("POR2X1_567/A") V("PAND2X1_114/B") V("PAND2X1_539/Y") V("PAND2X1_354/A") V("POR2X1_436/B") V("POR2X1_537/Y") V("POR2X1_592/Y") V("PAND2X1_592/Y") V("PAND2X1_643/A") V("PAND2X1_436/A") V("PAND2X1_593/Y") V("POR2X1_652/A") V("POR2X1_116/Y") V("POR2X1_88/Y") V("PAND2X1_717/A") V("POR2X1_761/A") V("POR2X1_373/Y") V("POR2X1_644/A") V("PAND2X1_216/B") V("POR2X1_717/B") V("PAND2X1_88/Y") V("POR2X1_483/B") V("POR2X1_544/B") V("POR2X1_252/Y") V("PAND2X1_267/Y") V("PAND2X1_631/A") V("PAND2X1_798/B") V("POR2X1_631/B") V("POR2X1_468/B") V("POR2X1_267/Y") 
    
    if ('showPlots' < 1)
        quit
    end
       
.endc

.end
