*** TEST 004 partitioning ***
*
* ngSPICE test for PLS experiments
*
* AES SBOX PLS test init file generator - protected dualRail SBOX area illuminated
*
* Author: Jan Belohoubek, 08/2020
* jan.belohoubek@fit.cvut.cz
*
* https://users.fit.cvut.cz/~belohja4/
*
*
* **************************************

.include ../../models.lib
.include ../../tsmc180nmcmos.lib
.include pDualRail.spice

* **************************************
* --- Test ---
* **************************************

* --- Settings
.param showPlots = 0
.param writeFile = 1
.param run_inputSet = 0

* redefine defaults ...
.include test00X_settings.inc

.csparam showPlots = {showPlots}
.csparam writeFile = {writeFile}
.csparam run_inputSet = {run_inputSet}

.global showPlots writeFile run_inputSet

* --- End of Settins

Vtrig LaserTrig 0 0 PWL(0ns 0V 20ns 0V 21ns SUPP)

.param beamDistanceTop = 0
.param beamDistanceBot = 0

.global LaserTrig beamDistanceTop beamDistanceBot

* --- inputs
Vvin0 INPUT_0 0 0 PWL(0ns 0V 5ns  0V 7ns  0V)
Vvin1 INPUT_1 0 0 PWL(0ns 0V 6ns  0V 8ns  0V)
Vvin2 INPUT_2 0 0 PWL(0ns 0V 7ns  0V 9ns  0V)
Vvin3 INPUT_3 0 0 PWL(0ns 0V 8ns  0V 10ns 0V)
Vvin4 INPUT_4 0 0 PWL(0ns 0V 9ns  0V 11ns 0V)
Vvin5 INPUT_5 0 0 PWL(0ns 0V 10ns 0V 12ns 0V)
Vvin6 INPUT_6 0 0 PWL(0ns 0V 11ns 0V 13ns 0V)
Vvin7 INPUT_7 0 0 PWL(0ns 0V 12ns 0V 14ns 0V)

Vvin0D D_INPUT_0 0 0 PWL(0ns 0V 5ns  0V 7ns  0V)
Vvin1D D_INPUT_1 0 0 PWL(0ns 0V 6ns  0V 8ns  0V)
Vvin2D D_INPUT_2 0 0 PWL(0ns 0V 7ns  0V 9ns  0V)
Vvin3D D_INPUT_3 0 0 PWL(0ns 0V 8ns  0V 10ns 0V)
Vvin4D D_INPUT_4 0 0 PWL(0ns 0V 9ns  0V 11ns 0V)
Vvin5D D_INPUT_5 0 0 PWL(0ns 0V 10ns 0V 12ns 0V)
Vvin6D D_INPUT_6 0 0 PWL(0ns 0V 11ns 0V 13ns 0V)
Vvin7D D_INPUT_7 0 0 PWL(0ns 0V 12ns 0V 14ns 0V)


* --- circuit layout model

Xsbox1 
+ POR2X1_452/A POR2X1_460/Y PAND2X1_635/Y POR2X1_152/Y POR2X1_612/B POR2X1_103/Y POR2X1_106/Y POR2X1_695/Y POR2X1_280/Y POR2X1_601/Y POR2X1_248/Y POR2X1_394/Y POR2X1_747/Y POR2X1_524/Y POR2X1_399/Y POR2X1_528/Y POR2X1_122/Y POR2X1_45/Y POR2X1_485/Y POR2X1_297/Y POR2X1_424/Y POR2X1_744/Y POR2X1_701/Y POR2X1_757/Y POR2X1_526/Y POR2X1_517/Y POR2X1_315/Y POR2X1_74/Y POR2X1_32/Y POR2X1_491/Y POR2X1_109/Y POR2X1_600/Y POR2X1_230/Y POR2X1_298/Y POR2X1_224/Y POR2X1_428/Y POR2X1_583/Y POR2X1_505/Y POR2X1_20/Y POR2X1_79/Y POR2X1_666/Y POR2X1_496/Y POR2X1_432/Y POR2X1_607/Y POR2X1_257/Y POR2X1_521/Y POR2X1_81/Y POR2X1_60/Y POR2X1_135/Y POR2X1_75/Y POR2X1_492/Y 
+ POR2X1_482/Y POR2X1_108/Y POR2X1_295/Y POR2X1_437/Y POR2X1_609/Y POR2X1_700/Y POR2X1_755/Y POR2X1_395/Y POR2X1_131/Y POR2X1_261/A POR2X1_679/A POR2X1_13/Y POR2X1_494/Y POR2X1_603/Y POR2X1_229/Y POR2X1_765/Y POR2X1_380/A POR2X1_707/Y POR2X1_307/Y POR2X1_197/Y POR2X1_379/Y POR2X1_334/B POR2X1_678/A POR2X1_84/A POR2X1_668/Y POR2X1_241/B POR2X1_34/B POR2X1_643/A POR2X1_538/A POR2X1_180/B POR2X1_844/B POR2X1_623/B POR2X1_33/A POR2X1_61/B POR2X1_523/A POR2X1_835/A POR2X1_709/B POR2X1_720/B POR2X1_343/B POR2X1_855/A POR2X1_832/B PAND2X1_65/Y POR2X1_593/B POR2X1_770/A POR2X1_324/A POR2X1_509/A POR2X1_703/A POR2X1_830/A POR2X1_520/B POR2X1_169/A PAND2X1_790/Y 
+ POR2X1_346/B POR2X1_443/A POR2X1_444/B POR2X1_620/A POR2X1_786/A POR2X1_267/B PAND2X1_41/Y POR2X1_610/Y POR2X1_769/A POR2X1_400/B POR2X1_781/B POR2X1_549/B POR2X1_391/A POR2X1_174/B POR2X1_540/A POR2X1_191/B POR2X1_169/B POR2X1_758/Y POR2X1_673/B POR2X1_835/B POR2X1_123/B POR2X1_123/A POR2X1_675/A POR2X1_501/B PAND2X1_72/Y POR2X1_605/A POR2X1_450/A POR2X1_544/A POR2X1_637/A POR2X1_174/A POR2X1_175/B POR2X1_180/A POR2X1_128/A POR2X1_555/A PAND2X1_7/Y POR2X1_719/B POR2X1_789/A POR2X1_194/B POR2X1_773/B POR2X1_402/B POR2X1_307/A POR2X1_311/Y POR2X1_176/Y POR2X1_83/Y POR2X1_669/A POR2X1_290/Y POR2X1_27/Y POR2X1_677/Y POR2X1_237/Y POR2X1_595/Y POR2X1_146/Y 
+ POR2X1_179/Y POR2X1_69/Y POR2X1_484/Y POR2X1_495/Y POR2X1_39/Y POR2X1_754/Y POR2X1_396/Y POR2X1_320/Y POR2X1_24/Y POR2X1_58/Y POR2X1_497/Y POR2X1_615/Y POR2X1_522/Y POR2X1_493/A POR2X1_483/A POR2X1_114/B POR2X1_84/B POR2X1_346/A POR2X1_61/A POR2X1_76/A POR2X1_440/B POR2X1_646/A POR2X1_710/B POR2X1_791/B POR2X1_401/B POR2X1_702/A POR2X1_558/A POR2X1_605/B POR2X1_260/Y POR2X1_678/Y POR2X1_193/A POR2X1_231/B POR2X1_770/B POR2X1_140/A POR2X1_447/A POR2X1_489/B POR2X1_98/A POR2X1_734/B POR2X1_653/B POR2X1_788/B POR2X1_456/B POR2X1_137/B POR2X1_768/A POR2X1_192/B POR2X1_128/B POR2X1_644/B POR2X1_448/Y POR2X1_356/A PAND2X1_565/A POR2X1_292/Y POR2X1_152/A 
+ POR2X1_173/Y PAND2X1_784/A PAND2X1_553/B PAND2X1_633/Y PAND2X1_640/B POR2X1_813/Y POR2X1_235/Y POR2X1_624/B POR2X1_711/B POR2X1_713/A PAND2X1_337/A PAND2X1_778/Y PAND2X1_198/Y POR2X1_72/Y POR2X1_184/Y POR2X1_335/Y POR2X1_784/A POR2X1_208/A POR2X1_202/A PAND2X1_673/Y POR2X1_65/Y POR2X1_117/Y POR2X1_262/Y PAND2X1_632/A PAND2X1_453/A POR2X1_789/Y PAND2X1_348/A POR2X1_707/A POR2X1_702/B POR2X1_776/A POR2X1_249/Y POR2X1_401/A POR2X1_507/A PAND2X1_561/A POR2X1_130/Y POR2X1_156/B POR2X1_231/A POR2X1_636/A POR2X1_247/Y POR2X1_620/B POR2X1_602/B POR2X1_345/A POR2X1_105/Y POR2X1_756/Y POR2X1_181/A PAND2X1_535/Y POR2X1_459/Y PAND2X1_454/B PAND2X1_506/Y PAND2X1_852/A PAND2X1_199/A 
+ PAND2X1_139/B POR2X1_132/Y POR2X1_305/Y POR2X1_384/A POR2X1_766/Y POR2X1_91/Y POR2X1_312/Y POR2X1_178/Y POR2X1_67/Y POR2X1_613/Y POR2X1_647/B POR2X1_670/Y POR2X1_822/Y POR2X1_420/Y POR2X1_591/A POR2X1_533/A POR2X1_239/Y POR2X1_172/Y PAND2X1_843/Y PAND2X1_287/Y POR2X1_602/A POR2X1_78/Y POR2X1_240/B POR2X1_446/A POR2X1_608/Y POR2X1_342/Y POR2X1_486/B POR2X1_546/B POR2X1_507/B POR2X1_720/A POR2X1_546/A POR2X1_848/Y PAND2X1_303/B PAND2X1_787/A PAND2X1_552/B PAND2X1_831/Y PAND2X1_716/B PAND2X1_392/B POR2X1_823/Y POR2X1_697/Y POR2X1_759/Y POR2X1_34/A POR2X1_250/A POR2X1_393/Y PAND2X1_156/A POR2X1_498/A POR2X1_134/Y POR2X1_679/B POR2X1_754/A POR2X1_427/Y PAND2X1_638/B 
+ PAND2X1_632/B POR2X1_416/Y POR2X1_481/Y POR2X1_509/B POR2X1_454/B POR2X1_704/Y POR2X1_333/Y POR2X1_557/B POR2X1_286/Y POR2X1_370/Y POR2X1_559/A POR2X1_834/Y POR2X1_783/B POR2X1_196/Y POR2X1_464/Y POR2X1_828/Y POR2X1_783/A POR2X1_832/Y POR2X1_841/B POR2X1_156/Y POR2X1_353/A POR2X1_149/B POR2X1_170/B POR2X1_785/A POR2X1_326/A POR2X1_638/Y POR2X1_712/A PAND2X1_656/A POR2X1_476/A POR2X1_362/A POR2X1_809/Y PAND2X1_472/A PAND2X1_243/B PAND2X1_839/B PAND2X1_338/B POR2X1_676/Y POR2X1_259/B POR2X1_614/Y POR2X1_545/A POR2X1_445/A PAND2X1_52/Y POR2X1_636/B POR2X1_523/B POR2X1_782/B POR2X1_836/B POR2X1_779/A POR2X1_542/B POR2X1_635/B POR2X1_710/A POR2X1_792/B POR2X1_383/Y 
+ POR2X1_131/A POR2X1_586/Y POR2X1_516/Y PAND2X1_793/A POR2X1_248/A POR2X1_423/Y POR2X1_584/Y POR2X1_7/Y POR2X1_183/Y POR2X1_33/B POR2X1_344/Y POR2X1_127/Y POR2X1_698/Y POR2X1_764/Y POR2X1_380/Y POR2X1_251/A POR2X1_125/Y POR2X1_442/Y POR2X1_261/Y POR2X1_757/A POR2X1_561/B POR2X1_112/Y POR2X1_332/Y POR2X1_550/A POR2X1_729/Y POR2X1_855/Y POR2X1_574/A POR2X1_503/Y POR2X1_142/Y POR2X1_518/Y POR2X1_167/Y POR2X1_667/Y POR2X1_250/Y POR2X1_829/Y POR2X1_591/Y POR2X1_321/Y POR2X1_189/Y POR2X1_96/Y POR2X1_487/Y POR2X1_406/Y POR2X1_759/A POR2X1_594/Y POR2X1_533/Y POR2X1_525/Y POR2X1_163/Y POR2X1_165/Y POR2X1_145/Y POR2X1_52/Y POR2X1_680/Y POR2X1_251/Y POR2X1_418/Y 
+ POR2X1_238/Y POR2X1_462/B POR2X1_259/A POR2X1_781/A POR2X1_181/B POR2X1_210/B POR2X1_719/A POR2X1_499/A POR2X1_435/B POR2X1_646/B PAND2X1_79/Y POR2X1_833/A POR2X1_194/A POR2X1_790/A POR2X1_324/B POR2X1_148/A PAND2X1_452/B POR2X1_769/Y POR2X1_635/Y PAND2X1_460/Y PAND2X1_197/Y PAND2X1_308/B POR2X1_554/B POR2X1_342/A POR2X1_400/A POR2X1_209/A POR2X1_113/B POR2X1_705/B POR2X1_347/B POR2X1_449/A POR2X1_780/A POR2X1_791/A POR2X1_403/B POR2X1_124/B POR2X1_493/B POR2X1_775/A POR2X1_302/B POR2X1_76/B POR2X1_227/B POR2X1_559/B POR2X1_97/A POR2X1_343/A POR2X1_506/B POR2X1_210/A POR2X1_168/A POR2X1_148/B POR2X1_728/A PAND2X1_452/A PAND2X1_707/Y POR2X1_793/A POR2X1_16/Y 
+ POR2X1_665/Y POR2X1_751/Y POR2X1_767/Y POR2X1_397/Y POR2X1_504/Y POR2X1_158/Y POR2X1_232/Y POR2X1_258/Y POR2X1_746/Y POR2X1_187/Y POR2X1_166/Y POR2X1_41/Y POR2X1_441/Y POR2X1_265/Y POR2X1_745/Y POR2X1_531/Y POR2X1_384/Y POR2X1_171/Y POR2X1_177/Y POR2X1_821/Y POR2X1_118/Y POR2X1_674/Y POR2X1_498/Y POR2X1_604/Y POR2X1_438/Y POR2X1_597/Y PAND2X1_356/B PAND2X1_389/Y PAND2X1_711/A PAND2X1_713/B POR2X1_665/A POR2X1_79/A POR2X1_151/Y POR2X1_188/Y POR2X1_590/Y POR2X1_777/Y POR2X1_633/Y POR2X1_553/A POR2X1_243/B POR2X1_664/Y POR2X1_640/A POR2X1_845/A POR2X1_460/B POR2X1_532/Y PAND2X1_624/A POR2X1_391/Y POR2X1_565/B POR2X1_673/Y POR2X1_158/B PAND2X1_783/B POR2X1_829/A 
+ PAND2X1_841/B PAND2X1_459/Y PAND2X1_651/A PAND2X1_712/B PAND2X1_308/Y PAND2X1_149/A PAND2X1_776/Y PAND2X1_168/Y PAND2X1_326/B POR2X1_552/A POR2X1_303/B POR2X1_450/Y POR2X1_302/Y POR2X1_638/A POR2X1_632/A POR2X1_389/Y POR2X1_632/B PAND2X1_840/B PAND2X1_779/Y PAND2X1_769/Y PAND2X1_199/B PAND2X1_642/B POR2X1_139/A POR2X1_567/B POR2X1_508/B POR2X1_454/A POR2X1_199/B POR2X1_852/B POR2X1_202/B POR2X1_612/Y PAND2X1_859/A PAND2X1_340/B PAND2X1_446/Y PAND2X1_714/B PAND2X1_333/Y PAND2X1_557/A PAND2X1_288/A PAND2X1_464/Y PAND2X1_349/A POR2X1_850/A POR2X1_288/A POR2X1_609/A POR2X1_669/Y PAND2X1_332/Y PAND2X1_115/B PAND2X1_550/B PAND2X1_856/B PAND2X1_730/B POR2X1_472/B POR2X1_243/A POR2X1_836/Y 
+ POR2X1_334/Y POR2X1_101/Y PAND2X1_473/Y PAND2X1_362/B PAND2X1_810/B PAND2X1_687/Y POR2X1_687/Y PAND2X1_254/Y POR2X1_254/Y PAND2X1_97/Y POR2X1_802/B POR2X1_802/A POR2X1_99/B PAND2X1_802/B PAND2X1_798/Y POR2X1_113/Y POR2X1_319/Y POR2X1_567/A PAND2X1_114/B PAND2X1_539/Y PAND2X1_354/A POR2X1_436/B POR2X1_537/Y POR2X1_592/Y PAND2X1_592/Y PAND2X1_643/A PAND2X1_436/A PAND2X1_593/Y POR2X1_652/A POR2X1_116/Y POR2X1_88/Y PAND2X1_717/A POR2X1_761/A POR2X1_373/Y POR2X1_644/A PAND2X1_216/B POR2X1_717/B PAND2X1_88/Y POR2X1_483/B POR2X1_544/B POR2X1_252/Y PAND2X1_267/Y PAND2X1_631/A PAND2X1_798/B POR2X1_631/B POR2X1_468/B POR2X1_267/Y 
+ VSS VDD 
+ PAND2X1_812/A PAND2X1_366/A PAND2X1_479/B POR2X1_660/A POR2X1_216/Y POR2X1_351/B POR2X1_852/A POR2X1_243/Y POR2X1_472/Y PAND2X1_739/B PAND2X1_863/A PAND2X1_550/Y PAND2X1_724/B PAND2X1_339/Y PAND2X1_721/B POR2X1_362/B POR2X1_858/B PAND2X1_359/B PAND2X1_477/B PAND2X1_362/A PAND2X1_773/B PAND2X1_351/A PAND2X1_714/Y PAND2X1_466/B PAND2X1_350/A PAND2X1_862/B PAND2X1_656/B POR2X1_206/A POR2X1_857/B POR2X1_207/B POR2X1_466/A POR2X1_856/B POR2X1_568/A POR2X1_139/Y PAND2X1_649/A PAND2X1_560/B PAND2X1_207/A PAND2X1_783/Y PAND2X1_840/Y POR2X1_632/Y POR2X1_392/B POR2X1_566/A POR2X1_452/Y POR2X1_723/B POR2X1_552/Y PAND2X1_717/Y PAND2X1_211/A PAND2X1_785/Y PAND2X1_209/A PAND2X1_353/Y PAND2X1_731/B 
+ PAND2X1_725/A PAND2X1_651/Y PAND2X1_472/B PAND2X1_841/Y POR2X1_734/A POR2X1_569/A POR2X1_860/A PAND2X1_658/A POR2X1_640/Y POR2X1_553/Y POR2X1_796/A PAND2X1_725/B PAND2X1_726/B PAND2X1_390/Y PAND2X1_365/A PAND2X1_644/Y PAND2X1_675/A PAND2X1_551/A PAND2X1_645/B PAND2X1_573/B PAND2X1_736/A PAND2X1_123/Y PAND2X1_835/Y PAND2X1_182/A PAND2X1_175/B PAND2X1_781/Y PAND2X1_641/Y PAND2X1_443/Y PAND2X1_545/Y PAND2X1_169/Y PAND2X1_191/Y PAND2X1_555/A PAND2X1_213/B PAND2X1_508/B PAND2X1_719/Y PAND2X1_200/B POR2X1_805/A PAND2X1_467/B POR2X1_730/B POR2X1_149/A POR2X1_467/Y POR2X1_210/Y POR2X1_244/B POR2X1_343/Y POR2X1_444/A POR2X1_785/B POR2X1_559/Y POR2X1_558/B POR2X1_572/B POR2X1_791/Y POR2X1_449/Y 
+ POR2X1_360/A POR2X1_556/A POR2X1_713/B POR2X1_768/Y POR2X1_213/B POR2X1_726/Y POR2X1_403/A POR2X1_554/Y POR2X1_639/Y POR2X1_324/Y POR2X1_644/Y POR2X1_200/A POR2X1_840/B POR2X1_500/A POR2X1_205/A POR2X1_646/Y POR2X1_722/A POR2X1_540/Y POR2X1_181/Y POR2X1_782/A POR2X1_555/B POR2X1_649/B PAND2X1_241/Y PAND2X1_349/B PAND2X1_730/A PAND2X1_341/A PAND2X1_148/Y PAND2X1_467/Y PAND2X1_546/Y PAND2X1_794/B PAND2X1_653/Y PAND2X1_479/A PAND2X1_737/B PAND2X1_192/Y PAND2X1_324/Y PAND2X1_718/Y PAND2X1_714/A PAND2X1_388/Y PAND2X1_830/Y POR2X1_574/Y POR2X1_863/B POR2X1_730/Y POR2X1_550/Y POR2X1_339/Y POR2X1_724/A POR2X1_561/Y PAND2X1_345/Y PAND2X1_444/Y PAND2X1_140/A POR2X1_359/B PAND2X1_553/A 
+ PAND2X1_190/Y PAND2X1_193/Y PAND2X1_639/B PAND2X1_449/Y PAND2X1_793/Y PAND2X1_575/B POR2X1_805/B POR2X1_710/Y POR2X1_542/Y POR2X1_797/A POR2X1_523/Y POR2X1_639/A POR2X1_228/Y POR2X1_551/A POR2X1_728/B PAND2X1_852/B PAND2X1_244/B PAND2X1_476/A POR2X1_812/B POR2X1_362/Y POR2X1_476/Y PAND2X1_660/B PAND2X1_218/A POR2X1_712/Y POR2X1_651/Y POR2X1_717/Y POR2X1_795/B POR2X1_566/B POR2X1_149/Y POR2X1_353/Y POR2X1_731/A POR2X1_851/A POR2X1_783/Y POR2X1_477/A POR2X1_840/Y POR2X1_794/B POR2X1_773/A POR2X1_724/B POR2X1_350/B PAND2X1_555/Y PAND2X1_658/B POR2X1_679/Y PAND2X1_137/Y PAND2X1_768/Y PAND2X1_403/B PAND2X1_805/A PAND2X1_474/A PAND2X1_723/A PAND2X1_303/Y PAND2X1_564/B PAND2X1_787/Y 
+ POR2X1_862/A POR2X1_550/B POR2X1_720/Y POR2X1_508/A POR2X1_349/Y POR2X1_788/A PAND2X1_850/Y PAND2X1_242/Y POR2X1_647/Y PAND2X1_620/Y PAND2X1_206/B PAND2X1_182/B PAND2X1_552/A PAND2X1_336/Y PAND2X1_785/A PAND2X1_771/B PAND2X1_139/Y PAND2X1_857/A POR2X1_463/Y PAND2X1_854/Y PAND2X1_568/B POR2X1_348/A POR2X1_623/A POR2X1_341/A PAND2X1_561/Y POR2X1_402/A POR2X1_241/Y POR2X1_715/A PAND2X1_348/Y PAND2X1_466/A PAND2X1_795/B PAND2X1_206/A PAND2X1_734/B POR2X1_208/Y POR2X1_337/Y PAND2X1_842/Y PAND2X1_205/A PAND2X1_214/B PAND2X1_796/B PAND2X1_352/B POR2X1_713/Y POR2X1_711/Y POR2X1_624/Y PAND2X1_650/A PAND2X1_563/A PAND2X1_853/B PAND2X1_346/Y PAND2X1_569/B POR2X1_356/Y POR2X1_453/Y POR2X1_140/B 
+ POR2X1_192/Y POR2X1_137/Y POR2X1_850/B POR2X1_190/Y POR2X1_788/Y POR2X1_661/B POR2X1_479/B POR2X1_737/A POR2X1_141/A POR2X1_771/A POR2X1_193/Y POR2X1_718/A POR2X1_558/Y POR2X1_440/Y POR2X1_61/Y POR2X1_347/A POR2X1_84/Y POR2X1_830/Y PAND2X1_844/B PAND2X1_623/Y PAND2X1_501/B PAND2X1_61/Y PAND2X1_402/B PAND2X1_840/A PAND2X1_499/Y PAND2X1_556/B PAND2X1_643/Y PAND2X1_84/Y POR2X1_562/B POR2X1_439/Y POR2X1_180/Y POR2X1_853/A POR2X1_175/A POR2X1_544/Y POR2X1_203/Y POR2X1_573/A POR2X1_675/Y POR2X1_123/Y POR2X1_835/Y POR2X1_169/Y POR2X1_191/Y POR2X1_650/A POR2X1_786/Y POR2X1_444/Y POR2X1_390/B POR2X1_703/Y POR2X1_337/A POR2X1_722/B POR2X1_201/Y POR2X1_623/Y POR2X1_500/Y 
+ POR2X1_643/Y PAND2X1_341/B PAND2X1_558/Y PAND2X1_140/Y PAND2X1_792/B PAND2X1_711/B PAND2X1_647/B PAND2X1_652/A PAND2X1_493/Y PAND2X1_715/B PAND2X1_205/B PAND2X1_602/Y PAND2X1_713/A PAND2X1_347/Y PAND2X1_124/Y PAND2X1_782/Y PAND2X1_563/B PAND2X1_213/A PAND2X1_731/A PAND2X1_639/Y POR2X1_802/B POR2X1_802/A PAND2X1_802/B PAND2X1_798/Y POR2X1_567/A PAND2X1_539/Y PAND2X1_810/A POR2X1_510/Y PAND2X1_657/B POR2X1_774/Y POR2X1_35/Y PAND2X1_35/Y PAND2X1_455/Y PAND2X1_404/Y POR2X1_465/B POR2X1_404/Y PAND2X1_267/Y PAND2X1_631/A PAND2X1_798/B POR2X1_652/A POR2X1_631/B POR2X1_468/B POR2X1_319/Y PAND2X1_593/Y POR2X1_267/Y PAND2X1_354/A 
+ AES_SBOX_2

.include outputs_1.plw

* **************************************
* --- Simulation Settings ---
* **************************************

.param SIM_LEN = 35ns
.csparam SIM_LEN = {SIM_LEN}

*.options abstol=0.000001 vntol=0.001 reltol=0.01

.tran 1ns 'SIM_LEN'
.param SIMSTEP = 'SIM_LEN/1ns'
.csparam SIMSTEP = {SIMSTEP}

* **************************************
* --- Simulation Control ---
* **************************************

.control
    .include ../inputsD.inc

    *stop when time = 8.500ns
    run
    
    if ('writeFile' > 0)   
      wrdata ivdd_2.out i(vvdd)
      wrdata ivss_2.out i(vvss)
      *snsave sim_2.snap
    end
    
    set wr_vecnames
    set wr_singlescale
    wrdata outputs_2.out V("PAND2X1_812/A") V("PAND2X1_366/A") V("PAND2X1_479/B") V("POR2X1_660/A") V("POR2X1_216/Y") V("POR2X1_351/B") V("POR2X1_852/A") V("POR2X1_243/Y") V("POR2X1_472/Y") V("PAND2X1_739/B") V("PAND2X1_863/A") V("PAND2X1_550/Y") V("PAND2X1_724/B") V("PAND2X1_339/Y") V("PAND2X1_721/B") V("POR2X1_362/B") V("POR2X1_858/B") V("PAND2X1_359/B") V("PAND2X1_477/B") V("PAND2X1_362/A") V("PAND2X1_773/B") V("PAND2X1_351/A") V("PAND2X1_714/Y") V("PAND2X1_466/B") V("PAND2X1_350/A") V("PAND2X1_862/B") V("PAND2X1_656/B") V("POR2X1_206/A") V("POR2X1_857/B") V("POR2X1_207/B") V("POR2X1_466/A") V("POR2X1_856/B") V("POR2X1_568/A") V("POR2X1_139/Y") V("PAND2X1_649/A") V("PAND2X1_560/B") V("PAND2X1_207/A") V("PAND2X1_783/Y") V("PAND2X1_840/Y") V("POR2X1_632/Y") V("POR2X1_392/B") V("POR2X1_566/A") V("POR2X1_452/Y") V("POR2X1_723/B") V("POR2X1_552/Y") V("PAND2X1_717/Y") V("PAND2X1_211/A") V("PAND2X1_785/Y") V("PAND2X1_209/A") V("PAND2X1_353/Y") V("PAND2X1_731/B") V("PAND2X1_725/A") V("PAND2X1_651/Y") V("PAND2X1_472/B") V("PAND2X1_841/Y") V("POR2X1_734/A") V("POR2X1_569/A") V("POR2X1_860/A") V("PAND2X1_658/A") V("POR2X1_640/Y") V("POR2X1_553/Y") V("POR2X1_796/A") V("PAND2X1_725/B") V("PAND2X1_726/B") V("PAND2X1_390/Y") V("PAND2X1_365/A") V("PAND2X1_644/Y") V("PAND2X1_675/A") V("PAND2X1_551/A") V("PAND2X1_645/B") V("PAND2X1_573/B") V("PAND2X1_736/A") V("PAND2X1_123/Y") V("PAND2X1_835/Y") V("PAND2X1_182/A") V("PAND2X1_175/B") V("PAND2X1_781/Y") V("PAND2X1_641/Y") V("PAND2X1_443/Y") V("PAND2X1_545/Y") V("PAND2X1_169/Y") V("PAND2X1_191/Y") V("PAND2X1_555/A") V("PAND2X1_213/B") V("PAND2X1_508/B") V("PAND2X1_719/Y") V("PAND2X1_200/B") V("POR2X1_805/A") V("PAND2X1_467/B") V("POR2X1_730/B") V("POR2X1_149/A") V("POR2X1_467/Y") V("POR2X1_210/Y") V("POR2X1_244/B") V("POR2X1_343/Y") V("POR2X1_444/A") V("POR2X1_785/B") V("POR2X1_559/Y") V("POR2X1_558/B") V("POR2X1_572/B") V("POR2X1_791/Y") V("POR2X1_449/Y") V("POR2X1_360/A") V("POR2X1_556/A") V("POR2X1_713/B") V("POR2X1_768/Y") V("POR2X1_213/B") V("POR2X1_726/Y") V("POR2X1_403/A") V("POR2X1_554/Y") V("POR2X1_639/Y") V("POR2X1_324/Y") V("POR2X1_644/Y") V("POR2X1_200/A") V("POR2X1_840/B") V("POR2X1_500/A") V("POR2X1_205/A") V("POR2X1_646/Y") V("POR2X1_722/A") V("POR2X1_540/Y") V("POR2X1_181/Y") V("POR2X1_782/A") V("POR2X1_555/B") V("POR2X1_649/B") V("PAND2X1_241/Y") V("PAND2X1_349/B") V("PAND2X1_730/A") V("PAND2X1_341/A") V("PAND2X1_148/Y") V("PAND2X1_467/Y") V("PAND2X1_546/Y") V("PAND2X1_794/B") V("PAND2X1_653/Y") V("PAND2X1_479/A") V("PAND2X1_737/B") V("PAND2X1_192/Y") V("PAND2X1_324/Y") V("PAND2X1_718/Y") V("PAND2X1_714/A") V("PAND2X1_388/Y") V("PAND2X1_830/Y") V("POR2X1_574/Y") V("POR2X1_863/B") V("POR2X1_730/Y") V("POR2X1_550/Y") V("POR2X1_339/Y") V("POR2X1_724/A") V("POR2X1_561/Y") V("PAND2X1_345/Y") V("PAND2X1_444/Y") V("PAND2X1_140/A") V("POR2X1_359/B") V("PAND2X1_553/A") V("PAND2X1_190/Y") V("PAND2X1_193/Y") V("PAND2X1_639/B") V("PAND2X1_449/Y") V("PAND2X1_793/Y") V("PAND2X1_575/B") V("POR2X1_805/B") V("POR2X1_710/Y") V("POR2X1_542/Y") V("POR2X1_797/A") V("POR2X1_523/Y") V("POR2X1_639/A") V("POR2X1_228/Y") V("POR2X1_551/A") V("POR2X1_728/B") V("PAND2X1_852/B") V("PAND2X1_244/B") V("PAND2X1_476/A") V("POR2X1_812/B") V("POR2X1_362/Y") V("POR2X1_476/Y") V("PAND2X1_660/B") V("PAND2X1_218/A") V("POR2X1_712/Y") V("POR2X1_651/Y") V("POR2X1_717/Y") V("POR2X1_795/B") V("POR2X1_566/B") V("POR2X1_149/Y") V("POR2X1_353/Y") V("POR2X1_731/A") V("POR2X1_851/A") V("POR2X1_783/Y") V("POR2X1_477/A") V("POR2X1_840/Y") V("POR2X1_794/B") V("POR2X1_773/A") V("POR2X1_724/B") V("POR2X1_350/B") V("PAND2X1_555/Y") V("PAND2X1_658/B") V("POR2X1_679/Y") V("PAND2X1_137/Y") V("PAND2X1_768/Y") V("PAND2X1_403/B") V("PAND2X1_805/A") V("PAND2X1_474/A") V("PAND2X1_723/A") V("PAND2X1_303/Y") V("PAND2X1_564/B") V("PAND2X1_787/Y") V("POR2X1_862/A") V("POR2X1_550/B") V("POR2X1_720/Y") V("POR2X1_508/A") V("POR2X1_349/Y") V("POR2X1_788/A") V("PAND2X1_850/Y") V("PAND2X1_242/Y") V("POR2X1_647/Y") V("PAND2X1_620/Y") V("PAND2X1_206/B") V("PAND2X1_182/B") V("PAND2X1_552/A") V("PAND2X1_336/Y") V("PAND2X1_785/A") V("PAND2X1_771/B") V("PAND2X1_139/Y") V("PAND2X1_857/A") V("POR2X1_463/Y") V("PAND2X1_854/Y") V("PAND2X1_568/B") V("POR2X1_348/A") V("POR2X1_623/A") V("POR2X1_341/A") V("PAND2X1_561/Y") V("POR2X1_402/A") V("POR2X1_241/Y") V("POR2X1_715/A") V("PAND2X1_348/Y") V("PAND2X1_466/A") V("PAND2X1_795/B") V("PAND2X1_206/A") V("PAND2X1_734/B") V("POR2X1_208/Y") V("POR2X1_337/Y") V("PAND2X1_842/Y") V("PAND2X1_205/A") V("PAND2X1_214/B") V("PAND2X1_796/B") V("PAND2X1_352/B") V("POR2X1_713/Y") V("POR2X1_711/Y") V("POR2X1_624/Y") V("PAND2X1_650/A") V("PAND2X1_563/A") V("PAND2X1_853/B") V("PAND2X1_346/Y") V("PAND2X1_569/B") V("POR2X1_356/Y") V("POR2X1_453/Y") V("POR2X1_140/B") V("POR2X1_192/Y") V("POR2X1_137/Y") V("POR2X1_850/B") V("POR2X1_190/Y") V("POR2X1_788/Y") V("POR2X1_661/B") V("POR2X1_479/B") V("POR2X1_737/A") V("POR2X1_141/A") V("POR2X1_771/A") V("POR2X1_193/Y") V("POR2X1_718/A") V("POR2X1_558/Y") V("POR2X1_440/Y") V("POR2X1_61/Y") V("POR2X1_347/A") V("POR2X1_84/Y") V("POR2X1_830/Y") V("PAND2X1_844/B") V("PAND2X1_623/Y") V("PAND2X1_501/B") V("PAND2X1_61/Y") V("PAND2X1_402/B") V("PAND2X1_840/A") V("PAND2X1_499/Y") V("PAND2X1_556/B") V("PAND2X1_643/Y") V("PAND2X1_84/Y") V("POR2X1_562/B") V("POR2X1_439/Y") V("POR2X1_180/Y") V("POR2X1_853/A") V("POR2X1_175/A") V("POR2X1_544/Y") V("POR2X1_203/Y") V("POR2X1_573/A") V("POR2X1_675/Y") V("POR2X1_123/Y") V("POR2X1_835/Y") V("POR2X1_169/Y") V("POR2X1_191/Y") V("POR2X1_650/A") V("POR2X1_786/Y") V("POR2X1_444/Y") V("POR2X1_390/B") V("POR2X1_703/Y") V("POR2X1_337/A") V("POR2X1_722/B") V("POR2X1_201/Y") V("POR2X1_623/Y") V("POR2X1_500/Y") V("POR2X1_643/Y") V("PAND2X1_341/B") V("PAND2X1_558/Y") V("PAND2X1_140/Y") V("PAND2X1_792/B") V("PAND2X1_711/B") V("PAND2X1_647/B") V("PAND2X1_652/A") V("PAND2X1_493/Y") V("PAND2X1_715/B") V("PAND2X1_205/B") V("PAND2X1_602/Y") V("PAND2X1_713/A") V("PAND2X1_347/Y") V("PAND2X1_124/Y") V("PAND2X1_782/Y") V("PAND2X1_563/B") V("PAND2X1_213/A") V("PAND2X1_731/A") V("PAND2X1_639/Y") V("POR2X1_802/B") V("POR2X1_802/A") V("PAND2X1_802/B") V("PAND2X1_798/Y") V("POR2X1_567/A") V("PAND2X1_539/Y") V("PAND2X1_810/A") V("POR2X1_510/Y") V("PAND2X1_657/B") V("POR2X1_774/Y") V("POR2X1_35/Y") V("PAND2X1_35/Y") V("PAND2X1_455/Y") V("PAND2X1_404/Y") V("POR2X1_465/B") V("POR2X1_404/Y") V("PAND2X1_267/Y") V("PAND2X1_631/A") V("PAND2X1_798/B") V("POR2X1_652/A") V("POR2X1_631/B") V("POR2X1_468/B") V("POR2X1_319/Y") V("PAND2X1_593/Y") V("POR2X1_267/Y") V("PAND2X1_354/A") 
    
    if ('showPlots' < 1)
        quit
    end
       
.endc

.end
