*** TEST 005 partitioning ***
*
* ngSPICE test for PLS experiments
*
* AES SBOX PLS test init file generator - protected dualRail SBOX area illuminated
*
* Author: Jan Belohoubek, 08/2020
* jan.belohoubek@fit.cvut.cz
*
* https://users.fit.cvut.cz/~belohja4/
*
*
* **************************************

.include ../../models.lib
.include ../../tsmc180nmcmos.lib
.include secLibDualRail.spice

* **************************************
* --- Test ---
* **************************************

* --- Settings
.param showPlots = 0
.param writeFile = 1
.param run_inputSet = 0

* redefine defaults ...
.include test00X_settings.inc

.csparam showPlots = {showPlots}
.csparam writeFile = {writeFile}
.csparam run_inputSet = {run_inputSet}

.global showPlots writeFile run_inputSet

* --- End of Settins

Vtrig LaserTrig 0 0 PWL(0ns 0V 40ns 0V 41ns SUPP)

.param beamDistanceTop = 0
.param beamDistanceBot = 0

.global LaserTrig beamDistanceTop beamDistanceBot

* --- inputs
Vvin0 INPUT_0 0 0 PWL(0ns 0V 5ns  0V 7ns  0V)
Vvin1 INPUT_1 0 0 PWL(0ns 0V 6ns  0V 8ns  0V)
Vvin2 INPUT_2 0 0 PWL(0ns 0V 7ns  0V 9ns  0V)
Vvin3 INPUT_3 0 0 PWL(0ns 0V 8ns  0V 10ns 0V)
Vvin4 INPUT_4 0 0 PWL(0ns 0V 9ns  0V 11ns 0V)
Vvin5 INPUT_5 0 0 PWL(0ns 0V 10ns 0V 12ns 0V)
Vvin6 INPUT_6 0 0 PWL(0ns 0V 11ns 0V 13ns 0V)
Vvin7 INPUT_7 0 0 PWL(0ns 0V 12ns 0V 14ns 0V)

Vvin0D D_INPUT_0 0 0 PWL(0ns 0V 5ns  0V 7ns  0V)
Vvin1D D_INPUT_1 0 0 PWL(0ns 0V 6ns  0V 8ns  0V)
Vvin2D D_INPUT_2 0 0 PWL(0ns 0V 7ns  0V 9ns  0V)
Vvin3D D_INPUT_3 0 0 PWL(0ns 0V 8ns  0V 10ns 0V)
Vvin4D D_INPUT_4 0 0 PWL(0ns 0V 9ns  0V 11ns 0V)
Vvin5D D_INPUT_5 0 0 PWL(0ns 0V 10ns 0V 12ns 0V)
Vvin6D D_INPUT_6 0 0 PWL(0ns 0V 11ns 0V 13ns 0V)
Vvin7D D_INPUT_7 0 0 PWL(0ns 0V 12ns 0V 14ns 0V)


* --- circuit layout model

Xsbox1 
+ INPUT_0 INPUT_1 INPUT_2 INPUT_3 INPUT_4 INPUT_5 INPUT_6 INPUT_7 D_INPUT_0 D_INPUT_1 D_INPUT_2 D_INPUT_3 D_INPUT_4 D_INPUT_5 D_INPUT_6 D_INPUT_7 
+ VSS VDD 
+ INVX1_1164/A INVX1_1506/A INVX1_1096/A INVX1_1095/A INVX1_1386/A INVX1_1385/A INVX1_526/A INVX1_300/A INVX1_114/A INVX1_136/A INVX1_620/A INVX1_142/A INVX1_135/A INVX1_1344/A INVX1_755/A INVX1_592/A INVX1_591/A INVX1_1654/A INVX1_86/A INVX1_838/A INVX1_1068/A INVX1_756/A INVX1_1170/A INVX1_588/A INVX1_829/A INVX1_1250/A INVX1_796/A INVX1_795/A INVX1_587/A INVX1_186/A INVX1_1256/A INVX1_844/A INVX1_600/A INVX1_242/A INVX1_598/A INVX1_241/A INVX1_1212/A INVX1_1211/A INVX1_738/A INVX1_1026/A INVX1_492/A INVX1_556/A INVX1_491/A INVX1_922/A INVX1_921/A INVX1_511/A INVX1_252/A INVX1_12/A INVX1_1496/A INVX1_979/A INVX1_46/A 
+ INVX1_512/A INVX1_38/A INVX1_980/A INVX1_199/A INVX1_200/A INVX1_187/A INVX1_1222/A INVX1_764/A INVX1_258/A INVX1_160/A INVX1_163/A INVX1_582/A INVX1_1648/A INVX1_468/A INVX1_860/A INVX1_859/A INVX1_1175/A INVX1_818/A INVX1_817/A INVX1_1163/A INVX1_1525/A INVX1_1505/A INVX1_112/A INVX1_111/A INVX1_607/A INVX1_608/A INVX1_852/A INVX1_1387/A INVX1_1388/A INVX1_851/A INVX1_774/A INVX1_773/A INVX1_658/A INVX1_1192/A INVX1_1191/A INVX1_842/A INVX1_657/A INVX1_841/A INVX1_525/A INVX1_257/A INVX1_251/A INVX1_299/A INVX1_37/A INVX1_11/A INVX1_619/A INVX1_141/A INVX1_159/A INVX1_113/A INVX1_1221/A INVX1_188/A INVX1_164/A 
+ INVX1_45/A INVX1_1238/A INVX1_830/A INVX1_1237/A INVX1_763/A INVX1_1343/A INVX1_916/A INVX1_915/A INVX1_752/A INVX1_1176/A INVX1_1003/A INVX1_328/A INVX1_1004/A INVX1_1392/A INVX1_288/A INVX1_578/A INVX1_1627/A INVX1_566/A INVX1_618/A INVX1_976/A INVX1_1628/A INVX1_452/A INVX1_751/A INVX1_327/A INVX1_287/A INVX1_1391/A INVX1_809/A INVX1_1038/A INVX1_810/A INVX1_96/A INVX1_1384/A INVX1_1526/A INVX1_1653/A INVX1_1067/A INVX1_837/A INVX1_85/A INVX1_1694/A INVX1_1693/A INVX1_1037/A INVX1_95/A INVX1_1383/A INVX1_1495/A INVX1_310/A INVX1_309/A INVX1_1486/A INVX1_866/A INVX1_185/A INVX1_1255/A INVX1_843/A INVX1_555/A INVX1_737/A 
+ INVX1_597/A INVX1_599/A INVX1_1485/A INVX1_865/A INVX1_451/A INVX1_577/A INVX1_617/A INVX1_565/A INVX1_975/A INVX1_1169/A INVX1_1249/A INVX1_1602/A INVX1_581/A INVX1_1647/A INVX1_467/A INVX1_1382/A INVX1_646/A INVX1_1053/A INVX1_645/A INVX1_1054/A INVX1_222/A INVX1_221/A INVX1_1025/A INVX1_1381/A INVX1_1030/A INVX1_1029/A INVX1_552/A INVX1_1500/A INVX1_551/A INVX1_1499/A INVX1_1601/A INVX1_51/Y INVX1_24/Y INVX1_23/Y INVX1_52/Y INVX1_741/Y INVX1_742/Y INVX1_1198/Y INVX1_272/Y INVX1_612/Y INVX1_271/Y INVX1_823/Y INVX1_824/Y INVX1_611/Y INVX1_548/Y INVX1_547/Y INVX1_170/Y INVX1_169/Y INVX1_1197/Y INVX1_176/Y INVX1_175/Y 
+ INVX1_822/Y INVX1_821/Y INVX1_317/Y INVX1_318/Y INVX1_541/Y INVX1_542/Y INVX1_833/Y INVX1_834/Y INVX1_61/Y INVX1_62/Y INVX1_127/Y INVX1_128/Y INVX1_189/Y INVX1_190/Y INVX1_1377/Y INVX1_1378/Y INVX1_1021/Y INVX1_1022/Y INVX1_94/Y INVX1_93/Y INVX1_72/Y INVX1_71/Y INVX1_76/Y INVX1_75/Y INVX1_30/Y INVX1_29/Y INVX1_131/Y INVX1_132/Y INVX1_20/Y INVX1_44/Y INVX1_19/Y INVX1_43/Y INVX1_35/Y INVX1_102/Y INVX1_314/Y INVX1_208/Y INVX1_207/Y INVX1_313/Y INVX1_101/Y INVX1_36/Y INVX1_747/Y INVX1_748/Y INVX1_1640/Y INVX1_1639/Y INVX1_140/Y INVX1_139/Y INVX1_6/Y INVX1_97/Y INVX1_5/Y 
+ INVX1_110/Y INVX1_98/Y INVX1_109/Y INVX1_204/Y INVX1_203/Y INVX1_239/Y INVX1_240/Y INVX1_118/Y INVX1_117/Y INVX1_554/Y INVX1_489/Y INVX1_490/Y INVX1_553/Y INVX1_509/Y INVX1_510/Y INVX1_1398/Y INVX1_1397/Y INVX1_653/Y INVX1_654/Y INVX1_754/Y INVX1_753/Y INVX1_750/Y INVX1_154/Y INVX1_153/Y INVX1_87/Y INVX1_749/Y INVX1_88/Y INVX1_1060/Y INVX1_1059/Y INVX1_124/Y INVX1_123/Y INVX1_79/Y INVX1_80/Y INVX1_180/Y INVX1_179/Y INVX1_471/Y INVX1_472/Y INVX1_265/Y INVX1_266/Y INVX1_369/Y INVX1_370/Y INVX1_814/Y INVX1_813/Y INVX1_1198/A INVX1_548/A INVX1_547/A INVX1_1197/A INVX1_176/A INVX1_175/A INVX1_822/A INVX1_821/A 
+ INVX1_541/A INVX1_542/A INVX1_1377/A INVX1_1378/A INVX1_131/A INVX1_132/A INVX1_747/A INVX1_748/A INVX1_1640/A INVX1_1639/A INVX1_239/A INVX1_240/A INVX1_653/A INVX1_654/A INVX1_750/A INVX1_749/A INVX1_1060/A INVX1_1059/A INVX1_369/A INVX1_370/A NOR3X1_175/B NOR3X1_821/B NOR3X1_1599/C NOR3X1_747/B NOR3X1_653/B INVX1_1196/Y INVX1_1195/Y INVX1_546/Y INVX1_544/Y INVX1_545/Y INVX1_543/Y INVX1_174/Y INVX1_173/Y INVX1_820/Y INVX1_819/Y INVX1_1520/Y INVX1_1373/Y INVX1_1519/Y INVX1_1374/Y INVX1_537/Y INVX1_539/Y INVX1_540/Y INVX1_538/Y INVX1_1375/Y INVX1_1376/Y INVX1_643/Y INVX1_745/Y INVX1_746/Y INVX1_644/Y 
+ INVX1_1637/Y INVX1_1636/Y INVX1_1638/Y INVX1_1635/Y INVX1_125/Y INVX1_528/Y INVX1_527/Y INVX1_126/Y INVX1_145/Y INVX1_146/Y INVX1_174/A INVX1_173/A INVX1_820/A INVX1_819/A INVX1_1520/A INVX1_1373/A INVX1_1519/A INVX1_1374/A INVX1_537/A INVX1_539/A INVX1_540/A INVX1_538/A INVX1_745/A INVX1_746/A INVX1_528/A INVX1_527/A NOR3X1_1519/B INVX1_58/Y INVX1_57/Y INVX1_1370/Y INVX1_1372/Y INVX1_1371/Y INVX1_1369/Y INVX1_535/Y INVX1_536/Y INVX1_1370/A INVX1_1372/A INVX1_1371/A INVX1_1369/A NOR3X1_1371/C NOR3X1_1369/B INVX1_1364/Y INVX1_1362/Y INVX1_1363/Y INVX1_1361/Y INVX1_1368/Y INVX1_1366/Y INVX1_1367/Y INVX1_1365/Y INVX1_1364/A INVX1_1363/A 
+ INVX1_1366/A INVX1_1365/A 
+ AES_SBOX_0


* **************************************
* --- Simulation Settings ---
* **************************************

.param SIM_LEN = 50ns
.csparam SIM_LEN = {SIM_LEN}

.tran 0.1ns 'SIM_LEN'
.param SIMSTEP = 'SIM_LEN/0.1ns'
.csparam SIMSTEP = {SIMSTEP}

* **************************************
* --- Simulation Control ---
* **************************************

.control
    .include ../inputsD.inc

    run
    
    if ('writeFile' > 0)   
      wrdata ivdd_0.out i(vvdd)
      wrdata ivss_0.out i(vvss)
      *snsave sim_0.snap
    end
    
    set wr_vecnames
    set wr_singlescale
    wrdata outputs_0.out V("INVX1_1164/A") V("INVX1_1506/A") V("INVX1_1096/A") V("INVX1_1095/A") V("INVX1_1386/A") V("INVX1_1385/A") V("INVX1_526/A") V("INVX1_300/A") V("INVX1_114/A") V("INVX1_136/A") V("INVX1_620/A") V("INVX1_142/A") V("INVX1_135/A") V("INVX1_1344/A") V("INVX1_755/A") V("INVX1_592/A") V("INVX1_591/A") V("INVX1_1654/A") V("INVX1_86/A") V("INVX1_838/A") V("INVX1_1068/A") V("INVX1_756/A") V("INVX1_1170/A") V("INVX1_588/A") V("INVX1_829/A") V("INVX1_1250/A") V("INVX1_796/A") V("INVX1_795/A") V("INVX1_587/A") V("INVX1_186/A") V("INVX1_1256/A") V("INVX1_844/A") V("INVX1_600/A") V("INVX1_242/A") V("INVX1_598/A") V("INVX1_241/A") V("INVX1_1212/A") V("INVX1_1211/A") V("INVX1_738/A") V("INVX1_1026/A") V("INVX1_492/A") V("INVX1_556/A") V("INVX1_491/A") V("INVX1_922/A") V("INVX1_921/A") V("INVX1_511/A") V("INVX1_252/A") V("INVX1_12/A") V("INVX1_1496/A") V("INVX1_979/A") V("INVX1_46/A") V("INVX1_512/A") V("INVX1_38/A") V("INVX1_980/A") V("INVX1_199/A") V("INVX1_200/A") V("INVX1_187/A") V("INVX1_1222/A") V("INVX1_764/A") V("INVX1_258/A") V("INVX1_160/A") V("INVX1_163/A") V("INVX1_582/A") V("INVX1_1648/A") V("INVX1_468/A") V("INVX1_860/A") V("INVX1_859/A") V("INVX1_1175/A") V("INVX1_818/A") V("INVX1_817/A") V("INVX1_1163/A") V("INVX1_1525/A") V("INVX1_1505/A") V("INVX1_112/A") V("INVX1_111/A") V("INVX1_607/A") V("INVX1_608/A") V("INVX1_852/A") V("INVX1_1387/A") V("INVX1_1388/A") V("INVX1_851/A") V("INVX1_774/A") V("INVX1_773/A") V("INVX1_658/A") V("INVX1_1192/A") V("INVX1_1191/A") V("INVX1_842/A") V("INVX1_657/A") V("INVX1_841/A") V("INVX1_525/A") V("INVX1_257/A") V("INVX1_251/A") V("INVX1_299/A") V("INVX1_37/A") V("INVX1_11/A") V("INVX1_619/A") V("INVX1_141/A") V("INVX1_159/A") V("INVX1_113/A") V("INVX1_1221/A") V("INVX1_188/A") V("INVX1_164/A") V("INVX1_45/A") V("INVX1_1238/A") V("INVX1_830/A") V("INVX1_1237/A") V("INVX1_763/A") V("INVX1_1343/A") V("INVX1_916/A") V("INVX1_915/A") V("INVX1_752/A") V("INVX1_1176/A") V("INVX1_1003/A") V("INVX1_328/A") V("INVX1_1004/A") V("INVX1_1392/A") V("INVX1_288/A") V("INVX1_578/A") V("INVX1_1627/A") V("INVX1_566/A") V("INVX1_618/A") V("INVX1_976/A") V("INVX1_1628/A") V("INVX1_452/A") V("INVX1_751/A") V("INVX1_327/A") V("INVX1_287/A") V("INVX1_1391/A") V("INVX1_809/A") V("INVX1_1038/A") V("INVX1_810/A") V("INVX1_96/A") V("INVX1_1384/A") V("INVX1_1526/A") V("INVX1_1653/A") V("INVX1_1067/A") V("INVX1_837/A") V("INVX1_85/A") V("INVX1_1694/A") V("INVX1_1693/A") V("INVX1_1037/A") V("INVX1_95/A") V("INVX1_1383/A") V("INVX1_1495/A") V("INVX1_310/A") V("INVX1_309/A") V("INVX1_1486/A") V("INVX1_866/A") V("INVX1_185/A") V("INVX1_1255/A") V("INVX1_843/A") V("INVX1_555/A") V("INVX1_737/A") V("INVX1_597/A") V("INVX1_599/A") V("INVX1_1485/A") V("INVX1_865/A") V("INVX1_451/A") V("INVX1_577/A") V("INVX1_617/A") V("INVX1_565/A") V("INVX1_975/A") V("INVX1_1169/A") V("INVX1_1249/A") V("INVX1_1602/A") V("INVX1_581/A") V("INVX1_1647/A") V("INVX1_467/A") V("INVX1_1382/A") V("INVX1_646/A") V("INVX1_1053/A") V("INVX1_645/A") V("INVX1_1054/A") V("INVX1_222/A") V("INVX1_221/A") V("INVX1_1025/A") V("INVX1_1381/A") V("INVX1_1030/A") V("INVX1_1029/A") V("INVX1_552/A") V("INVX1_1500/A") V("INVX1_551/A") V("INVX1_1499/A") V("INVX1_1601/A") V("INVX1_51/Y") V("INVX1_24/Y") V("INVX1_23/Y") V("INVX1_52/Y") V("INVX1_741/Y") V("INVX1_742/Y") V("INVX1_1198/Y") V("INVX1_272/Y") V("INVX1_612/Y") V("INVX1_271/Y") V("INVX1_823/Y") V("INVX1_824/Y") V("INVX1_611/Y") V("INVX1_548/Y") V("INVX1_547/Y") V("INVX1_170/Y") V("INVX1_169/Y") V("INVX1_1197/Y") V("INVX1_176/Y") V("INVX1_175/Y") V("INVX1_822/Y") V("INVX1_821/Y") V("INVX1_317/Y") V("INVX1_318/Y") V("INVX1_541/Y") V("INVX1_542/Y") V("INVX1_833/Y") V("INVX1_834/Y") V("INVX1_61/Y") V("INVX1_62/Y") V("INVX1_127/Y") V("INVX1_128/Y") V("INVX1_189/Y") V("INVX1_190/Y") V("INVX1_1377/Y") V("INVX1_1378/Y") V("INVX1_1021/Y") V("INVX1_1022/Y") V("INVX1_94/Y") V("INVX1_93/Y") V("INVX1_72/Y") V("INVX1_71/Y") V("INVX1_76/Y") V("INVX1_75/Y") V("INVX1_30/Y") V("INVX1_29/Y") V("INVX1_131/Y") V("INVX1_132/Y") V("INVX1_20/Y") V("INVX1_44/Y") V("INVX1_19/Y") V("INVX1_43/Y") V("INVX1_35/Y") V("INVX1_102/Y") V("INVX1_314/Y") V("INVX1_208/Y") V("INVX1_207/Y") V("INVX1_313/Y") V("INVX1_101/Y") V("INVX1_36/Y") V("INVX1_747/Y") V("INVX1_748/Y") V("INVX1_1640/Y") V("INVX1_1639/Y") V("INVX1_140/Y") V("INVX1_139/Y") V("INVX1_6/Y") V("INVX1_97/Y") V("INVX1_5/Y") V("INVX1_110/Y") V("INVX1_98/Y") V("INVX1_109/Y") V("INVX1_204/Y") V("INVX1_203/Y") V("INVX1_239/Y") V("INVX1_240/Y") V("INVX1_118/Y") V("INVX1_117/Y") V("INVX1_554/Y") V("INVX1_489/Y") V("INVX1_490/Y") V("INVX1_553/Y") V("INVX1_509/Y") V("INVX1_510/Y") V("INVX1_1398/Y") V("INVX1_1397/Y") V("INVX1_653/Y") V("INVX1_654/Y") V("INVX1_754/Y") V("INVX1_753/Y") V("INVX1_750/Y") V("INVX1_154/Y") V("INVX1_153/Y") V("INVX1_87/Y") V("INVX1_749/Y") V("INVX1_88/Y") V("INVX1_1060/Y") V("INVX1_1059/Y") V("INVX1_124/Y") V("INVX1_123/Y") V("INVX1_79/Y") V("INVX1_80/Y") V("INVX1_180/Y") V("INVX1_179/Y") V("INVX1_471/Y") V("INVX1_472/Y") V("INVX1_265/Y") V("INVX1_266/Y") V("INVX1_369/Y") V("INVX1_370/Y") V("INVX1_814/Y") V("INVX1_813/Y") V("INVX1_1198/A") V("INVX1_548/A") V("INVX1_547/A") V("INVX1_1197/A") V("INVX1_176/A") V("INVX1_175/A") V("INVX1_822/A") V("INVX1_821/A") V("INVX1_541/A") V("INVX1_1377/A") V("INVX1_1378/A") V("INVX1_131/A") V("INVX1_132/A") V("INVX1_747/A") V("INVX1_748/A") V("INVX1_1640/A") V("INVX1_1639/A") V("INVX1_239/A") V("INVX1_240/A") V("INVX1_653/A") V("INVX1_654/A") V("INVX1_750/A") V("INVX1_749/A") V("INVX1_1060/A") V("INVX1_1059/A") V("INVX1_369/A") V("INVX1_370/A") V("NOR3X1_175/B") V("NOR3X1_821/B") V("NOR3X1_1599/C") V("NOR3X1_747/B") V("NOR3X1_653/B") V("INVX1_1196/Y") V("INVX1_1195/Y") V("INVX1_546/Y") V("INVX1_544/Y") V("INVX1_545/Y") V("INVX1_543/Y") V("INVX1_174/Y") V("INVX1_173/Y") V("INVX1_820/Y") V("INVX1_819/Y") V("INVX1_1520/Y") V("INVX1_1373/Y") V("INVX1_1519/Y") V("INVX1_1374/Y") V("INVX1_537/Y") V("INVX1_539/Y") V("INVX1_540/Y") V("INVX1_538/Y") V("INVX1_1375/Y") V("INVX1_1376/Y") V("INVX1_643/Y") V("INVX1_745/Y") V("INVX1_746/Y") V("INVX1_644/Y") V("INVX1_1637/Y") V("INVX1_1636/Y") V("INVX1_1638/Y") V("INVX1_1635/Y") V("INVX1_125/Y") V("INVX1_528/Y") V("INVX1_527/Y") V("INVX1_126/Y") V("INVX1_145/Y") V("INVX1_146/Y") V("INVX1_174/A") V("INVX1_173/A") V("INVX1_820/A") V("INVX1_819/A") V("INVX1_1520/A") V("INVX1_1373/A") V("INVX1_1519/A") V("INVX1_1374/A") V("INVX1_537/A") V("INVX1_539/A") V("INVX1_540/A") V("INVX1_538/A") V("INVX1_745/A") V("INVX1_746/A") V("INVX1_528/A") V("INVX1_527/A") V("NOR3X1_1519/B") V("INVX1_58/Y") V("INVX1_57/Y") V("INVX1_1370/Y") V("INVX1_1372/Y") V("INVX1_1371/Y") V("INVX1_1369/Y") V("INVX1_535/Y") V("INVX1_536/Y") V("INVX1_1370/A") V("INVX1_1372/A") V("INVX1_1371/A") V("INVX1_1369/A") V("NOR3X1_1371/C") V("NOR3X1_1369/B") V("INVX1_1364/Y") V("INVX1_1362/Y") V("INVX1_1363/Y") V("INVX1_1361/Y") V("INVX1_1368/Y") V("INVX1_1366/Y") V("INVX1_1367/Y") V("INVX1_1365/Y") V("INVX1_1364/A") V("INVX1_1363/A") V("INVX1_1366/A") V("INVX1_1365/A") 
    
    if ('showPlots' < 1)
        quit
    end
       
.endc

.end
