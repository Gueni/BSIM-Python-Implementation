*** TEST 005 partitioning ***
*
* ngSPICE test for PLS experiments
*
* AES SBOX PLS test init file generator - protected dualRail SBOX area illuminated
*
* Author: Jan Belohoubek, 08/2020
* jan.belohoubek@fit.cvut.cz
*
* https://users.fit.cvut.cz/~belohja4/
*
*
* **************************************

.include ../../models.lib
.include ../../tsmc180nmcmos.lib
.include secLibDualRail.spice

* **************************************
* --- Test ---
* **************************************

* --- Settings
.param showPlots = 0
.param writeFile = 1
.param run_inputSet = 0

* redefine defaults ...
.include test00X_settings.inc

.csparam showPlots = {showPlots}
.csparam writeFile = {writeFile}
.csparam run_inputSet = {run_inputSet}

.global showPlots writeFile run_inputSet

* --- End of Settins

Vtrig LaserTrig 0 0 PWL(0ns 0V 40ns 0V 41ns SUPP)

.param beamDistanceTop = 0
.param beamDistanceBot = 0

.global LaserTrig beamDistanceTop beamDistanceBot

* --- inputs
Vvin0 INPUT_0 0 0 PWL(0ns 0V 5ns  0V 7ns  0V)
Vvin1 INPUT_1 0 0 PWL(0ns 0V 6ns  0V 8ns  0V)
Vvin2 INPUT_2 0 0 PWL(0ns 0V 7ns  0V 9ns  0V)
Vvin3 INPUT_3 0 0 PWL(0ns 0V 8ns  0V 10ns 0V)
Vvin4 INPUT_4 0 0 PWL(0ns 0V 9ns  0V 11ns 0V)
Vvin5 INPUT_5 0 0 PWL(0ns 0V 10ns 0V 12ns 0V)
Vvin6 INPUT_6 0 0 PWL(0ns 0V 11ns 0V 13ns 0V)
Vvin7 INPUT_7 0 0 PWL(0ns 0V 12ns 0V 14ns 0V)

Vvin0D D_INPUT_0 0 0 PWL(0ns 0V 5ns  0V 7ns  0V)
Vvin1D D_INPUT_1 0 0 PWL(0ns 0V 6ns  0V 8ns  0V)
Vvin2D D_INPUT_2 0 0 PWL(0ns 0V 7ns  0V 9ns  0V)
Vvin3D D_INPUT_3 0 0 PWL(0ns 0V 8ns  0V 10ns 0V)
Vvin4D D_INPUT_4 0 0 PWL(0ns 0V 9ns  0V 11ns 0V)
Vvin5D D_INPUT_5 0 0 PWL(0ns 0V 10ns 0V 12ns 0V)
Vvin6D D_INPUT_6 0 0 PWL(0ns 0V 11ns 0V 13ns 0V)
Vvin7D D_INPUT_7 0 0 PWL(0ns 0V 12ns 0V 14ns 0V)


* --- outputs
*C0 VSS GATE_222 10fF
*C1 VSS GATE_366 10fF
*C2 VSS GATE_479 10fF
*C3 VSS GATE_579 10fF
*C4 VSS GATE_662 10fF
*C5 VSS GATE_741 10fF
*C6 VSS GATE_811 10fF
*C7 VSS GATE_865 10fF
*
*C0d VSS D_GATE_222 10fF
*C1d VSS D_GATE_366 10fF
*C2d VSS D_GATE_479 10fF
*C3d VSS D_GATE_579 10fF
*C4d VSS D_GATE_662 10fF
*C5d VSS D_GATE_741 10fF
*C6d VSS D_GATE_811 10fF
*C7d VSS D_GATE_865 10fF

* --- circuit layout model

Xsbox1 
+ NOR3X1_1619/A NOR3X1_1619/B NOR3X1_1620/B NOR3X1_951/A NOR3X1_951/B NOR3X1_952/B NOR3X1_724/B NOR3X1_723/A NOR3X1_723/B NOR3X1_1577/B NOR3X1_952/A NOR3X1_952/C NOR3X1_724/A NOR3X1_724/C NOR3X1_1147/B NOR3X1_1148/B NOR3X1_1147/A NOR3X1_1459/A NOR3X1_1459/B NOR3X1_1460/B NOR3X1_1711/A NOR3X1_1711/B NOR3X1_1712/B NOR3X1_1148/A NOR3X1_1148/C NOR3X1_678/A NOR3X1_678/C NOR3X1_677/B NOR3X1_678/B NOR3X1_677/A NOR3X1_1429/C NOR3X1_1430/A NOR3X1_1430/B NOR3X1_1430/C NOR3X1_1429/A NOR3X1_1460/A NOR3X1_1460/C NOR3X1_1712/A NOR3X1_1712/C NOR3X1_485/A NOR3X1_485/B NOR3X1_486/B NOR3X1_486/A NOR3X1_486/C NOR3X1_675/B NOR3X1_676/A NOR3X1_676/C NOR3X1_675/A NOR3X1_676/B NOR3X1_1620/C NOR3X1_1620/A 
+ NOR3X1_1264/B NOR3X1_1263/A NOR3X1_1263/B NOR3X1_1264/A NOR3X1_1264/C NOR3X1_1275/B NOR3X1_1113/C NOR3X1_675/C NOR3X1_1427/B NOR3X1_1428/A NOR3X1_1428/C NOR3X1_907/C NOR3X1_908/C NOR3X1_907/A NOR3X1_1428/B NOR3X1_1427/A NOR3X1_908/A NOR3X1_908/B NOR3X1_679/A NOR3X1_679/B NOR3X1_680/B NOR3X1_680/A NOR3X1_680/C NOR3X1_1681/B NOR3X1_1682/A NOR3X1_1682/C NOR3X1_1681/A NOR3X1_1682/B NOR3X1_1565/B NOR3X1_1566/A NOR3X1_1566/C NOR3X1_1565/A NOR3X1_1566/B NOR3X1_1681/C NOR3X1_1431/A NOR3X1_1431/B NOR3X1_1432/B NOR3X1_1432/A NOR3X1_1432/C NOR3X1_1103/B NOR3X1_1104/B NOR3X1_1103/A NOR3X1_1104/A NOR3X1_1104/C NOR3X1_1573/C NOR3X1_1574/A NOR3X1_1574/B NOR3X1_1699/B NOR3X1_1700/B NOR3X1_1699/A NOR3X1_1700/A 
+ NOR3X1_1700/C NOR3X1_1263/C NOR3X1_315/C NOR3X1_1586/C NOR3X1_1585/A NOR3X1_1585/C NOR3X1_1586/B NOR3X1_1586/A NOR3X1_1679/B NOR3X1_1680/A NOR3X1_1680/C NOR3X1_1565/C NOR3X1_1679/A NOR3X1_1680/B NOR3X1_398/B NOR3X1_397/A NOR3X1_397/B NOR3X1_398/C NOR3X1_398/A NOR3X1_1283/B NOR3X1_1117/B NOR3X1_1118/A NOR3X1_1118/C NOR3X1_1284/A NOR3X1_1284/C NOR3X1_1283/A NOR3X1_1118/B NOR3X1_1117/A NOR3X1_1284/B NOR3X1_1717/C NOR3X1_1718/C NOR3X1_1717/A NOR3X1_1718/A NOR3X1_1718/B NOR3X1_277/B NOR3X1_278/B NOR3X1_277/A NOR3X1_278/A NOR3X1_278/C NOR3X1_397/C NOR3X1_907/B NOR3X1_1134/C NOR3X1_1133/A NOR3X1_1133/C NOR3X1_1134/A NOR3X1_1134/B NOR3X1_1704/C NOR3X1_1703/A NOR3X1_1703/C NOR3X1_1704/A NOR3X1_1704/B 
+ NOR3X1_1425/B NOR3X1_1426/A NOR3X1_1426/C NOR3X1_1287/A NOR3X1_1287/B NOR3X1_1288/B NOR3X1_1467/A NOR3X1_950/C NOR3X1_1467/C NOR3X1_1468/C NOR3X1_949/A NOR3X1_949/C NOR3X1_1424/B NOR3X1_1423/A NOR3X1_1423/B NOR3X1_1424/A NOR3X1_1424/C NOR3X1_1454/C NOR3X1_1453/A NOR3X1_1453/C NOR3X1_705/A NOR3X1_705/B NOR3X1_706/B NOR3X1_706/A NOR3X1_706/C NOR3X1_1454/A NOR3X1_1454/B NOR3X1_340/C NOR3X1_339/A NOR3X1_339/C NOR3X1_340/A NOR3X1_340/B NOR3X1_1569/A NOR3X1_1569/B NOR3X1_1570/B NOR3X1_1570/A NOR3X1_1570/C NOR3X1_1434/C NOR3X1_1433/A NOR3X1_1433/C NOR3X1_1434/A NOR3X1_1434/B NOR3X1_674/A NOR3X1_674/B NOR3X1_673/C NOR3X1_1573/A NOR3X1_1574/C NOR3X1_1301/A NOR3X1_1301/C NOR3X1_1302/C NOR3X1_941/A 
+ NOR3X1_941/C NOR3X1_942/C NOR3X1_942/A NOR3X1_942/B NOR3X1_1247/C NOR3X1_1248/A NOR3X1_1248/B NOR3X1_1248/C NOR3X1_1247/A NOR3X1_1347/B NOR3X1_1533/B NOR3X1_157/B NOR3X1_1229/B NOR3X1_1033/B NOR3X1_1333/B NOR3X1_404/A NOR3X1_404/B NOR3X1_403/C NOR3X1_415/A NOR3X1_415/B NOR3X1_416/B NOR3X1_416/A NOR3X1_416/C NOR3X1_674/C NOR3X1_673/A NOR3X1_1583/C NOR3X1_1584/A NOR3X1_1584/B NOR3X1_1513/B NOR3X1_1568/B NOR3X1_1567/A NOR3X1_1567/B NOR3X1_1568/A NOR3X1_1568/C NOR3X1_303/B NOR3X1_373/B NOR3X1_1187/B NOR3X1_1359/B NOR3X1_1105/B NOR3X1_1106/A NOR3X1_1106/C NOR3X1_1509/B NOR3X1_1329/B NOR3X1_1217/B NOR3X1_1331/B NOR3X1_499/B NOR3X1_1189/B NOR3X1_995/B NOR3X1_377/B NOR3X1_1567/C NOR3X1_1279/A 
+ NOR3X1_1279/C NOR3X1_1280/C NOR3X1_1280/A NOR3X1_1280/B NOR3X1_919/C NOR3X1_261/B NOR3X1_987/B NOR3X1_485/C NOR3X1_1279/B NOR3X1_905/C NOR3X1_906/A NOR3X1_906/B NOR3X1_711/B NOR3X1_712/A NOR3X1_712/C NOR3X1_711/A NOR3X1_712/B NOR3X1_905/A NOR3X1_906/C NOR3X1_1287/C NOR3X1_1288/A NOR3X1_1288/C NOR3X1_1423/C NOR3X1_615/B NOR3X1_395/B NOR3X1_1585/B NOR3X1_1437/B NOR3X1_1438/A NOR3X1_1438/C NOR3X1_407/C NOR3X1_408/A NOR3X1_408/B NOR3X1_1555/B NOR3X1_1093/B NOR3X1_391/C NOR3X1_1559/B NOR3X1_361/B NOR3X1_362/A NOR3X1_362/C NOR3X1_387/B NOR3X1_388/A NOR3X1_388/C NOR3X1_1579/B NOR3X1_1557/B NOR3X1_1415/B NOR3X1_479/C NOR3X1_1283/C NOR3X1_923/C NOR3X1_419/C NOR3X1_420/A NOR3X1_420/B 
+ NOR3X1_361/C NOR3X1_362/B NOR3X1_1302/A NOR3X1_1302/B NOR3X1_280/C NOR3X1_279/B NOR3X1_280/A NOR3X1_385/B NOR3X1_386/A NOR3X1_386/C NOR3X1_521/B NOR3X1_679/C NOR3X1_1553/B NOR3X1_1437/C NOR3X1_1438/B NOR3X1_387/C NOR3X1_388/B NOR3X1_385/C NOR3X1_386/B NOR3X1_1117/C NOR3X1_603/C NOR3X1_1085/C NOR3X1_1269/C NOR3X1_901/C NOR3X1_453/C NOR3X1_1087/B NOR3X1_1088/A NOR3X1_1088/C NOR3X1_1265/C NOR3X1_1349/A NOR3X1_1349/B NOR3X1_1350/B NOR3X1_349/C NOR3X1_350/A NOR3X1_350/B NOR3X1_1350/C NOR3X1_1350/A NOR3X1_360/C NOR3X1_359/B NOR3X1_360/A NOR3X1_1407/C NOR3X1_405/C NOR3X1_406/A NOR3X1_406/B NOR3X1_899/B NOR3X1_1001/C NOR3X1_1002/A NOR3X1_1002/B NOR3X1_1001/A NOR3X1_1002/C NOR3X1_401/B 
+ NOR3X1_402/A NOR3X1_402/C NOR3X1_1709/B NOR3X1_1435/C NOR3X1_1436/A NOR3X1_1436/B NOR3X1_1663/C NOR3X1_1417/C NOR3X1_293/C NOR3X1_1039/C NOR3X1_1468/A NOR3X1_1468/B NOR3X1_950/A NOR3X1_950/B NOR3X1_1575/C NOR3X1_1576/A NOR3X1_1576/B NOR3X1_1069/C NOR3X1_1305/C NOR3X1_1306/A NOR3X1_1306/B NOR3X1_893/B NOR3X1_384/A NOR3X1_384/B NOR3X1_383/C NOR3X1_1671/C NOR3X1_1551/B NOR3X1_335/B NOR3X1_933/C NOR3X1_420/C NOR3X1_419/B NOR3X1_934/A NOR3X1_934/B NOR3X1_891/B NOR3X1_1011/C NOR3X1_484/A NOR3X1_484/B NOR3X1_483/C NOR3X1_1685/C NOR3X1_1090/C NOR3X1_1089/B NOR3X1_1090/A NOR3X1_1451/C NOR3X1_1452/A NOR3X1_1452/B NOR3X1_417/B NOR3X1_418/A NOR3X1_418/C NOR3X1_683/B NOR3X1_1564/A NOR3X1_1564/B 
+ NOR3X1_1563/C NOR3X1_1107/C NOR3X1_1108/A NOR3X1_1108/B NOR3X1_1413/B NOR3X1_1345/C NOR3X1_1537/B NOR3X1_1572/A NOR3X1_1572/C NOR3X1_1571/B NOR3X1_1089/C NOR3X1_1090/B NOR3X1_665/C NOR3X1_1097/C NOR3X1_781/B NOR3X1_389/C NOR3X1_1223/C NOR3X1_1281/B NOR3X1_1282/A NOR3X1_1282/C NOR3X1_1517/B NOR3X1_601/C NOR3X1_275/C NOR3X1_663/B NOR3X1_1337/B NOR3X1_1267/C NOR3X1_667/C NOR3X1_1285/B NOR3X1_1286/A NOR3X1_1286/C NOR3X1_359/C NOR3X1_360/B NOR3X1_133/B NOR3X1_777/C NOR3X1_1667/B NOR3X1_1355/B NOR3X1_1087/C NOR3X1_1088/B NOR3X1_359/A NOR3X1_1089/A NOR3X1_1564/C NOR3X1_1563/A NOR3X1_387/A NOR3X1_1583/A NOR3X1_1584/C NOR3X1_404/C NOR3X1_403/A NOR3X1_361/A NOR3X1_484/C NOR3X1_483/A NOR3X1_1087/A 
+ NOR3X1_431/A NOR3X1_1311/A NOR3X1_431/C NOR3X1_1311/C NOR3X1_432/C NOR3X1_1312/C NOR3X1_432/A NOR3X1_432/B NOR3X1_1312/A NOR3X1_1312/B NOR3X1_1121/A NOR3X1_1121/C NOR3X1_1122/C NOR3X1_696/C NOR3X1_695/A NOR3X1_695/C NOR3X1_1122/A NOR3X1_1122/B NOR3X1_385/A NOR3X1_696/A NOR3X1_696/B NOR3X1_697/A NOR3X1_697/C NOR3X1_698/C NOR3X1_698/A NOR3X1_698/B NOR3X1_247/C NOR3X1_248/A NOR3X1_248/B NOR3X1_248/C NOR3X1_247/A NOR3X1_1110/C NOR3X1_1109/B NOR3X1_1110/A NOR3X1_1109/A NOR3X1_1110/B NOR3X1_1105/A NOR3X1_1106/B NOR3X1_693/C NOR3X1_694/A NOR3X1_694/B NOR3X1_693/A NOR3X1_694/C NOR3X1_403/B NOR3X1_405/A NOR3X1_406/C NOR3X1_350/C NOR3X1_349/A NOR3X1_401/A NOR3X1_402/B NOR3X1_1572/B 
+ NOR3X1_1571/A NOR3X1_1425/A NOR3X1_1426/B NOR3X1_1130/C NOR3X1_1129/A NOR3X1_1129/C NOR3X1_1130/A NOR3X1_1130/B NOR3X1_933/A NOR3X1_419/A NOR3X1_934/C NOR3X1_1451/A NOR3X1_1452/C NOR3X1_418/B NOR3X1_417/A NOR3X1_1107/A NOR3X1_1108/C NOR3X1_1435/A NOR3X1_1436/C NOR3X1_1285/A NOR3X1_1286/B NOR3X1_1282/B NOR3X1_1281/A NOR3X1_1437/A NOR3X1_408/C NOR3X1_407/A NOR3X1_279/A NOR3X1_280/B NOR3X1_1305/A NOR3X1_1306/C NOR3X1_1576/C NOR3X1_1575/A NOR3X1_384/C NOR3X1_383/A INVX1_965/Y INVX1_966/Y INVX1_534/Y INVX1_533/Y INVX1_323/A INVX1_324/A INVX1_1673/A INVX1_1674/A INVX1_965/A INVX1_966/A 
+ INVX1_1257/A INVX1_1258/A INVX1_567/A INVX1_568/A INVX1_508/A INVX1_507/A INVX1_197/A INVX1_198/A INVX1_662/A INVX1_661/A INVX1_1241/A INVX1_1242/A INVX1_913/A INVX1_914/A INVX1_569/A INVX1_570/A INVX1_1691/A INVX1_1692/A INVX1_534/A INVX1_533/A NOR3X1_197/C NOR3X1_232/A NOR3X1_232/B NOR3X1_232/C NOR3X1_231/A NOR3X1_231/B NOR3X1_231/C INVX1_194/Y INVX1_193/Y INVX1_229/Y INVX1_227/Y INVX1_230/Y INVX1_228/Y INVX1_194/A INVX1_193/A INVX1_229/A INVX1_227/A INVX1_230/A INVX1_228/A NOR3X1_1596/A NOR3X1_1596/B NOR3X1_1596/C NOR3X1_1598/A NOR3X1_1598/B NOR3X1_1598/C NOR3X1_1597/A NOR3X1_1597/B NOR3X1_1595/A NOR3X1_1595/B NOR3X1_227/B INVX1_871/Y 
+ INVX1_872/Y INVX1_226/Y INVX1_225/Y INVX1_871/A INVX1_872/A INVX1_1185/A INVX1_1186/A INVX1_226/A INVX1_225/A NOR3X1_871/C NOR3X1_637/A NOR3X1_637/B NOR3X1_637/C NOR3X1_638/A NOR3X1_638/B NOR3X1_638/C NOR3X1_1185/B NOR3X1_1077/A NOR3X1_1077/B NOR3X1_1077/C NOR3X1_1078/A NOR3X1_1078/B NOR3X1_1078/C INVX1_868/Y INVX1_867/Y INVX1_634/Y INVX1_636/Y INVX1_635/Y INVX1_633/Y INVX1_1184/Y INVX1_1183/Y INVX1_1074/Y INVX1_1076/Y INVX1_1075/Y INVX1_1073/Y INVX1_868/A INVX1_867/A INVX1_634/A INVX1_636/A INVX1_635/A INVX1_633/A INVX1_1184/A INVX1_1183/A INVX1_1074/A INVX1_1076/A INVX1_1075/A INVX1_1073/A INVX1_1548/Y INVX1_1547/Y INVX1_944/Y INVX1_943/Y 
+ INVX1_575/Y INVX1_576/Y INVX1_1019/Y INVX1_1020/Y INVX1_1456/Y INVX1_1455/Y INVX1_1708/Y INVX1_1707/Y INVX1_121/Y INVX1_122/Y INVX1_1403/Y INVX1_1404/Y INVX1_1092/Y INVX1_1091/Y INVX1_647/Y INVX1_648/Y INVX1_1669/Y INVX1_1670/Y INVX1_1535/Y INVX1_1536/Y INVX1_1405/Y INVX1_1406/Y INVX1_456/Y INVX1_455/Y INVX1_1083/Y INVX1_1084/Y INVX1_971/Y INVX1_972/Y INVX1_1683/Y INVX1_1684/Y INVX1_1665/Y INVX1_1666/Y INVX1_1697/Y INVX1_1698/Y INVX1_273/Y INVX1_274/Y INVX1_1014/Y INVX1_1013/Y INVX1_651/Y INVX1_652/Y INVX1_1677/Y INVX1_1678/Y INVX1_1540/Y INVX1_1539/Y INVX1_1409/Y INVX1_1410/Y INVX1_1442/Y INVX1_947/Y INVX1_1441/Y INVX1_948/Y INVX1_295/Y 
+ INVX1_296/Y INVX1_887/Y INVX1_888/Y INVX1_606/Y INVX1_605/Y INVX1_337/Y INVX1_338/Y INVX1_1550/Y INVX1_1549/Y INVX1_985/Y INVX1_986/Y INVX1_671/Y INVX1_672/Y INVX1_1278/Y INVX1_1277/Y INVX1_930/Y INVX1_929/Y INVX1_1440/Y INVX1_1439/Y INVX1_779/Y INVX1_780/Y INVX1_1245/Y INVX1_1246/Y INVX1_517/Y INVX1_518/Y INVX1_1291/Y INVX1_1292/Y INVX1_70/Y INVX1_69/Y INVX1_1581/Y INVX1_1582/Y INVX1_1079/Y INVX1_1080/Y INVX1_897/Y INVX1_898/Y INVX1_707/Y INVX1_708/Y INVX1_776/Y INVX1_775/Y INVX1_1271/Y INVX1_1272/Y INVX1_167/Y INVX1_168/Y INVX1_1046/Y INVX1_997/Y INVX1_998/Y INVX1_1045/Y INVX1_1239/Y INVX1_1240/Y INVX1_256/Y INVX1_255/Y 
+ INVX1_1543/Y INVX1_1544/Y INVX1_801/Y INVX1_802/Y INVX1_878/Y INVX1_877/Y INVX1_347/Y INVX1_348/Y INVX1_151/Y INVX1_152/Y INVX1_999/Y INVX1_1000/Y INVX1_1209/Y INVX1_1210/Y INVX1_1203/Y INVX1_1204/Y INVX1_1303/Y INVX1_1304/Y INVX1_1659/Y INVX1_1660/Y INVX1_381/Y INVX1_382/Y INVX1_1358/Y INVX1_1357/Y INVX1_903/Y INVX1_904/Y INVX1_481/Y INVX1_482/Y INVX1_1421/Y INVX1_1422/Y INVX1_297/Y INVX1_298/Y INVX1_1561/Y INVX1_1562/Y INVX1_885/Y INVX1_886/Y INVX1_379/Y INVX1_380/Y INVX1_461/Y INVX1_462/Y INVX1_1294/Y INVX1_1293/Y INVX1_1116/Y INVX1_1115/Y INVX1_689/Y INVX1_690/Y INVX1_925/Y INVX1_926/Y INVX1_686/Y INVX1_685/Y INVX1_245/Y 
+ INVX1_246/Y INVX1_799/Y INVX1_800/Y INVX1_691/Y INVX1_692/Y INVX1_1420/Y INVX1_1419/Y INVX1_1099/Y INVX1_1100/Y INVX1_944/A INVX1_943/A INVX1_575/A INVX1_576/A INVX1_1456/A INVX1_1455/A INVX1_1708/A INVX1_1707/A INVX1_121/A INVX1_122/A INVX1_1403/A INVX1_1404/A INVX1_1092/A INVX1_1091/A INVX1_647/A INVX1_648/A INVX1_1669/A INVX1_1670/A INVX1_1535/A INVX1_1536/A INVX1_1405/A INVX1_1406/A INVX1_456/A INVX1_455/A INVX1_1083/A INVX1_1084/A INVX1_971/A INVX1_972/A INVX1_1683/A INVX1_1684/A INVX1_1665/A INVX1_1666/A INVX1_273/A INVX1_274/A INVX1_1014/A INVX1_1013/A INVX1_651/A INVX1_652/A INVX1_1677/A INVX1_1678/A INVX1_1540/A INVX1_1539/A 
+ INVX1_1409/A INVX1_1410/A INVX1_1442/A INVX1_1441/A INVX1_295/A INVX1_296/A INVX1_887/A INVX1_888/A INVX1_606/A INVX1_605/A INVX1_337/A INVX1_338/A INVX1_1550/A INVX1_1549/A INVX1_985/A INVX1_986/A INVX1_671/A INVX1_672/A INVX1_1278/A INVX1_1277/A INVX1_1440/A INVX1_1439/A INVX1_779/A INVX1_780/A INVX1_1245/A INVX1_1246/A INVX1_517/A INVX1_518/A INVX1_1291/A INVX1_1292/A INVX1_1581/A INVX1_1582/A INVX1_1079/A INVX1_1080/A INVX1_897/A INVX1_898/A INVX1_776/A INVX1_775/A INVX1_1271/A INVX1_1272/A INVX1_167/A INVX1_168/A INVX1_1046/A INVX1_997/A INVX1_998/A INVX1_1045/A INVX1_1239/A INVX1_1240/A INVX1_256/A INVX1_255/A INVX1_1543/A 
+ INVX1_1544/A INVX1_801/A INVX1_802/A INVX1_878/A INVX1_877/A INVX1_347/A INVX1_348/A INVX1_151/A INVX1_152/A INVX1_999/A INVX1_1000/A INVX1_1209/A INVX1_1210/A INVX1_1203/A INVX1_1204/A INVX1_1659/A INVX1_1660/A INVX1_381/A INVX1_382/A INVX1_1358/A INVX1_1357/A INVX1_903/A INVX1_904/A INVX1_481/A INVX1_482/A INVX1_1421/A INVX1_1422/A INVX1_297/A INVX1_298/A INVX1_1561/A INVX1_1562/A INVX1_885/A INVX1_886/A INVX1_379/A INVX1_380/A INVX1_461/A INVX1_462/A INVX1_1294/A INVX1_1293/A INVX1_1116/A INVX1_1115/A INVX1_689/A INVX1_690/A INVX1_925/A INVX1_926/A INVX1_686/A INVX1_685/A INVX1_245/A INVX1_246/A INVX1_799/A INVX1_800/A 
+ INVX1_691/A INVX1_692/A INVX1_1420/A INVX1_1419/A INVX1_1099/A INVX1_1100/A NOR3X1_1548/A NOR3X1_1548/B NOR3X1_1548/C NOR3X1_1547/A NOR3X1_1547/B NOR3X1_1547/C NOR3X1_943/B NOR3X1_1019/A NOR3X1_1019/B NOR3X1_1019/C NOR3X1_1020/A NOR3X1_1020/B NOR3X1_1020/C NOR3X1_1455/C NOR3X1_1707/C NOR3X1_1683/B NOR3X1_1697/A NOR3X1_1697/B NOR3X1_1697/C NOR3X1_1698/A NOR3X1_1698/B NOR3X1_1698/C NOR3X1_651/C NOR3X1_1677/C NOR3X1_947/A NOR3X1_947/C NOR3X1_1441/B NOR3X1_948/A NOR3X1_948/B NOR3X1_948/C NOR3X1_887/B NOR3X1_1277/B NOR3X1_930/A NOR3X1_930/B NOR3X1_930/C NOR3X1_929/A NOR3X1_929/B NOR3X1_779/C NOR3X1_1245/B NOR3X1_70/A NOR3X1_70/B NOR3X1_70/C NOR3X1_69/A NOR3X1_69/B NOR3X1_69/C 
+ NOR3X1_707/A NOR3X1_707/B NOR3X1_708/A NOR3X1_708/B NOR3X1_708/C NOR3X1_1543/B NOR3X1_999/B NOR3X1_1303/A NOR3X1_1303/B NOR3X1_1303/C NOR3X1_1304/A NOR3X1_1304/B NOR3X1_1304/C NOR3X1_381/B NOR3X1_1421/B NOR3X1_297/B NOR3X1_1293/B NOR3X1_1115/C NOR3X1_689/C NOR3X1_1099/C INVX1_1545/Y INVX1_1541/Y INVX1_1546/Y INVX1_1542/Y INVX1_1016/Y INVX1_1018/Y INVX1_1017/Y INVX1_1015/Y INVX1_1688/Y INVX1_1690/Y INVX1_1689/Y INVX1_1687/Y INVX1_784/Y INVX1_808/Y INVX1_807/Y INVX1_783/Y INVX1_911/Y INVX1_909/Y INVX1_912/Y INVX1_910/Y INVX1_67/Y INVX1_65/Y INVX1_68/Y INVX1_66/Y INVX1_880/Y INVX1_879/Y INVX1_1545/A INVX1_1541/A INVX1_1546/A INVX1_1542/A INVX1_1016/A 
+ INVX1_1018/A INVX1_1017/A INVX1_1015/A INVX1_1688/A INVX1_1690/A INVX1_1689/A INVX1_1687/A INVX1_784/A INVX1_783/A INVX1_911/A INVX1_912/A INVX1_67/A INVX1_65/A INVX1_68/A INVX1_66/A INVX1_880/A INVX1_879/A NOR3X1_1545/B NOR3X1_1541/B NOR3X1_1015/B NOR3X1_1687/B NOR3X1_808/A NOR3X1_808/B NOR3X1_808/C NOR3X1_807/A NOR3X1_807/B NOR3X1_807/C NOR3X1_783/C NOR3X1_911/B NOR3X1_909/A NOR3X1_909/B NOR3X1_909/C NOR3X1_910/A NOR3X1_910/B NOR3X1_910/C NOR3X1_879/B INVX1_805/Y INVX1_803/Y INVX1_806/Y INVX1_804/Y INVX1_890/Y INVX1_889/Y INVX1_805/A INVX1_803/A INVX1_806/A INVX1_804/A INVX1_890/A INVX1_889/A NOR3X1_805/B NOR3X1_803/B INVX1_231/Y 
+ INVX1_232/Y INVX1_1186/Y INVX1_1185/Y INVX1_1077/Y INVX1_1078/Y INVX1_508/Y INVX1_507/Y INVX1_637/Y INVX1_638/Y INVX1_1374/Y INVX1_1373/Y 
+ VSS VDD 
+ INVX1_1624/A INVX1_732/A INVX1_957/A INVX1_731/A INVX1_1150/A INVX1_1726/A INVX1_1149/A INVX1_1447/A INVX1_1477/A INVX1_1725/A INVX1_1623/A INVX1_1448/A INVX1_1315/A INVX1_1724/A INVX1_1723/A INVX1_1136/A INVX1_1135/A INVX1_1474/A INVX1_958/A INVX1_1461/A INVX1_954/A INVX1_953/A INVX1_1316/A INVX1_1722/A INVX1_1721/A INVX1_428/A INVX1_427/A INVX1_730/A INVX1_729/A INVX1_1449/A INVX1_1472/A INVX1_1471/A INVX1_1473/A INVX1_1143/A INVX1_436/A INVX1_1320/A INVX1_435/A INVX1_1319/A INVX1_1142/A INVX1_1141/A INVX1_937/A INVX1_938/A INVX1_1144/A INVX1_1124/A INVX1_1123/A INVX1_1125/A INVX1_411/A INVX1_409/A INVX1_412/A INVX1_1450/A INVX1_1138/A 
+ INVX1_1137/A INVX1_1462/A INVX1_1126/A INVX1_410/A INVX1_1322/A INVX1_1321/A INVX1_1478/A INVX1_442/A INVX1_441/A INVX1_1548/Y INVX1_1547/Y INVX1_1019/Y INVX1_1020/Y INVX1_909/Y INVX1_910/Y INVX1_439/Y INVX1_440/Y INVX1_1308/Y INVX1_1307/Y INVX1_932/Y INVX1_931/Y INVX1_1127/Y INVX1_1128/Y INVX1_488/Y INVX1_487/Y INVX1_1111/Y INVX1_1112/Y INVX1_281/Y INVX1_282/Y INVX1_935/Y INVX1_936/Y INVX1_1120/Y INVX1_1119/Y INVX1_1310/Y INVX1_1309/Y INVX1_434/Y INVX1_433/Y INVX1_1465/Y INVX1_1466/Y 
+ INVX1_1470/Y INVX1_1469/Y INVX1_681/Y INVX1_682/Y INVX1_1299/Y INVX1_1300/Y INVX1_1289/Y INVX1_1290/Y INVX1_727/Y INVX1_728/Y INVX1_363/Y INVX1_364/Y INVX1_413/Y INVX1_414/Y INVX1_1719/Y INVX1_1720/Y INVX1_939/Y INVX1_940/Y INVX1_703/Y INVX1_704/Y INVX1_1705/Y INVX1_1706/Y INVX1_1132/Y INVX1_1131/Y INVX1_399/Y INVX1_400/Y INVX1_1715/Y INVX1_1716/Y INVX1_1702/Y INVX1_1701/Y INVX1_1101/Y INVX1_1102/Y INVX1_1621/Y INVX1_1622/Y INVX1_1714/Y INVX1_1713/Y INVX1_1146/Y INVX1_1145/Y INVX1_726/Y INVX1_725/Y INVX1_439/A INVX1_440/A INVX1_1310/A INVX1_1309/A INVX1_1465/A INVX1_1466/A INVX1_727/A INVX1_728/A INVX1_1621/A INVX1_1622/A INVX1_726/A 
+ INVX1_725/A NOR3X1_439/A NOR3X1_439/B NOR3X1_439/C NOR3X1_440/A NOR3X1_440/B NOR3X1_440/C NOR3X1_1310/A NOR3X1_1310/B NOR3X1_1310/C NOR3X1_1309/A NOR3X1_1309/B NOR3X1_1309/C NOR3X1_1465/A NOR3X1_1465/B NOR3X1_1465/C NOR3X1_1466/A NOR3X1_1466/B NOR3X1_1466/C NOR3X1_727/A NOR3X1_727/B NOR3X1_727/C NOR3X1_728/A NOR3X1_728/B NOR3X1_728/C NOR3X1_1621/A NOR3X1_1621/B NOR3X1_1621/C NOR3X1_1622/A NOR3X1_1622/B NOR3X1_1622/C NOR3X1_726/A NOR3X1_726/B NOR3X1_726/C NOR3X1_725/A NOR3X1_725/B NOR3X1_725/C INVX1_424/Y INVX1_426/Y INVX1_425/Y INVX1_423/Y INVX1_1297/Y INVX1_1295/Y INVX1_1298/Y INVX1_1296/Y INVX1_1444/Y INVX1_1446/Y INVX1_1445/Y INVX1_1443/Y INVX1_714/Y INVX1_716/Y 
+ INVX1_715/Y INVX1_713/Y INVX1_1614/Y INVX1_1616/Y INVX1_1615/Y INVX1_1613/Y INVX1_719/Y INVX1_717/Y INVX1_720/Y INVX1_718/Y INVX1_424/A INVX1_423/A INVX1_716/A INVX1_715/A INVX1_1614/A INVX1_1616/A INVX1_1615/A INVX1_1613/A NOR3X1_424/A NOR3X1_424/B NOR3X1_424/C NOR3X1_423/A NOR3X1_423/B NOR3X1_423/C NOR3X1_716/A NOR3X1_716/B NOR3X1_716/C NOR3X1_715/A NOR3X1_715/B NOR3X1_715/C NOR3X1_1614/A NOR3X1_1614/B NOR3X1_1614/C NOR3X1_1616/A NOR3X1_1616/B NOR3X1_1616/C NOR3X1_1615/A NOR3X1_1615/B NOR3X1_1615/C NOR3X1_1613/A NOR3X1_1613/B NOR3X1_1613/C INVX1_421/Y INVX1_422/Y INVX1_701/Y INVX1_699/Y INVX1_702/Y INVX1_700/Y INVX1_1611/Y INVX1_1609/Y INVX1_1612/Y 
+ INVX1_1610/Y INVX1_1607/Y INVX1_1605/Y INVX1_1608/Y INVX1_1606/Y INVX1_1607/A INVX1_1605/A INVX1_1608/A INVX1_1606/A NOR3X1_1607/A NOR3X1_1607/B NOR3X1_1607/C NOR3X1_1605/A NOR3X1_1605/B NOR3X1_1605/C NOR3X1_1608/A NOR3X1_1608/B NOR3X1_1608/C NOR3X1_1606/A NOR3X1_1606/B NOR3X1_1606/C INVX1_1588/Y INVX1_1590/Y INVX1_1589/Y INVX1_1587/Y INVX1_1592/Y INVX1_1594/Y INVX1_1593/Y INVX1_1591/Y INVX1_638/Y INVX1_637/Y INVX1_232/Y INVX1_231/Y INVX1_70/Y INVX1_69/Y INVX1_1077/Y INVX1_1078/Y INVX1_807/Y INVX1_808/Y 
+ AES_SBOX_3

.include outputs_2.plw

* **************************************
* --- Simulation Settings ---
* **************************************

.param SIM_LEN = 50ns
.csparam SIM_LEN = {SIM_LEN}

.tran 0.1ns 'SIM_LEN'
.param SIMSTEP = 'SIM_LEN/0.1ns'
.csparam SIMSTEP = {SIMSTEP}

* **************************************
* --- Simulation Control ---
* **************************************

.control
    .include ../inputsD.inc
    
    run
    
    if ('writeFile' > 0)   
      wrdata ivdd_3.out i(vvdd)
      wrdata ivss_3.out i(vvss)
      *snsave sim_3.snap
    end
    
    set wr_vecnames
    set wr_singlescale
    wrdata outputs_3.out V("INVX1_1624/A") V("INVX1_732/A") V("INVX1_957/A") V("INVX1_731/A") V("INVX1_1150/A") V("INVX1_1726/A") V("INVX1_1149/A") V("INVX1_1447/A") V("INVX1_1477/A") V("INVX1_1725/A") V("INVX1_1623/A") V("INVX1_1448/A") V("INVX1_1315/A") V("INVX1_1724/A") V("INVX1_1723/A") V("INVX1_1136/A") V("INVX1_1135/A") V("INVX1_1474/A") V("INVX1_958/A") V("INVX1_1461/A") V("INVX1_954/A") V("INVX1_953/A") V("INVX1_1316/A") V("INVX1_1722/A") V("INVX1_1721/A") V("INVX1_428/A") V("INVX1_427/A") V("INVX1_730/A") V("INVX1_729/A") V("INVX1_1449/A") V("INVX1_1472/A") V("INVX1_1471/A") V("INVX1_1473/A") V("INVX1_1143/A") V("INVX1_436/A") V("INVX1_1320/A") V("INVX1_435/A") V("INVX1_1319/A") V("INVX1_1142/A") V("INVX1_1141/A") V("INVX1_937/A") V("INVX1_938/A") V("INVX1_1144/A") V("INVX1_1124/A") V("INVX1_1123/A") V("INVX1_1125/A") V("INVX1_411/A") V("INVX1_409/A") V("INVX1_412/A") V("INVX1_1450/A") V("INVX1_1138/A") V("INVX1_1137/A") V("INVX1_1462/A") V("INVX1_1126/A") V("INVX1_410/A") V("INVX1_1322/A") V("INVX1_1321/A") V("INVX1_1478/A") V("INVX1_442/A") V("INVX1_441/A") V("INVX1_1548/Y") V("INVX1_1547/Y") V("INVX1_1019/Y") V("INVX1_1020/Y") V("INVX1_909/Y") V("INVX1_910/Y") V("INVX1_439/Y") V("INVX1_440/Y") V("INVX1_1308/Y") V("INVX1_1307/Y") V("INVX1_932/Y") V("INVX1_931/Y") V("INVX1_1127/Y") V("INVX1_1128/Y") V("INVX1_488/Y") V("INVX1_487/Y") V("INVX1_1111/Y") V("INVX1_1112/Y") V("INVX1_281/Y") V("INVX1_282/Y") V("INVX1_935/Y") V("INVX1_936/Y") V("INVX1_1120/Y") V("INVX1_1119/Y") V("INVX1_1310/Y") V("INVX1_1309/Y") V("INVX1_434/Y") V("INVX1_433/Y") V("INVX1_1465/Y") V("INVX1_1466/Y") V("INVX1_1470/Y") V("INVX1_1469/Y") V("INVX1_681/Y") V("INVX1_682/Y") V("INVX1_1299/Y") V("INVX1_1300/Y") V("INVX1_1289/Y") V("INVX1_1290/Y") V("INVX1_727/Y") V("INVX1_728/Y") V("INVX1_363/Y") V("INVX1_364/Y") V("INVX1_413/Y") V("INVX1_414/Y") V("INVX1_1719/Y") V("INVX1_1720/Y") V("INVX1_939/Y") V("INVX1_940/Y") V("INVX1_703/Y") V("INVX1_704/Y") V("INVX1_1705/Y") V("INVX1_1706/Y") V("INVX1_1132/Y") V("INVX1_1131/Y") V("INVX1_399/Y") V("INVX1_400/Y") V("INVX1_1715/Y") V("INVX1_1716/Y") V("INVX1_1702/Y") V("INVX1_1701/Y") V("INVX1_1101/Y") V("INVX1_1102/Y") V("INVX1_1621/Y") V("INVX1_1622/Y") V("INVX1_1714/Y") V("INVX1_1713/Y") V("INVX1_1146/Y") V("INVX1_1145/Y") V("INVX1_726/Y") V("INVX1_725/Y") V("INVX1_439/A") V("INVX1_440/A") V("INVX1_1310/A") V("INVX1_1309/A") V("INVX1_1465/A") V("INVX1_1466/A") V("INVX1_727/A") V("INVX1_728/A") V("INVX1_1621/A") V("INVX1_1622/A") V("INVX1_726/A") V("INVX1_725/A") V("NOR3X1_439/A") V("NOR3X1_439/B") V("NOR3X1_439/C") V("NOR3X1_440/A") V("NOR3X1_440/B") V("NOR3X1_440/C") V("NOR3X1_1310/A") V("NOR3X1_1310/B") V("NOR3X1_1310/C") V("NOR3X1_1309/A") V("NOR3X1_1309/B") V("NOR3X1_1309/C") V("NOR3X1_1465/A") V("NOR3X1_1465/B") V("NOR3X1_1465/C") V("NOR3X1_1466/A") V("NOR3X1_1466/B") V("NOR3X1_1466/C") V("NOR3X1_727/A") V("NOR3X1_727/B") V("NOR3X1_727/C") V("NOR3X1_728/A") V("NOR3X1_728/B") V("NOR3X1_728/C") V("NOR3X1_1621/A") V("NOR3X1_1621/B") V("NOR3X1_1621/C") V("NOR3X1_1622/A") V("NOR3X1_1622/B") V("NOR3X1_1622/C") V("NOR3X1_726/A") V("NOR3X1_726/B") V("NOR3X1_726/C") V("NOR3X1_725/A") V("NOR3X1_725/B") V("NOR3X1_725/C") V("INVX1_424/Y") V("INVX1_426/Y") V("INVX1_425/Y") V("INVX1_423/Y") V("INVX1_1297/Y") V("INVX1_1295/Y") V("INVX1_1298/Y") V("INVX1_1296/Y") V("INVX1_1444/Y") V("INVX1_1446/Y") V("INVX1_1445/Y") V("INVX1_1443/Y") V("INVX1_714/Y") V("INVX1_716/Y") V("INVX1_715/Y") V("INVX1_713/Y") V("INVX1_1614/Y") V("INVX1_1616/Y") V("INVX1_1615/Y") V("INVX1_1613/Y") V("INVX1_719/Y") V("INVX1_717/Y") V("INVX1_720/Y") V("INVX1_718/Y") V("INVX1_424/A") V("INVX1_423/A") V("INVX1_716/A") V("INVX1_715/A") V("INVX1_1614/A") V("INVX1_1616/A") V("INVX1_1615/A") V("INVX1_1613/A") V("NOR3X1_424/A") V("NOR3X1_424/B") V("NOR3X1_424/C") V("NOR3X1_423/A") V("NOR3X1_423/B") V("NOR3X1_423/C") V("NOR3X1_716/A") V("NOR3X1_716/B") V("NOR3X1_716/C") V("NOR3X1_715/A") V("NOR3X1_715/B") V("NOR3X1_715/C") V("NOR3X1_1614/A") V("NOR3X1_1614/B") V("NOR3X1_1614/C") V("NOR3X1_1616/A") V("NOR3X1_1616/B") V("NOR3X1_1616/C") V("NOR3X1_1615/A") V("NOR3X1_1615/B") V("NOR3X1_1615/C") V("NOR3X1_1613/A") V("NOR3X1_1613/B") V("NOR3X1_1613/C") V("INVX1_421/Y") V("INVX1_422/Y") V("INVX1_701/Y") V("INVX1_699/Y") V("INVX1_702/Y") V("INVX1_700/Y") V("INVX1_1611/Y") V("INVX1_1609/Y") V("INVX1_1612/Y") V("INVX1_1610/Y") V("INVX1_1607/Y") V("INVX1_1605/Y") V("INVX1_1608/Y") V("INVX1_1606/Y") V("INVX1_1607/A") V("INVX1_1605/A") V("INVX1_1608/A") V("INVX1_1606/A") V("NOR3X1_1607/A") V("NOR3X1_1607/B") V("NOR3X1_1607/C") V("NOR3X1_1605/A") V("NOR3X1_1605/B") V("NOR3X1_1605/C") V("NOR3X1_1608/A") V("NOR3X1_1608/B") V("NOR3X1_1608/C") V("NOR3X1_1606/A") V("NOR3X1_1606/B") V("NOR3X1_1606/C") V("INVX1_1588/Y") V("INVX1_1590/Y") V("INVX1_1589/Y") V("INVX1_1587/Y") V("INVX1_1592/Y") V("INVX1_1594/Y") V("INVX1_1593/Y") V("INVX1_1591/Y") V("INVX1_638/Y") V("INVX1_637/Y") V("INVX1_232/Y") V("INVX1_231/Y") V("INVX1_70/Y") V("INVX1_69/Y") V("INVX1_1077/Y") V("INVX1_1078/Y") V("INVX1_807/Y") V("INVX1_808/Y") 
    
    if ('showPlots' < 1)
        quit
    end
       
.endc

.end
