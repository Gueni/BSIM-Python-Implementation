*** TEST 005 partitioning ***
*
* ngSPICE test for PLS experiments
*
* AES SBOX PLS test init file generator - protected dualRail SBOX area illuminated
*
* Author: Jan Belohoubek, 08/2020
* jan.belohoubek@fit.cvut.cz
*
* https://users.fit.cvut.cz/~belohja4/
*
*
* **************************************

.include ../../models.lib
.include ../../tsmc180nmcmos.lib
.include secLibDualRail.spice

* **************************************
* --- Test ---
* **************************************

* --- Settings
.param showPlots = 0
.param writeFile = 1
.param run_inputSet = 0

* redefine defaults ...
.include test00X_settings.inc

.csparam showPlots = {showPlots}
.csparam writeFile = {writeFile}
.csparam run_inputSet = {run_inputSet}

.global showPlots writeFile run_inputSet

* --- End of Settins

Vtrig LaserTrig 0 0 PWL(0ns 0V 40ns 0V 41ns SUPP)

.param beamDistanceTop = 0
.param beamDistanceBot = 0

.global LaserTrig beamDistanceTop beamDistanceBot

* --- inputs
Vvin0 INPUT_0 0 0 PWL(0ns 0V 5ns  0V 7ns  0V)
Vvin1 INPUT_1 0 0 PWL(0ns 0V 6ns  0V 8ns  0V)
Vvin2 INPUT_2 0 0 PWL(0ns 0V 7ns  0V 9ns  0V)
Vvin3 INPUT_3 0 0 PWL(0ns 0V 8ns  0V 10ns 0V)
Vvin4 INPUT_4 0 0 PWL(0ns 0V 9ns  0V 11ns 0V)
Vvin5 INPUT_5 0 0 PWL(0ns 0V 10ns 0V 12ns 0V)
Vvin6 INPUT_6 0 0 PWL(0ns 0V 11ns 0V 13ns 0V)
Vvin7 INPUT_7 0 0 PWL(0ns 0V 12ns 0V 14ns 0V)

Vvin0D D_INPUT_0 0 0 PWL(0ns 0V 5ns  0V 7ns  0V)
Vvin1D D_INPUT_1 0 0 PWL(0ns 0V 6ns  0V 8ns  0V)
Vvin2D D_INPUT_2 0 0 PWL(0ns 0V 7ns  0V 9ns  0V)
Vvin3D D_INPUT_3 0 0 PWL(0ns 0V 8ns  0V 10ns 0V)
Vvin4D D_INPUT_4 0 0 PWL(0ns 0V 9ns  0V 11ns 0V)
Vvin5D D_INPUT_5 0 0 PWL(0ns 0V 10ns 0V 12ns 0V)
Vvin6D D_INPUT_6 0 0 PWL(0ns 0V 11ns 0V 13ns 0V)
Vvin7D D_INPUT_7 0 0 PWL(0ns 0V 12ns 0V 14ns 0V)


* --- circuit layout model

Xsbox1 
+ NOR3X1_1270/C NOR3X1_1269/B NOR3X1_1270/A NOR3X1_1579/C NOR3X1_1580/A NOR3X1_1580/B NOR3X1_377/C NOR3X1_367/B NOR3X1_267/C NOR3X1_378/C NOR3X1_368/B NOR3X1_268/C NOR3X1_377/A NOR3X1_264/B NOR3X1_1187/C NOR3X1_250/C NOR3X1_1188/C NOR3X1_263/A NOR3X1_263/B NOR3X1_267/A NOR3X1_367/A NOR3X1_249/A NOR3X1_1187/A NOR3X1_249/C NOR3X1_811/A NOR3X1_811/C NOR3X1_812/C NOR3X1_120/B NOR3X1_873/C NOR3X1_1217/C NOR3X1_984/C NOR3X1_1399/A NOR3X1_1509/A NOR3X1_1218/C NOR3X1_1399/C NOR3X1_161/A NOR3X1_1509/C NOR3X1_161/C NOR3X1_790/C NOR3X1_983/A NOR3X1_1217/A NOR3X1_162/C NOR3X1_983/C NOR3X1_789/A NOR3X1_789/C NOR3X1_1400/C NOR3X1_590/C NOR3X1_874/C NOR3X1_589/A NOR3X1_119/A NOR3X1_119/B 
+ NOR3X1_1510/C NOR3X1_589/C NOR3X1_873/A NOR3X1_1529/C NOR3X1_458/C NOR3X1_987/C NOR3X1_988/C NOR3X1_457/A NOR3X1_1205/A NOR3X1_1205/C NOR3X1_987/A NOR3X1_1206/C NOR3X1_261/A NOR3X1_261/C NOR3X1_262/C NOR3X1_1355/C NOR3X1_1356/A NOR3X1_1356/B NOR3X1_1530/C NOR3X1_457/C NOR3X1_1529/A NOR3X1_1214/C NOR3X1_39/A NOR3X1_513/A NOR3X1_39/C NOR3X1_513/C NOR3X1_157/C NOR3X1_1213/A NOR3X1_158/C NOR3X1_1331/A NOR3X1_1213/C NOR3X1_1010/C NOR3X1_1331/C NOR3X1_1332/C NOR3X1_157/A NOR3X1_1009/A NOR3X1_1009/C NOR3X1_1041/A NOR3X1_1041/C NOR3X1_40/C NOR3X1_514/C NOR3X1_1042/C NOR3X1_1533/C NOR3X1_1330/C NOR3X1_794/C NOR3X1_31/A NOR3X1_1329/A NOR3X1_793/A NOR3X1_31/C NOR3X1_1329/C NOR3X1_793/C 
+ NOR3X1_961/A NOR3X1_1534/C NOR3X1_32/C NOR3X1_14/C NOR3X1_961/C NOR3X1_254/C NOR3X1_962/C NOR3X1_13/A NOR3X1_253/A NOR3X1_13/C NOR3X1_253/C NOR3X1_1533/A NOR3X1_515/B NOR3X1_516/B NOR3X1_1007/B NOR3X1_1491/A NOR3X1_1491/B NOR3X1_1008/B NOR3X1_1492/B NOR3X1_315/A NOR3X1_1007/A NOR3X1_315/B NOR3X1_355/A NOR3X1_355/B NOR3X1_316/B NOR3X1_356/B NOR3X1_515/A NOR3X1_995/C NOR3X1_1207/C NOR3X1_996/A NOR3X1_1208/A NOR3X1_996/B NOR3X1_1208/B NOR3X1_233/B NOR3X1_144/A NOR3X1_144/B NOR3X1_143/C NOR3X1_354/A NOR3X1_354/C NOR3X1_1347/C NOR3X1_1348/A NOR3X1_234/A NOR3X1_1348/B NOR3X1_234/C NOR3X1_345/C NOR3X1_346/A NOR3X1_353/B NOR3X1_346/B NOR3X1_1641/B NOR3X1_875/B NOR3X1_1642/A 
+ NOR3X1_876/A NOR3X1_1642/C NOR3X1_876/C NOR3X1_583/A NOR3X1_1225/A NOR3X1_583/C NOR3X1_1225/C NOR3X1_1226/C NOR3X1_374/C NOR3X1_373/A NOR3X1_1490/C NOR3X1_785/A NOR3X1_373/C NOR3X1_785/B NOR3X1_331/A NOR3X1_331/B NOR3X1_786/B NOR3X1_332/B NOR3X1_1489/A NOR3X1_365/A NOR3X1_365/B NOR3X1_1489/C NOR3X1_366/B NOR3X1_881/A NOR3X1_884/C NOR3X1_881/C NOR3X1_584/C NOR3X1_882/C NOR3X1_883/A NOR3X1_883/C NOR3X1_53/A NOR3X1_53/B NOR3X1_165/A NOR3X1_165/C NOR3X1_166/C NOR3X1_1190/C NOR3X1_474/C NOR3X1_351/A NOR3X1_1189/A NOR3X1_351/C NOR3X1_1189/C NOR3X1_473/A NOR3X1_352/C NOR3X1_473/C NOR3X1_54/B NOR3X1_1043/A NOR3X1_994/C NOR3X1_116/C NOR3X1_1043/C NOR3X1_1229/A NOR3X1_1229/C 
+ NOR3X1_47/A NOR3X1_993/A NOR3X1_993/C NOR3X1_1044/C NOR3X1_115/A NOR3X1_1230/C NOR3X1_47/C NOR3X1_115/C NOR3X1_48/C NOR3X1_500/C NOR3X1_1643/C NOR3X1_624/B NOR3X1_623/A NOR3X1_623/B NOR3X1_499/A NOR3X1_1333/A NOR3X1_1005/A NOR3X1_499/C NOR3X1_1333/C NOR3X1_1005/C NOR3X1_333/A NOR3X1_1006/C NOR3X1_333/C NOR3X1_334/C NOR3X1_1334/C NOR3X1_641/A NOR3X1_1531/A NOR3X1_129/A NOR3X1_1644/C NOR3X1_641/B NOR3X1_129/B NOR3X1_1531/C NOR3X1_642/B NOR3X1_130/B NOR3X1_1532/C NOR3X1_1643/A NOR3X1_639/C NOR3X1_291/A NOR3X1_291/C NOR3X1_989/A NOR3X1_292/C NOR3X1_967/B NOR3X1_989/C NOR3X1_968/B NOR3X1_791/A NOR3X1_791/B NOR3X1_137/C NOR3X1_792/B NOR3X1_77/C NOR3X1_138/C NOR3X1_78/C 
+ NOR3X1_357/C NOR3X1_137/A NOR3X1_77/A NOR3X1_358/C NOR3X1_967/A NOR3X1_640/C NOR3X1_357/A NOR3X1_639/A NOR3X1_990/C NOR3X1_459/A NOR3X1_1165/A NOR3X1_459/B NOR3X1_981/A NOR3X1_1165/C NOR3X1_1200/C NOR3X1_981/C NOR3X1_460/B NOR3X1_1166/C NOR3X1_982/C NOR3X1_147/C NOR3X1_148/C NOR3X1_1033/A NOR3X1_1033/C NOR3X1_147/A NOR3X1_1199/A NOR3X1_1199/C NOR3X1_1051/A NOR3X1_64/B NOR3X1_1051/C NOR3X1_1052/C NOR3X1_1034/C NOR3X1_63/A NOR3X1_63/B NOR3X1_1513/A NOR3X1_970/C NOR3X1_1513/C NOR3X1_797/C NOR3X1_847/C NOR3X1_798/C NOR3X1_969/A NOR3X1_848/C NOR3X1_969/C NOR3X1_797/A NOR3X1_847/A NOR3X1_1401/A NOR3X1_244/C NOR3X1_1401/C NOR3X1_594/C NOR3X1_1402/C NOR3X1_243/A NOR3X1_243/C 
+ NOR3X1_593/A NOR3X1_1514/C NOR3X1_593/C NOR3X1_1047/A NOR3X1_1201/A NOR3X1_1201/B NOR3X1_1202/B NOR3X1_787/C NOR3X1_788/C NOR3X1_1494/C NOR3X1_787/A NOR3X1_1493/A NOR3X1_1493/C NOR3X1_304/C NOR3X1_1047/C NOR3X1_303/A NOR3X1_1048/C NOR3X1_303/C NOR3X1_1050/B NOR3X1_289/A NOR3X1_289/C NOR3X1_1167/A NOR3X1_325/A NOR3X1_1360/C NOR3X1_325/C NOR3X1_326/C NOR3X1_1167/B NOR3X1_1359/A NOR3X1_1359/C NOR3X1_1168/B NOR3X1_1049/A NOR3X1_1049/B NOR3X1_290/C NOR3X1_1097/B NOR3X1_1098/B NOR3X1_1097/A NOR3X1_1098/A NOR3X1_1098/C NOR3X1_1411/B NOR3X1_1412/A NOR3X1_1412/C NOR3X1_1417/B NOR3X1_1418/B NOR3X1_1417/A NOR3X1_1411/A NOR3X1_1412/B NOR3X1_1418/A NOR3X1_1418/C NOR3X1_233/A NOR3X1_233/C NOR3X1_130/C 
+ NOR3X1_129/C NOR3X1_1625/A NOR3X1_1625/B NOR3X1_1626/B NOR3X1_469/A NOR3X1_469/B NOR3X1_470/B NOR3X1_1267/B NOR3X1_1268/A NOR3X1_1268/C NOR3X1_1554/A NOR3X1_1554/B NOR3X1_1553/C NOR3X1_1265/B NOR3X1_1266/A NOR3X1_1266/C NOR3X1_1081/C NOR3X1_1082/A NOR3X1_1082/B NOR3X1_873/B NOR3X1_583/B NOR3X1_345/A NOR3X1_345/B NOR3X1_874/B NOR3X1_584/B NOR3X1_395/C NOR3X1_396/A NOR3X1_396/B NOR3X1_137/B NOR3X1_138/A NOR3X1_670/C NOR3X1_669/B NOR3X1_670/A NOR3X1_993/B NOR3X1_367/C NOR3X1_368/C NOR3X1_143/A NOR3X1_143/B NOR3X1_994/B NOR3X1_138/B NOR3X1_1555/C NOR3X1_1556/A NOR3X1_1556/B NOR3X1_1345/B NOR3X1_1346/A NOR3X1_1346/C NOR3X1_917/B NOR3X1_918/B NOR3X1_917/A NOR3X1_594/A NOR3X1_593/B 
+ NOR3X1_594/B NOR3X1_1675/C NOR3X1_1676/A NOR3X1_1676/B NOR3X1_389/B NOR3X1_390/A NOR3X1_390/C NOR3X1_1081/B NOR3X1_1082/C NOR3X1_1011/B NOR3X1_1012/A NOR3X1_1012/C NOR3X1_894/A NOR3X1_894/B NOR3X1_893/C NOR3X1_1070/C NOR3X1_1069/B NOR3X1_1070/A NOR3X1_275/B NOR3X1_276/A NOR3X1_276/C NOR3X1_918/A NOR3X1_918/C NOR3X1_961/B NOR3X1_962/A NOR3X1_589/B NOR3X1_590/A NOR3X1_1261/B NOR3X1_1262/A NOR3X1_1262/C NOR3X1_797/B NOR3X1_798/A NOR3X1_798/B NOR3X1_590/B NOR3X1_962/B NOR3X1_1259/C NOR3X1_1260/A NOR3X1_1260/B NOR3X1_895/B NOR3X1_896/A NOR3X1_896/C NOR3X1_601/B NOR3X1_602/A NOR3X1_602/C NOR3X1_1661/B NOR3X1_1662/A NOR3X1_1662/C NOR3X1_244/A NOR3X1_243/B NOR3X1_604/A NOR3X1_604/C 
+ NOR3X1_603/B NOR3X1_244/B NOR3X1_1214/A NOR3X1_1213/B NOR3X1_1214/B NOR3X1_1085/B NOR3X1_1086/A NOR3X1_1086/C NOR3X1_1031/C NOR3X1_1032/A NOR3X1_1032/B NOR3X1_967/C NOR3X1_968/C NOR3X1_1007/C NOR3X1_1008/C NOR3X1_1194/C NOR3X1_1193/A NOR3X1_1050/C NOR3X1_1193/C NOR3X1_1641/A NOR3X1_641/C NOR3X1_1641/C NOR3X1_642/C NOR3X1_1049/C NOR3X1_1337/A NOR3X1_1207/B NOR3X1_1207/A NOR3X1_1489/B NOR3X1_333/B NOR3X1_1490/B NOR3X1_1337/C NOR3X1_334/B NOR3X1_1051/B NOR3X1_1338/C NOR3X1_1052/B NOR3X1_1530/A NOR3X1_1201/C NOR3X1_1202/A NOR3X1_31/B NOR3X1_331/C NOR3X1_32/A NOR3X1_332/A NOR3X1_1529/B NOR3X1_683/C NOR3X1_684/A NOR3X1_684/B NOR3X1_1685/B NOR3X1_1686/A NOR3X1_573/C NOR3X1_1686/C NOR3X1_574/A 
+ NOR3X1_574/B NOR3X1_147/B NOR3X1_148/B NOR3X1_1491/C NOR3X1_1492/C NOR3X1_683/A NOR3X1_684/C NOR3X1_924/B NOR3X1_923/A NOR3X1_923/B NOR3X1_924/A NOR3X1_924/C NOR3X1_687/A NOR3X1_687/B NOR3X1_688/B NOR3X1_291/B NOR3X1_984/B NOR3X1_292/B NOR3X1_787/B NOR3X1_983/B NOR3X1_788/B NOR3X1_254/B NOR3X1_253/B NOR3X1_53/C NOR3X1_459/C NOR3X1_14/B NOR3X1_365/C NOR3X1_366/C NOR3X1_1167/C NOR3X1_13/B NOR3X1_1168/C NOR3X1_54/C NOR3X1_460/C NOR3X1_1577/C NOR3X1_1578/A NOR3X1_1578/B NOR3X1_522/C NOR3X1_789/B NOR3X1_790/B NOR3X1_357/B NOR3X1_1199/B NOR3X1_358/B NOR3X1_1200/B NOR3X1_884/B NOR3X1_249/B NOR3X1_250/B NOR3X1_521/A NOR3X1_883/B NOR3X1_521/C NOR3X1_1114/B NOR3X1_1113/A 
+ NOR3X1_1113/B NOR3X1_791/C NOR3X1_792/C NOR3X1_1009/B NOR3X1_1010/B NOR3X1_875/A NOR3X1_47/B NOR3X1_875/C NOR3X1_457/B NOR3X1_48/B NOR3X1_458/B NOR3X1_688/C NOR3X1_688/A NOR3X1_39/B NOR3X1_40/B NOR3X1_1114/A NOR3X1_1114/C NOR3X1_201/B NOR3X1_202/A NOR3X1_202/C NOR3X1_201/A NOR3X1_202/B NOR3X1_640/B NOR3X1_1399/B NOR3X1_1400/B NOR3X1_264/C NOR3X1_351/B NOR3X1_352/B NOR3X1_263/C NOR3X1_1531/B NOR3X1_1532/B NOR3X1_639/B NOR3X1_1625/C NOR3X1_1626/A NOR3X1_469/C NOR3X1_470/A NOR3X1_515/C NOR3X1_516/C NOR3X1_289/B NOR3X1_847/B NOR3X1_290/B NOR3X1_848/B NOR3X1_1643/B NOR3X1_1043/B NOR3X1_981/B NOR3X1_982/B NOR3X1_969/B NOR3X1_970/B NOR3X1_1644/B NOR3X1_1044/B NOR3X1_1223/A 
+ NOR3X1_1223/B NOR3X1_1224/B NOR3X1_1225/B NOR3X1_1226/B NOR3X1_989/B NOR3X1_624/C NOR3X1_990/B NOR3X1_134/C NOR3X1_623/C NOR3X1_355/C NOR3X1_356/C NOR3X1_133/A NOR3X1_133/C NOR3X1_63/C NOR3X1_64/C NOR3X1_781/C NOR3X1_782/A NOR3X1_782/B NOR3X1_513/B NOR3X1_267/B NOR3X1_268/B NOR3X1_1351/C NOR3X1_1352/A NOR3X1_1352/B NOR3X1_1047/B NOR3X1_1048/B NOR3X1_514/B NOR3X1_1518/C NOR3X1_1517/A NOR3X1_474/B NOR3X1_1401/B NOR3X1_473/B NOR3X1_1402/B NOR3X1_1517/C NOR3X1_77/B NOR3X1_785/C NOR3X1_78/B NOR3X1_786/C NOR3X1_120/C NOR3X1_119/C NOR3X1_161/B NOR3X1_162/B NOR3X1_165/B NOR3X1_794/A NOR3X1_166/A NOR3X1_793/B NOR3X1_1165/B NOR3X1_1166/B NOR3X1_1205/B NOR3X1_1206/B NOR3X1_1494/B 
+ NOR3X1_1493/B NOR3X1_881/B NOR3X1_353/A NOR3X1_882/B NOR3X1_353/C NOR3X1_1041/B NOR3X1_115/B NOR3X1_1042/B NOR3X1_116/B NOR3X1_667/B NOR3X1_668/A NOR3X1_668/C NOR3X1_1671/B NOR3X1_1672/A NOR3X1_1672/C NOR3X1_480/C NOR3X1_479/B NOR3X1_480/A NOR3X1_166/B NOR3X1_474/A NOR3X1_352/A NOR3X1_1190/A NOR3X1_1190/B NOR3X1_54/A NOR3X1_984/A NOR3X1_1218/A NOR3X1_1218/B NOR3X1_1400/A NOR3X1_1510/A NOR3X1_1510/B NOR3X1_162/A NOR3X1_790/A NOR3X1_874/A NOR3X1_120/A NOR3X1_1226/A NOR3X1_374/A NOR3X1_374/B NOR3X1_786/A NOR3X1_332/C NOR3X1_1490/A NOR3X1_366/A NOR3X1_884/A NOR3X1_584/A NOR3X1_882/A NOR3X1_1202/C NOR3X1_788/A NOR3X1_1494/A NOR3X1_304/A NOR3X1_304/B NOR3X1_1048/A NOR3X1_901/B 
+ NOR3X1_902/A NOR3X1_902/C NOR3X1_901/A NOR3X1_902/B NOR3X1_290/A NOR3X1_326/A NOR3X1_326/B NOR3X1_1168/A NOR3X1_1360/A NOR3X1_1360/B NOR3X1_1050/A NOR3X1_378/A NOR3X1_378/B NOR3X1_268/A NOR3X1_368/A NOR3X1_264/A NOR3X1_1188/A NOR3X1_1188/B NOR3X1_250/A NOR3X1_812/A NOR3X1_812/B NOR3X1_624/A NOR3X1_500/A NOR3X1_1006/A NOR3X1_500/B NOR3X1_1006/B NOR3X1_334/A NOR3X1_1334/A NOR3X1_1644/A NOR3X1_1334/B NOR3X1_642/A NOR3X1_1532/A NOR3X1_130/A NOR3X1_995/A NOR3X1_996/C NOR3X1_1208/C NOR3X1_144/C NOR3X1_354/B NOR3X1_234/B NOR3X1_1348/C NOR3X1_346/C NOR3X1_1347/A NOR3X1_1642/B NOR3X1_876/B NOR3X1_460/A NOR3X1_1166/A NOR3X1_982/A NOR3X1_148/A NOR3X1_1200/A NOR3X1_64/A NOR3X1_1052/A 
+ NOR3X1_1034/A NOR3X1_1034/B NOR3X1_794/B NOR3X1_1534/A NOR3X1_1534/B NOR3X1_1330/A NOR3X1_14/A NOR3X1_32/B NOR3X1_1330/B NOR3X1_254/A NOR3X1_1530/B NOR3X1_988/A NOR3X1_988/B NOR3X1_1206/A NOR3X1_262/A NOR3X1_262/B NOR3X1_1355/A NOR3X1_1356/C NOR3X1_458/A NOR3X1_1230/A NOR3X1_1230/B NOR3X1_1044/A NOR3X1_48/A NOR3X1_994/A NOR3X1_116/A NOR3X1_1275/A NOR3X1_1275/C NOR3X1_1276/C NOR3X1_516/A NOR3X1_1008/A NOR3X1_1492/A NOR3X1_316/A NOR3X1_356/A NOR3X1_316/C NOR3X1_640/A NOR3X1_292/A NOR3X1_968/A NOR3X1_990/A NOR3X1_792/A NOR3X1_78/A NOR3X1_358/A NOR3X1_848/A NOR3X1_970/A NOR3X1_1402/A NOR3X1_1514/A NOR3X1_1514/B NOR3X1_40/A NOR3X1_158/A NOR3X1_158/B NOR3X1_1332/A NOR3X1_1332/B 
+ NOR3X1_1010/A NOR3X1_514/A NOR3X1_1042/A NOR3X1_920/C NOR3X1_919/B NOR3X1_920/A NOR3X1_919/A NOR3X1_920/B NOR3X1_1269/A NOR3X1_1270/B NOR3X1_1537/C NOR3X1_1538/C NOR3X1_1537/A NOR3X1_1579/A NOR3X1_1580/C NOR3X1_899/C NOR3X1_900/A NOR3X1_900/B NOR3X1_1414/C NOR3X1_1413/A NOR3X1_1413/C NOR3X1_1414/A NOR3X1_1414/B NOR3X1_900/C NOR3X1_899/A NOR3X1_777/B NOR3X1_778/A NOR3X1_778/C NOR3X1_778/B NOR3X1_777/A NOR3X1_709/C NOR3X1_710/A NOR3X1_710/B NOR3X1_1194/A NOR3X1_1193/B NOR3X1_1194/B NOR3X1_895/C NOR3X1_896/B NOR3X1_710/C NOR3X1_709/A NOR3X1_895/A NOR3X1_1268/B NOR3X1_1267/A NOR3X1_470/C NOR3X1_1626/C NOR3X1_1265/A NOR3X1_1266/B NOR3X1_1554/C NOR3X1_1553/A NOR3X1_1081/A NOR3X1_1555/A 
+ NOR3X1_1556/C NOR3X1_1338/A NOR3X1_1338/B NOR3X1_1518/A NOR3X1_1518/B NOR3X1_669/A NOR3X1_670/B NOR3X1_395/A NOR3X1_396/C NOR3X1_1224/C NOR3X1_1224/A NOR3X1_134/A NOR3X1_134/B NOR3X1_1244/A NOR3X1_1244/B NOR3X1_1243/C NOR3X1_1351/A NOR3X1_1352/C NOR3X1_522/A NOR3X1_522/B NOR3X1_1244/C NOR3X1_1243/A NOR3X1_781/A NOR3X1_782/C NOR3X1_1345/A NOR3X1_1346/B NOR3X1_927/B NOR3X1_928/B NOR3X1_927/A NOR3X1_928/A NOR3X1_928/C NOR3X1_917/C NOR3X1_1276/A NOR3X1_1276/B NOR3X1_649/C NOR3X1_650/A NOR3X1_650/B NOR3X1_1005/B NOR3X1_1551/C NOR3X1_1552/A NOR3X1_1552/B NOR3X1_335/C NOR3X1_336/A NOR3X1_336/B NOR3X1_615/C NOR3X1_616/A NOR3X1_616/B NOR3X1_1415/C NOR3X1_1416/A NOR3X1_1416/B NOR3X1_294/C 
+ NOR3X1_293/B NOR3X1_294/A NOR3X1_665/B NOR3X1_666/A NOR3X1_666/C NOR3X1_572/A NOR3X1_572/B NOR3X1_571/C NOR3X1_1407/B NOR3X1_1408/A NOR3X1_891/C NOR3X1_1408/C NOR3X1_892/A NOR3X1_892/B NOR3X1_669/C NOR3X1_453/B NOR3X1_454/A NOR3X1_454/C NOR3X1_650/C NOR3X1_649/A NOR3X1_1551/A NOR3X1_1552/C NOR3X1_335/A NOR3X1_336/C NOR3X1_615/A NOR3X1_616/C NOR3X1_293/A NOR3X1_294/B NOR3X1_1415/A NOR3X1_1416/C NOR3X1_811/B NOR3X1_1039/B NOR3X1_1040/A NOR3X1_1040/C NOR3X1_1351/B NOR3X1_391/B NOR3X1_392/A NOR3X1_392/C NOR3X1_1667/C NOR3X1_1668/A NOR3X1_1668/B NOR3X1_1557/C NOR3X1_1558/A NOR3X1_1558/B NOR3X1_1411/C NOR3X1_1538/A NOR3X1_1538/B NOR3X1_1675/A NOR3X1_1676/C NOR3X1_1069/A NOR3X1_1070/B 
+ NOR3X1_1011/A NOR3X1_1012/B NOR3X1_894/C NOR3X1_893/A NOR3X1_389/A NOR3X1_390/B NOR3X1_275/A NOR3X1_276/B NOR3X1_1696/B NOR3X1_1695/A NOR3X1_1695/B NOR3X1_1696/A NOR3X1_1696/C NOR3X1_1040/B NOR3X1_1039/A NOR3X1_391/A NOR3X1_392/B NOR3X1_1668/C NOR3X1_1558/C NOR3X1_1557/A NOR3X1_1667/A NOR3X1_1577/A NOR3X1_1578/C NOR3X1_1559/C NOR3X1_1560/A NOR3X1_1560/B NOR3X1_1661/C NOR3X1_1662/B NOR3X1_1664/A NOR3X1_1664/C NOR3X1_1663/B NOR3X1_1260/C NOR3X1_1259/A NOR3X1_1685/A NOR3X1_573/A NOR3X1_1686/B NOR3X1_574/C NOR3X1_1085/A NOR3X1_1086/B NOR3X1_604/B NOR3X1_603/A NOR3X1_601/A NOR3X1_602/B NOR3X1_1661/A NOR3X1_1560/C NOR3X1_1559/A NOR3X1_1664/B NOR3X1_1663/A NOR3X1_453/A NOR3X1_454/B NOR3X1_891/A 
+ NOR3X1_1408/B NOR3X1_892/C NOR3X1_1407/A NOR3X1_665/A NOR3X1_666/B NOR3X1_572/C NOR3X1_571/A NOR3X1_1261/A NOR3X1_1262/B NOR3X1_1617/C NOR3X1_1618/C NOR3X1_1617/A NOR3X1_668/B NOR3X1_667/A NOR3X1_1671/A NOR3X1_1672/B NOR3X1_479/A NOR3X1_480/B NOR3X1_1458/B NOR3X1_1457/A NOR3X1_1710/C NOR3X1_1709/A NOR3X1_1709/C NOR3X1_1457/B NOR3X1_649/B NOR3X1_1094/C NOR3X1_1093/A NOR3X1_1093/C NOR3X1_1094/A NOR3X1_1094/B NOR3X1_664/A NOR3X1_664/B NOR3X1_663/C NOR3X1_664/C NOR3X1_663/A NOR3X1_1031/A NOR3X1_1032/C NOR3X1_1458/C NOR3X1_1710/A NOR3X1_1710/B NOR3X1_1458/A NOR3X1_1031/B NOR3X1_721/A NOR3X1_721/B NOR3X1_722/B NOR3X1_945/A NOR3X1_945/B NOR3X1_946/B NOR3X1_722/A NOR3X1_722/C NOR3X1_946/A 
+ NOR3X1_946/C NOR3X1_1618/A NOR3X1_1618/B INVX1_1198/Y INVX1_1197/Y INVX1_176/Y INVX1_175/Y INVX1_131/Y INVX1_132/Y INVX1_747/Y INVX1_748/Y INVX1_239/Y INVX1_240/Y INVX1_653/Y INVX1_654/Y INVX1_1198/A INVX1_548/A INVX1_547/A INVX1_1197/A INVX1_176/A INVX1_175/A INVX1_822/A INVX1_821/A INVX1_1377/A INVX1_1378/A INVX1_131/A INVX1_132/A INVX1_747/A INVX1_748/A INVX1_1640/A INVX1_1639/A INVX1_239/A INVX1_240/A INVX1_653/A INVX1_654/A INVX1_750/A INVX1_749/A INVX1_1060/A INVX1_1059/A INVX1_369/A INVX1_370/A NOR3X1_175/B NOR3X1_821/B NOR3X1_747/B NOR3X1_653/B INVX1_174/Y INVX1_173/Y INVX1_820/Y INVX1_819/Y INVX1_1520/Y INVX1_1519/Y 
+ INVX1_537/Y INVX1_538/Y INVX1_745/Y INVX1_746/Y INVX1_528/Y INVX1_527/Y INVX1_174/A INVX1_173/A INVX1_820/A INVX1_819/A INVX1_1520/A INVX1_1519/A INVX1_537/A INVX1_539/A INVX1_540/A INVX1_538/A INVX1_745/A INVX1_746/A INVX1_528/A INVX1_527/A NOR3X1_1519/B INVX1_1370/Y INVX1_1372/Y INVX1_1371/Y INVX1_1369/Y INVX1_1370/A INVX1_1372/A INVX1_1371/A INVX1_1369/A NOR3X1_1371/C NOR3X1_1369/B INVX1_1364/Y INVX1_1363/Y INVX1_1366/Y INVX1_1365/Y INVX1_1364/A INVX1_1363/A INVX1_1366/A INVX1_1365/A INVX1_855/Y INVX1_856/Y INVX1_1508/Y INVX1_1507/Y INVX1_376/Y INVX1_375/Y INVX1_372/Y INVX1_1063/Y INVX1_371/Y INVX1_1064/Y INVX1_1327/Y INVX1_1216/Y 
+ INVX1_1215/Y INVX1_1328/Y INVX1_766/Y INVX1_765/Y INVX1_259/Y INVX1_260/Y INVX1_1354/Y INVX1_1353/Y INVX1_156/Y INVX1_155/Y INVX1_311/Y INVX1_312/Y INVX1_498/Y INVX1_497/Y INVX1_1227/Y INVX1_1228/Y INVX1_1179/Y INVX1_1180/Y INVX1_1656/Y INVX1_1655/Y INVX1_1511/Y INVX1_1512/Y INVX1_209/Y INVX1_210/Y INVX1_493/Y INVX1_494/Y INVX1_302/Y INVX1_301/Y INVX1_323/Y INVX1_324/Y INVX1_1062/Y INVX1_1061/Y INVX1_1396/Y INVX1_1395/Y INVX1_524/Y INVX1_523/Y INVX1_580/Y INVX1_579/Y INVX1_610/Y INVX1_609/Y INVX1_236/Y INVX1_235/Y INVX1_393/Y INVX1_394/Y INVX1_992/Y INVX1_991/Y INVX1_1340/Y INVX1_1339/Y INVX1_1673/Y INVX1_1674/Y INVX1_82/Y 
+ INVX1_81/Y INVX1_478/Y INVX1_477/Y INVX1_840/Y INVX1_839/Y INVX1_1065/Y INVX1_1066/Y INVX1_270/Y INVX1_269/Y INVX1_1172/Y INVX1_1171/Y INVX1_965/Y INVX1_966/Y INVX1_192/Y INVX1_191/Y INVX1_1257/Y INVX1_1258/Y INVX1_150/Y INVX1_149/Y INVX1_596/Y INVX1_595/Y INVX1_630/Y INVX1_629/Y INVX1_1335/Y INVX1_1336/Y INVX1_496/Y INVX1_495/Y INVX1_502/Y INVX1_501/Y INVX1_567/Y INVX1_568/Y INVX1_832/Y INVX1_831/Y INVX1_508/Y INVX1_507/Y INVX1_758/Y INVX1_757/Y INVX1_1502/Y INVX1_1501/Y INVX1_520/Y INVX1_519/Y INVX1_977/Y INVX1_978/Y INVX1_197/Y INVX1_198/Y INVX1_1219/Y INVX1_1220/Y INVX1_768/Y INVX1_767/Y INVX1_1516/Y INVX1_1515/Y 
+ INVX1_1646/Y INVX1_1645/Y INVX1_463/Y INVX1_464/Y INVX1_1274/Y INVX1_1273/Y INVX1_759/Y INVX1_760/Y INVX1_1528/Y INVX1_1527/Y INVX1_103/Y INVX1_104/Y INVX1_854/Y INVX1_853/Y INVX1_1390/Y INVX1_1389/Y INVX1_770/Y INVX1_769/Y INVX1_662/Y INVX1_661/Y INVX1_1241/Y INVX1_1242/Y INVX1_913/Y INVX1_914/Y INVX1_476/Y INVX1_475/Y INVX1_330/Y INVX1_329/Y INVX1_613/Y INVX1_614/Y INVX1_1394/Y INVX1_1393/Y INVX1_283/Y INVX1_284/Y INVX1_342/Y INVX1_341/Y INVX1_569/Y INVX1_570/Y INVX1_626/Y INVX1_625/Y INVX1_836/Y INVX1_835/Y INVX1_974/Y INVX1_973/Y INVX1_448/Y INVX1_447/Y INVX1_1036/Y INVX1_1035/Y INVX1_90/Y INVX1_89/Y INVX1_1691/Y 
+ INVX1_1692/Y INVX1_308/Y INVX1_307/Y INVX1_1488/Y INVX1_1487/Y INVX1_864/Y INVX1_846/Y INVX1_845/Y INVX1_863/Y INVX1_1603/Y INVX1_1604/Y INVX1_1658/Y INVX1_1657/Y INVX1_1056/Y INVX1_1055/Y INVX1_218/Y INVX1_217/Y INVX1_534/Y INVX1_533/Y INVX1_232/Y INVX1_231/Y INVX1_855/A INVX1_856/A INVX1_1508/A INVX1_1507/A INVX1_376/A INVX1_375/A INVX1_372/A INVX1_1063/A INVX1_371/A INVX1_1064/A INVX1_1327/A INVX1_1216/A INVX1_1215/A INVX1_1328/A INVX1_766/A INVX1_765/A INVX1_259/A INVX1_260/A INVX1_1354/A INVX1_1353/A INVX1_156/A INVX1_155/A INVX1_311/A INVX1_312/A INVX1_498/A INVX1_497/A INVX1_1227/A INVX1_1228/A INVX1_1179/A INVX1_1180/A 
+ INVX1_1656/A INVX1_1655/A INVX1_1511/A INVX1_1512/A INVX1_209/A INVX1_210/A INVX1_493/A INVX1_494/A INVX1_302/A INVX1_301/A INVX1_323/A INVX1_324/A INVX1_1062/A INVX1_1061/A INVX1_1396/A INVX1_1395/A INVX1_524/A INVX1_523/A INVX1_580/A INVX1_579/A INVX1_610/A INVX1_609/A INVX1_236/A INVX1_235/A INVX1_393/A INVX1_394/A INVX1_992/A INVX1_991/A INVX1_1340/A INVX1_1339/A INVX1_1673/A INVX1_1674/A INVX1_82/A INVX1_81/A INVX1_478/A INVX1_477/A INVX1_840/A INVX1_839/A INVX1_1065/A INVX1_1066/A INVX1_270/A INVX1_269/A INVX1_1172/A INVX1_1171/A INVX1_965/A INVX1_966/A INVX1_192/A INVX1_191/A INVX1_1257/A INVX1_1258/A INVX1_150/A 
+ INVX1_149/A INVX1_596/A INVX1_595/A INVX1_630/A INVX1_629/A INVX1_1335/A INVX1_1336/A INVX1_496/A INVX1_495/A INVX1_502/A INVX1_501/A INVX1_567/A INVX1_568/A INVX1_832/A INVX1_831/A INVX1_508/A INVX1_507/A INVX1_758/A INVX1_757/A INVX1_1502/A INVX1_1501/A INVX1_520/A INVX1_519/A INVX1_977/A INVX1_978/A INVX1_197/A INVX1_198/A INVX1_1219/A INVX1_1220/A INVX1_768/A INVX1_767/A INVX1_1516/A INVX1_1515/A INVX1_1646/A INVX1_1645/A INVX1_463/A INVX1_464/A INVX1_1274/A INVX1_1273/A INVX1_759/A INVX1_760/A INVX1_1528/A INVX1_1527/A INVX1_103/A INVX1_104/A INVX1_854/A INVX1_853/A INVX1_1390/A INVX1_1389/A INVX1_770/A INVX1_769/A 
+ INVX1_662/A INVX1_661/A INVX1_1241/A INVX1_1242/A INVX1_913/A INVX1_914/A INVX1_476/A INVX1_475/A INVX1_330/A INVX1_329/A INVX1_613/A INVX1_614/A INVX1_1394/A INVX1_1393/A INVX1_283/A INVX1_284/A INVX1_342/A INVX1_341/A INVX1_569/A INVX1_570/A INVX1_626/A INVX1_625/A INVX1_836/A INVX1_835/A INVX1_974/A INVX1_973/A INVX1_448/A INVX1_447/A INVX1_1036/A INVX1_1035/A INVX1_90/A INVX1_89/A INVX1_1691/A INVX1_1692/A INVX1_308/A INVX1_307/A INVX1_1488/A INVX1_1487/A INVX1_864/A INVX1_846/A INVX1_845/A INVX1_863/A INVX1_1603/A INVX1_1604/A INVX1_1658/A INVX1_1657/A INVX1_1056/A INVX1_1055/A INVX1_218/A INVX1_217/A INVX1_534/A 
+ INVX1_533/A NOR3X1_1507/B NOR3X1_375/B NOR3X1_371/B NOR3X1_311/C NOR3X1_393/C NOR3X1_1065/B NOR3X1_495/B NOR3X1_501/B NOR3X1_977/C NOR3X1_197/C NOR3X1_767/B NOR3X1_1273/B NOR3X1_759/B NOR3X1_613/B NOR3X1_1603/A NOR3X1_1603/B NOR3X1_1603/C NOR3X1_1604/A NOR3X1_1604/B NOR3X1_1604/C NOR3X1_1657/B NOR3X1_232/A NOR3X1_232/B NOR3X1_232/C NOR3X1_231/A NOR3X1_231/B NOR3X1_231/C INVX1_320/Y INVX1_322/Y INVX1_321/Y INVX1_319/Y INVX1_1649/Y INVX1_1651/Y INVX1_1652/Y INVX1_1650/Y INVX1_503/Y INVX1_963/Y INVX1_964/Y INVX1_504/Y INVX1_1251/Y INVX1_1253/Y INVX1_1254/Y INVX1_1252/Y INVX1_557/Y INVX1_559/Y INVX1_560/Y INVX1_558/Y INVX1_506/Y INVX1_505/Y INVX1_194/Y 
+ INVX1_196/Y INVX1_195/Y INVX1_193/Y INVX1_660/Y INVX1_659/Y INVX1_1231/Y INVX1_1233/Y INVX1_1234/Y INVX1_1232/Y INVX1_735/Y INVX1_740/Y INVX1_739/Y INVX1_736/Y INVX1_561/Y INVX1_563/Y INVX1_564/Y INVX1_562/Y INVX1_1629/Y INVX1_1631/Y INVX1_1632/Y INVX1_1630/Y INVX1_1596/Y INVX1_1598/Y INVX1_1597/Y INVX1_1595/Y INVX1_531/Y INVX1_530/Y INVX1_532/Y INVX1_529/Y INVX1_229/Y INVX1_227/Y INVX1_230/Y INVX1_228/Y INVX1_320/A INVX1_322/A INVX1_321/A INVX1_319/A INVX1_1649/A INVX1_1651/A INVX1_1652/A INVX1_1650/A INVX1_503/A INVX1_963/A INVX1_964/A INVX1_504/A INVX1_1251/A INVX1_1253/A INVX1_1254/A INVX1_1252/A INVX1_557/A INVX1_559/A 
+ INVX1_560/A INVX1_558/A INVX1_506/A INVX1_505/A INVX1_194/A INVX1_196/A INVX1_195/A INVX1_193/A INVX1_660/A INVX1_659/A INVX1_1231/A INVX1_1233/A INVX1_1234/A INVX1_1232/A INVX1_735/A INVX1_740/A INVX1_739/A INVX1_736/A INVX1_561/A INVX1_563/A INVX1_564/A INVX1_562/A INVX1_1629/A INVX1_1631/A INVX1_1632/A INVX1_1630/A INVX1_531/A INVX1_530/A INVX1_532/A INVX1_529/A INVX1_229/A INVX1_227/A INVX1_230/A INVX1_228/A NOR3X1_195/B NOR3X1_735/B NOR3X1_1631/B NOR3X1_1596/A NOR3X1_1596/B NOR3X1_1596/C NOR3X1_1598/A NOR3X1_1598/B NOR3X1_1598/C NOR3X1_1597/A NOR3X1_1597/B NOR3X1_1595/A NOR3X1_1595/B NOR3X1_531/C NOR3X1_529/B NOR3X1_227/B INVX1_182/Y 
+ INVX1_178/Y INVX1_181/Y INVX1_177/Y INVX1_871/Y INVX1_637/Y INVX1_872/Y INVX1_638/Y INVX1_1185/Y INVX1_1077/Y INVX1_1186/Y INVX1_1078/Y INVX1_211/Y INVX1_224/Y INVX1_223/Y INVX1_212/Y INVX1_215/Y INVX1_226/Y INVX1_225/Y INVX1_216/Y INVX1_182/A INVX1_178/A INVX1_181/A INVX1_177/A INVX1_871/A INVX1_872/A INVX1_1185/A INVX1_1186/A INVX1_211/A INVX1_224/A INVX1_223/A INVX1_212/A INVX1_215/A INVX1_226/A INVX1_225/A INVX1_216/A NOR3X1_871/C NOR3X1_637/A NOR3X1_637/B NOR3X1_637/C NOR3X1_638/A NOR3X1_638/B NOR3X1_638/C NOR3X1_1185/B NOR3X1_1077/A NOR3X1_1077/B NOR3X1_1077/C NOR3X1_1078/A NOR3X1_1078/B NOR3X1_1078/C NOR3X1_211/B NOR3X1_223/C 
+ INVX1_868/Y INVX1_870/Y INVX1_869/Y INVX1_867/Y INVX1_634/Y INVX1_636/Y INVX1_635/Y INVX1_633/Y INVX1_1181/Y INVX1_1184/Y INVX1_1183/Y INVX1_1182/Y INVX1_1074/Y INVX1_1076/Y INVX1_1075/Y INVX1_1073/Y INVX1_214/Y INVX1_206/Y INVX1_213/Y INVX1_205/Y INVX1_868/A INVX1_870/A INVX1_869/A INVX1_867/A INVX1_634/A INVX1_636/A INVX1_635/A INVX1_633/A INVX1_1181/A INVX1_1184/A INVX1_1183/A INVX1_1182/A INVX1_1074/A INVX1_1076/A INVX1_1075/A INVX1_1073/A INVX1_214/A INVX1_206/A INVX1_213/A INVX1_205/A NOR3X1_869/C NOR3X1_1181/B INVX1_862/Y INVX1_344/Y INVX1_861/Y INVX1_343/Y INVX1_628/Y INVX1_627/Y INVX1_632/Y INVX1_631/Y INVX1_1178/Y 
+ INVX1_1177/Y INVX1_1072/Y INVX1_1071/Y INVX1_622/Y INVX1_26/Y INVX1_621/Y INVX1_25/Y INVX1_862/A INVX1_344/A INVX1_861/A INVX1_343/A INVX1_628/A INVX1_627/A INVX1_632/A INVX1_631/A INVX1_1178/A INVX1_1177/A INVX1_1072/A INVX1_1071/A INVX1_622/A INVX1_26/A INVX1_621/A INVX1_25/A INVX1_370/Y INVX1_369/Y INVX1_540/Y INVX1_539/Y INVX1_1374/Y INVX1_1373/Y 
+ VSS VDD 
+ NOR3X1_1619/A NOR3X1_1619/B NOR3X1_1620/B NOR3X1_951/A NOR3X1_951/B NOR3X1_952/B NOR3X1_724/B NOR3X1_723/A NOR3X1_723/B NOR3X1_1577/B NOR3X1_952/A NOR3X1_952/C NOR3X1_724/A NOR3X1_724/C NOR3X1_1147/B NOR3X1_1148/B NOR3X1_1147/A NOR3X1_1459/A NOR3X1_1459/B NOR3X1_1460/B NOR3X1_1711/A NOR3X1_1711/B NOR3X1_1712/B NOR3X1_1148/A NOR3X1_1148/C NOR3X1_678/A NOR3X1_678/C NOR3X1_677/B NOR3X1_678/B NOR3X1_677/A NOR3X1_1429/C NOR3X1_1430/A NOR3X1_1430/B NOR3X1_1430/C NOR3X1_1429/A NOR3X1_1460/A NOR3X1_1460/C NOR3X1_1712/A NOR3X1_1712/C NOR3X1_485/A NOR3X1_485/B NOR3X1_486/B NOR3X1_486/A NOR3X1_486/C NOR3X1_675/B NOR3X1_676/A NOR3X1_676/C NOR3X1_675/A NOR3X1_676/B NOR3X1_1620/C NOR3X1_1620/A 
+ NOR3X1_1264/B NOR3X1_1263/A NOR3X1_1263/B NOR3X1_1264/A NOR3X1_1264/C NOR3X1_1275/B NOR3X1_1113/C NOR3X1_675/C NOR3X1_1427/B NOR3X1_1428/A NOR3X1_1428/C NOR3X1_907/C NOR3X1_908/C NOR3X1_907/A NOR3X1_1428/B NOR3X1_1427/A NOR3X1_908/A NOR3X1_908/B NOR3X1_679/A NOR3X1_679/B NOR3X1_680/B NOR3X1_680/A NOR3X1_680/C NOR3X1_1681/B NOR3X1_1682/A NOR3X1_1682/C NOR3X1_1681/A NOR3X1_1682/B NOR3X1_1565/B NOR3X1_1566/A NOR3X1_1566/C NOR3X1_1565/A NOR3X1_1566/B NOR3X1_1681/C NOR3X1_1431/A NOR3X1_1431/B NOR3X1_1432/B NOR3X1_1432/A NOR3X1_1432/C NOR3X1_1103/B NOR3X1_1104/B NOR3X1_1103/A NOR3X1_1104/A NOR3X1_1104/C NOR3X1_1573/C NOR3X1_1574/A NOR3X1_1574/B NOR3X1_1699/B NOR3X1_1700/B NOR3X1_1699/A NOR3X1_1700/A 
+ NOR3X1_1700/C NOR3X1_1263/C NOR3X1_315/C NOR3X1_1586/C NOR3X1_1585/A NOR3X1_1585/C NOR3X1_1586/B NOR3X1_1586/A NOR3X1_1679/B NOR3X1_1680/A NOR3X1_1680/C NOR3X1_1565/C NOR3X1_1679/A NOR3X1_1680/B NOR3X1_398/B NOR3X1_397/A NOR3X1_397/B NOR3X1_398/C NOR3X1_398/A NOR3X1_1283/B NOR3X1_1117/B NOR3X1_1118/A NOR3X1_1118/C NOR3X1_1284/A NOR3X1_1284/C NOR3X1_1283/A NOR3X1_1118/B NOR3X1_1117/A NOR3X1_1284/B NOR3X1_1717/C NOR3X1_1718/C NOR3X1_1717/A NOR3X1_1718/A NOR3X1_1718/B NOR3X1_277/B NOR3X1_278/B NOR3X1_277/A NOR3X1_278/A NOR3X1_278/C NOR3X1_397/C NOR3X1_907/B NOR3X1_1134/C NOR3X1_1133/A NOR3X1_1133/C NOR3X1_1134/A NOR3X1_1134/B NOR3X1_1704/C NOR3X1_1703/A NOR3X1_1703/C NOR3X1_1704/A NOR3X1_1704/B 
+ NOR3X1_1425/B NOR3X1_1426/A NOR3X1_1426/C NOR3X1_1287/A NOR3X1_1287/B NOR3X1_1288/B NOR3X1_1467/A NOR3X1_950/C NOR3X1_1467/C NOR3X1_1468/C NOR3X1_949/A NOR3X1_949/C NOR3X1_1424/B NOR3X1_1423/A NOR3X1_1423/B NOR3X1_1424/A NOR3X1_1424/C NOR3X1_1454/C NOR3X1_1453/A NOR3X1_1453/C NOR3X1_705/A NOR3X1_705/B NOR3X1_706/B NOR3X1_706/A NOR3X1_706/C NOR3X1_1454/A NOR3X1_1454/B NOR3X1_340/C NOR3X1_339/A NOR3X1_339/C NOR3X1_340/A NOR3X1_340/B NOR3X1_1569/A NOR3X1_1569/B NOR3X1_1570/B NOR3X1_1570/A NOR3X1_1570/C NOR3X1_1434/C NOR3X1_1433/A NOR3X1_1433/C NOR3X1_1434/A NOR3X1_1434/B NOR3X1_674/A NOR3X1_674/B NOR3X1_673/C NOR3X1_1573/A NOR3X1_1574/C NOR3X1_1301/A NOR3X1_1301/C NOR3X1_1302/C NOR3X1_941/A 
+ NOR3X1_941/C NOR3X1_942/C NOR3X1_942/A NOR3X1_942/B NOR3X1_1247/C NOR3X1_1248/A NOR3X1_1248/B NOR3X1_1248/C NOR3X1_1247/A NOR3X1_1347/B NOR3X1_1533/B NOR3X1_157/B NOR3X1_1229/B NOR3X1_1033/B NOR3X1_1333/B NOR3X1_404/A NOR3X1_404/B NOR3X1_403/C NOR3X1_415/A NOR3X1_415/B NOR3X1_416/B NOR3X1_416/A NOR3X1_416/C NOR3X1_674/C NOR3X1_673/A NOR3X1_1583/C NOR3X1_1584/A NOR3X1_1584/B NOR3X1_1513/B NOR3X1_1568/B NOR3X1_1567/A NOR3X1_1567/B NOR3X1_1568/A NOR3X1_1568/C NOR3X1_303/B NOR3X1_373/B NOR3X1_1187/B NOR3X1_1359/B NOR3X1_1105/B NOR3X1_1106/A NOR3X1_1106/C NOR3X1_1509/B NOR3X1_1329/B NOR3X1_1217/B NOR3X1_1331/B NOR3X1_499/B NOR3X1_1189/B NOR3X1_995/B NOR3X1_377/B NOR3X1_1567/C NOR3X1_1279/A 
+ NOR3X1_1279/C NOR3X1_1280/C NOR3X1_1280/A NOR3X1_1280/B NOR3X1_919/C NOR3X1_261/B NOR3X1_987/B NOR3X1_485/C NOR3X1_1279/B NOR3X1_905/C NOR3X1_906/A NOR3X1_906/B NOR3X1_711/B NOR3X1_712/A NOR3X1_712/C NOR3X1_711/A NOR3X1_712/B NOR3X1_905/A NOR3X1_906/C NOR3X1_1287/C NOR3X1_1288/A NOR3X1_1288/C NOR3X1_1423/C NOR3X1_615/B NOR3X1_395/B NOR3X1_1585/B NOR3X1_1437/B NOR3X1_1438/A NOR3X1_1438/C NOR3X1_407/C NOR3X1_408/A NOR3X1_408/B NOR3X1_1555/B NOR3X1_1093/B NOR3X1_391/C NOR3X1_1559/B NOR3X1_361/B NOR3X1_362/A NOR3X1_362/C NOR3X1_387/B NOR3X1_388/A NOR3X1_388/C NOR3X1_1579/B NOR3X1_1557/B NOR3X1_1415/B NOR3X1_479/C NOR3X1_1283/C NOR3X1_923/C NOR3X1_419/C NOR3X1_420/A NOR3X1_420/B 
+ NOR3X1_361/C NOR3X1_362/B NOR3X1_1302/A NOR3X1_1302/B NOR3X1_280/C NOR3X1_279/B NOR3X1_280/A NOR3X1_385/B NOR3X1_386/A NOR3X1_386/C NOR3X1_521/B NOR3X1_679/C NOR3X1_1553/B NOR3X1_1437/C NOR3X1_1438/B NOR3X1_387/C NOR3X1_388/B NOR3X1_385/C NOR3X1_386/B NOR3X1_1117/C NOR3X1_603/C NOR3X1_1085/C NOR3X1_1269/C NOR3X1_901/C NOR3X1_453/C NOR3X1_1087/B NOR3X1_1088/A NOR3X1_1088/C NOR3X1_1265/C NOR3X1_1349/A NOR3X1_1349/B NOR3X1_1350/B NOR3X1_349/C NOR3X1_350/A NOR3X1_350/B NOR3X1_1350/C NOR3X1_1350/A NOR3X1_360/C NOR3X1_359/B NOR3X1_360/A NOR3X1_1407/C NOR3X1_405/C NOR3X1_406/A NOR3X1_406/B NOR3X1_899/B NOR3X1_1001/C NOR3X1_1002/A NOR3X1_1002/B NOR3X1_1001/A NOR3X1_1002/C NOR3X1_401/B 
+ NOR3X1_402/A NOR3X1_402/C NOR3X1_1709/B NOR3X1_1435/C NOR3X1_1436/A NOR3X1_1436/B NOR3X1_1663/C NOR3X1_1417/C NOR3X1_293/C NOR3X1_1039/C NOR3X1_1468/A NOR3X1_1468/B NOR3X1_950/A NOR3X1_950/B NOR3X1_1575/C NOR3X1_1576/A NOR3X1_1576/B NOR3X1_1069/C NOR3X1_1305/C NOR3X1_1306/A NOR3X1_1306/B NOR3X1_893/B NOR3X1_384/A NOR3X1_384/B NOR3X1_383/C NOR3X1_1671/C NOR3X1_1551/B NOR3X1_335/B NOR3X1_933/C NOR3X1_420/C NOR3X1_419/B NOR3X1_934/A NOR3X1_934/B NOR3X1_891/B NOR3X1_1011/C NOR3X1_484/A NOR3X1_484/B NOR3X1_483/C NOR3X1_1685/C NOR3X1_1090/C NOR3X1_1089/B NOR3X1_1090/A NOR3X1_1451/C NOR3X1_1452/A NOR3X1_1452/B NOR3X1_417/B NOR3X1_418/A NOR3X1_418/C NOR3X1_683/B NOR3X1_1564/A NOR3X1_1564/B 
+ NOR3X1_1563/C NOR3X1_1107/C NOR3X1_1108/A NOR3X1_1108/B NOR3X1_1413/B NOR3X1_1345/C NOR3X1_1537/B NOR3X1_1572/A NOR3X1_1572/C NOR3X1_1571/B NOR3X1_1089/C NOR3X1_1090/B NOR3X1_665/C NOR3X1_1097/C NOR3X1_781/B NOR3X1_389/C NOR3X1_1223/C NOR3X1_1281/B NOR3X1_1282/A NOR3X1_1282/C NOR3X1_1517/B NOR3X1_601/C NOR3X1_275/C NOR3X1_663/B NOR3X1_1337/B NOR3X1_1267/C NOR3X1_667/C NOR3X1_1285/B NOR3X1_1286/A NOR3X1_1286/C NOR3X1_359/C NOR3X1_360/B NOR3X1_133/B NOR3X1_777/C NOR3X1_1667/B NOR3X1_1355/B NOR3X1_1087/C NOR3X1_1088/B NOR3X1_359/A NOR3X1_1089/A NOR3X1_1564/C NOR3X1_1563/A NOR3X1_387/A NOR3X1_1583/A NOR3X1_1584/C NOR3X1_404/C NOR3X1_403/A NOR3X1_361/A NOR3X1_484/C NOR3X1_483/A NOR3X1_1087/A 
+ NOR3X1_431/A NOR3X1_1311/A NOR3X1_431/C NOR3X1_1311/C NOR3X1_432/C NOR3X1_1312/C NOR3X1_432/A NOR3X1_432/B NOR3X1_1312/A NOR3X1_1312/B NOR3X1_1121/A NOR3X1_1121/C NOR3X1_1122/C NOR3X1_696/C NOR3X1_695/A NOR3X1_695/C NOR3X1_1122/A NOR3X1_1122/B NOR3X1_385/A NOR3X1_696/A NOR3X1_696/B NOR3X1_697/A NOR3X1_697/C NOR3X1_698/C NOR3X1_698/A NOR3X1_698/B NOR3X1_247/C NOR3X1_248/A NOR3X1_248/B NOR3X1_248/C NOR3X1_247/A NOR3X1_1110/C NOR3X1_1109/B NOR3X1_1110/A NOR3X1_1109/A NOR3X1_1110/B NOR3X1_1105/A NOR3X1_1106/B NOR3X1_693/C NOR3X1_694/A NOR3X1_694/B NOR3X1_693/A NOR3X1_694/C NOR3X1_403/B NOR3X1_405/A NOR3X1_406/C NOR3X1_350/C NOR3X1_349/A NOR3X1_401/A NOR3X1_402/B NOR3X1_1572/B 
+ NOR3X1_1571/A NOR3X1_1425/A NOR3X1_1426/B NOR3X1_1130/C NOR3X1_1129/A NOR3X1_1129/C NOR3X1_1130/A NOR3X1_1130/B NOR3X1_933/A NOR3X1_419/A NOR3X1_934/C NOR3X1_1451/A NOR3X1_1452/C NOR3X1_418/B NOR3X1_417/A NOR3X1_1107/A NOR3X1_1108/C NOR3X1_1435/A NOR3X1_1436/C NOR3X1_1285/A NOR3X1_1286/B NOR3X1_1282/B NOR3X1_1281/A NOR3X1_1437/A NOR3X1_408/C NOR3X1_407/A NOR3X1_279/A NOR3X1_280/B NOR3X1_1305/A NOR3X1_1306/C NOR3X1_1576/C NOR3X1_1575/A NOR3X1_384/C NOR3X1_383/A INVX1_965/Y INVX1_966/Y INVX1_534/Y INVX1_533/Y INVX1_323/A INVX1_324/A INVX1_1673/A INVX1_1674/A INVX1_965/A INVX1_966/A 
+ INVX1_1257/A INVX1_1258/A INVX1_567/A INVX1_568/A INVX1_508/A INVX1_507/A INVX1_197/A INVX1_198/A INVX1_662/A INVX1_661/A INVX1_1241/A INVX1_1242/A INVX1_913/A INVX1_914/A INVX1_569/A INVX1_570/A INVX1_1691/A INVX1_1692/A INVX1_534/A INVX1_533/A NOR3X1_197/C NOR3X1_232/A NOR3X1_232/B NOR3X1_232/C NOR3X1_231/A NOR3X1_231/B NOR3X1_231/C INVX1_194/Y INVX1_193/Y INVX1_229/Y INVX1_227/Y INVX1_230/Y INVX1_228/Y INVX1_194/A INVX1_193/A INVX1_229/A INVX1_227/A INVX1_230/A INVX1_228/A NOR3X1_1596/A NOR3X1_1596/B NOR3X1_1596/C NOR3X1_1598/A NOR3X1_1598/B NOR3X1_1598/C NOR3X1_1597/A NOR3X1_1597/B NOR3X1_1595/A NOR3X1_1595/B NOR3X1_227/B INVX1_871/Y 
+ INVX1_872/Y INVX1_226/Y INVX1_225/Y INVX1_871/A INVX1_872/A INVX1_1185/A INVX1_1186/A INVX1_226/A INVX1_225/A NOR3X1_871/C NOR3X1_637/A NOR3X1_637/B NOR3X1_637/C NOR3X1_638/A NOR3X1_638/B NOR3X1_638/C NOR3X1_1185/B NOR3X1_1077/A NOR3X1_1077/B NOR3X1_1077/C NOR3X1_1078/A NOR3X1_1078/B NOR3X1_1078/C INVX1_868/Y INVX1_867/Y INVX1_634/Y INVX1_636/Y INVX1_635/Y INVX1_633/Y INVX1_1184/Y INVX1_1183/Y INVX1_1074/Y INVX1_1076/Y INVX1_1075/Y INVX1_1073/Y INVX1_868/A INVX1_867/A INVX1_634/A INVX1_636/A INVX1_635/A INVX1_633/A INVX1_1184/A INVX1_1183/A INVX1_1074/A INVX1_1076/A INVX1_1075/A INVX1_1073/A INVX1_1548/Y INVX1_1547/Y INVX1_944/Y INVX1_943/Y 
+ INVX1_575/Y INVX1_576/Y INVX1_1019/Y INVX1_1020/Y INVX1_1456/Y INVX1_1455/Y INVX1_1708/Y INVX1_1707/Y INVX1_121/Y INVX1_122/Y INVX1_1403/Y INVX1_1404/Y INVX1_1092/Y INVX1_1091/Y INVX1_647/Y INVX1_648/Y INVX1_1669/Y INVX1_1670/Y INVX1_1535/Y INVX1_1536/Y INVX1_1405/Y INVX1_1406/Y INVX1_456/Y INVX1_455/Y INVX1_1083/Y INVX1_1084/Y INVX1_971/Y INVX1_972/Y INVX1_1683/Y INVX1_1684/Y INVX1_1665/Y INVX1_1666/Y INVX1_1697/Y INVX1_1698/Y INVX1_273/Y INVX1_274/Y INVX1_1014/Y INVX1_1013/Y INVX1_651/Y INVX1_652/Y INVX1_1677/Y INVX1_1678/Y INVX1_1540/Y INVX1_1539/Y INVX1_1409/Y INVX1_1410/Y INVX1_1442/Y INVX1_947/Y INVX1_1441/Y INVX1_948/Y INVX1_295/Y 
+ INVX1_296/Y INVX1_887/Y INVX1_888/Y INVX1_606/Y INVX1_605/Y INVX1_337/Y INVX1_338/Y INVX1_1550/Y INVX1_1549/Y INVX1_985/Y INVX1_986/Y INVX1_671/Y INVX1_672/Y INVX1_1278/Y INVX1_1277/Y INVX1_930/Y INVX1_929/Y INVX1_1440/Y INVX1_1439/Y INVX1_779/Y INVX1_780/Y INVX1_1245/Y INVX1_1246/Y INVX1_517/Y INVX1_518/Y INVX1_1291/Y INVX1_1292/Y INVX1_70/Y INVX1_69/Y INVX1_1581/Y INVX1_1582/Y INVX1_1079/Y INVX1_1080/Y INVX1_897/Y INVX1_898/Y INVX1_707/Y INVX1_708/Y INVX1_776/Y INVX1_775/Y INVX1_1271/Y INVX1_1272/Y INVX1_167/Y INVX1_168/Y INVX1_1046/Y INVX1_997/Y INVX1_998/Y INVX1_1045/Y INVX1_1239/Y INVX1_1240/Y INVX1_256/Y INVX1_255/Y 
+ INVX1_1543/Y INVX1_1544/Y INVX1_801/Y INVX1_802/Y INVX1_878/Y INVX1_877/Y INVX1_347/Y INVX1_348/Y INVX1_151/Y INVX1_152/Y INVX1_999/Y INVX1_1000/Y INVX1_1209/Y INVX1_1210/Y INVX1_1203/Y INVX1_1204/Y INVX1_1303/Y INVX1_1304/Y INVX1_1659/Y INVX1_1660/Y INVX1_381/Y INVX1_382/Y INVX1_1358/Y INVX1_1357/Y INVX1_903/Y INVX1_904/Y INVX1_481/Y INVX1_482/Y INVX1_1421/Y INVX1_1422/Y INVX1_297/Y INVX1_298/Y INVX1_1561/Y INVX1_1562/Y INVX1_885/Y INVX1_886/Y INVX1_379/Y INVX1_380/Y INVX1_461/Y INVX1_462/Y INVX1_1294/Y INVX1_1293/Y INVX1_1116/Y INVX1_1115/Y INVX1_689/Y INVX1_690/Y INVX1_925/Y INVX1_926/Y INVX1_686/Y INVX1_685/Y INVX1_245/Y 
+ INVX1_246/Y INVX1_799/Y INVX1_800/Y INVX1_691/Y INVX1_692/Y INVX1_1420/Y INVX1_1419/Y INVX1_1099/Y INVX1_1100/Y INVX1_944/A INVX1_943/A INVX1_575/A INVX1_576/A INVX1_1456/A INVX1_1455/A INVX1_1708/A INVX1_1707/A INVX1_121/A INVX1_122/A INVX1_1403/A INVX1_1404/A INVX1_1092/A INVX1_1091/A INVX1_647/A INVX1_648/A INVX1_1669/A INVX1_1670/A INVX1_1535/A INVX1_1536/A INVX1_1405/A INVX1_1406/A INVX1_456/A INVX1_455/A INVX1_1083/A INVX1_1084/A INVX1_971/A INVX1_972/A INVX1_1683/A INVX1_1684/A INVX1_1665/A INVX1_1666/A INVX1_273/A INVX1_274/A INVX1_1014/A INVX1_1013/A INVX1_651/A INVX1_652/A INVX1_1677/A INVX1_1678/A INVX1_1540/A INVX1_1539/A 
+ INVX1_1409/A INVX1_1410/A INVX1_1442/A INVX1_1441/A INVX1_295/A INVX1_296/A INVX1_887/A INVX1_888/A INVX1_606/A INVX1_605/A INVX1_337/A INVX1_338/A INVX1_1550/A INVX1_1549/A INVX1_985/A INVX1_986/A INVX1_671/A INVX1_672/A INVX1_1278/A INVX1_1277/A INVX1_1440/A INVX1_1439/A INVX1_779/A INVX1_780/A INVX1_1245/A INVX1_1246/A INVX1_517/A INVX1_518/A INVX1_1291/A INVX1_1292/A INVX1_1581/A INVX1_1582/A INVX1_1079/A INVX1_1080/A INVX1_897/A INVX1_898/A INVX1_776/A INVX1_775/A INVX1_1271/A INVX1_1272/A INVX1_167/A INVX1_168/A INVX1_1046/A INVX1_997/A INVX1_998/A INVX1_1045/A INVX1_1239/A INVX1_1240/A INVX1_256/A INVX1_255/A INVX1_1543/A 
+ INVX1_1544/A INVX1_801/A INVX1_802/A INVX1_878/A INVX1_877/A INVX1_347/A INVX1_348/A INVX1_151/A INVX1_152/A INVX1_999/A INVX1_1000/A INVX1_1209/A INVX1_1210/A INVX1_1203/A INVX1_1204/A INVX1_1659/A INVX1_1660/A INVX1_381/A INVX1_382/A INVX1_1358/A INVX1_1357/A INVX1_903/A INVX1_904/A INVX1_481/A INVX1_482/A INVX1_1421/A INVX1_1422/A INVX1_297/A INVX1_298/A INVX1_1561/A INVX1_1562/A INVX1_885/A INVX1_886/A INVX1_379/A INVX1_380/A INVX1_461/A INVX1_462/A INVX1_1294/A INVX1_1293/A INVX1_1116/A INVX1_1115/A INVX1_689/A INVX1_690/A INVX1_925/A INVX1_926/A INVX1_686/A INVX1_685/A INVX1_245/A INVX1_246/A INVX1_799/A INVX1_800/A 
+ INVX1_691/A INVX1_692/A INVX1_1420/A INVX1_1419/A INVX1_1099/A INVX1_1100/A NOR3X1_1548/A NOR3X1_1548/B NOR3X1_1548/C NOR3X1_1547/A NOR3X1_1547/B NOR3X1_1547/C NOR3X1_943/B NOR3X1_1019/A NOR3X1_1019/B NOR3X1_1019/C NOR3X1_1020/A NOR3X1_1020/B NOR3X1_1020/C NOR3X1_1455/C NOR3X1_1707/C NOR3X1_1683/B NOR3X1_1697/A NOR3X1_1697/B NOR3X1_1697/C NOR3X1_1698/A NOR3X1_1698/B NOR3X1_1698/C NOR3X1_651/C NOR3X1_1677/C NOR3X1_947/A NOR3X1_947/C NOR3X1_1441/B NOR3X1_948/A NOR3X1_948/B NOR3X1_948/C NOR3X1_887/B NOR3X1_1277/B NOR3X1_930/A NOR3X1_930/B NOR3X1_930/C NOR3X1_929/A NOR3X1_929/B NOR3X1_779/C NOR3X1_1245/B NOR3X1_70/A NOR3X1_70/B NOR3X1_70/C NOR3X1_69/A NOR3X1_69/B NOR3X1_69/C 
+ NOR3X1_707/A NOR3X1_707/B NOR3X1_708/A NOR3X1_708/B NOR3X1_708/C NOR3X1_1543/B NOR3X1_999/B NOR3X1_1303/A NOR3X1_1303/B NOR3X1_1303/C NOR3X1_1304/A NOR3X1_1304/B NOR3X1_1304/C NOR3X1_381/B NOR3X1_1421/B NOR3X1_297/B NOR3X1_1293/B NOR3X1_1115/C NOR3X1_689/C NOR3X1_1099/C INVX1_1545/Y INVX1_1541/Y INVX1_1546/Y INVX1_1542/Y INVX1_1016/Y INVX1_1018/Y INVX1_1017/Y INVX1_1015/Y INVX1_1688/Y INVX1_1690/Y INVX1_1689/Y INVX1_1687/Y INVX1_784/Y INVX1_808/Y INVX1_807/Y INVX1_783/Y INVX1_911/Y INVX1_909/Y INVX1_912/Y INVX1_910/Y INVX1_67/Y INVX1_65/Y INVX1_68/Y INVX1_66/Y INVX1_880/Y INVX1_879/Y INVX1_1545/A INVX1_1541/A INVX1_1546/A INVX1_1542/A INVX1_1016/A 
+ INVX1_1018/A INVX1_1017/A INVX1_1015/A INVX1_1688/A INVX1_1690/A INVX1_1689/A INVX1_1687/A INVX1_784/A INVX1_783/A INVX1_911/A INVX1_912/A INVX1_67/A INVX1_65/A INVX1_68/A INVX1_66/A INVX1_880/A INVX1_879/A NOR3X1_1545/B NOR3X1_1541/B NOR3X1_1015/B NOR3X1_1687/B NOR3X1_808/A NOR3X1_808/B NOR3X1_808/C NOR3X1_807/A NOR3X1_807/B NOR3X1_807/C NOR3X1_783/C NOR3X1_911/B NOR3X1_909/A NOR3X1_909/B NOR3X1_909/C NOR3X1_910/A NOR3X1_910/B NOR3X1_910/C NOR3X1_879/B INVX1_805/Y INVX1_803/Y INVX1_806/Y INVX1_804/Y INVX1_890/Y INVX1_889/Y INVX1_805/A INVX1_803/A INVX1_806/A INVX1_804/A INVX1_890/A INVX1_889/A NOR3X1_805/B NOR3X1_803/B INVX1_231/Y 
+ INVX1_232/Y INVX1_1186/Y INVX1_1185/Y INVX1_1077/Y INVX1_1078/Y INVX1_508/Y INVX1_507/Y INVX1_637/Y INVX1_638/Y INVX1_1374/Y INVX1_1373/Y 
+ AES_SBOX_2

.include outputs_1.plw

* **************************************
* --- Simulation Settings ---
* **************************************

.param SIM_LEN = 50ns
.csparam SIM_LEN = {SIM_LEN}

*.options abstol=0.000001 vntol=0.001 reltol=0.01

.tran 1ns 'SIM_LEN'
.param SIMSTEP = 'SIM_LEN/1ns'
.csparam SIMSTEP = {SIMSTEP}

* **************************************
* --- Simulation Control ---
* **************************************

.control
    .include ../inputsD.inc

    run
    
    if ('writeFile' > 0)   
      wrdata ivdd_2.out i(vvdd)
      wrdata ivss_2.out i(vvss)
      *snsave sim_2.snap
    end
    
    set wr_vecnames
    set wr_singlescale
    wrdata outputs_2.out V("NOR3X1_1619/A") V("NOR3X1_1619/B") V("NOR3X1_1620/B") V("NOR3X1_951/A") V("NOR3X1_951/B") V("NOR3X1_952/B") V("NOR3X1_724/B") V("NOR3X1_723/A") V("NOR3X1_723/B") V("NOR3X1_1577/B") V("NOR3X1_952/A") V("NOR3X1_952/C") V("NOR3X1_724/A") V("NOR3X1_724/C") V("NOR3X1_1147/B") V("NOR3X1_1148/B") V("NOR3X1_1147/A") V("NOR3X1_1459/A") V("NOR3X1_1459/B") V("NOR3X1_1460/B") V("NOR3X1_1711/A") V("NOR3X1_1711/B") V("NOR3X1_1712/B") V("NOR3X1_1148/A") V("NOR3X1_1148/C") V("NOR3X1_678/A") V("NOR3X1_678/C") V("NOR3X1_677/B") V("NOR3X1_678/B") V("NOR3X1_677/A") V("NOR3X1_1429/C") V("NOR3X1_1430/A") V("NOR3X1_1430/B") V("NOR3X1_1430/C") V("NOR3X1_1429/A") V("NOR3X1_1460/A") V("NOR3X1_1460/C") V("NOR3X1_1712/A") V("NOR3X1_1712/C") V("NOR3X1_485/A") V("NOR3X1_485/B") V("NOR3X1_486/B") V("NOR3X1_486/A") V("NOR3X1_486/C") V("NOR3X1_675/B") V("NOR3X1_676/A") V("NOR3X1_676/C") V("NOR3X1_675/A") V("NOR3X1_676/B") V("NOR3X1_1620/C") V("NOR3X1_1620/A") V("NOR3X1_1264/B") V("NOR3X1_1263/A") V("NOR3X1_1263/B") V("NOR3X1_1264/A") V("NOR3X1_1264/C") V("NOR3X1_1275/B") V("NOR3X1_1113/C") V("NOR3X1_675/C") V("NOR3X1_1427/B") V("NOR3X1_1428/A") V("NOR3X1_1428/C") V("NOR3X1_907/C") V("NOR3X1_908/C") V("NOR3X1_907/A") V("NOR3X1_1428/B") V("NOR3X1_1427/A") V("NOR3X1_908/A") V("NOR3X1_908/B") V("NOR3X1_679/A") V("NOR3X1_679/B") V("NOR3X1_680/B") V("NOR3X1_680/A") V("NOR3X1_680/C") V("NOR3X1_1681/B") V("NOR3X1_1682/A") V("NOR3X1_1682/C") V("NOR3X1_1681/A") V("NOR3X1_1682/B") V("NOR3X1_1565/B") V("NOR3X1_1566/A") V("NOR3X1_1566/C") V("NOR3X1_1565/A") V("NOR3X1_1566/B") V("NOR3X1_1681/C") V("NOR3X1_1431/A") V("NOR3X1_1431/B") V("NOR3X1_1432/B") V("NOR3X1_1432/A") V("NOR3X1_1432/C") V("NOR3X1_1103/B") V("NOR3X1_1104/B") V("NOR3X1_1103/A") V("NOR3X1_1104/A") V("NOR3X1_1104/C") V("NOR3X1_1573/C") V("NOR3X1_1574/A") V("NOR3X1_1574/B") V("NOR3X1_1699/B") V("NOR3X1_1700/B") V("NOR3X1_1699/A") V("NOR3X1_1700/A") V("NOR3X1_1700/C") V("NOR3X1_1263/C") V("NOR3X1_315/C") V("NOR3X1_1586/C") V("NOR3X1_1585/A") V("NOR3X1_1585/C") V("NOR3X1_1586/B") V("NOR3X1_1586/A") V("NOR3X1_1679/B") V("NOR3X1_1680/A") V("NOR3X1_1680/C") V("NOR3X1_1565/C") V("NOR3X1_1679/A") V("NOR3X1_1680/B") V("NOR3X1_398/B") V("NOR3X1_397/A") V("NOR3X1_397/B") V("NOR3X1_398/C") V("NOR3X1_398/A") V("NOR3X1_1283/B") V("NOR3X1_1117/B") V("NOR3X1_1118/A") V("NOR3X1_1118/C") V("NOR3X1_1284/A") V("NOR3X1_1284/C") V("NOR3X1_1283/A") V("NOR3X1_1118/B") V("NOR3X1_1117/A") V("NOR3X1_1284/B") V("NOR3X1_1717/C") V("NOR3X1_1718/C") V("NOR3X1_1717/A") V("NOR3X1_1718/A") V("NOR3X1_1718/B") V("NOR3X1_277/B") V("NOR3X1_278/B") V("NOR3X1_277/A") V("NOR3X1_278/A") V("NOR3X1_278/C") V("NOR3X1_397/C") V("NOR3X1_907/B") V("NOR3X1_1134/C") V("NOR3X1_1133/A") V("NOR3X1_1133/C") V("NOR3X1_1134/A") V("NOR3X1_1134/B") V("NOR3X1_1704/C") V("NOR3X1_1703/A") V("NOR3X1_1703/C") V("NOR3X1_1704/A") V("NOR3X1_1704/B") V("NOR3X1_1425/B") V("NOR3X1_1426/A") V("NOR3X1_1426/C") V("NOR3X1_1287/A") V("NOR3X1_1287/B") V("NOR3X1_1288/B") V("NOR3X1_1467/A") V("NOR3X1_950/C") V("NOR3X1_1467/C") V("NOR3X1_1468/C") V("NOR3X1_949/A") V("NOR3X1_949/C") V("NOR3X1_1424/B") V("NOR3X1_1423/A") V("NOR3X1_1423/B") V("NOR3X1_1424/A") V("NOR3X1_1424/C") V("NOR3X1_1454/C") V("NOR3X1_1453/A") V("NOR3X1_1453/C") V("NOR3X1_705/A") V("NOR3X1_705/B") V("NOR3X1_706/B") V("NOR3X1_706/A") V("NOR3X1_706/C") V("NOR3X1_1454/A") V("NOR3X1_1454/B") V("NOR3X1_340/C") V("NOR3X1_339/A") V("NOR3X1_339/C") V("NOR3X1_340/A") V("NOR3X1_340/B") V("NOR3X1_1569/A") V("NOR3X1_1569/B") V("NOR3X1_1570/B") V("NOR3X1_1570/A") V("NOR3X1_1570/C") V("NOR3X1_1434/C") V("NOR3X1_1433/A") V("NOR3X1_1433/C") V("NOR3X1_1434/A") V("NOR3X1_1434/B") V("NOR3X1_674/A") V("NOR3X1_674/B") V("NOR3X1_673/C") V("NOR3X1_1573/A") V("NOR3X1_1574/C") V("NOR3X1_1301/A") V("NOR3X1_1301/C") V("NOR3X1_1302/C") V("NOR3X1_941/A") V("NOR3X1_941/C") V("NOR3X1_942/C") V("NOR3X1_942/A") V("NOR3X1_942/B") V("NOR3X1_1247/C") V("NOR3X1_1248/A") V("NOR3X1_1248/B") V("NOR3X1_1248/C") V("NOR3X1_1247/A") V("NOR3X1_1347/B") V("NOR3X1_1533/B") V("NOR3X1_157/B") V("NOR3X1_1229/B") V("NOR3X1_1033/B") V("NOR3X1_1333/B") V("NOR3X1_404/A") V("NOR3X1_404/B") V("NOR3X1_403/C") V("NOR3X1_415/A") V("NOR3X1_415/B") V("NOR3X1_416/B") V("NOR3X1_416/A") V("NOR3X1_416/C") V("NOR3X1_674/C") V("NOR3X1_673/A") V("NOR3X1_1583/C") V("NOR3X1_1584/A") V("NOR3X1_1584/B") V("NOR3X1_1513/B") V("NOR3X1_1568/B") V("NOR3X1_1567/A") V("NOR3X1_1567/B") V("NOR3X1_1568/A") V("NOR3X1_1568/C") V("NOR3X1_303/B") V("NOR3X1_373/B") V("NOR3X1_1187/B") V("NOR3X1_1359/B") V("NOR3X1_1105/B") V("NOR3X1_1106/A") V("NOR3X1_1106/C") V("NOR3X1_1509/B") V("NOR3X1_1329/B") V("NOR3X1_1217/B") V("NOR3X1_1331/B") V("NOR3X1_499/B") V("NOR3X1_1189/B") V("NOR3X1_995/B") V("NOR3X1_377/B") V("NOR3X1_1567/C") V("NOR3X1_1279/A") V("NOR3X1_1279/C") V("NOR3X1_1280/C") V("NOR3X1_1280/A") V("NOR3X1_1280/B") V("NOR3X1_919/C") V("NOR3X1_261/B") V("NOR3X1_987/B") V("NOR3X1_485/C") V("NOR3X1_1279/B") V("NOR3X1_905/C") V("NOR3X1_906/A") V("NOR3X1_906/B") V("NOR3X1_711/B") V("NOR3X1_712/A") V("NOR3X1_712/C") V("NOR3X1_711/A") V("NOR3X1_712/B") V("NOR3X1_905/A") V("NOR3X1_906/C") V("NOR3X1_1287/C") V("NOR3X1_1288/A") V("NOR3X1_1288/C") V("NOR3X1_1423/C") V("NOR3X1_615/B") V("NOR3X1_395/B") V("NOR3X1_1585/B") V("NOR3X1_1437/B") V("NOR3X1_1438/A") V("NOR3X1_1438/C") V("NOR3X1_407/C") V("NOR3X1_408/A") V("NOR3X1_408/B") V("NOR3X1_1555/B") V("NOR3X1_1093/B") V("NOR3X1_391/C") V("NOR3X1_1559/B") V("NOR3X1_361/B") V("NOR3X1_362/A") V("NOR3X1_362/C") V("NOR3X1_387/B") V("NOR3X1_388/A") V("NOR3X1_388/C") V("NOR3X1_1579/B") V("NOR3X1_1557/B") V("NOR3X1_1415/B") V("NOR3X1_479/C") V("NOR3X1_1283/C") V("NOR3X1_923/C") V("NOR3X1_419/C") V("NOR3X1_420/A") V("NOR3X1_420/B") V("NOR3X1_361/C") V("NOR3X1_362/B") V("NOR3X1_1302/A") V("NOR3X1_1302/B") V("NOR3X1_280/C") V("NOR3X1_279/B") V("NOR3X1_280/A") V("NOR3X1_385/B") V("NOR3X1_386/A") V("NOR3X1_386/C") V("NOR3X1_521/B") V("NOR3X1_679/C") V("NOR3X1_1553/B") V("NOR3X1_1437/C") V("NOR3X1_1438/B") V("NOR3X1_387/C") V("NOR3X1_388/B") V("NOR3X1_385/C") V("NOR3X1_386/B") V("NOR3X1_1117/C") V("NOR3X1_603/C") V("NOR3X1_1085/C") V("NOR3X1_1269/C") V("NOR3X1_901/C") V("NOR3X1_453/C") V("NOR3X1_1087/B") V("NOR3X1_1088/A") V("NOR3X1_1088/C") V("NOR3X1_1265/C") V("NOR3X1_1349/A") V("NOR3X1_1349/B") V("NOR3X1_1350/B") V("NOR3X1_349/C") V("NOR3X1_350/A") V("NOR3X1_350/B") V("NOR3X1_1350/C") V("NOR3X1_1350/A") V("NOR3X1_360/C") V("NOR3X1_359/B") V("NOR3X1_360/A") V("NOR3X1_1407/C") V("NOR3X1_405/C") V("NOR3X1_406/A") V("NOR3X1_406/B") V("NOR3X1_899/B") V("NOR3X1_1001/C") V("NOR3X1_1002/A") V("NOR3X1_1002/B") V("NOR3X1_1001/A") V("NOR3X1_1002/C") V("NOR3X1_401/B") V("NOR3X1_402/A") V("NOR3X1_402/C") V("NOR3X1_1709/B") V("NOR3X1_1435/C") V("NOR3X1_1436/A") V("NOR3X1_1436/B") V("NOR3X1_1663/C") V("NOR3X1_1417/C") V("NOR3X1_293/C") V("NOR3X1_1039/C") V("NOR3X1_1468/A") V("NOR3X1_1468/B") V("NOR3X1_950/A") V("NOR3X1_950/B") V("NOR3X1_1575/C") V("NOR3X1_1576/A") V("NOR3X1_1576/B") V("NOR3X1_1069/C") V("NOR3X1_1305/C") V("NOR3X1_1306/A") V("NOR3X1_1306/B") V("NOR3X1_893/B") V("NOR3X1_384/A") V("NOR3X1_384/B") V("NOR3X1_383/C") V("NOR3X1_1671/C") V("NOR3X1_1551/B") V("NOR3X1_335/B") V("NOR3X1_933/C") V("NOR3X1_420/C") V("NOR3X1_419/B") V("NOR3X1_934/A") V("NOR3X1_934/B") V("NOR3X1_891/B") V("NOR3X1_1011/C") V("NOR3X1_484/A") V("NOR3X1_484/B") V("NOR3X1_483/C") V("NOR3X1_1685/C") V("NOR3X1_1090/C") V("NOR3X1_1089/B") V("NOR3X1_1090/A") V("NOR3X1_1451/C") V("NOR3X1_1452/A") V("NOR3X1_1452/B") V("NOR3X1_417/B") V("NOR3X1_418/A") V("NOR3X1_418/C") V("NOR3X1_683/B") V("NOR3X1_1564/A") V("NOR3X1_1564/B") V("NOR3X1_1563/C") V("NOR3X1_1107/C") V("NOR3X1_1108/A") V("NOR3X1_1108/B") V("NOR3X1_1413/B") V("NOR3X1_1345/C") V("NOR3X1_1537/B") V("NOR3X1_1572/A") V("NOR3X1_1572/C") V("NOR3X1_1571/B") V("NOR3X1_1089/C") V("NOR3X1_1090/B") V("NOR3X1_665/C") V("NOR3X1_1097/C") V("NOR3X1_781/B") V("NOR3X1_389/C") V("NOR3X1_1223/C") V("NOR3X1_1281/B") V("NOR3X1_1282/A") V("NOR3X1_1282/C") V("NOR3X1_1517/B") V("NOR3X1_601/C") V("NOR3X1_275/C") V("NOR3X1_663/B") V("NOR3X1_1337/B") V("NOR3X1_1267/C") V("NOR3X1_667/C") V("NOR3X1_1285/B") V("NOR3X1_1286/A") V("NOR3X1_1286/C") V("NOR3X1_359/C") V("NOR3X1_360/B") V("NOR3X1_133/B") V("NOR3X1_777/C") V("NOR3X1_1667/B") V("NOR3X1_1355/B") V("NOR3X1_1087/C") V("NOR3X1_1088/B") V("NOR3X1_359/A") V("NOR3X1_1089/A") V("NOR3X1_1564/C") V("NOR3X1_1563/A") V("NOR3X1_387/A") V("NOR3X1_1583/A") V("NOR3X1_1584/C") V("NOR3X1_404/C") V("NOR3X1_403/A") V("NOR3X1_361/A") V("NOR3X1_484/C") V("NOR3X1_483/A") V("NOR3X1_1087/A") V("NOR3X1_431/A") V("NOR3X1_1311/A") V("NOR3X1_431/C") V("NOR3X1_1311/C") V("NOR3X1_432/C") V("NOR3X1_1312/C") V("NOR3X1_432/A") V("NOR3X1_432/B") V("NOR3X1_1312/A") V("NOR3X1_1312/B") V("NOR3X1_1121/A") V("NOR3X1_1121/C") V("NOR3X1_1122/C") V("NOR3X1_696/C") V("NOR3X1_695/A") V("NOR3X1_695/C") V("NOR3X1_1122/A") V("NOR3X1_1122/B") V("NOR3X1_385/A") V("NOR3X1_696/A") V("NOR3X1_696/B") V("NOR3X1_697/A") V("NOR3X1_697/C") V("NOR3X1_698/C") V("NOR3X1_698/A") V("NOR3X1_698/B") V("NOR3X1_247/C") V("NOR3X1_248/A") V("NOR3X1_248/B") V("NOR3X1_248/C") V("NOR3X1_247/A") V("NOR3X1_1110/C") V("NOR3X1_1109/B") V("NOR3X1_1110/A") V("NOR3X1_1109/A") V("NOR3X1_1110/B") V("NOR3X1_1105/A") V("NOR3X1_1106/B") V("NOR3X1_693/C") V("NOR3X1_694/A") V("NOR3X1_694/B") V("NOR3X1_693/A") V("NOR3X1_694/C") V("NOR3X1_403/B") V("NOR3X1_405/A") V("NOR3X1_406/C") V("NOR3X1_350/C") V("NOR3X1_349/A") V("NOR3X1_401/A") V("NOR3X1_402/B") V("NOR3X1_1572/B") V("NOR3X1_1571/A") V("NOR3X1_1425/A") V("NOR3X1_1426/B") V("NOR3X1_1130/C") V("NOR3X1_1129/A") V("NOR3X1_1129/C") V("NOR3X1_1130/A") V("NOR3X1_1130/B") V("NOR3X1_933/A") V("NOR3X1_419/A") V("NOR3X1_934/C") V("NOR3X1_1451/A") V("NOR3X1_1452/C") V("NOR3X1_418/B") V("NOR3X1_417/A") V("NOR3X1_1107/A") V("NOR3X1_1108/C") V("NOR3X1_1435/A") V("NOR3X1_1436/C") V("NOR3X1_1285/A") V("NOR3X1_1286/B") V("NOR3X1_1282/B") V("NOR3X1_1281/A") V("NOR3X1_1437/A") V("NOR3X1_408/C") V("NOR3X1_407/A") V("NOR3X1_279/A") V("NOR3X1_280/B") V("NOR3X1_1305/A") V("NOR3X1_1306/C") V("NOR3X1_1576/C") V("NOR3X1_1575/A") V("NOR3X1_384/C") V("NOR3X1_383/A") V("INVX1_965/Y") V("INVX1_966/Y") V("INVX1_534/Y") V("INVX1_533/Y") V("INVX1_323/A") V("INVX1_324/A") V("INVX1_1673/A") V("INVX1_1674/A") V("INVX1_965/A") V("INVX1_966/A") V("INVX1_1257/A") V("INVX1_1258/A") V("INVX1_567/A") V("INVX1_568/A") V("INVX1_508/A") V("INVX1_507/A") V("INVX1_197/A") V("INVX1_198/A") V("INVX1_662/A") V("INVX1_661/A") V("INVX1_1241/A") V("INVX1_1242/A") V("INVX1_913/A") V("INVX1_914/A") V("INVX1_569/A") V("INVX1_570/A") V("INVX1_1691/A") V("INVX1_1692/A") V("INVX1_534/A") V("INVX1_533/A") V("NOR3X1_197/C") V("NOR3X1_232/A") V("NOR3X1_232/B") V("NOR3X1_232/C") V("NOR3X1_231/A") V("NOR3X1_231/B") V("NOR3X1_231/C") V("INVX1_194/Y") V("INVX1_193/Y") V("INVX1_229/Y") V("INVX1_227/Y") V("INVX1_230/Y") V("INVX1_228/Y") V("INVX1_194/A") V("INVX1_193/A") V("INVX1_229/A") V("INVX1_227/A") V("INVX1_230/A") V("INVX1_228/A") V("NOR3X1_1596/A") V("NOR3X1_1596/B") V("NOR3X1_1596/C") V("NOR3X1_1598/A") V("NOR3X1_1598/B") V("NOR3X1_1598/C") V("NOR3X1_1597/A") V("NOR3X1_1597/B") V("NOR3X1_1595/A") V("NOR3X1_1595/B") V("NOR3X1_227/B") V("INVX1_871/Y") V("INVX1_872/Y") V("INVX1_226/Y") V("INVX1_225/Y") V("INVX1_871/A") V("INVX1_872/A") V("INVX1_1185/A") V("INVX1_1186/A") V("INVX1_226/A") V("INVX1_225/A") V("NOR3X1_871/C") V("NOR3X1_637/A") V("NOR3X1_637/B") V("NOR3X1_637/C") V("NOR3X1_638/A") V("NOR3X1_638/B") V("NOR3X1_638/C") V("NOR3X1_1185/B") V("NOR3X1_1077/A") V("NOR3X1_1077/B") V("NOR3X1_1077/C") V("NOR3X1_1078/A") V("NOR3X1_1078/B") V("NOR3X1_1078/C") V("INVX1_868/Y") V("INVX1_867/Y") V("INVX1_634/Y") V("INVX1_636/Y") V("INVX1_635/Y") V("INVX1_633/Y") V("INVX1_1184/Y") V("INVX1_1183/Y") V("INVX1_1074/Y") V("INVX1_1076/Y") V("INVX1_1075/Y") V("INVX1_1073/Y") V("INVX1_868/A") V("INVX1_867/A") V("INVX1_634/A") V("INVX1_636/A") V("INVX1_635/A") V("INVX1_633/A") V("INVX1_1184/A") V("INVX1_1183/A") V("INVX1_1074/A") V("INVX1_1076/A") V("INVX1_1075/A") V("INVX1_1073/A") V("INVX1_1548/Y") V("INVX1_1547/Y") V("INVX1_944/Y") V("INVX1_943/Y") V("INVX1_575/Y") V("INVX1_576/Y") V("INVX1_1019/Y") V("INVX1_1020/Y") V("INVX1_1456/Y") V("INVX1_1455/Y") V("INVX1_1708/Y") V("INVX1_1707/Y") V("INVX1_121/Y") V("INVX1_122/Y") V("INVX1_1403/Y") V("INVX1_1404/Y") V("INVX1_1092/Y") V("INVX1_1091/Y") V("INVX1_647/Y") V("INVX1_648/Y") V("INVX1_1669/Y") V("INVX1_1670/Y") V("INVX1_1535/Y") V("INVX1_1536/Y") V("INVX1_1405/Y") V("INVX1_1406/Y") V("INVX1_456/Y") V("INVX1_455/Y") V("INVX1_1083/Y") V("INVX1_1084/Y") V("INVX1_971/Y") V("INVX1_972/Y") V("INVX1_1683/Y") V("INVX1_1684/Y") V("INVX1_1665/Y") V("INVX1_1666/Y") V("INVX1_1697/Y") V("INVX1_1698/Y") V("INVX1_273/Y") V("INVX1_274/Y") V("INVX1_1014/Y") V("INVX1_1013/Y") V("INVX1_651/Y") V("INVX1_652/Y") V("INVX1_1677/Y") V("INVX1_1678/Y") V("INVX1_1540/Y") V("INVX1_1539/Y") V("INVX1_1409/Y") V("INVX1_1410/Y") V("INVX1_1442/Y") V("INVX1_947/Y") V("INVX1_1441/Y") V("INVX1_948/Y") V("INVX1_295/Y") V("INVX1_296/Y") V("INVX1_887/Y") V("INVX1_888/Y") V("INVX1_606/Y") V("INVX1_605/Y") V("INVX1_337/Y") V("INVX1_338/Y") V("INVX1_1550/Y") V("INVX1_1549/Y") V("INVX1_985/Y") V("INVX1_986/Y") V("INVX1_671/Y") V("INVX1_672/Y") V("INVX1_1278/Y") V("INVX1_1277/Y") V("INVX1_930/Y") V("INVX1_929/Y") V("INVX1_1440/Y") V("INVX1_1439/Y") V("INVX1_779/Y") V("INVX1_780/Y") V("INVX1_1245/Y") V("INVX1_1246/Y") V("INVX1_517/Y") V("INVX1_518/Y") V("INVX1_1291/Y") V("INVX1_1292/Y") V("INVX1_70/Y") V("INVX1_69/Y") V("INVX1_1581/Y") V("INVX1_1582/Y") V("INVX1_1079/Y") V("INVX1_1080/Y") V("INVX1_897/Y") V("INVX1_898/Y") V("INVX1_707/Y") V("INVX1_708/Y") V("INVX1_776/Y") V("INVX1_775/Y") V("INVX1_1271/Y") V("INVX1_1272/Y") V("INVX1_167/Y") V("INVX1_168/Y") V("INVX1_1046/Y") V("INVX1_997/Y") V("INVX1_998/Y") V("INVX1_1045/Y") V("INVX1_1239/Y") V("INVX1_1240/Y") V("INVX1_256/Y") V("INVX1_255/Y") V("INVX1_1543/Y") V("INVX1_1544/Y") V("INVX1_801/Y") V("INVX1_802/Y") V("INVX1_878/Y") V("INVX1_877/Y") V("INVX1_347/Y") V("INVX1_348/Y") V("INVX1_151/Y") V("INVX1_152/Y") V("INVX1_999/Y") V("INVX1_1000/Y") V("INVX1_1209/Y") V("INVX1_1210/Y") V("INVX1_1203/Y") V("INVX1_1204/Y") V("INVX1_1303/Y") V("INVX1_1304/Y") V("INVX1_1659/Y") V("INVX1_1660/Y") V("INVX1_381/Y") V("INVX1_382/Y") V("INVX1_1358/Y") V("INVX1_1357/Y") V("INVX1_903/Y") V("INVX1_904/Y") V("INVX1_481/Y") V("INVX1_482/Y") V("INVX1_1421/Y") V("INVX1_1422/Y") V("INVX1_297/Y") V("INVX1_298/Y") V("INVX1_1561/Y") V("INVX1_1562/Y") V("INVX1_885/Y") V("INVX1_886/Y") V("INVX1_379/Y") V("INVX1_380/Y") V("INVX1_461/Y") V("INVX1_462/Y") V("INVX1_1294/Y") V("INVX1_1293/Y") V("INVX1_1116/Y") V("INVX1_1115/Y") V("INVX1_689/Y") V("INVX1_690/Y") V("INVX1_925/Y") V("INVX1_926/Y") V("INVX1_686/Y") V("INVX1_685/Y") V("INVX1_245/Y") V("INVX1_246/Y") V("INVX1_799/Y") V("INVX1_800/Y") V("INVX1_691/Y") V("INVX1_692/Y") V("INVX1_1420/Y") V("INVX1_1419/Y") V("INVX1_1099/Y") V("INVX1_1100/Y") V("INVX1_944/A") V("INVX1_943/A") V("INVX1_575/A") V("INVX1_576/A") V("INVX1_1456/A") V("INVX1_1455/A") V("INVX1_1708/A") V("INVX1_1707/A") V("INVX1_121/A") V("INVX1_122/A") V("INVX1_1403/A") V("INVX1_1404/A") V("INVX1_1092/A") V("INVX1_1091/A") V("INVX1_647/A") V("INVX1_648/A") V("INVX1_1669/A") V("INVX1_1670/A") V("INVX1_1535/A") V("INVX1_1536/A") V("INVX1_1405/A") V("INVX1_1406/A") V("INVX1_456/A") V("INVX1_455/A") V("INVX1_1083/A") V("INVX1_1084/A") V("INVX1_971/A") V("INVX1_972/A") V("INVX1_1683/A") V("INVX1_1684/A") V("INVX1_1665/A") V("INVX1_1666/A") V("INVX1_273/A") V("INVX1_274/A") V("INVX1_1014/A") V("INVX1_1013/A") V("INVX1_651/A") V("INVX1_652/A") V("INVX1_1677/A") V("INVX1_1678/A") V("INVX1_1540/A") V("INVX1_1539/A") V("INVX1_1409/A") V("INVX1_1410/A") V("INVX1_1442/A") V("INVX1_1441/A") V("INVX1_295/A") V("INVX1_296/A") V("INVX1_887/A") V("INVX1_888/A") V("INVX1_606/A") V("INVX1_605/A") V("INVX1_337/A") V("INVX1_338/A") V("INVX1_1550/A") V("INVX1_1549/A") V("INVX1_985/A") V("INVX1_986/A") V("INVX1_671/A") V("INVX1_672/A") V("INVX1_1278/A") V("INVX1_1277/A") V("INVX1_1440/A") V("INVX1_1439/A") V("INVX1_779/A") V("INVX1_780/A") V("INVX1_1245/A") V("INVX1_1246/A") V("INVX1_517/A") V("INVX1_518/A") V("INVX1_1291/A") V("INVX1_1292/A") V("INVX1_1581/A") V("INVX1_1582/A") V("INVX1_1079/A") V("INVX1_1080/A") V("INVX1_897/A") V("INVX1_898/A") V("INVX1_776/A") V("INVX1_775/A") V("INVX1_1271/A") V("INVX1_1272/A") V("INVX1_167/A") V("INVX1_168/A") V("INVX1_1046/A") V("INVX1_997/A") V("INVX1_998/A") V("INVX1_1045/A") V("INVX1_1239/A") V("INVX1_1240/A") V("INVX1_256/A") V("INVX1_255/A") V("INVX1_1543/A") V("INVX1_1544/A") V("INVX1_801/A") V("INVX1_802/A") V("INVX1_878/A") V("INVX1_877/A") V("INVX1_347/A") V("INVX1_348/A") V("INVX1_151/A") V("INVX1_152/A") V("INVX1_999/A") V("INVX1_1000/A") V("INVX1_1209/A") V("INVX1_1210/A") V("INVX1_1203/A") V("INVX1_1204/A") V("INVX1_1659/A") V("INVX1_1660/A") V("INVX1_381/A") V("INVX1_382/A") V("INVX1_1358/A") V("INVX1_1357/A") V("INVX1_903/A") V("INVX1_904/A") V("INVX1_481/A") V("INVX1_482/A") V("INVX1_1421/A") V("INVX1_1422/A") V("INVX1_297/A") V("INVX1_298/A") V("INVX1_1561/A") V("INVX1_1562/A") V("INVX1_885/A") V("INVX1_886/A") V("INVX1_379/A") V("INVX1_380/A") V("INVX1_461/A") V("INVX1_462/A") V("INVX1_1294/A") V("INVX1_1293/A") V("INVX1_1116/A") V("INVX1_1115/A") V("INVX1_689/A") V("INVX1_690/A") V("INVX1_925/A") V("INVX1_926/A") V("INVX1_686/A") V("INVX1_685/A") V("INVX1_245/A") V("INVX1_246/A") V("INVX1_799/A") V("INVX1_800/A") V("INVX1_691/A") V("INVX1_692/A") V("INVX1_1420/A") V("INVX1_1419/A") V("INVX1_1099/A") V("INVX1_1100/A") V("NOR3X1_1548/A") V("NOR3X1_1548/B") V("NOR3X1_1548/C") V("NOR3X1_1547/A") V("NOR3X1_1547/B") V("NOR3X1_1547/C") V("NOR3X1_943/B") V("NOR3X1_1019/A") V("NOR3X1_1019/B") V("NOR3X1_1019/C") V("NOR3X1_1020/A") V("NOR3X1_1020/B") V("NOR3X1_1020/C") V("NOR3X1_1455/C") V("NOR3X1_1707/C") V("NOR3X1_1683/B") V("NOR3X1_1697/A") V("NOR3X1_1697/B") V("NOR3X1_1697/C") V("NOR3X1_1698/A") V("NOR3X1_1698/B") V("NOR3X1_1698/C") V("NOR3X1_651/C") V("NOR3X1_1677/C") V("NOR3X1_947/A") V("NOR3X1_947/C") V("NOR3X1_1441/B") V("NOR3X1_948/A") V("NOR3X1_948/B") V("NOR3X1_948/C") V("NOR3X1_887/B") V("NOR3X1_1277/B") V("NOR3X1_930/A") V("NOR3X1_930/B") V("NOR3X1_930/C") V("NOR3X1_929/A") V("NOR3X1_929/B") V("NOR3X1_779/C") V("NOR3X1_1245/B") V("NOR3X1_70/A") V("NOR3X1_70/B") V("NOR3X1_70/C") V("NOR3X1_69/A") V("NOR3X1_69/B") V("NOR3X1_69/C") V("NOR3X1_707/A") V("NOR3X1_707/B") V("NOR3X1_708/A") V("NOR3X1_708/B") V("NOR3X1_708/C") V("NOR3X1_1543/B") V("NOR3X1_999/B") V("NOR3X1_1303/A") V("NOR3X1_1303/B") V("NOR3X1_1303/C") V("NOR3X1_1304/A") V("NOR3X1_1304/B") V("NOR3X1_1304/C") V("NOR3X1_381/B") V("NOR3X1_1421/B") V("NOR3X1_297/B") V("NOR3X1_1293/B") V("NOR3X1_1115/C") V("NOR3X1_689/C") V("NOR3X1_1099/C") V("INVX1_1545/Y") V("INVX1_1541/Y") V("INVX1_1546/Y") V("INVX1_1542/Y") V("INVX1_1016/Y") V("INVX1_1018/Y") V("INVX1_1017/Y") V("INVX1_1015/Y") V("INVX1_1688/Y") V("INVX1_1690/Y") V("INVX1_1689/Y") V("INVX1_1687/Y") V("INVX1_784/Y") V("INVX1_808/Y") V("INVX1_807/Y") V("INVX1_783/Y") V("INVX1_911/Y") V("INVX1_909/Y") V("INVX1_912/Y") V("INVX1_910/Y") V("INVX1_67/Y") V("INVX1_65/Y") V("INVX1_68/Y") V("INVX1_66/Y") V("INVX1_880/Y") V("INVX1_879/Y") V("INVX1_1545/A") V("INVX1_1541/A") V("INVX1_1546/A") V("INVX1_1542/A") V("INVX1_1016/A") V("INVX1_1018/A") V("INVX1_1017/A") V("INVX1_1015/A") V("INVX1_1688/A") V("INVX1_1690/A") V("INVX1_1689/A") V("INVX1_1687/A") V("INVX1_784/A") V("INVX1_783/A") V("INVX1_911/A") V("INVX1_912/A") V("INVX1_67/A") V("INVX1_65/A") V("INVX1_68/A") V("INVX1_66/A") V("INVX1_880/A") V("INVX1_879/A") V("NOR3X1_1545/B") V("NOR3X1_1541/B") V("NOR3X1_1015/B") V("NOR3X1_1687/B") V("NOR3X1_808/A") V("NOR3X1_808/B") V("NOR3X1_808/C") V("NOR3X1_807/A") V("NOR3X1_807/B") V("NOR3X1_807/C") V("NOR3X1_783/C") V("NOR3X1_911/B") V("NOR3X1_909/A") V("NOR3X1_909/B") V("NOR3X1_909/C") V("NOR3X1_910/A") V("NOR3X1_910/B") V("NOR3X1_910/C") V("NOR3X1_879/B") V("INVX1_805/Y") V("INVX1_803/Y") V("INVX1_806/Y") V("INVX1_804/Y") V("INVX1_890/Y") V("INVX1_889/Y") V("INVX1_805/A") V("INVX1_803/A") V("INVX1_806/A") V("INVX1_804/A") V("INVX1_890/A") V("INVX1_889/A") V("NOR3X1_805/B") V("NOR3X1_803/B") V("INVX1_231/Y") V("INVX1_232/Y") V("INVX1_1186/Y") V("INVX1_1185/Y") V("INVX1_1077/Y") V("INVX1_1078/Y") V("INVX1_508/Y") V("INVX1_507/Y") V("INVX1_637/Y") V("INVX1_638/Y") V("INVX1_1374/Y") V("INVX1_1373/Y") 
    
    if ('showPlots' < 1)
       quit
    end
       
.endc

.end
