* SPICE3 file created from dualRail.ext - technology: scmos
*
* drain/source ordering enforced by hand
*

.subckt AND2X1_LOC a_36_24# Y a_8_24# VSS VDD A B
X0 Y a_8_24# VDD VDD PMOS_MAGIC ad=1p pd=5u as=2.2p ps=10.2u w=2u l=0.2u
X1 a_8_24# A a_36_24# VSS NMOS_MAGIC ad=0.6p pd=4.6u as=1p ps=5u w=2u l=0.2u
X2 Y a_8_24# VSS VSS NMOS_MAGIC ad=0.5p pd=3u as=1.1p ps=5.2u w=1u l=0.2u
X3 a_36_24# B VSS VSS NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=2u l=0.2u
X4 a_8_24# B VDD VDD PMOS_MAGIC ad=0p pd=0u as=1.2p ps=5.2u w=2u l=0.2u
X5 a_8_24# A VDD VDD PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=2u l=0.2u

C0 B a_8_24# 0.33fF
C1 a_8_24# Y 0.46fF
C2 a_8_24# a_36_24# 0.00fF
C3 VDD A 0.20fF
C4 VDD B 0.25fF
C5 A B 0.26fF
C6 VDD a_8_24# 0.82fF
C7 VDD Y 0.38fF
C8 A a_8_24# 0.06fF
C9 Y VSS 0.13fF
C10 a_8_24# VSS 0.48fF
C11 B VSS 0.19fF
C12 A VSS 0.25fF
C13 VDD VSS 2.08fF
.ends

.subckt OR2X1_LOC a_8_216# a_36_216# Y VSS VDD A B
X0 a_36_216# B VDD VDD PMOS_MAGIC ad=2.2p pd=9.2u as=1.2p ps=8.6u w=4u l=0.2u
X1 Y a_8_216# VDD VDD PMOS_MAGIC ad=1p pd=5u as=0p ps=0u w=2u l=0.2u
X2 a_8_216# B VSS VSS NMOS_MAGIC ad=1.1p pd=6.2u as=0.6p ps=3.2u w=1u l=0.2u
X3 a_8_216# A VSS VSS NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=1u l=0.2u
X4 a_8_216# A a_36_216# VDD PMOS_MAGIC ad=0p pd=0u as=2p ps=9u w=4u l=0.2u
X5 Y a_8_216# VSS VSS NMOS_MAGIC ad=0.5p pd=3u as=0p ps=0u w=1u l=0.2u

C0 VDD Y 0.41fF
C1 B a_8_216# 0.30fF
C2 a_8_216# Y 0.37fF
C3 VDD A 0.07fF
C4 VDD B 0.07fF
C5 A B 0.22fF
C6 VDD a_8_216# 0.45fF
C7 A a_8_216# 0.06fF
C8 Y VSS 0.29fF
C9 a_8_216# VSS 0.68fF
C10 B VSS 0.31fF
C11 A VSS 0.37fF
C12 VDD VSS 2.08fF
.ends

.subckt AES_SBOX INPUT_0 INPUT_1 INPUT_2 INPUT_3 INPUT_4 INPUT_5 INPUT_6 INPUT_7 
+ D_INPUT_0 D_INPUT_1 D_INPUT_2 D_INPUT_3 D_INPUT_4 D_INPUT_5 D_INPUT_6 D_INPUT_7 
+ GATE_222 GATE_366 GATE_479 GATE_579 GATE_662 GATE_741 GATE_811 GATE_865 
+ D_GATE_222 D_GATE_366 D_GATE_479 D_GATE_579 D_GATE_662 D_GATE_741 D_GATE_811 D_GATE_865 
+ VDD VSS 

XAND2X1_LOC_229 AND2X1_LOC_229/a_36_24# OR2X1_LOC_231/B AND2X1_LOC_229/a_8_24# VSS VDD
+ AND2X1_LOC_12/Y OR2X1_LOC_160/B AND2X1_LOC
XAND2X1_LOC_218 AND2X1_LOC_218/a_36_24# AND2X1_LOC_218/Y AND2X1_LOC_218/a_8_24# VSS VDD
+ AND2X1_LOC_216/Y AND2X1_LOC_217/Y AND2X1_LOC
XAND2X1_LOC_207 AND2X1_LOC_207/a_36_24# AND2X1_LOC_214/A AND2X1_LOC_207/a_8_24# VSS VDD
+ AND2X1_LOC_207/A AND2X1_LOC_207/B AND2X1_LOC
XAND2X1_LOC_741 AND2X1_LOC_741/a_36_24# AND2X1_LOC_741/Y AND2X1_LOC_741/a_8_24# VSS VDD
+ AND2X1_LOC_736/Y AND2X1_LOC_737/Y AND2X1_LOC
XAND2X1_LOC_730 AND2X1_LOC_730/a_36_24# AND2X1_LOC_739/B AND2X1_LOC_730/a_8_24# VSS VDD
+ AND2X1_LOC_728/Y AND2X1_LOC_729/Y AND2X1_LOC
XOR2X1_LOC_549 OR2X1_LOC_549/a_8_216# OR2X1_LOC_549/a_36_216# OR2X1_LOC_549/Y VSS VDD
+ OR2X1_LOC_549/A OR2X1_LOC_549/B OR2X1_LOC
XOR2X1_LOC_505 OR2X1_LOC_505/a_8_216# OR2X1_LOC_505/a_36_216# OR2X1_LOC_505/Y VSS VDD
+ OR2X1_LOC_45/B OR2X1_LOC_18/Y OR2X1_LOC
XOR2X1_LOC_527 OR2X1_LOC_527/a_8_216# OR2X1_LOC_527/a_36_216# OR2X1_LOC_527/Y VSS VDD
+ OR2X1_LOC_323/A OR2X1_LOC_64/Y OR2X1_LOC
XOR2X1_LOC_538 OR2X1_LOC_538/a_8_216# OR2X1_LOC_538/a_36_216# OR2X1_LOC_539/A VSS VDD
+ OR2X1_LOC_538/A OR2X1_LOC_193/A OR2X1_LOC
XOR2X1_LOC_516 OR2X1_LOC_516/a_8_216# OR2X1_LOC_516/a_36_216# OR2X1_LOC_516/Y VSS VDD
+ OR2X1_LOC_516/A OR2X1_LOC_516/B OR2X1_LOC
XAND2X1_LOC_785 AND2X1_LOC_785/a_36_24# AND2X1_LOC_785/Y AND2X1_LOC_785/a_8_24# VSS VDD
+ AND2X1_LOC_785/A AND2X1_LOC_776/Y AND2X1_LOC
XAND2X1_LOC_774 AND2X1_LOC_774/a_36_24# AND2X1_LOC_810/A AND2X1_LOC_774/a_8_24# VSS VDD
+ AND2X1_LOC_774/A AND2X1_LOC_773/Y AND2X1_LOC
XAND2X1_LOC_796 AND2X1_LOC_796/a_36_24# AND2X1_LOC_796/Y AND2X1_LOC_796/a_8_24# VSS VDD
+ AND2X1_LOC_796/A AND2X1_LOC_784/Y AND2X1_LOC
XAND2X1_LOC_763 AND2X1_LOC_763/a_36_24# OR2X1_LOC_769/B AND2X1_LOC_763/a_8_24# VSS VDD
+ AND2X1_LOC_48/A AND2X1_LOC_763/B AND2X1_LOC
XAND2X1_LOC_752 AND2X1_LOC_752/a_36_24# AND2X1_LOC_753/B AND2X1_LOC_752/a_8_24# VSS VDD
+ INPUT_5 AND2X1_LOC_50/Y AND2X1_LOC
XOR2X1_LOC_313 OR2X1_LOC_313/a_8_216# OR2X1_LOC_313/a_36_216# OR2X1_LOC_313/Y VSS VDD
+ OR2X1_LOC_91/A OR2X1_LOC_70/Y OR2X1_LOC
XAND2X1_LOC_560 AND2X1_LOC_560/a_36_24# AND2X1_LOC_571/A AND2X1_LOC_560/a_8_24# VSS VDD
+ AND2X1_LOC_523/Y AND2X1_LOC_560/B AND2X1_LOC
XAND2X1_LOC_571 AND2X1_LOC_571/a_36_24# AND2X1_LOC_571/Y AND2X1_LOC_571/a_8_24# VSS VDD
+ AND2X1_LOC_571/A AND2X1_LOC_571/B AND2X1_LOC
XAND2X1_LOC_593 AND2X1_LOC_593/a_36_24# AND2X1_LOC_593/Y AND2X1_LOC_593/a_8_24# VSS VDD
+ OR2X1_LOC_591/Y AND2X1_LOC_592/Y AND2X1_LOC
XAND2X1_LOC_582 AND2X1_LOC_582/a_36_24# OR2X1_LOC_635/A AND2X1_LOC_582/a_8_24# VSS VDD
+ OR2X1_LOC_161/B AND2X1_LOC_582/B AND2X1_LOC
XOR2X1_LOC_346 OR2X1_LOC_346/a_8_216# OR2X1_LOC_346/a_36_216# OR2X1_LOC_347/A VSS VDD
+ OR2X1_LOC_346/A OR2X1_LOC_346/B OR2X1_LOC
XOR2X1_LOC_335 OR2X1_LOC_335/a_8_216# OR2X1_LOC_335/a_36_216# OR2X1_LOC_335/Y VSS VDD
+ OR2X1_LOC_335/A OR2X1_LOC_335/B OR2X1_LOC
XOR2X1_LOC_357 OR2X1_LOC_357/a_8_216# OR2X1_LOC_357/a_36_216# OR2X1_LOC_364/B VSS VDD
+ OR2X1_LOC_357/A OR2X1_LOC_357/B OR2X1_LOC
XOR2X1_LOC_368 OR2X1_LOC_368/a_8_216# OR2X1_LOC_368/a_36_216# OR2X1_LOC_368/Y VSS VDD
+ OR2X1_LOC_368/A OR2X1_LOC_7/A OR2X1_LOC
XOR2X1_LOC_302 OR2X1_LOC_302/a_8_216# OR2X1_LOC_302/a_36_216# OR2X1_LOC_303/A VSS VDD
+ OR2X1_LOC_302/A OR2X1_LOC_302/B OR2X1_LOC
XOR2X1_LOC_324 OR2X1_LOC_324/a_8_216# OR2X1_LOC_324/a_36_216# OR2X1_LOC_326/B VSS VDD
+ OR2X1_LOC_324/A OR2X1_LOC_324/B OR2X1_LOC
XOR2X1_LOC_379 OR2X1_LOC_379/a_8_216# OR2X1_LOC_379/a_36_216# OR2X1_LOC_379/Y VSS VDD
+ OR2X1_LOC_66/A AND2X1_LOC_12/Y OR2X1_LOC
XOR2X1_LOC_110 OR2X1_LOC_110/a_8_216# OR2X1_LOC_110/a_36_216# OR2X1_LOC_323/A VSS VDD
+ OR2X1_LOC_46/A INPUT_0 OR2X1_LOC
XOR2X1_LOC_154 OR2X1_LOC_154/a_8_216# OR2X1_LOC_154/a_36_216# OR2X1_LOC_156/B VSS VDD
+ OR2X1_LOC_154/A AND2X1_LOC_7/B OR2X1_LOC
XAND2X1_LOC_390 AND2X1_LOC_390/a_36_24# AND2X1_LOC_392/A AND2X1_LOC_390/a_8_24# VSS VDD
+ AND2X1_LOC_388/Y AND2X1_LOC_390/B AND2X1_LOC
XOR2X1_LOC_187 OR2X1_LOC_187/a_8_216# OR2X1_LOC_187/a_36_216# OR2X1_LOC_187/Y VSS VDD
+ OR2X1_LOC_680/A OR2X1_LOC_40/Y OR2X1_LOC
XOR2X1_LOC_143 OR2X1_LOC_143/a_8_216# OR2X1_LOC_143/a_36_216# OR2X1_LOC_696/A VSS VDD
+ OR2X1_LOC_8/Y INPUT_1 OR2X1_LOC
XOR2X1_LOC_121 OR2X1_LOC_121/a_8_216# OR2X1_LOC_121/a_36_216# OR2X1_LOC_121/Y VSS VDD
+ OR2X1_LOC_121/A OR2X1_LOC_121/B OR2X1_LOC
XOR2X1_LOC_132 OR2X1_LOC_132/a_8_216# OR2X1_LOC_132/a_36_216# OR2X1_LOC_132/Y VSS VDD
+ OR2X1_LOC_95/Y OR2X1_LOC_91/A OR2X1_LOC
XOR2X1_LOC_165 OR2X1_LOC_165/a_8_216# OR2X1_LOC_165/a_36_216# OR2X1_LOC_165/Y VSS VDD
+ OR2X1_LOC_74/A OR2X1_LOC_51/Y OR2X1_LOC
XOR2X1_LOC_198 OR2X1_LOC_198/a_8_216# OR2X1_LOC_198/a_36_216# OR2X1_LOC_208/A VSS VDD
+ OR2X1_LOC_198/A AND2X1_LOC_57/Y OR2X1_LOC
XOR2X1_LOC_176 OR2X1_LOC_176/a_8_216# OR2X1_LOC_176/a_36_216# OR2X1_LOC_176/Y VSS VDD
+ OR2X1_LOC_91/A OR2X1_LOC_26/Y OR2X1_LOC
XOR2X1_LOC_709 OR2X1_LOC_709/a_8_216# OR2X1_LOC_709/a_36_216# OR2X1_LOC_711/B VSS VDD
+ OR2X1_LOC_709/A OR2X1_LOC_709/B OR2X1_LOC
XAND2X1_LOC_219 AND2X1_LOC_219/a_36_24# AND2X1_LOC_219/Y AND2X1_LOC_219/a_8_24# VSS VDD
+ AND2X1_LOC_219/A AND2X1_LOC_215/Y AND2X1_LOC
XAND2X1_LOC_208 AND2X1_LOC_208/a_36_24# AND2X1_LOC_208/Y AND2X1_LOC_208/a_8_24# VSS VDD
+ AND2X1_LOC_35/Y AND2X1_LOC_208/B AND2X1_LOC
XAND2X1_LOC_720 AND2X1_LOC_720/a_36_24# AND2X1_LOC_720/Y AND2X1_LOC_720/a_8_24# VSS VDD
+ OR2X1_LOC_667/Y OR2X1_LOC_669/Y AND2X1_LOC
XAND2X1_LOC_775 AND2X1_LOC_775/a_36_24# AND2X1_LOC_785/A AND2X1_LOC_775/a_8_24# VSS VDD
+ OR2X1_LOC_91/Y OR2X1_LOC_109/Y AND2X1_LOC
XAND2X1_LOC_731 AND2X1_LOC_731/a_36_24# AND2X1_LOC_731/Y AND2X1_LOC_731/a_8_24# VSS VDD
+ AND2X1_LOC_726/Y AND2X1_LOC_727/Y AND2X1_LOC
XAND2X1_LOC_742 AND2X1_LOC_742/a_36_24# GATE_741 AND2X1_LOC_742/a_8_24# VSS VDD
+ AND2X1_LOC_742/A AND2X1_LOC_741/Y AND2X1_LOC
XAND2X1_LOC_764 AND2X1_LOC_764/a_36_24# OR2X1_LOC_769/A AND2X1_LOC_764/a_8_24# VSS VDD
+ AND2X1_LOC_40/Y OR2X1_LOC_160/A AND2X1_LOC
XAND2X1_LOC_753 AND2X1_LOC_753/a_36_24# OR2X1_LOC_790/B AND2X1_LOC_753/a_8_24# VSS VDD
+ OR2X1_LOC_185/Y AND2X1_LOC_753/B AND2X1_LOC
XOR2X1_LOC_506 OR2X1_LOC_506/a_8_216# OR2X1_LOC_506/a_36_216# OR2X1_LOC_506/Y VSS VDD
+ OR2X1_LOC_506/A OR2X1_LOC_506/B OR2X1_LOC
XOR2X1_LOC_528 OR2X1_LOC_528/a_8_216# OR2X1_LOC_528/a_36_216# OR2X1_LOC_528/Y VSS VDD
+ OR2X1_LOC_44/Y OR2X1_LOC_7/A OR2X1_LOC
XOR2X1_LOC_517 OR2X1_LOC_517/a_8_216# OR2X1_LOC_517/a_36_216# OR2X1_LOC_517/Y VSS VDD
+ OR2X1_LOC_517/A OR2X1_LOC_31/Y OR2X1_LOC
XOR2X1_LOC_539 OR2X1_LOC_539/a_8_216# OR2X1_LOC_539/a_36_216# OR2X1_LOC_539/Y VSS VDD
+ OR2X1_LOC_539/A OR2X1_LOC_539/B OR2X1_LOC
XAND2X1_LOC_786 AND2X1_LOC_786/a_36_24# AND2X1_LOC_786/Y AND2X1_LOC_786/a_8_24# VSS VDD
+ AND2X1_LOC_84/Y OR2X1_LOC_262/Y AND2X1_LOC
XAND2X1_LOC_797 AND2X1_LOC_797/a_36_24# AND2X1_LOC_803/B AND2X1_LOC_797/a_8_24# VSS VDD
+ AND2X1_LOC_797/A AND2X1_LOC_797/B AND2X1_LOC
XOR2X1_LOC_314 OR2X1_LOC_314/a_8_216# OR2X1_LOC_314/a_36_216# OR2X1_LOC_314/Y VSS VDD
+ OR2X1_LOC_64/Y OR2X1_LOC_16/A OR2X1_LOC
XAND2X1_LOC_561 AND2X1_LOC_561/a_36_24# AND2X1_LOC_571/B AND2X1_LOC_561/a_8_24# VSS VDD
+ AND2X1_LOC_557/Y AND2X1_LOC_561/B AND2X1_LOC
XAND2X1_LOC_572 AND2X1_LOC_572/a_36_24# AND2X1_LOC_572/Y AND2X1_LOC_572/a_8_24# VSS VDD
+ AND2X1_LOC_572/A AND2X1_LOC_361/A AND2X1_LOC
XAND2X1_LOC_594 AND2X1_LOC_594/a_36_24# OR2X1_LOC_653/B AND2X1_LOC_594/a_8_24# VSS VDD
+ AND2X1_LOC_95/Y OR2X1_LOC_186/Y AND2X1_LOC
XAND2X1_LOC_550 AND2X1_LOC_550/a_36_24# AND2X1_LOC_565/B AND2X1_LOC_550/a_8_24# VSS VDD
+ AND2X1_LOC_550/A AND2X1_LOC_547/Y AND2X1_LOC
XAND2X1_LOC_583 AND2X1_LOC_583/a_36_24# OR2X1_LOC_636/B AND2X1_LOC_583/a_8_24# VSS VDD
+ AND2X1_LOC_31/Y OR2X1_LOC_87/A AND2X1_LOC
XOR2X1_LOC_347 OR2X1_LOC_347/a_8_216# OR2X1_LOC_347/a_36_216# OR2X1_LOC_347/Y VSS VDD
+ OR2X1_LOC_347/A OR2X1_LOC_347/B OR2X1_LOC
XOR2X1_LOC_358 OR2X1_LOC_358/a_8_216# OR2X1_LOC_358/a_36_216# OR2X1_LOC_364/A VSS VDD
+ OR2X1_LOC_358/A OR2X1_LOC_358/B OR2X1_LOC
XOR2X1_LOC_303 OR2X1_LOC_303/a_8_216# OR2X1_LOC_303/a_36_216# OR2X1_LOC_566/A VSS VDD
+ OR2X1_LOC_303/A OR2X1_LOC_303/B OR2X1_LOC
XOR2X1_LOC_336 OR2X1_LOC_336/a_8_216# OR2X1_LOC_336/a_36_216# OR2X1_LOC_337/A VSS VDD
+ OR2X1_LOC_703/A OR2X1_LOC_538/A OR2X1_LOC
XOR2X1_LOC_369 OR2X1_LOC_369/a_8_216# OR2X1_LOC_369/a_36_216# OR2X1_LOC_369/Y VSS VDD
+ OR2X1_LOC_426/B OR2X1_LOC_22/Y OR2X1_LOC
XOR2X1_LOC_325 OR2X1_LOC_325/a_8_216# OR2X1_LOC_325/a_36_216# OR2X1_LOC_325/Y VSS VDD
+ OR2X1_LOC_325/A OR2X1_LOC_325/B OR2X1_LOC
XOR2X1_LOC_144 OR2X1_LOC_144/a_8_216# OR2X1_LOC_144/a_36_216# OR2X1_LOC_144/Y VSS VDD
+ OR2X1_LOC_696/A OR2X1_LOC_59/Y OR2X1_LOC
XOR2X1_LOC_133 OR2X1_LOC_133/a_8_216# OR2X1_LOC_133/a_36_216# OR2X1_LOC_427/A VSS VDD
+ OR2X1_LOC_49/A OR2X1_LOC_8/Y OR2X1_LOC
XOR2X1_LOC_122 OR2X1_LOC_122/a_8_216# OR2X1_LOC_122/a_36_216# OR2X1_LOC_122/Y VSS VDD
+ OR2X1_LOC_122/A OR2X1_LOC_44/Y OR2X1_LOC
XOR2X1_LOC_100 OR2X1_LOC_100/a_8_216# OR2X1_LOC_100/a_36_216# OR2X1_LOC_100/Y VSS VDD
+ AND2X1_LOC_88/Y AND2X1_LOC_86/Y OR2X1_LOC
XOR2X1_LOC_111 OR2X1_LOC_111/a_8_216# OR2X1_LOC_111/a_36_216# OR2X1_LOC_111/Y VSS VDD
+ OR2X1_LOC_323/A OR2X1_LOC_31/Y OR2X1_LOC
XOR2X1_LOC_199 OR2X1_LOC_199/a_8_216# OR2X1_LOC_199/a_36_216# OR2X1_LOC_207/B VSS VDD
+ OR2X1_LOC_196/Y OR2X1_LOC_199/B OR2X1_LOC
XOR2X1_LOC_155 OR2X1_LOC_155/a_8_216# OR2X1_LOC_155/a_36_216# OR2X1_LOC_156/A VSS VDD
+ OR2X1_LOC_155/A OR2X1_LOC_87/A OR2X1_LOC
XOR2X1_LOC_166 OR2X1_LOC_166/a_8_216# OR2X1_LOC_166/a_36_216# OR2X1_LOC_166/Y VSS VDD
+ OR2X1_LOC_40/Y OR2X1_LOC_16/A OR2X1_LOC
XAND2X1_LOC_391 AND2X1_LOC_391/a_36_24# AND2X1_LOC_391/Y AND2X1_LOC_391/a_8_24# VSS VDD
+ OR2X1_LOC_382/Y OR2X1_LOC_384/Y AND2X1_LOC
XAND2X1_LOC_380 AND2X1_LOC_380/a_36_24# OR2X1_LOC_460/B AND2X1_LOC_380/a_8_24# VSS VDD
+ OR2X1_LOC_160/A OR2X1_LOC_379/Y AND2X1_LOC
XOR2X1_LOC_188 OR2X1_LOC_188/a_8_216# OR2X1_LOC_188/a_36_216# OR2X1_LOC_188/Y VSS VDD
+ OR2X1_LOC_185/Y OR2X1_LOC_154/A OR2X1_LOC
XOR2X1_LOC_177 OR2X1_LOC_177/a_8_216# OR2X1_LOC_177/a_36_216# OR2X1_LOC_177/Y VSS VDD
+ OR2X1_LOC_70/Y OR2X1_LOC_52/B OR2X1_LOC
XAND2X1_LOC_209 AND2X1_LOC_209/a_36_24# AND2X1_LOC_209/Y AND2X1_LOC_209/a_8_24# VSS VDD
+ AND2X1_LOC_797/A OR2X1_LOC_152/Y AND2X1_LOC
XAND2X1_LOC_721 AND2X1_LOC_721/a_36_24# AND2X1_LOC_721/Y AND2X1_LOC_721/a_8_24# VSS VDD
+ AND2X1_LOC_721/A AND2X1_LOC_720/Y AND2X1_LOC
XAND2X1_LOC_710 AND2X1_LOC_710/a_36_24# AND2X1_LOC_710/Y AND2X1_LOC_710/a_8_24# VSS VDD
+ OR2X1_LOC_700/Y OR2X1_LOC_701/Y AND2X1_LOC
XAND2X1_LOC_765 AND2X1_LOC_765/a_36_24# OR2X1_LOC_770/B AND2X1_LOC_765/a_8_24# VSS VDD
+ AND2X1_LOC_12/Y OR2X1_LOC_78/B AND2X1_LOC
XAND2X1_LOC_776 AND2X1_LOC_776/a_36_24# AND2X1_LOC_776/Y AND2X1_LOC_776/a_8_24# VSS VDD
+ OR2X1_LOC_164/Y OR2X1_LOC_238/Y AND2X1_LOC
XAND2X1_LOC_787 AND2X1_LOC_787/a_36_24# AND2X1_LOC_794/A AND2X1_LOC_787/a_8_24# VSS VDD
+ AND2X1_LOC_787/A AND2X1_LOC_486/Y AND2X1_LOC
XAND2X1_LOC_798 AND2X1_LOC_798/a_36_24# AND2X1_LOC_798/Y AND2X1_LOC_798/a_8_24# VSS VDD
+ AND2X1_LOC_798/A AND2X1_LOC_436/Y AND2X1_LOC
XAND2X1_LOC_743 AND2X1_LOC_743/a_36_24# OR2X1_LOC_780/B AND2X1_LOC_743/a_8_24# VSS VDD
+ AND2X1_LOC_3/Y OR2X1_LOC_155/A AND2X1_LOC
XAND2X1_LOC_754 AND2X1_LOC_754/a_36_24# OR2X1_LOC_790/A AND2X1_LOC_754/a_8_24# VSS VDD
+ AND2X1_LOC_36/Y OR2X1_LOC_614/Y AND2X1_LOC
XAND2X1_LOC_732 AND2X1_LOC_732/a_36_24# AND2X1_LOC_738/B AND2X1_LOC_732/a_8_24# VSS VDD
+ AND2X1_LOC_724/Y AND2X1_LOC_732/B AND2X1_LOC
XOR2X1_LOC_507 OR2X1_LOC_507/a_8_216# OR2X1_LOC_507/a_36_216# OR2X1_LOC_508/A VSS VDD
+ OR2X1_LOC_507/A OR2X1_LOC_507/B OR2X1_LOC
XOR2X1_LOC_529 OR2X1_LOC_529/a_8_216# OR2X1_LOC_529/a_36_216# OR2X1_LOC_529/Y VSS VDD
+ OR2X1_LOC_26/Y D_INPUT_3 OR2X1_LOC
XOR2X1_LOC_518 OR2X1_LOC_518/a_8_216# OR2X1_LOC_518/a_36_216# OR2X1_LOC_518/Y VSS VDD
+ OR2X1_LOC_74/A OR2X1_LOC_64/Y OR2X1_LOC
XOR2X1_LOC_304 OR2X1_LOC_304/a_8_216# OR2X1_LOC_304/a_36_216# OR2X1_LOC_304/Y VSS VDD
+ OR2X1_LOC_428/A OR2X1_LOC_53/Y OR2X1_LOC
XOR2X1_LOC_315 OR2X1_LOC_315/a_8_216# OR2X1_LOC_315/a_36_216# OR2X1_LOC_315/Y VSS VDD
+ OR2X1_LOC_427/A OR2X1_LOC_31/Y OR2X1_LOC
XOR2X1_LOC_326 OR2X1_LOC_326/a_8_216# OR2X1_LOC_326/a_36_216# OR2X1_LOC_354/A VSS VDD
+ OR2X1_LOC_325/Y OR2X1_LOC_326/B OR2X1_LOC
XAND2X1_LOC_573 AND2X1_LOC_573/a_36_24# AND2X1_LOC_573/Y AND2X1_LOC_573/a_8_24# VSS VDD
+ AND2X1_LOC_573/A AND2X1_LOC_501/Y AND2X1_LOC
XAND2X1_LOC_562 AND2X1_LOC_562/a_36_24# AND2X1_LOC_562/Y AND2X1_LOC_562/a_8_24# VSS VDD
+ AND2X1_LOC_555/Y AND2X1_LOC_562/B AND2X1_LOC
XAND2X1_LOC_595 AND2X1_LOC_595/a_36_24# OR2X1_LOC_643/A AND2X1_LOC_595/a_8_24# VSS VDD
+ OR2X1_LOC_66/A OR2X1_LOC_249/Y AND2X1_LOC
XAND2X1_LOC_540 AND2X1_LOC_540/a_36_24# AND2X1_LOC_553/A AND2X1_LOC_540/a_8_24# VSS VDD
+ OR2X1_LOC_178/Y OR2X1_LOC_183/Y AND2X1_LOC
XAND2X1_LOC_584 AND2X1_LOC_584/a_36_24# OR2X1_LOC_636/A AND2X1_LOC_584/a_8_24# VSS VDD
+ AND2X1_LOC_7/B AND2X1_LOC_51/Y AND2X1_LOC
XAND2X1_LOC_551 AND2X1_LOC_551/a_36_24# AND2X1_LOC_564/A AND2X1_LOC_551/a_8_24# VSS VDD
+ AND2X1_LOC_544/Y AND2X1_LOC_551/B AND2X1_LOC
XOR2X1_LOC_348 OR2X1_LOC_348/a_8_216# OR2X1_LOC_348/a_36_216# OR2X1_LOC_348/Y VSS VDD
+ OR2X1_LOC_345/Y OR2X1_LOC_348/B OR2X1_LOC
XOR2X1_LOC_359 OR2X1_LOC_359/a_8_216# OR2X1_LOC_359/a_36_216# OR2X1_LOC_363/B VSS VDD
+ OR2X1_LOC_359/A OR2X1_LOC_348/Y OR2X1_LOC
XOR2X1_LOC_337 OR2X1_LOC_337/a_8_216# OR2X1_LOC_337/a_36_216# OR2X1_LOC_352/A VSS VDD
+ OR2X1_LOC_337/A OR2X1_LOC_335/Y OR2X1_LOC
XOR2X1_LOC_860 OR2X1_LOC_860/a_8_216# OR2X1_LOC_860/a_36_216# OR2X1_LOC_860/Y VSS VDD
+ OR2X1_LOC_474/B OR2X1_LOC_244/Y OR2X1_LOC
XOR2X1_LOC_145 OR2X1_LOC_145/a_8_216# OR2X1_LOC_145/a_36_216# OR2X1_LOC_145/Y VSS VDD
+ OR2X1_LOC_89/A OR2X1_LOC_51/Y OR2X1_LOC
XOR2X1_LOC_156 OR2X1_LOC_156/a_8_216# OR2X1_LOC_156/a_36_216# OR2X1_LOC_156/Y VSS VDD
+ OR2X1_LOC_156/A OR2X1_LOC_156/B OR2X1_LOC
XOR2X1_LOC_167 OR2X1_LOC_167/a_8_216# OR2X1_LOC_167/a_36_216# OR2X1_LOC_167/Y VSS VDD
+ OR2X1_LOC_604/A OR2X1_LOC_64/Y OR2X1_LOC
XOR2X1_LOC_123 OR2X1_LOC_123/a_8_216# OR2X1_LOC_123/a_36_216# OR2X1_LOC_124/A VSS VDD
+ OR2X1_LOC_633/B OR2X1_LOC_123/B OR2X1_LOC
XOR2X1_LOC_101 OR2X1_LOC_101/a_8_216# OR2X1_LOC_101/a_36_216# OR2X1_LOC_656/B VSS VDD
+ OR2X1_LOC_100/Y OR2X1_LOC_99/Y OR2X1_LOC
XOR2X1_LOC_134 OR2X1_LOC_134/a_8_216# OR2X1_LOC_134/a_36_216# OR2X1_LOC_134/Y VSS VDD
+ OR2X1_LOC_427/A OR2X1_LOC_95/Y OR2X1_LOC
XOR2X1_LOC_112 OR2X1_LOC_112/a_8_216# OR2X1_LOC_112/a_36_216# OR2X1_LOC_715/B VSS VDD
+ OR2X1_LOC_112/A OR2X1_LOC_112/B OR2X1_LOC
XAND2X1_LOC_392 AND2X1_LOC_392/a_36_24# AND2X1_LOC_474/A AND2X1_LOC_392/a_8_24# VSS VDD
+ AND2X1_LOC_392/A AND2X1_LOC_391/Y AND2X1_LOC
XAND2X1_LOC_381 AND2X1_LOC_381/a_36_24# AND2X1_LOC_817/B AND2X1_LOC_381/a_8_24# VSS VDD
+ INPUT_3 AND2X1_LOC_12/Y AND2X1_LOC
XAND2X1_LOC_370 AND2X1_LOC_370/a_36_24# AND2X1_LOC_787/A AND2X1_LOC_370/a_8_24# VSS VDD
+ OR2X1_LOC_309/Y OR2X1_LOC_369/Y AND2X1_LOC
XOR2X1_LOC_178 OR2X1_LOC_178/a_8_216# OR2X1_LOC_178/a_36_216# OR2X1_LOC_178/Y VSS VDD
+ OR2X1_LOC_158/A OR2X1_LOC_56/A OR2X1_LOC
XOR2X1_LOC_189 OR2X1_LOC_189/a_8_216# OR2X1_LOC_189/a_36_216# OR2X1_LOC_189/Y VSS VDD
+ OR2X1_LOC_189/A OR2X1_LOC_95/Y OR2X1_LOC
XOR2X1_LOC_690 OR2X1_LOC_690/a_8_216# OR2X1_LOC_690/a_36_216# OR2X1_LOC_690/Y VSS VDD
+ OR2X1_LOC_690/A INPUT_0 OR2X1_LOC
XOR2X1_LOC_508 OR2X1_LOC_508/a_8_216# OR2X1_LOC_508/a_36_216# OR2X1_LOC_508/Y VSS VDD
+ OR2X1_LOC_508/A OR2X1_LOC_506/Y OR2X1_LOC
XAND2X1_LOC_711 AND2X1_LOC_711/a_36_24# AND2X1_LOC_711/Y AND2X1_LOC_711/a_8_24# VSS VDD
+ AND2X1_LOC_711/A AND2X1_LOC_710/Y AND2X1_LOC
XAND2X1_LOC_755 AND2X1_LOC_755/a_36_24# OR2X1_LOC_791/B AND2X1_LOC_755/a_8_24# VSS VDD
+ AND2X1_LOC_59/Y OR2X1_LOC_664/Y AND2X1_LOC
XAND2X1_LOC_766 AND2X1_LOC_766/a_36_24# OR2X1_LOC_770/A AND2X1_LOC_766/a_8_24# VSS VDD
+ AND2X1_LOC_64/Y AND2X1_LOC_91/B AND2X1_LOC
XAND2X1_LOC_722 AND2X1_LOC_722/a_36_24# AND2X1_LOC_722/Y AND2X1_LOC_722/a_8_24# VSS VDD
+ AND2X1_LOC_722/A AND2X1_LOC_719/Y AND2X1_LOC
XAND2X1_LOC_733 AND2X1_LOC_733/a_36_24# AND2X1_LOC_733/Y AND2X1_LOC_733/a_8_24# VSS VDD
+ AND2X1_LOC_722/Y AND2X1_LOC_723/Y AND2X1_LOC
XAND2X1_LOC_777 AND2X1_LOC_777/a_36_24# AND2X1_LOC_784/A AND2X1_LOC_777/a_8_24# VSS VDD
+ OR2X1_LOC_246/A OR2X1_LOC_305/Y AND2X1_LOC
XAND2X1_LOC_799 AND2X1_LOC_799/a_36_24# AND2X1_LOC_802/B AND2X1_LOC_799/a_8_24# VSS VDD
+ AND2X1_LOC_539/Y AND2X1_LOC_593/Y AND2X1_LOC
XAND2X1_LOC_788 AND2X1_LOC_788/a_36_24# AND2X1_LOC_794/B AND2X1_LOC_788/a_8_24# VSS VDD
+ OR2X1_LOC_533/Y AND2X1_LOC_645/A AND2X1_LOC
XAND2X1_LOC_700 AND2X1_LOC_700/a_36_24# OR2X1_LOC_710/B AND2X1_LOC_700/a_8_24# VSS VDD
+ AND2X1_LOC_59/Y AND2X1_LOC_91/B AND2X1_LOC
XAND2X1_LOC_744 AND2X1_LOC_744/a_36_24# OR2X1_LOC_780/A AND2X1_LOC_744/a_8_24# VSS VDD
+ AND2X1_LOC_44/Y OR2X1_LOC_160/A AND2X1_LOC
XOR2X1_LOC_519 OR2X1_LOC_519/a_8_216# OR2X1_LOC_519/a_36_216# OR2X1_LOC_519/Y VSS VDD
+ OR2X1_LOC_158/A OR2X1_LOC_48/B OR2X1_LOC
XOR2X1_LOC_305 OR2X1_LOC_305/a_8_216# OR2X1_LOC_305/a_36_216# OR2X1_LOC_305/Y VSS VDD
+ OR2X1_LOC_91/A OR2X1_LOC_3/Y OR2X1_LOC
XAND2X1_LOC_541 AND2X1_LOC_541/a_36_24# AND2X1_LOC_541/Y AND2X1_LOC_541/a_8_24# VSS VDD
+ OR2X1_LOC_256/A OR2X1_LOC_272/Y AND2X1_LOC
XAND2X1_LOC_530 AND2X1_LOC_530/a_36_24# OR2X1_LOC_548/A AND2X1_LOC_530/a_8_24# VSS VDD
+ AND2X1_LOC_36/Y OR2X1_LOC_532/B AND2X1_LOC
XOR2X1_LOC_349 OR2X1_LOC_349/a_8_216# OR2X1_LOC_349/a_36_216# OR2X1_LOC_359/A VSS VDD
+ OR2X1_LOC_349/A OR2X1_LOC_349/B OR2X1_LOC
XOR2X1_LOC_327 OR2X1_LOC_327/a_8_216# OR2X1_LOC_327/a_36_216# OR2X1_LOC_405/A VSS VDD
+ OR2X1_LOC_264/Y AND2X1_LOC_65/A OR2X1_LOC
XOR2X1_LOC_316 OR2X1_LOC_316/a_8_216# OR2X1_LOC_316/a_36_216# OR2X1_LOC_316/Y VSS VDD
+ OR2X1_LOC_80/Y OR2X1_LOC_12/Y OR2X1_LOC
XOR2X1_LOC_338 OR2X1_LOC_338/a_8_216# OR2X1_LOC_338/a_36_216# OR2X1_LOC_351/B VSS VDD
+ OR2X1_LOC_338/A OR2X1_LOC_338/B OR2X1_LOC
XAND2X1_LOC_574 AND2X1_LOC_574/a_36_24# AND2X1_LOC_574/Y AND2X1_LOC_574/a_8_24# VSS VDD
+ AND2X1_LOC_574/A OR2X1_LOC_516/Y AND2X1_LOC
XAND2X1_LOC_563 AND2X1_LOC_563/a_36_24# AND2X1_LOC_563/Y AND2X1_LOC_563/a_8_24# VSS VDD
+ AND2X1_LOC_563/A AND2X1_LOC_554/Y AND2X1_LOC
XAND2X1_LOC_552 AND2X1_LOC_552/a_36_24# AND2X1_LOC_564/B AND2X1_LOC_552/a_8_24# VSS VDD
+ AND2X1_LOC_552/A AND2X1_LOC_543/Y AND2X1_LOC
XAND2X1_LOC_585 AND2X1_LOC_585/a_36_24# OR2X1_LOC_637/B AND2X1_LOC_585/a_8_24# VSS VDD
+ AND2X1_LOC_22/Y OR2X1_LOC_598/A AND2X1_LOC
XAND2X1_LOC_596 AND2X1_LOC_596/a_36_24# OR2X1_LOC_597/A AND2X1_LOC_596/a_8_24# VSS VDD
+ OR2X1_LOC_44/Y OR2X1_LOC_421/A AND2X1_LOC
XOR2X1_LOC_850 OR2X1_LOC_850/a_8_216# OR2X1_LOC_850/a_36_216# OR2X1_LOC_858/B VSS VDD
+ OR2X1_LOC_850/A OR2X1_LOC_850/B OR2X1_LOC
XOR2X1_LOC_861 OR2X1_LOC_861/a_8_216# OR2X1_LOC_861/a_36_216# OR2X1_LOC_865/B VSS VDD
+ OR2X1_LOC_860/Y OR2X1_LOC_624/Y OR2X1_LOC
XOR2X1_LOC_157 OR2X1_LOC_157/a_8_216# OR2X1_LOC_157/a_36_216# OR2X1_LOC_158/A VSS VDD
+ OR2X1_LOC_17/Y OR2X1_LOC_2/Y OR2X1_LOC
XOR2X1_LOC_146 OR2X1_LOC_146/a_8_216# OR2X1_LOC_146/a_36_216# OR2X1_LOC_146/Y VSS VDD
+ OR2X1_LOC_744/A OR2X1_LOC_36/Y OR2X1_LOC
XOR2X1_LOC_135 OR2X1_LOC_135/a_8_216# OR2X1_LOC_135/a_36_216# OR2X1_LOC_135/Y VSS VDD
+ OR2X1_LOC_427/A OR2X1_LOC_59/Y OR2X1_LOC
XAND2X1_LOC_371 AND2X1_LOC_371/a_36_24# OR2X1_LOC_778/B AND2X1_LOC_371/a_8_24# VSS VDD
+ OR2X1_LOC_68/B AND2X1_LOC_31/Y AND2X1_LOC
XAND2X1_LOC_360 AND2X1_LOC_360/a_36_24# AND2X1_LOC_363/B AND2X1_LOC_360/a_8_24# VSS VDD
+ AND2X1_LOC_860/A AND2X1_LOC_347/Y AND2X1_LOC
XAND2X1_LOC_382 AND2X1_LOC_382/a_36_24# OR2X1_LOC_391/B AND2X1_LOC_382/a_8_24# VSS VDD
+ OR2X1_LOC_80/A AND2X1_LOC_817/B AND2X1_LOC
XOR2X1_LOC_113 OR2X1_LOC_113/a_8_216# OR2X1_LOC_113/a_36_216# OR2X1_LOC_113/Y VSS VDD
+ OR2X1_LOC_113/A OR2X1_LOC_113/B OR2X1_LOC
XOR2X1_LOC_102 OR2X1_LOC_102/a_8_216# OR2X1_LOC_102/a_36_216# OR2X1_LOC_485/A VSS VDD
+ OR2X1_LOC_54/Y OR2X1_LOC_8/Y OR2X1_LOC
XOR2X1_LOC_124 OR2X1_LOC_124/a_8_216# OR2X1_LOC_124/a_36_216# OR2X1_LOC_124/Y VSS VDD
+ OR2X1_LOC_124/A OR2X1_LOC_124/B OR2X1_LOC
XOR2X1_LOC_179 OR2X1_LOC_179/a_8_216# OR2X1_LOC_179/a_36_216# OR2X1_LOC_179/Y VSS VDD
+ OR2X1_LOC_600/A OR2X1_LOC_36/Y OR2X1_LOC
XOR2X1_LOC_168 OR2X1_LOC_168/a_8_216# OR2X1_LOC_168/a_36_216# OR2X1_LOC_168/Y VSS VDD
+ OR2X1_LOC_168/A OR2X1_LOC_168/B OR2X1_LOC
XAND2X1_LOC_393 AND2X1_LOC_393/a_36_24# OR2X1_LOC_400/B AND2X1_LOC_393/a_8_24# VSS VDD
+ OR2X1_LOC_154/A AND2X1_LOC_40/Y AND2X1_LOC
XOR2X1_LOC_680 OR2X1_LOC_680/a_8_216# OR2X1_LOC_680/a_36_216# OR2X1_LOC_680/Y VSS VDD
+ OR2X1_LOC_680/A OR2X1_LOC_51/Y OR2X1_LOC
XOR2X1_LOC_691 OR2X1_LOC_691/a_8_216# OR2X1_LOC_691/a_36_216# OR2X1_LOC_691/Y VSS VDD
+ OR2X1_LOC_691/A OR2X1_LOC_691/B OR2X1_LOC
XAND2X1_LOC_190 AND2X1_LOC_190/a_36_24# AND2X1_LOC_191/B AND2X1_LOC_190/a_8_24# VSS VDD
+ OR2X1_LOC_183/Y OR2X1_LOC_184/Y AND2X1_LOC
XAND2X1_LOC_723 AND2X1_LOC_723/a_36_24# AND2X1_LOC_723/Y AND2X1_LOC_723/a_8_24# VSS VDD
+ AND2X1_LOC_716/Y AND2X1_LOC_717/Y AND2X1_LOC
XAND2X1_LOC_701 AND2X1_LOC_701/a_36_24# OR2X1_LOC_710/A AND2X1_LOC_701/a_8_24# VSS VDD
+ AND2X1_LOC_44/Y OR2X1_LOC_269/B AND2X1_LOC
XAND2X1_LOC_712 AND2X1_LOC_712/a_36_24# AND2X1_LOC_712/Y AND2X1_LOC_712/a_8_24# VSS VDD
+ AND2X1_LOC_707/Y AND2X1_LOC_712/B AND2X1_LOC
XOR2X1_LOC_509 OR2X1_LOC_509/a_8_216# OR2X1_LOC_509/a_36_216# OR2X1_LOC_510/A VSS VDD
+ OR2X1_LOC_509/A OR2X1_LOC_227/Y OR2X1_LOC
XAND2X1_LOC_756 AND2X1_LOC_756/a_36_24# OR2X1_LOC_757/A AND2X1_LOC_756/a_8_24# VSS VDD
+ OR2X1_LOC_600/A OR2X1_LOC_604/A AND2X1_LOC
XAND2X1_LOC_789 AND2X1_LOC_789/a_36_24# AND2X1_LOC_789/Y AND2X1_LOC_789/a_8_24# VSS VDD
+ OR2X1_LOC_748/Y OR2X1_LOC_751/Y AND2X1_LOC
XAND2X1_LOC_767 AND2X1_LOC_767/a_36_24# OR2X1_LOC_773/B AND2X1_LOC_767/a_8_24# VSS VDD
+ AND2X1_LOC_3/Y OR2X1_LOC_78/Y AND2X1_LOC
XAND2X1_LOC_778 AND2X1_LOC_778/a_36_24# AND2X1_LOC_778/Y AND2X1_LOC_778/a_8_24# VSS VDD
+ OR2X1_LOC_371/Y OR2X1_LOC_496/Y AND2X1_LOC
XAND2X1_LOC_734 AND2X1_LOC_734/a_36_24# AND2X1_LOC_734/Y AND2X1_LOC_734/a_8_24# VSS VDD
+ OR2X1_LOC_406/Y AND2X1_LOC_721/Y AND2X1_LOC
XAND2X1_LOC_745 AND2X1_LOC_745/a_36_24# OR2X1_LOC_781/B AND2X1_LOC_745/a_8_24# VSS VDD
+ AND2X1_LOC_40/Y OR2X1_LOC_161/A AND2X1_LOC
XOR2X1_LOC_328 OR2X1_LOC_328/a_8_216# OR2X1_LOC_328/a_36_216# OR2X1_LOC_421/A VSS VDD
+ OR2X1_LOC_70/A INPUT_4 OR2X1_LOC
XOR2X1_LOC_306 OR2X1_LOC_306/a_8_216# OR2X1_LOC_306/a_36_216# OR2X1_LOC_306/Y VSS VDD
+ OR2X1_LOC_696/A OR2X1_LOC_22/Y OR2X1_LOC
XAND2X1_LOC_575 AND2X1_LOC_575/a_36_24# AND2X1_LOC_575/Y AND2X1_LOC_575/a_8_24# VSS VDD
+ AND2X1_LOC_573/Y AND2X1_LOC_574/Y AND2X1_LOC
XAND2X1_LOC_553 AND2X1_LOC_553/a_36_24# AND2X1_LOC_563/A AND2X1_LOC_553/a_8_24# VSS VDD
+ AND2X1_LOC_553/A AND2X1_LOC_541/Y AND2X1_LOC
XAND2X1_LOC_531 AND2X1_LOC_531/a_36_24# OR2X1_LOC_549/B AND2X1_LOC_531/a_8_24# VSS VDD
+ AND2X1_LOC_40/Y OR2X1_LOC_185/A AND2X1_LOC
XAND2X1_LOC_564 AND2X1_LOC_564/a_36_24# AND2X1_LOC_569/A AND2X1_LOC_564/a_8_24# VSS VDD
+ AND2X1_LOC_564/A AND2X1_LOC_564/B AND2X1_LOC
XAND2X1_LOC_520 AND2X1_LOC_520/a_36_24# AND2X1_LOC_520/Y AND2X1_LOC_520/a_8_24# VSS VDD
+ OR2X1_LOC_518/Y OR2X1_LOC_519/Y AND2X1_LOC
XAND2X1_LOC_542 AND2X1_LOC_542/a_36_24# AND2X1_LOC_552/A AND2X1_LOC_542/a_8_24# VSS VDD
+ OR2X1_LOC_280/Y OR2X1_LOC_312/Y AND2X1_LOC
XOR2X1_LOC_339 OR2X1_LOC_339/a_8_216# OR2X1_LOC_339/a_36_216# OR2X1_LOC_339/Y VSS VDD
+ OR2X1_LOC_339/A OR2X1_LOC_61/Y OR2X1_LOC
XOR2X1_LOC_317 OR2X1_LOC_317/a_8_216# OR2X1_LOC_317/a_36_216# OR2X1_LOC_319/B VSS VDD
+ OR2X1_LOC_317/A OR2X1_LOC_317/B OR2X1_LOC
XAND2X1_LOC_586 AND2X1_LOC_586/a_36_24# OR2X1_LOC_637/A AND2X1_LOC_586/a_8_24# VSS VDD
+ AND2X1_LOC_70/Y OR2X1_LOC_130/A AND2X1_LOC
XAND2X1_LOC_597 AND2X1_LOC_597/a_36_24# OR2X1_LOC_644/B AND2X1_LOC_597/a_8_24# VSS VDD
+ AND2X1_LOC_41/A OR2X1_LOC_596/Y AND2X1_LOC
XOR2X1_LOC_862 OR2X1_LOC_862/a_8_216# OR2X1_LOC_862/a_36_216# OR2X1_LOC_865/A VSS VDD
+ OR2X1_LOC_862/A OR2X1_LOC_862/B OR2X1_LOC
XOR2X1_LOC_840 OR2X1_LOC_840/a_8_216# OR2X1_LOC_840/a_36_216# OR2X1_LOC_851/B VSS VDD
+ OR2X1_LOC_840/A OR2X1_LOC_833/Y OR2X1_LOC
XOR2X1_LOC_851 OR2X1_LOC_851/a_8_216# OR2X1_LOC_851/a_36_216# OR2X1_LOC_858/A VSS VDD
+ OR2X1_LOC_851/A OR2X1_LOC_851/B OR2X1_LOC
XOR2X1_LOC_158 OR2X1_LOC_158/a_8_216# OR2X1_LOC_158/a_36_216# OR2X1_LOC_158/Y VSS VDD
+ OR2X1_LOC_158/A OR2X1_LOC_158/B OR2X1_LOC
XOR2X1_LOC_147 OR2X1_LOC_147/a_8_216# OR2X1_LOC_147/a_36_216# OR2X1_LOC_149/B VSS VDD
+ OR2X1_LOC_147/A OR2X1_LOC_147/B OR2X1_LOC
XAND2X1_LOC_361 AND2X1_LOC_361/a_36_24# AND2X1_LOC_362/B AND2X1_LOC_361/a_8_24# VSS VDD
+ AND2X1_LOC_361/A AND2X1_LOC_276/Y AND2X1_LOC
XAND2X1_LOC_372 AND2X1_LOC_372/a_36_24# OR2X1_LOC_458/B AND2X1_LOC_372/a_8_24# VSS VDD
+ D_INPUT_1 OR2X1_LOC_778/B AND2X1_LOC
XAND2X1_LOC_394 AND2X1_LOC_394/a_36_24# OR2X1_LOC_400/A AND2X1_LOC_394/a_8_24# VSS VDD
+ AND2X1_LOC_47/Y OR2X1_LOC_160/A AND2X1_LOC
XAND2X1_LOC_383 AND2X1_LOC_383/a_36_24# OR2X1_LOC_494/A AND2X1_LOC_383/a_8_24# VSS VDD
+ OR2X1_LOC_91/A OR2X1_LOC_428/A AND2X1_LOC
XAND2X1_LOC_350 AND2X1_LOC_350/a_36_24# AND2X1_LOC_350/Y AND2X1_LOC_350/a_8_24# VSS VDD
+ AND2X1_LOC_340/Y AND2X1_LOC_350/B AND2X1_LOC
XOR2X1_LOC_125 OR2X1_LOC_125/a_8_216# OR2X1_LOC_125/a_36_216# OR2X1_LOC_125/Y VSS VDD
+ OR2X1_LOC_600/A OR2X1_LOC_95/Y OR2X1_LOC
XOR2X1_LOC_114 OR2X1_LOC_114/a_8_216# OR2X1_LOC_114/a_36_216# OR2X1_LOC_114/Y VSS VDD
+ OR2X1_LOC_113/Y OR2X1_LOC_114/B OR2X1_LOC
XOR2X1_LOC_103 OR2X1_LOC_103/a_8_216# OR2X1_LOC_103/a_36_216# OR2X1_LOC_103/Y VSS VDD
+ OR2X1_LOC_485/A OR2X1_LOC_47/Y OR2X1_LOC
XOR2X1_LOC_169 OR2X1_LOC_169/a_8_216# OR2X1_LOC_169/a_36_216# OR2X1_LOC_170/A VSS VDD
+ OR2X1_LOC_703/B OR2X1_LOC_169/B OR2X1_LOC
XOR2X1_LOC_136 OR2X1_LOC_136/a_8_216# OR2X1_LOC_136/a_36_216# OR2X1_LOC_136/Y VSS VDD
+ OR2X1_LOC_43/A OR2X1_LOC_3/Y OR2X1_LOC
XAND2X1_LOC_90 AND2X1_LOC_90/a_36_24# AND2X1_LOC_91/B AND2X1_LOC_90/a_8_24# VSS VDD
+ AND2X1_LOC_42/B OR2X1_LOC_62/A AND2X1_LOC
XOR2X1_LOC_681 OR2X1_LOC_681/a_8_216# OR2X1_LOC_681/a_36_216# OR2X1_LOC_681/Y VSS VDD
+ OR2X1_LOC_743/A OR2X1_LOC_31/Y OR2X1_LOC
XOR2X1_LOC_692 OR2X1_LOC_692/a_8_216# OR2X1_LOC_692/a_36_216# OR2X1_LOC_692/Y VSS VDD
+ OR2X1_LOC_48/B OR2X1_LOC_18/Y OR2X1_LOC
XOR2X1_LOC_670 OR2X1_LOC_670/a_8_216# OR2X1_LOC_670/a_36_216# OR2X1_LOC_670/Y VSS VDD
+ OR2X1_LOC_485/A OR2X1_LOC_40/Y OR2X1_LOC
XAND2X1_LOC_191 AND2X1_LOC_191/a_36_24# AND2X1_LOC_191/Y AND2X1_LOC_191/a_8_24# VSS VDD
+ OR2X1_LOC_187/Y AND2X1_LOC_191/B AND2X1_LOC
XAND2X1_LOC_180 AND2X1_LOC_180/a_36_24# AND2X1_LOC_182/A AND2X1_LOC_180/a_8_24# VSS VDD
+ OR2X1_LOC_176/Y OR2X1_LOC_177/Y AND2X1_LOC
XAND2X1_LOC_735 AND2X1_LOC_735/a_36_24# AND2X1_LOC_735/Y AND2X1_LOC_735/a_8_24# VSS VDD
+ AND2X1_LOC_501/Y AND2X1_LOC_658/B AND2X1_LOC
XAND2X1_LOC_757 AND2X1_LOC_757/a_36_24# OR2X1_LOC_791/A AND2X1_LOC_757/a_8_24# VSS VDD
+ AND2X1_LOC_44/Y OR2X1_LOC_756/Y AND2X1_LOC
XAND2X1_LOC_702 AND2X1_LOC_702/a_36_24# AND2X1_LOC_702/Y AND2X1_LOC_702/a_8_24# VSS VDD
+ OR2X1_LOC_45/Y OR2X1_LOC_135/Y AND2X1_LOC
XAND2X1_LOC_746 AND2X1_LOC_746/a_36_24# OR2X1_LOC_781/A AND2X1_LOC_746/a_8_24# VSS VDD
+ OR2X1_LOC_185/A OR2X1_LOC_375/A AND2X1_LOC
XAND2X1_LOC_724 AND2X1_LOC_724/a_36_24# AND2X1_LOC_724/Y AND2X1_LOC_724/a_8_24# VSS VDD
+ AND2X1_LOC_724/A AND2X1_LOC_715/Y AND2X1_LOC
XAND2X1_LOC_713 AND2X1_LOC_713/a_36_24# AND2X1_LOC_713/Y AND2X1_LOC_713/a_8_24# VSS VDD
+ AND2X1_LOC_705/Y AND2X1_LOC_706/Y AND2X1_LOC
XAND2X1_LOC_768 AND2X1_LOC_768/a_36_24# AND2X1_LOC_772/B AND2X1_LOC_768/a_8_24# VSS VDD
+ OR2X1_LOC_103/Y OR2X1_LOC_134/Y AND2X1_LOC
XAND2X1_LOC_779 AND2X1_LOC_779/a_36_24# AND2X1_LOC_779/Y AND2X1_LOC_779/a_8_24# VSS VDD
+ OR2X1_LOC_511/Y OR2X1_LOC_697/Y AND2X1_LOC
XOR2X1_LOC_307 OR2X1_LOC_307/a_8_216# OR2X1_LOC_307/a_36_216# OR2X1_LOC_308/A VSS VDD
+ OR2X1_LOC_307/A OR2X1_LOC_307/B OR2X1_LOC
XOR2X1_LOC_329 OR2X1_LOC_329/a_8_216# OR2X1_LOC_329/a_36_216# OR2X1_LOC_329/Y VSS VDD
+ OR2X1_LOC_421/A OR2X1_LOC_329/B OR2X1_LOC
XAND2X1_LOC_510 AND2X1_LOC_510/a_36_24# AND2X1_LOC_574/A AND2X1_LOC_510/a_8_24# VSS VDD
+ AND2X1_LOC_510/A AND2X1_LOC_509/Y AND2X1_LOC
XAND2X1_LOC_576 AND2X1_LOC_576/a_36_24# AND2X1_LOC_576/Y AND2X1_LOC_576/a_8_24# VSS VDD
+ AND2X1_LOC_571/Y AND2X1_LOC_572/Y AND2X1_LOC
XAND2X1_LOC_554 AND2X1_LOC_554/a_36_24# AND2X1_LOC_554/Y AND2X1_LOC_554/a_8_24# VSS VDD
+ OR2X1_LOC_106/Y AND2X1_LOC_554/B AND2X1_LOC
XAND2X1_LOC_521 AND2X1_LOC_521/a_36_24# OR2X1_LOC_523/B AND2X1_LOC_521/a_8_24# VSS VDD
+ AND2X1_LOC_18/Y OR2X1_LOC_87/A AND2X1_LOC
XAND2X1_LOC_565 AND2X1_LOC_565/a_36_24# AND2X1_LOC_565/Y AND2X1_LOC_565/a_8_24# VSS VDD
+ AND2X1_LOC_549/Y AND2X1_LOC_565/B AND2X1_LOC
XAND2X1_LOC_543 AND2X1_LOC_543/a_36_24# AND2X1_LOC_543/Y AND2X1_LOC_543/a_8_24# VSS VDD
+ OR2X1_LOC_315/Y OR2X1_LOC_369/Y AND2X1_LOC
XAND2X1_LOC_532 AND2X1_LOC_532/a_36_24# OR2X1_LOC_533/A AND2X1_LOC_532/a_8_24# VSS VDD
+ OR2X1_LOC_485/A OR2X1_LOC_744/A AND2X1_LOC
XAND2X1_LOC_598 AND2X1_LOC_598/a_36_24# OR2X1_LOC_599/A AND2X1_LOC_598/a_8_24# VSS VDD
+ OR2X1_LOC_48/B OR2X1_LOC_585/A AND2X1_LOC
XAND2X1_LOC_587 AND2X1_LOC_587/a_36_24# AND2X1_LOC_588/B AND2X1_LOC_587/a_8_24# VSS VDD
+ D_INPUT_7 AND2X1_LOC_51/A AND2X1_LOC
XOR2X1_LOC_318 OR2X1_LOC_318/a_8_216# OR2X1_LOC_318/a_36_216# OR2X1_LOC_318/Y VSS VDD
+ OR2X1_LOC_318/A OR2X1_LOC_318/B OR2X1_LOC
XOR2X1_LOC_830 OR2X1_LOC_830/a_8_216# OR2X1_LOC_830/a_36_216# OR2X1_LOC_842/A VSS VDD
+ OR2X1_LOC_147/B OR2X1_LOC_114/B OR2X1_LOC
XOR2X1_LOC_841 OR2X1_LOC_841/a_8_216# OR2X1_LOC_841/a_36_216# OR2X1_LOC_851/A VSS VDD
+ OR2X1_LOC_841/A OR2X1_LOC_841/B OR2X1_LOC
XOR2X1_LOC_863 OR2X1_LOC_863/a_8_216# OR2X1_LOC_863/a_36_216# OR2X1_LOC_864/A VSS VDD
+ OR2X1_LOC_863/A OR2X1_LOC_863/B OR2X1_LOC
XOR2X1_LOC_852 OR2X1_LOC_852/a_8_216# OR2X1_LOC_852/a_36_216# OR2X1_LOC_857/B VSS VDD
+ OR2X1_LOC_852/A OR2X1_LOC_852/B OR2X1_LOC
XOR2X1_LOC_104 OR2X1_LOC_104/a_8_216# OR2X1_LOC_104/a_36_216# OR2X1_LOC_600/A VSS VDD
+ OR2X1_LOC_8/Y OR2X1_LOC_6/B OR2X1_LOC
XOR2X1_LOC_115 OR2X1_LOC_115/a_8_216# OR2X1_LOC_115/a_36_216# OR2X1_LOC_116/A VSS VDD
+ OR2X1_LOC_715/B OR2X1_LOC_115/B OR2X1_LOC
XOR2X1_LOC_126 OR2X1_LOC_126/a_8_216# OR2X1_LOC_126/a_36_216# OR2X1_LOC_744/A VSS VDD
+ OR2X1_LOC_85/A OR2X1_LOC_6/B OR2X1_LOC
XOR2X1_LOC_148 OR2X1_LOC_148/a_8_216# OR2X1_LOC_148/a_36_216# OR2X1_LOC_148/Y VSS VDD
+ OR2X1_LOC_148/A OR2X1_LOC_148/B OR2X1_LOC
XAND2X1_LOC_340 AND2X1_LOC_340/a_36_24# AND2X1_LOC_340/Y AND2X1_LOC_340/a_8_24# VSS VDD
+ OR2X1_LOC_88/Y AND2X1_LOC_227/Y AND2X1_LOC
XAND2X1_LOC_362 AND2X1_LOC_362/a_36_24# AND2X1_LOC_366/A AND2X1_LOC_362/a_8_24# VSS VDD
+ AND2X1_LOC_806/A AND2X1_LOC_362/B AND2X1_LOC
XAND2X1_LOC_384 AND2X1_LOC_384/a_36_24# OR2X1_LOC_391/A AND2X1_LOC_384/a_8_24# VSS VDD
+ AND2X1_LOC_40/Y OR2X1_LOC_383/Y AND2X1_LOC
XAND2X1_LOC_395 AND2X1_LOC_395/a_36_24# OR2X1_LOC_401/B AND2X1_LOC_395/a_8_24# VSS VDD
+ AND2X1_LOC_59/Y OR2X1_LOC_756/B AND2X1_LOC
XAND2X1_LOC_373 AND2X1_LOC_373/a_36_24# OR2X1_LOC_544/B AND2X1_LOC_373/a_8_24# VSS VDD
+ OR2X1_LOC_66/A OR2X1_LOC_78/A AND2X1_LOC
XAND2X1_LOC_351 AND2X1_LOC_351/a_36_24# AND2X1_LOC_351/Y AND2X1_LOC_351/a_8_24# VSS VDD
+ AND2X1_LOC_338/Y AND2X1_LOC_339/Y AND2X1_LOC
XOR2X1_LOC_159 OR2X1_LOC_159/a_8_216# OR2X1_LOC_159/a_36_216# OR2X1_LOC_604/A VSS VDD
+ OR2X1_LOC_9/Y OR2X1_LOC_6/A OR2X1_LOC
XOR2X1_LOC_137 OR2X1_LOC_137/a_8_216# OR2X1_LOC_137/a_36_216# OR2X1_LOC_137/Y VSS VDD
+ OR2X1_LOC_768/A OR2X1_LOC_137/B OR2X1_LOC
XAND2X1_LOC_80 AND2X1_LOC_80/a_36_24# AND2X1_LOC_81/B AND2X1_LOC_80/a_8_24# VSS VDD
+ OR2X1_LOC_68/B OR2X1_LOC_49/A AND2X1_LOC
XAND2X1_LOC_91 AND2X1_LOC_91/a_36_24# OR2X1_LOC_97/A AND2X1_LOC_91/a_8_24# VSS VDD
+ AND2X1_LOC_51/Y AND2X1_LOC_91/B AND2X1_LOC
XOR2X1_LOC_671 OR2X1_LOC_671/a_8_216# OR2X1_LOC_671/a_36_216# OR2X1_LOC_671/Y VSS VDD
+ OR2X1_LOC_6/B D_INPUT_2 OR2X1_LOC
XOR2X1_LOC_660 OR2X1_LOC_660/a_8_216# OR2X1_LOC_660/a_36_216# OR2X1_LOC_660/Y VSS VDD
+ OR2X1_LOC_656/Y OR2X1_LOC_660/B OR2X1_LOC
XOR2X1_LOC_682 OR2X1_LOC_682/a_8_216# OR2X1_LOC_682/a_36_216# OR2X1_LOC_682/Y VSS VDD
+ OR2X1_LOC_604/A OR2X1_LOC_36/Y OR2X1_LOC
XOR2X1_LOC_693 OR2X1_LOC_693/a_8_216# OR2X1_LOC_693/a_36_216# OR2X1_LOC_693/Y VSS VDD
+ OR2X1_LOC_36/Y OR2X1_LOC_46/A OR2X1_LOC
XAND2X1_LOC_181 AND2X1_LOC_181/a_36_24# AND2X1_LOC_181/Y AND2X1_LOC_181/a_8_24# VSS VDD
+ OR2X1_LOC_178/Y OR2X1_LOC_179/Y AND2X1_LOC
XAND2X1_LOC_170 AND2X1_LOC_170/a_36_24# AND2X1_LOC_170/Y AND2X1_LOC_170/a_8_24# VSS VDD
+ AND2X1_LOC_168/Y AND2X1_LOC_170/B AND2X1_LOC
XAND2X1_LOC_192 AND2X1_LOC_192/a_36_24# AND2X1_LOC_192/Y AND2X1_LOC_192/a_8_24# VSS VDD
+ OR2X1_LOC_189/Y AND2X1_LOC_191/Y AND2X1_LOC
XOR2X1_LOC_490 OR2X1_LOC_490/a_8_216# OR2X1_LOC_490/a_36_216# OR2X1_LOC_490/Y VSS VDD
+ OR2X1_LOC_86/A OR2X1_LOC_19/B OR2X1_LOC
XAND2X1_LOC_758 AND2X1_LOC_758/a_36_24# OR2X1_LOC_759/A AND2X1_LOC_758/a_8_24# VSS VDD
+ OR2X1_LOC_40/Y OR2X1_LOC_95/Y AND2X1_LOC
XAND2X1_LOC_736 AND2X1_LOC_736/a_36_24# AND2X1_LOC_736/Y AND2X1_LOC_736/a_8_24# VSS VDD
+ AND2X1_LOC_675/Y AND2X1_LOC_735/Y AND2X1_LOC
XAND2X1_LOC_703 AND2X1_LOC_703/a_36_24# AND2X1_LOC_703/Y AND2X1_LOC_703/a_8_24# VSS VDD
+ OR2X1_LOC_167/Y OR2X1_LOC_312/Y AND2X1_LOC
XAND2X1_LOC_747 AND2X1_LOC_747/a_36_24# OR2X1_LOC_782/B AND2X1_LOC_747/a_8_24# VSS VDD
+ AND2X1_LOC_47/Y OR2X1_LOC_87/A AND2X1_LOC
XAND2X1_LOC_769 AND2X1_LOC_769/a_36_24# AND2X1_LOC_769/Y AND2X1_LOC_769/a_8_24# VSS VDD
+ OR2X1_LOC_763/Y OR2X1_LOC_764/Y AND2X1_LOC
XAND2X1_LOC_714 AND2X1_LOC_714/a_36_24# AND2X1_LOC_724/A AND2X1_LOC_714/a_8_24# VSS VDD
+ AND2X1_LOC_703/Y AND2X1_LOC_714/B AND2X1_LOC
XAND2X1_LOC_725 AND2X1_LOC_725/a_36_24# AND2X1_LOC_732/B AND2X1_LOC_725/a_8_24# VSS VDD
+ AND2X1_LOC_712/Y AND2X1_LOC_713/Y AND2X1_LOC
XOR2X1_LOC_308 OR2X1_LOC_308/a_8_216# OR2X1_LOC_308/a_36_216# OR2X1_LOC_308/Y VSS VDD
+ OR2X1_LOC_308/A OR2X1_LOC_512/A OR2X1_LOC
XAND2X1_LOC_500 AND2X1_LOC_500/a_36_24# AND2X1_LOC_500/Y AND2X1_LOC_500/a_8_24# VSS VDD
+ OR2X1_LOC_497/Y AND2X1_LOC_500/B AND2X1_LOC
XAND2X1_LOC_522 AND2X1_LOC_522/a_36_24# OR2X1_LOC_523/A AND2X1_LOC_522/a_8_24# VSS VDD
+ AND2X1_LOC_22/Y OR2X1_LOC_532/B AND2X1_LOC
XAND2X1_LOC_555 AND2X1_LOC_555/a_36_24# AND2X1_LOC_555/Y AND2X1_LOC_555/a_8_24# VSS VDD
+ AND2X1_LOC_259/Y OR2X1_LOC_481/Y AND2X1_LOC
XAND2X1_LOC_577 AND2X1_LOC_577/a_36_24# AND2X1_LOC_577/Y AND2X1_LOC_577/a_8_24# VSS VDD
+ AND2X1_LOC_577/A AND2X1_LOC_570/Y AND2X1_LOC
XAND2X1_LOC_544 AND2X1_LOC_544/a_36_24# AND2X1_LOC_544/Y AND2X1_LOC_544/a_8_24# VSS VDD
+ OR2X1_LOC_373/Y OR2X1_LOC_438/Y AND2X1_LOC
XAND2X1_LOC_533 AND2X1_LOC_533/a_36_24# OR2X1_LOC_788/B AND2X1_LOC_533/a_8_24# VSS VDD
+ AND2X1_LOC_95/Y OR2X1_LOC_532/Y AND2X1_LOC
XAND2X1_LOC_566 AND2X1_LOC_566/a_36_24# AND2X1_LOC_566/Y AND2X1_LOC_566/a_8_24# VSS VDD
+ AND2X1_LOC_170/Y AND2X1_LOC_566/B AND2X1_LOC
XAND2X1_LOC_599 AND2X1_LOC_599/a_36_24# OR2X1_LOC_644/A AND2X1_LOC_599/a_8_24# VSS VDD
+ AND2X1_LOC_36/Y OR2X1_LOC_598/Y AND2X1_LOC
XAND2X1_LOC_511 AND2X1_LOC_511/a_36_24# OR2X1_LOC_779/B AND2X1_LOC_511/a_8_24# VSS VDD
+ AND2X1_LOC_31/Y AND2X1_LOC_48/A AND2X1_LOC
XAND2X1_LOC_588 AND2X1_LOC_588/a_36_24# OR2X1_LOC_638/B AND2X1_LOC_588/a_8_24# VSS VDD
+ OR2X1_LOC_502/A AND2X1_LOC_588/B AND2X1_LOC
XOR2X1_LOC_319 OR2X1_LOC_319/a_8_216# OR2X1_LOC_319/a_36_216# OR2X1_LOC_319/Y VSS VDD
+ OR2X1_LOC_318/Y OR2X1_LOC_319/B OR2X1_LOC
XOR2X1_LOC_864 OR2X1_LOC_864/a_8_216# OR2X1_LOC_864/a_36_216# OR2X1_LOC_866/B VSS VDD
+ OR2X1_LOC_864/A OR2X1_LOC_774/Y OR2X1_LOC
XOR2X1_LOC_820 OR2X1_LOC_820/a_8_216# OR2X1_LOC_820/a_36_216# OR2X1_LOC_820/Y VSS VDD
+ OR2X1_LOC_820/A OR2X1_LOC_820/B OR2X1_LOC
XOR2X1_LOC_842 OR2X1_LOC_842/a_8_216# OR2X1_LOC_842/a_36_216# OR2X1_LOC_850/B VSS VDD
+ OR2X1_LOC_842/A OR2X1_LOC_190/A OR2X1_LOC
XOR2X1_LOC_831 OR2X1_LOC_831/a_8_216# OR2X1_LOC_831/a_36_216# OR2X1_LOC_841/B VSS VDD
+ OR2X1_LOC_831/A OR2X1_LOC_831/B OR2X1_LOC
XOR2X1_LOC_853 OR2X1_LOC_853/a_8_216# OR2X1_LOC_853/a_36_216# OR2X1_LOC_857/A VSS VDD
+ OR2X1_LOC_175/Y OR2X1_LOC_35/Y OR2X1_LOC
XOR2X1_LOC_149 OR2X1_LOC_149/a_8_216# OR2X1_LOC_149/a_36_216# OR2X1_LOC_797/B VSS VDD
+ OR2X1_LOC_148/Y OR2X1_LOC_149/B OR2X1_LOC
XAND2X1_LOC_330 AND2X1_LOC_330/a_36_24# OR2X1_LOC_331/A AND2X1_LOC_330/a_8_24# VSS VDD
+ OR2X1_LOC_51/Y OR2X1_LOC_70/Y AND2X1_LOC
XOR2X1_LOC_105 OR2X1_LOC_105/a_8_216# OR2X1_LOC_105/a_36_216# OR2X1_LOC_105/Y VSS VDD
+ OR2X1_LOC_756/B OR2X1_LOC_78/A OR2X1_LOC
XOR2X1_LOC_127 OR2X1_LOC_127/a_8_216# OR2X1_LOC_127/a_36_216# OR2X1_LOC_127/Y VSS VDD
+ OR2X1_LOC_744/A OR2X1_LOC_3/Y OR2X1_LOC
XOR2X1_LOC_116 OR2X1_LOC_116/a_8_216# OR2X1_LOC_116/a_36_216# OR2X1_LOC_216/A VSS VDD
+ OR2X1_LOC_116/A OR2X1_LOC_114/Y OR2X1_LOC
XOR2X1_LOC_138 OR2X1_LOC_138/a_8_216# OR2X1_LOC_138/a_36_216# OR2X1_LOC_139/A VSS VDD
+ OR2X1_LOC_138/A OR2X1_LOC_702/A OR2X1_LOC
XAND2X1_LOC_363 AND2X1_LOC_363/a_36_24# AND2X1_LOC_363/Y AND2X1_LOC_363/a_8_24# VSS VDD
+ AND2X1_LOC_363/A AND2X1_LOC_363/B AND2X1_LOC
XAND2X1_LOC_396 AND2X1_LOC_396/a_36_24# OR2X1_LOC_401/A AND2X1_LOC_396/a_8_24# VSS VDD
+ OR2X1_LOC_160/B AND2X1_LOC_36/Y AND2X1_LOC
XAND2X1_LOC_374 AND2X1_LOC_374/a_36_24# AND2X1_LOC_374/Y AND2X1_LOC_374/a_8_24# VSS VDD
+ OR2X1_LOC_322/Y OR2X1_LOC_373/Y AND2X1_LOC
XAND2X1_LOC_385 AND2X1_LOC_385/a_36_24# OR2X1_LOC_389/B AND2X1_LOC_385/a_8_24# VSS VDD
+ OR2X1_LOC_66/A OR2X1_LOC_756/B AND2X1_LOC
XAND2X1_LOC_341 AND2X1_LOC_341/a_36_24# AND2X1_LOC_350/B AND2X1_LOC_341/a_8_24# VSS VDD
+ AND2X1_LOC_228/Y AND2X1_LOC_231/Y AND2X1_LOC
XAND2X1_LOC_352 AND2X1_LOC_352/a_36_24# AND2X1_LOC_357/A AND2X1_LOC_352/a_8_24# VSS VDD
+ AND2X1_LOC_212/A AND2X1_LOC_352/B AND2X1_LOC
XAND2X1_LOC_70 AND2X1_LOC_70/a_36_24# AND2X1_LOC_70/Y AND2X1_LOC_70/a_8_24# VSS VDD
+ AND2X1_LOC_2/Y AND2X1_LOC_50/Y AND2X1_LOC
XOR2X1_LOC_683 OR2X1_LOC_683/a_8_216# OR2X1_LOC_683/a_36_216# OR2X1_LOC_683/Y VSS VDD
+ OR2X1_LOC_22/Y OR2X1_LOC_16/A OR2X1_LOC
XOR2X1_LOC_694 OR2X1_LOC_694/a_8_216# OR2X1_LOC_694/a_36_216# OR2X1_LOC_694/Y VSS VDD
+ OR2X1_LOC_426/A OR2X1_LOC_427/A OR2X1_LOC
XAND2X1_LOC_81 AND2X1_LOC_81/a_36_24# OR2X1_LOC_84/B AND2X1_LOC_81/a_8_24# VSS VDD
+ AND2X1_LOC_59/Y AND2X1_LOC_81/B AND2X1_LOC
XAND2X1_LOC_92 AND2X1_LOC_92/a_36_24# AND2X1_LOC_92/Y AND2X1_LOC_92/a_8_24# VSS VDD
+ INPUT_1 AND2X1_LOC_8/Y AND2X1_LOC
XOR2X1_LOC_672 OR2X1_LOC_672/a_8_216# OR2X1_LOC_672/a_36_216# OR2X1_LOC_672/Y VSS VDD
+ OR2X1_LOC_671/Y OR2X1_LOC_158/A OR2X1_LOC
XOR2X1_LOC_650 OR2X1_LOC_650/a_8_216# OR2X1_LOC_650/a_36_216# OR2X1_LOC_650/Y VSS VDD
+ OR2X1_LOC_641/Y OR2X1_LOC_640/Y OR2X1_LOC
XOR2X1_LOC_661 OR2X1_LOC_661/a_8_216# OR2X1_LOC_661/a_36_216# OR2X1_LOC_662/A VSS VDD
+ OR2X1_LOC_661/A OR2X1_LOC_653/Y OR2X1_LOC
XAND2X1_LOC_171 AND2X1_LOC_171/a_36_24# OR2X1_LOC_333/B AND2X1_LOC_171/a_8_24# VSS VDD
+ OR2X1_LOC_160/B AND2X1_LOC_40/Y AND2X1_LOC
XAND2X1_LOC_182 AND2X1_LOC_182/a_36_24# AND2X1_LOC_212/A AND2X1_LOC_182/a_8_24# VSS VDD
+ AND2X1_LOC_182/A AND2X1_LOC_181/Y AND2X1_LOC
XAND2X1_LOC_160 AND2X1_LOC_160/a_36_24# AND2X1_LOC_160/Y AND2X1_LOC_160/a_8_24# VSS VDD
+ OR2X1_LOC_45/B OR2X1_LOC_744/A AND2X1_LOC
XAND2X1_LOC_193 AND2X1_LOC_193/a_36_24# AND2X1_LOC_193/Y AND2X1_LOC_193/a_8_24# VSS VDD
+ OR2X1_LOC_7/Y OR2X1_LOC_13/Y AND2X1_LOC
XOR2X1_LOC_480 OR2X1_LOC_480/a_8_216# OR2X1_LOC_480/a_36_216# D_GATE_479 VSS VDD
+ OR2X1_LOC_479/Y OR2X1_LOC_478/Y OR2X1_LOC
XOR2X1_LOC_491 OR2X1_LOC_491/a_8_216# OR2X1_LOC_491/a_36_216# OR2X1_LOC_491/Y VSS VDD
+ OR2X1_LOC_485/A OR2X1_LOC_31/Y OR2X1_LOC
XAND2X1_LOC_759 AND2X1_LOC_759/a_36_24# OR2X1_LOC_792/B AND2X1_LOC_759/a_8_24# VSS VDD
+ OR2X1_LOC_269/B OR2X1_LOC_758/Y AND2X1_LOC
XAND2X1_LOC_737 AND2X1_LOC_737/a_36_24# AND2X1_LOC_737/Y AND2X1_LOC_737/a_8_24# VSS VDD
+ AND2X1_LOC_733/Y AND2X1_LOC_734/Y AND2X1_LOC
XAND2X1_LOC_748 AND2X1_LOC_748/a_36_24# OR2X1_LOC_789/B AND2X1_LOC_748/a_8_24# VSS VDD
+ OR2X1_LOC_19/B OR2X1_LOC_709/A AND2X1_LOC
XAND2X1_LOC_715 AND2X1_LOC_715/a_36_24# AND2X1_LOC_715/Y AND2X1_LOC_715/a_8_24# VSS VDD
+ AND2X1_LOC_715/A AND2X1_LOC_702/Y AND2X1_LOC
XAND2X1_LOC_726 AND2X1_LOC_726/a_36_24# AND2X1_LOC_726/Y AND2X1_LOC_726/a_8_24# VSS VDD
+ OR2X1_LOC_152/Y AND2X1_LOC_711/Y AND2X1_LOC
XAND2X1_LOC_704 AND2X1_LOC_704/a_36_24# AND2X1_LOC_714/B AND2X1_LOC_704/a_8_24# VSS VDD
+ OR2X1_LOC_313/Y OR2X1_LOC_417/Y AND2X1_LOC
XAND2X1_LOC_501 AND2X1_LOC_501/a_36_24# AND2X1_LOC_501/Y AND2X1_LOC_501/a_8_24# VSS VDD
+ OR2X1_LOC_498/Y AND2X1_LOC_500/Y AND2X1_LOC
XAND2X1_LOC_523 AND2X1_LOC_523/a_36_24# AND2X1_LOC_523/Y AND2X1_LOC_523/a_8_24# VSS VDD
+ OR2X1_LOC_521/Y OR2X1_LOC_522/Y AND2X1_LOC
XAND2X1_LOC_512 AND2X1_LOC_512/a_36_24# AND2X1_LOC_512/Y AND2X1_LOC_512/a_8_24# VSS VDD
+ INPUT_0 OR2X1_LOC_306/Y AND2X1_LOC
XOR2X1_LOC_309 OR2X1_LOC_309/a_8_216# OR2X1_LOC_309/a_36_216# OR2X1_LOC_309/Y VSS VDD
+ OR2X1_LOC_417/A OR2X1_LOC_22/Y OR2X1_LOC
XAND2X1_LOC_556 AND2X1_LOC_556/a_36_24# AND2X1_LOC_562/B AND2X1_LOC_556/a_8_24# VSS VDD
+ AND2X1_LOC_483/Y AND2X1_LOC_486/Y AND2X1_LOC
XAND2X1_LOC_578 AND2X1_LOC_578/a_36_24# AND2X1_LOC_580/A AND2X1_LOC_578/a_8_24# VSS VDD
+ AND2X1_LOC_578/A AND2X1_LOC_577/Y AND2X1_LOC
XAND2X1_LOC_589 AND2X1_LOC_589/a_36_24# OR2X1_LOC_592/A AND2X1_LOC_589/a_8_24# VSS VDD
+ AND2X1_LOC_22/Y OR2X1_LOC_130/A AND2X1_LOC
XAND2X1_LOC_534 AND2X1_LOC_534/a_36_24# OR2X1_LOC_535/A AND2X1_LOC_534/a_8_24# VSS VDD
+ AND2X1_LOC_43/B AND2X1_LOC_59/Y AND2X1_LOC
XAND2X1_LOC_567 AND2X1_LOC_567/a_36_24# AND2X1_LOC_568/B AND2X1_LOC_567/a_8_24# VSS VDD
+ AND2X1_LOC_535/Y AND2X1_LOC_539/Y AND2X1_LOC
XAND2X1_LOC_545 AND2X1_LOC_545/a_36_24# AND2X1_LOC_551/B AND2X1_LOC_545/a_8_24# VSS VDD
+ OR2X1_LOC_441/Y OR2X1_LOC_524/Y AND2X1_LOC
XOR2X1_LOC_810 OR2X1_LOC_810/a_8_216# OR2X1_LOC_810/a_36_216# OR2X1_LOC_812/B VSS VDD
+ OR2X1_LOC_810/A OR2X1_LOC_774/Y OR2X1_LOC
XOR2X1_LOC_865 OR2X1_LOC_865/a_8_216# OR2X1_LOC_865/a_36_216# OR2X1_LOC_865/Y VSS VDD
+ OR2X1_LOC_865/A OR2X1_LOC_865/B OR2X1_LOC
XOR2X1_LOC_843 OR2X1_LOC_843/a_8_216# OR2X1_LOC_843/a_36_216# OR2X1_LOC_850/A VSS VDD
+ OR2X1_LOC_287/B OR2X1_LOC_843/B OR2X1_LOC
XOR2X1_LOC_821 OR2X1_LOC_821/a_8_216# OR2X1_LOC_821/a_36_216# OR2X1_LOC_821/Y VSS VDD
+ OR2X1_LOC_70/Y OR2X1_LOC_13/B OR2X1_LOC
XOR2X1_LOC_832 OR2X1_LOC_832/a_8_216# OR2X1_LOC_832/a_36_216# OR2X1_LOC_841/A VSS VDD
+ OR2X1_LOC_435/A OR2X1_LOC_449/B OR2X1_LOC
XOR2X1_LOC_854 OR2X1_LOC_854/a_8_216# OR2X1_LOC_854/a_36_216# OR2X1_LOC_856/B VSS VDD
+ OR2X1_LOC_854/A OR2X1_LOC_354/A OR2X1_LOC
XAND2X1_LOC_342 AND2X1_LOC_342/a_36_24# AND2X1_LOC_342/Y AND2X1_LOC_342/a_8_24# VSS VDD
+ OR2X1_LOC_246/Y OR2X1_LOC_248/Y AND2X1_LOC
XAND2X1_LOC_364 AND2X1_LOC_364/a_36_24# AND2X1_LOC_364/Y AND2X1_LOC_364/a_8_24# VSS VDD
+ AND2X1_LOC_364/A AND2X1_LOC_358/Y AND2X1_LOC
XAND2X1_LOC_353 AND2X1_LOC_353/a_36_24# AND2X1_LOC_357/B AND2X1_LOC_353/a_8_24# VSS VDD
+ AND2X1_LOC_566/B AND2X1_LOC_727/A AND2X1_LOC
XAND2X1_LOC_320 AND2X1_LOC_320/a_36_24# OR2X1_LOC_324/B AND2X1_LOC_320/a_8_24# VSS VDD
+ AND2X1_LOC_36/Y AND2X1_LOC_91/B AND2X1_LOC
XAND2X1_LOC_331 AND2X1_LOC_331/a_36_24# OR2X1_LOC_355/A AND2X1_LOC_331/a_8_24# VSS VDD
+ OR2X1_LOC_186/Y OR2X1_LOC_330/Y AND2X1_LOC
XOR2X1_LOC_128 OR2X1_LOC_128/a_8_216# OR2X1_LOC_128/a_36_216# OR2X1_LOC_140/B VSS VDD
+ OR2X1_LOC_128/A OR2X1_LOC_128/B OR2X1_LOC
XOR2X1_LOC_139 OR2X1_LOC_139/a_8_216# OR2X1_LOC_139/a_36_216# OR2X1_LOC_141/B VSS VDD
+ OR2X1_LOC_139/A OR2X1_LOC_137/Y OR2X1_LOC
XOR2X1_LOC_117 OR2X1_LOC_117/a_8_216# OR2X1_LOC_117/a_36_216# OR2X1_LOC_117/Y VSS VDD
+ OR2X1_LOC_70/Y OR2X1_LOC_65/B OR2X1_LOC
XOR2X1_LOC_106 OR2X1_LOC_106/a_8_216# OR2X1_LOC_106/a_36_216# OR2X1_LOC_106/Y VSS VDD
+ OR2X1_LOC_106/A OR2X1_LOC_47/Y OR2X1_LOC
XAND2X1_LOC_397 AND2X1_LOC_397/a_36_24# OR2X1_LOC_402/B AND2X1_LOC_397/a_8_24# VSS VDD
+ AND2X1_LOC_3/Y AND2X1_LOC_82/Y AND2X1_LOC
XAND2X1_LOC_375 AND2X1_LOC_375/a_36_24# OR2X1_LOC_376/A AND2X1_LOC_375/a_8_24# VSS VDD
+ OR2X1_LOC_31/Y OR2X1_LOC_158/A AND2X1_LOC
XAND2X1_LOC_386 AND2X1_LOC_386/a_36_24# AND2X1_LOC_387/B AND2X1_LOC_386/a_8_24# VSS VDD
+ D_INPUT_4 AND2X1_LOC_17/Y AND2X1_LOC
XAND2X1_LOC_93 AND2X1_LOC_93/a_36_24# OR2X1_LOC_98/B AND2X1_LOC_93/a_8_24# VSS VDD
+ OR2X1_LOC_66/A AND2X1_LOC_92/Y AND2X1_LOC
XAND2X1_LOC_71 AND2X1_LOC_71/a_36_24# AND2X1_LOC_72/B AND2X1_LOC_71/a_8_24# VSS VDD
+ OR2X1_LOC_68/B OR2X1_LOC_235/B AND2X1_LOC
XAND2X1_LOC_82 AND2X1_LOC_82/a_36_24# AND2X1_LOC_82/Y AND2X1_LOC_82/a_8_24# VSS VDD
+ OR2X1_LOC_377/A OR2X1_LOC_49/A AND2X1_LOC
XAND2X1_LOC_60 AND2X1_LOC_60/a_36_24# OR2X1_LOC_61/A AND2X1_LOC_60/a_8_24# VSS VDD
+ OR2X1_LOC_154/A AND2X1_LOC_59/Y AND2X1_LOC
XOR2X1_LOC_684 OR2X1_LOC_684/a_8_216# OR2X1_LOC_684/a_36_216# OR2X1_LOC_684/Y VSS VDD
+ OR2X1_LOC_43/A OR2X1_LOC_12/Y OR2X1_LOC
XOR2X1_LOC_695 OR2X1_LOC_695/a_8_216# OR2X1_LOC_695/a_36_216# OR2X1_LOC_695/Y VSS VDD
+ OR2X1_LOC_47/Y OR2X1_LOC_45/B OR2X1_LOC
XOR2X1_LOC_651 OR2X1_LOC_651/a_8_216# OR2X1_LOC_651/a_36_216# OR2X1_LOC_654/A VSS VDD
+ OR2X1_LOC_651/A OR2X1_LOC_651/B OR2X1_LOC
XOR2X1_LOC_673 OR2X1_LOC_673/a_8_216# OR2X1_LOC_673/a_36_216# OR2X1_LOC_673/Y VSS VDD
+ OR2X1_LOC_673/A OR2X1_LOC_673/B OR2X1_LOC
XOR2X1_LOC_662 OR2X1_LOC_662/a_8_216# OR2X1_LOC_662/a_36_216# OR2X1_LOC_663/A VSS VDD
+ OR2X1_LOC_662/A OR2X1_LOC_660/Y OR2X1_LOC
XOR2X1_LOC_640 OR2X1_LOC_640/a_8_216# OR2X1_LOC_640/a_36_216# OR2X1_LOC_640/Y VSS VDD
+ OR2X1_LOC_640/A OR2X1_LOC_633/Y OR2X1_LOC
XAND2X1_LOC_183 AND2X1_LOC_183/a_36_24# OR2X1_LOC_190/B AND2X1_LOC_183/a_8_24# VSS VDD
+ AND2X1_LOC_7/B AND2X1_LOC_40/Y AND2X1_LOC
XAND2X1_LOC_150 AND2X1_LOC_150/a_36_24# OR2X1_LOC_151/A AND2X1_LOC_150/a_8_24# VSS VDD
+ AND2X1_LOC_42/B OR2X1_LOC_235/B AND2X1_LOC
XAND2X1_LOC_172 AND2X1_LOC_172/a_36_24# OR2X1_LOC_174/A AND2X1_LOC_172/a_8_24# VSS VDD
+ AND2X1_LOC_70/Y OR2X1_LOC_532/B AND2X1_LOC
XAND2X1_LOC_194 AND2X1_LOC_194/a_36_24# AND2X1_LOC_194/Y AND2X1_LOC_194/a_8_24# VSS VDD
+ OR2X1_LOC_16/Y OR2X1_LOC_39/Y AND2X1_LOC
XAND2X1_LOC_161 AND2X1_LOC_161/a_36_24# AND2X1_LOC_161/Y AND2X1_LOC_161/a_8_24# VSS VDD
+ OR2X1_LOC_427/A OR2X1_LOC_604/A AND2X1_LOC
XOR2X1_LOC_470 OR2X1_LOC_470/a_8_216# OR2X1_LOC_470/a_36_216# OR2X1_LOC_477/B VSS VDD
+ OR2X1_LOC_470/A OR2X1_LOC_470/B OR2X1_LOC
XOR2X1_LOC_481 OR2X1_LOC_481/a_8_216# OR2X1_LOC_481/a_36_216# OR2X1_LOC_481/Y VSS VDD
+ OR2X1_LOC_481/A OR2X1_LOC_3/Y OR2X1_LOC
XOR2X1_LOC_492 OR2X1_LOC_492/a_8_216# OR2X1_LOC_492/a_36_216# OR2X1_LOC_492/Y VSS VDD
+ OR2X1_LOC_744/A OR2X1_LOC_59/Y OR2X1_LOC
XAND2X1_LOC_705 AND2X1_LOC_705/a_36_24# AND2X1_LOC_705/Y AND2X1_LOC_705/a_8_24# VSS VDD
+ OR2X1_LOC_485/Y OR2X1_LOC_526/Y AND2X1_LOC
XAND2X1_LOC_749 AND2X1_LOC_749/a_36_24# OR2X1_LOC_750/A AND2X1_LOC_749/a_8_24# VSS VDD
+ D_INPUT_0 AND2X1_LOC_8/Y AND2X1_LOC
XAND2X1_LOC_716 AND2X1_LOC_716/a_36_24# AND2X1_LOC_716/Y AND2X1_LOC_716/a_8_24# VSS VDD
+ AND2X1_LOC_228/Y AND2X1_LOC_303/A AND2X1_LOC
XAND2X1_LOC_727 AND2X1_LOC_727/a_36_24# AND2X1_LOC_727/Y AND2X1_LOC_727/a_8_24# VSS VDD
+ AND2X1_LOC_727/A AND2X1_LOC_727/B AND2X1_LOC
XAND2X1_LOC_738 AND2X1_LOC_738/a_36_24# AND2X1_LOC_738/Y AND2X1_LOC_738/a_8_24# VSS VDD
+ AND2X1_LOC_731/Y AND2X1_LOC_738/B AND2X1_LOC
XAND2X1_LOC_502 AND2X1_LOC_502/a_36_24# OR2X1_LOC_503/A AND2X1_LOC_502/a_8_24# VSS VDD
+ OR2X1_LOC_89/A OR2X1_LOC_696/A AND2X1_LOC
XAND2X1_LOC_557 AND2X1_LOC_557/a_36_24# AND2X1_LOC_557/Y AND2X1_LOC_557/a_8_24# VSS VDD
+ AND2X1_LOC_489/Y OR2X1_LOC_490/Y AND2X1_LOC
XAND2X1_LOC_524 AND2X1_LOC_524/a_36_24# OR2X1_LOC_545/A AND2X1_LOC_524/a_8_24# VSS VDD
+ AND2X1_LOC_47/Y OR2X1_LOC_161/B AND2X1_LOC
XAND2X1_LOC_535 AND2X1_LOC_535/a_36_24# AND2X1_LOC_535/Y AND2X1_LOC_535/a_8_24# VSS VDD
+ OR2X1_LOC_533/Y OR2X1_LOC_534/Y AND2X1_LOC
XAND2X1_LOC_513 AND2X1_LOC_513/a_36_24# OR2X1_LOC_516/B AND2X1_LOC_513/a_8_24# VSS VDD
+ OR2X1_LOC_511/Y AND2X1_LOC_512/Y AND2X1_LOC
XAND2X1_LOC_546 AND2X1_LOC_546/a_36_24# AND2X1_LOC_550/A AND2X1_LOC_546/a_8_24# VSS VDD
+ OR2X1_LOC_525/Y OR2X1_LOC_526/Y AND2X1_LOC
XAND2X1_LOC_579 AND2X1_LOC_579/a_36_24# AND2X1_LOC_580/B AND2X1_LOC_579/a_8_24# VSS VDD
+ AND2X1_LOC_575/Y AND2X1_LOC_576/Y AND2X1_LOC
XAND2X1_LOC_568 AND2X1_LOC_568/a_36_24# AND2X1_LOC_578/A AND2X1_LOC_568/a_8_24# VSS VDD
+ AND2X1_LOC_566/Y AND2X1_LOC_568/B AND2X1_LOC
XOR2X1_LOC_811 OR2X1_LOC_811/a_8_216# OR2X1_LOC_811/a_36_216# OR2X1_LOC_812/A VSS VDD
+ OR2X1_LOC_811/A OR2X1_LOC_807/Y OR2X1_LOC
XOR2X1_LOC_866 OR2X1_LOC_866/a_8_216# OR2X1_LOC_866/a_36_216# D_GATE_865 VSS VDD
+ OR2X1_LOC_865/Y OR2X1_LOC_866/B OR2X1_LOC
XOR2X1_LOC_844 OR2X1_LOC_844/a_8_216# OR2X1_LOC_844/a_36_216# OR2X1_LOC_844/Y VSS VDD
+ OR2X1_LOC_523/Y OR2X1_LOC_844/B OR2X1_LOC
XOR2X1_LOC_822 OR2X1_LOC_822/a_8_216# OR2X1_LOC_822/a_36_216# OR2X1_LOC_822/Y VSS VDD
+ OR2X1_LOC_485/A OR2X1_LOC_64/Y OR2X1_LOC
XOR2X1_LOC_833 OR2X1_LOC_833/a_8_216# OR2X1_LOC_833/a_36_216# OR2X1_LOC_833/Y VSS VDD
+ OR2X1_LOC_499/B OR2X1_LOC_833/B OR2X1_LOC
XOR2X1_LOC_800 OR2X1_LOC_800/a_8_216# OR2X1_LOC_800/a_36_216# OR2X1_LOC_800/Y VSS VDD
+ OR2X1_LOC_800/A OR2X1_LOC_687/Y OR2X1_LOC
XOR2X1_LOC_855 OR2X1_LOC_855/a_8_216# OR2X1_LOC_855/a_36_216# OR2X1_LOC_856/A VSS VDD
+ OR2X1_LOC_855/A OR2X1_LOC_691/Y OR2X1_LOC
XAND2X1_LOC_310 AND2X1_LOC_310/a_36_24# OR2X1_LOC_335/A AND2X1_LOC_310/a_8_24# VSS VDD
+ OR2X1_LOC_68/B AND2X1_LOC_40/Y AND2X1_LOC
XAND2X1_LOC_398 AND2X1_LOC_398/a_36_24# OR2X1_LOC_399/A AND2X1_LOC_398/a_8_24# VSS VDD
+ OR2X1_LOC_16/A OR2X1_LOC_585/A AND2X1_LOC
XAND2X1_LOC_343 AND2X1_LOC_343/a_36_24# AND2X1_LOC_349/B AND2X1_LOC_343/a_8_24# VSS VDD
+ OR2X1_LOC_250/Y OR2X1_LOC_251/Y AND2X1_LOC
XAND2X1_LOC_332 AND2X1_LOC_332/a_36_24# AND2X1_LOC_339/B AND2X1_LOC_332/a_8_24# VSS VDD
+ OR2X1_LOC_111/Y OR2X1_LOC_135/Y AND2X1_LOC
XAND2X1_LOC_387 AND2X1_LOC_387/a_36_24# OR2X1_LOC_389/A AND2X1_LOC_387/a_8_24# VSS VDD
+ AND2X1_LOC_92/Y AND2X1_LOC_387/B AND2X1_LOC
XAND2X1_LOC_365 AND2X1_LOC_365/a_36_24# AND2X1_LOC_367/A AND2X1_LOC_365/a_8_24# VSS VDD
+ AND2X1_LOC_365/A AND2X1_LOC_364/Y AND2X1_LOC
XAND2X1_LOC_321 AND2X1_LOC_321/a_36_24# OR2X1_LOC_324/A AND2X1_LOC_321/a_8_24# VSS VDD
+ AND2X1_LOC_41/A AND2X1_LOC_64/Y AND2X1_LOC
XAND2X1_LOC_354 AND2X1_LOC_354/a_36_24# AND2X1_LOC_354/Y AND2X1_LOC_354/a_8_24# VSS VDD
+ AND2X1_LOC_798/A AND2X1_LOC_354/B AND2X1_LOC
XAND2X1_LOC_376 AND2X1_LOC_376/a_36_24# OR2X1_LOC_459/B AND2X1_LOC_376/a_8_24# VSS VDD
+ OR2X1_LOC_502/A OR2X1_LOC_375/Y AND2X1_LOC
XOR2X1_LOC_118 OR2X1_LOC_118/a_8_216# OR2X1_LOC_118/a_36_216# OR2X1_LOC_118/Y VSS VDD
+ OR2X1_LOC_89/A OR2X1_LOC_70/Y OR2X1_LOC
XOR2X1_LOC_129 OR2X1_LOC_129/a_8_216# OR2X1_LOC_129/a_36_216# OR2X1_LOC_589/A VSS VDD
+ OR2X1_LOC_85/A OR2X1_LOC_80/A OR2X1_LOC
XOR2X1_LOC_107 OR2X1_LOC_107/a_8_216# OR2X1_LOC_107/a_36_216# OR2X1_LOC_107/Y VSS VDD
+ OR2X1_LOC_89/A OR2X1_LOC_64/Y OR2X1_LOC
XAND2X1_LOC_94 AND2X1_LOC_94/a_36_24# AND2X1_LOC_94/Y AND2X1_LOC_94/a_8_24# VSS VDD
+ OR2X1_LOC_377/A OR2X1_LOC_54/Y AND2X1_LOC
XAND2X1_LOC_72 AND2X1_LOC_72/a_36_24# AND2X1_LOC_72/Y AND2X1_LOC_72/a_8_24# VSS VDD
+ AND2X1_LOC_70/Y AND2X1_LOC_72/B AND2X1_LOC
XAND2X1_LOC_83 AND2X1_LOC_83/a_36_24# OR2X1_LOC_84/A AND2X1_LOC_83/a_8_24# VSS VDD
+ OR2X1_LOC_66/A AND2X1_LOC_82/Y AND2X1_LOC
XAND2X1_LOC_61 AND2X1_LOC_61/a_36_24# AND2X1_LOC_61/Y AND2X1_LOC_61/a_8_24# VSS VDD
+ OR2X1_LOC_58/Y OR2X1_LOC_60/Y AND2X1_LOC
XAND2X1_LOC_50 AND2X1_LOC_50/a_36_24# AND2X1_LOC_50/Y AND2X1_LOC_50/a_8_24# VSS VDD
+ D_INPUT_6 D_INPUT_7 AND2X1_LOC
XOR2X1_LOC_630 OR2X1_LOC_630/a_8_216# OR2X1_LOC_630/a_36_216# OR2X1_LOC_630/Y VSS VDD
+ OR2X1_LOC_629/Y OR2X1_LOC_630/B OR2X1_LOC
XOR2X1_LOC_685 OR2X1_LOC_685/a_8_216# OR2X1_LOC_685/a_36_216# OR2X1_LOC_687/B VSS VDD
+ OR2X1_LOC_685/A OR2X1_LOC_685/B OR2X1_LOC
XOR2X1_LOC_696 OR2X1_LOC_696/a_8_216# OR2X1_LOC_696/a_36_216# OR2X1_LOC_696/Y VSS VDD
+ OR2X1_LOC_696/A OR2X1_LOC_26/Y OR2X1_LOC
XOR2X1_LOC_663 OR2X1_LOC_663/a_8_216# OR2X1_LOC_663/a_36_216# D_GATE_662 VSS VDD
+ OR2X1_LOC_663/A OR2X1_LOC_659/Y OR2X1_LOC
XOR2X1_LOC_641 OR2X1_LOC_641/a_8_216# OR2X1_LOC_641/a_36_216# OR2X1_LOC_641/Y VSS VDD
+ OR2X1_LOC_641/A OR2X1_LOC_641/B OR2X1_LOC
XOR2X1_LOC_674 OR2X1_LOC_674/a_8_216# OR2X1_LOC_674/a_36_216# OR2X1_LOC_674/Y VSS VDD
+ OR2X1_LOC_329/B OR2X1_LOC_70/Y OR2X1_LOC
XOR2X1_LOC_652 OR2X1_LOC_652/a_8_216# OR2X1_LOC_652/a_36_216# OR2X1_LOC_653/A VSS VDD
+ OR2X1_LOC_799/A OR2X1_LOC_468/A OR2X1_LOC
XAND2X1_LOC_140 AND2X1_LOC_140/a_36_24# AND2X1_LOC_141/B AND2X1_LOC_140/a_8_24# VSS VDD
+ AND2X1_LOC_554/B OR2X1_LOC_131/Y AND2X1_LOC
XAND2X1_LOC_184 AND2X1_LOC_184/a_36_24# OR2X1_LOC_190/A AND2X1_LOC_184/a_8_24# VSS VDD
+ AND2X1_LOC_72/B AND2X1_LOC_95/Y AND2X1_LOC
XAND2X1_LOC_173 AND2X1_LOC_173/a_36_24# OR2X1_LOC_175/B AND2X1_LOC_173/a_8_24# VSS VDD
+ AND2X1_LOC_70/Y OR2X1_LOC_151/A AND2X1_LOC
XAND2X1_LOC_151 AND2X1_LOC_151/a_36_24# OR2X1_LOC_152/A AND2X1_LOC_151/a_8_24# VSS VDD
+ OR2X1_LOC_56/A OR2X1_LOC_437/A AND2X1_LOC
XAND2X1_LOC_195 AND2X1_LOC_195/a_36_24# AND2X1_LOC_199/A AND2X1_LOC_195/a_8_24# VSS VDD
+ OR2X1_LOC_41/Y OR2X1_LOC_43/Y AND2X1_LOC
XAND2X1_LOC_162 AND2X1_LOC_162/a_36_24# OR2X1_LOC_163/A AND2X1_LOC_162/a_8_24# VSS VDD
+ AND2X1_LOC_160/Y AND2X1_LOC_161/Y AND2X1_LOC
XOR2X1_LOC_471 OR2X1_LOC_471/a_8_216# OR2X1_LOC_471/a_36_216# OR2X1_LOC_471/Y VSS VDD
+ OR2X1_LOC_465/Y OR2X1_LOC_471/B OR2X1_LOC
XOR2X1_LOC_460 OR2X1_LOC_460/a_8_216# OR2X1_LOC_460/a_36_216# OR2X1_LOC_460/Y VSS VDD
+ OR2X1_LOC_460/A OR2X1_LOC_460/B OR2X1_LOC
XOR2X1_LOC_482 OR2X1_LOC_482/a_8_216# OR2X1_LOC_482/a_36_216# OR2X1_LOC_482/Y VSS VDD
+ OR2X1_LOC_59/Y OR2X1_LOC_7/A OR2X1_LOC
XOR2X1_LOC_493 OR2X1_LOC_493/a_8_216# OR2X1_LOC_493/a_36_216# OR2X1_LOC_493/Y VSS VDD
+ OR2X1_LOC_493/A OR2X1_LOC_493/B OR2X1_LOC
XOR2X1_LOC_290 OR2X1_LOC_290/a_8_216# OR2X1_LOC_290/a_36_216# OR2X1_LOC_290/Y VSS VDD
+ OR2X1_LOC_26/Y OR2X1_LOC_16/A OR2X1_LOC
XAND2X1_LOC_717 AND2X1_LOC_717/a_36_24# AND2X1_LOC_717/Y AND2X1_LOC_717/a_8_24# VSS VDD
+ AND2X1_LOC_374/Y AND2X1_LOC_717/B AND2X1_LOC
XAND2X1_LOC_739 AND2X1_LOC_739/a_36_24# AND2X1_LOC_740/B AND2X1_LOC_739/a_8_24# VSS VDD
+ AND2X1_LOC_192/Y AND2X1_LOC_739/B AND2X1_LOC
XAND2X1_LOC_728 AND2X1_LOC_728/a_36_24# AND2X1_LOC_728/Y AND2X1_LOC_728/a_8_24# VSS VDD
+ OR2X1_LOC_679/Y OR2X1_LOC_680/Y AND2X1_LOC
XAND2X1_LOC_706 AND2X1_LOC_706/a_36_24# AND2X1_LOC_706/Y AND2X1_LOC_706/a_8_24# VSS VDD
+ OR2X1_LOC_692/Y OR2X1_LOC_693/Y AND2X1_LOC
XAND2X1_LOC_558 AND2X1_LOC_558/a_36_24# AND2X1_LOC_561/B AND2X1_LOC_558/a_8_24# VSS VDD
+ AND2X1_LOC_717/B OR2X1_LOC_494/Y AND2X1_LOC
XAND2X1_LOC_503 AND2X1_LOC_503/a_36_24# OR2X1_LOC_509/A AND2X1_LOC_503/a_8_24# VSS VDD
+ AND2X1_LOC_64/Y OR2X1_LOC_502/Y AND2X1_LOC
XAND2X1_LOC_569 AND2X1_LOC_569/a_36_24# AND2X1_LOC_577/A AND2X1_LOC_569/a_8_24# VSS VDD
+ AND2X1_LOC_569/A AND2X1_LOC_565/Y AND2X1_LOC
XAND2X1_LOC_547 AND2X1_LOC_547/a_36_24# AND2X1_LOC_547/Y AND2X1_LOC_547/a_8_24# VSS VDD
+ OR2X1_LOC_527/Y OR2X1_LOC_528/Y AND2X1_LOC
XAND2X1_LOC_514 AND2X1_LOC_514/a_36_24# AND2X1_LOC_514/Y AND2X1_LOC_514/a_8_24# VSS VDD
+ D_INPUT_0 OR2X1_LOC_136/Y AND2X1_LOC
XAND2X1_LOC_536 AND2X1_LOC_536/a_36_24# OR2X1_LOC_537/A AND2X1_LOC_536/a_8_24# VSS VDD
+ AND2X1_LOC_12/Y OR2X1_LOC_532/B AND2X1_LOC
XAND2X1_LOC_525 AND2X1_LOC_525/a_36_24# OR2X1_LOC_546/B AND2X1_LOC_525/a_8_24# VSS VDD
+ AND2X1_LOC_41/A AND2X1_LOC_51/Y AND2X1_LOC
XOR2X1_LOC_812 OR2X1_LOC_812/a_8_216# OR2X1_LOC_812/a_36_216# D_GATE_811 VSS VDD
+ OR2X1_LOC_812/A OR2X1_LOC_812/B OR2X1_LOC
XOR2X1_LOC_801 OR2X1_LOC_801/a_8_216# OR2X1_LOC_801/a_36_216# OR2X1_LOC_809/B VSS VDD
+ OR2X1_LOC_800/Y OR2X1_LOC_801/B OR2X1_LOC
XOR2X1_LOC_834 OR2X1_LOC_834/a_8_216# OR2X1_LOC_834/a_36_216# OR2X1_LOC_840/A VSS VDD
+ OR2X1_LOC_834/A OR2X1_LOC_779/B OR2X1_LOC
XOR2X1_LOC_823 OR2X1_LOC_823/a_8_216# OR2X1_LOC_823/a_36_216# OR2X1_LOC_823/Y VSS VDD
+ OR2X1_LOC_428/A OR2X1_LOC_51/Y OR2X1_LOC
XOR2X1_LOC_845 OR2X1_LOC_845/a_8_216# OR2X1_LOC_845/a_36_216# OR2X1_LOC_849/A VSS VDD
+ OR2X1_LOC_845/A OR2X1_LOC_673/Y OR2X1_LOC
XOR2X1_LOC_856 OR2X1_LOC_856/a_8_216# OR2X1_LOC_856/a_36_216# OR2X1_LOC_863/B VSS VDD
+ OR2X1_LOC_856/A OR2X1_LOC_856/B OR2X1_LOC
XAND2X1_LOC_300 AND2X1_LOC_300/a_36_24# OR2X1_LOC_831/A AND2X1_LOC_300/a_8_24# VSS VDD
+ AND2X1_LOC_59/Y OR2X1_LOC_121/B AND2X1_LOC
XAND2X1_LOC_366 AND2X1_LOC_366/a_36_24# AND2X1_LOC_367/B AND2X1_LOC_366/a_8_24# VSS VDD
+ AND2X1_LOC_366/A AND2X1_LOC_363/Y AND2X1_LOC
XAND2X1_LOC_344 AND2X1_LOC_344/a_36_24# AND2X1_LOC_348/A AND2X1_LOC_344/a_8_24# VSS VDD
+ AND2X1_LOC_456/B OR2X1_LOC_256/Y AND2X1_LOC
XAND2X1_LOC_399 AND2X1_LOC_399/a_36_24# OR2X1_LOC_403/B AND2X1_LOC_399/a_8_24# VSS VDD
+ AND2X1_LOC_44/Y OR2X1_LOC_398/Y AND2X1_LOC
XAND2X1_LOC_333 AND2X1_LOC_333/a_36_24# AND2X1_LOC_338/A AND2X1_LOC_333/a_8_24# VSS VDD
+ OR2X1_LOC_171/Y OR2X1_LOC_289/Y AND2X1_LOC
XAND2X1_LOC_322 AND2X1_LOC_322/a_36_24# OR2X1_LOC_325/B AND2X1_LOC_322/a_8_24# VSS VDD
+ AND2X1_LOC_44/Y OR2X1_LOC_502/A AND2X1_LOC
XAND2X1_LOC_311 AND2X1_LOC_311/a_36_24# OR2X1_LOC_538/A AND2X1_LOC_311/a_8_24# VSS VDD
+ OR2X1_LOC_66/A OR2X1_LOC_532/B AND2X1_LOC
XAND2X1_LOC_377 AND2X1_LOC_377/a_36_24# AND2X1_LOC_377/Y AND2X1_LOC_377/a_8_24# VSS VDD
+ AND2X1_LOC_3/Y OR2X1_LOC_46/A AND2X1_LOC
XAND2X1_LOC_388 AND2X1_LOC_388/a_36_24# AND2X1_LOC_388/Y AND2X1_LOC_388/a_8_24# VSS VDD
+ OR2X1_LOC_167/Y OR2X1_LOC_176/Y AND2X1_LOC
XAND2X1_LOC_355 AND2X1_LOC_355/a_36_24# AND2X1_LOC_356/B AND2X1_LOC_355/a_8_24# VSS VDD
+ OR2X1_LOC_329/Y OR2X1_LOC_331/Y AND2X1_LOC
XOR2X1_LOC_119 OR2X1_LOC_119/a_8_216# OR2X1_LOC_119/a_36_216# OR2X1_LOC_426/B VSS VDD
+ OR2X1_LOC_46/A D_INPUT_1 OR2X1_LOC
XOR2X1_LOC_108 OR2X1_LOC_108/a_8_216# OR2X1_LOC_108/a_36_216# OR2X1_LOC_108/Y VSS VDD
+ OR2X1_LOC_485/A OR2X1_LOC_59/Y OR2X1_LOC
XAND2X1_LOC_73 AND2X1_LOC_73/a_36_24# OR2X1_LOC_185/A AND2X1_LOC_73/a_8_24# VSS VDD
+ OR2X1_LOC_62/B AND2X1_LOC_42/B AND2X1_LOC
XAND2X1_LOC_62 AND2X1_LOC_62/a_36_24# OR2X1_LOC_235/B AND2X1_LOC_62/a_8_24# VSS VDD
+ OR2X1_LOC_9/Y OR2X1_LOC_54/Y AND2X1_LOC
XAND2X1_LOC_84 AND2X1_LOC_84/a_36_24# AND2X1_LOC_84/Y AND2X1_LOC_84/a_8_24# VSS VDD
+ OR2X1_LOC_81/Y OR2X1_LOC_83/Y AND2X1_LOC
XAND2X1_LOC_40 AND2X1_LOC_40/a_36_24# AND2X1_LOC_40/Y AND2X1_LOC_40/a_8_24# VSS VDD
+ AND2X1_LOC_2/Y AND2X1_LOC_25/Y AND2X1_LOC
XAND2X1_LOC_95 AND2X1_LOC_95/a_36_24# AND2X1_LOC_95/Y AND2X1_LOC_95/a_8_24# VSS VDD
+ AND2X1_LOC_11/Y AND2X1_LOC_50/Y AND2X1_LOC
XAND2X1_LOC_51 AND2X1_LOC_51/a_36_24# AND2X1_LOC_51/Y AND2X1_LOC_51/a_8_24# VSS VDD
+ AND2X1_LOC_51/A AND2X1_LOC_50/Y AND2X1_LOC
XOR2X1_LOC_631 OR2X1_LOC_631/a_8_216# OR2X1_LOC_631/a_36_216# OR2X1_LOC_632/A VSS VDD
+ OR2X1_LOC_631/A OR2X1_LOC_631/B OR2X1_LOC
XOR2X1_LOC_642 OR2X1_LOC_642/a_8_216# OR2X1_LOC_642/a_36_216# OR2X1_LOC_649/B VSS VDD
+ OR2X1_LOC_520/Y OR2X1_LOC_462/B OR2X1_LOC
XOR2X1_LOC_653 OR2X1_LOC_653/a_8_216# OR2X1_LOC_653/a_36_216# OR2X1_LOC_653/Y VSS VDD
+ OR2X1_LOC_653/A OR2X1_LOC_653/B OR2X1_LOC
XOR2X1_LOC_620 OR2X1_LOC_620/a_8_216# OR2X1_LOC_620/a_36_216# OR2X1_LOC_620/Y VSS VDD
+ OR2X1_LOC_620/A OR2X1_LOC_620/B OR2X1_LOC
XOR2X1_LOC_686 OR2X1_LOC_686/a_8_216# OR2X1_LOC_686/a_36_216# OR2X1_LOC_687/A VSS VDD
+ OR2X1_LOC_686/A OR2X1_LOC_686/B OR2X1_LOC
XOR2X1_LOC_697 OR2X1_LOC_697/a_8_216# OR2X1_LOC_697/a_36_216# OR2X1_LOC_697/Y VSS VDD
+ OR2X1_LOC_428/A OR2X1_LOC_158/A OR2X1_LOC
XOR2X1_LOC_664 OR2X1_LOC_664/a_8_216# OR2X1_LOC_664/a_36_216# OR2X1_LOC_664/Y VSS VDD
+ OR2X1_LOC_78/A OR2X1_LOC_185/A OR2X1_LOC
XOR2X1_LOC_675 OR2X1_LOC_675/a_8_216# OR2X1_LOC_675/a_36_216# OR2X1_LOC_675/Y VSS VDD
+ OR2X1_LOC_675/A OR2X1_LOC_440/A OR2X1_LOC
XAND2X1_LOC_130 AND2X1_LOC_130/a_36_24# OR2X1_LOC_131/A AND2X1_LOC_130/a_8_24# VSS VDD
+ OR2X1_LOC_7/A OR2X1_LOC_589/A AND2X1_LOC
XAND2X1_LOC_141 AND2X1_LOC_141/a_36_24# AND2X1_LOC_657/A AND2X1_LOC_141/a_8_24# VSS VDD
+ AND2X1_LOC_141/A AND2X1_LOC_141/B AND2X1_LOC
XAND2X1_LOC_185 AND2X1_LOC_185/a_36_24# OR2X1_LOC_816/A AND2X1_LOC_185/a_8_24# VSS VDD
+ OR2X1_LOC_56/A OR2X1_LOC_74/A AND2X1_LOC
XAND2X1_LOC_174 AND2X1_LOC_174/a_36_24# AND2X1_LOC_175/B AND2X1_LOC_174/a_8_24# VSS VDD
+ OR2X1_LOC_171/Y OR2X1_LOC_172/Y AND2X1_LOC
XAND2X1_LOC_152 AND2X1_LOC_152/a_36_24# OR2X1_LOC_209/A AND2X1_LOC_152/a_8_24# VSS VDD
+ AND2X1_LOC_47/Y OR2X1_LOC_151/Y AND2X1_LOC
XAND2X1_LOC_196 AND2X1_LOC_196/a_36_24# AND2X1_LOC_196/Y AND2X1_LOC_196/a_8_24# VSS VDD
+ OR2X1_LOC_45/Y OR2X1_LOC_48/Y AND2X1_LOC
XAND2X1_LOC_163 AND2X1_LOC_163/a_36_24# OR2X1_LOC_467/B AND2X1_LOC_163/a_8_24# VSS VDD
+ AND2X1_LOC_51/Y OR2X1_LOC_162/Y AND2X1_LOC
XOR2X1_LOC_450 OR2X1_LOC_450/a_8_216# OR2X1_LOC_450/a_36_216# OR2X1_LOC_450/Y VSS VDD
+ OR2X1_LOC_450/A OR2X1_LOC_450/B OR2X1_LOC
XOR2X1_LOC_494 OR2X1_LOC_494/a_8_216# OR2X1_LOC_494/a_36_216# OR2X1_LOC_494/Y VSS VDD
+ OR2X1_LOC_494/A OR2X1_LOC_12/Y OR2X1_LOC
XOR2X1_LOC_483 OR2X1_LOC_483/a_8_216# OR2X1_LOC_483/a_36_216# OR2X1_LOC_631/B VSS VDD
+ OR2X1_LOC_833/B OR2X1_LOC_254/B OR2X1_LOC
XOR2X1_LOC_472 OR2X1_LOC_472/a_8_216# OR2X1_LOC_472/a_36_216# OR2X1_LOC_476/B VSS VDD
+ OR2X1_LOC_472/A OR2X1_LOC_472/B OR2X1_LOC
XOR2X1_LOC_461 OR2X1_LOC_461/a_8_216# OR2X1_LOC_461/a_36_216# OR2X1_LOC_461/Y VSS VDD
+ OR2X1_LOC_461/A OR2X1_LOC_461/B OR2X1_LOC
XOR2X1_LOC_291 OR2X1_LOC_291/a_8_216# OR2X1_LOC_291/a_36_216# OR2X1_LOC_291/Y VSS VDD
+ OR2X1_LOC_291/A OR2X1_LOC_36/Y OR2X1_LOC
XOR2X1_LOC_280 OR2X1_LOC_280/a_8_216# OR2X1_LOC_280/a_36_216# OR2X1_LOC_280/Y VSS VDD
+ OR2X1_LOC_428/A OR2X1_LOC_47/Y OR2X1_LOC
XAND2X1_LOC_729 AND2X1_LOC_729/a_36_24# AND2X1_LOC_729/Y AND2X1_LOC_729/a_8_24# VSS VDD
+ AND2X1_LOC_687/Y AND2X1_LOC_729/B AND2X1_LOC
XAND2X1_LOC_707 AND2X1_LOC_707/a_36_24# AND2X1_LOC_707/Y AND2X1_LOC_707/a_8_24# VSS VDD
+ OR2X1_LOC_694/Y OR2X1_LOC_695/Y AND2X1_LOC
XAND2X1_LOC_718 AND2X1_LOC_718/a_36_24# AND2X1_LOC_722/A AND2X1_LOC_718/a_8_24# VSS VDD
+ OR2X1_LOC_591/Y AND2X1_LOC_605/Y AND2X1_LOC
XAND2X1_LOC_504 AND2X1_LOC_504/a_36_24# OR2X1_LOC_507/B AND2X1_LOC_504/a_8_24# VSS VDD
+ AND2X1_LOC_41/A OR2X1_LOC_375/A AND2X1_LOC
XAND2X1_LOC_559 AND2X1_LOC_559/a_36_24# AND2X1_LOC_560/B AND2X1_LOC_559/a_8_24# VSS VDD
+ OR2X1_LOC_517/Y AND2X1_LOC_520/Y AND2X1_LOC
XAND2X1_LOC_548 AND2X1_LOC_548/a_36_24# AND2X1_LOC_548/Y AND2X1_LOC_548/a_8_24# VSS VDD
+ OR2X1_LOC_529/Y OR2X1_LOC_530/Y AND2X1_LOC
XAND2X1_LOC_515 AND2X1_LOC_515/a_36_24# OR2X1_LOC_516/A AND2X1_LOC_515/a_8_24# VSS VDD
+ OR2X1_LOC_417/Y AND2X1_LOC_514/Y AND2X1_LOC
XAND2X1_LOC_537 AND2X1_LOC_537/a_36_24# AND2X1_LOC_537/Y AND2X1_LOC_537/a_8_24# VSS VDD
+ OR2X1_LOC_385/Y OR2X1_LOC_536/Y AND2X1_LOC
XAND2X1_LOC_526 AND2X1_LOC_526/a_36_24# OR2X1_LOC_546/A AND2X1_LOC_526/a_8_24# VSS VDD
+ AND2X1_LOC_31/Y OR2X1_LOC_161/A AND2X1_LOC
XOR2X1_LOC_846 OR2X1_LOC_846/a_8_216# OR2X1_LOC_846/a_36_216# OR2X1_LOC_848/B VSS VDD
+ OR2X1_LOC_846/A OR2X1_LOC_846/B OR2X1_LOC
XOR2X1_LOC_824 OR2X1_LOC_824/a_8_216# OR2X1_LOC_824/a_36_216# OR2X1_LOC_824/Y VSS VDD
+ OR2X1_LOC_291/A OR2X1_LOC_26/Y OR2X1_LOC
XOR2X1_LOC_813 OR2X1_LOC_813/a_8_216# OR2X1_LOC_813/a_36_216# OR2X1_LOC_813/Y VSS VDD
+ OR2X1_LOC_813/A OR2X1_LOC_235/B OR2X1_LOC
XOR2X1_LOC_802 OR2X1_LOC_802/a_8_216# OR2X1_LOC_802/a_36_216# OR2X1_LOC_802/Y VSS VDD
+ OR2X1_LOC_802/A OR2X1_LOC_798/Y OR2X1_LOC
XOR2X1_LOC_835 OR2X1_LOC_835/a_8_216# OR2X1_LOC_835/a_36_216# OR2X1_LOC_835/Y VSS VDD
+ OR2X1_LOC_835/A OR2X1_LOC_835/B OR2X1_LOC
XOR2X1_LOC_857 OR2X1_LOC_857/a_8_216# OR2X1_LOC_857/a_36_216# OR2X1_LOC_863/A VSS VDD
+ OR2X1_LOC_857/A OR2X1_LOC_857/B OR2X1_LOC
XAND2X1_LOC_301 AND2X1_LOC_301/a_36_24# AND2X1_LOC_303/A AND2X1_LOC_301/a_8_24# VSS VDD
+ OR2X1_LOC_75/Y OR2X1_LOC_300/Y AND2X1_LOC
XAND2X1_LOC_312 AND2X1_LOC_312/a_36_24# OR2X1_LOC_703/A AND2X1_LOC_312/a_8_24# VSS VDD
+ AND2X1_LOC_56/B AND2X1_LOC_64/Y AND2X1_LOC
XOR2X1_LOC_109 OR2X1_LOC_109/a_8_216# OR2X1_LOC_109/a_36_216# OR2X1_LOC_109/Y VSS VDD
+ OR2X1_LOC_89/A OR2X1_LOC_31/Y OR2X1_LOC
XAND2X1_LOC_367 AND2X1_LOC_367/a_36_24# GATE_366 AND2X1_LOC_367/a_8_24# VSS VDD
+ AND2X1_LOC_367/A AND2X1_LOC_367/B AND2X1_LOC
XAND2X1_LOC_345 AND2X1_LOC_345/a_36_24# AND2X1_LOC_345/Y AND2X1_LOC_345/a_8_24# VSS VDD
+ AND2X1_LOC_259/Y OR2X1_LOC_261/Y AND2X1_LOC
XAND2X1_LOC_334 AND2X1_LOC_334/a_36_24# AND2X1_LOC_334/Y AND2X1_LOC_334/a_8_24# VSS VDD
+ OR2X1_LOC_290/Y OR2X1_LOC_291/Y AND2X1_LOC
XAND2X1_LOC_323 AND2X1_LOC_323/a_36_24# OR2X1_LOC_325/A AND2X1_LOC_323/a_8_24# VSS VDD
+ AND2X1_LOC_95/Y AND2X1_LOC_110/Y AND2X1_LOC
XAND2X1_LOC_378 AND2X1_LOC_378/a_36_24# OR2X1_LOC_459/A AND2X1_LOC_378/a_8_24# VSS VDD
+ OR2X1_LOC_43/A AND2X1_LOC_377/Y AND2X1_LOC
XAND2X1_LOC_356 AND2X1_LOC_356/a_36_24# AND2X1_LOC_365/A AND2X1_LOC_356/a_8_24# VSS VDD
+ AND2X1_LOC_354/Y AND2X1_LOC_356/B AND2X1_LOC
XAND2X1_LOC_389 AND2X1_LOC_389/a_36_24# AND2X1_LOC_390/B AND2X1_LOC_389/a_8_24# VSS VDD
+ OR2X1_LOC_385/Y OR2X1_LOC_387/Y AND2X1_LOC
XAND2X1_LOC_41 AND2X1_LOC_41/a_36_24# AND2X1_LOC_41/Y AND2X1_LOC_41/a_8_24# VSS VDD
+ AND2X1_LOC_41/A AND2X1_LOC_40/Y AND2X1_LOC
XAND2X1_LOC_52 AND2X1_LOC_52/a_36_24# AND2X1_LOC_52/Y AND2X1_LOC_52/a_8_24# VSS VDD
+ OR2X1_LOC_87/A AND2X1_LOC_51/Y AND2X1_LOC
XAND2X1_LOC_30 AND2X1_LOC_30/a_36_24# AND2X1_LOC_51/A AND2X1_LOC_30/a_8_24# VSS VDD
+ INPUT_4 INPUT_5 AND2X1_LOC
XOR2X1_LOC_687 OR2X1_LOC_687/a_8_216# OR2X1_LOC_687/a_36_216# OR2X1_LOC_687/Y VSS VDD
+ OR2X1_LOC_687/A OR2X1_LOC_687/B OR2X1_LOC
XOR2X1_LOC_676 OR2X1_LOC_676/a_8_216# OR2X1_LOC_676/a_36_216# OR2X1_LOC_676/Y VSS VDD
+ OR2X1_LOC_598/Y OR2X1_LOC_161/B OR2X1_LOC
XAND2X1_LOC_96 AND2X1_LOC_96/a_36_24# OR2X1_LOC_98/A AND2X1_LOC_96/a_8_24# VSS VDD
+ AND2X1_LOC_94/Y AND2X1_LOC_95/Y AND2X1_LOC
XAND2X1_LOC_74 AND2X1_LOC_74/a_36_24# OR2X1_LOC_76/B AND2X1_LOC_74/a_8_24# VSS VDD
+ AND2X1_LOC_31/Y OR2X1_LOC_185/A AND2X1_LOC
XAND2X1_LOC_63 AND2X1_LOC_63/a_36_24# AND2X1_LOC_65/A AND2X1_LOC_63/a_8_24# VSS VDD
+ AND2X1_LOC_8/Y OR2X1_LOC_235/B AND2X1_LOC
XAND2X1_LOC_85 AND2X1_LOC_85/a_36_24# AND2X1_LOC_86/B AND2X1_LOC_85/a_8_24# VSS VDD
+ AND2X1_LOC_18/Y AND2X1_LOC_42/B AND2X1_LOC
XOR2X1_LOC_665 OR2X1_LOC_665/a_8_216# OR2X1_LOC_665/a_36_216# OR2X1_LOC_665/Y VSS VDD
+ OR2X1_LOC_755/A OR2X1_LOC_3/Y OR2X1_LOC
XOR2X1_LOC_621 OR2X1_LOC_621/a_8_216# OR2X1_LOC_621/a_36_216# OR2X1_LOC_622/A VSS VDD
+ OR2X1_LOC_621/A OR2X1_LOC_621/B OR2X1_LOC
XOR2X1_LOC_632 OR2X1_LOC_632/a_8_216# OR2X1_LOC_632/a_36_216# OR2X1_LOC_632/Y VSS VDD
+ OR2X1_LOC_632/A OR2X1_LOC_630/Y OR2X1_LOC
XOR2X1_LOC_610 OR2X1_LOC_610/a_8_216# OR2X1_LOC_610/a_36_216# OR2X1_LOC_610/Y VSS VDD
+ AND2X1_LOC_47/Y AND2X1_LOC_40/Y OR2X1_LOC
XOR2X1_LOC_643 OR2X1_LOC_643/a_8_216# OR2X1_LOC_643/a_36_216# OR2X1_LOC_643/Y VSS VDD
+ OR2X1_LOC_643/A OR2X1_LOC_539/B OR2X1_LOC
XOR2X1_LOC_654 OR2X1_LOC_654/a_8_216# OR2X1_LOC_654/a_36_216# OR2X1_LOC_661/A VSS VDD
+ OR2X1_LOC_654/A OR2X1_LOC_650/Y OR2X1_LOC
XOR2X1_LOC_698 OR2X1_LOC_698/a_8_216# OR2X1_LOC_698/a_36_216# OR2X1_LOC_698/Y VSS VDD
+ OR2X1_LOC_744/A OR2X1_LOC_64/Y OR2X1_LOC
XAND2X1_LOC_153 AND2X1_LOC_153/a_36_24# OR2X1_LOC_155/A AND2X1_LOC_153/a_8_24# VSS VDD
+ D_INPUT_1 AND2X1_LOC_42/B AND2X1_LOC
XAND2X1_LOC_120 AND2X1_LOC_120/a_36_24# OR2X1_LOC_666/A AND2X1_LOC_120/a_8_24# VSS VDD
+ OR2X1_LOC_13/B OR2X1_LOC_39/A AND2X1_LOC
XAND2X1_LOC_131 AND2X1_LOC_131/a_36_24# OR2X1_LOC_140/A AND2X1_LOC_131/a_8_24# VSS VDD
+ AND2X1_LOC_12/Y OR2X1_LOC_130/Y AND2X1_LOC
XAND2X1_LOC_164 AND2X1_LOC_164/a_36_24# OR2X1_LOC_168/B AND2X1_LOC_164/a_8_24# VSS VDD
+ AND2X1_LOC_18/Y OR2X1_LOC_502/A AND2X1_LOC
XAND2X1_LOC_142 AND2X1_LOC_142/a_36_24# OR2X1_LOC_147/B AND2X1_LOC_142/a_8_24# VSS VDD
+ OR2X1_LOC_87/A AND2X1_LOC_64/Y AND2X1_LOC
XAND2X1_LOC_186 AND2X1_LOC_186/a_36_24# OR2X1_LOC_680/A AND2X1_LOC_186/a_8_24# VSS VDD
+ OR2X1_LOC_437/A OR2X1_LOC_816/A AND2X1_LOC
XAND2X1_LOC_175 AND2X1_LOC_175/a_36_24# AND2X1_LOC_211/B AND2X1_LOC_175/a_8_24# VSS VDD
+ OR2X1_LOC_173/Y AND2X1_LOC_175/B AND2X1_LOC
XAND2X1_LOC_197 AND2X1_LOC_197/a_36_24# AND2X1_LOC_197/Y AND2X1_LOC_197/a_8_24# VSS VDD
+ OR2X1_LOC_52/Y OR2X1_LOC_56/Y AND2X1_LOC
XOR2X1_LOC_451 OR2X1_LOC_451/a_8_216# OR2X1_LOC_451/a_36_216# OR2X1_LOC_452/A VSS VDD
+ OR2X1_LOC_451/A OR2X1_LOC_451/B OR2X1_LOC
XOR2X1_LOC_484 OR2X1_LOC_484/a_8_216# OR2X1_LOC_484/a_36_216# OR2X1_LOC_484/Y VSS VDD
+ OR2X1_LOC_36/Y OR2X1_LOC_13/B OR2X1_LOC
XOR2X1_LOC_473 OR2X1_LOC_473/a_8_216# OR2X1_LOC_473/a_36_216# OR2X1_LOC_473/Y VSS VDD
+ OR2X1_LOC_473/A OR2X1_LOC_216/A OR2X1_LOC
XOR2X1_LOC_495 OR2X1_LOC_495/a_8_216# OR2X1_LOC_495/a_36_216# OR2X1_LOC_495/Y VSS VDD
+ OR2X1_LOC_56/A OR2X1_LOC_36/Y OR2X1_LOC
XOR2X1_LOC_462 OR2X1_LOC_462/a_8_216# OR2X1_LOC_462/a_36_216# OR2X1_LOC_472/B VSS VDD
+ OR2X1_LOC_461/Y OR2X1_LOC_462/B OR2X1_LOC
XOR2X1_LOC_440 OR2X1_LOC_440/a_8_216# OR2X1_LOC_440/a_36_216# OR2X1_LOC_468/A VSS VDD
+ OR2X1_LOC_440/A OR2X1_LOC_440/B OR2X1_LOC
XOR2X1_LOC_292 OR2X1_LOC_292/a_8_216# OR2X1_LOC_292/a_36_216# OR2X1_LOC_292/Y VSS VDD
+ OR2X1_LOC_437/A OR2X1_LOC_40/Y OR2X1_LOC
XOR2X1_LOC_281 OR2X1_LOC_281/a_8_216# OR2X1_LOC_281/a_36_216# OR2X1_LOC_281/Y VSS VDD
+ OR2X1_LOC_428/A OR2X1_LOC_3/Y OR2X1_LOC
XOR2X1_LOC_270 OR2X1_LOC_270/a_8_216# OR2X1_LOC_270/a_36_216# OR2X1_LOC_270/Y VSS VDD
+ AND2X1_LOC_36/Y AND2X1_LOC_18/Y OR2X1_LOC
XAND2X1_LOC_719 AND2X1_LOC_719/a_36_24# AND2X1_LOC_719/Y AND2X1_LOC_719/a_8_24# VSS VDD
+ OR2X1_LOC_665/Y OR2X1_LOC_666/Y AND2X1_LOC
XAND2X1_LOC_708 AND2X1_LOC_708/a_36_24# AND2X1_LOC_712/B AND2X1_LOC_708/a_8_24# VSS VDD
+ OR2X1_LOC_696/Y OR2X1_LOC_697/Y AND2X1_LOC
XAND2X1_LOC_505 AND2X1_LOC_505/a_36_24# OR2X1_LOC_507/A AND2X1_LOC_505/a_8_24# VSS VDD
+ AND2X1_LOC_18/Y OR2X1_LOC_160/B AND2X1_LOC
XAND2X1_LOC_549 AND2X1_LOC_549/a_36_24# AND2X1_LOC_549/Y AND2X1_LOC_549/a_8_24# VSS VDD
+ OR2X1_LOC_531/Y AND2X1_LOC_548/Y AND2X1_LOC
XAND2X1_LOC_527 AND2X1_LOC_527/a_36_24# OR2X1_LOC_547/B AND2X1_LOC_527/a_8_24# VSS VDD
+ AND2X1_LOC_64/Y AND2X1_LOC_110/Y AND2X1_LOC
XAND2X1_LOC_516 AND2X1_LOC_516/a_36_24# OR2X1_LOC_574/A AND2X1_LOC_516/a_8_24# VSS VDD
+ OR2X1_LOC_513/Y OR2X1_LOC_515/Y AND2X1_LOC
XAND2X1_LOC_538 AND2X1_LOC_538/a_36_24# AND2X1_LOC_538/Y AND2X1_LOC_538/a_8_24# VSS VDD
+ OR2X1_LOC_13/Y OR2X1_LOC_311/Y AND2X1_LOC
XOR2X1_LOC_803 OR2X1_LOC_803/a_8_216# OR2X1_LOC_803/a_36_216# OR2X1_LOC_808/B VSS VDD
+ OR2X1_LOC_803/A OR2X1_LOC_803/B OR2X1_LOC
XOR2X1_LOC_847 OR2X1_LOC_847/a_8_216# OR2X1_LOC_847/a_36_216# OR2X1_LOC_848/A VSS VDD
+ OR2X1_LOC_847/A OR2X1_LOC_847/B OR2X1_LOC
XOR2X1_LOC_825 OR2X1_LOC_825/a_8_216# OR2X1_LOC_825/a_36_216# OR2X1_LOC_825/Y VSS VDD
+ OR2X1_LOC_96/B OR2X1_LOC_44/Y OR2X1_LOC
XOR2X1_LOC_858 OR2X1_LOC_858/a_8_216# OR2X1_LOC_858/a_36_216# OR2X1_LOC_862/B VSS VDD
+ OR2X1_LOC_858/A OR2X1_LOC_858/B OR2X1_LOC
XOR2X1_LOC_814 OR2X1_LOC_814/a_8_216# OR2X1_LOC_814/a_36_216# OR2X1_LOC_814/Y VSS VDD
+ OR2X1_LOC_814/A OR2X1_LOC_756/B OR2X1_LOC
XOR2X1_LOC_836 OR2X1_LOC_836/a_8_216# OR2X1_LOC_836/a_36_216# OR2X1_LOC_836/Y VSS VDD
+ OR2X1_LOC_836/A OR2X1_LOC_836/B OR2X1_LOC
XAND2X1_LOC_346 AND2X1_LOC_346/a_36_24# AND2X1_LOC_347/B AND2X1_LOC_346/a_8_24# VSS VDD
+ OR2X1_LOC_292/Y OR2X1_LOC_295/Y AND2X1_LOC
XAND2X1_LOC_335 AND2X1_LOC_335/a_36_24# AND2X1_LOC_335/Y AND2X1_LOC_335/a_8_24# VSS VDD
+ OR2X1_LOC_309/Y OR2X1_LOC_310/Y AND2X1_LOC
XAND2X1_LOC_302 AND2X1_LOC_302/a_36_24# AND2X1_LOC_303/B AND2X1_LOC_302/a_8_24# VSS VDD
+ OR2X1_LOC_298/Y OR2X1_LOC_299/Y AND2X1_LOC
XAND2X1_LOC_324 AND2X1_LOC_324/a_36_24# AND2X1_LOC_326/A AND2X1_LOC_324/a_8_24# VSS VDD
+ OR2X1_LOC_320/Y OR2X1_LOC_321/Y AND2X1_LOC
XAND2X1_LOC_313 AND2X1_LOC_313/a_36_24# OR2X1_LOC_317/B AND2X1_LOC_313/a_8_24# VSS VDD
+ AND2X1_LOC_70/Y AND2X1_LOC_91/B AND2X1_LOC
XAND2X1_LOC_368 AND2X1_LOC_368/a_36_24# OR2X1_LOC_457/B AND2X1_LOC_368/a_8_24# VSS VDD
+ AND2X1_LOC_7/B OR2X1_LOC_270/Y AND2X1_LOC
XAND2X1_LOC_357 AND2X1_LOC_357/a_36_24# AND2X1_LOC_364/A AND2X1_LOC_357/a_8_24# VSS VDD
+ AND2X1_LOC_357/A AND2X1_LOC_357/B AND2X1_LOC
XAND2X1_LOC_379 AND2X1_LOC_379/a_36_24# OR2X1_LOC_380/A AND2X1_LOC_379/a_8_24# VSS VDD
+ OR2X1_LOC_12/Y OR2X1_LOC_26/Y AND2X1_LOC
XAND2X1_LOC_42 AND2X1_LOC_42/a_36_24# AND2X1_LOC_43/B AND2X1_LOC_42/a_8_24# VSS VDD
+ INPUT_1 AND2X1_LOC_42/B AND2X1_LOC
XAND2X1_LOC_75 AND2X1_LOC_75/a_36_24# OR2X1_LOC_76/A AND2X1_LOC_75/a_8_24# VSS VDD
+ OR2X1_LOC_160/B AND2X1_LOC_59/Y AND2X1_LOC
XAND2X1_LOC_86 AND2X1_LOC_86/a_36_24# AND2X1_LOC_86/Y AND2X1_LOC_86/a_8_24# VSS VDD
+ INPUT_0 AND2X1_LOC_86/B AND2X1_LOC
XAND2X1_LOC_20 AND2X1_LOC_20/a_36_24# OR2X1_LOC_33/B AND2X1_LOC_20/a_8_24# VSS VDD
+ AND2X1_LOC_18/Y AND2X1_LOC_19/Y AND2X1_LOC
XAND2X1_LOC_53 AND2X1_LOC_53/a_36_24# AND2X1_LOC_53/Y AND2X1_LOC_53/a_8_24# VSS VDD
+ D_INPUT_5 AND2X1_LOC_50/Y AND2X1_LOC
XAND2X1_LOC_64 AND2X1_LOC_64/a_36_24# AND2X1_LOC_64/Y AND2X1_LOC_64/a_8_24# VSS VDD
+ AND2X1_LOC_21/Y AND2X1_LOC_50/Y AND2X1_LOC
XAND2X1_LOC_31 AND2X1_LOC_31/a_36_24# AND2X1_LOC_31/Y AND2X1_LOC_31/a_8_24# VSS VDD
+ AND2X1_LOC_1/Y AND2X1_LOC_51/A AND2X1_LOC
XOR2X1_LOC_600 OR2X1_LOC_600/a_8_216# OR2X1_LOC_600/a_36_216# OR2X1_LOC_600/Y VSS VDD
+ OR2X1_LOC_600/A OR2X1_LOC_31/Y OR2X1_LOC
XOR2X1_LOC_677 OR2X1_LOC_677/a_8_216# OR2X1_LOC_677/a_36_216# OR2X1_LOC_677/Y VSS VDD
+ OR2X1_LOC_427/A OR2X1_LOC_26/Y OR2X1_LOC
XAND2X1_LOC_97 AND2X1_LOC_97/a_36_24# AND2X1_LOC_99/A AND2X1_LOC_97/a_8_24# VSS VDD
+ OR2X1_LOC_89/Y OR2X1_LOC_91/Y AND2X1_LOC
XOR2X1_LOC_699 OR2X1_LOC_699/a_8_216# OR2X1_LOC_699/a_36_216# OR2X1_LOC_748/A VSS VDD
+ OR2X1_LOC_158/A OR2X1_LOC_46/A OR2X1_LOC
XOR2X1_LOC_622 OR2X1_LOC_622/a_8_216# OR2X1_LOC_622/a_36_216# OR2X1_LOC_624/B VSS VDD
+ OR2X1_LOC_622/A OR2X1_LOC_622/B OR2X1_LOC
XOR2X1_LOC_611 OR2X1_LOC_611/a_8_216# OR2X1_LOC_611/a_36_216# OR2X1_LOC_611/Y VSS VDD
+ OR2X1_LOC_62/A OR2X1_LOC_6/A OR2X1_LOC
XOR2X1_LOC_666 OR2X1_LOC_666/a_8_216# OR2X1_LOC_666/a_36_216# OR2X1_LOC_666/Y VSS VDD
+ OR2X1_LOC_666/A OR2X1_LOC_18/Y OR2X1_LOC
XOR2X1_LOC_633 OR2X1_LOC_633/a_8_216# OR2X1_LOC_633/a_36_216# OR2X1_LOC_633/Y VSS VDD
+ OR2X1_LOC_633/A OR2X1_LOC_633/B OR2X1_LOC
XOR2X1_LOC_655 OR2X1_LOC_655/a_8_216# OR2X1_LOC_655/a_36_216# OR2X1_LOC_660/B VSS VDD
+ OR2X1_LOC_655/A OR2X1_LOC_655/B OR2X1_LOC
XOR2X1_LOC_688 OR2X1_LOC_688/a_8_216# OR2X1_LOC_688/a_36_216# OR2X1_LOC_688/Y VSS VDD
+ OR2X1_LOC_598/A OR2X1_LOC_154/A OR2X1_LOC
XOR2X1_LOC_644 OR2X1_LOC_644/a_8_216# OR2X1_LOC_644/a_36_216# OR2X1_LOC_648/B VSS VDD
+ OR2X1_LOC_644/A OR2X1_LOC_644/B OR2X1_LOC
XAND2X1_LOC_121 AND2X1_LOC_121/a_36_24# OR2X1_LOC_122/A AND2X1_LOC_121/a_8_24# VSS VDD
+ OR2X1_LOC_426/B OR2X1_LOC_666/A AND2X1_LOC
XAND2X1_LOC_143 AND2X1_LOC_143/a_36_24# OR2X1_LOC_502/A AND2X1_LOC_143/a_8_24# VSS VDD
+ D_INPUT_1 AND2X1_LOC_8/Y AND2X1_LOC
XAND2X1_LOC_132 AND2X1_LOC_132/a_36_24# OR2X1_LOC_137/B AND2X1_LOC_132/a_8_24# VSS VDD
+ AND2X1_LOC_91/B AND2X1_LOC_95/Y AND2X1_LOC
XAND2X1_LOC_187 AND2X1_LOC_187/a_36_24# OR2X1_LOC_191/B AND2X1_LOC_187/a_8_24# VSS VDD
+ AND2X1_LOC_40/Y OR2X1_LOC_186/Y AND2X1_LOC
XAND2X1_LOC_176 AND2X1_LOC_176/a_36_24# OR2X1_LOC_180/B AND2X1_LOC_176/a_8_24# VSS VDD
+ OR2X1_LOC_66/A AND2X1_LOC_91/B AND2X1_LOC
XAND2X1_LOC_165 AND2X1_LOC_165/a_36_24# OR2X1_LOC_168/A AND2X1_LOC_165/a_8_24# VSS VDD
+ AND2X1_LOC_51/Y OR2X1_LOC_185/A AND2X1_LOC
XAND2X1_LOC_110 AND2X1_LOC_110/a_36_24# AND2X1_LOC_110/Y AND2X1_LOC_110/a_8_24# VSS VDD
+ D_INPUT_0 OR2X1_LOC_377/A AND2X1_LOC
XAND2X1_LOC_198 AND2X1_LOC_198/a_36_24# AND2X1_LOC_208/B AND2X1_LOC_198/a_8_24# VSS VDD
+ OR2X1_LOC_57/Y AND2X1_LOC_197/Y AND2X1_LOC
XAND2X1_LOC_154 AND2X1_LOC_154/a_36_24# AND2X1_LOC_154/Y AND2X1_LOC_154/a_8_24# VSS VDD
+ OR2X1_LOC_7/A OR2X1_LOC_39/A AND2X1_LOC
XOR2X1_LOC_430 OR2X1_LOC_430/a_8_216# OR2X1_LOC_430/a_36_216# OR2X1_LOC_430/Y VSS VDD
+ OR2X1_LOC_429/Y OR2X1_LOC_604/A OR2X1_LOC
XOR2X1_LOC_452 OR2X1_LOC_452/a_8_216# OR2X1_LOC_452/a_36_216# OR2X1_LOC_467/A VSS VDD
+ OR2X1_LOC_452/A OR2X1_LOC_450/Y OR2X1_LOC
XOR2X1_LOC_485 OR2X1_LOC_485/a_8_216# OR2X1_LOC_485/a_36_216# OR2X1_LOC_485/Y VSS VDD
+ OR2X1_LOC_485/A OR2X1_LOC_44/Y OR2X1_LOC
XOR2X1_LOC_463 OR2X1_LOC_463/a_8_216# OR2X1_LOC_463/a_36_216# OR2X1_LOC_472/A VSS VDD
+ OR2X1_LOC_460/Y OR2X1_LOC_463/B OR2X1_LOC
XOR2X1_LOC_474 OR2X1_LOC_474/a_8_216# OR2X1_LOC_474/a_36_216# OR2X1_LOC_474/Y VSS VDD
+ OR2X1_LOC_404/Y OR2X1_LOC_474/B OR2X1_LOC
XOR2X1_LOC_496 OR2X1_LOC_496/a_8_216# OR2X1_LOC_496/a_36_216# OR2X1_LOC_496/Y VSS VDD
+ OR2X1_LOC_56/A OR2X1_LOC_18/Y OR2X1_LOC
XOR2X1_LOC_441 OR2X1_LOC_441/a_8_216# OR2X1_LOC_441/a_36_216# OR2X1_LOC_441/Y VSS VDD
+ OR2X1_LOC_52/B OR2X1_LOC_40/Y OR2X1_LOC
XOR2X1_LOC_260 OR2X1_LOC_260/a_8_216# OR2X1_LOC_260/a_36_216# OR2X1_LOC_260/Y VSS VDD
+ OR2X1_LOC_375/A AND2X1_LOC_12/Y OR2X1_LOC
XOR2X1_LOC_271 OR2X1_LOC_271/a_8_216# OR2X1_LOC_271/a_36_216# OR2X1_LOC_271/Y VSS VDD
+ OR2X1_LOC_368/A OR2X1_LOC_271/B OR2X1_LOC
XOR2X1_LOC_282 OR2X1_LOC_282/a_8_216# OR2X1_LOC_282/a_36_216# OR2X1_LOC_282/Y VSS VDD
+ OR2X1_LOC_158/A OR2X1_LOC_485/A OR2X1_LOC
XOR2X1_LOC_293 OR2X1_LOC_293/a_8_216# OR2X1_LOC_293/a_36_216# OR2X1_LOC_585/A VSS VDD
+ OR2X1_LOC_6/A D_INPUT_1 OR2X1_LOC
XAND2X1_LOC_709 AND2X1_LOC_709/a_36_24# AND2X1_LOC_711/A AND2X1_LOC_709/a_8_24# VSS VDD
+ OR2X1_LOC_698/Y OR2X1_LOC_748/A AND2X1_LOC
XAND2X1_LOC_506 AND2X1_LOC_506/a_36_24# AND2X1_LOC_508/A AND2X1_LOC_506/a_8_24# VSS VDD
+ OR2X1_LOC_239/Y OR2X1_LOC_419/Y AND2X1_LOC
XAND2X1_LOC_517 AND2X1_LOC_517/a_36_24# OR2X1_LOC_559/B AND2X1_LOC_517/a_8_24# VSS VDD
+ AND2X1_LOC_31/Y OR2X1_LOC_264/Y AND2X1_LOC
XAND2X1_LOC_528 AND2X1_LOC_528/a_36_24# OR2X1_LOC_620/B AND2X1_LOC_528/a_8_24# VSS VDD
+ AND2X1_LOC_7/B AND2X1_LOC_44/Y AND2X1_LOC
XAND2X1_LOC_539 AND2X1_LOC_539/a_36_24# AND2X1_LOC_539/Y AND2X1_LOC_539/a_8_24# VSS VDD
+ AND2X1_LOC_537/Y AND2X1_LOC_538/Y AND2X1_LOC
XOR2X1_LOC_859 OR2X1_LOC_859/a_8_216# OR2X1_LOC_859/a_36_216# OR2X1_LOC_862/A VSS VDD
+ OR2X1_LOC_859/A OR2X1_LOC_859/B OR2X1_LOC
XOR2X1_LOC_848 OR2X1_LOC_848/a_8_216# OR2X1_LOC_848/a_36_216# OR2X1_LOC_859/B VSS VDD
+ OR2X1_LOC_848/A OR2X1_LOC_848/B OR2X1_LOC
XOR2X1_LOC_826 OR2X1_LOC_826/a_8_216# OR2X1_LOC_826/a_36_216# OR2X1_LOC_826/Y VSS VDD
+ OR2X1_LOC_95/Y OR2X1_LOC_56/A OR2X1_LOC
XOR2X1_LOC_815 OR2X1_LOC_815/a_8_216# OR2X1_LOC_815/a_36_216# OR2X1_LOC_815/Y VSS VDD
+ OR2X1_LOC_815/A OR2X1_LOC_3/Y OR2X1_LOC
XOR2X1_LOC_804 OR2X1_LOC_804/a_8_216# OR2X1_LOC_804/a_36_216# OR2X1_LOC_808/A VSS VDD
+ OR2X1_LOC_804/A OR2X1_LOC_804/B OR2X1_LOC
XOR2X1_LOC_837 OR2X1_LOC_837/a_8_216# OR2X1_LOC_837/a_36_216# OR2X1_LOC_837/Y VSS VDD
+ OR2X1_LOC_837/A OR2X1_LOC_837/B OR2X1_LOC
XAND2X1_LOC_369 AND2X1_LOC_369/a_36_24# OR2X1_LOC_543/A AND2X1_LOC_369/a_8_24# VSS VDD
+ AND2X1_LOC_22/Y OR2X1_LOC_121/B AND2X1_LOC
XAND2X1_LOC_347 AND2X1_LOC_347/a_36_24# AND2X1_LOC_347/Y AND2X1_LOC_347/a_8_24# VSS VDD
+ OR2X1_LOC_297/Y AND2X1_LOC_347/B AND2X1_LOC
XAND2X1_LOC_358 AND2X1_LOC_358/a_36_24# AND2X1_LOC_358/Y AND2X1_LOC_358/a_8_24# VSS VDD
+ AND2X1_LOC_350/Y AND2X1_LOC_351/Y AND2X1_LOC
XAND2X1_LOC_325 AND2X1_LOC_325/a_36_24# AND2X1_LOC_326/B AND2X1_LOC_325/a_8_24# VSS VDD
+ OR2X1_LOC_322/Y OR2X1_LOC_323/Y AND2X1_LOC
XAND2X1_LOC_303 AND2X1_LOC_303/a_36_24# AND2X1_LOC_566/B AND2X1_LOC_303/a_8_24# VSS VDD
+ AND2X1_LOC_303/A AND2X1_LOC_303/B AND2X1_LOC
XAND2X1_LOC_314 AND2X1_LOC_314/a_36_24# OR2X1_LOC_317/A AND2X1_LOC_314/a_8_24# VSS VDD
+ OR2X1_LOC_78/B AND2X1_LOC_64/Y AND2X1_LOC
XAND2X1_LOC_336 AND2X1_LOC_336/a_36_24# AND2X1_LOC_337/B AND2X1_LOC_336/a_8_24# VSS VDD
+ OR2X1_LOC_311/Y OR2X1_LOC_312/Y AND2X1_LOC
XOR2X1_LOC_601 OR2X1_LOC_601/a_8_216# OR2X1_LOC_601/a_36_216# OR2X1_LOC_601/Y VSS VDD
+ OR2X1_LOC_47/Y OR2X1_LOC_16/A OR2X1_LOC
XAND2X1_LOC_65 AND2X1_LOC_65/a_36_24# OR2X1_LOC_201/A AND2X1_LOC_65/a_8_24# VSS VDD
+ AND2X1_LOC_65/A AND2X1_LOC_64/Y AND2X1_LOC
XAND2X1_LOC_87 AND2X1_LOC_87/a_36_24# OR2X1_LOC_88/A AND2X1_LOC_87/a_8_24# VSS VDD
+ OR2X1_LOC_32/B OR2X1_LOC_52/B AND2X1_LOC
XAND2X1_LOC_10 AND2X1_LOC_10/a_36_24# AND2X1_LOC_41/A AND2X1_LOC_10/a_8_24# VSS VDD
+ AND2X1_LOC_8/Y OR2X1_LOC_62/B AND2X1_LOC
XAND2X1_LOC_98 AND2X1_LOC_98/a_36_24# AND2X1_LOC_98/Y AND2X1_LOC_98/a_8_24# VSS VDD
+ OR2X1_LOC_93/Y OR2X1_LOC_96/Y AND2X1_LOC
XAND2X1_LOC_54 AND2X1_LOC_54/a_36_24# OR2X1_LOC_62/A AND2X1_LOC_54/a_8_24# VSS VDD
+ INPUT_0 INPUT_1 AND2X1_LOC
XAND2X1_LOC_76 AND2X1_LOC_76/a_36_24# AND2X1_LOC_76/Y AND2X1_LOC_76/a_8_24# VSS VDD
+ OR2X1_LOC_74/Y OR2X1_LOC_75/Y AND2X1_LOC
XAND2X1_LOC_32 AND2X1_LOC_32/a_36_24# OR2X1_LOC_34/A AND2X1_LOC_32/a_8_24# VSS VDD
+ OR2X1_LOC_87/B AND2X1_LOC_31/Y AND2X1_LOC
XAND2X1_LOC_43 AND2X1_LOC_43/a_36_24# OR2X1_LOC_195/A AND2X1_LOC_43/a_8_24# VSS VDD
+ AND2X1_LOC_22/Y AND2X1_LOC_43/B AND2X1_LOC
XAND2X1_LOC_21 AND2X1_LOC_21/a_36_24# AND2X1_LOC_21/Y AND2X1_LOC_21/a_8_24# VSS VDD
+ INPUT_4 D_INPUT_5 AND2X1_LOC
XOR2X1_LOC_612 OR2X1_LOC_612/a_8_216# OR2X1_LOC_612/a_36_216# OR2X1_LOC_612/Y VSS VDD
+ OR2X1_LOC_611/Y OR2X1_LOC_612/B OR2X1_LOC
XOR2X1_LOC_678 OR2X1_LOC_678/a_8_216# OR2X1_LOC_678/a_36_216# OR2X1_LOC_678/Y VSS VDD
+ OR2X1_LOC_834/A AND2X1_LOC_12/Y OR2X1_LOC
XOR2X1_LOC_689 OR2X1_LOC_689/a_8_216# OR2X1_LOC_689/a_36_216# OR2X1_LOC_689/Y VSS VDD
+ OR2X1_LOC_689/A OR2X1_LOC_31/Y OR2X1_LOC
XOR2X1_LOC_667 OR2X1_LOC_667/a_8_216# OR2X1_LOC_667/a_36_216# OR2X1_LOC_667/Y VSS VDD
+ OR2X1_LOC_517/A OR2X1_LOC_64/Y OR2X1_LOC
XOR2X1_LOC_656 OR2X1_LOC_656/a_8_216# OR2X1_LOC_656/a_36_216# OR2X1_LOC_656/Y VSS VDD
+ OR2X1_LOC_647/Y OR2X1_LOC_656/B OR2X1_LOC
XOR2X1_LOC_645 OR2X1_LOC_645/a_8_216# OR2X1_LOC_645/a_36_216# OR2X1_LOC_648/A VSS VDD
+ OR2X1_LOC_605/Y OR2X1_LOC_602/Y OR2X1_LOC
XOR2X1_LOC_634 OR2X1_LOC_634/a_8_216# OR2X1_LOC_634/a_36_216# OR2X1_LOC_640/A VSS VDD
+ OR2X1_LOC_634/A OR2X1_LOC_334/B OR2X1_LOC
XOR2X1_LOC_623 OR2X1_LOC_623/a_8_216# OR2X1_LOC_623/a_36_216# OR2X1_LOC_624/A VSS VDD
+ OR2X1_LOC_620/Y OR2X1_LOC_623/B OR2X1_LOC
XAND2X1_LOC_100 AND2X1_LOC_100/a_36_24# AND2X1_LOC_101/B AND2X1_LOC_100/a_8_24# VSS VDD
+ OR2X1_LOC_86/Y OR2X1_LOC_88/Y AND2X1_LOC
XAND2X1_LOC_122 AND2X1_LOC_122/a_36_24# OR2X1_LOC_124/B AND2X1_LOC_122/a_8_24# VSS VDD
+ AND2X1_LOC_44/Y OR2X1_LOC_121/Y AND2X1_LOC
XAND2X1_LOC_133 AND2X1_LOC_133/a_36_24# OR2X1_LOC_161/B AND2X1_LOC_133/a_8_24# VSS VDD
+ AND2X1_LOC_8/Y OR2X1_LOC_80/A AND2X1_LOC
XAND2X1_LOC_188 AND2X1_LOC_188/a_36_24# OR2X1_LOC_189/A AND2X1_LOC_188/a_8_24# VSS VDD
+ OR2X1_LOC_39/A OR2X1_LOC_816/A AND2X1_LOC
XAND2X1_LOC_177 AND2X1_LOC_177/a_36_24# OR2X1_LOC_439/B AND2X1_LOC_177/a_8_24# VSS VDD
+ OR2X1_LOC_87/A AND2X1_LOC_70/Y AND2X1_LOC
XAND2X1_LOC_166 AND2X1_LOC_166/a_36_24# OR2X1_LOC_169/B AND2X1_LOC_166/a_8_24# VSS VDD
+ OR2X1_LOC_78/B AND2X1_LOC_40/Y AND2X1_LOC
XAND2X1_LOC_111 AND2X1_LOC_111/a_36_24# OR2X1_LOC_112/A AND2X1_LOC_111/a_8_24# VSS VDD
+ AND2X1_LOC_31/Y AND2X1_LOC_110/Y AND2X1_LOC
XAND2X1_LOC_199 AND2X1_LOC_199/a_36_24# AND2X1_LOC_207/A AND2X1_LOC_199/a_8_24# VSS VDD
+ AND2X1_LOC_199/A AND2X1_LOC_196/Y AND2X1_LOC
XAND2X1_LOC_144 AND2X1_LOC_144/a_36_24# OR2X1_LOC_147/A AND2X1_LOC_144/a_8_24# VSS VDD
+ AND2X1_LOC_59/Y OR2X1_LOC_502/A AND2X1_LOC
XAND2X1_LOC_155 AND2X1_LOC_155/a_36_24# AND2X1_LOC_155/Y AND2X1_LOC_155/a_8_24# VSS VDD
+ OR2X1_LOC_52/B OR2X1_LOC_743/A AND2X1_LOC
XOR2X1_LOC_453 OR2X1_LOC_453/a_8_216# OR2X1_LOC_453/a_36_216# OR2X1_LOC_453/Y VSS VDD
+ OR2X1_LOC_453/A OR2X1_LOC_448/Y OR2X1_LOC
XOR2X1_LOC_420 OR2X1_LOC_420/a_8_216# OR2X1_LOC_420/a_36_216# OR2X1_LOC_420/Y VSS VDD
+ OR2X1_LOC_485/A OR2X1_LOC_95/Y OR2X1_LOC
XOR2X1_LOC_431 OR2X1_LOC_431/a_8_216# OR2X1_LOC_431/a_36_216# OR2X1_LOC_431/Y VSS VDD
+ OR2X1_LOC_428/A OR2X1_LOC_70/Y OR2X1_LOC
XOR2X1_LOC_442 OR2X1_LOC_442/a_8_216# OR2X1_LOC_442/a_36_216# OR2X1_LOC_442/Y VSS VDD
+ OR2X1_LOC_600/A OR2X1_LOC_40/Y OR2X1_LOC
XOR2X1_LOC_464 OR2X1_LOC_464/a_8_216# OR2X1_LOC_464/a_36_216# OR2X1_LOC_471/B VSS VDD
+ OR2X1_LOC_464/A OR2X1_LOC_464/B OR2X1_LOC
XOR2X1_LOC_475 OR2X1_LOC_475/a_8_216# OR2X1_LOC_475/a_36_216# OR2X1_LOC_475/Y VSS VDD
+ OR2X1_LOC_474/Y OR2X1_LOC_475/B OR2X1_LOC
XOR2X1_LOC_497 OR2X1_LOC_497/a_8_216# OR2X1_LOC_497/a_36_216# OR2X1_LOC_497/Y VSS VDD
+ OR2X1_LOC_71/Y OR2X1_LOC_22/Y OR2X1_LOC
XOR2X1_LOC_486 OR2X1_LOC_486/a_8_216# OR2X1_LOC_486/a_36_216# OR2X1_LOC_486/Y VSS VDD
+ OR2X1_LOC_705/B OR2X1_LOC_486/B OR2X1_LOC
XOR2X1_LOC_261 OR2X1_LOC_261/a_8_216# OR2X1_LOC_261/a_36_216# OR2X1_LOC_261/Y VSS VDD
+ OR2X1_LOC_261/A OR2X1_LOC_600/A OR2X1_LOC
XOR2X1_LOC_294 OR2X1_LOC_294/a_8_216# OR2X1_LOC_294/a_36_216# OR2X1_LOC_294/Y VSS VDD
+ OR2X1_LOC_598/A AND2X1_LOC_41/A OR2X1_LOC
XOR2X1_LOC_250 OR2X1_LOC_250/a_8_216# OR2X1_LOC_250/a_36_216# OR2X1_LOC_250/Y VSS VDD
+ OR2X1_LOC_595/A OR2X1_LOC_64/Y OR2X1_LOC
XOR2X1_LOC_283 OR2X1_LOC_283/a_8_216# OR2X1_LOC_283/a_36_216# OR2X1_LOC_283/Y VSS VDD
+ OR2X1_LOC_417/A OR2X1_LOC_26/Y OR2X1_LOC
XOR2X1_LOC_272 OR2X1_LOC_272/a_8_216# OR2X1_LOC_272/a_36_216# OR2X1_LOC_272/Y VSS VDD
+ OR2X1_LOC_43/A OR2X1_LOC_31/Y OR2X1_LOC
XAND2X1_LOC_518 AND2X1_LOC_518/a_36_24# OR2X1_LOC_520/B AND2X1_LOC_518/a_8_24# VSS VDD
+ AND2X1_LOC_64/Y OR2X1_LOC_185/A AND2X1_LOC
XAND2X1_LOC_507 AND2X1_LOC_507/a_36_24# AND2X1_LOC_508/B AND2X1_LOC_507/a_8_24# VSS VDD
+ OR2X1_LOC_504/Y OR2X1_LOC_505/Y AND2X1_LOC
XAND2X1_LOC_529 AND2X1_LOC_529/a_36_24# OR2X1_LOC_548/B AND2X1_LOC_529/a_8_24# VSS VDD
+ INPUT_3 OR2X1_LOC_66/A AND2X1_LOC
XOR2X1_LOC_805 OR2X1_LOC_805/a_8_216# OR2X1_LOC_805/a_36_216# OR2X1_LOC_807/B VSS VDD
+ OR2X1_LOC_805/A OR2X1_LOC_792/Y OR2X1_LOC
XOR2X1_LOC_827 OR2X1_LOC_827/a_8_216# OR2X1_LOC_827/a_36_216# OR2X1_LOC_827/Y VSS VDD
+ OR2X1_LOC_158/A OR2X1_LOC_43/A OR2X1_LOC
XOR2X1_LOC_849 OR2X1_LOC_849/a_8_216# OR2X1_LOC_849/a_36_216# OR2X1_LOC_859/A VSS VDD
+ OR2X1_LOC_849/A OR2X1_LOC_844/Y OR2X1_LOC
XOR2X1_LOC_816 OR2X1_LOC_816/a_8_216# OR2X1_LOC_816/a_36_216# OR2X1_LOC_816/Y VSS VDD
+ OR2X1_LOC_816/A OR2X1_LOC_51/Y OR2X1_LOC
XOR2X1_LOC_838 OR2X1_LOC_838/a_8_216# OR2X1_LOC_838/a_36_216# OR2X1_LOC_852/B VSS VDD
+ OR2X1_LOC_837/Y OR2X1_LOC_838/B OR2X1_LOC
XAND2X1_LOC_315 AND2X1_LOC_315/a_36_24# OR2X1_LOC_318/B AND2X1_LOC_315/a_8_24# VSS VDD
+ AND2X1_LOC_31/Y OR2X1_LOC_161/B AND2X1_LOC
XAND2X1_LOC_359 AND2X1_LOC_359/a_36_24# AND2X1_LOC_363/A AND2X1_LOC_359/a_8_24# VSS VDD
+ AND2X1_LOC_348/Y AND2X1_LOC_359/B AND2X1_LOC
XAND2X1_LOC_348 AND2X1_LOC_348/a_36_24# AND2X1_LOC_348/Y AND2X1_LOC_348/a_8_24# VSS VDD
+ AND2X1_LOC_348/A AND2X1_LOC_345/Y AND2X1_LOC
XAND2X1_LOC_326 AND2X1_LOC_326/a_36_24# AND2X1_LOC_354/B AND2X1_LOC_326/a_8_24# VSS VDD
+ AND2X1_LOC_326/A AND2X1_LOC_326/B AND2X1_LOC
XAND2X1_LOC_337 AND2X1_LOC_337/a_36_24# AND2X1_LOC_352/B AND2X1_LOC_337/a_8_24# VSS VDD
+ AND2X1_LOC_335/Y AND2X1_LOC_337/B AND2X1_LOC
XAND2X1_LOC_304 AND2X1_LOC_304/a_36_24# OR2X1_LOC_307/B AND2X1_LOC_304/a_8_24# VSS VDD
+ AND2X1_LOC_53/Y OR2X1_LOC_269/B AND2X1_LOC
XOR2X1_LOC_635 OR2X1_LOC_635/a_8_216# OR2X1_LOC_635/a_36_216# OR2X1_LOC_639/B VSS VDD
+ OR2X1_LOC_635/A OR2X1_LOC_451/B OR2X1_LOC
XAND2X1_LOC_88 AND2X1_LOC_88/a_36_24# AND2X1_LOC_88/Y AND2X1_LOC_88/a_8_24# VSS VDD
+ AND2X1_LOC_3/Y OR2X1_LOC_87/Y AND2X1_LOC
XAND2X1_LOC_66 AND2X1_LOC_66/a_36_24# OR2X1_LOC_67/A AND2X1_LOC_66/a_8_24# VSS VDD
+ OR2X1_LOC_3/Y OR2X1_LOC_26/Y AND2X1_LOC
XAND2X1_LOC_99 AND2X1_LOC_99/a_36_24# AND2X1_LOC_99/Y AND2X1_LOC_99/a_8_24# VSS VDD
+ AND2X1_LOC_99/A AND2X1_LOC_98/Y AND2X1_LOC
XAND2X1_LOC_55 AND2X1_LOC_55/a_36_24# AND2X1_LOC_56/B AND2X1_LOC_55/a_8_24# VSS VDD
+ OR2X1_LOC_68/B OR2X1_LOC_62/A AND2X1_LOC
XAND2X1_LOC_77 AND2X1_LOC_77/a_36_24# OR2X1_LOC_78/A AND2X1_LOC_77/a_8_24# VSS VDD
+ OR2X1_LOC_377/A OR2X1_LOC_62/A AND2X1_LOC
XAND2X1_LOC_33 AND2X1_LOC_33/a_36_24# AND2X1_LOC_33/Y AND2X1_LOC_33/a_8_24# VSS VDD
+ OR2X1_LOC_20/Y OR2X1_LOC_24/Y AND2X1_LOC
XAND2X1_LOC_22 AND2X1_LOC_22/a_36_24# AND2X1_LOC_22/Y AND2X1_LOC_22/a_8_24# VSS VDD
+ AND2X1_LOC_1/Y AND2X1_LOC_21/Y AND2X1_LOC
XAND2X1_LOC_44 AND2X1_LOC_44/a_36_24# AND2X1_LOC_44/Y AND2X1_LOC_44/a_8_24# VSS VDD
+ AND2X1_LOC_17/Y AND2X1_LOC_51/A AND2X1_LOC
XAND2X1_LOC_11 AND2X1_LOC_11/a_36_24# AND2X1_LOC_11/Y AND2X1_LOC_11/a_8_24# VSS VDD
+ D_INPUT_4 INPUT_5 AND2X1_LOC
XOR2X1_LOC_624 OR2X1_LOC_624/a_8_216# OR2X1_LOC_624/a_36_216# OR2X1_LOC_624/Y VSS VDD
+ OR2X1_LOC_624/A OR2X1_LOC_624/B OR2X1_LOC
XOR2X1_LOC_613 OR2X1_LOC_613/a_8_216# OR2X1_LOC_613/a_36_216# OR2X1_LOC_613/Y VSS VDD
+ OR2X1_LOC_56/A OR2X1_LOC_40/Y OR2X1_LOC
XOR2X1_LOC_602 OR2X1_LOC_602/a_8_216# OR2X1_LOC_602/a_36_216# OR2X1_LOC_602/Y VSS VDD
+ OR2X1_LOC_602/A OR2X1_LOC_602/B OR2X1_LOC
XOR2X1_LOC_679 OR2X1_LOC_679/a_8_216# OR2X1_LOC_679/a_36_216# OR2X1_LOC_679/Y VSS VDD
+ OR2X1_LOC_679/A OR2X1_LOC_679/B OR2X1_LOC
XAND2X1_LOC_860 AND2X1_LOC_860/a_36_24# AND2X1_LOC_861/B AND2X1_LOC_860/a_8_24# VSS VDD
+ AND2X1_LOC_860/A AND2X1_LOC_474/A AND2X1_LOC
XOR2X1_LOC_668 OR2X1_LOC_668/a_8_216# OR2X1_LOC_668/a_36_216# OR2X1_LOC_668/Y VSS VDD
+ OR2X1_LOC_375/A OR2X1_LOC_66/A OR2X1_LOC
XOR2X1_LOC_657 OR2X1_LOC_657/a_8_216# OR2X1_LOC_657/a_36_216# OR2X1_LOC_659/B VSS VDD
+ OR2X1_LOC_510/Y OR2X1_LOC_217/A OR2X1_LOC
XOR2X1_LOC_646 OR2X1_LOC_646/a_8_216# OR2X1_LOC_646/a_36_216# OR2X1_LOC_647/A VSS VDD
+ OR2X1_LOC_646/A OR2X1_LOC_646/B OR2X1_LOC
XAND2X1_LOC_101 AND2X1_LOC_101/a_36_24# AND2X1_LOC_216/A AND2X1_LOC_101/a_8_24# VSS VDD
+ AND2X1_LOC_99/Y AND2X1_LOC_101/B AND2X1_LOC
XAND2X1_LOC_112 AND2X1_LOC_112/a_36_24# AND2X1_LOC_715/A AND2X1_LOC_112/a_8_24# VSS VDD
+ OR2X1_LOC_109/Y OR2X1_LOC_111/Y AND2X1_LOC
XAND2X1_LOC_189 AND2X1_LOC_189/a_36_24# OR2X1_LOC_192/B AND2X1_LOC_189/a_8_24# VSS VDD
+ AND2X1_LOC_95/Y OR2X1_LOC_188/Y AND2X1_LOC
XAND2X1_LOC_178 AND2X1_LOC_178/a_36_24# OR2X1_LOC_181/B AND2X1_LOC_178/a_8_24# VSS VDD
+ AND2X1_LOC_56/B OR2X1_LOC_375/A AND2X1_LOC
XAND2X1_LOC_123 AND2X1_LOC_123/a_36_24# AND2X1_LOC_123/Y AND2X1_LOC_123/a_8_24# VSS VDD
+ OR2X1_LOC_117/Y OR2X1_LOC_118/Y AND2X1_LOC
XAND2X1_LOC_134 AND2X1_LOC_134/a_36_24# OR2X1_LOC_768/A AND2X1_LOC_134/a_8_24# VSS VDD
+ AND2X1_LOC_95/Y OR2X1_LOC_161/B AND2X1_LOC
XAND2X1_LOC_167 AND2X1_LOC_167/a_36_24# OR2X1_LOC_703/B AND2X1_LOC_167/a_8_24# VSS VDD
+ AND2X1_LOC_64/Y OR2X1_LOC_161/A AND2X1_LOC
XAND2X1_LOC_145 AND2X1_LOC_145/a_36_24# OR2X1_LOC_148/B AND2X1_LOC_145/a_8_24# VSS VDD
+ AND2X1_LOC_51/Y OR2X1_LOC_78/A AND2X1_LOC
XAND2X1_LOC_156 AND2X1_LOC_156/a_36_24# OR2X1_LOC_158/B AND2X1_LOC_156/a_8_24# VSS VDD
+ AND2X1_LOC_154/Y AND2X1_LOC_155/Y AND2X1_LOC
XOR2X1_LOC_454 OR2X1_LOC_454/a_8_216# OR2X1_LOC_454/a_36_216# OR2X1_LOC_466/A VSS VDD
+ OR2X1_LOC_447/Y OR2X1_LOC_446/Y OR2X1_LOC
XOR2X1_LOC_421 OR2X1_LOC_421/a_8_216# OR2X1_LOC_421/a_36_216# OR2X1_LOC_421/Y VSS VDD
+ OR2X1_LOC_421/A OR2X1_LOC_91/A OR2X1_LOC
XOR2X1_LOC_432 OR2X1_LOC_432/a_8_216# OR2X1_LOC_432/a_36_216# OR2X1_LOC_432/Y VSS VDD
+ OR2X1_LOC_589/A OR2X1_LOC_18/Y OR2X1_LOC
XOR2X1_LOC_465 OR2X1_LOC_465/a_8_216# OR2X1_LOC_465/a_36_216# OR2X1_LOC_465/Y VSS VDD
+ OR2X1_LOC_456/Y OR2X1_LOC_465/B OR2X1_LOC
XOR2X1_LOC_487 OR2X1_LOC_487/a_8_216# OR2X1_LOC_487/a_36_216# OR2X1_LOC_487/Y VSS VDD
+ OR2X1_LOC_95/Y OR2X1_LOC_45/B OR2X1_LOC
XOR2X1_LOC_476 OR2X1_LOC_476/a_8_216# OR2X1_LOC_476/a_36_216# OR2X1_LOC_476/Y VSS VDD
+ OR2X1_LOC_473/Y OR2X1_LOC_476/B OR2X1_LOC
XOR2X1_LOC_443 OR2X1_LOC_443/a_8_216# OR2X1_LOC_443/a_36_216# OR2X1_LOC_443/Y VSS VDD
+ OR2X1_LOC_545/B OR2X1_LOC_97/A OR2X1_LOC
XOR2X1_LOC_410 OR2X1_LOC_410/a_8_216# OR2X1_LOC_410/a_36_216# OR2X1_LOC_410/Y VSS VDD
+ AND2X1_LOC_51/Y AND2X1_LOC_12/Y OR2X1_LOC
XAND2X1_LOC_690 AND2X1_LOC_690/a_36_24# OR2X1_LOC_691/A AND2X1_LOC_690/a_8_24# VSS VDD
+ D_INPUT_0 OR2X1_LOC_634/A AND2X1_LOC
XOR2X1_LOC_498 OR2X1_LOC_498/a_8_216# OR2X1_LOC_498/a_36_216# OR2X1_LOC_498/Y VSS VDD
+ OR2X1_LOC_189/A OR2X1_LOC_70/Y OR2X1_LOC
XOR2X1_LOC_295 OR2X1_LOC_295/a_8_216# OR2X1_LOC_295/a_36_216# OR2X1_LOC_295/Y VSS VDD
+ OR2X1_LOC_481/A OR2X1_LOC_59/Y OR2X1_LOC
XOR2X1_LOC_284 OR2X1_LOC_284/a_8_216# OR2X1_LOC_284/a_36_216# OR2X1_LOC_287/A VSS VDD
+ OR2X1_LOC_542/B OR2X1_LOC_284/B OR2X1_LOC
XOR2X1_LOC_251 OR2X1_LOC_251/a_8_216# OR2X1_LOC_251/a_36_216# OR2X1_LOC_251/Y VSS VDD
+ OR2X1_LOC_106/A OR2X1_LOC_51/Y OR2X1_LOC
XOR2X1_LOC_240 OR2X1_LOC_240/a_8_216# OR2X1_LOC_240/a_36_216# OR2X1_LOC_243/A VSS VDD
+ OR2X1_LOC_240/A OR2X1_LOC_240/B OR2X1_LOC
XOR2X1_LOC_262 OR2X1_LOC_262/a_8_216# OR2X1_LOC_262/a_36_216# OR2X1_LOC_262/Y VSS VDD
+ OR2X1_LOC_65/B OR2X1_LOC_40/Y OR2X1_LOC
XOR2X1_LOC_273 OR2X1_LOC_273/a_8_216# OR2X1_LOC_273/a_36_216# OR2X1_LOC_273/Y VSS VDD
+ OR2X1_LOC_743/A OR2X1_LOC_36/Y OR2X1_LOC
XAND2X1_LOC_519 AND2X1_LOC_519/a_36_24# OR2X1_LOC_520/A AND2X1_LOC_519/a_8_24# VSS VDD
+ AND2X1_LOC_48/A OR2X1_LOC_375/A AND2X1_LOC
XAND2X1_LOC_508 AND2X1_LOC_508/a_36_24# AND2X1_LOC_510/A AND2X1_LOC_508/a_8_24# VSS VDD
+ AND2X1_LOC_508/A AND2X1_LOC_508/B AND2X1_LOC
XOR2X1_LOC_828 OR2X1_LOC_828/a_8_216# OR2X1_LOC_828/a_36_216# OR2X1_LOC_828/Y VSS VDD
+ OR2X1_LOC_598/Y OR2X1_LOC_828/B OR2X1_LOC
XOR2X1_LOC_806 OR2X1_LOC_806/a_8_216# OR2X1_LOC_806/a_36_216# OR2X1_LOC_807/A VSS VDD
+ OR2X1_LOC_675/Y OR2X1_LOC_362/B OR2X1_LOC
XOR2X1_LOC_817 OR2X1_LOC_817/a_8_216# OR2X1_LOC_817/a_36_216# OR2X1_LOC_817/Y VSS VDD
+ OR2X1_LOC_382/A INPUT_1 OR2X1_LOC
XOR2X1_LOC_839 OR2X1_LOC_839/a_8_216# OR2X1_LOC_839/a_36_216# OR2X1_LOC_852/A VSS VDD
+ OR2X1_LOC_836/Y OR2X1_LOC_835/Y OR2X1_LOC
XAND2X1_LOC_316 AND2X1_LOC_316/a_36_24# OR2X1_LOC_318/A AND2X1_LOC_316/a_8_24# VSS VDD
+ AND2X1_LOC_12/Y AND2X1_LOC_81/B AND2X1_LOC
XAND2X1_LOC_349 AND2X1_LOC_349/a_36_24# AND2X1_LOC_359/B AND2X1_LOC_349/a_8_24# VSS VDD
+ AND2X1_LOC_342/Y AND2X1_LOC_349/B AND2X1_LOC
XAND2X1_LOC_327 AND2X1_LOC_327/a_36_24# OR2X1_LOC_329/B AND2X1_LOC_327/a_8_24# VSS VDD
+ OR2X1_LOC_65/B OR2X1_LOC_517/A AND2X1_LOC
XAND2X1_LOC_338 AND2X1_LOC_338/a_36_24# AND2X1_LOC_338/Y AND2X1_LOC_338/a_8_24# VSS VDD
+ AND2X1_LOC_338/A AND2X1_LOC_334/Y AND2X1_LOC
XAND2X1_LOC_305 AND2X1_LOC_305/a_36_24# OR2X1_LOC_307/A AND2X1_LOC_305/a_8_24# VSS VDD
+ AND2X1_LOC_3/Y AND2X1_LOC_91/B AND2X1_LOC
XAND2X1_LOC_34 AND2X1_LOC_34/a_36_24# AND2X1_LOC_34/Y AND2X1_LOC_34/a_8_24# VSS VDD
+ OR2X1_LOC_27/Y OR2X1_LOC_32/Y AND2X1_LOC
XAND2X1_LOC_23 AND2X1_LOC_23/a_36_24# OR2X1_LOC_160/B AND2X1_LOC_23/a_8_24# VSS VDD
+ OR2X1_LOC_19/B OR2X1_LOC_377/A AND2X1_LOC
XAND2X1_LOC_12 AND2X1_LOC_12/a_36_24# AND2X1_LOC_12/Y AND2X1_LOC_12/a_8_24# VSS VDD
+ AND2X1_LOC_1/Y AND2X1_LOC_11/Y AND2X1_LOC
XOR2X1_LOC_603 OR2X1_LOC_603/a_8_216# OR2X1_LOC_603/a_36_216# OR2X1_LOC_603/Y VSS VDD
+ OR2X1_LOC_52/B OR2X1_LOC_12/Y OR2X1_LOC
XOR2X1_LOC_636 OR2X1_LOC_636/a_8_216# OR2X1_LOC_636/a_36_216# OR2X1_LOC_639/A VSS VDD
+ OR2X1_LOC_636/A OR2X1_LOC_636/B OR2X1_LOC
XOR2X1_LOC_614 OR2X1_LOC_614/a_8_216# OR2X1_LOC_614/a_36_216# OR2X1_LOC_614/Y VSS VDD
+ OR2X1_LOC_161/B OR2X1_LOC_78/A OR2X1_LOC
XAND2X1_LOC_67 AND2X1_LOC_67/a_36_24# AND2X1_LOC_67/Y AND2X1_LOC_67/a_8_24# VSS VDD
+ AND2X1_LOC_56/B OR2X1_LOC_66/Y AND2X1_LOC
XAND2X1_LOC_850 AND2X1_LOC_850/a_36_24# AND2X1_LOC_850/Y AND2X1_LOC_850/a_8_24# VSS VDD
+ AND2X1_LOC_850/A AND2X1_LOC_843/Y AND2X1_LOC
XAND2X1_LOC_89 AND2X1_LOC_89/a_36_24# OR2X1_LOC_97/B AND2X1_LOC_89/a_8_24# VSS VDD
+ AND2X1_LOC_59/Y OR2X1_LOC_78/A AND2X1_LOC
XAND2X1_LOC_78 AND2X1_LOC_78/a_36_24# OR2X1_LOC_79/A AND2X1_LOC_78/a_8_24# VSS VDD
+ OR2X1_LOC_16/A OR2X1_LOC_89/A AND2X1_LOC
XAND2X1_LOC_45 AND2X1_LOC_45/a_36_24# OR2X1_LOC_196/B AND2X1_LOC_45/a_8_24# VSS VDD
+ OR2X1_LOC_160/B AND2X1_LOC_44/Y AND2X1_LOC
XAND2X1_LOC_56 AND2X1_LOC_56/a_36_24# OR2X1_LOC_197/A AND2X1_LOC_56/a_8_24# VSS VDD
+ AND2X1_LOC_53/Y AND2X1_LOC_56/B AND2X1_LOC
XOR2X1_LOC_658 OR2X1_LOC_658/a_8_216# OR2X1_LOC_658/a_36_216# OR2X1_LOC_659/A VSS VDD
+ OR2X1_LOC_632/Y OR2X1_LOC_624/Y OR2X1_LOC
XOR2X1_LOC_625 OR2X1_LOC_625/a_8_216# OR2X1_LOC_625/a_36_216# OR2X1_LOC_625/Y VSS VDD
+ OR2X1_LOC_585/A OR2X1_LOC_67/A OR2X1_LOC
XOR2X1_LOC_669 OR2X1_LOC_669/a_8_216# OR2X1_LOC_669/a_36_216# OR2X1_LOC_669/Y VSS VDD
+ OR2X1_LOC_669/A OR2X1_LOC_604/A OR2X1_LOC
XOR2X1_LOC_647 OR2X1_LOC_647/a_8_216# OR2X1_LOC_647/a_36_216# OR2X1_LOC_647/Y VSS VDD
+ OR2X1_LOC_647/A OR2X1_LOC_647/B OR2X1_LOC
XAND2X1_LOC_861 AND2X1_LOC_861/a_36_24# AND2X1_LOC_865/A AND2X1_LOC_861/a_8_24# VSS VDD
+ AND2X1_LOC_658/A AND2X1_LOC_861/B AND2X1_LOC
XAND2X1_LOC_113 AND2X1_LOC_113/a_36_24# AND2X1_LOC_113/Y AND2X1_LOC_113/a_8_24# VSS VDD
+ OR2X1_LOC_103/Y OR2X1_LOC_107/Y AND2X1_LOC
XAND2X1_LOC_124 AND2X1_LOC_124/a_36_24# AND2X1_LOC_572/A AND2X1_LOC_124/a_8_24# VSS VDD
+ OR2X1_LOC_122/Y AND2X1_LOC_123/Y AND2X1_LOC
XAND2X1_LOC_102 AND2X1_LOC_102/a_36_24# OR2X1_LOC_532/B AND2X1_LOC_102/a_8_24# VSS VDD
+ AND2X1_LOC_8/Y OR2X1_LOC_62/A AND2X1_LOC
XAND2X1_LOC_135 AND2X1_LOC_135/a_36_24# OR2X1_LOC_702/A AND2X1_LOC_135/a_8_24# VSS VDD
+ AND2X1_LOC_59/Y OR2X1_LOC_161/B AND2X1_LOC
XAND2X1_LOC_146 AND2X1_LOC_146/a_36_24# OR2X1_LOC_148/A AND2X1_LOC_146/a_8_24# VSS VDD
+ AND2X1_LOC_36/Y OR2X1_LOC_160/A AND2X1_LOC
XAND2X1_LOC_179 AND2X1_LOC_179/a_36_24# OR2X1_LOC_181/A AND2X1_LOC_179/a_8_24# VSS VDD
+ AND2X1_LOC_36/Y OR2X1_LOC_756/B AND2X1_LOC
XAND2X1_LOC_168 AND2X1_LOC_168/a_36_24# AND2X1_LOC_168/Y AND2X1_LOC_168/a_8_24# VSS VDD
+ OR2X1_LOC_164/Y OR2X1_LOC_165/Y AND2X1_LOC
XAND2X1_LOC_157 AND2X1_LOC_157/a_36_24# OR2X1_LOC_375/A AND2X1_LOC_157/a_8_24# VSS VDD
+ AND2X1_LOC_2/Y AND2X1_LOC_17/Y AND2X1_LOC
XOR2X1_LOC_466 OR2X1_LOC_466/a_8_216# OR2X1_LOC_466/a_36_216# OR2X1_LOC_470/B VSS VDD
+ OR2X1_LOC_466/A OR2X1_LOC_453/Y OR2X1_LOC
XOR2X1_LOC_477 OR2X1_LOC_477/a_8_216# OR2X1_LOC_477/a_36_216# OR2X1_LOC_477/Y VSS VDD
+ OR2X1_LOC_471/Y OR2X1_LOC_477/B OR2X1_LOC
XOR2X1_LOC_422 OR2X1_LOC_422/a_8_216# OR2X1_LOC_422/a_36_216# OR2X1_LOC_422/Y VSS VDD
+ OR2X1_LOC_92/Y OR2X1_LOC_12/Y OR2X1_LOC
XOR2X1_LOC_433 OR2X1_LOC_433/a_8_216# OR2X1_LOC_433/a_36_216# OR2X1_LOC_433/Y VSS VDD
+ OR2X1_LOC_743/A OR2X1_LOC_70/Y OR2X1_LOC
XAND2X1_LOC_680 AND2X1_LOC_680/a_36_24# OR2X1_LOC_728/A AND2X1_LOC_680/a_8_24# VSS VDD
+ AND2X1_LOC_51/Y OR2X1_LOC_186/Y AND2X1_LOC
XAND2X1_LOC_691 AND2X1_LOC_691/a_36_24# AND2X1_LOC_729/B AND2X1_LOC_691/a_8_24# VSS VDD
+ OR2X1_LOC_689/Y OR2X1_LOC_690/Y AND2X1_LOC
XOR2X1_LOC_400 OR2X1_LOC_400/a_8_216# OR2X1_LOC_400/a_36_216# OR2X1_LOC_403/A VSS VDD
+ OR2X1_LOC_400/A OR2X1_LOC_400/B OR2X1_LOC
XOR2X1_LOC_499 OR2X1_LOC_499/a_8_216# OR2X1_LOC_499/a_36_216# OR2X1_LOC_500/A VSS VDD
+ OR2X1_LOC_778/A OR2X1_LOC_499/B OR2X1_LOC
XOR2X1_LOC_455 OR2X1_LOC_455/a_8_216# OR2X1_LOC_455/a_36_216# OR2X1_LOC_465/B VSS VDD
+ OR2X1_LOC_455/A OR2X1_LOC_76/Y OR2X1_LOC
XOR2X1_LOC_488 OR2X1_LOC_488/a_8_216# OR2X1_LOC_488/a_36_216# OR2X1_LOC_488/Y VSS VDD
+ OR2X1_LOC_417/A OR2X1_LOC_158/A OR2X1_LOC
XOR2X1_LOC_444 OR2X1_LOC_444/a_8_216# OR2X1_LOC_444/a_36_216# OR2X1_LOC_469/B VSS VDD
+ OR2X1_LOC_443/Y OR2X1_LOC_444/B OR2X1_LOC
XOR2X1_LOC_411 OR2X1_LOC_411/a_8_216# OR2X1_LOC_411/a_36_216# OR2X1_LOC_411/Y VSS VDD
+ OR2X1_LOC_411/A OR2X1_LOC_600/A OR2X1_LOC
XOR2X1_LOC_285 OR2X1_LOC_285/a_8_216# OR2X1_LOC_285/a_36_216# OR2X1_LOC_285/Y VSS VDD
+ OR2X1_LOC_285/A OR2X1_LOC_285/B OR2X1_LOC
XOR2X1_LOC_252 OR2X1_LOC_252/a_8_216# OR2X1_LOC_252/a_36_216# OR2X1_LOC_252/Y VSS VDD
+ OR2X1_LOC_59/Y OR2X1_LOC_56/A OR2X1_LOC
XOR2X1_LOC_296 OR2X1_LOC_296/a_8_216# OR2X1_LOC_296/a_36_216# OR2X1_LOC_296/Y VSS VDD
+ AND2X1_LOC_56/B AND2X1_LOC_43/B OR2X1_LOC
XOR2X1_LOC_263 OR2X1_LOC_263/a_8_216# OR2X1_LOC_263/a_36_216# OR2X1_LOC_813/A VSS VDD
+ OR2X1_LOC_85/A OR2X1_LOC_22/Y OR2X1_LOC
XOR2X1_LOC_274 OR2X1_LOC_274/a_8_216# OR2X1_LOC_274/a_36_216# OR2X1_LOC_274/Y VSS VDD
+ OR2X1_LOC_831/B OR2X1_LOC_541/A OR2X1_LOC
XOR2X1_LOC_241 OR2X1_LOC_241/a_8_216# OR2X1_LOC_241/a_36_216# OR2X1_LOC_241/Y VSS VDD
+ OR2X1_LOC_776/A OR2X1_LOC_241/B OR2X1_LOC
XOR2X1_LOC_230 OR2X1_LOC_230/a_8_216# OR2X1_LOC_230/a_36_216# OR2X1_LOC_230/Y VSS VDD
+ OR2X1_LOC_31/Y OR2X1_LOC_7/A OR2X1_LOC
XAND2X1_LOC_509 AND2X1_LOC_509/a_36_24# AND2X1_LOC_509/Y AND2X1_LOC_509/a_8_24# VSS VDD
+ AND2X1_LOC_227/Y OR2X1_LOC_503/Y AND2X1_LOC
XOR2X1_LOC_829 OR2X1_LOC_829/a_8_216# OR2X1_LOC_829/a_36_216# OR2X1_LOC_829/Y VSS VDD
+ OR2X1_LOC_829/A OR2X1_LOC_64/Y OR2X1_LOC
XOR2X1_LOC_807 OR2X1_LOC_807/a_8_216# OR2X1_LOC_807/a_36_216# OR2X1_LOC_807/Y VSS VDD
+ OR2X1_LOC_807/A OR2X1_LOC_807/B OR2X1_LOC
XOR2X1_LOC_818 OR2X1_LOC_818/a_8_216# OR2X1_LOC_818/a_36_216# OR2X1_LOC_818/Y VSS VDD
+ OR2X1_LOC_502/A OR2X1_LOC_68/B OR2X1_LOC
XAND2X1_LOC_306 AND2X1_LOC_306/a_36_24# OR2X1_LOC_512/A AND2X1_LOC_306/a_8_24# VSS VDD
+ AND2X1_LOC_22/Y OR2X1_LOC_502/A AND2X1_LOC
XAND2X1_LOC_328 AND2X1_LOC_328/a_36_24# OR2X1_LOC_596/A AND2X1_LOC_328/a_8_24# VSS VDD
+ D_INPUT_4 AND2X1_LOC_50/Y AND2X1_LOC
XAND2X1_LOC_317 AND2X1_LOC_317/a_36_24# AND2X1_LOC_319/A AND2X1_LOC_317/a_8_24# VSS VDD
+ OR2X1_LOC_313/Y OR2X1_LOC_314/Y AND2X1_LOC
XAND2X1_LOC_339 AND2X1_LOC_339/a_36_24# AND2X1_LOC_339/Y AND2X1_LOC_339/a_8_24# VSS VDD
+ AND2X1_LOC_61/Y AND2X1_LOC_339/B AND2X1_LOC
XAND2X1_LOC_46 AND2X1_LOC_46/a_36_24# AND2X1_LOC_48/A AND2X1_LOC_46/a_8_24# VSS VDD
+ D_INPUT_1 OR2X1_LOC_377/A AND2X1_LOC
XAND2X1_LOC_68 AND2X1_LOC_68/a_36_24# OR2X1_LOC_69/A AND2X1_LOC_68/a_8_24# VSS VDD
+ OR2X1_LOC_6/A OR2X1_LOC_52/B AND2X1_LOC
XAND2X1_LOC_24 AND2X1_LOC_24/a_36_24# OR2X1_LOC_33/A AND2X1_LOC_24/a_8_24# VSS VDD
+ AND2X1_LOC_22/Y OR2X1_LOC_160/B AND2X1_LOC
XAND2X1_LOC_57 AND2X1_LOC_57/a_36_24# AND2X1_LOC_57/Y AND2X1_LOC_57/a_8_24# VSS VDD
+ OR2X1_LOC_68/B AND2X1_LOC_44/Y AND2X1_LOC
XAND2X1_LOC_35 AND2X1_LOC_35/a_36_24# AND2X1_LOC_35/Y AND2X1_LOC_35/a_8_24# VSS VDD
+ AND2X1_LOC_33/Y AND2X1_LOC_34/Y AND2X1_LOC
XAND2X1_LOC_13 AND2X1_LOC_13/a_36_24# OR2X1_LOC_193/A AND2X1_LOC_13/a_8_24# VSS VDD
+ AND2X1_LOC_41/A AND2X1_LOC_12/Y AND2X1_LOC
XOR2X1_LOC_604 OR2X1_LOC_604/a_8_216# OR2X1_LOC_604/a_36_216# OR2X1_LOC_604/Y VSS VDD
+ OR2X1_LOC_604/A OR2X1_LOC_70/Y OR2X1_LOC
XOR2X1_LOC_637 OR2X1_LOC_637/a_8_216# OR2X1_LOC_637/a_36_216# OR2X1_LOC_637/Y VSS VDD
+ OR2X1_LOC_637/A OR2X1_LOC_637/B OR2X1_LOC
XAND2X1_LOC_862 AND2X1_LOC_862/a_36_24# AND2X1_LOC_862/Y AND2X1_LOC_862/a_8_24# VSS VDD
+ AND2X1_LOC_862/A AND2X1_LOC_859/Y AND2X1_LOC
XAND2X1_LOC_79 AND2X1_LOC_79/a_36_24# AND2X1_LOC_79/Y AND2X1_LOC_79/a_8_24# VSS VDD
+ AND2X1_LOC_18/Y OR2X1_LOC_78/Y AND2X1_LOC
XAND2X1_LOC_851 AND2X1_LOC_851/a_36_24# AND2X1_LOC_858/B AND2X1_LOC_851/a_8_24# VSS VDD
+ AND2X1_LOC_851/A AND2X1_LOC_851/B AND2X1_LOC
XAND2X1_LOC_840 AND2X1_LOC_840/a_36_24# AND2X1_LOC_851/A AND2X1_LOC_840/a_8_24# VSS VDD
+ AND2X1_LOC_840/A AND2X1_LOC_840/B AND2X1_LOC
XOR2X1_LOC_659 OR2X1_LOC_659/a_8_216# OR2X1_LOC_659/a_36_216# OR2X1_LOC_659/Y VSS VDD
+ OR2X1_LOC_659/A OR2X1_LOC_659/B OR2X1_LOC
XOR2X1_LOC_626 OR2X1_LOC_626/a_8_216# OR2X1_LOC_626/a_36_216# OR2X1_LOC_626/Y VSS VDD
+ OR2X1_LOC_604/A OR2X1_LOC_95/Y OR2X1_LOC
XOR2X1_LOC_615 OR2X1_LOC_615/a_8_216# OR2X1_LOC_615/a_36_216# OR2X1_LOC_615/Y VSS VDD
+ OR2X1_LOC_754/A OR2X1_LOC_22/Y OR2X1_LOC
XOR2X1_LOC_648 OR2X1_LOC_648/a_8_216# OR2X1_LOC_648/a_36_216# OR2X1_LOC_655/B VSS VDD
+ OR2X1_LOC_648/A OR2X1_LOC_648/B OR2X1_LOC
XAND2X1_LOC_103 AND2X1_LOC_103/a_36_24# OR2X1_LOC_113/B AND2X1_LOC_103/a_8_24# VSS VDD
+ AND2X1_LOC_47/Y OR2X1_LOC_532/B AND2X1_LOC
XAND2X1_LOC_125 AND2X1_LOC_125/a_36_24# OR2X1_LOC_128/B AND2X1_LOC_125/a_8_24# VSS VDD
+ AND2X1_LOC_95/Y OR2X1_LOC_756/B AND2X1_LOC
XAND2X1_LOC_114 AND2X1_LOC_114/a_36_24# AND2X1_LOC_114/Y AND2X1_LOC_114/a_8_24# VSS VDD
+ OR2X1_LOC_108/Y AND2X1_LOC_113/Y AND2X1_LOC
XAND2X1_LOC_136 AND2X1_LOC_136/a_36_24# OR2X1_LOC_138/A AND2X1_LOC_136/a_8_24# VSS VDD
+ AND2X1_LOC_3/Y AND2X1_LOC_43/B AND2X1_LOC
XAND2X1_LOC_169 AND2X1_LOC_169/a_36_24# AND2X1_LOC_170/B AND2X1_LOC_169/a_8_24# VSS VDD
+ OR2X1_LOC_166/Y OR2X1_LOC_167/Y AND2X1_LOC
XAND2X1_LOC_147 AND2X1_LOC_147/a_36_24# AND2X1_LOC_147/Y AND2X1_LOC_147/a_8_24# VSS VDD
+ OR2X1_LOC_142/Y OR2X1_LOC_144/Y AND2X1_LOC
XAND2X1_LOC_158 AND2X1_LOC_158/a_36_24# OR2X1_LOC_210/B AND2X1_LOC_158/a_8_24# VSS VDD
+ OR2X1_LOC_156/Y OR2X1_LOC_375/A AND2X1_LOC
XOR2X1_LOC_401 OR2X1_LOC_401/a_8_216# OR2X1_LOC_401/a_36_216# OR2X1_LOC_401/Y VSS VDD
+ OR2X1_LOC_401/A OR2X1_LOC_401/B OR2X1_LOC
XOR2X1_LOC_90 OR2X1_LOC_90/a_8_216# OR2X1_LOC_90/a_36_216# OR2X1_LOC_91/A VSS VDD
+ OR2X1_LOC_54/Y OR2X1_LOC_85/A OR2X1_LOC
XOR2X1_LOC_478 OR2X1_LOC_478/a_8_216# OR2X1_LOC_478/a_36_216# OR2X1_LOC_478/Y VSS VDD
+ OR2X1_LOC_477/Y OR2X1_LOC_469/Y OR2X1_LOC
XOR2X1_LOC_467 OR2X1_LOC_467/a_8_216# OR2X1_LOC_467/a_36_216# OR2X1_LOC_470/A VSS VDD
+ OR2X1_LOC_467/A OR2X1_LOC_467/B OR2X1_LOC
XOR2X1_LOC_423 OR2X1_LOC_423/a_8_216# OR2X1_LOC_423/a_36_216# OR2X1_LOC_423/Y VSS VDD
+ OR2X1_LOC_64/Y OR2X1_LOC_7/A OR2X1_LOC
XAND2X1_LOC_670 AND2X1_LOC_670/a_36_24# OR2X1_LOC_673/B AND2X1_LOC_670/a_8_24# VSS VDD
+ AND2X1_LOC_40/Y OR2X1_LOC_532/B AND2X1_LOC
XAND2X1_LOC_692 AND2X1_LOC_692/a_36_24# OR2X1_LOC_706/B AND2X1_LOC_692/a_8_24# VSS VDD
+ AND2X1_LOC_18/Y AND2X1_LOC_48/A AND2X1_LOC
XAND2X1_LOC_681 AND2X1_LOC_681/a_36_24# OR2X1_LOC_685/B AND2X1_LOC_681/a_8_24# VSS VDD
+ AND2X1_LOC_31/Y OR2X1_LOC_155/A AND2X1_LOC
XOR2X1_LOC_489 OR2X1_LOC_489/a_8_216# OR2X1_LOC_489/a_36_216# OR2X1_LOC_772/B VSS VDD
+ OR2X1_LOC_489/A OR2X1_LOC_489/B OR2X1_LOC
XOR2X1_LOC_456 OR2X1_LOC_456/a_8_216# OR2X1_LOC_456/a_36_216# OR2X1_LOC_456/Y VSS VDD
+ OR2X1_LOC_456/A OR2X1_LOC_190/A OR2X1_LOC
XOR2X1_LOC_445 OR2X1_LOC_445/a_8_216# OR2X1_LOC_445/a_36_216# OR2X1_LOC_455/A VSS VDD
+ OR2X1_LOC_318/B OR2X1_LOC_241/B OR2X1_LOC
XOR2X1_LOC_412 OR2X1_LOC_412/a_8_216# OR2X1_LOC_412/a_36_216# OR2X1_LOC_690/A VSS VDD
+ OR2X1_LOC_44/Y OR2X1_LOC_85/A OR2X1_LOC
XOR2X1_LOC_434 OR2X1_LOC_434/a_8_216# OR2X1_LOC_434/a_36_216# OR2X1_LOC_436/B VSS VDD
+ OR2X1_LOC_434/A OR2X1_LOC_174/A OR2X1_LOC
XAND2X1_LOC_1 AND2X1_LOC_1/a_36_24# AND2X1_LOC_1/Y AND2X1_LOC_1/a_8_24# VSS VDD D_INPUT_6
+ INPUT_7 AND2X1_LOC
XOR2X1_LOC_253 OR2X1_LOC_253/a_8_216# OR2X1_LOC_253/a_36_216# OR2X1_LOC_253/Y VSS VDD
+ OR2X1_LOC_427/A OR2X1_LOC_64/Y OR2X1_LOC
XOR2X1_LOC_242 OR2X1_LOC_242/a_8_216# OR2X1_LOC_242/a_36_216# OR2X1_LOC_244/B VSS VDD
+ OR2X1_LOC_241/Y OR2X1_LOC_506/B OR2X1_LOC
XOR2X1_LOC_231 OR2X1_LOC_231/a_8_216# OR2X1_LOC_231/a_36_216# OR2X1_LOC_641/B VSS VDD
+ OR2X1_LOC_231/A OR2X1_LOC_231/B OR2X1_LOC
XOR2X1_LOC_220 OR2X1_LOC_220/a_8_216# OR2X1_LOC_220/a_36_216# OR2X1_LOC_221/A VSS VDD
+ OR2X1_LOC_220/A OR2X1_LOC_220/B OR2X1_LOC
XOR2X1_LOC_286 OR2X1_LOC_286/a_8_216# OR2X1_LOC_286/a_36_216# OR2X1_LOC_286/Y VSS VDD
+ OR2X1_LOC_285/Y OR2X1_LOC_286/B OR2X1_LOC
XOR2X1_LOC_297 OR2X1_LOC_297/a_8_216# OR2X1_LOC_297/a_36_216# OR2X1_LOC_297/Y VSS VDD
+ OR2X1_LOC_297/A OR2X1_LOC_44/Y OR2X1_LOC
XOR2X1_LOC_264 OR2X1_LOC_264/a_8_216# OR2X1_LOC_264/a_36_216# OR2X1_LOC_264/Y VSS VDD
+ OR2X1_LOC_78/A AND2X1_LOC_41/A OR2X1_LOC
XOR2X1_LOC_275 OR2X1_LOC_275/a_8_216# OR2X1_LOC_275/a_36_216# OR2X1_LOC_275/Y VSS VDD
+ OR2X1_LOC_275/A INPUT_0 OR2X1_LOC
XOR2X1_LOC_819 OR2X1_LOC_819/a_8_216# OR2X1_LOC_819/a_36_216# OR2X1_LOC_820/A VSS VDD
+ OR2X1_LOC_62/A OR2X1_LOC_47/Y OR2X1_LOC
XOR2X1_LOC_808 OR2X1_LOC_808/a_8_216# OR2X1_LOC_808/a_36_216# OR2X1_LOC_811/A VSS VDD
+ OR2X1_LOC_808/A OR2X1_LOC_808/B OR2X1_LOC
XAND2X1_LOC_318 AND2X1_LOC_318/a_36_24# AND2X1_LOC_318/Y AND2X1_LOC_318/a_8_24# VSS VDD
+ OR2X1_LOC_315/Y OR2X1_LOC_316/Y AND2X1_LOC
XAND2X1_LOC_329 AND2X1_LOC_329/a_36_24# OR2X1_LOC_355/B AND2X1_LOC_329/a_8_24# VSS VDD
+ OR2X1_LOC_405/A OR2X1_LOC_596/A AND2X1_LOC
XAND2X1_LOC_307 AND2X1_LOC_307/a_36_24# AND2X1_LOC_307/Y AND2X1_LOC_307/a_8_24# VSS VDD
+ OR2X1_LOC_304/Y OR2X1_LOC_305/Y AND2X1_LOC
XAND2X1_LOC_69 AND2X1_LOC_69/a_36_24# AND2X1_LOC_69/Y AND2X1_LOC_69/a_8_24# VSS VDD
+ AND2X1_LOC_36/Y OR2X1_LOC_68/Y AND2X1_LOC
XAND2X1_LOC_14 AND2X1_LOC_14/a_36_24# OR2X1_LOC_377/A AND2X1_LOC_14/a_8_24# VSS VDD
+ D_INPUT_2 D_INPUT_3 AND2X1_LOC
XAND2X1_LOC_58 AND2X1_LOC_58/a_36_24# OR2X1_LOC_61/B AND2X1_LOC_58/a_8_24# VSS VDD
+ AND2X1_LOC_22/Y OR2X1_LOC_87/A AND2X1_LOC
XAND2X1_LOC_47 AND2X1_LOC_47/a_36_24# AND2X1_LOC_47/Y AND2X1_LOC_47/a_8_24# VSS VDD
+ AND2X1_LOC_25/Y AND2X1_LOC_51/A AND2X1_LOC
XAND2X1_LOC_36 AND2X1_LOC_36/a_36_24# AND2X1_LOC_36/Y AND2X1_LOC_36/a_8_24# VSS VDD
+ AND2X1_LOC_17/Y AND2X1_LOC_21/Y AND2X1_LOC
XAND2X1_LOC_25 AND2X1_LOC_25/a_36_24# AND2X1_LOC_25/Y AND2X1_LOC_25/a_8_24# VSS VDD
+ INPUT_6 D_INPUT_7 AND2X1_LOC
XOR2X1_LOC_638 OR2X1_LOC_638/a_8_216# OR2X1_LOC_638/a_36_216# OR2X1_LOC_651/B VSS VDD
+ OR2X1_LOC_637/Y OR2X1_LOC_638/B OR2X1_LOC
XAND2X1_LOC_852 AND2X1_LOC_852/a_36_24# AND2X1_LOC_852/Y AND2X1_LOC_852/a_8_24# VSS VDD
+ AND2X1_LOC_838/Y AND2X1_LOC_852/B AND2X1_LOC
XAND2X1_LOC_830 AND2X1_LOC_830/a_36_24# AND2X1_LOC_842/B AND2X1_LOC_830/a_8_24# VSS VDD
+ OR2X1_LOC_108/Y OR2X1_LOC_142/Y AND2X1_LOC
XAND2X1_LOC_841 AND2X1_LOC_841/a_36_24# AND2X1_LOC_851/B AND2X1_LOC_841/a_8_24# VSS VDD
+ AND2X1_LOC_831/Y AND2X1_LOC_841/B AND2X1_LOC
XAND2X1_LOC_863 AND2X1_LOC_863/a_36_24# AND2X1_LOC_863/Y AND2X1_LOC_863/a_8_24# VSS VDD
+ AND2X1_LOC_863/A AND2X1_LOC_857/Y AND2X1_LOC
XOR2X1_LOC_616 OR2X1_LOC_616/a_8_216# OR2X1_LOC_616/a_36_216# OR2X1_LOC_616/Y VSS VDD
+ OR2X1_LOC_600/A OR2X1_LOC_18/Y OR2X1_LOC
XOR2X1_LOC_627 OR2X1_LOC_627/a_8_216# OR2X1_LOC_627/a_36_216# OR2X1_LOC_627/Y VSS VDD
+ OR2X1_LOC_36/Y OR2X1_LOC_7/A OR2X1_LOC
XOR2X1_LOC_605 OR2X1_LOC_605/a_8_216# OR2X1_LOC_605/a_36_216# OR2X1_LOC_605/Y VSS VDD
+ OR2X1_LOC_605/A OR2X1_LOC_605/B OR2X1_LOC
XOR2X1_LOC_649 OR2X1_LOC_649/a_8_216# OR2X1_LOC_649/a_36_216# OR2X1_LOC_655/A VSS VDD
+ OR2X1_LOC_643/Y OR2X1_LOC_649/B OR2X1_LOC
XAND2X1_LOC_137 AND2X1_LOC_137/a_36_24# AND2X1_LOC_139/A AND2X1_LOC_137/a_8_24# VSS VDD
+ OR2X1_LOC_132/Y OR2X1_LOC_134/Y AND2X1_LOC
XAND2X1_LOC_126 AND2X1_LOC_126/a_36_24# OR2X1_LOC_160/A AND2X1_LOC_126/a_8_24# VSS VDD
+ OR2X1_LOC_19/B AND2X1_LOC_42/B AND2X1_LOC
XAND2X1_LOC_104 AND2X1_LOC_104/a_36_24# OR2X1_LOC_756/B AND2X1_LOC_104/a_8_24# VSS VDD
+ OR2X1_LOC_19/B AND2X1_LOC_8/Y AND2X1_LOC
XAND2X1_LOC_159 AND2X1_LOC_159/a_36_24# OR2X1_LOC_161/A AND2X1_LOC_159/a_8_24# VSS VDD
+ OR2X1_LOC_68/B OR2X1_LOC_62/B AND2X1_LOC
XAND2X1_LOC_115 AND2X1_LOC_115/a_36_24# AND2X1_LOC_116/B AND2X1_LOC_115/a_8_24# VSS VDD
+ OR2X1_LOC_106/Y AND2X1_LOC_715/A AND2X1_LOC
XAND2X1_LOC_148 AND2X1_LOC_148/a_36_24# AND2X1_LOC_148/Y AND2X1_LOC_148/a_8_24# VSS VDD
+ OR2X1_LOC_145/Y OR2X1_LOC_146/Y AND2X1_LOC
XOR2X1_LOC_424 OR2X1_LOC_424/a_8_216# OR2X1_LOC_424/a_36_216# OR2X1_LOC_424/Y VSS VDD
+ OR2X1_LOC_89/A OR2X1_LOC_44/Y OR2X1_LOC
XOR2X1_LOC_402 OR2X1_LOC_402/a_8_216# OR2X1_LOC_402/a_36_216# OR2X1_LOC_402/Y VSS VDD
+ OR2X1_LOC_401/Y OR2X1_LOC_402/B OR2X1_LOC
XOR2X1_LOC_80 OR2X1_LOC_80/a_8_216# OR2X1_LOC_80/a_36_216# OR2X1_LOC_80/Y VSS VDD
+ OR2X1_LOC_80/A OR2X1_LOC_6/A OR2X1_LOC
XOR2X1_LOC_435 OR2X1_LOC_435/a_8_216# OR2X1_LOC_435/a_36_216# OR2X1_LOC_435/Y VSS VDD
+ OR2X1_LOC_435/A OR2X1_LOC_435/B OR2X1_LOC
XOR2X1_LOC_413 OR2X1_LOC_413/a_8_216# OR2X1_LOC_413/a_36_216# OR2X1_LOC_413/Y VSS VDD
+ OR2X1_LOC_690/A D_INPUT_0 OR2X1_LOC
XOR2X1_LOC_91 OR2X1_LOC_91/a_8_216# OR2X1_LOC_91/a_36_216# OR2X1_LOC_91/Y VSS VDD
+ OR2X1_LOC_91/A OR2X1_LOC_51/Y OR2X1_LOC
XOR2X1_LOC_446 OR2X1_LOC_446/a_8_216# OR2X1_LOC_446/a_36_216# OR2X1_LOC_446/Y VSS VDD
+ OR2X1_LOC_446/A OR2X1_LOC_446/B OR2X1_LOC
XAND2X1_LOC_671 AND2X1_LOC_671/a_36_24# AND2X1_LOC_672/B AND2X1_LOC_671/a_8_24# VSS VDD
+ INPUT_2 OR2X1_LOC_19/B AND2X1_LOC
XAND2X1_LOC_660 AND2X1_LOC_660/a_36_24# AND2X1_LOC_660/Y AND2X1_LOC_660/a_8_24# VSS VDD
+ AND2X1_LOC_660/A AND2X1_LOC_656/Y AND2X1_LOC
XAND2X1_LOC_693 AND2X1_LOC_693/a_36_24# OR2X1_LOC_706/A AND2X1_LOC_693/a_8_24# VSS VDD
+ OR2X1_LOC_377/A AND2X1_LOC_36/Y AND2X1_LOC
XAND2X1_LOC_682 AND2X1_LOC_682/a_36_24# OR2X1_LOC_685/A AND2X1_LOC_682/a_8_24# VSS VDD
+ AND2X1_LOC_36/Y OR2X1_LOC_161/A AND2X1_LOC
XOR2X1_LOC_457 OR2X1_LOC_457/a_8_216# OR2X1_LOC_457/a_36_216# OR2X1_LOC_464/B VSS VDD
+ OR2X1_LOC_787/B OR2X1_LOC_457/B OR2X1_LOC
XOR2X1_LOC_479 OR2X1_LOC_479/a_8_216# OR2X1_LOC_479/a_36_216# OR2X1_LOC_479/Y VSS VDD
+ OR2X1_LOC_476/Y OR2X1_LOC_475/Y OR2X1_LOC
XOR2X1_LOC_468 OR2X1_LOC_468/a_8_216# OR2X1_LOC_468/a_36_216# OR2X1_LOC_468/Y VSS VDD
+ OR2X1_LOC_468/A OR2X1_LOC_436/Y OR2X1_LOC
XAND2X1_LOC_2 AND2X1_LOC_2/a_36_24# AND2X1_LOC_2/Y AND2X1_LOC_2/a_8_24# VSS VDD D_INPUT_4
+ D_INPUT_5 AND2X1_LOC
XOR2X1_LOC_210 OR2X1_LOC_210/a_8_216# OR2X1_LOC_210/a_36_216# OR2X1_LOC_213/A VSS VDD
+ OR2X1_LOC_467/B OR2X1_LOC_210/B OR2X1_LOC
XOR2X1_LOC_232 OR2X1_LOC_232/a_8_216# OR2X1_LOC_232/a_36_216# OR2X1_LOC_232/Y VSS VDD
+ OR2X1_LOC_158/A OR2X1_LOC_16/A OR2X1_LOC
XOR2X1_LOC_254 OR2X1_LOC_254/a_8_216# OR2X1_LOC_254/a_36_216# OR2X1_LOC_456/A VSS VDD
+ OR2X1_LOC_254/A OR2X1_LOC_254/B OR2X1_LOC
XOR2X1_LOC_243 OR2X1_LOC_243/a_8_216# OR2X1_LOC_243/a_36_216# OR2X1_LOC_244/A VSS VDD
+ OR2X1_LOC_243/A OR2X1_LOC_243/B OR2X1_LOC
XOR2X1_LOC_276 OR2X1_LOC_276/a_8_216# OR2X1_LOC_276/a_36_216# OR2X1_LOC_473/A VSS VDD
+ OR2X1_LOC_276/A OR2X1_LOC_276/B OR2X1_LOC
XOR2X1_LOC_265 OR2X1_LOC_265/a_8_216# OR2X1_LOC_265/a_36_216# OR2X1_LOC_265/Y VSS VDD
+ OR2X1_LOC_517/A OR2X1_LOC_40/Y OR2X1_LOC
XOR2X1_LOC_221 OR2X1_LOC_221/a_8_216# OR2X1_LOC_221/a_36_216# OR2X1_LOC_223/B VSS VDD
+ OR2X1_LOC_221/A OR2X1_LOC_739/B OR2X1_LOC
XAND2X1_LOC_490 AND2X1_LOC_490/a_36_24# OR2X1_LOC_557/A AND2X1_LOC_490/a_8_24# VSS VDD
+ OR2X1_LOC_6/B AND2X1_LOC_86/B AND2X1_LOC
XOR2X1_LOC_287 OR2X1_LOC_287/a_8_216# OR2X1_LOC_287/a_36_216# OR2X1_LOC_288/A VSS VDD
+ OR2X1_LOC_287/A OR2X1_LOC_287/B OR2X1_LOC
XOR2X1_LOC_298 OR2X1_LOC_298/a_8_216# OR2X1_LOC_298/a_36_216# OR2X1_LOC_298/Y VSS VDD
+ OR2X1_LOC_56/A OR2X1_LOC_31/Y OR2X1_LOC
XOR2X1_LOC_809 OR2X1_LOC_809/a_8_216# OR2X1_LOC_809/a_36_216# OR2X1_LOC_810/A VSS VDD
+ OR2X1_LOC_802/Y OR2X1_LOC_809/B OR2X1_LOC
XAND2X1_LOC_308 AND2X1_LOC_308/a_36_24# AND2X1_LOC_727/A AND2X1_LOC_308/a_8_24# VSS VDD
+ OR2X1_LOC_306/Y AND2X1_LOC_307/Y AND2X1_LOC
XAND2X1_LOC_319 AND2X1_LOC_319/a_36_24# AND2X1_LOC_798/A AND2X1_LOC_319/a_8_24# VSS VDD
+ AND2X1_LOC_319/A AND2X1_LOC_318/Y AND2X1_LOC
XOR2X1_LOC_1 OR2X1_LOC_1/a_8_216# OR2X1_LOC_1/a_36_216# OR2X1_LOC_3/B VSS VDD D_INPUT_7
+ INPUT_6 OR2X1_LOC
XAND2X1_LOC_37 AND2X1_LOC_37/a_36_24# AND2X1_LOC_42/B AND2X1_LOC_37/a_8_24# VSS VDD
+ INPUT_2 INPUT_3 AND2X1_LOC
XAND2X1_LOC_15 AND2X1_LOC_15/a_36_24# OR2X1_LOC_78/B AND2X1_LOC_15/a_8_24# VSS VDD
+ OR2X1_LOC_62/B OR2X1_LOC_377/A AND2X1_LOC
XAND2X1_LOC_48 AND2X1_LOC_48/a_36_24# AND2X1_LOC_48/Y AND2X1_LOC_48/a_8_24# VSS VDD
+ AND2X1_LOC_48/A AND2X1_LOC_47/Y AND2X1_LOC
XAND2X1_LOC_59 AND2X1_LOC_59/a_36_24# AND2X1_LOC_59/Y AND2X1_LOC_59/a_8_24# VSS VDD
+ AND2X1_LOC_11/Y AND2X1_LOC_25/Y AND2X1_LOC
XAND2X1_LOC_26 AND2X1_LOC_26/a_36_24# OR2X1_LOC_66/A AND2X1_LOC_26/a_8_24# VSS VDD
+ AND2X1_LOC_21/Y AND2X1_LOC_25/Y AND2X1_LOC
XOR2X1_LOC_617 OR2X1_LOC_617/a_8_216# OR2X1_LOC_617/a_36_216# OR2X1_LOC_617/Y VSS VDD
+ OR2X1_LOC_51/Y OR2X1_LOC_39/A OR2X1_LOC
XOR2X1_LOC_606 OR2X1_LOC_606/a_8_216# OR2X1_LOC_606/a_36_216# OR2X1_LOC_606/Y VSS VDD
+ OR2X1_LOC_121/B OR2X1_LOC_532/B OR2X1_LOC
XOR2X1_LOC_639 OR2X1_LOC_639/a_8_216# OR2X1_LOC_639/a_36_216# OR2X1_LOC_651/A VSS VDD
+ OR2X1_LOC_639/A OR2X1_LOC_639/B OR2X1_LOC
XAND2X1_LOC_842 AND2X1_LOC_842/a_36_24# AND2X1_LOC_850/A AND2X1_LOC_842/a_8_24# VSS VDD
+ OR2X1_LOC_184/Y AND2X1_LOC_842/B AND2X1_LOC
XAND2X1_LOC_820 AND2X1_LOC_820/a_36_24# OR2X1_LOC_847/A AND2X1_LOC_820/a_8_24# VSS VDD
+ OR2X1_LOC_818/Y AND2X1_LOC_820/B AND2X1_LOC
XAND2X1_LOC_831 AND2X1_LOC_831/a_36_24# AND2X1_LOC_831/Y AND2X1_LOC_831/a_8_24# VSS VDD
+ OR2X1_LOC_273/Y OR2X1_LOC_300/Y AND2X1_LOC
XAND2X1_LOC_853 AND2X1_LOC_853/a_36_24# AND2X1_LOC_853/Y AND2X1_LOC_853/a_8_24# VSS VDD
+ AND2X1_LOC_35/Y AND2X1_LOC_211/B AND2X1_LOC
XAND2X1_LOC_864 AND2X1_LOC_864/a_36_24# AND2X1_LOC_866/A AND2X1_LOC_864/a_8_24# VSS VDD
+ AND2X1_LOC_810/A AND2X1_LOC_863/Y AND2X1_LOC
XOR2X1_LOC_628 OR2X1_LOC_628/a_8_216# OR2X1_LOC_628/a_36_216# OR2X1_LOC_628/Y VSS VDD
+ OR2X1_LOC_92/Y OR2X1_LOC_47/Y OR2X1_LOC
XAND2X1_LOC_105 AND2X1_LOC_105/a_36_24# OR2X1_LOC_106/A AND2X1_LOC_105/a_8_24# VSS VDD
+ OR2X1_LOC_89/A OR2X1_LOC_600/A AND2X1_LOC
XAND2X1_LOC_127 AND2X1_LOC_127/a_36_24# OR2X1_LOC_128/A AND2X1_LOC_127/a_8_24# VSS VDD
+ AND2X1_LOC_3/Y OR2X1_LOC_160/A AND2X1_LOC
XAND2X1_LOC_116 AND2X1_LOC_116/a_36_24# AND2X1_LOC_116/Y AND2X1_LOC_116/a_8_24# VSS VDD
+ AND2X1_LOC_114/Y AND2X1_LOC_116/B AND2X1_LOC
XAND2X1_LOC_138 AND2X1_LOC_138/a_36_24# AND2X1_LOC_139/B AND2X1_LOC_138/a_8_24# VSS VDD
+ OR2X1_LOC_135/Y OR2X1_LOC_136/Y AND2X1_LOC
XAND2X1_LOC_149 AND2X1_LOC_149/a_36_24# AND2X1_LOC_797/A AND2X1_LOC_149/a_8_24# VSS VDD
+ AND2X1_LOC_147/Y AND2X1_LOC_148/Y AND2X1_LOC
XOR2X1_LOC_70 OR2X1_LOC_70/a_8_216# OR2X1_LOC_70/a_36_216# OR2X1_LOC_70/Y VSS VDD
+ OR2X1_LOC_70/A OR2X1_LOC_2/Y OR2X1_LOC
XOR2X1_LOC_425 OR2X1_LOC_425/a_8_216# OR2X1_LOC_425/a_36_216# OR2X1_LOC_426/A VSS VDD
+ OR2X1_LOC_17/Y INPUT_5 OR2X1_LOC
XOR2X1_LOC_447 OR2X1_LOC_447/a_8_216# OR2X1_LOC_447/a_36_216# OR2X1_LOC_447/Y VSS VDD
+ OR2X1_LOC_447/A OR2X1_LOC_506/A OR2X1_LOC
XOR2X1_LOC_469 OR2X1_LOC_469/a_8_216# OR2X1_LOC_469/a_36_216# OR2X1_LOC_469/Y VSS VDD
+ OR2X1_LOC_468/Y OR2X1_LOC_469/B OR2X1_LOC
XAND2X1_LOC_650 AND2X1_LOC_650/a_36_24# AND2X1_LOC_650/Y AND2X1_LOC_650/a_8_24# VSS VDD
+ AND2X1_LOC_640/Y AND2X1_LOC_641/Y AND2X1_LOC
XOR2X1_LOC_403 OR2X1_LOC_403/a_8_216# OR2X1_LOC_403/a_36_216# OR2X1_LOC_404/A VSS VDD
+ OR2X1_LOC_403/A OR2X1_LOC_403/B OR2X1_LOC
XOR2X1_LOC_92 OR2X1_LOC_92/a_8_216# OR2X1_LOC_92/a_36_216# OR2X1_LOC_92/Y VSS VDD
+ OR2X1_LOC_8/Y D_INPUT_1 OR2X1_LOC
XOR2X1_LOC_458 OR2X1_LOC_458/a_8_216# OR2X1_LOC_458/a_36_216# OR2X1_LOC_464/A VSS VDD
+ OR2X1_LOC_374/Y OR2X1_LOC_458/B OR2X1_LOC
XOR2X1_LOC_414 OR2X1_LOC_414/a_8_216# OR2X1_LOC_414/a_36_216# OR2X1_LOC_414/Y VSS VDD
+ OR2X1_LOC_6/B D_INPUT_3 OR2X1_LOC
XOR2X1_LOC_81 OR2X1_LOC_81/a_8_216# OR2X1_LOC_81/a_36_216# OR2X1_LOC_81/Y VSS VDD
+ OR2X1_LOC_80/Y OR2X1_LOC_59/Y OR2X1_LOC
XOR2X1_LOC_436 OR2X1_LOC_436/a_8_216# OR2X1_LOC_436/a_36_216# OR2X1_LOC_436/Y VSS VDD
+ OR2X1_LOC_435/Y OR2X1_LOC_436/B OR2X1_LOC
XAND2X1_LOC_672 AND2X1_LOC_672/a_36_24# OR2X1_LOC_673/A AND2X1_LOC_672/a_8_24# VSS VDD
+ OR2X1_LOC_375/A AND2X1_LOC_672/B AND2X1_LOC
XAND2X1_LOC_661 AND2X1_LOC_661/a_36_24# AND2X1_LOC_662/B AND2X1_LOC_661/a_8_24# VSS VDD
+ AND2X1_LOC_661/A AND2X1_LOC_654/Y AND2X1_LOC
XAND2X1_LOC_683 AND2X1_LOC_683/a_36_24# OR2X1_LOC_686/B AND2X1_LOC_683/a_8_24# VSS VDD
+ OR2X1_LOC_78/B AND2X1_LOC_22/Y AND2X1_LOC
XAND2X1_LOC_694 AND2X1_LOC_694/a_36_24# OR2X1_LOC_707/B AND2X1_LOC_694/a_8_24# VSS VDD
+ OR2X1_LOC_161/B AND2X1_LOC_425/Y AND2X1_LOC
XAND2X1_LOC_3 AND2X1_LOC_3/a_36_24# AND2X1_LOC_3/Y AND2X1_LOC_3/a_8_24# VSS VDD AND2X1_LOC_1/Y
+ AND2X1_LOC_2/Y AND2X1_LOC
XOR2X1_LOC_200 OR2X1_LOC_200/a_8_216# OR2X1_LOC_200/a_36_216# OR2X1_LOC_200/Y VSS VDD
+ OR2X1_LOC_194/Y OR2X1_LOC_193/Y OR2X1_LOC
XAND2X1_LOC_491 AND2X1_LOC_491/a_36_24# OR2X1_LOC_493/B AND2X1_LOC_491/a_8_24# VSS VDD
+ AND2X1_LOC_31/Y OR2X1_LOC_532/B AND2X1_LOC
XAND2X1_LOC_480 AND2X1_LOC_480/a_36_24# GATE_479 AND2X1_LOC_480/a_8_24# VSS VDD
+ AND2X1_LOC_480/A AND2X1_LOC_479/Y AND2X1_LOC
XOR2X1_LOC_288 OR2X1_LOC_288/a_8_216# OR2X1_LOC_288/a_36_216# OR2X1_LOC_362/B VSS VDD
+ OR2X1_LOC_288/A OR2X1_LOC_286/Y OR2X1_LOC
XOR2X1_LOC_233 OR2X1_LOC_233/a_8_216# OR2X1_LOC_233/a_36_216# OR2X1_LOC_291/A VSS VDD
+ OR2X1_LOC_46/A D_INPUT_0 OR2X1_LOC
XOR2X1_LOC_255 OR2X1_LOC_255/a_8_216# OR2X1_LOC_255/a_36_216# OR2X1_LOC_256/A VSS VDD
+ OR2X1_LOC_158/A OR2X1_LOC_85/A OR2X1_LOC
XOR2X1_LOC_244 OR2X1_LOC_244/a_8_216# OR2X1_LOC_244/a_36_216# OR2X1_LOC_244/Y VSS VDD
+ OR2X1_LOC_244/A OR2X1_LOC_244/B OR2X1_LOC
XOR2X1_LOC_266 OR2X1_LOC_266/a_8_216# OR2X1_LOC_266/a_36_216# OR2X1_LOC_267/A VSS VDD
+ OR2X1_LOC_266/A OR2X1_LOC_786/A OR2X1_LOC
XOR2X1_LOC_277 OR2X1_LOC_277/a_8_216# OR2X1_LOC_277/a_36_216# OR2X1_LOC_278/A VSS VDD
+ OR2X1_LOC_47/Y OR2X1_LOC_85/A OR2X1_LOC
XOR2X1_LOC_222 OR2X1_LOC_222/a_8_216# OR2X1_LOC_222/a_36_216# OR2X1_LOC_223/A VSS VDD
+ OR2X1_LOC_222/A OR2X1_LOC_218/Y OR2X1_LOC
XOR2X1_LOC_211 OR2X1_LOC_211/a_8_216# OR2X1_LOC_211/a_36_216# OR2X1_LOC_212/A VSS VDD
+ OR2X1_LOC_175/Y OR2X1_LOC_170/Y OR2X1_LOC
XOR2X1_LOC_299 OR2X1_LOC_299/a_8_216# OR2X1_LOC_299/a_36_216# OR2X1_LOC_299/Y VSS VDD
+ OR2X1_LOC_426/B OR2X1_LOC_12/Y OR2X1_LOC
XAND2X1_LOC_309 AND2X1_LOC_309/a_36_24# OR2X1_LOC_335/B AND2X1_LOC_309/a_8_24# VSS VDD
+ AND2X1_LOC_22/Y OR2X1_LOC_814/A AND2X1_LOC
XOR2X1_LOC_2 OR2X1_LOC_2/a_8_216# OR2X1_LOC_2/a_36_216# OR2X1_LOC_2/Y VSS VDD INPUT_5
+ INPUT_4 OR2X1_LOC
XAND2X1_LOC_16 AND2X1_LOC_16/a_36_24# OR2X1_LOC_194/B AND2X1_LOC_16/a_8_24# VSS VDD
+ AND2X1_LOC_3/Y OR2X1_LOC_78/B AND2X1_LOC
XAND2X1_LOC_49 AND2X1_LOC_49/a_36_24# OR2X1_LOC_87/A AND2X1_LOC_49/a_8_24# VSS VDD
+ OR2X1_LOC_377/A OR2X1_LOC_80/A AND2X1_LOC
XAND2X1_LOC_38 AND2X1_LOC_38/a_36_24# OR2X1_LOC_154/A AND2X1_LOC_38/a_8_24# VSS VDD
+ OR2X1_LOC_80/A AND2X1_LOC_42/B AND2X1_LOC
XAND2X1_LOC_27 AND2X1_LOC_27/a_36_24# OR2X1_LOC_34/B AND2X1_LOC_27/a_8_24# VSS VDD
+ AND2X1_LOC_7/B OR2X1_LOC_66/A AND2X1_LOC
XAND2X1_LOC_821 AND2X1_LOC_821/a_36_24# OR2X1_LOC_835/B AND2X1_LOC_821/a_8_24# VSS VDD
+ AND2X1_LOC_41/A AND2X1_LOC_70/Y AND2X1_LOC
XAND2X1_LOC_810 AND2X1_LOC_810/a_36_24# AND2X1_LOC_810/Y AND2X1_LOC_810/a_8_24# VSS VDD
+ AND2X1_LOC_810/A AND2X1_LOC_810/B AND2X1_LOC
XAND2X1_LOC_832 AND2X1_LOC_832/a_36_24# AND2X1_LOC_841/B AND2X1_LOC_832/a_8_24# VSS VDD
+ OR2X1_LOC_423/Y OR2X1_LOC_433/Y AND2X1_LOC
XOR2X1_LOC_618 OR2X1_LOC_618/a_8_216# OR2X1_LOC_618/a_36_216# OR2X1_LOC_618/Y VSS VDD
+ OR2X1_LOC_49/A INPUT_3 OR2X1_LOC
XOR2X1_LOC_629 OR2X1_LOC_629/a_8_216# OR2X1_LOC_629/a_36_216# OR2X1_LOC_629/Y VSS VDD
+ OR2X1_LOC_629/A OR2X1_LOC_629/B OR2X1_LOC
XOR2X1_LOC_607 OR2X1_LOC_607/a_8_216# OR2X1_LOC_607/a_36_216# OR2X1_LOC_607/Y VSS VDD
+ OR2X1_LOC_607/A OR2X1_LOC_18/Y OR2X1_LOC
XAND2X1_LOC_865 AND2X1_LOC_865/a_36_24# AND2X1_LOC_866/B AND2X1_LOC_865/a_8_24# VSS VDD
+ AND2X1_LOC_865/A AND2X1_LOC_862/Y AND2X1_LOC
XAND2X1_LOC_843 AND2X1_LOC_843/a_36_24# AND2X1_LOC_843/Y AND2X1_LOC_843/a_8_24# VSS VDD
+ OR2X1_LOC_251/Y OR2X1_LOC_278/Y AND2X1_LOC
XAND2X1_LOC_854 AND2X1_LOC_854/a_36_24# AND2X1_LOC_856/A AND2X1_LOC_854/a_8_24# VSS VDD
+ AND2X1_LOC_354/B AND2X1_LOC_535/Y AND2X1_LOC
XAND2X1_LOC_117 AND2X1_LOC_117/a_36_24# OR2X1_LOC_123/B AND2X1_LOC_117/a_8_24# VSS VDD
+ AND2X1_LOC_65/A AND2X1_LOC_70/Y AND2X1_LOC
XAND2X1_LOC_128 AND2X1_LOC_128/a_36_24# AND2X1_LOC_554/B AND2X1_LOC_128/a_8_24# VSS VDD
+ OR2X1_LOC_125/Y OR2X1_LOC_127/Y AND2X1_LOC
XAND2X1_LOC_106 AND2X1_LOC_106/a_36_24# OR2X1_LOC_115/B AND2X1_LOC_106/a_8_24# VSS VDD
+ AND2X1_LOC_47/Y OR2X1_LOC_105/Y AND2X1_LOC
XAND2X1_LOC_139 AND2X1_LOC_139/a_36_24# AND2X1_LOC_141/A AND2X1_LOC_139/a_8_24# VSS VDD
+ AND2X1_LOC_139/A AND2X1_LOC_139/B AND2X1_LOC
XOR2X1_LOC_71 OR2X1_LOC_71/a_8_216# OR2X1_LOC_71/a_36_216# OR2X1_LOC_71/Y VSS VDD
+ OR2X1_LOC_71/A OR2X1_LOC_6/A OR2X1_LOC
XOR2X1_LOC_82 OR2X1_LOC_82/a_8_216# OR2X1_LOC_82/a_36_216# OR2X1_LOC_83/A VSS VDD
+ OR2X1_LOC_80/A OR2X1_LOC_46/A OR2X1_LOC
XOR2X1_LOC_60 OR2X1_LOC_60/a_8_216# OR2X1_LOC_60/a_36_216# OR2X1_LOC_60/Y VSS VDD
+ OR2X1_LOC_59/Y OR2X1_LOC_39/A OR2X1_LOC
XOR2X1_LOC_426 OR2X1_LOC_426/a_8_216# OR2X1_LOC_426/a_36_216# OR2X1_LOC_426/Y VSS VDD
+ OR2X1_LOC_426/A OR2X1_LOC_426/B OR2X1_LOC
XOR2X1_LOC_448 OR2X1_LOC_448/a_8_216# OR2X1_LOC_448/a_36_216# OR2X1_LOC_448/Y VSS VDD
+ OR2X1_LOC_448/A OR2X1_LOC_448/B OR2X1_LOC
XOR2X1_LOC_459 OR2X1_LOC_459/a_8_216# OR2X1_LOC_459/a_36_216# OR2X1_LOC_463/B VSS VDD
+ OR2X1_LOC_459/A OR2X1_LOC_459/B OR2X1_LOC
XAND2X1_LOC_673 AND2X1_LOC_673/a_36_24# AND2X1_LOC_721/A AND2X1_LOC_673/a_8_24# VSS VDD
+ OR2X1_LOC_670/Y OR2X1_LOC_672/Y AND2X1_LOC
XAND2X1_LOC_662 AND2X1_LOC_662/a_36_24# AND2X1_LOC_663/B AND2X1_LOC_662/a_8_24# VSS VDD
+ AND2X1_LOC_660/Y AND2X1_LOC_662/B AND2X1_LOC
XAND2X1_LOC_640 AND2X1_LOC_640/a_36_24# AND2X1_LOC_640/Y AND2X1_LOC_640/a_8_24# VSS VDD
+ AND2X1_LOC_633/Y AND2X1_LOC_634/Y AND2X1_LOC
XAND2X1_LOC_684 AND2X1_LOC_684/a_36_24# OR2X1_LOC_686/A AND2X1_LOC_684/a_8_24# VSS VDD
+ AND2X1_LOC_12/Y AND2X1_LOC_43/B AND2X1_LOC
XAND2X1_LOC_651 AND2X1_LOC_651/a_36_24# AND2X1_LOC_654/B AND2X1_LOC_651/a_8_24# VSS VDD
+ AND2X1_LOC_638/Y AND2X1_LOC_651/B AND2X1_LOC
XOR2X1_LOC_404 OR2X1_LOC_404/a_8_216# OR2X1_LOC_404/a_36_216# OR2X1_LOC_404/Y VSS VDD
+ OR2X1_LOC_404/A OR2X1_LOC_402/Y OR2X1_LOC
XOR2X1_LOC_93 OR2X1_LOC_93/a_8_216# OR2X1_LOC_93/a_36_216# OR2X1_LOC_93/Y VSS VDD
+ OR2X1_LOC_92/Y OR2X1_LOC_26/Y OR2X1_LOC
XOR2X1_LOC_415 OR2X1_LOC_415/a_8_216# OR2X1_LOC_415/a_36_216# OR2X1_LOC_415/Y VSS VDD
+ OR2X1_LOC_415/A OR2X1_LOC_598/A OR2X1_LOC
XOR2X1_LOC_437 OR2X1_LOC_437/a_8_216# OR2X1_LOC_437/a_36_216# OR2X1_LOC_437/Y VSS VDD
+ OR2X1_LOC_437/A OR2X1_LOC_59/Y OR2X1_LOC
XAND2X1_LOC_695 AND2X1_LOC_695/a_36_24# OR2X1_LOC_707/A AND2X1_LOC_695/a_8_24# VSS VDD
+ OR2X1_LOC_160/B AND2X1_LOC_47/Y AND2X1_LOC
XAND2X1_LOC_4 AND2X1_LOC_4/a_36_24# OR2X1_LOC_19/B AND2X1_LOC_4/a_8_24# VSS VDD INPUT_0
+ D_INPUT_1 AND2X1_LOC
XOR2X1_LOC_201 OR2X1_LOC_201/a_8_216# OR2X1_LOC_201/a_36_216# OR2X1_LOC_201/Y VSS VDD
+ OR2X1_LOC_201/A OR2X1_LOC_61/Y OR2X1_LOC
XAND2X1_LOC_492 AND2X1_LOC_492/a_36_24# OR2X1_LOC_493/A AND2X1_LOC_492/a_8_24# VSS VDD
+ AND2X1_LOC_59/Y OR2X1_LOC_160/A AND2X1_LOC
XAND2X1_LOC_481 AND2X1_LOC_481/a_36_24# OR2X1_LOC_555/A AND2X1_LOC_481/a_8_24# VSS VDD
+ AND2X1_LOC_3/Y OR2X1_LOC_294/Y AND2X1_LOC
XAND2X1_LOC_470 AND2X1_LOC_470/a_36_24# AND2X1_LOC_477/A AND2X1_LOC_470/a_8_24# VSS VDD
+ AND2X1_LOC_470/A AND2X1_LOC_470/B AND2X1_LOC
XOR2X1_LOC_234 OR2X1_LOC_234/a_8_216# OR2X1_LOC_234/a_36_216# OR2X1_LOC_234/Y VSS VDD
+ OR2X1_LOC_291/A OR2X1_LOC_47/Y OR2X1_LOC
XOR2X1_LOC_256 OR2X1_LOC_256/a_8_216# OR2X1_LOC_256/a_36_216# OR2X1_LOC_256/Y VSS VDD
+ OR2X1_LOC_256/A OR2X1_LOC_19/B OR2X1_LOC
XOR2X1_LOC_267 OR2X1_LOC_267/a_8_216# OR2X1_LOC_267/a_36_216# OR2X1_LOC_267/Y VSS VDD
+ OR2X1_LOC_267/A OR2X1_LOC_641/A OR2X1_LOC
XOR2X1_LOC_278 OR2X1_LOC_278/a_8_216# OR2X1_LOC_278/a_36_216# OR2X1_LOC_278/Y VSS VDD
+ OR2X1_LOC_278/A OR2X1_LOC_62/B OR2X1_LOC
XOR2X1_LOC_245 OR2X1_LOC_245/a_8_216# OR2X1_LOC_245/a_36_216# OR2X1_LOC_246/A VSS VDD
+ OR2X1_LOC_85/A OR2X1_LOC_26/Y OR2X1_LOC
XOR2X1_LOC_223 OR2X1_LOC_223/a_8_216# OR2X1_LOC_223/a_36_216# D_GATE_222 VSS VDD
+ OR2X1_LOC_223/A OR2X1_LOC_223/B OR2X1_LOC
XOR2X1_LOC_289 OR2X1_LOC_289/a_8_216# OR2X1_LOC_289/a_36_216# OR2X1_LOC_289/Y VSS VDD
+ OR2X1_LOC_417/A OR2X1_LOC_51/Y OR2X1_LOC
XOR2X1_LOC_212 OR2X1_LOC_212/a_8_216# OR2X1_LOC_212/a_36_216# OR2X1_LOC_220/B VSS VDD
+ OR2X1_LOC_212/A OR2X1_LOC_212/B OR2X1_LOC
XOR2X1_LOC_790 OR2X1_LOC_790/a_8_216# OR2X1_LOC_790/a_36_216# OR2X1_LOC_793/A VSS VDD
+ OR2X1_LOC_790/A OR2X1_LOC_790/B OR2X1_LOC
XOR2X1_LOC_3 OR2X1_LOC_3/a_8_216# OR2X1_LOC_3/a_36_216# OR2X1_LOC_3/Y VSS VDD OR2X1_LOC_2/Y
+ OR2X1_LOC_3/B OR2X1_LOC
XAND2X1_LOC_28 AND2X1_LOC_28/a_36_24# OR2X1_LOC_80/A AND2X1_LOC_28/a_8_24# VSS VDD
+ D_INPUT_0 INPUT_1 AND2X1_LOC
XAND2X1_LOC_39 AND2X1_LOC_39/a_36_24# AND2X1_LOC_39/Y AND2X1_LOC_39/a_8_24# VSS VDD
+ AND2X1_LOC_36/Y OR2X1_LOC_154/A AND2X1_LOC
XAND2X1_LOC_17 AND2X1_LOC_17/a_36_24# AND2X1_LOC_17/Y AND2X1_LOC_17/a_8_24# VSS VDD
+ INPUT_6 INPUT_7 AND2X1_LOC
XAND2X1_LOC_844 AND2X1_LOC_844/a_36_24# AND2X1_LOC_849/A AND2X1_LOC_844/a_8_24# VSS VDD
+ OR2X1_LOC_497/Y AND2X1_LOC_523/Y AND2X1_LOC
XAND2X1_LOC_866 AND2X1_LOC_866/a_36_24# GATE_865 AND2X1_LOC_866/a_8_24# VSS VDD
+ AND2X1_LOC_866/A AND2X1_LOC_866/B AND2X1_LOC
XAND2X1_LOC_833 AND2X1_LOC_833/a_36_24# AND2X1_LOC_840/A AND2X1_LOC_833/a_8_24# VSS VDD
+ OR2X1_LOC_482/Y OR2X1_LOC_495/Y AND2X1_LOC
XAND2X1_LOC_811 AND2X1_LOC_811/a_36_24# AND2X1_LOC_811/Y AND2X1_LOC_811/a_8_24# VSS VDD
+ AND2X1_LOC_807/Y AND2X1_LOC_811/B AND2X1_LOC
XAND2X1_LOC_822 AND2X1_LOC_822/a_36_24# OR2X1_LOC_835/A AND2X1_LOC_822/a_8_24# VSS VDD
+ AND2X1_LOC_64/Y OR2X1_LOC_532/B AND2X1_LOC
XAND2X1_LOC_855 AND2X1_LOC_855/a_36_24# AND2X1_LOC_856/B AND2X1_LOC_855/a_8_24# VSS VDD
+ AND2X1_LOC_729/B OR2X1_LOC_829/Y AND2X1_LOC
XAND2X1_LOC_800 AND2X1_LOC_800/a_36_24# AND2X1_LOC_801/B AND2X1_LOC_800/a_8_24# VSS VDD
+ AND2X1_LOC_687/Y OR2X1_LOC_760/Y AND2X1_LOC
XOR2X1_LOC_619 OR2X1_LOC_619/a_8_216# OR2X1_LOC_619/a_36_216# OR2X1_LOC_619/Y VSS VDD
+ OR2X1_LOC_618/Y OR2X1_LOC_36/Y OR2X1_LOC
XOR2X1_LOC_608 OR2X1_LOC_608/a_8_216# OR2X1_LOC_608/a_36_216# OR2X1_LOC_608/Y VSS VDD
+ OR2X1_LOC_185/A OR2X1_LOC_78/B OR2X1_LOC
XAND2X1_LOC_129 AND2X1_LOC_129/a_36_24# OR2X1_LOC_130/A AND2X1_LOC_129/a_8_24# VSS VDD
+ OR2X1_LOC_49/A AND2X1_LOC_42/B AND2X1_LOC
XAND2X1_LOC_118 AND2X1_LOC_118/a_36_24# OR2X1_LOC_633/B AND2X1_LOC_118/a_8_24# VSS VDD
+ AND2X1_LOC_70/Y OR2X1_LOC_78/A AND2X1_LOC
XAND2X1_LOC_107 AND2X1_LOC_107/a_36_24# OR2X1_LOC_113/A AND2X1_LOC_107/a_8_24# VSS VDD
+ AND2X1_LOC_64/Y OR2X1_LOC_78/A AND2X1_LOC
XOR2X1_LOC_50 OR2X1_LOC_50/a_8_216# OR2X1_LOC_50/a_36_216# OR2X1_LOC_70/A VSS VDD
+ INPUT_7 INPUT_6 OR2X1_LOC
XOR2X1_LOC_94 OR2X1_LOC_94/a_8_216# OR2X1_LOC_94/a_36_216# OR2X1_LOC_96/B VSS VDD
+ OR2X1_LOC_62/A OR2X1_LOC_46/A OR2X1_LOC
XOR2X1_LOC_83 OR2X1_LOC_83/a_8_216# OR2X1_LOC_83/a_36_216# OR2X1_LOC_83/Y VSS VDD
+ OR2X1_LOC_83/A OR2X1_LOC_26/Y OR2X1_LOC
XOR2X1_LOC_72 OR2X1_LOC_72/a_8_216# OR2X1_LOC_72/a_36_216# OR2X1_LOC_72/Y VSS VDD
+ OR2X1_LOC_71/Y OR2X1_LOC_70/Y OR2X1_LOC
XOR2X1_LOC_61 OR2X1_LOC_61/a_8_216# OR2X1_LOC_61/a_36_216# OR2X1_LOC_61/Y VSS VDD
+ OR2X1_LOC_61/A OR2X1_LOC_61/B OR2X1_LOC
XOR2X1_LOC_427 OR2X1_LOC_427/a_8_216# OR2X1_LOC_427/a_36_216# OR2X1_LOC_427/Y VSS VDD
+ OR2X1_LOC_427/A OR2X1_LOC_70/Y OR2X1_LOC
XOR2X1_LOC_449 OR2X1_LOC_449/a_8_216# OR2X1_LOC_449/a_36_216# OR2X1_LOC_453/A VSS VDD
+ OR2X1_LOC_449/A OR2X1_LOC_449/B OR2X1_LOC
XAND2X1_LOC_674 AND2X1_LOC_674/a_36_24# OR2X1_LOC_675/A AND2X1_LOC_674/a_8_24# VSS VDD
+ AND2X1_LOC_70/Y OR2X1_LOC_405/A AND2X1_LOC
XAND2X1_LOC_630 AND2X1_LOC_630/a_36_24# AND2X1_LOC_632/A AND2X1_LOC_630/a_8_24# VSS VDD
+ OR2X1_LOC_628/Y AND2X1_LOC_629/Y AND2X1_LOC
XAND2X1_LOC_663 AND2X1_LOC_663/a_36_24# GATE_662 AND2X1_LOC_663/a_8_24# VSS VDD
+ AND2X1_LOC_663/A AND2X1_LOC_663/B AND2X1_LOC
XAND2X1_LOC_641 AND2X1_LOC_641/a_36_24# AND2X1_LOC_641/Y AND2X1_LOC_641/a_8_24# VSS VDD
+ AND2X1_LOC_231/Y OR2X1_LOC_265/Y AND2X1_LOC
XAND2X1_LOC_652 AND2X1_LOC_652/a_36_24# AND2X1_LOC_653/B AND2X1_LOC_652/a_8_24# VSS VDD
+ AND2X1_LOC_468/B AND2X1_LOC_593/Y AND2X1_LOC
XAND2X1_LOC_696 AND2X1_LOC_696/a_36_24# OR2X1_LOC_708/B AND2X1_LOC_696/a_8_24# VSS VDD
+ OR2X1_LOC_66/A OR2X1_LOC_502/A AND2X1_LOC
XAND2X1_LOC_685 AND2X1_LOC_685/a_36_24# AND2X1_LOC_687/A AND2X1_LOC_685/a_8_24# VSS VDD
+ OR2X1_LOC_681/Y OR2X1_LOC_682/Y AND2X1_LOC
XOR2X1_LOC_416 OR2X1_LOC_416/a_8_216# OR2X1_LOC_416/a_36_216# OR2X1_LOC_416/Y VSS VDD
+ OR2X1_LOC_416/A OR2X1_LOC_158/A OR2X1_LOC
XOR2X1_LOC_405 OR2X1_LOC_405/a_8_216# OR2X1_LOC_405/a_36_216# OR2X1_LOC_405/Y VSS VDD
+ OR2X1_LOC_405/A AND2X1_LOC_48/A OR2X1_LOC
XOR2X1_LOC_438 OR2X1_LOC_438/a_8_216# OR2X1_LOC_438/a_36_216# OR2X1_LOC_438/Y VSS VDD
+ OR2X1_LOC_70/Y OR2X1_LOC_45/B OR2X1_LOC
XAND2X1_LOC_5 AND2X1_LOC_5/a_36_24# OR2X1_LOC_68/B AND2X1_LOC_5/a_8_24# VSS VDD D_INPUT_2
+ INPUT_3 AND2X1_LOC
XOR2X1_LOC_213 OR2X1_LOC_213/a_8_216# OR2X1_LOC_213/a_36_216# OR2X1_LOC_220/A VSS VDD
+ OR2X1_LOC_213/A OR2X1_LOC_213/B OR2X1_LOC
XOR2X1_LOC_235 OR2X1_LOC_235/a_8_216# OR2X1_LOC_235/a_36_216# OR2X1_LOC_235/Y VSS VDD
+ OR2X1_LOC_86/A OR2X1_LOC_235/B OR2X1_LOC
XOR2X1_LOC_202 OR2X1_LOC_202/a_8_216# OR2X1_LOC_202/a_36_216# OR2X1_LOC_206/A VSS VDD
+ AND2X1_LOC_69/Y AND2X1_LOC_67/Y OR2X1_LOC
XOR2X1_LOC_224 OR2X1_LOC_224/a_8_216# OR2X1_LOC_224/a_36_216# OR2X1_LOC_224/Y VSS VDD
+ OR2X1_LOC_744/A OR2X1_LOC_31/Y OR2X1_LOC
XAND2X1_LOC_482 AND2X1_LOC_482/a_36_24# OR2X1_LOC_833/B AND2X1_LOC_482/a_8_24# VSS VDD
+ AND2X1_LOC_7/B AND2X1_LOC_59/Y AND2X1_LOC
XAND2X1_LOC_493 AND2X1_LOC_493/a_36_24# AND2X1_LOC_717/B AND2X1_LOC_493/a_8_24# VSS VDD
+ OR2X1_LOC_491/Y OR2X1_LOC_492/Y AND2X1_LOC
XAND2X1_LOC_471 AND2X1_LOC_471/a_36_24# AND2X1_LOC_471/Y AND2X1_LOC_471/a_8_24# VSS VDD
+ AND2X1_LOC_464/Y AND2X1_LOC_465/Y AND2X1_LOC
XAND2X1_LOC_460 AND2X1_LOC_460/a_36_24# AND2X1_LOC_463/B AND2X1_LOC_460/a_8_24# VSS VDD
+ OR2X1_LOC_380/Y OR2X1_LOC_409/Y AND2X1_LOC
XOR2X1_LOC_257 OR2X1_LOC_257/a_8_216# OR2X1_LOC_257/a_36_216# OR2X1_LOC_257/Y VSS VDD
+ OR2X1_LOC_427/A OR2X1_LOC_18/Y OR2X1_LOC
XOR2X1_LOC_246 OR2X1_LOC_246/a_8_216# OR2X1_LOC_246/a_36_216# OR2X1_LOC_246/Y VSS VDD
+ OR2X1_LOC_246/A OR2X1_LOC_9/Y OR2X1_LOC
XOR2X1_LOC_279 OR2X1_LOC_279/a_8_216# OR2X1_LOC_279/a_36_216# OR2X1_LOC_279/Y VSS VDD
+ OR2X1_LOC_427/A OR2X1_LOC_44/Y OR2X1_LOC
XOR2X1_LOC_268 OR2X1_LOC_268/a_8_216# OR2X1_LOC_268/a_36_216# OR2X1_LOC_268/Y VSS VDD
+ OR2X1_LOC_92/Y OR2X1_LOC_36/Y OR2X1_LOC
XOR2X1_LOC_780 OR2X1_LOC_780/a_8_216# OR2X1_LOC_780/a_36_216# OR2X1_LOC_783/A VSS VDD
+ OR2X1_LOC_780/A OR2X1_LOC_780/B OR2X1_LOC
XOR2X1_LOC_791 OR2X1_LOC_791/a_8_216# OR2X1_LOC_791/a_36_216# OR2X1_LOC_792/A VSS VDD
+ OR2X1_LOC_791/A OR2X1_LOC_791/B OR2X1_LOC
XAND2X1_LOC_290 AND2X1_LOC_290/a_36_24# OR2X1_LOC_334/B AND2X1_LOC_290/a_8_24# VSS VDD
+ OR2X1_LOC_78/B OR2X1_LOC_66/A AND2X1_LOC
XAND2X1_LOC_29 AND2X1_LOC_29/a_36_24# OR2X1_LOC_87/B AND2X1_LOC_29/a_8_24# VSS VDD
+ AND2X1_LOC_8/Y OR2X1_LOC_49/A AND2X1_LOC
XAND2X1_LOC_18 AND2X1_LOC_18/a_36_24# AND2X1_LOC_18/Y AND2X1_LOC_18/a_8_24# VSS VDD
+ AND2X1_LOC_11/Y AND2X1_LOC_17/Y AND2X1_LOC
XOR2X1_LOC_4 OR2X1_LOC_4/a_8_216# OR2X1_LOC_4/a_36_216# OR2X1_LOC_6/B VSS VDD INPUT_1
+ D_INPUT_0 OR2X1_LOC
XAND2X1_LOC_845 AND2X1_LOC_845/a_36_24# AND2X1_LOC_845/Y AND2X1_LOC_845/a_8_24# VSS VDD
+ AND2X1_LOC_721/A OR2X1_LOC_813/Y AND2X1_LOC
XAND2X1_LOC_823 AND2X1_LOC_823/a_36_24# OR2X1_LOC_836/B AND2X1_LOC_823/a_8_24# VSS VDD
+ AND2X1_LOC_51/Y OR2X1_LOC_269/B AND2X1_LOC
XAND2X1_LOC_856 AND2X1_LOC_856/a_36_24# AND2X1_LOC_863/A AND2X1_LOC_856/a_8_24# VSS VDD
+ AND2X1_LOC_856/A AND2X1_LOC_856/B AND2X1_LOC
XAND2X1_LOC_812 AND2X1_LOC_812/a_36_24# GATE_811 AND2X1_LOC_812/a_8_24# VSS VDD
+ AND2X1_LOC_810/Y AND2X1_LOC_811/Y AND2X1_LOC
XAND2X1_LOC_801 AND2X1_LOC_801/a_36_24# AND2X1_LOC_809/A AND2X1_LOC_801/a_8_24# VSS VDD
+ OR2X1_LOC_761/Y AND2X1_LOC_801/B AND2X1_LOC
XAND2X1_LOC_834 AND2X1_LOC_834/a_36_24# AND2X1_LOC_840/B AND2X1_LOC_834/a_8_24# VSS VDD
+ OR2X1_LOC_511/Y OR2X1_LOC_677/Y AND2X1_LOC
XOR2X1_LOC_609 OR2X1_LOC_609/a_8_216# OR2X1_LOC_609/a_36_216# OR2X1_LOC_609/Y VSS VDD
+ OR2X1_LOC_609/A OR2X1_LOC_59/Y OR2X1_LOC
XAND2X1_LOC_119 AND2X1_LOC_119/a_36_24# OR2X1_LOC_121/B AND2X1_LOC_119/a_8_24# VSS VDD
+ INPUT_1 OR2X1_LOC_377/A AND2X1_LOC
XAND2X1_LOC_108 AND2X1_LOC_108/a_36_24# OR2X1_LOC_114/B AND2X1_LOC_108/a_8_24# VSS VDD
+ AND2X1_LOC_59/Y OR2X1_LOC_532/B AND2X1_LOC
XOR2X1_LOC_51 OR2X1_LOC_51/a_8_216# OR2X1_LOC_51/a_36_216# OR2X1_LOC_51/Y VSS VDD
+ OR2X1_LOC_70/A OR2X1_LOC_51/B OR2X1_LOC
XOR2X1_LOC_40 OR2X1_LOC_40/a_8_216# OR2X1_LOC_40/a_36_216# OR2X1_LOC_40/Y VSS VDD
+ OR2X1_LOC_25/Y OR2X1_LOC_2/Y OR2X1_LOC
XOR2X1_LOC_95 OR2X1_LOC_95/a_8_216# OR2X1_LOC_95/a_36_216# OR2X1_LOC_95/Y VSS VDD
+ OR2X1_LOC_70/A OR2X1_LOC_11/Y OR2X1_LOC
XOR2X1_LOC_73 OR2X1_LOC_73/a_8_216# OR2X1_LOC_73/a_36_216# OR2X1_LOC_74/A VSS VDD
+ OR2X1_LOC_85/A OR2X1_LOC_9/Y OR2X1_LOC
XOR2X1_LOC_62 OR2X1_LOC_62/a_8_216# OR2X1_LOC_62/a_36_216# OR2X1_LOC_71/A VSS VDD
+ OR2X1_LOC_62/A OR2X1_LOC_62/B OR2X1_LOC
XOR2X1_LOC_84 OR2X1_LOC_84/a_8_216# OR2X1_LOC_84/a_36_216# OR2X1_LOC_84/Y VSS VDD
+ OR2X1_LOC_84/A OR2X1_LOC_84/B OR2X1_LOC
XOR2X1_LOC_406 OR2X1_LOC_406/a_8_216# OR2X1_LOC_406/a_36_216# OR2X1_LOC_406/Y VSS VDD
+ OR2X1_LOC_406/A OR2X1_LOC_95/Y OR2X1_LOC
XOR2X1_LOC_417 OR2X1_LOC_417/a_8_216# OR2X1_LOC_417/a_36_216# OR2X1_LOC_417/Y VSS VDD
+ OR2X1_LOC_417/A OR2X1_LOC_47/Y OR2X1_LOC
XOR2X1_LOC_428 OR2X1_LOC_428/a_8_216# OR2X1_LOC_428/a_36_216# OR2X1_LOC_428/Y VSS VDD
+ OR2X1_LOC_428/A OR2X1_LOC_31/Y OR2X1_LOC
XAND2X1_LOC_631 AND2X1_LOC_631/a_36_24# AND2X1_LOC_631/Y AND2X1_LOC_631/a_8_24# VSS VDD
+ AND2X1_LOC_483/Y OR2X1_LOC_625/Y AND2X1_LOC
XAND2X1_LOC_620 AND2X1_LOC_620/a_36_24# AND2X1_LOC_620/Y AND2X1_LOC_620/a_8_24# VSS VDD
+ OR2X1_LOC_528/Y OR2X1_LOC_613/Y AND2X1_LOC
XAND2X1_LOC_664 AND2X1_LOC_664/a_36_24# OR2X1_LOC_755/A AND2X1_LOC_664/a_8_24# VSS VDD
+ OR2X1_LOC_74/A OR2X1_LOC_89/A AND2X1_LOC
XAND2X1_LOC_675 AND2X1_LOC_675/a_36_24# AND2X1_LOC_675/Y AND2X1_LOC_675/a_8_24# VSS VDD
+ AND2X1_LOC_675/A OR2X1_LOC_674/Y AND2X1_LOC
XAND2X1_LOC_642 AND2X1_LOC_642/a_36_24# AND2X1_LOC_642/Y AND2X1_LOC_642/a_8_24# VSS VDD
+ OR2X1_LOC_416/Y AND2X1_LOC_520/Y AND2X1_LOC
XAND2X1_LOC_653 AND2X1_LOC_653/a_36_24# AND2X1_LOC_661/A AND2X1_LOC_653/a_8_24# VSS VDD
+ OR2X1_LOC_594/Y AND2X1_LOC_653/B AND2X1_LOC
XAND2X1_LOC_697 AND2X1_LOC_697/a_36_24# OR2X1_LOC_779/A AND2X1_LOC_697/a_8_24# VSS VDD
+ OR2X1_LOC_375/A OR2X1_LOC_269/B AND2X1_LOC
XAND2X1_LOC_686 AND2X1_LOC_686/a_36_24# AND2X1_LOC_687/B AND2X1_LOC_686/a_8_24# VSS VDD
+ OR2X1_LOC_683/Y OR2X1_LOC_684/Y AND2X1_LOC
XOR2X1_LOC_439 OR2X1_LOC_439/a_8_216# OR2X1_LOC_439/a_36_216# OR2X1_LOC_440/A VSS VDD
+ OR2X1_LOC_544/A OR2X1_LOC_439/B OR2X1_LOC
XAND2X1_LOC_6 AND2X1_LOC_6/a_36_24# AND2X1_LOC_7/B AND2X1_LOC_6/a_8_24# VSS VDD OR2X1_LOC_19/B
+ OR2X1_LOC_68/B AND2X1_LOC
XAND2X1_LOC_450 AND2X1_LOC_450/a_36_24# AND2X1_LOC_450/Y AND2X1_LOC_450/a_8_24# VSS VDD
+ OR2X1_LOC_426/Y OR2X1_LOC_427/Y AND2X1_LOC
XOR2X1_LOC_236 OR2X1_LOC_236/a_8_216# OR2X1_LOC_236/a_36_216# OR2X1_LOC_428/A VSS VDD
+ OR2X1_LOC_49/A OR2X1_LOC_6/A OR2X1_LOC
XOR2X1_LOC_258 OR2X1_LOC_258/a_8_216# OR2X1_LOC_258/a_36_216# OR2X1_LOC_258/Y VSS VDD
+ OR2X1_LOC_158/A OR2X1_LOC_89/A OR2X1_LOC
XOR2X1_LOC_225 OR2X1_LOC_225/a_8_216# OR2X1_LOC_225/a_36_216# OR2X1_LOC_417/A VSS VDD
+ OR2X1_LOC_6/A INPUT_1 OR2X1_LOC
XOR2X1_LOC_247 OR2X1_LOC_247/a_8_216# OR2X1_LOC_247/a_36_216# OR2X1_LOC_247/Y VSS VDD
+ AND2X1_LOC_41/A AND2X1_LOC_7/B OR2X1_LOC
XOR2X1_LOC_203 OR2X1_LOC_203/a_8_216# OR2X1_LOC_203/a_36_216# OR2X1_LOC_203/Y VSS VDD
+ OR2X1_LOC_76/Y AND2X1_LOC_72/Y OR2X1_LOC
XOR2X1_LOC_214 OR2X1_LOC_214/a_8_216# OR2X1_LOC_214/a_36_216# OR2X1_LOC_219/B VSS VDD
+ OR2X1_LOC_214/A OR2X1_LOC_214/B OR2X1_LOC
XAND2X1_LOC_483 AND2X1_LOC_483/a_36_24# AND2X1_LOC_483/Y AND2X1_LOC_483/a_8_24# VSS VDD
+ OR2X1_LOC_252/Y OR2X1_LOC_482/Y AND2X1_LOC
XAND2X1_LOC_494 AND2X1_LOC_494/a_36_24# OR2X1_LOC_558/A AND2X1_LOC_494/a_8_24# VSS VDD
+ AND2X1_LOC_12/Y OR2X1_LOC_383/Y AND2X1_LOC
XAND2X1_LOC_472 AND2X1_LOC_472/a_36_24# AND2X1_LOC_476/A AND2X1_LOC_472/a_8_24# VSS VDD
+ AND2X1_LOC_462/Y AND2X1_LOC_472/B AND2X1_LOC
XAND2X1_LOC_461 AND2X1_LOC_461/a_36_24# AND2X1_LOC_462/B AND2X1_LOC_461/a_8_24# VSS VDD
+ OR2X1_LOC_411/Y OR2X1_LOC_413/Y AND2X1_LOC
XOR2X1_LOC_269 OR2X1_LOC_269/a_8_216# OR2X1_LOC_269/a_36_216# OR2X1_LOC_269/Y VSS VDD
+ OR2X1_LOC_269/A OR2X1_LOC_269/B OR2X1_LOC
XOR2X1_LOC_781 OR2X1_LOC_781/a_8_216# OR2X1_LOC_781/a_36_216# OR2X1_LOC_781/Y VSS VDD
+ OR2X1_LOC_781/A OR2X1_LOC_781/B OR2X1_LOC
XOR2X1_LOC_792 OR2X1_LOC_792/a_8_216# OR2X1_LOC_792/a_36_216# OR2X1_LOC_792/Y VSS VDD
+ OR2X1_LOC_792/A OR2X1_LOC_792/B OR2X1_LOC
XOR2X1_LOC_770 OR2X1_LOC_770/a_8_216# OR2X1_LOC_770/a_36_216# OR2X1_LOC_770/Y VSS VDD
+ OR2X1_LOC_770/A OR2X1_LOC_770/B OR2X1_LOC
XAND2X1_LOC_280 AND2X1_LOC_280/a_36_24# OR2X1_LOC_542/B AND2X1_LOC_280/a_8_24# VSS VDD
+ AND2X1_LOC_47/Y OR2X1_LOC_269/B AND2X1_LOC
XAND2X1_LOC_291 AND2X1_LOC_291/a_36_24# OR2X1_LOC_334/A AND2X1_LOC_291/a_8_24# VSS VDD
+ AND2X1_LOC_36/Y AND2X1_LOC_824/B AND2X1_LOC
XAND2X1_LOC_19 AND2X1_LOC_19/a_36_24# AND2X1_LOC_19/Y AND2X1_LOC_19/a_8_24# VSS VDD
+ OR2X1_LOC_6/B OR2X1_LOC_68/B AND2X1_LOC
XOR2X1_LOC_5 OR2X1_LOC_5/a_8_216# OR2X1_LOC_5/a_36_216# OR2X1_LOC_6/A VSS VDD D_INPUT_3
+ INPUT_2 OR2X1_LOC
XAND2X1_LOC_835 AND2X1_LOC_835/a_36_24# AND2X1_LOC_839/A AND2X1_LOC_835/a_8_24# VSS VDD
+ OR2X1_LOC_821/Y OR2X1_LOC_822/Y AND2X1_LOC
XAND2X1_LOC_813 AND2X1_LOC_813/a_36_24# OR2X1_LOC_845/A AND2X1_LOC_813/a_8_24# VSS VDD
+ OR2X1_LOC_71/A OR2X1_LOC_266/A AND2X1_LOC
XAND2X1_LOC_846 AND2X1_LOC_846/a_36_24# AND2X1_LOC_848/A AND2X1_LOC_846/a_8_24# VSS VDD
+ OR2X1_LOC_815/Y OR2X1_LOC_816/Y AND2X1_LOC
XAND2X1_LOC_824 AND2X1_LOC_824/a_36_24# OR2X1_LOC_836/A AND2X1_LOC_824/a_8_24# VSS VDD
+ OR2X1_LOC_66/A AND2X1_LOC_824/B AND2X1_LOC
XAND2X1_LOC_857 AND2X1_LOC_857/a_36_24# AND2X1_LOC_857/Y AND2X1_LOC_857/a_8_24# VSS VDD
+ AND2X1_LOC_852/Y AND2X1_LOC_853/Y AND2X1_LOC
XAND2X1_LOC_802 AND2X1_LOC_802/a_36_24# AND2X1_LOC_802/Y AND2X1_LOC_802/a_8_24# VSS VDD
+ AND2X1_LOC_798/Y AND2X1_LOC_802/B AND2X1_LOC
XAND2X1_LOC_109 AND2X1_LOC_109/a_36_24# OR2X1_LOC_112/B AND2X1_LOC_109/a_8_24# VSS VDD
+ AND2X1_LOC_31/Y OR2X1_LOC_78/A AND2X1_LOC
XOR2X1_LOC_30 OR2X1_LOC_30/a_8_216# OR2X1_LOC_30/a_36_216# OR2X1_LOC_51/B VSS VDD
+ D_INPUT_5 D_INPUT_4 OR2X1_LOC
XOR2X1_LOC_418 OR2X1_LOC_418/a_8_216# OR2X1_LOC_418/a_36_216# OR2X1_LOC_418/Y VSS VDD
+ OR2X1_LOC_51/Y OR2X1_LOC_16/A OR2X1_LOC
XOR2X1_LOC_429 OR2X1_LOC_429/a_8_216# OR2X1_LOC_429/a_36_216# OR2X1_LOC_429/Y VSS VDD
+ OR2X1_LOC_11/Y INPUT_7 OR2X1_LOC
XOR2X1_LOC_41 OR2X1_LOC_41/a_8_216# OR2X1_LOC_41/a_36_216# OR2X1_LOC_41/Y VSS VDD
+ OR2X1_LOC_40/Y OR2X1_LOC_13/B OR2X1_LOC
XOR2X1_LOC_407 OR2X1_LOC_407/a_8_216# OR2X1_LOC_407/a_36_216# OR2X1_LOC_828/B VSS VDD
+ OR2X1_LOC_155/A AND2X1_LOC_56/B OR2X1_LOC
XAND2X1_LOC_610 AND2X1_LOC_610/a_36_24# OR2X1_LOC_612/B AND2X1_LOC_610/a_8_24# VSS VDD
+ OR2X1_LOC_40/Y OR2X1_LOC_47/Y AND2X1_LOC
XAND2X1_LOC_632 AND2X1_LOC_632/a_36_24# AND2X1_LOC_658/B AND2X1_LOC_632/a_8_24# VSS VDD
+ AND2X1_LOC_632/A AND2X1_LOC_631/Y AND2X1_LOC
XAND2X1_LOC_621 AND2X1_LOC_621/a_36_24# AND2X1_LOC_621/Y AND2X1_LOC_621/a_8_24# VSS VDD
+ OR2X1_LOC_616/Y OR2X1_LOC_617/Y AND2X1_LOC
XOR2X1_LOC_96 OR2X1_LOC_96/a_8_216# OR2X1_LOC_96/a_36_216# OR2X1_LOC_96/Y VSS VDD
+ OR2X1_LOC_95/Y OR2X1_LOC_96/B OR2X1_LOC
XOR2X1_LOC_85 OR2X1_LOC_85/a_8_216# OR2X1_LOC_85/a_36_216# OR2X1_LOC_86/A VSS VDD
+ OR2X1_LOC_85/A OR2X1_LOC_18/Y OR2X1_LOC
XOR2X1_LOC_63 OR2X1_LOC_63/a_8_216# OR2X1_LOC_63/a_36_216# OR2X1_LOC_65/B VSS VDD
+ OR2X1_LOC_71/A OR2X1_LOC_8/Y OR2X1_LOC
XOR2X1_LOC_74 OR2X1_LOC_74/a_8_216# OR2X1_LOC_74/a_36_216# OR2X1_LOC_74/Y VSS VDD
+ OR2X1_LOC_74/A OR2X1_LOC_31/Y OR2X1_LOC
XOR2X1_LOC_52 OR2X1_LOC_52/a_8_216# OR2X1_LOC_52/a_36_216# OR2X1_LOC_52/Y VSS VDD
+ OR2X1_LOC_51/Y OR2X1_LOC_52/B OR2X1_LOC
XAND2X1_LOC_665 AND2X1_LOC_665/a_36_24# OR2X1_LOC_719/B AND2X1_LOC_665/a_8_24# VSS VDD
+ AND2X1_LOC_3/Y OR2X1_LOC_664/Y AND2X1_LOC
XAND2X1_LOC_643 AND2X1_LOC_643/a_36_24# AND2X1_LOC_649/B AND2X1_LOC_643/a_8_24# VSS VDD
+ AND2X1_LOC_537/Y OR2X1_LOC_595/Y AND2X1_LOC
XAND2X1_LOC_654 AND2X1_LOC_654/a_36_24# AND2X1_LOC_654/Y AND2X1_LOC_654/a_8_24# VSS VDD
+ AND2X1_LOC_650/Y AND2X1_LOC_654/B AND2X1_LOC
XAND2X1_LOC_698 AND2X1_LOC_698/a_36_24# OR2X1_LOC_709/B AND2X1_LOC_698/a_8_24# VSS VDD
+ AND2X1_LOC_64/Y OR2X1_LOC_160/A AND2X1_LOC
XAND2X1_LOC_687 AND2X1_LOC_687/a_36_24# AND2X1_LOC_687/Y AND2X1_LOC_687/a_8_24# VSS VDD
+ AND2X1_LOC_687/A AND2X1_LOC_687/B AND2X1_LOC
XAND2X1_LOC_676 AND2X1_LOC_676/a_36_24# OR2X1_LOC_679/B AND2X1_LOC_676/a_8_24# VSS VDD
+ OR2X1_LOC_427/A OR2X1_LOC_599/A AND2X1_LOC
XAND2X1_LOC_7 AND2X1_LOC_7/a_36_24# AND2X1_LOC_7/Y AND2X1_LOC_7/a_8_24# VSS VDD AND2X1_LOC_3/Y
+ AND2X1_LOC_7/B AND2X1_LOC
XAND2X1_LOC_473 AND2X1_LOC_473/a_36_24# AND2X1_LOC_473/Y AND2X1_LOC_473/a_8_24# VSS VDD
+ AND2X1_LOC_116/Y AND2X1_LOC_276/Y AND2X1_LOC
XAND2X1_LOC_462 AND2X1_LOC_462/a_36_24# AND2X1_LOC_462/Y AND2X1_LOC_462/a_8_24# VSS VDD
+ OR2X1_LOC_416/Y AND2X1_LOC_462/B AND2X1_LOC
XAND2X1_LOC_440 AND2X1_LOC_440/a_36_24# AND2X1_LOC_468/B AND2X1_LOC_440/a_8_24# VSS VDD
+ OR2X1_LOC_437/Y AND2X1_LOC_675/A AND2X1_LOC
XAND2X1_LOC_451 AND2X1_LOC_451/a_36_24# AND2X1_LOC_451/Y AND2X1_LOC_451/a_8_24# VSS VDD
+ OR2X1_LOC_428/Y OR2X1_LOC_430/Y AND2X1_LOC
XOR2X1_LOC_259 OR2X1_LOC_259/a_8_216# OR2X1_LOC_259/a_36_216# OR2X1_LOC_555/B VSS VDD
+ OR2X1_LOC_259/A OR2X1_LOC_259/B OR2X1_LOC
XOR2X1_LOC_248 OR2X1_LOC_248/a_8_216# OR2X1_LOC_248/a_36_216# OR2X1_LOC_248/Y VSS VDD
+ OR2X1_LOC_248/A OR2X1_LOC_47/Y OR2X1_LOC
XOR2X1_LOC_204 OR2X1_LOC_204/a_8_216# OR2X1_LOC_204/a_36_216# OR2X1_LOC_204/Y VSS VDD
+ OR2X1_LOC_84/Y AND2X1_LOC_79/Y OR2X1_LOC
XOR2X1_LOC_226 OR2X1_LOC_226/a_8_216# OR2X1_LOC_226/a_36_216# OR2X1_LOC_226/Y VSS VDD
+ OR2X1_LOC_417/A OR2X1_LOC_18/Y OR2X1_LOC
XOR2X1_LOC_215 OR2X1_LOC_215/a_8_216# OR2X1_LOC_215/a_36_216# OR2X1_LOC_215/Y VSS VDD
+ OR2X1_LOC_215/A OR2X1_LOC_205/Y OR2X1_LOC
XOR2X1_LOC_237 OR2X1_LOC_237/a_8_216# OR2X1_LOC_237/a_36_216# OR2X1_LOC_237/Y VSS VDD
+ OR2X1_LOC_428/A OR2X1_LOC_26/Y OR2X1_LOC
XAND2X1_LOC_495 AND2X1_LOC_495/a_36_24# OR2X1_LOC_499/B AND2X1_LOC_495/a_8_24# VSS VDD
+ AND2X1_LOC_36/Y AND2X1_LOC_56/B AND2X1_LOC
XAND2X1_LOC_484 AND2X1_LOC_484/a_36_24# OR2X1_LOC_486/B AND2X1_LOC_484/a_8_24# VSS VDD
+ AND2X1_LOC_41/A AND2X1_LOC_36/Y AND2X1_LOC
XOR2X1_LOC_782 OR2X1_LOC_782/a_8_216# OR2X1_LOC_782/a_36_216# OR2X1_LOC_797/A VSS VDD
+ OR2X1_LOC_781/Y OR2X1_LOC_782/B OR2X1_LOC
XOR2X1_LOC_760 OR2X1_LOC_760/a_8_216# OR2X1_LOC_760/a_36_216# OR2X1_LOC_760/Y VSS VDD
+ OR2X1_LOC_329/B OR2X1_LOC_64/Y OR2X1_LOC
XOR2X1_LOC_771 OR2X1_LOC_771/a_8_216# OR2X1_LOC_771/a_36_216# OR2X1_LOC_774/B VSS VDD
+ OR2X1_LOC_770/Y OR2X1_LOC_771/B OR2X1_LOC
XOR2X1_LOC_793 OR2X1_LOC_793/a_8_216# OR2X1_LOC_793/a_36_216# OR2X1_LOC_805/A VSS VDD
+ OR2X1_LOC_793/A OR2X1_LOC_793/B OR2X1_LOC
XAND2X1_LOC_292 AND2X1_LOC_292/a_36_24# OR2X1_LOC_346/B AND2X1_LOC_292/a_8_24# VSS VDD
+ AND2X1_LOC_40/Y OR2X1_LOC_151/A AND2X1_LOC
XAND2X1_LOC_281 AND2X1_LOC_281/a_36_24# OR2X1_LOC_285/B AND2X1_LOC_281/a_8_24# VSS VDD
+ AND2X1_LOC_3/Y OR2X1_LOC_269/B AND2X1_LOC
XAND2X1_LOC_270 AND2X1_LOC_270/a_36_24# OR2X1_LOC_368/A AND2X1_LOC_270/a_8_24# VSS VDD
+ OR2X1_LOC_18/Y OR2X1_LOC_36/Y AND2X1_LOC
XOR2X1_LOC_590 OR2X1_LOC_590/a_8_216# OR2X1_LOC_590/a_36_216# OR2X1_LOC_590/Y VSS VDD
+ OR2X1_LOC_532/B OR2X1_LOC_154/A OR2X1_LOC
XOR2X1_LOC_6 OR2X1_LOC_6/a_8_216# OR2X1_LOC_6/a_36_216# OR2X1_LOC_7/A VSS VDD OR2X1_LOC_6/A
+ OR2X1_LOC_6/B OR2X1_LOC
XAND2X1_LOC_814 AND2X1_LOC_814/a_36_24# OR2X1_LOC_815/A AND2X1_LOC_814/a_8_24# VSS VDD
+ OR2X1_LOC_600/A OR2X1_LOC_417/A AND2X1_LOC
XAND2X1_LOC_803 AND2X1_LOC_803/a_36_24# AND2X1_LOC_808/A AND2X1_LOC_803/a_8_24# VSS VDD
+ AND2X1_LOC_796/Y AND2X1_LOC_803/B AND2X1_LOC
XAND2X1_LOC_858 AND2X1_LOC_858/a_36_24# AND2X1_LOC_862/A AND2X1_LOC_858/a_8_24# VSS VDD
+ AND2X1_LOC_850/Y AND2X1_LOC_858/B AND2X1_LOC
XAND2X1_LOC_836 AND2X1_LOC_836/a_36_24# AND2X1_LOC_839/B AND2X1_LOC_836/a_8_24# VSS VDD
+ OR2X1_LOC_823/Y OR2X1_LOC_824/Y AND2X1_LOC
XAND2X1_LOC_847 AND2X1_LOC_847/a_36_24# AND2X1_LOC_847/Y AND2X1_LOC_847/a_8_24# VSS VDD
+ OR2X1_LOC_817/Y OR2X1_LOC_820/Y AND2X1_LOC
XAND2X1_LOC_825 AND2X1_LOC_825/a_36_24# OR2X1_LOC_837/B AND2X1_LOC_825/a_8_24# VSS VDD
+ AND2X1_LOC_44/Y AND2X1_LOC_94/Y AND2X1_LOC
XOR2X1_LOC_64 OR2X1_LOC_64/a_8_216# OR2X1_LOC_64/a_36_216# OR2X1_LOC_64/Y VSS VDD
+ OR2X1_LOC_70/A OR2X1_LOC_22/A OR2X1_LOC
XOR2X1_LOC_31 OR2X1_LOC_31/a_8_216# OR2X1_LOC_31/a_36_216# OR2X1_LOC_31/Y VSS VDD
+ OR2X1_LOC_51/B OR2X1_LOC_3/B OR2X1_LOC
XOR2X1_LOC_53 OR2X1_LOC_53/a_8_216# OR2X1_LOC_53/a_36_216# OR2X1_LOC_53/Y VSS VDD
+ OR2X1_LOC_70/A INPUT_5 OR2X1_LOC
XOR2X1_LOC_42 OR2X1_LOC_42/a_8_216# OR2X1_LOC_42/a_36_216# OR2X1_LOC_43/A VSS VDD
+ OR2X1_LOC_85/A D_INPUT_1 OR2X1_LOC
XOR2X1_LOC_20 OR2X1_LOC_20/a_8_216# OR2X1_LOC_20/a_36_216# OR2X1_LOC_20/Y VSS VDD
+ OR2X1_LOC_20/A OR2X1_LOC_18/Y OR2X1_LOC
XOR2X1_LOC_408 OR2X1_LOC_408/a_8_216# OR2X1_LOC_408/a_36_216# OR2X1_LOC_408/Y VSS VDD
+ OR2X1_LOC_22/A INPUT_6 OR2X1_LOC
XOR2X1_LOC_419 OR2X1_LOC_419/a_8_216# OR2X1_LOC_419/a_36_216# OR2X1_LOC_419/Y VSS VDD
+ OR2X1_LOC_43/A OR2X1_LOC_36/Y OR2X1_LOC
XAND2X1_LOC_633 AND2X1_LOC_633/a_36_24# AND2X1_LOC_633/Y AND2X1_LOC_633/a_8_24# VSS VDD
+ OR2X1_LOC_118/Y OR2X1_LOC_278/A AND2X1_LOC
XAND2X1_LOC_611 AND2X1_LOC_611/a_36_24# AND2X1_LOC_612/B AND2X1_LOC_611/a_8_24# VSS VDD
+ OR2X1_LOC_68/B OR2X1_LOC_54/Y AND2X1_LOC
XAND2X1_LOC_666 AND2X1_LOC_666/a_36_24# OR2X1_LOC_719/A AND2X1_LOC_666/a_8_24# VSS VDD
+ AND2X1_LOC_18/Y OR2X1_LOC_121/A AND2X1_LOC
XAND2X1_LOC_600 AND2X1_LOC_600/a_36_24# OR2X1_LOC_602/B AND2X1_LOC_600/a_8_24# VSS VDD
+ AND2X1_LOC_31/Y OR2X1_LOC_756/B AND2X1_LOC
XAND2X1_LOC_655 AND2X1_LOC_655/a_36_24# AND2X1_LOC_660/A AND2X1_LOC_655/a_8_24# VSS VDD
+ AND2X1_LOC_655/A AND2X1_LOC_649/Y AND2X1_LOC
XAND2X1_LOC_644 AND2X1_LOC_644/a_36_24# AND2X1_LOC_644/Y AND2X1_LOC_644/a_8_24# VSS VDD
+ OR2X1_LOC_597/Y OR2X1_LOC_599/Y AND2X1_LOC
XAND2X1_LOC_622 AND2X1_LOC_622/a_36_24# AND2X1_LOC_624/A AND2X1_LOC_622/a_8_24# VSS VDD
+ OR2X1_LOC_619/Y AND2X1_LOC_621/Y AND2X1_LOC
XOR2X1_LOC_86 OR2X1_LOC_86/a_8_216# OR2X1_LOC_86/a_36_216# OR2X1_LOC_86/Y VSS VDD
+ OR2X1_LOC_86/A D_INPUT_0 OR2X1_LOC
XOR2X1_LOC_97 OR2X1_LOC_97/a_8_216# OR2X1_LOC_97/a_36_216# OR2X1_LOC_99/B VSS VDD
+ OR2X1_LOC_97/A OR2X1_LOC_97/B OR2X1_LOC
XOR2X1_LOC_75 OR2X1_LOC_75/a_8_216# OR2X1_LOC_75/a_36_216# OR2X1_LOC_75/Y VSS VDD
+ OR2X1_LOC_59/Y OR2X1_LOC_45/B OR2X1_LOC
XAND2X1_LOC_699 AND2X1_LOC_699/a_36_24# OR2X1_LOC_709/A AND2X1_LOC_699/a_8_24# VSS VDD
+ OR2X1_LOC_377/A OR2X1_LOC_375/A AND2X1_LOC
XAND2X1_LOC_688 AND2X1_LOC_688/a_36_24# OR2X1_LOC_689/A AND2X1_LOC_688/a_8_24# VSS VDD
+ OR2X1_LOC_39/A OR2X1_LOC_585/A AND2X1_LOC
XAND2X1_LOC_677 AND2X1_LOC_677/a_36_24# OR2X1_LOC_834/A AND2X1_LOC_677/a_8_24# VSS VDD
+ OR2X1_LOC_66/A OR2X1_LOC_161/B AND2X1_LOC
XAND2X1_LOC_8 AND2X1_LOC_8/a_36_24# AND2X1_LOC_8/Y AND2X1_LOC_8/a_8_24# VSS VDD INPUT_2
+ D_INPUT_3 AND2X1_LOC
XAND2X1_LOC_474 AND2X1_LOC_474/a_36_24# AND2X1_LOC_474/Y AND2X1_LOC_474/a_8_24# VSS VDD
+ AND2X1_LOC_474/A AND2X1_LOC_573/A AND2X1_LOC
XAND2X1_LOC_496 AND2X1_LOC_496/a_36_24# OR2X1_LOC_778/A AND2X1_LOC_496/a_8_24# VSS VDD
+ AND2X1_LOC_18/Y AND2X1_LOC_56/B AND2X1_LOC
XAND2X1_LOC_441 AND2X1_LOC_441/a_36_24# OR2X1_LOC_545/B AND2X1_LOC_441/a_8_24# VSS VDD
+ AND2X1_LOC_40/Y OR2X1_LOC_87/A AND2X1_LOC
XAND2X1_LOC_485 AND2X1_LOC_485/a_36_24# OR2X1_LOC_705/B AND2X1_LOC_485/a_8_24# VSS VDD
+ AND2X1_LOC_44/Y OR2X1_LOC_532/B AND2X1_LOC
XAND2X1_LOC_463 AND2X1_LOC_463/a_36_24# AND2X1_LOC_472/B AND2X1_LOC_463/a_8_24# VSS VDD
+ AND2X1_LOC_459/Y AND2X1_LOC_463/B AND2X1_LOC
XAND2X1_LOC_430 AND2X1_LOC_430/a_36_24# OR2X1_LOC_451/A AND2X1_LOC_430/a_8_24# VSS VDD
+ OR2X1_LOC_161/A AND2X1_LOC_430/B AND2X1_LOC
XAND2X1_LOC_452 AND2X1_LOC_452/a_36_24# AND2X1_LOC_452/Y AND2X1_LOC_452/a_8_24# VSS VDD
+ AND2X1_LOC_450/Y AND2X1_LOC_451/Y AND2X1_LOC
XOR2X1_LOC_249 OR2X1_LOC_249/a_8_216# OR2X1_LOC_249/a_36_216# OR2X1_LOC_249/Y VSS VDD
+ OR2X1_LOC_154/A OR2X1_LOC_160/B OR2X1_LOC
XOR2X1_LOC_205 OR2X1_LOC_205/a_8_216# OR2X1_LOC_205/a_36_216# OR2X1_LOC_205/Y VSS VDD
+ OR2X1_LOC_204/Y OR2X1_LOC_203/Y OR2X1_LOC
XOR2X1_LOC_216 OR2X1_LOC_216/a_8_216# OR2X1_LOC_216/a_36_216# OR2X1_LOC_216/Y VSS VDD
+ OR2X1_LOC_216/A OR2X1_LOC_656/B OR2X1_LOC
XOR2X1_LOC_227 OR2X1_LOC_227/a_8_216# OR2X1_LOC_227/a_36_216# OR2X1_LOC_227/Y VSS VDD
+ OR2X1_LOC_227/A OR2X1_LOC_227/B OR2X1_LOC
XOR2X1_LOC_238 OR2X1_LOC_238/a_8_216# OR2X1_LOC_238/a_36_216# OR2X1_LOC_238/Y VSS VDD
+ OR2X1_LOC_51/Y OR2X1_LOC_45/B OR2X1_LOC
XOR2X1_LOC_783 OR2X1_LOC_783/a_8_216# OR2X1_LOC_783/a_36_216# OR2X1_LOC_796/B VSS VDD
+ OR2X1_LOC_783/A OR2X1_LOC_779/Y OR2X1_LOC
XOR2X1_LOC_761 OR2X1_LOC_761/a_8_216# OR2X1_LOC_761/a_36_216# OR2X1_LOC_761/Y VSS VDD
+ OR2X1_LOC_599/Y INPUT_0 OR2X1_LOC
XOR2X1_LOC_772 OR2X1_LOC_772/a_8_216# OR2X1_LOC_772/a_36_216# OR2X1_LOC_772/Y VSS VDD
+ OR2X1_LOC_772/A OR2X1_LOC_772/B OR2X1_LOC
XOR2X1_LOC_794 OR2X1_LOC_794/a_8_216# OR2X1_LOC_794/a_36_216# OR2X1_LOC_804/B VSS VDD
+ OR2X1_LOC_794/A OR2X1_LOC_787/Y OR2X1_LOC
XOR2X1_LOC_750 OR2X1_LOC_750/a_8_216# OR2X1_LOC_750/a_36_216# OR2X1_LOC_750/Y VSS VDD
+ OR2X1_LOC_750/A OR2X1_LOC_161/A OR2X1_LOC
XAND2X1_LOC_271 AND2X1_LOC_271/a_36_24# OR2X1_LOC_276/B AND2X1_LOC_271/a_8_24# VSS VDD
+ OR2X1_LOC_269/Y OR2X1_LOC_270/Y AND2X1_LOC
XAND2X1_LOC_282 AND2X1_LOC_282/a_36_24# OR2X1_LOC_285/A AND2X1_LOC_282/a_8_24# VSS VDD
+ OR2X1_LOC_532/B OR2X1_LOC_375/A AND2X1_LOC
XAND2X1_LOC_260 AND2X1_LOC_260/a_36_24# OR2X1_LOC_261/A AND2X1_LOC_260/a_8_24# VSS VDD
+ OR2X1_LOC_12/Y OR2X1_LOC_158/A AND2X1_LOC
XAND2X1_LOC_293 AND2X1_LOC_293/a_36_24# OR2X1_LOC_598/A AND2X1_LOC_293/a_8_24# VSS VDD
+ INPUT_1 OR2X1_LOC_68/B AND2X1_LOC
XOR2X1_LOC_580 OR2X1_LOC_580/a_8_216# OR2X1_LOC_580/a_36_216# D_GATE_579 VSS VDD
+ OR2X1_LOC_580/A OR2X1_LOC_580/B OR2X1_LOC
XOR2X1_LOC_591 OR2X1_LOC_591/a_8_216# OR2X1_LOC_591/a_36_216# OR2X1_LOC_591/Y VSS VDD
+ OR2X1_LOC_591/A OR2X1_LOC_64/Y OR2X1_LOC
XOR2X1_LOC_7 OR2X1_LOC_7/a_8_216# OR2X1_LOC_7/a_36_216# OR2X1_LOC_7/Y VSS VDD OR2X1_LOC_7/A
+ OR2X1_LOC_3/Y OR2X1_LOC
XAND2X1_LOC_837 AND2X1_LOC_837/a_36_24# AND2X1_LOC_838/B AND2X1_LOC_837/a_8_24# VSS VDD
+ OR2X1_LOC_825/Y OR2X1_LOC_826/Y AND2X1_LOC
XAND2X1_LOC_848 AND2X1_LOC_848/a_36_24# AND2X1_LOC_848/Y AND2X1_LOC_848/a_8_24# VSS VDD
+ AND2X1_LOC_848/A AND2X1_LOC_847/Y AND2X1_LOC
XAND2X1_LOC_815 AND2X1_LOC_815/a_36_24# OR2X1_LOC_846/B AND2X1_LOC_815/a_8_24# VSS VDD
+ AND2X1_LOC_3/Y OR2X1_LOC_814/Y AND2X1_LOC
XAND2X1_LOC_826 AND2X1_LOC_826/a_36_24# OR2X1_LOC_837/A AND2X1_LOC_826/a_8_24# VSS VDD
+ AND2X1_LOC_56/B AND2X1_LOC_95/Y AND2X1_LOC
XAND2X1_LOC_804 AND2X1_LOC_804/a_36_24# AND2X1_LOC_804/Y AND2X1_LOC_804/a_8_24# VSS VDD
+ AND2X1_LOC_804/A AND2X1_LOC_795/Y AND2X1_LOC
XAND2X1_LOC_859 AND2X1_LOC_859/a_36_24# AND2X1_LOC_859/Y AND2X1_LOC_859/a_8_24# VSS VDD
+ AND2X1_LOC_848/Y AND2X1_LOC_859/B AND2X1_LOC
XOR2X1_LOC_21 OR2X1_LOC_21/a_8_216# OR2X1_LOC_21/a_36_216# OR2X1_LOC_22/A VSS VDD
+ INPUT_5 D_INPUT_4 OR2X1_LOC
XOR2X1_LOC_43 OR2X1_LOC_43/a_8_216# OR2X1_LOC_43/a_36_216# OR2X1_LOC_43/Y VSS VDD
+ OR2X1_LOC_43/A OR2X1_LOC_22/Y OR2X1_LOC
XOR2X1_LOC_54 OR2X1_LOC_54/a_8_216# OR2X1_LOC_54/a_36_216# OR2X1_LOC_54/Y VSS VDD
+ D_INPUT_1 D_INPUT_0 OR2X1_LOC
XOR2X1_LOC_10 OR2X1_LOC_10/a_8_216# OR2X1_LOC_10/a_36_216# OR2X1_LOC_13/B VSS VDD
+ OR2X1_LOC_9/Y OR2X1_LOC_8/Y OR2X1_LOC
XOR2X1_LOC_76 OR2X1_LOC_76/a_8_216# OR2X1_LOC_76/a_36_216# OR2X1_LOC_76/Y VSS VDD
+ OR2X1_LOC_76/A OR2X1_LOC_76/B OR2X1_LOC
XOR2X1_LOC_87 OR2X1_LOC_87/a_8_216# OR2X1_LOC_87/a_36_216# OR2X1_LOC_87/Y VSS VDD
+ OR2X1_LOC_87/A OR2X1_LOC_87/B OR2X1_LOC
XOR2X1_LOC_32 OR2X1_LOC_32/a_8_216# OR2X1_LOC_32/a_36_216# OR2X1_LOC_32/Y VSS VDD
+ OR2X1_LOC_31/Y OR2X1_LOC_32/B OR2X1_LOC
XOR2X1_LOC_65 OR2X1_LOC_65/a_8_216# OR2X1_LOC_65/a_36_216# OR2X1_LOC_65/Y VSS VDD
+ OR2X1_LOC_64/Y OR2X1_LOC_65/B OR2X1_LOC
XOR2X1_LOC_409 OR2X1_LOC_409/a_8_216# OR2X1_LOC_409/a_36_216# OR2X1_LOC_409/Y VSS VDD
+ OR2X1_LOC_408/Y OR2X1_LOC_409/B OR2X1_LOC
XAND2X1_LOC_656 AND2X1_LOC_656/a_36_24# AND2X1_LOC_656/Y AND2X1_LOC_656/a_8_24# VSS VDD
+ AND2X1_LOC_216/A AND2X1_LOC_647/Y AND2X1_LOC
XAND2X1_LOC_612 AND2X1_LOC_612/a_36_24# OR2X1_LOC_647/B AND2X1_LOC_612/a_8_24# VSS VDD
+ OR2X1_LOC_610/Y AND2X1_LOC_612/B AND2X1_LOC
XAND2X1_LOC_667 AND2X1_LOC_667/a_36_24# OR2X1_LOC_720/B AND2X1_LOC_667/a_8_24# VSS VDD
+ AND2X1_LOC_64/Y OR2X1_LOC_264/Y AND2X1_LOC
XAND2X1_LOC_623 AND2X1_LOC_623/a_36_24# AND2X1_LOC_624/B AND2X1_LOC_623/a_8_24# VSS VDD
+ OR2X1_LOC_615/Y AND2X1_LOC_620/Y AND2X1_LOC
XAND2X1_LOC_601 AND2X1_LOC_601/a_36_24# OR2X1_LOC_602/A AND2X1_LOC_601/a_8_24# VSS VDD
+ OR2X1_LOC_78/B AND2X1_LOC_47/Y AND2X1_LOC
XAND2X1_LOC_634 AND2X1_LOC_634/a_36_24# AND2X1_LOC_634/Y AND2X1_LOC_634/a_8_24# VSS VDD
+ OR2X1_LOC_290/Y OR2X1_LOC_690/A AND2X1_LOC
XAND2X1_LOC_689 AND2X1_LOC_689/a_36_24# OR2X1_LOC_691/B AND2X1_LOC_689/a_8_24# VSS VDD
+ AND2X1_LOC_31/Y OR2X1_LOC_688/Y AND2X1_LOC
XAND2X1_LOC_678 AND2X1_LOC_678/a_36_24# OR2X1_LOC_679/A AND2X1_LOC_678/a_8_24# VSS VDD
+ OR2X1_LOC_12/Y OR2X1_LOC_677/Y AND2X1_LOC
XAND2X1_LOC_645 AND2X1_LOC_645/a_36_24# AND2X1_LOC_648/B AND2X1_LOC_645/a_8_24# VSS VDD
+ AND2X1_LOC_645/A AND2X1_LOC_605/Y AND2X1_LOC
XOR2X1_LOC_98 OR2X1_LOC_98/a_8_216# OR2X1_LOC_98/a_36_216# OR2X1_LOC_99/A VSS VDD
+ OR2X1_LOC_98/A OR2X1_LOC_98/B OR2X1_LOC
XAND2X1_LOC_9 AND2X1_LOC_9/a_36_24# OR2X1_LOC_62/B AND2X1_LOC_9/a_8_24# VSS VDD D_INPUT_0
+ D_INPUT_1 AND2X1_LOC
XOR2X1_LOC_217 OR2X1_LOC_217/a_8_216# OR2X1_LOC_217/a_36_216# OR2X1_LOC_217/Y VSS VDD
+ OR2X1_LOC_217/A OR2X1_LOC_124/Y OR2X1_LOC
XOR2X1_LOC_206 OR2X1_LOC_206/a_8_216# OR2X1_LOC_206/a_36_216# OR2X1_LOC_215/A VSS VDD
+ OR2X1_LOC_206/A OR2X1_LOC_201/Y OR2X1_LOC
XOR2X1_LOC_228 OR2X1_LOC_228/a_8_216# OR2X1_LOC_228/a_36_216# OR2X1_LOC_228/Y VSS VDD
+ AND2X1_LOC_52/Y AND2X1_LOC_7/Y OR2X1_LOC
XAND2X1_LOC_497 AND2X1_LOC_497/a_36_24# OR2X1_LOC_844/B AND2X1_LOC_497/a_8_24# VSS VDD
+ AND2X1_LOC_22/Y AND2X1_LOC_72/B AND2X1_LOC
XAND2X1_LOC_464 AND2X1_LOC_464/a_36_24# AND2X1_LOC_464/Y AND2X1_LOC_464/a_8_24# VSS VDD
+ AND2X1_LOC_464/A AND2X1_LOC_458/Y AND2X1_LOC
XAND2X1_LOC_475 AND2X1_LOC_475/a_36_24# AND2X1_LOC_475/Y AND2X1_LOC_475/a_8_24# VSS VDD
+ OR2X1_LOC_406/Y AND2X1_LOC_474/Y AND2X1_LOC
XAND2X1_LOC_442 AND2X1_LOC_442/a_36_24# OR2X1_LOC_444/B AND2X1_LOC_442/a_8_24# VSS VDD
+ AND2X1_LOC_40/Y OR2X1_LOC_756/B AND2X1_LOC
XAND2X1_LOC_431 AND2X1_LOC_431/a_36_24# OR2X1_LOC_434/A AND2X1_LOC_431/a_8_24# VSS VDD
+ AND2X1_LOC_70/Y OR2X1_LOC_269/B AND2X1_LOC
XAND2X1_LOC_420 AND2X1_LOC_420/a_36_24# OR2X1_LOC_447/A AND2X1_LOC_420/a_8_24# VSS VDD
+ AND2X1_LOC_95/Y OR2X1_LOC_532/B AND2X1_LOC
XAND2X1_LOC_486 AND2X1_LOC_486/a_36_24# AND2X1_LOC_486/Y AND2X1_LOC_486/a_8_24# VSS VDD
+ OR2X1_LOC_484/Y OR2X1_LOC_485/Y AND2X1_LOC
XAND2X1_LOC_453 AND2X1_LOC_453/a_36_24# AND2X1_LOC_453/Y AND2X1_LOC_453/a_8_24# VSS VDD
+ AND2X1_LOC_448/Y AND2X1_LOC_449/Y AND2X1_LOC
XOR2X1_LOC_239 OR2X1_LOC_239/a_8_216# OR2X1_LOC_239/a_36_216# OR2X1_LOC_239/Y VSS VDD
+ OR2X1_LOC_485/A OR2X1_LOC_51/Y OR2X1_LOC
XOR2X1_LOC_762 OR2X1_LOC_762/a_8_216# OR2X1_LOC_762/a_36_216# OR2X1_LOC_762/Y VSS VDD
+ OR2X1_LOC_11/Y D_INPUT_6 OR2X1_LOC
XOR2X1_LOC_751 OR2X1_LOC_751/a_8_216# OR2X1_LOC_751/a_36_216# OR2X1_LOC_751/Y VSS VDD
+ OR2X1_LOC_751/A OR2X1_LOC_3/Y OR2X1_LOC
XOR2X1_LOC_740 OR2X1_LOC_740/a_8_216# OR2X1_LOC_740/a_36_216# OR2X1_LOC_742/B VSS VDD
+ OR2X1_LOC_739/Y OR2X1_LOC_740/B OR2X1_LOC
XOR2X1_LOC_784 OR2X1_LOC_784/a_8_216# OR2X1_LOC_784/a_36_216# OR2X1_LOC_784/Y VSS VDD
+ OR2X1_LOC_778/Y OR2X1_LOC_784/B OR2X1_LOC
XOR2X1_LOC_773 OR2X1_LOC_773/a_8_216# OR2X1_LOC_773/a_36_216# OR2X1_LOC_773/Y VSS VDD
+ OR2X1_LOC_772/Y OR2X1_LOC_773/B OR2X1_LOC
XOR2X1_LOC_795 OR2X1_LOC_795/a_8_216# OR2X1_LOC_795/a_36_216# OR2X1_LOC_804/A VSS VDD
+ OR2X1_LOC_786/Y OR2X1_LOC_795/B OR2X1_LOC
XAND2X1_LOC_272 AND2X1_LOC_272/a_36_24# OR2X1_LOC_541/A AND2X1_LOC_272/a_8_24# VSS VDD
+ AND2X1_LOC_31/Y AND2X1_LOC_43/B AND2X1_LOC
XAND2X1_LOC_294 AND2X1_LOC_294/a_36_24# OR2X1_LOC_481/A AND2X1_LOC_294/a_8_24# VSS VDD
+ OR2X1_LOC_13/B OR2X1_LOC_585/A AND2X1_LOC
XAND2X1_LOC_261 AND2X1_LOC_261/a_36_24# OR2X1_LOC_345/A AND2X1_LOC_261/a_8_24# VSS VDD
+ OR2X1_LOC_756/B OR2X1_LOC_260/Y AND2X1_LOC
XAND2X1_LOC_283 AND2X1_LOC_283/a_36_24# OR2X1_LOC_286/B AND2X1_LOC_283/a_8_24# VSS VDD
+ OR2X1_LOC_66/A OR2X1_LOC_814/A AND2X1_LOC
XAND2X1_LOC_250 AND2X1_LOC_250/a_36_24# OR2X1_LOC_343/B AND2X1_LOC_250/a_8_24# VSS VDD
+ AND2X1_LOC_64/Y OR2X1_LOC_249/Y AND2X1_LOC
XOR2X1_LOC_581 OR2X1_LOC_581/a_8_216# OR2X1_LOC_581/a_36_216# OR2X1_LOC_581/Y VSS VDD
+ OR2X1_LOC_2/Y D_INPUT_6 OR2X1_LOC
XOR2X1_LOC_570 OR2X1_LOC_570/a_8_216# OR2X1_LOC_570/a_36_216# OR2X1_LOC_570/Y VSS VDD
+ OR2X1_LOC_570/A OR2X1_LOC_562/Y OR2X1_LOC
XOR2X1_LOC_592 OR2X1_LOC_592/a_8_216# OR2X1_LOC_592/a_36_216# OR2X1_LOC_593/A VSS VDD
+ OR2X1_LOC_592/A OR2X1_LOC_449/B OR2X1_LOC
XOR2X1_LOC_8 OR2X1_LOC_8/a_8_216# OR2X1_LOC_8/a_36_216# OR2X1_LOC_8/Y VSS VDD INPUT_3
+ D_INPUT_2 OR2X1_LOC
XAND2X1_LOC_849 AND2X1_LOC_849/a_36_24# AND2X1_LOC_859/B AND2X1_LOC_849/a_8_24# VSS VDD
+ AND2X1_LOC_849/A AND2X1_LOC_845/Y AND2X1_LOC
XAND2X1_LOC_805 AND2X1_LOC_805/a_36_24# AND2X1_LOC_805/Y AND2X1_LOC_805/a_8_24# VSS VDD
+ AND2X1_LOC_792/Y AND2X1_LOC_793/Y AND2X1_LOC
XAND2X1_LOC_838 AND2X1_LOC_838/a_36_24# AND2X1_LOC_838/Y AND2X1_LOC_838/a_8_24# VSS VDD
+ OR2X1_LOC_827/Y AND2X1_LOC_838/B AND2X1_LOC
XAND2X1_LOC_816 AND2X1_LOC_816/a_36_24# OR2X1_LOC_846/A AND2X1_LOC_816/a_8_24# VSS VDD
+ AND2X1_LOC_51/Y OR2X1_LOC_185/Y AND2X1_LOC
XAND2X1_LOC_827 AND2X1_LOC_827/a_36_24# OR2X1_LOC_838/B AND2X1_LOC_827/a_8_24# VSS VDD
+ AND2X1_LOC_43/B OR2X1_LOC_375/A AND2X1_LOC
XOR2X1_LOC_11 OR2X1_LOC_11/a_8_216# OR2X1_LOC_11/a_36_216# OR2X1_LOC_11/Y VSS VDD
+ D_INPUT_5 INPUT_4 OR2X1_LOC
XOR2X1_LOC_22 OR2X1_LOC_22/a_8_216# OR2X1_LOC_22/a_36_216# OR2X1_LOC_22/Y VSS VDD
+ OR2X1_LOC_22/A OR2X1_LOC_3/B OR2X1_LOC
XOR2X1_LOC_44 OR2X1_LOC_44/a_8_216# OR2X1_LOC_44/a_36_216# OR2X1_LOC_44/Y VSS VDD
+ OR2X1_LOC_51/B OR2X1_LOC_17/Y OR2X1_LOC
XOR2X1_LOC_77 OR2X1_LOC_77/a_8_216# OR2X1_LOC_77/a_36_216# OR2X1_LOC_89/A VSS VDD
+ OR2X1_LOC_54/Y OR2X1_LOC_46/A OR2X1_LOC
XOR2X1_LOC_55 OR2X1_LOC_55/a_8_216# OR2X1_LOC_55/a_36_216# OR2X1_LOC_56/A VSS VDD
+ OR2X1_LOC_54/Y OR2X1_LOC_6/A OR2X1_LOC
XOR2X1_LOC_66 OR2X1_LOC_66/a_8_216# OR2X1_LOC_66/a_36_216# OR2X1_LOC_66/Y VSS VDD
+ OR2X1_LOC_66/A AND2X1_LOC_3/Y OR2X1_LOC
XOR2X1_LOC_88 OR2X1_LOC_88/a_8_216# OR2X1_LOC_88/a_36_216# OR2X1_LOC_88/Y VSS VDD
+ OR2X1_LOC_88/A OR2X1_LOC_3/Y OR2X1_LOC
XOR2X1_LOC_99 OR2X1_LOC_99/a_8_216# OR2X1_LOC_99/a_36_216# OR2X1_LOC_99/Y VSS VDD
+ OR2X1_LOC_99/A OR2X1_LOC_99/B OR2X1_LOC
XOR2X1_LOC_33 OR2X1_LOC_33/a_8_216# OR2X1_LOC_33/a_36_216# OR2X1_LOC_35/B VSS VDD
+ OR2X1_LOC_33/A OR2X1_LOC_33/B OR2X1_LOC
XAND2X1_LOC_657 AND2X1_LOC_657/a_36_24# AND2X1_LOC_657/Y AND2X1_LOC_657/a_8_24# VSS VDD
+ AND2X1_LOC_657/A AND2X1_LOC_574/A AND2X1_LOC
XAND2X1_LOC_646 AND2X1_LOC_646/a_36_24# AND2X1_LOC_647/B AND2X1_LOC_646/a_8_24# VSS VDD
+ OR2X1_LOC_607/Y OR2X1_LOC_609/Y AND2X1_LOC
XAND2X1_LOC_668 AND2X1_LOC_668/a_36_24# OR2X1_LOC_669/A AND2X1_LOC_668/a_8_24# VSS VDD
+ OR2X1_LOC_26/Y OR2X1_LOC_158/A AND2X1_LOC
XAND2X1_LOC_624 AND2X1_LOC_624/a_36_24# AND2X1_LOC_658/A AND2X1_LOC_624/a_8_24# VSS VDD
+ AND2X1_LOC_624/A AND2X1_LOC_624/B AND2X1_LOC
XAND2X1_LOC_613 AND2X1_LOC_613/a_36_24# OR2X1_LOC_620/A AND2X1_LOC_613/a_8_24# VSS VDD
+ AND2X1_LOC_40/Y AND2X1_LOC_56/B AND2X1_LOC
XAND2X1_LOC_679 AND2X1_LOC_679/a_36_24# OR2X1_LOC_728/B AND2X1_LOC_679/a_8_24# VSS VDD
+ OR2X1_LOC_676/Y OR2X1_LOC_678/Y AND2X1_LOC
XAND2X1_LOC_602 AND2X1_LOC_602/a_36_24# AND2X1_LOC_645/A AND2X1_LOC_602/a_8_24# VSS VDD
+ OR2X1_LOC_600/Y OR2X1_LOC_601/Y AND2X1_LOC
XAND2X1_LOC_635 AND2X1_LOC_635/a_36_24# AND2X1_LOC_639/A AND2X1_LOC_635/a_8_24# VSS VDD
+ OR2X1_LOC_428/Y OR2X1_LOC_582/Y AND2X1_LOC
XOR2X1_LOC_207 OR2X1_LOC_207/a_8_216# OR2X1_LOC_207/a_36_216# OR2X1_LOC_214/B VSS VDD
+ OR2X1_LOC_200/Y OR2X1_LOC_207/B OR2X1_LOC
XAND2X1_LOC_432 AND2X1_LOC_432/a_36_24# OR2X1_LOC_435/B AND2X1_LOC_432/a_8_24# VSS VDD
+ AND2X1_LOC_18/Y OR2X1_LOC_130/A AND2X1_LOC
XAND2X1_LOC_410 AND2X1_LOC_410/a_36_24# OR2X1_LOC_411/A AND2X1_LOC_410/a_8_24# VSS VDD
+ OR2X1_LOC_12/Y OR2X1_LOC_51/Y AND2X1_LOC
XAND2X1_LOC_421 AND2X1_LOC_421/a_36_24# OR2X1_LOC_448/B AND2X1_LOC_421/a_8_24# VSS VDD
+ AND2X1_LOC_91/B OR2X1_LOC_596/A AND2X1_LOC
XOR2X1_LOC_218 OR2X1_LOC_218/a_8_216# OR2X1_LOC_218/a_36_216# OR2X1_LOC_218/Y VSS VDD
+ OR2X1_LOC_217/Y OR2X1_LOC_216/Y OR2X1_LOC
XOR2X1_LOC_229 OR2X1_LOC_229/a_8_216# OR2X1_LOC_229/a_36_216# OR2X1_LOC_229/Y VSS VDD
+ OR2X1_LOC_45/B OR2X1_LOC_12/Y OR2X1_LOC
XAND2X1_LOC_498 AND2X1_LOC_498/a_36_24# OR2X1_LOC_501/B AND2X1_LOC_498/a_8_24# VSS VDD
+ AND2X1_LOC_70/Y OR2X1_LOC_188/Y AND2X1_LOC
XAND2X1_LOC_487 AND2X1_LOC_487/a_36_24# OR2X1_LOC_489/B AND2X1_LOC_487/a_8_24# VSS VDD
+ OR2X1_LOC_160/B AND2X1_LOC_95/Y AND2X1_LOC
XAND2X1_LOC_465 AND2X1_LOC_465/a_36_24# AND2X1_LOC_465/Y AND2X1_LOC_465/a_8_24# VSS VDD
+ AND2X1_LOC_465/A AND2X1_LOC_456/Y AND2X1_LOC
XAND2X1_LOC_476 AND2X1_LOC_476/a_36_24# AND2X1_LOC_476/Y AND2X1_LOC_476/a_8_24# VSS VDD
+ AND2X1_LOC_476/A AND2X1_LOC_473/Y AND2X1_LOC
XAND2X1_LOC_443 AND2X1_LOC_443/a_36_24# AND2X1_LOC_443/Y AND2X1_LOC_443/a_8_24# VSS VDD
+ OR2X1_LOC_91/Y OR2X1_LOC_441/Y AND2X1_LOC
XAND2X1_LOC_454 AND2X1_LOC_454/a_36_24# AND2X1_LOC_454/Y AND2X1_LOC_454/a_8_24# VSS VDD
+ AND2X1_LOC_454/A AND2X1_LOC_447/Y AND2X1_LOC
XOR2X1_LOC_763 OR2X1_LOC_763/a_8_216# OR2X1_LOC_763/a_36_216# OR2X1_LOC_763/Y VSS VDD
+ OR2X1_LOC_762/Y OR2X1_LOC_48/B OR2X1_LOC
XOR2X1_LOC_796 OR2X1_LOC_796/a_8_216# OR2X1_LOC_796/a_36_216# OR2X1_LOC_803/B VSS VDD
+ OR2X1_LOC_784/Y OR2X1_LOC_796/B OR2X1_LOC
XOR2X1_LOC_752 OR2X1_LOC_752/a_8_216# OR2X1_LOC_752/a_36_216# OR2X1_LOC_753/A VSS VDD
+ OR2X1_LOC_70/A D_INPUT_5 OR2X1_LOC
XOR2X1_LOC_774 OR2X1_LOC_774/a_8_216# OR2X1_LOC_774/a_36_216# OR2X1_LOC_774/Y VSS VDD
+ OR2X1_LOC_773/Y OR2X1_LOC_774/B OR2X1_LOC
XOR2X1_LOC_741 OR2X1_LOC_741/a_8_216# OR2X1_LOC_741/a_36_216# OR2X1_LOC_741/Y VSS VDD
+ OR2X1_LOC_741/A OR2X1_LOC_736/Y OR2X1_LOC
XOR2X1_LOC_785 OR2X1_LOC_785/a_8_216# OR2X1_LOC_785/a_36_216# OR2X1_LOC_795/B VSS VDD
+ OR2X1_LOC_776/Y OR2X1_LOC_785/B OR2X1_LOC
XOR2X1_LOC_730 OR2X1_LOC_730/a_8_216# OR2X1_LOC_730/a_36_216# OR2X1_LOC_739/A VSS VDD
+ OR2X1_LOC_730/A OR2X1_LOC_730/B OR2X1_LOC
XAND2X1_LOC_273 AND2X1_LOC_273/a_36_24# OR2X1_LOC_831/B AND2X1_LOC_273/a_8_24# VSS VDD
+ AND2X1_LOC_36/Y OR2X1_LOC_155/A AND2X1_LOC
XAND2X1_LOC_262 AND2X1_LOC_262/a_36_24# OR2X1_LOC_786/A AND2X1_LOC_262/a_8_24# VSS VDD
+ AND2X1_LOC_40/Y AND2X1_LOC_65/A AND2X1_LOC
XAND2X1_LOC_240 AND2X1_LOC_240/a_36_24# AND2X1_LOC_240/Y AND2X1_LOC_240/a_8_24# VSS VDD
+ OR2X1_LOC_232/Y OR2X1_LOC_234/Y AND2X1_LOC
XAND2X1_LOC_251 AND2X1_LOC_251/a_36_24# OR2X1_LOC_843/B AND2X1_LOC_251/a_8_24# VSS VDD
+ AND2X1_LOC_51/Y OR2X1_LOC_105/Y AND2X1_LOC
XAND2X1_LOC_284 AND2X1_LOC_284/a_36_24# AND2X1_LOC_287/B AND2X1_LOC_284/a_8_24# VSS VDD
+ OR2X1_LOC_279/Y OR2X1_LOC_280/Y AND2X1_LOC
XAND2X1_LOC_295 AND2X1_LOC_295/a_36_24# OR2X1_LOC_346/A AND2X1_LOC_295/a_8_24# VSS VDD
+ AND2X1_LOC_59/Y OR2X1_LOC_294/Y AND2X1_LOC
XOR2X1_LOC_582 OR2X1_LOC_582/a_8_216# OR2X1_LOC_582/a_36_216# OR2X1_LOC_582/Y VSS VDD
+ OR2X1_LOC_581/Y OR2X1_LOC_427/A OR2X1_LOC
XOR2X1_LOC_571 OR2X1_LOC_571/a_8_216# OR2X1_LOC_571/a_36_216# OR2X1_LOC_571/Y VSS VDD
+ OR2X1_LOC_561/Y OR2X1_LOC_571/B OR2X1_LOC
XOR2X1_LOC_560 OR2X1_LOC_560/a_8_216# OR2X1_LOC_560/a_36_216# OR2X1_LOC_571/B VSS VDD
+ OR2X1_LOC_560/A OR2X1_LOC_523/Y OR2X1_LOC
XOR2X1_LOC_593 OR2X1_LOC_593/a_8_216# OR2X1_LOC_593/a_36_216# OR2X1_LOC_799/A VSS VDD
+ OR2X1_LOC_593/A OR2X1_LOC_593/B OR2X1_LOC
XOR2X1_LOC_390 OR2X1_LOC_390/a_8_216# OR2X1_LOC_390/a_36_216# OR2X1_LOC_392/B VSS VDD
+ OR2X1_LOC_390/A OR2X1_LOC_390/B OR2X1_LOC
XOR2X1_LOC_9 OR2X1_LOC_9/a_8_216# OR2X1_LOC_9/a_36_216# OR2X1_LOC_9/Y VSS VDD INPUT_1
+ INPUT_0 OR2X1_LOC
XAND2X1_LOC_806 AND2X1_LOC_806/a_36_24# AND2X1_LOC_807/B AND2X1_LOC_806/a_8_24# VSS VDD
+ AND2X1_LOC_806/A AND2X1_LOC_675/Y AND2X1_LOC
XAND2X1_LOC_839 AND2X1_LOC_839/a_36_24# AND2X1_LOC_852/B AND2X1_LOC_839/a_8_24# VSS VDD
+ AND2X1_LOC_839/A AND2X1_LOC_839/B AND2X1_LOC
XAND2X1_LOC_817 AND2X1_LOC_817/a_36_24# OR2X1_LOC_847/B AND2X1_LOC_817/a_8_24# VSS VDD
+ D_INPUT_1 AND2X1_LOC_817/B AND2X1_LOC
XAND2X1_LOC_828 AND2X1_LOC_828/a_36_24# OR2X1_LOC_829/A AND2X1_LOC_828/a_8_24# VSS VDD
+ OR2X1_LOC_409/B OR2X1_LOC_599/A AND2X1_LOC
XOR2X1_LOC_12 OR2X1_LOC_12/a_8_216# OR2X1_LOC_12/a_36_216# OR2X1_LOC_12/Y VSS VDD
+ OR2X1_LOC_11/Y OR2X1_LOC_3/B OR2X1_LOC
XOR2X1_LOC_45 OR2X1_LOC_45/a_8_216# OR2X1_LOC_45/a_36_216# OR2X1_LOC_45/Y VSS VDD
+ OR2X1_LOC_44/Y OR2X1_LOC_45/B OR2X1_LOC
XOR2X1_LOC_56 OR2X1_LOC_56/a_8_216# OR2X1_LOC_56/a_36_216# OR2X1_LOC_56/Y VSS VDD
+ OR2X1_LOC_56/A OR2X1_LOC_53/Y OR2X1_LOC
XAND2X1_LOC_603 AND2X1_LOC_603/a_36_24# OR2X1_LOC_605/B AND2X1_LOC_603/a_8_24# VSS VDD
+ AND2X1_LOC_12/Y OR2X1_LOC_87/A AND2X1_LOC
XAND2X1_LOC_614 AND2X1_LOC_614/a_36_24# OR2X1_LOC_754/A AND2X1_LOC_614/a_8_24# VSS VDD
+ OR2X1_LOC_89/A OR2X1_LOC_427/A AND2X1_LOC
XOR2X1_LOC_78 OR2X1_LOC_78/a_8_216# OR2X1_LOC_78/a_36_216# OR2X1_LOC_78/Y VSS VDD
+ OR2X1_LOC_78/A OR2X1_LOC_78/B OR2X1_LOC
XOR2X1_LOC_23 OR2X1_LOC_23/a_8_216# OR2X1_LOC_23/a_36_216# OR2X1_LOC_45/B VSS VDD
+ OR2X1_LOC_46/A OR2X1_LOC_6/B OR2X1_LOC
XOR2X1_LOC_67 OR2X1_LOC_67/a_8_216# OR2X1_LOC_67/a_36_216# OR2X1_LOC_67/Y VSS VDD
+ OR2X1_LOC_67/A OR2X1_LOC_56/A OR2X1_LOC
XOR2X1_LOC_89 OR2X1_LOC_89/a_8_216# OR2X1_LOC_89/a_36_216# OR2X1_LOC_89/Y VSS VDD
+ OR2X1_LOC_89/A OR2X1_LOC_59/Y OR2X1_LOC
XOR2X1_LOC_34 OR2X1_LOC_34/a_8_216# OR2X1_LOC_34/a_36_216# OR2X1_LOC_35/A VSS VDD
+ OR2X1_LOC_34/A OR2X1_LOC_34/B OR2X1_LOC
XAND2X1_LOC_625 AND2X1_LOC_625/a_36_24# OR2X1_LOC_631/A AND2X1_LOC_625/a_8_24# VSS VDD
+ OR2X1_LOC_66/Y OR2X1_LOC_598/A AND2X1_LOC
XAND2X1_LOC_647 AND2X1_LOC_647/a_36_24# AND2X1_LOC_647/Y AND2X1_LOC_647/a_8_24# VSS VDD
+ OR2X1_LOC_612/Y AND2X1_LOC_647/B AND2X1_LOC
XAND2X1_LOC_669 AND2X1_LOC_669/a_36_24# OR2X1_LOC_720/A AND2X1_LOC_669/a_8_24# VSS VDD
+ OR2X1_LOC_161/A OR2X1_LOC_668/Y AND2X1_LOC
XAND2X1_LOC_636 AND2X1_LOC_636/a_36_24# AND2X1_LOC_639/B AND2X1_LOC_636/a_8_24# VSS VDD
+ OR2X1_LOC_583/Y OR2X1_LOC_584/Y AND2X1_LOC
XAND2X1_LOC_658 AND2X1_LOC_658/a_36_24# AND2X1_LOC_658/Y AND2X1_LOC_658/a_8_24# VSS VDD
+ AND2X1_LOC_658/A AND2X1_LOC_658/B AND2X1_LOC
XAND2X1_LOC_400 AND2X1_LOC_400/a_36_24# AND2X1_LOC_403/B AND2X1_LOC_400/a_8_24# VSS VDD
+ OR2X1_LOC_393/Y OR2X1_LOC_394/Y AND2X1_LOC
XAND2X1_LOC_455 AND2X1_LOC_455/a_36_24# AND2X1_LOC_465/A AND2X1_LOC_455/a_8_24# VSS VDD
+ AND2X1_LOC_76/Y AND2X1_LOC_455/B AND2X1_LOC
XAND2X1_LOC_433 AND2X1_LOC_433/a_36_24# OR2X1_LOC_435/A AND2X1_LOC_433/a_8_24# VSS VDD
+ AND2X1_LOC_70/Y OR2X1_LOC_155/A AND2X1_LOC
XAND2X1_LOC_411 AND2X1_LOC_411/a_36_24# OR2X1_LOC_461/B AND2X1_LOC_411/a_8_24# VSS VDD
+ OR2X1_LOC_756/B OR2X1_LOC_410/Y AND2X1_LOC
XAND2X1_LOC_444 AND2X1_LOC_444/a_36_24# AND2X1_LOC_727/B AND2X1_LOC_444/a_8_24# VSS VDD
+ OR2X1_LOC_442/Y AND2X1_LOC_443/Y AND2X1_LOC
XAND2X1_LOC_422 AND2X1_LOC_422/a_36_24# OR2X1_LOC_448/A AND2X1_LOC_422/a_8_24# VSS VDD
+ AND2X1_LOC_12/Y AND2X1_LOC_92/Y AND2X1_LOC
XOR2X1_LOC_219 OR2X1_LOC_219/a_8_216# OR2X1_LOC_219/a_36_216# OR2X1_LOC_222/A VSS VDD
+ OR2X1_LOC_215/Y OR2X1_LOC_219/B OR2X1_LOC
XOR2X1_LOC_208 OR2X1_LOC_208/a_8_216# OR2X1_LOC_208/a_36_216# OR2X1_LOC_214/A VSS VDD
+ OR2X1_LOC_208/A OR2X1_LOC_35/Y OR2X1_LOC
XAND2X1_LOC_488 AND2X1_LOC_488/a_36_24# OR2X1_LOC_489/A AND2X1_LOC_488/a_8_24# VSS VDD
+ OR2X1_LOC_375/A OR2X1_LOC_814/A AND2X1_LOC
XAND2X1_LOC_499 AND2X1_LOC_499/a_36_24# AND2X1_LOC_500/B AND2X1_LOC_499/a_8_24# VSS VDD
+ OR2X1_LOC_495/Y OR2X1_LOC_496/Y AND2X1_LOC
XAND2X1_LOC_477 AND2X1_LOC_477/a_36_24# AND2X1_LOC_477/Y AND2X1_LOC_477/a_8_24# VSS VDD
+ AND2X1_LOC_477/A AND2X1_LOC_471/Y AND2X1_LOC
XAND2X1_LOC_466 AND2X1_LOC_466/a_36_24# AND2X1_LOC_470/A AND2X1_LOC_466/a_8_24# VSS VDD
+ AND2X1_LOC_453/Y AND2X1_LOC_454/Y AND2X1_LOC
XOR2X1_LOC_764 OR2X1_LOC_764/a_8_216# OR2X1_LOC_764/a_36_216# OR2X1_LOC_764/Y VSS VDD
+ OR2X1_LOC_744/A OR2X1_LOC_40/Y OR2X1_LOC
XOR2X1_LOC_797 OR2X1_LOC_797/a_8_216# OR2X1_LOC_797/a_36_216# OR2X1_LOC_803/A VSS VDD
+ OR2X1_LOC_797/A OR2X1_LOC_797/B OR2X1_LOC
XOR2X1_LOC_731 OR2X1_LOC_731/a_8_216# OR2X1_LOC_731/a_36_216# OR2X1_LOC_738/B VSS VDD
+ OR2X1_LOC_731/A OR2X1_LOC_731/B OR2X1_LOC
XOR2X1_LOC_720 OR2X1_LOC_720/a_8_216# OR2X1_LOC_720/a_36_216# OR2X1_LOC_720/Y VSS VDD
+ OR2X1_LOC_720/A OR2X1_LOC_720/B OR2X1_LOC
XOR2X1_LOC_753 OR2X1_LOC_753/a_8_216# OR2X1_LOC_753/a_36_216# OR2X1_LOC_753/Y VSS VDD
+ OR2X1_LOC_753/A OR2X1_LOC_816/A OR2X1_LOC
XOR2X1_LOC_786 OR2X1_LOC_786/a_8_216# OR2X1_LOC_786/a_36_216# OR2X1_LOC_786/Y VSS VDD
+ OR2X1_LOC_786/A OR2X1_LOC_84/Y OR2X1_LOC
XOR2X1_LOC_742 OR2X1_LOC_742/a_8_216# OR2X1_LOC_742/a_36_216# D_GATE_741 VSS VDD
+ OR2X1_LOC_741/Y OR2X1_LOC_742/B OR2X1_LOC
XOR2X1_LOC_775 OR2X1_LOC_775/a_8_216# OR2X1_LOC_775/a_36_216# OR2X1_LOC_785/B VSS VDD
+ OR2X1_LOC_112/B OR2X1_LOC_97/A OR2X1_LOC
XAND2X1_LOC_230 AND2X1_LOC_230/a_36_24# OR2X1_LOC_231/A AND2X1_LOC_230/a_8_24# VSS VDD
+ AND2X1_LOC_7/B AND2X1_LOC_31/Y AND2X1_LOC
XAND2X1_LOC_252 AND2X1_LOC_252/a_36_24# OR2X1_LOC_254/B AND2X1_LOC_252/a_8_24# VSS VDD
+ AND2X1_LOC_56/B AND2X1_LOC_59/Y AND2X1_LOC
XAND2X1_LOC_263 AND2X1_LOC_263/a_36_24# OR2X1_LOC_266/A AND2X1_LOC_263/a_8_24# VSS VDD
+ AND2X1_LOC_22/Y AND2X1_LOC_42/B AND2X1_LOC
XAND2X1_LOC_285 AND2X1_LOC_285/a_36_24# AND2X1_LOC_285/Y AND2X1_LOC_285/a_8_24# VSS VDD
+ OR2X1_LOC_281/Y OR2X1_LOC_282/Y AND2X1_LOC
XAND2X1_LOC_296 AND2X1_LOC_296/a_36_24# OR2X1_LOC_297/A AND2X1_LOC_296/a_8_24# VSS VDD
+ OR2X1_LOC_43/A OR2X1_LOC_56/A AND2X1_LOC
XAND2X1_LOC_274 AND2X1_LOC_274/a_36_24# OR2X1_LOC_275/A AND2X1_LOC_274/a_8_24# VSS VDD
+ OR2X1_LOC_272/Y OR2X1_LOC_273/Y AND2X1_LOC
XAND2X1_LOC_241 AND2X1_LOC_241/a_36_24# AND2X1_LOC_242/B AND2X1_LOC_241/a_8_24# VSS VDD
+ OR2X1_LOC_237/Y OR2X1_LOC_238/Y AND2X1_LOC
XOR2X1_LOC_583 OR2X1_LOC_583/a_8_216# OR2X1_LOC_583/a_36_216# OR2X1_LOC_583/Y VSS VDD
+ OR2X1_LOC_52/B OR2X1_LOC_31/Y OR2X1_LOC
XOR2X1_LOC_594 OR2X1_LOC_594/a_8_216# OR2X1_LOC_594/a_36_216# OR2X1_LOC_594/Y VSS VDD
+ OR2X1_LOC_680/A OR2X1_LOC_95/Y OR2X1_LOC
XOR2X1_LOC_561 OR2X1_LOC_561/a_8_216# OR2X1_LOC_561/a_36_216# OR2X1_LOC_561/Y VSS VDD
+ OR2X1_LOC_561/A OR2X1_LOC_561/B OR2X1_LOC
XOR2X1_LOC_572 OR2X1_LOC_572/a_8_216# OR2X1_LOC_572/a_36_216# OR2X1_LOC_576/A VSS VDD
+ OR2X1_LOC_267/Y OR2X1_LOC_124/Y OR2X1_LOC
XOR2X1_LOC_550 OR2X1_LOC_550/a_8_216# OR2X1_LOC_550/a_36_216# OR2X1_LOC_565/A VSS VDD
+ OR2X1_LOC_550/A OR2X1_LOC_550/B OR2X1_LOC
XOR2X1_LOC_380 OR2X1_LOC_380/a_8_216# OR2X1_LOC_380/a_36_216# OR2X1_LOC_380/Y VSS VDD
+ OR2X1_LOC_380/A OR2X1_LOC_744/A OR2X1_LOC
XOR2X1_LOC_391 OR2X1_LOC_391/a_8_216# OR2X1_LOC_391/a_36_216# OR2X1_LOC_392/A VSS VDD
+ OR2X1_LOC_391/A OR2X1_LOC_391/B OR2X1_LOC
XAND2X1_LOC_807 AND2X1_LOC_807/a_36_24# AND2X1_LOC_807/Y AND2X1_LOC_807/a_8_24# VSS VDD
+ AND2X1_LOC_805/Y AND2X1_LOC_807/B AND2X1_LOC
XAND2X1_LOC_818 AND2X1_LOC_818/a_36_24# OR2X1_LOC_820/B AND2X1_LOC_818/a_8_24# VSS VDD
+ OR2X1_LOC_6/A OR2X1_LOC_696/A AND2X1_LOC
XAND2X1_LOC_829 AND2X1_LOC_829/a_36_24# OR2X1_LOC_855/A AND2X1_LOC_829/a_8_24# VSS VDD
+ AND2X1_LOC_64/Y OR2X1_LOC_828/Y AND2X1_LOC
XOR2X1_LOC_13 OR2X1_LOC_13/a_8_216# OR2X1_LOC_13/a_36_216# OR2X1_LOC_13/Y VSS VDD
+ OR2X1_LOC_12/Y OR2X1_LOC_13/B OR2X1_LOC
XOR2X1_LOC_35 OR2X1_LOC_35/a_8_216# OR2X1_LOC_35/a_36_216# OR2X1_LOC_35/Y VSS VDD
+ OR2X1_LOC_35/A OR2X1_LOC_35/B OR2X1_LOC
XOR2X1_LOC_46 OR2X1_LOC_46/a_8_216# OR2X1_LOC_46/a_36_216# OR2X1_LOC_48/B VSS VDD
+ OR2X1_LOC_46/A INPUT_1 OR2X1_LOC
XOR2X1_LOC_24 OR2X1_LOC_24/a_8_216# OR2X1_LOC_24/a_36_216# OR2X1_LOC_24/Y VSS VDD
+ OR2X1_LOC_45/B OR2X1_LOC_22/Y OR2X1_LOC
XAND2X1_LOC_604 AND2X1_LOC_604/a_36_24# OR2X1_LOC_605/A AND2X1_LOC_604/a_8_24# VSS VDD
+ AND2X1_LOC_70/Y OR2X1_LOC_161/A AND2X1_LOC
XAND2X1_LOC_626 AND2X1_LOC_626/a_36_24# OR2X1_LOC_629/B AND2X1_LOC_626/a_8_24# VSS VDD
+ AND2X1_LOC_95/Y OR2X1_LOC_161/A AND2X1_LOC
XAND2X1_LOC_637 AND2X1_LOC_637/a_36_24# AND2X1_LOC_637/Y AND2X1_LOC_637/a_8_24# VSS VDD
+ OR2X1_LOC_585/Y OR2X1_LOC_586/Y AND2X1_LOC
XAND2X1_LOC_615 AND2X1_LOC_615/a_36_24# OR2X1_LOC_623/B AND2X1_LOC_615/a_8_24# VSS VDD
+ AND2X1_LOC_22/Y OR2X1_LOC_614/Y AND2X1_LOC
XAND2X1_LOC_648 AND2X1_LOC_648/a_36_24# AND2X1_LOC_655/A AND2X1_LOC_648/a_8_24# VSS VDD
+ AND2X1_LOC_644/Y AND2X1_LOC_648/B AND2X1_LOC
XOR2X1_LOC_68 OR2X1_LOC_68/a_8_216# OR2X1_LOC_68/a_36_216# OR2X1_LOC_68/Y VSS VDD
+ OR2X1_LOC_87/A OR2X1_LOC_68/B OR2X1_LOC
XOR2X1_LOC_79 OR2X1_LOC_79/a_8_216# OR2X1_LOC_79/a_36_216# OR2X1_LOC_79/Y VSS VDD
+ OR2X1_LOC_79/A OR2X1_LOC_18/Y OR2X1_LOC
XOR2X1_LOC_57 OR2X1_LOC_57/a_8_216# OR2X1_LOC_57/a_36_216# OR2X1_LOC_57/Y VSS VDD
+ OR2X1_LOC_44/Y OR2X1_LOC_6/A OR2X1_LOC
XAND2X1_LOC_659 AND2X1_LOC_659/a_36_24# AND2X1_LOC_663/A AND2X1_LOC_659/a_8_24# VSS VDD
+ AND2X1_LOC_657/Y AND2X1_LOC_658/Y AND2X1_LOC
XOR2X1_LOC_209 OR2X1_LOC_209/a_8_216# OR2X1_LOC_209/a_36_216# OR2X1_LOC_213/B VSS VDD
+ OR2X1_LOC_209/A OR2X1_LOC_797/B OR2X1_LOC
XAND2X1_LOC_456 AND2X1_LOC_456/a_36_24# AND2X1_LOC_456/Y AND2X1_LOC_456/a_8_24# VSS VDD
+ OR2X1_LOC_184/Y AND2X1_LOC_456/B AND2X1_LOC
XAND2X1_LOC_489 AND2X1_LOC_489/a_36_24# AND2X1_LOC_489/Y AND2X1_LOC_489/a_8_24# VSS VDD
+ OR2X1_LOC_487/Y OR2X1_LOC_488/Y AND2X1_LOC
XAND2X1_LOC_401 AND2X1_LOC_401/a_36_24# AND2X1_LOC_401/Y AND2X1_LOC_401/a_8_24# VSS VDD
+ OR2X1_LOC_395/Y OR2X1_LOC_396/Y AND2X1_LOC
XAND2X1_LOC_412 AND2X1_LOC_412/a_36_24# OR2X1_LOC_634/A AND2X1_LOC_412/a_8_24# VSS VDD
+ AND2X1_LOC_42/B AND2X1_LOC_44/Y AND2X1_LOC
XAND2X1_LOC_445 AND2X1_LOC_445/a_36_24# AND2X1_LOC_455/B AND2X1_LOC_445/a_8_24# VSS VDD
+ OR2X1_LOC_237/Y OR2X1_LOC_315/Y AND2X1_LOC
XAND2X1_LOC_478 AND2X1_LOC_478/a_36_24# AND2X1_LOC_480/A AND2X1_LOC_478/a_8_24# VSS VDD
+ AND2X1_LOC_469/Y AND2X1_LOC_477/Y AND2X1_LOC
XAND2X1_LOC_434 AND2X1_LOC_434/a_36_24# AND2X1_LOC_434/Y AND2X1_LOC_434/a_8_24# VSS VDD
+ OR2X1_LOC_172/Y OR2X1_LOC_431/Y AND2X1_LOC
XAND2X1_LOC_423 AND2X1_LOC_423/a_36_24# OR2X1_LOC_449/B AND2X1_LOC_423/a_8_24# VSS VDD
+ AND2X1_LOC_7/B AND2X1_LOC_64/Y AND2X1_LOC
XAND2X1_LOC_467 AND2X1_LOC_467/a_36_24# AND2X1_LOC_470/B AND2X1_LOC_467/a_8_24# VSS VDD
+ OR2X1_LOC_163/Y AND2X1_LOC_452/Y AND2X1_LOC
XOR2X1_LOC_710 OR2X1_LOC_710/a_8_216# OR2X1_LOC_710/a_36_216# OR2X1_LOC_711/A VSS VDD
+ OR2X1_LOC_710/A OR2X1_LOC_710/B OR2X1_LOC
XOR2X1_LOC_721 OR2X1_LOC_721/a_8_216# OR2X1_LOC_721/a_36_216# OR2X1_LOC_721/Y VSS VDD
+ OR2X1_LOC_720/Y OR2X1_LOC_673/Y OR2X1_LOC
XOR2X1_LOC_765 OR2X1_LOC_765/a_8_216# OR2X1_LOC_765/a_36_216# OR2X1_LOC_765/Y VSS VDD
+ OR2X1_LOC_16/A OR2X1_LOC_12/Y OR2X1_LOC
XOR2X1_LOC_743 OR2X1_LOC_743/a_8_216# OR2X1_LOC_743/a_36_216# OR2X1_LOC_743/Y VSS VDD
+ OR2X1_LOC_743/A OR2X1_LOC_3/Y OR2X1_LOC
XOR2X1_LOC_732 OR2X1_LOC_732/a_8_216# OR2X1_LOC_732/a_36_216# OR2X1_LOC_738/A VSS VDD
+ OR2X1_LOC_732/A OR2X1_LOC_732/B OR2X1_LOC
XOR2X1_LOC_754 OR2X1_LOC_754/a_8_216# OR2X1_LOC_754/a_36_216# OR2X1_LOC_754/Y VSS VDD
+ OR2X1_LOC_754/A OR2X1_LOC_36/Y OR2X1_LOC
XOR2X1_LOC_787 OR2X1_LOC_787/a_8_216# OR2X1_LOC_787/a_36_216# OR2X1_LOC_787/Y VSS VDD
+ OR2X1_LOC_486/Y OR2X1_LOC_787/B OR2X1_LOC
XOR2X1_LOC_776 OR2X1_LOC_776/a_8_216# OR2X1_LOC_776/a_36_216# OR2X1_LOC_776/Y VSS VDD
+ OR2X1_LOC_776/A OR2X1_LOC_168/B OR2X1_LOC
XOR2X1_LOC_798 OR2X1_LOC_798/a_8_216# OR2X1_LOC_798/a_36_216# OR2X1_LOC_798/Y VSS VDD
+ OR2X1_LOC_436/Y OR2X1_LOC_319/Y OR2X1_LOC
XAND2X1_LOC_242 AND2X1_LOC_242/a_36_24# AND2X1_LOC_244/A AND2X1_LOC_242/a_8_24# VSS VDD
+ OR2X1_LOC_239/Y AND2X1_LOC_242/B AND2X1_LOC
XAND2X1_LOC_275 AND2X1_LOC_275/a_36_24# OR2X1_LOC_276/A AND2X1_LOC_275/a_8_24# VSS VDD
+ D_INPUT_0 OR2X1_LOC_274/Y AND2X1_LOC
XAND2X1_LOC_286 AND2X1_LOC_286/a_36_24# AND2X1_LOC_286/Y AND2X1_LOC_286/a_8_24# VSS VDD
+ OR2X1_LOC_283/Y AND2X1_LOC_285/Y AND2X1_LOC
XAND2X1_LOC_253 AND2X1_LOC_253/a_36_24# OR2X1_LOC_254/A AND2X1_LOC_253/a_8_24# VSS VDD
+ AND2X1_LOC_64/Y OR2X1_LOC_161/B AND2X1_LOC
XAND2X1_LOC_297 AND2X1_LOC_297/a_36_24# OR2X1_LOC_347/B AND2X1_LOC_297/a_8_24# VSS VDD
+ AND2X1_LOC_44/Y OR2X1_LOC_296/Y AND2X1_LOC
XAND2X1_LOC_264 AND2X1_LOC_264/a_36_24# OR2X1_LOC_517/A AND2X1_LOC_264/a_8_24# VSS VDD
+ OR2X1_LOC_13/B OR2X1_LOC_89/A AND2X1_LOC
XAND2X1_LOC_231 AND2X1_LOC_231/a_36_24# AND2X1_LOC_231/Y AND2X1_LOC_231/a_8_24# VSS VDD
+ OR2X1_LOC_229/Y OR2X1_LOC_230/Y AND2X1_LOC
XAND2X1_LOC_220 AND2X1_LOC_220/a_36_24# AND2X1_LOC_220/Y AND2X1_LOC_220/a_8_24# VSS VDD
+ AND2X1_LOC_212/Y AND2X1_LOC_220/B AND2X1_LOC
XOR2X1_LOC_562 OR2X1_LOC_562/a_8_216# OR2X1_LOC_562/a_36_216# OR2X1_LOC_562/Y VSS VDD
+ OR2X1_LOC_562/A OR2X1_LOC_562/B OR2X1_LOC
XOR2X1_LOC_540 OR2X1_LOC_540/a_8_216# OR2X1_LOC_540/a_36_216# OR2X1_LOC_553/B VSS VDD
+ OR2X1_LOC_190/B OR2X1_LOC_181/B OR2X1_LOC
XOR2X1_LOC_551 OR2X1_LOC_551/a_8_216# OR2X1_LOC_551/a_36_216# OR2X1_LOC_564/B VSS VDD
+ OR2X1_LOC_551/A OR2X1_LOC_551/B OR2X1_LOC
XOR2X1_LOC_584 OR2X1_LOC_584/a_8_216# OR2X1_LOC_584/a_36_216# OR2X1_LOC_584/Y VSS VDD
+ OR2X1_LOC_51/Y OR2X1_LOC_7/A OR2X1_LOC
XOR2X1_LOC_573 OR2X1_LOC_573/a_8_216# OR2X1_LOC_573/a_36_216# OR2X1_LOC_573/Y VSS VDD
+ OR2X1_LOC_735/B OR2X1_LOC_404/Y OR2X1_LOC
XOR2X1_LOC_595 OR2X1_LOC_595/a_8_216# OR2X1_LOC_595/a_36_216# OR2X1_LOC_595/Y VSS VDD
+ OR2X1_LOC_595/A OR2X1_LOC_26/Y OR2X1_LOC
XOR2X1_LOC_392 OR2X1_LOC_392/a_8_216# OR2X1_LOC_392/a_36_216# OR2X1_LOC_474/B VSS VDD
+ OR2X1_LOC_392/A OR2X1_LOC_392/B OR2X1_LOC
XOR2X1_LOC_381 OR2X1_LOC_381/a_8_216# OR2X1_LOC_381/a_36_216# OR2X1_LOC_382/A VSS VDD
+ OR2X1_LOC_12/Y D_INPUT_3 OR2X1_LOC
XOR2X1_LOC_370 OR2X1_LOC_370/a_8_216# OR2X1_LOC_370/a_36_216# OR2X1_LOC_787/B VSS VDD
+ OR2X1_LOC_543/A OR2X1_LOC_335/B OR2X1_LOC
XAND2X1_LOC_819 AND2X1_LOC_819/a_36_24# AND2X1_LOC_820/B AND2X1_LOC_819/a_8_24# VSS VDD
+ AND2X1_LOC_47/Y OR2X1_LOC_54/Y AND2X1_LOC
XAND2X1_LOC_808 AND2X1_LOC_808/a_36_24# AND2X1_LOC_811/B AND2X1_LOC_808/a_8_24# VSS VDD
+ AND2X1_LOC_808/A AND2X1_LOC_804/Y AND2X1_LOC
XOR2X1_LOC_25 OR2X1_LOC_25/a_8_216# OR2X1_LOC_25/a_36_216# OR2X1_LOC_25/Y VSS VDD
+ INPUT_7 D_INPUT_6 OR2X1_LOC
XOR2X1_LOC_47 OR2X1_LOC_47/a_8_216# OR2X1_LOC_47/a_36_216# OR2X1_LOC_47/Y VSS VDD
+ OR2X1_LOC_51/B OR2X1_LOC_25/Y OR2X1_LOC
XOR2X1_LOC_36 OR2X1_LOC_36/a_8_216# OR2X1_LOC_36/a_36_216# OR2X1_LOC_36/Y VSS VDD
+ OR2X1_LOC_22/A OR2X1_LOC_17/Y OR2X1_LOC
XOR2X1_LOC_14 OR2X1_LOC_14/a_8_216# OR2X1_LOC_14/a_36_216# OR2X1_LOC_46/A VSS VDD
+ INPUT_3 INPUT_2 OR2X1_LOC
XOR2X1_LOC_58 OR2X1_LOC_58/a_8_216# OR2X1_LOC_58/a_36_216# OR2X1_LOC_58/Y VSS VDD
+ OR2X1_LOC_52/B OR2X1_LOC_22/Y OR2X1_LOC
XOR2X1_LOC_69 OR2X1_LOC_69/a_8_216# OR2X1_LOC_69/a_36_216# OR2X1_LOC_69/Y VSS VDD
+ OR2X1_LOC_69/A OR2X1_LOC_36/Y OR2X1_LOC
XAND2X1_LOC_627 AND2X1_LOC_627/a_36_24# OR2X1_LOC_629/A AND2X1_LOC_627/a_8_24# VSS VDD
+ AND2X1_LOC_7/B AND2X1_LOC_36/Y AND2X1_LOC
XAND2X1_LOC_616 AND2X1_LOC_616/a_36_24# OR2X1_LOC_621/B AND2X1_LOC_616/a_8_24# VSS VDD
+ AND2X1_LOC_18/Y OR2X1_LOC_756/B AND2X1_LOC
XAND2X1_LOC_649 AND2X1_LOC_649/a_36_24# AND2X1_LOC_649/Y AND2X1_LOC_649/a_8_24# VSS VDD
+ AND2X1_LOC_642/Y AND2X1_LOC_649/B AND2X1_LOC
XAND2X1_LOC_638 AND2X1_LOC_638/a_36_24# AND2X1_LOC_638/Y AND2X1_LOC_638/a_8_24# VSS VDD
+ OR2X1_LOC_588/Y AND2X1_LOC_637/Y AND2X1_LOC
XAND2X1_LOC_605 AND2X1_LOC_605/a_36_24# AND2X1_LOC_605/Y AND2X1_LOC_605/a_8_24# VSS VDD
+ OR2X1_LOC_603/Y OR2X1_LOC_604/Y AND2X1_LOC
XAND2X1_LOC_402 AND2X1_LOC_402/a_36_24# AND2X1_LOC_404/A AND2X1_LOC_402/a_8_24# VSS VDD
+ OR2X1_LOC_397/Y AND2X1_LOC_401/Y AND2X1_LOC
XAND2X1_LOC_413 AND2X1_LOC_413/a_36_24# OR2X1_LOC_461/A AND2X1_LOC_413/a_8_24# VSS VDD
+ INPUT_0 OR2X1_LOC_634/A AND2X1_LOC
XAND2X1_LOC_457 AND2X1_LOC_457/a_36_24# AND2X1_LOC_464/A AND2X1_LOC_457/a_8_24# VSS VDD
+ OR2X1_LOC_368/Y AND2X1_LOC_787/A AND2X1_LOC
XAND2X1_LOC_479 AND2X1_LOC_479/a_36_24# AND2X1_LOC_479/Y AND2X1_LOC_479/a_8_24# VSS VDD
+ AND2X1_LOC_475/Y AND2X1_LOC_476/Y AND2X1_LOC
XAND2X1_LOC_468 AND2X1_LOC_468/a_36_24# AND2X1_LOC_469/B AND2X1_LOC_468/a_8_24# VSS VDD
+ AND2X1_LOC_436/Y AND2X1_LOC_468/B AND2X1_LOC
XAND2X1_LOC_424 AND2X1_LOC_424/a_36_24# OR2X1_LOC_449/A AND2X1_LOC_424/a_8_24# VSS VDD
+ AND2X1_LOC_44/Y OR2X1_LOC_78/A AND2X1_LOC
XAND2X1_LOC_435 AND2X1_LOC_435/a_36_24# AND2X1_LOC_436/B AND2X1_LOC_435/a_8_24# VSS VDD
+ OR2X1_LOC_432/Y OR2X1_LOC_433/Y AND2X1_LOC
XAND2X1_LOC_446 AND2X1_LOC_446/a_36_24# AND2X1_LOC_454/A AND2X1_LOC_446/a_8_24# VSS VDD
+ OR2X1_LOC_417/Y OR2X1_LOC_418/Y AND2X1_LOC
XOR2X1_LOC_744 OR2X1_LOC_744/a_8_216# OR2X1_LOC_744/a_36_216# OR2X1_LOC_744/Y VSS VDD
+ OR2X1_LOC_744/A OR2X1_LOC_44/Y OR2X1_LOC
XOR2X1_LOC_711 OR2X1_LOC_711/a_8_216# OR2X1_LOC_711/a_36_216# OR2X1_LOC_726/A VSS VDD
+ OR2X1_LOC_711/A OR2X1_LOC_711/B OR2X1_LOC
XOR2X1_LOC_700 OR2X1_LOC_700/a_8_216# OR2X1_LOC_700/a_36_216# OR2X1_LOC_700/Y VSS VDD
+ OR2X1_LOC_91/A OR2X1_LOC_59/Y OR2X1_LOC
XOR2X1_LOC_733 OR2X1_LOC_733/a_8_216# OR2X1_LOC_733/a_36_216# OR2X1_LOC_733/Y VSS VDD
+ OR2X1_LOC_733/A OR2X1_LOC_733/B OR2X1_LOC
XOR2X1_LOC_722 OR2X1_LOC_722/a_8_216# OR2X1_LOC_722/a_36_216# OR2X1_LOC_733/B VSS VDD
+ OR2X1_LOC_719/Y OR2X1_LOC_722/B OR2X1_LOC
XOR2X1_LOC_766 OR2X1_LOC_766/a_8_216# OR2X1_LOC_766/a_36_216# OR2X1_LOC_766/Y VSS VDD
+ OR2X1_LOC_91/A OR2X1_LOC_64/Y OR2X1_LOC
XOR2X1_LOC_777 OR2X1_LOC_777/a_8_216# OR2X1_LOC_777/a_36_216# OR2X1_LOC_784/B VSS VDD
+ OR2X1_LOC_307/A OR2X1_LOC_777/B OR2X1_LOC
XOR2X1_LOC_755 OR2X1_LOC_755/a_8_216# OR2X1_LOC_755/a_36_216# OR2X1_LOC_755/Y VSS VDD
+ OR2X1_LOC_755/A OR2X1_LOC_59/Y OR2X1_LOC
XOR2X1_LOC_788 OR2X1_LOC_788/a_8_216# OR2X1_LOC_788/a_36_216# OR2X1_LOC_794/A VSS VDD
+ OR2X1_LOC_602/Y OR2X1_LOC_788/B OR2X1_LOC
XOR2X1_LOC_799 OR2X1_LOC_799/a_8_216# OR2X1_LOC_799/a_36_216# OR2X1_LOC_802/A VSS VDD
+ OR2X1_LOC_799/A OR2X1_LOC_539/Y OR2X1_LOC
XAND2X1_LOC_221 AND2X1_LOC_221/a_36_24# AND2X1_LOC_223/A AND2X1_LOC_221/a_8_24# VSS VDD
+ AND2X1_LOC_192/Y AND2X1_LOC_220/Y AND2X1_LOC
XAND2X1_LOC_210 AND2X1_LOC_210/a_36_24# AND2X1_LOC_213/B AND2X1_LOC_210/a_8_24# VSS VDD
+ OR2X1_LOC_158/Y OR2X1_LOC_163/Y AND2X1_LOC
XAND2X1_LOC_265 AND2X1_LOC_265/a_36_24# OR2X1_LOC_641/A AND2X1_LOC_265/a_8_24# VSS VDD
+ AND2X1_LOC_40/Y OR2X1_LOC_264/Y AND2X1_LOC
XAND2X1_LOC_232 AND2X1_LOC_232/a_36_24# OR2X1_LOC_240/B AND2X1_LOC_232/a_8_24# VSS VDD
+ OR2X1_LOC_78/B OR2X1_LOC_375/A AND2X1_LOC
XAND2X1_LOC_287 AND2X1_LOC_287/a_36_24# AND2X1_LOC_287/Y AND2X1_LOC_287/a_8_24# VSS VDD
+ OR2X1_LOC_278/Y AND2X1_LOC_287/B AND2X1_LOC
XAND2X1_LOC_243 AND2X1_LOC_243/a_36_24# AND2X1_LOC_243/Y AND2X1_LOC_243/a_8_24# VSS VDD
+ OR2X1_LOC_235/Y AND2X1_LOC_240/Y AND2X1_LOC
XAND2X1_LOC_254 AND2X1_LOC_254/a_36_24# AND2X1_LOC_456/B AND2X1_LOC_254/a_8_24# VSS VDD
+ OR2X1_LOC_252/Y OR2X1_LOC_253/Y AND2X1_LOC
XAND2X1_LOC_276 AND2X1_LOC_276/a_36_24# AND2X1_LOC_276/Y AND2X1_LOC_276/a_8_24# VSS VDD
+ OR2X1_LOC_271/Y OR2X1_LOC_275/Y AND2X1_LOC
XAND2X1_LOC_298 AND2X1_LOC_298/a_36_24# OR2X1_LOC_302/B AND2X1_LOC_298/a_8_24# VSS VDD
+ AND2X1_LOC_31/Y AND2X1_LOC_56/B AND2X1_LOC
XOR2X1_LOC_585 OR2X1_LOC_585/a_8_216# OR2X1_LOC_585/a_36_216# OR2X1_LOC_585/Y VSS VDD
+ OR2X1_LOC_585/A OR2X1_LOC_22/Y OR2X1_LOC
XOR2X1_LOC_596 OR2X1_LOC_596/a_8_216# OR2X1_LOC_596/a_36_216# OR2X1_LOC_596/Y VSS VDD
+ OR2X1_LOC_596/A AND2X1_LOC_44/Y OR2X1_LOC
XOR2X1_LOC_563 OR2X1_LOC_563/a_8_216# OR2X1_LOC_563/a_36_216# OR2X1_LOC_570/A VSS VDD
+ OR2X1_LOC_563/A OR2X1_LOC_563/B OR2X1_LOC
XOR2X1_LOC_574 OR2X1_LOC_574/a_8_216# OR2X1_LOC_574/a_36_216# OR2X1_LOC_575/A VSS VDD
+ OR2X1_LOC_574/A OR2X1_LOC_510/Y OR2X1_LOC
XOR2X1_LOC_541 OR2X1_LOC_541/a_8_216# OR2X1_LOC_541/a_36_216# OR2X1_LOC_553/A VSS VDD
+ OR2X1_LOC_541/A OR2X1_LOC_541/B OR2X1_LOC
XOR2X1_LOC_552 OR2X1_LOC_552/a_8_216# OR2X1_LOC_552/a_36_216# OR2X1_LOC_564/A VSS VDD
+ OR2X1_LOC_552/A OR2X1_LOC_552/B OR2X1_LOC
XOR2X1_LOC_530 OR2X1_LOC_530/a_8_216# OR2X1_LOC_530/a_36_216# OR2X1_LOC_530/Y VSS VDD
+ OR2X1_LOC_485/A OR2X1_LOC_36/Y OR2X1_LOC
XOR2X1_LOC_382 OR2X1_LOC_382/a_8_216# OR2X1_LOC_382/a_36_216# OR2X1_LOC_382/Y VSS VDD
+ OR2X1_LOC_382/A OR2X1_LOC_49/A OR2X1_LOC
XOR2X1_LOC_360 OR2X1_LOC_360/a_8_216# OR2X1_LOC_360/a_36_216# OR2X1_LOC_363/A VSS VDD
+ OR2X1_LOC_347/Y OR2X1_LOC_244/Y OR2X1_LOC
XOR2X1_LOC_393 OR2X1_LOC_393/a_8_216# OR2X1_LOC_393/a_36_216# OR2X1_LOC_393/Y VSS VDD
+ OR2X1_LOC_40/Y OR2X1_LOC_39/A OR2X1_LOC
XOR2X1_LOC_371 OR2X1_LOC_371/a_8_216# OR2X1_LOC_371/a_36_216# OR2X1_LOC_371/Y VSS VDD
+ OR2X1_LOC_31/Y OR2X1_LOC_6/A OR2X1_LOC
XAND2X1_LOC_809 AND2X1_LOC_809/a_36_24# AND2X1_LOC_810/B AND2X1_LOC_809/a_8_24# VSS VDD
+ AND2X1_LOC_809/A AND2X1_LOC_802/Y AND2X1_LOC
XOR2X1_LOC_190 OR2X1_LOC_190/a_8_216# OR2X1_LOC_190/a_36_216# OR2X1_LOC_190/Y VSS VDD
+ OR2X1_LOC_190/A OR2X1_LOC_190/B OR2X1_LOC
XOR2X1_LOC_26 OR2X1_LOC_26/a_8_216# OR2X1_LOC_26/a_36_216# OR2X1_LOC_26/Y VSS VDD
+ OR2X1_LOC_25/Y OR2X1_LOC_22/A OR2X1_LOC
XOR2X1_LOC_59 OR2X1_LOC_59/a_8_216# OR2X1_LOC_59/a_36_216# OR2X1_LOC_59/Y VSS VDD
+ OR2X1_LOC_25/Y OR2X1_LOC_11/Y OR2X1_LOC
XOR2X1_LOC_48 OR2X1_LOC_48/a_8_216# OR2X1_LOC_48/a_36_216# OR2X1_LOC_48/Y VSS VDD
+ OR2X1_LOC_47/Y OR2X1_LOC_48/B OR2X1_LOC
XOR2X1_LOC_37 OR2X1_LOC_37/a_8_216# OR2X1_LOC_37/a_36_216# OR2X1_LOC_85/A VSS VDD
+ D_INPUT_3 D_INPUT_2 OR2X1_LOC
XOR2X1_LOC_15 OR2X1_LOC_15/a_8_216# OR2X1_LOC_15/a_36_216# OR2X1_LOC_16/A VSS VDD
+ OR2X1_LOC_46/A OR2X1_LOC_9/Y OR2X1_LOC
XAND2X1_LOC_606 AND2X1_LOC_606/a_36_24# OR2X1_LOC_607/A AND2X1_LOC_606/a_8_24# VSS VDD
+ OR2X1_LOC_485/A OR2X1_LOC_426/B AND2X1_LOC
XAND2X1_LOC_628 AND2X1_LOC_628/a_36_24# OR2X1_LOC_630/B AND2X1_LOC_628/a_8_24# VSS VDD
+ AND2X1_LOC_47/Y AND2X1_LOC_92/Y AND2X1_LOC
XAND2X1_LOC_617 AND2X1_LOC_617/a_36_24# OR2X1_LOC_621/A AND2X1_LOC_617/a_8_24# VSS VDD
+ OR2X1_LOC_154/A AND2X1_LOC_51/Y AND2X1_LOC
XAND2X1_LOC_639 AND2X1_LOC_639/a_36_24# AND2X1_LOC_651/B AND2X1_LOC_639/a_8_24# VSS VDD
+ AND2X1_LOC_639/A AND2X1_LOC_639/B AND2X1_LOC
XAND2X1_LOC_403 AND2X1_LOC_403/a_36_24# AND2X1_LOC_404/B AND2X1_LOC_403/a_8_24# VSS VDD
+ OR2X1_LOC_399/Y AND2X1_LOC_403/B AND2X1_LOC
XAND2X1_LOC_414 AND2X1_LOC_414/a_36_24# OR2X1_LOC_415/A AND2X1_LOC_414/a_8_24# VSS VDD
+ INPUT_3 OR2X1_LOC_19/B AND2X1_LOC
XAND2X1_LOC_458 AND2X1_LOC_458/a_36_24# AND2X1_LOC_458/Y AND2X1_LOC_458/a_8_24# VSS VDD
+ OR2X1_LOC_372/Y AND2X1_LOC_374/Y AND2X1_LOC
XAND2X1_LOC_469 AND2X1_LOC_469/a_36_24# AND2X1_LOC_469/Y AND2X1_LOC_469/a_8_24# VSS VDD
+ AND2X1_LOC_727/B AND2X1_LOC_469/B AND2X1_LOC
XAND2X1_LOC_436 AND2X1_LOC_436/a_36_24# AND2X1_LOC_436/Y AND2X1_LOC_436/a_8_24# VSS VDD
+ AND2X1_LOC_434/Y AND2X1_LOC_436/B AND2X1_LOC
XAND2X1_LOC_447 AND2X1_LOC_447/a_36_24# AND2X1_LOC_447/Y AND2X1_LOC_447/a_8_24# VSS VDD
+ OR2X1_LOC_419/Y OR2X1_LOC_420/Y AND2X1_LOC
XAND2X1_LOC_425 AND2X1_LOC_425/a_36_24# AND2X1_LOC_425/Y AND2X1_LOC_425/a_8_24# VSS VDD
+ D_INPUT_5 AND2X1_LOC_17/Y AND2X1_LOC
XOR2X1_LOC_745 OR2X1_LOC_745/a_8_216# OR2X1_LOC_745/a_36_216# OR2X1_LOC_745/Y VSS VDD
+ OR2X1_LOC_604/A OR2X1_LOC_40/Y OR2X1_LOC
XOR2X1_LOC_712 OR2X1_LOC_712/a_8_216# OR2X1_LOC_712/a_36_216# OR2X1_LOC_725/B VSS VDD
+ OR2X1_LOC_708/Y OR2X1_LOC_712/B OR2X1_LOC
XOR2X1_LOC_701 OR2X1_LOC_701/a_8_216# OR2X1_LOC_701/a_36_216# OR2X1_LOC_701/Y VSS VDD
+ OR2X1_LOC_428/A OR2X1_LOC_44/Y OR2X1_LOC
XOR2X1_LOC_756 OR2X1_LOC_756/a_8_216# OR2X1_LOC_756/a_36_216# OR2X1_LOC_756/Y VSS VDD
+ OR2X1_LOC_161/A OR2X1_LOC_756/B OR2X1_LOC
XOR2X1_LOC_723 OR2X1_LOC_723/a_8_216# OR2X1_LOC_723/a_36_216# OR2X1_LOC_733/A VSS VDD
+ OR2X1_LOC_723/A OR2X1_LOC_723/B OR2X1_LOC
XOR2X1_LOC_778 OR2X1_LOC_778/a_8_216# OR2X1_LOC_778/a_36_216# OR2X1_LOC_778/Y VSS VDD
+ OR2X1_LOC_778/A OR2X1_LOC_778/B OR2X1_LOC
XOR2X1_LOC_734 OR2X1_LOC_734/a_8_216# OR2X1_LOC_734/a_36_216# OR2X1_LOC_737/A VSS VDD
+ OR2X1_LOC_721/Y OR2X1_LOC_475/B OR2X1_LOC
XOR2X1_LOC_767 OR2X1_LOC_767/a_8_216# OR2X1_LOC_767/a_36_216# OR2X1_LOC_767/Y VSS VDD
+ OR2X1_LOC_79/A OR2X1_LOC_3/Y OR2X1_LOC
XOR2X1_LOC_789 OR2X1_LOC_789/a_8_216# OR2X1_LOC_789/a_36_216# OR2X1_LOC_793/B VSS VDD
+ OR2X1_LOC_789/A OR2X1_LOC_789/B OR2X1_LOC
XAND2X1_LOC_255 AND2X1_LOC_255/a_36_24# OR2X1_LOC_541/B AND2X1_LOC_255/a_8_24# VSS VDD
+ AND2X1_LOC_42/B OR2X1_LOC_375/A AND2X1_LOC
XAND2X1_LOC_244 AND2X1_LOC_244/a_36_24# AND2X1_LOC_860/A AND2X1_LOC_244/a_8_24# VSS VDD
+ AND2X1_LOC_244/A AND2X1_LOC_243/Y AND2X1_LOC
XAND2X1_LOC_222 AND2X1_LOC_222/a_36_24# AND2X1_LOC_222/Y AND2X1_LOC_222/a_8_24# VSS VDD
+ AND2X1_LOC_218/Y AND2X1_LOC_219/Y AND2X1_LOC
XAND2X1_LOC_233 AND2X1_LOC_233/a_36_24# AND2X1_LOC_824/B AND2X1_LOC_233/a_8_24# VSS VDD
+ INPUT_0 OR2X1_LOC_377/A AND2X1_LOC
XAND2X1_LOC_211 AND2X1_LOC_211/a_36_24# AND2X1_LOC_212/B AND2X1_LOC_211/a_8_24# VSS VDD
+ AND2X1_LOC_170/Y AND2X1_LOC_211/B AND2X1_LOC
XAND2X1_LOC_200 AND2X1_LOC_200/a_36_24# AND2X1_LOC_207/B AND2X1_LOC_200/a_8_24# VSS VDD
+ AND2X1_LOC_193/Y AND2X1_LOC_194/Y AND2X1_LOC
XAND2X1_LOC_266 AND2X1_LOC_266/a_36_24# AND2X1_LOC_266/Y AND2X1_LOC_266/a_8_24# VSS VDD
+ OR2X1_LOC_262/Y OR2X1_LOC_813/A AND2X1_LOC
XAND2X1_LOC_288 AND2X1_LOC_288/a_36_24# AND2X1_LOC_806/A AND2X1_LOC_288/a_8_24# VSS VDD
+ AND2X1_LOC_286/Y AND2X1_LOC_287/Y AND2X1_LOC
XAND2X1_LOC_277 AND2X1_LOC_277/a_36_24# OR2X1_LOC_633/A AND2X1_LOC_277/a_8_24# VSS VDD
+ AND2X1_LOC_42/B AND2X1_LOC_47/Y AND2X1_LOC
XAND2X1_LOC_299 AND2X1_LOC_299/a_36_24# OR2X1_LOC_302/A AND2X1_LOC_299/a_8_24# VSS VDD
+ AND2X1_LOC_12/Y OR2X1_LOC_121/B AND2X1_LOC
XOR2X1_LOC_597 OR2X1_LOC_597/a_8_216# OR2X1_LOC_597/a_36_216# OR2X1_LOC_597/Y VSS VDD
+ OR2X1_LOC_597/A OR2X1_LOC_13/B OR2X1_LOC
XOR2X1_LOC_586 OR2X1_LOC_586/a_8_216# OR2X1_LOC_586/a_36_216# OR2X1_LOC_586/Y VSS VDD
+ OR2X1_LOC_589/A OR2X1_LOC_70/Y OR2X1_LOC
XOR2X1_LOC_575 OR2X1_LOC_575/a_8_216# OR2X1_LOC_575/a_36_216# OR2X1_LOC_579/B VSS VDD
+ OR2X1_LOC_575/A OR2X1_LOC_573/Y OR2X1_LOC
XOR2X1_LOC_553 OR2X1_LOC_553/a_8_216# OR2X1_LOC_553/a_36_216# OR2X1_LOC_563/B VSS VDD
+ OR2X1_LOC_553/A OR2X1_LOC_553/B OR2X1_LOC
XOR2X1_LOC_564 OR2X1_LOC_564/a_8_216# OR2X1_LOC_564/a_36_216# OR2X1_LOC_569/B VSS VDD
+ OR2X1_LOC_564/A OR2X1_LOC_564/B OR2X1_LOC
XOR2X1_LOC_542 OR2X1_LOC_542/a_8_216# OR2X1_LOC_542/a_36_216# OR2X1_LOC_552/B VSS VDD
+ OR2X1_LOC_703/A OR2X1_LOC_542/B OR2X1_LOC
XOR2X1_LOC_520 OR2X1_LOC_520/a_8_216# OR2X1_LOC_520/a_36_216# OR2X1_LOC_520/Y VSS VDD
+ OR2X1_LOC_520/A OR2X1_LOC_520/B OR2X1_LOC
XOR2X1_LOC_531 OR2X1_LOC_531/a_8_216# OR2X1_LOC_531/a_36_216# OR2X1_LOC_531/Y VSS VDD
+ OR2X1_LOC_74/A OR2X1_LOC_40/Y OR2X1_LOC
XOR2X1_LOC_383 OR2X1_LOC_383/a_8_216# OR2X1_LOC_383/a_36_216# OR2X1_LOC_383/Y VSS VDD
+ OR2X1_LOC_269/B AND2X1_LOC_91/B OR2X1_LOC
XOR2X1_LOC_361 OR2X1_LOC_361/a_8_216# OR2X1_LOC_361/a_36_216# OR2X1_LOC_362/A VSS VDD
+ OR2X1_LOC_473/A OR2X1_LOC_267/Y OR2X1_LOC
XOR2X1_LOC_394 OR2X1_LOC_394/a_8_216# OR2X1_LOC_394/a_36_216# OR2X1_LOC_394/Y VSS VDD
+ OR2X1_LOC_744/A OR2X1_LOC_47/Y OR2X1_LOC
XOR2X1_LOC_350 OR2X1_LOC_350/a_8_216# OR2X1_LOC_350/a_36_216# OR2X1_LOC_358/B VSS VDD
+ OR2X1_LOC_341/Y OR2X1_LOC_340/Y OR2X1_LOC
XOR2X1_LOC_372 OR2X1_LOC_372/a_8_216# OR2X1_LOC_372/a_36_216# OR2X1_LOC_372/Y VSS VDD
+ OR2X1_LOC_371/Y INPUT_1 OR2X1_LOC
XOR2X1_LOC_180 OR2X1_LOC_180/a_8_216# OR2X1_LOC_180/a_36_216# OR2X1_LOC_182/B VSS VDD
+ OR2X1_LOC_439/B OR2X1_LOC_180/B OR2X1_LOC
XOR2X1_LOC_191 OR2X1_LOC_191/a_8_216# OR2X1_LOC_191/a_36_216# OR2X1_LOC_192/A VSS VDD
+ OR2X1_LOC_190/Y OR2X1_LOC_191/B OR2X1_LOC
XOR2X1_LOC_16 OR2X1_LOC_16/a_8_216# OR2X1_LOC_16/a_36_216# OR2X1_LOC_16/Y VSS VDD
+ OR2X1_LOC_16/A OR2X1_LOC_3/Y OR2X1_LOC
XOR2X1_LOC_38 OR2X1_LOC_38/a_8_216# OR2X1_LOC_38/a_36_216# OR2X1_LOC_39/A VSS VDD
+ OR2X1_LOC_85/A OR2X1_LOC_49/A OR2X1_LOC
XOR2X1_LOC_49 OR2X1_LOC_49/a_8_216# OR2X1_LOC_49/a_36_216# OR2X1_LOC_52/B VSS VDD
+ OR2X1_LOC_49/A OR2X1_LOC_46/A OR2X1_LOC
XOR2X1_LOC_27 OR2X1_LOC_27/a_8_216# OR2X1_LOC_27/a_36_216# OR2X1_LOC_27/Y VSS VDD
+ OR2X1_LOC_26/Y OR2X1_LOC_7/A OR2X1_LOC
XAND2X1_LOC_607 AND2X1_LOC_607/a_36_24# OR2X1_LOC_646/B AND2X1_LOC_607/a_8_24# VSS VDD
+ AND2X1_LOC_18/Y OR2X1_LOC_606/Y AND2X1_LOC
XAND2X1_LOC_629 AND2X1_LOC_629/a_36_24# AND2X1_LOC_629/Y AND2X1_LOC_629/a_8_24# VSS VDD
+ OR2X1_LOC_626/Y OR2X1_LOC_627/Y AND2X1_LOC
XAND2X1_LOC_618 AND2X1_LOC_618/a_36_24# AND2X1_LOC_619/B AND2X1_LOC_618/a_8_24# VSS VDD
+ D_INPUT_3 OR2X1_LOC_80/A AND2X1_LOC
XAND2X1_LOC_404 AND2X1_LOC_404/a_36_24# AND2X1_LOC_573/A AND2X1_LOC_404/a_8_24# VSS VDD
+ AND2X1_LOC_404/A AND2X1_LOC_404/B AND2X1_LOC
XAND2X1_LOC_415 AND2X1_LOC_415/a_36_24# OR2X1_LOC_416/A AND2X1_LOC_415/a_8_24# VSS VDD
+ OR2X1_LOC_585/A OR2X1_LOC_414/Y AND2X1_LOC
XAND2X1_LOC_437 AND2X1_LOC_437/a_36_24# OR2X1_LOC_440/B AND2X1_LOC_437/a_8_24# VSS VDD
+ AND2X1_LOC_59/Y OR2X1_LOC_151/A AND2X1_LOC
XAND2X1_LOC_426 AND2X1_LOC_426/a_36_24# OR2X1_LOC_450/B AND2X1_LOC_426/a_8_24# VSS VDD
+ OR2X1_LOC_121/B AND2X1_LOC_425/Y AND2X1_LOC
XAND2X1_LOC_459 AND2X1_LOC_459/a_36_24# AND2X1_LOC_459/Y AND2X1_LOC_459/a_8_24# VSS VDD
+ OR2X1_LOC_376/Y OR2X1_LOC_378/Y AND2X1_LOC
XAND2X1_LOC_448 AND2X1_LOC_448/a_36_24# AND2X1_LOC_448/Y AND2X1_LOC_448/a_8_24# VSS VDD
+ OR2X1_LOC_421/Y OR2X1_LOC_422/Y AND2X1_LOC
XOR2X1_LOC_746 OR2X1_LOC_746/a_8_216# OR2X1_LOC_746/a_36_216# OR2X1_LOC_746/Y VSS VDD
+ OR2X1_LOC_158/A OR2X1_LOC_74/A OR2X1_LOC
XOR2X1_LOC_779 OR2X1_LOC_779/a_8_216# OR2X1_LOC_779/a_36_216# OR2X1_LOC_779/Y VSS VDD
+ OR2X1_LOC_779/A OR2X1_LOC_779/B OR2X1_LOC
XOR2X1_LOC_713 OR2X1_LOC_713/a_8_216# OR2X1_LOC_713/a_36_216# OR2X1_LOC_725/A VSS VDD
+ OR2X1_LOC_713/A OR2X1_LOC_705/Y OR2X1_LOC
XOR2X1_LOC_702 OR2X1_LOC_702/a_8_216# OR2X1_LOC_702/a_36_216# OR2X1_LOC_715/A VSS VDD
+ OR2X1_LOC_702/A OR2X1_LOC_196/B OR2X1_LOC
XOR2X1_LOC_724 OR2X1_LOC_724/a_8_216# OR2X1_LOC_724/a_36_216# OR2X1_LOC_732/B VSS VDD
+ OR2X1_LOC_724/A OR2X1_LOC_714/Y OR2X1_LOC
XOR2X1_LOC_757 OR2X1_LOC_757/a_8_216# OR2X1_LOC_757/a_36_216# OR2X1_LOC_757/Y VSS VDD
+ OR2X1_LOC_757/A OR2X1_LOC_44/Y OR2X1_LOC
XOR2X1_LOC_768 OR2X1_LOC_768/a_8_216# OR2X1_LOC_768/a_36_216# OR2X1_LOC_772/A VSS VDD
+ OR2X1_LOC_768/A OR2X1_LOC_113/B OR2X1_LOC
XOR2X1_LOC_735 OR2X1_LOC_735/a_8_216# OR2X1_LOC_735/a_36_216# OR2X1_LOC_736/A VSS VDD
+ OR2X1_LOC_632/Y OR2X1_LOC_735/B OR2X1_LOC
XAND2X1_LOC_267 AND2X1_LOC_267/a_36_24# AND2X1_LOC_361/A AND2X1_LOC_267/a_8_24# VSS VDD
+ OR2X1_LOC_265/Y AND2X1_LOC_266/Y AND2X1_LOC
XAND2X1_LOC_256 AND2X1_LOC_256/a_36_24# OR2X1_LOC_344/A AND2X1_LOC_256/a_8_24# VSS VDD
+ OR2X1_LOC_6/B OR2X1_LOC_541/B AND2X1_LOC
XAND2X1_LOC_245 AND2X1_LOC_245/a_36_24# OR2X1_LOC_777/B AND2X1_LOC_245/a_8_24# VSS VDD
+ OR2X1_LOC_66/A AND2X1_LOC_42/B AND2X1_LOC
XAND2X1_LOC_278 AND2X1_LOC_278/a_36_24# OR2X1_LOC_287/B AND2X1_LOC_278/a_8_24# VSS VDD
+ OR2X1_LOC_9/Y OR2X1_LOC_633/A AND2X1_LOC
XAND2X1_LOC_234 AND2X1_LOC_234/a_36_24# OR2X1_LOC_240/A AND2X1_LOC_234/a_8_24# VSS VDD
+ AND2X1_LOC_47/Y AND2X1_LOC_824/B AND2X1_LOC
XAND2X1_LOC_201 AND2X1_LOC_201/a_36_24# AND2X1_LOC_201/Y AND2X1_LOC_201/a_8_24# VSS VDD
+ AND2X1_LOC_61/Y OR2X1_LOC_65/Y AND2X1_LOC
XAND2X1_LOC_289 AND2X1_LOC_289/a_36_24# OR2X1_LOC_333/A AND2X1_LOC_289/a_8_24# VSS VDD
+ AND2X1_LOC_51/Y OR2X1_LOC_814/A AND2X1_LOC
XAND2X1_LOC_223 AND2X1_LOC_223/a_36_24# GATE_222 AND2X1_LOC_223/a_8_24# VSS VDD
+ AND2X1_LOC_223/A AND2X1_LOC_222/Y AND2X1_LOC
XAND2X1_LOC_212 AND2X1_LOC_212/a_36_24# AND2X1_LOC_212/Y AND2X1_LOC_212/a_8_24# VSS VDD
+ AND2X1_LOC_212/A AND2X1_LOC_212/B AND2X1_LOC
XOR2X1_LOC_510 OR2X1_LOC_510/a_8_216# OR2X1_LOC_510/a_36_216# OR2X1_LOC_510/Y VSS VDD
+ OR2X1_LOC_510/A OR2X1_LOC_508/Y OR2X1_LOC
XOR2X1_LOC_587 OR2X1_LOC_587/a_8_216# OR2X1_LOC_587/a_36_216# OR2X1_LOC_588/A VSS VDD
+ OR2X1_LOC_51/B INPUT_7 OR2X1_LOC
XAND2X1_LOC_790 AND2X1_LOC_790/a_36_24# AND2X1_LOC_793/B AND2X1_LOC_790/a_8_24# VSS VDD
+ OR2X1_LOC_753/Y OR2X1_LOC_754/Y AND2X1_LOC
XOR2X1_LOC_576 OR2X1_LOC_576/a_8_216# OR2X1_LOC_576/a_36_216# OR2X1_LOC_579/A VSS VDD
+ OR2X1_LOC_576/A OR2X1_LOC_571/Y OR2X1_LOC
XOR2X1_LOC_554 OR2X1_LOC_554/a_8_216# OR2X1_LOC_554/a_36_216# OR2X1_LOC_563/A VSS VDD
+ OR2X1_LOC_140/B OR2X1_LOC_115/B OR2X1_LOC
XOR2X1_LOC_565 OR2X1_LOC_565/a_8_216# OR2X1_LOC_565/a_36_216# OR2X1_LOC_569/A VSS VDD
+ OR2X1_LOC_565/A OR2X1_LOC_549/Y OR2X1_LOC
XOR2X1_LOC_543 OR2X1_LOC_543/a_8_216# OR2X1_LOC_543/a_36_216# OR2X1_LOC_552/A VSS VDD
+ OR2X1_LOC_543/A OR2X1_LOC_318/B OR2X1_LOC
XOR2X1_LOC_521 OR2X1_LOC_521/a_8_216# OR2X1_LOC_521/a_36_216# OR2X1_LOC_521/Y VSS VDD
+ OR2X1_LOC_52/B OR2X1_LOC_18/Y OR2X1_LOC
XOR2X1_LOC_532 OR2X1_LOC_532/a_8_216# OR2X1_LOC_532/a_36_216# OR2X1_LOC_532/Y VSS VDD
+ OR2X1_LOC_160/A OR2X1_LOC_532/B OR2X1_LOC
XOR2X1_LOC_598 OR2X1_LOC_598/a_8_216# OR2X1_LOC_598/a_36_216# OR2X1_LOC_598/Y VSS VDD
+ OR2X1_LOC_598/A AND2X1_LOC_48/A OR2X1_LOC
XOR2X1_LOC_362 OR2X1_LOC_362/a_8_216# OR2X1_LOC_362/a_36_216# OR2X1_LOC_366/B VSS VDD
+ OR2X1_LOC_362/A OR2X1_LOC_362/B OR2X1_LOC
XOR2X1_LOC_340 OR2X1_LOC_340/a_8_216# OR2X1_LOC_340/a_36_216# OR2X1_LOC_340/Y VSS VDD
+ OR2X1_LOC_227/Y AND2X1_LOC_88/Y OR2X1_LOC
XOR2X1_LOC_351 OR2X1_LOC_351/a_8_216# OR2X1_LOC_351/a_36_216# OR2X1_LOC_358/A VSS VDD
+ OR2X1_LOC_339/Y OR2X1_LOC_351/B OR2X1_LOC
XOR2X1_LOC_384 OR2X1_LOC_384/a_8_216# OR2X1_LOC_384/a_36_216# OR2X1_LOC_384/Y VSS VDD
+ OR2X1_LOC_494/A OR2X1_LOC_40/Y OR2X1_LOC
XOR2X1_LOC_395 OR2X1_LOC_395/a_8_216# OR2X1_LOC_395/a_36_216# OR2X1_LOC_395/Y VSS VDD
+ OR2X1_LOC_600/A OR2X1_LOC_59/Y OR2X1_LOC
XOR2X1_LOC_373 OR2X1_LOC_373/a_8_216# OR2X1_LOC_373/a_36_216# OR2X1_LOC_373/Y VSS VDD
+ OR2X1_LOC_89/A OR2X1_LOC_26/Y OR2X1_LOC
XOR2X1_LOC_192 OR2X1_LOC_192/a_8_216# OR2X1_LOC_192/a_36_216# OR2X1_LOC_739/B VSS VDD
+ OR2X1_LOC_192/A OR2X1_LOC_192/B OR2X1_LOC
XOR2X1_LOC_181 OR2X1_LOC_181/a_8_216# OR2X1_LOC_181/a_36_216# OR2X1_LOC_181/Y VSS VDD
+ OR2X1_LOC_181/A OR2X1_LOC_181/B OR2X1_LOC
XOR2X1_LOC_170 OR2X1_LOC_170/a_8_216# OR2X1_LOC_170/a_36_216# OR2X1_LOC_170/Y VSS VDD
+ OR2X1_LOC_170/A OR2X1_LOC_168/Y OR2X1_LOC
XOR2X1_LOC_17 OR2X1_LOC_17/a_8_216# OR2X1_LOC_17/a_36_216# OR2X1_LOC_17/Y VSS VDD
+ D_INPUT_7 D_INPUT_6 OR2X1_LOC
XOR2X1_LOC_28 OR2X1_LOC_28/a_8_216# OR2X1_LOC_28/a_36_216# OR2X1_LOC_49/A VSS VDD
+ D_INPUT_1 INPUT_0 OR2X1_LOC
XOR2X1_LOC_39 OR2X1_LOC_39/a_8_216# OR2X1_LOC_39/a_36_216# OR2X1_LOC_39/Y VSS VDD
+ OR2X1_LOC_39/A OR2X1_LOC_36/Y OR2X1_LOC
XAND2X1_LOC_608 AND2X1_LOC_608/a_36_24# OR2X1_LOC_609/A AND2X1_LOC_608/a_8_24# VSS VDD
+ OR2X1_LOC_16/A OR2X1_LOC_74/A AND2X1_LOC
XAND2X1_LOC_619 AND2X1_LOC_619/a_36_24# OR2X1_LOC_622/B AND2X1_LOC_619/a_8_24# VSS VDD
+ AND2X1_LOC_36/Y AND2X1_LOC_619/B AND2X1_LOC
XAND2X1_LOC_416 AND2X1_LOC_416/a_36_24# OR2X1_LOC_462/B AND2X1_LOC_416/a_8_24# VSS VDD
+ OR2X1_LOC_375/A OR2X1_LOC_415/Y AND2X1_LOC
XAND2X1_LOC_438 AND2X1_LOC_438/a_36_24# OR2X1_LOC_544/A AND2X1_LOC_438/a_8_24# VSS VDD
+ OR2X1_LOC_160/B AND2X1_LOC_70/Y AND2X1_LOC
XAND2X1_LOC_405 AND2X1_LOC_405/a_36_24# OR2X1_LOC_406/A AND2X1_LOC_405/a_8_24# VSS VDD
+ OR2X1_LOC_48/B OR2X1_LOC_329/B AND2X1_LOC
XAND2X1_LOC_427 AND2X1_LOC_427/a_36_24# OR2X1_LOC_450/A AND2X1_LOC_427/a_8_24# VSS VDD
+ AND2X1_LOC_70/Y OR2X1_LOC_161/B AND2X1_LOC
XAND2X1_LOC_449 AND2X1_LOC_449/a_36_24# AND2X1_LOC_449/Y AND2X1_LOC_449/a_8_24# VSS VDD
+ OR2X1_LOC_423/Y OR2X1_LOC_424/Y AND2X1_LOC
XOR2X1_LOC_703 OR2X1_LOC_703/a_8_216# OR2X1_LOC_703/a_36_216# OR2X1_LOC_703/Y VSS VDD
+ OR2X1_LOC_703/A OR2X1_LOC_703/B OR2X1_LOC
XOR2X1_LOC_747 OR2X1_LOC_747/a_8_216# OR2X1_LOC_747/a_36_216# OR2X1_LOC_747/Y VSS VDD
+ OR2X1_LOC_52/B OR2X1_LOC_47/Y OR2X1_LOC
XOR2X1_LOC_725 OR2X1_LOC_725/a_8_216# OR2X1_LOC_725/a_36_216# OR2X1_LOC_732/A VSS VDD
+ OR2X1_LOC_725/A OR2X1_LOC_725/B OR2X1_LOC
XOR2X1_LOC_714 OR2X1_LOC_714/a_8_216# OR2X1_LOC_714/a_36_216# OR2X1_LOC_714/Y VSS VDD
+ OR2X1_LOC_714/A OR2X1_LOC_703/Y OR2X1_LOC
XOR2X1_LOC_758 OR2X1_LOC_758/a_8_216# OR2X1_LOC_758/a_36_216# OR2X1_LOC_758/Y VSS VDD
+ AND2X1_LOC_95/Y AND2X1_LOC_40/Y OR2X1_LOC
XOR2X1_LOC_736 OR2X1_LOC_736/a_8_216# OR2X1_LOC_736/a_36_216# OR2X1_LOC_736/Y VSS VDD
+ OR2X1_LOC_736/A OR2X1_LOC_675/Y OR2X1_LOC
XOR2X1_LOC_769 OR2X1_LOC_769/a_8_216# OR2X1_LOC_769/a_36_216# OR2X1_LOC_771/B VSS VDD
+ OR2X1_LOC_769/A OR2X1_LOC_769/B OR2X1_LOC
XAND2X1_LOC_224 AND2X1_LOC_224/a_36_24# OR2X1_LOC_227/B AND2X1_LOC_224/a_8_24# VSS VDD
+ AND2X1_LOC_31/Y OR2X1_LOC_160/A AND2X1_LOC
XAND2X1_LOC_202 AND2X1_LOC_202/a_36_24# AND2X1_LOC_202/Y AND2X1_LOC_202/a_8_24# VSS VDD
+ OR2X1_LOC_67/Y OR2X1_LOC_69/Y AND2X1_LOC
XAND2X1_LOC_268 AND2X1_LOC_268/a_36_24# OR2X1_LOC_269/A AND2X1_LOC_268/a_8_24# VSS VDD
+ AND2X1_LOC_36/Y AND2X1_LOC_92/Y AND2X1_LOC
XAND2X1_LOC_235 AND2X1_LOC_235/a_36_24# OR2X1_LOC_243/B AND2X1_LOC_235/a_8_24# VSS VDD
+ OR2X1_LOC_71/A AND2X1_LOC_86/B AND2X1_LOC
XAND2X1_LOC_279 AND2X1_LOC_279/a_36_24# OR2X1_LOC_284/B AND2X1_LOC_279/a_8_24# VSS VDD
+ AND2X1_LOC_44/Y OR2X1_LOC_161/B AND2X1_LOC
XAND2X1_LOC_257 AND2X1_LOC_257/a_36_24# OR2X1_LOC_259/B AND2X1_LOC_257/a_8_24# VSS VDD
+ AND2X1_LOC_18/Y OR2X1_LOC_161/B AND2X1_LOC
XAND2X1_LOC_246 AND2X1_LOC_246/a_36_24# OR2X1_LOC_342/B AND2X1_LOC_246/a_8_24# VSS VDD
+ OR2X1_LOC_62/B OR2X1_LOC_777/B AND2X1_LOC
XAND2X1_LOC_213 AND2X1_LOC_213/a_36_24# AND2X1_LOC_220/B AND2X1_LOC_213/a_8_24# VSS VDD
+ AND2X1_LOC_209/Y AND2X1_LOC_213/B AND2X1_LOC
XOR2X1_LOC_511 OR2X1_LOC_511/a_8_216# OR2X1_LOC_511/a_36_216# OR2X1_LOC_511/Y VSS VDD
+ OR2X1_LOC_48/B OR2X1_LOC_31/Y OR2X1_LOC
XOR2X1_LOC_533 OR2X1_LOC_533/a_8_216# OR2X1_LOC_533/a_36_216# OR2X1_LOC_533/Y VSS VDD
+ OR2X1_LOC_533/A OR2X1_LOC_95/Y OR2X1_LOC
XOR2X1_LOC_500 OR2X1_LOC_500/a_8_216# OR2X1_LOC_500/a_36_216# OR2X1_LOC_501/A VSS VDD
+ OR2X1_LOC_500/A OR2X1_LOC_844/B OR2X1_LOC
XOR2X1_LOC_522 OR2X1_LOC_522/a_8_216# OR2X1_LOC_522/a_36_216# OR2X1_LOC_522/Y VSS VDD
+ OR2X1_LOC_485/A OR2X1_LOC_22/Y OR2X1_LOC
XOR2X1_LOC_544 OR2X1_LOC_544/a_8_216# OR2X1_LOC_544/a_36_216# OR2X1_LOC_551/B VSS VDD
+ OR2X1_LOC_544/A OR2X1_LOC_544/B OR2X1_LOC
XOR2X1_LOC_588 OR2X1_LOC_588/a_8_216# OR2X1_LOC_588/a_36_216# OR2X1_LOC_588/Y VSS VDD
+ OR2X1_LOC_588/A OR2X1_LOC_696/A OR2X1_LOC
XOR2X1_LOC_599 OR2X1_LOC_599/a_8_216# OR2X1_LOC_599/a_36_216# OR2X1_LOC_599/Y VSS VDD
+ OR2X1_LOC_599/A OR2X1_LOC_36/Y OR2X1_LOC
XAND2X1_LOC_791 AND2X1_LOC_791/a_36_24# AND2X1_LOC_792/B AND2X1_LOC_791/a_8_24# VSS VDD
+ OR2X1_LOC_755/Y OR2X1_LOC_757/Y AND2X1_LOC
XAND2X1_LOC_780 AND2X1_LOC_780/a_36_24# AND2X1_LOC_783/B AND2X1_LOC_780/a_8_24# VSS VDD
+ OR2X1_LOC_743/Y OR2X1_LOC_744/Y AND2X1_LOC
XOR2X1_LOC_555 OR2X1_LOC_555/a_8_216# OR2X1_LOC_555/a_36_216# OR2X1_LOC_562/B VSS VDD
+ OR2X1_LOC_555/A OR2X1_LOC_555/B OR2X1_LOC
XOR2X1_LOC_577 OR2X1_LOC_577/a_8_216# OR2X1_LOC_577/a_36_216# OR2X1_LOC_577/Y VSS VDD
+ OR2X1_LOC_570/Y OR2X1_LOC_577/B OR2X1_LOC
XOR2X1_LOC_566 OR2X1_LOC_566/a_8_216# OR2X1_LOC_566/a_36_216# OR2X1_LOC_566/Y VSS VDD
+ OR2X1_LOC_566/A OR2X1_LOC_170/Y OR2X1_LOC
XOR2X1_LOC_385 OR2X1_LOC_385/a_8_216# OR2X1_LOC_385/a_36_216# OR2X1_LOC_385/Y VSS VDD
+ OR2X1_LOC_600/A OR2X1_LOC_26/Y OR2X1_LOC
XOR2X1_LOC_363 OR2X1_LOC_363/a_8_216# OR2X1_LOC_363/a_36_216# OR2X1_LOC_366/A VSS VDD
+ OR2X1_LOC_363/A OR2X1_LOC_363/B OR2X1_LOC
XOR2X1_LOC_396 OR2X1_LOC_396/a_8_216# OR2X1_LOC_396/a_36_216# OR2X1_LOC_396/Y VSS VDD
+ OR2X1_LOC_36/Y OR2X1_LOC_45/B OR2X1_LOC
XOR2X1_LOC_341 OR2X1_LOC_341/a_8_216# OR2X1_LOC_341/a_36_216# OR2X1_LOC_341/Y VSS VDD
+ OR2X1_LOC_641/B OR2X1_LOC_228/Y OR2X1_LOC
XOR2X1_LOC_374 OR2X1_LOC_374/a_8_216# OR2X1_LOC_374/a_36_216# OR2X1_LOC_374/Y VSS VDD
+ OR2X1_LOC_544/B OR2X1_LOC_325/B OR2X1_LOC
XOR2X1_LOC_352 OR2X1_LOC_352/a_8_216# OR2X1_LOC_352/a_36_216# OR2X1_LOC_357/B VSS VDD
+ OR2X1_LOC_352/A OR2X1_LOC_212/B OR2X1_LOC
XOR2X1_LOC_330 OR2X1_LOC_330/a_8_216# OR2X1_LOC_330/a_36_216# OR2X1_LOC_330/Y VSS VDD
+ AND2X1_LOC_70/Y AND2X1_LOC_51/Y OR2X1_LOC
XOR2X1_LOC_160 OR2X1_LOC_160/a_8_216# OR2X1_LOC_160/a_36_216# OR2X1_LOC_160/Y VSS VDD
+ OR2X1_LOC_160/A OR2X1_LOC_160/B OR2X1_LOC
XOR2X1_LOC_193 OR2X1_LOC_193/a_8_216# OR2X1_LOC_193/a_36_216# OR2X1_LOC_193/Y VSS VDD
+ OR2X1_LOC_193/A AND2X1_LOC_7/Y OR2X1_LOC
XOR2X1_LOC_182 OR2X1_LOC_182/a_8_216# OR2X1_LOC_182/a_36_216# OR2X1_LOC_212/B VSS VDD
+ OR2X1_LOC_181/Y OR2X1_LOC_182/B OR2X1_LOC
XOR2X1_LOC_171 OR2X1_LOC_171/a_8_216# OR2X1_LOC_171/a_36_216# OR2X1_LOC_171/Y VSS VDD
+ OR2X1_LOC_40/Y OR2X1_LOC_45/B OR2X1_LOC
XOR2X1_LOC_18 OR2X1_LOC_18/a_8_216# OR2X1_LOC_18/a_36_216# OR2X1_LOC_18/Y VSS VDD
+ OR2X1_LOC_17/Y OR2X1_LOC_11/Y OR2X1_LOC
XOR2X1_LOC_29 OR2X1_LOC_29/a_8_216# OR2X1_LOC_29/a_36_216# OR2X1_LOC_32/B VSS VDD
+ OR2X1_LOC_80/A OR2X1_LOC_8/Y OR2X1_LOC
XAND2X1_LOC_609 AND2X1_LOC_609/a_36_24# OR2X1_LOC_646/A AND2X1_LOC_609/a_8_24# VSS VDD
+ AND2X1_LOC_59/Y OR2X1_LOC_608/Y AND2X1_LOC
XAND2X1_LOC_406 AND2X1_LOC_406/a_36_24# OR2X1_LOC_475/B AND2X1_LOC_406/a_8_24# VSS VDD
+ AND2X1_LOC_95/Y OR2X1_LOC_405/Y AND2X1_LOC
XAND2X1_LOC_439 AND2X1_LOC_439/a_36_24# AND2X1_LOC_675/A AND2X1_LOC_439/a_8_24# VSS VDD
+ OR2X1_LOC_177/Y OR2X1_LOC_438/Y AND2X1_LOC
XAND2X1_LOC_417 AND2X1_LOC_417/a_36_24# OR2X1_LOC_446/B AND2X1_LOC_417/a_8_24# VSS VDD
+ AND2X1_LOC_47/Y OR2X1_LOC_814/A AND2X1_LOC
XAND2X1_LOC_428 AND2X1_LOC_428/a_36_24# OR2X1_LOC_451/B AND2X1_LOC_428/a_8_24# VSS VDD
+ AND2X1_LOC_31/Y OR2X1_LOC_269/B AND2X1_LOC
XOR2X1_LOC_715 OR2X1_LOC_715/a_8_216# OR2X1_LOC_715/a_36_216# OR2X1_LOC_724/A VSS VDD
+ OR2X1_LOC_715/A OR2X1_LOC_715/B OR2X1_LOC
XOR2X1_LOC_704 OR2X1_LOC_704/a_8_216# OR2X1_LOC_704/a_36_216# OR2X1_LOC_714/A VSS VDD
+ OR2X1_LOC_446/B OR2X1_LOC_317/B OR2X1_LOC
XOR2X1_LOC_726 OR2X1_LOC_726/a_8_216# OR2X1_LOC_726/a_36_216# OR2X1_LOC_731/B VSS VDD
+ OR2X1_LOC_726/A OR2X1_LOC_209/A OR2X1_LOC
XOR2X1_LOC_748 OR2X1_LOC_748/a_8_216# OR2X1_LOC_748/a_36_216# OR2X1_LOC_748/Y VSS VDD
+ OR2X1_LOC_748/A OR2X1_LOC_6/B OR2X1_LOC
XOR2X1_LOC_759 OR2X1_LOC_759/a_8_216# OR2X1_LOC_759/a_36_216# OR2X1_LOC_759/Y VSS VDD
+ OR2X1_LOC_759/A OR2X1_LOC_428/A OR2X1_LOC
XOR2X1_LOC_737 OR2X1_LOC_737/a_8_216# OR2X1_LOC_737/a_36_216# OR2X1_LOC_741/A VSS VDD
+ OR2X1_LOC_737/A OR2X1_LOC_733/Y OR2X1_LOC
XAND2X1_LOC_203 AND2X1_LOC_203/a_36_24# AND2X1_LOC_203/Y AND2X1_LOC_203/a_8_24# VSS VDD
+ OR2X1_LOC_72/Y AND2X1_LOC_76/Y AND2X1_LOC
XAND2X1_LOC_247 AND2X1_LOC_247/a_36_24# OR2X1_LOC_248/A AND2X1_LOC_247/a_8_24# VSS VDD
+ OR2X1_LOC_7/A OR2X1_LOC_13/B AND2X1_LOC
XAND2X1_LOC_258 AND2X1_LOC_258/a_36_24# OR2X1_LOC_259/A AND2X1_LOC_258/a_8_24# VSS VDD
+ OR2X1_LOC_78/A OR2X1_LOC_375/A AND2X1_LOC
XAND2X1_LOC_225 AND2X1_LOC_225/a_36_24# OR2X1_LOC_814/A AND2X1_LOC_225/a_8_24# VSS VDD
+ D_INPUT_1 OR2X1_LOC_68/B AND2X1_LOC
XAND2X1_LOC_236 AND2X1_LOC_236/a_36_24# OR2X1_LOC_269/B AND2X1_LOC_236/a_8_24# VSS VDD
+ OR2X1_LOC_68/B OR2X1_LOC_80/A AND2X1_LOC
XAND2X1_LOC_269 AND2X1_LOC_269/a_36_24# OR2X1_LOC_271/B AND2X1_LOC_269/a_8_24# VSS VDD
+ OR2X1_LOC_428/A OR2X1_LOC_268/Y AND2X1_LOC
XAND2X1_LOC_214 AND2X1_LOC_214/a_36_24# AND2X1_LOC_219/A AND2X1_LOC_214/a_8_24# VSS VDD
+ AND2X1_LOC_214/A AND2X1_LOC_208/Y AND2X1_LOC
XOR2X1_LOC_512 OR2X1_LOC_512/a_8_216# OR2X1_LOC_512/a_36_216# OR2X1_LOC_512/Y VSS VDD
+ OR2X1_LOC_512/A D_INPUT_0 OR2X1_LOC
XOR2X1_LOC_534 OR2X1_LOC_534/a_8_216# OR2X1_LOC_534/a_36_216# OR2X1_LOC_534/Y VSS VDD
+ OR2X1_LOC_59/Y OR2X1_LOC_43/A OR2X1_LOC
XOR2X1_LOC_501 OR2X1_LOC_501/a_8_216# OR2X1_LOC_501/a_36_216# OR2X1_LOC_735/B VSS VDD
+ OR2X1_LOC_501/A OR2X1_LOC_501/B OR2X1_LOC
XOR2X1_LOC_523 OR2X1_LOC_523/a_8_216# OR2X1_LOC_523/a_36_216# OR2X1_LOC_523/Y VSS VDD
+ OR2X1_LOC_523/A OR2X1_LOC_523/B OR2X1_LOC
XOR2X1_LOC_556 OR2X1_LOC_556/a_8_216# OR2X1_LOC_556/a_36_216# OR2X1_LOC_562/A VSS VDD
+ OR2X1_LOC_486/Y OR2X1_LOC_631/B OR2X1_LOC
XOR2X1_LOC_578 OR2X1_LOC_578/a_8_216# OR2X1_LOC_578/a_36_216# OR2X1_LOC_580/B VSS VDD
+ OR2X1_LOC_577/Y OR2X1_LOC_578/B OR2X1_LOC
XOR2X1_LOC_545 OR2X1_LOC_545/a_8_216# OR2X1_LOC_545/a_36_216# OR2X1_LOC_551/A VSS VDD
+ OR2X1_LOC_545/A OR2X1_LOC_545/B OR2X1_LOC
XOR2X1_LOC_567 OR2X1_LOC_567/a_8_216# OR2X1_LOC_567/a_36_216# OR2X1_LOC_568/A VSS VDD
+ OR2X1_LOC_539/Y OR2X1_LOC_854/A OR2X1_LOC
XOR2X1_LOC_589 OR2X1_LOC_589/a_8_216# OR2X1_LOC_589/a_36_216# OR2X1_LOC_589/Y VSS VDD
+ OR2X1_LOC_589/A OR2X1_LOC_22/Y OR2X1_LOC
XAND2X1_LOC_792 AND2X1_LOC_792/a_36_24# AND2X1_LOC_792/Y AND2X1_LOC_792/a_8_24# VSS VDD
+ OR2X1_LOC_759/Y AND2X1_LOC_792/B AND2X1_LOC
XAND2X1_LOC_770 AND2X1_LOC_770/a_36_24# AND2X1_LOC_771/B AND2X1_LOC_770/a_8_24# VSS VDD
+ OR2X1_LOC_765/Y OR2X1_LOC_766/Y AND2X1_LOC
XAND2X1_LOC_781 AND2X1_LOC_781/a_36_24# AND2X1_LOC_781/Y AND2X1_LOC_781/a_8_24# VSS VDD
+ OR2X1_LOC_745/Y OR2X1_LOC_746/Y AND2X1_LOC
XOR2X1_LOC_386 OR2X1_LOC_386/a_8_216# OR2X1_LOC_386/a_36_216# OR2X1_LOC_387/A VSS VDD
+ OR2X1_LOC_17/Y INPUT_4 OR2X1_LOC
XOR2X1_LOC_375 OR2X1_LOC_375/a_8_216# OR2X1_LOC_375/a_36_216# OR2X1_LOC_375/Y VSS VDD
+ OR2X1_LOC_375/A AND2X1_LOC_31/Y OR2X1_LOC
XOR2X1_LOC_331 OR2X1_LOC_331/a_8_216# OR2X1_LOC_331/a_36_216# OR2X1_LOC_331/Y VSS VDD
+ OR2X1_LOC_331/A OR2X1_LOC_680/A OR2X1_LOC
XOR2X1_LOC_342 OR2X1_LOC_342/a_8_216# OR2X1_LOC_342/a_36_216# OR2X1_LOC_349/B VSS VDD
+ OR2X1_LOC_342/A OR2X1_LOC_342/B OR2X1_LOC
XOR2X1_LOC_397 OR2X1_LOC_397/a_8_216# OR2X1_LOC_397/a_36_216# OR2X1_LOC_397/Y VSS VDD
+ OR2X1_LOC_83/A OR2X1_LOC_3/Y OR2X1_LOC
XOR2X1_LOC_364 OR2X1_LOC_364/a_8_216# OR2X1_LOC_364/a_36_216# OR2X1_LOC_364/Y VSS VDD
+ OR2X1_LOC_364/A OR2X1_LOC_364/B OR2X1_LOC
XOR2X1_LOC_353 OR2X1_LOC_353/a_8_216# OR2X1_LOC_353/a_36_216# OR2X1_LOC_357/A VSS VDD
+ OR2X1_LOC_308/Y OR2X1_LOC_566/A OR2X1_LOC
XOR2X1_LOC_320 OR2X1_LOC_320/a_8_216# OR2X1_LOC_320/a_36_216# OR2X1_LOC_320/Y VSS VDD
+ OR2X1_LOC_91/A OR2X1_LOC_36/Y OR2X1_LOC
XOR2X1_LOC_161 OR2X1_LOC_161/a_8_216# OR2X1_LOC_161/a_36_216# OR2X1_LOC_162/A VSS VDD
+ OR2X1_LOC_161/A OR2X1_LOC_161/B OR2X1_LOC
XOR2X1_LOC_194 OR2X1_LOC_194/a_8_216# OR2X1_LOC_194/a_36_216# OR2X1_LOC_194/Y VSS VDD
+ AND2X1_LOC_39/Y OR2X1_LOC_194/B OR2X1_LOC
XOR2X1_LOC_172 OR2X1_LOC_172/a_8_216# OR2X1_LOC_172/a_36_216# OR2X1_LOC_172/Y VSS VDD
+ OR2X1_LOC_485/A OR2X1_LOC_70/Y OR2X1_LOC
XOR2X1_LOC_150 OR2X1_LOC_150/a_8_216# OR2X1_LOC_150/a_36_216# OR2X1_LOC_437/A VSS VDD
+ OR2X1_LOC_71/A OR2X1_LOC_85/A OR2X1_LOC
XOR2X1_LOC_183 OR2X1_LOC_183/a_8_216# OR2X1_LOC_183/a_36_216# OR2X1_LOC_183/Y VSS VDD
+ OR2X1_LOC_40/Y OR2X1_LOC_7/A OR2X1_LOC
XOR2X1_LOC_19 OR2X1_LOC_19/a_8_216# OR2X1_LOC_19/a_36_216# OR2X1_LOC_20/A VSS VDD
+ OR2X1_LOC_6/A OR2X1_LOC_19/B OR2X1_LOC
XAND2X1_LOC_407 AND2X1_LOC_407/a_36_24# OR2X1_LOC_409/B AND2X1_LOC_407/a_8_24# VSS VDD
+ OR2X1_LOC_56/A OR2X1_LOC_743/A AND2X1_LOC
XAND2X1_LOC_418 AND2X1_LOC_418/a_36_24# OR2X1_LOC_446/A AND2X1_LOC_418/a_8_24# VSS VDD
+ OR2X1_LOC_78/B AND2X1_LOC_51/Y AND2X1_LOC
XAND2X1_LOC_429 AND2X1_LOC_429/a_36_24# AND2X1_LOC_430/B AND2X1_LOC_429/a_8_24# VSS VDD
+ D_INPUT_7 AND2X1_LOC_11/Y AND2X1_LOC
XOR2X1_LOC_705 OR2X1_LOC_705/a_8_216# OR2X1_LOC_705/a_36_216# OR2X1_LOC_705/Y VSS VDD
+ OR2X1_LOC_546/A OR2X1_LOC_705/B OR2X1_LOC
XOR2X1_LOC_727 OR2X1_LOC_727/a_8_216# OR2X1_LOC_727/a_36_216# OR2X1_LOC_731/A VSS VDD
+ OR2X1_LOC_469/B OR2X1_LOC_308/Y OR2X1_LOC
XOR2X1_LOC_738 OR2X1_LOC_738/a_8_216# OR2X1_LOC_738/a_36_216# OR2X1_LOC_740/B VSS VDD
+ OR2X1_LOC_738/A OR2X1_LOC_738/B OR2X1_LOC
XOR2X1_LOC_749 OR2X1_LOC_749/a_8_216# OR2X1_LOC_749/a_36_216# OR2X1_LOC_749/Y VSS VDD
+ OR2X1_LOC_8/Y INPUT_0 OR2X1_LOC
XOR2X1_LOC_716 OR2X1_LOC_716/a_8_216# OR2X1_LOC_716/a_36_216# OR2X1_LOC_723/B VSS VDD
+ OR2X1_LOC_303/B OR2X1_LOC_228/Y OR2X1_LOC
XAND2X1_LOC_226 AND2X1_LOC_226/a_36_24# OR2X1_LOC_227/A AND2X1_LOC_226/a_8_24# VSS VDD
+ AND2X1_LOC_18/Y OR2X1_LOC_814/A AND2X1_LOC
XAND2X1_LOC_237 AND2X1_LOC_237/a_36_24# OR2X1_LOC_241/B AND2X1_LOC_237/a_8_24# VSS VDD
+ OR2X1_LOC_66/A OR2X1_LOC_269/B AND2X1_LOC
XAND2X1_LOC_215 AND2X1_LOC_215/a_36_24# AND2X1_LOC_215/Y AND2X1_LOC_215/a_8_24# VSS VDD
+ AND2X1_LOC_215/A AND2X1_LOC_206/Y AND2X1_LOC
XAND2X1_LOC_204 AND2X1_LOC_204/a_36_24# AND2X1_LOC_204/Y AND2X1_LOC_204/a_8_24# VSS VDD
+ OR2X1_LOC_79/Y AND2X1_LOC_84/Y AND2X1_LOC
XAND2X1_LOC_248 AND2X1_LOC_248/a_36_24# OR2X1_LOC_342/A AND2X1_LOC_248/a_8_24# VSS VDD
+ AND2X1_LOC_47/Y OR2X1_LOC_247/Y AND2X1_LOC
XAND2X1_LOC_259 AND2X1_LOC_259/a_36_24# AND2X1_LOC_259/Y AND2X1_LOC_259/a_8_24# VSS VDD
+ OR2X1_LOC_257/Y OR2X1_LOC_258/Y AND2X1_LOC
XOR2X1_LOC_513 OR2X1_LOC_513/a_8_216# OR2X1_LOC_513/a_36_216# OR2X1_LOC_513/Y VSS VDD
+ OR2X1_LOC_512/Y OR2X1_LOC_779/B OR2X1_LOC
XOR2X1_LOC_546 OR2X1_LOC_546/a_8_216# OR2X1_LOC_546/a_36_216# OR2X1_LOC_550/B VSS VDD
+ OR2X1_LOC_546/A OR2X1_LOC_546/B OR2X1_LOC
XAND2X1_LOC_793 AND2X1_LOC_793/a_36_24# AND2X1_LOC_793/Y AND2X1_LOC_793/a_8_24# VSS VDD
+ AND2X1_LOC_789/Y AND2X1_LOC_793/B AND2X1_LOC
XAND2X1_LOC_760 AND2X1_LOC_760/a_36_24# OR2X1_LOC_800/A AND2X1_LOC_760/a_8_24# VSS VDD
+ AND2X1_LOC_64/Y OR2X1_LOC_405/A AND2X1_LOC
XAND2X1_LOC_771 AND2X1_LOC_771/a_36_24# AND2X1_LOC_774/A AND2X1_LOC_771/a_8_24# VSS VDD
+ AND2X1_LOC_769/Y AND2X1_LOC_771/B AND2X1_LOC
XAND2X1_LOC_782 AND2X1_LOC_782/a_36_24# AND2X1_LOC_797/B AND2X1_LOC_782/a_8_24# VSS VDD
+ OR2X1_LOC_747/Y AND2X1_LOC_781/Y AND2X1_LOC
XOR2X1_LOC_557 OR2X1_LOC_557/a_8_216# OR2X1_LOC_557/a_36_216# OR2X1_LOC_561/B VSS VDD
+ OR2X1_LOC_557/A OR2X1_LOC_772/B OR2X1_LOC
XOR2X1_LOC_579 OR2X1_LOC_579/a_8_216# OR2X1_LOC_579/a_36_216# OR2X1_LOC_580/A VSS VDD
+ OR2X1_LOC_579/A OR2X1_LOC_579/B OR2X1_LOC
XOR2X1_LOC_502 OR2X1_LOC_502/a_8_216# OR2X1_LOC_502/a_36_216# OR2X1_LOC_502/Y VSS VDD
+ OR2X1_LOC_502/A OR2X1_LOC_78/A OR2X1_LOC
XOR2X1_LOC_524 OR2X1_LOC_524/a_8_216# OR2X1_LOC_524/a_36_216# OR2X1_LOC_524/Y VSS VDD
+ OR2X1_LOC_427/A OR2X1_LOC_47/Y OR2X1_LOC
XOR2X1_LOC_568 OR2X1_LOC_568/a_8_216# OR2X1_LOC_568/a_36_216# OR2X1_LOC_578/B VSS VDD
+ OR2X1_LOC_568/A OR2X1_LOC_566/Y OR2X1_LOC
XOR2X1_LOC_535 OR2X1_LOC_535/a_8_216# OR2X1_LOC_535/a_36_216# OR2X1_LOC_854/A VSS VDD
+ OR2X1_LOC_535/A OR2X1_LOC_788/B OR2X1_LOC
XOR2X1_LOC_310 OR2X1_LOC_310/a_8_216# OR2X1_LOC_310/a_36_216# OR2X1_LOC_310/Y VSS VDD
+ OR2X1_LOC_40/Y OR2X1_LOC_6/A OR2X1_LOC
XOR2X1_LOC_387 OR2X1_LOC_387/a_8_216# OR2X1_LOC_387/a_36_216# OR2X1_LOC_387/Y VSS VDD
+ OR2X1_LOC_387/A OR2X1_LOC_92/Y OR2X1_LOC
XOR2X1_LOC_376 OR2X1_LOC_376/a_8_216# OR2X1_LOC_376/a_36_216# OR2X1_LOC_376/Y VSS VDD
+ OR2X1_LOC_376/A OR2X1_LOC_696/A OR2X1_LOC
XAND2X1_LOC_590 AND2X1_LOC_590/a_36_24# OR2X1_LOC_591/A AND2X1_LOC_590/a_8_24# VSS VDD
+ OR2X1_LOC_39/A OR2X1_LOC_485/A AND2X1_LOC
XOR2X1_LOC_343 OR2X1_LOC_343/a_8_216# OR2X1_LOC_343/a_36_216# OR2X1_LOC_349/A VSS VDD
+ OR2X1_LOC_843/B OR2X1_LOC_343/B OR2X1_LOC
XOR2X1_LOC_398 OR2X1_LOC_398/a_8_216# OR2X1_LOC_398/a_36_216# OR2X1_LOC_398/Y VSS VDD
+ OR2X1_LOC_598/A OR2X1_LOC_78/B OR2X1_LOC
XOR2X1_LOC_365 OR2X1_LOC_365/a_8_216# OR2X1_LOC_365/a_36_216# OR2X1_LOC_367/B VSS VDD
+ OR2X1_LOC_364/Y OR2X1_LOC_365/B OR2X1_LOC
XOR2X1_LOC_332 OR2X1_LOC_332/a_8_216# OR2X1_LOC_332/a_36_216# OR2X1_LOC_339/A VSS VDD
+ OR2X1_LOC_702/A OR2X1_LOC_112/A OR2X1_LOC
XOR2X1_LOC_354 OR2X1_LOC_354/a_8_216# OR2X1_LOC_354/a_36_216# OR2X1_LOC_356/B VSS VDD
+ OR2X1_LOC_354/A OR2X1_LOC_319/Y OR2X1_LOC
XOR2X1_LOC_321 OR2X1_LOC_321/a_8_216# OR2X1_LOC_321/a_36_216# OR2X1_LOC_321/Y VSS VDD
+ OR2X1_LOC_64/Y OR2X1_LOC_13/B OR2X1_LOC
XOR2X1_LOC_162 OR2X1_LOC_162/a_8_216# OR2X1_LOC_162/a_36_216# OR2X1_LOC_162/Y VSS VDD
+ OR2X1_LOC_162/A OR2X1_LOC_160/Y OR2X1_LOC
XOR2X1_LOC_140 OR2X1_LOC_140/a_8_216# OR2X1_LOC_140/a_36_216# OR2X1_LOC_140/Y VSS VDD
+ OR2X1_LOC_140/A OR2X1_LOC_140/B OR2X1_LOC
XOR2X1_LOC_151 OR2X1_LOC_151/a_8_216# OR2X1_LOC_151/a_36_216# OR2X1_LOC_151/Y VSS VDD
+ OR2X1_LOC_151/A AND2X1_LOC_56/B OR2X1_LOC
XOR2X1_LOC_195 OR2X1_LOC_195/a_8_216# OR2X1_LOC_195/a_36_216# OR2X1_LOC_199/B VSS VDD
+ OR2X1_LOC_195/A AND2X1_LOC_41/Y OR2X1_LOC
XOR2X1_LOC_184 OR2X1_LOC_184/a_8_216# OR2X1_LOC_184/a_36_216# OR2X1_LOC_184/Y VSS VDD
+ OR2X1_LOC_95/Y OR2X1_LOC_71/Y OR2X1_LOC
XOR2X1_LOC_173 OR2X1_LOC_173/a_8_216# OR2X1_LOC_173/a_36_216# OR2X1_LOC_173/Y VSS VDD
+ OR2X1_LOC_437/A OR2X1_LOC_70/Y OR2X1_LOC
XAND2X1_LOC_419 AND2X1_LOC_419/a_36_24# OR2X1_LOC_506/A AND2X1_LOC_419/a_8_24# VSS VDD
+ AND2X1_LOC_36/Y AND2X1_LOC_43/B AND2X1_LOC
XAND2X1_LOC_408 AND2X1_LOC_408/a_36_24# AND2X1_LOC_409/B AND2X1_LOC_408/a_8_24# VSS VDD
+ D_INPUT_6 AND2X1_LOC_21/Y AND2X1_LOC
XOR2X1_LOC_706 OR2X1_LOC_706/a_8_216# OR2X1_LOC_706/a_36_216# OR2X1_LOC_713/A VSS VDD
+ OR2X1_LOC_706/A OR2X1_LOC_706/B OR2X1_LOC
XOR2X1_LOC_717 OR2X1_LOC_717/a_8_216# OR2X1_LOC_717/a_36_216# OR2X1_LOC_723/A VSS VDD
+ OR2X1_LOC_493/Y OR2X1_LOC_374/Y OR2X1_LOC
XOR2X1_LOC_739 OR2X1_LOC_739/a_8_216# OR2X1_LOC_739/a_36_216# OR2X1_LOC_739/Y VSS VDD
+ OR2X1_LOC_739/A OR2X1_LOC_739/B OR2X1_LOC
XOR2X1_LOC_728 OR2X1_LOC_728/a_8_216# OR2X1_LOC_728/a_36_216# OR2X1_LOC_730/B VSS VDD
+ OR2X1_LOC_728/A OR2X1_LOC_728/B OR2X1_LOC
XAND2X1_LOC_238 AND2X1_LOC_238/a_36_24# OR2X1_LOC_776/A AND2X1_LOC_238/a_8_24# VSS VDD
+ OR2X1_LOC_160/B AND2X1_LOC_51/Y AND2X1_LOC
XAND2X1_LOC_227 AND2X1_LOC_227/a_36_24# AND2X1_LOC_227/Y AND2X1_LOC_227/a_8_24# VSS VDD
+ OR2X1_LOC_224/Y OR2X1_LOC_226/Y AND2X1_LOC
XAND2X1_LOC_249 AND2X1_LOC_249/a_36_24# OR2X1_LOC_595/A AND2X1_LOC_249/a_8_24# VSS VDD
+ OR2X1_LOC_45/B OR2X1_LOC_39/A AND2X1_LOC
XAND2X1_LOC_205 AND2X1_LOC_205/a_36_24# AND2X1_LOC_215/A AND2X1_LOC_205/a_8_24# VSS VDD
+ AND2X1_LOC_203/Y AND2X1_LOC_204/Y AND2X1_LOC
XAND2X1_LOC_216 AND2X1_LOC_216/a_36_24# AND2X1_LOC_216/Y AND2X1_LOC_216/a_8_24# VSS VDD
+ AND2X1_LOC_216/A AND2X1_LOC_116/Y AND2X1_LOC
XOR2X1_LOC_536 OR2X1_LOC_536/a_8_216# OR2X1_LOC_536/a_36_216# OR2X1_LOC_536/Y VSS VDD
+ OR2X1_LOC_485/A OR2X1_LOC_12/Y OR2X1_LOC
XOR2X1_LOC_525 OR2X1_LOC_525/a_8_216# OR2X1_LOC_525/a_36_216# OR2X1_LOC_525/Y VSS VDD
+ OR2X1_LOC_51/Y OR2X1_LOC_13/B OR2X1_LOC
XOR2X1_LOC_514 OR2X1_LOC_514/a_8_216# OR2X1_LOC_514/a_36_216# OR2X1_LOC_515/A VSS VDD
+ OR2X1_LOC_138/A INPUT_0 OR2X1_LOC
XAND2X1_LOC_772 AND2X1_LOC_772/a_36_24# AND2X1_LOC_772/Y AND2X1_LOC_772/a_8_24# VSS VDD
+ AND2X1_LOC_489/Y AND2X1_LOC_772/B AND2X1_LOC
XAND2X1_LOC_750 AND2X1_LOC_750/a_36_24# OR2X1_LOC_751/A AND2X1_LOC_750/a_8_24# VSS VDD
+ OR2X1_LOC_604/A OR2X1_LOC_749/Y AND2X1_LOC
XAND2X1_LOC_794 AND2X1_LOC_794/a_36_24# AND2X1_LOC_804/A AND2X1_LOC_794/a_8_24# VSS VDD
+ AND2X1_LOC_794/A AND2X1_LOC_794/B AND2X1_LOC
XAND2X1_LOC_761 AND2X1_LOC_761/a_36_24# OR2X1_LOC_801/B AND2X1_LOC_761/a_8_24# VSS VDD
+ D_INPUT_0 OR2X1_LOC_644/A AND2X1_LOC
XAND2X1_LOC_783 AND2X1_LOC_783/a_36_24# AND2X1_LOC_796/A AND2X1_LOC_783/a_8_24# VSS VDD
+ AND2X1_LOC_779/Y AND2X1_LOC_783/B AND2X1_LOC
XOR2X1_LOC_558 OR2X1_LOC_558/a_8_216# OR2X1_LOC_558/a_36_216# OR2X1_LOC_561/A VSS VDD
+ OR2X1_LOC_558/A OR2X1_LOC_493/Y OR2X1_LOC
XOR2X1_LOC_569 OR2X1_LOC_569/a_8_216# OR2X1_LOC_569/a_36_216# OR2X1_LOC_577/B VSS VDD
+ OR2X1_LOC_569/A OR2X1_LOC_569/B OR2X1_LOC
XOR2X1_LOC_503 OR2X1_LOC_503/a_8_216# OR2X1_LOC_503/a_36_216# OR2X1_LOC_503/Y VSS VDD
+ OR2X1_LOC_503/A OR2X1_LOC_64/Y OR2X1_LOC
XOR2X1_LOC_547 OR2X1_LOC_547/a_8_216# OR2X1_LOC_547/a_36_216# OR2X1_LOC_550/A VSS VDD
+ OR2X1_LOC_620/B OR2X1_LOC_547/B OR2X1_LOC
XOR2X1_LOC_311 OR2X1_LOC_311/a_8_216# OR2X1_LOC_311/a_36_216# OR2X1_LOC_311/Y VSS VDD
+ OR2X1_LOC_485/A OR2X1_LOC_26/Y OR2X1_LOC
XOR2X1_LOC_344 OR2X1_LOC_344/a_8_216# OR2X1_LOC_344/a_36_216# OR2X1_LOC_348/B VSS VDD
+ OR2X1_LOC_344/A OR2X1_LOC_456/A OR2X1_LOC
XOR2X1_LOC_300 OR2X1_LOC_300/a_8_216# OR2X1_LOC_300/a_36_216# OR2X1_LOC_300/Y VSS VDD
+ OR2X1_LOC_426/B OR2X1_LOC_59/Y OR2X1_LOC
XOR2X1_LOC_333 OR2X1_LOC_333/a_8_216# OR2X1_LOC_333/a_36_216# OR2X1_LOC_338/B VSS VDD
+ OR2X1_LOC_333/A OR2X1_LOC_333/B OR2X1_LOC
XOR2X1_LOC_322 OR2X1_LOC_322/a_8_216# OR2X1_LOC_322/a_36_216# OR2X1_LOC_322/Y VSS VDD
+ OR2X1_LOC_696/A OR2X1_LOC_44/Y OR2X1_LOC
XOR2X1_LOC_377 OR2X1_LOC_377/a_8_216# OR2X1_LOC_377/a_36_216# OR2X1_LOC_378/A VSS VDD
+ OR2X1_LOC_377/A OR2X1_LOC_3/Y OR2X1_LOC
XAND2X1_LOC_591 AND2X1_LOC_591/a_36_24# OR2X1_LOC_593/B AND2X1_LOC_591/a_8_24# VSS VDD
+ AND2X1_LOC_64/Y OR2X1_LOC_590/Y AND2X1_LOC
XAND2X1_LOC_580 AND2X1_LOC_580/a_36_24# GATE_579 AND2X1_LOC_580/a_8_24# VSS VDD
+ AND2X1_LOC_580/A AND2X1_LOC_580/B AND2X1_LOC
XOR2X1_LOC_366 OR2X1_LOC_366/a_8_216# OR2X1_LOC_366/a_36_216# OR2X1_LOC_366/Y VSS VDD
+ OR2X1_LOC_366/A OR2X1_LOC_366/B OR2X1_LOC
XOR2X1_LOC_399 OR2X1_LOC_399/a_8_216# OR2X1_LOC_399/a_36_216# OR2X1_LOC_399/Y VSS VDD
+ OR2X1_LOC_399/A OR2X1_LOC_44/Y OR2X1_LOC
XOR2X1_LOC_388 OR2X1_LOC_388/a_8_216# OR2X1_LOC_388/a_36_216# OR2X1_LOC_390/B VSS VDD
+ OR2X1_LOC_180/B OR2X1_LOC_703/B OR2X1_LOC
XOR2X1_LOC_355 OR2X1_LOC_355/a_8_216# OR2X1_LOC_355/a_36_216# OR2X1_LOC_356/A VSS VDD
+ OR2X1_LOC_355/A OR2X1_LOC_355/B OR2X1_LOC
XOR2X1_LOC_163 OR2X1_LOC_163/a_8_216# OR2X1_LOC_163/a_36_216# OR2X1_LOC_163/Y VSS VDD
+ OR2X1_LOC_163/A OR2X1_LOC_51/Y OR2X1_LOC
XOR2X1_LOC_152 OR2X1_LOC_152/a_8_216# OR2X1_LOC_152/a_36_216# OR2X1_LOC_152/Y VSS VDD
+ OR2X1_LOC_152/A OR2X1_LOC_47/Y OR2X1_LOC
XOR2X1_LOC_141 OR2X1_LOC_141/a_8_216# OR2X1_LOC_141/a_36_216# OR2X1_LOC_217/A VSS VDD
+ OR2X1_LOC_140/Y OR2X1_LOC_141/B OR2X1_LOC
XOR2X1_LOC_130 OR2X1_LOC_130/a_8_216# OR2X1_LOC_130/a_36_216# OR2X1_LOC_130/Y VSS VDD
+ OR2X1_LOC_130/A AND2X1_LOC_7/B OR2X1_LOC
XOR2X1_LOC_174 OR2X1_LOC_174/a_8_216# OR2X1_LOC_174/a_36_216# OR2X1_LOC_174/Y VSS VDD
+ OR2X1_LOC_174/A OR2X1_LOC_333/B OR2X1_LOC
XOR2X1_LOC_185 OR2X1_LOC_185/a_8_216# OR2X1_LOC_185/a_36_216# OR2X1_LOC_185/Y VSS VDD
+ OR2X1_LOC_185/A AND2X1_LOC_56/B OR2X1_LOC
XOR2X1_LOC_196 OR2X1_LOC_196/a_8_216# OR2X1_LOC_196/a_36_216# OR2X1_LOC_196/Y VSS VDD
+ AND2X1_LOC_48/Y OR2X1_LOC_196/B OR2X1_LOC
XAND2X1_LOC_409 AND2X1_LOC_409/a_36_24# OR2X1_LOC_460/A AND2X1_LOC_409/a_8_24# VSS VDD
+ OR2X1_LOC_828/B AND2X1_LOC_409/B AND2X1_LOC
XOR2X1_LOC_707 OR2X1_LOC_707/a_8_216# OR2X1_LOC_707/a_36_216# OR2X1_LOC_712/B VSS VDD
+ OR2X1_LOC_707/A OR2X1_LOC_707/B OR2X1_LOC
XOR2X1_LOC_718 OR2X1_LOC_718/a_8_216# OR2X1_LOC_718/a_36_216# OR2X1_LOC_722/B VSS VDD
+ OR2X1_LOC_605/Y OR2X1_LOC_593/B OR2X1_LOC
XOR2X1_LOC_729 OR2X1_LOC_729/a_8_216# OR2X1_LOC_729/a_36_216# OR2X1_LOC_730/A VSS VDD
+ OR2X1_LOC_691/Y OR2X1_LOC_687/Y OR2X1_LOC
XAND2X1_LOC_217 AND2X1_LOC_217/a_36_24# AND2X1_LOC_217/Y AND2X1_LOC_217/a_8_24# VSS VDD
+ AND2X1_LOC_572/A AND2X1_LOC_657/A AND2X1_LOC
XAND2X1_LOC_239 AND2X1_LOC_239/a_36_24# OR2X1_LOC_506/B AND2X1_LOC_239/a_8_24# VSS VDD
+ AND2X1_LOC_51/Y OR2X1_LOC_532/B AND2X1_LOC
XAND2X1_LOC_206 AND2X1_LOC_206/a_36_24# AND2X1_LOC_206/Y AND2X1_LOC_206/a_8_24# VSS VDD
+ AND2X1_LOC_201/Y AND2X1_LOC_202/Y AND2X1_LOC
XAND2X1_LOC_228 AND2X1_LOC_228/a_36_24# AND2X1_LOC_228/Y AND2X1_LOC_228/a_8_24# VSS VDD
+ OR2X1_LOC_7/Y OR2X1_LOC_52/Y AND2X1_LOC
XOR2X1_LOC_526 OR2X1_LOC_526/a_8_216# OR2X1_LOC_526/a_36_216# OR2X1_LOC_526/Y VSS VDD
+ OR2X1_LOC_604/A OR2X1_LOC_31/Y OR2X1_LOC
XOR2X1_LOC_515 OR2X1_LOC_515/a_8_216# OR2X1_LOC_515/a_36_216# OR2X1_LOC_515/Y VSS VDD
+ OR2X1_LOC_515/A OR2X1_LOC_446/B OR2X1_LOC
XOR2X1_LOC_504 OR2X1_LOC_504/a_8_216# OR2X1_LOC_504/a_36_216# OR2X1_LOC_504/Y VSS VDD
+ OR2X1_LOC_158/A OR2X1_LOC_13/B OR2X1_LOC
XAND2X1_LOC_773 AND2X1_LOC_773/a_36_24# AND2X1_LOC_773/Y AND2X1_LOC_773/a_8_24# VSS VDD
+ OR2X1_LOC_767/Y AND2X1_LOC_772/Y AND2X1_LOC
XAND2X1_LOC_795 AND2X1_LOC_795/a_36_24# AND2X1_LOC_795/Y AND2X1_LOC_795/a_8_24# VSS VDD
+ AND2X1_LOC_785/Y AND2X1_LOC_786/Y AND2X1_LOC
XAND2X1_LOC_784 AND2X1_LOC_784/a_36_24# AND2X1_LOC_784/Y AND2X1_LOC_784/a_8_24# VSS VDD
+ AND2X1_LOC_784/A AND2X1_LOC_778/Y AND2X1_LOC
XAND2X1_LOC_751 AND2X1_LOC_751/a_36_24# OR2X1_LOC_789/A AND2X1_LOC_751/a_8_24# VSS VDD
+ AND2X1_LOC_3/Y OR2X1_LOC_750/Y AND2X1_LOC
XAND2X1_LOC_740 AND2X1_LOC_740/a_36_24# AND2X1_LOC_742/A AND2X1_LOC_740/a_8_24# VSS VDD
+ AND2X1_LOC_738/Y AND2X1_LOC_740/B AND2X1_LOC
XAND2X1_LOC_762 AND2X1_LOC_762/a_36_24# AND2X1_LOC_763/B AND2X1_LOC_762/a_8_24# VSS VDD
+ INPUT_6 AND2X1_LOC_11/Y AND2X1_LOC
XOR2X1_LOC_548 OR2X1_LOC_548/a_8_216# OR2X1_LOC_548/a_36_216# OR2X1_LOC_549/A VSS VDD
+ OR2X1_LOC_548/A OR2X1_LOC_548/B OR2X1_LOC
XOR2X1_LOC_559 OR2X1_LOC_559/a_8_216# OR2X1_LOC_559/a_36_216# OR2X1_LOC_560/A VSS VDD
+ OR2X1_LOC_520/Y OR2X1_LOC_559/B OR2X1_LOC
XOR2X1_LOC_537 OR2X1_LOC_537/a_8_216# OR2X1_LOC_537/a_36_216# OR2X1_LOC_539/B VSS VDD
+ OR2X1_LOC_537/A OR2X1_LOC_389/B OR2X1_LOC
XOR2X1_LOC_312 OR2X1_LOC_312/a_8_216# OR2X1_LOC_312/a_36_216# OR2X1_LOC_312/Y VSS VDD
+ OR2X1_LOC_64/Y OR2X1_LOC_56/A OR2X1_LOC
XOR2X1_LOC_378 OR2X1_LOC_378/a_8_216# OR2X1_LOC_378/a_36_216# OR2X1_LOC_378/Y VSS VDD
+ OR2X1_LOC_378/A AND2X1_LOC_43/B OR2X1_LOC
XOR2X1_LOC_345 OR2X1_LOC_345/a_8_216# OR2X1_LOC_345/a_36_216# OR2X1_LOC_345/Y VSS VDD
+ OR2X1_LOC_345/A OR2X1_LOC_555/B OR2X1_LOC
XOR2X1_LOC_367 OR2X1_LOC_367/a_8_216# OR2X1_LOC_367/a_36_216# D_GATE_366 VSS VDD
+ OR2X1_LOC_366/Y OR2X1_LOC_367/B OR2X1_LOC
XOR2X1_LOC_301 OR2X1_LOC_301/a_8_216# OR2X1_LOC_301/a_36_216# OR2X1_LOC_303/B VSS VDD
+ OR2X1_LOC_831/A OR2X1_LOC_76/A OR2X1_LOC
XOR2X1_LOC_334 OR2X1_LOC_334/a_8_216# OR2X1_LOC_334/a_36_216# OR2X1_LOC_338/A VSS VDD
+ OR2X1_LOC_334/A OR2X1_LOC_334/B OR2X1_LOC
XOR2X1_LOC_323 OR2X1_LOC_323/a_8_216# OR2X1_LOC_323/a_36_216# OR2X1_LOC_323/Y VSS VDD
+ OR2X1_LOC_323/A OR2X1_LOC_95/Y OR2X1_LOC
XOR2X1_LOC_356 OR2X1_LOC_356/a_8_216# OR2X1_LOC_356/a_36_216# OR2X1_LOC_365/B VSS VDD
+ OR2X1_LOC_356/A OR2X1_LOC_356/B OR2X1_LOC
XAND2X1_LOC_570 AND2X1_LOC_570/a_36_24# AND2X1_LOC_570/Y AND2X1_LOC_570/a_8_24# VSS VDD
+ AND2X1_LOC_562/Y AND2X1_LOC_563/Y AND2X1_LOC
XAND2X1_LOC_592 AND2X1_LOC_592/a_36_24# AND2X1_LOC_592/Y AND2X1_LOC_592/a_8_24# VSS VDD
+ OR2X1_LOC_423/Y OR2X1_LOC_589/Y AND2X1_LOC
XAND2X1_LOC_581 AND2X1_LOC_581/a_36_24# AND2X1_LOC_582/B AND2X1_LOC_581/a_8_24# VSS VDD
+ INPUT_6 AND2X1_LOC_2/Y AND2X1_LOC
XOR2X1_LOC_389 OR2X1_LOC_389/a_8_216# OR2X1_LOC_389/a_36_216# OR2X1_LOC_390/A VSS VDD
+ OR2X1_LOC_389/A OR2X1_LOC_389/B OR2X1_LOC
XOR2X1_LOC_197 OR2X1_LOC_197/a_8_216# OR2X1_LOC_197/a_36_216# OR2X1_LOC_198/A VSS VDD
+ OR2X1_LOC_197/A AND2X1_LOC_52/Y OR2X1_LOC
XOR2X1_LOC_142 OR2X1_LOC_142/a_8_216# OR2X1_LOC_142/a_36_216# OR2X1_LOC_142/Y VSS VDD
+ OR2X1_LOC_64/Y OR2X1_LOC_52/B OR2X1_LOC
XOR2X1_LOC_120 OR2X1_LOC_120/a_8_216# OR2X1_LOC_120/a_36_216# OR2X1_LOC_121/A VSS VDD
+ OR2X1_LOC_154/A AND2X1_LOC_41/A OR2X1_LOC
XOR2X1_LOC_131 OR2X1_LOC_131/a_8_216# OR2X1_LOC_131/a_36_216# OR2X1_LOC_131/Y VSS VDD
+ OR2X1_LOC_131/A OR2X1_LOC_12/Y OR2X1_LOC
XOR2X1_LOC_153 OR2X1_LOC_153/a_8_216# OR2X1_LOC_153/a_36_216# OR2X1_LOC_743/A VSS VDD
+ OR2X1_LOC_85/A INPUT_1 OR2X1_LOC
XOR2X1_LOC_164 OR2X1_LOC_164/a_8_216# OR2X1_LOC_164/a_36_216# OR2X1_LOC_164/Y VSS VDD
+ OR2X1_LOC_696/A OR2X1_LOC_18/Y OR2X1_LOC
XOR2X1_LOC_175 OR2X1_LOC_175/a_8_216# OR2X1_LOC_175/a_36_216# OR2X1_LOC_175/Y VSS VDD
+ OR2X1_LOC_174/Y OR2X1_LOC_175/B OR2X1_LOC
XOR2X1_LOC_186 OR2X1_LOC_186/a_8_216# OR2X1_LOC_186/a_36_216# OR2X1_LOC_186/Y VSS VDD
+ OR2X1_LOC_185/Y OR2X1_LOC_151/A OR2X1_LOC
XOR2X1_LOC_708 OR2X1_LOC_708/a_8_216# OR2X1_LOC_708/a_36_216# OR2X1_LOC_708/Y VSS VDD
+ OR2X1_LOC_779/A OR2X1_LOC_708/B OR2X1_LOC
XOR2X1_LOC_719 OR2X1_LOC_719/a_8_216# OR2X1_LOC_719/a_36_216# OR2X1_LOC_719/Y VSS VDD
+ OR2X1_LOC_719/A OR2X1_LOC_719/B OR2X1_LOC
C0 VDD OR2X1_LOC_620/A -0.00fF
C1 OR2X1_LOC_246/Y OR2X1_LOC_585/A 0.09fF
C2 OR2X1_LOC_84/Y OR2X1_LOC_549/A 0.00fF
C3 AND2X1_LOC_729/Y AND2X1_LOC_191/Y 0.03fF
C4 AND2X1_LOC_363/A OR2X1_LOC_44/Y 0.94fF
C5 OR2X1_LOC_633/A OR2X1_LOC_598/A 0.32fF
C6 OR2X1_LOC_680/A OR2X1_LOC_89/A 0.03fF
C7 OR2X1_LOC_667/a_8_216# OR2X1_LOC_26/Y 0.01fF
C8 OR2X1_LOC_605/B OR2X1_LOC_161/A 0.01fF
C9 AND2X1_LOC_525/a_8_24# OR2X1_LOC_375/A 0.01fF
C10 OR2X1_LOC_639/A AND2X1_LOC_11/Y 0.06fF
C11 AND2X1_LOC_40/Y AND2X1_LOC_48/A 0.42fF
C12 AND2X1_LOC_548/a_36_24# AND2X1_LOC_624/A 0.01fF
C13 AND2X1_LOC_22/Y OR2X1_LOC_560/A 0.21fF
C14 OR2X1_LOC_155/A OR2X1_LOC_269/B 0.10fF
C15 OR2X1_LOC_88/A OR2X1_LOC_74/A 0.96fF
C16 OR2X1_LOC_263/a_8_216# OR2X1_LOC_92/Y 0.01fF
C17 OR2X1_LOC_755/A AND2X1_LOC_621/Y 0.10fF
C18 AND2X1_LOC_729/Y OR2X1_LOC_70/Y 0.04fF
C19 AND2X1_LOC_22/Y OR2X1_LOC_198/A 0.12fF
C20 AND2X1_LOC_214/A OR2X1_LOC_31/Y 0.02fF
C21 OR2X1_LOC_631/B OR2X1_LOC_574/A 0.02fF
C22 AND2X1_LOC_95/Y OR2X1_LOC_476/a_8_216# 0.01fF
C23 OR2X1_LOC_405/A OR2X1_LOC_121/B 0.11fF
C24 OR2X1_LOC_185/Y OR2X1_LOC_702/A 0.02fF
C25 OR2X1_LOC_43/A OR2X1_LOC_73/a_8_216# 0.03fF
C26 AND2X1_LOC_354/Y OR2X1_LOC_311/Y 0.00fF
C27 OR2X1_LOC_807/a_8_216# OR2X1_LOC_269/B 0.02fF
C28 OR2X1_LOC_648/A OR2X1_LOC_112/B 0.03fF
C29 OR2X1_LOC_856/B AND2X1_LOC_23/a_8_24# 0.06fF
C30 AND2X1_LOC_656/Y OR2X1_LOC_517/A 0.27fF
C31 OR2X1_LOC_375/A AND2X1_LOC_51/Y 1.52fF
C32 AND2X1_LOC_220/Y AND2X1_LOC_221/a_8_24# 0.00fF
C33 AND2X1_LOC_601/a_36_24# AND2X1_LOC_51/Y 0.00fF
C34 OR2X1_LOC_779/B OR2X1_LOC_713/A 0.22fF
C35 OR2X1_LOC_814/Y OR2X1_LOC_814/A 0.01fF
C36 OR2X1_LOC_64/Y OR2X1_LOC_265/Y 0.03fF
C37 AND2X1_LOC_687/Y OR2X1_LOC_48/B 0.02fF
C38 OR2X1_LOC_19/B AND2X1_LOC_233/a_8_24# 0.17fF
C39 AND2X1_LOC_717/B OR2X1_LOC_238/Y 0.03fF
C40 OR2X1_LOC_862/B AND2X1_LOC_225/a_8_24# 0.04fF
C41 AND2X1_LOC_784/A OR2X1_LOC_70/Y 0.07fF
C42 OR2X1_LOC_246/A OR2X1_LOC_595/a_8_216# 0.11fF
C43 AND2X1_LOC_727/A OR2X1_LOC_39/A 0.03fF
C44 OR2X1_LOC_18/Y AND2X1_LOC_687/Y 0.06fF
C45 OR2X1_LOC_411/Y AND2X1_LOC_461/a_8_24# 0.01fF
C46 OR2X1_LOC_43/A AND2X1_LOC_260/a_8_24# 0.01fF
C47 OR2X1_LOC_18/Y AND2X1_LOC_630/a_8_24# 0.03fF
C48 AND2X1_LOC_12/Y AND2X1_LOC_494/a_8_24# 0.02fF
C49 OR2X1_LOC_593/B OR2X1_LOC_390/B 0.02fF
C50 AND2X1_LOC_663/B OR2X1_LOC_701/a_8_216# 0.01fF
C51 INPUT_0 OR2X1_LOC_214/B 0.07fF
C52 OR2X1_LOC_36/Y AND2X1_LOC_856/a_8_24# 0.05fF
C53 OR2X1_LOC_364/A OR2X1_LOC_476/B 0.01fF
C54 OR2X1_LOC_836/Y OR2X1_LOC_375/A 0.02fF
C55 OR2X1_LOC_416/Y OR2X1_LOC_6/A 0.02fF
C56 OR2X1_LOC_813/A AND2X1_LOC_573/A 0.05fF
C57 AND2X1_LOC_769/a_8_24# OR2X1_LOC_70/Y 0.06fF
C58 OR2X1_LOC_419/Y AND2X1_LOC_663/A 0.05fF
C59 OR2X1_LOC_532/B AND2X1_LOC_617/a_8_24# 0.01fF
C60 AND2X1_LOC_784/A AND2X1_LOC_514/Y 0.04fF
C61 OR2X1_LOC_600/A OR2X1_LOC_749/a_36_216# 0.00fF
C62 OR2X1_LOC_193/A AND2X1_LOC_3/Y 0.23fF
C63 AND2X1_LOC_53/Y AND2X1_LOC_43/B 1.01fF
C64 OR2X1_LOC_485/A OR2X1_LOC_481/A 0.01fF
C65 AND2X1_LOC_124/a_8_24# AND2X1_LOC_845/Y 0.03fF
C66 OR2X1_LOC_673/Y OR2X1_LOC_62/B 0.02fF
C67 OR2X1_LOC_685/a_36_216# AND2X1_LOC_425/Y 0.00fF
C68 AND2X1_LOC_91/B OR2X1_LOC_703/Y 0.00fF
C69 AND2X1_LOC_64/Y OR2X1_LOC_714/a_8_216# 0.01fF
C70 OR2X1_LOC_36/Y OR2X1_LOC_7/Y 0.01fF
C71 AND2X1_LOC_508/B AND2X1_LOC_657/A 0.00fF
C72 OR2X1_LOC_109/Y AND2X1_LOC_318/Y 0.02fF
C73 AND2X1_LOC_348/a_8_24# OR2X1_LOC_481/A 0.17fF
C74 OR2X1_LOC_95/Y OR2X1_LOC_39/A 0.14fF
C75 AND2X1_LOC_440/a_8_24# OR2X1_LOC_39/A 0.14fF
C76 AND2X1_LOC_866/A AND2X1_LOC_848/Y 0.08fF
C77 AND2X1_LOC_508/a_8_24# AND2X1_LOC_657/A 0.02fF
C78 AND2X1_LOC_738/B AND2X1_LOC_796/A 0.10fF
C79 OR2X1_LOC_431/a_36_216# OR2X1_LOC_304/Y 0.00fF
C80 OR2X1_LOC_849/A OR2X1_LOC_532/B 0.02fF
C81 OR2X1_LOC_223/A AND2X1_LOC_43/B 0.03fF
C82 OR2X1_LOC_59/Y OR2X1_LOC_172/Y 0.01fF
C83 AND2X1_LOC_849/a_8_24# AND2X1_LOC_806/A 0.01fF
C84 OR2X1_LOC_736/A OR2X1_LOC_675/Y 0.04fF
C85 OR2X1_LOC_12/Y D_INPUT_6 0.41fF
C86 AND2X1_LOC_663/A OR2X1_LOC_152/A 0.03fF
C87 AND2X1_LOC_55/a_8_24# D_INPUT_3 0.26fF
C88 OR2X1_LOC_8/Y OR2X1_LOC_71/A 0.32fF
C89 OR2X1_LOC_244/B OR2X1_LOC_560/A 0.02fF
C90 D_INPUT_0 AND2X1_LOC_3/Y 0.54fF
C91 AND2X1_LOC_386/a_8_24# AND2X1_LOC_7/Y 0.21fF
C92 OR2X1_LOC_362/A OR2X1_LOC_349/B 0.02fF
C93 OR2X1_LOC_94/a_8_216# D_INPUT_1 0.01fF
C94 OR2X1_LOC_70/Y AND2X1_LOC_639/A 0.04fF
C95 OR2X1_LOC_485/A OR2X1_LOC_71/Y 0.09fF
C96 AND2X1_LOC_850/A AND2X1_LOC_657/A 0.07fF
C97 OR2X1_LOC_31/Y AND2X1_LOC_645/A 0.00fF
C98 OR2X1_LOC_92/Y AND2X1_LOC_562/Y 0.05fF
C99 AND2X1_LOC_348/Y OR2X1_LOC_47/Y 0.03fF
C100 OR2X1_LOC_151/A OR2X1_LOC_308/Y 0.07fF
C101 OR2X1_LOC_185/A OR2X1_LOC_192/B 0.31fF
C102 OR2X1_LOC_619/Y AND2X1_LOC_647/Y 0.03fF
C103 OR2X1_LOC_476/B OR2X1_LOC_472/B 0.01fF
C104 VDD OR2X1_LOC_217/A 0.00fF
C105 OR2X1_LOC_47/Y OR2X1_LOC_753/A 0.05fF
C106 OR2X1_LOC_685/B AND2X1_LOC_418/a_8_24# 0.20fF
C107 OR2X1_LOC_680/A AND2X1_LOC_804/a_8_24# 0.03fF
C108 AND2X1_LOC_784/A OR2X1_LOC_437/Y 0.31fF
C109 OR2X1_LOC_617/Y AND2X1_LOC_866/A 0.02fF
C110 OR2X1_LOC_47/Y OR2X1_LOC_754/a_8_216# 0.01fF
C111 AND2X1_LOC_544/Y AND2X1_LOC_212/Y 0.19fF
C112 OR2X1_LOC_696/A OR2X1_LOC_6/B 0.07fF
C113 AND2X1_LOC_110/Y OR2X1_LOC_354/a_8_216# 0.01fF
C114 OR2X1_LOC_502/A AND2X1_LOC_406/a_36_24# 0.01fF
C115 AND2X1_LOC_74/a_36_24# OR2X1_LOC_578/B 0.01fF
C116 AND2X1_LOC_56/B AND2X1_LOC_699/a_8_24# 0.01fF
C117 OR2X1_LOC_696/A AND2X1_LOC_713/Y 0.01fF
C118 OR2X1_LOC_808/B OR2X1_LOC_303/B 0.05fF
C119 OR2X1_LOC_589/A AND2X1_LOC_773/a_8_24# 0.17fF
C120 AND2X1_LOC_130/a_8_24# AND2X1_LOC_772/Y 0.14fF
C121 OR2X1_LOC_485/A D_INPUT_1 0.02fF
C122 OR2X1_LOC_448/Y AND2X1_LOC_31/Y 0.01fF
C123 AND2X1_LOC_91/B OR2X1_LOC_596/A 0.56fF
C124 AND2X1_LOC_707/Y OR2X1_LOC_12/Y 0.13fF
C125 AND2X1_LOC_56/B OR2X1_LOC_675/Y 0.02fF
C126 AND2X1_LOC_22/Y OR2X1_LOC_435/A 0.08fF
C127 OR2X1_LOC_778/Y OR2X1_LOC_374/Y 0.02fF
C128 OR2X1_LOC_158/A OR2X1_LOC_56/Y 0.03fF
C129 AND2X1_LOC_64/Y OR2X1_LOC_6/B 0.16fF
C130 AND2X1_LOC_785/Y AND2X1_LOC_795/a_8_24# -0.00fF
C131 OR2X1_LOC_22/Y AND2X1_LOC_293/a_8_24# 0.03fF
C132 AND2X1_LOC_196/Y AND2X1_LOC_199/a_8_24# 0.03fF
C133 OR2X1_LOC_709/A OR2X1_LOC_691/Y 0.00fF
C134 AND2X1_LOC_340/Y OR2X1_LOC_16/A 0.03fF
C135 OR2X1_LOC_804/a_36_216# OR2X1_LOC_593/B 0.00fF
C136 OR2X1_LOC_792/Y OR2X1_LOC_580/A 0.01fF
C137 AND2X1_LOC_477/A OR2X1_LOC_31/Y 0.10fF
C138 AND2X1_LOC_849/A OR2X1_LOC_224/Y 0.14fF
C139 AND2X1_LOC_706/Y AND2X1_LOC_714/a_8_24# 0.02fF
C140 OR2X1_LOC_215/Y AND2X1_LOC_406/a_8_24# 0.10fF
C141 AND2X1_LOC_773/Y OR2X1_LOC_589/A 1.48fF
C142 OR2X1_LOC_625/Y OR2X1_LOC_437/A 0.24fF
C143 AND2X1_LOC_633/Y AND2X1_LOC_476/A 0.01fF
C144 OR2X1_LOC_6/A OR2X1_LOC_80/A 0.14fF
C145 OR2X1_LOC_532/B OR2X1_LOC_440/A 0.03fF
C146 D_INPUT_0 AND2X1_LOC_476/A 0.07fF
C147 OR2X1_LOC_97/A OR2X1_LOC_832/a_8_216# 0.01fF
C148 OR2X1_LOC_161/A OR2X1_LOC_515/Y 0.16fF
C149 OR2X1_LOC_175/Y AND2X1_LOC_70/Y 0.10fF
C150 OR2X1_LOC_193/Y OR2X1_LOC_193/a_8_216# 0.01fF
C151 AND2X1_LOC_460/a_8_24# OR2X1_LOC_22/A 0.01fF
C152 OR2X1_LOC_160/B OR2X1_LOC_61/A 0.10fF
C153 OR2X1_LOC_319/B OR2X1_LOC_354/a_36_216# 0.01fF
C154 OR2X1_LOC_6/B AND2X1_LOC_82/Y 0.02fF
C155 OR2X1_LOC_40/Y OR2X1_LOC_135/Y 0.01fF
C156 OR2X1_LOC_464/B OR2X1_LOC_367/B 0.01fF
C157 OR2X1_LOC_426/B AND2X1_LOC_636/a_8_24# 0.17fF
C158 AND2X1_LOC_191/B GATE_579 0.01fF
C159 OR2X1_LOC_47/Y AND2X1_LOC_845/Y 0.02fF
C160 OR2X1_LOC_628/Y AND2X1_LOC_624/B 0.15fF
C161 AND2X1_LOC_469/B AND2X1_LOC_794/a_8_24# 0.01fF
C162 OR2X1_LOC_833/B AND2X1_LOC_36/Y 0.08fF
C163 OR2X1_LOC_95/Y OR2X1_LOC_760/a_8_216# 0.01fF
C164 AND2X1_LOC_59/Y OR2X1_LOC_535/a_8_216# 0.14fF
C165 OR2X1_LOC_160/B OR2X1_LOC_659/Y 0.04fF
C166 AND2X1_LOC_70/Y OR2X1_LOC_691/Y 0.05fF
C167 OR2X1_LOC_599/A OR2X1_LOC_536/a_8_216# 0.00fF
C168 OR2X1_LOC_479/Y OR2X1_LOC_353/a_8_216# 0.03fF
C169 OR2X1_LOC_59/Y AND2X1_LOC_206/a_8_24# 0.17fF
C170 OR2X1_LOC_84/B OR2X1_LOC_71/A 0.00fF
C171 OR2X1_LOC_517/A AND2X1_LOC_772/Y 0.51fF
C172 OR2X1_LOC_34/B OR2X1_LOC_598/A 0.10fF
C173 OR2X1_LOC_70/Y OR2X1_LOC_88/Y 0.02fF
C174 AND2X1_LOC_454/A OR2X1_LOC_423/Y 0.01fF
C175 AND2X1_LOC_69/Y OR2X1_LOC_68/B 0.04fF
C176 AND2X1_LOC_181/Y OR2X1_LOC_108/Y 0.81fF
C177 AND2X1_LOC_474/A AND2X1_LOC_287/B 0.01fF
C178 OR2X1_LOC_70/Y OR2X1_LOC_172/Y 0.31fF
C179 OR2X1_LOC_608/a_8_216# OR2X1_LOC_502/Y 0.39fF
C180 OR2X1_LOC_189/Y AND2X1_LOC_738/Y 0.11fF
C181 AND2X1_LOC_218/Y AND2X1_LOC_786/Y 0.04fF
C182 AND2X1_LOC_339/B AND2X1_LOC_61/Y 0.23fF
C183 OR2X1_LOC_507/B OR2X1_LOC_508/Y 0.01fF
C184 OR2X1_LOC_62/A AND2X1_LOC_14/a_8_24# 0.20fF
C185 OR2X1_LOC_6/B AND2X1_LOC_86/a_8_24# 0.11fF
C186 OR2X1_LOC_254/B AND2X1_LOC_36/Y 0.01fF
C187 OR2X1_LOC_326/B AND2X1_LOC_64/Y 0.03fF
C188 OR2X1_LOC_51/Y AND2X1_LOC_605/a_8_24# 0.01fF
C189 OR2X1_LOC_604/A OR2X1_LOC_96/Y 0.07fF
C190 OR2X1_LOC_40/Y OR2X1_LOC_815/a_8_216# 0.01fF
C191 OR2X1_LOC_750/A OR2X1_LOC_228/Y 0.10fF
C192 OR2X1_LOC_648/B OR2X1_LOC_66/A 0.11fF
C193 OR2X1_LOC_97/A OR2X1_LOC_634/a_36_216# 0.00fF
C194 OR2X1_LOC_40/Y AND2X1_LOC_98/a_8_24# 0.01fF
C195 OR2X1_LOC_177/Y AND2X1_LOC_663/A 0.03fF
C196 AND2X1_LOC_285/a_8_24# OR2X1_LOC_56/A 0.00fF
C197 VDD OR2X1_LOC_450/Y -0.00fF
C198 OR2X1_LOC_696/A AND2X1_LOC_436/B 0.00fF
C199 AND2X1_LOC_548/a_8_24# OR2X1_LOC_437/A 0.03fF
C200 OR2X1_LOC_185/A OR2X1_LOC_502/Y 0.22fF
C201 AND2X1_LOC_486/Y AND2X1_LOC_721/Y 0.03fF
C202 OR2X1_LOC_814/A OR2X1_LOC_641/B 0.00fF
C203 AND2X1_LOC_91/B OR2X1_LOC_732/a_8_216# 0.04fF
C204 AND2X1_LOC_388/Y AND2X1_LOC_434/Y 0.13fF
C205 AND2X1_LOC_565/B AND2X1_LOC_565/a_8_24# 0.01fF
C206 VDD AND2X1_LOC_508/B 0.27fF
C207 AND2X1_LOC_3/Y OR2X1_LOC_339/A 1.32fF
C208 VDD OR2X1_LOC_679/Y -0.00fF
C209 OR2X1_LOC_566/A OR2X1_LOC_212/A 0.02fF
C210 AND2X1_LOC_12/Y OR2X1_LOC_308/A 0.03fF
C211 OR2X1_LOC_40/Y AND2X1_LOC_443/Y 0.00fF
C212 OR2X1_LOC_132/a_8_216# VDD 0.21fF
C213 OR2X1_LOC_646/A AND2X1_LOC_36/Y 0.06fF
C214 OR2X1_LOC_45/B OR2X1_LOC_427/A 0.15fF
C215 OR2X1_LOC_668/a_8_216# AND2X1_LOC_44/Y 0.01fF
C216 OR2X1_LOC_382/Y OR2X1_LOC_158/A 0.01fF
C217 OR2X1_LOC_604/A AND2X1_LOC_663/A 0.14fF
C218 OR2X1_LOC_56/A OR2X1_LOC_627/Y 0.01fF
C219 AND2X1_LOC_64/Y OR2X1_LOC_579/B 0.18fF
C220 AND2X1_LOC_12/Y OR2X1_LOC_866/B 0.16fF
C221 OR2X1_LOC_160/B AND2X1_LOC_24/a_8_24# 0.00fF
C222 AND2X1_LOC_715/Y AND2X1_LOC_436/B 0.02fF
C223 OR2X1_LOC_502/A OR2X1_LOC_356/A 0.20fF
C224 OR2X1_LOC_858/B OR2X1_LOC_362/A 0.02fF
C225 AND2X1_LOC_51/Y OR2X1_LOC_515/Y 0.65fF
C226 OR2X1_LOC_329/B AND2X1_LOC_112/a_8_24# 0.05fF
C227 OR2X1_LOC_8/Y OR2X1_LOC_59/Y 0.04fF
C228 OR2X1_LOC_124/A AND2X1_LOC_70/Y 0.28fF
C229 OR2X1_LOC_48/B OR2X1_LOC_373/Y 0.02fF
C230 OR2X1_LOC_379/Y OR2X1_LOC_855/a_8_216# 0.01fF
C231 AND2X1_LOC_716/Y OR2X1_LOC_309/a_8_216# 0.03fF
C232 AND2X1_LOC_374/a_8_24# AND2X1_LOC_476/Y 0.02fF
C233 AND2X1_LOC_810/A OR2X1_LOC_619/Y 0.05fF
C234 OR2X1_LOC_18/Y OR2X1_LOC_373/Y 0.00fF
C235 AND2X1_LOC_486/Y OR2X1_LOC_482/Y 0.07fF
C236 OR2X1_LOC_92/Y AND2X1_LOC_448/a_8_24# 0.02fF
C237 OR2X1_LOC_106/Y AND2X1_LOC_361/A 0.74fF
C238 OR2X1_LOC_696/A OR2X1_LOC_529/Y 0.03fF
C239 AND2X1_LOC_655/A OR2X1_LOC_428/A 0.10fF
C240 OR2X1_LOC_709/A AND2X1_LOC_699/a_36_24# 0.00fF
C241 VDD AND2X1_LOC_850/A 0.17fF
C242 OR2X1_LOC_427/A OR2X1_LOC_382/A 0.17fF
C243 AND2X1_LOC_550/A AND2X1_LOC_212/Y 0.07fF
C244 AND2X1_LOC_194/Y OR2X1_LOC_16/Y 0.00fF
C245 OR2X1_LOC_185/A AND2X1_LOC_603/a_36_24# 0.00fF
C246 OR2X1_LOC_121/a_8_216# OR2X1_LOC_375/A 0.01fF
C247 VDD OR2X1_LOC_708/Y -0.00fF
C248 GATE_479 GATE_222 0.03fF
C249 OR2X1_LOC_45/B AND2X1_LOC_464/a_8_24# 0.00fF
C250 D_INPUT_2 OR2X1_LOC_80/A 0.16fF
C251 AND2X1_LOC_91/B AND2X1_LOC_399/a_36_24# 0.01fF
C252 OR2X1_LOC_808/A OR2X1_LOC_645/a_8_216# 0.01fF
C253 OR2X1_LOC_240/B OR2X1_LOC_549/A 0.03fF
C254 OR2X1_LOC_643/A OR2X1_LOC_392/B 0.05fF
C255 AND2X1_LOC_228/Y OR2X1_LOC_16/A 0.13fF
C256 OR2X1_LOC_85/A OR2X1_LOC_79/Y 0.04fF
C257 OR2X1_LOC_697/Y OR2X1_LOC_743/a_8_216# 0.01fF
C258 OR2X1_LOC_45/B OR2X1_LOC_271/a_8_216# 0.01fF
C259 AND2X1_LOC_82/a_8_24# OR2X1_LOC_633/A 0.03fF
C260 OR2X1_LOC_161/A OR2X1_LOC_549/A 0.03fF
C261 OR2X1_LOC_87/A AND2X1_LOC_44/Y 0.48fF
C262 VDD OR2X1_LOC_608/a_8_216# 0.00fF
C263 OR2X1_LOC_158/A AND2X1_LOC_375/a_36_24# 0.01fF
C264 AND2X1_LOC_91/B AND2X1_LOC_85/a_8_24# 0.01fF
C265 OR2X1_LOC_848/A OR2X1_LOC_489/A 0.01fF
C266 OR2X1_LOC_857/B AND2X1_LOC_824/a_8_24# 0.01fF
C267 OR2X1_LOC_255/a_36_216# OR2X1_LOC_13/B 0.00fF
C268 OR2X1_LOC_691/A OR2X1_LOC_835/B 0.01fF
C269 OR2X1_LOC_631/B AND2X1_LOC_627/a_8_24# 0.03fF
C270 OR2X1_LOC_292/Y OR2X1_LOC_91/A 0.08fF
C271 AND2X1_LOC_773/Y OR2X1_LOC_43/A 0.17fF
C272 AND2X1_LOC_696/a_8_24# AND2X1_LOC_44/Y 0.01fF
C273 OR2X1_LOC_496/Y AND2X1_LOC_785/Y 0.27fF
C274 AND2X1_LOC_94/Y AND2X1_LOC_402/a_8_24# 0.20fF
C275 OR2X1_LOC_128/a_36_216# OR2X1_LOC_151/A 0.01fF
C276 AND2X1_LOC_555/Y OR2X1_LOC_282/Y 0.01fF
C277 OR2X1_LOC_684/a_8_216# OR2X1_LOC_427/A 0.01fF
C278 OR2X1_LOC_406/Y AND2X1_LOC_475/a_8_24# -0.00fF
C279 OR2X1_LOC_223/A OR2X1_LOC_367/B 0.03fF
C280 AND2X1_LOC_56/B OR2X1_LOC_736/Y 0.03fF
C281 OR2X1_LOC_40/Y AND2X1_LOC_175/B 0.12fF
C282 OR2X1_LOC_475/a_8_216# OR2X1_LOC_78/A 0.02fF
C283 OR2X1_LOC_666/a_8_216# OR2X1_LOC_18/Y 0.07fF
C284 AND2X1_LOC_19/a_8_24# AND2X1_LOC_44/Y 0.05fF
C285 VDD OR2X1_LOC_185/A 1.01fF
C286 OR2X1_LOC_510/Y AND2X1_LOC_625/a_8_24# 0.00fF
C287 OR2X1_LOC_40/Y AND2X1_LOC_848/Y 0.15fF
C288 OR2X1_LOC_585/A OR2X1_LOC_16/A 0.21fF
C289 OR2X1_LOC_604/A AND2X1_LOC_449/Y 0.00fF
C290 AND2X1_LOC_59/Y AND2X1_LOC_313/a_8_24# 0.02fF
C291 VDD OR2X1_LOC_249/Y 0.24fF
C292 OR2X1_LOC_643/A OR2X1_LOC_113/B 1.62fF
C293 AND2X1_LOC_568/B AND2X1_LOC_365/A 0.00fF
C294 AND2X1_LOC_76/Y OR2X1_LOC_59/Y 0.04fF
C295 OR2X1_LOC_848/A OR2X1_LOC_772/A 0.01fF
C296 AND2X1_LOC_337/B AND2X1_LOC_802/Y 0.04fF
C297 OR2X1_LOC_135/Y OR2X1_LOC_7/A 0.07fF
C298 OR2X1_LOC_774/B AND2X1_LOC_236/a_8_24# 0.27fF
C299 AND2X1_LOC_729/Y AND2X1_LOC_658/B 0.03fF
C300 OR2X1_LOC_112/B OR2X1_LOC_112/A 0.10fF
C301 AND2X1_LOC_162/a_8_24# OR2X1_LOC_619/Y 0.00fF
C302 AND2X1_LOC_578/A AND2X1_LOC_786/Y 0.07fF
C303 OR2X1_LOC_474/Y OR2X1_LOC_475/B 0.00fF
C304 OR2X1_LOC_754/A OR2X1_LOC_753/a_36_216# 0.00fF
C305 OR2X1_LOC_43/A AND2X1_LOC_243/Y 0.07fF
C306 AND2X1_LOC_706/Y OR2X1_LOC_743/A 0.05fF
C307 OR2X1_LOC_770/A OR2X1_LOC_401/B 0.05fF
C308 AND2X1_LOC_766/a_36_24# OR2X1_LOC_401/A 0.00fF
C309 AND2X1_LOC_303/A OR2X1_LOC_426/B 0.13fF
C310 AND2X1_LOC_217/Y OR2X1_LOC_26/Y 0.03fF
C311 AND2X1_LOC_65/a_36_24# OR2X1_LOC_61/Y -0.02fF
C312 OR2X1_LOC_113/Y OR2X1_LOC_161/A 0.00fF
C313 OR2X1_LOC_533/a_8_216# OR2X1_LOC_331/a_8_216# 0.47fF
C314 OR2X1_LOC_492/Y OR2X1_LOC_485/A 0.01fF
C315 AND2X1_LOC_64/Y OR2X1_LOC_68/Y 0.03fF
C316 OR2X1_LOC_810/A AND2X1_LOC_625/a_8_24# 0.18fF
C317 OR2X1_LOC_482/Y OR2X1_LOC_666/Y 0.02fF
C318 AND2X1_LOC_95/Y OR2X1_LOC_634/A 0.18fF
C319 OR2X1_LOC_646/a_8_216# OR2X1_LOC_646/B 0.02fF
C320 AND2X1_LOC_83/a_8_24# OR2X1_LOC_624/B 0.02fF
C321 OR2X1_LOC_405/A OR2X1_LOC_317/a_8_216# 0.01fF
C322 OR2X1_LOC_219/a_36_216# AND2X1_LOC_92/Y 0.00fF
C323 OR2X1_LOC_814/A OR2X1_LOC_227/A 0.01fF
C324 OR2X1_LOC_377/A AND2X1_LOC_41/A 0.84fF
C325 AND2X1_LOC_168/Y OR2X1_LOC_165/Y 0.80fF
C326 VDD OR2X1_LOC_117/Y 0.04fF
C327 AND2X1_LOC_732/a_8_24# OR2X1_LOC_44/Y 0.01fF
C328 OR2X1_LOC_326/a_36_216# AND2X1_LOC_59/Y 0.00fF
C329 OR2X1_LOC_34/B OR2X1_LOC_34/A 0.16fF
C330 VDD OR2X1_LOC_498/Y 0.18fF
C331 OR2X1_LOC_598/Y AND2X1_LOC_3/Y 0.04fF
C332 OR2X1_LOC_863/a_8_216# OR2X1_LOC_35/Y 0.01fF
C333 OR2X1_LOC_78/A OR2X1_LOC_779/a_8_216# 0.01fF
C334 OR2X1_LOC_466/A OR2X1_LOC_449/A 0.14fF
C335 OR2X1_LOC_108/a_8_216# OR2X1_LOC_485/A 0.01fF
C336 OR2X1_LOC_641/Y AND2X1_LOC_8/Y 0.15fF
C337 AND2X1_LOC_217/Y OR2X1_LOC_89/A 0.03fF
C338 OR2X1_LOC_832/a_36_216# OR2X1_LOC_155/A 0.00fF
C339 AND2X1_LOC_729/B OR2X1_LOC_829/A 0.10fF
C340 AND2X1_LOC_191/Y AND2X1_LOC_478/a_36_24# 0.01fF
C341 AND2X1_LOC_64/Y AND2X1_LOC_47/Y 0.57fF
C342 OR2X1_LOC_45/B AND2X1_LOC_687/B 0.04fF
C343 OR2X1_LOC_51/Y AND2X1_LOC_853/Y 0.31fF
C344 OR2X1_LOC_354/A OR2X1_LOC_161/A 0.63fF
C345 AND2X1_LOC_593/a_36_24# OR2X1_LOC_89/A 0.00fF
C346 AND2X1_LOC_42/B OR2X1_LOC_641/A 0.03fF
C347 AND2X1_LOC_51/Y OR2X1_LOC_549/A 0.07fF
C348 OR2X1_LOC_235/B OR2X1_LOC_720/A 0.01fF
C349 OR2X1_LOC_683/a_8_216# AND2X1_LOC_452/Y 0.01fF
C350 AND2X1_LOC_727/A AND2X1_LOC_727/B 0.33fF
C351 AND2X1_LOC_702/Y OR2X1_LOC_91/A 0.03fF
C352 AND2X1_LOC_38/a_8_24# AND2X1_LOC_18/Y 0.01fF
C353 OR2X1_LOC_604/A OR2X1_LOC_617/a_8_216# 0.15fF
C354 OR2X1_LOC_405/A OR2X1_LOC_856/B 0.07fF
C355 OR2X1_LOC_502/A AND2X1_LOC_43/B 0.26fF
C356 AND2X1_LOC_392/A AND2X1_LOC_276/Y 0.03fF
C357 OR2X1_LOC_40/Y OR2X1_LOC_617/Y 0.06fF
C358 AND2X1_LOC_41/A OR2X1_LOC_203/Y 0.07fF
C359 AND2X1_LOC_377/Y OR2X1_LOC_43/A 0.10fF
C360 OR2X1_LOC_323/A AND2X1_LOC_270/a_36_24# 0.00fF
C361 OR2X1_LOC_59/Y OR2X1_LOC_52/B 0.27fF
C362 OR2X1_LOC_706/B AND2X1_LOC_44/Y 0.01fF
C363 OR2X1_LOC_574/A OR2X1_LOC_648/A 0.10fF
C364 OR2X1_LOC_7/A AND2X1_LOC_454/a_36_24# 0.00fF
C365 AND2X1_LOC_527/a_36_24# OR2X1_LOC_620/Y 0.00fF
C366 OR2X1_LOC_426/B OR2X1_LOC_485/A 0.06fF
C367 OR2X1_LOC_849/A OR2X1_LOC_624/Y 0.01fF
C368 AND2X1_LOC_40/Y OR2X1_LOC_350/a_8_216# 0.14fF
C369 OR2X1_LOC_693/Y OR2X1_LOC_22/Y 0.11fF
C370 AND2X1_LOC_634/Y OR2X1_LOC_16/A 0.01fF
C371 OR2X1_LOC_532/B OR2X1_LOC_721/a_8_216# 0.01fF
C372 AND2X1_LOC_194/a_8_24# OR2X1_LOC_36/Y 0.01fF
C373 OR2X1_LOC_859/a_8_216# OR2X1_LOC_859/B 0.00fF
C374 OR2X1_LOC_637/a_8_216# OR2X1_LOC_828/B 0.01fF
C375 VDD OR2X1_LOC_435/Y 0.12fF
C376 OR2X1_LOC_808/B AND2X1_LOC_56/B 0.10fF
C377 AND2X1_LOC_266/a_8_24# AND2X1_LOC_266/Y 0.03fF
C378 OR2X1_LOC_757/A OR2X1_LOC_89/A 0.73fF
C379 OR2X1_LOC_51/Y OR2X1_LOC_17/Y 1.58fF
C380 OR2X1_LOC_154/A AND2X1_LOC_173/a_8_24# 0.06fF
C381 OR2X1_LOC_756/B OR2X1_LOC_389/B 0.00fF
C382 AND2X1_LOC_139/a_8_24# AND2X1_LOC_361/A 0.03fF
C383 OR2X1_LOC_3/Y AND2X1_LOC_434/Y 0.00fF
C384 AND2X1_LOC_703/Y OR2X1_LOC_31/Y 0.00fF
C385 OR2X1_LOC_61/a_36_216# OR2X1_LOC_358/B 0.00fF
C386 OR2X1_LOC_3/Y AND2X1_LOC_219/Y 0.07fF
C387 VDD AND2X1_LOC_523/Y 0.37fF
C388 OR2X1_LOC_113/A OR2X1_LOC_113/B 0.00fF
C389 OR2X1_LOC_235/B OR2X1_LOC_278/a_8_216# 0.01fF
C390 AND2X1_LOC_176/a_8_24# OR2X1_LOC_78/A 0.01fF
C391 OR2X1_LOC_185/A OR2X1_LOC_223/B 0.13fF
C392 OR2X1_LOC_214/B OR2X1_LOC_214/A 0.06fF
C393 VDD AND2X1_LOC_119/a_8_24# -0.00fF
C394 AND2X1_LOC_784/A AND2X1_LOC_357/a_8_24# 0.04fF
C395 AND2X1_LOC_453/a_8_24# AND2X1_LOC_452/Y 0.02fF
C396 OR2X1_LOC_358/a_8_216# OR2X1_LOC_624/A 0.11fF
C397 OR2X1_LOC_755/A OR2X1_LOC_59/Y 0.05fF
C398 OR2X1_LOC_283/Y AND2X1_LOC_843/Y 0.80fF
C399 INPUT_0 OR2X1_LOC_193/A 0.04fF
C400 OR2X1_LOC_684/a_8_216# AND2X1_LOC_687/B 0.47fF
C401 OR2X1_LOC_436/Y OR2X1_LOC_390/A 0.01fF
C402 AND2X1_LOC_348/Y OR2X1_LOC_625/Y 0.02fF
C403 OR2X1_LOC_70/Y OR2X1_LOC_674/a_36_216# 0.02fF
C404 AND2X1_LOC_40/Y AND2X1_LOC_3/Y 0.20fF
C405 AND2X1_LOC_40/Y OR2X1_LOC_647/B 0.78fF
C406 VDD OR2X1_LOC_815/A -0.00fF
C407 AND2X1_LOC_64/Y OR2X1_LOC_598/A 0.15fF
C408 OR2X1_LOC_625/Y OR2X1_LOC_753/A 0.17fF
C409 AND2X1_LOC_724/A AND2X1_LOC_648/B 0.00fF
C410 AND2X1_LOC_91/B OR2X1_LOC_374/Y 0.08fF
C411 OR2X1_LOC_589/A OR2X1_LOC_72/a_36_216# 0.00fF
C412 AND2X1_LOC_7/B OR2X1_LOC_241/B 2.12fF
C413 OR2X1_LOC_201/A OR2X1_LOC_475/Y 0.02fF
C414 AND2X1_LOC_100/a_8_24# OR2X1_LOC_18/Y 0.03fF
C415 OR2X1_LOC_647/a_8_216# OR2X1_LOC_78/B 0.02fF
C416 AND2X1_LOC_70/Y OR2X1_LOC_750/a_8_216# 0.00fF
C417 VDD AND2X1_LOC_431/a_8_24# 0.00fF
C418 OR2X1_LOC_633/A D_INPUT_1 0.04fF
C419 AND2X1_LOC_12/Y OR2X1_LOC_847/B 0.04fF
C420 OR2X1_LOC_744/A AND2X1_LOC_465/Y 0.02fF
C421 AND2X1_LOC_392/A AND2X1_LOC_831/Y 0.07fF
C422 AND2X1_LOC_365/a_8_24# AND2X1_LOC_514/Y 0.03fF
C423 OR2X1_LOC_117/a_36_216# OR2X1_LOC_67/Y 0.00fF
C424 OR2X1_LOC_625/Y OR2X1_LOC_754/a_8_216# 0.02fF
C425 OR2X1_LOC_354/A AND2X1_LOC_51/Y 0.09fF
C426 OR2X1_LOC_164/Y OR2X1_LOC_64/Y 0.40fF
C427 OR2X1_LOC_536/Y OR2X1_LOC_95/Y 0.02fF
C428 AND2X1_LOC_175/B OR2X1_LOC_7/A 0.00fF
C429 OR2X1_LOC_440/B OR2X1_LOC_440/A 0.16fF
C430 OR2X1_LOC_280/a_8_216# OR2X1_LOC_237/a_8_216# 0.47fF
C431 OR2X1_LOC_155/A OR2X1_LOC_539/Y 0.03fF
C432 OR2X1_LOC_673/a_8_216# D_INPUT_1 0.01fF
C433 OR2X1_LOC_305/a_8_216# OR2X1_LOC_305/Y 0.00fF
C434 OR2X1_LOC_430/a_8_216# OR2X1_LOC_427/A 0.01fF
C435 AND2X1_LOC_56/B OR2X1_LOC_82/a_8_216# 0.06fF
C436 OR2X1_LOC_455/a_8_216# OR2X1_LOC_457/B 0.05fF
C437 OR2X1_LOC_70/Y AND2X1_LOC_76/Y 0.03fF
C438 OR2X1_LOC_7/A AND2X1_LOC_848/Y 0.07fF
C439 AND2X1_LOC_120/a_8_24# AND2X1_LOC_850/Y 0.03fF
C440 INPUT_0 D_INPUT_0 0.59fF
C441 AND2X1_LOC_12/Y OR2X1_LOC_557/A 0.11fF
C442 OR2X1_LOC_714/A OR2X1_LOC_308/Y 0.03fF
C443 AND2X1_LOC_547/Y OR2X1_LOC_47/Y 0.02fF
C444 AND2X1_LOC_3/Y OR2X1_LOC_87/Y 0.00fF
C445 AND2X1_LOC_154/a_36_24# OR2X1_LOC_7/A 0.01fF
C446 OR2X1_LOC_299/a_8_216# OR2X1_LOC_6/A 0.01fF
C447 OR2X1_LOC_406/A AND2X1_LOC_795/a_36_24# 0.00fF
C448 AND2X1_LOC_673/a_36_24# OR2X1_LOC_6/A 0.00fF
C449 OR2X1_LOC_789/B OR2X1_LOC_193/A 0.13fF
C450 OR2X1_LOC_377/A AND2X1_LOC_135/a_8_24# 0.01fF
C451 AND2X1_LOC_367/a_8_24# OR2X1_LOC_485/A 0.01fF
C452 AND2X1_LOC_355/a_8_24# OR2X1_LOC_43/A 0.01fF
C453 AND2X1_LOC_349/B AND2X1_LOC_359/B 0.31fF
C454 AND2X1_LOC_359/B OR2X1_LOC_89/A 0.03fF
C455 AND2X1_LOC_47/Y AND2X1_LOC_819/a_8_24# 0.10fF
C456 OR2X1_LOC_164/Y OR2X1_LOC_417/A 0.07fF
C457 OR2X1_LOC_315/Y AND2X1_LOC_523/Y 0.02fF
C458 OR2X1_LOC_788/B OR2X1_LOC_605/Y 0.02fF
C459 OR2X1_LOC_473/Y OR2X1_LOC_805/A 0.00fF
C460 OR2X1_LOC_18/Y AND2X1_LOC_849/A 0.04fF
C461 OR2X1_LOC_748/A AND2X1_LOC_347/a_8_24# 0.01fF
C462 OR2X1_LOC_553/a_8_216# OR2X1_LOC_563/B 0.00fF
C463 OR2X1_LOC_479/Y OR2X1_LOC_469/a_8_216# 0.03fF
C464 OR2X1_LOC_306/Y AND2X1_LOC_856/a_8_24# 0.00fF
C465 OR2X1_LOC_512/A AND2X1_LOC_47/Y 0.01fF
C466 AND2X1_LOC_727/A AND2X1_LOC_593/Y 0.01fF
C467 OR2X1_LOC_774/Y OR2X1_LOC_864/a_36_216# 0.00fF
C468 AND2X1_LOC_733/a_8_24# OR2X1_LOC_95/Y 0.04fF
C469 AND2X1_LOC_95/Y OR2X1_LOC_335/B 0.36fF
C470 OR2X1_LOC_377/A OR2X1_LOC_403/a_8_216# 0.04fF
C471 AND2X1_LOC_662/B INPUT_1 0.07fF
C472 AND2X1_LOC_48/A AND2X1_LOC_43/B 0.13fF
C473 OR2X1_LOC_70/Y OR2X1_LOC_52/B 0.16fF
C474 AND2X1_LOC_91/B OR2X1_LOC_532/a_36_216# 0.00fF
C475 OR2X1_LOC_485/A OR2X1_LOC_743/A 2.04fF
C476 OR2X1_LOC_557/A AND2X1_LOC_79/Y 0.00fF
C477 AND2X1_LOC_831/a_8_24# OR2X1_LOC_416/Y 0.01fF
C478 AND2X1_LOC_788/a_36_24# OR2X1_LOC_533/A 0.00fF
C479 OR2X1_LOC_417/Y OR2X1_LOC_418/Y 0.34fF
C480 OR2X1_LOC_605/B OR2X1_LOC_787/Y 0.01fF
C481 OR2X1_LOC_291/Y OR2X1_LOC_69/Y 0.03fF
C482 OR2X1_LOC_416/Y OR2X1_LOC_44/Y 0.03fF
C483 OR2X1_LOC_611/a_36_216# OR2X1_LOC_6/A 0.03fF
C484 AND2X1_LOC_51/Y OR2X1_LOC_68/a_36_216# 0.00fF
C485 AND2X1_LOC_51/Y OR2X1_LOC_711/A 0.01fF
C486 OR2X1_LOC_427/A AND2X1_LOC_811/Y 0.10fF
C487 AND2X1_LOC_216/A OR2X1_LOC_59/Y 0.16fF
C488 OR2X1_LOC_305/Y AND2X1_LOC_537/Y 0.07fF
C489 OR2X1_LOC_427/A OR2X1_LOC_428/Y 0.01fF
C490 AND2X1_LOC_489/Y AND2X1_LOC_557/a_36_24# 0.00fF
C491 AND2X1_LOC_371/a_8_24# OR2X1_LOC_68/B 0.11fF
C492 AND2X1_LOC_593/Y OR2X1_LOC_95/Y 0.03fF
C493 AND2X1_LOC_18/Y OR2X1_LOC_68/B 0.61fF
C494 OR2X1_LOC_97/A OR2X1_LOC_771/B 0.05fF
C495 OR2X1_LOC_596/A OR2X1_LOC_446/B 0.04fF
C496 OR2X1_LOC_756/B OR2X1_LOC_339/Y 0.01fF
C497 AND2X1_LOC_425/Y OR2X1_LOC_449/B 0.01fF
C498 OR2X1_LOC_3/Y OR2X1_LOC_119/a_8_216# 0.01fF
C499 AND2X1_LOC_706/Y OR2X1_LOC_589/a_36_216# -0.00fF
C500 AND2X1_LOC_196/Y OR2X1_LOC_36/Y 0.01fF
C501 OR2X1_LOC_654/A OR2X1_LOC_476/B 0.01fF
C502 AND2X1_LOC_711/Y OR2X1_LOC_755/A 0.00fF
C503 OR2X1_LOC_814/A OR2X1_LOC_269/B 0.11fF
C504 OR2X1_LOC_742/B OR2X1_LOC_191/a_8_216# 0.01fF
C505 OR2X1_LOC_337/a_36_216# OR2X1_LOC_365/B 0.02fF
C506 AND2X1_LOC_657/Y AND2X1_LOC_657/A 0.01fF
C507 OR2X1_LOC_493/A OR2X1_LOC_786/Y 0.01fF
C508 OR2X1_LOC_833/B OR2X1_LOC_269/Y 0.01fF
C509 AND2X1_LOC_191/B AND2X1_LOC_657/A 0.07fF
C510 OR2X1_LOC_844/Y AND2X1_LOC_42/B 0.05fF
C511 AND2X1_LOC_687/Y OR2X1_LOC_585/A 0.01fF
C512 OR2X1_LOC_173/Y D_INPUT_0 0.03fF
C513 OR2X1_LOC_643/A OR2X1_LOC_532/B 0.03fF
C514 D_INPUT_0 OR2X1_LOC_690/A 0.11fF
C515 INPUT_1 AND2X1_LOC_634/a_8_24# 0.00fF
C516 OR2X1_LOC_95/Y OR2X1_LOC_85/A 0.15fF
C517 OR2X1_LOC_485/A OR2X1_LOC_246/A 0.03fF
C518 AND2X1_LOC_44/Y OR2X1_LOC_844/B 0.01fF
C519 OR2X1_LOC_320/Y AND2X1_LOC_863/A 0.10fF
C520 OR2X1_LOC_524/Y OR2X1_LOC_746/Y 0.03fF
C521 OR2X1_LOC_532/B OR2X1_LOC_778/Y 0.10fF
C522 AND2X1_LOC_397/a_36_24# OR2X1_LOC_68/B 0.01fF
C523 OR2X1_LOC_117/Y OR2X1_LOC_256/A 0.07fF
C524 AND2X1_LOC_571/a_8_24# AND2X1_LOC_571/B 0.19fF
C525 AND2X1_LOC_729/Y OR2X1_LOC_47/Y 0.13fF
C526 AND2X1_LOC_22/Y OR2X1_LOC_605/Y 0.01fF
C527 AND2X1_LOC_319/A AND2X1_LOC_319/a_8_24# 0.03fF
C528 OR2X1_LOC_22/Y AND2X1_LOC_650/a_8_24# 0.03fF
C529 OR2X1_LOC_151/A OR2X1_LOC_535/a_36_216# 0.02fF
C530 VDD OR2X1_LOC_399/Y 0.12fF
C531 OR2X1_LOC_95/Y AND2X1_LOC_602/a_8_24# 0.01fF
C532 OR2X1_LOC_91/Y OR2X1_LOC_437/a_8_216# 0.03fF
C533 OR2X1_LOC_487/a_36_216# OR2X1_LOC_71/Y 0.00fF
C534 AND2X1_LOC_91/B OR2X1_LOC_392/B 0.10fF
C535 OR2X1_LOC_647/A OR2X1_LOC_532/B 0.02fF
C536 OR2X1_LOC_273/Y INPUT_1 0.03fF
C537 OR2X1_LOC_805/A OR2X1_LOC_241/B 0.07fF
C538 AND2X1_LOC_91/B AND2X1_LOC_263/a_8_24# 0.01fF
C539 AND2X1_LOC_784/A OR2X1_LOC_47/Y 0.09fF
C540 OR2X1_LOC_744/A OR2X1_LOC_589/a_8_216# 0.01fF
C541 OR2X1_LOC_188/Y AND2X1_LOC_7/B 0.05fF
C542 OR2X1_LOC_810/A OR2X1_LOC_223/A 0.03fF
C543 OR2X1_LOC_121/B AND2X1_LOC_425/Y 0.00fF
C544 OR2X1_LOC_311/Y AND2X1_LOC_537/Y 0.02fF
C545 OR2X1_LOC_484/Y OR2X1_LOC_437/A 0.01fF
C546 OR2X1_LOC_509/A OR2X1_LOC_560/A 0.04fF
C547 AND2X1_LOC_794/a_8_24# AND2X1_LOC_804/A 0.00fF
C548 OR2X1_LOC_64/Y D_INPUT_0 0.07fF
C549 AND2X1_LOC_537/Y AND2X1_LOC_538/Y 0.11fF
C550 OR2X1_LOC_19/B INPUT_1 0.08fF
C551 OR2X1_LOC_808/A OR2X1_LOC_303/B 0.26fF
C552 OR2X1_LOC_117/Y OR2X1_LOC_67/Y 0.80fF
C553 OR2X1_LOC_375/A AND2X1_LOC_52/Y 0.05fF
C554 OR2X1_LOC_827/Y D_INPUT_1 0.04fF
C555 OR2X1_LOC_47/Y OR2X1_LOC_3/a_8_216# 0.01fF
C556 OR2X1_LOC_646/a_8_216# D_INPUT_1 0.03fF
C557 OR2X1_LOC_157/a_36_216# OR2X1_LOC_70/A 0.00fF
C558 AND2X1_LOC_128/a_36_24# INPUT_1 0.01fF
C559 AND2X1_LOC_231/Y OR2X1_LOC_12/Y 0.01fF
C560 OR2X1_LOC_486/Y OR2X1_LOC_563/A 0.01fF
C561 AND2X1_LOC_364/a_8_24# OR2X1_LOC_12/Y 0.03fF
C562 OR2X1_LOC_31/Y AND2X1_LOC_465/Y 0.01fF
C563 OR2X1_LOC_32/Y OR2X1_LOC_598/A 0.00fF
C564 OR2X1_LOC_286/a_8_216# OR2X1_LOC_286/B 0.08fF
C565 AND2X1_LOC_22/Y AND2X1_LOC_511/a_8_24# 0.02fF
C566 OR2X1_LOC_528/Y AND2X1_LOC_580/a_8_24# 0.01fF
C567 D_INPUT_0 OR2X1_LOC_417/A 0.07fF
C568 OR2X1_LOC_186/Y OR2X1_LOC_355/a_8_216# 0.01fF
C569 AND2X1_LOC_47/Y AND2X1_LOC_600/a_8_24# 0.01fF
C570 OR2X1_LOC_12/Y AND2X1_LOC_770/a_8_24# 0.17fF
C571 AND2X1_LOC_413/a_8_24# OR2X1_LOC_68/B 0.01fF
C572 OR2X1_LOC_105/a_36_216# OR2X1_LOC_579/A 0.01fF
C573 AND2X1_LOC_53/Y AND2X1_LOC_56/a_8_24# 0.21fF
C574 OR2X1_LOC_766/Y AND2X1_LOC_770/a_8_24# 0.01fF
C575 OR2X1_LOC_371/Y OR2X1_LOC_406/A 0.01fF
C576 OR2X1_LOC_589/A OR2X1_LOC_12/Y 0.33fF
C577 INPUT_1 OR2X1_LOC_75/Y 0.26fF
C578 OR2X1_LOC_721/Y OR2X1_LOC_523/a_8_216# 0.29fF
C579 OR2X1_LOC_70/Y AND2X1_LOC_216/A 0.02fF
C580 AND2X1_LOC_534/a_8_24# OR2X1_LOC_151/A 0.02fF
C581 OR2X1_LOC_95/Y OR2X1_LOC_226/Y 0.01fF
C582 OR2X1_LOC_47/Y AND2X1_LOC_639/A 0.08fF
C583 OR2X1_LOC_648/A OR2X1_LOC_390/a_8_216# -0.06fF
C584 VDD OR2X1_LOC_577/Y 0.00fF
C585 OR2X1_LOC_579/B OR2X1_LOC_579/a_8_216# 0.04fF
C586 OR2X1_LOC_51/Y AND2X1_LOC_287/B 0.04fF
C587 OR2X1_LOC_389/A AND2X1_LOC_44/Y 0.03fF
C588 AND2X1_LOC_539/Y INPUT_0 0.01fF
C589 OR2X1_LOC_160/B OR2X1_LOC_706/a_8_216# -0.02fF
C590 OR2X1_LOC_246/Y OR2X1_LOC_437/A 0.02fF
C591 OR2X1_LOC_511/Y OR2X1_LOC_13/B 0.25fF
C592 OR2X1_LOC_51/Y OR2X1_LOC_816/A 0.26fF
C593 OR2X1_LOC_538/A OR2X1_LOC_703/a_8_216# 0.00fF
C594 OR2X1_LOC_378/Y OR2X1_LOC_378/A 0.01fF
C595 OR2X1_LOC_44/Y AND2X1_LOC_592/a_8_24# 0.02fF
C596 OR2X1_LOC_555/A OR2X1_LOC_348/B 0.28fF
C597 AND2X1_LOC_576/Y OR2X1_LOC_437/A 0.07fF
C598 AND2X1_LOC_61/Y AND2X1_LOC_219/A 0.01fF
C599 AND2X1_LOC_835/a_8_24# D_INPUT_1 0.00fF
C600 AND2X1_LOC_561/B OR2X1_LOC_428/A 0.14fF
C601 OR2X1_LOC_190/A OR2X1_LOC_580/B 0.03fF
C602 OR2X1_LOC_471/B AND2X1_LOC_7/B 0.01fF
C603 AND2X1_LOC_22/Y AND2X1_LOC_20/a_8_24# 0.03fF
C604 OR2X1_LOC_248/a_8_216# OR2X1_LOC_13/B 0.01fF
C605 OR2X1_LOC_49/A OR2X1_LOC_56/A 1.94fF
C606 OR2X1_LOC_151/A AND2X1_LOC_110/Y 0.05fF
C607 OR2X1_LOC_329/B OR2X1_LOC_310/a_8_216# 0.12fF
C608 OR2X1_LOC_139/A AND2X1_LOC_65/a_8_24# 0.02fF
C609 OR2X1_LOC_696/A OR2X1_LOC_103/a_36_216# 0.00fF
C610 OR2X1_LOC_62/A OR2X1_LOC_47/Y 3.63fF
C611 AND2X1_LOC_322/a_8_24# AND2X1_LOC_110/Y 0.01fF
C612 AND2X1_LOC_141/a_36_24# OR2X1_LOC_595/A 0.00fF
C613 OR2X1_LOC_851/A OR2X1_LOC_831/B 0.20fF
C614 AND2X1_LOC_561/a_8_24# AND2X1_LOC_572/Y 0.01fF
C615 AND2X1_LOC_294/a_8_24# OR2X1_LOC_13/B 0.02fF
C616 OR2X1_LOC_485/A OR2X1_LOC_599/a_8_216# 0.01fF
C617 AND2X1_LOC_32/a_8_24# AND2X1_LOC_36/Y 0.01fF
C618 AND2X1_LOC_663/A AND2X1_LOC_212/Y 0.10fF
C619 OR2X1_LOC_421/A AND2X1_LOC_596/a_8_24# 0.01fF
C620 OR2X1_LOC_539/A OR2X1_LOC_175/Y 0.02fF
C621 OR2X1_LOC_281/Y OR2X1_LOC_59/Y 0.03fF
C622 AND2X1_LOC_423/a_8_24# AND2X1_LOC_7/B 0.01fF
C623 AND2X1_LOC_794/B AND2X1_LOC_469/B 0.22fF
C624 OR2X1_LOC_787/a_8_216# OR2X1_LOC_787/B 0.05fF
C625 AND2X1_LOC_778/a_36_24# OR2X1_LOC_18/Y 0.00fF
C626 AND2X1_LOC_64/Y OR2X1_LOC_506/A 0.09fF
C627 AND2X1_LOC_30/a_8_24# INPUT_6 0.02fF
C628 OR2X1_LOC_576/A OR2X1_LOC_721/Y 0.07fF
C629 AND2X1_LOC_769/a_36_24# OR2X1_LOC_48/B 0.01fF
C630 OR2X1_LOC_369/Y OR2X1_LOC_309/Y 0.32fF
C631 AND2X1_LOC_555/Y OR2X1_LOC_127/a_36_216# 0.01fF
C632 AND2X1_LOC_857/Y OR2X1_LOC_16/A 4.09fF
C633 OR2X1_LOC_499/a_36_216# OR2X1_LOC_140/B 0.00fF
C634 OR2X1_LOC_47/Y OR2X1_LOC_234/a_36_216# 0.03fF
C635 AND2X1_LOC_769/a_36_24# OR2X1_LOC_18/Y 0.00fF
C636 VDD AND2X1_LOC_657/Y 3.89fF
C637 AND2X1_LOC_64/Y AND2X1_LOC_129/a_8_24# 0.02fF
C638 AND2X1_LOC_738/B OR2X1_LOC_526/Y 0.06fF
C639 OR2X1_LOC_598/Y INPUT_0 0.03fF
C640 AND2X1_LOC_654/B OR2X1_LOC_12/Y 0.32fF
C641 AND2X1_LOC_191/B VDD 0.58fF
C642 AND2X1_LOC_707/a_8_24# OR2X1_LOC_51/Y 0.01fF
C643 AND2X1_LOC_734/Y AND2X1_LOC_476/Y 0.07fF
C644 VDD AND2X1_LOC_469/B 0.27fF
C645 OR2X1_LOC_161/A OR2X1_LOC_161/a_8_216# 0.01fF
C646 OR2X1_LOC_155/A OR2X1_LOC_319/Y 0.13fF
C647 OR2X1_LOC_405/Y AND2X1_LOC_7/B 0.06fF
C648 OR2X1_LOC_6/B OR2X1_LOC_756/B 0.02fF
C649 OR2X1_LOC_641/Y AND2X1_LOC_92/Y 0.01fF
C650 OR2X1_LOC_188/Y OR2X1_LOC_805/A 0.03fF
C651 AND2X1_LOC_326/B INPUT_0 0.03fF
C652 OR2X1_LOC_114/B AND2X1_LOC_71/a_8_24# 0.01fF
C653 OR2X1_LOC_651/A AND2X1_LOC_31/Y 0.06fF
C654 AND2X1_LOC_59/Y AND2X1_LOC_60/a_8_24# 0.00fF
C655 OR2X1_LOC_139/A OR2X1_LOC_130/A 0.07fF
C656 OR2X1_LOC_633/Y OR2X1_LOC_633/A 0.00fF
C657 OR2X1_LOC_375/A OR2X1_LOC_576/A 0.03fF
C658 OR2X1_LOC_680/A OR2X1_LOC_816/A 0.03fF
C659 OR2X1_LOC_207/B AND2X1_LOC_43/B 0.03fF
C660 OR2X1_LOC_36/Y OR2X1_LOC_321/a_8_216# 0.02fF
C661 OR2X1_LOC_87/A OR2X1_LOC_352/a_8_216# 0.01fF
C662 OR2X1_LOC_329/B AND2X1_LOC_434/Y 0.07fF
C663 OR2X1_LOC_121/B OR2X1_LOC_723/B 0.00fF
C664 OR2X1_LOC_158/A OR2X1_LOC_427/A 0.37fF
C665 AND2X1_LOC_663/B AND2X1_LOC_791/a_8_24# 0.01fF
C666 OR2X1_LOC_310/Y OR2X1_LOC_56/A 0.03fF
C667 AND2X1_LOC_704/a_36_24# OR2X1_LOC_427/A 0.00fF
C668 AND2X1_LOC_320/a_8_24# OR2X1_LOC_324/B 0.01fF
C669 OR2X1_LOC_624/A AND2X1_LOC_65/A 0.05fF
C670 OR2X1_LOC_109/a_8_216# AND2X1_LOC_476/Y 0.03fF
C671 VDD OR2X1_LOC_833/a_8_216# 0.21fF
C672 AND2X1_LOC_535/Y OR2X1_LOC_761/Y 0.01fF
C673 OR2X1_LOC_677/Y AND2X1_LOC_657/Y 0.28fF
C674 AND2X1_LOC_32/a_36_24# OR2X1_LOC_34/A 0.00fF
C675 OR2X1_LOC_660/Y OR2X1_LOC_662/a_8_216# 0.01fF
C676 AND2X1_LOC_22/Y OR2X1_LOC_845/a_8_216# 0.04fF
C677 AND2X1_LOC_537/a_8_24# OR2X1_LOC_92/Y 0.03fF
C678 AND2X1_LOC_29/a_8_24# AND2X1_LOC_44/Y 0.01fF
C679 OR2X1_LOC_244/A OR2X1_LOC_140/Y 0.20fF
C680 OR2X1_LOC_51/Y OR2X1_LOC_251/a_8_216# 0.04fF
C681 AND2X1_LOC_231/Y AND2X1_LOC_650/Y 0.26fF
C682 OR2X1_LOC_40/Y OR2X1_LOC_291/a_8_216# 0.01fF
C683 OR2X1_LOC_687/Y OR2X1_LOC_161/B 0.03fF
C684 AND2X1_LOC_41/A OR2X1_LOC_78/B 0.14fF
C685 OR2X1_LOC_294/a_8_216# OR2X1_LOC_78/A 0.01fF
C686 AND2X1_LOC_304/a_8_24# OR2X1_LOC_78/A 0.01fF
C687 OR2X1_LOC_696/A OR2X1_LOC_481/A 0.02fF
C688 OR2X1_LOC_49/A AND2X1_LOC_56/B 0.07fF
C689 OR2X1_LOC_31/Y OR2X1_LOC_589/a_8_216# 0.01fF
C690 OR2X1_LOC_122/Y AND2X1_LOC_474/A 0.01fF
C691 AND2X1_LOC_266/Y OR2X1_LOC_595/A 0.27fF
C692 OR2X1_LOC_648/A AND2X1_LOC_58/a_8_24# 0.02fF
C693 OR2X1_LOC_744/A AND2X1_LOC_141/A 0.00fF
C694 OR2X1_LOC_821/Y OR2X1_LOC_85/A 0.06fF
C695 AND2X1_LOC_852/Y AND2X1_LOC_219/A 0.46fF
C696 AND2X1_LOC_160/a_36_24# OR2X1_LOC_744/A 0.00fF
C697 OR2X1_LOC_49/A AND2X1_LOC_8/Y 0.62fF
C698 OR2X1_LOC_528/Y OR2X1_LOC_252/Y 0.12fF
C699 OR2X1_LOC_151/A OR2X1_LOC_664/Y 0.03fF
C700 AND2X1_LOC_562/B OR2X1_LOC_698/a_8_216# 0.00fF
C701 OR2X1_LOC_43/A OR2X1_LOC_12/Y 0.41fF
C702 AND2X1_LOC_447/Y OR2X1_LOC_48/B 0.03fF
C703 AND2X1_LOC_40/Y INPUT_0 0.07fF
C704 AND2X1_LOC_358/Y AND2X1_LOC_211/B 0.04fF
C705 OR2X1_LOC_780/B OR2X1_LOC_712/B 0.00fF
C706 OR2X1_LOC_675/Y OR2X1_LOC_736/a_8_216# 0.14fF
C707 AND2X1_LOC_56/B OR2X1_LOC_596/A 0.02fF
C708 AND2X1_LOC_22/Y AND2X1_LOC_43/a_36_24# 0.00fF
C709 OR2X1_LOC_490/a_8_216# AND2X1_LOC_101/B 0.47fF
C710 OR2X1_LOC_56/A AND2X1_LOC_805/Y 0.00fF
C711 OR2X1_LOC_811/A OR2X1_LOC_78/A 0.03fF
C712 AND2X1_LOC_41/A OR2X1_LOC_721/Y 0.05fF
C713 AND2X1_LOC_352/B AND2X1_LOC_662/B 0.82fF
C714 OR2X1_LOC_45/B AND2X1_LOC_640/Y 3.61fF
C715 OR2X1_LOC_335/A OR2X1_LOC_121/B 0.00fF
C716 OR2X1_LOC_51/Y AND2X1_LOC_843/a_8_24# 0.01fF
C717 AND2X1_LOC_539/Y OR2X1_LOC_64/Y 0.02fF
C718 AND2X1_LOC_528/a_36_24# AND2X1_LOC_44/Y 0.01fF
C719 OR2X1_LOC_193/A AND2X1_LOC_7/B 0.03fF
C720 OR2X1_LOC_728/B OR2X1_LOC_715/a_8_216# 0.47fF
C721 OR2X1_LOC_161/A OR2X1_LOC_360/a_8_216# 0.01fF
C722 OR2X1_LOC_798/Y OR2X1_LOC_802/a_8_216# 0.01fF
C723 AND2X1_LOC_486/Y AND2X1_LOC_850/A 0.23fF
C724 AND2X1_LOC_70/Y OR2X1_LOC_639/B 0.01fF
C725 OR2X1_LOC_421/A OR2X1_LOC_36/Y 0.05fF
C726 OR2X1_LOC_669/A AND2X1_LOC_860/A 0.01fF
C727 AND2X1_LOC_191/B OR2X1_LOC_616/Y 0.00fF
C728 AND2X1_LOC_533/a_8_24# OR2X1_LOC_78/A 0.06fF
C729 OR2X1_LOC_508/A OR2X1_LOC_721/Y 0.45fF
C730 OR2X1_LOC_45/B OR2X1_LOC_681/Y 0.06fF
C731 OR2X1_LOC_696/A OR2X1_LOC_71/Y 0.04fF
C732 OR2X1_LOC_402/Y OR2X1_LOC_78/a_8_216# 0.01fF
C733 OR2X1_LOC_597/A OR2X1_LOC_599/A 0.02fF
C734 OR2X1_LOC_662/A OR2X1_LOC_78/B 0.01fF
C735 OR2X1_LOC_323/A INPUT_1 0.03fF
C736 OR2X1_LOC_847/A AND2X1_LOC_820/B 0.02fF
C737 OR2X1_LOC_814/A OR2X1_LOC_718/a_36_216# 0.01fF
C738 OR2X1_LOC_639/A AND2X1_LOC_44/Y 0.02fF
C739 OR2X1_LOC_517/A OR2X1_LOC_278/Y 0.00fF
C740 AND2X1_LOC_863/a_8_24# AND2X1_LOC_654/Y 0.04fF
C741 AND2X1_LOC_212/Y AND2X1_LOC_212/B 0.02fF
C742 OR2X1_LOC_610/a_8_216# OR2X1_LOC_502/A 0.01fF
C743 OR2X1_LOC_303/B OR2X1_LOC_374/Y 0.57fF
C744 OR2X1_LOC_352/A AND2X1_LOC_95/Y 0.03fF
C745 OR2X1_LOC_103/Y OR2X1_LOC_427/A 0.01fF
C746 AND2X1_LOC_436/B AND2X1_LOC_436/a_8_24# 0.06fF
C747 VDD AND2X1_LOC_158/a_8_24# -0.00fF
C748 OR2X1_LOC_580/A OR2X1_LOC_493/Y 0.03fF
C749 OR2X1_LOC_45/B OR2X1_LOC_416/Y 0.06fF
C750 OR2X1_LOC_60/a_8_216# OR2X1_LOC_12/Y 0.01fF
C751 OR2X1_LOC_9/Y AND2X1_LOC_37/a_8_24# 0.00fF
C752 OR2X1_LOC_589/A OR2X1_LOC_272/Y 0.02fF
C753 OR2X1_LOC_59/Y AND2X1_LOC_286/Y 0.17fF
C754 AND2X1_LOC_240/Y AND2X1_LOC_243/Y 0.01fF
C755 AND2X1_LOC_538/a_36_24# OR2X1_LOC_485/A 0.00fF
C756 AND2X1_LOC_95/Y OR2X1_LOC_434/a_36_216# 0.00fF
C757 AND2X1_LOC_41/A OR2X1_LOC_375/A 1.98fF
C758 VDD AND2X1_LOC_638/a_8_24# -0.00fF
C759 AND2X1_LOC_658/B OR2X1_LOC_52/B 0.09fF
C760 AND2X1_LOC_91/B OR2X1_LOC_532/B 0.53fF
C761 OR2X1_LOC_139/A OR2X1_LOC_62/B 0.00fF
C762 OR2X1_LOC_92/Y OR2X1_LOC_71/a_8_216# 0.01fF
C763 OR2X1_LOC_154/A OR2X1_LOC_235/B -0.03fF
C764 OR2X1_LOC_70/Y OR2X1_LOC_584/Y 0.03fF
C765 AND2X1_LOC_794/B OR2X1_LOC_417/a_36_216# 0.01fF
C766 AND2X1_LOC_703/a_8_24# AND2X1_LOC_841/B 0.06fF
C767 OR2X1_LOC_649/a_8_216# AND2X1_LOC_44/Y 0.03fF
C768 AND2X1_LOC_22/Y OR2X1_LOC_335/B 0.05fF
C769 D_INPUT_7 VDD 0.36fF
C770 AND2X1_LOC_510/a_8_24# AND2X1_LOC_580/A 0.03fF
C771 D_INPUT_0 AND2X1_LOC_7/B 0.04fF
C772 AND2X1_LOC_191/B OR2X1_LOC_251/Y 0.03fF
C773 OR2X1_LOC_756/B OR2X1_LOC_579/B 0.00fF
C774 OR2X1_LOC_64/Y AND2X1_LOC_771/B 0.03fF
C775 AND2X1_LOC_642/a_8_24# AND2X1_LOC_649/a_8_24# 0.23fF
C776 AND2X1_LOC_642/a_36_24# AND2X1_LOC_642/Y 0.00fF
C777 OR2X1_LOC_147/B OR2X1_LOC_739/A 0.10fF
C778 OR2X1_LOC_643/A OR2X1_LOC_624/Y 0.03fF
C779 OR2X1_LOC_702/A VDD 0.23fF
C780 AND2X1_LOC_510/A AND2X1_LOC_474/Y 0.89fF
C781 AND2X1_LOC_570/Y AND2X1_LOC_456/Y 0.34fF
C782 OR2X1_LOC_502/A OR2X1_LOC_510/Y 0.01fF
C783 OR2X1_LOC_508/A OR2X1_LOC_375/A 0.00fF
C784 OR2X1_LOC_235/B OR2X1_LOC_267/A 0.03fF
C785 OR2X1_LOC_604/A OR2X1_LOC_279/Y 0.10fF
C786 AND2X1_LOC_259/Y OR2X1_LOC_56/A 0.00fF
C787 OR2X1_LOC_848/B OR2X1_LOC_392/A 0.71fF
C788 AND2X1_LOC_337/B AND2X1_LOC_352/B 0.15fF
C789 AND2X1_LOC_456/B OR2X1_LOC_36/Y 0.16fF
C790 OR2X1_LOC_333/B AND2X1_LOC_70/Y 0.06fF
C791 OR2X1_LOC_109/Y OR2X1_LOC_48/B 0.02fF
C792 OR2X1_LOC_696/A D_INPUT_1 0.95fF
C793 OR2X1_LOC_784/a_8_216# OR2X1_LOC_78/A 0.01fF
C794 AND2X1_LOC_570/Y OR2X1_LOC_74/A 0.03fF
C795 AND2X1_LOC_64/Y OR2X1_LOC_227/Y 0.08fF
C796 AND2X1_LOC_666/a_8_24# AND2X1_LOC_18/Y 0.03fF
C797 OR2X1_LOC_311/Y OR2X1_LOC_13/Y 1.09fF
C798 OR2X1_LOC_317/A OR2X1_LOC_739/A 0.01fF
C799 OR2X1_LOC_808/a_36_216# OR2X1_LOC_375/A 0.00fF
C800 OR2X1_LOC_840/A OR2X1_LOC_468/Y 0.03fF
C801 OR2X1_LOC_109/Y OR2X1_LOC_18/Y 0.01fF
C802 OR2X1_LOC_280/Y OR2X1_LOC_59/Y 0.03fF
C803 OR2X1_LOC_678/Y OR2X1_LOC_155/A 0.01fF
C804 AND2X1_LOC_559/a_36_24# OR2X1_LOC_517/A 0.00fF
C805 OR2X1_LOC_848/A OR2X1_LOC_772/B 0.03fF
C806 OR2X1_LOC_448/Y OR2X1_LOC_784/Y 0.18fF
C807 OR2X1_LOC_324/a_8_216# AND2X1_LOC_56/B 0.03fF
C808 AND2X1_LOC_64/Y D_INPUT_1 0.05fF
C809 AND2X1_LOC_47/Y OR2X1_LOC_342/A 0.01fF
C810 AND2X1_LOC_304/a_8_24# OR2X1_LOC_155/A 0.06fF
C811 AND2X1_LOC_654/B AND2X1_LOC_650/Y 0.00fF
C812 AND2X1_LOC_191/B AND2X1_LOC_624/a_8_24# 0.01fF
C813 OR2X1_LOC_744/A AND2X1_LOC_651/B 0.00fF
C814 AND2X1_LOC_160/a_8_24# OR2X1_LOC_7/A 0.05fF
C815 AND2X1_LOC_621/Y OR2X1_LOC_39/A 0.15fF
C816 AND2X1_LOC_326/B OR2X1_LOC_64/Y 0.03fF
C817 OR2X1_LOC_451/a_36_216# AND2X1_LOC_425/Y 0.00fF
C818 AND2X1_LOC_562/B OR2X1_LOC_7/A 0.03fF
C819 VDD OR2X1_LOC_476/B 1.07fF
C820 OR2X1_LOC_502/A OR2X1_LOC_810/A 0.07fF
C821 OR2X1_LOC_160/B OR2X1_LOC_750/A 0.03fF
C822 OR2X1_LOC_32/B OR2X1_LOC_69/A 0.03fF
C823 OR2X1_LOC_307/a_8_216# OR2X1_LOC_502/A 0.03fF
C824 AND2X1_LOC_583/a_8_24# OR2X1_LOC_636/A 0.09fF
C825 AND2X1_LOC_40/Y OR2X1_LOC_592/a_36_216# 0.00fF
C826 OR2X1_LOC_485/A AND2X1_LOC_842/a_36_24# 0.00fF
C827 OR2X1_LOC_604/A OR2X1_LOC_77/a_8_216# 0.02fF
C828 AND2X1_LOC_39/a_8_24# AND2X1_LOC_3/Y 0.01fF
C829 OR2X1_LOC_603/a_8_216# AND2X1_LOC_453/Y 0.47fF
C830 AND2X1_LOC_135/a_8_24# OR2X1_LOC_78/B 0.04fF
C831 VDD OR2X1_LOC_650/Y 0.39fF
C832 AND2X1_LOC_124/a_8_24# OR2X1_LOC_67/A 0.02fF
C833 OR2X1_LOC_452/a_8_216# AND2X1_LOC_425/Y 0.01fF
C834 OR2X1_LOC_680/A AND2X1_LOC_807/Y 0.10fF
C835 AND2X1_LOC_64/Y OR2X1_LOC_356/a_36_216# 0.03fF
C836 OR2X1_LOC_489/B OR2X1_LOC_848/A 0.01fF
C837 OR2X1_LOC_51/Y AND2X1_LOC_727/A 0.02fF
C838 OR2X1_LOC_71/Y OR2X1_LOC_131/a_36_216# 0.00fF
C839 AND2X1_LOC_165/a_8_24# OR2X1_LOC_66/A 0.01fF
C840 AND2X1_LOC_500/Y AND2X1_LOC_574/A 0.00fF
C841 OR2X1_LOC_203/a_8_216# OR2X1_LOC_203/Y 0.00fF
C842 OR2X1_LOC_64/Y AND2X1_LOC_471/Y 0.05fF
C843 OR2X1_LOC_121/Y OR2X1_LOC_276/a_36_216# 0.01fF
C844 OR2X1_LOC_295/a_36_216# OR2X1_LOC_59/Y 0.03fF
C845 OR2X1_LOC_807/a_8_216# OR2X1_LOC_811/A 0.14fF
C846 OR2X1_LOC_694/a_8_216# OR2X1_LOC_43/A 0.06fF
C847 OR2X1_LOC_161/B OR2X1_LOC_364/a_36_216# 0.00fF
C848 AND2X1_LOC_737/Y AND2X1_LOC_711/Y 0.04fF
C849 OR2X1_LOC_836/A AND2X1_LOC_824/a_36_24# 0.00fF
C850 AND2X1_LOC_97/a_8_24# OR2X1_LOC_89/A 0.12fF
C851 OR2X1_LOC_22/Y OR2X1_LOC_59/Y 0.21fF
C852 AND2X1_LOC_94/Y AND2X1_LOC_825/a_8_24# 0.09fF
C853 AND2X1_LOC_72/B AND2X1_LOC_248/a_8_24# 0.01fF
C854 AND2X1_LOC_82/Y D_INPUT_1 0.03fF
C855 OR2X1_LOC_154/A AND2X1_LOC_393/a_8_24# 0.14fF
C856 OR2X1_LOC_185/Y OR2X1_LOC_194/Y 0.52fF
C857 OR2X1_LOC_697/Y AND2X1_LOC_708/a_8_24# 0.12fF
C858 OR2X1_LOC_697/a_36_216# AND2X1_LOC_712/B 0.00fF
C859 VDD OR2X1_LOC_111/Y 0.25fF
C860 OR2X1_LOC_632/A OR2X1_LOC_574/A 0.04fF
C861 AND2X1_LOC_326/B OR2X1_LOC_417/A 0.15fF
C862 AND2X1_LOC_17/Y OR2X1_LOC_639/B 0.16fF
C863 AND2X1_LOC_44/Y OR2X1_LOC_493/Y 0.01fF
C864 OR2X1_LOC_615/a_8_216# OR2X1_LOC_92/Y 0.01fF
C865 OR2X1_LOC_185/Y OR2X1_LOC_114/Y 0.05fF
C866 OR2X1_LOC_6/A OR2X1_LOC_44/Y 1.81fF
C867 OR2X1_LOC_520/Y OR2X1_LOC_99/Y 0.02fF
C868 OR2X1_LOC_715/B OR2X1_LOC_223/A 0.05fF
C869 OR2X1_LOC_375/A OR2X1_LOC_217/a_36_216# 0.00fF
C870 OR2X1_LOC_246/Y OR2X1_LOC_753/A 0.08fF
C871 AND2X1_LOC_580/B OR2X1_LOC_613/Y 0.04fF
C872 OR2X1_LOC_19/B OR2X1_LOC_517/A 0.05fF
C873 AND2X1_LOC_3/Y AND2X1_LOC_43/B 0.35fF
C874 OR2X1_LOC_369/Y OR2X1_LOC_31/Y -0.00fF
C875 OR2X1_LOC_562/A OR2X1_LOC_344/a_8_216# 0.01fF
C876 AND2X1_LOC_31/Y OR2X1_LOC_338/A 0.02fF
C877 OR2X1_LOC_51/Y OR2X1_LOC_95/Y 3.67fF
C878 OR2X1_LOC_223/A OR2X1_LOC_543/A 0.01fF
C879 AND2X1_LOC_8/Y OR2X1_LOC_87/B 0.11fF
C880 AND2X1_LOC_656/Y AND2X1_LOC_218/Y 0.01fF
C881 AND2X1_LOC_729/B OR2X1_LOC_48/B 0.03fF
C882 AND2X1_LOC_59/Y OR2X1_LOC_557/A 0.02fF
C883 AND2X1_LOC_218/a_36_24# AND2X1_LOC_660/A 0.00fF
C884 OR2X1_LOC_64/Y AND2X1_LOC_840/A 0.03fF
C885 INPUT_0 AND2X1_LOC_826/a_8_24# 0.05fF
C886 OR2X1_LOC_62/B OR2X1_LOC_244/a_8_216# 0.01fF
C887 AND2X1_LOC_810/Y OR2X1_LOC_56/A 0.01fF
C888 OR2X1_LOC_26/Y OR2X1_LOC_588/Y 0.04fF
C889 OR2X1_LOC_405/A AND2X1_LOC_674/a_8_24# 0.00fF
C890 AND2X1_LOC_86/a_8_24# D_INPUT_1 0.05fF
C891 AND2X1_LOC_512/a_8_24# OR2X1_LOC_36/Y 0.03fF
C892 VDD OR2X1_LOC_146/Y 0.08fF
C893 OR2X1_LOC_218/Y AND2X1_LOC_92/Y 0.02fF
C894 OR2X1_LOC_18/Y AND2X1_LOC_729/B 0.03fF
C895 OR2X1_LOC_252/Y AND2X1_LOC_483/a_8_24# 0.09fF
C896 OR2X1_LOC_600/A AND2X1_LOC_837/a_8_24# 0.01fF
C897 AND2X1_LOC_683/a_8_24# OR2X1_LOC_87/A 0.02fF
C898 AND2X1_LOC_803/B AND2X1_LOC_803/a_8_24# 0.11fF
C899 AND2X1_LOC_95/Y OR2X1_LOC_479/a_8_216# 0.04fF
C900 OR2X1_LOC_36/Y AND2X1_LOC_717/B 0.04fF
C901 OR2X1_LOC_703/A OR2X1_LOC_443/a_8_216# 0.04fF
C902 OR2X1_LOC_8/Y OR2X1_LOC_47/Y 0.06fF
C903 OR2X1_LOC_751/Y INPUT_1 0.01fF
C904 OR2X1_LOC_154/A OR2X1_LOC_844/a_8_216# -0.02fF
C905 OR2X1_LOC_269/B OR2X1_LOC_383/a_8_216# 0.01fF
C906 OR2X1_LOC_319/B D_INPUT_0 0.06fF
C907 OR2X1_LOC_231/B OR2X1_LOC_641/B 0.01fF
C908 OR2X1_LOC_756/B AND2X1_LOC_47/Y 0.17fF
C909 OR2X1_LOC_329/B AND2X1_LOC_851/B 0.00fF
C910 OR2X1_LOC_485/A OR2X1_LOC_497/Y 0.03fF
C911 AND2X1_LOC_59/Y OR2X1_LOC_675/A 0.00fF
C912 AND2X1_LOC_56/B OR2X1_LOC_33/B 0.22fF
C913 AND2X1_LOC_95/Y OR2X1_LOC_34/B 0.01fF
C914 AND2X1_LOC_85/a_8_24# AND2X1_LOC_8/Y 0.01fF
C915 OR2X1_LOC_45/B OR2X1_LOC_80/A 0.05fF
C916 AND2X1_LOC_387/B OR2X1_LOC_269/B 0.02fF
C917 OR2X1_LOC_87/A AND2X1_LOC_69/Y 0.03fF
C918 OR2X1_LOC_186/Y AND2X1_LOC_31/Y 0.11fF
C919 OR2X1_LOC_655/a_8_216# AND2X1_LOC_48/A 0.01fF
C920 OR2X1_LOC_185/Y OR2X1_LOC_201/Y 0.08fF
C921 OR2X1_LOC_84/B OR2X1_LOC_633/B 0.00fF
C922 OR2X1_LOC_318/Y D_INPUT_0 0.20fF
C923 OR2X1_LOC_272/Y OR2X1_LOC_43/A 0.03fF
C924 AND2X1_LOC_95/Y AND2X1_LOC_107/a_8_24# 0.01fF
C925 OR2X1_LOC_256/Y AND2X1_LOC_866/A 0.03fF
C926 OR2X1_LOC_357/a_36_216# OR2X1_LOC_578/B 0.02fF
C927 OR2X1_LOC_404/Y OR2X1_LOC_720/A 0.01fF
C928 OR2X1_LOC_160/A OR2X1_LOC_227/a_36_216# 0.00fF
C929 AND2X1_LOC_191/B AND2X1_LOC_624/B 0.03fF
C930 AND2X1_LOC_717/B AND2X1_LOC_493/a_36_24# 0.00fF
C931 OR2X1_LOC_680/A AND2X1_LOC_727/A 0.03fF
C932 AND2X1_LOC_143/a_8_24# OR2X1_LOC_62/A 0.09fF
C933 OR2X1_LOC_757/A AND2X1_LOC_792/Y 0.07fF
C934 OR2X1_LOC_185/Y OR2X1_LOC_844/Y 0.05fF
C935 AND2X1_LOC_838/Y OR2X1_LOC_46/A 0.02fF
C936 AND2X1_LOC_211/B AND2X1_LOC_650/a_8_24# 0.01fF
C937 OR2X1_LOC_814/A OR2X1_LOC_539/Y 0.13fF
C938 OR2X1_LOC_70/Y AND2X1_LOC_356/B 0.03fF
C939 OR2X1_LOC_486/Y OR2X1_LOC_365/a_36_216# 0.02fF
C940 OR2X1_LOC_17/Y AND2X1_LOC_639/a_8_24# 0.01fF
C941 D_INPUT_0 OR2X1_LOC_805/A 0.03fF
C942 AND2X1_LOC_554/B AND2X1_LOC_140/a_8_24# 0.01fF
C943 OR2X1_LOC_175/Y OR2X1_LOC_771/B 0.12fF
C944 AND2X1_LOC_7/B OR2X1_LOC_339/A 0.12fF
C945 OR2X1_LOC_3/Y AND2X1_LOC_196/a_8_24# 0.06fF
C946 AND2X1_LOC_497/a_8_24# OR2X1_LOC_632/Y -0.00fF
C947 OR2X1_LOC_16/A OR2X1_LOC_437/A 0.07fF
C948 AND2X1_LOC_512/Y OR2X1_LOC_599/Y 0.13fF
C949 OR2X1_LOC_433/a_8_216# OR2X1_LOC_22/Y 0.01fF
C950 OR2X1_LOC_66/A OR2X1_LOC_228/Y 0.03fF
C951 OR2X1_LOC_532/a_8_216# AND2X1_LOC_44/Y 0.02fF
C952 VDD OR2X1_LOC_588/a_8_216# 0.21fF
C953 OR2X1_LOC_841/A OR2X1_LOC_228/Y 0.01fF
C954 OR2X1_LOC_287/B AND2X1_LOC_816/a_8_24# 0.01fF
C955 OR2X1_LOC_836/A D_INPUT_0 0.01fF
C956 OR2X1_LOC_485/A AND2X1_LOC_844/a_8_24# 0.10fF
C957 OR2X1_LOC_161/B OR2X1_LOC_181/Y 0.02fF
C958 OR2X1_LOC_743/Y AND2X1_LOC_780/a_8_24# 0.23fF
C959 AND2X1_LOC_8/Y OR2X1_LOC_649/a_36_216# 0.03fF
C960 OR2X1_LOC_542/a_8_216# OR2X1_LOC_367/B 0.31fF
C961 OR2X1_LOC_97/A OR2X1_LOC_593/B 0.02fF
C962 OR2X1_LOC_756/B OR2X1_LOC_598/A 0.07fF
C963 VDD AND2X1_LOC_206/Y 0.01fF
C964 OR2X1_LOC_680/A OR2X1_LOC_95/Y 0.37fF
C965 AND2X1_LOC_512/Y OR2X1_LOC_331/a_8_216# 0.03fF
C966 OR2X1_LOC_80/a_36_216# OR2X1_LOC_6/A 0.03fF
C967 OR2X1_LOC_43/A AND2X1_LOC_801/B 0.00fF
C968 OR2X1_LOC_428/A OR2X1_LOC_268/Y 0.06fF
C969 OR2X1_LOC_287/B OR2X1_LOC_859/A 0.02fF
C970 OR2X1_LOC_22/A OR2X1_LOC_21/a_8_216# -0.00fF
C971 OR2X1_LOC_481/A AND2X1_LOC_663/B 0.00fF
C972 OR2X1_LOC_151/A OR2X1_LOC_550/B 0.07fF
C973 OR2X1_LOC_428/A OR2X1_LOC_183/Y 0.02fF
C974 OR2X1_LOC_837/B AND2X1_LOC_462/B 0.65fF
C975 OR2X1_LOC_436/Y OR2X1_LOC_798/a_36_216# 0.00fF
C976 OR2X1_LOC_222/a_8_216# OR2X1_LOC_222/A 0.04fF
C977 OR2X1_LOC_380/A OR2X1_LOC_64/a_36_216# 0.00fF
C978 AND2X1_LOC_114/a_8_24# AND2X1_LOC_114/Y 0.00fF
C979 OR2X1_LOC_744/A AND2X1_LOC_793/B 0.60fF
C980 OR2X1_LOC_154/A OR2X1_LOC_276/B 0.10fF
C981 VDD OR2X1_LOC_164/a_8_216# 0.21fF
C982 OR2X1_LOC_185/Y OR2X1_LOC_201/a_8_216# 0.01fF
C983 OR2X1_LOC_47/Y OR2X1_LOC_67/A 0.02fF
C984 D_INPUT_7 AND2X1_LOC_25/a_8_24# 0.09fF
C985 OR2X1_LOC_235/B OR2X1_LOC_560/A 0.02fF
C986 OR2X1_LOC_744/A OR2X1_LOC_533/A 0.01fF
C987 OR2X1_LOC_108/Y OR2X1_LOC_437/A 1.05fF
C988 OR2X1_LOC_506/B OR2X1_LOC_87/A 0.03fF
C989 OR2X1_LOC_375/A OR2X1_LOC_207/a_8_216# 0.01fF
C990 OR2X1_LOC_70/Y OR2X1_LOC_22/Y 2.22fF
C991 OR2X1_LOC_696/A OR2X1_LOC_585/a_8_216# 0.02fF
C992 AND2X1_LOC_324/a_8_24# OR2X1_LOC_46/A 0.05fF
C993 OR2X1_LOC_32/Y AND2X1_LOC_462/Y 0.00fF
C994 AND2X1_LOC_159/a_36_24# AND2X1_LOC_47/Y 0.00fF
C995 OR2X1_LOC_190/A OR2X1_LOC_367/a_8_216# 0.05fF
C996 AND2X1_LOC_51/Y OR2X1_LOC_846/A 0.01fF
C997 OR2X1_LOC_813/A OR2X1_LOC_74/A 0.00fF
C998 OR2X1_LOC_502/A AND2X1_LOC_609/a_36_24# 0.00fF
C999 AND2X1_LOC_798/A AND2X1_LOC_354/B 0.00fF
C1000 OR2X1_LOC_64/Y AND2X1_LOC_687/A 0.03fF
C1001 OR2X1_LOC_696/A AND2X1_LOC_714/a_8_24# 0.03fF
C1002 OR2X1_LOC_476/B OR2X1_LOC_476/a_36_216# 0.03fF
C1003 OR2X1_LOC_31/Y OR2X1_LOC_47/a_8_216# 0.01fF
C1004 OR2X1_LOC_47/Y AND2X1_LOC_374/Y 0.01fF
C1005 AND2X1_LOC_514/Y OR2X1_LOC_22/Y 0.07fF
C1006 OR2X1_LOC_31/Y AND2X1_LOC_651/B 0.01fF
C1007 OR2X1_LOC_47/Y OR2X1_LOC_52/B 0.22fF
C1008 AND2X1_LOC_663/B OR2X1_LOC_71/Y 0.01fF
C1009 OR2X1_LOC_78/A OR2X1_LOC_777/B 0.11fF
C1010 OR2X1_LOC_364/A OR2X1_LOC_544/a_8_216# 0.02fF
C1011 AND2X1_LOC_538/a_8_24# OR2X1_LOC_22/Y 0.01fF
C1012 AND2X1_LOC_564/B OR2X1_LOC_373/Y 0.00fF
C1013 OR2X1_LOC_548/A OR2X1_LOC_415/Y 0.01fF
C1014 AND2X1_LOC_489/Y OR2X1_LOC_47/Y 0.02fF
C1015 AND2X1_LOC_12/Y OR2X1_LOC_641/B 0.07fF
C1016 AND2X1_LOC_476/A OR2X1_LOC_27/a_8_216# 0.04fF
C1017 OR2X1_LOC_648/A OR2X1_LOC_539/B 0.03fF
C1018 OR2X1_LOC_276/B OR2X1_LOC_778/A 0.00fF
C1019 AND2X1_LOC_157/a_8_24# AND2X1_LOC_430/B 0.00fF
C1020 OR2X1_LOC_231/a_36_216# AND2X1_LOC_31/Y 0.00fF
C1021 AND2X1_LOC_47/a_8_24# AND2X1_LOC_31/Y 0.01fF
C1022 OR2X1_LOC_458/B OR2X1_LOC_777/B 0.03fF
C1023 AND2X1_LOC_712/a_36_24# OR2X1_LOC_428/A 0.00fF
C1024 AND2X1_LOC_554/B AND2X1_LOC_721/A 0.02fF
C1025 AND2X1_LOC_520/a_8_24# AND2X1_LOC_339/B 0.19fF
C1026 OR2X1_LOC_161/A OR2X1_LOC_348/B 0.03fF
C1027 OR2X1_LOC_269/B OR2X1_LOC_318/B 0.03fF
C1028 OR2X1_LOC_91/Y AND2X1_LOC_563/Y 0.03fF
C1029 OR2X1_LOC_3/a_8_216# OR2X1_LOC_3/B 0.03fF
C1030 OR2X1_LOC_160/A OR2X1_LOC_80/A 0.06fF
C1031 AND2X1_LOC_727/a_8_24# AND2X1_LOC_727/B 0.11fF
C1032 AND2X1_LOC_81/B AND2X1_LOC_31/Y 0.03fF
C1033 OR2X1_LOC_12/Y AND2X1_LOC_771/a_8_24# 0.01fF
C1034 OR2X1_LOC_696/A OR2X1_LOC_426/B 0.17fF
C1035 AND2X1_LOC_339/Y AND2X1_LOC_339/B 0.21fF
C1036 AND2X1_LOC_717/B OR2X1_LOC_419/Y 0.05fF
C1037 OR2X1_LOC_448/B OR2X1_LOC_777/B 0.04fF
C1038 OR2X1_LOC_323/A AND2X1_LOC_325/a_8_24# 0.09fF
C1039 AND2X1_LOC_7/B OR2X1_LOC_515/A 0.03fF
C1040 OR2X1_LOC_479/Y OR2X1_LOC_804/A 0.02fF
C1041 AND2X1_LOC_168/Y OR2X1_LOC_437/A 0.08fF
C1042 OR2X1_LOC_436/B OR2X1_LOC_174/Y 0.11fF
C1043 OR2X1_LOC_39/A OR2X1_LOC_71/A 0.86fF
C1044 OR2X1_LOC_74/A OR2X1_LOC_406/A 0.03fF
C1045 AND2X1_LOC_731/Y AND2X1_LOC_220/B 0.03fF
C1046 OR2X1_LOC_44/Y AND2X1_LOC_783/a_36_24# 0.00fF
C1047 AND2X1_LOC_92/Y OR2X1_LOC_120/a_8_216# 0.05fF
C1048 AND2X1_LOC_785/a_36_24# OR2X1_LOC_56/A 0.00fF
C1049 OR2X1_LOC_22/Y OR2X1_LOC_184/Y 0.19fF
C1050 AND2X1_LOC_390/B OR2X1_LOC_761/a_8_216# 0.03fF
C1051 AND2X1_LOC_321/a_8_24# OR2X1_LOC_469/B 0.04fF
C1052 OR2X1_LOC_614/Y OR2X1_LOC_790/A 0.01fF
C1053 OR2X1_LOC_3/B AND2X1_LOC_639/A 0.01fF
C1054 AND2X1_LOC_91/B OR2X1_LOC_624/Y 0.02fF
C1055 OR2X1_LOC_436/Y OR2X1_LOC_468/a_8_216# 0.02fF
C1056 OR2X1_LOC_97/A OR2X1_LOC_645/a_36_216# 0.00fF
C1057 AND2X1_LOC_707/Y AND2X1_LOC_454/a_36_24# 0.01fF
C1058 OR2X1_LOC_30/a_8_216# D_INPUT_6 0.03fF
C1059 D_GATE_479 OR2X1_LOC_467/A 0.01fF
C1060 OR2X1_LOC_22/Y AND2X1_LOC_641/a_8_24# 0.04fF
C1061 AND2X1_LOC_86/B OR2X1_LOC_80/A 0.27fF
C1062 OR2X1_LOC_528/Y AND2X1_LOC_475/Y 0.05fF
C1063 AND2X1_LOC_91/B OR2X1_LOC_391/A 0.62fF
C1064 AND2X1_LOC_227/Y OR2X1_LOC_224/Y 0.02fF
C1065 OR2X1_LOC_467/A OR2X1_LOC_161/B 0.03fF
C1066 OR2X1_LOC_244/B OR2X1_LOC_267/Y 0.47fF
C1067 OR2X1_LOC_842/A OR2X1_LOC_294/Y 0.01fF
C1068 OR2X1_LOC_114/B AND2X1_LOC_295/a_36_24# 0.00fF
C1069 OR2X1_LOC_624/B OR2X1_LOC_80/A 0.13fF
C1070 OR2X1_LOC_40/Y AND2X1_LOC_443/a_36_24# 0.02fF
C1071 OR2X1_LOC_591/Y VDD 0.04fF
C1072 OR2X1_LOC_134/Y OR2X1_LOC_92/Y 0.03fF
C1073 OR2X1_LOC_647/Y OR2X1_LOC_68/B 0.05fF
C1074 OR2X1_LOC_375/A INPUT_6 0.09fF
C1075 OR2X1_LOC_756/B OR2X1_LOC_34/A 0.01fF
C1076 OR2X1_LOC_22/Y OR2X1_LOC_70/A 0.97fF
C1077 AND2X1_LOC_43/B OR2X1_LOC_388/a_8_216# 0.02fF
C1078 OR2X1_LOC_124/B OR2X1_LOC_6/B 0.11fF
C1079 OR2X1_LOC_671/Y OR2X1_LOC_56/A 0.11fF
C1080 OR2X1_LOC_777/a_8_216# OR2X1_LOC_784/B -0.00fF
C1081 AND2X1_LOC_91/B OR2X1_LOC_714/Y 0.01fF
C1082 AND2X1_LOC_40/Y AND2X1_LOC_7/B 0.20fF
C1083 OR2X1_LOC_678/a_8_216# OR2X1_LOC_713/A 0.01fF
C1084 OR2X1_LOC_196/B AND2X1_LOC_31/Y 0.72fF
C1085 OR2X1_LOC_813/A AND2X1_LOC_647/Y 0.01fF
C1086 OR2X1_LOC_596/A AND2X1_LOC_92/Y 0.03fF
C1087 AND2X1_LOC_549/Y AND2X1_LOC_565/a_8_24# 0.19fF
C1088 OR2X1_LOC_106/a_8_216# OR2X1_LOC_56/A 0.00fF
C1089 AND2X1_LOC_64/Y AND2X1_LOC_95/Y 0.73fF
C1090 AND2X1_LOC_83/a_36_24# OR2X1_LOC_78/B 0.01fF
C1091 OR2X1_LOC_855/a_8_216# OR2X1_LOC_637/A 0.47fF
C1092 OR2X1_LOC_36/Y OR2X1_LOC_395/Y 0.09fF
C1093 OR2X1_LOC_160/A OR2X1_LOC_115/B 0.15fF
C1094 AND2X1_LOC_41/A OR2X1_LOC_549/A 0.14fF
C1095 AND2X1_LOC_768/a_8_24# VDD 0.00fF
C1096 AND2X1_LOC_721/Y OR2X1_LOC_427/A 0.03fF
C1097 OR2X1_LOC_516/B AND2X1_LOC_212/Y 0.01fF
C1098 OR2X1_LOC_134/Y OR2X1_LOC_65/B 0.14fF
C1099 OR2X1_LOC_167/Y OR2X1_LOC_331/Y 0.02fF
C1100 AND2X1_LOC_69/a_8_24# OR2X1_LOC_68/B 0.01fF
C1101 OR2X1_LOC_485/Y OR2X1_LOC_59/Y 0.43fF
C1102 OR2X1_LOC_524/Y AND2X1_LOC_469/a_36_24# 0.09fF
C1103 AND2X1_LOC_773/Y AND2X1_LOC_364/A 0.10fF
C1104 AND2X1_LOC_59/Y OR2X1_LOC_703/a_8_216# 0.01fF
C1105 OR2X1_LOC_641/Y OR2X1_LOC_650/a_8_216# 0.03fF
C1106 OR2X1_LOC_471/a_8_216# AND2X1_LOC_7/B 0.06fF
C1107 OR2X1_LOC_537/A AND2X1_LOC_7/B 0.03fF
C1108 OR2X1_LOC_194/B AND2X1_LOC_44/Y 0.01fF
C1109 OR2X1_LOC_851/B OR2X1_LOC_840/A 0.25fF
C1110 OR2X1_LOC_122/a_8_216# OR2X1_LOC_426/B 0.03fF
C1111 OR2X1_LOC_616/Y AND2X1_LOC_580/a_36_24# 0.00fF
C1112 OR2X1_LOC_604/A AND2X1_LOC_456/B 0.06fF
C1113 OR2X1_LOC_715/B OR2X1_LOC_502/A 0.10fF
C1114 AND2X1_LOC_64/Y OR2X1_LOC_99/Y 0.03fF
C1115 OR2X1_LOC_666/A AND2X1_LOC_858/B 0.02fF
C1116 OR2X1_LOC_744/A AND2X1_LOC_468/a_8_24# 0.01fF
C1117 OR2X1_LOC_648/A OR2X1_LOC_78/B 0.38fF
C1118 AND2X1_LOC_721/Y AND2X1_LOC_464/a_8_24# 0.01fF
C1119 OR2X1_LOC_719/Y OR2X1_LOC_722/B 0.07fF
C1120 OR2X1_LOC_417/A OR2X1_LOC_384/a_36_216# 0.01fF
C1121 AND2X1_LOC_22/Y OR2X1_LOC_520/Y 0.07fF
C1122 OR2X1_LOC_319/B OR2X1_LOC_356/a_8_216# 0.01fF
C1123 AND2X1_LOC_663/B AND2X1_LOC_789/Y 0.07fF
C1124 OR2X1_LOC_121/B OR2X1_LOC_712/B 0.03fF
C1125 OR2X1_LOC_419/a_36_216# OR2X1_LOC_419/Y 0.00fF
C1126 OR2X1_LOC_696/A OR2X1_LOC_743/A 2.59fF
C1127 AND2X1_LOC_92/a_8_24# OR2X1_LOC_462/B 0.01fF
C1128 OR2X1_LOC_532/B OR2X1_LOC_446/B 0.03fF
C1129 AND2X1_LOC_181/a_8_24# OR2X1_LOC_744/A 0.01fF
C1130 OR2X1_LOC_155/A OR2X1_LOC_831/B 0.11fF
C1131 OR2X1_LOC_112/B AND2X1_LOC_31/Y 0.06fF
C1132 AND2X1_LOC_364/Y OR2X1_LOC_329/B 0.03fF
C1133 VDD OR2X1_LOC_802/a_8_216# 0.00fF
C1134 AND2X1_LOC_675/Y AND2X1_LOC_549/a_8_24# 0.11fF
C1135 AND2X1_LOC_861/B OR2X1_LOC_56/A 0.07fF
C1136 AND2X1_LOC_181/Y OR2X1_LOC_109/Y 0.04fF
C1137 OR2X1_LOC_45/B OR2X1_LOC_6/A 0.09fF
C1138 OR2X1_LOC_329/B OR2X1_LOC_674/a_8_216# 0.18fF
C1139 OR2X1_LOC_181/B OR2X1_LOC_565/A 0.13fF
C1140 AND2X1_LOC_593/a_8_24# OR2X1_LOC_48/B 0.03fF
C1141 OR2X1_LOC_204/Y OR2X1_LOC_161/B 0.08fF
C1142 OR2X1_LOC_205/a_8_216# AND2X1_LOC_44/Y 0.01fF
C1143 AND2X1_LOC_2/Y D_INPUT_5 0.03fF
C1144 AND2X1_LOC_737/Y AND2X1_LOC_658/B 0.03fF
C1145 OR2X1_LOC_668/a_8_216# AND2X1_LOC_18/Y 0.02fF
C1146 OR2X1_LOC_709/A OR2X1_LOC_154/A 0.09fF
C1147 OR2X1_LOC_3/Y AND2X1_LOC_773/a_8_24# 0.01fF
C1148 OR2X1_LOC_409/B OR2X1_LOC_385/a_8_216# 0.01fF
C1149 OR2X1_LOC_739/Y OR2X1_LOC_740/a_8_216# 0.39fF
C1150 INPUT_0 AND2X1_LOC_39/a_8_24# 0.01fF
C1151 OR2X1_LOC_517/a_8_216# OR2X1_LOC_275/Y 0.40fF
C1152 OR2X1_LOC_186/Y OR2X1_LOC_809/a_8_216# 0.01fF
C1153 AND2X1_LOC_486/Y AND2X1_LOC_469/B 0.22fF
C1154 OR2X1_LOC_753/A OR2X1_LOC_16/A 0.59fF
C1155 AND2X1_LOC_70/Y OR2X1_LOC_620/Y 0.07fF
C1156 OR2X1_LOC_506/A OR2X1_LOC_776/Y 0.14fF
C1157 OR2X1_LOC_599/A OR2X1_LOC_829/A 0.02fF
C1158 OR2X1_LOC_270/Y OR2X1_LOC_367/B 0.03fF
C1159 OR2X1_LOC_78/A OR2X1_LOC_575/A 0.01fF
C1160 OR2X1_LOC_6/A OR2X1_LOC_382/A 0.10fF
C1161 AND2X1_LOC_716/Y OR2X1_LOC_91/A 0.15fF
C1162 OR2X1_LOC_181/B OR2X1_LOC_190/Y 0.06fF
C1163 AND2X1_LOC_657/Y AND2X1_LOC_811/B 0.42fF
C1164 OR2X1_LOC_409/B OR2X1_LOC_376/Y 0.00fF
C1165 AND2X1_LOC_573/a_8_24# AND2X1_LOC_501/Y 0.15fF
C1166 OR2X1_LOC_696/A OR2X1_LOC_125/Y 0.01fF
C1167 OR2X1_LOC_659/B OR2X1_LOC_113/B 0.00fF
C1168 AND2X1_LOC_721/a_8_24# AND2X1_LOC_366/A 0.04fF
C1169 AND2X1_LOC_572/A AND2X1_LOC_243/Y 0.02fF
C1170 AND2X1_LOC_42/B OR2X1_LOC_572/a_8_216# 0.01fF
C1171 AND2X1_LOC_250/a_8_24# OR2X1_LOC_580/A 0.00fF
C1172 OR2X1_LOC_155/a_8_216# OR2X1_LOC_87/A 0.04fF
C1173 AND2X1_LOC_811/B AND2X1_LOC_469/B 0.01fF
C1174 OR2X1_LOC_756/B OR2X1_LOC_400/a_36_216# 0.01fF
C1175 OR2X1_LOC_475/Y AND2X1_LOC_7/B 0.02fF
C1176 OR2X1_LOC_91/A AND2X1_LOC_654/Y 0.09fF
C1177 AND2X1_LOC_857/Y OR2X1_LOC_298/a_36_216# 0.00fF
C1178 AND2X1_LOC_773/Y OR2X1_LOC_3/Y 2.21fF
C1179 OR2X1_LOC_347/B OR2X1_LOC_244/Y 0.10fF
C1180 D_GATE_479 OR2X1_LOC_466/a_8_216# 0.01fF
C1181 OR2X1_LOC_478/Y OR2X1_LOC_470/B 0.02fF
C1182 OR2X1_LOC_505/a_8_216# OR2X1_LOC_74/A 0.03fF
C1183 AND2X1_LOC_345/Y OR2X1_LOC_428/A 0.12fF
C1184 OR2X1_LOC_820/a_8_216# OR2X1_LOC_820/B 0.05fF
C1185 AND2X1_LOC_486/Y AND2X1_LOC_733/Y 0.42fF
C1186 AND2X1_LOC_12/Y AND2X1_LOC_2/Y 1.05fF
C1187 AND2X1_LOC_225/a_8_24# OR2X1_LOC_558/A 0.09fF
C1188 AND2X1_LOC_719/Y OR2X1_LOC_26/Y 0.02fF
C1189 OR2X1_LOC_566/Y OR2X1_LOC_568/a_8_216# 0.03fF
C1190 OR2X1_LOC_466/a_8_216# OR2X1_LOC_161/B 0.02fF
C1191 OR2X1_LOC_299/Y OR2X1_LOC_12/Y 0.01fF
C1192 OR2X1_LOC_696/A OR2X1_LOC_225/a_8_216# 0.01fF
C1193 OR2X1_LOC_87/A AND2X1_LOC_18/Y 0.16fF
C1194 OR2X1_LOC_133/a_8_216# OR2X1_LOC_74/A 0.40fF
C1195 AND2X1_LOC_302/a_8_24# OR2X1_LOC_426/B 0.03fF
C1196 OR2X1_LOC_703/A OR2X1_LOC_620/Y 0.07fF
C1197 VDD OR2X1_LOC_264/a_8_216# 0.21fF
C1198 OR2X1_LOC_154/A AND2X1_LOC_70/Y 0.26fF
C1199 OR2X1_LOC_652/a_8_216# OR2X1_LOC_78/A 0.01fF
C1200 OR2X1_LOC_160/B OR2X1_LOC_719/Y 0.02fF
C1201 AND2X1_LOC_861/B AND2X1_LOC_850/Y 0.00fF
C1202 OR2X1_LOC_518/a_8_216# OR2X1_LOC_417/A 0.03fF
C1203 OR2X1_LOC_59/Y OR2X1_LOC_39/A 6.03fF
C1204 OR2X1_LOC_62/A AND2X1_LOC_36/Y 0.09fF
C1205 OR2X1_LOC_92/Y OR2X1_LOC_586/a_8_216# 0.01fF
C1206 OR2X1_LOC_464/A OR2X1_LOC_737/A 0.15fF
C1207 OR2X1_LOC_114/B OR2X1_LOC_269/B 0.03fF
C1208 AND2X1_LOC_513/a_8_24# OR2X1_LOC_48/B 0.03fF
C1209 OR2X1_LOC_61/B OR2X1_LOC_61/a_8_216# 0.05fF
C1210 OR2X1_LOC_648/A AND2X1_LOC_601/a_36_24# 0.01fF
C1211 OR2X1_LOC_11/Y AND2X1_LOC_637/a_8_24# 0.01fF
C1212 OR2X1_LOC_139/A OR2X1_LOC_121/B 0.03fF
C1213 INPUT_0 AND2X1_LOC_43/B 0.29fF
C1214 AND2X1_LOC_40/Y OR2X1_LOC_318/Y 0.03fF
C1215 OR2X1_LOC_756/B OR2X1_LOC_506/A 0.03fF
C1216 AND2X1_LOC_719/Y OR2X1_LOC_89/A 0.03fF
C1217 AND2X1_LOC_311/a_36_24# OR2X1_LOC_161/A 0.01fF
C1218 AND2X1_LOC_59/Y AND2X1_LOC_437/a_36_24# 0.00fF
C1219 AND2X1_LOC_732/B OR2X1_LOC_52/B 0.03fF
C1220 OR2X1_LOC_410/a_8_216# OR2X1_LOC_375/A 0.06fF
C1221 OR2X1_LOC_696/A OR2X1_LOC_409/B 0.05fF
C1222 AND2X1_LOC_95/Y OR2X1_LOC_464/A 0.03fF
C1223 OR2X1_LOC_74/Y AND2X1_LOC_76/a_8_24# 0.23fF
C1224 OR2X1_LOC_42/a_8_216# OR2X1_LOC_56/A 0.04fF
C1225 AND2X1_LOC_753/B AND2X1_LOC_53/a_36_24# 0.00fF
C1226 AND2X1_LOC_22/Y AND2X1_LOC_107/a_8_24# 0.06fF
C1227 OR2X1_LOC_604/A AND2X1_LOC_717/B 0.14fF
C1228 OR2X1_LOC_87/B AND2X1_LOC_92/Y 0.03fF
C1229 AND2X1_LOC_47/Y OR2X1_LOC_140/B 0.04fF
C1230 OR2X1_LOC_850/A OR2X1_LOC_362/A 0.02fF
C1231 OR2X1_LOC_3/Y AND2X1_LOC_243/Y 0.08fF
C1232 OR2X1_LOC_684/Y OR2X1_LOC_16/A 0.39fF
C1233 OR2X1_LOC_348/Y AND2X1_LOC_3/Y 0.03fF
C1234 OR2X1_LOC_160/A OR2X1_LOC_840/A 0.10fF
C1235 OR2X1_LOC_287/B OR2X1_LOC_66/A 0.03fF
C1236 AND2X1_LOC_555/a_8_24# OR2X1_LOC_481/Y 0.04fF
C1237 OR2X1_LOC_744/A AND2X1_LOC_859/Y 0.07fF
C1238 GATE_366 OR2X1_LOC_91/A 0.06fF
C1239 VDD OR2X1_LOC_438/a_8_216# 0.21fF
C1240 OR2X1_LOC_759/A OR2X1_LOC_258/a_8_216# 0.01fF
C1241 OR2X1_LOC_40/Y OR2X1_LOC_258/Y 0.61fF
C1242 OR2X1_LOC_792/Y OR2X1_LOC_807/B 0.04fF
C1243 AND2X1_LOC_40/Y OR2X1_LOC_407/a_8_216# 0.01fF
C1244 OR2X1_LOC_502/A OR2X1_LOC_215/Y 0.03fF
C1245 AND2X1_LOC_738/B AND2X1_LOC_645/A 0.01fF
C1246 AND2X1_LOC_40/Y OR2X1_LOC_805/A 0.03fF
C1247 OR2X1_LOC_70/Y OR2X1_LOC_485/Y 0.07fF
C1248 AND2X1_LOC_568/B AND2X1_LOC_568/a_8_24# 0.00fF
C1249 OR2X1_LOC_178/Y OR2X1_LOC_7/A 0.04fF
C1250 OR2X1_LOC_805/a_8_216# OR2X1_LOC_362/B 0.01fF
C1251 OR2X1_LOC_538/A OR2X1_LOC_269/B 0.03fF
C1252 AND2X1_LOC_845/Y AND2X1_LOC_244/A 0.03fF
C1253 OR2X1_LOC_837/A AND2X1_LOC_34/Y 0.02fF
C1254 AND2X1_LOC_211/B OR2X1_LOC_59/Y 0.03fF
C1255 OR2X1_LOC_158/A OR2X1_LOC_416/Y 0.03fF
C1256 VDD OR2X1_LOC_863/B 0.12fF
C1257 OR2X1_LOC_312/Y OR2X1_LOC_91/A 0.07fF
C1258 AND2X1_LOC_70/Y OR2X1_LOC_856/a_8_216# 0.01fF
C1259 OR2X1_LOC_856/B AND2X1_LOC_536/a_36_24# 0.01fF
C1260 AND2X1_LOC_190/a_36_24# OR2X1_LOC_485/A 0.00fF
C1261 OR2X1_LOC_405/A OR2X1_LOC_624/A 0.24fF
C1262 OR2X1_LOC_663/A OR2X1_LOC_849/A 0.03fF
C1263 OR2X1_LOC_54/Y OR2X1_LOC_382/a_8_216# -0.03fF
C1264 AND2X1_LOC_41/A OR2X1_LOC_711/A 0.01fF
C1265 AND2X1_LOC_70/Y OR2X1_LOC_778/A 0.01fF
C1266 OR2X1_LOC_859/a_8_216# OR2X1_LOC_810/A 0.09fF
C1267 OR2X1_LOC_6/B OR2X1_LOC_611/a_8_216# 0.00fF
C1268 OR2X1_LOC_656/Y OR2X1_LOC_99/Y 0.02fF
C1269 OR2X1_LOC_485/a_8_216# OR2X1_LOC_44/Y 0.07fF
C1270 AND2X1_LOC_112/a_8_24# OR2X1_LOC_64/Y 0.01fF
C1271 OR2X1_LOC_76/A OR2X1_LOC_66/A 0.14fF
C1272 OR2X1_LOC_3/Y AND2X1_LOC_377/Y 0.16fF
C1273 OR2X1_LOC_426/B AND2X1_LOC_663/B 0.10fF
C1274 OR2X1_LOC_215/Y AND2X1_LOC_230/a_8_24# 0.23fF
C1275 AND2X1_LOC_136/a_8_24# OR2X1_LOC_78/B 0.03fF
C1276 AND2X1_LOC_141/B AND2X1_LOC_141/a_36_24# 0.00fF
C1277 OR2X1_LOC_160/B OR2X1_LOC_474/a_8_216# 0.02fF
C1278 OR2X1_LOC_774/Y OR2X1_LOC_862/A 0.14fF
C1279 AND2X1_LOC_33/Y AND2X1_LOC_35/a_8_24# 0.18fF
C1280 OR2X1_LOC_256/Y OR2X1_LOC_7/A 0.04fF
C1281 OR2X1_LOC_49/A D_INPUT_3 0.04fF
C1282 AND2X1_LOC_466/a_8_24# AND2X1_LOC_452/Y 0.04fF
C1283 OR2X1_LOC_698/Y OR2X1_LOC_258/a_8_216# 0.01fF
C1284 OR2X1_LOC_462/B OR2X1_LOC_185/A 0.01fF
C1285 AND2X1_LOC_648/B OR2X1_LOC_428/A 0.03fF
C1286 OR2X1_LOC_748/A OR2X1_LOC_427/A 0.01fF
C1287 OR2X1_LOC_185/A OR2X1_LOC_483/a_8_216# 0.02fF
C1288 AND2X1_LOC_56/B AND2X1_LOC_16/a_36_24# 0.00fF
C1289 OR2X1_LOC_648/B D_INPUT_0 0.03fF
C1290 OR2X1_LOC_669/a_8_216# OR2X1_LOC_278/Y 0.01fF
C1291 OR2X1_LOC_160/B OR2X1_LOC_859/A 0.00fF
C1292 AND2X1_LOC_361/a_8_24# AND2X1_LOC_227/Y 0.01fF
C1293 OR2X1_LOC_140/B OR2X1_LOC_598/A 0.04fF
C1294 OR2X1_LOC_590/a_8_216# OR2X1_LOC_718/a_8_216# 0.47fF
C1295 OR2X1_LOC_648/a_8_216# AND2X1_LOC_18/Y 0.01fF
C1296 OR2X1_LOC_45/a_8_216# OR2X1_LOC_44/Y 0.05fF
C1297 AND2X1_LOC_665/a_8_24# OR2X1_LOC_719/B 0.01fF
C1298 OR2X1_LOC_701/Y OR2X1_LOC_44/Y 0.10fF
C1299 OR2X1_LOC_700/Y OR2X1_LOC_701/a_8_216# 0.02fF
C1300 AND2X1_LOC_403/B OR2X1_LOC_44/Y 0.23fF
C1301 OR2X1_LOC_724/A OR2X1_LOC_308/Y 0.21fF
C1302 AND2X1_LOC_215/Y AND2X1_LOC_640/a_8_24# 0.01fF
C1303 D_INPUT_3 OR2X1_LOC_381/a_36_216# 0.03fF
C1304 AND2X1_LOC_334/Y AND2X1_LOC_634/Y 0.00fF
C1305 OR2X1_LOC_275/A OR2X1_LOC_517/A 0.24fF
C1306 AND2X1_LOC_392/A OR2X1_LOC_71/Y 0.03fF
C1307 OR2X1_LOC_610/a_8_216# OR2X1_LOC_647/B 0.03fF
C1308 OR2X1_LOC_368/a_8_216# OR2X1_LOC_31/Y 0.09fF
C1309 AND2X1_LOC_12/Y OR2X1_LOC_269/B 0.28fF
C1310 OR2X1_LOC_349/B OR2X1_LOC_580/A 0.00fF
C1311 AND2X1_LOC_738/B AND2X1_LOC_477/A 1.00fF
C1312 OR2X1_LOC_649/a_36_216# AND2X1_LOC_92/Y 0.00fF
C1313 AND2X1_LOC_217/Y OR2X1_LOC_95/Y 0.16fF
C1314 AND2X1_LOC_112/a_8_24# OR2X1_LOC_417/A 0.01fF
C1315 OR2X1_LOC_719/Y OR2X1_LOC_553/A 0.01fF
C1316 OR2X1_LOC_379/Y OR2X1_LOC_654/A 0.03fF
C1317 OR2X1_LOC_169/a_8_216# OR2X1_LOC_468/Y 0.01fF
C1318 OR2X1_LOC_476/B OR2X1_LOC_334/B 0.01fF
C1319 OR2X1_LOC_773/B OR2X1_LOC_774/Y 0.09fF
C1320 OR2X1_LOC_40/Y AND2X1_LOC_318/Y 0.02fF
C1321 AND2X1_LOC_95/Y OR2X1_LOC_445/a_36_216# 0.02fF
C1322 OR2X1_LOC_47/Y OR2X1_LOC_584/Y 0.01fF
C1323 OR2X1_LOC_864/A AND2X1_LOC_81/B 0.03fF
C1324 AND2X1_LOC_121/a_8_24# AND2X1_LOC_845/Y 0.03fF
C1325 AND2X1_LOC_40/Y OR2X1_LOC_436/a_8_216# 0.01fF
C1326 OR2X1_LOC_759/A AND2X1_LOC_866/A 0.01fF
C1327 OR2X1_LOC_306/Y AND2X1_LOC_512/a_8_24# 0.03fF
C1328 OR2X1_LOC_436/Y OR2X1_LOC_66/A 0.03fF
C1329 VDD OR2X1_LOC_276/A 0.21fF
C1330 OR2X1_LOC_304/Y OR2X1_LOC_427/A 0.00fF
C1331 AND2X1_LOC_286/Y AND2X1_LOC_288/a_36_24# 0.01fF
C1332 OR2X1_LOC_510/Y AND2X1_LOC_3/Y 0.09fF
C1333 OR2X1_LOC_82/a_8_216# OR2X1_LOC_83/A 0.02fF
C1334 OR2X1_LOC_817/Y AND2X1_LOC_847/Y 0.05fF
C1335 AND2X1_LOC_81/B OR2X1_LOC_633/B 0.02fF
C1336 AND2X1_LOC_49/a_8_24# OR2X1_LOC_633/B 0.01fF
C1337 OR2X1_LOC_757/A OR2X1_LOC_95/Y 0.02fF
C1338 OR2X1_LOC_816/A AND2X1_LOC_790/a_8_24# 0.03fF
C1339 AND2X1_LOC_70/Y AND2X1_LOC_684/a_8_24# 0.01fF
C1340 OR2X1_LOC_70/Y OR2X1_LOC_39/A 1.89fF
C1341 OR2X1_LOC_479/Y OR2X1_LOC_130/A 0.03fF
C1342 AND2X1_LOC_589/a_36_24# OR2X1_LOC_130/A 0.01fF
C1343 AND2X1_LOC_384/a_8_24# OR2X1_LOC_383/Y 0.24fF
C1344 OR2X1_LOC_475/Y OR2X1_LOC_805/A 0.01fF
C1345 AND2X1_LOC_476/A AND2X1_LOC_219/Y -0.08fF
C1346 AND2X1_LOC_12/Y OR2X1_LOC_215/A 0.41fF
C1347 AND2X1_LOC_719/a_8_24# AND2X1_LOC_859/Y 0.03fF
C1348 AND2X1_LOC_658/B AND2X1_LOC_808/A 0.03fF
C1349 OR2X1_LOC_40/Y OR2X1_LOC_815/Y 0.02fF
C1350 AND2X1_LOC_191/Y AND2X1_LOC_569/a_8_24# 0.05fF
C1351 OR2X1_LOC_46/A OR2X1_LOC_48/B 0.04fF
C1352 OR2X1_LOC_154/A OR2X1_LOC_206/a_8_216# 0.01fF
C1353 OR2X1_LOC_604/A OR2X1_LOC_419/a_36_216# 0.00fF
C1354 OR2X1_LOC_811/A OR2X1_LOC_814/A 0.04fF
C1355 OR2X1_LOC_810/A AND2X1_LOC_3/Y 0.03fF
C1356 OR2X1_LOC_321/Y OR2X1_LOC_36/Y 0.00fF
C1357 AND2X1_LOC_40/Y AND2X1_LOC_441/a_8_24# 0.04fF
C1358 OR2X1_LOC_643/A AND2X1_LOC_42/B 0.04fF
C1359 OR2X1_LOC_812/B OR2X1_LOC_383/Y 0.06fF
C1360 AND2X1_LOC_788/a_8_24# OR2X1_LOC_331/Y 0.02fF
C1361 OR2X1_LOC_833/Y AND2X1_LOC_31/Y 0.02fF
C1362 OR2X1_LOC_631/B OR2X1_LOC_629/a_8_216# 0.01fF
C1363 OR2X1_LOC_18/Y OR2X1_LOC_46/A 0.04fF
C1364 AND2X1_LOC_42/B OR2X1_LOC_124/Y 0.03fF
C1365 OR2X1_LOC_154/A OR2X1_LOC_404/Y 0.15fF
C1366 AND2X1_LOC_647/Y AND2X1_LOC_606/a_8_24# 0.01fF
C1367 OR2X1_LOC_235/B AND2X1_LOC_813/a_8_24# 0.03fF
C1368 AND2X1_LOC_42/B OR2X1_LOC_778/Y 0.02fF
C1369 OR2X1_LOC_70/Y AND2X1_LOC_569/a_8_24# 0.17fF
C1370 AND2X1_LOC_173/a_36_24# D_INPUT_0 0.00fF
C1371 OR2X1_LOC_804/B OR2X1_LOC_269/B 0.12fF
C1372 AND2X1_LOC_120/a_8_24# AND2X1_LOC_806/A 0.01fF
C1373 OR2X1_LOC_524/Y AND2X1_LOC_803/a_8_24# 0.29fF
C1374 OR2X1_LOC_795/a_8_216# AND2X1_LOC_92/Y 0.06fF
C1375 OR2X1_LOC_124/B OR2X1_LOC_598/A 0.02fF
C1376 OR2X1_LOC_690/A OR2X1_LOC_27/a_8_216# 0.01fF
C1377 AND2X1_LOC_13/a_8_24# OR2X1_LOC_155/A 0.04fF
C1378 AND2X1_LOC_562/B OR2X1_LOC_615/Y 0.01fF
C1379 OR2X1_LOC_70/Y AND2X1_LOC_211/B 0.03fF
C1380 OR2X1_LOC_417/Y AND2X1_LOC_661/A 0.03fF
C1381 OR2X1_LOC_756/B D_INPUT_1 0.22fF
C1382 AND2X1_LOC_729/B OR2X1_LOC_585/A 0.06fF
C1383 OR2X1_LOC_243/A OR2X1_LOC_244/A 0.01fF
C1384 OR2X1_LOC_70/Y OR2X1_LOC_429/Y 0.06fF
C1385 OR2X1_LOC_504/Y OR2X1_LOC_39/A 0.43fF
C1386 VDD OR2X1_LOC_512/Y 0.00fF
C1387 AND2X1_LOC_326/a_8_24# AND2X1_LOC_354/B 0.04fF
C1388 AND2X1_LOC_227/Y OR2X1_LOC_18/Y 0.05fF
C1389 AND2X1_LOC_737/Y OR2X1_LOC_47/Y 0.02fF
C1390 INPUT_5 OR2X1_LOC_2/a_8_216# 0.06fF
C1391 AND2X1_LOC_61/Y OR2X1_LOC_72/Y 0.01fF
C1392 AND2X1_LOC_514/Y AND2X1_LOC_211/B 0.08fF
C1393 OR2X1_LOC_160/A OR2X1_LOC_241/Y 0.07fF
C1394 OR2X1_LOC_115/B OR2X1_LOC_130/Y 0.00fF
C1395 OR2X1_LOC_344/A D_GATE_366 0.13fF
C1396 AND2X1_LOC_70/Y OR2X1_LOC_560/A 0.02fF
C1397 AND2X1_LOC_56/B OR2X1_LOC_532/B 0.27fF
C1398 AND2X1_LOC_53/Y OR2X1_LOC_793/A 0.02fF
C1399 AND2X1_LOC_70/Y OR2X1_LOC_198/A 0.17fF
C1400 OR2X1_LOC_47/Y OR2X1_LOC_394/Y 0.37fF
C1401 OR2X1_LOC_151/A OR2X1_LOC_140/Y 0.87fF
C1402 OR2X1_LOC_659/B OR2X1_LOC_532/B 0.02fF
C1403 OR2X1_LOC_436/Y OR2X1_LOC_799/a_36_216# 0.00fF
C1404 AND2X1_LOC_554/Y OR2X1_LOC_47/Y 0.03fF
C1405 AND2X1_LOC_8/Y OR2X1_LOC_532/B 0.07fF
C1406 OR2X1_LOC_364/A OR2X1_LOC_440/A 0.11fF
C1407 OR2X1_LOC_13/B OR2X1_LOC_131/a_8_216# 0.02fF
C1408 OR2X1_LOC_532/B OR2X1_LOC_720/a_36_216# 0.00fF
C1409 OR2X1_LOC_62/B AND2X1_LOC_4/a_8_24# 0.01fF
C1410 OR2X1_LOC_47/Y OR2X1_LOC_48/a_8_216# 0.07fF
C1411 AND2X1_LOC_65/a_8_24# OR2X1_LOC_68/B 0.01fF
C1412 OR2X1_LOC_18/Y OR2X1_LOC_813/Y 0.01fF
C1413 AND2X1_LOC_42/B OR2X1_LOC_113/A 0.00fF
C1414 OR2X1_LOC_710/A AND2X1_LOC_7/B 0.13fF
C1415 OR2X1_LOC_41/Y OR2X1_LOC_48/B 0.12fF
C1416 OR2X1_LOC_626/a_8_216# OR2X1_LOC_95/Y 0.17fF
C1417 OR2X1_LOC_437/Y OR2X1_LOC_39/A 0.38fF
C1418 AND2X1_LOC_64/Y AND2X1_LOC_22/Y 0.43fF
C1419 AND2X1_LOC_778/Y OR2X1_LOC_142/Y 0.07fF
C1420 AND2X1_LOC_727/A AND2X1_LOC_802/a_8_24# 0.01fF
C1421 OR2X1_LOC_809/a_8_216# OR2X1_LOC_112/B 0.02fF
C1422 AND2X1_LOC_47/Y AND2X1_LOC_18/a_8_24# 0.01fF
C1423 OR2X1_LOC_444/B AND2X1_LOC_442/a_8_24# 0.01fF
C1424 OR2X1_LOC_123/B D_INPUT_0 0.05fF
C1425 OR2X1_LOC_280/a_8_216# AND2X1_LOC_851/B 0.06fF
C1426 OR2X1_LOC_629/B AND2X1_LOC_36/Y 0.01fF
C1427 AND2X1_LOC_259/Y D_INPUT_3 0.00fF
C1428 AND2X1_LOC_465/A OR2X1_LOC_428/A 0.05fF
C1429 AND2X1_LOC_391/Y OR2X1_LOC_13/B 0.03fF
C1430 OR2X1_LOC_599/A OR2X1_LOC_597/Y 0.01fF
C1431 AND2X1_LOC_858/B OR2X1_LOC_13/B 0.01fF
C1432 OR2X1_LOC_70/Y OR2X1_LOC_428/a_8_216# 0.01fF
C1433 OR2X1_LOC_91/A OR2X1_LOC_13/B 3.20fF
C1434 OR2X1_LOC_136/Y AND2X1_LOC_358/Y 0.56fF
C1435 OR2X1_LOC_78/B OR2X1_LOC_112/A 0.37fF
C1436 OR2X1_LOC_231/A OR2X1_LOC_68/B 0.28fF
C1437 AND2X1_LOC_812/a_8_24# OR2X1_LOC_74/A 0.05fF
C1438 AND2X1_LOC_722/Y OR2X1_LOC_437/A 0.01fF
C1439 OR2X1_LOC_36/Y AND2X1_LOC_646/a_36_24# 0.00fF
C1440 AND2X1_LOC_48/A AND2X1_LOC_519/a_8_24# 0.10fF
C1441 OR2X1_LOC_280/Y OR2X1_LOC_47/Y 0.02fF
C1442 AND2X1_LOC_91/a_8_24# OR2X1_LOC_161/B 0.01fF
C1443 OR2X1_LOC_97/A AND2X1_LOC_44/Y 0.03fF
C1444 OR2X1_LOC_858/B OR2X1_LOC_580/A 0.02fF
C1445 OR2X1_LOC_70/Y OR2X1_LOC_760/a_8_216# 0.14fF
C1446 OR2X1_LOC_539/Y OR2X1_LOC_854/A 0.20fF
C1447 AND2X1_LOC_59/Y OR2X1_LOC_641/B 0.01fF
C1448 AND2X1_LOC_45/a_8_24# AND2X1_LOC_53/Y 0.03fF
C1449 OR2X1_LOC_847/A OR2X1_LOC_80/A 0.03fF
C1450 OR2X1_LOC_208/A OR2X1_LOC_648/B 0.04fF
C1451 AND2X1_LOC_81/B OR2X1_LOC_608/Y 0.01fF
C1452 OR2X1_LOC_233/a_36_216# D_INPUT_1 0.00fF
C1453 OR2X1_LOC_417/Y AND2X1_LOC_810/Y 0.72fF
C1454 AND2X1_LOC_784/A AND2X1_LOC_784/a_36_24# 0.01fF
C1455 OR2X1_LOC_400/A OR2X1_LOC_398/Y 0.01fF
C1456 OR2X1_LOC_340/Y OR2X1_LOC_68/B 0.02fF
C1457 AND2X1_LOC_211/B AND2X1_LOC_641/a_8_24# 0.01fF
C1458 OR2X1_LOC_212/A OR2X1_LOC_353/a_36_216# 0.00fF
C1459 AND2X1_LOC_18/Y OR2X1_LOC_390/B 0.01fF
C1460 AND2X1_LOC_191/Y AND2X1_LOC_781/Y 0.03fF
C1461 OR2X1_LOC_654/a_8_216# AND2X1_LOC_7/B 0.01fF
C1462 AND2X1_LOC_278/a_36_24# OR2X1_LOC_80/A 0.01fF
C1463 OR2X1_LOC_447/A AND2X1_LOC_419/a_8_24# 0.17fF
C1464 OR2X1_LOC_130/A OR2X1_LOC_68/B 0.25fF
C1465 OR2X1_LOC_793/B OR2X1_LOC_801/B 0.04fF
C1466 OR2X1_LOC_377/A OR2X1_LOC_71/A 0.03fF
C1467 AND2X1_LOC_776/Y AND2X1_LOC_776/a_8_24# 0.09fF
C1468 OR2X1_LOC_756/B OR2X1_LOC_180/B 0.06fF
C1469 OR2X1_LOC_44/Y AND2X1_LOC_570/a_8_24# 0.14fF
C1470 OR2X1_LOC_116/a_8_216# OR2X1_LOC_560/A 0.00fF
C1471 OR2X1_LOC_190/A OR2X1_LOC_562/A 0.03fF
C1472 OR2X1_LOC_479/Y OR2X1_LOC_365/B 0.03fF
C1473 OR2X1_LOC_135/Y OR2X1_LOC_589/A 0.02fF
C1474 OR2X1_LOC_429/Y OR2X1_LOC_70/A 0.17fF
C1475 AND2X1_LOC_8/a_8_24# OR2X1_LOC_54/Y 0.03fF
C1476 AND2X1_LOC_573/A OR2X1_LOC_13/B 0.07fF
C1477 OR2X1_LOC_22/Y OR2X1_LOC_47/Y 0.14fF
C1478 OR2X1_LOC_156/a_8_216# OR2X1_LOC_803/A 0.01fF
C1479 OR2X1_LOC_85/A OR2X1_LOC_71/A 0.85fF
C1480 AND2X1_LOC_592/Y AND2X1_LOC_705/Y 0.00fF
C1481 OR2X1_LOC_574/A AND2X1_LOC_31/Y 0.06fF
C1482 OR2X1_LOC_271/Y OR2X1_LOC_521/a_8_216# 0.19fF
C1483 AND2X1_LOC_612/a_8_24# OR2X1_LOC_68/B 0.01fF
C1484 AND2X1_LOC_229/a_8_24# OR2X1_LOC_160/B 0.03fF
C1485 AND2X1_LOC_64/Y OR2X1_LOC_244/B 0.00fF
C1486 OR2X1_LOC_185/A AND2X1_LOC_591/a_8_24# 0.00fF
C1487 OR2X1_LOC_549/B OR2X1_LOC_756/B 0.00fF
C1488 OR2X1_LOC_392/B AND2X1_LOC_92/Y 0.07fF
C1489 OR2X1_LOC_22/Y AND2X1_LOC_461/a_8_24# 0.05fF
C1490 AND2X1_LOC_719/Y AND2X1_LOC_552/A 0.03fF
C1491 OR2X1_LOC_111/Y AND2X1_LOC_660/A 0.08fF
C1492 OR2X1_LOC_696/A AND2X1_LOC_374/a_8_24# 0.02fF
C1493 OR2X1_LOC_447/Y OR2X1_LOC_779/Y 0.10fF
C1494 AND2X1_LOC_43/B OR2X1_LOC_195/a_36_216# 0.01fF
C1495 OR2X1_LOC_449/B OR2X1_LOC_728/A 0.04fF
C1496 VDD OR2X1_LOC_294/Y 0.41fF
C1497 OR2X1_LOC_473/Y OR2X1_LOC_228/Y 0.01fF
C1498 AND2X1_LOC_70/Y OR2X1_LOC_435/A 0.26fF
C1499 OR2X1_LOC_598/Y OR2X1_LOC_648/B 0.01fF
C1500 OR2X1_LOC_338/a_36_216# OR2X1_LOC_160/B 0.00fF
C1501 OR2X1_LOC_78/A OR2X1_LOC_161/B 0.54fF
C1502 VDD OR2X1_LOC_550/a_8_216# 0.00fF
C1503 OR2X1_LOC_404/Y OR2X1_LOC_560/A 0.03fF
C1504 OR2X1_LOC_500/A OR2X1_LOC_844/B 0.14fF
C1505 AND2X1_LOC_232/a_8_24# OR2X1_LOC_633/A 0.03fF
C1506 AND2X1_LOC_744/a_8_24# AND2X1_LOC_44/Y 0.01fF
C1507 AND2X1_LOC_541/Y VDD 0.19fF
C1508 AND2X1_LOC_39/a_8_24# AND2X1_LOC_7/B 0.01fF
C1509 AND2X1_LOC_200/a_8_24# AND2X1_LOC_207/B 0.01fF
C1510 VDD OR2X1_LOC_641/A 0.14fF
C1511 OR2X1_LOC_40/Y OR2X1_LOC_759/A 0.05fF
C1512 OR2X1_LOC_512/A AND2X1_LOC_22/Y 0.01fF
C1513 AND2X1_LOC_64/Y OR2X1_LOC_630/a_8_216# 0.01fF
C1514 VDD OR2X1_LOC_733/A 0.12fF
C1515 OR2X1_LOC_47/Y AND2X1_LOC_808/A 0.05fF
C1516 OR2X1_LOC_97/A OR2X1_LOC_61/a_8_216# 0.01fF
C1517 OR2X1_LOC_160/B OR2X1_LOC_66/A 0.42fF
C1518 AND2X1_LOC_64/Y OR2X1_LOC_664/a_8_216# 0.01fF
C1519 OR2X1_LOC_62/B OR2X1_LOC_68/B 0.08fF
C1520 OR2X1_LOC_139/A OR2X1_LOC_856/B 0.07fF
C1521 AND2X1_LOC_392/A OR2X1_LOC_426/B 0.26fF
C1522 AND2X1_LOC_47/Y OR2X1_LOC_675/Y 0.02fF
C1523 AND2X1_LOC_564/B OR2X1_LOC_109/Y 0.00fF
C1524 OR2X1_LOC_653/Y AND2X1_LOC_60/a_8_24# 0.03fF
C1525 AND2X1_LOC_64/Y AND2X1_LOC_153/a_8_24# 0.01fF
C1526 AND2X1_LOC_40/Y OR2X1_LOC_580/B 0.20fF
C1527 AND2X1_LOC_84/Y OR2X1_LOC_32/B 0.03fF
C1528 OR2X1_LOC_319/B OR2X1_LOC_356/A 0.15fF
C1529 OR2X1_LOC_109/Y OR2X1_LOC_368/Y 0.01fF
C1530 OR2X1_LOC_696/A OR2X1_LOC_497/Y 0.22fF
C1531 OR2X1_LOC_149/B OR2X1_LOC_375/A 0.72fF
C1532 AND2X1_LOC_523/a_8_24# OR2X1_LOC_428/A 0.01fF
C1533 VDD OR2X1_LOC_107/a_8_216# 0.00fF
C1534 OR2X1_LOC_715/B OR2X1_LOC_201/A 0.08fF
C1535 AND2X1_LOC_364/A OR2X1_LOC_12/Y 0.23fF
C1536 AND2X1_LOC_43/B AND2X1_LOC_7/B 0.37fF
C1537 OR2X1_LOC_139/A OR2X1_LOC_793/a_8_216# 0.40fF
C1538 AND2X1_LOC_849/A OR2X1_LOC_437/A 0.14fF
C1539 OR2X1_LOC_456/A D_GATE_366 0.00fF
C1540 OR2X1_LOC_45/B OR2X1_LOC_45/a_8_216# 0.08fF
C1541 AND2X1_LOC_95/Y OR2X1_LOC_342/A 0.00fF
C1542 OR2X1_LOC_866/B OR2X1_LOC_848/B 0.09fF
C1543 AND2X1_LOC_662/B AND2X1_LOC_786/Y 0.07fF
C1544 OR2X1_LOC_664/Y OR2X1_LOC_563/A 0.03fF
C1545 OR2X1_LOC_40/Y OR2X1_LOC_698/Y 0.01fF
C1546 OR2X1_LOC_106/Y OR2X1_LOC_271/Y 0.00fF
C1547 AND2X1_LOC_362/a_8_24# OR2X1_LOC_666/A 0.01fF
C1548 OR2X1_LOC_158/A OR2X1_LOC_281/a_8_216# 0.01fF
C1549 AND2X1_LOC_95/Y OR2X1_LOC_185/a_8_216# 0.01fF
C1550 OR2X1_LOC_486/B OR2X1_LOC_726/a_8_216# 0.47fF
C1551 OR2X1_LOC_237/Y OR2X1_LOC_428/A 0.01fF
C1552 INPUT_1 OR2X1_LOC_300/a_8_216# 0.01fF
C1553 INPUT_0 AND2X1_LOC_434/Y 0.17fF
C1554 INPUT_0 AND2X1_LOC_219/Y 0.00fF
C1555 AND2X1_LOC_22/Y AND2X1_LOC_369/a_8_24# 0.09fF
C1556 AND2X1_LOC_729/Y OR2X1_LOC_16/A 0.03fF
C1557 OR2X1_LOC_602/A OR2X1_LOC_161/B 0.02fF
C1558 AND2X1_LOC_474/A OR2X1_LOC_59/Y 0.03fF
C1559 AND2X1_LOC_64/Y OR2X1_LOC_296/a_8_216# 0.01fF
C1560 AND2X1_LOC_587/a_8_24# AND2X1_LOC_51/A 0.01fF
C1561 OR2X1_LOC_45/B AND2X1_LOC_831/a_8_24# 0.01fF
C1562 OR2X1_LOC_814/A OR2X1_LOC_777/B 0.07fF
C1563 OR2X1_LOC_678/Y OR2X1_LOC_715/A 0.00fF
C1564 AND2X1_LOC_572/A OR2X1_LOC_12/Y 0.68fF
C1565 OR2X1_LOC_45/B OR2X1_LOC_44/Y 0.19fF
C1566 AND2X1_LOC_12/Y OR2X1_LOC_338/a_8_216# 0.01fF
C1567 OR2X1_LOC_203/a_8_216# OR2X1_LOC_549/A 0.03fF
C1568 OR2X1_LOC_435/B OR2X1_LOC_78/A 0.23fF
C1569 OR2X1_LOC_493/a_8_216# OR2X1_LOC_473/a_8_216# 0.47fF
C1570 AND2X1_LOC_48/a_8_24# OR2X1_LOC_78/A 0.01fF
C1571 AND2X1_LOC_731/a_8_24# AND2X1_LOC_191/Y 0.05fF
C1572 OR2X1_LOC_188/Y OR2X1_LOC_564/A 0.04fF
C1573 OR2X1_LOC_176/Y AND2X1_LOC_566/a_8_24# 0.17fF
C1574 AND2X1_LOC_706/Y AND2X1_LOC_319/A 0.07fF
C1575 AND2X1_LOC_810/A AND2X1_LOC_702/Y 0.02fF
C1576 AND2X1_LOC_544/Y AND2X1_LOC_148/Y 0.03fF
C1577 AND2X1_LOC_91/B AND2X1_LOC_42/B 0.11fF
C1578 OR2X1_LOC_738/A OR2X1_LOC_726/A 0.11fF
C1579 AND2X1_LOC_40/Y OR2X1_LOC_742/a_8_216# 0.14fF
C1580 OR2X1_LOC_696/A AND2X1_LOC_844/a_8_24# 0.01fF
C1581 AND2X1_LOC_504/a_8_24# OR2X1_LOC_507/A 0.20fF
C1582 OR2X1_LOC_49/A OR2X1_LOC_83/A 0.03fF
C1583 AND2X1_LOC_785/a_8_24# OR2X1_LOC_70/Y 0.04fF
C1584 OR2X1_LOC_216/Y AND2X1_LOC_65/A 0.40fF
C1585 AND2X1_LOC_86/Y OR2X1_LOC_66/A 0.01fF
C1586 OR2X1_LOC_135/Y OR2X1_LOC_43/A 0.03fF
C1587 OR2X1_LOC_604/A AND2X1_LOC_452/Y 1.12fF
C1588 OR2X1_LOC_379/Y VDD 0.14fF
C1589 OR2X1_LOC_114/B OR2X1_LOC_347/B 0.03fF
C1590 OR2X1_LOC_244/B OR2X1_LOC_244/a_36_216# 0.00fF
C1591 OR2X1_LOC_155/A OR2X1_LOC_161/B 0.15fF
C1592 OR2X1_LOC_61/Y OR2X1_LOC_78/A 0.46fF
C1593 OR2X1_LOC_158/A AND2X1_LOC_35/a_36_24# 0.01fF
C1594 INPUT_3 OR2X1_LOC_66/A 0.50fF
C1595 AND2X1_LOC_91/B OR2X1_LOC_705/Y 0.00fF
C1596 OR2X1_LOC_158/A OR2X1_LOC_6/A 1.94fF
C1597 OR2X1_LOC_382/A OR2X1_LOC_44/Y 0.00fF
C1598 AND2X1_LOC_564/A AND2X1_LOC_711/Y 9.83fF
C1599 AND2X1_LOC_566/a_8_24# AND2X1_LOC_212/Y 0.01fF
C1600 OR2X1_LOC_691/a_36_216# OR2X1_LOC_269/B 0.00fF
C1601 OR2X1_LOC_154/A OR2X1_LOC_362/A 0.07fF
C1602 AND2X1_LOC_564/A OR2X1_LOC_70/Y 0.03fF
C1603 OR2X1_LOC_584/a_8_216# OR2X1_LOC_52/B 0.03fF
C1604 OR2X1_LOC_670/a_8_216# OR2X1_LOC_9/Y 0.12fF
C1605 AND2X1_LOC_539/Y OR2X1_LOC_829/Y 0.02fF
C1606 VDD OR2X1_LOC_316/Y 0.62fF
C1607 OR2X1_LOC_51/Y AND2X1_LOC_621/Y 0.23fF
C1608 AND2X1_LOC_658/B OR2X1_LOC_39/A 1.64fF
C1609 OR2X1_LOC_264/Y OR2X1_LOC_663/A 4.05fF
C1610 AND2X1_LOC_714/B AND2X1_LOC_446/a_8_24# 0.20fF
C1611 AND2X1_LOC_357/B OR2X1_LOC_36/Y 0.01fF
C1612 OR2X1_LOC_553/A OR2X1_LOC_66/A 0.25fF
C1613 OR2X1_LOC_3/Y OR2X1_LOC_12/Y 1.68fF
C1614 AND2X1_LOC_556/a_36_24# OR2X1_LOC_92/Y 0.00fF
C1615 AND2X1_LOC_593/Y OR2X1_LOC_59/Y 0.02fF
C1616 OR2X1_LOC_651/A AND2X1_LOC_36/Y 0.03fF
C1617 VDD OR2X1_LOC_194/Y 0.11fF
C1618 OR2X1_LOC_3/Y OR2X1_LOC_766/Y 0.02fF
C1619 OR2X1_LOC_8/Y OR2X1_LOC_246/Y 0.10fF
C1620 AND2X1_LOC_621/Y AND2X1_LOC_444/a_8_24# 0.03fF
C1621 OR2X1_LOC_273/Y AND2X1_LOC_786/Y 0.03fF
C1622 OR2X1_LOC_51/Y AND2X1_LOC_668/a_8_24# 0.00fF
C1623 OR2X1_LOC_326/B OR2X1_LOC_808/B 0.10fF
C1624 VDD AND2X1_LOC_354/B 0.10fF
C1625 OR2X1_LOC_114/Y VDD 0.12fF
C1626 AND2X1_LOC_520/Y OR2X1_LOC_275/Y 0.00fF
C1627 OR2X1_LOC_756/B AND2X1_LOC_95/Y 2.12fF
C1628 AND2X1_LOC_722/A OR2X1_LOC_48/B 0.04fF
C1629 OR2X1_LOC_89/A OR2X1_LOC_382/a_8_216# 0.01fF
C1630 OR2X1_LOC_814/A OR2X1_LOC_831/B 0.07fF
C1631 OR2X1_LOC_403/B AND2X1_LOC_18/Y 0.01fF
C1632 AND2X1_LOC_95/Y OR2X1_LOC_735/a_36_216# 0.00fF
C1633 OR2X1_LOC_715/B AND2X1_LOC_3/Y 0.47fF
C1634 OR2X1_LOC_864/A OR2X1_LOC_641/a_36_216# 0.00fF
C1635 OR2X1_LOC_809/B OR2X1_LOC_802/Y 0.10fF
C1636 AND2X1_LOC_798/Y AND2X1_LOC_810/B 0.04fF
C1637 OR2X1_LOC_241/Y OR2X1_LOC_130/Y 0.00fF
C1638 AND2X1_LOC_719/Y AND2X1_LOC_719/a_36_24# 0.00fF
C1639 OR2X1_LOC_85/A OR2X1_LOC_59/Y 2.47fF
C1640 OR2X1_LOC_517/A OR2X1_LOC_118/Y 0.03fF
C1641 OR2X1_LOC_656/B OR2X1_LOC_502/A 0.07fF
C1642 OR2X1_LOC_219/B OR2X1_LOC_66/A 0.01fF
C1643 AND2X1_LOC_561/B OR2X1_LOC_26/Y 0.25fF
C1644 AND2X1_LOC_656/Y AND2X1_LOC_772/Y 0.09fF
C1645 OR2X1_LOC_160/A OR2X1_LOC_216/A 0.01fF
C1646 OR2X1_LOC_53/Y AND2X1_LOC_199/a_8_24# 0.01fF
C1647 AND2X1_LOC_366/A AND2X1_LOC_367/a_8_24# 0.01fF
C1648 AND2X1_LOC_512/Y OR2X1_LOC_511/Y 0.10fF
C1649 OR2X1_LOC_319/B AND2X1_LOC_43/B 0.02fF
C1650 AND2X1_LOC_573/A AND2X1_LOC_266/a_8_24# 0.04fF
C1651 AND2X1_LOC_175/B AND2X1_LOC_654/B 0.01fF
C1652 AND2X1_LOC_141/a_36_24# OR2X1_LOC_26/Y 0.01fF
C1653 AND2X1_LOC_340/Y OR2X1_LOC_46/A 0.03fF
C1654 OR2X1_LOC_235/B OR2X1_LOC_845/a_8_216# 0.01fF
C1655 AND2X1_LOC_154/Y AND2X1_LOC_658/a_8_24# 0.03fF
C1656 OR2X1_LOC_702/A OR2X1_LOC_676/Y 0.01fF
C1657 AND2X1_LOC_714/B OR2X1_LOC_417/Y 0.15fF
C1658 AND2X1_LOC_98/Y OR2X1_LOC_6/A 0.03fF
C1659 OR2X1_LOC_778/Y OR2X1_LOC_778/a_8_216# 0.01fF
C1660 OR2X1_LOC_680/A AND2X1_LOC_865/a_8_24# 0.03fF
C1661 OR2X1_LOC_154/A OR2X1_LOC_474/Y 0.10fF
C1662 VDD AND2X1_LOC_390/B 1.08fF
C1663 AND2X1_LOC_570/Y OR2X1_LOC_239/Y 0.01fF
C1664 AND2X1_LOC_561/B OR2X1_LOC_89/A 0.03fF
C1665 OR2X1_LOC_347/a_8_216# OR2X1_LOC_161/A 0.01fF
C1666 OR2X1_LOC_32/B OR2X1_LOC_393/a_8_216# 0.05fF
C1667 OR2X1_LOC_539/A OR2X1_LOC_154/A 0.01fF
C1668 VDD OR2X1_LOC_201/Y 0.12fF
C1669 OR2X1_LOC_53/Y OR2X1_LOC_689/Y 0.01fF
C1670 OR2X1_LOC_499/B OR2X1_LOC_631/B 0.00fF
C1671 OR2X1_LOC_405/A OR2X1_LOC_730/a_36_216# 0.00fF
C1672 OR2X1_LOC_46/A AND2X1_LOC_415/a_36_24# 0.00fF
C1673 AND2X1_LOC_141/a_36_24# OR2X1_LOC_89/A 0.00fF
C1674 INPUT_5 OR2X1_LOC_36/Y 0.01fF
C1675 OR2X1_LOC_405/A OR2X1_LOC_161/A 0.19fF
C1676 OR2X1_LOC_639/B AND2X1_LOC_11/Y 0.22fF
C1677 OR2X1_LOC_140/B D_INPUT_1 0.03fF
C1678 AND2X1_LOC_189/a_8_24# OR2X1_LOC_564/A 0.24fF
C1679 AND2X1_LOC_55/a_8_24# AND2X1_LOC_414/a_8_24# 0.23fF
C1680 OR2X1_LOC_728/B AND2X1_LOC_36/Y 0.01fF
C1681 OR2X1_LOC_697/a_8_216# OR2X1_LOC_7/A -0.04fF
C1682 AND2X1_LOC_318/Y AND2X1_LOC_476/a_8_24# 0.00fF
C1683 OR2X1_LOC_131/Y OR2X1_LOC_744/A 0.49fF
C1684 OR2X1_LOC_739/B OR2X1_LOC_739/A 0.14fF
C1685 AND2X1_LOC_644/Y AND2X1_LOC_648/a_8_24# 0.09fF
C1686 OR2X1_LOC_235/B OR2X1_LOC_485/A 0.09fF
C1687 VDD OR2X1_LOC_431/Y 0.09fF
C1688 OR2X1_LOC_65/B AND2X1_LOC_656/a_36_24# 0.00fF
C1689 AND2X1_LOC_452/Y AND2X1_LOC_467/a_8_24# 0.05fF
C1690 AND2X1_LOC_59/Y OR2X1_LOC_739/A 0.03fF
C1691 OR2X1_LOC_273/a_36_216# AND2X1_LOC_219/Y 0.01fF
C1692 AND2X1_LOC_340/Y AND2X1_LOC_227/Y 0.10fF
C1693 VDD OR2X1_LOC_844/Y 0.05fF
C1694 OR2X1_LOC_810/A OR2X1_LOC_775/a_8_216# 0.05fF
C1695 AND2X1_LOC_851/B AND2X1_LOC_445/a_8_24# 0.04fF
C1696 OR2X1_LOC_315/Y OR2X1_LOC_316/Y 0.05fF
C1697 VDD AND2X1_LOC_101/a_8_24# -0.00fF
C1698 AND2X1_LOC_47/Y OR2X1_LOC_736/Y 0.01fF
C1699 AND2X1_LOC_318/a_36_24# OR2X1_LOC_18/Y 0.00fF
C1700 OR2X1_LOC_75/Y AND2X1_LOC_786/Y 0.01fF
C1701 OR2X1_LOC_680/A AND2X1_LOC_621/Y 0.03fF
C1702 OR2X1_LOC_805/A AND2X1_LOC_43/B 0.22fF
C1703 OR2X1_LOC_599/A OR2X1_LOC_48/B 0.79fF
C1704 OR2X1_LOC_184/Y AND2X1_LOC_456/a_8_24# 0.10fF
C1705 OR2X1_LOC_614/Y AND2X1_LOC_47/Y 0.16fF
C1706 AND2X1_LOC_784/A AND2X1_LOC_168/Y 0.05fF
C1707 AND2X1_LOC_715/A OR2X1_LOC_268/a_8_216# 0.09fF
C1708 AND2X1_LOC_702/a_8_24# OR2X1_LOC_36/Y 0.01fF
C1709 OR2X1_LOC_64/Y AND2X1_LOC_434/Y 0.01fF
C1710 OR2X1_LOC_854/A OR2X1_LOC_319/Y 0.33fF
C1711 OR2X1_LOC_62/A OR2X1_LOC_16/A 0.23fF
C1712 AND2X1_LOC_42/B AND2X1_LOC_819/a_36_24# 0.00fF
C1713 OR2X1_LOC_733/a_8_216# OR2X1_LOC_722/a_8_216# 0.47fF
C1714 OR2X1_LOC_160/A OR2X1_LOC_802/Y 0.03fF
C1715 AND2X1_LOC_727/A AND2X1_LOC_436/Y 0.01fF
C1716 OR2X1_LOC_599/A OR2X1_LOC_18/Y 0.02fF
C1717 AND2X1_LOC_56/B OR2X1_LOC_269/a_36_216# 0.00fF
C1718 AND2X1_LOC_95/Y OR2X1_LOC_76/Y 0.03fF
C1719 AND2X1_LOC_741/Y GATE_811 0.00fF
C1720 AND2X1_LOC_211/B AND2X1_LOC_357/a_8_24# 0.04fF
C1721 OR2X1_LOC_539/Y OR2X1_LOC_802/A 0.01fF
C1722 OR2X1_LOC_864/a_8_216# OR2X1_LOC_772/B 0.01fF
C1723 AND2X1_LOC_164/a_36_24# AND2X1_LOC_51/Y 0.00fF
C1724 OR2X1_LOC_160/A OR2X1_LOC_468/Y 0.00fF
C1725 AND2X1_LOC_833/a_8_24# OR2X1_LOC_238/Y 0.01fF
C1726 AND2X1_LOC_435/a_8_24# OR2X1_LOC_44/Y 0.01fF
C1727 OR2X1_LOC_502/A AND2X1_LOC_612/a_36_24# 0.00fF
C1728 OR2X1_LOC_858/a_36_216# OR2X1_LOC_814/A -0.00fF
C1729 OR2X1_LOC_3/Y OR2X1_LOC_422/a_8_216# 0.00fF
C1730 OR2X1_LOC_31/Y OR2X1_LOC_583/a_8_216# 0.01fF
C1731 AND2X1_LOC_465/Y OR2X1_LOC_56/A 0.00fF
C1732 VDD OR2X1_LOC_286/a_8_216# 0.00fF
C1733 OR2X1_LOC_210/a_8_216# OR2X1_LOC_87/A 0.01fF
C1734 OR2X1_LOC_437/A OR2X1_LOC_142/a_36_216# 0.00fF
C1735 OR2X1_LOC_617/Y AND2X1_LOC_866/B 0.97fF
C1736 OR2X1_LOC_189/a_8_216# AND2X1_LOC_578/A 0.03fF
C1737 OR2X1_LOC_244/A OR2X1_LOC_66/A 0.19fF
C1738 AND2X1_LOC_59/Y OR2X1_LOC_269/B 1.36fF
C1739 VDD AND2X1_LOC_863/Y 0.21fF
C1740 AND2X1_LOC_592/Y AND2X1_LOC_648/B 0.01fF
C1741 AND2X1_LOC_102/a_8_24# OR2X1_LOC_375/A 0.01fF
C1742 AND2X1_LOC_753/B AND2X1_LOC_51/Y 0.00fF
C1743 AND2X1_LOC_70/Y AND2X1_LOC_821/a_8_24# 0.11fF
C1744 OR2X1_LOC_26/Y AND2X1_LOC_266/Y 0.03fF
C1745 OR2X1_LOC_185/Y OR2X1_LOC_643/A 0.05fF
C1746 OR2X1_LOC_865/a_8_216# OR2X1_LOC_269/B 0.00fF
C1747 AND2X1_LOC_808/A AND2X1_LOC_469/Y 0.02fF
C1748 AND2X1_LOC_390/B OR2X1_LOC_829/a_8_216# 0.04fF
C1749 OR2X1_LOC_532/B AND2X1_LOC_92/Y 0.14fF
C1750 OR2X1_LOC_364/A OR2X1_LOC_778/Y 0.10fF
C1751 OR2X1_LOC_95/Y AND2X1_LOC_436/Y 0.02fF
C1752 OR2X1_LOC_426/A OR2X1_LOC_684/Y 0.16fF
C1753 OR2X1_LOC_786/Y AND2X1_LOC_625/a_8_24# 0.03fF
C1754 OR2X1_LOC_694/a_8_216# OR2X1_LOC_3/Y 0.02fF
C1755 AND2X1_LOC_8/Y OR2X1_LOC_99/a_8_216# 0.03fF
C1756 AND2X1_LOC_149/a_8_24# OR2X1_LOC_679/B 0.20fF
C1757 OR2X1_LOC_70/Y AND2X1_LOC_593/Y 0.12fF
C1758 AND2X1_LOC_795/Y AND2X1_LOC_476/Y 0.12fF
C1759 OR2X1_LOC_405/A AND2X1_LOC_51/Y 0.45fF
C1760 OR2X1_LOC_485/A AND2X1_LOC_319/A 0.02fF
C1761 OR2X1_LOC_599/A OR2X1_LOC_385/Y 0.00fF
C1762 AND2X1_LOC_571/a_8_24# AND2X1_LOC_657/A 0.01fF
C1763 OR2X1_LOC_75/a_36_216# AND2X1_LOC_219/Y 0.00fF
C1764 AND2X1_LOC_489/Y AND2X1_LOC_576/Y 0.15fF
C1765 OR2X1_LOC_261/Y OR2X1_LOC_44/Y 0.26fF
C1766 OR2X1_LOC_83/A AND2X1_LOC_612/B 0.23fF
C1767 OR2X1_LOC_661/a_8_216# OR2X1_LOC_476/B 0.02fF
C1768 AND2X1_LOC_472/B OR2X1_LOC_378/Y 0.06fF
C1769 OR2X1_LOC_106/A OR2X1_LOC_585/A 0.03fF
C1770 AND2X1_LOC_578/A AND2X1_LOC_565/Y 0.01fF
C1771 AND2X1_LOC_59/Y AND2X1_LOC_75/a_8_24# 0.11fF
C1772 OR2X1_LOC_8/Y OR2X1_LOC_29/a_8_216# 0.06fF
C1773 VDD OR2X1_LOC_796/B -0.00fF
C1774 OR2X1_LOC_70/Y OR2X1_LOC_85/A 0.35fF
C1775 AND2X1_LOC_371/a_8_24# OR2X1_LOC_493/Y 0.02fF
C1776 OR2X1_LOC_808/B AND2X1_LOC_47/Y 0.02fF
C1777 AND2X1_LOC_7/B OR2X1_LOC_367/B 0.03fF
C1778 OR2X1_LOC_625/Y OR2X1_LOC_22/Y 0.02fF
C1779 OR2X1_LOC_12/Y AND2X1_LOC_772/a_8_24# 0.01fF
C1780 AND2X1_LOC_18/Y OR2X1_LOC_493/Y 0.10fF
C1781 AND2X1_LOC_500/a_36_24# OR2X1_LOC_485/A 0.00fF
C1782 AND2X1_LOC_18/Y OR2X1_LOC_801/B 0.07fF
C1783 VDD OR2X1_LOC_544/a_8_216# 0.21fF
C1784 AND2X1_LOC_36/Y OR2X1_LOC_622/B 0.05fF
C1785 OR2X1_LOC_703/Y OR2X1_LOC_714/a_8_216# 0.06fF
C1786 OR2X1_LOC_592/A OR2X1_LOC_592/a_8_216# 0.47fF
C1787 OR2X1_LOC_647/Y OR2X1_LOC_87/A 0.11fF
C1788 VDD OR2X1_LOC_741/A -0.00fF
C1789 OR2X1_LOC_384/Y OR2X1_LOC_428/A 0.68fF
C1790 AND2X1_LOC_823/a_8_24# AND2X1_LOC_51/Y 0.01fF
C1791 OR2X1_LOC_652/a_8_216# OR2X1_LOC_814/A 0.16fF
C1792 AND2X1_LOC_729/Y AND2X1_LOC_687/Y 0.01fF
C1793 OR2X1_LOC_462/B OR2X1_LOC_650/Y 0.13fF
C1794 OR2X1_LOC_43/A AND2X1_LOC_856/B 0.01fF
C1795 AND2X1_LOC_714/a_8_24# OR2X1_LOC_589/Y 0.01fF
C1796 AND2X1_LOC_724/A OR2X1_LOC_423/Y 0.09fF
C1797 OR2X1_LOC_837/B AND2X1_LOC_476/A 0.07fF
C1798 OR2X1_LOC_837/A AND2X1_LOC_472/a_36_24# 0.00fF
C1799 OR2X1_LOC_3/Y OR2X1_LOC_272/Y 0.11fF
C1800 AND2X1_LOC_48/A OR2X1_LOC_793/A 0.01fF
C1801 OR2X1_LOC_223/A OR2X1_LOC_785/B 0.02fF
C1802 D_INPUT_3 AND2X1_LOC_820/a_8_24# 0.01fF
C1803 AND2X1_LOC_36/Y OR2X1_LOC_338/A 0.07fF
C1804 OR2X1_LOC_18/Y AND2X1_LOC_866/A 0.03fF
C1805 AND2X1_LOC_831/Y AND2X1_LOC_138/a_8_24# 0.01fF
C1806 OR2X1_LOC_764/Y OR2X1_LOC_64/Y 0.02fF
C1807 OR2X1_LOC_687/A AND2X1_LOC_430/B 0.01fF
C1808 AND2X1_LOC_841/a_8_24# AND2X1_LOC_662/B 0.03fF
C1809 AND2X1_LOC_69/a_8_24# OR2X1_LOC_87/A 0.01fF
C1810 OR2X1_LOC_472/B OR2X1_LOC_472/A 0.43fF
C1811 AND2X1_LOC_86/Y OR2X1_LOC_84/A 0.04fF
C1812 OR2X1_LOC_687/Y AND2X1_LOC_53/Y 0.46fF
C1813 OR2X1_LOC_585/A OR2X1_LOC_46/A 0.27fF
C1814 OR2X1_LOC_589/A OR2X1_LOC_536/a_8_216# 0.01fF
C1815 OR2X1_LOC_479/Y OR2X1_LOC_121/B 0.10fF
C1816 OR2X1_LOC_744/A AND2X1_LOC_657/A 0.41fF
C1817 AND2X1_LOC_345/Y OR2X1_LOC_54/Y 0.23fF
C1818 OR2X1_LOC_779/Y OR2X1_LOC_161/A 0.01fF
C1819 OR2X1_LOC_47/Y OR2X1_LOC_39/A 0.19fF
C1820 AND2X1_LOC_123/a_8_24# AND2X1_LOC_845/Y 0.02fF
C1821 OR2X1_LOC_62/B OR2X1_LOC_74/A 0.02fF
C1822 OR2X1_LOC_186/Y AND2X1_LOC_36/Y 0.07fF
C1823 OR2X1_LOC_334/A OR2X1_LOC_338/A 0.09fF
C1824 OR2X1_LOC_56/A OR2X1_LOC_521/a_36_216# 0.01fF
C1825 OR2X1_LOC_472/A OR2X1_LOC_852/A 0.01fF
C1826 OR2X1_LOC_160/A OR2X1_LOC_205/Y 0.09fF
C1827 AND2X1_LOC_716/Y AND2X1_LOC_222/Y 0.00fF
C1828 OR2X1_LOC_78/B OR2X1_LOC_71/A 0.03fF
C1829 OR2X1_LOC_474/Y OR2X1_LOC_560/A 0.03fF
C1830 OR2X1_LOC_726/A AND2X1_LOC_36/Y 0.40fF
C1831 OR2X1_LOC_596/A OR2X1_LOC_714/a_8_216# 0.04fF
C1832 AND2X1_LOC_213/B AND2X1_LOC_209/Y 0.01fF
C1833 OR2X1_LOC_323/A AND2X1_LOC_786/Y 0.04fF
C1834 AND2X1_LOC_476/Y AND2X1_LOC_439/a_8_24# 0.04fF
C1835 OR2X1_LOC_244/Y OR2X1_LOC_777/B 0.05fF
C1836 AND2X1_LOC_48/A AND2X1_LOC_45/a_8_24# 0.01fF
C1837 OR2X1_LOC_417/Y AND2X1_LOC_477/A 0.57fF
C1838 OR2X1_LOC_224/Y OR2X1_LOC_7/A 0.00fF
C1839 AND2X1_LOC_721/A OR2X1_LOC_248/a_36_216# 0.00fF
C1840 OR2X1_LOC_211/a_8_216# OR2X1_LOC_566/a_8_216# 0.47fF
C1841 OR2X1_LOC_175/Y AND2X1_LOC_44/Y 0.05fF
C1842 AND2X1_LOC_362/a_8_24# OR2X1_LOC_13/B 0.03fF
C1843 AND2X1_LOC_211/B OR2X1_LOC_47/Y 0.02fF
C1844 OR2X1_LOC_74/A AND2X1_LOC_796/Y 0.03fF
C1845 OR2X1_LOC_87/A AND2X1_LOC_428/a_8_24# 0.02fF
C1846 OR2X1_LOC_36/Y AND2X1_LOC_204/Y 0.01fF
C1847 OR2X1_LOC_444/B OR2X1_LOC_444/a_8_216# 0.47fF
C1848 OR2X1_LOC_644/B OR2X1_LOC_644/A 0.04fF
C1849 AND2X1_LOC_849/A AND2X1_LOC_845/Y 0.02fF
C1850 OR2X1_LOC_377/A AND2X1_LOC_31/Y 0.07fF
C1851 OR2X1_LOC_405/Y OR2X1_LOC_228/Y 0.01fF
C1852 OR2X1_LOC_212/a_8_216# OR2X1_LOC_357/A 0.40fF
C1853 OR2X1_LOC_833/Y OR2X1_LOC_121/A 0.02fF
C1854 OR2X1_LOC_691/Y AND2X1_LOC_44/Y 0.03fF
C1855 OR2X1_LOC_756/B OR2X1_LOC_788/B 0.00fF
C1856 AND2X1_LOC_461/a_36_24# OR2X1_LOC_690/A 0.02fF
C1857 OR2X1_LOC_522/a_8_216# OR2X1_LOC_428/A 0.01fF
C1858 OR2X1_LOC_114/Y OR2X1_LOC_140/a_8_216# 0.01fF
C1859 OR2X1_LOC_16/A OR2X1_LOC_312/a_36_216# 0.00fF
C1860 OR2X1_LOC_116/A OR2X1_LOC_560/A 0.01fF
C1861 OR2X1_LOC_485/A AND2X1_LOC_721/A 0.02fF
C1862 OR2X1_LOC_655/B OR2X1_LOC_655/A 0.07fF
C1863 OR2X1_LOC_64/Y AND2X1_LOC_851/B 0.06fF
C1864 OR2X1_LOC_516/Y OR2X1_LOC_56/A 0.03fF
C1865 OR2X1_LOC_52/B AND2X1_LOC_784/a_36_24# 0.00fF
C1866 AND2X1_LOC_44/Y OR2X1_LOC_713/A 0.44fF
C1867 AND2X1_LOC_70/Y OR2X1_LOC_605/Y 0.05fF
C1868 OR2X1_LOC_196/Y AND2X1_LOC_754/a_8_24# 0.24fF
C1869 OR2X1_LOC_217/Y OR2X1_LOC_560/A 0.46fF
C1870 AND2X1_LOC_719/Y AND2X1_LOC_287/B 0.00fF
C1871 OR2X1_LOC_485/A AND2X1_LOC_644/a_36_24# 0.00fF
C1872 AND2X1_LOC_719/Y OR2X1_LOC_816/A 0.03fF
C1873 OR2X1_LOC_538/A OR2X1_LOC_319/Y 0.22fF
C1874 AND2X1_LOC_620/Y AND2X1_LOC_624/a_36_24# 0.00fF
C1875 OR2X1_LOC_312/Y AND2X1_LOC_222/Y 0.03fF
C1876 OR2X1_LOC_109/Y OR2X1_LOC_437/A 0.10fF
C1877 OR2X1_LOC_375/A OR2X1_LOC_71/A 0.03fF
C1878 OR2X1_LOC_191/B OR2X1_LOC_742/B 0.06fF
C1879 AND2X1_LOC_51/Y OR2X1_LOC_330/a_8_216# 0.09fF
C1880 OR2X1_LOC_778/Y OR2X1_LOC_568/A 0.10fF
C1881 OR2X1_LOC_317/A OR2X1_LOC_777/B 0.13fF
C1882 AND2X1_LOC_41/A OR2X1_LOC_510/a_8_216# 0.01fF
C1883 AND2X1_LOC_555/Y OR2X1_LOC_59/Y 0.03fF
C1884 AND2X1_LOC_472/B OR2X1_LOC_378/A 0.12fF
C1885 AND2X1_LOC_22/Y OR2X1_LOC_776/Y 0.20fF
C1886 OR2X1_LOC_49/A OR2X1_LOC_6/B 0.21fF
C1887 OR2X1_LOC_76/A OR2X1_LOC_241/B 0.23fF
C1888 OR2X1_LOC_65/a_8_216# AND2X1_LOC_204/Y 0.48fF
C1889 OR2X1_LOC_337/A OR2X1_LOC_182/B 0.02fF
C1890 OR2X1_LOC_595/A OR2X1_LOC_131/a_8_216# 0.01fF
C1891 AND2X1_LOC_56/B AND2X1_LOC_268/a_8_24# 0.01fF
C1892 OR2X1_LOC_473/A D_INPUT_0 0.15fF
C1893 OR2X1_LOC_22/Y OR2X1_LOC_3/B 0.02fF
C1894 AND2X1_LOC_851/B OR2X1_LOC_417/A 0.53fF
C1895 AND2X1_LOC_542/a_8_24# AND2X1_LOC_476/Y 0.01fF
C1896 OR2X1_LOC_244/A OR2X1_LOC_84/A 0.04fF
C1897 OR2X1_LOC_600/A AND2X1_LOC_219/A 0.07fF
C1898 VDD AND2X1_LOC_639/B 0.06fF
C1899 OR2X1_LOC_43/Y OR2X1_LOC_600/A 0.08fF
C1900 OR2X1_LOC_853/a_8_216# OR2X1_LOC_35/Y 0.03fF
C1901 OR2X1_LOC_188/Y AND2X1_LOC_498/a_8_24# 0.00fF
C1902 OR2X1_LOC_596/A OR2X1_LOC_596/a_8_216# 0.13fF
C1903 AND2X1_LOC_544/Y AND2X1_LOC_545/a_8_24# 0.04fF
C1904 AND2X1_LOC_725/a_36_24# OR2X1_LOC_12/Y 0.00fF
C1905 OR2X1_LOC_161/A AND2X1_LOC_246/a_36_24# 0.01fF
C1906 OR2X1_LOC_76/Y OR2X1_LOC_269/A 0.21fF
C1907 AND2X1_LOC_658/B AND2X1_LOC_727/B 0.06fF
C1908 OR2X1_LOC_691/B OR2X1_LOC_66/A 0.01fF
C1909 OR2X1_LOC_124/A AND2X1_LOC_44/Y 0.05fF
C1910 OR2X1_LOC_235/B OR2X1_LOC_267/Y 0.00fF
C1911 OR2X1_LOC_8/Y OR2X1_LOC_16/A 0.08fF
C1912 AND2X1_LOC_515/a_8_24# OR2X1_LOC_600/A 0.01fF
C1913 OR2X1_LOC_184/Y OR2X1_LOC_226/Y 0.00fF
C1914 VDD OR2X1_LOC_604/Y 0.06fF
C1915 OR2X1_LOC_154/A OR2X1_LOC_771/B 0.14fF
C1916 AND2X1_LOC_391/Y OR2X1_LOC_428/A 0.01fF
C1917 AND2X1_LOC_712/Y AND2X1_LOC_713/Y 0.08fF
C1918 OR2X1_LOC_91/A OR2X1_LOC_428/A 2.36fF
C1919 OR2X1_LOC_62/B AND2X1_LOC_647/Y 0.01fF
C1920 OR2X1_LOC_40/Y AND2X1_LOC_357/A 0.09fF
C1921 AND2X1_LOC_22/Y OR2X1_LOC_756/B 0.08fF
C1922 AND2X1_LOC_64/Y OR2X1_LOC_509/A 0.01fF
C1923 OR2X1_LOC_316/Y AND2X1_LOC_269/a_8_24# 0.01fF
C1924 OR2X1_LOC_47/Y OR2X1_LOC_760/a_8_216# 0.01fF
C1925 OR2X1_LOC_155/A OR2X1_LOC_707/a_8_216# 0.01fF
C1926 AND2X1_LOC_866/A AND2X1_LOC_620/Y 0.01fF
C1927 OR2X1_LOC_738/A OR2X1_LOC_727/a_8_216# 0.01fF
C1928 AND2X1_LOC_150/a_8_24# OR2X1_LOC_244/Y 0.23fF
C1929 OR2X1_LOC_235/B OR2X1_LOC_633/A 0.08fF
C1930 OR2X1_LOC_91/A OR2X1_LOC_595/A 0.07fF
C1931 OR2X1_LOC_121/B OR2X1_LOC_68/B 0.06fF
C1932 OR2X1_LOC_223/A OR2X1_LOC_786/Y 0.00fF
C1933 VDD OR2X1_LOC_309/Y 0.12fF
C1934 OR2X1_LOC_417/A OR2X1_LOC_595/Y 0.02fF
C1935 AND2X1_LOC_229/a_36_24# AND2X1_LOC_41/A 0.01fF
C1936 OR2X1_LOC_154/A OR2X1_LOC_776/A 0.00fF
C1937 AND2X1_LOC_95/Y OR2X1_LOC_140/B 0.01fF
C1938 OR2X1_LOC_114/B AND2X1_LOC_184/a_8_24# 0.01fF
C1939 AND2X1_LOC_794/B OR2X1_LOC_744/A 0.03fF
C1940 OR2X1_LOC_174/A OR2X1_LOC_390/A 0.03fF
C1941 AND2X1_LOC_721/A OR2X1_LOC_10/a_8_216# 0.19fF
C1942 OR2X1_LOC_324/B OR2X1_LOC_151/A 0.05fF
C1943 AND2X1_LOC_706/Y AND2X1_LOC_605/Y 0.23fF
C1944 OR2X1_LOC_139/A OR2X1_LOC_175/B 0.27fF
C1945 OR2X1_LOC_610/a_8_216# AND2X1_LOC_7/B 0.16fF
C1946 OR2X1_LOC_235/B OR2X1_LOC_673/a_8_216# 0.02fF
C1947 OR2X1_LOC_621/A AND2X1_LOC_616/a_36_24# 0.01fF
C1948 AND2X1_LOC_41/A AND2X1_LOC_65/A 0.07fF
C1949 AND2X1_LOC_810/Y AND2X1_LOC_486/a_8_24# 0.03fF
C1950 D_INPUT_0 OR2X1_LOC_228/Y 0.02fF
C1951 OR2X1_LOC_600/A AND2X1_LOC_658/A 0.12fF
C1952 AND2X1_LOC_26/a_8_24# AND2X1_LOC_762/a_8_24# 0.23fF
C1953 OR2X1_LOC_47/Y AND2X1_LOC_781/Y 0.10fF
C1954 AND2X1_LOC_728/Y AND2X1_LOC_544/Y 0.03fF
C1955 AND2X1_LOC_507/a_8_24# OR2X1_LOC_56/A 0.09fF
C1956 AND2X1_LOC_717/B OR2X1_LOC_183/a_8_216# 0.00fF
C1957 OR2X1_LOC_756/B OR2X1_LOC_621/A 0.07fF
C1958 OR2X1_LOC_186/Y OR2X1_LOC_325/a_8_216# 0.10fF
C1959 AND2X1_LOC_865/A AND2X1_LOC_807/B 0.24fF
C1960 VDD OR2X1_LOC_744/A 1.19fF
C1961 OR2X1_LOC_510/A AND2X1_LOC_41/A 0.06fF
C1962 OR2X1_LOC_643/A OR2X1_LOC_510/a_36_216# 0.01fF
C1963 AND2X1_LOC_756/a_36_24# OR2X1_LOC_600/A 0.00fF
C1964 OR2X1_LOC_147/B OR2X1_LOC_344/A 0.03fF
C1965 AND2X1_LOC_699/a_36_24# AND2X1_LOC_44/Y -0.02fF
C1966 OR2X1_LOC_774/B D_INPUT_1 0.01fF
C1967 OR2X1_LOC_40/Y AND2X1_LOC_508/A 0.02fF
C1968 AND2X1_LOC_76/Y OR2X1_LOC_16/A 0.02fF
C1969 OR2X1_LOC_364/A AND2X1_LOC_91/B 0.08fF
C1970 OR2X1_LOC_51/Y OR2X1_LOC_59/Y 4.85fF
C1971 OR2X1_LOC_40/Y AND2X1_LOC_303/a_36_24# 0.00fF
C1972 OR2X1_LOC_252/Y OR2X1_LOC_816/A 0.00fF
C1973 OR2X1_LOC_185/Y AND2X1_LOC_91/B 0.10fF
C1974 OR2X1_LOC_151/A AND2X1_LOC_142/a_8_24# 0.04fF
C1975 OR2X1_LOC_456/Y AND2X1_LOC_7/B 0.16fF
C1976 AND2X1_LOC_555/Y OR2X1_LOC_820/B 0.03fF
C1977 OR2X1_LOC_773/B AND2X1_LOC_488/a_8_24# 0.20fF
C1978 OR2X1_LOC_158/A AND2X1_LOC_155/a_36_24# 0.00fF
C1979 OR2X1_LOC_53/Y OR2X1_LOC_36/Y 0.06fF
C1980 AND2X1_LOC_793/Y AND2X1_LOC_805/a_8_24# 0.05fF
C1981 OR2X1_LOC_551/B OR2X1_LOC_545/a_8_216# 0.01fF
C1982 AND2X1_LOC_573/A OR2X1_LOC_595/A 0.09fF
C1983 OR2X1_LOC_505/a_36_216# OR2X1_LOC_39/A 0.00fF
C1984 OR2X1_LOC_151/A AND2X1_LOC_314/a_8_24# 0.03fF
C1985 OR2X1_LOC_92/Y AND2X1_LOC_614/a_8_24# 0.01fF
C1986 OR2X1_LOC_78/A OR2X1_LOC_630/B 0.03fF
C1987 OR2X1_LOC_774/Y OR2X1_LOC_773/Y 0.74fF
C1988 OR2X1_LOC_538/a_8_216# AND2X1_LOC_70/Y 0.01fF
C1989 AND2X1_LOC_283/a_8_24# OR2X1_LOC_580/A 0.04fF
C1990 AND2X1_LOC_364/Y INPUT_0 0.03fF
C1991 OR2X1_LOC_61/B AND2X1_LOC_18/Y 0.03fF
C1992 OR2X1_LOC_464/A OR2X1_LOC_741/Y 0.54fF
C1993 AND2X1_LOC_658/A AND2X1_LOC_862/Y 0.21fF
C1994 D_INPUT_1 OR2X1_LOC_557/a_8_216# 0.01fF
C1995 OR2X1_LOC_506/Y AND2X1_LOC_81/B 0.01fF
C1996 OR2X1_LOC_40/Y OR2X1_LOC_48/B 6.64fF
C1997 OR2X1_LOC_114/B OR2X1_LOC_811/A 0.03fF
C1998 OR2X1_LOC_207/B OR2X1_LOC_793/A 0.02fF
C1999 OR2X1_LOC_810/A AND2X1_LOC_7/B 3.52fF
C2000 OR2X1_LOC_196/B AND2X1_LOC_36/Y 0.03fF
C2001 AND2X1_LOC_719/Y AND2X1_LOC_843/a_8_24# 0.02fF
C2002 OR2X1_LOC_323/A AND2X1_LOC_578/A 0.03fF
C2003 AND2X1_LOC_362/B AND2X1_LOC_572/Y 0.10fF
C2004 OR2X1_LOC_744/A OR2X1_LOC_677/Y 0.03fF
C2005 OR2X1_LOC_406/Y OR2X1_LOC_189/Y 0.03fF
C2006 AND2X1_LOC_84/Y OR2X1_LOC_74/A 0.03fF
C2007 OR2X1_LOC_40/Y OR2X1_LOC_18/Y 1.17fF
C2008 OR2X1_LOC_310/Y AND2X1_LOC_335/a_8_24# 0.01fF
C2009 AND2X1_LOC_749/a_8_24# OR2X1_LOC_78/B 0.01fF
C2010 OR2X1_LOC_575/A OR2X1_LOC_244/Y 0.02fF
C2011 OR2X1_LOC_194/B AND2X1_LOC_18/Y 0.10fF
C2012 OR2X1_LOC_427/A AND2X1_LOC_657/Y 0.06fF
C2013 OR2X1_LOC_92/Y OR2X1_LOC_597/a_8_216# 0.03fF
C2014 AND2X1_LOC_95/Y OR2X1_LOC_370/a_8_216# 0.02fF
C2015 OR2X1_LOC_600/A AND2X1_LOC_847/Y 0.01fF
C2016 AND2X1_LOC_794/B AND2X1_LOC_840/B 0.10fF
C2017 AND2X1_LOC_705/Y OR2X1_LOC_26/Y 0.03fF
C2018 OR2X1_LOC_16/A OR2X1_LOC_52/B 0.21fF
C2019 AND2X1_LOC_191/B OR2X1_LOC_427/A 0.03fF
C2020 AND2X1_LOC_56/B OR2X1_LOC_729/a_8_216# 0.03fF
C2021 VDD OR2X1_LOC_1/a_8_216# 0.21fF
C2022 OR2X1_LOC_441/a_8_216# OR2X1_LOC_441/Y 0.01fF
C2023 VDD OR2X1_LOC_541/B 0.30fF
C2024 OR2X1_LOC_801/B OR2X1_LOC_789/A 1.08fF
C2025 OR2X1_LOC_158/A OR2X1_LOC_44/Y 1.17fF
C2026 OR2X1_LOC_501/B OR2X1_LOC_575/A 0.07fF
C2027 OR2X1_LOC_427/A AND2X1_LOC_469/B 0.03fF
C2028 OR2X1_LOC_797/B OR2X1_LOC_87/A 0.02fF
C2029 AND2X1_LOC_716/Y AND2X1_LOC_367/A 0.03fF
C2030 AND2X1_LOC_658/A OR2X1_LOC_619/Y 0.03fF
C2031 OR2X1_LOC_158/A AND2X1_LOC_288/a_8_24# 0.01fF
C2032 OR2X1_LOC_114/Y OR2X1_LOC_361/a_36_216# 0.00fF
C2033 OR2X1_LOC_348/Y OR2X1_LOC_805/A 0.07fF
C2034 OR2X1_LOC_62/B AND2X1_LOC_235/a_8_24# 0.01fF
C2035 OR2X1_LOC_781/B OR2X1_LOC_781/a_8_216# 0.01fF
C2036 OR2X1_LOC_406/Y OR2X1_LOC_527/Y 0.18fF
C2037 AND2X1_LOC_705/Y OR2X1_LOC_89/A 0.02fF
C2038 OR2X1_LOC_6/B OR2X1_LOC_87/B 0.10fF
C2039 AND2X1_LOC_82/Y AND2X1_LOC_490/a_8_24# 0.01fF
C2040 OR2X1_LOC_190/A OR2X1_LOC_553/A 0.07fF
C2041 AND2X1_LOC_365/a_8_24# AND2X1_LOC_661/a_8_24# 0.23fF
C2042 OR2X1_LOC_223/A OR2X1_LOC_181/Y 0.01fF
C2043 AND2X1_LOC_47/Y OR2X1_LOC_500/a_8_216# 0.05fF
C2044 OR2X1_LOC_604/A OR2X1_LOC_236/a_36_216# 0.01fF
C2045 OR2X1_LOC_188/Y OR2X1_LOC_76/A 0.04fF
C2046 AND2X1_LOC_576/a_8_24# AND2X1_LOC_561/B 0.01fF
C2047 OR2X1_LOC_757/A AND2X1_LOC_621/Y 0.03fF
C2048 AND2X1_LOC_121/a_8_24# OR2X1_LOC_67/A 0.21fF
C2049 OR2X1_LOC_426/B OR2X1_LOC_67/a_8_216# 0.01fF
C2050 OR2X1_LOC_506/B AND2X1_LOC_239/a_8_24# 0.01fF
C2051 OR2X1_LOC_261/Y OR2X1_LOC_382/A 0.01fF
C2052 VDD AND2X1_LOC_840/B 1.59fF
C2053 OR2X1_LOC_502/A OR2X1_LOC_785/B 0.01fF
C2054 OR2X1_LOC_147/B OR2X1_LOC_254/A 0.10fF
C2055 OR2X1_LOC_858/A OR2X1_LOC_375/A 0.02fF
C2056 OR2X1_LOC_47/Y AND2X1_LOC_247/a_36_24# 0.00fF
C2057 OR2X1_LOC_358/a_8_216# OR2X1_LOC_648/A 0.03fF
C2058 OR2X1_LOC_364/A OR2X1_LOC_645/a_8_216# 0.01fF
C2059 AND2X1_LOC_533/a_8_24# OR2X1_LOC_538/A 0.00fF
C2060 OR2X1_LOC_680/A OR2X1_LOC_59/Y 0.11fF
C2061 AND2X1_LOC_475/a_36_24# AND2X1_LOC_475/Y 0.00fF
C2062 OR2X1_LOC_158/A AND2X1_LOC_116/Y 0.09fF
C2063 OR2X1_LOC_585/A INPUT_2 0.08fF
C2064 AND2X1_LOC_12/Y OR2X1_LOC_678/Y 0.01fF
C2065 VDD OR2X1_LOC_849/A 0.12fF
C2066 INPUT_1 OR2X1_LOC_748/Y 0.01fF
C2067 OR2X1_LOC_40/Y OR2X1_LOC_385/Y 0.03fF
C2068 OR2X1_LOC_6/B AND2X1_LOC_85/a_8_24# 0.14fF
C2069 AND2X1_LOC_474/A AND2X1_LOC_124/a_8_24# 0.01fF
C2070 AND2X1_LOC_535/Y AND2X1_LOC_356/B 0.01fF
C2071 OR2X1_LOC_516/A AND2X1_LOC_477/a_8_24# 0.01fF
C2072 AND2X1_LOC_99/A OR2X1_LOC_92/Y 0.08fF
C2073 OR2X1_LOC_50/a_8_216# D_INPUT_6 0.01fF
C2074 OR2X1_LOC_223/A OR2X1_LOC_301/a_36_216# 0.00fF
C2075 AND2X1_LOC_47/Y OR2X1_LOC_120/a_8_216# 0.04fF
C2076 OR2X1_LOC_318/B OR2X1_LOC_777/B 0.03fF
C2077 OR2X1_LOC_502/A OR2X1_LOC_459/B 0.01fF
C2078 OR2X1_LOC_744/A OR2X1_LOC_491/Y 0.01fF
C2079 OR2X1_LOC_323/A AND2X1_LOC_841/a_8_24# 0.08fF
C2080 OR2X1_LOC_287/B OR2X1_LOC_862/B 0.00fF
C2081 AND2X1_LOC_65/a_8_24# OR2X1_LOC_87/A 0.05fF
C2082 OR2X1_LOC_448/Y OR2X1_LOC_712/a_8_216# 0.03fF
C2083 AND2X1_LOC_566/B AND2X1_LOC_326/A 0.02fF
C2084 AND2X1_LOC_719/Y OR2X1_LOC_488/Y 0.07fF
C2085 OR2X1_LOC_101/a_36_216# OR2X1_LOC_656/B 0.00fF
C2086 AND2X1_LOC_367/B OR2X1_LOC_7/A 0.02fF
C2087 OR2X1_LOC_814/A OR2X1_LOC_161/B 0.03fF
C2088 AND2X1_LOC_843/Y OR2X1_LOC_18/Y 0.03fF
C2089 AND2X1_LOC_802/B AND2X1_LOC_170/B 0.07fF
C2090 OR2X1_LOC_48/B AND2X1_LOC_644/Y 0.02fF
C2091 D_GATE_741 OR2X1_LOC_564/B 0.02fF
C2092 AND2X1_LOC_12/Y OR2X1_LOC_811/A 0.04fF
C2093 AND2X1_LOC_861/B AND2X1_LOC_806/A 0.01fF
C2094 OR2X1_LOC_590/a_8_216# OR2X1_LOC_593/B 0.02fF
C2095 OR2X1_LOC_687/Y OR2X1_LOC_502/A 0.07fF
C2096 AND2X1_LOC_736/Y AND2X1_LOC_580/A 0.29fF
C2097 OR2X1_LOC_18/Y AND2X1_LOC_644/Y 0.05fF
C2098 OR2X1_LOC_424/a_8_216# OR2X1_LOC_48/B 0.04fF
C2099 OR2X1_LOC_459/A AND2X1_LOC_688/a_8_24# 0.20fF
C2100 OR2X1_LOC_476/B OR2X1_LOC_661/A 0.02fF
C2101 OR2X1_LOC_103/Y OR2X1_LOC_44/Y 0.03fF
C2102 OR2X1_LOC_834/a_8_216# OR2X1_LOC_449/B 0.05fF
C2103 D_INPUT_4 AND2X1_LOC_25/Y 0.01fF
C2104 AND2X1_LOC_289/a_36_24# OR2X1_LOC_333/A 0.00fF
C2105 AND2X1_LOC_99/A OR2X1_LOC_65/B 0.06fF
C2106 OR2X1_LOC_70/Y OR2X1_LOC_51/Y 0.93fF
C2107 AND2X1_LOC_70/Y OR2X1_LOC_602/a_8_216# 0.01fF
C2108 OR2X1_LOC_618/a_8_216# AND2X1_LOC_852/B 0.01fF
C2109 AND2X1_LOC_731/a_8_24# OR2X1_LOC_47/Y 0.04fF
C2110 OR2X1_LOC_527/Y OR2X1_LOC_496/a_8_216# 0.03fF
C2111 OR2X1_LOC_49/A AND2X1_LOC_47/Y 0.10fF
C2112 OR2X1_LOC_379/a_8_216# AND2X1_LOC_95/Y 0.02fF
C2113 AND2X1_LOC_42/B OR2X1_LOC_573/a_8_216# 0.01fF
C2114 OR2X1_LOC_433/Y AND2X1_LOC_436/B 0.01fF
C2115 AND2X1_LOC_508/A OR2X1_LOC_7/A 0.00fF
C2116 OR2X1_LOC_91/A AND2X1_LOC_211/a_8_24# 0.09fF
C2117 AND2X1_LOC_553/A OR2X1_LOC_26/Y 0.03fF
C2118 OR2X1_LOC_623/B OR2X1_LOC_269/B 0.01fF
C2119 AND2X1_LOC_717/Y OR2X1_LOC_372/Y 0.81fF
C2120 OR2X1_LOC_545/A OR2X1_LOC_545/B 0.16fF
C2121 AND2X1_LOC_564/A OR2X1_LOC_47/Y 0.06fF
C2122 OR2X1_LOC_231/A OR2X1_LOC_87/A 0.14fF
C2123 AND2X1_LOC_535/Y OR2X1_LOC_22/Y 0.03fF
C2124 AND2X1_LOC_773/Y AND2X1_LOC_476/A 0.10fF
C2125 OR2X1_LOC_532/B OR2X1_LOC_741/a_36_216# 0.02fF
C2126 OR2X1_LOC_837/A AND2X1_LOC_472/B 0.01fF
C2127 OR2X1_LOC_517/A AND2X1_LOC_105/a_36_24# 0.00fF
C2128 AND2X1_LOC_333/a_8_24# OR2X1_LOC_51/Y 0.01fF
C2129 AND2X1_LOC_559/a_8_24# AND2X1_LOC_76/Y 0.01fF
C2130 AND2X1_LOC_570/Y AND2X1_LOC_842/B 0.02fF
C2131 OR2X1_LOC_600/A AND2X1_LOC_814/a_8_24# 0.07fF
C2132 OR2X1_LOC_641/a_8_216# AND2X1_LOC_48/A 0.01fF
C2133 OR2X1_LOC_154/A OR2X1_LOC_402/Y 0.01fF
C2134 AND2X1_LOC_40/Y OR2X1_LOC_564/A 0.02fF
C2135 OR2X1_LOC_405/A OR2X1_LOC_216/Y 0.85fF
C2136 AND2X1_LOC_514/Y OR2X1_LOC_51/Y 0.02fF
C2137 AND2X1_LOC_47/Y OR2X1_LOC_596/A 0.04fF
C2138 AND2X1_LOC_553/A OR2X1_LOC_89/A 0.00fF
C2139 AND2X1_LOC_723/Y AND2X1_LOC_578/A 0.07fF
C2140 OR2X1_LOC_426/B AND2X1_LOC_537/Y 0.07fF
C2141 AND2X1_LOC_363/a_8_24# AND2X1_LOC_866/A 0.17fF
C2142 OR2X1_LOC_689/a_36_216# OR2X1_LOC_585/A 0.00fF
C2143 AND2X1_LOC_840/a_8_24# OR2X1_LOC_89/A 0.02fF
C2144 AND2X1_LOC_638/Y AND2X1_LOC_651/B 0.01fF
C2145 AND2X1_LOC_145/a_36_24# OR2X1_LOC_375/A 0.01fF
C2146 OR2X1_LOC_377/A OR2X1_LOC_461/A 0.70fF
C2147 OR2X1_LOC_841/a_8_216# OR2X1_LOC_479/Y 0.09fF
C2148 AND2X1_LOC_789/a_8_24# OR2X1_LOC_3/Y 0.01fF
C2149 OR2X1_LOC_87/A OR2X1_LOC_340/Y 0.02fF
C2150 AND2X1_LOC_716/Y OR2X1_LOC_74/A 0.65fF
C2151 AND2X1_LOC_364/Y OR2X1_LOC_64/Y 0.03fF
C2152 AND2X1_LOC_857/a_8_24# OR2X1_LOC_48/B 0.12fF
C2153 OR2X1_LOC_3/Y AND2X1_LOC_404/A 0.01fF
C2154 OR2X1_LOC_250/a_8_216# OR2X1_LOC_585/A 0.15fF
C2155 AND2X1_LOC_719/Y OR2X1_LOC_95/Y 0.14fF
C2156 OR2X1_LOC_680/Y AND2X1_LOC_147/a_8_24# 0.01fF
C2157 OR2X1_LOC_87/A OR2X1_LOC_707/A 0.05fF
C2158 OR2X1_LOC_831/B OR2X1_LOC_318/B 0.35fF
C2159 OR2X1_LOC_89/A AND2X1_LOC_804/Y 0.03fF
C2160 OR2X1_LOC_864/A OR2X1_LOC_377/A 0.12fF
C2161 OR2X1_LOC_458/a_8_216# OR2X1_LOC_675/A 0.49fF
C2162 OR2X1_LOC_7/A OR2X1_LOC_48/B 0.91fF
C2163 OR2X1_LOC_18/Y AND2X1_LOC_857/a_8_24# 0.01fF
C2164 OR2X1_LOC_87/A OR2X1_LOC_130/A 1.12fF
C2165 AND2X1_LOC_34/Y AND2X1_LOC_472/B 0.14fF
C2166 AND2X1_LOC_316/a_8_24# AND2X1_LOC_51/Y 0.01fF
C2167 OR2X1_LOC_656/B AND2X1_LOC_3/Y 1.15fF
C2168 OR2X1_LOC_18/Y OR2X1_LOC_7/A 0.31fF
C2169 OR2X1_LOC_124/A OR2X1_LOC_720/B 0.09fF
C2170 OR2X1_LOC_377/A OR2X1_LOC_240/A 7.16fF
C2171 OR2X1_LOC_504/Y OR2X1_LOC_51/Y 0.04fF
C2172 VDD OR2X1_LOC_31/Y 1.18fF
C2173 OR2X1_LOC_810/A OR2X1_LOC_805/A 0.15fF
C2174 OR2X1_LOC_26/Y OR2X1_LOC_511/Y 0.34fF
C2175 OR2X1_LOC_377/A OR2X1_LOC_633/B 0.04fF
C2176 OR2X1_LOC_235/B AND2X1_LOC_107/a_8_24# 0.01fF
C2177 OR2X1_LOC_604/A OR2X1_LOC_96/a_8_216# 0.47fF
C2178 D_INPUT_4 AND2X1_LOC_51/Y 0.02fF
C2179 AND2X1_LOC_705/Y OR2X1_LOC_419/a_8_216# 0.05fF
C2180 AND2X1_LOC_767/a_8_24# AND2X1_LOC_3/Y 0.04fF
C2181 AND2X1_LOC_729/B OR2X1_LOC_761/Y 0.00fF
C2182 AND2X1_LOC_339/B OR2X1_LOC_289/Y 0.04fF
C2183 VDD OR2X1_LOC_440/A 0.10fF
C2184 OR2X1_LOC_87/A AND2X1_LOC_7/a_8_24# 0.17fF
C2185 OR2X1_LOC_160/A AND2X1_LOC_86/B 0.01fF
C2186 AND2X1_LOC_41/A AND2X1_LOC_23/a_8_24# 0.04fF
C2187 AND2X1_LOC_70/Y OR2X1_LOC_439/a_8_216# 0.01fF
C2188 AND2X1_LOC_824/B OR2X1_LOC_240/A 0.02fF
C2189 OR2X1_LOC_49/A OR2X1_LOC_598/A 0.03fF
C2190 AND2X1_LOC_91/B OR2X1_LOC_568/A 0.07fF
C2191 AND2X1_LOC_857/Y OR2X1_LOC_46/A 0.03fF
C2192 OR2X1_LOC_435/B OR2X1_LOC_814/A 0.10fF
C2193 OR2X1_LOC_821/Y OR2X1_LOC_86/A 0.01fF
C2194 OR2X1_LOC_511/Y OR2X1_LOC_89/A 0.02fF
C2195 AND2X1_LOC_559/a_8_24# OR2X1_LOC_52/B 0.02fF
C2196 AND2X1_LOC_548/a_8_24# OR2X1_LOC_39/A 0.01fF
C2197 OR2X1_LOC_137/a_36_216# OR2X1_LOC_720/B 0.00fF
C2198 OR2X1_LOC_744/A OR2X1_LOC_256/A 0.03fF
C2199 OR2X1_LOC_40/Y AND2X1_LOC_620/Y 0.06fF
C2200 OR2X1_LOC_599/A OR2X1_LOC_585/A 0.01fF
C2201 OR2X1_LOC_614/Y AND2X1_LOC_48/Y 0.01fF
C2202 OR2X1_LOC_426/A AND2X1_LOC_639/A 0.13fF
C2203 AND2X1_LOC_59/Y AND2X1_LOC_176/a_8_24# 0.02fF
C2204 OR2X1_LOC_865/A OR2X1_LOC_561/B 0.10fF
C2205 OR2X1_LOC_793/A AND2X1_LOC_3/Y 1.81fF
C2206 OR2X1_LOC_756/B OR2X1_LOC_434/A 0.01fF
C2207 AND2X1_LOC_711/Y OR2X1_LOC_680/A 0.00fF
C2208 AND2X1_LOC_576/Y OR2X1_LOC_280/Y 0.07fF
C2209 OR2X1_LOC_305/a_8_216# OR2X1_LOC_743/A 0.05fF
C2210 OR2X1_LOC_70/Y OR2X1_LOC_680/A 0.11fF
C2211 OR2X1_LOC_160/B OR2X1_LOC_214/B 0.03fF
C2212 AND2X1_LOC_56/B AND2X1_LOC_42/B 0.05fF
C2213 AND2X1_LOC_43/a_8_24# OR2X1_LOC_269/B 0.00fF
C2214 OR2X1_LOC_61/Y OR2X1_LOC_814/A 0.00fF
C2215 OR2X1_LOC_97/A OR2X1_LOC_364/Y 0.01fF
C2216 OR2X1_LOC_659/B AND2X1_LOC_42/B 0.01fF
C2217 OR2X1_LOC_160/B OR2X1_LOC_241/B 0.92fF
C2218 OR2X1_LOC_11/Y OR2X1_LOC_762/a_8_216# 0.02fF
C2219 AND2X1_LOC_208/B OR2X1_LOC_31/Y 0.00fF
C2220 VDD OR2X1_LOC_257/Y 0.12fF
C2221 AND2X1_LOC_36/Y OR2X1_LOC_727/a_8_216# 0.01fF
C2222 OR2X1_LOC_385/Y OR2X1_LOC_7/A 0.68fF
C2223 AND2X1_LOC_8/Y AND2X1_LOC_42/B 0.43fF
C2224 OR2X1_LOC_689/A OR2X1_LOC_31/Y 0.23fF
C2225 OR2X1_LOC_312/Y OR2X1_LOC_74/A 0.03fF
C2226 AND2X1_LOC_474/A OR2X1_LOC_47/Y 0.02fF
C2227 AND2X1_LOC_425/Y OR2X1_LOC_161/A 0.00fF
C2228 OR2X1_LOC_831/A OR2X1_LOC_228/Y 0.04fF
C2229 AND2X1_LOC_727/A AND2X1_LOC_655/A 0.08fF
C2230 OR2X1_LOC_47/Y AND2X1_LOC_240/a_8_24# 0.04fF
C2231 OR2X1_LOC_813/A OR2X1_LOC_71/a_8_216# 0.41fF
C2232 OR2X1_LOC_744/A OR2X1_LOC_67/Y 0.03fF
C2233 OR2X1_LOC_364/a_8_216# OR2X1_LOC_578/B 0.05fF
C2234 AND2X1_LOC_345/Y OR2X1_LOC_89/A 0.03fF
C2235 AND2X1_LOC_389/a_36_24# OR2X1_LOC_585/A 0.00fF
C2236 OR2X1_LOC_598/Y OR2X1_LOC_228/Y 0.03fF
C2237 AND2X1_LOC_86/B OR2X1_LOC_624/B 0.07fF
C2238 INPUT_4 AND2X1_LOC_639/A 0.17fF
C2239 OR2X1_LOC_687/Y AND2X1_LOC_48/A 0.03fF
C2240 OR2X1_LOC_680/A AND2X1_LOC_657/a_8_24# 0.04fF
C2241 OR2X1_LOC_31/Y AND2X1_LOC_274/a_8_24# 0.01fF
C2242 OR2X1_LOC_51/Y OR2X1_LOC_70/A 0.10fF
C2243 AND2X1_LOC_576/Y OR2X1_LOC_22/Y 0.96fF
C2244 AND2X1_LOC_563/a_8_24# OR2X1_LOC_71/Y 0.01fF
C2245 OR2X1_LOC_62/B OR2X1_LOC_87/A 0.03fF
C2246 OR2X1_LOC_851/A OR2X1_LOC_223/A 0.01fF
C2247 OR2X1_LOC_315/Y OR2X1_LOC_31/Y 0.14fF
C2248 OR2X1_LOC_680/A OR2X1_LOC_504/Y 0.03fF
C2249 OR2X1_LOC_146/Y OR2X1_LOC_427/A 0.01fF
C2250 OR2X1_LOC_36/Y INPUT_1 0.22fF
C2251 AND2X1_LOC_339/a_8_24# OR2X1_LOC_416/Y 0.01fF
C2252 OR2X1_LOC_95/Y AND2X1_LOC_655/A 0.02fF
C2253 OR2X1_LOC_614/a_8_216# OR2X1_LOC_375/A 0.05fF
C2254 OR2X1_LOC_827/a_36_216# OR2X1_LOC_46/A 0.00fF
C2255 AND2X1_LOC_640/a_8_24# OR2X1_LOC_26/Y 0.02fF
C2256 INPUT_0 OR2X1_LOC_749/a_8_216# 0.06fF
C2257 AND2X1_LOC_786/Y OR2X1_LOC_142/Y 0.07fF
C2258 OR2X1_LOC_834/A OR2X1_LOC_512/Y 0.01fF
C2259 OR2X1_LOC_472/B AND2X1_LOC_34/a_8_24# 0.23fF
C2260 AND2X1_LOC_687/Y OR2X1_LOC_52/B -0.11fF
C2261 OR2X1_LOC_795/B OR2X1_LOC_228/Y 0.01fF
C2262 OR2X1_LOC_3/Y OR2X1_LOC_278/A 0.01fF
C2263 OR2X1_LOC_56/A AND2X1_LOC_793/B 0.07fF
C2264 D_INPUT_5 OR2X1_LOC_378/a_8_216# 0.02fF
C2265 OR2X1_LOC_87/A OR2X1_LOC_780/B 0.01fF
C2266 AND2X1_LOC_31/Y OR2X1_LOC_78/B 0.35fF
C2267 OR2X1_LOC_316/Y AND2X1_LOC_660/A 0.03fF
C2268 AND2X1_LOC_738/B OR2X1_LOC_533/A 0.02fF
C2269 AND2X1_LOC_537/Y OR2X1_LOC_743/A 0.02fF
C2270 OR2X1_LOC_256/a_8_216# AND2X1_LOC_721/A 0.00fF
C2271 OR2X1_LOC_48/B OR2X1_LOC_511/a_8_216# 0.02fF
C2272 AND2X1_LOC_560/B AND2X1_LOC_660/a_8_24# 0.02fF
C2273 AND2X1_LOC_859/Y AND2X1_LOC_859/B 0.01fF
C2274 OR2X1_LOC_186/Y OR2X1_LOC_469/B 0.12fF
C2275 OR2X1_LOC_64/Y OR2X1_LOC_762/a_8_216# 0.01fF
C2276 OR2X1_LOC_833/Y AND2X1_LOC_36/Y 0.01fF
C2277 AND2X1_LOC_399/a_36_24# AND2X1_LOC_47/Y 0.00fF
C2278 OR2X1_LOC_409/Y OR2X1_LOC_11/Y 0.01fF
C2279 OR2X1_LOC_481/A OR2X1_LOC_295/Y 0.01fF
C2280 AND2X1_LOC_40/Y D_GATE_579 0.01fF
C2281 AND2X1_LOC_753/B AND2X1_LOC_52/Y 0.10fF
C2282 OR2X1_LOC_391/A OR2X1_LOC_561/B 0.02fF
C2283 OR2X1_LOC_599/A AND2X1_LOC_645/a_8_24# 0.00fF
C2284 OR2X1_LOC_114/B OR2X1_LOC_777/B 0.06fF
C2285 OR2X1_LOC_47/Y OR2X1_LOC_85/A 1.67fF
C2286 AND2X1_LOC_151/a_36_24# AND2X1_LOC_810/Y 0.01fF
C2287 AND2X1_LOC_85/a_8_24# AND2X1_LOC_47/Y 0.01fF
C2288 AND2X1_LOC_40/Y OR2X1_LOC_228/Y 0.23fF
C2289 OR2X1_LOC_711/a_8_216# OR2X1_LOC_308/Y 0.04fF
C2290 OR2X1_LOC_726/A OR2X1_LOC_469/B 0.09fF
C2291 OR2X1_LOC_244/Y OR2X1_LOC_735/B 0.02fF
C2292 AND2X1_LOC_499/a_36_24# OR2X1_LOC_142/Y 0.01fF
C2293 INPUT_1 AND2X1_LOC_847/a_36_24# 0.00fF
C2294 OR2X1_LOC_448/a_8_216# AND2X1_LOC_31/Y 0.01fF
C2295 OR2X1_LOC_553/A OR2X1_LOC_241/B 0.15fF
C2296 OR2X1_LOC_66/A AND2X1_LOC_246/a_8_24# 0.02fF
C2297 AND2X1_LOC_95/Y OR2X1_LOC_675/Y 0.03fF
C2298 AND2X1_LOC_705/Y AND2X1_LOC_590/a_8_24# 0.21fF
C2299 AND2X1_LOC_48/A OR2X1_LOC_643/Y 0.00fF
C2300 VDD OR2X1_LOC_320/a_8_216# 0.21fF
C2301 OR2X1_LOC_89/A AND2X1_LOC_648/B 0.10fF
C2302 OR2X1_LOC_703/B OR2X1_LOC_365/B 0.17fF
C2303 OR2X1_LOC_430/a_8_216# OR2X1_LOC_428/Y 0.40fF
C2304 AND2X1_LOC_367/A OR2X1_LOC_13/B 0.08fF
C2305 OR2X1_LOC_7/A AND2X1_LOC_620/Y 0.08fF
C2306 OR2X1_LOC_538/A OR2X1_LOC_777/B 0.03fF
C2307 OR2X1_LOC_87/A OR2X1_LOC_365/B 0.66fF
C2308 OR2X1_LOC_850/B OR2X1_LOC_366/Y 0.02fF
C2309 OR2X1_LOC_65/B OR2X1_LOC_72/Y 0.02fF
C2310 OR2X1_LOC_185/A OR2X1_LOC_80/A 0.15fF
C2311 OR2X1_LOC_375/A AND2X1_LOC_31/Y 0.97fF
C2312 AND2X1_LOC_407/a_8_24# AND2X1_LOC_774/A 0.13fF
C2313 OR2X1_LOC_427/A OR2X1_LOC_164/a_8_216# 0.04fF
C2314 OR2X1_LOC_62/B AND2X1_LOC_15/a_36_24# 0.01fF
C2315 AND2X1_LOC_564/A AND2X1_LOC_469/Y 0.03fF
C2316 OR2X1_LOC_715/B AND2X1_LOC_7/B 0.53fF
C2317 OR2X1_LOC_6/B OR2X1_LOC_392/B 0.10fF
C2318 OR2X1_LOC_45/B OR2X1_LOC_158/A 0.35fF
C2319 AND2X1_LOC_787/A AND2X1_LOC_476/Y 0.02fF
C2320 AND2X1_LOC_626/a_8_24# AND2X1_LOC_7/B 0.04fF
C2321 OR2X1_LOC_691/B OR2X1_LOC_691/a_8_216# 0.07fF
C2322 OR2X1_LOC_53/Y AND2X1_LOC_207/B 0.01fF
C2323 OR2X1_LOC_40/Y OR2X1_LOC_764/a_8_216# 0.09fF
C2324 OR2X1_LOC_49/A OR2X1_LOC_646/B 0.03fF
C2325 AND2X1_LOC_100/a_8_24# OR2X1_LOC_88/Y 0.00fF
C2326 D_INPUT_5 D_INPUT_6 1.12fF
C2327 OR2X1_LOC_188/Y OR2X1_LOC_160/B 0.05fF
C2328 OR2X1_LOC_49/A OR2X1_LOC_672/a_8_216# 0.01fF
C2329 OR2X1_LOC_502/A OR2X1_LOC_199/B 0.02fF
C2330 OR2X1_LOC_808/B OR2X1_LOC_180/B 0.05fF
C2331 AND2X1_LOC_457/a_36_24# AND2X1_LOC_476/Y 0.01fF
C2332 OR2X1_LOC_696/A OR2X1_LOC_235/B 0.79fF
C2333 AND2X1_LOC_47/Y OR2X1_LOC_223/a_8_216# 0.01fF
C2334 OR2X1_LOC_217/a_8_216# OR2X1_LOC_560/A 0.01fF
C2335 AND2X1_LOC_244/A AND2X1_LOC_244/a_8_24# 0.10fF
C2336 AND2X1_LOC_776/Y OR2X1_LOC_329/B 0.48fF
C2337 OR2X1_LOC_379/Y OR2X1_LOC_769/a_36_216# 0.00fF
C2338 OR2X1_LOC_97/A AND2X1_LOC_18/Y 0.04fF
C2339 VDD OR2X1_LOC_572/a_8_216# 0.00fF
C2340 AND2X1_LOC_340/Y OR2X1_LOC_40/Y 0.03fF
C2341 AND2X1_LOC_12/Y OR2X1_LOC_777/B 0.05fF
C2342 AND2X1_LOC_64/Y OR2X1_LOC_235/B 0.11fF
C2343 OR2X1_LOC_158/A OR2X1_LOC_382/A 0.05fF
C2344 OR2X1_LOC_40/Y AND2X1_LOC_810/B 0.42fF
C2345 OR2X1_LOC_364/A OR2X1_LOC_303/B 0.07fF
C2346 OR2X1_LOC_348/Y OR2X1_LOC_580/B 0.10fF
C2347 OR2X1_LOC_161/A OR2X1_LOC_723/B 0.04fF
C2348 VDD AND2X1_LOC_213/B 0.19fF
C2349 OR2X1_LOC_160/A OR2X1_LOC_532/Y 0.03fF
C2350 OR2X1_LOC_566/A OR2X1_LOC_538/A 0.03fF
C2351 OR2X1_LOC_700/Y AND2X1_LOC_789/Y 0.02fF
C2352 AND2X1_LOC_48/A OR2X1_LOC_644/A 0.00fF
C2353 OR2X1_LOC_40/Y AND2X1_LOC_363/a_8_24# 0.01fF
C2354 OR2X1_LOC_6/B OR2X1_LOC_671/Y 0.06fF
C2355 OR2X1_LOC_363/A OR2X1_LOC_366/B 0.27fF
C2356 OR2X1_LOC_421/A AND2X1_LOC_771/B 0.61fF
C2357 OR2X1_LOC_40/Y AND2X1_LOC_181/Y 0.00fF
C2358 OR2X1_LOC_475/Y OR2X1_LOC_228/Y 0.01fF
C2359 OR2X1_LOC_244/Y OR2X1_LOC_161/B 0.01fF
C2360 OR2X1_LOC_196/B OR2X1_LOC_196/a_8_216# 0.07fF
C2361 OR2X1_LOC_426/a_8_216# AND2X1_LOC_451/Y 0.01fF
C2362 AND2X1_LOC_401/Y OR2X1_LOC_397/Y 0.01fF
C2363 OR2X1_LOC_488/a_8_216# AND2X1_LOC_657/A 0.02fF
C2364 OR2X1_LOC_597/A OR2X1_LOC_589/A 0.07fF
C2365 AND2X1_LOC_362/a_8_24# OR2X1_LOC_428/A 0.17fF
C2366 AND2X1_LOC_40/Y OR2X1_LOC_562/A 0.04fF
C2367 OR2X1_LOC_151/A OR2X1_LOC_66/A 0.19fF
C2368 OR2X1_LOC_154/A OR2X1_LOC_593/B 0.00fF
C2369 AND2X1_LOC_91/B OR2X1_LOC_814/a_8_216# 0.02fF
C2370 OR2X1_LOC_501/B OR2X1_LOC_161/B 0.07fF
C2371 OR2X1_LOC_426/B OR2X1_LOC_13/Y 0.03fF
C2372 VDD OR2X1_LOC_129/a_8_216# 0.21fF
C2373 OR2X1_LOC_858/A OR2X1_LOC_549/A 0.02fF
C2374 OR2X1_LOC_95/Y OR2X1_LOC_599/Y 0.25fF
C2375 OR2X1_LOC_630/a_8_216# OR2X1_LOC_140/B 0.01fF
C2376 OR2X1_LOC_516/Y OR2X1_LOC_91/Y 0.42fF
C2377 AND2X1_LOC_47/Y OR2X1_LOC_374/Y 0.25fF
C2378 OR2X1_LOC_186/Y AND2X1_LOC_167/a_8_24# 0.17fF
C2379 OR2X1_LOC_51/Y AND2X1_LOC_499/a_8_24# 0.01fF
C2380 OR2X1_LOC_377/A OR2X1_LOC_397/a_8_216# 0.05fF
C2381 OR2X1_LOC_74/A OR2X1_LOC_13/B 0.21fF
C2382 OR2X1_LOC_850/A OR2X1_LOC_580/A 0.04fF
C2383 OR2X1_LOC_335/A OR2X1_LOC_161/A 0.04fF
C2384 OR2X1_LOC_151/A AND2X1_LOC_311/a_8_24# 0.01fF
C2385 OR2X1_LOC_60/Y AND2X1_LOC_61/a_8_24# 0.23fF
C2386 OR2X1_LOC_696/A AND2X1_LOC_319/A 0.19fF
C2387 OR2X1_LOC_270/Y AND2X1_LOC_271/a_8_24# 0.05fF
C2388 OR2X1_LOC_130/A OR2X1_LOC_390/B 0.02fF
C2389 AND2X1_LOC_95/Y OR2X1_LOC_174/a_36_216# 0.00fF
C2390 OR2X1_LOC_666/A AND2X1_LOC_860/A 0.24fF
C2391 OR2X1_LOC_122/A AND2X1_LOC_243/Y 0.05fF
C2392 OR2X1_LOC_102/a_8_216# AND2X1_LOC_98/Y 0.14fF
C2393 OR2X1_LOC_158/A OR2X1_LOC_292/a_8_216# 0.01fF
C2394 AND2X1_LOC_12/Y OR2X1_LOC_831/B 0.03fF
C2395 OR2X1_LOC_95/Y OR2X1_LOC_331/a_8_216# 0.06fF
C2396 AND2X1_LOC_17/a_36_24# INPUT_6 0.00fF
C2397 OR2X1_LOC_506/a_36_216# AND2X1_LOC_12/Y 0.02fF
C2398 OR2X1_LOC_804/B OR2X1_LOC_777/B 0.12fF
C2399 OR2X1_LOC_566/A AND2X1_LOC_12/Y 0.15fF
C2400 AND2X1_LOC_217/Y OR2X1_LOC_59/Y 0.09fF
C2401 INPUT_5 OR2X1_LOC_36/a_36_216# 0.00fF
C2402 OR2X1_LOC_71/Y AND2X1_LOC_563/Y 1.62fF
C2403 OR2X1_LOC_147/B OR2X1_LOC_161/B 15.77fF
C2404 OR2X1_LOC_574/A AND2X1_LOC_36/Y 0.01fF
C2405 AND2X1_LOC_363/Y AND2X1_LOC_366/a_8_24# 0.09fF
C2406 OR2X1_LOC_485/Y OR2X1_LOC_484/Y 0.29fF
C2407 OR2X1_LOC_178/a_36_216# OR2X1_LOC_56/A 0.00fF
C2408 AND2X1_LOC_70/Y AND2X1_LOC_110/a_8_24# 0.01fF
C2409 OR2X1_LOC_535/A OR2X1_LOC_502/A 0.00fF
C2410 OR2X1_LOC_18/Y AND2X1_LOC_284/a_36_24# 0.00fF
C2411 AND2X1_LOC_571/a_8_24# AND2X1_LOC_571/Y 0.00fF
C2412 AND2X1_LOC_12/Y OR2X1_LOC_770/A 0.00fF
C2413 OR2X1_LOC_139/A OR2X1_LOC_624/A 0.17fF
C2414 AND2X1_LOC_578/A OR2X1_LOC_142/Y 0.12fF
C2415 OR2X1_LOC_215/Y AND2X1_LOC_7/B 0.25fF
C2416 AND2X1_LOC_330/a_36_24# OR2X1_LOC_51/Y 0.00fF
C2417 OR2X1_LOC_541/A AND2X1_LOC_18/Y 0.05fF
C2418 OR2X1_LOC_188/Y OR2X1_LOC_553/A 0.00fF
C2419 OR2X1_LOC_748/A AND2X1_LOC_792/a_36_24# 0.00fF
C2420 OR2X1_LOC_17/Y OR2X1_LOC_386/a_8_216# 0.00fF
C2421 AND2X1_LOC_715/Y AND2X1_LOC_319/A 0.01fF
C2422 OR2X1_LOC_186/Y OR2X1_LOC_211/a_8_216# 0.08fF
C2423 OR2X1_LOC_46/A OR2X1_LOC_437/A 0.07fF
C2424 OR2X1_LOC_40/Y OR2X1_LOC_165/Y 0.01fF
C2425 OR2X1_LOC_264/Y AND2X1_LOC_265/a_8_24# 0.05fF
C2426 OR2X1_LOC_639/B AND2X1_LOC_44/Y 0.11fF
C2427 AND2X1_LOC_181/a_8_24# OR2X1_LOC_56/A 0.01fF
C2428 OR2X1_LOC_523/Y OR2X1_LOC_113/B 0.01fF
C2429 OR2X1_LOC_109/Y OR2X1_LOC_323/Y 0.27fF
C2430 OR2X1_LOC_591/Y OR2X1_LOC_427/A 0.08fF
C2431 OR2X1_LOC_26/Y AND2X1_LOC_465/A 1.50fF
C2432 OR2X1_LOC_756/B OR2X1_LOC_741/Y 0.02fF
C2433 OR2X1_LOC_653/B AND2X1_LOC_95/Y 0.01fF
C2434 OR2X1_LOC_49/A AND2X1_LOC_129/a_8_24# 0.03fF
C2435 OR2X1_LOC_507/a_8_216# VDD 0.00fF
C2436 OR2X1_LOC_743/A OR2X1_LOC_743/Y 0.02fF
C2437 AND2X1_LOC_548/Y AND2X1_LOC_549/a_8_24# 0.03fF
C2438 OR2X1_LOC_296/a_8_216# OR2X1_LOC_140/B 0.01fF
C2439 AND2X1_LOC_244/A AND2X1_LOC_286/Y 0.00fF
C2440 OR2X1_LOC_49/A AND2X1_LOC_82/a_8_24# 0.00fF
C2441 AND2X1_LOC_721/Y OR2X1_LOC_44/Y 0.02fF
C2442 OR2X1_LOC_160/B OR2X1_LOC_469/Y 0.03fF
C2443 AND2X1_LOC_21/a_8_24# D_INPUT_6 0.01fF
C2444 VDD OR2X1_LOC_144/Y 0.19fF
C2445 AND2X1_LOC_73/a_8_24# AND2X1_LOC_529/a_8_24# 0.23fF
C2446 OR2X1_LOC_720/A AND2X1_LOC_44/Y 0.06fF
C2447 OR2X1_LOC_87/B OR2X1_LOC_34/A 0.00fF
C2448 OR2X1_LOC_516/Y OR2X1_LOC_527/Y 0.07fF
C2449 OR2X1_LOC_114/B OR2X1_LOC_575/A 0.02fF
C2450 AND2X1_LOC_539/Y AND2X1_LOC_512/a_8_24# 0.01fF
C2451 OR2X1_LOC_264/Y VDD 0.12fF
C2452 AND2X1_LOC_377/Y INPUT_0 0.06fF
C2453 OR2X1_LOC_506/A OR2X1_LOC_596/A 0.29fF
C2454 OR2X1_LOC_111/a_8_216# OR2X1_LOC_74/A 0.05fF
C2455 AND2X1_LOC_363/B VDD 0.24fF
C2456 OR2X1_LOC_427/A OR2X1_LOC_583/a_36_216# 0.02fF
C2457 AND2X1_LOC_468/B AND2X1_LOC_477/Y 0.01fF
C2458 OR2X1_LOC_158/A AND2X1_LOC_435/a_8_24# 0.06fF
C2459 OR2X1_LOC_6/A AND2X1_LOC_214/a_36_24# 0.00fF
C2460 AND2X1_LOC_227/Y OR2X1_LOC_437/A 0.03fF
C2461 OR2X1_LOC_528/Y AND2X1_LOC_573/A 0.03fF
C2462 OR2X1_LOC_447/Y OR2X1_LOC_712/B 0.03fF
C2463 OR2X1_LOC_446/Y OR2X1_LOC_707/a_36_216# 0.00fF
C2464 AND2X1_LOC_348/A OR2X1_LOC_56/A 0.03fF
C2465 AND2X1_LOC_99/A OR2X1_LOC_600/A 0.03fF
C2466 OR2X1_LOC_136/a_36_216# OR2X1_LOC_3/Y 0.04fF
C2467 AND2X1_LOC_374/Y OR2X1_LOC_373/Y 0.00fF
C2468 OR2X1_LOC_715/B OR2X1_LOC_805/A 0.07fF
C2469 AND2X1_LOC_768/a_8_24# OR2X1_LOC_427/A 0.04fF
C2470 OR2X1_LOC_62/B OR2X1_LOC_844/B 0.00fF
C2471 OR2X1_LOC_269/a_8_216# AND2X1_LOC_18/Y 0.01fF
C2472 AND2X1_LOC_554/a_36_24# AND2X1_LOC_489/Y 0.00fF
C2473 OR2X1_LOC_334/B OR2X1_LOC_634/a_8_216# 0.08fF
C2474 OR2X1_LOC_516/Y AND2X1_LOC_574/A 0.01fF
C2475 AND2X1_LOC_486/Y OR2X1_LOC_744/A 4.95fF
C2476 OR2X1_LOC_143/a_36_216# OR2X1_LOC_54/Y 0.00fF
C2477 OR2X1_LOC_40/Y AND2X1_LOC_228/Y 0.07fF
C2478 OR2X1_LOC_680/A AND2X1_LOC_499/a_8_24# 0.03fF
C2479 AND2X1_LOC_22/Y AND2X1_LOC_18/a_8_24# 0.01fF
C2480 AND2X1_LOC_810/A OR2X1_LOC_312/Y 0.03fF
C2481 OR2X1_LOC_691/Y OR2X1_LOC_793/B 0.01fF
C2482 OR2X1_LOC_238/Y AND2X1_LOC_786/Y 0.01fF
C2483 OR2X1_LOC_333/B AND2X1_LOC_44/Y 0.09fF
C2484 OR2X1_LOC_482/Y OR2X1_LOC_44/Y 0.03fF
C2485 AND2X1_LOC_12/Y OR2X1_LOC_858/a_36_216# 0.02fF
C2486 AND2X1_LOC_753/B AND2X1_LOC_41/A 0.91fF
C2487 AND2X1_LOC_773/Y OR2X1_LOC_272/a_8_216# 0.47fF
C2488 D_INPUT_0 OR2X1_LOC_395/Y 0.03fF
C2489 OR2X1_LOC_7/A AND2X1_LOC_810/B 0.07fF
C2490 AND2X1_LOC_387/B OR2X1_LOC_161/B 0.07fF
C2491 AND2X1_LOC_729/Y AND2X1_LOC_447/Y 0.01fF
C2492 OR2X1_LOC_677/Y OR2X1_LOC_144/Y 0.12fF
C2493 AND2X1_LOC_772/B AND2X1_LOC_573/A 0.01fF
C2494 INPUT_5 AND2X1_LOC_50/Y 0.87fF
C2495 OR2X1_LOC_691/A OR2X1_LOC_688/Y 0.00fF
C2496 OR2X1_LOC_703/B OR2X1_LOC_468/A 0.02fF
C2497 AND2X1_LOC_658/B OR2X1_LOC_680/A 5.47fF
C2498 OR2X1_LOC_493/a_8_216# OR2X1_LOC_130/A 0.06fF
C2499 OR2X1_LOC_3/Y OR2X1_LOC_135/Y 0.75fF
C2500 OR2X1_LOC_676/Y OR2X1_LOC_194/Y 0.19fF
C2501 AND2X1_LOC_181/Y OR2X1_LOC_7/A 0.03fF
C2502 AND2X1_LOC_56/B AND2X1_LOC_411/a_36_24# 0.00fF
C2503 OR2X1_LOC_502/A AND2X1_LOC_404/A 0.01fF
C2504 OR2X1_LOC_49/A OR2X1_LOC_481/A 0.42fF
C2505 OR2X1_LOC_484/Y OR2X1_LOC_39/A 0.23fF
C2506 AND2X1_LOC_330/a_36_24# OR2X1_LOC_680/A 0.00fF
C2507 OR2X1_LOC_40/Y OR2X1_LOC_585/A 0.20fF
C2508 VDD OR2X1_LOC_643/A 0.29fF
C2509 OR2X1_LOC_99/B AND2X1_LOC_44/Y 0.01fF
C2510 AND2X1_LOC_773/Y OR2X1_LOC_64/Y 0.26fF
C2511 AND2X1_LOC_391/Y AND2X1_LOC_342/Y 0.12fF
C2512 OR2X1_LOC_666/A AND2X1_LOC_287/Y 0.15fF
C2513 OR2X1_LOC_9/Y OR2X1_LOC_485/A 0.11fF
C2514 AND2X1_LOC_713/Y AND2X1_LOC_645/A 0.09fF
C2515 OR2X1_LOC_227/a_8_216# OR2X1_LOC_227/B 0.01fF
C2516 OR2X1_LOC_527/Y AND2X1_LOC_547/a_8_24# -0.00fF
C2517 VDD OR2X1_LOC_778/Y 2.81fF
C2518 OR2X1_LOC_250/Y OR2X1_LOC_517/A 0.01fF
C2519 AND2X1_LOC_342/Y OR2X1_LOC_91/A 0.12fF
C2520 AND2X1_LOC_95/Y OR2X1_LOC_808/B 0.03fF
C2521 OR2X1_LOC_624/B OR2X1_LOC_768/a_8_216# 0.01fF
C2522 OR2X1_LOC_744/A AND2X1_LOC_834/a_8_24# 0.02fF
C2523 OR2X1_LOC_624/A OR2X1_LOC_244/a_8_216# 0.10fF
C2524 VDD OR2X1_LOC_472/A 0.34fF
C2525 OR2X1_LOC_799/A OR2X1_LOC_798/Y 0.25fF
C2526 AND2X1_LOC_334/a_8_24# AND2X1_LOC_219/A 0.04fF
C2527 OR2X1_LOC_840/A OR2X1_LOC_185/A 0.11fF
C2528 AND2X1_LOC_506/a_36_24# AND2X1_LOC_807/Y 0.07fF
C2529 AND2X1_LOC_647/Y OR2X1_LOC_13/B 0.03fF
C2530 OR2X1_LOC_108/Y OR2X1_LOC_280/Y 0.07fF
C2531 OR2X1_LOC_22/Y AND2X1_LOC_244/A 0.03fF
C2532 INPUT_0 OR2X1_LOC_793/A 0.07fF
C2533 OR2X1_LOC_604/A AND2X1_LOC_154/Y 0.01fF
C2534 VDD OR2X1_LOC_420/Y 0.15fF
C2535 OR2X1_LOC_809/a_8_216# OR2X1_LOC_78/B 0.00fF
C2536 OR2X1_LOC_744/A OR2X1_LOC_248/Y 0.19fF
C2537 OR2X1_LOC_165/a_8_216# AND2X1_LOC_168/Y 0.01fF
C2538 OR2X1_LOC_3/Y OR2X1_LOC_815/a_8_216# 0.02fF
C2539 OR2X1_LOC_864/A OR2X1_LOC_78/B 0.10fF
C2540 OR2X1_LOC_496/Y AND2X1_LOC_663/A 0.43fF
C2541 AND2X1_LOC_866/A AND2X1_LOC_455/a_8_24# 0.04fF
C2542 OR2X1_LOC_22/Y OR2X1_LOC_16/A 0.30fF
C2543 OR2X1_LOC_831/A OR2X1_LOC_76/A 0.05fF
C2544 VDD OR2X1_LOC_647/A 0.06fF
C2545 OR2X1_LOC_502/A OR2X1_LOC_828/B 0.31fF
C2546 OR2X1_LOC_316/Y AND2X1_LOC_642/Y 0.01fF
C2547 AND2X1_LOC_95/Y OR2X1_LOC_668/a_36_216# 0.00fF
C2548 AND2X1_LOC_47/Y OR2X1_LOC_392/B 0.03fF
C2549 AND2X1_LOC_36/Y AND2X1_LOC_761/a_8_24# 0.02fF
C2550 AND2X1_LOC_333/a_36_24# OR2X1_LOC_46/A 0.00fF
C2551 OR2X1_LOC_600/A OR2X1_LOC_417/a_8_216# 0.01fF
C2552 OR2X1_LOC_682/Y OR2X1_LOC_91/A 0.01fF
C2553 OR2X1_LOC_545/B OR2X1_LOC_161/B 0.01fF
C2554 OR2X1_LOC_630/Y OR2X1_LOC_574/A 0.02fF
C2555 AND2X1_LOC_47/Y AND2X1_LOC_263/a_8_24# 0.01fF
C2556 OR2X1_LOC_64/Y AND2X1_LOC_243/Y 0.08fF
C2557 OR2X1_LOC_160/B OR2X1_LOC_193/A 0.02fF
C2558 VDD OR2X1_LOC_488/a_8_216# 0.21fF
C2559 OR2X1_LOC_633/B OR2X1_LOC_78/B 0.03fF
C2560 OR2X1_LOC_696/A AND2X1_LOC_721/A 0.04fF
C2561 AND2X1_LOC_59/Y OR2X1_LOC_811/A 0.03fF
C2562 OR2X1_LOC_303/B OR2X1_LOC_578/B 0.11fF
C2563 AND2X1_LOC_31/Y OR2X1_LOC_515/Y 0.34fF
C2564 AND2X1_LOC_773/Y OR2X1_LOC_417/A 0.10fF
C2565 AND2X1_LOC_727/Y GATE_811 0.01fF
C2566 AND2X1_LOC_42/B AND2X1_LOC_92/Y 0.15fF
C2567 AND2X1_LOC_863/a_36_24# AND2X1_LOC_354/B 0.01fF
C2568 AND2X1_LOC_486/Y AND2X1_LOC_840/B 0.07fF
C2569 OR2X1_LOC_315/a_8_216# INPUT_1 0.02fF
C2570 AND2X1_LOC_317/a_8_24# OR2X1_LOC_427/A 0.01fF
C2571 AND2X1_LOC_64/a_8_24# OR2X1_LOC_502/A 0.01fF
C2572 AND2X1_LOC_858/B OR2X1_LOC_279/a_8_216# 0.01fF
C2573 OR2X1_LOC_757/A AND2X1_LOC_711/Y 0.00fF
C2574 OR2X1_LOC_265/a_8_216# OR2X1_LOC_26/Y 0.01fF
C2575 OR2X1_LOC_507/B OR2X1_LOC_510/Y 0.01fF
C2576 OR2X1_LOC_44/Y OR2X1_LOC_586/Y 0.03fF
C2577 AND2X1_LOC_536/a_36_24# OR2X1_LOC_161/A 0.00fF
C2578 AND2X1_LOC_59/Y AND2X1_LOC_533/a_8_24# 0.01fF
C2579 OR2X1_LOC_651/a_8_216# OR2X1_LOC_651/B 0.06fF
C2580 OR2X1_LOC_76/B AND2X1_LOC_56/B 0.12fF
C2581 OR2X1_LOC_426/A OR2X1_LOC_52/B 0.01fF
C2582 OR2X1_LOC_367/B OR2X1_LOC_367/a_8_216# 0.33fF
C2583 OR2X1_LOC_403/B OR2X1_LOC_403/A 0.07fF
C2584 AND2X1_LOC_395/a_8_24# OR2X1_LOC_402/Y 0.03fF
C2585 AND2X1_LOC_141/B OR2X1_LOC_91/A 0.19fF
C2586 OR2X1_LOC_547/B AND2X1_LOC_56/B 1.61fF
C2587 OR2X1_LOC_108/Y OR2X1_LOC_22/Y 0.94fF
C2588 OR2X1_LOC_185/A OR2X1_LOC_222/A 0.01fF
C2589 OR2X1_LOC_829/Y AND2X1_LOC_434/Y 0.01fF
C2590 AND2X1_LOC_713/a_8_24# OR2X1_LOC_31/Y 0.01fF
C2591 AND2X1_LOC_476/A OR2X1_LOC_12/Y 0.14fF
C2592 OR2X1_LOC_619/Y AND2X1_LOC_466/a_36_24# 0.00fF
C2593 AND2X1_LOC_47/Y OR2X1_LOC_113/B 0.08fF
C2594 OR2X1_LOC_145/a_8_216# AND2X1_LOC_621/Y 0.14fF
C2595 OR2X1_LOC_604/A INPUT_1 0.09fF
C2596 OR2X1_LOC_6/B OR2X1_LOC_532/B 0.09fF
C2597 OR2X1_LOC_833/B OR2X1_LOC_269/B 0.02fF
C2598 AND2X1_LOC_12/Y OR2X1_LOC_772/a_8_216# 0.01fF
C2599 AND2X1_LOC_554/B OR2X1_LOC_92/Y 0.06fF
C2600 AND2X1_LOC_583/a_8_24# AND2X1_LOC_51/Y 0.01fF
C2601 AND2X1_LOC_675/A AND2X1_LOC_476/Y 0.05fF
C2602 OR2X1_LOC_417/A AND2X1_LOC_243/Y 0.07fF
C2603 OR2X1_LOC_160/B D_INPUT_0 0.14fF
C2604 OR2X1_LOC_36/Y AND2X1_LOC_624/A 0.03fF
C2605 OR2X1_LOC_18/Y OR2X1_LOC_86/a_8_216# 0.01fF
C2606 OR2X1_LOC_701/Y OR2X1_LOC_748/A 0.00fF
C2607 OR2X1_LOC_49/A D_INPUT_1 0.47fF
C2608 INPUT_1 OR2X1_LOC_66/A 5.99fF
C2609 OR2X1_LOC_624/B OR2X1_LOC_400/a_8_216# 0.01fF
C2610 OR2X1_LOC_411/Y OR2X1_LOC_46/A 0.01fF
C2611 OR2X1_LOC_770/B D_INPUT_1 0.02fF
C2612 D_INPUT_4 OR2X1_LOC_17/Y 0.01fF
C2613 OR2X1_LOC_160/A OR2X1_LOC_835/a_36_216# 0.00fF
C2614 OR2X1_LOC_585/A AND2X1_LOC_644/Y 0.01fF
C2615 OR2X1_LOC_438/a_8_216# OR2X1_LOC_427/A 0.01fF
C2616 AND2X1_LOC_59/Y OR2X1_LOC_649/B 0.10fF
C2617 OR2X1_LOC_91/A OR2X1_LOC_54/Y 3.49fF
C2618 OR2X1_LOC_90/a_36_216# OR2X1_LOC_46/A 0.00fF
C2619 OR2X1_LOC_392/B OR2X1_LOC_598/A 0.10fF
C2620 OR2X1_LOC_864/A OR2X1_LOC_375/A 0.03fF
C2621 AND2X1_LOC_86/B OR2X1_LOC_847/A 1.50fF
C2622 AND2X1_LOC_578/a_8_24# AND2X1_LOC_577/A 0.20fF
C2623 OR2X1_LOC_26/Y OR2X1_LOC_237/Y 0.04fF
C2624 OR2X1_LOC_254/B OR2X1_LOC_269/B 0.03fF
C2625 OR2X1_LOC_450/A AND2X1_LOC_47/Y 0.00fF
C2626 OR2X1_LOC_60/Y OR2X1_LOC_31/Y 0.01fF
C2627 OR2X1_LOC_185/Y AND2X1_LOC_56/B 0.04fF
C2628 OR2X1_LOC_442/a_8_216# OR2X1_LOC_56/A 0.20fF
C2629 OR2X1_LOC_848/B OR2X1_LOC_269/B 0.01fF
C2630 OR2X1_LOC_703/B OR2X1_LOC_449/B 0.15fF
C2631 VDD AND2X1_LOC_270/a_8_24# -0.00fF
C2632 AND2X1_LOC_123/a_8_24# OR2X1_LOC_67/A 0.09fF
C2633 OR2X1_LOC_624/B OR2X1_LOC_847/A 0.00fF
C2634 AND2X1_LOC_53/Y OR2X1_LOC_78/A 0.00fF
C2635 OR2X1_LOC_748/A OR2X1_LOC_44/Y 0.04fF
C2636 AND2X1_LOC_228/Y OR2X1_LOC_7/A 0.00fF
C2637 AND2X1_LOC_73/a_8_24# OR2X1_LOC_532/B 0.03fF
C2638 OR2X1_LOC_87/A OR2X1_LOC_449/B 0.07fF
C2639 OR2X1_LOC_146/a_8_216# AND2X1_LOC_796/A 0.47fF
C2640 OR2X1_LOC_633/B OR2X1_LOC_375/A 1.75fF
C2641 OR2X1_LOC_137/Y OR2X1_LOC_204/Y 0.02fF
C2642 AND2X1_LOC_487/a_36_24# AND2X1_LOC_3/Y 0.00fF
C2643 OR2X1_LOC_318/B OR2X1_LOC_161/B 0.10fF
C2644 AND2X1_LOC_580/A OR2X1_LOC_239/a_8_216# 0.02fF
C2645 OR2X1_LOC_3/Y AND2X1_LOC_848/Y 0.03fF
C2646 AND2X1_LOC_337/a_8_24# AND2X1_LOC_318/Y 0.16fF
C2647 OR2X1_LOC_687/Y AND2X1_LOC_3/Y 0.03fF
C2648 OR2X1_LOC_484/a_8_216# AND2X1_LOC_810/Y 0.05fF
C2649 AND2X1_LOC_141/B AND2X1_LOC_573/A 0.03fF
C2650 AND2X1_LOC_222/Y OR2X1_LOC_428/A 0.03fF
C2651 AND2X1_LOC_12/Y AND2X1_LOC_13/a_8_24# 0.04fF
C2652 OR2X1_LOC_81/Y OR2X1_LOC_83/Y 0.01fF
C2653 OR2X1_LOC_644/B OR2X1_LOC_155/A 0.06fF
C2654 OR2X1_LOC_246/a_36_216# OR2X1_LOC_585/A 0.00fF
C2655 OR2X1_LOC_161/B OR2X1_LOC_854/A 0.14fF
C2656 AND2X1_LOC_191/Y OR2X1_LOC_498/a_8_216# 0.06fF
C2657 OR2X1_LOC_51/Y OR2X1_LOC_47/Y 0.17fF
C2658 OR2X1_LOC_506/B OR2X1_LOC_242/a_8_216# 0.06fF
C2659 AND2X1_LOC_688/a_36_24# AND2X1_LOC_472/B 0.01fF
C2660 AND2X1_LOC_729/Y AND2X1_LOC_729/B 0.03fF
C2661 AND2X1_LOC_798/A OR2X1_LOC_56/A 0.03fF
C2662 OR2X1_LOC_636/A OR2X1_LOC_87/A 0.02fF
C2663 OR2X1_LOC_777/B OR2X1_LOC_356/B 0.96fF
C2664 OR2X1_LOC_223/A OR2X1_LOC_78/A 0.03fF
C2665 OR2X1_LOC_22/Y AND2X1_LOC_661/a_8_24# 0.04fF
C2666 OR2X1_LOC_7/A OR2X1_LOC_585/A 0.15fF
C2667 OR2X1_LOC_18/Y AND2X1_LOC_115/a_8_24# 0.00fF
C2668 AND2X1_LOC_62/a_36_24# OR2X1_LOC_54/Y 0.01fF
C2669 OR2X1_LOC_85/A OR2X1_LOC_8/a_8_216# 0.40fF
C2670 OR2X1_LOC_223/A D_GATE_741 0.01fF
C2671 OR2X1_LOC_70/Y OR2X1_LOC_498/a_8_216# 0.07fF
C2672 AND2X1_LOC_347/Y AND2X1_LOC_866/A 0.07fF
C2673 AND2X1_LOC_356/B AND2X1_LOC_336/a_8_24# 0.01fF
C2674 OR2X1_LOC_837/Y AND2X1_LOC_476/A 0.82fF
C2675 OR2X1_LOC_326/B OR2X1_LOC_532/B 0.00fF
C2676 OR2X1_LOC_160/A AND2X1_LOC_127/a_8_24# 0.05fF
C2677 AND2X1_LOC_86/Y D_INPUT_0 0.02fF
C2678 AND2X1_LOC_40/Y OR2X1_LOC_436/Y 0.10fF
C2679 OR2X1_LOC_532/B OR2X1_LOC_523/Y 0.01fF
C2680 OR2X1_LOC_643/Y OR2X1_LOC_350/a_8_216# 0.00fF
C2681 OR2X1_LOC_428/A OR2X1_LOC_423/Y 0.01fF
C2682 AND2X1_LOC_48/A OR2X1_LOC_828/B 0.00fF
C2683 INPUT_3 D_INPUT_0 4.74fF
C2684 AND2X1_LOC_578/A OR2X1_LOC_238/Y 0.04fF
C2685 OR2X1_LOC_121/B OR2X1_LOC_87/A 0.23fF
C2686 OR2X1_LOC_222/a_36_216# OR2X1_LOC_475/B 0.00fF
C2687 OR2X1_LOC_472/B AND2X1_LOC_56/B 0.03fF
C2688 OR2X1_LOC_300/a_8_216# AND2X1_LOC_786/Y 0.02fF
C2689 AND2X1_LOC_259/Y OR2X1_LOC_481/A 0.04fF
C2690 OR2X1_LOC_542/B OR2X1_LOC_552/A 0.12fF
C2691 AND2X1_LOC_559/a_8_24# OR2X1_LOC_22/Y 0.01fF
C2692 AND2X1_LOC_95/Y OR2X1_LOC_218/Y 0.04fF
C2693 AND2X1_LOC_753/B OR2X1_LOC_207/a_8_216# 0.01fF
C2694 OR2X1_LOC_315/Y AND2X1_LOC_270/a_8_24# 0.25fF
C2695 OR2X1_LOC_46/A OR2X1_LOC_753/A 0.18fF
C2696 AND2X1_LOC_473/Y OR2X1_LOC_268/Y 0.03fF
C2697 OR2X1_LOC_666/A AND2X1_LOC_562/Y 0.03fF
C2698 OR2X1_LOC_855/A AND2X1_LOC_36/Y 0.28fF
C2699 OR2X1_LOC_78/B OR2X1_LOC_608/Y 0.01fF
C2700 OR2X1_LOC_401/B AND2X1_LOC_3/Y 0.01fF
C2701 AND2X1_LOC_627/a_8_24# AND2X1_LOC_36/Y 0.03fF
C2702 OR2X1_LOC_49/A AND2X1_LOC_789/Y 0.18fF
C2703 AND2X1_LOC_336/a_8_24# OR2X1_LOC_22/Y 0.04fF
C2704 OR2X1_LOC_121/B OR2X1_LOC_216/a_8_216# 0.01fF
C2705 OR2X1_LOC_207/B OR2X1_LOC_199/B 0.72fF
C2706 OR2X1_LOC_811/A OR2X1_LOC_733/Y 0.17fF
C2707 D_INPUT_0 OR2X1_LOC_219/B 0.16fF
C2708 OR2X1_LOC_106/A AND2X1_LOC_845/Y 0.01fF
C2709 OR2X1_LOC_462/B OR2X1_LOC_416/a_8_216# 0.02fF
C2710 AND2X1_LOC_95/Y AND2X1_LOC_289/a_8_24# 0.01fF
C2711 OR2X1_LOC_114/B OR2X1_LOC_735/B 0.03fF
C2712 OR2X1_LOC_680/A OR2X1_LOC_47/Y 0.03fF
C2713 OR2X1_LOC_65/Y AND2X1_LOC_201/a_8_24# 0.01fF
C2714 OR2X1_LOC_343/B OR2X1_LOC_579/B 0.13fF
C2715 AND2X1_LOC_27/a_8_24# AND2X1_LOC_51/Y 0.01fF
C2716 AND2X1_LOC_860/A OR2X1_LOC_13/B 0.28fF
C2717 AND2X1_LOC_151/a_8_24# AND2X1_LOC_796/Y 0.20fF
C2718 AND2X1_LOC_59/Y AND2X1_LOC_237/a_8_24# 0.01fF
C2719 OR2X1_LOC_366/B OR2X1_LOC_366/A 0.08fF
C2720 OR2X1_LOC_512/A OR2X1_LOC_779/B 0.01fF
C2721 AND2X1_LOC_67/Y OR2X1_LOC_814/A 0.02fF
C2722 OR2X1_LOC_404/Y AND2X1_LOC_107/a_8_24# 0.01fF
C2723 OR2X1_LOC_387/Y OR2X1_LOC_95/Y 0.02fF
C2724 OR2X1_LOC_791/A OR2X1_LOC_345/a_8_216# 0.18fF
C2725 OR2X1_LOC_87/B D_INPUT_1 0.18fF
C2726 OR2X1_LOC_419/Y AND2X1_LOC_624/A 0.03fF
C2727 OR2X1_LOC_223/A OR2X1_LOC_155/A 0.03fF
C2728 OR2X1_LOC_709/A AND2X1_LOC_64/Y 0.06fF
C2729 AND2X1_LOC_359/a_8_24# AND2X1_LOC_721/A 0.01fF
C2730 D_INPUT_3 AND2X1_LOC_42/B 0.03fF
C2731 OR2X1_LOC_45/B AND2X1_LOC_721/Y 0.99fF
C2732 OR2X1_LOC_118/Y OR2X1_LOC_88/a_8_216# 0.01fF
C2733 OR2X1_LOC_415/Y OR2X1_LOC_548/a_36_216# 0.00fF
C2734 OR2X1_LOC_525/Y AND2X1_LOC_796/A 0.10fF
C2735 OR2X1_LOC_619/Y OR2X1_LOC_72/Y 0.07fF
C2736 AND2X1_LOC_3/Y OR2X1_LOC_786/Y 0.09fF
C2737 OR2X1_LOC_798/Y OR2X1_LOC_446/B 0.22fF
C2738 OR2X1_LOC_22/Y AND2X1_LOC_687/Y 0.02fF
C2739 AND2X1_LOC_722/A OR2X1_LOC_437/A 0.07fF
C2740 OR2X1_LOC_605/A OR2X1_LOC_223/A 0.01fF
C2741 AND2X1_LOC_85/a_8_24# D_INPUT_1 0.02fF
C2742 AND2X1_LOC_43/B OR2X1_LOC_228/Y 0.08fF
C2743 AND2X1_LOC_521/a_8_24# OR2X1_LOC_392/B 0.22fF
C2744 AND2X1_LOC_100/a_8_24# AND2X1_LOC_216/A 0.17fF
C2745 OR2X1_LOC_49/A OR2X1_LOC_15/a_8_216# 0.01fF
C2746 OR2X1_LOC_412/a_36_216# INPUT_1 0.02fF
C2747 AND2X1_LOC_624/A OR2X1_LOC_152/A 0.03fF
C2748 AND2X1_LOC_211/B OR2X1_LOC_173/a_36_216# 0.00fF
C2749 AND2X1_LOC_56/B OR2X1_LOC_552/A 0.02fF
C2750 AND2X1_LOC_43/B OR2X1_LOC_513/Y 0.02fF
C2751 AND2X1_LOC_3/Y OR2X1_LOC_644/A 0.02fF
C2752 OR2X1_LOC_208/A OR2X1_LOC_160/B 1.16fF
C2753 OR2X1_LOC_653/B AND2X1_LOC_22/Y 0.01fF
C2754 AND2X1_LOC_560/a_8_24# VDD 0.00fF
C2755 OR2X1_LOC_89/a_36_216# AND2X1_LOC_243/Y 0.01fF
C2756 OR2X1_LOC_88/A OR2X1_LOC_72/Y 0.01fF
C2757 OR2X1_LOC_614/Y AND2X1_LOC_22/Y 0.27fF
C2758 OR2X1_LOC_468/A OR2X1_LOC_390/B 0.00fF
C2759 OR2X1_LOC_571/a_8_216# OR2X1_LOC_579/A 0.03fF
C2760 OR2X1_LOC_325/A OR2X1_LOC_532/Y 0.23fF
C2761 AND2X1_LOC_564/B OR2X1_LOC_40/Y 0.02fF
C2762 AND2X1_LOC_53/Y OR2X1_LOC_228/a_8_216# 0.04fF
C2763 AND2X1_LOC_91/B VDD 4.07fF
C2764 OR2X1_LOC_696/A OR2X1_LOC_107/a_36_216# 0.00fF
C2765 AND2X1_LOC_64/Y AND2X1_LOC_70/Y 0.70fF
C2766 AND2X1_LOC_56/B OR2X1_LOC_578/B 0.03fF
C2767 OR2X1_LOC_175/Y AND2X1_LOC_18/Y 0.03fF
C2768 OR2X1_LOC_48/B OR2X1_LOC_424/Y 0.03fF
C2769 AND2X1_LOC_243/a_36_24# AND2X1_LOC_243/Y 0.01fF
C2770 AND2X1_LOC_47/Y OR2X1_LOC_532/B 0.88fF
C2771 OR2X1_LOC_754/a_8_216# OR2X1_LOC_753/Y 0.01fF
C2772 AND2X1_LOC_663/B AND2X1_LOC_721/A 0.03fF
C2773 AND2X1_LOC_56/B OR2X1_LOC_151/a_8_216# 0.02fF
C2774 OR2X1_LOC_471/Y OR2X1_LOC_620/A 0.12fF
C2775 AND2X1_LOC_828/a_8_24# AND2X1_LOC_771/B 0.01fF
C2776 OR2X1_LOC_9/Y OR2X1_LOC_633/A 0.04fF
C2777 OR2X1_LOC_696/A AND2X1_LOC_605/Y 0.01fF
C2778 OR2X1_LOC_589/A OR2X1_LOC_829/A 0.80fF
C2779 OR2X1_LOC_154/A OR2X1_LOC_317/B 0.03fF
C2780 OR2X1_LOC_40/Y AND2X1_LOC_341/a_36_24# 0.00fF
C2781 OR2X1_LOC_691/Y AND2X1_LOC_18/Y 0.03fF
C2782 AND2X1_LOC_22/Y OR2X1_LOC_641/Y 0.46fF
C2783 OR2X1_LOC_209/a_8_216# OR2X1_LOC_550/B 0.40fF
C2784 AND2X1_LOC_59/Y OR2X1_LOC_777/B 0.17fF
C2785 OR2X1_LOC_161/A OR2X1_LOC_712/B 0.04fF
C2786 OR2X1_LOC_45/B OR2X1_LOC_496/a_36_216# 0.00fF
C2787 OR2X1_LOC_177/Y AND2X1_LOC_778/Y 0.12fF
C2788 OR2X1_LOC_160/B AND2X1_LOC_438/a_8_24# 0.04fF
C2789 OR2X1_LOC_31/Y AND2X1_LOC_660/A 0.05fF
C2790 VDD OR2X1_LOC_821/a_8_216# 0.00fF
C2791 OR2X1_LOC_18/Y D_INPUT_6 1.63fF
C2792 AND2X1_LOC_287/Y OR2X1_LOC_13/B 0.19fF
C2793 AND2X1_LOC_110/Y OR2X1_LOC_486/Y 0.03fF
C2794 AND2X1_LOC_95/Y OR2X1_LOC_703/Y 0.01fF
C2795 VDD OR2X1_LOC_522/Y 0.04fF
C2796 OR2X1_LOC_377/A AND2X1_LOC_36/Y 8.97fF
C2797 AND2X1_LOC_95/Y OR2X1_LOC_500/a_8_216# 0.01fF
C2798 OR2X1_LOC_62/B OR2X1_LOC_493/Y 0.03fF
C2799 AND2X1_LOC_201/a_8_24# OR2X1_LOC_72/Y 0.06fF
C2800 INPUT_1 OR2X1_LOC_98/B 0.10fF
C2801 OR2X1_LOC_89/A OR2X1_LOC_384/Y 0.13fF
C2802 OR2X1_LOC_648/A AND2X1_LOC_433/a_8_24# 0.02fF
C2803 VDD OR2X1_LOC_364/a_8_216# 0.00fF
C2804 OR2X1_LOC_813/Y AND2X1_LOC_845/Y 0.01fF
C2805 AND2X1_LOC_736/Y AND2X1_LOC_544/Y 1.68fF
C2806 AND2X1_LOC_276/Y OR2X1_LOC_521/a_36_216# 0.00fF
C2807 OR2X1_LOC_474/Y OR2X1_LOC_267/Y 0.05fF
C2808 AND2X1_LOC_367/A OR2X1_LOC_428/A 0.05fF
C2809 AND2X1_LOC_592/Y AND2X1_LOC_724/Y 0.00fF
C2810 INPUT_0 OR2X1_LOC_12/Y 0.02fF
C2811 OR2X1_LOC_538/A OR2X1_LOC_161/B 0.04fF
C2812 AND2X1_LOC_663/B AND2X1_LOC_217/a_8_24# 0.13fF
C2813 AND2X1_LOC_22/Y OR2X1_LOC_808/B 0.03fF
C2814 OR2X1_LOC_160/B AND2X1_LOC_505/a_8_24# 0.03fF
C2815 OR2X1_LOC_532/B OR2X1_LOC_598/A 0.31fF
C2816 OR2X1_LOC_203/Y AND2X1_LOC_36/Y 0.06fF
C2817 OR2X1_LOC_155/a_8_216# OR2X1_LOC_803/A 0.01fF
C2818 OR2X1_LOC_337/A OR2X1_LOC_337/a_8_216# 0.18fF
C2819 OR2X1_LOC_532/B OR2X1_LOC_717/a_36_216# 0.00fF
C2820 AND2X1_LOC_367/A OR2X1_LOC_595/A 0.10fF
C2821 AND2X1_LOC_787/A AND2X1_LOC_168/a_8_24# 0.01fF
C2822 OR2X1_LOC_615/Y AND2X1_LOC_620/Y 1.01fF
C2823 AND2X1_LOC_443/Y AND2X1_LOC_477/Y 0.04fF
C2824 AND2X1_LOC_758/a_36_24# OR2X1_LOC_600/A 0.00fF
C2825 OR2X1_LOC_450/A OR2X1_LOC_450/a_8_216# 0.01fF
C2826 AND2X1_LOC_259/Y AND2X1_LOC_789/Y 0.02fF
C2827 AND2X1_LOC_824/B OR2X1_LOC_334/A 0.01fF
C2828 OR2X1_LOC_78/A OR2X1_LOC_777/a_8_216# 0.01fF
C2829 OR2X1_LOC_18/Y AND2X1_LOC_242/B 0.82fF
C2830 AND2X1_LOC_59/Y OR2X1_LOC_831/B 0.10fF
C2831 OR2X1_LOC_609/Y AND2X1_LOC_647/B 0.78fF
C2832 AND2X1_LOC_586/a_8_24# OR2X1_LOC_855/A 0.05fF
C2833 AND2X1_LOC_539/Y OR2X1_LOC_306/a_36_216# 0.00fF
C2834 OR2X1_LOC_49/A AND2X1_LOC_414/a_8_24# 0.03fF
C2835 AND2X1_LOC_621/Y AND2X1_LOC_580/a_8_24# 0.01fF
C2836 OR2X1_LOC_620/Y AND2X1_LOC_44/Y 0.14fF
C2837 OR2X1_LOC_178/a_8_216# OR2X1_LOC_59/Y 0.01fF
C2838 OR2X1_LOC_188/a_8_216# AND2X1_LOC_59/Y 0.01fF
C2839 AND2X1_LOC_729/Y AND2X1_LOC_220/B 0.03fF
C2840 AND2X1_LOC_570/Y AND2X1_LOC_658/A 0.03fF
C2841 OR2X1_LOC_139/A OR2X1_LOC_161/A 0.07fF
C2842 OR2X1_LOC_375/A OR2X1_LOC_121/A 0.73fF
C2843 OR2X1_LOC_130/A OR2X1_LOC_390/a_36_216# -0.01fF
C2844 OR2X1_LOC_49/A AND2X1_LOC_95/Y 0.02fF
C2845 AND2X1_LOC_784/Y OR2X1_LOC_516/B 0.16fF
C2846 OR2X1_LOC_449/B OR2X1_LOC_390/B 0.05fF
C2847 OR2X1_LOC_335/Y OR2X1_LOC_160/B 0.10fF
C2848 AND2X1_LOC_347/Y OR2X1_LOC_40/Y 0.00fF
C2849 OR2X1_LOC_49/A OR2X1_LOC_633/Y 0.07fF
C2850 OR2X1_LOC_40/Y AND2X1_LOC_857/Y 0.07fF
C2851 AND2X1_LOC_244/A OR2X1_LOC_39/A 0.02fF
C2852 AND2X1_LOC_574/a_8_24# AND2X1_LOC_500/Y 0.01fF
C2853 OR2X1_LOC_310/Y OR2X1_LOC_426/B 0.01fF
C2854 OR2X1_LOC_212/a_36_216# OR2X1_LOC_486/Y 0.02fF
C2855 AND2X1_LOC_12/Y OR2X1_LOC_161/B 1.33fF
C2856 OR2X1_LOC_179/a_8_216# VDD 0.00fF
C2857 AND2X1_LOC_670/a_8_24# AND2X1_LOC_36/Y 0.00fF
C2858 OR2X1_LOC_170/A OR2X1_LOC_175/Y 0.07fF
C2859 AND2X1_LOC_203/Y AND2X1_LOC_215/A 0.01fF
C2860 AND2X1_LOC_204/Y AND2X1_LOC_205/a_8_24# 0.03fF
C2861 AND2X1_LOC_164/a_36_24# OR2X1_LOC_648/A 0.01fF
C2862 OR2X1_LOC_467/a_8_216# OR2X1_LOC_161/B 0.02fF
C2863 OR2X1_LOC_793/A AND2X1_LOC_7/B 0.15fF
C2864 OR2X1_LOC_694/a_8_216# OR2X1_LOC_766/a_8_216# 0.47fF
C2865 OR2X1_LOC_427/A OR2X1_LOC_765/a_8_216# 0.01fF
C2866 OR2X1_LOC_16/A OR2X1_LOC_39/A 0.10fF
C2867 OR2X1_LOC_154/A AND2X1_LOC_44/Y 0.37fF
C2868 OR2X1_LOC_858/A AND2X1_LOC_498/a_36_24# 0.01fF
C2869 AND2X1_LOC_40/Y OR2X1_LOC_160/B 0.38fF
C2870 OR2X1_LOC_759/A AND2X1_LOC_866/B 0.02fF
C2871 AND2X1_LOC_863/Y AND2X1_LOC_212/a_8_24# 0.04fF
C2872 OR2X1_LOC_335/A OR2X1_LOC_787/Y 0.01fF
C2873 AND2X1_LOC_541/Y OR2X1_LOC_427/A 0.01fF
C2874 AND2X1_LOC_59/Y OR2X1_LOC_344/A 0.04fF
C2875 OR2X1_LOC_11/Y OR2X1_LOC_12/Y 0.18fF
C2876 OR2X1_LOC_501/B OR2X1_LOC_630/B 1.11fF
C2877 OR2X1_LOC_858/A OR2X1_LOC_499/B 0.11fF
C2878 OR2X1_LOC_325/a_36_216# AND2X1_LOC_110/Y 0.00fF
C2879 OR2X1_LOC_40/Y AND2X1_LOC_833/a_36_24# 0.00fF
C2880 INPUT_0 AND2X1_LOC_54/a_8_24# 0.14fF
C2881 AND2X1_LOC_719/Y AND2X1_LOC_621/Y 0.03fF
C2882 INPUT_0 OR2X1_LOC_837/Y 0.07fF
C2883 OR2X1_LOC_36/Y AND2X1_LOC_774/A 0.21fF
C2884 OR2X1_LOC_7/A OR2X1_LOC_230/Y 0.02fF
C2885 OR2X1_LOC_756/B OR2X1_LOC_235/B 0.00fF
C2886 OR2X1_LOC_154/A OR2X1_LOC_514/a_8_216# 0.03fF
C2887 AND2X1_LOC_866/A OR2X1_LOC_437/A 0.19fF
C2888 OR2X1_LOC_7/A OR2X1_LOC_368/Y 0.18fF
C2889 OR2X1_LOC_49/A OR2X1_LOC_99/Y 0.03fF
C2890 OR2X1_LOC_502/A OR2X1_LOC_78/A 1.30fF
C2891 OR2X1_LOC_653/Y AND2X1_LOC_172/a_8_24# -0.05fF
C2892 AND2X1_LOC_64/Y OR2X1_LOC_206/a_8_216# 0.01fF
C2893 VDD AND2X1_LOC_809/A 0.25fF
C2894 AND2X1_LOC_673/a_8_24# OR2X1_LOC_428/A 0.01fF
C2895 OR2X1_LOC_378/Y OR2X1_LOC_375/a_8_216# 0.39fF
C2896 AND2X1_LOC_566/B AND2X1_LOC_303/A 0.01fF
C2897 AND2X1_LOC_787/A OR2X1_LOC_485/A 0.03fF
C2898 OR2X1_LOC_160/B OR2X1_LOC_537/A 0.01fF
C2899 OR2X1_LOC_519/a_8_216# OR2X1_LOC_426/B 0.03fF
C2900 VDD OR2X1_LOC_799/A 0.15fF
C2901 AND2X1_LOC_720/a_8_24# OR2X1_LOC_51/Y 0.01fF
C2902 AND2X1_LOC_64/Y OR2X1_LOC_404/Y 0.09fF
C2903 OR2X1_LOC_604/A AND2X1_LOC_624/A 0.10fF
C2904 OR2X1_LOC_43/A OR2X1_LOC_829/A 0.27fF
C2905 OR2X1_LOC_108/Y OR2X1_LOC_39/A 0.19fF
C2906 AND2X1_LOC_729/Y AND2X1_LOC_209/a_8_24# 0.01fF
C2907 OR2X1_LOC_51/Y OR2X1_LOC_625/Y 0.12fF
C2908 OR2X1_LOC_748/A OR2X1_LOC_382/A 0.57fF
C2909 OR2X1_LOC_107/a_8_216# OR2X1_LOC_427/A 0.03fF
C2910 OR2X1_LOC_678/Y OR2X1_LOC_623/B 0.03fF
C2911 AND2X1_LOC_211/B OR2X1_LOC_16/A 0.49fF
C2912 OR2X1_LOC_864/A OR2X1_LOC_549/A 0.07fF
C2913 OR2X1_LOC_450/A AND2X1_LOC_695/a_8_24# 0.24fF
C2914 OR2X1_LOC_74/A OR2X1_LOC_428/A 0.07fF
C2915 OR2X1_LOC_405/A OR2X1_LOC_648/A 0.31fF
C2916 OR2X1_LOC_229/a_8_216# OR2X1_LOC_7/A -0.03fF
C2917 AND2X1_LOC_588/B AND2X1_LOC_51/Y 0.00fF
C2918 AND2X1_LOC_79/Y OR2X1_LOC_161/B 0.00fF
C2919 OR2X1_LOC_280/Y OR2X1_LOC_373/Y 0.00fF
C2920 OR2X1_LOC_329/a_8_216# OR2X1_LOC_312/Y 0.57fF
C2921 OR2X1_LOC_756/B OR2X1_LOC_814/a_36_216# 0.00fF
C2922 OR2X1_LOC_240/A OR2X1_LOC_549/A 0.09fF
C2923 OR2X1_LOC_45/B OR2X1_LOC_304/Y 0.09fF
C2924 AND2X1_LOC_310/a_36_24# OR2X1_LOC_185/A 0.00fF
C2925 OR2X1_LOC_492/a_8_216# OR2X1_LOC_529/Y 0.01fF
C2926 OR2X1_LOC_490/Y OR2X1_LOC_595/A 0.01fF
C2927 OR2X1_LOC_139/A AND2X1_LOC_51/Y 0.01fF
C2928 AND2X1_LOC_43/B OR2X1_LOC_702/a_36_216# 0.00fF
C2929 OR2X1_LOC_74/A OR2X1_LOC_595/A 0.15fF
C2930 OR2X1_LOC_633/B OR2X1_LOC_549/A 0.01fF
C2931 OR2X1_LOC_86/A OR2X1_LOC_71/A 0.00fF
C2932 OR2X1_LOC_662/A AND2X1_LOC_19/Y 0.07fF
C2933 AND2X1_LOC_50/Y OR2X1_LOC_651/B 0.01fF
C2934 VDD AND2X1_LOC_303/B 0.02fF
C2935 OR2X1_LOC_865/B OR2X1_LOC_571/a_8_216# 0.06fF
C2936 AND2X1_LOC_101/B AND2X1_LOC_243/Y 0.00fF
C2937 OR2X1_LOC_753/A INPUT_2 0.02fF
C2938 AND2X1_LOC_508/B OR2X1_LOC_44/Y 0.00fF
C2939 INPUT_0 OR2X1_LOC_459/B 0.40fF
C2940 AND2X1_LOC_570/Y OR2X1_LOC_497/a_8_216# 0.01fF
C2941 OR2X1_LOC_377/A OR2X1_LOC_633/a_8_216# 0.02fF
C2942 OR2X1_LOC_532/B OR2X1_LOC_186/a_8_216# 0.01fF
C2943 OR2X1_LOC_831/A OR2X1_LOC_794/a_8_216# 0.01fF
C2944 OR2X1_LOC_89/A OR2X1_LOC_131/a_8_216# 0.01fF
C2945 OR2X1_LOC_822/a_8_216# OR2X1_LOC_585/A 0.01fF
C2946 AND2X1_LOC_859/Y AND2X1_LOC_285/Y 0.02fF
C2947 AND2X1_LOC_508/a_8_24# OR2X1_LOC_44/Y 0.01fF
C2948 OR2X1_LOC_364/A AND2X1_LOC_92/Y 0.07fF
C2949 AND2X1_LOC_712/Y OR2X1_LOC_743/A 0.01fF
C2950 AND2X1_LOC_594/a_36_24# OR2X1_LOC_435/Y 0.00fF
C2951 AND2X1_LOC_86/Y AND2X1_LOC_40/Y 0.09fF
C2952 OR2X1_LOC_185/Y AND2X1_LOC_92/Y 0.53fF
C2953 OR2X1_LOC_64/Y OR2X1_LOC_12/Y 0.23fF
C2954 OR2X1_LOC_36/Y AND2X1_LOC_434/a_8_24# 0.01fF
C2955 AND2X1_LOC_447/Y OR2X1_LOC_52/B 0.01fF
C2956 OR2X1_LOC_448/a_8_216# OR2X1_LOC_784/Y 0.43fF
C2957 AND2X1_LOC_40/a_8_24# AND2X1_LOC_1/Y 0.01fF
C2958 AND2X1_LOC_736/Y AND2X1_LOC_550/A 0.03fF
C2959 OR2X1_LOC_850/B OR2X1_LOC_161/A 0.01fF
C2960 OR2X1_LOC_45/B AND2X1_LOC_471/a_8_24# 0.01fF
C2961 OR2X1_LOC_160/A AND2X1_LOC_424/a_8_24# 0.02fF
C2962 OR2X1_LOC_151/A OR2X1_LOC_473/Y 0.03fF
C2963 AND2X1_LOC_841/B OR2X1_LOC_48/B 0.19fF
C2964 AND2X1_LOC_554/B OR2X1_LOC_600/A 0.04fF
C2965 OR2X1_LOC_26/Y AND2X1_LOC_637/a_36_24# -0.00fF
C2966 OR2X1_LOC_31/Y OR2X1_LOC_56/Y 0.24fF
C2967 OR2X1_LOC_91/A OR2X1_LOC_26/Y 0.32fF
C2968 OR2X1_LOC_182/a_8_216# OR2X1_LOC_365/B 0.12fF
C2969 OR2X1_LOC_123/a_36_216# OR2X1_LOC_633/B 0.00fF
C2970 AND2X1_LOC_321/a_8_24# OR2X1_LOC_739/A 0.01fF
C2971 OR2X1_LOC_564/B OR2X1_LOC_192/A 0.31fF
C2972 AND2X1_LOC_393/a_8_24# OR2X1_LOC_756/B 0.02fF
C2973 AND2X1_LOC_12/Y OR2X1_LOC_61/Y 0.11fF
C2974 OR2X1_LOC_529/a_8_216# OR2X1_LOC_427/A 0.03fF
C2975 OR2X1_LOC_13/B AND2X1_LOC_562/Y 0.10fF
C2976 AND2X1_LOC_40/Y OR2X1_LOC_553/A 0.09fF
C2977 AND2X1_LOC_850/A OR2X1_LOC_44/Y 0.12fF
C2978 AND2X1_LOC_72/a_8_24# OR2X1_LOC_78/A 0.01fF
C2979 OR2X1_LOC_405/A OR2X1_LOC_405/a_8_216# 0.16fF
C2980 AND2X1_LOC_191/B AND2X1_LOC_465/a_8_24# 0.19fF
C2981 OR2X1_LOC_154/A OR2X1_LOC_61/a_8_216# 0.01fF
C2982 AND2X1_LOC_858/B OR2X1_LOC_89/A 0.03fF
C2983 OR2X1_LOC_157/a_8_216# OR2X1_LOC_2/Y 0.04fF
C2984 OR2X1_LOC_494/a_36_216# AND2X1_LOC_359/B 0.00fF
C2985 OR2X1_LOC_91/A OR2X1_LOC_89/A 0.13fF
C2986 OR2X1_LOC_70/Y AND2X1_LOC_436/Y 0.01fF
C2987 AND2X1_LOC_59/Y OR2X1_LOC_493/A 0.20fF
C2988 AND2X1_LOC_91/B OR2X1_LOC_845/A 0.17fF
C2989 OR2X1_LOC_31/Y AND2X1_LOC_457/a_8_24# 0.01fF
C2990 AND2X1_LOC_12/Y AND2X1_LOC_536/a_8_24# 0.01fF
C2991 OR2X1_LOC_189/a_8_216# AND2X1_LOC_565/Y 0.49fF
C2992 AND2X1_LOC_305/a_8_24# OR2X1_LOC_375/A 0.00fF
C2993 OR2X1_LOC_863/B OR2X1_LOC_35/Y 0.00fF
C2994 OR2X1_LOC_417/A OR2X1_LOC_12/Y 0.07fF
C2995 OR2X1_LOC_656/B OR2X1_LOC_805/A 0.01fF
C2996 AND2X1_LOC_849/A AND2X1_LOC_244/a_8_24# 0.09fF
C2997 OR2X1_LOC_791/B OR2X1_LOC_555/B 0.06fF
C2998 OR2X1_LOC_252/Y AND2X1_LOC_621/Y 0.03fF
C2999 AND2X1_LOC_785/A OR2X1_LOC_406/A 0.01fF
C3000 AND2X1_LOC_667/a_36_24# AND2X1_LOC_65/A 0.00fF
C3001 AND2X1_LOC_421/a_8_24# OR2X1_LOC_269/B 0.01fF
C3002 AND2X1_LOC_737/a_8_24# OR2X1_LOC_52/B 0.01fF
C3003 AND2X1_LOC_86/B OR2X1_LOC_78/Y 0.03fF
C3004 OR2X1_LOC_235/B OR2X1_LOC_233/a_36_216# 0.01fF
C3005 AND2X1_LOC_521/a_8_24# OR2X1_LOC_532/B 0.01fF
C3006 AND2X1_LOC_107/a_8_24# OR2X1_LOC_362/A 0.01fF
C3007 AND2X1_LOC_12/Y OR2X1_LOC_846/a_8_216# 0.01fF
C3008 AND2X1_LOC_354/Y AND2X1_LOC_319/A 0.31fF
C3009 AND2X1_LOC_857/Y OR2X1_LOC_7/A 0.11fF
C3010 OR2X1_LOC_502/A OR2X1_LOC_155/A 0.20fF
C3011 OR2X1_LOC_574/A OR2X1_LOC_274/Y 0.05fF
C3012 AND2X1_LOC_705/Y OR2X1_LOC_95/Y 0.15fF
C3013 OR2X1_LOC_493/a_8_216# OR2X1_LOC_121/B 0.01fF
C3014 OR2X1_LOC_759/A AND2X1_LOC_664/a_8_24# 0.01fF
C3015 AND2X1_LOC_40/Y OR2X1_LOC_219/B 0.07fF
C3016 OR2X1_LOC_624/B OR2X1_LOC_78/Y 0.02fF
C3017 OR2X1_LOC_532/B OR2X1_LOC_646/B 0.43fF
C3018 AND2X1_LOC_160/a_8_24# OR2X1_LOC_3/Y 0.01fF
C3019 AND2X1_LOC_324/a_36_24# OR2X1_LOC_56/A 0.00fF
C3020 AND2X1_LOC_562/B OR2X1_LOC_3/Y 0.40fF
C3021 OR2X1_LOC_760/a_8_216# OR2X1_LOC_16/A 0.01fF
C3022 AND2X1_LOC_271/a_8_24# AND2X1_LOC_7/B 0.02fF
C3023 OR2X1_LOC_320/Y AND2X1_LOC_857/Y 0.10fF
C3024 OR2X1_LOC_823/a_8_216# OR2X1_LOC_26/Y 0.01fF
C3025 OR2X1_LOC_109/Y AND2X1_LOC_374/Y 0.02fF
C3026 AND2X1_LOC_391/a_8_24# AND2X1_LOC_348/a_8_24# 0.23fF
C3027 OR2X1_LOC_271/B AND2X1_LOC_318/a_8_24# 0.06fF
C3028 AND2X1_LOC_848/a_8_24# OR2X1_LOC_44/Y 0.01fF
C3029 AND2X1_LOC_559/a_8_24# OR2X1_LOC_39/A 0.03fF
C3030 AND2X1_LOC_22/Y AND2X1_LOC_289/a_8_24# 0.02fF
C3031 OR2X1_LOC_26/Y AND2X1_LOC_573/A 0.09fF
C3032 AND2X1_LOC_48/A OR2X1_LOC_78/A 0.01fF
C3033 OR2X1_LOC_743/A OR2X1_LOC_422/Y 0.21fF
C3034 AND2X1_LOC_70/Y AND2X1_LOC_600/a_8_24# 0.01fF
C3035 OR2X1_LOC_246/Y OR2X1_LOC_85/A 0.40fF
C3036 AND2X1_LOC_532/a_8_24# OR2X1_LOC_485/A 0.03fF
C3037 AND2X1_LOC_448/Y OR2X1_LOC_52/B 0.05fF
C3038 OR2X1_LOC_46/A AND2X1_LOC_222/a_8_24# 0.09fF
C3039 OR2X1_LOC_804/a_36_216# OR2X1_LOC_121/B 0.00fF
C3040 AND2X1_LOC_392/A AND2X1_LOC_170/B 0.03fF
C3041 AND2X1_LOC_51/A AND2X1_LOC_47/a_8_24# 0.01fF
C3042 AND2X1_LOC_390/B OR2X1_LOC_427/A 0.07fF
C3043 AND2X1_LOC_337/B AND2X1_LOC_662/B 0.01fF
C3044 OR2X1_LOC_64/Y OR2X1_LOC_763/a_36_216# 0.00fF
C3045 AND2X1_LOC_36/Y OR2X1_LOC_732/A 0.03fF
C3046 AND2X1_LOC_390/B AND2X1_LOC_801/a_8_24# 0.01fF
C3047 AND2X1_LOC_94/Y INPUT_1 0.17fF
C3048 VDD AND2X1_LOC_859/B 0.01fF
C3049 OR2X1_LOC_89/A AND2X1_LOC_573/A 0.09fF
C3050 OR2X1_LOC_671/Y D_INPUT_1 0.25fF
C3051 AND2X1_LOC_95/Y OR2X1_LOC_33/B 0.00fF
C3052 AND2X1_LOC_34/Y OR2X1_LOC_24/Y 0.04fF
C3053 OR2X1_LOC_589/A OR2X1_LOC_597/Y 0.04fF
C3054 OR2X1_LOC_467/A OR2X1_LOC_780/a_36_216# 0.00fF
C3055 OR2X1_LOC_473/A AND2X1_LOC_625/a_36_24# 0.01fF
C3056 AND2X1_LOC_303/a_8_24# D_INPUT_0 0.03fF
C3057 AND2X1_LOC_40/Y OR2X1_LOC_647/a_36_216# 0.02fF
C3058 OR2X1_LOC_703/Y OR2X1_LOC_788/B 0.81fF
C3059 AND2X1_LOC_692/a_36_24# OR2X1_LOC_706/A 0.00fF
C3060 AND2X1_LOC_647/Y OR2X1_LOC_595/A 0.00fF
C3061 OR2X1_LOC_563/A OR2X1_LOC_344/a_8_216# 0.03fF
C3062 AND2X1_LOC_548/a_8_24# OR2X1_LOC_680/A 0.02fF
C3063 OR2X1_LOC_624/Y AND2X1_LOC_47/Y 0.03fF
C3064 OR2X1_LOC_654/A AND2X1_LOC_56/B 0.03fF
C3065 AND2X1_LOC_326/A OR2X1_LOC_619/Y 0.01fF
C3066 OR2X1_LOC_91/A AND2X1_LOC_864/a_8_24# 0.08fF
C3067 OR2X1_LOC_669/Y OR2X1_LOC_26/Y 0.21fF
C3068 OR2X1_LOC_173/Y AND2X1_LOC_175/a_8_24# 0.23fF
C3069 OR2X1_LOC_358/A OR2X1_LOC_390/A 1.67fF
C3070 AND2X1_LOC_392/A AND2X1_LOC_721/A 0.15fF
C3071 OR2X1_LOC_261/Y OR2X1_LOC_748/A 0.01fF
C3072 OR2X1_LOC_19/B OR2X1_LOC_278/Y 0.02fF
C3073 OR2X1_LOC_837/B AND2X1_LOC_825/a_8_24# 0.01fF
C3074 AND2X1_LOC_44/Y OR2X1_LOC_560/A 0.02fF
C3075 OR2X1_LOC_691/Y OR2X1_LOC_789/A 0.01fF
C3076 D_INPUT_0 AND2X1_LOC_839/a_8_24# 0.17fF
C3077 AND2X1_LOC_866/A OR2X1_LOC_755/Y 0.04fF
C3078 OR2X1_LOC_574/A OR2X1_LOC_592/a_8_216# 0.11fF
C3079 OR2X1_LOC_694/a_8_216# OR2X1_LOC_64/Y 0.01fF
C3080 AND2X1_LOC_40/Y OR2X1_LOC_244/A 0.07fF
C3081 OR2X1_LOC_68/B OR2X1_LOC_548/B 0.01fF
C3082 OR2X1_LOC_51/Y OR2X1_LOC_3/B 0.69fF
C3083 AND2X1_LOC_122/a_8_24# OR2X1_LOC_203/Y 0.01fF
C3084 AND2X1_LOC_560/B OR2X1_LOC_272/Y 0.09fF
C3085 AND2X1_LOC_206/Y AND2X1_LOC_206/a_36_24# 0.00fF
C3086 AND2X1_LOC_42/B OR2X1_LOC_83/A 0.02fF
C3087 OR2X1_LOC_31/Y AND2X1_LOC_642/Y 0.03fF
C3088 AND2X1_LOC_553/A OR2X1_LOC_95/Y 0.02fF
C3089 AND2X1_LOC_95/Y OR2X1_LOC_287/a_8_216# 0.02fF
C3090 OR2X1_LOC_593/B OR2X1_LOC_605/Y 0.08fF
C3091 OR2X1_LOC_417/Y OR2X1_LOC_603/a_36_216# 0.00fF
C3092 OR2X1_LOC_185/A OR2X1_LOC_471/Y 0.03fF
C3093 AND2X1_LOC_840/a_8_24# OR2X1_LOC_95/Y 0.01fF
C3094 AND2X1_LOC_523/Y OR2X1_LOC_44/Y 0.03fF
C3095 OR2X1_LOC_121/B AND2X1_LOC_29/a_8_24# 0.05fF
C3096 AND2X1_LOC_663/B AND2X1_LOC_361/A 0.10fF
C3097 OR2X1_LOC_185/A OR2X1_LOC_655/B 0.67fF
C3098 AND2X1_LOC_729/B OR2X1_LOC_52/B 0.15fF
C3099 AND2X1_LOC_366/A AND2X1_LOC_721/A 0.08fF
C3100 AND2X1_LOC_658/A OR2X1_LOC_406/A 0.19fF
C3101 OR2X1_LOC_506/A OR2X1_LOC_532/B 0.47fF
C3102 AND2X1_LOC_392/A OR2X1_LOC_331/Y 0.01fF
C3103 OR2X1_LOC_696/A OR2X1_LOC_387/A 0.02fF
C3104 OR2X1_LOC_272/a_8_216# OR2X1_LOC_272/Y 0.01fF
C3105 INPUT_1 OR2X1_LOC_265/Y 0.03fF
C3106 AND2X1_LOC_51/Y OR2X1_LOC_208/a_8_216# 0.06fF
C3107 AND2X1_LOC_647/B AND2X1_LOC_647/a_8_24# 0.01fF
C3108 AND2X1_LOC_729/Y OR2X1_LOC_679/A 0.01fF
C3109 AND2X1_LOC_656/Y OR2X1_LOC_118/Y 0.01fF
C3110 OR2X1_LOC_19/B AND2X1_LOC_472/B 0.05fF
C3111 OR2X1_LOC_787/B OR2X1_LOC_552/A 0.72fF
C3112 AND2X1_LOC_738/B OR2X1_LOC_331/a_36_216# 0.01fF
C3113 AND2X1_LOC_784/A OR2X1_LOC_46/A 0.07fF
C3114 OR2X1_LOC_185/A OR2X1_LOC_222/a_8_216# 0.01fF
C3115 OR2X1_LOC_12/Y AND2X1_LOC_247/a_8_24# 0.03fF
C3116 OR2X1_LOC_541/A OR2X1_LOC_723/A 0.01fF
C3117 AND2X1_LOC_48/A OR2X1_LOC_155/A 0.07fF
C3118 OR2X1_LOC_267/A OR2X1_LOC_720/B 0.03fF
C3119 AND2X1_LOC_21/a_36_24# AND2X1_LOC_21/Y 0.01fF
C3120 OR2X1_LOC_574/A AND2X1_LOC_491/a_36_24# 0.08fF
C3121 AND2X1_LOC_685/a_36_24# OR2X1_LOC_7/A 0.01fF
C3122 OR2X1_LOC_272/Y OR2X1_LOC_64/Y 0.05fF
C3123 AND2X1_LOC_509/a_8_24# AND2X1_LOC_657/A 0.01fF
C3124 OR2X1_LOC_111/Y OR2X1_LOC_6/A 0.16fF
C3125 OR2X1_LOC_56/A AND2X1_LOC_657/A 0.02fF
C3126 OR2X1_LOC_787/B OR2X1_LOC_578/B 0.07fF
C3127 AND2X1_LOC_576/Y OR2X1_LOC_226/Y 0.01fF
C3128 AND2X1_LOC_92/Y OR2X1_LOC_568/A 0.07fF
C3129 OR2X1_LOC_427/a_8_216# AND2X1_LOC_451/Y 0.49fF
C3130 OR2X1_LOC_233/a_8_216# OR2X1_LOC_54/Y 0.01fF
C3131 OR2X1_LOC_529/Y AND2X1_LOC_465/Y 0.00fF
C3132 AND2X1_LOC_436/a_8_24# OR2X1_LOC_331/Y 0.01fF
C3133 OR2X1_LOC_31/Y OR2X1_LOC_591/A 0.00fF
C3134 OR2X1_LOC_40/Y OR2X1_LOC_437/A 0.60fF
C3135 OR2X1_LOC_596/A AND2X1_LOC_41/Y 0.16fF
C3136 OR2X1_LOC_206/A OR2X1_LOC_206/a_8_216# 0.08fF
C3137 VDD OR2X1_LOC_446/B 0.13fF
C3138 AND2X1_LOC_348/Y AND2X1_LOC_866/A 0.68fF
C3139 OR2X1_LOC_510/Y OR2X1_LOC_473/A 0.04fF
C3140 OR2X1_LOC_662/a_36_216# AND2X1_LOC_31/Y 0.00fF
C3141 OR2X1_LOC_737/A OR2X1_LOC_374/Y 0.10fF
C3142 VDD OR2X1_LOC_303/B 0.08fF
C3143 OR2X1_LOC_401/A OR2X1_LOC_401/B 0.08fF
C3144 AND2X1_LOC_866/A OR2X1_LOC_753/A 0.07fF
C3145 OR2X1_LOC_251/Y AND2X1_LOC_859/B 0.00fF
C3146 OR2X1_LOC_63/a_36_216# OR2X1_LOC_67/Y 0.01fF
C3147 OR2X1_LOC_76/Y OR2X1_LOC_276/B 0.02fF
C3148 OR2X1_LOC_161/B OR2X1_LOC_356/B 0.08fF
C3149 AND2X1_LOC_359/B OR2X1_LOC_47/Y 0.15fF
C3150 OR2X1_LOC_53/Y OR2X1_LOC_304/a_8_216# 0.07fF
C3151 AND2X1_LOC_472/B OR2X1_LOC_838/B 0.12fF
C3152 OR2X1_LOC_42/a_8_216# D_INPUT_1 0.07fF
C3153 OR2X1_LOC_696/A AND2X1_LOC_542/a_8_24# 0.10fF
C3154 OR2X1_LOC_22/Y AND2X1_LOC_849/A 0.00fF
C3155 OR2X1_LOC_473/A OR2X1_LOC_810/A 0.29fF
C3156 OR2X1_LOC_375/A OR2X1_LOC_451/B 0.11fF
C3157 OR2X1_LOC_696/A AND2X1_LOC_713/a_36_24# 0.01fF
C3158 OR2X1_LOC_606/a_8_216# OR2X1_LOC_606/Y 0.00fF
C3159 AND2X1_LOC_110/Y OR2X1_LOC_308/Y 0.03fF
C3160 OR2X1_LOC_43/A OR2X1_LOC_597/Y 0.01fF
C3161 OR2X1_LOC_64/Y AND2X1_LOC_801/B 0.00fF
C3162 OR2X1_LOC_696/A OR2X1_LOC_9/Y 1.74fF
C3163 OR2X1_LOC_743/A OR2X1_LOC_760/Y 0.09fF
C3164 AND2X1_LOC_313/a_36_24# OR2X1_LOC_308/Y 0.01fF
C3165 OR2X1_LOC_816/A OR2X1_LOC_530/a_36_216# 0.00fF
C3166 AND2X1_LOC_56/B OR2X1_LOC_192/B 0.09fF
C3167 OR2X1_LOC_47/Y AND2X1_LOC_639/a_8_24# 0.01fF
C3168 OR2X1_LOC_624/A OR2X1_LOC_68/B 0.01fF
C3169 AND2X1_LOC_555/Y AND2X1_LOC_555/a_8_24# 0.02fF
C3170 AND2X1_LOC_166/a_8_24# OR2X1_LOC_568/A 0.02fF
C3171 OR2X1_LOC_112/a_8_216# OR2X1_LOC_175/Y 0.01fF
C3172 AND2X1_LOC_64/Y OR2X1_LOC_362/A 0.22fF
C3173 AND2X1_LOC_810/A OR2X1_LOC_428/A 0.06fF
C3174 OR2X1_LOC_78/B AND2X1_LOC_36/Y 0.44fF
C3175 OR2X1_LOC_113/a_36_216# OR2X1_LOC_113/B 0.00fF
C3176 AND2X1_LOC_802/Y AND2X1_LOC_809/a_8_24# 0.03fF
C3177 OR2X1_LOC_70/A OR2X1_LOC_588/Y 0.02fF
C3178 AND2X1_LOC_721/Y OR2X1_LOC_158/A 0.27fF
C3179 AND2X1_LOC_22/Y OR2X1_LOC_596/A 0.01fF
C3180 AND2X1_LOC_28/a_8_24# D_INPUT_0 0.04fF
C3181 AND2X1_LOC_817/B AND2X1_LOC_236/a_8_24# 0.01fF
C3182 OR2X1_LOC_62/A OR2X1_LOC_46/A 0.50fF
C3183 OR2X1_LOC_19/B OR2X1_LOC_838/B 0.01fF
C3184 AND2X1_LOC_714/a_8_24# AND2X1_LOC_714/B 0.00fF
C3185 OR2X1_LOC_138/a_8_216# OR2X1_LOC_160/B 0.06fF
C3186 OR2X1_LOC_70/Y OR2X1_LOC_86/A 0.50fF
C3187 OR2X1_LOC_810/A OR2X1_LOC_228/Y 0.07fF
C3188 AND2X1_LOC_687/A AND2X1_LOC_687/a_8_24# 0.10fF
C3189 AND2X1_LOC_403/B OR2X1_LOC_399/Y 0.13fF
C3190 AND2X1_LOC_866/A AND2X1_LOC_845/Y 0.07fF
C3191 OR2X1_LOC_433/Y OR2X1_LOC_589/a_36_216# -0.00fF
C3192 AND2X1_LOC_436/B OR2X1_LOC_589/a_8_216# 0.47fF
C3193 OR2X1_LOC_66/A OR2X1_LOC_563/A 0.07fF
C3194 OR2X1_LOC_478/Y VDD -0.00fF
C3195 OR2X1_LOC_405/A OR2X1_LOC_730/B 0.07fF
C3196 OR2X1_LOC_223/A OR2X1_LOC_814/A 0.03fF
C3197 AND2X1_LOC_40/Y OR2X1_LOC_731/B 0.11fF
C3198 VDD OR2X1_LOC_366/B 0.06fF
C3199 D_INPUT_4 INPUT_6 0.90fF
C3200 AND2X1_LOC_860/A OR2X1_LOC_428/A 0.00fF
C3201 OR2X1_LOC_555/A OR2X1_LOC_259/B 0.09fF
C3202 OR2X1_LOC_307/A OR2X1_LOC_713/A 0.03fF
C3203 OR2X1_LOC_45/B AND2X1_LOC_508/B 0.03fF
C3204 OR2X1_LOC_121/B OR2X1_LOC_493/Y 0.26fF
C3205 OR2X1_LOC_663/a_8_216# OR2X1_LOC_772/A 0.40fF
C3206 OR2X1_LOC_158/A OR2X1_LOC_482/Y 0.03fF
C3207 OR2X1_LOC_536/Y OR2X1_LOC_16/A 0.01fF
C3208 AND2X1_LOC_340/a_8_24# OR2X1_LOC_595/A 0.20fF
C3209 OR2X1_LOC_532/B AND2X1_LOC_420/a_8_24# 0.00fF
C3210 INPUT_0 AND2X1_LOC_829/a_8_24# 0.01fF
C3211 OR2X1_LOC_190/A AND2X1_LOC_279/a_8_24# 0.00fF
C3212 OR2X1_LOC_532/B D_INPUT_1 0.11fF
C3213 AND2X1_LOC_64/Y OR2X1_LOC_474/Y 1.26fF
C3214 AND2X1_LOC_788/a_8_24# OR2X1_LOC_600/A 0.02fF
C3215 OR2X1_LOC_609/A OR2X1_LOC_71/A 0.02fF
C3216 OR2X1_LOC_520/Y OR2X1_LOC_771/B 0.01fF
C3217 AND2X1_LOC_643/a_8_24# OR2X1_LOC_46/A 0.01fF
C3218 AND2X1_LOC_95/Y OR2X1_LOC_333/A 0.01fF
C3219 OR2X1_LOC_750/A OR2X1_LOC_358/A 0.07fF
C3220 OR2X1_LOC_143/a_8_216# INPUT_3 0.01fF
C3221 OR2X1_LOC_51/Y OR2X1_LOC_584/a_8_216# 0.01fF
C3222 OR2X1_LOC_375/A AND2X1_LOC_36/Y 8.48fF
C3223 AND2X1_LOC_362/B OR2X1_LOC_600/A 0.07fF
C3224 AND2X1_LOC_474/A AND2X1_LOC_244/A 1.37fF
C3225 OR2X1_LOC_600/A AND2X1_LOC_476/Y 0.07fF
C3226 OR2X1_LOC_311/Y OR2X1_LOC_761/a_8_216# 0.02fF
C3227 VDD OR2X1_LOC_719/B 0.17fF
C3228 OR2X1_LOC_769/A AND2X1_LOC_585/a_8_24# 0.09fF
C3229 OR2X1_LOC_204/a_8_216# OR2X1_LOC_71/A 0.09fF
C3230 AND2X1_LOC_22/Y OR2X1_LOC_808/A 0.05fF
C3231 OR2X1_LOC_814/A OR2X1_LOC_351/a_36_216# 0.00fF
C3232 OR2X1_LOC_7/A OR2X1_LOC_437/A 2.05fF
C3233 AND2X1_LOC_322/a_8_24# OR2X1_LOC_325/B 0.01fF
C3234 AND2X1_LOC_738/B AND2X1_LOC_794/B 0.03fF
C3235 OR2X1_LOC_106/a_8_216# OR2X1_LOC_426/B 0.02fF
C3236 OR2X1_LOC_696/A AND2X1_LOC_572/Y 0.03fF
C3237 AND2X1_LOC_677/a_8_24# OR2X1_LOC_779/B 0.01fF
C3238 OR2X1_LOC_40/Y AND2X1_LOC_715/A 0.03fF
C3239 OR2X1_LOC_323/A AND2X1_LOC_662/B 0.03fF
C3240 AND2X1_LOC_352/a_8_24# AND2X1_LOC_352/B 0.00fF
C3241 OR2X1_LOC_54/Y OR2X1_LOC_68/B 0.10fF
C3242 OR2X1_LOC_364/B OR2X1_LOC_756/B 0.00fF
C3243 OR2X1_LOC_118/Y AND2X1_LOC_772/Y 0.01fF
C3244 AND2X1_LOC_719/Y OR2X1_LOC_59/Y 1.05fF
C3245 VDD OR2X1_LOC_542/B 0.07fF
C3246 OR2X1_LOC_658/a_36_216# OR2X1_LOC_113/B 0.00fF
C3247 OR2X1_LOC_506/Y OR2X1_LOC_721/Y 0.06fF
C3248 AND2X1_LOC_51/Y OR2X1_LOC_728/A 0.04fF
C3249 OR2X1_LOC_40/Y AND2X1_LOC_851/a_8_24# 0.02fF
C3250 AND2X1_LOC_95/Y OR2X1_LOC_392/B 0.08fF
C3251 AND2X1_LOC_738/B VDD 1.29fF
C3252 OR2X1_LOC_186/Y OR2X1_LOC_330/Y 0.12fF
C3253 OR2X1_LOC_6/B AND2X1_LOC_14/a_36_24# 0.01fF
C3254 VDD OR2X1_LOC_56/A 1.17fF
C3255 AND2X1_LOC_543/a_8_24# AND2X1_LOC_476/Y 0.03fF
C3256 OR2X1_LOC_9/Y AND2X1_LOC_819/a_8_24# 0.01fF
C3257 OR2X1_LOC_486/a_8_216# OR2X1_LOC_550/B 0.06fF
C3258 OR2X1_LOC_328/a_36_216# OR2X1_LOC_40/Y 0.00fF
C3259 AND2X1_LOC_710/Y VDD 0.11fF
C3260 AND2X1_LOC_706/Y OR2X1_LOC_92/Y 0.10fF
C3261 AND2X1_LOC_64/Y OR2X1_LOC_217/Y 0.03fF
C3262 OR2X1_LOC_696/A AND2X1_LOC_852/Y 0.01fF
C3263 AND2X1_LOC_231/Y OR2X1_LOC_18/Y 0.28fF
C3264 VDD OR2X1_LOC_819/a_8_216# 0.00fF
C3265 VDD OR2X1_LOC_573/a_8_216# 0.21fF
C3266 AND2X1_LOC_227/Y OR2X1_LOC_88/Y 0.24fF
C3267 AND2X1_LOC_841/B AND2X1_LOC_810/B 0.07fF
C3268 OR2X1_LOC_696/A OR2X1_LOC_6/a_36_216# 0.00fF
C3269 OR2X1_LOC_516/Y OR2X1_LOC_529/Y 0.03fF
C3270 AND2X1_LOC_40/Y OR2X1_LOC_180/a_8_216# 0.01fF
C3271 AND2X1_LOC_564/B OR2X1_LOC_406/a_36_216# 0.01fF
C3272 OR2X1_LOC_427/A OR2X1_LOC_604/Y 0.01fF
C3273 AND2X1_LOC_706/a_8_24# OR2X1_LOC_48/B 0.03fF
C3274 OR2X1_LOC_687/Y AND2X1_LOC_7/B 0.07fF
C3275 AND2X1_LOC_91/B OR2X1_LOC_845/a_36_216# 0.00fF
C3276 OR2X1_LOC_97/A OR2X1_LOC_130/A 0.12fF
C3277 OR2X1_LOC_199/a_36_216# OR2X1_LOC_375/A 0.02fF
C3278 OR2X1_LOC_589/A OR2X1_LOC_48/B 0.35fF
C3279 AND2X1_LOC_59/Y OR2X1_LOC_161/B 0.18fF
C3280 AND2X1_LOC_341/a_8_24# OR2X1_LOC_265/Y 0.02fF
C3281 OR2X1_LOC_632/a_8_216# OR2X1_LOC_78/A 0.01fF
C3282 VDD AND2X1_LOC_638/Y -0.00fF
C3283 AND2X1_LOC_706/a_8_24# OR2X1_LOC_18/Y 0.04fF
C3284 AND2X1_LOC_121/a_8_24# AND2X1_LOC_474/A 0.01fF
C3285 OR2X1_LOC_666/A AND2X1_LOC_860/a_8_24# 0.20fF
C3286 OR2X1_LOC_756/B AND2X1_LOC_70/Y 1.42fF
C3287 VDD OR2X1_LOC_736/A 0.03fF
C3288 OR2X1_LOC_39/A OR2X1_LOC_373/Y 0.05fF
C3289 OR2X1_LOC_47/Y AND2X1_LOC_790/a_8_24# 0.02fF
C3290 AND2X1_LOC_95/Y OR2X1_LOC_113/B 0.23fF
C3291 OR2X1_LOC_306/Y AND2X1_LOC_774/A 0.00fF
C3292 OR2X1_LOC_506/Y OR2X1_LOC_375/A 0.01fF
C3293 AND2X1_LOC_83/a_8_24# AND2X1_LOC_617/a_8_24# 0.23fF
C3294 OR2X1_LOC_589/A OR2X1_LOC_18/Y 0.20fF
C3295 AND2X1_LOC_624/A AND2X1_LOC_212/Y 0.07fF
C3296 OR2X1_LOC_851/B OR2X1_LOC_185/A 0.24fF
C3297 OR2X1_LOC_633/a_8_216# OR2X1_LOC_78/B 0.01fF
C3298 OR2X1_LOC_633/a_36_216# OR2X1_LOC_78/A 0.00fF
C3299 AND2X1_LOC_738/B OR2X1_LOC_677/Y 0.08fF
C3300 OR2X1_LOC_152/Y AND2X1_LOC_209/Y 0.01fF
C3301 OR2X1_LOC_456/a_36_216# OR2X1_LOC_549/A 0.00fF
C3302 OR2X1_LOC_9/Y OR2X1_LOC_823/a_36_216# 0.00fF
C3303 OR2X1_LOC_201/A OR2X1_LOC_78/A 0.04fF
C3304 VDD OR2X1_LOC_426/Y 0.12fF
C3305 OR2X1_LOC_36/Y AND2X1_LOC_786/Y 0.07fF
C3306 OR2X1_LOC_85/A OR2X1_LOC_16/A 0.06fF
C3307 OR2X1_LOC_856/B OR2X1_LOC_389/A 0.07fF
C3308 OR2X1_LOC_526/Y OR2X1_LOC_525/Y 0.07fF
C3309 OR2X1_LOC_346/a_8_216# OR2X1_LOC_346/A 0.05fF
C3310 VDD OR2X1_LOC_631/a_8_216# 0.00fF
C3311 AND2X1_LOC_425/Y INPUT_6 0.03fF
C3312 OR2X1_LOC_635/A OR2X1_LOC_78/B 0.01fF
C3313 OR2X1_LOC_224/a_8_216# OR2X1_LOC_437/A 0.01fF
C3314 VDD AND2X1_LOC_850/Y 0.21fF
C3315 OR2X1_LOC_756/B OR2X1_LOC_703/A 0.03fF
C3316 OR2X1_LOC_857/B OR2X1_LOC_836/A 0.79fF
C3317 OR2X1_LOC_559/B AND2X1_LOC_18/Y 0.01fF
C3318 OR2X1_LOC_45/B AND2X1_LOC_339/a_8_24# 0.01fF
C3319 AND2X1_LOC_541/a_8_24# OR2X1_LOC_272/Y 0.00fF
C3320 AND2X1_LOC_724/a_36_24# OR2X1_LOC_485/A 0.00fF
C3321 AND2X1_LOC_711/Y AND2X1_LOC_580/a_8_24# 0.01fF
C3322 AND2X1_LOC_776/Y OR2X1_LOC_64/Y 0.20fF
C3323 OR2X1_LOC_91/Y AND2X1_LOC_722/a_8_24# -0.00fF
C3324 AND2X1_LOC_22/Y OR2X1_LOC_33/B 0.09fF
C3325 OR2X1_LOC_585/A AND2X1_LOC_415/a_8_24# 0.03fF
C3326 OR2X1_LOC_160/B AND2X1_LOC_43/B 0.14fF
C3327 AND2X1_LOC_865/A AND2X1_LOC_805/Y 0.08fF
C3328 OR2X1_LOC_158/A OR2X1_LOC_748/A 0.03fF
C3329 OR2X1_LOC_744/A OR2X1_LOC_427/A 0.23fF
C3330 OR2X1_LOC_137/B OR2X1_LOC_66/A 0.03fF
C3331 OR2X1_LOC_429/Y INPUT_7 0.17fF
C3332 OR2X1_LOC_528/Y AND2X1_LOC_564/a_8_24# 0.01fF
C3333 AND2X1_LOC_348/A OR2X1_LOC_494/a_8_216# 0.00fF
C3334 OR2X1_LOC_663/a_8_216# AND2X1_LOC_3/Y 0.03fF
C3335 AND2X1_LOC_104/a_8_24# OR2X1_LOC_78/A 0.03fF
C3336 OR2X1_LOC_40/Y AND2X1_LOC_348/Y 0.01fF
C3337 OR2X1_LOC_720/A AND2X1_LOC_18/Y 0.02fF
C3338 AND2X1_LOC_595/a_36_24# OR2X1_LOC_154/A 0.01fF
C3339 OR2X1_LOC_477/Y OR2X1_LOC_469/Y 0.19fF
C3340 OR2X1_LOC_368/a_36_216# OR2X1_LOC_44/Y 0.02fF
C3341 AND2X1_LOC_723/Y AND2X1_LOC_723/a_8_24# 0.04fF
C3342 OR2X1_LOC_589/A OR2X1_LOC_385/Y 0.01fF
C3343 OR2X1_LOC_210/a_8_216# OR2X1_LOC_803/A 0.01fF
C3344 OR2X1_LOC_847/A OR2X1_LOC_78/Y 0.03fF
C3345 OR2X1_LOC_40/Y OR2X1_LOC_753/A 0.03fF
C3346 AND2X1_LOC_392/A AND2X1_LOC_170/Y 0.17fF
C3347 VDD AND2X1_LOC_56/B 1.30fF
C3348 OR2X1_LOC_604/A OR2X1_LOC_669/a_8_216# 0.10fF
C3349 AND2X1_LOC_842/B AND2X1_LOC_242/a_8_24# 0.01fF
C3350 VDD OR2X1_LOC_659/B 0.18fF
C3351 AND2X1_LOC_392/A AND2X1_LOC_361/A 0.07fF
C3352 AND2X1_LOC_799/a_8_24# AND2X1_LOC_727/A 0.01fF
C3353 AND2X1_LOC_480/A AND2X1_LOC_220/Y 0.05fF
C3354 AND2X1_LOC_81/a_36_24# OR2X1_LOC_786/A 0.00fF
C3355 AND2X1_LOC_12/Y OR2X1_LOC_630/B 0.01fF
C3356 AND2X1_LOC_714/B OR2X1_LOC_743/A 0.03fF
C3357 OR2X1_LOC_653/A OR2X1_LOC_648/A 0.08fF
C3358 AND2X1_LOC_576/Y OR2X1_LOC_51/Y 0.00fF
C3359 INPUT_0 OR2X1_LOC_828/B 0.07fF
C3360 OR2X1_LOC_157/a_8_216# OR2X1_LOC_25/Y 0.02fF
C3361 VDD AND2X1_LOC_8/Y 0.62fF
C3362 OR2X1_LOC_161/A OR2X1_LOC_735/a_8_216# 0.01fF
C3363 OR2X1_LOC_574/A OR2X1_LOC_730/A 0.15fF
C3364 OR2X1_LOC_160/A OR2X1_LOC_114/a_36_216# 0.01fF
C3365 OR2X1_LOC_231/A OR2X1_LOC_475/B 0.13fF
C3366 OR2X1_LOC_421/A OR2X1_LOC_764/Y 0.01fF
C3367 OR2X1_LOC_633/a_8_216# OR2X1_LOC_375/A 0.01fF
C3368 OR2X1_LOC_791/B OR2X1_LOC_756/B 0.03fF
C3369 AND2X1_LOC_191/B OR2X1_LOC_44/Y 0.07fF
C3370 AND2X1_LOC_654/B OR2X1_LOC_48/B 0.02fF
C3371 OR2X1_LOC_36/Y AND2X1_LOC_218/Y 0.02fF
C3372 OR2X1_LOC_528/Y OR2X1_LOC_74/A 10.35fF
C3373 OR2X1_LOC_348/Y OR2X1_LOC_287/B 0.02fF
C3374 AND2X1_LOC_729/B OR2X1_LOC_13/a_8_216# 0.01fF
C3375 OR2X1_LOC_81/a_8_216# OR2X1_LOC_59/Y 0.07fF
C3376 OR2X1_LOC_6/B AND2X1_LOC_42/B 1.13fF
C3377 OR2X1_LOC_18/Y AND2X1_LOC_654/B 0.01fF
C3378 OR2X1_LOC_40/Y AND2X1_LOC_243/a_8_24# 0.01fF
C3379 OR2X1_LOC_349/a_8_216# OR2X1_LOC_287/B 0.01fF
C3380 AND2X1_LOC_729/Y AND2X1_LOC_722/A 0.07fF
C3381 VDD AND2X1_LOC_21/Y 0.53fF
C3382 OR2X1_LOC_333/B AND2X1_LOC_18/Y 0.03fF
C3383 AND2X1_LOC_724/Y OR2X1_LOC_89/A 0.02fF
C3384 OR2X1_LOC_251/Y OR2X1_LOC_56/A 0.07fF
C3385 OR2X1_LOC_18/Y OR2X1_LOC_495/Y 0.03fF
C3386 AND2X1_LOC_722/a_36_24# OR2X1_LOC_74/A 0.01fF
C3387 OR2X1_LOC_811/A OR2X1_LOC_833/B 0.03fF
C3388 AND2X1_LOC_48/A OR2X1_LOC_706/a_36_216# 0.00fF
C3389 OR2X1_LOC_95/Y AND2X1_LOC_465/A 1.81fF
C3390 OR2X1_LOC_635/A OR2X1_LOC_375/A 0.07fF
C3391 VDD AND2X1_LOC_641/Y 0.21fF
C3392 OR2X1_LOC_411/Y OR2X1_LOC_7/A 0.03fF
C3393 AND2X1_LOC_512/a_8_24# AND2X1_LOC_434/Y 0.01fF
C3394 OR2X1_LOC_530/Y AND2X1_LOC_658/A 0.03fF
C3395 VDD OR2X1_LOC_291/A 0.03fF
C3396 OR2X1_LOC_130/A OR2X1_LOC_475/B 0.03fF
C3397 AND2X1_LOC_59/Y OR2X1_LOC_61/Y 0.03fF
C3398 OR2X1_LOC_609/A OR2X1_LOC_59/Y 0.00fF
C3399 AND2X1_LOC_95/Y OR2X1_LOC_286/Y -0.00fF
C3400 AND2X1_LOC_568/B AND2X1_LOC_212/B 0.01fF
C3401 AND2X1_LOC_772/B OR2X1_LOC_490/Y 0.01fF
C3402 AND2X1_LOC_3/Y OR2X1_LOC_78/A 5.41fF
C3403 OR2X1_LOC_274/Y OR2X1_LOC_203/Y 0.02fF
C3404 OR2X1_LOC_647/B OR2X1_LOC_78/A 0.19fF
C3405 OR2X1_LOC_11/Y OR2X1_LOC_59/a_8_216# 0.01fF
C3406 AND2X1_LOC_784/A AND2X1_LOC_722/A 0.07fF
C3407 OR2X1_LOC_528/a_8_216# AND2X1_LOC_574/A 0.48fF
C3408 OR2X1_LOC_18/Y AND2X1_LOC_858/a_8_24# 0.02fF
C3409 AND2X1_LOC_99/A AND2X1_LOC_123/Y 0.01fF
C3410 OR2X1_LOC_160/A OR2X1_LOC_185/A 0.31fF
C3411 AND2X1_LOC_73/a_8_24# AND2X1_LOC_42/B 0.09fF
C3412 AND2X1_LOC_59/Y AND2X1_LOC_536/a_8_24# 0.01fF
C3413 OR2X1_LOC_100/Y OR2X1_LOC_99/Y 0.00fF
C3414 OR2X1_LOC_227/a_36_216# OR2X1_LOC_641/A 0.02fF
C3415 AND2X1_LOC_576/a_8_24# AND2X1_LOC_573/A 0.02fF
C3416 OR2X1_LOC_826/a_8_216# OR2X1_LOC_56/A 0.04fF
C3417 OR2X1_LOC_151/A D_INPUT_0 0.27fF
C3418 OR2X1_LOC_147/B OR2X1_LOC_464/B 0.11fF
C3419 OR2X1_LOC_427/A AND2X1_LOC_840/B 0.10fF
C3420 AND2X1_LOC_81/B AND2X1_LOC_504/a_8_24# 0.01fF
C3421 OR2X1_LOC_786/Y AND2X1_LOC_7/B 0.10fF
C3422 OR2X1_LOC_797/B OR2X1_LOC_797/A 0.11fF
C3423 OR2X1_LOC_97/A AND2X1_LOC_438/a_36_24# 0.00fF
C3424 OR2X1_LOC_865/A D_INPUT_1 0.09fF
C3425 OR2X1_LOC_346/a_8_216# OR2X1_LOC_161/A 0.01fF
C3426 OR2X1_LOC_43/A OR2X1_LOC_48/B 0.32fF
C3427 AND2X1_LOC_76/Y AND2X1_LOC_264/a_8_24# 0.01fF
C3428 OR2X1_LOC_385/Y AND2X1_LOC_654/B 0.29fF
C3429 AND2X1_LOC_359/B OR2X1_LOC_625/Y 0.70fF
C3430 OR2X1_LOC_3/Y OR2X1_LOC_256/Y 0.03fF
C3431 OR2X1_LOC_8/Y OR2X1_LOC_46/A 0.23fF
C3432 AND2X1_LOC_97/a_36_24# OR2X1_LOC_44/Y 0.01fF
C3433 AND2X1_LOC_350/Y OR2X1_LOC_59/Y 0.03fF
C3434 OR2X1_LOC_485/A OR2X1_LOC_92/Y 0.24fF
C3435 OR2X1_LOC_429/Y OR2X1_LOC_426/A 0.05fF
C3436 AND2X1_LOC_22/Y OR2X1_LOC_795/a_8_216# 0.01fF
C3437 OR2X1_LOC_43/A OR2X1_LOC_18/Y 0.25fF
C3438 OR2X1_LOC_449/B AND2X1_LOC_426/a_8_24# 0.01fF
C3439 AND2X1_LOC_729/Y OR2X1_LOC_599/A 0.11fF
C3440 AND2X1_LOC_576/Y OR2X1_LOC_680/A 0.07fF
C3441 AND2X1_LOC_528/a_8_24# OR2X1_LOC_220/B 0.01fF
C3442 OR2X1_LOC_32/B OR2X1_LOC_26/Y 0.34fF
C3443 OR2X1_LOC_520/Y OR2X1_LOC_642/a_8_216# 0.01fF
C3444 AND2X1_LOC_22/Y OR2X1_LOC_374/Y 0.03fF
C3445 AND2X1_LOC_42/B OR2X1_LOC_523/Y 0.01fF
C3446 OR2X1_LOC_711/A OR2X1_LOC_738/A 0.13fF
C3447 OR2X1_LOC_307/a_36_216# OR2X1_LOC_161/A 0.01fF
C3448 OR2X1_LOC_280/Y OR2X1_LOC_109/Y 0.02fF
C3449 OR2X1_LOC_97/A OR2X1_LOC_365/B 0.02fF
C3450 OR2X1_LOC_106/A OR2X1_LOC_67/A 0.02fF
C3451 OR2X1_LOC_185/A AND2X1_LOC_86/B 0.01fF
C3452 OR2X1_LOC_600/a_8_216# OR2X1_LOC_95/Y 0.01fF
C3453 OR2X1_LOC_419/Y AND2X1_LOC_786/Y 0.10fF
C3454 AND2X1_LOC_345/a_8_24# AND2X1_LOC_847/Y 0.02fF
C3455 AND2X1_LOC_719/Y OR2X1_LOC_184/Y 0.31fF
C3456 OR2X1_LOC_485/A OR2X1_LOC_65/B 0.09fF
C3457 OR2X1_LOC_125/a_8_216# D_INPUT_3 0.00fF
C3458 AND2X1_LOC_36/Y OR2X1_LOC_515/Y 0.01fF
C3459 OR2X1_LOC_479/Y OR2X1_LOC_161/A 0.16fF
C3460 OR2X1_LOC_391/B OR2X1_LOC_864/A 0.01fF
C3461 OR2X1_LOC_512/a_8_216# OR2X1_LOC_713/A 0.01fF
C3462 OR2X1_LOC_316/Y AND2X1_LOC_640/Y 0.01fF
C3463 AND2X1_LOC_316/a_36_24# OR2X1_LOC_206/A 0.00fF
C3464 AND2X1_LOC_703/a_8_24# OR2X1_LOC_64/Y 0.01fF
C3465 OR2X1_LOC_246/a_36_216# OR2X1_LOC_753/A 0.01fF
C3466 INPUT_4 OR2X1_LOC_429/Y 0.01fF
C3467 OR2X1_LOC_391/B OR2X1_LOC_774/Y 0.25fF
C3468 AND2X1_LOC_638/a_8_24# OR2X1_LOC_44/Y 0.00fF
C3469 AND2X1_LOC_264/a_8_24# OR2X1_LOC_52/B 0.03fF
C3470 OR2X1_LOC_70/Y OR2X1_LOC_313/Y 0.01fF
C3471 AND2X1_LOC_348/Y OR2X1_LOC_7/A 0.08fF
C3472 AND2X1_LOC_12/Y AND2X1_LOC_67/Y 0.03fF
C3473 OR2X1_LOC_502/A OR2X1_LOC_814/A 0.13fF
C3474 AND2X1_LOC_122/a_8_24# OR2X1_LOC_375/A 0.01fF
C3475 AND2X1_LOC_42/B OR2X1_LOC_579/B 0.01fF
C3476 OR2X1_LOC_64/Y AND2X1_LOC_468/B 3.57fF
C3477 OR2X1_LOC_260/Y OR2X1_LOC_345/A 0.01fF
C3478 OR2X1_LOC_47/Y AND2X1_LOC_436/Y 0.03fF
C3479 AND2X1_LOC_744/a_8_24# OR2X1_LOC_780/B 0.27fF
C3480 OR2X1_LOC_121/B AND2X1_LOC_426/a_8_24# 0.03fF
C3481 OR2X1_LOC_154/A AND2X1_LOC_69/Y 0.02fF
C3482 OR2X1_LOC_7/A OR2X1_LOC_753/A 0.10fF
C3483 AND2X1_LOC_756/a_8_24# GATE_662 0.01fF
C3484 OR2X1_LOC_837/a_8_216# OR2X1_LOC_46/A 0.01fF
C3485 OR2X1_LOC_287/B OR2X1_LOC_810/A 0.05fF
C3486 OR2X1_LOC_683/Y AND2X1_LOC_452/Y 0.01fF
C3487 OR2X1_LOC_223/A OR2X1_LOC_192/A 0.00fF
C3488 OR2X1_LOC_277/a_8_216# OR2X1_LOC_39/A 0.01fF
C3489 AND2X1_LOC_580/A OR2X1_LOC_617/Y 0.02fF
C3490 OR2X1_LOC_26/Y OR2X1_LOC_371/Y 0.07fF
C3491 AND2X1_LOC_3/Y OR2X1_LOC_155/A 0.15fF
C3492 OR2X1_LOC_316/Y OR2X1_LOC_416/Y 2.98fF
C3493 AND2X1_LOC_31/Y AND2X1_LOC_65/A 0.02fF
C3494 OR2X1_LOC_7/A OR2X1_LOC_754/a_8_216# 0.03fF
C3495 OR2X1_LOC_426/A OR2X1_LOC_428/a_8_216# 0.01fF
C3496 AND2X1_LOC_46/a_36_24# OR2X1_LOC_375/A 0.00fF
C3497 OR2X1_LOC_532/B OR2X1_LOC_737/A 0.09fF
C3498 OR2X1_LOC_814/A OR2X1_LOC_571/B 0.02fF
C3499 OR2X1_LOC_185/A OR2X1_LOC_655/A 0.02fF
C3500 AND2X1_LOC_624/B OR2X1_LOC_56/A 0.00fF
C3501 AND2X1_LOC_64/Y OR2X1_LOC_771/B 0.03fF
C3502 OR2X1_LOC_89/A OR2X1_LOC_371/Y 0.07fF
C3503 OR2X1_LOC_715/B OR2X1_LOC_228/Y 0.10fF
C3504 OR2X1_LOC_835/A OR2X1_LOC_19/B 0.04fF
C3505 AND2X1_LOC_95/Y OR2X1_LOC_532/B 3.08fF
C3506 OR2X1_LOC_31/Y OR2X1_LOC_427/A 1.92fF
C3507 OR2X1_LOC_391/A D_INPUT_1 0.25fF
C3508 OR2X1_LOC_646/a_36_216# OR2X1_LOC_647/A 0.00fF
C3509 AND2X1_LOC_154/Y AND2X1_LOC_155/Y 0.22fF
C3510 OR2X1_LOC_633/Y OR2X1_LOC_532/B 0.01fF
C3511 AND2X1_LOC_63/a_8_24# OR2X1_LOC_62/B 0.01fF
C3512 AND2X1_LOC_486/a_8_24# AND2X1_LOC_468/a_8_24# 0.23fF
C3513 AND2X1_LOC_344/a_8_24# OR2X1_LOC_47/Y 0.02fF
C3514 OR2X1_LOC_715/B OR2X1_LOC_513/Y 0.00fF
C3515 AND2X1_LOC_56/B OR2X1_LOC_444/B 0.01fF
C3516 OR2X1_LOC_404/Y AND2X1_LOC_159/a_36_24# 0.00fF
C3517 OR2X1_LOC_78/A OR2X1_LOC_196/a_36_216# 0.00fF
C3518 OR2X1_LOC_490/Y AND2X1_LOC_141/B 0.02fF
C3519 OR2X1_LOC_147/B OR2X1_LOC_223/A 0.03fF
C3520 OR2X1_LOC_864/A OR2X1_LOC_772/Y 0.00fF
C3521 D_INPUT_7 AND2X1_LOC_1/Y 0.01fF
C3522 AND2X1_LOC_520/Y AND2X1_LOC_476/A 0.04fF
C3523 OR2X1_LOC_787/a_36_216# OR2X1_LOC_578/B 0.02fF
C3524 AND2X1_LOC_64/Y OR2X1_LOC_776/A 0.03fF
C3525 OR2X1_LOC_487/a_8_216# OR2X1_LOC_488/Y 0.40fF
C3526 AND2X1_LOC_866/B AND2X1_LOC_620/Y 0.02fF
C3527 AND2X1_LOC_661/A AND2X1_LOC_802/a_36_24# 0.00fF
C3528 AND2X1_LOC_832/a_8_24# AND2X1_LOC_648/B 0.01fF
C3529 OR2X1_LOC_59/Y OR2X1_LOC_331/a_8_216# 0.01fF
C3530 AND2X1_LOC_708/a_36_24# OR2X1_LOC_52/B 0.01fF
C3531 OR2X1_LOC_774/Y OR2X1_LOC_772/Y 0.17fF
C3532 OR2X1_LOC_756/B OR2X1_LOC_544/a_36_216# 0.00fF
C3533 OR2X1_LOC_774/Y OR2X1_LOC_846/A 0.74fF
C3534 OR2X1_LOC_96/B OR2X1_LOC_54/a_8_216# 0.01fF
C3535 OR2X1_LOC_46/A OR2X1_LOC_52/B 0.03fF
C3536 OR2X1_LOC_672/Y OR2X1_LOC_46/A 0.01fF
C3537 OR2X1_LOC_479/Y AND2X1_LOC_51/Y 0.10fF
C3538 OR2X1_LOC_273/Y OR2X1_LOC_275/A 0.01fF
C3539 OR2X1_LOC_291/Y OR2X1_LOC_609/a_8_216# 0.02fF
C3540 OR2X1_LOC_66/A OR2X1_LOC_724/A 0.07fF
C3541 INPUT_4 OR2X1_LOC_428/a_8_216# 0.00fF
C3542 OR2X1_LOC_79/A OR2X1_LOC_64/Y 0.01fF
C3543 AND2X1_LOC_681/a_8_24# OR2X1_LOC_161/A 0.01fF
C3544 AND2X1_LOC_658/B OR2X1_LOC_152/a_8_216# 0.06fF
C3545 OR2X1_LOC_377/A AND2X1_LOC_827/a_8_24# 0.03fF
C3546 OR2X1_LOC_62/a_36_216# OR2X1_LOC_585/A 0.00fF
C3547 OR2X1_LOC_70/Y AND2X1_LOC_350/Y 0.03fF
C3548 OR2X1_LOC_74/A OR2X1_LOC_54/Y 0.02fF
C3549 AND2X1_LOC_22/Y OR2X1_LOC_333/A 0.20fF
C3550 OR2X1_LOC_532/B OR2X1_LOC_99/Y 0.00fF
C3551 OR2X1_LOC_73/a_36_216# OR2X1_LOC_46/A 0.00fF
C3552 D_INPUT_3 AND2X1_LOC_852/a_8_24# 0.00fF
C3553 OR2X1_LOC_805/A OR2X1_LOC_786/Y 0.10fF
C3554 OR2X1_LOC_743/A AND2X1_LOC_477/A 0.03fF
C3555 AND2X1_LOC_727/Y AND2X1_LOC_544/Y 0.03fF
C3556 OR2X1_LOC_147/B OR2X1_LOC_705/B 0.02fF
C3557 OR2X1_LOC_696/A AND2X1_LOC_787/A 0.01fF
C3558 AND2X1_LOC_784/A AND2X1_LOC_866/A 0.07fF
C3559 AND2X1_LOC_36/Y OR2X1_LOC_549/A 0.29fF
C3560 OR2X1_LOC_436/Y OR2X1_LOC_810/A 0.23fF
C3561 AND2X1_LOC_387/B AND2X1_LOC_53/Y 0.07fF
C3562 OR2X1_LOC_261/A OR2X1_LOC_54/Y -0.04fF
C3563 AND2X1_LOC_307/Y AND2X1_LOC_308/a_8_24# 0.01fF
C3564 OR2X1_LOC_22/Y AND2X1_LOC_729/B 0.08fF
C3565 AND2X1_LOC_196/a_8_24# AND2X1_LOC_196/Y 0.01fF
C3566 OR2X1_LOC_144/a_8_216# OR2X1_LOC_12/Y 0.06fF
C3567 OR2X1_LOC_793/a_8_216# OR2X1_LOC_801/B 0.04fF
C3568 OR2X1_LOC_47/Y OR2X1_LOC_588/Y 0.02fF
C3569 OR2X1_LOC_32/B AND2X1_LOC_202/a_8_24# 0.03fF
C3570 OR2X1_LOC_99/a_8_216# D_INPUT_1 0.06fF
C3571 AND2X1_LOC_42/B AND2X1_LOC_47/Y 1.43fF
C3572 OR2X1_LOC_62/B OR2X1_LOC_415/A 0.01fF
C3573 AND2X1_LOC_851/B AND2X1_LOC_717/B 0.07fF
C3574 AND2X1_LOC_22/Y OR2X1_LOC_392/B 0.17fF
C3575 OR2X1_LOC_406/Y AND2X1_LOC_734/a_8_24# 0.01fF
C3576 AND2X1_LOC_539/Y AND2X1_LOC_802/Y 0.10fF
C3577 OR2X1_LOC_440/B OR2X1_LOC_180/B 0.01fF
C3578 OR2X1_LOC_696/A AND2X1_LOC_566/B 0.03fF
C3579 AND2X1_LOC_22/Y AND2X1_LOC_263/a_8_24# 0.05fF
C3580 OR2X1_LOC_625/Y AND2X1_LOC_790/a_8_24# 0.06fF
C3581 OR2X1_LOC_139/A OR2X1_LOC_576/A 0.01fF
C3582 OR2X1_LOC_476/B OR2X1_LOC_655/B 0.03fF
C3583 AND2X1_LOC_48/A OR2X1_LOC_814/A 0.09fF
C3584 AND2X1_LOC_860/a_8_24# OR2X1_LOC_13/B 0.01fF
C3585 AND2X1_LOC_43/B OR2X1_LOC_197/a_8_216# 0.03fF
C3586 AND2X1_LOC_7/B AND2X1_LOC_255/a_8_24# 0.01fF
C3587 OR2X1_LOC_161/A OR2X1_LOC_259/B 0.02fF
C3588 AND2X1_LOC_633/Y INPUT_1 0.02fF
C3589 OR2X1_LOC_215/Y OR2X1_LOC_228/Y 0.01fF
C3590 AND2X1_LOC_848/A OR2X1_LOC_44/Y 0.09fF
C3591 OR2X1_LOC_155/A OR2X1_LOC_194/a_8_216# 0.04fF
C3592 OR2X1_LOC_161/A OR2X1_LOC_68/B 0.04fF
C3593 OR2X1_LOC_18/Y OR2X1_LOC_384/a_8_216# 0.14fF
C3594 AND2X1_LOC_681/a_8_24# AND2X1_LOC_51/Y 0.01fF
C3595 AND2X1_LOC_703/Y AND2X1_LOC_714/a_8_24# 0.09fF
C3596 INPUT_1 D_INPUT_0 1.88fF
C3597 OR2X1_LOC_31/Y AND2X1_LOC_687/B 0.79fF
C3598 OR2X1_LOC_91/Y AND2X1_LOC_657/A 0.07fF
C3599 OR2X1_LOC_36/Y OR2X1_LOC_88/a_8_216# 0.02fF
C3600 OR2X1_LOC_78/A OR2X1_LOC_388/a_8_216# 0.01fF
C3601 AND2X1_LOC_191/Y OR2X1_LOC_747/a_36_216# 0.02fF
C3602 OR2X1_LOC_26/Y AND2X1_LOC_222/Y 0.06fF
C3603 OR2X1_LOC_36/Y OR2X1_LOC_172/a_8_216# -0.00fF
C3604 OR2X1_LOC_329/a_8_216# OR2X1_LOC_428/A 0.04fF
C3605 OR2X1_LOC_44/Y OR2X1_LOC_588/a_8_216# 0.19fF
C3606 OR2X1_LOC_160/A OR2X1_LOC_705/a_8_216# 0.04fF
C3607 AND2X1_LOC_171/a_36_24# OR2X1_LOC_339/Y 0.00fF
C3608 OR2X1_LOC_315/a_8_216# AND2X1_LOC_786/Y 0.04fF
C3609 AND2X1_LOC_59/Y AND2X1_LOC_406/a_8_24# 0.01fF
C3610 OR2X1_LOC_66/A OR2X1_LOC_415/Y 0.05fF
C3611 OR2X1_LOC_417/A OR2X1_LOC_226/a_36_216# 0.00fF
C3612 AND2X1_LOC_578/A OR2X1_LOC_419/Y 0.10fF
C3613 AND2X1_LOC_340/Y OR2X1_LOC_589/A 0.03fF
C3614 OR2X1_LOC_479/Y OR2X1_LOC_551/B 0.03fF
C3615 AND2X1_LOC_42/B OR2X1_LOC_598/A 0.14fF
C3616 OR2X1_LOC_36/Y OR2X1_LOC_378/A 0.07fF
C3617 OR2X1_LOC_553/A OR2X1_LOC_367/B 0.10fF
C3618 AND2X1_LOC_448/a_8_24# OR2X1_LOC_428/A 0.01fF
C3619 OR2X1_LOC_833/B OR2X1_LOC_777/B 0.07fF
C3620 OR2X1_LOC_89/A AND2X1_LOC_222/Y 0.03fF
C3621 AND2X1_LOC_351/Y OR2X1_LOC_289/Y 0.21fF
C3622 OR2X1_LOC_492/a_8_216# OR2X1_LOC_492/Y 0.01fF
C3623 OR2X1_LOC_190/A OR2X1_LOC_563/A 0.07fF
C3624 OR2X1_LOC_131/Y AND2X1_LOC_656/a_8_24# 0.24fF
C3625 OR2X1_LOC_70/Y OR2X1_LOC_331/a_8_216# 0.01fF
C3626 OR2X1_LOC_604/A AND2X1_LOC_786/Y 0.10fF
C3627 AND2X1_LOC_721/Y OR2X1_LOC_496/a_36_216# 0.00fF
C3628 OR2X1_LOC_121/Y AND2X1_LOC_625/a_8_24# 0.04fF
C3629 OR2X1_LOC_696/A AND2X1_LOC_391/a_8_24# 0.18fF
C3630 AND2X1_LOC_181/Y OR2X1_LOC_322/Y 0.03fF
C3631 OR2X1_LOC_45/B AND2X1_LOC_657/Y 0.01fF
C3632 AND2X1_LOC_534/a_8_24# AND2X1_LOC_110/Y 0.01fF
C3633 AND2X1_LOC_70/Y OR2X1_LOC_355/A 0.01fF
C3634 AND2X1_LOC_364/Y OR2X1_LOC_321/a_8_216# 0.03fF
C3635 OR2X1_LOC_244/B OR2X1_LOC_392/B 0.03fF
C3636 AND2X1_LOC_454/a_8_24# OR2X1_LOC_12/Y 0.03fF
C3637 AND2X1_LOC_858/B OR2X1_LOC_816/A 0.07fF
C3638 OR2X1_LOC_51/Y OR2X1_LOC_16/A 0.61fF
C3639 OR2X1_LOC_179/Y AND2X1_LOC_465/A 0.06fF
C3640 OR2X1_LOC_461/Y OR2X1_LOC_68/B 0.01fF
C3641 OR2X1_LOC_139/A AND2X1_LOC_41/A 0.29fF
C3642 AND2X1_LOC_51/Y OR2X1_LOC_68/B 3.59fF
C3643 OR2X1_LOC_634/A AND2X1_LOC_44/Y 0.09fF
C3644 OR2X1_LOC_696/A OR2X1_LOC_127/a_8_216# 0.01fF
C3645 AND2X1_LOC_363/B OR2X1_LOC_494/A 0.01fF
C3646 OR2X1_LOC_124/a_8_216# OR2X1_LOC_641/A 0.06fF
C3647 OR2X1_LOC_244/a_8_216# OR2X1_LOC_576/A 0.01fF
C3648 OR2X1_LOC_508/A OR2X1_LOC_139/A 0.10fF
C3649 OR2X1_LOC_363/B OR2X1_LOC_362/A 0.38fF
C3650 OR2X1_LOC_100/Y AND2X1_LOC_22/Y 1.97fF
C3651 OR2X1_LOC_58/Y OR2X1_LOC_600/A 0.03fF
C3652 OR2X1_LOC_8/Y INPUT_2 1.74fF
C3653 AND2X1_LOC_48/A OR2X1_LOC_341/a_8_216# 0.01fF
C3654 AND2X1_LOC_64/Y OR2X1_LOC_402/Y 0.09fF
C3655 AND2X1_LOC_727/Y AND2X1_LOC_550/A 0.01fF
C3656 AND2X1_LOC_574/A AND2X1_LOC_657/A 0.16fF
C3657 AND2X1_LOC_212/A OR2X1_LOC_91/A 0.04fF
C3658 AND2X1_LOC_22/Y AND2X1_LOC_58/a_36_24# 0.01fF
C3659 OR2X1_LOC_633/a_8_216# OR2X1_LOC_549/A 0.03fF
C3660 AND2X1_LOC_227/Y AND2X1_LOC_216/A 0.02fF
C3661 VDD AND2X1_LOC_285/Y 0.19fF
C3662 OR2X1_LOC_711/A AND2X1_LOC_36/Y 0.27fF
C3663 OR2X1_LOC_623/B OR2X1_LOC_161/B 0.03fF
C3664 VDD OR2X1_LOC_787/B 0.16fF
C3665 OR2X1_LOC_124/B AND2X1_LOC_70/Y 0.05fF
C3666 OR2X1_LOC_478/a_8_216# OR2X1_LOC_161/B 0.01fF
C3667 OR2X1_LOC_220/B AND2X1_LOC_7/B 0.02fF
C3668 AND2X1_LOC_329/a_8_24# OR2X1_LOC_703/Y 0.17fF
C3669 OR2X1_LOC_319/B OR2X1_LOC_535/A 0.01fF
C3670 OR2X1_LOC_158/A AND2X1_LOC_850/A 0.03fF
C3671 VDD AND2X1_LOC_92/Y 1.85fF
C3672 OR2X1_LOC_427/A AND2X1_LOC_464/A 0.03fF
C3673 OR2X1_LOC_756/B OR2X1_LOC_362/A 0.04fF
C3674 OR2X1_LOC_794/A OR2X1_LOC_161/B 0.00fF
C3675 OR2X1_LOC_427/A AND2X1_LOC_213/B 0.00fF
C3676 OR2X1_LOC_48/B AND2X1_LOC_771/a_8_24# 0.02fF
C3677 OR2X1_LOC_524/Y OR2X1_LOC_745/a_8_216# 0.09fF
C3678 OR2X1_LOC_185/A OR2X1_LOC_266/A 0.01fF
C3679 OR2X1_LOC_223/A OR2X1_LOC_318/B 0.01fF
C3680 AND2X1_LOC_64/Y OR2X1_LOC_642/a_8_216# 0.05fF
C3681 AND2X1_LOC_573/A OR2X1_LOC_816/A 0.03fF
C3682 OR2X1_LOC_269/B OR2X1_LOC_170/a_8_216# 0.06fF
C3683 AND2X1_LOC_40/Y OR2X1_LOC_151/A 0.32fF
C3684 OR2X1_LOC_632/Y OR2X1_LOC_66/A 0.06fF
C3685 OR2X1_LOC_6/B OR2X1_LOC_663/A 0.07fF
C3686 OR2X1_LOC_175/Y OR2X1_LOC_130/A 0.03fF
C3687 OR2X1_LOC_18/Y AND2X1_LOC_771/a_8_24# 0.02fF
C3688 AND2X1_LOC_707/a_8_24# OR2X1_LOC_91/A 0.03fF
C3689 OR2X1_LOC_833/B OR2X1_LOC_344/A 0.02fF
C3690 AND2X1_LOC_231/Y AND2X1_LOC_228/Y 0.07fF
C3691 OR2X1_LOC_178/Y OR2X1_LOC_329/B 0.00fF
C3692 D_INPUT_3 AND2X1_LOC_657/A 0.02fF
C3693 OR2X1_LOC_842/a_8_216# OR2X1_LOC_190/A 0.05fF
C3694 AND2X1_LOC_706/Y OR2X1_LOC_619/Y 0.01fF
C3695 AND2X1_LOC_21/Y AND2X1_LOC_762/a_36_24# 0.00fF
C3696 OR2X1_LOC_36/Y AND2X1_LOC_202/Y 0.00fF
C3697 AND2X1_LOC_82/Y OR2X1_LOC_402/Y 0.01fF
C3698 OR2X1_LOC_813/Y AND2X1_LOC_216/A 0.01fF
C3699 INPUT_0 OR2X1_LOC_78/A 0.03fF
C3700 OR2X1_LOC_691/Y OR2X1_LOC_130/A 0.02fF
C3701 AND2X1_LOC_449/Y OR2X1_LOC_12/Y 0.02fF
C3702 OR2X1_LOC_62/B OR2X1_LOC_141/a_8_216# 0.01fF
C3703 OR2X1_LOC_377/A OR2X1_LOC_856/A 0.02fF
C3704 VDD OR2X1_LOC_290/Y 0.15fF
C3705 AND2X1_LOC_365/A AND2X1_LOC_810/B 0.07fF
C3706 AND2X1_LOC_464/a_8_24# AND2X1_LOC_464/A -0.00fF
C3707 AND2X1_LOC_40/Y AND2X1_LOC_41/a_36_24# 0.01fF
C3708 AND2X1_LOC_729/Y OR2X1_LOC_167/a_36_216# 0.01fF
C3709 AND2X1_LOC_861/B AND2X1_LOC_865/A 0.01fF
C3710 AND2X1_LOC_786/a_8_24# OR2X1_LOC_262/Y 0.11fF
C3711 OR2X1_LOC_254/B OR2X1_LOC_344/A 0.01fF
C3712 OR2X1_LOC_232/Y OR2X1_LOC_234/Y 0.09fF
C3713 OR2X1_LOC_669/Y AND2X1_LOC_287/B 0.03fF
C3714 OR2X1_LOC_47/Y OR2X1_LOC_152/a_8_216# 0.05fF
C3715 OR2X1_LOC_97/A OR2X1_LOC_449/B 0.00fF
C3716 OR2X1_LOC_624/Y OR2X1_LOC_658/a_36_216# 0.03fF
C3717 AND2X1_LOC_509/Y AND2X1_LOC_508/A 0.00fF
C3718 AND2X1_LOC_804/a_8_24# AND2X1_LOC_222/Y 0.01fF
C3719 OR2X1_LOC_753/A OR2X1_LOC_753/a_8_216# 0.12fF
C3720 AND2X1_LOC_486/Y OR2X1_LOC_56/A 0.03fF
C3721 AND2X1_LOC_12/Y AND2X1_LOC_625/a_8_24# 0.02fF
C3722 OR2X1_LOC_43/A AND2X1_LOC_810/B 0.15fF
C3723 OR2X1_LOC_308/a_8_216# OR2X1_LOC_834/A 0.00fF
C3724 AND2X1_LOC_729/Y OR2X1_LOC_40/Y 0.03fF
C3725 AND2X1_LOC_736/Y AND2X1_LOC_675/Y 0.00fF
C3726 AND2X1_LOC_168/Y OR2X1_LOC_51/Y 0.01fF
C3727 AND2X1_LOC_741/Y AND2X1_LOC_220/Y 0.11fF
C3728 AND2X1_LOC_722/Y AND2X1_LOC_733/a_8_24# 0.18fF
C3729 AND2X1_LOC_776/a_8_24# OR2X1_LOC_18/Y 0.01fF
C3730 OR2X1_LOC_591/Y OR2X1_LOC_44/Y 0.04fF
C3731 VDD AND2X1_LOC_166/a_8_24# -0.00fF
C3732 OR2X1_LOC_864/A AND2X1_LOC_65/A 0.03fF
C3733 OR2X1_LOC_571/B OR2X1_LOC_244/Y 0.00fF
C3734 AND2X1_LOC_765/a_8_24# OR2X1_LOC_557/A 0.19fF
C3735 OR2X1_LOC_108/Y OR2X1_LOC_680/A 0.05fF
C3736 OR2X1_LOC_405/A OR2X1_LOC_858/A 0.02fF
C3737 OR2X1_LOC_7/A OR2X1_LOC_323/Y 0.08fF
C3738 OR2X1_LOC_185/Y OR2X1_LOC_6/B 0.10fF
C3739 OR2X1_LOC_170/Y OR2X1_LOC_568/a_8_216# 0.40fF
C3740 INPUT_0 AND2X1_LOC_520/Y 0.16fF
C3741 OR2X1_LOC_154/A AND2X1_LOC_18/Y 3.07fF
C3742 OR2X1_LOC_820/B OR2X1_LOC_382/a_8_216# 0.01fF
C3743 OR2X1_LOC_589/A OR2X1_LOC_585/A 0.03fF
C3744 OR2X1_LOC_91/Y VDD 0.50fF
C3745 OR2X1_LOC_235/B OR2X1_LOC_668/a_36_216# 0.00fF
C3746 AND2X1_LOC_402/a_8_24# AND2X1_LOC_404/A 0.00fF
C3747 OR2X1_LOC_270/Y D_GATE_366 0.74fF
C3748 AND2X1_LOC_329/a_8_24# OR2X1_LOC_596/A 0.06fF
C3749 OR2X1_LOC_633/B AND2X1_LOC_65/A 0.03fF
C3750 AND2X1_LOC_748/a_8_24# OR2X1_LOC_78/B 0.04fF
C3751 AND2X1_LOC_784/A OR2X1_LOC_40/Y 0.10fF
C3752 AND2X1_LOC_571/B OR2X1_LOC_71/Y 0.01fF
C3753 AND2X1_LOC_729/a_8_24# OR2X1_LOC_485/A 0.02fF
C3754 OR2X1_LOC_570/Y D_GATE_366 0.00fF
C3755 OR2X1_LOC_822/a_8_216# OR2X1_LOC_753/A 0.01fF
C3756 OR2X1_LOC_743/a_36_216# OR2X1_LOC_39/A 0.00fF
C3757 AND2X1_LOC_521/a_8_24# AND2X1_LOC_42/B 0.03fF
C3758 OR2X1_LOC_464/A OR2X1_LOC_733/a_8_216# 0.01fF
C3759 OR2X1_LOC_267/A AND2X1_LOC_18/Y 0.13fF
C3760 AND2X1_LOC_191/Y AND2X1_LOC_475/Y 0.03fF
C3761 OR2X1_LOC_305/Y VDD 0.16fF
C3762 OR2X1_LOC_168/a_36_216# OR2X1_LOC_756/B 0.00fF
C3763 OR2X1_LOC_177/Y AND2X1_LOC_578/A 0.03fF
C3764 AND2X1_LOC_738/B AND2X1_LOC_834/a_8_24# 0.04fF
C3765 OR2X1_LOC_97/A OR2X1_LOC_121/B 0.21fF
C3766 OR2X1_LOC_160/B AND2X1_LOC_159/a_8_24# 0.03fF
C3767 OR2X1_LOC_580/A OR2X1_LOC_366/a_8_216# 0.03fF
C3768 AND2X1_LOC_711/Y AND2X1_LOC_220/a_8_24# 0.05fF
C3769 VDD OR2X1_LOC_551/a_8_216# 0.00fF
C3770 OR2X1_LOC_144/Y OR2X1_LOC_427/A 0.03fF
C3771 OR2X1_LOC_160/B OR2X1_LOC_810/A 0.10fF
C3772 AND2X1_LOC_122/a_8_24# OR2X1_LOC_549/A 0.01fF
C3773 AND2X1_LOC_555/Y OR2X1_LOC_225/a_36_216# 0.00fF
C3774 OR2X1_LOC_734/a_8_216# OR2X1_LOC_737/A 0.03fF
C3775 AND2X1_LOC_344/a_8_24# OR2X1_LOC_625/Y 0.02fF
C3776 OR2X1_LOC_602/Y OR2X1_LOC_778/Y 0.23fF
C3777 AND2X1_LOC_721/Y AND2X1_LOC_471/a_8_24# 0.01fF
C3778 OR2X1_LOC_665/Y OR2X1_LOC_600/A 0.09fF
C3779 OR2X1_LOC_70/Y AND2X1_LOC_475/Y 0.18fF
C3780 OR2X1_LOC_251/Y AND2X1_LOC_285/Y 0.02fF
C3781 OR2X1_LOC_467/B OR2X1_LOC_470/B 0.28fF
C3782 OR2X1_LOC_151/A OR2X1_LOC_475/Y 0.15fF
C3783 AND2X1_LOC_486/Y AND2X1_LOC_850/Y 0.10fF
C3784 OR2X1_LOC_189/Y VDD 0.35fF
C3785 OR2X1_LOC_40/Y OR2X1_LOC_3/a_8_216# 0.40fF
C3786 VDD OR2X1_LOC_563/B 0.21fF
C3787 INPUT_5 AND2X1_LOC_43/B 0.02fF
C3788 OR2X1_LOC_485/A OR2X1_LOC_600/A 0.25fF
C3789 OR2X1_LOC_290/a_36_216# OR2X1_LOC_316/Y 0.00fF
C3790 OR2X1_LOC_822/Y AND2X1_LOC_240/Y 0.00fF
C3791 OR2X1_LOC_178/a_36_216# OR2X1_LOC_529/Y 0.00fF
C3792 OR2X1_LOC_274/Y OR2X1_LOC_375/A 0.01fF
C3793 VDD OR2X1_LOC_757/Y 0.00fF
C3794 OR2X1_LOC_158/A AND2X1_LOC_523/Y 0.10fF
C3795 OR2X1_LOC_279/a_8_216# AND2X1_LOC_860/A 0.01fF
C3796 OR2X1_LOC_279/Y AND2X1_LOC_243/Y 0.29fF
C3797 OR2X1_LOC_604/A AND2X1_LOC_578/A 2.96fF
C3798 VDD OR2X1_LOC_152/Y 0.39fF
C3799 AND2X1_LOC_794/B OR2X1_LOC_417/Y 0.02fF
C3800 OR2X1_LOC_759/A OR2X1_LOC_3/Y 0.02fF
C3801 OR2X1_LOC_254/B OR2X1_LOC_254/A 0.09fF
C3802 OR2X1_LOC_334/B AND2X1_LOC_56/B 0.02fF
C3803 AND2X1_LOC_22/Y OR2X1_LOC_532/B 0.11fF
C3804 OR2X1_LOC_46/A OR2X1_LOC_9/a_8_216# 0.01fF
C3805 AND2X1_LOC_228/Y AND2X1_LOC_654/B 0.00fF
C3806 AND2X1_LOC_341/a_8_24# D_INPUT_0 0.02fF
C3807 OR2X1_LOC_621/A AND2X1_LOC_670/a_36_24# 0.01fF
C3808 OR2X1_LOC_624/A OR2X1_LOC_668/a_8_216# 0.15fF
C3809 OR2X1_LOC_814/A OR2X1_LOC_489/A 0.01fF
C3810 AND2X1_LOC_621/Y AND2X1_LOC_804/Y 0.03fF
C3811 VDD AND2X1_LOC_183/a_8_24# -0.00fF
C3812 OR2X1_LOC_467/A OR2X1_LOC_453/Y 0.01fF
C3813 INPUT_0 OR2X1_LOC_155/A 0.02fF
C3814 OR2X1_LOC_152/Y AND2X1_LOC_738/a_8_24# 0.17fF
C3815 AND2X1_LOC_367/A OR2X1_LOC_26/Y 0.05fF
C3816 OR2X1_LOC_40/Y AND2X1_LOC_632/a_36_24# 0.01fF
C3817 AND2X1_LOC_736/Y OR2X1_LOC_189/A 0.04fF
C3818 OR2X1_LOC_660/a_8_216# OR2X1_LOC_520/Y 0.04fF
C3819 VDD OR2X1_LOC_527/Y 0.04fF
C3820 AND2X1_LOC_181/a_8_24# OR2X1_LOC_529/Y 0.01fF
C3821 AND2X1_LOC_710/Y AND2X1_LOC_347/a_8_24# 0.05fF
C3822 OR2X1_LOC_544/A OR2X1_LOC_161/B 0.04fF
C3823 OR2X1_LOC_482/Y OR2X1_LOC_628/Y 0.02fF
C3824 OR2X1_LOC_109/Y OR2X1_LOC_39/A 0.05fF
C3825 OR2X1_LOC_135/Y OR2X1_LOC_417/A 0.01fF
C3826 AND2X1_LOC_367/A OR2X1_LOC_89/A 0.17fF
C3827 VDD OR2X1_LOC_417/Y 0.46fF
C3828 VDD OR2X1_LOC_291/Y 0.38fF
C3829 AND2X1_LOC_807/Y AND2X1_LOC_573/A 0.03fF
C3830 OR2X1_LOC_185/Y OR2X1_LOC_523/Y 0.43fF
C3831 OR2X1_LOC_3/Y OR2X1_LOC_697/a_8_216# -0.00fF
C3832 AND2X1_LOC_363/B AND2X1_LOC_363/A 0.10fF
C3833 AND2X1_LOC_130/a_8_24# D_INPUT_0 0.03fF
C3834 OR2X1_LOC_40/Y AND2X1_LOC_639/A 0.00fF
C3835 OR2X1_LOC_31/Y OR2X1_LOC_322/a_8_216# 0.01fF
C3836 AND2X1_LOC_654/B OR2X1_LOC_585/A 0.03fF
C3837 VDD OR2X1_LOC_311/Y 0.11fF
C3838 OR2X1_LOC_814/A OR2X1_LOC_772/A 0.02fF
C3839 OR2X1_LOC_694/Y AND2X1_LOC_687/B 0.01fF
C3840 AND2X1_LOC_339/B OR2X1_LOC_75/a_8_216# 0.01fF
C3841 AND2X1_LOC_715/A AND2X1_LOC_115/a_8_24# 0.00fF
C3842 OR2X1_LOC_91/Y OR2X1_LOC_315/Y 0.27fF
C3843 OR2X1_LOC_3/Y OR2X1_LOC_698/Y 0.01fF
C3844 AND2X1_LOC_794/A AND2X1_LOC_784/A -0.01fF
C3845 VDD AND2X1_LOC_574/A 0.01fF
C3846 OR2X1_LOC_621/A OR2X1_LOC_532/B 0.21fF
C3847 OR2X1_LOC_624/A OR2X1_LOC_87/A 0.10fF
C3848 VDD AND2X1_LOC_538/Y 0.23fF
C3849 AND2X1_LOC_387/B OR2X1_LOC_502/A 0.01fF
C3850 OR2X1_LOC_3/Y D_INPUT_5 0.00fF
C3851 OR2X1_LOC_456/Y OR2X1_LOC_553/A 0.04fF
C3852 OR2X1_LOC_154/A OR2X1_LOC_500/A 0.06fF
C3853 OR2X1_LOC_448/Y OR2X1_LOC_779/a_8_216# 0.43fF
C3854 OR2X1_LOC_476/a_36_216# AND2X1_LOC_92/Y -0.01fF
C3855 INPUT_0 AND2X1_LOC_856/B 0.01fF
C3856 AND2X1_LOC_398/a_8_24# OR2X1_LOC_585/A 0.01fF
C3857 OR2X1_LOC_316/Y OR2X1_LOC_6/A 0.00fF
C3858 OR2X1_LOC_693/Y AND2X1_LOC_648/B 0.01fF
C3859 AND2X1_LOC_12/Y OR2X1_LOC_644/B 0.03fF
C3860 OR2X1_LOC_715/B OR2X1_LOC_436/Y 0.04fF
C3861 INPUT_0 AND2X1_LOC_863/A 0.03fF
C3862 OR2X1_LOC_51/Y AND2X1_LOC_687/Y -0.01fF
C3863 OR2X1_LOC_860/Y OR2X1_LOC_392/a_8_216# 0.01fF
C3864 AND2X1_LOC_474/A AND2X1_LOC_849/A 0.02fF
C3865 INPUT_4 AND2X1_LOC_30/a_8_24# 0.10fF
C3866 OR2X1_LOC_175/Y OR2X1_LOC_365/B 0.00fF
C3867 OR2X1_LOC_91/A AND2X1_LOC_727/A 0.01fF
C3868 OR2X1_LOC_269/Y OR2X1_LOC_549/A 0.01fF
C3869 AND2X1_LOC_454/Y OR2X1_LOC_52/B 0.08fF
C3870 OR2X1_LOC_103/Y AND2X1_LOC_523/Y 0.16fF
C3871 AND2X1_LOC_354/B OR2X1_LOC_6/A 0.17fF
C3872 OR2X1_LOC_485/A OR2X1_LOC_619/Y 0.03fF
C3873 INPUT_0 AND2X1_LOC_825/a_36_24# 0.01fF
C3874 AND2X1_LOC_191/Y OR2X1_LOC_616/a_8_216# 0.03fF
C3875 AND2X1_LOC_719/Y OR2X1_LOC_47/Y 0.03fF
C3876 AND2X1_LOC_732/a_8_24# OR2X1_LOC_31/Y 0.10fF
C3877 AND2X1_LOC_729/Y OR2X1_LOC_7/A 0.07fF
C3878 OR2X1_LOC_624/A OR2X1_LOC_216/a_8_216# 0.14fF
C3879 OR2X1_LOC_121/B OR2X1_LOC_475/B 0.01fF
C3880 VDD D_INPUT_3 1.12fF
C3881 OR2X1_LOC_74/A AND2X1_LOC_274/a_36_24# 0.01fF
C3882 OR2X1_LOC_749/Y AND2X1_LOC_750/a_8_24# 0.01fF
C3883 AND2X1_LOC_554/B AND2X1_LOC_123/Y 0.04fF
C3884 AND2X1_LOC_811/Y AND2X1_LOC_657/Y 0.34fF
C3885 AND2X1_LOC_106/a_8_24# OR2X1_LOC_244/Y 0.00fF
C3886 OR2X1_LOC_599/A OR2X1_LOC_52/B 0.07fF
C3887 OR2X1_LOC_158/B OR2X1_LOC_619/Y 0.01fF
C3888 AND2X1_LOC_30/a_8_24# AND2X1_LOC_51/A 0.00fF
C3889 OR2X1_LOC_103/a_8_216# AND2X1_LOC_523/Y 0.03fF
C3890 OR2X1_LOC_779/B OR2X1_LOC_779/A 0.37fF
C3891 OR2X1_LOC_590/Y OR2X1_LOC_593/B 0.01fF
C3892 OR2X1_LOC_244/B OR2X1_LOC_532/B 0.01fF
C3893 OR2X1_LOC_709/A AND2X1_LOC_699/a_8_24# 0.00fF
C3894 AND2X1_LOC_658/A AND2X1_LOC_796/Y 0.03fF
C3895 AND2X1_LOC_42/B AND2X1_LOC_129/a_8_24# 0.00fF
C3896 OR2X1_LOC_43/A OR2X1_LOC_585/A 0.10fF
C3897 AND2X1_LOC_842/a_8_24# OR2X1_LOC_71/Y 0.08fF
C3898 AND2X1_LOC_858/B OR2X1_LOC_95/Y 0.09fF
C3899 AND2X1_LOC_811/Y AND2X1_LOC_469/B 0.02fF
C3900 OR2X1_LOC_517/A D_INPUT_0 0.22fF
C3901 OR2X1_LOC_91/A OR2X1_LOC_95/Y 0.08fF
C3902 OR2X1_LOC_32/a_8_216# OR2X1_LOC_753/A 0.30fF
C3903 OR2X1_LOC_831/a_8_216# OR2X1_LOC_479/Y 0.02fF
C3904 OR2X1_LOC_488/Y AND2X1_LOC_573/A 0.02fF
C3905 AND2X1_LOC_673/a_8_24# OR2X1_LOC_26/Y 0.01fF
C3906 AND2X1_LOC_59/Y AND2X1_LOC_67/Y 0.05fF
C3907 AND2X1_LOC_784/A OR2X1_LOC_7/A 0.07fF
C3908 AND2X1_LOC_717/B OR2X1_LOC_372/Y 0.15fF
C3909 OR2X1_LOC_486/B OR2X1_LOC_738/A 0.01fF
C3910 AND2X1_LOC_141/A OR2X1_LOC_71/Y 0.00fF
C3911 OR2X1_LOC_629/Y OR2X1_LOC_62/B 0.01fF
C3912 OR2X1_LOC_709/A AND2X1_LOC_679/a_36_24# 0.00fF
C3913 OR2X1_LOC_663/A AND2X1_LOC_47/Y 0.57fF
C3914 OR2X1_LOC_70/Y AND2X1_LOC_266/Y 0.03fF
C3915 OR2X1_LOC_311/Y OR2X1_LOC_829/a_8_216# 0.01fF
C3916 OR2X1_LOC_48/Y OR2X1_LOC_36/Y 0.01fF
C3917 AND2X1_LOC_31/Y AND2X1_LOC_433/a_8_24# 0.01fF
C3918 OR2X1_LOC_351/B OR2X1_LOC_351/a_36_216# 0.02fF
C3919 OR2X1_LOC_46/A OR2X1_LOC_394/Y 0.08fF
C3920 OR2X1_LOC_160/A OR2X1_LOC_476/B 0.07fF
C3921 OR2X1_LOC_26/Y OR2X1_LOC_74/A 0.27fF
C3922 OR2X1_LOC_863/a_8_216# OR2X1_LOC_863/B 0.05fF
C3923 OR2X1_LOC_291/a_36_216# OR2X1_LOC_62/B 0.00fF
C3924 VDD AND2X1_LOC_483/Y -0.00fF
C3925 AND2X1_LOC_17/Y AND2X1_LOC_18/a_8_24# 0.06fF
C3926 OR2X1_LOC_854/a_36_216# OR2X1_LOC_532/B 0.00fF
C3927 OR2X1_LOC_160/A OR2X1_LOC_650/Y 0.07fF
C3928 AND2X1_LOC_456/Y OR2X1_LOC_89/A 0.02fF
C3929 OR2X1_LOC_277/a_8_216# OR2X1_LOC_85/A 0.08fF
C3930 OR2X1_LOC_490/Y OR2X1_LOC_89/A 0.00fF
C3931 OR2X1_LOC_74/A OR2X1_LOC_89/A 0.14fF
C3932 AND2X1_LOC_520/Y OR2X1_LOC_417/A 0.04fF
C3933 OR2X1_LOC_283/Y OR2X1_LOC_64/Y 0.05fF
C3934 OR2X1_LOC_479/Y OR2X1_LOC_787/Y 0.19fF
C3935 AND2X1_LOC_64/Y OR2X1_LOC_593/B 0.01fF
C3936 OR2X1_LOC_453/Y OR2X1_LOC_466/a_8_216# 0.39fF
C3937 OR2X1_LOC_60/a_8_216# OR2X1_LOC_585/A 0.02fF
C3938 OR2X1_LOC_604/A OR2X1_LOC_746/Y 0.16fF
C3939 OR2X1_LOC_745/a_8_216# OR2X1_LOC_746/Y 0.39fF
C3940 AND2X1_LOC_12/Y AND2X1_LOC_53/Y 0.09fF
C3941 OR2X1_LOC_59/Y AND2X1_LOC_205/a_36_24# 0.00fF
C3942 OR2X1_LOC_427/Y AND2X1_LOC_451/Y 0.01fF
C3943 AND2X1_LOC_587/a_8_24# D_INPUT_6 0.01fF
C3944 OR2X1_LOC_510/Y OR2X1_LOC_244/A 0.01fF
C3945 AND2X1_LOC_18/Y OR2X1_LOC_560/A 0.06fF
C3946 OR2X1_LOC_89/A OR2X1_LOC_261/A 0.79fF
C3947 OR2X1_LOC_95/Y AND2X1_LOC_573/A 0.11fF
C3948 OR2X1_LOC_417/A AND2X1_LOC_848/Y 0.06fF
C3949 AND2X1_LOC_571/A OR2X1_LOC_696/A 0.01fF
C3950 OR2X1_LOC_22/Y AND2X1_LOC_264/a_8_24# 0.03fF
C3951 AND2X1_LOC_588/B INPUT_6 -0.01fF
C3952 VDD OR2X1_LOC_561/B 0.03fF
C3953 OR2X1_LOC_447/Y OR2X1_LOC_87/A 0.07fF
C3954 AND2X1_LOC_339/B OR2X1_LOC_13/B 0.03fF
C3955 OR2X1_LOC_663/A OR2X1_LOC_598/A 0.07fF
C3956 AND2X1_LOC_171/a_8_24# AND2X1_LOC_48/A 0.03fF
C3957 OR2X1_LOC_364/A AND2X1_LOC_47/Y 0.21fF
C3958 OR2X1_LOC_185/Y AND2X1_LOC_47/Y 0.16fF
C3959 OR2X1_LOC_506/a_8_216# AND2X1_LOC_64/Y 0.06fF
C3960 AND2X1_LOC_12/Y OR2X1_LOC_223/A 0.03fF
C3961 OR2X1_LOC_283/Y OR2X1_LOC_417/A 0.07fF
C3962 OR2X1_LOC_611/Y OR2X1_LOC_612/B 0.06fF
C3963 AND2X1_LOC_387/B AND2X1_LOC_48/A 0.08fF
C3964 OR2X1_LOC_831/A OR2X1_LOC_716/a_8_216# 0.01fF
C3965 OR2X1_LOC_605/a_8_216# OR2X1_LOC_121/B 0.01fF
C3966 AND2X1_LOC_3/Y OR2X1_LOC_814/A 0.22fF
C3967 AND2X1_LOC_313/a_8_24# OR2X1_LOC_732/A 0.08fF
C3968 OR2X1_LOC_676/Y OR2X1_LOC_446/B 0.05fF
C3969 OR2X1_LOC_744/A OR2X1_LOC_80/A 0.23fF
C3970 OR2X1_LOC_416/a_8_216# OR2X1_LOC_6/A 0.08fF
C3971 AND2X1_LOC_137/a_8_24# AND2X1_LOC_361/A 0.02fF
C3972 OR2X1_LOC_62/B OR2X1_LOC_629/a_36_216# 0.00fF
C3973 AND2X1_LOC_543/Y AND2X1_LOC_564/B 0.02fF
C3974 OR2X1_LOC_502/A OR2X1_LOC_854/A 0.03fF
C3975 OR2X1_LOC_440/B OR2X1_LOC_788/B 0.10fF
C3976 OR2X1_LOC_64/Y AND2X1_LOC_863/A 0.17fF
C3977 OR2X1_LOC_277/a_36_216# OR2X1_LOC_278/A 0.01fF
C3978 AND2X1_LOC_640/Y AND2X1_LOC_640/a_36_24# 0.01fF
C3979 AND2X1_LOC_543/Y OR2X1_LOC_368/Y 0.78fF
C3980 OR2X1_LOC_834/A OR2X1_LOC_446/B 0.03fF
C3981 OR2X1_LOC_841/B OR2X1_LOC_223/A 0.01fF
C3982 OR2X1_LOC_251/Y D_INPUT_3 0.19fF
C3983 OR2X1_LOC_640/A OR2X1_LOC_68/B 0.01fF
C3984 OR2X1_LOC_280/Y AND2X1_LOC_227/Y 0.03fF
C3985 AND2X1_LOC_753/B AND2X1_LOC_31/Y 0.04fF
C3986 OR2X1_LOC_639/B AND2X1_LOC_428/a_8_24# 0.25fF
C3987 AND2X1_LOC_853/a_8_24# D_INPUT_0 0.01fF
C3988 AND2X1_LOC_489/Y AND2X1_LOC_866/A 0.03fF
C3989 OR2X1_LOC_245/a_8_216# OR2X1_LOC_246/A 0.01fF
C3990 OR2X1_LOC_728/B OR2X1_LOC_739/A 0.12fF
C3991 AND2X1_LOC_231/Y OR2X1_LOC_230/Y 0.79fF
C3992 OR2X1_LOC_267/Y AND2X1_LOC_44/Y 0.03fF
C3993 OR2X1_LOC_47/Y OR2X1_LOC_609/A 0.03fF
C3994 OR2X1_LOC_22/Y OR2X1_LOC_46/A 0.05fF
C3995 OR2X1_LOC_615/Y OR2X1_LOC_754/a_8_216# 0.41fF
C3996 OR2X1_LOC_405/A AND2X1_LOC_31/Y 0.57fF
C3997 OR2X1_LOC_78/B OR2X1_LOC_535/a_8_216# 0.01fF
C3998 OR2X1_LOC_185/Y OR2X1_LOC_598/A 0.10fF
C3999 AND2X1_LOC_572/a_8_24# OR2X1_LOC_595/A 0.03fF
C4000 OR2X1_LOC_755/A AND2X1_LOC_866/A 0.01fF
C4001 OR2X1_LOC_223/A OR2X1_LOC_804/B 0.09fF
C4002 OR2X1_LOC_551/a_8_216# OR2X1_LOC_551/A 0.39fF
C4003 AND2X1_LOC_341/a_8_24# AND2X1_LOC_350/B 0.04fF
C4004 OR2X1_LOC_362/A OR2X1_LOC_140/B 0.01fF
C4005 OR2X1_LOC_31/Y OR2X1_LOC_416/Y 0.03fF
C4006 OR2X1_LOC_174/A OR2X1_LOC_339/A 0.11fF
C4007 AND2X1_LOC_42/B D_INPUT_1 0.67fF
C4008 OR2X1_LOC_756/B OR2X1_LOC_771/B 0.14fF
C4009 OR2X1_LOC_66/A OR2X1_LOC_168/Y 1.10fF
C4010 OR2X1_LOC_59/Y OR2X1_LOC_183/Y 0.04fF
C4011 OR2X1_LOC_123/B OR2X1_LOC_786/Y 0.01fF
C4012 AND2X1_LOC_711/Y AND2X1_LOC_623/a_8_24# 0.07fF
C4013 OR2X1_LOC_36/Y AND2X1_LOC_779/Y 0.03fF
C4014 AND2X1_LOC_421/a_8_24# OR2X1_LOC_777/B 0.17fF
C4015 AND2X1_LOC_40/Y OR2X1_LOC_716/a_8_216# 0.03fF
C4016 OR2X1_LOC_22/Y AND2X1_LOC_227/Y 0.07fF
C4017 AND2X1_LOC_464/A OR2X1_LOC_322/a_8_216# 0.47fF
C4018 VDD OR2X1_LOC_171/Y 0.27fF
C4019 OR2X1_LOC_368/Y OR2X1_LOC_322/Y 0.01fF
C4020 AND2X1_LOC_841/B OR2X1_LOC_437/A 0.07fF
C4021 OR2X1_LOC_74/A AND2X1_LOC_804/a_8_24# 0.01fF
C4022 OR2X1_LOC_499/B AND2X1_LOC_36/Y 0.01fF
C4023 OR2X1_LOC_89/A AND2X1_LOC_647/Y 0.00fF
C4024 AND2X1_LOC_91/B OR2X1_LOC_602/Y 0.11fF
C4025 OR2X1_LOC_736/Y AND2X1_LOC_295/a_8_24# 0.01fF
C4026 OR2X1_LOC_175/Y OR2X1_LOC_468/A 0.07fF
C4027 OR2X1_LOC_132/a_36_216# OR2X1_LOC_134/Y 0.00fF
C4028 AND2X1_LOC_727/Y AND2X1_LOC_663/A 0.45fF
C4029 OR2X1_LOC_408/Y OR2X1_LOC_409/B 0.14fF
C4030 OR2X1_LOC_151/A OR2X1_LOC_356/A 0.02fF
C4031 OR2X1_LOC_673/Y OR2X1_LOC_71/A 0.01fF
C4032 OR2X1_LOC_454/a_8_216# OR2X1_LOC_783/A 0.39fF
C4033 AND2X1_LOC_95/Y OR2X1_LOC_174/Y 0.03fF
C4034 AND2X1_LOC_300/a_8_24# OR2X1_LOC_831/A 0.02fF
C4035 OR2X1_LOC_140/A OR2X1_LOC_161/B 0.01fF
C4036 OR2X1_LOC_89/A AND2X1_LOC_783/a_8_24# 0.01fF
C4037 OR2X1_LOC_7/A OR2X1_LOC_172/Y 0.00fF
C4038 OR2X1_LOC_279/a_8_216# AND2X1_LOC_562/Y 0.10fF
C4039 OR2X1_LOC_711/B OR2X1_LOC_711/a_8_216# 0.04fF
C4040 OR2X1_LOC_117/a_8_216# OR2X1_LOC_426/B 0.01fF
C4041 OR2X1_LOC_139/A OR2X1_LOC_648/A 0.07fF
C4042 OR2X1_LOC_78/A AND2X1_LOC_7/B 0.27fF
C4043 OR2X1_LOC_696/A OR2X1_LOC_92/Y 14.46fF
C4044 OR2X1_LOC_389/A OR2X1_LOC_389/a_8_216# 0.01fF
C4045 AND2X1_LOC_130/a_8_24# OR2X1_LOC_131/A 0.14fF
C4046 OR2X1_LOC_435/A AND2X1_LOC_18/Y 0.01fF
C4047 AND2X1_LOC_739/a_8_24# AND2X1_LOC_742/A 0.20fF
C4048 AND2X1_LOC_740/B AND2X1_LOC_740/a_8_24# 0.05fF
C4049 OR2X1_LOC_472/B OR2X1_LOC_598/A 0.01fF
C4050 OR2X1_LOC_22/Y OR2X1_LOC_41/Y 0.28fF
C4051 AND2X1_LOC_392/A AND2X1_LOC_566/B 0.07fF
C4052 AND2X1_LOC_778/Y AND2X1_LOC_784/a_8_24# 0.11fF
C4053 AND2X1_LOC_560/a_8_24# OR2X1_LOC_427/A 0.02fF
C4054 OR2X1_LOC_653/B AND2X1_LOC_70/Y 0.00fF
C4055 OR2X1_LOC_696/A AND2X1_LOC_801/a_36_24# 0.01fF
C4056 OR2X1_LOC_22/Y OR2X1_LOC_753/Y 0.02fF
C4057 AND2X1_LOC_705/Y OR2X1_LOC_59/Y 0.07fF
C4058 OR2X1_LOC_614/Y AND2X1_LOC_70/Y 0.01fF
C4059 OR2X1_LOC_49/A OR2X1_LOC_235/B 0.11fF
C4060 AND2X1_LOC_715/Y OR2X1_LOC_92/Y 1.05fF
C4061 AND2X1_LOC_191/B OR2X1_LOC_158/A 0.18fF
C4062 AND2X1_LOC_231/Y AND2X1_LOC_857/Y 0.01fF
C4063 OR2X1_LOC_647/a_8_216# OR2X1_LOC_68/B 0.01fF
C4064 OR2X1_LOC_8/Y OR2X1_LOC_40/Y 0.07fF
C4065 OR2X1_LOC_524/Y AND2X1_LOC_212/Y 0.10fF
C4066 AND2X1_LOC_60/a_8_24# AND2X1_LOC_58/a_8_24# 0.23fF
C4067 AND2X1_LOC_535/Y AND2X1_LOC_436/Y 1.13fF
C4068 OR2X1_LOC_186/Y AND2X1_LOC_312/a_36_24# 0.00fF
C4069 OR2X1_LOC_666/a_8_216# OR2X1_LOC_51/Y 0.01fF
C4070 OR2X1_LOC_92/a_8_216# AND2X1_LOC_647/Y 0.01fF
C4071 OR2X1_LOC_711/A OR2X1_LOC_469/B 0.04fF
C4072 AND2X1_LOC_715/Y AND2X1_LOC_801/a_36_24# 0.01fF
C4073 OR2X1_LOC_47/Y OR2X1_LOC_599/Y 0.02fF
C4074 OR2X1_LOC_276/a_36_216# OR2X1_LOC_66/Y 0.02fF
C4075 OR2X1_LOC_709/A OR2X1_LOC_808/B 0.10fF
C4076 OR2X1_LOC_602/Y OR2X1_LOC_645/a_8_216# 0.01fF
C4077 OR2X1_LOC_243/a_8_216# OR2X1_LOC_68/B 0.01fF
C4078 OR2X1_LOC_274/Y OR2X1_LOC_549/A 0.07fF
C4079 OR2X1_LOC_185/Y OR2X1_LOC_186/a_8_216# 0.19fF
C4080 OR2X1_LOC_589/A AND2X1_LOC_857/Y 0.03fF
C4081 VDD OR2X1_LOC_402/B 0.04fF
C4082 OR2X1_LOC_131/A OR2X1_LOC_517/A 0.10fF
C4083 AND2X1_LOC_47/Y AND2X1_LOC_432/a_8_24# 0.01fF
C4084 AND2X1_LOC_142/a_8_24# OR2X1_LOC_486/Y 0.25fF
C4085 OR2X1_LOC_18/Y AND2X1_LOC_785/Y 0.04fF
C4086 OR2X1_LOC_833/B OR2X1_LOC_161/B 0.00fF
C4087 OR2X1_LOC_484/Y AND2X1_LOC_436/Y 0.13fF
C4088 AND2X1_LOC_47/Y OR2X1_LOC_578/B 0.03fF
C4089 OR2X1_LOC_485/Y AND2X1_LOC_513/a_8_24# 0.17fF
C4090 OR2X1_LOC_186/Y OR2X1_LOC_739/A 0.04fF
C4091 OR2X1_LOC_520/Y AND2X1_LOC_44/Y 0.03fF
C4092 OR2X1_LOC_121/a_8_216# OR2X1_LOC_241/a_8_216# 0.47fF
C4093 OR2X1_LOC_254/B OR2X1_LOC_161/B 0.04fF
C4094 AND2X1_LOC_95/Y OR2X1_LOC_729/a_8_216# 0.01fF
C4095 OR2X1_LOC_175/Y OR2X1_LOC_449/B 0.07fF
C4096 OR2X1_LOC_176/a_8_216# AND2X1_LOC_784/A 0.03fF
C4097 OR2X1_LOC_680/A OR2X1_LOC_373/Y 0.07fF
C4098 OR2X1_LOC_382/Y OR2X1_LOC_56/A 0.01fF
C4099 OR2X1_LOC_779/Y AND2X1_LOC_31/Y 0.01fF
C4100 AND2X1_LOC_70/Y OR2X1_LOC_808/B 0.11fF
C4101 AND2X1_LOC_812/a_36_24# OR2X1_LOC_152/A 0.00fF
C4102 OR2X1_LOC_814/A OR2X1_LOC_576/a_8_216# 0.01fF
C4103 OR2X1_LOC_31/Y AND2X1_LOC_592/a_8_24# 0.01fF
C4104 OR2X1_LOC_186/Y OR2X1_LOC_798/a_8_216# -0.00fF
C4105 OR2X1_LOC_499/B OR2X1_LOC_630/Y 0.00fF
C4106 OR2X1_LOC_155/A AND2X1_LOC_7/B 0.14fF
C4107 OR2X1_LOC_51/Y OR2X1_LOC_426/A 0.02fF
C4108 OR2X1_LOC_151/A AND2X1_LOC_43/B 4.32fF
C4109 OR2X1_LOC_690/A AND2X1_LOC_214/a_8_24# 0.17fF
C4110 AND2X1_LOC_12/Y AND2X1_LOC_275/a_36_24# 0.00fF
C4111 AND2X1_LOC_863/a_36_24# OR2X1_LOC_56/A 0.00fF
C4112 AND2X1_LOC_759/a_8_24# OR2X1_LOC_792/Y 0.01fF
C4113 AND2X1_LOC_553/A OR2X1_LOC_59/Y 0.01fF
C4114 OR2X1_LOC_186/Y OR2X1_LOC_269/B 0.03fF
C4115 OR2X1_LOC_318/Y OR2X1_LOC_78/A 0.07fF
C4116 OR2X1_LOC_354/A AND2X1_LOC_167/a_8_24# 0.01fF
C4117 OR2X1_LOC_538/A OR2X1_LOC_502/A 0.03fF
C4118 OR2X1_LOC_45/B OR2X1_LOC_438/a_8_216# 0.06fF
C4119 OR2X1_LOC_449/B OR2X1_LOC_713/A 0.07fF
C4120 OR2X1_LOC_177/a_8_216# OR2X1_LOC_52/B 0.02fF
C4121 OR2X1_LOC_751/A OR2X1_LOC_749/Y 0.01fF
C4122 OR2X1_LOC_703/A OR2X1_LOC_808/B 0.03fF
C4123 AND2X1_LOC_40/Y OR2X1_LOC_174/A 0.01fF
C4124 AND2X1_LOC_593/Y AND2X1_LOC_447/Y 0.07fF
C4125 AND2X1_LOC_41/a_36_24# AND2X1_LOC_43/B 0.00fF
C4126 AND2X1_LOC_182/A OR2X1_LOC_91/a_8_216# 0.48fF
C4127 AND2X1_LOC_40/Y OR2X1_LOC_435/a_8_216# 0.01fF
C4128 AND2X1_LOC_857/Y AND2X1_LOC_654/B 0.34fF
C4129 D_INPUT_5 OR2X1_LOC_502/A 0.06fF
C4130 OR2X1_LOC_124/B OR2X1_LOC_217/Y 0.02fF
C4131 AND2X1_LOC_721/Y AND2X1_LOC_523/Y 0.37fF
C4132 OR2X1_LOC_656/Y OR2X1_LOC_660/a_8_216# 0.18fF
C4133 INPUT_4 OR2X1_LOC_51/Y 0.06fF
C4134 AND2X1_LOC_339/B AND2X1_LOC_339/a_36_24# 0.01fF
C4135 VDD OR2X1_LOC_457/a_8_216# 0.21fF
C4136 OR2X1_LOC_8/Y OR2X1_LOC_618/a_8_216# 0.01fF
C4137 AND2X1_LOC_59/Y OR2X1_LOC_520/a_8_216# 0.01fF
C4138 OR2X1_LOC_676/Y AND2X1_LOC_56/B 0.01fF
C4139 OR2X1_LOC_495/a_8_216# OR2X1_LOC_600/A 0.06fF
C4140 OR2X1_LOC_653/B OR2X1_LOC_653/a_8_216# 0.05fF
C4141 OR2X1_LOC_114/a_8_216# AND2X1_LOC_95/Y 0.01fF
C4142 OR2X1_LOC_805/A OR2X1_LOC_78/A 0.10fF
C4143 OR2X1_LOC_40/Y OR2X1_LOC_52/B 0.96fF
C4144 AND2X1_LOC_578/A AND2X1_LOC_212/Y 0.01fF
C4145 OR2X1_LOC_26/Y AND2X1_LOC_860/A 0.04fF
C4146 OR2X1_LOC_40/Y OR2X1_LOC_672/Y 0.00fF
C4147 OR2X1_LOC_600/A AND2X1_LOC_838/a_8_24# 0.01fF
C4148 VDD OR2X1_LOC_701/a_8_216# 0.21fF
C4149 AND2X1_LOC_526/a_8_24# OR2X1_LOC_161/A 0.01fF
C4150 VDD AND2X1_LOC_806/A 0.31fF
C4151 OR2X1_LOC_511/Y OR2X1_LOC_59/Y 0.03fF
C4152 AND2X1_LOC_99/A AND2X1_LOC_99/a_8_24# 0.05fF
C4153 OR2X1_LOC_756/B OR2X1_LOC_402/Y 0.21fF
C4154 VDD OR2X1_LOC_83/A 0.00fF
C4155 AND2X1_LOC_566/a_8_24# AND2X1_LOC_568/B 0.01fF
C4156 OR2X1_LOC_389/B VDD 0.00fF
C4157 OR2X1_LOC_168/a_8_216# OR2X1_LOC_840/A 0.33fF
C4158 OR2X1_LOC_11/Y OR2X1_LOC_26/a_8_216# 0.01fF
C4159 AND2X1_LOC_91/B OR2X1_LOC_602/B 0.04fF
C4160 OR2X1_LOC_527/a_8_216# OR2X1_LOC_485/A 0.06fF
C4161 AND2X1_LOC_602/a_8_24# AND2X1_LOC_447/Y 0.04fF
C4162 OR2X1_LOC_653/Y OR2X1_LOC_61/Y 0.01fF
C4163 OR2X1_LOC_39/Y OR2X1_LOC_39/A 0.06fF
C4164 AND2X1_LOC_833/a_8_24# AND2X1_LOC_840/A 0.01fF
C4165 OR2X1_LOC_495/a_36_216# OR2X1_LOC_56/A 0.02fF
C4166 OR2X1_LOC_107/a_8_216# OR2X1_LOC_44/Y 0.02fF
C4167 OR2X1_LOC_744/A OR2X1_LOC_6/A 0.33fF
C4168 OR2X1_LOC_89/A AND2X1_LOC_860/A 4.36fF
C4169 OR2X1_LOC_184/Y OR2X1_LOC_183/Y 0.14fF
C4170 OR2X1_LOC_458/B OR2X1_LOC_805/A 0.10fF
C4171 OR2X1_LOC_600/A OR2X1_LOC_827/Y 0.00fF
C4172 OR2X1_LOC_100/a_8_216# OR2X1_LOC_502/A 0.01fF
C4173 OR2X1_LOC_604/A OR2X1_LOC_418/a_8_216# 0.01fF
C4174 OR2X1_LOC_405/A OR2X1_LOC_473/a_36_216# 0.00fF
C4175 OR2X1_LOC_49/A OR2X1_LOC_293/a_36_216# 0.00fF
C4176 AND2X1_LOC_107/a_8_24# AND2X1_LOC_44/Y 0.01fF
C4177 AND2X1_LOC_364/A OR2X1_LOC_48/B 0.01fF
C4178 AND2X1_LOC_126/a_8_24# OR2X1_LOC_375/A 0.04fF
C4179 OR2X1_LOC_8/Y OR2X1_LOC_7/A 0.03fF
C4180 OR2X1_LOC_585/A OR2X1_LOC_585/Y 0.01fF
C4181 OR2X1_LOC_121/B OR2X1_LOC_713/A 0.07fF
C4182 AND2X1_LOC_12/Y OR2X1_LOC_502/A 0.16fF
C4183 AND2X1_LOC_693/a_36_24# OR2X1_LOC_375/A 0.00fF
C4184 OR2X1_LOC_651/B AND2X1_LOC_43/B 0.01fF
C4185 OR2X1_LOC_6/B AND2X1_LOC_496/a_36_24# 0.01fF
C4186 AND2X1_LOC_801/a_8_24# AND2X1_LOC_809/A 0.00fF
C4187 VDD AND2X1_LOC_276/Y 0.46fF
C4188 OR2X1_LOC_54/Y OR2X1_LOC_381/a_8_216# 0.03fF
C4189 OR2X1_LOC_668/a_8_216# OR2X1_LOC_161/A 0.01fF
C4190 OR2X1_LOC_40/Y OR2X1_LOC_755/A 0.93fF
C4191 OR2X1_LOC_91/Y AND2X1_LOC_486/Y 0.07fF
C4192 AND2X1_LOC_347/Y OR2X1_LOC_43/A 0.06fF
C4193 OR2X1_LOC_297/Y OR2X1_LOC_59/Y 0.01fF
C4194 AND2X1_LOC_712/B AND2X1_LOC_448/a_8_24# 0.02fF
C4195 OR2X1_LOC_501/B AND2X1_LOC_3/Y 0.03fF
C4196 OR2X1_LOC_625/Y OR2X1_LOC_252/Y 0.00fF
C4197 OR2X1_LOC_43/A AND2X1_LOC_857/Y 0.03fF
C4198 AND2X1_LOC_465/a_8_24# OR2X1_LOC_744/A 0.02fF
C4199 OR2X1_LOC_296/Y OR2X1_LOC_78/A 0.01fF
C4200 OR2X1_LOC_235/B AND2X1_LOC_85/a_8_24# 0.01fF
C4201 OR2X1_LOC_227/Y AND2X1_LOC_224/a_8_24# 0.23fF
C4202 OR2X1_LOC_862/A OR2X1_LOC_269/B 0.01fF
C4203 OR2X1_LOC_307/a_8_216# OR2X1_LOC_307/B 0.06fF
C4204 AND2X1_LOC_557/a_8_24# OR2X1_LOC_744/A 0.02fF
C4205 AND2X1_LOC_359/a_8_24# OR2X1_LOC_92/Y 0.01fF
C4206 AND2X1_LOC_12/Y AND2X1_LOC_230/a_8_24# 0.01fF
C4207 OR2X1_LOC_154/A OR2X1_LOC_560/a_8_216# 0.03fF
C4208 OR2X1_LOC_319/B OR2X1_LOC_155/A 0.19fF
C4209 AND2X1_LOC_578/A AND2X1_LOC_549/a_8_24# 0.01fF
C4210 AND2X1_LOC_377/a_8_24# AND2X1_LOC_472/B 0.07fF
C4211 AND2X1_LOC_301/a_8_24# OR2X1_LOC_416/Y 0.01fF
C4212 OR2X1_LOC_91/Y AND2X1_LOC_571/Y 0.08fF
C4213 AND2X1_LOC_364/Y OR2X1_LOC_321/Y 0.02fF
C4214 OR2X1_LOC_703/B OR2X1_LOC_161/A 0.03fF
C4215 OR2X1_LOC_520/B OR2X1_LOC_66/A 0.17fF
C4216 OR2X1_LOC_479/Y AND2X1_LOC_41/A 0.07fF
C4217 AND2X1_LOC_376/a_8_24# OR2X1_LOC_502/A 0.01fF
C4218 OR2X1_LOC_185/Y OR2X1_LOC_506/A 0.15fF
C4219 OR2X1_LOC_87/A OR2X1_LOC_161/A 0.28fF
C4220 AND2X1_LOC_359/a_36_24# OR2X1_LOC_427/A 0.01fF
C4221 OR2X1_LOC_154/A AND2X1_LOC_394/a_8_24# 0.20fF
C4222 OR2X1_LOC_196/B OR2X1_LOC_702/a_8_216# 0.02fF
C4223 AND2X1_LOC_794/A OR2X1_LOC_52/B 0.03fF
C4224 OR2X1_LOC_147/B AND2X1_LOC_3/Y 0.02fF
C4225 OR2X1_LOC_87/a_36_216# OR2X1_LOC_87/Y 0.00fF
C4226 OR2X1_LOC_26/Y AND2X1_LOC_400/a_8_24# 0.01fF
C4227 OR2X1_LOC_316/Y AND2X1_LOC_831/a_8_24# 0.01fF
C4228 OR2X1_LOC_358/a_36_216# OR2X1_LOC_130/A 0.01fF
C4229 OR2X1_LOC_68/B AND2X1_LOC_238/a_36_24# 0.00fF
C4230 OR2X1_LOC_316/Y OR2X1_LOC_44/Y 0.11fF
C4231 AND2X1_LOC_76/Y OR2X1_LOC_7/A 0.03fF
C4232 AND2X1_LOC_67/a_36_24# AND2X1_LOC_67/Y 0.01fF
C4233 OR2X1_LOC_748/A AND2X1_LOC_848/a_8_24# 0.01fF
C4234 AND2X1_LOC_696/a_8_24# OR2X1_LOC_161/A 0.02fF
C4235 OR2X1_LOC_644/B AND2X1_LOC_59/Y 0.14fF
C4236 OR2X1_LOC_602/Y AND2X1_LOC_600/a_36_24# 0.00fF
C4237 AND2X1_LOC_264/a_8_24# OR2X1_LOC_39/A 0.03fF
C4238 AND2X1_LOC_517/a_8_24# AND2X1_LOC_3/Y 0.01fF
C4239 OR2X1_LOC_773/B OR2X1_LOC_269/B 0.02fF
C4240 AND2X1_LOC_562/B OR2X1_LOC_64/Y 0.03fF
C4241 OR2X1_LOC_462/B AND2X1_LOC_56/B 0.03fF
C4242 AND2X1_LOC_42/B OR2X1_LOC_737/A 0.02fF
C4243 AND2X1_LOC_348/A OR2X1_LOC_481/A 0.02fF
C4244 OR2X1_LOC_3/Y OR2X1_LOC_48/B 0.15fF
C4245 OR2X1_LOC_47/Y AND2X1_LOC_475/Y 0.00fF
C4246 OR2X1_LOC_219/B OR2X1_LOC_215/Y 0.05fF
C4247 OR2X1_LOC_107/Y OR2X1_LOC_22/Y 0.03fF
C4248 AND2X1_LOC_767/a_8_24# OR2X1_LOC_287/B 0.01fF
C4249 OR2X1_LOC_460/Y OR2X1_LOC_463/a_8_216# 0.39fF
C4250 OR2X1_LOC_842/A AND2X1_LOC_47/Y 0.00fF
C4251 OR2X1_LOC_92/Y AND2X1_LOC_663/B 0.10fF
C4252 AND2X1_LOC_486/Y OR2X1_LOC_527/Y 0.07fF
C4253 OR2X1_LOC_262/a_8_216# OR2X1_LOC_85/A 0.01fF
C4254 AND2X1_LOC_724/Y OR2X1_LOC_95/Y 0.01fF
C4255 OR2X1_LOC_271/B OR2X1_LOC_271/Y 0.02fF
C4256 AND2X1_LOC_95/Y AND2X1_LOC_42/B 0.08fF
C4257 OR2X1_LOC_3/Y OR2X1_LOC_18/Y 9.00fF
C4258 OR2X1_LOC_462/B AND2X1_LOC_8/Y 0.02fF
C4259 OR2X1_LOC_116/a_36_216# OR2X1_LOC_87/A 0.02fF
C4260 OR2X1_LOC_26/Y AND2X1_LOC_287/Y 0.01fF
C4261 OR2X1_LOC_377/A OR2X1_LOC_557/A 0.00fF
C4262 OR2X1_LOC_633/Y AND2X1_LOC_42/B 0.03fF
C4263 OR2X1_LOC_532/B AND2X1_LOC_232/a_8_24# 0.00fF
C4264 AND2X1_LOC_813/a_8_24# AND2X1_LOC_18/Y 0.01fF
C4265 OR2X1_LOC_759/A GATE_662 0.01fF
C4266 AND2X1_LOC_852/Y OR2X1_LOC_69/Y 0.03fF
C4267 OR2X1_LOC_400/B OR2X1_LOC_403/B 0.00fF
C4268 OR2X1_LOC_643/A OR2X1_LOC_720/a_8_216# 0.02fF
C4269 OR2X1_LOC_174/Y OR2X1_LOC_175/a_8_216# 0.18fF
C4270 OR2X1_LOC_741/a_8_216# OR2X1_LOC_741/A 0.39fF
C4271 OR2X1_LOC_43/A OR2X1_LOC_827/a_36_216# 0.01fF
C4272 OR2X1_LOC_264/Y AND2X1_LOC_667/a_8_24# 0.03fF
C4273 AND2X1_LOC_363/A AND2X1_LOC_359/a_36_24# 0.00fF
C4274 OR2X1_LOC_814/A OR2X1_LOC_775/a_8_216# 0.11fF
C4275 AND2X1_LOC_525/a_8_24# OR2X1_LOC_87/A 0.05fF
C4276 AND2X1_LOC_64/Y OR2X1_LOC_317/B 0.03fF
C4277 OR2X1_LOC_486/a_36_216# OR2X1_LOC_739/A 0.00fF
C4278 OR2X1_LOC_158/A AND2X1_LOC_848/A 0.16fF
C4279 OR2X1_LOC_860/Y OR2X1_LOC_814/A 0.01fF
C4280 AND2X1_LOC_663/B OR2X1_LOC_65/B 0.01fF
C4281 AND2X1_LOC_569/A AND2X1_LOC_475/a_8_24# 0.19fF
C4282 AND2X1_LOC_476/Y OR2X1_LOC_406/A 0.01fF
C4283 D_INPUT_7 AND2X1_LOC_30/a_36_24# 0.00fF
C4284 OR2X1_LOC_695/a_36_216# AND2X1_LOC_687/B 0.00fF
C4285 AND2X1_LOC_366/a_36_24# OR2X1_LOC_47/Y 0.00fF
C4286 OR2X1_LOC_7/A OR2X1_LOC_52/B 4.28fF
C4287 AND2X1_LOC_390/B OR2X1_LOC_44/Y 0.07fF
C4288 OR2X1_LOC_427/A AND2X1_LOC_686/a_36_24# 0.00fF
C4289 VDD OR2X1_LOC_215/a_8_216# 0.00fF
C4290 AND2X1_LOC_543/Y OR2X1_LOC_437/A 0.02fF
C4291 AND2X1_LOC_64/Y OR2X1_LOC_580/A 0.00fF
C4292 OR2X1_LOC_585/A AND2X1_LOC_240/Y 0.01fF
C4293 AND2X1_LOC_173/a_8_24# OR2X1_LOC_532/B 0.00fF
C4294 OR2X1_LOC_168/B OR2X1_LOC_223/A 0.03fF
C4295 AND2X1_LOC_212/A AND2X1_LOC_222/Y 0.01fF
C4296 AND2X1_LOC_345/Y OR2X1_LOC_820/B 0.01fF
C4297 OR2X1_LOC_825/a_8_216# OR2X1_LOC_44/Y 0.00fF
C4298 AND2X1_LOC_91/B OR2X1_LOC_561/A 0.03fF
C4299 AND2X1_LOC_62/a_8_24# D_INPUT_0 0.01fF
C4300 VDD OR2X1_LOC_339/Y 0.12fF
C4301 AND2X1_LOC_12/Y AND2X1_LOC_48/A 0.22fF
C4302 OR2X1_LOC_87/A AND2X1_LOC_51/Y 0.55fF
C4303 OR2X1_LOC_158/A OR2X1_LOC_588/a_8_216# 0.05fF
C4304 AND2X1_LOC_387/B AND2X1_LOC_3/Y 0.04fF
C4305 OR2X1_LOC_46/A OR2X1_LOC_39/A 0.19fF
C4306 AND2X1_LOC_702/Y AND2X1_LOC_326/A 0.01fF
C4307 OR2X1_LOC_663/A OR2X1_LOC_227/Y 0.08fF
C4308 OR2X1_LOC_158/A AND2X1_LOC_203/a_8_24# 0.01fF
C4309 OR2X1_LOC_489/B OR2X1_LOC_814/A 0.00fF
C4310 AND2X1_LOC_95/Y OR2X1_LOC_286/B 0.36fF
C4311 AND2X1_LOC_434/Y OR2X1_LOC_311/a_8_216# 0.03fF
C4312 OR2X1_LOC_158/A AND2X1_LOC_206/Y 0.02fF
C4313 INPUT_1 AND2X1_LOC_43/B 0.04fF
C4314 OR2X1_LOC_139/A OR2X1_LOC_112/A 0.03fF
C4315 AND2X1_LOC_56/B AND2X1_LOC_27/a_36_24# 0.00fF
C4316 AND2X1_LOC_364/a_8_24# OR2X1_LOC_437/A 0.04fF
C4317 OR2X1_LOC_154/A AND2X1_LOC_79/a_36_24# 0.01fF
C4318 AND2X1_LOC_59/Y AND2X1_LOC_53/Y 0.07fF
C4319 OR2X1_LOC_129/a_8_216# OR2X1_LOC_80/A 0.01fF
C4320 OR2X1_LOC_53/a_8_216# OR2X1_LOC_409/B 0.00fF
C4321 OR2X1_LOC_599/A OR2X1_LOC_22/Y 0.09fF
C4322 OR2X1_LOC_154/A AND2X1_LOC_69/a_8_24# 0.01fF
C4323 OR2X1_LOC_196/B OR2X1_LOC_269/B 0.00fF
C4324 AND2X1_LOC_22/Y OR2X1_LOC_174/Y 0.37fF
C4325 OR2X1_LOC_147/B OR2X1_LOC_270/Y 0.03fF
C4326 AND2X1_LOC_227/Y OR2X1_LOC_39/A 0.00fF
C4327 AND2X1_LOC_611/a_8_24# OR2X1_LOC_54/Y 0.01fF
C4328 OR2X1_LOC_476/Y OR2X1_LOC_475/Y 0.06fF
C4329 OR2X1_LOC_62/a_36_216# OR2X1_LOC_753/A 0.00fF
C4330 AND2X1_LOC_211/B OR2X1_LOC_46/A 0.07fF
C4331 OR2X1_LOC_437/A OR2X1_LOC_322/Y 0.19fF
C4332 OR2X1_LOC_559/B AND2X1_LOC_88/Y 0.03fF
C4333 OR2X1_LOC_31/Y OR2X1_LOC_6/A 0.83fF
C4334 AND2X1_LOC_59/Y OR2X1_LOC_223/A 0.04fF
C4335 AND2X1_LOC_170/B AND2X1_LOC_661/A 0.11fF
C4336 OR2X1_LOC_19/B OR2X1_LOC_83/a_8_216# 0.09fF
C4337 OR2X1_LOC_62/B OR2X1_LOC_278/a_8_216# 0.03fF
C4338 OR2X1_LOC_485/A AND2X1_LOC_539/a_8_24# 0.01fF
C4339 AND2X1_LOC_329/a_8_24# OR2X1_LOC_532/B 0.01fF
C4340 OR2X1_LOC_139/a_36_216# OR2X1_LOC_244/A 0.00fF
C4341 OR2X1_LOC_600/A OR2X1_LOC_385/a_8_216# 0.14fF
C4342 AND2X1_LOC_394/a_36_24# OR2X1_LOC_84/A 0.01fF
C4343 AND2X1_LOC_41/A OR2X1_LOC_68/B 0.06fF
C4344 OR2X1_LOC_709/A OR2X1_LOC_703/Y 0.04fF
C4345 AND2X1_LOC_66/a_36_24# OR2X1_LOC_13/B 0.00fF
C4346 AND2X1_LOC_731/a_8_24# AND2X1_LOC_220/B 0.07fF
C4347 OR2X1_LOC_413/Y AND2X1_LOC_461/a_8_24# 0.01fF
C4348 AND2X1_LOC_316/a_8_24# AND2X1_LOC_31/Y 0.01fF
C4349 OR2X1_LOC_433/a_8_216# AND2X1_LOC_648/B 0.00fF
C4350 D_INPUT_3 OR2X1_LOC_6/a_8_216# 0.01fF
C4351 INPUT_1 OR2X1_LOC_27/a_8_216# 0.01fF
C4352 AND2X1_LOC_564/A AND2X1_LOC_220/B 0.03fF
C4353 D_INPUT_4 AND2X1_LOC_31/Y 0.02fF
C4354 OR2X1_LOC_185/Y D_INPUT_1 0.07fF
C4355 AND2X1_LOC_64/Y AND2X1_LOC_44/Y 0.98fF
C4356 OR2X1_LOC_711/B OR2X1_LOC_308/Y 0.04fF
C4357 AND2X1_LOC_465/a_8_24# OR2X1_LOC_31/Y 0.02fF
C4358 OR2X1_LOC_785/B OR2X1_LOC_228/Y 0.00fF
C4359 OR2X1_LOC_45/B AND2X1_LOC_227/a_8_24# 0.17fF
C4360 OR2X1_LOC_19/B OR2X1_LOC_750/A 0.05fF
C4361 OR2X1_LOC_95/Y OR2X1_LOC_371/Y 0.10fF
C4362 AND2X1_LOC_423/a_8_24# OR2X1_LOC_724/A 0.03fF
C4363 AND2X1_LOC_86/Y OR2X1_LOC_398/Y 0.03fF
C4364 AND2X1_LOC_382/a_36_24# D_INPUT_1 0.00fF
C4365 OR2X1_LOC_175/Y OR2X1_LOC_857/A 0.18fF
C4366 AND2X1_LOC_671/a_36_24# OR2X1_LOC_54/Y 0.01fF
C4367 AND2X1_LOC_597/a_36_24# OR2X1_LOC_214/B 0.01fF
C4368 AND2X1_LOC_293/a_8_24# OR2X1_LOC_27/Y 0.25fF
C4369 OR2X1_LOC_78/B OR2X1_LOC_537/a_8_216# 0.04fF
C4370 AND2X1_LOC_59/Y AND2X1_LOC_609/a_8_24# 0.10fF
C4371 AND2X1_LOC_807/Y AND2X1_LOC_222/Y 0.16fF
C4372 OR2X1_LOC_70/Y AND2X1_LOC_451/Y 0.01fF
C4373 OR2X1_LOC_819/a_8_216# OR2X1_LOC_749/Y 0.40fF
C4374 AND2X1_LOC_22/Y OR2X1_LOC_855/a_8_216# 0.03fF
C4375 OR2X1_LOC_269/B AND2X1_LOC_225/a_36_24# 0.00fF
C4376 OR2X1_LOC_820/a_8_216# OR2X1_LOC_748/a_8_216# 0.47fF
C4377 OR2X1_LOC_338/a_8_216# OR2X1_LOC_338/A 0.06fF
C4378 OR2X1_LOC_70/Y AND2X1_LOC_648/B 0.02fF
C4379 OR2X1_LOC_696/A OR2X1_LOC_600/A 10.88fF
C4380 OR2X1_LOC_662/A OR2X1_LOC_68/B 0.07fF
C4381 OR2X1_LOC_3/Y AND2X1_LOC_620/Y 0.03fF
C4382 OR2X1_LOC_696/A AND2X1_LOC_335/Y 0.12fF
C4383 VDD OR2X1_LOC_731/A 0.12fF
C4384 OR2X1_LOC_74/A AND2X1_LOC_792/Y 0.14fF
C4385 AND2X1_LOC_631/Y AND2X1_LOC_620/Y 0.01fF
C4386 AND2X1_LOC_632/a_36_24# OR2X1_LOC_615/Y 0.00fF
C4387 OR2X1_LOC_324/B OR2X1_LOC_308/Y 0.14fF
C4388 OR2X1_LOC_653/A AND2X1_LOC_31/Y 0.03fF
C4389 OR2X1_LOC_160/B OR2X1_LOC_338/B 0.01fF
C4390 OR2X1_LOC_756/B OR2X1_LOC_593/B 0.00fF
C4391 OR2X1_LOC_7/A AND2X1_LOC_216/A 0.15fF
C4392 OR2X1_LOC_186/Y OR2X1_LOC_337/A 0.01fF
C4393 OR2X1_LOC_22/Y AND2X1_LOC_866/A 0.07fF
C4394 OR2X1_LOC_654/A OR2X1_LOC_598/A 0.03fF
C4395 OR2X1_LOC_866/a_8_216# OR2X1_LOC_561/B 0.02fF
C4396 OR2X1_LOC_516/Y AND2X1_LOC_574/a_8_24# 0.00fF
C4397 OR2X1_LOC_26/Y AND2X1_LOC_562/Y 0.03fF
C4398 AND2X1_LOC_110/Y OR2X1_LOC_703/a_36_216# 0.00fF
C4399 OR2X1_LOC_703/A OR2X1_LOC_703/Y 0.01fF
C4400 OR2X1_LOC_375/A OR2X1_LOC_725/a_8_216# 0.01fF
C4401 AND2X1_LOC_771/B AND2X1_LOC_774/A -0.00fF
C4402 OR2X1_LOC_631/B OR2X1_LOC_68/B 0.03fF
C4403 AND2X1_LOC_776/a_8_24# AND2X1_LOC_564/B 0.01fF
C4404 OR2X1_LOC_843/B OR2X1_LOC_349/A 0.03fF
C4405 OR2X1_LOC_89/A AND2X1_LOC_562/Y 0.10fF
C4406 AND2X1_LOC_388/Y AND2X1_LOC_810/B 0.01fF
C4407 OR2X1_LOC_709/A OR2X1_LOC_596/A 0.08fF
C4408 OR2X1_LOC_696/A AND2X1_LOC_543/a_8_24# 0.02fF
C4409 OR2X1_LOC_375/A OR2X1_LOC_546/a_8_216# 0.01fF
C4410 AND2X1_LOC_465/A OR2X1_LOC_59/Y 0.07fF
C4411 AND2X1_LOC_721/Y AND2X1_LOC_657/Y 0.03fF
C4412 AND2X1_LOC_469/Y AND2X1_LOC_220/a_8_24# 0.20fF
C4413 OR2X1_LOC_494/A OR2X1_LOC_56/A 0.08fF
C4414 OR2X1_LOC_421/A OR2X1_LOC_12/Y 0.02fF
C4415 OR2X1_LOC_53/Y AND2X1_LOC_434/Y 0.02fF
C4416 OR2X1_LOC_181/B AND2X1_LOC_36/Y 0.18fF
C4417 OR2X1_LOC_502/A OR2X1_LOC_356/B 0.63fF
C4418 OR2X1_LOC_13/Y AND2X1_LOC_193/Y 0.01fF
C4419 OR2X1_LOC_235/B OR2X1_LOC_392/B 0.03fF
C4420 OR2X1_LOC_43/A OR2X1_LOC_437/A 0.22fF
C4421 AND2X1_LOC_318/Y AND2X1_LOC_476/A 0.26fF
C4422 AND2X1_LOC_60/a_8_24# OR2X1_LOC_78/B 0.03fF
C4423 OR2X1_LOC_161/A OR2X1_LOC_844/B 0.02fF
C4424 OR2X1_LOC_235/B AND2X1_LOC_263/a_8_24# 0.02fF
C4425 AND2X1_LOC_802/Y AND2X1_LOC_434/Y 0.02fF
C4426 OR2X1_LOC_114/a_8_216# AND2X1_LOC_22/Y 0.07fF
C4427 OR2X1_LOC_78/A OR2X1_LOC_580/B 0.03fF
C4428 AND2X1_LOC_745/a_8_24# VDD 0.00fF
C4429 OR2X1_LOC_406/Y AND2X1_LOC_734/Y 0.01fF
C4430 OR2X1_LOC_696/A OR2X1_LOC_619/Y 0.15fF
C4431 VDD OR2X1_LOC_596/a_8_216# 0.21fF
C4432 OR2X1_LOC_696/A AND2X1_LOC_356/a_8_24# 0.03fF
C4433 OR2X1_LOC_643/Y OR2X1_LOC_228/Y 0.02fF
C4434 OR2X1_LOC_6/B VDD 0.85fF
C4435 AND2X1_LOC_40/Y OR2X1_LOC_563/A 0.11fF
C4436 AND2X1_LOC_713/Y VDD 0.38fF
C4437 OR2X1_LOC_178/a_8_216# OR2X1_LOC_108/Y -0.01fF
C4438 OR2X1_LOC_96/Y AND2X1_LOC_98/a_8_24# 0.00fF
C4439 OR2X1_LOC_656/Y AND2X1_LOC_44/Y 0.02fF
C4440 OR2X1_LOC_164/Y AND2X1_LOC_786/Y 0.01fF
C4441 OR2X1_LOC_512/A AND2X1_LOC_44/Y 0.01fF
C4442 AND2X1_LOC_40/Y OR2X1_LOC_357/B 0.23fF
C4443 OR2X1_LOC_8/Y OR2X1_LOC_822/a_8_216# 0.01fF
C4444 OR2X1_LOC_93/Y OR2X1_LOC_51/Y 0.01fF
C4445 OR2X1_LOC_287/B OR2X1_LOC_576/a_36_216# 0.00fF
C4446 OR2X1_LOC_604/A AND2X1_LOC_160/Y 0.01fF
C4447 AND2X1_LOC_460/a_8_24# OR2X1_LOC_588/A 0.10fF
C4448 OR2X1_LOC_244/A OR2X1_LOC_398/Y 0.03fF
C4449 OR2X1_LOC_516/Y OR2X1_LOC_497/Y 0.02fF
C4450 AND2X1_LOC_212/A AND2X1_LOC_367/A 0.42fF
C4451 OR2X1_LOC_40/Y AND2X1_LOC_514/a_8_24# 0.02fF
C4452 AND2X1_LOC_217/Y OR2X1_LOC_132/Y 0.01fF
C4453 AND2X1_LOC_778/a_36_24# OR2X1_LOC_680/A 0.01fF
C4454 OR2X1_LOC_372/a_36_216# OR2X1_LOC_437/A 0.15fF
C4455 AND2X1_LOC_508/B AND2X1_LOC_508/a_8_24# 0.00fF
C4456 OR2X1_LOC_308/A OR2X1_LOC_375/A 0.00fF
C4457 OR2X1_LOC_51/Y AND2X1_LOC_334/Y 0.03fF
C4458 AND2X1_LOC_566/B AND2X1_LOC_365/a_36_24# 0.00fF
C4459 AND2X1_LOC_357/B AND2X1_LOC_364/Y 0.01fF
C4460 OR2X1_LOC_122/a_8_216# OR2X1_LOC_600/A 0.05fF
C4461 OR2X1_LOC_95/Y AND2X1_LOC_222/Y 0.03fF
C4462 AND2X1_LOC_321/a_36_24# AND2X1_LOC_44/Y 0.00fF
C4463 AND2X1_LOC_20/a_8_24# AND2X1_LOC_18/Y -0.00fF
C4464 AND2X1_LOC_440/a_8_24# AND2X1_LOC_222/Y 0.01fF
C4465 OR2X1_LOC_563/B OR2X1_LOC_577/B 0.88fF
C4466 OR2X1_LOC_3/a_8_216# D_INPUT_6 0.01fF
C4467 OR2X1_LOC_555/B AND2X1_LOC_44/Y 0.09fF
C4468 AND2X1_LOC_841/B OR2X1_LOC_323/Y 0.00fF
C4469 OR2X1_LOC_555/B OR2X1_LOC_555/a_8_216# 0.07fF
C4470 OR2X1_LOC_51/Y OR2X1_LOC_743/a_36_216# 0.00fF
C4471 OR2X1_LOC_643/A OR2X1_LOC_115/B 0.83fF
C4472 OR2X1_LOC_691/Y OR2X1_LOC_793/a_8_216# 0.01fF
C4473 OR2X1_LOC_45/B OR2X1_LOC_316/Y 0.06fF
C4474 OR2X1_LOC_709/A OR2X1_LOC_732/a_8_216# 0.04fF
C4475 OR2X1_LOC_421/A OR2X1_LOC_763/a_36_216# 0.00fF
C4476 AND2X1_LOC_12/Y OR2X1_LOC_34/a_8_216# 0.01fF
C4477 AND2X1_LOC_51/Y OR2X1_LOC_579/A 0.26fF
C4478 AND2X1_LOC_12/Y OR2X1_LOC_489/A 0.00fF
C4479 AND2X1_LOC_764/a_8_24# OR2X1_LOC_637/Y 0.24fF
C4480 OR2X1_LOC_345/Y AND2X1_LOC_12/Y 0.01fF
C4481 VDD OR2X1_LOC_441/Y 0.48fF
C4482 AND2X1_LOC_786/a_8_24# OR2X1_LOC_36/Y 0.02fF
C4483 AND2X1_LOC_737/Y OR2X1_LOC_40/Y 0.01fF
C4484 OR2X1_LOC_756/B OR2X1_LOC_645/a_36_216# 0.00fF
C4485 OR2X1_LOC_786/Y OR2X1_LOC_228/Y 0.01fF
C4486 AND2X1_LOC_392/A OR2X1_LOC_92/Y 0.14fF
C4487 AND2X1_LOC_70/Y OR2X1_LOC_808/A 0.46fF
C4488 OR2X1_LOC_48/B AND2X1_LOC_477/Y 0.07fF
C4489 OR2X1_LOC_186/Y OR2X1_LOC_539/Y 0.05fF
C4490 AND2X1_LOC_571/a_8_24# OR2X1_LOC_44/Y 0.03fF
C4491 OR2X1_LOC_404/Y OR2X1_LOC_500/a_8_216# 0.02fF
C4492 OR2X1_LOC_249/Y OR2X1_LOC_343/a_8_216# 0.13fF
C4493 OR2X1_LOC_165/a_8_216# OR2X1_LOC_40/Y 0.01fF
C4494 OR2X1_LOC_375/A OR2X1_LOC_160/Y 0.00fF
C4495 OR2X1_LOC_326/B OR2X1_LOC_302/A 0.01fF
C4496 OR2X1_LOC_36/Y AND2X1_LOC_455/B 0.07fF
C4497 AND2X1_LOC_300/a_8_24# AND2X1_LOC_43/B 0.04fF
C4498 OR2X1_LOC_326/B VDD 0.08fF
C4499 OR2X1_LOC_667/Y VDD 0.12fF
C4500 OR2X1_LOC_151/A OR2X1_LOC_510/Y 0.15fF
C4501 AND2X1_LOC_639/A D_INPUT_6 0.10fF
C4502 OR2X1_LOC_656/B OR2X1_LOC_160/B 0.07fF
C4503 OR2X1_LOC_160/A OR2X1_LOC_641/A 0.03fF
C4504 AND2X1_LOC_51/Y OR2X1_LOC_390/B 0.29fF
C4505 OR2X1_LOC_156/a_36_216# OR2X1_LOC_479/Y 0.02fF
C4506 AND2X1_LOC_465/a_36_24# AND2X1_LOC_465/A 0.01fF
C4507 AND2X1_LOC_12/Y OR2X1_LOC_772/A 0.00fF
C4508 OR2X1_LOC_834/a_8_216# AND2X1_LOC_41/A 0.01fF
C4509 OR2X1_LOC_434/A OR2X1_LOC_174/Y 0.12fF
C4510 OR2X1_LOC_168/B OR2X1_LOC_502/A 0.00fF
C4511 OR2X1_LOC_519/Y VDD 0.09fF
C4512 AND2X1_LOC_851/a_8_24# OR2X1_LOC_495/Y 0.01fF
C4513 AND2X1_LOC_738/B OR2X1_LOC_427/A 0.09fF
C4514 OR2X1_LOC_679/a_8_216# OR2X1_LOC_679/B 0.01fF
C4515 AND2X1_LOC_767/a_8_24# OR2X1_LOC_160/B 0.04fF
C4516 AND2X1_LOC_392/A OR2X1_LOC_65/B 2.46fF
C4517 OR2X1_LOC_427/A OR2X1_LOC_56/A 5.92fF
C4518 AND2X1_LOC_366/A OR2X1_LOC_92/Y 0.00fF
C4519 OR2X1_LOC_389/A OR2X1_LOC_161/A 0.01fF
C4520 AND2X1_LOC_338/Y AND2X1_LOC_640/Y 0.00fF
C4521 AND2X1_LOC_99/A OR2X1_LOC_666/A 0.37fF
C4522 OR2X1_LOC_499/B OR2X1_LOC_274/Y 0.05fF
C4523 OR2X1_LOC_74/A OR2X1_LOC_816/A 0.04fF
C4524 AND2X1_LOC_22/Y AND2X1_LOC_42/B 0.52fF
C4525 OR2X1_LOC_109/Y OR2X1_LOC_51/Y 0.07fF
C4526 OR2X1_LOC_677/Y OR2X1_LOC_441/Y 0.03fF
C4527 AND2X1_LOC_719/Y AND2X1_LOC_576/Y 0.10fF
C4528 VDD AND2X1_LOC_436/B 0.39fF
C4529 OR2X1_LOC_778/a_8_216# OR2X1_LOC_737/A 0.03fF
C4530 OR2X1_LOC_696/A OR2X1_LOC_22/A 0.00fF
C4531 OR2X1_LOC_45/B AND2X1_LOC_390/B 0.07fF
C4532 OR2X1_LOC_329/B OR2X1_LOC_48/B 0.14fF
C4533 VDD AND2X1_LOC_139/B 0.30fF
C4534 OR2X1_LOC_51/Y AND2X1_LOC_448/Y 0.03fF
C4535 AND2X1_LOC_95/Y OR2X1_LOC_363/A 0.09fF
C4536 OR2X1_LOC_121/Y AND2X1_LOC_3/Y 0.08fF
C4537 AND2X1_LOC_504/a_8_24# OR2X1_LOC_78/B 0.18fF
C4538 AND2X1_LOC_340/Y OR2X1_LOC_3/Y 0.01fF
C4539 OR2X1_LOC_89/A OR2X1_LOC_381/a_8_216# 0.01fF
C4540 OR2X1_LOC_151/A OR2X1_LOC_810/A 0.10fF
C4541 OR2X1_LOC_759/A AND2X1_LOC_580/A 0.03fF
C4542 OR2X1_LOC_129/a_36_216# OR2X1_LOC_69/Y 0.00fF
C4543 VDD OR2X1_LOC_579/B 0.06fF
C4544 AND2X1_LOC_84/Y OR2X1_LOC_65/Y 0.01fF
C4545 OR2X1_LOC_329/B OR2X1_LOC_18/Y 0.12fF
C4546 AND2X1_LOC_858/B AND2X1_LOC_621/Y 0.03fF
C4547 OR2X1_LOC_744/A AND2X1_LOC_403/B 0.01fF
C4548 OR2X1_LOC_663/a_36_216# OR2X1_LOC_557/A 0.00fF
C4549 AND2X1_LOC_799/a_36_24# OR2X1_LOC_417/Y 0.01fF
C4550 OR2X1_LOC_845/a_8_216# AND2X1_LOC_18/Y 0.02fF
C4551 OR2X1_LOC_604/A AND2X1_LOC_580/B 0.02fF
C4552 AND2X1_LOC_172/a_8_24# OR2X1_LOC_358/B 0.01fF
C4553 AND2X1_LOC_758/a_8_24# AND2X1_LOC_580/B 0.01fF
C4554 AND2X1_LOC_363/a_8_24# OR2X1_LOC_3/Y 0.01fF
C4555 AND2X1_LOC_464/a_8_24# OR2X1_LOC_56/A 0.01fF
C4556 VDD OR2X1_LOC_235/Y 0.12fF
C4557 OR2X1_LOC_45/B OR2X1_LOC_431/Y 0.02fF
C4558 AND2X1_LOC_387/a_8_24# OR2X1_LOC_269/B 0.01fF
C4559 OR2X1_LOC_862/B OR2X1_LOC_561/a_8_216# 0.03fF
C4560 OR2X1_LOC_7/A OR2X1_LOC_253/Y 0.00fF
C4561 AND2X1_LOC_95/Y OR2X1_LOC_663/A 0.05fF
C4562 OR2X1_LOC_844/a_8_216# OR2X1_LOC_113/B 0.01fF
C4563 OR2X1_LOC_114/B AND2X1_LOC_292/a_36_24# 0.00fF
C4564 OR2X1_LOC_462/B AND2X1_LOC_92/Y 0.35fF
C4565 D_INPUT_0 OR2X1_LOC_415/Y 0.00fF
C4566 OR2X1_LOC_377/A OR2X1_LOC_39/Y 0.14fF
C4567 OR2X1_LOC_47/Y OR2X1_LOC_386/a_8_216# 0.01fF
C4568 AND2X1_LOC_12/Y OR2X1_LOC_859/a_8_216# 0.01fF
C4569 AND2X1_LOC_354/Y OR2X1_LOC_92/Y 0.11fF
C4570 OR2X1_LOC_47/Y OR2X1_LOC_183/Y 0.23fF
C4571 AND2X1_LOC_12/Y OR2X1_LOC_201/A 0.01fF
C4572 AND2X1_LOC_191/B OR2X1_LOC_748/A 0.08fF
C4573 OR2X1_LOC_114/B AND2X1_LOC_3/Y 0.06fF
C4574 OR2X1_LOC_814/A AND2X1_LOC_7/B 0.45fF
C4575 OR2X1_LOC_427/A OR2X1_LOC_426/Y 0.01fF
C4576 AND2X1_LOC_41/A OR2X1_LOC_219/a_8_216# 0.03fF
C4577 AND2X1_LOC_856/a_36_24# OR2X1_LOC_428/A 0.01fF
C4578 AND2X1_LOC_501/Y AND2X1_LOC_474/Y 0.02fF
C4579 AND2X1_LOC_41/A OR2X1_LOC_241/a_8_216# 0.01fF
C4580 OR2X1_LOC_744/A OR2X1_LOC_44/Y 0.89fF
C4581 AND2X1_LOC_624/A OR2X1_LOC_746/a_8_216# 0.01fF
C4582 OR2X1_LOC_154/A AND2X1_LOC_65/a_8_24# 0.03fF
C4583 AND2X1_LOC_363/A OR2X1_LOC_56/A 0.03fF
C4584 OR2X1_LOC_2/Y OR2X1_LOC_30/a_8_216# 0.02fF
C4585 VDD OR2X1_LOC_529/Y 0.57fF
C4586 AND2X1_LOC_396/a_8_24# AND2X1_LOC_3/Y 0.02fF
C4587 AND2X1_LOC_570/Y AND2X1_LOC_474/Y 0.03fF
C4588 OR2X1_LOC_139/A AND2X1_LOC_667/a_36_24# 0.00fF
C4589 AND2X1_LOC_59/Y OR2X1_LOC_502/A 0.62fF
C4590 OR2X1_LOC_660/a_8_216# OR2X1_LOC_660/B 0.05fF
C4591 OR2X1_LOC_756/B OR2X1_LOC_270/a_36_216# 0.00fF
C4592 OR2X1_LOC_220/A OR2X1_LOC_375/A 0.05fF
C4593 OR2X1_LOC_6/B OR2X1_LOC_826/a_8_216# 0.07fF
C4594 AND2X1_LOC_570/Y OR2X1_LOC_485/A 0.05fF
C4595 OR2X1_LOC_250/Y OR2X1_LOC_278/Y 0.18fF
C4596 OR2X1_LOC_497/Y AND2X1_LOC_842/a_8_24# 0.02fF
C4597 OR2X1_LOC_331/A OR2X1_LOC_485/A 0.06fF
C4598 D_INPUT_0 AND2X1_LOC_786/Y 0.07fF
C4599 AND2X1_LOC_329/a_36_24# OR2X1_LOC_78/A 0.01fF
C4600 AND2X1_LOC_474/A OR2X1_LOC_106/A 0.00fF
C4601 OR2X1_LOC_160/A OR2X1_LOC_730/a_8_216# 0.03fF
C4602 AND2X1_LOC_729/Y AND2X1_LOC_841/B 0.07fF
C4603 OR2X1_LOC_154/A OR2X1_LOC_403/A 0.07fF
C4604 AND2X1_LOC_566/B AND2X1_LOC_537/Y 0.16fF
C4605 OR2X1_LOC_379/Y OR2X1_LOC_160/A 0.16fF
C4606 OR2X1_LOC_600/A AND2X1_LOC_663/B 6.90fF
C4607 OR2X1_LOC_391/B OR2X1_LOC_392/A 0.05fF
C4608 OR2X1_LOC_604/A OR2X1_LOC_295/a_8_216# 0.11fF
C4609 OR2X1_LOC_557/A OR2X1_LOC_78/B 0.06fF
C4610 OR2X1_LOC_538/A AND2X1_LOC_3/Y 0.03fF
C4611 AND2X1_LOC_33/Y OR2X1_LOC_18/Y 0.02fF
C4612 OR2X1_LOC_597/A OR2X1_LOC_64/Y 0.01fF
C4613 AND2X1_LOC_387/B INPUT_0 0.07fF
C4614 AND2X1_LOC_621/Y AND2X1_LOC_573/A 0.03fF
C4615 OR2X1_LOC_184/Y AND2X1_LOC_465/A 0.06fF
C4616 AND2X1_LOC_31/Y OR2X1_LOC_723/B 0.03fF
C4617 AND2X1_LOC_504/a_8_24# OR2X1_LOC_375/A 0.11fF
C4618 OR2X1_LOC_51/Y AND2X1_LOC_729/B 0.03fF
C4619 OR2X1_LOC_185/Y OR2X1_LOC_737/A 0.07fF
C4620 AND2X1_LOC_486/Y AND2X1_LOC_806/A 0.01fF
C4621 OR2X1_LOC_40/Y OR2X1_LOC_22/Y 0.25fF
C4622 OR2X1_LOC_160/B AND2X1_LOC_45/a_8_24# 0.09fF
C4623 OR2X1_LOC_617/Y AND2X1_LOC_663/A 0.17fF
C4624 AND2X1_LOC_302/a_8_24# OR2X1_LOC_619/Y 0.02fF
C4625 OR2X1_LOC_43/A OR2X1_LOC_761/Y 0.01fF
C4626 AND2X1_LOC_563/a_8_24# AND2X1_LOC_572/Y 0.02fF
C4627 OR2X1_LOC_244/B AND2X1_LOC_42/B 0.06fF
C4628 AND2X1_LOC_672/B INPUT_2 0.01fF
C4629 AND2X1_LOC_41/A AND2X1_LOC_697/a_8_24# 0.04fF
C4630 AND2X1_LOC_474/A OR2X1_LOC_279/a_36_216# 0.00fF
C4631 OR2X1_LOC_36/Y OR2X1_LOC_278/Y 0.03fF
C4632 OR2X1_LOC_364/A AND2X1_LOC_95/Y 0.26fF
C4633 AND2X1_LOC_784/A AND2X1_LOC_841/B 0.07fF
C4634 OR2X1_LOC_154/A OR2X1_LOC_447/a_8_216# 0.04fF
C4635 OR2X1_LOC_185/Y AND2X1_LOC_95/Y 0.08fF
C4636 D_INPUT_5 AND2X1_LOC_3/Y 0.09fF
C4637 AND2X1_LOC_787/A OR2X1_LOC_437/a_8_216# 0.10fF
C4638 AND2X1_LOC_214/A OR2X1_LOC_52/a_8_216# 0.01fF
C4639 AND2X1_LOC_711/a_8_24# AND2X1_LOC_663/B 0.01fF
C4640 OR2X1_LOC_36/Y AND2X1_LOC_662/B 0.03fF
C4641 OR2X1_LOC_479/a_36_216# AND2X1_LOC_92/Y 0.01fF
C4642 OR2X1_LOC_70/Y AND2X1_LOC_477/a_8_24# 0.04fF
C4643 AND2X1_LOC_857/Y OR2X1_LOC_299/Y 0.21fF
C4644 OR2X1_LOC_667/Y OR2X1_LOC_251/Y 0.01fF
C4645 D_INPUT_0 OR2X1_LOC_631/A 0.00fF
C4646 AND2X1_LOC_578/A OR2X1_LOC_164/Y 0.13fF
C4647 AND2X1_LOC_41/A AND2X1_LOC_666/a_8_24# 0.10fF
C4648 VDD OR2X1_LOC_68/Y 0.16fF
C4649 OR2X1_LOC_578/B OR2X1_LOC_180/B 0.00fF
C4650 OR2X1_LOC_160/A OR2X1_LOC_114/Y 0.04fF
C4651 OR2X1_LOC_861/a_8_216# OR2X1_LOC_287/B 0.01fF
C4652 OR2X1_LOC_318/a_8_216# OR2X1_LOC_223/A 0.01fF
C4653 OR2X1_LOC_154/A OR2X1_LOC_130/A 0.17fF
C4654 OR2X1_LOC_517/A AND2X1_LOC_660/Y 0.01fF
C4655 OR2X1_LOC_26/Y AND2X1_LOC_287/a_8_24# 0.02fF
C4656 OR2X1_LOC_599/A OR2X1_LOC_39/A 0.07fF
C4657 OR2X1_LOC_262/Y OR2X1_LOC_118/Y 0.00fF
C4658 OR2X1_LOC_160/A OR2X1_LOC_449/A 0.01fF
C4659 AND2X1_LOC_177/a_8_24# AND2X1_LOC_51/Y 0.03fF
C4660 AND2X1_LOC_502/a_36_24# OR2X1_LOC_36/Y 0.01fF
C4661 OR2X1_LOC_70/Y OR2X1_LOC_265/a_8_216# 0.01fF
C4662 OR2X1_LOC_285/a_8_216# OR2X1_LOC_285/B 0.03fF
C4663 AND2X1_LOC_65/A OR2X1_LOC_340/a_8_216# 0.06fF
C4664 AND2X1_LOC_11/Y AND2X1_LOC_18/a_8_24# 0.11fF
C4665 VDD AND2X1_LOC_47/Y 1.73fF
C4666 OR2X1_LOC_643/A OR2X1_LOC_222/A 0.00fF
C4667 OR2X1_LOC_643/a_8_216# OR2X1_LOC_215/Y 0.01fF
C4668 OR2X1_LOC_467/A OR2X1_LOC_446/Y 0.00fF
C4669 VDD D_GATE_222 0.04fF
C4670 INPUT_1 AND2X1_LOC_219/Y 0.01fF
C4671 AND2X1_LOC_12/Y AND2X1_LOC_3/Y 1.25fF
C4672 AND2X1_LOC_500/a_8_24# AND2X1_LOC_576/Y 0.02fF
C4673 AND2X1_LOC_84/Y OR2X1_LOC_72/Y 0.03fF
C4674 AND2X1_LOC_573/a_36_24# AND2X1_LOC_474/Y 0.00fF
C4675 OR2X1_LOC_669/Y AND2X1_LOC_668/a_8_24# 0.01fF
C4676 OR2X1_LOC_774/Y OR2X1_LOC_865/Y 0.01fF
C4677 AND2X1_LOC_514/Y AND2X1_LOC_863/a_8_24# 0.01fF
C4678 AND2X1_LOC_141/a_8_24# AND2X1_LOC_656/Y 0.23fF
C4679 OR2X1_LOC_864/A OR2X1_LOC_673/Y 0.03fF
C4680 OR2X1_LOC_36/Y AND2X1_LOC_472/B 5.47fF
C4681 AND2X1_LOC_807/Y OR2X1_LOC_74/A 3.12fF
C4682 OR2X1_LOC_557/A OR2X1_LOC_375/A 0.03fF
C4683 AND2X1_LOC_148/Y AND2X1_LOC_624/A 0.11fF
C4684 OR2X1_LOC_43/A OR2X1_LOC_753/A 0.10fF
C4685 OR2X1_LOC_40/Y AND2X1_LOC_808/A 0.03fF
C4686 OR2X1_LOC_235/B OR2X1_LOC_532/B 0.06fF
C4687 AND2X1_LOC_91/B OR2X1_LOC_80/A 0.12fF
C4688 OR2X1_LOC_865/B AND2X1_LOC_51/Y 0.04fF
C4689 AND2X1_LOC_731/Y GATE_811 0.02fF
C4690 OR2X1_LOC_639/B OR2X1_LOC_636/A 0.08fF
C4691 OR2X1_LOC_160/A OR2X1_LOC_201/Y 0.00fF
C4692 AND2X1_LOC_153/a_8_24# AND2X1_LOC_42/B 0.11fF
C4693 OR2X1_LOC_45/B OR2X1_LOC_153/a_8_216# 0.06fF
C4694 OR2X1_LOC_87/A OR2X1_LOC_787/Y 0.07fF
C4695 AND2X1_LOC_117/a_8_24# OR2X1_LOC_375/A 0.01fF
C4696 AND2X1_LOC_76/Y AND2X1_LOC_115/a_8_24# 0.00fF
C4697 OR2X1_LOC_32/a_8_216# OR2X1_LOC_52/B 0.01fF
C4698 AND2X1_LOC_367/A OR2X1_LOC_95/Y 0.05fF
C4699 OR2X1_LOC_216/Y OR2X1_LOC_216/a_8_216# 0.02fF
C4700 OR2X1_LOC_559/B OR2X1_LOC_121/B 0.01fF
C4701 OR2X1_LOC_26/Y AND2X1_LOC_634/a_36_24# 0.00fF
C4702 OR2X1_LOC_856/B OR2X1_LOC_750/a_8_216# 0.03fF
C4703 OR2X1_LOC_529/Y OR2X1_LOC_491/Y 0.01fF
C4704 AND2X1_LOC_95/Y OR2X1_LOC_472/B 0.02fF
C4705 OR2X1_LOC_598/a_36_216# OR2X1_LOC_771/B 0.01fF
C4706 AND2X1_LOC_53/Y OR2X1_LOC_623/B 0.51fF
C4707 OR2X1_LOC_66/a_8_216# OR2X1_LOC_66/A 0.04fF
C4708 OR2X1_LOC_273/Y OR2X1_LOC_36/Y 0.73fF
C4709 AND2X1_LOC_59/Y AND2X1_LOC_518/a_8_24# 0.03fF
C4710 OR2X1_LOC_455/a_8_216# OR2X1_LOC_455/A 0.39fF
C4711 OR2X1_LOC_243/A OR2X1_LOC_19/B 0.00fF
C4712 OR2X1_LOC_377/A OR2X1_LOC_46/A 0.14fF
C4713 OR2X1_LOC_723/a_8_216# OR2X1_LOC_723/A 0.39fF
C4714 OR2X1_LOC_3/Y OR2X1_LOC_585/A 0.21fF
C4715 OR2X1_LOC_280/Y OR2X1_LOC_7/A 0.07fF
C4716 OR2X1_LOC_485/a_8_216# OR2X1_LOC_31/Y 0.01fF
C4717 AND2X1_LOC_59/Y AND2X1_LOC_48/A 2.09fF
C4718 VDD OR2X1_LOC_598/A 0.98fF
C4719 OR2X1_LOC_362/a_8_216# OR2X1_LOC_580/A 0.02fF
C4720 AND2X1_LOC_824/B OR2X1_LOC_46/A 0.10fF
C4721 OR2X1_LOC_275/A AND2X1_LOC_264/a_36_24# 0.00fF
C4722 AND2X1_LOC_70/Y OR2X1_LOC_374/Y 0.56fF
C4723 OR2X1_LOC_253/a_8_216# OR2X1_LOC_36/Y 0.01fF
C4724 OR2X1_LOC_791/B OR2X1_LOC_287/a_8_216# 0.48fF
C4725 OR2X1_LOC_623/a_36_216# OR2X1_LOC_532/B 0.00fF
C4726 OR2X1_LOC_403/B AND2X1_LOC_51/Y 0.00fF
C4727 OR2X1_LOC_305/Y AND2X1_LOC_307/Y 0.91fF
C4728 OR2X1_LOC_805/A OR2X1_LOC_814/A 0.10fF
C4729 OR2X1_LOC_36/Y OR2X1_LOC_19/B 0.08fF
C4730 OR2X1_LOC_85/A OR2X1_LOC_46/A 1.17fF
C4731 OR2X1_LOC_154/A OR2X1_LOC_62/B 0.08fF
C4732 OR2X1_LOC_43/A OR2X1_LOC_684/Y 0.01fF
C4733 OR2X1_LOC_618/Y AND2X1_LOC_852/B 0.34fF
C4734 AND2X1_LOC_553/A OR2X1_LOC_47/Y 0.33fF
C4735 OR2X1_LOC_617/a_8_216# OR2X1_LOC_617/Y 0.01fF
C4736 OR2X1_LOC_287/B OR2X1_LOC_401/B 0.01fF
C4737 OR2X1_LOC_223/A OR2X1_LOC_794/A 0.02fF
C4738 OR2X1_LOC_62/B OR2X1_LOC_267/A 0.04fF
C4739 OR2X1_LOC_223/B AND2X1_LOC_47/Y 0.00fF
C4740 OR2X1_LOC_160/A OR2X1_LOC_201/a_8_216# 0.01fF
C4741 AND2X1_LOC_34/a_8_24# OR2X1_LOC_416/Y 0.01fF
C4742 AND2X1_LOC_866/A OR2X1_LOC_39/A 0.07fF
C4743 OR2X1_LOC_22/Y AND2X1_LOC_857/a_8_24# 0.00fF
C4744 OR2X1_LOC_19/B AND2X1_LOC_822/a_8_24# 0.02fF
C4745 OR2X1_LOC_18/Y GATE_662 0.02fF
C4746 AND2X1_LOC_393/a_8_24# OR2X1_LOC_532/B 0.01fF
C4747 OR2X1_LOC_779/Y OR2X1_LOC_784/Y 0.11fF
C4748 OR2X1_LOC_22/Y OR2X1_LOC_7/A 0.62fF
C4749 AND2X1_LOC_227/Y OR2X1_LOC_85/A 0.05fF
C4750 OR2X1_LOC_769/B AND2X1_LOC_31/Y 0.05fF
C4751 AND2X1_LOC_270/a_8_24# OR2X1_LOC_6/A 0.01fF
C4752 OR2X1_LOC_31/Y OR2X1_LOC_44/Y 2.63fF
C4753 OR2X1_LOC_537/a_36_216# OR2X1_LOC_390/A 0.00fF
C4754 AND2X1_LOC_486/Y AND2X1_LOC_405/a_8_24# 0.06fF
C4755 AND2X1_LOC_583/a_8_24# AND2X1_LOC_31/Y 0.01fF
C4756 OR2X1_LOC_112/B OR2X1_LOC_539/Y 0.02fF
C4757 OR2X1_LOC_639/A AND2X1_LOC_51/Y 0.01fF
C4758 AND2X1_LOC_76/Y AND2X1_LOC_203/Y 0.03fF
C4759 AND2X1_LOC_91/B OR2X1_LOC_115/B 0.34fF
C4760 AND2X1_LOC_64/Y OR2X1_LOC_554/a_8_216# 0.05fF
C4761 OR2X1_LOC_85/a_8_216# OR2X1_LOC_278/Y 0.01fF
C4762 OR2X1_LOC_62/B OR2X1_LOC_204/a_36_216# 0.00fF
C4763 OR2X1_LOC_629/B OR2X1_LOC_777/B 0.01fF
C4764 OR2X1_LOC_599/A OR2X1_LOC_760/a_8_216# 0.00fF
C4765 AND2X1_LOC_856/B AND2X1_LOC_856/a_8_24# 0.01fF
C4766 OR2X1_LOC_160/A OR2X1_LOC_796/B 0.01fF
C4767 OR2X1_LOC_620/Y OR2X1_LOC_365/B 0.00fF
C4768 OR2X1_LOC_121/B OR2X1_LOC_99/B 0.02fF
C4769 OR2X1_LOC_62/B OR2X1_LOC_778/A 0.00fF
C4770 AND2X1_LOC_817/B D_INPUT_1 0.26fF
C4771 AND2X1_LOC_12/Y AND2X1_LOC_225/a_8_24# 0.01fF
C4772 OR2X1_LOC_186/Y OR2X1_LOC_319/Y 0.02fF
C4773 AND2X1_LOC_856/a_8_24# AND2X1_LOC_863/A 0.02fF
C4774 AND2X1_LOC_12/Y OR2X1_LOC_194/a_8_216# 0.01fF
C4775 OR2X1_LOC_131/Y OR2X1_LOC_71/Y 0.43fF
C4776 OR2X1_LOC_161/A OR2X1_LOC_493/Y 0.01fF
C4777 OR2X1_LOC_47/Y OR2X1_LOC_248/a_8_216# 0.08fF
C4778 OR2X1_LOC_363/B OR2X1_LOC_580/A 0.01fF
C4779 AND2X1_LOC_211/B AND2X1_LOC_866/A 0.07fF
C4780 AND2X1_LOC_456/Y OR2X1_LOC_95/Y 0.03fF
C4781 AND2X1_LOC_852/a_8_24# D_INPUT_1 0.01fF
C4782 OR2X1_LOC_726/A OR2X1_LOC_726/a_36_216# 0.00fF
C4783 OR2X1_LOC_851/A OR2X1_LOC_228/Y 0.02fF
C4784 OR2X1_LOC_490/Y OR2X1_LOC_95/Y 0.07fF
C4785 OR2X1_LOC_74/A OR2X1_LOC_95/Y 0.16fF
C4786 OR2X1_LOC_436/a_8_216# OR2X1_LOC_814/A 0.02fF
C4787 OR2X1_LOC_106/Y OR2X1_LOC_428/A 0.02fF
C4788 OR2X1_LOC_74/A AND2X1_LOC_440/a_8_24# 0.01fF
C4789 OR2X1_LOC_280/Y OR2X1_LOC_224/a_8_216# 0.03fF
C4790 OR2X1_LOC_813/Y OR2X1_LOC_85/A 0.10fF
C4791 OR2X1_LOC_641/Y OR2X1_LOC_771/B 0.10fF
C4792 AND2X1_LOC_95/Y OR2X1_LOC_552/A 0.03fF
C4793 OR2X1_LOC_597/a_8_216# OR2X1_LOC_13/B 0.02fF
C4794 OR2X1_LOC_405/Y OR2X1_LOC_358/A 0.09fF
C4795 OR2X1_LOC_675/a_8_216# OR2X1_LOC_440/A 0.07fF
C4796 OR2X1_LOC_47/Y AND2X1_LOC_294/a_8_24# 0.02fF
C4797 AND2X1_LOC_564/B AND2X1_LOC_785/Y 0.01fF
C4798 OR2X1_LOC_631/B OR2X1_LOC_247/a_8_216# 0.06fF
C4799 OR2X1_LOC_680/Y AND2X1_LOC_796/Y -0.00fF
C4800 OR2X1_LOC_106/Y OR2X1_LOC_595/A 0.09fF
C4801 OR2X1_LOC_781/Y OR2X1_LOC_782/a_8_216# 0.02fF
C4802 OR2X1_LOC_756/B OR2X1_LOC_580/A 0.25fF
C4803 OR2X1_LOC_66/A OR2X1_LOC_308/Y 0.07fF
C4804 OR2X1_LOC_95/Y OR2X1_LOC_261/A 0.01fF
C4805 AND2X1_LOC_580/B AND2X1_LOC_805/a_8_24# 0.01fF
C4806 AND2X1_LOC_572/Y AND2X1_LOC_563/Y 0.54fF
C4807 AND2X1_LOC_95/Y OR2X1_LOC_578/B 8.49fF
C4808 AND2X1_LOC_44/Y OR2X1_LOC_342/A 0.01fF
C4809 OR2X1_LOC_748/A AND2X1_LOC_848/A 0.04fF
C4810 OR2X1_LOC_87/A AND2X1_LOC_52/Y 0.22fF
C4811 AND2X1_LOC_832/a_8_24# OR2X1_LOC_423/Y 0.04fF
C4812 OR2X1_LOC_685/A AND2X1_LOC_430/B 0.00fF
C4813 OR2X1_LOC_256/Y AND2X1_LOC_247/a_8_24# 0.01fF
C4814 OR2X1_LOC_64/Y AND2X1_LOC_318/Y 0.05fF
C4815 AND2X1_LOC_828/a_8_24# OR2X1_LOC_12/Y 0.01fF
C4816 OR2X1_LOC_578/a_36_216# OR2X1_LOC_549/A 0.00fF
C4817 AND2X1_LOC_719/Y AND2X1_LOC_244/A 0.05fF
C4818 AND2X1_LOC_99/A OR2X1_LOC_13/B 0.01fF
C4819 AND2X1_LOC_500/B OR2X1_LOC_530/a_8_216# 0.18fF
C4820 OR2X1_LOC_49/A OR2X1_LOC_9/Y 0.06fF
C4821 AND2X1_LOC_287/B AND2X1_LOC_860/A 0.01fF
C4822 AND2X1_LOC_141/a_8_24# AND2X1_LOC_772/Y 0.02fF
C4823 AND2X1_LOC_645/A OR2X1_LOC_331/Y 0.26fF
C4824 OR2X1_LOC_134/Y AND2X1_LOC_772/B 0.01fF
C4825 AND2X1_LOC_851/B INPUT_1 0.07fF
C4826 OR2X1_LOC_743/A OR2X1_LOC_761/a_8_216# 0.01fF
C4827 AND2X1_LOC_227/Y OR2X1_LOC_226/Y 0.80fF
C4828 OR2X1_LOC_176/a_36_216# AND2X1_LOC_568/B 0.01fF
C4829 OR2X1_LOC_322/Y OR2X1_LOC_323/Y 0.78fF
C4830 AND2X1_LOC_282/a_8_24# OR2X1_LOC_366/Y 0.02fF
C4831 AND2X1_LOC_795/a_8_24# AND2X1_LOC_778/Y 0.19fF
C4832 D_INPUT_3 AND2X1_LOC_839/A 0.00fF
C4833 AND2X1_LOC_70/Y OR2X1_LOC_392/B 0.01fF
C4834 OR2X1_LOC_62/B OR2X1_LOC_84/a_8_216# 0.01fF
C4835 OR2X1_LOC_502/A AND2X1_LOC_762/a_8_24# 0.01fF
C4836 AND2X1_LOC_215/Y AND2X1_LOC_219/A 0.00fF
C4837 OR2X1_LOC_808/A OR2X1_LOC_718/a_8_216# 0.04fF
C4838 OR2X1_LOC_135/a_8_216# VDD 0.21fF
C4839 AND2X1_LOC_831/Y AND2X1_LOC_660/A 0.04fF
C4840 OR2X1_LOC_715/B OR2X1_LOC_151/A 0.10fF
C4841 OR2X1_LOC_405/A AND2X1_LOC_36/Y 0.07fF
C4842 AND2X1_LOC_7/B OR2X1_LOC_715/A 0.02fF
C4843 OR2X1_LOC_624/A AND2X1_LOC_239/a_8_24# 0.25fF
C4844 AND2X1_LOC_47/Y OR2X1_LOC_845/A 0.21fF
C4845 OR2X1_LOC_364/A OR2X1_LOC_788/B 0.07fF
C4846 OR2X1_LOC_45/B OR2X1_LOC_744/A 1.58fF
C4847 OR2X1_LOC_574/a_8_216# OR2X1_LOC_140/B 0.01fF
C4848 AND2X1_LOC_521/a_8_24# VDD 0.00fF
C4849 OR2X1_LOC_437/a_8_216# AND2X1_LOC_675/A 0.07fF
C4850 OR2X1_LOC_185/Y AND2X1_LOC_41/Y 0.00fF
C4851 AND2X1_LOC_91/B OR2X1_LOC_840/A 0.10fF
C4852 AND2X1_LOC_719/Y OR2X1_LOC_108/Y 0.10fF
C4853 VDD OR2X1_LOC_646/B 0.02fF
C4854 INPUT_1 OR2X1_LOC_595/Y 0.11fF
C4855 AND2X1_LOC_22/Y OR2X1_LOC_663/A 0.07fF
C4856 OR2X1_LOC_52/B OR2X1_LOC_424/Y -0.01fF
C4857 OR2X1_LOC_863/A OR2X1_LOC_35/Y 0.01fF
C4858 AND2X1_LOC_471/Y AND2X1_LOC_786/Y 0.01fF
C4859 OR2X1_LOC_756/B AND2X1_LOC_44/Y 0.07fF
C4860 OR2X1_LOC_329/B AND2X1_LOC_810/B 1.53fF
C4861 OR2X1_LOC_47/Y AND2X1_LOC_648/B 0.03fF
C4862 OR2X1_LOC_494/Y AND2X1_LOC_243/Y 0.07fF
C4863 D_INPUT_0 OR2X1_LOC_358/A 0.07fF
C4864 AND2X1_LOC_47/Y OR2X1_LOC_551/A 0.01fF
C4865 INPUT_0 OR2X1_LOC_829/A 0.10fF
C4866 OR2X1_LOC_175/Y OR2X1_LOC_175/B 0.09fF
C4867 AND2X1_LOC_392/A AND2X1_LOC_335/Y 0.01fF
C4868 AND2X1_LOC_181/Y OR2X1_LOC_329/B 0.01fF
C4869 OR2X1_LOC_147/B AND2X1_LOC_7/B 0.03fF
C4870 AND2X1_LOC_477/A OR2X1_LOC_331/Y 0.07fF
C4871 OR2X1_LOC_62/B OR2X1_LOC_560/A 0.02fF
C4872 OR2X1_LOC_776/Y OR2X1_LOC_785/a_8_216# 0.02fF
C4873 OR2X1_LOC_348/Y OR2X1_LOC_287/A 0.08fF
C4874 OR2X1_LOC_165/a_36_216# AND2X1_LOC_787/A 0.00fF
C4875 OR2X1_LOC_696/A AND2X1_LOC_818/a_8_24# 0.06fF
C4876 OR2X1_LOC_71/Y AND2X1_LOC_657/A 0.28fF
C4877 OR2X1_LOC_602/Y AND2X1_LOC_92/Y 0.42fF
C4878 AND2X1_LOC_43/B OR2X1_LOC_563/A 0.00fF
C4879 OR2X1_LOC_97/A OR2X1_LOC_624/A 0.03fF
C4880 OR2X1_LOC_323/A OR2X1_LOC_36/Y 0.04fF
C4881 AND2X1_LOC_293/a_8_24# OR2X1_LOC_68/B -0.01fF
C4882 AND2X1_LOC_847/Y OR2X1_LOC_428/A 0.01fF
C4883 OR2X1_LOC_660/B AND2X1_LOC_44/Y 0.03fF
C4884 AND2X1_LOC_541/Y OR2X1_LOC_103/Y 0.19fF
C4885 OR2X1_LOC_148/a_36_216# OR2X1_LOC_161/A 0.00fF
C4886 AND2X1_LOC_452/Y OR2X1_LOC_12/Y 0.01fF
C4887 OR2X1_LOC_773/Y OR2X1_LOC_269/B 0.01fF
C4888 AND2X1_LOC_858/B OR2X1_LOC_59/Y 0.10fF
C4889 OR2X1_LOC_448/Y OR2X1_LOC_161/B 0.02fF
C4890 OR2X1_LOC_506/A AND2X1_LOC_433/a_36_24# 0.00fF
C4891 AND2X1_LOC_656/a_36_24# OR2X1_LOC_595/A 0.01fF
C4892 OR2X1_LOC_364/A AND2X1_LOC_22/Y 0.07fF
C4893 OR2X1_LOC_313/Y OR2X1_LOC_16/A 0.08fF
C4894 OR2X1_LOC_91/A OR2X1_LOC_59/Y 0.08fF
C4895 OR2X1_LOC_185/Y AND2X1_LOC_22/Y 5.21fF
C4896 OR2X1_LOC_116/a_8_216# OR2X1_LOC_392/B 0.12fF
C4897 VDD OR2X1_LOC_828/a_8_216# 0.21fF
C4898 OR2X1_LOC_148/Y OR2X1_LOC_161/A 0.01fF
C4899 AND2X1_LOC_655/A OR2X1_LOC_16/A 0.11fF
C4900 AND2X1_LOC_513/a_8_24# OR2X1_LOC_51/Y 0.08fF
C4901 AND2X1_LOC_88/Y OR2X1_LOC_560/A 0.01fF
C4902 OR2X1_LOC_45/B AND2X1_LOC_840/B 0.03fF
C4903 OR2X1_LOC_87/A OR2X1_LOC_576/A 0.94fF
C4904 OR2X1_LOC_49/A OR2X1_LOC_96/B 0.21fF
C4905 OR2X1_LOC_130/A OR2X1_LOC_435/A 0.02fF
C4906 AND2X1_LOC_40/Y AND2X1_LOC_616/a_8_24# 0.01fF
C4907 AND2X1_LOC_125/a_8_24# OR2X1_LOC_66/A 0.02fF
C4908 AND2X1_LOC_464/A OR2X1_LOC_44/Y 0.05fF
C4909 AND2X1_LOC_729/Y OR2X1_LOC_589/A 0.03fF
C4910 AND2X1_LOC_213/B OR2X1_LOC_44/Y 0.02fF
C4911 AND2X1_LOC_707/Y OR2X1_LOC_52/B 0.03fF
C4912 OR2X1_LOC_604/A OR2X1_LOC_278/Y 0.05fF
C4913 OR2X1_LOC_158/A OR2X1_LOC_316/Y 0.04fF
C4914 AND2X1_LOC_572/a_8_24# OR2X1_LOC_89/A 0.01fF
C4915 AND2X1_LOC_784/A AND2X1_LOC_364/a_8_24# 0.01fF
C4916 AND2X1_LOC_64/Y AND2X1_LOC_69/Y 0.01fF
C4917 OR2X1_LOC_107/a_8_216# OR2X1_LOC_103/Y 0.01fF
C4918 OR2X1_LOC_49/A AND2X1_LOC_852/Y 0.03fF
C4919 AND2X1_LOC_191/Y AND2X1_LOC_192/a_36_24# 0.01fF
C4920 AND2X1_LOC_392/A OR2X1_LOC_619/Y 3.24fF
C4921 OR2X1_LOC_427/A AND2X1_LOC_285/Y 0.02fF
C4922 AND2X1_LOC_552/a_8_24# AND2X1_LOC_578/A 0.02fF
C4923 OR2X1_LOC_24/Y AND2X1_LOC_208/Y 0.80fF
C4924 OR2X1_LOC_653/a_8_216# OR2X1_LOC_392/B 0.40fF
C4925 OR2X1_LOC_40/Y OR2X1_LOC_39/A 0.18fF
C4926 VDD OR2X1_LOC_506/A 0.85fF
C4927 OR2X1_LOC_87/A OR2X1_LOC_439/B 0.03fF
C4928 AND2X1_LOC_22/Y AND2X1_LOC_171/a_36_24# 0.00fF
C4929 OR2X1_LOC_114/B OR2X1_LOC_128/a_8_216# 0.01fF
C4930 OR2X1_LOC_158/A AND2X1_LOC_354/B 0.11fF
C4931 OR2X1_LOC_528/Y AND2X1_LOC_186/a_36_24# 0.01fF
C4932 VDD AND2X1_LOC_695/a_8_24# -0.00fF
C4933 OR2X1_LOC_609/A OR2X1_LOC_16/A 0.48fF
C4934 OR2X1_LOC_19/B OR2X1_LOC_19/a_8_216# 0.09fF
C4935 VDD AND2X1_LOC_129/a_8_24# -0.00fF
C4936 OR2X1_LOC_39/Y OR2X1_LOC_16/Y 0.05fF
C4937 OR2X1_LOC_520/Y AND2X1_LOC_18/Y 0.03fF
C4938 OR2X1_LOC_85/A INPUT_2 0.02fF
C4939 OR2X1_LOC_404/Y OR2X1_LOC_392/B 0.05fF
C4940 AND2X1_LOC_365/a_8_24# AND2X1_LOC_841/B 0.07fF
C4941 AND2X1_LOC_154/a_8_24# AND2X1_LOC_658/A 0.03fF
C4942 OR2X1_LOC_160/B OR2X1_LOC_687/Y 0.07fF
C4943 OR2X1_LOC_805/A OR2X1_LOC_244/Y 0.03fF
C4944 AND2X1_LOC_573/A OR2X1_LOC_59/Y 0.03fF
C4945 OR2X1_LOC_223/A OR2X1_LOC_716/a_36_216# 0.00fF
C4946 AND2X1_LOC_390/a_8_24# OR2X1_LOC_43/A 0.01fF
C4947 AND2X1_LOC_724/a_8_24# OR2X1_LOC_417/Y 0.07fF
C4948 OR2X1_LOC_496/Y AND2X1_LOC_778/Y 0.01fF
C4949 OR2X1_LOC_821/Y OR2X1_LOC_74/A 0.01fF
C4950 OR2X1_LOC_6/B OR2X1_LOC_6/a_8_216# 0.08fF
C4951 OR2X1_LOC_502/A OR2X1_LOC_623/B 0.01fF
C4952 OR2X1_LOC_599/A OR2X1_LOC_536/Y 0.01fF
C4953 OR2X1_LOC_744/A AND2X1_LOC_435/a_8_24# 0.01fF
C4954 AND2X1_LOC_70/Y OR2X1_LOC_685/A 0.01fF
C4955 OR2X1_LOC_86/a_36_216# AND2X1_LOC_243/Y 0.01fF
C4956 AND2X1_LOC_12/Y INPUT_0 0.04fF
C4957 INPUT_3 AND2X1_LOC_54/a_8_24# 0.01fF
C4958 OR2X1_LOC_650/a_8_216# OR2X1_LOC_462/B 0.01fF
C4959 OR2X1_LOC_641/Y OR2X1_LOC_642/a_8_216# 0.03fF
C4960 OR2X1_LOC_441/Y AND2X1_LOC_811/B 0.06fF
C4961 OR2X1_LOC_136/Y OR2X1_LOC_46/A 0.00fF
C4962 OR2X1_LOC_40/Y AND2X1_LOC_211/B 0.53fF
C4963 AND2X1_LOC_675/Y AND2X1_LOC_186/a_8_24# 0.08fF
C4964 OR2X1_LOC_158/A OR2X1_LOC_824/a_8_216# 0.14fF
C4965 INPUT_0 AND2X1_LOC_838/Y 0.16fF
C4966 OR2X1_LOC_158/A AND2X1_LOC_390/B 0.07fF
C4967 AND2X1_LOC_354/a_8_24# OR2X1_LOC_329/B 0.06fF
C4968 AND2X1_LOC_56/B OR2X1_LOC_35/Y 0.04fF
C4969 AND2X1_LOC_576/Y AND2X1_LOC_561/B 0.84fF
C4970 AND2X1_LOC_633/Y AND2X1_LOC_202/Y 0.16fF
C4971 AND2X1_LOC_117/a_8_24# OR2X1_LOC_549/A 0.03fF
C4972 OR2X1_LOC_329/Y OR2X1_LOC_485/A 0.01fF
C4973 AND2X1_LOC_95/Y OR2X1_LOC_798/Y 0.09fF
C4974 AND2X1_LOC_715/Y OR2X1_LOC_601/a_36_216# 0.01fF
C4975 AND2X1_LOC_95/Y AND2X1_LOC_52/a_8_24# 0.08fF
C4976 OR2X1_LOC_485/A AND2X1_LOC_606/a_8_24# 0.03fF
C4977 OR2X1_LOC_529/a_8_216# OR2X1_LOC_103/Y 0.01fF
C4978 OR2X1_LOC_181/B OR2X1_LOC_540/a_8_216# 0.02fF
C4979 OR2X1_LOC_593/A OR2X1_LOC_66/A 0.01fF
C4980 OR2X1_LOC_545/B AND2X1_LOC_7/B 0.03fF
C4981 OR2X1_LOC_64/Y OR2X1_LOC_829/A 0.01fF
C4982 OR2X1_LOC_134/a_36_216# AND2X1_LOC_227/Y 0.00fF
C4983 OR2X1_LOC_70/Y OR2X1_LOC_131/a_8_216# 0.15fF
C4984 OR2X1_LOC_404/Y OR2X1_LOC_113/B 0.00fF
C4985 OR2X1_LOC_624/A OR2X1_LOC_475/B 0.03fF
C4986 OR2X1_LOC_51/Y OR2X1_LOC_106/A 0.01fF
C4987 AND2X1_LOC_810/A AND2X1_LOC_727/A 3.08fF
C4988 AND2X1_LOC_513/a_8_24# OR2X1_LOC_680/A -0.06fF
C4989 OR2X1_LOC_154/A OR2X1_LOC_659/A 0.19fF
C4990 AND2X1_LOC_580/A AND2X1_LOC_508/A 0.03fF
C4991 AND2X1_LOC_41/A OR2X1_LOC_87/A 0.23fF
C4992 OR2X1_LOC_467/A OR2X1_LOC_453/A 0.01fF
C4993 OR2X1_LOC_656/B OR2X1_LOC_327/a_8_216# 0.01fF
C4994 AND2X1_LOC_12/Y OR2X1_LOC_772/B 0.60fF
C4995 OR2X1_LOC_865/a_8_216# OR2X1_LOC_859/a_8_216# 0.47fF
C4996 OR2X1_LOC_91/A OR2X1_LOC_820/B 0.61fF
C4997 AND2X1_LOC_91/B OR2X1_LOC_241/Y 0.10fF
C4998 AND2X1_LOC_64/Y OR2X1_LOC_506/B 0.15fF
C4999 OR2X1_LOC_669/Y OR2X1_LOC_59/Y 0.82fF
C5000 AND2X1_LOC_705/a_36_24# OR2X1_LOC_485/A 0.00fF
C5001 OR2X1_LOC_329/B OR2X1_LOC_585/A 0.21fF
C5002 AND2X1_LOC_332/a_8_24# OR2X1_LOC_46/A 0.07fF
C5003 OR2X1_LOC_358/A OR2X1_LOC_339/A 0.72fF
C5004 OR2X1_LOC_185/A AND2X1_LOC_74/a_36_24# 0.01fF
C5005 OR2X1_LOC_92/Y OR2X1_LOC_67/a_8_216# 0.05fF
C5006 OR2X1_LOC_742/B OR2X1_LOC_550/B 0.33fF
C5007 AND2X1_LOC_354/Y AND2X1_LOC_356/a_8_24# 0.10fF
C5008 AND2X1_LOC_376/a_8_24# INPUT_0 0.01fF
C5009 OR2X1_LOC_629/A OR2X1_LOC_78/A 0.01fF
C5010 VDD OR2X1_LOC_481/A 0.36fF
C5011 OR2X1_LOC_508/A OR2X1_LOC_87/A 0.07fF
C5012 OR2X1_LOC_45/B OR2X1_LOC_31/Y 0.59fF
C5013 OR2X1_LOC_260/Y OR2X1_LOC_555/B 0.02fF
C5014 OR2X1_LOC_756/B OR2X1_LOC_465/B 0.06fF
C5015 OR2X1_LOC_446/B AND2X1_LOC_419/a_8_24# 0.01fF
C5016 OR2X1_LOC_568/A OR2X1_LOC_788/B 0.13fF
C5017 AND2X1_LOC_724/A OR2X1_LOC_167/Y 0.05fF
C5018 OR2X1_LOC_377/A OR2X1_LOC_240/a_8_216# 0.01fF
C5019 OR2X1_LOC_604/A OR2X1_LOC_253/a_8_216# 0.03fF
C5020 OR2X1_LOC_47/Y AND2X1_LOC_465/A 0.02fF
C5021 AND2X1_LOC_605/Y AND2X1_LOC_645/A 0.00fF
C5022 AND2X1_LOC_31/Y OR2X1_LOC_712/B 0.03fF
C5023 OR2X1_LOC_91/Y OR2X1_LOC_427/A 0.10fF
C5024 AND2X1_LOC_597/a_36_24# AND2X1_LOC_40/Y 0.00fF
C5025 OR2X1_LOC_808/a_36_216# OR2X1_LOC_87/A 0.00fF
C5026 AND2X1_LOC_12/Y OR2X1_LOC_489/B 0.00fF
C5027 AND2X1_LOC_476/A AND2X1_LOC_476/a_36_24# 0.00fF
C5028 OR2X1_LOC_154/A OR2X1_LOC_724/a_36_216# 0.00fF
C5029 OR2X1_LOC_451/B AND2X1_LOC_581/a_36_24# 0.00fF
C5030 OR2X1_LOC_160/B OR2X1_LOC_643/Y 0.02fF
C5031 OR2X1_LOC_648/B OR2X1_LOC_814/A 0.16fF
C5032 OR2X1_LOC_502/A OR2X1_LOC_585/A 0.03fF
C5033 AND2X1_LOC_721/a_8_24# OR2X1_LOC_251/Y 0.01fF
C5034 OR2X1_LOC_70/Y OR2X1_LOC_91/A 0.69fF
C5035 OR2X1_LOC_19/B OR2X1_LOC_66/A 0.86fF
C5036 AND2X1_LOC_580/A OR2X1_LOC_18/Y 0.03fF
C5037 AND2X1_LOC_107/a_8_24# AND2X1_LOC_18/Y 0.02fF
C5038 AND2X1_LOC_59/Y OR2X1_LOC_350/a_8_216# 0.01fF
C5039 OR2X1_LOC_625/Y OR2X1_LOC_248/a_8_216# -0.00fF
C5040 AND2X1_LOC_347/Y OR2X1_LOC_3/Y 0.00fF
C5041 OR2X1_LOC_158/A AND2X1_LOC_863/Y 0.07fF
C5042 AND2X1_LOC_64/Y OR2X1_LOC_247/Y 0.01fF
C5043 OR2X1_LOC_845/A AND2X1_LOC_263/a_36_24# 0.01fF
C5044 OR2X1_LOC_620/Y OR2X1_LOC_449/B 0.07fF
C5045 OR2X1_LOC_3/Y AND2X1_LOC_857/Y 0.03fF
C5046 OR2X1_LOC_502/A AND2X1_LOC_43/a_8_24# 0.01fF
C5047 AND2X1_LOC_144/a_8_24# AND2X1_LOC_51/Y 0.01fF
C5048 OR2X1_LOC_427/A AND2X1_LOC_446/a_8_24# 0.01fF
C5049 OR2X1_LOC_599/A AND2X1_LOC_593/Y 0.04fF
C5050 OR2X1_LOC_662/A OR2X1_LOC_87/A 0.28fF
C5051 OR2X1_LOC_51/Y OR2X1_LOC_46/A 0.01fF
C5052 AND2X1_LOC_486/Y OR2X1_LOC_529/Y 0.03fF
C5053 OR2X1_LOC_426/B AND2X1_LOC_326/a_8_24# 0.03fF
C5054 OR2X1_LOC_189/Y OR2X1_LOC_427/A 0.03fF
C5055 AND2X1_LOC_779/a_8_24# OR2X1_LOC_89/A 0.01fF
C5056 OR2X1_LOC_377/A OR2X1_LOC_269/B 1.58fF
C5057 AND2X1_LOC_1/Y AND2X1_LOC_12/a_8_24# 0.09fF
C5058 AND2X1_LOC_514/Y OR2X1_LOC_91/A 0.02fF
C5059 OR2X1_LOC_81/Y OR2X1_LOC_69/A 0.01fF
C5060 OR2X1_LOC_625/Y AND2X1_LOC_294/a_8_24# 0.02fF
C5061 VDD OR2X1_LOC_71/Y 0.53fF
C5062 AND2X1_LOC_729/Y OR2X1_LOC_43/A 0.04fF
C5063 OR2X1_LOC_759/A OR2X1_LOC_417/A 0.02fF
C5064 AND2X1_LOC_165/a_8_24# OR2X1_LOC_78/A 0.03fF
C5065 VDD OR2X1_LOC_780/A 0.21fF
C5066 AND2X1_LOC_95/Y OR2X1_LOC_654/A 0.03fF
C5067 AND2X1_LOC_303/B OR2X1_LOC_6/A 1.52fF
C5068 AND2X1_LOC_70/Y OR2X1_LOC_532/B 2.58fF
C5069 AND2X1_LOC_578/A AND2X1_LOC_840/A 0.03fF
C5070 AND2X1_LOC_7/B OR2X1_LOC_318/B 0.00fF
C5071 AND2X1_LOC_40/Y OR2X1_LOC_285/B 0.17fF
C5072 OR2X1_LOC_599/Y OR2X1_LOC_16/A 0.04fF
C5073 AND2X1_LOC_705/a_8_24# OR2X1_LOC_31/Y 0.07fF
C5074 OR2X1_LOC_95/Y OR2X1_LOC_626/Y 0.06fF
C5075 AND2X1_LOC_716/Y AND2X1_LOC_326/A 0.00fF
C5076 OR2X1_LOC_154/A OR2X1_LOC_449/B 0.07fF
C5077 OR2X1_LOC_375/A OR2X1_LOC_552/a_36_216# 0.00fF
C5078 OR2X1_LOC_7/A OR2X1_LOC_39/A 0.13fF
C5079 OR2X1_LOC_574/A OR2X1_LOC_539/Y 0.15fF
C5080 AND2X1_LOC_86/B AND2X1_LOC_617/a_8_24# 0.03fF
C5081 OR2X1_LOC_169/a_8_216# OR2X1_LOC_778/Y 0.35fF
C5082 AND2X1_LOC_59/Y AND2X1_LOC_3/Y 0.09fF
C5083 OR2X1_LOC_85/A AND2X1_LOC_267/a_36_24# 0.00fF
C5084 OR2X1_LOC_446/Y OR2X1_LOC_78/A 0.01fF
C5085 AND2X1_LOC_605/Y AND2X1_LOC_477/A 0.03fF
C5086 AND2X1_LOC_326/B AND2X1_LOC_841/a_8_24# 0.01fF
C5087 OR2X1_LOC_504/Y AND2X1_LOC_858/B 0.01fF
C5088 OR2X1_LOC_468/Y OR2X1_LOC_778/Y 0.05fF
C5089 AND2X1_LOC_784/A OR2X1_LOC_43/A 0.07fF
C5090 OR2X1_LOC_659/B OR2X1_LOC_720/a_8_216# 0.14fF
C5091 AND2X1_LOC_326/A AND2X1_LOC_654/Y 0.01fF
C5092 AND2X1_LOC_41/A OR2X1_LOC_706/B 0.04fF
C5093 AND2X1_LOC_287/B AND2X1_LOC_562/Y 0.11fF
C5094 OR2X1_LOC_624/B AND2X1_LOC_617/a_8_24# 0.01fF
C5095 VDD OR2X1_LOC_227/Y 0.19fF
C5096 AND2X1_LOC_537/Y OR2X1_LOC_92/Y 0.01fF
C5097 OR2X1_LOC_70/Y AND2X1_LOC_573/A 0.04fF
C5098 OR2X1_LOC_139/A AND2X1_LOC_31/Y 0.03fF
C5099 OR2X1_LOC_160/B OR2X1_LOC_786/Y 0.03fF
C5100 OR2X1_LOC_816/A AND2X1_LOC_562/Y 0.10fF
C5101 OR2X1_LOC_417/Y OR2X1_LOC_427/A 0.04fF
C5102 AND2X1_LOC_48/A OR2X1_LOC_623/B 0.03fF
C5103 OR2X1_LOC_620/Y OR2X1_LOC_121/B 0.02fF
C5104 VDD D_INPUT_1 1.93fF
C5105 OR2X1_LOC_311/Y OR2X1_LOC_427/A 0.03fF
C5106 OR2X1_LOC_161/B AND2X1_LOC_257/a_8_24# 0.00fF
C5107 AND2X1_LOC_474/A AND2X1_LOC_866/A 0.03fF
C5108 OR2X1_LOC_311/Y AND2X1_LOC_801/a_8_24# 0.01fF
C5109 AND2X1_LOC_78/a_8_24# OR2X1_LOC_36/Y 0.01fF
C5110 OR2X1_LOC_753/A AND2X1_LOC_240/Y 0.01fF
C5111 OR2X1_LOC_185/A OR2X1_LOC_476/B 0.00fF
C5112 AND2X1_LOC_211/B AND2X1_LOC_857/a_8_24# 0.01fF
C5113 OR2X1_LOC_473/A OR2X1_LOC_78/A 0.10fF
C5114 OR2X1_LOC_682/a_8_216# OR2X1_LOC_743/A 0.01fF
C5115 AND2X1_LOC_642/a_8_24# OR2X1_LOC_46/A 0.02fF
C5116 OR2X1_LOC_837/B INPUT_1 0.03fF
C5117 OR2X1_LOC_754/A OR2X1_LOC_36/Y 0.14fF
C5118 VDD OR2X1_LOC_173/a_8_216# 0.21fF
C5119 OR2X1_LOC_357/B OR2X1_LOC_357/A 0.15fF
C5120 AND2X1_LOC_211/B OR2X1_LOC_7/A 0.07fF
C5121 OR2X1_LOC_275/A OR2X1_LOC_36/Y 0.02fF
C5122 OR2X1_LOC_849/A OR2X1_LOC_624/B 0.00fF
C5123 D_INPUT_3 AND2X1_LOC_820/B 0.03fF
C5124 AND2X1_LOC_858/B OR2X1_LOC_184/Y 0.08fF
C5125 AND2X1_LOC_177/a_36_24# OR2X1_LOC_440/A 0.00fF
C5126 OR2X1_LOC_158/A OR2X1_LOC_153/a_8_216# 0.01fF
C5127 OR2X1_LOC_154/A OR2X1_LOC_121/B 0.14fF
C5128 AND2X1_LOC_328/a_8_24# AND2X1_LOC_47/Y 0.01fF
C5129 OR2X1_LOC_835/a_8_216# AND2X1_LOC_51/Y 0.01fF
C5130 OR2X1_LOC_401/Y OR2X1_LOC_557/A 0.01fF
C5131 AND2X1_LOC_573/A AND2X1_LOC_657/a_8_24# 0.01fF
C5132 OR2X1_LOC_375/A OR2X1_LOC_46/A 0.07fF
C5133 OR2X1_LOC_223/A OR2X1_LOC_776/a_8_216# 0.01fF
C5134 AND2X1_LOC_240/Y AND2X1_LOC_243/a_8_24# 0.11fF
C5135 AND2X1_LOC_56/B OR2X1_LOC_416/Y 0.16fF
C5136 AND2X1_LOC_640/Y AND2X1_LOC_641/Y 0.23fF
C5137 AND2X1_LOC_34/Y D_INPUT_0 0.00fF
C5138 OR2X1_LOC_699/a_8_216# OR2X1_LOC_54/Y 0.03fF
C5139 OR2X1_LOC_521/Y AND2X1_LOC_851/B 0.01fF
C5140 OR2X1_LOC_791/B OR2X1_LOC_532/B 0.04fF
C5141 D_INPUT_3 OR2X1_LOC_427/A 0.02fF
C5142 OR2X1_LOC_62/B OR2X1_LOC_267/a_8_216# 0.01fF
C5143 OR2X1_LOC_615/a_8_216# OR2X1_LOC_89/A 0.01fF
C5144 OR2X1_LOC_31/Y AND2X1_LOC_435/a_8_24# 0.01fF
C5145 OR2X1_LOC_507/a_8_216# OR2X1_LOC_205/Y 0.05fF
C5146 OR2X1_LOC_791/A OR2X1_LOC_792/A 0.95fF
C5147 OR2X1_LOC_643/Y OR2X1_LOC_219/B 0.00fF
C5148 OR2X1_LOC_18/Y AND2X1_LOC_476/A 0.07fF
C5149 AND2X1_LOC_476/A AND2X1_LOC_649/a_36_24# 0.01fF
C5150 OR2X1_LOC_264/Y OR2X1_LOC_205/Y 0.06fF
C5151 AND2X1_LOC_821/a_8_24# OR2X1_LOC_130/A 0.13fF
C5152 OR2X1_LOC_70/A AND2X1_LOC_637/a_36_24# 0.00fF
C5153 OR2X1_LOC_823/Y D_INPUT_3 0.01fF
C5154 OR2X1_LOC_186/Y OR2X1_LOC_777/B 0.02fF
C5155 OR2X1_LOC_49/A OR2X1_LOC_771/B 0.10fF
C5156 OR2X1_LOC_334/B OR2X1_LOC_598/A 0.42fF
C5157 OR2X1_LOC_22/Y OR2X1_LOC_32/a_8_216# 0.01fF
C5158 AND2X1_LOC_86/Y OR2X1_LOC_786/Y 0.02fF
C5159 OR2X1_LOC_78/A OR2X1_LOC_228/Y 0.07fF
C5160 OR2X1_LOC_78/B OR2X1_LOC_641/B 0.03fF
C5161 AND2X1_LOC_67/Y OR2X1_LOC_202/a_36_216# 0.03fF
C5162 AND2X1_LOC_324/a_8_24# OR2X1_LOC_64/Y 0.01fF
C5163 OR2X1_LOC_184/Y AND2X1_LOC_573/A 0.02fF
C5164 AND2X1_LOC_500/B OR2X1_LOC_437/A 0.01fF
C5165 OR2X1_LOC_637/Y AND2X1_LOC_31/Y 0.02fF
C5166 OR2X1_LOC_427/A AND2X1_LOC_483/Y 0.03fF
C5167 OR2X1_LOC_312/Y OR2X1_LOC_167/Y 0.09fF
C5168 AND2X1_LOC_59/Y OR2X1_LOC_270/Y 0.28fF
C5169 OR2X1_LOC_47/Y OR2X1_LOC_237/Y 0.02fF
C5170 OR2X1_LOC_446/Y OR2X1_LOC_155/A 1.17fF
C5171 AND2X1_LOC_40/Y OR2X1_LOC_358/A 0.00fF
C5172 AND2X1_LOC_489/a_8_24# OR2X1_LOC_437/A 0.02fF
C5173 OR2X1_LOC_319/B OR2X1_LOC_854/A 0.02fF
C5174 OR2X1_LOC_318/Y OR2X1_LOC_318/B 0.00fF
C5175 AND2X1_LOC_192/Y GATE_811 0.09fF
C5176 OR2X1_LOC_458/a_36_216# AND2X1_LOC_31/Y 0.00fF
C5177 OR2X1_LOC_43/A OR2X1_LOC_62/A 0.18fF
C5178 OR2X1_LOC_653/a_8_216# OR2X1_LOC_532/B 0.01fF
C5179 AND2X1_LOC_580/A AND2X1_LOC_620/Y 0.03fF
C5180 OR2X1_LOC_87/A OR2X1_LOC_207/a_8_216# 0.01fF
C5181 OR2X1_LOC_140/B AND2X1_LOC_44/Y 0.01fF
C5182 AND2X1_LOC_224/a_8_24# OR2X1_LOC_227/B 0.02fF
C5183 AND2X1_LOC_654/B OR2X1_LOC_172/Y 0.74fF
C5184 AND2X1_LOC_848/A AND2X1_LOC_848/a_8_24# 0.02fF
C5185 OR2X1_LOC_22/Y AND2X1_LOC_115/a_8_24# -0.01fF
C5186 OR2X1_LOC_643/A OR2X1_LOC_205/Y 0.19fF
C5187 OR2X1_LOC_404/Y OR2X1_LOC_532/B 0.03fF
C5188 AND2X1_LOC_621/Y AND2X1_LOC_222/Y 0.03fF
C5189 OR2X1_LOC_205/Y OR2X1_LOC_124/Y 0.01fF
C5190 OR2X1_LOC_186/Y OR2X1_LOC_566/A 0.02fF
C5191 OR2X1_LOC_323/A OR2X1_LOC_315/a_8_216# 0.00fF
C5192 VDD OR2X1_LOC_180/B 0.09fF
C5193 OR2X1_LOC_45/B OR2X1_LOC_79/a_8_216# 0.02fF
C5194 OR2X1_LOC_840/A OR2X1_LOC_446/B 0.01fF
C5195 OR2X1_LOC_175/Y OR2X1_LOC_389/a_8_216# 0.01fF
C5196 OR2X1_LOC_45/B AND2X1_LOC_464/A 0.00fF
C5197 AND2X1_LOC_100/a_8_24# OR2X1_LOC_86/A 0.05fF
C5198 OR2X1_LOC_121/Y AND2X1_LOC_7/B 0.01fF
C5199 OR2X1_LOC_188/Y OR2X1_LOC_486/Y 0.03fF
C5200 OR2X1_LOC_847/a_8_216# OR2X1_LOC_68/B 0.01fF
C5201 OR2X1_LOC_323/A OR2X1_LOC_604/A 0.03fF
C5202 AND2X1_LOC_43/B OR2X1_LOC_724/A 0.11fF
C5203 OR2X1_LOC_64/Y OR2X1_LOC_224/Y 0.01fF
C5204 AND2X1_LOC_64/Y AND2X1_LOC_18/Y 0.48fF
C5205 AND2X1_LOC_364/A OR2X1_LOC_437/A 0.31fF
C5206 OR2X1_LOC_43/A OR2X1_LOC_88/Y 0.03fF
C5207 OR2X1_LOC_256/A OR2X1_LOC_71/Y 0.03fF
C5208 OR2X1_LOC_691/B OR2X1_LOC_857/B 0.01fF
C5209 AND2X1_LOC_56/B OR2X1_LOC_80/A 0.08fF
C5210 OR2X1_LOC_155/A OR2X1_LOC_228/Y 0.08fF
C5211 OR2X1_LOC_860/a_8_216# OR2X1_LOC_576/a_8_216# 0.47fF
C5212 OR2X1_LOC_64/Y OR2X1_LOC_597/Y 0.01fF
C5213 OR2X1_LOC_604/A OR2X1_LOC_744/a_8_216# 0.01fF
C5214 D_INPUT_4 AND2X1_LOC_36/Y 0.48fF
C5215 AND2X1_LOC_719/Y OR2X1_LOC_373/Y 0.03fF
C5216 OR2X1_LOC_523/Y OR2X1_LOC_523/A 0.95fF
C5217 AND2X1_LOC_8/Y OR2X1_LOC_80/A 0.07fF
C5218 AND2X1_LOC_734/a_8_24# VDD -0.00fF
C5219 OR2X1_LOC_629/B OR2X1_LOC_161/B 0.00fF
C5220 OR2X1_LOC_155/A OR2X1_LOC_513/Y 0.02fF
C5221 OR2X1_LOC_45/B OR2X1_LOC_694/Y 0.05fF
C5222 OR2X1_LOC_161/A OR2X1_LOC_349/B 0.01fF
C5223 OR2X1_LOC_45/B AND2X1_LOC_301/a_8_24# 0.02fF
C5224 OR2X1_LOC_124/B AND2X1_LOC_44/Y 0.28fF
C5225 VDD OR2X1_LOC_585/a_8_216# 0.00fF
C5226 OR2X1_LOC_31/Y OR2X1_LOC_428/Y 0.00fF
C5227 OR2X1_LOC_160/B AND2X1_LOC_255/a_8_24# 0.01fF
C5228 OR2X1_LOC_9/Y OR2X1_LOC_671/Y 0.02fF
C5229 AND2X1_LOC_568/B AND2X1_LOC_802/Y 0.01fF
C5230 AND2X1_LOC_535/Y AND2X1_LOC_809/a_36_24# 0.00fF
C5231 AND2X1_LOC_564/B OR2X1_LOC_329/B 0.02fF
C5232 AND2X1_LOC_40/Y OR2X1_LOC_168/Y 0.07fF
C5233 OR2X1_LOC_22/Y AND2X1_LOC_203/Y 0.08fF
C5234 AND2X1_LOC_363/Y OR2X1_LOC_12/Y 0.14fF
C5235 OR2X1_LOC_269/B OR2X1_LOC_732/A 0.01fF
C5236 OR2X1_LOC_468/A OR2X1_LOC_435/A 0.00fF
C5237 AND2X1_LOC_425/Y OR2X1_LOC_451/B 0.01fF
C5238 OR2X1_LOC_488/a_36_216# AND2X1_LOC_563/Y -0.00fF
C5239 OR2X1_LOC_188/Y AND2X1_LOC_368/a_36_24# 0.00fF
C5240 OR2X1_LOC_354/A OR2X1_LOC_703/a_8_216# 0.04fF
C5241 VDD OR2X1_LOC_492/Y 0.17fF
C5242 OR2X1_LOC_71/Y OR2X1_LOC_67/Y 0.01fF
C5243 AND2X1_LOC_434/Y AND2X1_LOC_774/A 0.10fF
C5244 OR2X1_LOC_158/A AND2X1_LOC_61/a_8_24# -0.01fF
C5245 AND2X1_LOC_719/Y OR2X1_LOC_666/a_8_216# 0.00fF
C5246 OR2X1_LOC_663/A OR2X1_LOC_227/B 0.01fF
C5247 OR2X1_LOC_87/B OR2X1_LOC_771/B 0.07fF
C5248 OR2X1_LOC_528/Y OR2X1_LOC_505/Y 0.04fF
C5249 OR2X1_LOC_334/B OR2X1_LOC_34/A 1.10fF
C5250 OR2X1_LOC_36/Y OR2X1_LOC_142/Y 0.02fF
C5251 AND2X1_LOC_4/a_8_24# OR2X1_LOC_71/A 0.00fF
C5252 OR2X1_LOC_676/Y OR2X1_LOC_596/a_8_216# 0.01fF
C5253 OR2X1_LOC_44/Y AND2X1_LOC_750/a_8_24# 0.01fF
C5254 AND2X1_LOC_59/Y OR2X1_LOC_388/a_8_216# 0.17fF
C5255 OR2X1_LOC_121/B OR2X1_LOC_560/A 0.03fF
C5256 D_INPUT_0 AND2X1_LOC_679/a_8_24# 0.17fF
C5257 VDD OR2X1_LOC_108/a_8_216# 0.21fF
C5258 AND2X1_LOC_362/B OR2X1_LOC_666/A 0.84fF
C5259 OR2X1_LOC_631/a_8_216# OR2X1_LOC_115/B 0.03fF
C5260 OR2X1_LOC_631/a_36_216# OR2X1_LOC_140/B 0.00fF
C5261 OR2X1_LOC_51/B OR2X1_LOC_587/a_8_216# 0.01fF
C5262 OR2X1_LOC_834/a_36_216# AND2X1_LOC_44/Y 0.00fF
C5263 OR2X1_LOC_3/Y OR2X1_LOC_437/A 0.09fF
C5264 INPUT_1 OR2X1_LOC_749/a_8_216# 0.01fF
C5265 OR2X1_LOC_528/Y AND2X1_LOC_658/A 0.03fF
C5266 AND2X1_LOC_110/Y OR2X1_LOC_66/A 0.03fF
C5267 AND2X1_LOC_554/B OR2X1_LOC_13/B 0.02fF
C5268 OR2X1_LOC_269/B OR2X1_LOC_539/B 0.27fF
C5269 OR2X1_LOC_158/A OR2X1_LOC_744/A 1.01fF
C5270 OR2X1_LOC_259/a_8_216# OR2X1_LOC_259/A 0.47fF
C5271 OR2X1_LOC_78/A OR2X1_LOC_786/a_36_216# 0.00fF
C5272 VDD OR2X1_LOC_426/B 2.02fF
C5273 AND2X1_LOC_64/Y OR2X1_LOC_500/A 0.01fF
C5274 AND2X1_LOC_43/B OR2X1_LOC_415/Y 0.08fF
C5275 OR2X1_LOC_175/Y OR2X1_LOC_624/A 0.29fF
C5276 OR2X1_LOC_67/Y D_INPUT_1 0.04fF
C5277 OR2X1_LOC_865/B OR2X1_LOC_576/A 0.02fF
C5278 AND2X1_LOC_311/a_8_24# AND2X1_LOC_110/Y 0.01fF
C5279 OR2X1_LOC_474/Y OR2X1_LOC_113/B 0.26fF
C5280 OR2X1_LOC_195/A AND2X1_LOC_36/Y 0.01fF
C5281 OR2X1_LOC_506/a_36_216# AND2X1_LOC_81/B 0.00fF
C5282 OR2X1_LOC_303/A OR2X1_LOC_302/A 0.86fF
C5283 AND2X1_LOC_12/Y AND2X1_LOC_7/B 0.24fF
C5284 OR2X1_LOC_97/A OR2X1_LOC_161/A 0.03fF
C5285 AND2X1_LOC_657/Y AND2X1_LOC_469/B 0.03fF
C5286 OR2X1_LOC_469/Y OR2X1_LOC_711/a_8_216# 0.40fF
C5287 OR2X1_LOC_574/A OR2X1_LOC_319/Y 0.15fF
C5288 OR2X1_LOC_709/A OR2X1_LOC_714/Y -0.02fF
C5289 OR2X1_LOC_624/A AND2X1_LOC_417/a_8_24# 0.03fF
C5290 AND2X1_LOC_786/a_8_24# OR2X1_LOC_265/Y 0.03fF
C5291 AND2X1_LOC_91/B OR2X1_LOC_468/Y 0.03fF
C5292 AND2X1_LOC_723/Y OR2X1_LOC_604/A 0.10fF
C5293 AND2X1_LOC_99/A OR2X1_LOC_595/A 0.03fF
C5294 OR2X1_LOC_389/A AND2X1_LOC_41/A 0.01fF
C5295 OR2X1_LOC_770/B OR2X1_LOC_402/Y 0.03fF
C5296 AND2X1_LOC_733/a_8_24# OR2X1_LOC_40/Y 0.02fF
C5297 AND2X1_LOC_543/Y AND2X1_LOC_374/Y 0.02fF
C5298 D_GATE_741 OR2X1_LOC_191/a_8_216# 0.39fF
C5299 AND2X1_LOC_364/Y AND2X1_LOC_352/B 0.04fF
C5300 OR2X1_LOC_290/a_8_216# OR2X1_LOC_600/A 0.05fF
C5301 OR2X1_LOC_134/Y OR2X1_LOC_26/Y 0.01fF
C5302 AND2X1_LOC_51/Y AND2X1_LOC_239/a_8_24# 0.03fF
C5303 OR2X1_LOC_589/A AND2X1_LOC_76/Y 0.02fF
C5304 OR2X1_LOC_656/Y AND2X1_LOC_18/Y 0.01fF
C5305 AND2X1_LOC_283/a_8_24# OR2X1_LOC_366/Y 0.27fF
C5306 OR2X1_LOC_391/B OR2X1_LOC_866/B 0.27fF
C5307 OR2X1_LOC_154/A OR2X1_LOC_857/A 0.08fF
C5308 OR2X1_LOC_507/A OR2X1_LOC_502/A 0.01fF
C5309 OR2X1_LOC_862/a_8_216# OR2X1_LOC_269/B 0.01fF
C5310 OR2X1_LOC_519/a_8_216# AND2X1_LOC_566/B 0.01fF
C5311 AND2X1_LOC_722/A OR2X1_LOC_51/Y 0.03fF
C5312 OR2X1_LOC_858/A OR2X1_LOC_735/a_8_216# 0.27fF
C5313 OR2X1_LOC_516/A AND2X1_LOC_515/a_8_24# 0.01fF
C5314 OR2X1_LOC_167/Y OR2X1_LOC_13/B 0.02fF
C5315 OR2X1_LOC_114/a_8_216# OR2X1_LOC_235/B 0.01fF
C5316 OR2X1_LOC_113/Y AND2X1_LOC_71/a_8_24# 0.08fF
C5317 OR2X1_LOC_276/B AND2X1_LOC_268/a_8_24# 0.02fF
C5318 VDD OR2X1_LOC_737/A 0.12fF
C5319 OR2X1_LOC_22/Y D_INPUT_6 0.00fF
C5320 AND2X1_LOC_231/Y OR2X1_LOC_52/B 0.01fF
C5321 OR2X1_LOC_744/A OR2X1_LOC_103/Y 0.03fF
C5322 OR2X1_LOC_7/A AND2X1_LOC_456/a_8_24# 0.01fF
C5323 OR2X1_LOC_375/A OR2X1_LOC_786/a_8_216# 0.01fF
C5324 OR2X1_LOC_76/B OR2X1_LOC_741/Y 0.79fF
C5325 AND2X1_LOC_22/Y OR2X1_LOC_654/A 0.19fF
C5326 OR2X1_LOC_671/Y OR2X1_LOC_96/B 0.19fF
C5327 OR2X1_LOC_744/A OR2X1_LOC_594/Y 0.10fF
C5328 VDD AND2X1_LOC_95/Y 2.04fF
C5329 OR2X1_LOC_319/B OR2X1_LOC_538/A 0.00fF
C5330 AND2X1_LOC_91/B OR2X1_LOC_846/B 0.00fF
C5331 OR2X1_LOC_186/Y AND2X1_LOC_187/a_8_24# 0.00fF
C5332 OR2X1_LOC_84/B OR2X1_LOC_161/B 0.13fF
C5333 OR2X1_LOC_281/a_8_216# OR2X1_LOC_56/A 0.01fF
C5334 OR2X1_LOC_7/A OR2X1_LOC_744/Y 0.01fF
C5335 OR2X1_LOC_449/B OR2X1_LOC_435/A 0.14fF
C5336 OR2X1_LOC_239/Y OR2X1_LOC_816/A 0.06fF
C5337 OR2X1_LOC_250/a_8_216# OR2X1_LOC_51/Y 0.01fF
C5338 VDD OR2X1_LOC_633/Y 0.25fF
C5339 AND2X1_LOC_361/a_8_24# AND2X1_LOC_560/B 0.02fF
C5340 OR2X1_LOC_114/B OR2X1_LOC_805/A 0.03fF
C5341 OR2X1_LOC_52/B AND2X1_LOC_770/a_8_24# 0.01fF
C5342 OR2X1_LOC_141/B OR2X1_LOC_161/B 0.03fF
C5343 AND2X1_LOC_658/B AND2X1_LOC_573/A 0.36fF
C5344 AND2X1_LOC_22/Y OR2X1_LOC_856/a_36_216# 0.01fF
C5345 OR2X1_LOC_97/A OR2X1_LOC_653/a_36_216# 0.00fF
C5346 OR2X1_LOC_812/a_8_216# OR2X1_LOC_269/B 0.02fF
C5347 AND2X1_LOC_728/Y AND2X1_LOC_803/B 0.00fF
C5348 OR2X1_LOC_318/Y OR2X1_LOC_538/A 0.12fF
C5349 AND2X1_LOC_566/B AND2X1_LOC_661/A 0.00fF
C5350 OR2X1_LOC_674/a_36_216# OR2X1_LOC_495/Y 0.00fF
C5351 OR2X1_LOC_158/A OR2X1_LOC_74/a_8_216# 0.02fF
C5352 OR2X1_LOC_40/Y OR2X1_LOC_85/A 1.52fF
C5353 OR2X1_LOC_849/A OR2X1_LOC_768/a_8_216# 0.01fF
C5354 OR2X1_LOC_851/B OR2X1_LOC_778/Y 0.19fF
C5355 INPUT_0 OR2X1_LOC_48/B 4.08fF
C5356 AND2X1_LOC_41/A AND2X1_LOC_422/a_8_24# 0.02fF
C5357 OR2X1_LOC_589/A OR2X1_LOC_52/B 0.08fF
C5358 AND2X1_LOC_474/A AND2X1_LOC_843/Y 0.00fF
C5359 OR2X1_LOC_664/Y OR2X1_LOC_66/A 0.05fF
C5360 OR2X1_LOC_51/Y AND2X1_LOC_454/Y 0.02fF
C5361 OR2X1_LOC_663/A OR2X1_LOC_509/A 0.02fF
C5362 OR2X1_LOC_160/B OR2X1_LOC_204/Y 0.03fF
C5363 VDD OR2X1_LOC_517/Y 0.12fF
C5364 INPUT_0 OR2X1_LOC_18/Y 0.06fF
C5365 AND2X1_LOC_2/Y OR2X1_LOC_375/A 0.01fF
C5366 OR2X1_LOC_739/A OR2X1_LOC_78/B 0.03fF
C5367 OR2X1_LOC_857/B OR2X1_LOC_688/a_36_216# 0.00fF
C5368 OR2X1_LOC_312/Y AND2X1_LOC_476/Y 0.01fF
C5369 OR2X1_LOC_97/A AND2X1_LOC_51/Y 0.03fF
C5370 OR2X1_LOC_32/B OR2X1_LOC_59/Y 0.11fF
C5371 OR2X1_LOC_604/A OR2X1_LOC_601/Y 0.01fF
C5372 OR2X1_LOC_52/Y AND2X1_LOC_208/Y 0.11fF
C5373 AND2X1_LOC_76/Y OR2X1_LOC_275/Y 0.01fF
C5374 OR2X1_LOC_866/B OR2X1_LOC_846/A 0.10fF
C5375 OR2X1_LOC_67/a_36_216# OR2X1_LOC_56/A 0.03fF
C5376 AND2X1_LOC_59/Y INPUT_0 0.07fF
C5377 OR2X1_LOC_756/B OR2X1_LOC_260/Y 0.07fF
C5378 OR2X1_LOC_22/Y AND2X1_LOC_242/B 0.02fF
C5379 D_INPUT_0 AND2X1_LOC_772/Y 0.82fF
C5380 AND2X1_LOC_19/Y AND2X1_LOC_129/a_36_24# 0.01fF
C5381 OR2X1_LOC_45/B AND2X1_LOC_308/a_8_24# 0.02fF
C5382 OR2X1_LOC_599/A OR2X1_LOC_51/Y 0.02fF
C5383 AND2X1_LOC_365/a_8_24# AND2X1_LOC_365/A 0.03fF
C5384 OR2X1_LOC_600/A AND2X1_LOC_458/a_8_24# 0.02fF
C5385 OR2X1_LOC_158/A OR2X1_LOC_282/a_8_216# 0.19fF
C5386 OR2X1_LOC_8/Y OR2X1_LOC_43/A 0.04fF
C5387 OR2X1_LOC_538/A OR2X1_LOC_805/A 0.03fF
C5388 OR2X1_LOC_56/A OR2X1_LOC_6/A 0.77fF
C5389 OR2X1_LOC_78/B OR2X1_LOC_798/a_8_216# 0.01fF
C5390 OR2X1_LOC_648/A OR2X1_LOC_87/A 0.01fF
C5391 OR2X1_LOC_837/Y AND2X1_LOC_233/a_8_24# 0.05fF
C5392 OR2X1_LOC_544/a_8_216# OR2X1_LOC_544/B 0.03fF
C5393 OR2X1_LOC_536/Y OR2X1_LOC_7/A 0.03fF
C5394 AND2X1_LOC_456/B AND2X1_LOC_848/Y 0.03fF
C5395 OR2X1_LOC_51/Y OR2X1_LOC_93/a_8_216# 0.01fF
C5396 OR2X1_LOC_856/B OR2X1_LOC_620/Y 0.41fF
C5397 AND2X1_LOC_736/a_8_24# OR2X1_LOC_189/A 0.22fF
C5398 OR2X1_LOC_380/Y OR2X1_LOC_588/Y 0.73fF
C5399 D_GATE_662 AND2X1_LOC_51/Y 0.14fF
C5400 OR2X1_LOC_675/Y OR2X1_LOC_580/A 0.07fF
C5401 OR2X1_LOC_80/A AND2X1_LOC_236/a_8_24# 0.02fF
C5402 AND2X1_LOC_555/Y AND2X1_LOC_866/A 0.05fF
C5403 OR2X1_LOC_769/a_36_216# OR2X1_LOC_598/A 0.00fF
C5404 OR2X1_LOC_114/B OR2X1_LOC_296/Y 0.00fF
C5405 AND2X1_LOC_722/A OR2X1_LOC_680/A 0.05fF
C5406 AND2X1_LOC_743/a_8_24# OR2X1_LOC_707/B 0.03fF
C5407 AND2X1_LOC_717/Y OR2X1_LOC_18/Y 0.09fF
C5408 OR2X1_LOC_68/B OR2X1_LOC_71/A 0.08fF
C5409 OR2X1_LOC_78/B OR2X1_LOC_269/B 5.09fF
C5410 VDD OR2X1_LOC_743/A 0.87fF
C5411 OR2X1_LOC_691/a_8_216# OR2X1_LOC_19/B 0.01fF
C5412 OR2X1_LOC_448/a_36_216# OR2X1_LOC_161/A 0.00fF
C5413 OR2X1_LOC_299/a_8_216# OR2X1_LOC_56/A 0.01fF
C5414 OR2X1_LOC_604/A OR2X1_LOC_754/A 0.40fF
C5415 OR2X1_LOC_807/Y OR2X1_LOC_807/B 0.84fF
C5416 AND2X1_LOC_550/a_8_24# AND2X1_LOC_711/Y 0.04fF
C5417 AND2X1_LOC_773/Y INPUT_1 0.10fF
C5418 AND2X1_LOC_550/a_8_24# OR2X1_LOC_70/Y 0.09fF
C5419 OR2X1_LOC_179/a_8_216# OR2X1_LOC_44/Y 0.02fF
C5420 OR2X1_LOC_287/B OR2X1_LOC_78/A 0.86fF
C5421 AND2X1_LOC_456/B OR2X1_LOC_283/Y 0.01fF
C5422 AND2X1_LOC_394/a_36_24# AND2X1_LOC_40/Y 0.01fF
C5423 OR2X1_LOC_840/A AND2X1_LOC_56/B 0.10fF
C5424 AND2X1_LOC_357/A OR2X1_LOC_64/Y 0.01fF
C5425 OR2X1_LOC_36/Y OR2X1_LOC_16/a_8_216# 0.01fF
C5426 OR2X1_LOC_847/A AND2X1_LOC_617/a_8_24# 0.01fF
C5427 OR2X1_LOC_561/B OR2X1_LOC_561/A 0.06fF
C5428 OR2X1_LOC_45/B AND2X1_LOC_270/a_8_24# 0.01fF
C5429 OR2X1_LOC_376/Y OR2X1_LOC_377/a_8_216# 0.01fF
C5430 AND2X1_LOC_474/A OR2X1_LOC_7/A 0.02fF
C5431 OR2X1_LOC_850/a_8_216# OR2X1_LOC_287/B 0.01fF
C5432 OR2X1_LOC_59/Y OR2X1_LOC_371/Y 0.07fF
C5433 OR2X1_LOC_121/B AND2X1_LOC_299/a_8_24# 0.03fF
C5434 OR2X1_LOC_62/B OR2X1_LOC_361/a_8_216# 0.01fF
C5435 OR2X1_LOC_154/A OR2X1_LOC_856/B 0.07fF
C5436 OR2X1_LOC_421/a_8_216# OR2X1_LOC_7/A 0.04fF
C5437 OR2X1_LOC_275/Y OR2X1_LOC_52/B 0.03fF
C5438 OR2X1_LOC_447/Y OR2X1_LOC_713/A 0.65fF
C5439 AND2X1_LOC_530/a_36_24# INPUT_1 0.01fF
C5440 OR2X1_LOC_548/A D_INPUT_0 0.01fF
C5441 OR2X1_LOC_665/a_8_216# OR2X1_LOC_600/A 0.01fF
C5442 AND2X1_LOC_59/Y OR2X1_LOC_732/B 0.03fF
C5443 OR2X1_LOC_681/a_8_216# AND2X1_LOC_687/A 0.03fF
C5444 AND2X1_LOC_47/Y AND2X1_LOC_277/a_36_24# 0.00fF
C5445 AND2X1_LOC_81/B OR2X1_LOC_493/A 0.05fF
C5446 OR2X1_LOC_18/Y OR2X1_LOC_11/Y 0.17fF
C5447 OR2X1_LOC_524/Y AND2X1_LOC_148/Y 0.03fF
C5448 AND2X1_LOC_753/a_36_24# OR2X1_LOC_375/A 0.00fF
C5449 OR2X1_LOC_97/a_8_216# OR2X1_LOC_78/A 0.01fF
C5450 OR2X1_LOC_611/a_8_216# OR2X1_LOC_600/A 0.02fF
C5451 OR2X1_LOC_235/B AND2X1_LOC_42/B 0.15fF
C5452 AND2X1_LOC_12/Y OR2X1_LOC_805/A 0.13fF
C5453 AND2X1_LOC_654/B OR2X1_LOC_52/B 0.00fF
C5454 AND2X1_LOC_86/Y OR2X1_LOC_204/Y 0.04fF
C5455 OR2X1_LOC_152/A OR2X1_LOC_142/Y 0.03fF
C5456 OR2X1_LOC_472/A OR2X1_LOC_852/B 0.05fF
C5457 VDD OR2X1_LOC_125/Y 0.12fF
C5458 AND2X1_LOC_340/Y AND2X1_LOC_476/A 0.07fF
C5459 AND2X1_LOC_319/a_8_24# OR2X1_LOC_428/A 0.03fF
C5460 OR2X1_LOC_502/A OR2X1_LOC_646/A 0.58fF
C5461 VDD OR2X1_LOC_246/A 1.15fF
C5462 OR2X1_LOC_427/A AND2X1_LOC_806/A 0.12fF
C5463 AND2X1_LOC_76/Y OR2X1_LOC_43/A 0.03fF
C5464 OR2X1_LOC_438/Y OR2X1_LOC_74/A 0.03fF
C5465 OR2X1_LOC_158/A OR2X1_LOC_31/Y 4.59fF
C5466 OR2X1_LOC_329/a_8_216# OR2X1_LOC_95/Y 0.01fF
C5467 AND2X1_LOC_453/a_8_24# AND2X1_LOC_466/a_8_24# 0.23fF
C5468 OR2X1_LOC_532/B OR2X1_LOC_362/A 0.10fF
C5469 OR2X1_LOC_36/Y OR2X1_LOC_118/Y 0.03fF
C5470 AND2X1_LOC_560/B OR2X1_LOC_18/Y 0.07fF
C5471 OR2X1_LOC_404/Y OR2X1_LOC_624/Y 0.00fF
C5472 AND2X1_LOC_94/Y OR2X1_LOC_19/B 0.03fF
C5473 OR2X1_LOC_173/Y OR2X1_LOC_18/Y 0.02fF
C5474 OR2X1_LOC_160/A OR2X1_LOC_643/A 0.07fF
C5475 OR2X1_LOC_18/Y OR2X1_LOC_690/A 0.03fF
C5476 AND2X1_LOC_356/B AND2X1_LOC_841/B 0.11fF
C5477 OR2X1_LOC_450/B OR2X1_LOC_707/B 0.01fF
C5478 OR2X1_LOC_504/Y AND2X1_LOC_806/a_8_24# 0.01fF
C5479 OR2X1_LOC_276/a_36_216# OR2X1_LOC_549/A 0.01fF
C5480 OR2X1_LOC_844/Y OR2X1_LOC_658/a_8_216# 0.01fF
C5481 AND2X1_LOC_763/a_8_24# AND2X1_LOC_48/A 0.03fF
C5482 AND2X1_LOC_43/B AND2X1_LOC_413/a_36_24# 0.01fF
C5483 OR2X1_LOC_160/A OR2X1_LOC_778/Y 0.10fF
C5484 AND2X1_LOC_217/Y AND2X1_LOC_227/Y 0.03fF
C5485 OR2X1_LOC_200/a_8_216# OR2X1_LOC_375/A 0.01fF
C5486 OR2X1_LOC_266/a_8_216# OR2X1_LOC_204/Y 0.39fF
C5487 AND2X1_LOC_571/A AND2X1_LOC_563/Y 0.00fF
C5488 OR2X1_LOC_696/a_8_216# OR2X1_LOC_427/A 0.02fF
C5489 AND2X1_LOC_390/B OR2X1_LOC_586/Y 0.79fF
C5490 OR2X1_LOC_856/B OR2X1_LOC_856/a_8_216# 0.05fF
C5491 OR2X1_LOC_375/A OR2X1_LOC_269/B 1.86fF
C5492 AND2X1_LOC_56/B OR2X1_LOC_241/a_36_216# 0.02fF
C5493 AND2X1_LOC_631/a_8_24# AND2X1_LOC_483/a_8_24# 0.23fF
C5494 OR2X1_LOC_676/Y AND2X1_LOC_47/Y 0.07fF
C5495 OR2X1_LOC_97/A OR2X1_LOC_551/B 0.08fF
C5496 OR2X1_LOC_427/A AND2X1_LOC_276/Y 0.01fF
C5497 OR2X1_LOC_32/a_8_216# OR2X1_LOC_39/A 0.01fF
C5498 OR2X1_LOC_26/Y AND2X1_LOC_859/a_8_24# 0.01fF
C5499 OR2X1_LOC_743/A OR2X1_LOC_829/a_8_216# 0.01fF
C5500 AND2X1_LOC_558/a_8_24# OR2X1_LOC_417/A 0.02fF
C5501 OR2X1_LOC_604/A OR2X1_LOC_55/a_36_216# 0.01fF
C5502 OR2X1_LOC_148/A OR2X1_LOC_78/A 0.01fF
C5503 OR2X1_LOC_743/A AND2X1_LOC_274/a_8_24# 0.24fF
C5504 OR2X1_LOC_426/B OR2X1_LOC_256/A 0.07fF
C5505 AND2X1_LOC_699/a_8_24# AND2X1_LOC_44/Y -0.01fF
C5506 OR2X1_LOC_272/a_8_216# OR2X1_LOC_18/Y 0.10fF
C5507 AND2X1_LOC_367/B OR2X1_LOC_417/A 0.08fF
C5508 OR2X1_LOC_343/B OR2X1_LOC_362/A 0.01fF
C5509 OR2X1_LOC_442/a_36_216# AND2X1_LOC_469/B 0.00fF
C5510 AND2X1_LOC_43/B OR2X1_LOC_378/Y 0.06fF
C5511 OR2X1_LOC_74/A AND2X1_LOC_621/Y 0.12fF
C5512 AND2X1_LOC_193/a_8_24# OR2X1_LOC_585/A 0.01fF
C5513 OR2X1_LOC_290/Y OR2X1_LOC_416/Y 0.01fF
C5514 AND2X1_LOC_729/Y AND2X1_LOC_147/Y 0.01fF
C5515 OR2X1_LOC_160/A OR2X1_LOC_647/A 0.06fF
C5516 OR2X1_LOC_262/Y OR2X1_LOC_36/Y 0.00fF
C5517 OR2X1_LOC_675/Y AND2X1_LOC_44/Y 0.02fF
C5518 OR2X1_LOC_51/Y AND2X1_LOC_866/A 0.03fF
C5519 OR2X1_LOC_7/A OR2X1_LOC_85/A 0.08fF
C5520 OR2X1_LOC_605/a_8_216# OR2X1_LOC_161/A 0.01fF
C5521 AND2X1_LOC_554/a_8_24# AND2X1_LOC_657/A 0.01fF
C5522 OR2X1_LOC_158/A OR2X1_LOC_257/Y 0.01fF
C5523 OR2X1_LOC_546/B OR2X1_LOC_375/A 0.01fF
C5524 AND2X1_LOC_54/a_8_24# AND2X1_LOC_28/a_8_24# 0.23fF
C5525 OR2X1_LOC_43/A OR2X1_LOC_52/B 0.21fF
C5526 OR2X1_LOC_64/Y OR2X1_LOC_48/B 0.26fF
C5527 OR2X1_LOC_635/A AND2X1_LOC_425/Y 0.01fF
C5528 OR2X1_LOC_43/A OR2X1_LOC_672/Y 0.01fF
C5529 OR2X1_LOC_36/Y OR2X1_LOC_238/Y 0.01fF
C5530 OR2X1_LOC_699/a_8_216# OR2X1_LOC_89/A 0.01fF
C5531 OR2X1_LOC_64/Y OR2X1_LOC_18/Y 0.38fF
C5532 OR2X1_LOC_653/Y AND2X1_LOC_48/A 0.42fF
C5533 OR2X1_LOC_474/Y OR2X1_LOC_532/B 0.06fF
C5534 OR2X1_LOC_3/Y AND2X1_LOC_348/Y 0.01fF
C5535 OR2X1_LOC_391/B OR2X1_LOC_557/A 0.01fF
C5536 AND2X1_LOC_59/Y OR2X1_LOC_401/A 0.09fF
C5537 OR2X1_LOC_648/A AND2X1_LOC_109/a_36_24# 0.01fF
C5538 OR2X1_LOC_539/A OR2X1_LOC_532/B 0.01fF
C5539 AND2X1_LOC_660/a_8_24# OR2X1_LOC_517/A 0.01fF
C5540 OR2X1_LOC_722/a_8_216# OR2X1_LOC_733/B 0.01fF
C5541 AND2X1_LOC_537/Y OR2X1_LOC_619/Y 0.07fF
C5542 OR2X1_LOC_3/Y OR2X1_LOC_753/A 0.13fF
C5543 AND2X1_LOC_486/Y OR2X1_LOC_71/Y 0.17fF
C5544 OR2X1_LOC_643/A OR2X1_LOC_624/B 0.03fF
C5545 AND2X1_LOC_391/Y OR2X1_LOC_47/Y 0.03fF
C5546 OR2X1_LOC_401/a_36_216# OR2X1_LOC_402/Y 0.01fF
C5547 OR2X1_LOC_513/a_8_216# OR2X1_LOC_713/A 0.01fF
C5548 AND2X1_LOC_116/a_8_24# OR2X1_LOC_59/Y 0.00fF
C5549 OR2X1_LOC_91/A OR2X1_LOC_47/Y 0.83fF
C5550 OR2X1_LOC_496/a_8_216# AND2X1_LOC_795/Y 0.47fF
C5551 OR2X1_LOC_426/B OR2X1_LOC_67/Y 0.89fF
C5552 AND2X1_LOC_115/a_8_24# OR2X1_LOC_39/A 0.02fF
C5553 AND2X1_LOC_43/a_8_24# AND2X1_LOC_3/Y 0.01fF
C5554 OR2X1_LOC_411/Y AND2X1_LOC_462/B 0.01fF
C5555 OR2X1_LOC_287/B OR2X1_LOC_392/a_8_216# 0.01fF
C5556 OR2X1_LOC_18/Y AND2X1_LOC_632/A 0.03fF
C5557 OR2X1_LOC_160/A OR2X1_LOC_113/A 0.05fF
C5558 OR2X1_LOC_18/Y AND2X1_LOC_471/a_36_24# 0.02fF
C5559 OR2X1_LOC_797/A OR2X1_LOC_161/A 0.13fF
C5560 AND2X1_LOC_571/Y OR2X1_LOC_71/Y 0.01fF
C5561 OR2X1_LOC_18/Y OR2X1_LOC_417/A 1.28fF
C5562 AND2X1_LOC_191/B AND2X1_LOC_848/A 0.07fF
C5563 AND2X1_LOC_532/a_8_24# AND2X1_LOC_810/Y 0.07fF
C5564 OR2X1_LOC_844/a_8_216# AND2X1_LOC_42/B 0.01fF
C5565 AND2X1_LOC_727/A AND2X1_LOC_653/a_8_24# 0.01fF
C5566 OR2X1_LOC_245/a_8_216# AND2X1_LOC_361/A 0.03fF
C5567 OR2X1_LOC_70/Y OR2X1_LOC_371/Y 0.03fF
C5568 AND2X1_LOC_151/a_8_24# AND2X1_LOC_727/A 0.01fF
C5569 AND2X1_LOC_685/a_8_24# OR2X1_LOC_52/B 0.03fF
C5570 AND2X1_LOC_390/a_8_24# OR2X1_LOC_534/Y 0.02fF
C5571 AND2X1_LOC_572/A AND2X1_LOC_845/Y 0.01fF
C5572 AND2X1_LOC_41/A OR2X1_LOC_493/Y 0.01fF
C5573 OR2X1_LOC_687/B AND2X1_LOC_425/Y 0.01fF
C5574 AND2X1_LOC_41/A OR2X1_LOC_801/B 0.07fF
C5575 OR2X1_LOC_403/B OR2X1_LOC_403/a_8_216# 0.05fF
C5576 OR2X1_LOC_50/a_8_216# OR2X1_LOC_2/Y 0.02fF
C5577 OR2X1_LOC_244/A OR2X1_LOC_204/Y 0.03fF
C5578 OR2X1_LOC_59/Y AND2X1_LOC_222/Y 0.03fF
C5579 OR2X1_LOC_804/A OR2X1_LOC_776/a_36_216# 0.00fF
C5580 AND2X1_LOC_788/a_8_24# OR2X1_LOC_13/B 0.04fF
C5581 OR2X1_LOC_833/Y OR2X1_LOC_777/B 0.11fF
C5582 OR2X1_LOC_291/Y AND2X1_LOC_640/Y 0.01fF
C5583 OR2X1_LOC_462/B AND2X1_LOC_47/Y 0.02fF
C5584 OR2X1_LOC_76/A OR2X1_LOC_605/A 0.19fF
C5585 OR2X1_LOC_741/Y OR2X1_LOC_578/B 0.03fF
C5586 AND2X1_LOC_510/A AND2X1_LOC_657/A 0.03fF
C5587 OR2X1_LOC_680/A AND2X1_LOC_866/A 0.02fF
C5588 AND2X1_LOC_477/Y OR2X1_LOC_437/A 0.46fF
C5589 OR2X1_LOC_858/A OR2X1_LOC_68/B 0.01fF
C5590 AND2X1_LOC_362/B OR2X1_LOC_13/B 0.00fF
C5591 OR2X1_LOC_75/Y OR2X1_LOC_265/Y 0.15fF
C5592 OR2X1_LOC_47/Y AND2X1_LOC_573/A 0.02fF
C5593 AND2X1_LOC_37/a_8_24# OR2X1_LOC_54/Y 0.01fF
C5594 OR2X1_LOC_751/A OR2X1_LOC_44/Y 0.28fF
C5595 OR2X1_LOC_615/Y OR2X1_LOC_39/A 0.03fF
C5596 OR2X1_LOC_431/Y OR2X1_LOC_304/Y 0.73fF
C5597 AND2X1_LOC_859/B OR2X1_LOC_44/Y 0.01fF
C5598 OR2X1_LOC_177/Y OR2X1_LOC_142/Y 0.03fF
C5599 OR2X1_LOC_421/Y AND2X1_LOC_449/a_8_24# 0.01fF
C5600 AND2X1_LOC_56/B OR2X1_LOC_241/Y 0.09fF
C5601 OR2X1_LOC_140/B OR2X1_LOC_554/a_8_216# 0.03fF
C5602 VDD OR2X1_LOC_269/A -0.00fF
C5603 OR2X1_LOC_415/Y AND2X1_LOC_416/a_8_24# 0.11fF
C5604 OR2X1_LOC_427/A AND2X1_LOC_405/a_8_24# 0.01fF
C5605 OR2X1_LOC_226/Y OR2X1_LOC_7/A 0.03fF
C5606 OR2X1_LOC_66/A OR2X1_LOC_342/a_8_216# 0.02fF
C5607 OR2X1_LOC_436/Y OR2X1_LOC_155/A 0.03fF
C5608 OR2X1_LOC_6/B OR2X1_LOC_749/Y 0.01fF
C5609 OR2X1_LOC_3/Y AND2X1_LOC_845/Y 0.04fF
C5610 OR2X1_LOC_756/B OR2X1_LOC_364/Y 0.01fF
C5611 OR2X1_LOC_291/Y OR2X1_LOC_416/Y 0.02fF
C5612 VDD OR2X1_LOC_788/B 0.02fF
C5613 AND2X1_LOC_749/a_8_24# OR2X1_LOC_68/B 0.03fF
C5614 OR2X1_LOC_39/A AND2X1_LOC_203/Y 0.01fF
C5615 AND2X1_LOC_476/A OR2X1_LOC_585/A 0.07fF
C5616 OR2X1_LOC_866/a_8_216# D_INPUT_1 0.01fF
C5617 OR2X1_LOC_476/B OR2X1_LOC_650/Y 0.07fF
C5618 OR2X1_LOC_848/A OR2X1_LOC_770/Y 0.03fF
C5619 OR2X1_LOC_702/a_8_216# OR2X1_LOC_515/Y 0.55fF
C5620 OR2X1_LOC_329/B OR2X1_LOC_437/A 0.11fF
C5621 OR2X1_LOC_151/A OR2X1_LOC_388/a_36_216# 0.02fF
C5622 OR2X1_LOC_856/B OR2X1_LOC_198/A 0.04fF
C5623 OR2X1_LOC_108/Y OR2X1_LOC_183/Y 0.01fF
C5624 AND2X1_LOC_172/a_8_24# OR2X1_LOC_539/B 0.17fF
C5625 OR2X1_LOC_276/B AND2X1_LOC_42/B 0.07fF
C5626 AND2X1_LOC_44/Y OR2X1_LOC_779/A 0.06fF
C5627 OR2X1_LOC_462/B OR2X1_LOC_598/A 0.00fF
C5628 AND2X1_LOC_462/B OR2X1_LOC_753/A 0.10fF
C5629 OR2X1_LOC_111/a_8_216# AND2X1_LOC_476/Y 0.10fF
C5630 OR2X1_LOC_631/B OR2X1_LOC_493/Y 0.03fF
C5631 AND2X1_LOC_110/Y OR2X1_LOC_354/a_36_216# 0.00fF
C5632 OR2X1_LOC_769/B AND2X1_LOC_36/Y 0.07fF
C5633 OR2X1_LOC_49/A OR2X1_LOC_414/Y 0.01fF
C5634 OR2X1_LOC_778/Y OR2X1_LOC_717/a_8_216# 0.01fF
C5635 AND2X1_LOC_555/Y OR2X1_LOC_40/Y 0.02fF
C5636 AND2X1_LOC_786/Y AND2X1_LOC_795/a_8_24# 0.08fF
C5637 AND2X1_LOC_43/B OR2X1_LOC_378/A 0.50fF
C5638 OR2X1_LOC_419/Y OR2X1_LOC_238/Y 0.05fF
C5639 OR2X1_LOC_696/A AND2X1_LOC_705/a_36_24# 0.01fF
C5640 OR2X1_LOC_736/Y AND2X1_LOC_44/Y 0.43fF
C5641 OR2X1_LOC_186/Y OR2X1_LOC_161/B 0.06fF
C5642 AND2X1_LOC_715/Y OR2X1_LOC_329/Y 0.01fF
C5643 OR2X1_LOC_808/A OR2X1_LOC_593/B 0.19fF
C5644 AND2X1_LOC_539/Y AND2X1_LOC_567/a_8_24# 0.04fF
C5645 AND2X1_LOC_712/a_8_24# OR2X1_LOC_421/Y 0.01fF
C5646 OR2X1_LOC_136/Y OR2X1_LOC_40/Y 0.01fF
C5647 OR2X1_LOC_648/A OR2X1_LOC_390/B 1.20fF
C5648 AND2X1_LOC_706/Y AND2X1_LOC_724/A 0.02fF
C5649 AND2X1_LOC_774/a_8_24# OR2X1_LOC_589/A 0.03fF
C5650 AND2X1_LOC_573/Y AND2X1_LOC_501/a_8_24# 0.09fF
C5651 AND2X1_LOC_41/A OR2X1_LOC_130/a_8_216# 0.01fF
C5652 OR2X1_LOC_158/A AND2X1_LOC_213/B 0.12fF
C5653 AND2X1_LOC_634/Y AND2X1_LOC_476/A 0.03fF
C5654 OR2X1_LOC_36/Y OR2X1_LOC_39/a_8_216# 0.01fF
C5655 OR2X1_LOC_187/Y VDD 0.12fF
C5656 OR2X1_LOC_784/Y OR2X1_LOC_712/B 0.05fF
C5657 AND2X1_LOC_191/Y AND2X1_LOC_222/Y 0.03fF
C5658 OR2X1_LOC_469/Y OR2X1_LOC_308/Y 0.02fF
C5659 AND2X1_LOC_22/Y VDD 0.73fF
C5660 AND2X1_LOC_423/a_8_24# OR2X1_LOC_308/Y 0.03fF
C5661 OR2X1_LOC_19/B OR2X1_LOC_214/B 0.07fF
C5662 OR2X1_LOC_802/Y OR2X1_LOC_446/B 0.90fF
C5663 AND2X1_LOC_711/Y AND2X1_LOC_222/Y 0.03fF
C5664 AND2X1_LOC_619/B AND2X1_LOC_619/a_8_24# 0.19fF
C5665 OR2X1_LOC_786/a_8_216# OR2X1_LOC_549/A 0.01fF
C5666 OR2X1_LOC_114/B OR2X1_LOC_580/B 0.03fF
C5667 OR2X1_LOC_70/Y AND2X1_LOC_222/Y 0.03fF
C5668 OR2X1_LOC_641/Y AND2X1_LOC_44/Y 0.03fF
C5669 OR2X1_LOC_319/B OR2X1_LOC_356/B 0.23fF
C5670 OR2X1_LOC_246/A OR2X1_LOC_67/Y 0.07fF
C5671 OR2X1_LOC_468/Y OR2X1_LOC_303/B 0.03fF
C5672 OR2X1_LOC_479/Y AND2X1_LOC_31/Y 0.19fF
C5673 AND2X1_LOC_632/A AND2X1_LOC_620/Y 0.01fF
C5674 AND2X1_LOC_469/B AND2X1_LOC_804/A 0.01fF
C5675 AND2X1_LOC_721/Y OR2X1_LOC_744/A 0.02fF
C5676 OR2X1_LOC_160/B OR2X1_LOC_663/a_8_216# 0.02fF
C5677 AND2X1_LOC_70/Y OR2X1_LOC_855/a_8_216# 0.01fF
C5678 OR2X1_LOC_351/B OR2X1_LOC_648/B 0.10fF
C5679 OR2X1_LOC_319/a_8_216# OR2X1_LOC_319/Y -0.00fF
C5680 AND2X1_LOC_383/a_8_24# OR2X1_LOC_292/Y 0.23fF
C5681 AND2X1_LOC_388/Y AND2X1_LOC_390/a_8_24# 0.01fF
C5682 D_INPUT_0 OR2X1_LOC_66/a_8_216# 0.02fF
C5683 VDD OR2X1_LOC_467/B 0.04fF
C5684 OR2X1_LOC_600/A OR2X1_LOC_13/Y 0.03fF
C5685 AND2X1_LOC_219/Y AND2X1_LOC_786/Y 0.02fF
C5686 AND2X1_LOC_733/Y AND2X1_LOC_804/A 0.02fF
C5687 OR2X1_LOC_604/A AND2X1_LOC_347/B 0.04fF
C5688 OR2X1_LOC_74/A OR2X1_LOC_71/A 0.04fF
C5689 VDD OR2X1_LOC_621/A 0.21fF
C5690 OR2X1_LOC_176/Y AND2X1_LOC_723/Y 0.08fF
C5691 OR2X1_LOC_97/A OR2X1_LOC_640/A 0.09fF
C5692 OR2X1_LOC_580/a_8_216# OR2X1_LOC_286/B 0.01fF
C5693 AND2X1_LOC_43/B OR2X1_LOC_168/Y 0.03fF
C5694 OR2X1_LOC_291/Y OR2X1_LOC_80/A 0.07fF
C5695 OR2X1_LOC_808/B AND2X1_LOC_44/Y 0.02fF
C5696 OR2X1_LOC_696/A AND2X1_LOC_435/a_36_24# 0.01fF
C5697 AND2X1_LOC_41/A AND2X1_LOC_255/a_36_24# 0.01fF
C5698 OR2X1_LOC_40/Y OR2X1_LOC_51/Y 3.05fF
C5699 OR2X1_LOC_814/A OR2X1_LOC_228/Y 0.11fF
C5700 OR2X1_LOC_482/Y OR2X1_LOC_744/A 0.10fF
C5701 AND2X1_LOC_658/B AND2X1_LOC_806/a_8_24# 0.00fF
C5702 OR2X1_LOC_516/a_36_216# OR2X1_LOC_26/Y 0.02fF
C5703 AND2X1_LOC_91/B OR2X1_LOC_160/A 0.37fF
C5704 AND2X1_LOC_59/Y OR2X1_LOC_214/A 0.01fF
C5705 AND2X1_LOC_785/A OR2X1_LOC_26/Y 0.01fF
C5706 OR2X1_LOC_375/A OR2X1_LOC_718/a_36_216# 0.00fF
C5707 AND2X1_LOC_561/a_8_24# OR2X1_LOC_26/Y 0.17fF
C5708 OR2X1_LOC_160/B OR2X1_LOC_78/A 0.12fF
C5709 OR2X1_LOC_45/B OR2X1_LOC_695/a_36_216# 0.02fF
C5710 OR2X1_LOC_175/Y OR2X1_LOC_161/A 0.07fF
C5711 OR2X1_LOC_429/Y D_INPUT_6 0.04fF
C5712 AND2X1_LOC_347/a_8_24# AND2X1_LOC_789/Y 0.02fF
C5713 AND2X1_LOC_242/B OR2X1_LOC_39/A 0.03fF
C5714 AND2X1_LOC_40/Y OR2X1_LOC_486/Y 0.07fF
C5715 OR2X1_LOC_759/A AND2X1_LOC_663/A 0.03fF
C5716 AND2X1_LOC_59/Y AND2X1_LOC_7/B 0.38fF
C5717 OR2X1_LOC_329/B AND2X1_LOC_715/A 0.09fF
C5718 AND2X1_LOC_172/a_8_24# OR2X1_LOC_78/B 0.01fF
C5719 AND2X1_LOC_785/A OR2X1_LOC_89/A 0.09fF
C5720 AND2X1_LOC_486/Y OR2X1_LOC_492/Y 0.03fF
C5721 OR2X1_LOC_149/B OR2X1_LOC_87/A 0.07fF
C5722 AND2X1_LOC_561/a_8_24# OR2X1_LOC_89/A 0.01fF
C5723 VDD OR2X1_LOC_244/B 0.12fF
C5724 OR2X1_LOC_517/A AND2X1_LOC_243/Y 0.07fF
C5725 OR2X1_LOC_512/A OR2X1_LOC_307/A 0.25fF
C5726 AND2X1_LOC_716/Y AND2X1_LOC_182/a_8_24# 0.02fF
C5727 OR2X1_LOC_756/B AND2X1_LOC_18/Y 0.59fF
C5728 OR2X1_LOC_691/Y OR2X1_LOC_161/A 0.03fF
C5729 AND2X1_LOC_712/Y OR2X1_LOC_92/Y 0.03fF
C5730 VDD OR2X1_LOC_706/A 0.21fF
C5731 OR2X1_LOC_691/A OR2X1_LOC_377/A 0.01fF
C5732 AND2X1_LOC_218/Y AND2X1_LOC_219/Y 0.11fF
C5733 OR2X1_LOC_106/Y OR2X1_LOC_26/Y 0.03fF
C5734 VDD OR2X1_LOC_298/a_8_216# 0.21fF
C5735 AND2X1_LOC_47/a_36_24# AND2X1_LOC_44/Y 0.00fF
C5736 OR2X1_LOC_744/A OR2X1_LOC_816/Y 0.14fF
C5737 AND2X1_LOC_12/Y OR2X1_LOC_580/B 0.05fF
C5738 OR2X1_LOC_329/B AND2X1_LOC_851/a_8_24# 0.01fF
C5739 OR2X1_LOC_604/A OR2X1_LOC_683/a_8_216# 0.01fF
C5740 AND2X1_LOC_721/Y AND2X1_LOC_840/B 0.03fF
C5741 AND2X1_LOC_553/A OR2X1_LOC_108/Y 0.00fF
C5742 GATE_479 AND2X1_LOC_223/a_36_24# 0.00fF
C5743 D_INPUT_3 OR2X1_LOC_80/A 0.23fF
C5744 OR2X1_LOC_240/a_8_216# OR2X1_LOC_549/A 0.40fF
C5745 OR2X1_LOC_448/A OR2X1_LOC_66/A 0.03fF
C5746 AND2X1_LOC_367/A OR2X1_LOC_59/Y 0.05fF
C5747 OR2X1_LOC_670/a_8_216# OR2X1_LOC_428/A 0.01fF
C5748 OR2X1_LOC_437/Y AND2X1_LOC_222/Y -0.01fF
C5749 OR2X1_LOC_45/B OR2X1_LOC_271/a_36_216# 0.00fF
C5750 OR2X1_LOC_849/A OR2X1_LOC_474/B 0.00fF
C5751 AND2X1_LOC_640/Y OR2X1_LOC_171/Y 0.02fF
C5752 OR2X1_LOC_106/Y OR2X1_LOC_89/A 0.18fF
C5753 AND2X1_LOC_719/Y OR2X1_LOC_109/Y 0.10fF
C5754 AND2X1_LOC_543/Y OR2X1_LOC_280/Y 0.01fF
C5755 AND2X1_LOC_144/a_8_24# AND2X1_LOC_41/A 0.04fF
C5756 AND2X1_LOC_91/B AND2X1_LOC_86/B 0.01fF
C5757 OR2X1_LOC_524/Y AND2X1_LOC_545/a_8_24# 0.07fF
C5758 OR2X1_LOC_405/A OR2X1_LOC_730/A 0.01fF
C5759 OR2X1_LOC_691/B OR2X1_LOC_835/B 0.01fF
C5760 OR2X1_LOC_510/A AND2X1_LOC_504/a_8_24# 0.01fF
C5761 OR2X1_LOC_185/A OR2X1_LOC_641/A 0.23fF
C5762 OR2X1_LOC_840/A AND2X1_LOC_92/Y 0.17fF
C5763 VDD OR2X1_LOC_525/Y 0.05fF
C5764 OR2X1_LOC_708/B AND2X1_LOC_44/Y 0.03fF
C5765 OR2X1_LOC_26/Y AND2X1_LOC_219/A 0.67fF
C5766 OR2X1_LOC_235/B OR2X1_LOC_663/A 0.03fF
C5767 AND2X1_LOC_91/B OR2X1_LOC_624/B 0.07fF
C5768 AND2X1_LOC_586/a_36_24# OR2X1_LOC_598/Y 0.00fF
C5769 AND2X1_LOC_12/Y OR2X1_LOC_648/B 0.02fF
C5770 AND2X1_LOC_778/a_8_24# AND2X1_LOC_785/Y 0.23fF
C5771 OR2X1_LOC_496/Y AND2X1_LOC_786/Y 0.04fF
C5772 AND2X1_LOC_93/a_36_24# OR2X1_LOC_633/Y 0.01fF
C5773 OR2X1_LOC_813/a_36_216# OR2X1_LOC_278/Y 0.00fF
C5774 OR2X1_LOC_477/B OR2X1_LOC_161/B 0.01fF
C5775 OR2X1_LOC_532/B OR2X1_LOC_771/B 0.06fF
C5776 OR2X1_LOC_689/a_8_216# OR2X1_LOC_690/Y 0.40fF
C5777 OR2X1_LOC_493/B OR2X1_LOC_493/A 0.02fF
C5778 OR2X1_LOC_474/Y OR2X1_LOC_624/Y 0.01fF
C5779 OR2X1_LOC_863/a_8_216# OR2X1_LOC_863/A 0.39fF
C5780 OR2X1_LOC_43/A OR2X1_LOC_9/a_8_216# 0.02fF
C5781 OR2X1_LOC_121/B OR2X1_LOC_605/Y 0.01fF
C5782 OR2X1_LOC_51/Y AND2X1_LOC_843/Y 0.01fF
C5783 AND2X1_LOC_60/a_36_24# OR2X1_LOC_219/B 0.01fF
C5784 OR2X1_LOC_485/A AND2X1_LOC_242/a_8_24# 0.02fF
C5785 OR2X1_LOC_160/A AND2X1_LOC_86/a_36_24# 0.00fF
C5786 OR2X1_LOC_532/B OR2X1_LOC_209/A 0.09fF
C5787 OR2X1_LOC_440/A OR2X1_LOC_544/B 0.88fF
C5788 VDD OR2X1_LOC_664/a_8_216# 0.21fF
C5789 OR2X1_LOC_310/Y OR2X1_LOC_92/Y 0.13fF
C5790 OR2X1_LOC_43/A OR2X1_LOC_13/a_8_216# 0.04fF
C5791 OR2X1_LOC_40/Y OR2X1_LOC_680/A 10.75fF
C5792 OR2X1_LOC_604/A AND2X1_LOC_453/a_8_24# 0.01fF
C5793 AND2X1_LOC_334/a_36_24# OR2X1_LOC_26/Y 0.00fF
C5794 OR2X1_LOC_482/Y AND2X1_LOC_840/B 0.02fF
C5795 OR2X1_LOC_269/B OR2X1_LOC_549/A 0.07fF
C5796 AND2X1_LOC_554/B OR2X1_LOC_428/A 0.01fF
C5797 AND2X1_LOC_27/a_8_24# OR2X1_LOC_334/A 0.01fF
C5798 AND2X1_LOC_86/Y OR2X1_LOC_78/A 0.02fF
C5799 AND2X1_LOC_41/A OR2X1_LOC_61/B 0.09fF
C5800 VDD AND2X1_LOC_153/a_8_24# -0.00fF
C5801 AND2X1_LOC_76/a_36_24# OR2X1_LOC_59/Y 0.00fF
C5802 AND2X1_LOC_668/a_8_24# AND2X1_LOC_860/A 0.01fF
C5803 OR2X1_LOC_175/Y AND2X1_LOC_51/Y 0.14fF
C5804 OR2X1_LOC_45/a_8_216# OR2X1_LOC_56/A 0.03fF
C5805 OR2X1_LOC_822/a_8_216# OR2X1_LOC_85/A 0.01fF
C5806 OR2X1_LOC_532/B OR2X1_LOC_776/A 0.03fF
C5807 AND2X1_LOC_724/A OR2X1_LOC_485/A 0.21fF
C5808 AND2X1_LOC_173/a_36_24# OR2X1_LOC_538/A 0.00fF
C5809 AND2X1_LOC_554/B OR2X1_LOC_595/A 0.02fF
C5810 OR2X1_LOC_615/a_8_216# OR2X1_LOC_816/A 0.03fF
C5811 OR2X1_LOC_542/B OR2X1_LOC_457/B 0.14fF
C5812 OR2X1_LOC_64/Y OR2X1_LOC_764/a_8_216# 0.01fF
C5813 AND2X1_LOC_182/a_8_24# OR2X1_LOC_312/Y 0.02fF
C5814 AND2X1_LOC_593/a_36_24# OR2X1_LOC_599/A 0.00fF
C5815 OR2X1_LOC_770/A OR2X1_LOC_401/a_8_216# 0.47fF
C5816 OR2X1_LOC_228/Y OR2X1_LOC_341/a_8_216# 0.03fF
C5817 D_INPUT_5 OR2X1_LOC_2/Y 0.02fF
C5818 OR2X1_LOC_525/Y OR2X1_LOC_677/Y 0.01fF
C5819 AND2X1_LOC_842/B OR2X1_LOC_816/A 0.12fF
C5820 VDD OR2X1_LOC_86/Y 0.12fF
C5821 OR2X1_LOC_76/Y AND2X1_LOC_18/Y 0.02fF
C5822 OR2X1_LOC_441/Y OR2X1_LOC_427/A 0.06fF
C5823 OR2X1_LOC_691/Y AND2X1_LOC_51/Y 0.03fF
C5824 OR2X1_LOC_78/B OR2X1_LOC_539/Y 1.55fF
C5825 AND2X1_LOC_31/Y OR2X1_LOC_68/B 0.71fF
C5826 AND2X1_LOC_647/Y OR2X1_LOC_71/A 0.03fF
C5827 AND2X1_LOC_95/Y OR2X1_LOC_334/B 0.00fF
C5828 AND2X1_LOC_64/Y AND2X1_LOC_69/a_8_24# 0.02fF
C5829 VDD OR2X1_LOC_497/Y 0.39fF
C5830 OR2X1_LOC_482/Y AND2X1_LOC_719/a_8_24# 0.23fF
C5831 OR2X1_LOC_810/A OR2X1_LOC_631/A 0.03fF
C5832 OR2X1_LOC_533/A OR2X1_LOC_331/Y 0.01fF
C5833 AND2X1_LOC_66/a_36_24# OR2X1_LOC_26/Y 0.01fF
C5834 OR2X1_LOC_646/a_36_216# OR2X1_LOC_646/B 0.00fF
C5835 AND2X1_LOC_728/Y OR2X1_LOC_524/Y 0.06fF
C5836 OR2X1_LOC_422/Y OR2X1_LOC_92/Y 0.01fF
C5837 OR2X1_LOC_222/A AND2X1_LOC_92/Y 0.02fF
C5838 AND2X1_LOC_117/a_8_24# AND2X1_LOC_65/A 0.10fF
C5839 OR2X1_LOC_62/B OR2X1_LOC_267/Y 0.01fF
C5840 AND2X1_LOC_738/B OR2X1_LOC_44/Y 0.04fF
C5841 OR2X1_LOC_160/B OR2X1_LOC_155/A 0.21fF
C5842 AND2X1_LOC_509/a_8_24# OR2X1_LOC_44/Y 0.01fF
C5843 AND2X1_LOC_340/Y OR2X1_LOC_64/Y 0.03fF
C5844 OR2X1_LOC_604/A OR2X1_LOC_238/Y 0.03fF
C5845 OR2X1_LOC_56/A OR2X1_LOC_44/Y 0.26fF
C5846 AND2X1_LOC_51/Y OR2X1_LOC_713/A 0.19fF
C5847 OR2X1_LOC_78/A OR2X1_LOC_779/a_36_216# 0.00fF
C5848 OR2X1_LOC_140/A AND2X1_LOC_3/Y 0.03fF
C5849 AND2X1_LOC_710/Y OR2X1_LOC_44/Y 0.01fF
C5850 AND2X1_LOC_658/A OR2X1_LOC_26/Y 0.03fF
C5851 OR2X1_LOC_640/Y AND2X1_LOC_8/Y 0.03fF
C5852 AND2X1_LOC_231/Y OR2X1_LOC_22/Y 0.00fF
C5853 OR2X1_LOC_158/A OR2X1_LOC_488/a_8_216# 0.02fF
C5854 OR2X1_LOC_819/a_8_216# OR2X1_LOC_44/Y 0.01fF
C5855 AND2X1_LOC_392/A AND2X1_LOC_566/Y 0.67fF
C5856 OR2X1_LOC_92/Y OR2X1_LOC_433/Y 0.20fF
C5857 AND2X1_LOC_787/A AND2X1_LOC_477/A 0.15fF
C5858 AND2X1_LOC_514/a_8_24# OR2X1_LOC_43/A 0.03fF
C5859 OR2X1_LOC_185/Y OR2X1_LOC_235/B 0.05fF
C5860 OR2X1_LOC_319/B AND2X1_LOC_59/Y 0.05fF
C5861 OR2X1_LOC_683/a_36_216# AND2X1_LOC_452/Y 0.00fF
C5862 OR2X1_LOC_8/Y AND2X1_LOC_240/Y 0.05fF
C5863 OR2X1_LOC_490/a_8_216# OR2X1_LOC_19/B 0.01fF
C5864 OR2X1_LOC_51/Y OR2X1_LOC_7/A 2.92fF
C5865 AND2X1_LOC_658/A OR2X1_LOC_89/A 0.03fF
C5866 VDD OR2X1_LOC_229/Y 0.12fF
C5867 OR2X1_LOC_62/B OR2X1_LOC_633/A 0.03fF
C5868 AND2X1_LOC_159/a_8_24# OR2X1_LOC_632/Y 0.02fF
C5869 OR2X1_LOC_339/a_8_216# OR2X1_LOC_333/B 0.01fF
C5870 AND2X1_LOC_40/Y AND2X1_LOC_80/a_8_24# 0.01fF
C5871 AND2X1_LOC_41/A OR2X1_LOC_205/a_8_216# 0.07fF
C5872 AND2X1_LOC_378/a_8_24# OR2X1_LOC_43/A 0.04fF
C5873 OR2X1_LOC_374/Y OR2X1_LOC_593/B 0.03fF
C5874 D_GATE_865 OR2X1_LOC_391/A 0.02fF
C5875 OR2X1_LOC_666/A OR2X1_LOC_485/A 0.03fF
C5876 OR2X1_LOC_810/A OR2X1_LOC_632/Y 0.10fF
C5877 OR2X1_LOC_612/B OR2X1_LOC_612/Y 0.01fF
C5878 INPUT_0 OR2X1_LOC_585/A 0.03fF
C5879 AND2X1_LOC_59/Y OR2X1_LOC_318/Y 0.01fF
C5880 AND2X1_LOC_721/Y OR2X1_LOC_31/Y 0.18fF
C5881 AND2X1_LOC_706/a_8_24# OR2X1_LOC_22/Y 0.02fF
C5882 AND2X1_LOC_640/a_8_24# OR2X1_LOC_16/A 0.01fF
C5883 OR2X1_LOC_532/B OR2X1_LOC_721/a_36_216# 0.00fF
C5884 AND2X1_LOC_716/Y AND2X1_LOC_303/A 0.01fF
C5885 AND2X1_LOC_456/Y OR2X1_LOC_59/Y 0.00fF
C5886 AND2X1_LOC_70/Y AND2X1_LOC_42/B 0.03fF
C5887 INPUT_1 OR2X1_LOC_12/Y 0.17fF
C5888 AND2X1_LOC_638/Y OR2X1_LOC_44/Y 0.04fF
C5889 AND2X1_LOC_116/Y OR2X1_LOC_56/A 0.04fF
C5890 OR2X1_LOC_481/a_8_216# OR2X1_LOC_700/a_8_216# 0.47fF
C5891 OR2X1_LOC_589/A OR2X1_LOC_22/Y 0.49fF
C5892 OR2X1_LOC_348/Y OR2X1_LOC_285/B 0.01fF
C5893 OR2X1_LOC_154/A OR2X1_LOC_175/B 0.02fF
C5894 AND2X1_LOC_139/a_8_24# OR2X1_LOC_26/Y 0.01fF
C5895 OR2X1_LOC_101/a_8_216# OR2X1_LOC_520/Y 0.02fF
C5896 OR2X1_LOC_74/A OR2X1_LOC_59/Y 0.31fF
C5897 AND2X1_LOC_141/A AND2X1_LOC_361/A 0.04fF
C5898 OR2X1_LOC_160/A OR2X1_LOC_799/A 0.05fF
C5899 OR2X1_LOC_354/A OR2X1_LOC_269/B 0.05fF
C5900 AND2X1_LOC_798/Y AND2X1_LOC_436/Y 0.00fF
C5901 OR2X1_LOC_61/Y OR2X1_LOC_358/B 0.04fF
C5902 D_INPUT_7 AND2X1_LOC_50/a_8_24# 0.12fF
C5903 OR2X1_LOC_502/A OR2X1_LOC_753/A 0.05fF
C5904 AND2X1_LOC_711/A OR2X1_LOC_295/a_8_216# 0.47fF
C5905 OR2X1_LOC_377/A OR2X1_LOC_404/a_8_216# 0.04fF
C5906 OR2X1_LOC_235/B OR2X1_LOC_278/a_36_216# 0.00fF
C5907 OR2X1_LOC_434/a_8_216# AND2X1_LOC_3/Y 0.04fF
C5908 OR2X1_LOC_46/A AND2X1_LOC_411/a_8_24# 0.04fF
C5909 AND2X1_LOC_51/Y OR2X1_LOC_803/A 0.02fF
C5910 AND2X1_LOC_196/a_36_24# OR2X1_LOC_59/Y 0.00fF
C5911 AND2X1_LOC_64/Y OR2X1_LOC_804/A 0.07fF
C5912 AND2X1_LOC_22/Y OR2X1_LOC_845/A 0.05fF
C5913 AND2X1_LOC_363/a_8_24# OR2X1_LOC_417/A 0.02fF
C5914 AND2X1_LOC_784/A AND2X1_LOC_364/A 0.08fF
C5915 AND2X1_LOC_181/Y OR2X1_LOC_417/A 0.02fF
C5916 AND2X1_LOC_59/Y OR2X1_LOC_805/A 0.15fF
C5917 OR2X1_LOC_600/A OR2X1_LOC_295/Y 0.01fF
C5918 AND2X1_LOC_851/B AND2X1_LOC_786/Y 0.07fF
C5919 OR2X1_LOC_147/a_8_216# OR2X1_LOC_147/B 0.10fF
C5920 OR2X1_LOC_242/a_8_216# AND2X1_LOC_51/Y 0.01fF
C5921 AND2X1_LOC_850/Y AND2X1_LOC_288/a_8_24# 0.20fF
C5922 OR2X1_LOC_574/A OR2X1_LOC_575/A 0.01fF
C5923 OR2X1_LOC_520/Y OR2X1_LOC_130/A 0.05fF
C5924 AND2X1_LOC_720/a_8_24# OR2X1_LOC_669/Y 0.06fF
C5925 OR2X1_LOC_114/a_8_216# OR2X1_LOC_404/Y 0.02fF
C5926 OR2X1_LOC_382/Y OR2X1_LOC_481/A 0.41fF
C5927 AND2X1_LOC_211/B AND2X1_LOC_841/B 0.07fF
C5928 AND2X1_LOC_101/B OR2X1_LOC_18/Y 0.71fF
C5929 AND2X1_LOC_1/Y AND2X1_LOC_3/a_8_24# 0.09fF
C5930 OR2X1_LOC_653/Y AND2X1_LOC_3/Y 0.07fF
C5931 OR2X1_LOC_529/Y OR2X1_LOC_427/A 0.04fF
C5932 OR2X1_LOC_600/A OR2X1_LOC_80/a_8_216# 0.01fF
C5933 OR2X1_LOC_91/Y OR2X1_LOC_6/A 0.03fF
C5934 AND2X1_LOC_795/Y OR2X1_LOC_373/a_8_216# 0.11fF
C5935 VDD OR2X1_LOC_434/A -0.00fF
C5936 AND2X1_LOC_259/Y OR2X1_LOC_257/a_8_216# 0.01fF
C5937 AND2X1_LOC_817/B AND2X1_LOC_817/a_8_24# 0.20fF
C5938 AND2X1_LOC_702/Y AND2X1_LOC_302/a_8_24# 0.01fF
C5939 AND2X1_LOC_367/A AND2X1_LOC_514/Y 0.03fF
C5940 AND2X1_LOC_537/a_8_24# OR2X1_LOC_95/Y 0.01fF
C5941 OR2X1_LOC_602/Y AND2X1_LOC_47/Y 0.15fF
C5942 OR2X1_LOC_151/A OR2X1_LOC_786/Y 0.03fF
C5943 OR2X1_LOC_703/Y OR2X1_LOC_317/B 0.00fF
C5944 OR2X1_LOC_89/A AND2X1_LOC_656/a_36_24# 0.00fF
C5945 OR2X1_LOC_11/Y OR2X1_LOC_585/A 0.04fF
C5946 OR2X1_LOC_305/a_36_216# OR2X1_LOC_305/Y 0.00fF
C5947 AND2X1_LOC_339/a_8_24# OR2X1_LOC_316/Y 0.01fF
C5948 OR2X1_LOC_244/A OR2X1_LOC_78/A 0.07fF
C5949 AND2X1_LOC_356/B AND2X1_LOC_365/A 0.01fF
C5950 OR2X1_LOC_595/Y AND2X1_LOC_786/Y 0.02fF
C5951 AND2X1_LOC_193/a_36_24# OR2X1_LOC_43/A 0.00fF
C5952 OR2X1_LOC_70/Y AND2X1_LOC_76/a_36_24# 0.01fF
C5953 AND2X1_LOC_502/a_8_24# OR2X1_LOC_485/A 0.02fF
C5954 OR2X1_LOC_62/B AND2X1_LOC_647/a_8_24# 0.01fF
C5955 AND2X1_LOC_235/a_8_24# OR2X1_LOC_71/A 0.01fF
C5956 OR2X1_LOC_820/Y AND2X1_LOC_847/Y 0.92fF
C5957 OR2X1_LOC_22/Y OR2X1_LOC_275/Y 0.14fF
C5958 AND2X1_LOC_54/a_8_24# INPUT_1 0.08fF
C5959 AND2X1_LOC_727/A OR2X1_LOC_594/a_36_216# 0.00fF
C5960 OR2X1_LOC_30/a_36_216# OR2X1_LOC_17/Y 0.00fF
C5961 OR2X1_LOC_831/a_36_216# OR2X1_LOC_155/A 0.00fF
C5962 AND2X1_LOC_12/Y AND2X1_LOC_425/a_8_24# 0.01fF
C5963 AND2X1_LOC_550/a_8_24# OR2X1_LOC_47/Y 0.01fF
C5964 OR2X1_LOC_22/Y AND2X1_LOC_654/B 2.15fF
C5965 AND2X1_LOC_306/a_8_24# AND2X1_LOC_47/Y 0.07fF
C5966 OR2X1_LOC_757/A AND2X1_LOC_866/A 0.02fF
C5967 OR2X1_LOC_690/A OR2X1_LOC_585/A 0.03fF
C5968 GATE_366 OR2X1_LOC_485/A 0.01fF
C5969 OR2X1_LOC_463/a_8_216# AND2X1_LOC_3/Y 0.01fF
C5970 AND2X1_LOC_569/A OR2X1_LOC_189/Y 0.32fF
C5971 AND2X1_LOC_356/B OR2X1_LOC_43/A 0.01fF
C5972 AND2X1_LOC_729/B AND2X1_LOC_655/A 0.44fF
C5973 OR2X1_LOC_165/Y OR2X1_LOC_417/A 0.02fF
C5974 AND2X1_LOC_784/A OR2X1_LOC_3/Y 0.41fF
C5975 AND2X1_LOC_564/a_8_24# AND2X1_LOC_711/Y 0.03fF
C5976 AND2X1_LOC_784/A AND2X1_LOC_568/a_8_24# 0.03fF
C5977 OR2X1_LOC_815/a_8_216# AND2X1_LOC_793/Y 0.04fF
C5978 OR2X1_LOC_763/Y OR2X1_LOC_764/Y 0.21fF
C5979 OR2X1_LOC_299/Y OR2X1_LOC_52/B 0.13fF
C5980 OR2X1_LOC_479/Y OR2X1_LOC_469/a_36_216# 0.02fF
C5981 OR2X1_LOC_485/A OR2X1_LOC_312/Y 0.00fF
C5982 AND2X1_LOC_727/A AND2X1_LOC_652/a_8_24# 0.01fF
C5983 OR2X1_LOC_646/A OR2X1_LOC_647/B 0.01fF
C5984 OR2X1_LOC_496/Y AND2X1_LOC_578/A 0.01fF
C5985 OR2X1_LOC_675/a_36_216# OR2X1_LOC_76/Y 0.00fF
C5986 OR2X1_LOC_532/B OR2X1_LOC_733/a_8_216# 0.01fF
C5987 OR2X1_LOC_378/Y AND2X1_LOC_459/a_8_24# 0.01fF
C5988 OR2X1_LOC_750/a_8_216# OR2X1_LOC_161/A 0.07fF
C5989 OR2X1_LOC_377/A OR2X1_LOC_403/a_36_216# 0.01fF
C5990 AND2X1_LOC_365/A OR2X1_LOC_22/Y 0.07fF
C5991 OR2X1_LOC_435/B OR2X1_LOC_112/B 0.04fF
C5992 AND2X1_LOC_569/A OR2X1_LOC_527/Y 0.00fF
C5993 AND2X1_LOC_711/Y OR2X1_LOC_757/a_8_216# 0.01fF
C5994 OR2X1_LOC_18/Y OR2X1_LOC_226/a_8_216# 0.09fF
C5995 OR2X1_LOC_160/A AND2X1_LOC_698/a_36_24# 0.01fF
C5996 OR2X1_LOC_261/A OR2X1_LOC_820/B -0.00fF
C5997 AND2X1_LOC_91/B OR2X1_LOC_532/Y 0.01fF
C5998 OR2X1_LOC_402/Y OR2X1_LOC_532/B 0.16fF
C5999 OR2X1_LOC_92/Y OR2X1_LOC_760/Y 0.03fF
C6000 OR2X1_LOC_605/a_8_216# OR2X1_LOC_787/Y 0.01fF
C6001 OR2X1_LOC_64/Y OR2X1_LOC_585/A 0.88fF
C6002 OR2X1_LOC_70/Y OR2X1_LOC_490/Y 0.09fF
C6003 OR2X1_LOC_70/Y OR2X1_LOC_74/A 0.17fF
C6004 AND2X1_LOC_658/B AND2X1_LOC_222/Y 0.03fF
C6005 OR2X1_LOC_3/Y OR2X1_LOC_481/Y 0.01fF
C6006 AND2X1_LOC_1/Y AND2X1_LOC_21/Y 0.90fF
C6007 OR2X1_LOC_43/A OR2X1_LOC_22/Y 0.21fF
C6008 AND2X1_LOC_56/B OR2X1_LOC_471/Y 0.06fF
C6009 AND2X1_LOC_345/a_8_24# AND2X1_LOC_663/B 0.01fF
C6010 OR2X1_LOC_596/A OR2X1_LOC_317/B 0.07fF
C6011 AND2X1_LOC_348/A AND2X1_LOC_721/A 0.00fF
C6012 OR2X1_LOC_404/Y AND2X1_LOC_42/B 0.03fF
C6013 AND2X1_LOC_694/a_8_24# OR2X1_LOC_449/B 0.01fF
C6014 OR2X1_LOC_139/A AND2X1_LOC_36/Y 0.04fF
C6015 AND2X1_LOC_180/a_8_24# OR2X1_LOC_437/A 0.04fF
C6016 OR2X1_LOC_742/B OR2X1_LOC_191/a_36_216# 0.02fF
C6017 OR2X1_LOC_352/A OR2X1_LOC_365/B 0.00fF
C6018 OR2X1_LOC_483/a_36_216# OR2X1_LOC_532/B 0.03fF
C6019 D_INPUT_0 AND2X1_LOC_472/B 0.03fF
C6020 OR2X1_LOC_833/B OR2X1_LOC_270/Y 0.01fF
C6021 OR2X1_LOC_89/A AND2X1_LOC_814/a_8_24# 0.01fF
C6022 AND2X1_LOC_8/Y OR2X1_LOC_655/B 0.05fF
C6023 OR2X1_LOC_287/B OR2X1_LOC_814/A 0.06fF
C6024 AND2X1_LOC_212/Y OR2X1_LOC_142/Y 0.07fF
C6025 AND2X1_LOC_44/Y OR2X1_LOC_500/a_8_216# 0.01fF
C6026 OR2X1_LOC_32/B OR2X1_LOC_47/Y 0.10fF
C6027 OR2X1_LOC_715/A OR2X1_LOC_513/Y 0.15fF
C6028 OR2X1_LOC_3/Y AND2X1_LOC_639/A 0.02fF
C6029 AND2X1_LOC_359/B AND2X1_LOC_866/A 0.08fF
C6030 D_INPUT_3 OR2X1_LOC_6/A 0.08fF
C6031 OR2X1_LOC_520/Y AND2X1_LOC_88/Y 0.14fF
C6032 OR2X1_LOC_254/B OR2X1_LOC_270/Y 0.01fF
C6033 AND2X1_LOC_319/A AND2X1_LOC_798/A 0.17fF
C6034 OR2X1_LOC_66/A OR2X1_LOC_140/Y 0.02fF
C6035 OR2X1_LOC_504/Y OR2X1_LOC_74/A 0.19fF
C6036 OR2X1_LOC_487/Y OR2X1_LOC_71/Y 0.01fF
C6037 OR2X1_LOC_22/Y OR2X1_LOC_60/a_8_216# 0.01fF
C6038 AND2X1_LOC_357/a_8_24# AND2X1_LOC_222/Y 0.01fF
C6039 AND2X1_LOC_91/B OR2X1_LOC_266/A 0.22fF
C6040 OR2X1_LOC_76/A OR2X1_LOC_814/A 0.07fF
C6041 OR2X1_LOC_85/A AND2X1_LOC_203/Y 0.01fF
C6042 AND2X1_LOC_43/B AND2X1_LOC_679/a_8_24# 0.01fF
C6043 OR2X1_LOC_121/B OR2X1_LOC_335/B 0.00fF
C6044 OR2X1_LOC_582/Y AND2X1_LOC_639/A 0.87fF
C6045 OR2X1_LOC_86/Y OR2X1_LOC_67/Y 0.01fF
C6046 AND2X1_LOC_537/Y AND2X1_LOC_539/a_8_24# 0.09fF
C6047 AND2X1_LOC_557/a_8_24# D_INPUT_3 0.16fF
C6048 AND2X1_LOC_578/A AND2X1_LOC_851/B 0.08fF
C6049 AND2X1_LOC_456/Y OR2X1_LOC_184/Y 0.60fF
C6050 OR2X1_LOC_19/B D_INPUT_0 0.81fF
C6051 AND2X1_LOC_315/a_8_24# AND2X1_LOC_31/Y 0.01fF
C6052 AND2X1_LOC_721/Y AND2X1_LOC_464/A 0.00fF
C6053 OR2X1_LOC_47/Y OR2X1_LOC_371/Y 0.04fF
C6054 AND2X1_LOC_179/a_8_24# AND2X1_LOC_36/Y 0.08fF
C6055 OR2X1_LOC_646/a_36_216# D_INPUT_1 0.02fF
C6056 AND2X1_LOC_831/Y OR2X1_LOC_416/Y 0.01fF
C6057 OR2X1_LOC_49/A AND2X1_LOC_44/Y 0.84fF
C6058 AND2X1_LOC_773/Y AND2X1_LOC_774/A 0.01fF
C6059 OR2X1_LOC_437/Y OR2X1_LOC_74/A -0.02fF
C6060 OR2X1_LOC_64/Y AND2X1_LOC_645/a_8_24# 0.01fF
C6061 AND2X1_LOC_18/Y OR2X1_LOC_140/B 0.03fF
C6062 AND2X1_LOC_41/A AND2X1_LOC_239/a_8_24# 0.01fF
C6063 OR2X1_LOC_161/A OR2X1_LOC_546/A 0.01fF
C6064 OR2X1_LOC_97/A OR2X1_LOC_439/B 0.02fF
C6065 OR2X1_LOC_78/B OR2X1_LOC_319/Y 0.00fF
C6066 OR2X1_LOC_108/Y AND2X1_LOC_465/A 0.15fF
C6067 OR2X1_LOC_436/Y OR2X1_LOC_814/A 0.04fF
C6068 AND2X1_LOC_47/Y OR2X1_LOC_602/B 0.05fF
C6069 OR2X1_LOC_596/A AND2X1_LOC_44/Y 0.20fF
C6070 AND2X1_LOC_362/B OR2X1_LOC_428/A 0.06fF
C6071 OR2X1_LOC_160/A OR2X1_LOC_446/B 0.21fF
C6072 AND2X1_LOC_476/Y OR2X1_LOC_428/A 2.04fF
C6073 OR2X1_LOC_461/A OR2X1_LOC_68/B 0.04fF
C6074 OR2X1_LOC_617/Y AND2X1_LOC_793/Y 0.01fF
C6075 OR2X1_LOC_3/Y AND2X1_LOC_643/a_8_24# 0.07fF
C6076 OR2X1_LOC_105/Y OR2X1_LOC_579/A 0.24fF
C6077 AND2X1_LOC_729/B OR2X1_LOC_599/Y 0.03fF
C6078 OR2X1_LOC_550/a_8_216# OR2X1_LOC_550/A 0.39fF
C6079 OR2X1_LOC_508/A AND2X1_LOC_239/a_8_24# 0.06fF
C6080 AND2X1_LOC_53/Y OR2X1_LOC_197/A 0.03fF
C6081 OR2X1_LOC_864/A OR2X1_LOC_68/B 0.10fF
C6082 AND2X1_LOC_130/a_8_24# OR2X1_LOC_12/Y 0.07fF
C6083 AND2X1_LOC_687/Y AND2X1_LOC_648/B 0.02fF
C6084 OR2X1_LOC_415/A OR2X1_LOC_396/Y 0.09fF
C6085 OR2X1_LOC_70/Y AND2X1_LOC_647/Y 0.02fF
C6086 OR2X1_LOC_160/A OR2X1_LOC_728/a_8_216# 0.02fF
C6087 AND2X1_LOC_362/B OR2X1_LOC_595/A 0.31fF
C6088 OR2X1_LOC_83/A OR2X1_LOC_80/A 0.29fF
C6089 OR2X1_LOC_596/A OR2X1_LOC_514/a_8_216# 0.01fF
C6090 OR2X1_LOC_176/a_8_216# OR2X1_LOC_51/Y 0.14fF
C6091 OR2X1_LOC_633/B OR2X1_LOC_68/B 0.00fF
C6092 VDD OR2X1_LOC_162/A -0.00fF
C6093 AND2X1_LOC_95/Y OR2X1_LOC_523/A 0.01fF
C6094 OR2X1_LOC_49/A OR2X1_LOC_600/A 0.59fF
C6095 D_INPUT_0 OR2X1_LOC_838/B 0.03fF
C6096 AND2X1_LOC_387/a_36_24# AND2X1_LOC_44/Y 0.01fF
C6097 AND2X1_LOC_188/a_8_24# OR2X1_LOC_816/A 0.00fF
C6098 AND2X1_LOC_64/Y AND2X1_LOC_65/a_8_24# 0.11fF
C6099 AND2X1_LOC_580/A OR2X1_LOC_437/A 0.07fF
C6100 OR2X1_LOC_3/Y OR2X1_LOC_88/Y 0.03fF
C6101 AND2X1_LOC_560/a_8_24# OR2X1_LOC_103/Y 0.24fF
C6102 AND2X1_LOC_459/a_8_24# OR2X1_LOC_378/A 0.04fF
C6103 OR2X1_LOC_3/Y OR2X1_LOC_172/Y 0.27fF
C6104 OR2X1_LOC_323/A OR2X1_LOC_164/Y 0.02fF
C6105 OR2X1_LOC_696/A AND2X1_LOC_113/a_8_24# 0.01fF
C6106 OR2X1_LOC_45/B OR2X1_LOC_56/A 0.82fF
C6107 AND2X1_LOC_814/a_36_24# AND2X1_LOC_624/B 0.01fF
C6108 D_INPUT_2 D_INPUT_3 0.28fF
C6109 AND2X1_LOC_839/A D_INPUT_1 0.00fF
C6110 OR2X1_LOC_70/A OR2X1_LOC_762/a_36_216# 0.00fF
C6111 OR2X1_LOC_66/A OR2X1_LOC_548/a_36_216# 0.02fF
C6112 OR2X1_LOC_248/a_36_216# OR2X1_LOC_13/B 0.00fF
C6113 OR2X1_LOC_66/A OR2X1_LOC_390/A 0.09fF
C6114 OR2X1_LOC_203/Y OR2X1_LOC_777/B 0.07fF
C6115 AND2X1_LOC_525/a_8_24# OR2X1_LOC_546/A 0.02fF
C6116 AND2X1_LOC_707/Y OR2X1_LOC_421/a_8_216# 0.03fF
C6117 OR2X1_LOC_62/A OR2X1_LOC_673/A 0.04fF
C6118 AND2X1_LOC_91/B OR2X1_LOC_400/a_8_216# 0.05fF
C6119 AND2X1_LOC_64/Y OR2X1_LOC_403/A 0.01fF
C6120 OR2X1_LOC_97/A AND2X1_LOC_41/A 0.03fF
C6121 INPUT_4 OR2X1_LOC_386/a_8_216# 0.07fF
C6122 OR2X1_LOC_442/Y AND2X1_LOC_212/Y 0.03fF
C6123 OR2X1_LOC_820/a_36_216# OR2X1_LOC_600/A 0.00fF
C6124 OR2X1_LOC_147/B OR2X1_LOC_562/A 0.03fF
C6125 OR2X1_LOC_325/B AND2X1_LOC_110/Y 0.01fF
C6126 AND2X1_LOC_571/B AND2X1_LOC_572/Y 0.02fF
C6127 OR2X1_LOC_56/A OR2X1_LOC_382/A 0.10fF
C6128 OR2X1_LOC_421/A OR2X1_LOC_597/A 0.01fF
C6129 OR2X1_LOC_623/B AND2X1_LOC_7/B 0.07fF
C6130 OR2X1_LOC_485/A OR2X1_LOC_13/B 0.28fF
C6131 OR2X1_LOC_53/Y OR2X1_LOC_59/a_8_216# 0.40fF
C6132 AND2X1_LOC_51/Y OR2X1_LOC_546/A 0.02fF
C6133 OR2X1_LOC_135/Y AND2X1_LOC_303/a_8_24# 0.15fF
C6134 OR2X1_LOC_690/Y AND2X1_LOC_194/Y 0.05fF
C6135 AND2X1_LOC_724/Y AND2X1_LOC_732/B 0.01fF
C6136 AND2X1_LOC_64/Y OR2X1_LOC_447/a_8_216# 0.09fF
C6137 AND2X1_LOC_22/Y AND2X1_LOC_328/a_8_24# 0.01fF
C6138 OR2X1_LOC_517/A OR2X1_LOC_12/Y 0.13fF
C6139 OR2X1_LOC_324/a_8_216# AND2X1_LOC_44/Y 0.02fF
C6140 OR2X1_LOC_500/A OR2X1_LOC_140/B 0.01fF
C6141 VDD OR2X1_LOC_741/Y 0.06fF
C6142 D_INPUT_4 INPUT_7 0.02fF
C6143 OR2X1_LOC_757/A OR2X1_LOC_40/Y 0.07fF
C6144 VDD AND2X1_LOC_658/Y 0.26fF
C6145 AND2X1_LOC_64/Y OR2X1_LOC_130/A 0.03fF
C6146 VDD OR2X1_LOC_743/a_8_216# 0.21fF
C6147 OR2X1_LOC_179/a_8_216# OR2X1_LOC_158/A 0.01fF
C6148 OR2X1_LOC_59/Y AND2X1_LOC_860/A 0.17fF
C6149 OR2X1_LOC_114/a_8_216# OR2X1_LOC_362/A 0.02fF
C6150 OR2X1_LOC_59/Y OR2X1_LOC_626/Y 0.08fF
C6151 OR2X1_LOC_6/A OR2X1_LOC_171/Y 0.02fF
C6152 OR2X1_LOC_135/a_8_216# OR2X1_LOC_427/A 0.02fF
C6153 OR2X1_LOC_738/B OR2X1_LOC_738/a_8_216# 0.39fF
C6154 OR2X1_LOC_640/Y AND2X1_LOC_92/Y 0.01fF
C6155 OR2X1_LOC_137/a_8_216# OR2X1_LOC_160/B 0.05fF
C6156 AND2X1_LOC_714/B OR2X1_LOC_92/Y 0.04fF
C6157 AND2X1_LOC_44/a_36_24# INPUT_6 0.00fF
C6158 OR2X1_LOC_97/A OR2X1_LOC_662/A 0.01fF
C6159 OR2X1_LOC_310/Y AND2X1_LOC_335/Y 0.79fF
C6160 OR2X1_LOC_406/Y OR2X1_LOC_406/a_8_216# 0.01fF
C6161 OR2X1_LOC_191/a_8_216# OR2X1_LOC_192/A -0.00fF
C6162 AND2X1_LOC_859/a_8_24# AND2X1_LOC_287/B 0.01fF
C6163 AND2X1_LOC_702/a_8_24# OR2X1_LOC_135/Y 0.01fF
C6164 OR2X1_LOC_813/Y OR2X1_LOC_86/A 0.02fF
C6165 OR2X1_LOC_47/Y AND2X1_LOC_222/Y 0.05fF
C6166 VDD AND2X1_LOC_734/Y 0.05fF
C6167 OR2X1_LOC_87/A OR2X1_LOC_352/a_36_216# 0.00fF
C6168 AND2X1_LOC_763/a_8_24# INPUT_0 0.04fF
C6169 OR2X1_LOC_52/B AND2X1_LOC_780/a_36_24# 0.01fF
C6170 OR2X1_LOC_292/a_8_216# OR2X1_LOC_56/A 0.02fF
C6171 AND2X1_LOC_663/B AND2X1_LOC_792/B 0.01fF
C6172 AND2X1_LOC_70/Y OR2X1_LOC_663/A 0.03fF
C6173 OR2X1_LOC_113/a_8_216# OR2X1_LOC_643/A 0.01fF
C6174 AND2X1_LOC_722/A AND2X1_LOC_436/Y 0.03fF
C6175 OR2X1_LOC_175/Y OR2X1_LOC_214/a_8_216# 0.01fF
C6176 OR2X1_LOC_643/A OR2X1_LOC_474/B 0.02fF
C6177 OR2X1_LOC_154/A OR2X1_LOC_389/a_8_216# 0.01fF
C6178 OR2X1_LOC_51/Y OR2X1_LOC_251/a_36_216# 0.02fF
C6179 OR2X1_LOC_87/B AND2X1_LOC_44/Y 0.18fF
C6180 OR2X1_LOC_467/A OR2X1_LOC_477/Y 0.16fF
C6181 AND2X1_LOC_508/A AND2X1_LOC_663/A 0.05fF
C6182 AND2X1_LOC_712/Y OR2X1_LOC_619/Y 0.09fF
C6183 OR2X1_LOC_744/A AND2X1_LOC_850/A 0.24fF
C6184 AND2X1_LOC_539/Y AND2X1_LOC_337/B 0.01fF
C6185 OR2X1_LOC_307/B OR2X1_LOC_78/A 0.01fF
C6186 OR2X1_LOC_589/A OR2X1_LOC_39/A 0.02fF
C6187 AND2X1_LOC_802/B OR2X1_LOC_312/Y 0.03fF
C6188 OR2X1_LOC_268/a_8_216# OR2X1_LOC_268/Y 0.01fF
C6189 AND2X1_LOC_41/A OR2X1_LOC_541/A 0.09fF
C6190 OR2X1_LOC_372/Y AND2X1_LOC_786/Y 0.04fF
C6191 OR2X1_LOC_364/B OR2X1_LOC_364/A 0.18fF
C6192 OR2X1_LOC_3/Y OR2X1_LOC_397/Y 0.34fF
C6193 OR2X1_LOC_600/A AND2X1_LOC_805/Y 0.01fF
C6194 D_INPUT_5 OR2X1_LOC_25/Y 0.05fF
C6195 OR2X1_LOC_51/Y OR2X1_LOC_46/a_8_216# 0.01fF
C6196 OR2X1_LOC_709/A OR2X1_LOC_185/Y 0.03fF
C6197 INPUT_0 AND2X1_LOC_857/Y 0.03fF
C6198 OR2X1_LOC_648/A OR2X1_LOC_61/B 0.20fF
C6199 OR2X1_LOC_203/Y OR2X1_LOC_344/A -0.01fF
C6200 VDD OR2X1_LOC_109/a_8_216# 0.21fF
C6201 AND2X1_LOC_231/Y AND2X1_LOC_211/B 0.26fF
C6202 AND2X1_LOC_562/B OR2X1_LOC_698/a_36_216# 0.00fF
C6203 AND2X1_LOC_807/B AND2X1_LOC_807/a_8_24# 0.01fF
C6204 AND2X1_LOC_326/B AND2X1_LOC_662/B 0.03fF
C6205 AND2X1_LOC_364/a_8_24# AND2X1_LOC_211/B 0.01fF
C6206 OR2X1_LOC_532/B OR2X1_LOC_593/B 0.03fF
C6207 AND2X1_LOC_723/Y OR2X1_LOC_164/Y 0.14fF
C6208 AND2X1_LOC_456/B OR2X1_LOC_256/Y 0.23fF
C6209 OR2X1_LOC_318/B OR2X1_LOC_228/Y 0.01fF
C6210 OR2X1_LOC_327/a_8_216# OR2X1_LOC_78/A 0.02fF
C6211 AND2X1_LOC_155/Y OR2X1_LOC_744/a_8_216# 0.49fF
C6212 OR2X1_LOC_574/A OR2X1_LOC_161/B 0.30fF
C6213 OR2X1_LOC_208/A OR2X1_LOC_19/B 0.01fF
C6214 OR2X1_LOC_494/A OR2X1_LOC_481/A 0.31fF
C6215 OR2X1_LOC_45/B AND2X1_LOC_641/Y 0.05fF
C6216 OR2X1_LOC_696/A OR2X1_LOC_62/B 0.01fF
C6217 AND2X1_LOC_784/A AND2X1_LOC_477/Y 0.02fF
C6218 AND2X1_LOC_141/a_8_24# OR2X1_LOC_118/Y 0.01fF
C6219 OR2X1_LOC_813/a_8_216# OR2X1_LOC_85/A 0.05fF
C6220 AND2X1_LOC_363/Y AND2X1_LOC_848/Y 0.08fF
C6221 AND2X1_LOC_564/B OR2X1_LOC_64/Y 0.08fF
C6222 OR2X1_LOC_18/Y AND2X1_LOC_663/A 0.05fF
C6223 OR2X1_LOC_614/Y AND2X1_LOC_683/a_8_24# 0.23fF
C6224 AND2X1_LOC_64/Y OR2X1_LOC_62/B 0.10fF
C6225 OR2X1_LOC_746/Y AND2X1_LOC_781/a_8_24# 0.00fF
C6226 OR2X1_LOC_538/a_8_216# OR2X1_LOC_856/B 0.06fF
C6227 OR2X1_LOC_158/A AND2X1_LOC_34/a_8_24# 0.03fF
C6228 OR2X1_LOC_457/B OR2X1_LOC_787/B 0.14fF
C6229 OR2X1_LOC_431/a_8_216# OR2X1_LOC_428/A 0.04fF
C6230 OR2X1_LOC_402/Y OR2X1_LOC_78/a_36_216# 0.00fF
C6231 VDD AND2X1_LOC_817/a_8_24# -0.00fF
C6232 OR2X1_LOC_40/Y OR2X1_LOC_626/a_8_216# 0.02fF
C6233 AND2X1_LOC_729/Y OR2X1_LOC_329/B 0.43fF
C6234 OR2X1_LOC_364/A AND2X1_LOC_70/Y 0.49fF
C6235 AND2X1_LOC_186/a_8_24# AND2X1_LOC_548/Y 0.00fF
C6236 OR2X1_LOC_185/Y AND2X1_LOC_70/Y 0.04fF
C6237 OR2X1_LOC_814/A OR2X1_LOC_722/B 0.01fF
C6238 AND2X1_LOC_2/a_8_24# AND2X1_LOC_11/Y 0.22fF
C6239 OR2X1_LOC_506/a_8_216# OR2X1_LOC_532/B 0.05fF
C6240 OR2X1_LOC_756/B OR2X1_LOC_456/a_8_216# 0.01fF
C6241 OR2X1_LOC_169/a_8_216# AND2X1_LOC_92/Y 0.02fF
C6242 VDD OR2X1_LOC_24/a_8_216# 0.21fF
C6243 VDD OR2X1_LOC_210/B 0.00fF
C6244 AND2X1_LOC_662/B AND2X1_LOC_276/a_8_24# 0.01fF
C6245 OR2X1_LOC_858/A OR2X1_LOC_87/A 0.03fF
C6246 OR2X1_LOC_9/Y AND2X1_LOC_42/B 0.01fF
C6247 OR2X1_LOC_678/Y OR2X1_LOC_375/A 0.01fF
C6248 OR2X1_LOC_59/Y AND2X1_LOC_287/Y 0.03fF
C6249 OR2X1_LOC_468/Y AND2X1_LOC_92/Y 0.03fF
C6250 OR2X1_LOC_89/A AND2X1_LOC_614/a_8_24# 0.01fF
C6251 AND2X1_LOC_259/Y OR2X1_LOC_600/A 1.28fF
C6252 AND2X1_LOC_42/B OR2X1_LOC_362/A 0.03fF
C6253 OR2X1_LOC_40/Y AND2X1_LOC_639/a_8_24# 0.01fF
C6254 OR2X1_LOC_275/Y OR2X1_LOC_39/A 0.04fF
C6255 OR2X1_LOC_160/A OR2X1_LOC_736/A 0.25fF
C6256 AND2X1_LOC_576/Y AND2X1_LOC_858/B 0.10fF
C6257 AND2X1_LOC_810/A AND2X1_LOC_514/Y 0.05fF
C6258 OR2X1_LOC_92/Y OR2X1_LOC_71/a_36_216# 0.00fF
C6259 OR2X1_LOC_649/a_36_216# AND2X1_LOC_44/Y 0.01fF
C6260 AND2X1_LOC_784/A OR2X1_LOC_329/B 0.07fF
C6261 AND2X1_LOC_564/B OR2X1_LOC_417/A 0.07fF
C6262 OR2X1_LOC_134/Y OR2X1_LOC_95/Y 0.21fF
C6263 OR2X1_LOC_287/B OR2X1_LOC_244/Y 0.02fF
C6264 AND2X1_LOC_866/B OR2X1_LOC_39/A 0.18fF
C6265 OR2X1_LOC_187/a_8_216# OR2X1_LOC_680/A 0.01fF
C6266 OR2X1_LOC_656/Y OR2X1_LOC_130/A 0.16fF
C6267 AND2X1_LOC_59/Y AND2X1_LOC_331/a_8_24# 0.02fF
C6268 OR2X1_LOC_643/A OR2X1_LOC_658/a_8_216# 0.01fF
C6269 AND2X1_LOC_711/Y OR2X1_LOC_626/Y 0.03fF
C6270 AND2X1_LOC_508/a_36_24# AND2X1_LOC_474/Y 0.00fF
C6271 OR2X1_LOC_620/Y OR2X1_LOC_624/A 0.52fF
C6272 OR2X1_LOC_495/Y OR2X1_LOC_39/A 0.07fF
C6273 AND2X1_LOC_259/Y AND2X1_LOC_296/a_8_24# 0.01fF
C6274 INPUT_4 D_INPUT_4 0.06fF
C6275 AND2X1_LOC_719/a_36_24# AND2X1_LOC_658/A 0.01fF
C6276 OR2X1_LOC_585/A OR2X1_LOC_232/Y 0.01fF
C6277 AND2X1_LOC_772/B AND2X1_LOC_554/B 0.00fF
C6278 AND2X1_LOC_64/Y AND2X1_LOC_88/Y 0.00fF
C6279 AND2X1_LOC_701/a_8_24# AND2X1_LOC_526/a_8_24# 0.23fF
C6280 OR2X1_LOC_811/A OR2X1_LOC_375/A 0.01fF
C6281 AND2X1_LOC_677/a_8_24# OR2X1_LOC_307/A 0.10fF
C6282 AND2X1_LOC_700/a_8_24# AND2X1_LOC_51/Y 0.04fF
C6283 OR2X1_LOC_598/Y OR2X1_LOC_19/B 0.00fF
C6284 AND2X1_LOC_486/Y OR2X1_LOC_497/Y 0.10fF
C6285 OR2X1_LOC_525/Y AND2X1_LOC_834/a_8_24# 0.02fF
C6286 AND2X1_LOC_858/a_8_24# OR2X1_LOC_39/A 0.01fF
C6287 OR2X1_LOC_452/A AND2X1_LOC_425/Y 0.02fF
C6288 OR2X1_LOC_6/B AND2X1_LOC_667/a_8_24# 0.04fF
C6289 AND2X1_LOC_86/a_8_24# OR2X1_LOC_62/B 0.01fF
C6290 AND2X1_LOC_95/Y OR2X1_LOC_462/B 0.72fF
C6291 AND2X1_LOC_578/A OR2X1_LOC_674/a_8_216# 0.03fF
C6292 AND2X1_LOC_51/A D_INPUT_4 0.05fF
C6293 AND2X1_LOC_583/a_8_24# OR2X1_LOC_636/B 0.02fF
C6294 OR2X1_LOC_154/A OR2X1_LOC_624/A 0.47fF
C6295 AND2X1_LOC_40/Y OR2X1_LOC_593/A 0.01fF
C6296 OR2X1_LOC_750/A OR2X1_LOC_66/A 0.03fF
C6297 OR2X1_LOC_633/Y OR2X1_LOC_462/B 0.00fF
C6298 OR2X1_LOC_604/A OR2X1_LOC_77/a_36_216# 0.01fF
C6299 AND2X1_LOC_824/B AND2X1_LOC_824/a_8_24# 0.01fF
C6300 AND2X1_LOC_572/A OR2X1_LOC_67/A 0.01fF
C6301 OR2X1_LOC_744/A AND2X1_LOC_523/Y 0.07fF
C6302 OR2X1_LOC_703/B OR2X1_LOC_169/B 0.24fF
C6303 OR2X1_LOC_160/B OR2X1_LOC_814/A 17.61fF
C6304 OR2X1_LOC_272/Y OR2X1_LOC_517/A 0.18fF
C6305 AND2X1_LOC_110/Y D_INPUT_0 0.03fF
C6306 OR2X1_LOC_756/B OR2X1_LOC_35/B 0.01fF
C6307 AND2X1_LOC_99/A OR2X1_LOC_26/Y 0.02fF
C6308 AND2X1_LOC_576/Y AND2X1_LOC_573/A 0.02fF
C6309 OR2X1_LOC_158/A AND2X1_LOC_859/B 0.01fF
C6310 OR2X1_LOC_474/Y AND2X1_LOC_42/B 0.22fF
C6311 AND2X1_LOC_661/A OR2X1_LOC_619/Y 0.07fF
C6312 OR2X1_LOC_160/A AND2X1_LOC_56/B 1.56fF
C6313 AND2X1_LOC_166/a_8_24# OR2X1_LOC_468/Y 0.01fF
C6314 AND2X1_LOC_143/a_8_24# AND2X1_LOC_4/a_8_24# 0.23fF
C6315 OR2X1_LOC_168/A OR2X1_LOC_66/A 0.01fF
C6316 AND2X1_LOC_719/Y AND2X1_LOC_227/Y 0.03fF
C6317 OR2X1_LOC_22/Y OR2X1_LOC_585/Y 0.08fF
C6318 AND2X1_LOC_654/a_8_24# OR2X1_LOC_619/Y 0.06fF
C6319 AND2X1_LOC_178/a_8_24# OR2X1_LOC_564/A 0.01fF
C6320 OR2X1_LOC_121/Y OR2X1_LOC_473/A 0.03fF
C6321 OR2X1_LOC_283/Y AND2X1_LOC_843/a_36_24# 0.00fF
C6322 OR2X1_LOC_160/A AND2X1_LOC_8/Y 0.63fF
C6323 OR2X1_LOC_43/A OR2X1_LOC_39/A 0.37fF
C6324 OR2X1_LOC_663/A OR2X1_LOC_404/Y 0.03fF
C6325 AND2X1_LOC_741/a_8_24# AND2X1_LOC_711/Y 0.05fF
C6326 OR2X1_LOC_91/Y OR2X1_LOC_44/Y 11.98fF
C6327 AND2X1_LOC_99/A OR2X1_LOC_89/A 0.01fF
C6328 OR2X1_LOC_856/B AND2X1_LOC_111/a_8_24# 0.02fF
C6329 OR2X1_LOC_3/Y AND2X1_LOC_76/Y 0.03fF
C6330 OR2X1_LOC_520/A OR2X1_LOC_520/a_8_216# 0.47fF
C6331 OR2X1_LOC_64/Y AND2X1_LOC_857/Y 0.02fF
C6332 OR2X1_LOC_154/A OR2X1_LOC_400/B 0.02fF
C6333 OR2X1_LOC_185/Y OR2X1_LOC_193/Y 0.16fF
C6334 OR2X1_LOC_697/Y AND2X1_LOC_712/B 0.79fF
C6335 OR2X1_LOC_145/a_8_216# OR2X1_LOC_599/A 0.01fF
C6336 OR2X1_LOC_634/A AND2X1_LOC_119/a_36_24# 0.01fF
C6337 OR2X1_LOC_811/A OR2X1_LOC_605/B 0.80fF
C6338 OR2X1_LOC_262/Y OR2X1_LOC_265/Y 0.02fF
C6339 OR2X1_LOC_600/A AND2X1_LOC_810/Y 0.07fF
C6340 AND2X1_LOC_621/Y OR2X1_LOC_239/Y 0.03fF
C6341 AND2X1_LOC_44/Y AND2X1_LOC_761/a_36_24# 0.02fF
C6342 OR2X1_LOC_655/B AND2X1_LOC_92/Y 0.23fF
C6343 OR2X1_LOC_496/a_8_216# AND2X1_LOC_675/A 0.18fF
C6344 OR2X1_LOC_70/Y OR2X1_LOC_432/a_8_216# 0.14fF
C6345 OR2X1_LOC_121/B OR2X1_LOC_776/a_36_216# 0.00fF
C6346 OR2X1_LOC_481/A OR2X1_LOC_427/A 0.11fF
C6347 OR2X1_LOC_613/Y AND2X1_LOC_620/a_8_24# 0.05fF
C6348 AND2X1_LOC_573/a_8_24# AND2X1_LOC_711/Y 0.06fF
C6349 AND2X1_LOC_715/A AND2X1_LOC_476/A 0.02fF
C6350 OR2X1_LOC_562/A OR2X1_LOC_344/a_36_216# 0.00fF
C6351 OR2X1_LOC_391/B OR2X1_LOC_269/B 0.06fF
C6352 AND2X1_LOC_8/Y AND2X1_LOC_29/a_36_24# 0.01fF
C6353 OR2X1_LOC_3/Y OR2X1_LOC_67/A 0.55fF
C6354 AND2X1_LOC_660/a_8_24# AND2X1_LOC_218/Y 0.20fF
C6355 AND2X1_LOC_489/Y AND2X1_LOC_572/A 0.37fF
C6356 OR2X1_LOC_479/Y OR2X1_LOC_738/A 0.07fF
C6357 AND2X1_LOC_554/B AND2X1_LOC_342/Y 0.02fF
C6358 OR2X1_LOC_68/B OR2X1_LOC_121/A 0.03fF
C6359 OR2X1_LOC_64/Y AND2X1_LOC_833/a_36_24# 0.01fF
C6360 OR2X1_LOC_62/B OR2X1_LOC_244/a_36_216# 0.00fF
C6361 OR2X1_LOC_26/Y AND2X1_LOC_637/Y 0.01fF
C6362 AND2X1_LOC_856/a_8_24# OR2X1_LOC_48/B 0.01fF
C6363 OR2X1_LOC_222/a_8_216# AND2X1_LOC_92/Y 0.04fF
C6364 AND2X1_LOC_512/Y OR2X1_LOC_167/Y 0.12fF
C6365 OR2X1_LOC_486/B OR2X1_LOC_739/A 0.00fF
C6366 AND2X1_LOC_314/a_36_24# AND2X1_LOC_51/Y 0.00fF
C6367 AND2X1_LOC_359/B OR2X1_LOC_7/A 0.03fF
C6368 AND2X1_LOC_211/B OR2X1_LOC_43/A 0.08fF
C6369 OR2X1_LOC_51/Y OR2X1_LOC_615/Y 0.02fF
C6370 OR2X1_LOC_92/Y AND2X1_LOC_477/A 0.07fF
C6371 OR2X1_LOC_364/A OR2X1_LOC_653/a_8_216# 0.03fF
C6372 AND2X1_LOC_789/a_8_24# INPUT_1 0.02fF
C6373 AND2X1_LOC_229/a_36_24# OR2X1_LOC_641/B 0.00fF
C6374 OR2X1_LOC_44/Y OR2X1_LOC_757/Y 0.37fF
C6375 AND2X1_LOC_347/Y OR2X1_LOC_417/A 0.02fF
C6376 AND2X1_LOC_50/Y AND2X1_LOC_7/Y 0.00fF
C6377 AND2X1_LOC_473/Y OR2X1_LOC_521/a_8_216# 0.18fF
C6378 OR2X1_LOC_60/a_8_216# OR2X1_LOC_39/A 0.03fF
C6379 OR2X1_LOC_639/B AND2X1_LOC_51/Y 0.03fF
C6380 AND2X1_LOC_99/Y AND2X1_LOC_845/Y 0.88fF
C6381 OR2X1_LOC_524/Y AND2X1_LOC_479/Y 0.80fF
C6382 AND2X1_LOC_56/B OR2X1_LOC_33/a_8_216# 0.01fF
C6383 AND2X1_LOC_86/B AND2X1_LOC_8/Y 0.04fF
C6384 OR2X1_LOC_624/B OR2X1_LOC_659/B 0.00fF
C6385 OR2X1_LOC_423/a_8_216# OR2X1_LOC_7/A 0.10fF
C6386 OR2X1_LOC_804/A OR2X1_LOC_776/Y 0.02fF
C6387 OR2X1_LOC_3/Y OR2X1_LOC_52/B 0.23fF
C6388 AND2X1_LOC_658/A AND2X1_LOC_792/Y 0.07fF
C6389 AND2X1_LOC_470/a_36_24# OR2X1_LOC_427/A 0.00fF
C6390 OR2X1_LOC_287/B OR2X1_LOC_843/a_8_216# 0.19fF
C6391 AND2X1_LOC_620/Y AND2X1_LOC_663/A 0.03fF
C6392 AND2X1_LOC_139/B OR2X1_LOC_416/Y 0.03fF
C6393 OR2X1_LOC_364/B OR2X1_LOC_578/B 0.00fF
C6394 OR2X1_LOC_130/A OR2X1_LOC_206/A 0.14fF
C6395 AND2X1_LOC_492/a_8_24# OR2X1_LOC_532/B 0.04fF
C6396 OR2X1_LOC_185/Y OR2X1_LOC_404/Y 0.10fF
C6397 OR2X1_LOC_520/Y OR2X1_LOC_121/B 0.00fF
C6398 OR2X1_LOC_71/Y OR2X1_LOC_427/A 0.06fF
C6399 OR2X1_LOC_95/Y OR2X1_LOC_586/a_8_216# 0.01fF
C6400 AND2X1_LOC_367/A OR2X1_LOC_47/Y 0.03fF
C6401 OR2X1_LOC_36/Y OR2X1_LOC_65/a_8_216# 0.02fF
C6402 OR2X1_LOC_351/B OR2X1_LOC_228/Y 0.33fF
C6403 OR2X1_LOC_46/A AND2X1_LOC_655/A 0.00fF
C6404 OR2X1_LOC_185/A AND2X1_LOC_309/a_36_24# 0.00fF
C6405 AND2X1_LOC_18/Y OR2X1_LOC_675/Y 0.02fF
C6406 OR2X1_LOC_417/Y OR2X1_LOC_44/Y 0.07fF
C6407 OR2X1_LOC_426/A AND2X1_LOC_451/Y 0.57fF
C6408 OR2X1_LOC_502/A OR2X1_LOC_62/A 0.31fF
C6409 AND2X1_LOC_59/a_36_24# AND2X1_LOC_7/Y 0.00fF
C6410 OR2X1_LOC_656/Y AND2X1_LOC_88/Y 0.01fF
C6411 OR2X1_LOC_486/Y OR2X1_LOC_367/B 0.39fF
C6412 AND2X1_LOC_554/B AND2X1_LOC_141/B 0.02fF
C6413 OR2X1_LOC_131/Y AND2X1_LOC_140/a_8_24# 0.00fF
C6414 AND2X1_LOC_574/A OR2X1_LOC_44/Y 0.09fF
C6415 OR2X1_LOC_576/A OR2X1_LOC_141/a_8_216# 0.01fF
C6416 OR2X1_LOC_772/Y OR2X1_LOC_269/B 0.01fF
C6417 OR2X1_LOC_6/B OR2X1_LOC_80/A 0.29fF
C6418 AND2X1_LOC_72/B OR2X1_LOC_735/a_8_216# 0.01fF
C6419 OR2X1_LOC_846/A OR2X1_LOC_269/B 0.03fF
C6420 AND2X1_LOC_810/Y OR2X1_LOC_619/Y 0.07fF
C6421 OR2X1_LOC_185/A OR2X1_LOC_440/A 0.03fF
C6422 OR2X1_LOC_154/A OR2X1_LOC_447/Y 0.45fF
C6423 OR2X1_LOC_601/a_8_216# OR2X1_LOC_44/Y 0.05fF
C6424 AND2X1_LOC_375/a_36_24# OR2X1_LOC_409/B 0.00fF
C6425 OR2X1_LOC_333/B AND2X1_LOC_51/Y 0.11fF
C6426 AND2X1_LOC_22/Y OR2X1_LOC_523/A 0.33fF
C6427 AND2X1_LOC_802/a_8_24# OR2X1_LOC_7/A 0.02fF
C6428 OR2X1_LOC_3/Y OR2X1_LOC_755/A 0.00fF
C6429 AND2X1_LOC_68/a_8_24# OR2X1_LOC_6/A 0.01fF
C6430 AND2X1_LOC_70/Y AND2X1_LOC_432/a_8_24# 0.02fF
C6431 OR2X1_LOC_743/A AND2X1_LOC_307/Y 0.05fF
C6432 AND2X1_LOC_8/Y OR2X1_LOC_655/A 0.01fF
C6433 OR2X1_LOC_84/B AND2X1_LOC_133/a_8_24# 0.03fF
C6434 OR2X1_LOC_59/Y AND2X1_LOC_562/Y 0.01fF
C6435 AND2X1_LOC_92/Y OR2X1_LOC_750/Y 0.10fF
C6436 OR2X1_LOC_609/A OR2X1_LOC_46/A 0.05fF
C6437 OR2X1_LOC_219/B OR2X1_LOC_814/A 0.12fF
C6438 AND2X1_LOC_12/Y OR2X1_LOC_473/A 0.18fF
C6439 OR2X1_LOC_614/a_8_216# OR2X1_LOC_87/A 0.01fF
C6440 INPUT_4 AND2X1_LOC_451/Y 0.00fF
C6441 AND2X1_LOC_472/B AND2X1_LOC_826/a_8_24# 0.01fF
C6442 AND2X1_LOC_36/Y OR2X1_LOC_138/A 0.01fF
C6443 OR2X1_LOC_703/A OR2X1_LOC_552/A 0.00fF
C6444 OR2X1_LOC_63/a_8_216# D_INPUT_1 0.01fF
C6445 OR2X1_LOC_680/A OR2X1_LOC_615/Y 0.03fF
C6446 OR2X1_LOC_599/A OR2X1_LOC_145/Y 0.01fF
C6447 OR2X1_LOC_243/B AND2X1_LOC_42/B 0.05fF
C6448 AND2X1_LOC_476/A OR2X1_LOC_753/A 0.10fF
C6449 OR2X1_LOC_76/A AND2X1_LOC_75/a_36_24# 0.00fF
C6450 AND2X1_LOC_339/a_8_24# OR2X1_LOC_31/Y 0.04fF
C6451 OR2X1_LOC_696/A AND2X1_LOC_724/A 0.01fF
C6452 OR2X1_LOC_64/Y AND2X1_LOC_685/a_36_24# 0.00fF
C6453 OR2X1_LOC_335/a_8_216# AND2X1_LOC_22/Y 0.01fF
C6454 AND2X1_LOC_91/B OR2X1_LOC_474/B 0.03fF
C6455 AND2X1_LOC_350/Y OR2X1_LOC_46/A 0.39fF
C6456 OR2X1_LOC_275/A D_INPUT_0 0.03fF
C6457 AND2X1_LOC_38/a_36_24# AND2X1_LOC_47/Y 0.00fF
C6458 AND2X1_LOC_41/A OR2X1_LOC_193/a_8_216# 0.02fF
C6459 AND2X1_LOC_201/Y AND2X1_LOC_206/a_8_24# 0.07fF
C6460 INPUT_0 OR2X1_LOC_437/A 0.07fF
C6461 OR2X1_LOC_392/B AND2X1_LOC_44/Y 0.05fF
C6462 OR2X1_LOC_779/A OR2X1_LOC_708/a_8_216# 0.01fF
C6463 OR2X1_LOC_36/Y OR2X1_LOC_419/Y 1.82fF
C6464 OR2X1_LOC_51/Y D_INPUT_6 0.90fF
C6465 AND2X1_LOC_715/Y AND2X1_LOC_724/A 0.01fF
C6466 OR2X1_LOC_149/B OR2X1_LOC_148/Y 0.14fF
C6467 OR2X1_LOC_490/Y OR2X1_LOC_47/Y 0.05fF
C6468 OR2X1_LOC_47/Y OR2X1_LOC_74/A 0.12fF
C6469 AND2X1_LOC_12/Y OR2X1_LOC_228/Y 0.12fF
C6470 OR2X1_LOC_624/A OR2X1_LOC_560/A 0.05fF
C6471 AND2X1_LOC_220/a_8_24# AND2X1_LOC_220/B 0.01fF
C6472 AND2X1_LOC_47/Y OR2X1_LOC_416/Y 0.08fF
C6473 AND2X1_LOC_627/a_8_24# OR2X1_LOC_161/B 0.01fF
C6474 AND2X1_LOC_159/a_8_24# AND2X1_LOC_497/a_8_24# 0.23fF
C6475 AND2X1_LOC_773/Y AND2X1_LOC_786/Y 0.21fF
C6476 AND2X1_LOC_12/Y OR2X1_LOC_513/Y 0.01fF
C6477 OR2X1_LOC_6/B OR2X1_LOC_115/B 0.03fF
C6478 OR2X1_LOC_244/A OR2X1_LOC_814/A 0.07fF
C6479 AND2X1_LOC_717/Y OR2X1_LOC_437/A 0.01fF
C6480 AND2X1_LOC_706/Y OR2X1_LOC_428/A 0.07fF
C6481 OR2X1_LOC_12/Y AND2X1_LOC_774/A 0.01fF
C6482 OR2X1_LOC_447/A OR2X1_LOC_446/B 0.02fF
C6483 OR2X1_LOC_598/Y OR2X1_LOC_828/Y 0.00fF
C6484 OR2X1_LOC_87/A AND2X1_LOC_31/Y 0.21fF
C6485 OR2X1_LOC_323/A AND2X1_LOC_326/B 0.01fF
C6486 OR2X1_LOC_841/B OR2X1_LOC_228/Y 0.02fF
C6487 AND2X1_LOC_64/Y OR2X1_LOC_468/A 0.03fF
C6488 OR2X1_LOC_26/Y OR2X1_LOC_72/Y 0.01fF
C6489 AND2X1_LOC_40/Y OR2X1_LOC_535/a_36_216# -0.00fF
C6490 OR2X1_LOC_3/Y AND2X1_LOC_216/A 0.22fF
C6491 OR2X1_LOC_256/a_8_216# OR2X1_LOC_13/B 0.00fF
C6492 AND2X1_LOC_696/a_8_24# AND2X1_LOC_31/Y 0.01fF
C6493 AND2X1_LOC_67/Y OR2X1_LOC_66/Y 0.02fF
C6494 AND2X1_LOC_53/Y OR2X1_LOC_651/A 1.36fF
C6495 OR2X1_LOC_235/a_8_216# OR2X1_LOC_71/A 0.01fF
C6496 OR2X1_LOC_7/A AND2X1_LOC_790/a_8_24# 0.03fF
C6497 OR2X1_LOC_51/Y AND2X1_LOC_242/B 0.03fF
C6498 OR2X1_LOC_354/A OR2X1_LOC_319/Y 0.13fF
C6499 OR2X1_LOC_323/A AND2X1_LOC_471/Y 0.18fF
C6500 OR2X1_LOC_427/A AND2X1_LOC_789/Y 0.09fF
C6501 AND2X1_LOC_390/B OR2X1_LOC_761/a_36_216# 0.01fF
C6502 AND2X1_LOC_707/Y OR2X1_LOC_51/Y 0.01fF
C6503 AND2X1_LOC_814/a_8_24# AND2X1_LOC_792/Y 0.01fF
C6504 AND2X1_LOC_658/A OR2X1_LOC_816/A 0.10fF
C6505 AND2X1_LOC_489/Y AND2X1_LOC_772/a_8_24# 0.03fF
C6506 OR2X1_LOC_599/Y OR2X1_LOC_46/A 0.06fF
C6507 OR2X1_LOC_375/A OR2X1_LOC_777/B 5.11fF
C6508 AND2X1_LOC_91/B OR2X1_LOC_561/Y 0.33fF
C6509 OR2X1_LOC_696/A AND2X1_LOC_716/Y 0.07fF
C6510 AND2X1_LOC_91/B OR2X1_LOC_78/Y 0.06fF
C6511 OR2X1_LOC_770/A OR2X1_LOC_78/B 0.01fF
C6512 OR2X1_LOC_97/A OR2X1_LOC_648/A 0.02fF
C6513 OR2X1_LOC_76/A OR2X1_LOC_318/B 0.03fF
C6514 OR2X1_LOC_421/A OR2X1_LOC_829/A 0.05fF
C6515 AND2X1_LOC_22/Y OR2X1_LOC_834/A 0.08fF
C6516 OR2X1_LOC_736/Y AND2X1_LOC_18/Y 0.03fF
C6517 OR2X1_LOC_416/Y OR2X1_LOC_598/A 0.22fF
C6518 AND2X1_LOC_351/a_8_24# OR2X1_LOC_51/Y 0.01fF
C6519 AND2X1_LOC_85/a_36_24# OR2X1_LOC_80/A 0.00fF
C6520 OR2X1_LOC_653/B AND2X1_LOC_18/Y 0.01fF
C6521 AND2X1_LOC_140/a_8_24# AND2X1_LOC_657/A 0.01fF
C6522 OR2X1_LOC_131/Y AND2X1_LOC_217/a_8_24# 0.02fF
C6523 AND2X1_LOC_705/Y AND2X1_LOC_447/Y 0.18fF
C6524 OR2X1_LOC_185/A AND2X1_LOC_238/a_8_24# 0.01fF
C6525 OR2X1_LOC_175/Y AND2X1_LOC_41/A 0.03fF
C6526 OR2X1_LOC_696/A AND2X1_LOC_654/Y 0.07fF
C6527 OR2X1_LOC_671/Y OR2X1_LOC_600/A 0.68fF
C6528 OR2X1_LOC_589/A OR2X1_LOC_536/Y 0.01fF
C6529 AND2X1_LOC_858/B AND2X1_LOC_244/A 0.03fF
C6530 OR2X1_LOC_62/A OR2X1_LOC_618/Y 0.12fF
C6531 OR2X1_LOC_846/B OR2X1_LOC_561/B 0.07fF
C6532 OR2X1_LOC_133/a_36_216# OR2X1_LOC_8/Y 0.02fF
C6533 AND2X1_LOC_43/B OR2X1_LOC_308/Y 0.07fF
C6534 AND2X1_LOC_667/a_8_24# OR2X1_LOC_598/A 0.02fF
C6535 AND2X1_LOC_56/B OR2X1_LOC_532/Y 0.01fF
C6536 OR2X1_LOC_502/A OR2X1_LOC_397/Y 0.34fF
C6537 AND2X1_LOC_40/Y OR2X1_LOC_828/Y 0.01fF
C6538 OR2X1_LOC_691/Y AND2X1_LOC_41/A 0.03fF
C6539 OR2X1_LOC_91/A OR2X1_LOC_16/A 0.05fF
C6540 AND2X1_LOC_110/Y OR2X1_LOC_356/a_8_216# 0.01fF
C6541 OR2X1_LOC_465/a_8_216# AND2X1_LOC_36/Y 0.05fF
C6542 OR2X1_LOC_840/a_8_216# OR2X1_LOC_858/A 0.40fF
C6543 OR2X1_LOC_124/Y OR2X1_LOC_217/A 0.16fF
C6544 OR2X1_LOC_198/a_8_216# OR2X1_LOC_377/A 0.02fF
C6545 AND2X1_LOC_541/Y AND2X1_LOC_768/a_8_24# 0.02fF
C6546 OR2X1_LOC_443/a_8_216# OR2X1_LOC_551/B 0.05fF
C6547 OR2X1_LOC_158/A OR2X1_LOC_56/A 19.94fF
C6548 OR2X1_LOC_696/A AND2X1_LOC_502/a_8_24# 0.00fF
C6549 OR2X1_LOC_124/a_8_216# OR2X1_LOC_6/B 0.03fF
C6550 AND2X1_LOC_91/B OR2X1_LOC_724/a_8_216# 0.01fF
C6551 OR2X1_LOC_151/A OR2X1_LOC_78/A 0.31fF
C6552 OR2X1_LOC_40/Y AND2X1_LOC_436/Y 0.16fF
C6553 AND2X1_LOC_41/A OR2X1_LOC_713/A 1.05fF
C6554 OR2X1_LOC_653/Y AND2X1_LOC_7/B 0.07fF
C6555 OR2X1_LOC_8/Y OR2X1_LOC_671/a_8_216# 0.40fF
C6556 OR2X1_LOC_104/a_8_216# OR2X1_LOC_6/B 0.09fF
C6557 AND2X1_LOC_631/a_8_24# OR2X1_LOC_816/A 0.01fF
C6558 AND2X1_LOC_788/a_8_24# AND2X1_LOC_512/Y 0.02fF
C6559 OR2X1_LOC_160/B OR2X1_LOC_244/Y 0.05fF
C6560 AND2X1_LOC_501/Y AND2X1_LOC_500/Y 0.01fF
C6561 OR2X1_LOC_347/Y OR2X1_LOC_66/A 0.02fF
C6562 AND2X1_LOC_727/Y AND2X1_LOC_624/A 0.03fF
C6563 OR2X1_LOC_833/B AND2X1_LOC_7/B 1.07fF
C6564 OR2X1_LOC_686/A OR2X1_LOC_78/B 0.02fF
C6565 OR2X1_LOC_506/a_36_216# OR2X1_LOC_375/A 0.00fF
C6566 AND2X1_LOC_42/B OR2X1_LOC_771/B 0.08fF
C6567 OR2X1_LOC_375/A OR2X1_LOC_831/B 0.00fF
C6568 OR2X1_LOC_64/Y OR2X1_LOC_437/A 0.25fF
C6569 OR2X1_LOC_108/Y AND2X1_LOC_858/B 0.07fF
C6570 AND2X1_LOC_539/Y AND2X1_LOC_388/a_8_24# 0.01fF
C6571 OR2X1_LOC_638/B VDD 0.21fF
C6572 AND2X1_LOC_570/Y AND2X1_LOC_500/Y -0.00fF
C6573 OR2X1_LOC_97/A OR2X1_LOC_405/a_8_216# 0.01fF
C6574 OR2X1_LOC_188/a_8_216# OR2X1_LOC_375/A 0.01fF
C6575 OR2X1_LOC_640/Y OR2X1_LOC_650/a_8_216# 0.39fF
C6576 OR2X1_LOC_436/Y OR2X1_LOC_854/A 0.03fF
C6577 AND2X1_LOC_719/Y AND2X1_LOC_722/A 0.00fF
C6578 AND2X1_LOC_16/a_36_24# AND2X1_LOC_44/Y 0.00fF
C6579 AND2X1_LOC_16/a_8_24# OR2X1_LOC_161/B 0.02fF
C6580 OR2X1_LOC_156/Y OR2X1_LOC_375/A 0.10fF
C6581 OR2X1_LOC_319/a_8_216# OR2X1_LOC_161/B 0.01fF
C6582 OR2X1_LOC_47/Y AND2X1_LOC_647/Y 0.08fF
C6583 OR2X1_LOC_479/Y AND2X1_LOC_36/Y 0.04fF
C6584 AND2X1_LOC_573/A AND2X1_LOC_244/A 0.03fF
C6585 OR2X1_LOC_241/a_8_216# OR2X1_LOC_121/A 0.01fF
C6586 OR2X1_LOC_696/A OR2X1_LOC_312/Y 0.01fF
C6587 VDD OR2X1_LOC_235/B 2.18fF
C6588 OR2X1_LOC_866/B OR2X1_LOC_865/Y 0.06fF
C6589 AND2X1_LOC_47/Y OR2X1_LOC_80/A 0.23fF
C6590 AND2X1_LOC_191/B OR2X1_LOC_744/A 0.02fF
C6591 AND2X1_LOC_397/a_8_24# OR2X1_LOC_402/B 0.01fF
C6592 OR2X1_LOC_811/A OR2X1_LOC_549/A 0.07fF
C6593 AND2X1_LOC_64/Y OR2X1_LOC_449/B 0.06fF
C6594 AND2X1_LOC_331/a_36_24# OR2X1_LOC_151/A 0.01fF
C6595 OR2X1_LOC_377/A OR2X1_LOC_161/B 0.03fF
C6596 AND2X1_LOC_383/a_8_24# GATE_366 0.01fF
C6597 OR2X1_LOC_858/B OR2X1_LOC_858/a_8_216# 0.39fF
C6598 OR2X1_LOC_287/B OR2X1_LOC_363/a_8_216# 0.00fF
C6599 OR2X1_LOC_744/A AND2X1_LOC_469/B 0.01fF
C6600 AND2X1_LOC_573/A OR2X1_LOC_16/A 0.03fF
C6601 OR2X1_LOC_45/B OR2X1_LOC_91/Y 0.03fF
C6602 OR2X1_LOC_158/A AND2X1_LOC_850/Y 0.04fF
C6603 OR2X1_LOC_532/B OR2X1_LOC_317/B 0.00fF
C6604 AND2X1_LOC_354/a_36_24# OR2X1_LOC_428/A 0.01fF
C6605 OR2X1_LOC_52/B AND2X1_LOC_201/Y 0.01fF
C6606 AND2X1_LOC_64/Y AND2X1_LOC_88/a_8_24# 0.02fF
C6607 AND2X1_LOC_41/A OR2X1_LOC_242/a_8_216# 0.00fF
C6608 OR2X1_LOC_45/B OR2X1_LOC_305/Y 0.02fF
C6609 OR2X1_LOC_417/A OR2X1_LOC_437/A 1.39fF
C6610 AND2X1_LOC_715/Y OR2X1_LOC_312/Y 0.06fF
C6611 OR2X1_LOC_70/A OR2X1_LOC_581/a_8_216# 0.01fF
C6612 OR2X1_LOC_192/B OR2X1_LOC_192/a_8_216# 0.07fF
C6613 OR2X1_LOC_516/a_8_216# AND2X1_LOC_212/Y 0.01fF
C6614 AND2X1_LOC_8/Y OR2X1_LOC_266/A 0.03fF
C6615 AND2X1_LOC_698/a_8_24# OR2X1_LOC_308/Y 0.04fF
C6616 OR2X1_LOC_49/A AND2X1_LOC_818/a_8_24# 0.03fF
C6617 OR2X1_LOC_709/B OR2X1_LOC_154/A 0.01fF
C6618 OR2X1_LOC_708/B OR2X1_LOC_708/a_8_216# 0.03fF
C6619 OR2X1_LOC_95/Y OR2X1_LOC_536/a_36_216# 0.00fF
C6620 OR2X1_LOC_45/B OR2X1_LOC_371/a_8_216# 0.01fF
C6621 AND2X1_LOC_314/a_8_24# OR2X1_LOC_66/A 0.03fF
C6622 OR2X1_LOC_856/B AND2X1_LOC_110/a_8_24# 0.01fF
C6623 OR2X1_LOC_517/a_8_216# OR2X1_LOC_517/A 0.01fF
C6624 AND2X1_LOC_202/a_8_24# OR2X1_LOC_72/Y 0.05fF
C6625 OR2X1_LOC_426/B OR2X1_LOC_427/A 0.02fF
C6626 OR2X1_LOC_589/A OR2X1_LOC_85/A 0.02fF
C6627 AND2X1_LOC_72/B OR2X1_LOC_68/B 0.05fF
C6628 OR2X1_LOC_421/A AND2X1_LOC_648/a_8_24# 0.01fF
C6629 OR2X1_LOC_23/a_8_216# OR2X1_LOC_59/Y -0.00fF
C6630 AND2X1_LOC_3/Y AND2X1_LOC_248/a_8_24# 0.01fF
C6631 AND2X1_LOC_861/B AND2X1_LOC_862/Y 0.01fF
C6632 OR2X1_LOC_599/A AND2X1_LOC_828/a_36_24# 0.01fF
C6633 OR2X1_LOC_820/B OR2X1_LOC_381/a_8_216# 0.01fF
C6634 AND2X1_LOC_736/Y OR2X1_LOC_524/Y 0.07fF
C6635 AND2X1_LOC_573/a_8_24# AND2X1_LOC_658/B 0.01fF
C6636 OR2X1_LOC_485/A OR2X1_LOC_428/A 0.42fF
C6637 AND2X1_LOC_514/a_8_24# AND2X1_LOC_364/A 0.04fF
C6638 AND2X1_LOC_789/a_36_24# OR2X1_LOC_820/A 0.00fF
C6639 OR2X1_LOC_604/A AND2X1_LOC_466/a_8_24# 0.01fF
C6640 AND2X1_LOC_784/A AND2X1_LOC_180/a_8_24# 0.01fF
C6641 OR2X1_LOC_426/B OR2X1_LOC_63/a_8_216# 0.02fF
C6642 OR2X1_LOC_343/B OR2X1_LOC_580/A 0.01fF
C6643 AND2X1_LOC_64/Y OR2X1_LOC_121/B 2.88fF
C6644 OR2X1_LOC_243/A OR2X1_LOC_66/A 0.00fF
C6645 AND2X1_LOC_666/a_8_24# OR2X1_LOC_121/A 0.04fF
C6646 OR2X1_LOC_185/Y OR2X1_LOC_362/A 0.06fF
C6647 AND2X1_LOC_481/a_8_24# OR2X1_LOC_294/Y 0.00fF
C6648 OR2X1_LOC_329/B AND2X1_LOC_76/Y 0.03fF
C6649 OR2X1_LOC_6/B OR2X1_LOC_6/A 0.56fF
C6650 OR2X1_LOC_80/A OR2X1_LOC_598/A 0.17fF
C6651 OR2X1_LOC_756/B OR2X1_LOC_403/A 0.02fF
C6652 OR2X1_LOC_130/A OR2X1_LOC_776/Y 0.19fF
C6653 OR2X1_LOC_200/Y AND2X1_LOC_41/Y 0.01fF
C6654 OR2X1_LOC_91/A AND2X1_LOC_661/a_8_24# 0.04fF
C6655 OR2X1_LOC_668/Y OR2X1_LOC_66/A 0.01fF
C6656 D_GATE_479 OR2X1_LOC_466/a_36_216# 0.00fF
C6657 OR2X1_LOC_480/a_8_216# OR2X1_LOC_470/B 0.01fF
C6658 AND2X1_LOC_168/Y OR2X1_LOC_91/A 0.02fF
C6659 OR2X1_LOC_505/a_36_216# OR2X1_LOC_74/A 0.02fF
C6660 AND2X1_LOC_348/a_8_24# OR2X1_LOC_428/A 0.01fF
C6661 OR2X1_LOC_364/A OR2X1_LOC_832/a_8_216# 0.01fF
C6662 AND2X1_LOC_658/A AND2X1_LOC_807/Y 0.00fF
C6663 D_INPUT_1 OR2X1_LOC_561/A 0.02fF
C6664 OR2X1_LOC_151/A OR2X1_LOC_155/A 0.07fF
C6665 OR2X1_LOC_59/Y AND2X1_LOC_287/a_8_24# 0.01fF
C6666 OR2X1_LOC_604/A OR2X1_LOC_36/Y 0.36fF
C6667 VDD AND2X1_LOC_319/A 0.29fF
C6668 OR2X1_LOC_160/A AND2X1_LOC_92/Y 0.17fF
C6669 AND2X1_LOC_675/Y OR2X1_LOC_18/Y 0.00fF
C6670 AND2X1_LOC_477/Y OR2X1_LOC_52/B 0.07fF
C6671 OR2X1_LOC_45/B OR2X1_LOC_527/Y 0.11fF
C6672 AND2X1_LOC_12/Y AND2X1_LOC_498/a_8_24# 0.00fF
C6673 OR2X1_LOC_516/Y AND2X1_LOC_675/A 0.07fF
C6674 AND2X1_LOC_367/A OR2X1_LOC_625/Y 0.24fF
C6675 OR2X1_LOC_3/Y OR2X1_LOC_281/Y 0.33fF
C6676 AND2X1_LOC_393/a_8_24# VDD -0.00fF
C6677 OR2X1_LOC_769/A OR2X1_LOC_828/B 0.15fF
C6678 AND2X1_LOC_860/a_36_24# AND2X1_LOC_850/Y 0.00fF
C6679 OR2X1_LOC_45/B OR2X1_LOC_417/Y 0.07fF
C6680 OR2X1_LOC_516/B OR2X1_LOC_48/B 0.03fF
C6681 OR2X1_LOC_719/Y OR2X1_LOC_66/A 0.01fF
C6682 OR2X1_LOC_830/a_8_216# OR2X1_LOC_269/B 0.05fF
C6683 AND2X1_LOC_509/Y OR2X1_LOC_39/A 0.04fF
C6684 OR2X1_LOC_45/B OR2X1_LOC_291/Y 0.03fF
C6685 OR2X1_LOC_3/Y OR2X1_LOC_584/Y 0.00fF
C6686 AND2X1_LOC_725/a_36_24# OR2X1_LOC_52/B 0.01fF
C6687 OR2X1_LOC_158/A OR2X1_LOC_291/A 0.02fF
C6688 OR2X1_LOC_837/A OR2X1_LOC_837/B 0.12fF
C6689 OR2X1_LOC_45/B OR2X1_LOC_311/Y 0.03fF
C6690 AND2X1_LOC_657/A AND2X1_LOC_217/a_8_24# 0.02fF
C6691 OR2X1_LOC_136/a_8_216# D_INPUT_0 0.01fF
C6692 AND2X1_LOC_840/B AND2X1_LOC_469/B 0.03fF
C6693 OR2X1_LOC_600/A AND2X1_LOC_645/A 0.19fF
C6694 OR2X1_LOC_51/Y OR2X1_LOC_22/a_8_216# 0.01fF
C6695 OR2X1_LOC_74/Y AND2X1_LOC_76/Y 0.01fF
C6696 OR2X1_LOC_178/a_8_216# OR2X1_LOC_7/A 0.01fF
C6697 OR2X1_LOC_160/B AND2X1_LOC_171/a_8_24# 0.03fF
C6698 OR2X1_LOC_45/B AND2X1_LOC_574/A 0.03fF
C6699 AND2X1_LOC_47/Y OR2X1_LOC_115/B 0.02fF
C6700 OR2X1_LOC_215/A AND2X1_LOC_65/A 0.17fF
C6701 AND2X1_LOC_533/a_8_24# OR2X1_LOC_354/A 0.26fF
C6702 OR2X1_LOC_434/a_8_216# OR2X1_LOC_805/A 0.05fF
C6703 OR2X1_LOC_756/B OR2X1_LOC_130/A 0.04fF
C6704 OR2X1_LOC_74/A OR2X1_LOC_607/A 0.11fF
C6705 OR2X1_LOC_280/Y AND2X1_LOC_489/a_8_24# 0.17fF
C6706 AND2X1_LOC_396/a_8_24# OR2X1_LOC_287/B 0.01fF
C6707 AND2X1_LOC_559/a_8_24# OR2X1_LOC_91/A 0.03fF
C6708 OR2X1_LOC_160/B AND2X1_LOC_387/B 0.12fF
C6709 OR2X1_LOC_411/Y OR2X1_LOC_690/A 0.10fF
C6710 OR2X1_LOC_7/A AND2X1_LOC_436/Y 0.03fF
C6711 OR2X1_LOC_106/Y OR2X1_LOC_95/Y 0.03fF
C6712 OR2X1_LOC_759/A OR2X1_LOC_258/a_36_216# 0.00fF
C6713 OR2X1_LOC_666/A OR2X1_LOC_89/a_8_216# 0.01fF
C6714 INPUT_0 OR2X1_LOC_753/A 0.08fF
C6715 AND2X1_LOC_733/Y AND2X1_LOC_840/B 0.23fF
C6716 OR2X1_LOC_191/B D_GATE_741 0.02fF
C6717 OR2X1_LOC_329/B OR2X1_LOC_52/B 0.19fF
C6718 OR2X1_LOC_744/A AND2X1_LOC_638/a_8_24# 0.00fF
C6719 D_INPUT_5 AND2X1_LOC_1/a_8_24# 0.01fF
C6720 OR2X1_LOC_620/Y OR2X1_LOC_161/A 0.10fF
C6721 OR2X1_LOC_532/B AND2X1_LOC_44/Y 1.17fF
C6722 AND2X1_LOC_866/A AND2X1_LOC_580/a_8_24# 0.02fF
C6723 VDD OR2X1_LOC_52/a_8_216# 0.21fF
C6724 OR2X1_LOC_147/B OR2X1_LOC_553/A 0.07fF
C6725 OR2X1_LOC_653/Y OR2X1_LOC_805/A 0.46fF
C6726 AND2X1_LOC_70/Y OR2X1_LOC_856/a_36_216# 0.00fF
C6727 OR2X1_LOC_493/B AND2X1_LOC_67/Y 0.16fF
C6728 AND2X1_LOC_675/A OR2X1_LOC_373/a_8_216# 0.01fF
C6729 OR2X1_LOC_362/B OR2X1_LOC_806/a_8_216# 0.09fF
C6730 OR2X1_LOC_377/A AND2X1_LOC_536/a_8_24# 0.03fF
C6731 OR2X1_LOC_485/A AND2X1_LOC_468/a_36_24# 0.00fF
C6732 AND2X1_LOC_302/a_8_24# AND2X1_LOC_654/Y 0.04fF
C6733 OR2X1_LOC_833/B OR2X1_LOC_805/A 0.03fF
C6734 OR2X1_LOC_203/a_8_216# OR2X1_LOC_269/a_8_216# 0.47fF
C6735 OR2X1_LOC_6/B OR2X1_LOC_611/a_36_216# 0.01fF
C6736 AND2X1_LOC_715/A OR2X1_LOC_64/Y 0.04fF
C6737 OR2X1_LOC_313/a_8_216# AND2X1_LOC_452/Y -0.02fF
C6738 AND2X1_LOC_710/a_8_24# AND2X1_LOC_847/Y 0.02fF
C6739 AND2X1_LOC_181/a_36_24# OR2X1_LOC_485/A 0.00fF
C6740 OR2X1_LOC_160/B AND2X1_LOC_75/a_36_24# 0.01fF
C6741 OR2X1_LOC_697/Y OR2X1_LOC_89/A 0.00fF
C6742 AND2X1_LOC_367/a_8_24# OR2X1_LOC_427/A 0.01fF
C6743 OR2X1_LOC_3/Y AND2X1_LOC_378/a_8_24# 0.17fF
C6744 OR2X1_LOC_164/Y OR2X1_LOC_238/Y 0.00fF
C6745 OR2X1_LOC_629/Y OR2X1_LOC_631/B 0.01fF
C6746 OR2X1_LOC_837/B OR2X1_LOC_49/a_8_216# 0.01fF
C6747 AND2X1_LOC_554/Y AND2X1_LOC_572/A 0.17fF
C6748 OR2X1_LOC_474/a_8_216# OR2X1_LOC_66/A 0.08fF
C6749 AND2X1_LOC_34/Y AND2X1_LOC_35/a_8_24# 0.06fF
C6750 OR2X1_LOC_660/B OR2X1_LOC_130/A 0.24fF
C6751 AND2X1_LOC_344/a_8_24# OR2X1_LOC_7/A 0.04fF
C6752 OR2X1_LOC_74/Y OR2X1_LOC_52/B 0.03fF
C6753 AND2X1_LOC_515/a_8_24# OR2X1_LOC_95/Y 0.05fF
C6754 AND2X1_LOC_56/B OR2X1_LOC_447/A 0.01fF
C6755 AND2X1_LOC_470/A AND2X1_LOC_452/Y 0.09fF
C6756 OR2X1_LOC_154/A OR2X1_LOC_161/A 0.27fF
C6757 OR2X1_LOC_698/Y OR2X1_LOC_258/a_36_216# 0.00fF
C6758 AND2X1_LOC_36/Y OR2X1_LOC_68/B 0.25fF
C6759 OR2X1_LOC_656/Y AND2X1_LOC_88/a_8_24# 0.24fF
C6760 OR2X1_LOC_519/Y OR2X1_LOC_6/A 0.01fF
C6761 OR2X1_LOC_433/a_8_216# OR2X1_LOC_432/Y 0.42fF
C6762 OR2X1_LOC_600/A AND2X1_LOC_477/A 0.13fF
C6763 OR2X1_LOC_859/A OR2X1_LOC_66/A 0.01fF
C6764 OR2X1_LOC_538/a_36_216# OR2X1_LOC_702/A 0.00fF
C6765 OR2X1_LOC_115/B OR2X1_LOC_598/A 0.11fF
C6766 OR2X1_LOC_185/A OR2X1_LOC_643/A 0.18fF
C6767 AND2X1_LOC_98/a_8_24# INPUT_1 0.06fF
C6768 OR2X1_LOC_43/A AND2X1_LOC_593/Y 0.35fF
C6769 OR2X1_LOC_701/Y OR2X1_LOC_701/a_8_216# 0.05fF
C6770 AND2X1_LOC_219/a_8_24# AND2X1_LOC_640/a_8_24# 0.23fF
C6771 D_INPUT_3 OR2X1_LOC_382/A 0.02fF
C6772 OR2X1_LOC_185/A OR2X1_LOC_778/Y 0.05fF
C6773 AND2X1_LOC_334/Y AND2X1_LOC_640/a_8_24# 0.00fF
C6774 AND2X1_LOC_247/a_8_24# OR2X1_LOC_437/A 0.01fF
C6775 OR2X1_LOC_306/Y OR2X1_LOC_36/Y 0.10fF
C6776 AND2X1_LOC_736/Y AND2X1_LOC_578/A 0.07fF
C6777 OR2X1_LOC_599/A AND2X1_LOC_655/A 0.02fF
C6778 OR2X1_LOC_69/A OR2X1_LOC_69/Y 0.01fF
C6779 AND2X1_LOC_31/Y OR2X1_LOC_390/B 0.13fF
C6780 OR2X1_LOC_457/B OR2X1_LOC_457/a_8_216# 0.07fF
C6781 OR2X1_LOC_619/Y AND2X1_LOC_645/A 0.02fF
C6782 AND2X1_LOC_391/Y AND2X1_LOC_128/a_8_24# 0.01fF
C6783 OR2X1_LOC_743/A OR2X1_LOC_427/A 0.13fF
C6784 OR2X1_LOC_6/B D_INPUT_2 0.05fF
C6785 OR2X1_LOC_68/B OR2X1_LOC_333/a_8_216# 0.05fF
C6786 OR2X1_LOC_655/A AND2X1_LOC_92/Y 0.01fF
C6787 OR2X1_LOC_743/A AND2X1_LOC_801/a_8_24# 0.01fF
C6788 AND2X1_LOC_715/A OR2X1_LOC_417/A 0.02fF
C6789 AND2X1_LOC_87/a_36_24# OR2X1_LOC_85/A 0.00fF
C6790 OR2X1_LOC_91/A AND2X1_LOC_128/a_8_24# 0.02fF
C6791 OR2X1_LOC_505/Y OR2X1_LOC_95/Y 0.03fF
C6792 OR2X1_LOC_532/B OR2X1_LOC_785/a_8_216# 0.03fF
C6793 AND2X1_LOC_516/a_8_24# AND2X1_LOC_43/B 0.01fF
C6794 VDD AND2X1_LOC_170/B 0.12fF
C6795 OR2X1_LOC_169/a_36_216# OR2X1_LOC_468/Y 0.00fF
C6796 OR2X1_LOC_476/B OR2X1_LOC_634/a_8_216# 0.03fF
C6797 AND2X1_LOC_12/Y OR2X1_LOC_287/B 0.05fF
C6798 OR2X1_LOC_68/B OR2X1_LOC_334/A 0.01fF
C6799 OR2X1_LOC_91/A AND2X1_LOC_687/Y 0.11fF
C6800 OR2X1_LOC_43/A OR2X1_LOC_85/A 1.61fF
C6801 OR2X1_LOC_178/a_8_216# OR2X1_LOC_224/a_8_216# 0.47fF
C6802 OR2X1_LOC_656/Y OR2X1_LOC_121/B 0.01fF
C6803 OR2X1_LOC_122/A AND2X1_LOC_845/Y 0.03fF
C6804 OR2X1_LOC_666/A AND2X1_LOC_849/a_8_24# 0.00fF
C6805 AND2X1_LOC_41/A OR2X1_LOC_750/a_8_216# 0.01fF
C6806 OR2X1_LOC_44/Y OR2X1_LOC_701/a_8_216# 0.01fF
C6807 OR2X1_LOC_864/A OR2X1_LOC_87/A 0.03fF
C6808 AND2X1_LOC_367/a_8_24# AND2X1_LOC_363/A 0.20fF
C6809 OR2X1_LOC_670/a_8_216# OR2X1_LOC_26/Y 0.01fF
C6810 AND2X1_LOC_658/A OR2X1_LOC_95/Y 0.06fF
C6811 AND2X1_LOC_191/B OR2X1_LOC_31/Y 0.00fF
C6812 OR2X1_LOC_44/Y AND2X1_LOC_806/A 0.04fF
C6813 VDD OR2X1_LOC_276/B 0.02fF
C6814 AND2X1_LOC_288/a_8_24# AND2X1_LOC_806/A 0.01fF
C6815 AND2X1_LOC_127/a_8_24# OR2X1_LOC_736/A 0.01fF
C6816 OR2X1_LOC_620/Y AND2X1_LOC_51/Y 0.07fF
C6817 OR2X1_LOC_70/Y OR2X1_LOC_432/Y 0.18fF
C6818 AND2X1_LOC_662/B AND2X1_LOC_660/Y 0.00fF
C6819 OR2X1_LOC_18/Y OR2X1_LOC_279/Y 0.19fF
C6820 OR2X1_LOC_177/Y OR2X1_LOC_419/Y 0.03fF
C6821 OR2X1_LOC_8/Y OR2X1_LOC_618/Y 0.01fF
C6822 OR2X1_LOC_47/Y AND2X1_LOC_860/A 0.03fF
C6823 AND2X1_LOC_385/a_8_24# OR2X1_LOC_389/B 0.02fF
C6824 OR2X1_LOC_690/A OR2X1_LOC_753/A 0.03fF
C6825 AND2X1_LOC_648/B AND2X1_LOC_447/Y 0.02fF
C6826 OR2X1_LOC_3/Y OR2X1_LOC_48/a_8_216# 0.05fF
C6827 OR2X1_LOC_87/A OR2X1_LOC_633/B 0.82fF
C6828 OR2X1_LOC_696/A OR2X1_LOC_13/B 1.19fF
C6829 AND2X1_LOC_259/Y AND2X1_LOC_818/a_8_24# 0.01fF
C6830 OR2X1_LOC_696/a_8_216# OR2X1_LOC_44/Y 0.02fF
C6831 AND2X1_LOC_476/A AND2X1_LOC_222/a_8_24# 0.02fF
C6832 OR2X1_LOC_66/Y AND2X1_LOC_625/a_8_24# 0.01fF
C6833 VDD AND2X1_LOC_721/A 0.60fF
C6834 AND2X1_LOC_12/Y OR2X1_LOC_76/A 0.03fF
C6835 OR2X1_LOC_705/B OR2X1_LOC_726/A 0.02fF
C6836 OR2X1_LOC_40/Y OR2X1_LOC_86/A 0.00fF
C6837 OR2X1_LOC_502/A OR2X1_LOC_818/a_36_216# 0.02fF
C6838 OR2X1_LOC_715/B AND2X1_LOC_679/a_8_24# 0.02fF
C6839 AND2X1_LOC_171/a_8_24# OR2X1_LOC_219/B 0.06fF
C6840 OR2X1_LOC_456/A OR2X1_LOC_375/A 0.03fF
C6841 OR2X1_LOC_680/Y OR2X1_LOC_26/Y 0.00fF
C6842 OR2X1_LOC_604/A OR2X1_LOC_419/Y 0.17fF
C6843 OR2X1_LOC_840/A AND2X1_LOC_47/Y 1.25fF
C6844 OR2X1_LOC_154/A AND2X1_LOC_51/Y 0.34fF
C6845 OR2X1_LOC_812/B AND2X1_LOC_494/a_8_24# 0.02fF
C6846 AND2X1_LOC_794/B OR2X1_LOC_331/Y 0.00fF
C6847 OR2X1_LOC_631/B OR2X1_LOC_629/a_36_216# 0.01fF
C6848 OR2X1_LOC_19/B AND2X1_LOC_43/B 0.18fF
C6849 INPUT_1 AND2X1_LOC_520/Y 0.02fF
C6850 OR2X1_LOC_60/a_8_216# OR2X1_LOC_85/A 0.01fF
C6851 AND2X1_LOC_647/Y OR2X1_LOC_607/A 0.01fF
C6852 OR2X1_LOC_235/B OR2X1_LOC_845/A 0.06fF
C6853 AND2X1_LOC_196/Y OR2X1_LOC_48/B 0.01fF
C6854 OR2X1_LOC_413/Y OR2X1_LOC_46/A 0.01fF
C6855 OR2X1_LOC_70/Y AND2X1_LOC_577/A 0.32fF
C6856 OR2X1_LOC_40/Y AND2X1_LOC_804/a_36_24# 0.00fF
C6857 AND2X1_LOC_477/A OR2X1_LOC_619/Y 0.11fF
C6858 GATE_366 AND2X1_LOC_663/B 0.03fF
C6859 AND2X1_LOC_715/Y OR2X1_LOC_13/B 0.10fF
C6860 OR2X1_LOC_160/B OR2X1_LOC_318/B 0.03fF
C6861 OR2X1_LOC_502/A OR2X1_LOC_651/A 0.07fF
C6862 AND2X1_LOC_554/B OR2X1_LOC_89/A 0.01fF
C6863 AND2X1_LOC_465/a_8_24# OR2X1_LOC_529/Y 0.01fF
C6864 OR2X1_LOC_680/Y OR2X1_LOC_89/A 0.15fF
C6865 OR2X1_LOC_690/A OR2X1_LOC_27/a_36_216# 0.00fF
C6866 OR2X1_LOC_124/a_8_216# OR2X1_LOC_598/A 0.02fF
C6867 VDD OR2X1_LOC_580/a_8_216# 0.00fF
C6868 OR2X1_LOC_130/A OR2X1_LOC_227/a_8_216# 0.03fF
C6869 OR2X1_LOC_154/A OR2X1_LOC_849/a_8_216# 0.03fF
C6870 OR2X1_LOC_865/A OR2X1_LOC_580/A 0.09fF
C6871 AND2X1_LOC_369/a_8_24# OR2X1_LOC_121/B 0.04fF
C6872 D_INPUT_0 OR2X1_LOC_118/Y 0.03fF
C6873 OR2X1_LOC_858/A OR2X1_LOC_493/Y 0.08fF
C6874 AND2X1_LOC_8/Y AND2X1_LOC_46/a_8_24# 0.10fF
C6875 OR2X1_LOC_64/Y OR2X1_LOC_753/A 0.02fF
C6876 OR2X1_LOC_427/A OR2X1_LOC_409/B 0.03fF
C6877 AND2X1_LOC_116/Y AND2X1_LOC_276/Y 0.06fF
C6878 AND2X1_LOC_55/a_8_24# OR2X1_LOC_62/B 0.01fF
C6879 OR2X1_LOC_657/a_8_216# OR2X1_LOC_62/B 0.01fF
C6880 AND2X1_LOC_702/Y AND2X1_LOC_537/Y 0.03fF
C6881 AND2X1_LOC_649/B AND2X1_LOC_649/Y 0.00fF
C6882 VDD OR2X1_LOC_331/Y 0.12fF
C6883 VDD AND2X1_LOC_430/B 0.47fF
C6884 OR2X1_LOC_696/Y OR2X1_LOC_89/A 0.01fF
C6885 VDD OR2X1_LOC_779/B 0.21fF
C6886 OR2X1_LOC_48/Y AND2X1_LOC_196/a_8_24# 0.01fF
C6887 AND2X1_LOC_571/A AND2X1_LOC_571/B 0.10fF
C6888 OR2X1_LOC_40/Y OR2X1_LOC_152/a_8_216# 0.02fF
C6889 OR2X1_LOC_696/A OR2X1_LOC_111/a_8_216# 0.01fF
C6890 AND2X1_LOC_23/a_8_24# OR2X1_LOC_269/B 0.02fF
C6891 OR2X1_LOC_856/a_8_216# AND2X1_LOC_51/Y 0.01fF
C6892 OR2X1_LOC_756/B OR2X1_LOC_365/B 0.00fF
C6893 OR2X1_LOC_47/Y AND2X1_LOC_400/a_8_24# 0.01fF
C6894 AND2X1_LOC_150/a_36_24# OR2X1_LOC_140/Y -0.00fF
C6895 AND2X1_LOC_831/Y AND2X1_LOC_831/a_8_24# 0.00fF
C6896 AND2X1_LOC_348/Y OR2X1_LOC_417/A 0.01fF
C6897 OR2X1_LOC_777/B OR2X1_LOC_549/A 0.07fF
C6898 OR2X1_LOC_7/Y OR2X1_LOC_585/A 0.00fF
C6899 OR2X1_LOC_436/Y OR2X1_LOC_802/A 0.01fF
C6900 AND2X1_LOC_227/Y AND2X1_LOC_266/Y 0.09fF
C6901 AND2X1_LOC_139/A AND2X1_LOC_139/B 0.03fF
C6902 OR2X1_LOC_168/B OR2X1_LOC_228/Y 0.07fF
C6903 OR2X1_LOC_630/Y OR2X1_LOC_68/B 0.07fF
C6904 OR2X1_LOC_240/B AND2X1_LOC_6/a_8_24# 0.20fF
C6905 OR2X1_LOC_417/A OR2X1_LOC_753/A 0.07fF
C6906 OR2X1_LOC_477/B OR2X1_LOC_477/a_8_216# 0.02fF
C6907 AND2X1_LOC_59/Y OR2X1_LOC_473/A 0.00fF
C6908 OR2X1_LOC_3/Y OR2X1_LOC_22/Y 2.56fF
C6909 D_INPUT_0 OR2X1_LOC_24/Y 0.01fF
C6910 OR2X1_LOC_633/a_8_216# OR2X1_LOC_68/B 0.01fF
C6911 OR2X1_LOC_45/B OR2X1_LOC_171/Y 2.76fF
C6912 AND2X1_LOC_64/Y OR2X1_LOC_857/A 0.05fF
C6913 OR2X1_LOC_510/Y OR2X1_LOC_66/a_8_216# 0.01fF
C6914 AND2X1_LOC_41/A OR2X1_LOC_546/A 0.26fF
C6915 OR2X1_LOC_602/Y OR2X1_LOC_788/B 0.06fF
C6916 OR2X1_LOC_809/a_36_216# OR2X1_LOC_112/B 0.03fF
C6917 AND2X1_LOC_390/B AND2X1_LOC_169/a_8_24# 0.02fF
C6918 AND2X1_LOC_373/a_36_24# OR2X1_LOC_440/A 0.00fF
C6919 OR2X1_LOC_193/A AND2X1_LOC_7/Y 0.14fF
C6920 AND2X1_LOC_140/a_8_24# OR2X1_LOC_256/A 0.09fF
C6921 AND2X1_LOC_626/a_36_24# AND2X1_LOC_36/Y 0.01fF
C6922 AND2X1_LOC_455/a_36_24# OR2X1_LOC_428/A 0.00fF
C6923 AND2X1_LOC_838/Y OR2X1_LOC_28/a_8_216# 0.14fF
C6924 OR2X1_LOC_599/A OR2X1_LOC_599/Y 0.01fF
C6925 OR2X1_LOC_64/Y AND2X1_LOC_845/Y 0.02fF
C6926 OR2X1_LOC_136/Y AND2X1_LOC_364/a_8_24# 0.12fF
C6927 OR2X1_LOC_78/B OR2X1_LOC_332/a_8_216# 0.01fF
C6928 OR2X1_LOC_553/A OR2X1_LOC_318/B 0.02fF
C6929 OR2X1_LOC_251/Y AND2X1_LOC_721/A 0.02fF
C6930 AND2X1_LOC_48/A OR2X1_LOC_520/A 0.01fF
C6931 OR2X1_LOC_6/A OR2X1_LOC_598/A 0.12fF
C6932 AND2X1_LOC_59/Y OR2X1_LOC_228/Y 3.56fF
C6933 OR2X1_LOC_161/A OR2X1_LOC_560/A 0.02fF
C6934 OR2X1_LOC_196/B AND2X1_LOC_53/Y 0.18fF
C6935 AND2X1_LOC_554/Y AND2X1_LOC_772/a_8_24# 0.20fF
C6936 AND2X1_LOC_81/B AND2X1_LOC_609/a_8_24# 0.01fF
C6937 AND2X1_LOC_462/Y OR2X1_LOC_416/Y 0.01fF
C6938 AND2X1_LOC_684/a_8_24# AND2X1_LOC_51/Y 0.01fF
C6939 OR2X1_LOC_136/Y OR2X1_LOC_589/A 0.84fF
C6940 OR2X1_LOC_354/A OR2X1_LOC_777/B 0.07fF
C6941 OR2X1_LOC_714/Y OR2X1_LOC_317/B 0.00fF
C6942 AND2X1_LOC_40/Y OR2X1_LOC_550/B 0.03fF
C6943 AND2X1_LOC_53/Y AND2X1_LOC_692/a_8_24# 0.02fF
C6944 OR2X1_LOC_86/A OR2X1_LOC_7/A 0.05fF
C6945 OR2X1_LOC_12/Y AND2X1_LOC_786/Y 0.07fF
C6946 OR2X1_LOC_604/A AND2X1_LOC_590/a_36_24# 0.00fF
C6947 OR2X1_LOC_506/A AND2X1_LOC_419/a_8_24# 0.01fF
C6948 OR2X1_LOC_71/a_8_216# OR2X1_LOC_71/A 0.01fF
C6949 OR2X1_LOC_532/B OR2X1_LOC_720/B 0.02fF
C6950 AND2X1_LOC_358/Y AND2X1_LOC_339/B 0.32fF
C6951 OR2X1_LOC_323/A AND2X1_LOC_112/a_8_24# 0.01fF
C6952 OR2X1_LOC_416/A OR2X1_LOC_46/A 0.26fF
C6953 AND2X1_LOC_18/Y OR2X1_LOC_120/a_8_216# 0.01fF
C6954 AND2X1_LOC_483/a_36_24# AND2X1_LOC_620/Y 0.00fF
C6955 OR2X1_LOC_712/a_8_216# OR2X1_LOC_712/B 0.02fF
C6956 OR2X1_LOC_417/A AND2X1_LOC_845/Y 0.07fF
C6957 AND2X1_LOC_785/a_8_24# AND2X1_LOC_776/a_8_24# 0.23fF
C6958 AND2X1_LOC_543/Y OR2X1_LOC_51/Y 0.01fF
C6959 AND2X1_LOC_361/A AND2X1_LOC_657/A 0.02fF
C6960 OR2X1_LOC_116/a_36_216# OR2X1_LOC_560/A 0.00fF
C6961 OR2X1_LOC_794/a_8_216# OR2X1_LOC_318/B 0.01fF
C6962 OR2X1_LOC_344/A OR2X1_LOC_549/A 0.08fF
C6963 OR2X1_LOC_111/Y OR2X1_LOC_31/Y 0.48fF
C6964 OR2X1_LOC_61/Y OR2X1_LOC_539/B 0.02fF
C6965 AND2X1_LOC_656/Y AND2X1_LOC_660/a_8_24# 0.04fF
C6966 AND2X1_LOC_636/a_8_24# OR2X1_LOC_583/Y 0.23fF
C6967 AND2X1_LOC_562/a_8_24# OR2X1_LOC_56/A 0.04fF
C6968 OR2X1_LOC_750/A OR2X1_LOC_214/B 0.06fF
C6969 AND2X1_LOC_592/Y AND2X1_LOC_706/Y 0.16fF
C6970 OR2X1_LOC_271/Y OR2X1_LOC_521/a_36_216# 0.00fF
C6971 AND2X1_LOC_564/B AND2X1_LOC_663/A 0.10fF
C6972 AND2X1_LOC_721/Y OR2X1_LOC_56/A 0.05fF
C6973 OR2X1_LOC_549/a_8_216# OR2X1_LOC_756/B 0.01fF
C6974 OR2X1_LOC_122/Y OR2X1_LOC_106/Y 0.15fF
C6975 OR2X1_LOC_22/Y AND2X1_LOC_462/B 0.72fF
C6976 OR2X1_LOC_486/Y OR2X1_LOC_543/A 0.03fF
C6977 OR2X1_LOC_177/Y OR2X1_LOC_604/A 0.03fF
C6978 OR2X1_LOC_447/Y OR2X1_LOC_783/a_8_216# 0.02fF
C6979 AND2X1_LOC_110/Y OR2X1_LOC_356/A 0.12fF
C6980 AND2X1_LOC_657/Y AND2X1_LOC_213/B 0.03fF
C6981 OR2X1_LOC_709/A VDD 0.21fF
C6982 AND2X1_LOC_22/Y AND2X1_LOC_306/a_8_24# 0.04fF
C6983 AND2X1_LOC_719/Y OR2X1_LOC_40/Y 0.03fF
C6984 AND2X1_LOC_18/Y OR2X1_LOC_596/A 0.03fF
C6985 OR2X1_LOC_51/Y AND2X1_LOC_770/a_8_24# 0.09fF
C6986 AND2X1_LOC_70/Y AND2X1_LOC_433/a_36_24# 0.00fF
C6987 OR2X1_LOC_639/A AND2X1_LOC_31/Y 0.01fF
C6988 OR2X1_LOC_78/B OR2X1_LOC_161/B 4.66fF
C6989 OR2X1_LOC_351/B OR2X1_LOC_160/B 0.17fF
C6990 OR2X1_LOC_256/A AND2X1_LOC_721/A 0.04fF
C6991 AND2X1_LOC_51/Y OR2X1_LOC_198/A 0.35fF
C6992 OR2X1_LOC_753/A AND2X1_LOC_247/a_8_24# 0.01fF
C6993 OR2X1_LOC_500/A OR2X1_LOC_500/a_8_216# 0.18fF
C6994 AND2X1_LOC_64/Y OR2X1_LOC_856/B 0.09fF
C6995 OR2X1_LOC_158/A AND2X1_LOC_285/Y 0.29fF
C6996 OR2X1_LOC_89/a_8_216# OR2X1_LOC_13/B 0.03fF
C6997 AND2X1_LOC_347/B AND2X1_LOC_711/A 0.05fF
C6998 OR2X1_LOC_604/A OR2X1_LOC_745/a_8_216# 0.12fF
C6999 OR2X1_LOC_51/Y OR2X1_LOC_322/Y 0.01fF
C7000 OR2X1_LOC_40/Y OR2X1_LOC_745/a_36_216# 0.02fF
C7001 OR2X1_LOC_146/a_8_216# OR2X1_LOC_427/A 0.01fF
C7002 OR2X1_LOC_114/B OR2X1_LOC_160/B 0.03fF
C7003 OR2X1_LOC_160/A AND2X1_LOC_235/a_36_24# 0.00fF
C7004 AND2X1_LOC_360/a_8_24# OR2X1_LOC_428/A 0.01fF
C7005 OR2X1_LOC_185/Y OR2X1_LOC_776/A 0.13fF
C7006 OR2X1_LOC_117/a_8_216# OR2X1_LOC_92/Y 0.04fF
C7007 OR2X1_LOC_97/A OR2X1_LOC_61/a_36_216# 0.00fF
C7008 AND2X1_LOC_91/B OR2X1_LOC_185/A 0.03fF
C7009 AND2X1_LOC_40/Y OR2X1_LOC_61/A 0.13fF
C7010 OR2X1_LOC_721/Y OR2X1_LOC_161/B 0.03fF
C7011 OR2X1_LOC_600/a_8_216# AND2X1_LOC_447/Y 0.03fF
C7012 VDD OR2X1_LOC_758/Y 0.15fF
C7013 OR2X1_LOC_629/a_8_216# OR2X1_LOC_777/B 0.04fF
C7014 VDD AND2X1_LOC_70/Y 1.07fF
C7015 AND2X1_LOC_12/Y OR2X1_LOC_722/B 0.01fF
C7016 OR2X1_LOC_186/Y OR2X1_LOC_502/A 0.19fF
C7017 AND2X1_LOC_711/a_36_24# AND2X1_LOC_347/B 0.00fF
C7018 AND2X1_LOC_663/B OR2X1_LOC_13/B 0.03fF
C7019 OR2X1_LOC_205/Y OR2X1_LOC_215/a_8_216# 0.06fF
C7020 OR2X1_LOC_475/a_8_216# AND2X1_LOC_65/A 0.18fF
C7021 OR2X1_LOC_31/Y OR2X1_LOC_588/a_8_216# 0.03fF
C7022 OR2X1_LOC_479/Y OR2X1_LOC_469/B 0.09fF
C7023 OR2X1_LOC_160/B OR2X1_LOC_538/A 0.00fF
C7024 OR2X1_LOC_850/B OR2X1_LOC_349/A 0.03fF
C7025 OR2X1_LOC_31/Y AND2X1_LOC_203/a_8_24# 0.01fF
C7026 AND2X1_LOC_311/a_8_24# OR2X1_LOC_66/A 0.09fF
C7027 AND2X1_LOC_47/Y OR2X1_LOC_739/a_8_216# 0.05fF
C7028 AND2X1_LOC_555/Y OR2X1_LOC_43/A 0.07fF
C7029 OR2X1_LOC_52/B OR2X1_LOC_525/a_8_216# 0.06fF
C7030 OR2X1_LOC_117/a_8_216# OR2X1_LOC_65/B 0.02fF
C7031 OR2X1_LOC_6/B OR2X1_LOC_216/A 0.03fF
C7032 OR2X1_LOC_816/Y OR2X1_LOC_56/A 0.02fF
C7033 OR2X1_LOC_31/Y AND2X1_LOC_206/Y 0.02fF
C7034 OR2X1_LOC_815/Y AND2X1_LOC_793/Y 0.02fF
C7035 AND2X1_LOC_700/a_8_24# AND2X1_LOC_41/A 0.02fF
C7036 VDD AND2X1_LOC_605/Y 0.29fF
C7037 OR2X1_LOC_287/A OR2X1_LOC_78/A -0.00fF
C7038 VDD OR2X1_LOC_703/A 0.06fF
C7039 AND2X1_LOC_32/a_8_24# AND2X1_LOC_7/B 0.01fF
C7040 OR2X1_LOC_756/B OR2X1_LOC_468/A 0.02fF
C7041 AND2X1_LOC_366/A OR2X1_LOC_666/A 0.01fF
C7042 AND2X1_LOC_95/Y OR2X1_LOC_185/a_36_216# 0.02fF
C7043 OR2X1_LOC_47/Y AND2X1_LOC_562/Y 0.05fF
C7044 OR2X1_LOC_615/Y AND2X1_LOC_790/a_8_24# 0.03fF
C7045 OR2X1_LOC_132/Y OR2X1_LOC_91/A 0.26fF
C7046 OR2X1_LOC_32/B OR2X1_LOC_16/A 5.66fF
C7047 OR2X1_LOC_375/A OR2X1_LOC_161/B 0.41fF
C7048 OR2X1_LOC_136/Y OR2X1_LOC_43/A 0.07fF
C7049 AND2X1_LOC_719/Y AND2X1_LOC_843/Y -0.05fF
C7050 OR2X1_LOC_494/Y OR2X1_LOC_256/Y 0.01fF
C7051 AND2X1_LOC_392/A AND2X1_LOC_716/Y 0.07fF
C7052 OR2X1_LOC_653/Y OR2X1_LOC_648/B 0.18fF
C7053 INPUT_0 AND2X1_LOC_222/a_8_24# 0.01fF
C7054 OR2X1_LOC_254/B OR2X1_LOC_580/B 1.57fF
C7055 AND2X1_LOC_363/Y OR2X1_LOC_256/Y 0.28fF
C7056 OR2X1_LOC_482/Y AND2X1_LOC_850/Y 0.07fF
C7057 AND2X1_LOC_534/a_8_24# AND2X1_LOC_43/B 0.22fF
C7058 OR2X1_LOC_31/Y OR2X1_LOC_164/a_8_216# 0.01fF
C7059 AND2X1_LOC_588/B AND2X1_LOC_51/A 0.01fF
C7060 AND2X1_LOC_509/Y AND2X1_LOC_474/A 0.15fF
C7061 OR2X1_LOC_306/a_36_216# OR2X1_LOC_829/A 0.13fF
C7062 OR2X1_LOC_203/a_36_216# OR2X1_LOC_549/A 0.01fF
C7063 OR2X1_LOC_435/a_8_216# OR2X1_LOC_78/A 0.01fF
C7064 OR2X1_LOC_51/Y AND2X1_LOC_866/B 0.02fF
C7065 OR2X1_LOC_421/A OR2X1_LOC_48/B 0.09fF
C7066 OR2X1_LOC_529/a_8_216# AND2X1_LOC_541/Y 0.01fF
C7067 OR2X1_LOC_45/B AND2X1_LOC_806/A 0.03fF
C7068 OR2X1_LOC_131/A OR2X1_LOC_118/Y 0.00fF
C7069 OR2X1_LOC_526/Y OR2X1_LOC_485/a_36_216# 0.00fF
C7070 AND2X1_LOC_392/A AND2X1_LOC_654/Y 0.01fF
C7071 AND2X1_LOC_849/a_8_24# OR2X1_LOC_13/B 0.00fF
C7072 AND2X1_LOC_777/a_8_24# OR2X1_LOC_12/Y 0.01fF
C7073 AND2X1_LOC_720/a_8_24# AND2X1_LOC_860/A 0.01fF
C7074 AND2X1_LOC_707/Y OR2X1_LOC_423/a_8_216# 0.03fF
C7075 D_INPUT_1 OR2X1_LOC_80/A 0.34fF
C7076 AND2X1_LOC_50/Y AND2X1_LOC_70/a_8_24# 0.24fF
C7077 OR2X1_LOC_51/Y OR2X1_LOC_495/Y 0.01fF
C7078 OR2X1_LOC_421/A OR2X1_LOC_18/Y 0.01fF
C7079 OR2X1_LOC_445/a_8_216# AND2X1_LOC_7/B 0.01fF
C7080 OR2X1_LOC_625/Y AND2X1_LOC_860/A 0.07fF
C7081 AND2X1_LOC_810/A AND2X1_LOC_715/a_8_24# 0.01fF
C7082 OR2X1_LOC_161/A OR2X1_LOC_723/a_8_216# 0.14fF
C7083 OR2X1_LOC_6/B AND2X1_LOC_403/B 0.12fF
C7084 AND2X1_LOC_690/a_36_24# OR2X1_LOC_66/A 0.00fF
C7085 AND2X1_LOC_560/a_8_24# AND2X1_LOC_523/Y 0.01fF
C7086 OR2X1_LOC_604/A OR2X1_LOC_252/a_8_216# 0.07fF
C7087 OR2X1_LOC_91/Y OR2X1_LOC_158/A 0.03fF
C7088 OR2X1_LOC_105/a_8_216# OR2X1_LOC_561/Y 0.01fF
C7089 OR2X1_LOC_756/B OR2X1_LOC_571/a_8_216# 0.01fF
C7090 OR2X1_LOC_507/B OR2X1_LOC_507/A 0.18fF
C7091 OR2X1_LOC_185/A AND2X1_LOC_86/a_36_24# 0.01fF
C7092 AND2X1_LOC_31/Y OR2X1_LOC_493/Y 0.02fF
C7093 OR2X1_LOC_91/A OR2X1_LOC_426/A 0.16fF
C7094 AND2X1_LOC_500/B OR2X1_LOC_39/A 0.02fF
C7095 OR2X1_LOC_40/Y AND2X1_LOC_655/A 0.03fF
C7096 OR2X1_LOC_604/A AND2X1_LOC_467/a_8_24# 0.01fF
C7097 AND2X1_LOC_110/Y AND2X1_LOC_43/B 0.02fF
C7098 OR2X1_LOC_114/B AND2X1_LOC_297/a_36_24# 0.00fF
C7099 OR2X1_LOC_596/Y OR2X1_LOC_596/A 0.04fF
C7100 AND2X1_LOC_12/Y OR2X1_LOC_160/B 5.76fF
C7101 OR2X1_LOC_61/Y OR2X1_LOC_78/B 0.03fF
C7102 OR2X1_LOC_9/Y AND2X1_LOC_852/a_8_24# 0.01fF
C7103 AND2X1_LOC_532/a_36_24# AND2X1_LOC_436/Y 0.00fF
C7104 OR2X1_LOC_797/B OR2X1_LOC_213/B 0.01fF
C7105 OR2X1_LOC_763/Y OR2X1_LOC_12/Y 0.01fF
C7106 OR2X1_LOC_791/B VDD 0.09fF
C7107 AND2X1_LOC_95/Y OR2X1_LOC_35/Y 0.04fF
C7108 AND2X1_LOC_539/Y AND2X1_LOC_855/a_8_24# 0.01fF
C7109 AND2X1_LOC_362/B OR2X1_LOC_26/Y 0.16fF
C7110 OR2X1_LOC_26/Y AND2X1_LOC_476/Y 0.09fF
C7111 AND2X1_LOC_361/a_36_24# AND2X1_LOC_361/A 0.02fF
C7112 OR2X1_LOC_6/B OR2X1_LOC_44/Y 0.01fF
C7113 AND2X1_LOC_713/Y OR2X1_LOC_44/Y 0.01fF
C7114 AND2X1_LOC_353/a_36_24# OR2X1_LOC_36/Y 0.00fF
C7115 OR2X1_LOC_471/Y OR2X1_LOC_731/A 0.07fF
C7116 AND2X1_LOC_373/a_8_24# OR2X1_LOC_439/B 0.20fF
C7117 OR2X1_LOC_62/B OR2X1_LOC_140/B 2.28fF
C7118 OR2X1_LOC_351/B OR2X1_LOC_219/B 0.10fF
C7119 VDD OR2X1_LOC_193/Y 0.12fF
C7120 OR2X1_LOC_750/Y AND2X1_LOC_751/a_8_24# 0.00fF
C7121 AND2X1_LOC_719/Y OR2X1_LOC_7/A 0.07fF
C7122 AND2X1_LOC_362/B OR2X1_LOC_89/A 0.10fF
C7123 AND2X1_LOC_82/Y OR2X1_LOC_402/a_36_216# 0.00fF
C7124 OR2X1_LOC_89/A AND2X1_LOC_476/Y 0.11fF
C7125 OR2X1_LOC_517/A AND2X1_LOC_520/Y 0.00fF
C7126 OR2X1_LOC_528/Y AND2X1_LOC_474/Y 0.14fF
C7127 AND2X1_LOC_718/a_36_24# OR2X1_LOC_48/B 0.01fF
C7128 VDD AND2X1_LOC_361/A 0.01fF
C7129 OR2X1_LOC_756/B AND2X1_LOC_487/a_8_24# 0.01fF
C7130 AND2X1_LOC_456/B OR2X1_LOC_18/Y 0.04fF
C7131 OR2X1_LOC_89/A OR2X1_LOC_382/a_36_216# -0.00fF
C7132 OR2X1_LOC_40/Y OR2X1_LOC_609/A 0.03fF
C7133 OR2X1_LOC_820/a_8_216# OR2X1_LOC_3/Y 0.01fF
C7134 AND2X1_LOC_374/a_8_24# OR2X1_LOC_427/A 0.01fF
C7135 AND2X1_LOC_845/Y OR2X1_LOC_89/a_36_216# 0.01fF
C7136 AND2X1_LOC_3/Y OR2X1_LOC_629/B 0.02fF
C7137 AND2X1_LOC_392/A OR2X1_LOC_312/Y 0.07fF
C7138 VDD AND2X1_LOC_17/Y 0.93fF
C7139 AND2X1_LOC_704/a_8_24# OR2X1_LOC_70/Y 0.01fF
C7140 OR2X1_LOC_43/A OR2X1_LOC_51/Y 0.19fF
C7141 OR2X1_LOC_297/a_8_216# AND2X1_LOC_847/Y 0.03fF
C7142 OR2X1_LOC_840/A OR2X1_LOC_506/A 0.05fF
C7143 AND2X1_LOC_523/Y OR2X1_LOC_522/Y 0.79fF
C7144 OR2X1_LOC_768/A OR2X1_LOC_673/Y 0.01fF
C7145 OR2X1_LOC_748/A OR2X1_LOC_56/A 0.00fF
C7146 OR2X1_LOC_458/a_8_216# OR2X1_LOC_805/A 0.05fF
C7147 AND2X1_LOC_85/a_8_24# AND2X1_LOC_18/Y 0.10fF
C7148 AND2X1_LOC_710/Y OR2X1_LOC_748/A 0.01fF
C7149 AND2X1_LOC_141/A OR2X1_LOC_65/B 0.03fF
C7150 OR2X1_LOC_848/a_8_216# OR2X1_LOC_391/A 0.03fF
C7151 OR2X1_LOC_203/Y OR2X1_LOC_630/B 0.03fF
C7152 OR2X1_LOC_456/A OR2X1_LOC_549/A 0.01fF
C7153 OR2X1_LOC_264/Y AND2X1_LOC_517/a_36_24# 0.01fF
C7154 AND2X1_LOC_366/A GATE_366 0.01fF
C7155 AND2X1_LOC_784/A INPUT_0 0.07fF
C7156 D_INPUT_0 AND2X1_LOC_208/Y 0.01fF
C7157 VDD OR2X1_LOC_653/a_8_216# 0.00fF
C7158 OR2X1_LOC_160/B AND2X1_LOC_496/a_8_24# 0.06fF
C7159 OR2X1_LOC_753/A OR2X1_LOC_232/Y 0.01fF
C7160 OR2X1_LOC_158/A OR2X1_LOC_417/Y 0.03fF
C7161 OR2X1_LOC_235/B OR2X1_LOC_845/a_36_216# 0.00fF
C7162 OR2X1_LOC_318/A OR2X1_LOC_814/A 0.03fF
C7163 OR2X1_LOC_756/B AND2X1_LOC_282/a_36_24# 0.00fF
C7164 OR2X1_LOC_91/Y OR2X1_LOC_103/Y 0.03fF
C7165 OR2X1_LOC_158/A OR2X1_LOC_291/Y 0.07fF
C7166 AND2X1_LOC_843/Y AND2X1_LOC_850/a_36_24# 0.00fF
C7167 OR2X1_LOC_680/A AND2X1_LOC_866/B 2.26fF
C7168 AND2X1_LOC_86/Y OR2X1_LOC_100/a_8_216# 0.18fF
C7169 AND2X1_LOC_81/B OR2X1_LOC_502/A -0.01fF
C7170 OR2X1_LOC_158/A OR2X1_LOC_311/Y 0.03fF
C7171 OR2X1_LOC_756/B OR2X1_LOC_449/B 0.03fF
C7172 AND2X1_LOC_337/B AND2X1_LOC_434/Y 0.03fF
C7173 OR2X1_LOC_45/B AND2X1_LOC_831/Y 0.01fF
C7174 OR2X1_LOC_502/A OR2X1_LOC_358/B 0.05fF
C7175 OR2X1_LOC_405/A OR2X1_LOC_739/A 0.01fF
C7176 OR2X1_LOC_799/A OR2X1_LOC_185/A 0.07fF
C7177 D_INPUT_5 AND2X1_LOC_17/a_8_24# 0.01fF
C7178 OR2X1_LOC_329/B OR2X1_LOC_280/Y 0.09fF
C7179 OR2X1_LOC_506/B OR2X1_LOC_392/B 0.03fF
C7180 INPUT_3 AND2X1_LOC_12/Y 0.10fF
C7181 AND2X1_LOC_293/a_8_24# AND2X1_LOC_219/A 0.05fF
C7182 OR2X1_LOC_272/Y AND2X1_LOC_218/Y 0.01fF
C7183 OR2X1_LOC_151/A OR2X1_LOC_814/A 0.07fF
C7184 OR2X1_LOC_705/B OR2X1_LOC_727/a_8_216# 0.14fF
C7185 AND2X1_LOC_191/B OR2X1_LOC_488/a_8_216# 0.02fF
C7186 OR2X1_LOC_326/B OR2X1_LOC_468/Y 0.33fF
C7187 OR2X1_LOC_304/Y OR2X1_LOC_56/A 0.13fF
C7188 AND2X1_LOC_753/B OR2X1_LOC_200/a_8_216# 0.02fF
C7189 AND2X1_LOC_349/a_36_24# OR2X1_LOC_92/Y 0.01fF
C7190 OR2X1_LOC_333/B AND2X1_LOC_41/A 0.03fF
C7191 D_INPUT_7 AND2X1_LOC_12/a_8_24# 0.01fF
C7192 INPUT_3 AND2X1_LOC_838/Y 0.00fF
C7193 AND2X1_LOC_753/B OR2X1_LOC_269/B 0.16fF
C7194 AND2X1_LOC_452/Y AND2X1_LOC_470/B 0.23fF
C7195 OR2X1_LOC_273/Y AND2X1_LOC_219/Y 0.02fF
C7196 AND2X1_LOC_79/a_8_24# AND2X1_LOC_18/Y 0.06fF
C7197 AND2X1_LOC_512/Y OR2X1_LOC_485/A 0.02fF
C7198 OR2X1_LOC_87/A OR2X1_LOC_784/Y 0.16fF
C7199 AND2X1_LOC_851/B AND2X1_LOC_455/B 0.05fF
C7200 OR2X1_LOC_49/A AND2X1_LOC_672/a_8_24# 0.04fF
C7201 OR2X1_LOC_497/Y OR2X1_LOC_427/A 0.07fF
C7202 OR2X1_LOC_51/Y AND2X1_LOC_685/a_8_24# 0.05fF
C7203 AND2X1_LOC_186/a_8_24# AND2X1_LOC_624/A 0.05fF
C7204 OR2X1_LOC_805/A AND2X1_LOC_272/a_8_24# 0.00fF
C7205 OR2X1_LOC_426/B OR2X1_LOC_416/Y 0.01fF
C7206 AND2X1_LOC_754/a_8_24# AND2X1_LOC_47/Y 0.01fF
C7207 OR2X1_LOC_591/Y OR2X1_LOC_31/Y 0.29fF
C7208 OR2X1_LOC_209/A OR2X1_LOC_151/a_8_216# 0.01fF
C7209 AND2X1_LOC_715/A OR2X1_LOC_268/a_36_216# 0.03fF
C7210 OR2X1_LOC_146/Y AND2X1_LOC_213/B 0.31fF
C7211 AND2X1_LOC_856/A OR2X1_LOC_48/B 0.04fF
C7212 OR2X1_LOC_405/A OR2X1_LOC_269/B 0.42fF
C7213 OR2X1_LOC_87/A OR2X1_LOC_738/A 0.07fF
C7214 AND2X1_LOC_742/a_8_24# GATE_811 0.05fF
C7215 AND2X1_LOC_211/B AND2X1_LOC_364/A 0.31fF
C7216 OR2X1_LOC_460/Y OR2X1_LOC_375/A 0.02fF
C7217 AND2X1_LOC_95/Y OR2X1_LOC_720/a_8_216# 0.01fF
C7218 OR2X1_LOC_865/B OR2X1_LOC_774/Y 0.06fF
C7219 AND2X1_LOC_840/A OR2X1_LOC_238/Y 0.28fF
C7220 AND2X1_LOC_436/B OR2X1_LOC_44/Y 0.00fF
C7221 OR2X1_LOC_860/a_8_216# OR2X1_LOC_287/B 0.00fF
C7222 OR2X1_LOC_628/Y OR2X1_LOC_56/A 0.09fF
C7223 OR2X1_LOC_158/A D_INPUT_3 0.04fF
C7224 AND2X1_LOC_471/a_8_24# OR2X1_LOC_56/A 0.01fF
C7225 OR2X1_LOC_26/Y OR2X1_LOC_595/a_8_216# 0.07fF
C7226 OR2X1_LOC_210/a_36_216# OR2X1_LOC_87/A 0.00fF
C7227 OR2X1_LOC_36/Y OR2X1_LOC_265/Y 0.03fF
C7228 OR2X1_LOC_123/a_8_216# D_INPUT_0 0.02fF
C7229 OR2X1_LOC_756/B OR2X1_LOC_121/B 0.03fF
C7230 OR2X1_LOC_329/B OR2X1_LOC_22/Y 0.94fF
C7231 OR2X1_LOC_329/a_8_216# OR2X1_LOC_47/Y 0.01fF
C7232 AND2X1_LOC_86/Y AND2X1_LOC_79/Y 0.15fF
C7233 AND2X1_LOC_12/Y OR2X1_LOC_219/B 0.06fF
C7234 OR2X1_LOC_18/Y AND2X1_LOC_717/B 0.16fF
C7235 OR2X1_LOC_715/B AND2X1_LOC_109/a_8_24# 0.13fF
C7236 OR2X1_LOC_252/Y OR2X1_LOC_7/A 0.17fF
C7237 OR2X1_LOC_154/A OR2X1_LOC_214/a_8_216# 0.03fF
C7238 AND2X1_LOC_59/Y OR2X1_LOC_287/B 0.04fF
C7239 OR2X1_LOC_640/Y AND2X1_LOC_47/Y 0.05fF
C7240 OR2X1_LOC_292/Y OR2X1_LOC_295/Y 0.04fF
C7241 AND2X1_LOC_852/a_8_24# AND2X1_LOC_852/Y 0.03fF
C7242 AND2X1_LOC_267/a_8_24# AND2X1_LOC_361/A -0.03fF
C7243 OR2X1_LOC_185/A OR2X1_LOC_455/A 0.13fF
C7244 AND2X1_LOC_808/A AND2X1_LOC_477/Y 0.01fF
C7245 OR2X1_LOC_516/A OR2X1_LOC_485/A 0.03fF
C7246 AND2X1_LOC_555/Y OR2X1_LOC_384/a_8_216# 0.01fF
C7247 AND2X1_LOC_192/Y AND2X1_LOC_220/Y 0.12fF
C7248 OR2X1_LOC_419/Y AND2X1_LOC_212/Y 0.10fF
C7249 AND2X1_LOC_823/a_8_24# OR2X1_LOC_269/B 0.05fF
C7250 OR2X1_LOC_3/Y OR2X1_LOC_39/A 0.18fF
C7251 OR2X1_LOC_502/A OR2X1_LOC_196/B 0.01fF
C7252 AND2X1_LOC_561/B AND2X1_LOC_866/A 0.07fF
C7253 OR2X1_LOC_485/A AND2X1_LOC_342/Y 0.23fF
C7254 AND2X1_LOC_8/Y OR2X1_LOC_99/a_36_216# 0.02fF
C7255 AND2X1_LOC_8/a_8_24# INPUT_2 0.01fF
C7256 OR2X1_LOC_84/A OR2X1_LOC_66/A 0.02fF
C7257 OR2X1_LOC_405/A OR2X1_LOC_215/A 0.03fF
C7258 OR2X1_LOC_440/A AND2X1_LOC_437/a_8_24# -0.00fF
C7259 OR2X1_LOC_85/A AND2X1_LOC_240/Y 0.01fF
C7260 OR2X1_LOC_320/Y AND2X1_LOC_655/A 0.10fF
C7261 OR2X1_LOC_95/Y OR2X1_LOC_597/a_8_216# 0.01fF
C7262 OR2X1_LOC_6/B OR2X1_LOC_205/Y 0.00fF
C7263 AND2X1_LOC_456/Y AND2X1_LOC_576/Y 0.02fF
C7264 OR2X1_LOC_246/Y OR2X1_LOC_74/A 0.03fF
C7265 AND2X1_LOC_631/Y OR2X1_LOC_39/A 0.03fF
C7266 OR2X1_LOC_74/Y OR2X1_LOC_22/Y 0.06fF
C7267 OR2X1_LOC_529/Y OR2X1_LOC_44/Y 0.03fF
C7268 OR2X1_LOC_75/Y AND2X1_LOC_219/Y 0.03fF
C7269 OR2X1_LOC_656/B OR2X1_LOC_656/a_8_216# 0.02fF
C7270 OR2X1_LOC_277/a_8_216# AND2X1_LOC_573/A 0.02fF
C7271 VDD OR2X1_LOC_430/Y 0.16fF
C7272 AND2X1_LOC_576/Y OR2X1_LOC_74/A 0.07fF
C7273 OR2X1_LOC_661/a_36_216# OR2X1_LOC_476/B 0.01fF
C7274 AND2X1_LOC_40/Y AND2X1_LOC_7/Y 0.03fF
C7275 AND2X1_LOC_472/B AND2X1_LOC_459/a_8_24# 0.14fF
C7276 INPUT_0 OR2X1_LOC_62/A 0.06fF
C7277 OR2X1_LOC_318/a_8_216# OR2X1_LOC_228/Y 0.02fF
C7278 AND2X1_LOC_849/A AND2X1_LOC_573/A 0.02fF
C7279 AND2X1_LOC_729/Y OR2X1_LOC_64/Y 0.51fF
C7280 AND2X1_LOC_18/a_8_24# AND2X1_LOC_7/a_8_24# 0.23fF
C7281 AND2X1_LOC_59/Y OR2X1_LOC_76/A 0.01fF
C7282 OR2X1_LOC_414/a_8_216# OR2X1_LOC_46/A 0.01fF
C7283 VDD AND2X1_LOC_795/Y 0.06fF
C7284 OR2X1_LOC_759/A AND2X1_LOC_793/Y 0.01fF
C7285 AND2X1_LOC_758/a_8_24# AND2X1_LOC_805/a_8_24# 0.23fF
C7286 OR2X1_LOC_481/A OR2X1_LOC_6/A 0.04fF
C7287 AND2X1_LOC_580/A OR2X1_LOC_755/A 0.04fF
C7288 AND2X1_LOC_98/Y D_INPUT_3 0.01fF
C7289 OR2X1_LOC_98/B OR2X1_LOC_66/A 0.23fF
C7290 OR2X1_LOC_598/a_8_216# AND2X1_LOC_36/Y 0.06fF
C7291 OR2X1_LOC_141/B AND2X1_LOC_3/Y 0.03fF
C7292 OR2X1_LOC_804/a_8_216# OR2X1_LOC_223/A 0.01fF
C7293 OR2X1_LOC_792/Y OR2X1_LOC_288/A 0.01fF
C7294 AND2X1_LOC_553/A AND2X1_LOC_227/Y 0.55fF
C7295 OR2X1_LOC_687/Y OR2X1_LOC_687/a_8_216# 0.01fF
C7296 OR2X1_LOC_3/Y AND2X1_LOC_211/B 0.07fF
C7297 OR2X1_LOC_22/Y AND2X1_LOC_113/Y 0.06fF
C7298 OR2X1_LOC_103/Y D_INPUT_3 0.00fF
C7299 AND2X1_LOC_72/a_36_24# AND2X1_LOC_3/Y 0.00fF
C7300 OR2X1_LOC_431/a_8_216# OR2X1_LOC_26/Y 0.14fF
C7301 OR2X1_LOC_175/Y OR2X1_LOC_112/A 0.03fF
C7302 OR2X1_LOC_665/Y AND2X1_LOC_483/a_8_24# 0.03fF
C7303 AND2X1_LOC_784/A OR2X1_LOC_64/Y 0.14fF
C7304 OR2X1_LOC_485/A OR2X1_LOC_279/a_8_216# 0.03fF
C7305 OR2X1_LOC_11/Y AND2X1_LOC_639/A 0.01fF
C7306 AND2X1_LOC_456/B AND2X1_LOC_620/Y 0.39fF
C7307 OR2X1_LOC_43/A AND2X1_LOC_855/a_36_24# 0.00fF
C7308 AND2X1_LOC_724/A OR2X1_LOC_589/Y 0.01fF
C7309 AND2X1_LOC_714/a_36_24# OR2X1_LOC_423/Y 0.00fF
C7310 AND2X1_LOC_48/A OR2X1_LOC_358/B 0.00fF
C7311 AND2X1_LOC_99/A OR2X1_LOC_95/Y 0.03fF
C7312 OR2X1_LOC_502/A OR2X1_LOC_112/B 0.03fF
C7313 AND2X1_LOC_185/a_36_24# OR2X1_LOC_615/Y 0.00fF
C7314 OR2X1_LOC_794/a_8_216# OR2X1_LOC_804/B 0.01fF
C7315 OR2X1_LOC_840/A D_INPUT_1 0.00fF
C7316 OR2X1_LOC_743/A OR2X1_LOC_681/Y 0.02fF
C7317 OR2X1_LOC_241/Y OR2X1_LOC_506/A 0.01fF
C7318 D_INPUT_3 OR2X1_LOC_847/A 0.54fF
C7319 OR2X1_LOC_476/B OR2X1_LOC_472/A 0.01fF
C7320 AND2X1_LOC_769/a_8_24# OR2X1_LOC_64/Y 0.01fF
C7321 OR2X1_LOC_864/A OR2X1_LOC_649/a_8_216# 0.01fF
C7322 OR2X1_LOC_698/Y AND2X1_LOC_793/Y 0.01fF
C7323 OR2X1_LOC_620/a_8_216# OR2X1_LOC_550/B 0.06fF
C7324 OR2X1_LOC_285/Y OR2X1_LOC_269/B 0.01fF
C7325 OR2X1_LOC_97/B INPUT_1 0.22fF
C7326 OR2X1_LOC_321/Y AND2X1_LOC_324/a_8_24# 0.23fF
C7327 OR2X1_LOC_244/A OR2X1_LOC_266/a_36_216# 0.01fF
C7328 OR2X1_LOC_802/Y AND2X1_LOC_47/Y 0.18fF
C7329 OR2X1_LOC_743/A OR2X1_LOC_416/Y 0.03fF
C7330 OR2X1_LOC_429/Y OR2X1_LOC_582/Y 0.13fF
C7331 OR2X1_LOC_485/A OR2X1_LOC_54/Y 0.05fF
C7332 OR2X1_LOC_216/A OR2X1_LOC_598/A 0.02fF
C7333 AND2X1_LOC_57/Y OR2X1_LOC_175/Y 0.05fF
C7334 AND2X1_LOC_784/A OR2X1_LOC_417/A 0.25fF
C7335 OR2X1_LOC_339/A OR2X1_LOC_390/A 0.07fF
C7336 AND2X1_LOC_196/Y OR2X1_LOC_585/A 0.03fF
C7337 OR2X1_LOC_515/A OR2X1_LOC_515/a_8_216# 0.39fF
C7338 OR2X1_LOC_256/A AND2X1_LOC_361/A 0.02fF
C7339 AND2X1_LOC_772/Y AND2X1_LOC_773/a_8_24# 0.07fF
C7340 AND2X1_LOC_56/B OR2X1_LOC_620/A 0.01fF
C7341 OR2X1_LOC_599/Y AND2X1_LOC_644/Y 0.79fF
C7342 AND2X1_LOC_392/A OR2X1_LOC_13/B 0.01fF
C7343 OR2X1_LOC_739/A OR2X1_LOC_330/a_8_216# 0.01fF
C7344 OR2X1_LOC_696/A OR2X1_LOC_428/A 0.50fF
C7345 OR2X1_LOC_160/A OR2X1_LOC_215/a_8_216# 0.04fF
C7346 OR2X1_LOC_244/A AND2X1_LOC_79/Y 0.08fF
C7347 OR2X1_LOC_617/Y AND2X1_LOC_621/a_8_24# 0.09fF
C7348 AND2X1_LOC_476/A OR2X1_LOC_52/B 0.07fF
C7349 OR2X1_LOC_274/Y OR2X1_LOC_68/B 1.56fF
C7350 AND2X1_LOC_557/a_8_24# OR2X1_LOC_71/Y 0.01fF
C7351 OR2X1_LOC_6/A D_INPUT_1 0.13fF
C7352 OR2X1_LOC_696/A OR2X1_LOC_595/A 0.07fF
C7353 OR2X1_LOC_419/Y AND2X1_LOC_447/a_8_24# 0.01fF
C7354 OR2X1_LOC_92/Y AND2X1_LOC_793/B 0.02fF
C7355 AND2X1_LOC_785/a_8_24# AND2X1_LOC_785/Y 0.11fF
C7356 AND2X1_LOC_776/Y AND2X1_LOC_786/Y 0.02fF
C7357 AND2X1_LOC_773/Y AND2X1_LOC_772/Y 0.17fF
C7358 OR2X1_LOC_246/A OR2X1_LOC_416/Y 0.01fF
C7359 OR2X1_LOC_499/a_8_216# OR2X1_LOC_598/A 0.03fF
C7360 AND2X1_LOC_663/A OR2X1_LOC_437/A 0.10fF
C7361 AND2X1_LOC_168/Y AND2X1_LOC_222/Y 0.01fF
C7362 OR2X1_LOC_623/B OR2X1_LOC_513/Y 0.13fF
C7363 OR2X1_LOC_244/Y AND2X1_LOC_246/a_8_24# 0.00fF
C7364 AND2X1_LOC_383/a_8_24# OR2X1_LOC_428/A 0.04fF
C7365 AND2X1_LOC_48/A OR2X1_LOC_196/B 0.61fF
C7366 OR2X1_LOC_611/a_8_216# OR2X1_LOC_62/B 0.01fF
C7367 AND2X1_LOC_715/Y OR2X1_LOC_428/A 0.08fF
C7368 OR2X1_LOC_625/Y AND2X1_LOC_562/Y 0.10fF
C7369 OR2X1_LOC_574/A OR2X1_LOC_223/A 0.03fF
C7370 AND2X1_LOC_721/A OR2X1_LOC_248/Y 0.00fF
C7371 OR2X1_LOC_34/a_8_216# OR2X1_LOC_338/A 0.01fF
C7372 AND2X1_LOC_436/a_8_24# OR2X1_LOC_13/B 0.01fF
C7373 OR2X1_LOC_719/Y OR2X1_LOC_241/B 0.02fF
C7374 AND2X1_LOC_366/A OR2X1_LOC_13/B 0.01fF
C7375 AND2X1_LOC_721/A OR2X1_LOC_6/a_8_216# 0.47fF
C7376 OR2X1_LOC_449/A OR2X1_LOC_796/B 0.02fF
C7377 AND2X1_LOC_821/a_8_24# AND2X1_LOC_51/Y 0.01fF
C7378 OR2X1_LOC_201/a_8_216# OR2X1_LOC_201/Y 0.02fF
C7379 AND2X1_LOC_1/Y AND2X1_LOC_47/Y 0.20fF
C7380 OR2X1_LOC_87/A OR2X1_LOC_451/B 0.02fF
C7381 OR2X1_LOC_158/A AND2X1_LOC_780/a_8_24# 0.01fF
C7382 AND2X1_LOC_48/A AND2X1_LOC_692/a_8_24# 0.04fF
C7383 OR2X1_LOC_516/Y OR2X1_LOC_600/A 0.11fF
C7384 D_INPUT_0 OR2X1_LOC_750/A 0.43fF
C7385 AND2X1_LOC_687/a_36_24# OR2X1_LOC_7/A 0.01fF
C7386 OR2X1_LOC_86/A OR2X1_LOC_86/a_8_216# 0.01fF
C7387 VDD OR2X1_LOC_387/A 0.06fF
C7388 AND2X1_LOC_49/a_36_24# OR2X1_LOC_598/A 0.00fF
C7389 AND2X1_LOC_572/Y AND2X1_LOC_657/A 0.00fF
C7390 AND2X1_LOC_593/Y OR2X1_LOC_534/Y 0.21fF
C7391 OR2X1_LOC_235/B OR2X1_LOC_523/A 0.01fF
C7392 OR2X1_LOC_114/Y OR2X1_LOC_140/a_36_216# 0.00fF
C7393 OR2X1_LOC_633/A OR2X1_LOC_548/B 0.01fF
C7394 OR2X1_LOC_459/B OR2X1_LOC_460/A 0.88fF
C7395 OR2X1_LOC_22/A OR2X1_LOC_408/Y 0.02fF
C7396 OR2X1_LOC_49/A OR2X1_LOC_133/a_8_216# 0.01fF
C7397 OR2X1_LOC_196/Y OR2X1_LOC_790/A 0.16fF
C7398 OR2X1_LOC_199/a_8_216# OR2X1_LOC_614/Y 0.10fF
C7399 OR2X1_LOC_471/Y AND2X1_LOC_47/Y 0.03fF
C7400 OR2X1_LOC_185/A OR2X1_LOC_446/B 0.03fF
C7401 AND2X1_LOC_649/Y OR2X1_LOC_46/A 0.02fF
C7402 OR2X1_LOC_161/B OR2X1_LOC_549/A 0.07fF
C7403 AND2X1_LOC_354/Y OR2X1_LOC_13/B 0.06fF
C7404 OR2X1_LOC_589/A AND2X1_LOC_407/a_36_24# 0.00fF
C7405 AND2X1_LOC_727/A AND2X1_LOC_319/a_8_24# 0.01fF
C7406 OR2X1_LOC_74/A AND2X1_LOC_784/a_36_24# 0.01fF
C7407 OR2X1_LOC_538/A OR2X1_LOC_354/a_8_216# 0.01fF
C7408 OR2X1_LOC_10/a_8_216# OR2X1_LOC_54/Y 0.01fF
C7409 OR2X1_LOC_421/A OR2X1_LOC_764/a_8_216# 0.01fF
C7410 AND2X1_LOC_787/A AND2X1_LOC_722/a_8_24# 0.00fF
C7411 AND2X1_LOC_672/B OR2X1_LOC_673/A 0.02fF
C7412 AND2X1_LOC_648/B OR2X1_LOC_46/A 0.00fF
C7413 OR2X1_LOC_392/B AND2X1_LOC_18/Y 0.10fF
C7414 OR2X1_LOC_45/B OR2X1_LOC_6/B 1.16fF
C7415 AND2X1_LOC_562/a_8_24# AND2X1_LOC_285/Y 0.00fF
C7416 OR2X1_LOC_45/B AND2X1_LOC_713/Y 0.01fF
C7417 AND2X1_LOC_187/a_36_24# OR2X1_LOC_742/B 0.01fF
C7418 AND2X1_LOC_727/A AND2X1_LOC_810/a_8_24# 0.01fF
C7419 OR2X1_LOC_273/Y OR2X1_LOC_595/Y 0.01fF
C7420 AND2X1_LOC_263/a_8_24# AND2X1_LOC_18/Y 0.03fF
C7421 AND2X1_LOC_645/A OR2X1_LOC_534/a_8_216# 0.04fF
C7422 OR2X1_LOC_506/B OR2X1_LOC_532/B 0.01fF
C7423 AND2X1_LOC_810/A AND2X1_LOC_535/Y 0.01fF
C7424 INPUT_0 OR2X1_LOC_397/Y 0.03fF
C7425 OR2X1_LOC_533/Y OR2X1_LOC_604/A 0.03fF
C7426 AND2X1_LOC_727/Y OR2X1_LOC_524/Y 0.03fF
C7427 OR2X1_LOC_336/a_8_216# VDD 0.00fF
C7428 AND2X1_LOC_552/A AND2X1_LOC_476/Y 0.04fF
C7429 AND2X1_LOC_22/Y OR2X1_LOC_35/Y 0.03fF
C7430 OR2X1_LOC_78/A OR2X1_LOC_563/A 0.09fF
C7431 OR2X1_LOC_604/A AND2X1_LOC_212/Y 0.10fF
C7432 OR2X1_LOC_853/a_36_216# OR2X1_LOC_35/Y 0.03fF
C7433 OR2X1_LOC_47/Y AND2X1_LOC_800/a_36_24# 0.00fF
C7434 OR2X1_LOC_596/A OR2X1_LOC_596/a_36_216# 0.00fF
C7435 AND2X1_LOC_544/Y AND2X1_LOC_551/B 0.10fF
C7436 AND2X1_LOC_727/a_8_24# AND2X1_LOC_658/A 0.03fF
C7437 OR2X1_LOC_443/Y OR2X1_LOC_551/B 0.01fF
C7438 AND2X1_LOC_817/B OR2X1_LOC_771/B 0.00fF
C7439 AND2X1_LOC_338/A AND2X1_LOC_338/a_8_24# 0.01fF
C7440 AND2X1_LOC_712/Y AND2X1_LOC_725/a_8_24# 0.18fF
C7441 OR2X1_LOC_64/Y OR2X1_LOC_88/Y 0.03fF
C7442 AND2X1_LOC_732/B AND2X1_LOC_448/a_8_24# 0.19fF
C7443 OR2X1_LOC_329/B AND2X1_LOC_445/a_36_24# 0.01fF
C7444 OR2X1_LOC_114/a_8_216# AND2X1_LOC_44/Y 0.01fF
C7445 OR2X1_LOC_160/A OR2X1_LOC_500/a_36_216# 0.01fF
C7446 OR2X1_LOC_9/Y VDD 0.72fF
C7447 VDD AND2X1_LOC_193/Y 0.25fF
C7448 OR2X1_LOC_674/Y AND2X1_LOC_675/a_8_24# 0.01fF
C7449 VDD OR2X1_LOC_362/A 0.39fF
C7450 AND2X1_LOC_339/B OR2X1_LOC_59/Y 0.07fF
C7451 OR2X1_LOC_161/A OR2X1_LOC_605/Y 0.01fF
C7452 OR2X1_LOC_87/A AND2X1_LOC_36/Y 0.13fF
C7453 OR2X1_LOC_36/Y OR2X1_LOC_183/a_8_216# 0.06fF
C7454 OR2X1_LOC_97/A AND2X1_LOC_749/a_8_24# 0.01fF
C7455 OR2X1_LOC_44/Y AND2X1_LOC_791/a_8_24# 0.01fF
C7456 OR2X1_LOC_482/a_8_216# OR2X1_LOC_59/Y 0.01fF
C7457 GATE_811 AND2X1_LOC_808/A 0.09fF
C7458 OR2X1_LOC_417/A AND2X1_LOC_643/a_8_24# 0.02fF
C7459 VDD OR2X1_LOC_832/a_8_216# 0.21fF
C7460 AND2X1_LOC_95/Y OR2X1_LOC_115/B 0.06fF
C7461 OR2X1_LOC_501/B OR2X1_LOC_151/A 0.07fF
C7462 OR2X1_LOC_354/A OR2X1_LOC_161/B 0.07fF
C7463 OR2X1_LOC_415/a_8_216# OR2X1_LOC_80/A 0.06fF
C7464 AND2X1_LOC_721/A OR2X1_LOC_10/a_36_216# 0.00fF
C7465 AND2X1_LOC_705/Y AND2X1_LOC_722/A 0.15fF
C7466 AND2X1_LOC_320/a_36_24# OR2X1_LOC_151/A 0.01fF
C7467 AND2X1_LOC_713/a_8_24# AND2X1_LOC_605/Y 0.00fF
C7468 OR2X1_LOC_654/A OR2X1_LOC_771/B 0.02fF
C7469 AND2X1_LOC_541/Y OR2X1_LOC_744/A 0.15fF
C7470 AND2X1_LOC_477/A OR2X1_LOC_534/a_8_216# 0.04fF
C7471 VDD AND2X1_LOC_61/Y 0.15fF
C7472 OR2X1_LOC_415/A OR2X1_LOC_71/A 0.01fF
C7473 OR2X1_LOC_624/A OR2X1_LOC_267/Y 0.05fF
C7474 AND2X1_LOC_729/Y AND2X1_LOC_544/Y 0.03fF
C7475 OR2X1_LOC_93/Y OR2X1_LOC_91/A 0.12fF
C7476 OR2X1_LOC_440/a_8_216# AND2X1_LOC_92/Y 0.05fF
C7477 AND2X1_LOC_508/B OR2X1_LOC_56/A 0.01fF
C7478 AND2X1_LOC_665/a_36_24# OR2X1_LOC_675/Y 0.01fF
C7479 OR2X1_LOC_220/A OR2X1_LOC_740/B 0.03fF
C7480 AND2X1_LOC_40/Y OR2X1_LOC_390/A 0.07fF
C7481 OR2X1_LOC_506/a_8_216# OR2X1_LOC_185/Y 0.09fF
C7482 AND2X1_LOC_94/Y OR2X1_LOC_66/A 0.03fF
C7483 AND2X1_LOC_367/A OR2X1_LOC_108/Y 0.06fF
C7484 OR2X1_LOC_8/Y INPUT_0 0.02fF
C7485 OR2X1_LOC_711/B OR2X1_LOC_469/Y 0.05fF
C7486 OR2X1_LOC_841/A AND2X1_LOC_164/a_8_24# 0.23fF
C7487 AND2X1_LOC_828/a_8_24# OR2X1_LOC_48/B 0.01fF
C7488 OR2X1_LOC_151/A OR2X1_LOC_147/B 0.14fF
C7489 AND2X1_LOC_573/Y OR2X1_LOC_498/Y 0.15fF
C7490 AND2X1_LOC_509/Y OR2X1_LOC_51/Y 0.02fF
C7491 AND2X1_LOC_787/a_8_24# AND2X1_LOC_794/B 0.02fF
C7492 OR2X1_LOC_805/A AND2X1_LOC_248/a_8_24# 0.06fF
C7493 AND2X1_LOC_84/Y OR2X1_LOC_69/Y 0.80fF
C7494 OR2X1_LOC_205/Y OR2X1_LOC_598/A 0.14fF
C7495 OR2X1_LOC_45/B AND2X1_LOC_139/B 0.03fF
C7496 OR2X1_LOC_18/Y AND2X1_LOC_828/a_8_24# 0.01fF
C7497 AND2X1_LOC_712/a_36_24# AND2X1_LOC_454/Y 0.00fF
C7498 OR2X1_LOC_304/a_8_216# OR2X1_LOC_36/Y 0.01fF
C7499 OR2X1_LOC_270/a_8_216# OR2X1_LOC_577/Y 0.01fF
C7500 OR2X1_LOC_154/A OR2X1_LOC_576/A 0.07fF
C7501 AND2X1_LOC_796/Y AND2X1_LOC_796/A 0.23fF
C7502 OR2X1_LOC_188/Y OR2X1_LOC_719/Y 0.02fF
C7503 OR2X1_LOC_858/A OR2X1_LOC_541/A 0.29fF
C7504 VDD OR2X1_LOC_474/Y 1.02fF
C7505 OR2X1_LOC_369/Y AND2X1_LOC_543/a_8_24# 0.09fF
C7506 OR2X1_LOC_100/Y AND2X1_LOC_18/Y 0.08fF
C7507 OR2X1_LOC_151/A OR2X1_LOC_317/A 0.09fF
C7508 OR2X1_LOC_154/a_8_216# OR2X1_LOC_87/A 0.02fF
C7509 OR2X1_LOC_537/A OR2X1_LOC_390/A 0.00fF
C7510 AND2X1_LOC_50/Y OR2X1_LOC_66/A 0.00fF
C7511 AND2X1_LOC_509/a_8_24# AND2X1_LOC_850/A 0.03fF
C7512 OR2X1_LOC_858/B OR2X1_LOC_858/A 0.46fF
C7513 OR2X1_LOC_286/B OR2X1_LOC_580/A 0.08fF
C7514 OR2X1_LOC_438/Y AND2X1_LOC_658/A 0.11fF
C7515 AND2X1_LOC_658/A AND2X1_LOC_865/a_8_24# 0.01fF
C7516 OR2X1_LOC_6/A OR2X1_LOC_15/a_8_216# 0.14fF
C7517 OR2X1_LOC_842/a_8_216# OR2X1_LOC_78/A 0.01fF
C7518 AND2X1_LOC_22/Y OR2X1_LOC_720/a_8_216# 0.06fF
C7519 OR2X1_LOC_653/B OR2X1_LOC_130/A 0.01fF
C7520 OR2X1_LOC_506/Y OR2X1_LOC_87/A 0.04fF
C7521 AND2X1_LOC_2/Y D_INPUT_4 0.04fF
C7522 AND2X1_LOC_51/Y OR2X1_LOC_605/Y 0.37fF
C7523 OR2X1_LOC_427/A OR2X1_LOC_582/a_8_216# 0.05fF
C7524 AND2X1_LOC_477/Y OR2X1_LOC_39/A 0.10fF
C7525 AND2X1_LOC_705/Y OR2X1_LOC_599/A 0.02fF
C7526 AND2X1_LOC_547/Y AND2X1_LOC_550/A 0.14fF
C7527 OR2X1_LOC_160/A OR2X1_LOC_6/B 0.14fF
C7528 OR2X1_LOC_757/A AND2X1_LOC_866/B 0.11fF
C7529 AND2X1_LOC_508/B AND2X1_LOC_850/Y 0.00fF
C7530 AND2X1_LOC_841/B AND2X1_LOC_436/Y 0.03fF
C7531 OR2X1_LOC_604/A AND2X1_LOC_447/a_8_24# 0.08fF
C7532 OR2X1_LOC_766/a_8_216# OR2X1_LOC_52/B 0.03fF
C7533 OR2X1_LOC_45/B OR2X1_LOC_529/Y 0.02fF
C7534 AND2X1_LOC_553/A OR2X1_LOC_107/Y 0.01fF
C7535 AND2X1_LOC_95/Y OR2X1_LOC_370/a_36_216# 0.02fF
C7536 OR2X1_LOC_185/A OR2X1_LOC_542/B 0.03fF
C7537 AND2X1_LOC_292/a_8_24# OR2X1_LOC_736/Y 0.03fF
C7538 OR2X1_LOC_441/a_36_216# OR2X1_LOC_441/Y 0.00fF
C7539 AND2X1_LOC_59/Y OR2X1_LOC_160/B 0.48fF
C7540 AND2X1_LOC_572/Y VDD 0.33fF
C7541 OR2X1_LOC_859/a_8_216# OR2X1_LOC_862/A 0.04fF
C7542 OR2X1_LOC_801/B AND2X1_LOC_751/a_36_24# 0.01fF
C7543 OR2X1_LOC_116/A VDD -0.00fF
C7544 AND2X1_LOC_658/A AND2X1_LOC_621/Y 31.40fF
C7545 OR2X1_LOC_40/Y AND2X1_LOC_266/Y 0.03fF
C7546 OR2X1_LOC_158/A AND2X1_LOC_806/A 0.06fF
C7547 AND2X1_LOC_42/B AND2X1_LOC_44/Y 0.45fF
C7548 OR2X1_LOC_348/Y OR2X1_LOC_664/Y 0.02fF
C7549 INPUT_0 AND2X1_LOC_76/Y 0.02fF
C7550 OR2X1_LOC_203/Y AND2X1_LOC_625/a_8_24# 0.02fF
C7551 INPUT_5 D_INPUT_5 1.38fF
C7552 OR2X1_LOC_418/a_8_216# OR2X1_LOC_12/Y 0.01fF
C7553 AND2X1_LOC_721/Y OR2X1_LOC_527/Y 0.02fF
C7554 AND2X1_LOC_52/Y OR2X1_LOC_198/A 0.01fF
C7555 AND2X1_LOC_706/Y OR2X1_LOC_89/A 0.01fF
C7556 OR2X1_LOC_837/A OR2X1_LOC_837/Y 0.02fF
C7557 OR2X1_LOC_74/A OR2X1_LOC_16/A 0.09fF
C7558 OR2X1_LOC_529/a_8_216# OR2X1_LOC_744/A 0.05fF
C7559 OR2X1_LOC_629/a_8_216# OR2X1_LOC_161/B 0.01fF
C7560 OR2X1_LOC_641/Y OR2X1_LOC_130/A 0.02fF
C7561 VDD OR2X1_LOC_217/Y 0.06fF
C7562 AND2X1_LOC_364/Y AND2X1_LOC_662/B 0.01fF
C7563 VDD OR2X1_LOC_96/B -0.00fF
C7564 AND2X1_LOC_710/Y AND2X1_LOC_848/a_8_24# 0.01fF
C7565 OR2X1_LOC_705/Y AND2X1_LOC_44/Y 0.03fF
C7566 OR2X1_LOC_122/Y AND2X1_LOC_99/A 0.02fF
C7567 OR2X1_LOC_715/B AND2X1_LOC_516/a_8_24# 0.02fF
C7568 OR2X1_LOC_122/A OR2X1_LOC_67/A 0.03fF
C7569 AND2X1_LOC_348/A OR2X1_LOC_92/Y 0.50fF
C7570 AND2X1_LOC_734/Y OR2X1_LOC_427/A 3.32fF
C7571 OR2X1_LOC_744/A OR2X1_LOC_316/Y 0.03fF
C7572 AND2X1_LOC_663/B OR2X1_LOC_428/A 0.08fF
C7573 OR2X1_LOC_329/B OR2X1_LOC_39/A 0.12fF
C7574 AND2X1_LOC_850/A AND2X1_LOC_850/Y 0.00fF
C7575 VDD D_GATE_865 0.06fF
C7576 OR2X1_LOC_58/Y OR2X1_LOC_26/Y 0.03fF
C7577 OR2X1_LOC_426/B OR2X1_LOC_6/A 0.17fF
C7578 OR2X1_LOC_421/A OR2X1_LOC_585/A 0.00fF
C7579 VDD AND2X1_LOC_852/Y 0.61fF
C7580 AND2X1_LOC_859/a_8_24# OR2X1_LOC_59/Y 0.00fF
C7581 OR2X1_LOC_70/Y AND2X1_LOC_339/B 0.03fF
C7582 OR2X1_LOC_158/A AND2X1_LOC_276/Y 0.14fF
C7583 AND2X1_LOC_95/Y OR2X1_LOC_840/A 0.01fF
C7584 OR2X1_LOC_40/Y OR2X1_LOC_387/Y 0.11fF
C7585 VDD OR2X1_LOC_83/Y 0.24fF
C7586 OR2X1_LOC_6/B AND2X1_LOC_86/B 0.61fF
C7587 AND2X1_LOC_663/B OR2X1_LOC_595/A 0.10fF
C7588 OR2X1_LOC_538/a_8_216# OR2X1_LOC_161/A 0.04fF
C7589 AND2X1_LOC_474/A AND2X1_LOC_572/A 0.03fF
C7590 AND2X1_LOC_535/Y AND2X1_LOC_355/a_36_24# 0.00fF
C7591 AND2X1_LOC_456/Y OR2X1_LOC_108/Y 0.00fF
C7592 OR2X1_LOC_837/Y AND2X1_LOC_34/Y 0.03fF
C7593 OR2X1_LOC_380/A OR2X1_LOC_26/a_8_216# 0.01fF
C7594 OR2X1_LOC_405/A OR2X1_LOC_475/a_8_216# 0.04fF
C7595 OR2X1_LOC_71/Y OR2X1_LOC_184/a_8_216# 0.08fF
C7596 OR2X1_LOC_117/Y OR2X1_LOC_56/A 0.02fF
C7597 OR2X1_LOC_154/A AND2X1_LOC_41/A 0.46fF
C7598 AND2X1_LOC_208/a_8_24# AND2X1_LOC_35/Y 0.26fF
C7599 AND2X1_LOC_511/a_8_24# AND2X1_LOC_51/Y 0.06fF
C7600 OR2X1_LOC_426/B OR2X1_LOC_299/a_8_216# 0.03fF
C7601 OR2X1_LOC_109/a_8_216# OR2X1_LOC_427/A 0.03fF
C7602 INPUT_3 AND2X1_LOC_852/B 0.22fF
C7603 AND2X1_LOC_42/a_36_24# OR2X1_LOC_66/A 0.01fF
C7604 AND2X1_LOC_631/a_8_24# AND2X1_LOC_621/Y 0.02fF
C7605 OR2X1_LOC_323/A AND2X1_LOC_851/B 0.11fF
C7606 OR2X1_LOC_850/A OR2X1_LOC_858/a_8_216# 0.02fF
C7607 AND2X1_LOC_787/a_36_24# OR2X1_LOC_48/B 0.01fF
C7608 AND2X1_LOC_72/B OR2X1_LOC_844/B 0.84fF
C7609 OR2X1_LOC_347/a_8_216# OR2X1_LOC_347/B 0.01fF
C7610 OR2X1_LOC_74/Y OR2X1_LOC_39/A 0.04fF
C7611 INPUT_0 OR2X1_LOC_52/B 0.04fF
C7612 AND2X1_LOC_41/A OR2X1_LOC_267/A 0.05fF
C7613 AND2X1_LOC_805/Y AND2X1_LOC_807/a_8_24# 0.01fF
C7614 OR2X1_LOC_329/B AND2X1_LOC_211/B 0.07fF
C7615 OR2X1_LOC_635/A OR2X1_LOC_87/A 0.01fF
C7616 OR2X1_LOC_264/Y OR2X1_LOC_264/a_8_216# 0.05fF
C7617 AND2X1_LOC_86/Y AND2X1_LOC_59/Y 0.13fF
C7618 AND2X1_LOC_364/Y AND2X1_LOC_337/B 0.34fF
C7619 AND2X1_LOC_566/B AND2X1_LOC_326/a_8_24# 0.00fF
C7620 OR2X1_LOC_405/A OR2X1_LOC_539/Y 0.03fF
C7621 AND2X1_LOC_390/B OR2X1_LOC_744/A 0.07fF
C7622 AND2X1_LOC_342/Y OR2X1_LOC_256/a_8_216# 0.04fF
C7623 AND2X1_LOC_572/a_8_24# OR2X1_LOC_47/Y 0.17fF
C7624 AND2X1_LOC_656/Y OR2X1_LOC_12/Y 0.03fF
C7625 AND2X1_LOC_259/Y OR2X1_LOC_292/Y 0.14fF
C7626 AND2X1_LOC_50/Y OR2X1_LOC_651/a_8_216# 0.01fF
C7627 OR2X1_LOC_3/Y AND2X1_LOC_474/A 0.03fF
C7628 OR2X1_LOC_8/Y OR2X1_LOC_64/Y 0.00fF
C7629 OR2X1_LOC_3/Y OR2X1_LOC_421/a_8_216# 0.05fF
C7630 OR2X1_LOC_69/Y OR2X1_LOC_393/a_8_216# 0.04fF
C7631 AND2X1_LOC_524/a_36_24# OR2X1_LOC_545/B 0.00fF
C7632 AND2X1_LOC_95/Y OR2X1_LOC_222/A 0.06fF
C7633 AND2X1_LOC_132/a_8_24# OR2X1_LOC_375/A 0.03fF
C7634 AND2X1_LOC_523/Y OR2X1_LOC_56/A 0.03fF
C7635 OR2X1_LOC_856/a_8_216# AND2X1_LOC_41/A 0.05fF
C7636 AND2X1_LOC_318/Y AND2X1_LOC_802/Y 0.00fF
C7637 AND2X1_LOC_387/a_8_24# AND2X1_LOC_48/A 0.03fF
C7638 AND2X1_LOC_560/B AND2X1_LOC_76/Y 0.01fF
C7639 OR2X1_LOC_464/A OR2X1_LOC_733/B 1.01fF
C7640 AND2X1_LOC_344/a_36_24# AND2X1_LOC_363/A 0.00fF
C7641 AND2X1_LOC_95/Y OR2X1_LOC_6/A 0.04fF
C7642 OR2X1_LOC_574/A OR2X1_LOC_502/A 0.10fF
C7643 OR2X1_LOC_91/A AND2X1_LOC_729/B 0.07fF
C7644 AND2X1_LOC_59/Y OR2X1_LOC_553/A 0.13fF
C7645 OR2X1_LOC_158/A AND2X1_LOC_831/Y 0.07fF
C7646 OR2X1_LOC_185/A AND2X1_LOC_56/B 1.45fF
C7647 OR2X1_LOC_654/A OR2X1_LOC_637/B 0.11fF
C7648 OR2X1_LOC_506/A OR2X1_LOC_468/Y 0.03fF
C7649 AND2X1_LOC_41/A OR2X1_LOC_778/A 0.02fF
C7650 VDD OR2X1_LOC_243/B 0.02fF
C7651 OR2X1_LOC_103/Y AND2X1_LOC_276/Y 0.17fF
C7652 AND2X1_LOC_371/a_8_24# OR2X1_LOC_532/B 0.01fF
C7653 OR2X1_LOC_634/A AND2X1_LOC_51/Y 0.02fF
C7654 AND2X1_LOC_2/Y AND2X1_LOC_425/Y 0.10fF
C7655 OR2X1_LOC_185/A AND2X1_LOC_8/Y 0.11fF
C7656 OR2X1_LOC_493/Y OR2X1_LOC_121/A 0.03fF
C7657 AND2X1_LOC_785/a_36_24# OR2X1_LOC_406/A 0.01fF
C7658 OR2X1_LOC_532/B AND2X1_LOC_18/Y 0.24fF
C7659 OR2X1_LOC_757/A AND2X1_LOC_664/a_8_24# 0.01fF
C7660 AND2X1_LOC_641/Y AND2X1_LOC_641/a_36_24# 0.00fF
C7661 OR2X1_LOC_666/A AND2X1_LOC_66/a_8_24# 0.01fF
C7662 OR2X1_LOC_87/A AND2X1_LOC_129/a_36_24# 0.00fF
C7663 OR2X1_LOC_599/A OR2X1_LOC_511/Y 0.02fF
C7664 OR2X1_LOC_70/Y OR2X1_LOC_586/a_8_216# 0.09fF
C7665 AND2X1_LOC_168/Y OR2X1_LOC_74/A 0.39fF
C7666 OR2X1_LOC_154/A OR2X1_LOC_631/B 0.03fF
C7667 AND2X1_LOC_59/Y OR2X1_LOC_219/B 0.05fF
C7668 OR2X1_LOC_440/A OR2X1_LOC_733/A 0.04fF
C7669 OR2X1_LOC_124/A AND2X1_LOC_667/a_36_24# 0.01fF
C7670 INPUT_5 AND2X1_LOC_21/a_8_24# 0.09fF
C7671 OR2X1_LOC_413/Y OR2X1_LOC_7/A 0.14fF
C7672 OR2X1_LOC_865/Y OR2X1_LOC_269/B 0.00fF
C7673 OR2X1_LOC_391/B OR2X1_LOC_772/a_8_216# 0.02fF
C7674 OR2X1_LOC_158/A OR2X1_LOC_51/a_8_216# 0.02fF
C7675 OR2X1_LOC_604/A OR2X1_LOC_96/a_36_216# 0.01fF
C7676 OR2X1_LOC_683/a_8_216# OR2X1_LOC_683/Y -0.00fF
C7677 OR2X1_LOC_773/B AND2X1_LOC_3/Y 0.01fF
C7678 OR2X1_LOC_699/a_8_216# OR2X1_LOC_820/B 0.01fF
C7679 OR2X1_LOC_377/A OR2X1_LOC_3/Y 0.28fF
C7680 OR2X1_LOC_174/A OR2X1_LOC_814/A 0.02fF
C7681 OR2X1_LOC_809/B AND2X1_LOC_47/Y 0.05fF
C7682 AND2X1_LOC_70/Y OR2X1_LOC_439/a_36_216# 0.00fF
C7683 AND2X1_LOC_111/a_8_24# OR2X1_LOC_161/A 0.03fF
C7684 AND2X1_LOC_191/B AND2X1_LOC_859/B 0.02fF
C7685 OR2X1_LOC_140/A OR2X1_LOC_473/A 0.37fF
C7686 OR2X1_LOC_318/A OR2X1_LOC_318/B 0.23fF
C7687 OR2X1_LOC_154/A OR2X1_LOC_688/a_8_216# 0.01fF
C7688 OR2X1_LOC_744/A AND2X1_LOC_863/Y 0.07fF
C7689 OR2X1_LOC_81/Y OR2X1_LOC_26/Y 0.05fF
C7690 OR2X1_LOC_435/a_8_216# OR2X1_LOC_814/A 0.07fF
C7691 AND2X1_LOC_81/B AND2X1_LOC_3/Y 0.03fF
C7692 AND2X1_LOC_647/Y OR2X1_LOC_16/A 0.01fF
C7693 OR2X1_LOC_6/B AND2X1_LOC_838/B 0.02fF
C7694 AND2X1_LOC_560/B OR2X1_LOC_52/B 0.10fF
C7695 OR2X1_LOC_502/A AND2X1_LOC_672/B 0.03fF
C7696 AND2X1_LOC_81/B OR2X1_LOC_647/B 0.01fF
C7697 AND2X1_LOC_3/Y OR2X1_LOC_358/B 0.03fF
C7698 OR2X1_LOC_97/A AND2X1_LOC_31/Y 0.10fF
C7699 OR2X1_LOC_482/Y AND2X1_LOC_483/Y 0.00fF
C7700 OR2X1_LOC_149/B OR2X1_LOC_546/A 0.13fF
C7701 OR2X1_LOC_690/A OR2X1_LOC_52/B 0.06fF
C7702 AND2X1_LOC_598/a_8_24# OR2X1_LOC_485/A 0.02fF
C7703 OR2X1_LOC_3/Y OR2X1_LOC_85/A 0.05fF
C7704 OR2X1_LOC_743/A OR2X1_LOC_6/A 0.03fF
C7705 AND2X1_LOC_537/Y AND2X1_LOC_654/Y 0.07fF
C7706 AND2X1_LOC_67/Y OR2X1_LOC_375/A 0.12fF
C7707 OR2X1_LOC_612/B AND2X1_LOC_610/a_36_24# 0.00fF
C7708 OR2X1_LOC_329/B OR2X1_LOC_760/a_8_216# 0.05fF
C7709 AND2X1_LOC_559/a_8_24# OR2X1_LOC_74/A 0.07fF
C7710 OR2X1_LOC_485/A OR2X1_LOC_26/Y 0.74fF
C7711 VDD AND2X1_LOC_647/B 0.03fF
C7712 OR2X1_LOC_214/B OR2X1_LOC_66/A 0.02fF
C7713 OR2X1_LOC_195/A OR2X1_LOC_269/B 0.03fF
C7714 OR2X1_LOC_64/Y OR2X1_LOC_67/A 0.03fF
C7715 OR2X1_LOC_473/a_8_216# OR2X1_LOC_532/B 0.01fF
C7716 OR2X1_LOC_613/Y OR2X1_LOC_617/Y 0.03fF
C7717 OR2X1_LOC_813/a_8_216# OR2X1_LOC_86/A 0.00fF
C7718 OR2X1_LOC_66/A OR2X1_LOC_241/B 0.54fF
C7719 OR2X1_LOC_665/Y OR2X1_LOC_89/A 0.01fF
C7720 AND2X1_LOC_70/Y AND2X1_LOC_418/a_8_24# 0.01fF
C7721 OR2X1_LOC_485/A AND2X1_LOC_493/a_8_24# 0.01fF
C7722 AND2X1_LOC_343/a_36_24# OR2X1_LOC_585/A 0.00fF
C7723 OR2X1_LOC_280/a_8_216# OR2X1_LOC_280/Y 0.01fF
C7724 OR2X1_LOC_151/A OR2X1_LOC_854/A 0.01fF
C7725 OR2X1_LOC_481/A OR2X1_LOC_44/Y 0.03fF
C7726 OR2X1_LOC_441/Y AND2X1_LOC_811/Y 0.13fF
C7727 OR2X1_LOC_631/B OR2X1_LOC_778/A 0.00fF
C7728 AND2X1_LOC_227/Y OR2X1_LOC_265/a_8_216# 0.01fF
C7729 AND2X1_LOC_349/B OR2X1_LOC_485/A 0.00fF
C7730 OR2X1_LOC_485/A OR2X1_LOC_89/A 1.49fF
C7731 AND2X1_LOC_553/A AND2X1_LOC_866/A 0.03fF
C7732 AND2X1_LOC_259/Y AND2X1_LOC_345/a_8_24# 0.10fF
C7733 AND2X1_LOC_86/B AND2X1_LOC_85/a_36_24# 0.00fF
C7734 OR2X1_LOC_696/Y OR2X1_LOC_591/a_8_216# 0.57fF
C7735 OR2X1_LOC_813/A OR2X1_LOC_71/a_36_216# 0.00fF
C7736 AND2X1_LOC_792/a_36_24# AND2X1_LOC_789/Y 0.01fF
C7737 OR2X1_LOC_125/Y OR2X1_LOC_6/A 0.01fF
C7738 OR2X1_LOC_154/A OR2X1_LOC_403/a_8_216# 0.05fF
C7739 OR2X1_LOC_231/A OR2X1_LOC_218/Y 0.16fF
C7740 OR2X1_LOC_243/A D_INPUT_0 0.00fF
C7741 OR2X1_LOC_377/A AND2X1_LOC_53/Y 0.01fF
C7742 D_INPUT_5 OR2X1_LOC_17/a_8_216# 0.01fF
C7743 OR2X1_LOC_246/A OR2X1_LOC_6/A 0.01fF
C7744 AND2X1_LOC_7/Y AND2X1_LOC_43/B 0.04fF
C7745 OR2X1_LOC_64/Y OR2X1_LOC_52/B 0.32fF
C7746 AND2X1_LOC_798/A OR2X1_LOC_92/Y 0.03fF
C7747 AND2X1_LOC_76/a_8_24# OR2X1_LOC_75/Y 0.00fF
C7748 AND2X1_LOC_59/Y OR2X1_LOC_244/A 0.03fF
C7749 OR2X1_LOC_354/a_8_216# OR2X1_LOC_356/B 0.03fF
C7750 OR2X1_LOC_36/Y AND2X1_LOC_633/Y 0.02fF
C7751 OR2X1_LOC_160/A AND2X1_LOC_47/Y 0.14fF
C7752 OR2X1_LOC_600/A AND2X1_LOC_793/B 0.00fF
C7753 OR2X1_LOC_316/Y OR2X1_LOC_31/Y 0.07fF
C7754 AND2X1_LOC_489/Y OR2X1_LOC_64/Y 0.02fF
C7755 OR2X1_LOC_225/a_8_216# OR2X1_LOC_6/A 0.18fF
C7756 OR2X1_LOC_600/A OR2X1_LOC_533/A 0.16fF
C7757 OR2X1_LOC_36/Y D_INPUT_0 0.37fF
C7758 OR2X1_LOC_164/Y OR2X1_LOC_419/Y 0.05fF
C7759 AND2X1_LOC_703/a_36_24# OR2X1_LOC_47/Y 0.00fF
C7760 OR2X1_LOC_71/Y OR2X1_LOC_44/Y 0.03fF
C7761 OR2X1_LOC_602/a_8_216# AND2X1_LOC_51/Y 0.01fF
C7762 OR2X1_LOC_377/A OR2X1_LOC_673/A 0.03fF
C7763 OR2X1_LOC_302/B AND2X1_LOC_31/Y 0.00fF
C7764 OR2X1_LOC_51/Y OR2X1_LOC_534/Y 0.00fF
C7765 OR2X1_LOC_834/A OR2X1_LOC_779/B 0.17fF
C7766 OR2X1_LOC_808/B OR2X1_LOC_365/B 0.03fF
C7767 OR2X1_LOC_252/Y OR2X1_LOC_615/Y 0.02fF
C7768 AND2X1_LOC_722/Y AND2X1_LOC_222/Y 0.01fF
C7769 OR2X1_LOC_541/A AND2X1_LOC_31/Y 0.01fF
C7770 OR2X1_LOC_78/A OR2X1_LOC_724/A 0.07fF
C7771 OR2X1_LOC_256/a_36_216# AND2X1_LOC_721/A 0.00fF
C7772 AND2X1_LOC_566/Y AND2X1_LOC_477/A 0.00fF
C7773 OR2X1_LOC_404/A AND2X1_LOC_79/Y 0.80fF
C7774 OR2X1_LOC_561/Y OR2X1_LOC_561/B 0.00fF
C7775 OR2X1_LOC_574/A AND2X1_LOC_69/a_36_24# 0.06fF
C7776 AND2X1_LOC_41/A OR2X1_LOC_560/A 0.25fF
C7777 OR2X1_LOC_776/a_8_216# OR2X1_LOC_228/Y 0.01fF
C7778 AND2X1_LOC_41/A OR2X1_LOC_198/A 0.04fF
C7779 AND2X1_LOC_42/B OR2X1_LOC_720/B 0.03fF
C7780 AND2X1_LOC_784/Y OR2X1_LOC_142/Y 0.03fF
C7781 AND2X1_LOC_537/Y AND2X1_LOC_307/a_8_24# 0.06fF
C7782 OR2X1_LOC_599/A AND2X1_LOC_648/B 0.00fF
C7783 AND2X1_LOC_489/Y OR2X1_LOC_417/A 0.20fF
C7784 AND2X1_LOC_126/a_8_24# OR2X1_LOC_68/B 0.00fF
C7785 AND2X1_LOC_22/Y OR2X1_LOC_115/B 0.02fF
C7786 OR2X1_LOC_779/Y OR2X1_LOC_779/a_8_216# 0.00fF
C7787 AND2X1_LOC_40/Y OR2X1_LOC_742/B 0.14fF
C7788 AND2X1_LOC_86/B AND2X1_LOC_47/Y 0.01fF
C7789 AND2X1_LOC_31/Y OR2X1_LOC_475/B 0.03fF
C7790 AND2X1_LOC_554/B OR2X1_LOC_95/Y 0.03fF
C7791 OR2X1_LOC_485/A OR2X1_LOC_92/a_8_216# 0.01fF
C7792 OR2X1_LOC_297/Y AND2X1_LOC_866/A 0.04fF
C7793 OR2X1_LOC_160/A OR2X1_LOC_598/A 0.30fF
C7794 VDD OR2X1_LOC_771/B 1.94fF
C7795 OR2X1_LOC_624/B AND2X1_LOC_47/Y 1.06fF
C7796 OR2X1_LOC_272/Y AND2X1_LOC_656/Y 0.40fF
C7797 OR2X1_LOC_40/Y OR2X1_LOC_386/a_8_216# 0.03fF
C7798 OR2X1_LOC_604/A OR2X1_LOC_183/a_8_216# 0.30fF
C7799 OR2X1_LOC_363/A OR2X1_LOC_580/A 0.04fF
C7800 OR2X1_LOC_653/Y OR2X1_LOC_228/Y 0.02fF
C7801 AND2X1_LOC_675/Y OR2X1_LOC_437/A 0.08fF
C7802 OR2X1_LOC_40/Y OR2X1_LOC_183/Y 0.00fF
C7803 VDD OR2X1_LOC_209/A 0.04fF
C7804 OR2X1_LOC_59/Y OR2X1_LOC_300/Y 0.08fF
C7805 OR2X1_LOC_12/Y AND2X1_LOC_772/Y 0.28fF
C7806 OR2X1_LOC_755/A OR2X1_LOC_417/A 0.00fF
C7807 AND2X1_LOC_592/Y OR2X1_LOC_696/A 0.02fF
C7808 OR2X1_LOC_89/A AND2X1_LOC_645/a_36_24# 0.00fF
C7809 OR2X1_LOC_6/B OR2X1_LOC_130/Y 0.02fF
C7810 OR2X1_LOC_18/a_8_216# OR2X1_LOC_428/A 0.01fF
C7811 OR2X1_LOC_161/B OR2X1_LOC_161/a_8_216# 0.03fF
C7812 VDD OR2X1_LOC_776/A 0.16fF
C7813 AND2X1_LOC_835/a_8_24# OR2X1_LOC_54/Y 0.00fF
C7814 OR2X1_LOC_516/B OR2X1_LOC_437/A 0.03fF
C7815 OR2X1_LOC_167/Y AND2X1_LOC_727/A 0.00fF
C7816 OR2X1_LOC_45/B OR2X1_LOC_135/a_8_216# 0.01fF
C7817 AND2X1_LOC_64/Y OR2X1_LOC_786/A 0.03fF
C7818 OR2X1_LOC_485/A OR2X1_LOC_419/a_8_216# 0.01fF
C7819 OR2X1_LOC_176/Y AND2X1_LOC_212/Y 0.04fF
C7820 AND2X1_LOC_3/Y OR2X1_LOC_66/Y 0.01fF
C7821 OR2X1_LOC_291/a_36_216# OR2X1_LOC_71/A 0.01fF
C7822 OR2X1_LOC_615/a_8_216# OR2X1_LOC_47/Y 0.01fF
C7823 OR2X1_LOC_846/B D_INPUT_1 0.02fF
C7824 AND2X1_LOC_564/A AND2X1_LOC_477/Y 0.07fF
C7825 AND2X1_LOC_787/A AND2X1_LOC_794/B 0.01fF
C7826 OR2X1_LOC_22/Y AND2X1_LOC_476/A 0.07fF
C7827 OR2X1_LOC_272/a_8_216# AND2X1_LOC_216/A 0.03fF
C7828 OR2X1_LOC_326/B OR2X1_LOC_532/Y 0.01fF
C7829 OR2X1_LOC_167/Y OR2X1_LOC_95/Y 0.01fF
C7830 OR2X1_LOC_603/Y AND2X1_LOC_605/a_8_24# 0.23fF
C7831 AND2X1_LOC_318/Y INPUT_1 0.00fF
C7832 AND2X1_LOC_477/Y AND2X1_LOC_727/B 0.11fF
C7833 OR2X1_LOC_188/Y OR2X1_LOC_66/A 0.00fF
C7834 OR2X1_LOC_121/Y OR2X1_LOC_151/A 0.07fF
C7835 OR2X1_LOC_275/A OR2X1_LOC_595/Y 0.81fF
C7836 OR2X1_LOC_217/a_36_216# OR2X1_LOC_560/A 0.00fF
C7837 AND2X1_LOC_43/B OR2X1_LOC_515/a_8_216# 0.01fF
C7838 OR2X1_LOC_696/A AND2X1_LOC_512/Y 0.07fF
C7839 AND2X1_LOC_244/A AND2X1_LOC_860/A 0.05fF
C7840 AND2X1_LOC_392/A OR2X1_LOC_428/A 0.07fF
C7841 AND2X1_LOC_787/A VDD 0.28fF
C7842 OR2X1_LOC_106/Y OR2X1_LOC_59/Y 0.03fF
C7843 OR2X1_LOC_542/B OR2X1_LOC_577/Y 0.03fF
C7844 OR2X1_LOC_64/Y AND2X1_LOC_216/A 0.00fF
C7845 OR2X1_LOC_710/B AND2X1_LOC_44/Y 0.13fF
C7846 AND2X1_LOC_392/A OR2X1_LOC_595/A 0.07fF
C7847 AND2X1_LOC_92/a_8_24# AND2X1_LOC_92/Y 0.01fF
C7848 OR2X1_LOC_628/Y AND2X1_LOC_483/Y 0.86fF
C7849 OR2X1_LOC_701/Y AND2X1_LOC_789/Y -0.02fF
C7850 AND2X1_LOC_48/A AND2X1_LOC_761/a_8_24# 0.03fF
C7851 AND2X1_LOC_810/Y AND2X1_LOC_812/a_8_24# 0.03fF
C7852 OR2X1_LOC_6/B OR2X1_LOC_158/A 0.03fF
C7853 OR2X1_LOC_709/A OR2X1_LOC_676/Y 0.01fF
C7854 AND2X1_LOC_596/a_8_24# AND2X1_LOC_771/B 0.01fF
C7855 AND2X1_LOC_713/Y OR2X1_LOC_158/A 0.00fF
C7856 OR2X1_LOC_693/a_8_216# VDD 0.21fF
C7857 OR2X1_LOC_40/Y OR2X1_LOC_309/a_8_216# 0.01fF
C7858 OR2X1_LOC_426/a_36_216# AND2X1_LOC_451/Y 0.00fF
C7859 AND2X1_LOC_715/Y AND2X1_LOC_512/Y 0.10fF
C7860 OR2X1_LOC_539/a_8_216# OR2X1_LOC_539/B 0.40fF
C7861 OR2X1_LOC_114/B OR2X1_LOC_151/A 0.00fF
C7862 AND2X1_LOC_402/a_8_24# OR2X1_LOC_397/Y 0.03fF
C7863 AND2X1_LOC_157/a_8_24# INPUT_6 0.01fF
C7864 OR2X1_LOC_715/B AND2X1_LOC_110/Y 0.03fF
C7865 AND2X1_LOC_357/A AND2X1_LOC_357/B 1.32fF
C7866 AND2X1_LOC_366/A OR2X1_LOC_428/A 0.25fF
C7867 AND2X1_LOC_857/Y OR2X1_LOC_321/a_8_216# 0.01fF
C7868 VDD AND2X1_LOC_566/B 0.01fF
C7869 OR2X1_LOC_502/A OR2X1_LOC_390/a_8_216# 0.03fF
C7870 AND2X1_LOC_93/a_8_24# OR2X1_LOC_66/A 0.01fF
C7871 AND2X1_LOC_12/Y AND2X1_LOC_581/a_8_24# 0.01fF
C7872 OR2X1_LOC_532/B AND2X1_LOC_485/a_8_24# 0.01fF
C7873 OR2X1_LOC_702/A OR2X1_LOC_446/B 0.01fF
C7874 AND2X1_LOC_463/B OR2X1_LOC_409/B 0.00fF
C7875 OR2X1_LOC_44/Y AND2X1_LOC_789/Y 0.09fF
C7876 INPUT_0 OR2X1_LOC_9/a_8_216# 0.08fF
C7877 OR2X1_LOC_87/A OR2X1_LOC_469/B 0.01fF
C7878 AND2X1_LOC_22/Y OR2X1_LOC_840/A 0.03fF
C7879 OR2X1_LOC_663/A AND2X1_LOC_44/Y 0.04fF
C7880 OR2X1_LOC_496/Y OR2X1_LOC_142/Y 0.03fF
C7881 OR2X1_LOC_630/a_36_216# OR2X1_LOC_140/B 0.00fF
C7882 AND2X1_LOC_729/Y OR2X1_LOC_144/a_8_216# 0.01fF
C7883 OR2X1_LOC_499/B OR2X1_LOC_161/B 0.01fF
C7884 INPUT_0 OR2X1_LOC_13/a_8_216# 0.01fF
C7885 OR2X1_LOC_160/A OR2X1_LOC_186/a_8_216# 0.04fF
C7886 OR2X1_LOC_136/Y AND2X1_LOC_364/A 0.02fF
C7887 OR2X1_LOC_51/Y AND2X1_LOC_500/B 0.03fF
C7888 OR2X1_LOC_630/B OR2X1_LOC_549/A 0.01fF
C7889 AND2X1_LOC_64/Y OR2X1_LOC_624/A 0.05fF
C7890 OR2X1_LOC_121/Y AND2X1_LOC_67/a_8_24# 0.23fF
C7891 OR2X1_LOC_403/B AND2X1_LOC_36/Y 0.03fF
C7892 OR2X1_LOC_279/Y OR2X1_LOC_437/A 0.19fF
C7893 VDD OR2X1_LOC_695/Y 0.16fF
C7894 OR2X1_LOC_151/A OR2X1_LOC_538/A 0.08fF
C7895 AND2X1_LOC_724/Y AND2X1_LOC_447/Y 0.05fF
C7896 OR2X1_LOC_78/A OR2X1_LOC_631/A 0.02fF
C7897 OR2X1_LOC_309/Y OR2X1_LOC_744/A 0.03fF
C7898 OR2X1_LOC_177/Y OR2X1_LOC_164/Y 0.03fF
C7899 OR2X1_LOC_158/A AND2X1_LOC_335/a_8_24# 0.05fF
C7900 AND2X1_LOC_658/B AND2X1_LOC_188/a_8_24# 0.03fF
C7901 OR2X1_LOC_494/Y AND2X1_LOC_558/a_8_24# 0.09fF
C7902 AND2X1_LOC_218/a_8_24# OR2X1_LOC_59/Y 0.01fF
C7903 OR2X1_LOC_71/Y AND2X1_LOC_570/a_8_24# 0.03fF
C7904 OR2X1_LOC_254/B OR2X1_LOC_562/A 0.12fF
C7905 AND2X1_LOC_363/Y AND2X1_LOC_367/B 0.21fF
C7906 OR2X1_LOC_7/A OR2X1_LOC_183/Y 0.35fF
C7907 AND2X1_LOC_354/Y OR2X1_LOC_428/A 0.05fF
C7908 AND2X1_LOC_322/a_8_24# OR2X1_LOC_538/A 0.01fF
C7909 OR2X1_LOC_547/B AND2X1_LOC_44/Y 0.02fF
C7910 OR2X1_LOC_31/Y OR2X1_LOC_153/a_8_216# 0.01fF
C7911 OR2X1_LOC_375/A OR2X1_LOC_259/A 0.01fF
C7912 AND2X1_LOC_738/B AND2X1_LOC_657/Y 0.10fF
C7913 AND2X1_LOC_181/a_8_24# OR2X1_LOC_600/A 0.01fF
C7914 OR2X1_LOC_622/a_8_216# AND2X1_LOC_36/Y 0.01fF
C7915 AND2X1_LOC_620/Y AND2X1_LOC_793/Y 0.07fF
C7916 AND2X1_LOC_520/Y AND2X1_LOC_786/Y 0.05fF
C7917 OR2X1_LOC_175/Y OR2X1_LOC_169/B 0.01fF
C7918 AND2X1_LOC_647/B OR2X1_LOC_67/Y 0.06fF
C7919 OR2X1_LOC_78/A AND2X1_LOC_616/a_8_24# 0.07fF
C7920 VDD OR2X1_LOC_678/a_8_216# 0.00fF
C7921 AND2X1_LOC_528/a_36_24# AND2X1_LOC_36/Y 0.01fF
C7922 AND2X1_LOC_191/B OR2X1_LOC_56/A 0.07fF
C7923 OR2X1_LOC_166/Y AND2X1_LOC_436/Y 0.01fF
C7924 OR2X1_LOC_323/A OR2X1_LOC_372/Y 0.01fF
C7925 AND2X1_LOC_658/A OR2X1_LOC_59/Y 0.07fF
C7926 OR2X1_LOC_56/A AND2X1_LOC_469/B 0.02fF
C7927 AND2X1_LOC_43/B OR2X1_LOC_375/a_8_216# 0.04fF
C7928 OR2X1_LOC_335/A OR2X1_LOC_269/B 0.14fF
C7929 AND2X1_LOC_539/Y OR2X1_LOC_36/Y 0.03fF
C7930 OR2X1_LOC_240/B OR2X1_LOC_633/A 0.01fF
C7931 AND2X1_LOC_537/Y OR2X1_LOC_13/B 0.01fF
C7932 OR2X1_LOC_604/A OR2X1_LOC_164/Y 0.07fF
C7933 OR2X1_LOC_404/Y OR2X1_LOC_523/A 0.16fF
C7934 AND2X1_LOC_514/a_36_24# OR2X1_LOC_426/B 0.01fF
C7935 AND2X1_LOC_12/Y OR2X1_LOC_318/A 0.01fF
C7936 OR2X1_LOC_787/Y OR2X1_LOC_605/Y 0.01fF
C7937 OR2X1_LOC_264/Y OR2X1_LOC_641/A 0.04fF
C7938 AND2X1_LOC_72/B OR2X1_LOC_493/Y 0.03fF
C7939 AND2X1_LOC_794/B AND2X1_LOC_532/a_8_24# 0.06fF
C7940 OR2X1_LOC_560/a_8_216# OR2X1_LOC_113/B 0.01fF
C7941 OR2X1_LOC_40/Y AND2X1_LOC_840/a_8_24# 0.02fF
C7942 OR2X1_LOC_78/A OR2X1_LOC_632/Y 0.02fF
C7943 OR2X1_LOC_485/A AND2X1_LOC_590/a_8_24# 0.16fF
C7944 OR2X1_LOC_680/A AND2X1_LOC_785/Y 0.09fF
C7945 AND2X1_LOC_544/Y OR2X1_LOC_52/B 0.05fF
C7946 AND2X1_LOC_785/A OR2X1_LOC_70/Y 0.06fF
C7947 AND2X1_LOC_594/a_36_24# AND2X1_LOC_95/Y 0.01fF
C7948 AND2X1_LOC_66/a_8_24# OR2X1_LOC_13/B 0.04fF
C7949 OR2X1_LOC_110/a_8_216# OR2X1_LOC_74/A 0.06fF
C7950 OR2X1_LOC_296/a_36_216# OR2X1_LOC_140/B 0.00fF
C7951 OR2X1_LOC_160/B OR2X1_LOC_623/B 0.07fF
C7952 AND2X1_LOC_733/Y OR2X1_LOC_56/A 0.46fF
C7953 AND2X1_LOC_244/A AND2X1_LOC_287/Y 0.00fF
C7954 VDD OR2X1_LOC_637/B 0.21fF
C7955 OR2X1_LOC_185/Y AND2X1_LOC_44/Y 0.12fF
C7956 AND2X1_LOC_721/Y AND2X1_LOC_806/A 0.02fF
C7957 OR2X1_LOC_40/Y AND2X1_LOC_804/Y 0.03fF
C7958 OR2X1_LOC_519/Y OR2X1_LOC_158/A 0.01fF
C7959 AND2X1_LOC_170/B AND2X1_LOC_212/a_8_24# 0.04fF
C7960 AND2X1_LOC_378/a_8_24# INPUT_0 0.01fF
C7961 OR2X1_LOC_447/a_8_216# OR2X1_LOC_596/A 0.01fF
C7962 OR2X1_LOC_278/Y AND2X1_LOC_243/Y 0.80fF
C7963 AND2X1_LOC_555/Y OR2X1_LOC_3/Y 0.50fF
C7964 OR2X1_LOC_6/B OR2X1_LOC_847/A 0.02fF
C7965 VDD OR2X1_LOC_808/a_8_216# 0.00fF
C7966 OR2X1_LOC_864/A OR2X1_LOC_97/A 0.03fF
C7967 AND2X1_LOC_12/Y OR2X1_LOC_151/A 0.92fF
C7968 OR2X1_LOC_160/A OR2X1_LOC_646/B 0.11fF
C7969 OR2X1_LOC_374/Y OR2X1_LOC_723/A 0.02fF
C7970 OR2X1_LOC_158/A AND2X1_LOC_436/B 0.65fF
C7971 AND2X1_LOC_412/a_8_24# AND2X1_LOC_44/Y 0.02fF
C7972 AND2X1_LOC_564/B AND2X1_LOC_717/B 0.10fF
C7973 AND2X1_LOC_714/a_8_24# OR2X1_LOC_44/Y 0.02fF
C7974 OR2X1_LOC_272/Y AND2X1_LOC_772/Y 0.11fF
C7975 AND2X1_LOC_807/Y AND2X1_LOC_476/Y 0.02fF
C7976 OR2X1_LOC_158/A AND2X1_LOC_139/B 0.07fF
C7977 VDD AND2X1_LOC_11/Y 0.90fF
C7978 OR2X1_LOC_136/Y OR2X1_LOC_3/Y 0.05fF
C7979 OR2X1_LOC_154/A AND2X1_LOC_83/a_36_24# 0.00fF
C7980 AND2X1_LOC_797/A AND2X1_LOC_213/a_8_24# 0.20fF
C7981 OR2X1_LOC_858/A OR2X1_LOC_629/Y 0.03fF
C7982 OR2X1_LOC_494/Y OR2X1_LOC_18/Y 0.05fF
C7983 OR2X1_LOC_634/A OR2X1_LOC_640/A 0.01fF
C7984 VDD OR2X1_LOC_402/Y 0.62fF
C7985 AND2X1_LOC_765/a_8_24# AND2X1_LOC_3/Y 0.02fF
C7986 AND2X1_LOC_363/Y OR2X1_LOC_18/Y 0.02fF
C7987 OR2X1_LOC_696/A OR2X1_LOC_54/Y 0.14fF
C7988 AND2X1_LOC_711/Y AND2X1_LOC_726/a_8_24# 0.04fF
C7989 OR2X1_LOC_152/Y AND2X1_LOC_726/a_36_24# 0.00fF
C7990 OR2X1_LOC_280/Y AND2X1_LOC_445/a_8_24# 0.23fF
C7991 OR2X1_LOC_680/A AND2X1_LOC_500/B 0.02fF
C7992 AND2X1_LOC_712/a_36_24# OR2X1_LOC_7/A 0.01fF
C7993 OR2X1_LOC_185/A OR2X1_LOC_787/B 0.67fF
C7994 AND2X1_LOC_520/Y AND2X1_LOC_218/Y 0.82fF
C7995 AND2X1_LOC_301/a_8_24# OR2X1_LOC_316/Y 0.01fF
C7996 OR2X1_LOC_203/Y AND2X1_LOC_275/a_36_24# 0.01fF
C7997 AND2X1_LOC_110/a_8_24# OR2X1_LOC_161/A 0.02fF
C7998 OR2X1_LOC_186/Y AND2X1_LOC_528/a_8_24# 0.07fF
C7999 OR2X1_LOC_482/Y AND2X1_LOC_806/A 0.03fF
C8000 OR2X1_LOC_774/Y D_GATE_662 0.25fF
C8001 OR2X1_LOC_185/A AND2X1_LOC_92/Y 0.11fF
C8002 OR2X1_LOC_9/Y OR2X1_LOC_6/a_8_216# 0.03fF
C8003 OR2X1_LOC_167/a_8_216# OR2X1_LOC_485/A 0.01fF
C8004 INPUT_5 AND2X1_LOC_752/a_8_24# 0.10fF
C8005 AND2X1_LOC_847/Y OR2X1_LOC_59/Y 0.01fF
C8006 OR2X1_LOC_671/a_8_216# OR2X1_LOC_85/A 0.01fF
C8007 D_INPUT_5 OR2X1_LOC_651/B 0.01fF
C8008 AND2X1_LOC_773/Y OR2X1_LOC_273/Y 0.12fF
C8009 VDD OR2X1_LOC_642/a_8_216# 0.21fF
C8010 OR2X1_LOC_502/A AND2X1_LOC_402/a_36_24# 0.00fF
C8011 OR2X1_LOC_326/B OR2X1_LOC_325/A 0.52fF
C8012 OR2X1_LOC_224/a_8_216# OR2X1_LOC_183/Y 0.01fF
C8013 OR2X1_LOC_158/A OR2X1_LOC_529/Y 0.03fF
C8014 OR2X1_LOC_216/A OR2X1_LOC_737/A 0.01fF
C8015 AND2X1_LOC_326/B OR2X1_LOC_36/Y 0.03fF
C8016 AND2X1_LOC_729/Y AND2X1_LOC_663/A 0.05fF
C8017 OR2X1_LOC_154/A OR2X1_LOC_648/A 0.08fF
C8018 OR2X1_LOC_539/a_8_216# OR2X1_LOC_78/B 0.01fF
C8019 OR2X1_LOC_185/Y OR2X1_LOC_785/a_8_216# 0.05fF
C8020 OR2X1_LOC_585/A AND2X1_LOC_200/a_8_24# 0.01fF
C8021 AND2X1_LOC_64/Y OR2X1_LOC_447/Y 0.01fF
C8022 OR2X1_LOC_137/a_8_216# OR2X1_LOC_137/B 0.02fF
C8023 OR2X1_LOC_426/B OR2X1_LOC_44/Y 0.24fF
C8024 AND2X1_LOC_48/A OR2X1_LOC_855/A 0.09fF
C8025 AND2X1_LOC_774/a_8_24# OR2X1_LOC_64/Y 0.17fF
C8026 AND2X1_LOC_486/Y AND2X1_LOC_787/a_8_24# 0.05fF
C8027 VDD OR2X1_LOC_217/a_8_216# 0.21fF
C8028 OR2X1_LOC_43/A AND2X1_LOC_436/Y 0.01fF
C8029 OR2X1_LOC_379/Y OR2X1_LOC_637/A 0.01fF
C8030 AND2X1_LOC_464/Y AND2X1_LOC_786/Y 0.02fF
C8031 OR2X1_LOC_502/A AND2X1_LOC_278/a_8_24# 0.08fF
C8032 OR2X1_LOC_744/A AND2X1_LOC_840/B 0.05fF
C8033 AND2X1_LOC_862/a_8_24# OR2X1_LOC_56/A 0.03fF
C8034 OR2X1_LOC_296/Y OR2X1_LOC_629/B 0.00fF
C8035 OR2X1_LOC_347/a_8_216# OR2X1_LOC_811/A 0.13fF
C8036 OR2X1_LOC_377/A OR2X1_LOC_502/A 0.07fF
C8037 OR2X1_LOC_40/Y AND2X1_LOC_345/Y 0.00fF
C8038 OR2X1_LOC_189/Y OR2X1_LOC_679/Y 0.14fF
C8039 OR2X1_LOC_604/A AND2X1_LOC_155/Y 0.01fF
C8040 OR2X1_LOC_303/A OR2X1_LOC_468/Y 0.09fF
C8041 OR2X1_LOC_318/B OR2X1_LOC_716/a_8_216# 0.01fF
C8042 OR2X1_LOC_477/Y OR2X1_LOC_467/a_8_216# 0.01fF
C8043 OR2X1_LOC_49/A OR2X1_LOC_62/B 0.03fF
C8044 OR2X1_LOC_840/A AND2X1_LOC_153/a_8_24# 0.02fF
C8045 AND2X1_LOC_41/A OR2X1_LOC_267/a_8_216# 0.01fF
C8046 AND2X1_LOC_392/A AND2X1_LOC_211/a_8_24# 0.04fF
C8047 AND2X1_LOC_711/Y OR2X1_LOC_505/Y 0.08fF
C8048 OR2X1_LOC_3/Y OR2X1_LOC_815/a_36_216# 0.03fF
C8049 AND2X1_LOC_709/a_8_24# OR2X1_LOC_258/Y 0.24fF
C8050 AND2X1_LOC_36/Y OR2X1_LOC_493/Y 0.06fF
C8051 OR2X1_LOC_152/Y OR2X1_LOC_679/Y 0.01fF
C8052 OR2X1_LOC_298/a_8_216# OR2X1_LOC_6/A 0.02fF
C8053 AND2X1_LOC_702/a_8_24# OR2X1_LOC_48/B 0.01fF
C8054 OR2X1_LOC_45/B OR2X1_LOC_71/Y 0.04fF
C8055 OR2X1_LOC_528/Y AND2X1_LOC_663/B 0.00fF
C8056 AND2X1_LOC_36/Y OR2X1_LOC_801/B 0.10fF
C8057 OR2X1_LOC_196/Y AND2X1_LOC_47/Y 0.01fF
C8058 OR2X1_LOC_3/Y OR2X1_LOC_51/Y 0.21fF
C8059 VDD OR2X1_LOC_817/Y 0.12fF
C8060 AND2X1_LOC_378/a_8_24# OR2X1_LOC_690/A 0.08fF
C8061 OR2X1_LOC_632/a_8_216# OR2X1_LOC_574/A 0.02fF
C8062 OR2X1_LOC_833/a_8_216# AND2X1_LOC_56/B 0.01fF
C8063 AND2X1_LOC_47/Y OR2X1_LOC_266/A 0.01fF
C8064 AND2X1_LOC_711/Y AND2X1_LOC_658/A 0.01fF
C8065 AND2X1_LOC_736/Y AND2X1_LOC_565/Y 0.14fF
C8066 OR2X1_LOC_70/Y AND2X1_LOC_658/A 0.03fF
C8067 OR2X1_LOC_74/Y OR2X1_LOC_85/A 0.01fF
C8068 OR2X1_LOC_160/A OR2X1_LOC_506/A 0.10fF
C8069 OR2X1_LOC_31/Y AND2X1_LOC_639/B 0.04fF
C8070 AND2X1_LOC_120/a_8_24# OR2X1_LOC_666/A 0.01fF
C8071 AND2X1_LOC_571/Y AND2X1_LOC_572/Y 0.12fF
C8072 OR2X1_LOC_19/B AND2X1_LOC_243/Y 0.07fF
C8073 AND2X1_LOC_319/A OR2X1_LOC_427/A 0.03fF
C8074 AND2X1_LOC_564/A GATE_811 0.03fF
C8075 OR2X1_LOC_682/a_8_216# OR2X1_LOC_92/Y 0.03fF
C8076 AND2X1_LOC_858/B OR2X1_LOC_279/a_36_216# 0.01fF
C8077 AND2X1_LOC_756/a_36_24# AND2X1_LOC_711/Y 0.01fF
C8078 OR2X1_LOC_598/A OR2X1_LOC_130/Y 0.10fF
C8079 AND2X1_LOC_722/Y OR2X1_LOC_74/A 0.05fF
C8080 OR2X1_LOC_154/A OR2X1_LOC_405/a_8_216# 0.02fF
C8081 AND2X1_LOC_64/Y OR2X1_LOC_84/Y 0.06fF
C8082 AND2X1_LOC_384/a_8_24# OR2X1_LOC_269/B 0.01fF
C8083 OR2X1_LOC_160/A AND2X1_LOC_129/a_8_24# 0.01fF
C8084 OR2X1_LOC_400/A OR2X1_LOC_377/A 0.02fF
C8085 AND2X1_LOC_95/Y OR2X1_LOC_468/Y 0.03fF
C8086 AND2X1_LOC_855/a_8_24# AND2X1_LOC_434/Y 0.02fF
C8087 AND2X1_LOC_553/A OR2X1_LOC_7/A 0.00fF
C8088 OR2X1_LOC_529/Y OR2X1_LOC_103/Y 0.01fF
C8089 OR2X1_LOC_494/A AND2X1_LOC_721/A 0.00fF
C8090 AND2X1_LOC_47/Y OR2X1_LOC_768/a_8_216# 0.01fF
C8091 AND2X1_LOC_580/A OR2X1_LOC_39/A 0.06fF
C8092 OR2X1_LOC_45/B D_INPUT_1 0.02fF
C8093 OR2X1_LOC_812/B OR2X1_LOC_269/B 0.03fF
C8094 OR2X1_LOC_417/A OR2X1_LOC_253/Y 0.04fF
C8095 OR2X1_LOC_95/Y AND2X1_LOC_476/Y 0.22fF
C8096 AND2X1_LOC_362/B OR2X1_LOC_95/Y 0.01fF
C8097 AND2X1_LOC_629/Y OR2X1_LOC_627/Y 0.00fF
C8098 OR2X1_LOC_36/Y OR2X1_LOC_237/a_8_216# 0.01fF
C8099 AND2X1_LOC_847/Y OR2X1_LOC_820/B 0.01fF
C8100 OR2X1_LOC_3/Y OR2X1_LOC_16/Y 0.34fF
C8101 OR2X1_LOC_391/B OR2X1_LOC_846/a_8_216# 0.09fF
C8102 OR2X1_LOC_368/A AND2X1_LOC_476/Y 0.05fF
C8103 OR2X1_LOC_504/Y OR2X1_LOC_505/Y 0.01fF
C8104 AND2X1_LOC_550/A OR2X1_LOC_52/B 0.03fF
C8105 OR2X1_LOC_627/a_8_216# AND2X1_LOC_621/Y 0.06fF
C8106 D_INPUT_0 OR2X1_LOC_66/A 0.51fF
C8107 OR2X1_LOC_160/B OR2X1_LOC_544/A 0.00fF
C8108 AND2X1_LOC_382/a_8_24# OR2X1_LOC_848/A 0.02fF
C8109 OR2X1_LOC_406/Y OR2X1_LOC_406/A 0.01fF
C8110 OR2X1_LOC_794/a_8_216# OR2X1_LOC_794/A 0.18fF
C8111 OR2X1_LOC_91/A OR2X1_LOC_46/A 0.11fF
C8112 INPUT_0 OR2X1_LOC_22/Y 1.46fF
C8113 OR2X1_LOC_504/Y AND2X1_LOC_658/A 0.03fF
C8114 AND2X1_LOC_95/a_8_24# AND2X1_LOC_47/Y 0.01fF
C8115 OR2X1_LOC_604/A AND2X1_LOC_450/Y -0.00fF
C8116 AND2X1_LOC_571/A AND2X1_LOC_657/A 0.03fF
C8117 OR2X1_LOC_555/A OR2X1_LOC_555/B 0.04fF
C8118 AND2X1_LOC_379/a_8_24# OR2X1_LOC_588/Y 0.06fF
C8119 AND2X1_LOC_580/A AND2X1_LOC_569/a_8_24# 0.01fF
C8120 VDD AND2X1_LOC_675/A 0.82fF
C8121 AND2X1_LOC_61/a_8_24# OR2X1_LOC_31/Y 0.00fF
C8122 OR2X1_LOC_54/Y AND2X1_LOC_819/a_8_24# 0.01fF
C8123 OR2X1_LOC_280/a_8_216# OR2X1_LOC_39/A 0.04fF
C8124 AND2X1_LOC_59/Y OR2X1_LOC_643/a_8_216# 0.01fF
C8125 OR2X1_LOC_3/Y AND2X1_LOC_94/a_8_24# 0.01fF
C8126 OR2X1_LOC_728/B AND2X1_LOC_7/B 0.01fF
C8127 OR2X1_LOC_808/B OR2X1_LOC_121/B 0.04fF
C8128 OR2X1_LOC_306/a_8_216# OR2X1_LOC_485/A 0.03fF
C8129 AND2X1_LOC_311/a_8_24# D_INPUT_0 0.01fF
C8130 AND2X1_LOC_53/Y OR2X1_LOC_78/B 0.07fF
C8131 OR2X1_LOC_571/Y OR2X1_LOC_579/A 0.89fF
C8132 OR2X1_LOC_748/A OR2X1_LOC_701/a_8_216# 0.01fF
C8133 OR2X1_LOC_526/Y AND2X1_LOC_796/Y 0.00fF
C8134 OR2X1_LOC_175/Y AND2X1_LOC_31/Y 0.03fF
C8135 AND2X1_LOC_193/a_36_24# OR2X1_LOC_690/A 0.02fF
C8136 OR2X1_LOC_596/A AND2X1_LOC_39/Y 0.01fF
C8137 OR2X1_LOC_131/Y OR2X1_LOC_65/B 0.15fF
C8138 OR2X1_LOC_139/a_8_216# OR2X1_LOC_204/Y 0.00fF
C8139 OR2X1_LOC_45/Y OR2X1_LOC_431/a_8_216# 0.03fF
C8140 AND2X1_LOC_749/a_36_24# OR2X1_LOC_750/A 0.00fF
C8141 OR2X1_LOC_744/A OR2X1_LOC_31/Y 0.11fF
C8142 OR2X1_LOC_543/a_8_216# OR2X1_LOC_161/B 0.02fF
C8143 OR2X1_LOC_625/Y OR2X1_LOC_615/a_8_216# 0.01fF
C8144 AND2X1_LOC_352/B AND2X1_LOC_318/Y 0.06fF
C8145 AND2X1_LOC_93/a_8_24# OR2X1_LOC_98/B 0.01fF
C8146 OR2X1_LOC_663/A OR2X1_LOC_720/B 3.11fF
C8147 AND2X1_LOC_227/Y AND2X1_LOC_858/B 0.03fF
C8148 AND2X1_LOC_244/A AND2X1_LOC_562/Y 0.06fF
C8149 OR2X1_LOC_130/A OR2X1_LOC_33/B 0.02fF
C8150 OR2X1_LOC_248/a_8_216# OR2X1_LOC_7/A 0.01fF
C8151 AND2X1_LOC_597/a_36_24# OR2X1_LOC_155/A 0.01fF
C8152 AND2X1_LOC_227/Y OR2X1_LOC_91/A 0.03fF
C8153 AND2X1_LOC_41/A AND2X1_LOC_821/a_8_24# 0.03fF
C8154 AND2X1_LOC_576/Y OR2X1_LOC_239/Y 0.15fF
C8155 OR2X1_LOC_119/a_8_216# OR2X1_LOC_118/Y 0.01fF
C8156 AND2X1_LOC_224/a_36_24# OR2X1_LOC_68/B 0.00fF
C8157 OR2X1_LOC_691/Y AND2X1_LOC_31/Y 0.03fF
C8158 OR2X1_LOC_158/A OR2X1_LOC_598/A 0.10fF
C8159 AND2X1_LOC_300/a_8_24# OR2X1_LOC_318/B 0.01fF
C8160 OR2X1_LOC_680/A AND2X1_LOC_631/Y 0.03fF
C8161 OR2X1_LOC_6/A OR2X1_LOC_229/Y 0.01fF
C8162 OR2X1_LOC_485/A OR2X1_LOC_246/a_8_216# 0.01fF
C8163 OR2X1_LOC_702/A AND2X1_LOC_56/B 0.84fF
C8164 OR2X1_LOC_154/A AND2X1_LOC_136/a_8_24# 0.02fF
C8165 OR2X1_LOC_743/A OR2X1_LOC_44/Y 0.21fF
C8166 AND2X1_LOC_31/Y OR2X1_LOC_375/Y 0.01fF
C8167 OR2X1_LOC_636/B OR2X1_LOC_87/A 0.02fF
C8168 AND2X1_LOC_612/B AND2X1_LOC_612/a_8_24# 0.03fF
C8169 OR2X1_LOC_366/A OR2X1_LOC_580/A 0.04fF
C8170 AND2X1_LOC_342/Y AND2X1_LOC_663/B 0.07fF
C8171 OR2X1_LOC_7/A AND2X1_LOC_294/a_8_24# 0.04fF
C8172 AND2X1_LOC_95/Y AND2X1_LOC_134/a_8_24# 0.05fF
C8173 AND2X1_LOC_31/Y OR2X1_LOC_713/A 0.03fF
C8174 OR2X1_LOC_432/a_8_216# AND2X1_LOC_687/Y 0.18fF
C8175 OR2X1_LOC_18/Y AND2X1_LOC_116/B 0.01fF
C8176 OR2X1_LOC_91/Y AND2X1_LOC_523/Y 5.61fF
C8177 OR2X1_LOC_161/B OR2X1_LOC_348/B 0.09fF
C8178 OR2X1_LOC_275/a_36_216# AND2X1_LOC_139/B 0.01fF
C8179 OR2X1_LOC_574/A AND2X1_LOC_3/Y 0.03fF
C8180 OR2X1_LOC_846/a_8_216# OR2X1_LOC_846/A 0.14fF
C8181 AND2X1_LOC_355/a_8_24# AND2X1_LOC_337/B 0.20fF
C8182 OR2X1_LOC_377/A AND2X1_LOC_48/A 0.10fF
C8183 D_INPUT_7 AND2X1_LOC_21/Y 0.01fF
C8184 AND2X1_LOC_573/A OR2X1_LOC_46/A 0.08fF
C8185 AND2X1_LOC_727/a_36_24# OR2X1_LOC_152/A 0.00fF
C8186 OR2X1_LOC_600/A AND2X1_LOC_846/a_8_24# 0.01fF
C8187 AND2X1_LOC_95/Y OR2X1_LOC_471/Y 0.06fF
C8188 AND2X1_LOC_107/a_8_24# OR2X1_LOC_161/A 0.01fF
C8189 OR2X1_LOC_165/a_8_216# OR2X1_LOC_417/A 0.03fF
C8190 AND2X1_LOC_40/Y OR2X1_LOC_468/a_8_216# 0.01fF
C8191 OR2X1_LOC_496/a_8_216# OR2X1_LOC_406/A 0.02fF
C8192 OR2X1_LOC_503/A OR2X1_LOC_22/Y 0.01fF
C8193 OR2X1_LOC_22/Y OR2X1_LOC_11/Y 0.78fF
C8194 OR2X1_LOC_604/a_8_216# OR2X1_LOC_427/A 0.02fF
C8195 AND2X1_LOC_59/Y OR2X1_LOC_404/A 0.04fF
C8196 OR2X1_LOC_91/A OR2X1_LOC_813/Y 0.19fF
C8197 OR2X1_LOC_847/A AND2X1_LOC_47/Y 0.00fF
C8198 OR2X1_LOC_643/A OR2X1_LOC_844/Y 0.67fF
C8199 OR2X1_LOC_630/Y OR2X1_LOC_493/Y 0.10fF
C8200 OR2X1_LOC_36/Y AND2X1_LOC_687/A 0.04fF
C8201 OR2X1_LOC_112/B OR2X1_LOC_775/a_8_216# 0.47fF
C8202 AND2X1_LOC_838/Y INPUT_1 0.01fF
C8203 AND2X1_LOC_710/Y AND2X1_LOC_848/A 0.03fF
C8204 OR2X1_LOC_300/a_36_216# AND2X1_LOC_786/Y 0.01fF
C8205 OR2X1_LOC_160/A OR2X1_LOC_780/A 0.01fF
C8206 OR2X1_LOC_476/B AND2X1_LOC_8/Y 0.01fF
C8207 OR2X1_LOC_419/Y AND2X1_LOC_471/Y 0.59fF
C8208 AND2X1_LOC_53/Y OR2X1_LOC_375/A 0.44fF
C8209 AND2X1_LOC_560/B OR2X1_LOC_22/Y 0.09fF
C8210 AND2X1_LOC_95/Y OR2X1_LOC_222/a_8_216# 0.01fF
C8211 AND2X1_LOC_227/Y AND2X1_LOC_573/A 0.01fF
C8212 OR2X1_LOC_650/Y AND2X1_LOC_8/Y 0.27fF
C8213 OR2X1_LOC_859/B OR2X1_LOC_859/A 0.35fF
C8214 OR2X1_LOC_114/Y OR2X1_LOC_113/A 0.81fF
C8215 OR2X1_LOC_280/Y OR2X1_LOC_64/Y 0.03fF
C8216 OR2X1_LOC_22/Y OR2X1_LOC_690/A 0.40fF
C8217 OR2X1_LOC_18/Y AND2X1_LOC_270/a_36_24# 0.00fF
C8218 AND2X1_LOC_476/a_8_24# OR2X1_LOC_268/Y 0.01fF
C8219 OR2X1_LOC_401/a_8_216# AND2X1_LOC_3/Y 0.02fF
C8220 OR2X1_LOC_78/B AND2X1_LOC_609/a_8_24# 0.02fF
C8221 OR2X1_LOC_417/A AND2X1_LOC_286/Y 0.01fF
C8222 AND2X1_LOC_648/B AND2X1_LOC_644/Y 0.00fF
C8223 AND2X1_LOC_141/B AND2X1_LOC_663/B 0.10fF
C8224 OR2X1_LOC_92/Y AND2X1_LOC_644/a_8_24# 0.02fF
C8225 OR2X1_LOC_13/Y OR2X1_LOC_13/B 0.05fF
C8226 OR2X1_LOC_160/A OR2X1_LOC_227/Y 0.00fF
C8227 OR2X1_LOC_427/A AND2X1_LOC_721/A 0.03fF
C8228 OR2X1_LOC_424/a_8_216# AND2X1_LOC_648/B 0.48fF
C8229 OR2X1_LOC_31/Y AND2X1_LOC_840/B 0.20fF
C8230 AND2X1_LOC_18/Y AND2X1_LOC_268/a_8_24# 0.01fF
C8231 AND2X1_LOC_64/Y OR2X1_LOC_556/a_8_216# 0.01fF
C8232 OR2X1_LOC_160/A AND2X1_LOC_420/a_8_24# 0.00fF
C8233 AND2X1_LOC_306/a_8_24# OR2X1_LOC_779/B 0.01fF
C8234 OR2X1_LOC_673/A OR2X1_LOC_375/A 0.02fF
C8235 OR2X1_LOC_335/B OR2X1_LOC_787/Y 0.00fF
C8236 OR2X1_LOC_409/B OR2X1_LOC_44/Y 0.03fF
C8237 OR2X1_LOC_31/Y OR2X1_LOC_74/a_8_216# 0.02fF
C8238 OR2X1_LOC_47/Y AND2X1_LOC_633/a_8_24# 0.16fF
C8239 OR2X1_LOC_160/A D_INPUT_1 0.10fF
C8240 OR2X1_LOC_618/Y OR2X1_LOC_85/A 0.03fF
C8241 OR2X1_LOC_26/Y OR2X1_LOC_238/a_8_216# 0.01fF
C8242 AND2X1_LOC_737/a_8_24# AND2X1_LOC_222/Y 0.01fF
C8243 OR2X1_LOC_382/A AND2X1_LOC_789/Y 0.07fF
C8244 OR2X1_LOC_34/B AND2X1_LOC_51/Y 0.05fF
C8245 AND2X1_LOC_244/a_36_24# OR2X1_LOC_13/B 0.01fF
C8246 AND2X1_LOC_663/B OR2X1_LOC_54/Y 0.07fF
C8247 OR2X1_LOC_595/Y AND2X1_LOC_643/a_36_24# 0.01fF
C8248 OR2X1_LOC_497/a_8_216# OR2X1_LOC_184/Y 0.16fF
C8249 OR2X1_LOC_280/Y OR2X1_LOC_417/A 0.74fF
C8250 AND2X1_LOC_107/a_8_24# AND2X1_LOC_51/Y 0.03fF
C8251 OR2X1_LOC_202/a_8_216# OR2X1_LOC_814/A 0.03fF
C8252 OR2X1_LOC_22/Y OR2X1_LOC_64/Y 1.30fF
C8253 AND2X1_LOC_7/B OR2X1_LOC_338/A 0.34fF
C8254 OR2X1_LOC_511/Y OR2X1_LOC_511/a_8_216# -0.00fF
C8255 OR2X1_LOC_279/Y AND2X1_LOC_845/Y 0.16fF
C8256 AND2X1_LOC_40/Y OR2X1_LOC_344/a_8_216# 0.01fF
C8257 OR2X1_LOC_92/Y AND2X1_LOC_657/A 0.10fF
C8258 AND2X1_LOC_219/Y OR2X1_LOC_300/a_8_216# 0.03fF
C8259 OR2X1_LOC_66/A OR2X1_LOC_339/A 0.01fF
C8260 AND2X1_LOC_851/B OR2X1_LOC_238/Y 0.04fF
C8261 OR2X1_LOC_705/B OR2X1_LOC_375/A 0.53fF
C8262 VDD OR2X1_LOC_593/B 0.38fF
C8263 OR2X1_LOC_7/A AND2X1_LOC_648/B 0.03fF
C8264 OR2X1_LOC_151/A OR2X1_LOC_356/B 0.10fF
C8265 OR2X1_LOC_756/B OR2X1_LOC_366/Y 0.01fF
C8266 OR2X1_LOC_709/B AND2X1_LOC_64/Y 0.00fF
C8267 AND2X1_LOC_363/A AND2X1_LOC_721/A 0.00fF
C8268 OR2X1_LOC_45/B AND2X1_LOC_734/a_8_24# 0.16fF
C8269 OR2X1_LOC_118/Y OR2X1_LOC_88/a_36_216# 0.00fF
C8270 AND2X1_LOC_456/B OR2X1_LOC_437/A 0.04fF
C8271 AND2X1_LOC_291/a_36_24# OR2X1_LOC_598/A 0.00fF
C8272 OR2X1_LOC_802/a_8_216# OR2X1_LOC_446/B 0.01fF
C8273 OR2X1_LOC_696/A AND2X1_LOC_553/a_8_24# 0.00fF
C8274 OR2X1_LOC_17/Y OR2X1_LOC_587/a_8_216# 0.01fF
C8275 OR2X1_LOC_143/a_36_216# INPUT_2 0.03fF
C8276 OR2X1_LOC_43/A OR2X1_LOC_86/A 0.03fF
C8277 OR2X1_LOC_177/Y AND2X1_LOC_552/a_8_24# 0.01fF
C8278 OR2X1_LOC_54/a_8_216# OR2X1_LOC_54/Y 0.01fF
C8279 AND2X1_LOC_86/B D_INPUT_1 4.06fF
C8280 OR2X1_LOC_186/Y AND2X1_LOC_7/B 0.01fF
C8281 OR2X1_LOC_605/B OR2X1_LOC_223/A 0.00fF
C8282 OR2X1_LOC_665/Y AND2X1_LOC_792/Y 0.02fF
C8283 OR2X1_LOC_562/Y OR2X1_LOC_570/a_8_216# 0.02fF
C8284 OR2X1_LOC_65/B AND2X1_LOC_657/A 0.16fF
C8285 OR2X1_LOC_121/B OR2X1_LOC_218/Y 0.01fF
C8286 OR2X1_LOC_516/Y AND2X1_LOC_570/Y 0.03fF
C8287 OR2X1_LOC_523/B OR2X1_LOC_392/B 0.04fF
C8288 OR2X1_LOC_624/B D_INPUT_1 0.07fF
C8289 OR2X1_LOC_22/Y OR2X1_LOC_417/A 0.31fF
C8290 AND2X1_LOC_100/a_8_24# AND2X1_LOC_647/Y 0.09fF
C8291 AND2X1_LOC_101/B AND2X1_LOC_216/A 0.46fF
C8292 OR2X1_LOC_49/A OR2X1_LOC_15/a_36_216# 0.00fF
C8293 AND2X1_LOC_127/a_8_24# AND2X1_LOC_47/Y -0.00fF
C8294 AND2X1_LOC_3/Y AND2X1_LOC_761/a_8_24# 0.01fF
C8295 AND2X1_LOC_594/a_36_24# AND2X1_LOC_22/Y 0.00fF
C8296 OR2X1_LOC_89/Y AND2X1_LOC_243/Y 0.02fF
C8297 OR2X1_LOC_208/A OR2X1_LOC_66/A 0.04fF
C8298 OR2X1_LOC_40/Y AND2X1_LOC_465/A 0.02fF
C8299 AND2X1_LOC_754/a_8_24# AND2X1_LOC_22/Y 0.17fF
C8300 OR2X1_LOC_506/a_8_216# VDD 0.00fF
C8301 OR2X1_LOC_571/a_36_216# OR2X1_LOC_579/A 0.01fF
C8302 AND2X1_LOC_552/a_8_24# OR2X1_LOC_604/A 0.12fF
C8303 OR2X1_LOC_78/A OR2X1_LOC_168/Y 0.42fF
C8304 AND2X1_LOC_65/A OR2X1_LOC_161/B 0.03fF
C8305 OR2X1_LOC_156/a_8_216# VDD 0.00fF
C8306 OR2X1_LOC_329/a_8_216# OR2X1_LOC_16/A 0.01fF
C8307 OR2X1_LOC_12/Y OR2X1_LOC_421/Y 0.00fF
C8308 OR2X1_LOC_865/B OR2X1_LOC_571/Y 0.07fF
C8309 AND2X1_LOC_817/a_8_24# OR2X1_LOC_80/A 0.02fF
C8310 OR2X1_LOC_847/B OR2X1_LOC_68/B 0.05fF
C8311 AND2X1_LOC_56/B OR2X1_LOC_151/a_36_216# 0.03fF
C8312 OR2X1_LOC_600/A AND2X1_LOC_794/a_8_24# 0.01fF
C8313 OR2X1_LOC_600/A GATE_579 0.76fF
C8314 OR2X1_LOC_405/A OR2X1_LOC_777/B 0.11fF
C8315 OR2X1_LOC_188/Y OR2X1_LOC_190/A 1.02fF
C8316 OR2X1_LOC_696/A AND2X1_LOC_718/a_8_24# 0.02fF
C8317 AND2X1_LOC_199/A OR2X1_LOC_13/Y 0.01fF
C8318 OR2X1_LOC_154/A OR2X1_LOC_704/a_8_216# 0.04fF
C8319 AND2X1_LOC_339/Y VDD 0.01fF
C8320 OR2X1_LOC_842/A AND2X1_LOC_44/Y 0.00fF
C8321 OR2X1_LOC_45/B OR2X1_LOC_426/B 0.13fF
C8322 OR2X1_LOC_158/A OR2X1_LOC_672/a_8_216# 0.03fF
C8323 VDD OR2X1_LOC_414/Y 0.19fF
C8324 OR2X1_LOC_113/B OR2X1_LOC_768/a_36_216# 0.00fF
C8325 AND2X1_LOC_625/a_8_24# OR2X1_LOC_549/A 0.04fF
C8326 OR2X1_LOC_154/A OR2X1_LOC_112/A 0.11fF
C8327 AND2X1_LOC_810/Y AND2X1_LOC_796/Y 0.01fF
C8328 OR2X1_LOC_501/B OR2X1_LOC_563/A 0.46fF
C8329 OR2X1_LOC_541/A OR2X1_LOC_121/A 0.01fF
C8330 OR2X1_LOC_703/B OR2X1_LOC_535/a_8_216# 0.19fF
C8331 OR2X1_LOC_169/a_8_216# OR2X1_LOC_788/B 0.02fF
C8332 OR2X1_LOC_26/Y OR2X1_LOC_385/a_8_216# 0.03fF
C8333 AND2X1_LOC_65/a_8_24# OR2X1_LOC_392/B 0.11fF
C8334 OR2X1_LOC_468/Y OR2X1_LOC_788/B 0.03fF
C8335 OR2X1_LOC_212/A OR2X1_LOC_308/Y 0.00fF
C8336 INPUT_1 OR2X1_LOC_98/a_8_216# 0.18fF
C8337 OR2X1_LOC_744/A AND2X1_LOC_213/B 0.05fF
C8338 OR2X1_LOC_648/A OR2X1_LOC_435/A 0.13fF
C8339 AND2X1_LOC_363/a_8_24# AND2X1_LOC_363/Y 0.02fF
C8340 AND2X1_LOC_845/a_8_24# AND2X1_LOC_845/Y 0.00fF
C8341 OR2X1_LOC_278/a_8_216# OR2X1_LOC_71/A 0.03fF
C8342 OR2X1_LOC_506/A OR2X1_LOC_130/Y 0.09fF
C8343 AND2X1_LOC_737/Y AND2X1_LOC_544/Y 0.05fF
C8344 AND2X1_LOC_717/B OR2X1_LOC_437/A 0.14fF
C8345 OR2X1_LOC_528/Y AND2X1_LOC_565/B 0.02fF
C8346 OR2X1_LOC_598/Y OR2X1_LOC_66/A 0.23fF
C8347 OR2X1_LOC_185/A AND2X1_LOC_235/a_36_24# 0.01fF
C8348 OR2X1_LOC_160/B OR2X1_LOC_507/A 0.10fF
C8349 OR2X1_LOC_147/B OR2X1_LOC_563/A 0.07fF
C8350 OR2X1_LOC_66/A OR2X1_LOC_356/a_8_216# 0.05fF
C8351 OR2X1_LOC_177/Y AND2X1_LOC_471/Y 0.03fF
C8352 OR2X1_LOC_532/B OR2X1_LOC_723/A 0.01fF
C8353 OR2X1_LOC_8/Y OR2X1_LOC_96/Y 0.03fF
C8354 OR2X1_LOC_125/a_8_216# OR2X1_LOC_600/A 0.07fF
C8355 OR2X1_LOC_759/A AND2X1_LOC_709/a_8_24# 0.18fF
C8356 OR2X1_LOC_405/A OR2X1_LOC_831/B 0.07fF
C8357 OR2X1_LOC_615/Y AND2X1_LOC_623/a_8_24# 0.03fF
C8358 AND2X1_LOC_658/B OR2X1_LOC_505/Y 0.13fF
C8359 AND2X1_LOC_486/Y AND2X1_LOC_787/A 0.05fF
C8360 AND2X1_LOC_64/Y OR2X1_LOC_161/A 0.60fF
C8361 AND2X1_LOC_57/Y OR2X1_LOC_154/A 0.03fF
C8362 OR2X1_LOC_53/Y OR2X1_LOC_48/B 0.00fF
C8363 OR2X1_LOC_763/a_8_216# OR2X1_LOC_12/Y 0.01fF
C8364 AND2X1_LOC_444/a_8_24# AND2X1_LOC_477/Y 0.03fF
C8365 AND2X1_LOC_120/a_8_24# OR2X1_LOC_13/B 0.01fF
C8366 OR2X1_LOC_186/Y OR2X1_LOC_319/B 0.02fF
C8367 OR2X1_LOC_396/a_8_216# OR2X1_LOC_396/Y -0.00fF
C8368 OR2X1_LOC_786/Y OR2X1_LOC_66/a_8_216# 0.04fF
C8369 OR2X1_LOC_122/Y AND2X1_LOC_362/B 0.01fF
C8370 OR2X1_LOC_53/Y OR2X1_LOC_18/Y 0.03fF
C8371 OR2X1_LOC_261/Y AND2X1_LOC_789/Y 0.02fF
C8372 OR2X1_LOC_78/A OR2X1_LOC_777/a_36_216# 0.00fF
C8373 AND2X1_LOC_614/a_8_24# OR2X1_LOC_59/Y 0.06fF
C8374 OR2X1_LOC_790/A AND2X1_LOC_693/a_8_24# 0.09fF
C8375 AND2X1_LOC_658/B AND2X1_LOC_658/A 0.28fF
C8376 AND2X1_LOC_70/Y OR2X1_LOC_602/Y 0.01fF
C8377 AND2X1_LOC_646/a_8_24# AND2X1_LOC_647/B 0.01fF
C8378 OR2X1_LOC_106/Y AND2X1_LOC_124/a_8_24# 0.23fF
C8379 AND2X1_LOC_539/Y OR2X1_LOC_306/Y 0.02fF
C8380 OR2X1_LOC_6/B OR2X1_LOC_78/Y 0.11fF
C8381 OR2X1_LOC_696/A OR2X1_LOC_26/Y 2.03fF
C8382 OR2X1_LOC_186/Y OR2X1_LOC_318/Y 0.03fF
C8383 AND2X1_LOC_22/a_36_24# AND2X1_LOC_44/Y 0.00fF
C8384 AND2X1_LOC_190/a_8_24# OR2X1_LOC_59/Y 0.00fF
C8385 OR2X1_LOC_186/Y OR2X1_LOC_212/a_8_216# 0.03fF
C8386 OR2X1_LOC_12/Y OR2X1_LOC_278/Y 0.03fF
C8387 OR2X1_LOC_114/a_8_216# AND2X1_LOC_18/Y 0.02fF
C8388 OR2X1_LOC_130/A OR2X1_LOC_392/B 0.00fF
C8389 OR2X1_LOC_61/Y AND2X1_LOC_65/A 0.00fF
C8390 OR2X1_LOC_329/B OR2X1_LOC_51/Y 0.14fF
C8391 AND2X1_LOC_392/A AND2X1_LOC_512/Y 0.02fF
C8392 OR2X1_LOC_509/a_8_216# AND2X1_LOC_40/Y 0.01fF
C8393 AND2X1_LOC_81/B AND2X1_LOC_7/B 1.22fF
C8394 OR2X1_LOC_696/A OR2X1_LOC_89/A 0.28fF
C8395 AND2X1_LOC_445/a_8_24# OR2X1_LOC_39/A 0.03fF
C8396 AND2X1_LOC_715/Y AND2X1_LOC_598/a_8_24# 0.02fF
C8397 AND2X1_LOC_701/a_36_24# OR2X1_LOC_269/B 0.01fF
C8398 AND2X1_LOC_719/Y OR2X1_LOC_495/Y 0.01fF
C8399 OR2X1_LOC_497/Y OR2X1_LOC_184/a_8_216# 0.04fF
C8400 AND2X1_LOC_7/B OR2X1_LOC_358/B 0.73fF
C8401 OR2X1_LOC_40/Y OR2X1_LOC_265/a_8_216# 0.03fF
C8402 OR2X1_LOC_339/a_8_216# OR2X1_LOC_756/B 0.09fF
C8403 OR2X1_LOC_318/A AND2X1_LOC_59/Y 0.00fF
C8404 AND2X1_LOC_204/Y AND2X1_LOC_215/A 0.00fF
C8405 OR2X1_LOC_739/A OR2X1_LOC_740/B 0.03fF
C8406 OR2X1_LOC_175/Y OR2X1_LOC_809/a_8_216# 0.01fF
C8407 AND2X1_LOC_570/Y AND2X1_LOC_842/a_8_24# 0.01fF
C8408 OR2X1_LOC_863/a_8_216# AND2X1_LOC_22/Y 0.06fF
C8409 OR2X1_LOC_864/A OR2X1_LOC_175/Y 0.03fF
C8410 OR2X1_LOC_305/a_8_216# OR2X1_LOC_428/A 0.06fF
C8411 OR2X1_LOC_696/A OR2X1_LOC_824/a_36_216# 0.00fF
C8412 VDD OR2X1_LOC_92/Y 3.25fF
C8413 AND2X1_LOC_40/Y OR2X1_LOC_66/A 1.06fF
C8414 AND2X1_LOC_866/A OR2X1_LOC_384/Y 0.03fF
C8415 OR2X1_LOC_7/A AND2X1_LOC_465/A 0.75fF
C8416 OR2X1_LOC_121/B OR2X1_LOC_703/Y 0.27fF
C8417 OR2X1_LOC_175/Y AND2X1_LOC_385/a_36_24# 0.00fF
C8418 AND2X1_LOC_48/A OR2X1_LOC_539/B 0.02fF
C8419 OR2X1_LOC_160/B OR2X1_LOC_653/Y 0.07fF
C8420 OR2X1_LOC_802/Y AND2X1_LOC_417/a_36_24# 0.00fF
C8421 OR2X1_LOC_589/A AND2X1_LOC_655/A 0.02fF
C8422 OR2X1_LOC_539/a_36_216# OR2X1_LOC_390/A 0.01fF
C8423 AND2X1_LOC_59/Y OR2X1_LOC_151/A 0.17fF
C8424 AND2X1_LOC_555/Y AND2X1_LOC_345/a_36_24# 0.00fF
C8425 VDD AND2X1_LOC_492/a_8_24# 0.00fF
C8426 AND2X1_LOC_512/Y AND2X1_LOC_436/a_8_24# 0.03fF
C8427 OR2X1_LOC_499/B OR2X1_LOC_630/B 0.02fF
C8428 OR2X1_LOC_833/a_8_216# AND2X1_LOC_92/Y 0.01fF
C8429 OR2X1_LOC_269/B OR2X1_LOC_758/a_8_216# 0.01fF
C8430 OR2X1_LOC_7/A AND2X1_LOC_231/a_8_24# 0.03fF
C8431 AND2X1_LOC_3/Y OR2X1_LOC_855/A 0.00fF
C8432 OR2X1_LOC_665/Y OR2X1_LOC_816/A 0.03fF
C8433 AND2X1_LOC_47/Y OR2X1_LOC_544/B 0.09fF
C8434 AND2X1_LOC_474/Y OR2X1_LOC_816/A 0.14fF
C8435 OR2X1_LOC_502/A OR2X1_LOC_78/B 1.39fF
C8436 AND2X1_LOC_721/Y OR2X1_LOC_529/Y 0.02fF
C8437 OR2X1_LOC_355/B OR2X1_LOC_355/A 0.04fF
C8438 VDD OR2X1_LOC_257/a_8_216# 0.21fF
C8439 OR2X1_LOC_563/B OR2X1_LOC_577/Y 0.02fF
C8440 OR2X1_LOC_680/A AND2X1_LOC_477/Y 0.07fF
C8441 AND2X1_LOC_64/Y AND2X1_LOC_51/Y 10.19fF
C8442 AND2X1_LOC_3/Y AND2X1_LOC_627/a_8_24# 0.01fF
C8443 OR2X1_LOC_485/A OR2X1_LOC_816/A 3.42fF
C8444 OR2X1_LOC_40/Y OR2X1_LOC_237/Y 0.00fF
C8445 OR2X1_LOC_516/a_8_216# AND2X1_LOC_784/Y 0.14fF
C8446 AND2X1_LOC_716/Y OR2X1_LOC_310/Y 0.02fF
C8447 AND2X1_LOC_573/A AND2X1_LOC_403/a_8_24# 0.01fF
C8448 OR2X1_LOC_45/B OR2X1_LOC_743/A 0.29fF
C8449 OR2X1_LOC_537/A OR2X1_LOC_66/A 0.03fF
C8450 AND2X1_LOC_730/a_8_24# AND2X1_LOC_209/a_8_24# 0.23fF
C8451 VDD OR2X1_LOC_65/B 0.79fF
C8452 OR2X1_LOC_759/A AND2X1_LOC_624/A 0.03fF
C8453 OR2X1_LOC_450/A OR2X1_LOC_707/A 0.05fF
C8454 AND2X1_LOC_161/a_8_24# AND2X1_LOC_161/Y 0.01fF
C8455 OR2X1_LOC_449/B OR2X1_LOC_596/A 0.04fF
C8456 OR2X1_LOC_204/a_8_216# OR2X1_LOC_161/B 0.49fF
C8457 OR2X1_LOC_6/B OR2X1_LOC_748/A 0.14fF
C8458 OR2X1_LOC_87/Y OR2X1_LOC_66/A 0.16fF
C8459 OR2X1_LOC_139/A OR2X1_LOC_215/A 0.05fF
C8460 AND2X1_LOC_22/Y AND2X1_LOC_1/Y 0.00fF
C8461 AND2X1_LOC_523/a_36_24# OR2X1_LOC_744/A 0.01fF
C8462 AND2X1_LOC_12/Y OR2X1_LOC_287/A 0.03fF
C8463 AND2X1_LOC_605/Y OR2X1_LOC_427/A 0.01fF
C8464 AND2X1_LOC_720/Y AND2X1_LOC_721/a_8_24# 0.19fF
C8465 OR2X1_LOC_492/a_36_216# OR2X1_LOC_529/Y 0.00fF
C8466 AND2X1_LOC_773/Y OR2X1_LOC_275/A 0.16fF
C8467 AND2X1_LOC_512/Y AND2X1_LOC_354/Y 0.02fF
C8468 AND2X1_LOC_367/A OR2X1_LOC_109/Y 0.08fF
C8469 OR2X1_LOC_100/Y OR2X1_LOC_101/a_8_216# 0.00fF
C8470 OR2X1_LOC_482/Y OR2X1_LOC_529/Y 0.03fF
C8471 INPUT_0 OR2X1_LOC_39/A 0.40fF
C8472 VDD OR2X1_LOC_271/Y 0.28fF
C8473 OR2X1_LOC_491/a_8_216# OR2X1_LOC_485/A 0.01fF
C8474 INPUT_0 OR2X1_LOC_459/a_8_216# -0.00fF
C8475 OR2X1_LOC_96/Y OR2X1_LOC_672/Y 0.02fF
C8476 OR2X1_LOC_756/B OR2X1_LOC_624/A 0.03fF
C8477 OR2X1_LOC_196/B AND2X1_LOC_7/B 0.23fF
C8478 OR2X1_LOC_43/A AND2X1_LOC_200/a_36_24# 0.00fF
C8479 AND2X1_LOC_508/B AND2X1_LOC_806/A 0.00fF
C8480 OR2X1_LOC_532/B OR2X1_LOC_186/a_36_216# 0.00fF
C8481 OR2X1_LOC_863/B OR2X1_LOC_863/A 0.07fF
C8482 OR2X1_LOC_822/a_36_216# OR2X1_LOC_585/A 0.00fF
C8483 OR2X1_LOC_865/B OR2X1_LOC_392/A 0.02fF
C8484 OR2X1_LOC_62/B OR2X1_LOC_392/B 0.03fF
C8485 AND2X1_LOC_859/Y AND2X1_LOC_286/a_8_24# 0.01fF
C8486 OR2X1_LOC_49/A OR2X1_LOC_121/B 0.18fF
C8487 AND2X1_LOC_510/A OR2X1_LOC_44/Y 0.29fF
C8488 AND2X1_LOC_22/Y AND2X1_LOC_134/a_8_24# 0.03fF
C8489 OR2X1_LOC_519/a_8_216# AND2X1_LOC_716/Y 0.01fF
C8490 AND2X1_LOC_82/Y AND2X1_LOC_51/Y 0.02fF
C8491 AND2X1_LOC_94/a_8_24# OR2X1_LOC_502/A 0.01fF
C8492 AND2X1_LOC_537/Y OR2X1_LOC_428/A 0.07fF
C8493 OR2X1_LOC_45/B OR2X1_LOC_246/A 0.01fF
C8494 AND2X1_LOC_454/a_8_24# OR2X1_LOC_52/B 0.02fF
C8495 AND2X1_LOC_744/a_36_24# OR2X1_LOC_160/A 0.00fF
C8496 AND2X1_LOC_716/Y AND2X1_LOC_723/a_36_24# 0.01fF
C8497 OR2X1_LOC_561/Y OR2X1_LOC_579/B 0.00fF
C8498 OR2X1_LOC_158/A OR2X1_LOC_481/A 0.06fF
C8499 OR2X1_LOC_124/A OR2X1_LOC_864/A 0.03fF
C8500 OR2X1_LOC_512/A OR2X1_LOC_161/A 0.00fF
C8501 OR2X1_LOC_649/B AND2X1_LOC_19/Y 0.01fF
C8502 AND2X1_LOC_785/A OR2X1_LOC_47/Y 0.01fF
C8503 OR2X1_LOC_91/Y AND2X1_LOC_733/Y 0.03fF
C8504 OR2X1_LOC_599/A OR2X1_LOC_91/A 0.03fF
C8505 AND2X1_LOC_832/a_36_24# OR2X1_LOC_48/B 0.01fF
C8506 AND2X1_LOC_22/Y OR2X1_LOC_655/B 0.08fF
C8507 AND2X1_LOC_42/B AND2X1_LOC_18/Y 2.19fF
C8508 AND2X1_LOC_755/a_36_24# OR2X1_LOC_850/B 0.00fF
C8509 AND2X1_LOC_663/A OR2X1_LOC_52/B 0.04fF
C8510 OR2X1_LOC_502/A OR2X1_LOC_375/A 0.20fF
C8511 OR2X1_LOC_121/B OR2X1_LOC_596/A 2.49fF
C8512 AND2X1_LOC_588/a_8_24# AND2X1_LOC_21/Y 0.01fF
C8513 OR2X1_LOC_224/a_8_216# AND2X1_LOC_465/A 0.01fF
C8514 OR2X1_LOC_405/A OR2X1_LOC_493/A 0.08fF
C8515 OR2X1_LOC_124/A OR2X1_LOC_633/B 0.26fF
C8516 AND2X1_LOC_456/B AND2X1_LOC_348/Y 0.37fF
C8517 OR2X1_LOC_113/a_8_216# AND2X1_LOC_47/Y 0.01fF
C8518 OR2X1_LOC_154/A OR2X1_LOC_105/Y 0.01fF
C8519 OR2X1_LOC_400/B OR2X1_LOC_756/B 0.03fF
C8520 OR2X1_LOC_324/A OR2X1_LOC_739/A 0.01fF
C8521 OR2X1_LOC_160/A OR2X1_LOC_737/A 0.14fF
C8522 OR2X1_LOC_235/B OR2X1_LOC_720/a_8_216# 0.00fF
C8523 AND2X1_LOC_47/Y OR2X1_LOC_474/B 0.04fF
C8524 AND2X1_LOC_191/B OR2X1_LOC_757/Y 0.38fF
C8525 AND2X1_LOC_524/a_8_24# OR2X1_LOC_443/Y 0.23fF
C8526 OR2X1_LOC_447/A OR2X1_LOC_506/A 0.07fF
C8527 OR2X1_LOC_711/B AND2X1_LOC_698/a_8_24# 0.01fF
C8528 AND2X1_LOC_211/B INPUT_0 0.07fF
C8529 AND2X1_LOC_850/A AND2X1_LOC_806/A 0.03fF
C8530 OR2X1_LOC_837/Y AND2X1_LOC_472/B 0.17fF
C8531 AND2X1_LOC_456/B OR2X1_LOC_753/A 0.00fF
C8532 OR2X1_LOC_756/B OR2X1_LOC_552/a_8_216# 0.14fF
C8533 OR2X1_LOC_393/a_36_216# OR2X1_LOC_39/A 0.03fF
C8534 OR2X1_LOC_485/Y OR2X1_LOC_64/Y 0.28fF
C8535 AND2X1_LOC_456/B OR2X1_LOC_669/a_36_216# 0.00fF
C8536 OR2X1_LOC_160/A AND2X1_LOC_95/Y 0.22fF
C8537 OR2X1_LOC_858/A OR2X1_LOC_850/A 0.03fF
C8538 OR2X1_LOC_555/B OR2X1_LOC_161/A 0.24fF
C8539 OR2X1_LOC_402/B OR2X1_LOC_402/a_8_216# 0.02fF
C8540 OR2X1_LOC_757/A OR2X1_LOC_3/Y 0.09fF
C8541 OR2X1_LOC_31/Y AND2X1_LOC_464/A 0.01fF
C8542 OR2X1_LOC_516/Y OR2X1_LOC_406/A 0.07fF
C8543 OR2X1_LOC_467/B OR2X1_LOC_471/Y 0.09fF
C8544 OR2X1_LOC_527/Y AND2X1_LOC_657/Y 0.10fF
C8545 AND2X1_LOC_544/Y AND2X1_LOC_808/A 3.01fF
C8546 AND2X1_LOC_849/A AND2X1_LOC_860/A 0.13fF
C8547 OR2X1_LOC_604/A AND2X1_LOC_687/A 0.22fF
C8548 OR2X1_LOC_523/B OR2X1_LOC_532/B 0.01fF
C8549 AND2X1_LOC_726/a_8_24# OR2X1_LOC_47/Y 0.02fF
C8550 OR2X1_LOC_416/A AND2X1_LOC_415/a_8_24# 0.01fF
C8551 OR2X1_LOC_158/A OR2X1_LOC_71/Y 0.05fF
C8552 AND2X1_LOC_654/Y AND2X1_LOC_661/A 0.09fF
C8553 OR2X1_LOC_774/a_8_216# D_INPUT_1 0.01fF
C8554 OR2X1_LOC_427/A AND2X1_LOC_361/A 0.33fF
C8555 OR2X1_LOC_9/Y AND2X1_LOC_839/A 0.00fF
C8556 OR2X1_LOC_439/a_8_216# OR2X1_LOC_439/B 0.08fF
C8557 OR2X1_LOC_417/Y AND2X1_LOC_469/B 0.00fF
C8558 AND2X1_LOC_737/a_8_24# OR2X1_LOC_74/A 0.01fF
C8559 OR2X1_LOC_760/a_36_216# OR2X1_LOC_16/A 0.00fF
C8560 OR2X1_LOC_653/Y OR2X1_LOC_219/B 0.07fF
C8561 OR2X1_LOC_158/A AND2X1_LOC_462/Y 0.03fF
C8562 OR2X1_LOC_213/A OR2X1_LOC_375/A 0.00fF
C8563 OR2X1_LOC_476/B AND2X1_LOC_92/Y 0.10fF
C8564 AND2X1_LOC_717/a_8_24# OR2X1_LOC_26/Y 0.05fF
C8565 AND2X1_LOC_574/A AND2X1_LOC_657/Y 0.15fF
C8566 OR2X1_LOC_188/Y OR2X1_LOC_241/B 0.03fF
C8567 OR2X1_LOC_321/Y AND2X1_LOC_857/Y 0.02fF
C8568 AND2X1_LOC_389/a_8_24# OR2X1_LOC_92/Y 0.01fF
C8569 OR2X1_LOC_650/Y AND2X1_LOC_92/Y 0.16fF
C8570 OR2X1_LOC_271/Y OR2X1_LOC_315/Y 0.15fF
C8571 OR2X1_LOC_66/Y AND2X1_LOC_7/B 0.02fF
C8572 AND2X1_LOC_847/Y OR2X1_LOC_701/a_36_216# 0.01fF
C8573 OR2X1_LOC_800/A OR2X1_LOC_687/Y 0.09fF
C8574 AND2X1_LOC_560/B OR2X1_LOC_39/A 0.02fF
C8575 OR2X1_LOC_160/A OR2X1_LOC_99/Y 0.03fF
C8576 OR2X1_LOC_796/a_8_216# OR2X1_LOC_155/A 0.01fF
C8577 AND2X1_LOC_16/a_8_24# AND2X1_LOC_3/Y 0.10fF
C8578 OR2X1_LOC_693/a_36_216# AND2X1_LOC_648/B 0.00fF
C8579 AND2X1_LOC_57/Y OR2X1_LOC_198/A 0.17fF
C8580 AND2X1_LOC_48/A OR2X1_LOC_78/B 0.40fF
C8581 OR2X1_LOC_43/A AND2X1_LOC_655/A 1.03fF
C8582 AND2X1_LOC_461/a_8_24# AND2X1_LOC_219/A 0.03fF
C8583 AND2X1_LOC_70/Y OR2X1_LOC_602/B 0.01fF
C8584 OR2X1_LOC_45/Y OR2X1_LOC_485/A 0.23fF
C8585 OR2X1_LOC_685/B OR2X1_LOC_685/a_8_216# 0.07fF
C8586 OR2X1_LOC_690/A OR2X1_LOC_39/A 0.11fF
C8587 AND2X1_LOC_449/Y OR2X1_LOC_52/B 0.10fF
C8588 OR2X1_LOC_694/Y OR2X1_LOC_31/Y 0.09fF
C8589 OR2X1_LOC_756/B AND2X1_LOC_442/a_36_24# 0.01fF
C8590 OR2X1_LOC_808/A OR2X1_LOC_121/B 0.04fF
C8591 OR2X1_LOC_837/Y OR2X1_LOC_19/B 0.02fF
C8592 OR2X1_LOC_377/A AND2X1_LOC_3/Y 0.48fF
C8593 AND2X1_LOC_807/Y AND2X1_LOC_474/Y 0.03fF
C8594 OR2X1_LOC_377/A OR2X1_LOC_647/B 0.07fF
C8595 AND2X1_LOC_390/B AND2X1_LOC_809/A 0.04fF
C8596 OR2X1_LOC_109/Y OR2X1_LOC_74/A 0.11fF
C8597 AND2X1_LOC_529/a_8_24# OR2X1_LOC_62/B 0.01fF
C8598 OR2X1_LOC_158/A D_INPUT_1 0.81fF
C8599 AND2X1_LOC_246/a_8_24# OR2X1_LOC_342/B 0.01fF
C8600 AND2X1_LOC_95/Y OR2X1_LOC_624/B 0.04fF
C8601 OR2X1_LOC_680/Y AND2X1_LOC_621/Y 0.03fF
C8602 AND2X1_LOC_95/Y OR2X1_LOC_33/a_8_216# 0.01fF
C8603 AND2X1_LOC_35/a_8_24# OR2X1_LOC_24/Y 0.01fF
C8604 OR2X1_LOC_151/Y AND2X1_LOC_152/a_8_24# 0.01fF
C8605 OR2X1_LOC_589/A OR2X1_LOC_599/Y 0.03fF
C8606 OR2X1_LOC_467/A OR2X1_LOC_783/A 0.01fF
C8607 OR2X1_LOC_849/A OR2X1_LOC_643/A 0.03fF
C8608 OR2X1_LOC_545/A OR2X1_LOC_545/a_8_216# 0.47fF
C8609 OR2X1_LOC_182/a_8_216# OR2X1_LOC_469/B 0.40fF
C8610 OR2X1_LOC_185/Y OR2X1_LOC_793/B 0.21fF
C8611 OR2X1_LOC_312/Y AND2X1_LOC_661/A 0.03fF
C8612 OR2X1_LOC_203/Y AND2X1_LOC_3/Y 0.26fF
C8613 OR2X1_LOC_352/a_8_216# OR2X1_LOC_578/B 0.01fF
C8614 OR2X1_LOC_658/a_8_216# AND2X1_LOC_47/Y 0.01fF
C8615 OR2X1_LOC_91/A AND2X1_LOC_866/A 0.12fF
C8616 AND2X1_LOC_658/A OR2X1_LOC_47/Y 0.12fF
C8617 OR2X1_LOC_173/Y AND2X1_LOC_211/B 0.01fF
C8618 AND2X1_LOC_190/a_8_24# OR2X1_LOC_184/Y 0.11fF
C8619 OR2X1_LOC_610/Y AND2X1_LOC_612/a_8_24# 0.23fF
C8620 AND2X1_LOC_359/a_8_24# OR2X1_LOC_89/A 0.03fF
C8621 OR2X1_LOC_229/Y OR2X1_LOC_44/Y 0.02fF
C8622 OR2X1_LOC_3/Y AND2X1_LOC_359/B 0.23fF
C8623 OR2X1_LOC_262/a_8_216# OR2X1_LOC_74/A 0.06fF
C8624 OR2X1_LOC_64/Y OR2X1_LOC_39/A 0.10fF
C8625 AND2X1_LOC_319/A OR2X1_LOC_681/Y 0.01fF
C8626 OR2X1_LOC_403/A OR2X1_LOC_532/B 0.01fF
C8627 OR2X1_LOC_89/A OR2X1_LOC_89/a_8_216# 0.05fF
C8628 OR2X1_LOC_92/Y OR2X1_LOC_256/A 0.07fF
C8629 OR2X1_LOC_3/Y OR2X1_LOC_423/a_8_216# 0.01fF
C8630 OR2X1_LOC_32/B OR2X1_LOC_46/A 0.51fF
C8631 AND2X1_LOC_486/Y AND2X1_LOC_675/A 0.07fF
C8632 OR2X1_LOC_18/Y INPUT_1 0.21fF
C8633 AND2X1_LOC_576/Y AND2X1_LOC_842/B 0.02fF
C8634 AND2X1_LOC_48/A OR2X1_LOC_375/A 0.87fF
C8635 OR2X1_LOC_413/a_8_216# D_INPUT_0 0.06fF
C8636 AND2X1_LOC_851/A OR2X1_LOC_95/Y 0.03fF
C8637 OR2X1_LOC_600/A AND2X1_LOC_805/a_36_24# 0.00fF
C8638 OR2X1_LOC_246/A OR2X1_LOC_767/a_8_216# 0.16fF
C8639 OR2X1_LOC_45/B OR2X1_LOC_599/a_8_216# 0.02fF
C8640 OR2X1_LOC_837/Y OR2X1_LOC_838/B 0.07fF
C8641 AND2X1_LOC_663/B OR2X1_LOC_26/Y 0.09fF
C8642 OR2X1_LOC_121/B OR2X1_LOC_87/B 0.72fF
C8643 OR2X1_LOC_3/Y AND2X1_LOC_639/a_8_24# 0.02fF
C8644 AND2X1_LOC_581/a_8_24# AND2X1_LOC_582/B 0.01fF
C8645 AND2X1_LOC_556/a_36_24# OR2X1_LOC_47/Y 0.00fF
C8646 AND2X1_LOC_40/Y OR2X1_LOC_84/A 0.23fF
C8647 OR2X1_LOC_814/A AND2X1_LOC_251/a_8_24# 0.01fF
C8648 OR2X1_LOC_100/Y AND2X1_LOC_88/Y 0.01fF
C8649 OR2X1_LOC_272/a_36_216# OR2X1_LOC_272/Y 0.00fF
C8650 D_INPUT_0 OR2X1_LOC_265/Y 0.01fF
C8651 AND2X1_LOC_211/B OR2X1_LOC_64/Y 0.07fF
C8652 OR2X1_LOC_417/A OR2X1_LOC_39/A 0.07fF
C8653 OR2X1_LOC_278/A OR2X1_LOC_612/B 0.05fF
C8654 OR2X1_LOC_256/A OR2X1_LOC_65/B 0.02fF
C8655 AND2X1_LOC_663/B OR2X1_LOC_89/A 0.11fF
C8656 AND2X1_LOC_84/Y AND2X1_LOC_204/a_8_24# 0.01fF
C8657 OR2X1_LOC_600/A AND2X1_LOC_657/A 0.07fF
C8658 OR2X1_LOC_130/A OR2X1_LOC_532/B 0.21fF
C8659 AND2X1_LOC_866/A AND2X1_LOC_573/A 0.07fF
C8660 OR2X1_LOC_78/B OR2X1_LOC_398/a_8_216# 0.05fF
C8661 OR2X1_LOC_274/Y OR2X1_LOC_493/Y 0.25fF
C8662 OR2X1_LOC_92/Y OR2X1_LOC_67/Y 0.39fF
C8663 OR2X1_LOC_97/A AND2X1_LOC_36/Y 0.03fF
C8664 OR2X1_LOC_40/Y OR2X1_LOC_384/Y 0.01fF
C8665 OR2X1_LOC_7/Y OR2X1_LOC_52/B 0.01fF
C8666 OR2X1_LOC_59/Y OR2X1_LOC_72/Y 0.02fF
C8667 OR2X1_LOC_426/A OR2X1_LOC_581/a_8_216# 0.40fF
C8668 OR2X1_LOC_427/A OR2X1_LOC_430/Y 0.01fF
C8669 OR2X1_LOC_72/a_8_216# OR2X1_LOC_85/A 0.01fF
C8670 OR2X1_LOC_485/A AND2X1_LOC_727/A 0.03fF
C8671 AND2X1_LOC_31/Y OR2X1_LOC_778/B 0.42fF
C8672 OR2X1_LOC_847/A D_INPUT_1 0.20fF
C8673 OR2X1_LOC_427/a_36_216# AND2X1_LOC_451/Y 0.00fF
C8674 OR2X1_LOC_233/a_8_216# OR2X1_LOC_46/A 0.01fF
C8675 OR2X1_LOC_532/B AND2X1_LOC_292/a_8_24# 0.17fF
C8676 OR2X1_LOC_331/A OR2X1_LOC_533/A 0.15fF
C8677 AND2X1_LOC_514/Y OR2X1_LOC_417/a_8_216# 0.03fF
C8678 OR2X1_LOC_417/Y OR2X1_LOC_417/a_36_216# 0.00fF
C8679 OR2X1_LOC_680/A GATE_662 0.20fF
C8680 OR2X1_LOC_427/A AND2X1_LOC_795/Y 0.02fF
C8681 VDD OR2X1_LOC_317/B 0.03fF
C8682 OR2X1_LOC_185/Y OR2X1_LOC_506/B 0.11fF
C8683 OR2X1_LOC_206/A AND2X1_LOC_51/Y 0.01fF
C8684 AND2X1_LOC_211/B OR2X1_LOC_417/A 0.16fF
C8685 OR2X1_LOC_737/A OR2X1_LOC_717/a_8_216# 0.03fF
C8686 OR2X1_LOC_158/A AND2X1_LOC_789/Y 0.29fF
C8687 OR2X1_LOC_235/B OR2X1_LOC_80/A 0.11fF
C8688 AND2X1_LOC_71/a_8_24# OR2X1_LOC_68/B 0.02fF
C8689 OR2X1_LOC_6/B OR2X1_LOC_217/A 0.04fF
C8690 VDD OR2X1_LOC_580/A 0.12fF
C8691 OR2X1_LOC_65/B OR2X1_LOC_67/Y 0.05fF
C8692 OR2X1_LOC_95/Y AND2X1_LOC_474/Y 0.03fF
C8693 OR2X1_LOC_97/A OR2X1_LOC_334/A 0.01fF
C8694 AND2X1_LOC_748/a_8_24# OR2X1_LOC_801/B -0.01fF
C8695 OR2X1_LOC_691/Y AND2X1_LOC_760/a_8_24# 0.01fF
C8696 OR2X1_LOC_485/A OR2X1_LOC_95/Y 0.94fF
C8697 OR2X1_LOC_176/Y AND2X1_LOC_539/Y 0.00fF
C8698 AND2X1_LOC_600/a_8_24# AND2X1_LOC_51/Y 0.02fF
C8699 OR2X1_LOC_19/B AND2X1_LOC_671/a_8_24# 0.09fF
C8700 OR2X1_LOC_42/a_36_216# D_INPUT_1 0.03fF
C8701 INPUT_4 OR2X1_LOC_581/a_8_216# 0.00fF
C8702 AND2X1_LOC_74/a_8_24# AND2X1_LOC_31/Y 0.01fF
C8703 OR2X1_LOC_696/A AND2X1_LOC_552/A 0.03fF
C8704 OR2X1_LOC_267/Y OR2X1_LOC_576/A 0.74fF
C8705 AND2X1_LOC_135/a_36_24# D_INPUT_0 0.00fF
C8706 OR2X1_LOC_606/a_36_216# OR2X1_LOC_606/Y 0.00fF
C8707 OR2X1_LOC_43/A OR2X1_LOC_599/Y 0.31fF
C8708 AND2X1_LOC_787/A AND2X1_LOC_457/a_8_24# 0.11fF
C8709 OR2X1_LOC_167/a_8_216# AND2X1_LOC_715/Y 0.04fF
C8710 OR2X1_LOC_22/Y OR2X1_LOC_226/a_8_216# 0.02fF
C8711 OR2X1_LOC_639/B AND2X1_LOC_31/Y 0.13fF
C8712 OR2X1_LOC_617/Y AND2X1_LOC_663/a_36_24# 0.00fF
C8713 OR2X1_LOC_62/B OR2X1_LOC_532/B 0.34fF
C8714 OR2X1_LOC_64/Y OR2X1_LOC_760/a_8_216# 0.01fF
C8715 AND2X1_LOC_774/a_36_24# OR2X1_LOC_428/A 0.01fF
C8716 OR2X1_LOC_585/A AND2X1_LOC_228/a_8_24# 0.03fF
C8717 OR2X1_LOC_730/a_8_216# OR2X1_LOC_446/B 0.06fF
C8718 AND2X1_LOC_679/a_8_24# OR2X1_LOC_155/A 0.04fF
C8719 AND2X1_LOC_802/Y AND2X1_LOC_810/B 0.32fF
C8720 OR2X1_LOC_70/A AND2X1_LOC_637/Y 0.03fF
C8721 OR2X1_LOC_51/Y OR2X1_LOC_525/a_8_216# 0.01fF
C8722 AND2X1_LOC_285/a_8_24# OR2X1_LOC_428/A 0.08fF
C8723 AND2X1_LOC_46/a_8_24# D_INPUT_1 0.03fF
C8724 OR2X1_LOC_13/Y OR2X1_LOC_428/A 0.03fF
C8725 OR2X1_LOC_739/A OR2X1_LOC_728/A 0.01fF
C8726 OR2X1_LOC_532/B AND2X1_LOC_108/a_36_24# 0.01fF
C8727 AND2X1_LOC_31/Y OR2X1_LOC_722/a_8_216# 0.01fF
C8728 OR2X1_LOC_19/B AND2X1_LOC_827/a_36_24# 0.00fF
C8729 AND2X1_LOC_755/a_8_24# OR2X1_LOC_580/A 0.03fF
C8730 D_INPUT_4 D_INPUT_6 1.24fF
C8731 AND2X1_LOC_138/a_8_24# OR2X1_LOC_13/B 0.03fF
C8732 AND2X1_LOC_95/Y OR2X1_LOC_532/Y 0.02fF
C8733 VDD AND2X1_LOC_44/Y 1.80fF
C8734 OR2X1_LOC_19/B OR2X1_LOC_644/A -0.01fF
C8735 AND2X1_LOC_40/Y OR2X1_LOC_502/a_8_216# 0.01fF
C8736 AND2X1_LOC_290/a_8_24# AND2X1_LOC_36/Y 0.01fF
C8737 OR2X1_LOC_121/B OR2X1_LOC_374/Y 0.03fF
C8738 AND2X1_LOC_537/a_8_24# OR2X1_LOC_16/A 0.02fF
C8739 AND2X1_LOC_491/a_36_24# OR2X1_LOC_493/Y 0.00fF
C8740 OR2X1_LOC_427/A AND2X1_LOC_439/a_8_24# 0.03fF
C8741 OR2X1_LOC_269/a_8_216# AND2X1_LOC_36/Y 0.01fF
C8742 OR2X1_LOC_158/A OR2X1_LOC_108/a_8_216# 0.02fF
C8743 INPUT_0 OR2X1_LOC_855/A 0.01fF
C8744 D_INPUT_0 OR2X1_LOC_214/B 2.72fF
C8745 OR2X1_LOC_269/B OR2X1_LOC_558/a_8_216# 0.01fF
C8746 OR2X1_LOC_188/Y AND2X1_LOC_189/a_8_24# 0.00fF
C8747 AND2X1_LOC_41/A OR2X1_LOC_267/Y 0.01fF
C8748 OR2X1_LOC_542/B OR2X1_LOC_294/Y 0.03fF
C8749 VDD AND2X1_LOC_729/a_8_24# -0.00fF
C8750 AND2X1_LOC_794/B OR2X1_LOC_600/A 0.00fF
C8751 AND2X1_LOC_716/a_36_24# OR2X1_LOC_437/A 0.00fF
C8752 OR2X1_LOC_659/A OR2X1_LOC_392/B 0.10fF
C8753 OR2X1_LOC_66/A OR2X1_LOC_356/A 0.06fF
C8754 OR2X1_LOC_462/B OR2X1_LOC_771/B 0.05fF
C8755 OR2X1_LOC_335/A OR2X1_LOC_811/A 0.01fF
C8756 OR2X1_LOC_3/Y OR2X1_LOC_399/a_8_216# 0.01fF
C8757 OR2X1_LOC_158/A OR2X1_LOC_426/B 0.14fF
C8758 AND2X1_LOC_180/a_8_24# OR2X1_LOC_51/Y 0.01fF
C8759 OR2X1_LOC_744/A OR2X1_LOC_522/Y 0.07fF
C8760 OR2X1_LOC_814/A OR2X1_LOC_358/A 1.37fF
C8761 OR2X1_LOC_696/A OR2X1_LOC_306/a_8_216# 0.09fF
C8762 OR2X1_LOC_46/A AND2X1_LOC_222/Y 0.03fF
C8763 AND2X1_LOC_388/Y AND2X1_LOC_436/Y 0.06fF
C8764 AND2X1_LOC_571/A AND2X1_LOC_571/Y 0.26fF
C8765 AND2X1_LOC_471/Y AND2X1_LOC_212/Y 0.01fF
C8766 OR2X1_LOC_139/A OR2X1_LOC_475/a_8_216# 0.25fF
C8767 OR2X1_LOC_291/Y AND2X1_LOC_206/Y 0.17fF
C8768 AND2X1_LOC_41/A OR2X1_LOC_725/A 0.06fF
C8769 AND2X1_LOC_541/Y OR2X1_LOC_56/A 0.04fF
C8770 VDD OR2X1_LOC_600/A 1.35fF
C8771 OR2X1_LOC_46/A OR2X1_LOC_68/B 0.03fF
C8772 OR2X1_LOC_680/A OR2X1_LOC_525/a_8_216# 0.03fF
C8773 AND2X1_LOC_51/Y OR2X1_LOC_579/a_8_216# 0.01fF
C8774 OR2X1_LOC_294/Y OR2X1_LOC_736/A 0.00fF
C8775 OR2X1_LOC_659/A OR2X1_LOC_113/B 0.01fF
C8776 OR2X1_LOC_753/A OR2X1_LOC_395/Y 0.05fF
C8777 AND2X1_LOC_391/Y OR2X1_LOC_40/Y 0.01fF
C8778 OR2X1_LOC_40/Y AND2X1_LOC_858/B 0.18fF
C8779 OR2X1_LOC_604/A OR2X1_LOC_90/a_8_216# 0.06fF
C8780 OR2X1_LOC_40/Y OR2X1_LOC_91/A 0.27fF
C8781 OR2X1_LOC_186/Y AND2X1_LOC_331/a_8_24# 0.01fF
C8782 OR2X1_LOC_9/Y AND2X1_LOC_820/B 0.01fF
C8783 VDD AND2X1_LOC_296/a_8_24# 0.00fF
C8784 AND2X1_LOC_12/Y OR2X1_LOC_563/A 0.07fF
C8785 OR2X1_LOC_438/Y AND2X1_LOC_476/Y 0.02fF
C8786 OR2X1_LOC_160/A AND2X1_LOC_22/Y 0.12fF
C8787 AND2X1_LOC_341/a_8_24# OR2X1_LOC_18/Y 0.01fF
C8788 OR2X1_LOC_700/Y OR2X1_LOC_428/A 0.02fF
C8789 AND2X1_LOC_706/Y AND2X1_LOC_832/a_8_24# 0.02fF
C8790 OR2X1_LOC_151/A OR2X1_LOC_623/B 0.20fF
C8791 OR2X1_LOC_858/A AND2X1_LOC_245/a_8_24# 0.15fF
C8792 OR2X1_LOC_405/A OR2X1_LOC_161/B 0.10fF
C8793 OR2X1_LOC_139/A OR2X1_LOC_539/Y 0.03fF
C8794 OR2X1_LOC_244/Y OR2X1_LOC_632/Y 0.06fF
C8795 OR2X1_LOC_161/A OR2X1_LOC_342/A 0.02fF
C8796 AND2X1_LOC_305/a_8_24# OR2X1_LOC_713/A 0.00fF
C8797 OR2X1_LOC_604/A OR2X1_LOC_746/a_8_216# 0.01fF
C8798 OR2X1_LOC_91/Y AND2X1_LOC_804/A 0.25fF
C8799 OR2X1_LOC_663/A AND2X1_LOC_18/Y 0.10fF
C8800 AND2X1_LOC_542/a_8_24# OR2X1_LOC_427/A 0.04fF
C8801 AND2X1_LOC_91/B OR2X1_LOC_849/A 0.09fF
C8802 AND2X1_LOC_732/a_8_24# AND2X1_LOC_605/Y 0.01fF
C8803 OR2X1_LOC_207/B OR2X1_LOC_375/A 0.03fF
C8804 VDD AND2X1_LOC_862/Y 0.02fF
C8805 AND2X1_LOC_350/B OR2X1_LOC_265/Y 0.06fF
C8806 OR2X1_LOC_122/A AND2X1_LOC_474/A 0.01fF
C8807 OR2X1_LOC_87/A AND2X1_LOC_224/a_36_24# 0.00fF
C8808 OR2X1_LOC_345/Y OR2X1_LOC_375/A 0.16fF
C8809 AND2X1_LOC_354/a_8_24# AND2X1_LOC_802/Y 0.04fF
C8810 AND2X1_LOC_563/a_8_24# OR2X1_LOC_595/A 0.03fF
C8811 OR2X1_LOC_501/B OR2X1_LOC_632/Y 0.08fF
C8812 OR2X1_LOC_36/Y OR2X1_LOC_310/a_8_216# 0.04fF
C8813 OR2X1_LOC_852/a_36_216# AND2X1_LOC_824/B 0.00fF
C8814 VDD OR2X1_LOC_61/a_8_216# 0.00fF
C8815 OR2X1_LOC_833/Y OR2X1_LOC_805/A 0.02fF
C8816 AND2X1_LOC_40/Y OR2X1_LOC_190/A 1.00fF
C8817 OR2X1_LOC_53/Y OR2X1_LOC_585/A 0.05fF
C8818 OR2X1_LOC_124/Y OR2X1_LOC_572/a_8_216# 0.07fF
C8819 OR2X1_LOC_45/B OR2X1_LOC_497/Y 0.02fF
C8820 AND2X1_LOC_621/Y AND2X1_LOC_476/Y 0.07fF
C8821 OR2X1_LOC_325/Y OR2X1_LOC_502/A 0.01fF
C8822 OR2X1_LOC_179/a_8_216# OR2X1_LOC_744/A 0.02fF
C8823 AND2X1_LOC_59/Y AND2X1_LOC_300/a_8_24# 0.03fF
C8824 OR2X1_LOC_9/Y OR2X1_LOC_823/Y 0.01fF
C8825 OR2X1_LOC_18/Y AND2X1_LOC_778/Y 0.20fF
C8826 OR2X1_LOC_6/B OR2X1_LOC_185/A 0.14fF
C8827 OR2X1_LOC_856/B AND2X1_LOC_387/a_36_24# 0.01fF
C8828 OR2X1_LOC_574/A AND2X1_LOC_7/B 0.11fF
C8829 OR2X1_LOC_782/B OR2X1_LOC_160/Y 0.08fF
C8830 OR2X1_LOC_579/B OR2X1_LOC_343/a_8_216# 0.05fF
C8831 OR2X1_LOC_87/A OR2X1_LOC_160/Y 0.03fF
C8832 OR2X1_LOC_118/Y AND2X1_LOC_243/Y 0.04fF
C8833 OR2X1_LOC_40/Y AND2X1_LOC_573/A 0.09fF
C8834 AND2X1_LOC_810/Y OR2X1_LOC_13/B 0.05fF
C8835 OR2X1_LOC_589/A AND2X1_LOC_266/Y 0.15fF
C8836 OR2X1_LOC_375/A OR2X1_LOC_542/a_8_216# 0.01fF
C8837 OR2X1_LOC_158/A OR2X1_LOC_517/Y 0.08fF
C8838 VDD OR2X1_LOC_619/Y 1.53fF
C8839 AND2X1_LOC_737/Y AND2X1_LOC_663/A 0.30fF
C8840 AND2X1_LOC_729/Y OR2X1_LOC_421/A 0.02fF
C8841 OR2X1_LOC_84/a_8_216# OR2X1_LOC_71/A 0.01fF
C8842 OR2X1_LOC_769/B OR2X1_LOC_637/a_8_216# 0.47fF
C8843 AND2X1_LOC_91/B OR2X1_LOC_602/a_36_216# 0.01fF
C8844 OR2X1_LOC_625/Y AND2X1_LOC_658/A 0.42fF
C8845 OR2X1_LOC_600/A OR2X1_LOC_616/Y 0.83fF
C8846 INPUT_0 OR2X1_LOC_818/Y 0.02fF
C8847 AND2X1_LOC_843/Y AND2X1_LOC_858/B 0.01fF
C8848 AND2X1_LOC_43/B OR2X1_LOC_66/A 0.11fF
C8849 OR2X1_LOC_99/Y AND2X1_LOC_607/a_8_24# 0.01fF
C8850 AND2X1_LOC_648/B OR2X1_LOC_424/Y 0.02fF
C8851 OR2X1_LOC_493/B OR2X1_LOC_805/A 0.05fF
C8852 OR2X1_LOC_43/A OR2X1_LOC_382/a_8_216# 0.01fF
C8853 INPUT_0 AND2X1_LOC_16/a_8_24# 0.01fF
C8854 OR2X1_LOC_354/A OR2X1_LOC_502/A 0.04fF
C8855 AND2X1_LOC_73/a_8_24# OR2X1_LOC_185/A 0.02fF
C8856 OR2X1_LOC_364/A AND2X1_LOC_18/Y 0.78fF
C8857 OR2X1_LOC_663/a_36_216# AND2X1_LOC_3/Y 0.02fF
C8858 OR2X1_LOC_821/Y OR2X1_LOC_485/A 0.40fF
C8859 INPUT_0 AND2X1_LOC_278/a_8_24# 0.01fF
C8860 OR2X1_LOC_185/Y AND2X1_LOC_18/Y 0.20fF
C8861 AND2X1_LOC_50/Y AND2X1_LOC_40/Y 0.07fF
C8862 OR2X1_LOC_316/Y OR2X1_LOC_56/A 0.03fF
C8863 OR2X1_LOC_461/B OR2X1_LOC_461/A 0.32fF
C8864 OR2X1_LOC_121/B OR2X1_LOC_392/B 0.03fF
C8865 OR2X1_LOC_641/B OR2X1_LOC_68/B 0.01fF
C8866 OR2X1_LOC_377/A INPUT_0 0.25fF
C8867 OR2X1_LOC_457/B OR2X1_LOC_741/Y 0.00fF
C8868 AND2X1_LOC_10/a_8_24# OR2X1_LOC_161/B 0.01fF
C8869 AND2X1_LOC_580/A OR2X1_LOC_51/Y 0.03fF
C8870 OR2X1_LOC_135/a_8_216# OR2X1_LOC_304/Y 0.01fF
C8871 AND2X1_LOC_486/Y OR2X1_LOC_92/Y 0.00fF
C8872 AND2X1_LOC_724/Y OR2X1_LOC_599/A 0.33fF
C8873 AND2X1_LOC_392/A OR2X1_LOC_26/Y 0.03fF
C8874 OR2X1_LOC_405/A OR2X1_LOC_435/B 1.33fF
C8875 OR2X1_LOC_275/A OR2X1_LOC_12/Y 0.03fF
C8876 AND2X1_LOC_842/B AND2X1_LOC_244/A 0.01fF
C8877 AND2X1_LOC_802/B AND2X1_LOC_727/A 0.01fF
C8878 OR2X1_LOC_158/A OR2X1_LOC_743/A 0.10fF
C8879 AND2X1_LOC_480/A AND2X1_LOC_221/a_8_24# 0.20fF
C8880 OR2X1_LOC_154/A OR2X1_LOC_858/A 0.30fF
C8881 AND2X1_LOC_12/Y AND2X1_LOC_628/a_36_24# 0.00fF
C8882 OR2X1_LOC_380/a_8_216# OR2X1_LOC_44/Y 0.01fF
C8883 OR2X1_LOC_450/A OR2X1_LOC_449/B 0.46fF
C8884 INPUT_0 AND2X1_LOC_824/B 0.04fF
C8885 OR2X1_LOC_756/B OR2X1_LOC_161/A 0.18fF
C8886 OR2X1_LOC_251/Y OR2X1_LOC_600/A 0.30fF
C8887 OR2X1_LOC_18/Y OR2X1_LOC_517/A 0.15fF
C8888 OR2X1_LOC_161/A OR2X1_LOC_735/a_36_216# 0.00fF
C8889 AND2X1_LOC_354/B OR2X1_LOC_56/A 0.03fF
C8890 AND2X1_LOC_543/a_8_24# OR2X1_LOC_315/Y 0.08fF
C8891 OR2X1_LOC_325/A AND2X1_LOC_95/Y 0.16fF
C8892 VDD OR2X1_LOC_465/B -0.00fF
C8893 OR2X1_LOC_629/A OR2X1_LOC_629/B 0.39fF
C8894 OR2X1_LOC_421/A AND2X1_LOC_769/a_8_24# 0.01fF
C8895 AND2X1_LOC_508/A AND2X1_LOC_624/A 0.07fF
C8896 OR2X1_LOC_633/a_36_216# OR2X1_LOC_375/A 0.00fF
C8897 OR2X1_LOC_36/Y AND2X1_LOC_434/Y 0.08fF
C8898 OR2X1_LOC_621/A OR2X1_LOC_624/B 0.01fF
C8899 AND2X1_LOC_191/B AND2X1_LOC_806/A 0.03fF
C8900 INPUT_0 OR2X1_LOC_85/A 0.03fF
C8901 AND2X1_LOC_392/A OR2X1_LOC_89/A 0.03fF
C8902 OR2X1_LOC_295/Y OR2X1_LOC_428/A 0.04fF
C8903 OR2X1_LOC_36/Y AND2X1_LOC_219/Y 0.09fF
C8904 OR2X1_LOC_359/a_8_216# OR2X1_LOC_287/B 0.00fF
C8905 AND2X1_LOC_729/B OR2X1_LOC_13/a_36_216# 0.00fF
C8906 OR2X1_LOC_625/Y AND2X1_LOC_631/a_8_24# 0.00fF
C8907 OR2X1_LOC_18/Y AND2X1_LOC_651/a_36_24# 0.00fF
C8908 OR2X1_LOC_235/B OR2X1_LOC_6/A 1.01fF
C8909 OR2X1_LOC_405/A OR2X1_LOC_61/Y 0.10fF
C8910 OR2X1_LOC_521/Y OR2X1_LOC_18/Y 0.32fF
C8911 OR2X1_LOC_598/A OR2X1_LOC_217/A 0.01fF
C8912 AND2X1_LOC_721/Y OR2X1_LOC_71/Y 0.02fF
C8913 AND2X1_LOC_312/a_8_24# AND2X1_LOC_56/B 0.12fF
C8914 AND2X1_LOC_366/A OR2X1_LOC_26/Y 0.03fF
C8915 OR2X1_LOC_770/A OR2X1_LOC_770/a_8_216# 0.01fF
C8916 OR2X1_LOC_696/A OR2X1_LOC_588/A 0.04fF
C8917 AND2X1_LOC_340/Y INPUT_1 0.11fF
C8918 AND2X1_LOC_548/a_8_24# AND2X1_LOC_658/A 0.05fF
C8919 AND2X1_LOC_391/Y OR2X1_LOC_7/A 0.07fF
C8920 AND2X1_LOC_92/a_8_24# AND2X1_LOC_47/Y 0.01fF
C8921 AND2X1_LOC_572/Y OR2X1_LOC_427/A 0.07fF
C8922 OR2X1_LOC_158/A OR2X1_LOC_125/Y 0.00fF
C8923 AND2X1_LOC_95/Y OR2X1_LOC_288/a_8_216# 0.01fF
C8924 AND2X1_LOC_858/B OR2X1_LOC_7/A 0.49fF
C8925 AND2X1_LOC_3/Y OR2X1_LOC_78/B 1.04fF
C8926 AND2X1_LOC_59/Y AND2X1_LOC_482/a_8_24# 0.11fF
C8927 OR2X1_LOC_5/a_8_216# INPUT_2 0.05fF
C8928 OR2X1_LOC_826/a_8_216# OR2X1_LOC_600/A 0.01fF
C8929 OR2X1_LOC_91/A OR2X1_LOC_7/A 0.28fF
C8930 OR2X1_LOC_803/a_8_216# OR2X1_LOC_155/A 0.01fF
C8931 OR2X1_LOC_647/B OR2X1_LOC_78/B 0.07fF
C8932 OR2X1_LOC_158/A OR2X1_LOC_246/A 0.10fF
C8933 AND2X1_LOC_390/B OR2X1_LOC_56/A 0.14fF
C8934 D_INPUT_5 OR2X1_LOC_752/a_8_216# 0.03fF
C8935 AND2X1_LOC_367/A OR2X1_LOC_106/A 0.05fF
C8936 OR2X1_LOC_604/A OR2X1_LOC_683/Y 0.02fF
C8937 AND2X1_LOC_366/A OR2X1_LOC_89/A 0.27fF
C8938 OR2X1_LOC_18/Y AND2X1_LOC_862/A 0.01fF
C8939 OR2X1_LOC_648/A OR2X1_LOC_602/a_8_216# 0.03fF
C8940 AND2X1_LOC_99/A AND2X1_LOC_124/a_8_24# 0.01fF
C8941 OR2X1_LOC_264/Y OR2X1_LOC_643/A 0.03fF
C8942 OR2X1_LOC_18/Y AND2X1_LOC_624/A 0.03fF
C8943 OR2X1_LOC_516/B OR2X1_LOC_52/B 0.03fF
C8944 AND2X1_LOC_181/Y INPUT_1 0.07fF
C8945 OR2X1_LOC_92/Y OR2X1_LOC_248/Y 0.08fF
C8946 D_INPUT_7 AND2X1_LOC_51/a_8_24# 0.02fF
C8947 AND2X1_LOC_344/a_36_24# OR2X1_LOC_44/Y 0.01fF
C8948 OR2X1_LOC_320/Y OR2X1_LOC_91/A 0.01fF
C8949 OR2X1_LOC_686/A AND2X1_LOC_425/Y 0.00fF
C8950 AND2X1_LOC_56/B OR2X1_LOC_730/a_8_216# -0.02fF
C8951 AND2X1_LOC_81/B OR2X1_LOC_507/B 0.01fF
C8952 OR2X1_LOC_319/B OR2X1_LOC_574/A 0.03fF
C8953 OR2X1_LOC_421/A AND2X1_LOC_639/A 0.12fF
C8954 AND2X1_LOC_318/Y AND2X1_LOC_786/Y 0.02fF
C8955 OR2X1_LOC_114/Y OR2X1_LOC_631/a_8_216# 0.13fF
C8956 OR2X1_LOC_379/Y AND2X1_LOC_56/B 0.03fF
C8957 OR2X1_LOC_662/A OR2X1_LOC_520/Y 0.75fF
C8958 OR2X1_LOC_431/Y OR2X1_LOC_56/A 0.02fF
C8959 OR2X1_LOC_179/Y OR2X1_LOC_485/A 0.01fF
C8960 OR2X1_LOC_249/Y OR2X1_LOC_579/B 0.02fF
C8961 AND2X1_LOC_3/Y OR2X1_LOC_721/Y 0.06fF
C8962 VDD OR2X1_LOC_22/A 0.27fF
C8963 OR2X1_LOC_92/Y AND2X1_LOC_294/a_36_24# 0.00fF
C8964 AND2X1_LOC_351/Y OR2X1_LOC_59/Y 0.07fF
C8965 OR2X1_LOC_790/a_8_216# OR2X1_LOC_375/A 0.02fF
C8966 OR2X1_LOC_650/a_8_216# OR2X1_LOC_650/Y 0.01fF
C8967 OR2X1_LOC_158/A OR2X1_LOC_409/B 0.03fF
C8968 AND2X1_LOC_474/A OR2X1_LOC_64/Y 0.04fF
C8969 VDD OR2X1_LOC_720/B 0.09fF
C8970 AND2X1_LOC_580/A OR2X1_LOC_680/A 0.03fF
C8971 AND2X1_LOC_216/Y AND2X1_LOC_656/Y 0.00fF
C8972 OR2X1_LOC_421/a_8_216# OR2X1_LOC_64/Y 0.02fF
C8973 OR2X1_LOC_756/B AND2X1_LOC_51/Y 0.87fF
C8974 AND2X1_LOC_70/Y AND2X1_LOC_667/a_8_24# 0.01fF
C8975 OR2X1_LOC_471/Y OR2X1_LOC_741/Y 0.02fF
C8976 OR2X1_LOC_181/B OR2X1_LOC_564/B 0.15fF
C8977 OR2X1_LOC_651/a_8_216# AND2X1_LOC_43/B 0.04fF
C8978 OR2X1_LOC_462/B OR2X1_LOC_642/a_8_216# 0.03fF
C8979 AND2X1_LOC_56/B OR2X1_LOC_194/Y 0.00fF
C8980 AND2X1_LOC_392/A AND2X1_LOC_864/a_8_24# 0.06fF
C8981 AND2X1_LOC_733/a_8_24# OR2X1_LOC_64/Y 0.05fF
C8982 OR2X1_LOC_7/A AND2X1_LOC_573/A 0.11fF
C8983 AND2X1_LOC_42/B OR2X1_LOC_560/a_8_216# 0.01fF
C8984 OR2X1_LOC_777/B OR2X1_LOC_723/B 0.03fF
C8985 OR2X1_LOC_448/Y OR2X1_LOC_453/A 0.06fF
C8986 OR2X1_LOC_574/A OR2X1_LOC_805/A 0.10fF
C8987 AND2X1_LOC_863/Y OR2X1_LOC_56/A 0.08fF
C8988 OR2X1_LOC_100/Y OR2X1_LOC_121/B 0.16fF
C8989 OR2X1_LOC_375/A AND2X1_LOC_3/Y 0.31fF
C8990 OR2X1_LOC_68/B OR2X1_LOC_227/A 0.04fF
C8991 OR2X1_LOC_479/Y OR2X1_LOC_739/A 0.03fF
C8992 OR2X1_LOC_375/A OR2X1_LOC_647/B 0.03fF
C8993 OR2X1_LOC_445/a_8_216# OR2X1_LOC_553/A 0.04fF
C8994 OR2X1_LOC_125/a_36_216# D_INPUT_3 0.00fF
C8995 OR2X1_LOC_24/a_8_216# OR2X1_LOC_44/Y 0.06fF
C8996 OR2X1_LOC_47/Y AND2X1_LOC_614/a_8_24# 0.02fF
C8997 OR2X1_LOC_643/A OR2X1_LOC_124/Y 0.03fF
C8998 OR2X1_LOC_18/Y AND2X1_LOC_853/a_8_24# 0.01fF
C8999 OR2X1_LOC_544/B OR2X1_LOC_180/B 0.01fF
C9000 AND2X1_LOC_394/a_8_24# AND2X1_LOC_42/B 0.01fF
C9001 OR2X1_LOC_259/A OR2X1_LOC_348/B 0.11fF
C9002 AND2X1_LOC_474/A OR2X1_LOC_417/A 0.03fF
C9003 OR2X1_LOC_18/Y AND2X1_LOC_650/a_36_24# 0.01fF
C9004 OR2X1_LOC_598/Y OR2X1_LOC_214/B 0.08fF
C9005 AND2X1_LOC_557/Y AND2X1_LOC_489/Y 0.01fF
C9006 AND2X1_LOC_59/Y OR2X1_LOC_476/Y 0.01fF
C9007 AND2X1_LOC_369/a_8_24# OR2X1_LOC_787/Y 0.04fF
C9008 OR2X1_LOC_428/A AND2X1_LOC_563/Y 0.02fF
C9009 OR2X1_LOC_36/Y AND2X1_LOC_459/a_8_24# 0.02fF
C9010 AND2X1_LOC_12/Y OR2X1_LOC_202/a_8_216# 0.01fF
C9011 OR2X1_LOC_113/Y AND2X1_LOC_106/a_8_24# 0.23fF
C9012 OR2X1_LOC_64/Y AND2X1_LOC_593/Y 0.01fF
C9013 OR2X1_LOC_506/A AND2X1_LOC_491/a_8_24# 0.17fF
C9014 AND2X1_LOC_523/a_8_24# AND2X1_LOC_115/a_8_24# 0.23fF
C9015 AND2X1_LOC_367/A AND2X1_LOC_227/Y 0.05fF
C9016 OR2X1_LOC_757/A GATE_662 0.15fF
C9017 OR2X1_LOC_600/A AND2X1_LOC_624/B 0.28fF
C9018 OR2X1_LOC_684/Y AND2X1_LOC_452/Y 0.10fF
C9019 OR2X1_LOC_74/A AND2X1_LOC_264/a_8_24# 0.02fF
C9020 OR2X1_LOC_277/a_36_216# OR2X1_LOC_39/A 0.00fF
C9021 OR2X1_LOC_595/A AND2X1_LOC_563/Y 0.11fF
C9022 OR2X1_LOC_3/Y OR2X1_LOC_588/Y 0.03fF
C9023 OR2X1_LOC_780/A AND2X1_LOC_424/a_8_24# 0.20fF
C9024 OR2X1_LOC_52/a_8_216# OR2X1_LOC_6/A 0.01fF
C9025 AND2X1_LOC_677/a_8_24# OR2X1_LOC_161/A 0.02fF
C9026 OR2X1_LOC_479/Y OR2X1_LOC_269/B 0.07fF
C9027 AND2X1_LOC_580/B OR2X1_LOC_617/Y 0.05fF
C9028 OR2X1_LOC_748/A OR2X1_LOC_481/A 0.06fF
C9029 OR2X1_LOC_64/Y OR2X1_LOC_85/A 0.11fF
C9030 OR2X1_LOC_185/A OR2X1_LOC_68/Y 0.01fF
C9031 OR2X1_LOC_561/Y D_INPUT_1 0.00fF
C9032 OR2X1_LOC_78/Y D_INPUT_1 0.03fF
C9033 OR2X1_LOC_835/B OR2X1_LOC_19/B 0.10fF
C9034 OR2X1_LOC_274/a_8_216# D_INPUT_1 0.04fF
C9035 OR2X1_LOC_78/B OR2X1_LOC_194/a_8_216# 0.03fF
C9036 OR2X1_LOC_404/Y OR2X1_LOC_720/a_8_216# 0.01fF
C9037 AND2X1_LOC_95/Y AND2X1_LOC_108/a_8_24# 0.01fF
C9038 OR2X1_LOC_709/A AND2X1_LOC_419/a_8_24# 0.02fF
C9039 AND2X1_LOC_675/A OR2X1_LOC_531/a_8_216# 0.18fF
C9040 OR2X1_LOC_472/B AND2X1_LOC_413/a_8_24# 0.03fF
C9041 OR2X1_LOC_335/A AND2X1_LOC_591/a_36_24# 0.00fF
C9042 OR2X1_LOC_557/A AND2X1_LOC_815/a_8_24# 0.06fF
C9043 OR2X1_LOC_272/Y AND2X1_LOC_78/a_8_24# 0.16fF
C9044 OR2X1_LOC_256/a_8_216# OR2X1_LOC_95/Y 0.03fF
C9045 OR2X1_LOC_7/A OR2X1_LOC_27/Y 0.15fF
C9046 OR2X1_LOC_824/a_8_216# OR2X1_LOC_291/A 0.01fF
C9047 OR2X1_LOC_185/A AND2X1_LOC_47/Y 0.17fF
C9048 AND2X1_LOC_56/B OR2X1_LOC_444/a_8_216# 0.06fF
C9049 AND2X1_LOC_432/a_8_24# AND2X1_LOC_18/Y 0.02fF
C9050 AND2X1_LOC_642/a_8_24# AND2X1_LOC_476/A 0.01fF
C9051 OR2X1_LOC_529/Y AND2X1_LOC_523/Y 0.68fF
C9052 OR2X1_LOC_487/a_36_216# OR2X1_LOC_488/Y 0.00fF
C9053 AND2X1_LOC_841/B AND2X1_LOC_648/B 0.00fF
C9054 OR2X1_LOC_97/A OR2X1_LOC_374/a_8_216# 0.02fF
C9055 AND2X1_LOC_18/Y OR2X1_LOC_578/B 0.27fF
C9056 AND2X1_LOC_40/Y OR2X1_LOC_214/B 0.03fF
C9057 AND2X1_LOC_566/B AND2X1_LOC_212/a_8_24# 0.00fF
C9058 OR2X1_LOC_756/B OR2X1_LOC_551/B 0.29fF
C9059 OR2X1_LOC_643/A OR2X1_LOC_113/A 0.00fF
C9060 AND2X1_LOC_99/A OR2X1_LOC_47/Y 0.02fF
C9061 OR2X1_LOC_291/Y OR2X1_LOC_609/a_36_216# 0.02fF
C9062 OR2X1_LOC_473/Y OR2X1_LOC_475/Y 0.02fF
C9063 OR2X1_LOC_269/a_8_216# OR2X1_LOC_269/Y -0.00fF
C9064 OR2X1_LOC_691/Y AND2X1_LOC_36/Y 0.01fF
C9065 INPUT_1 OR2X1_LOC_585/A 0.03fF
C9066 OR2X1_LOC_532/B OR2X1_LOC_449/B 0.03fF
C9067 OR2X1_LOC_6/B OR2X1_LOC_399/Y 0.02fF
C9068 OR2X1_LOC_70/Y AND2X1_LOC_351/Y 0.15fF
C9069 OR2X1_LOC_74/A OR2X1_LOC_46/A 0.01fF
C9070 AND2X1_LOC_357/B OR2X1_LOC_437/A 0.02fF
C9071 AND2X1_LOC_726/Y AND2X1_LOC_727/Y 0.11fF
C9072 AND2X1_LOC_722/A AND2X1_LOC_222/Y 0.00fF
C9073 AND2X1_LOC_624/A AND2X1_LOC_620/Y 0.23fF
C9074 AND2X1_LOC_142/a_36_24# OR2X1_LOC_705/B 0.01fF
C9075 AND2X1_LOC_851/B OR2X1_LOC_36/Y 0.07fF
C9076 OR2X1_LOC_619/Y OR2X1_LOC_67/Y 0.07fF
C9077 AND2X1_LOC_377/Y OR2X1_LOC_39/a_8_216# 0.03fF
C9078 VDD AND2X1_LOC_742/A 0.21fF
C9079 AND2X1_LOC_514/Y AND2X1_LOC_326/A 0.01fF
C9080 OR2X1_LOC_494/Y OR2X1_LOC_437/A 0.01fF
C9081 OR2X1_LOC_670/a_36_216# D_INPUT_3 0.00fF
C9082 AND2X1_LOC_363/Y OR2X1_LOC_437/A 0.02fF
C9083 AND2X1_LOC_465/A AND2X1_LOC_242/B 0.06fF
C9084 OR2X1_LOC_679/A OR2X1_LOC_74/A 0.03fF
C9085 OR2X1_LOC_840/A OR2X1_LOC_779/B 0.01fF
C9086 OR2X1_LOC_420/a_8_216# OR2X1_LOC_95/Y 0.03fF
C9087 OR2X1_LOC_783/A OR2X1_LOC_155/A 0.02fF
C9088 AND2X1_LOC_260/a_36_24# OR2X1_LOC_54/Y 0.01fF
C9089 OR2X1_LOC_261/A OR2X1_LOC_46/A 0.00fF
C9090 OR2X1_LOC_22/Y OR2X1_LOC_829/Y 0.01fF
C9091 AND2X1_LOC_456/Y AND2X1_LOC_227/Y 0.02fF
C9092 OR2X1_LOC_828/Y AND2X1_LOC_829/a_8_24# 0.00fF
C9093 OR2X1_LOC_19/B OR2X1_LOC_278/A 0.07fF
C9094 OR2X1_LOC_185/A OR2X1_LOC_598/A 0.10fF
C9095 AND2X1_LOC_729/Y OR2X1_LOC_419/a_36_216# 0.01fF
C9096 OR2X1_LOC_70/Y OR2X1_LOC_167/Y 0.16fF
C9097 OR2X1_LOC_193/A D_INPUT_0 0.26fF
C9098 OR2X1_LOC_287/B OR2X1_LOC_62/A 0.02fF
C9099 AND2X1_LOC_548/Y OR2X1_LOC_437/A 0.01fF
C9100 AND2X1_LOC_721/A OR2X1_LOC_6/A 0.16fF
C9101 OR2X1_LOC_619/Y OR2X1_LOC_163/Y 0.01fF
C9102 OR2X1_LOC_620/Y AND2X1_LOC_31/Y 0.02fF
C9103 OR2X1_LOC_696/A AND2X1_LOC_212/A 0.03fF
C9104 OR2X1_LOC_196/Y AND2X1_LOC_22/Y 0.35fF
C9105 AND2X1_LOC_721/Y AND2X1_LOC_734/a_8_24# 0.09fF
C9106 AND2X1_LOC_539/Y AND2X1_LOC_809/a_8_24# 0.01fF
C9107 AND2X1_LOC_7/B AND2X1_LOC_627/a_8_24# 0.10fF
C9108 AND2X1_LOC_303/a_8_24# OR2X1_LOC_437/A 0.03fF
C9109 OR2X1_LOC_440/a_8_216# OR2X1_LOC_180/B 0.01fF
C9110 OR2X1_LOC_121/B OR2X1_LOC_532/B 0.30fF
C9111 OR2X1_LOC_64/Y OR2X1_LOC_226/Y 0.01fF
C9112 AND2X1_LOC_861/B OR2X1_LOC_13/B 0.01fF
C9113 OR2X1_LOC_36/Y OR2X1_LOC_595/Y 0.84fF
C9114 OR2X1_LOC_326/a_8_216# OR2X1_LOC_532/Y 0.03fF
C9115 OR2X1_LOC_51/B OR2X1_LOC_47/a_8_216# 0.00fF
C9116 AND2X1_LOC_634/Y INPUT_1 0.01fF
C9117 OR2X1_LOC_302/B OR2X1_LOC_469/B 0.03fF
C9118 OR2X1_LOC_49/A OR2X1_LOC_428/A 0.22fF
C9119 AND2X1_LOC_91/B OR2X1_LOC_673/a_36_216# 0.00fF
C9120 OR2X1_LOC_831/A AND2X1_LOC_273/a_36_24# 0.01fF
C9121 OR2X1_LOC_45/B AND2X1_LOC_249/a_8_24# 0.11fF
C9122 OR2X1_LOC_78/A OR2X1_LOC_308/Y 0.07fF
C9123 OR2X1_LOC_405/A AND2X1_LOC_406/a_8_24# 0.26fF
C9124 OR2X1_LOC_154/A AND2X1_LOC_31/Y 0.58fF
C9125 OR2X1_LOC_154/A OR2X1_LOC_715/a_8_216# 0.03fF
C9126 OR2X1_LOC_813/Y OR2X1_LOC_74/A 0.15fF
C9127 OR2X1_LOC_3/Y OR2X1_LOC_86/A 0.00fF
C9128 OR2X1_LOC_170/A OR2X1_LOC_568/A 0.05fF
C9129 OR2X1_LOC_333/B OR2X1_LOC_351/a_8_216# 0.48fF
C9130 AND2X1_LOC_171/a_8_24# OR2X1_LOC_358/A 0.01fF
C9131 OR2X1_LOC_315/a_36_216# AND2X1_LOC_786/Y 0.01fF
C9132 AND2X1_LOC_339/B OR2X1_LOC_16/A 0.05fF
C9133 OR2X1_LOC_732/B OR2X1_LOC_732/A 0.13fF
C9134 AND2X1_LOC_70/Y OR2X1_LOC_115/B 0.00fF
C9135 OR2X1_LOC_417/A OR2X1_LOC_226/Y 0.05fF
C9136 AND2X1_LOC_712/Y OR2X1_LOC_428/A 0.01fF
C9137 OR2X1_LOC_182/B OR2X1_LOC_357/B 0.01fF
C9138 AND2X1_LOC_663/B AND2X1_LOC_792/Y 0.01fF
C9139 OR2X1_LOC_111/Y AND2X1_LOC_831/Y 0.09fF
C9140 OR2X1_LOC_269/B OR2X1_LOC_68/B 0.03fF
C9141 AND2X1_LOC_95/Y OR2X1_LOC_544/B 0.07fF
C9142 AND2X1_LOC_22/Y AND2X1_LOC_95/a_8_24# 0.02fF
C9143 OR2X1_LOC_492/a_36_216# OR2X1_LOC_492/Y 0.00fF
C9144 OR2X1_LOC_486/B OR2X1_LOC_705/B 0.14fF
C9145 VDD AND2X1_LOC_769/Y 0.25fF
C9146 OR2X1_LOC_696/A OR2X1_LOC_251/a_8_216# 0.05fF
C9147 AND2X1_LOC_621/a_8_24# AND2X1_LOC_620/Y 0.00fF
C9148 OR2X1_LOC_599/A OR2X1_LOC_423/Y 0.01fF
C9149 AND2X1_LOC_183/a_36_24# OR2X1_LOC_190/A 0.01fF
C9150 AND2X1_LOC_474/A OR2X1_LOC_89/a_36_216# 0.00fF
C9151 AND2X1_LOC_64/Y AND2X1_LOC_41/A 1.61fF
C9152 OR2X1_LOC_492/Y OR2X1_LOC_482/Y 0.19fF
C9153 OR2X1_LOC_121/Y OR2X1_LOC_631/A 0.02fF
C9154 OR2X1_LOC_154/a_8_216# OR2X1_LOC_803/A 0.01fF
C9155 OR2X1_LOC_535/A AND2X1_LOC_110/Y 0.01fF
C9156 OR2X1_LOC_176/a_8_216# OR2X1_LOC_91/A 0.01fF
C9157 AND2X1_LOC_364/Y OR2X1_LOC_321/a_36_216# 0.00fF
C9158 OR2X1_LOC_778/A AND2X1_LOC_31/Y 0.00fF
C9159 OR2X1_LOC_51/Y OR2X1_LOC_766/a_8_216# 0.01fF
C9160 OR2X1_LOC_151/A OR2X1_LOC_140/A 0.01fF
C9161 OR2X1_LOC_508/A AND2X1_LOC_64/Y 0.13fF
C9162 AND2X1_LOC_647/Y OR2X1_LOC_46/A 0.06fF
C9163 OR2X1_LOC_118/a_8_216# OR2X1_LOC_744/A 0.01fF
C9164 INPUT_5 AND2X1_LOC_587/a_8_24# 0.01fF
C9165 OR2X1_LOC_215/A OR2X1_LOC_68/B 0.08fF
C9166 OR2X1_LOC_506/Y OR2X1_LOC_242/a_8_216# 0.41fF
C9167 AND2X1_LOC_645/A OR2X1_LOC_13/B 0.02fF
C9168 OR2X1_LOC_45/B AND2X1_LOC_734/Y 0.15fF
C9169 OR2X1_LOC_40/Y AND2X1_LOC_806/a_8_24# 0.04fF
C9170 OR2X1_LOC_696/A OR2X1_LOC_127/a_36_216# 0.00fF
C9171 AND2X1_LOC_110/Y AND2X1_LOC_323/a_8_24# 0.09fF
C9172 OR2X1_LOC_510/Y OR2X1_LOC_508/Y 0.01fF
C9173 OR2X1_LOC_528/Y OR2X1_LOC_627/Y 0.03fF
C9174 AND2X1_LOC_788/a_8_24# OR2X1_LOC_59/Y 0.01fF
C9175 AND2X1_LOC_58/a_8_24# AND2X1_LOC_7/B 0.01fF
C9176 OR2X1_LOC_748/A AND2X1_LOC_789/Y 0.28fF
C9177 AND2X1_LOC_360/a_36_24# OR2X1_LOC_494/A 0.00fF
C9178 AND2X1_LOC_357/B AND2X1_LOC_715/A 0.10fF
C9179 AND2X1_LOC_91/B AND2X1_LOC_384/a_36_24# 0.01fF
C9180 OR2X1_LOC_528/Y AND2X1_LOC_500/Y 0.03fF
C9181 OR2X1_LOC_124/a_36_216# OR2X1_LOC_641/A 0.01fF
C9182 OR2X1_LOC_620/B OR2X1_LOC_550/B 0.04fF
C9183 OR2X1_LOC_244/a_36_216# OR2X1_LOC_576/A 0.00fF
C9184 AND2X1_LOC_810/a_8_24# OR2X1_LOC_47/Y 0.04fF
C9185 OR2X1_LOC_450/a_8_216# OR2X1_LOC_450/Y -0.00fF
C9186 AND2X1_LOC_362/B OR2X1_LOC_59/Y 0.00fF
C9187 AND2X1_LOC_476/Y OR2X1_LOC_59/Y 0.07fF
C9188 OR2X1_LOC_161/A OR2X1_LOC_140/B 0.46fF
C9189 OR2X1_LOC_359/A OR2X1_LOC_362/A 0.02fF
C9190 OR2X1_LOC_348/Y OR2X1_LOC_66/A 0.17fF
C9191 OR2X1_LOC_633/a_36_216# OR2X1_LOC_549/A 0.00fF
C9192 OR2X1_LOC_641/A AND2X1_LOC_92/Y 0.00fF
C9193 AND2X1_LOC_16/a_8_24# AND2X1_LOC_7/B 0.01fF
C9194 OR2X1_LOC_683/a_8_216# OR2X1_LOC_12/Y 0.01fF
C9195 OR2X1_LOC_422/Y OR2X1_LOC_428/A 0.01fF
C9196 AND2X1_LOC_353/a_8_24# OR2X1_LOC_91/A 0.01fF
C9197 AND2X1_LOC_787/A OR2X1_LOC_427/A 0.00fF
C9198 OR2X1_LOC_709/A OR2X1_LOC_840/A 0.10fF
C9199 OR2X1_LOC_124/a_8_216# AND2X1_LOC_70/Y 0.01fF
C9200 OR2X1_LOC_696/A OR2X1_LOC_824/Y 0.16fF
C9201 OR2X1_LOC_355/B OR2X1_LOC_703/Y 0.04fF
C9202 OR2X1_LOC_377/A AND2X1_LOC_7/B 0.12fF
C9203 OR2X1_LOC_114/B OR2X1_LOC_632/Y 0.01fF
C9204 AND2X1_LOC_866/A AND2X1_LOC_222/Y 0.03fF
C9205 OR2X1_LOC_703/B OR2X1_LOC_703/a_8_216# 0.07fF
C9206 OR2X1_LOC_160/A OR2X1_LOC_227/B 0.01fF
C9207 OR2X1_LOC_828/B OR2X1_LOC_828/Y 1.00fF
C9208 OR2X1_LOC_696/A OR2X1_LOC_591/a_8_216# 0.03fF
C9209 OR2X1_LOC_427/A AND2X1_LOC_457/a_36_24# 0.00fF
C9210 AND2X1_LOC_59/Y OR2X1_LOC_563/A 0.02fF
C9211 AND2X1_LOC_586/a_8_24# OR2X1_LOC_691/Y 0.01fF
C9212 OR2X1_LOC_48/B AND2X1_LOC_774/A 0.02fF
C9213 OR2X1_LOC_433/Y OR2X1_LOC_428/A 0.03fF
C9214 OR2X1_LOC_651/A OR2X1_LOC_228/Y 0.03fF
C9215 AND2X1_LOC_824/B AND2X1_LOC_7/B 0.03fF
C9216 OR2X1_LOC_278/A AND2X1_LOC_608/a_8_24# 0.01fF
C9217 OR2X1_LOC_97/A OR2X1_LOC_640/a_8_216# 0.04fF
C9218 OR2X1_LOC_134/a_36_216# AND2X1_LOC_560/B 0.01fF
C9219 AND2X1_LOC_64/Y OR2X1_LOC_631/B 0.06fF
C9220 AND2X1_LOC_738/B OR2X1_LOC_744/A 0.07fF
C9221 AND2X1_LOC_550/A AND2X1_LOC_727/B 0.03fF
C9222 INPUT_0 OR2X1_LOC_51/Y 0.03fF
C9223 OR2X1_LOC_18/Y AND2X1_LOC_774/A 0.00fF
C9224 OR2X1_LOC_744/A OR2X1_LOC_56/A 0.17fF
C9225 OR2X1_LOC_6/B OR2X1_LOC_833/a_8_216# 0.07fF
C9226 AND2X1_LOC_174/a_8_24# OR2X1_LOC_12/Y 0.01fF
C9227 AND2X1_LOC_91/B OR2X1_LOC_643/A 0.34fF
C9228 OR2X1_LOC_118/Y OR2X1_LOC_12/Y 0.00fF
C9229 OR2X1_LOC_833/B AND2X1_LOC_256/a_36_24# 0.01fF
C9230 OR2X1_LOC_653/Y OR2X1_LOC_151/A 0.01fF
C9231 AND2X1_LOC_684/a_8_24# AND2X1_LOC_31/Y 0.01fF
C9232 AND2X1_LOC_341/a_8_24# AND2X1_LOC_228/Y 0.03fF
C9233 AND2X1_LOC_91/B OR2X1_LOC_778/Y 0.14fF
C9234 OR2X1_LOC_203/Y AND2X1_LOC_7/B 0.09fF
C9235 AND2X1_LOC_40/Y OR2X1_LOC_325/B 0.03fF
C9236 AND2X1_LOC_477/A OR2X1_LOC_13/B 0.07fF
C9237 INPUT_0 OR2X1_LOC_78/B 0.08fF
C9238 AND2X1_LOC_574/Y AND2X1_LOC_474/Y 0.05fF
C9239 OR2X1_LOC_62/B OR2X1_LOC_141/a_36_216# 0.00fF
C9240 OR2X1_LOC_441/Y AND2X1_LOC_657/Y 0.60fF
C9241 OR2X1_LOC_621/A OR2X1_LOC_847/A 0.01fF
C9242 AND2X1_LOC_486/Y OR2X1_LOC_600/A 0.03fF
C9243 AND2X1_LOC_70/Y OR2X1_LOC_840/A 0.03fF
C9244 AND2X1_LOC_533/a_36_24# OR2X1_LOC_356/A 0.06fF
C9245 OR2X1_LOC_232/Y AND2X1_LOC_240/a_8_24# 0.23fF
C9246 AND2X1_LOC_555/a_8_24# AND2X1_LOC_847/Y 0.02fF
C9247 OR2X1_LOC_441/Y AND2X1_LOC_469/B 0.03fF
C9248 OR2X1_LOC_673/Y OR2X1_LOC_161/B 0.00fF
C9249 OR2X1_LOC_95/Y OR2X1_LOC_385/a_8_216# 0.39fF
C9250 OR2X1_LOC_744/A AND2X1_LOC_638/Y 0.36fF
C9251 OR2X1_LOC_624/Y OR2X1_LOC_659/A 0.14fF
C9252 OR2X1_LOC_47/Y OR2X1_LOC_152/a_36_216# 0.03fF
C9253 OR2X1_LOC_625/Y AND2X1_LOC_614/a_8_24# 0.06fF
C9254 OR2X1_LOC_440/A OR2X1_LOC_303/B 0.03fF
C9255 AND2X1_LOC_717/Y OR2X1_LOC_51/Y 4.61fF
C9256 AND2X1_LOC_448/Y AND2X1_LOC_448/a_8_24# 0.05fF
C9257 OR2X1_LOC_426/B OR2X1_LOC_586/Y 0.91fF
C9258 OR2X1_LOC_164/Y AND2X1_LOC_471/Y 0.16fF
C9259 AND2X1_LOC_773/Y AND2X1_LOC_264/a_36_24# 0.01fF
C9260 OR2X1_LOC_377/A OR2X1_LOC_621/a_8_216# 0.05fF
C9261 AND2X1_LOC_440/a_36_24# OR2X1_LOC_437/A 0.01fF
C9262 AND2X1_LOC_12/Y OR2X1_LOC_631/A 0.01fF
C9263 AND2X1_LOC_705/Y OR2X1_LOC_43/A 0.06fF
C9264 OR2X1_LOC_40/Y OR2X1_LOC_32/B 0.20fF
C9265 AND2X1_LOC_51/Y OR2X1_LOC_140/B 0.03fF
C9266 OR2X1_LOC_43/A AND2X1_LOC_809/a_36_24# 0.00fF
C9267 AND2X1_LOC_391/a_36_24# OR2X1_LOC_91/A 0.00fF
C9268 AND2X1_LOC_259/Y OR2X1_LOC_428/A 0.02fF
C9269 OR2X1_LOC_404/Y OR2X1_LOC_115/B 0.02fF
C9270 AND2X1_LOC_733/Y OR2X1_LOC_441/Y 0.00fF
C9271 VDD OR2X1_LOC_260/Y 0.06fF
C9272 AND2X1_LOC_736/Y AND2X1_LOC_735/Y 0.00fF
C9273 AND2X1_LOC_810/Y OR2X1_LOC_142/a_8_216# 0.07fF
C9274 AND2X1_LOC_775/a_8_24# AND2X1_LOC_476/Y 0.03fF
C9275 OR2X1_LOC_696/A AND2X1_LOC_727/A 0.03fF
C9276 OR2X1_LOC_512/A AND2X1_LOC_41/A 0.04fF
C9277 AND2X1_LOC_741/Y AND2X1_LOC_221/a_8_24# 0.14fF
C9278 OR2X1_LOC_6/A OR2X1_LOC_57/a_8_216# 0.07fF
C9279 OR2X1_LOC_160/B OR2X1_LOC_448/Y 0.11fF
C9280 AND2X1_LOC_40/Y AND2X1_LOC_189/a_8_24# 0.17fF
C9281 OR2X1_LOC_48/B AND2X1_LOC_434/a_8_24# 0.01fF
C9282 OR2X1_LOC_158/A OR2X1_LOC_497/Y 0.06fF
C9283 OR2X1_LOC_385/Y AND2X1_LOC_774/A 0.10fF
C9284 OR2X1_LOC_296/Y AND2X1_LOC_627/a_8_24# 0.01fF
C9285 OR2X1_LOC_17/Y OR2X1_LOC_18/a_8_216# 0.03fF
C9286 OR2X1_LOC_709/A OR2X1_LOC_789/a_8_216# 0.01fF
C9287 OR2X1_LOC_605/A AND2X1_LOC_604/a_8_24# 0.10fF
C9288 OR2X1_LOC_744/A AND2X1_LOC_850/Y 0.07fF
C9289 VDD OR2X1_LOC_613/a_8_216# 0.21fF
C9290 OR2X1_LOC_510/Y OR2X1_LOC_66/A 0.02fF
C9291 AND2X1_LOC_443/a_8_24# OR2X1_LOC_52/B 0.01fF
C9292 VDD OR2X1_LOC_148/B -0.00fF
C9293 AND2X1_LOC_40/Y OR2X1_LOC_285/a_8_216# 0.01fF
C9294 INPUT_0 AND2X1_LOC_642/a_8_24# 0.01fF
C9295 OR2X1_LOC_751/Y AND2X1_LOC_789/a_8_24# 0.01fF
C9296 OR2X1_LOC_820/B OR2X1_LOC_382/a_36_216# 0.00fF
C9297 AND2X1_LOC_94/a_8_24# INPUT_0 0.04fF
C9298 AND2X1_LOC_500/a_8_24# AND2X1_LOC_500/B 0.00fF
C9299 AND2X1_LOC_64/Y OR2X1_LOC_403/a_8_216# 0.06fF
C9300 OR2X1_LOC_51/Y OR2X1_LOC_11/Y 0.07fF
C9301 AND2X1_LOC_3/Y OR2X1_LOC_549/A 0.12fF
C9302 OR2X1_LOC_471/a_8_216# OR2X1_LOC_471/B 0.39fF
C9303 AND2X1_LOC_51/Y OR2X1_LOC_355/A 0.04fF
C9304 AND2X1_LOC_94/Y AND2X1_LOC_43/B 0.09fF
C9305 AND2X1_LOC_391/Y OR2X1_LOC_127/Y 0.06fF
C9306 AND2X1_LOC_12/Y OR2X1_LOC_632/Y 1.49fF
C9307 AND2X1_LOC_663/A OR2X1_LOC_39/A 0.06fF
C9308 OR2X1_LOC_306/Y AND2X1_LOC_434/Y 0.03fF
C9309 AND2X1_LOC_715/Y AND2X1_LOC_727/A 0.00fF
C9310 OR2X1_LOC_494/Y AND2X1_LOC_348/Y 0.01fF
C9311 OR2X1_LOC_127/Y OR2X1_LOC_91/A 0.10fF
C9312 OR2X1_LOC_690/a_8_216# VDD 0.21fF
C9313 OR2X1_LOC_421/A OR2X1_LOC_52/B 0.04fF
C9314 OR2X1_LOC_822/a_36_216# OR2X1_LOC_753/A 0.00fF
C9315 VDD AND2X1_LOC_818/a_8_24# 0.00fF
C9316 OR2X1_LOC_850/B OR2X1_LOC_811/A 0.03fF
C9317 AND2X1_LOC_810/A AND2X1_LOC_798/Y 0.01fF
C9318 AND2X1_LOC_363/Y AND2X1_LOC_348/Y 1.02fF
C9319 AND2X1_LOC_840/a_8_24# OR2X1_LOC_495/Y 0.01fF
C9320 OR2X1_LOC_91/Y OR2X1_LOC_107/a_8_216# 0.05fF
C9321 AND2X1_LOC_191/Y AND2X1_LOC_476/Y 1.50fF
C9322 AND2X1_LOC_576/Y AND2X1_LOC_658/A 0.07fF
C9323 OR2X1_LOC_185/A AND2X1_LOC_529/a_36_24# 0.01fF
C9324 INPUT_0 OR2X1_LOC_375/A 0.12fF
C9325 OR2X1_LOC_319/B OR2X1_LOC_319/a_8_216# 0.02fF
C9326 AND2X1_LOC_738/B AND2X1_LOC_840/B 0.03fF
C9327 OR2X1_LOC_696/A OR2X1_LOC_95/Y 1.22fF
C9328 AND2X1_LOC_788/a_8_24# OR2X1_LOC_70/Y 0.01fF
C9329 OR2X1_LOC_494/Y OR2X1_LOC_753/A 0.03fF
C9330 AND2X1_LOC_840/B OR2X1_LOC_56/A 0.05fF
C9331 OR2X1_LOC_757/A AND2X1_LOC_580/A 0.03fF
C9332 AND2X1_LOC_147/a_8_24# OR2X1_LOC_427/A 0.03fF
C9333 AND2X1_LOC_363/Y OR2X1_LOC_753/A 0.02fF
C9334 OR2X1_LOC_696/A OR2X1_LOC_368/A 0.01fF
C9335 AND2X1_LOC_555/Y OR2X1_LOC_417/A 0.01fF
C9336 AND2X1_LOC_711/Y AND2X1_LOC_476/Y 0.07fF
C9337 OR2X1_LOC_810/A OR2X1_LOC_66/A 0.18fF
C9338 OR2X1_LOC_85/A OR2X1_LOC_232/Y 0.02fF
C9339 OR2X1_LOC_70/Y AND2X1_LOC_476/Y 0.14fF
C9340 OR2X1_LOC_318/Y OR2X1_LOC_319/a_8_216# 0.02fF
C9341 AND2X1_LOC_563/A AND2X1_LOC_489/Y 0.02fF
C9342 AND2X1_LOC_756/a_8_24# AND2X1_LOC_580/B 0.01fF
C9343 OR2X1_LOC_251/Y AND2X1_LOC_286/a_8_24# 0.01fF
C9344 VDD OR2X1_LOC_793/B -0.00fF
C9345 AND2X1_LOC_364/Y OR2X1_LOC_36/Y 0.06fF
C9346 AND2X1_LOC_50/Y AND2X1_LOC_43/B 0.02fF
C9347 OR2X1_LOC_290/Y OR2X1_LOC_316/Y 0.02fF
C9348 OR2X1_LOC_447/Y OR2X1_LOC_779/A 0.03fF
C9349 AND2X1_LOC_425/Y OR2X1_LOC_161/B 0.01fF
C9350 OR2X1_LOC_136/Y OR2X1_LOC_417/A 0.00fF
C9351 OR2X1_LOC_653/A OR2X1_LOC_435/B 0.01fF
C9352 AND2X1_LOC_810/A OR2X1_LOC_46/A 0.02fF
C9353 OR2X1_LOC_158/A AND2X1_LOC_844/a_8_24# 0.02fF
C9354 OR2X1_LOC_279/Y AND2X1_LOC_244/a_8_24# 0.03fF
C9355 AND2X1_LOC_589/a_8_24# OR2X1_LOC_66/A 0.01fF
C9356 AND2X1_LOC_658/B OR2X1_LOC_680/Y 0.03fF
C9357 OR2X1_LOC_254/B AND2X1_LOC_253/a_36_24# 0.00fF
C9358 AND2X1_LOC_715/Y OR2X1_LOC_95/Y 0.00fF
C9359 OR2X1_LOC_593/A OR2X1_LOC_78/A 0.01fF
C9360 OR2X1_LOC_46/A OR2X1_LOC_9/a_36_216# 0.00fF
C9361 AND2X1_LOC_40/Y OR2X1_LOC_652/a_36_216# 0.00fF
C9362 OR2X1_LOC_358/a_8_216# OR2X1_LOC_502/A 0.01fF
C9363 AND2X1_LOC_191/B OR2X1_LOC_529/Y 0.02fF
C9364 AND2X1_LOC_350/B D_INPUT_0 0.01fF
C9365 AND2X1_LOC_768/a_8_24# AND2X1_LOC_276/Y 0.11fF
C9366 OR2X1_LOC_624/A OR2X1_LOC_668/a_36_216# 0.12fF
C9367 OR2X1_LOC_621/B AND2X1_LOC_670/a_36_24# 0.01fF
C9368 AND2X1_LOC_496/a_36_24# AND2X1_LOC_18/Y 0.01fF
C9369 AND2X1_LOC_364/A AND2X1_LOC_655/A 0.10fF
C9370 OR2X1_LOC_185/A OR2X1_LOC_506/A 0.02fF
C9371 OR2X1_LOC_834/a_8_216# OR2X1_LOC_269/B 0.01fF
C9372 AND2X1_LOC_198/a_36_24# OR2X1_LOC_6/A 0.00fF
C9373 OR2X1_LOC_282/a_8_216# OR2X1_LOC_56/A 0.05fF
C9374 OR2X1_LOC_290/a_8_216# OR2X1_LOC_26/Y 0.07fF
C9375 OR2X1_LOC_791/B OR2X1_LOC_260/a_8_216# 0.01fF
C9376 AND2X1_LOC_848/Y OR2X1_LOC_278/Y 0.03fF
C9377 OR2X1_LOC_185/A OR2X1_LOC_341/Y 0.01fF
C9378 OR2X1_LOC_426/B OR2X1_LOC_304/Y 0.45fF
C9379 OR2X1_LOC_690/a_8_216# OR2X1_LOC_689/A -0.00fF
C9380 OR2X1_LOC_517/A OR2X1_LOC_585/A 0.75fF
C9381 OR2X1_LOC_8/Y OR2X1_LOC_825/Y 0.03fF
C9382 AND2X1_LOC_332/a_8_24# OR2X1_LOC_417/A 0.03fF
C9383 OR2X1_LOC_857/a_8_216# OR2X1_LOC_66/A 0.01fF
C9384 VDD AND2X1_LOC_430/a_8_24# 0.00fF
C9385 OR2X1_LOC_377/A OR2X1_LOC_805/A 0.83fF
C9386 OR2X1_LOC_51/Y OR2X1_LOC_64/Y 2.25fF
C9387 OR2X1_LOC_185/Y OR2X1_LOC_560/a_8_216# 0.15fF
C9388 OR2X1_LOC_131/A D_INPUT_0 0.85fF
C9389 AND2X1_LOC_95/Y OR2X1_LOC_285/A 0.27fF
C9390 AND2X1_LOC_61/Y OR2X1_LOC_416/Y 0.03fF
C9391 OR2X1_LOC_431/a_8_216# OR2X1_LOC_59/Y 0.01fF
C9392 D_INPUT_5 OR2X1_LOC_378/Y 0.15fF
C9393 AND2X1_LOC_722/A OR2X1_LOC_74/A 0.09fF
C9394 OR2X1_LOC_283/Y OR2X1_LOC_278/Y 0.05fF
C9395 OR2X1_LOC_695/Y AND2X1_LOC_687/B 0.02fF
C9396 AND2X1_LOC_715/A AND2X1_LOC_116/B 0.01fF
C9397 AND2X1_LOC_557/Y AND2X1_LOC_554/Y 0.20fF
C9398 OR2X1_LOC_401/A OR2X1_LOC_78/B 0.01fF
C9399 AND2X1_LOC_787/a_36_24# AND2X1_LOC_784/A 0.00fF
C9400 AND2X1_LOC_131/a_8_24# D_INPUT_0 0.03fF
C9401 OR2X1_LOC_621/B OR2X1_LOC_532/B 0.20fF
C9402 OR2X1_LOC_377/A OR2X1_LOC_836/A 0.02fF
C9403 AND2X1_LOC_56/B OR2X1_LOC_541/B 0.04fF
C9404 AND2X1_LOC_174/a_8_24# AND2X1_LOC_650/Y 0.01fF
C9405 AND2X1_LOC_12/Y OR2X1_LOC_561/a_8_216# 0.01fF
C9406 OR2X1_LOC_395/a_8_216# OR2X1_LOC_80/A 0.09fF
C9407 OR2X1_LOC_19/B OR2X1_LOC_78/A 1.94fF
C9408 OR2X1_LOC_448/Y OR2X1_LOC_779/a_36_216# 0.00fF
C9409 OR2X1_LOC_805/A OR2X1_LOC_203/Y 0.07fF
C9410 AND2X1_LOC_318/a_8_24# OR2X1_LOC_6/A 0.01fF
C9411 AND2X1_LOC_36/Y OR2X1_LOC_546/A 0.53fF
C9412 OR2X1_LOC_429/Y OR2X1_LOC_2/Y 0.29fF
C9413 AND2X1_LOC_706/a_8_24# AND2X1_LOC_648/B 0.01fF
C9414 OR2X1_LOC_836/A AND2X1_LOC_824/B 0.01fF
C9415 OR2X1_LOC_835/A OR2X1_LOC_835/B 0.14fF
C9416 OR2X1_LOC_494/Y AND2X1_LOC_845/Y 0.12fF
C9417 OR2X1_LOC_22/Y OR2X1_LOC_25/Y 0.24fF
C9418 OR2X1_LOC_589/A AND2X1_LOC_648/B 0.01fF
C9419 AND2X1_LOC_541/Y D_INPUT_3 0.01fF
C9420 AND2X1_LOC_340/a_8_24# AND2X1_LOC_227/Y 0.03fF
C9421 AND2X1_LOC_59/Y AND2X1_LOC_252/a_8_24# 0.00fF
C9422 OR2X1_LOC_665/Y AND2X1_LOC_621/Y 0.07fF
C9423 INPUT_3 OR2X1_LOC_37/a_8_216# 0.02fF
C9424 AND2X1_LOC_621/Y AND2X1_LOC_474/Y 0.03fF
C9425 OR2X1_LOC_160/A AND2X1_LOC_329/a_8_24# 0.03fF
C9426 AND2X1_LOC_576/Y OR2X1_LOC_497/a_8_216# 0.03fF
C9427 AND2X1_LOC_319/A OR2X1_LOC_44/Y 0.07fF
C9428 OR2X1_LOC_36/Y OR2X1_LOC_69/a_8_216# 0.01fF
C9429 OR2X1_LOC_270/Y OR2X1_LOC_549/A 0.05fF
C9430 AND2X1_LOC_584/a_8_24# OR2X1_LOC_87/A 0.01fF
C9431 OR2X1_LOC_235/B AND2X1_LOC_134/a_8_24# 0.00fF
C9432 OR2X1_LOC_51/Y OR2X1_LOC_417/A 1.54fF
C9433 OR2X1_LOC_814/Y AND2X1_LOC_815/a_8_24# 0.23fF
C9434 OR2X1_LOC_154/A OR2X1_LOC_864/A 0.10fF
C9435 OR2X1_LOC_485/A AND2X1_LOC_621/Y 0.05fF
C9436 OR2X1_LOC_604/A AND2X1_LOC_851/B 0.10fF
C9437 AND2X1_LOC_191/Y OR2X1_LOC_616/a_36_216# 0.02fF
C9438 AND2X1_LOC_101/B OR2X1_LOC_85/A 0.21fF
C9439 AND2X1_LOC_738/B OR2X1_LOC_31/Y 0.15fF
C9440 OR2X1_LOC_251/Y OR2X1_LOC_669/A 0.01fF
C9441 OR2X1_LOC_849/A OR2X1_LOC_659/B 0.02fF
C9442 OR2X1_LOC_31/Y OR2X1_LOC_56/A 0.09fF
C9443 OR2X1_LOC_624/A OR2X1_LOC_216/a_36_216# 0.15fF
C9444 OR2X1_LOC_26/Y OR2X1_LOC_69/Y 0.00fF
C9445 OR2X1_LOC_121/B OR2X1_LOC_734/a_8_216# 0.01fF
C9446 OR2X1_LOC_405/A AND2X1_LOC_67/Y 0.02fF
C9447 OR2X1_LOC_864/A OR2X1_LOC_267/A 0.03fF
C9448 AND2X1_LOC_491/a_8_24# OR2X1_LOC_737/A 0.03fF
C9449 OR2X1_LOC_103/a_36_216# AND2X1_LOC_523/Y 0.01fF
C9450 AND2X1_LOC_591/a_8_24# OR2X1_LOC_593/B 0.01fF
C9451 OR2X1_LOC_41/a_36_216# OR2X1_LOC_13/Y 0.00fF
C9452 OR2X1_LOC_317/a_8_216# OR2X1_LOC_532/B 0.01fF
C9453 AND2X1_LOC_810/Y AND2X1_LOC_468/a_36_24# 0.00fF
C9454 AND2X1_LOC_12/Y OR2X1_LOC_285/B 0.01fF
C9455 AND2X1_LOC_717/B AND2X1_LOC_374/Y 0.13fF
C9456 AND2X1_LOC_516/a_8_24# OR2X1_LOC_155/A 0.03fF
C9457 OR2X1_LOC_294/Y OR2X1_LOC_736/a_8_216# 0.01fF
C9458 OR2X1_LOC_379/a_8_216# AND2X1_LOC_51/Y 0.14fF
C9459 AND2X1_LOC_40/Y D_INPUT_0 0.10fF
C9460 OR2X1_LOC_599/A OR2X1_LOC_74/A 0.03fF
C9461 AND2X1_LOC_367/A AND2X1_LOC_866/A 0.10fF
C9462 VDD OR2X1_LOC_289/Y 0.12fF
C9463 AND2X1_LOC_710/a_8_24# AND2X1_LOC_663/B 0.01fF
C9464 AND2X1_LOC_196/a_8_24# OR2X1_LOC_36/Y 0.01fF
C9465 AND2X1_LOC_31/Y OR2X1_LOC_435/A 0.01fF
C9466 OR2X1_LOC_403/B OR2X1_LOC_557/A 0.00fF
C9467 AND2X1_LOC_640/Y AND2X1_LOC_852/Y 2.74fF
C9468 OR2X1_LOC_351/B OR2X1_LOC_358/A 0.08fF
C9469 OR2X1_LOC_291/Y OR2X1_LOC_316/Y 0.02fF
C9470 OR2X1_LOC_43/A AND2X1_LOC_345/Y 0.07fF
C9471 AND2X1_LOC_697/a_8_24# OR2X1_LOC_269/B 0.11fF
C9472 OR2X1_LOC_46/A AND2X1_LOC_400/a_8_24# 0.01fF
C9473 OR2X1_LOC_680/A OR2X1_LOC_64/Y 1.55fF
C9474 OR2X1_LOC_52/a_8_216# OR2X1_LOC_44/Y 0.01fF
C9475 OR2X1_LOC_401/Y AND2X1_LOC_3/Y 0.79fF
C9476 OR2X1_LOC_856/B OR2X1_LOC_532/B 0.12fF
C9477 VDD OR2X1_LOC_247/Y 0.33fF
C9478 AND2X1_LOC_7/B OR2X1_LOC_732/A 0.03fF
C9479 AND2X1_LOC_489/Y AND2X1_LOC_717/B 0.09fF
C9480 AND2X1_LOC_86/B AND2X1_LOC_490/a_8_24# 0.04fF
C9481 AND2X1_LOC_666/a_8_24# OR2X1_LOC_269/B 0.01fF
C9482 OR2X1_LOC_40/Y AND2X1_LOC_222/Y 0.02fF
C9483 OR2X1_LOC_667/a_8_216# OR2X1_LOC_64/Y 0.07fF
C9484 OR2X1_LOC_629/a_8_216# AND2X1_LOC_3/Y 0.02fF
C9485 AND2X1_LOC_727/Y OR2X1_LOC_142/Y 0.06fF
C9486 OR2X1_LOC_409/B OR2X1_LOC_586/Y 0.00fF
C9487 OR2X1_LOC_537/A D_INPUT_0 0.01fF
C9488 OR2X1_LOC_427/A AND2X1_LOC_675/A 0.02fF
C9489 AND2X1_LOC_78/a_8_24# OR2X1_LOC_79/A 0.09fF
C9490 AND2X1_LOC_31/Y OR2X1_LOC_723/a_8_216# 0.01fF
C9491 OR2X1_LOC_26/Y OR2X1_LOC_43/a_8_216# 0.06fF
C9492 OR2X1_LOC_519/Y OR2X1_LOC_111/Y 0.00fF
C9493 OR2X1_LOC_280/Y OR2X1_LOC_279/Y 0.08fF
C9494 OR2X1_LOC_9/Y OR2X1_LOC_80/A 0.61fF
C9495 AND2X1_LOC_717/a_8_24# OR2X1_LOC_95/Y 0.03fF
C9496 AND2X1_LOC_852/Y OR2X1_LOC_416/Y 0.03fF
C9497 AND2X1_LOC_196/Y OR2X1_LOC_48/a_8_216# 0.47fF
C9498 AND2X1_LOC_679/a_8_24# OR2X1_LOC_715/A 0.02fF
C9499 OR2X1_LOC_331/A OR2X1_LOC_331/a_36_216# 0.00fF
C9500 AND2X1_LOC_450/a_8_24# AND2X1_LOC_451/Y 0.01fF
C9501 AND2X1_LOC_588/B D_INPUT_6 0.00fF
C9502 OR2X1_LOC_624/A OR2X1_LOC_218/Y 0.76fF
C9503 AND2X1_LOC_7/B OR2X1_LOC_539/B 0.02fF
C9504 OR2X1_LOC_16/A OR2X1_LOC_536/a_36_216# 0.00fF
C9505 VDD OR2X1_LOC_534/a_8_216# 0.21fF
C9506 OR2X1_LOC_665/a_8_216# OR2X1_LOC_89/A 0.00fF
C9507 OR2X1_LOC_16/A OR2X1_LOC_300/Y 0.10fF
C9508 OR2X1_LOC_529/a_8_216# D_INPUT_3 0.06fF
C9509 AND2X1_LOC_587/a_36_24# INPUT_6 0.00fF
C9510 INPUT_3 OR2X1_LOC_62/A 0.53fF
C9511 AND2X1_LOC_44/Y OR2X1_LOC_523/A 0.01fF
C9512 OR2X1_LOC_181/B OR2X1_LOC_223/A 0.00fF
C9513 AND2X1_LOC_66/a_8_24# OR2X1_LOC_26/Y 0.17fF
C9514 OR2X1_LOC_95/Y AND2X1_LOC_458/Y 0.00fF
C9515 AND2X1_LOC_570/Y AND2X1_LOC_657/A 0.00fF
C9516 OR2X1_LOC_417/Y AND2X1_LOC_390/B 0.07fF
C9517 OR2X1_LOC_70/Y OR2X1_LOC_431/a_8_216# 0.08fF
C9518 OR2X1_LOC_516/Y AND2X1_LOC_242/a_8_24# 0.02fF
C9519 AND2X1_LOC_170/B OR2X1_LOC_44/Y 0.03fF
C9520 AND2X1_LOC_390/B OR2X1_LOC_311/Y 0.06fF
C9521 OR2X1_LOC_185/A D_INPUT_1 0.07fF
C9522 OR2X1_LOC_349/B OR2X1_LOC_349/A 0.10fF
C9523 OR2X1_LOC_605/a_36_216# OR2X1_LOC_121/B 0.00fF
C9524 AND2X1_LOC_66/a_8_24# OR2X1_LOC_89/A 0.09fF
C9525 OR2X1_LOC_190/A OR2X1_LOC_367/B 0.31fF
C9526 AND2X1_LOC_42/B OR2X1_LOC_62/B 0.22fF
C9527 AND2X1_LOC_390/B AND2X1_LOC_538/Y 0.02fF
C9528 OR2X1_LOC_22/Y OR2X1_LOC_279/Y 0.16fF
C9529 OR2X1_LOC_43/A AND2X1_LOC_649/Y 0.12fF
C9530 AND2X1_LOC_137/a_8_24# OR2X1_LOC_26/Y 0.04fF
C9531 AND2X1_LOC_43/B OR2X1_LOC_214/B 0.00fF
C9532 AND2X1_LOC_139/A AND2X1_LOC_361/A 0.04fF
C9533 OR2X1_LOC_36/Y OR2X1_LOC_619/a_8_216# 0.03fF
C9534 AND2X1_LOC_43/B OR2X1_LOC_241/B 0.04fF
C9535 AND2X1_LOC_866/A OR2X1_LOC_757/a_8_216# 0.02fF
C9536 OR2X1_LOC_613/Y AND2X1_LOC_620/Y 0.01fF
C9537 OR2X1_LOC_362/B OR2X1_LOC_580/a_8_216# 0.01fF
C9538 OR2X1_LOC_702/A AND2X1_LOC_47/Y 0.03fF
C9539 D_INPUT_5 OR2X1_LOC_378/A 0.30fF
C9540 OR2X1_LOC_639/B OR2X1_LOC_451/B 0.19fF
C9541 AND2X1_LOC_866/A OR2X1_LOC_74/A 0.07fF
C9542 AND2X1_LOC_721/A OR2X1_LOC_44/Y 0.03fF
C9543 OR2X1_LOC_161/A OR2X1_LOC_675/Y 0.06fF
C9544 OR2X1_LOC_245/a_36_216# OR2X1_LOC_246/A 0.07fF
C9545 AND2X1_LOC_12/Y OR2X1_LOC_358/A 0.36fF
C9546 OR2X1_LOC_91/A AND2X1_LOC_212/a_36_24# 0.01fF
C9547 OR2X1_LOC_100/a_36_216# OR2X1_LOC_608/Y 0.00fF
C9548 OR2X1_LOC_824/a_8_216# D_INPUT_3 0.01fF
C9549 OR2X1_LOC_35/Y OR2X1_LOC_771/B 0.03fF
C9550 AND2X1_LOC_554/B OR2X1_LOC_47/Y 0.02fF
C9551 AND2X1_LOC_663/B OR2X1_LOC_95/Y 0.17fF
C9552 OR2X1_LOC_56/A OR2X1_LOC_320/a_8_216# 0.01fF
C9553 OR2X1_LOC_69/Y AND2X1_LOC_202/a_8_24# 0.00fF
C9554 AND2X1_LOC_191/B AND2X1_LOC_791/a_8_24# 0.01fF
C9555 OR2X1_LOC_16/A AND2X1_LOC_219/A 0.11fF
C9556 OR2X1_LOC_87/A OR2X1_LOC_641/B 0.39fF
C9557 OR2X1_LOC_139/A AND2X1_LOC_150/a_8_24# 0.11fF
C9558 OR2X1_LOC_358/B OR2X1_LOC_228/Y 0.02fF
C9559 OR2X1_LOC_607/Y OR2X1_LOC_46/A 0.02fF
C9560 OR2X1_LOC_44/Y OR2X1_LOC_331/Y 0.07fF
C9561 VDD AND2X1_LOC_783/B 0.06fF
C9562 AND2X1_LOC_564/B AND2X1_LOC_778/Y 0.02fF
C9563 AND2X1_LOC_714/B OR2X1_LOC_428/A 0.12fF
C9564 AND2X1_LOC_40/Y OR2X1_LOC_339/A 0.12fF
C9565 AND2X1_LOC_71/a_8_24# OR2X1_LOC_844/B 0.00fF
C9566 VDD AND2X1_LOC_258/a_8_24# -0.00fF
C9567 OR2X1_LOC_599/A AND2X1_LOC_783/a_8_24# 0.03fF
C9568 OR2X1_LOC_220/B OR2X1_LOC_550/B 0.00fF
C9569 AND2X1_LOC_64/Y OR2X1_LOC_648/A 0.07fF
C9570 AND2X1_LOC_91/B OR2X1_LOC_645/a_8_216# 0.03fF
C9571 OR2X1_LOC_864/A OR2X1_LOC_560/A 0.14fF
C9572 OR2X1_LOC_7/A AND2X1_LOC_222/Y 0.03fF
C9573 OR2X1_LOC_736/Y OR2X1_LOC_346/A 0.79fF
C9574 OR2X1_LOC_26/Y AND2X1_LOC_796/A 0.10fF
C9575 AND2X1_LOC_674/a_8_24# OR2X1_LOC_374/Y 0.02fF
C9576 AND2X1_LOC_852/Y OR2X1_LOC_80/A 0.07fF
C9577 OR2X1_LOC_132/Y OR2X1_LOC_134/Y 0.11fF
C9578 OR2X1_LOC_676/a_8_216# OR2X1_LOC_161/B 0.03fF
C9579 OR2X1_LOC_676/Y AND2X1_LOC_44/Y 0.09fF
C9580 VDD OR2X1_LOC_708/a_8_216# 0.21fF
C9581 OR2X1_LOC_89/A AND2X1_LOC_796/A 0.03fF
C9582 OR2X1_LOC_502/A OR2X1_LOC_510/a_8_216# 0.01fF
C9583 AND2X1_LOC_858/B AND2X1_LOC_242/B 0.83fF
C9584 OR2X1_LOC_167/Y OR2X1_LOC_47/Y 0.01fF
C9585 OR2X1_LOC_78/B AND2X1_LOC_7/B 0.16fF
C9586 OR2X1_LOC_476/B OR2X1_LOC_598/A 0.01fF
C9587 OR2X1_LOC_778/Y OR2X1_LOC_446/B 0.14fF
C9588 AND2X1_LOC_740/B AND2X1_LOC_742/A 0.01fF
C9589 AND2X1_LOC_848/a_8_24# AND2X1_LOC_789/Y 0.01fF
C9590 OR2X1_LOC_56/A AND2X1_LOC_464/A 0.03fF
C9591 OR2X1_LOC_6/B AND2X1_LOC_262/a_8_24# 0.06fF
C9592 OR2X1_LOC_834/A AND2X1_LOC_44/Y 0.01fF
C9593 OR2X1_LOC_696/A AND2X1_LOC_832/a_8_24# 0.03fF
C9594 AND2X1_LOC_707/Y OR2X1_LOC_91/A 0.03fF
C9595 OR2X1_LOC_778/Y OR2X1_LOC_303/B 0.05fF
C9596 OR2X1_LOC_585/A OR2X1_LOC_150/a_8_216# 0.01fF
C9597 OR2X1_LOC_676/Y OR2X1_LOC_514/a_8_216# 0.03fF
C9598 AND2X1_LOC_1/Y AND2X1_LOC_430/B 0.09fF
C9599 OR2X1_LOC_7/A OR2X1_LOC_423/Y 0.05fF
C9600 AND2X1_LOC_392/A AND2X1_LOC_212/A 0.04fF
C9601 OR2X1_LOC_485/A OR2X1_LOC_71/A 0.54fF
C9602 AND2X1_LOC_663/A AND2X1_LOC_727/B 0.73fF
C9603 AND2X1_LOC_571/A OR2X1_LOC_427/A 0.01fF
C9604 AND2X1_LOC_18/Y AND2X1_LOC_265/a_8_24# 0.13fF
C9605 OR2X1_LOC_756/B OR2X1_LOC_576/A 0.02fF
C9606 AND2X1_LOC_658/B AND2X1_LOC_476/Y 0.07fF
C9607 OR2X1_LOC_715/B OR2X1_LOC_66/A 0.08fF
C9608 OR2X1_LOC_494/A OR2X1_LOC_92/Y 0.02fF
C9609 OR2X1_LOC_158/A OR2X1_LOC_743/a_8_216# 0.01fF
C9610 OR2X1_LOC_335/Y AND2X1_LOC_438/a_8_24# 0.03fF
C9611 D_INPUT_3 AND2X1_LOC_8/a_36_24# 0.01fF
C9612 AND2X1_LOC_371/a_8_24# VDD 0.00fF
C9613 OR2X1_LOC_756/Y OR2X1_LOC_756/a_8_216# 0.01fF
C9614 VDD AND2X1_LOC_18/Y 1.16fF
C9615 OR2X1_LOC_154/A OR2X1_LOC_714/a_36_216# 0.00fF
C9616 OR2X1_LOC_784/B OR2X1_LOC_66/A 0.01fF
C9617 AND2X1_LOC_60/a_8_24# OR2X1_LOC_61/B 0.01fF
C9618 AND2X1_LOC_501/Y VDD 0.01fF
C9619 AND2X1_LOC_719/Y OR2X1_LOC_329/B 0.10fF
C9620 AND2X1_LOC_454/A AND2X1_LOC_449/a_36_24# 0.00fF
C9621 OR2X1_LOC_273/a_8_216# OR2X1_LOC_300/Y 0.39fF
C9622 OR2X1_LOC_756/B OR2X1_LOC_439/B 0.00fF
C9623 OR2X1_LOC_666/a_36_216# OR2X1_LOC_51/Y 0.00fF
C9624 AND2X1_LOC_110/Y OR2X1_LOC_78/A 0.03fF
C9625 AND2X1_LOC_570/Y VDD 0.52fF
C9626 OR2X1_LOC_92/a_36_216# AND2X1_LOC_647/Y 0.00fF
C9627 OR2X1_LOC_473/A OR2X1_LOC_66/Y 0.02fF
C9628 OR2X1_LOC_331/A VDD 0.03fF
C9629 AND2X1_LOC_40/Y OR2X1_LOC_673/B 0.03fF
C9630 OR2X1_LOC_58/Y OR2X1_LOC_59/Y 0.01fF
C9631 OR2X1_LOC_858/B OR2X1_LOC_349/A 0.02fF
C9632 OR2X1_LOC_197/A OR2X1_LOC_197/a_8_216# 0.47fF
C9633 AND2X1_LOC_92/a_8_24# AND2X1_LOC_95/Y 0.17fF
C9634 AND2X1_LOC_564/B AND2X1_LOC_624/A 0.07fF
C9635 OR2X1_LOC_502/A AND2X1_LOC_65/A 0.06fF
C9636 OR2X1_LOC_161/A OR2X1_LOC_779/A 0.03fF
C9637 AND2X1_LOC_456/B OR2X1_LOC_253/Y 0.79fF
C9638 OR2X1_LOC_40/Y AND2X1_LOC_367/A 0.05fF
C9639 OR2X1_LOC_130/A AND2X1_LOC_224/a_8_24# 0.03fF
C9640 OR2X1_LOC_589/A OR2X1_LOC_265/a_8_216# 0.01fF
C9641 AND2X1_LOC_130/a_36_24# OR2X1_LOC_517/A 0.00fF
C9642 OR2X1_LOC_147/B OR2X1_LOC_486/Y 0.08fF
C9643 AND2X1_LOC_40/Y OR2X1_LOC_831/A 0.03fF
C9644 OR2X1_LOC_375/A AND2X1_LOC_7/B 0.25fF
C9645 OR2X1_LOC_619/Y AND2X1_LOC_210/a_8_24# 0.01fF
C9646 AND2X1_LOC_748/a_8_24# OR2X1_LOC_691/Y 0.01fF
C9647 OR2X1_LOC_18/Y AND2X1_LOC_786/Y 0.24fF
C9648 OR2X1_LOC_87/A OR2X1_LOC_227/A 0.03fF
C9649 OR2X1_LOC_154/A OR2X1_LOC_121/A 0.03fF
C9650 AND2X1_LOC_830/a_8_24# OR2X1_LOC_142/Y 0.03fF
C9651 OR2X1_LOC_147/B OR2X1_LOC_711/a_8_216# 0.14fF
C9652 OR2X1_LOC_30/a_36_216# INPUT_7 0.00fF
C9653 OR2X1_LOC_382/Y OR2X1_LOC_600/A 0.03fF
C9654 OR2X1_LOC_485/Y OR2X1_LOC_516/B 0.24fF
C9655 OR2X1_LOC_287/a_8_216# OR2X1_LOC_366/Y 0.02fF
C9656 OR2X1_LOC_151/A AND2X1_LOC_321/a_8_24# 0.04fF
C9657 AND2X1_LOC_40/Y OR2X1_LOC_598/Y 0.01fF
C9658 OR2X1_LOC_510/A OR2X1_LOC_502/A 0.16fF
C9659 AND2X1_LOC_40/Y AND2X1_LOC_505/a_8_24# 0.10fF
C9660 AND2X1_LOC_484/a_36_24# AND2X1_LOC_36/Y 0.01fF
C9661 INPUT_1 OR2X1_LOC_437/A 0.39fF
C9662 OR2X1_LOC_45/B AND2X1_LOC_319/A 0.07fF
C9663 OR2X1_LOC_333/B OR2X1_LOC_333/a_8_216# 0.03fF
C9664 AND2X1_LOC_776/Y OR2X1_LOC_238/Y 0.02fF
C9665 OR2X1_LOC_462/B AND2X1_LOC_44/Y 0.01fF
C9666 OR2X1_LOC_659/B OR2X1_LOC_572/a_8_216# 0.40fF
C9667 OR2X1_LOC_657/a_8_216# OR2X1_LOC_576/A 0.01fF
C9668 OR2X1_LOC_53/Y OR2X1_LOC_753/A 0.03fF
C9669 AND2X1_LOC_721/Y OR2X1_LOC_497/Y 0.04fF
C9670 OR2X1_LOC_614/Y OR2X1_LOC_161/A 0.03fF
C9671 OR2X1_LOC_528/Y AND2X1_LOC_805/Y 0.15fF
C9672 AND2X1_LOC_70/Y OR2X1_LOC_216/A 0.01fF
C9673 AND2X1_LOC_773/Y OR2X1_LOC_36/Y 0.03fF
C9674 GATE_811 OR2X1_LOC_152/a_8_216# 0.48fF
C9675 AND2X1_LOC_349/a_8_24# OR2X1_LOC_12/Y 0.05fF
C9676 OR2X1_LOC_369/Y AND2X1_LOC_716/Y -0.02fF
C9677 OR2X1_LOC_391/B OR2X1_LOC_489/A 0.00fF
C9678 OR2X1_LOC_377/A OR2X1_LOC_648/B 0.10fF
C9679 OR2X1_LOC_319/B OR2X1_LOC_78/B 0.04fF
C9680 AND2X1_LOC_363/B OR2X1_LOC_56/A 0.02fF
C9681 OR2X1_LOC_756/B AND2X1_LOC_41/A 0.18fF
C9682 AND2X1_LOC_31/Y OR2X1_LOC_737/a_8_216# 0.01fF
C9683 OR2X1_LOC_174/A OR2X1_LOC_434/a_8_216# 0.00fF
C9684 AND2X1_LOC_810/A AND2X1_LOC_854/a_8_24# 0.01fF
C9685 AND2X1_LOC_706/Y OR2X1_LOC_433/a_8_216# 0.04fF
C9686 OR2X1_LOC_792/B OR2X1_LOC_792/Y 0.89fF
C9687 VDD OR2X1_LOC_807/B -0.00fF
C9688 AND2X1_LOC_554/Y AND2X1_LOC_563/A 0.01fF
C9689 OR2X1_LOC_78/A OR2X1_LOC_712/a_36_216# 0.00fF
C9690 OR2X1_LOC_585/A AND2X1_LOC_774/A 0.03fF
C9691 OR2X1_LOC_160/B OR2X1_LOC_803/B 0.03fF
C9692 AND2X1_LOC_264/a_36_24# OR2X1_LOC_12/Y 0.01fF
C9693 AND2X1_LOC_828/a_8_24# OR2X1_LOC_52/B 0.02fF
C9694 OR2X1_LOC_686/B AND2X1_LOC_43/B 0.01fF
C9695 OR2X1_LOC_335/Y AND2X1_LOC_40/Y 0.03fF
C9696 INPUT_3 OR2X1_LOC_8/Y 0.05fF
C9697 OR2X1_LOC_318/Y OR2X1_LOC_78/B 0.03fF
C9698 AND2X1_LOC_161/a_8_24# OR2X1_LOC_51/Y 0.00fF
C9699 OR2X1_LOC_778/A OR2X1_LOC_121/A 0.02fF
C9700 OR2X1_LOC_486/Y AND2X1_LOC_298/a_36_24# 0.01fF
C9701 OR2X1_LOC_177/a_36_216# OR2X1_LOC_52/B 0.03fF
C9702 OR2X1_LOC_9/Y OR2X1_LOC_6/A 0.48fF
C9703 OR2X1_LOC_751/A AND2X1_LOC_750/a_8_24# 0.10fF
C9704 OR2X1_LOC_753/Y AND2X1_LOC_562/Y 0.10fF
C9705 OR2X1_LOC_447/Y OR2X1_LOC_703/Y 0.00fF
C9706 OR2X1_LOC_57/a_8_216# OR2X1_LOC_44/Y 0.01fF
C9707 OR2X1_LOC_323/A AND2X1_LOC_464/Y 0.01fF
C9708 VDD AND2X1_LOC_123/Y 0.02fF
C9709 AND2X1_LOC_807/Y AND2X1_LOC_807/B 0.13fF
C9710 VDD OR2X1_LOC_500/A 0.07fF
C9711 OR2X1_LOC_143/a_8_216# D_INPUT_0 0.01fF
C9712 OR2X1_LOC_482/Y OR2X1_LOC_497/Y 0.01fF
C9713 OR2X1_LOC_91/A AND2X1_LOC_841/B 0.07fF
C9714 OR2X1_LOC_26/Y OR2X1_LOC_13/Y 0.02fF
C9715 OR2X1_LOC_96/Y OR2X1_LOC_85/A 0.03fF
C9716 OR2X1_LOC_70/Y AND2X1_LOC_636/a_8_24# 0.05fF
C9717 AND2X1_LOC_40/Y OR2X1_LOC_435/a_36_216# 0.00fF
C9718 OR2X1_LOC_673/a_36_216# AND2X1_LOC_8/Y 0.00fF
C9719 OR2X1_LOC_18/Y AND2X1_LOC_218/Y 0.00fF
C9720 OR2X1_LOC_653/Y OR2X1_LOC_174/A 0.00fF
C9721 OR2X1_LOC_190/A OR2X1_LOC_456/Y 0.03fF
C9722 OR2X1_LOC_541/B AND2X1_LOC_92/Y 0.02fF
C9723 OR2X1_LOC_391/B OR2X1_LOC_772/A 0.01fF
C9724 OR2X1_LOC_177/a_8_216# OR2X1_LOC_74/A 0.02fF
C9725 AND2X1_LOC_550/A AND2X1_LOC_444/a_8_24# 0.07fF
C9726 AND2X1_LOC_784/A AND2X1_LOC_357/B 0.02fF
C9727 AND2X1_LOC_803/B AND2X1_LOC_192/Y 0.03fF
C9728 AND2X1_LOC_721/Y AND2X1_LOC_844/a_8_24# 0.17fF
C9729 OR2X1_LOC_596/Y VDD 0.16fF
C9730 OR2X1_LOC_170/A VDD -0.00fF
C9731 OR2X1_LOC_114/a_36_216# AND2X1_LOC_95/Y 0.00fF
C9732 OR2X1_LOC_805/A OR2X1_LOC_78/B 0.03fF
C9733 AND2X1_LOC_675/Y OR2X1_LOC_39/A 0.00fF
C9734 OR2X1_LOC_664/Y OR2X1_LOC_78/A 0.07fF
C9735 OR2X1_LOC_160/A OR2X1_LOC_235/B 0.19fF
C9736 VDD OR2X1_LOC_469/a_8_216# 0.21fF
C9737 OR2X1_LOC_40/Y AND2X1_LOC_673/a_8_24# 0.01fF
C9738 AND2X1_LOC_110/Y OR2X1_LOC_155/A 0.03fF
C9739 AND2X1_LOC_706/Y OR2X1_LOC_70/Y 0.05fF
C9740 OR2X1_LOC_45/B AND2X1_LOC_708/a_8_24# 0.01fF
C9741 OR2X1_LOC_476/B OR2X1_LOC_34/A -0.00fF
C9742 OR2X1_LOC_377/A AND2X1_LOC_232/a_36_24# 0.00fF
C9743 AND2X1_LOC_219/Y OR2X1_LOC_265/Y 0.07fF
C9744 AND2X1_LOC_70/Y OR2X1_LOC_468/Y 0.03fF
C9745 OR2X1_LOC_600/a_8_216# OR2X1_LOC_43/A 0.15fF
C9746 OR2X1_LOC_91/Y OR2X1_LOC_744/A 0.07fF
C9747 AND2X1_LOC_303/A OR2X1_LOC_59/Y 4.37fF
C9748 OR2X1_LOC_92/Y OR2X1_LOC_427/A 0.69fF
C9749 OR2X1_LOC_3/Y OR2X1_LOC_382/a_8_216# 0.06fF
C9750 OR2X1_LOC_466/A OR2X1_LOC_449/B 0.21fF
C9751 OR2X1_LOC_11/Y OR2X1_LOC_26/a_36_216# 0.00fF
C9752 OR2X1_LOC_426/B OR2X1_LOC_117/Y 0.42fF
C9753 AND2X1_LOC_541/Y AND2X1_LOC_276/Y 0.17fF
C9754 OR2X1_LOC_604/A OR2X1_LOC_73/a_8_216# 0.02fF
C9755 OR2X1_LOC_808/B OR2X1_LOC_161/A 0.04fF
C9756 OR2X1_LOC_160/B OR2X1_LOC_141/B 0.12fF
C9757 OR2X1_LOC_40/Y OR2X1_LOC_74/A 1.74fF
C9758 OR2X1_LOC_107/a_36_216# OR2X1_LOC_44/Y 0.02fF
C9759 OR2X1_LOC_49/A OR2X1_LOC_54/Y 0.60fF
C9760 OR2X1_LOC_772/Y OR2X1_LOC_489/A 0.21fF
C9761 OR2X1_LOC_516/B OR2X1_LOC_39/A 0.28fF
C9762 OR2X1_LOC_81/Y OR2X1_LOC_59/Y 0.03fF
C9763 OR2X1_LOC_614/Y AND2X1_LOC_51/Y 0.01fF
C9764 OR2X1_LOC_417/Y OR2X1_LOC_604/Y 0.23fF
C9765 AND2X1_LOC_377/Y OR2X1_LOC_36/Y 0.08fF
C9766 OR2X1_LOC_663/A OR2X1_LOC_130/A 0.01fF
C9767 OR2X1_LOC_369/Y OR2X1_LOC_312/Y 0.05fF
C9768 AND2X1_LOC_477/A OR2X1_LOC_428/A 0.12fF
C9769 OR2X1_LOC_235/B OR2X1_LOC_235/a_36_216# 0.03fF
C9770 AND2X1_LOC_456/B AND2X1_LOC_286/Y 0.58fF
C9771 AND2X1_LOC_43/B AND2X1_LOC_423/a_8_24# 0.01fF
C9772 OR2X1_LOC_805/A OR2X1_LOC_721/Y 0.02fF
C9773 OR2X1_LOC_261/a_8_216# OR2X1_LOC_817/a_8_216# 0.47fF
C9774 OR2X1_LOC_600/A OR2X1_LOC_817/a_36_216# 0.00fF
C9775 OR2X1_LOC_427/A OR2X1_LOC_257/a_8_216# 0.00fF
C9776 AND2X1_LOC_605/Y OR2X1_LOC_44/Y 0.02fF
C9777 OR2X1_LOC_703/A OR2X1_LOC_468/Y 0.03fF
C9778 OR2X1_LOC_665/Y OR2X1_LOC_59/Y 0.00fF
C9779 OR2X1_LOC_604/A AND2X1_LOC_260/a_8_24# 0.05fF
C9780 OR2X1_LOC_282/a_8_216# AND2X1_LOC_285/Y 0.00fF
C9781 AND2X1_LOC_312/a_36_24# OR2X1_LOC_87/A 0.01fF
C9782 OR2X1_LOC_495/Y OR2X1_LOC_237/Y 0.24fF
C9783 OR2X1_LOC_668/a_36_216# OR2X1_LOC_161/A 0.00fF
C9784 AND2X1_LOC_95/Y OR2X1_LOC_185/A 0.12fF
C9785 AND2X1_LOC_56/B OR2X1_LOC_637/A 0.17fF
C9786 OR2X1_LOC_485/A OR2X1_LOC_59/Y 1.11fF
C9787 AND2X1_LOC_712/Y AND2X1_LOC_712/B 0.06fF
C9788 OR2X1_LOC_429/Y OR2X1_LOC_25/Y 0.01fF
C9789 AND2X1_LOC_689/a_8_24# OR2X1_LOC_66/A 0.17fF
C9790 AND2X1_LOC_593/a_36_24# OR2X1_LOC_64/Y 0.00fF
C9791 AND2X1_LOC_367/A OR2X1_LOC_7/A 3.62fF
C9792 OR2X1_LOC_63/a_8_216# OR2X1_LOC_65/B 0.02fF
C9793 OR2X1_LOC_235/B AND2X1_LOC_86/B 0.02fF
C9794 OR2X1_LOC_662/A OR2X1_LOC_660/B 0.03fF
C9795 OR2X1_LOC_654/a_8_216# D_INPUT_0 0.02fF
C9796 AND2X1_LOC_70/Y AND2X1_LOC_1/Y 0.00fF
C9797 OR2X1_LOC_499/B AND2X1_LOC_3/Y 0.02fF
C9798 AND2X1_LOC_363/A OR2X1_LOC_92/Y 0.39fF
C9799 OR2X1_LOC_447/Y OR2X1_LOC_596/A 0.08fF
C9800 OR2X1_LOC_421/A OR2X1_LOC_22/Y 0.11fF
C9801 AND2X1_LOC_392/A AND2X1_LOC_727/A 0.03fF
C9802 OR2X1_LOC_186/Y OR2X1_LOC_436/Y 0.02fF
C9803 OR2X1_LOC_792/Y OR2X1_LOC_269/B 0.19fF
C9804 OR2X1_LOC_771/B OR2X1_LOC_80/A 0.03fF
C9805 OR2X1_LOC_762/Y AND2X1_LOC_651/B 0.13fF
C9806 OR2X1_LOC_659/A AND2X1_LOC_42/B 0.08fF
C9807 OR2X1_LOC_805/A OR2X1_LOC_375/A 0.07fF
C9808 OR2X1_LOC_847/A AND2X1_LOC_817/a_8_24# 0.01fF
C9809 AND2X1_LOC_207/a_8_24# AND2X1_LOC_729/B 0.01fF
C9810 OR2X1_LOC_154/A OR2X1_LOC_738/A 0.31fF
C9811 OR2X1_LOC_87/A OR2X1_LOC_739/A 0.03fF
C9812 OR2X1_LOC_417/Y OR2X1_LOC_744/A 0.03fF
C9813 OR2X1_LOC_165/a_36_216# OR2X1_LOC_26/Y 0.02fF
C9814 OR2X1_LOC_673/Y AND2X1_LOC_132/a_8_24# 0.01fF
C9815 OR2X1_LOC_291/Y OR2X1_LOC_744/A 0.03fF
C9816 AND2X1_LOC_31/Y AND2X1_LOC_409/B 0.03fF
C9817 OR2X1_LOC_196/B OR2X1_LOC_702/a_36_216# 0.02fF
C9818 OR2X1_LOC_846/a_36_216# OR2X1_LOC_848/A 0.00fF
C9819 OR2X1_LOC_20/Y D_INPUT_0 0.02fF
C9820 AND2X1_LOC_86/Y OR2X1_LOC_84/B 1.40fF
C9821 OR2X1_LOC_763/Y OR2X1_LOC_48/B 0.01fF
C9822 OR2X1_LOC_364/A OR2X1_LOC_130/A 0.03fF
C9823 OR2X1_LOC_185/Y OR2X1_LOC_130/A 0.08fF
C9824 VDD OR2X1_LOC_813/A 0.12fF
C9825 OR2X1_LOC_91/Y AND2X1_LOC_840/B 0.10fF
C9826 OR2X1_LOC_708/B OR2X1_LOC_161/A 0.10fF
C9827 AND2X1_LOC_452/Y OR2X1_LOC_52/B 0.01fF
C9828 AND2X1_LOC_490/a_8_24# OR2X1_LOC_847/A 0.06fF
C9829 OR2X1_LOC_763/Y OR2X1_LOC_18/Y 0.00fF
C9830 OR2X1_LOC_808/B AND2X1_LOC_51/Y 0.03fF
C9831 OR2X1_LOC_648/A AND2X1_LOC_600/a_8_24# 0.24fF
C9832 OR2X1_LOC_297/a_8_216# AND2X1_LOC_663/B 0.01fF
C9833 OR2X1_LOC_6/B OR2X1_LOC_276/A 0.04fF
C9834 OR2X1_LOC_96/B OR2X1_LOC_6/A 0.01fF
C9835 AND2X1_LOC_392/A OR2X1_LOC_95/Y 0.03fF
C9836 OR2X1_LOC_19/B OR2X1_LOC_394/a_8_216# 0.04fF
C9837 OR2X1_LOC_32/B OR2X1_LOC_32/a_8_216# 0.03fF
C9838 AND2X1_LOC_191/B OR2X1_LOC_71/Y 0.03fF
C9839 OR2X1_LOC_47/Y AND2X1_LOC_476/Y 0.16fF
C9840 AND2X1_LOC_565/B OR2X1_LOC_95/Y 0.01fF
C9841 AND2X1_LOC_362/B OR2X1_LOC_47/Y 0.24fF
C9842 OR2X1_LOC_95/Y AND2X1_LOC_807/B 1.05fF
C9843 OR2X1_LOC_773/B OR2X1_LOC_287/B 0.00fF
C9844 AND2X1_LOC_350/a_8_24# OR2X1_LOC_289/Y 0.24fF
C9845 OR2X1_LOC_200/a_8_216# OR2X1_LOC_87/A 0.07fF
C9846 OR2X1_LOC_102/a_8_216# AND2X1_LOC_721/A 0.01fF
C9847 OR2X1_LOC_756/B OR2X1_LOC_403/a_8_216# 0.02fF
C9848 OR2X1_LOC_383/Y OR2X1_LOC_391/A 0.05fF
C9849 AND2X1_LOC_456/B OR2X1_LOC_22/Y 0.06fF
C9850 OR2X1_LOC_87/A OR2X1_LOC_269/B 0.08fF
C9851 AND2X1_LOC_563/a_8_24# OR2X1_LOC_89/A 0.01fF
C9852 OR2X1_LOC_643/A OR2X1_LOC_659/B 0.06fF
C9853 AND2X1_LOC_578/A OR2X1_LOC_18/Y 0.10fF
C9854 AND2X1_LOC_56/B OR2X1_LOC_778/Y 0.10fF
C9855 OR2X1_LOC_418/a_36_216# AND2X1_LOC_452/Y 0.01fF
C9856 AND2X1_LOC_95/Y OR2X1_LOC_435/Y 0.13fF
C9857 OR2X1_LOC_757/A OR2X1_LOC_417/A 0.02fF
C9858 OR2X1_LOC_663/A OR2X1_LOC_62/B 0.03fF
C9859 OR2X1_LOC_838/a_8_216# OR2X1_LOC_46/A 0.02fF
C9860 AND2X1_LOC_35/Y OR2X1_LOC_7/A 0.51fF
C9861 OR2X1_LOC_83/Y OR2X1_LOC_6/A 0.00fF
C9862 OR2X1_LOC_358/a_8_216# AND2X1_LOC_3/Y 0.05fF
C9863 AND2X1_LOC_106/a_36_24# OR2X1_LOC_66/A 0.00fF
C9864 AND2X1_LOC_572/Y AND2X1_LOC_557/a_8_24# 0.19fF
C9865 OR2X1_LOC_472/A AND2X1_LOC_56/B 0.03fF
C9866 OR2X1_LOC_845/A AND2X1_LOC_18/Y 0.07fF
C9867 AND2X1_LOC_712/B OR2X1_LOC_422/Y 0.12fF
C9868 OR2X1_LOC_6/B OR2X1_LOC_84/a_36_216# 0.00fF
C9869 OR2X1_LOC_46/A OR2X1_LOC_23/a_8_216# 0.01fF
C9870 OR2X1_LOC_3/Y AND2X1_LOC_266/Y 0.15fF
C9871 OR2X1_LOC_486/Y OR2X1_LOC_318/B 0.12fF
C9872 OR2X1_LOC_123/a_8_216# OR2X1_LOC_786/Y 0.01fF
C9873 OR2X1_LOC_193/A AND2X1_LOC_43/B 0.01fF
C9874 OR2X1_LOC_744/A D_INPUT_3 0.09fF
C9875 AND2X1_LOC_354/Y AND2X1_LOC_727/A 0.01fF
C9876 AND2X1_LOC_64/Y OR2X1_LOC_704/a_8_216# 0.01fF
C9877 AND2X1_LOC_91/B OR2X1_LOC_446/B 0.03fF
C9878 AND2X1_LOC_262/a_8_24# OR2X1_LOC_598/A 0.02fF
C9879 AND2X1_LOC_476/Y AND2X1_LOC_405/a_36_24# 0.00fF
C9880 AND2X1_LOC_749/a_36_24# D_INPUT_0 0.00fF
C9881 OR2X1_LOC_188/Y OR2X1_LOC_367/B 0.03fF
C9882 OR2X1_LOC_278/A OR2X1_LOC_118/Y 0.38fF
C9883 AND2X1_LOC_393/a_8_24# OR2X1_LOC_624/B 0.02fF
C9884 AND2X1_LOC_753/B AND2X1_LOC_53/Y 0.12fF
C9885 AND2X1_LOC_70/Y OR2X1_LOC_205/Y 0.10fF
C9886 OR2X1_LOC_114/B AND2X1_LOC_497/a_8_24# 0.01fF
C9887 OR2X1_LOC_647/A AND2X1_LOC_8/Y 0.03fF
C9888 OR2X1_LOC_175/B OR2X1_LOC_532/B 0.00fF
C9889 OR2X1_LOC_542/a_8_216# OR2X1_LOC_543/a_8_216# 0.47fF
C9890 AND2X1_LOC_456/Y OR2X1_LOC_7/A 0.01fF
C9891 OR2X1_LOC_40/Y AND2X1_LOC_647/Y 0.33fF
C9892 AND2X1_LOC_345/Y AND2X1_LOC_818/a_36_24# 0.01fF
C9893 OR2X1_LOC_345/Y OR2X1_LOC_348/B 0.00fF
C9894 OR2X1_LOC_527/Y AND2X1_LOC_840/B 0.10fF
C9895 AND2X1_LOC_191/Y AND2X1_LOC_474/Y 9.02fF
C9896 OR2X1_LOC_87/A OR2X1_LOC_215/A 0.06fF
C9897 AND2X1_LOC_511/a_8_24# AND2X1_LOC_31/Y 0.01fF
C9898 OR2X1_LOC_280/Y AND2X1_LOC_717/B 0.10fF
C9899 VDD OR2X1_LOC_406/A 0.21fF
C9900 OR2X1_LOC_74/A OR2X1_LOC_7/A 0.25fF
C9901 AND2X1_LOC_711/Y AND2X1_LOC_474/Y 0.03fF
C9902 OR2X1_LOC_663/A AND2X1_LOC_88/Y 0.03fF
C9903 AND2X1_LOC_95/Y AND2X1_LOC_431/a_8_24# 0.01fF
C9904 OR2X1_LOC_70/Y AND2X1_LOC_474/Y 0.14fF
C9905 OR2X1_LOC_633/A OR2X1_LOC_71/A 0.09fF
C9906 AND2X1_LOC_7/B OR2X1_LOC_515/Y 0.13fF
C9907 AND2X1_LOC_17/Y AND2X1_LOC_1/Y 0.02fF
C9908 VDD OR2X1_LOC_745/Y 0.12fF
C9909 OR2X1_LOC_473/Y OR2X1_LOC_810/A 0.01fF
C9910 D_INPUT_0 AND2X1_LOC_43/B 0.05fF
C9911 OR2X1_LOC_175/Y OR2X1_LOC_535/a_8_216# 0.05fF
C9912 AND2X1_LOC_465/a_36_24# OR2X1_LOC_485/A 0.00fF
C9913 OR2X1_LOC_158/A AND2X1_LOC_215/a_8_24# 0.01fF
C9914 OR2X1_LOC_654/A OR2X1_LOC_35/B 0.03fF
C9915 OR2X1_LOC_70/Y OR2X1_LOC_485/A 9.68fF
C9916 OR2X1_LOC_66/A OR2X1_LOC_398/Y 0.00fF
C9917 OR2X1_LOC_185/Y OR2X1_LOC_62/B 0.05fF
C9918 OR2X1_LOC_527/Y AND2X1_LOC_475/a_8_24# 0.01fF
C9919 VDD OR2X1_LOC_377/a_8_216# 0.21fF
C9920 AND2X1_LOC_169/a_8_24# AND2X1_LOC_436/B 0.03fF
C9921 OR2X1_LOC_316/Y AND2X1_LOC_831/Y 0.00fF
C9922 AND2X1_LOC_70/Y OR2X1_LOC_750/Y 0.15fF
C9923 OR2X1_LOC_744/A AND2X1_LOC_656/a_8_24# 0.01fF
C9924 AND2X1_LOC_612/B OR2X1_LOC_54/Y 0.01fF
C9925 OR2X1_LOC_161/B OR2X1_LOC_712/B 0.01fF
C9926 OR2X1_LOC_91/Y OR2X1_LOC_31/Y 0.03fF
C9927 AND2X1_LOC_259/Y OR2X1_LOC_54/Y 0.00fF
C9928 INPUT_1 OR2X1_LOC_753/A 0.01fF
C9929 AND2X1_LOC_512/a_8_24# OR2X1_LOC_22/Y 0.01fF
C9930 AND2X1_LOC_42/B OR2X1_LOC_121/B 0.04fF
C9931 OR2X1_LOC_295/a_8_216# OR2X1_LOC_258/Y 0.01fF
C9932 OR2X1_LOC_22/Y AND2X1_LOC_717/B 0.07fF
C9933 AND2X1_LOC_474/Y AND2X1_LOC_657/a_8_24# 0.00fF
C9934 AND2X1_LOC_538/a_8_24# OR2X1_LOC_485/A 0.02fF
C9935 OR2X1_LOC_80/a_8_216# OR2X1_LOC_26/Y 0.01fF
C9936 OR2X1_LOC_84/B OR2X1_LOC_244/A 0.01fF
C9937 OR2X1_LOC_62/B OR2X1_LOC_278/a_36_216# 0.03fF
C9938 OR2X1_LOC_355/B OR2X1_LOC_532/B 0.01fF
C9939 OR2X1_LOC_141/B OR2X1_LOC_244/A 0.18fF
C9940 OR2X1_LOC_862/B OR2X1_LOC_558/A 0.36fF
C9941 AND2X1_LOC_785/A OR2X1_LOC_373/Y 0.01fF
C9942 OR2X1_LOC_532/B OR2X1_LOC_733/B 0.01fF
C9943 AND2X1_LOC_12/Y OR2X1_LOC_770/Y 0.01fF
C9944 OR2X1_LOC_413/Y AND2X1_LOC_462/B 0.79fF
C9945 OR2X1_LOC_549/B OR2X1_LOC_577/Y 0.02fF
C9946 OR2X1_LOC_404/Y AND2X1_LOC_134/a_8_24# 0.01fF
C9947 AND2X1_LOC_157/a_8_24# OR2X1_LOC_451/B 0.01fF
C9948 OR2X1_LOC_600/A OR2X1_LOC_749/Y 0.46fF
C9949 AND2X1_LOC_647/a_8_24# OR2X1_LOC_71/A 0.05fF
C9950 OR2X1_LOC_154/A AND2X1_LOC_72/B 0.03fF
C9951 AND2X1_LOC_674/a_8_24# OR2X1_LOC_532/B 0.01fF
C9952 AND2X1_LOC_687/a_8_24# OR2X1_LOC_52/B 0.01fF
C9953 AND2X1_LOC_425/Y OR2X1_LOC_451/A 0.01fF
C9954 OR2X1_LOC_48/B OR2X1_LOC_172/a_8_216# 0.01fF
C9955 OR2X1_LOC_574/A OR2X1_LOC_473/A 0.15fF
C9956 AND2X1_LOC_59/Y OR2X1_LOC_358/A 1.10fF
C9957 OR2X1_LOC_527/Y OR2X1_LOC_31/Y 0.09fF
C9958 OR2X1_LOC_97/A AND2X1_LOC_60/a_8_24# 0.01fF
C9959 AND2X1_LOC_191/B AND2X1_LOC_789/Y 0.07fF
C9960 OR2X1_LOC_485/A OR2X1_LOC_184/Y 0.01fF
C9961 OR2X1_LOC_351/B OR2X1_LOC_333/a_36_216# 0.00fF
C9962 OR2X1_LOC_139/A OR2X1_LOC_161/B 0.22fF
C9963 OR2X1_LOC_70/Y AND2X1_LOC_452/a_8_24# 0.02fF
C9964 OR2X1_LOC_819/a_36_216# OR2X1_LOC_749/Y 0.00fF
C9965 OR2X1_LOC_417/Y OR2X1_LOC_31/Y 0.03fF
C9966 OR2X1_LOC_291/Y OR2X1_LOC_31/Y 0.06fF
C9967 AND2X1_LOC_11/a_8_24# AND2X1_LOC_25/a_8_24# 0.23fF
C9968 OR2X1_LOC_866/B D_GATE_662 0.14fF
C9969 OR2X1_LOC_518/a_8_216# AND2X1_LOC_326/B 0.01fF
C9970 AND2X1_LOC_7/B OR2X1_LOC_549/A 0.15fF
C9971 AND2X1_LOC_340/Y AND2X1_LOC_786/Y 2.01fF
C9972 OR2X1_LOC_130/A AND2X1_LOC_432/a_8_24# 0.03fF
C9973 OR2X1_LOC_144/a_8_216# OR2X1_LOC_51/Y 0.14fF
C9974 AND2X1_LOC_632/a_8_24# AND2X1_LOC_620/Y 0.01fF
C9975 OR2X1_LOC_691/Y OR2X1_LOC_856/A 0.01fF
C9976 OR2X1_LOC_619/Y AND2X1_LOC_212/a_8_24# 0.05fF
C9977 OR2X1_LOC_799/A OR2X1_LOC_446/B 0.09fF
C9978 OR2X1_LOC_151/A AND2X1_LOC_248/a_8_24# 0.01fF
C9979 OR2X1_LOC_696/A AND2X1_LOC_732/a_36_24# 0.01fF
C9980 OR2X1_LOC_659/Y OR2X1_LOC_663/a_8_216# 0.03fF
C9981 AND2X1_LOC_181/Y AND2X1_LOC_786/Y 0.07fF
C9982 OR2X1_LOC_160/B OR2X1_LOC_338/A 0.01fF
C9983 OR2X1_LOC_26/Y AND2X1_LOC_563/Y 0.02fF
C9984 AND2X1_LOC_181/Y OR2X1_LOC_323/a_8_216# 0.14fF
C9985 OR2X1_LOC_744/A AND2X1_LOC_780/a_8_24# 0.02fF
C9986 OR2X1_LOC_755/A AND2X1_LOC_793/Y 0.08fF
C9987 OR2X1_LOC_665/a_8_216# AND2X1_LOC_792/Y 0.01fF
C9988 AND2X1_LOC_624/A OR2X1_LOC_437/A 0.09fF
C9989 OR2X1_LOC_574/A OR2X1_LOC_228/Y 0.10fF
C9990 OR2X1_LOC_481/A AND2X1_LOC_848/A 0.03fF
C9991 OR2X1_LOC_89/A AND2X1_LOC_563/Y 0.04fF
C9992 AND2X1_LOC_810/A OR2X1_LOC_40/Y 0.06fF
C9993 OR2X1_LOC_375/A OR2X1_LOC_546/a_36_216# 0.00fF
C9994 OR2X1_LOC_147/B OR2X1_LOC_308/Y 0.10fF
C9995 AND2X1_LOC_477/Y AND2X1_LOC_220/a_8_24# 0.01fF
C9996 AND2X1_LOC_596/a_8_24# OR2X1_LOC_12/Y 0.18fF
C9997 OR2X1_LOC_356/A OR2X1_LOC_356/a_8_216# 0.17fF
C9998 OR2X1_LOC_602/a_8_216# AND2X1_LOC_31/Y -0.00fF
C9999 OR2X1_LOC_13/Y AND2X1_LOC_194/Y 0.01fF
C10000 AND2X1_LOC_91/B OR2X1_LOC_105/a_8_216# 0.01fF
C10001 OR2X1_LOC_436/Y OR2X1_LOC_112/B 0.02fF
C10002 OR2X1_LOC_161/A OR2X1_LOC_500/a_8_216# 0.48fF
C10003 OR2X1_LOC_813/A OR2X1_LOC_67/Y 0.01fF
C10004 AND2X1_LOC_359/B AND2X1_LOC_247/a_8_24# 0.03fF
C10005 OR2X1_LOC_6/B OR2X1_LOC_641/A 0.07fF
C10006 OR2X1_LOC_235/B OR2X1_LOC_266/A 0.06fF
C10007 OR2X1_LOC_64/Y AND2X1_LOC_790/a_8_24# 0.17fF
C10008 AND2X1_LOC_809/a_8_24# AND2X1_LOC_434/Y 0.01fF
C10009 OR2X1_LOC_781/B VDD -0.00fF
C10010 AND2X1_LOC_721/Y AND2X1_LOC_734/Y 0.01fF
C10011 OR2X1_LOC_154/A AND2X1_LOC_36/Y 2.56fF
C10012 OR2X1_LOC_45/B AND2X1_LOC_605/Y 0.02fF
C10013 OR2X1_LOC_16/A OR2X1_LOC_597/a_8_216# 0.01fF
C10014 VDD OR2X1_LOC_307/A 0.21fF
C10015 OR2X1_LOC_40/Y AND2X1_LOC_860/A 0.06fF
C10016 OR2X1_LOC_623/a_8_216# OR2X1_LOC_186/a_8_216# 0.47fF
C10017 AND2X1_LOC_529/a_8_24# OR2X1_LOC_548/B 0.00fF
C10018 OR2X1_LOC_329/Y VDD 0.17fF
C10019 OR2X1_LOC_673/A AND2X1_LOC_8/a_8_24# 0.19fF
C10020 OR2X1_LOC_40/Y OR2X1_LOC_626/Y 0.03fF
C10021 VDD AND2X1_LOC_606/a_8_24# 0.00fF
C10022 AND2X1_LOC_59/Y OR2X1_LOC_168/Y 0.02fF
C10023 OR2X1_LOC_2/a_36_216# INPUT_7 0.00fF
C10024 AND2X1_LOC_22/Y OR2X1_LOC_608/a_8_216# 0.03fF
C10025 OR2X1_LOC_589/A OR2X1_LOC_91/A 4.15fF
C10026 OR2X1_LOC_244/a_8_216# OR2X1_LOC_161/B 0.01fF
C10027 AND2X1_LOC_190/a_8_24# OR2X1_LOC_108/Y 0.01fF
C10028 OR2X1_LOC_139/A OR2X1_LOC_61/Y 0.07fF
C10029 OR2X1_LOC_96/Y OR2X1_LOC_51/Y 0.00fF
C10030 VDD OR2X1_LOC_411/A -0.00fF
C10031 OR2X1_LOC_160/A AND2X1_LOC_226/a_8_24# 0.03fF
C10032 AND2X1_LOC_326/B AND2X1_LOC_112/a_8_24# 0.01fF
C10033 OR2X1_LOC_666/a_8_216# AND2X1_LOC_658/A 0.01fF
C10034 OR2X1_LOC_479/Y OR2X1_LOC_777/B 0.07fF
C10035 OR2X1_LOC_44/Y OR2X1_LOC_387/A 0.02fF
C10036 AND2X1_LOC_12/Y OR2X1_LOC_334/a_8_216# 0.01fF
C10037 OR2X1_LOC_756/B AND2X1_LOC_524/a_8_24# 0.18fF
C10038 OR2X1_LOC_648/B OR2X1_LOC_78/B 0.35fF
C10039 OR2X1_LOC_833/B OR2X1_LOC_563/A 0.01fF
C10040 OR2X1_LOC_502/A AND2X1_LOC_433/a_8_24# 0.01fF
C10041 AND2X1_LOC_352/a_8_24# AND2X1_LOC_364/Y 0.01fF
C10042 AND2X1_LOC_352/a_36_24# OR2X1_LOC_329/B 0.01fF
C10043 AND2X1_LOC_508/B AND2X1_LOC_510/A 0.00fF
C10044 AND2X1_LOC_22/Y OR2X1_LOC_185/A 0.16fF
C10045 AND2X1_LOC_70/Y OR2X1_LOC_809/B 0.24fF
C10046 OR2X1_LOC_651/A OR2X1_LOC_197/a_8_216# 0.04fF
C10047 AND2X1_LOC_508/a_8_24# AND2X1_LOC_510/A 0.00fF
C10048 OR2X1_LOC_3/Y OR2X1_LOC_386/a_8_216# 0.02fF
C10049 AND2X1_LOC_334/Y AND2X1_LOC_338/a_36_24# 0.01fF
C10050 OR2X1_LOC_87/A OR2X1_LOC_718/a_36_216# 0.00fF
C10051 OR2X1_LOC_188/Y OR2X1_LOC_456/Y 0.00fF
C10052 OR2X1_LOC_631/B OR2X1_LOC_140/B 1.39fF
C10053 OR2X1_LOC_254/B OR2X1_LOC_563/A 0.15fF
C10054 AND2X1_LOC_853/Y OR2X1_LOC_171/a_8_216# 0.48fF
C10055 OR2X1_LOC_51/Y AND2X1_LOC_663/A 0.03fF
C10056 AND2X1_LOC_91/B AND2X1_LOC_56/B 0.16fF
C10057 OR2X1_LOC_231/B OR2X1_LOC_231/a_8_216# 0.47fF
C10058 AND2X1_LOC_337/a_8_24# OR2X1_LOC_91/A 0.05fF
C10059 OR2X1_LOC_124/B AND2X1_LOC_41/A 0.01fF
C10060 AND2X1_LOC_580/A AND2X1_LOC_580/a_8_24# 0.10fF
C10061 AND2X1_LOC_339/B AND2X1_LOC_649/B 0.01fF
C10062 AND2X1_LOC_861/a_8_24# AND2X1_LOC_865/A 0.01fF
C10063 OR2X1_LOC_778/A AND2X1_LOC_36/Y 0.01fF
C10064 OR2X1_LOC_756/B OR2X1_LOC_858/a_8_216# 0.02fF
C10065 OR2X1_LOC_691/Y OR2X1_LOC_793/a_36_216# 0.00fF
C10066 OR2X1_LOC_84/A OR2X1_LOC_398/Y 0.43fF
C10067 OR2X1_LOC_45/B AND2X1_LOC_318/a_8_24# 0.01fF
C10068 VDD OR2X1_LOC_292/Y 0.31fF
C10069 AND2X1_LOC_6/a_36_24# OR2X1_LOC_598/A 0.00fF
C10070 AND2X1_LOC_773/Y OR2X1_LOC_306/Y 0.00fF
C10071 OR2X1_LOC_154/a_8_216# OR2X1_LOC_154/A 0.04fF
C10072 AND2X1_LOC_91/B AND2X1_LOC_8/Y 0.28fF
C10073 AND2X1_LOC_51/Y OR2X1_LOC_703/Y 0.02fF
C10074 OR2X1_LOC_532/B OR2X1_LOC_366/Y 0.04fF
C10075 OR2X1_LOC_756/B OR2X1_LOC_648/A 0.07fF
C10076 OR2X1_LOC_624/A OR2X1_LOC_113/B 0.00fF
C10077 OR2X1_LOC_186/Y OR2X1_LOC_799/a_8_216# 0.01fF
C10078 OR2X1_LOC_179/a_8_216# OR2X1_LOC_56/A 0.01fF
C10079 OR2X1_LOC_741/Y OR2X1_LOC_190/B 0.12fF
C10080 AND2X1_LOC_72/Y OR2X1_LOC_719/B 1.05fF
C10081 AND2X1_LOC_70/Y AND2X1_LOC_177/a_36_24# 0.01fF
C10082 OR2X1_LOC_161/A OR2X1_LOC_596/A 0.03fF
C10083 OR2X1_LOC_8/Y AND2X1_LOC_839/a_8_24# 0.00fF
C10084 OR2X1_LOC_336/a_8_216# OR2X1_LOC_468/Y 0.01fF
C10085 OR2X1_LOC_45/B AND2X1_LOC_361/A 0.30fF
C10086 OR2X1_LOC_805/A OR2X1_LOC_549/A 0.07fF
C10087 OR2X1_LOC_362/B OR2X1_LOC_362/A 0.04fF
C10088 OR2X1_LOC_756/B OR2X1_LOC_410/a_8_216# 0.03fF
C10089 AND2X1_LOC_843/Y AND2X1_LOC_860/A 0.02fF
C10090 OR2X1_LOC_831/A AND2X1_LOC_43/B 0.03fF
C10091 OR2X1_LOC_337/A OR2X1_LOC_87/A 0.02fF
C10092 OR2X1_LOC_521/Y AND2X1_LOC_715/A 0.01fF
C10093 OR2X1_LOC_600/A OR2X1_LOC_427/A 0.36fF
C10094 OR2X1_LOC_91/A OR2X1_LOC_275/Y 0.03fF
C10095 OR2X1_LOC_36/Y OR2X1_LOC_12/Y 0.30fF
C10096 AND2X1_LOC_125/a_8_24# OR2X1_LOC_244/Y 0.01fF
C10097 AND2X1_LOC_486/Y AND2X1_LOC_570/Y 0.03fF
C10098 OR2X1_LOC_763/Y OR2X1_LOC_764/a_8_216# 0.39fF
C10099 OR2X1_LOC_479/Y OR2X1_LOC_831/B 0.02fF
C10100 OR2X1_LOC_448/A OR2X1_LOC_78/A 0.00fF
C10101 AND2X1_LOC_43/B OR2X1_LOC_515/A 0.01fF
C10102 OR2X1_LOC_51/Y OR2X1_LOC_2/Y 0.07fF
C10103 OR2X1_LOC_566/A OR2X1_LOC_479/Y 0.05fF
C10104 VDD OR2X1_LOC_560/a_8_216# 0.00fF
C10105 AND2X1_LOC_737/a_36_24# AND2X1_LOC_443/Y 0.00fF
C10106 AND2X1_LOC_347/B AND2X1_LOC_848/Y 0.04fF
C10107 AND2X1_LOC_765/a_8_24# OR2X1_LOC_287/B 0.00fF
C10108 AND2X1_LOC_575/a_36_24# AND2X1_LOC_191/Y 0.01fF
C10109 AND2X1_LOC_164/a_36_24# OR2X1_LOC_502/A 0.01fF
C10110 AND2X1_LOC_719/Y AND2X1_LOC_580/A 0.03fF
C10111 AND2X1_LOC_858/B OR2X1_LOC_495/Y 0.01fF
C10112 AND2X1_LOC_546/a_8_24# AND2X1_LOC_658/A 0.04fF
C10113 AND2X1_LOC_566/B OR2X1_LOC_6/A 0.03fF
C10114 OR2X1_LOC_189/Y AND2X1_LOC_213/B 0.05fF
C10115 OR2X1_LOC_773/B OR2X1_LOC_160/B 0.03fF
C10116 OR2X1_LOC_427/A AND2X1_LOC_296/a_8_24# 0.10fF
C10117 OR2X1_LOC_49/A OR2X1_LOC_89/A 0.07fF
C10118 AND2X1_LOC_387/a_36_24# OR2X1_LOC_161/A 0.00fF
C10119 OR2X1_LOC_568/A OR2X1_LOC_365/B 0.00fF
C10120 AND2X1_LOC_810/A OR2X1_LOC_7/A 0.03fF
C10121 AND2X1_LOC_99/A AND2X1_LOC_121/a_8_24# 0.01fF
C10122 AND2X1_LOC_22/Y OR2X1_LOC_435/Y 0.34fF
C10123 OR2X1_LOC_216/A OR2X1_LOC_474/Y 0.21fF
C10124 OR2X1_LOC_319/B OR2X1_LOC_354/A 0.21fF
C10125 OR2X1_LOC_160/A AND2X1_LOC_70/Y 0.22fF
C10126 OR2X1_LOC_578/B OR2X1_LOC_365/B 0.06fF
C10127 OR2X1_LOC_6/B AND2X1_LOC_404/a_8_24# 0.01fF
C10128 AND2X1_LOC_81/B OR2X1_LOC_160/B 0.03fF
C10129 OR2X1_LOC_6/B OR2X1_LOC_114/Y 0.03fF
C10130 OR2X1_LOC_51/Y AND2X1_LOC_449/Y 0.02fF
C10131 OR2X1_LOC_682/Y AND2X1_LOC_714/B 0.01fF
C10132 OR2X1_LOC_160/B OR2X1_LOC_358/B 0.09fF
C10133 AND2X1_LOC_3/Y AND2X1_LOC_65/A 0.35fF
C10134 OR2X1_LOC_89/A OR2X1_LOC_381/a_36_216# 0.00fF
C10135 OR2X1_LOC_448/A OR2X1_LOC_448/B 0.26fF
C10136 AND2X1_LOC_753/B OR2X1_LOC_502/A 0.03fF
C10137 OR2X1_LOC_744/A AND2X1_LOC_400/a_36_24# 0.00fF
C10138 AND2X1_LOC_592/Y AND2X1_LOC_645/A 0.00fF
C10139 D_GATE_662 OR2X1_LOC_557/A 0.04fF
C10140 VDD AND2X1_LOC_702/Y 0.28fF
C10141 OR2X1_LOC_241/Y OR2X1_LOC_776/A 0.01fF
C10142 OR2X1_LOC_759/A AND2X1_LOC_580/B 0.61fF
C10143 AND2X1_LOC_365/A OR2X1_LOC_91/A 0.29fF
C10144 AND2X1_LOC_86/a_36_24# AND2X1_LOC_8/Y 0.01fF
C10145 OR2X1_LOC_368/a_8_216# OR2X1_LOC_312/Y 0.01fF
C10146 OR2X1_LOC_526/Y OR2X1_LOC_26/Y 0.00fF
C10147 OR2X1_LOC_283/a_8_216# OR2X1_LOC_51/Y 0.01fF
C10148 OR2X1_LOC_756/Y OR2X1_LOC_555/B 0.07fF
C10149 OR2X1_LOC_680/A AND2X1_LOC_663/A 0.03fF
C10150 AND2X1_LOC_303/B OR2X1_LOC_56/A 0.21fF
C10151 OR2X1_LOC_854/a_8_216# OR2X1_LOC_856/B 0.01fF
C10152 OR2X1_LOC_389/A OR2X1_LOC_269/B 0.01fF
C10153 AND2X1_LOC_542/a_36_24# OR2X1_LOC_280/Y 0.02fF
C10154 OR2X1_LOC_461/a_8_216# OR2X1_LOC_461/A 0.47fF
C10155 AND2X1_LOC_541/Y OR2X1_LOC_529/Y 0.02fF
C10156 OR2X1_LOC_7/A AND2X1_LOC_254/a_8_24# 0.07fF
C10157 OR2X1_LOC_154/A OR2X1_LOC_630/Y 0.10fF
C10158 AND2X1_LOC_339/Y OR2X1_LOC_416/Y 0.01fF
C10159 OR2X1_LOC_808/A OR2X1_LOC_161/A 0.98fF
C10160 OR2X1_LOC_76/A AND2X1_LOC_604/a_36_24# 0.01fF
C10161 OR2X1_LOC_691/A AND2X1_LOC_689/a_36_24# 0.00fF
C10162 OR2X1_LOC_666/A AND2X1_LOC_859/Y 0.01fF
C10163 OR2X1_LOC_8/Y AND2X1_LOC_839/B 0.00fF
C10164 OR2X1_LOC_325/a_8_216# OR2X1_LOC_620/Y 0.02fF
C10165 OR2X1_LOC_282/Y AND2X1_LOC_285/a_8_24# 0.01fF
C10166 OR2X1_LOC_7/A AND2X1_LOC_860/A 0.07fF
C10167 OR2X1_LOC_375/A AND2X1_LOC_232/a_36_24# 0.01fF
C10168 OR2X1_LOC_405/A OR2X1_LOC_502/A 3.75fF
C10169 OR2X1_LOC_31/Y OR2X1_LOC_171/Y 0.17fF
C10170 AND2X1_LOC_6/a_8_24# AND2X1_LOC_36/Y 0.01fF
C10171 OR2X1_LOC_830/a_8_216# AND2X1_LOC_3/Y 0.01fF
C10172 OR2X1_LOC_643/A AND2X1_LOC_92/Y 0.02fF
C10173 OR2X1_LOC_526/Y OR2X1_LOC_89/A 0.03fF
C10174 AND2X1_LOC_658/B AND2X1_LOC_474/Y 0.03fF
C10175 AND2X1_LOC_707/a_36_24# OR2X1_LOC_52/B 0.01fF
C10176 OR2X1_LOC_744/A AND2X1_LOC_806/A 0.03fF
C10177 OR2X1_LOC_778/Y AND2X1_LOC_92/Y 0.25fF
C10178 AND2X1_LOC_51/Y OR2X1_LOC_596/A 0.14fF
C10179 OR2X1_LOC_245/a_8_216# OR2X1_LOC_595/A 0.05fF
C10180 VDD OR2X1_LOC_530/Y 0.16fF
C10181 AND2X1_LOC_489/Y OR2X1_LOC_494/Y 0.00fF
C10182 OR2X1_LOC_6/B OR2X1_LOC_825/a_8_216# 0.04fF
C10183 AND2X1_LOC_40/Y AND2X1_LOC_43/B 0.10fF
C10184 OR2X1_LOC_744/A OR2X1_LOC_83/A 0.27fF
C10185 OR2X1_LOC_43/A OR2X1_LOC_91/A 10.31fF
C10186 AND2X1_LOC_22/Y AND2X1_LOC_431/a_8_24# -0.00fF
C10187 OR2X1_LOC_185/Y OR2X1_LOC_571/a_8_216# 0.02fF
C10188 OR2X1_LOC_715/B OR2X1_LOC_473/Y 0.03fF
C10189 AND2X1_LOC_516/a_8_24# OR2X1_LOC_715/A 0.27fF
C10190 OR2X1_LOC_427/A OR2X1_LOC_619/Y 0.03fF
C10191 AND2X1_LOC_848/A AND2X1_LOC_789/Y 0.21fF
C10192 OR2X1_LOC_497/Y AND2X1_LOC_850/A 0.01fF
C10193 AND2X1_LOC_398/a_8_24# AND2X1_LOC_573/A 0.01fF
C10194 OR2X1_LOC_382/Y AND2X1_LOC_818/a_8_24# 0.01fF
C10195 OR2X1_LOC_671/Y OR2X1_LOC_54/Y 0.01fF
C10196 VDD OR2X1_LOC_35/B 0.00fF
C10197 OR2X1_LOC_129/a_8_216# OR2X1_LOC_291/Y 0.02fF
C10198 OR2X1_LOC_532/B OR2X1_LOC_548/B 0.00fF
C10199 OR2X1_LOC_797/A OR2X1_LOC_160/Y 0.01fF
C10200 OR2X1_LOC_531/Y OR2X1_LOC_74/A 0.01fF
C10201 OR2X1_LOC_475/a_8_216# OR2X1_LOC_87/A 0.05fF
C10202 OR2X1_LOC_185/A OR2X1_LOC_664/a_8_216# 0.02fF
C10203 AND2X1_LOC_76/a_8_24# OR2X1_LOC_265/Y 0.02fF
C10204 OR2X1_LOC_634/A OR2X1_LOC_240/A 0.12fF
C10205 AND2X1_LOC_12/Y OR2X1_LOC_231/a_8_216# 0.01fF
C10206 OR2X1_LOC_777/B OR2X1_LOC_68/B 0.03fF
C10207 AND2X1_LOC_380/a_8_24# OR2X1_LOC_160/A 0.03fF
C10208 OR2X1_LOC_533/A OR2X1_LOC_13/B 0.02fF
C10209 AND2X1_LOC_490/a_8_24# OR2X1_LOC_78/Y 0.24fF
C10210 AND2X1_LOC_512/Y AND2X1_LOC_645/A 0.62fF
C10211 AND2X1_LOC_34/Y OR2X1_LOC_18/Y 0.00fF
C10212 OR2X1_LOC_391/B OR2X1_LOC_772/B 0.29fF
C10213 OR2X1_LOC_185/A AND2X1_LOC_153/a_8_24# 0.01fF
C10214 AND2X1_LOC_56/B AND2X1_LOC_39/a_36_24# 0.00fF
C10215 AND2X1_LOC_86/Y AND2X1_LOC_81/B 0.02fF
C10216 AND2X1_LOC_592/Y AND2X1_LOC_477/A 0.03fF
C10217 OR2X1_LOC_630/Y OR2X1_LOC_778/A 0.01fF
C10218 OR2X1_LOC_64/Y AND2X1_LOC_436/Y 0.06fF
C10219 AND2X1_LOC_47/Y OR2X1_LOC_294/Y 0.01fF
C10220 OR2X1_LOC_160/B OR2X1_LOC_196/B 0.07fF
C10221 AND2X1_LOC_422/a_8_24# OR2X1_LOC_269/B 0.01fF
C10222 OR2X1_LOC_808/B OR2X1_LOC_787/Y 0.10fF
C10223 AND2X1_LOC_474/A OR2X1_LOC_279/Y 0.01fF
C10224 OR2X1_LOC_47/Y AND2X1_LOC_636/a_8_24# 0.01fF
C10225 OR2X1_LOC_316/Y AND2X1_LOC_139/B 0.03fF
C10226 AND2X1_LOC_36/Y OR2X1_LOC_198/A 0.02fF
C10227 OR2X1_LOC_424/Y OR2X1_LOC_423/Y 0.61fF
C10228 OR2X1_LOC_154/A OR2X1_LOC_447/a_36_216# 0.00fF
C10229 AND2X1_LOC_56/B AND2X1_LOC_72/Y 0.00fF
C10230 OR2X1_LOC_127/a_8_216# OR2X1_LOC_6/A 0.01fF
C10231 AND2X1_LOC_580/A OR2X1_LOC_252/Y 0.03fF
C10232 OR2X1_LOC_599/A OR2X1_LOC_432/Y 0.00fF
C10233 OR2X1_LOC_865/B OR2X1_LOC_269/B 0.03fF
C10234 OR2X1_LOC_160/B AND2X1_LOC_692/a_8_24# 0.05fF
C10235 OR2X1_LOC_19/B AND2X1_LOC_403/a_36_24# 0.01fF
C10236 AND2X1_LOC_155/a_8_24# OR2X1_LOC_7/A -0.00fF
C10237 OR2X1_LOC_656/B OR2X1_LOC_218/a_8_216# 0.02fF
C10238 AND2X1_LOC_535/Y OR2X1_LOC_167/Y 0.02fF
C10239 AND2X1_LOC_572/Y OR2X1_LOC_44/Y 0.03fF
C10240 OR2X1_LOC_91/A AND2X1_LOC_685/a_8_24# 0.01fF
C10241 OR2X1_LOC_475/a_8_216# OR2X1_LOC_216/a_8_216# 0.47fF
C10242 OR2X1_LOC_861/a_36_216# OR2X1_LOC_287/B 0.00fF
C10243 OR2X1_LOC_391/B OR2X1_LOC_489/B 0.03fF
C10244 OR2X1_LOC_43/A AND2X1_LOC_573/A 0.07fF
C10245 OR2X1_LOC_462/a_36_216# INPUT_0 0.01fF
C10246 OR2X1_LOC_318/a_36_216# OR2X1_LOC_223/A 0.00fF
C10247 AND2X1_LOC_662/a_8_24# OR2X1_LOC_275/Y 0.01fF
C10248 OR2X1_LOC_51/Y OR2X1_LOC_7/Y 0.16fF
C10249 OR2X1_LOC_45/B AND2X1_LOC_795/Y 0.00fF
C10250 OR2X1_LOC_83/Y AND2X1_LOC_403/B 0.81fF
C10251 OR2X1_LOC_11/Y OR2X1_LOC_588/Y 0.01fF
C10252 OR2X1_LOC_663/A OR2X1_LOC_121/B 0.03fF
C10253 OR2X1_LOC_96/B OR2X1_LOC_44/Y 0.04fF
C10254 OR2X1_LOC_48/Y OR2X1_LOC_48/B 0.28fF
C10255 AND2X1_LOC_811/a_8_24# OR2X1_LOC_52/B 0.17fF
C10256 OR2X1_LOC_467/A OR2X1_LOC_454/a_8_216# 0.01fF
C10257 OR2X1_LOC_652/a_36_216# OR2X1_LOC_810/A 0.02fF
C10258 INPUT_1 AND2X1_LOC_222/a_8_24# 0.01fF
C10259 OR2X1_LOC_121/Y OR2X1_LOC_66/a_8_216# 0.02fF
C10260 D_INPUT_0 AND2X1_LOC_219/Y 0.07fF
C10261 OR2X1_LOC_364/A OR2X1_LOC_449/B 0.01fF
C10262 OR2X1_LOC_497/a_36_216# OR2X1_LOC_497/Y 0.01fF
C10263 AND2X1_LOC_717/B OR2X1_LOC_39/A 0.07fF
C10264 OR2X1_LOC_831/B OR2X1_LOC_68/B 0.03fF
C10265 AND2X1_LOC_604/a_8_24# OR2X1_LOC_318/B 0.01fF
C10266 OR2X1_LOC_419/Y OR2X1_LOC_12/Y 0.00fF
C10267 OR2X1_LOC_158/A AND2X1_LOC_721/A 0.00fF
C10268 OR2X1_LOC_219/B OR2X1_LOC_358/B 0.01fF
C10269 AND2X1_LOC_512/Y AND2X1_LOC_477/A 0.07fF
C10270 AND2X1_LOC_520/a_36_24# AND2X1_LOC_222/Y 0.00fF
C10271 OR2X1_LOC_772/B OR2X1_LOC_772/Y 0.73fF
C10272 AND2X1_LOC_390/B AND2X1_LOC_436/B 0.46fF
C10273 OR2X1_LOC_83/Y OR2X1_LOC_44/Y 0.02fF
C10274 OR2X1_LOC_53/Y OR2X1_LOC_172/Y 0.09fF
C10275 OR2X1_LOC_770/A OR2X1_LOC_68/B 0.00fF
C10276 AND2X1_LOC_51/Y OR2X1_LOC_732/a_8_216# 0.14fF
C10277 AND2X1_LOC_97/a_8_24# OR2X1_LOC_64/Y 0.26fF
C10278 OR2X1_LOC_26/Y AND2X1_LOC_654/a_8_24# 0.02fF
C10279 OR2X1_LOC_844/Y OR2X1_LOC_523/Y 0.01fF
C10280 OR2X1_LOC_639/B OR2X1_LOC_636/B 0.06fF
C10281 OR2X1_LOC_160/A OR2X1_LOC_206/a_8_216# 0.01fF
C10282 AND2X1_LOC_753/B AND2X1_LOC_48/A 0.15fF
C10283 AND2X1_LOC_64/Y OR2X1_LOC_71/A 0.08fF
C10284 OR2X1_LOC_696/A AND2X1_LOC_592/a_36_24# 0.01fF
C10285 OR2X1_LOC_517/A AND2X1_LOC_845/Y 0.17fF
C10286 AND2X1_LOC_606/a_8_24# OR2X1_LOC_67/Y 0.04fF
C10287 AND2X1_LOC_663/B AND2X1_LOC_621/Y 0.01fF
C10288 AND2X1_LOC_64/Y AND2X1_LOC_419/a_36_24# -0.00fF
C10289 OR2X1_LOC_123/B OR2X1_LOC_375/A 0.02fF
C10290 AND2X1_LOC_95/Y OR2X1_LOC_476/B 0.03fF
C10291 OR2X1_LOC_609/A AND2X1_LOC_610/a_8_24# 0.01fF
C10292 AND2X1_LOC_76/Y AND2X1_LOC_116/B 0.01fF
C10293 OR2X1_LOC_272/Y OR2X1_LOC_36/Y 0.02fF
C10294 OR2X1_LOC_405/A AND2X1_LOC_48/A 0.22fF
C10295 VDD OR2X1_LOC_804/A 0.30fF
C10296 OR2X1_LOC_641/A OR2X1_LOC_598/A 0.07fF
C10297 OR2X1_LOC_489/B OR2X1_LOC_772/Y 0.12fF
C10298 OR2X1_LOC_12/Y OR2X1_LOC_526/a_8_216# 0.08fF
C10299 AND2X1_LOC_59/Y OR2X1_LOC_520/B 0.01fF
C10300 AND2X1_LOC_707/Y OR2X1_LOC_423/Y 0.03fF
C10301 OR2X1_LOC_446/a_8_216# OR2X1_LOC_155/A 0.05fF
C10302 OR2X1_LOC_22/Y AND2X1_LOC_452/Y 0.00fF
C10303 OR2X1_LOC_364/A OR2X1_LOC_121/B 0.07fF
C10304 OR2X1_LOC_497/Y AND2X1_LOC_523/Y 0.19fF
C10305 OR2X1_LOC_185/Y OR2X1_LOC_121/B 0.09fF
C10306 VDD OR2X1_LOC_723/A -0.00fF
C10307 OR2X1_LOC_635/A AND2X1_LOC_684/a_8_24# 0.04fF
C10308 OR2X1_LOC_516/A AND2X1_LOC_477/A 0.31fF
C10309 AND2X1_LOC_81/B OR2X1_LOC_647/a_36_216# 0.00fF
C10310 OR2X1_LOC_428/A OR2X1_LOC_589/a_8_216# 0.04fF
C10311 OR2X1_LOC_64/Y OR2X1_LOC_588/Y 0.26fF
C10312 OR2X1_LOC_175/Y OR2X1_LOC_537/a_8_216# 0.01fF
C10313 OR2X1_LOC_624/A OR2X1_LOC_532/B 0.33fF
C10314 OR2X1_LOC_3/Y AND2X1_LOC_345/Y 0.11fF
C10315 OR2X1_LOC_18/Y AND2X1_LOC_656/Y 0.01fF
C10316 OR2X1_LOC_296/Y OR2X1_LOC_629/a_8_216# 0.01fF
C10317 AND2X1_LOC_98/Y AND2X1_LOC_721/A 0.02fF
C10318 OR2X1_LOC_510/Y D_INPUT_0 0.07fF
C10319 OR2X1_LOC_744/A AND2X1_LOC_486/a_8_24# 0.01fF
C10320 OR2X1_LOC_502/A AND2X1_LOC_8/a_8_24# 0.03fF
C10321 OR2X1_LOC_617/a_36_216# OR2X1_LOC_617/Y 0.00fF
C10322 AND2X1_LOC_720/Y AND2X1_LOC_721/A 0.11fF
C10323 AND2X1_LOC_318/Y AND2X1_LOC_662/B 0.03fF
C10324 OR2X1_LOC_287/B OR2X1_LOC_401/a_8_216# 0.01fF
C10325 OR2X1_LOC_502/A OR2X1_LOC_330/a_8_216# 0.02fF
C10326 AND2X1_LOC_51/Y OR2X1_LOC_33/B 0.03fF
C10327 OR2X1_LOC_126/a_8_216# OR2X1_LOC_278/A 0.40fF
C10328 OR2X1_LOC_624/B OR2X1_LOC_404/Y 0.03fF
C10329 OR2X1_LOC_95/Y OR2X1_LOC_67/a_8_216# 0.04fF
C10330 AND2X1_LOC_86/a_8_24# OR2X1_LOC_71/A 0.01fF
C10331 OR2X1_LOC_616/a_8_216# GATE_662 0.01fF
C10332 AND2X1_LOC_387/B OR2X1_LOC_19/B 0.07fF
C10333 OR2X1_LOC_45/B OR2X1_LOC_395/a_8_216# 0.01fF
C10334 OR2X1_LOC_400/B OR2X1_LOC_532/B 0.03fF
C10335 OR2X1_LOC_599/A AND2X1_LOC_800/a_36_24# 0.00fF
C10336 OR2X1_LOC_810/A D_INPUT_0 0.10fF
C10337 OR2X1_LOC_216/Y OR2X1_LOC_218/Y 0.03fF
C10338 INPUT_1 OR2X1_LOC_37/a_8_216# 0.01fF
C10339 OR2X1_LOC_364/B OR2X1_LOC_212/B 0.01fF
C10340 AND2X1_LOC_76/Y AND2X1_LOC_204/Y 0.03fF
C10341 AND2X1_LOC_523/Y AND2X1_LOC_844/a_8_24# 0.09fF
C10342 OR2X1_LOC_85/a_36_216# OR2X1_LOC_278/Y 0.00fF
C10343 OR2X1_LOC_64/a_8_216# OR2X1_LOC_588/Y 0.01fF
C10344 OR2X1_LOC_91/A OR2X1_LOC_384/a_8_216# 0.06fF
C10345 OR2X1_LOC_26/Y AND2X1_LOC_810/Y 0.07fF
C10346 OR2X1_LOC_95/Y AND2X1_LOC_458/a_8_24# 0.04fF
C10347 AND2X1_LOC_798/a_8_24# OR2X1_LOC_428/A 0.05fF
C10348 AND2X1_LOC_79/a_8_24# AND2X1_LOC_51/Y 0.01fF
C10349 OR2X1_LOC_473/A OR2X1_LOC_203/Y 0.20fF
C10350 AND2X1_LOC_58/a_8_24# OR2X1_LOC_228/Y 0.17fF
C10351 AND2X1_LOC_12/Y OR2X1_LOC_194/a_36_216# 0.00fF
C10352 OR2X1_LOC_379/Y OR2X1_LOC_598/A 0.39fF
C10353 OR2X1_LOC_574/A OR2X1_LOC_436/Y 0.03fF
C10354 OR2X1_LOC_161/A OR2X1_LOC_374/Y 0.05fF
C10355 OR2X1_LOC_696/a_8_216# OR2X1_LOC_31/Y 0.01fF
C10356 AND2X1_LOC_810/Y OR2X1_LOC_89/A 0.15fF
C10357 OR2X1_LOC_217/Y OR2X1_LOC_205/Y 0.03fF
C10358 AND2X1_LOC_841/B AND2X1_LOC_222/Y 0.03fF
C10359 AND2X1_LOC_18/Y OR2X1_LOC_523/A 0.04fF
C10360 OR2X1_LOC_359/A OR2X1_LOC_580/A 0.05fF
C10361 OR2X1_LOC_575/A OR2X1_LOC_68/B 1.46fF
C10362 OR2X1_LOC_12/Y AND2X1_LOC_590/a_36_24# 0.00fF
C10363 AND2X1_LOC_337/B AND2X1_LOC_318/Y 0.19fF
C10364 AND2X1_LOC_70/Y OR2X1_LOC_532/Y 0.09fF
C10365 OR2X1_LOC_656/B OR2X1_LOC_559/a_8_216# 0.03fF
C10366 AND2X1_LOC_712/B AND2X1_LOC_477/A 0.01fF
C10367 OR2X1_LOC_597/a_36_216# OR2X1_LOC_13/B 0.03fF
C10368 AND2X1_LOC_40/Y OR2X1_LOC_357/A 0.02fF
C10369 OR2X1_LOC_220/B OR2X1_LOC_742/B 0.03fF
C10370 AND2X1_LOC_564/B AND2X1_LOC_786/Y 0.02fF
C10371 OR2X1_LOC_234/a_8_216# OR2X1_LOC_585/A 0.01fF
C10372 VDD AND2X1_LOC_792/B 0.01fF
C10373 OR2X1_LOC_308/A OR2X1_LOC_713/A 0.01fF
C10374 OR2X1_LOC_735/a_8_216# OR2X1_LOC_735/B 0.39fF
C10375 OR2X1_LOC_485/A OR2X1_LOC_47/Y 5.49fF
C10376 OR2X1_LOC_74/A OR2X1_LOC_615/Y 0.03fF
C10377 OR2X1_LOC_839/a_8_216# OR2X1_LOC_19/B 0.02fF
C10378 OR2X1_LOC_377/A OR2X1_LOC_228/Y 0.26fF
C10379 OR2X1_LOC_22/Y OR2X1_LOC_412/a_8_216# 0.04fF
C10380 OR2X1_LOC_105/Y OR2X1_LOC_579/a_8_216# 0.40fF
C10381 AND2X1_LOC_227/Y AND2X1_LOC_842/B 0.29fF
C10382 AND2X1_LOC_404/a_8_24# OR2X1_LOC_598/A 0.17fF
C10383 OR2X1_LOC_114/Y OR2X1_LOC_598/A 0.00fF
C10384 OR2X1_LOC_844/Y AND2X1_LOC_47/Y 0.03fF
C10385 OR2X1_LOC_269/B OR2X1_LOC_493/Y 0.01fF
C10386 OR2X1_LOC_532/B OR2X1_LOC_54/Y 0.07fF
C10387 OR2X1_LOC_52/B AND2X1_LOC_204/Y 0.03fF
C10388 OR2X1_LOC_269/B OR2X1_LOC_801/B 0.07fF
C10389 AND2X1_LOC_576/a_8_24# AND2X1_LOC_563/Y 0.01fF
C10390 AND2X1_LOC_437/a_8_24# OR2X1_LOC_180/B 0.01fF
C10391 OR2X1_LOC_329/B OR2X1_LOC_268/Y 0.03fF
C10392 OR2X1_LOC_52/B AND2X1_LOC_228/a_8_24# 0.04fF
C10393 AND2X1_LOC_841/B OR2X1_LOC_423/Y 0.15fF
C10394 AND2X1_LOC_832/a_8_24# OR2X1_LOC_589/Y 0.24fF
C10395 OR2X1_LOC_86/a_8_216# AND2X1_LOC_647/Y 0.01fF
C10396 OR2X1_LOC_631/B OR2X1_LOC_675/Y 0.02fF
C10397 OR2X1_LOC_703/A OR2X1_LOC_532/Y 0.00fF
C10398 OR2X1_LOC_520/Y AND2X1_LOC_31/Y 0.01fF
C10399 OR2X1_LOC_685/B AND2X1_LOC_430/B 0.00fF
C10400 OR2X1_LOC_419/Y OR2X1_LOC_239/a_8_216# 0.01fF
C10401 AND2X1_LOC_70/Y OR2X1_LOC_130/Y 0.00fF
C10402 AND2X1_LOC_348/A OR2X1_LOC_13/B 0.00fF
C10403 AND2X1_LOC_537/Y OR2X1_LOC_95/Y 0.01fF
C10404 OR2X1_LOC_825/Y OR2X1_LOC_826/Y 0.21fF
C10405 OR2X1_LOC_703/A OR2X1_LOC_212/B 0.00fF
C10406 AND2X1_LOC_7/Y OR2X1_LOC_228/a_8_216# 0.07fF
C10407 OR2X1_LOC_528/Y OR2X1_LOC_406/Y 0.01fF
C10408 OR2X1_LOC_696/A OR2X1_LOC_59/Y 0.04fF
C10409 AND2X1_LOC_649/B OR2X1_LOC_300/Y 0.01fF
C10410 OR2X1_LOC_840/A OR2X1_LOC_593/B 0.01fF
C10411 OR2X1_LOC_580/B OR2X1_LOC_549/A -0.00fF
C10412 OR2X1_LOC_485/A AND2X1_LOC_486/a_36_24# 0.00fF
C10413 OR2X1_LOC_691/Y OR2X1_LOC_644/a_36_216# 0.00fF
C10414 OR2X1_LOC_175/B OR2X1_LOC_174/Y 0.04fF
C10415 OR2X1_LOC_449/B OR2X1_LOC_568/A 0.55fF
C10416 AND2X1_LOC_64/Y OR2X1_LOC_858/A 0.04fF
C10417 AND2X1_LOC_831/Y OR2X1_LOC_31/Y 0.15fF
C10418 OR2X1_LOC_293/a_8_216# D_INPUT_1 0.10fF
C10419 OR2X1_LOC_62/A INPUT_1 2.58fF
C10420 OR2X1_LOC_7/A AND2X1_LOC_562/Y 0.12fF
C10421 OR2X1_LOC_743/A OR2X1_LOC_761/a_36_216# 0.00fF
C10422 AND2X1_LOC_91/B AND2X1_LOC_92/Y 0.20fF
C10423 AND2X1_LOC_539/Y AND2X1_LOC_434/Y 0.04fF
C10424 OR2X1_LOC_739/A OR2X1_LOC_532/a_8_216# 0.01fF
C10425 OR2X1_LOC_176/Y AND2X1_LOC_568/B 0.03fF
C10426 AND2X1_LOC_51/Y OR2X1_LOC_374/Y 0.01fF
C10427 AND2X1_LOC_191/B OR2X1_LOC_187/Y 0.01fF
C10428 OR2X1_LOC_64/Y OR2X1_LOC_86/A 0.10fF
C10429 OR2X1_LOC_620/Y OR2X1_LOC_469/B 0.03fF
C10430 AND2X1_LOC_56/B OR2X1_LOC_446/B 0.07fF
C10431 OR2X1_LOC_45/B AND2X1_LOC_61/Y 0.12fF
C10432 AND2X1_LOC_137/a_8_24# OR2X1_LOC_95/Y 0.08fF
C10433 OR2X1_LOC_604/A OR2X1_LOC_12/Y 0.21fF
C10434 OR2X1_LOC_486/Y OR2X1_LOC_182/B 0.03fF
C10435 OR2X1_LOC_615/a_8_216# OR2X1_LOC_753/Y 0.40fF
C10436 AND2X1_LOC_219/a_8_24# AND2X1_LOC_219/A 0.07fF
C10437 AND2X1_LOC_831/Y AND2X1_LOC_655/a_36_24# 0.00fF
C10438 AND2X1_LOC_334/Y AND2X1_LOC_219/A 0.17fF
C10439 OR2X1_LOC_35/Y AND2X1_LOC_44/Y 0.05fF
C10440 OR2X1_LOC_753/A OR2X1_LOC_150/a_8_216# 0.04fF
C10441 AND2X1_LOC_706/Y AND2X1_LOC_732/B 0.09fF
C10442 AND2X1_LOC_56/B OR2X1_LOC_728/a_8_216# 0.03fF
C10443 AND2X1_LOC_325/a_8_24# OR2X1_LOC_323/Y 0.07fF
C10444 AND2X1_LOC_568/B AND2X1_LOC_212/Y 0.01fF
C10445 OR2X1_LOC_840/A AND2X1_LOC_273/a_8_24# 0.14fF
C10446 AND2X1_LOC_122/a_8_24# OR2X1_LOC_560/A 0.01fF
C10447 AND2X1_LOC_47/Y AND2X1_LOC_813/a_36_24# 0.00fF
C10448 OR2X1_LOC_857/B OR2X1_LOC_66/A 0.04fF
C10449 OR2X1_LOC_574/a_36_216# OR2X1_LOC_140/B 0.00fF
C10450 OR2X1_LOC_523/B VDD -0.00fF
C10451 AND2X1_LOC_41/A OR2X1_LOC_779/A 0.03fF
C10452 AND2X1_LOC_12/Y OR2X1_LOC_308/Y 0.01fF
C10453 OR2X1_LOC_803/A OR2X1_LOC_160/Y 0.01fF
C10454 AND2X1_LOC_789/a_8_24# OR2X1_LOC_748/Y 0.23fF
C10455 OR2X1_LOC_155/A OR2X1_LOC_515/a_8_216# -0.02fF
C10456 AND2X1_LOC_456/B AND2X1_LOC_456/a_8_24# 0.11fF
C10457 OR2X1_LOC_797/B VDD 0.19fF
C10458 OR2X1_LOC_428/Y OR2X1_LOC_430/Y 0.19fF
C10459 OR2X1_LOC_47/Y OR2X1_LOC_10/a_8_216# 0.00fF
C10460 AND2X1_LOC_40/Y AND2X1_LOC_258/a_36_24# 0.01fF
C10461 AND2X1_LOC_47/Y OR2X1_LOC_544/a_8_216# 0.01fF
C10462 OR2X1_LOC_121/B OR2X1_LOC_578/B 0.03fF
C10463 OR2X1_LOC_160/B AND2X1_LOC_387/a_8_24# 0.01fF
C10464 OR2X1_LOC_47/Y OR2X1_LOC_609/Y 0.06fF
C10465 OR2X1_LOC_676/Y AND2X1_LOC_18/Y 0.07fF
C10466 AND2X1_LOC_727/A AND2X1_LOC_796/A 0.00fF
C10467 OR2X1_LOC_18/Y AND2X1_LOC_772/Y 0.08fF
C10468 AND2X1_LOC_462/B AND2X1_LOC_293/a_36_24# 0.01fF
C10469 AND2X1_LOC_232/a_36_24# OR2X1_LOC_549/A 0.00fF
C10470 AND2X1_LOC_141/A OR2X1_LOC_595/A 0.00fF
C10471 AND2X1_LOC_566/B AND2X1_LOC_514/a_36_24# 0.00fF
C10472 AND2X1_LOC_91/B AND2X1_LOC_166/a_8_24# 0.05fF
C10473 OR2X1_LOC_6/B OR2X1_LOC_744/A 0.19fF
C10474 AND2X1_LOC_753/B OR2X1_LOC_207/B 0.18fF
C10475 OR2X1_LOC_158/A AND2X1_LOC_605/Y 0.05fF
C10476 OR2X1_LOC_392/B OR2X1_LOC_161/A 0.03fF
C10477 OR2X1_LOC_808/B OR2X1_LOC_439/B 0.53fF
C10478 OR2X1_LOC_696/A OR2X1_LOC_820/B 0.04fF
C10479 AND2X1_LOC_806/a_36_24# OR2X1_LOC_56/A 0.00fF
C10480 OR2X1_LOC_421/A OR2X1_LOC_421/a_8_216# 0.18fF
C10481 OR2X1_LOC_309/Y AND2X1_LOC_335/a_8_24# 0.23fF
C10482 OR2X1_LOC_645/a_8_216# AND2X1_LOC_92/Y 0.05fF
C10483 OR2X1_LOC_158/A AND2X1_LOC_198/a_36_24# 0.01fF
C10484 OR2X1_LOC_51/Y OR2X1_LOC_25/Y 0.07fF
C10485 AND2X1_LOC_675/Y OR2X1_LOC_51/Y 0.01fF
C10486 OR2X1_LOC_709/A OR2X1_LOC_447/A 0.02fF
C10487 AND2X1_LOC_284/a_8_24# OR2X1_LOC_44/Y 0.01fF
C10488 OR2X1_LOC_757/A AND2X1_LOC_663/A 0.03fF
C10489 AND2X1_LOC_477/Y AND2X1_LOC_804/Y 0.01fF
C10490 AND2X1_LOC_865/a_8_24# AND2X1_LOC_807/B 0.09fF
C10491 OR2X1_LOC_762/a_36_216# D_INPUT_6 0.01fF
C10492 OR2X1_LOC_116/a_36_216# OR2X1_LOC_392/B 0.14fF
C10493 AND2X1_LOC_22/Y AND2X1_LOC_669/a_36_24# 0.01fF
C10494 OR2X1_LOC_306/Y OR2X1_LOC_12/Y 0.05fF
C10495 AND2X1_LOC_110/Y OR2X1_LOC_147/B 0.03fF
C10496 AND2X1_LOC_787/A OR2X1_LOC_44/Y 0.03fF
C10497 AND2X1_LOC_572/a_36_24# AND2X1_LOC_361/A 0.01fF
C10498 OR2X1_LOC_516/B OR2X1_LOC_51/Y 0.01fF
C10499 OR2X1_LOC_340/a_8_216# OR2X1_LOC_560/A 0.39fF
C10500 OR2X1_LOC_696/A OR2X1_LOC_70/Y 0.05fF
C10501 AND2X1_LOC_737/a_8_24# AND2X1_LOC_658/A 0.04fF
C10502 AND2X1_LOC_51/Y OR2X1_LOC_333/A 0.05fF
C10503 VDD OR2X1_LOC_403/A -0.00fF
C10504 OR2X1_LOC_6/A OR2X1_LOC_414/Y 0.00fF
C10505 OR2X1_LOC_755/a_8_216# OR2X1_LOC_755/Y -0.00fF
C10506 AND2X1_LOC_57/a_8_24# OR2X1_LOC_66/A 0.02fF
C10507 OR2X1_LOC_80/Y OR2X1_LOC_12/Y 0.00fF
C10508 OR2X1_LOC_589/A OR2X1_LOC_32/B 0.21fF
C10509 OR2X1_LOC_585/A OR2X1_LOC_312/a_8_216# 0.01fF
C10510 OR2X1_LOC_101/a_8_216# VDD 0.21fF
C10511 OR2X1_LOC_45/B AND2X1_LOC_852/Y 0.22fF
C10512 OR2X1_LOC_3/Y OR2X1_LOC_56/a_8_216# 0.01fF
C10513 AND2X1_LOC_456/Y AND2X1_LOC_242/B 0.02fF
C10514 VDD OR2X1_LOC_231/A 0.21fF
C10515 AND2X1_LOC_456/B AND2X1_LOC_474/A 0.02fF
C10516 OR2X1_LOC_6/B OR2X1_LOC_541/B 0.01fF
C10517 OR2X1_LOC_160/A OR2X1_LOC_362/A 0.15fF
C10518 OR2X1_LOC_471/Y OR2X1_LOC_209/A 0.09fF
C10519 OR2X1_LOC_107/a_36_216# OR2X1_LOC_103/Y 0.00fF
C10520 AND2X1_LOC_265/a_8_24# OR2X1_LOC_340/Y 0.00fF
C10521 OR2X1_LOC_6/B AND2X1_LOC_617/a_8_24# 0.17fF
C10522 OR2X1_LOC_693/a_8_216# OR2X1_LOC_44/Y 0.00fF
C10523 OR2X1_LOC_756/Y OR2X1_LOC_756/B 0.02fF
C10524 AND2X1_LOC_564/B AND2X1_LOC_578/A 0.07fF
C10525 OR2X1_LOC_696/A AND2X1_LOC_514/Y 0.07fF
C10526 OR2X1_LOC_631/B OR2X1_LOC_736/Y 0.19fF
C10527 OR2X1_LOC_329/B AND2X1_LOC_840/a_8_24# 0.01fF
C10528 OR2X1_LOC_808/B AND2X1_LOC_41/A 0.07fF
C10529 OR2X1_LOC_113/a_8_216# OR2X1_LOC_844/a_8_216# 0.47fF
C10530 VDD OR2X1_LOC_447/a_8_216# 0.21fF
C10531 AND2X1_LOC_131/a_8_24# OR2X1_LOC_510/Y 0.01fF
C10532 AND2X1_LOC_715/Y OR2X1_LOC_70/Y 0.01fF
C10533 AND2X1_LOC_56/B OR2X1_LOC_719/B 0.02fF
C10534 OR2X1_LOC_325/A OR2X1_LOC_703/A 0.01fF
C10535 OR2X1_LOC_756/B OR2X1_LOC_105/Y 0.00fF
C10536 OR2X1_LOC_185/A OR2X1_LOC_741/Y 0.04fF
C10537 OR2X1_LOC_633/A OR2X1_LOC_240/A 0.01fF
C10538 AND2X1_LOC_566/B OR2X1_LOC_44/Y 0.03fF
C10539 VDD OR2X1_LOC_340/Y 0.20fF
C10540 OR2X1_LOC_121/a_36_216# OR2X1_LOC_574/A 0.17fF
C10541 OR2X1_LOC_641/Y OR2X1_LOC_662/A 0.30fF
C10542 OR2X1_LOC_40/Y OR2X1_LOC_235/a_8_216# 0.01fF
C10543 AND2X1_LOC_651/B OR2X1_LOC_428/A 0.01fF
C10544 AND2X1_LOC_500/Y AND2X1_LOC_807/Y 0.01fF
C10545 VDD OR2X1_LOC_130/A 1.43fF
C10546 AND2X1_LOC_397/a_8_24# OR2X1_LOC_402/Y 0.23fF
C10547 AND2X1_LOC_51/Y OR2X1_LOC_392/B 0.17fF
C10548 OR2X1_LOC_479/Y OR2X1_LOC_161/B 0.24fF
C10549 AND2X1_LOC_784/A AND2X1_LOC_778/Y 0.02fF
C10550 AND2X1_LOC_367/A AND2X1_LOC_841/B 2.23fF
C10551 OR2X1_LOC_620/Y AND2X1_LOC_167/a_8_24# 0.01fF
C10552 VDD AND2X1_LOC_575/Y 0.25fF
C10553 OR2X1_LOC_502/A D_INPUT_4 0.11fF
C10554 OR2X1_LOC_223/A OR2X1_LOC_723/B 0.01fF
C10555 OR2X1_LOC_644/B OR2X1_LOC_676/a_8_216# 0.00fF
C10556 OR2X1_LOC_596/Y OR2X1_LOC_676/Y 0.04fF
C10557 AND2X1_LOC_778/a_8_24# AND2X1_LOC_778/Y 0.08fF
C10558 OR2X1_LOC_756/B OR2X1_LOC_465/Y 0.42fF
C10559 AND2X1_LOC_509/Y AND2X1_LOC_573/A 0.57fF
C10560 OR2X1_LOC_624/A OR2X1_LOC_624/Y 0.00fF
C10561 OR2X1_LOC_599/A AND2X1_LOC_537/a_8_24# 0.01fF
C10562 OR2X1_LOC_744/A AND2X1_LOC_436/B 0.10fF
C10563 AND2X1_LOC_56/B OR2X1_LOC_542/B 0.12fF
C10564 OR2X1_LOC_502/A AND2X1_LOC_423/a_36_24# 0.01fF
C10565 AND2X1_LOC_70/Y OR2X1_LOC_685/B 0.01fF
C10566 OR2X1_LOC_849/a_8_216# OR2X1_LOC_392/B 0.10fF
C10567 OR2X1_LOC_43/Y AND2X1_LOC_729/B 0.02fF
C10568 AND2X1_LOC_22/Y OR2X1_LOC_476/B 0.09fF
C10569 AND2X1_LOC_399/a_8_24# OR2X1_LOC_66/A 0.01fF
C10570 OR2X1_LOC_7/A AND2X1_LOC_448/a_8_24# 0.05fF
C10571 INPUT_0 AND2X1_LOC_655/A 0.03fF
C10572 AND2X1_LOC_302/a_8_24# OR2X1_LOC_59/Y 0.04fF
C10573 INPUT_1 OR2X1_LOC_397/Y 0.13fF
C10574 OR2X1_LOC_40/Y AND2X1_LOC_175/a_36_24# 0.00fF
C10575 AND2X1_LOC_675/Y OR2X1_LOC_680/A 0.23fF
C10576 OR2X1_LOC_850/A OR2X1_LOC_349/A 0.28fF
C10577 VDD AND2X1_LOC_688/a_8_24# 0.00fF
C10578 OR2X1_LOC_40/Y OR2X1_LOC_239/Y 0.06fF
C10579 OR2X1_LOC_123/B OR2X1_LOC_549/A 0.04fF
C10580 AND2X1_LOC_191/B OR2X1_LOC_497/Y 0.07fF
C10581 AND2X1_LOC_95/Y OR2X1_LOC_802/a_8_216# 0.02fF
C10582 AND2X1_LOC_89/a_8_24# OR2X1_LOC_78/A 0.03fF
C10583 AND2X1_LOC_498/a_8_24# OR2X1_LOC_203/Y 0.01fF
C10584 OR2X1_LOC_792/Y OR2X1_LOC_811/A 0.02fF
C10585 OR2X1_LOC_529/a_36_216# OR2X1_LOC_103/Y 0.00fF
C10586 OR2X1_LOC_154/A OR2X1_LOC_624/a_8_216# 0.08fF
C10587 AND2X1_LOC_580/A AND2X1_LOC_549/a_36_24# 0.00fF
C10588 OR2X1_LOC_813/a_8_216# OR2X1_LOC_74/A 0.01fF
C10589 AND2X1_LOC_51/Y OR2X1_LOC_113/B 0.52fF
C10590 OR2X1_LOC_506/a_8_216# OR2X1_LOC_241/Y 0.01fF
C10591 OR2X1_LOC_91/Y OR2X1_LOC_179/a_8_216# 0.05fF
C10592 AND2X1_LOC_667/a_8_24# AND2X1_LOC_44/Y 0.00fF
C10593 OR2X1_LOC_134/Y AND2X1_LOC_227/Y 0.02fF
C10594 OR2X1_LOC_761/a_8_216# OR2X1_LOC_13/B 0.05fF
C10595 OR2X1_LOC_600/A AND2X1_LOC_640/Y 0.03fF
C10596 OR2X1_LOC_516/B OR2X1_LOC_680/A 0.03fF
C10597 AND2X1_LOC_158/a_36_24# OR2X1_LOC_803/A 0.00fF
C10598 AND2X1_LOC_553/A AND2X1_LOC_113/Y 0.25fF
C10599 OR2X1_LOC_36/Y OR2X1_LOC_234/Y 0.02fF
C10600 OR2X1_LOC_533/A OR2X1_LOC_533/a_8_216# 0.01fF
C10601 OR2X1_LOC_323/A AND2X1_LOC_318/Y 0.02fF
C10602 AND2X1_LOC_144/a_8_24# OR2X1_LOC_269/B 0.01fF
C10603 OR2X1_LOC_696/A OR2X1_LOC_184/Y 0.15fF
C10604 AND2X1_LOC_719/Y OR2X1_LOC_64/Y 0.04fF
C10605 AND2X1_LOC_40/Y OR2X1_LOC_456/Y 0.02fF
C10606 OR2X1_LOC_89/a_8_216# OR2X1_LOC_59/Y 0.07fF
C10607 AND2X1_LOC_797/a_8_24# AND2X1_LOC_797/A 0.09fF
C10608 AND2X1_LOC_95/Y OR2X1_LOC_623/a_8_216# 0.06fF
C10609 OR2X1_LOC_335/A OR2X1_LOC_223/A 0.00fF
C10610 OR2X1_LOC_849/a_8_216# OR2X1_LOC_113/B 0.01fF
C10611 AND2X1_LOC_207/A AND2X1_LOC_729/B 0.01fF
C10612 AND2X1_LOC_339/B OR2X1_LOC_46/A 0.07fF
C10613 AND2X1_LOC_737/Y AND2X1_LOC_811/a_8_24# 0.19fF
C10614 AND2X1_LOC_777/a_8_24# AND2X1_LOC_857/Y 0.01fF
C10615 OR2X1_LOC_92/Y OR2X1_LOC_67/a_36_216# 0.00fF
C10616 OR2X1_LOC_325/a_36_216# AND2X1_LOC_59/Y 0.00fF
C10617 OR2X1_LOC_653/A OR2X1_LOC_502/A 0.02fF
C10618 OR2X1_LOC_529/Y OR2X1_LOC_744/A 0.04fF
C10619 OR2X1_LOC_92/Y OR2X1_LOC_6/A 0.14fF
C10620 OR2X1_LOC_479/Y OR2X1_LOC_785/a_36_216# 0.00fF
C10621 OR2X1_LOC_167/Y OR2X1_LOC_16/A 0.03fF
C10622 OR2X1_LOC_318/B OR2X1_LOC_301/a_8_216# 0.01fF
C10623 OR2X1_LOC_103/Y AND2X1_LOC_361/A 0.17fF
C10624 OR2X1_LOC_553/B OR2X1_LOC_553/A 0.10fF
C10625 D_INPUT_5 AND2X1_LOC_472/B 0.11fF
C10626 OR2X1_LOC_51/Y AND2X1_LOC_483/a_36_24# 0.01fF
C10627 AND2X1_LOC_360/a_36_24# OR2X1_LOC_44/Y 0.01fF
C10628 AND2X1_LOC_148/a_8_24# AND2X1_LOC_148/Y 0.00fF
C10629 OR2X1_LOC_185/Y OR2X1_LOC_856/B 0.14fF
C10630 OR2X1_LOC_228/Y OR2X1_LOC_539/B 0.02fF
C10631 OR2X1_LOC_811/A OR2X1_LOC_87/A 0.01fF
C10632 OR2X1_LOC_600/A OR2X1_LOC_416/Y 0.03fF
C10633 AND2X1_LOC_802/B OR2X1_LOC_47/Y 0.03fF
C10634 OR2X1_LOC_405/Y OR2X1_LOC_215/Y 0.00fF
C10635 OR2X1_LOC_689/A AND2X1_LOC_688/a_8_24# 0.01fF
C10636 AND2X1_LOC_779/a_8_24# OR2X1_LOC_599/A 0.03fF
C10637 OR2X1_LOC_808/A OR2X1_LOC_787/Y 0.00fF
C10638 AND2X1_LOC_40/Y OR2X1_LOC_810/A 0.03fF
C10639 AND2X1_LOC_729/Y AND2X1_LOC_624/A 0.03fF
C10640 OR2X1_LOC_80/Y OR2X1_LOC_393/Y 0.18fF
C10641 AND2X1_LOC_143/a_36_24# OR2X1_LOC_585/A 0.01fF
C10642 OR2X1_LOC_715/B D_INPUT_0 0.11fF
C10643 OR2X1_LOC_427/A AND2X1_LOC_818/a_8_24# 0.01fF
C10644 OR2X1_LOC_685/A OR2X1_LOC_161/A 0.01fF
C10645 AND2X1_LOC_681/a_8_24# OR2X1_LOC_161/B 0.01fF
C10646 AND2X1_LOC_663/B OR2X1_LOC_59/Y 0.04fF
C10647 OR2X1_LOC_696/A OR2X1_LOC_70/A 0.02fF
C10648 OR2X1_LOC_673/A AND2X1_LOC_277/a_8_24# 0.01fF
C10649 OR2X1_LOC_625/Y OR2X1_LOC_248/a_36_216# 0.03fF
C10650 AND2X1_LOC_719/Y OR2X1_LOC_417/A 3.68fF
C10651 OR2X1_LOC_358/a_8_216# OR2X1_LOC_805/A 0.05fF
C10652 OR2X1_LOC_606/Y OR2X1_LOC_66/A 0.07fF
C10653 VDD OR2X1_LOC_62/B 1.24fF
C10654 OR2X1_LOC_194/B OR2X1_LOC_269/B 0.05fF
C10655 OR2X1_LOC_502/A OR2X1_LOC_195/A 0.02fF
C10656 OR2X1_LOC_185/Y OR2X1_LOC_793/a_8_216# 0.01fF
C10657 OR2X1_LOC_810/a_8_216# OR2X1_LOC_810/A 0.06fF
C10658 AND2X1_LOC_753/B AND2X1_LOC_3/Y 0.04fF
C10659 OR2X1_LOC_147/A AND2X1_LOC_51/Y 0.01fF
C10660 OR2X1_LOC_427/A AND2X1_LOC_454/A 0.03fF
C10661 AND2X1_LOC_580/B OR2X1_LOC_18/Y 0.02fF
C10662 AND2X1_LOC_40/Y AND2X1_LOC_589/a_8_24# 0.01fF
C10663 OR2X1_LOC_274/Y OR2X1_LOC_778/A 0.08fF
C10664 AND2X1_LOC_99/A AND2X1_LOC_123/a_8_24# 0.01fF
C10665 OR2X1_LOC_8/Y INPUT_1 1.48fF
C10666 OR2X1_LOC_665/Y OR2X1_LOC_625/Y 0.03fF
C10667 AND2X1_LOC_19/Y AND2X1_LOC_48/A 0.03fF
C10668 AND2X1_LOC_713/Y OR2X1_LOC_31/Y 0.01fF
C10669 OR2X1_LOC_294/Y OR2X1_LOC_284/B 0.01fF
C10670 OR2X1_LOC_49/A OR2X1_LOC_396/Y 0.03fF
C10671 AND2X1_LOC_338/a_36_24# OR2X1_LOC_46/A 0.00fF
C10672 OR2X1_LOC_400/A OR2X1_LOC_673/Y 0.01fF
C10673 OR2X1_LOC_50/a_36_216# INPUT_7 0.00fF
C10674 AND2X1_LOC_841/B OR2X1_LOC_74/A 0.00fF
C10675 AND2X1_LOC_549/Y OR2X1_LOC_95/Y 0.03fF
C10676 OR2X1_LOC_405/A AND2X1_LOC_3/Y 2.06fF
C10677 OR2X1_LOC_168/A OR2X1_LOC_78/A 0.05fF
C10678 OR2X1_LOC_485/A OR2X1_LOC_625/Y 0.11fF
C10679 VDD OR2X1_LOC_780/B 0.21fF
C10680 OR2X1_LOC_287/B OR2X1_LOC_377/A 0.04fF
C10681 AND2X1_LOC_64/Y AND2X1_LOC_31/Y 1.54fF
C10682 OR2X1_LOC_147/a_8_216# OR2X1_LOC_375/A 0.00fF
C10683 OR2X1_LOC_95/Y OR2X1_LOC_627/Y 0.02fF
C10684 OR2X1_LOC_271/Y OR2X1_LOC_6/A 0.01fF
C10685 OR2X1_LOC_375/A OR2X1_LOC_564/A 0.01fF
C10686 AND2X1_LOC_500/Y OR2X1_LOC_95/Y 0.03fF
C10687 AND2X1_LOC_727/Y OR2X1_LOC_152/A 0.01fF
C10688 OR2X1_LOC_574/A OR2X1_LOC_799/a_8_216# 0.06fF
C10689 AND2X1_LOC_364/Y D_INPUT_0 0.16fF
C10690 OR2X1_LOC_835/a_8_216# OR2X1_LOC_269/B -0.03fF
C10691 OR2X1_LOC_357/a_8_216# OR2X1_LOC_365/B 0.01fF
C10692 OR2X1_LOC_462/B AND2X1_LOC_234/a_8_24# 0.01fF
C10693 AND2X1_LOC_91/B OR2X1_LOC_561/B 0.00fF
C10694 VDD AND2X1_LOC_796/Y 0.21fF
C10695 OR2X1_LOC_137/Y OR2X1_LOC_673/Y 0.00fF
C10696 AND2X1_LOC_1/Y AND2X1_LOC_11/Y 0.07fF
C10697 AND2X1_LOC_326/B AND2X1_LOC_851/B 0.83fF
C10698 AND2X1_LOC_544/Y OR2X1_LOC_152/a_8_216# 0.05fF
C10699 OR2X1_LOC_835/B AND2X1_LOC_822/a_8_24# 0.04fF
C10700 OR2X1_LOC_859/B OR2X1_LOC_810/A 0.03fF
C10701 OR2X1_LOC_864/a_8_216# OR2X1_LOC_848/A 0.01fF
C10702 OR2X1_LOC_377/A OR2X1_LOC_97/a_8_216# 0.01fF
C10703 AND2X1_LOC_716/Y AND2X1_LOC_326/a_8_24# 0.01fF
C10704 OR2X1_LOC_585/A OR2X1_LOC_49/a_8_216# 0.01fF
C10705 OR2X1_LOC_786/Y OR2X1_LOC_66/A 0.02fF
C10706 OR2X1_LOC_32/B OR2X1_LOC_60/a_8_216# 0.03fF
C10707 OR2X1_LOC_311/Y AND2X1_LOC_809/A 0.03fF
C10708 OR2X1_LOC_79/A OR2X1_LOC_36/Y 0.47fF
C10709 OR2X1_LOC_416/Y OR2X1_LOC_619/Y 0.03fF
C10710 OR2X1_LOC_562/Y OR2X1_LOC_562/B 0.00fF
C10711 OR2X1_LOC_161/B OR2X1_LOC_68/B 0.07fF
C10712 OR2X1_LOC_160/A AND2X1_LOC_680/a_8_24# 0.04fF
C10713 OR2X1_LOC_64/Y AND2X1_LOC_655/A 0.05fF
C10714 OR2X1_LOC_817/Y OR2X1_LOC_44/Y 0.02fF
C10715 OR2X1_LOC_685/A AND2X1_LOC_51/Y 0.01fF
C10716 AND2X1_LOC_12/Y OR2X1_LOC_19/B 0.10fF
C10717 OR2X1_LOC_89/A AND2X1_LOC_645/A 0.02fF
C10718 AND2X1_LOC_154/Y OR2X1_LOC_52/B 0.58fF
C10719 INPUT_3 AND2X1_LOC_672/B 0.02fF
C10720 AND2X1_LOC_76/Y INPUT_1 0.20fF
C10721 OR2X1_LOC_447/Y OR2X1_LOC_714/Y 0.04fF
C10722 D_INPUT_3 AND2X1_LOC_819/a_36_24# 0.01fF
C10723 AND2X1_LOC_830/a_8_24# OR2X1_LOC_36/Y 0.01fF
C10724 OR2X1_LOC_626/a_8_216# OR2X1_LOC_617/a_8_216# 0.47fF
C10725 OR2X1_LOC_825/Y OR2X1_LOC_85/A 0.10fF
C10726 OR2X1_LOC_48/Y OR2X1_LOC_585/A 0.03fF
C10727 OR2X1_LOC_677/Y AND2X1_LOC_796/Y 0.09fF
C10728 OR2X1_LOC_51/Y AND2X1_LOC_845/a_8_24# 0.04fF
C10729 OR2X1_LOC_687/A OR2X1_LOC_451/B 0.01fF
C10730 VDD OR2X1_LOC_365/B 0.30fF
C10731 AND2X1_LOC_633/a_8_24# OR2X1_LOC_46/A 0.12fF
C10732 AND2X1_LOC_36/Y AND2X1_LOC_763/B 0.01fF
C10733 OR2X1_LOC_401/Y AND2X1_LOC_490/a_36_24# 0.00fF
C10734 OR2X1_LOC_377/A OR2X1_LOC_835/Y 0.34fF
C10735 OR2X1_LOC_160/A OR2X1_LOC_243/B 0.95fF
C10736 OR2X1_LOC_3/Y OR2X1_LOC_817/a_8_216# 0.01fF
C10737 AND2X1_LOC_663/B OR2X1_LOC_820/B 0.03fF
C10738 OR2X1_LOC_240/B OR2X1_LOC_532/B 0.01fF
C10739 AND2X1_LOC_110/Y OR2X1_LOC_854/A 0.00fF
C10740 OR2X1_LOC_412/a_8_216# OR2X1_LOC_39/A 0.01fF
C10741 INPUT_0 OR2X1_LOC_599/Y 0.11fF
C10742 OR2X1_LOC_36/Y OR2X1_LOC_278/A 0.08fF
C10743 OR2X1_LOC_62/A AND2X1_LOC_619/B 0.03fF
C10744 OR2X1_LOC_532/B OR2X1_LOC_161/A 0.24fF
C10745 AND2X1_LOC_147/Y AND2X1_LOC_149/a_8_24# 0.09fF
C10746 OR2X1_LOC_437/A AND2X1_LOC_786/Y 0.10fF
C10747 AND2X1_LOC_35/a_8_24# D_INPUT_0 0.01fF
C10748 OR2X1_LOC_699/a_8_216# OR2X1_LOC_46/A 0.01fF
C10749 AND2X1_LOC_191/Y AND2X1_LOC_797/A 0.03fF
C10750 OR2X1_LOC_519/Y OR2X1_LOC_31/Y 0.00fF
C10751 AND2X1_LOC_280/a_8_24# OR2X1_LOC_78/A 0.02fF
C10752 OR2X1_LOC_744/A OR2X1_LOC_598/A 0.04fF
C10753 OR2X1_LOC_62/B OR2X1_LOC_267/a_36_216# 0.00fF
C10754 OR2X1_LOC_417/A AND2X1_LOC_655/A 0.01fF
C10755 OR2X1_LOC_31/Y AND2X1_LOC_436/B 0.01fF
C10756 AND2X1_LOC_811/Y AND2X1_LOC_808/a_36_24# 0.00fF
C10757 OR2X1_LOC_600/A OR2X1_LOC_80/A 0.50fF
C10758 AND2X1_LOC_139/B OR2X1_LOC_31/Y 0.13fF
C10759 OR2X1_LOC_263/a_8_216# OR2X1_LOC_86/a_8_216# 0.47fF
C10760 OR2X1_LOC_26/Y AND2X1_LOC_477/A 0.04fF
C10761 OR2X1_LOC_549/A OR2X1_LOC_367/a_8_216# 0.04fF
C10762 AND2X1_LOC_711/Y AND2X1_LOC_663/B 2.31fF
C10763 OR2X1_LOC_47/Y OR2X1_LOC_256/a_8_216# 0.01fF
C10764 OR2X1_LOC_634/a_8_216# OR2X1_LOC_598/A 0.01fF
C10765 AND2X1_LOC_851/B OR2X1_LOC_237/a_8_216# 0.06fF
C10766 OR2X1_LOC_72/a_36_216# OR2X1_LOC_265/Y 0.00fF
C10767 OR2X1_LOC_720/B OR2X1_LOC_720/a_8_216# 0.02fF
C10768 OR2X1_LOC_78/B OR2X1_LOC_228/Y 0.11fF
C10769 INPUT_1 OR2X1_LOC_52/B 0.50fF
C10770 OR2X1_LOC_470/B AND2X1_LOC_51/Y 0.10fF
C10771 AND2X1_LOC_81/a_8_24# D_INPUT_0 0.02fF
C10772 OR2X1_LOC_742/B D_GATE_741 0.18fF
C10773 AND2X1_LOC_792/Y AND2X1_LOC_805/Y 0.01fF
C10774 AND2X1_LOC_477/A OR2X1_LOC_89/A 0.03fF
C10775 OR2X1_LOC_473/A OR2X1_LOC_375/A 0.02fF
C10776 OR2X1_LOC_849/A AND2X1_LOC_47/Y 0.03fF
C10777 OR2X1_LOC_70/Y AND2X1_LOC_686/a_8_24# 0.02fF
C10778 AND2X1_LOC_717/B OR2X1_LOC_226/Y 0.13fF
C10779 OR2X1_LOC_464/A AND2X1_LOC_31/Y 0.03fF
C10780 AND2X1_LOC_468/B OR2X1_LOC_419/Y 0.03fF
C10781 AND2X1_LOC_338/Y OR2X1_LOC_171/Y 0.16fF
C10782 OR2X1_LOC_653/Y OR2X1_LOC_358/A 0.01fF
C10783 OR2X1_LOC_512/A AND2X1_LOC_31/Y 0.01fF
C10784 OR2X1_LOC_429/Y OR2X1_LOC_70/a_8_216# 0.05fF
C10785 OR2X1_LOC_244/Y OR2X1_LOC_342/a_8_216# 0.01fF
C10786 OR2X1_LOC_653/a_36_216# OR2X1_LOC_532/B 0.00fF
C10787 OR2X1_LOC_529/Y OR2X1_LOC_31/Y 0.01fF
C10788 OR2X1_LOC_115/B AND2X1_LOC_44/Y 0.05fF
C10789 AND2X1_LOC_92/Y OR2X1_LOC_303/B 0.02fF
C10790 OR2X1_LOC_541/B OR2X1_LOC_598/A 0.00fF
C10791 AND2X1_LOC_618/a_8_24# OR2X1_LOC_68/B 0.03fF
C10792 OR2X1_LOC_416/Y AND2X1_LOC_462/a_8_24# 0.01fF
C10793 AND2X1_LOC_70/Y OR2X1_LOC_544/B 0.01fF
C10794 AND2X1_LOC_102/a_36_24# OR2X1_LOC_62/A 0.01fF
C10795 OR2X1_LOC_61/Y OR2X1_LOC_68/B 0.24fF
C10796 AND2X1_LOC_437/a_8_24# OR2X1_LOC_788/B 0.02fF
C10797 OR2X1_LOC_516/Y OR2X1_LOC_528/Y 0.03fF
C10798 OR2X1_LOC_532/B AND2X1_LOC_51/Y 0.13fF
C10799 OR2X1_LOC_22/Y AND2X1_LOC_116/B 0.01fF
C10800 OR2X1_LOC_205/Y OR2X1_LOC_217/a_8_216# 0.07fF
C10801 AND2X1_LOC_208/Y AND2X1_LOC_214/a_8_24# 0.02fF
C10802 AND2X1_LOC_350/Y OR2X1_LOC_417/A 0.13fF
C10803 OR2X1_LOC_45/B OR2X1_LOC_79/a_36_216# 0.02fF
C10804 AND2X1_LOC_101/B OR2X1_LOC_86/A 0.16fF
C10805 OR2X1_LOC_375/A OR2X1_LOC_228/Y 0.01fF
C10806 AND2X1_LOC_65/A AND2X1_LOC_7/B 0.04fF
C10807 OR2X1_LOC_87/a_8_216# OR2X1_LOC_68/B 0.04fF
C10808 OR2X1_LOC_45/B OR2X1_LOC_693/a_8_216# 0.02fF
C10809 AND2X1_LOC_259/Y AND2X1_LOC_259/a_8_24# 0.01fF
C10810 OR2X1_LOC_375/A OR2X1_LOC_513/Y 0.01fF
C10811 AND2X1_LOC_280/a_36_24# OR2X1_LOC_366/Y 0.01fF
C10812 OR2X1_LOC_787/Y OR2X1_LOC_374/Y 0.68fF
C10813 AND2X1_LOC_357/a_36_24# OR2X1_LOC_437/A 0.00fF
C10814 AND2X1_LOC_22/Y AND2X1_LOC_262/a_8_24# 0.04fF
C10815 AND2X1_LOC_84/Y VDD 0.01fF
C10816 OR2X1_LOC_64/Y AND2X1_LOC_687/a_36_24# 0.00fF
C10817 OR2X1_LOC_186/Y OR2X1_LOC_151/A 0.13fF
C10818 AND2X1_LOC_55/a_8_24# OR2X1_LOC_71/A 0.02fF
C10819 OR2X1_LOC_64/Y OR2X1_LOC_599/Y 0.21fF
C10820 OR2X1_LOC_604/A OR2X1_LOC_744/a_36_216# 0.00fF
C10821 AND2X1_LOC_47/Y OR2X1_LOC_440/A 0.04fF
C10822 OR2X1_LOC_201/a_36_216# OR2X1_LOC_532/B 0.01fF
C10823 OR2X1_LOC_528/Y AND2X1_LOC_547/a_8_24# 0.00fF
C10824 OR2X1_LOC_329/B AND2X1_LOC_465/A 0.72fF
C10825 OR2X1_LOC_45/B OR2X1_LOC_695/Y 0.02fF
C10826 OR2X1_LOC_619/a_8_216# D_INPUT_0 0.01fF
C10827 OR2X1_LOC_634/A OR2X1_LOC_334/A 0.09fF
C10828 OR2X1_LOC_490/a_8_216# AND2X1_LOC_243/Y 0.02fF
C10829 OR2X1_LOC_124/a_8_216# AND2X1_LOC_44/Y 0.01fF
C10830 OR2X1_LOC_624/A OR2X1_LOC_174/Y 0.04fF
C10831 OR2X1_LOC_47/Y AND2X1_LOC_835/a_8_24# 0.01fF
C10832 AND2X1_LOC_41/A OR2X1_LOC_120/a_8_216# 0.05fF
C10833 OR2X1_LOC_160/A OR2X1_LOC_771/B 0.05fF
C10834 OR2X1_LOC_852/a_8_216# VDD -0.00fF
C10835 OR2X1_LOC_9/Y OR2X1_LOC_158/A 0.29fF
C10836 AND2X1_LOC_715/A AND2X1_LOC_786/Y 0.02fF
C10837 OR2X1_LOC_703/B OR2X1_LOC_777/B 0.06fF
C10838 AND2X1_LOC_567/a_8_24# AND2X1_LOC_810/B 0.03fF
C10839 OR2X1_LOC_64/Y OR2X1_LOC_331/a_8_216# 0.04fF
C10840 AND2X1_LOC_724/A VDD 0.21fF
C10841 AND2X1_LOC_91/a_36_24# AND2X1_LOC_70/Y 0.01fF
C10842 OR2X1_LOC_22/Y AND2X1_LOC_204/Y 0.04fF
C10843 OR2X1_LOC_22/Y OR2X1_LOC_311/a_8_216# 0.03fF
C10844 OR2X1_LOC_87/A OR2X1_LOC_777/B 0.07fF
C10845 OR2X1_LOC_488/Y AND2X1_LOC_563/Y 0.32fF
C10846 AND2X1_LOC_141/a_8_24# OR2X1_LOC_12/Y 0.01fF
C10847 AND2X1_LOC_59/Y OR2X1_LOC_308/Y 0.07fF
C10848 OR2X1_LOC_62/B OR2X1_LOC_140/a_8_216# 0.01fF
C10849 OR2X1_LOC_3/Y OR2X1_LOC_384/Y 0.79fF
C10850 AND2X1_LOC_47/a_36_24# INPUT_6 0.00fF
C10851 OR2X1_LOC_653/B OR2X1_LOC_648/A 0.02fF
C10852 OR2X1_LOC_158/A AND2X1_LOC_61/Y 0.08fF
C10853 OR2X1_LOC_516/A OR2X1_LOC_516/Y 0.01fF
C10854 OR2X1_LOC_206/A AND2X1_LOC_31/Y 0.01fF
C10855 OR2X1_LOC_427/A AND2X1_LOC_783/B 0.01fF
C10856 OR2X1_LOC_676/Y OR2X1_LOC_596/a_36_216# 0.01fF
C10857 AND2X1_LOC_534/a_8_24# OR2X1_LOC_538/A 0.01fF
C10858 AND2X1_LOC_362/B AND2X1_LOC_121/a_8_24# 0.04fF
C10859 OR2X1_LOC_632/A OR2X1_LOC_140/B 0.01fF
C10860 OR2X1_LOC_3/B OR2X1_LOC_587/a_8_216# 0.01fF
C10861 OR2X1_LOC_840/A AND2X1_LOC_44/Y 0.01fF
C10862 AND2X1_LOC_578/A OR2X1_LOC_437/A 0.02fF
C10863 OR2X1_LOC_441/Y AND2X1_LOC_213/B 0.03fF
C10864 OR2X1_LOC_31/Y OR2X1_LOC_598/A 0.06fF
C10865 OR2X1_LOC_421/A OR2X1_LOC_51/Y 0.01fF
C10866 OR2X1_LOC_834/A OR2X1_LOC_307/A 0.03fF
C10867 AND2X1_LOC_348/A OR2X1_LOC_428/A 0.00fF
C10868 VDD OR2X1_LOC_468/A 0.26fF
C10869 AND2X1_LOC_600/a_8_24# AND2X1_LOC_31/Y 0.01fF
C10870 OR2X1_LOC_511/Y OR2X1_LOC_525/a_8_216# 0.03fF
C10871 OR2X1_LOC_181/B AND2X1_LOC_7/B 0.03fF
C10872 AND2X1_LOC_41/A OR2X1_LOC_596/A 0.11fF
C10873 OR2X1_LOC_95/Y OR2X1_LOC_387/a_36_216# 0.00fF
C10874 AND2X1_LOC_367/A OR2X1_LOC_322/Y 0.49fF
C10875 VDD OR2X1_LOC_666/A 0.37fF
C10876 OR2X1_LOC_104/a_8_216# OR2X1_LOC_600/A 0.02fF
C10877 AND2X1_LOC_43/B AND2X1_LOC_416/a_8_24# 0.04fF
C10878 OR2X1_LOC_375/A OR2X1_LOC_562/A 0.03fF
C10879 AND2X1_LOC_477/a_8_24# AND2X1_LOC_477/Y 0.02fF
C10880 AND2X1_LOC_392/A OR2X1_LOC_59/Y 0.03fF
C10881 OR2X1_LOC_624/B OR2X1_LOC_771/B 0.07fF
C10882 OR2X1_LOC_33/a_8_216# OR2X1_LOC_771/B 0.05fF
C10883 AND2X1_LOC_571/A OR2X1_LOC_44/Y 0.03fF
C10884 OR2X1_LOC_538/A AND2X1_LOC_110/Y 0.02fF
C10885 OR2X1_LOC_56/A AND2X1_LOC_285/Y 0.03fF
C10886 AND2X1_LOC_810/A AND2X1_LOC_841/B 0.03fF
C10887 OR2X1_LOC_181/B OR2X1_LOC_564/a_8_216# 0.47fF
C10888 OR2X1_LOC_176/Y AND2X1_LOC_170/a_8_24# 0.29fF
C10889 OR2X1_LOC_95/Y AND2X1_LOC_563/Y 0.00fF
C10890 OR2X1_LOC_303/a_8_216# OR2X1_LOC_468/Y 0.01fF
C10891 OR2X1_LOC_87/A OR2X1_LOC_831/B 0.07fF
C10892 OR2X1_LOC_709/A OR2X1_LOC_724/a_8_216# 0.06fF
C10893 AND2X1_LOC_315/a_8_24# OR2X1_LOC_161/B 0.05fF
C10894 OR2X1_LOC_715/B AND2X1_LOC_40/Y 0.01fF
C10895 VDD OR2X1_LOC_762/Y 0.17fF
C10896 AND2X1_LOC_64/Y OR2X1_LOC_864/A 0.03fF
C10897 OR2X1_LOC_744/A OR2X1_LOC_484/a_8_216# 0.01fF
C10898 OR2X1_LOC_156/Y OR2X1_LOC_87/A 0.09fF
C10899 VDD OR2X1_LOC_659/A 0.00fF
C10900 AND2X1_LOC_95/Y OR2X1_LOC_294/Y 0.03fF
C10901 OR2X1_LOC_45/B OR2X1_LOC_406/a_8_216# 0.01fF
C10902 OR2X1_LOC_53/Y AND2X1_LOC_193/a_36_24# 0.00fF
C10903 OR2X1_LOC_12/Y AND2X1_LOC_447/a_8_24# -0.00fF
C10904 AND2X1_LOC_170/a_8_24# AND2X1_LOC_212/Y 0.02fF
C10905 OR2X1_LOC_286/B OR2X1_LOC_366/Y 0.03fF
C10906 AND2X1_LOC_456/B OR2X1_LOC_51/Y 0.05fF
C10907 AND2X1_LOC_734/Y AND2X1_LOC_657/Y 0.03fF
C10908 AND2X1_LOC_366/A OR2X1_LOC_59/Y 0.06fF
C10909 AND2X1_LOC_505/a_36_24# OR2X1_LOC_502/A 0.00fF
C10910 AND2X1_LOC_64/Y OR2X1_LOC_633/B 0.03fF
C10911 OR2X1_LOC_9/Y OR2X1_LOC_847/A 0.02fF
C10912 AND2X1_LOC_716/Y VDD -0.00fF
C10913 OR2X1_LOC_858/A OR2X1_LOC_756/B 0.14fF
C10914 AND2X1_LOC_598/a_8_24# AND2X1_LOC_703/Y 0.20fF
C10915 OR2X1_LOC_733/A OR2X1_LOC_737/A 0.04fF
C10916 AND2X1_LOC_735/Y AND2X1_LOC_736/a_8_24# 0.11fF
C10917 OR2X1_LOC_97/A OR2X1_LOC_269/B 0.03fF
C10918 AND2X1_LOC_543/Y OR2X1_LOC_74/A 0.04fF
C10919 OR2X1_LOC_114/a_36_216# OR2X1_LOC_235/B 0.00fF
C10920 OR2X1_LOC_725/B OR2X1_LOC_66/A 0.01fF
C10921 VDD AND2X1_LOC_654/Y 0.80fF
C10922 OR2X1_LOC_851/A OR2X1_LOC_841/A 0.01fF
C10923 OR2X1_LOC_135/Y OR2X1_LOC_36/Y 0.01fF
C10924 OR2X1_LOC_604/A AND2X1_LOC_468/B 0.01fF
C10925 AND2X1_LOC_81/B OR2X1_LOC_151/A 0.03fF
C10926 OR2X1_LOC_375/A OR2X1_LOC_786/a_36_216# 0.00fF
C10927 AND2X1_LOC_12/Y AND2X1_LOC_110/Y 0.00fF
C10928 OR2X1_LOC_440/B OR2X1_LOC_161/A 0.04fF
C10929 AND2X1_LOC_570/Y OR2X1_LOC_427/A 0.14fF
C10930 AND2X1_LOC_573/A AND2X1_LOC_489/a_8_24# 0.01fF
C10931 AND2X1_LOC_150/a_8_24# OR2X1_LOC_87/A 0.03fF
C10932 OR2X1_LOC_158/A OR2X1_LOC_96/B 0.03fF
C10933 OR2X1_LOC_160/B OR2X1_LOC_377/A 0.02fF
C10934 AND2X1_LOC_340/a_36_24# OR2X1_LOC_65/B 0.00fF
C10935 D_GATE_662 OR2X1_LOC_269/B 0.02fF
C10936 AND2X1_LOC_212/A AND2X1_LOC_661/A 0.02fF
C10937 OR2X1_LOC_114/B OR2X1_LOC_664/Y 0.03fF
C10938 AND2X1_LOC_364/A OR2X1_LOC_91/A 0.46fF
C10939 AND2X1_LOC_729/Y AND2X1_LOC_803/B 0.00fF
C10940 OR2X1_LOC_158/A AND2X1_LOC_852/Y 0.08fF
C10941 OR2X1_LOC_154/A AND2X1_LOC_313/a_8_24# 0.02fF
C10942 OR2X1_LOC_828/B OR2X1_LOC_66/A 0.14fF
C10943 OR2X1_LOC_674/a_8_216# AND2X1_LOC_840/A 0.47fF
C10944 OR2X1_LOC_686/A OR2X1_LOC_87/A 0.02fF
C10945 OR2X1_LOC_426/B OR2X1_LOC_316/Y 0.03fF
C10946 AND2X1_LOC_42/B OR2X1_LOC_548/B 0.04fF
C10947 OR2X1_LOC_404/Y OR2X1_LOC_474/B 0.07fF
C10948 OR2X1_LOC_6/B OR2X1_LOC_643/A 0.07fF
C10949 OR2X1_LOC_600/A OR2X1_LOC_6/A 5.32fF
C10950 OR2X1_LOC_160/B OR2X1_LOC_203/Y 0.07fF
C10951 OR2X1_LOC_6/B OR2X1_LOC_124/Y 0.05fF
C10952 AND2X1_LOC_476/A OR2X1_LOC_268/Y 0.02fF
C10953 OR2X1_LOC_52/B AND2X1_LOC_778/Y 0.00fF
C10954 VDD GATE_366 0.17fF
C10955 OR2X1_LOC_856/A OR2X1_LOC_856/a_8_216# 0.18fF
C10956 AND2X1_LOC_548/Y OR2X1_LOC_39/A 0.01fF
C10957 OR2X1_LOC_52/Y AND2X1_LOC_214/a_8_24# 0.24fF
C10958 AND2X1_LOC_76/Y OR2X1_LOC_517/A 0.01fF
C10959 OR2X1_LOC_216/A AND2X1_LOC_492/a_8_24# 0.05fF
C10960 OR2X1_LOC_91/Y OR2X1_LOC_56/A 0.03fF
C10961 OR2X1_LOC_763/a_8_216# OR2X1_LOC_48/B 0.10fF
C10962 OR2X1_LOC_589/A OR2X1_LOC_74/A 0.03fF
C10963 AND2X1_LOC_56/B OR2X1_LOC_787/B 0.01fF
C10964 OR2X1_LOC_426/B AND2X1_LOC_354/B 0.12fF
C10965 OR2X1_LOC_329/B OR2X1_LOC_237/Y 0.05fF
C10966 OR2X1_LOC_53/Y OR2X1_LOC_22/Y 0.07fF
C10967 OR2X1_LOC_687/B OR2X1_LOC_687/A 0.15fF
C10968 AND2X1_LOC_357/B AND2X1_LOC_211/B 0.07fF
C10969 VDD OR2X1_LOC_449/B 0.27fF
C10970 OR2X1_LOC_74/A OR2X1_LOC_322/Y 0.10fF
C10971 OR2X1_LOC_18/Y OR2X1_LOC_763/a_8_216# 0.01fF
C10972 OR2X1_LOC_484/a_8_216# AND2X1_LOC_840/B 0.27fF
C10973 OR2X1_LOC_3/Y OR2X1_LOC_131/a_8_216# 0.01fF
C10974 AND2X1_LOC_56/B AND2X1_LOC_92/Y 1.27fF
C10975 OR2X1_LOC_305/Y OR2X1_LOC_56/A 0.00fF
C10976 OR2X1_LOC_302/B AND2X1_LOC_298/a_8_24# 0.02fF
C10977 OR2X1_LOC_405/A OR2X1_LOC_775/a_8_216# 0.01fF
C10978 VDD OR2X1_LOC_312/Y 0.48fF
C10979 AND2X1_LOC_42/B OR2X1_LOC_786/A 0.05fF
C10980 AND2X1_LOC_358/Y AND2X1_LOC_537/Y 0.09fF
C10981 OR2X1_LOC_521/Y AND2X1_LOC_76/Y 0.01fF
C10982 AND2X1_LOC_537/a_8_24# OR2X1_LOC_7/A 0.05fF
C10983 AND2X1_LOC_347/B OR2X1_LOC_258/Y 0.01fF
C10984 OR2X1_LOC_517/A OR2X1_LOC_67/A 0.02fF
C10985 OR2X1_LOC_46/A AND2X1_LOC_219/A 0.03fF
C10986 OR2X1_LOC_160/A OR2X1_LOC_637/B 0.25fF
C10987 AND2X1_LOC_8/Y AND2X1_LOC_92/Y 2.07fF
C10988 AND2X1_LOC_191/Y AND2X1_LOC_807/B 0.03fF
C10989 OR2X1_LOC_106/Y AND2X1_LOC_227/Y 0.03fF
C10990 OR2X1_LOC_22/Y AND2X1_LOC_802/Y 0.15fF
C10991 OR2X1_LOC_696/A OR2X1_LOC_47/Y 0.26fF
C10992 OR2X1_LOC_51/Y AND2X1_LOC_717/B 0.03fF
C10993 OR2X1_LOC_756/B OR2X1_LOC_593/a_8_216# 0.01fF
C10994 AND2X1_LOC_571/a_8_24# OR2X1_LOC_71/Y 0.01fF
C10995 AND2X1_LOC_557/a_8_24# OR2X1_LOC_600/A 0.04fF
C10996 OR2X1_LOC_581/a_8_216# D_INPUT_6 0.07fF
C10997 AND2X1_LOC_776/a_8_24# OR2X1_LOC_371/Y 0.01fF
C10998 AND2X1_LOC_711/Y AND2X1_LOC_807/B 0.03fF
C10999 AND2X1_LOC_565/B AND2X1_LOC_711/Y 0.08fF
C11000 AND2X1_LOC_392/A OR2X1_LOC_70/Y 0.01fF
C11001 AND2X1_LOC_95/Y OR2X1_LOC_730/a_8_216# 0.01fF
C11002 AND2X1_LOC_773/Y D_INPUT_0 2.03fF
C11003 OR2X1_LOC_18/Y OR2X1_LOC_278/Y 0.02fF
C11004 AND2X1_LOC_738/B OR2X1_LOC_152/Y 0.04fF
C11005 AND2X1_LOC_565/B OR2X1_LOC_70/Y 0.03fF
C11006 OR2X1_LOC_179/a_36_216# OR2X1_LOC_44/Y 0.02fF
C11007 OR2X1_LOC_287/B OR2X1_LOC_78/B 0.06fF
C11008 AND2X1_LOC_390/B OR2X1_LOC_426/B 0.72fF
C11009 OR2X1_LOC_121/B AND2X1_LOC_265/a_8_24# 0.01fF
C11010 OR2X1_LOC_814/A OR2X1_LOC_390/A 0.07fF
C11011 AND2X1_LOC_807/Y AND2X1_LOC_805/Y 0.01fF
C11012 OR2X1_LOC_692/a_8_216# OR2X1_LOC_44/Y 0.01fF
C11013 OR2X1_LOC_45/B AND2X1_LOC_675/A 0.02fF
C11014 OR2X1_LOC_484/Y OR2X1_LOC_485/A 0.56fF
C11015 INPUT_3 OR2X1_LOC_377/A 0.01fF
C11016 OR2X1_LOC_92/Y OR2X1_LOC_44/Y 0.13fF
C11017 AND2X1_LOC_211/B AND2X1_LOC_303/a_8_24# 0.01fF
C11018 AND2X1_LOC_391/Y OR2X1_LOC_3/Y 0.04fF
C11019 OR2X1_LOC_850/a_36_216# OR2X1_LOC_287/B 0.00fF
C11020 OR2X1_LOC_517/A OR2X1_LOC_52/B 0.19fF
C11021 OR2X1_LOC_62/B OR2X1_LOC_361/a_36_216# 0.00fF
C11022 OR2X1_LOC_513/Y OR2X1_LOC_515/Y 0.15fF
C11023 OR2X1_LOC_477/B OR2X1_LOC_477/Y 0.72fF
C11024 OR2X1_LOC_3/Y OR2X1_LOC_91/A 4.30fF
C11025 AND2X1_LOC_578/A AND2X1_LOC_851/a_8_24# 0.03fF
C11026 OR2X1_LOC_49/A OR2X1_LOC_95/Y 0.02fF
C11027 AND2X1_LOC_715/Y OR2X1_LOC_47/Y 0.09fF
C11028 AND2X1_LOC_568/a_8_24# OR2X1_LOC_91/A 0.08fF
C11029 AND2X1_LOC_392/A AND2X1_LOC_514/Y 0.07fF
C11030 VDD OR2X1_LOC_121/B 0.60fF
C11031 OR2X1_LOC_527/Y OR2X1_LOC_56/A 0.03fF
C11032 OR2X1_LOC_139/A OR2X1_LOC_223/A 0.03fF
C11033 OR2X1_LOC_18/Y OR2X1_LOC_95/a_8_216# 0.02fF
C11034 OR2X1_LOC_36/Y AND2X1_LOC_520/Y 0.28fF
C11035 AND2X1_LOC_572/A AND2X1_LOC_573/A 0.06fF
C11036 AND2X1_LOC_561/B OR2X1_LOC_64/Y 0.02fF
C11037 AND2X1_LOC_719/Y OR2X1_LOC_226/a_8_216# 0.16fF
C11038 OR2X1_LOC_70/Y AND2X1_LOC_436/a_8_24# 0.01fF
C11039 OR2X1_LOC_643/A OR2X1_LOC_523/Y 0.01fF
C11040 AND2X1_LOC_12/Y OR2X1_LOC_664/Y 0.09fF
C11041 OR2X1_LOC_74/A OR2X1_LOC_275/Y 0.06fF
C11042 INPUT_3 OR2X1_LOC_85/A 0.10fF
C11043 OR2X1_LOC_619/Y OR2X1_LOC_6/A 0.03fF
C11044 AND2X1_LOC_798/A OR2X1_LOC_428/A 0.07fF
C11045 AND2X1_LOC_543/a_36_24# OR2X1_LOC_74/A 0.00fF
C11046 OR2X1_LOC_83/a_8_216# OR2X1_LOC_394/a_8_216# 0.47fF
C11047 OR2X1_LOC_603/a_8_216# AND2X1_LOC_449/Y 0.00fF
C11048 INPUT_5 OR2X1_LOC_429/Y 0.02fF
C11049 OR2X1_LOC_114/Y AND2X1_LOC_95/Y 0.01fF
C11050 OR2X1_LOC_405/a_36_216# OR2X1_LOC_358/B 0.00fF
C11051 D_INPUT_0 AND2X1_LOC_243/Y 0.16fF
C11052 OR2X1_LOC_673/Y AND2X1_LOC_104/a_8_24# 0.28fF
C11053 OR2X1_LOC_791/B OR2X1_LOC_285/A 0.01fF
C11054 OR2X1_LOC_624/Y AND2X1_LOC_51/Y 0.03fF
C11055 VDD AND2X1_LOC_629/Y 0.01fF
C11056 AND2X1_LOC_866/B OR2X1_LOC_74/A 0.04fF
C11057 OR2X1_LOC_311/Y OR2X1_LOC_56/A 0.06fF
C11058 OR2X1_LOC_92/Y AND2X1_LOC_116/Y 0.05fF
C11059 OR2X1_LOC_269/a_8_216# OR2X1_LOC_269/B 0.04fF
C11060 AND2X1_LOC_721/Y AND2X1_LOC_795/Y 0.00fF
C11061 AND2X1_LOC_141/B AND2X1_LOC_141/A 0.14fF
C11062 OR2X1_LOC_702/A AND2X1_LOC_173/a_8_24# 0.02fF
C11063 AND2X1_LOC_64/Y OR2X1_LOC_608/Y 0.04fF
C11064 AND2X1_LOC_538/Y OR2X1_LOC_56/A 0.09fF
C11065 AND2X1_LOC_746/a_8_24# OR2X1_LOC_375/A 0.00fF
C11066 OR2X1_LOC_450/a_8_216# OR2X1_LOC_707/B 0.47fF
C11067 OR2X1_LOC_413/Y OR2X1_LOC_690/A 0.09fF
C11068 OR2X1_LOC_504/Y AND2X1_LOC_807/B 0.01fF
C11069 OR2X1_LOC_849/a_8_216# OR2X1_LOC_624/Y 0.01fF
C11070 OR2X1_LOC_844/Y OR2X1_LOC_658/a_36_216# 0.00fF
C11071 AND2X1_LOC_650/Y OR2X1_LOC_265/Y 0.02fF
C11072 OR2X1_LOC_473/A OR2X1_LOC_549/A 0.03fF
C11073 OR2X1_LOC_299/a_8_216# OR2X1_LOC_619/Y 0.01fF
C11074 OR2X1_LOC_189/A OR2X1_LOC_498/a_8_216# 0.01fF
C11075 OR2X1_LOC_115/a_8_216# AND2X1_LOC_3/Y 0.01fF
C11076 OR2X1_LOC_247/a_8_216# OR2X1_LOC_161/B 0.01fF
C11077 AND2X1_LOC_624/A OR2X1_LOC_52/B 0.06fF
C11078 OR2X1_LOC_328/a_8_216# AND2X1_LOC_639/A 0.09fF
C11079 OR2X1_LOC_312/Y OR2X1_LOC_315/Y 0.00fF
C11080 AND2X1_LOC_342/Y AND2X1_LOC_349/a_36_24# 0.01fF
C11081 OR2X1_LOC_215/A OR2X1_LOC_475/B 0.05fF
C11082 VDD OR2X1_LOC_75/a_8_216# 0.21fF
C11083 AND2X1_LOC_546/a_8_24# OR2X1_LOC_680/Y 0.23fF
C11084 OR2X1_LOC_32/a_36_216# OR2X1_LOC_39/A 0.00fF
C11085 AND2X1_LOC_89/a_8_24# OR2X1_LOC_97/B 0.02fF
C11086 AND2X1_LOC_86/B OR2X1_LOC_402/Y 0.15fF
C11087 AND2X1_LOC_561/B OR2X1_LOC_417/A 0.05fF
C11088 AND2X1_LOC_175/a_8_24# OR2X1_LOC_265/Y 0.01fF
C11089 OR2X1_LOC_43/Y OR2X1_LOC_41/Y 0.23fF
C11090 OR2X1_LOC_287/B OR2X1_LOC_375/A 0.03fF
C11091 OR2X1_LOC_70/Y AND2X1_LOC_354/Y 0.00fF
C11092 OR2X1_LOC_744/A OR2X1_LOC_71/Y 0.12fF
C11093 OR2X1_LOC_3/Y AND2X1_LOC_573/A 0.09fF
C11094 OR2X1_LOC_624/A AND2X1_LOC_42/B 0.05fF
C11095 AND2X1_LOC_728/a_8_24# OR2X1_LOC_679/B 0.09fF
C11096 OR2X1_LOC_624/B OR2X1_LOC_402/Y 0.07fF
C11097 OR2X1_LOC_65/B AND2X1_LOC_116/Y 0.01fF
C11098 OR2X1_LOC_155/A OR2X1_LOC_798/a_36_216# 0.02fF
C11099 OR2X1_LOC_662/A OR2X1_LOC_33/B 0.81fF
C11100 OR2X1_LOC_743/A OR2X1_LOC_316/Y 0.03fF
C11101 AND2X1_LOC_576/Y AND2X1_LOC_474/Y 0.07fF
C11102 OR2X1_LOC_246/Y OR2X1_LOC_485/A 0.26fF
C11103 OR2X1_LOC_151/A OR2X1_LOC_66/Y 0.03fF
C11104 AND2X1_LOC_158/a_8_24# OR2X1_LOC_210/B 0.01fF
C11105 OR2X1_LOC_436/Y OR2X1_LOC_78/B 0.04fF
C11106 D_INPUT_3 OR2X1_LOC_56/A 0.10fF
C11107 OR2X1_LOC_673/Y AND2X1_LOC_3/Y 0.03fF
C11108 OR2X1_LOC_699/a_36_216# OR2X1_LOC_89/A 0.00fF
C11109 AND2X1_LOC_576/Y OR2X1_LOC_485/A 0.09fF
C11110 OR2X1_LOC_145/Y AND2X1_LOC_663/A 0.38fF
C11111 OR2X1_LOC_97/a_8_216# OR2X1_LOC_375/A 0.01fF
C11112 AND2X1_LOC_522/a_8_24# OR2X1_LOC_560/A 0.21fF
C11113 OR2X1_LOC_263/a_36_216# OR2X1_LOC_92/Y 0.00fF
C11114 OR2X1_LOC_755/A AND2X1_LOC_624/A 0.05fF
C11115 AND2X1_LOC_179/a_8_24# OR2X1_LOC_223/A 0.01fF
C11116 OR2X1_LOC_18/Y OR2X1_LOC_19/B 0.89fF
C11117 OR2X1_LOC_43/A OR2X1_LOC_74/A 0.17fF
C11118 AND2X1_LOC_637/Y AND2X1_LOC_638/a_36_24# 0.00fF
C11119 OR2X1_LOC_578/a_8_216# OR2X1_LOC_578/B 0.02fF
C11120 OR2X1_LOC_51/Y AND2X1_LOC_675/a_36_24# 0.00fF
C11121 AND2X1_LOC_227/Y AND2X1_LOC_139/a_8_24# 0.01fF
C11122 OR2X1_LOC_113/A OR2X1_LOC_523/Y 0.28fF
C11123 OR2X1_LOC_76/A OR2X1_LOC_375/A 0.03fF
C11124 AND2X1_LOC_59/Y OR2X1_LOC_19/B 3.84fF
C11125 AND2X1_LOC_554/B AND2X1_LOC_123/a_8_24# 0.17fF
C11126 OR2X1_LOC_744/A D_INPUT_1 0.02fF
C11127 AND2X1_LOC_470/a_8_24# AND2X1_LOC_452/Y 0.02fF
C11128 OR2X1_LOC_856/A OR2X1_LOC_198/A 1.07fF
C11129 OR2X1_LOC_64/Y AND2X1_LOC_266/Y 0.13fF
C11130 AND2X1_LOC_116/B OR2X1_LOC_39/A 0.01fF
C11131 OR2X1_LOC_195/A AND2X1_LOC_3/Y 0.01fF
C11132 OR2X1_LOC_316/Y OR2X1_LOC_246/A 0.03fF
C11133 AND2X1_LOC_95/Y OR2X1_LOC_286/a_8_216# 0.01fF
C11134 OR2X1_LOC_36/Y AND2X1_LOC_856/B 0.26fF
C11135 OR2X1_LOC_43/A OR2X1_LOC_261/A 0.00fF
C11136 AND2X1_LOC_853/a_8_24# OR2X1_LOC_52/B 0.06fF
C11137 AND2X1_LOC_12/Y AND2X1_LOC_494/a_36_24# 0.01fF
C11138 OR2X1_LOC_675/A OR2X1_LOC_722/a_8_216# 0.01fF
C11139 AND2X1_LOC_663/B OR2X1_LOC_701/a_36_216# 0.00fF
C11140 OR2X1_LOC_36/Y AND2X1_LOC_863/A 0.11fF
C11141 OR2X1_LOC_629/A OR2X1_LOC_629/a_8_216# 0.51fF
C11142 AND2X1_LOC_390/B OR2X1_LOC_743/A 0.07fF
C11143 OR2X1_LOC_834/A OR2X1_LOC_512/a_8_216# -0.00fF
C11144 OR2X1_LOC_95/Y AND2X1_LOC_805/Y 0.02fF
C11145 OR2X1_LOC_835/Y OR2X1_LOC_375/A 0.16fF
C11146 OR2X1_LOC_615/a_8_216# OR2X1_LOC_7/A 0.03fF
C11147 OR2X1_LOC_148/A OR2X1_LOC_375/A 0.03fF
C11148 AND2X1_LOC_727/A AND2X1_LOC_661/A 0.03fF
C11149 OR2X1_LOC_26/Y OR2X1_LOC_245/a_8_216# 0.11fF
C11150 OR2X1_LOC_412/a_8_216# OR2X1_LOC_85/A 0.05fF
C11151 AND2X1_LOC_56/a_8_24# AND2X1_LOC_43/B 0.04fF
C11152 OR2X1_LOC_649/B OR2X1_LOC_649/a_8_216# 0.06fF
C11153 AND2X1_LOC_67/a_8_24# OR2X1_LOC_66/Y 0.11fF
C11154 OR2X1_LOC_695/a_8_216# OR2X1_LOC_47/Y 0.06fF
C11155 AND2X1_LOC_91/B OR2X1_LOC_714/a_8_216# 0.01fF
C11156 D_INPUT_3 AND2X1_LOC_9/a_8_24# 0.01fF
C11157 AND2X1_LOC_794/B OR2X1_LOC_13/B 0.01fF
C11158 AND2X1_LOC_334/a_8_24# AND2X1_LOC_640/Y 0.01fF
C11159 OR2X1_LOC_76/A OR2X1_LOC_605/B 1.93fF
C11160 OR2X1_LOC_497/a_8_216# AND2X1_LOC_227/Y 0.01fF
C11161 AND2X1_LOC_434/a_8_24# OR2X1_LOC_172/Y 0.04fF
C11162 OR2X1_LOC_562/Y OR2X1_LOC_570/A 0.06fF
C11163 OR2X1_LOC_633/A AND2X1_LOC_36/Y 0.03fF
C11164 OR2X1_LOC_264/Y OR2X1_LOC_598/A 0.01fF
C11165 AND2X1_LOC_42/B OR2X1_LOC_54/Y 0.03fF
C11166 OR2X1_LOC_643/A AND2X1_LOC_47/Y 0.03fF
C11167 OR2X1_LOC_115/B OR2X1_LOC_554/a_8_216# 0.18fF
C11168 OR2X1_LOC_523/B OR2X1_LOC_523/A 0.16fF
C11169 AND2X1_LOC_859/B AND2X1_LOC_806/A 0.01fF
C11170 AND2X1_LOC_47/Y OR2X1_LOC_778/Y 0.12fF
C11171 AND2X1_LOC_834/a_8_24# AND2X1_LOC_796/Y 0.01fF
C11172 AND2X1_LOC_56/B D_INPUT_3 0.04fF
C11173 OR2X1_LOC_756/B AND2X1_LOC_31/Y 0.16fF
C11174 OR2X1_LOC_736/A OR2X1_LOC_736/a_8_216# 0.04fF
C11175 OR2X1_LOC_8/Y OR2X1_LOC_150/a_8_216# 0.01fF
C11176 OR2X1_LOC_246/Y OR2X1_LOC_10/a_8_216# 0.06fF
C11177 AND2X1_LOC_387/B AND2X1_LOC_7/Y 0.12fF
C11178 OR2X1_LOC_427/A OR2X1_LOC_406/A -0.04fF
C11179 VDD OR2X1_LOC_13/B 0.79fF
C11180 AND2X1_LOC_40/Y OR2X1_LOC_398/Y 0.03fF
C11181 AND2X1_LOC_8/Y D_INPUT_3 0.02fF
C11182 AND2X1_LOC_512/Y OR2X1_LOC_533/A 0.01fF
C11183 OR2X1_LOC_244/Y OR2X1_LOC_140/Y 0.01fF
C11184 OR2X1_LOC_6/B AND2X1_LOC_750/a_8_24# -0.03fF
C11185 OR2X1_LOC_70/Y AND2X1_LOC_635/a_36_24# -0.00fF
C11186 AND2X1_LOC_334/a_8_24# OR2X1_LOC_416/Y 0.01fF
C11187 OR2X1_LOC_39/A AND2X1_LOC_204/Y 0.00fF
C11188 VDD OR2X1_LOC_195/a_8_216# 0.21fF
C11189 OR2X1_LOC_647/A AND2X1_LOC_47/Y 0.08fF
C11190 AND2X1_LOC_359/a_8_24# OR2X1_LOC_47/Y 0.02fF
C11191 AND2X1_LOC_534/a_8_24# OR2X1_LOC_356/B -0.01fF
C11192 OR2X1_LOC_185/A OR2X1_LOC_192/a_8_216# 0.05fF
C11193 OR2X1_LOC_447/Y OR2X1_LOC_705/Y 0.09fF
C11194 AND2X1_LOC_70/Y OR2X1_LOC_217/A 0.00fF
C11195 OR2X1_LOC_234/a_8_216# OR2X1_LOC_753/A 0.03fF
C11196 OR2X1_LOC_392/B OR2X1_LOC_576/A 0.03fF
C11197 OR2X1_LOC_750/A OR2X1_LOC_814/A 0.09fF
C11198 D_INPUT_3 OR2X1_LOC_291/A 0.00fF
C11199 OR2X1_LOC_45/B AND2X1_LOC_339/Y 0.01fF
C11200 OR2X1_LOC_22/Y INPUT_1 3.08fF
C11201 AND2X1_LOC_110/Y OR2X1_LOC_356/B 0.01fF
C11202 OR2X1_LOC_696/A AND2X1_LOC_732/B 0.01fF
C11203 AND2X1_LOC_573/A AND2X1_LOC_772/a_8_24# 0.01fF
C11204 OR2X1_LOC_643/A OR2X1_LOC_598/A 0.07fF
C11205 AND2X1_LOC_335/a_36_24# OR2X1_LOC_437/A 0.00fF
C11206 OR2X1_LOC_43/A AND2X1_LOC_647/Y 0.03fF
C11207 OR2X1_LOC_124/Y OR2X1_LOC_598/A 0.03fF
C11208 OR2X1_LOC_355/A OR2X1_LOC_355/a_8_216# 0.47fF
C11209 AND2X1_LOC_711/A AND2X1_LOC_792/a_8_24# 0.05fF
C11210 AND2X1_LOC_797/A OR2X1_LOC_47/Y 0.03fF
C11211 AND2X1_LOC_712/a_8_24# OR2X1_LOC_12/Y 0.02fF
C11212 OR2X1_LOC_158/A AND2X1_LOC_284/a_8_24# 0.04fF
C11213 AND2X1_LOC_91/B OR2X1_LOC_6/B 0.11fF
C11214 OR2X1_LOC_472/A OR2X1_LOC_598/A 0.03fF
C11215 AND2X1_LOC_727/A AND2X1_LOC_810/Y 0.01fF
C11216 OR2X1_LOC_111/a_8_216# VDD 0.21fF
C11217 OR2X1_LOC_473/Y OR2X1_LOC_786/Y 0.41fF
C11218 AND2X1_LOC_663/B OR2X1_LOC_47/Y 0.03fF
C11219 OR2X1_LOC_323/a_8_216# OR2X1_LOC_323/Y 0.02fF
C11220 AND2X1_LOC_726/Y AND2X1_LOC_731/Y 0.02fF
C11221 AND2X1_LOC_47/Y OR2X1_LOC_113/A 0.00fF
C11222 OR2X1_LOC_576/A OR2X1_LOC_113/B 0.03fF
C11223 OR2X1_LOC_262/a_8_216# OR2X1_LOC_72/Y 0.01fF
C11224 OR2X1_LOC_400/a_8_216# OR2X1_LOC_771/B 0.06fF
C11225 OR2X1_LOC_629/B OR2X1_LOC_563/A 0.01fF
C11226 OR2X1_LOC_215/Y AND2X1_LOC_406/a_36_24# 0.00fF
C11227 OR2X1_LOC_481/A OR2X1_LOC_257/Y 0.01fF
C11228 AND2X1_LOC_574/Y AND2X1_LOC_500/Y 0.24fF
C11229 OR2X1_LOC_829/a_8_216# OR2X1_LOC_13/B 0.04fF
C11230 AND2X1_LOC_462/B OR2X1_LOC_27/Y 0.21fF
C11231 OR2X1_LOC_362/B OR2X1_LOC_580/A 0.01fF
C11232 OR2X1_LOC_858/A OR2X1_LOC_140/B 0.03fF
C11233 AND2X1_LOC_640/a_8_24# AND2X1_LOC_476/A 0.03fF
C11234 AND2X1_LOC_753/a_8_24# AND2X1_LOC_41/Y 0.01fF
C11235 AND2X1_LOC_476/Y OR2X1_LOC_373/Y 0.05fF
C11236 OR2X1_LOC_97/A OR2X1_LOC_832/a_36_216# 0.00fF
C11237 OR2X1_LOC_575/A OR2X1_LOC_844/B 0.00fF
C11238 OR2X1_LOC_857/A VDD 0.00fF
C11239 OR2X1_LOC_125/a_8_216# OR2X1_LOC_428/A 0.01fF
C11240 AND2X1_LOC_810/Y OR2X1_LOC_95/Y 0.02fF
C11241 OR2X1_LOC_97/A AND2X1_LOC_172/a_8_24# 0.01fF
C11242 OR2X1_LOC_200/a_8_216# OR2X1_LOC_193/a_8_216# 0.47fF
C11243 AND2X1_LOC_463/B OR2X1_LOC_22/A 0.26fF
C11244 OR2X1_LOC_47/Y OR2X1_LOC_54/a_8_216# 0.06fF
C11245 OR2X1_LOC_58/Y OR2X1_LOC_16/A 0.03fF
C11246 OR2X1_LOC_158/A AND2X1_LOC_566/B 0.03fF
C11247 OR2X1_LOC_786/a_36_216# OR2X1_LOC_549/A 0.00fF
C11248 OR2X1_LOC_426/B AND2X1_LOC_639/B 0.14fF
C11249 OR2X1_LOC_586/Y OR2X1_LOC_387/A 0.01fF
C11250 AND2X1_LOC_632/A AND2X1_LOC_623/a_8_24# 0.01fF
C11251 OR2X1_LOC_95/Y OR2X1_LOC_760/Y 0.04fF
C11252 AND2X1_LOC_476/A AND2X1_LOC_649/Y 0.05fF
C11253 OR2X1_LOC_154/A OR2X1_LOC_537/a_8_216# 0.03fF
C11254 OR2X1_LOC_18/Y OR2X1_LOC_504/a_8_216# 0.01fF
C11255 OR2X1_LOC_194/Y AND2X1_LOC_41/Y 0.08fF
C11256 VDD AND2X1_LOC_199/A 0.25fF
C11257 OR2X1_LOC_479/Y OR2X1_LOC_353/a_36_216# 0.02fF
C11258 AND2X1_LOC_476/A AND2X1_LOC_293/a_36_24# 0.00fF
C11259 AND2X1_LOC_41/A OR2X1_LOC_392/B 0.03fF
C11260 AND2X1_LOC_67/Y OR2X1_LOC_68/B 0.00fF
C11261 OR2X1_LOC_696/A OR2X1_LOC_625/Y 0.07fF
C11262 OR2X1_LOC_251/Y OR2X1_LOC_13/B 0.07fF
C11263 AND2X1_LOC_70/Y AND2X1_LOC_40/a_8_24# 0.01fF
C11264 AND2X1_LOC_222/a_8_24# AND2X1_LOC_786/Y 0.05fF
C11265 OR2X1_LOC_507/B OR2X1_LOC_510/a_8_216# 0.49fF
C11266 AND2X1_LOC_861/B OR2X1_LOC_816/A 0.80fF
C11267 AND2X1_LOC_588/B OR2X1_LOC_502/A 0.05fF
C11268 OR2X1_LOC_474/Y OR2X1_LOC_474/B 0.03fF
C11269 OR2X1_LOC_508/A OR2X1_LOC_392/B 0.10fF
C11270 AND2X1_LOC_677/a_8_24# AND2X1_LOC_31/Y 0.01fF
C11271 AND2X1_LOC_498/a_8_24# OR2X1_LOC_549/A 0.01fF
C11272 AND2X1_LOC_3/Y OR2X1_LOC_769/a_8_216# 0.01fF
C11273 OR2X1_LOC_227/a_8_216# AND2X1_LOC_31/Y 0.01fF
C11274 OR2X1_LOC_139/A OR2X1_LOC_502/A 0.07fF
C11275 AND2X1_LOC_753/B AND2X1_LOC_7/B 0.04fF
C11276 OR2X1_LOC_323/A OR2X1_LOC_18/Y 0.05fF
C11277 OR2X1_LOC_492/Y OR2X1_LOC_744/A 0.04fF
C11278 OR2X1_LOC_309/Y OR2X1_LOC_426/B 0.01fF
C11279 OR2X1_LOC_45/B OR2X1_LOC_92/Y 0.96fF
C11280 OR2X1_LOC_509/a_8_216# OR2X1_LOC_78/A 0.01fF
C11281 OR2X1_LOC_18/Y OR2X1_LOC_89/Y 0.09fF
C11282 AND2X1_LOC_719/Y AND2X1_LOC_663/A 0.52fF
C11283 AND2X1_LOC_64/Y OR2X1_LOC_738/A 0.03fF
C11284 AND2X1_LOC_91/B OR2X1_LOC_732/a_36_216# 0.03fF
C11285 OR2X1_LOC_108/a_8_216# OR2X1_LOC_744/A 0.03fF
C11286 OR2X1_LOC_156/a_8_216# OR2X1_LOC_160/A 0.02fF
C11287 OR2X1_LOC_516/Y OR2X1_LOC_26/Y 0.03fF
C11288 AND2X1_LOC_306/a_8_24# OR2X1_LOC_307/A 0.01fF
C11289 OR2X1_LOC_405/A AND2X1_LOC_7/B 0.10fF
C11290 OR2X1_LOC_611/a_8_216# OR2X1_LOC_71/A 0.02fF
C11291 OR2X1_LOC_379/Y AND2X1_LOC_22/Y 0.03fF
C11292 OR2X1_LOC_375/A OR2X1_LOC_722/B 0.01fF
C11293 OR2X1_LOC_348/a_8_216# AND2X1_LOC_40/Y 0.05fF
C11294 OR2X1_LOC_646/a_8_216# AND2X1_LOC_36/Y 0.04fF
C11295 OR2X1_LOC_318/Y AND2X1_LOC_433/a_8_24# 0.02fF
C11296 OR2X1_LOC_160/B OR2X1_LOC_78/B 0.38fF
C11297 AND2X1_LOC_738/B AND2X1_LOC_330/a_8_24# 0.01fF
C11298 OR2X1_LOC_78/A OR2X1_LOC_66/A 0.55fF
C11299 AND2X1_LOC_547/Y OR2X1_LOC_524/Y 0.06fF
C11300 AND2X1_LOC_91/B OR2X1_LOC_579/B 0.40fF
C11301 OR2X1_LOC_214/B OR2X1_LOC_644/A 0.03fF
C11302 OR2X1_LOC_516/Y OR2X1_LOC_89/A 0.03fF
C11303 OR2X1_LOC_329/B AND2X1_LOC_112/a_36_24# 0.01fF
C11304 OR2X1_LOC_744/A OR2X1_LOC_426/B 0.17fF
C11305 OR2X1_LOC_175/Y OR2X1_LOC_798/a_8_216# 0.04fF
C11306 OR2X1_LOC_494/Y AND2X1_LOC_474/A 0.05fF
C11307 AND2X1_LOC_775/a_36_24# OR2X1_LOC_89/A 0.00fF
C11308 OR2X1_LOC_45/B OR2X1_LOC_65/B 0.13fF
C11309 OR2X1_LOC_497/Y AND2X1_LOC_227/a_8_24# 0.01fF
C11310 AND2X1_LOC_571/B OR2X1_LOC_89/A 0.01fF
C11311 OR2X1_LOC_379/Y OR2X1_LOC_855/a_36_216# 0.00fF
C11312 AND2X1_LOC_12/Y OR2X1_LOC_61/A 0.02fF
C11313 AND2X1_LOC_468/B AND2X1_LOC_212/Y 0.07fF
C11314 OR2X1_LOC_589/A OR2X1_LOC_432/a_8_216# 0.03fF
C11315 OR2X1_LOC_691/B OR2X1_LOC_377/A 0.00fF
C11316 OR2X1_LOC_154/A AND2X1_LOC_60/a_8_24# 0.04fF
C11317 AND2X1_LOC_218/Y AND2X1_LOC_222/a_8_24# 0.11fF
C11318 AND2X1_LOC_810/A AND2X1_LOC_365/A 0.03fF
C11319 OR2X1_LOC_329/B AND2X1_LOC_858/B 0.09fF
C11320 OR2X1_LOC_604/A OR2X1_LOC_683/a_36_216# 0.00fF
C11321 OR2X1_LOC_121/a_36_216# OR2X1_LOC_375/A 0.00fF
C11322 OR2X1_LOC_329/B OR2X1_LOC_91/A 0.07fF
C11323 OR2X1_LOC_703/B OR2X1_LOC_161/B 0.04fF
C11324 AND2X1_LOC_22/Y OR2X1_LOC_114/Y 0.03fF
C11325 OR2X1_LOC_175/Y OR2X1_LOC_269/B 0.10fF
C11326 AND2X1_LOC_866/B OR2X1_LOC_626/Y 0.19fF
C11327 AND2X1_LOC_59/Y AND2X1_LOC_534/a_8_24# 0.03fF
C11328 AND2X1_LOC_539/Y AND2X1_LOC_355/a_8_24# 0.18fF
C11329 OR2X1_LOC_494/a_8_216# OR2X1_LOC_56/A 0.05fF
C11330 OR2X1_LOC_468/Y AND2X1_LOC_44/Y 0.02fF
C11331 OR2X1_LOC_448/B OR2X1_LOC_66/A 0.02fF
C11332 AND2X1_LOC_303/A OR2X1_LOC_16/A 0.06fF
C11333 OR2X1_LOC_697/Y OR2X1_LOC_743/a_36_216# 0.00fF
C11334 OR2X1_LOC_45/B OR2X1_LOC_271/Y 0.01fF
C11335 OR2X1_LOC_87/A OR2X1_LOC_161/B 0.16fF
C11336 OR2X1_LOC_26/Y OR2X1_LOC_373/a_8_216# 0.04fF
C11337 AND2X1_LOC_641/Y OR2X1_LOC_171/Y 0.13fF
C11338 OR2X1_LOC_254/B OR2X1_LOC_486/Y 0.26fF
C11339 OR2X1_LOC_139/A OR2X1_LOC_137/Y 0.07fF
C11340 OR2X1_LOC_147/A AND2X1_LOC_41/A 0.15fF
C11341 OR2X1_LOC_682/a_8_216# OR2X1_LOC_428/A 0.05fF
C11342 VDD OR2X1_LOC_856/B 0.27fF
C11343 OR2X1_LOC_256/A OR2X1_LOC_13/B 0.04fF
C11344 OR2X1_LOC_691/Y OR2X1_LOC_269/B 0.03fF
C11345 OR2X1_LOC_691/a_8_216# OR2X1_LOC_835/B 0.02fF
C11346 OR2X1_LOC_510/A OR2X1_LOC_507/B 0.36fF
C11347 AND2X1_LOC_486/Y OR2X1_LOC_666/A 0.03fF
C11348 OR2X1_LOC_692/Y OR2X1_LOC_44/Y 0.14fF
C11349 OR2X1_LOC_715/B AND2X1_LOC_43/B 0.00fF
C11350 AND2X1_LOC_810/A OR2X1_LOC_43/A 0.03fF
C11351 OR2X1_LOC_8/Y AND2X1_LOC_62/a_8_24# 0.01fF
C11352 AND2X1_LOC_778/a_8_24# AND2X1_LOC_786/Y 0.02fF
C11353 OR2X1_LOC_496/Y AND2X1_LOC_795/a_8_24# 0.01fF
C11354 OR2X1_LOC_689/a_36_216# OR2X1_LOC_690/Y 0.00fF
C11355 OR2X1_LOC_89/A OR2X1_LOC_373/a_8_216# 0.01fF
C11356 OR2X1_LOC_493/a_8_216# OR2X1_LOC_493/A 0.01fF
C11357 OR2X1_LOC_52/B AND2X1_LOC_774/A 0.42fF
C11358 OR2X1_LOC_269/B OR2X1_LOC_713/A 0.09fF
C11359 AND2X1_LOC_59/Y AND2X1_LOC_110/Y 0.03fF
C11360 OR2X1_LOC_502/A OR2X1_LOC_637/Y 0.03fF
C11361 VDD OR2X1_LOC_679/B 0.21fF
C11362 OR2X1_LOC_485/A AND2X1_LOC_244/A 0.04fF
C11363 VDD OR2X1_LOC_793/a_8_216# 0.00fF
C11364 OR2X1_LOC_604/A AND2X1_LOC_848/Y 0.20fF
C11365 OR2X1_LOC_510/Y AND2X1_LOC_625/a_36_24# 0.00fF
C11366 OR2X1_LOC_532/B OR2X1_LOC_523/a_8_216# 0.01fF
C11367 AND2X1_LOC_70/Y OR2X1_LOC_185/A 0.10fF
C11368 AND2X1_LOC_719/Y OR2X1_LOC_283/a_8_216# 0.04fF
C11369 OR2X1_LOC_287/B OR2X1_LOC_843/B 0.27fF
C11370 AND2X1_LOC_500/Y AND2X1_LOC_621/Y 0.03fF
C11371 OR2X1_LOC_160/B OR2X1_LOC_375/A 3.67fF
C11372 AND2X1_LOC_17/Y AND2X1_LOC_40/a_8_24# 0.01fF
C11373 OR2X1_LOC_181/B OR2X1_LOC_742/a_8_216# 0.01fF
C11374 OR2X1_LOC_371/Y AND2X1_LOC_785/Y 0.33fF
C11375 OR2X1_LOC_51/Y AND2X1_LOC_452/Y 0.01fF
C11376 AND2X1_LOC_86/Y OR2X1_LOC_78/B 0.32fF
C11377 OR2X1_LOC_485/A OR2X1_LOC_16/A 0.07fF
C11378 OR2X1_LOC_813/a_8_216# OR2X1_LOC_235/a_8_216# 0.47fF
C11379 OR2X1_LOC_528/Y AND2X1_LOC_859/Y 0.14fF
C11380 AND2X1_LOC_337/B AND2X1_LOC_810/B 0.03fF
C11381 OR2X1_LOC_482/a_8_216# OR2X1_LOC_7/A 0.09fF
C11382 OR2X1_LOC_131/Y OR2X1_LOC_595/A 0.01fF
C11383 OR2X1_LOC_440/A OR2X1_LOC_180/B 0.00fF
C11384 AND2X1_LOC_12/Y AND2X1_LOC_24/a_8_24# 0.01fF
C11385 OR2X1_LOC_475/a_8_216# OR2X1_LOC_475/B 0.03fF
C11386 OR2X1_LOC_151/A OR2X1_LOC_574/A 0.09fF
C11387 OR2X1_LOC_600/A OR2X1_LOC_44/Y 2.13fF
C11388 OR2X1_LOC_252/Y AND2X1_LOC_663/A 0.03fF
C11389 AND2X1_LOC_1/Y AND2X1_LOC_44/Y 0.04fF
C11390 OR2X1_LOC_67/Y OR2X1_LOC_13/B 0.07fF
C11391 OR2X1_LOC_228/Y OR2X1_LOC_341/a_36_216# 0.03fF
C11392 AND2X1_LOC_550/A OR2X1_LOC_677/a_8_216# 0.47fF
C11393 OR2X1_LOC_230/a_8_216# OR2X1_LOC_12/Y 0.01fF
C11394 OR2X1_LOC_78/B OR2X1_LOC_799/a_8_216# 0.01fF
C11395 OR2X1_LOC_114/a_8_216# OR2X1_LOC_161/A 0.01fF
C11396 OR2X1_LOC_720/a_8_216# AND2X1_LOC_18/Y 0.01fF
C11397 AND2X1_LOC_91/B OR2X1_LOC_68/Y 0.19fF
C11398 OR2X1_LOC_185/A OR2X1_LOC_703/A 0.06fF
C11399 AND2X1_LOC_561/a_8_24# AND2X1_LOC_866/A 0.04fF
C11400 OR2X1_LOC_599/A AND2X1_LOC_658/A 0.03fF
C11401 OR2X1_LOC_647/A OR2X1_LOC_646/B 0.67fF
C11402 AND2X1_LOC_729/Y OR2X1_LOC_524/Y 0.03fF
C11403 OR2X1_LOC_166/a_8_216# OR2X1_LOC_44/Y 0.05fF
C11404 OR2X1_LOC_405/A OR2X1_LOC_319/B 0.09fF
C11405 AND2X1_LOC_168/Y AND2X1_LOC_168/a_8_24# 0.01fF
C11406 OR2X1_LOC_123/B AND2X1_LOC_65/A 0.04fF
C11407 AND2X1_LOC_861/B AND2X1_LOC_807/Y 0.00fF
C11408 AND2X1_LOC_532/a_8_24# OR2X1_LOC_594/Y 0.25fF
C11409 OR2X1_LOC_132/a_8_216# AND2X1_LOC_361/A 0.01fF
C11410 AND2X1_LOC_136/a_8_24# OR2X1_LOC_596/A 0.01fF
C11411 AND2X1_LOC_203/a_8_24# AND2X1_LOC_215/a_8_24# 0.23fF
C11412 OR2X1_LOC_863/a_36_216# OR2X1_LOC_35/Y 0.00fF
C11413 OR2X1_LOC_656/B AND2X1_LOC_40/Y 0.08fF
C11414 AND2X1_LOC_296/a_8_24# OR2X1_LOC_44/Y 0.04fF
C11415 OR2X1_LOC_155/A OR2X1_LOC_66/A 0.03fF
C11416 AND2X1_LOC_705/Y OR2X1_LOC_64/Y 0.05fF
C11417 OR2X1_LOC_466/A OR2X1_LOC_449/a_8_216# 0.40fF
C11418 OR2X1_LOC_162/Y AND2X1_LOC_51/Y 0.10fF
C11419 AND2X1_LOC_711/a_8_24# OR2X1_LOC_44/Y 0.01fF
C11420 OR2X1_LOC_108/Y OR2X1_LOC_485/A 0.19fF
C11421 OR2X1_LOC_650/a_8_216# AND2X1_LOC_8/Y 0.04fF
C11422 OR2X1_LOC_56/A AND2X1_LOC_806/A 0.00fF
C11423 OR2X1_LOC_69/Y OR2X1_LOC_59/Y 0.02fF
C11424 OR2X1_LOC_841/A OR2X1_LOC_155/A 0.03fF
C11425 OR2X1_LOC_421/A AND2X1_LOC_639/a_8_24# 0.23fF
C11426 OR2X1_LOC_158/A OR2X1_LOC_488/a_36_216# 0.03fF
C11427 AND2X1_LOC_37/a_8_24# INPUT_2 0.09fF
C11428 AND2X1_LOC_206/Y AND2X1_LOC_215/a_8_24# 0.03fF
C11429 OR2X1_LOC_218/a_8_216# OR2X1_LOC_78/A 0.02fF
C11430 AND2X1_LOC_91/B AND2X1_LOC_47/Y 0.21fF
C11431 AND2X1_LOC_51/Y OR2X1_LOC_729/a_8_216# 0.02fF
C11432 OR2X1_LOC_588/Y OR2X1_LOC_25/Y 0.03fF
C11433 OR2X1_LOC_854/a_8_216# OR2X1_LOC_161/A 0.01fF
C11434 OR2X1_LOC_92/Y AND2X1_LOC_435/a_8_24# 0.28fF
C11435 OR2X1_LOC_174/A OR2X1_LOC_358/B 0.00fF
C11436 OR2X1_LOC_114/Y OR2X1_LOC_244/B 0.16fF
C11437 OR2X1_LOC_471/Y AND2X1_LOC_44/Y 0.03fF
C11438 OR2X1_LOC_160/A OR2X1_LOC_660/a_8_216# 0.01fF
C11439 AND2X1_LOC_737/Y AND2X1_LOC_624/A 0.03fF
C11440 OR2X1_LOC_309/a_8_216# OR2X1_LOC_64/Y 0.06fF
C11441 OR2X1_LOC_604/A OR2X1_LOC_617/Y 0.06fF
C11442 OR2X1_LOC_655/B AND2X1_LOC_44/Y 1.97fF
C11443 OR2X1_LOC_219/B OR2X1_LOC_78/B 0.08fF
C11444 OR2X1_LOC_339/a_36_216# OR2X1_LOC_333/B 0.00fF
C11445 OR2X1_LOC_575/A OR2X1_LOC_573/Y 0.12fF
C11446 OR2X1_LOC_532/B OR2X1_LOC_576/A 0.03fF
C11447 OR2X1_LOC_160/A AND2X1_LOC_492/a_8_24# 0.11fF
C11448 OR2X1_LOC_256/Y AND2X1_LOC_349/a_8_24# 0.04fF
C11449 AND2X1_LOC_562/B OR2X1_LOC_36/Y 0.03fF
C11450 AND2X1_LOC_456/B AND2X1_LOC_359/B 0.02fF
C11451 AND2X1_LOC_280/a_36_24# OR2X1_LOC_161/A 0.00fF
C11452 OR2X1_LOC_864/A OR2X1_LOC_756/B 0.11fF
C11453 OR2X1_LOC_847/A OR2X1_LOC_402/Y 0.07fF
C11454 OR2X1_LOC_687/Y AND2X1_LOC_615/a_8_24# 0.06fF
C11455 INPUT_5 AND2X1_LOC_30/a_8_24# 0.01fF
C11456 AND2X1_LOC_706/Y AND2X1_LOC_687/Y 0.17fF
C11457 OR2X1_LOC_769/B AND2X1_LOC_3/Y 0.00fF
C11458 D_INPUT_0 OR2X1_LOC_12/Y 2.67fF
C11459 OR2X1_LOC_637/a_36_216# OR2X1_LOC_828/B 0.00fF
C11460 AND2X1_LOC_276/Y OR2X1_LOC_56/A 0.06fF
C11461 OR2X1_LOC_744/A OR2X1_LOC_743/A 0.14fF
C11462 AND2X1_LOC_141/A OR2X1_LOC_26/Y 0.01fF
C11463 AND2X1_LOC_86/Y OR2X1_LOC_375/A 0.02fF
C11464 AND2X1_LOC_139/a_36_24# AND2X1_LOC_361/A 0.01fF
C11465 AND2X1_LOC_50/Y AND2X1_LOC_64/a_8_24# 0.04fF
C11466 AND2X1_LOC_553/A AND2X1_LOC_560/B 0.02fF
C11467 OR2X1_LOC_857/B D_INPUT_0 0.46fF
C11468 OR2X1_LOC_405/A OR2X1_LOC_805/A 1.63fF
C11469 OR2X1_LOC_377/A AND2X1_LOC_233/a_8_24# 0.02fF
C11470 OR2X1_LOC_87/A OR2X1_LOC_61/Y 0.63fF
C11471 AND2X1_LOC_714/a_8_24# OR2X1_LOC_31/Y 0.01fF
C11472 OR2X1_LOC_661/a_8_216# OR2X1_LOC_130/A 0.14fF
C11473 OR2X1_LOC_656/B OR2X1_LOC_87/Y 0.03fF
C11474 OR2X1_LOC_377/A OR2X1_LOC_404/a_36_216# 0.00fF
C11475 OR2X1_LOC_820/a_8_216# INPUT_1 0.01fF
C11476 OR2X1_LOC_179/a_8_216# OR2X1_LOC_529/Y 0.01fF
C11477 OR2X1_LOC_291/a_8_216# OR2X1_LOC_36/Y 0.10fF
C11478 OR2X1_LOC_837/A OR2X1_LOC_753/A 0.14fF
C11479 OR2X1_LOC_46/A OR2X1_LOC_461/B 0.03fF
C11480 AND2X1_LOC_64/Y AND2X1_LOC_72/B 0.04fF
C11481 AND2X1_LOC_516/a_8_24# OR2X1_LOC_623/B 0.03fF
C11482 AND2X1_LOC_141/A OR2X1_LOC_89/A 0.02fF
C11483 AND2X1_LOC_340/Y OR2X1_LOC_75/Y 0.01fF
C11484 OR2X1_LOC_47/Y OR2X1_LOC_18/a_8_216# 0.01fF
C11485 AND2X1_LOC_47/Y OR2X1_LOC_364/a_8_216# 0.01fF
C11486 OR2X1_LOC_364/A OR2X1_LOC_624/A 0.07fF
C11487 AND2X1_LOC_59/Y OR2X1_LOC_664/Y 0.19fF
C11488 VDD OR2X1_LOC_383/Y 0.20fF
C11489 OR2X1_LOC_185/Y OR2X1_LOC_624/A 0.07fF
C11490 OR2X1_LOC_831/B OR2X1_LOC_493/Y 0.07fF
C11491 OR2X1_LOC_619/Y OR2X1_LOC_44/Y 0.14fF
C11492 OR2X1_LOC_375/A OR2X1_LOC_553/A 0.07fF
C11493 AND2X1_LOC_145/a_8_24# OR2X1_LOC_148/B 0.01fF
C11494 AND2X1_LOC_850/Y AND2X1_LOC_806/A 0.01fF
C11495 OR2X1_LOC_671/Y OR2X1_LOC_95/Y 0.02fF
C11496 AND2X1_LOC_359/a_8_24# OR2X1_LOC_625/Y 0.04fF
C11497 OR2X1_LOC_756/B AND2X1_LOC_281/a_8_24# 0.00fF
C11498 AND2X1_LOC_95/Y OR2X1_LOC_849/A 0.02fF
C11499 OR2X1_LOC_585/A OR2X1_LOC_278/Y 0.04fF
C11500 AND2X1_LOC_584/a_8_24# OR2X1_LOC_639/B 0.04fF
C11501 OR2X1_LOC_462/B OR2X1_LOC_130/A 0.52fF
C11502 AND2X1_LOC_91/B OR2X1_LOC_598/A 0.10fF
C11503 OR2X1_LOC_87/A OR2X1_LOC_87/a_8_216# 0.05fF
C11504 AND2X1_LOC_99/A OR2X1_LOC_106/A 0.00fF
C11505 OR2X1_LOC_205/Y AND2X1_LOC_44/Y 0.02fF
C11506 OR2X1_LOC_6/B OR2X1_LOC_751/A 0.04fF
C11507 OR2X1_LOC_744/A OR2X1_LOC_246/A 0.02fF
C11508 AND2X1_LOC_70/Y OR2X1_LOC_750/a_36_216# 0.00fF
C11509 OR2X1_LOC_600/A OR2X1_LOC_80/a_36_216# 0.02fF
C11510 OR2X1_LOC_585/A OR2X1_LOC_38/a_8_216# 0.01fF
C11511 AND2X1_LOC_70/Y AND2X1_LOC_431/a_8_24# 0.09fF
C11512 AND2X1_LOC_255/a_8_24# OR2X1_LOC_241/B 0.06fF
C11513 OR2X1_LOC_625/Y OR2X1_LOC_754/a_36_216# 0.01fF
C11514 OR2X1_LOC_510/Y OR2X1_LOC_810/A 0.03fF
C11515 OR2X1_LOC_836/A AND2X1_LOC_823/a_8_24# 0.08fF
C11516 OR2X1_LOC_645/a_8_216# AND2X1_LOC_47/Y 0.01fF
C11517 AND2X1_LOC_78/a_8_24# OR2X1_LOC_18/Y 0.03fF
C11518 OR2X1_LOC_290/Y OR2X1_LOC_291/Y 0.05fF
C11519 AND2X1_LOC_553/A OR2X1_LOC_64/Y 0.00fF
C11520 OR2X1_LOC_6/A AND2X1_LOC_818/a_8_24# 0.01fF
C11521 OR2X1_LOC_426/B OR2X1_LOC_31/Y 0.13fF
C11522 OR2X1_LOC_280/a_8_216# OR2X1_LOC_237/Y 0.01fF
C11523 OR2X1_LOC_95/a_8_216# OR2X1_LOC_585/A 0.03fF
C11524 AND2X1_LOC_80/a_8_24# OR2X1_LOC_646/A 0.09fF
C11525 OR2X1_LOC_673/a_36_216# D_INPUT_1 0.00fF
C11526 AND2X1_LOC_831/Y OR2X1_LOC_56/A 0.07fF
C11527 OR2X1_LOC_244/A OR2X1_LOC_78/B 0.08fF
C11528 AND2X1_LOC_56/B OR2X1_LOC_83/A 0.03fF
C11529 OR2X1_LOC_465/B OR2X1_LOC_457/B 0.82fF
C11530 AND2X1_LOC_42/B OR2X1_LOC_161/A 0.06fF
C11531 OR2X1_LOC_22/Y OR2X1_LOC_517/A 0.20fF
C11532 AND2X1_LOC_658/A AND2X1_LOC_866/A 0.01fF
C11533 AND2X1_LOC_154/Y OR2X1_LOC_39/A 0.04fF
C11534 AND2X1_LOC_847/a_8_24# AND2X1_LOC_847/Y 0.02fF
C11535 OR2X1_LOC_3/Y OR2X1_LOC_32/B 0.03fF
C11536 OR2X1_LOC_252/a_8_216# OR2X1_LOC_617/Y 0.01fF
C11537 AND2X1_LOC_54/a_8_24# D_INPUT_0 0.02fF
C11538 AND2X1_LOC_392/A OR2X1_LOC_47/Y 0.03fF
C11539 AND2X1_LOC_41/A OR2X1_LOC_532/B 0.07fF
C11540 OR2X1_LOC_837/Y D_INPUT_0 0.18fF
C11541 AND2X1_LOC_565/B OR2X1_LOC_47/Y 0.01fF
C11542 OR2X1_LOC_154/A OR2X1_LOC_557/A 0.00fF
C11543 OR2X1_LOC_744/A OR2X1_LOC_409/B 0.83fF
C11544 AND2X1_LOC_472/B OR2X1_LOC_585/A 0.07fF
C11545 AND2X1_LOC_44/Y OR2X1_LOC_750/Y 0.68fF
C11546 OR2X1_LOC_521/Y OR2X1_LOC_22/Y 0.03fF
C11547 OR2X1_LOC_51/Y AND2X1_LOC_687/a_8_24# 0.01fF
C11548 AND2X1_LOC_861/B OR2X1_LOC_95/Y 0.07fF
C11549 OR2X1_LOC_829/Y AND2X1_LOC_655/A 0.14fF
C11550 OR2X1_LOC_676/Y AND2X1_LOC_39/Y 0.01fF
C11551 OR2X1_LOC_508/A OR2X1_LOC_532/B 0.01fF
C11552 AND2X1_LOC_777/a_36_24# OR2X1_LOC_3/Y 0.01fF
C11553 OR2X1_LOC_306/Y AND2X1_LOC_856/B 0.16fF
C11554 OR2X1_LOC_437/a_8_216# OR2X1_LOC_59/Y 0.04fF
C11555 AND2X1_LOC_784/A AND2X1_LOC_578/A 0.05fF
C11556 OR2X1_LOC_815/a_36_216# AND2X1_LOC_793/Y 0.00fF
C11557 OR2X1_LOC_287/B OR2X1_LOC_401/Y 0.01fF
C11558 OR2X1_LOC_748/A AND2X1_LOC_347/a_36_24# 0.00fF
C11559 OR2X1_LOC_595/A AND2X1_LOC_657/A 0.09fF
C11560 OR2X1_LOC_70/Y OR2X1_LOC_418/Y 0.01fF
C11561 OR2X1_LOC_230/a_8_216# AND2X1_LOC_650/Y 0.01fF
C11562 OR2X1_LOC_306/Y AND2X1_LOC_863/A 0.09fF
C11563 AND2X1_LOC_366/A OR2X1_LOC_47/Y 0.00fF
C11564 AND2X1_LOC_727/A AND2X1_LOC_653/B 0.01fF
C11565 OR2X1_LOC_189/Y OR2X1_LOC_152/Y 0.03fF
C11566 OR2X1_LOC_532/B OR2X1_LOC_733/a_36_216# 0.00fF
C11567 AND2X1_LOC_95/Y AND2X1_LOC_309/a_36_24# 0.00fF
C11568 OR2X1_LOC_833/a_8_216# OR2X1_LOC_276/B 0.02fF
C11569 OR2X1_LOC_74/A AND2X1_LOC_240/Y 0.03fF
C11570 OR2X1_LOC_377/A OR2X1_LOC_404/A 0.12fF
C11571 OR2X1_LOC_435/a_8_216# OR2X1_LOC_112/B 0.15fF
C11572 AND2X1_LOC_711/Y OR2X1_LOC_757/a_36_216# 0.00fF
C11573 OR2X1_LOC_440/A OR2X1_LOC_737/A 0.02fF
C11574 INPUT_1 OR2X1_LOC_39/A 0.06fF
C11575 AND2X1_LOC_64/Y AND2X1_LOC_36/Y 2.36fF
C11576 OR2X1_LOC_264/Y OR2X1_LOC_227/Y 0.07fF
C11577 OR2X1_LOC_380/A OR2X1_LOC_22/Y 0.05fF
C11578 OR2X1_LOC_189/Y OR2X1_LOC_527/Y 0.07fF
C11579 OR2X1_LOC_417/Y AND2X1_LOC_446/a_8_24# 0.01fF
C11580 OR2X1_LOC_605/a_36_216# OR2X1_LOC_787/Y 0.01fF
C11581 OR2X1_LOC_595/Y AND2X1_LOC_219/Y 0.02fF
C11582 AND2X1_LOC_580/A AND2X1_LOC_664/a_36_24# 0.01fF
C11583 OR2X1_LOC_244/A OR2X1_LOC_375/A 0.14fF
C11584 OR2X1_LOC_22/A OR2X1_LOC_44/Y 0.06fF
C11585 OR2X1_LOC_653/Y AND2X1_LOC_109/a_8_24# 0.23fF
C11586 OR2X1_LOC_427/A AND2X1_LOC_812/a_8_24# 0.02fF
C11587 AND2X1_LOC_866/A AND2X1_LOC_847/Y 0.01fF
C11588 OR2X1_LOC_416/Y AND2X1_LOC_234/a_8_24# 0.23fF
C11589 OR2X1_LOC_19/B OR2X1_LOC_585/A 0.09fF
C11590 OR2X1_LOC_506/a_8_216# OR2X1_LOC_130/Y 0.40fF
C11591 AND2X1_LOC_18/Y OR2X1_LOC_80/A 0.06fF
C11592 OR2X1_LOC_750/a_8_216# OR2X1_LOC_269/B -0.06fF
C11593 AND2X1_LOC_42/B AND2X1_LOC_51/Y 0.03fF
C11594 D_INPUT_0 AND2X1_LOC_650/Y 0.02fF
C11595 AND2X1_LOC_599/a_8_24# AND2X1_LOC_36/Y 0.04fF
C11596 OR2X1_LOC_596/A OR2X1_LOC_704/a_8_216# 0.01fF
C11597 OR2X1_LOC_756/B OR2X1_LOC_351/a_8_216# 0.01fF
C11598 AND2X1_LOC_182/A OR2X1_LOC_437/A 0.02fF
C11599 OR2X1_LOC_631/B OR2X1_LOC_532/B 0.07fF
C11600 AND2X1_LOC_51/Y OR2X1_LOC_705/Y 0.01fF
C11601 AND2X1_LOC_512/Y OR2X1_LOC_761/a_8_216# 0.01fF
C11602 OR2X1_LOC_849/a_8_216# AND2X1_LOC_42/B 0.03fF
C11603 AND2X1_LOC_800/a_8_24# OR2X1_LOC_585/A 0.01fF
C11604 OR2X1_LOC_575/A OR2X1_LOC_493/Y 0.01fF
C11605 OR2X1_LOC_59/Y AND2X1_LOC_796/A 0.03fF
C11606 AND2X1_LOC_175/a_8_24# D_INPUT_0 0.01fF
C11607 OR2X1_LOC_220/A OR2X1_LOC_739/Y 0.02fF
C11608 AND2X1_LOC_209/Y AND2X1_LOC_213/a_8_24# 0.09fF
C11609 OR2X1_LOC_631/B AND2X1_LOC_665/a_8_24# 0.04fF
C11610 OR2X1_LOC_812/B AND2X1_LOC_225/a_8_24# 0.02fF
C11611 OR2X1_LOC_485/A AND2X1_LOC_687/Y 0.02fF
C11612 AND2X1_LOC_99/A OR2X1_LOC_813/Y 0.00fF
C11613 AND2X1_LOC_82/Y AND2X1_LOC_36/Y 0.00fF
C11614 AND2X1_LOC_808/A AND2X1_LOC_624/A 0.03fF
C11615 OR2X1_LOC_22/Y AND2X1_LOC_853/a_8_24# 0.04fF
C11616 OR2X1_LOC_22/Y AND2X1_LOC_650/a_36_24# 0.00fF
C11617 OR2X1_LOC_95/Y AND2X1_LOC_645/A 0.01fF
C11618 OR2X1_LOC_272/Y D_INPUT_0 0.03fF
C11619 OR2X1_LOC_161/B OR2X1_LOC_390/B 0.54fF
C11620 OR2X1_LOC_743/A OR2X1_LOC_31/Y 1.42fF
C11621 AND2X1_LOC_345/Y OR2X1_LOC_417/A 0.18fF
C11622 OR2X1_LOC_805/A AND2X1_LOC_237/a_36_24# 0.01fF
C11623 OR2X1_LOC_488/a_8_216# OR2X1_LOC_71/Y 0.01fF
C11624 AND2X1_LOC_455/a_8_24# AND2X1_LOC_455/B -0.01fF
C11625 AND2X1_LOC_721/Y AND2X1_LOC_284/a_8_24# 0.17fF
C11626 OR2X1_LOC_506/Y AND2X1_LOC_64/Y 0.05fF
C11627 AND2X1_LOC_135/a_8_24# OR2X1_LOC_532/B 0.01fF
C11628 OR2X1_LOC_814/A AND2X1_LOC_816/a_8_24# 0.01fF
C11629 OR2X1_LOC_85/A AND2X1_LOC_204/Y 0.02fF
C11630 OR2X1_LOC_778/Y D_INPUT_1 0.33fF
C11631 OR2X1_LOC_311/Y AND2X1_LOC_538/Y 0.02fF
C11632 AND2X1_LOC_539/Y OR2X1_LOC_12/Y 0.03fF
C11633 AND2X1_LOC_635/a_8_24# AND2X1_LOC_639/A 0.05fF
C11634 AND2X1_LOC_191/Y AND2X1_LOC_480/a_8_24# 0.03fF
C11635 AND2X1_LOC_727/A AND2X1_LOC_477/A 0.03fF
C11636 OR2X1_LOC_426/B OR2X1_LOC_320/a_8_216# 0.11fF
C11637 OR2X1_LOC_188/Y AND2X1_LOC_255/a_8_24# 0.24fF
C11638 OR2X1_LOC_323/A AND2X1_LOC_181/Y 0.03fF
C11639 AND2X1_LOC_504/a_8_24# OR2X1_LOC_560/A 0.03fF
C11640 OR2X1_LOC_696/A AND2X1_LOC_535/Y 0.03fF
C11641 OR2X1_LOC_859/A OR2X1_LOC_814/A 0.03fF
C11642 AND2X1_LOC_134/a_8_24# OR2X1_LOC_720/B 0.01fF
C11643 AND2X1_LOC_672/B INPUT_1 0.10fF
C11644 OR2X1_LOC_479/Y OR2X1_LOC_223/A 1.05fF
C11645 OR2X1_LOC_804/a_8_216# OR2X1_LOC_716/a_8_216# 0.47fF
C11646 OR2X1_LOC_375/A OR2X1_LOC_197/a_8_216# 0.02fF
C11647 OR2X1_LOC_647/A D_INPUT_1 0.03fF
C11648 OR2X1_LOC_403/a_8_216# OR2X1_LOC_532/B 0.01fF
C11649 OR2X1_LOC_78/Y OR2X1_LOC_771/B 0.03fF
C11650 OR2X1_LOC_45/B OR2X1_LOC_692/Y 0.01fF
C11651 OR2X1_LOC_246/A OR2X1_LOC_31/Y 0.01fF
C11652 AND2X1_LOC_774/a_8_24# AND2X1_LOC_774/A 0.04fF
C11653 AND2X1_LOC_486/Y OR2X1_LOC_13/B 0.01fF
C11654 OR2X1_LOC_64/Y AND2X1_LOC_648/B 0.01fF
C11655 AND2X1_LOC_18/Y OR2X1_LOC_115/B 0.02fF
C11656 AND2X1_LOC_364/a_36_24# OR2X1_LOC_12/Y 0.01fF
C11657 AND2X1_LOC_34/a_8_24# OR2X1_LOC_598/A 0.01fF
C11658 OR2X1_LOC_78/A OR2X1_LOC_502/a_8_216# 0.03fF
C11659 AND2X1_LOC_715/Y AND2X1_LOC_535/Y 0.13fF
C11660 AND2X1_LOC_555/Y AND2X1_LOC_363/Y 0.01fF
C11661 AND2X1_LOC_477/A OR2X1_LOC_95/Y 0.06fF
C11662 OR2X1_LOC_552/a_8_216# OR2X1_LOC_552/A 0.04fF
C11663 OR2X1_LOC_641/A OR2X1_LOC_227/B 0.08fF
C11664 OR2X1_LOC_528/Y GATE_579 0.04fF
C11665 OR2X1_LOC_12/Y AND2X1_LOC_771/B 0.26fF
C11666 OR2X1_LOC_160/A OR2X1_LOC_317/B 0.01fF
C11667 OR2X1_LOC_160/A OR2X1_LOC_501/a_8_216# 0.05fF
C11668 OR2X1_LOC_617/Y AND2X1_LOC_805/a_8_24# 0.01fF
C11669 AND2X1_LOC_53/Y AND2X1_LOC_56/a_36_24# 0.00fF
C11670 OR2X1_LOC_766/Y AND2X1_LOC_771/B 0.78fF
C11671 AND2X1_LOC_64/Y OR2X1_LOC_630/Y 0.16fF
C11672 OR2X1_LOC_131/A OR2X1_LOC_12/Y 1.45fF
C11673 OR2X1_LOC_146/a_8_216# OR2X1_LOC_744/A 0.18fF
C11674 OR2X1_LOC_45/B OR2X1_LOC_600/A 0.20fF
C11675 OR2X1_LOC_31/Y OR2X1_LOC_409/B 0.03fF
C11676 OR2X1_LOC_417/A AND2X1_LOC_649/Y 0.01fF
C11677 INPUT_1 OR2X1_LOC_826/Y 0.01fF
C11678 OR2X1_LOC_435/B OR2X1_LOC_390/B 0.01fF
C11679 VDD OR2X1_LOC_428/A 1.89fF
C11680 OR2X1_LOC_648/A OR2X1_LOC_392/B 0.01fF
C11681 OR2X1_LOC_89/A AND2X1_LOC_793/B 0.34fF
C11682 OR2X1_LOC_579/B OR2X1_LOC_579/a_36_216# 0.02fF
C11683 OR2X1_LOC_18/Y OR2X1_LOC_142/Y 0.03fF
C11684 D_INPUT_0 OR2X1_LOC_786/Y 0.01fF
C11685 OR2X1_LOC_362/A OR2X1_LOC_343/a_8_216# 0.01fF
C11686 AND2X1_LOC_554/a_8_24# OR2X1_LOC_744/A 0.01fF
C11687 AND2X1_LOC_19/Y AND2X1_LOC_7/B 0.02fF
C11688 AND2X1_LOC_776/Y OR2X1_LOC_164/Y 0.04fF
C11689 AND2X1_LOC_571/A OR2X1_LOC_103/Y 0.01fF
C11690 OR2X1_LOC_241/Y OR2X1_LOC_506/B 0.09fF
C11691 OR2X1_LOC_87/A OR2X1_LOC_707/a_8_216# 0.02fF
C11692 OR2X1_LOC_528/a_8_216# OR2X1_LOC_528/Y 0.15fF
C11693 VDD OR2X1_LOC_595/A 0.34fF
C11694 OR2X1_LOC_136/Y AND2X1_LOC_303/a_8_24# 0.23fF
C11695 OR2X1_LOC_160/B OR2X1_LOC_549/A 0.14fF
C11696 OR2X1_LOC_208/A AND2X1_LOC_57/a_8_24# 0.17fF
C11697 AND2X1_LOC_22/Y AND2X1_LOC_20/a_36_24# 0.01fF
C11698 OR2X1_LOC_217/Y OR2X1_LOC_217/A 0.00fF
C11699 OR2X1_LOC_600/A OR2X1_LOC_382/A 0.13fF
C11700 OR2X1_LOC_248/Y OR2X1_LOC_13/B 0.13fF
C11701 D_INPUT_0 OR2X1_LOC_644/A 0.17fF
C11702 OR2X1_LOC_546/B OR2X1_LOC_546/A 0.16fF
C11703 OR2X1_LOC_624/Y OR2X1_LOC_576/A 0.03fF
C11704 AND2X1_LOC_707/Y OR2X1_LOC_421/a_36_216# 0.01fF
C11705 OR2X1_LOC_583/a_8_216# OR2X1_LOC_583/Y -0.00fF
C11706 OR2X1_LOC_3/Y OR2X1_LOC_423/Y 0.01fF
C11707 AND2X1_LOC_316/a_8_24# AND2X1_LOC_7/B 0.03fF
C11708 OR2X1_LOC_40/Y OR2X1_LOC_505/Y 0.01fF
C11709 AND2X1_LOC_443/Y AND2X1_LOC_212/Y 0.02fF
C11710 AND2X1_LOC_370/a_8_24# AND2X1_LOC_716/Y 0.01fF
C11711 OR2X1_LOC_851/A AND2X1_LOC_273/a_36_24# 0.00fF
C11712 AND2X1_LOC_294/a_8_24# AND2X1_LOC_247/a_8_24# 0.23fF
C11713 D_INPUT_5 OR2X1_LOC_375/a_8_216# 0.01fF
C11714 OR2X1_LOC_620/Y OR2X1_LOC_703/a_8_216# 0.01fF
C11715 AND2X1_LOC_410/a_8_24# OR2X1_LOC_600/A 0.01fF
C11716 OR2X1_LOC_185/A OR2X1_LOC_718/a_8_216# 0.01fF
C11717 AND2X1_LOC_64/Y AND2X1_LOC_586/a_8_24# 0.02fF
C11718 AND2X1_LOC_647/a_8_24# OR2X1_LOC_16/A 0.01fF
C11719 OR2X1_LOC_13/Y OR2X1_LOC_59/Y 0.03fF
C11720 OR2X1_LOC_40/Y AND2X1_LOC_658/A 0.19fF
C11721 AND2X1_LOC_691/a_8_24# AND2X1_LOC_194/Y 0.01fF
C11722 AND2X1_LOC_3/Y OR2X1_LOC_712/B 0.09fF
C11723 AND2X1_LOC_215/Y VDD 0.19fF
C11724 OR2X1_LOC_6/B OR2X1_LOC_56/A 0.21fF
C11725 AND2X1_LOC_91/B OR2X1_LOC_506/A 0.09fF
C11726 OR2X1_LOC_643/a_8_216# OR2X1_LOC_539/B 0.02fF
C11727 OR2X1_LOC_778/Y OR2X1_LOC_180/B 0.05fF
C11728 OR2X1_LOC_437/a_8_216# OR2X1_LOC_437/Y 0.05fF
C11729 OR2X1_LOC_6/B OR2X1_LOC_819/a_8_216# 0.04fF
C11730 OR2X1_LOC_696/A AND2X1_LOC_576/Y 0.01fF
C11731 OR2X1_LOC_122/Y OR2X1_LOC_106/a_8_216# 0.40fF
C11732 AND2X1_LOC_756/a_8_24# OR2X1_LOC_604/A 0.11fF
C11733 OR2X1_LOC_494/Y OR2X1_LOC_51/Y 0.03fF
C11734 OR2X1_LOC_289/a_8_216# OR2X1_LOC_289/Y -0.00fF
C11735 OR2X1_LOC_347/Y OR2X1_LOC_244/Y 0.06fF
C11736 OR2X1_LOC_676/a_8_216# INPUT_0 0.01fF
C11737 AND2X1_LOC_95/Y OR2X1_LOC_721/a_8_216# 0.01fF
C11738 OR2X1_LOC_114/a_36_216# OR2X1_LOC_362/A 0.00fF
C11739 AND2X1_LOC_707/a_36_24# OR2X1_LOC_51/Y 0.00fF
C11740 AND2X1_LOC_76/Y AND2X1_LOC_786/Y 0.34fF
C11741 OR2X1_LOC_175/Y OR2X1_LOC_539/Y 0.10fF
C11742 OR2X1_LOC_190/A OR2X1_LOC_78/A 0.02fF
C11743 OR2X1_LOC_59/Y OR2X1_LOC_627/Y 0.00fF
C11744 OR2X1_LOC_113/Y OR2X1_LOC_160/B 0.00fF
C11745 OR2X1_LOC_45/B OR2X1_LOC_619/Y 0.13fF
C11746 OR2X1_LOC_406/Y AND2X1_LOC_807/Y 0.06fF
C11747 OR2X1_LOC_516/A AND2X1_LOC_794/a_8_24# 0.01fF
C11748 AND2X1_LOC_146/a_8_24# OR2X1_LOC_546/A 0.20fF
C11749 AND2X1_LOC_729/Y OR2X1_LOC_312/a_8_216# 0.04fF
C11750 OR2X1_LOC_158/A OR2X1_LOC_92/Y 0.24fF
C11751 OR2X1_LOC_650/a_8_216# AND2X1_LOC_92/Y 0.01fF
C11752 OR2X1_LOC_160/A AND2X1_LOC_44/Y 0.69fF
C11753 OR2X1_LOC_604/A AND2X1_LOC_160/a_8_24# 0.01fF
C11754 AND2X1_LOC_321/a_8_24# OR2X1_LOC_486/Y 0.02fF
C11755 OR2X1_LOC_137/a_8_216# OR2X1_LOC_66/A 0.01fF
C11756 AND2X1_LOC_721/Y OR2X1_LOC_406/a_8_216# 0.01fF
C11757 OR2X1_LOC_315/Y OR2X1_LOC_428/A 0.00fF
C11758 OR2X1_LOC_604/A AND2X1_LOC_562/B 0.08fF
C11759 AND2X1_LOC_714/B AND2X1_LOC_832/a_8_24# 0.04fF
C11760 AND2X1_LOC_12/Y OR2X1_LOC_706/a_8_216# 0.01fF
C11761 OR2X1_LOC_539/Y AND2X1_LOC_417/a_8_24# 0.04fF
C11762 AND2X1_LOC_86/Y OR2X1_LOC_549/A 0.02fF
C11763 AND2X1_LOC_110/Y OR2X1_LOC_623/B 0.03fF
C11764 OR2X1_LOC_319/a_8_216# OR2X1_LOC_151/A 0.03fF
C11765 OR2X1_LOC_45/B OR2X1_LOC_88/A 0.00fF
C11766 OR2X1_LOC_673/A OR2X1_LOC_68/B 0.14fF
C11767 OR2X1_LOC_769/B INPUT_0 0.03fF
C11768 OR2X1_LOC_158/A OR2X1_LOC_257/a_8_216# 0.02fF
C11769 AND2X1_LOC_12/Y OR2X1_LOC_390/A 0.03fF
C11770 OR2X1_LOC_589/A OR2X1_LOC_432/Y 0.02fF
C11771 AND2X1_LOC_335/a_8_24# OR2X1_LOC_56/A 0.03fF
C11772 AND2X1_LOC_47/Y OR2X1_LOC_446/B 0.12fF
C11773 AND2X1_LOC_388/a_8_24# AND2X1_LOC_810/B 0.02fF
C11774 OR2X1_LOC_113/a_36_216# OR2X1_LOC_643/A 0.00fF
C11775 INPUT_5 OR2X1_LOC_51/Y 0.05fF
C11776 OR2X1_LOC_44/Y AND2X1_LOC_769/Y 0.03fF
C11777 OR2X1_LOC_109/Y AND2X1_LOC_476/Y 0.19fF
C11778 AND2X1_LOC_738/B OR2X1_LOC_441/Y 0.07fF
C11779 AND2X1_LOC_663/B OR2X1_LOC_759/Y 0.01fF
C11780 OR2X1_LOC_441/Y OR2X1_LOC_56/A 0.06fF
C11781 AND2X1_LOC_498/a_8_24# OR2X1_LOC_499/B 0.09fF
C11782 AND2X1_LOC_70/Y OR2X1_LOC_833/a_8_216# 0.01fF
C11783 AND2X1_LOC_22/Y OR2X1_LOC_849/A 0.01fF
C11784 AND2X1_LOC_47/Y OR2X1_LOC_303/B 0.03fF
C11785 OR2X1_LOC_467/A OR2X1_LOC_469/Y 0.00fF
C11786 OR2X1_LOC_268/a_36_216# OR2X1_LOC_268/Y 0.00fF
C11787 AND2X1_LOC_374/Y AND2X1_LOC_786/Y 0.02fF
C11788 OR2X1_LOC_249/Y OR2X1_LOC_362/A 0.22fF
C11789 OR2X1_LOC_251/Y OR2X1_LOC_428/A 0.02fF
C11790 OR2X1_LOC_51/Y OR2X1_LOC_46/a_36_216# 0.00fF
C11791 OR2X1_LOC_139/A AND2X1_LOC_3/Y 0.10fF
C11792 AND2X1_LOC_462/B OR2X1_LOC_68/B 0.05fF
C11793 OR2X1_LOC_648/A AND2X1_LOC_58/a_36_24# 0.01fF
C11794 OR2X1_LOC_203/Y AND2X1_LOC_256/a_36_24# 0.00fF
C11795 OR2X1_LOC_52/B AND2X1_LOC_786/Y 0.02fF
C11796 OR2X1_LOC_312/Y AND2X1_LOC_457/a_8_24# 0.01fF
C11797 OR2X1_LOC_715/B OR2X1_LOC_510/Y 0.00fF
C11798 AND2X1_LOC_99/Y OR2X1_LOC_91/A 0.06fF
C11799 AND2X1_LOC_341/a_8_24# AND2X1_LOC_211/B 0.00fF
C11800 OR2X1_LOC_49/A AND2X1_LOC_102/a_8_24# 0.04fF
C11801 OR2X1_LOC_47/Y AND2X1_LOC_738/Y 0.04fF
C11802 OR2X1_LOC_795/B OR2X1_LOC_785/B 0.01fF
C11803 OR2X1_LOC_43/A OR2X1_LOC_381/a_8_216# 0.01fF
C11804 OR2X1_LOC_526/Y AND2X1_LOC_621/Y 0.08fF
C11805 OR2X1_LOC_440/A OR2X1_LOC_788/B 0.11fF
C11806 OR2X1_LOC_151/A OR2X1_LOC_203/Y 0.07fF
C11807 OR2X1_LOC_7/A AND2X1_LOC_219/A 0.09fF
C11808 OR2X1_LOC_251/Y OR2X1_LOC_595/A 0.01fF
C11809 AND2X1_LOC_76/Y AND2X1_LOC_218/Y 0.02fF
C11810 AND2X1_LOC_723/Y OR2X1_LOC_165/Y 0.02fF
C11811 OR2X1_LOC_525/Y OR2X1_LOC_744/A 0.19fF
C11812 AND2X1_LOC_56/B OR2X1_LOC_596/a_8_216# 0.01fF
C11813 OR2X1_LOC_158/A OR2X1_LOC_271/Y 0.11fF
C11814 OR2X1_LOC_335/a_8_216# OR2X1_LOC_121/B 0.01fF
C11815 OR2X1_LOC_6/B AND2X1_LOC_56/B 0.03fF
C11816 OR2X1_LOC_485/A OR2X1_LOC_373/Y 0.03fF
C11817 OR2X1_LOC_170/Y OR2X1_LOC_566/a_8_216# 0.01fF
C11818 OR2X1_LOC_743/A AND2X1_LOC_213/B 0.03fF
C11819 OR2X1_LOC_222/A AND2X1_LOC_18/Y 0.03fF
C11820 AND2X1_LOC_842/B AND2X1_LOC_242/B 0.33fF
C11821 AND2X1_LOC_366/a_8_24# AND2X1_LOC_848/Y 0.03fF
C11822 OR2X1_LOC_45/B OR2X1_LOC_372/a_8_216# 0.01fF
C11823 OR2X1_LOC_700/Y OR2X1_LOC_59/Y 0.01fF
C11824 OR2X1_LOC_161/A OR2X1_LOC_363/A 0.01fF
C11825 AND2X1_LOC_366/A OR2X1_LOC_625/Y 0.09fF
C11826 OR2X1_LOC_715/B OR2X1_LOC_810/A 0.01fF
C11827 OR2X1_LOC_6/B AND2X1_LOC_8/Y 0.12fF
C11828 OR2X1_LOC_709/A OR2X1_LOC_702/A 1.01fF
C11829 OR2X1_LOC_405/A AND2X1_LOC_372/a_8_24# 0.01fF
C11830 OR2X1_LOC_172/a_8_216# OR2X1_LOC_172/Y 0.00fF
C11831 OR2X1_LOC_457/a_8_216# OR2X1_LOC_787/B 0.07fF
C11832 OR2X1_LOC_402/Y OR2X1_LOC_78/Y 0.12fF
C11833 OR2X1_LOC_494/Y OR2X1_LOC_667/a_8_216# 0.01fF
C11834 OR2X1_LOC_40/Y OR2X1_LOC_626/a_36_216# 0.02fF
C11835 OR2X1_LOC_168/B AND2X1_LOC_601/a_8_24# 0.20fF
C11836 OR2X1_LOC_680/A AND2X1_LOC_548/Y 0.89fF
C11837 AND2X1_LOC_700/a_8_24# OR2X1_LOC_269/B 0.01fF
C11838 OR2X1_LOC_154/A OR2X1_LOC_768/A 0.01fF
C11839 OR2X1_LOC_178/Y OR2X1_LOC_36/Y 0.00fF
C11840 OR2X1_LOC_756/B OR2X1_LOC_456/a_36_216# 0.00fF
C11841 AND2X1_LOC_286/a_36_24# AND2X1_LOC_286/Y 0.00fF
C11842 OR2X1_LOC_169/a_36_216# AND2X1_LOC_92/Y 0.02fF
C11843 AND2X1_LOC_113/a_8_24# OR2X1_LOC_427/A 0.02fF
C11844 AND2X1_LOC_539/Y AND2X1_LOC_801/B 0.02fF
C11845 AND2X1_LOC_73/a_8_24# AND2X1_LOC_56/B 0.00fF
C11846 OR2X1_LOC_70/Y OR2X1_LOC_13/Y 0.02fF
C11847 VDD OR2X1_LOC_355/B -0.00fF
C11848 AND2X1_LOC_95/Y OR2X1_LOC_436/B 0.01fF
C11849 AND2X1_LOC_719/Y OR2X1_LOC_279/Y 0.10fF
C11850 OR2X1_LOC_417/A AND2X1_LOC_465/A 0.07fF
C11851 OR2X1_LOC_517/A OR2X1_LOC_39/A 0.03fF
C11852 OR2X1_LOC_599/A OR2X1_LOC_597/a_8_216# 0.01fF
C11853 OR2X1_LOC_744/A OR2X1_LOC_497/Y 0.07fF
C11854 VDD OR2X1_LOC_733/B -0.00fF
C11855 AND2X1_LOC_61/Y AND2X1_LOC_339/a_8_24# -0.00fF
C11856 OR2X1_LOC_834/A OR2X1_LOC_449/B 0.03fF
C11857 INPUT_5 OR2X1_LOC_375/A 0.02fF
C11858 AND2X1_LOC_658/A OR2X1_LOC_7/A 0.15fF
C11859 AND2X1_LOC_191/Y OR2X1_LOC_627/Y 0.08fF
C11860 AND2X1_LOC_181/a_8_24# OR2X1_LOC_26/Y 0.02fF
C11861 OR2X1_LOC_22/Y AND2X1_LOC_774/A 0.03fF
C11862 AND2X1_LOC_550/A AND2X1_LOC_804/Y 0.03fF
C11863 AND2X1_LOC_555/a_8_24# AND2X1_LOC_663/B 0.01fF
C11864 OR2X1_LOC_811/A OR2X1_LOC_269/a_8_216# 0.02fF
C11865 OR2X1_LOC_643/A OR2X1_LOC_658/a_36_216# 0.00fF
C11866 OR2X1_LOC_521/Y OR2X1_LOC_39/A 0.02fF
C11867 OR2X1_LOC_529/Y OR2X1_LOC_56/A 0.00fF
C11868 AND2X1_LOC_711/Y OR2X1_LOC_627/Y 0.03fF
C11869 OR2X1_LOC_406/Y OR2X1_LOC_95/Y 0.03fF
C11870 AND2X1_LOC_833/a_8_24# OR2X1_LOC_39/A 0.03fF
C11871 OR2X1_LOC_524/Y OR2X1_LOC_52/B 0.11fF
C11872 OR2X1_LOC_702/A AND2X1_LOC_70/Y 0.03fF
C11873 AND2X1_LOC_721/Y AND2X1_LOC_675/A 0.02fF
C11874 OR2X1_LOC_793/A AND2X1_LOC_39/a_8_24# 0.05fF
C11875 AND2X1_LOC_711/Y AND2X1_LOC_500/Y 0.08fF
C11876 OR2X1_LOC_784/a_36_216# OR2X1_LOC_78/A 0.00fF
C11877 OR2X1_LOC_351/B OR2X1_LOC_750/A 0.46fF
C11878 OR2X1_LOC_799/A OR2X1_LOC_506/A 0.03fF
C11879 VDD AND2X1_LOC_674/a_8_24# 0.00fF
C11880 OR2X1_LOC_18/Y OR2X1_LOC_118/Y 0.03fF
C11881 AND2X1_LOC_22/Y OR2X1_LOC_440/A 0.03fF
C11882 OR2X1_LOC_491/a_8_216# AND2X1_LOC_465/Y 0.47fF
C11883 OR2X1_LOC_329/B OR2X1_LOC_371/Y 0.09fF
C11884 AND2X1_LOC_703/Y OR2X1_LOC_95/Y 0.01fF
C11885 OR2X1_LOC_710/B AND2X1_LOC_51/Y 0.01fF
C11886 OR2X1_LOC_35/B OR2X1_LOC_35/Y 0.73fF
C11887 OR2X1_LOC_326/B AND2X1_LOC_56/B 0.00fF
C11888 AND2X1_LOC_91/B D_INPUT_1 0.51fF
C11889 AND2X1_LOC_47/Y AND2X1_LOC_248/a_36_24# 0.00fF
C11890 OR2X1_LOC_40/Y AND2X1_LOC_814/a_8_24# 0.01fF
C11891 AND2X1_LOC_120/a_8_24# OR2X1_LOC_59/Y 0.03fF
C11892 AND2X1_LOC_727/a_8_24# AND2X1_LOC_810/Y 0.02fF
C11893 OR2X1_LOC_256/A OR2X1_LOC_595/A 0.02fF
C11894 AND2X1_LOC_139/a_8_24# OR2X1_LOC_7/A 0.02fF
C11895 OR2X1_LOC_525/Y AND2X1_LOC_840/B 0.84fF
C11896 AND2X1_LOC_862/A OR2X1_LOC_39/A 0.01fF
C11897 OR2X1_LOC_3/Y AND2X1_LOC_367/A 0.05fF
C11898 AND2X1_LOC_624/A OR2X1_LOC_39/A 0.06fF
C11899 AND2X1_LOC_175/B OR2X1_LOC_265/Y 0.01fF
C11900 OR2X1_LOC_473/Y OR2X1_LOC_78/A 0.03fF
C11901 AND2X1_LOC_583/a_36_24# OR2X1_LOC_636/A 0.00fF
C11902 AND2X1_LOC_70/Y OR2X1_LOC_476/B 0.38fF
C11903 AND2X1_LOC_580/A AND2X1_LOC_573/A 0.03fF
C11904 OR2X1_LOC_778/Y OR2X1_LOC_737/A 0.54fF
C11905 INPUT_7 OR2X1_LOC_587/a_8_216# 0.05fF
C11906 OR2X1_LOC_474/a_8_216# OR2X1_LOC_244/Y 0.01fF
C11907 OR2X1_LOC_364/A OR2X1_LOC_161/A 0.07fF
C11908 AND2X1_LOC_124/a_36_24# OR2X1_LOC_67/A 0.00fF
C11909 OR2X1_LOC_452/a_36_216# AND2X1_LOC_425/Y 0.00fF
C11910 OR2X1_LOC_185/Y OR2X1_LOC_161/A 0.07fF
C11911 OR2X1_LOC_668/Y AND2X1_LOC_669/a_8_24# 0.23fF
C11912 AND2X1_LOC_95/Y OR2X1_LOC_643/A 0.03fF
C11913 AND2X1_LOC_91/B OR2X1_LOC_356/a_36_216# 0.01fF
C11914 OR2X1_LOC_814/A OR2X1_LOC_66/A 2.38fF
C11915 AND2X1_LOC_466/a_8_24# AND2X1_LOC_470/A 0.00fF
C11916 AND2X1_LOC_454/Y AND2X1_LOC_466/a_36_24# 0.01fF
C11917 OR2X1_LOC_502/A AND2X1_LOC_4/a_8_24# 0.01fF
C11918 AND2X1_LOC_95/Y OR2X1_LOC_778/Y 0.03fF
C11919 OR2X1_LOC_859/A OR2X1_LOC_244/Y 0.43fF
C11920 OR2X1_LOC_170/a_8_216# OR2X1_LOC_170/Y 0.00fF
C11921 AND2X1_LOC_95/Y OR2X1_LOC_472/A 0.03fF
C11922 OR2X1_LOC_22/Y AND2X1_LOC_434/a_8_24# 0.02fF
C11923 OR2X1_LOC_181/B OR2X1_LOC_564/A 0.12fF
C11924 OR2X1_LOC_663/A AND2X1_LOC_51/Y 0.00fF
C11925 OR2X1_LOC_639/B OR2X1_LOC_269/B 0.05fF
C11926 OR2X1_LOC_235/B OR2X1_LOC_293/a_8_216# 0.05fF
C11927 OR2X1_LOC_18/Y OR2X1_LOC_238/Y 0.03fF
C11928 OR2X1_LOC_342/B OR2X1_LOC_342/a_8_216# 0.01fF
C11929 OR2X1_LOC_18/Y OR2X1_LOC_24/Y 0.65fF
C11930 AND2X1_LOC_72/B OR2X1_LOC_342/A 0.01fF
C11931 OR2X1_LOC_542/B AND2X1_LOC_47/Y 0.03fF
C11932 OR2X1_LOC_64/Y AND2X1_LOC_863/a_8_24# 0.01fF
C11933 OR2X1_LOC_154/A AND2X1_LOC_393/a_36_24# 0.00fF
C11934 OR2X1_LOC_648/A OR2X1_LOC_532/B 0.08fF
C11935 OR2X1_LOC_161/B OR2X1_LOC_493/Y 0.10fF
C11936 OR2X1_LOC_64/Y OR2X1_LOC_265/a_8_216# 0.06fF
C11937 OR2X1_LOC_161/B OR2X1_LOC_801/B 0.07fF
C11938 AND2X1_LOC_859/Y OR2X1_LOC_26/Y 0.01fF
C11939 AND2X1_LOC_131/a_8_24# OR2X1_LOC_786/Y 0.01fF
C11940 OR2X1_LOC_31/Y OR2X1_LOC_12/a_8_216# 0.01fF
C11941 D_INPUT_0 OR2X1_LOC_234/Y 0.03fF
C11942 AND2X1_LOC_40/Y OR2X1_LOC_643/Y 0.03fF
C11943 OR2X1_LOC_562/A OR2X1_LOC_348/B 0.03fF
C11944 AND2X1_LOC_31/Y OR2X1_LOC_779/A 0.01fF
C11945 OR2X1_LOC_490/Y AND2X1_LOC_572/A 0.03fF
C11946 OR2X1_LOC_756/B OR2X1_LOC_288/A 0.01fF
C11947 OR2X1_LOC_682/a_8_216# OR2X1_LOC_682/Y 0.01fF
C11948 OR2X1_LOC_600/A AND2X1_LOC_838/B 0.02fF
C11949 OR2X1_LOC_837/Y AND2X1_LOC_826/a_8_24# 0.01fF
C11950 OR2X1_LOC_598/Y OR2X1_LOC_644/A 0.01fF
C11951 OR2X1_LOC_91/A AND2X1_LOC_476/A 0.07fF
C11952 OR2X1_LOC_298/a_8_216# OR2X1_LOC_31/Y 0.01fF
C11953 AND2X1_LOC_473/Y OR2X1_LOC_521/a_36_216# 0.12fF
C11954 D_INPUT_7 AND2X1_LOC_17/Y 0.01fF
C11955 OR2X1_LOC_333/B OR2X1_LOC_269/B 0.12fF
C11956 AND2X1_LOC_47/Y OR2X1_LOC_736/A 0.46fF
C11957 OR2X1_LOC_786/Y OR2X1_LOC_795/B 0.12fF
C11958 AND2X1_LOC_31/Y OR2X1_LOC_736/Y 0.00fF
C11959 OR2X1_LOC_87/A AND2X1_LOC_67/Y 0.00fF
C11960 OR2X1_LOC_748/A OR2X1_LOC_817/Y 0.01fF
C11961 AND2X1_LOC_12/Y OR2X1_LOC_750/A 0.03fF
C11962 AND2X1_LOC_374/a_8_24# OR2X1_LOC_31/Y 0.02fF
C11963 OR2X1_LOC_364/A AND2X1_LOC_51/Y 0.22fF
C11964 OR2X1_LOC_329/B AND2X1_LOC_116/a_8_24# 0.01fF
C11965 OR2X1_LOC_614/Y AND2X1_LOC_31/Y 0.01fF
C11966 AND2X1_LOC_95/Y OR2X1_LOC_113/A 0.01fF
C11967 OR2X1_LOC_185/Y AND2X1_LOC_51/Y 4.12fF
C11968 OR2X1_LOC_287/B OR2X1_LOC_843/a_36_216# 0.00fF
C11969 OR2X1_LOC_185/A OR2X1_LOC_243/B 0.15fF
C11970 INPUT_1 AND2X1_LOC_278/a_8_24# 0.17fF
C11971 OR2X1_LOC_404/Y AND2X1_LOC_669/a_36_24# 0.00fF
C11972 OR2X1_LOC_216/A OR2X1_LOC_506/B 0.02fF
C11973 OR2X1_LOC_49/A OR2X1_LOC_71/A 0.19fF
C11974 OR2X1_LOC_95/Y OR2X1_LOC_586/a_36_216# 0.00fF
C11975 OR2X1_LOC_377/A INPUT_1 0.27fF
C11976 OR2X1_LOC_51/Y AND2X1_LOC_228/a_8_24# 0.08fF
C11977 OR2X1_LOC_405/a_8_216# OR2X1_LOC_532/B 0.01fF
C11978 OR2X1_LOC_426/A AND2X1_LOC_452/a_8_24# 0.01fF
C11979 OR2X1_LOC_3/Y OR2X1_LOC_490/Y 0.01fF
C11980 OR2X1_LOC_3/Y OR2X1_LOC_74/A 0.10fF
C11981 OR2X1_LOC_757/A AND2X1_LOC_793/Y 0.55fF
C11982 AND2X1_LOC_92/Y OR2X1_LOC_339/Y 0.03fF
C11983 AND2X1_LOC_64/Y OR2X1_LOC_469/B 0.12fF
C11984 OR2X1_LOC_17/Y OR2X1_LOC_47/a_8_216# 0.00fF
C11985 AND2X1_LOC_211/B AND2X1_LOC_853/a_8_24# 0.01fF
C11986 OR2X1_LOC_528/Y AND2X1_LOC_657/A 0.12fF
C11987 INPUT_1 AND2X1_LOC_824/B 0.01fF
C11988 AND2X1_LOC_59/Y AND2X1_LOC_7/Y 0.11fF
C11989 OR2X1_LOC_97/A OR2X1_LOC_777/B 0.03fF
C11990 AND2X1_LOC_99/A AND2X1_LOC_866/A 0.03fF
C11991 AND2X1_LOC_40/Y OR2X1_LOC_786/Y 0.02fF
C11992 OR2X1_LOC_74/A AND2X1_LOC_631/Y 0.08fF
C11993 OR2X1_LOC_17/Y AND2X1_LOC_651/B 0.09fF
C11994 OR2X1_LOC_427/A AND2X1_LOC_796/Y 0.03fF
C11995 OR2X1_LOC_853/a_8_216# OR2X1_LOC_771/B 0.05fF
C11996 AND2X1_LOC_91/B OR2X1_LOC_180/B 0.03fF
C11997 OR2X1_LOC_131/Y AND2X1_LOC_141/B 0.28fF
C11998 OR2X1_LOC_576/A OR2X1_LOC_141/a_36_216# 0.00fF
C11999 D_INPUT_5 OR2X1_LOC_2/a_8_216# 0.01fF
C12000 AND2X1_LOC_733/Y AND2X1_LOC_795/Y 0.00fF
C12001 INPUT_1 OR2X1_LOC_85/A 1.41fF
C12002 AND2X1_LOC_72/B OR2X1_LOC_735/a_36_216# 0.00fF
C12003 AND2X1_LOC_810/Y AND2X1_LOC_621/Y 0.03fF
C12004 OR2X1_LOC_168/Y OR2X1_LOC_170/a_8_216# 0.02fF
C12005 D_INPUT_0 OR2X1_LOC_204/Y 0.02fF
C12006 OR2X1_LOC_532/Y AND2X1_LOC_44/Y 0.07fF
C12007 OR2X1_LOC_3/Y OR2X1_LOC_261/A 0.00fF
C12008 OR2X1_LOC_813/A OR2X1_LOC_6/A 0.00fF
C12009 OR2X1_LOC_287/B OR2X1_LOC_846/A 0.00fF
C12010 OR2X1_LOC_329/B AND2X1_LOC_222/Y 0.03fF
C12011 OR2X1_LOC_485/A AND2X1_LOC_849/A 0.01fF
C12012 AND2X1_LOC_449/a_36_24# OR2X1_LOC_428/A 0.00fF
C12013 AND2X1_LOC_772/B AND2X1_LOC_657/A 0.02fF
C12014 AND2X1_LOC_40/Y OR2X1_LOC_644/A 0.14fF
C12015 AND2X1_LOC_315/a_8_24# OR2X1_LOC_223/A 0.01fF
C12016 OR2X1_LOC_175/Y OR2X1_LOC_319/Y 0.03fF
C12017 AND2X1_LOC_56/B AND2X1_LOC_47/Y 0.12fF
C12018 OR2X1_LOC_659/B AND2X1_LOC_47/Y 0.04fF
C12019 AND2X1_LOC_512/Y OR2X1_LOC_331/a_36_216# 0.01fF
C12020 OR2X1_LOC_428/A AND2X1_LOC_269/a_8_24# 0.10fF
C12021 OR2X1_LOC_516/Y OR2X1_LOC_816/A 0.07fF
C12022 AND2X1_LOC_8/Y AND2X1_LOC_47/Y 0.07fF
C12023 VDD OR2X1_LOC_366/Y 0.65fF
C12024 AND2X1_LOC_307/a_8_24# AND2X1_LOC_307/Y 0.01fF
C12025 OR2X1_LOC_323/A AND2X1_LOC_564/B 0.11fF
C12026 OR2X1_LOC_36/Y AND2X1_LOC_318/Y 0.01fF
C12027 OR2X1_LOC_461/Y OR2X1_LOC_472/B 0.01fF
C12028 OR2X1_LOC_243/a_8_216# AND2X1_LOC_42/B 0.01fF
C12029 OR2X1_LOC_808/B AND2X1_LOC_31/Y 0.02fF
C12030 OR2X1_LOC_487/a_8_216# OR2X1_LOC_417/A 0.01fF
C12031 OR2X1_LOC_680/Y OR2X1_LOC_679/A 0.01fF
C12032 AND2X1_LOC_21/Y AND2X1_LOC_47/Y 0.07fF
C12033 D_INPUT_3 OR2X1_LOC_83/A 0.02fF
C12034 OR2X1_LOC_631/a_8_216# OR2X1_LOC_598/A 0.03fF
C12035 OR2X1_LOC_696/A OR2X1_LOC_16/A 4.44fF
C12036 AND2X1_LOC_34/a_8_24# AND2X1_LOC_462/Y 0.11fF
C12037 OR2X1_LOC_190/A D_GATE_366 0.04fF
C12038 OR2X1_LOC_696/A AND2X1_LOC_714/a_36_24# 0.01fF
C12039 OR2X1_LOC_502/A OR2X1_LOC_68/B 0.43fF
C12040 OR2X1_LOC_31/Y OR2X1_LOC_229/Y 0.01fF
C12041 AND2X1_LOC_351/Y OR2X1_LOC_46/A 0.01fF
C12042 OR2X1_LOC_278/A AND2X1_LOC_633/Y 0.02fF
C12043 OR2X1_LOC_146/a_8_216# AND2X1_LOC_213/B 0.01fF
C12044 AND2X1_LOC_202/Y AND2X1_LOC_206/a_8_24# 0.11fF
C12045 AND2X1_LOC_345/Y OR2X1_LOC_55/a_8_216# 0.03fF
C12046 AND2X1_LOC_22/Y OR2X1_LOC_721/a_8_216# 0.06fF
C12047 OR2X1_LOC_364/A OR2X1_LOC_551/B 0.10fF
C12048 AND2X1_LOC_715/Y OR2X1_LOC_16/A 0.05fF
C12049 OR2X1_LOC_214/B OR2X1_LOC_155/A 0.07fF
C12050 OR2X1_LOC_541/A OR2X1_LOC_777/B 0.03fF
C12051 AND2X1_LOC_56/B OR2X1_LOC_598/A 0.08fF
C12052 AND2X1_LOC_724/a_8_24# AND2X1_LOC_724/A 0.03fF
C12053 OR2X1_LOC_696/A OR2X1_LOC_108/Y 0.07fF
C12054 AND2X1_LOC_476/A OR2X1_LOC_27/Y 0.04fF
C12055 OR2X1_LOC_161/A OR2X1_LOC_568/A 0.07fF
C12056 AND2X1_LOC_230/a_8_24# OR2X1_LOC_68/B 0.01fF
C12057 AND2X1_LOC_8/Y OR2X1_LOC_598/A 0.10fF
C12058 AND2X1_LOC_785/a_8_24# AND2X1_LOC_778/Y 0.01fF
C12059 AND2X1_LOC_465/Y OR2X1_LOC_95/Y 0.10fF
C12060 AND2X1_LOC_723/a_8_24# OR2X1_LOC_437/A 0.20fF
C12061 AND2X1_LOC_40/Y OR2X1_LOC_181/Y 0.00fF
C12062 OR2X1_LOC_756/B AND2X1_LOC_36/Y 0.26fF
C12063 OR2X1_LOC_89/A AND2X1_LOC_846/a_8_24# 0.01fF
C12064 OR2X1_LOC_506/A OR2X1_LOC_446/B 0.03fF
C12065 OR2X1_LOC_598/Y AND2X1_LOC_829/a_8_24# 0.08fF
C12066 OR2X1_LOC_278/Y OR2X1_LOC_437/A 0.03fF
C12067 OR2X1_LOC_323/A AND2X1_LOC_325/a_36_24# 0.00fF
C12068 OR2X1_LOC_468/Y OR2X1_LOC_353/a_8_216# 0.03fF
C12069 AND2X1_LOC_755/a_8_24# OR2X1_LOC_366/Y 0.03fF
C12070 OR2X1_LOC_52/B OR2X1_LOC_746/Y 0.01fF
C12071 OR2X1_LOC_3/Y AND2X1_LOC_647/Y 0.00fF
C12072 OR2X1_LOC_708/B AND2X1_LOC_31/Y 0.03fF
C12073 OR2X1_LOC_45/B OR2X1_LOC_527/a_8_216# 0.01fF
C12074 OR2X1_LOC_256/a_36_216# OR2X1_LOC_13/B 0.00fF
C12075 OR2X1_LOC_506/A OR2X1_LOC_728/a_8_216# 0.03fF
C12076 OR2X1_LOC_774/Y OR2X1_LOC_557/a_8_216# 0.01fF
C12077 AND2X1_LOC_810/A AND2X1_LOC_388/Y 0.01fF
C12078 AND2X1_LOC_2/a_8_24# INPUT_6 0.02fF
C12079 OR2X1_LOC_53/Y OR2X1_LOC_51/Y 0.03fF
C12080 OR2X1_LOC_756/B OR2X1_LOC_333/a_8_216# 0.02fF
C12081 OR2X1_LOC_51/Y AND2X1_LOC_241/a_36_24# 0.00fF
C12082 OR2X1_LOC_354/A OR2X1_LOC_354/a_8_216# 0.01fF
C12083 OR2X1_LOC_185/A OR2X1_LOC_771/B 0.07fF
C12084 AND2X1_LOC_321/a_36_24# OR2X1_LOC_469/B 0.01fF
C12085 AND2X1_LOC_64/Y AND2X1_LOC_167/a_8_24# 0.04fF
C12086 OR2X1_LOC_756/B OR2X1_LOC_334/A 0.01fF
C12087 OR2X1_LOC_541/A OR2X1_LOC_831/B 0.50fF
C12088 OR2X1_LOC_185/A OR2X1_LOC_209/A 0.15fF
C12089 VDD OR2X1_LOC_389/a_8_216# 0.00fF
C12090 OR2X1_LOC_490/Y AND2X1_LOC_772/a_8_24# 0.02fF
C12091 OR2X1_LOC_535/A OR2X1_LOC_356/a_8_216# 0.47fF
C12092 OR2X1_LOC_436/Y OR2X1_LOC_468/a_36_216# 0.03fF
C12093 AND2X1_LOC_766/a_8_24# OR2X1_LOC_78/Y 0.01fF
C12094 AND2X1_LOC_596/a_8_24# OR2X1_LOC_829/A 0.20fF
C12095 OR2X1_LOC_30/a_36_216# D_INPUT_6 0.03fF
C12096 OR2X1_LOC_805/A OR2X1_LOC_723/B 0.09fF
C12097 OR2X1_LOC_276/A OR2X1_LOC_276/B 0.01fF
C12098 OR2X1_LOC_348/a_8_216# OR2X1_LOC_348/Y -0.00fF
C12099 AND2X1_LOC_372/a_36_24# OR2X1_LOC_831/B 0.01fF
C12100 AND2X1_LOC_141/B AND2X1_LOC_657/A 0.18fF
C12101 AND2X1_LOC_706/Y AND2X1_LOC_447/Y 0.02fF
C12102 OR2X1_LOC_135/a_8_216# OR2X1_LOC_56/A 0.08fF
C12103 OR2X1_LOC_185/A OR2X1_LOC_776/A 0.02fF
C12104 AND2X1_LOC_773/Y AND2X1_LOC_219/Y 0.24fF
C12105 OR2X1_LOC_589/A AND2X1_LOC_537/a_8_24# 0.01fF
C12106 OR2X1_LOC_158/A OR2X1_LOC_600/A 3.65fF
C12107 OR2X1_LOC_158/A AND2X1_LOC_335/Y 0.01fF
C12108 AND2X1_LOC_51/Y OR2X1_LOC_568/A 0.44fF
C12109 AND2X1_LOC_153/a_8_24# AND2X1_LOC_238/a_8_24# 0.23fF
C12110 OR2X1_LOC_744/A AND2X1_LOC_249/a_8_24# 0.01fF
C12111 AND2X1_LOC_592/Y VDD 0.08fF
C12112 OR2X1_LOC_778/Y OR2X1_LOC_788/B 0.03fF
C12113 OR2X1_LOC_516/Y AND2X1_LOC_807/Y 0.10fF
C12114 OR2X1_LOC_91/A OR2X1_LOC_766/a_8_216# 0.10fF
C12115 OR2X1_LOC_369/Y AND2X1_LOC_212/A 0.79fF
C12116 OR2X1_LOC_528/Y VDD 0.90fF
C12117 AND2X1_LOC_40/Y AND2X1_LOC_829/a_8_24# 0.01fF
C12118 OR2X1_LOC_375/A AND2X1_LOC_581/a_8_24# 0.20fF
C12119 OR2X1_LOC_53/Y OR2X1_LOC_16/Y 0.00fF
C12120 AND2X1_LOC_70/Y AND2X1_LOC_262/a_8_24# 0.01fF
C12121 OR2X1_LOC_756/B AND2X1_LOC_488/a_8_24# 0.01fF
C12122 AND2X1_LOC_91/B OR2X1_LOC_737/A 0.10fF
C12123 AND2X1_LOC_22/Y OR2X1_LOC_637/A 0.01fF
C12124 OR2X1_LOC_158/A AND2X1_LOC_296/a_8_24# 0.02fF
C12125 OR2X1_LOC_672/a_8_216# OR2X1_LOC_56/A 0.02fF
C12126 AND2X1_LOC_22/Y OR2X1_LOC_436/B 0.01fF
C12127 VDD OR2X1_LOC_583/Y 0.12fF
C12128 OR2X1_LOC_325/A AND2X1_LOC_44/Y 0.94fF
C12129 AND2X1_LOC_190/a_8_24# OR2X1_LOC_40/Y 0.08fF
C12130 AND2X1_LOC_93/a_8_24# OR2X1_LOC_78/A 0.07fF
C12131 OR2X1_LOC_678/Y OR2X1_LOC_713/A 0.73fF
C12132 AND2X1_LOC_23/a_8_24# OR2X1_LOC_228/Y 0.04fF
C12133 OR2X1_LOC_76/Y AND2X1_LOC_36/Y 0.03fF
C12134 OR2X1_LOC_151/A OR2X1_LOC_78/B 5.67fF
C12135 AND2X1_LOC_739/B AND2X1_LOC_739/a_8_24# 0.01fF
C12136 AND2X1_LOC_658/B AND2X1_LOC_549/Y 0.03fF
C12137 AND2X1_LOC_48/A OR2X1_LOC_68/B 0.03fF
C12138 AND2X1_LOC_91/B AND2X1_LOC_95/Y 0.21fF
C12139 OR2X1_LOC_6/B AND2X1_LOC_92/Y 0.01fF
C12140 OR2X1_LOC_339/a_8_216# VDD 0.21fF
C12141 AND2X1_LOC_794/B AND2X1_LOC_512/Y 0.00fF
C12142 OR2X1_LOC_591/Y AND2X1_LOC_605/Y 0.17fF
C12143 AND2X1_LOC_772/B VDD 0.04fF
C12144 OR2X1_LOC_244/Y OR2X1_LOC_66/A 0.85fF
C12145 AND2X1_LOC_658/B AND2X1_LOC_500/Y 0.03fF
C12146 AND2X1_LOC_169/a_8_24# OR2X1_LOC_331/Y 0.01fF
C12147 AND2X1_LOC_69/a_36_24# OR2X1_LOC_68/B 0.00fF
C12148 AND2X1_LOC_40/Y OR2X1_LOC_535/A 0.00fF
C12149 AND2X1_LOC_535/Y AND2X1_LOC_436/a_8_24# 0.00fF
C12150 OR2X1_LOC_526/Y OR2X1_LOC_59/Y 0.01fF
C12151 OR2X1_LOC_18/Y AND2X1_LOC_208/Y 0.01fF
C12152 AND2X1_LOC_59/Y OR2X1_LOC_703/a_36_216# 0.00fF
C12153 AND2X1_LOC_570/Y AND2X1_LOC_501/a_8_24# 0.01fF
C12154 OR2X1_LOC_188/a_36_216# OR2X1_LOC_375/A 0.00fF
C12155 AND2X1_LOC_655/A OR2X1_LOC_321/a_8_216# 0.12fF
C12156 AND2X1_LOC_307/Y OR2X1_LOC_13/B 0.03fF
C12157 OR2X1_LOC_468/a_8_216# OR2X1_LOC_854/A 0.01fF
C12158 OR2X1_LOC_151/A OR2X1_LOC_721/Y 0.17fF
C12159 OR2X1_LOC_44/Y AND2X1_LOC_783/B 0.04fF
C12160 AND2X1_LOC_536/a_36_24# AND2X1_LOC_7/B 0.01fF
C12161 OR2X1_LOC_19/B OR2X1_LOC_437/A 0.00fF
C12162 OR2X1_LOC_218/Y AND2X1_LOC_31/Y 0.06fF
C12163 OR2X1_LOC_744/A OR2X1_LOC_380/a_8_216# 0.05fF
C12164 AND2X1_LOC_426/a_8_24# OR2X1_LOC_161/B 0.01fF
C12165 AND2X1_LOC_676/a_8_24# AND2X1_LOC_213/B 0.01fF
C12166 AND2X1_LOC_474/a_8_24# AND2X1_LOC_244/A 0.10fF
C12167 OR2X1_LOC_600/A AND2X1_LOC_98/Y 0.22fF
C12168 OR2X1_LOC_851/A OR2X1_LOC_831/A 0.02fF
C12169 OR2X1_LOC_160/B OR2X1_LOC_499/B 0.09fF
C12170 OR2X1_LOC_744/A OR2X1_LOC_743/a_8_216# 0.02fF
C12171 AND2X1_LOC_40/a_8_24# AND2X1_LOC_11/Y 0.01fF
C12172 AND2X1_LOC_340/Y OR2X1_LOC_118/Y 0.01fF
C12173 VDD AND2X1_LOC_512/Y 0.85fF
C12174 AND2X1_LOC_190/a_36_24# OR2X1_LOC_744/A 0.01fF
C12175 AND2X1_LOC_64/Y OR2X1_LOC_592/a_8_216# 0.05fF
C12176 OR2X1_LOC_287/B OR2X1_LOC_363/a_36_216# 0.00fF
C12177 OR2X1_LOC_269/a_8_216# OR2X1_LOC_344/A 0.01fF
C12178 AND2X1_LOC_624/A AND2X1_LOC_727/B 0.03fF
C12179 OR2X1_LOC_417/A OR2X1_LOC_384/Y 0.41fF
C12180 OR2X1_LOC_298/Y OR2X1_LOC_12/Y 0.10fF
C12181 OR2X1_LOC_600/A OR2X1_LOC_103/Y 0.03fF
C12182 AND2X1_LOC_56/B OR2X1_LOC_34/A 0.03fF
C12183 INPUT_0 OR2X1_LOC_91/A 0.13fF
C12184 OR2X1_LOC_600/A OR2X1_LOC_594/Y 0.07fF
C12185 OR2X1_LOC_158/A OR2X1_LOC_619/Y 0.21fF
C12186 AND2X1_LOC_22/Y OR2X1_LOC_643/A 0.07fF
C12187 INPUT_0 OR2X1_LOC_637/Y 0.03fF
C12188 OR2X1_LOC_121/a_8_216# OR2X1_LOC_185/Y 0.03fF
C12189 OR2X1_LOC_158/A AND2X1_LOC_356/a_8_24# 0.06fF
C12190 AND2X1_LOC_675/Y AND2X1_LOC_549/a_36_24# 0.07fF
C12191 AND2X1_LOC_367/A OR2X1_LOC_329/B 0.23fF
C12192 OR2X1_LOC_52/B AND2X1_LOC_202/Y 0.03fF
C12193 AND2X1_LOC_22/Y OR2X1_LOC_778/Y 0.05fF
C12194 OR2X1_LOC_516/A AND2X1_LOC_794/B 0.01fF
C12195 AND2X1_LOC_535/Y AND2X1_LOC_354/Y 0.03fF
C12196 OR2X1_LOC_532/B OR2X1_LOC_112/A 0.00fF
C12197 OR2X1_LOC_6/a_8_216# OR2X1_LOC_428/A 0.02fF
C12198 OR2X1_LOC_49/A OR2X1_LOC_820/B 0.03fF
C12199 OR2X1_LOC_151/A OR2X1_LOC_375/A 0.03fF
C12200 OR2X1_LOC_709/a_8_216# OR2X1_LOC_154/A 0.04fF
C12201 OR2X1_LOC_78/A AND2X1_LOC_615/a_8_24# 0.01fF
C12202 OR2X1_LOC_45/B AND2X1_LOC_454/A 0.02fF
C12203 AND2X1_LOC_792/Y AND2X1_LOC_793/B 0.02fF
C12204 OR2X1_LOC_469/Y OR2X1_LOC_78/A 0.03fF
C12205 OR2X1_LOC_708/B OR2X1_LOC_708/a_36_216# 0.01fF
C12206 AND2X1_LOC_474/A OR2X1_LOC_517/A 0.03fF
C12207 OR2X1_LOC_528/Y OR2X1_LOC_616/Y 0.97fF
C12208 OR2X1_LOC_45/B OR2X1_LOC_371/a_36_216# 0.00fF
C12209 AND2X1_LOC_340/Y OR2X1_LOC_262/Y 0.46fF
C12210 OR2X1_LOC_385/Y AND2X1_LOC_407/a_8_24# 0.02fF
C12211 AND2X1_LOC_715/A AND2X1_LOC_662/B 0.02fF
C12212 OR2X1_LOC_598/Y OR2X1_LOC_828/B 0.00fF
C12213 OR2X1_LOC_676/a_8_216# OR2X1_LOC_407/a_8_216# 0.47fF
C12214 OR2X1_LOC_313/a_8_216# OR2X1_LOC_604/A 0.01fF
C12215 OR2X1_LOC_666/A OR2X1_LOC_427/A 0.07fF
C12216 VDD OR2X1_LOC_624/A 2.15fF
C12217 OR2X1_LOC_499/a_8_216# AND2X1_LOC_18/Y 0.05fF
C12218 OR2X1_LOC_421/A AND2X1_LOC_655/A 0.01fF
C12219 AND2X1_LOC_787/a_8_24# AND2X1_LOC_469/B 0.01fF
C12220 AND2X1_LOC_861/B AND2X1_LOC_865/a_8_24# 0.01fF
C12221 OR2X1_LOC_820/B OR2X1_LOC_381/a_36_216# 0.00fF
C12222 AND2X1_LOC_798/a_8_24# AND2X1_LOC_727/A 0.01fF
C12223 AND2X1_LOC_737/Y OR2X1_LOC_524/Y 0.05fF
C12224 AND2X1_LOC_663/A AND2X1_LOC_804/Y 0.05fF
C12225 OR2X1_LOC_842/A OR2X1_LOC_161/A 0.02fF
C12226 OR2X1_LOC_696/A AND2X1_LOC_128/a_8_24# 0.01fF
C12227 AND2X1_LOC_805/Y OR2X1_LOC_59/Y 0.00fF
C12228 OR2X1_LOC_280/Y AND2X1_LOC_786/Y 0.07fF
C12229 AND2X1_LOC_42/B OR2X1_LOC_576/A 0.07fF
C12230 OR2X1_LOC_551/B OR2X1_LOC_578/B 0.68fF
C12231 AND2X1_LOC_41/a_36_24# OR2X1_LOC_375/A 0.00fF
C12232 AND2X1_LOC_784/A AND2X1_LOC_182/A 0.04fF
C12233 OR2X1_LOC_604/A AND2X1_LOC_470/A 0.01fF
C12234 AND2X1_LOC_250/a_36_24# OR2X1_LOC_580/A 0.00fF
C12235 OR2X1_LOC_834/a_8_216# OR2X1_LOC_502/A 0.08fF
C12236 OR2X1_LOC_156/A OR2X1_LOC_87/A 0.13fF
C12237 VDD AND2X1_LOC_342/Y 0.02fF
C12238 AND2X1_LOC_2/Y AND2X1_LOC_157/a_8_24# 0.01fF
C12239 AND2X1_LOC_220/a_8_24# AND2X1_LOC_220/Y 0.00fF
C12240 AND2X1_LOC_669/a_8_24# OR2X1_LOC_66/A 0.01fF
C12241 OR2X1_LOC_620/a_8_216# OR2X1_LOC_620/B 0.05fF
C12242 OR2X1_LOC_216/A OR2X1_LOC_473/a_8_216# 0.04fF
C12243 AND2X1_LOC_786/a_36_24# OR2X1_LOC_70/Y 0.00fF
C12244 OR2X1_LOC_106/Y AND2X1_LOC_115/a_8_24# 0.09fF
C12245 OR2X1_LOC_512/Y OR2X1_LOC_779/B 0.08fF
C12246 AND2X1_LOC_57/Y OR2X1_LOC_532/B 0.00fF
C12247 OR2X1_LOC_696/A OR2X1_LOC_225/a_36_216# -0.00fF
C12248 AND2X1_LOC_468/B AND2X1_LOC_471/Y 0.23fF
C12249 OR2X1_LOC_130/A OR2X1_LOC_35/Y 0.02fF
C12250 AND2X1_LOC_27/a_8_24# AND2X1_LOC_7/B 0.08fF
C12251 OR2X1_LOC_516/Y OR2X1_LOC_95/Y 0.03fF
C12252 OR2X1_LOC_154/A OR2X1_LOC_702/a_8_216# 0.01fF
C12253 AND2X1_LOC_303/B OR2X1_LOC_426/B -0.00fF
C12254 AND2X1_LOC_46/a_8_24# AND2X1_LOC_44/Y 0.01fF
C12255 AND2X1_LOC_555/Y INPUT_1 0.00fF
C12256 OR2X1_LOC_400/B VDD 0.00fF
C12257 AND2X1_LOC_719/Y AND2X1_LOC_717/B 0.03fF
C12258 OR2X1_LOC_494/Y AND2X1_LOC_359/B 0.01fF
C12259 AND2X1_LOC_557/Y AND2X1_LOC_561/B 0.15fF
C12260 OR2X1_LOC_681/a_8_216# OR2X1_LOC_52/B 0.03fF
C12261 D_INPUT_4 OR2X1_LOC_2/Y 0.09fF
C12262 OR2X1_LOC_92/Y OR2X1_LOC_586/Y 0.08fF
C12263 OR2X1_LOC_518/Y OR2X1_LOC_417/A -0.05fF
C12264 AND2X1_LOC_363/Y AND2X1_LOC_359/B 0.02fF
C12265 AND2X1_LOC_861/B AND2X1_LOC_621/Y 0.07fF
C12266 OR2X1_LOC_45/B AND2X1_LOC_334/a_8_24# 0.03fF
C12267 AND2X1_LOC_768/a_8_24# AND2X1_LOC_361/A 0.03fF
C12268 AND2X1_LOC_570/Y OR2X1_LOC_44/Y 0.20fF
C12269 AND2X1_LOC_367/A AND2X1_LOC_113/Y 0.05fF
C12270 OR2X1_LOC_74/A AND2X1_LOC_477/Y 0.07fF
C12271 OR2X1_LOC_803/a_8_216# OR2X1_LOC_448/Y 0.10fF
C12272 OR2X1_LOC_864/A OR2X1_LOC_641/Y 0.00fF
C12273 VDD OR2X1_LOC_552/a_8_216# 0.00fF
C12274 OR2X1_LOC_329/B AND2X1_LOC_114/a_36_24# 0.00fF
C12275 VDD AND2X1_LOC_105/a_8_24# -0.00fF
C12276 OR2X1_LOC_7/A AND2X1_LOC_614/a_8_24# 0.01fF
C12277 AND2X1_LOC_40/Y OR2X1_LOC_220/B 0.03fF
C12278 OR2X1_LOC_837/A OR2X1_LOC_837/a_8_216# 0.02fF
C12279 OR2X1_LOC_682/Y VDD 0.05fF
C12280 OR2X1_LOC_683/Y OR2X1_LOC_12/Y 0.02fF
C12281 OR2X1_LOC_40/Y OR2X1_LOC_278/a_8_216# 0.01fF
C12282 AND2X1_LOC_67/a_8_24# OR2X1_LOC_375/A 0.01fF
C12283 AND2X1_LOC_127/a_8_24# AND2X1_LOC_44/Y 0.01fF
C12284 AND2X1_LOC_522/a_8_24# AND2X1_LOC_107/a_8_24# 0.23fF
C12285 AND2X1_LOC_22/Y OR2X1_LOC_113/A 0.03fF
C12286 AND2X1_LOC_340/a_8_24# OR2X1_LOC_3/Y 0.01fF
C12287 VDD OR2X1_LOC_555/A 0.21fF
C12288 OR2X1_LOC_3/Y AND2X1_LOC_860/A 0.00fF
C12289 AND2X1_LOC_686/a_8_24# OR2X1_LOC_16/A 0.01fF
C12290 OR2X1_LOC_185/A OR2X1_LOC_808/a_8_216# 0.01fF
C12291 OR2X1_LOC_22/Y AND2X1_LOC_786/Y 0.12fF
C12292 OR2X1_LOC_114/Y OR2X1_LOC_235/B 0.16fF
C12293 OR2X1_LOC_604/A OR2X1_LOC_258/Y 0.02fF
C12294 OR2X1_LOC_528/Y AND2X1_LOC_624/a_8_24# 0.01fF
C12295 AND2X1_LOC_207/a_8_24# OR2X1_LOC_43/A 0.01fF
C12296 OR2X1_LOC_485/A AND2X1_LOC_447/Y 0.12fF
C12297 AND2X1_LOC_40/Y OR2X1_LOC_828/B 0.04fF
C12298 AND2X1_LOC_306/a_8_24# OR2X1_LOC_449/B 0.05fF
C12299 OR2X1_LOC_651/B OR2X1_LOC_375/A 0.04fF
C12300 OR2X1_LOC_517/A OR2X1_LOC_85/A 0.29fF
C12301 AND2X1_LOC_355/a_8_24# AND2X1_LOC_434/Y 0.01fF
C12302 OR2X1_LOC_599/A OR2X1_LOC_697/Y 0.01fF
C12303 OR2X1_LOC_698/Y OR2X1_LOC_36/Y 0.01fF
C12304 AND2X1_LOC_678/a_8_24# OR2X1_LOC_12/Y 0.07fF
C12305 VDD AND2X1_LOC_483/a_8_24# 0.00fF
C12306 OR2X1_LOC_807/B OR2X1_LOC_362/B 0.01fF
C12307 OR2X1_LOC_792/Y OR2X1_LOC_807/A 0.04fF
C12308 VDD AND2X1_LOC_141/B 0.01fF
C12309 AND2X1_LOC_56/B OR2X1_LOC_828/a_8_216# 0.01fF
C12310 AND2X1_LOC_849/a_8_24# AND2X1_LOC_244/A 0.01fF
C12311 OR2X1_LOC_118/a_8_216# OR2X1_LOC_71/Y 0.01fF
C12312 AND2X1_LOC_95/Y OR2X1_LOC_799/A 0.00fF
C12313 D_INPUT_5 OR2X1_LOC_36/Y 0.03fF
C12314 AND2X1_LOC_17/Y AND2X1_LOC_50/a_8_24# 0.20fF
C12315 OR2X1_LOC_135/Y D_INPUT_0 0.13fF
C12316 AND2X1_LOC_70/Y OR2X1_LOC_863/B 0.01fF
C12317 AND2X1_LOC_392/A AND2X1_LOC_327/a_8_24# 0.05fF
C12318 OR2X1_LOC_158/A OR2X1_LOC_22/A 0.03fF
C12319 OR2X1_LOC_493/a_8_216# AND2X1_LOC_67/Y 0.15fF
C12320 OR2X1_LOC_634/A AND2X1_LOC_412/a_36_24# 0.00fF
C12321 OR2X1_LOC_329/B OR2X1_LOC_74/A 0.07fF
C12322 OR2X1_LOC_664/Y OR2X1_LOC_833/B 0.08fF
C12323 OR2X1_LOC_481/A OR2X1_LOC_56/A 0.20fF
C12324 AND2X1_LOC_228/Y AND2X1_LOC_174/a_8_24# 0.00fF
C12325 OR2X1_LOC_313/a_36_216# AND2X1_LOC_452/Y 0.01fF
C12326 VDD AND2X1_LOC_712/B 0.05fF
C12327 OR2X1_LOC_620/Y AND2X1_LOC_298/a_8_24# 0.00fF
C12328 OR2X1_LOC_503/A AND2X1_LOC_573/A 0.02fF
C12329 AND2X1_LOC_72/B OR2X1_LOC_140/B 0.01fF
C12330 GATE_366 OR2X1_LOC_427/A 0.01fF
C12331 OR2X1_LOC_3/Y OR2X1_LOC_459/A 0.04fF
C12332 AND2X1_LOC_41/A AND2X1_LOC_42/B 0.74fF
C12333 OR2X1_LOC_603/a_8_216# AND2X1_LOC_452/Y 0.03fF
C12334 AND2X1_LOC_134/a_8_24# AND2X1_LOC_18/Y 0.02fF
C12335 VDD OR2X1_LOC_54/Y 0.48fF
C12336 OR2X1_LOC_620/Y OR2X1_LOC_269/B 0.07fF
C12337 AND2X1_LOC_56/B OR2X1_LOC_506/A 0.07fF
C12338 OR2X1_LOC_642/a_8_216# OR2X1_LOC_185/A 0.01fF
C12339 AND2X1_LOC_391/Y OR2X1_LOC_64/Y 0.00fF
C12340 AND2X1_LOC_858/B OR2X1_LOC_64/Y 0.04fF
C12341 AND2X1_LOC_12/Y AND2X1_LOC_382/a_8_24# 0.01fF
C12342 OR2X1_LOC_687/Y AND2X1_LOC_43/B 0.03fF
C12343 AND2X1_LOC_41/A OR2X1_LOC_705/Y 0.08fF
C12344 OR2X1_LOC_669/a_36_216# OR2X1_LOC_278/Y 0.00fF
C12345 OR2X1_LOC_91/A OR2X1_LOC_64/Y 1.71fF
C12346 AND2X1_LOC_362/B AND2X1_LOC_227/Y 0.01fF
C12347 OR2X1_LOC_539/A OR2X1_LOC_702/A 0.78fF
C12348 OR2X1_LOC_312/Y OR2X1_LOC_427/A 0.00fF
C12349 OR2X1_LOC_6/A OR2X1_LOC_69/A 0.01fF
C12350 OR2X1_LOC_36/Y AND2X1_LOC_648/a_8_24# 0.08fF
C12351 OR2X1_LOC_655/B AND2X1_LOC_18/Y 0.01fF
C12352 OR2X1_LOC_74/Y OR2X1_LOC_74/A 0.02fF
C12353 OR2X1_LOC_753/A OR2X1_LOC_38/a_8_216# 0.03fF
C12354 VDD OR2X1_LOC_447/Y 0.08fF
C12355 OR2X1_LOC_51/Y INPUT_1 0.15fF
C12356 AND2X1_LOC_191/Y AND2X1_LOC_805/Y 0.03fF
C12357 AND2X1_LOC_479/Y AND2X1_LOC_480/A 0.00fF
C12358 AND2X1_LOC_52/a_8_24# AND2X1_LOC_51/Y 0.14fF
C12359 OR2X1_LOC_6/B D_INPUT_3 0.92fF
C12360 OR2X1_LOC_743/A AND2X1_LOC_809/A 0.00fF
C12361 AND2X1_LOC_112/a_36_24# OR2X1_LOC_417/A 0.01fF
C12362 OR2X1_LOC_278/Y AND2X1_LOC_243/a_8_24# 0.01fF
C12363 OR2X1_LOC_47/Y OR2X1_LOC_13/Y 0.02fF
C12364 OR2X1_LOC_109/Y OR2X1_LOC_485/A 0.24fF
C12365 AND2X1_LOC_711/Y AND2X1_LOC_805/Y 5.87fF
C12366 OR2X1_LOC_154/A OR2X1_LOC_269/B 0.29fF
C12367 OR2X1_LOC_71/Y OR2X1_LOC_56/A 0.02fF
C12368 OR2X1_LOC_170/A OR2X1_LOC_468/Y 0.01fF
C12369 OR2X1_LOC_476/B OR2X1_LOC_634/a_36_216# 0.01fF
C12370 D_INPUT_0 OR2X1_LOC_78/A 0.16fF
C12371 OR2X1_LOC_168/B OR2X1_LOC_168/A 0.04fF
C12372 OR2X1_LOC_303/B OR2X1_LOC_180/B 0.03fF
C12373 OR2X1_LOC_402/a_8_216# OR2X1_LOC_402/Y 0.01fF
C12374 AND2X1_LOC_40/Y OR2X1_LOC_436/a_36_216# 0.00fF
C12375 OR2X1_LOC_369/Y OR2X1_LOC_95/Y 0.00fF
C12376 AND2X1_LOC_190/a_36_24# OR2X1_LOC_31/Y 0.00fF
C12377 AND2X1_LOC_47/Y AND2X1_LOC_92/Y 0.26fF
C12378 VDD OR2X1_LOC_276/a_8_216# 0.21fF
C12379 AND2X1_LOC_391/Y OR2X1_LOC_417/A 1.09fF
C12380 AND2X1_LOC_307/a_8_24# OR2X1_LOC_427/A 0.08fF
C12381 AND2X1_LOC_858/B OR2X1_LOC_417/A 4.53fF
C12382 OR2X1_LOC_40/Y AND2X1_LOC_810/a_8_24# 0.02fF
C12383 AND2X1_LOC_70/Y OR2X1_LOC_276/A 0.01fF
C12384 OR2X1_LOC_91/Y OR2X1_LOC_529/Y 0.03fF
C12385 OR2X1_LOC_91/A OR2X1_LOC_417/A 0.77fF
C12386 INPUT_1 OR2X1_LOC_58/a_8_216# 0.02fF
C12387 AND2X1_LOC_654/a_36_24# OR2X1_LOC_6/A 0.00fF
C12388 AND2X1_LOC_702/Y OR2X1_LOC_299/a_8_216# 0.01fF
C12389 AND2X1_LOC_810/Y OR2X1_LOC_59/Y 0.07fF
C12390 OR2X1_LOC_670/Y OR2X1_LOC_672/Y 0.08fF
C12391 OR2X1_LOC_528/Y AND2X1_LOC_624/B 0.05fF
C12392 OR2X1_LOC_542/B OR2X1_LOC_284/B 0.61fF
C12393 AND2X1_LOC_658/A OR2X1_LOC_615/Y 0.19fF
C12394 OR2X1_LOC_251/Y AND2X1_LOC_105/a_8_24# 0.01fF
C12395 OR2X1_LOC_816/A AND2X1_LOC_793/B 0.01fF
C12396 AND2X1_LOC_259/Y OR2X1_LOC_820/B 0.00fF
C12397 OR2X1_LOC_186/Y OR2X1_LOC_170/Y 0.01fF
C12398 OR2X1_LOC_205/Y AND2X1_LOC_18/Y 0.18fF
C12399 OR2X1_LOC_565/A OR2X1_LOC_192/B 0.03fF
C12400 OR2X1_LOC_64/Y AND2X1_LOC_573/A 0.11fF
C12401 OR2X1_LOC_323/A OR2X1_LOC_437/A 0.05fF
C12402 OR2X1_LOC_66/Y OR2X1_LOC_631/A 0.01fF
C12403 OR2X1_LOC_631/B AND2X1_LOC_42/B 0.15fF
C12404 VDD OR2X1_LOC_84/Y 0.12fF
C12405 AND2X1_LOC_797/a_8_24# AND2X1_LOC_797/B 0.01fF
C12406 OR2X1_LOC_56/A D_INPUT_1 0.04fF
C12407 OR2X1_LOC_131/Y OR2X1_LOC_26/Y 0.03fF
C12408 OR2X1_LOC_154/A OR2X1_LOC_215/A 0.04fF
C12409 OR2X1_LOC_856/a_8_216# OR2X1_LOC_269/B 0.01fF
C12410 AND2X1_LOC_180/a_8_24# AND2X1_LOC_222/Y 0.01fF
C12411 AND2X1_LOC_324/a_8_24# OR2X1_LOC_36/Y 0.05fF
C12412 OR2X1_LOC_311/Y AND2X1_LOC_436/B 0.01fF
C12413 AND2X1_LOC_59/Y OR2X1_LOC_750/A 5.93fF
C12414 INPUT_1 AND2X1_LOC_642/a_8_24# 0.01fF
C12415 OR2X1_LOC_599/A OR2X1_LOC_696/Y 0.01fF
C12416 AND2X1_LOC_91/B OR2X1_LOC_788/B 0.04fF
C12417 AND2X1_LOC_31/Y OR2X1_LOC_596/A 0.03fF
C12418 AND2X1_LOC_845/Y OR2X1_LOC_278/Y 0.01fF
C12419 AND2X1_LOC_12/Y OR2X1_LOC_859/A 0.08fF
C12420 OR2X1_LOC_524/Y AND2X1_LOC_808/A 0.03fF
C12421 OR2X1_LOC_795/a_36_216# AND2X1_LOC_92/Y 0.01fF
C12422 OR2X1_LOC_596/A OR2X1_LOC_715/a_8_216# 0.01fF
C12423 OR2X1_LOC_190/Y OR2X1_LOC_192/B 0.35fF
C12424 OR2X1_LOC_131/Y OR2X1_LOC_89/A 0.01fF
C12425 OR2X1_LOC_43/A OR2X1_LOC_275/a_8_216# 0.06fF
C12426 OR2X1_LOC_690/A OR2X1_LOC_27/Y 0.03fF
C12427 OR2X1_LOC_175/Y OR2X1_LOC_777/B 0.07fF
C12428 OR2X1_LOC_725/A OR2X1_LOC_725/a_8_216# 0.39fF
C12429 AND2X1_LOC_175/B D_INPUT_0 0.01fF
C12430 OR2X1_LOC_46/A AND2X1_LOC_233/a_36_24# 0.00fF
C12431 OR2X1_LOC_193/A OR2X1_LOC_155/A 0.08fF
C12432 OR2X1_LOC_841/A OR2X1_LOC_318/B 0.00fF
C12433 OR2X1_LOC_40/Y OR2X1_LOC_72/Y 0.01fF
C12434 OR2X1_LOC_109/a_8_216# OR2X1_LOC_31/Y 0.09fF
C12435 AND2X1_LOC_556/a_36_24# OR2X1_LOC_615/Y 0.01fF
C12436 AND2X1_LOC_578/A OR2X1_LOC_280/Y 0.07fF
C12437 AND2X1_LOC_136/a_36_24# OR2X1_LOC_155/A 0.01fF
C12438 INPUT_1 OR2X1_LOC_375/A 0.58fF
C12439 AND2X1_LOC_514/Y AND2X1_LOC_661/A 0.02fF
C12440 AND2X1_LOC_564/B OR2X1_LOC_142/Y 0.07fF
C12441 AND2X1_LOC_116/Y AND2X1_LOC_473/a_8_24# 0.20fF
C12442 OR2X1_LOC_417/A AND2X1_LOC_573/A 0.08fF
C12443 OR2X1_LOC_657/a_36_216# OR2X1_LOC_62/B 0.00fF
C12444 OR2X1_LOC_19/B OR2X1_LOC_753/A 0.20fF
C12445 AND2X1_LOC_631/a_8_24# OR2X1_LOC_615/Y 0.02fF
C12446 OR2X1_LOC_654/A AND2X1_LOC_51/Y 0.06fF
C12447 OR2X1_LOC_485/A AND2X1_LOC_729/B 0.08fF
C12448 VDD OR2X1_LOC_513/a_8_216# 0.00fF
C12449 OR2X1_LOC_352/a_8_216# OR2X1_LOC_212/B 0.01fF
C12450 OR2X1_LOC_40/Y OR2X1_LOC_152/a_36_216# 0.02fF
C12451 AND2X1_LOC_342/Y OR2X1_LOC_256/A 0.33fF
C12452 AND2X1_LOC_61/Y AND2X1_LOC_203/a_8_24# 0.01fF
C12453 OR2X1_LOC_840/A OR2X1_LOC_804/A 0.10fF
C12454 AND2X1_LOC_53/Y OR2X1_LOC_87/A 0.02fF
C12455 OR2X1_LOC_777/B OR2X1_LOC_713/A 0.03fF
C12456 OR2X1_LOC_405/A OR2X1_LOC_473/A 0.01fF
C12457 AND2X1_LOC_61/Y AND2X1_LOC_206/Y 0.00fF
C12458 D_INPUT_0 OR2X1_LOC_155/A 0.19fF
C12459 AND2X1_LOC_47/Y OR2X1_LOC_551/a_8_216# 0.01fF
C12460 AND2X1_LOC_9/a_8_24# D_INPUT_1 0.07fF
C12461 AND2X1_LOC_43/B AND2X1_LOC_827/a_36_24# 0.01fF
C12462 OR2X1_LOC_669/Y OR2X1_LOC_417/A 0.18fF
C12463 OR2X1_LOC_633/a_36_216# OR2X1_LOC_68/B 0.00fF
C12464 OR2X1_LOC_223/A OR2X1_LOC_87/A 0.03fF
C12465 OR2X1_LOC_201/A OR2X1_LOC_68/B 0.29fF
C12466 OR2X1_LOC_566/A OR2X1_LOC_175/Y 0.27fF
C12467 AND2X1_LOC_56/B AND2X1_LOC_420/a_8_24# 0.03fF
C12468 OR2X1_LOC_696/A OR2X1_LOC_373/Y 0.00fF
C12469 AND2X1_LOC_753/B OR2X1_LOC_228/Y 0.01fF
C12470 AND2X1_LOC_91/B AND2X1_LOC_22/Y 0.25fF
C12471 AND2X1_LOC_56/B D_INPUT_1 0.03fF
C12472 AND2X1_LOC_529/a_8_24# OR2X1_LOC_71/A 0.01fF
C12473 AND2X1_LOC_390/B AND2X1_LOC_170/B 0.00fF
C12474 OR2X1_LOC_280/a_36_216# AND2X1_LOC_851/B 0.01fF
C12475 OR2X1_LOC_139/A AND2X1_LOC_7/B 0.07fF
C12476 AND2X1_LOC_681/a_8_24# AND2X1_LOC_3/Y 0.02fF
C12477 AND2X1_LOC_141/B OR2X1_LOC_256/A 0.12fF
C12478 AND2X1_LOC_8/Y D_INPUT_1 13.54fF
C12479 AND2X1_LOC_627/a_8_24# OR2X1_LOC_563/A 0.01fF
C12480 OR2X1_LOC_405/A OR2X1_LOC_228/Y 0.10fF
C12481 OR2X1_LOC_70/Y AND2X1_LOC_810/Y 0.07fF
C12482 OR2X1_LOC_520/B OR2X1_LOC_520/A 0.05fF
C12483 OR2X1_LOC_561/Y OR2X1_LOC_580/A 0.35fF
C12484 AND2X1_LOC_723/Y OR2X1_LOC_437/A 0.28fF
C12485 OR2X1_LOC_87/A OR2X1_LOC_705/B 0.15fF
C12486 AND2X1_LOC_710/Y AND2X1_LOC_789/Y 0.01fF
C12487 OR2X1_LOC_19/B AND2X1_LOC_845/Y 0.16fF
C12488 OR2X1_LOC_358/B OR2X1_LOC_358/A 0.00fF
C12489 OR2X1_LOC_97/A OR2X1_LOC_161/B 0.01fF
C12490 OR2X1_LOC_756/B OR2X1_LOC_571/Y 0.01fF
C12491 OR2X1_LOC_70/Y OR2X1_LOC_760/Y 0.04fF
C12492 AND2X1_LOC_512/a_8_24# OR2X1_LOC_599/Y 0.09fF
C12493 AND2X1_LOC_45/a_36_24# AND2X1_LOC_53/Y 0.01fF
C12494 AND2X1_LOC_229/a_8_24# OR2X1_LOC_231/B 0.01fF
C12495 OR2X1_LOC_291/A D_INPUT_1 0.04fF
C12496 OR2X1_LOC_756/B OR2X1_LOC_374/a_8_216# 0.01fF
C12497 OR2X1_LOC_174/A OR2X1_LOC_539/B 0.23fF
C12498 OR2X1_LOC_212/A OR2X1_LOC_357/A 0.14fF
C12499 AND2X1_LOC_64/Y AND2X1_LOC_313/a_8_24# 0.01fF
C12500 OR2X1_LOC_724/a_8_216# OR2X1_LOC_317/B 0.01fF
C12501 AND2X1_LOC_53/Y OR2X1_LOC_706/B 0.04fF
C12502 OR2X1_LOC_654/a_36_216# AND2X1_LOC_7/B 0.00fF
C12503 AND2X1_LOC_95/Y OR2X1_LOC_446/B 0.06fF
C12504 VDD OR2X1_LOC_556/a_8_216# 0.00fF
C12505 OR2X1_LOC_323/A AND2X1_LOC_715/A 0.32fF
C12506 OR2X1_LOC_427/A OR2X1_LOC_13/B 0.93fF
C12507 AND2X1_LOC_72/Y OR2X1_LOC_269/A 0.15fF
C12508 AND2X1_LOC_95/Y OR2X1_LOC_303/B 0.03fF
C12509 AND2X1_LOC_801/a_8_24# OR2X1_LOC_13/B 0.04fF
C12510 OR2X1_LOC_294/Y AND2X1_LOC_295/a_8_24# 0.07fF
C12511 AND2X1_LOC_95/Y OR2X1_LOC_728/a_8_216# 0.01fF
C12512 OR2X1_LOC_26/Y AND2X1_LOC_657/A 0.02fF
C12513 OR2X1_LOC_269/B OR2X1_LOC_198/A 0.01fF
C12514 AND2X1_LOC_67/Y OR2X1_LOC_493/Y 0.10fF
C12515 OR2X1_LOC_535/A OR2X1_LOC_356/A 0.08fF
C12516 OR2X1_LOC_630/Y OR2X1_LOC_140/B 0.07fF
C12517 AND2X1_LOC_721/Y OR2X1_LOC_600/A 0.05fF
C12518 AND2X1_LOC_170/B AND2X1_LOC_863/Y 0.00fF
C12519 AND2X1_LOC_803/B AND2X1_LOC_564/A 0.03fF
C12520 AND2X1_LOC_339/B OR2X1_LOC_589/A 0.02fF
C12521 AND2X1_LOC_741/Y AND2X1_LOC_480/A 0.10fF
C12522 OR2X1_LOC_156/Y OR2X1_LOC_803/A 0.01fF
C12523 OR2X1_LOC_151/A OR2X1_LOC_549/A 0.12fF
C12524 OR2X1_LOC_85/A OR2X1_LOC_150/a_8_216# 0.05fF
C12525 OR2X1_LOC_3/Y AND2X1_LOC_562/Y 0.01fF
C12526 AND2X1_LOC_3/Y OR2X1_LOC_68/B 0.11fF
C12527 AND2X1_LOC_592/Y AND2X1_LOC_713/a_8_24# 0.01fF
C12528 OR2X1_LOC_89/A AND2X1_LOC_657/A 0.09fF
C12529 AND2X1_LOC_390/B OR2X1_LOC_331/Y 0.02fF
C12530 D_INPUT_3 AND2X1_LOC_47/Y 0.81fF
C12531 OR2X1_LOC_647/B OR2X1_LOC_68/B 0.39fF
C12532 AND2X1_LOC_229/a_36_24# OR2X1_LOC_160/B 0.01fF
C12533 OR2X1_LOC_45/B AND2X1_LOC_570/Y 0.03fF
C12534 OR2X1_LOC_185/A OR2X1_LOC_593/B 0.04fF
C12535 OR2X1_LOC_80/a_8_216# OR2X1_LOC_47/Y 0.01fF
C12536 OR2X1_LOC_549/a_36_216# OR2X1_LOC_756/B 0.00fF
C12537 OR2X1_LOC_118/a_8_216# OR2X1_LOC_426/B 0.27fF
C12538 AND2X1_LOC_787/A AND2X1_LOC_469/B 0.00fF
C12539 OR2X1_LOC_160/B AND2X1_LOC_65/A 3.31fF
C12540 OR2X1_LOC_447/Y OR2X1_LOC_783/a_36_216# 0.02fF
C12541 OR2X1_LOC_121/Y OR2X1_LOC_66/A 0.01fF
C12542 AND2X1_LOC_43/B OR2X1_LOC_199/B 0.03fF
C12543 OR2X1_LOC_379/a_8_216# AND2X1_LOC_36/Y 0.01fF
C12544 AND2X1_LOC_70/Y OR2X1_LOC_294/Y 0.01fF
C12545 AND2X1_LOC_773/Y AND2X1_LOC_364/Y 0.39fF
C12546 OR2X1_LOC_12/Y AND2X1_LOC_434/Y 0.03fF
C12547 AND2X1_LOC_810/A OR2X1_LOC_329/B 0.03fF
C12548 OR2X1_LOC_12/Y AND2X1_LOC_219/Y 0.07fF
C12549 AND2X1_LOC_787/A AND2X1_LOC_733/Y 0.03fF
C12550 VDD OR2X1_LOC_565/A 0.16fF
C12551 INPUT_0 OR2X1_LOC_138/A 0.04fF
C12552 OR2X1_LOC_97/A OR2X1_LOC_435/B 0.00fF
C12553 VDD OR2X1_LOC_765/Y -0.00fF
C12554 OR2X1_LOC_510/A OR2X1_LOC_160/B 0.30fF
C12555 OR2X1_LOC_382/Y OR2X1_LOC_428/A 0.02fF
C12556 AND2X1_LOC_553/a_8_24# VDD 0.00fF
C12557 AND2X1_LOC_758/a_8_24# OR2X1_LOC_759/A 0.01fF
C12558 OR2X1_LOC_40/Y AND2X1_LOC_758/a_36_24# 0.01fF
C12559 OR2X1_LOC_114/B OR2X1_LOC_66/A 0.03fF
C12560 AND2X1_LOC_70/Y OR2X1_LOC_641/A 0.03fF
C12561 OR2X1_LOC_108/a_8_216# OR2X1_LOC_56/A 0.01fF
C12562 AND2X1_LOC_727/A OR2X1_LOC_533/A 0.01fF
C12563 OR2X1_LOC_117/a_36_216# OR2X1_LOC_92/Y 0.00fF
C12564 AND2X1_LOC_70/Y OR2X1_LOC_733/A 0.12fF
C12565 OR2X1_LOC_97/A OR2X1_LOC_61/Y 0.04fF
C12566 VDD OR2X1_LOC_190/Y 0.07fF
C12567 OR2X1_LOC_784/Y OR2X1_LOC_779/A 0.01fF
C12568 OR2X1_LOC_62/B OR2X1_LOC_80/A 0.05fF
C12569 AND2X1_LOC_505/a_8_24# OR2X1_LOC_78/A 0.02fF
C12570 D_INPUT_3 OR2X1_LOC_598/A 0.02fF
C12571 AND2X1_LOC_47/Y OR2X1_LOC_736/a_8_216# 0.01fF
C12572 OR2X1_LOC_653/Y OR2X1_LOC_61/A 0.02fF
C12573 OR2X1_LOC_600/A OR2X1_LOC_816/Y 0.00fF
C12574 OR2X1_LOC_757/Y AND2X1_LOC_791/a_8_24# 0.04fF
C12575 AND2X1_LOC_22/Y OR2X1_LOC_799/A 0.17fF
C12576 OR2X1_LOC_426/B OR2X1_LOC_56/A 0.48fF
C12577 OR2X1_LOC_354/A OR2X1_LOC_151/A 0.23fF
C12578 AND2X1_LOC_18/a_8_24# AND2X1_LOC_36/Y 0.01fF
C12579 OR2X1_LOC_604/A OR2X1_LOC_697/a_8_216# 0.14fF
C12580 AND2X1_LOC_347/Y AND2X1_LOC_347/B 0.11fF
C12581 OR2X1_LOC_31/Y OR2X1_LOC_588/a_36_216# 0.00fF
C12582 AND2X1_LOC_476/A AND2X1_LOC_222/Y 0.04fF
C12583 AND2X1_LOC_568/B AND2X1_LOC_364/Y 0.09fF
C12584 OR2X1_LOC_770/Y OR2X1_LOC_771/a_8_216# 0.39fF
C12585 OR2X1_LOC_139/A OR2X1_LOC_805/A 0.10fF
C12586 OR2X1_LOC_538/A OR2X1_LOC_66/A 0.05fF
C12587 OR2X1_LOC_45/B OR2X1_LOC_45/a_36_216# 0.00fF
C12588 AND2X1_LOC_350/B AND2X1_LOC_175/B 0.00fF
C12589 OR2X1_LOC_497/a_8_216# AND2X1_LOC_242/B 0.01fF
C12590 OR2X1_LOC_604/A OR2X1_LOC_698/Y 0.01fF
C12591 AND2X1_LOC_229/a_8_24# AND2X1_LOC_12/Y 0.09fF
C12592 OR2X1_LOC_117/a_36_216# OR2X1_LOC_65/B 0.03fF
C12593 OR2X1_LOC_128/B OR2X1_LOC_342/A 0.37fF
C12594 OR2X1_LOC_95/Y OR2X1_LOC_533/A 0.07fF
C12595 OR2X1_LOC_31/Y AND2X1_LOC_215/a_8_24# 0.01fF
C12596 OR2X1_LOC_710/B AND2X1_LOC_41/A 0.03fF
C12597 AND2X1_LOC_846/a_8_24# AND2X1_LOC_792/Y 0.02fF
C12598 OR2X1_LOC_532/B OR2X1_LOC_71/A 0.02fF
C12599 AND2X1_LOC_476/A OR2X1_LOC_68/B 0.01fF
C12600 AND2X1_LOC_658/B OR2X1_LOC_441/a_8_216# 0.05fF
C12601 OR2X1_LOC_39/A AND2X1_LOC_786/Y 0.17fF
C12602 OR2X1_LOC_476/B OR2X1_LOC_771/B 0.10fF
C12603 AND2X1_LOC_859/Y AND2X1_LOC_287/B 0.12fF
C12604 AND2X1_LOC_214/A OR2X1_LOC_59/Y 0.12fF
C12605 AND2X1_LOC_67/Y OR2X1_LOC_130/a_8_216# 0.47fF
C12606 OR2X1_LOC_650/Y OR2X1_LOC_771/B 0.18fF
C12607 AND2X1_LOC_63/a_8_24# OR2X1_LOC_161/B 0.01fF
C12608 OR2X1_LOC_51/Y OR2X1_LOC_517/A 0.01fF
C12609 OR2X1_LOC_185/Y OR2X1_LOC_576/A 0.02fF
C12610 AND2X1_LOC_363/Y AND2X1_LOC_344/a_8_24# 0.01fF
C12611 OR2X1_LOC_535/A AND2X1_LOC_43/B 0.05fF
C12612 AND2X1_LOC_72/B OR2X1_LOC_675/Y 0.02fF
C12613 AND2X1_LOC_311/a_8_24# OR2X1_LOC_538/A 0.00fF
C12614 AND2X1_LOC_859/Y OR2X1_LOC_816/A 0.07fF
C12615 AND2X1_LOC_861/B OR2X1_LOC_59/Y 0.36fF
C12616 AND2X1_LOC_588/B AND2X1_LOC_44/a_8_24# 0.19fF
C12617 OR2X1_LOC_306/Y OR2X1_LOC_829/A 0.15fF
C12618 OR2X1_LOC_600/A OR2X1_LOC_586/Y 0.05fF
C12619 AND2X1_LOC_564/B OR2X1_LOC_238/Y 0.01fF
C12620 OR2X1_LOC_190/A OR2X1_LOC_147/B 0.03fF
C12621 AND2X1_LOC_596/a_8_24# OR2X1_LOC_48/B 0.02fF
C12622 OR2X1_LOC_155/a_8_216# OR2X1_LOC_160/A 0.02fF
C12623 OR2X1_LOC_529/a_36_216# AND2X1_LOC_541/Y 0.01fF
C12624 AND2X1_LOC_392/A AND2X1_LOC_661/a_8_24# 0.04fF
C12625 AND2X1_LOC_731/a_36_24# AND2X1_LOC_191/Y 0.01fF
C12626 AND2X1_LOC_707/Y OR2X1_LOC_423/a_36_216# 0.01fF
C12627 OR2X1_LOC_585/A AND2X1_LOC_407/a_8_24# 0.01fF
C12628 AND2X1_LOC_40/Y OR2X1_LOC_78/A 0.20fF
C12629 OR2X1_LOC_51/Y AND2X1_LOC_833/a_8_24# 0.01fF
C12630 D_INPUT_1 AND2X1_LOC_236/a_8_24# 0.02fF
C12631 AND2X1_LOC_596/a_8_24# OR2X1_LOC_18/Y 0.02fF
C12632 AND2X1_LOC_326/B AND2X1_LOC_520/Y 0.00fF
C12633 OR2X1_LOC_663/A AND2X1_LOC_41/A 0.03fF
C12634 AND2X1_LOC_571/A AND2X1_LOC_523/Y 0.03fF
C12635 OR2X1_LOC_364/A OR2X1_LOC_439/B 0.01fF
C12636 OR2X1_LOC_756/B OR2X1_LOC_571/a_36_216# 0.00fF
C12637 AND2X1_LOC_40/Y D_GATE_741 0.04fF
C12638 AND2X1_LOC_339/Y AND2X1_LOC_339/a_8_24# 0.00fF
C12639 OR2X1_LOC_696/A AND2X1_LOC_849/A 0.01fF
C12640 VDD OR2X1_LOC_240/B 0.21fF
C12641 OR2X1_LOC_790/B VDD 0.00fF
C12642 AND2X1_LOC_785/a_36_24# OR2X1_LOC_70/Y 0.01fF
C12643 AND2X1_LOC_31/Y OR2X1_LOC_374/Y 0.04fF
C12644 OR2X1_LOC_158/A OR2X1_LOC_669/A 0.41fF
C12645 AND2X1_LOC_48/A OR2X1_LOC_598/a_8_216# 0.09fF
C12646 AND2X1_LOC_95/Y OR2X1_LOC_542/B 0.00fF
C12647 OR2X1_LOC_49/A OR2X1_LOC_240/A 0.07fF
C12648 OR2X1_LOC_160/A AND2X1_LOC_18/Y 0.54fF
C12649 AND2X1_LOC_339/B OR2X1_LOC_43/A 0.03fF
C12650 OR2X1_LOC_680/A AND2X1_LOC_778/Y 0.46fF
C12651 OR2X1_LOC_460/B VDD 0.00fF
C12652 VDD OR2X1_LOC_161/A 2.66fF
C12653 OR2X1_LOC_604/A AND2X1_LOC_470/B 0.01fF
C12654 VDD AND2X1_LOC_453/Y -0.00fF
C12655 OR2X1_LOC_379/Y AND2X1_LOC_70/Y 0.02fF
C12656 OR2X1_LOC_496/a_8_216# AND2X1_LOC_621/Y 0.04fF
C12657 OR2X1_LOC_756/B OR2X1_LOC_392/A 0.00fF
C12658 OR2X1_LOC_160/B OR2X1_LOC_659/a_8_216# 0.01fF
C12659 AND2X1_LOC_12/Y OR2X1_LOC_66/A 0.27fF
C12660 OR2X1_LOC_158/A AND2X1_LOC_818/a_8_24# 0.02fF
C12661 OR2X1_LOC_764/Y OR2X1_LOC_12/Y 0.01fF
C12662 OR2X1_LOC_312/Y OR2X1_LOC_322/a_8_216# 0.01fF
C12663 OR2X1_LOC_670/a_36_216# OR2X1_LOC_9/Y 0.00fF
C12664 AND2X1_LOC_539/Y AND2X1_LOC_856/B 0.01fF
C12665 OR2X1_LOC_670/a_8_216# OR2X1_LOC_40/Y 0.08fF
C12666 OR2X1_LOC_506/A AND2X1_LOC_92/Y 0.03fF
C12667 AND2X1_LOC_357/A OR2X1_LOC_36/Y 0.04fF
C12668 OR2X1_LOC_132/a_8_216# OR2X1_LOC_65/B 0.02fF
C12669 OR2X1_LOC_51/Y AND2X1_LOC_624/A 0.13fF
C12670 AND2X1_LOC_541/Y AND2X1_LOC_361/A 0.03fF
C12671 OR2X1_LOC_158/A AND2X1_LOC_454/A 0.04fF
C12672 OR2X1_LOC_831/A OR2X1_LOC_155/A 0.17fF
C12673 OR2X1_LOC_158/A OR2X1_LOC_232/a_8_216# 0.07fF
C12674 AND2X1_LOC_92/Y OR2X1_LOC_341/Y 0.03fF
C12675 OR2X1_LOC_406/a_8_216# AND2X1_LOC_657/Y 0.28fF
C12676 OR2X1_LOC_154/A AND2X1_LOC_172/a_8_24# 0.00fF
C12677 VDD AND2X1_LOC_25/Y 0.33fF
C12678 OR2X1_LOC_6/B OR2X1_LOC_83/A 0.02fF
C12679 OR2X1_LOC_62/B OR2X1_LOC_115/B 0.02fF
C12680 AND2X1_LOC_218/Y OR2X1_LOC_39/A 0.02fF
C12681 OR2X1_LOC_155/A OR2X1_LOC_515/A 0.03fF
C12682 OR2X1_LOC_3/Y OR2X1_LOC_381/a_8_216# 0.11fF
C12683 OR2X1_LOC_748/A OR2X1_LOC_600/A 0.06fF
C12684 OR2X1_LOC_380/A OR2X1_LOC_51/Y 0.03fF
C12685 OR2X1_LOC_598/Y OR2X1_LOC_155/A 0.30fF
C12686 OR2X1_LOC_750/Y OR2X1_LOC_789/A 0.00fF
C12687 AND2X1_LOC_180/a_8_24# OR2X1_LOC_74/A 0.04fF
C12688 OR2X1_LOC_61/Y OR2X1_LOC_475/B 0.10fF
C12689 OR2X1_LOC_803/a_8_216# OR2X1_LOC_803/B 0.02fF
C12690 AND2X1_LOC_307/Y OR2X1_LOC_428/A 0.05fF
C12691 VDD OR2X1_LOC_26/Y 1.48fF
C12692 OR2X1_LOC_841/B OR2X1_LOC_841/A 0.20fF
C12693 OR2X1_LOC_114/Y AND2X1_LOC_70/Y 0.00fF
C12694 OR2X1_LOC_574/A OR2X1_LOC_631/A 0.04fF
C12695 AND2X1_LOC_95/Y OR2X1_LOC_736/A 0.04fF
C12696 OR2X1_LOC_744/A AND2X1_LOC_319/A 0.03fF
C12697 AND2X1_LOC_802/a_8_24# AND2X1_LOC_802/Y 0.03fF
C12698 AND2X1_LOC_174/a_8_24# AND2X1_LOC_857/Y 0.01fF
C12699 OR2X1_LOC_239/Y AND2X1_LOC_500/B 0.00fF
C12700 AND2X1_LOC_845/Y OR2X1_LOC_89/Y 0.07fF
C12701 AND2X1_LOC_711/a_36_24# AND2X1_LOC_848/Y 0.01fF
C12702 AND2X1_LOC_714/B OR2X1_LOC_70/Y 0.01fF
C12703 OR2X1_LOC_3/Y AND2X1_LOC_448/a_8_24# 0.00fF
C12704 OR2X1_LOC_662/A OR2X1_LOC_663/A 0.01fF
C12705 OR2X1_LOC_40/Y AND2X1_LOC_554/B 0.01fF
C12706 OR2X1_LOC_40/Y OR2X1_LOC_680/Y 0.03fF
C12707 AND2X1_LOC_160/Y OR2X1_LOC_52/B 0.13fF
C12708 AND2X1_LOC_577/a_8_24# AND2X1_LOC_577/A 0.07fF
C12709 OR2X1_LOC_458/a_36_216# OR2X1_LOC_805/A 0.02fF
C12710 VDD AND2X1_LOC_349/B 0.08fF
C12711 AND2X1_LOC_86/B AND2X1_LOC_18/Y 0.01fF
C12712 AND2X1_LOC_711/a_8_24# OR2X1_LOC_748/A 0.00fF
C12713 VDD OR2X1_LOC_89/A 0.78fF
C12714 OR2X1_LOC_857/B OR2X1_LOC_857/a_8_216# 0.00fF
C12715 OR2X1_LOC_160/A OR2X1_LOC_473/a_8_216# 0.06fF
C12716 OR2X1_LOC_850/B OR2X1_LOC_805/A 0.23fF
C12717 OR2X1_LOC_203/Y AND2X1_LOC_628/a_36_24# 0.01fF
C12718 VDD AND2X1_LOC_525/a_8_24# -0.00fF
C12719 OR2X1_LOC_185/Y AND2X1_LOC_41/A 0.16fF
C12720 AND2X1_LOC_79/Y OR2X1_LOC_66/A 0.03fF
C12721 OR2X1_LOC_624/B AND2X1_LOC_18/Y 0.18fF
C12722 OR2X1_LOC_516/A AND2X1_LOC_486/Y 0.03fF
C12723 VDD OR2X1_LOC_820/Y 0.06fF
C12724 OR2X1_LOC_703/B OR2X1_LOC_502/A 0.01fF
C12725 OR2X1_LOC_235/B OR2X1_LOC_849/A 0.01fF
C12726 AND2X1_LOC_645/A OR2X1_LOC_59/Y 0.02fF
C12727 OR2X1_LOC_40/Y AND2X1_LOC_326/A 0.02fF
C12728 AND2X1_LOC_699/a_8_24# AND2X1_LOC_36/Y 0.02fF
C12729 OR2X1_LOC_743/A OR2X1_LOC_56/A 0.06fF
C12730 AND2X1_LOC_80/a_36_24# OR2X1_LOC_502/A 0.00fF
C12731 VDD OR2X1_LOC_461/Y 0.00fF
C12732 OR2X1_LOC_756/B OR2X1_LOC_592/a_8_216# 0.01fF
C12733 OR2X1_LOC_502/A OR2X1_LOC_87/A 0.14fF
C12734 OR2X1_LOC_677/Y OR2X1_LOC_26/Y 0.02fF
C12735 AND2X1_LOC_36/Y OR2X1_LOC_675/Y 0.02fF
C12736 VDD AND2X1_LOC_51/Y 2.52fF
C12737 OR2X1_LOC_532/B OR2X1_LOC_355/a_8_216# 0.01fF
C12738 INPUT_5 OR2X1_LOC_588/Y 0.03fF
C12739 OR2X1_LOC_651/a_8_216# D_INPUT_5 0.01fF
C12740 AND2X1_LOC_724/Y OR2X1_LOC_64/Y 0.02fF
C12741 OR2X1_LOC_36/Y AND2X1_LOC_852/B 0.17fF
C12742 OR2X1_LOC_502/A AND2X1_LOC_696/a_8_24# 0.03fF
C12743 OR2X1_LOC_697/Y OR2X1_LOC_7/A 0.03fF
C12744 OR2X1_LOC_117/Y OR2X1_LOC_92/Y 0.15fF
C12745 INPUT_0 AND2X1_LOC_4/a_8_24# 0.04fF
C12746 OR2X1_LOC_313/Y AND2X1_LOC_452/Y 0.17fF
C12747 AND2X1_LOC_191/B OR2X1_LOC_488/a_36_216# 0.01fF
C12748 AND2X1_LOC_140/a_8_24# OR2X1_LOC_744/A 0.01fF
C12749 OR2X1_LOC_244/A AND2X1_LOC_65/A 0.01fF
C12750 OR2X1_LOC_475/Y OR2X1_LOC_78/A 0.01fF
C12751 OR2X1_LOC_160/A OR2X1_LOC_500/A 0.01fF
C12752 AND2X1_LOC_40/Y OR2X1_LOC_155/A 2.28fF
C12753 OR2X1_LOC_677/Y OR2X1_LOC_89/A 0.03fF
C12754 AND2X1_LOC_753/a_8_24# OR2X1_LOC_193/Y 0.23fF
C12755 AND2X1_LOC_467/a_8_24# AND2X1_LOC_470/B 0.01fF
C12756 AND2X1_LOC_741/Y AND2X1_LOC_479/Y 0.00fF
C12757 OR2X1_LOC_36/Y OR2X1_LOC_48/B 0.15fF
C12758 OR2X1_LOC_810/A OR2X1_LOC_785/B 0.07fF
C12759 OR2X1_LOC_316/Y AND2X1_LOC_318/a_8_24# 0.11fF
C12760 AND2X1_LOC_95/Y AND2X1_LOC_56/B 9.31fF
C12761 OR2X1_LOC_132/Y AND2X1_LOC_663/B 0.11fF
C12762 AND2X1_LOC_711/Y AND2X1_LOC_861/B 0.39fF
C12763 OR2X1_LOC_680/A AND2X1_LOC_624/A 0.08fF
C12764 OR2X1_LOC_160/B AND2X1_LOC_23/a_8_24# 0.01fF
C12765 AND2X1_LOC_40/Y OR2X1_LOC_807/a_8_216# 0.01fF
C12766 AND2X1_LOC_95/Y OR2X1_LOC_659/B 0.02fF
C12767 OR2X1_LOC_18/Y OR2X1_LOC_36/Y 1.09fF
C12768 VDD OR2X1_LOC_836/Y -0.00fF
C12769 OR2X1_LOC_154/A OR2X1_LOC_539/Y 0.06fF
C12770 OR2X1_LOC_181/Y OR2X1_LOC_367/B 0.80fF
C12771 INPUT_0 OR2X1_LOC_5/a_8_216# 0.01fF
C12772 AND2X1_LOC_784/A AND2X1_LOC_662/B 0.07fF
C12773 OR2X1_LOC_49/A OR2X1_LOC_47/Y 0.07fF
C12774 OR2X1_LOC_790/A AND2X1_LOC_47/Y 0.01fF
C12775 OR2X1_LOC_87/A AND2X1_LOC_230/a_8_24# 0.02fF
C12776 AND2X1_LOC_216/A AND2X1_LOC_772/Y 0.01fF
C12777 AND2X1_LOC_859/Y AND2X1_LOC_843/a_8_24# 0.01fF
C12778 AND2X1_LOC_792/Y GATE_579 0.00fF
C12779 AND2X1_LOC_95/Y AND2X1_LOC_8/Y 0.04fF
C12780 AND2X1_LOC_727/A AND2X1_LOC_468/a_8_24# 0.01fF
C12781 AND2X1_LOC_866/A AND2X1_LOC_476/Y 0.07fF
C12782 GATE_741 GATE_811 0.28fF
C12783 OR2X1_LOC_246/A OR2X1_LOC_56/A 0.01fF
C12784 OR2X1_LOC_130/A OR2X1_LOC_222/A 0.21fF
C12785 AND2X1_LOC_362/B AND2X1_LOC_866/A 0.15fF
C12786 OR2X1_LOC_69/A OR2X1_LOC_44/Y 0.02fF
C12787 AND2X1_LOC_95/Y OR2X1_LOC_720/a_36_216# 0.00fF
C12788 OR2X1_LOC_160/A OR2X1_LOC_469/a_8_216# 0.01fF
C12789 OR2X1_LOC_633/Y AND2X1_LOC_8/Y 0.03fF
C12790 AND2X1_LOC_859/Y AND2X1_LOC_807/Y 0.02fF
C12791 OR2X1_LOC_860/a_36_216# OR2X1_LOC_287/B 0.00fF
C12792 OR2X1_LOC_862/B OR2X1_LOC_814/A 0.33fF
C12793 AND2X1_LOC_717/Y OR2X1_LOC_371/Y 0.00fF
C12794 AND2X1_LOC_59/Y OR2X1_LOC_719/Y 0.01fF
C12795 D_INPUT_7 AND2X1_LOC_11/Y 0.27fF
C12796 OR2X1_LOC_315/Y OR2X1_LOC_26/Y 0.00fF
C12797 OR2X1_LOC_368/a_8_216# OR2X1_LOC_95/Y 0.00fF
C12798 OR2X1_LOC_213/A OR2X1_LOC_87/A 0.01fF
C12799 OR2X1_LOC_32/B OR2X1_LOC_690/A 0.01fF
C12800 OR2X1_LOC_437/A OR2X1_LOC_142/Y 0.06fF
C12801 OR2X1_LOC_194/Y OR2X1_LOC_193/Y 0.12fF
C12802 AND2X1_LOC_342/Y OR2X1_LOC_248/Y 0.17fF
C12803 AND2X1_LOC_477/A OR2X1_LOC_59/Y 0.03fF
C12804 AND2X1_LOC_86/Y OR2X1_LOC_204/a_8_216# 0.03fF
C12805 OR2X1_LOC_112/A OR2X1_LOC_174/Y 0.27fF
C12806 OR2X1_LOC_634/A OR2X1_LOC_46/A 0.35fF
C12807 OR2X1_LOC_45/B OR2X1_LOC_406/A 0.00fF
C12808 OR2X1_LOC_858/A OR2X1_LOC_532/B 0.02fF
C12809 AND2X1_LOC_801/B AND2X1_LOC_434/Y 0.01fF
C12810 OR2X1_LOC_699/a_8_216# OR2X1_LOC_43/A 0.03fF
C12811 AND2X1_LOC_858/B OR2X1_LOC_226/a_8_216# 0.25fF
C12812 OR2X1_LOC_114/Y OR2X1_LOC_116/a_8_216# 0.07fF
C12813 OR2X1_LOC_26/Y AND2X1_LOC_267/a_8_24# 0.01fF
C12814 AND2X1_LOC_63/a_36_24# AND2X1_LOC_8/Y 0.00fF
C12815 AND2X1_LOC_72/B OR2X1_LOC_736/Y 0.04fF
C12816 AND2X1_LOC_390/B OR2X1_LOC_829/a_36_216# 0.01fF
C12817 AND2X1_LOC_31/Y OR2X1_LOC_392/B 0.03fF
C12818 OR2X1_LOC_95/Y AND2X1_LOC_468/a_8_24# 0.04fF
C12819 AND2X1_LOC_170/a_36_24# AND2X1_LOC_566/Y 0.01fF
C12820 AND2X1_LOC_362/a_8_24# OR2X1_LOC_417/A 0.03fF
C12821 OR2X1_LOC_744/A AND2X1_LOC_170/B 0.03fF
C12822 AND2X1_LOC_578/A OR2X1_LOC_39/A 0.14fF
C12823 OR2X1_LOC_185/A OR2X1_LOC_254/a_8_216# 0.01fF
C12824 OR2X1_LOC_251/Y OR2X1_LOC_26/Y 0.01fF
C12825 AND2X1_LOC_580/A OR2X1_LOC_74/A 5.55fF
C12826 OR2X1_LOC_95/Y OR2X1_LOC_597/a_36_216# 0.00fF
C12827 OR2X1_LOC_256/Y OR2X1_LOC_255/a_8_216# 0.48fF
C12828 OR2X1_LOC_48/Y OR2X1_LOC_48/a_8_216# 0.01fF
C12829 OR2X1_LOC_491/Y AND2X1_LOC_493/a_8_24# 0.23fF
C12830 OR2X1_LOC_491/Y OR2X1_LOC_89/A 0.07fF
C12831 OR2X1_LOC_656/B OR2X1_LOC_656/a_36_216# 0.00fF
C12832 OR2X1_LOC_277/a_36_216# AND2X1_LOC_573/A 0.01fF
C12833 AND2X1_LOC_345/a_8_24# OR2X1_LOC_44/Y 0.01fF
C12834 AND2X1_LOC_733/Y AND2X1_LOC_675/A 0.00fF
C12835 OR2X1_LOC_860/a_8_216# OR2X1_LOC_859/A 0.10fF
C12836 OR2X1_LOC_251/Y OR2X1_LOC_89/A 0.05fF
C12837 AND2X1_LOC_578/A AND2X1_LOC_569/a_8_24# 0.03fF
C12838 AND2X1_LOC_638/Y OR2X1_LOC_409/B 0.31fF
C12839 OR2X1_LOC_136/a_8_216# OR2X1_LOC_437/A 0.03fF
C12840 OR2X1_LOC_759/A AND2X1_LOC_805/a_8_24# 0.01fF
C12841 OR2X1_LOC_98/a_8_216# OR2X1_LOC_66/A -0.00fF
C12842 AND2X1_LOC_22/Y OR2X1_LOC_446/B 0.03fF
C12843 OR2X1_LOC_754/A OR2X1_LOC_753/A 0.17fF
C12844 VDD OR2X1_LOC_551/B 0.05fF
C12845 OR2X1_LOC_804/a_36_216# OR2X1_LOC_223/A 0.00fF
C12846 OR2X1_LOC_114/Y OR2X1_LOC_404/Y 0.01fF
C12847 OR2X1_LOC_744/A AND2X1_LOC_721/A 0.03fF
C12848 AND2X1_LOC_580/B OR2X1_LOC_755/A 0.13fF
C12849 AND2X1_LOC_22/Y OR2X1_LOC_303/B 0.57fF
C12850 OR2X1_LOC_441/a_8_216# OR2X1_LOC_47/Y 0.14fF
C12851 OR2X1_LOC_94/a_8_216# OR2X1_LOC_46/A 0.03fF
C12852 OR2X1_LOC_271/Y AND2X1_LOC_523/Y 0.00fF
C12853 OR2X1_LOC_500/a_8_216# OR2X1_LOC_501/A -0.00fF
C12854 OR2X1_LOC_439/B OR2X1_LOC_578/B 0.36fF
C12855 OR2X1_LOC_70/Y AND2X1_LOC_645/A 0.12fF
C12856 OR2X1_LOC_836/B AND2X1_LOC_51/Y 0.34fF
C12857 OR2X1_LOC_175/Y OR2X1_LOC_332/a_8_216# 0.39fF
C12858 AND2X1_LOC_303/A OR2X1_LOC_46/A 0.12fF
C12859 OR2X1_LOC_754/A OR2X1_LOC_754/a_8_216# 0.13fF
C12860 OR2X1_LOC_471/Y OR2X1_LOC_210/a_8_216# 0.14fF
C12861 OR2X1_LOC_485/A OR2X1_LOC_279/a_36_216# 0.01fF
C12862 OR2X1_LOC_22/A AND2X1_LOC_459/Y 0.00fF
C12863 OR2X1_LOC_652/a_36_216# OR2X1_LOC_814/A 0.05fF
C12864 AND2X1_LOC_729/Y AND2X1_LOC_800/a_8_24# 0.01fF
C12865 OR2X1_LOC_519/Y AND2X1_LOC_831/Y 0.01fF
C12866 AND2X1_LOC_48/A OR2X1_LOC_87/A 0.02fF
C12867 AND2X1_LOC_724/A AND2X1_LOC_592/a_8_24# 0.20fF
C12868 OR2X1_LOC_52/Y OR2X1_LOC_585/A 0.07fF
C12869 OR2X1_LOC_696/Y OR2X1_LOC_7/A 0.01fF
C12870 AND2X1_LOC_185/a_8_24# AND2X1_LOC_620/Y 0.01fF
C12871 OR2X1_LOC_405/A OR2X1_LOC_436/Y 0.03fF
C12872 OR2X1_LOC_62/B OR2X1_LOC_6/A 0.02fF
C12873 OR2X1_LOC_287/B AND2X1_LOC_77/a_8_24# -0.00fF
C12874 OR2X1_LOC_248/Y OR2X1_LOC_54/Y 0.00fF
C12875 OR2X1_LOC_91/Y OR2X1_LOC_71/Y 0.03fF
C12876 AND2X1_LOC_44/Y OR2X1_LOC_217/A 0.17fF
C12877 OR2X1_LOC_161/B OR2X1_LOC_141/a_8_216# 0.01fF
C12878 AND2X1_LOC_25/a_8_24# AND2X1_LOC_25/Y 0.00fF
C12879 D_INPUT_3 AND2X1_LOC_820/a_36_24# 0.00fF
C12880 AND2X1_LOC_831/Y AND2X1_LOC_139/B 0.08fF
C12881 AND2X1_LOC_508/A OR2X1_LOC_419/Y 0.00fF
C12882 OR2X1_LOC_864/A OR2X1_LOC_649/a_36_216# 0.00fF
C12883 OR2X1_LOC_201/Y OR2X1_LOC_206/a_8_216# 0.00fF
C12884 OR2X1_LOC_835/Y AND2X1_LOC_823/a_8_24# 0.02fF
C12885 OR2X1_LOC_64/Y OR2X1_LOC_371/Y 0.15fF
C12886 OR2X1_LOC_269/A OR2X1_LOC_719/B 0.02fF
C12887 OR2X1_LOC_276/B OR2X1_LOC_541/B 0.01fF
C12888 OR2X1_LOC_580/A OR2X1_LOC_343/a_8_216# 0.01fF
C12889 AND2X1_LOC_69/a_36_24# OR2X1_LOC_87/A 0.00fF
C12890 OR2X1_LOC_62/A OR2X1_LOC_38/a_8_216# -0.03fF
C12891 INPUT_0 AND2X1_LOC_222/Y 0.01fF
C12892 OR2X1_LOC_744/A OR2X1_LOC_331/Y 0.03fF
C12893 AND2X1_LOC_319/A OR2X1_LOC_31/Y 0.03fF
C12894 OR2X1_LOC_241/Y OR2X1_LOC_130/A 0.01fF
C12895 OR2X1_LOC_589/A OR2X1_LOC_300/Y 0.04fF
C12896 OR2X1_LOC_429/Y AND2X1_LOC_635/a_8_24# 0.02fF
C12897 OR2X1_LOC_485/A OR2X1_LOC_46/A 0.02fF
C12898 AND2X1_LOC_821/a_8_24# OR2X1_LOC_269/B 0.03fF
C12899 INPUT_0 OR2X1_LOC_68/B 1.35fF
C12900 OR2X1_LOC_256/A OR2X1_LOC_26/Y 0.03fF
C12901 OR2X1_LOC_744/A AND2X1_LOC_217/a_8_24# 0.01fF
C12902 AND2X1_LOC_52/a_8_24# AND2X1_LOC_52/Y 0.01fF
C12903 OR2X1_LOC_510/Y OR2X1_LOC_786/Y 0.03fF
C12904 OR2X1_LOC_736/Y AND2X1_LOC_36/Y 0.03fF
C12905 OR2X1_LOC_334/a_8_216# OR2X1_LOC_338/A 0.01fF
C12906 OR2X1_LOC_18/Y OR2X1_LOC_85/a_8_216# 0.03fF
C12907 OR2X1_LOC_120/a_8_216# OR2X1_LOC_121/A 0.01fF
C12908 OR2X1_LOC_614/Y AND2X1_LOC_36/Y 0.26fF
C12909 OR2X1_LOC_739/A OR2X1_LOC_330/a_36_216# 0.00fF
C12910 OR2X1_LOC_70/Y AND2X1_LOC_477/A 0.06fF
C12911 OR2X1_LOC_256/A OR2X1_LOC_89/A 0.05fF
C12912 OR2X1_LOC_18/Y OR2X1_LOC_419/Y 0.05fF
C12913 OR2X1_LOC_689/Y OR2X1_LOC_585/A 0.01fF
C12914 OR2X1_LOC_244/A OR2X1_LOC_204/a_8_216# 0.04fF
C12915 AND2X1_LOC_717/Y AND2X1_LOC_222/Y 0.03fF
C12916 OR2X1_LOC_417/A OR2X1_LOC_371/Y 0.07fF
C12917 OR2X1_LOC_47/Y AND2X1_LOC_661/A 0.03fF
C12918 OR2X1_LOC_485/A AND2X1_LOC_227/Y 0.03fF
C12919 OR2X1_LOC_36/Y AND2X1_LOC_620/Y 0.03fF
C12920 OR2X1_LOC_51/B OR2X1_LOC_44/Y 0.01fF
C12921 OR2X1_LOC_92/Y AND2X1_LOC_790/a_36_24# 0.00fF
C12922 AND2X1_LOC_785/a_8_24# AND2X1_LOC_786/Y 0.02fF
C12923 AND2X1_LOC_773/Y AND2X1_LOC_773/a_8_24# 0.00fF
C12924 OR2X1_LOC_323/A OR2X1_LOC_323/Y 0.02fF
C12925 OR2X1_LOC_810/A OR2X1_LOC_786/Y 0.12fF
C12926 OR2X1_LOC_74/A AND2X1_LOC_476/A 0.07fF
C12927 OR2X1_LOC_31/Y OR2X1_LOC_52/a_8_216# 0.01fF
C12928 AND2X1_LOC_514/Y AND2X1_LOC_477/A 0.16fF
C12929 OR2X1_LOC_611/a_36_216# OR2X1_LOC_62/B 0.00fF
C12930 OR2X1_LOC_494/A OR2X1_LOC_428/A 0.01fF
C12931 OR2X1_LOC_393/a_8_216# OR2X1_LOC_80/A 0.10fF
C12932 OR2X1_LOC_475/B AND2X1_LOC_406/a_8_24# 0.01fF
C12933 AND2X1_LOC_362/a_36_24# OR2X1_LOC_13/B 0.00fF
C12934 OR2X1_LOC_641/Y AND2X1_LOC_36/Y 0.19fF
C12935 OR2X1_LOC_175/Y OR2X1_LOC_161/B 0.07fF
C12936 OR2X1_LOC_26/Y OR2X1_LOC_67/Y 0.06fF
C12937 OR2X1_LOC_201/a_8_216# OR2X1_LOC_206/a_8_216# 0.47fF
C12938 AND2X1_LOC_7/B OR2X1_LOC_138/A 0.02fF
C12939 AND2X1_LOC_48/A OR2X1_LOC_706/B 0.01fF
C12940 OR2X1_LOC_158/A AND2X1_LOC_783/B 0.01fF
C12941 OR2X1_LOC_696/A OR2X1_LOC_93/Y 0.01fF
C12942 OR2X1_LOC_88/a_8_216# OR2X1_LOC_39/A 0.01fF
C12943 OR2X1_LOC_45/B OR2X1_LOC_505/a_8_216# 0.05fF
C12944 OR2X1_LOC_247/a_8_216# AND2X1_LOC_3/Y 0.01fF
C12945 D_INPUT_0 OR2X1_LOC_814/A 0.16fF
C12946 OR2X1_LOC_89/A AND2X1_LOC_624/B 0.02fF
C12947 OR2X1_LOC_416/Y OR2X1_LOC_75/a_8_216# 0.01fF
C12948 AND2X1_LOC_92/Y OR2X1_LOC_180/B 0.03fF
C12949 OR2X1_LOC_691/Y OR2X1_LOC_161/B 0.03fF
C12950 AND2X1_LOC_576/a_8_24# AND2X1_LOC_657/A 0.02fF
C12951 OR2X1_LOC_83/A OR2X1_LOC_598/A 0.02fF
C12952 AND2X1_LOC_387/B OR2X1_LOC_214/B 4.29fF
C12953 OR2X1_LOC_696/A AND2X1_LOC_447/Y 0.02fF
C12954 AND2X1_LOC_610/a_8_24# AND2X1_LOC_647/Y 0.20fF
C12955 OR2X1_LOC_66/A OR2X1_LOC_356/B 0.07fF
C12956 VDD AND2X1_LOC_590/a_8_24# -0.00fF
C12957 OR2X1_LOC_685/A AND2X1_LOC_31/Y 0.09fF
C12958 AND2X1_LOC_40/Y D_GATE_366 0.11fF
C12959 AND2X1_LOC_118/a_8_24# OR2X1_LOC_598/A 0.07fF
C12960 AND2X1_LOC_40/a_8_24# AND2X1_LOC_44/Y 0.01fF
C12961 OR2X1_LOC_62/A OR2X1_LOC_19/B 0.08fF
C12962 OR2X1_LOC_161/B OR2X1_LOC_713/A 0.15fF
C12963 OR2X1_LOC_696/A OR2X1_LOC_380/Y 0.12fF
C12964 OR2X1_LOC_196/Y AND2X1_LOC_754/a_36_24# 0.00fF
C12965 OR2X1_LOC_527/a_8_216# AND2X1_LOC_721/Y 0.01fF
C12966 AND2X1_LOC_655/a_8_24# OR2X1_LOC_46/A 0.01fF
C12967 OR2X1_LOC_808/B AND2X1_LOC_36/Y 0.03fF
C12968 OR2X1_LOC_186/Y OR2X1_LOC_486/Y 0.07fF
C12969 AND2X1_LOC_727/A AND2X1_LOC_798/A 0.01fF
C12970 OR2X1_LOC_485/A OR2X1_LOC_753/Y 0.02fF
C12971 OR2X1_LOC_710/A OR2X1_LOC_78/A 0.01fF
C12972 AND2X1_LOC_715/Y AND2X1_LOC_447/Y 0.02fF
C12973 OR2X1_LOC_690/A OR2X1_LOC_68/B 0.28fF
C12974 OR2X1_LOC_45/B AND2X1_LOC_725/a_8_24# 0.02fF
C12975 OR2X1_LOC_177/a_8_216# AND2X1_LOC_476/Y 0.04fF
C12976 OR2X1_LOC_249/Y OR2X1_LOC_580/A 0.00fF
C12977 OR2X1_LOC_46/A OR2X1_LOC_609/Y 0.01fF
C12978 OR2X1_LOC_266/A AND2X1_LOC_18/Y 0.01fF
C12979 D_INPUT_3 OR2X1_LOC_71/Y 0.17fF
C12980 OR2X1_LOC_831/B OR2X1_LOC_778/B 0.08fF
C12981 AND2X1_LOC_645/A OR2X1_LOC_534/a_36_216# 0.00fF
C12982 AND2X1_LOC_56/B OR2X1_LOC_269/A 0.01fF
C12983 OR2X1_LOC_160/B AND2X1_LOC_603/a_8_24# 0.05fF
C12984 AND2X1_LOC_841/a_36_24# OR2X1_LOC_417/A -0.01fF
C12985 OR2X1_LOC_571/B OR2X1_LOC_579/A 0.02fF
C12986 OR2X1_LOC_857/A OR2X1_LOC_35/Y 0.04fF
C12987 AND2X1_LOC_570/Y AND2X1_LOC_456/a_36_24# 0.00fF
C12988 OR2X1_LOC_158/A AND2X1_LOC_285/a_36_24# 0.00fF
C12989 OR2X1_LOC_502/A OR2X1_LOC_390/B 0.08fF
C12990 AND2X1_LOC_436/Y AND2X1_LOC_802/Y 0.03fF
C12991 OR2X1_LOC_620/Y OR2X1_LOC_319/Y 0.01fF
C12992 AND2X1_LOC_564/A OR2X1_LOC_524/Y 0.07fF
C12993 OR2X1_LOC_40/Y AND2X1_LOC_476/Y 0.03fF
C12994 OR2X1_LOC_64/Y AND2X1_LOC_222/Y 0.06fF
C12995 AND2X1_LOC_18/Y AND2X1_LOC_607/a_8_24# 0.03fF
C12996 AND2X1_LOC_515/a_36_24# OR2X1_LOC_600/A 0.00fF
C12997 OR2X1_LOC_308/A OR2X1_LOC_512/A 0.47fF
C12998 VDD AND2X1_LOC_605/a_8_24# 0.00fF
C12999 AND2X1_LOC_552/A VDD 0.25fF
C13000 OR2X1_LOC_235/B OR2X1_LOC_721/a_8_216# 0.01fF
C13001 OR2X1_LOC_516/Y AND2X1_LOC_621/Y 0.07fF
C13002 OR2X1_LOC_696/A OR2X1_LOC_109/Y 0.06fF
C13003 OR2X1_LOC_112/a_8_216# OR2X1_LOC_809/B 0.03fF
C13004 D_INPUT_3 D_INPUT_1 0.04fF
C13005 OR2X1_LOC_47/Y OR2X1_LOC_760/Y 0.01fF
C13006 VDD AND2X1_LOC_194/Y 0.01fF
C13007 OR2X1_LOC_155/A OR2X1_LOC_707/a_36_216# 0.00fF
C13008 OR2X1_LOC_492/a_8_216# OR2X1_LOC_59/Y 0.06fF
C13009 OR2X1_LOC_19/B OR2X1_LOC_88/Y 0.01fF
C13010 OR2X1_LOC_78/A OR2X1_LOC_356/A 0.07fF
C13011 OR2X1_LOC_92/a_8_216# OR2X1_LOC_67/Y 0.05fF
C13012 OR2X1_LOC_708/Y AND2X1_LOC_44/Y 0.01fF
C13013 OR2X1_LOC_607/a_8_216# AND2X1_LOC_647/Y 0.01fF
C13014 OR2X1_LOC_188/Y OR2X1_LOC_147/B 0.03fF
C13015 AND2X1_LOC_64/Y AND2X1_LOC_504/a_8_24# 0.01fF
C13016 OR2X1_LOC_44/Y AND2X1_LOC_792/B 0.21fF
C13017 OR2X1_LOC_329/a_8_216# OR2X1_LOC_329/B 0.04fF
C13018 OR2X1_LOC_190/A OR2X1_LOC_190/a_8_216# 0.03fF
C13019 OR2X1_LOC_114/B OR2X1_LOC_190/A 0.03fF
C13020 OR2X1_LOC_290/a_8_216# OR2X1_LOC_16/A 0.01fF
C13021 OR2X1_LOC_71/Y AND2X1_LOC_656/a_8_24# 0.01fF
C13022 AND2X1_LOC_605/Y OR2X1_LOC_604/Y 0.80fF
C13023 OR2X1_LOC_377/A OR2X1_LOC_415/Y 0.03fF
C13024 OR2X1_LOC_434/a_8_216# OR2X1_LOC_390/A 0.01fF
C13025 OR2X1_LOC_235/B OR2X1_LOC_673/a_36_216# 0.00fF
C13026 OR2X1_LOC_417/A AND2X1_LOC_222/Y 0.22fF
C13027 OR2X1_LOC_158/A AND2X1_LOC_162/a_36_24# 0.00fF
C13028 AND2X1_LOC_810/Y AND2X1_LOC_486/a_36_24# 0.00fF
C13029 OR2X1_LOC_532/B AND2X1_LOC_31/Y 7.61fF
C13030 OR2X1_LOC_151/A OR2X1_LOC_499/B 0.01fF
C13031 OR2X1_LOC_757/Y AND2X1_LOC_789/Y 0.02fF
C13032 OR2X1_LOC_756/B OR2X1_LOC_349/A 0.79fF
C13033 OR2X1_LOC_427/A OR2X1_LOC_428/A 0.28fF
C13034 OR2X1_LOC_629/Y OR2X1_LOC_161/B 0.02fF
C13035 OR2X1_LOC_96/Y OR2X1_LOC_91/A 0.05fF
C13036 AND2X1_LOC_76/Y AND2X1_LOC_455/B 0.04fF
C13037 AND2X1_LOC_507/a_36_24# OR2X1_LOC_56/A 0.00fF
C13038 AND2X1_LOC_717/B OR2X1_LOC_183/Y 0.07fF
C13039 OR2X1_LOC_269/B OR2X1_LOC_605/Y 0.03fF
C13040 OR2X1_LOC_635/A OR2X1_LOC_614/Y 0.02fF
C13041 OR2X1_LOC_614/a_36_216# OR2X1_LOC_78/A 0.03fF
C13042 OR2X1_LOC_185/A AND2X1_LOC_44/Y 0.17fF
C13043 OR2X1_LOC_375/A OR2X1_LOC_563/A 0.07fF
C13044 OR2X1_LOC_687/Y AND2X1_LOC_760/a_36_24# 0.00fF
C13045 AND2X1_LOC_160/Y AND2X1_LOC_161/Y 0.10fF
C13046 OR2X1_LOC_168/B OR2X1_LOC_66/A 0.03fF
C13047 OR2X1_LOC_416/Y OR2X1_LOC_13/B 0.03fF
C13048 AND2X1_LOC_3/Y OR2X1_LOC_598/a_8_216# 0.01fF
C13049 OR2X1_LOC_328/a_8_216# OR2X1_LOC_51/Y 0.01fF
C13050 OR2X1_LOC_653/Y OR2X1_LOC_390/A 0.01fF
C13051 AND2X1_LOC_84/Y OR2X1_LOC_6/A 0.10fF
C13052 OR2X1_LOC_269/Y OR2X1_LOC_675/Y 0.01fF
C13053 AND2X1_LOC_217/Y OR2X1_LOC_517/A 0.07fF
C13054 OR2X1_LOC_841/A OR2X1_LOC_168/B 0.01fF
C13055 OR2X1_LOC_327/a_8_216# AND2X1_LOC_65/A 0.01fF
C13056 OR2X1_LOC_177/Y OR2X1_LOC_48/B 0.02fF
C13057 OR2X1_LOC_98/B OR2X1_LOC_98/a_8_216# 0.01fF
C13058 AND2X1_LOC_482/a_8_24# OR2X1_LOC_549/A 0.01fF
C13059 OR2X1_LOC_151/A AND2X1_LOC_142/a_36_24# 0.00fF
C13060 OR2X1_LOC_689/A AND2X1_LOC_194/Y 0.03fF
C13061 OR2X1_LOC_67/Y AND2X1_LOC_202/a_8_24# 0.09fF
C13062 OR2X1_LOC_465/a_8_216# AND2X1_LOC_7/B 0.01fF
C13063 AND2X1_LOC_443/a_8_24# AND2X1_LOC_804/Y 0.20fF
C13064 AND2X1_LOC_612/B OR2X1_LOC_397/a_8_216# 0.47fF
C13065 OR2X1_LOC_177/Y OR2X1_LOC_18/Y 0.00fF
C13066 AND2X1_LOC_22/Y AND2X1_LOC_56/B 0.10fF
C13067 OR2X1_LOC_315/a_8_216# OR2X1_LOC_18/Y 0.01fF
C13068 VDD OR2X1_LOC_640/A 0.06fF
C13069 OR2X1_LOC_318/B OR2X1_LOC_241/B 0.18fF
C13070 OR2X1_LOC_7/A OR2X1_LOC_503/a_8_216# 0.01fF
C13071 OR2X1_LOC_549/B OR2X1_LOC_563/B 0.42fF
C13072 AND2X1_LOC_22/Y OR2X1_LOC_659/B 0.02fF
C13073 OR2X1_LOC_551/B OR2X1_LOC_551/A 0.08fF
C13074 OR2X1_LOC_840/A OR2X1_LOC_468/A 0.03fF
C13075 AND2X1_LOC_367/A OR2X1_LOC_122/A 0.08fF
C13076 OR2X1_LOC_92/Y AND2X1_LOC_614/a_36_24# 0.00fF
C13077 OR2X1_LOC_45/B AND2X1_LOC_702/Y 0.00fF
C13078 OR2X1_LOC_154/A OR2X1_LOC_691/A 0.00fF
C13079 OR2X1_LOC_85/A AND2X1_LOC_786/Y 0.06fF
C13080 AND2X1_LOC_64/Y OR2X1_LOC_557/A 0.03fF
C13081 OR2X1_LOC_538/a_36_216# AND2X1_LOC_70/Y 0.00fF
C13082 AND2X1_LOC_283/a_36_24# OR2X1_LOC_580/A 0.01fF
C13083 AND2X1_LOC_22/Y AND2X1_LOC_8/Y 0.06fF
C13084 OR2X1_LOC_207/B OR2X1_LOC_87/A 0.23fF
C13085 AND2X1_LOC_544/a_8_24# AND2X1_LOC_658/A 0.04fF
C13086 OR2X1_LOC_814/A OR2X1_LOC_339/A 0.08fF
C13087 AND2X1_LOC_540/a_8_24# OR2X1_LOC_178/Y 0.24fF
C13088 AND2X1_LOC_658/A AND2X1_LOC_866/B 0.01fF
C13089 OR2X1_LOC_696/A AND2X1_LOC_729/B 0.08fF
C13090 OR2X1_LOC_604/A OR2X1_LOC_48/B 0.05fF
C13091 OR2X1_LOC_508/a_8_216# AND2X1_LOC_81/B 0.01fF
C13092 D_INPUT_1 OR2X1_LOC_561/B 0.09fF
C13093 AND2X1_LOC_340/Y OR2X1_LOC_36/Y 0.03fF
C13094 OR2X1_LOC_528/a_8_216# AND2X1_LOC_807/Y 0.12fF
C13095 AND2X1_LOC_363/A OR2X1_LOC_428/A 0.00fF
C13096 OR2X1_LOC_823/a_8_216# OR2X1_LOC_96/Y 0.01fF
C13097 AND2X1_LOC_191/B OR2X1_LOC_92/Y 0.03fF
C13098 OR2X1_LOC_43/Y OR2X1_LOC_43/A 0.01fF
C13099 OR2X1_LOC_485/A AND2X1_LOC_227/a_36_24# 0.00fF
C13100 AND2X1_LOC_719/Y AND2X1_LOC_843/a_36_24# 0.01fF
C13101 OR2X1_LOC_847/A AND2X1_LOC_18/Y 0.00fF
C13102 OR2X1_LOC_179/Y AND2X1_LOC_181/a_8_24# 0.23fF
C13103 OR2X1_LOC_604/A OR2X1_LOC_18/Y 0.06fF
C13104 OR2X1_LOC_405/A OR2X1_LOC_160/B 0.07fF
C13105 AND2X1_LOC_706/Y OR2X1_LOC_599/A 0.00fF
C13106 AND2X1_LOC_550/a_8_24# AND2X1_LOC_550/A 0.03fF
C13107 OR2X1_LOC_8/Y OR2X1_LOC_278/Y 0.04fF
C13108 AND2X1_LOC_738/B OR2X1_LOC_525/Y 0.31fF
C13109 VDD AND2X1_LOC_297/a_8_24# 0.00fF
C13110 AND2X1_LOC_181/Y OR2X1_LOC_36/Y 0.03fF
C13111 OR2X1_LOC_406/Y AND2X1_LOC_711/Y 0.04fF
C13112 AND2X1_LOC_92/Y OR2X1_LOC_737/A 0.07fF
C13113 OR2X1_LOC_715/B OR2X1_LOC_687/Y 0.10fF
C13114 AND2X1_LOC_95/Y OR2X1_LOC_787/B 0.01fF
C13115 OR2X1_LOC_261/a_8_216# AND2X1_LOC_847/Y 0.01fF
C13116 OR2X1_LOC_346/B OR2X1_LOC_736/Y 0.01fF
C13117 OR2X1_LOC_185/A OR2X1_LOC_785/a_8_216# 0.01fF
C13118 OR2X1_LOC_377/A AND2X1_LOC_616/a_8_24# 0.03fF
C13119 AND2X1_LOC_70/Y OR2X1_LOC_541/B 0.08fF
C13120 AND2X1_LOC_511/a_8_24# OR2X1_LOC_269/B 0.01fF
C13121 AND2X1_LOC_59/Y OR2X1_LOC_66/A 1.00fF
C13122 AND2X1_LOC_658/A AND2X1_LOC_858/a_8_24# 0.04fF
C13123 AND2X1_LOC_658/A AND2X1_LOC_622/a_8_24# 0.01fF
C13124 AND2X1_LOC_95/Y AND2X1_LOC_92/Y 0.22fF
C13125 OR2X1_LOC_114/Y OR2X1_LOC_362/A 0.01fF
C13126 OR2X1_LOC_619/Y AND2X1_LOC_658/a_36_24# 0.00fF
C13127 AND2X1_LOC_61/Y OR2X1_LOC_316/Y 0.03fF
C13128 OR2X1_LOC_52/B OR2X1_LOC_421/Y 0.01fF
C13129 AND2X1_LOC_59/Y OR2X1_LOC_841/A 0.06fF
C13130 OR2X1_LOC_203/Y OR2X1_LOC_631/A 0.04fF
C13131 AND2X1_LOC_50/Y D_INPUT_5 1.38fF
C13132 OR2X1_LOC_831/a_8_216# VDD 0.21fF
C13133 AND2X1_LOC_570/Y AND2X1_LOC_577/Y 0.00fF
C13134 OR2X1_LOC_633/Y AND2X1_LOC_92/Y 0.23fF
C13135 AND2X1_LOC_734/a_8_24# OR2X1_LOC_527/Y 0.01fF
C13136 AND2X1_LOC_713/a_8_24# OR2X1_LOC_89/A 0.01fF
C13137 AND2X1_LOC_82/Y OR2X1_LOC_557/A 0.05fF
C13138 AND2X1_LOC_573/A AND2X1_LOC_663/A 0.05fF
C13139 OR2X1_LOC_629/a_36_216# OR2X1_LOC_161/B 0.00fF
C13140 AND2X1_LOC_847/Y OR2X1_LOC_297/A 0.01fF
C13141 VDD OR2X1_LOC_216/Y 0.34fF
C13142 AND2X1_LOC_207/A OR2X1_LOC_43/A 0.01fF
C13143 AND2X1_LOC_43/B OR2X1_LOC_78/A 0.23fF
C13144 OR2X1_LOC_188/Y AND2X1_LOC_75/a_36_24# 0.00fF
C13145 OR2X1_LOC_757/A AND2X1_LOC_624/A 0.03fF
C13146 OR2X1_LOC_7/A AND2X1_LOC_476/Y 1.28fF
C13147 AND2X1_LOC_121/a_36_24# OR2X1_LOC_67/A 0.00fF
C13148 OR2X1_LOC_648/B OR2X1_LOC_208/a_8_216# 0.33fF
C13149 OR2X1_LOC_744/A AND2X1_LOC_318/a_8_24# 0.06fF
C13150 AND2X1_LOC_663/B OR2X1_LOC_759/a_8_216# 0.01fF
C13151 AND2X1_LOC_500/Y AND2X1_LOC_576/Y 0.00fF
C13152 OR2X1_LOC_364/A OR2X1_LOC_648/A 0.02fF
C13153 VDD OR2X1_LOC_214/a_8_216# 0.00fF
C13154 OR2X1_LOC_185/Y OR2X1_LOC_648/A 0.07fF
C13155 OR2X1_LOC_305/Y OR2X1_LOC_426/B 0.00fF
C13156 AND2X1_LOC_533/a_36_24# OR2X1_LOC_538/A 0.00fF
C13157 OR2X1_LOC_762/a_8_216# OR2X1_LOC_12/Y 0.19fF
C13158 VDD AND2X1_LOC_853/Y 0.05fF
C13159 AND2X1_LOC_119/a_8_24# AND2X1_LOC_44/Y 0.00fF
C13160 AND2X1_LOC_392/A AND2X1_LOC_123/a_8_24# 0.03fF
C13161 OR2X1_LOC_9/Y OR2X1_LOC_824/a_8_216# 0.01fF
C13162 OR2X1_LOC_158/A AND2X1_LOC_473/a_8_24# 0.02fF
C13163 OR2X1_LOC_51/Y OR2X1_LOC_669/a_8_216# 0.01fF
C13164 OR2X1_LOC_43/A OR2X1_LOC_690/Y 0.01fF
C13165 OR2X1_LOC_458/B AND2X1_LOC_43/B 0.12fF
C13166 OR2X1_LOC_6/B AND2X1_LOC_85/a_36_24# 0.01fF
C13167 OR2X1_LOC_857/B AND2X1_LOC_689/a_8_24# 0.01fF
C13168 OR2X1_LOC_154/A OR2X1_LOC_678/Y 0.02fF
C13169 OR2X1_LOC_380/A OR2X1_LOC_26/a_36_216# 0.00fF
C13170 OR2X1_LOC_405/A OR2X1_LOC_475/a_36_216# -0.02fF
C13171 OR2X1_LOC_611/a_8_216# OR2X1_LOC_16/A 0.07fF
C13172 OR2X1_LOC_151/A OR2X1_LOC_486/B 0.02fF
C13173 VDD OR2X1_LOC_787/Y 0.35fF
C13174 OR2X1_LOC_744/A AND2X1_LOC_361/A 0.07fF
C13175 AND2X1_LOC_537/Y OR2X1_LOC_16/A 0.03fF
C13176 OR2X1_LOC_235/B OR2X1_LOC_643/A 0.03fF
C13177 AND2X1_LOC_76/Y AND2X1_LOC_662/B 0.02fF
C13178 AND2X1_LOC_367/A AND2X1_LOC_560/B 0.10fF
C13179 OR2X1_LOC_688/Y OR2X1_LOC_66/A 0.01fF
C13180 AND2X1_LOC_520/a_8_24# OR2X1_LOC_111/Y 0.02fF
C13181 VDD OR2X1_LOC_17/Y 0.05fF
C13182 OR2X1_LOC_201/A OR2X1_LOC_87/A 0.09fF
C13183 OR2X1_LOC_865/B OR2X1_LOC_571/B 0.02fF
C13184 OR2X1_LOC_448/Y OR2X1_LOC_712/a_36_216# 0.00fF
C13185 AND2X1_LOC_72/B OR2X1_LOC_500/a_8_216# 0.01fF
C13186 AND2X1_LOC_533/a_8_24# OR2X1_LOC_620/Y -0.03fF
C13187 AND2X1_LOC_851/a_8_24# OR2X1_LOC_238/Y 0.01fF
C13188 VDD OR2X1_LOC_282/Y 0.04fF
C13189 AND2X1_LOC_850/a_8_24# OR2X1_LOC_18/Y -0.01fF
C13190 D_INPUT_4 AND2X1_LOC_1/a_8_24# 0.02fF
C13191 AND2X1_LOC_723/Y AND2X1_LOC_784/A 0.54fF
C13192 AND2X1_LOC_675/A AND2X1_LOC_804/A 0.02fF
C13193 OR2X1_LOC_95/Y GATE_579 0.00fF
C13194 AND2X1_LOC_842/B AND2X1_LOC_500/B 0.53fF
C13195 AND2X1_LOC_716/Y OR2X1_LOC_6/A 0.09fF
C13196 OR2X1_LOC_538/a_8_216# OR2X1_LOC_269/B 0.01fF
C13197 OR2X1_LOC_67/A OR2X1_LOC_278/Y 0.00fF
C13198 OR2X1_LOC_600/A AND2X1_LOC_523/Y 0.03fF
C13199 OR2X1_LOC_306/Y OR2X1_LOC_48/B 0.00fF
C13200 OR2X1_LOC_760/a_8_216# OR2X1_LOC_312/a_8_216# 0.47fF
C13201 OR2X1_LOC_228/Y OR2X1_LOC_723/B 0.01fF
C13202 OR2X1_LOC_753/A OR2X1_LOC_16/a_8_216# 0.38fF
C13203 OR2X1_LOC_840/A OR2X1_LOC_449/B 0.79fF
C13204 INPUT_0 OR2X1_LOC_74/A 0.01fF
C13205 AND2X1_LOC_70/Y OR2X1_LOC_602/a_36_216# 0.00fF
C13206 AND2X1_LOC_207/a_8_24# OR2X1_LOC_3/Y 0.03fF
C13207 AND2X1_LOC_39/a_8_24# OR2X1_LOC_155/A 0.03fF
C13208 AND2X1_LOC_654/Y OR2X1_LOC_6/A 0.01fF
C13209 AND2X1_LOC_486/Y OR2X1_LOC_26/Y 0.06fF
C13210 OR2X1_LOC_502/A AND2X1_LOC_611/a_8_24# 0.01fF
C13211 OR2X1_LOC_91/A AND2X1_LOC_212/B 0.03fF
C13212 AND2X1_LOC_392/A OR2X1_LOC_268/a_8_216# 0.04fF
C13213 AND2X1_LOC_722/A OR2X1_LOC_485/A 0.08fF
C13214 OR2X1_LOC_8/Y OR2X1_LOC_19/B 0.06fF
C13215 AND2X1_LOC_505/a_8_24# OR2X1_LOC_814/A 0.04fF
C13216 OR2X1_LOC_389/A AND2X1_LOC_48/A 0.03fF
C13217 AND2X1_LOC_486/Y AND2X1_LOC_493/a_8_24# 0.08fF
C13218 OR2X1_LOC_600/A OR2X1_LOC_815/A 0.03fF
C13219 OR2X1_LOC_311/Y OR2X1_LOC_426/B 0.03fF
C13220 AND2X1_LOC_386/a_8_24# D_INPUT_4 0.01fF
C13221 OR2X1_LOC_154/A OR2X1_LOC_404/a_8_216# 0.08fF
C13222 OR2X1_LOC_91/A OR2X1_LOC_829/Y 0.10fF
C13223 AND2X1_LOC_779/a_36_24# OR2X1_LOC_44/Y 0.02fF
C13224 AND2X1_LOC_486/Y OR2X1_LOC_89/A 0.03fF
C13225 OR2X1_LOC_105/Y AND2X1_LOC_42/B 0.00fF
C13226 AND2X1_LOC_654/Y OR2X1_LOC_299/a_8_216# 0.03fF
C13227 OR2X1_LOC_494/a_8_216# OR2X1_LOC_481/A 0.47fF
C13228 VDD OR2X1_LOC_243/a_8_216# 0.21fF
C13229 OR2X1_LOC_116/A OR2X1_LOC_114/Y 0.06fF
C13230 OR2X1_LOC_6/B AND2X1_LOC_47/Y 0.09fF
C13231 AND2X1_LOC_651/a_8_24# AND2X1_LOC_651/B 0.00fF
C13232 AND2X1_LOC_662/B OR2X1_LOC_52/B 0.02fF
C13233 OR2X1_LOC_334/B AND2X1_LOC_51/Y 0.03fF
C13234 OR2X1_LOC_841/a_36_216# OR2X1_LOC_479/Y 0.01fF
C13235 AND2X1_LOC_717/Y OR2X1_LOC_74/A 0.02fF
C13236 OR2X1_LOC_680/A OR2X1_LOC_613/Y 0.00fF
C13237 AND2X1_LOC_367/A OR2X1_LOC_64/Y 0.05fF
C13238 OR2X1_LOC_250/Y OR2X1_LOC_585/A 0.15fF
C13239 AND2X1_LOC_465/Y OR2X1_LOC_59/Y 0.01fF
C13240 AND2X1_LOC_273/a_36_24# OR2X1_LOC_318/B 0.00fF
C13241 AND2X1_LOC_729/Y OR2X1_LOC_601/Y 0.13fF
C13242 OR2X1_LOC_316/Y AND2X1_LOC_852/Y 0.03fF
C13243 OR2X1_LOC_318/Y OR2X1_LOC_479/Y 0.01fF
C13244 OR2X1_LOC_464/A OR2X1_LOC_675/A 0.01fF
C13245 OR2X1_LOC_188/Y OR2X1_LOC_318/B 0.03fF
C13246 OR2X1_LOC_671/Y OR2X1_LOC_47/Y 0.07fF
C13247 AND2X1_LOC_544/Y AND2X1_LOC_222/Y 0.03fF
C13248 AND2X1_LOC_43/B OR2X1_LOC_155/A 0.04fF
C13249 OR2X1_LOC_814/A OR2X1_LOC_795/B 0.03fF
C13250 AND2X1_LOC_571/Y OR2X1_LOC_89/A 0.07fF
C13251 OR2X1_LOC_125/a_8_216# OR2X1_LOC_95/Y 0.10fF
C13252 OR2X1_LOC_400/A OR2X1_LOC_403/B 1.20fF
C13253 OR2X1_LOC_106/a_8_216# OR2X1_LOC_47/Y 0.07fF
C13254 D_INPUT_0 OR2X1_LOC_715/A 0.06fF
C13255 OR2X1_LOC_382/Y OR2X1_LOC_54/Y 0.01fF
C13256 OR2X1_LOC_840/A OR2X1_LOC_121/B 0.01fF
C13257 OR2X1_LOC_26/Y AND2X1_LOC_834/a_8_24# 0.02fF
C13258 AND2X1_LOC_76/Y OR2X1_LOC_273/Y 0.02fF
C13259 OR2X1_LOC_715/B OR2X1_LOC_786/Y 0.03fF
C13260 OR2X1_LOC_235/B OR2X1_LOC_113/A 0.00fF
C13261 OR2X1_LOC_156/Y OR2X1_LOC_160/a_8_216# 0.38fF
C13262 OR2X1_LOC_421/A AND2X1_LOC_648/B 1.51fF
C13263 AND2X1_LOC_767/a_36_24# AND2X1_LOC_3/Y 0.00fF
C13264 AND2X1_LOC_456/Y OR2X1_LOC_503/A 0.15fF
C13265 OR2X1_LOC_127/Y AND2X1_LOC_554/B 0.79fF
C13266 OR2X1_LOC_699/a_36_216# OR2X1_LOC_820/B 0.00fF
C13267 AND2X1_LOC_70/Y OR2X1_LOC_440/A 0.08fF
C13268 OR2X1_LOC_36/Y OR2X1_LOC_585/A 0.16fF
C13269 OR2X1_LOC_26/Y OR2X1_LOC_248/Y 0.18fF
C13270 OR2X1_LOC_426/B D_INPUT_3 0.07fF
C13271 OR2X1_LOC_435/a_36_216# OR2X1_LOC_814/A 0.01fF
C13272 OR2X1_LOC_26/Y OR2X1_LOC_6/a_8_216# 0.01fF
C13273 AND2X1_LOC_559/a_36_24# OR2X1_LOC_52/B 0.01fF
C13274 AND2X1_LOC_7/B OR2X1_LOC_68/B 0.29fF
C13275 OR2X1_LOC_604/A AND2X1_LOC_620/Y 0.07fF
C13276 AND2X1_LOC_56/B OR2X1_LOC_296/a_8_216# 0.07fF
C13277 OR2X1_LOC_87/A AND2X1_LOC_3/Y 0.26fF
C13278 OR2X1_LOC_160/B OR2X1_LOC_779/Y 0.03fF
C13279 AND2X1_LOC_367/A OR2X1_LOC_417/A 0.12fF
C13280 OR2X1_LOC_87/A OR2X1_LOC_647/B 0.39fF
C13281 OR2X1_LOC_614/Y OR2X1_LOC_196/a_8_216# 0.01fF
C13282 OR2X1_LOC_653/Y OR2X1_LOC_750/A 0.00fF
C13283 AND2X1_LOC_40/Y OR2X1_LOC_814/A 2.78fF
C13284 OR2X1_LOC_816/A AND2X1_LOC_657/A 0.07fF
C13285 VDD OR2X1_LOC_588/A 0.09fF
C13286 OR2X1_LOC_599/A OR2X1_LOC_485/A 0.04fF
C13287 AND2X1_LOC_59/Y AND2X1_LOC_176/a_36_24# 0.00fF
C13288 AND2X1_LOC_12/Y OR2X1_LOC_473/Y 0.05fF
C13289 AND2X1_LOC_605/Y OR2X1_LOC_31/Y 0.76fF
C13290 AND2X1_LOC_349/B OR2X1_LOC_248/Y 0.28fF
C13291 OR2X1_LOC_753/A OR2X1_LOC_24/Y 0.05fF
C13292 OR2X1_LOC_305/Y OR2X1_LOC_743/A 0.03fF
C13293 OR2X1_LOC_329/B OR2X1_LOC_760/a_36_216# 0.02fF
C13294 AND2X1_LOC_560/B OR2X1_LOC_74/A 0.14fF
C13295 AND2X1_LOC_36/Y OR2X1_LOC_703/Y 0.04fF
C13296 VDD OR2X1_LOC_396/Y 0.00fF
C13297 OR2X1_LOC_844/a_8_216# OR2X1_LOC_643/A 0.01fF
C13298 AND2X1_LOC_43/a_36_24# OR2X1_LOC_269/B 0.01fF
C13299 OR2X1_LOC_97/A OR2X1_LOC_365/a_8_216# 0.01fF
C13300 OR2X1_LOC_6/B OR2X1_LOC_598/A 0.26fF
C13301 OR2X1_LOC_473/a_36_216# OR2X1_LOC_532/B 0.00fF
C13302 OR2X1_LOC_111/Y OR2X1_LOC_92/Y 0.00fF
C13303 OR2X1_LOC_11/Y OR2X1_LOC_762/a_36_216# 0.00fF
C13304 AND2X1_LOC_70/Y OR2X1_LOC_446/A 0.01fF
C13305 OR2X1_LOC_643/Y OR2X1_LOC_215/Y 0.09fF
C13306 AND2X1_LOC_102/a_8_24# AND2X1_LOC_42/B 0.17fF
C13307 AND2X1_LOC_227/Y OR2X1_LOC_265/a_36_216# 0.00fF
C13308 OR2X1_LOC_499/a_8_216# OR2X1_LOC_62/B 0.01fF
C13309 OR2X1_LOC_273/Y OR2X1_LOC_52/B 0.02fF
C13310 OR2X1_LOC_261/Y AND2X1_LOC_345/a_8_24# 0.00fF
C13311 AND2X1_LOC_47/Y OR2X1_LOC_523/Y 0.03fF
C13312 OR2X1_LOC_849/A OR2X1_LOC_404/Y 2.15fF
C13313 AND2X1_LOC_3/Y AND2X1_LOC_815/a_8_24# 0.07fF
C13314 OR2X1_LOC_118/Y AND2X1_LOC_845/Y 0.01fF
C13315 OR2X1_LOC_676/a_8_216# OR2X1_LOC_228/Y 0.06fF
C13316 INPUT_4 AND2X1_LOC_635/a_36_24# -0.00fF
C13317 OR2X1_LOC_228/a_8_216# AND2X1_LOC_43/B 0.03fF
C13318 AND2X1_LOC_76/Y OR2X1_LOC_75/Y 0.04fF
C13319 OR2X1_LOC_305/Y OR2X1_LOC_246/A 0.02fF
C13320 AND2X1_LOC_456/Y OR2X1_LOC_64/Y 0.02fF
C13321 OR2X1_LOC_64/Y OR2X1_LOC_74/A 0.12fF
C13322 OR2X1_LOC_417/Y OR2X1_LOC_743/A 0.03fF
C13323 OR2X1_LOC_648/A AND2X1_LOC_432/a_8_24# 0.03fF
C13324 OR2X1_LOC_827/Y OR2X1_LOC_46/A 0.01fF
C13325 OR2X1_LOC_809/a_8_216# OR2X1_LOC_532/B 0.02fF
C13326 OR2X1_LOC_222/a_8_216# OR2X1_LOC_130/A 0.30fF
C13327 OR2X1_LOC_311/Y OR2X1_LOC_743/A 0.03fF
C13328 OR2X1_LOC_834/A OR2X1_LOC_513/a_8_216# 0.01fF
C13329 OR2X1_LOC_231/A OR2X1_LOC_205/Y 0.00fF
C13330 OR2X1_LOC_49/A AND2X1_LOC_36/Y 0.17fF
C13331 OR2X1_LOC_864/A OR2X1_LOC_532/B 0.03fF
C13332 INPUT_3 AND2X1_LOC_8/a_8_24# 0.02fF
C13333 AND2X1_LOC_538/Y OR2X1_LOC_743/A 0.01fF
C13334 OR2X1_LOC_70/Y OR2X1_LOC_245/a_8_216# 0.01fF
C13335 OR2X1_LOC_532/B OR2X1_LOC_240/A 0.02fF
C13336 AND2X1_LOC_639/B OR2X1_LOC_387/A 0.01fF
C13337 OR2X1_LOC_369/a_8_216# OR2X1_LOC_437/A 0.03fF
C13338 OR2X1_LOC_186/Y OR2X1_LOC_308/Y 0.15fF
C13339 OR2X1_LOC_100/Y OR2X1_LOC_608/Y 0.27fF
C13340 OR2X1_LOC_64/Y OR2X1_LOC_762/a_36_216# 0.00fF
C13341 OR2X1_LOC_633/B OR2X1_LOC_532/B 0.04fF
C13342 AND2X1_LOC_12/Y OR2X1_LOC_214/B 0.03fF
C13343 OR2X1_LOC_161/A AND2X1_LOC_418/a_8_24# 0.01fF
C13344 AND2X1_LOC_387/B D_INPUT_0 2.06fF
C13345 OR2X1_LOC_119/a_8_216# OR2X1_LOC_278/A 0.03fF
C13346 OR2X1_LOC_36/Y AND2X1_LOC_645/a_8_24# 0.01fF
C13347 AND2X1_LOC_460/a_8_24# OR2X1_LOC_11/Y 0.01fF
C13348 AND2X1_LOC_216/A OR2X1_LOC_278/Y 0.02fF
C13349 OR2X1_LOC_616/Y AND2X1_LOC_792/Y 0.00fF
C13350 OR2X1_LOC_596/A AND2X1_LOC_36/Y 0.08fF
C13351 OR2X1_LOC_160/A OR2X1_LOC_804/A 0.13fF
C13352 AND2X1_LOC_796/a_8_24# OR2X1_LOC_142/Y 0.24fF
C13353 AND2X1_LOC_753/B OR2X1_LOC_197/a_8_216# 0.03fF
C13354 OR2X1_LOC_599/A AND2X1_LOC_645/a_36_24# 0.00fF
C13355 OR2X1_LOC_75/Y OR2X1_LOC_52/B 0.00fF
C13356 OR2X1_LOC_391/a_8_216# OR2X1_LOC_561/B 0.02fF
C13357 OR2X1_LOC_74/A OR2X1_LOC_417/A 0.75fF
C13358 OR2X1_LOC_130/A OR2X1_LOC_205/Y 0.00fF
C13359 OR2X1_LOC_234/a_8_216# OR2X1_LOC_85/A 0.01fF
C13360 OR2X1_LOC_779/Y OR2X1_LOC_779/a_36_216# 0.01fF
C13361 AND2X1_LOC_85/a_36_24# AND2X1_LOC_47/Y 0.00fF
C13362 OR2X1_LOC_726/A OR2X1_LOC_308/Y 0.01fF
C13363 AND2X1_LOC_10/a_8_24# OR2X1_LOC_244/A 0.02fF
C13364 OR2X1_LOC_485/A AND2X1_LOC_866/A 0.04fF
C13365 OR2X1_LOC_532/B AND2X1_LOC_281/a_8_24# 0.01fF
C13366 OR2X1_LOC_131/Y OR2X1_LOC_95/Y 0.03fF
C13367 AND2X1_LOC_11/Y AND2X1_LOC_429/a_8_24# 0.03fF
C13368 OR2X1_LOC_553/A AND2X1_LOC_237/a_36_24# 0.00fF
C13369 OR2X1_LOC_66/A OR2X1_LOC_342/B 0.01fF
C13370 AND2X1_LOC_245/a_8_24# OR2X1_LOC_777/B 0.00fF
C13371 AND2X1_LOC_81/a_8_24# OR2X1_LOC_786/Y 0.24fF
C13372 AND2X1_LOC_550/A AND2X1_LOC_222/Y 0.03fF
C13373 AND2X1_LOC_92/Y OR2X1_LOC_788/B 0.03fF
C13374 OR2X1_LOC_12/Y AND2X1_LOC_773/a_8_24# 0.04fF
C13375 AND2X1_LOC_48/A OR2X1_LOC_649/a_8_216# 0.01fF
C13376 AND2X1_LOC_593/a_8_24# OR2X1_LOC_696/A 0.04fF
C13377 OR2X1_LOC_169/a_8_216# OR2X1_LOC_365/B 0.00fF
C13378 OR2X1_LOC_468/Y OR2X1_LOC_365/B 0.02fF
C13379 AND2X1_LOC_839/A OR2X1_LOC_54/Y 0.05fF
C13380 AND2X1_LOC_807/Y AND2X1_LOC_657/A 0.10fF
C13381 OR2X1_LOC_377/A OR2X1_LOC_378/A 0.32fF
C13382 OR2X1_LOC_241/Y OR2X1_LOC_121/B 0.02fF
C13383 OR2X1_LOC_805/A OR2X1_LOC_68/B 0.07fF
C13384 AND2X1_LOC_773/Y OR2X1_LOC_12/Y 0.17fF
C13385 AND2X1_LOC_826/a_36_24# OR2X1_LOC_46/A 0.00fF
C13386 AND2X1_LOC_399/a_8_24# OR2X1_LOC_398/Y 0.09fF
C13387 AND2X1_LOC_719/Y AND2X1_LOC_241/a_36_24# 0.06fF
C13388 AND2X1_LOC_153/a_36_24# OR2X1_LOC_68/B 0.00fF
C13389 AND2X1_LOC_576/Y AND2X1_LOC_563/Y 0.01fF
C13390 D_INPUT_3 OR2X1_LOC_125/Y 0.01fF
C13391 OR2X1_LOC_744/A OR2X1_LOC_387/A 0.18fF
C13392 OR2X1_LOC_574/A AND2X1_LOC_679/a_8_24# 0.20fF
C13393 INPUT_0 AND2X1_LOC_235/a_8_24# 0.02fF
C13394 OR2X1_LOC_188/Y OR2X1_LOC_190/a_8_216# 0.18fF
C13395 AND2X1_LOC_626/a_36_24# AND2X1_LOC_7/B 0.01fF
C13396 OR2X1_LOC_620/Y OR2X1_LOC_777/B 0.07fF
C13397 OR2X1_LOC_778/Y OR2X1_LOC_779/B 0.17fF
C13398 AND2X1_LOC_51/Y AND2X1_LOC_418/a_8_24# 0.02fF
C13399 OR2X1_LOC_607/a_8_216# OR2X1_LOC_607/Y -0.00fF
C13400 OR2X1_LOC_53/Y AND2X1_LOC_200/a_36_24# 0.00fF
C13401 OR2X1_LOC_40/Y OR2X1_LOC_764/a_36_216# 0.03fF
C13402 VDD AND2X1_LOC_473/Y 0.21fF
C13403 VDD AND2X1_LOC_287/B 0.29fF
C13404 D_INPUT_3 OR2X1_LOC_225/a_8_216# 0.01fF
C13405 OR2X1_LOC_133/a_8_216# OR2X1_LOC_158/A 0.02fF
C13406 OR2X1_LOC_406/Y AND2X1_LOC_658/B 0.03fF
C13407 AND2X1_LOC_47/Y D_GATE_222 0.09fF
C13408 AND2X1_LOC_477/A OR2X1_LOC_47/Y 0.42fF
C13409 AND2X1_LOC_43/B OR2X1_LOC_515/a_36_216# 0.00fF
C13410 VDD OR2X1_LOC_816/A 0.32fF
C13411 AND2X1_LOC_166/a_8_24# OR2X1_LOC_788/B 0.02fF
C13412 OR2X1_LOC_379/Y OR2X1_LOC_771/B 0.01fF
C13413 VDD OR2X1_LOC_576/A 0.19fF
C13414 OR2X1_LOC_12/Y AND2X1_LOC_243/Y 0.07fF
C13415 VDD OR2X1_LOC_79/Y 0.06fF
C13416 AND2X1_LOC_91/B OR2X1_LOC_235/B 0.01fF
C13417 AND2X1_LOC_64/Y AND2X1_LOC_71/a_8_24# 0.01fF
C13418 AND2X1_LOC_349/a_8_24# OR2X1_LOC_437/A 0.01fF
C13419 OR2X1_LOC_64/Y AND2X1_LOC_647/Y 0.03fF
C13420 OR2X1_LOC_732/a_8_216# AND2X1_LOC_36/Y 0.01fF
C13421 OR2X1_LOC_161/A OR2X1_LOC_523/A 0.01fF
C13422 AND2X1_LOC_22/Y AND2X1_LOC_92/Y 0.17fF
C13423 OR2X1_LOC_154/A OR2X1_LOC_777/B 0.10fF
C13424 OR2X1_LOC_6/A OR2X1_LOC_13/B 0.03fF
C13425 OR2X1_LOC_51/Y AND2X1_LOC_786/Y 0.03fF
C13426 OR2X1_LOC_19/B AND2X1_LOC_216/A 0.02fF
C13427 AND2X1_LOC_729/Y OR2X1_LOC_142/Y 0.02fF
C13428 OR2X1_LOC_562/a_8_216# OR2X1_LOC_562/B 0.39fF
C13429 AND2X1_LOC_48/A OR2X1_LOC_801/B 0.39fF
C13430 AND2X1_LOC_811/Y AND2X1_LOC_812/a_8_24# 0.06fF
C13431 OR2X1_LOC_597/A AND2X1_LOC_771/B 0.01fF
C13432 AND2X1_LOC_725/a_8_24# OR2X1_LOC_158/A 0.01fF
C13433 OR2X1_LOC_40/Y AND2X1_LOC_182/a_8_24# 0.02fF
C13434 VDD OR2X1_LOC_439/B 0.23fF
C13435 OR2X1_LOC_488/Y AND2X1_LOC_657/A 0.00fF
C13436 AND2X1_LOC_857/Y OR2X1_LOC_321/a_36_216# 0.00fF
C13437 AND2X1_LOC_42/B OR2X1_LOC_71/A 1.29fF
C13438 AND2X1_LOC_810/A INPUT_0 0.03fF
C13439 OR2X1_LOC_502/A OR2X1_LOC_390/a_36_216# -0.02fF
C13440 AND2X1_LOC_570/Y OR2X1_LOC_482/Y 0.03fF
C13441 AND2X1_LOC_463/B OR2X1_LOC_409/a_8_216# 0.01fF
C13442 OR2X1_LOC_701/a_8_216# AND2X1_LOC_789/Y 0.02fF
C13443 OR2X1_LOC_87/B AND2X1_LOC_36/Y 5.54fF
C13444 OR2X1_LOC_703/B OR2X1_LOC_388/a_8_216# 0.18fF
C13445 OR2X1_LOC_95/Y AND2X1_LOC_644/a_8_24# 0.01fF
C13446 AND2X1_LOC_778/a_8_24# OR2X1_LOC_142/Y 0.02fF
C13447 OR2X1_LOC_589/A OR2X1_LOC_597/a_8_216# 0.11fF
C13448 AND2X1_LOC_47/Y OR2X1_LOC_598/A 0.14fF
C13449 OR2X1_LOC_51/Y AND2X1_LOC_499/a_36_24# 0.00fF
C13450 OR2X1_LOC_542/B OR2X1_LOC_741/Y 0.03fF
C13451 AND2X1_LOC_191/B OR2X1_LOC_600/A 0.03fF
C13452 OR2X1_LOC_158/A OR2X1_LOC_292/Y 0.00fF
C13453 OR2X1_LOC_600/A AND2X1_LOC_469/B 0.00fF
C13454 OR2X1_LOC_188/Y AND2X1_LOC_12/Y 0.01fF
C13455 OR2X1_LOC_154/A OR2X1_LOC_831/B 0.32fF
C13456 OR2X1_LOC_325/B OR2X1_LOC_538/A 0.04fF
C13457 AND2X1_LOC_624/B AND2X1_LOC_792/Y 0.02fF
C13458 AND2X1_LOC_642/a_8_24# AND2X1_LOC_786/Y 0.06fF
C13459 OR2X1_LOC_188/a_8_216# OR2X1_LOC_154/A 0.05fF
C13460 AND2X1_LOC_571/a_8_24# AND2X1_LOC_572/Y 0.01fF
C13461 OR2X1_LOC_78/Y AND2X1_LOC_18/Y 0.01fF
C13462 OR2X1_LOC_696/A OR2X1_LOC_106/A 0.03fF
C13463 OR2X1_LOC_36/Y AND2X1_LOC_455/a_8_24# 0.14fF
C13464 OR2X1_LOC_323/A AND2X1_LOC_374/Y 0.02fF
C13465 OR2X1_LOC_95/Y AND2X1_LOC_657/A 0.08fF
C13466 OR2X1_LOC_274/a_8_216# AND2X1_LOC_18/Y 0.18fF
C13467 OR2X1_LOC_241/a_8_216# AND2X1_LOC_7/B 0.03fF
C13468 OR2X1_LOC_349/a_8_216# OR2X1_LOC_850/a_8_216# 0.47fF
C13469 OR2X1_LOC_48/B AND2X1_LOC_212/Y 0.07fF
C13470 VDD AND2X1_LOC_41/A 1.00fF
C13471 AND2X1_LOC_509/Y AND2X1_LOC_658/A 0.03fF
C13472 OR2X1_LOC_240/a_8_216# OR2X1_LOC_633/A 0.03fF
C13473 OR2X1_LOC_85/A AND2X1_LOC_202/Y 0.01fF
C13474 AND2X1_LOC_784/A OR2X1_LOC_136/a_8_216# 0.13fF
C13475 OR2X1_LOC_40/Y AND2X1_LOC_168/a_8_24# 0.02fF
C13476 VDD OR2X1_LOC_251/a_8_216# 0.21fF
C13477 OR2X1_LOC_516/Y OR2X1_LOC_70/Y 0.03fF
C13478 OR2X1_LOC_560/a_36_216# OR2X1_LOC_113/B 0.00fF
C13479 OR2X1_LOC_680/A AND2X1_LOC_786/Y 0.07fF
C13480 AND2X1_LOC_164/a_8_24# OR2X1_LOC_168/B 0.01fF
C13481 OR2X1_LOC_40/Y AND2X1_LOC_851/A 0.01fF
C13482 AND2X1_LOC_775/a_36_24# OR2X1_LOC_70/Y 0.01fF
C13483 AND2X1_LOC_706/Y OR2X1_LOC_424/a_8_216# 0.03fF
C13484 OR2X1_LOC_743/A AND2X1_LOC_780/a_8_24# 0.01fF
C13485 AND2X1_LOC_548/Y AND2X1_LOC_549/a_36_24# 0.01fF
C13486 AND2X1_LOC_842/a_8_24# OR2X1_LOC_59/Y 0.02fF
C13487 OR2X1_LOC_638/B OR2X1_LOC_638/a_8_216# 0.05fF
C13488 AND2X1_LOC_70/Y OR2X1_LOC_637/A 0.01fF
C13489 AND2X1_LOC_717/B AND2X1_LOC_465/A 0.21fF
C13490 OR2X1_LOC_753/A AND2X1_LOC_208/Y 0.54fF
C13491 OR2X1_LOC_251/Y AND2X1_LOC_287/B 0.08fF
C13492 OR2X1_LOC_459/A INPUT_0 0.34fF
C13493 OR2X1_LOC_447/a_36_216# OR2X1_LOC_596/A 0.02fF
C13494 AND2X1_LOC_79/a_8_24# AND2X1_LOC_36/Y 0.14fF
C13495 OR2X1_LOC_264/Y AND2X1_LOC_70/Y 0.09fF
C13496 OR2X1_LOC_865/A OR2X1_LOC_774/Y 0.06fF
C13497 OR2X1_LOC_717/a_8_216# OR2X1_LOC_723/A -0.00fF
C13498 OR2X1_LOC_744/a_8_216# OR2X1_LOC_52/B 0.03fF
C13499 OR2X1_LOC_148/Y OR2X1_LOC_213/A 0.28fF
C13500 AND2X1_LOC_544/Y OR2X1_LOC_74/A 0.03fF
C13501 AND2X1_LOC_724/A OR2X1_LOC_44/Y 0.08fF
C13502 OR2X1_LOC_272/Y AND2X1_LOC_773/a_8_24# 0.01fF
C13503 OR2X1_LOC_45/Y VDD 0.26fF
C13504 AND2X1_LOC_506/a_8_24# AND2X1_LOC_508/A 0.01fF
C13505 OR2X1_LOC_446/Y OR2X1_LOC_712/B 0.01fF
C13506 OR2X1_LOC_502/A AND2X1_LOC_144/a_8_24# 0.07fF
C13507 OR2X1_LOC_269/B OR2X1_LOC_725/A 0.01fF
C13508 AND2X1_LOC_772/B OR2X1_LOC_427/A 0.09fF
C13509 AND2X1_LOC_12/Y OR2X1_LOC_686/B 0.94fF
C13510 AND2X1_LOC_170/a_8_24# AND2X1_LOC_568/B 0.02fF
C13511 AND2X1_LOC_797/A AND2X1_LOC_220/B 0.45fF
C13512 OR2X1_LOC_223/A OR2X1_LOC_181/a_8_216# 0.01fF
C13513 OR2X1_LOC_629/a_8_216# OR2X1_LOC_563/A 0.02fF
C13514 OR2X1_LOC_676/Y OR2X1_LOC_161/A 0.07fF
C13515 OR2X1_LOC_335/A OR2X1_LOC_76/A 0.03fF
C13516 AND2X1_LOC_716/Y AND2X1_LOC_514/a_36_24# 0.01fF
C13517 OR2X1_LOC_610/a_8_216# OR2X1_LOC_78/A 0.03fF
C13518 OR2X1_LOC_709/A OR2X1_LOC_778/Y 0.10fF
C13519 OR2X1_LOC_662/A VDD 0.09fF
C13520 AND2X1_LOC_566/B AND2X1_LOC_354/B 0.04fF
C13521 OR2X1_LOC_696/A OR2X1_LOC_46/A 0.03fF
C13522 OR2X1_LOC_40/Y AND2X1_LOC_303/A 0.31fF
C13523 OR2X1_LOC_680/A AND2X1_LOC_499/a_36_24# 0.01fF
C13524 VDD AND2X1_LOC_807/Y 1.36fF
C13525 OR2X1_LOC_629/Y OR2X1_LOC_630/B 0.07fF
C13526 AND2X1_LOC_252/a_8_24# OR2X1_LOC_549/A 0.01fF
C13527 AND2X1_LOC_710/a_8_24# VDD -0.00fF
C13528 AND2X1_LOC_520/Y AND2X1_LOC_219/Y 0.12fF
C13529 AND2X1_LOC_12/Y OR2X1_LOC_862/B 0.25fF
C13530 OR2X1_LOC_70/Y OR2X1_LOC_373/a_8_216# 0.01fF
C13531 AND2X1_LOC_706/Y OR2X1_LOC_7/A 0.07fF
C13532 OR2X1_LOC_634/A AND2X1_LOC_690/a_8_24# 0.11fF
C13533 AND2X1_LOC_773/Y OR2X1_LOC_272/Y 0.01fF
C13534 AND2X1_LOC_120/a_8_24# AND2X1_LOC_244/A 0.00fF
C13535 OR2X1_LOC_834/A OR2X1_LOC_161/A 0.00fF
C13536 AND2X1_LOC_535/Y AND2X1_LOC_661/A 0.02fF
C13537 AND2X1_LOC_50/Y AND2X1_LOC_752/a_8_24# 0.04fF
C13538 OR2X1_LOC_160/B OR2X1_LOC_673/Y 0.03fF
C13539 AND2X1_LOC_182/A AND2X1_LOC_211/B 0.11fF
C13540 AND2X1_LOC_572/Y OR2X1_LOC_744/A 0.00fF
C13541 OR2X1_LOC_404/Y OR2X1_LOC_721/a_8_216# 0.01fF
C13542 AND2X1_LOC_512/Y AND2X1_LOC_801/a_8_24# 0.01fF
C13543 AND2X1_LOC_675/Y AND2X1_LOC_573/A 0.02fF
C13544 AND2X1_LOC_153/a_8_24# AND2X1_LOC_92/Y 0.06fF
C13545 OR2X1_LOC_3/Y AND2X1_LOC_339/B 0.03fF
C13546 OR2X1_LOC_31/Y OR2X1_LOC_387/A 0.01fF
C13547 AND2X1_LOC_40/Y OR2X1_LOC_147/B 0.06fF
C13548 OR2X1_LOC_702/A OR2X1_LOC_514/a_8_216# 0.01fF
C13549 OR2X1_LOC_510/Y OR2X1_LOC_78/A 0.10fF
C13550 OR2X1_LOC_468/A OR2X1_LOC_468/Y 0.02fF
C13551 VDD OR2X1_LOC_824/Y 0.00fF
C13552 AND2X1_LOC_56/B OR2X1_LOC_741/Y 0.05fF
C13553 VDD OR2X1_LOC_631/B 0.63fF
C13554 OR2X1_LOC_40/Y OR2X1_LOC_665/Y 0.01fF
C13555 OR2X1_LOC_40/Y AND2X1_LOC_474/Y 0.02fF
C13556 OR2X1_LOC_808/B OR2X1_LOC_211/a_8_216# 0.35fF
C13557 OR2X1_LOC_696/A AND2X1_LOC_227/Y 2.18fF
C13558 OR2X1_LOC_160/A AND2X1_LOC_65/a_8_24# 0.01fF
C13559 OR2X1_LOC_585/A AND2X1_LOC_207/B 0.18fF
C13560 OR2X1_LOC_476/B AND2X1_LOC_44/Y 0.07fF
C13561 OR2X1_LOC_666/A OR2X1_LOC_44/Y 0.05fF
C13562 AND2X1_LOC_47/Y OR2X1_LOC_186/a_8_216# 0.05fF
C13563 AND2X1_LOC_70/Y OR2X1_LOC_643/A 0.03fF
C13564 AND2X1_LOC_810/A OR2X1_LOC_64/Y 0.04fF
C13565 OR2X1_LOC_666/A AND2X1_LOC_288/a_8_24# 0.01fF
C13566 OR2X1_LOC_756/B OR2X1_LOC_570/a_8_216# 0.06fF
C13567 OR2X1_LOC_40/Y OR2X1_LOC_485/A 0.88fF
C13568 AND2X1_LOC_351/a_8_24# AND2X1_LOC_351/Y 0.01fF
C13569 OR2X1_LOC_757/A OR2X1_LOC_613/Y 0.00fF
C13570 AND2X1_LOC_70/Y OR2X1_LOC_124/Y 0.01fF
C13571 OR2X1_LOC_379/Y OR2X1_LOC_637/B 0.01fF
C13572 AND2X1_LOC_70/Y OR2X1_LOC_778/Y 0.03fF
C13573 VDD OR2X1_LOC_688/a_8_216# 0.21fF
C13574 OR2X1_LOC_347/a_36_216# OR2X1_LOC_811/A 0.17fF
C13575 OR2X1_LOC_647/Y AND2X1_LOC_607/a_8_24# 0.13fF
C13576 OR2X1_LOC_40/Y AND2X1_LOC_348/a_8_24# 0.01fF
C13577 AND2X1_LOC_50/Y AND2X1_LOC_59/Y 0.01fF
C13578 OR2X1_LOC_744/A AND2X1_LOC_852/Y 0.03fF
C13579 AND2X1_LOC_215/Y AND2X1_LOC_640/Y 0.01fF
C13580 OR2X1_LOC_810/A OR2X1_LOC_78/A 0.12fF
C13581 OR2X1_LOC_307/a_8_216# OR2X1_LOC_78/A 0.01fF
C13582 OR2X1_LOC_762/Y OR2X1_LOC_44/Y 0.04fF
C13583 OR2X1_LOC_83/Y OR2X1_LOC_744/A 0.01fF
C13584 AND2X1_LOC_711/Y AND2X1_LOC_507/a_8_24# 0.05fF
C13585 AND2X1_LOC_209/a_8_24# AND2X1_LOC_797/A 0.03fF
C13586 AND2X1_LOC_866/A AND2X1_LOC_455/a_36_24# 0.01fF
C13587 AND2X1_LOC_711/A OR2X1_LOC_258/Y 0.01fF
C13588 AND2X1_LOC_91/B OR2X1_LOC_276/B 0.10fF
C13589 AND2X1_LOC_36/Y AND2X1_LOC_761/a_36_24# 0.00fF
C13590 OR2X1_LOC_160/A OR2X1_LOC_231/A 0.03fF
C13591 AND2X1_LOC_794/B AND2X1_LOC_727/A 0.03fF
C13592 AND2X1_LOC_857/Y OR2X1_LOC_36/Y 0.04fF
C13593 OR2X1_LOC_3/Y OR2X1_LOC_816/a_8_216# 0.03fF
C13594 OR2X1_LOC_358/A OR2X1_LOC_539/B 0.02fF
C13595 OR2X1_LOC_703/A OR2X1_LOC_778/Y 0.14fF
C13596 OR2X1_LOC_154/A OR2X1_LOC_575/A 0.01fF
C13597 VDD AND2X1_LOC_135/a_8_24# 0.00fF
C13598 OR2X1_LOC_443/a_8_216# OR2X1_LOC_161/B 0.01fF
C13599 AND2X1_LOC_47/Y AND2X1_LOC_263/a_36_24# 0.00fF
C13600 AND2X1_LOC_589/a_8_24# OR2X1_LOC_78/A 0.02fF
C13601 AND2X1_LOC_862/a_8_24# AND2X1_LOC_862/Y 0.01fF
C13602 OR2X1_LOC_774/Y OR2X1_LOC_391/A 0.10fF
C13603 AND2X1_LOC_371/a_8_24# AND2X1_LOC_491/a_8_24# 0.23fF
C13604 VDD OR2X1_LOC_488/Y 0.08fF
C13605 OR2X1_LOC_121/Y D_INPUT_0 0.01fF
C13606 OR2X1_LOC_858/A AND2X1_LOC_42/B 3.92fF
C13607 OR2X1_LOC_64/Y AND2X1_LOC_860/A 0.02fF
C13608 OR2X1_LOC_676/Y AND2X1_LOC_51/Y 0.46fF
C13609 AND2X1_LOC_716/Y OR2X1_LOC_44/Y 0.07fF
C13610 OR2X1_LOC_80/a_8_216# OR2X1_LOC_16/A 0.07fF
C13611 OR2X1_LOC_849/A OR2X1_LOC_474/Y 0.17fF
C13612 D_INPUT_4 AND2X1_LOC_17/a_8_24# 0.02fF
C13613 OR2X1_LOC_251/Y OR2X1_LOC_251/a_8_216# 0.08fF
C13614 AND2X1_LOC_571/Y AND2X1_LOC_576/a_8_24# 0.18fF
C13615 AND2X1_LOC_317/a_36_24# OR2X1_LOC_427/A 0.00fF
C13616 OR2X1_LOC_278/Y AND2X1_LOC_286/Y 0.01fF
C13617 OR2X1_LOC_382/Y OR2X1_LOC_89/A 0.01fF
C13618 OR2X1_LOC_18/Y OR2X1_LOC_265/Y 0.00fF
C13619 AND2X1_LOC_858/B OR2X1_LOC_279/Y 0.03fF
C13620 AND2X1_LOC_215/Y OR2X1_LOC_416/Y 0.02fF
C13621 OR2X1_LOC_756/B OR2X1_LOC_557/A 0.06fF
C13622 OR2X1_LOC_351/B D_INPUT_0 0.39fF
C13623 AND2X1_LOC_40/Y OR2X1_LOC_383/a_8_216# 0.01fF
C13624 VDD AND2X1_LOC_727/A 0.60fF
C13625 OR2X1_LOC_160/A OR2X1_LOC_130/A 9.11fF
C13626 OR2X1_LOC_834/A AND2X1_LOC_51/Y 0.03fF
C13627 AND2X1_LOC_542/a_8_24# OR2X1_LOC_31/Y 0.01fF
C13628 AND2X1_LOC_40/Y AND2X1_LOC_171/a_8_24# 0.14fF
C13629 AND2X1_LOC_557/Y AND2X1_LOC_573/A 0.03fF
C13630 VDD OR2X1_LOC_403/a_8_216# 0.00fF
C13631 AND2X1_LOC_856/B AND2X1_LOC_434/Y 0.01fF
C13632 AND2X1_LOC_703/Y OR2X1_LOC_47/Y 0.03fF
C13633 AND2X1_LOC_566/B AND2X1_LOC_863/Y 0.09fF
C13634 AND2X1_LOC_794/B OR2X1_LOC_95/Y 0.07fF
C13635 OR2X1_LOC_247/a_8_216# AND2X1_LOC_7/B 0.07fF
C13636 AND2X1_LOC_40/Y AND2X1_LOC_387/B 0.27fF
C13637 OR2X1_LOC_6/B AND2X1_LOC_5/a_36_24# 0.01fF
C13638 AND2X1_LOC_859/Y AND2X1_LOC_621/Y 0.07fF
C13639 AND2X1_LOC_564/B OR2X1_LOC_419/Y 0.10fF
C13640 OR2X1_LOC_7/a_8_216# OR2X1_LOC_56/A 0.02fF
C13641 OR2X1_LOC_333/B OR2X1_LOC_61/Y 0.00fF
C13642 OR2X1_LOC_504/Y AND2X1_LOC_507/a_8_24# 0.01fF
C13643 OR2X1_LOC_417/A AND2X1_LOC_860/A 0.11fF
C13644 OR2X1_LOC_624/B OR2X1_LOC_403/A 0.02fF
C13645 OR2X1_LOC_612/B OR2X1_LOC_39/A 0.03fF
C13646 AND2X1_LOC_721/Y OR2X1_LOC_406/A 0.00fF
C13647 OR2X1_LOC_427/A OR2X1_LOC_279/a_8_216# 0.05fF
C13648 OR2X1_LOC_91/A OR2X1_LOC_77/a_8_216# 0.43fF
C13649 AND2X1_LOC_574/a_8_24# AND2X1_LOC_574/A 0.09fF
C13650 OR2X1_LOC_485/A AND2X1_LOC_644/Y 0.01fF
C13651 OR2X1_LOC_34/A OR2X1_LOC_598/A 0.05fF
C13652 VDD OR2X1_LOC_95/Y 1.41fF
C13653 AND2X1_LOC_580/A AND2X1_LOC_577/A 0.02fF
C13654 GATE_366 OR2X1_LOC_44/Y 0.03fF
C13655 OR2X1_LOC_380/A OR2X1_LOC_588/Y 0.06fF
C13656 AND2X1_LOC_550/A OR2X1_LOC_74/A 0.10fF
C13657 OR2X1_LOC_686/A AND2X1_LOC_684/a_8_24# 0.01fF
C13658 OR2X1_LOC_600/A OR2X1_LOC_411/a_8_216# 0.03fF
C13659 AND2X1_LOC_61/Y OR2X1_LOC_31/Y 0.68fF
C13660 OR2X1_LOC_216/A OR2X1_LOC_121/B 0.23fF
C13661 OR2X1_LOC_54/Y AND2X1_LOC_820/B 0.01fF
C13662 OR2X1_LOC_670/Y OR2X1_LOC_85/A 0.01fF
C13663 OR2X1_LOC_158/A OR2X1_LOC_51/B 0.06fF
C13664 AND2X1_LOC_349/a_8_24# OR2X1_LOC_753/A 0.01fF
C13665 AND2X1_LOC_76/Y OR2X1_LOC_275/A 0.01fF
C13666 OR2X1_LOC_375/A OR2X1_LOC_378/Y 0.21fF
C13667 AND2X1_LOC_717/B OR2X1_LOC_237/Y 0.03fF
C13668 OR2X1_LOC_80/Y OR2X1_LOC_585/A 0.02fF
C13669 OR2X1_LOC_468/Y OR2X1_LOC_449/B 0.03fF
C13670 OR2X1_LOC_538/A D_INPUT_0 0.84fF
C13671 OR2X1_LOC_476/B OR2X1_LOC_61/a_8_216# 0.04fF
C13672 OR2X1_LOC_185/A AND2X1_LOC_69/Y 0.01fF
C13673 OR2X1_LOC_576/a_8_216# OR2X1_LOC_579/A 0.01fF
C13674 AND2X1_LOC_326/B AND2X1_LOC_318/Y 0.02fF
C13675 OR2X1_LOC_135/Y OR2X1_LOC_595/Y 0.02fF
C13676 OR2X1_LOC_6/B D_INPUT_1 0.25fF
C13677 AND2X1_LOC_56/B AND2X1_LOC_329/a_8_24# 0.04fF
C13678 OR2X1_LOC_40/Y OR2X1_LOC_609/Y 0.15fF
C13679 OR2X1_LOC_3/Y AND2X1_LOC_633/a_8_24# 0.01fF
C13680 AND2X1_LOC_627/a_36_24# OR2X1_LOC_598/A 0.00fF
C13681 OR2X1_LOC_139/A OR2X1_LOC_228/Y 0.07fF
C13682 OR2X1_LOC_45/Y OR2X1_LOC_431/a_36_216# 0.00fF
C13683 OR2X1_LOC_312/Y OR2X1_LOC_44/Y 0.03fF
C13684 OR2X1_LOC_543/a_36_216# OR2X1_LOC_161/B 0.02fF
C13685 OR2X1_LOC_625/Y OR2X1_LOC_615/a_36_216# 0.01fF
C13686 AND2X1_LOC_580/A OR2X1_LOC_239/Y 0.03fF
C13687 AND2X1_LOC_337/a_36_24# AND2X1_LOC_318/Y 0.01fF
C13688 AND2X1_LOC_48/A OR2X1_LOC_61/B 0.05fF
C13689 AND2X1_LOC_712/B OR2X1_LOC_427/A 0.94fF
C13690 OR2X1_LOC_484/Y AND2X1_LOC_810/Y 0.26fF
C13691 VDD OR2X1_LOC_207/a_8_216# 0.00fF
C13692 AND2X1_LOC_578/A OR2X1_LOC_680/A 0.07fF
C13693 AND2X1_LOC_12/Y OR2X1_LOC_193/A 0.05fF
C13694 OR2X1_LOC_89/A OR2X1_LOC_591/A 0.02fF
C13695 OR2X1_LOC_119/a_36_216# OR2X1_LOC_118/Y 0.00fF
C13696 OR2X1_LOC_427/A OR2X1_LOC_54/Y 0.41fF
C13697 AND2X1_LOC_40/Y OR2X1_LOC_545/B 0.31fF
C13698 AND2X1_LOC_59/Y OR2X1_LOC_473/Y 0.01fF
C13699 OR2X1_LOC_19/B OR2X1_LOC_394/Y 0.07fF
C13700 OR2X1_LOC_831/A OR2X1_LOC_318/B 0.76fF
C13701 OR2X1_LOC_680/A AND2X1_LOC_632/a_8_24# 0.07fF
C13702 OR2X1_LOC_22/Y OR2X1_LOC_278/Y 0.03fF
C13703 AND2X1_LOC_512/a_36_24# OR2X1_LOC_43/A 0.00fF
C13704 OR2X1_LOC_462/B OR2X1_LOC_461/Y 0.06fF
C13705 OR2X1_LOC_665/Y OR2X1_LOC_7/A 0.03fF
C13706 OR2X1_LOC_7/A AND2X1_LOC_474/Y 0.01fF
C13707 AND2X1_LOC_611/a_8_24# OR2X1_LOC_647/B 0.19fF
C13708 OR2X1_LOC_22/Y AND2X1_LOC_662/B 0.01fF
C13709 OR2X1_LOC_308/Y OR2X1_LOC_727/a_8_216# 0.05fF
C13710 OR2X1_LOC_589/A OR2X1_LOC_72/Y 0.22fF
C13711 OR2X1_LOC_485/A OR2X1_LOC_7/A 0.34fF
C13712 OR2X1_LOC_487/a_8_216# AND2X1_LOC_717/B 0.05fF
C13713 AND2X1_LOC_356/B AND2X1_LOC_337/B 0.01fF
C13714 OR2X1_LOC_600/A AND2X1_LOC_848/A 0.18fF
C13715 OR2X1_LOC_160/A OR2X1_LOC_62/B 0.16fF
C13716 OR2X1_LOC_76/Y OR2X1_LOC_675/A 0.00fF
C13717 OR2X1_LOC_275/A OR2X1_LOC_52/B 0.10fF
C13718 OR2X1_LOC_643/A OR2X1_LOC_404/Y 0.03fF
C13719 AND2X1_LOC_43/B OR2X1_LOC_814/A 0.07fF
C13720 OR2X1_LOC_121/B OR2X1_LOC_468/Y 0.03fF
C13721 OR2X1_LOC_288/A OR2X1_LOC_286/Y 0.12fF
C13722 OR2X1_LOC_22/Y OR2X1_LOC_95/a_8_216# 0.01fF
C13723 AND2X1_LOC_12/Y D_INPUT_0 0.35fF
C13724 OR2X1_LOC_52/Y OR2X1_LOC_753/A 0.20fF
C13725 INPUT_3 OR2X1_LOC_4/a_8_216# 0.01fF
C13726 OR2X1_LOC_223/A OR2X1_LOC_475/B 0.13fF
C13727 OR2X1_LOC_506/A AND2X1_LOC_47/Y 0.02fF
C13728 AND2X1_LOC_838/Y D_INPUT_0 0.03fF
C13729 OR2X1_LOC_160/A OR2X1_LOC_780/B 0.15fF
C13730 AND2X1_LOC_47/Y AND2X1_LOC_695/a_8_24# 0.11fF
C13731 OR2X1_LOC_315/Y OR2X1_LOC_95/Y 0.00fF
C13732 OR2X1_LOC_78/B OR2X1_LOC_358/A 0.07fF
C13733 OR2X1_LOC_276/B AND2X1_LOC_72/Y 0.01fF
C13734 OR2X1_LOC_616/Y OR2X1_LOC_95/Y 0.00fF
C13735 OR2X1_LOC_315/Y OR2X1_LOC_368/A 0.10fF
C13736 OR2X1_LOC_335/Y OR2X1_LOC_318/B 0.00fF
C13737 AND2X1_LOC_1/Y OR2X1_LOC_636/A 0.31fF
C13738 AND2X1_LOC_663/A AND2X1_LOC_222/Y 0.03fF
C13739 OR2X1_LOC_417/A AND2X1_LOC_287/Y 0.01fF
C13740 OR2X1_LOC_26/Y AND2X1_LOC_839/A 0.00fF
C13741 AND2X1_LOC_337/B OR2X1_LOC_22/Y 0.03fF
C13742 OR2X1_LOC_424/a_36_216# AND2X1_LOC_648/B 0.00fF
C13743 AND2X1_LOC_86/B OR2X1_LOC_62/B 0.02fF
C13744 OR2X1_LOC_335/A OR2X1_LOC_722/B 0.02fF
C13745 AND2X1_LOC_40/Y OR2X1_LOC_318/B 0.03fF
C13746 OR2X1_LOC_59/Y OR2X1_LOC_533/A 0.44fF
C13747 OR2X1_LOC_31/Y AND2X1_LOC_852/Y 0.04fF
C13748 AND2X1_LOC_785/A AND2X1_LOC_785/Y 0.51fF
C13749 OR2X1_LOC_31/Y OR2X1_LOC_74/a_36_216# 0.02fF
C13750 OR2X1_LOC_624/B OR2X1_LOC_62/B 0.05fF
C13751 OR2X1_LOC_26/Y OR2X1_LOC_238/a_36_216# 0.02fF
C13752 OR2X1_LOC_689/Y OR2X1_LOC_753/A 0.00fF
C13753 OR2X1_LOC_273/Y OR2X1_LOC_22/Y 0.14fF
C13754 AND2X1_LOC_59/Y OR2X1_LOC_214/B 0.05fF
C13755 AND2X1_LOC_40/Y OR2X1_LOC_854/A 0.01fF
C13756 AND2X1_LOC_95/Y OR2X1_LOC_339/Y 0.01fF
C13757 OR2X1_LOC_213/a_8_216# OR2X1_LOC_375/A 0.01fF
C13758 OR2X1_LOC_247/a_8_216# OR2X1_LOC_805/A 0.02fF
C13759 OR2X1_LOC_579/B D_INPUT_1 2.01fF
C13760 AND2X1_LOC_663/B OR2X1_LOC_46/A 0.07fF
C13761 AND2X1_LOC_59/Y OR2X1_LOC_241/B 0.05fF
C13762 OR2X1_LOC_6/B AND2X1_LOC_789/Y 0.08fF
C13763 OR2X1_LOC_308/a_8_216# OR2X1_LOC_779/B 0.01fF
C13764 AND2X1_LOC_245/a_8_24# OR2X1_LOC_735/B 0.08fF
C13765 OR2X1_LOC_404/Y OR2X1_LOC_113/A 0.03fF
C13766 AND2X1_LOC_389/a_8_24# OR2X1_LOC_95/Y 0.01fF
C13767 AND2X1_LOC_40/Y OR2X1_LOC_344/a_36_216# 0.02fF
C13768 OR2X1_LOC_70/A OR2X1_LOC_53/a_8_216# 0.08fF
C13769 AND2X1_LOC_476/A AND2X1_LOC_634/a_36_24# 0.01fF
C13770 AND2X1_LOC_219/Y OR2X1_LOC_300/a_36_216# 0.01fF
C13771 OR2X1_LOC_485/A OR2X1_LOC_224/a_8_216# 0.01fF
C13772 OR2X1_LOC_22/Y OR2X1_LOC_19/B 0.03fF
C13773 AND2X1_LOC_30/a_36_24# OR2X1_LOC_51/B 0.00fF
C13774 OR2X1_LOC_516/Y AND2X1_LOC_499/a_8_24# 0.02fF
C13775 OR2X1_LOC_685/A OR2X1_LOC_451/B 0.03fF
C13776 VDD INPUT_6 0.46fF
C13777 OR2X1_LOC_709/a_8_216# AND2X1_LOC_64/Y 0.02fF
C13778 OR2X1_LOC_709/A AND2X1_LOC_91/B 0.16fF
C13779 OR2X1_LOC_507/A OR2X1_LOC_508/Y 0.02fF
C13780 OR2X1_LOC_506/Y OR2X1_LOC_392/B 0.09fF
C13781 OR2X1_LOC_118/Y OR2X1_LOC_88/Y 1.25fF
C13782 AND2X1_LOC_227/Y AND2X1_LOC_663/B 0.03fF
C13783 OR2X1_LOC_415/Y OR2X1_LOC_549/A 0.01fF
C13784 AND2X1_LOC_539/Y OR2X1_LOC_829/A 0.01fF
C13785 AND2X1_LOC_174/a_8_24# OR2X1_LOC_172/Y 0.00fF
C13786 OR2X1_LOC_516/Y AND2X1_LOC_658/B 0.05fF
C13787 OR2X1_LOC_177/Y AND2X1_LOC_564/B 0.01fF
C13788 OR2X1_LOC_54/a_8_216# OR2X1_LOC_46/A 0.01fF
C13789 OR2X1_LOC_605/a_8_216# OR2X1_LOC_223/A 0.01fF
C13790 OR2X1_LOC_562/Y OR2X1_LOC_570/a_36_216# 0.03fF
C13791 OR2X1_LOC_176/Y AND2X1_LOC_810/B 0.01fF
C13792 OR2X1_LOC_296/Y OR2X1_LOC_247/a_8_216# 0.01fF
C13793 OR2X1_LOC_49/A OR2X1_LOC_16/A 0.10fF
C13794 OR2X1_LOC_147/A AND2X1_LOC_36/Y 0.00fF
C13795 AND2X1_LOC_3/Y OR2X1_LOC_493/Y 0.01fF
C13796 AND2X1_LOC_3/Y OR2X1_LOC_801/B 0.09fF
C13797 OR2X1_LOC_790/A AND2X1_LOC_22/Y 0.01fF
C13798 OR2X1_LOC_12/Y OR2X1_LOC_766/Y 0.06fF
C13799 AND2X1_LOC_564/B OR2X1_LOC_604/A 0.10fF
C13800 OR2X1_LOC_22/Y OR2X1_LOC_75/Y 0.02fF
C13801 OR2X1_LOC_288/A OR2X1_LOC_532/B 0.01fF
C13802 AND2X1_LOC_802/B OR2X1_LOC_40/Y 0.03fF
C13803 AND2X1_LOC_262/a_8_24# AND2X1_LOC_44/Y 0.01fF
C13804 AND2X1_LOC_571/A OR2X1_LOC_107/a_8_216# 0.47fF
C13805 OR2X1_LOC_262/Y OR2X1_LOC_88/Y 0.01fF
C13806 OR2X1_LOC_696/A OR2X1_LOC_107/Y 0.01fF
C13807 AND2X1_LOC_91/B AND2X1_LOC_70/Y 0.35fF
C13808 OR2X1_LOC_364/B OR2X1_LOC_364/a_8_216# 0.05fF
C13809 AND2X1_LOC_663/B OR2X1_LOC_813/Y 0.05fF
C13810 OR2X1_LOC_208/a_8_216# OR2X1_LOC_228/Y 0.00fF
C13811 OR2X1_LOC_754/a_36_216# OR2X1_LOC_753/Y 0.00fF
C13812 OR2X1_LOC_865/B OR2X1_LOC_576/a_8_216# 0.04fF
C13813 OR2X1_LOC_121/B OR2X1_LOC_205/Y 0.03fF
C13814 OR2X1_LOC_600/A AND2X1_LOC_804/A 0.03fF
C13815 OR2X1_LOC_829/A AND2X1_LOC_771/B 0.00fF
C13816 OR2X1_LOC_6/B OR2X1_LOC_15/a_8_216# 0.02fF
C13817 AND2X1_LOC_50/Y AND2X1_LOC_408/a_8_24# 0.17fF
C13818 OR2X1_LOC_256/A OR2X1_LOC_95/Y 9.35fF
C13819 OR2X1_LOC_70/A AND2X1_LOC_651/B 0.02fF
C13820 OR2X1_LOC_696/A AND2X1_LOC_722/A 0.01fF
C13821 OR2X1_LOC_154/A OR2X1_LOC_704/a_36_216# 0.00fF
C13822 AND2X1_LOC_50/Y AND2X1_LOC_762/a_8_24# 0.01fF
C13823 OR2X1_LOC_186/Y AND2X1_LOC_110/Y 0.13fF
C13824 OR2X1_LOC_121/Y AND2X1_LOC_131/a_8_24# 0.01fF
C13825 AND2X1_LOC_42/B AND2X1_LOC_31/Y 0.02fF
C13826 OR2X1_LOC_456/Y D_GATE_366 0.01fF
C13827 OR2X1_LOC_36/Y OR2X1_LOC_437/A 0.38fF
C13828 OR2X1_LOC_91/A OR2X1_LOC_321/a_8_216# 0.03fF
C13829 OR2X1_LOC_775/a_8_216# OR2X1_LOC_390/B -0.02fF
C13830 OR2X1_LOC_631/A OR2X1_LOC_549/A 0.01fF
C13831 OR2X1_LOC_91/a_8_216# OR2X1_LOC_437/A 0.03fF
C13832 AND2X1_LOC_831/a_8_24# OR2X1_LOC_13/B 0.03fF
C13833 AND2X1_LOC_64/Y AND2X1_LOC_312/a_36_24# 0.01fF
C13834 OR2X1_LOC_154/A OR2X1_LOC_332/a_8_216# 0.05fF
C13835 OR2X1_LOC_674/Y OR2X1_LOC_95/Y 0.01fF
C13836 AND2X1_LOC_47/Y OR2X1_LOC_284/B 0.09fF
C13837 VDD OR2X1_LOC_821/Y 0.12fF
C13838 OR2X1_LOC_44/Y OR2X1_LOC_13/B 0.15fF
C13839 AND2X1_LOC_288/a_8_24# OR2X1_LOC_13/B 0.01fF
C13840 AND2X1_LOC_47/Y D_INPUT_1 12.92fF
C13841 VDD AND2X1_LOC_524/a_8_24# -0.00fF
C13842 AND2X1_LOC_95/Y OR2X1_LOC_500/a_36_216# 0.00fF
C13843 OR2X1_LOC_70/Y OR2X1_LOC_533/A 0.00fF
C13844 OR2X1_LOC_499/B OR2X1_LOC_563/A 0.12fF
C13845 OR2X1_LOC_532/B AND2X1_LOC_72/B 0.02fF
C13846 OR2X1_LOC_648/A AND2X1_LOC_433/a_36_24# 0.01fF
C13847 OR2X1_LOC_278/a_36_216# OR2X1_LOC_71/A 0.00fF
C13848 OR2X1_LOC_693/a_8_216# OR2X1_LOC_744/A 0.01fF
C13849 OR2X1_LOC_95/Y AND2X1_LOC_624/B 0.02fF
C13850 OR2X1_LOC_269/B OR2X1_LOC_590/Y 0.02fF
C13851 AND2X1_LOC_47/Y AND2X1_LOC_48/Y 0.01fF
C13852 AND2X1_LOC_592/Y AND2X1_LOC_732/a_8_24# 0.01fF
C13853 OR2X1_LOC_712/a_8_216# OR2X1_LOC_779/A 0.01fF
C13854 OR2X1_LOC_708/Y OR2X1_LOC_708/a_8_216# -0.00fF
C13855 OR2X1_LOC_691/A OR2X1_LOC_634/A 0.00fF
C13856 OR2X1_LOC_52/B OR2X1_LOC_142/Y 0.03fF
C13857 OR2X1_LOC_97/A OR2X1_LOC_502/A 0.08fF
C13858 OR2X1_LOC_160/B AND2X1_LOC_505/a_36_24# 0.01fF
C13859 OR2X1_LOC_22/A OR2X1_LOC_588/a_8_216# 0.01fF
C13860 OR2X1_LOC_156/A OR2X1_LOC_803/A 0.09fF
C13861 AND2X1_LOC_64/Y OR2X1_LOC_739/A 0.24fF
C13862 OR2X1_LOC_337/A OR2X1_LOC_352/A 0.37fF
C13863 AND2X1_LOC_566/B OR2X1_LOC_744/A 0.03fF
C13864 OR2X1_LOC_3/Y OR2X1_LOC_300/Y 0.03fF
C13865 OR2X1_LOC_759/A AND2X1_LOC_711/A 0.42fF
C13866 OR2X1_LOC_715/B OR2X1_LOC_78/A 2.84fF
C13867 AND2X1_LOC_462/Y OR2X1_LOC_598/A 0.30fF
C13868 AND2X1_LOC_486/Y OR2X1_LOC_816/A 0.47fF
C13869 OR2X1_LOC_681/a_8_216# OR2X1_LOC_51/Y 0.01fF
C13870 OR2X1_LOC_304/a_8_216# OR2X1_LOC_48/B 0.04fF
C13871 OR2X1_LOC_852/a_8_216# OR2X1_LOC_852/B 0.39fF
C13872 OR2X1_LOC_422/a_8_216# OR2X1_LOC_12/Y 0.04fF
C13873 OR2X1_LOC_281/a_8_216# OR2X1_LOC_428/A 0.15fF
C13874 OR2X1_LOC_417/A AND2X1_LOC_562/Y 0.08fF
C13875 OR2X1_LOC_696/A OR2X1_LOC_599/A 0.12fF
C13876 VDD OR2X1_LOC_648/A 0.12fF
C13877 OR2X1_LOC_786/Y OR2X1_LOC_66/a_36_216# 0.01fF
C13878 OR2X1_LOC_78/A OR2X1_LOC_784/B 0.01fF
C13879 OR2X1_LOC_741/Y OR2X1_LOC_787/B 0.02fF
C13880 OR2X1_LOC_790/A OR2X1_LOC_706/A 0.28fF
C13881 OR2X1_LOC_421/A OR2X1_LOC_91/A 0.10fF
C13882 AND2X1_LOC_70/Y OR2X1_LOC_645/a_8_216# 0.01fF
C13883 OR2X1_LOC_106/Y AND2X1_LOC_572/A 0.27fF
C13884 AND2X1_LOC_586/a_36_24# OR2X1_LOC_855/A 0.00fF
C13885 OR2X1_LOC_620/Y OR2X1_LOC_161/B 0.07fF
C13886 OR2X1_LOC_538/A OR2X1_LOC_356/a_8_216# 0.01fF
C13887 OR2X1_LOC_188/Y AND2X1_LOC_59/Y 0.01fF
C13888 AND2X1_LOC_675/Y AND2X1_LOC_806/a_8_24# 0.11fF
C13889 OR2X1_LOC_696/A OR2X1_LOC_93/a_8_216# 0.01fF
C13890 OR2X1_LOC_539/a_8_216# OR2X1_LOC_175/Y 0.01fF
C13891 D_INPUT_1 OR2X1_LOC_598/A 1.05fF
C13892 AND2X1_LOC_693/a_8_24# AND2X1_LOC_18/Y 0.01fF
C13893 OR2X1_LOC_814/A OR2X1_LOC_558/A 0.83fF
C13894 AND2X1_LOC_347/Y OR2X1_LOC_604/A 0.12fF
C13895 AND2X1_LOC_64/Y OR2X1_LOC_269/B 0.15fF
C13896 AND2X1_LOC_339/Y OR2X1_LOC_316/Y 0.00fF
C13897 AND2X1_LOC_541/Y OR2X1_LOC_92/Y 0.05fF
C13898 AND2X1_LOC_360/a_8_24# OR2X1_LOC_40/Y 0.01fF
C13899 AND2X1_LOC_455/B OR2X1_LOC_39/A 0.04fF
C13900 AND2X1_LOC_715/Y OR2X1_LOC_599/A 0.02fF
C13901 AND2X1_LOC_53/Y OR2X1_LOC_193/a_8_216# 0.02fF
C13902 OR2X1_LOC_87/A AND2X1_LOC_7/B 0.61fF
C13903 OR2X1_LOC_497/Y OR2X1_LOC_184/a_36_216# 0.01fF
C13904 AND2X1_LOC_181/a_8_24# OR2X1_LOC_59/Y 0.01fF
C13905 AND2X1_LOC_335/a_8_24# OR2X1_LOC_426/B 0.01fF
C13906 AND2X1_LOC_841/B AND2X1_LOC_476/Y 0.04fF
C13907 OR2X1_LOC_179/Y VDD 0.16fF
C13908 AND2X1_LOC_40/Y OR2X1_LOC_190/a_8_216# 0.14fF
C13909 VDD AND2X1_LOC_253/a_8_24# -0.00fF
C13910 OR2X1_LOC_114/B AND2X1_LOC_40/Y 0.00fF
C13911 AND2X1_LOC_204/Y AND2X1_LOC_205/a_36_24# 0.01fF
C13912 AND2X1_LOC_205/a_8_24# AND2X1_LOC_215/A 0.01fF
C13913 OR2X1_LOC_198/a_8_216# OR2X1_LOC_856/a_8_216# 0.47fF
C13914 AND2X1_LOC_715/Y AND2X1_LOC_854/a_8_24# 0.20fF
C13915 OR2X1_LOC_470/A OR2X1_LOC_161/B 0.02fF
C13916 AND2X1_LOC_570/Y AND2X1_LOC_850/A 0.00fF
C13917 AND2X1_LOC_340/Y OR2X1_LOC_265/Y 0.07fF
C13918 OR2X1_LOC_405/A OR2X1_LOC_151/A 0.25fF
C13919 OR2X1_LOC_652/a_8_216# OR2X1_LOC_435/A 0.01fF
C13920 OR2X1_LOC_113/Y OR2X1_LOC_632/Y 0.01fF
C13921 OR2X1_LOC_427/A OR2X1_LOC_765/Y 0.03fF
C13922 OR2X1_LOC_608/a_8_216# AND2X1_LOC_18/Y 0.04fF
C13923 OR2X1_LOC_323/A OR2X1_LOC_280/Y 0.06fF
C13924 OR2X1_LOC_6/A OR2X1_LOC_428/A 0.23fF
C13925 AND2X1_LOC_251/a_8_24# OR2X1_LOC_843/B 0.00fF
C13926 OR2X1_LOC_154/A OR2X1_LOC_161/B 0.20fF
C13927 OR2X1_LOC_335/a_8_216# OR2X1_LOC_787/Y 0.03fF
C13928 AND2X1_LOC_553/a_8_24# OR2X1_LOC_427/A 0.04fF
C13929 OR2X1_LOC_644/B OR2X1_LOC_691/Y 0.00fF
C13930 OR2X1_LOC_6/B AND2X1_LOC_95/Y 0.51fF
C13931 OR2X1_LOC_106/Y OR2X1_LOC_3/Y 0.01fF
C13932 AND2X1_LOC_719/Y AND2X1_LOC_862/A 0.25fF
C13933 OR2X1_LOC_494/A OR2X1_LOC_89/A 0.03fF
C13934 AND2X1_LOC_650/Y OR2X1_LOC_12/Y 0.00fF
C13935 AND2X1_LOC_541/Y OR2X1_LOC_65/B 0.04fF
C13936 OR2X1_LOC_267/A OR2X1_LOC_161/B 0.01fF
C13937 AND2X1_LOC_719/Y AND2X1_LOC_624/A 0.03fF
C13938 OR2X1_LOC_499/B AND2X1_LOC_628/a_36_24# 0.00fF
C13939 AND2X1_LOC_12/Y OR2X1_LOC_598/Y 0.02fF
C13940 OR2X1_LOC_154/A OR2X1_LOC_514/a_36_216# 0.00fF
C13941 OR2X1_LOC_185/A AND2X1_LOC_18/Y 6.66fF
C13942 AND2X1_LOC_12/Y AND2X1_LOC_131/a_8_24# 0.07fF
C13943 OR2X1_LOC_666/Y OR2X1_LOC_816/A 0.12fF
C13944 OR2X1_LOC_833/B OR2X1_LOC_66/A 0.03fF
C13945 AND2X1_LOC_43/B OR2X1_LOC_410/Y 0.03fF
C13946 AND2X1_LOC_481/a_8_24# AND2X1_LOC_44/Y 0.03fF
C13947 AND2X1_LOC_199/A OR2X1_LOC_44/Y 0.10fF
C13948 AND2X1_LOC_64/Y OR2X1_LOC_215/A 0.01fF
C13949 AND2X1_LOC_563/A AND2X1_LOC_573/A 0.01fF
C13950 AND2X1_LOC_98/Y AND2X1_LOC_99/a_8_24# 0.06fF
C13951 AND2X1_LOC_59/Y OR2X1_LOC_325/B 0.00fF
C13952 AND2X1_LOC_25/a_8_24# INPUT_6 0.04fF
C13953 OR2X1_LOC_485/A OR2X1_LOC_753/a_8_216# -0.00fF
C13954 OR2X1_LOC_532/B AND2X1_LOC_36/Y 3.45fF
C13955 OR2X1_LOC_519/Y OR2X1_LOC_426/B 0.02fF
C13956 AND2X1_LOC_91/B OR2X1_LOC_404/Y 0.10fF
C13957 OR2X1_LOC_602/Y OR2X1_LOC_161/A 0.08fF
C13958 OR2X1_LOC_160/A OR2X1_LOC_468/A 0.07fF
C13959 OR2X1_LOC_303/A OR2X1_LOC_326/B 0.17fF
C13960 AND2X1_LOC_532/a_8_24# OR2X1_LOC_744/A 0.01fF
C13961 OR2X1_LOC_643/A OR2X1_LOC_362/A 0.03fF
C13962 INPUT_5 D_INPUT_4 1.83fF
C13963 OR2X1_LOC_103/Y AND2X1_LOC_113/a_8_24# 0.01fF
C13964 OR2X1_LOC_6/B OR2X1_LOC_99/Y 0.03fF
C13965 OR2X1_LOC_502/A OR2X1_LOC_475/B 0.03fF
C13966 OR2X1_LOC_272/Y OR2X1_LOC_12/Y 0.03fF
C13967 OR2X1_LOC_756/B OR2X1_LOC_814/Y 0.02fF
C13968 OR2X1_LOC_715/B OR2X1_LOC_155/A 0.49fF
C13969 AND2X1_LOC_718/a_8_24# OR2X1_LOC_427/A -0.01fF
C13970 OR2X1_LOC_165/a_8_216# AND2X1_LOC_723/Y 0.02fF
C13971 OR2X1_LOC_778/A OR2X1_LOC_161/B 0.01fF
C13972 OR2X1_LOC_45/B AND2X1_LOC_307/a_8_24# 0.01fF
C13973 OR2X1_LOC_492/Y OR2X1_LOC_529/Y 0.01fF
C13974 AND2X1_LOC_557/a_8_24# OR2X1_LOC_595/A 0.02fF
C13975 AND2X1_LOC_43/B OR2X1_LOC_715/A 0.01fF
C13976 AND2X1_LOC_306/a_8_24# OR2X1_LOC_161/A 0.01fF
C13977 AND2X1_LOC_753/B OR2X1_LOC_651/B 0.00fF
C13978 OR2X1_LOC_369/a_8_216# AND2X1_LOC_784/A 0.04fF
C13979 AND2X1_LOC_715/A OR2X1_LOC_36/Y 2.69fF
C13980 OR2X1_LOC_501/B AND2X1_LOC_43/B 1.05fF
C13981 AND2X1_LOC_319/A OR2X1_LOC_56/A 0.42fF
C13982 OR2X1_LOC_419/Y OR2X1_LOC_437/A 0.19fF
C13983 AND2X1_LOC_375/a_8_24# D_INPUT_5 0.02fF
C13984 OR2X1_LOC_96/Y AND2X1_LOC_673/a_8_24# 0.00fF
C13985 AND2X1_LOC_570/Y OR2X1_LOC_497/a_36_216# 0.00fF
C13986 OR2X1_LOC_164/Y OR2X1_LOC_18/Y 1.16fF
C13987 OR2X1_LOC_58/Y OR2X1_LOC_32/a_8_216# 0.01fF
C13988 AND2X1_LOC_456/B AND2X1_LOC_573/A 0.04fF
C13989 AND2X1_LOC_621/a_8_24# AND2X1_LOC_580/a_8_24# 0.23fF
C13990 OR2X1_LOC_108/a_8_216# OR2X1_LOC_529/Y 0.01fF
C13991 OR2X1_LOC_696/A AND2X1_LOC_866/A 0.10fF
C13992 OR2X1_LOC_831/A OR2X1_LOC_804/B 0.01fF
C13993 OR2X1_LOC_51/Y OR2X1_LOC_670/Y 0.01fF
C13994 OR2X1_LOC_753/A AND2X1_LOC_404/B 0.05fF
C13995 OR2X1_LOC_97/A AND2X1_LOC_48/A 0.03fF
C13996 AND2X1_LOC_83/a_8_24# AND2X1_LOC_51/Y 0.01fF
C13997 OR2X1_LOC_860/Y OR2X1_LOC_865/B 0.14fF
C13998 AND2X1_LOC_713/Y OR2X1_LOC_743/A 0.02fF
C13999 OR2X1_LOC_648/a_8_216# AND2X1_LOC_7/B 0.01fF
C14000 AND2X1_LOC_570/Y OR2X1_LOC_498/Y 0.02fF
C14001 OR2X1_LOC_822/a_8_216# OR2X1_LOC_485/A 0.01fF
C14002 OR2X1_LOC_100/a_8_216# AND2X1_LOC_40/Y 0.01fF
C14003 OR2X1_LOC_585/Y AND2X1_LOC_637/Y 0.82fF
C14004 OR2X1_LOC_516/Y OR2X1_LOC_47/Y 0.03fF
C14005 AND2X1_LOC_859/Y OR2X1_LOC_59/Y 0.02fF
C14006 OR2X1_LOC_62/B OR2X1_LOC_266/A 0.02fF
C14007 OR2X1_LOC_96/Y OR2X1_LOC_74/A 0.02fF
C14008 OR2X1_LOC_3/Y AND2X1_LOC_207/A 0.03fF
C14009 AND2X1_LOC_40/a_36_24# AND2X1_LOC_1/Y 0.00fF
C14010 OR2X1_LOC_446/B OR2X1_LOC_779/B 0.03fF
C14011 OR2X1_LOC_326/B AND2X1_LOC_95/Y 0.09fF
C14012 AND2X1_LOC_12/Y AND2X1_LOC_40/Y 1.34fF
C14013 OR2X1_LOC_235/B OR2X1_LOC_659/B 0.03fF
C14014 OR2X1_LOC_329/a_8_216# OR2X1_LOC_64/Y 0.01fF
C14015 AND2X1_LOC_81/a_8_24# OR2X1_LOC_78/A 0.01fF
C14016 OR2X1_LOC_319/B OR2X1_LOC_703/B 0.03fF
C14017 OR2X1_LOC_316/Y OR2X1_LOC_92/Y 0.03fF
C14018 OR2X1_LOC_160/A AND2X1_LOC_424/a_36_24# 0.00fF
C14019 AND2X1_LOC_95/Y OR2X1_LOC_523/Y 0.01fF
C14020 OR2X1_LOC_70/Y OR2X1_LOC_581/Y 0.28fF
C14021 OR2X1_LOC_599/A AND2X1_LOC_148/a_36_24# 0.00fF
C14022 AND2X1_LOC_566/a_8_24# OR2X1_LOC_91/A 0.01fF
C14023 OR2X1_LOC_51/Y OR2X1_LOC_418/a_8_216# 0.01fF
C14024 OR2X1_LOC_462/B OR2X1_LOC_640/A 0.02fF
C14025 OR2X1_LOC_235/B AND2X1_LOC_8/Y 0.16fF
C14026 OR2X1_LOC_3/Y AND2X1_LOC_658/A 0.03fF
C14027 VDD AND2X1_LOC_136/a_8_24# 0.00fF
C14028 AND2X1_LOC_588/a_8_24# AND2X1_LOC_36/a_8_24# 0.23fF
C14029 OR2X1_LOC_638/B AND2X1_LOC_21/Y 0.01fF
C14030 OR2X1_LOC_212/B OR2X1_LOC_365/B 0.36fF
C14031 OR2X1_LOC_235/B OR2X1_LOC_720/a_36_216# 0.00fF
C14032 AND2X1_LOC_12/Y OR2X1_LOC_810/a_8_216# 0.01fF
C14033 AND2X1_LOC_743/a_8_24# OR2X1_LOC_780/B 0.01fF
C14034 OR2X1_LOC_427/A AND2X1_LOC_453/Y 0.01fF
C14035 OR2X1_LOC_264/Y OR2X1_LOC_217/Y 0.37fF
C14036 AND2X1_LOC_787/A OR2X1_LOC_31/Y 0.00fF
C14037 OR2X1_LOC_48/Y OR2X1_LOC_51/Y 0.03fF
C14038 AND2X1_LOC_858/B AND2X1_LOC_717/B 0.03fF
C14039 OR2X1_LOC_139/A OR2X1_LOC_436/Y 0.15fF
C14040 AND2X1_LOC_807/Y AND2X1_LOC_811/B 0.04fF
C14041 OR2X1_LOC_154/A OR2X1_LOC_61/Y 0.32fF
C14042 OR2X1_LOC_45/B OR2X1_LOC_75/a_8_216# 0.03fF
C14043 OR2X1_LOC_506/Y OR2X1_LOC_532/B 0.01fF
C14044 OR2X1_LOC_643/A OR2X1_LOC_474/Y 0.01fF
C14045 OR2X1_LOC_114/Y OR2X1_LOC_574/a_8_216# 0.01fF
C14046 AND2X1_LOC_456/B OR2X1_LOC_669/Y 0.01fF
C14047 OR2X1_LOC_74/A AND2X1_LOC_663/A 1.74fF
C14048 AND2X1_LOC_140/a_8_24# OR2X1_LOC_56/A 0.17fF
C14049 AND2X1_LOC_662/B OR2X1_LOC_39/A 0.09fF
C14050 OR2X1_LOC_512/A OR2X1_LOC_269/B 0.01fF
C14051 OR2X1_LOC_602/Y AND2X1_LOC_51/Y 0.36fF
C14052 OR2X1_LOC_160/A OR2X1_LOC_128/A 0.05fF
C14053 AND2X1_LOC_53/Y OR2X1_LOC_713/A 0.03fF
C14054 OR2X1_LOC_31/Y AND2X1_LOC_457/a_36_24# 0.00fF
C14055 AND2X1_LOC_12/Y OR2X1_LOC_537/A 0.13fF
C14056 OR2X1_LOC_189/a_36_216# AND2X1_LOC_565/Y 0.00fF
C14057 OR2X1_LOC_118/Y OR2X1_LOC_67/A 0.00fF
C14058 AND2X1_LOC_849/A AND2X1_LOC_244/a_36_24# 0.00fF
C14059 OR2X1_LOC_252/Y AND2X1_LOC_624/A 0.09fF
C14060 OR2X1_LOC_641/a_8_216# OR2X1_LOC_643/Y 0.01fF
C14061 AND2X1_LOC_59/Y OR2X1_LOC_405/Y 0.00fF
C14062 AND2X1_LOC_80/a_8_24# OR2X1_LOC_377/A 0.03fF
C14063 AND2X1_LOC_737/a_36_24# OR2X1_LOC_52/B 0.00fF
C14064 OR2X1_LOC_235/B OR2X1_LOC_291/A 0.05fF
C14065 OR2X1_LOC_113/A OR2X1_LOC_362/A 0.01fF
C14066 OR2X1_LOC_850/B OR2X1_LOC_287/B 0.63fF
C14067 OR2X1_LOC_47/Y OR2X1_LOC_373/a_8_216# 0.01fF
C14068 AND2X1_LOC_577/Y AND2X1_LOC_578/a_8_24# 0.03fF
C14069 OR2X1_LOC_375/A OR2X1_LOC_209/a_8_216# 0.00fF
C14070 AND2X1_LOC_684/a_8_24# OR2X1_LOC_161/B 0.01fF
C14071 OR2X1_LOC_624/B OR2X1_LOC_659/A 0.01fF
C14072 OR2X1_LOC_26/Y OR2X1_LOC_427/A 0.63fF
C14073 OR2X1_LOC_807/Y OR2X1_LOC_269/B 0.01fF
C14074 AND2X1_LOC_228/Y OR2X1_LOC_265/Y 0.01fF
C14075 AND2X1_LOC_817/B OR2X1_LOC_847/a_8_216# 0.01fF
C14076 AND2X1_LOC_12/Y OR2X1_LOC_848/A 0.46fF
C14077 OR2X1_LOC_348/Y OR2X1_LOC_814/A 0.02fF
C14078 OR2X1_LOC_760/Y OR2X1_LOC_16/A 0.01fF
C14079 OR2X1_LOC_349/a_8_216# OR2X1_LOC_814/A 0.01fF
C14080 OR2X1_LOC_87/A OR2X1_LOC_805/A 0.14fF
C14081 AND2X1_LOC_12/Y OR2X1_LOC_859/B 0.50fF
C14082 AND2X1_LOC_390/B OR2X1_LOC_92/Y 0.08fF
C14083 OR2X1_LOC_823/Y OR2X1_LOC_26/Y 0.02fF
C14084 AND2X1_LOC_734/Y OR2X1_LOC_527/Y 0.00fF
C14085 OR2X1_LOC_427/A OR2X1_LOC_89/A 15.38fF
C14086 AND2X1_LOC_174/a_8_24# OR2X1_LOC_52/B 0.02fF
C14087 OR2X1_LOC_276/B OR2X1_LOC_719/B 0.02fF
C14088 OR2X1_LOC_160/A OR2X1_LOC_449/B 0.07fF
C14089 OR2X1_LOC_271/Y OR2X1_LOC_316/Y 0.59fF
C14090 AND2X1_LOC_364/Y AND2X1_LOC_863/A 0.16fF
C14091 OR2X1_LOC_271/B AND2X1_LOC_318/a_36_24# 0.00fF
C14092 OR2X1_LOC_256/a_8_216# OR2X1_LOC_7/A 0.01fF
C14093 AND2X1_LOC_22/Y AND2X1_LOC_289/a_36_24# 0.00fF
C14094 AND2X1_LOC_211/B AND2X1_LOC_662/B 0.07fF
C14095 AND2X1_LOC_472/B OR2X1_LOC_39/A 0.03fF
C14096 OR2X1_LOC_194/B AND2X1_LOC_3/Y 0.01fF
C14097 OR2X1_LOC_198/a_8_216# OR2X1_LOC_198/A 0.13fF
C14098 AND2X1_LOC_22/Y OR2X1_LOC_339/Y 0.49fF
C14099 AND2X1_LOC_462/B AND2X1_LOC_219/A 0.15fF
C14100 AND2X1_LOC_392/A AND2X1_LOC_227/Y 0.03fF
C14101 OR2X1_LOC_695/Y OR2X1_LOC_31/Y 0.01fF
C14102 OR2X1_LOC_217/Y OR2X1_LOC_643/A 3.01fF
C14103 AND2X1_LOC_717/B AND2X1_LOC_573/A 0.01fF
C14104 OR2X1_LOC_217/Y OR2X1_LOC_124/Y 0.00fF
C14105 OR2X1_LOC_646/B D_INPUT_1 0.09fF
C14106 OR2X1_LOC_502/A OR2X1_LOC_415/A 0.01fF
C14107 OR2X1_LOC_3/Y AND2X1_LOC_847/Y 0.01fF
C14108 OR2X1_LOC_166/Y OR2X1_LOC_167/Y 0.20fF
C14109 OR2X1_LOC_36/Y OR2X1_LOC_753/A 0.06fF
C14110 AND2X1_LOC_387/B AND2X1_LOC_43/B 0.07fF
C14111 AND2X1_LOC_95/Y OR2X1_LOC_33/a_36_216# 0.00fF
C14112 AND2X1_LOC_31/Y AND2X1_LOC_224/a_8_24# 0.01fF
C14113 OR2X1_LOC_866/B OR2X1_LOC_557/a_8_216# 0.42fF
C14114 OR2X1_LOC_151/A OR2X1_LOC_330/a_8_216# 0.02fF
C14115 OR2X1_LOC_633/a_8_216# OR2X1_LOC_532/B 0.01fF
C14116 OR2X1_LOC_805/A OR2X1_LOC_216/a_8_216# 0.01fF
C14117 AND2X1_LOC_486/Y AND2X1_LOC_727/A 0.03fF
C14118 AND2X1_LOC_12/Y OR2X1_LOC_475/Y 0.02fF
C14119 AND2X1_LOC_44/Y OR2X1_LOC_512/Y 0.01fF
C14120 OR2X1_LOC_273/Y OR2X1_LOC_39/A 0.03fF
C14121 OR2X1_LOC_36/Y OR2X1_LOC_754/a_8_216# 0.03fF
C14122 OR2X1_LOC_563/A OR2X1_LOC_348/B 0.03fF
C14123 OR2X1_LOC_523/A OR2X1_LOC_523/a_8_216# 0.01fF
C14124 AND2X1_LOC_791/a_8_24# AND2X1_LOC_789/Y 0.04fF
C14125 OR2X1_LOC_352/a_36_216# OR2X1_LOC_578/B 0.00fF
C14126 AND2X1_LOC_548/a_36_24# OR2X1_LOC_680/A 0.00fF
C14127 OR2X1_LOC_205/a_8_216# AND2X1_LOC_3/Y 0.02fF
C14128 AND2X1_LOC_363/A OR2X1_LOC_89/A 0.04fF
C14129 AND2X1_LOC_345/a_8_24# OR2X1_LOC_748/A 0.00fF
C14130 OR2X1_LOC_160/A OR2X1_LOC_121/B 0.17fF
C14131 D_INPUT_0 AND2X1_LOC_852/B 0.13fF
C14132 OR2X1_LOC_574/A OR2X1_LOC_593/A 0.08fF
C14133 OR2X1_LOC_80/A OR2X1_LOC_548/B 0.03fF
C14134 OR2X1_LOC_864/A AND2X1_LOC_42/B 0.03fF
C14135 AND2X1_LOC_863/Y OR2X1_LOC_92/Y 0.07fF
C14136 AND2X1_LOC_122/a_36_24# OR2X1_LOC_203/Y 0.01fF
C14137 OR2X1_LOC_19/B OR2X1_LOC_39/A 0.98fF
C14138 AND2X1_LOC_702/Y OR2X1_LOC_304/Y 0.01fF
C14139 AND2X1_LOC_721/A OR2X1_LOC_56/A 0.03fF
C14140 D_INPUT_0 OR2X1_LOC_48/B 0.07fF
C14141 OR2X1_LOC_64/Y OR2X1_LOC_235/a_8_216# 0.18fF
C14142 AND2X1_LOC_486/Y OR2X1_LOC_95/Y 0.03fF
C14143 AND2X1_LOC_42/B OR2X1_LOC_240/A 0.16fF
C14144 AND2X1_LOC_47/Y OR2X1_LOC_737/A 0.07fF
C14145 OR2X1_LOC_70/A OR2X1_LOC_581/Y 0.09fF
C14146 AND2X1_LOC_95/Y OR2X1_LOC_287/a_36_216# 0.01fF
C14147 OR2X1_LOC_18/Y D_INPUT_0 1.81fF
C14148 OR2X1_LOC_808/a_8_216# OR2X1_LOC_440/A 0.06fF
C14149 OR2X1_LOC_246/A OR2X1_LOC_767/a_36_216# 0.15fF
C14150 OR2X1_LOC_377/A AND2X1_LOC_15/a_8_24# 0.05fF
C14151 OR2X1_LOC_440/A OR2X1_LOC_733/a_8_216# 0.14fF
C14152 OR2X1_LOC_45/B OR2X1_LOC_13/B 0.17fF
C14153 AND2X1_LOC_95/Y AND2X1_LOC_47/Y 0.21fF
C14154 AND2X1_LOC_59/Y D_INPUT_0 0.61fF
C14155 OR2X1_LOC_417/A AND2X1_LOC_287/a_8_24# 0.01fF
C14156 OR2X1_LOC_709/A OR2X1_LOC_446/B 0.40fF
C14157 OR2X1_LOC_633/Y AND2X1_LOC_47/Y 7.73fF
C14158 OR2X1_LOC_426/a_8_216# OR2X1_LOC_427/A 0.01fF
C14159 D_INPUT_4 OR2X1_LOC_17/a_8_216# 0.02fF
C14160 AND2X1_LOC_660/A AND2X1_LOC_649/a_8_24# 0.05fF
C14161 OR2X1_LOC_786/Y OR2X1_LOC_785/B 0.03fF
C14162 OR2X1_LOC_92/a_8_216# OR2X1_LOC_63/a_8_216# 0.47fF
C14163 OR2X1_LOC_186/Y OR2X1_LOC_550/B 0.05fF
C14164 AND2X1_LOC_738/B OR2X1_LOC_331/Y 0.27fF
C14165 OR2X1_LOC_177/Y OR2X1_LOC_437/A 0.05fF
C14166 OR2X1_LOC_78/B OR2X1_LOC_398/a_36_216# 0.02fF
C14167 AND2X1_LOC_706/Y OR2X1_LOC_424/Y 0.01fF
C14168 OR2X1_LOC_102/a_8_216# OR2X1_LOC_13/B 0.01fF
C14169 OR2X1_LOC_87/A AND2X1_LOC_441/a_8_24# 0.01fF
C14170 OR2X1_LOC_75/Y OR2X1_LOC_39/A 0.03fF
C14171 OR2X1_LOC_12/Y OR2X1_LOC_248/A 0.05fF
C14172 OR2X1_LOC_810/A OR2X1_LOC_814/A 2.23fF
C14173 OR2X1_LOC_506/A AND2X1_LOC_420/a_8_24# 0.05fF
C14174 OR2X1_LOC_43/A OR2X1_LOC_167/Y 0.02fF
C14175 OR2X1_LOC_280/Y AND2X1_LOC_844/a_36_24# 0.01fF
C14176 OR2X1_LOC_427/A AND2X1_LOC_451/a_8_24# 0.01fF
C14177 AND2X1_LOC_31/Y OR2X1_LOC_778/a_8_216# 0.01fF
C14178 AND2X1_LOC_840/B AND2X1_LOC_675/A 0.10fF
C14179 OR2X1_LOC_255/a_8_216# OR2X1_LOC_585/A 0.01fF
C14180 OR2X1_LOC_3/Y AND2X1_LOC_814/a_8_24# 0.01fF
C14181 OR2X1_LOC_532/B OR2X1_LOC_346/B 0.23fF
C14182 OR2X1_LOC_726/A OR2X1_LOC_550/B 0.11fF
C14183 AND2X1_LOC_729/B OR2X1_LOC_43/a_8_216# 0.01fF
C14184 OR2X1_LOC_811/A OR2X1_LOC_366/a_8_216# 0.11fF
C14185 OR2X1_LOC_604/A OR2X1_LOC_437/A 0.19fF
C14186 AND2X1_LOC_3/a_8_24# AND2X1_LOC_430/B 0.19fF
C14187 OR2X1_LOC_95/Y OR2X1_LOC_248/Y 0.04fF
C14188 AND2X1_LOC_56/B OR2X1_LOC_276/B 0.16fF
C14189 OR2X1_LOC_194/B OR2X1_LOC_194/a_8_216# 0.06fF
C14190 OR2X1_LOC_22/Y OR2X1_LOC_754/A 0.44fF
C14191 AND2X1_LOC_70/Y OR2X1_LOC_446/B 0.02fF
C14192 OR2X1_LOC_663/A AND2X1_LOC_31/Y 0.06fF
C14193 AND2X1_LOC_571/A AND2X1_LOC_571/a_8_24# 0.00fF
C14194 AND2X1_LOC_537/Y AND2X1_LOC_729/B 0.02fF
C14195 OR2X1_LOC_22/Y OR2X1_LOC_275/A 0.07fF
C14196 OR2X1_LOC_672/a_8_216# AND2X1_LOC_789/Y 0.01fF
C14197 AND2X1_LOC_70/Y OR2X1_LOC_303/B 0.06fF
C14198 VDD OR2X1_LOC_112/A 0.21fF
C14199 AND2X1_LOC_95/Y OR2X1_LOC_598/A 0.22fF
C14200 VDD OR2X1_LOC_730/B 0.05fF
C14201 OR2X1_LOC_789/B OR2X1_LOC_801/B 0.04fF
C14202 OR2X1_LOC_160/B OR2X1_LOC_712/B 0.01fF
C14203 OR2X1_LOC_118/Y AND2X1_LOC_216/A 0.02fF
C14204 OR2X1_LOC_633/Y OR2X1_LOC_598/A 0.03fF
C14205 OR2X1_LOC_602/B AND2X1_LOC_51/Y 0.01fF
C14206 OR2X1_LOC_856/B OR2X1_LOC_750/Y 0.02fF
C14207 OR2X1_LOC_19/B AND2X1_LOC_672/B 0.02fF
C14208 OR2X1_LOC_665/Y OR2X1_LOC_615/Y 0.03fF
C14209 OR2X1_LOC_76/B AND2X1_LOC_31/Y 0.01fF
C14210 OR2X1_LOC_203/Y OR2X1_LOC_66/a_8_216# 0.02fF
C14211 AND2X1_LOC_43/B OR2X1_LOC_318/B 0.03fF
C14212 OR2X1_LOC_703/A OR2X1_LOC_303/B 0.01fF
C14213 OR2X1_LOC_485/A OR2X1_LOC_615/Y 0.20fF
C14214 OR2X1_LOC_696/A OR2X1_LOC_40/Y 0.16fF
C14215 OR2X1_LOC_147/B OR2X1_LOC_367/B 0.54fF
C14216 AND2X1_LOC_866/A AND2X1_LOC_663/B 0.02fF
C14217 OR2X1_LOC_167/a_36_216# AND2X1_LOC_715/Y 0.01fF
C14218 AND2X1_LOC_621/Y AND2X1_LOC_657/A 0.07fF
C14219 OR2X1_LOC_356/B OR2X1_LOC_356/a_8_216# 0.08fF
C14220 AND2X1_LOC_543/Y AND2X1_LOC_476/Y 0.04fF
C14221 OR2X1_LOC_47/Y AND2X1_LOC_651/B 0.01fF
C14222 D_INPUT_5 OR2X1_LOC_376/a_8_216# 0.01fF
C14223 AND2X1_LOC_57/Y VDD 0.00fF
C14224 AND2X1_LOC_56/B OR2X1_LOC_740/a_8_216# 0.03fF
C14225 AND2X1_LOC_555/Y AND2X1_LOC_555/a_36_24# 0.00fF
C14226 OR2X1_LOC_169/B OR2X1_LOC_568/A 0.06fF
C14227 AND2X1_LOC_91/B OR2X1_LOC_362/A 0.03fF
C14228 AND2X1_LOC_773/Y OR2X1_LOC_135/Y 0.03fF
C14229 OR2X1_LOC_294/Y AND2X1_LOC_44/Y 0.01fF
C14230 OR2X1_LOC_364/A AND2X1_LOC_31/Y 0.34fF
C14231 OR2X1_LOC_185/Y AND2X1_LOC_31/Y 0.22fF
C14232 AND2X1_LOC_809/a_8_24# AND2X1_LOC_810/B 0.00fF
C14233 AND2X1_LOC_802/Y AND2X1_LOC_809/a_36_24# 0.01fF
C14234 AND2X1_LOC_91/B OR2X1_LOC_832/a_8_216# 0.28fF
C14235 AND2X1_LOC_383/a_8_24# OR2X1_LOC_40/Y 0.01fF
C14236 AND2X1_LOC_574/Y VDD 0.05fF
C14237 AND2X1_LOC_28/a_36_24# INPUT_1 0.01fF
C14238 OR2X1_LOC_149/B VDD 0.12fF
C14239 OR2X1_LOC_416/A INPUT_1 0.03fF
C14240 OR2X1_LOC_6/B AND2X1_LOC_22/Y 0.07fF
C14241 OR2X1_LOC_641/A AND2X1_LOC_44/Y 0.03fF
C14242 OR2X1_LOC_139/A OR2X1_LOC_160/B 0.74fF
C14243 OR2X1_LOC_651/A AND2X1_LOC_7/Y 0.12fF
C14244 AND2X1_LOC_18/Y OR2X1_LOC_577/Y 0.02fF
C14245 OR2X1_LOC_106/Y OR2X1_LOC_329/B 0.17fF
C14246 OR2X1_LOC_714/Y AND2X1_LOC_36/Y 0.02fF
C14247 VDD AND2X1_LOC_358/Y 0.46fF
C14248 AND2X1_LOC_24/a_8_24# OR2X1_LOC_338/A 0.10fF
C14249 OR2X1_LOC_555/A AND2X1_LOC_257/a_36_24# 0.00fF
C14250 OR2X1_LOC_479/Y OR2X1_LOC_228/Y 0.01fF
C14251 OR2X1_LOC_505/a_8_216# AND2X1_LOC_508/B 0.01fF
C14252 OR2X1_LOC_19/B AND2X1_LOC_761/a_8_24# 0.01fF
C14253 AND2X1_LOC_476/Y OR2X1_LOC_322/Y 0.12fF
C14254 VDD OR2X1_LOC_693/Y 0.16fF
C14255 OR2X1_LOC_415/a_8_216# OR2X1_LOC_598/A 0.03fF
C14256 OR2X1_LOC_6/B OR2X1_LOC_621/A 0.04fF
C14257 AND2X1_LOC_633/Y AND2X1_LOC_215/A 0.02fF
C14258 AND2X1_LOC_64/Y OR2X1_LOC_475/a_8_216# 0.04fF
C14259 OR2X1_LOC_318/Y OR2X1_LOC_390/B 0.07fF
C14260 OR2X1_LOC_39/A OR2X1_LOC_504/a_8_216# 0.01fF
C14261 AND2X1_LOC_541/Y OR2X1_LOC_600/A 0.04fF
C14262 AND2X1_LOC_849/A AND2X1_LOC_563/Y 0.02fF
C14263 OR2X1_LOC_392/B OR2X1_LOC_392/A 0.05fF
C14264 OR2X1_LOC_175/Y OR2X1_LOC_502/A 0.07fF
C14265 OR2X1_LOC_769/A AND2X1_LOC_585/a_36_24# 0.00fF
C14266 OR2X1_LOC_227/a_8_216# OR2X1_LOC_641/B 0.00fF
C14267 AND2X1_LOC_70/Y OR2X1_LOC_719/B 0.10fF
C14268 AND2X1_LOC_182/A OR2X1_LOC_51/Y 0.01fF
C14269 OR2X1_LOC_158/A OR2X1_LOC_666/A 0.06fF
C14270 AND2X1_LOC_214/A OR2X1_LOC_16/A 0.33fF
C14271 OR2X1_LOC_696/A OR2X1_LOC_424/a_8_216# 0.03fF
C14272 AND2X1_LOC_658/A AND2X1_LOC_477/Y 0.07fF
C14273 OR2X1_LOC_686/B OR2X1_LOC_686/a_8_216# 0.00fF
C14274 OR2X1_LOC_291/Y AND2X1_LOC_215/a_8_24# 0.13fF
C14275 OR2X1_LOC_748/A AND2X1_LOC_792/B 0.00fF
C14276 OR2X1_LOC_538/A OR2X1_LOC_356/A 0.00fF
C14277 OR2X1_LOC_435/B OR2X1_LOC_435/A 1.13fF
C14278 AND2X1_LOC_719/Y AND2X1_LOC_286/a_36_24# 0.01fF
C14279 OR2X1_LOC_694/Y OR2X1_LOC_695/Y 0.21fF
C14280 OR2X1_LOC_54/Y OR2X1_LOC_80/A 0.10fF
C14281 OR2X1_LOC_696/A OR2X1_LOC_618/a_8_216# 0.01fF
C14282 OR2X1_LOC_624/a_8_216# OR2X1_LOC_113/B 0.01fF
C14283 OR2X1_LOC_502/A OR2X1_LOC_375/Y 0.00fF
C14284 OR2X1_LOC_421/a_8_216# OR2X1_LOC_421/Y 0.00fF
C14285 AND2X1_LOC_64/Y OR2X1_LOC_539/Y 0.09fF
C14286 AND2X1_LOC_22/Y OR2X1_LOC_523/Y 0.01fF
C14287 AND2X1_LOC_501/Y AND2X1_LOC_657/Y 0.04fF
C14288 OR2X1_LOC_40/Y AND2X1_LOC_851/a_36_24# 0.00fF
C14289 OR2X1_LOC_604/A OR2X1_LOC_90/a_36_216# 0.01fF
C14290 OR2X1_LOC_502/A OR2X1_LOC_713/A 0.07fF
C14291 OR2X1_LOC_335/Y OR2X1_LOC_182/B 0.00fF
C14292 OR2X1_LOC_6/B OR2X1_LOC_244/B 0.03fF
C14293 OR2X1_LOC_792/Y OR2X1_LOC_580/B 0.26fF
C14294 AND2X1_LOC_95/Y OR2X1_LOC_34/A 0.00fF
C14295 AND2X1_LOC_570/Y AND2X1_LOC_657/Y 0.05fF
C14296 AND2X1_LOC_160/Y OR2X1_LOC_51/Y 0.07fF
C14297 AND2X1_LOC_543/a_36_24# AND2X1_LOC_476/Y 0.00fF
C14298 AND2X1_LOC_48/A OR2X1_LOC_193/a_8_216# 0.01fF
C14299 AND2X1_LOC_716/Y OR2X1_LOC_158/A 0.07fF
C14300 AND2X1_LOC_544/a_8_24# AND2X1_LOC_476/Y 0.02fF
C14301 AND2X1_LOC_350/B OR2X1_LOC_18/Y 0.01fF
C14302 OR2X1_LOC_744/a_8_216# OR2X1_LOC_39/A 0.01fF
C14303 OR2X1_LOC_701/Y OR2X1_LOC_428/A 0.00fF
C14304 AND2X1_LOC_706/Y AND2X1_LOC_841/B 0.02fF
C14305 OR2X1_LOC_481/A AND2X1_LOC_789/Y 0.07fF
C14306 OR2X1_LOC_676/Y AND2X1_LOC_41/A 0.12fF
C14307 OR2X1_LOC_696/A OR2X1_LOC_7/A 0.36fF
C14308 OR2X1_LOC_545/B OR2X1_LOC_367/B 0.08fF
C14309 OR2X1_LOC_613/Y AND2X1_LOC_580/a_8_24# 0.01fF
C14310 AND2X1_LOC_40/Y OR2X1_LOC_182/B 0.03fF
C14311 OR2X1_LOC_541/B AND2X1_LOC_256/a_8_24# 0.00fF
C14312 OR2X1_LOC_756/Y VDD 0.05fF
C14313 OR2X1_LOC_48/B AND2X1_LOC_771/B 0.01fF
C14314 OR2X1_LOC_158/A AND2X1_LOC_654/Y 0.07fF
C14315 OR2X1_LOC_427/A AND2X1_LOC_605/a_8_24# 0.02fF
C14316 OR2X1_LOC_121/B OR2X1_LOC_532/Y 0.28fF
C14317 AND2X1_LOC_552/A OR2X1_LOC_427/A 0.01fF
C14318 OR2X1_LOC_703/A OR2X1_LOC_542/B 0.00fF
C14319 AND2X1_LOC_706/a_36_24# OR2X1_LOC_48/B 0.01fF
C14320 AND2X1_LOC_521/a_8_24# AND2X1_LOC_95/Y 0.01fF
C14321 AND2X1_LOC_738/B AND2X1_LOC_605/Y 0.01fF
C14322 OR2X1_LOC_438/Y VDD 0.10fF
C14323 OR2X1_LOC_864/A AND2X1_LOC_224/a_8_24# 0.03fF
C14324 OR2X1_LOC_18/Y AND2X1_LOC_771/B 0.00fF
C14325 OR2X1_LOC_105/Y VDD 0.13fF
C14326 AND2X1_LOC_706/a_36_24# OR2X1_LOC_18/Y 0.00fF
C14327 OR2X1_LOC_194/Y AND2X1_LOC_44/Y 0.01fF
C14328 OR2X1_LOC_121/B OR2X1_LOC_212/B 0.08fF
C14329 AND2X1_LOC_207/a_8_24# INPUT_0 0.01fF
C14330 OR2X1_LOC_834/A AND2X1_LOC_41/A 0.02fF
C14331 OR2X1_LOC_47/Y AND2X1_LOC_793/B 0.01fF
C14332 AND2X1_LOC_421/a_8_24# OR2X1_LOC_66/A 0.03fF
C14333 OR2X1_LOC_61/A OR2X1_LOC_358/B 0.02fF
C14334 AND2X1_LOC_42/B OR2X1_LOC_397/a_8_216# 0.12fF
C14335 OR2X1_LOC_508/a_8_216# OR2X1_LOC_375/A 0.01fF
C14336 OR2X1_LOC_114/Y AND2X1_LOC_44/Y 0.01fF
C14337 OR2X1_LOC_44/Y OR2X1_LOC_428/A 0.23fF
C14338 OR2X1_LOC_375/A OR2X1_LOC_486/Y 0.03fF
C14339 OR2X1_LOC_267/a_8_216# OR2X1_LOC_161/B 0.15fF
C14340 AND2X1_LOC_715/Y OR2X1_LOC_7/A 0.07fF
C14341 AND2X1_LOC_59/Y OR2X1_LOC_831/A 0.01fF
C14342 VDD OR2X1_LOC_427/Y 0.00fF
C14343 OR2X1_LOC_485/A AND2X1_LOC_242/B 0.02fF
C14344 OR2X1_LOC_709/A AND2X1_LOC_56/B 0.06fF
C14345 OR2X1_LOC_692/a_8_216# OR2X1_LOC_744/A 0.01fF
C14346 VDD OR2X1_LOC_465/Y 0.12fF
C14347 OR2X1_LOC_44/Y OR2X1_LOC_595/A 0.03fF
C14348 AND2X1_LOC_47/Y OR2X1_LOC_788/B 0.00fF
C14349 OR2X1_LOC_526/Y AND2X1_LOC_546/a_8_24# 0.00fF
C14350 OR2X1_LOC_744/A OR2X1_LOC_92/Y 0.17fF
C14351 AND2X1_LOC_47/Y AND2X1_LOC_41/Y 0.00fF
C14352 AND2X1_LOC_191/Y GATE_579 0.17fF
C14353 AND2X1_LOC_59/Y OR2X1_LOC_598/Y 0.03fF
C14354 OR2X1_LOC_529/a_8_216# OR2X1_LOC_600/A 0.03fF
C14355 OR2X1_LOC_97/A AND2X1_LOC_3/Y 0.03fF
C14356 INPUT_1 OR2X1_LOC_268/Y 0.01fF
C14357 AND2X1_LOC_42/B OR2X1_LOC_121/A 0.03fF
C14358 OR2X1_LOC_856/B OR2X1_LOC_809/B 0.07fF
C14359 OR2X1_LOC_151/A OR2X1_LOC_653/A 0.69fF
C14360 VDD OR2X1_LOC_632/A -0.00fF
C14361 OR2X1_LOC_375/A OR2X1_LOC_542/a_36_216# 0.00fF
C14362 AND2X1_LOC_848/Y AND2X1_LOC_243/Y 0.00fF
C14363 OR2X1_LOC_84/Y OR2X1_LOC_80/A 0.02fF
C14364 AND2X1_LOC_59/Y OR2X1_LOC_356/a_8_216# 0.01fF
C14365 AND2X1_LOC_517/a_36_24# AND2X1_LOC_18/Y 0.00fF
C14366 AND2X1_LOC_425/Y AND2X1_LOC_581/a_8_24# 0.01fF
C14367 VDD AND2X1_LOC_621/Y 0.98fF
C14368 OR2X1_LOC_158/A GATE_366 0.03fF
C14369 OR2X1_LOC_532/B OR2X1_LOC_469/B 0.03fF
C14370 AND2X1_LOC_711/Y GATE_579 0.04fF
C14371 OR2X1_LOC_600/A OR2X1_LOC_316/Y 0.03fF
C14372 OR2X1_LOC_99/Y OR2X1_LOC_646/B 0.01fF
C14373 OR2X1_LOC_656/B OR2X1_LOC_78/A 0.01fF
C14374 AND2X1_LOC_31/Y OR2X1_LOC_552/A 0.13fF
C14375 OR2X1_LOC_493/a_8_216# OR2X1_LOC_805/A 0.04fF
C14376 OR2X1_LOC_330/Y OR2X1_LOC_808/B 0.35fF
C14377 OR2X1_LOC_190/A OR2X1_LOC_254/B 0.09fF
C14378 OR2X1_LOC_43/A OR2X1_LOC_382/a_36_216# -0.01fF
C14379 INPUT_0 OR2X1_LOC_194/B 0.00fF
C14380 AND2X1_LOC_474/A OR2X1_LOC_278/Y 0.01fF
C14381 OR2X1_LOC_637/A OR2X1_LOC_637/B 0.14fF
C14382 OR2X1_LOC_528/Y AND2X1_LOC_569/A 0.01fF
C14383 OR2X1_LOC_705/B OR2X1_LOC_546/A 0.00fF
C14384 AND2X1_LOC_104/a_36_24# OR2X1_LOC_78/A 0.01fF
C14385 OR2X1_LOC_227/a_8_216# OR2X1_LOC_227/A 0.47fF
C14386 OR2X1_LOC_18/Y AND2X1_LOC_471/Y 0.04fF
C14387 OR2X1_LOC_744/A OR2X1_LOC_65/B 0.04fF
C14388 AND2X1_LOC_810/A AND2X1_LOC_212/B 0.15fF
C14389 AND2X1_LOC_12/a_8_24# AND2X1_LOC_11/Y 0.01fF
C14390 OR2X1_LOC_469/Y OR2X1_LOC_478/a_8_216# 0.06fF
C14391 OR2X1_LOC_91/A AND2X1_LOC_452/Y 0.02fF
C14392 OR2X1_LOC_405/A OR2X1_LOC_174/A 0.13fF
C14393 AND2X1_LOC_31/Y AND2X1_LOC_432/a_8_24# 0.01fF
C14394 OR2X1_LOC_604/A OR2X1_LOC_753/A 0.10fF
C14395 AND2X1_LOC_59/Y OR2X1_LOC_795/B 0.01fF
C14396 OR2X1_LOC_213/A OR2X1_LOC_803/A 0.73fF
C14397 OR2X1_LOC_457/a_8_216# OR2X1_LOC_741/Y 0.01fF
C14398 AND2X1_LOC_80/a_8_24# OR2X1_LOC_78/B 0.05fF
C14399 AND2X1_LOC_70/Y AND2X1_LOC_56/B 1.47fF
C14400 OR2X1_LOC_175/Y AND2X1_LOC_48/A 0.03fF
C14401 OR2X1_LOC_538/A AND2X1_LOC_43/B 0.18fF
C14402 AND2X1_LOC_31/Y OR2X1_LOC_578/B 0.03fF
C14403 AND2X1_LOC_480/A AND2X1_LOC_223/A 0.10fF
C14404 OR2X1_LOC_450/B OR2X1_LOC_449/B 0.39fF
C14405 AND2X1_LOC_110/Y OR2X1_LOC_574/A 0.03fF
C14406 AND2X1_LOC_642/Y AND2X1_LOC_649/a_8_24# 0.03fF
C14407 OR2X1_LOC_677/Y AND2X1_LOC_621/Y 0.03fF
C14408 OR2X1_LOC_317/a_8_216# OR2X1_LOC_160/A 0.02fF
C14409 OR2X1_LOC_160/B OR2X1_LOC_208/a_8_216# 0.02fF
C14410 AND2X1_LOC_810/A AND2X1_LOC_856/a_8_24# 0.01fF
C14411 OR2X1_LOC_56/A AND2X1_LOC_361/A 0.02fF
C14412 AND2X1_LOC_755/a_36_24# OR2X1_LOC_756/B 0.00fF
C14413 OR2X1_LOC_621/B OR2X1_LOC_624/B 0.27fF
C14414 AND2X1_LOC_12/Y AND2X1_LOC_39/a_8_24# 0.01fF
C14415 OR2X1_LOC_691/Y AND2X1_LOC_48/A 0.05fF
C14416 OR2X1_LOC_36/Y AND2X1_LOC_222/a_8_24# 0.01fF
C14417 OR2X1_LOC_810/A OR2X1_LOC_244/Y 0.05fF
C14418 OR2X1_LOC_359/a_36_216# OR2X1_LOC_287/B 0.00fF
C14419 AND2X1_LOC_729/B OR2X1_LOC_13/Y 1.99fF
C14420 OR2X1_LOC_443/Y OR2X1_LOC_161/B 0.01fF
C14421 OR2X1_LOC_744/A OR2X1_LOC_271/Y 0.03fF
C14422 D_INPUT_5 AND2X1_LOC_43/B 0.93fF
C14423 AND2X1_LOC_557/Y AND2X1_LOC_367/A 0.40fF
C14424 VDD OR2X1_LOC_220/a_8_216# 0.00fF
C14425 OR2X1_LOC_702/A AND2X1_LOC_18/Y 0.13fF
C14426 OR2X1_LOC_349/a_36_216# OR2X1_LOC_287/B 0.00fF
C14427 AND2X1_LOC_40/Y AND2X1_LOC_59/Y 1.88fF
C14428 OR2X1_LOC_506/A OR2X1_LOC_737/A 0.02fF
C14429 AND2X1_LOC_732/a_8_24# OR2X1_LOC_89/A 0.01fF
C14430 OR2X1_LOC_139/A OR2X1_LOC_244/A 0.02fF
C14431 OR2X1_LOC_703/A AND2X1_LOC_56/B 0.00fF
C14432 OR2X1_LOC_121/B AND2X1_LOC_607/a_8_24# 0.01fF
C14433 OR2X1_LOC_617/a_8_216# OR2X1_LOC_626/Y 0.01fF
C14434 AND2X1_LOC_48/A OR2X1_LOC_713/A 0.05fF
C14435 OR2X1_LOC_276/a_8_216# OR2X1_LOC_115/B 0.00fF
C14436 OR2X1_LOC_160/A OR2X1_LOC_856/B 0.07fF
C14437 AND2X1_LOC_520/a_8_24# OR2X1_LOC_31/Y 0.01fF
C14438 OR2X1_LOC_825/a_8_216# OR2X1_LOC_600/A 0.01fF
C14439 OR2X1_LOC_40/Y AND2X1_LOC_663/B 0.03fF
C14440 AND2X1_LOC_22/Y AND2X1_LOC_47/Y 0.45fF
C14441 OR2X1_LOC_756/B OR2X1_LOC_269/B 0.05fF
C14442 AND2X1_LOC_95/Y OR2X1_LOC_506/A 0.03fF
C14443 INPUT_3 AND2X1_LOC_62/a_36_24# 0.00fF
C14444 AND2X1_LOC_576/a_8_24# OR2X1_LOC_427/A 0.04fF
C14445 OR2X1_LOC_609/a_8_216# OR2X1_LOC_59/Y 0.02fF
C14446 OR2X1_LOC_166/a_8_216# AND2X1_LOC_390/B 0.03fF
C14447 OR2X1_LOC_864/A OR2X1_LOC_663/A 14.17fF
C14448 AND2X1_LOC_339/Y OR2X1_LOC_31/Y 0.08fF
C14449 OR2X1_LOC_5/a_36_216# INPUT_2 0.03fF
C14450 AND2X1_LOC_346/a_8_24# OR2X1_LOC_295/Y 0.01fF
C14451 AND2X1_LOC_3/Y OR2X1_LOC_78/a_8_216# 0.02fF
C14452 OR2X1_LOC_604/A OR2X1_LOC_684/Y 0.02fF
C14453 AND2X1_LOC_675/Y OR2X1_LOC_74/A 0.93fF
C14454 OR2X1_LOC_316/Y OR2X1_LOC_619/Y 0.03fF
C14455 OR2X1_LOC_18/Y AND2X1_LOC_858/a_36_24# 0.00fF
C14456 OR2X1_LOC_368/A AND2X1_LOC_457/a_8_24# 0.17fF
C14457 AND2X1_LOC_99/A AND2X1_LOC_572/A 0.01fF
C14458 OR2X1_LOC_476/B AND2X1_LOC_18/Y 0.08fF
C14459 OR2X1_LOC_616/Y AND2X1_LOC_621/Y 0.14fF
C14460 AND2X1_LOC_47/Y AND2X1_LOC_417/a_36_24# 0.01fF
C14461 AND2X1_LOC_59/Y OR2X1_LOC_537/A 0.01fF
C14462 AND2X1_LOC_12/Y AND2X1_LOC_43/B 0.41fF
C14463 OR2X1_LOC_715/B OR2X1_LOC_814/A 0.10fF
C14464 OR2X1_LOC_85/A OR2X1_LOC_278/Y 0.02fF
C14465 OR2X1_LOC_321/Y OR2X1_LOC_91/A 0.00fF
C14466 AND2X1_LOC_51/Y OR2X1_LOC_35/Y 0.04fF
C14467 OR2X1_LOC_648/B OR2X1_LOC_648/a_8_216# 0.01fF
C14468 OR2X1_LOC_85/A OR2X1_LOC_38/a_8_216# 0.00fF
C14469 AND2X1_LOC_354/B OR2X1_LOC_619/Y 0.07fF
C14470 OR2X1_LOC_404/Y OR2X1_LOC_573/a_8_216# 0.05fF
C14471 AND2X1_LOC_3/Y OR2X1_LOC_475/B 0.03fF
C14472 AND2X1_LOC_59/Y OR2X1_LOC_87/Y 0.03fF
C14473 INPUT_0 OR2X1_LOC_275/a_8_216# 0.02fF
C14474 AND2X1_LOC_339/B AND2X1_LOC_476/A 0.14fF
C14475 OR2X1_LOC_604/A AND2X1_LOC_845/Y 0.10fF
C14476 OR2X1_LOC_695/a_8_216# OR2X1_LOC_7/A 0.04fF
C14477 OR2X1_LOC_15/a_8_216# D_INPUT_1 0.01fF
C14478 AND2X1_LOC_729/Y OR2X1_LOC_36/Y 0.04fF
C14479 OR2X1_LOC_377/A AND2X1_LOC_472/B 6.12fF
C14480 AND2X1_LOC_217/Y AND2X1_LOC_656/Y 3.33fF
C14481 OR2X1_LOC_235/B OR2X1_LOC_291/Y 0.00fF
C14482 AND2X1_LOC_7/B OR2X1_LOC_493/Y 0.10fF
C14483 AND2X1_LOC_7/B OR2X1_LOC_801/B 0.07fF
C14484 OR2X1_LOC_485/A AND2X1_LOC_841/B 0.03fF
C14485 AND2X1_LOC_36/Y AND2X1_LOC_268/a_8_24# 0.01fF
C14486 AND2X1_LOC_335/Y AND2X1_LOC_863/Y 0.01fF
C14487 AND2X1_LOC_580/B OR2X1_LOC_680/A 0.03fF
C14488 AND2X1_LOC_824/B AND2X1_LOC_472/B 0.01fF
C14489 OR2X1_LOC_620/B OR2X1_LOC_220/B 0.01fF
C14490 OR2X1_LOC_426/B OR2X1_LOC_71/Y 0.08fF
C14491 OR2X1_LOC_462/B OR2X1_LOC_642/a_36_216# 0.03fF
C14492 OR2X1_LOC_520/Y OR2X1_LOC_649/B 0.01fF
C14493 AND2X1_LOC_22/Y OR2X1_LOC_598/A 0.11fF
C14494 AND2X1_LOC_392/A AND2X1_LOC_866/A 0.07fF
C14495 OR2X1_LOC_3/Y AND2X1_LOC_99/A 0.12fF
C14496 OR2X1_LOC_865/a_8_216# OR2X1_LOC_859/B 0.04fF
C14497 OR2X1_LOC_7/A AND2X1_LOC_474/a_8_24# 0.01fF
C14498 OR2X1_LOC_483/a_8_216# OR2X1_LOC_631/B 0.03fF
C14499 OR2X1_LOC_732/A OR2X1_LOC_308/Y 0.02fF
C14500 OR2X1_LOC_185/Y OR2X1_LOC_809/a_8_216# 0.04fF
C14501 OR2X1_LOC_325/A OR2X1_LOC_121/B 0.01fF
C14502 OR2X1_LOC_562/Y OR2X1_LOC_562/A 0.14fF
C14503 OR2X1_LOC_251/Y AND2X1_LOC_668/a_8_24# 0.01fF
C14504 AND2X1_LOC_784/A OR2X1_LOC_36/Y 0.07fF
C14505 AND2X1_LOC_390/B OR2X1_LOC_619/Y 0.07fF
C14506 AND2X1_LOC_784/A OR2X1_LOC_91/a_8_216# 0.03fF
C14507 OR2X1_LOC_600/Y OR2X1_LOC_95/Y 0.02fF
C14508 AND2X1_LOC_356/a_8_24# AND2X1_LOC_390/B 0.01fF
C14509 AND2X1_LOC_302/a_8_24# OR2X1_LOC_7/A 0.02fF
C14510 OR2X1_LOC_221/A OR2X1_LOC_739/B 0.90fF
C14511 OR2X1_LOC_76/Y OR2X1_LOC_269/B 0.44fF
C14512 OR2X1_LOC_793/A OR2X1_LOC_155/A 0.07fF
C14513 OR2X1_LOC_271/B OR2X1_LOC_7/A 0.01fF
C14514 AND2X1_LOC_621/Y AND2X1_LOC_624/a_8_24# 0.20fF
C14515 AND2X1_LOC_167/a_8_24# OR2X1_LOC_532/B 0.01fF
C14516 OR2X1_LOC_124/Y OR2X1_LOC_217/a_8_216# 0.05fF
C14517 OR2X1_LOC_64/Y OR2X1_LOC_71/a_8_216# 0.05fF
C14518 OR2X1_LOC_275/A OR2X1_LOC_39/A 0.04fF
C14519 AND2X1_LOC_59/Y OR2X1_LOC_475/Y 0.00fF
C14520 OR2X1_LOC_276/B AND2X1_LOC_92/Y 0.02fF
C14521 OR2X1_LOC_70/Y OR2X1_LOC_314/Y 0.01fF
C14522 AND2X1_LOC_264/a_36_24# OR2X1_LOC_52/B 0.01fF
C14523 AND2X1_LOC_412/a_8_24# OR2X1_LOC_240/A 0.05fF
C14524 OR2X1_LOC_244/A OR2X1_LOC_244/a_8_216# 0.06fF
C14525 AND2X1_LOC_359/a_8_24# OR2X1_LOC_7/A 0.01fF
C14526 AND2X1_LOC_228/Y OR2X1_LOC_230/a_8_216# 0.01fF
C14527 OR2X1_LOC_22/Y OR2X1_LOC_40/a_8_216# 0.40fF
C14528 D_INPUT_0 OR2X1_LOC_623/B 0.03fF
C14529 OR2X1_LOC_426/B D_INPUT_1 0.21fF
C14530 OR2X1_LOC_44/Y AND2X1_LOC_211/a_8_24# 0.04fF
C14531 AND2X1_LOC_17/Y AND2X1_LOC_21/Y 0.09fF
C14532 OR2X1_LOC_154/A AND2X1_LOC_67/Y 0.03fF
C14533 OR2X1_LOC_235/B D_INPUT_3 0.01fF
C14534 AND2X1_LOC_640/Y OR2X1_LOC_26/Y 0.01fF
C14535 OR2X1_LOC_377/A OR2X1_LOC_19/B 0.32fF
C14536 AND2X1_LOC_443/a_8_24# AND2X1_LOC_222/Y 0.01fF
C14537 OR2X1_LOC_780/B AND2X1_LOC_424/a_8_24# 0.04fF
C14538 OR2X1_LOC_91/A AND2X1_LOC_687/a_8_24# 0.01fF
C14539 OR2X1_LOC_22/Y OR2X1_LOC_118/Y 0.03fF
C14540 OR2X1_LOC_92/Y OR2X1_LOC_31/Y 0.06fF
C14541 OR2X1_LOC_19/B AND2X1_LOC_824/B 1.76fF
C14542 OR2X1_LOC_404/Y OR2X1_LOC_659/B 0.02fF
C14543 AND2X1_LOC_795/Y OR2X1_LOC_56/A 0.13fF
C14544 AND2X1_LOC_717/B OR2X1_LOC_371/Y 0.01fF
C14545 OR2X1_LOC_185/A AND2X1_LOC_69/a_8_24# 0.00fF
C14546 OR2X1_LOC_311/Y AND2X1_LOC_319/A 0.16fF
C14547 OR2X1_LOC_207/B OR2X1_LOC_193/a_8_216# 0.05fF
C14548 OR2X1_LOC_680/Y AND2X1_LOC_147/Y 0.01fF
C14549 AND2X1_LOC_75/a_8_24# OR2X1_LOC_76/Y 0.01fF
C14550 OR2X1_LOC_176/Y OR2X1_LOC_437/A 0.02fF
C14551 AND2X1_LOC_657/Y OR2X1_LOC_406/A 0.14fF
C14552 OR2X1_LOC_476/B AND2X1_LOC_413/a_8_24# 0.23fF
C14553 OR2X1_LOC_19/B OR2X1_LOC_85/A 0.04fF
C14554 AND2X1_LOC_91/B OR2X1_LOC_771/B 0.03fF
C14555 OR2X1_LOC_78/B OR2X1_LOC_194/a_36_216# 0.01fF
C14556 OR2X1_LOC_336/a_8_216# OR2X1_LOC_303/B 0.01fF
C14557 OR2X1_LOC_95/Y OR2X1_LOC_531/a_8_216# 0.01fF
C14558 OR2X1_LOC_54/Y OR2X1_LOC_6/A 0.48fF
C14559 AND2X1_LOC_863/Y OR2X1_LOC_619/Y 0.04fF
C14560 OR2X1_LOC_782/B OR2X1_LOC_781/Y 0.45fF
C14561 OR2X1_LOC_52/Y OR2X1_LOC_52/B 0.01fF
C14562 OR2X1_LOC_391/a_8_216# D_INPUT_1 0.01fF
C14563 OR2X1_LOC_87/A OR2X1_LOC_781/Y 0.11fF
C14564 OR2X1_LOC_472/B OR2X1_LOC_461/A 0.15fF
C14565 AND2X1_LOC_154/Y AND2X1_LOC_156/a_8_24# 0.03fF
C14566 AND2X1_LOC_228/Y D_INPUT_0 0.02fF
C14567 OR2X1_LOC_272/Y OR2X1_LOC_79/A 0.19fF
C14568 OR2X1_LOC_26/Y OR2X1_LOC_416/Y 0.04fF
C14569 OR2X1_LOC_256/a_36_216# OR2X1_LOC_95/Y 0.01fF
C14570 AND2X1_LOC_348/A OR2X1_LOC_47/Y 0.01fF
C14571 AND2X1_LOC_663/B OR2X1_LOC_7/A 0.07fF
C14572 OR2X1_LOC_70/Y OR2X1_LOC_131/Y 0.04fF
C14573 OR2X1_LOC_46/A OR2X1_LOC_69/Y 0.00fF
C14574 AND2X1_LOC_212/Y OR2X1_LOC_437/A 0.07fF
C14575 AND2X1_LOC_64/Y OR2X1_LOC_319/Y 0.58fF
C14576 AND2X1_LOC_212/A AND2X1_LOC_212/a_8_24# 0.09fF
C14577 AND2X1_LOC_91/B OR2X1_LOC_776/A 0.10fF
C14578 OR2X1_LOC_244/B OR2X1_LOC_598/A 0.02fF
C14579 AND2X1_LOC_153/a_8_24# AND2X1_LOC_47/Y 0.03fF
C14580 OR2X1_LOC_487/Y OR2X1_LOC_488/Y 0.08fF
C14581 OR2X1_LOC_737/A D_INPUT_1 0.04fF
C14582 OR2X1_LOC_427/A AND2X1_LOC_452/a_36_24# 0.00fF
C14583 OR2X1_LOC_479/Y OR2X1_LOC_76/A 0.02fF
C14584 AND2X1_LOC_95/Y AND2X1_LOC_420/a_8_24# 0.03fF
C14585 OR2X1_LOC_158/A OR2X1_LOC_13/B 1.19fF
C14586 AND2X1_LOC_839/A OR2X1_LOC_824/Y 0.03fF
C14587 AND2X1_LOC_7/B OR2X1_LOC_130/a_8_216# 0.05fF
C14588 OR2X1_LOC_59/Y AND2X1_LOC_657/A 0.07fF
C14589 AND2X1_LOC_95/Y D_INPUT_1 0.03fF
C14590 OR2X1_LOC_855/a_8_216# AND2X1_LOC_36/Y 0.01fF
C14591 D_INPUT_7 AND2X1_LOC_11/a_8_24# 0.01fF
C14592 OR2X1_LOC_377/A OR2X1_LOC_838/B 0.01fF
C14593 D_INPUT_0 OR2X1_LOC_585/A 0.11fF
C14594 VDD OR2X1_LOC_71/A 1.12fF
C14595 OR2X1_LOC_633/Y D_INPUT_1 0.03fF
C14596 OR2X1_LOC_2/Y OR2X1_LOC_581/a_8_216# 0.01fF
C14597 OR2X1_LOC_85/A OR2X1_LOC_75/Y 0.00fF
C14598 AND2X1_LOC_363/Y OR2X1_LOC_384/Y 0.01fF
C14599 AND2X1_LOC_726/Y AND2X1_LOC_731/a_8_24# 0.18fF
C14600 OR2X1_LOC_461/Y OR2X1_LOC_416/Y 0.00fF
C14601 AND2X1_LOC_46/a_8_24# OR2X1_LOC_121/B 0.01fF
C14602 OR2X1_LOC_62/A OR2X1_LOC_36/Y 0.00fF
C14603 AND2X1_LOC_621/Y AND2X1_LOC_624/B 0.03fF
C14604 OR2X1_LOC_185/A OR2X1_LOC_804/A 0.19fF
C14605 OR2X1_LOC_524/Y OR2X1_LOC_152/a_8_216# 0.15fF
C14606 OR2X1_LOC_53/Y OR2X1_LOC_56/a_8_216# 0.07fF
C14607 OR2X1_LOC_204/Y OR2X1_LOC_786/Y 0.00fF
C14608 OR2X1_LOC_161/B OR2X1_LOC_605/Y 0.02fF
C14609 OR2X1_LOC_630/a_8_216# OR2X1_LOC_598/A 0.03fF
C14610 AND2X1_LOC_366/a_8_24# OR2X1_LOC_437/A 0.02fF
C14611 OR2X1_LOC_420/a_36_216# OR2X1_LOC_95/Y 0.03fF
C14612 OR2X1_LOC_375/A OR2X1_LOC_66/a_8_216# 0.01fF
C14613 AND2X1_LOC_260/a_36_24# OR2X1_LOC_46/A 0.00fF
C14614 AND2X1_LOC_307/Y AND2X1_LOC_727/A 0.01fF
C14615 OR2X1_LOC_22/Y AND2X1_LOC_855/a_8_24# 0.01fF
C14616 AND2X1_LOC_196/a_36_24# AND2X1_LOC_196/Y 0.00fF
C14617 AND2X1_LOC_729/Y OR2X1_LOC_419/Y 0.48fF
C14618 OR2X1_LOC_805/A OR2X1_LOC_493/Y 0.05fF
C14619 OR2X1_LOC_805/A OR2X1_LOC_801/B 0.02fF
C14620 AND2X1_LOC_64/Y OR2X1_LOC_691/A 0.00fF
C14621 OR2X1_LOC_356/B OR2X1_LOC_356/A 0.78fF
C14622 AND2X1_LOC_537/Y OR2X1_LOC_46/A 0.00fF
C14623 AND2X1_LOC_539/Y AND2X1_LOC_810/B 0.26fF
C14624 OR2X1_LOC_440/a_36_216# OR2X1_LOC_180/B 0.00fF
C14625 OR2X1_LOC_111/a_8_216# OR2X1_LOC_158/A 0.03fF
C14626 AND2X1_LOC_22/Y AND2X1_LOC_263/a_36_24# 0.01fF
C14627 OR2X1_LOC_625/Y AND2X1_LOC_793/B -0.02fF
C14628 AND2X1_LOC_633/Y AND2X1_LOC_634/Y 0.19fF
C14629 AND2X1_LOC_98/Y OR2X1_LOC_13/B 0.02fF
C14630 OR2X1_LOC_417/Y OR2X1_LOC_604/a_8_216# 0.01fF
C14631 OR2X1_LOC_45/B OR2X1_LOC_428/A 0.20fF
C14632 AND2X1_LOC_784/A OR2X1_LOC_419/Y 0.10fF
C14633 OR2X1_LOC_417/Y AND2X1_LOC_170/B 0.31fF
C14634 OR2X1_LOC_246/A OR2X1_LOC_71/Y 0.02fF
C14635 OR2X1_LOC_3/B OR2X1_LOC_47/a_8_216# 0.05fF
C14636 OR2X1_LOC_70/A OR2X1_LOC_25/a_8_216# 0.01fF
C14637 AND2X1_LOC_640/a_8_24# INPUT_1 0.01fF
C14638 OR2X1_LOC_219/a_8_216# OR2X1_LOC_228/Y 0.01fF
C14639 AND2X1_LOC_150/a_8_24# OR2X1_LOC_267/Y 0.01fF
C14640 OR2X1_LOC_348/Y OR2X1_LOC_363/a_8_216# 0.02fF
C14641 AND2X1_LOC_703/Y OR2X1_LOC_16/A 0.01fF
C14642 OR2X1_LOC_56/A AND2X1_LOC_439/a_8_24# 0.04fF
C14643 OR2X1_LOC_45/B OR2X1_LOC_595/A 0.03fF
C14644 AND2X1_LOC_521/a_8_24# AND2X1_LOC_22/Y 0.03fF
C14645 AND2X1_LOC_729/Y OR2X1_LOC_526/a_8_216# 0.01fF
C14646 AND2X1_LOC_217/Y AND2X1_LOC_772/Y 0.02fF
C14647 OR2X1_LOC_154/A OR2X1_LOC_715/a_36_216# 0.01fF
C14648 OR2X1_LOC_296/a_8_216# OR2X1_LOC_598/A -0.02fF
C14649 OR2X1_LOC_135/Y OR2X1_LOC_12/Y 0.48fF
C14650 AND2X1_LOC_42/B AND2X1_LOC_72/B 0.03fF
C14651 OR2X1_LOC_288/A OR2X1_LOC_286/B 0.02fF
C14652 OR2X1_LOC_482/Y AND2X1_LOC_242/a_8_24# 0.04fF
C14653 OR2X1_LOC_36/Y OR2X1_LOC_172/Y 0.04fF
C14654 AND2X1_LOC_12/Y OR2X1_LOC_558/A 0.33fF
C14655 OR2X1_LOC_333/B OR2X1_LOC_351/a_36_216# 0.00fF
C14656 OR2X1_LOC_361/a_8_216# OR2X1_LOC_161/B 0.02fF
C14657 OR2X1_LOC_40/Y OR2X1_LOC_18/a_8_216# 0.01fF
C14658 INPUT_1 AND2X1_LOC_649/Y 0.01fF
C14659 AND2X1_LOC_719/Y AND2X1_LOC_786/Y 0.10fF
C14660 AND2X1_LOC_706/Y OR2X1_LOC_589/A 0.11fF
C14661 OR2X1_LOC_486/Y OR2X1_LOC_549/A 0.07fF
C14662 OR2X1_LOC_26/Y OR2X1_LOC_80/A 0.72fF
C14663 OR2X1_LOC_654/A AND2X1_LOC_31/Y 8.99fF
C14664 OR2X1_LOC_287/B OR2X1_LOC_68/B 0.04fF
C14665 OR2X1_LOC_45/B AND2X1_LOC_215/Y 0.45fF
C14666 OR2X1_LOC_41/Y OR2X1_LOC_43/a_8_216# 0.42fF
C14667 OR2X1_LOC_70/Y OR2X1_LOC_331/a_36_216# 0.00fF
C14668 AND2X1_LOC_721/Y OR2X1_LOC_666/A 0.02fF
C14669 AND2X1_LOC_227/Y AND2X1_LOC_137/a_8_24# 0.01fF
C14670 OR2X1_LOC_160/B OR2X1_LOC_138/A 0.06fF
C14671 OR2X1_LOC_599/A OR2X1_LOC_589/Y 0.00fF
C14672 AND2X1_LOC_474/A OR2X1_LOC_89/Y 0.01fF
C14673 AND2X1_LOC_64/Y OR2X1_LOC_294/a_8_216# 0.01fF
C14674 OR2X1_LOC_492/a_8_216# OR2X1_LOC_108/Y 0.06fF
C14675 OR2X1_LOC_39/A OR2X1_LOC_142/Y 0.02fF
C14676 AND2X1_LOC_851/B AND2X1_LOC_318/Y 0.23fF
C14677 AND2X1_LOC_3/Y OR2X1_LOC_193/a_8_216# 0.04fF
C14678 AND2X1_LOC_564/B OR2X1_LOC_164/Y 0.01fF
C14679 OR2X1_LOC_417/Y OR2X1_LOC_331/Y 0.07fF
C14680 AND2X1_LOC_262/a_8_24# AND2X1_LOC_18/Y 0.03fF
C14681 OR2X1_LOC_118/a_36_216# OR2X1_LOC_744/A 0.00fF
C14682 OR2X1_LOC_659/A OR2X1_LOC_474/B 0.00fF
C14683 INPUT_5 AND2X1_LOC_588/B 0.01fF
C14684 OR2X1_LOC_292/a_8_216# OR2X1_LOC_428/A 0.02fF
C14685 OR2X1_LOC_375/A OR2X1_LOC_308/Y 0.01fF
C14686 OR2X1_LOC_692/Y OR2X1_LOC_744/A 0.01fF
C14687 OR2X1_LOC_709/A AND2X1_LOC_92/Y 0.07fF
C14688 AND2X1_LOC_64/Y OR2X1_LOC_811/A 0.03fF
C14689 AND2X1_LOC_392/A OR2X1_LOC_40/Y 0.10fF
C14690 OR2X1_LOC_829/A AND2X1_LOC_434/Y 0.10fF
C14691 OR2X1_LOC_200/Y OR2X1_LOC_207/a_8_216# 0.39fF
C14692 AND2X1_LOC_22/Y OR2X1_LOC_828/a_8_216# 0.03fF
C14693 OR2X1_LOC_40/Y AND2X1_LOC_807/B 0.01fF
C14694 OR2X1_LOC_696/A OR2X1_LOC_127/Y 0.22fF
C14695 AND2X1_LOC_794/B OR2X1_LOC_59/Y 0.10fF
C14696 D_INPUT_3 AND2X1_LOC_721/A 0.04fF
C14697 AND2X1_LOC_339/B INPUT_0 0.14fF
C14698 OR2X1_LOC_61/B AND2X1_LOC_7/B 0.01fF
C14699 AND2X1_LOC_43/B OR2X1_LOC_356/B 0.02fF
C14700 OR2X1_LOC_97/A OR2X1_LOC_775/a_8_216# 0.03fF
C14701 OR2X1_LOC_9/Y OR2X1_LOC_56/A 0.07fF
C14702 OR2X1_LOC_538/a_8_216# OR2X1_LOC_161/B 0.01fF
C14703 OR2X1_LOC_778/Y OR2X1_LOC_593/B 0.03fF
C14704 OR2X1_LOC_516/Y AND2X1_LOC_576/Y 0.02fF
C14705 OR2X1_LOC_161/A OR2X1_LOC_115/B 0.12fF
C14706 AND2X1_LOC_392/A AND2X1_LOC_535/a_8_24# 0.20fF
C14707 OR2X1_LOC_715/B OR2X1_LOC_715/A 0.21fF
C14708 AND2X1_LOC_91/B OR2X1_LOC_402/Y 0.46fF
C14709 OR2X1_LOC_35/a_8_216# OR2X1_LOC_66/A 0.14fF
C14710 OR2X1_LOC_338/a_8_216# OR2X1_LOC_756/B 0.01fF
C14711 OR2X1_LOC_194/B AND2X1_LOC_7/B 0.05fF
C14712 OR2X1_LOC_427/A OR2X1_LOC_816/A 2.22fF
C14713 AND2X1_LOC_357/B OR2X1_LOC_91/A 0.00fF
C14714 OR2X1_LOC_858/A VDD 1.33fF
C14715 AND2X1_LOC_22/Y OR2X1_LOC_506/A 0.02fF
C14716 OR2X1_LOC_744/A OR2X1_LOC_600/A 6.00fF
C14717 OR2X1_LOC_696/A AND2X1_LOC_836/a_8_24# 0.01fF
C14718 VDD OR2X1_LOC_59/Y 1.25fF
C14719 OR2X1_LOC_185/Y AND2X1_LOC_760/a_8_24# 0.24fF
C14720 D_GATE_662 OR2X1_LOC_772/B 0.02fF
C14721 OR2X1_LOC_828/B AND2X1_LOC_829/a_8_24# 0.01fF
C14722 OR2X1_LOC_456/a_8_216# OR2X1_LOC_577/Y 0.01fF
C14723 AND2X1_LOC_42/B AND2X1_LOC_36/Y 0.16fF
C14724 OR2X1_LOC_739/A OR2X1_LOC_355/A 0.01fF
C14725 AND2X1_LOC_70/Y AND2X1_LOC_92/Y 0.07fF
C14726 OR2X1_LOC_48/B AND2X1_LOC_771/a_36_24# 0.01fF
C14727 OR2X1_LOC_524/Y OR2X1_LOC_745/a_36_216# 0.16fF
C14728 AND2X1_LOC_363/Y OR2X1_LOC_91/A 0.09fF
C14729 OR2X1_LOC_196/B OR2X1_LOC_515/a_8_216# 0.01fF
C14730 AND2X1_LOC_291/a_8_24# AND2X1_LOC_7/B 0.01fF
C14731 OR2X1_LOC_121/B OR2X1_LOC_544/B 0.27fF
C14732 OR2X1_LOC_134/Y AND2X1_LOC_560/B 0.15fF
C14733 OR2X1_LOC_18/Y AND2X1_LOC_771/a_36_24# 0.00fF
C14734 AND2X1_LOC_707/a_36_24# OR2X1_LOC_91/A 0.00fF
C14735 OR2X1_LOC_185/Y OR2X1_LOC_121/A 0.13fF
C14736 AND2X1_LOC_175/B OR2X1_LOC_12/Y 0.01fF
C14737 OR2X1_LOC_831/A OR2X1_LOC_794/A 0.16fF
C14738 OR2X1_LOC_255/a_8_216# OR2X1_LOC_437/A 0.03fF
C14739 OR2X1_LOC_36/Y AND2X1_LOC_206/a_8_24# 0.01fF
C14740 OR2X1_LOC_147/B OR2X1_LOC_543/A 0.05fF
C14741 AND2X1_LOC_90/a_8_24# OR2X1_LOC_375/A 0.01fF
C14742 AND2X1_LOC_700/a_8_24# OR2X1_LOC_502/A 0.00fF
C14743 OR2X1_LOC_62/B OR2X1_LOC_217/A 0.01fF
C14744 OR2X1_LOC_703/A AND2X1_LOC_92/Y 0.03fF
C14745 OR2X1_LOC_441/Y AND2X1_LOC_658/Y 0.02fF
C14746 OR2X1_LOC_136/a_8_216# AND2X1_LOC_211/B 0.03fF
C14747 OR2X1_LOC_767/a_8_216# OR2X1_LOC_595/A 0.01fF
C14748 OR2X1_LOC_121/Y OR2X1_LOC_510/Y 0.24fF
C14749 OR2X1_LOC_184/Y AND2X1_LOC_657/A 0.03fF
C14750 OR2X1_LOC_621/B OR2X1_LOC_847/A 0.01fF
C14751 AND2X1_LOC_59/Y OR2X1_LOC_356/A 0.21fF
C14752 OR2X1_LOC_624/a_8_216# OR2X1_LOC_624/Y 0.01fF
C14753 OR2X1_LOC_319/a_8_216# AND2X1_LOC_110/Y 0.01fF
C14754 OR2X1_LOC_9/Y AND2X1_LOC_9/a_8_24# 0.01fF
C14755 OR2X1_LOC_175/Y AND2X1_LOC_3/Y 0.03fF
C14756 AND2X1_LOC_712/Y AND2X1_LOC_448/Y 0.01fF
C14757 AND2X1_LOC_723/a_8_24# OR2X1_LOC_51/Y 0.01fF
C14758 AND2X1_LOC_367/A AND2X1_LOC_456/B 0.01fF
C14759 OR2X1_LOC_20/Y OR2X1_LOC_18/Y 0.02fF
C14760 OR2X1_LOC_377/A OR2X1_LOC_621/a_36_216# 0.01fF
C14761 AND2X1_LOC_12/Y AND2X1_LOC_625/a_36_24# 0.00fF
C14762 OR2X1_LOC_51/Y OR2X1_LOC_278/Y 2.61fF
C14763 AND2X1_LOC_51/Y OR2X1_LOC_115/B 0.03fF
C14764 OR2X1_LOC_177/Y AND2X1_LOC_784/A 0.02fF
C14765 AND2X1_LOC_566/B AND2X1_LOC_303/B 0.14fF
C14766 AND2X1_LOC_729/Y OR2X1_LOC_604/A 0.07fF
C14767 OR2X1_LOC_691/Y AND2X1_LOC_3/Y 0.05fF
C14768 AND2X1_LOC_476/A OR2X1_LOC_300/Y 0.01fF
C14769 OR2X1_LOC_348/Y AND2X1_LOC_12/Y 0.29fF
C14770 AND2X1_LOC_734/Y OR2X1_LOC_441/Y 0.17fF
C14771 OR2X1_LOC_156/A OR2X1_LOC_154/A 0.14fF
C14772 AND2X1_LOC_736/Y AND2X1_LOC_736/a_8_24# 0.01fF
C14773 OR2X1_LOC_494/Y AND2X1_LOC_573/A 0.02fF
C14774 OR2X1_LOC_95/Y OR2X1_LOC_749/Y 0.01fF
C14775 OR2X1_LOC_121/Y OR2X1_LOC_810/A 0.10fF
C14776 AND2X1_LOC_741/Y AND2X1_LOC_223/A 0.00fF
C14777 AND2X1_LOC_12/Y OR2X1_LOC_349/a_8_216# 0.01fF
C14778 AND2X1_LOC_592/Y OR2X1_LOC_44/Y 0.05fF
C14779 OR2X1_LOC_448/Y OR2X1_LOC_66/A 0.01fF
C14780 VDD OR2X1_LOC_169/B 0.00fF
C14781 OR2X1_LOC_411/Y OR2X1_LOC_413/a_8_216# 0.40fF
C14782 OR2X1_LOC_67/Y OR2X1_LOC_71/A 0.03fF
C14783 OR2X1_LOC_605/B AND2X1_LOC_604/a_8_24# 0.02fF
C14784 AND2X1_LOC_3/Y OR2X1_LOC_713/A 0.01fF
C14785 AND2X1_LOC_111/a_8_24# OR2X1_LOC_161/B 0.01fF
C14786 OR2X1_LOC_744/A OR2X1_LOC_619/Y 0.13fF
C14787 OR2X1_LOC_600/A AND2X1_LOC_840/B 0.05fF
C14788 OR2X1_LOC_602/a_8_216# OR2X1_LOC_161/B 0.03fF
C14789 OR2X1_LOC_65/Y AND2X1_LOC_201/Y 0.80fF
C14790 AND2X1_LOC_784/A OR2X1_LOC_604/A 0.10fF
C14791 AND2X1_LOC_259/Y AND2X1_LOC_346/a_8_24# 0.20fF
C14792 AND2X1_LOC_748/a_36_24# OR2X1_LOC_78/B 0.01fF
C14793 OR2X1_LOC_589/A OR2X1_LOC_485/A 0.18fF
C14794 VDD OR2X1_LOC_433/a_8_216# 0.00fF
C14795 AND2X1_LOC_580/A AND2X1_LOC_658/A 11.83fF
C14796 OR2X1_LOC_811/A OR2X1_LOC_464/A 0.12fF
C14797 OR2X1_LOC_8/Y OR2X1_LOC_36/Y 0.04fF
C14798 OR2X1_LOC_114/B AND2X1_LOC_159/a_8_24# 0.01fF
C14799 OR2X1_LOC_74/A AND2X1_LOC_443/a_8_24# 0.03fF
C14800 OR2X1_LOC_577/a_8_216# D_GATE_366 0.01fF
C14801 VDD OR2X1_LOC_820/B 0.11fF
C14802 AND2X1_LOC_521/a_36_24# AND2X1_LOC_42/B 0.01fF
C14803 OR2X1_LOC_96/B OR2X1_LOC_56/A 0.04fF
C14804 AND2X1_LOC_191/Y AND2X1_LOC_479/a_8_24# 0.05fF
C14805 AND2X1_LOC_840/a_8_24# AND2X1_LOC_833/a_8_24# 0.23fF
C14806 AND2X1_LOC_851/A OR2X1_LOC_495/Y 0.01fF
C14807 AND2X1_LOC_468/B OR2X1_LOC_594/a_8_216# 0.03fF
C14808 OR2X1_LOC_6/B AND2X1_LOC_490/a_8_24# 0.11fF
C14809 OR2X1_LOC_687/Y OR2X1_LOC_78/A 0.03fF
C14810 OR2X1_LOC_744/A OR2X1_LOC_88/A 0.00fF
C14811 AND2X1_LOC_794/B OR2X1_LOC_70/Y 0.08fF
C14812 AND2X1_LOC_711/Y AND2X1_LOC_220/a_36_24# 0.01fF
C14813 AND2X1_LOC_481/a_8_24# AND2X1_LOC_18/Y 0.14fF
C14814 AND2X1_LOC_366/a_8_24# OR2X1_LOC_753/A 0.03fF
C14815 AND2X1_LOC_392/A OR2X1_LOC_7/A 0.07fF
C14816 OR2X1_LOC_22/Y AND2X1_LOC_208/Y 0.00fF
C14817 AND2X1_LOC_122/a_36_24# OR2X1_LOC_549/A 0.01fF
C14818 OR2X1_LOC_494/Y OR2X1_LOC_669/Y 0.07fF
C14819 OR2X1_LOC_9/Y OR2X1_LOC_291/A 0.00fF
C14820 OR2X1_LOC_216/A OR2X1_LOC_624/A 0.33fF
C14821 AND2X1_LOC_719/Y AND2X1_LOC_578/A 0.10fF
C14822 AND2X1_LOC_348/A OR2X1_LOC_625/Y 0.02fF
C14823 OR2X1_LOC_840/A OR2X1_LOC_161/A 0.10fF
C14824 OR2X1_LOC_70/Y AND2X1_LOC_479/a_8_24# 0.02fF
C14825 OR2X1_LOC_807/Y OR2X1_LOC_811/A 0.04fF
C14826 OR2X1_LOC_757/A AND2X1_LOC_580/B 0.03fF
C14827 OR2X1_LOC_491/Y OR2X1_LOC_59/Y 0.03fF
C14828 AND2X1_LOC_554/a_8_24# OR2X1_LOC_71/Y 0.01fF
C14829 AND2X1_LOC_191/Y VDD 0.69fF
C14830 OR2X1_LOC_40/Y OR2X1_LOC_3/a_36_216# 0.00fF
C14831 AND2X1_LOC_752/a_8_24# AND2X1_LOC_43/B 0.04fF
C14832 OR2X1_LOC_160/B OR2X1_LOC_479/Y 0.10fF
C14833 OR2X1_LOC_251/Y OR2X1_LOC_59/Y 0.03fF
C14834 AND2X1_LOC_694/a_8_24# OR2X1_LOC_161/B 0.10fF
C14835 OR2X1_LOC_653/A OR2X1_LOC_435/a_8_216# 0.39fF
C14836 AND2X1_LOC_576/Y AND2X1_LOC_842/a_8_24# 0.01fF
C14837 OR2X1_LOC_279/Y AND2X1_LOC_860/A 0.31fF
C14838 AND2X1_LOC_512/Y OR2X1_LOC_44/Y 0.07fF
C14839 VDD AND2X1_LOC_711/Y 0.92fF
C14840 AND2X1_LOC_794/B AND2X1_LOC_514/Y 0.17fF
C14841 OR2X1_LOC_592/A OR2X1_LOC_66/A 0.01fF
C14842 OR2X1_LOC_426/B OR2X1_LOC_743/A 6.55fF
C14843 OR2X1_LOC_422/Y AND2X1_LOC_448/Y 0.80fF
C14844 OR2X1_LOC_676/Y AND2X1_LOC_136/a_8_24# 0.02fF
C14845 AND2X1_LOC_724/a_8_24# OR2X1_LOC_95/Y 0.01fF
C14846 OR2X1_LOC_653/Y OR2X1_LOC_405/Y 0.01fF
C14847 AND2X1_LOC_522/a_8_24# OR2X1_LOC_532/B 0.01fF
C14848 VDD OR2X1_LOC_70/Y 2.03fF
C14849 OR2X1_LOC_358/a_36_216# OR2X1_LOC_502/A 0.00fF
C14850 OR2X1_LOC_47/Y AND2X1_LOC_209/Y 0.14fF
C14851 AND2X1_LOC_138/a_8_24# AND2X1_LOC_649/B 0.20fF
C14852 OR2X1_LOC_467/A OR2X1_LOC_466/a_8_216# 0.01fF
C14853 AND2X1_LOC_807/Y OR2X1_LOC_427/A 0.07fF
C14854 OR2X1_LOC_58/Y OR2X1_LOC_60/a_8_216# 0.01fF
C14855 OR2X1_LOC_239/Y AND2X1_LOC_663/A 0.42fF
C14856 OR2X1_LOC_427/a_8_216# OR2X1_LOC_427/A 0.01fF
C14857 AND2X1_LOC_580/A AND2X1_LOC_631/a_8_24# 0.07fF
C14858 AND2X1_LOC_366/A OR2X1_LOC_7/A 0.01fF
C14859 OR2X1_LOC_834/a_36_216# OR2X1_LOC_269/B 0.00fF
C14860 OR2X1_LOC_791/B OR2X1_LOC_260/a_36_216# 0.00fF
C14861 OR2X1_LOC_544/A AND2X1_LOC_438/a_8_24# 0.09fF
C14862 OR2X1_LOC_185/A OR2X1_LOC_340/Y 0.02fF
C14863 AND2X1_LOC_567/a_8_24# AND2X1_LOC_802/a_8_24# 0.23fF
C14864 OR2X1_LOC_409/B OR2X1_LOC_585/a_8_216# 0.01fF
C14865 OR2X1_LOC_439/a_8_216# OR2X1_LOC_161/B 0.03fF
C14866 OR2X1_LOC_856/A OR2X1_LOC_532/B 0.02fF
C14867 OR2X1_LOC_118/Y OR2X1_LOC_39/A 0.02fF
C14868 AND2X1_LOC_456/Y AND2X1_LOC_456/B 0.00fF
C14869 OR2X1_LOC_428/Y OR2X1_LOC_428/A 0.00fF
C14870 AND2X1_LOC_145/a_8_24# OR2X1_LOC_161/A 0.01fF
C14871 OR2X1_LOC_185/A OR2X1_LOC_130/A 0.23fF
C14872 AND2X1_LOC_339/B OR2X1_LOC_417/A 0.03fF
C14873 VDD AND2X1_LOC_514/Y 0.72fF
C14874 AND2X1_LOC_76/Y OR2X1_LOC_36/Y 0.02fF
C14875 AND2X1_LOC_59/Y AND2X1_LOC_43/B 5.75fF
C14876 AND2X1_LOC_476/A AND2X1_LOC_219/A 0.78fF
C14877 OR2X1_LOC_108/Y AND2X1_LOC_465/Y 0.00fF
C14878 AND2X1_LOC_12/Y OR2X1_LOC_510/Y 0.00fF
C14879 OR2X1_LOC_51/Y OR2X1_LOC_253/a_8_216# 0.01fF
C14880 OR2X1_LOC_816/a_8_216# OR2X1_LOC_64/Y 0.01fF
C14881 OR2X1_LOC_185/Y OR2X1_LOC_560/a_36_216# 0.14fF
C14882 OR2X1_LOC_3/Y OR2X1_LOC_697/Y 0.01fF
C14883 OR2X1_LOC_377/A OR2X1_LOC_835/A 0.02fF
C14884 OR2X1_LOC_369/a_8_216# OR2X1_LOC_22/Y 0.00fF
C14885 OR2X1_LOC_667/a_8_216# OR2X1_LOC_278/Y 0.01fF
C14886 AND2X1_LOC_388/Y OR2X1_LOC_167/Y 0.07fF
C14887 OR2X1_LOC_624/A OR2X1_LOC_802/Y 0.03fF
C14888 D_INPUT_5 AND2X1_LOC_459/a_8_24# 0.02fF
C14889 OR2X1_LOC_427/A OR2X1_LOC_591/a_8_216# 0.02fF
C14890 OR2X1_LOC_756/B AND2X1_LOC_176/a_8_24# 0.13fF
C14891 AND2X1_LOC_707/a_8_24# AND2X1_LOC_687/B 0.01fF
C14892 OR2X1_LOC_485/A AND2X1_LOC_654/B 0.02fF
C14893 OR2X1_LOC_426/B OR2X1_LOC_246/A 0.97fF
C14894 OR2X1_LOC_539/a_8_216# OR2X1_LOC_154/A 0.05fF
C14895 OR2X1_LOC_140/A D_INPUT_0 0.01fF
C14896 AND2X1_LOC_175/B AND2X1_LOC_650/Y 0.15fF
C14897 AND2X1_LOC_334/a_36_24# AND2X1_LOC_476/A 0.00fF
C14898 OR2X1_LOC_823/Y OR2X1_LOC_824/Y 0.04fF
C14899 OR2X1_LOC_485/A OR2X1_LOC_495/Y 0.03fF
C14900 INPUT_0 OR2X1_LOC_415/A 0.01fF
C14901 OR2X1_LOC_629/Y AND2X1_LOC_3/Y 0.16fF
C14902 OR2X1_LOC_465/a_8_216# OR2X1_LOC_553/A 0.04fF
C14903 OR2X1_LOC_19/B OR2X1_LOC_78/B 0.01fF
C14904 OR2X1_LOC_230/a_8_216# AND2X1_LOC_857/Y 0.01fF
C14905 OR2X1_LOC_399/A OR2X1_LOC_585/A 0.01fF
C14906 AND2X1_LOC_605/Y OR2X1_LOC_417/Y 0.13fF
C14907 VDD OR2X1_LOC_504/Y 0.12fF
C14908 AND2X1_LOC_22/Y AND2X1_LOC_48/Y 0.04fF
C14909 OR2X1_LOC_744/A OR2X1_LOC_22/A 0.01fF
C14910 OR2X1_LOC_43/A OR2X1_LOC_94/a_8_216# 0.43fF
C14911 OR2X1_LOC_861/a_8_216# OR2X1_LOC_392/a_8_216# 0.47fF
C14912 AND2X1_LOC_175/B AND2X1_LOC_175/a_8_24# 0.01fF
C14913 OR2X1_LOC_262/Y OR2X1_LOC_39/A 0.00fF
C14914 AND2X1_LOC_12/Y OR2X1_LOC_810/A 0.17fF
C14915 OR2X1_LOC_840/A AND2X1_LOC_51/Y 0.06fF
C14916 OR2X1_LOC_600/A OR2X1_LOC_31/Y 0.50fF
C14917 OR2X1_LOC_666/Y AND2X1_LOC_621/Y 0.03fF
C14918 OR2X1_LOC_160/A OR2X1_LOC_355/B 0.06fF
C14919 OR2X1_LOC_437/A OR2X1_LOC_183/a_8_216# 0.03fF
C14920 AND2X1_LOC_12/Y OR2X1_LOC_864/a_8_216# 0.01fF
C14921 OR2X1_LOC_238/Y OR2X1_LOC_39/A 0.06fF
C14922 GATE_366 OR2X1_LOC_748/A 0.03fF
C14923 OR2X1_LOC_47/Y OR2X1_LOC_583/a_8_216# 0.01fF
C14924 OR2X1_LOC_411/A OR2X1_LOC_411/a_8_216# 0.47fF
C14925 OR2X1_LOC_83/a_8_216# OR2X1_LOC_394/Y 0.01fF
C14926 OR2X1_LOC_26/Y OR2X1_LOC_6/A 0.14fF
C14927 AND2X1_LOC_191/Y OR2X1_LOC_616/Y 0.03fF
C14928 AND2X1_LOC_722/a_8_24# OR2X1_LOC_47/Y 0.03fF
C14929 OR2X1_LOC_72/Y AND2X1_LOC_201/Y 0.12fF
C14930 OR2X1_LOC_621/A D_INPUT_1 0.14fF
C14931 OR2X1_LOC_426/B OR2X1_LOC_409/B 0.03fF
C14932 OR2X1_LOC_66/a_8_216# OR2X1_LOC_549/A 0.06fF
C14933 OR2X1_LOC_687/Y OR2X1_LOC_155/A 0.53fF
C14934 AND2X1_LOC_326/A AND2X1_LOC_364/A 0.06fF
C14935 OR2X1_LOC_36/Y OR2X1_LOC_52/B 7.04fF
C14936 OR2X1_LOC_247/Y OR2X1_LOC_294/Y 0.02fF
C14937 OR2X1_LOC_18/Y AND2X1_LOC_660/Y 0.03fF
C14938 OR2X1_LOC_788/B OR2X1_LOC_180/B 0.03fF
C14939 AND2X1_LOC_554/B AND2X1_LOC_572/A 0.34fF
C14940 AND2X1_LOC_711/Y OR2X1_LOC_616/Y 0.03fF
C14941 OR2X1_LOC_335/Y OR2X1_LOC_544/A 0.02fF
C14942 OR2X1_LOC_601/Y AND2X1_LOC_602/a_8_24# -0.00fF
C14943 AND2X1_LOC_106/a_36_24# OR2X1_LOC_244/Y 0.00fF
C14944 OR2X1_LOC_89/A OR2X1_LOC_6/A 0.78fF
C14945 VDD OR2X1_LOC_184/Y 0.36fF
C14946 INPUT_3 OR2X1_LOC_5/a_8_216# 0.02fF
C14947 OR2X1_LOC_791/B OR2X1_LOC_792/a_8_216# 0.03fF
C14948 AND2X1_LOC_857/Y D_INPUT_0 0.07fF
C14949 OR2X1_LOC_41/Y OR2X1_LOC_13/Y 0.13fF
C14950 OR2X1_LOC_317/a_36_216# OR2X1_LOC_532/B 0.00fF
C14951 OR2X1_LOC_696/A OR2X1_LOC_424/Y 0.01fF
C14952 AND2X1_LOC_543/a_8_24# OR2X1_LOC_31/Y 0.01fF
C14953 OR2X1_LOC_831/a_36_216# OR2X1_LOC_479/Y 0.01fF
C14954 OR2X1_LOC_485/A OR2X1_LOC_43/A 0.53fF
C14955 AND2X1_LOC_145/a_8_24# AND2X1_LOC_51/Y 0.16fF
C14956 VDD OR2X1_LOC_437/Y 0.12fF
C14957 AND2X1_LOC_364/Y AND2X1_LOC_318/Y 0.02fF
C14958 OR2X1_LOC_279/a_8_216# OR2X1_LOC_44/Y 0.03fF
C14959 OR2X1_LOC_186/Y OR2X1_LOC_742/B 0.42fF
C14960 OR2X1_LOC_600/A OR2X1_LOC_257/Y 0.01fF
C14961 OR2X1_LOC_786/Y OR2X1_LOC_78/A 0.06fF
C14962 OR2X1_LOC_70/Y AND2X1_LOC_267/a_8_24# 0.01fF
C14963 OR2X1_LOC_311/Y OR2X1_LOC_829/a_36_216# 0.00fF
C14964 OR2X1_LOC_653/Y D_INPUT_0 0.30fF
C14965 AND2X1_LOC_334/a_8_24# OR2X1_LOC_316/Y 0.01fF
C14966 AND2X1_LOC_64/Y OR2X1_LOC_777/B 1.88fF
C14967 OR2X1_LOC_656/B OR2X1_LOC_814/A 0.07fF
C14968 AND2X1_LOC_456/Y AND2X1_LOC_717/B 0.00fF
C14969 OR2X1_LOC_185/A OR2X1_LOC_62/B 0.03fF
C14970 OR2X1_LOC_543/A OR2X1_LOC_318/B 0.20fF
C14971 OR2X1_LOC_19/B OR2X1_LOC_375/A 0.07fF
C14972 AND2X1_LOC_788/a_8_24# OR2X1_LOC_534/Y 0.23fF
C14973 AND2X1_LOC_624/B OR2X1_LOC_59/Y 0.00fF
C14974 OR2X1_LOC_719/A OR2X1_LOC_269/B 0.01fF
C14975 AND2X1_LOC_721/Y OR2X1_LOC_13/B 0.02fF
C14976 AND2X1_LOC_170/Y OR2X1_LOC_417/Y 0.15fF
C14977 AND2X1_LOC_56/B AND2X1_LOC_680/a_8_24# 0.03fF
C14978 OR2X1_LOC_32/B OR2X1_LOC_412/a_8_216# -0.01fF
C14979 AND2X1_LOC_557/a_8_24# OR2X1_LOC_89/A 0.01fF
C14980 OR2X1_LOC_3/Y AND2X1_LOC_554/B 0.02fF
C14981 VDD OR2X1_LOC_70/A 0.27fF
C14982 AND2X1_LOC_211/B AND2X1_LOC_211/a_36_24# 0.01fF
C14983 OR2X1_LOC_427/A OR2X1_LOC_95/Y 0.96fF
C14984 OR2X1_LOC_479/Y OR2X1_LOC_794/a_8_216# -0.03fF
C14985 OR2X1_LOC_65/a_8_216# OR2X1_LOC_52/B 0.06fF
C14986 AND2X1_LOC_31/Y OR2X1_LOC_723/a_36_216# 0.00fF
C14987 OR2X1_LOC_427/A OR2X1_LOC_368/A 0.40fF
C14988 AND2X1_LOC_31/Y OR2X1_LOC_302/A 0.14fF
C14989 OR2X1_LOC_31/Y OR2X1_LOC_619/Y 0.10fF
C14990 OR2X1_LOC_599/A AND2X1_LOC_537/Y 0.00fF
C14991 OR2X1_LOC_494/a_8_216# AND2X1_LOC_721/A 0.01fF
C14992 OR2X1_LOC_70/Y AND2X1_LOC_389/a_8_24# 0.11fF
C14993 OR2X1_LOC_60/a_36_216# OR2X1_LOC_585/A 0.02fF
C14994 OR2X1_LOC_12/Y OR2X1_LOC_536/a_8_216# 0.09fF
C14995 OR2X1_LOC_745/a_36_216# OR2X1_LOC_746/Y 0.00fF
C14996 OR2X1_LOC_82/a_8_216# OR2X1_LOC_46/A 0.01fF
C14997 AND2X1_LOC_372/a_8_24# OR2X1_LOC_493/Y 0.05fF
C14998 AND2X1_LOC_232/a_8_24# OR2X1_LOC_598/A 0.04fF
C14999 VDD AND2X1_LOC_31/Y 1.48fF
C15000 OR2X1_LOC_160/B OR2X1_LOC_68/B 12.78fF
C15001 AND2X1_LOC_330/a_8_24# OR2X1_LOC_331/Y 0.23fF
C15002 AND2X1_LOC_587/a_36_24# D_INPUT_6 0.00fF
C15003 OR2X1_LOC_182/B OR2X1_LOC_357/A 0.02fF
C15004 OR2X1_LOC_624/A OR2X1_LOC_222/a_8_216# 0.12fF
C15005 AND2X1_LOC_711/Y AND2X1_LOC_624/a_8_24# 0.01fF
C15006 OR2X1_LOC_3/Y OR2X1_LOC_696/Y 0.01fF
C15007 OR2X1_LOC_665/a_36_216# OR2X1_LOC_89/A 0.00fF
C15008 AND2X1_LOC_658/B AND2X1_LOC_657/A 0.37fF
C15009 OR2X1_LOC_417/A AND2X1_LOC_859/a_8_24# 0.00fF
C15010 OR2X1_LOC_292/Y AND2X1_LOC_848/A 0.00fF
C15011 OR2X1_LOC_446/Y OR2X1_LOC_87/A 0.29fF
C15012 OR2X1_LOC_95/Y AND2X1_LOC_464/a_8_24# 0.03fF
C15013 OR2X1_LOC_255/a_8_216# OR2X1_LOC_753/A 0.01fF
C15014 AND2X1_LOC_727/B OR2X1_LOC_142/Y 0.00fF
C15015 OR2X1_LOC_497/Y OR2X1_LOC_71/Y 0.03fF
C15016 OR2X1_LOC_185/A AND2X1_LOC_88/Y 0.03fF
C15017 AND2X1_LOC_79/a_8_24# OR2X1_LOC_557/A 0.01fF
C15018 OR2X1_LOC_482/Y OR2X1_LOC_13/B 0.03fF
C15019 AND2X1_LOC_463/a_8_24# OR2X1_LOC_408/Y 0.24fF
C15020 OR2X1_LOC_696/A AND2X1_LOC_242/B 1.99fF
C15021 OR2X1_LOC_333/B AND2X1_LOC_48/A 0.03fF
C15022 OR2X1_LOC_743/A OR2X1_LOC_246/A 2.92fF
C15023 OR2X1_LOC_516/Y AND2X1_LOC_244/A 0.04fF
C15024 AND2X1_LOC_64/Y OR2X1_LOC_831/B 0.03fF
C15025 OR2X1_LOC_271/a_8_216# OR2X1_LOC_368/A 0.47fF
C15026 OR2X1_LOC_817/a_8_216# INPUT_1 0.05fF
C15027 OR2X1_LOC_154/A OR2X1_LOC_223/A 0.03fF
C15028 AND2X1_LOC_390/B AND2X1_LOC_539/a_8_24# 0.03fF
C15029 OR2X1_LOC_134/Y AND2X1_LOC_541/a_8_24# 0.01fF
C15030 AND2X1_LOC_91/B AND2X1_LOC_766/a_8_24# 0.05fF
C15031 OR2X1_LOC_416/a_36_216# OR2X1_LOC_6/A 0.03fF
C15032 OR2X1_LOC_43/A AND2X1_LOC_655/a_8_24# 0.02fF
C15033 AND2X1_LOC_139/A OR2X1_LOC_26/Y 0.29fF
C15034 OR2X1_LOC_121/B AND2X1_LOC_491/a_8_24# 0.03fF
C15035 AND2X1_LOC_137/a_36_24# AND2X1_LOC_361/A 0.01fF
C15036 OR2X1_LOC_792/Y D_GATE_579 0.01fF
C15037 AND2X1_LOC_48/A OR2X1_LOC_99/B 0.81fF
C15038 OR2X1_LOC_91/Y AND2X1_LOC_795/Y 0.00fF
C15039 OR2X1_LOC_639/B AND2X1_LOC_428/a_36_24# 0.01fF
C15040 OR2X1_LOC_97/A AND2X1_LOC_7/B 2.92fF
C15041 OR2X1_LOC_516/Y OR2X1_LOC_108/Y 0.17fF
C15042 OR2X1_LOC_267/Y OR2X1_LOC_161/B 0.06fF
C15043 AND2X1_LOC_338/Y AND2X1_LOC_339/Y 0.14fF
C15044 OR2X1_LOC_628/Y AND2X1_LOC_629/Y 0.04fF
C15045 D_INPUT_7 OR2X1_LOC_51/B 0.05fF
C15046 OR2X1_LOC_164/Y OR2X1_LOC_437/A 0.00fF
C15047 INPUT_3 OR2X1_LOC_68/B 3.84fF
C15048 OR2X1_LOC_241/Y AND2X1_LOC_51/Y 0.16fF
C15049 OR2X1_LOC_51/Y OR2X1_LOC_504/a_8_216# 0.14fF
C15050 AND2X1_LOC_191/B AND2X1_LOC_792/B 0.18fF
C15051 OR2X1_LOC_774/B OR2X1_LOC_269/B 0.03fF
C15052 OR2X1_LOC_78/A OR2X1_LOC_199/B 0.00fF
C15053 AND2X1_LOC_572/a_36_24# OR2X1_LOC_595/A -0.02fF
C15054 OR2X1_LOC_80/a_8_216# OR2X1_LOC_46/A 0.02fF
C15055 OR2X1_LOC_434/a_8_216# OR2X1_LOC_339/A 0.10fF
C15056 OR2X1_LOC_39/A OR2X1_LOC_39/a_8_216# 0.09fF
C15057 OR2X1_LOC_69/A AND2X1_LOC_206/Y 0.13fF
C15058 OR2X1_LOC_269/B OR2X1_LOC_675/Y 0.50fF
C15059 OR2X1_LOC_31/Y OR2X1_LOC_22/A 0.05fF
C15060 OR2X1_LOC_87/A OR2X1_LOC_228/Y 1.13fF
C15061 AND2X1_LOC_711/Y AND2X1_LOC_624/B 0.03fF
C15062 AND2X1_LOC_40/Y OR2X1_LOC_716/a_36_216# 0.02fF
C15063 OR2X1_LOC_158/A OR2X1_LOC_428/A 1.02fF
C15064 OR2X1_LOC_70/Y OR2X1_LOC_67/Y 0.00fF
C15065 OR2X1_LOC_323/A OR2X1_LOC_51/Y 0.03fF
C15066 AND2X1_LOC_66/a_8_24# AND2X1_LOC_866/A 0.06fF
C15067 OR2X1_LOC_599/A AND2X1_LOC_796/A 0.11fF
C15068 OR2X1_LOC_269/B OR2X1_LOC_557/a_8_216# 0.01fF
C15069 OR2X1_LOC_45/B OR2X1_LOC_528/Y 0.25fF
C15070 OR2X1_LOC_527/Y AND2X1_LOC_795/Y 0.19fF
C15071 AND2X1_LOC_91/B OR2X1_LOC_645/a_36_216# 0.01fF
C15072 AND2X1_LOC_95/Y OR2X1_LOC_788/B 0.01fF
C15073 OR2X1_LOC_158/A OR2X1_LOC_595/A 0.01fF
C15074 OR2X1_LOC_675/A OR2X1_LOC_374/Y 0.26fF
C15075 OR2X1_LOC_121/Y OR2X1_LOC_715/B 0.08fF
C15076 AND2X1_LOC_390/a_8_24# OR2X1_LOC_533/Y 0.01fF
C15077 OR2X1_LOC_600/A AND2X1_LOC_464/A 0.03fF
C15078 OR2X1_LOC_51/Y OR2X1_LOC_744/a_8_216# 0.01fF
C15079 OR2X1_LOC_547/B AND2X1_LOC_36/Y 1.46fF
C15080 OR2X1_LOC_89/A AND2X1_LOC_783/a_36_24# 0.00fF
C15081 AND2X1_LOC_554/B AND2X1_LOC_772/a_8_24# 0.11fF
C15082 OR2X1_LOC_619/Y OR2X1_LOC_320/a_8_216# 0.01fF
C15083 OR2X1_LOC_279/Y AND2X1_LOC_562/Y 0.11fF
C15084 OR2X1_LOC_799/A OR2X1_LOC_593/B 0.17fF
C15085 AND2X1_LOC_564/B AND2X1_LOC_471/Y 0.00fF
C15086 AND2X1_LOC_110/a_8_24# OR2X1_LOC_161/B 0.01fF
C15087 OR2X1_LOC_541/A AND2X1_LOC_7/B 0.08fF
C15088 OR2X1_LOC_744/A AND2X1_LOC_769/Y 0.01fF
C15089 OR2X1_LOC_696/A AND2X1_LOC_841/B 0.02fF
C15090 OR2X1_LOC_585/A OR2X1_LOC_150/a_36_216# 0.00fF
C15091 OR2X1_LOC_7/A OR2X1_LOC_589/Y 0.03fF
C15092 AND2X1_LOC_64/Y OR2X1_LOC_575/A 0.07fF
C15093 AND2X1_LOC_215/Y OR2X1_LOC_158/A 0.01fF
C15094 AND2X1_LOC_56/B OR2X1_LOC_771/B 0.03fF
C15095 INPUT_0 OR2X1_LOC_375/Y 0.00fF
C15096 OR2X1_LOC_43/Y INPUT_0 0.01fF
C15097 OR2X1_LOC_45/B AND2X1_LOC_512/Y 0.03fF
C15098 AND2X1_LOC_595/a_8_24# OR2X1_LOC_160/B 0.04fF
C15099 AND2X1_LOC_18/Y OR2X1_LOC_641/A 0.05fF
C15100 AND2X1_LOC_56/B OR2X1_LOC_209/A 0.03fF
C15101 AND2X1_LOC_98/Y OR2X1_LOC_428/A 0.00fF
C15102 AND2X1_LOC_505/a_8_24# OR2X1_LOC_507/A 0.01fF
C15103 OR2X1_LOC_185/Y AND2X1_LOC_36/Y 0.10fF
C15104 AND2X1_LOC_8/Y OR2X1_LOC_771/B 0.09fF
C15105 AND2X1_LOC_7/B OR2X1_LOC_475/B 0.10fF
C15106 AND2X1_LOC_566/B OR2X1_LOC_56/A 0.58fF
C15107 OR2X1_LOC_756/Y OR2X1_LOC_756/a_36_216# 0.00fF
C15108 OR2X1_LOC_103/Y OR2X1_LOC_428/A 0.04fF
C15109 AND2X1_LOC_720/Y OR2X1_LOC_428/A 0.03fF
C15110 OR2X1_LOC_8/Y OR2X1_LOC_604/A 0.08fF
C15111 AND2X1_LOC_56/B OR2X1_LOC_776/A 0.00fF
C15112 AND2X1_LOC_715/Y AND2X1_LOC_841/B 0.07fF
C15113 OR2X1_LOC_264/Y AND2X1_LOC_44/Y 0.00fF
C15114 AND2X1_LOC_567/a_8_24# AND2X1_LOC_436/Y 0.00fF
C15115 AND2X1_LOC_658/B VDD 0.87fF
C15116 OR2X1_LOC_524/Y AND2X1_LOC_475/Y 0.01fF
C15117 OR2X1_LOC_97/A OR2X1_LOC_318/Y 0.02fF
C15118 OR2X1_LOC_273/a_36_216# OR2X1_LOC_300/Y 0.00fF
C15119 AND2X1_LOC_290/a_8_24# AND2X1_LOC_7/B 0.01fF
C15120 AND2X1_LOC_181/a_36_24# OR2X1_LOC_158/A 0.00fF
C15121 OR2X1_LOC_715/B OR2X1_LOC_538/A 0.01fF
C15122 AND2X1_LOC_110/Y OR2X1_LOC_78/B 0.03fF
C15123 OR2X1_LOC_711/A OR2X1_LOC_308/Y 0.02fF
C15124 OR2X1_LOC_269/a_8_216# AND2X1_LOC_7/B 0.01fF
C15125 AND2X1_LOC_22/Y AND2X1_LOC_95/Y 0.26fF
C15126 OR2X1_LOC_103/a_8_216# OR2X1_LOC_428/A 0.14fF
C15127 OR2X1_LOC_6/B OR2X1_LOC_235/B 0.07fF
C15128 INPUT_0 AND2X1_LOC_207/A 0.03fF
C15129 OR2X1_LOC_602/Y OR2X1_LOC_648/A 0.40fF
C15130 OR2X1_LOC_244/A OR2X1_LOC_68/B 0.04fF
C15131 OR2X1_LOC_60/Y OR2X1_LOC_59/Y 0.01fF
C15132 AND2X1_LOC_53/Y OR2X1_LOC_198/A 0.02fF
C15133 AND2X1_LOC_362/a_8_24# OR2X1_LOC_494/Y 0.11fF
C15134 OR2X1_LOC_589/A OR2X1_LOC_265/a_36_216# 0.00fF
C15135 OR2X1_LOC_186/Y AND2X1_LOC_314/a_8_24# 0.01fF
C15136 OR2X1_LOC_619/Y AND2X1_LOC_213/B 0.11fF
C15137 OR2X1_LOC_789/B OR2X1_LOC_691/Y 0.01fF
C15138 AND2X1_LOC_456/B AND2X1_LOC_860/A 0.08fF
C15139 OR2X1_LOC_97/A OR2X1_LOC_805/A 0.03fF
C15140 OR2X1_LOC_18/Y AND2X1_LOC_795/a_8_24# 0.02fF
C15141 OR2X1_LOC_106/Y AND2X1_LOC_560/B 0.07fF
C15142 INPUT_0 OR2X1_LOC_690/Y 0.01fF
C15143 OR2X1_LOC_769/B OR2X1_LOC_769/A 0.05fF
C15144 OR2X1_LOC_151/A OR2X1_LOC_324/A 0.07fF
C15145 OR2X1_LOC_600/A AND2X1_LOC_477/a_36_24# 0.00fF
C15146 OR2X1_LOC_85/a_8_216# AND2X1_LOC_216/A 0.47fF
C15147 D_INPUT_0 OR2X1_LOC_437/A 0.01fF
C15148 OR2X1_LOC_426/B OR2X1_LOC_298/a_8_216# 0.05fF
C15149 AND2X1_LOC_723/Y OR2X1_LOC_51/Y 0.17fF
C15150 OR2X1_LOC_666/A AND2X1_LOC_850/A 0.12fF
C15151 OR2X1_LOC_657/a_36_216# OR2X1_LOC_576/A 0.00fF
C15152 OR2X1_LOC_47/Y AND2X1_LOC_657/A 0.02fF
C15153 OR2X1_LOC_269/B OR2X1_LOC_779/A 0.01fF
C15154 AND2X1_LOC_600/a_8_24# OR2X1_LOC_777/B 0.03fF
C15155 OR2X1_LOC_176/Y AND2X1_LOC_784/A 0.06fF
C15156 AND2X1_LOC_22/Y OR2X1_LOC_99/Y 0.05fF
C15157 OR2X1_LOC_421/A OR2X1_LOC_432/a_8_216# 0.00fF
C15158 OR2X1_LOC_89/A OR2X1_LOC_184/a_8_216# 0.01fF
C15159 OR2X1_LOC_643/A AND2X1_LOC_44/Y 0.03fF
C15160 AND2X1_LOC_774/a_8_24# OR2X1_LOC_36/Y 0.01fF
C15161 OR2X1_LOC_158/A AND2X1_LOC_154/a_8_24# 0.09fF
C15162 OR2X1_LOC_102/a_8_216# AND2X1_LOC_342/Y 0.54fF
C15163 OR2X1_LOC_335/Y OR2X1_LOC_337/a_8_216# 0.07fF
C15164 OR2X1_LOC_124/Y AND2X1_LOC_44/Y 0.51fF
C15165 OR2X1_LOC_188/Y OR2X1_LOC_445/a_8_216# 0.01fF
C15166 OR2X1_LOC_715/B AND2X1_LOC_12/Y 0.03fF
C15167 AND2X1_LOC_753/a_8_24# AND2X1_LOC_18/Y 0.01fF
C15168 OR2X1_LOC_778/Y AND2X1_LOC_44/Y 0.36fF
C15169 AND2X1_LOC_763/a_8_24# AND2X1_LOC_40/Y 0.01fF
C15170 OR2X1_LOC_45/B OR2X1_LOC_682/Y 0.04fF
C15171 OR2X1_LOC_690/A AND2X1_LOC_219/A 0.45fF
C15172 AND2X1_LOC_31/Y OR2X1_LOC_737/a_36_216# 0.00fF
C15173 OR2X1_LOC_271/Y OR2X1_LOC_522/Y 0.01fF
C15174 AND2X1_LOC_486/Y OR2X1_LOC_59/Y 0.07fF
C15175 OR2X1_LOC_396/Y OR2X1_LOC_80/A 0.03fF
C15176 AND2X1_LOC_810/A AND2X1_LOC_856/A 0.01fF
C15177 OR2X1_LOC_736/Y OR2X1_LOC_269/B 0.07fF
C15178 OR2X1_LOC_78/A OR2X1_LOC_725/B 0.01fF
C15179 OR2X1_LOC_177/Y AND2X1_LOC_374/Y 0.01fF
C15180 OR2X1_LOC_185/A OR2X1_LOC_468/A 0.03fF
C15181 OR2X1_LOC_337/a_8_216# AND2X1_LOC_40/Y 0.01fF
C15182 OR2X1_LOC_348/Y AND2X1_LOC_59/Y 0.07fF
C15183 OR2X1_LOC_614/Y OR2X1_LOC_269/B 0.01fF
C15184 OR2X1_LOC_48/B AND2X1_LOC_434/Y 0.08fF
C15185 OR2X1_LOC_160/B OR2X1_LOC_219/a_8_216# 0.12fF
C15186 AND2X1_LOC_40/Y OR2X1_LOC_434/a_8_216# 0.01fF
C15187 OR2X1_LOC_36/Y OR2X1_LOC_253/Y 0.01fF
C15188 OR2X1_LOC_809/B OR2X1_LOC_624/A 0.28fF
C15189 OR2X1_LOC_235/B OR2X1_LOC_523/Y 0.00fF
C15190 OR2X1_LOC_326/a_8_216# AND2X1_LOC_95/Y 0.02fF
C15191 OR2X1_LOC_194/Y AND2X1_LOC_18/Y 0.50fF
C15192 OR2X1_LOC_18/Y AND2X1_LOC_219/Y 0.07fF
C15193 OR2X1_LOC_423/a_8_216# OR2X1_LOC_421/Y 0.44fF
C15194 OR2X1_LOC_40/Y OR2X1_LOC_69/Y 0.01fF
C15195 OR2X1_LOC_756/B OR2X1_LOC_811/A 0.01fF
C15196 OR2X1_LOC_114/Y AND2X1_LOC_18/Y 0.01fF
C15197 AND2X1_LOC_464/A OR2X1_LOC_372/a_8_216# 0.05fF
C15198 OR2X1_LOC_450/Y OR2X1_LOC_449/B 0.27fF
C15199 VDD OR2X1_LOC_461/A 0.01fF
C15200 OR2X1_LOC_557/A OR2X1_LOC_113/B 0.01fF
C15201 VDD OR2X1_LOC_809/a_8_216# 0.00fF
C15202 OR2X1_LOC_604/A OR2X1_LOC_52/B 0.14fF
C15203 OR2X1_LOC_745/a_8_216# OR2X1_LOC_52/B 0.02fF
C15204 OR2X1_LOC_604/A OR2X1_LOC_672/Y 0.07fF
C15205 OR2X1_LOC_864/A VDD 0.37fF
C15206 AND2X1_LOC_350/a_8_24# OR2X1_LOC_70/Y 0.06fF
C15207 OR2X1_LOC_502/A OR2X1_LOC_620/Y 0.07fF
C15208 OR2X1_LOC_426/B OR2X1_LOC_86/Y 0.05fF
C15209 OR2X1_LOC_45/B AND2X1_LOC_712/B 0.15fF
C15210 OR2X1_LOC_541/A OR2X1_LOC_805/A 0.02fF
C15211 AND2X1_LOC_362/B OR2X1_LOC_3/Y 0.00fF
C15212 AND2X1_LOC_716/a_8_24# OR2X1_LOC_59/Y 0.05fF
C15213 AND2X1_LOC_99/A AND2X1_LOC_99/Y 0.37fF
C15214 OR2X1_LOC_774/Y VDD 0.11fF
C15215 OR2X1_LOC_808/B OR2X1_LOC_739/A 0.05fF
C15216 OR2X1_LOC_369/a_8_216# AND2X1_LOC_211/B 0.04fF
C15217 OR2X1_LOC_389/B AND2X1_LOC_70/Y 0.02fF
C15218 VDD OR2X1_LOC_240/A 0.11fF
C15219 OR2X1_LOC_660/Y OR2X1_LOC_87/A 0.01fF
C15220 OR2X1_LOC_604/A OR2X1_LOC_73/a_36_216# 0.01fF
C15221 OR2X1_LOC_690/Y OR2X1_LOC_690/A 0.01fF
C15222 AND2X1_LOC_645/A AND2X1_LOC_447/Y 0.07fF
C15223 AND2X1_LOC_515/a_8_24# OR2X1_LOC_64/Y 0.07fF
C15224 VDD OR2X1_LOC_633/B 0.16fF
C15225 AND2X1_LOC_216/Y OR2X1_LOC_272/Y 0.01fF
C15226 OR2X1_LOC_49/A OR2X1_LOC_46/A 0.38fF
C15227 OR2X1_LOC_604/A OR2X1_LOC_418/a_36_216# 0.00fF
C15228 AND2X1_LOC_574/a_36_24# OR2X1_LOC_680/A 0.01fF
C15229 OR2X1_LOC_720/B OR2X1_LOC_721/a_8_216# 0.01fF
C15230 OR2X1_LOC_113/A AND2X1_LOC_44/Y 0.01fF
C15231 AND2X1_LOC_126/a_36_24# OR2X1_LOC_375/A 0.01fF
C15232 AND2X1_LOC_43/B OR2X1_LOC_623/B 0.03fF
C15233 OR2X1_LOC_585/A AND2X1_LOC_637/a_8_24# 0.01fF
C15234 OR2X1_LOC_235/B OR2X1_LOC_235/Y 0.01fF
C15235 AND2X1_LOC_456/B AND2X1_LOC_287/Y 0.48fF
C15236 OR2X1_LOC_805/A OR2X1_LOC_475/B 5.79fF
C15237 OR2X1_LOC_656/B AND2X1_LOC_517/a_8_24# 0.01fF
C15238 AND2X1_LOC_40/Y OR2X1_LOC_254/B 0.55fF
C15239 OR2X1_LOC_427/A OR2X1_LOC_257/a_36_216# 0.02fF
C15240 OR2X1_LOC_19/B OR2X1_LOC_549/A 0.02fF
C15241 AND2X1_LOC_718/a_8_24# OR2X1_LOC_44/Y -0.01fF
C15242 OR2X1_LOC_666/Y OR2X1_LOC_59/Y 0.09fF
C15243 OR2X1_LOC_154/A OR2X1_LOC_502/A 0.21fF
C15244 AND2X1_LOC_621/Y OR2X1_LOC_531/a_8_216# 0.04fF
C15245 OR2X1_LOC_54/Y OR2X1_LOC_382/A 0.10fF
C15246 AND2X1_LOC_509/Y AND2X1_LOC_474/Y 0.01fF
C15247 OR2X1_LOC_160/B AND2X1_LOC_666/a_8_24# 0.01fF
C15248 OR2X1_LOC_40/Y OR2X1_LOC_665/a_8_216# 0.01fF
C15249 OR2X1_LOC_71/Y AND2X1_LOC_249/a_8_24# 0.01fF
C15250 AND2X1_LOC_59/Y OR2X1_LOC_655/a_8_216# 0.00fF
C15251 OR2X1_LOC_808/B OR2X1_LOC_269/B 0.03fF
C15252 AND2X1_LOC_347/a_8_24# OR2X1_LOC_59/Y 0.02fF
C15253 OR2X1_LOC_160/A OR2X1_LOC_624/A 0.10fF
C15254 OR2X1_LOC_290/Y AND2X1_LOC_852/Y 0.06fF
C15255 AND2X1_LOC_663/a_8_24# GATE_579 0.20fF
C15256 OR2X1_LOC_40/Y AND2X1_LOC_537/Y 0.02fF
C15257 OR2X1_LOC_227/Y OR2X1_LOC_227/B 0.00fF
C15258 OR2X1_LOC_121/a_8_216# OR2X1_LOC_241/Y 0.05fF
C15259 AND2X1_LOC_12/Y OR2X1_LOC_215/Y 0.01fF
C15260 AND2X1_LOC_729/Y AND2X1_LOC_447/a_8_24# 0.02fF
C15261 AND2X1_LOC_359/a_36_24# OR2X1_LOC_92/Y 0.00fF
C15262 OR2X1_LOC_154/A OR2X1_LOC_571/B 0.01fF
C15263 AND2X1_LOC_658/A OR2X1_LOC_64/Y 0.09fF
C15264 AND2X1_LOC_61/Y OR2X1_LOC_291/Y 0.02fF
C15265 AND2X1_LOC_228/Y OR2X1_LOC_298/Y 0.00fF
C15266 OR2X1_LOC_76/Y OR2X1_LOC_811/A 0.03fF
C15267 OR2X1_LOC_186/Y OR2X1_LOC_468/a_8_216# 0.01fF
C15268 AND2X1_LOC_40/Y OR2X1_LOC_646/A 0.01fF
C15269 OR2X1_LOC_91/Y AND2X1_LOC_572/Y 0.03fF
C15270 OR2X1_LOC_635/a_8_216# OR2X1_LOC_87/A 0.01fF
C15271 AND2X1_LOC_364/Y AND2X1_LOC_324/a_8_24# 0.01fF
C15272 OR2X1_LOC_85/A OR2X1_LOC_118/Y 0.06fF
C15273 AND2X1_LOC_793/B AND2X1_LOC_793/a_8_24# 0.01fF
C15274 OR2X1_LOC_169/a_8_216# OR2X1_LOC_161/A 0.06fF
C15275 OR2X1_LOC_851/A OR2X1_LOC_155/A 0.17fF
C15276 OR2X1_LOC_641/a_8_216# OR2X1_LOC_814/A 0.14fF
C15277 AND2X1_LOC_214/A AND2X1_LOC_729/B 0.01fF
C15278 AND2X1_LOC_36/Y OR2X1_LOC_578/B 0.03fF
C15279 OR2X1_LOC_468/Y OR2X1_LOC_161/A 0.03fF
C15280 OR2X1_LOC_496/Y OR2X1_LOC_18/Y 0.00fF
C15281 OR2X1_LOC_673/Y OR2X1_LOC_137/B 0.03fF
C15282 AND2X1_LOC_477/A AND2X1_LOC_447/Y 0.15fF
C15283 OR2X1_LOC_185/A OR2X1_LOC_449/B 0.01fF
C15284 OR2X1_LOC_154/A OR2X1_LOC_400/A 0.06fF
C15285 OR2X1_LOC_527/a_8_216# OR2X1_LOC_31/Y 0.14fF
C15286 OR2X1_LOC_649/B OR2X1_LOC_660/B 0.72fF
C15287 OR2X1_LOC_276/A AND2X1_LOC_275/a_8_24# 0.09fF
C15288 OR2X1_LOC_848/B OR2X1_LOC_848/A 0.47fF
C15289 OR2X1_LOC_26/Y AND2X1_LOC_403/B 0.01fF
C15290 AND2X1_LOC_21/Y AND2X1_LOC_11/Y 0.17fF
C15291 OR2X1_LOC_764/Y OR2X1_LOC_48/B 0.02fF
C15292 OR2X1_LOC_314/a_8_216# OR2X1_LOC_70/Y 0.02fF
C15293 OR2X1_LOC_36/Y OR2X1_LOC_48/a_8_216# 0.01fF
C15294 OR2X1_LOC_9/Y D_INPUT_3 0.90fF
C15295 AND2X1_LOC_486/Y OR2X1_LOC_70/Y 0.03fF
C15296 OR2X1_LOC_216/A AND2X1_LOC_51/Y 0.36fF
C15297 OR2X1_LOC_36/Y AND2X1_LOC_286/Y 0.03fF
C15298 OR2X1_LOC_764/Y OR2X1_LOC_18/Y 0.01fF
C15299 AND2X1_LOC_794/B OR2X1_LOC_47/Y 0.02fF
C15300 OR2X1_LOC_648/A OR2X1_LOC_602/B 0.05fF
C15301 OR2X1_LOC_559/B AND2X1_LOC_3/Y 0.03fF
C15302 OR2X1_LOC_844/a_8_216# OR2X1_LOC_523/Y 0.01fF
C15303 AND2X1_LOC_59/Y OR2X1_LOC_810/A 0.04fF
C15304 OR2X1_LOC_6/B OR2X1_LOC_276/B 0.02fF
C15305 OR2X1_LOC_303/B OR2X1_LOC_593/B 0.03fF
C15306 OR2X1_LOC_411/Y D_INPUT_0 0.12fF
C15307 AND2X1_LOC_577/A OR2X1_LOC_189/A 0.07fF
C15308 AND2X1_LOC_658/A OR2X1_LOC_417/A 0.02fF
C15309 OR2X1_LOC_674/Y AND2X1_LOC_499/a_8_24# 0.24fF
C15310 AND2X1_LOC_391/Y INPUT_1 0.09fF
C15311 OR2X1_LOC_47/Y AND2X1_LOC_479/a_8_24# 0.01fF
C15312 OR2X1_LOC_219/B OR2X1_LOC_219/a_8_216# 0.02fF
C15313 AND2X1_LOC_580/A OR2X1_LOC_627/a_8_216# 0.06fF
C15314 OR2X1_LOC_91/A INPUT_1 0.15fF
C15315 AND2X1_LOC_43/a_8_24# AND2X1_LOC_43/B 0.10fF
C15316 OR2X1_LOC_639/B AND2X1_LOC_3/Y 0.16fF
C15317 OR2X1_LOC_262/Y OR2X1_LOC_85/A 0.04fF
C15318 OR2X1_LOC_126/a_8_216# OR2X1_LOC_39/A 0.03fF
C15319 OR2X1_LOC_80/Y OR2X1_LOC_52/B 0.02fF
C15320 OR2X1_LOC_102/a_36_216# AND2X1_LOC_721/A 0.00fF
C15321 OR2X1_LOC_756/B OR2X1_LOC_403/a_36_216# 0.01fF
C15322 AND2X1_LOC_494/a_8_24# OR2X1_LOC_391/A 0.23fF
C15323 OR2X1_LOC_651/A OR2X1_LOC_66/A 0.04fF
C15324 OR2X1_LOC_313/Y OR2X1_LOC_418/a_8_216# 0.01fF
C15325 OR2X1_LOC_3/Y OR2X1_LOC_595/a_8_216# 0.02fF
C15326 OR2X1_LOC_26/Y OR2X1_LOC_44/Y 0.60fF
C15327 OR2X1_LOC_642/a_8_216# AND2X1_LOC_8/Y 0.01fF
C15328 OR2X1_LOC_40/Y OR2X1_LOC_437/a_8_216# 0.01fF
C15329 AND2X1_LOC_675/A OR2X1_LOC_56/A 0.22fF
C15330 OR2X1_LOC_838/a_36_216# OR2X1_LOC_46/A 0.02fF
C15331 AND2X1_LOC_84/a_8_24# OR2X1_LOC_6/A 0.10fF
C15332 AND2X1_LOC_796/Y AND2X1_LOC_657/Y 0.03fF
C15333 OR2X1_LOC_137/Y OR2X1_LOC_267/A 0.02fF
C15334 VDD OR2X1_LOC_47/Y 2.54fF
C15335 OR2X1_LOC_6/B AND2X1_LOC_721/A 0.02fF
C15336 OR2X1_LOC_235/B AND2X1_LOC_47/Y 0.10fF
C15337 OR2X1_LOC_416/Y AND2X1_LOC_649/a_8_24# 0.01fF
C15338 OR2X1_LOC_89/A OR2X1_LOC_44/Y 0.47fF
C15339 OR2X1_LOC_280/Y OR2X1_LOC_36/Y 0.51fF
C15340 OR2X1_LOC_814/A OR2X1_LOC_785/B 0.35fF
C15341 AND2X1_LOC_191/Y AND2X1_LOC_740/B 0.09fF
C15342 AND2X1_LOC_660/A OR2X1_LOC_59/Y 0.00fF
C15343 OR2X1_LOC_185/A OR2X1_LOC_121/B 1.76fF
C15344 OR2X1_LOC_303/a_8_216# OR2X1_LOC_303/B 0.01fF
C15345 AND2X1_LOC_666/a_8_24# OR2X1_LOC_553/A 0.25fF
C15346 AND2X1_LOC_91/B OR2X1_LOC_317/B 0.03fF
C15347 OR2X1_LOC_330/Y OR2X1_LOC_532/B 0.02fF
C15348 OR2X1_LOC_861/a_8_216# OR2X1_LOC_814/A 0.01fF
C15349 OR2X1_LOC_820/Y OR2X1_LOC_44/Y 0.01fF
C15350 OR2X1_LOC_400/B OR2X1_LOC_624/B 0.05fF
C15351 AND2X1_LOC_276/Y AND2X1_LOC_361/A 0.04fF
C15352 AND2X1_LOC_91/B OR2X1_LOC_580/A 0.06fF
C15353 AND2X1_LOC_1/Y AND2X1_LOC_25/Y 0.31fF
C15354 OR2X1_LOC_476/B OR2X1_LOC_130/A 0.05fF
C15355 OR2X1_LOC_497/a_8_216# OR2X1_LOC_64/Y 0.06fF
C15356 AND2X1_LOC_661/A AND2X1_LOC_798/Y 0.02fF
C15357 AND2X1_LOC_138/a_8_24# OR2X1_LOC_46/A 0.01fF
C15358 OR2X1_LOC_468/Y AND2X1_LOC_51/Y 0.03fF
C15359 AND2X1_LOC_535/Y OR2X1_LOC_761/a_8_216# 0.00fF
C15360 OR2X1_LOC_76/A OR2X1_LOC_87/A 0.03fF
C15361 OR2X1_LOC_471/Y OR2X1_LOC_161/A 0.02fF
C15362 AND2X1_LOC_357/B AND2X1_LOC_222/Y 0.00fF
C15363 OR2X1_LOC_287/B AND2X1_LOC_815/a_8_24# 0.01fF
C15364 AND2X1_LOC_477/A AND2X1_LOC_448/Y 0.04fF
C15365 OR2X1_LOC_663/A OR2X1_LOC_340/a_8_216# 0.05fF
C15366 AND2X1_LOC_95/Y OR2X1_LOC_434/A 0.01fF
C15367 OR2X1_LOC_154/A AND2X1_LOC_48/A 0.19fF
C15368 VDD OR2X1_LOC_608/Y 0.06fF
C15369 OR2X1_LOC_160/A OR2X1_LOC_447/Y 0.03fF
C15370 OR2X1_LOC_291/Y AND2X1_LOC_852/Y 0.36fF
C15371 AND2X1_LOC_22/Y AND2X1_LOC_41/Y 0.02fF
C15372 OR2X1_LOC_509/A OR2X1_LOC_227/Y 0.11fF
C15373 OR2X1_LOC_22/Y OR2X1_LOC_36/Y 2.68fF
C15374 AND2X1_LOC_364/a_36_24# OR2X1_LOC_437/A 0.00fF
C15375 OR2X1_LOC_641/a_8_216# OR2X1_LOC_341/a_8_216# 0.47fF
C15376 AND2X1_LOC_486/Y OR2X1_LOC_184/Y 0.25fF
C15377 AND2X1_LOC_32/a_8_24# D_INPUT_0 0.04fF
C15378 AND2X1_LOC_170/B AND2X1_LOC_436/B 0.01fF
C15379 OR2X1_LOC_3/Y OR2X1_LOC_431/a_8_216# 0.01fF
C15380 OR2X1_LOC_148/A OR2X1_LOC_87/A 0.03fF
C15381 AND2X1_LOC_851/B OR2X1_LOC_18/Y 0.10fF
C15382 OR2X1_LOC_643/A OR2X1_LOC_720/B 0.03fF
C15383 OR2X1_LOC_696/A AND2X1_LOC_543/Y 0.03fF
C15384 AND2X1_LOC_572/Y D_INPUT_3 0.31fF
C15385 OR2X1_LOC_503/Y OR2X1_LOC_39/A 0.01fF
C15386 AND2X1_LOC_486/Y OR2X1_LOC_437/Y 0.23fF
C15387 AND2X1_LOC_537/Y OR2X1_LOC_7/A 4.03fF
C15388 D_INPUT_0 OR2X1_LOC_753/A 0.27fF
C15389 OR2X1_LOC_846/B AND2X1_LOC_51/Y 0.13fF
C15390 OR2X1_LOC_486/a_8_216# OR2X1_LOC_486/B 0.05fF
C15391 OR2X1_LOC_268/Y AND2X1_LOC_786/Y 0.06fF
C15392 OR2X1_LOC_154/A AND2X1_LOC_106/a_8_24# 0.04fF
C15393 AND2X1_LOC_1/Y AND2X1_LOC_51/Y 0.01fF
C15394 AND2X1_LOC_456/B AND2X1_LOC_562/Y 0.03fF
C15395 OR2X1_LOC_334/B AND2X1_LOC_31/Y 0.02fF
C15396 OR2X1_LOC_19/B OR2X1_LOC_83/a_36_216# 0.01fF
C15397 OR2X1_LOC_516/Y OR2X1_LOC_373/Y 0.07fF
C15398 AND2X1_LOC_392/A AND2X1_LOC_212/a_36_24# 0.01fF
C15399 AND2X1_LOC_326/B OR2X1_LOC_437/A 0.01fF
C15400 OR2X1_LOC_175/Y OR2X1_LOC_214/A 0.01fF
C15401 OR2X1_LOC_709/A OR2X1_LOC_714/a_8_216# 0.04fF
C15402 D_INPUT_3 AND2X1_LOC_852/Y 0.01fF
C15403 OR2X1_LOC_557/A OR2X1_LOC_532/B 0.00fF
C15404 OR2X1_LOC_136/a_8_216# OR2X1_LOC_136/Y 0.01fF
C15405 OR2X1_LOC_549/a_8_216# OR2X1_LOC_577/Y 0.01fF
C15406 OR2X1_LOC_285/Y OR2X1_LOC_285/B 0.03fF
C15407 OR2X1_LOC_433/a_36_216# AND2X1_LOC_648/B 0.00fF
C15408 D_INPUT_3 OR2X1_LOC_6/a_36_216# 0.00fF
C15409 OR2X1_LOC_502/A OR2X1_LOC_560/A 0.62fF
C15410 INPUT_1 OR2X1_LOC_27/Y 0.20fF
C15411 OR2X1_LOC_175/Y AND2X1_LOC_7/B 0.03fF
C15412 OR2X1_LOC_471/Y AND2X1_LOC_51/Y 0.00fF
C15413 OR2X1_LOC_405/A OR2X1_LOC_358/A 0.25fF
C15414 OR2X1_LOC_844/a_8_216# AND2X1_LOC_47/Y 0.01fF
C15415 AND2X1_LOC_817/a_8_24# D_INPUT_1 0.07fF
C15416 OR2X1_LOC_600/A AND2X1_LOC_750/a_8_24# 0.01fF
C15417 AND2X1_LOC_91/B AND2X1_LOC_44/Y 0.22fF
C15418 AND2X1_LOC_64/Y OR2X1_LOC_161/B 2.43fF
C15419 OR2X1_LOC_84/B OR2X1_LOC_84/A 0.04fF
C15420 AND2X1_LOC_687/A AND2X1_LOC_685/a_36_24# 0.00fF
C15421 OR2X1_LOC_696/A OR2X1_LOC_589/A 0.36fF
C15422 OR2X1_LOC_347/B OR2X1_LOC_675/Y 0.09fF
C15423 OR2X1_LOC_675/A OR2X1_LOC_532/B -0.00fF
C15424 OR2X1_LOC_696/A OR2X1_LOC_322/Y 0.16fF
C15425 AND2X1_LOC_401/a_8_24# OR2X1_LOC_80/A 0.07fF
C15426 OR2X1_LOC_51/Y OR2X1_LOC_142/Y 0.02fF
C15427 OR2X1_LOC_643/Y OR2X1_LOC_814/A 0.02fF
C15428 OR2X1_LOC_48/B OR2X1_LOC_172/a_36_216# 0.00fF
C15429 OR2X1_LOC_691/Y AND2X1_LOC_7/B 0.03fF
C15430 OR2X1_LOC_853/a_8_216# OR2X1_LOC_857/A 0.01fF
C15431 AND2X1_LOC_92/Y OR2X1_LOC_771/B 0.05fF
C15432 AND2X1_LOC_490/a_8_24# D_INPUT_1 0.02fF
C15433 OR2X1_LOC_218/Y OR2X1_LOC_215/A 0.24fF
C15434 AND2X1_LOC_436/B OR2X1_LOC_331/Y 0.02fF
C15435 OR2X1_LOC_78/B OR2X1_LOC_537/a_36_216# 0.02fF
C15436 AND2X1_LOC_850/A OR2X1_LOC_13/B 0.28fF
C15437 AND2X1_LOC_811/a_8_24# AND2X1_LOC_222/Y 0.01fF
C15438 OR2X1_LOC_756/B OR2X1_LOC_777/B 0.05fF
C15439 OR2X1_LOC_40/Y OR2X1_LOC_171/a_8_216# 0.01fF
C15440 OR2X1_LOC_351/B OR2X1_LOC_338/B 0.74fF
C15441 OR2X1_LOC_820/A OR2X1_LOC_749/Y 0.01fF
C15442 OR2X1_LOC_373/a_8_216# OR2X1_LOC_373/Y 0.03fF
C15443 VDD OR2X1_LOC_501/A -0.00fF
C15444 OR2X1_LOC_417/A AND2X1_LOC_814/a_8_24# 0.11fF
C15445 OR2X1_LOC_759/A AND2X1_LOC_792/a_8_24# 0.08fF
C15446 OR2X1_LOC_696/A AND2X1_LOC_337/a_8_24# 0.02fF
C15447 OR2X1_LOC_518/a_36_216# AND2X1_LOC_326/B 0.00fF
C15448 AND2X1_LOC_92/Y OR2X1_LOC_776/A 0.02fF
C15449 OR2X1_LOC_74/A AND2X1_LOC_793/Y 0.09fF
C15450 VDD AND2X1_LOC_760/a_8_24# -0.00fF
C15451 AND2X1_LOC_632/a_8_24# AND2X1_LOC_623/a_8_24# 0.23fF
C15452 OR2X1_LOC_476/a_8_216# OR2X1_LOC_223/A 0.42fF
C15453 AND2X1_LOC_195/a_8_24# AND2X1_LOC_199/A 0.00fF
C15454 OR2X1_LOC_97/A OR2X1_LOC_648/B 0.00fF
C15455 D_GATE_865 OR2X1_LOC_561/B 0.02fF
C15456 OR2X1_LOC_786/A OR2X1_LOC_266/A 0.17fF
C15457 OR2X1_LOC_66/A OR2X1_LOC_338/A 0.01fF
C15458 OR2X1_LOC_375/A OR2X1_LOC_725/a_36_216# 0.00fF
C15459 VDD OR2X1_LOC_121/A 0.12fF
C15460 OR2X1_LOC_237/a_8_216# OR2X1_LOC_437/A 0.15fF
C15461 OR2X1_LOC_744/A AND2X1_LOC_783/B 0.01fF
C15462 AND2X1_LOC_116/B AND2X1_LOC_116/a_8_24# 0.01fF
C15463 OR2X1_LOC_291/Y AND2X1_LOC_647/B 0.09fF
C15464 OR2X1_LOC_85/A AND2X1_LOC_215/a_36_24# 0.00fF
C15465 OR2X1_LOC_49/A INPUT_2 0.01fF
C15466 OR2X1_LOC_786/Y OR2X1_LOC_814/A 0.03fF
C15467 AND2X1_LOC_94/Y OR2X1_LOC_397/Y 0.09fF
C15468 OR2X1_LOC_375/A OR2X1_LOC_550/B 0.01fF
C15469 OR2X1_LOC_803/A AND2X1_LOC_7/B 0.00fF
C15470 OR2X1_LOC_773/a_8_216# D_INPUT_1 0.01fF
C15471 OR2X1_LOC_276/B AND2X1_LOC_47/Y 0.08fF
C15472 OR2X1_LOC_597/A OR2X1_LOC_12/Y 0.32fF
C15473 OR2X1_LOC_696/A AND2X1_LOC_654/B 0.12fF
C15474 OR2X1_LOC_604/A OR2X1_LOC_281/Y 0.09fF
C15475 OR2X1_LOC_696/A OR2X1_LOC_495/Y 0.03fF
C15476 OR2X1_LOC_186/Y OR2X1_LOC_66/A 0.44fF
C15477 OR2X1_LOC_256/A OR2X1_LOC_47/Y 0.04fF
C15478 OR2X1_LOC_22/Y OR2X1_LOC_419/Y 0.03fF
C15479 OR2X1_LOC_40/Y OR2X1_LOC_13/Y 0.03fF
C15480 OR2X1_LOC_739/A OR2X1_LOC_703/Y 0.02fF
C15481 OR2X1_LOC_866/B OR2X1_LOC_391/A 0.09fF
C15482 OR2X1_LOC_185/Y OR2X1_LOC_571/Y 0.03fF
C15483 OR2X1_LOC_680/A OR2X1_LOC_142/Y 14.00fF
C15484 OR2X1_LOC_61/A OR2X1_LOC_78/B 0.03fF
C15485 OR2X1_LOC_364/A OR2X1_LOC_374/a_8_216# 0.05fF
C15486 OR2X1_LOC_471/Y OR2X1_LOC_551/B 0.19fF
C15487 AND2X1_LOC_340/Y AND2X1_LOC_219/Y 0.07fF
C15488 VDD AND2X1_LOC_469/Y 0.21fF
C15489 OR2X1_LOC_604/A OR2X1_LOC_253/Y 0.02fF
C15490 AND2X1_LOC_64/Y OR2X1_LOC_61/Y 0.00fF
C15491 OR2X1_LOC_289/Y OR2X1_LOC_31/Y 0.03fF
C15492 AND2X1_LOC_810/B AND2X1_LOC_434/Y 0.00fF
C15493 OR2X1_LOC_16/A OR2X1_LOC_597/a_36_216# 0.00fF
C15494 AND2X1_LOC_539/Y OR2X1_LOC_761/Y 0.02fF
C15495 OR2X1_LOC_450/Y OR2X1_LOC_452/a_8_216# 0.01fF
C15496 OR2X1_LOC_186/Y AND2X1_LOC_311/a_8_24# 0.23fF
C15497 OR2X1_LOC_596/A OR2X1_LOC_702/a_8_216# 0.01fF
C15498 OR2X1_LOC_40/Y OR2X1_LOC_627/Y 0.03fF
C15499 OR2X1_LOC_768/A OR2X1_LOC_113/B 0.16fF
C15500 OR2X1_LOC_643/Y OR2X1_LOC_341/a_8_216# 0.01fF
C15501 OR2X1_LOC_318/Y OR2X1_LOC_175/Y 0.07fF
C15502 AND2X1_LOC_81/B OR2X1_LOC_508/Y 0.65fF
C15503 OR2X1_LOC_40/Y AND2X1_LOC_500/Y 0.02fF
C15504 AND2X1_LOC_732/B VDD 0.41fF
C15505 OR2X1_LOC_6/B AND2X1_LOC_70/Y 0.50fF
C15506 AND2X1_LOC_521/a_8_24# OR2X1_LOC_235/B 0.02fF
C15507 AND2X1_LOC_22/Y OR2X1_LOC_608/a_36_216# 0.02fF
C15508 OR2X1_LOC_464/A OR2X1_LOC_161/B 0.03fF
C15509 OR2X1_LOC_325/Y AND2X1_LOC_110/Y 0.01fF
C15510 OR2X1_LOC_329/B AND2X1_LOC_476/Y 0.04fF
C15511 OR2X1_LOC_269/B OR2X1_LOC_703/Y 0.15fF
C15512 OR2X1_LOC_308/a_8_216# AND2X1_LOC_44/Y 0.01fF
C15513 OR2X1_LOC_512/A OR2X1_LOC_161/B 0.01fF
C15514 AND2X1_LOC_12/Y OR2X1_LOC_338/B 0.01fF
C15515 OR2X1_LOC_256/Y OR2X1_LOC_12/Y 0.07fF
C15516 AND2X1_LOC_326/B AND2X1_LOC_715/A 0.02fF
C15517 OR2X1_LOC_287/B OR2X1_LOC_579/A 0.01fF
C15518 OR2X1_LOC_666/a_36_216# AND2X1_LOC_658/A 0.02fF
C15519 OR2X1_LOC_47/Y OR2X1_LOC_67/Y 0.03fF
C15520 OR2X1_LOC_756/B OR2X1_LOC_545/A 0.13fF
C15521 OR2X1_LOC_586/Y OR2X1_LOC_428/A 0.07fF
C15522 AND2X1_LOC_534/a_8_24# OR2X1_LOC_354/A 0.02fF
C15523 OR2X1_LOC_151/A OR2X1_LOC_735/a_8_216# 0.02fF
C15524 AND2X1_LOC_39/a_36_24# AND2X1_LOC_44/Y 0.00fF
C15525 AND2X1_LOC_463/B OR2X1_LOC_588/A 0.32fF
C15526 OR2X1_LOC_502/A OR2X1_LOC_435/A 0.01fF
C15527 OR2X1_LOC_158/A AND2X1_LOC_512/Y 0.07fF
C15528 AND2X1_LOC_357/A AND2X1_LOC_364/Y 0.01fF
C15529 OR2X1_LOC_654/A AND2X1_LOC_36/Y 0.05fF
C15530 OR2X1_LOC_696/A OR2X1_LOC_43/A 0.61fF
C15531 AND2X1_LOC_181/a_8_24# OR2X1_LOC_108/Y 0.01fF
C15532 INPUT_0 OR2X1_LOC_461/B 0.13fF
C15533 AND2X1_LOC_338/Y OR2X1_LOC_619/Y 0.03fF
C15534 AND2X1_LOC_47/Y OR2X1_LOC_779/B 0.01fF
C15535 OR2X1_LOC_51/Y AND2X1_LOC_338/a_8_24# 0.01fF
C15536 OR2X1_LOC_175/Y OR2X1_LOC_805/A 0.03fF
C15537 AND2X1_LOC_713/Y AND2X1_LOC_605/Y 0.00fF
C15538 AND2X1_LOC_191/B OR2X1_LOC_666/A 0.03fF
C15539 AND2X1_LOC_866/A AND2X1_LOC_563/Y 0.03fF
C15540 OR2X1_LOC_87/A OR2X1_LOC_722/B 0.01fF
C15541 AND2X1_LOC_570/Y OR2X1_LOC_744/A 0.03fF
C15542 OR2X1_LOC_631/B OR2X1_LOC_115/B 0.05fF
C15543 AND2X1_LOC_852/Y OR2X1_LOC_171/Y 0.02fF
C15544 AND2X1_LOC_853/Y OR2X1_LOC_171/a_36_216# 0.00fF
C15545 AND2X1_LOC_352/B OR2X1_LOC_91/A 0.04fF
C15546 OR2X1_LOC_179/a_8_216# OR2X1_LOC_600/A 0.01fF
C15547 AND2X1_LOC_367/A OR2X1_LOC_494/Y 0.01fF
C15548 OR2X1_LOC_7/A OR2X1_LOC_743/Y 0.02fF
C15549 OR2X1_LOC_118/a_8_216# OR2X1_LOC_65/B 0.00fF
C15550 AND2X1_LOC_392/A AND2X1_LOC_392/a_36_24# 0.01fF
C15551 OR2X1_LOC_354/A AND2X1_LOC_110/Y 0.01fF
C15552 AND2X1_LOC_367/A AND2X1_LOC_363/Y 0.11fF
C15553 OR2X1_LOC_691/Y OR2X1_LOC_805/A 0.01fF
C15554 OR2X1_LOC_91/Y AND2X1_LOC_787/A 0.85fF
C15555 AND2X1_LOC_473/Y OR2X1_LOC_6/A 0.00fF
C15556 OR2X1_LOC_779/a_8_216# OR2X1_LOC_779/A 0.01fF
C15557 OR2X1_LOC_442/Y AND2X1_LOC_444/a_8_24# 0.23fF
C15558 AND2X1_LOC_774/a_8_24# OR2X1_LOC_306/Y 0.01fF
C15559 OR2X1_LOC_313/a_8_216# OR2X1_LOC_12/Y 0.01fF
C15560 AND2X1_LOC_12/Y OR2X1_LOC_35/A 0.01fF
C15561 AND2X1_LOC_580/B AND2X1_LOC_580/a_8_24# 0.03fF
C15562 AND2X1_LOC_715/Y OR2X1_LOC_43/A 0.01fF
C15563 OR2X1_LOC_769/A OR2X1_LOC_637/Y 0.05fF
C15564 OR2X1_LOC_348/a_8_216# AND2X1_LOC_12/Y 0.01fF
C15565 AND2X1_LOC_715/A AND2X1_LOC_276/a_8_24# 0.11fF
C15566 OR2X1_LOC_739/A OR2X1_LOC_596/A 0.00fF
C15567 OR2X1_LOC_179/a_36_216# OR2X1_LOC_56/A 0.00fF
C15568 AND2X1_LOC_372/a_8_24# OR2X1_LOC_541/A 0.01fF
C15569 OR2X1_LOC_748/A OR2X1_LOC_428/A 0.04fF
C15570 OR2X1_LOC_336/a_36_216# OR2X1_LOC_468/Y 0.00fF
C15571 OR2X1_LOC_45/B OR2X1_LOC_26/Y 0.22fF
C15572 AND2X1_LOC_56/B AND2X1_LOC_256/a_8_24# 0.01fF
C15573 AND2X1_LOC_392/A AND2X1_LOC_841/B 0.07fF
C15574 OR2X1_LOC_850/B OR2X1_LOC_287/A 0.22fF
C15575 AND2X1_LOC_391/Y OR2X1_LOC_517/A 0.00fF
C15576 OR2X1_LOC_36/Y AND2X1_LOC_445/a_36_24# 0.01fF
C15577 OR2X1_LOC_92/Y OR2X1_LOC_56/A 0.54fF
C15578 OR2X1_LOC_421/A OR2X1_LOC_432/Y 0.01fF
C15579 OR2X1_LOC_91/A OR2X1_LOC_517/A 4.66fF
C15580 OR2X1_LOC_158/A AND2X1_LOC_342/Y 0.05fF
C15581 OR2X1_LOC_326/B AND2X1_LOC_70/Y 0.39fF
C15582 VDD OR2X1_LOC_784/Y 0.08fF
C15583 AND2X1_LOC_712/Y AND2X1_LOC_454/Y 0.01fF
C15584 OR2X1_LOC_715/B AND2X1_LOC_59/Y 0.08fF
C15585 OR2X1_LOC_448/B OR2X1_LOC_78/A 0.11fF
C15586 OR2X1_LOC_51/Y OR2X1_LOC_40/a_8_216# 0.01fF
C15587 VDD OR2X1_LOC_625/Y 1.30fF
C15588 OR2X1_LOC_76/Y OR2X1_LOC_344/A 0.02fF
C15589 AND2X1_LOC_18/Y OR2X1_LOC_541/B 0.06fF
C15590 OR2X1_LOC_45/B OR2X1_LOC_89/A 0.05fF
C15591 OR2X1_LOC_509/a_8_216# AND2X1_LOC_81/B 0.00fF
C15592 OR2X1_LOC_840/A AND2X1_LOC_41/A 0.01fF
C15593 AND2X1_LOC_95/Y OR2X1_LOC_741/Y 0.17fF
C15594 AND2X1_LOC_212/Y OR2X1_LOC_52/B 0.07fF
C15595 OR2X1_LOC_3/Y AND2X1_LOC_636/a_8_24# 0.01fF
C15596 AND2X1_LOC_550/A AND2X1_LOC_658/A 9.73fF
C15597 OR2X1_LOC_679/Y OR2X1_LOC_679/B 0.20fF
C15598 AND2X1_LOC_767/a_8_24# AND2X1_LOC_396/a_8_24# 0.23fF
C15599 VDD OR2X1_LOC_738/A 0.05fF
C15600 AND2X1_LOC_819/a_8_24# AND2X1_LOC_618/a_8_24# 0.23fF
C15601 OR2X1_LOC_154/A OR2X1_LOC_772/A 0.01fF
C15602 AND2X1_LOC_99/A OR2X1_LOC_122/A 0.01fF
C15603 OR2X1_LOC_596/A OR2X1_LOC_269/B 0.05fF
C15604 AND2X1_LOC_364/Y OR2X1_LOC_48/B 0.03fF
C15605 OR2X1_LOC_809/B OR2X1_LOC_161/A 0.07fF
C15606 OR2X1_LOC_326/B OR2X1_LOC_703/A 0.00fF
C15607 OR2X1_LOC_318/A OR2X1_LOC_479/Y 0.00fF
C15608 OR2X1_LOC_6/B OR2X1_LOC_116/a_8_216# -0.01fF
C15609 OR2X1_LOC_485/Y OR2X1_LOC_36/Y 0.06fF
C15610 OR2X1_LOC_65/B OR2X1_LOC_56/A 0.04fF
C15611 OR2X1_LOC_51/Y AND2X1_LOC_453/a_8_24# 0.01fF
C15612 OR2X1_LOC_682/Y OR2X1_LOC_158/A 0.35fF
C15613 OR2X1_LOC_304/Y OR2X1_LOC_428/A 0.53fF
C15614 OR2X1_LOC_160/B OR2X1_LOC_87/A 6.33fF
C15615 OR2X1_LOC_244/A AND2X1_LOC_235/a_8_24# 0.01fF
C15616 OR2X1_LOC_177/Y OR2X1_LOC_280/Y 0.00fF
C15617 OR2X1_LOC_89/A OR2X1_LOC_382/A 0.26fF
C15618 AND2X1_LOC_53/Y AND2X1_LOC_763/B 0.12fF
C15619 AND2X1_LOC_858/B AND2X1_LOC_624/A 0.42fF
C15620 AND2X1_LOC_601/a_8_24# OR2X1_LOC_78/B 0.08fF
C15621 OR2X1_LOC_849/A AND2X1_LOC_18/Y 0.01fF
C15622 OR2X1_LOC_438/Y OR2X1_LOC_427/A 0.04fF
C15623 OR2X1_LOC_368/a_36_216# OR2X1_LOC_312/Y 0.00fF
C15624 AND2X1_LOC_456/B AND2X1_LOC_287/a_8_24# 0.01fF
C15625 AND2X1_LOC_464/a_36_24# OR2X1_LOC_56/A 0.00fF
C15626 OR2X1_LOC_158/A OR2X1_LOC_279/a_8_216# 0.01fF
C15627 OR2X1_LOC_283/a_36_216# OR2X1_LOC_51/Y 0.00fF
C15628 OR2X1_LOC_653/Y AND2X1_LOC_749/a_36_24# 0.00fF
C15629 OR2X1_LOC_479/Y OR2X1_LOC_151/A 0.07fF
C15630 OR2X1_LOC_844/a_36_216# OR2X1_LOC_113/B 0.00fF
C15631 OR2X1_LOC_517/A AND2X1_LOC_573/A 0.07fF
C15632 OR2X1_LOC_756/B OR2X1_LOC_652/a_8_216# 0.01fF
C15633 OR2X1_LOC_642/a_8_216# AND2X1_LOC_92/Y 0.01fF
C15634 OR2X1_LOC_485/A AND2X1_LOC_500/B 0.24fF
C15635 OR2X1_LOC_271/Y OR2X1_LOC_56/A 0.03fF
C15636 OR2X1_LOC_473/A OR2X1_LOC_130/a_8_216# 0.18fF
C15637 OR2X1_LOC_604/A OR2X1_LOC_280/Y 0.10fF
C15638 OR2X1_LOC_329/Y AND2X1_LOC_390/B 0.02fF
C15639 AND2X1_LOC_98/Y AND2X1_LOC_342/Y 0.03fF
C15640 OR2X1_LOC_298/Y AND2X1_LOC_857/Y 0.01fF
C15641 AND2X1_LOC_41/A OR2X1_LOC_222/A 0.03fF
C15642 OR2X1_LOC_427/A OR2X1_LOC_427/Y 0.01fF
C15643 OR2X1_LOC_324/a_8_216# OR2X1_LOC_739/A 0.01fF
C15644 OR2X1_LOC_223/A OR2X1_LOC_605/Y 0.15fF
C15645 OR2X1_LOC_51/Y OR2X1_LOC_238/Y 0.01fF
C15646 OR2X1_LOC_154/A OR2X1_LOC_201/A 0.01fF
C15647 OR2X1_LOC_448/A OR2X1_LOC_375/A 0.09fF
C15648 OR2X1_LOC_856/B OR2X1_LOC_185/A 0.07fF
C15649 AND2X1_LOC_396/a_36_24# AND2X1_LOC_3/Y 0.00fF
C15650 OR2X1_LOC_155/A OR2X1_LOC_78/A 0.54fF
C15651 AND2X1_LOC_337/B AND2X1_LOC_436/Y 0.54fF
C15652 AND2X1_LOC_22/Y OR2X1_LOC_434/A 0.31fF
C15653 OR2X1_LOC_185/Y OR2X1_LOC_571/a_36_216# 0.17fF
C15654 AND2X1_LOC_600/a_8_24# OR2X1_LOC_161/B 0.01fF
C15655 OR2X1_LOC_158/A AND2X1_LOC_712/B 0.29fF
C15656 OR2X1_LOC_427/A AND2X1_LOC_621/Y 0.09fF
C15657 OR2X1_LOC_185/Y OR2X1_LOC_274/Y 0.02fF
C15658 OR2X1_LOC_743/A OR2X1_LOC_743/a_8_216# 0.09fF
C15659 OR2X1_LOC_158/A OR2X1_LOC_54/Y 0.36fF
C15660 OR2X1_LOC_382/Y OR2X1_LOC_820/B 0.90fF
C15661 OR2X1_LOC_671/Y OR2X1_LOC_46/A 0.06fF
C15662 OR2X1_LOC_185/Y OR2X1_LOC_392/A 0.00fF
C15663 OR2X1_LOC_808/A OR2X1_LOC_269/B 0.07fF
C15664 OR2X1_LOC_532/B OR2X1_LOC_548/a_8_216# 0.01fF
C15665 AND2X1_LOC_548/Y OR2X1_LOC_74/A 0.11fF
C15666 OR2X1_LOC_542/B OR2X1_LOC_254/a_8_216# 0.05fF
C15667 AND2X1_LOC_76/Y OR2X1_LOC_265/Y 0.03fF
C15668 OR2X1_LOC_400/B OR2X1_LOC_400/a_8_216# 0.47fF
C15669 OR2X1_LOC_160/A OR2X1_LOC_161/A 3.92fF
C15670 OR2X1_LOC_261/a_8_216# AND2X1_LOC_663/B 0.03fF
C15671 OR2X1_LOC_604/A OR2X1_LOC_295/a_36_216# 0.01fF
C15672 AND2X1_LOC_35/a_8_24# OR2X1_LOC_18/Y 0.01fF
C15673 AND2X1_LOC_624/A AND2X1_LOC_573/A 0.03fF
C15674 OR2X1_LOC_40/Y OR2X1_LOC_295/Y 0.07fF
C15675 OR2X1_LOC_446/B OR2X1_LOC_317/B 0.14fF
C15676 OR2X1_LOC_364/B AND2X1_LOC_47/Y 0.00fF
C15677 OR2X1_LOC_709/A AND2X1_LOC_47/Y 0.03fF
C15678 AND2X1_LOC_649/Y AND2X1_LOC_786/Y 0.01fF
C15679 AND2X1_LOC_59/Y OR2X1_LOC_215/Y 0.31fF
C15680 OR2X1_LOC_604/A OR2X1_LOC_22/Y 0.10fF
C15681 AND2X1_LOC_47/Y AND2X1_LOC_295/a_8_24# 0.01fF
C15682 OR2X1_LOC_160/B AND2X1_LOC_45/a_36_24# 0.00fF
C15683 AND2X1_LOC_303/B OR2X1_LOC_619/Y -0.03fF
C15684 AND2X1_LOC_87/a_8_24# OR2X1_LOC_65/B 0.17fF
C15685 AND2X1_LOC_375/a_8_24# OR2X1_LOC_753/A 0.23fF
C15686 AND2X1_LOC_126/a_8_24# AND2X1_LOC_42/B 0.00fF
C15687 OR2X1_LOC_424/Y OR2X1_LOC_589/Y 0.07fF
C15688 AND2X1_LOC_663/B OR2X1_LOC_297/A 0.00fF
C15689 AND2X1_LOC_728/Y AND2X1_LOC_192/Y 0.06fF
C15690 OR2X1_LOC_64/Y OR2X1_LOC_597/a_8_216# 0.15fF
C15691 AND2X1_LOC_214/A OR2X1_LOC_52/a_36_216# 0.00fF
C15692 AND2X1_LOC_787/A OR2X1_LOC_437/a_36_216# 0.01fF
C15693 OR2X1_LOC_18/Y OR2X1_LOC_372/Y 0.01fF
C15694 OR2X1_LOC_599/A OR2X1_LOC_433/Y 0.01fF
C15695 AND2X1_LOC_12/Y OR2X1_LOC_793/A 0.11fF
C15696 OR2X1_LOC_160/B OR2X1_LOC_706/B 0.01fF
C15697 AND2X1_LOC_449/Y AND2X1_LOC_453/a_36_24# 0.01fF
C15698 AND2X1_LOC_720/a_8_24# OR2X1_LOC_251/Y 0.01fF
C15699 OR2X1_LOC_36/Y OR2X1_LOC_39/A 0.82fF
C15700 AND2X1_LOC_181/Y AND2X1_LOC_851/B 0.07fF
C15701 OR2X1_LOC_413/a_8_216# OR2X1_LOC_52/B 0.03fF
C15702 OR2X1_LOC_865/B OR2X1_LOC_287/B 0.00fF
C15703 OR2X1_LOC_756/B OR2X1_LOC_456/A 0.00fF
C15704 AND2X1_LOC_578/A AND2X1_LOC_840/a_8_24# 0.03fF
C15705 OR2X1_LOC_629/Y OR2X1_LOC_296/Y 0.75fF
C15706 OR2X1_LOC_630/a_8_216# OR2X1_LOC_296/a_8_216# 0.47fF
C15707 AND2X1_LOC_409/B AND2X1_LOC_409/a_8_24# 0.03fF
C15708 AND2X1_LOC_663/B OR2X1_LOC_275/Y 0.01fF
C15709 AND2X1_LOC_147/a_36_24# OR2X1_LOC_74/A 0.01fF
C15710 VDD OR2X1_LOC_288/A 0.12fF
C15711 AND2X1_LOC_139/B AND2X1_LOC_361/A 0.02fF
C15712 AND2X1_LOC_59/Y AND2X1_LOC_81/a_8_24# 0.06fF
C15713 OR2X1_LOC_600/A OR2X1_LOC_751/A 0.01fF
C15714 OR2X1_LOC_26/Y OR2X1_LOC_767/a_8_216# 0.14fF
C15715 OR2X1_LOC_11/Y AND2X1_LOC_637/Y 0.01fF
C15716 AND2X1_LOC_190/a_8_24# OR2X1_LOC_417/A 0.03fF
C15717 OR2X1_LOC_52/B OR2X1_LOC_265/Y 0.07fF
C15718 OR2X1_LOC_291/Y AND2X1_LOC_647/a_36_24# 0.01fF
C15719 AND2X1_LOC_702/Y AND2X1_LOC_354/B 0.06fF
C15720 OR2X1_LOC_824/Y OR2X1_LOC_6/A 0.16fF
C15721 AND2X1_LOC_196/a_8_24# OR2X1_LOC_48/B 0.01fF
C15722 AND2X1_LOC_70/Y AND2X1_LOC_47/Y 3.37fF
C15723 OR2X1_LOC_744/A OR2X1_LOC_813/A 0.03fF
C15724 OR2X1_LOC_121/Y OR2X1_LOC_66/a_36_216# 0.01fF
C15725 OR2X1_LOC_768/A OR2X1_LOC_532/B 0.01fF
C15726 OR2X1_LOC_89/A OR2X1_LOC_767/a_8_216# 0.05fF
C15727 OR2X1_LOC_404/Y OR2X1_LOC_523/Y 0.14fF
C15728 OR2X1_LOC_774/Y OR2X1_LOC_866/a_8_216# 0.01fF
C15729 AND2X1_LOC_58/a_8_24# OR2X1_LOC_750/A 0.00fF
C15730 OR2X1_LOC_154/A AND2X1_LOC_3/Y 0.26fF
C15731 OR2X1_LOC_61/Y OR2X1_LOC_206/A 0.11fF
C15732 AND2X1_LOC_84/Y AND2X1_LOC_206/Y 0.01fF
C15733 AND2X1_LOC_811/a_8_24# OR2X1_LOC_74/A 0.04fF
C15734 AND2X1_LOC_211/B OR2X1_LOC_36/Y 0.07fF
C15735 OR2X1_LOC_304/a_8_216# OR2X1_LOC_172/Y 0.18fF
C15736 OR2X1_LOC_40/Y AND2X1_LOC_803/a_36_24# 0.01fF
C15737 AND2X1_LOC_211/B OR2X1_LOC_91/a_8_216# 0.11fF
C15738 OR2X1_LOC_112/B OR2X1_LOC_66/A 0.20fF
C15739 AND2X1_LOC_99/A OR2X1_LOC_64/Y 0.12fF
C15740 OR2X1_LOC_18/Y OR2X1_LOC_762/a_8_216# 0.04fF
C15741 OR2X1_LOC_844/Y OR2X1_LOC_560/a_8_216# 0.41fF
C15742 OR2X1_LOC_160/A OR2X1_LOC_206/a_36_216# 0.00fF
C15743 OR2X1_LOC_291/a_8_216# OR2X1_LOC_278/A 0.01fF
C15744 OR2X1_LOC_160/A AND2X1_LOC_51/Y 0.30fF
C15745 OR2X1_LOC_703/A AND2X1_LOC_47/Y 0.03fF
C15746 VDD OR2X1_LOC_3/B 0.00fF
C15747 OR2X1_LOC_607/A OR2X1_LOC_67/Y 0.03fF
C15748 AND2X1_LOC_11/a_36_24# D_INPUT_4 0.01fF
C15749 OR2X1_LOC_851/A OR2X1_LOC_814/A 0.02fF
C15750 OR2X1_LOC_609/A OR2X1_LOC_612/B 1.33fF
C15751 OR2X1_LOC_847/A OR2X1_LOC_54/Y 0.00fF
C15752 OR2X1_LOC_527/Y OR2X1_LOC_406/a_8_216# 0.01fF
C15753 AND2X1_LOC_41/A OR2X1_LOC_241/Y 0.26fF
C15754 OR2X1_LOC_318/A OR2X1_LOC_68/B 0.01fF
C15755 OR2X1_LOC_17/Y OR2X1_LOC_44/Y 0.00fF
C15756 AND2X1_LOC_517/a_36_24# OR2X1_LOC_121/B 0.00fF
C15757 OR2X1_LOC_485/Y OR2X1_LOC_419/Y 0.14fF
C15758 AND2X1_LOC_722/A AND2X1_LOC_810/Y 0.07fF
C15759 OR2X1_LOC_377/A OR2X1_LOC_750/A 0.02fF
C15760 VDD AND2X1_LOC_72/B 0.48fF
C15761 OR2X1_LOC_140/B OR2X1_LOC_777/B 0.03fF
C15762 VDD OR2X1_LOC_451/B 0.21fF
C15763 OR2X1_LOC_3/Y OR2X1_LOC_665/Y 0.02fF
C15764 AND2X1_LOC_50/Y OR2X1_LOC_651/A 0.05fF
C15765 OR2X1_LOC_446/a_36_216# OR2X1_LOC_155/A 0.01fF
C15766 AND2X1_LOC_391/a_8_24# D_INPUT_3 0.05fF
C15767 OR2X1_LOC_235/B D_INPUT_1 1.10fF
C15768 AND2X1_LOC_44/Y OR2X1_LOC_446/B 0.03fF
C15769 OR2X1_LOC_306/Y OR2X1_LOC_22/Y 0.03fF
C15770 OR2X1_LOC_151/A OR2X1_LOC_68/B 0.10fF
C15771 OR2X1_LOC_43/A AND2X1_LOC_663/B 0.15fF
C15772 OR2X1_LOC_3/Y OR2X1_LOC_485/A 0.04fF
C15773 AND2X1_LOC_59/Y AND2X1_LOC_519/a_8_24# 0.01fF
C15774 OR2X1_LOC_366/B OR2X1_LOC_580/A 0.02fF
C15775 OR2X1_LOC_497/Y AND2X1_LOC_844/a_8_24# 0.04fF
C15776 OR2X1_LOC_32/B INPUT_1 0.24fF
C15777 AND2X1_LOC_70/Y OR2X1_LOC_598/A 1.43fF
C15778 OR2X1_LOC_64/Y AND2X1_LOC_637/Y 0.03fF
C15779 OR2X1_LOC_778/A AND2X1_LOC_3/Y 0.03fF
C15780 OR2X1_LOC_791/B OR2X1_LOC_287/a_36_216# 0.00fF
C15781 OR2X1_LOC_325/B OR2X1_LOC_566/a_8_216# 0.06fF
C15782 OR2X1_LOC_22/Y OR2X1_LOC_80/Y 0.01fF
C15783 OR2X1_LOC_3/Y AND2X1_LOC_348/a_8_24# 0.01fF
C15784 OR2X1_LOC_18/Y AND2X1_LOC_660/a_8_24# -0.05fF
C15785 OR2X1_LOC_296/Y OR2X1_LOC_629/a_36_216# 0.00fF
C15786 OR2X1_LOC_375/A AND2X1_LOC_7/Y 0.04fF
C15787 OR2X1_LOC_42/a_8_216# OR2X1_LOC_46/A 0.01fF
C15788 OR2X1_LOC_204/Y OR2X1_LOC_814/A 0.03fF
C15789 AND2X1_LOC_486/Y OR2X1_LOC_47/Y 0.03fF
C15790 OR2X1_LOC_619/a_8_216# AND2X1_LOC_852/B 0.03fF
C15791 OR2X1_LOC_676/Y AND2X1_LOC_31/Y 0.07fF
C15792 OR2X1_LOC_485/Y OR2X1_LOC_526/a_8_216# 0.39fF
C15793 OR2X1_LOC_688/Y AND2X1_LOC_689/a_8_24# 0.23fF
C15794 AND2X1_LOC_721/a_8_24# AND2X1_LOC_721/A -0.00fF
C15795 OR2X1_LOC_127/a_8_216# D_INPUT_3 0.02fF
C15796 OR2X1_LOC_624/B AND2X1_LOC_51/Y 0.01fF
C15797 AND2X1_LOC_51/Y OR2X1_LOC_33/a_8_216# 0.01fF
C15798 OR2X1_LOC_502/A OR2X1_LOC_330/a_36_216# 0.02fF
C15799 OR2X1_LOC_91/Y AND2X1_LOC_675/A 0.32fF
C15800 AND2X1_LOC_784/A D_INPUT_0 0.08fF
C15801 OR2X1_LOC_160/A OR2X1_LOC_201/a_36_216# 0.03fF
C15802 OR2X1_LOC_834/A AND2X1_LOC_31/Y 0.01fF
C15803 OR2X1_LOC_22/Y AND2X1_LOC_857/a_36_24# -0.01fF
C15804 OR2X1_LOC_19/B AND2X1_LOC_822/a_36_24# 0.00fF
C15805 OR2X1_LOC_616/a_36_216# GATE_662 0.00fF
C15806 OR2X1_LOC_43/A OR2X1_LOC_54/a_8_216# 0.04fF
C15807 AND2X1_LOC_702/Y AND2X1_LOC_863/Y 0.01fF
C15808 OR2X1_LOC_95/Y OR2X1_LOC_6/A 0.06fF
C15809 OR2X1_LOC_368/A OR2X1_LOC_6/A 0.01fF
C15810 OR2X1_LOC_539/B OR2X1_LOC_390/A 0.04fF
C15811 D_INPUT_0 OR2X1_LOC_37/a_8_216# 0.02fF
C15812 AND2X1_LOC_17/Y AND2X1_LOC_47/Y 0.08fF
C15813 AND2X1_LOC_76/Y AND2X1_LOC_205/a_8_24# 0.01fF
C15814 OR2X1_LOC_416/A OR2X1_LOC_49/a_8_216# 0.47fF
C15815 AND2X1_LOC_835/a_8_24# AND2X1_LOC_240/Y 0.06fF
C15816 AND2X1_LOC_91/B OR2X1_LOC_554/a_8_216# 0.27fF
C15817 INPUT_1 OR2X1_LOC_371/Y 0.38fF
C15818 OR2X1_LOC_86/A OR2X1_LOC_278/Y 0.01fF
C15819 AND2X1_LOC_582/a_8_24# AND2X1_LOC_430/B 0.01fF
C15820 OR2X1_LOC_599/A OR2X1_LOC_760/Y 0.01fF
C15821 AND2X1_LOC_856/B AND2X1_LOC_863/A 0.05fF
C15822 OR2X1_LOC_811/A OR2X1_LOC_675/Y 2.04fF
C15823 OR2X1_LOC_61/B OR2X1_LOC_228/Y 0.06fF
C15824 AND2X1_LOC_259/Y AND2X1_LOC_866/A 0.05fF
C15825 AND2X1_LOC_140/a_8_24# OR2X1_LOC_71/Y 0.01fF
C15826 OR2X1_LOC_47/Y OR2X1_LOC_248/Y 0.70fF
C15827 AND2X1_LOC_191/B OR2X1_LOC_13/B 0.07fF
C15828 OR2X1_LOC_44/Y OR2X1_LOC_588/A 0.00fF
C15829 OR2X1_LOC_687/a_8_216# AND2X1_LOC_425/Y 0.01fF
C15830 AND2X1_LOC_465/a_8_24# OR2X1_LOC_95/Y 0.01fF
C15831 OR2X1_LOC_419/Y OR2X1_LOC_39/A 0.11fF
C15832 AND2X1_LOC_213/B AND2X1_LOC_783/B 0.10fF
C15833 OR2X1_LOC_216/Y OR2X1_LOC_205/Y 0.07fF
C15834 OR2X1_LOC_417/a_8_216# OR2X1_LOC_417/A 0.02fF
C15835 OR2X1_LOC_478/Y OR2X1_LOC_480/a_8_216# 0.39fF
C15836 AND2X1_LOC_684/a_8_24# AND2X1_LOC_3/Y 0.02fF
C15837 OR2X1_LOC_436/a_36_216# OR2X1_LOC_814/A 0.01fF
C15838 AND2X1_LOC_792/Y OR2X1_LOC_44/Y 0.01fF
C15839 OR2X1_LOC_74/A AND2X1_LOC_440/a_36_24# 0.01fF
C15840 OR2X1_LOC_280/Y OR2X1_LOC_224/a_36_216# 0.02fF
C15841 VDD AND2X1_LOC_36/Y 1.73fF
C15842 OR2X1_LOC_160/B OR2X1_LOC_844/B 0.06fF
C15843 AND2X1_LOC_564/B AND2X1_LOC_795/a_8_24# 0.02fF
C15844 OR2X1_LOC_47/Y AND2X1_LOC_294/a_36_24# 0.00fF
C15845 OR2X1_LOC_527/Y AND2X1_LOC_675/A 0.02fF
C15846 OR2X1_LOC_631/B OR2X1_LOC_247/a_36_216# 0.01fF
C15847 OR2X1_LOC_404/Y AND2X1_LOC_47/Y 0.04fF
C15848 AND2X1_LOC_840/B OR2X1_LOC_406/A 0.45fF
C15849 VDD OR2X1_LOC_759/Y 0.12fF
C15850 GATE_366 AND2X1_LOC_848/A 2.01fF
C15851 AND2X1_LOC_92/Y OR2X1_LOC_593/B 0.03fF
C15852 OR2X1_LOC_116/a_8_216# OR2X1_LOC_598/A -0.01fF
C15853 OR2X1_LOC_269/B OR2X1_LOC_374/Y 4.83fF
C15854 OR2X1_LOC_416/Y AND2X1_LOC_293/a_8_24# 0.01fF
C15855 OR2X1_LOC_52/B AND2X1_LOC_205/a_8_24# 0.01fF
C15856 OR2X1_LOC_721/Y OR2X1_LOC_140/Y 0.34fF
C15857 OR2X1_LOC_518/a_8_216# AND2X1_LOC_715/A 0.47fF
C15858 VDD OR2X1_LOC_333/a_8_216# 0.21fF
C15859 OR2X1_LOC_287/B OR2X1_LOC_493/Y 0.03fF
C15860 AND2X1_LOC_841/B OR2X1_LOC_589/Y 0.01fF
C15861 AND2X1_LOC_832/a_36_24# OR2X1_LOC_423/Y 0.00fF
C15862 OR2X1_LOC_86/a_36_216# AND2X1_LOC_647/Y 0.00fF
C15863 OR2X1_LOC_419/Y OR2X1_LOC_239/a_36_216# 0.00fF
C15864 AND2X1_LOC_387/B OR2X1_LOC_644/A 0.03fF
C15865 OR2X1_LOC_685/a_8_216# AND2X1_LOC_430/B 0.01fF
C15866 VDD OR2X1_LOC_767/Y 0.12fF
C15867 OR2X1_LOC_256/Y OR2X1_LOC_248/A 0.01fF
C15868 AND2X1_LOC_388/Y AND2X1_LOC_802/B 0.01fF
C15869 OR2X1_LOC_696/A OR2X1_LOC_585/Y 0.04fF
C15870 AND2X1_LOC_57/Y OR2X1_LOC_35/Y 0.01fF
C15871 OR2X1_LOC_74/A AND2X1_LOC_204/Y 0.21fF
C15872 OR2X1_LOC_175/Y OR2X1_LOC_648/B 0.10fF
C15873 OR2X1_LOC_481/A AND2X1_LOC_721/A 0.00fF
C15874 AND2X1_LOC_576/Y AND2X1_LOC_657/A 0.01fF
C15875 OR2X1_LOC_528/Y AND2X1_LOC_721/Y 0.06fF
C15876 OR2X1_LOC_147/B OR2X1_LOC_181/Y 0.05fF
C15877 OR2X1_LOC_829/A OR2X1_LOC_12/Y 0.04fF
C15878 OR2X1_LOC_719/A AND2X1_LOC_237/a_8_24# 0.21fF
C15879 OR2X1_LOC_691/Y OR2X1_LOC_648/B 0.01fF
C15880 AND2X1_LOC_273/a_8_24# AND2X1_LOC_92/Y 0.06fF
C15881 AND2X1_LOC_97/a_36_24# OR2X1_LOC_13/B 0.00fF
C15882 OR2X1_LOC_49/A OR2X1_LOC_159/a_8_216# 0.04fF
C15883 AND2X1_LOC_141/a_36_24# AND2X1_LOC_772/Y 0.01fF
C15884 OR2X1_LOC_293/a_36_216# D_INPUT_1 0.03fF
C15885 OR2X1_LOC_223/A OR2X1_LOC_335/B 0.00fF
C15886 OR2X1_LOC_62/A D_INPUT_0 0.11fF
C15887 OR2X1_LOC_7/A AND2X1_LOC_563/Y 0.00fF
C15888 OR2X1_LOC_721/a_8_216# AND2X1_LOC_18/Y 0.01fF
C15889 OR2X1_LOC_375/A OR2X1_LOC_140/Y 0.03fF
C15890 OR2X1_LOC_154/a_8_216# VDD 0.00fF
C15891 AND2X1_LOC_64/Y OR2X1_LOC_630/B 0.00fF
C15892 OR2X1_LOC_739/A OR2X1_LOC_532/a_36_216# 0.00fF
C15893 AND2X1_LOC_3/Y OR2X1_LOC_560/A 0.06fF
C15894 OR2X1_LOC_502/A AND2X1_LOC_409/B 0.09fF
C15895 AND2X1_LOC_3/Y OR2X1_LOC_198/A 0.02fF
C15896 OR2X1_LOC_542/B AND2X1_LOC_44/Y 0.03fF
C15897 AND2X1_LOC_56/B OR2X1_LOC_317/B 0.00fF
C15898 OR2X1_LOC_62/B OR2X1_LOC_84/a_36_216# 0.00fF
C15899 OR2X1_LOC_852/A AND2X1_LOC_827/a_8_24# 0.23fF
C15900 OR2X1_LOC_19/B OR2X1_LOC_86/A 0.01fF
C15901 OR2X1_LOC_506/Y VDD 0.00fF
C15902 OR2X1_LOC_502/A AND2X1_LOC_763/B 0.01fF
C15903 OR2X1_LOC_719/B OR2X1_LOC_719/a_8_216# 0.02fF
C15904 OR2X1_LOC_615/a_36_216# OR2X1_LOC_753/Y 0.00fF
C15905 OR2X1_LOC_272/Y AND2X1_LOC_216/a_8_24# 0.24fF
C15906 VDD OR2X1_LOC_584/a_8_216# 0.21fF
C15907 OR2X1_LOC_753/A OR2X1_LOC_150/a_36_216# 0.00fF
C15908 OR2X1_LOC_671/Y INPUT_2 0.02fF
C15909 OR2X1_LOC_9/Y OR2X1_LOC_6/B 0.18fF
C15910 OR2X1_LOC_230/a_8_216# OR2X1_LOC_172/Y 0.04fF
C15911 AND2X1_LOC_92/Y AND2X1_LOC_256/a_8_24# 0.01fF
C15912 OR2X1_LOC_575/A OR2X1_LOC_140/B 0.03fF
C15913 OR2X1_LOC_437/a_36_216# AND2X1_LOC_675/A 0.00fF
C15914 OR2X1_LOC_235/B OR2X1_LOC_15/a_8_216# 0.01fF
C15915 OR2X1_LOC_91/A AND2X1_LOC_774/A 0.22fF
C15916 OR2X1_LOC_276/B D_INPUT_1 0.07fF
C15917 OR2X1_LOC_604/A OR2X1_LOC_485/Y 0.09fF
C15918 OR2X1_LOC_78/B OR2X1_LOC_390/A 0.03fF
C15919 OR2X1_LOC_52/B AND2X1_LOC_449/a_8_24# 0.02fF
C15920 VDD AND2X1_LOC_535/Y 0.01fF
C15921 OR2X1_LOC_705/Y OR2X1_LOC_725/a_8_216# 0.01fF
C15922 OR2X1_LOC_756/B OR2X1_LOC_161/B 0.55fF
C15923 OR2X1_LOC_756/B OR2X1_LOC_562/B 0.00fF
C15924 OR2X1_LOC_736/A AND2X1_LOC_44/Y 1.03fF
C15925 INPUT_1 AND2X1_LOC_222/Y 0.01fF
C15926 OR2X1_LOC_494/Y AND2X1_LOC_860/A 0.10fF
C15927 OR2X1_LOC_160/B OR2X1_LOC_389/A 0.01fF
C15928 AND2X1_LOC_363/Y AND2X1_LOC_860/A 0.03fF
C15929 AND2X1_LOC_81/B OR2X1_LOC_502/a_8_216# 0.01fF
C15930 OR2X1_LOC_47/Y AND2X1_LOC_646/a_8_24# 0.17fF
C15931 OR2X1_LOC_18/Y AND2X1_LOC_773/a_8_24# 0.06fF
C15932 OR2X1_LOC_39/A OR2X1_LOC_19/a_8_216# 0.06fF
C15933 AND2X1_LOC_392/A AND2X1_LOC_337/a_8_24# 0.02fF
C15934 AND2X1_LOC_112/a_8_24# AND2X1_LOC_715/A 0.00fF
C15935 OR2X1_LOC_479/Y OR2X1_LOC_716/a_8_216# 0.02fF
C15936 AND2X1_LOC_571/A OR2X1_LOC_91/Y 0.05fF
C15937 AND2X1_LOC_738/B OR2X1_LOC_600/A 0.13fF
C15938 D_INPUT_0 OR2X1_LOC_88/Y 0.03fF
C15939 INPUT_1 OR2X1_LOC_68/B 0.35fF
C15940 OR2X1_LOC_600/A OR2X1_LOC_56/A 6.28fF
C15941 AND2X1_LOC_335/Y OR2X1_LOC_56/A 0.02fF
C15942 AND2X1_LOC_514/Y AND2X1_LOC_212/a_8_24# 0.04fF
C15943 OR2X1_LOC_40/Y OR2X1_LOC_310/Y 0.01fF
C15944 OR2X1_LOC_624/A OR2X1_LOC_474/B 0.02fF
C15945 AND2X1_LOC_773/Y OR2X1_LOC_48/B 0.05fF
C15946 OR2X1_LOC_600/A OR2X1_LOC_819/a_8_216# 0.01fF
C15947 VDD OR2X1_LOC_630/Y 0.37fF
C15948 OR2X1_LOC_71/Y AND2X1_LOC_217/a_8_24# 0.01fF
C15949 AND2X1_LOC_511/a_8_24# OR2X1_LOC_502/A 0.01fF
C15950 OR2X1_LOC_639/B AND2X1_LOC_7/B 0.02fF
C15951 OR2X1_LOC_40/Y OR2X1_LOC_441/a_8_216# 0.03fF
C15952 AND2X1_LOC_658/A AND2X1_LOC_663/A 0.03fF
C15953 OR2X1_LOC_56/A AND2X1_LOC_296/a_8_24# 0.01fF
C15954 AND2X1_LOC_51/Y OR2X1_LOC_532/Y 0.01fF
C15955 OR2X1_LOC_6/B OR2X1_LOC_474/Y 0.07fF
C15956 AND2X1_LOC_675/Y AND2X1_LOC_188/a_8_24# 0.05fF
C15957 OR2X1_LOC_837/B AND2X1_LOC_415/a_36_24# 0.00fF
C15958 AND2X1_LOC_392/A OR2X1_LOC_275/Y 0.03fF
C15959 OR2X1_LOC_375/A OR2X1_LOC_375/a_8_216# 0.02fF
C15960 AND2X1_LOC_710/Y AND2X1_LOC_711/a_8_24# 0.01fF
C15961 OR2X1_LOC_715/B OR2X1_LOC_623/B 0.07fF
C15962 OR2X1_LOC_158/A OR2X1_LOC_689/a_8_216# 0.01fF
C15963 AND2X1_LOC_553/a_8_24# OR2X1_LOC_103/Y 0.01fF
C15964 OR2X1_LOC_709/A OR2X1_LOC_506/A 0.03fF
C15965 D_GATE_479 OR2X1_LOC_453/a_8_216# 0.02fF
C15966 OR2X1_LOC_426/A OR2X1_LOC_581/Y 0.34fF
C15967 OR2X1_LOC_375/A OR2X1_LOC_706/a_8_216# 0.01fF
C15968 AND2X1_LOC_287/B OR2X1_LOC_44/Y 0.00fF
C15969 OR2X1_LOC_36/Y AND2X1_LOC_456/a_8_24# 0.04fF
C15970 OR2X1_LOC_166/Y AND2X1_LOC_436/a_8_24# 0.01fF
C15971 AND2X1_LOC_477/Y AND2X1_LOC_808/a_8_24# 0.01fF
C15972 AND2X1_LOC_564/B OR2X1_LOC_496/Y 0.02fF
C15973 OR2X1_LOC_264/Y AND2X1_LOC_18/Y 0.22fF
C15974 AND2X1_LOC_284/a_8_24# AND2X1_LOC_806/A 0.01fF
C15975 OR2X1_LOC_453/a_8_216# OR2X1_LOC_161/B 0.01fF
C15976 AND2X1_LOC_719/Y OR2X1_LOC_278/Y 0.01fF
C15977 OR2X1_LOC_314/Y OR2X1_LOC_16/A 0.05fF
C15978 OR2X1_LOC_49/A OR2X1_LOC_618/a_8_216# 0.18fF
C15979 OR2X1_LOC_816/A OR2X1_LOC_44/Y 0.03fF
C15980 OR2X1_LOC_185/Y AND2X1_LOC_522/a_8_24# 0.28fF
C15981 AND2X1_LOC_56/B AND2X1_LOC_44/Y 0.47fF
C15982 OR2X1_LOC_149/a_8_216# OR2X1_LOC_161/A 0.01fF
C15983 OR2X1_LOC_177/Y OR2X1_LOC_39/A 0.05fF
C15984 AND2X1_LOC_513/a_36_24# OR2X1_LOC_51/Y 0.00fF
C15985 OR2X1_LOC_657/a_8_216# OR2X1_LOC_161/B 0.01fF
C15986 OR2X1_LOC_40/Y AND2X1_LOC_805/Y 0.04fF
C15987 OR2X1_LOC_92/Y AND2X1_LOC_285/Y 0.02fF
C15988 OR2X1_LOC_519/a_8_216# OR2X1_LOC_40/Y 0.01fF
C15989 OR2X1_LOC_840/A OR2X1_LOC_648/A 0.10fF
C15990 AND2X1_LOC_51/Y OR2X1_LOC_130/Y 0.13fF
C15991 OR2X1_LOC_545/B OR2X1_LOC_181/Y 0.17fF
C15992 AND2X1_LOC_723/a_36_24# OR2X1_LOC_40/Y 0.00fF
C15993 OR2X1_LOC_45/B AND2X1_LOC_853/Y 0.01fF
C15994 AND2X1_LOC_8/Y AND2X1_LOC_44/Y 0.29fF
C15995 OR2X1_LOC_18/Y AND2X1_LOC_243/Y 0.10fF
C15996 AND2X1_LOC_125/a_36_24# OR2X1_LOC_66/A 0.00fF
C15997 OR2X1_LOC_821/Y OR2X1_LOC_6/A 0.02fF
C15998 AND2X1_LOC_712/a_8_24# OR2X1_LOC_52/B 0.02fF
C15999 AND2X1_LOC_572/a_36_24# OR2X1_LOC_89/A -0.00fF
C16000 AND2X1_LOC_217/Y OR2X1_LOC_118/Y 0.01fF
C16001 OR2X1_LOC_538/A AND2X1_LOC_167/a_36_24# 0.00fF
C16002 OR2X1_LOC_756/B OR2X1_LOC_435/B 0.09fF
C16003 AND2X1_LOC_64/Y AND2X1_LOC_67/Y 0.02fF
C16004 OR2X1_LOC_471/Y OR2X1_LOC_726/a_8_216# 0.04fF
C16005 OR2X1_LOC_641/A OR2X1_LOC_340/Y 1.22fF
C16006 OR2X1_LOC_116/A OR2X1_LOC_6/B 0.05fF
C16007 OR2X1_LOC_333/B AND2X1_LOC_7/B 0.03fF
C16008 AND2X1_LOC_56/B OR2X1_LOC_514/a_8_216# 0.02fF
C16009 AND2X1_LOC_116/Y AND2X1_LOC_473/Y 0.09fF
C16010 AND2X1_LOC_586/a_8_24# VDD -0.00fF
C16011 OR2X1_LOC_216/A AND2X1_LOC_41/A 0.03fF
C16012 AND2X1_LOC_70/Y AND2X1_LOC_682/a_8_24# 0.01fF
C16013 AND2X1_LOC_21/Y AND2X1_LOC_44/Y 0.02fF
C16014 AND2X1_LOC_292/a_8_24# OR2X1_LOC_294/Y 0.01fF
C16015 OR2X1_LOC_604/A OR2X1_LOC_39/A 0.42fF
C16016 OR2X1_LOC_329/B AND2X1_LOC_851/A 0.03fF
C16017 OR2X1_LOC_130/A OR2X1_LOC_641/A 0.07fF
C16018 OR2X1_LOC_599/A AND2X1_LOC_714/B 0.00fF
C16019 AND2X1_LOC_392/A AND2X1_LOC_365/A 0.02fF
C16020 OR2X1_LOC_579/B OR2X1_LOC_362/A 0.03fF
C16021 OR2X1_LOC_697/a_8_216# OR2X1_LOC_422/a_8_216# 0.47fF
C16022 OR2X1_LOC_87/A OR2X1_LOC_180/a_8_216# 0.01fF
C16023 OR2X1_LOC_140/A OR2X1_LOC_510/Y 0.03fF
C16024 OR2X1_LOC_427/A OR2X1_LOC_59/Y 0.35fF
C16025 AND2X1_LOC_70/Y OR2X1_LOC_506/A 0.02fF
C16026 OR2X1_LOC_507/A OR2X1_LOC_510/Y 0.09fF
C16027 INPUT_4 OR2X1_LOC_581/Y 0.01fF
C16028 AND2X1_LOC_192/Y AND2X1_LOC_480/A 0.08fF
C16029 OR2X1_LOC_369/Y OR2X1_LOC_109/Y 0.01fF
C16030 OR2X1_LOC_6/B OR2X1_LOC_217/Y 0.03fF
C16031 OR2X1_LOC_6/B OR2X1_LOC_96/B 0.03fF
C16032 AND2X1_LOC_48/A AND2X1_LOC_763/B 0.04fF
C16033 OR2X1_LOC_619/Y OR2X1_LOC_56/A 0.16fF
C16034 OR2X1_LOC_158/A OR2X1_LOC_26/Y 0.42fF
C16035 OR2X1_LOC_215/A OR2X1_LOC_392/B 0.08fF
C16036 OR2X1_LOC_467/B OR2X1_LOC_210/B 0.16fF
C16037 AND2X1_LOC_356/a_8_24# OR2X1_LOC_56/A 0.03fF
C16038 OR2X1_LOC_19/B OR2X1_LOC_20/A 0.01fF
C16039 OR2X1_LOC_756/B OR2X1_LOC_61/Y 0.01fF
C16040 OR2X1_LOC_123/a_8_216# OR2X1_LOC_375/A 0.01fF
C16041 OR2X1_LOC_508/A OR2X1_LOC_216/A 0.03fF
C16042 AND2X1_LOC_639/a_36_24# OR2X1_LOC_428/A 0.00fF
C16043 OR2X1_LOC_402/B OR2X1_LOC_402/Y 0.17fF
C16044 AND2X1_LOC_388/a_8_24# AND2X1_LOC_436/Y 0.02fF
C16045 VDD OR2X1_LOC_246/Y 0.03fF
C16046 OR2X1_LOC_40/Y AND2X1_LOC_661/A 0.03fF
C16047 AND2X1_LOC_784/A AND2X1_LOC_784/a_8_24# 0.01fF
C16048 OR2X1_LOC_99/B AND2X1_LOC_7/B 0.02fF
C16049 AND2X1_LOC_95/Y OR2X1_LOC_235/B 0.03fF
C16050 AND2X1_LOC_95/a_8_24# AND2X1_LOC_25/Y 0.01fF
C16051 VDD AND2X1_LOC_576/Y 0.02fF
C16052 OR2X1_LOC_158/A OR2X1_LOC_89/A 0.36fF
C16053 OR2X1_LOC_666/a_8_216# AND2X1_LOC_859/Y 0.03fF
C16054 AND2X1_LOC_392/A OR2X1_LOC_43/A 0.01fF
C16055 AND2X1_LOC_597/a_8_24# OR2X1_LOC_676/Y 0.04fF
C16056 OR2X1_LOC_643/A AND2X1_LOC_18/Y 0.15fF
C16057 OR2X1_LOC_538/A OR2X1_LOC_212/A 0.00fF
C16058 AND2X1_LOC_523/Y OR2X1_LOC_428/A 0.06fF
C16059 AND2X1_LOC_509/Y AND2X1_LOC_474/a_8_24# 0.20fF
C16060 OR2X1_LOC_805/A OR2X1_LOC_778/B 0.15fF
C16061 VDD OR2X1_LOC_687/B -0.00fF
C16062 OR2X1_LOC_744/A AND2X1_LOC_435/a_36_24# 0.00fF
C16063 AND2X1_LOC_712/Y OR2X1_LOC_7/A 0.01fF
C16064 OR2X1_LOC_485/A AND2X1_LOC_477/Y 0.14fF
C16065 AND2X1_LOC_784/A AND2X1_LOC_326/B 0.05fF
C16066 OR2X1_LOC_479/Y AND2X1_LOC_300/a_8_24# 0.02fF
C16067 OR2X1_LOC_650/a_36_216# OR2X1_LOC_462/B 0.00fF
C16068 OR2X1_LOC_641/Y OR2X1_LOC_649/B 0.01fF
C16069 VDD OR2X1_LOC_346/B 0.21fF
C16070 OR2X1_LOC_154/A INPUT_0 0.35fF
C16071 AND2X1_LOC_675/Y AND2X1_LOC_186/a_36_24# 0.01fF
C16072 OR2X1_LOC_389/A OR2X1_LOC_219/B 0.08fF
C16073 OR2X1_LOC_371/Y AND2X1_LOC_778/Y 0.00fF
C16074 OR2X1_LOC_542/B OR2X1_LOC_465/B 0.03fF
C16075 AND2X1_LOC_521/a_8_24# OR2X1_LOC_404/Y 0.01fF
C16076 OR2X1_LOC_97/B OR2X1_LOC_78/A 0.08fF
C16077 OR2X1_LOC_482/Y AND2X1_LOC_483/a_8_24# 0.00fF
C16078 OR2X1_LOC_604/A OR2X1_LOC_429/Y 0.23fF
C16079 AND2X1_LOC_486/Y OR2X1_LOC_625/Y 0.33fF
C16080 AND2X1_LOC_677/a_8_24# OR2X1_LOC_161/B 0.04fF
C16081 OR2X1_LOC_147/B OR2X1_LOC_220/B 0.14fF
C16082 OR2X1_LOC_574/A OR2X1_LOC_66/A 0.03fF
C16083 OR2X1_LOC_181/B OR2X1_LOC_540/a_36_216# 0.03fF
C16084 AND2X1_LOC_474/A OR2X1_LOC_36/Y 0.03fF
C16085 AND2X1_LOC_51/Y OR2X1_LOC_768/a_8_216# 0.01fF
C16086 AND2X1_LOC_784/A AND2X1_LOC_471/Y 0.03fF
C16087 OR2X1_LOC_95/Y OR2X1_LOC_184/a_8_216# 0.18fF
C16088 OR2X1_LOC_600/A AND2X1_LOC_641/Y 0.03fF
C16089 OR2X1_LOC_43/A AND2X1_LOC_436/a_8_24# 0.01fF
C16090 AND2X1_LOC_513/a_36_24# OR2X1_LOC_680/A 0.01fF
C16091 OR2X1_LOC_147/A OR2X1_LOC_269/B 0.24fF
C16092 AND2X1_LOC_851/B AND2X1_LOC_455/a_8_24# 0.03fF
C16093 AND2X1_LOC_385/a_8_24# AND2X1_LOC_41/A 0.03fF
C16094 OR2X1_LOC_45/Y OR2X1_LOC_45/a_8_216# 0.03fF
C16095 AND2X1_LOC_332/a_36_24# OR2X1_LOC_46/A 0.01fF
C16096 AND2X1_LOC_511/a_8_24# AND2X1_LOC_48/A 0.03fF
C16097 OR2X1_LOC_838/B OR2X1_LOC_20/A 1.11fF
C16098 OR2X1_LOC_329/B OR2X1_LOC_485/A 0.19fF
C16099 OR2X1_LOC_656/B AND2X1_LOC_59/Y 0.03fF
C16100 AND2X1_LOC_95/a_8_24# AND2X1_LOC_51/Y 0.17fF
C16101 OR2X1_LOC_103/Y OR2X1_LOC_26/Y 0.10fF
C16102 AND2X1_LOC_12/Y OR2X1_LOC_212/A 0.03fF
C16103 AND2X1_LOC_720/Y OR2X1_LOC_26/Y 0.01fF
C16104 OR2X1_LOC_568/A OR2X1_LOC_535/a_8_216# 0.03fF
C16105 OR2X1_LOC_528/Y OR2X1_LOC_628/Y 0.07fF
C16106 OR2X1_LOC_124/A OR2X1_LOC_123/B 0.81fF
C16107 OR2X1_LOC_377/A OR2X1_LOC_243/A 0.00fF
C16108 OR2X1_LOC_379/Y OR2X1_LOC_130/A 0.03fF
C16109 AND2X1_LOC_775/a_8_24# OR2X1_LOC_427/A 0.02fF
C16110 AND2X1_LOC_710/a_8_24# OR2X1_LOC_701/Y 0.00fF
C16111 OR2X1_LOC_62/B OR2X1_LOC_641/A 0.00fF
C16112 OR2X1_LOC_51/Y OR2X1_LOC_52/Y 0.02fF
C16113 AND2X1_LOC_87/a_8_24# OR2X1_LOC_619/Y 0.03fF
C16114 AND2X1_LOC_108/a_8_24# OR2X1_LOC_346/A 0.08fF
C16115 OR2X1_LOC_812/B OR2X1_LOC_561/a_8_216# 0.02fF
C16116 AND2X1_LOC_43/B AND2X1_LOC_272/a_8_24# 0.06fF
C16117 OR2X1_LOC_154/A OR2X1_LOC_732/B 0.10fF
C16118 OR2X1_LOC_45/Y OR2X1_LOC_44/Y 0.08fF
C16119 OR2X1_LOC_103/Y OR2X1_LOC_89/A 0.32fF
C16120 OR2X1_LOC_427/A OR2X1_LOC_820/B 0.02fF
C16121 OR2X1_LOC_685/B OR2X1_LOC_161/A 0.01fF
C16122 AND2X1_LOC_354/Y OR2X1_LOC_43/A 0.02fF
C16123 OR2X1_LOC_47/Y AND2X1_LOC_457/a_8_24# 0.10fF
C16124 AND2X1_LOC_12/Y OR2X1_LOC_687/Y 0.08fF
C16125 OR2X1_LOC_837/B OR2X1_LOC_585/A 0.15fF
C16126 AND2X1_LOC_326/A INPUT_0 0.12fF
C16127 OR2X1_LOC_673/A OR2X1_LOC_633/A 0.04fF
C16128 OR2X1_LOC_113/A AND2X1_LOC_18/Y 0.01fF
C16129 OR2X1_LOC_36/Y AND2X1_LOC_593/Y 0.01fF
C16130 OR2X1_LOC_625/Y OR2X1_LOC_248/Y 0.22fF
C16131 AND2X1_LOC_360/a_8_24# OR2X1_LOC_3/Y 0.01fF
C16132 OR2X1_LOC_377/A OR2X1_LOC_36/Y 5.35fF
C16133 OR2X1_LOC_9/Y AND2X1_LOC_47/Y 0.00fF
C16134 OR2X1_LOC_80/Y OR2X1_LOC_39/A 0.00fF
C16135 OR2X1_LOC_286/Y OR2X1_LOC_269/B 0.01fF
C16136 OR2X1_LOC_516/a_8_216# OR2X1_LOC_680/A 0.02fF
C16137 OR2X1_LOC_422/Y OR2X1_LOC_7/A 0.01fF
C16138 AND2X1_LOC_47/Y OR2X1_LOC_362/A 0.03fF
C16139 OR2X1_LOC_427/A AND2X1_LOC_446/a_36_24# 0.00fF
C16140 AND2X1_LOC_338/Y OR2X1_LOC_289/Y 0.17fF
C16141 AND2X1_LOC_580/B OR2X1_LOC_616/a_8_216# 0.01fF
C16142 AND2X1_LOC_40/Y OR2X1_LOC_592/A 0.01fF
C16143 OR2X1_LOC_515/a_8_216# OR2X1_LOC_515/Y 0.01fF
C16144 OR2X1_LOC_631/B OR2X1_LOC_499/a_8_216# 0.01fF
C16145 AND2X1_LOC_89/a_8_24# OR2X1_LOC_375/A 0.04fF
C16146 OR2X1_LOC_426/B AND2X1_LOC_326/a_36_24# 0.01fF
C16147 OR2X1_LOC_750/A OR2X1_LOC_78/B 0.01fF
C16148 AND2X1_LOC_710/a_8_24# OR2X1_LOC_44/Y 0.01fF
C16149 AND2X1_LOC_476/A AND2X1_LOC_476/Y 0.19fF
C16150 OR2X1_LOC_103/a_8_216# OR2X1_LOC_89/A 0.01fF
C16151 OR2X1_LOC_121/Y OR2X1_LOC_786/Y 0.56fF
C16152 OR2X1_LOC_8/Y D_INPUT_0 0.26fF
C16153 OR2X1_LOC_673/a_8_216# OR2X1_LOC_673/A 0.08fF
C16154 AND2X1_LOC_191/Y OR2X1_LOC_427/A 0.03fF
C16155 OR2X1_LOC_832/a_8_216# AND2X1_LOC_47/Y 0.01fF
C16156 OR2X1_LOC_702/A OR2X1_LOC_856/B 0.03fF
C16157 AND2X1_LOC_808/A AND2X1_LOC_212/Y 0.06fF
C16158 OR2X1_LOC_814/A OR2X1_LOC_78/A 0.15fF
C16159 OR2X1_LOC_36/Y OR2X1_LOC_85/A 0.07fF
C16160 OR2X1_LOC_375/A OR2X1_LOC_710/a_8_216# 0.01fF
C16161 OR2X1_LOC_168/A OR2X1_LOC_78/B 0.02fF
C16162 OR2X1_LOC_400/a_8_216# AND2X1_LOC_51/Y 0.01fF
C16163 AND2X1_LOC_711/Y OR2X1_LOC_427/A 0.03fF
C16164 VDD OR2X1_LOC_780/a_8_216# 0.21fF
C16165 OR2X1_LOC_377/A AND2X1_LOC_822/a_8_24# 0.02fF
C16166 AND2X1_LOC_302/a_36_24# OR2X1_LOC_6/A 0.00fF
C16167 AND2X1_LOC_376/a_8_24# OR2X1_LOC_459/B 0.02fF
C16168 OR2X1_LOC_70/Y OR2X1_LOC_427/A 4.74fF
C16169 AND2X1_LOC_99/a_8_24# AND2X1_LOC_101/a_8_24# 0.23fF
C16170 OR2X1_LOC_417/Y OR2X1_LOC_92/Y 0.07fF
C16171 AND2X1_LOC_644/a_8_24# OR2X1_LOC_16/A 0.01fF
C16172 OR2X1_LOC_850/a_8_216# OR2X1_LOC_814/A 0.01fF
C16173 OR2X1_LOC_291/A OR2X1_LOC_619/Y 0.40fF
C16174 OR2X1_LOC_574/A OR2X1_LOC_799/a_36_216# 0.16fF
C16175 AND2X1_LOC_367/A INPUT_1 0.10fF
C16176 OR2X1_LOC_591/a_8_216# OR2X1_LOC_44/Y 0.02fF
C16177 AND2X1_LOC_395/a_8_24# AND2X1_LOC_3/Y 0.02fF
C16178 OR2X1_LOC_357/a_36_216# OR2X1_LOC_365/B 0.00fF
C16179 OR2X1_LOC_462/B OR2X1_LOC_240/A 0.24fF
C16180 OR2X1_LOC_311/Y OR2X1_LOC_92/Y 0.03fF
C16181 AND2X1_LOC_722/A AND2X1_LOC_477/A 0.03fF
C16182 OR2X1_LOC_847/A AND2X1_LOC_51/Y 0.00fF
C16183 OR2X1_LOC_97/A OR2X1_LOC_228/Y 0.02fF
C16184 OR2X1_LOC_447/A AND2X1_LOC_51/Y 0.01fF
C16185 OR2X1_LOC_599/A AND2X1_LOC_645/A 0.03fF
C16186 AND2X1_LOC_302/a_8_24# OR2X1_LOC_299/Y 0.01fF
C16187 VDD OR2X1_LOC_269/Y 0.12fF
C16188 OR2X1_LOC_669/a_8_216# OR2X1_LOC_669/Y 0.01fF
C16189 OR2X1_LOC_743/A AND2X1_LOC_319/A 0.01fF
C16190 AND2X1_LOC_578/A OR2X1_LOC_237/Y 0.08fF
C16191 OR2X1_LOC_344/A OR2X1_LOC_675/Y 0.02fF
C16192 AND2X1_LOC_744/a_8_24# OR2X1_LOC_446/Y 0.05fF
C16193 AND2X1_LOC_661/A OR2X1_LOC_7/A 0.03fF
C16194 AND2X1_LOC_244/A AND2X1_LOC_657/A 0.07fF
C16195 AND2X1_LOC_654/a_8_24# OR2X1_LOC_7/A 0.02fF
C16196 AND2X1_LOC_538/a_8_24# OR2X1_LOC_427/A 0.06fF
C16197 AND2X1_LOC_70/Y D_INPUT_1 0.03fF
C16198 AND2X1_LOC_76/Y AND2X1_LOC_633/Y 0.06fF
C16199 AND2X1_LOC_78/a_36_24# OR2X1_LOC_36/Y 0.00fF
C16200 OR2X1_LOC_474/Y AND2X1_LOC_47/Y 0.18fF
C16201 AND2X1_LOC_727/B OR2X1_LOC_152/A 0.00fF
C16202 OR2X1_LOC_160/A OR2X1_LOC_647/a_8_216# 0.05fF
C16203 AND2X1_LOC_81/B OR2X1_LOC_473/Y 0.33fF
C16204 OR2X1_LOC_160/B OR2X1_LOC_493/Y 0.17fF
C16205 AND2X1_LOC_12/Y OR2X1_LOC_643/Y 0.03fF
C16206 OR2X1_LOC_682/a_36_216# OR2X1_LOC_743/A 0.00fF
C16207 OR2X1_LOC_160/B OR2X1_LOC_801/B 0.07fF
C16208 OR2X1_LOC_685/B AND2X1_LOC_51/Y 0.01fF
C16209 AND2X1_LOC_155/Y OR2X1_LOC_52/B 0.02fF
C16210 AND2X1_LOC_76/Y D_INPUT_0 0.03fF
C16211 OR2X1_LOC_447/Y OR2X1_LOC_724/a_8_216# 0.01fF
C16212 AND2X1_LOC_21/Y AND2X1_LOC_36/a_8_24# 0.01fF
C16213 D_INPUT_4 OR2X1_LOC_639/a_8_216# 0.14fF
C16214 OR2X1_LOC_209/A OR2X1_LOC_731/A 0.07fF
C16215 AND2X1_LOC_196/a_8_24# OR2X1_LOC_585/A 0.03fF
C16216 AND2X1_LOC_222/Y AND2X1_LOC_778/Y 0.02fF
C16217 OR2X1_LOC_264/a_8_216# OR2X1_LOC_121/B 0.01fF
C16218 OR2X1_LOC_131/A OR2X1_LOC_88/Y 0.00fF
C16219 OR2X1_LOC_230/a_8_216# OR2X1_LOC_52/B 0.04fF
C16220 D_INPUT_3 OR2X1_LOC_92/Y 0.03fF
C16221 OR2X1_LOC_437/A OR2X1_LOC_310/a_8_216# 0.03fF
C16222 OR2X1_LOC_22/Y OR2X1_LOC_265/Y 0.07fF
C16223 OR2X1_LOC_223/A OR2X1_LOC_776/a_36_216# 0.00fF
C16224 OR2X1_LOC_240/a_8_216# OR2X1_LOC_532/B 0.01fF
C16225 OR2X1_LOC_532/B OR2X1_LOC_739/A 0.03fF
C16226 OR2X1_LOC_412/a_36_216# OR2X1_LOC_39/A 0.00fF
C16227 OR2X1_LOC_662/A OR2X1_LOC_655/B 0.24fF
C16228 AND2X1_LOC_41/A OR2X1_LOC_205/Y 0.03fF
C16229 AND2X1_LOC_108/a_8_24# OR2X1_LOC_161/A 0.01fF
C16230 AND2X1_LOC_727/A OR2X1_LOC_44/Y 0.03fF
C16231 AND2X1_LOC_640/Y AND2X1_LOC_650/a_8_24# 0.04fF
C16232 OR2X1_LOC_748/A OR2X1_LOC_54/Y 0.01fF
C16233 OR2X1_LOC_114/Y OR2X1_LOC_62/B 0.02fF
C16234 OR2X1_LOC_602/Y AND2X1_LOC_31/Y 0.06fF
C16235 OR2X1_LOC_599/A AND2X1_LOC_477/A 0.07fF
C16236 AND2X1_LOC_95/Y OR2X1_LOC_276/B 0.01fF
C16237 OR2X1_LOC_659/B OR2X1_LOC_720/B 0.54fF
C16238 AND2X1_LOC_554/B OR2X1_LOC_64/Y 0.02fF
C16239 OR2X1_LOC_405/A AND2X1_LOC_109/a_8_24# 0.01fF
C16240 OR2X1_LOC_19/B OR2X1_LOC_609/A 0.01fF
C16241 AND2X1_LOC_633/Y OR2X1_LOC_52/B 0.02fF
C16242 OR2X1_LOC_184/Y OR2X1_LOC_427/A 0.18fF
C16243 AND2X1_LOC_708/a_8_24# OR2X1_LOC_743/A 0.01fF
C16244 AND2X1_LOC_821/a_36_24# OR2X1_LOC_130/A 0.01fF
C16245 OR2X1_LOC_549/A OR2X1_LOC_367/a_36_216# 0.01fF
C16246 OR2X1_LOC_836/a_8_216# OR2X1_LOC_835/Y 0.05fF
C16247 OR2X1_LOC_92/Y AND2X1_LOC_483/Y 0.01fF
C16248 OR2X1_LOC_814/A OR2X1_LOC_155/A 0.03fF
C16249 AND2X1_LOC_851/B OR2X1_LOC_237/a_36_216# 0.01fF
C16250 OR2X1_LOC_71/Y AND2X1_LOC_361/A 0.28fF
C16251 OR2X1_LOC_720/B OR2X1_LOC_720/a_36_216# 0.03fF
C16252 OR2X1_LOC_474/Y OR2X1_LOC_598/A 0.07fF
C16253 AND2X1_LOC_784/Y OR2X1_LOC_437/A 0.02fF
C16254 OR2X1_LOC_532/B OR2X1_LOC_269/B 0.26fF
C16255 D_INPUT_0 OR2X1_LOC_52/B 3.70fF
C16256 OR2X1_LOC_84/B D_INPUT_0 0.00fF
C16257 AND2X1_LOC_306/a_8_24# AND2X1_LOC_31/Y 0.01fF
C16258 AND2X1_LOC_12/Y OR2X1_LOC_786/Y 0.15fF
C16259 OR2X1_LOC_95/Y OR2X1_LOC_44/Y 2.17fF
C16260 OR2X1_LOC_1/a_8_216# OR2X1_LOC_51/B 0.03fF
C16261 INPUT_0 OR2X1_LOC_198/A 0.02fF
C16262 OR2X1_LOC_696/Y OR2X1_LOC_64/Y 0.09fF
C16263 AND2X1_LOC_326/A OR2X1_LOC_64/Y 0.01fF
C16264 AND2X1_LOC_41/A OR2X1_LOC_750/Y 0.04fF
C16265 OR2X1_LOC_368/A OR2X1_LOC_44/Y 0.03fF
C16266 OR2X1_LOC_70/Y AND2X1_LOC_687/B 0.22fF
C16267 OR2X1_LOC_814/A OR2X1_LOC_392/a_8_216# 0.01fF
C16268 INPUT_1 OR2X1_LOC_74/A 0.09fF
C16269 OR2X1_LOC_628/Y AND2X1_LOC_483/a_8_24# 0.01fF
C16270 OR2X1_LOC_851/A OR2X1_LOC_318/B 0.12fF
C16271 OR2X1_LOC_312/Y AND2X1_LOC_169/a_8_24# 0.14fF
C16272 AND2X1_LOC_59/Y AND2X1_LOC_271/a_8_24# 0.17fF
C16273 OR2X1_LOC_683/Y OR2X1_LOC_684/Y 0.01fF
C16274 OR2X1_LOC_31/Y AND2X1_LOC_654/a_36_24# 0.01fF
C16275 OR2X1_LOC_6/B OR2X1_LOC_771/B 3.69fF
C16276 AND2X1_LOC_739/a_8_24# GATE_811 0.01fF
C16277 AND2X1_LOC_12/Y OR2X1_LOC_644/A 0.02fF
C16278 AND2X1_LOC_92/Y OR2X1_LOC_317/B 0.11fF
C16279 AND2X1_LOC_593/Y OR2X1_LOC_419/Y 0.01fF
C16280 OR2X1_LOC_475/B OR2X1_LOC_228/Y 0.08fF
C16281 VDD OR2X1_LOC_571/Y -0.00fF
C16282 OR2X1_LOC_140/B OR2X1_LOC_161/B 0.03fF
C16283 VDD OR2X1_LOC_374/a_8_216# 0.00fF
C16284 OR2X1_LOC_116/A OR2X1_LOC_598/A 0.01fF
C16285 OR2X1_LOC_287/B AND2X1_LOC_250/a_8_24# 0.01fF
C16286 OR2X1_LOC_85/a_8_216# OR2X1_LOC_85/A 0.01fF
C16287 AND2X1_LOC_280/a_8_24# OR2X1_LOC_375/A 0.07fF
C16288 AND2X1_LOC_23/a_8_24# OR2X1_LOC_19/B 0.04fF
C16289 OR2X1_LOC_45/B AND2X1_LOC_473/Y 0.02fF
C16290 VDD OR2X1_LOC_469/B 0.14fF
C16291 OR2X1_LOC_167/Y OR2X1_LOC_64/Y 0.02fF
C16292 OR2X1_LOC_65/B AND2X1_LOC_656/a_8_24# 0.01fF
C16293 OR2X1_LOC_217/Y OR2X1_LOC_598/A 0.02fF
C16294 AND2X1_LOC_624/A AND2X1_LOC_222/Y 0.03fF
C16295 OR2X1_LOC_45/B OR2X1_LOC_816/A 0.03fF
C16296 AND2X1_LOC_351/Y OR2X1_LOC_417/A 0.02fF
C16297 OR2X1_LOC_85/A AND2X1_LOC_202/a_36_24# 0.00fF
C16298 AND2X1_LOC_70/Y OR2X1_LOC_180/B 0.03fF
C16299 OR2X1_LOC_323/A AND2X1_LOC_719/Y 0.03fF
C16300 AND2X1_LOC_100/a_36_24# OR2X1_LOC_86/A 0.00fF
C16301 AND2X1_LOC_227/Y OR2X1_LOC_245/a_8_216# 0.01fF
C16302 AND2X1_LOC_810/A AND2X1_LOC_802/Y 0.01fF
C16303 OR2X1_LOC_479/a_8_216# OR2X1_LOC_223/A 0.01fF
C16304 OR2X1_LOC_847/a_8_216# OR2X1_LOC_80/A 0.02fF
C16305 AND2X1_LOC_91/B AND2X1_LOC_371/a_8_24# 0.15fF
C16306 OR2X1_LOC_334/B AND2X1_LOC_36/Y 0.01fF
C16307 AND2X1_LOC_91/B AND2X1_LOC_18/Y 0.32fF
C16308 OR2X1_LOC_404/Y D_INPUT_1 0.07fF
C16309 OR2X1_LOC_185/A OR2X1_LOC_366/Y 0.03fF
C16310 OR2X1_LOC_736/Y OR2X1_LOC_344/A 0.03fF
C16311 OR2X1_LOC_604/A OR2X1_LOC_744/Y 0.21fF
C16312 AND2X1_LOC_328/a_8_24# AND2X1_LOC_36/Y 0.01fF
C16313 VDD AND2X1_LOC_244/A 0.28fF
C16314 AND2X1_LOC_715/A OR2X1_LOC_310/a_8_216# 0.16fF
C16315 OR2X1_LOC_45/B AND2X1_LOC_707/a_8_24# 0.03fF
C16316 OR2X1_LOC_334/B OR2X1_LOC_334/A 0.48fF
C16317 OR2X1_LOC_186/Y OR2X1_LOC_325/B 1.76fF
C16318 OR2X1_LOC_490/a_36_216# AND2X1_LOC_243/Y 0.01fF
C16319 OR2X1_LOC_47/Y AND2X1_LOC_839/A 0.01fF
C16320 VDD OR2X1_LOC_16/A 1.24fF
C16321 OR2X1_LOC_159/a_8_216# OR2X1_LOC_671/Y 0.02fF
C16322 OR2X1_LOC_158/A AND2X1_LOC_194/Y 0.03fF
C16323 AND2X1_LOC_568/B AND2X1_LOC_810/B 0.03fF
C16324 OR2X1_LOC_22/Y AND2X1_LOC_205/a_8_24# 0.04fF
C16325 AND2X1_LOC_92/Y AND2X1_LOC_44/Y 1.81fF
C16326 OR2X1_LOC_566/A OR2X1_LOC_808/B 0.05fF
C16327 AND2X1_LOC_533/a_8_24# OR2X1_LOC_703/Y 0.10fF
C16328 AND2X1_LOC_22/Y OR2X1_LOC_235/B 0.16fF
C16329 OR2X1_LOC_31/Y OR2X1_LOC_51/B 0.01fF
C16330 OR2X1_LOC_715/B OR2X1_LOC_140/A 0.17fF
C16331 OR2X1_LOC_123/a_8_216# OR2X1_LOC_549/A 0.01fF
C16332 OR2X1_LOC_91/A AND2X1_LOC_786/Y 0.07fF
C16333 OR2X1_LOC_62/B OR2X1_LOC_140/a_36_216# 0.00fF
C16334 OR2X1_LOC_528/Y AND2X1_LOC_508/B 0.02fF
C16335 OR2X1_LOC_475/a_8_216# OR2X1_LOC_392/B 0.12fF
C16336 AND2X1_LOC_702/Y OR2X1_LOC_320/a_8_216# 0.01fF
C16337 OR2X1_LOC_287/B OR2X1_LOC_349/B 0.02fF
C16338 D_INPUT_0 OR2X1_LOC_728/B 0.52fF
C16339 VDD OR2X1_LOC_108/Y 0.06fF
C16340 OR2X1_LOC_535/A OR2X1_LOC_538/A 0.02fF
C16341 AND2X1_LOC_362/B OR2X1_LOC_122/A 0.05fF
C16342 OR2X1_LOC_632/A OR2X1_LOC_115/B 0.01fF
C16343 OR2X1_LOC_527/a_8_216# OR2X1_LOC_56/A 0.01fF
C16344 AND2X1_LOC_557/Y AND2X1_LOC_561/a_8_24# -0.00fF
C16345 OR2X1_LOC_3/Y OR2X1_LOC_376/Y 0.02fF
C16346 OR2X1_LOC_678/Y OR2X1_LOC_596/A 0.02fF
C16347 OR2X1_LOC_602/B AND2X1_LOC_31/Y 0.05fF
C16348 OR2X1_LOC_511/Y OR2X1_LOC_525/a_36_216# 0.02fF
C16349 OR2X1_LOC_482/a_8_216# AND2X1_LOC_456/B 0.02fF
C16350 OR2X1_LOC_45/B AND2X1_LOC_649/a_8_24# 0.01fF
C16351 AND2X1_LOC_521/a_8_24# OR2X1_LOC_474/Y 0.13fF
C16352 OR2X1_LOC_549/Y OR2X1_LOC_577/a_8_216# 0.00fF
C16353 VDD AND2X1_LOC_121/a_8_24# 0.00fF
C16354 OR2X1_LOC_45/B OR2X1_LOC_45/Y 0.47fF
C16355 OR2X1_LOC_486/B OR2X1_LOC_550/B 0.34fF
C16356 AND2X1_LOC_675/Y OR2X1_LOC_505/Y 0.02fF
C16357 AND2X1_LOC_722/a_8_24# AND2X1_LOC_722/Y 0.01fF
C16358 AND2X1_LOC_719/Y AND2X1_LOC_723/Y 0.15fF
C16359 OR2X1_LOC_154/A OR2X1_LOC_214/A 0.03fF
C16360 OR2X1_LOC_604/A AND2X1_LOC_474/A 0.05fF
C16361 OR2X1_LOC_40/Y AND2X1_LOC_861/B 0.07fF
C16362 OR2X1_LOC_538/A AND2X1_LOC_323/a_8_24# 0.00fF
C16363 AND2X1_LOC_555/Y OR2X1_LOC_36/Y 0.00fF
C16364 OR2X1_LOC_785/a_8_216# AND2X1_LOC_92/Y 0.06fF
C16365 OR2X1_LOC_78/A OR2X1_LOC_244/Y 0.02fF
C16366 OR2X1_LOC_48/B OR2X1_LOC_12/Y 3.68fF
C16367 OR2X1_LOC_303/a_36_216# OR2X1_LOC_468/Y 0.00fF
C16368 OR2X1_LOC_747/a_8_216# AND2X1_LOC_781/Y 0.48fF
C16369 VDD OR2X1_LOC_624/a_8_216# 0.00fF
C16370 OR2X1_LOC_185/A OR2X1_LOC_548/B 0.05fF
C16371 AND2X1_LOC_675/Y AND2X1_LOC_658/A 0.03fF
C16372 AND2X1_LOC_367/A AND2X1_LOC_325/a_8_24# 0.16fF
C16373 OR2X1_LOC_45/B AND2X1_LOC_807/Y 3.10fF
C16374 OR2X1_LOC_154/A AND2X1_LOC_7/B 8.44fF
C16375 AND2X1_LOC_274/a_8_24# OR2X1_LOC_16/A 0.17fF
C16376 OR2X1_LOC_18/Y OR2X1_LOC_12/Y 2.67fF
C16377 AND2X1_LOC_717/Y AND2X1_LOC_476/Y 0.07fF
C16378 OR2X1_LOC_744/A OR2X1_LOC_484/a_36_216# 0.00fF
C16379 AND2X1_LOC_564/B OR2X1_LOC_372/Y 0.04fF
C16380 D_GATE_741 OR2X1_LOC_192/A 0.01fF
C16381 OR2X1_LOC_91/A AND2X1_LOC_218/Y 0.06fF
C16382 OR2X1_LOC_501/B OR2X1_LOC_78/A 0.12fF
C16383 OR2X1_LOC_696/A OR2X1_LOC_3/Y 0.56fF
C16384 VDD OR2X1_LOC_274/Y 0.09fF
C16385 AND2X1_LOC_1/Y INPUT_6 0.29fF
C16386 AND2X1_LOC_212/Y OR2X1_LOC_39/A 0.10fF
C16387 OR2X1_LOC_190/B OR2X1_LOC_190/Y 0.10fF
C16388 OR2X1_LOC_160/B OR2X1_LOC_61/B 0.03fF
C16389 AND2X1_LOC_704/a_8_24# AND2X1_LOC_452/Y 0.02fF
C16390 AND2X1_LOC_358/Y OR2X1_LOC_6/A 0.00fF
C16391 OR2X1_LOC_865/A OR2X1_LOC_269/B 0.70fF
C16392 AND2X1_LOC_721/Y OR2X1_LOC_26/Y 0.09fF
C16393 OR2X1_LOC_49/A OR2X1_LOC_236/a_8_216# 0.13fF
C16394 OR2X1_LOC_519/Y AND2X1_LOC_566/B 0.00fF
C16395 AND2X1_LOC_741/Y AND2X1_LOC_192/Y 0.14fF
C16396 OR2X1_LOC_833/B AND2X1_LOC_626/a_8_24# 0.02fF
C16397 OR2X1_LOC_862/B OR2X1_LOC_862/A 0.56fF
C16398 OR2X1_LOC_599/A AND2X1_LOC_703/Y 0.02fF
C16399 OR2X1_LOC_25/a_8_216# INPUT_7 0.08fF
C16400 AND2X1_LOC_2/Y AND2X1_LOC_2/a_8_24# 0.01fF
C16401 OR2X1_LOC_318/A OR2X1_LOC_87/A 0.05fF
C16402 OR2X1_LOC_235/B OR2X1_LOC_244/B 0.03fF
C16403 OR2X1_LOC_756/B OR2X1_LOC_570/A 0.02fF
C16404 AND2X1_LOC_798/a_8_24# AND2X1_LOC_798/Y 0.01fF
C16405 OR2X1_LOC_185/A OR2X1_LOC_786/A 0.02fF
C16406 AND2X1_LOC_169/a_8_24# OR2X1_LOC_13/B 0.01fF
C16407 AND2X1_LOC_544/Y OR2X1_LOC_680/Y 0.09fF
C16408 OR2X1_LOC_303/A OR2X1_LOC_703/A 0.03fF
C16409 OR2X1_LOC_368/a_8_216# OR2X1_LOC_109/Y 0.03fF
C16410 OR2X1_LOC_6/B OR2X1_LOC_402/Y 0.04fF
C16411 OR2X1_LOC_276/B OR2X1_LOC_269/A 0.02fF
C16412 OR2X1_LOC_703/B OR2X1_LOC_151/A 0.08fF
C16413 AND2X1_LOC_383/a_8_24# OR2X1_LOC_3/Y 0.01fF
C16414 AND2X1_LOC_721/Y OR2X1_LOC_89/A 0.05fF
C16415 AND2X1_LOC_658/B OR2X1_LOC_427/A 0.08fF
C16416 AND2X1_LOC_364/Y AND2X1_LOC_857/Y 0.12fF
C16417 OR2X1_LOC_832/a_8_216# OR2X1_LOC_506/A 0.00fF
C16418 OR2X1_LOC_83/A OR2X1_LOC_414/Y 0.73fF
C16419 AND2X1_LOC_70/Y OR2X1_LOC_737/A 0.14fF
C16420 OR2X1_LOC_604/A AND2X1_LOC_593/Y 0.03fF
C16421 AND2X1_LOC_72/Y AND2X1_LOC_18/Y 0.00fF
C16422 AND2X1_LOC_367/A OR2X1_LOC_517/A 0.05fF
C16423 AND2X1_LOC_851/B OR2X1_LOC_437/A 0.10fF
C16424 OR2X1_LOC_761/Y AND2X1_LOC_434/Y 0.03fF
C16425 AND2X1_LOC_486/Y OR2X1_LOC_484/Y 0.78fF
C16426 VDD AND2X1_LOC_748/a_8_24# -0.00fF
C16427 OR2X1_LOC_440/a_8_216# OR2X1_LOC_161/A 0.03fF
C16428 OR2X1_LOC_329/B AND2X1_LOC_276/a_36_24# 0.01fF
C16429 OR2X1_LOC_151/A OR2X1_LOC_87/A 11.18fF
C16430 AND2X1_LOC_47/Y OR2X1_LOC_771/B 0.03fF
C16431 AND2X1_LOC_208/a_8_24# AND2X1_LOC_208/B 0.00fF
C16432 OR2X1_LOC_68/Y OR2X1_LOC_776/A 0.00fF
C16433 OR2X1_LOC_64/Y OR2X1_LOC_503/a_8_216# 0.06fF
C16434 AND2X1_LOC_70/Y AND2X1_LOC_95/Y 1.30fF
C16435 AND2X1_LOC_59/Y OR2X1_LOC_641/a_8_216# 0.01fF
C16436 OR2X1_LOC_589/A OR2X1_LOC_69/Y 0.30fF
C16437 OR2X1_LOC_377/A OR2X1_LOC_66/A 0.22fF
C16438 OR2X1_LOC_250/Y OR2X1_LOC_51/Y 0.19fF
C16439 VDD OR2X1_LOC_640/a_8_216# 0.21fF
C16440 OR2X1_LOC_778/A AND2X1_LOC_7/B 0.02fF
C16441 OR2X1_LOC_479/Y OR2X1_LOC_357/B 0.03fF
C16442 AND2X1_LOC_362/B AND2X1_LOC_560/B 0.01fF
C16443 OR2X1_LOC_834/A AND2X1_LOC_305/a_8_24# 0.08fF
C16444 AND2X1_LOC_211/B AND2X1_LOC_212/Y 0.00fF
C16445 OR2X1_LOC_52/B AND2X1_LOC_771/B 0.06fF
C16446 OR2X1_LOC_494/a_8_216# OR2X1_LOC_92/Y -0.00fF
C16447 OR2X1_LOC_91/Y OR2X1_LOC_600/A 0.12fF
C16448 D_GATE_811 OR2X1_LOC_269/B 0.09fF
C16449 AND2X1_LOC_730/a_8_24# AND2X1_LOC_803/B 0.01fF
C16450 OR2X1_LOC_604/A OR2X1_LOC_85/A 0.11fF
C16451 OR2X1_LOC_270/a_8_216# AND2X1_LOC_18/Y 0.08fF
C16452 OR2X1_LOC_441/Y AND2X1_LOC_147/a_8_24# 0.07fF
C16453 OR2X1_LOC_467/A OR2X1_LOC_467/a_8_216# 0.04fF
C16454 OR2X1_LOC_287/B D_GATE_662 0.02fF
C16455 AND2X1_LOC_42/B OR2X1_LOC_548/a_8_216# 0.05fF
C16456 AND2X1_LOC_51/Y OR2X1_LOC_474/B 0.26fF
C16457 AND2X1_LOC_474/A AND2X1_LOC_850/a_8_24# 0.01fF
C16458 OR2X1_LOC_51/Y AND2X1_LOC_466/a_8_24# 0.01fF
C16459 AND2X1_LOC_714/B OR2X1_LOC_7/A 0.23fF
C16460 OR2X1_LOC_482/Y AND2X1_LOC_493/a_8_24# 0.12fF
C16461 OR2X1_LOC_45/B OR2X1_LOC_488/Y 0.00fF
C16462 OR2X1_LOC_6/B OR2X1_LOC_217/a_8_216# 0.07fF
C16463 AND2X1_LOC_3/Y OR2X1_LOC_361/a_8_216# 0.01fF
C16464 OR2X1_LOC_47/Y OR2X1_LOC_749/Y 0.04fF
C16465 OR2X1_LOC_243/A OR2X1_LOC_78/B 0.08fF
C16466 OR2X1_LOC_108/Y OR2X1_LOC_491/Y 0.02fF
C16467 OR2X1_LOC_203/Y OR2X1_LOC_66/A 0.02fF
C16468 OR2X1_LOC_52/B AND2X1_LOC_784/a_8_24# 0.02fF
C16469 OR2X1_LOC_857/B OR2X1_LOC_688/Y 0.02fF
C16470 OR2X1_LOC_41/a_8_216# OR2X1_LOC_13/B 0.08fF
C16471 OR2X1_LOC_6/B AND2X1_LOC_838/a_36_24# -0.01fF
C16472 OR2X1_LOC_482/Y OR2X1_LOC_89/A 0.17fF
C16473 OR2X1_LOC_319/B OR2X1_LOC_620/Y 0.00fF
C16474 AND2X1_LOC_95/Y OR2X1_LOC_703/A 1.86fF
C16475 OR2X1_LOC_604/A AND2X1_LOC_602/a_8_24# 0.01fF
C16476 AND2X1_LOC_76/Y AND2X1_LOC_276/a_8_24# 0.01fF
C16477 OR2X1_LOC_837/Y OR2X1_LOC_18/Y 0.09fF
C16478 OR2X1_LOC_51/Y OR2X1_LOC_36/Y 0.68fF
C16479 OR2X1_LOC_160/A AND2X1_LOC_41/A 0.93fF
C16480 AND2X1_LOC_64/Y AND2X1_LOC_53/Y 0.17fF
C16481 OR2X1_LOC_158/A OR2X1_LOC_17/Y 0.10fF
C16482 OR2X1_LOC_333/B OR2X1_LOC_648/B 0.03fF
C16483 OR2X1_LOC_426/B AND2X1_LOC_361/A 0.10fF
C16484 OR2X1_LOC_45/B AND2X1_LOC_727/A 0.00fF
C16485 OR2X1_LOC_158/A OR2X1_LOC_282/Y 0.01fF
C16486 D_INPUT_0 OR2X1_LOC_338/A 0.07fF
C16487 OR2X1_LOC_74/A AND2X1_LOC_778/Y 0.00fF
C16488 OR2X1_LOC_56/A AND2X1_LOC_818/a_8_24# 0.03fF
C16489 OR2X1_LOC_318/Y OR2X1_LOC_620/Y 0.07fF
C16490 AND2X1_LOC_56/B AND2X1_LOC_628/a_8_24# 0.01fF
C16491 AND2X1_LOC_777/a_8_24# OR2X1_LOC_91/A 0.12fF
C16492 OR2X1_LOC_329/B OR2X1_LOC_495/a_8_216# 0.02fF
C16493 AND2X1_LOC_456/B AND2X1_LOC_859/a_8_24# 0.01fF
C16494 OR2X1_LOC_856/B OR2X1_LOC_623/a_8_216# 0.02fF
C16495 AND2X1_LOC_736/a_36_24# OR2X1_LOC_189/A 0.00fF
C16496 AND2X1_LOC_325/a_8_24# OR2X1_LOC_74/A 0.03fF
C16497 OR2X1_LOC_771/B OR2X1_LOC_598/A 0.40fF
C16498 OR2X1_LOC_668/Y OR2X1_LOC_721/Y 0.04fF
C16499 OR2X1_LOC_64/Y AND2X1_LOC_476/Y 0.14fF
C16500 AND2X1_LOC_362/B OR2X1_LOC_64/Y 0.02fF
C16501 OR2X1_LOC_80/A OR2X1_LOC_71/A 0.05fF
C16502 OR2X1_LOC_155/A OR2X1_LOC_715/A 0.07fF
C16503 OR2X1_LOC_56/A AND2X1_LOC_458/a_36_24# 0.01fF
C16504 OR2X1_LOC_756/B OR2X1_LOC_593/a_36_216# 0.00fF
C16505 AND2X1_LOC_59/Y OR2X1_LOC_785/B 0.02fF
C16506 AND2X1_LOC_12/Y OR2X1_LOC_851/A 0.00fF
C16507 AND2X1_LOC_520/a_8_24# AND2X1_LOC_831/Y 0.02fF
C16508 VDD OR2X1_LOC_273/a_8_216# 0.00fF
C16509 AND2X1_LOC_550/a_36_24# AND2X1_LOC_711/Y 0.01fF
C16510 AND2X1_LOC_64/Y OR2X1_LOC_223/A 0.03fF
C16511 AND2X1_LOC_377/Y OR2X1_LOC_585/A 0.06fF
C16512 OR2X1_LOC_816/Y OR2X1_LOC_89/A 0.04fF
C16513 OR2X1_LOC_391/A OR2X1_LOC_269/B 0.44fF
C16514 OR2X1_LOC_589/A AND2X1_LOC_537/Y 0.01fF
C16515 OR2X1_LOC_297/a_8_216# OR2X1_LOC_44/Y 0.03fF
C16516 AND2X1_LOC_550/a_36_24# OR2X1_LOC_70/Y 0.00fF
C16517 OR2X1_LOC_287/B OR2X1_LOC_78/a_8_216# 0.01fF
C16518 OR2X1_LOC_186/Y D_INPUT_0 0.01fF
C16519 OR2X1_LOC_121/B OR2X1_LOC_641/A 0.04fF
C16520 OR2X1_LOC_185/A OR2X1_LOC_624/A 0.03fF
C16521 OR2X1_LOC_464/B OR2X1_LOC_464/A 0.15fF
C16522 OR2X1_LOC_122/a_8_216# OR2X1_LOC_3/Y 0.01fF
C16523 AND2X1_LOC_214/A OR2X1_LOC_7/A 0.05fF
C16524 AND2X1_LOC_716/Y AND2X1_LOC_354/B 0.08fF
C16525 OR2X1_LOC_45/B OR2X1_LOC_95/Y 0.56fF
C16526 OR2X1_LOC_791/B AND2X1_LOC_95/Y 0.03fF
C16527 D_INPUT_5 AND2X1_LOC_64/a_8_24# 0.09fF
C16528 OR2X1_LOC_36/Y OR2X1_LOC_16/Y 0.02fF
C16529 AND2X1_LOC_486/Y AND2X1_LOC_576/Y 0.10fF
C16530 OR2X1_LOC_417/Y OR2X1_LOC_600/A 0.04fF
C16531 OR2X1_LOC_45/B OR2X1_LOC_368/A 0.01fF
C16532 AND2X1_LOC_508/A OR2X1_LOC_239/a_8_216# 0.01fF
C16533 AND2X1_LOC_861/B OR2X1_LOC_7/A 0.02fF
C16534 OR2X1_LOC_858/B OR2X1_LOC_287/B 0.01fF
C16535 OR2X1_LOC_121/B AND2X1_LOC_299/a_36_24# 0.01fF
C16536 AND2X1_LOC_276/a_8_24# OR2X1_LOC_52/B 0.13fF
C16537 OR2X1_LOC_160/A OR2X1_LOC_662/A 0.00fF
C16538 AND2X1_LOC_578/A AND2X1_LOC_858/B 0.08fF
C16539 OR2X1_LOC_494/A OR2X1_LOC_47/Y 0.03fF
C16540 OR2X1_LOC_851/A OR2X1_LOC_841/B 0.86fF
C16541 AND2X1_LOC_832/a_8_24# OR2X1_LOC_44/Y 0.02fF
C16542 AND2X1_LOC_654/Y AND2X1_LOC_354/B 0.07fF
C16543 AND2X1_LOC_605/Y OR2X1_LOC_743/A 0.06fF
C16544 AND2X1_LOC_40/Y OR2X1_LOC_84/B 0.47fF
C16545 INPUT_5 OR2X1_LOC_21/a_8_216# 0.18fF
C16546 OR2X1_LOC_604/A AND2X1_LOC_470/a_8_24# 0.01fF
C16547 OR2X1_LOC_18/Y OR2X1_LOC_95/a_36_216# 0.02fF
C16548 OR2X1_LOC_26/Y OR2X1_LOC_586/Y 0.04fF
C16549 OR2X1_LOC_97/a_36_216# OR2X1_LOC_78/A 0.01fF
C16550 OR2X1_LOC_663/A OR2X1_LOC_557/A 0.00fF
C16551 OR2X1_LOC_61/B OR2X1_LOC_219/B 0.03fF
C16552 OR2X1_LOC_36/Y AND2X1_LOC_642/a_8_24# 0.01fF
C16553 OR2X1_LOC_490/Y OR2X1_LOC_517/A 1.24fF
C16554 OR2X1_LOC_39/A OR2X1_LOC_265/Y 0.07fF
C16555 OR2X1_LOC_517/A OR2X1_LOC_74/A 0.06fF
C16556 OR2X1_LOC_643/A OR2X1_LOC_560/a_8_216# 0.01fF
C16557 AND2X1_LOC_362/B OR2X1_LOC_417/A 0.03fF
C16558 OR2X1_LOC_417/A AND2X1_LOC_476/Y 0.21fF
C16559 OR2X1_LOC_502/A OR2X1_LOC_646/a_8_216# 0.01fF
C16560 OR2X1_LOC_18/Y AND2X1_LOC_650/Y 0.17fF
C16561 OR2X1_LOC_154/A OR2X1_LOC_805/A 0.17fF
C16562 OR2X1_LOC_305/Y OR2X1_LOC_619/Y 0.01fF
C16563 AND2X1_LOC_64/Y OR2X1_LOC_705/B 0.01fF
C16564 OR2X1_LOC_405/Y OR2X1_LOC_358/B 0.02fF
C16565 VDD AND2X1_LOC_687/Y 0.04fF
C16566 AND2X1_LOC_51/Y OR2X1_LOC_561/Y 0.01fF
C16567 OR2X1_LOC_416/Y OR2X1_LOC_59/Y 0.04fF
C16568 AND2X1_LOC_51/Y OR2X1_LOC_78/Y 0.02fF
C16569 OR2X1_LOC_92/Y AND2X1_LOC_276/Y 0.05fF
C16570 AND2X1_LOC_155/a_8_24# AND2X1_LOC_154/Y 0.23fF
C16571 OR2X1_LOC_269/a_36_216# OR2X1_LOC_269/B 0.03fF
C16572 INPUT_4 OR2X1_LOC_25/a_8_216# 0.01fF
C16573 OR2X1_LOC_185/A OR2X1_LOC_552/a_8_216# 0.01fF
C16574 OR2X1_LOC_604/A OR2X1_LOC_226/Y 0.01fF
C16575 OR2X1_LOC_702/A OR2X1_LOC_175/B 0.00fF
C16576 AND2X1_LOC_175/a_8_24# OR2X1_LOC_18/Y 0.01fF
C16577 OR2X1_LOC_680/A OR2X1_LOC_36/Y 0.33fF
C16578 OR2X1_LOC_80/Y OR2X1_LOC_85/A 0.02fF
C16579 OR2X1_LOC_695/a_8_216# OR2X1_LOC_3/Y 0.02fF
C16580 OR2X1_LOC_99/A AND2X1_LOC_7/B 0.05fF
C16581 AND2X1_LOC_172/a_8_24# OR2X1_LOC_532/B 0.01fF
C16582 OR2X1_LOC_844/Y OR2X1_LOC_659/A 0.03fF
C16583 AND2X1_LOC_763/a_36_24# AND2X1_LOC_48/A 0.01fF
C16584 OR2X1_LOC_246/Y OR2X1_LOC_248/Y 0.09fF
C16585 AND2X1_LOC_95/Y OR2X1_LOC_653/a_8_216# 0.06fF
C16586 AND2X1_LOC_848/A OR2X1_LOC_428/A 0.02fF
C16587 AND2X1_LOC_654/B OR2X1_LOC_43/a_8_216# 0.17fF
C16588 OR2X1_LOC_26/Y AND2X1_LOC_859/a_36_24# 0.00fF
C16589 OR2X1_LOC_833/Y OR2X1_LOC_241/B 0.01fF
C16590 OR2X1_LOC_743/A OR2X1_LOC_829/a_36_216# 0.00fF
C16591 OR2X1_LOC_600/A D_INPUT_3 11.43fF
C16592 AND2X1_LOC_211/B OR2X1_LOC_265/Y 0.19fF
C16593 OR2X1_LOC_9/Y D_INPUT_1 0.71fF
C16594 OR2X1_LOC_272/Y OR2X1_LOC_18/Y 0.08fF
C16595 OR2X1_LOC_175/Y OR2X1_LOC_228/Y 0.22fF
C16596 OR2X1_LOC_362/A D_INPUT_1 0.03fF
C16597 OR2X1_LOC_74/A AND2X1_LOC_624/A 0.07fF
C16598 AND2X1_LOC_580/A AND2X1_LOC_474/Y 0.06fF
C16599 OR2X1_LOC_158/A AND2X1_LOC_792/Y 0.09fF
C16600 OR2X1_LOC_675/Y OR2X1_LOC_161/B 0.02fF
C16601 OR2X1_LOC_736/a_8_216# AND2X1_LOC_44/Y 0.01fF
C16602 AND2X1_LOC_342/a_8_24# OR2X1_LOC_585/A 0.01fF
C16603 AND2X1_LOC_259/Y OR2X1_LOC_236/a_8_216# 0.00fF
C16604 OR2X1_LOC_449/A OR2X1_LOC_449/B 0.00fF
C16605 AND2X1_LOC_22/Y OR2X1_LOC_779/B 0.01fF
C16606 OR2X1_LOC_329/B OR2X1_LOC_238/a_8_216# 0.02fF
C16607 OR2X1_LOC_563/A OR2X1_LOC_68/B 0.05fF
C16608 OR2X1_LOC_258/Y AND2X1_LOC_848/Y 0.03fF
C16609 AND2X1_LOC_95/Y OR2X1_LOC_404/Y 0.02fF
C16610 OR2X1_LOC_158/A AND2X1_LOC_259/a_8_24# 0.02fF
C16611 AND2X1_LOC_525/a_36_24# OR2X1_LOC_375/A 0.01fF
C16612 OR2X1_LOC_468/a_8_216# OR2X1_LOC_78/B 0.01fF
C16613 OR2X1_LOC_805/A OR2X1_LOC_778/A 0.01fF
C16614 OR2X1_LOC_691/Y OR2X1_LOC_228/Y 0.03fF
C16615 AND2X1_LOC_851/a_8_24# AND2X1_LOC_851/B 0.01fF
C16616 OR2X1_LOC_748/A OR2X1_LOC_89/A 0.01fF
C16617 OR2X1_LOC_417/Y OR2X1_LOC_619/Y 13.69fF
C16618 OR2X1_LOC_744/A AND2X1_LOC_796/Y 0.11fF
C16619 OR2X1_LOC_291/Y OR2X1_LOC_619/Y 0.07fF
C16620 AND2X1_LOC_680/a_8_24# OR2X1_LOC_506/A 0.01fF
C16621 AND2X1_LOC_227/Y AND2X1_LOC_842/a_8_24# 0.09fF
C16622 AND2X1_LOC_35/Y AND2X1_LOC_853/a_8_24# 0.06fF
C16623 OR2X1_LOC_815/a_8_216# OR2X1_LOC_815/Y -0.00fF
C16624 OR2X1_LOC_185/A OR2X1_LOC_54/Y 0.07fF
C16625 OR2X1_LOC_271/Y AND2X1_LOC_276/Y 0.02fF
C16626 AND2X1_LOC_572/A AND2X1_LOC_663/B 0.06fF
C16627 OR2X1_LOC_748/A OR2X1_LOC_820/Y 0.01fF
C16628 AND2X1_LOC_356/a_8_24# OR2X1_LOC_311/Y 0.01fF
C16629 AND2X1_LOC_395/a_8_24# OR2X1_LOC_401/A 0.21fF
C16630 OR2X1_LOC_578/a_36_216# OR2X1_LOC_578/B 0.00fF
C16631 AND2X1_LOC_227/Y AND2X1_LOC_141/A 0.01fF
C16632 AND2X1_LOC_387/B OR2X1_LOC_155/A 0.07fF
C16633 AND2X1_LOC_831/Y OR2X1_LOC_92/Y 0.07fF
C16634 OR2X1_LOC_154/A OR2X1_LOC_436/a_8_216# 0.05fF
C16635 AND2X1_LOC_59/Y OR2X1_LOC_643/Y 0.01fF
C16636 OR2X1_LOC_513/Y OR2X1_LOC_713/A 0.01fF
C16637 AND2X1_LOC_390/B OR2X1_LOC_312/Y 0.02fF
C16638 OR2X1_LOC_520/Y AND2X1_LOC_518/a_8_24# 0.10fF
C16639 OR2X1_LOC_304/Y OR2X1_LOC_26/Y 0.02fF
C16640 AND2X1_LOC_40/Y OR2X1_LOC_651/A 3.28fF
C16641 OR2X1_LOC_862/B AND2X1_LOC_225/a_36_24# 0.00fF
C16642 INPUT_3 AND2X1_LOC_5/a_8_24# 0.11fF
C16643 AND2X1_LOC_863/Y AND2X1_LOC_654/Y 0.04fF
C16644 OR2X1_LOC_51/Y OR2X1_LOC_419/Y 0.06fF
C16645 OR2X1_LOC_577/Y OR2X1_LOC_366/Y 0.47fF
C16646 OR2X1_LOC_662/A OR2X1_LOC_655/A 0.00fF
C16647 AND2X1_LOC_11/Y AND2X1_LOC_47/Y 0.08fF
C16648 OR2X1_LOC_520/Y AND2X1_LOC_48/A 0.54fF
C16649 OR2X1_LOC_43/A OR2X1_LOC_43/a_8_216# 0.01fF
C16650 AND2X1_LOC_729/Y AND2X1_LOC_678/a_8_24# 0.01fF
C16651 AND2X1_LOC_572/Y OR2X1_LOC_71/Y 0.20fF
C16652 OR2X1_LOC_19/B AND2X1_LOC_823/a_8_24# 0.02fF
C16653 OR2X1_LOC_532/B OR2X1_LOC_539/Y 0.07fF
C16654 AND2X1_LOC_537/Y OR2X1_LOC_43/A 0.01fF
C16655 AND2X1_LOC_532/a_36_24# AND2X1_LOC_810/Y 0.01fF
C16656 OR2X1_LOC_246/A AND2X1_LOC_361/A 0.03fF
C16657 AND2X1_LOC_81/B D_INPUT_0 0.01fF
C16658 AND2X1_LOC_687/A OR2X1_LOC_52/B 0.26fF
C16659 AND2X1_LOC_392/A OR2X1_LOC_534/Y 0.01fF
C16660 OR2X1_LOC_197/A AND2X1_LOC_43/B 0.05fF
C16661 AND2X1_LOC_49/a_8_24# D_INPUT_0 0.03fF
C16662 OR2X1_LOC_316/Y OR2X1_LOC_75/a_8_216# 0.01fF
C16663 D_INPUT_3 OR2X1_LOC_619/Y 0.00fF
C16664 OR2X1_LOC_849/A OR2X1_LOC_62/B 0.02fF
C16665 OR2X1_LOC_3/Y AND2X1_LOC_663/B 0.05fF
C16666 OR2X1_LOC_47/Y OR2X1_LOC_427/A 1.44fF
C16667 AND2X1_LOC_807/Y AND2X1_LOC_811/Y 0.03fF
C16668 OR2X1_LOC_814/A OR2X1_LOC_68/a_8_216# 0.03fF
C16669 OR2X1_LOC_247/Y OR2X1_LOC_736/A 0.04fF
C16670 OR2X1_LOC_377/A OR2X1_LOC_84/A 0.03fF
C16671 OR2X1_LOC_76/A OR2X1_LOC_605/a_8_216# 0.01fF
C16672 AND2X1_LOC_293/a_8_24# OR2X1_LOC_44/Y 0.02fF
C16673 OR2X1_LOC_596/A OR2X1_LOC_777/B 0.72fF
C16674 AND2X1_LOC_477/A OR2X1_LOC_7/A 0.07fF
C16675 OR2X1_LOC_637/B OR2X1_LOC_598/A 0.00fF
C16676 AND2X1_LOC_303/A AND2X1_LOC_476/A 0.03fF
C16677 OR2X1_LOC_70/Y OR2X1_LOC_416/Y 0.03fF
C16678 AND2X1_LOC_42/B OR2X1_LOC_46/A 0.00fF
C16679 OR2X1_LOC_59/Y OR2X1_LOC_80/A 0.04fF
C16680 AND2X1_LOC_59/Y OR2X1_LOC_786/Y 0.21fF
C16681 OR2X1_LOC_624/B OR2X1_LOC_403/a_8_216# 0.01fF
C16682 OR2X1_LOC_140/B OR2X1_LOC_554/a_36_216# 0.02fF
C16683 OR2X1_LOC_653/A AND2X1_LOC_109/a_8_24# 0.01fF
C16684 OR2X1_LOC_185/A OR2X1_LOC_84/Y 0.10fF
C16685 OR2X1_LOC_312/Y AND2X1_LOC_863/Y 0.07fF
C16686 OR2X1_LOC_22/Y OR2X1_LOC_230/a_8_216# 0.04fF
C16687 AND2X1_LOC_369/a_8_24# OR2X1_LOC_223/A 0.01fF
C16688 AND2X1_LOC_386/a_36_24# AND2X1_LOC_7/Y 0.00fF
C16689 OR2X1_LOC_9/Y AND2X1_LOC_789/Y 0.01fF
C16690 OR2X1_LOC_427/A AND2X1_LOC_405/a_36_24# 0.01fF
C16691 OR2X1_LOC_96/B D_INPUT_1 0.33fF
C16692 AND2X1_LOC_59/Y OR2X1_LOC_644/A 0.13fF
C16693 OR2X1_LOC_756/B OR2X1_LOC_365/a_8_216# 0.01fF
C16694 VDD OR2X1_LOC_535/a_8_216# 0.21fF
C16695 OR2X1_LOC_39/A AND2X1_LOC_205/a_8_24# 0.03fF
C16696 AND2X1_LOC_70/Y OR2X1_LOC_788/B 0.00fF
C16697 D_GATE_865 D_INPUT_1 0.00fF
C16698 AND2X1_LOC_363/A OR2X1_LOC_47/Y 0.01fF
C16699 OR2X1_LOC_535/A OR2X1_LOC_356/B 0.00fF
C16700 OR2X1_LOC_447/Y OR2X1_LOC_713/a_8_216# 0.03fF
C16701 OR2X1_LOC_680/A OR2X1_LOC_419/Y 0.10fF
C16702 AND2X1_LOC_852/Y D_INPUT_1 0.04fF
C16703 OR2X1_LOC_848/A OR2X1_LOC_771/a_8_216# 0.02fF
C16704 AND2X1_LOC_364/Y OR2X1_LOC_437/A 0.01fF
C16705 OR2X1_LOC_66/A OR2X1_LOC_539/B 0.01fF
C16706 OR2X1_LOC_676/Y AND2X1_LOC_36/Y 0.09fF
C16707 OR2X1_LOC_151/A OR2X1_LOC_390/B 0.72fF
C16708 OR2X1_LOC_22/Y AND2X1_LOC_633/Y 0.03fF
C16709 AND2X1_LOC_573/A OR2X1_LOC_88/a_8_216# 0.02fF
C16710 OR2X1_LOC_770/B OR2X1_LOC_770/A 0.22fF
C16711 OR2X1_LOC_778/Y OR2X1_LOC_804/A 0.09fF
C16712 OR2X1_LOC_22/Y D_INPUT_0 0.23fF
C16713 OR2X1_LOC_188/Y OR2X1_LOC_833/Y 0.02fF
C16714 OR2X1_LOC_764/a_8_216# OR2X1_LOC_12/Y 0.01fF
C16715 AND2X1_LOC_362/B OR2X1_LOC_89/a_36_216# 0.00fF
C16716 OR2X1_LOC_143/a_8_216# OR2X1_LOC_8/Y 0.18fF
C16717 OR2X1_LOC_703/A OR2X1_LOC_788/B 0.03fF
C16718 AND2X1_LOC_544/Y AND2X1_LOC_476/Y 0.02fF
C16719 AND2X1_LOC_91/B OR2X1_LOC_307/A 0.09fF
C16720 OR2X1_LOC_217/a_8_216# OR2X1_LOC_598/A 0.02fF
C16721 OR2X1_LOC_375/A OR2X1_LOC_344/a_8_216# 0.02fF
C16722 OR2X1_LOC_158/A AND2X1_LOC_473/Y 0.10fF
C16723 OR2X1_LOC_110/a_8_216# VDD 0.21fF
C16724 AND2X1_LOC_555/Y OR2X1_LOC_604/A 0.12fF
C16725 OR2X1_LOC_181/B OR2X1_LOC_181/A 0.09fF
C16726 AND2X1_LOC_170/B AND2X1_LOC_802/a_36_24# 0.00fF
C16727 OR2X1_LOC_49/A AND2X1_LOC_415/a_8_24# 0.04fF
C16728 OR2X1_LOC_778/Y OR2X1_LOC_723/A 0.03fF
C16729 OR2X1_LOC_158/A AND2X1_LOC_287/B 0.00fF
C16730 OR2X1_LOC_600/A OR2X1_LOC_171/Y 2.75fF
C16731 OR2X1_LOC_155/A OR2X1_LOC_318/B 0.03fF
C16732 OR2X1_LOC_848/a_8_216# OR2X1_LOC_561/B 0.01fF
C16733 AND2X1_LOC_573/Y AND2X1_LOC_501/Y 0.01fF
C16734 OR2X1_LOC_736/Y OR2X1_LOC_161/B 0.03fF
C16735 OR2X1_LOC_158/A OR2X1_LOC_816/A 0.03fF
C16736 AND2X1_LOC_212/Y AND2X1_LOC_727/B 0.08fF
C16737 AND2X1_LOC_727/Y AND2X1_LOC_731/Y 0.26fF
C16738 INPUT_0 AND2X1_LOC_409/B 0.00fF
C16739 OR2X1_LOC_262/a_36_216# OR2X1_LOC_72/Y 0.01fF
C16740 OR2X1_LOC_696/A OR2X1_LOC_329/B 0.21fF
C16741 AND2X1_LOC_680/a_8_24# AND2X1_LOC_420/a_8_24# 0.23fF
C16742 OR2X1_LOC_614/Y OR2X1_LOC_161/B 0.01fF
C16743 AND2X1_LOC_573/Y AND2X1_LOC_570/Y 0.00fF
C16744 OR2X1_LOC_9/Y OR2X1_LOC_15/a_8_216# 0.05fF
C16745 INPUT_0 AND2X1_LOC_763/B 0.02fF
C16746 AND2X1_LOC_574/Y AND2X1_LOC_501/a_8_24# 0.01fF
C16747 OR2X1_LOC_47/Y AND2X1_LOC_687/B 0.07fF
C16748 OR2X1_LOC_605/A OR2X1_LOC_318/B 0.21fF
C16749 AND2X1_LOC_41/A OR2X1_LOC_130/Y 0.01fF
C16750 OR2X1_LOC_97/A OR2X1_LOC_160/B 0.12fF
C16751 OR2X1_LOC_6/A OR2X1_LOC_71/A 0.04fF
C16752 OR2X1_LOC_6/B AND2X1_LOC_256/a_8_24# 0.07fF
C16753 OR2X1_LOC_630/B OR2X1_LOC_140/B 0.00fF
C16754 OR2X1_LOC_316/Y OR2X1_LOC_13/B 0.03fF
C16755 AND2X1_LOC_423/a_36_24# OR2X1_LOC_308/Y 0.00fF
C16756 OR2X1_LOC_575/A OR2X1_LOC_500/a_8_216# 0.01fF
C16757 OR2X1_LOC_121/B OR2X1_LOC_544/a_8_216# 0.03fF
C16758 AND2X1_LOC_22/Y AND2X1_LOC_70/Y 8.99fF
C16759 AND2X1_LOC_212/A OR2X1_LOC_158/A 0.03fF
C16760 AND2X1_LOC_715/Y OR2X1_LOC_329/B 0.07fF
C16761 OR2X1_LOC_147/a_8_216# OR2X1_LOC_546/A 0.02fF
C16762 VDD INPUT_7 0.23fF
C16763 AND2X1_LOC_729/B OR2X1_LOC_761/a_8_216# 0.02fF
C16764 OR2X1_LOC_599/A OR2X1_LOC_589/a_8_216# 0.01fF
C16765 VDD OR2X1_LOC_373/Y 0.39fF
C16766 OR2X1_LOC_60/Y OR2X1_LOC_16/A 0.09fF
C16767 AND2X1_LOC_662/B OR2X1_LOC_268/Y 0.07fF
C16768 OR2X1_LOC_174/A OR2X1_LOC_174/a_8_216# 0.01fF
C16769 AND2X1_LOC_630/a_8_24# AND2X1_LOC_624/B 0.20fF
C16770 VDD OR2X1_LOC_856/A 0.06fF
C16771 OR2X1_LOC_160/B D_GATE_662 0.01fF
C16772 AND2X1_LOC_64/Y OR2X1_LOC_502/A 0.39fF
C16773 AND2X1_LOC_784/Y AND2X1_LOC_796/a_8_24# 0.11fF
C16774 OR2X1_LOC_193/Y AND2X1_LOC_41/Y 0.01fF
C16775 AND2X1_LOC_229/a_8_24# OR2X1_LOC_78/B 0.13fF
C16776 AND2X1_LOC_18/Y OR2X1_LOC_719/B 0.02fF
C16777 AND2X1_LOC_388/Y AND2X1_LOC_392/A 0.01fF
C16778 OR2X1_LOC_202/a_8_216# OR2X1_LOC_68/B 0.02fF
C16779 D_INPUT_0 OR2X1_LOC_66/Y 0.06fF
C16780 OR2X1_LOC_177/Y OR2X1_LOC_51/Y 0.03fF
C16781 OR2X1_LOC_121/Y OR2X1_LOC_78/A 0.07fF
C16782 OR2X1_LOC_462/B AND2X1_LOC_36/Y 0.03fF
C16783 AND2X1_LOC_736/Y AND2X1_LOC_564/B 0.19fF
C16784 OR2X1_LOC_74/A OR2X1_LOC_150/a_8_216# 0.14fF
C16785 OR2X1_LOC_375/A OR2X1_LOC_508/Y 0.04fF
C16786 VDD OR2X1_LOC_452/A -0.00fF
C16787 OR2X1_LOC_696/A AND2X1_LOC_113/Y 0.01fF
C16788 OR2X1_LOC_40/Y OR2X1_LOC_496/a_8_216# 0.14fF
C16789 OR2X1_LOC_528/Y AND2X1_LOC_657/Y 0.15fF
C16790 OR2X1_LOC_619/Y OR2X1_LOC_171/Y 1.75fF
C16791 AND2X1_LOC_773/Y AND2X1_LOC_857/Y 0.05fF
C16792 AND2X1_LOC_776/Y OR2X1_LOC_18/Y 0.09fF
C16793 OR2X1_LOC_227/a_36_216# AND2X1_LOC_31/Y 0.00fF
C16794 OR2X1_LOC_185/A OR2X1_LOC_556/a_8_216# 0.13fF
C16795 OR2X1_LOC_759/A OR2X1_LOC_815/a_8_216# 0.01fF
C16796 OR2X1_LOC_348/Y OR2X1_LOC_359/a_8_216# 0.05fF
C16797 OR2X1_LOC_528/Y AND2X1_LOC_191/B 0.00fF
C16798 AND2X1_LOC_390/B OR2X1_LOC_13/B 0.09fF
C16799 OR2X1_LOC_808/B OR2X1_LOC_161/B 0.10fF
C16800 OR2X1_LOC_542/B AND2X1_LOC_18/Y 0.03fF
C16801 OR2X1_LOC_604/A OR2X1_LOC_51/Y 1.48fF
C16802 AND2X1_LOC_486/Y AND2X1_LOC_244/A 0.03fF
C16803 OR2X1_LOC_509/a_8_216# OR2X1_LOC_78/B 0.03fF
C16804 OR2X1_LOC_51/Y AND2X1_LOC_207/B 0.13fF
C16805 OR2X1_LOC_494/A OR2X1_LOC_625/Y 0.01fF
C16806 AND2X1_LOC_388/Y AND2X1_LOC_436/a_8_24# 0.10fF
C16807 OR2X1_LOC_314/a_8_216# OR2X1_LOC_16/A 0.05fF
C16808 OR2X1_LOC_186/Y AND2X1_LOC_40/Y 0.49fF
C16809 OR2X1_LOC_114/B OR2X1_LOC_78/A 0.04fF
C16810 OR2X1_LOC_614/Y AND2X1_LOC_48/a_8_24# 0.01fF
C16811 OR2X1_LOC_519/Y AND2X1_LOC_520/a_8_24# 0.01fF
C16812 AND2X1_LOC_285/Y AND2X1_LOC_286/a_8_24# 0.11fF
C16813 AND2X1_LOC_91/B AND2X1_LOC_394/a_8_24# 0.01fF
C16814 OR2X1_LOC_611/a_36_216# OR2X1_LOC_71/A 0.00fF
C16815 OR2X1_LOC_681/a_8_216# OR2X1_LOC_91/A 0.01fF
C16816 OR2X1_LOC_132/Y VDD 0.17fF
C16817 OR2X1_LOC_318/Y OR2X1_LOC_435/A 0.04fF
C16818 AND2X1_LOC_738/B OR2X1_LOC_331/A 0.13fF
C16819 OR2X1_LOC_78/B OR2X1_LOC_66/A 10.24fF
C16820 OR2X1_LOC_176/Y AND2X1_LOC_593/Y 0.03fF
C16821 OR2X1_LOC_160/B OR2X1_LOC_541/A 0.02fF
C16822 AND2X1_LOC_347/a_36_24# AND2X1_LOC_789/Y 0.01fF
C16823 AND2X1_LOC_550/a_8_24# OR2X1_LOC_524/Y 0.03fF
C16824 AND2X1_LOC_654/B OR2X1_LOC_13/Y 0.02fF
C16825 AND2X1_LOC_364/Y AND2X1_LOC_715/A 0.03fF
C16826 AND2X1_LOC_744/a_8_24# OR2X1_LOC_160/B 0.01fF
C16827 OR2X1_LOC_326/a_8_216# AND2X1_LOC_70/Y 0.05fF
C16828 OR2X1_LOC_316/a_8_216# OR2X1_LOC_52/B 0.02fF
C16829 OR2X1_LOC_744/A OR2X1_LOC_666/A 0.03fF
C16830 OR2X1_LOC_461/a_8_216# INPUT_0 0.01fF
C16831 AND2X1_LOC_722/Y VDD 0.21fF
C16832 AND2X1_LOC_561/a_36_24# OR2X1_LOC_89/A 0.00fF
C16833 AND2X1_LOC_92/Y AND2X1_LOC_628/a_8_24# 0.02fF
C16834 AND2X1_LOC_70/Y OR2X1_LOC_244/B 0.02fF
C16835 OR2X1_LOC_533/Y AND2X1_LOC_593/Y 0.11fF
C16836 AND2X1_LOC_716/Y OR2X1_LOC_309/Y 0.03fF
C16837 AND2X1_LOC_713/Y OR2X1_LOC_92/Y 0.01fF
C16838 VDD AND2X1_LOC_401/Y 0.38fF
C16839 AND2X1_LOC_59/Y AND2X1_LOC_255/a_8_24# 0.01fF
C16840 OR2X1_LOC_691/a_8_216# OR2X1_LOC_377/A 0.02fF
C16841 AND2X1_LOC_219/Y AND2X1_LOC_222/a_8_24# 0.01fF
C16842 AND2X1_LOC_456/B AND2X1_LOC_658/A 0.03fF
C16843 OR2X1_LOC_538/A OR2X1_LOC_78/A 0.03fF
C16844 AND2X1_LOC_64/Y AND2X1_LOC_72/a_8_24# 0.01fF
C16845 OR2X1_LOC_329/B AND2X1_LOC_851/a_36_24# 0.01fF
C16846 OR2X1_LOC_659/Y OR2X1_LOC_659/a_8_216# 0.00fF
C16847 AND2X1_LOC_486/Y OR2X1_LOC_108/Y 0.07fF
C16848 AND2X1_LOC_228/Y OR2X1_LOC_12/Y 0.03fF
C16849 VDD OR2X1_LOC_426/A 0.08fF
C16850 OR2X1_LOC_721/Y OR2X1_LOC_66/A 0.01fF
C16851 AND2X1_LOC_866/B OR2X1_LOC_627/Y 0.02fF
C16852 OR2X1_LOC_309/a_8_216# AND2X1_LOC_662/B 0.04fF
C16853 AND2X1_LOC_14/a_8_24# OR2X1_LOC_80/A 0.02fF
C16854 OR2X1_LOC_744/A OR2X1_LOC_762/Y 0.26fF
C16855 AND2X1_LOC_59/Y OR2X1_LOC_535/A 0.01fF
C16856 AND2X1_LOC_550/A AND2X1_LOC_476/Y 0.02fF
C16857 OR2X1_LOC_243/A OR2X1_LOC_549/A 0.03fF
C16858 AND2X1_LOC_539/Y AND2X1_LOC_356/B 0.55fF
C16859 AND2X1_LOC_784/A OR2X1_LOC_310/a_8_216# 0.04fF
C16860 OR2X1_LOC_185/A OR2X1_LOC_565/A 6.13fF
C16861 OR2X1_LOC_448/a_8_216# OR2X1_LOC_66/A 0.01fF
C16862 INPUT_0 OR2X1_LOC_634/A 0.09fF
C16863 AND2X1_LOC_95/Y OR2X1_LOC_362/A 0.49fF
C16864 OR2X1_LOC_326/a_8_216# OR2X1_LOC_703/A 0.01fF
C16865 OR2X1_LOC_768/A OR2X1_LOC_663/A 0.03fF
C16866 OR2X1_LOC_177/Y OR2X1_LOC_680/A 0.03fF
C16867 AND2X1_LOC_22/Y AND2X1_LOC_17/Y 0.29fF
C16868 OR2X1_LOC_415/A OR2X1_LOC_395/Y 0.00fF
C16869 AND2X1_LOC_552/a_8_24# OR2X1_LOC_280/Y 0.03fF
C16870 OR2X1_LOC_858/A OR2X1_LOC_840/A 0.09fF
C16871 OR2X1_LOC_139/A OR2X1_LOC_139/a_8_216# 0.08fF
C16872 AND2X1_LOC_3/Y OR2X1_LOC_267/Y 0.03fF
C16873 OR2X1_LOC_389/B AND2X1_LOC_44/Y 0.09fF
C16874 OR2X1_LOC_405/A AND2X1_LOC_110/Y 0.03fF
C16875 OR2X1_LOC_97/A OR2X1_LOC_219/B 0.03fF
C16876 OR2X1_LOC_524/Y AND2X1_LOC_545/a_36_24# 0.01fF
C16877 AND2X1_LOC_545/a_8_24# AND2X1_LOC_551/B 0.00fF
C16878 OR2X1_LOC_693/Y OR2X1_LOC_44/Y 0.01fF
C16879 AND2X1_LOC_40/a_8_24# AND2X1_LOC_25/Y 0.14fF
C16880 AND2X1_LOC_716/Y OR2X1_LOC_744/A 0.07fF
C16881 AND2X1_LOC_624/A AND2X1_LOC_254/a_8_24# 0.02fF
C16882 OR2X1_LOC_168/a_8_216# OR2X1_LOC_468/A 0.01fF
C16883 OR2X1_LOC_805/A OR2X1_LOC_723/a_8_216# 0.04fF
C16884 AND2X1_LOC_703/Y OR2X1_LOC_7/A 0.12fF
C16885 OR2X1_LOC_585/A OR2X1_LOC_12/Y 0.19fF
C16886 OR2X1_LOC_185/A OR2X1_LOC_190/Y 0.02fF
C16887 OR2X1_LOC_154/A OR2X1_LOC_648/B 0.10fF
C16888 OR2X1_LOC_3/Y OR2X1_LOC_18/a_8_216# 0.01fF
C16889 OR2X1_LOC_281/a_8_216# OR2X1_LOC_59/Y 0.03fF
C16890 OR2X1_LOC_851/A OR2X1_LOC_168/B 0.06fF
C16891 OR2X1_LOC_485/A AND2X1_LOC_242/a_36_24# 0.00fF
C16892 OR2X1_LOC_502/A AND2X1_LOC_819/a_8_24# 0.03fF
C16893 OR2X1_LOC_158/A OR2X1_LOC_824/Y 0.07fF
C16894 OR2X1_LOC_51/Y OR2X1_LOC_252/a_8_216# 0.01fF
C16895 OR2X1_LOC_604/A OR2X1_LOC_680/A 0.07fF
C16896 AND2X1_LOC_47/Y OR2X1_LOC_593/B 0.05fF
C16897 OR2X1_LOC_532/B OR2X1_LOC_523/a_36_216# 0.00fF
C16898 OR2X1_LOC_43/A OR2X1_LOC_13/Y 0.05fF
C16899 AND2X1_LOC_81/B AND2X1_LOC_505/a_8_24# 0.01fF
C16900 AND2X1_LOC_758/a_8_24# OR2X1_LOC_680/A 0.02fF
C16901 AND2X1_LOC_392/A AND2X1_LOC_572/A 0.03fF
C16902 AND2X1_LOC_33/a_8_24# AND2X1_LOC_33/Y 0.00fF
C16903 OR2X1_LOC_371/Y AND2X1_LOC_786/Y 0.07fF
C16904 OR2X1_LOC_375/A OR2X1_LOC_66/A 0.36fF
C16905 VDD INPUT_4 0.04fF
C16906 OR2X1_LOC_51/Y AND2X1_LOC_467/a_8_24# 0.01fF
C16907 OR2X1_LOC_754/Y AND2X1_LOC_790/a_8_24# 0.23fF
C16908 OR2X1_LOC_160/A OR2X1_LOC_648/A 0.07fF
C16909 OR2X1_LOC_670/a_8_216# OR2X1_LOC_96/Y 0.01fF
C16910 OR2X1_LOC_532/B OR2X1_LOC_319/Y 0.01fF
C16911 OR2X1_LOC_512/A OR2X1_LOC_502/A 0.00fF
C16912 AND2X1_LOC_64/Y AND2X1_LOC_48/A 0.13fF
C16913 OR2X1_LOC_528/Y AND2X1_LOC_862/a_8_24# 0.17fF
C16914 OR2X1_LOC_377/A AND2X1_LOC_94/Y 0.46fF
C16915 AND2X1_LOC_123/Y OR2X1_LOC_56/A 0.01fF
C16916 AND2X1_LOC_56/B AND2X1_LOC_18/Y 1.46fF
C16917 AND2X1_LOC_22/Y OR2X1_LOC_404/Y 0.02fF
C16918 AND2X1_LOC_12/Y OR2X1_LOC_78/A 0.10fF
C16919 OR2X1_LOC_711/B OR2X1_LOC_711/A 0.48fF
C16920 AND2X1_LOC_593/a_36_24# OR2X1_LOC_36/Y 0.01fF
C16921 OR2X1_LOC_516/A AND2X1_LOC_469/B 0.01fF
C16922 OR2X1_LOC_482/a_36_216# OR2X1_LOC_7/A 0.03fF
C16923 AND2X1_LOC_539/Y OR2X1_LOC_22/Y 0.07fF
C16924 OR2X1_LOC_475/a_36_216# OR2X1_LOC_475/B 0.01fF
C16925 AND2X1_LOC_719/Y OR2X1_LOC_238/Y 0.20fF
C16926 OR2X1_LOC_64/Y OR2X1_LOC_764/a_36_216# 0.00fF
C16927 OR2X1_LOC_309/Y OR2X1_LOC_312/Y 0.03fF
C16928 AND2X1_LOC_8/Y AND2X1_LOC_18/Y 0.04fF
C16929 OR2X1_LOC_771/B D_INPUT_1 0.02fF
C16930 OR2X1_LOC_810/a_8_216# OR2X1_LOC_862/A 0.41fF
C16931 OR2X1_LOC_409/B OR2X1_LOC_387/A 0.16fF
C16932 OR2X1_LOC_58/Y OR2X1_LOC_690/A 0.01fF
C16933 AND2X1_LOC_12/Y OR2X1_LOC_850/a_8_216# 0.00fF
C16934 OR2X1_LOC_149/B OR2X1_LOC_471/Y 0.12fF
C16935 AND2X1_LOC_546/a_8_24# OR2X1_LOC_677/Y 0.10fF
C16936 INPUT_0 OR2X1_LOC_94/a_8_216# 0.01fF
C16937 OR2X1_LOC_114/a_36_216# OR2X1_LOC_161/A 0.00fF
C16938 AND2X1_LOC_64/Y AND2X1_LOC_69/a_36_24# 0.01fF
C16939 OR2X1_LOC_154/A AND2X1_LOC_103/a_8_24# -0.04fF
C16940 OR2X1_LOC_625/a_8_216# OR2X1_LOC_92/Y 0.02fF
C16941 AND2X1_LOC_95/Y OR2X1_LOC_474/Y 0.05fF
C16942 D_INPUT_5 OR2X1_LOC_30/a_8_216# 0.01fF
C16943 VDD AND2X1_LOC_51/A 0.37fF
C16944 AND2X1_LOC_599/a_8_24# AND2X1_LOC_48/A 0.02fF
C16945 OR2X1_LOC_161/A OR2X1_LOC_708/Y 0.03fF
C16946 OR2X1_LOC_6/A OR2X1_LOC_59/Y 0.07fF
C16947 AND2X1_LOC_13/a_8_24# OR2X1_LOC_596/A 0.09fF
C16948 AND2X1_LOC_47/Y AND2X1_LOC_273/a_8_24# 0.02fF
C16949 OR2X1_LOC_132/a_8_216# OR2X1_LOC_26/Y 0.01fF
C16950 AND2X1_LOC_117/a_36_24# AND2X1_LOC_65/A 0.00fF
C16951 OR2X1_LOC_62/B OR2X1_LOC_572/a_8_216# 0.01fF
C16952 OR2X1_LOC_176/a_8_216# AND2X1_LOC_477/A 0.01fF
C16953 OR2X1_LOC_34/B OR2X1_LOC_34/a_8_216# 0.47fF
C16954 OR2X1_LOC_777/B OR2X1_LOC_374/Y 0.03fF
C16955 AND2X1_LOC_40/a_8_24# AND2X1_LOC_51/Y 0.01fF
C16956 OR2X1_LOC_864/A OR2X1_LOC_35/Y 0.03fF
C16957 OR2X1_LOC_164/Y OR2X1_LOC_39/A 0.01fF
C16958 AND2X1_LOC_706/Y OR2X1_LOC_64/Y 0.00fF
C16959 OR2X1_LOC_696/A OR2X1_LOC_618/Y 0.01fF
C16960 AND2X1_LOC_163/a_8_24# AND2X1_LOC_51/Y 0.01fF
C16961 AND2X1_LOC_392/A OR2X1_LOC_3/Y 0.03fF
C16962 AND2X1_LOC_12/Y OR2X1_LOC_448/B 0.18fF
C16963 AND2X1_LOC_720/a_8_24# OR2X1_LOC_427/A 0.04fF
C16964 OR2X1_LOC_820/A OR2X1_LOC_44/Y 0.01fF
C16965 OR2X1_LOC_264/Y OR2X1_LOC_340/Y 0.00fF
C16966 AND2X1_LOC_110/a_8_24# AND2X1_LOC_3/Y 0.02fF
C16967 OR2X1_LOC_625/Y OR2X1_LOC_427/A 0.28fF
C16968 OR2X1_LOC_527/a_8_216# OR2X1_LOC_527/Y 0.03fF
C16969 OR2X1_LOC_744/A OR2X1_LOC_312/Y 0.06fF
C16970 AND2X1_LOC_634/Y OR2X1_LOC_12/Y 0.13fF
C16971 OR2X1_LOC_851/A AND2X1_LOC_59/Y 0.01fF
C16972 OR2X1_LOC_759/A OR2X1_LOC_617/Y 0.03fF
C16973 OR2X1_LOC_175/Y OR2X1_LOC_436/Y 0.13fF
C16974 AND2X1_LOC_40/Y AND2X1_LOC_81/B 0.05fF
C16975 OR2X1_LOC_563/a_8_216# OR2X1_LOC_563/B 0.06fF
C16976 AND2X1_LOC_378/a_36_24# OR2X1_LOC_43/A 0.01fF
C16977 OR2X1_LOC_538/A OR2X1_LOC_155/A 0.03fF
C16978 OR2X1_LOC_158/A AND2X1_LOC_727/A 0.03fF
C16979 OR2X1_LOC_849/A OR2X1_LOC_659/A 0.15fF
C16980 OR2X1_LOC_687/Y OR2X1_LOC_623/B 0.33fF
C16981 AND2X1_LOC_40/Y OR2X1_LOC_358/B 0.26fF
C16982 OR2X1_LOC_739/B OR2X1_LOC_220/B 0.14fF
C16983 AND2X1_LOC_465/a_8_24# OR2X1_LOC_59/Y 0.01fF
C16984 AND2X1_LOC_651/a_8_24# OR2X1_LOC_44/Y 0.01fF
C16985 OR2X1_LOC_691/A OR2X1_LOC_532/B 0.00fF
C16986 OR2X1_LOC_185/A OR2X1_LOC_161/A 0.09fF
C16987 OR2X1_LOC_485/A INPUT_0 1.06fF
C16988 OR2X1_LOC_196/B OR2X1_LOC_515/A 0.09fF
C16989 AND2X1_LOC_473/a_8_24# OR2X1_LOC_56/A 0.05fF
C16990 OR2X1_LOC_9/Y OR2X1_LOC_246/A 0.14fF
C16991 OR2X1_LOC_680/Y AND2X1_LOC_663/A 0.05fF
C16992 AND2X1_LOC_266/a_36_24# AND2X1_LOC_266/Y 0.02fF
C16993 OR2X1_LOC_52/B OR2X1_LOC_746/a_8_216# 0.02fF
C16994 OR2X1_LOC_436/Y AND2X1_LOC_417/a_8_24# 0.01fF
C16995 OR2X1_LOC_40/Y AND2X1_LOC_465/Y 0.02fF
C16996 AND2X1_LOC_724/A OR2X1_LOC_31/Y 0.01fF
C16997 VDD AND2X1_LOC_849/A 0.38fF
C16998 AND2X1_LOC_728/Y AND2X1_LOC_729/Y 0.42fF
C16999 OR2X1_LOC_179/a_36_216# OR2X1_LOC_529/Y 0.00fF
C17000 AND2X1_LOC_841/B AND2X1_LOC_661/A 0.03fF
C17001 OR2X1_LOC_643/A OR2X1_LOC_231/A 0.03fF
C17002 VDD OR2X1_LOC_268/a_8_216# 0.21fF
C17003 AND2X1_LOC_91/B OR2X1_LOC_804/A 0.10fF
C17004 AND2X1_LOC_372/a_8_24# OR2X1_LOC_778/A 0.08fF
C17005 OR2X1_LOC_270/a_8_216# OR2X1_LOC_456/a_8_216# 0.47fF
C17006 AND2X1_LOC_182/a_8_24# OR2X1_LOC_417/A 0.04fF
C17007 OR2X1_LOC_247/a_8_216# OR2X1_LOC_563/A 0.02fF
C17008 OR2X1_LOC_773/B OR2X1_LOC_848/A 0.01fF
C17009 OR2X1_LOC_168/a_8_216# OR2X1_LOC_449/B 0.01fF
C17010 OR2X1_LOC_158/A OR2X1_LOC_95/Y 3.15fF
C17011 AND2X1_LOC_621/Y OR2X1_LOC_44/Y 0.03fF
C17012 AND2X1_LOC_59/Y OR2X1_LOC_204/Y 0.04fF
C17013 AND2X1_LOC_363/A OR2X1_LOC_625/Y 0.01fF
C17014 AND2X1_LOC_387/a_8_24# D_INPUT_0 0.01fF
C17015 OR2X1_LOC_85/A OR2X1_LOC_265/Y 0.06fF
C17016 OR2X1_LOC_569/B OR2X1_LOC_549/Y 0.70fF
C17017 OR2X1_LOC_814/A OR2X1_LOC_244/Y 0.02fF
C17018 AND2X1_LOC_228/Y AND2X1_LOC_650/Y 0.46fF
C17019 OR2X1_LOC_47/Y OR2X1_LOC_322/a_8_216# 0.01fF
C17020 OR2X1_LOC_298/Y OR2X1_LOC_52/B 0.02fF
C17021 OR2X1_LOC_643/A OR2X1_LOC_130/A 0.07fF
C17022 AND2X1_LOC_12/Y OR2X1_LOC_155/A 0.06fF
C17023 AND2X1_LOC_795/Y OR2X1_LOC_373/a_36_216# 0.03fF
C17024 OR2X1_LOC_585/A OR2X1_LOC_38/a_36_216# 0.00fF
C17025 OR2X1_LOC_651/a_8_216# OR2X1_LOC_375/A 0.01fF
C17026 AND2X1_LOC_817/B OR2X1_LOC_847/B 0.01fF
C17027 AND2X1_LOC_702/Y AND2X1_LOC_303/B 0.00fF
C17028 OR2X1_LOC_596/Y AND2X1_LOC_56/B 0.01fF
C17029 AND2X1_LOC_76/Y AND2X1_LOC_660/Y 0.00fF
C17030 OR2X1_LOC_79/A OR2X1_LOC_18/Y 0.15fF
C17031 OR2X1_LOC_6/A OR2X1_LOC_820/B 0.03fF
C17032 OR2X1_LOC_702/A OR2X1_LOC_624/A 0.05fF
C17033 OR2X1_LOC_290/Y AND2X1_LOC_334/a_8_24# -0.00fF
C17034 OR2X1_LOC_415/Y OR2X1_LOC_68/B 0.04fF
C17035 OR2X1_LOC_714/a_8_216# OR2X1_LOC_317/B 0.16fF
C17036 OR2X1_LOC_175/Y OR2X1_LOC_566/Y 0.09fF
C17037 OR2X1_LOC_280/Y OR2X1_LOC_237/a_8_216# 0.01fF
C17038 OR2X1_LOC_755/A AND2X1_LOC_846/a_36_24# 0.00fF
C17039 AND2X1_LOC_256/a_8_24# OR2X1_LOC_598/A 0.01fF
C17040 OR2X1_LOC_369/Y AND2X1_LOC_866/A 0.14fF
C17041 OR2X1_LOC_503/A OR2X1_LOC_485/A 0.01fF
C17042 OR2X1_LOC_132/Y OR2X1_LOC_256/A 0.08fF
C17043 OR2X1_LOC_520/Y AND2X1_LOC_3/Y 0.09fF
C17044 AND2X1_LOC_155/Y OR2X1_LOC_39/A 0.01fF
C17045 OR2X1_LOC_223/A OR2X1_LOC_776/Y 0.01fF
C17046 OR2X1_LOC_22/Y AND2X1_LOC_276/a_8_24# 0.01fF
C17047 AND2X1_LOC_120/a_36_24# AND2X1_LOC_850/Y 0.01fF
C17048 AND2X1_LOC_54/a_36_24# INPUT_1 0.01fF
C17049 AND2X1_LOC_727/A OR2X1_LOC_594/Y 0.01fF
C17050 OR2X1_LOC_841/B OR2X1_LOC_155/A 0.01fF
C17051 OR2X1_LOC_91/A AND2X1_LOC_656/Y 2.01fF
C17052 OR2X1_LOC_496/Y AND2X1_LOC_778/a_8_24# 0.11fF
C17053 OR2X1_LOC_151/A OR2X1_LOC_493/Y 0.10fF
C17054 OR2X1_LOC_185/A AND2X1_LOC_51/Y 0.04fF
C17055 AND2X1_LOC_222/Y AND2X1_LOC_786/Y 0.04fF
C17056 AND2X1_LOC_34/Y OR2X1_LOC_27/Y 0.01fF
C17057 AND2X1_LOC_339/a_8_24# OR2X1_LOC_26/Y 0.04fF
C17058 AND2X1_LOC_95/Y AND2X1_LOC_680/a_8_24# 0.01fF
C17059 OR2X1_LOC_19/B OR2X1_LOC_414/a_8_216# 0.06fF
C17060 AND2X1_LOC_131/a_8_24# OR2X1_LOC_66/Y 0.01fF
C17061 OR2X1_LOC_476/B OR2X1_LOC_624/A 0.01fF
C17062 AND2X1_LOC_855/a_8_24# AND2X1_LOC_655/A 0.27fF
C17063 OR2X1_LOC_70/Y OR2X1_LOC_6/A 0.03fF
C17064 AND2X1_LOC_168/a_8_24# OR2X1_LOC_417/A 0.04fF
C17065 AND2X1_LOC_784/A AND2X1_LOC_568/a_36_24# 0.01fF
C17066 OR2X1_LOC_103/Y OR2X1_LOC_95/Y 1.03fF
C17067 OR2X1_LOC_289/a_8_216# OR2X1_LOC_59/Y 0.06fF
C17068 OR2X1_LOC_764/Y AND2X1_LOC_769/a_8_24# 0.23fF
C17069 OR2X1_LOC_811/A OR2X1_LOC_532/B 0.02fF
C17070 OR2X1_LOC_756/B OR2X1_LOC_223/A 0.02fF
C17071 OR2X1_LOC_646/a_8_216# OR2X1_LOC_647/B 0.01fF
C17072 OR2X1_LOC_816/Y AND2X1_LOC_792/Y 0.01fF
C17073 OR2X1_LOC_269/B OR2X1_LOC_705/Y 0.02fF
C17074 OR2X1_LOC_52/B OR2X1_LOC_27/a_8_216# 0.03fF
C17075 AND2X1_LOC_660/Y OR2X1_LOC_52/B 0.05fF
C17076 AND2X1_LOC_633/Y OR2X1_LOC_39/A 0.03fF
C17077 AND2X1_LOC_197/a_8_24# OR2X1_LOC_753/A 0.17fF
C17078 AND2X1_LOC_654/Y OR2X1_LOC_31/Y 0.01fF
C17079 OR2X1_LOC_811/A AND2X1_LOC_665/a_8_24# 0.03fF
C17080 OR2X1_LOC_26/Y AND2X1_LOC_523/Y 0.03fF
C17081 AND2X1_LOC_514/Y OR2X1_LOC_6/A 0.01fF
C17082 OR2X1_LOC_18/Y OR2X1_LOC_226/a_36_216# 0.03fF
C17083 OR2X1_LOC_323/A OR2X1_LOC_268/Y 0.70fF
C17084 OR2X1_LOC_103/a_8_216# OR2X1_LOC_95/Y 0.01fF
C17085 OR2X1_LOC_673/Y OR2X1_LOC_19/B 0.15fF
C17086 AND2X1_LOC_773/Y OR2X1_LOC_437/A 0.10fF
C17087 OR2X1_LOC_56/A OR2X1_LOC_406/A 0.29fF
C17088 D_INPUT_0 OR2X1_LOC_39/A 0.10fF
C17089 AND2X1_LOC_578/A OR2X1_LOC_371/Y 0.07fF
C17090 AND2X1_LOC_216/Y AND2X1_LOC_216/a_8_24# 0.00fF
C17091 OR2X1_LOC_264/Y AND2X1_LOC_88/Y 0.02fF
C17092 AND2X1_LOC_40/Y OR2X1_LOC_112/B 0.02fF
C17093 OR2X1_LOC_404/a_8_216# OR2X1_LOC_532/B 0.01fF
C17094 OR2X1_LOC_417/Y AND2X1_LOC_454/A 0.01fF
C17095 AND2X1_LOC_656/Y AND2X1_LOC_573/A 0.03fF
C17096 AND2X1_LOC_523/Y OR2X1_LOC_89/A 0.02fF
C17097 AND2X1_LOC_392/A AND2X1_LOC_772/a_8_24# 0.06fF
C17098 OR2X1_LOC_46/A AND2X1_LOC_412/a_8_24# 0.02fF
C17099 AND2X1_LOC_63/a_8_24# OR2X1_LOC_244/A 0.02fF
C17100 OR2X1_LOC_255/a_8_216# OR2X1_LOC_85/A 0.02fF
C17101 OR2X1_LOC_643/A OR2X1_LOC_62/B 0.03fF
C17102 OR2X1_LOC_829/A OR2X1_LOC_536/a_8_216# 0.28fF
C17103 OR2X1_LOC_485/A OR2X1_LOC_64/Y 5.80fF
C17104 OR2X1_LOC_62/B OR2X1_LOC_124/Y 0.00fF
C17105 AND2X1_LOC_671/a_8_24# OR2X1_LOC_585/A 0.23fF
C17106 AND2X1_LOC_303/A OR2X1_LOC_417/A 0.00fF
C17107 OR2X1_LOC_651/A AND2X1_LOC_43/B 0.01fF
C17108 OR2X1_LOC_596/A OR2X1_LOC_704/a_36_216# 0.00fF
C17109 OR2X1_LOC_707/B OR2X1_LOC_449/B 0.01fF
C17110 OR2X1_LOC_524/Y AND2X1_LOC_222/Y 0.05fF
C17111 AND2X1_LOC_180/a_36_24# OR2X1_LOC_437/A 0.01fF
C17112 OR2X1_LOC_286/B OR2X1_LOC_269/B 0.35fF
C17113 VDD OR2X1_LOC_725/a_8_216# 0.00fF
C17114 OR2X1_LOC_439/B OR2X1_LOC_544/B 0.49fF
C17115 OR2X1_LOC_308/a_8_216# OR2X1_LOC_512/a_8_216# 0.47fF
C17116 OR2X1_LOC_833/B AND2X1_LOC_271/a_8_24# 0.01fF
C17117 OR2X1_LOC_89/A OR2X1_LOC_815/A 0.01fF
C17118 AND2X1_LOC_434/Y OR2X1_LOC_172/Y 0.01fF
C17119 AND2X1_LOC_171/a_8_24# OR2X1_LOC_814/A 0.01fF
C17120 AND2X1_LOC_243/Y OR2X1_LOC_437/A 0.07fF
C17121 OR2X1_LOC_151/A OR2X1_LOC_532/a_8_216# 0.06fF
C17122 AND2X1_LOC_512/Y OR2X1_LOC_761/a_36_216# 0.00fF
C17123 OR2X1_LOC_574/a_8_216# OR2X1_LOC_598/A 0.02fF
C17124 OR2X1_LOC_402/Y D_INPUT_1 0.19fF
C17125 AND2X1_LOC_801/B OR2X1_LOC_585/A 0.01fF
C17126 OR2X1_LOC_632/Y OR2X1_LOC_68/B 0.09fF
C17127 AND2X1_LOC_211/B D_INPUT_0 0.40fF
C17128 OR2X1_LOC_287/B AND2X1_LOC_283/a_8_24# 0.01fF
C17129 OR2X1_LOC_843/a_8_216# OR2X1_LOC_814/A 0.01fF
C17130 OR2X1_LOC_574/A D_INPUT_0 0.03fF
C17131 AND2X1_LOC_324/a_8_24# AND2X1_LOC_863/A 0.11fF
C17132 AND2X1_LOC_83/a_8_24# AND2X1_LOC_36/Y 0.01fF
C17133 OR2X1_LOC_377/A OR2X1_LOC_214/B 0.12fF
C17134 OR2X1_LOC_312/Y OR2X1_LOC_31/Y 0.00fF
C17135 OR2X1_LOC_840/A AND2X1_LOC_31/Y 0.03fF
C17136 OR2X1_LOC_485/A OR2X1_LOC_417/A 0.12fF
C17137 AND2X1_LOC_8/Y AND2X1_LOC_672/a_8_24# 0.01fF
C17138 OR2X1_LOC_291/Y AND2X1_LOC_334/a_8_24# 0.11fF
C17139 AND2X1_LOC_722/A OR2X1_LOC_533/A 0.05fF
C17140 OR2X1_LOC_375/A OR2X1_LOC_98/B 0.09fF
C17141 AND2X1_LOC_192/Y OR2X1_LOC_747/Y 0.02fF
C17142 AND2X1_LOC_348/a_8_24# OR2X1_LOC_417/A 0.01fF
C17143 OR2X1_LOC_809/B OR2X1_LOC_112/A 0.23fF
C17144 OR2X1_LOC_488/a_36_216# OR2X1_LOC_71/Y -0.00fF
C17145 AND2X1_LOC_721/Y AND2X1_LOC_287/B 0.05fF
C17146 AND2X1_LOC_465/A AND2X1_LOC_455/B 0.83fF
C17147 OR2X1_LOC_472/B OR2X1_LOC_46/A 0.07fF
C17148 OR2X1_LOC_744/A OR2X1_LOC_13/B 0.17fF
C17149 OR2X1_LOC_748/A AND2X1_LOC_792/Y 0.14fF
C17150 OR2X1_LOC_516/Y OR2X1_LOC_40/Y 0.07fF
C17151 AND2X1_LOC_43/B OR2X1_LOC_728/B 0.01fF
C17152 OR2X1_LOC_311/Y AND2X1_LOC_539/a_8_24# 0.01fF
C17153 OR2X1_LOC_85/A AND2X1_LOC_205/a_8_24# 0.01fF
C17154 OR2X1_LOC_576/A OR2X1_LOC_474/B 0.15fF
C17155 AND2X1_LOC_100/a_8_24# OR2X1_LOC_67/Y 0.01fF
C17156 AND2X1_LOC_739/B VDD 0.13fF
C17157 AND2X1_LOC_538/Y AND2X1_LOC_539/a_8_24# 0.19fF
C17158 OR2X1_LOC_230/Y OR2X1_LOC_12/Y 0.21fF
C17159 AND2X1_LOC_672/B D_INPUT_0 0.15fF
C17160 OR2X1_LOC_121/B OR2X1_LOC_440/A 0.03fF
C17161 OR2X1_LOC_778/Y OR2X1_LOC_365/B 0.05fF
C17162 AND2X1_LOC_150/a_8_24# OR2X1_LOC_392/B 0.12fF
C17163 OR2X1_LOC_677/a_8_216# OR2X1_LOC_142/Y 0.18fF
C17164 AND2X1_LOC_90/a_8_24# AND2X1_LOC_277/a_8_24# 0.23fF
C17165 AND2X1_LOC_707/Y AND2X1_LOC_714/B 0.07fF
C17166 OR2X1_LOC_64/Y AND2X1_LOC_645/a_36_24# 0.00fF
C17167 OR2X1_LOC_229/a_8_216# OR2X1_LOC_12/Y 0.01fF
C17168 OR2X1_LOC_78/B OR2X1_LOC_502/a_8_216# 0.05fF
C17169 OR2X1_LOC_482/Y OR2X1_LOC_816/A 10.04fF
C17170 AND2X1_LOC_22/Y OR2X1_LOC_362/A 0.07fF
C17171 AND2X1_LOC_22/Y AND2X1_LOC_511/a_36_24# 0.00fF
C17172 OR2X1_LOC_175/Y OR2X1_LOC_160/B 0.30fF
C17173 OR2X1_LOC_596/A OR2X1_LOC_161/B 0.06fF
C17174 OR2X1_LOC_596/a_8_216# AND2X1_LOC_44/Y 0.16fF
C17175 OR2X1_LOC_186/Y OR2X1_LOC_356/A 0.01fF
C17176 OR2X1_LOC_562/a_8_216# OR2X1_LOC_562/A 0.18fF
C17177 OR2X1_LOC_866/B VDD 0.08fF
C17178 OR2X1_LOC_6/B AND2X1_LOC_44/Y 11.35fF
C17179 OR2X1_LOC_160/A OR2X1_LOC_501/a_36_216# 0.01fF
C17180 OR2X1_LOC_59/Y AND2X1_LOC_792/a_36_24# 0.00fF
C17181 VDD AND2X1_LOC_60/a_8_24# -0.00fF
C17182 OR2X1_LOC_91/A AND2X1_LOC_772/Y 0.07fF
C17183 AND2X1_LOC_654/Y OR2X1_LOC_320/a_8_216# 0.03fF
C17184 AND2X1_LOC_95/Y OR2X1_LOC_771/B 0.03fF
C17185 OR2X1_LOC_160/A OR2X1_LOC_730/B 0.28fF
C17186 OR2X1_LOC_160/B OR2X1_LOC_691/Y 0.03fF
C17187 OR2X1_LOC_333/B OR2X1_LOC_228/Y 0.16fF
C17188 OR2X1_LOC_417/A AND2X1_LOC_655/a_8_24# 0.02fF
C17189 INPUT_1 AND2X1_LOC_837/a_8_24# 0.01fF
C17190 AND2X1_LOC_578/A AND2X1_LOC_222/Y 0.03fF
C17191 OR2X1_LOC_596/A OR2X1_LOC_514/a_36_216# 0.00fF
C17192 OR2X1_LOC_240/A OR2X1_LOC_80/A 0.08fF
C17193 VDD OR2X1_LOC_759/a_8_216# 0.21fF
C17194 OR2X1_LOC_176/Y OR2X1_LOC_51/Y 0.04fF
C17195 OR2X1_LOC_579/B OR2X1_LOC_580/A 0.01fF
C17196 OR2X1_LOC_633/B OR2X1_LOC_80/A 0.00fF
C17197 OR2X1_LOC_737/A OR2X1_LOC_776/A 0.07fF
C17198 OR2X1_LOC_362/A OR2X1_LOC_343/a_36_216# 0.00fF
C17199 OR2X1_LOC_506/A OR2X1_LOC_593/B 0.02fF
C17200 AND2X1_LOC_20/a_8_24# AND2X1_LOC_7/B 0.01fF
C17201 AND2X1_LOC_64/Y OR2X1_LOC_201/A 0.01fF
C17202 AND2X1_LOC_207/a_8_24# OR2X1_LOC_53/Y 0.01fF
C17203 OR2X1_LOC_160/B OR2X1_LOC_713/A 0.01fF
C17204 OR2X1_LOC_539/Y OR2X1_LOC_174/Y 0.02fF
C17205 AND2X1_LOC_342/a_8_24# OR2X1_LOC_437/A 0.02fF
C17206 AND2X1_LOC_840/B OR2X1_LOC_13/B 0.08fF
C17207 VDD OR2X1_LOC_160/Y 0.12fF
C17208 OR2X1_LOC_505/a_8_216# OR2X1_LOC_56/A 0.00fF
C17209 OR2X1_LOC_533/Y OR2X1_LOC_51/Y 0.01fF
C17210 D_INPUT_2 AND2X1_LOC_14/a_8_24# 0.02fF
C17211 OR2X1_LOC_634/A AND2X1_LOC_7/B 0.03fF
C17212 OR2X1_LOC_66/A OR2X1_LOC_549/A 0.12fF
C17213 OR2X1_LOC_51/Y AND2X1_LOC_212/Y 0.02fF
C17214 OR2X1_LOC_123/a_8_216# AND2X1_LOC_65/A 0.01fF
C17215 OR2X1_LOC_133/a_8_216# OR2X1_LOC_56/A 0.02fF
C17216 OR2X1_LOC_6/B OR2X1_LOC_612/a_8_216# 0.03fF
C17217 INPUT_0 OR2X1_LOC_633/A 0.58fF
C17218 OR2X1_LOC_6/B OR2X1_LOC_600/A 9.11fF
C17219 AND2X1_LOC_367/A AND2X1_LOC_786/Y 0.10fF
C17220 AND2X1_LOC_22/Y OR2X1_LOC_474/Y 0.10fF
C17221 OR2X1_LOC_40/Y AND2X1_LOC_507/a_8_24# 0.01fF
C17222 AND2X1_LOC_566/B OR2X1_LOC_426/B 0.04fF
C17223 OR2X1_LOC_99/Y OR2X1_LOC_771/B 0.05fF
C17224 AND2X1_LOC_444/a_8_24# AND2X1_LOC_212/Y 0.03fF
C17225 VDD OR2X1_LOC_93/Y 0.12fF
C17226 AND2X1_LOC_114/Y AND2X1_LOC_116/a_8_24# 0.19fF
C17227 OR2X1_LOC_485/A AND2X1_LOC_247/a_8_24# 0.01fF
C17228 AND2X1_LOC_663/A AND2X1_LOC_476/Y 0.10fF
C17229 AND2X1_LOC_51/Y OR2X1_LOC_705/a_8_216# 0.01fF
C17230 OR2X1_LOC_369/Y OR2X1_LOC_40/Y 0.00fF
C17231 AND2X1_LOC_573/A AND2X1_LOC_772/Y 0.02fF
C17232 AND2X1_LOC_182/A OR2X1_LOC_91/A 0.19fF
C17233 AND2X1_LOC_857/Y OR2X1_LOC_12/Y 0.04fF
C17234 AND2X1_LOC_732/a_8_24# AND2X1_LOC_732/B 0.00fF
C17235 VDD AND2X1_LOC_447/Y 0.19fF
C17236 AND2X1_LOC_91/B OR2X1_LOC_447/a_8_216# 0.02fF
C17237 AND2X1_LOC_30/a_36_24# INPUT_6 0.00fF
C17238 VDD AND2X1_LOC_334/Y 0.01fF
C17239 AND2X1_LOC_22/Y AND2X1_LOC_328/a_36_24# 0.00fF
C17240 OR2X1_LOC_643/a_36_216# OR2X1_LOC_539/B 0.03fF
C17241 OR2X1_LOC_831/A OR2X1_LOC_804/a_8_216# 0.01fF
C17242 OR2X1_LOC_326/B AND2X1_LOC_44/Y 0.14fF
C17243 OR2X1_LOC_160/B OR2X1_LOC_803/A 0.01fF
C17244 OR2X1_LOC_124/A OR2X1_LOC_160/B 0.03fF
C17245 AND2X1_LOC_486/Y OR2X1_LOC_373/Y 0.19fF
C17246 AND2X1_LOC_18/Y AND2X1_LOC_92/Y 0.17fF
C17247 OR2X1_LOC_523/Y AND2X1_LOC_44/Y 0.01fF
C17248 OR2X1_LOC_833/Y AND2X1_LOC_40/Y 0.03fF
C17249 AND2X1_LOC_768/a_8_24# AND2X1_LOC_772/B 0.00fF
C17250 OR2X1_LOC_757/A AND2X1_LOC_758/a_8_24# 0.01fF
C17251 AND2X1_LOC_392/A OR2X1_LOC_329/B 10.44fF
C17252 OR2X1_LOC_347/Y OR2X1_LOC_360/a_8_216# 0.39fF
C17253 OR2X1_LOC_179/Y OR2X1_LOC_158/A 0.01fF
C17254 OR2X1_LOC_32/B AND2X1_LOC_202/Y 0.15fF
C17255 AND2X1_LOC_95/Y OR2X1_LOC_721/a_36_216# 0.00fF
C17256 OR2X1_LOC_175/Y OR2X1_LOC_799/a_8_216# 0.03fF
C17257 AND2X1_LOC_721/Y AND2X1_LOC_807/Y 0.02fF
C17258 OR2X1_LOC_45/B AND2X1_LOC_621/Y 0.03fF
C17259 OR2X1_LOC_817/Y AND2X1_LOC_789/Y 0.02fF
C17260 OR2X1_LOC_516/A AND2X1_LOC_804/A 0.01fF
C17261 OR2X1_LOC_113/Y OR2X1_LOC_66/A 0.01fF
C17262 OR2X1_LOC_135/Y OR2X1_LOC_48/B 0.36fF
C17263 OR2X1_LOC_316/Y OR2X1_LOC_428/A 0.02fF
C17264 OR2X1_LOC_114/B AND2X1_LOC_71/a_36_24# 0.00fF
C17265 AND2X1_LOC_714/B AND2X1_LOC_841/B 0.07fF
C17266 OR2X1_LOC_188/Y OR2X1_LOC_203/Y 0.00fF
C17267 OR2X1_LOC_49/A OR2X1_LOC_87/a_8_216# 0.02fF
C17268 OR2X1_LOC_168/B OR2X1_LOC_78/A 0.02fF
C17269 OR2X1_LOC_186/Y AND2X1_LOC_43/B 0.02fF
C17270 OR2X1_LOC_354/A OR2X1_LOC_66/A 0.07fF
C17271 AND2X1_LOC_40/Y AND2X1_LOC_387/a_8_24# 0.17fF
C17272 OR2X1_LOC_87/A OR2X1_LOC_357/B 0.01fF
C17273 AND2X1_LOC_64/Y AND2X1_LOC_3/Y 0.26fF
C17274 VDD OR2X1_LOC_330/Y 0.16fF
C17275 OR2X1_LOC_292/Y OR2X1_LOC_56/A 0.00fF
C17276 VDD OR2X1_LOC_220/A 0.26fF
C17277 OR2X1_LOC_589/A OR2X1_LOC_433/Y 0.03fF
C17278 AND2X1_LOC_354/B OR2X1_LOC_428/A 0.03fF
C17279 OR2X1_LOC_595/Y AND2X1_LOC_643/a_8_24# 0.07fF
C17280 OR2X1_LOC_175/Y OR2X1_LOC_219/B 0.01fF
C17281 AND2X1_LOC_47/Y OR2X1_LOC_501/a_8_216# 0.01fF
C17282 OR2X1_LOC_680/A AND2X1_LOC_212/Y 0.07fF
C17283 AND2X1_LOC_535/Y AND2X1_LOC_801/a_8_24# 0.00fF
C17284 OR2X1_LOC_589/A AND2X1_LOC_138/a_8_24# 0.17fF
C17285 OR2X1_LOC_47/Y OR2X1_LOC_80/A 0.40fF
C17286 OR2X1_LOC_244/A OR2X1_LOC_141/a_8_216# 0.03fF
C17287 OR2X1_LOC_532/B OR2X1_LOC_777/B 0.05fF
C17288 OR2X1_LOC_467/A OR2X1_LOC_478/a_8_216# 0.01fF
C17289 AND2X1_LOC_70/Y AND2X1_LOC_173/a_8_24# 0.00fF
C17290 OR2X1_LOC_49/A OR2X1_LOC_43/A 0.91fF
C17291 VDD AND2X1_LOC_649/B 0.23fF
C17292 OR2X1_LOC_31/Y OR2X1_LOC_13/B 0.20fF
C17293 AND2X1_LOC_41/A OR2X1_LOC_274/a_8_216# 0.01fF
C17294 OR2X1_LOC_744/A AND2X1_LOC_266/a_8_24# 0.01fF
C17295 AND2X1_LOC_599/a_8_24# AND2X1_LOC_3/Y 0.01fF
C17296 OR2X1_LOC_160/B OR2X1_LOC_249/a_8_216# 0.07fF
C17297 OR2X1_LOC_485/a_8_216# OR2X1_LOC_59/Y 0.01fF
C17298 VDD AND2X1_LOC_504/a_8_24# -0.00fF
C17299 OR2X1_LOC_474/Y OR2X1_LOC_244/B 0.05fF
C17300 VDD OR2X1_LOC_109/Y 0.62fF
C17301 OR2X1_LOC_312/Y AND2X1_LOC_464/A 0.01fF
C17302 AND2X1_LOC_350/B AND2X1_LOC_211/B 0.89fF
C17303 OR2X1_LOC_852/a_8_216# OR2X1_LOC_472/A 0.03fF
C17304 AND2X1_LOC_562/B OR2X1_LOC_698/Y 0.01fF
C17305 OR2X1_LOC_43/A OR2X1_LOC_381/a_36_216# 0.00fF
C17306 OR2X1_LOC_756/B OR2X1_LOC_502/A 0.03fF
C17307 OR2X1_LOC_783/A OR2X1_LOC_712/B 0.00fF
C17308 VDD OR2X1_LOC_570/a_8_216# 0.00fF
C17309 AND2X1_LOC_733/a_8_24# OR2X1_LOC_164/Y 0.10fF
C17310 AND2X1_LOC_215/Y OR2X1_LOC_316/Y 0.55fF
C17311 AND2X1_LOC_390/B OR2X1_LOC_428/A 0.07fF
C17312 OR2X1_LOC_74/A AND2X1_LOC_786/Y 0.09fF
C17313 OR2X1_LOC_316/a_8_216# OR2X1_LOC_22/Y 0.05fF
C17314 AND2X1_LOC_764/a_8_24# OR2X1_LOC_160/A 0.02fF
C17315 OR2X1_LOC_74/A OR2X1_LOC_323/a_8_216# 0.03fF
C17316 AND2X1_LOC_82/Y AND2X1_LOC_3/Y 0.00fF
C17317 OR2X1_LOC_190/A OR2X1_LOC_375/A 0.07fF
C17318 OR2X1_LOC_45/B AND2X1_LOC_650/a_8_24# 0.07fF
C17319 OR2X1_LOC_335/a_36_216# OR2X1_LOC_121/B 0.00fF
C17320 OR2X1_LOC_814/A OR2X1_LOC_363/a_8_216# 0.01fF
C17321 AND2X1_LOC_721/Y OR2X1_LOC_488/Y 0.11fF
C17322 OR2X1_LOC_45/a_8_216# OR2X1_LOC_59/Y 0.02fF
C17323 OR2X1_LOC_701/Y OR2X1_LOC_59/Y 0.01fF
C17324 OR2X1_LOC_51/Y OR2X1_LOC_265/Y 0.03fF
C17325 AND2X1_LOC_784/Y OR2X1_LOC_52/B 0.17fF
C17326 OR2X1_LOC_446/B OR2X1_LOC_512/a_8_216# 0.03fF
C17327 OR2X1_LOC_739/B D_GATE_741 0.01fF
C17328 AND2X1_LOC_59/Y OR2X1_LOC_78/A 0.25fF
C17329 OR2X1_LOC_804/A OR2X1_LOC_303/B 0.18fF
C17330 OR2X1_LOC_669/a_8_216# AND2X1_LOC_860/A 0.03fF
C17331 AND2X1_LOC_91/B OR2X1_LOC_62/B 0.03fF
C17332 OR2X1_LOC_756/B OR2X1_LOC_571/B 0.02fF
C17333 AND2X1_LOC_571/A OR2X1_LOC_71/Y 0.00fF
C17334 OR2X1_LOC_612/Y OR2X1_LOC_39/A 0.01fF
C17335 OR2X1_LOC_604/A OR2X1_LOC_626/a_8_216# 0.05fF
C17336 OR2X1_LOC_431/Y OR2X1_LOC_428/A 0.02fF
C17337 VDD OR2X1_LOC_847/B 0.00fF
C17338 AND2X1_LOC_566/B OR2X1_LOC_743/A 0.03fF
C17339 OR2X1_LOC_116/A OR2X1_LOC_244/B 0.31fF
C17340 AND2X1_LOC_866/B AND2X1_LOC_805/Y 0.02fF
C17341 OR2X1_LOC_710/B OR2X1_LOC_269/B 0.24fF
C17342 AND2X1_LOC_702/Y OR2X1_LOC_56/A 0.03fF
C17343 OR2X1_LOC_468/A OR2X1_LOC_778/Y 0.47fF
C17344 OR2X1_LOC_532/B OR2X1_LOC_831/B 0.03fF
C17345 OR2X1_LOC_111/a_8_216# OR2X1_LOC_31/Y 0.02fF
C17346 AND2X1_LOC_307/Y OR2X1_LOC_16/A 0.14fF
C17347 OR2X1_LOC_628/Y OR2X1_LOC_816/A 0.04fF
C17348 OR2X1_LOC_59/Y OR2X1_LOC_44/Y 2.89fF
C17349 OR2X1_LOC_733/a_8_216# OR2X1_LOC_737/A 0.01fF
C17350 OR2X1_LOC_733/B OR2X1_LOC_733/A 0.08fF
C17351 AND2X1_LOC_191/B OR2X1_LOC_26/Y 0.03fF
C17352 OR2X1_LOC_802/a_8_216# OR2X1_LOC_624/A 0.01fF
C17353 AND2X1_LOC_211/B AND2X1_LOC_326/B 0.07fF
C17354 OR2X1_LOC_529/Y OR2X1_LOC_600/A 0.00fF
C17355 AND2X1_LOC_243/a_8_24# AND2X1_LOC_243/Y 0.00fF
C17356 OR2X1_LOC_400/A OR2X1_LOC_756/B 0.01fF
C17357 OR2X1_LOC_26/Y AND2X1_LOC_469/B 0.03fF
C17358 OR2X1_LOC_40/Y AND2X1_LOC_651/B 0.01fF
C17359 AND2X1_LOC_276/a_8_24# OR2X1_LOC_39/A 0.03fF
C17360 AND2X1_LOC_190/a_8_24# AND2X1_LOC_717/B 0.03fF
C17361 VDD OR2X1_LOC_557/A 0.53fF
C17362 AND2X1_LOC_434/Y OR2X1_LOC_52/B 0.07fF
C17363 AND2X1_LOC_784/A AND2X1_LOC_364/Y 0.00fF
C17364 AND2X1_LOC_50/Y OR2X1_LOC_375/A 0.04fF
C17365 OR2X1_LOC_369/Y OR2X1_LOC_7/A 0.03fF
C17366 AND2X1_LOC_191/B OR2X1_LOC_89/A 0.06fF
C17367 OR2X1_LOC_168/B OR2X1_LOC_155/A 0.03fF
C17368 OR2X1_LOC_89/A AND2X1_LOC_469/B 0.03fF
C17369 AND2X1_LOC_674/a_8_24# OR2X1_LOC_733/A 0.24fF
C17370 VDD AND2X1_LOC_117/a_8_24# 0.00fF
C17371 OR2X1_LOC_643/A OR2X1_LOC_659/A 0.01fF
C17372 AND2X1_LOC_733/Y OR2X1_LOC_26/Y 0.07fF
C17373 OR2X1_LOC_623/a_8_216# OR2X1_LOC_624/A 0.02fF
C17374 AND2X1_LOC_721/Y OR2X1_LOC_95/Y 0.07fF
C17375 AND2X1_LOC_840/A OR2X1_LOC_39/A 0.02fF
C17376 AND2X1_LOC_857/Y AND2X1_LOC_650/Y 0.00fF
C17377 AND2X1_LOC_259/Y OR2X1_LOC_297/A 0.02fF
C17378 OR2X1_LOC_585/A OR2X1_LOC_234/Y 0.35fF
C17379 INPUT_0 OR2X1_LOC_827/Y 0.01fF
C17380 AND2X1_LOC_863/Y OR2X1_LOC_428/A 0.07fF
C17381 AND2X1_LOC_711/Y AND2X1_LOC_501/a_8_24# 0.05fF
C17382 OR2X1_LOC_74/A AND2X1_LOC_218/Y 0.02fF
C17383 VDD AND2X1_LOC_729/B 0.76fF
C17384 AND2X1_LOC_47/Y AND2X1_LOC_44/Y 0.31fF
C17385 AND2X1_LOC_175/B OR2X1_LOC_18/Y 0.16fF
C17386 AND2X1_LOC_116/Y OR2X1_LOC_59/Y 1.06fF
C17387 AND2X1_LOC_566/B OR2X1_LOC_246/A 0.01fF
C17388 OR2X1_LOC_109/Y OR2X1_LOC_315/Y 0.01fF
C17389 OR2X1_LOC_532/B OR2X1_LOC_344/A 0.03fF
C17390 AND2X1_LOC_357/a_8_24# OR2X1_LOC_6/A 0.01fF
C17391 OR2X1_LOC_289/Y OR2X1_LOC_171/Y 0.29fF
C17392 OR2X1_LOC_184/Y OR2X1_LOC_184/a_8_216# 0.00fF
C17393 AND2X1_LOC_733/Y OR2X1_LOC_89/A 0.42fF
C17394 OR2X1_LOC_351/B OR2X1_LOC_814/A 0.35fF
C17395 AND2X1_LOC_576/Y OR2X1_LOC_427/A 0.07fF
C17396 OR2X1_LOC_799/A OR2X1_LOC_130/A 0.02fF
C17397 OR2X1_LOC_237/a_8_216# OR2X1_LOC_39/A 0.04fF
C17398 AND2X1_LOC_141/A OR2X1_LOC_7/A 0.04fF
C17399 AND2X1_LOC_160/a_36_24# OR2X1_LOC_7/A 0.00fF
C17400 OR2X1_LOC_656/Y AND2X1_LOC_3/Y 0.09fF
C17401 OR2X1_LOC_643/a_8_216# OR2X1_LOC_475/B 0.47fF
C17402 OR2X1_LOC_6/B OR2X1_LOC_720/B -0.02fF
C17403 OR2X1_LOC_118/Y AND2X1_LOC_266/Y 0.81fF
C17404 AND2X1_LOC_40/Y OR2X1_LOC_574/A 0.03fF
C17405 OR2X1_LOC_160/B OR2X1_LOC_750/a_8_216# 0.01fF
C17406 AND2X1_LOC_583/a_36_24# OR2X1_LOC_636/B 0.00fF
C17407 OR2X1_LOC_640/a_8_216# OR2X1_LOC_462/B 0.01fF
C17408 AND2X1_LOC_845/Y AND2X1_LOC_243/Y 1.38fF
C17409 AND2X1_LOC_135/a_36_24# OR2X1_LOC_78/B 0.01fF
C17410 OR2X1_LOC_703/B AND2X1_LOC_166/a_36_24# 0.00fF
C17411 OR2X1_LOC_169/a_8_216# OR2X1_LOC_169/B 0.47fF
C17412 OR2X1_LOC_482/Y OR2X1_LOC_95/Y 0.00fF
C17413 AND2X1_LOC_570/Y AND2X1_LOC_574/A 0.00fF
C17414 OR2X1_LOC_460/Y OR2X1_LOC_463/B 0.07fF
C17415 OR2X1_LOC_169/B OR2X1_LOC_468/Y 0.01fF
C17416 OR2X1_LOC_87/B OR2X1_LOC_87/a_8_216# 0.00fF
C17417 AND2X1_LOC_365/A AND2X1_LOC_661/A 0.18fF
C17418 OR2X1_LOC_22/Y AND2X1_LOC_637/a_8_24# 0.00fF
C17419 AND2X1_LOC_710/a_8_24# OR2X1_LOC_748/A 0.01fF
C17420 AND2X1_LOC_12/Y OR2X1_LOC_68/a_8_216# 0.01fF
C17421 OR2X1_LOC_481/A OR2X1_LOC_92/Y 0.03fF
C17422 OR2X1_LOC_235/B OR2X1_LOC_293/a_36_216# 0.00fF
C17423 AND2X1_LOC_741/a_36_24# AND2X1_LOC_711/Y 0.01fF
C17424 OR2X1_LOC_201/A OR2X1_LOC_206/A 0.34fF
C17425 AND2X1_LOC_59/Y OR2X1_LOC_155/A 0.09fF
C17426 AND2X1_LOC_97/a_36_24# OR2X1_LOC_89/A 0.00fF
C17427 AND2X1_LOC_99/Y AND2X1_LOC_663/B 0.42fF
C17428 AND2X1_LOC_382/a_8_24# OR2X1_LOC_391/B 0.01fF
C17429 OR2X1_LOC_756/B AND2X1_LOC_48/A 0.07fF
C17430 OR2X1_LOC_433/a_8_216# OR2X1_LOC_44/Y 0.01fF
C17431 INPUT_3 AND2X1_LOC_37/a_8_24# 0.14fF
C17432 OR2X1_LOC_13/B OR2X1_LOC_320/a_8_216# 0.03fF
C17433 AND2X1_LOC_44/Y OR2X1_LOC_598/A 0.08fF
C17434 OR2X1_LOC_364/A OR2X1_LOC_269/B 0.07fF
C17435 OR2X1_LOC_161/B OR2X1_LOC_374/Y 0.19fF
C17436 OR2X1_LOC_262/Y AND2X1_LOC_266/Y 0.06fF
C17437 OR2X1_LOC_185/Y OR2X1_LOC_269/B 3.79fF
C17438 AND2X1_LOC_624/A OR2X1_LOC_239/Y 0.03fF
C17439 OR2X1_LOC_264/Y OR2X1_LOC_121/B 1.38fF
C17440 OR2X1_LOC_141/B OR2X1_LOC_510/Y 0.00fF
C17441 OR2X1_LOC_702/A OR2X1_LOC_161/A 0.03fF
C17442 OR2X1_LOC_820/B OR2X1_LOC_44/Y 0.00fF
C17443 OR2X1_LOC_45/Y OR2X1_LOC_304/Y 0.31fF
C17444 OR2X1_LOC_193/A AND2X1_LOC_16/a_8_24# 0.37fF
C17445 AND2X1_LOC_342/a_8_24# OR2X1_LOC_753/A 0.01fF
C17446 OR2X1_LOC_18/Y OR2X1_LOC_617/Y 0.04fF
C17447 OR2X1_LOC_481/A OR2X1_LOC_257/a_8_216# 0.01fF
C17448 OR2X1_LOC_140/A OR2X1_LOC_786/Y 0.01fF
C17449 OR2X1_LOC_70/Y OR2X1_LOC_45/a_8_216# 0.01fF
C17450 D_INPUT_0 AND2X1_LOC_240/a_8_24# 0.05fF
C17451 OR2X1_LOC_829/a_8_216# AND2X1_LOC_729/B 0.01fF
C17452 AND2X1_LOC_382/a_36_24# OR2X1_LOC_269/B 0.00fF
C17453 OR2X1_LOC_3/Y OR2X1_LOC_67/a_8_216# 0.01fF
C17454 D_INPUT_7 AND2X1_LOC_25/Y 0.01fF
C17455 AND2X1_LOC_856/B OR2X1_LOC_48/B 0.00fF
C17456 OR2X1_LOC_377/A OR2X1_LOC_193/A 0.01fF
C17457 INPUT_0 AND2X1_LOC_826/a_36_24# 0.01fF
C17458 AND2X1_LOC_181/a_8_24# AND2X1_LOC_866/A 0.06fF
C17459 AND2X1_LOC_863/A OR2X1_LOC_48/B 0.06fF
C17460 AND2X1_LOC_749/a_8_24# OR2X1_LOC_655/B 0.23fF
C17461 OR2X1_LOC_222/a_36_216# AND2X1_LOC_92/Y 0.01fF
C17462 AND2X1_LOC_259/Y OR2X1_LOC_43/A 0.00fF
C17463 OR2X1_LOC_305/a_8_216# OR2X1_LOC_3/Y 0.02fF
C17464 AND2X1_LOC_512/Y AND2X1_LOC_169/a_8_24# 0.02fF
C17465 AND2X1_LOC_664/a_8_24# AND2X1_LOC_805/Y 0.19fF
C17466 OR2X1_LOC_18/Y AND2X1_LOC_464/Y 0.03fF
C17467 AND2X1_LOC_58/a_8_24# D_INPUT_0 0.04fF
C17468 AND2X1_LOC_789/a_36_24# INPUT_1 0.00fF
C17469 AND2X1_LOC_360/a_8_24# OR2X1_LOC_417/A 0.02fF
C17470 OR2X1_LOC_92/Y OR2X1_LOC_71/Y 0.76fF
C17471 AND2X1_LOC_711/Y OR2X1_LOC_44/Y 0.01fF
C17472 AND2X1_LOC_753/B AND2X1_LOC_7/Y 0.10fF
C17473 OR2X1_LOC_60/a_36_216# OR2X1_LOC_39/A 0.02fF
C17474 AND2X1_LOC_56/B OR2X1_LOC_35/B 0.23fF
C17475 OR2X1_LOC_818/Y D_INPUT_0 0.02fF
C17476 OR2X1_LOC_70/Y OR2X1_LOC_44/Y 0.13fF
C17477 AND2X1_LOC_31/Y OR2X1_LOC_741/a_8_216# 0.01fF
C17478 AND2X1_LOC_580/A AND2X1_LOC_663/B 0.00fF
C17479 OR2X1_LOC_87/A OR2X1_LOC_202/a_8_216# 0.03fF
C17480 OR2X1_LOC_660/B AND2X1_LOC_48/A 0.01fF
C17481 OR2X1_LOC_196/B AND2X1_LOC_43/B 0.15fF
C17482 OR2X1_LOC_319/a_8_216# D_INPUT_0 0.02fF
C17483 AND2X1_LOC_658/A AND2X1_LOC_793/Y 0.07fF
C17484 OR2X1_LOC_287/B OR2X1_LOC_850/A 0.01fF
C17485 AND2X1_LOC_348/A AND2X1_LOC_866/A 0.03fF
C17486 OR2X1_LOC_185/A OR2X1_LOC_243/a_8_216# 0.02fF
C17487 OR2X1_LOC_493/A OR2X1_LOC_532/B 0.18fF
C17488 AND2X1_LOC_12/Y OR2X1_LOC_814/A 1.72fF
C17489 OR2X1_LOC_127/a_8_216# OR2X1_LOC_225/a_8_216# 0.47fF
C17490 OR2X1_LOC_95/Y OR2X1_LOC_586/Y 0.09fF
C17491 OR2X1_LOC_51/Y OR2X1_LOC_163/A 0.05fF
C17492 AND2X1_LOC_692/a_8_24# AND2X1_LOC_43/B 0.04fF
C17493 AND2X1_LOC_158/a_8_24# AND2X1_LOC_51/Y 0.17fF
C17494 OR2X1_LOC_377/A D_INPUT_0 0.39fF
C17495 AND2X1_LOC_514/Y OR2X1_LOC_44/Y 0.07fF
C17496 OR2X1_LOC_643/A OR2X1_LOC_121/B 0.03fF
C17497 OR2X1_LOC_757/A AND2X1_LOC_805/a_8_24# 0.01fF
C17498 OR2X1_LOC_44/a_8_216# OR2X1_LOC_47/a_8_216# 0.47fF
C17499 AND2X1_LOC_578/A OR2X1_LOC_74/A 0.12fF
C17500 AND2X1_LOC_633/Y OR2X1_LOC_85/A 0.04fF
C17501 OR2X1_LOC_40/Y AND2X1_LOC_793/B 0.00fF
C17502 OR2X1_LOC_71/Y OR2X1_LOC_65/B 0.08fF
C17503 OR2X1_LOC_121/B OR2X1_LOC_778/Y 0.05fF
C17504 D_INPUT_0 AND2X1_LOC_824/B 0.00fF
C17505 OR2X1_LOC_12/Y OR2X1_LOC_437/A 0.11fF
C17506 OR2X1_LOC_294/Y OR2X1_LOC_366/Y 0.03fF
C17507 OR2X1_LOC_420/a_8_216# OR2X1_LOC_64/Y 0.02fF
C17508 D_INPUT_7 AND2X1_LOC_51/Y 0.09fF
C17509 AND2X1_LOC_76/Y AND2X1_LOC_851/B 0.14fF
C17510 AND2X1_LOC_22/Y OR2X1_LOC_771/B 0.01fF
C17511 OR2X1_LOC_17/Y AND2X1_LOC_639/a_36_24# 0.00fF
C17512 AND2X1_LOC_733/Y AND2X1_LOC_804/a_8_24# 0.03fF
C17513 OR2X1_LOC_576/A OR2X1_LOC_217/A 0.01fF
C17514 D_INPUT_0 OR2X1_LOC_85/A 0.22fF
C17515 AND2X1_LOC_566/Y OR2X1_LOC_417/Y 0.01fF
C17516 D_INPUT_0 OR2X1_LOC_203/Y 0.04fF
C17517 OR2X1_LOC_3/Y OR2X1_LOC_665/a_8_216# 0.01fF
C17518 AND2X1_LOC_40/Y AND2X1_LOC_761/a_8_24# 0.17fF
C17519 AND2X1_LOC_22/Y OR2X1_LOC_776/A 0.00fF
C17520 OR2X1_LOC_84/B AND2X1_LOC_133/a_36_24# 0.00fF
C17521 OR2X1_LOC_609/a_8_216# OR2X1_LOC_46/A 0.01fF
C17522 OR2X1_LOC_3/Y AND2X1_LOC_537/Y 0.07fF
C17523 OR2X1_LOC_65/B D_INPUT_1 0.01fF
C17524 OR2X1_LOC_698/a_8_216# AND2X1_LOC_793/B 0.02fF
C17525 AND2X1_LOC_776/Y AND2X1_LOC_564/B 0.18fF
C17526 OR2X1_LOC_3/Y AND2X1_LOC_66/a_8_24# 0.01fF
C17527 OR2X1_LOC_485/A OR2X1_LOC_226/a_8_216# 0.01fF
C17528 OR2X1_LOC_22/Y AND2X1_LOC_660/Y 0.01fF
C17529 AND2X1_LOC_76/Y OR2X1_LOC_595/Y 0.01fF
C17530 OR2X1_LOC_243/a_36_216# AND2X1_LOC_42/B 0.00fF
C17531 OR2X1_LOC_375/A OR2X1_LOC_214/B 0.01fF
C17532 OR2X1_LOC_47/Y OR2X1_LOC_6/A 0.11fF
C17533 AND2X1_LOC_728/a_8_24# OR2X1_LOC_679/A 0.09fF
C17534 AND2X1_LOC_324/a_36_24# OR2X1_LOC_46/A 0.01fF
C17535 AND2X1_LOC_339/a_36_24# OR2X1_LOC_31/Y 0.01fF
C17536 OR2X1_LOC_375/A OR2X1_LOC_241/B 0.06fF
C17537 OR2X1_LOC_184/Y OR2X1_LOC_44/Y 0.03fF
C17538 OR2X1_LOC_293/a_8_216# OR2X1_LOC_54/Y 0.01fF
C17539 AND2X1_LOC_358/a_8_24# OR2X1_LOC_46/A 0.01fF
C17540 OR2X1_LOC_146/a_36_216# AND2X1_LOC_213/B 0.00fF
C17541 AND2X1_LOC_841/a_8_24# OR2X1_LOC_74/A -0.01fF
C17542 AND2X1_LOC_23/a_8_24# OR2X1_LOC_750/A 0.08fF
C17543 AND2X1_LOC_191/Y AND2X1_LOC_866/a_8_24# 0.20fF
C17544 OR2X1_LOC_146/Y OR2X1_LOC_89/A 0.08fF
C17545 AND2X1_LOC_326/a_8_24# OR2X1_LOC_46/A 0.06fF
C17546 OR2X1_LOC_91/Y OR2X1_LOC_406/A 0.08fF
C17547 OR2X1_LOC_181/B OR2X1_LOC_742/B 0.14fF
C17548 AND2X1_LOC_345/Y OR2X1_LOC_55/a_36_216# 0.02fF
C17549 OR2X1_LOC_744/A OR2X1_LOC_142/a_8_216# 0.01fF
C17550 OR2X1_LOC_807/A OR2X1_LOC_675/Y 0.16fF
C17551 OR2X1_LOC_392/B OR2X1_LOC_161/B 0.03fF
C17552 AND2X1_LOC_7/B OR2X1_LOC_633/A 0.11fF
C17553 OR2X1_LOC_35/Y AND2X1_LOC_36/Y 0.03fF
C17554 OR2X1_LOC_149/B OR2X1_LOC_149/a_8_216# 0.00fF
C17555 AND2X1_LOC_639/B OR2X1_LOC_428/A 1.33fF
C17556 AND2X1_LOC_34/Y OR2X1_LOC_68/B 0.01fF
C17557 OR2X1_LOC_739/A OR2X1_LOC_151/a_8_216# 0.01fF
C17558 AND2X1_LOC_5/a_8_24# INPUT_1 0.01fF
C17559 OR2X1_LOC_70/A OR2X1_LOC_44/Y 0.09fF
C17560 OR2X1_LOC_595/Y OR2X1_LOC_52/B 0.02fF
C17561 OR2X1_LOC_154/A OR2X1_LOC_228/Y 0.14fF
C17562 OR2X1_LOC_628/Y OR2X1_LOC_95/Y 0.19fF
C17563 OR2X1_LOC_802/Y AND2X1_LOC_31/Y 0.02fF
C17564 AND2X1_LOC_521/a_8_24# AND2X1_LOC_44/Y 0.01fF
C17565 AND2X1_LOC_471/a_8_24# OR2X1_LOC_95/Y 0.06fF
C17566 OR2X1_LOC_97/A OR2X1_LOC_151/A 0.03fF
C17567 OR2X1_LOC_154/A OR2X1_LOC_513/Y 0.01fF
C17568 OR2X1_LOC_160/A OR2X1_LOC_71/A 0.04fF
C17569 OR2X1_LOC_89/A AND2X1_LOC_848/A 0.01fF
C17570 OR2X1_LOC_447/a_8_216# OR2X1_LOC_446/B 0.01fF
C17571 OR2X1_LOC_598/Y OR2X1_LOC_855/A 0.45fF
C17572 OR2X1_LOC_696/A INPUT_0 0.11fF
C17573 VDD AND2X1_LOC_220/B 0.40fF
C17574 AND2X1_LOC_91/B OR2X1_LOC_468/A 0.03fF
C17575 OR2X1_LOC_269/B OR2X1_LOC_568/A 0.46fF
C17576 OR2X1_LOC_52/B AND2X1_LOC_781/a_8_24# 0.02fF
C17577 OR2X1_LOC_45/B OR2X1_LOC_527/a_36_216# 0.00fF
C17578 OR2X1_LOC_309/Y OR2X1_LOC_428/A 0.12fF
C17579 OR2X1_LOC_506/A OR2X1_LOC_728/a_36_216# 0.02fF
C17580 OR2X1_LOC_774/Y OR2X1_LOC_557/a_36_216# 0.00fF
C17581 AND2X1_LOC_64/Y INPUT_0 0.16fF
C17582 OR2X1_LOC_527/Y OR2X1_LOC_406/A 0.01fF
C17583 OR2X1_LOC_74/A OR2X1_LOC_88/a_8_216# 0.05fF
C17584 AND2X1_LOC_56/a_8_24# OR2X1_LOC_651/A 0.02fF
C17585 OR2X1_LOC_235/a_36_216# OR2X1_LOC_71/A 0.00fF
C17586 OR2X1_LOC_62/a_8_216# D_INPUT_1 0.01fF
C17587 OR2X1_LOC_7/A AND2X1_LOC_793/B 0.01fF
C17588 OR2X1_LOC_854/a_8_216# OR2X1_LOC_319/Y 0.06fF
C17589 OR2X1_LOC_450/A OR2X1_LOC_161/B 0.24fF
C17590 AND2X1_LOC_814/a_8_24# AND2X1_LOC_793/Y 0.01fF
C17591 OR2X1_LOC_815/A AND2X1_LOC_792/Y 0.02fF
C17592 OR2X1_LOC_26/Y OR2X1_LOC_164/a_8_216# 0.01fF
C17593 AND2X1_LOC_91/B OR2X1_LOC_571/a_8_216# 0.01fF
C17594 OR2X1_LOC_696/A AND2X1_LOC_717/Y 0.19fF
C17595 OR2X1_LOC_35/A OR2X1_LOC_35/a_8_216# 0.39fF
C17596 OR2X1_LOC_45/B OR2X1_LOC_59/Y 5.59fF
C17597 D_INPUT_3 AND2X1_LOC_672/a_8_24# 0.07fF
C17598 AND2X1_LOC_462/a_8_24# OR2X1_LOC_598/A 0.21fF
C17599 OR2X1_LOC_744/A OR2X1_LOC_428/A 0.12fF
C17600 AND2X1_LOC_140/a_8_24# AND2X1_LOC_217/a_8_24# 0.23fF
C17601 AND2X1_LOC_1/Y AND2X1_LOC_31/Y 0.07fF
C17602 OR2X1_LOC_185/A AND2X1_LOC_238/a_36_24# 0.00fF
C17603 OR2X1_LOC_190/A OR2X1_LOC_549/A 0.07fF
C17604 AND2X1_LOC_86/B OR2X1_LOC_71/A 0.08fF
C17605 OR2X1_LOC_790/A AND2X1_LOC_18/Y 0.00fF
C17606 OR2X1_LOC_62/A OR2X1_LOC_619/a_8_216# 0.09fF
C17607 OR2X1_LOC_720/B OR2X1_LOC_598/A -0.02fF
C17608 OR2X1_LOC_744/A OR2X1_LOC_595/A 0.08fF
C17609 OR2X1_LOC_656/a_8_216# OR2X1_LOC_68/B 0.18fF
C17610 AND2X1_LOC_40/Y OR2X1_LOC_855/A 0.01fF
C17611 OR2X1_LOC_13/a_8_216# AND2X1_LOC_434/Y 0.03fF
C17612 OR2X1_LOC_756/B OR2X1_LOC_34/a_8_216# 0.01fF
C17613 OR2X1_LOC_851/B OR2X1_LOC_858/A 0.03fF
C17614 OR2X1_LOC_756/B OR2X1_LOC_489/A 0.01fF
C17615 AND2X1_LOC_22/Y OR2X1_LOC_637/B 0.00fF
C17616 OR2X1_LOC_208/A OR2X1_LOC_377/A 0.02fF
C17617 AND2X1_LOC_541/Y AND2X1_LOC_772/B 0.01fF
C17618 OR2X1_LOC_345/Y OR2X1_LOC_756/B 0.34fF
C17619 OR2X1_LOC_61/Y OR2X1_LOC_392/B 0.10fF
C17620 OR2X1_LOC_696/A OR2X1_LOC_11/Y 0.05fF
C17621 AND2X1_LOC_91/B OR2X1_LOC_724/a_36_216# 0.00fF
C17622 AND2X1_LOC_64/Y OR2X1_LOC_732/B 0.01fF
C17623 OR2X1_LOC_316/a_8_216# OR2X1_LOC_39/A 0.01fF
C17624 OR2X1_LOC_604/A AND2X1_LOC_436/Y 0.08fF
C17625 AND2X1_LOC_739/B AND2X1_LOC_740/B 0.05fF
C17626 INPUT_5 OR2X1_LOC_375/Y 0.09fF
C17627 AND2X1_LOC_91/a_8_24# OR2X1_LOC_794/A 0.23fF
C17628 OR2X1_LOC_97/A OR2X1_LOC_788/a_8_216# 0.01fF
C17629 AND2X1_LOC_91/B AND2X1_LOC_487/a_8_24# 0.02fF
C17630 AND2X1_LOC_539/Y AND2X1_LOC_593/Y 0.09fF
C17631 OR2X1_LOC_6/B AND2X1_LOC_628/a_8_24# 0.03fF
C17632 AND2X1_LOC_22/Y AND2X1_LOC_11/Y 0.01fF
C17633 OR2X1_LOC_818/a_8_216# OR2X1_LOC_68/B 0.01fF
C17634 OR2X1_LOC_591/Y AND2X1_LOC_718/a_8_24# 0.00fF
C17635 OR2X1_LOC_427/A AND2X1_LOC_244/A 0.03fF
C17636 AND2X1_LOC_86/a_8_24# INPUT_0 0.03fF
C17637 OR2X1_LOC_696/A AND2X1_LOC_560/B 0.12fF
C17638 OR2X1_LOC_360/a_8_216# OR2X1_LOC_66/A 0.01fF
C17639 AND2X1_LOC_703/Y AND2X1_LOC_841/B 0.15fF
C17640 AND2X1_LOC_482/a_36_24# AND2X1_LOC_7/B 0.00fF
C17641 OR2X1_LOC_160/B OR2X1_LOC_778/B 0.03fF
C17642 OR2X1_LOC_686/B OR2X1_LOC_78/B 0.20fF
C17643 AND2X1_LOC_170/B OR2X1_LOC_331/Y 0.01fF
C17644 OR2X1_LOC_768/A VDD -0.00fF
C17645 OR2X1_LOC_114/B OR2X1_LOC_501/B 0.00fF
C17646 AND2X1_LOC_330/a_8_24# OR2X1_LOC_331/A 0.02fF
C17647 AND2X1_LOC_705/a_8_24# OR2X1_LOC_59/Y 0.01fF
C17648 OR2X1_LOC_641/Y OR2X1_LOC_520/a_8_216# 0.06fF
C17649 OR2X1_LOC_756/B OR2X1_LOC_772/A 0.02fF
C17650 OR2X1_LOC_427/A OR2X1_LOC_16/A 0.12fF
C17651 OR2X1_LOC_97/A OR2X1_LOC_405/a_36_216# 0.00fF
C17652 OR2X1_LOC_188/Y OR2X1_LOC_375/A 0.09fF
C17653 AND2X1_LOC_655/A OR2X1_LOC_321/a_36_216# 0.14fF
C17654 OR2X1_LOC_848/A OR2X1_LOC_773/Y 0.03fF
C17655 OR2X1_LOC_468/a_8_216# OR2X1_LOC_567/a_8_216# 0.47fF
C17656 AND2X1_LOC_722/a_8_24# AND2X1_LOC_722/A 0.00fF
C17657 OR2X1_LOC_151/A OR2X1_LOC_475/B 0.03fF
C17658 AND2X1_LOC_227/Y AND2X1_LOC_657/A 0.01fF
C17659 OR2X1_LOC_319/a_36_216# OR2X1_LOC_161/B 0.00fF
C17660 INPUT_0 AND2X1_LOC_33/a_8_24# 0.05fF
C17661 OR2X1_LOC_679/B AND2X1_LOC_213/B 0.01fF
C17662 OR2X1_LOC_241/a_36_216# OR2X1_LOC_121/A 0.00fF
C17663 OR2X1_LOC_122/a_8_216# OR2X1_LOC_122/A 0.47fF
C17664 OR2X1_LOC_866/B OR2X1_LOC_866/a_8_216# 0.06fF
C17665 VDD OR2X1_LOC_39/Y 0.07fF
C17666 AND2X1_LOC_129/a_8_24# AND2X1_LOC_44/Y 0.01fF
C17667 OR2X1_LOC_405/A OR2X1_LOC_390/A 0.02fF
C17668 AND2X1_LOC_91/B OR2X1_LOC_449/B 0.00fF
C17669 OR2X1_LOC_160/A OR2X1_LOC_355/a_8_216# 0.03fF
C17670 OR2X1_LOC_40/Y AND2X1_LOC_348/A 0.03fF
C17671 OR2X1_LOC_377/A OR2X1_LOC_673/B 0.03fF
C17672 OR2X1_LOC_269/a_36_216# OR2X1_LOC_344/A 0.00fF
C17673 OR2X1_LOC_722/a_8_216# OR2X1_LOC_722/B 0.18fF
C17674 OR2X1_LOC_473/A OR2X1_LOC_560/A 0.23fF
C17675 AND2X1_LOC_449/Y OR2X1_LOC_603/Y 0.00fF
C17676 OR2X1_LOC_114/B OR2X1_LOC_147/B 0.14fF
C17677 OR2X1_LOC_685/A OR2X1_LOC_161/B 0.03fF
C17678 AND2X1_LOC_181/a_36_24# OR2X1_LOC_744/A 0.01fF
C17679 OR2X1_LOC_158/A AND2X1_LOC_621/Y 0.02fF
C17680 OR2X1_LOC_108/Y OR2X1_LOC_427/A 0.07fF
C17681 OR2X1_LOC_426/B OR2X1_LOC_92/Y 1.38fF
C17682 OR2X1_LOC_205/Y AND2X1_LOC_31/Y 0.06fF
C17683 AND2X1_LOC_773/Y AND2X1_LOC_784/A 0.10fF
C17684 AND2X1_LOC_216/Y OR2X1_LOC_18/Y 0.02fF
C17685 AND2X1_LOC_348/Y OR2X1_LOC_12/Y 0.09fF
C17686 AND2X1_LOC_41/A AND2X1_LOC_693/a_8_24# 0.01fF
C17687 OR2X1_LOC_770/Y OR2X1_LOC_68/B 0.01fF
C17688 OR2X1_LOC_696/A OR2X1_LOC_64/Y 0.41fF
C17689 VDD OR2X1_LOC_814/Y 0.16fF
C17690 OR2X1_LOC_49/A AND2X1_LOC_818/a_36_24# 0.00fF
C17691 OR2X1_LOC_709/a_36_216# OR2X1_LOC_154/A 0.01fF
C17692 OR2X1_LOC_158/A AND2X1_LOC_668/a_8_24# 0.14fF
C17693 OR2X1_LOC_78/A OR2X1_LOC_623/B 0.01fF
C17694 GATE_811 AND2X1_LOC_738/Y 0.01fF
C17695 OR2X1_LOC_753/A OR2X1_LOC_12/Y 0.04fF
C17696 OR2X1_LOC_151/Y OR2X1_LOC_740/B 0.06fF
C17697 OR2X1_LOC_856/B AND2X1_LOC_110/a_36_24# 0.01fF
C17698 AND2X1_LOC_64/Y OR2X1_LOC_401/A 0.00fF
C17699 OR2X1_LOC_313/a_36_216# OR2X1_LOC_604/A 0.00fF
C17700 OR2X1_LOC_442/Y AND2X1_LOC_804/Y -0.00fF
C17701 AND2X1_LOC_497/a_8_24# OR2X1_LOC_68/B 0.02fF
C17702 OR2X1_LOC_186/Y OR2X1_LOC_810/A 0.00fF
C17703 OR2X1_LOC_799/A OR2X1_LOC_468/A 0.11fF
C17704 AND2X1_LOC_3/Y OR2X1_LOC_342/A 0.09fF
C17705 INPUT_5 OR2X1_LOC_2/a_36_216# 0.00fF
C17706 OR2X1_LOC_20/Y OR2X1_LOC_39/A 0.10fF
C17707 OR2X1_LOC_671/Y OR2X1_LOC_43/A 0.43fF
C17708 AND2X1_LOC_861/B AND2X1_LOC_866/B 0.00fF
C17709 OR2X1_LOC_820/B OR2X1_LOC_382/A 0.02fF
C17710 OR2X1_LOC_604/A OR2X1_LOC_603/a_8_216# 0.01fF
C17711 AND2X1_LOC_719/Y OR2X1_LOC_36/Y 0.08fF
C17712 AND2X1_LOC_508/B AND2X1_LOC_807/Y 0.03fF
C17713 AND2X1_LOC_391/Y OR2X1_LOC_278/Y 0.12fF
C17714 AND2X1_LOC_12/Y OR2X1_LOC_244/Y 0.03fF
C17715 OR2X1_LOC_156/B OR2X1_LOC_479/Y 0.05fF
C17716 OR2X1_LOC_426/B OR2X1_LOC_65/B 0.28fF
C17717 OR2X1_LOC_834/a_36_216# OR2X1_LOC_502/A 0.02fF
C17718 AND2X1_LOC_91/B OR2X1_LOC_121/B 0.06fF
C17719 OR2X1_LOC_91/A OR2X1_LOC_278/Y 0.03fF
C17720 OR2X1_LOC_45/B OR2X1_LOC_70/Y 0.29fF
C17721 AND2X1_LOC_131/a_8_24# OR2X1_LOC_203/Y 0.01fF
C17722 D_INPUT_1 OR2X1_LOC_580/A 0.03fF
C17723 AND2X1_LOC_715/Y OR2X1_LOC_64/Y 0.03fF
C17724 AND2X1_LOC_110/a_8_24# OR2X1_LOC_805/A 0.03fF
C17725 OR2X1_LOC_858/A OR2X1_LOC_160/A 0.10fF
C17726 OR2X1_LOC_91/A AND2X1_LOC_662/B 0.01fF
C17727 AND2X1_LOC_565/B AND2X1_LOC_580/A 0.00fF
C17728 OR2X1_LOC_549/Y D_GATE_366 0.01fF
C17729 D_GATE_479 OR2X1_LOC_470/B 0.75fF
C17730 AND2X1_LOC_861/a_8_24# AND2X1_LOC_807/Y 0.04fF
C17731 OR2X1_LOC_106/Y AND2X1_LOC_116/B 0.03fF
C17732 OR2X1_LOC_512/Y OR2X1_LOC_513/a_8_216# 0.39fF
C17733 OR2X1_LOC_591/Y OR2X1_LOC_89/A 0.01fF
C17734 OR2X1_LOC_198/a_8_216# OR2X1_LOC_532/B 0.01fF
C17735 OR2X1_LOC_470/B OR2X1_LOC_161/B 0.82fF
C17736 OR2X1_LOC_696/A OR2X1_LOC_417/A 0.41fF
C17737 AND2X1_LOC_12/Y OR2X1_LOC_501/B 0.01fF
C17738 OR2X1_LOC_185/A AND2X1_LOC_41/A 0.03fF
C17739 AND2X1_LOC_763/a_8_24# OR2X1_LOC_828/B 0.01fF
C17740 OR2X1_LOC_154/A OR2X1_LOC_702/a_36_216# 0.00fF
C17741 AND2X1_LOC_784/A AND2X1_LOC_568/B 0.02fF
C17742 OR2X1_LOC_59/Y OR2X1_LOC_767/a_8_216# 0.01fF
C17743 OR2X1_LOC_756/B AND2X1_LOC_104/a_8_24# 0.00fF
C17744 OR2X1_LOC_3/Y AND2X1_LOC_285/a_8_24# 0.00fF
C17745 OR2X1_LOC_3/Y OR2X1_LOC_13/Y 0.03fF
C17746 OR2X1_LOC_303/B OR2X1_LOC_365/B 0.02fF
C17747 OR2X1_LOC_368/a_8_216# OR2X1_LOC_7/A 0.03fF
C17748 OR2X1_LOC_62/A AND2X1_LOC_619/a_8_24# 0.15fF
C17749 OR2X1_LOC_673/B AND2X1_LOC_670/a_8_24# 0.04fF
C17750 AND2X1_LOC_768/a_8_24# OR2X1_LOC_26/Y 0.01fF
C17751 AND2X1_LOC_367/A AND2X1_LOC_114/a_8_24# 0.15fF
C17752 AND2X1_LOC_189/a_8_24# OR2X1_LOC_375/A 0.01fF
C17753 OR2X1_LOC_837/B OR2X1_LOC_837/a_8_216# 0.02fF
C17754 AND2X1_LOC_492/a_8_24# OR2X1_LOC_737/A 0.25fF
C17755 OR2X1_LOC_485/A OR2X1_LOC_96/Y 0.00fF
C17756 OR2X1_LOC_684/Y OR2X1_LOC_12/Y 0.39fF
C17757 OR2X1_LOC_136/Y D_INPUT_0 0.07fF
C17758 AND2X1_LOC_76/a_8_24# AND2X1_LOC_76/Y 0.02fF
C17759 OR2X1_LOC_160/B OR2X1_LOC_333/B 0.26fF
C17760 AND2X1_LOC_40/Y OR2X1_LOC_377/A 0.23fF
C17761 AND2X1_LOC_486/Y OR2X1_LOC_109/Y 0.03fF
C17762 AND2X1_LOC_383/a_8_24# OR2X1_LOC_417/A 0.08fF
C17763 AND2X1_LOC_22/Y AND2X1_LOC_107/a_36_24# 0.00fF
C17764 AND2X1_LOC_533/a_36_24# OR2X1_LOC_354/A 0.01fF
C17765 AND2X1_LOC_687/B OR2X1_LOC_16/A 0.13fF
C17766 OR2X1_LOC_469/Y OR2X1_LOC_375/A 0.03fF
C17767 AND2X1_LOC_214/A OR2X1_LOC_43/A 0.03fF
C17768 OR2X1_LOC_759/A OR2X1_LOC_258/Y 0.03fF
C17769 OR2X1_LOC_45/B OR2X1_LOC_504/Y 0.32fF
C17770 AND2X1_LOC_474/Y AND2X1_LOC_663/A 0.05fF
C17771 AND2X1_LOC_356/B AND2X1_LOC_434/Y 0.01fF
C17772 OR2X1_LOC_70/Y OR2X1_LOC_684/a_8_216# 0.02fF
C17773 OR2X1_LOC_51/Y AND2X1_LOC_155/Y 0.01fF
C17774 OR2X1_LOC_241/Y OR2X1_LOC_121/A 0.04fF
C17775 OR2X1_LOC_600/A OR2X1_LOC_481/A 0.03fF
C17776 OR2X1_LOC_780/A AND2X1_LOC_44/Y 0.09fF
C17777 AND2X1_LOC_181/a_8_24# OR2X1_LOC_7/A 0.01fF
C17778 AND2X1_LOC_716/Y AND2X1_LOC_303/B 0.52fF
C17779 OR2X1_LOC_623/a_8_216# OR2X1_LOC_161/A 0.03fF
C17780 VDD AND2X1_LOC_798/Y -0.00fF
C17781 OR2X1_LOC_118/a_36_216# OR2X1_LOC_71/Y 0.00fF
C17782 AND2X1_LOC_367/a_8_24# OR2X1_LOC_92/Y 0.01fF
C17783 OR2X1_LOC_748/A OR2X1_LOC_297/a_8_216# 0.01fF
C17784 OR2X1_LOC_532/B OR2X1_LOC_161/B 1.81fF
C17785 AND2X1_LOC_866/A GATE_579 0.01fF
C17786 AND2X1_LOC_845/Y OR2X1_LOC_12/Y 0.07fF
C17787 OR2X1_LOC_31/Y OR2X1_LOC_428/A 0.66fF
C17788 OR2X1_LOC_317/a_8_216# OR2X1_LOC_778/Y 0.33fF
C17789 AND2X1_LOC_337/B OR2X1_LOC_91/A 0.01fF
C17790 AND2X1_LOC_339/B INPUT_1 0.02fF
C17791 AND2X1_LOC_191/B OR2X1_LOC_282/Y 0.03fF
C17792 OR2X1_LOC_662/A OR2X1_LOC_185/A 0.45fF
C17793 AND2X1_LOC_675/A OR2X1_LOC_373/a_36_216# 0.02fF
C17794 OR2X1_LOC_377/A OR2X1_LOC_537/A 0.01fF
C17795 AND2X1_LOC_665/a_8_24# OR2X1_LOC_161/B 0.01fF
C17796 AND2X1_LOC_303/B AND2X1_LOC_654/Y -0.07fF
C17797 OR2X1_LOC_756/B AND2X1_LOC_3/Y 0.06fF
C17798 OR2X1_LOC_862/A OR2X1_LOC_810/A 0.77fF
C17799 OR2X1_LOC_481/A AND2X1_LOC_296/a_8_24# 0.00fF
C17800 OR2X1_LOC_31/Y OR2X1_LOC_595/A 0.03fF
C17801 AND2X1_LOC_228/Y AND2X1_LOC_175/B 0.02fF
C17802 OR2X1_LOC_459/a_8_216# AND2X1_LOC_43/B 0.06fF
C17803 AND2X1_LOC_843/Y AND2X1_LOC_859/Y 0.00fF
C17804 AND2X1_LOC_72/B OR2X1_LOC_115/B 0.26fF
C17805 OR2X1_LOC_155/A OR2X1_LOC_623/B 0.07fF
C17806 OR2X1_LOC_193/A OR2X1_LOC_78/B 0.44fF
C17807 AND2X1_LOC_512/Y AND2X1_LOC_390/B 1.38fF
C17808 VDD OR2X1_LOC_46/A 1.61fF
C17809 OR2X1_LOC_837/B OR2X1_LOC_52/B 0.03fF
C17810 AND2X1_LOC_348/A OR2X1_LOC_7/A 0.03fF
C17811 AND2X1_LOC_44/Y OR2X1_LOC_284/B 0.01fF
C17812 OR2X1_LOC_40/Y OR2X1_LOC_442/a_8_216# 0.07fF
C17813 AND2X1_LOC_840/a_8_24# OR2X1_LOC_238/Y 0.01fF
C17814 AND2X1_LOC_76/a_8_24# OR2X1_LOC_52/B 0.02fF
C17815 AND2X1_LOC_470/A AND2X1_LOC_470/B 0.09fF
C17816 AND2X1_LOC_515/a_36_24# OR2X1_LOC_95/Y 0.01fF
C17817 OR2X1_LOC_698/Y OR2X1_LOC_258/Y 0.23fF
C17818 AND2X1_LOC_36/Y OR2X1_LOC_80/A 0.15fF
C17819 AND2X1_LOC_44/Y D_INPUT_1 0.15fF
C17820 AND2X1_LOC_81/B OR2X1_LOC_510/Y 0.03fF
C17821 OR2X1_LOC_185/A OR2X1_LOC_631/B 0.39fF
C17822 OR2X1_LOC_235/B OR2X1_LOC_404/Y 0.00fF
C17823 OR2X1_LOC_502/A AND2X1_LOC_18/a_8_24# 0.02fF
C17824 OR2X1_LOC_743/A OR2X1_LOC_92/Y 0.12fF
C17825 OR2X1_LOC_252/Y OR2X1_LOC_36/Y 0.07fF
C17826 AND2X1_LOC_41/A OR2X1_LOC_713/a_8_216# 0.05fF
C17827 OR2X1_LOC_433/a_36_216# OR2X1_LOC_432/Y 0.00fF
C17828 OR2X1_LOC_669/Y OR2X1_LOC_278/Y 0.02fF
C17829 OR2X1_LOC_185/Y OR2X1_LOC_539/Y 0.07fF
C17830 OR2X1_LOC_554/a_8_216# OR2X1_LOC_598/A -0.01fF
C17831 OR2X1_LOC_799/A OR2X1_LOC_449/B 0.25fF
C17832 AND2X1_LOC_59/Y OR2X1_LOC_97/B 0.05fF
C17833 OR2X1_LOC_36/Y AND2X1_LOC_655/A 0.04fF
C17834 OR2X1_LOC_563/A OR2X1_LOC_493/Y 0.03fF
C17835 OR2X1_LOC_600/A OR2X1_LOC_71/Y 0.03fF
C17836 VDD OR2X1_LOC_679/A 0.21fF
C17837 AND2X1_LOC_36/Y AND2X1_LOC_419/a_8_24# 0.01fF
C17838 AND2X1_LOC_56/B OR2X1_LOC_130/A 0.07fF
C17839 OR2X1_LOC_91/A OR2X1_LOC_19/B 0.03fF
C17840 AND2X1_LOC_804/a_8_24# AND2X1_LOC_804/A -0.00fF
C17841 OR2X1_LOC_753/A OR2X1_LOC_38/a_36_216# 0.00fF
C17842 OR2X1_LOC_701/Y OR2X1_LOC_701/a_36_216# 0.00fF
C17843 OR2X1_LOC_22/Y AND2X1_LOC_434/Y 0.44fF
C17844 OR2X1_LOC_213/A OR2X1_LOC_213/B 0.13fF
C17845 OR2X1_LOC_248/A OR2X1_LOC_437/A 0.01fF
C17846 OR2X1_LOC_51/Y D_INPUT_0 0.04fF
C17847 OR2X1_LOC_358/A OR2X1_LOC_174/a_8_216# 0.05fF
C17848 OR2X1_LOC_275/a_8_216# OR2X1_LOC_517/A 0.48fF
C17849 AND2X1_LOC_40/Y AND2X1_LOC_670/a_8_24# 0.04fF
C17850 AND2X1_LOC_817/B OR2X1_LOC_269/B 0.05fF
C17851 AND2X1_LOC_215/Y OR2X1_LOC_31/Y 0.01fF
C17852 AND2X1_LOC_391/Y AND2X1_LOC_128/a_36_24# 0.05fF
C17853 AND2X1_LOC_8/Y OR2X1_LOC_130/A 0.02fF
C17854 OR2X1_LOC_223/A OR2X1_LOC_787/a_8_216# 0.01fF
C17855 VDD AND2X1_LOC_227/Y 0.44fF
C17856 AND2X1_LOC_508/B OR2X1_LOC_95/Y 0.03fF
C17857 OR2X1_LOC_802/Y OR2X1_LOC_809/a_8_216# 0.11fF
C17858 AND2X1_LOC_12/Y AND2X1_LOC_171/a_8_24# 0.01fF
C17859 OR2X1_LOC_532/B OR2X1_LOC_785/a_36_216# 0.02fF
C17860 OR2X1_LOC_574/A AND2X1_LOC_43/B 0.01fF
C17861 OR2X1_LOC_634/A AND2X1_LOC_825/a_8_24# 0.20fF
C17862 AND2X1_LOC_392/A AND2X1_LOC_476/A 0.07fF
C17863 D_INPUT_0 OR2X1_LOC_78/B 0.54fF
C17864 OR2X1_LOC_476/B OR2X1_LOC_640/A 0.01fF
C17865 OR2X1_LOC_305/Y AND2X1_LOC_702/Y 0.02fF
C17866 OR2X1_LOC_792/Y OR2X1_LOC_285/B 0.03fF
C17867 AND2X1_LOC_81/B OR2X1_LOC_810/A 0.06fF
C17868 AND2X1_LOC_12/Y AND2X1_LOC_387/B 0.03fF
C17869 OR2X1_LOC_43/A OR2X1_LOC_42/a_8_216# 0.03fF
C17870 OR2X1_LOC_69/a_8_216# OR2X1_LOC_52/B 0.01fF
C17871 OR2X1_LOC_132/a_8_216# OR2X1_LOC_95/Y 0.02fF
C17872 OR2X1_LOC_372/Y AND2X1_LOC_374/Y 0.21fF
C17873 OR2X1_LOC_666/A AND2X1_LOC_859/B 0.01fF
C17874 OR2X1_LOC_611/a_8_216# OR2X1_LOC_502/A 0.47fF
C17875 OR2X1_LOC_695/a_8_216# OR2X1_LOC_64/Y 0.02fF
C17876 OR2X1_LOC_339/A OR2X1_LOC_539/B 0.03fF
C17877 OR2X1_LOC_62/B OR2X1_LOC_736/A 0.03fF
C17878 AND2X1_LOC_47/Y AND2X1_LOC_628/a_8_24# 0.03fF
C17879 AND2X1_LOC_70/Y OR2X1_LOC_276/B 0.36fF
C17880 OR2X1_LOC_92/Y OR2X1_LOC_246/A 0.03fF
C17881 AND2X1_LOC_662/B AND2X1_LOC_662/a_8_24# 0.08fF
C17882 OR2X1_LOC_36/Y OR2X1_LOC_609/A 0.03fF
C17883 AND2X1_LOC_738/B AND2X1_LOC_796/Y 0.02fF
C17884 OR2X1_LOC_8/Y OR2X1_LOC_619/a_8_216# 0.01fF
C17885 OR2X1_LOC_600/A D_INPUT_1 0.06fF
C17886 AND2X1_LOC_796/Y OR2X1_LOC_56/A 0.14fF
C17887 AND2X1_LOC_660/Y OR2X1_LOC_39/A 0.02fF
C17888 OR2X1_LOC_43/A AND2X1_LOC_645/A 0.04fF
C17889 AND2X1_LOC_859/Y OR2X1_LOC_7/A 0.02fF
C17890 OR2X1_LOC_670/Y AND2X1_LOC_673/a_8_24# 0.23fF
C17891 D_INPUT_0 OR2X1_LOC_721/Y 0.10fF
C17892 OR2X1_LOC_251/Y OR2X1_LOC_106/A 0.03fF
C17893 OR2X1_LOC_193/A OR2X1_LOC_375/A 0.03fF
C17894 AND2X1_LOC_259/Y AND2X1_LOC_818/a_36_24# 0.00fF
C17895 OR2X1_LOC_654/A OR2X1_LOC_269/B 0.07fF
C17896 OR2X1_LOC_696/A AND2X1_LOC_247/a_8_24# 0.19fF
C17897 D_INPUT_4 AND2X1_LOC_7/Y 0.09fF
C17898 OR2X1_LOC_672/Y OR2X1_LOC_73/a_8_216# 0.45fF
C17899 VDD OR2X1_LOC_813/Y 0.00fF
C17900 OR2X1_LOC_631/a_8_216# OR2X1_LOC_62/B 0.01fF
C17901 OR2X1_LOC_759/A OR2X1_LOC_815/Y 0.02fF
C17902 OR2X1_LOC_40/Y AND2X1_LOC_846/a_8_24# 0.01fF
C17903 OR2X1_LOC_860/a_8_216# OR2X1_LOC_814/A 0.01fF
C17904 OR2X1_LOC_19/B AND2X1_LOC_573/A 0.03fF
C17905 AND2X1_LOC_191/Y AND2X1_LOC_569/a_36_24# 0.01fF
C17906 OR2X1_LOC_333/B OR2X1_LOC_219/B 0.25fF
C17907 OR2X1_LOC_856/a_36_216# OR2X1_LOC_269/B 0.00fF
C17908 AND2X1_LOC_182/A AND2X1_LOC_222/Y 0.01fF
C17909 OR2X1_LOC_337/A OR2X1_LOC_578/B 0.02fF
C17910 OR2X1_LOC_61/Y OR2X1_LOC_532/B 0.86fF
C17911 VDD OR2X1_LOC_41/Y 0.21fF
C17912 OR2X1_LOC_266/A OR2X1_LOC_71/A 0.14fF
C17913 AND2X1_LOC_191/B AND2X1_LOC_792/Y 0.01fF
C17914 OR2X1_LOC_246/A OR2X1_LOC_65/B 0.03fF
C17915 OR2X1_LOC_92/Y OR2X1_LOC_409/B 0.03fF
C17916 OR2X1_LOC_379/a_8_216# AND2X1_LOC_48/A 0.01fF
C17917 AND2X1_LOC_560/B AND2X1_LOC_663/B 4.54fF
C17918 AND2X1_LOC_42/a_8_24# AND2X1_LOC_42/B 0.06fF
C17919 AND2X1_LOC_470/a_36_24# OR2X1_LOC_619/Y 0.00fF
C17920 OR2X1_LOC_804/A AND2X1_LOC_92/Y 0.75fF
C17921 OR2X1_LOC_756/B OR2X1_LOC_270/Y 0.10fF
C17922 OR2X1_LOC_774/Y OR2X1_LOC_846/B 0.19fF
C17923 OR2X1_LOC_808/B OR2X1_LOC_223/A 0.03fF
C17924 AND2X1_LOC_59/Y OR2X1_LOC_814/A 0.17fF
C17925 OR2X1_LOC_596/A OR2X1_LOC_715/a_36_216# 0.00fF
C17926 D_INPUT_7 OR2X1_LOC_17/Y 0.01fF
C17927 AND2X1_LOC_536/a_8_24# OR2X1_LOC_532/B 0.01fF
C17928 OR2X1_LOC_508/Y OR2X1_LOC_510/a_8_216# 0.02fF
C17929 VDD OR2X1_LOC_753/Y 0.23fF
C17930 OR2X1_LOC_88/Y AND2X1_LOC_243/Y 0.01fF
C17931 AND2X1_LOC_13/a_36_24# OR2X1_LOC_155/A 0.01fF
C17932 OR2X1_LOC_344/A AND2X1_LOC_268/a_8_24# 0.20fF
C17933 D_INPUT_0 OR2X1_LOC_375/A 0.27fF
C17934 AND2X1_LOC_489/a_8_24# AND2X1_LOC_563/Y 0.01fF
C17935 AND2X1_LOC_276/Y AND2X1_LOC_473/a_8_24# 0.14fF
C17936 D_INPUT_5 OR2X1_LOC_50/a_8_216# 0.01fF
C17937 AND2X1_LOC_56/B OR2X1_LOC_62/B 0.01fF
C17938 OR2X1_LOC_659/B OR2X1_LOC_62/B 0.02fF
C17939 OR2X1_LOC_821/a_8_216# OR2X1_LOC_13/B 0.01fF
C17940 AND2X1_LOC_671/a_8_24# OR2X1_LOC_753/A 0.04fF
C17941 OR2X1_LOC_70/Y OR2X1_LOC_430/a_8_216# 0.02fF
C17942 AND2X1_LOC_824/B AND2X1_LOC_826/a_8_24# 0.20fF
C17943 OR2X1_LOC_417/A AND2X1_LOC_458/Y 0.03fF
C17944 AND2X1_LOC_22/Y OR2X1_LOC_593/B 0.03fF
C17945 OR2X1_LOC_43/A AND2X1_LOC_477/A 0.03fF
C17946 AND2X1_LOC_8/Y OR2X1_LOC_62/B 0.21fF
C17947 OR2X1_LOC_809/B AND2X1_LOC_31/Y 0.07fF
C17948 OR2X1_LOC_516/Y AND2X1_LOC_242/B 0.09fF
C17949 OR2X1_LOC_863/B AND2X1_LOC_51/Y 0.01fF
C17950 OR2X1_LOC_487/Y AND2X1_LOC_849/A 0.23fF
C17951 AND2X1_LOC_61/Y AND2X1_LOC_215/a_8_24# 0.04fF
C17952 OR2X1_LOC_154/A OR2X1_LOC_436/Y 0.03fF
C17953 OR2X1_LOC_864/A OR2X1_LOC_655/B 0.02fF
C17954 OR2X1_LOC_447/Y OR2X1_LOC_449/A 0.07fF
C17955 OR2X1_LOC_538/A OR2X1_LOC_854/A 0.02fF
C17956 OR2X1_LOC_47/Y AND2X1_LOC_403/B 0.01fF
C17957 AND2X1_LOC_831/Y AND2X1_LOC_831/a_36_24# 0.01fF
C17958 OR2X1_LOC_619/Y D_INPUT_1 0.14fF
C17959 AND2X1_LOC_170/Y AND2X1_LOC_170/B 0.01fF
C17960 AND2X1_LOC_227/Y AND2X1_LOC_267/a_8_24# 0.01fF
C17961 OR2X1_LOC_64/Y AND2X1_LOC_663/B 0.05fF
C17962 OR2X1_LOC_477/B OR2X1_LOC_477/a_36_216# 0.00fF
C17963 OR2X1_LOC_117/Y OR2X1_LOC_95/Y 0.07fF
C17964 AND2X1_LOC_1/Y AND2X1_LOC_31/a_8_24# -0.00fF
C17965 OR2X1_LOC_62/B OR2X1_LOC_291/A 0.03fF
C17966 OR2X1_LOC_223/a_8_216# OR2X1_LOC_564/B 0.40fF
C17967 AND2X1_LOC_64/Y AND2X1_LOC_7/B 0.32fF
C17968 OR2X1_LOC_450/A OR2X1_LOC_707/a_8_216# 0.03fF
C17969 AND2X1_LOC_22/Y AND2X1_LOC_273/a_8_24# 0.01fF
C17970 OR2X1_LOC_848/a_8_216# D_INPUT_1 0.01fF
C17971 OR2X1_LOC_47/Y OR2X1_LOC_44/Y 9.11fF
C17972 AND2X1_LOC_564/A AND2X1_LOC_192/a_8_24# 0.20fF
C17973 OR2X1_LOC_440/A OR2X1_LOC_733/B 0.20fF
C17974 OR2X1_LOC_510/Y OR2X1_LOC_66/Y 0.01fF
C17975 AND2X1_LOC_41/A OR2X1_LOC_705/a_8_216# 0.01fF
C17976 AND2X1_LOC_56/B AND2X1_LOC_39/Y 0.04fF
C17977 OR2X1_LOC_600/A AND2X1_LOC_789/Y 0.15fF
C17978 AND2X1_LOC_12/Y OR2X1_LOC_318/B 0.03fF
C17979 OR2X1_LOC_280/Y AND2X1_LOC_851/B 0.16fF
C17980 OR2X1_LOC_36/Y OR2X1_LOC_599/Y 0.03fF
C17981 OR2X1_LOC_510/A OR2X1_LOC_508/Y 0.01fF
C17982 OR2X1_LOC_53/Y OR2X1_LOC_43/Y 0.00fF
C17983 OR2X1_LOC_599/A AND2X1_LOC_644/a_8_24# 0.00fF
C17984 OR2X1_LOC_26/Y OR2X1_LOC_41/a_8_216# 0.01fF
C17985 AND2X1_LOC_687/Y AND2X1_LOC_687/B 0.01fF
C17986 OR2X1_LOC_70/Y OR2X1_LOC_428/Y 0.01fF
C17987 OR2X1_LOC_78/B OR2X1_LOC_339/A 0.19fF
C17988 D_INPUT_2 OR2X1_LOC_8/a_8_216# 0.03fF
C17989 AND2X1_LOC_500/a_8_24# OR2X1_LOC_419/Y 0.01fF
C17990 AND2X1_LOC_812/a_36_24# OR2X1_LOC_74/A 0.01fF
C17991 OR2X1_LOC_231/a_8_216# OR2X1_LOC_68/B 0.02fF
C17992 AND2X1_LOC_523/Y OR2X1_LOC_95/Y 0.01fF
C17993 OR2X1_LOC_160/A AND2X1_LOC_31/Y 5.25fF
C17994 AND2X1_LOC_711/a_8_24# AND2X1_LOC_789/Y 0.01fF
C17995 OR2X1_LOC_810/A OR2X1_LOC_66/Y 0.05fF
C17996 OR2X1_LOC_92/Y OR2X1_LOC_599/a_8_216# 0.03fF
C17997 OR2X1_LOC_841/B OR2X1_LOC_318/B 0.01fF
C17998 OR2X1_LOC_756/B OR2X1_LOC_576/a_8_216# 0.01fF
C17999 AND2X1_LOC_59/Y OR2X1_LOC_341/a_8_216# 0.06fF
C18000 OR2X1_LOC_188/Y OR2X1_LOC_549/A 0.03fF
C18001 AND2X1_LOC_80/a_8_24# OR2X1_LOC_68/B 0.01fF
C18002 OR2X1_LOC_175/Y OR2X1_LOC_151/A 0.10fF
C18003 AND2X1_LOC_858/B OR2X1_LOC_504/a_8_216# 0.04fF
C18004 OR2X1_LOC_632/Y OR2X1_LOC_844/B 0.02fF
C18005 AND2X1_LOC_53/Y AND2X1_LOC_692/a_36_24# 0.01fF
C18006 OR2X1_LOC_323/A AND2X1_LOC_112/a_36_24# 0.00fF
C18007 AND2X1_LOC_95/Y OR2X1_LOC_501/a_8_216# 0.01fF
C18008 OR2X1_LOC_53/Y AND2X1_LOC_207/A 0.01fF
C18009 AND2X1_LOC_82/a_36_24# OR2X1_LOC_68/B 0.00fF
C18010 OR2X1_LOC_22/Y AND2X1_LOC_851/B 0.01fF
C18011 OR2X1_LOC_712/a_36_216# OR2X1_LOC_712/B 0.03fF
C18012 OR2X1_LOC_40/Y GATE_579 0.02fF
C18013 AND2X1_LOC_809/A OR2X1_LOC_13/B 0.10fF
C18014 AND2X1_LOC_468/B OR2X1_LOC_437/A 0.00fF
C18015 AND2X1_LOC_17/Y AND2X1_LOC_430/B 0.01fF
C18016 OR2X1_LOC_840/A AND2X1_LOC_36/Y 0.14fF
C18017 AND2X1_LOC_40/Y OR2X1_LOC_539/B 0.02fF
C18018 OR2X1_LOC_139/A AND2X1_LOC_110/Y 0.06fF
C18019 OR2X1_LOC_756/B OR2X1_LOC_388/a_8_216# 0.01fF
C18020 OR2X1_LOC_294/Y OR2X1_LOC_346/A 0.01fF
C18021 OR2X1_LOC_804/B OR2X1_LOC_318/B 0.01fF
C18022 OR2X1_LOC_680/a_8_216# OR2X1_LOC_51/Y 0.16fF
C18023 OR2X1_LOC_630/Y OR2X1_LOC_115/B 0.12fF
C18024 OR2X1_LOC_632/a_8_216# OR2X1_LOC_140/B 0.01fF
C18025 AND2X1_LOC_227/Y OR2X1_LOC_256/A 0.00fF
C18026 OR2X1_LOC_308/A OR2X1_LOC_834/A 0.04fF
C18027 OR2X1_LOC_186/Y OR2X1_LOC_715/B 0.19fF
C18028 OR2X1_LOC_53/Y OR2X1_LOC_690/Y 0.00fF
C18029 AND2X1_LOC_8/a_36_24# OR2X1_LOC_54/Y 0.00fF
C18030 OR2X1_LOC_177/Y AND2X1_LOC_719/Y 0.03fF
C18031 OR2X1_LOC_600/A OR2X1_LOC_15/a_8_216# 0.02fF
C18032 AND2X1_LOC_191/B AND2X1_LOC_287/B 0.01fF
C18033 OR2X1_LOC_45/B AND2X1_LOC_658/B 0.03fF
C18034 OR2X1_LOC_509/a_8_216# AND2X1_LOC_65/A 0.03fF
C18035 OR2X1_LOC_85/A OR2X1_LOC_150/a_36_216# 0.03fF
C18036 OR2X1_LOC_176/Y AND2X1_LOC_436/Y 0.00fF
C18037 OR2X1_LOC_816/A AND2X1_LOC_657/Y 0.03fF
C18038 OR2X1_LOC_800/Y OR2X1_LOC_138/A 0.00fF
C18039 OR2X1_LOC_46/A OR2X1_LOC_67/Y 0.10fF
C18040 AND2X1_LOC_191/B OR2X1_LOC_816/A 0.98fF
C18041 OR2X1_LOC_449/B OR2X1_LOC_446/B 0.06fF
C18042 AND2X1_LOC_350/B OR2X1_LOC_51/Y 0.50fF
C18043 AND2X1_LOC_64/Y OR2X1_LOC_319/B 0.18fF
C18044 OR2X1_LOC_22/Y AND2X1_LOC_461/a_36_24# 0.01fF
C18045 OR2X1_LOC_134/Y OR2X1_LOC_517/A 0.05fF
C18046 AND2X1_LOC_332/a_8_24# AND2X1_LOC_326/B 0.00fF
C18047 AND2X1_LOC_842/a_8_24# AND2X1_LOC_242/B 0.01fF
C18048 OR2X1_LOC_22/Y OR2X1_LOC_595/Y 0.02fF
C18049 AND2X1_LOC_91/B OR2X1_LOC_841/a_8_216# 0.28fF
C18050 AND2X1_LOC_541/Y AND2X1_LOC_553/a_8_24# 0.05fF
C18051 OR2X1_LOC_347/A AND2X1_LOC_95/Y 0.01fF
C18052 OR2X1_LOC_709/A AND2X1_LOC_70/Y 0.04fF
C18053 OR2X1_LOC_585/A OR2X1_LOC_536/a_8_216# 0.01fF
C18054 AND2X1_LOC_22/Y AND2X1_LOC_306/a_36_24# 0.00fF
C18055 AND2X1_LOC_722/a_8_24# OR2X1_LOC_40/Y 0.02fF
C18056 OR2X1_LOC_369/a_8_216# OR2X1_LOC_309/a_8_216# 0.47fF
C18057 OR2X1_LOC_97/A OR2X1_LOC_174/A 0.01fF
C18058 AND2X1_LOC_64/Y OR2X1_LOC_318/Y 7.13fF
C18059 OR2X1_LOC_51/Y AND2X1_LOC_771/B 0.01fF
C18060 OR2X1_LOC_476/a_8_216# OR2X1_LOC_228/Y 0.01fF
C18061 VDD OR2X1_LOC_786/a_8_216# 0.21fF
C18062 OR2X1_LOC_256/A OR2X1_LOC_813/Y 0.03fF
C18063 OR2X1_LOC_6/B AND2X1_LOC_18/Y 0.64fF
C18064 OR2X1_LOC_345/A OR2X1_LOC_345/a_8_216# 0.47fF
C18065 OR2X1_LOC_108/a_8_216# OR2X1_LOC_600/A 0.01fF
C18066 OR2X1_LOC_753/A OR2X1_LOC_248/A 0.01fF
C18067 OR2X1_LOC_125/a_8_216# OR2X1_LOC_40/Y 0.01fF
C18068 AND2X1_LOC_232/a_36_24# OR2X1_LOC_633/A 0.01fF
C18069 AND2X1_LOC_47/Y OR2X1_LOC_247/Y 0.02fF
C18070 VDD INPUT_2 0.23fF
C18071 AND2X1_LOC_12/Y OR2X1_LOC_363/a_8_216# 0.01fF
C18072 OR2X1_LOC_158/A OR2X1_LOC_59/Y 0.22fF
C18073 OR2X1_LOC_660/a_8_216# AND2X1_LOC_22/Y 0.05fF
C18074 OR2X1_LOC_703/B OR2X1_LOC_168/Y 0.04fF
C18075 AND2X1_LOC_363/B OR2X1_LOC_428/A 0.01fF
C18076 OR2X1_LOC_108/a_36_216# OR2X1_LOC_56/A 0.00fF
C18077 OR2X1_LOC_135/Y AND2X1_LOC_857/Y 0.03fF
C18078 OR2X1_LOC_426/B OR2X1_LOC_600/A 0.07fF
C18079 AND2X1_LOC_794/A AND2X1_LOC_794/a_8_24# 0.19fF
C18080 OR2X1_LOC_426/B AND2X1_LOC_335/Y 0.03fF
C18081 AND2X1_LOC_64/Y OR2X1_LOC_805/A 0.10fF
C18082 OR2X1_LOC_9/Y OR2X1_LOC_235/B 0.34fF
C18083 OR2X1_LOC_789/a_8_216# AND2X1_LOC_36/Y 0.02fF
C18084 AND2X1_LOC_830/a_8_24# OR2X1_LOC_437/A 0.01fF
C18085 AND2X1_LOC_2/Y VDD 0.52fF
C18086 OR2X1_LOC_140/A OR2X1_LOC_78/A 0.02fF
C18087 OR2X1_LOC_316/a_8_216# OR2X1_LOC_85/A 0.01fF
C18088 OR2X1_LOC_235/B OR2X1_LOC_362/A 0.02fF
C18089 AND2X1_LOC_794/B AND2X1_LOC_722/A 0.07fF
C18090 OR2X1_LOC_600/Y AND2X1_LOC_447/Y 0.05fF
C18091 AND2X1_LOC_505/a_8_24# OR2X1_LOC_78/B 0.03fF
C18092 OR2X1_LOC_507/A OR2X1_LOC_78/A 0.01fF
C18093 VDD OR2X1_LOC_792/B 0.00fF
C18094 AND2X1_LOC_773/Y AND2X1_LOC_76/Y 0.03fF
C18095 OR2X1_LOC_653/Y AND2X1_LOC_60/a_36_24# 0.00fF
C18096 OR2X1_LOC_653/B OR2X1_LOC_502/A 0.02fF
C18097 AND2X1_LOC_721/Y AND2X1_LOC_621/Y 0.03fF
C18098 OR2X1_LOC_121/B OR2X1_LOC_303/B 0.07fF
C18099 OR2X1_LOC_614/Y OR2X1_LOC_502/A 0.02fF
C18100 AND2X1_LOC_95/Y AND2X1_LOC_44/Y 2.93fF
C18101 AND2X1_LOC_40/Y OR2X1_LOC_812/a_8_216# 0.01fF
C18102 OR2X1_LOC_427/A OR2X1_LOC_373/Y 0.03fF
C18103 OR2X1_LOC_109/Y AND2X1_LOC_457/a_8_24# 0.02fF
C18104 OR2X1_LOC_666/A OR2X1_LOC_56/A 0.00fF
C18105 AND2X1_LOC_523/a_36_24# OR2X1_LOC_428/A 0.00fF
C18106 VDD OR2X1_LOC_107/Y 0.16fF
C18107 OR2X1_LOC_633/Y AND2X1_LOC_44/Y 0.03fF
C18108 AND2X1_LOC_568/B AND2X1_LOC_365/a_8_24# 0.01fF
C18109 AND2X1_LOC_772/B OR2X1_LOC_744/A 0.05fF
C18110 OR2X1_LOC_479/Y OR2X1_LOC_308/Y 0.07fF
C18111 AND2X1_LOC_866/A AND2X1_LOC_657/A 0.07fF
C18112 AND2X1_LOC_47/Y OR2X1_LOC_364/Y 0.01fF
C18113 OR2X1_LOC_11/Y OR2X1_LOC_18/a_8_216# 0.02fF
C18114 AND2X1_LOC_721/Y AND2X1_LOC_668/a_8_24# 0.20fF
C18115 OR2X1_LOC_151/A OR2X1_LOC_629/Y 0.14fF
C18116 OR2X1_LOC_231/B AND2X1_LOC_12/Y 0.05fF
C18117 OR2X1_LOC_759/A OR2X1_LOC_698/Y 0.55fF
C18118 AND2X1_LOC_740/B AND2X1_LOC_220/B 0.03fF
C18119 VDD AND2X1_LOC_722/A 0.10fF
C18120 AND2X1_LOC_848/A AND2X1_LOC_792/Y 0.08fF
C18121 AND2X1_LOC_611/a_8_24# OR2X1_LOC_415/Y 0.13fF
C18122 AND2X1_LOC_70/Y OR2X1_LOC_703/A 0.03fF
C18123 AND2X1_LOC_364/Y AND2X1_LOC_514/a_8_24# 0.20fF
C18124 AND2X1_LOC_315/a_8_24# OR2X1_LOC_486/Y 0.05fF
C18125 AND2X1_LOC_729/Y OR2X1_LOC_12/Y 0.00fF
C18126 OR2X1_LOC_121/Y AND2X1_LOC_12/Y 0.08fF
C18127 AND2X1_LOC_3/Y OR2X1_LOC_140/B 0.04fF
C18128 OR2X1_LOC_615/Y AND2X1_LOC_793/B 0.00fF
C18129 INPUT_1 OR2X1_LOC_300/Y 0.54fF
C18130 OR2X1_LOC_673/B OR2X1_LOC_375/A 0.06fF
C18131 OR2X1_LOC_89/A AND2X1_LOC_227/a_8_24# 0.01fF
C18132 AND2X1_LOC_534/a_36_24# AND2X1_LOC_43/B 0.01fF
C18133 AND2X1_LOC_512/Y OR2X1_LOC_744/A 0.07fF
C18134 OR2X1_LOC_490/Y AND2X1_LOC_772/Y 0.02fF
C18135 AND2X1_LOC_64/Y OR2X1_LOC_296/Y 0.01fF
C18136 OR2X1_LOC_523/Y AND2X1_LOC_18/Y 0.01fF
C18137 OR2X1_LOC_99/Y AND2X1_LOC_44/Y 0.03fF
C18138 AND2X1_LOC_12/Y OR2X1_LOC_351/B 0.03fF
C18139 AND2X1_LOC_42/B OR2X1_LOC_831/B 0.06fF
C18140 AND2X1_LOC_716/Y OR2X1_LOC_56/A 0.07fF
C18141 OR2X1_LOC_597/A OR2X1_LOC_48/B 0.12fF
C18142 OR2X1_LOC_505/a_8_216# AND2X1_LOC_806/A 0.01fF
C18143 AND2X1_LOC_720/Y OR2X1_LOC_59/Y 0.01fF
C18144 OR2X1_LOC_188/a_8_216# AND2X1_LOC_42/B 0.00fF
C18145 AND2X1_LOC_773/Y OR2X1_LOC_52/B 0.02fF
C18146 AND2X1_LOC_784/A OR2X1_LOC_12/Y 0.19fF
C18147 AND2X1_LOC_658/A OR2X1_LOC_628/a_8_216# 0.03fF
C18148 AND2X1_LOC_211/B OR2X1_LOC_310/a_8_216# 0.03fF
C18149 AND2X1_LOC_50/Y AND2X1_LOC_70/a_36_24# 0.00fF
C18150 AND2X1_LOC_40/Y OR2X1_LOC_78/B 0.91fF
C18151 OR2X1_LOC_51/Y AND2X1_LOC_840/A -0.01fF
C18152 OR2X1_LOC_597/A OR2X1_LOC_18/Y 0.01fF
C18153 OR2X1_LOC_235/B OR2X1_LOC_474/Y 0.07fF
C18154 OR2X1_LOC_161/A OR2X1_LOC_733/A 0.14fF
C18155 OR2X1_LOC_67/A AND2X1_LOC_243/Y 0.04fF
C18156 OR2X1_LOC_860/a_8_216# OR2X1_LOC_244/Y 0.02fF
C18157 AND2X1_LOC_638/Y OR2X1_LOC_762/Y 0.14fF
C18158 OR2X1_LOC_604/A OR2X1_LOC_252/Y 0.01fF
C18159 AND2X1_LOC_12/Y OR2X1_LOC_114/B 0.03fF
C18160 OR2X1_LOC_461/B AND2X1_LOC_233/a_8_24# 0.20fF
C18161 OR2X1_LOC_105/a_8_216# OR2X1_LOC_571/a_8_216# 0.47fF
C18162 OR2X1_LOC_105/Y OR2X1_LOC_561/Y 0.01fF
C18163 AND2X1_LOC_654/Y OR2X1_LOC_56/A 0.16fF
C18164 OR2X1_LOC_604/A OR2X1_LOC_313/Y 0.02fF
C18165 VDD OR2X1_LOC_739/A 0.49fF
C18166 AND2X1_LOC_31/Y OR2X1_LOC_717/a_8_216# 0.01fF
C18167 OR2X1_LOC_715/B AND2X1_LOC_81/B 0.03fF
C18168 OR2X1_LOC_653/Y OR2X1_LOC_78/A 0.10fF
C18169 OR2X1_LOC_218/a_8_216# AND2X1_LOC_65/A 0.03fF
C18170 OR2X1_LOC_666/A AND2X1_LOC_850/Y 0.02fF
C18171 OR2X1_LOC_426/B OR2X1_LOC_619/Y 0.08fF
C18172 VDD AND2X1_LOC_454/Y 0.21fF
C18173 OR2X1_LOC_158/A OR2X1_LOC_820/B 0.05fF
C18174 OR2X1_LOC_185/A OR2X1_LOC_648/A 0.07fF
C18175 AND2X1_LOC_388/Y AND2X1_LOC_661/A 0.03fF
C18176 AND2X1_LOC_541/a_8_24# AND2X1_LOC_663/B 0.05fF
C18177 OR2X1_LOC_49/A OR2X1_LOC_3/Y 0.32fF
C18178 OR2X1_LOC_860/Y OR2X1_LOC_756/B 0.01fF
C18179 AND2X1_LOC_769/a_8_24# OR2X1_LOC_12/Y 0.01fF
C18180 OR2X1_LOC_479/Y AND2X1_LOC_604/a_8_24# 0.06fF
C18181 OR2X1_LOC_154/A OR2X1_LOC_160/B 2.91fF
C18182 OR2X1_LOC_808/B OR2X1_LOC_502/A 0.01fF
C18183 AND2X1_LOC_541/Y OR2X1_LOC_26/Y 0.01fF
C18184 AND2X1_LOC_640/Y OR2X1_LOC_16/A 0.01fF
C18185 AND2X1_LOC_298/a_8_24# OR2X1_LOC_302/A 0.08fF
C18186 AND2X1_LOC_165/a_36_24# OR2X1_LOC_449/B 0.00fF
C18187 OR2X1_LOC_696/A OR2X1_LOC_226/a_8_216# 0.04fF
C18188 OR2X1_LOC_241/Y AND2X1_LOC_36/Y 0.07fF
C18189 AND2X1_LOC_564/B AND2X1_LOC_464/Y 0.01fF
C18190 AND2X1_LOC_779/Y AND2X1_LOC_783/a_8_24# 0.19fF
C18191 AND2X1_LOC_732/B OR2X1_LOC_44/Y 0.01fF
C18192 AND2X1_LOC_392/A AND2X1_LOC_560/B 0.07fF
C18193 OR2X1_LOC_206/A AND2X1_LOC_7/B 0.01fF
C18194 OR2X1_LOC_426/B OR2X1_LOC_88/A 0.25fF
C18195 AND2X1_LOC_91/B OR2X1_LOC_383/Y 0.05fF
C18196 OR2X1_LOC_599/A VDD 0.02fF
C18197 OR2X1_LOC_160/B OR2X1_LOC_267/A 0.01fF
C18198 OR2X1_LOC_130/A AND2X1_LOC_92/Y 0.18fF
C18199 OR2X1_LOC_8/Y AND2X1_LOC_342/a_8_24# 0.01fF
C18200 AND2X1_LOC_150/a_8_24# AND2X1_LOC_42/B 0.03fF
C18201 OR2X1_LOC_744/A AND2X1_LOC_342/Y 0.39fF
C18202 AND2X1_LOC_751/a_8_24# OR2X1_LOC_789/A 0.01fF
C18203 VDD OR2X1_LOC_269/B 2.36fF
C18204 AND2X1_LOC_182/A OR2X1_LOC_74/A 0.07fF
C18205 OR2X1_LOC_426/A OR2X1_LOC_427/A 0.42fF
C18206 AND2X1_LOC_308/a_8_24# OR2X1_LOC_428/A 0.04fF
C18207 OR2X1_LOC_528/Y AND2X1_LOC_475/a_8_24# 0.01fF
C18208 VDD OR2X1_LOC_93/a_8_216# 0.00fF
C18209 OR2X1_LOC_116/a_8_216# AND2X1_LOC_70/Y 0.01fF
C18210 OR2X1_LOC_90/a_8_216# OR2X1_LOC_85/A 0.02fF
C18211 OR2X1_LOC_756/B OR2X1_LOC_489/B 0.00fF
C18212 GATE_366 OR2X1_LOC_56/A 0.07fF
C18213 AND2X1_LOC_649/B AND2X1_LOC_642/Y 0.01fF
C18214 AND2X1_LOC_710/Y GATE_366 0.03fF
C18215 AND2X1_LOC_712/Y OR2X1_LOC_3/Y 0.01fF
C18216 OR2X1_LOC_185/A AND2X1_LOC_253/a_8_24# 0.01fF
C18217 INPUT_0 AND2X1_LOC_55/a_8_24# 0.02fF
C18218 OR2X1_LOC_128/A OR2X1_LOC_736/A 0.01fF
C18219 OR2X1_LOC_158/A OR2X1_LOC_70/Y 0.10fF
C18220 AND2X1_LOC_175/B AND2X1_LOC_857/Y 0.01fF
C18221 OR2X1_LOC_809/B OR2X1_LOC_809/a_8_216# 0.02fF
C18222 AND2X1_LOC_704/a_36_24# OR2X1_LOC_70/Y -0.00fF
C18223 OR2X1_LOC_377/A AND2X1_LOC_39/a_8_24# 0.01fF
C18224 AND2X1_LOC_70/Y AND2X1_LOC_17/Y 0.42fF
C18225 OR2X1_LOC_297/a_36_216# AND2X1_LOC_847/Y 0.01fF
C18226 OR2X1_LOC_124/B AND2X1_LOC_3/Y 0.03fF
C18227 AND2X1_LOC_347/Y AND2X1_LOC_848/Y 0.80fF
C18228 OR2X1_LOC_416/Y OR2X1_LOC_16/A 0.05fF
C18229 OR2X1_LOC_40/Y AND2X1_LOC_728/a_8_24# 0.06fF
C18230 AND2X1_LOC_12/Y D_INPUT_5 0.01fF
C18231 AND2X1_LOC_734/Y OR2X1_LOC_406/a_8_216# 0.48fF
C18232 OR2X1_LOC_519/a_8_216# AND2X1_LOC_364/A 0.02fF
C18233 OR2X1_LOC_798/Y OR2X1_LOC_539/Y 0.44fF
C18234 VDD OR2X1_LOC_258/a_8_216# 0.21fF
C18235 OR2X1_LOC_848/a_8_216# OR2X1_LOC_391/a_8_216# 0.47fF
C18236 OR2X1_LOC_748/A OR2X1_LOC_820/A 0.39fF
C18237 VDD OR2X1_LOC_546/B 0.00fF
C18238 OR2X1_LOC_850/B OR2X1_LOC_664/Y 0.00fF
C18239 AND2X1_LOC_40/Y OR2X1_LOC_375/A 6.37fF
C18240 AND2X1_LOC_570/Y OR2X1_LOC_529/Y 0.97fF
C18241 OR2X1_LOC_405/A AND2X1_LOC_314/a_8_24# 0.02fF
C18242 OR2X1_LOC_235/B AND2X1_LOC_852/Y 0.07fF
C18243 AND2X1_LOC_639/A OR2X1_LOC_12/Y 0.02fF
C18244 INPUT_1 AND2X1_LOC_219/A 0.04fF
C18245 OR2X1_LOC_160/B OR2X1_LOC_778/A 0.10fF
C18246 AND2X1_LOC_753/a_8_24# OR2X1_LOC_790/B 0.01fF
C18247 AND2X1_LOC_154/Y AND2X1_LOC_658/A 0.57fF
C18248 AND2X1_LOC_350/a_8_24# OR2X1_LOC_46/A 0.01fF
C18249 OR2X1_LOC_589/A OR2X1_LOC_245/a_8_216# 0.01fF
C18250 OR2X1_LOC_753/A OR2X1_LOC_234/Y 0.05fF
C18251 OR2X1_LOC_158/A AND2X1_LOC_514/Y 0.07fF
C18252 AND2X1_LOC_156/a_8_24# AND2X1_LOC_658/a_8_24# 0.23fF
C18253 AND2X1_LOC_70/Y OR2X1_LOC_653/a_8_216# 0.00fF
C18254 AND2X1_LOC_675/Y AND2X1_LOC_474/Y 0.02fF
C18255 OR2X1_LOC_614/Y AND2X1_LOC_48/A 0.00fF
C18256 OR2X1_LOC_807/Y OR2X1_LOC_805/A 0.02fF
C18257 OR2X1_LOC_756/B OR2X1_LOC_592/a_36_216# 0.00fF
C18258 OR2X1_LOC_715/B OR2X1_LOC_196/B 0.00fF
C18259 AND2X1_LOC_392/A OR2X1_LOC_64/Y 0.22fF
C18260 INPUT_4 OR2X1_LOC_427/A 1.20fF
C18261 OR2X1_LOC_86/Y OR2X1_LOC_92/Y 0.01fF
C18262 D_INPUT_0 OR2X1_LOC_549/A 0.26fF
C18263 OR2X1_LOC_377/A AND2X1_LOC_43/B 0.24fF
C18264 OR2X1_LOC_502/A OR2X1_LOC_708/B 0.00fF
C18265 OR2X1_LOC_471/a_8_216# OR2X1_LOC_375/A 0.03fF
C18266 OR2X1_LOC_40/Y AND2X1_LOC_326/a_8_24# 0.02fF
C18267 AND2X1_LOC_318/Y AND2X1_LOC_476/a_36_24# 0.01fF
C18268 AND2X1_LOC_141/B OR2X1_LOC_744/A 0.04fF
C18269 AND2X1_LOC_31/Y OR2X1_LOC_212/B 0.17fF
C18270 OR2X1_LOC_600/A OR2X1_LOC_125/Y 0.03fF
C18271 OR2X1_LOC_506/Y OR2X1_LOC_241/Y 0.10fF
C18272 AND2X1_LOC_53/Y OR2X1_LOC_596/A 0.07fF
C18273 OR2X1_LOC_469/Y OR2X1_LOC_711/A 0.17fF
C18274 OR2X1_LOC_641/Y AND2X1_LOC_518/a_8_24# 0.01fF
C18275 OR2X1_LOC_516/B OR2X1_LOC_485/A 0.23fF
C18276 AND2X1_LOC_824/B AND2X1_LOC_43/B 0.07fF
C18277 OR2X1_LOC_306/Y AND2X1_LOC_655/A 0.05fF
C18278 OR2X1_LOC_87/A OR2X1_LOC_796/a_8_216# 0.05fF
C18279 OR2X1_LOC_45/B OR2X1_LOC_47/Y 5.07fF
C18280 OR2X1_LOC_49/A OR2X1_LOC_673/A 0.05fF
C18281 OR2X1_LOC_625/Y OR2X1_LOC_44/Y 0.07fF
C18282 OR2X1_LOC_51/Y AND2X1_LOC_687/A 0.19fF
C18283 AND2X1_LOC_186/a_36_24# AND2X1_LOC_624/A 0.00fF
C18284 OR2X1_LOC_641/Y AND2X1_LOC_48/A 0.35fF
C18285 OR2X1_LOC_114/Y OR2X1_LOC_161/A 0.03fF
C18286 AND2X1_LOC_592/Y OR2X1_LOC_31/Y 0.01fF
C18287 OR2X1_LOC_251/Y OR2X1_LOC_250/a_8_216# 0.03fF
C18288 AND2X1_LOC_784/A AND2X1_LOC_170/a_8_24# 0.03fF
C18289 OR2X1_LOC_600/A OR2X1_LOC_225/a_8_216# -0.01fF
C18290 AND2X1_LOC_647/Y AND2X1_LOC_772/Y 0.01fF
C18291 OR2X1_LOC_516/A AND2X1_LOC_840/B 0.03fF
C18292 OR2X1_LOC_468/Y OR2X1_LOC_738/A 0.01fF
C18293 OR2X1_LOC_529/a_8_216# OR2X1_LOC_26/Y 0.01fF
C18294 OR2X1_LOC_203/Y AND2X1_LOC_43/B 0.07fF
C18295 AND2X1_LOC_727/A AND2X1_LOC_469/B 0.03fF
C18296 OR2X1_LOC_849/A OR2X1_LOC_624/A 0.01fF
C18297 AND2X1_LOC_742/a_36_24# GATE_811 0.00fF
C18298 OR2X1_LOC_756/B OR2X1_LOC_401/A 0.01fF
C18299 OR2X1_LOC_160/A OR2X1_LOC_864/A 0.03fF
C18300 AND2X1_LOC_392/A OR2X1_LOC_417/A 0.07fF
C18301 OR2X1_LOC_160/A OR2X1_LOC_469/a_36_216# 0.00fF
C18302 AND2X1_LOC_42/B OR2X1_LOC_575/A 0.00fF
C18303 AND2X1_LOC_862/a_8_24# AND2X1_LOC_807/Y 0.00fF
C18304 OR2X1_LOC_3/Y OR2X1_LOC_422/Y 0.00fF
C18305 OR2X1_LOC_475/Y OR2X1_LOC_721/Y 0.09fF
C18306 OR2X1_LOC_316/Y OR2X1_LOC_26/Y 0.04fF
C18307 OR2X1_LOC_476/B AND2X1_LOC_41/A 0.07fF
C18308 AND2X1_LOC_47/Y AND2X1_LOC_18/Y 1.11fF
C18309 OR2X1_LOC_31/Y OR2X1_LOC_583/Y 0.02fF
C18310 AND2X1_LOC_2/Y AND2X1_LOC_25/a_8_24# 0.18fF
C18311 OR2X1_LOC_102/a_8_216# OR2X1_LOC_47/Y 0.01fF
C18312 OR2X1_LOC_473/A OR2X1_LOC_361/a_8_216# 0.03fF
C18313 OR2X1_LOC_80/Y OR2X1_LOC_81/a_8_216# 0.18fF
C18314 AND2X1_LOC_364/Y OR2X1_LOC_22/Y 0.03fF
C18315 AND2X1_LOC_490/a_8_24# OR2X1_LOC_402/Y 0.03fF
C18316 OR2X1_LOC_600/A OR2X1_LOC_409/B 0.00fF
C18317 D_INPUT_5 AND2X1_LOC_21/a_8_24# 0.19fF
C18318 OR2X1_LOC_160/A OR2X1_LOC_633/B 0.14fF
C18319 OR2X1_LOC_743/A OR2X1_LOC_619/Y 0.10fF
C18320 VDD AND2X1_LOC_866/A 0.62fF
C18321 OR2X1_LOC_715/B OR2X1_LOC_112/B 0.14fF
C18322 AND2X1_LOC_857/Y AND2X1_LOC_863/A 0.06fF
C18323 AND2X1_LOC_81/B AND2X1_LOC_81/a_8_24# 0.11fF
C18324 OR2X1_LOC_379/a_8_216# AND2X1_LOC_3/Y 0.01fF
C18325 OR2X1_LOC_154/A OR2X1_LOC_219/B 0.04fF
C18326 OR2X1_LOC_237/Y OR2X1_LOC_238/Y 0.06fF
C18327 OR2X1_LOC_95/Y AND2X1_LOC_657/Y 0.27fF
C18328 OR2X1_LOC_574/A OR2X1_LOC_510/Y 0.34fF
C18329 OR2X1_LOC_699/a_36_216# OR2X1_LOC_43/A 0.01fF
C18330 AND2X1_LOC_395/a_8_24# OR2X1_LOC_287/B 0.00fF
C18331 AND2X1_LOC_56/B OR2X1_LOC_449/B 0.07fF
C18332 AND2X1_LOC_59/Y AND2X1_LOC_387/B 0.00fF
C18333 OR2X1_LOC_189/A AND2X1_LOC_474/Y 0.03fF
C18334 OR2X1_LOC_506/A AND2X1_LOC_69/Y 0.13fF
C18335 AND2X1_LOC_191/B OR2X1_LOC_95/Y 0.36fF
C18336 AND2X1_LOC_12/Y AND2X1_LOC_496/a_8_24# 0.01fF
C18337 OR2X1_LOC_9/Y AND2X1_LOC_721/A 0.18fF
C18338 AND2X1_LOC_555/Y OR2X1_LOC_384/a_36_216# 0.00fF
C18339 OR2X1_LOC_95/Y AND2X1_LOC_469/B 0.04fF
C18340 AND2X1_LOC_51/Y OR2X1_LOC_730/a_8_216# 0.00fF
C18341 OR2X1_LOC_426/A AND2X1_LOC_687/B 1.00fF
C18342 OR2X1_LOC_836/B OR2X1_LOC_269/B 0.00fF
C18343 AND2X1_LOC_366/A OR2X1_LOC_417/A 3.54fF
C18344 OR2X1_LOC_379/Y AND2X1_LOC_51/Y 0.04fF
C18345 OR2X1_LOC_185/A OR2X1_LOC_254/a_36_216# 0.00fF
C18346 OR2X1_LOC_495/Y AND2X1_LOC_465/Y 0.02fF
C18347 OR2X1_LOC_354/A D_INPUT_0 0.05fF
C18348 OR2X1_LOC_715/B OR2X1_LOC_66/Y 0.03fF
C18349 OR2X1_LOC_48/Y OR2X1_LOC_48/a_36_216# 0.00fF
C18350 OR2X1_LOC_682/a_8_216# OR2X1_LOC_7/A 0.04fF
C18351 OR2X1_LOC_837/B OR2X1_LOC_22/Y 0.03fF
C18352 OR2X1_LOC_280/Y OR2X1_LOC_372/Y 0.03fF
C18353 AND2X1_LOC_76/a_8_24# OR2X1_LOC_22/Y 0.04fF
C18354 OR2X1_LOC_119/a_8_216# OR2X1_LOC_39/A 0.01fF
C18355 AND2X1_LOC_733/Y AND2X1_LOC_440/a_8_24# 0.01fF
C18356 OR2X1_LOC_88/Y OR2X1_LOC_12/Y 0.00fF
C18357 AND2X1_LOC_580/B OR2X1_LOC_74/A 0.03fF
C18358 OR2X1_LOC_574/A OR2X1_LOC_810/A 0.19fF
C18359 OR2X1_LOC_158/A OR2X1_LOC_70/A 0.20fF
C18360 OR2X1_LOC_662/A OR2X1_LOC_476/B 0.01fF
C18361 OR2X1_LOC_246/A OR2X1_LOC_619/Y 0.01fF
C18362 OR2X1_LOC_12/Y OR2X1_LOC_172/Y 0.00fF
C18363 OR2X1_LOC_864/A OR2X1_LOC_624/B 0.07fF
C18364 AND2X1_LOC_578/A AND2X1_LOC_577/A 0.11fF
C18365 OR2X1_LOC_32/B OR2X1_LOC_19/B 0.01fF
C18366 OR2X1_LOC_628/Y AND2X1_LOC_621/Y 0.07fF
C18367 OR2X1_LOC_290/a_8_216# AND2X1_LOC_476/A 0.04fF
C18368 OR2X1_LOC_16/A OR2X1_LOC_80/A 5.77fF
C18369 AND2X1_LOC_371/a_36_24# OR2X1_LOC_493/Y 0.00fF
C18370 AND2X1_LOC_18/Y OR2X1_LOC_598/A 0.14fF
C18371 OR2X1_LOC_481/A AND2X1_LOC_818/a_8_24# 0.01fF
C18372 OR2X1_LOC_502/A OR2X1_LOC_218/Y 0.03fF
C18373 OR2X1_LOC_114/Y AND2X1_LOC_51/Y 0.03fF
C18374 AND2X1_LOC_95/Y OR2X1_LOC_720/B 0.02fF
C18375 AND2X1_LOC_486/Y AND2X1_LOC_227/Y 0.03fF
C18376 AND2X1_LOC_619/a_8_24# OR2X1_LOC_622/B 0.01fF
C18377 OR2X1_LOC_3/Y AND2X1_LOC_259/Y 0.06fF
C18378 OR2X1_LOC_131/Y OR2X1_LOC_7/A 0.03fF
C18379 OR2X1_LOC_808/A OR2X1_LOC_223/A 0.20fF
C18380 AND2X1_LOC_18/a_8_24# AND2X1_LOC_3/Y 0.03fF
C18381 INPUT_1 AND2X1_LOC_847/Y 0.03fF
C18382 AND2X1_LOC_56/B OR2X1_LOC_121/B 0.10fF
C18383 OR2X1_LOC_471/Y OR2X1_LOC_738/A 0.07fF
C18384 AND2X1_LOC_51/a_8_24# OR2X1_LOC_51/B 0.01fF
C18385 OR2X1_LOC_431/Y OR2X1_LOC_26/Y 0.18fF
C18386 OR2X1_LOC_665/Y AND2X1_LOC_483/a_36_24# 0.01fF
C18387 OR2X1_LOC_632/Y OR2X1_LOC_493/Y 0.10fF
C18388 AND2X1_LOC_68/a_8_24# OR2X1_LOC_69/A 0.01fF
C18389 AND2X1_LOC_92/Y OR2X1_LOC_365/B 0.03fF
C18390 AND2X1_LOC_8/Y OR2X1_LOC_121/B 0.46fF
C18391 AND2X1_LOC_729/Y AND2X1_LOC_801/B 0.01fF
C18392 AND2X1_LOC_101/a_8_24# OR2X1_LOC_26/Y 0.06fF
C18393 OR2X1_LOC_135/Y OR2X1_LOC_437/A 0.10fF
C18394 AND2X1_LOC_44/Y AND2X1_LOC_41/Y 0.02fF
C18395 OR2X1_LOC_160/B OR2X1_LOC_560/A 0.04fF
C18396 OR2X1_LOC_421/Y OR2X1_LOC_423/Y 0.05fF
C18397 OR2X1_LOC_168/Y OR2X1_LOC_390/B 0.71fF
C18398 OR2X1_LOC_218/Y AND2X1_LOC_230/a_8_24# 0.17fF
C18399 OR2X1_LOC_168/B OR2X1_LOC_318/B 0.00fF
C18400 D_INPUT_4 OR2X1_LOC_2/a_8_216# 0.02fF
C18401 OR2X1_LOC_500/A AND2X1_LOC_47/Y 0.06fF
C18402 OR2X1_LOC_315/Y AND2X1_LOC_866/A 1.75fF
C18403 AND2X1_LOC_831/Y AND2X1_LOC_138/a_36_24# 0.02fF
C18404 OR2X1_LOC_616/Y AND2X1_LOC_866/A 0.03fF
C18405 OR2X1_LOC_864/A OR2X1_LOC_655/A 0.01fF
C18406 AND2X1_LOC_841/a_36_24# AND2X1_LOC_662/B 0.01fF
C18407 AND2X1_LOC_851/B OR2X1_LOC_39/A 0.09fF
C18408 AND2X1_LOC_86/Y OR2X1_LOC_84/a_8_216# 0.03fF
C18409 OR2X1_LOC_244/A OR2X1_LOC_267/A 0.12fF
C18410 OR2X1_LOC_273/a_8_216# OR2X1_LOC_416/Y 0.01fF
C18411 OR2X1_LOC_19/B AND2X1_LOC_4/a_8_24# 0.14fF
C18412 OR2X1_LOC_338/B OR2X1_LOC_338/A 0.06fF
C18413 OR2X1_LOC_844/Y AND2X1_LOC_51/Y 0.13fF
C18414 OR2X1_LOC_485/A AND2X1_LOC_196/Y 0.15fF
C18415 AND2X1_LOC_37/a_8_24# INPUT_1 0.01fF
C18416 AND2X1_LOC_47/Y AND2X1_LOC_234/a_8_24# 0.01fF
C18417 OR2X1_LOC_251/Y AND2X1_LOC_866/A 0.07fF
C18418 AND2X1_LOC_754/a_8_24# AND2X1_LOC_36/Y 0.01fF
C18419 OR2X1_LOC_160/A OR2X1_LOC_215/a_36_216# 0.01fF
C18420 OR2X1_LOC_244/A OR2X1_LOC_204/a_36_216# 0.00fF
C18421 OR2X1_LOC_617/Y AND2X1_LOC_621/a_36_24# 0.00fF
C18422 OR2X1_LOC_306/Y OR2X1_LOC_599/Y 0.02fF
C18423 OR2X1_LOC_844/Y OR2X1_LOC_849/a_8_216# 0.02fF
C18424 AND2X1_LOC_723/a_8_24# AND2X1_LOC_222/Y 0.01fF
C18425 OR2X1_LOC_56/A OR2X1_LOC_13/B 0.33fF
C18426 OR2X1_LOC_6/A OR2X1_LOC_29/a_8_216# 0.03fF
C18427 OR2X1_LOC_3/B OR2X1_LOC_44/Y 0.01fF
C18428 OR2X1_LOC_595/Y OR2X1_LOC_39/A 0.05fF
C18429 OR2X1_LOC_291/Y OR2X1_LOC_62/B 0.01fF
C18430 AND2X1_LOC_67/Y OR2X1_LOC_532/B 0.02fF
C18431 AND2X1_LOC_64/Y OR2X1_LOC_580/B 0.05fF
C18432 AND2X1_LOC_662/B AND2X1_LOC_222/Y 0.03fF
C18433 OR2X1_LOC_500/A OR2X1_LOC_598/A 0.00fF
C18434 AND2X1_LOC_59/Y OR2X1_LOC_318/B 0.04fF
C18435 AND2X1_LOC_213/B AND2X1_LOC_213/a_8_24# 0.00fF
C18436 AND2X1_LOC_476/Y AND2X1_LOC_439/a_36_24# 0.00fF
C18437 OR2X1_LOC_244/Y OR2X1_LOC_342/B 0.01fF
C18438 AND2X1_LOC_383/a_36_24# OR2X1_LOC_428/A 0.02fF
C18439 OR2X1_LOC_232/a_8_216# D_INPUT_1 0.01fF
C18440 AND2X1_LOC_22/Y AND2X1_LOC_44/Y 0.21fF
C18441 OR2X1_LOC_35/A OR2X1_LOC_338/A 0.02fF
C18442 AND2X1_LOC_866/A AND2X1_LOC_624/a_8_24# 0.02fF
C18443 OR2X1_LOC_521/Y OR2X1_LOC_521/a_8_216# -0.00fF
C18444 AND2X1_LOC_413/a_8_24# OR2X1_LOC_598/A 0.01fF
C18445 AND2X1_LOC_59/Y OR2X1_LOC_854/A 0.04fF
C18446 OR2X1_LOC_18/Y AND2X1_LOC_216/a_8_24# 0.04fF
C18447 OR2X1_LOC_696/A OR2X1_LOC_96/Y 0.04fF
C18448 AND2X1_LOC_48/A AND2X1_LOC_692/a_36_24# 0.01fF
C18449 OR2X1_LOC_88/a_36_216# OR2X1_LOC_39/A 0.00fF
C18450 OR2X1_LOC_235/B OR2X1_LOC_771/B 0.07fF
C18451 AND2X1_LOC_773/Y AND2X1_LOC_774/a_8_24# 0.11fF
C18452 OR2X1_LOC_856/B OR2X1_LOC_446/B 1.17fF
C18453 OR2X1_LOC_522/Y OR2X1_LOC_428/A 0.01fF
C18454 OR2X1_LOC_612/B AND2X1_LOC_647/Y 0.17fF
C18455 AND2X1_LOC_741/Y AND2X1_LOC_742/a_8_24# 0.11fF
C18456 AND2X1_LOC_699/a_8_24# AND2X1_LOC_3/Y 0.01fF
C18457 OR2X1_LOC_22/A OR2X1_LOC_409/B 0.00fF
C18458 OR2X1_LOC_162/Y OR2X1_LOC_161/B 0.01fF
C18459 OR2X1_LOC_199/a_8_216# OR2X1_LOC_790/A 0.47fF
C18460 AND2X1_LOC_650/Y OR2X1_LOC_172/Y 0.00fF
C18461 OR2X1_LOC_111/a_8_216# OR2X1_LOC_56/A 0.02fF
C18462 OR2X1_LOC_527/a_36_216# AND2X1_LOC_721/Y 0.00fF
C18463 AND2X1_LOC_850/Y OR2X1_LOC_13/B 0.01fF
C18464 AND2X1_LOC_3/Y OR2X1_LOC_675/Y 0.20fF
C18465 D_INPUT_3 OR2X1_LOC_62/B 0.03fF
C18466 AND2X1_LOC_660/A OR2X1_LOC_46/A 0.03fF
C18467 OR2X1_LOC_549/B OR2X1_LOC_563/a_8_216# 0.49fF
C18468 OR2X1_LOC_538/A OR2X1_LOC_356/B 0.09fF
C18469 OR2X1_LOC_421/A OR2X1_LOC_764/a_36_216# 0.00fF
C18470 OR2X1_LOC_502/A OR2X1_LOC_703/Y 0.03fF
C18471 AND2X1_LOC_624/B AND2X1_LOC_624/a_36_24# 0.01fF
C18472 AND2X1_LOC_724/a_8_24# AND2X1_LOC_447/Y 0.04fF
C18473 AND2X1_LOC_863/Y AND2X1_LOC_864/a_8_24# 0.04fF
C18474 AND2X1_LOC_848/Y OR2X1_LOC_437/A 5.95fF
C18475 OR2X1_LOC_45/B AND2X1_LOC_732/B 0.01fF
C18476 AND2X1_LOC_1/Y OR2X1_LOC_451/B 0.07fF
C18477 AND2X1_LOC_186/a_8_24# OR2X1_LOC_437/A 0.04fF
C18478 OR2X1_LOC_46/A AND2X1_LOC_646/a_8_24# 0.03fF
C18479 OR2X1_LOC_7/A AND2X1_LOC_657/A 0.13fF
C18480 AND2X1_LOC_645/A OR2X1_LOC_534/Y 0.01fF
C18481 AND2X1_LOC_672/a_8_24# AND2X1_LOC_47/Y 0.02fF
C18482 OR2X1_LOC_516/Y OR2X1_LOC_495/Y 0.03fF
C18483 D_GATE_479 OR2X1_LOC_466/A 0.00fF
C18484 AND2X1_LOC_810/A AND2X1_LOC_567/a_8_24# 0.01fF
C18485 AND2X1_LOC_745/a_8_24# OR2X1_LOC_781/B 0.01fF
C18486 OR2X1_LOC_421/A AND2X1_LOC_706/Y 0.08fF
C18487 OR2X1_LOC_223/A OR2X1_LOC_223/a_8_216# 0.18fF
C18488 OR2X1_LOC_337/A VDD 0.06fF
C18489 AND2X1_LOC_542/a_36_24# AND2X1_LOC_476/Y -0.02fF
C18490 AND2X1_LOC_721/Y OR2X1_LOC_59/Y 0.08fF
C18491 OR2X1_LOC_466/A OR2X1_LOC_161/B 0.51fF
C18492 AND2X1_LOC_131/a_8_24# OR2X1_LOC_549/A 0.03fF
C18493 OR2X1_LOC_244/A OR2X1_LOC_84/a_8_216# 0.04fF
C18494 OR2X1_LOC_6/B AND2X1_LOC_275/a_8_24# 0.04fF
C18495 AND2X1_LOC_521/a_8_24# AND2X1_LOC_18/Y 0.05fF
C18496 OR2X1_LOC_364/A OR2X1_LOC_777/B 0.07fF
C18497 OR2X1_LOC_620/Y OR2X1_LOC_354/a_8_216# 0.01fF
C18498 AND2X1_LOC_551/a_8_24# AND2X1_LOC_551/B 0.19fF
C18499 AND2X1_LOC_338/A OR2X1_LOC_51/Y 0.01fF
C18500 AND2X1_LOC_658/B AND2X1_LOC_469/a_8_24# 0.03fF
C18501 OR2X1_LOC_338/a_8_216# VDD 0.21fF
C18502 OR2X1_LOC_756/B AND2X1_LOC_7/B 0.28fF
C18503 OR2X1_LOC_188/Y OR2X1_LOC_499/B 0.00fF
C18504 OR2X1_LOC_604/A OR2X1_LOC_382/a_8_216# 0.04fF
C18505 OR2X1_LOC_235/B OR2X1_LOC_721/a_36_216# 0.00fF
C18506 OR2X1_LOC_106/Y OR2X1_LOC_521/Y 0.18fF
C18507 OR2X1_LOC_706/A AND2X1_LOC_44/Y 0.01fF
C18508 OR2X1_LOC_160/A OR2X1_LOC_501/A 0.03fF
C18509 OR2X1_LOC_40/Y VDD 2.02fF
C18510 OR2X1_LOC_336/a_8_216# OR2X1_LOC_703/A 0.01fF
C18511 OR2X1_LOC_369/Y OR2X1_LOC_322/Y 0.06fF
C18512 AND2X1_LOC_866/A AND2X1_LOC_624/B 0.02fF
C18513 OR2X1_LOC_468/Y AND2X1_LOC_36/Y 0.00fF
C18514 OR2X1_LOC_36/Y OR2X1_LOC_268/Y 0.60fF
C18515 OR2X1_LOC_92/a_36_216# OR2X1_LOC_67/Y 0.01fF
C18516 OR2X1_LOC_19/B OR2X1_LOC_68/B 1.64fF
C18517 OR2X1_LOC_654/a_8_216# OR2X1_LOC_78/B 0.01fF
C18518 OR2X1_LOC_36/Y OR2X1_LOC_183/Y 0.01fF
C18519 AND2X1_LOC_64/Y OR2X1_LOC_507/B 0.40fF
C18520 OR2X1_LOC_223/A OR2X1_LOC_795/a_8_216# 0.01fF
C18521 AND2X1_LOC_42/B OR2X1_LOC_735/B 0.00fF
C18522 OR2X1_LOC_482/Y OR2X1_LOC_59/Y 0.29fF
C18523 OR2X1_LOC_830/a_8_216# OR2X1_LOC_190/A 0.01fF
C18524 OR2X1_LOC_114/B AND2X1_LOC_184/a_36_24# 0.00fF
C18525 OR2X1_LOC_51/a_8_216# OR2X1_LOC_51/B 0.07fF
C18526 AND2X1_LOC_70/Y OR2X1_LOC_832/a_8_216# 0.01fF
C18527 OR2X1_LOC_49/A OR2X1_LOC_502/A 8.26fF
C18528 OR2X1_LOC_44/Y OR2X1_LOC_759/Y 0.22fF
C18529 VDD AND2X1_LOC_172/a_8_24# -0.00fF
C18530 OR2X1_LOC_710/A OR2X1_LOC_375/A 0.00fF
C18531 VDD AND2X1_LOC_535/a_8_24# 0.00fF
C18532 OR2X1_LOC_854/a_8_216# OR2X1_LOC_161/B 0.01fF
C18533 AND2X1_LOC_477/A OR2X1_LOC_534/Y 0.03fF
C18534 OR2X1_LOC_223/A OR2X1_LOC_374/Y 0.03fF
C18535 AND2X1_LOC_130/a_8_24# AND2X1_LOC_139/a_8_24# 0.23fF
C18536 D_INPUT_7 INPUT_6 0.61fF
C18537 AND2X1_LOC_728/Y AND2X1_LOC_564/A 0.03fF
C18538 OR2X1_LOC_51/Y OR2X1_LOC_411/a_36_216# 0.00fF
C18539 AND2X1_LOC_40/Y OR2X1_LOC_549/A 0.08fF
C18540 OR2X1_LOC_805/A OR2X1_LOC_362/a_8_216# 0.02fF
C18541 AND2X1_LOC_76/Y OR2X1_LOC_12/Y 0.03fF
C18542 OR2X1_LOC_502/A OR2X1_LOC_596/A 0.04fF
C18543 OR2X1_LOC_185/Y OR2X1_LOC_831/B 0.04fF
C18544 OR2X1_LOC_506/a_36_216# OR2X1_LOC_185/Y 0.15fF
C18545 AND2X1_LOC_160/Y AND2X1_LOC_162/a_8_24# 0.09fF
C18546 OR2X1_LOC_479/Y OR2X1_LOC_301/a_8_216# 0.01fF
C18547 AND2X1_LOC_576/Y OR2X1_LOC_184/a_8_216# 0.01fF
C18548 OR2X1_LOC_158/A AND2X1_LOC_357/a_8_24# 0.01fF
C18549 OR2X1_LOC_829/A OR2X1_LOC_48/B 0.02fF
C18550 OR2X1_LOC_354/A OR2X1_LOC_356/a_8_216# 0.03fF
C18551 AND2X1_LOC_574/Y OR2X1_LOC_498/Y 0.06fF
C18552 AND2X1_LOC_794/A AND2X1_LOC_794/B 0.11fF
C18553 OR2X1_LOC_294/Y AND2X1_LOC_297/a_8_24# 0.01fF
C18554 OR2X1_LOC_65/B AND2X1_LOC_249/a_8_24# -0.00fF
C18555 OR2X1_LOC_18/Y OR2X1_LOC_829/A 0.01fF
C18556 OR2X1_LOC_67/A OR2X1_LOC_12/Y 0.03fF
C18557 OR2X1_LOC_76/Y AND2X1_LOC_7/B 0.15fF
C18558 OR2X1_LOC_549/a_8_216# OR2X1_LOC_563/B 0.14fF
C18559 AND2X1_LOC_70/Y OR2X1_LOC_474/Y 0.03fF
C18560 OR2X1_LOC_151/A AND2X1_LOC_314/a_36_24# 0.01fF
C18561 OR2X1_LOC_156/B OR2X1_LOC_87/A 0.02fF
C18562 OR2X1_LOC_95/Y OR2X1_LOC_164/a_8_216# 0.02fF
C18563 OR2X1_LOC_323/A OR2X1_LOC_371/Y 0.02fF
C18564 AND2X1_LOC_753/B OR2X1_LOC_66/A 0.07fF
C18565 OR2X1_LOC_154/A OR2X1_LOC_691/B 0.01fF
C18566 OR2X1_LOC_318/Y OR2X1_LOC_776/Y 0.73fF
C18567 AND2X1_LOC_377/Y AND2X1_LOC_378/a_8_24# 0.00fF
C18568 OR2X1_LOC_539/A AND2X1_LOC_70/Y 0.01fF
C18569 AND2X1_LOC_861/a_8_24# AND2X1_LOC_865/a_8_24# 0.23fF
C18570 AND2X1_LOC_865/A AND2X1_LOC_862/Y 0.02fF
C18571 OR2X1_LOC_6/A OR2X1_LOC_16/A 5.46fF
C18572 OR2X1_LOC_118/Y OR2X1_LOC_131/a_8_216# 0.01fF
C18573 OR2X1_LOC_696/A OR2X1_LOC_829/Y 0.02fF
C18574 OR2X1_LOC_347/a_8_216# OR2X1_LOC_66/A 0.08fF
C18575 VDD AND2X1_LOC_843/Y 0.01fF
C18576 OR2X1_LOC_351/B AND2X1_LOC_59/Y 0.07fF
C18577 AND2X1_LOC_781/a_8_24# AND2X1_LOC_781/Y 0.01fF
C18578 AND2X1_LOC_39/a_8_24# OR2X1_LOC_78/B 0.02fF
C18579 AND2X1_LOC_705/Y OR2X1_LOC_36/Y 0.10fF
C18580 OR2X1_LOC_508/a_8_216# OR2X1_LOC_87/A 0.03fF
C18581 AND2X1_LOC_12/Y OR2X1_LOC_182/B 0.03fF
C18582 AND2X1_LOC_794/A VDD 0.25fF
C18583 OR2X1_LOC_76/A OR2X1_LOC_605/Y 0.01fF
C18584 OR2X1_LOC_329/Y AND2X1_LOC_436/B 0.02fF
C18585 AND2X1_LOC_571/a_8_24# OR2X1_LOC_89/A 0.01fF
C18586 OR2X1_LOC_87/A OR2X1_LOC_486/Y 0.32fF
C18587 OR2X1_LOC_506/A AND2X1_LOC_18/Y 0.00fF
C18588 OR2X1_LOC_471/Y AND2X1_LOC_36/Y 3.66fF
C18589 OR2X1_LOC_623/B OR2X1_LOC_715/A 0.04fF
C18590 AND2X1_LOC_193/a_8_24# OR2X1_LOC_13/Y 0.01fF
C18591 OR2X1_LOC_458/B OR2X1_LOC_458/a_8_216# 0.13fF
C18592 OR2X1_LOC_40/Y OR2X1_LOC_616/Y 0.44fF
C18593 OR2X1_LOC_405/A OR2X1_LOC_66/A 0.10fF
C18594 AND2X1_LOC_713/a_8_24# OR2X1_LOC_599/A 0.00fF
C18595 OR2X1_LOC_12/Y OR2X1_LOC_52/B 0.58fF
C18596 OR2X1_LOC_840/A AND2X1_LOC_167/a_8_24# 0.12fF
C18597 OR2X1_LOC_114/B AND2X1_LOC_59/Y 0.02fF
C18598 AND2X1_LOC_508/B AND2X1_LOC_621/Y 0.03fF
C18599 OR2X1_LOC_517/A AND2X1_LOC_139/a_8_24# 0.03fF
C18600 OR2X1_LOC_766/Y OR2X1_LOC_52/B 0.03fF
C18601 OR2X1_LOC_299/a_8_216# OR2X1_LOC_16/A 0.06fF
C18602 OR2X1_LOC_261/a_36_216# AND2X1_LOC_847/Y 0.00fF
C18603 AND2X1_LOC_721/Y OR2X1_LOC_70/Y 0.03fF
C18604 OR2X1_LOC_691/A OR2X1_LOC_654/A 0.03fF
C18605 VDD OR2X1_LOC_539/Y 0.27fF
C18606 AND2X1_LOC_555/a_8_24# OR2X1_LOC_44/Y 0.01fF
C18607 AND2X1_LOC_549/Y AND2X1_LOC_580/A 0.01fF
C18608 AND2X1_LOC_489/Y OR2X1_LOC_12/Y 0.00fF
C18609 AND2X1_LOC_658/A AND2X1_LOC_862/A 0.00fF
C18610 AND2X1_LOC_539/Y AND2X1_LOC_802/a_8_24# 0.01fF
C18611 AND2X1_LOC_658/A AND2X1_LOC_624/A 0.10fF
C18612 AND2X1_LOC_84/Y OR2X1_LOC_291/Y 0.03fF
C18613 OR2X1_LOC_116/A AND2X1_LOC_70/Y 0.01fF
C18614 OR2X1_LOC_318/Y OR2X1_LOC_756/B 0.03fF
C18615 OR2X1_LOC_40/Y AND2X1_LOC_267/a_8_24# 0.00fF
C18616 OR2X1_LOC_363/B OR2X1_LOC_805/A 0.03fF
C18617 OR2X1_LOC_467/A OR2X1_LOC_448/Y 0.00fF
C18618 AND2X1_LOC_42/B OR2X1_LOC_161/B 0.05fF
C18619 AND2X1_LOC_3/Y OR2X1_LOC_736/Y 0.01fF
C18620 OR2X1_LOC_385/Y OR2X1_LOC_829/A 0.06fF
C18621 AND2X1_LOC_535/Y OR2X1_LOC_44/Y 0.03fF
C18622 OR2X1_LOC_203/Y AND2X1_LOC_625/a_36_24# 0.00fF
C18623 VDD OR2X1_LOC_618/a_8_216# 0.21fF
C18624 AND2X1_LOC_752/a_8_24# D_INPUT_5 0.01fF
C18625 AND2X1_LOC_367/A OR2X1_LOC_278/Y 0.05fF
C18626 OR2X1_LOC_614/Y AND2X1_LOC_3/Y 0.01fF
C18627 OR2X1_LOC_630/Y OR2X1_LOC_499/a_8_216# 0.01fF
C18628 AND2X1_LOC_83/a_8_24# OR2X1_LOC_557/A 0.00fF
C18629 OR2X1_LOC_91/A OR2X1_LOC_118/Y 0.03fF
C18630 AND2X1_LOC_388/Y AND2X1_LOC_645/A 0.09fF
C18631 AND2X1_LOC_500/Y AND2X1_LOC_580/A 0.03fF
C18632 OR2X1_LOC_91/Y OR2X1_LOC_666/A 0.02fF
C18633 AND2X1_LOC_43/B OR2X1_LOC_78/B 0.11fF
C18634 AND2X1_LOC_736/Y AND2X1_LOC_737/Y 0.05fF
C18635 OR2X1_LOC_217/Y AND2X1_LOC_70/Y 0.01fF
C18636 OR2X1_LOC_715/B OR2X1_LOC_574/A 0.01fF
C18637 AND2X1_LOC_344/a_36_24# OR2X1_LOC_92/Y 0.00fF
C18638 AND2X1_LOC_714/B OR2X1_LOC_3/Y 0.07fF
C18639 AND2X1_LOC_724/Y OR2X1_LOC_601/Y 0.01fF
C18640 AND2X1_LOC_663/B OR2X1_LOC_759/a_36_216# 0.00fF
C18641 OR2X1_LOC_298/a_8_216# OR2X1_LOC_619/Y 0.02fF
C18642 AND2X1_LOC_59/Y OR2X1_LOC_538/A 0.02fF
C18643 OR2X1_LOC_674/a_8_216# OR2X1_LOC_39/A 0.06fF
C18644 AND2X1_LOC_501/a_8_24# AND2X1_LOC_576/Y 0.03fF
C18645 OR2X1_LOC_106/a_8_216# OR2X1_LOC_3/Y -0.00fF
C18646 OR2X1_LOC_597/A OR2X1_LOC_585/A 0.00fF
C18647 AND2X1_LOC_859/a_36_24# OR2X1_LOC_59/Y 0.00fF
C18648 OR2X1_LOC_502/A OR2X1_LOC_732/a_8_216# 0.02fF
C18649 OR2X1_LOC_280/Y AND2X1_LOC_243/Y 0.02fF
C18650 OR2X1_LOC_756/B OR2X1_LOC_805/A 0.06fF
C18651 AND2X1_LOC_598/a_8_24# OR2X1_LOC_744/A 0.04fF
C18652 OR2X1_LOC_421/A OR2X1_LOC_485/A 0.03fF
C18653 OR2X1_LOC_43/A AND2X1_LOC_691/a_8_24# 0.01fF
C18654 OR2X1_LOC_458/B AND2X1_LOC_272/a_8_24# 0.20fF
C18655 OR2X1_LOC_40/Y AND2X1_LOC_389/a_8_24# 0.03fF
C18656 OR2X1_LOC_70/Y OR2X1_LOC_482/Y 0.00fF
C18657 VDD OR2X1_LOC_7/A 0.91fF
C18658 AND2X1_LOC_465/a_8_24# OR2X1_LOC_108/Y 0.04fF
C18659 OR2X1_LOC_748/A OR2X1_LOC_59/Y 0.02fF
C18660 OR2X1_LOC_624/A OR2X1_LOC_436/B 0.08fF
C18661 AND2X1_LOC_773/Y OR2X1_LOC_22/Y 0.12fF
C18662 OR2X1_LOC_49/A AND2X1_LOC_48/A 0.00fF
C18663 AND2X1_LOC_22/Y OR2X1_LOC_720/B 0.01fF
C18664 OR2X1_LOC_523/Y OR2X1_LOC_560/a_8_216# 0.08fF
C18665 OR2X1_LOC_479/Y AND2X1_LOC_110/Y 0.03fF
C18666 OR2X1_LOC_841/B OR2X1_LOC_168/B 0.03fF
C18667 OR2X1_LOC_744/A OR2X1_LOC_26/Y 3.43fF
C18668 OR2X1_LOC_803/a_8_216# OR2X1_LOC_87/A 0.01fF
C18669 AND2X1_LOC_41/A OR2X1_LOC_264/a_8_216# 0.09fF
C18670 AND2X1_LOC_208/a_36_24# AND2X1_LOC_35/Y 0.00fF
C18671 OR2X1_LOC_109/Y OR2X1_LOC_427/A 0.02fF
C18672 OR2X1_LOC_317/a_8_216# AND2X1_LOC_56/B 0.03fF
C18673 VDD OR2X1_LOC_320/Y 0.04fF
C18674 OR2X1_LOC_404/Y OR2X1_LOC_362/A 0.07fF
C18675 OR2X1_LOC_502/A OR2X1_LOC_463/B 0.08fF
C18676 OR2X1_LOC_744/A AND2X1_LOC_493/a_8_24# 0.01fF
C18677 AND2X1_LOC_724/A OR2X1_LOC_601/a_8_216# 0.03fF
C18678 OR2X1_LOC_323/A AND2X1_LOC_841/a_36_24# -0.00fF
C18679 OR2X1_LOC_91/Y AND2X1_LOC_716/Y 0.01fF
C18680 OR2X1_LOC_448/Y OR2X1_LOC_725/B 0.01fF
C18681 VDD AND2X1_LOC_176/a_8_24# 0.00fF
C18682 OR2X1_LOC_837/B OR2X1_LOC_39/A 0.03fF
C18683 AND2X1_LOC_497/a_8_24# OR2X1_LOC_844/B 0.01fF
C18684 AND2X1_LOC_349/B OR2X1_LOC_744/A 0.06fF
C18685 OR2X1_LOC_427/A AND2X1_LOC_448/Y 0.03fF
C18686 AND2X1_LOC_858/B OR2X1_LOC_238/Y 0.01fF
C18687 AND2X1_LOC_76/a_8_24# OR2X1_LOC_39/A 0.03fF
C18688 AND2X1_LOC_838/Y AND2X1_LOC_852/B 0.26fF
C18689 AND2X1_LOC_729/Y AND2X1_LOC_703/a_8_24# 0.03fF
C18690 OR2X1_LOC_744/A OR2X1_LOC_89/A 0.13fF
C18691 OR2X1_LOC_160/A OR2X1_LOC_784/Y 0.03fF
C18692 AND2X1_LOC_364/Y AND2X1_LOC_211/B 0.00fF
C18693 OR2X1_LOC_48/B AND2X1_LOC_648/a_8_24# 0.04fF
C18694 AND2X1_LOC_48/A OR2X1_LOC_596/A 0.03fF
C18695 OR2X1_LOC_116/a_8_216# OR2X1_LOC_474/Y 0.05fF
C18696 OR2X1_LOC_777/B OR2X1_LOC_568/A 0.07fF
C18697 OR2X1_LOC_290/a_8_216# OR2X1_LOC_690/A 0.01fF
C18698 OR2X1_LOC_264/Y OR2X1_LOC_264/a_36_216# 0.00fF
C18699 OR2X1_LOC_118/Y AND2X1_LOC_573/A 0.04fF
C18700 OR2X1_LOC_161/A OR2X1_LOC_541/B 0.02fF
C18701 OR2X1_LOC_409/B AND2X1_LOC_769/Y 0.01fF
C18702 OR2X1_LOC_18/Y AND2X1_LOC_648/a_8_24# 0.02fF
C18703 OR2X1_LOC_473/A OR2X1_LOC_267/Y 0.04fF
C18704 OR2X1_LOC_223/A OR2X1_LOC_392/B 0.12fF
C18705 OR2X1_LOC_256/Y OR2X1_LOC_585/A 0.13fF
C18706 AND2X1_LOC_566/B AND2X1_LOC_326/a_36_24# 0.00fF
C18707 AND2X1_LOC_214/A OR2X1_LOC_3/Y 0.02fF
C18708 OR2X1_LOC_160/A OR2X1_LOC_738/A 0.05fF
C18709 OR2X1_LOC_22/Y AND2X1_LOC_243/Y 0.09fF
C18710 AND2X1_LOC_12/Y AND2X1_LOC_59/Y 0.39fF
C18711 OR2X1_LOC_304/Y OR2X1_LOC_59/Y 0.21fF
C18712 OR2X1_LOC_422/a_8_216# OR2X1_LOC_52/B 0.03fF
C18713 AND2X1_LOC_456/B OR2X1_LOC_485/A 0.06fF
C18714 AND2X1_LOC_50/Y OR2X1_LOC_651/a_36_216# 0.00fF
C18715 AND2X1_LOC_753/B OR2X1_LOC_651/a_8_216# 0.01fF
C18716 OR2X1_LOC_305/Y AND2X1_LOC_654/Y 0.04fF
C18717 OR2X1_LOC_185/Y OR2X1_LOC_493/A 0.14fF
C18718 AND2X1_LOC_36/Y OR2X1_LOC_750/Y 0.00fF
C18719 OR2X1_LOC_502/A AND2X1_LOC_612/B 0.40fF
C18720 OR2X1_LOC_375/A AND2X1_LOC_43/B 0.54fF
C18721 OR2X1_LOC_91/A AND2X1_LOC_211/a_36_24# 0.00fF
C18722 OR2X1_LOC_69/Y OR2X1_LOC_393/a_36_216# 0.00fF
C18723 OR2X1_LOC_358/a_8_216# OR2X1_LOC_405/Y 0.40fF
C18724 OR2X1_LOC_231/a_8_216# OR2X1_LOC_87/A 0.02fF
C18725 OR2X1_LOC_863/B AND2X1_LOC_41/A 0.09fF
C18726 AND2X1_LOC_663/B AND2X1_LOC_663/A 0.00fF
C18727 AND2X1_LOC_319/a_8_24# AND2X1_LOC_802/Y 0.01fF
C18728 AND2X1_LOC_318/Y AND2X1_LOC_810/B 0.00fF
C18729 OR2X1_LOC_476/B OR2X1_LOC_648/A 0.02fF
C18730 OR2X1_LOC_600/A AND2X1_LOC_814/a_36_24# 0.00fF
C18731 AND2X1_LOC_12/Y OR2X1_LOC_865/a_8_216# 0.01fF
C18732 OR2X1_LOC_121/B AND2X1_LOC_92/Y 0.10fF
C18733 AND2X1_LOC_784/A AND2X1_LOC_468/B 0.12fF
C18734 OR2X1_LOC_654/A OR2X1_LOC_637/a_8_216# 0.02fF
C18735 AND2X1_LOC_566/B AND2X1_LOC_170/B 0.00fF
C18736 OR2X1_LOC_69/a_8_216# OR2X1_LOC_39/A 0.03fF
C18737 INPUT_0 OR2X1_LOC_43/a_8_216# 0.01fF
C18738 AND2X1_LOC_47/Y OR2X1_LOC_307/A 0.00fF
C18739 OR2X1_LOC_643/A OR2X1_LOC_624/A 0.00fF
C18740 OR2X1_LOC_31/Y OR2X1_LOC_765/Y 0.00fF
C18741 AND2X1_LOC_42/B AND2X1_LOC_618/a_8_24# 0.01fF
C18742 OR2X1_LOC_510/Y OR2X1_LOC_203/Y 0.18fF
C18743 AND2X1_LOC_59/Y OR2X1_LOC_841/B 0.01fF
C18744 OR2X1_LOC_116/A OR2X1_LOC_116/a_8_216# 0.39fF
C18745 OR2X1_LOC_756/B OR2X1_LOC_436/a_8_216# 0.01fF
C18746 OR2X1_LOC_262/Y AND2X1_LOC_573/A 0.02fF
C18747 OR2X1_LOC_628/Y OR2X1_LOC_59/Y 0.07fF
C18748 OR2X1_LOC_47/Y AND2X1_LOC_469/a_8_24# 0.18fF
C18749 AND2X1_LOC_723/a_8_24# OR2X1_LOC_74/A 0.12fF
C18750 OR2X1_LOC_36/Y OR2X1_LOC_511/Y 0.16fF
C18751 OR2X1_LOC_270/Y OR2X1_LOC_736/Y 0.03fF
C18752 AND2X1_LOC_537/Y INPUT_0 0.03fF
C18753 AND2X1_LOC_12/Y AND2X1_LOC_495/a_8_24# 0.02fF
C18754 OR2X1_LOC_404/Y OR2X1_LOC_474/Y 0.05fF
C18755 AND2X1_LOC_848/Y OR2X1_LOC_753/A 0.07fF
C18756 OR2X1_LOC_694/a_8_216# OR2X1_LOC_52/B 0.02fF
C18757 OR2X1_LOC_74/A OR2X1_LOC_278/Y 0.89fF
C18758 AND2X1_LOC_570/Y OR2X1_LOC_71/Y 0.02fF
C18759 OR2X1_LOC_158/A OR2X1_LOC_47/Y 0.14fF
C18760 OR2X1_LOC_70/Y OR2X1_LOC_586/Y 0.09fF
C18761 OR2X1_LOC_185/A OR2X1_LOC_220/a_8_216# 0.06fF
C18762 AND2X1_LOC_76/Y OR2X1_LOC_272/Y 0.00fF
C18763 OR2X1_LOC_315/Y OR2X1_LOC_7/A 0.49fF
C18764 AND2X1_LOC_662/B OR2X1_LOC_74/A 0.16fF
C18765 OR2X1_LOC_125/a_36_216# OR2X1_LOC_95/Y 0.03fF
C18766 OR2X1_LOC_377/A AND2X1_LOC_459/a_8_24# 0.08fF
C18767 OR2X1_LOC_40/Y OR2X1_LOC_674/Y 0.01fF
C18768 AND2X1_LOC_768/a_8_24# OR2X1_LOC_95/Y 0.01fF
C18769 OR2X1_LOC_106/a_36_216# OR2X1_LOC_47/Y 0.03fF
C18770 OR2X1_LOC_866/a_8_216# OR2X1_LOC_269/B 0.01fF
C18771 OR2X1_LOC_91/Y OR2X1_LOC_312/Y 0.03fF
C18772 OR2X1_LOC_26/Y AND2X1_LOC_840/B 0.05fF
C18773 AND2X1_LOC_729/B OR2X1_LOC_427/A 0.03fF
C18774 OR2X1_LOC_306/a_8_216# AND2X1_LOC_390/B 0.04fF
C18775 OR2X1_LOC_156/Y OR2X1_LOC_160/a_36_216# 0.00fF
C18776 AND2X1_LOC_59/Y AND2X1_LOC_79/Y 0.16fF
C18777 AND2X1_LOC_705/Y OR2X1_LOC_419/Y 0.00fF
C18778 OR2X1_LOC_748/A OR2X1_LOC_820/B 0.40fF
C18779 AND2X1_LOC_18/Y OR2X1_LOC_227/Y 0.03fF
C18780 AND2X1_LOC_216/A OR2X1_LOC_12/Y 0.02fF
C18781 OR2X1_LOC_810/A OR2X1_LOC_203/Y 0.10fF
C18782 AND2X1_LOC_564/A AND2X1_LOC_781/a_8_24# 0.07fF
C18783 OR2X1_LOC_434/a_8_216# OR2X1_LOC_814/A 0.02fF
C18784 AND2X1_LOC_650/Y OR2X1_LOC_52/B 0.00fF
C18785 OR2X1_LOC_453/a_8_216# OR2X1_LOC_453/Y 0.01fF
C18786 OR2X1_LOC_157/a_8_216# OR2X1_LOC_429/Y 0.03fF
C18787 AND2X1_LOC_42/B OR2X1_LOC_87/a_8_216# 0.01fF
C18788 OR2X1_LOC_318/a_8_216# OR2X1_LOC_318/B 0.08fF
C18789 OR2X1_LOC_46/A AND2X1_LOC_642/Y 0.17fF
C18790 OR2X1_LOC_6/B AND2X1_LOC_837/a_36_24# 0.00fF
C18791 AND2X1_LOC_840/B OR2X1_LOC_89/A 0.23fF
C18792 AND2X1_LOC_18/Y D_INPUT_1 5.02fF
C18793 OR2X1_LOC_759/A AND2X1_LOC_620/Y 0.03fF
C18794 OR2X1_LOC_40/Y AND2X1_LOC_624/B 0.05fF
C18795 OR2X1_LOC_160/B OR2X1_LOC_783/a_8_216# 0.01fF
C18796 OR2X1_LOC_779/Y OR2X1_LOC_66/A 0.01fF
C18797 OR2X1_LOC_614/Y OR2X1_LOC_196/a_36_216# 0.00fF
C18798 OR2X1_LOC_40/Y OR2X1_LOC_67/Y 3.78fF
C18799 OR2X1_LOC_476/B OR2X1_LOC_405/a_8_216# 0.03fF
C18800 AND2X1_LOC_598/a_36_24# OR2X1_LOC_485/A 0.00fF
C18801 AND2X1_LOC_718/a_8_24# OR2X1_LOC_31/Y 0.00fF
C18802 OR2X1_LOC_653/Y OR2X1_LOC_814/A 0.02fF
C18803 AND2X1_LOC_559/a_36_24# OR2X1_LOC_74/A 0.01fF
C18804 OR2X1_LOC_160/B OR2X1_LOC_737/a_8_216# 0.06fF
C18805 AND2X1_LOC_711/Y OR2X1_LOC_748/A 0.00fF
C18806 AND2X1_LOC_355/a_8_24# AND2X1_LOC_356/B 0.01fF
C18807 OR2X1_LOC_743/A AND2X1_LOC_454/A 0.00fF
C18808 AND2X1_LOC_350/Y OR2X1_LOC_265/Y 0.13fF
C18809 OR2X1_LOC_274/Y OR2X1_LOC_241/Y 0.78fF
C18810 OR2X1_LOC_272/Y OR2X1_LOC_52/B 0.05fF
C18811 AND2X1_LOC_814/a_8_24# AND2X1_LOC_624/A 0.01fF
C18812 OR2X1_LOC_344/A OR2X1_LOC_578/B 0.03fF
C18813 OR2X1_LOC_485/A AND2X1_LOC_717/B 1.11fF
C18814 OR2X1_LOC_441/Y AND2X1_LOC_812/a_8_24# 0.06fF
C18815 OR2X1_LOC_305/Y AND2X1_LOC_307/a_8_24# 0.01fF
C18816 OR2X1_LOC_529/Y OR2X1_LOC_530/Y 0.21fF
C18817 AND2X1_LOC_98/Y OR2X1_LOC_47/Y 0.02fF
C18818 OR2X1_LOC_689/a_8_216# OR2X1_LOC_31/Y 0.09fF
C18819 OR2X1_LOC_499/a_36_216# OR2X1_LOC_62/B 0.01fF
C18820 OR2X1_LOC_139/A OR2X1_LOC_140/Y 0.01fF
C18821 OR2X1_LOC_282/a_8_216# OR2X1_LOC_89/A 0.02fF
C18822 AND2X1_LOC_47/Y OR2X1_LOC_560/a_8_216# 0.01fF
C18823 OR2X1_LOC_462/B OR2X1_LOC_46/A 0.94fF
C18824 OR2X1_LOC_103/Y OR2X1_LOC_47/Y 0.03fF
C18825 AND2X1_LOC_128/a_8_24# OR2X1_LOC_6/A 0.01fF
C18826 OR2X1_LOC_154/A OR2X1_LOC_404/A 0.10fF
C18827 AND2X1_LOC_48/A OR2X1_LOC_87/B 0.21fF
C18828 OR2X1_LOC_702/A AND2X1_LOC_136/a_8_24# 0.01fF
C18829 OR2X1_LOC_273/Y OR2X1_LOC_74/A 0.02fF
C18830 INPUT_0 AND2X1_LOC_699/a_8_24# 0.02fF
C18831 OR2X1_LOC_680/A AND2X1_LOC_657/a_36_24# 0.01fF
C18832 OR2X1_LOC_147/A OR2X1_LOC_705/B 0.21fF
C18833 AND2X1_LOC_394/a_8_24# AND2X1_LOC_47/Y 0.04fF
C18834 OR2X1_LOC_440/A OR2X1_LOC_161/A 0.03fF
C18835 OR2X1_LOC_311/Y OR2X1_LOC_312/Y 0.11fF
C18836 AND2X1_LOC_327/a_8_24# AND2X1_LOC_116/Y 0.01fF
C18837 OR2X1_LOC_70/Y OR2X1_LOC_304/Y 0.32fF
C18838 OR2X1_LOC_103/a_8_216# OR2X1_LOC_47/Y 0.01fF
C18839 OR2X1_LOC_244/A OR2X1_LOC_267/a_8_216# 0.01fF
C18840 OR2X1_LOC_490/Y OR2X1_LOC_19/B 0.01fF
C18841 OR2X1_LOC_19/B OR2X1_LOC_74/A 0.07fF
C18842 OR2X1_LOC_809/a_36_216# OR2X1_LOC_532/B 0.01fF
C18843 AND2X1_LOC_640/a_36_24# OR2X1_LOC_26/Y 0.00fF
C18844 OR2X1_LOC_447/Y OR2X1_LOC_778/Y 0.03fF
C18845 AND2X1_LOC_840/a_8_24# OR2X1_LOC_419/Y 0.13fF
C18846 OR2X1_LOC_231/A OR2X1_LOC_215/a_8_216# 0.01fF
C18847 AND2X1_LOC_41/A OR2X1_LOC_512/Y 0.03fF
C18848 OR2X1_LOC_87/A OR2X1_LOC_783/A 0.02fF
C18849 AND2X1_LOC_723/Y AND2X1_LOC_222/Y 0.01fF
C18850 OR2X1_LOC_26/Y OR2X1_LOC_31/Y 8.00fF
C18851 AND2X1_LOC_711/Y OR2X1_LOC_628/Y 0.03fF
C18852 AND2X1_LOC_738/B OR2X1_LOC_533/a_8_216# 0.04fF
C18853 AND2X1_LOC_539/a_8_24# OR2X1_LOC_743/A 0.01fF
C18854 OR2X1_LOC_36/Y AND2X1_LOC_649/Y 0.01fF
C18855 OR2X1_LOC_3/Y AND2X1_LOC_477/A 0.03fF
C18856 AND2X1_LOC_568/a_8_24# AND2X1_LOC_477/A 0.01fF
C18857 OR2X1_LOC_500/A D_INPUT_1 0.10fF
C18858 OR2X1_LOC_100/Y AND2X1_LOC_609/a_8_24# 0.23fF
C18859 OR2X1_LOC_161/A OR2X1_LOC_446/A 0.02fF
C18860 OR2X1_LOC_36/Y AND2X1_LOC_648/B 0.03fF
C18861 OR2X1_LOC_256/A OR2X1_LOC_7/A 0.32fF
C18862 OR2X1_LOC_794/A OR2X1_LOC_318/B 0.00fF
C18863 OR2X1_LOC_70/A OR2X1_LOC_586/Y 0.01fF
C18864 OR2X1_LOC_160/A AND2X1_LOC_72/B 0.08fF
C18865 OR2X1_LOC_31/Y OR2X1_LOC_89/A 0.17fF
C18866 AND2X1_LOC_537/Y AND2X1_LOC_307/a_36_24# 0.01fF
C18867 OR2X1_LOC_130/A OR2X1_LOC_215/a_8_216# 0.03fF
C18868 OR2X1_LOC_218/Y AND2X1_LOC_3/Y 0.35fF
C18869 AND2X1_LOC_401/Y OR2X1_LOC_80/A 0.03fF
C18870 AND2X1_LOC_347/a_8_24# AND2X1_LOC_866/A 0.02fF
C18871 AND2X1_LOC_463/B AND2X1_LOC_463/a_8_24# 0.11fF
C18872 OR2X1_LOC_84/B OR2X1_LOC_786/Y 0.00fF
C18873 OR2X1_LOC_66/A AND2X1_LOC_246/a_36_24# 0.00fF
C18874 AND2X1_LOC_70/Y OR2X1_LOC_771/B 0.03fF
C18875 OR2X1_LOC_604/A OR2X1_LOC_183/Y 0.03fF
C18876 AND2X1_LOC_705/Y AND2X1_LOC_590/a_36_24# 0.00fF
C18877 OR2X1_LOC_74/A OR2X1_LOC_75/Y 0.00fF
C18878 OR2X1_LOC_639/A OR2X1_LOC_639/a_8_216# 0.39fF
C18879 OR2X1_LOC_244/a_8_216# OR2X1_LOC_140/Y 0.01fF
C18880 OR2X1_LOC_440/A AND2X1_LOC_51/Y 0.03fF
C18881 AND2X1_LOC_835/a_36_24# OR2X1_LOC_54/Y 0.00fF
C18882 OR2X1_LOC_7/A AND2X1_LOC_624/B 0.00fF
C18883 AND2X1_LOC_537/Y OR2X1_LOC_417/A 0.00fF
C18884 OR2X1_LOC_68/Y AND2X1_LOC_69/a_8_24# 0.23fF
C18885 OR2X1_LOC_7/A OR2X1_LOC_67/Y 0.03fF
C18886 OR2X1_LOC_139/A OR2X1_LOC_390/A 0.06fF
C18887 OR2X1_LOC_287/B OR2X1_LOC_366/a_8_216# 0.01fF
C18888 OR2X1_LOC_368/a_8_216# AND2X1_LOC_543/Y 0.01fF
C18889 OR2X1_LOC_118/a_8_216# OR2X1_LOC_595/A 0.07fF
C18890 OR2X1_LOC_399/A OR2X1_LOC_399/a_8_216# 0.47fF
C18891 OR2X1_LOC_185/A OR2X1_LOC_71/A 0.02fF
C18892 AND2X1_LOC_122/a_8_24# OR2X1_LOC_205/Y 0.03fF
C18893 OR2X1_LOC_813/A OR2X1_LOC_71/Y 0.35fF
C18894 AND2X1_LOC_50/a_8_24# INPUT_6 0.02fF
C18895 OR2X1_LOC_696/A OR2X1_LOC_25/Y 0.01fF
C18896 OR2X1_LOC_375/A OR2X1_LOC_367/B 0.03fF
C18897 OR2X1_LOC_272/Y AND2X1_LOC_216/A 0.30fF
C18898 AND2X1_LOC_539/Y AND2X1_LOC_436/Y 0.02fF
C18899 OR2X1_LOC_176/a_8_216# VDD 0.21fF
C18900 OR2X1_LOC_604/Y AND2X1_LOC_605/a_8_24# 0.01fF
C18901 OR2X1_LOC_216/A AND2X1_LOC_239/a_36_24# 0.01fF
C18902 AND2X1_LOC_721/Y AND2X1_LOC_658/B 0.03fF
C18903 AND2X1_LOC_469/Y AND2X1_LOC_469/a_8_24# 0.01fF
C18904 AND2X1_LOC_43/B OR2X1_LOC_515/Y 0.20fF
C18905 OR2X1_LOC_673/A OR2X1_LOC_532/B 0.61fF
C18906 OR2X1_LOC_323/A AND2X1_LOC_367/A 0.05fF
C18907 OR2X1_LOC_91/Y OR2X1_LOC_13/B 0.00fF
C18908 AND2X1_LOC_555/a_8_24# OR2X1_LOC_382/A 0.02fF
C18909 OR2X1_LOC_223/A OR2X1_LOC_532/B 0.03fF
C18910 AND2X1_LOC_745/a_8_24# OR2X1_LOC_797/B 0.23fF
C18911 AND2X1_LOC_705/Y OR2X1_LOC_604/A 0.71fF
C18912 OR2X1_LOC_691/A VDD 0.21fF
C18913 OR2X1_LOC_56/A OR2X1_LOC_428/A 1.21fF
C18914 OR2X1_LOC_482/Y AND2X1_LOC_499/a_8_24# 0.04fF
C18915 OR2X1_LOC_19/B AND2X1_LOC_647/Y 0.07fF
C18916 OR2X1_LOC_160/A AND2X1_LOC_36/Y 0.27fF
C18917 OR2X1_LOC_368/a_8_216# OR2X1_LOC_322/Y 0.03fF
C18918 AND2X1_LOC_732/B OR2X1_LOC_158/A 0.01fF
C18919 OR2X1_LOC_479/a_8_216# OR2X1_LOC_228/Y 0.01fF
C18920 OR2X1_LOC_56/A OR2X1_LOC_595/A 1.51fF
C18921 D_INPUT_0 OR2X1_LOC_86/A 0.19fF
C18922 AND2X1_LOC_362/B OR2X1_LOC_494/Y 0.07fF
C18923 AND2X1_LOC_672/a_8_24# D_INPUT_1 0.00fF
C18924 AND2X1_LOC_47/Y OR2X1_LOC_804/A 0.07fF
C18925 OR2X1_LOC_25/a_8_216# D_INPUT_6 0.01fF
C18926 OR2X1_LOC_502/A OR2X1_LOC_392/B 0.01fF
C18927 AND2X1_LOC_12/Y AND2X1_LOC_582/B 0.14fF
C18928 OR2X1_LOC_468/Y OR2X1_LOC_469/B 0.05fF
C18929 OR2X1_LOC_532/B OR2X1_LOC_705/B 0.01fF
C18930 VDD OR2X1_LOC_822/a_8_216# 0.00fF
C18931 OR2X1_LOC_756/B OR2X1_LOC_580/B 0.05fF
C18932 OR2X1_LOC_87/A OR2X1_LOC_308/Y 0.65fF
C18933 OR2X1_LOC_663/A OR2X1_LOC_161/B 0.03fF
C18934 AND2X1_LOC_59/Y OR2X1_LOC_356/B 0.11fF
C18935 AND2X1_LOC_41/A OR2X1_LOC_294/Y 0.09fF
C18936 OR2X1_LOC_629/Y OR2X1_LOC_563/A 0.02fF
C18937 VDD AND2X1_LOC_184/a_8_24# 0.00fF
C18938 AND2X1_LOC_729/Y OR2X1_LOC_144/a_36_216# 0.00fF
C18939 INPUT_0 OR2X1_LOC_13/Y 0.04fF
C18940 AND2X1_LOC_803/B OR2X1_LOC_679/a_8_216# 0.01fF
C18941 OR2X1_LOC_702/A OR2X1_LOC_112/A 0.03fF
C18942 OR2X1_LOC_7/A AND2X1_LOC_449/a_36_24# 0.01fF
C18943 OR2X1_LOC_676/Y OR2X1_LOC_702/a_8_216# 0.01fF
C18944 OR2X1_LOC_371/Y OR2X1_LOC_142/Y 0.06fF
C18945 OR2X1_LOC_354/A OR2X1_LOC_356/A 0.37fF
C18946 OR2X1_LOC_375/A AND2X1_LOC_416/a_8_24# 0.10fF
C18947 AND2X1_LOC_86/B AND2X1_LOC_36/Y 0.03fF
C18948 VDD OR2X1_LOC_531/Y 0.12fF
C18949 OR2X1_LOC_756/B OR2X1_LOC_648/B 0.10fF
C18950 AND2X1_LOC_41/A OR2X1_LOC_641/A 0.02fF
C18951 OR2X1_LOC_417/Y OR2X1_LOC_13/B 0.07fF
C18952 AND2X1_LOC_719/Y OR2X1_LOC_164/Y 0.09fF
C18953 OR2X1_LOC_316/Y AND2X1_LOC_473/Y 0.02fF
C18954 AND2X1_LOC_322/a_36_24# OR2X1_LOC_538/A 0.00fF
C18955 OR2X1_LOC_154/a_8_216# OR2X1_LOC_160/A 0.02fF
C18956 OR2X1_LOC_624/B AND2X1_LOC_36/Y 0.45fF
C18957 AND2X1_LOC_817/B OR2X1_LOC_770/A 0.00fF
C18958 OR2X1_LOC_36/Y OR2X1_LOC_56/a_8_216# 0.01fF
C18959 OR2X1_LOC_175/Y AND2X1_LOC_166/a_36_24# 0.00fF
C18960 VDD OR2X1_LOC_678/Y 0.14fF
C18961 OR2X1_LOC_311/Y OR2X1_LOC_13/B 0.10fF
C18962 OR2X1_LOC_36/Y AND2X1_LOC_465/A 0.08fF
C18963 VDD OR2X1_LOC_294/a_8_216# 0.21fF
C18964 OR2X1_LOC_538/a_8_216# OR2X1_LOC_160/B 0.01fF
C18965 AND2X1_LOC_773/Y OR2X1_LOC_39/A 0.07fF
C18966 VDD AND2X1_LOC_304/a_8_24# 0.00fF
C18967 AND2X1_LOC_554/Y OR2X1_LOC_12/Y 0.18fF
C18968 AND2X1_LOC_538/Y OR2X1_LOC_13/B -0.01fF
C18969 OR2X1_LOC_151/A OR2X1_LOC_620/Y 0.09fF
C18970 OR2X1_LOC_186/Y OR2X1_LOC_212/A 0.18fF
C18971 OR2X1_LOC_109/Y OR2X1_LOC_322/a_8_216# 0.02fF
C18972 AND2X1_LOC_784/A OR2X1_LOC_136/a_36_216# 0.00fF
C18973 AND2X1_LOC_452/Y OR2X1_LOC_603/Y 0.02fF
C18974 OR2X1_LOC_264/Y AND2X1_LOC_265/a_36_24# 0.00fF
C18975 AND2X1_LOC_486/Y OR2X1_LOC_40/Y 0.06fF
C18976 OR2X1_LOC_158/A OR2X1_LOC_625/Y 0.03fF
C18977 OR2X1_LOC_571/B OR2X1_LOC_113/B 0.01fF
C18978 AND2X1_LOC_51/Y AND2X1_LOC_238/a_8_24# 0.07fF
C18979 OR2X1_LOC_40/Y AND2X1_LOC_840/a_36_24# 0.00fF
C18980 OR2X1_LOC_45/B AND2X1_LOC_576/Y 0.09fF
C18981 OR2X1_LOC_154/A OR2X1_LOC_318/A 0.00fF
C18982 AND2X1_LOC_706/Y OR2X1_LOC_424/a_36_216# 0.01fF
C18983 AND2X1_LOC_64/Y OR2X1_LOC_629/A 0.18fF
C18984 OR2X1_LOC_438/Y AND2X1_LOC_657/Y 0.03fF
C18985 AND2X1_LOC_371/a_8_24# OR2X1_LOC_737/A 0.01fF
C18986 AND2X1_LOC_244/A OR2X1_LOC_44/Y 0.12fF
C18987 OR2X1_LOC_743/A AND2X1_LOC_783/B 0.01fF
C18988 AND2X1_LOC_322/a_8_24# OR2X1_LOC_620/Y 0.02fF
C18989 OR2X1_LOC_323/A OR2X1_LOC_74/A 0.15fF
C18990 OR2X1_LOC_296/Y OR2X1_LOC_140/B 0.03fF
C18991 OR2X1_LOC_317/a_8_216# AND2X1_LOC_92/Y 0.02fF
C18992 AND2X1_LOC_707/Y OR2X1_LOC_682/a_8_216# 0.01fF
C18993 OR2X1_LOC_364/A OR2X1_LOC_161/B 0.45fF
C18994 AND2X1_LOC_244/A AND2X1_LOC_288/a_8_24# 0.01fF
C18995 AND2X1_LOC_43/B OR2X1_LOC_549/A 0.07fF
C18996 AND2X1_LOC_850/A OR2X1_LOC_59/Y 0.07fF
C18997 OR2X1_LOC_185/Y OR2X1_LOC_161/B 0.12fF
C18998 OR2X1_LOC_40/Y AND2X1_LOC_811/B 0.02fF
C18999 VDD OR2X1_LOC_46/a_8_216# 0.21fF
C19000 OR2X1_LOC_278/Y AND2X1_LOC_860/A 0.03fF
C19001 OR2X1_LOC_841/a_8_216# AND2X1_LOC_92/Y 0.04fF
C19002 VDD OR2X1_LOC_811/A 0.64fF
C19003 OR2X1_LOC_16/A OR2X1_LOC_44/Y 0.06fF
C19004 OR2X1_LOC_26/Y AND2X1_LOC_464/A 0.03fF
C19005 AND2X1_LOC_95/Y AND2X1_LOC_18/Y 0.21fF
C19006 AND2X1_LOC_22/Y AND2X1_LOC_683/a_8_24# 0.11fF
C19007 OR2X1_LOC_154/A OR2X1_LOC_151/A 0.17fF
C19008 OR2X1_LOC_631/B OR2X1_LOC_294/Y 0.03fF
C19009 AND2X1_LOC_18/a_8_24# AND2X1_LOC_7/B 0.01fF
C19010 AND2X1_LOC_70/Y AND2X1_LOC_11/Y 0.77fF
C19011 AND2X1_LOC_784/Y OR2X1_LOC_680/A 0.13fF
C19012 AND2X1_LOC_773/Y AND2X1_LOC_211/B 0.10fF
C19013 D_INPUT_3 OR2X1_LOC_13/B 0.05fF
C19014 OR2X1_LOC_856/B AND2X1_LOC_92/Y 0.14fF
C19015 OR2X1_LOC_9/Y OR2X1_LOC_96/B 0.73fF
C19016 OR2X1_LOC_538/A OR2X1_LOC_623/B 0.00fF
C19017 OR2X1_LOC_127/Y VDD 0.00fF
C19018 OR2X1_LOC_287/B OR2X1_LOC_633/A 0.05fF
C19019 OR2X1_LOC_89/A AND2X1_LOC_213/B 0.00fF
C19020 OR2X1_LOC_49/A OR2X1_LOC_647/B 0.01fF
C19021 VDD OR2X1_LOC_404/a_8_216# 0.21fF
C19022 OR2X1_LOC_770/B AND2X1_LOC_3/Y 0.01fF
C19023 AND2X1_LOC_170/Y AND2X1_LOC_566/B 0.17fF
C19024 OR2X1_LOC_604/A OR2X1_LOC_511/Y 0.17fF
C19025 OR2X1_LOC_619/Y AND2X1_LOC_658/Y 0.09fF
C19026 OR2X1_LOC_715/B OR2X1_LOC_203/Y 0.00fF
C19027 OR2X1_LOC_348/Y OR2X1_LOC_375/A 0.01fF
C19028 OR2X1_LOC_40/Y AND2X1_LOC_716/a_8_24# 0.02fF
C19029 OR2X1_LOC_585/A OR2X1_LOC_829/A 0.05fF
C19030 OR2X1_LOC_203/Y AND2X1_LOC_626/a_8_24# 0.01fF
C19031 AND2X1_LOC_810/A AND2X1_LOC_337/B 0.02fF
C19032 AND2X1_LOC_191/B AND2X1_LOC_621/Y 0.01fF
C19033 AND2X1_LOC_520/Y AND2X1_LOC_222/a_8_24# 0.27fF
C19034 AND2X1_LOC_642/a_8_24# AND2X1_LOC_219/Y 0.01fF
C19035 OR2X1_LOC_640/Y OR2X1_LOC_640/a_8_216# -0.00fF
C19036 OR2X1_LOC_858/A OR2X1_LOC_185/A 0.00fF
C19037 OR2X1_LOC_690/A OR2X1_LOC_13/Y 0.02fF
C19038 OR2X1_LOC_17/Y AND2X1_LOC_639/B 0.26fF
C19039 OR2X1_LOC_426/B AND2X1_LOC_123/Y 0.03fF
C19040 OR2X1_LOC_9/Y AND2X1_LOC_852/Y 0.19fF
C19041 AND2X1_LOC_110/a_36_24# OR2X1_LOC_161/A 0.01fF
C19042 OR2X1_LOC_186/Y OR2X1_LOC_620/B 0.07fF
C19043 AND2X1_LOC_621/Y AND2X1_LOC_469/B 0.03fF
C19044 OR2X1_LOC_517/a_8_216# AND2X1_LOC_76/Y 0.01fF
C19045 OR2X1_LOC_129/a_8_216# OR2X1_LOC_26/Y 0.01fF
C19046 OR2X1_LOC_108/Y OR2X1_LOC_44/Y 0.07fF
C19047 OR2X1_LOC_100/Y OR2X1_LOC_502/A 0.04fF
C19048 AND2X1_LOC_753/a_8_24# AND2X1_LOC_41/A 0.03fF
C19049 OR2X1_LOC_653/A OR2X1_LOC_66/A 0.07fF
C19050 AND2X1_LOC_50/Y AND2X1_LOC_753/B 0.03fF
C19051 OR2X1_LOC_40/Y OR2X1_LOC_6/a_8_216# 0.01fF
C19052 AND2X1_LOC_848/a_8_24# OR2X1_LOC_59/Y 0.02fF
C19053 OR2X1_LOC_448/Y OR2X1_LOC_78/A 0.21fF
C19054 AND2X1_LOC_3/Y OR2X1_LOC_596/A 0.04fF
C19055 OR2X1_LOC_673/Y OR2X1_LOC_66/A 1.16fF
C19056 AND2X1_LOC_512/Y AND2X1_LOC_809/A 0.07fF
C19057 OR2X1_LOC_99/Y AND2X1_LOC_18/Y 0.20fF
C19058 OR2X1_LOC_613/Y AND2X1_LOC_658/A 0.01fF
C19059 AND2X1_LOC_59/Y OR2X1_LOC_168/B 0.22fF
C19060 AND2X1_LOC_555/a_8_24# OR2X1_LOC_261/Y 0.01fF
C19061 OR2X1_LOC_224/a_36_216# OR2X1_LOC_183/Y 0.00fF
C19062 AND2X1_LOC_99/A OR2X1_LOC_517/A 0.03fF
C19063 OR2X1_LOC_676/Y OR2X1_LOC_269/B 0.07fF
C19064 AND2X1_LOC_377/Y OR2X1_LOC_39/A 0.03fF
C19065 OR2X1_LOC_473/a_8_216# OR2X1_LOC_737/A 0.01fF
C19066 OR2X1_LOC_844/Y OR2X1_LOC_576/A 0.03fF
C19067 AND2X1_LOC_733/Y AND2X1_LOC_621/Y 0.05fF
C19068 D_INPUT_0 OR2X1_LOC_20/A 0.00fF
C19069 AND2X1_LOC_720/a_8_24# AND2X1_LOC_720/Y 0.00fF
C19070 AND2X1_LOC_61/Y AND2X1_LOC_852/Y 0.06fF
C19071 AND2X1_LOC_91/B OR2X1_LOC_447/Y 0.24fF
C19072 AND2X1_LOC_486/Y AND2X1_LOC_843/Y 0.39fF
C19073 AND2X1_LOC_121/a_8_24# OR2X1_LOC_44/Y 0.01fF
C19074 OR2X1_LOC_137/a_36_216# OR2X1_LOC_137/B 0.02fF
C19075 OR2X1_LOC_808/B OR2X1_LOC_732/B 0.10fF
C19076 OR2X1_LOC_496/Y OR2X1_LOC_51/Y 0.00fF
C19077 OR2X1_LOC_666/A AND2X1_LOC_806/A 1.62fF
C19078 OR2X1_LOC_151/A OR2X1_LOC_778/A 0.01fF
C19079 AND2X1_LOC_568/B AND2X1_LOC_211/B 0.01fF
C19080 AND2X1_LOC_70/Y OR2X1_LOC_217/a_8_216# 0.01fF
C19081 AND2X1_LOC_380/a_8_24# OR2X1_LOC_637/B 0.20fF
C19082 OR2X1_LOC_395/Y OR2X1_LOC_396/a_8_216# 0.40fF
C19083 OR2X1_LOC_354/A AND2X1_LOC_43/B 0.00fF
C19084 OR2X1_LOC_834/A OR2X1_LOC_269/B 0.02fF
C19085 AND2X1_LOC_41/A OR2X1_LOC_194/Y 0.08fF
C19086 OR2X1_LOC_95/Y AND2X1_LOC_227/a_8_24# 0.01fF
C19087 INPUT_0 OR2X1_LOC_82/a_8_216# 0.03fF
C19088 OR2X1_LOC_604/A AND2X1_LOC_345/Y 0.07fF
C19089 AND2X1_LOC_12/Y OR2X1_LOC_623/B 0.03fF
C19090 AND2X1_LOC_109/a_8_24# OR2X1_LOC_390/B 0.05fF
C19091 OR2X1_LOC_364/A OR2X1_LOC_435/B 0.01fF
C19092 OR2X1_LOC_22/Y OR2X1_LOC_12/Y 0.51fF
C19093 OR2X1_LOC_185/Y OR2X1_LOC_435/B 0.20fF
C19094 OR2X1_LOC_510/Y OR2X1_LOC_721/Y 0.03fF
C19095 OR2X1_LOC_478/a_8_216# OR2X1_LOC_467/a_8_216# 0.47fF
C19096 OR2X1_LOC_477/Y OR2X1_LOC_470/A 0.01fF
C19097 OR2X1_LOC_810/A OR2X1_LOC_78/B 0.00fF
C19098 AND2X1_LOC_392/A AND2X1_LOC_212/B 0.05fF
C19099 AND2X1_LOC_334/Y AND2X1_LOC_640/Y 1.13fF
C19100 OR2X1_LOC_18/Y OR2X1_LOC_48/B 1.89fF
C19101 OR2X1_LOC_394/Y OR2X1_LOC_393/Y 0.10fF
C19102 OR2X1_LOC_459/A AND2X1_LOC_472/B 0.03fF
C19103 OR2X1_LOC_753/A OR2X1_LOC_394/a_8_216# 0.33fF
C19104 AND2X1_LOC_64/Y OR2X1_LOC_473/A 0.07fF
C19105 OR2X1_LOC_254/B OR2X1_LOC_147/B 0.03fF
C19106 OR2X1_LOC_517/a_8_216# OR2X1_LOC_52/B 0.03fF
C19107 AND2X1_LOC_319/A OR2X1_LOC_92/Y 0.06fF
C19108 AND2X1_LOC_370/a_8_24# AND2X1_LOC_866/A 0.08fF
C19109 OR2X1_LOC_316/Y AND2X1_LOC_649/a_8_24# 0.01fF
C19110 AND2X1_LOC_863/a_8_24# OR2X1_LOC_36/Y 0.02fF
C19111 OR2X1_LOC_199/a_8_216# AND2X1_LOC_47/Y 0.01fF
C19112 OR2X1_LOC_3/Y OR2X1_LOC_816/a_36_216# 0.03fF
C19113 AND2X1_LOC_222/Y OR2X1_LOC_142/Y 0.03fF
C19114 OR2X1_LOC_443/a_36_216# OR2X1_LOC_161/B 0.00fF
C19115 AND2X1_LOC_711/Y AND2X1_LOC_861/a_8_24# 0.07fF
C19116 OR2X1_LOC_833/a_36_216# AND2X1_LOC_56/B 0.00fF
C19117 OR2X1_LOC_592/A OR2X1_LOC_78/A 0.02fF
C19118 AND2X1_LOC_95/Y OR2X1_LOC_500/A 0.02fF
C19119 D_INPUT_0 AND2X1_LOC_65/A 0.09fF
C19120 AND2X1_LOC_76/a_8_24# OR2X1_LOC_85/A 0.01fF
C19121 OR2X1_LOC_251/Y OR2X1_LOC_251/a_36_216# 0.00fF
C19122 OR2X1_LOC_502/A OR2X1_LOC_610/Y 0.01fF
C19123 OR2X1_LOC_541/B OR2X1_LOC_541/a_8_216# 0.49fF
C19124 AND2X1_LOC_477/A AND2X1_LOC_477/Y 0.23fF
C19125 OR2X1_LOC_333/B OR2X1_LOC_174/A 0.08fF
C19126 OR2X1_LOC_6/B OR2X1_LOC_62/B 0.30fF
C19127 OR2X1_LOC_278/Y AND2X1_LOC_287/Y 0.01fF
C19128 AND2X1_LOC_429/a_8_24# INPUT_6 0.00fF
C19129 AND2X1_LOC_219/a_8_24# OR2X1_LOC_416/Y 0.01fF
C19130 VDD AND2X1_LOC_115/a_8_24# 0.00fF
C19131 OR2X1_LOC_468/Y OR2X1_LOC_211/a_8_216# 0.01fF
C19132 AND2X1_LOC_334/Y OR2X1_LOC_416/Y 0.01fF
C19133 AND2X1_LOC_723/Y OR2X1_LOC_74/A 0.04fF
C19134 OR2X1_LOC_276/B AND2X1_LOC_256/a_8_24# 0.01fF
C19135 AND2X1_LOC_95/Y AND2X1_LOC_413/a_8_24# 0.17fF
C19136 AND2X1_LOC_212/A AND2X1_LOC_863/Y 0.13fF
C19137 AND2X1_LOC_523/Y OR2X1_LOC_59/Y 0.03fF
C19138 OR2X1_LOC_144/Y OR2X1_LOC_89/A 0.10fF
C19139 OR2X1_LOC_185/A OR2X1_LOC_593/a_8_216# 0.01fF
C19140 OR2X1_LOC_510/Y OR2X1_LOC_375/A 0.08fF
C19141 AND2X1_LOC_552/A OR2X1_LOC_31/Y 0.01fF
C19142 OR2X1_LOC_58/Y OR2X1_LOC_412/a_8_216# 0.01fF
C19143 AND2X1_LOC_658/B OR2X1_LOC_628/Y 0.00fF
C19144 AND2X1_LOC_486/Y OR2X1_LOC_7/A 0.05fF
C19145 OR2X1_LOC_160/B OR2X1_LOC_335/B 0.03fF
C19146 AND2X1_LOC_17/Y AND2X1_LOC_11/Y 0.98fF
C19147 OR2X1_LOC_292/Y OR2X1_LOC_481/A 0.02fF
C19148 OR2X1_LOC_45/B OR2X1_LOC_29/a_8_216# 0.01fF
C19149 OR2X1_LOC_22/A OR2X1_LOC_380/a_8_216# 0.01fF
C19150 OR2X1_LOC_265/Y AND2X1_LOC_266/Y 0.55fF
C19151 OR2X1_LOC_31/Y AND2X1_LOC_194/Y 0.02fF
C19152 AND2X1_LOC_541/Y OR2X1_LOC_95/Y 0.01fF
C19153 AND2X1_LOC_629/Y AND2X1_LOC_629/a_8_24# 0.00fF
C19154 OR2X1_LOC_385/Y OR2X1_LOC_48/B 0.03fF
C19155 OR2X1_LOC_36/Y OR2X1_LOC_237/Y 0.08fF
C19156 OR2X1_LOC_778/Y OR2X1_LOC_161/A 0.04fF
C19157 OR2X1_LOC_504/Y AND2X1_LOC_508/B 0.01fF
C19158 AND2X1_LOC_699/a_8_24# AND2X1_LOC_7/B 0.02fF
C19159 AND2X1_LOC_73/a_8_24# OR2X1_LOC_62/B 0.00fF
C19160 OR2X1_LOC_426/B OR2X1_LOC_813/A 0.03fF
C19161 AND2X1_LOC_64/Y OR2X1_LOC_228/Y 0.07fF
C19162 OR2X1_LOC_448/Y OR2X1_LOC_155/A 0.02fF
C19163 OR2X1_LOC_496/Y OR2X1_LOC_680/A 0.12fF
C19164 OR2X1_LOC_391/B OR2X1_LOC_848/A 0.40fF
C19165 OR2X1_LOC_810/A OR2X1_LOC_375/A 0.05fF
C19166 AND2X1_LOC_7/B OR2X1_LOC_675/Y 0.02fF
C19167 OR2X1_LOC_126/a_8_216# AND2X1_LOC_573/A 0.01fF
C19168 OR2X1_LOC_235/B OR2X1_LOC_62/a_8_216# 0.02fF
C19169 OR2X1_LOC_599/A OR2X1_LOC_591/A 0.05fF
C19170 OR2X1_LOC_604/A AND2X1_LOC_451/Y 0.81fF
C19171 OR2X1_LOC_114/Y OR2X1_LOC_631/B 0.10fF
C19172 OR2X1_LOC_280/a_36_216# OR2X1_LOC_39/A 0.00fF
C19173 OR2X1_LOC_97/A OR2X1_LOC_358/A 0.00fF
C19174 OR2X1_LOC_158/A OR2X1_LOC_3/B 0.07fF
C19175 AND2X1_LOC_123/a_36_24# OR2X1_LOC_67/A 0.00fF
C19176 OR2X1_LOC_84/B OR2X1_LOC_204/Y 0.01fF
C19177 OR2X1_LOC_463/B AND2X1_LOC_3/Y 0.00fF
C19178 AND2X1_LOC_311/a_36_24# D_INPUT_0 0.00fF
C19179 OR2X1_LOC_476/B OR2X1_LOC_61/a_36_216# 0.01fF
C19180 OR2X1_LOC_135/Y AND2X1_LOC_643/a_8_24# 0.03fF
C19181 OR2X1_LOC_107/a_8_216# OR2X1_LOC_95/Y 0.01fF
C19182 AND2X1_LOC_606/a_8_24# D_INPUT_1 0.01fF
C19183 AND2X1_LOC_711/Y AND2X1_LOC_848/a_8_24# 0.19fF
C19184 OR2X1_LOC_596/A OR2X1_LOC_194/a_8_216# 0.01fF
C19185 AND2X1_LOC_56/B OR2X1_LOC_355/B 0.03fF
C19186 OR2X1_LOC_51/Y AND2X1_LOC_851/B 0.05fF
C19187 OR2X1_LOC_141/B OR2X1_LOC_204/Y 0.20fF
C19188 OR2X1_LOC_405/A OR2X1_LOC_473/Y 0.00fF
C19189 OR2X1_LOC_73/a_8_216# OR2X1_LOC_85/A 0.08fF
C19190 OR2X1_LOC_45/Y OR2X1_LOC_431/Y 0.16fF
C19191 OR2X1_LOC_552/A OR2X1_LOC_161/B 0.03fF
C19192 AND2X1_LOC_649/B OR2X1_LOC_416/Y 0.04fF
C19193 OR2X1_LOC_495/a_8_216# AND2X1_LOC_717/B 0.04fF
C19194 AND2X1_LOC_12/Y AND2X1_LOC_13/a_36_24# 0.01fF
C19195 OR2X1_LOC_248/Y OR2X1_LOC_7/A 0.78fF
C19196 OR2X1_LOC_62/A OR2X1_LOC_78/A 0.02fF
C19197 AND2X1_LOC_791/a_8_24# AND2X1_LOC_792/B 0.01fF
C19198 VDD AND2X1_LOC_237/a_8_24# -0.00fF
C19199 OR2X1_LOC_427/A OR2X1_LOC_46/A 0.27fF
C19200 OR2X1_LOC_805/A OR2X1_LOC_719/A 0.03fF
C19201 OR2X1_LOC_161/B OR2X1_LOC_568/A 0.07fF
C19202 OR2X1_LOC_824/a_8_216# OR2X1_LOC_824/Y 0.01fF
C19203 OR2X1_LOC_502/A OR2X1_LOC_532/B 0.18fF
C19204 OR2X1_LOC_285/B AND2X1_LOC_282/a_8_24# 0.20fF
C19205 OR2X1_LOC_506/B OR2X1_LOC_244/B 0.01fF
C19206 VDD AND2X1_LOC_203/Y 0.25fF
C19207 OR2X1_LOC_161/B OR2X1_LOC_578/B 0.16fF
C19208 OR2X1_LOC_666/Y OR2X1_LOC_7/A 0.02fF
C19209 AND2X1_LOC_612/B OR2X1_LOC_647/B 0.03fF
C19210 AND2X1_LOC_40/a_8_24# AND2X1_LOC_31/Y 0.01fF
C19211 AND2X1_LOC_84/a_36_24# OR2X1_LOC_585/A 0.01fF
C19212 OR2X1_LOC_679/A OR2X1_LOC_427/A 0.03fF
C19213 OR2X1_LOC_600/a_8_216# OR2X1_LOC_419/Y 0.39fF
C19214 OR2X1_LOC_441/Y AND2X1_LOC_796/Y 0.03fF
C19215 OR2X1_LOC_846/a_36_216# OR2X1_LOC_846/A 0.01fF
C19216 OR2X1_LOC_238/Y OR2X1_LOC_371/Y 0.02fF
C19217 AND2X1_LOC_69/a_8_24# OR2X1_LOC_506/A 0.17fF
C19218 OR2X1_LOC_113/A OR2X1_LOC_161/A 0.01fF
C19219 OR2X1_LOC_151/A OR2X1_LOC_560/A 0.03fF
C19220 OR2X1_LOC_643/A AND2X1_LOC_51/Y 0.03fF
C19221 OR2X1_LOC_848/A OR2X1_LOC_772/Y 0.04fF
C19222 AND2X1_LOC_40/Y OR2X1_LOC_468/a_36_216# 0.00fF
C19223 OR2X1_LOC_848/A OR2X1_LOC_846/A 0.09fF
C19224 OR2X1_LOC_778/Y AND2X1_LOC_51/Y 0.04fF
C19225 OR2X1_LOC_643/Y OR2X1_LOC_358/B 0.00fF
C19226 OR2X1_LOC_687/Y OR2X1_LOC_196/B 0.65fF
C19227 AND2X1_LOC_227/Y OR2X1_LOC_427/A 0.03fF
C19228 OR2X1_LOC_268/a_8_216# OR2X1_LOC_6/A 0.06fF
C19229 AND2X1_LOC_727/A AND2X1_LOC_354/B 0.04fF
C19230 AND2X1_LOC_12/Y OR2X1_LOC_544/A 0.05fF
C19231 OR2X1_LOC_643/A OR2X1_LOC_849/a_8_216# 0.01fF
C19232 OR2X1_LOC_367/B OR2X1_LOC_549/A 0.12fF
C19233 OR2X1_LOC_529/a_8_216# OR2X1_LOC_95/Y 0.01fF
C19234 OR2X1_LOC_22/Y AND2X1_LOC_650/Y 0.12fF
C19235 OR2X1_LOC_275/A OR2X1_LOC_74/A 0.08fF
C19236 OR2X1_LOC_300/Y AND2X1_LOC_786/Y 0.04fF
C19237 OR2X1_LOC_419/Y AND2X1_LOC_477/a_8_24# 0.12fF
C19238 OR2X1_LOC_400/A OR2X1_LOC_532/B 0.00fF
C19239 AND2X1_LOC_687/Y OR2X1_LOC_44/Y 0.02fF
C19240 AND2X1_LOC_56/a_8_24# OR2X1_LOC_375/A 0.02fF
C19241 OR2X1_LOC_92/Y AND2X1_LOC_721/A 0.06fF
C19242 OR2X1_LOC_503/Y AND2X1_LOC_573/A 0.01fF
C19243 OR2X1_LOC_196/Y AND2X1_LOC_36/Y 0.09fF
C19244 AND2X1_LOC_47/Y OR2X1_LOC_130/A 0.05fF
C19245 AND2X1_LOC_753/B OR2X1_LOC_214/B 0.00fF
C19246 AND2X1_LOC_1/Y OR2X1_LOC_636/B 0.01fF
C19247 OR2X1_LOC_78/B AND2X1_LOC_609/a_36_24# 0.00fF
C19248 OR2X1_LOC_146/Y AND2X1_LOC_621/Y 0.02fF
C19249 OR2X1_LOC_776/a_8_216# OR2X1_LOC_318/B 0.01fF
C19250 OR2X1_LOC_133/a_8_216# AND2X1_LOC_789/Y 0.11fF
C19251 AND2X1_LOC_365/A AND2X1_LOC_798/A 0.26fF
C19252 AND2X1_LOC_336/a_36_24# OR2X1_LOC_22/Y 0.01fF
C19253 AND2X1_LOC_47/Y AND2X1_LOC_7/a_8_24# 0.01fF
C19254 OR2X1_LOC_486/Y OR2X1_LOC_182/a_8_216# 0.03fF
C19255 AND2X1_LOC_18/Y OR2X1_LOC_269/A 0.01fF
C19256 AND2X1_LOC_64/Y OR2X1_LOC_562/A 0.09fF
C19257 AND2X1_LOC_47/Y AND2X1_LOC_292/a_8_24# 0.02fF
C19258 OR2X1_LOC_516/Y AND2X1_LOC_785/Y 0.11fF
C19259 OR2X1_LOC_272/Y OR2X1_LOC_22/Y 0.05fF
C19260 AND2X1_LOC_785/A AND2X1_LOC_786/Y 0.01fF
C19261 OR2X1_LOC_542/B OR2X1_LOC_366/Y 0.06fF
C19262 AND2X1_LOC_554/B INPUT_1 0.03fF
C19263 OR2X1_LOC_435/B AND2X1_LOC_432/a_8_24# 0.00fF
C19264 AND2X1_LOC_81/B OR2X1_LOC_786/Y 0.14fF
C19265 AND2X1_LOC_31/Y OR2X1_LOC_708/Y 0.01fF
C19266 OR2X1_LOC_673/Y OR2X1_LOC_84/A 0.01fF
C19267 AND2X1_LOC_18/Y AND2X1_LOC_41/Y 0.06fF
C19268 VDD OR2X1_LOC_424/Y 0.09fF
C19269 AND2X1_LOC_40/Y OR2X1_LOC_567/a_8_216# 0.01fF
C19270 VDD OR2X1_LOC_777/B 0.99fF
C19271 OR2X1_LOC_427/A OR2X1_LOC_753/Y 0.33fF
C19272 AND2X1_LOC_330/a_8_24# OR2X1_LOC_13/B 0.01fF
C19273 OR2X1_LOC_497/a_36_216# OR2X1_LOC_184/Y 0.00fF
C19274 OR2X1_LOC_440/A OR2X1_LOC_787/Y 0.07fF
C19275 AND2X1_LOC_779/a_8_24# AND2X1_LOC_779/Y 0.00fF
C19276 OR2X1_LOC_202/a_36_216# OR2X1_LOC_814/A 0.01fF
C19277 OR2X1_LOC_404/Y AND2X1_LOC_107/a_36_24# 0.00fF
C19278 OR2X1_LOC_31/Y OR2X1_LOC_17/Y 0.06fF
C19279 OR2X1_LOC_279/Y AND2X1_LOC_849/a_8_24# 0.00fF
C19280 AND2X1_LOC_390/B OR2X1_LOC_95/Y 0.01fF
C19281 AND2X1_LOC_40/Y OR2X1_LOC_348/B 0.09fF
C19282 OR2X1_LOC_278/Y AND2X1_LOC_562/Y 0.03fF
C19283 OR2X1_LOC_263/a_8_216# OR2X1_LOC_19/B 0.01fF
C19284 VDD D_INPUT_6 0.24fF
C19285 OR2X1_LOC_825/a_8_216# OR2X1_LOC_95/Y 0.01fF
C19286 OR2X1_LOC_516/Y AND2X1_LOC_500/B 0.04fF
C19287 AND2X1_LOC_95/a_8_24# AND2X1_LOC_36/Y 0.01fF
C19288 OR2X1_LOC_685/B OR2X1_LOC_451/B 0.16fF
C19289 AND2X1_LOC_70/Y OR2X1_LOC_593/B 2.91fF
C19290 OR2X1_LOC_185/A AND2X1_LOC_31/Y 0.39fF
C19291 OR2X1_LOC_86/a_8_216# OR2X1_LOC_67/Y 0.01fF
C19292 OR2X1_LOC_597/Y OR2X1_LOC_585/A 0.01fF
C19293 OR2X1_LOC_622/A OR2X1_LOC_622/B 0.16fF
C19294 OR2X1_LOC_696/A OR2X1_LOC_421/A 0.07fF
C19295 OR2X1_LOC_256/Y OR2X1_LOC_437/A 0.03fF
C19296 OR2X1_LOC_696/A AND2X1_LOC_563/A 0.00fF
C19297 AND2X1_LOC_48/A OR2X1_LOC_532/B 0.04fF
C19298 OR2X1_LOC_54/a_36_216# OR2X1_LOC_46/A 0.00fF
C19299 OR2X1_LOC_736/Y AND2X1_LOC_7/B 3.53fF
C19300 AND2X1_LOC_727/A AND2X1_LOC_863/Y 0.00fF
C19301 OR2X1_LOC_605/a_36_216# OR2X1_LOC_223/A 0.00fF
C19302 OR2X1_LOC_665/Y AND2X1_LOC_793/Y 0.01fF
C19303 OR2X1_LOC_45/B OR2X1_LOC_16/A 0.24fF
C19304 OR2X1_LOC_19/B OR2X1_LOC_607/Y 0.05fF
C19305 OR2X1_LOC_65/B AND2X1_LOC_217/a_8_24# 0.17fF
C19306 OR2X1_LOC_43/A OR2X1_LOC_761/a_8_216# 0.02fF
C19307 OR2X1_LOC_62/B AND2X1_LOC_47/Y 0.27fF
C19308 OR2X1_LOC_604/A AND2X1_LOC_465/A 0.10fF
C19309 OR2X1_LOC_624/A OR2X1_LOC_446/B 0.10fF
C19310 OR2X1_LOC_421/A AND2X1_LOC_715/Y 0.01fF
C19311 AND2X1_LOC_754/a_36_24# AND2X1_LOC_22/Y 0.00fF
C19312 VDD OR2X1_LOC_831/B 0.25fF
C19313 AND2X1_LOC_370/a_8_24# OR2X1_LOC_40/Y 0.02fF
C19314 OR2X1_LOC_566/A VDD 0.00fF
C19315 OR2X1_LOC_325/a_8_216# OR2X1_LOC_532/Y 0.03fF
C19316 OR2X1_LOC_188/a_8_216# VDD -0.00fF
C19317 OR2X1_LOC_78/A OR2X1_LOC_170/a_8_216# 0.03fF
C19318 OR2X1_LOC_156/Y VDD 0.06fF
C19319 VDD AND2X1_LOC_242/B 0.23fF
C19320 OR2X1_LOC_400/a_8_216# AND2X1_LOC_36/Y 0.01fF
C19321 OR2X1_LOC_329/a_36_216# OR2X1_LOC_16/A 0.00fF
C19322 AND2X1_LOC_22/Y AND2X1_LOC_18/Y 13.06fF
C19323 OR2X1_LOC_720/Y OR2X1_LOC_66/A 0.01fF
C19324 AND2X1_LOC_521/a_8_24# OR2X1_LOC_523/B 0.01fF
C19325 OR2X1_LOC_45/B OR2X1_LOC_108/Y 0.02fF
C19326 OR2X1_LOC_847/B OR2X1_LOC_80/A 0.05fF
C19327 AND2X1_LOC_707/Y VDD 0.74fF
C19328 OR2X1_LOC_641/Y AND2X1_LOC_7/B 0.06fF
C19329 INPUT_5 AND2X1_LOC_409/B 0.26fF
C19330 OR2X1_LOC_696/A AND2X1_LOC_718/a_36_24# 0.01fF
C19331 OR2X1_LOC_485/Y OR2X1_LOC_12/Y 0.03fF
C19332 OR2X1_LOC_154/A OR2X1_LOC_714/A 0.03fF
C19333 OR2X1_LOC_847/A AND2X1_LOC_36/Y 0.00fF
C19334 OR2X1_LOC_303/a_8_216# OR2X1_LOC_703/A 0.01fF
C19335 OR2X1_LOC_121/Y OR2X1_LOC_140/A 0.00fF
C19336 OR2X1_LOC_447/A AND2X1_LOC_36/Y 0.03fF
C19337 AND2X1_LOC_127/a_8_24# AND2X1_LOC_72/B 0.01fF
C19338 OR2X1_LOC_421/Y AND2X1_LOC_448/a_8_24# -0.00fF
C19339 OR2X1_LOC_684/a_8_216# OR2X1_LOC_16/A 0.02fF
C19340 OR2X1_LOC_136/Y AND2X1_LOC_364/Y 0.01fF
C19341 OR2X1_LOC_113/B OR2X1_LOC_772/A 0.01fF
C19342 AND2X1_LOC_212/A OR2X1_LOC_309/Y 0.01fF
C19343 OR2X1_LOC_435/Y AND2X1_LOC_31/Y 0.14fF
C19344 VDD OR2X1_LOC_344/A 0.35fF
C19345 OR2X1_LOC_158/A AND2X1_LOC_535/Y 0.03fF
C19346 OR2X1_LOC_744/A OR2X1_LOC_816/A 0.07fF
C19347 OR2X1_LOC_160/A OR2X1_LOC_469/B 0.00fF
C19348 OR2X1_LOC_215/Y OR2X1_LOC_539/B 0.03fF
C19349 AND2X1_LOC_70/Y AND2X1_LOC_256/a_8_24# 0.02fF
C19350 AND2X1_LOC_47/Y AND2X1_LOC_279/a_36_24# 0.00fF
C19351 OR2X1_LOC_274/a_8_216# OR2X1_LOC_121/A 0.01fF
C19352 OR2X1_LOC_170/A OR2X1_LOC_788/B 0.03fF
C19353 AND2X1_LOC_806/A OR2X1_LOC_13/B 0.02fF
C19354 OR2X1_LOC_26/Y OR2X1_LOC_385/a_36_216# 0.03fF
C19355 OR2X1_LOC_31/Y OR2X1_LOC_588/A 0.00fF
C19356 OR2X1_LOC_62/B OR2X1_LOC_598/A 0.00fF
C19357 OR2X1_LOC_201/A OR2X1_LOC_392/B 0.03fF
C19358 OR2X1_LOC_64/Y AND2X1_LOC_563/Y 0.02fF
C19359 OR2X1_LOC_468/Y OR2X1_LOC_535/a_8_216# 0.01fF
C19360 OR2X1_LOC_235/B AND2X1_LOC_44/Y 0.09fF
C19361 OR2X1_LOC_621/A AND2X1_LOC_18/Y 0.17fF
C19362 OR2X1_LOC_49/A INPUT_0 0.22fF
C19363 OR2X1_LOC_510/A AND2X1_LOC_505/a_8_24# 0.24fF
C19364 OR2X1_LOC_808/B AND2X1_LOC_7/B 0.03fF
C19365 AND2X1_LOC_363/a_36_24# AND2X1_LOC_363/Y 0.02fF
C19366 VDD OR2X1_LOC_686/A 0.21fF
C19367 AND2X1_LOC_675/A AND2X1_LOC_795/Y 0.48fF
C19368 OR2X1_LOC_269/B AND2X1_LOC_591/a_8_24# -0.01fF
C19369 AND2X1_LOC_866/B GATE_579 0.03fF
C19370 AND2X1_LOC_592/Y AND2X1_LOC_738/B 0.01fF
C19371 OR2X1_LOC_604/A OR2X1_LOC_600/a_8_216# 0.01fF
C19372 OR2X1_LOC_426/B AND2X1_LOC_606/a_8_24# 0.11fF
C19373 AND2X1_LOC_212/A OR2X1_LOC_744/A 0.03fF
C19374 AND2X1_LOC_47/Y OR2X1_LOC_365/B 0.00fF
C19375 OR2X1_LOC_491/a_8_216# OR2X1_LOC_744/A 0.02fF
C19376 OR2X1_LOC_528/Y OR2X1_LOC_56/A 0.32fF
C19377 OR2X1_LOC_22/A OR2X1_LOC_588/a_36_216# 0.00fF
C19378 INPUT_0 OR2X1_LOC_596/A 0.03fF
C19379 OR2X1_LOC_715/B OR2X1_LOC_78/B 0.10fF
C19380 OR2X1_LOC_160/B AND2X1_LOC_110/a_8_24# 0.01fF
C19381 OR2X1_LOC_800/Y OR2X1_LOC_801/a_8_216# 0.39fF
C19382 AND2X1_LOC_658/B AND2X1_LOC_508/B 0.03fF
C19383 AND2X1_LOC_91/B OR2X1_LOC_161/A 0.11fF
C19384 AND2X1_LOC_787/a_8_24# AND2X1_LOC_787/A 0.03fF
C19385 OR2X1_LOC_78/A OR2X1_LOC_629/B 0.02fF
C19386 OR2X1_LOC_764/a_8_216# OR2X1_LOC_48/B 0.02fF
C19387 OR2X1_LOC_304/a_36_216# OR2X1_LOC_48/B 0.00fF
C19388 OR2X1_LOC_74/A OR2X1_LOC_142/Y 0.07fF
C19389 OR2X1_LOC_422/a_36_216# OR2X1_LOC_12/Y 0.02fF
C19390 OR2X1_LOC_417/A AND2X1_LOC_563/Y 0.03fF
C19391 AND2X1_LOC_539/Y AND2X1_LOC_655/A 0.01fF
C19392 OR2X1_LOC_18/Y OR2X1_LOC_764/a_8_216# 0.01fF
C19393 AND2X1_LOC_474/A AND2X1_LOC_243/Y 0.07fF
C19394 OR2X1_LOC_786/Y OR2X1_LOC_66/Y 0.91fF
C19395 AND2X1_LOC_345/a_8_24# AND2X1_LOC_789/Y 0.01fF
C19396 AND2X1_LOC_70/Y OR2X1_LOC_645/a_36_216# 0.00fF
C19397 AND2X1_LOC_40/Y AND2X1_LOC_65/A 0.55fF
C19398 OR2X1_LOC_235/B OR2X1_LOC_600/A 0.07fF
C19399 AND2X1_LOC_212/Y AND2X1_LOC_804/Y 0.02fF
C19400 OR2X1_LOC_382/Y OR2X1_LOC_40/Y 0.01fF
C19401 OR2X1_LOC_696/A AND2X1_LOC_512/a_8_24# 0.02fF
C19402 OR2X1_LOC_409/B OR2X1_LOC_377/a_8_216# 0.02fF
C19403 AND2X1_LOC_191/B OR2X1_LOC_59/Y 0.07fF
C19404 OR2X1_LOC_706/A AND2X1_LOC_18/Y 0.01fF
C19405 OR2X1_LOC_186/Y OR2X1_LOC_220/B 0.05fF
C19406 OR2X1_LOC_696/A AND2X1_LOC_717/B 0.06fF
C19407 AND2X1_LOC_469/B OR2X1_LOC_59/Y 0.03fF
C19408 OR2X1_LOC_674/a_8_216# OR2X1_LOC_51/Y 0.01fF
C19409 AND2X1_LOC_574/a_8_24# AND2X1_LOC_570/Y 0.01fF
C19410 OR2X1_LOC_510/A AND2X1_LOC_40/Y 0.01fF
C19411 OR2X1_LOC_257/Y AND2X1_LOC_259/a_8_24# 0.23fF
C19412 AND2X1_LOC_560/a_8_24# OR2X1_LOC_89/A 0.01fF
C19413 OR2X1_LOC_447/Y OR2X1_LOC_446/B 0.09fF
C19414 OR2X1_LOC_91/Y OR2X1_LOC_428/A 0.03fF
C19415 AND2X1_LOC_46/a_8_24# AND2X1_LOC_36/Y 0.03fF
C19416 AND2X1_LOC_64/Y OR2X1_LOC_287/B 0.07fF
C19417 OR2X1_LOC_12/Y OR2X1_LOC_39/A 1.16fF
C19418 AND2X1_LOC_705/Y AND2X1_LOC_447/a_8_24# 0.05fF
C19419 AND2X1_LOC_810/A AND2X1_LOC_388/a_8_24# 0.01fF
C19420 AND2X1_LOC_738/B AND2X1_LOC_512/Y 1.11fF
C19421 AND2X1_LOC_215/Y OR2X1_LOC_290/Y 0.07fF
C19422 OR2X1_LOC_318/a_8_216# AND2X1_LOC_59/Y 0.01fF
C19423 AND2X1_LOC_181/Y OR2X1_LOC_18/Y 0.03fF
C19424 AND2X1_LOC_512/Y OR2X1_LOC_56/A 0.07fF
C19425 OR2X1_LOC_482/Y OR2X1_LOC_625/Y 0.21fF
C19426 AND2X1_LOC_733/Y OR2X1_LOC_59/Y 0.03fF
C19427 OR2X1_LOC_305/Y OR2X1_LOC_428/A 0.04fF
C19428 OR2X1_LOC_703/B AND2X1_LOC_534/a_8_24# 0.20fF
C19429 OR2X1_LOC_40/Y OR2X1_LOC_531/a_8_216# 0.15fF
C19430 VDD OR2X1_LOC_575/A 0.33fF
C19431 OR2X1_LOC_163/A OR2X1_LOC_163/a_8_216# 0.47fF
C19432 AND2X1_LOC_338/Y OR2X1_LOC_26/Y 0.06fF
C19433 OR2X1_LOC_335/a_36_216# OR2X1_LOC_787/Y 0.00fF
C19434 OR2X1_LOC_510/Y OR2X1_LOC_549/A 0.07fF
C19435 OR2X1_LOC_456/Y OR2X1_LOC_549/A 0.12fF
C19436 AND2X1_LOC_831/Y OR2X1_LOC_13/B 0.06fF
C19437 AND2X1_LOC_3/Y OR2X1_LOC_392/B 0.01fF
C19438 VDD AND2X1_LOC_841/B 0.51fF
C19439 AND2X1_LOC_17/Y AND2X1_LOC_425/a_36_24# 0.01fF
C19440 VDD OR2X1_LOC_493/A 0.02fF
C19441 OR2X1_LOC_379/a_8_216# OR2X1_LOC_648/B 0.40fF
C19442 OR2X1_LOC_833/a_36_216# AND2X1_LOC_92/Y 0.00fF
C19443 OR2X1_LOC_715/B OR2X1_LOC_375/A 0.03fF
C19444 AND2X1_LOC_43/B AND2X1_LOC_411/a_8_24# 0.05fF
C19445 OR2X1_LOC_653/Y AND2X1_LOC_172/a_36_24# 0.00fF
C19446 OR2X1_LOC_158/A AND2X1_LOC_576/Y 0.07fF
C19447 OR2X1_LOC_135/Y OR2X1_LOC_52/B 0.07fF
C19448 OR2X1_LOC_375/A OR2X1_LOC_543/A 0.01fF
C19449 AND2X1_LOC_91/B AND2X1_LOC_51/Y 1.08fF
C19450 OR2X1_LOC_604/A OR2X1_LOC_237/Y 0.03fF
C19451 OR2X1_LOC_703/B AND2X1_LOC_110/Y 0.01fF
C19452 OR2X1_LOC_117/a_8_216# OR2X1_LOC_3/Y 0.01fF
C19453 AND2X1_LOC_211/B OR2X1_LOC_12/Y 0.10fF
C19454 AND2X1_LOC_605/Y OR2X1_LOC_92/Y 0.02fF
C19455 AND2X1_LOC_716/Y AND2X1_LOC_335/a_8_24# 0.03fF
C19456 VDD OR2X1_LOC_652/a_8_216# 0.21fF
C19457 OR2X1_LOC_645/a_8_216# OR2X1_LOC_161/A 0.03fF
C19458 AND2X1_LOC_573/A AND2X1_LOC_404/B 0.91fF
C19459 OR2X1_LOC_85/A AND2X1_LOC_243/Y 0.04fF
C19460 OR2X1_LOC_45/B OR2X1_LOC_273/a_8_216# 0.01fF
C19461 OR2X1_LOC_287/B AND2X1_LOC_82/Y 1.06fF
C19462 OR2X1_LOC_810/A OR2X1_LOC_549/A 0.10fF
C19463 OR2X1_LOC_93/Y OR2X1_LOC_6/A 0.01fF
C19464 OR2X1_LOC_107/Y OR2X1_LOC_427/A 0.01fF
C19465 OR2X1_LOC_450/A AND2X1_LOC_695/a_36_24# 0.01fF
C19466 AND2X1_LOC_565/B OR2X1_LOC_189/A 0.00fF
C19467 OR2X1_LOC_516/A OR2X1_LOC_56/A 0.10fF
C19468 AND2X1_LOC_50/Y D_INPUT_4 0.36fF
C19469 AND2X1_LOC_8/Y OR2X1_LOC_786/A 0.02fF
C19470 AND2X1_LOC_3/Y OR2X1_LOC_113/B 0.03fF
C19471 OR2X1_LOC_325/A OR2X1_LOC_325/a_8_216# 0.02fF
C19472 OR2X1_LOC_235/B OR2X1_LOC_619/Y 0.07fF
C19473 AND2X1_LOC_675/A AND2X1_LOC_439/a_8_24# 0.01fF
C19474 AND2X1_LOC_722/A OR2X1_LOC_427/A 0.01fF
C19475 OR2X1_LOC_377/A AND2X1_LOC_377/Y 0.03fF
C19476 OR2X1_LOC_417/Y OR2X1_LOC_428/A 0.03fF
C19477 AND2X1_LOC_1/Y INPUT_7 0.01fF
C19478 AND2X1_LOC_41/A OR2X1_LOC_541/B 0.02fF
C19479 AND2X1_LOC_664/a_8_24# GATE_579 0.01fF
C19480 AND2X1_LOC_702/Y OR2X1_LOC_426/B 0.00fF
C19481 VDD AND2X1_LOC_187/a_8_24# 0.00fF
C19482 AND2X1_LOC_350/B AND2X1_LOC_350/Y 0.01fF
C19483 OR2X1_LOC_51/Y OR2X1_LOC_372/Y 0.06fF
C19484 INPUT_0 OR2X1_LOC_463/B 0.01fF
C19485 AND2X1_LOC_321/a_8_24# OR2X1_LOC_147/B 0.22fF
C19486 OR2X1_LOC_111/a_8_216# AND2X1_LOC_831/Y 0.01fF
C19487 AND2X1_LOC_570/Y OR2X1_LOC_497/Y 0.05fF
C19488 OR2X1_LOC_58/Y OR2X1_LOC_32/a_36_216# 0.00fF
C19489 OR2X1_LOC_311/Y OR2X1_LOC_428/A 0.06fF
C19490 OR2X1_LOC_108/a_36_216# OR2X1_LOC_529/Y 0.00fF
C19491 AND2X1_LOC_40/Y OR2X1_LOC_181/B 0.02fF
C19492 OR2X1_LOC_499/B AND2X1_LOC_43/B 0.03fF
C19493 OR2X1_LOC_822/Y OR2X1_LOC_585/A 0.02fF
C19494 OR2X1_LOC_837/Y OR2X1_LOC_39/A 0.07fF
C19495 OR2X1_LOC_604/A OR2X1_LOC_487/a_8_216# 0.30fF
C19496 OR2X1_LOC_533/A OR2X1_LOC_534/Y 0.19fF
C19497 OR2X1_LOC_49/A OR2X1_LOC_606/a_8_216# 0.11fF
C19498 OR2X1_LOC_519/Y AND2X1_LOC_716/Y 0.00fF
C19499 AND2X1_LOC_858/B OR2X1_LOC_36/Y 0.10fF
C19500 OR2X1_LOC_134/Y AND2X1_LOC_656/Y 0.03fF
C19501 AND2X1_LOC_725/a_8_24# OR2X1_LOC_743/A 0.01fF
C19502 AND2X1_LOC_303/A AND2X1_LOC_303/a_8_24# 0.01fF
C19503 OR2X1_LOC_653/B OR2X1_LOC_436/a_8_216# 0.47fF
C19504 OR2X1_LOC_154/A OR2X1_LOC_174/A 0.01fF
C19505 OR2X1_LOC_648/a_36_216# AND2X1_LOC_7/B 0.00fF
C19506 OR2X1_LOC_822/a_36_216# OR2X1_LOC_485/A 0.02fF
C19507 OR2X1_LOC_450/A AND2X1_LOC_3/Y 0.01fF
C19508 OR2X1_LOC_91/A OR2X1_LOC_36/Y 0.73fF
C19509 AND2X1_LOC_64/Y OR2X1_LOC_436/Y 0.03fF
C19510 AND2X1_LOC_862/a_8_24# OR2X1_LOC_59/Y 0.01fF
C19511 OR2X1_LOC_244/A OR2X1_LOC_267/Y 0.13fF
C19512 AND2X1_LOC_454/a_36_24# OR2X1_LOC_52/B 0.01fF
C19513 AND2X1_LOC_580/A AND2X1_LOC_861/B 0.07fF
C19514 OR2X1_LOC_45/B AND2X1_LOC_687/Y 0.01fF
C19515 AND2X1_LOC_76/Y AND2X1_LOC_520/Y 0.02fF
C19516 OR2X1_LOC_494/Y OR2X1_LOC_485/A 0.01fF
C19517 AND2X1_LOC_363/Y OR2X1_LOC_485/A 0.02fF
C19518 AND2X1_LOC_443/Y OR2X1_LOC_52/B 0.17fF
C19519 OR2X1_LOC_84/B OR2X1_LOC_78/A 0.00fF
C19520 AND2X1_LOC_12/Y OR2X1_LOC_653/Y 0.07fF
C19521 OR2X1_LOC_278/Y AND2X1_LOC_287/a_8_24# 0.01fF
C19522 OR2X1_LOC_494/A AND2X1_LOC_866/A 0.03fF
C19523 OR2X1_LOC_224/a_36_216# AND2X1_LOC_465/A 0.00fF
C19524 OR2X1_LOC_256/Y AND2X1_LOC_348/Y 0.03fF
C19525 OR2X1_LOC_732/a_8_216# OR2X1_LOC_732/B 0.04fF
C19526 AND2X1_LOC_578/A AND2X1_LOC_658/A 0.07fF
C19527 OR2X1_LOC_427/A AND2X1_LOC_454/Y 0.02fF
C19528 OR2X1_LOC_106/Y AND2X1_LOC_114/Y 0.00fF
C19529 OR2X1_LOC_609/A OR2X1_LOC_612/Y 0.00fF
C19530 OR2X1_LOC_755/A OR2X1_LOC_815/a_8_216# 0.02fF
C19531 OR2X1_LOC_264/Y OR2X1_LOC_216/Y 0.02fF
C19532 OR2X1_LOC_6/B OR2X1_LOC_121/B 0.03fF
C19533 OR2X1_LOC_244/A OR2X1_LOC_633/A 0.19fF
C19534 OR2X1_LOC_506/A OR2X1_LOC_447/a_8_216# 0.08fF
C19535 OR2X1_LOC_70/Y AND2X1_LOC_657/Y 0.12fF
C19536 AND2X1_LOC_72/a_36_24# OR2X1_LOC_78/A 0.00fF
C19537 AND2X1_LOC_191/B AND2X1_LOC_711/Y 0.00fF
C19538 OR2X1_LOC_405/A OR2X1_LOC_405/Y 0.14fF
C19539 AND2X1_LOC_228/Y OR2X1_LOC_48/B 0.03fF
C19540 OR2X1_LOC_838/a_8_216# AND2X1_LOC_472/B 0.06fF
C19541 OR2X1_LOC_256/Y OR2X1_LOC_753/A 0.01fF
C19542 OR2X1_LOC_114/Y OR2X1_LOC_574/a_36_216# 0.00fF
C19543 OR2X1_LOC_756/B OR2X1_LOC_564/A 0.04fF
C19544 AND2X1_LOC_727/Y AND2X1_LOC_808/A 0.03fF
C19545 AND2X1_LOC_530/a_8_24# OR2X1_LOC_532/B 0.01fF
C19546 VDD OR2X1_LOC_456/A -0.00fF
C19547 AND2X1_LOC_141/B OR2X1_LOC_56/A 0.18fF
C19548 OR2X1_LOC_402/B OR2X1_LOC_402/a_36_216# 0.01fF
C19549 OR2X1_LOC_92/Y AND2X1_LOC_361/A 0.10fF
C19550 OR2X1_LOC_645/a_8_216# AND2X1_LOC_51/Y 0.02fF
C19551 OR2X1_LOC_160/A OR2X1_LOC_128/B 0.02fF
C19552 OR2X1_LOC_70/Y AND2X1_LOC_469/B 0.03fF
C19553 AND2X1_LOC_228/Y OR2X1_LOC_18/Y 0.04fF
C19554 AND2X1_LOC_215/Y OR2X1_LOC_291/Y 0.54fF
C19555 OR2X1_LOC_341/Y OR2X1_LOC_340/Y 0.06fF
C19556 OR2X1_LOC_472/A OR2X1_LOC_640/A 0.11fF
C19557 INPUT_1 AND2X1_LOC_476/Y 0.01fF
C19558 OR2X1_LOC_235/a_8_216# OR2X1_LOC_278/Y 0.01fF
C19559 D_INPUT_3 OR2X1_LOC_428/A 0.03fF
C19560 OR2X1_LOC_506/A OR2X1_LOC_130/A 0.11fF
C19561 AND2X1_LOC_27/a_8_24# OR2X1_LOC_66/A 0.11fF
C19562 OR2X1_LOC_459/B OR2X1_LOC_459/a_8_216# 0.02fF
C19563 OR2X1_LOC_103/a_8_216# AND2X1_LOC_576/Y 0.01fF
C19564 OR2X1_LOC_599/A OR2X1_LOC_427/A 0.08fF
C19565 OR2X1_LOC_624/B OR2X1_LOC_624/a_8_216# 0.01fF
C19566 AND2X1_LOC_12/Y OR2X1_LOC_848/B 0.28fF
C19567 AND2X1_LOC_726/a_36_24# OR2X1_LOC_47/Y 0.00fF
C19568 AND2X1_LOC_539/Y OR2X1_LOC_599/Y 0.03fF
C19569 AND2X1_LOC_554/B OR2X1_LOC_517/A 0.02fF
C19570 OR2X1_LOC_100/Y AND2X1_LOC_3/Y 0.00fF
C19571 OR2X1_LOC_3/Y AND2X1_LOC_141/A 0.11fF
C19572 D_INPUT_3 OR2X1_LOC_595/A 0.02fF
C19573 AND2X1_LOC_733/Y OR2X1_LOC_70/Y 0.03fF
C19574 OR2X1_LOC_811/a_8_216# OR2X1_LOC_269/B 0.02fF
C19575 OR2X1_LOC_377/A OR2X1_LOC_793/A 0.07fF
C19576 OR2X1_LOC_491/a_8_216# OR2X1_LOC_31/Y 0.08fF
C19577 OR2X1_LOC_36/Y AND2X1_LOC_573/A 0.14fF
C19578 AND2X1_LOC_817/B OR2X1_LOC_847/a_36_216# 0.00fF
C19579 OR2X1_LOC_359/a_8_216# OR2X1_LOC_814/A 0.01fF
C19580 OR2X1_LOC_440/A OR2X1_LOC_439/B 0.50fF
C19581 AND2X1_LOC_520/Y OR2X1_LOC_52/B 0.01fF
C19582 OR2X1_LOC_448/A AND2X1_LOC_697/a_8_24# 0.20fF
C19583 AND2X1_LOC_514/Y AND2X1_LOC_469/B 0.09fF
C19584 OR2X1_LOC_585/A OR2X1_LOC_48/B 0.10fF
C19585 AND2X1_LOC_737/a_36_24# OR2X1_LOC_74/A 0.01fF
C19586 AND2X1_LOC_271/a_36_24# AND2X1_LOC_7/B 0.00fF
C19587 OR2X1_LOC_54/Y OR2X1_LOC_56/A 0.29fF
C19588 OR2X1_LOC_864/A OR2X1_LOC_185/A 0.03fF
C19589 OR2X1_LOC_158/A AND2X1_LOC_472/a_8_24# 0.05fF
C19590 OR2X1_LOC_188/Y AND2X1_LOC_237/a_36_24# 0.00fF
C19591 AND2X1_LOC_657/a_8_24# AND2X1_LOC_657/Y 0.01fF
C19592 AND2X1_LOC_324/a_8_24# AND2X1_LOC_857/Y 0.01fF
C19593 OR2X1_LOC_744/A AND2X1_LOC_727/A 0.03fF
C19594 OR2X1_LOC_434/A AND2X1_LOC_18/Y 0.52fF
C19595 OR2X1_LOC_65/B AND2X1_LOC_361/A 0.25fF
C19596 OR2X1_LOC_18/Y OR2X1_LOC_585/A 0.10fF
C19597 AND2X1_LOC_175/B OR2X1_LOC_52/B 0.00fF
C19598 OR2X1_LOC_271/Y AND2X1_LOC_318/a_8_24# 0.23fF
C19599 OR2X1_LOC_329/B AND2X1_LOC_465/Y 0.02fF
C19600 OR2X1_LOC_800/A OR2X1_LOC_800/a_8_216# 0.47fF
C19601 OR2X1_LOC_803/B OR2X1_LOC_155/A 0.01fF
C19602 OR2X1_LOC_185/A OR2X1_LOC_633/B 0.03fF
C19603 OR2X1_LOC_76/A OR2X1_LOC_464/A 0.03fF
C19604 AND2X1_LOC_81/a_8_24# OR2X1_LOC_375/A 0.01fF
C19605 AND2X1_LOC_342/a_8_24# OR2X1_LOC_85/A 0.02fF
C19606 AND2X1_LOC_753/B OR2X1_LOC_193/A 0.02fF
C19607 OR2X1_LOC_312/Y AND2X1_LOC_436/B 1.06fF
C19608 OR2X1_LOC_517/a_8_216# OR2X1_LOC_22/Y 0.01fF
C19609 AND2X1_LOC_707/a_8_24# OR2X1_LOC_31/Y 0.01fF
C19610 OR2X1_LOC_46/A AND2X1_LOC_222/a_36_24# 0.00fF
C19611 AND2X1_LOC_749/a_8_24# OR2X1_LOC_476/B 0.02fF
C19612 OR2X1_LOC_216/Y OR2X1_LOC_643/A 0.48fF
C19613 OR2X1_LOC_175/Y OR2X1_LOC_170/Y 0.09fF
C19614 OR2X1_LOC_490/Y OR2X1_LOC_118/Y 0.03fF
C19615 OR2X1_LOC_74/A OR2X1_LOC_118/Y 0.03fF
C19616 OR2X1_LOC_217/Y OR2X1_LOC_217/a_8_216# 0.01fF
C19617 AND2X1_LOC_154/a_36_24# OR2X1_LOC_52/B 0.00fF
C19618 OR2X1_LOC_756/B AND2X1_LOC_165/a_8_24# 0.01fF
C19619 AND2X1_LOC_96/a_8_24# INPUT_1 0.01fF
C19620 OR2X1_LOC_235/B OR2X1_LOC_720/B 0.79fF
C19621 OR2X1_LOC_481/a_8_216# AND2X1_LOC_847/Y 0.03fF
C19622 AND2X1_LOC_56/B OR2X1_LOC_552/a_8_216# 0.01fF
C19623 OR2X1_LOC_680/Y AND2X1_LOC_624/A 0.03fF
C19624 AND2X1_LOC_95/Y OR2X1_LOC_35/B 0.01fF
C19625 AND2X1_LOC_35/Y OR2X1_LOC_24/Y 0.00fF
C19626 OR2X1_LOC_685/A AND2X1_LOC_3/Y 0.01fF
C19627 OR2X1_LOC_326/B OR2X1_LOC_121/B 0.02fF
C19628 OR2X1_LOC_272/Y OR2X1_LOC_39/A 0.02fF
C19629 OR2X1_LOC_19/B OR2X1_LOC_23/a_8_216# -0.04fF
C19630 OR2X1_LOC_744/A OR2X1_LOC_95/Y 0.40fF
C19631 OR2X1_LOC_589/A AND2X1_LOC_644/a_8_24# 0.04fF
C19632 OR2X1_LOC_805/A OR2X1_LOC_216/a_36_216# 0.02fF
C19633 AND2X1_LOC_211/B AND2X1_LOC_650/Y 0.01fF
C19634 OR2X1_LOC_799/A AND2X1_LOC_51/Y 0.22fF
C19635 OR2X1_LOC_551/B OR2X1_LOC_364/a_8_216# 0.40fF
C19636 AND2X1_LOC_44/Y OR2X1_LOC_779/B 0.79fF
C19637 OR2X1_LOC_22/Y OR2X1_LOC_59/a_8_216# 0.01fF
C19638 AND2X1_LOC_656/a_8_24# OR2X1_LOC_595/A 0.01fF
C19639 AND2X1_LOC_792/B AND2X1_LOC_789/Y 0.03fF
C19640 OR2X1_LOC_600/A AND2X1_LOC_721/A 0.03fF
C19641 OR2X1_LOC_659/A AND2X1_LOC_47/Y 0.10fF
C19642 AND2X1_LOC_702/Y OR2X1_LOC_743/A 0.03fF
C19643 OR2X1_LOC_145/Y AND2X1_LOC_148/a_8_24# 0.23fF
C19644 OR2X1_LOC_183/a_8_216# OR2X1_LOC_183/Y 0.01fF
C19645 AND2X1_LOC_191/B OR2X1_LOC_184/Y 0.11fF
C19646 AND2X1_LOC_175/a_8_24# AND2X1_LOC_211/B 0.01fF
C19647 OR2X1_LOC_610/Y OR2X1_LOC_647/B 0.04fF
C19648 OR2X1_LOC_385/Y OR2X1_LOC_585/A 0.47fF
C19649 OR2X1_LOC_131/Y OR2X1_LOC_43/A 0.12fF
C19650 OR2X1_LOC_625/Y OR2X1_LOC_628/Y 0.11fF
C19651 OR2X1_LOC_185/Y AND2X1_LOC_67/Y 0.17fF
C19652 OR2X1_LOC_800/Y OR2X1_LOC_801/B 0.06fF
C19653 OR2X1_LOC_80/A OR2X1_LOC_548/a_8_216# 0.05fF
C19654 AND2X1_LOC_632/A AND2X1_LOC_805/Y 0.03fF
C19655 AND2X1_LOC_862/a_36_24# OR2X1_LOC_74/A 0.01fF
C19656 OR2X1_LOC_405/A D_INPUT_0 0.05fF
C19657 INPUT_5 OR2X1_LOC_587/a_8_216# 0.01fF
C19658 OR2X1_LOC_64/Y AND2X1_LOC_661/A 0.03fF
C19659 OR2X1_LOC_593/B OR2X1_LOC_718/a_8_216# 0.01fF
C19660 OR2X1_LOC_647/Y OR2X1_LOC_99/Y 0.00fF
C19661 AND2X1_LOC_519/a_8_24# OR2X1_LOC_375/A 0.03fF
C19662 AND2X1_LOC_849/A OR2X1_LOC_44/Y 0.02fF
C19663 OR2X1_LOC_838/a_8_216# OR2X1_LOC_838/B 0.05fF
C19664 AND2X1_LOC_1/Y AND2X1_LOC_51/A 0.01fF
C19665 OR2X1_LOC_369/a_8_216# AND2X1_LOC_222/Y 0.01fF
C19666 OR2X1_LOC_3/Y AND2X1_LOC_42/B 0.08fF
C19667 AND2X1_LOC_727/A AND2X1_LOC_840/B 0.05fF
C19668 AND2X1_LOC_866/A OR2X1_LOC_427/A 0.17fF
C19669 AND2X1_LOC_56/B OR2X1_LOC_54/Y 0.18fF
C19670 OR2X1_LOC_440/A OR2X1_LOC_733/a_36_216# 0.01fF
C19671 OR2X1_LOC_600/A OR2X1_LOC_331/Y 0.07fF
C19672 OR2X1_LOC_3/Y AND2X1_LOC_651/B 0.01fF
C19673 AND2X1_LOC_733/Y OR2X1_LOC_437/Y 0.15fF
C19674 AND2X1_LOC_170/B OR2X1_LOC_619/Y 0.07fF
C19675 OR2X1_LOC_807/A OR2X1_LOC_286/B 0.01fF
C19676 OR2X1_LOC_776/Y OR2X1_LOC_228/Y 0.01fF
C19677 AND2X1_LOC_702/Y OR2X1_LOC_246/A 0.00fF
C19678 AND2X1_LOC_486/Y OR2X1_LOC_615/Y 0.01fF
C19679 OR2X1_LOC_128/A AND2X1_LOC_47/Y 0.04fF
C19680 AND2X1_LOC_848/A OR2X1_LOC_59/Y 0.05fF
C19681 OR2X1_LOC_709/A OR2X1_LOC_317/B 0.08fF
C19682 AND2X1_LOC_138/a_8_24# OR2X1_LOC_417/A 0.02fF
C19683 AND2X1_LOC_8/Y OR2X1_LOC_54/Y 0.07fF
C19684 AND2X1_LOC_645/a_8_24# OR2X1_LOC_48/B 0.02fF
C19685 OR2X1_LOC_166/a_8_216# OR2X1_LOC_331/Y 0.01fF
C19686 OR2X1_LOC_218/Y OR2X1_LOC_805/A 0.09fF
C19687 AND2X1_LOC_7/B OR2X1_LOC_703/Y 0.00fF
C19688 OR2X1_LOC_102/a_36_216# OR2X1_LOC_13/B 0.00fF
C19689 OR2X1_LOC_12/Y AND2X1_LOC_247/a_36_24# 0.00fF
C19690 OR2X1_LOC_647/A OR2X1_LOC_647/a_8_216# 0.08fF
C19691 OR2X1_LOC_59/Y AND2X1_LOC_203/a_8_24# 0.01fF
C19692 OR2X1_LOC_139/A OR2X1_LOC_508/Y 0.36fF
C19693 OR2X1_LOC_175/Y OR2X1_LOC_168/Y 0.01fF
C19694 AND2X1_LOC_840/B OR2X1_LOC_95/Y 0.12fF
C19695 AND2X1_LOC_31/Y OR2X1_LOC_778/a_36_216# 0.00fF
C19696 AND2X1_LOC_640/Y OR2X1_LOC_46/A 0.06fF
C19697 OR2X1_LOC_715/B OR2X1_LOC_515/Y 0.01fF
C19698 OR2X1_LOC_59/Y AND2X1_LOC_206/Y 0.51fF
C19699 OR2X1_LOC_291/A OR2X1_LOC_54/Y 0.11fF
C19700 AND2X1_LOC_108/a_8_24# OR2X1_LOC_346/B 0.01fF
C19701 OR2X1_LOC_130/A OR2X1_LOC_227/Y -0.00fF
C19702 AND2X1_LOC_729/B OR2X1_LOC_43/a_36_216# 0.00fF
C19703 AND2X1_LOC_47/Y OR2X1_LOC_449/B 0.11fF
C19704 OR2X1_LOC_31/Y OR2X1_LOC_591/a_8_216# 0.01fF
C19705 OR2X1_LOC_112/a_8_216# OR2X1_LOC_175/a_8_216# 0.47fF
C19706 OR2X1_LOC_26/Y AND2X1_LOC_859/B 0.02fF
C19707 AND2X1_LOC_514/Y OR2X1_LOC_417/a_36_216# 0.01fF
C19708 OR2X1_LOC_532/B AND2X1_LOC_3/Y 0.17fF
C19709 OR2X1_LOC_532/B OR2X1_LOC_647/B 0.02fF
C19710 OR2X1_LOC_45/B OR2X1_LOC_110/a_8_216# 0.01fF
C19711 OR2X1_LOC_737/A OR2X1_LOC_723/A 0.04fF
C19712 AND2X1_LOC_7/B OR2X1_LOC_120/a_8_216# 0.01fF
C19713 OR2X1_LOC_158/A AND2X1_LOC_793/a_8_24# 0.08fF
C19714 AND2X1_LOC_665/a_8_24# AND2X1_LOC_3/Y 0.04fF
C19715 VDD OR2X1_LOC_332/a_8_216# 0.00fF
C19716 AND2X1_LOC_748/a_36_24# OR2X1_LOC_801/B 0.01fF
C19717 OR2X1_LOC_66/A OR2X1_LOC_712/B 0.00fF
C19718 OR2X1_LOC_118/Y AND2X1_LOC_647/Y 0.02fF
C19719 OR2X1_LOC_832/a_8_216# OR2X1_LOC_593/B 0.14fF
C19720 OR2X1_LOC_516/Y AND2X1_LOC_477/Y 0.00fF
C19721 OR2X1_LOC_176/Y AND2X1_LOC_799/a_8_24# 0.11fF
C19722 AND2X1_LOC_600/a_36_24# AND2X1_LOC_51/Y 0.00fF
C19723 OR2X1_LOC_619/Y OR2X1_LOC_331/Y 0.07fF
C19724 AND2X1_LOC_773/Y OR2X1_LOC_136/Y 0.02fF
C19725 OR2X1_LOC_572/a_8_216# OR2X1_LOC_576/A 0.01fF
C19726 OR2X1_LOC_49/A AND2X1_LOC_7/B 0.07fF
C19727 AND2X1_LOC_8/Y OR2X1_LOC_84/Y 0.27fF
C19728 AND2X1_LOC_42/B OR2X1_LOC_673/A 0.02fF
C19729 OR2X1_LOC_43/A AND2X1_LOC_644/a_8_24# 0.02fF
C19730 OR2X1_LOC_121/B AND2X1_LOC_47/Y 0.25fF
C19731 OR2X1_LOC_555/B OR2X1_LOC_345/a_8_216# 0.02fF
C19732 OR2X1_LOC_64/Y AND2X1_LOC_810/Y 0.09fF
C19733 OR2X1_LOC_97/A OR2X1_LOC_486/Y 0.03fF
C19734 OR2X1_LOC_709/A AND2X1_LOC_44/Y 0.46fF
C19735 AND2X1_LOC_7/B OR2X1_LOC_596/A 0.07fF
C19736 OR2X1_LOC_64/Y OR2X1_LOC_760/Y 0.06fF
C19737 OR2X1_LOC_585/A AND2X1_LOC_228/a_36_24# 0.01fF
C19738 AND2X1_LOC_64/Y OR2X1_LOC_160/B 0.18fF
C19739 AND2X1_LOC_295/a_8_24# AND2X1_LOC_44/Y 0.01fF
C19740 OR2X1_LOC_78/Y AND2X1_LOC_36/Y 0.11fF
C19741 OR2X1_LOC_485/A OR2X1_LOC_311/a_8_216# 0.01fF
C19742 OR2X1_LOC_47/Y AND2X1_LOC_523/Y 0.03fF
C19743 OR2X1_LOC_833/Y AND2X1_LOC_255/a_8_24# 0.17fF
C19744 OR2X1_LOC_728/B OR2X1_LOC_155/A 0.00fF
C19745 AND2X1_LOC_543/Y VDD 0.10fF
C19746 OR2X1_LOC_158/A AND2X1_LOC_244/A 0.05fF
C19747 OR2X1_LOC_494/A OR2X1_LOC_40/Y 0.01fF
C19748 OR2X1_LOC_70/A AND2X1_LOC_638/a_8_24# 0.01fF
C19749 OR2X1_LOC_161/A OR2X1_LOC_446/B 1.34fF
C19750 AND2X1_LOC_22/Y OR2X1_LOC_307/A 0.28fF
C19751 AND2X1_LOC_28/a_36_24# D_INPUT_0 0.00fF
C19752 OR2X1_LOC_161/A OR2X1_LOC_303/B 0.06fF
C19753 OR2X1_LOC_780/A OR2X1_LOC_780/B 0.04fF
C19754 OR2X1_LOC_709/A OR2X1_LOC_514/a_8_216# 0.01fF
C19755 OR2X1_LOC_730/a_8_216# OR2X1_LOC_730/B 0.01fF
C19756 OR2X1_LOC_319/B OR2X1_LOC_703/Y 0.01fF
C19757 AND2X1_LOC_540/a_8_24# OR2X1_LOC_183/Y 0.04fF
C19758 OR2X1_LOC_158/A OR2X1_LOC_16/A 0.14fF
C19759 AND2X1_LOC_711/Y AND2X1_LOC_848/A 0.08fF
C19760 AND2X1_LOC_31/Y OR2X1_LOC_722/a_36_216# 0.00fF
C19761 OR2X1_LOC_651/A OR2X1_LOC_228/a_8_216# 0.03fF
C19762 OR2X1_LOC_139/A OR2X1_LOC_66/A 0.05fF
C19763 AND2X1_LOC_436/B OR2X1_LOC_13/B -0.01fF
C19764 OR2X1_LOC_31/Y OR2X1_LOC_95/Y 0.15fF
C19765 AND2X1_LOC_231/Y VDD 0.06fF
C19766 OR2X1_LOC_62/B D_INPUT_1 0.11fF
C19767 D_GATE_479 VDD 0.11fF
C19768 OR2X1_LOC_31/Y OR2X1_LOC_368/A 0.11fF
C19769 OR2X1_LOC_724/a_8_216# AND2X1_LOC_36/Y 0.01fF
C19770 OR2X1_LOC_151/A OR2X1_LOC_361/a_8_216# 0.02fF
C19771 OR2X1_LOC_92/Y OR2X1_LOC_387/A 0.00fF
C19772 OR2X1_LOC_402/Y OR2X1_LOC_771/B 0.07fF
C19773 OR2X1_LOC_715/B OR2X1_LOC_549/A 0.31fF
C19774 OR2X1_LOC_702/A AND2X1_LOC_31/Y 0.05fF
C19775 VDD OR2X1_LOC_161/B 2.21fF
C19776 AND2X1_LOC_626/a_8_24# OR2X1_LOC_549/A 0.02fF
C19777 OR2X1_LOC_754/A AND2X1_LOC_562/Y 0.03fF
C19778 OR2X1_LOC_3/Y AND2X1_LOC_793/B 0.03fF
C19779 AND2X1_LOC_70/Y AND2X1_LOC_44/Y 1.74fF
C19780 OR2X1_LOC_505/a_36_216# AND2X1_LOC_508/B 0.00fF
C19781 VDD OR2X1_LOC_562/B -0.00fF
C19782 OR2X1_LOC_19/B OR2X1_LOC_801/B 0.02fF
C19783 OR2X1_LOC_756/B OR2X1_LOC_562/A 0.14fF
C19784 OR2X1_LOC_532/B OR2X1_LOC_270/Y 0.03fF
C19785 AND2X1_LOC_544/Y OR2X1_LOC_441/a_8_216# 0.03fF
C19786 OR2X1_LOC_788/a_8_216# OR2X1_LOC_605/Y 0.01fF
C19787 AND2X1_LOC_476/Y AND2X1_LOC_778/Y 0.07fF
C19788 OR2X1_LOC_1/a_8_216# INPUT_6 0.07fF
C19789 OR2X1_LOC_158/A OR2X1_LOC_108/Y 0.17fF
C19790 OR2X1_LOC_464/A OR2X1_LOC_722/B 0.04fF
C19791 OR2X1_LOC_415/a_36_216# OR2X1_LOC_598/A 0.03fF
C19792 OR2X1_LOC_269/B OR2X1_LOC_561/A 0.01fF
C19793 OR2X1_LOC_7/A AND2X1_LOC_212/a_8_24# 0.02fF
C19794 VDD OR2X1_LOC_589/A 0.85fF
C19795 AND2X1_LOC_92/Y OR2X1_LOC_389/a_8_216# 0.06fF
C19796 AND2X1_LOC_64/Y OR2X1_LOC_475/a_36_216# 0.02fF
C19797 OR2X1_LOC_287/B OR2X1_LOC_579/a_8_216# 0.01fF
C19798 OR2X1_LOC_865/A OR2X1_LOC_859/a_8_216# 0.01fF
C19799 VDD OR2X1_LOC_322/Y 0.49fF
C19800 AND2X1_LOC_325/a_8_24# AND2X1_LOC_476/Y 0.06fF
C19801 OR2X1_LOC_39/A OR2X1_LOC_504/a_36_216# 0.00fF
C19802 OR2X1_LOC_186/Y OR2X1_LOC_78/A 0.03fF
C19803 OR2X1_LOC_696/A INPUT_3 0.01fF
C19804 OR2X1_LOC_476/B AND2X1_LOC_31/Y 0.01fF
C19805 OR2X1_LOC_227/Y AND2X1_LOC_88/Y 0.06fF
C19806 OR2X1_LOC_703/A AND2X1_LOC_44/Y 0.00fF
C19807 OR2X1_LOC_302/B OR2X1_LOC_486/Y 0.03fF
C19808 AND2X1_LOC_474/A OR2X1_LOC_12/Y 2.23fF
C19809 AND2X1_LOC_86/Y AND2X1_LOC_64/Y 0.11fF
C19810 AND2X1_LOC_486/Y AND2X1_LOC_242/B 0.03fF
C19811 OR2X1_LOC_860/Y OR2X1_LOC_392/B 0.10fF
C19812 OR2X1_LOC_750/A OR2X1_LOC_68/B 0.04fF
C19813 AND2X1_LOC_571/A AND2X1_LOC_572/Y 0.20fF
C19814 OR2X1_LOC_671/Y INPUT_0 0.05fF
C19815 AND2X1_LOC_477/a_8_24# AND2X1_LOC_212/Y 0.01fF
C19816 OR2X1_LOC_435/a_8_216# OR2X1_LOC_435/A 0.08fF
C19817 AND2X1_LOC_51/Y OR2X1_LOC_446/B 0.06fF
C19818 OR2X1_LOC_46/A OR2X1_LOC_80/A 0.56fF
C19819 OR2X1_LOC_748/A OR2X1_LOC_759/Y 0.01fF
C19820 AND2X1_LOC_564/B OR2X1_LOC_18/Y 0.19fF
C19821 OR2X1_LOC_404/Y OR2X1_LOC_501/a_8_216# 0.02fF
C19822 AND2X1_LOC_568/B OR2X1_LOC_51/Y 0.03fF
C19823 AND2X1_LOC_64/Y OR2X1_LOC_799/a_8_216# 0.02fF
C19824 OR2X1_LOC_732/a_8_216# AND2X1_LOC_7/B 0.01fF
C19825 OR2X1_LOC_18/Y OR2X1_LOC_230/Y 0.07fF
C19826 AND2X1_LOC_658/B AND2X1_LOC_657/Y 0.44fF
C19827 AND2X1_LOC_51/Y OR2X1_LOC_728/a_8_216# 0.02fF
C19828 OR2X1_LOC_604/A OR2X1_LOC_91/A 0.23fF
C19829 OR2X1_LOC_337/a_8_216# OR2X1_LOC_182/B 0.01fF
C19830 AND2X1_LOC_658/B AND2X1_LOC_469/B 0.03fF
C19831 OR2X1_LOC_747/Y AND2X1_LOC_781/Y 0.09fF
C19832 AND2X1_LOC_663/A OR2X1_LOC_627/Y 0.27fF
C19833 AND2X1_LOC_48/A OR2X1_LOC_193/a_36_216# 0.00fF
C19834 OR2X1_LOC_177/a_8_216# OR2X1_LOC_427/A 0.01fF
C19835 AND2X1_LOC_500/Y AND2X1_LOC_663/A 0.03fF
C19836 OR2X1_LOC_676/Y OR2X1_LOC_678/Y 0.14fF
C19837 OR2X1_LOC_744/a_36_216# OR2X1_LOC_39/A 0.00fF
C19838 OR2X1_LOC_154/A OR2X1_LOC_563/A 0.01fF
C19839 OR2X1_LOC_574/a_8_216# OR2X1_LOC_362/A 0.40fF
C19840 AND2X1_LOC_35/Y AND2X1_LOC_208/Y 0.01fF
C19841 VDD OR2X1_LOC_275/Y 0.00fF
C19842 OR2X1_LOC_160/B OR2X1_LOC_464/A 0.03fF
C19843 OR2X1_LOC_471/Y OR2X1_LOC_546/a_8_216# 0.10fF
C19844 VDD AND2X1_LOC_48/a_8_24# -0.00fF
C19845 OR2X1_LOC_604/A OR2X1_LOC_746/a_36_216# 0.00fF
C19846 OR2X1_LOC_87/B AND2X1_LOC_7/B 0.03fF
C19847 AND2X1_LOC_721/Y AND2X1_LOC_576/Y 0.02fF
C19848 OR2X1_LOC_512/A OR2X1_LOC_160/B 0.18fF
C19849 OR2X1_LOC_523/B AND2X1_LOC_95/Y 0.01fF
C19850 OR2X1_LOC_244/a_8_216# OR2X1_LOC_66/A 0.14fF
C19851 OR2X1_LOC_589/A OR2X1_LOC_829/a_8_216# 0.05fF
C19852 OR2X1_LOC_850/B OR2X1_LOC_66/A 0.00fF
C19853 OR2X1_LOC_834/A OR2X1_LOC_678/Y 0.00fF
C19854 OR2X1_LOC_684/a_8_216# OR2X1_LOC_426/A 0.01fF
C19855 OR2X1_LOC_64/Y AND2X1_LOC_204/a_8_24# 0.01fF
C19856 AND2X1_LOC_491/a_8_24# AND2X1_LOC_36/Y 0.03fF
C19857 VDD AND2X1_LOC_866/B 0.39fF
C19858 OR2X1_LOC_629/A OR2X1_LOC_140/B 0.21fF
C19859 OR2X1_LOC_122/Y OR2X1_LOC_744/A 0.06fF
C19860 VDD AND2X1_LOC_654/B 0.24fF
C19861 AND2X1_LOC_214/A INPUT_0 0.01fF
C19862 INPUT_0 AND2X1_LOC_529/a_8_24# 0.02fF
C19863 OR2X1_LOC_47/Y AND2X1_LOC_790/a_36_24# 0.00fF
C19864 OR2X1_LOC_40/Y OR2X1_LOC_427/A 0.11fF
C19865 AND2X1_LOC_354/a_8_24# AND2X1_LOC_810/B 0.02fF
C19866 AND2X1_LOC_354/a_36_24# AND2X1_LOC_802/Y 0.01fF
C19867 VDD OR2X1_LOC_495/Y 0.26fF
C19868 OR2X1_LOC_643/A OR2X1_LOC_576/A 0.06fF
C19869 AND2X1_LOC_86/Y AND2X1_LOC_86/a_8_24# 0.01fF
C19870 OR2X1_LOC_857/B AND2X1_LOC_824/B 0.21fF
C19871 VDD OR2X1_LOC_61/Y 0.23fF
C19872 OR2X1_LOC_44/Y OR2X1_LOC_759/a_8_216# 0.01fF
C19873 OR2X1_LOC_85/A OR2X1_LOC_12/Y 0.00fF
C19874 OR2X1_LOC_287/B OR2X1_LOC_362/a_8_216# 0.01fF
C19875 OR2X1_LOC_315/Y OR2X1_LOC_322/Y 0.02fF
C19876 OR2X1_LOC_124/Y OR2X1_LOC_576/A 0.00fF
C19877 OR2X1_LOC_494/A OR2X1_LOC_7/A 0.01fF
C19878 AND2X1_LOC_624/A AND2X1_LOC_476/Y 0.07fF
C19879 AND2X1_LOC_366/A AND2X1_LOC_456/B 0.03fF
C19880 OR2X1_LOC_179/Y OR2X1_LOC_744/A 0.01fF
C19881 OR2X1_LOC_168/B OR2X1_LOC_776/a_8_216# 0.01fF
C19882 OR2X1_LOC_53/Y OR2X1_LOC_485/A 0.02fF
C19883 AND2X1_LOC_17/Y AND2X1_LOC_44/Y 0.75fF
C19884 VDD AND2X1_LOC_398/a_8_24# -0.00fF
C19885 OR2X1_LOC_160/A OR2X1_LOC_730/A 0.02fF
C19886 AND2X1_LOC_340/a_8_24# OR2X1_LOC_118/Y 0.01fF
C19887 OR2X1_LOC_859/a_8_216# OR2X1_LOC_391/A 0.02fF
C19888 OR2X1_LOC_604/A AND2X1_LOC_573/A 0.10fF
C19889 AND2X1_LOC_47/Y OR2X1_LOC_195/a_8_216# 0.01fF
C19890 OR2X1_LOC_529/a_36_216# OR2X1_LOC_600/A 0.02fF
C19891 OR2X1_LOC_507/a_8_216# AND2X1_LOC_41/A 0.01fF
C19892 OR2X1_LOC_147/a_36_216# AND2X1_LOC_51/Y 0.00fF
C19893 OR2X1_LOC_33/B AND2X1_LOC_7/B 0.01fF
C19894 OR2X1_LOC_589/A AND2X1_LOC_267/a_8_24# 0.01fF
C19895 OR2X1_LOC_468/A OR2X1_LOC_506/A 0.03fF
C19896 OR2X1_LOC_224/Y OR2X1_LOC_437/A 0.08fF
C19897 OR2X1_LOC_375/A OR2X1_LOC_552/B 0.01fF
C19898 AND2X1_LOC_848/Y AND2X1_LOC_244/a_8_24# 0.01fF
C19899 OR2X1_LOC_158/A AND2X1_LOC_559/a_8_24# 0.03fF
C19900 OR2X1_LOC_744/A AND2X1_LOC_832/a_8_24# 0.02fF
C19901 OR2X1_LOC_866/B OR2X1_LOC_846/B 0.02fF
C19902 OR2X1_LOC_186/Y OR2X1_LOC_155/A 0.03fF
C19903 OR2X1_LOC_264/Y AND2X1_LOC_41/A 0.17fF
C19904 OR2X1_LOC_542/B OR2X1_LOC_161/A 0.03fF
C19905 VDD OR2X1_LOC_846/a_8_216# 0.00fF
C19906 AND2X1_LOC_576/Y OR2X1_LOC_482/Y 0.07fF
C19907 OR2X1_LOC_778/A OR2X1_LOC_563/A 0.14fF
C19908 OR2X1_LOC_84/a_36_216# OR2X1_LOC_71/A 0.00fF
C19909 VDD AND2X1_LOC_365/A 0.24fF
C19910 AND2X1_LOC_81/a_8_24# OR2X1_LOC_549/A 0.02fF
C19911 VDD OR2X1_LOC_87/a_8_216# 0.21fF
C19912 AND2X1_LOC_555/a_8_24# OR2X1_LOC_748/A 0.02fF
C19913 INPUT_0 AND2X1_LOC_820/a_8_24# 0.01fF
C19914 OR2X1_LOC_656/B OR2X1_LOC_78/B 0.10fF
C19915 AND2X1_LOC_850/a_8_24# AND2X1_LOC_858/B 0.03fF
C19916 VDD AND2X1_LOC_379/a_8_24# 0.00fF
C19917 OR2X1_LOC_624/A AND2X1_LOC_92/Y 0.10fF
C19918 OR2X1_LOC_493/a_36_216# OR2X1_LOC_805/A 0.01fF
C19919 VDD OR2X1_LOC_460/Y 0.00fF
C19920 AND2X1_LOC_73/a_36_24# OR2X1_LOC_185/A 0.00fF
C19921 AND2X1_LOC_767/a_8_24# OR2X1_LOC_78/B 0.01fF
C19922 OR2X1_LOC_40/Y AND2X1_LOC_363/A 0.17fF
C19923 AND2X1_LOC_753/B AND2X1_LOC_40/Y 0.07fF
C19924 AND2X1_LOC_724/Y OR2X1_LOC_36/Y 0.03fF
C19925 OR2X1_LOC_45/B OR2X1_LOC_277/a_8_216# 0.01fF
C19926 AND2X1_LOC_56/B OR2X1_LOC_190/Y 0.09fF
C19927 AND2X1_LOC_340/a_8_24# OR2X1_LOC_262/Y 0.02fF
C19928 AND2X1_LOC_605/Y OR2X1_LOC_619/Y 0.03fF
C19929 INPUT_3 AND2X1_LOC_819/a_8_24# 0.03fF
C19930 AND2X1_LOC_447/Y OR2X1_LOC_44/Y 0.71fF
C19931 AND2X1_LOC_857/Y OR2X1_LOC_48/B 0.08fF
C19932 VDD OR2X1_LOC_43/A 1.08fF
C19933 AND2X1_LOC_392/A AND2X1_LOC_566/a_8_24# 0.04fF
C19934 OR2X1_LOC_528/Y OR2X1_LOC_189/Y 0.03fF
C19935 OR2X1_LOC_306/Y OR2X1_LOC_91/A 0.03fF
C19936 OR2X1_LOC_604/A OR2X1_LOC_669/Y 1.05fF
C19937 AND2X1_LOC_732/a_8_24# OR2X1_LOC_599/A 0.01fF
C19938 AND2X1_LOC_81/B OR2X1_LOC_78/A 0.08fF
C19939 AND2X1_LOC_64/Y OR2X1_LOC_244/A 0.07fF
C19940 OR2X1_LOC_151/A AND2X1_LOC_111/a_8_24# 0.02fF
C19941 OR2X1_LOC_517/a_8_216# OR2X1_LOC_39/A 0.02fF
C19942 OR2X1_LOC_377/A OR2X1_LOC_837/Y 3.02fF
C19943 AND2X1_LOC_49/a_8_24# OR2X1_LOC_78/A 0.01fF
C19944 OR2X1_LOC_711/B OR2X1_LOC_479/Y 0.03fF
C19945 AND2X1_LOC_857/Y OR2X1_LOC_18/Y 0.07fF
C19946 OR2X1_LOC_380/Y OR2X1_LOC_44/Y 0.30fF
C19947 OR2X1_LOC_450/a_8_216# OR2X1_LOC_449/B 0.01fF
C19948 OR2X1_LOC_45/B OR2X1_LOC_268/a_8_216# 0.01fF
C19949 OR2X1_LOC_405/A AND2X1_LOC_40/Y 0.03fF
C19950 OR2X1_LOC_160/B OR2X1_LOC_208/a_36_216# 0.02fF
C19951 OR2X1_LOC_161/A OR2X1_LOC_736/A 0.03fF
C19952 OR2X1_LOC_793/A OR2X1_LOC_78/B 0.02fF
C19953 AND2X1_LOC_738/B OR2X1_LOC_26/Y 0.08fF
C19954 OR2X1_LOC_208/a_8_216# OR2X1_LOC_66/A 0.02fF
C19955 AND2X1_LOC_59/Y OR2X1_LOC_776/a_8_216# 0.01fF
C19956 OR2X1_LOC_26/Y OR2X1_LOC_56/A 0.07fF
C19957 OR2X1_LOC_837/Y AND2X1_LOC_824/B 0.00fF
C19958 INPUT_0 OR2X1_LOC_42/a_8_216# 0.01fF
C19959 OR2X1_LOC_855/a_8_216# AND2X1_LOC_48/A 0.01fF
C19960 AND2X1_LOC_12/Y AND2X1_LOC_421/a_8_24# 0.02fF
C19961 OR2X1_LOC_363/B OR2X1_LOC_287/B -0.00fF
C19962 OR2X1_LOC_616/Y AND2X1_LOC_866/B 0.03fF
C19963 AND2X1_LOC_714/B OR2X1_LOC_64/Y 0.03fF
C19964 AND2X1_LOC_803/B OR2X1_LOC_680/Y 0.27fF
C19965 OR2X1_LOC_528/Y OR2X1_LOC_527/Y 0.01fF
C19966 AND2X1_LOC_738/B OR2X1_LOC_89/A 0.17fF
C19967 OR2X1_LOC_643/A AND2X1_LOC_41/A 0.03fF
C19968 OR2X1_LOC_265/a_8_216# OR2X1_LOC_265/Y 0.01fF
C19969 OR2X1_LOC_121/B OR2X1_LOC_646/B 0.16fF
C19970 OR2X1_LOC_617/a_8_216# OR2X1_LOC_627/Y 0.01fF
C19971 OR2X1_LOC_89/A OR2X1_LOC_56/A 0.67fF
C19972 AND2X1_LOC_592/Y OR2X1_LOC_417/Y 0.03fF
C19973 AND2X1_LOC_702/Y OR2X1_LOC_298/a_8_216# 0.05fF
C19974 OR2X1_LOC_473/A OR2X1_LOC_140/B 0.00fF
C19975 AND2X1_LOC_41/A OR2X1_LOC_124/Y 0.03fF
C19976 AND2X1_LOC_41/A OR2X1_LOC_778/Y 0.10fF
C19977 AND2X1_LOC_59/Y OR2X1_LOC_653/Y 0.07fF
C19978 OR2X1_LOC_471/Y OR2X1_LOC_160/Y 0.02fF
C19979 AND2X1_LOC_787/A AND2X1_LOC_675/A 0.08fF
C19980 AND2X1_LOC_831/Y OR2X1_LOC_428/A 0.12fF
C19981 AND2X1_LOC_548/a_36_24# AND2X1_LOC_658/A 0.01fF
C19982 OR2X1_LOC_130/A OR2X1_LOC_737/A 0.07fF
C19983 OR2X1_LOC_609/a_36_216# OR2X1_LOC_59/Y 0.03fF
C19984 OR2X1_LOC_158/A AND2X1_LOC_128/a_8_24# 0.01fF
C19985 OR2X1_LOC_166/a_36_216# AND2X1_LOC_390/B 0.01fF
C19986 AND2X1_LOC_160/a_8_24# OR2X1_LOC_52/B 0.04fF
C19987 AND2X1_LOC_59/Y OR2X1_LOC_833/B 0.02fF
C19988 VDD OR2X1_LOC_60/a_8_216# 0.00fF
C19989 OR2X1_LOC_826/a_36_216# OR2X1_LOC_600/A 0.00fF
C19990 OR2X1_LOC_185/A OR2X1_LOC_738/A 0.06fF
C19991 D_INPUT_5 OR2X1_LOC_753/A 0.01fF
C19992 OR2X1_LOC_756/B OR2X1_LOC_287/B 0.09fF
C19993 OR2X1_LOC_689/A OR2X1_LOC_43/A 0.39fF
C19994 OR2X1_LOC_95/Y AND2X1_LOC_464/A 0.02fF
C19995 OR2X1_LOC_528/Y AND2X1_LOC_574/A 0.09fF
C19996 OR2X1_LOC_479/Y OR2X1_LOC_324/B 0.03fF
C19997 AND2X1_LOC_95/Y OR2X1_LOC_130/A 0.15fF
C19998 OR2X1_LOC_49/A OR2X1_LOC_55/a_8_216# 0.03fF
C19999 AND2X1_LOC_831/a_8_24# AND2X1_LOC_649/B 0.01fF
C20000 OR2X1_LOC_97/A AND2X1_LOC_109/a_8_24# 0.01fF
C20001 D_INPUT_7 AND2X1_LOC_51/a_36_24# 0.00fF
C20002 OR2X1_LOC_101/a_8_216# OR2X1_LOC_99/Y 0.03fF
C20003 VDD AND2X1_LOC_664/a_8_24# 0.00fF
C20004 OR2X1_LOC_686/B AND2X1_LOC_425/Y 0.00fF
C20005 OR2X1_LOC_109/Y OR2X1_LOC_44/Y 0.08fF
C20006 AND2X1_LOC_170/Y OR2X1_LOC_619/Y 0.04fF
C20007 AND2X1_LOC_56/B OR2X1_LOC_161/A 0.07fF
C20008 OR2X1_LOC_43/A OR2X1_LOC_829/a_8_216# 0.06fF
C20009 OR2X1_LOC_58/Y INPUT_1 0.04fF
C20010 AND2X1_LOC_86/a_8_24# OR2X1_LOC_244/A 0.01fF
C20011 OR2X1_LOC_502/A AND2X1_LOC_42/B 0.05fF
C20012 OR2X1_LOC_32/B OR2X1_LOC_36/Y 0.01fF
C20013 OR2X1_LOC_506/A OR2X1_LOC_449/B 0.29fF
C20014 OR2X1_LOC_3/Y AND2X1_LOC_348/A 0.00fF
C20015 AND2X1_LOC_45/a_8_24# OR2X1_LOC_78/B 0.05fF
C20016 OR2X1_LOC_196/B OR2X1_LOC_78/A 0.00fF
C20017 OR2X1_LOC_793/A OR2X1_LOC_375/A 0.01fF
C20018 OR2X1_LOC_427/A OR2X1_LOC_7/A 0.36fF
C20019 OR2X1_LOC_430/a_8_216# OR2X1_LOC_426/A 0.01fF
C20020 AND2X1_LOC_22/Y OR2X1_LOC_804/A 0.07fF
C20021 OR2X1_LOC_15/a_36_216# D_INPUT_1 0.00fF
C20022 AND2X1_LOC_218/a_8_24# AND2X1_LOC_656/Y 0.01fF
C20023 AND2X1_LOC_70/Y OR2X1_LOC_720/B -0.00fF
C20024 OR2X1_LOC_105/a_8_216# AND2X1_LOC_51/Y 0.06fF
C20025 AND2X1_LOC_512/Y OR2X1_LOC_417/Y 0.07fF
C20026 AND2X1_LOC_695/a_8_24# OR2X1_LOC_449/B 0.04fF
C20027 OR2X1_LOC_502/A OR2X1_LOC_705/Y 0.02fF
C20028 AND2X1_LOC_87/a_8_24# OR2X1_LOC_26/Y 0.01fF
C20029 OR2X1_LOC_283/Y AND2X1_LOC_286/Y 0.10fF
C20030 AND2X1_LOC_512/Y OR2X1_LOC_311/Y 0.26fF
C20031 AND2X1_LOC_19/Y D_INPUT_0 0.00fF
C20032 OR2X1_LOC_447/Y AND2X1_LOC_92/Y 0.42fF
C20033 OR2X1_LOC_865/a_36_216# OR2X1_LOC_859/B 0.00fF
C20034 AND2X1_LOC_42/B OR2X1_LOC_571/B 0.01fF
C20035 OR2X1_LOC_453/a_8_216# OR2X1_LOC_453/A 0.39fF
C20036 AND2X1_LOC_784/A OR2X1_LOC_91/a_36_216# 0.01fF
C20037 INPUT_0 OR2X1_LOC_532/B 2.01fF
C20038 OR2X1_LOC_634/A INPUT_1 0.53fF
C20039 OR2X1_LOC_589/A OR2X1_LOC_67/Y 0.00fF
C20040 OR2X1_LOC_405/A OR2X1_LOC_475/Y 0.01fF
C20041 OR2X1_LOC_161/B OR2X1_LOC_140/a_8_216# 0.01fF
C20042 OR2X1_LOC_221/A OR2X1_LOC_221/a_8_216# 0.18fF
C20043 OR2X1_LOC_68/B AND2X1_LOC_226/a_36_24# 0.00fF
C20044 OR2X1_LOC_445/a_36_216# OR2X1_LOC_553/A 0.00fF
C20045 OR2X1_LOC_47/Y AND2X1_LOC_614/a_36_24# 0.00fF
C20046 AND2X1_LOC_21/Y AND2X1_LOC_25/Y 0.96fF
C20047 AND2X1_LOC_40/Y OR2X1_LOC_285/Y 0.01fF
C20048 OR2X1_LOC_648/B AND2X1_LOC_289/a_8_24# 0.14fF
C20049 OR2X1_LOC_400/A AND2X1_LOC_42/B 0.01fF
C20050 AND2X1_LOC_861/B OR2X1_LOC_417/A 0.10fF
C20051 INPUT_4 OR2X1_LOC_430/a_8_216# 0.01fF
C20052 OR2X1_LOC_391/B OR2X1_LOC_864/a_8_216# 0.01fF
C20053 OR2X1_LOC_47/Y AND2X1_LOC_657/Y 0.03fF
C20054 OR2X1_LOC_276/B AND2X1_LOC_628/a_8_24# 0.02fF
C20055 OR2X1_LOC_70/Y AND2X1_LOC_317/a_8_24# 0.02fF
C20056 AND2X1_LOC_830/a_8_24# OR2X1_LOC_39/A 0.01fF
C20057 OR2X1_LOC_62/B AND2X1_LOC_414/a_8_24# 0.01fF
C20058 OR2X1_LOC_121/B OR2X1_LOC_506/A 0.47fF
C20059 OR2X1_LOC_446/a_8_216# OR2X1_LOC_87/A 0.02fF
C20060 AND2X1_LOC_363/A OR2X1_LOC_7/A 0.00fF
C20061 AND2X1_LOC_191/B OR2X1_LOC_47/Y 0.03fF
C20062 OR2X1_LOC_19/B OR2X1_LOC_71/a_8_216# 0.02fF
C20063 OR2X1_LOC_756/B OR2X1_LOC_436/Y 0.01fF
C20064 OR2X1_LOC_22/Y AND2X1_LOC_520/Y 0.01fF
C20065 AND2X1_LOC_744/a_36_24# OR2X1_LOC_780/B 0.00fF
C20066 OR2X1_LOC_47/Y AND2X1_LOC_469/B 0.14fF
C20067 OR2X1_LOC_154/A OR2X1_LOC_202/a_8_216# 0.02fF
C20068 GATE_366 OR2X1_LOC_481/A 0.03fF
C20069 AND2X1_LOC_686/a_8_24# AND2X1_LOC_452/Y 0.01fF
C20070 AND2X1_LOC_784/Y AND2X1_LOC_804/a_36_24# 0.00fF
C20071 OR2X1_LOC_461/Y AND2X1_LOC_56/B 0.01fF
C20072 OR2X1_LOC_74/A AND2X1_LOC_264/a_36_24# 0.00fF
C20073 OR2X1_LOC_278/A OR2X1_LOC_39/A 0.32fF
C20074 AND2X1_LOC_95/Y OR2X1_LOC_62/B 0.21fF
C20075 OR2X1_LOC_291/A OR2X1_LOC_26/Y 0.01fF
C20076 OR2X1_LOC_137/Y AND2X1_LOC_42/B 0.04fF
C20077 OR2X1_LOC_616/Y AND2X1_LOC_664/a_8_24# 0.03fF
C20078 AND2X1_LOC_729/B OR2X1_LOC_44/Y 0.03fF
C20079 OR2X1_LOC_377/A OR2X1_LOC_606/Y 0.15fF
C20080 OR2X1_LOC_128/B AND2X1_LOC_127/a_8_24# 0.00fF
C20081 AND2X1_LOC_56/B AND2X1_LOC_51/Y 1.94fF
C20082 AND2X1_LOC_45/a_8_24# OR2X1_LOC_375/A 0.01fF
C20083 OR2X1_LOC_115/a_8_216# D_INPUT_0 0.02fF
C20084 OR2X1_LOC_856/B AND2X1_LOC_47/Y 0.07fF
C20085 AND2X1_LOC_832/a_8_24# OR2X1_LOC_31/Y 0.01fF
C20086 OR2X1_LOC_426/A OR2X1_LOC_428/Y 0.58fF
C20087 AND2X1_LOC_728/a_8_24# AND2X1_LOC_147/Y 0.00fF
C20088 OR2X1_LOC_76/A OR2X1_LOC_76/Y 0.01fF
C20089 OR2X1_LOC_66/Y OR2X1_LOC_78/A 0.03fF
C20090 OR2X1_LOC_835/a_8_216# OR2X1_LOC_19/B 0.01fF
C20091 OR2X1_LOC_70/Y OR2X1_LOC_438/a_8_216# 0.01fF
C20092 AND2X1_LOC_502/a_8_24# OR2X1_LOC_71/Y 0.01fF
C20093 OR2X1_LOC_46/A OR2X1_LOC_6/A 0.16fF
C20094 OR2X1_LOC_864/A OR2X1_LOC_476/B 0.07fF
C20095 OR2X1_LOC_495/Y OR2X1_LOC_674/Y 0.24fF
C20096 AND2X1_LOC_465/A OR2X1_LOC_183/a_8_216# 0.03fF
C20097 OR2X1_LOC_391/A AND2X1_LOC_225/a_8_24# 0.03fF
C20098 OR2X1_LOC_557/A OR2X1_LOC_846/B 0.09fF
C20099 AND2X1_LOC_155/Y AND2X1_LOC_156/a_8_24# 0.03fF
C20100 AND2X1_LOC_303/A INPUT_1 0.00fF
C20101 OR2X1_LOC_64/Y AND2X1_LOC_645/A 0.02fF
C20102 AND2X1_LOC_21/Y AND2X1_LOC_51/Y 0.04fF
C20103 OR2X1_LOC_489/a_8_216# D_INPUT_1 0.01fF
C20104 AND2X1_LOC_550/A AND2X1_LOC_810/Y 0.03fF
C20105 OR2X1_LOC_836/a_8_216# OR2X1_LOC_19/B 0.02fF
C20106 AND2X1_LOC_578/A OR2X1_LOC_417/a_8_216# 0.47fF
C20107 AND2X1_LOC_64/Y OR2X1_LOC_354/a_8_216# 0.02fF
C20108 OR2X1_LOC_196/B OR2X1_LOC_155/A 0.02fF
C20109 AND2X1_LOC_866/B AND2X1_LOC_624/B 0.02fF
C20110 OR2X1_LOC_87/A AND2X1_LOC_7/Y 0.19fF
C20111 OR2X1_LOC_185/Y AND2X1_LOC_53/Y 0.01fF
C20112 AND2X1_LOC_734/Y OR2X1_LOC_406/A 0.39fF
C20113 AND2X1_LOC_40/Y OR2X1_LOC_545/a_8_216# 0.14fF
C20114 AND2X1_LOC_687/B OR2X1_LOC_7/A 0.08fF
C20115 OR2X1_LOC_421/A OR2X1_LOC_589/Y 0.01fF
C20116 INPUT_4 OR2X1_LOC_428/Y 0.01fF
C20117 OR2X1_LOC_549/B OR2X1_LOC_549/a_8_216# 0.07fF
C20118 OR2X1_LOC_476/a_8_216# OR2X1_LOC_476/Y -0.00fF
C20119 OR2X1_LOC_141/B OR2X1_LOC_814/A 0.03fF
C20120 OR2X1_LOC_427/A OR2X1_LOC_511/a_8_216# 0.02fF
C20121 AND2X1_LOC_776/Y AND2X1_LOC_785/a_8_24# 0.03fF
C20122 AND2X1_LOC_357/A OR2X1_LOC_437/A 0.00fF
C20123 OR2X1_LOC_362/A OR2X1_LOC_580/A 0.07fF
C20124 OR2X1_LOC_780/A OR2X1_LOC_449/B 0.00fF
C20125 AND2X1_LOC_509/Y AND2X1_LOC_657/A 0.02fF
C20126 AND2X1_LOC_48/A AND2X1_LOC_42/B 0.01fF
C20127 AND2X1_LOC_727/Y AND2X1_LOC_731/a_8_24# 0.00fF
C20128 OR2X1_LOC_604/a_8_216# AND2X1_LOC_454/A 0.47fF
C20129 OR2X1_LOC_185/Y OR2X1_LOC_223/A 0.03fF
C20130 AND2X1_LOC_784/A AND2X1_LOC_318/Y 0.02fF
C20131 OR2X1_LOC_756/B OR2X1_LOC_345/a_8_216# 0.02fF
C20132 AND2X1_LOC_727/Y AND2X1_LOC_564/A 0.03fF
C20133 OR2X1_LOC_524/Y OR2X1_LOC_152/a_36_216# 0.17fF
C20134 OR2X1_LOC_417/Y AND2X1_LOC_712/B 0.01fF
C20135 AND2X1_LOC_95/Y OR2X1_LOC_365/B 0.04fF
C20136 OR2X1_LOC_203/Y OR2X1_LOC_786/Y 0.00fF
C20137 OR2X1_LOC_420/Y OR2X1_LOC_95/Y 0.01fF
C20138 AND2X1_LOC_259/Y OR2X1_LOC_55/a_8_216# 0.01fF
C20139 OR2X1_LOC_375/A OR2X1_LOC_66/a_36_216# 0.00fF
C20140 AND2X1_LOC_308/a_8_24# AND2X1_LOC_727/A 0.01fF
C20141 OR2X1_LOC_22/Y AND2X1_LOC_856/B 0.01fF
C20142 OR2X1_LOC_99/Y AND2X1_LOC_88/Y 0.23fF
C20143 OR2X1_LOC_392/B AND2X1_LOC_7/B 0.10fF
C20144 AND2X1_LOC_91/B OR2X1_LOC_576/A 0.01fF
C20145 OR2X1_LOC_484/a_8_216# OR2X1_LOC_13/B 0.08fF
C20146 OR2X1_LOC_64/Y AND2X1_LOC_477/A 0.06fF
C20147 OR2X1_LOC_805/A OR2X1_LOC_374/Y 0.10fF
C20148 OR2X1_LOC_404/Y OR2X1_LOC_720/B 0.00fF
C20149 OR2X1_LOC_70/Y AND2X1_LOC_169/a_8_24# 0.01fF
C20150 AND2X1_LOC_727/Y AND2X1_LOC_727/B 0.01fF
C20151 AND2X1_LOC_64/Y OR2X1_LOC_691/B 0.03fF
C20152 OR2X1_LOC_32/B AND2X1_LOC_202/a_36_24# 0.01fF
C20153 AND2X1_LOC_42/B AND2X1_LOC_106/a_8_24# 0.01fF
C20154 OR2X1_LOC_623/a_8_216# AND2X1_LOC_31/Y 0.05fF
C20155 OR2X1_LOC_43/A OR2X1_LOC_67/Y 0.46fF
C20156 OR2X1_LOC_199/a_8_216# AND2X1_LOC_22/Y 0.00fF
C20157 AND2X1_LOC_802/B AND2X1_LOC_802/Y 0.11fF
C20158 AND2X1_LOC_56/B OR2X1_LOC_551/B 0.07fF
C20159 AND2X1_LOC_303/a_36_24# OR2X1_LOC_437/A 0.01fF
C20160 OR2X1_LOC_468/A OR2X1_LOC_180/B 0.83fF
C20161 OR2X1_LOC_111/a_36_216# OR2X1_LOC_158/A 0.02fF
C20162 OR2X1_LOC_136/Y OR2X1_LOC_12/Y 0.14fF
C20163 OR2X1_LOC_174/a_8_216# OR2X1_LOC_390/A 0.03fF
C20164 OR2X1_LOC_121/B OR2X1_LOC_780/A 0.14fF
C20165 AND2X1_LOC_633/Y AND2X1_LOC_640/a_8_24# 0.11fF
C20166 OR2X1_LOC_606/a_8_216# OR2X1_LOC_532/B 0.07fF
C20167 OR2X1_LOC_326/a_36_216# OR2X1_LOC_532/Y 0.00fF
C20168 OR2X1_LOC_144/a_8_216# OR2X1_LOC_526/Y 0.41fF
C20169 OR2X1_LOC_240/a_8_216# OR2X1_LOC_80/A 0.04fF
C20170 OR2X1_LOC_243/A OR2X1_LOC_68/B 0.00fF
C20171 OR2X1_LOC_70/A OR2X1_LOC_25/a_36_216# 0.00fF
C20172 OR2X1_LOC_151/A OR2X1_LOC_267/Y 0.04fF
C20173 OR2X1_LOC_36/Y AND2X1_LOC_222/Y 0.04fF
C20174 OR2X1_LOC_523/B AND2X1_LOC_22/Y 0.01fF
C20175 OR2X1_LOC_564/B OR2X1_LOC_192/B 0.02fF
C20176 OR2X1_LOC_91/a_8_216# AND2X1_LOC_222/Y 0.01fF
C20177 AND2X1_LOC_729/Y OR2X1_LOC_526/a_36_216# 0.00fF
C20178 AND2X1_LOC_477/A OR2X1_LOC_417/A 0.00fF
C20179 OR2X1_LOC_405/A AND2X1_LOC_406/a_36_24# 0.06fF
C20180 AND2X1_LOC_693/a_8_24# AND2X1_LOC_36/Y 0.14fF
C20181 D_INPUT_0 OR2X1_LOC_4/a_8_216# 0.01fF
C20182 OR2X1_LOC_121/B OR2X1_LOC_227/Y 0.02fF
C20183 D_INPUT_3 OR2X1_LOC_54/Y 0.16fF
C20184 OR2X1_LOC_154/A OR2X1_LOC_724/A 0.47fF
C20185 OR2X1_LOC_48/B OR2X1_LOC_437/A 0.04fF
C20186 OR2X1_LOC_419/Y OR2X1_LOC_371/Y 0.10fF
C20187 AND2X1_LOC_12/a_8_24# INPUT_6 0.01fF
C20188 AND2X1_LOC_483/Y AND2X1_LOC_483/a_8_24# 0.02fF
C20189 OR2X1_LOC_18/Y OR2X1_LOC_437/A 0.08fF
C20190 OR2X1_LOC_121/B D_INPUT_1 0.01fF
C20191 AND2X1_LOC_721/Y OR2X1_LOC_108/Y 0.02fF
C20192 OR2X1_LOC_362/A AND2X1_LOC_44/Y 0.51fF
C20193 OR2X1_LOC_333/B OR2X1_LOC_358/A 0.10fF
C20194 OR2X1_LOC_40/Y OR2X1_LOC_18/a_36_216# 0.00fF
C20195 OR2X1_LOC_6/B OR2X1_LOC_428/A 0.08fF
C20196 AND2X1_LOC_713/Y OR2X1_LOC_428/A 0.00fF
C20197 OR2X1_LOC_114/B AND2X1_LOC_248/a_8_24# 0.01fF
C20198 OR2X1_LOC_269/B OR2X1_LOC_80/A 0.09fF
C20199 AND2X1_LOC_448/a_36_24# OR2X1_LOC_428/A 0.00fF
C20200 OR2X1_LOC_289/a_8_216# OR2X1_LOC_46/A 0.01fF
C20201 OR2X1_LOC_49/A OR2X1_LOC_96/Y 0.01fF
C20202 OR2X1_LOC_36/Y OR2X1_LOC_423/Y 0.53fF
C20203 AND2X1_LOC_270/a_8_24# OR2X1_LOC_368/A 0.01fF
C20204 INPUT_5 OR2X1_LOC_696/A 0.20fF
C20205 OR2X1_LOC_45/B AND2X1_LOC_447/Y 0.01fF
C20206 OR2X1_LOC_45/B AND2X1_LOC_219/a_8_24# 0.01fF
C20207 OR2X1_LOC_45/B AND2X1_LOC_334/Y 0.01fF
C20208 OR2X1_LOC_41/Y OR2X1_LOC_43/a_36_216# 0.00fF
C20209 AND2X1_LOC_227/Y AND2X1_LOC_139/A 0.01fF
C20210 OR2X1_LOC_599/A AND2X1_LOC_592/a_8_24# 0.01fF
C20211 OR2X1_LOC_696/A AND2X1_LOC_839/a_8_24# 0.01fF
C20212 OR2X1_LOC_87/A OR2X1_LOC_140/Y 0.03fF
C20213 AND2X1_LOC_91/B AND2X1_LOC_41/A 0.06fF
C20214 AND2X1_LOC_450/Y AND2X1_LOC_451/Y 0.10fF
C20215 OR2X1_LOC_185/A AND2X1_LOC_36/Y 0.67fF
C20216 OR2X1_LOC_156/B OR2X1_LOC_803/A 0.01fF
C20217 OR2X1_LOC_147/A AND2X1_LOC_7/B 0.03fF
C20218 OR2X1_LOC_51/Y OR2X1_LOC_12/Y 1.44fF
C20219 OR2X1_LOC_176/Y OR2X1_LOC_91/A 0.04fF
C20220 AND2X1_LOC_540/a_8_24# AND2X1_LOC_465/A 0.01fF
C20221 OR2X1_LOC_482/Y OR2X1_LOC_108/Y 0.11fF
C20222 OR2X1_LOC_51/Y OR2X1_LOC_766/Y 0.01fF
C20223 OR2X1_LOC_856/B OR2X1_LOC_186/a_8_216# 0.03fF
C20224 OR2X1_LOC_9/Y OR2X1_LOC_600/A 0.08fF
C20225 AND2X1_LOC_430/a_8_24# AND2X1_LOC_430/B 0.10fF
C20226 OR2X1_LOC_462/a_8_216# OR2X1_LOC_68/B 0.01fF
C20227 OR2X1_LOC_787/Y OR2X1_LOC_303/B 0.08fF
C20228 GATE_366 AND2X1_LOC_789/Y 0.07fF
C20229 OR2X1_LOC_693/Y OR2X1_LOC_744/A 0.01fF
C20230 AND2X1_LOC_151/a_8_24# OR2X1_LOC_142/Y 0.01fF
C20231 OR2X1_LOC_91/A AND2X1_LOC_212/Y 0.15fF
C20232 AND2X1_LOC_357/A AND2X1_LOC_715/A 0.03fF
C20233 OR2X1_LOC_474/Y AND2X1_LOC_44/Y 0.05fF
C20234 OR2X1_LOC_516/Y AND2X1_LOC_580/A 0.07fF
C20235 AND2X1_LOC_788/a_36_24# OR2X1_LOC_59/Y 0.00fF
C20236 AND2X1_LOC_724/Y OR2X1_LOC_604/A 0.01fF
C20237 OR2X1_LOC_97/A OR2X1_LOC_775/a_36_216# 0.03fF
C20238 AND2X1_LOC_601/a_8_24# OR2X1_LOC_390/B 0.04fF
C20239 OR2X1_LOC_833/Y OR2X1_LOC_458/B 0.02fF
C20240 AND2X1_LOC_810/a_36_24# OR2X1_LOC_47/Y 0.01fF
C20241 AND2X1_LOC_656/a_36_24# AND2X1_LOC_772/Y 0.01fF
C20242 OR2X1_LOC_101/a_8_216# AND2X1_LOC_22/Y 0.03fF
C20243 AND2X1_LOC_3/Y OR2X1_LOC_174/Y 0.01fF
C20244 OR2X1_LOC_104/a_8_216# INPUT_2 0.14fF
C20245 AND2X1_LOC_766/a_8_24# OR2X1_LOC_402/Y 0.03fF
C20246 AND2X1_LOC_352/a_8_24# OR2X1_LOC_91/A 0.06fF
C20247 VDD OR2X1_LOC_585/Y -0.00fF
C20248 OR2X1_LOC_45/B AND2X1_LOC_649/B 0.09fF
C20249 OR2X1_LOC_427/A OR2X1_LOC_753/a_8_216# 0.01fF
C20250 AND2X1_LOC_353/a_36_24# OR2X1_LOC_91/A 0.01fF
C20251 AND2X1_LOC_122/a_8_24# OR2X1_LOC_217/A 0.08fF
C20252 OR2X1_LOC_426/B OR2X1_LOC_666/A 0.18fF
C20253 OR2X1_LOC_696/A AND2X1_LOC_839/B 0.02fF
C20254 OR2X1_LOC_805/A OR2X1_LOC_392/B 0.10fF
C20255 AND2X1_LOC_228/Y OR2X1_LOC_230/Y 0.01fF
C20256 AND2X1_LOC_509/Y VDD 0.27fF
C20257 OR2X1_LOC_235/B AND2X1_LOC_18/Y 0.05fF
C20258 VDD OR2X1_LOC_570/A -0.00fF
C20259 OR2X1_LOC_828/B OR2X1_LOC_855/A 0.01fF
C20260 AND2X1_LOC_70/Y AND2X1_LOC_628/a_8_24# 0.01fF
C20261 AND2X1_LOC_566/B OR2X1_LOC_92/Y 0.03fF
C20262 OR2X1_LOC_45/B AND2X1_LOC_448/Y 0.01fF
C20263 OR2X1_LOC_756/B OR2X1_LOC_160/B 0.24fF
C20264 AND2X1_LOC_675/Y AND2X1_LOC_500/Y 0.02fF
C20265 AND2X1_LOC_22/Y OR2X1_LOC_130/A 0.42fF
C20266 AND2X1_LOC_436/B OR2X1_LOC_428/A 0.72fF
C20267 OR2X1_LOC_278/A AND2X1_LOC_608/a_36_24# 0.00fF
C20268 AND2X1_LOC_91/B OR2X1_LOC_631/B 0.03fF
C20269 AND2X1_LOC_330/a_8_24# AND2X1_LOC_512/Y 0.03fF
C20270 AND2X1_LOC_341/a_36_24# AND2X1_LOC_228/Y 0.01fF
C20271 AND2X1_LOC_181/a_8_24# OR2X1_LOC_329/B 0.03fF
C20272 OR2X1_LOC_217/Y AND2X1_LOC_44/Y 0.00fF
C20273 OR2X1_LOC_229/a_8_216# AND2X1_LOC_228/Y 0.48fF
C20274 OR2X1_LOC_223/A OR2X1_LOC_578/B 0.03fF
C20275 AND2X1_LOC_22/Y AND2X1_LOC_7/a_8_24# 0.02fF
C20276 OR2X1_LOC_710/B OR2X1_LOC_502/A 0.07fF
C20277 OR2X1_LOC_121/a_8_216# AND2X1_LOC_56/B 0.01fF
C20278 OR2X1_LOC_71/Y OR2X1_LOC_13/B 0.03fF
C20279 AND2X1_LOC_575/a_8_24# AND2X1_LOC_474/Y 0.03fF
C20280 OR2X1_LOC_9/Y OR2X1_LOC_619/Y 0.01fF
C20281 OR2X1_LOC_136/a_36_216# AND2X1_LOC_211/B 0.00fF
C20282 OR2X1_LOC_857/B OR2X1_LOC_375/A 0.14fF
C20283 AND2X1_LOC_787/a_8_24# OR2X1_LOC_600/A 0.01fF
C20284 AND2X1_LOC_716/Y OR2X1_LOC_426/B 0.83fF
C20285 OR2X1_LOC_419/Y AND2X1_LOC_222/Y 0.03fF
C20286 OR2X1_LOC_234/Y AND2X1_LOC_240/a_8_24# 0.00fF
C20287 OR2X1_LOC_95/Y OR2X1_LOC_385/a_36_216# 0.00fF
C20288 OR2X1_LOC_158/A INPUT_4 0.04fF
C20289 OR2X1_LOC_744/A AND2X1_LOC_651/a_8_24# 0.01fF
C20290 OR2X1_LOC_426/B AND2X1_LOC_654/Y 0.09fF
C20291 OR2X1_LOC_389/B OR2X1_LOC_389/a_8_216# 0.01fF
C20292 OR2X1_LOC_47/Y OR2X1_LOC_164/a_8_216# 0.01fF
C20293 OR2X1_LOC_377/A OR2X1_LOC_622/A 0.03fF
C20294 AND2X1_LOC_50/Y OR2X1_LOC_637/Y 0.02fF
C20295 AND2X1_LOC_95/Y OR2X1_LOC_468/A 0.05fF
C20296 AND2X1_LOC_715/A OR2X1_LOC_18/Y 0.37fF
C20297 AND2X1_LOC_572/Y OR2X1_LOC_600/A 0.05fF
C20298 OR2X1_LOC_529/Y OR2X1_LOC_428/A 0.02fF
C20299 OR2X1_LOC_812/B OR2X1_LOC_862/B 0.12fF
C20300 AND2X1_LOC_61/Y OR2X1_LOC_619/Y 0.07fF
C20301 VDD AND2X1_LOC_132/a_8_24# 0.00fF
C20302 OR2X1_LOC_855/a_8_216# AND2X1_LOC_3/Y 0.01fF
C20303 OR2X1_LOC_359/a_8_216# AND2X1_LOC_12/Y 0.01fF
C20304 AND2X1_LOC_191/B OR2X1_LOC_625/Y 0.07fF
C20305 AND2X1_LOC_12/Y OR2X1_LOC_35/a_8_216# 0.01fF
C20306 OR2X1_LOC_95/Y AND2X1_LOC_750/a_8_24# 0.00fF
C20307 OR2X1_LOC_135/Y AND2X1_LOC_211/B 0.10fF
C20308 OR2X1_LOC_308/a_8_216# AND2X1_LOC_41/A 0.02fF
C20309 AND2X1_LOC_741/Y AND2X1_LOC_221/a_36_24# 0.01fF
C20310 OR2X1_LOC_663/A OR2X1_LOC_502/A 0.03fF
C20311 OR2X1_LOC_512/A OR2X1_LOC_307/B 0.00fF
C20312 AND2X1_LOC_593/a_8_24# OR2X1_LOC_44/Y 0.02fF
C20313 AND2X1_LOC_141/a_8_24# AND2X1_LOC_573/A 0.03fF
C20314 OR2X1_LOC_694/a_8_216# OR2X1_LOC_51/Y 0.01fF
C20315 OR2X1_LOC_709/A OR2X1_LOC_793/B 0.01fF
C20316 OR2X1_LOC_6/A INPUT_2 0.18fF
C20317 OR2X1_LOC_605/A AND2X1_LOC_604/a_36_24# 0.01fF
C20318 OR2X1_LOC_161/A AND2X1_LOC_92/Y 9.54fF
C20319 OR2X1_LOC_600/A OR2X1_LOC_96/B 0.00fF
C20320 OR2X1_LOC_528/Y AND2X1_LOC_806/A 0.02fF
C20321 OR2X1_LOC_139/A OR2X1_LOC_473/Y 0.05fF
C20322 AND2X1_LOC_443/a_36_24# OR2X1_LOC_52/B 0.00fF
C20323 OR2X1_LOC_45/B AND2X1_LOC_729/B 0.03fF
C20324 OR2X1_LOC_534/a_8_216# OR2X1_LOC_331/Y 0.01fF
C20325 AND2X1_LOC_503/a_8_24# OR2X1_LOC_502/A 0.09fF
C20326 AND2X1_LOC_40/Y D_INPUT_4 0.07fF
C20327 AND2X1_LOC_573/a_8_24# AND2X1_LOC_735/Y 0.00fF
C20328 OR2X1_LOC_394/Y OR2X1_LOC_394/a_8_216# 0.01fF
C20329 OR2X1_LOC_87/A OR2X1_LOC_797/a_8_216# 0.01fF
C20330 OR2X1_LOC_316/Y OR2X1_LOC_59/Y 0.04fF
C20331 AND2X1_LOC_655/A AND2X1_LOC_434/Y 0.10fF
C20332 AND2X1_LOC_367/A OR2X1_LOC_250/Y 0.10fF
C20333 AND2X1_LOC_329/a_36_24# OR2X1_LOC_596/A 0.01fF
C20334 OR2X1_LOC_633/B AND2X1_LOC_262/a_8_24# 0.01fF
C20335 OR2X1_LOC_160/B OR2X1_LOC_76/Y 0.00fF
C20336 AND2X1_LOC_118/a_8_24# OR2X1_LOC_786/A 0.08fF
C20337 OR2X1_LOC_600/A AND2X1_LOC_852/Y 0.03fF
C20338 AND2X1_LOC_486/Y OR2X1_LOC_495/Y 0.03fF
C20339 AND2X1_LOC_703/Y OR2X1_LOC_64/Y 0.01fF
C20340 AND2X1_LOC_729/a_36_24# OR2X1_LOC_485/A 0.00fF
C20341 AND2X1_LOC_19/Y OR2X1_LOC_87/Y 0.00fF
C20342 OR2X1_LOC_577/a_36_216# D_GATE_366 0.00fF
C20343 OR2X1_LOC_822/Y OR2X1_LOC_753/A 0.04fF
C20344 AND2X1_LOC_363/Y AND2X1_LOC_359/a_8_24# 0.01fF
C20345 AND2X1_LOC_560/a_8_24# OR2X1_LOC_95/Y 0.01fF
C20346 OR2X1_LOC_26/Y AND2X1_LOC_285/Y 0.00fF
C20347 OR2X1_LOC_687/Y OR2X1_LOC_78/B 0.19fF
C20348 OR2X1_LOC_319/B OR2X1_LOC_319/a_36_216# 0.02fF
C20349 OR2X1_LOC_154/A OR2X1_LOC_632/Y 0.12fF
C20350 OR2X1_LOC_160/B AND2X1_LOC_159/a_36_24# 0.01fF
C20351 AND2X1_LOC_297/a_8_24# OR2X1_LOC_736/A 0.01fF
C20352 OR2X1_LOC_3/Y OR2X1_LOC_583/a_8_216# 0.02fF
C20353 VDD OR2X1_LOC_564/B 0.08fF
C20354 AND2X1_LOC_22/Y OR2X1_LOC_62/B 0.05fF
C20355 OR2X1_LOC_840/A OR2X1_LOC_739/A 0.05fF
C20356 OR2X1_LOC_70/Y OR2X1_LOC_765/a_8_216# 0.01fF
C20357 AND2X1_LOC_367/B OR2X1_LOC_753/A 0.04fF
C20358 OR2X1_LOC_40/Y AND2X1_LOC_640/Y 0.00fF
C20359 OR2X1_LOC_756/B OR2X1_LOC_553/A 0.03fF
C20360 OR2X1_LOC_788/B OR2X1_LOC_365/B 0.16fF
C20361 OR2X1_LOC_604/A OR2X1_LOC_371/Y 0.10fF
C20362 OR2X1_LOC_648/A OR2X1_LOC_778/Y 0.40fF
C20363 VDD AND2X1_LOC_240/Y 0.07fF
C20364 OR2X1_LOC_85/A OR2X1_LOC_234/Y 0.01fF
C20365 OR2X1_LOC_160/A OR2X1_LOC_330/Y 0.02fF
C20366 AND2X1_LOC_228/Y AND2X1_LOC_857/Y 0.03fF
C20367 OR2X1_LOC_49/A AND2X1_LOC_825/a_8_24# 0.03fF
C20368 OR2X1_LOC_51/Y OR2X1_LOC_239/a_8_216# 0.11fF
C20369 OR2X1_LOC_89/A AND2X1_LOC_285/Y 0.03fF
C20370 OR2X1_LOC_532/B AND2X1_LOC_7/B 0.25fF
C20371 OR2X1_LOC_757/A AND2X1_LOC_620/a_8_24# 0.12fF
C20372 AND2X1_LOC_367/A OR2X1_LOC_36/Y 0.01fF
C20373 AND2X1_LOC_70/Y AND2X1_LOC_683/a_8_24# 0.01fF
C20374 VDD OR2X1_LOC_299/Y 0.04fF
C20375 AND2X1_LOC_227/Y OR2X1_LOC_184/a_8_216# 0.01fF
C20376 AND2X1_LOC_38/a_8_24# OR2X1_LOC_66/A 0.04fF
C20377 AND2X1_LOC_753/B AND2X1_LOC_43/B 0.91fF
C20378 AND2X1_LOC_576/Y AND2X1_LOC_850/A 0.01fF
C20379 OR2X1_LOC_706/B OR2X1_LOC_706/a_8_216# 0.47fF
C20380 OR2X1_LOC_158/A AND2X1_LOC_849/A 0.08fF
C20381 OR2X1_LOC_574/A OR2X1_LOC_78/A 0.29fF
C20382 OR2X1_LOC_676/Y AND2X1_LOC_13/a_8_24# 0.02fF
C20383 OR2X1_LOC_186/Y OR2X1_LOC_814/A 0.03fF
C20384 OR2X1_LOC_472/A OR2X1_LOC_410/a_8_216# 0.06fF
C20385 AND2X1_LOC_859/B AND2X1_LOC_287/B 0.12fF
C20386 INPUT_1 OR2X1_LOC_633/A 0.09fF
C20387 OR2X1_LOC_479/Y OR2X1_LOC_841/A 0.04fF
C20388 AND2X1_LOC_40/Y OR2X1_LOC_653/A 0.01fF
C20389 OR2X1_LOC_364/A OR2X1_LOC_502/A 0.09fF
C20390 AND2X1_LOC_95/Y AND2X1_LOC_487/a_8_24# 0.11fF
C20391 VDD AND2X1_LOC_67/Y 0.27fF
C20392 OR2X1_LOC_185/Y OR2X1_LOC_502/A 0.07fF
C20393 AND2X1_LOC_95/Y OR2X1_LOC_128/A 0.02fF
C20394 OR2X1_LOC_467/A OR2X1_LOC_466/a_36_216# 0.00fF
C20395 AND2X1_LOC_520/Y OR2X1_LOC_39/A 0.05fF
C20396 AND2X1_LOC_468/B AND2X1_LOC_593/Y 0.04fF
C20397 AND2X1_LOC_605/Y AND2X1_LOC_454/A 0.02fF
C20398 AND2X1_LOC_40/Y OR2X1_LOC_673/Y 0.07fF
C20399 OR2X1_LOC_756/B OR2X1_LOC_219/B 0.07fF
C20400 OR2X1_LOC_137/Y OR2X1_LOC_663/A 0.12fF
C20401 OR2X1_LOC_405/A AND2X1_LOC_43/B 0.12fF
C20402 OR2X1_LOC_840/A OR2X1_LOC_269/B 0.01fF
C20403 OR2X1_LOC_282/Y OR2X1_LOC_56/A 0.05fF
C20404 OR2X1_LOC_290/Y OR2X1_LOC_26/Y 0.01fF
C20405 OR2X1_LOC_640/A AND2X1_LOC_8/Y 0.02fF
C20406 OR2X1_LOC_791/B OR2X1_LOC_260/Y 0.24fF
C20407 AND2X1_LOC_859/a_8_24# OR2X1_LOC_278/Y 0.00fF
C20408 OR2X1_LOC_439/a_36_216# OR2X1_LOC_161/B 0.01fF
C20409 OR2X1_LOC_524/Y OR2X1_LOC_680/Y 0.03fF
C20410 OR2X1_LOC_427/A OR2X1_LOC_236/a_8_216# 0.01fF
C20411 AND2X1_LOC_196/Y OR2X1_LOC_13/Y 0.00fF
C20412 AND2X1_LOC_22/Y AND2X1_LOC_88/Y 0.03fF
C20413 AND2X1_LOC_332/a_36_24# OR2X1_LOC_417/A 0.00fF
C20414 OR2X1_LOC_459/B OR2X1_LOC_375/A 0.03fF
C20415 OR2X1_LOC_442/a_8_216# AND2X1_LOC_477/Y 0.05fF
C20416 INPUT_3 AND2X1_LOC_55/a_8_24# 0.03fF
C20417 AND2X1_LOC_51/Y AND2X1_LOC_92/Y 0.13fF
C20418 VDD OR2X1_LOC_451/A -0.00fF
C20419 AND2X1_LOC_186/a_8_24# OR2X1_LOC_39/A 0.01fF
C20420 OR2X1_LOC_816/a_8_216# OR2X1_LOC_253/a_8_216# 0.47fF
C20421 OR2X1_LOC_185/Y OR2X1_LOC_571/B 0.16fF
C20422 OR2X1_LOC_377/A OR2X1_LOC_835/B 0.31fF
C20423 AND2X1_LOC_185/a_8_24# OR2X1_LOC_74/A 0.08fF
C20424 OR2X1_LOC_431/Y OR2X1_LOC_59/Y 0.01fF
C20425 OR2X1_LOC_32/B OR2X1_LOC_80/Y 0.03fF
C20426 AND2X1_LOC_339/B OR2X1_LOC_75/Y 0.01fF
C20427 AND2X1_LOC_557/Y AND2X1_LOC_563/a_8_24# 0.20fF
C20428 OR2X1_LOC_631/B AND2X1_LOC_72/Y 0.03fF
C20429 OR2X1_LOC_401/B OR2X1_LOC_78/B 0.01fF
C20430 AND2X1_LOC_716/Y OR2X1_LOC_743/A 0.07fF
C20431 AND2X1_LOC_95/Y OR2X1_LOC_449/B 0.03fF
C20432 OR2X1_LOC_687/Y OR2X1_LOC_375/A 0.03fF
C20433 OR2X1_LOC_18/Y OR2X1_LOC_753/A 0.06fF
C20434 AND2X1_LOC_174/a_36_24# AND2X1_LOC_650/Y 0.00fF
C20435 OR2X1_LOC_823/Y AND2X1_LOC_836/a_8_24# 0.23fF
C20436 OR2X1_LOC_465/a_36_216# OR2X1_LOC_553/A 0.00fF
C20437 OR2X1_LOC_643/Y OR2X1_LOC_78/B 0.03fF
C20438 OR2X1_LOC_230/a_36_216# AND2X1_LOC_857/Y 0.00fF
C20439 AND2X1_LOC_310/a_8_24# OR2X1_LOC_814/A 0.01fF
C20440 OR2X1_LOC_743/A AND2X1_LOC_654/Y 0.07fF
C20441 AND2X1_LOC_719/Y AND2X1_LOC_851/B 0.10fF
C20442 OR2X1_LOC_161/B AND2X1_LOC_418/a_8_24# 0.01fF
C20443 AND2X1_LOC_459/Y AND2X1_LOC_463/a_8_24# 0.09fF
C20444 OR2X1_LOC_835/A OR2X1_LOC_835/a_8_216# 0.47fF
C20445 OR2X1_LOC_76/Y OR2X1_LOC_553/A 0.06fF
C20446 OR2X1_LOC_865/Y OR2X1_LOC_859/B 0.01fF
C20447 AND2X1_LOC_175/B AND2X1_LOC_211/B 0.36fF
C20448 OR2X1_LOC_204/Y OR2X1_LOC_203/Y 0.29fF
C20449 OR2X1_LOC_210/B OR2X1_LOC_210/a_8_216# 0.47fF
C20450 OR2X1_LOC_91/Y OR2X1_LOC_26/Y 0.16fF
C20451 AND2X1_LOC_340/a_36_24# AND2X1_LOC_227/Y 0.02fF
C20452 OR2X1_LOC_617/a_8_216# AND2X1_LOC_805/Y 0.01fF
C20453 AND2X1_LOC_719/a_8_24# AND2X1_LOC_621/Y 0.03fF
C20454 OR2X1_LOC_665/Y AND2X1_LOC_624/A 6.13fF
C20455 AND2X1_LOC_624/A AND2X1_LOC_474/Y 0.03fF
C20456 AND2X1_LOC_271/a_8_24# OR2X1_LOC_549/A 0.01fF
C20457 OR2X1_LOC_244/B OR2X1_LOC_62/B 0.00fF
C20458 AND2X1_LOC_391/Y OR2X1_LOC_255/a_8_216# 0.08fF
C20459 OR2X1_LOC_276/B AND2X1_LOC_18/Y 0.21fF
C20460 OR2X1_LOC_485/A AND2X1_LOC_624/A 0.03fF
C20461 AND2X1_LOC_576/Y OR2X1_LOC_498/Y 0.07fF
C20462 OR2X1_LOC_93/a_8_216# OR2X1_LOC_6/A 0.01fF
C20463 OR2X1_LOC_72/Y AND2X1_LOC_202/Y 0.04fF
C20464 OR2X1_LOC_91/Y OR2X1_LOC_89/A 2.32fF
C20465 OR2X1_LOC_235/B OR2X1_LOC_813/A 0.04fF
C20466 AND2X1_LOC_716/Y OR2X1_LOC_246/A 0.10fF
C20467 OR2X1_LOC_121/B OR2X1_LOC_737/A 0.08fF
C20468 OR2X1_LOC_131/Y AND2X1_LOC_572/A 0.13fF
C20469 OR2X1_LOC_70/Y OR2X1_LOC_316/Y 0.03fF
C20470 AND2X1_LOC_456/Y OR2X1_LOC_36/Y 0.03fF
C20471 OR2X1_LOC_617/Y OR2X1_LOC_39/A 0.00fF
C20472 AND2X1_LOC_191/B AND2X1_LOC_663/a_8_24# 0.01fF
C20473 AND2X1_LOC_810/Y AND2X1_LOC_663/A 0.03fF
C20474 AND2X1_LOC_156/a_36_24# OR2X1_LOC_619/Y 0.00fF
C20475 OR2X1_LOC_789/a_8_216# OR2X1_LOC_269/B 0.05fF
C20476 AND2X1_LOC_95/Y OR2X1_LOC_121/B 0.04fF
C20477 AND2X1_LOC_654/Y OR2X1_LOC_246/A 0.02fF
C20478 OR2X1_LOC_36/Y OR2X1_LOC_74/A 0.36fF
C20479 OR2X1_LOC_319/B OR2X1_LOC_532/B 0.13fF
C20480 AND2X1_LOC_364/A AND2X1_LOC_326/a_8_24# 0.06fF
C20481 OR2X1_LOC_91/a_8_216# OR2X1_LOC_74/A 0.16fF
C20482 OR2X1_LOC_409/B OR2X1_LOC_762/Y 0.20fF
C20483 AND2X1_LOC_52/a_8_24# AND2X1_LOC_53/Y 0.03fF
C20484 AND2X1_LOC_229/a_8_24# OR2X1_LOC_68/B 0.01fF
C20485 OR2X1_LOC_633/Y OR2X1_LOC_121/B 0.22fF
C20486 AND2X1_LOC_88/a_8_24# OR2X1_LOC_99/Y 0.07fF
C20487 OR2X1_LOC_417/Y AND2X1_LOC_453/Y 0.18fF
C20488 OR2X1_LOC_177/Y AND2X1_LOC_222/Y 0.02fF
C20489 AND2X1_LOC_717/B AND2X1_LOC_458/a_8_24# 0.03fF
C20490 OR2X1_LOC_71/Y AND2X1_LOC_266/a_8_24# 0.01fF
C20491 OR2X1_LOC_235/B AND2X1_LOC_672/a_8_24# 0.01fF
C20492 OR2X1_LOC_574/A OR2X1_LOC_155/A 0.21fF
C20493 OR2X1_LOC_279/a_36_216# OR2X1_LOC_44/Y 0.03fF
C20494 OR2X1_LOC_294/Y OR2X1_LOC_736/a_36_216# 0.00fF
C20495 OR2X1_LOC_682/a_8_216# OR2X1_LOC_3/Y 0.02fF
C20496 OR2X1_LOC_329/B AND2X1_LOC_798/A 0.03fF
C20497 OR2X1_LOC_279/a_8_216# AND2X1_LOC_806/A 0.49fF
C20498 OR2X1_LOC_630/a_8_216# OR2X1_LOC_62/B 0.01fF
C20499 AND2X1_LOC_53/a_8_24# AND2X1_LOC_53/Y 0.00fF
C20500 OR2X1_LOC_318/Y OR2X1_LOC_532/B 0.00fF
C20501 OR2X1_LOC_46/A AND2X1_LOC_403/B 0.01fF
C20502 AND2X1_LOC_584/a_8_24# AND2X1_LOC_1/Y 0.01fF
C20503 OR2X1_LOC_543/A OR2X1_LOC_543/a_8_216# 0.01fF
C20504 AND2X1_LOC_660/A OR2X1_LOC_275/Y 0.03fF
C20505 AND2X1_LOC_576/Y AND2X1_LOC_523/Y 0.01fF
C20506 AND2X1_LOC_70/Y OR2X1_LOC_247/Y 0.09fF
C20507 OR2X1_LOC_599/Y AND2X1_LOC_434/Y 0.08fF
C20508 AND2X1_LOC_42/B AND2X1_LOC_3/Y 0.06fF
C20509 OR2X1_LOC_278/A OR2X1_LOC_85/A 0.10fF
C20510 OR2X1_LOC_18/Y AND2X1_LOC_845/Y 0.00fF
C20511 OR2X1_LOC_604/A AND2X1_LOC_222/Y 0.03fF
C20512 AND2X1_LOC_273/a_8_24# OR2X1_LOC_593/B 0.01fF
C20513 AND2X1_LOC_514/Y AND2X1_LOC_354/B 0.85fF
C20514 AND2X1_LOC_31/Y OR2X1_LOC_641/A 0.03fF
C20515 OR2X1_LOC_3/Y OR2X1_LOC_131/Y 0.04fF
C20516 OR2X1_LOC_417/Y OR2X1_LOC_26/Y 0.00fF
C20517 AND2X1_LOC_536/a_36_24# D_INPUT_0 0.00fF
C20518 OR2X1_LOC_291/Y OR2X1_LOC_26/Y 0.03fF
C20519 OR2X1_LOC_185/Y AND2X1_LOC_48/A 0.02fF
C20520 OR2X1_LOC_681/Y OR2X1_LOC_7/A 0.02fF
C20521 OR2X1_LOC_121/B OR2X1_LOC_99/Y 0.04fF
C20522 AND2X1_LOC_81/B OR2X1_LOC_814/A 0.03fF
C20523 OR2X1_LOC_479/Y OR2X1_LOC_794/a_36_216# 0.00fF
C20524 OR2X1_LOC_79/A AND2X1_LOC_78/a_36_24# 0.00fF
C20525 AND2X1_LOC_31/Y OR2X1_LOC_733/A 0.01fF
C20526 OR2X1_LOC_786/Y OR2X1_LOC_721/Y 0.03fF
C20527 OR2X1_LOC_527/Y OR2X1_LOC_89/A 0.84fF
C20528 OR2X1_LOC_46/A OR2X1_LOC_44/Y 0.03fF
C20529 OR2X1_LOC_532/B OR2X1_LOC_805/A 0.19fF
C20530 OR2X1_LOC_525/Y AND2X1_LOC_796/Y 0.00fF
C20531 OR2X1_LOC_70/Y AND2X1_LOC_390/B 0.58fF
C20532 AND2X1_LOC_717/a_36_24# OR2X1_LOC_95/Y 0.00fF
C20533 OR2X1_LOC_40/Y OR2X1_LOC_80/A 0.01fF
C20534 AND2X1_LOC_489/a_8_24# AND2X1_LOC_657/A 0.01fF
C20535 OR2X1_LOC_83/A OR2X1_LOC_54/Y 0.00fF
C20536 OR2X1_LOC_417/Y OR2X1_LOC_89/A 0.03fF
C20537 OR2X1_LOC_728/B OR2X1_LOC_715/A 0.14fF
C20538 OR2X1_LOC_427/A OR2X1_LOC_615/Y 0.24fF
C20539 OR2X1_LOC_771/B AND2X1_LOC_44/Y 0.03fF
C20540 OR2X1_LOC_331/A OR2X1_LOC_331/Y 0.11fF
C20541 OR2X1_LOC_66/A OR2X1_LOC_68/B 0.21fF
C20542 OR2X1_LOC_639/B OR2X1_LOC_639/a_8_216# 0.07fF
C20543 OR2X1_LOC_657/a_8_216# OR2X1_LOC_244/A 0.03fF
C20544 VDD OR2X1_LOC_534/Y 0.12fF
C20545 OR2X1_LOC_11/Y OR2X1_LOC_408/Y 0.02fF
C20546 OR2X1_LOC_439/B OR2X1_LOC_303/B 0.13fF
C20547 OR2X1_LOC_416/Y OR2X1_LOC_7/A 0.00fF
C20548 AND2X1_LOC_342/a_36_24# OR2X1_LOC_54/Y 0.00fF
C20549 AND2X1_LOC_181/Y OR2X1_LOC_437/A 0.01fF
C20550 OR2X1_LOC_754/A OR2X1_LOC_615/a_8_216# 0.13fF
C20551 AND2X1_LOC_44/Y OR2X1_LOC_209/A 0.28fF
C20552 AND2X1_LOC_36/Y OR2X1_LOC_577/Y 0.04fF
C20553 INPUT_1 AND2X1_LOC_838/a_8_24# 0.01fF
C20554 OR2X1_LOC_59/Y OR2X1_LOC_153/a_8_216# 0.02fF
C20555 OR2X1_LOC_848/A OR2X1_LOC_770/a_8_216# 0.41fF
C20556 VDD OR2X1_LOC_365/a_8_216# 0.00fF
C20557 OR2X1_LOC_296/a_8_216# OR2X1_LOC_62/B 0.01fF
C20558 OR2X1_LOC_70/Y OR2X1_LOC_431/Y 0.01fF
C20559 AND2X1_LOC_171/a_36_24# AND2X1_LOC_48/A 0.01fF
C20560 AND2X1_LOC_227/Y OR2X1_LOC_44/Y 0.06fF
C20561 AND2X1_LOC_866/A OR2X1_LOC_6/A 0.23fF
C20562 OR2X1_LOC_827/Y INPUT_1 0.03fF
C20563 AND2X1_LOC_390/B AND2X1_LOC_538/a_8_24# 0.03fF
C20564 OR2X1_LOC_375/A OR2X1_LOC_786/Y 0.57fF
C20565 OR2X1_LOC_831/A OR2X1_LOC_723/B 0.86fF
C20566 OR2X1_LOC_308/Y OR2X1_LOC_713/A 0.02fF
C20567 OR2X1_LOC_703/A OR2X1_LOC_353/a_8_216# 0.01fF
C20568 D_INPUT_3 OR2X1_LOC_26/Y 0.08fF
C20569 AND2X1_LOC_539/Y AND2X1_LOC_799/a_8_24# 0.01fF
C20570 OR2X1_LOC_696/A AND2X1_LOC_802/Y 0.05fF
C20571 OR2X1_LOC_19/B OR2X1_LOC_415/A 0.83fF
C20572 OR2X1_LOC_426/B OR2X1_LOC_13/B 0.67fF
C20573 OR2X1_LOC_502/A AND2X1_LOC_432/a_8_24# 0.04fF
C20574 OR2X1_LOC_602/Y OR2X1_LOC_777/B 0.46fF
C20575 AND2X1_LOC_566/Y AND2X1_LOC_170/B 0.02fF
C20576 AND2X1_LOC_543/Y AND2X1_LOC_457/a_8_24# 0.01fF
C20577 AND2X1_LOC_64/Y OR2X1_LOC_318/A 0.01fF
C20578 D_INPUT_3 OR2X1_LOC_89/A 0.04fF
C20579 AND2X1_LOC_41/A OR2X1_LOC_446/B 0.07fF
C20580 OR2X1_LOC_91/Y AND2X1_LOC_804/a_8_24# 0.01fF
C20581 OR2X1_LOC_390/B OR2X1_LOC_390/A 0.23fF
C20582 OR2X1_LOC_648/B OR2X1_LOC_333/A 0.19fF
C20583 OR2X1_LOC_484/a_8_216# OR2X1_LOC_142/a_8_216# 0.47fF
C20584 AND2X1_LOC_715/Y AND2X1_LOC_802/Y 0.00fF
C20585 OR2X1_LOC_648/a_8_216# OR2X1_LOC_750/A 0.01fF
C20586 OR2X1_LOC_379/Y AND2X1_LOC_31/Y 0.03fF
C20587 OR2X1_LOC_47/Y OR2X1_LOC_438/a_8_216# 0.03fF
C20588 OR2X1_LOC_824/a_36_216# D_INPUT_3 0.00fF
C20589 AND2X1_LOC_64/Y OR2X1_LOC_151/A 0.43fF
C20590 OR2X1_LOC_154/A OR2X1_LOC_358/A 0.03fF
C20591 OR2X1_LOC_165/Y OR2X1_LOC_437/A 0.02fF
C20592 OR2X1_LOC_36/Y AND2X1_LOC_647/Y 0.06fF
C20593 AND2X1_LOC_514/Y AND2X1_LOC_863/Y 0.81fF
C20594 OR2X1_LOC_739/A OR2X1_LOC_739/a_8_216# 0.18fF
C20595 OR2X1_LOC_135/a_8_216# OR2X1_LOC_428/A 0.03fF
C20596 AND2X1_LOC_572/A AND2X1_LOC_657/A 0.14fF
C20597 OR2X1_LOC_160/B OR2X1_LOC_140/B 0.03fF
C20598 AND2X1_LOC_557/Y AND2X1_LOC_563/Y 0.09fF
C20599 AND2X1_LOC_477/Y AND2X1_LOC_794/a_8_24# 0.02fF
C20600 OR2X1_LOC_74/A OR2X1_LOC_419/Y 0.17fF
C20601 OR2X1_LOC_36/Y AND2X1_LOC_783/a_8_24# 0.01fF
C20602 AND2X1_LOC_40/Y OR2X1_LOC_723/B 1.16fF
C20603 OR2X1_LOC_287/B OR2X1_LOC_675/Y 0.03fF
C20604 OR2X1_LOC_693/a_8_216# OR2X1_LOC_692/Y 0.02fF
C20605 AND2X1_LOC_457/a_8_24# OR2X1_LOC_322/Y 0.02fF
C20606 OR2X1_LOC_599/A AND2X1_LOC_783/a_36_24# 0.01fF
C20607 AND2X1_LOC_476/Y AND2X1_LOC_786/Y 0.04fF
C20608 OR2X1_LOC_833/a_8_216# AND2X1_LOC_36/Y 0.01fF
C20609 OR2X1_LOC_89/A AND2X1_LOC_656/a_8_24# 0.01fF
C20610 AND2X1_LOC_476/Y OR2X1_LOC_323/a_8_216# 0.05fF
C20611 OR2X1_LOC_755/A OR2X1_LOC_815/Y 0.01fF
C20612 AND2X1_LOC_91/B OR2X1_LOC_648/A 0.16fF
C20613 AND2X1_LOC_787/A OR2X1_LOC_600/A 0.05fF
C20614 AND2X1_LOC_228/Y OR2X1_LOC_437/A 0.16fF
C20615 OR2X1_LOC_95/Y OR2X1_LOC_751/A 0.04fF
C20616 AND2X1_LOC_22/Y OR2X1_LOC_468/A 0.09fF
C20617 AND2X1_LOC_674/a_36_24# OR2X1_LOC_374/Y 0.00fF
C20618 OR2X1_LOC_691/Y OR2X1_LOC_800/Y 0.01fF
C20619 AND2X1_LOC_473/Y OR2X1_LOC_56/A 1.10fF
C20620 AND2X1_LOC_217/Y OR2X1_LOC_12/Y 0.00fF
C20621 VDD AND2X1_LOC_785/Y 0.21fF
C20622 AND2X1_LOC_96/a_8_24# OR2X1_LOC_415/Y 0.17fF
C20623 OR2X1_LOC_158/A AND2X1_LOC_346/a_8_24# 0.02fF
C20624 OR2X1_LOC_676/Y OR2X1_LOC_161/B 0.01fF
C20625 OR2X1_LOC_409/B OR2X1_LOC_409/a_8_216# 0.07fF
C20626 OR2X1_LOC_51/Y OR2X1_LOC_744/a_36_216# 0.00fF
C20627 AND2X1_LOC_593/a_36_24# OR2X1_LOC_12/Y 0.01fF
C20628 OR2X1_LOC_831/A AND2X1_LOC_300/a_36_24# 0.00fF
C20629 OR2X1_LOC_74/A OR2X1_LOC_152/A 0.03fF
C20630 OR2X1_LOC_816/A OR2X1_LOC_56/A 0.01fF
C20631 OR2X1_LOC_709/A AND2X1_LOC_18/Y 0.03fF
C20632 OR2X1_LOC_619/Y OR2X1_LOC_320/a_36_216# 0.01fF
C20633 OR2X1_LOC_201/Y AND2X1_LOC_31/Y 0.01fF
C20634 OR2X1_LOC_687/Y OR2X1_LOC_515/Y 0.12fF
C20635 OR2X1_LOC_76/A OR2X1_LOC_675/Y 0.81fF
C20636 OR2X1_LOC_671/Y OR2X1_LOC_96/Y 0.09fF
C20637 OR2X1_LOC_78/A AND2X1_LOC_627/a_8_24# 0.01fF
C20638 OR2X1_LOC_389/A OR2X1_LOC_390/A 0.01fF
C20639 OR2X1_LOC_778/Y OR2X1_LOC_704/a_8_216# 0.30fF
C20640 AND2X1_LOC_592/Y AND2X1_LOC_713/Y 0.01fF
C20641 OR2X1_LOC_375/A OR2X1_LOC_199/B 0.05fF
C20642 OR2X1_LOC_6/B OR2X1_LOC_786/A 0.06fF
C20643 OR2X1_LOC_678/a_8_216# AND2X1_LOC_44/Y 0.01fF
C20644 OR2X1_LOC_834/A OR2X1_LOC_161/B 0.01fF
C20645 OR2X1_LOC_696/A AND2X1_LOC_832/a_36_24# 0.01fF
C20646 OR2X1_LOC_585/A OR2X1_LOC_437/A 0.26fF
C20647 OR2X1_LOC_676/Y OR2X1_LOC_514/a_36_216# 0.01fF
C20648 OR2X1_LOC_482/Y OR2X1_LOC_666/a_8_216# 0.01fF
C20649 AND2X1_LOC_566/B AND2X1_LOC_335/Y 0.02fF
C20650 AND2X1_LOC_857/Y OR2X1_LOC_230/Y 0.21fF
C20651 AND2X1_LOC_388/Y VDD 0.06fF
C20652 OR2X1_LOC_158/A AND2X1_LOC_447/Y 0.00fF
C20653 OR2X1_LOC_485/A OR2X1_LOC_150/a_8_216# 0.01fF
C20654 AND2X1_LOC_850/A AND2X1_LOC_244/A 1.35fF
C20655 VDD AND2X1_LOC_625/a_8_24# 0.00fF
C20656 OR2X1_LOC_535/A OR2X1_LOC_78/B 0.12fF
C20657 AND2X1_LOC_212/A OR2X1_LOC_56/A 0.03fF
C20658 VDD AND2X1_LOC_500/B 0.17fF
C20659 AND2X1_LOC_595/a_8_24# OR2X1_LOC_66/A 0.05fF
C20660 OR2X1_LOC_158/A OR2X1_LOC_380/Y 0.03fF
C20661 AND2X1_LOC_103/a_8_24# OR2X1_LOC_113/B 0.01fF
C20662 OR2X1_LOC_285/a_8_216# OR2X1_LOC_758/a_8_216# 0.47fF
C20663 OR2X1_LOC_743/A OR2X1_LOC_13/B 0.18fF
C20664 OR2X1_LOC_427/A AND2X1_LOC_242/B 0.07fF
C20665 AND2X1_LOC_7/B OR2X1_LOC_714/Y 0.01fF
C20666 AND2X1_LOC_721/a_8_24# OR2X1_LOC_428/A 0.16fF
C20667 OR2X1_LOC_229/a_8_216# AND2X1_LOC_857/Y 0.04fF
C20668 AND2X1_LOC_70/Y AND2X1_LOC_18/Y 3.98fF
C20669 OR2X1_LOC_61/A OR2X1_LOC_61/B 0.07fF
C20670 AND2X1_LOC_568/B AND2X1_LOC_436/Y 0.00fF
C20671 OR2X1_LOC_524/Y AND2X1_LOC_476/Y 0.15fF
C20672 OR2X1_LOC_302/B AND2X1_LOC_110/Y 0.01fF
C20673 OR2X1_LOC_273/Y OR2X1_LOC_300/Y 0.01fF
C20674 AND2X1_LOC_11/Y AND2X1_LOC_44/Y 0.03fF
C20675 AND2X1_LOC_850/Y OR2X1_LOC_816/A 0.07fF
C20676 OR2X1_LOC_186/Y OR2X1_LOC_147/B 0.07fF
C20677 AND2X1_LOC_61/a_8_24# OR2X1_LOC_59/Y 0.01fF
C20678 OR2X1_LOC_702/A AND2X1_LOC_36/Y 0.00fF
C20679 OR2X1_LOC_218/Y OR2X1_LOC_228/Y 0.01fF
C20680 OR2X1_LOC_44/Y OR2X1_LOC_748/a_8_216# 0.01fF
C20681 OR2X1_LOC_663/A OR2X1_LOC_772/A 0.09fF
C20682 OR2X1_LOC_286/Y OR2X1_LOC_580/B 0.03fF
C20683 OR2X1_LOC_201/a_8_216# AND2X1_LOC_31/Y 0.01fF
C20684 AND2X1_LOC_74/a_8_24# OR2X1_LOC_486/Y 0.03fF
C20685 AND2X1_LOC_366/A OR2X1_LOC_494/Y 0.03fF
C20686 OR2X1_LOC_121/B OR2X1_LOC_788/B 0.01fF
C20687 OR2X1_LOC_130/A OR2X1_LOC_227/B 0.02fF
C20688 OR2X1_LOC_186/Y OR2X1_LOC_317/A 0.01fF
C20689 AND2X1_LOC_366/A AND2X1_LOC_363/Y 0.19fF
C20690 AND2X1_LOC_621/Y AND2X1_LOC_213/B 0.02fF
C20691 OR2X1_LOC_619/Y AND2X1_LOC_210/a_36_24# 0.00fF
C20692 OR2X1_LOC_246/A OR2X1_LOC_13/B 0.18fF
C20693 OR2X1_LOC_87/A AND2X1_LOC_226/a_36_24# 0.02fF
C20694 INPUT_0 AND2X1_LOC_691/a_8_24# 0.01fF
C20695 OR2X1_LOC_147/B OR2X1_LOC_726/A 0.05fF
C20696 OR2X1_LOC_744/A OR2X1_LOC_59/Y 10.06fF
C20697 AND2X1_LOC_391/a_8_24# OR2X1_LOC_600/A 0.03fF
C20698 OR2X1_LOC_287/a_36_216# OR2X1_LOC_366/Y 0.01fF
C20699 OR2X1_LOC_151/A AND2X1_LOC_321/a_36_24# 0.01fF
C20700 AND2X1_LOC_40/Y OR2X1_LOC_676/a_8_216# 0.01fF
C20701 OR2X1_LOC_99/a_8_216# AND2X1_LOC_7/B 0.06fF
C20702 OR2X1_LOC_375/A AND2X1_LOC_255/a_8_24# 0.02fF
C20703 OR2X1_LOC_800/A OR2X1_LOC_691/Y 0.01fF
C20704 OR2X1_LOC_158/A OR2X1_LOC_109/Y 0.03fF
C20705 OR2X1_LOC_333/B OR2X1_LOC_333/a_36_216# 0.02fF
C20706 OR2X1_LOC_476/B AND2X1_LOC_36/Y 0.08fF
C20707 OR2X1_LOC_497/Y AND2X1_LOC_242/a_8_24# 0.05fF
C20708 OR2X1_LOC_659/B OR2X1_LOC_576/A 0.02fF
C20709 AND2X1_LOC_47/Y OR2X1_LOC_366/Y 0.03fF
C20710 AND2X1_LOC_566/B OR2X1_LOC_619/Y 0.03fF
C20711 OR2X1_LOC_205/Y OR2X1_LOC_641/B 0.04fF
C20712 AND2X1_LOC_861/B AND2X1_LOC_663/A 0.10fF
C20713 AND2X1_LOC_97/a_8_24# AND2X1_LOC_243/Y 0.02fF
C20714 OR2X1_LOC_483/a_8_216# OR2X1_LOC_161/B 0.01fF
C20715 OR2X1_LOC_207/B OR2X1_LOC_185/Y 0.03fF
C20716 AND2X1_LOC_22/Y OR2X1_LOC_449/B 0.03fF
C20717 OR2X1_LOC_158/A AND2X1_LOC_448/Y 0.01fF
C20718 AND2X1_LOC_776/a_8_24# AND2X1_LOC_486/Y 0.03fF
C20719 OR2X1_LOC_421/A OR2X1_LOC_432/a_36_216# 0.00fF
C20720 OR2X1_LOC_650/Y AND2X1_LOC_36/Y 1.03fF
C20721 AND2X1_LOC_471/Y AND2X1_LOC_477/a_8_24# 0.06fF
C20722 AND2X1_LOC_810/A OR2X1_LOC_36/Y 0.04fF
C20723 VDD AND2X1_LOC_364/A 0.03fF
C20724 OR2X1_LOC_640/A AND2X1_LOC_92/Y 0.02fF
C20725 OR2X1_LOC_6/B OR2X1_LOC_624/A 0.10fF
C20726 OR2X1_LOC_102/a_36_216# AND2X1_LOC_342/Y 0.01fF
C20727 AND2X1_LOC_359/B OR2X1_LOC_12/Y 0.01fF
C20728 OR2X1_LOC_644/a_8_216# AND2X1_LOC_36/Y 0.01fF
C20729 OR2X1_LOC_769/B AND2X1_LOC_40/Y 0.01fF
C20730 AND2X1_LOC_634/a_8_24# AND2X1_LOC_219/A 0.04fF
C20731 OR2X1_LOC_127/a_8_216# OR2X1_LOC_600/A 0.02fF
C20732 AND2X1_LOC_31/Y OR2X1_LOC_741/A 0.01fF
C20733 AND2X1_LOC_363/a_8_24# AND2X1_LOC_348/Y 0.01fF
C20734 AND2X1_LOC_706/Y OR2X1_LOC_433/a_36_216# 0.01fF
C20735 OR2X1_LOC_45/Y OR2X1_LOC_56/A 0.52fF
C20736 AND2X1_LOC_563/a_8_24# AND2X1_LOC_563/A 0.10fF
C20737 AND2X1_LOC_403/B AND2X1_LOC_403/a_8_24# 0.04fF
C20738 AND2X1_LOC_339/a_8_24# OR2X1_LOC_16/A 0.01fF
C20739 OR2X1_LOC_476/B OR2X1_LOC_334/A 0.00fF
C20740 OR2X1_LOC_354/A AND2X1_LOC_167/a_36_24# 0.00fF
C20741 OR2X1_LOC_631/B OR2X1_LOC_719/B 0.03fF
C20742 VDD OR2X1_LOC_807/A 0.04fF
C20743 AND2X1_LOC_754/a_8_24# OR2X1_LOC_269/B 0.01fF
C20744 OR2X1_LOC_539/a_8_216# VDD 0.00fF
C20745 OR2X1_LOC_159/a_8_216# OR2X1_LOC_6/A 0.02fF
C20746 OR2X1_LOC_447/Y OR2X1_LOC_714/a_8_216# 0.01fF
C20747 OR2X1_LOC_485/A AND2X1_LOC_774/A 0.01fF
C20748 OR2X1_LOC_40/Y OR2X1_LOC_6/A 0.13fF
C20749 VDD AND2X1_LOC_572/A 0.15fF
C20750 OR2X1_LOC_36/Y AND2X1_LOC_254/a_8_24# 0.08fF
C20751 OR2X1_LOC_8/Y AND2X1_LOC_838/Y 0.01fF
C20752 OR2X1_LOC_696/A INPUT_1 0.03fF
C20753 AND2X1_LOC_784/A AND2X1_LOC_357/A 0.02fF
C20754 OR2X1_LOC_377/A OR2X1_LOC_78/A 0.33fF
C20755 OR2X1_LOC_36/Y AND2X1_LOC_860/A 0.07fF
C20756 OR2X1_LOC_193/Y AND2X1_LOC_18/Y 0.18fF
C20757 OR2X1_LOC_423/a_36_216# OR2X1_LOC_421/Y 0.01fF
C20758 OR2X1_LOC_481/A OR2X1_LOC_428/A 0.06fF
C20759 AND2X1_LOC_807/Y OR2X1_LOC_56/A 0.07fF
C20760 OR2X1_LOC_864/A OR2X1_LOC_641/A 0.05fF
C20761 OR2X1_LOC_298/a_8_216# AND2X1_LOC_654/Y 0.03fF
C20762 AND2X1_LOC_710/a_8_24# AND2X1_LOC_710/Y 0.01fF
C20763 OR2X1_LOC_177/Y OR2X1_LOC_74/A 0.02fF
C20764 AND2X1_LOC_721/Y AND2X1_LOC_849/A 1.01fF
C20765 AND2X1_LOC_22/Y OR2X1_LOC_121/B 0.07fF
C20766 OR2X1_LOC_644/B VDD 0.00fF
C20767 VDD OR2X1_LOC_464/B -0.00fF
C20768 OR2X1_LOC_557/A OR2X1_LOC_768/a_8_216# 0.01fF
C20769 AND2X1_LOC_576/Y AND2X1_LOC_657/Y 0.10fF
C20770 OR2X1_LOC_831/a_8_216# AND2X1_LOC_92/Y 0.03fF
C20771 AND2X1_LOC_772/a_8_24# AND2X1_LOC_657/A 0.01fF
C20772 AND2X1_LOC_364/Y AND2X1_LOC_655/A 0.48fF
C20773 AND2X1_LOC_191/B AND2X1_LOC_576/Y 0.07fF
C20774 AND2X1_LOC_394/a_8_24# OR2X1_LOC_235/B 0.03fF
C20775 OR2X1_LOC_160/A AND2X1_LOC_71/a_8_24# 0.04fF
C20776 AND2X1_LOC_707/Y AND2X1_LOC_687/B 0.16fF
C20777 AND2X1_LOC_578/A AND2X1_LOC_476/Y 0.07fF
C20778 AND2X1_LOC_512/Y AND2X1_LOC_436/B 0.03fF
C20779 AND2X1_LOC_40/Y OR2X1_LOC_812/B 0.14fF
C20780 AND2X1_LOC_840/B OR2X1_LOC_59/Y 0.07fF
C20781 OR2X1_LOC_203/Y OR2X1_LOC_78/A 0.07fF
C20782 AND2X1_LOC_330/a_8_24# OR2X1_LOC_26/Y 0.03fF
C20783 OR2X1_LOC_691/Y OR2X1_LOC_19/B 0.04fF
C20784 OR2X1_LOC_318/A OR2X1_LOC_206/A 0.98fF
C20785 AND2X1_LOC_99/A AND2X1_LOC_99/a_36_24# 0.01fF
C20786 OR2X1_LOC_45/B OR2X1_LOC_46/A 0.24fF
C20787 OR2X1_LOC_744/A OR2X1_LOC_433/a_8_216# 0.01fF
C20788 OR2X1_LOC_144/Y AND2X1_LOC_621/Y 0.19fF
C20789 OR2X1_LOC_604/A OR2X1_LOC_74/A 0.23fF
C20790 OR2X1_LOC_662/a_8_216# OR2X1_LOC_87/A 0.01fF
C20791 AND2X1_LOC_691/a_8_24# OR2X1_LOC_690/A 0.02fF
C20792 AND2X1_LOC_602/a_36_24# AND2X1_LOC_447/Y 0.01fF
C20793 OR2X1_LOC_74/a_8_216# OR2X1_LOC_59/Y 0.02fF
C20794 OR2X1_LOC_840/A OR2X1_LOC_539/Y 0.16fF
C20795 OR2X1_LOC_653/a_8_216# AND2X1_LOC_18/Y 0.01fF
C20796 AND2X1_LOC_217/Y OR2X1_LOC_272/Y 0.16fF
C20797 OR2X1_LOC_139/A D_INPUT_0 0.16fF
C20798 AND2X1_LOC_484/a_8_24# OR2X1_LOC_726/A 0.01fF
C20799 OR2X1_LOC_49/A OR2X1_LOC_77/a_8_216# 0.01fF
C20800 AND2X1_LOC_95/Y OR2X1_LOC_856/B 0.14fF
C20801 OR2X1_LOC_92/Y OR2X1_LOC_65/B 0.02fF
C20802 AND2X1_LOC_41/A AND2X1_LOC_56/B 1.56fF
C20803 VDD OR2X1_LOC_3/Y 1.01fF
C20804 OR2X1_LOC_417/Y AND2X1_LOC_605/a_8_24# 0.01fF
C20805 OR2X1_LOC_589/A AND2X1_LOC_307/Y 0.03fF
C20806 OR2X1_LOC_459/A OR2X1_LOC_36/Y 0.03fF
C20807 OR2X1_LOC_720/B OR2X1_LOC_721/a_36_216# 0.00fF
C20808 OR2X1_LOC_805/A OR2X1_LOC_734/a_8_216# 0.06fF
C20809 OR2X1_LOC_600/A OR2X1_LOC_817/Y 0.01fF
C20810 OR2X1_LOC_71/Y OR2X1_LOC_428/A 0.02fF
C20811 OR2X1_LOC_167/a_8_216# OR2X1_LOC_601/a_8_216# 0.47fF
C20812 AND2X1_LOC_722/A OR2X1_LOC_44/Y 0.01fF
C20813 VDD AND2X1_LOC_631/Y 0.04fF
C20814 OR2X1_LOC_485/A AND2X1_LOC_434/a_8_24# 0.01fF
C20815 OR2X1_LOC_697/a_8_216# OR2X1_LOC_52/B 0.04fF
C20816 AND2X1_LOC_719/a_8_24# OR2X1_LOC_59/Y 0.01fF
C20817 OR2X1_LOC_382/Y OR2X1_LOC_43/A 0.00fF
C20818 OR2X1_LOC_375/A OR2X1_LOC_725/B 0.00fF
C20819 OR2X1_LOC_833/Y OR2X1_LOC_814/A 0.01fF
C20820 OR2X1_LOC_604/A OR2X1_LOC_261/A -0.01fF
C20821 OR2X1_LOC_282/Y AND2X1_LOC_285/Y 0.80fF
C20822 OR2X1_LOC_108/Y AND2X1_LOC_523/Y 0.07fF
C20823 OR2X1_LOC_160/B OR2X1_LOC_719/A 0.02fF
C20824 OR2X1_LOC_404/Y AND2X1_LOC_18/Y 0.00fF
C20825 OR2X1_LOC_759/A OR2X1_LOC_755/A 0.01fF
C20826 OR2X1_LOC_532/B OR2X1_LOC_580/B 0.03fF
C20827 AND2X1_LOC_729/Y OR2X1_LOC_48/B 0.05fF
C20828 OR2X1_LOC_45/B AND2X1_LOC_227/Y 0.11fF
C20829 AND2X1_LOC_142/a_8_24# OR2X1_LOC_87/A 0.04fF
C20830 AND2X1_LOC_713/Y AND2X1_LOC_712/B 0.01fF
C20831 AND2X1_LOC_72/Y OR2X1_LOC_203/a_8_216# 0.05fF
C20832 OR2X1_LOC_105/Y OR2X1_LOC_643/A 0.02fF
C20833 OR2X1_LOC_71/Y OR2X1_LOC_595/A 0.04fF
C20834 OR2X1_LOC_768/A OR2X1_LOC_624/B 0.00fF
C20835 OR2X1_LOC_6/B OR2X1_LOC_54/Y 0.30fF
C20836 OR2X1_LOC_271/Y OR2X1_LOC_92/Y 0.06fF
C20837 AND2X1_LOC_689/a_36_24# OR2X1_LOC_66/A 0.00fF
C20838 INPUT_0 AND2X1_LOC_42/B 0.08fF
C20839 GATE_662 GATE_579 0.02fF
C20840 AND2X1_LOC_12/Y AND2X1_LOC_305/a_36_24# 0.00fF
C20841 AND2X1_LOC_465/a_36_24# OR2X1_LOC_744/A 0.01fF
C20842 OR2X1_LOC_181/A OR2X1_LOC_181/a_8_216# 0.47fF
C20843 OR2X1_LOC_70/Y OR2X1_LOC_744/A 0.34fF
C20844 AND2X1_LOC_2/Y AND2X1_LOC_1/Y 0.11fF
C20845 OR2X1_LOC_663/A AND2X1_LOC_3/Y 0.03fF
C20846 OR2X1_LOC_680/A AND2X1_LOC_468/B 0.00fF
C20847 OR2X1_LOC_432/a_8_216# OR2X1_LOC_36/Y 0.01fF
C20848 VDD OR2X1_LOC_582/Y 0.04fF
C20849 AND2X1_LOC_410/a_8_24# OR2X1_LOC_46/A 0.01fF
C20850 AND2X1_LOC_658/A OR2X1_LOC_253/a_8_216# 0.03fF
C20851 AND2X1_LOC_374/a_8_24# OR2X1_LOC_312/Y 0.01fF
C20852 OR2X1_LOC_237/a_8_216# OR2X1_LOC_237/Y 0.01fF
C20853 D_INPUT_0 OR2X1_LOC_131/a_8_216# 0.04fF
C20854 AND2X1_LOC_784/A OR2X1_LOC_48/B 0.09fF
C20855 OR2X1_LOC_631/a_8_216# OR2X1_LOC_631/B 0.02fF
C20856 OR2X1_LOC_805/a_8_216# OR2X1_LOC_269/B 0.02fF
C20857 VDD AND2X1_LOC_133/a_8_24# -0.00fF
C20858 OR2X1_LOC_648/B OR2X1_LOC_532/B 0.08fF
C20859 OR2X1_LOC_468/Y OR2X1_LOC_739/A 0.03fF
C20860 OR2X1_LOC_847/A OR2X1_LOC_847/B 0.17fF
C20861 OR2X1_LOC_400/a_8_216# OR2X1_LOC_557/A 0.01fF
C20862 OR2X1_LOC_3/Y OR2X1_LOC_689/A 0.02fF
C20863 AND2X1_LOC_727/A OR2X1_LOC_56/A 0.06fF
C20864 AND2X1_LOC_16/a_8_24# OR2X1_LOC_155/A 0.01fF
C20865 OR2X1_LOC_326/a_8_216# OR2X1_LOC_121/B 0.01fF
C20866 OR2X1_LOC_362/B OR2X1_LOC_269/B 0.02fF
C20867 AND2X1_LOC_514/Y OR2X1_LOC_744/A 0.07fF
C20868 OR2X1_LOC_204/Y OR2X1_LOC_375/A 0.03fF
C20869 AND2X1_LOC_452/Y OR2X1_LOC_418/Y 0.05fF
C20870 OR2X1_LOC_405/A OR2X1_LOC_810/A 0.13fF
C20871 AND2X1_LOC_778/a_8_24# OR2X1_LOC_18/Y 0.02fF
C20872 AND2X1_LOC_502/a_8_24# OR2X1_LOC_497/Y 0.01fF
C20873 OR2X1_LOC_185/A OR2X1_LOC_592/a_8_216# 0.06fF
C20874 AND2X1_LOC_73/a_8_24# OR2X1_LOC_54/Y 0.06fF
C20875 AND2X1_LOC_841/a_8_24# AND2X1_LOC_476/Y 0.00fF
C20876 AND2X1_LOC_640/Y OR2X1_LOC_46/a_8_216# 0.06fF
C20877 OR2X1_LOC_276/B AND2X1_LOC_275/a_8_24# 0.02fF
C20878 OR2X1_LOC_662/A AND2X1_LOC_8/Y 0.03fF
C20879 VDD AND2X1_LOC_53/Y 0.21fF
C20880 AND2X1_LOC_769/a_8_24# OR2X1_LOC_48/B 0.02fF
C20881 OR2X1_LOC_468/Y OR2X1_LOC_798/a_8_216# 0.39fF
C20882 OR2X1_LOC_377/A OR2X1_LOC_155/A 0.01fF
C20883 OR2X1_LOC_786/Y OR2X1_LOC_549/A 0.01fF
C20884 OR2X1_LOC_748/A AND2X1_LOC_848/a_36_24# 0.00fF
C20885 OR2X1_LOC_557/A OR2X1_LOC_847/A 0.05fF
C20886 AND2X1_LOC_580/A AND2X1_LOC_859/Y 0.07fF
C20887 AND2X1_LOC_769/a_8_24# OR2X1_LOC_18/Y 0.02fF
C20888 OR2X1_LOC_808/B OR2X1_LOC_76/A 0.11fF
C20889 OR2X1_LOC_36/Y AND2X1_LOC_287/Y 0.03fF
C20890 OR2X1_LOC_648/A AND2X1_LOC_600/a_36_24# 0.00fF
C20891 OR2X1_LOC_297/a_36_216# AND2X1_LOC_663/B 0.00fF
C20892 OR2X1_LOC_6/B OR2X1_LOC_276/a_8_216# 0.04fF
C20893 AND2X1_LOC_41/Y OR2X1_LOC_195/a_8_216# 0.07fF
C20894 OR2X1_LOC_369/Y OR2X1_LOC_417/A -0.00fF
C20895 OR2X1_LOC_19/B OR2X1_LOC_394/a_36_216# 0.01fF
C20896 OR2X1_LOC_599/A OR2X1_LOC_44/Y 0.09fF
C20897 OR2X1_LOC_674/Y AND2X1_LOC_500/B 0.01fF
C20898 AND2X1_LOC_541/Y OR2X1_LOC_47/Y 0.00fF
C20899 OR2X1_LOC_631/B AND2X1_LOC_56/B 0.00fF
C20900 OR2X1_LOC_553/A OR2X1_LOC_553/a_8_216# 0.04fF
C20901 AND2X1_LOC_214/A OR2X1_LOC_7/Y 0.02fF
C20902 OR2X1_LOC_219/B OR2X1_LOC_219/a_36_216# 0.01fF
C20903 AND2X1_LOC_103/a_8_24# OR2X1_LOC_532/B 0.03fF
C20904 OR2X1_LOC_468/Y OR2X1_LOC_269/B 0.03fF
C20905 OR2X1_LOC_598/A OR2X1_LOC_548/B 0.00fF
C20906 OR2X1_LOC_195/A AND2X1_LOC_43/B 0.14fF
C20907 AND2X1_LOC_738/B OR2X1_LOC_95/Y 0.05fF
C20908 OR2X1_LOC_95/Y OR2X1_LOC_56/A 0.45fF
C20909 OR2X1_LOC_642/a_36_216# AND2X1_LOC_8/Y 0.00fF
C20910 INPUT_1 AND2X1_LOC_819/a_8_24# 0.01fF
C20911 OR2X1_LOC_176/Y AND2X1_LOC_222/Y 0.00fF
C20912 OR2X1_LOC_31/Y OR2X1_LOC_59/Y 2.28fF
C20913 OR2X1_LOC_70/A AND2X1_LOC_639/B 0.07fF
C20914 VDD OR2X1_LOC_673/A 0.26fF
C20915 VDD OR2X1_LOC_223/A 0.41fF
C20916 AND2X1_LOC_372/a_8_24# OR2X1_LOC_532/B 0.01fF
C20917 OR2X1_LOC_7/A OR2X1_LOC_6/A 0.26fF
C20918 AND2X1_LOC_576/a_36_24# AND2X1_LOC_489/Y 0.00fF
C20919 OR2X1_LOC_819/a_8_216# OR2X1_LOC_95/Y 0.01fF
C20920 OR2X1_LOC_139/a_8_216# OR2X1_LOC_267/A 0.04fF
C20921 OR2X1_LOC_185/Y AND2X1_LOC_3/Y 0.09fF
C20922 OR2X1_LOC_585/A OR2X1_LOC_753/A 0.45fF
C20923 OR2X1_LOC_6/B OR2X1_LOC_84/Y 0.17fF
C20924 AND2X1_LOC_342/a_36_24# OR2X1_LOC_26/Y 0.01fF
C20925 AND2X1_LOC_170/Y AND2X1_LOC_566/Y 0.83fF
C20926 OR2X1_LOC_186/Y OR2X1_LOC_854/A 0.39fF
C20927 OR2X1_LOC_123/a_36_216# OR2X1_LOC_786/Y 0.00fF
C20928 OR2X1_LOC_86/A AND2X1_LOC_243/Y 0.03fF
C20929 OR2X1_LOC_404/Y OR2X1_LOC_500/A 0.00fF
C20930 OR2X1_LOC_696/a_8_216# OR2X1_LOC_26/Y 0.03fF
C20931 OR2X1_LOC_680/A AND2X1_LOC_830/a_8_24# 0.01fF
C20932 OR2X1_LOC_107/a_8_216# OR2X1_LOC_47/Y 0.01fF
C20933 OR2X1_LOC_719/A OR2X1_LOC_553/A 0.21fF
C20934 AND2X1_LOC_64/Y OR2X1_LOC_714/A 0.02fF
C20935 AND2X1_LOC_91/B OR2X1_LOC_704/a_8_216# 0.01fF
C20936 OR2X1_LOC_786/A OR2X1_LOC_598/A 0.08fF
C20937 OR2X1_LOC_70/Y AND2X1_LOC_840/B 0.03fF
C20938 AND2X1_LOC_331/a_8_24# OR2X1_LOC_532/B 0.01fF
C20939 VDD AND2X1_LOC_462/B 0.02fF
C20940 AND2X1_LOC_847/a_8_24# OR2X1_LOC_44/Y 0.01fF
C20941 OR2X1_LOC_306/a_8_216# OR2X1_LOC_311/Y 0.01fF
C20942 OR2X1_LOC_299/a_8_216# OR2X1_LOC_7/A 0.02fF
C20943 OR2X1_LOC_291/A OR2X1_LOC_824/Y 0.02fF
C20944 AND2X1_LOC_7/B AND2X1_LOC_268/a_8_24# 0.02fF
C20945 OR2X1_LOC_26/Y AND2X1_LOC_276/Y 0.00fF
C20946 OR2X1_LOC_675/a_8_216# OR2X1_LOC_269/B 0.01fF
C20947 OR2X1_LOC_744/A OR2X1_LOC_184/Y 0.07fF
C20948 OR2X1_LOC_84/B AND2X1_LOC_79/Y 0.00fF
C20949 AND2X1_LOC_753/B AND2X1_LOC_56/a_8_24# 0.04fF
C20950 OR2X1_LOC_18/Y AND2X1_LOC_639/A 0.01fF
C20951 OR2X1_LOC_709/A OR2X1_LOC_789/A 0.22fF
C20952 OR2X1_LOC_542/a_8_216# OR2X1_LOC_552/A 0.01fF
C20953 AND2X1_LOC_633/Y AND2X1_LOC_573/A 0.00fF
C20954 D_INPUT_5 OR2X1_LOC_651/A 0.26fF
C20955 OR2X1_LOC_846/B OR2X1_LOC_269/B 0.02fF
C20956 OR2X1_LOC_474/Y OR2X1_LOC_506/B 0.03fF
C20957 VDD OR2X1_LOC_705/B 0.27fF
C20958 OR2X1_LOC_696/a_8_216# OR2X1_LOC_89/A 0.01fF
C20959 AND2X1_LOC_191/Y AND2X1_LOC_475/a_8_24# 0.05fF
C20960 OR2X1_LOC_348/a_8_216# OR2X1_LOC_348/B 0.06fF
C20961 OR2X1_LOC_471/Y OR2X1_LOC_739/A 0.03fF
C20962 OR2X1_LOC_329/Y OR2X1_LOC_331/Y 0.09fF
C20963 OR2X1_LOC_160/B OR2X1_LOC_675/Y 0.00fF
C20964 OR2X1_LOC_307/A OR2X1_LOC_779/B 0.35fF
C20965 OR2X1_LOC_530/a_8_216# OR2X1_LOC_437/A 0.05fF
C20966 D_INPUT_0 AND2X1_LOC_573/A 0.07fF
C20967 OR2X1_LOC_596/A OR2X1_LOC_513/Y 0.02fF
C20968 OR2X1_LOC_43/A AND2X1_LOC_307/Y 0.03fF
C20969 OR2X1_LOC_70/Y AND2X1_LOC_475/a_8_24# 0.17fF
C20970 OR2X1_LOC_62/A AND2X1_LOC_852/B 0.03fF
C20971 OR2X1_LOC_624/A AND2X1_LOC_47/Y 0.17fF
C20972 AND2X1_LOC_334/a_8_24# AND2X1_LOC_852/Y 0.03fF
C20973 AND2X1_LOC_22/Y OR2X1_LOC_195/a_8_216# 0.01fF
C20974 OR2X1_LOC_271/B INPUT_1 0.05fF
C20975 OR2X1_LOC_701/Y AND2X1_LOC_866/A 0.01fF
C20976 OR2X1_LOC_744/A OR2X1_LOC_70/A 0.28fF
C20977 AND2X1_LOC_572/A OR2X1_LOC_256/A 0.06fF
C20978 AND2X1_LOC_733/Y AND2X1_LOC_784/a_36_24# 0.00fF
C20979 OR2X1_LOC_428/A AND2X1_LOC_789/Y 0.04fF
C20980 OR2X1_LOC_64/Y AND2X1_LOC_651/B 0.04fF
C20981 OR2X1_LOC_476/Y OR2X1_LOC_479/a_8_216# 0.39fF
C20982 OR2X1_LOC_529/a_8_216# OR2X1_LOC_47/Y 0.01fF
C20983 OR2X1_LOC_32/Y INPUT_1 0.01fF
C20984 OR2X1_LOC_134/a_8_216# OR2X1_LOC_134/Y 0.01fF
C20985 OR2X1_LOC_574/A OR2X1_LOC_814/A 0.10fF
C20986 OR2X1_LOC_433/a_8_216# OR2X1_LOC_31/Y 0.19fF
C20987 OR2X1_LOC_36/Y OR2X1_LOC_607/Y 0.01fF
C20988 OR2X1_LOC_223/B OR2X1_LOC_223/A 0.17fF
C20989 AND2X1_LOC_866/A OR2X1_LOC_44/Y 0.39fF
C20990 AND2X1_LOC_726/Y AND2X1_LOC_726/a_8_24# 0.00fF
C20991 OR2X1_LOC_862/B OR2X1_LOC_558/a_8_216# 0.02fF
C20992 AND2X1_LOC_12/Y OR2X1_LOC_771/a_8_216# 0.01fF
C20993 OR2X1_LOC_136/a_36_216# OR2X1_LOC_136/Y 0.00fF
C20994 OR2X1_LOC_624/A OR2X1_LOC_598/A 0.10fF
C20995 OR2X1_LOC_3/Y OR2X1_LOC_256/A 0.03fF
C20996 AND2X1_LOC_139/A OR2X1_LOC_7/A 0.19fF
C20997 AND2X1_LOC_663/B INPUT_1 3.05fF
C20998 OR2X1_LOC_437/Y AND2X1_LOC_840/B 0.44fF
C20999 AND2X1_LOC_465/a_36_24# OR2X1_LOC_31/Y 0.00fF
C21000 OR2X1_LOC_70/Y OR2X1_LOC_31/Y 0.28fF
C21001 OR2X1_LOC_185/Y OR2X1_LOC_194/a_8_216# 0.04fF
C21002 OR2X1_LOC_154/A AND2X1_LOC_679/a_8_24# 0.01fF
C21003 OR2X1_LOC_48/B OR2X1_LOC_172/Y 0.44fF
C21004 OR2X1_LOC_160/A OR2X1_LOC_641/B 0.03fF
C21005 OR2X1_LOC_553/A OR2X1_LOC_675/Y 0.01fF
C21006 OR2X1_LOC_18/Y OR2X1_LOC_88/Y 0.00fF
C21007 OR2X1_LOC_136/Y OR2X1_LOC_135/Y 0.00fF
C21008 OR2X1_LOC_97/A OR2X1_LOC_61/A 0.01fF
C21009 OR2X1_LOC_18/Y OR2X1_LOC_172/Y 0.07fF
C21010 AND2X1_LOC_390/B OR2X1_LOC_47/Y 0.07fF
C21011 OR2X1_LOC_26/Y AND2X1_LOC_405/a_8_24# 0.01fF
C21012 OR2X1_LOC_820/A AND2X1_LOC_750/a_8_24# -0.02fF
C21013 OR2X1_LOC_696/A AND2X1_LOC_325/a_8_24# 0.03fF
C21014 OR2X1_LOC_66/A AND2X1_LOC_235/a_8_24# 0.01fF
C21015 AND2X1_LOC_47/Y OR2X1_LOC_54/Y 0.05fF
C21016 OR2X1_LOC_3/Y AND2X1_LOC_624/B 0.03fF
C21017 OR2X1_LOC_696/A AND2X1_LOC_352/B 0.03fF
C21018 OR2X1_LOC_518/Y AND2X1_LOC_326/B -0.00fF
C21019 OR2X1_LOC_3/Y OR2X1_LOC_67/Y 0.07fF
C21020 OR2X1_LOC_36/Y AND2X1_LOC_562/Y 0.52fF
C21021 OR2X1_LOC_89/A AND2X1_LOC_405/a_8_24# 0.12fF
C21022 AND2X1_LOC_632/a_36_24# AND2X1_LOC_620/Y 0.00fF
C21023 AND2X1_LOC_3/a_8_24# INPUT_6 0.01fF
C21024 OR2X1_LOC_476/a_36_216# OR2X1_LOC_223/A -0.00fF
C21025 OR2X1_LOC_205/Y OR2X1_LOC_215/A 0.31fF
C21026 OR2X1_LOC_376/A OR2X1_LOC_376/a_8_216# 0.47fF
C21027 OR2X1_LOC_269/B OR2X1_LOC_750/Y 0.29fF
C21028 OR2X1_LOC_151/A OR2X1_LOC_342/A 0.01fF
C21029 OR2X1_LOC_805/A AND2X1_LOC_268/a_8_24# 0.04fF
C21030 OR2X1_LOC_659/Y D_GATE_662 0.74fF
C21031 AND2X1_LOC_181/Y OR2X1_LOC_323/Y 0.12fF
C21032 OR2X1_LOC_237/a_36_216# OR2X1_LOC_437/A 0.15fF
C21033 OR2X1_LOC_665/a_8_216# AND2X1_LOC_793/Y -0.06fF
C21034 AND2X1_LOC_717/B AND2X1_LOC_563/Y 0.00fF
C21035 OR2X1_LOC_696/A OR2X1_LOC_517/A 0.03fF
C21036 OR2X1_LOC_816/A AND2X1_LOC_285/Y 0.03fF
C21037 AND2X1_LOC_539/Y OR2X1_LOC_91/A 0.03fF
C21038 AND2X1_LOC_794/B AND2X1_LOC_477/Y 0.01fF
C21039 OR2X1_LOC_318/A OR2X1_LOC_776/Y 0.06fF
C21040 OR2X1_LOC_11/a_8_216# OR2X1_LOC_17/Y 0.01fF
C21041 AND2X1_LOC_42/a_8_24# OR2X1_LOC_80/A 0.09fF
C21042 OR2X1_LOC_634/A OR2X1_LOC_415/Y 0.00fF
C21043 OR2X1_LOC_426/B OR2X1_LOC_428/A 0.10fF
C21044 OR2X1_LOC_602/Y OR2X1_LOC_161/B 0.02fF
C21045 AND2X1_LOC_191/B AND2X1_LOC_244/A 0.03fF
C21046 OR2X1_LOC_805/A OR2X1_LOC_174/Y 0.03fF
C21047 OR2X1_LOC_79/a_8_216# OR2X1_LOC_59/Y 0.01fF
C21048 OR2X1_LOC_131/A OR2X1_LOC_131/a_8_216# 0.11fF
C21049 AND2X1_LOC_866/A AND2X1_LOC_866/a_8_24# -0.00fF
C21050 OR2X1_LOC_502/A OR2X1_LOC_502/Y 0.01fF
C21051 OR2X1_LOC_621/A OR2X1_LOC_621/B 0.62fF
C21052 OR2X1_LOC_54/Y OR2X1_LOC_598/A 0.19fF
C21053 OR2X1_LOC_184/Y OR2X1_LOC_31/Y 0.00fF
C21054 OR2X1_LOC_13/Y AND2X1_LOC_200/a_8_24# 0.01fF
C21055 OR2X1_LOC_426/B OR2X1_LOC_595/A 1.27fF
C21056 OR2X1_LOC_808/B OR2X1_LOC_722/B 0.02fF
C21057 OR2X1_LOC_185/Y OR2X1_LOC_576/a_8_216# 0.01fF
C21058 AND2X1_LOC_91/B OR2X1_LOC_105/Y 0.03fF
C21059 OR2X1_LOC_473/Y OR2X1_LOC_68/B 0.02fF
C21060 OR2X1_LOC_161/A OR2X1_LOC_500/a_36_216# 0.00fF
C21061 OR2X1_LOC_452/A OR2X1_LOC_450/Y 0.06fF
C21062 AND2X1_LOC_359/B OR2X1_LOC_248/A 0.04fF
C21063 AND2X1_LOC_18/Y OR2X1_LOC_362/A 0.07fF
C21064 VDD AND2X1_LOC_477/Y 0.03fF
C21065 OR2X1_LOC_604/A AND2X1_LOC_254/a_8_24# -0.04fF
C21066 AND2X1_LOC_306/a_8_24# OR2X1_LOC_161/B 0.01fF
C21067 OR2X1_LOC_64/Y AND2X1_LOC_793/B 0.35fF
C21068 AND2X1_LOC_70/Y AND2X1_LOC_275/a_8_24# 0.01fF
C21069 OR2X1_LOC_841/a_8_216# AND2X1_LOC_22/Y 0.01fF
C21070 OR2X1_LOC_604/A AND2X1_LOC_860/A 0.50fF
C21071 AND2X1_LOC_543/Y OR2X1_LOC_427/A 0.00fF
C21072 OR2X1_LOC_596/A OR2X1_LOC_702/a_36_216# 0.00fF
C21073 VDD OR2X1_LOC_777/a_8_216# 0.21fF
C21074 OR2X1_LOC_186/Y OR2X1_LOC_538/A 1.59fF
C21075 OR2X1_LOC_832/a_8_216# AND2X1_LOC_18/Y 0.01fF
C21076 AND2X1_LOC_529/a_36_24# OR2X1_LOC_548/B 0.00fF
C21077 OR2X1_LOC_604/A OR2X1_LOC_626/Y 0.03fF
C21078 AND2X1_LOC_40/Y OR2X1_LOC_139/A 0.03fF
C21079 D_INPUT_3 OR2X1_LOC_396/Y 0.14fF
C21080 OR2X1_LOC_671/a_8_216# VDD 0.00fF
C21081 OR2X1_LOC_523/B OR2X1_LOC_235/B 0.01fF
C21082 AND2X1_LOC_40/Y OR2X1_LOC_758/a_8_216# 0.04fF
C21083 AND2X1_LOC_22/Y OR2X1_LOC_856/B 0.20fF
C21084 OR2X1_LOC_129/a_8_216# OR2X1_LOC_59/Y 0.14fF
C21085 OR2X1_LOC_660/a_8_216# AND2X1_LOC_44/Y 0.01fF
C21086 OR2X1_LOC_308/a_36_216# AND2X1_LOC_44/Y 0.00fF
C21087 AND2X1_LOC_191/B OR2X1_LOC_108/Y 0.00fF
C21088 OR2X1_LOC_8/Y OR2X1_LOC_822/Y 0.01fF
C21089 AND2X1_LOC_98/a_8_24# OR2X1_LOC_51/Y 0.02fF
C21090 AND2X1_LOC_555/Y AND2X1_LOC_848/Y 0.03fF
C21091 OR2X1_LOC_31/Y OR2X1_LOC_70/A 0.05fF
C21092 OR2X1_LOC_160/A OR2X1_LOC_227/A 0.03fF
C21093 OR2X1_LOC_756/B OR2X1_LOC_151/A 0.29fF
C21094 OR2X1_LOC_535/A OR2X1_LOC_354/A 0.00fF
C21095 AND2X1_LOC_710/a_36_24# OR2X1_LOC_748/A 0.00fF
C21096 AND2X1_LOC_12/Y OR2X1_LOC_338/A 0.01fF
C21097 OR2X1_LOC_151/A OR2X1_LOC_735/a_36_216# 0.01fF
C21098 AND2X1_LOC_460/a_36_24# OR2X1_LOC_588/A 0.00fF
C21099 OR2X1_LOC_40/Y AND2X1_LOC_514/a_36_24# 0.00fF
C21100 AND2X1_LOC_21/Y INPUT_6 1.02fF
C21101 AND2X1_LOC_301/a_8_24# OR2X1_LOC_59/Y 0.14fF
C21102 AND2X1_LOC_729/a_8_24# OR2X1_LOC_92/Y 0.02fF
C21103 VDD OR2X1_LOC_329/B 0.42fF
C21104 AND2X1_LOC_354/Y AND2X1_LOC_802/Y 0.01fF
C21105 AND2X1_LOC_326/B OR2X1_LOC_91/A 0.03fF
C21106 OR2X1_LOC_132/a_8_216# OR2X1_LOC_132/Y 0.05fF
C21107 OR2X1_LOC_440/A AND2X1_LOC_31/Y 0.11fF
C21108 AND2X1_LOC_510/A AND2X1_LOC_508/a_36_24# 0.00fF
C21109 OR2X1_LOC_45/B AND2X1_LOC_454/Y 0.01fF
C21110 OR2X1_LOC_97/A AND2X1_LOC_601/a_8_24# 0.01fF
C21111 OR2X1_LOC_620/Y OR2X1_LOC_486/Y 0.03fF
C21112 OR2X1_LOC_188/Y OR2X1_LOC_465/a_8_216# 0.01fF
C21113 AND2X1_LOC_853/Y OR2X1_LOC_171/Y 0.04fF
C21114 OR2X1_LOC_436/a_8_216# OR2X1_LOC_174/Y 0.18fF
C21115 AND2X1_LOC_337/a_36_24# OR2X1_LOC_91/A 0.00fF
C21116 AND2X1_LOC_580/A GATE_579 0.05fF
C21117 OR2X1_LOC_589/A OR2X1_LOC_427/A 0.03fF
C21118 AND2X1_LOC_865/A AND2X1_LOC_861/a_36_24# 0.00fF
C21119 OR2X1_LOC_160/B OR2X1_LOC_808/B 0.01fF
C21120 OR2X1_LOC_78/A OR2X1_LOC_78/B 1.11fF
C21121 OR2X1_LOC_474/Y AND2X1_LOC_18/Y 0.37fF
C21122 AND2X1_LOC_476/a_8_24# OR2X1_LOC_6/A 0.01fF
C21123 OR2X1_LOC_656/B AND2X1_LOC_65/A 0.53fF
C21124 OR2X1_LOC_84/Y OR2X1_LOC_598/A 0.00fF
C21125 OR2X1_LOC_186/Y AND2X1_LOC_12/Y 0.07fF
C21126 AND2X1_LOC_443/Y AND2X1_LOC_444/a_8_24# 0.03fF
C21127 AND2X1_LOC_795/Y OR2X1_LOC_406/A 0.22fF
C21128 OR2X1_LOC_427/A OR2X1_LOC_322/Y 0.01fF
C21129 OR2X1_LOC_122/Y OR2X1_LOC_56/A 0.01fF
C21130 AND2X1_LOC_810/A OR2X1_LOC_306/Y 0.01fF
C21131 AND2X1_LOC_160/Y OR2X1_LOC_697/Y 0.01fF
C21132 OR2X1_LOC_600/A OR2X1_LOC_92/Y 0.03fF
C21133 AND2X1_LOC_442/a_8_24# AND2X1_LOC_36/Y 0.07fF
C21134 AND2X1_LOC_41/A AND2X1_LOC_92/Y 0.33fF
C21135 VDD OR2X1_LOC_502/A 1.23fF
C21136 OR2X1_LOC_604/A AND2X1_LOC_155/a_8_24# 0.01fF
C21137 AND2X1_LOC_303/A AND2X1_LOC_786/Y -0.03fF
C21138 AND2X1_LOC_367/a_8_24# OR2X1_LOC_428/A 0.17fF
C21139 OR2X1_LOC_603/a_8_216# OR2X1_LOC_12/Y 0.08fF
C21140 OR2X1_LOC_45/B OR2X1_LOC_599/A 0.03fF
C21141 AND2X1_LOC_229/a_8_24# OR2X1_LOC_87/A 0.04fF
C21142 OR2X1_LOC_715/B OR2X1_LOC_405/A 0.11fF
C21143 AND2X1_LOC_745/a_8_24# OR2X1_LOC_161/A 0.11fF
C21144 OR2X1_LOC_795/a_8_216# OR2X1_LOC_228/Y 0.01fF
C21145 VDD OR2X1_LOC_74/Y 0.12fF
C21146 AND2X1_LOC_554/B AND2X1_LOC_772/Y 0.01fF
C21147 OR2X1_LOC_736/Y OR2X1_LOC_553/A 0.07fF
C21148 OR2X1_LOC_186/Y OR2X1_LOC_802/A 0.01fF
C21149 OR2X1_LOC_179/Y OR2X1_LOC_56/A 0.02fF
C21150 AND2X1_LOC_710/Y OR2X1_LOC_297/a_8_216# 0.49fF
C21151 OR2X1_LOC_131/A AND2X1_LOC_573/A 0.02fF
C21152 OR2X1_LOC_203/a_8_216# OR2X1_LOC_719/B 0.14fF
C21153 OR2X1_LOC_270/Y OR2X1_LOC_578/B 0.03fF
C21154 OR2X1_LOC_748/A OR2X1_LOC_759/a_8_216# 0.00fF
C21155 OR2X1_LOC_8/Y AND2X1_LOC_852/B 0.48fF
C21156 OR2X1_LOC_337/A OR2X1_LOC_468/Y 0.01fF
C21157 OR2X1_LOC_859/A OR2X1_LOC_579/A 0.07fF
C21158 OR2X1_LOC_45/B AND2X1_LOC_267/a_36_24# 0.01fF
C21159 AND2X1_LOC_850/a_8_24# AND2X1_LOC_860/A 0.01fF
C21160 OR2X1_LOC_668/a_8_216# OR2X1_LOC_66/A 0.10fF
C21161 AND2X1_LOC_300/a_36_24# AND2X1_LOC_43/B 0.01fF
C21162 OR2X1_LOC_78/A OR2X1_LOC_721/Y 0.14fF
C21163 OR2X1_LOC_6/B OR2X1_LOC_161/A 0.04fF
C21164 OR2X1_LOC_421/A OR2X1_LOC_433/Y 0.04fF
C21165 OR2X1_LOC_600/A OR2X1_LOC_257/a_8_216# 0.01fF
C21166 AND2X1_LOC_125/a_36_24# OR2X1_LOC_244/Y 0.00fF
C21167 OR2X1_LOC_68/B OR2X1_LOC_241/B 0.07fF
C21168 OR2X1_LOC_763/Y OR2X1_LOC_764/a_36_216# 0.00fF
C21169 OR2X1_LOC_204/Y OR2X1_LOC_549/A 0.02fF
C21170 OR2X1_LOC_12/Y OR2X1_LOC_588/Y 0.12fF
C21171 OR2X1_LOC_512/a_8_216# OR2X1_LOC_779/B 0.01fF
C21172 OR2X1_LOC_448/a_8_216# OR2X1_LOC_78/A 0.03fF
C21173 VDD OR2X1_LOC_571/B 0.20fF
C21174 OR2X1_LOC_252/a_8_216# OR2X1_LOC_626/Y 0.39fF
C21175 AND2X1_LOC_42/B AND2X1_LOC_7/B 0.06fF
C21176 OR2X1_LOC_49/A OR2X1_LOC_287/B 0.03fF
C21177 AND2X1_LOC_40/Y OR2X1_LOC_637/Y 0.09fF
C21178 OR2X1_LOC_8/Y OR2X1_LOC_18/Y 0.04fF
C21179 OR2X1_LOC_509/a_36_216# AND2X1_LOC_81/B 0.00fF
C21180 OR2X1_LOC_770/B OR2X1_LOC_287/B -0.00fF
C21181 OR2X1_LOC_176/Y OR2X1_LOC_74/A 0.05fF
C21182 VDD AND2X1_LOC_33/Y 0.21fF
C21183 AND2X1_LOC_784/A AND2X1_LOC_181/Y 0.05fF
C21184 OR2X1_LOC_743/A OR2X1_LOC_428/A 0.11fF
C21185 VDD AND2X1_LOC_113/Y 0.33fF
C21186 OR2X1_LOC_485/A AND2X1_LOC_786/Y 0.07fF
C21187 AND2X1_LOC_191/Y AND2X1_LOC_213/B 0.04fF
C21188 OR2X1_LOC_158/A AND2X1_LOC_264/a_8_24# 0.01fF
C21189 AND2X1_LOC_19/Y OR2X1_LOC_655/a_8_216# 0.04fF
C21190 OR2X1_LOC_427/A OR2X1_LOC_297/A 0.01fF
C21191 AND2X1_LOC_7/B OR2X1_LOC_705/Y 0.03fF
C21192 OR2X1_LOC_708/Y OR2X1_LOC_712/a_8_216# 0.39fF
C21193 OR2X1_LOC_756/B OR2X1_LOC_788/a_8_216# 0.01fF
C21194 AND2X1_LOC_12/Y AND2X1_LOC_310/a_8_24# 0.01fF
C21195 OR2X1_LOC_40/Y OR2X1_LOC_44/Y 0.10fF
C21196 OR2X1_LOC_703/B OR2X1_LOC_66/A 0.29fF
C21197 OR2X1_LOC_822/a_8_216# OR2X1_LOC_6/A 0.14fF
C21198 VDD OR2X1_LOC_213/A 0.08fF
C21199 AND2X1_LOC_707/Y OR2X1_LOC_681/Y 0.05fF
C21200 OR2X1_LOC_216/A OR2X1_LOC_475/a_8_216# 0.03fF
C21201 OR2X1_LOC_319/B OR2X1_LOC_854/a_8_216# 0.06fF
C21202 OR2X1_LOC_51/Y AND2X1_LOC_848/Y 0.03fF
C21203 OR2X1_LOC_662/A AND2X1_LOC_92/Y 0.06fF
C21204 OR2X1_LOC_276/A AND2X1_LOC_36/Y 0.16fF
C21205 OR2X1_LOC_6/B OR2X1_LOC_26/Y 0.03fF
C21206 OR2X1_LOC_74/A AND2X1_LOC_212/Y 0.07fF
C21207 OR2X1_LOC_49/A OR2X1_LOC_97/a_8_216# 0.01fF
C21208 OR2X1_LOC_329/B OR2X1_LOC_315/Y 0.00fF
C21209 OR2X1_LOC_87/A OR2X1_LOC_66/A 0.11fF
C21210 OR2X1_LOC_448/B OR2X1_LOC_448/a_8_216# 0.07fF
C21211 OR2X1_LOC_375/A OR2X1_LOC_78/A 1.89fF
C21212 AND2X1_LOC_472/B OR2X1_LOC_461/B 0.05fF
C21213 OR2X1_LOC_744/A AND2X1_LOC_124/a_8_24# 0.02fF
C21214 AND2X1_LOC_544/a_8_24# OR2X1_LOC_427/A 0.01fF
C21215 AND2X1_LOC_696/a_8_24# OR2X1_LOC_66/A 0.03fF
C21216 OR2X1_LOC_185/A AND2X1_LOC_126/a_8_24# 0.03fF
C21217 VDD OR2X1_LOC_137/Y 0.06fF
C21218 AND2X1_LOC_713/Y OR2X1_LOC_89/A 0.01fF
C21219 OR2X1_LOC_283/Y OR2X1_LOC_51/Y 0.54fF
C21220 AND2X1_LOC_757/a_8_24# OR2X1_LOC_555/B 0.41fF
C21221 AND2X1_LOC_302/a_36_24# OR2X1_LOC_56/A 0.00fF
C21222 OR2X1_LOC_125/Y OR2X1_LOC_428/A 0.04fF
C21223 OR2X1_LOC_495/Y OR2X1_LOC_427/A 0.03fF
C21224 OR2X1_LOC_642/a_36_216# AND2X1_LOC_92/Y 0.00fF
C21225 OR2X1_LOC_458/B OR2X1_LOC_375/A 0.03fF
C21226 OR2X1_LOC_185/Y INPUT_0 0.07fF
C21227 OR2X1_LOC_92/Y OR2X1_LOC_619/Y 0.14fF
C21228 AND2X1_LOC_56/B OR2X1_LOC_410/a_8_216# 0.02fF
C21229 AND2X1_LOC_12/Y OR2X1_LOC_862/A 0.17fF
C21230 AND2X1_LOC_387/B AND2X1_LOC_387/a_8_24# 0.04fF
C21231 OR2X1_LOC_858/A OR2X1_LOC_778/Y 0.03fF
C21232 OR2X1_LOC_842/A AND2X1_LOC_3/Y 0.06fF
C21233 OR2X1_LOC_427/A AND2X1_LOC_450/a_8_24# 0.02fF
C21234 OR2X1_LOC_324/a_36_216# OR2X1_LOC_739/A 0.00fF
C21235 AND2X1_LOC_520/Y AND2X1_LOC_642/a_8_24# 0.01fF
C21236 AND2X1_LOC_99/A OR2X1_LOC_278/Y 0.00fF
C21237 OR2X1_LOC_466/A OR2X1_LOC_453/Y 0.15fF
C21238 OR2X1_LOC_246/A OR2X1_LOC_595/A 0.31fF
C21239 OR2X1_LOC_225/a_8_216# OR2X1_LOC_428/A 0.01fF
C21240 OR2X1_LOC_448/B OR2X1_LOC_375/A 0.01fF
C21241 AND2X1_LOC_489/Y AND2X1_LOC_558/a_8_24# 0.22fF
C21242 AND2X1_LOC_76/Y OR2X1_LOC_18/Y 0.07fF
C21243 OR2X1_LOC_155/A OR2X1_LOC_78/B 0.19fF
C21244 OR2X1_LOC_6/B AND2X1_LOC_51/Y 0.21fF
C21245 AND2X1_LOC_22/Y AND2X1_LOC_431/a_36_24# 0.00fF
C21246 OR2X1_LOC_523/Y OR2X1_LOC_161/A 0.01fF
C21247 OR2X1_LOC_602/B OR2X1_LOC_161/B 0.02fF
C21248 OR2X1_LOC_574/A OR2X1_LOC_715/A 0.01fF
C21249 OR2X1_LOC_22/Y OR2X1_LOC_829/A 0.17fF
C21250 AND2X1_LOC_22/a_8_24# AND2X1_LOC_47/a_8_24# 0.23fF
C21251 OR2X1_LOC_364/A OR2X1_LOC_775/a_8_216# 0.01fF
C21252 AND2X1_LOC_848/A AND2X1_LOC_793/a_8_24# 0.06fF
C21253 OR2X1_LOC_399/A AND2X1_LOC_573/A 0.01fF
C21254 OR2X1_LOC_158/A OR2X1_LOC_46/A 0.25fF
C21255 OR2X1_LOC_51/Y OR2X1_LOC_617/Y 0.00fF
C21256 OR2X1_LOC_405/A OR2X1_LOC_215/Y 0.10fF
C21257 OR2X1_LOC_185/Y OR2X1_LOC_860/Y 0.01fF
C21258 OR2X1_LOC_45/B AND2X1_LOC_866/A 0.03fF
C21259 OR2X1_LOC_409/B OR2X1_LOC_428/A 0.03fF
C21260 OR2X1_LOC_160/A OR2X1_LOC_739/A 0.00fF
C21261 AND2X1_LOC_549/a_8_24# OR2X1_LOC_74/A 0.04fF
C21262 OR2X1_LOC_36/Y OR2X1_LOC_23/a_8_216# -0.00fF
C21263 OR2X1_LOC_115/a_8_216# OR2X1_LOC_510/Y 0.01fF
C21264 AND2X1_LOC_316/a_8_24# OR2X1_LOC_810/A 0.05fF
C21265 OR2X1_LOC_261/a_36_216# AND2X1_LOC_663/B 0.01fF
C21266 AND2X1_LOC_160/Y OR2X1_LOC_696/Y 0.15fF
C21267 OR2X1_LOC_557/A OR2X1_LOC_78/Y 0.03fF
C21268 AND2X1_LOC_12/Y OR2X1_LOC_773/B 0.00fF
C21269 AND2X1_LOC_506/a_8_24# OR2X1_LOC_74/A 0.04fF
C21270 OR2X1_LOC_441/Y OR2X1_LOC_89/A 0.03fF
C21271 OR2X1_LOC_100/a_8_216# AND2X1_LOC_81/B 0.02fF
C21272 OR2X1_LOC_411/a_8_216# OR2X1_LOC_16/A 0.06fF
C21273 OR2X1_LOC_80/Y AND2X1_LOC_400/a_8_24# 0.23fF
C21274 OR2X1_LOC_667/Y OR2X1_LOC_26/Y 0.01fF
C21275 OR2X1_LOC_64/Y AND2X1_LOC_468/a_8_24# 0.05fF
C21276 AND2X1_LOC_47/Y OR2X1_LOC_346/A 0.01fF
C21277 OR2X1_LOC_43/A OR2X1_LOC_427/A 1.26fF
C21278 VDD AND2X1_LOC_48/A 0.42fF
C21279 OR2X1_LOC_164/Y OR2X1_LOC_371/Y 0.05fF
C21280 OR2X1_LOC_43/A AND2X1_LOC_801/a_8_24# -0.00fF
C21281 AND2X1_LOC_12/Y AND2X1_LOC_81/B 0.03fF
C21282 OR2X1_LOC_36/Y OR2X1_LOC_432/Y 0.02fF
C21283 OR2X1_LOC_88/A OR2X1_LOC_65/B 0.43fF
C21284 AND2X1_LOC_644/Y OR2X1_LOC_44/Y 0.00fF
C21285 OR2X1_LOC_446/B OR2X1_LOC_730/B 0.43fF
C21286 OR2X1_LOC_47/Y AND2X1_LOC_639/B 0.35fF
C21287 OR2X1_LOC_228/Y OR2X1_LOC_333/A 0.06fF
C21288 AND2X1_LOC_186/a_8_24# OR2X1_LOC_680/A 0.02fF
C21289 AND2X1_LOC_12/Y OR2X1_LOC_358/B 0.03fF
C21290 OR2X1_LOC_185/Y OR2X1_LOC_789/B 0.02fF
C21291 OR2X1_LOC_814/a_8_216# AND2X1_LOC_3/Y 0.02fF
C21292 AND2X1_LOC_47/Y OR2X1_LOC_565/A 0.03fF
C21293 OR2X1_LOC_158/A AND2X1_LOC_227/Y 0.03fF
C21294 AND2X1_LOC_392/A INPUT_1 0.07fF
C21295 AND2X1_LOC_729/Y AND2X1_LOC_192/Y 0.03fF
C21296 AND2X1_LOC_449/a_8_24# OR2X1_LOC_423/Y 0.23fF
C21297 OR2X1_LOC_424/Y AND2X1_LOC_592/a_8_24# 0.10fF
C21298 AND2X1_LOC_56/B OR2X1_LOC_203/a_8_216# 0.01fF
C21299 OR2X1_LOC_127/Y OR2X1_LOC_6/A 0.01fF
C21300 OR2X1_LOC_48/B OR2X1_LOC_52/B 0.20fF
C21301 OR2X1_LOC_802/Y OR2X1_LOC_539/Y 0.05fF
C21302 OR2X1_LOC_18/Y AND2X1_LOC_374/Y 0.02fF
C21303 OR2X1_LOC_377/A OR2X1_LOC_97/B 0.00fF
C21304 OR2X1_LOC_599/A AND2X1_LOC_435/a_8_24# 0.01fF
C21305 OR2X1_LOC_160/B AND2X1_LOC_692/a_36_24# 0.00fF
C21306 OR2X1_LOC_424/a_8_216# OR2X1_LOC_44/Y 0.05fF
C21307 AND2X1_LOC_155/a_36_24# OR2X1_LOC_7/A 0.01fF
C21308 OR2X1_LOC_479/Y OR2X1_LOC_469/Y 7.71fF
C21309 AND2X1_LOC_197/a_8_24# AND2X1_LOC_197/Y 0.01fF
C21310 OR2X1_LOC_667/Y OR2X1_LOC_89/A 0.02fF
C21311 OR2X1_LOC_468/Y OR2X1_LOC_539/Y 0.01fF
C21312 OR2X1_LOC_733/B OR2X1_LOC_737/A 0.12fF
C21313 AND2X1_LOC_535/Y AND2X1_LOC_169/a_8_24# 0.01fF
C21314 AND2X1_LOC_578/A AND2X1_LOC_168/a_8_24# 0.10fF
C21315 OR2X1_LOC_18/Y OR2X1_LOC_52/B 0.38fF
C21316 OR2X1_LOC_160/A OR2X1_LOC_269/B 0.14fF
C21317 AND2X1_LOC_41/A AND2X1_LOC_666/a_36_24# 0.01fF
C21318 OR2X1_LOC_547/B AND2X1_LOC_528/a_8_24# 0.04fF
C21319 OR2X1_LOC_413/a_36_216# OR2X1_LOC_52/B 0.02fF
C21320 OR2X1_LOC_91/A AND2X1_LOC_687/A 0.03fF
C21321 OR2X1_LOC_97/B AND2X1_LOC_824/B 0.04fF
C21322 OR2X1_LOC_472/B INPUT_0 0.24fF
C21323 AND2X1_LOC_483/Y OR2X1_LOC_816/A 0.11fF
C21324 OR2X1_LOC_517/A AND2X1_LOC_663/B 1.99fF
C21325 OR2X1_LOC_450/A OR2X1_LOC_446/Y 0.01fF
C21326 OR2X1_LOC_470/a_8_216# OR2X1_LOC_470/A 0.39fF
C21327 AND2X1_LOC_578/A AND2X1_LOC_851/A 0.06fF
C21328 OR2X1_LOC_76/A OR2X1_LOC_808/A 0.08fF
C21329 OR2X1_LOC_26/Y AND2X1_LOC_287/a_36_24# 0.00fF
C21330 OR2X1_LOC_169/B OR2X1_LOC_778/Y 0.05fF
C21331 AND2X1_LOC_139/B OR2X1_LOC_26/Y 0.00fF
C21332 AND2X1_LOC_59/Y OR2X1_LOC_84/B 0.28fF
C21333 AND2X1_LOC_729/Y OR2X1_LOC_585/A 0.59fF
C21334 AND2X1_LOC_537/Y AND2X1_LOC_303/a_8_24# 0.17fF
C21335 AND2X1_LOC_772/B OR2X1_LOC_71/Y 0.00fF
C21336 OR2X1_LOC_375/A OR2X1_LOC_155/A 0.04fF
C21337 OR2X1_LOC_235/B OR2X1_LOC_62/B 0.45fF
C21338 AND2X1_LOC_715/a_8_24# AND2X1_LOC_354/B 0.01fF
C21339 AND2X1_LOC_674/a_8_24# OR2X1_LOC_737/A 0.04fF
C21340 AND2X1_LOC_836/a_8_24# OR2X1_LOC_6/A 0.17fF
C21341 AND2X1_LOC_811/a_36_24# OR2X1_LOC_52/B 0.00fF
C21342 AND2X1_LOC_72/B OR2X1_LOC_294/Y 1.19fF
C21343 OR2X1_LOC_121/Y OR2X1_LOC_66/Y 0.01fF
C21344 OR2X1_LOC_392/B OR2X1_LOC_228/Y 0.07fF
C21345 AND2X1_LOC_214/A AND2X1_LOC_196/Y 0.18fF
C21346 OR2X1_LOC_54/Y AND2X1_LOC_240/a_36_24# 0.00fF
C21347 VDD OR2X1_LOC_618/Y 0.00fF
C21348 AND2X1_LOC_51/Y OR2X1_LOC_523/Y 0.03fF
C21349 AND2X1_LOC_604/a_36_24# OR2X1_LOC_318/B 0.00fF
C21350 OR2X1_LOC_89/A OR2X1_LOC_767/a_36_216# 0.00fF
C21351 VDD GATE_662 0.07fF
C21352 OR2X1_LOC_864/A OR2X1_LOC_849/A 0.03fF
C21353 OR2X1_LOC_61/B OR2X1_LOC_750/A 0.13fF
C21354 AND2X1_LOC_42/B OR2X1_LOC_805/A 0.02fF
C21355 OR2X1_LOC_74/A OR2X1_LOC_265/Y 0.07fF
C21356 OR2X1_LOC_516/B AND2X1_LOC_477/A 0.10fF
C21357 OR2X1_LOC_489/a_8_216# OR2X1_LOC_773/a_8_216# 0.47fF
C21358 OR2X1_LOC_7/A OR2X1_LOC_44/Y 9.23fF
C21359 OR2X1_LOC_820/A OR2X1_LOC_751/A 0.82fF
C21360 OR2X1_LOC_494/A OR2X1_LOC_384/a_8_216# 0.48fF
C21361 OR2X1_LOC_861/a_8_216# OR2X1_LOC_846/A 0.00fF
C21362 OR2X1_LOC_770/A OR2X1_LOC_80/A 0.01fF
C21363 OR2X1_LOC_844/Y OR2X1_LOC_560/a_36_216# 0.00fF
C21364 AND2X1_LOC_738/a_8_24# GATE_811 0.00fF
C21365 OR2X1_LOC_639/B OR2X1_LOC_636/a_8_216# 0.06fF
C21366 AND2X1_LOC_649/Y AND2X1_LOC_219/Y 0.00fF
C21367 OR2X1_LOC_160/A OR2X1_LOC_215/A 0.03fF
C21368 OR2X1_LOC_680/A OR2X1_LOC_617/Y 0.03fF
C21369 AND2X1_LOC_91/B OR2X1_LOC_71/A 0.02fF
C21370 AND2X1_LOC_99/A OR2X1_LOC_19/B 0.03fF
C21371 AND2X1_LOC_663/B AND2X1_LOC_624/A 0.00fF
C21372 OR2X1_LOC_529/Y OR2X1_LOC_26/Y 0.04fF
C21373 AND2X1_LOC_340/Y OR2X1_LOC_88/Y 0.84fF
C21374 OR2X1_LOC_385/Y OR2X1_LOC_52/B 0.72fF
C21375 OR2X1_LOC_160/B AND2X1_LOC_289/a_8_24# 0.04fF
C21376 OR2X1_LOC_609/A AND2X1_LOC_610/a_36_24# 0.00fF
C21377 OR2X1_LOC_3/Y OR2X1_LOC_248/Y 0.02fF
C21378 AND2X1_LOC_56/B AND2X1_LOC_136/a_8_24# 0.02fF
C21379 OR2X1_LOC_865/B OR2X1_LOC_859/A 0.20fF
C21380 OR2X1_LOC_744/A OR2X1_LOC_47/Y 0.29fF
C21381 OR2X1_LOC_529/Y AND2X1_LOC_493/a_8_24# 0.01fF
C21382 AND2X1_LOC_348/A OR2X1_LOC_417/A 0.01fF
C21383 AND2X1_LOC_51/Y OR2X1_LOC_579/B 0.16fF
C21384 OR2X1_LOC_103/Y AND2X1_LOC_227/Y 0.02fF
C21385 AND2X1_LOC_12/Y OR2X1_LOC_196/B 0.43fF
C21386 OR2X1_LOC_654/A AND2X1_LOC_3/Y 0.03fF
C21387 OR2X1_LOC_251/a_8_216# D_INPUT_3 0.06fF
C21388 OR2X1_LOC_529/Y OR2X1_LOC_89/A 0.03fF
C21389 AND2X1_LOC_807/Y AND2X1_LOC_574/A 0.03fF
C21390 AND2X1_LOC_70/Y AND2X1_LOC_428/a_8_24# 0.01fF
C21391 OR2X1_LOC_32/B AND2X1_LOC_633/Y 0.02fF
C21392 AND2X1_LOC_578/A AND2X1_LOC_474/Y 0.07fF
C21393 AND2X1_LOC_12/Y AND2X1_LOC_692/a_8_24# 0.02fF
C21394 AND2X1_LOC_859/Y OR2X1_LOC_64/Y 0.02fF
C21395 OR2X1_LOC_160/A AND2X1_LOC_146/a_8_24# 0.00fF
C21396 OR2X1_LOC_837/B OR2X1_LOC_416/A 0.43fF
C21397 AND2X1_LOC_44/Y OR2X1_LOC_501/a_8_216# 0.01fF
C21398 AND2X1_LOC_59/Y OR2X1_LOC_520/A 0.01fF
C21399 AND2X1_LOC_578/A OR2X1_LOC_485/A 0.07fF
C21400 OR2X1_LOC_103/a_8_216# AND2X1_LOC_227/Y 0.01fF
C21401 D_INPUT_3 AND2X1_LOC_401/a_8_24# 0.17fF
C21402 OR2X1_LOC_604/A AND2X1_LOC_562/Y 0.22fF
C21403 OR2X1_LOC_296/Y AND2X1_LOC_42/B 0.03fF
C21404 OR2X1_LOC_605/A OR2X1_LOC_605/B 0.61fF
C21405 AND2X1_LOC_47/Y OR2X1_LOC_161/A 11.54fF
C21406 AND2X1_LOC_55/a_8_24# INPUT_1 0.03fF
C21407 AND2X1_LOC_98/Y OR2X1_LOC_813/Y 0.00fF
C21408 OR2X1_LOC_375/A OR2X1_LOC_228/a_8_216# 0.01fF
C21409 OR2X1_LOC_154/A AND2X1_LOC_15/a_8_24# 0.07fF
C21410 OR2X1_LOC_42/a_36_216# OR2X1_LOC_46/A 0.00fF
C21411 OR2X1_LOC_43/A AND2X1_LOC_687/B 1.51fF
C21412 OR2X1_LOC_127/a_36_216# D_INPUT_3 0.00fF
C21413 OR2X1_LOC_804/a_8_216# OR2X1_LOC_318/B 0.01fF
C21414 AND2X1_LOC_59/Y OR2X1_LOC_651/A 0.24fF
C21415 OR2X1_LOC_287/B OR2X1_LOC_401/a_36_216# 0.00fF
C21416 OR2X1_LOC_862/B OR2X1_LOC_68/B 0.20fF
C21417 OR2X1_LOC_91/Y OR2X1_LOC_95/Y 0.13fF
C21418 OR2X1_LOC_91/Y AND2X1_LOC_440/a_8_24# 0.03fF
C21419 AND2X1_LOC_25/Y AND2X1_LOC_47/Y 0.06fF
C21420 OR2X1_LOC_91/Y OR2X1_LOC_368/A 0.03fF
C21421 AND2X1_LOC_859/Y OR2X1_LOC_417/A 0.03fF
C21422 OR2X1_LOC_616/Y GATE_662 0.03fF
C21423 OR2X1_LOC_287/B OR2X1_LOC_287/a_8_216# 0.02fF
C21424 AND2X1_LOC_573/Y AND2X1_LOC_574/Y 0.01fF
C21425 OR2X1_LOC_796/B OR2X1_LOC_784/Y 0.21fF
C21426 OR2X1_LOC_164/Y AND2X1_LOC_222/Y 0.02fF
C21427 OR2X1_LOC_49/A OR2X1_LOC_395/Y 0.03fF
C21428 OR2X1_LOC_233/a_8_216# D_INPUT_0 0.08fF
C21429 OR2X1_LOC_481/A OR2X1_LOC_54/Y 0.07fF
C21430 AND2X1_LOC_839/A AND2X1_LOC_240/Y 0.83fF
C21431 AND2X1_LOC_76/Y AND2X1_LOC_215/A 0.37fF
C21432 D_INPUT_3 OR2X1_LOC_824/Y 0.01fF
C21433 AND2X1_LOC_64/Y OR2X1_LOC_563/A 0.60fF
C21434 AND2X1_LOC_715/A OR2X1_LOC_437/A 0.07fF
C21435 OR2X1_LOC_95/Y OR2X1_LOC_371/a_8_216# 0.03fF
C21436 OR2X1_LOC_47/Y AND2X1_LOC_840/B 0.05fF
C21437 OR2X1_LOC_637/A AND2X1_LOC_31/Y 0.06fF
C21438 OR2X1_LOC_696/A AND2X1_LOC_774/A 0.12fF
C21439 OR2X1_LOC_417/Y AND2X1_LOC_727/A 0.03fF
C21440 OR2X1_LOC_264/Y AND2X1_LOC_31/Y 0.26fF
C21441 AND2X1_LOC_12/Y OR2X1_LOC_66/Y 0.21fF
C21442 OR2X1_LOC_240/B OR2X1_LOC_598/A 0.03fF
C21443 OR2X1_LOC_18/Y AND2X1_LOC_216/A 0.27fF
C21444 OR2X1_LOC_62/A OR2X1_LOC_585/A 1.25fF
C21445 AND2X1_LOC_663/B AND2X1_LOC_621/a_8_24# 0.01fF
C21446 AND2X1_LOC_18/Y OR2X1_LOC_771/B 0.06fF
C21447 OR2X1_LOC_68/Y AND2X1_LOC_51/Y 0.01fF
C21448 OR2X1_LOC_241/a_8_216# OR2X1_LOC_241/B 0.05fF
C21449 OR2X1_LOC_161/A OR2X1_LOC_598/A 0.02fF
C21450 AND2X1_LOC_141/B OR2X1_LOC_71/Y 0.01fF
C21451 OR2X1_LOC_687/a_36_216# AND2X1_LOC_425/Y 0.00fF
C21452 OR2X1_LOC_44/Y OR2X1_LOC_511/a_8_216# 0.05fF
C21453 AND2X1_LOC_658/A OR2X1_LOC_142/Y 0.03fF
C21454 AND2X1_LOC_371/a_8_24# OR2X1_LOC_776/A 0.05fF
C21455 AND2X1_LOC_543/Y OR2X1_LOC_322/a_8_216# 0.07fF
C21456 OR2X1_LOC_656/B OR2X1_LOC_559/a_36_216# 0.00fF
C21457 AND2X1_LOC_47/Y AND2X1_LOC_51/Y 0.19fF
C21458 OR2X1_LOC_527/Y OR2X1_LOC_95/Y 0.03fF
C21459 OR2X1_LOC_66/A OR2X1_LOC_844/B 0.02fF
C21460 OR2X1_LOC_234/a_36_216# OR2X1_LOC_585/A 0.00fF
C21461 OR2X1_LOC_151/A OR2X1_LOC_140/B 0.11fF
C21462 OR2X1_LOC_427/A OR2X1_LOC_384/a_8_216# 0.02fF
C21463 AND2X1_LOC_554/a_8_24# OR2X1_LOC_595/A 0.02fF
C21464 OR2X1_LOC_417/Y OR2X1_LOC_95/Y 0.03fF
C21465 AND2X1_LOC_17/Y AND2X1_LOC_428/a_8_24# 0.01fF
C21466 OR2X1_LOC_105/Y OR2X1_LOC_579/a_36_216# 0.00fF
C21467 AND2X1_LOC_810/A OR2X1_LOC_176/Y 0.17fF
C21468 OR2X1_LOC_849/a_8_216# AND2X1_LOC_47/Y 0.01fF
C21469 OR2X1_LOC_52/B AND2X1_LOC_215/A -0.01fF
C21470 VDD OR2X1_LOC_525/a_8_216# 0.21fF
C21471 AND2X1_LOC_228/Y OR2X1_LOC_172/Y 0.00fF
C21472 OR2X1_LOC_97/A OR2X1_LOC_390/A 0.00fF
C21473 OR2X1_LOC_52/B AND2X1_LOC_228/a_36_24# 0.00fF
C21474 OR2X1_LOC_66/A OR2X1_LOC_390/B 0.01fF
C21475 OR2X1_LOC_812/B OR2X1_LOC_558/A 0.03fF
C21476 OR2X1_LOC_516/Y AND2X1_LOC_663/A 0.10fF
C21477 OR2X1_LOC_419/Y OR2X1_LOC_239/Y 0.49fF
C21478 OR2X1_LOC_685/a_36_216# AND2X1_LOC_430/B 0.00fF
C21479 OR2X1_LOC_841/A OR2X1_LOC_390/B 0.03fF
C21480 OR2X1_LOC_160/B OR2X1_LOC_120/a_8_216# 0.01fF
C21481 AND2X1_LOC_580/A AND2X1_LOC_657/A 0.07fF
C21482 OR2X1_LOC_755/A AND2X1_LOC_620/Y 0.03fF
C21483 OR2X1_LOC_601/a_8_216# OR2X1_LOC_95/Y 0.01fF
C21484 AND2X1_LOC_810/A AND2X1_LOC_212/Y 0.05fF
C21485 OR2X1_LOC_574/A OR2X1_LOC_318/B 0.03fF
C21486 AND2X1_LOC_95/Y OR2X1_LOC_366/Y 0.07fF
C21487 OR2X1_LOC_151/A OR2X1_LOC_355/A 0.09fF
C21488 OR2X1_LOC_643/A AND2X1_LOC_31/Y 0.03fF
C21489 AND2X1_LOC_547/Y AND2X1_LOC_564/B 0.02fF
C21490 OR2X1_LOC_528/Y AND2X1_LOC_734/a_8_24# 0.01fF
C21491 AND2X1_LOC_666/a_8_24# OR2X1_LOC_241/B 0.03fF
C21492 OR2X1_LOC_778/Y AND2X1_LOC_31/Y 0.09fF
C21493 OR2X1_LOC_22/Y OR2X1_LOC_224/Y 0.03fF
C21494 OR2X1_LOC_45/B OR2X1_LOC_40/Y 1.46fF
C21495 OR2X1_LOC_175/B OR2X1_LOC_175/a_8_216# 0.06fF
C21496 OR2X1_LOC_54/Y D_INPUT_1 0.34fF
C21497 OR2X1_LOC_710/B AND2X1_LOC_7/B 0.03fF
C21498 OR2X1_LOC_322/a_8_216# OR2X1_LOC_322/Y 0.01fF
C21499 OR2X1_LOC_461/Y OR2X1_LOC_598/A 0.01fF
C21500 OR2X1_LOC_7/A AND2X1_LOC_570/a_8_24# 0.01fF
C21501 OR2X1_LOC_485/A OR2X1_LOC_172/a_8_216# 0.01fF
C21502 AND2X1_LOC_51/Y OR2X1_LOC_598/A 2.38fF
C21503 OR2X1_LOC_739/A OR2X1_LOC_532/Y 0.03fF
C21504 OR2X1_LOC_375/A D_GATE_366 0.03fF
C21505 OR2X1_LOC_473/A OR2X1_LOC_532/B 0.72fF
C21506 OR2X1_LOC_620/Y OR2X1_LOC_308/Y 0.03fF
C21507 D_INPUT_3 OR2X1_LOC_95/Y 0.02fF
C21508 OR2X1_LOC_379/Y AND2X1_LOC_36/Y 0.04fF
C21509 AND2X1_LOC_742/a_8_24# AND2X1_LOC_731/Y 0.19fF
C21510 AND2X1_LOC_555/Y AND2X1_LOC_562/B 0.07fF
C21511 OR2X1_LOC_604/A OR2X1_LOC_381/a_8_216# 0.03fF
C21512 AND2X1_LOC_658/B AND2X1_LOC_213/B 0.03fF
C21513 OR2X1_LOC_837/Y OR2X1_LOC_20/A 0.18fF
C21514 AND2X1_LOC_348/Y OR2X1_LOC_437/A 0.16fF
C21515 OR2X1_LOC_719/B OR2X1_LOC_719/a_36_216# 0.03fF
C21516 AND2X1_LOC_530/a_8_24# VDD 0.00fF
C21517 OR2X1_LOC_106/Y AND2X1_LOC_116/a_36_24# 0.00fF
C21518 OR2X1_LOC_808/A OR2X1_LOC_722/B 0.10fF
C21519 OR2X1_LOC_421/A AND2X1_LOC_714/B 0.08fF
C21520 OR2X1_LOC_47/Y OR2X1_LOC_31/Y 3.32fF
C21521 OR2X1_LOC_753/A OR2X1_LOC_437/A 0.19fF
C21522 OR2X1_LOC_671/Y OR2X1_LOC_14/a_8_216# 0.01fF
C21523 AND2X1_LOC_56/B OR2X1_LOC_730/B 0.02fF
C21524 OR2X1_LOC_840/A OR2X1_LOC_831/B 0.08fF
C21525 OR2X1_LOC_696/A AND2X1_LOC_62/a_8_24# 0.01fF
C21526 OR2X1_LOC_160/B OR2X1_LOC_596/A 0.03fF
C21527 AND2X1_LOC_180/a_8_24# VDD -0.00fF
C21528 OR2X1_LOC_575/A OR2X1_LOC_115/B 0.03fF
C21529 OR2X1_LOC_155/A OR2X1_LOC_515/Y 0.04fF
C21530 OR2X1_LOC_235/B OR2X1_LOC_15/a_36_216# 0.00fF
C21531 OR2X1_LOC_154/A OR2X1_LOC_308/Y 0.07fF
C21532 OR2X1_LOC_269/B OR2X1_LOC_532/Y 0.02fF
C21533 VDD OR2X1_LOC_772/A 0.08fF
C21534 OR2X1_LOC_78/A OR2X1_LOC_549/A 1.50fF
C21535 OR2X1_LOC_161/A OR2X1_LOC_186/a_8_216# 0.01fF
C21536 AND2X1_LOC_47/Y OR2X1_LOC_551/B 0.60fF
C21537 OR2X1_LOC_389/A OR2X1_LOC_66/A 0.03fF
C21538 AND2X1_LOC_392/A AND2X1_LOC_352/B 0.05fF
C21539 OR2X1_LOC_340/Y AND2X1_LOC_226/a_8_24# 0.17fF
C21540 OR2X1_LOC_547/B AND2X1_LOC_7/B 0.03fF
C21541 AND2X1_LOC_266/a_8_24# AND2X1_LOC_249/a_8_24# 0.23fF
C21542 OR2X1_LOC_532/B OR2X1_LOC_228/Y 0.10fF
C21543 OR2X1_LOC_790/A AND2X1_LOC_41/A 0.02fF
C21544 OR2X1_LOC_448/A OR2X1_LOC_713/A 0.01fF
C21545 OR2X1_LOC_696/A OR2X1_LOC_752/a_8_216# 0.03fF
C21546 D_INPUT_0 OR2X1_LOC_68/B 0.33fF
C21547 OR2X1_LOC_130/A AND2X1_LOC_226/a_8_24# 0.03fF
C21548 OR2X1_LOC_542/B OR2X1_LOC_284/a_8_216# 0.47fF
C21549 OR2X1_LOC_541/B OR2X1_LOC_121/A 0.48fF
C21550 OR2X1_LOC_600/A AND2X1_LOC_296/a_8_24# 0.01fF
C21551 OR2X1_LOC_757/A OR2X1_LOC_815/a_8_216# 0.03fF
C21552 OR2X1_LOC_40/Y OR2X1_LOC_292/a_8_216# 0.03fF
C21553 OR2X1_LOC_427/A AND2X1_LOC_771/a_8_24# 0.06fF
C21554 AND2X1_LOC_774/a_8_24# OR2X1_LOC_48/B 0.01fF
C21555 OR2X1_LOC_600/A OR2X1_LOC_819/a_36_216# 0.00fF
C21556 AND2X1_LOC_340/Y AND2X1_LOC_76/Y 0.03fF
C21557 OR2X1_LOC_808/B OR2X1_LOC_180/a_8_216# 0.29fF
C21558 VDD OR2X1_LOC_632/a_8_216# 0.00fF
C21559 AND2X1_LOC_576/Y AND2X1_LOC_227/a_8_24# 0.01fF
C21560 OR2X1_LOC_49/A INPUT_3 0.41fF
C21561 OR2X1_LOC_648/A AND2X1_LOC_92/Y 0.07fF
C21562 AND2X1_LOC_765/a_8_24# AND2X1_LOC_12/Y 0.02fF
C21563 AND2X1_LOC_486/Y AND2X1_LOC_477/Y 0.13fF
C21564 AND2X1_LOC_392/A OR2X1_LOC_517/A 0.20fF
C21565 AND2X1_LOC_7/Y OR2X1_LOC_193/a_8_216# 0.07fF
C21566 AND2X1_LOC_181/Y AND2X1_LOC_76/Y 0.03fF
C21567 OR2X1_LOC_158/A OR2X1_LOC_689/a_36_216# 0.01fF
C21568 OR2X1_LOC_185/Y AND2X1_LOC_7/B 0.19fF
C21569 AND2X1_LOC_177/a_8_24# OR2X1_LOC_66/A 0.01fF
C21570 OR2X1_LOC_709/A OR2X1_LOC_447/a_8_216# 0.02fF
C21571 OR2X1_LOC_313/Y OR2X1_LOC_12/Y 0.51fF
C21572 AND2X1_LOC_160/a_8_24# OR2X1_LOC_51/Y 0.18fF
C21573 OR2X1_LOC_186/Y AND2X1_LOC_59/Y 0.77fF
C21574 AND2X1_LOC_12/Y OR2X1_LOC_833/Y 0.04fF
C21575 AND2X1_LOC_521/a_8_24# OR2X1_LOC_161/A 0.01fF
C21576 OR2X1_LOC_594/a_8_216# AND2X1_LOC_436/Y -0.00fF
C21577 AND2X1_LOC_477/Y AND2X1_LOC_811/B 0.00fF
C21578 AND2X1_LOC_564/B AND2X1_LOC_778/a_8_24# 0.02fF
C21579 AND2X1_LOC_287/B AND2X1_LOC_806/A 0.01fF
C21580 OR2X1_LOC_774/a_8_216# OR2X1_LOC_269/B 0.01fF
C21581 AND2X1_LOC_845/Y OR2X1_LOC_437/A 0.07fF
C21582 OR2X1_LOC_756/B OR2X1_LOC_287/A 0.26fF
C21583 AND2X1_LOC_317/a_8_24# OR2X1_LOC_16/A 0.04fF
C21584 OR2X1_LOC_196/Y OR2X1_LOC_269/B 0.01fF
C21585 OR2X1_LOC_54/Y AND2X1_LOC_789/Y 0.21fF
C21586 OR2X1_LOC_816/A AND2X1_LOC_806/A 0.03fF
C21587 OR2X1_LOC_149/a_36_216# OR2X1_LOC_161/A 0.00fF
C21588 OR2X1_LOC_179/a_8_216# OR2X1_LOC_59/Y 0.01fF
C21589 AND2X1_LOC_110/Y AND2X1_LOC_527/a_8_24# 0.08fF
C21590 OR2X1_LOC_438/Y OR2X1_LOC_56/A 0.07fF
C21591 AND2X1_LOC_737/a_36_24# AND2X1_LOC_658/A 0.01fF
C21592 OR2X1_LOC_158/A AND2X1_LOC_454/Y 0.01fF
C21593 OR2X1_LOC_287/B OR2X1_LOC_392/B 0.05fF
C21594 AND2X1_LOC_347/B AND2X1_LOC_847/Y 0.01fF
C21595 OR2X1_LOC_847/A INPUT_2 0.00fF
C21596 OR2X1_LOC_354/A OR2X1_LOC_78/A 0.03fF
C21597 OR2X1_LOC_6/A AND2X1_LOC_415/a_8_24# 0.01fF
C21598 AND2X1_LOC_57/a_36_24# OR2X1_LOC_66/A 0.00fF
C21599 OR2X1_LOC_585/A OR2X1_LOC_312/a_36_216# 0.00fF
C21600 OR2X1_LOC_814/A OR2X1_LOC_539/B 0.02fF
C21601 OR2X1_LOC_45/B AND2X1_LOC_857/a_8_24# 0.01fF
C21602 OR2X1_LOC_756/B OR2X1_LOC_174/A 0.26fF
C21603 OR2X1_LOC_18/Y AND2X1_LOC_244/a_8_24# 0.01fF
C21604 OR2X1_LOC_3/Y OR2X1_LOC_56/Y 0.01fF
C21605 OR2X1_LOC_66/a_8_216# OR2X1_LOC_560/A 0.01fF
C21606 OR2X1_LOC_455/a_8_216# OR2X1_LOC_161/B 0.06fF
C21607 OR2X1_LOC_485/A OR2X1_LOC_312/a_8_216# 0.02fF
C21608 OR2X1_LOC_45/B OR2X1_LOC_7/A 0.96fF
C21609 OR2X1_LOC_756/B OR2X1_LOC_435/a_8_216# 0.01fF
C21610 AND2X1_LOC_64/Y OR2X1_LOC_202/a_8_216# 0.01fF
C21611 OR2X1_LOC_107/Y OR2X1_LOC_103/Y 0.23fF
C21612 AND2X1_LOC_340/Y OR2X1_LOC_52/B 0.07fF
C21613 AND2X1_LOC_335/Y OR2X1_LOC_619/Y 0.02fF
C21614 AND2X1_LOC_276/Y AND2X1_LOC_473/Y 0.12fF
C21615 AND2X1_LOC_486/Y OR2X1_LOC_329/B 0.06fF
C21616 AND2X1_LOC_824/B OR2X1_LOC_410/Y 0.11fF
C21617 OR2X1_LOC_339/a_8_216# AND2X1_LOC_95/Y 0.01fF
C21618 OR2X1_LOC_346/B OR2X1_LOC_294/Y 0.01fF
C21619 OR2X1_LOC_599/A OR2X1_LOC_158/A 0.03fF
C21620 OR2X1_LOC_715/B OR2X1_LOC_653/A 0.03fF
C21621 OR2X1_LOC_24/Y AND2X1_LOC_219/A 0.21fF
C21622 AND2X1_LOC_468/B AND2X1_LOC_436/Y 0.01fF
C21623 OR2X1_LOC_329/B AND2X1_LOC_840/a_36_24# 0.01fF
C21624 D_INPUT_7 INPUT_7 0.85fF
C21625 OR2X1_LOC_87/A OR2X1_LOC_180/a_36_216# 0.00fF
C21626 AND2X1_LOC_131/a_36_24# OR2X1_LOC_510/Y 0.00fF
C21627 OR2X1_LOC_188/Y AND2X1_LOC_666/a_8_24# 0.01fF
C21628 OR2X1_LOC_573/Y OR2X1_LOC_66/A 0.01fF
C21629 AND2X1_LOC_738/B AND2X1_LOC_621/Y 0.07fF
C21630 AND2X1_LOC_638/Y AND2X1_LOC_651/a_8_24# 0.10fF
C21631 AND2X1_LOC_621/Y OR2X1_LOC_56/A 0.12fF
C21632 OR2X1_LOC_744/A OR2X1_LOC_625/Y 0.99fF
C21633 AND2X1_LOC_535/Y AND2X1_LOC_354/B 0.27fF
C21634 OR2X1_LOC_53/Y OR2X1_LOC_43/a_8_216# 0.01fF
C21635 VDD OR2X1_LOC_790/a_8_216# 0.21fF
C21636 OR2X1_LOC_102/a_8_216# OR2X1_LOC_7/A 0.01fF
C21637 VDD AND2X1_LOC_580/A 0.31fF
C21638 OR2X1_LOC_809/B OR2X1_LOC_539/Y 0.01fF
C21639 AND2X1_LOC_70/Y OR2X1_LOC_130/A 0.98fF
C21640 AND2X1_LOC_51/Y OR2X1_LOC_34/A 0.00fF
C21641 OR2X1_LOC_821/a_8_216# OR2X1_LOC_70/Y 0.07fF
C21642 AND2X1_LOC_338/Y AND2X1_LOC_333/a_8_24# 0.01fF
C21643 OR2X1_LOC_502/A AND2X1_LOC_328/a_8_24# 0.02fF
C21644 OR2X1_LOC_666/a_36_216# AND2X1_LOC_859/Y 0.01fF
C21645 OR2X1_LOC_158/A OR2X1_LOC_258/a_8_216# 0.20fF
C21646 OR2X1_LOC_644/B OR2X1_LOC_676/Y 0.76fF
C21647 OR2X1_LOC_805/A OR2X1_LOC_778/a_8_216# 0.03fF
C21648 AND2X1_LOC_510/a_8_24# AND2X1_LOC_573/A 0.01fF
C21649 OR2X1_LOC_599/A AND2X1_LOC_537/a_36_24# 0.00fF
C21650 AND2X1_LOC_3/Y AND2X1_LOC_265/a_8_24# 0.01fF
C21651 OR2X1_LOC_637/Y AND2X1_LOC_43/B 0.03fF
C21652 OR2X1_LOC_462/B OR2X1_LOC_520/a_8_216# 0.01fF
C21653 AND2X1_LOC_195/a_8_24# AND2X1_LOC_729/B 0.01fF
C21654 OR2X1_LOC_856/B AND2X1_LOC_173/a_8_24# -0.02fF
C21655 OR2X1_LOC_479/Y OR2X1_LOC_831/A 0.05fF
C21656 OR2X1_LOC_403/B OR2X1_LOC_66/A 0.01fF
C21657 OR2X1_LOC_97/A OR2X1_LOC_750/A 0.01fF
C21658 OR2X1_LOC_426/Y OR2X1_LOC_427/Y 0.05fF
C21659 OR2X1_LOC_8/Y OR2X1_LOC_585/A 0.21fF
C21660 OR2X1_LOC_185/A OR2X1_LOC_220/A 8.56fF
C21661 OR2X1_LOC_54/Y OR2X1_LOC_15/a_8_216# 0.04fF
C21662 AND2X1_LOC_95/Y OR2X1_LOC_802/a_36_216# 0.02fF
C21663 AND2X1_LOC_89/a_36_24# OR2X1_LOC_78/A 0.01fF
C21664 OR2X1_LOC_523/B OR2X1_LOC_404/Y 0.01fF
C21665 VDD AND2X1_LOC_3/Y 1.04fF
C21666 OR2X1_LOC_501/B OR2X1_LOC_203/Y 0.01fF
C21667 OR2X1_LOC_805/a_8_216# OR2X1_LOC_811/A 0.06fF
C21668 AND2X1_LOC_535/Y AND2X1_LOC_390/B 0.02fF
C21669 AND2X1_LOC_95/Y AND2X1_LOC_52/a_36_24# 0.01fF
C21670 OR2X1_LOC_293/a_8_216# OR2X1_LOC_16/A 0.43fF
C21671 VDD OR2X1_LOC_647/B 0.23fF
C21672 OR2X1_LOC_487/Y AND2X1_LOC_489/a_8_24# 0.23fF
C21673 OR2X1_LOC_160/B OR2X1_LOC_33/B 0.00fF
C21674 OR2X1_LOC_813/a_36_216# OR2X1_LOC_74/A 0.00fF
C21675 OR2X1_LOC_506/a_8_216# OR2X1_LOC_506/B 0.03fF
C21676 AND2X1_LOC_485/a_8_24# OR2X1_LOC_209/A 0.04fF
C21677 OR2X1_LOC_720/B AND2X1_LOC_44/Y -0.00fF
C21678 OR2X1_LOC_362/B OR2X1_LOC_811/A 0.12fF
C21679 OR2X1_LOC_589/A OR2X1_LOC_416/Y 0.02fF
C21680 OR2X1_LOC_256/Y OR2X1_LOC_85/A 0.05fF
C21681 OR2X1_LOC_656/B OR2X1_LOC_405/A 0.12fF
C21682 AND2X1_LOC_851/B AND2X1_LOC_465/A 0.03fF
C21683 OR2X1_LOC_401/Y OR2X1_LOC_78/A 0.16fF
C21684 OR2X1_LOC_379/Y AND2X1_LOC_586/a_8_24# 0.01fF
C21685 AND2X1_LOC_721/Y AND2X1_LOC_227/Y 0.02fF
C21686 OR2X1_LOC_389/B AND2X1_LOC_41/A 0.03fF
C21687 AND2X1_LOC_682/a_8_24# OR2X1_LOC_161/A 0.01fF
C21688 AND2X1_LOC_850/Y AND2X1_LOC_621/Y 0.05fF
C21689 AND2X1_LOC_95/Y OR2X1_LOC_624/A 1.02fF
C21690 AND2X1_LOC_803/B AND2X1_LOC_797/A 0.00fF
C21691 OR2X1_LOC_335/a_8_216# OR2X1_LOC_223/A 0.01fF
C21692 OR2X1_LOC_447/A OR2X1_LOC_739/A 0.01fF
C21693 OR2X1_LOC_849/a_36_216# OR2X1_LOC_113/B -0.00fF
C21694 OR2X1_LOC_286/B OR2X1_LOC_580/B 0.05fF
C21695 OR2X1_LOC_654/A INPUT_0 0.07fF
C21696 AND2X1_LOC_784/A AND2X1_LOC_857/Y 0.01fF
C21697 OR2X1_LOC_538/A OR2X1_LOC_574/A 0.03fF
C21698 OR2X1_LOC_506/A OR2X1_LOC_161/A 0.07fF
C21699 OR2X1_LOC_364/A OR2X1_LOC_318/Y 0.07fF
C21700 OR2X1_LOC_629/a_8_216# OR2X1_LOC_78/A 0.01fF
C21701 OR2X1_LOC_479/Y OR2X1_LOC_795/B 0.02fF
C21702 OR2X1_LOC_48/B OR2X1_LOC_48/a_8_216# 0.03fF
C21703 AND2X1_LOC_471/Y OR2X1_LOC_371/Y 0.13fF
C21704 OR2X1_LOC_264/Y OR2X1_LOC_864/A 0.03fF
C21705 AND2X1_LOC_721/a_8_24# OR2X1_LOC_26/Y 0.02fF
C21706 OR2X1_LOC_446/B AND2X1_LOC_419/a_36_24# -0.00fF
C21707 OR2X1_LOC_354/A OR2X1_LOC_155/A 0.02fF
C21708 OR2X1_LOC_757/A OR2X1_LOC_617/Y 0.03fF
C21709 AND2X1_LOC_779/a_8_24# OR2X1_LOC_36/Y 0.01fF
C21710 OR2X1_LOC_160/A OR2X1_LOC_539/Y 0.07fF
C21711 AND2X1_LOC_372/a_8_24# AND2X1_LOC_42/B 0.17fF
C21712 OR2X1_LOC_335/Y OR2X1_LOC_479/Y 0.04fF
C21713 AND2X1_LOC_512/Y OR2X1_LOC_743/A 0.00fF
C21714 OR2X1_LOC_92/Y AND2X1_LOC_454/A 0.09fF
C21715 OR2X1_LOC_18/Y AND2X1_LOC_286/Y 0.02fF
C21716 OR2X1_LOC_808/A OR2X1_LOC_794/a_8_216# 0.03fF
C21717 OR2X1_LOC_804/a_8_216# OR2X1_LOC_804/B 0.01fF
C21718 OR2X1_LOC_382/Y OR2X1_LOC_3/Y 0.03fF
C21719 OR2X1_LOC_812/B OR2X1_LOC_561/a_36_216# 0.00fF
C21720 OR2X1_LOC_164/Y OR2X1_LOC_74/A 0.02fF
C21721 OR2X1_LOC_799/A OR2X1_LOC_593/a_8_216# 0.01fF
C21722 AND2X1_LOC_59/Y AND2X1_LOC_81/B 0.46fF
C21723 OR2X1_LOC_47/Y AND2X1_LOC_464/A 0.42fF
C21724 AND2X1_LOC_580/A OR2X1_LOC_616/Y 1.25fF
C21725 AND2X1_LOC_663/B OR2X1_LOC_755/a_8_216# 0.01fF
C21726 OR2X1_LOC_47/Y AND2X1_LOC_213/B 0.14fF
C21727 OR2X1_LOC_300/a_8_216# OR2X1_LOC_300/Y 0.01fF
C21728 AND2X1_LOC_59/Y OR2X1_LOC_358/B 0.01fF
C21729 AND2X1_LOC_722/a_8_24# OR2X1_LOC_417/A 0.05fF
C21730 OR2X1_LOC_288/a_8_216# OR2X1_LOC_269/B 0.01fF
C21731 OR2X1_LOC_158/A AND2X1_LOC_866/A 0.08fF
C21732 OR2X1_LOC_185/Y OR2X1_LOC_805/A 0.08fF
C21733 AND2X1_LOC_95/Y OR2X1_LOC_552/a_8_216# 0.01fF
C21734 AND2X1_LOC_40/Y OR2X1_LOC_479/Y 0.10fF
C21735 OR2X1_LOC_797/A OR2X1_LOC_797/a_8_216# 0.39fF
C21736 AND2X1_LOC_339/Y OR2X1_LOC_289/Y 0.02fF
C21737 AND2X1_LOC_580/B OR2X1_LOC_616/a_36_216# 0.00fF
C21738 OR2X1_LOC_631/B OR2X1_LOC_499/a_36_216# 0.00fF
C21739 OR2X1_LOC_97/B OR2X1_LOC_375/A 1.60fF
C21740 AND2X1_LOC_807/Y AND2X1_LOC_806/A 0.03fF
C21741 AND2X1_LOC_852/Y OR2X1_LOC_69/A 0.05fF
C21742 AND2X1_LOC_732/B OR2X1_LOC_31/Y 0.00fF
C21743 OR2X1_LOC_786/Y AND2X1_LOC_65/A 0.04fF
C21744 AND2X1_LOC_554/B OR2X1_LOC_278/Y 0.02fF
C21745 INPUT_0 AND2X1_LOC_326/a_8_24# 0.02fF
C21746 OR2X1_LOC_40/Y AND2X1_LOC_811/Y 0.01fF
C21747 OR2X1_LOC_675/a_8_216# OR2X1_LOC_811/A 0.05fF
C21748 AND2X1_LOC_107/a_8_24# OR2X1_LOC_632/Y 0.02fF
C21749 OR2X1_LOC_208/A OR2X1_LOC_68/B 0.03fF
C21750 OR2X1_LOC_83/Y OR2X1_LOC_69/A 0.00fF
C21751 OR2X1_LOC_814/A OR2X1_LOC_78/B 0.33fF
C21752 OR2X1_LOC_585/A OR2X1_LOC_67/A 0.16fF
C21753 AND2X1_LOC_228/Y OR2X1_LOC_52/B 0.00fF
C21754 OR2X1_LOC_375/A OR2X1_LOC_710/a_36_216# 0.00fF
C21755 AND2X1_LOC_565/a_8_24# OR2X1_LOC_95/Y 0.01fF
C21756 OR2X1_LOC_280/Y OR2X1_LOC_18/Y 0.03fF
C21757 AND2X1_LOC_12/Y OR2X1_LOC_574/A 0.04fF
C21758 OR2X1_LOC_400/a_36_216# AND2X1_LOC_51/Y 0.00fF
C21759 OR2X1_LOC_303/a_8_216# OR2X1_LOC_353/a_8_216# 0.47fF
C21760 AND2X1_LOC_91/B AND2X1_LOC_31/Y 0.16fF
C21761 AND2X1_LOC_387/B OR2X1_LOC_377/A 0.02fF
C21762 OR2X1_LOC_834/A AND2X1_LOC_53/Y 0.39fF
C21763 AND2X1_LOC_12/Y OR2X1_LOC_33/A 0.01fF
C21764 AND2X1_LOC_7/B OR2X1_LOC_552/A 0.06fF
C21765 OR2X1_LOC_129/a_8_216# OR2X1_LOC_47/Y 0.02fF
C21766 AND2X1_LOC_64/Y OR2X1_LOC_724/A 0.13fF
C21767 OR2X1_LOC_154/A AND2X1_LOC_516/a_8_24# 0.01fF
C21768 AND2X1_LOC_320/a_8_24# OR2X1_LOC_532/B 0.01fF
C21769 VDD AND2X1_LOC_476/A -0.00fF
C21770 OR2X1_LOC_850/a_36_216# OR2X1_LOC_814/A 0.00fF
C21771 AND2X1_LOC_348/Y OR2X1_LOC_753/A 0.00fF
C21772 OR2X1_LOC_485/A AND2X1_LOC_114/a_8_24# 0.08fF
C21773 D_INPUT_7 INPUT_4 0.29fF
C21774 AND2X1_LOC_620/Y OR2X1_LOC_253/Y 0.03fF
C21775 OR2X1_LOC_185/A AND2X1_LOC_117/a_8_24# 0.02fF
C21776 AND2X1_LOC_727/Y OR2X1_LOC_152/a_8_216# 0.01fF
C21777 AND2X1_LOC_682/a_8_24# AND2X1_LOC_51/Y 0.01fF
C21778 OR2X1_LOC_835/a_36_216# OR2X1_LOC_269/B 0.01fF
C21779 OR2X1_LOC_364/B OR2X1_LOC_365/B 0.01fF
C21780 AND2X1_LOC_859/B OR2X1_LOC_59/Y 0.02fF
C21781 OR2X1_LOC_694/Y OR2X1_LOC_47/Y 0.13fF
C21782 OR2X1_LOC_290/a_8_216# INPUT_1 0.01fF
C21783 OR2X1_LOC_653/a_8_216# OR2X1_LOC_130/A 0.03fF
C21784 OR2X1_LOC_506/A AND2X1_LOC_51/Y 0.59fF
C21785 OR2X1_LOC_13/Y OR2X1_LOC_311/a_8_216# 0.01fF
C21786 VDD OR2X1_LOC_270/Y 0.24fF
C21787 OR2X1_LOC_671/Y OR2X1_LOC_28/a_8_216# -0.04fF
C21788 AND2X1_LOC_731/Y AND2X1_LOC_808/A 0.32fF
C21789 OR2X1_LOC_377/A OR2X1_LOC_97/a_36_216# 0.00fF
C21790 AND2X1_LOC_8/Y AND2X1_LOC_102/a_8_24# 0.01fF
C21791 AND2X1_LOC_7/B OR2X1_LOC_578/B 0.03fF
C21792 AND2X1_LOC_716/Y AND2X1_LOC_326/a_36_24# 0.01fF
C21793 OR2X1_LOC_585/A OR2X1_LOC_52/B 0.62fF
C21794 OR2X1_LOC_472/a_8_216# AND2X1_LOC_824/B 0.01fF
C21795 OR2X1_LOC_22/Y OR2X1_LOC_48/B 0.37fF
C21796 AND2X1_LOC_11/a_8_24# AND2X1_LOC_11/Y 0.00fF
C21797 AND2X1_LOC_327/a_36_24# OR2X1_LOC_18/Y 0.00fF
C21798 OR2X1_LOC_151/A OR2X1_LOC_675/Y 0.02fF
C21799 D_INPUT_7 AND2X1_LOC_51/A 0.34fF
C21800 OR2X1_LOC_122/Y D_INPUT_3 0.13fF
C21801 OR2X1_LOC_640/A AND2X1_LOC_47/Y 0.02fF
C21802 OR2X1_LOC_22/Y OR2X1_LOC_18/Y 0.92fF
C21803 OR2X1_LOC_682/Y OR2X1_LOC_743/A 0.38fF
C21804 OR2X1_LOC_103/Y AND2X1_LOC_866/A 0.03fF
C21805 OR2X1_LOC_274/Y OR2X1_LOC_276/A 0.01fF
C21806 OR2X1_LOC_613/Y AND2X1_LOC_663/B 0.01fF
C21807 OR2X1_LOC_66/A OR2X1_LOC_493/Y 0.01fF
C21808 OR2X1_LOC_473/Y OR2X1_LOC_87/A 0.08fF
C21809 OR2X1_LOC_726/a_8_216# OR2X1_LOC_731/A 0.03fF
C21810 AND2X1_LOC_842/B OR2X1_LOC_36/Y 0.00fF
C21811 OR2X1_LOC_626/a_8_216# OR2X1_LOC_617/Y 0.01fF
C21812 AND2X1_LOC_222/Y AND2X1_LOC_784/a_8_24# 0.01fF
C21813 OR2X1_LOC_589/A OR2X1_LOC_80/A 0.11fF
C21814 AND2X1_LOC_70/Y OR2X1_LOC_365/B 0.03fF
C21815 AND2X1_LOC_470/a_8_24# AND2X1_LOC_470/A 0.19fF
C21816 OR2X1_LOC_682/a_8_216# OR2X1_LOC_64/Y 0.02fF
C21817 OR2X1_LOC_377/A OR2X1_LOC_839/a_8_216# 0.03fF
C21818 OR2X1_LOC_327/a_8_216# OR2X1_LOC_218/Y 0.40fF
C21819 OR2X1_LOC_375/A OR2X1_LOC_814/A 0.51fF
C21820 OR2X1_LOC_373/Y OR2X1_LOC_164/a_8_216# 0.01fF
C21821 OR2X1_LOC_481/A OR2X1_LOC_89/A 0.06fF
C21822 OR2X1_LOC_43/A OR2X1_LOC_416/Y 0.03fF
C21823 AND2X1_LOC_47/Y AND2X1_LOC_297/a_8_24# 0.02fF
C21824 AND2X1_LOC_326/B AND2X1_LOC_222/Y 0.03fF
C21825 AND2X1_LOC_148/Y AND2X1_LOC_149/a_8_24# 0.00fF
C21826 OR2X1_LOC_550/B OR2X1_LOC_547/a_8_216# 0.01fF
C21827 AND2X1_LOC_641/Y AND2X1_LOC_650/a_8_24# 0.04fF
C21828 AND2X1_LOC_35/Y D_INPUT_0 0.35fF
C21829 AND2X1_LOC_523/a_8_24# AND2X1_LOC_851/B 0.01fF
C21830 OR2X1_LOC_494/Y AND2X1_LOC_563/Y 0.02fF
C21831 OR2X1_LOC_703/A OR2X1_LOC_365/B 0.35fF
C21832 OR2X1_LOC_3/Y AND2X1_LOC_307/Y 0.15fF
C21833 AND2X1_LOC_660/Y AND2X1_LOC_662/a_8_24# 0.09fF
C21834 AND2X1_LOC_712/B OR2X1_LOC_743/A 0.26fF
C21835 OR2X1_LOC_649/B OR2X1_LOC_655/B 0.04fF
C21836 OR2X1_LOC_549/A D_GATE_366 0.11fF
C21837 OR2X1_LOC_385/Y OR2X1_LOC_22/Y 0.04fF
C21838 AND2X1_LOC_471/Y AND2X1_LOC_222/Y 0.11fF
C21839 OR2X1_LOC_640/A OR2X1_LOC_598/A 0.01fF
C21840 AND2X1_LOC_851/B OR2X1_LOC_237/Y 0.06fF
C21841 OR2X1_LOC_26/Y OR2X1_LOC_71/Y 0.05fF
C21842 OR2X1_LOC_161/A OR2X1_LOC_284/B 0.03fF
C21843 OR2X1_LOC_856/a_8_216# OR2X1_LOC_19/B 0.07fF
C21844 AND2X1_LOC_796/a_8_24# OR2X1_LOC_437/A 0.01fF
C21845 OR2X1_LOC_161/A D_INPUT_1 0.13fF
C21846 OR2X1_LOC_681/Y AND2X1_LOC_685/a_8_24# 0.23fF
C21847 AND2X1_LOC_793/Y AND2X1_LOC_805/Y 0.01fF
C21848 OR2X1_LOC_287/B OR2X1_LOC_532/B 0.05fF
C21849 AND2X1_LOC_41/A AND2X1_LOC_751/a_8_24# 0.03fF
C21850 AND2X1_LOC_388/a_8_24# AND2X1_LOC_810/a_8_24# 0.23fF
C21851 OR2X1_LOC_638/a_8_216# AND2X1_LOC_31/Y 0.01fF
C21852 OR2X1_LOC_71/Y OR2X1_LOC_89/A 0.04fF
C21853 OR2X1_LOC_70/Y AND2X1_LOC_686/a_36_24# 0.00fF
C21854 D_INPUT_0 OR2X1_LOC_74/A 0.10fF
C21855 OR2X1_LOC_605/B OR2X1_LOC_814/A 0.02fF
C21856 OR2X1_LOC_312/Y AND2X1_LOC_170/B 0.04fF
C21857 OR2X1_LOC_696/A AND2X1_LOC_786/Y 0.07fF
C21858 OR2X1_LOC_48/B OR2X1_LOC_387/a_8_216# 0.05fF
C21859 OR2X1_LOC_696/A OR2X1_LOC_323/a_8_216# 0.01fF
C21860 AND2X1_LOC_242/B OR2X1_LOC_184/a_8_216# 0.05fF
C21861 AND2X1_LOC_740/B GATE_811 0.00fF
C21862 AND2X1_LOC_857/Y OR2X1_LOC_172/Y 0.02fF
C21863 AND2X1_LOC_12/Y AND2X1_LOC_761/a_8_24# 0.01fF
C21864 OR2X1_LOC_404/Y OR2X1_LOC_62/B 0.02fF
C21865 AND2X1_LOC_92/Y OR2X1_LOC_704/a_8_216# 0.02fF
C21866 OR2X1_LOC_429/Y OR2X1_LOC_70/a_36_216# 0.01fF
C21867 AND2X1_LOC_40/Y OR2X1_LOC_68/B 0.77fF
C21868 AND2X1_LOC_580/A AND2X1_LOC_624/B 0.03fF
C21869 OR2X1_LOC_87/A OR2X1_LOC_214/B 0.01fF
C21870 OR2X1_LOC_115/B OR2X1_LOC_161/B 0.08fF
C21871 OR2X1_LOC_95/Y AND2X1_LOC_276/Y 0.00fF
C21872 AND2X1_LOC_618/a_8_24# OR2X1_LOC_80/A 0.11fF
C21873 OR2X1_LOC_246/A OR2X1_LOC_54/Y 0.00fF
C21874 OR2X1_LOC_287/B OR2X1_LOC_343/B 0.01fF
C21875 OR2X1_LOC_406/a_8_216# OR2X1_LOC_406/A 0.01fF
C21876 OR2X1_LOC_45/B AND2X1_LOC_476/a_8_24# 0.01fF
C21877 OR2X1_LOC_76/A OR2X1_LOC_532/B 0.03fF
C21878 OR2X1_LOC_160/B OR2X1_LOC_333/A 0.01fF
C21879 AND2X1_LOC_208/Y AND2X1_LOC_219/A 0.16fF
C21880 VDD OR2X1_LOC_388/a_8_216# 0.21fF
C21881 AND2X1_LOC_358/a_8_24# OR2X1_LOC_417/A 0.10fF
C21882 OR2X1_LOC_375/a_8_216# OR2X1_LOC_375/Y 0.02fF
C21883 OR2X1_LOC_175/Y OR2X1_LOC_390/A 0.01fF
C21884 OR2X1_LOC_503/A AND2X1_LOC_657/A 0.01fF
C21885 AND2X1_LOC_227/Y OR2X1_LOC_245/a_36_216# 0.00fF
C21886 OR2X1_LOC_53/Y OR2X1_LOC_13/Y 0.16fF
C21887 OR2X1_LOC_673/Y OR2X1_LOC_398/Y 0.01fF
C21888 AND2X1_LOC_420/a_8_24# AND2X1_LOC_51/Y 0.02fF
C21889 OR2X1_LOC_87/Y OR2X1_LOC_68/B 0.02fF
C21890 OR2X1_LOC_479/a_36_216# OR2X1_LOC_223/A 0.00fF
C21891 OR2X1_LOC_45/B OR2X1_LOC_693/a_36_216# 0.02fF
C21892 AND2X1_LOC_259/Y AND2X1_LOC_259/a_36_24# 0.00fF
C21893 OR2X1_LOC_848/A OR2X1_LOC_68/B 0.01fF
C21894 OR2X1_LOC_385/Y OR2X1_LOC_387/a_8_216# 0.40fF
C21895 AND2X1_LOC_249/a_8_24# OR2X1_LOC_595/A 0.00fF
C21896 OR2X1_LOC_794/a_8_216# OR2X1_LOC_374/Y 0.04fF
C21897 AND2X1_LOC_51/a_8_24# INPUT_6 0.01fF
C21898 OR2X1_LOC_449/B OR2X1_LOC_779/B 0.03fF
C21899 OR2X1_LOC_160/B OR2X1_LOC_392/B 0.10fF
C21900 OR2X1_LOC_312/Y OR2X1_LOC_331/Y 0.51fF
C21901 AND2X1_LOC_164/a_8_24# OR2X1_LOC_390/B 0.03fF
C21902 OR2X1_LOC_436/Y OR2X1_LOC_532/B 0.03fF
C21903 OR2X1_LOC_765/a_8_216# OR2X1_LOC_16/A 0.06fF
C21904 OR2X1_LOC_19/B AND2X1_LOC_6/a_8_24# 0.09fF
C21905 OR2X1_LOC_516/Y OR2X1_LOC_516/B 0.01fF
C21906 OR2X1_LOC_151/A OR2X1_LOC_736/Y 0.49fF
C21907 AND2X1_LOC_41/A OR2X1_LOC_731/A 0.27fF
C21908 AND2X1_LOC_64/Y OR2X1_LOC_632/Y 0.15fF
C21909 AND2X1_LOC_56/B OR2X1_LOC_71/A 0.01fF
C21910 OR2X1_LOC_64/Y AND2X1_LOC_644/a_8_24# 0.01fF
C21911 AND2X1_LOC_772/B AND2X1_LOC_554/a_8_24# 0.03fF
C21912 OR2X1_LOC_339/a_8_216# AND2X1_LOC_22/Y 0.01fF
C21913 AND2X1_LOC_842/B OR2X1_LOC_419/Y 0.03fF
C21914 AND2X1_LOC_53/Y OR2X1_LOC_200/Y 0.03fF
C21915 AND2X1_LOC_18/Y AND2X1_LOC_256/a_8_24# 0.05fF
C21916 OR2X1_LOC_40/Y AND2X1_LOC_469/a_8_24# 0.04fF
C21917 AND2X1_LOC_319/A OR2X1_LOC_13/B 0.02fF
C21918 OR2X1_LOC_634/a_8_216# OR2X1_LOC_334/A 0.47fF
C21919 AND2X1_LOC_8/Y OR2X1_LOC_71/A 0.13fF
C21920 AND2X1_LOC_182/A AND2X1_LOC_182/a_8_24# 0.10fF
C21921 OR2X1_LOC_624/A OR2X1_LOC_175/a_8_216# 0.03fF
C21922 OR2X1_LOC_159/a_8_216# OR2X1_LOC_158/A 0.02fF
C21923 AND2X1_LOC_784/A OR2X1_LOC_437/A 0.16fF
C21924 OR2X1_LOC_536/Y OR2X1_LOC_829/A 0.11fF
C21925 OR2X1_LOC_604/A AND2X1_LOC_704/a_8_24# 0.02fF
C21926 OR2X1_LOC_40/Y OR2X1_LOC_158/A 1.67fF
C21927 OR2X1_LOC_45/B OR2X1_LOC_531/Y 0.02fF
C21928 OR2X1_LOC_541/B AND2X1_LOC_36/Y 0.00fF
C21929 AND2X1_LOC_727/A AND2X1_LOC_486/a_8_24# 0.01fF
C21930 AND2X1_LOC_617/a_8_24# AND2X1_LOC_36/Y 0.01fF
C21931 OR2X1_LOC_22/Y AND2X1_LOC_215/A 0.06fF
C21932 OR2X1_LOC_161/A OR2X1_LOC_180/B 0.03fF
C21933 OR2X1_LOC_44/Y OR2X1_LOC_424/Y 0.02fF
C21934 AND2X1_LOC_531/a_8_24# OR2X1_LOC_562/A 0.01fF
C21935 OR2X1_LOC_160/B OR2X1_LOC_113/B 0.20fF
C21936 OR2X1_LOC_475/Y OR2X1_LOC_68/B 0.02fF
C21937 OR2X1_LOC_468/Y OR2X1_LOC_777/B 0.03fF
C21938 OR2X1_LOC_607/a_8_216# OR2X1_LOC_67/Y 0.02fF
C21939 OR2X1_LOC_31/Y OR2X1_LOC_3/B 0.07fF
C21940 AND2X1_LOC_216/Y AND2X1_LOC_217/Y 0.01fF
C21941 OR2X1_LOC_92/a_8_216# D_INPUT_1 0.07fF
C21942 OR2X1_LOC_121/B OR2X1_LOC_779/B 0.03fF
C21943 OR2X1_LOC_64/Y AND2X1_LOC_657/A 0.03fF
C21944 OR2X1_LOC_291/A OR2X1_LOC_71/A 0.08fF
C21945 D_INPUT_0 AND2X1_LOC_647/Y 0.03fF
C21946 OR2X1_LOC_44/Y D_INPUT_6 0.02fF
C21947 AND2X1_LOC_702/Y OR2X1_LOC_320/a_36_216# 0.00fF
C21948 AND2X1_LOC_95/Y OR2X1_LOC_556/a_8_216# 0.02fF
C21949 OR2X1_LOC_19/B OR2X1_LOC_198/A 0.03fF
C21950 OR2X1_LOC_160/B OR2X1_LOC_450/A 0.11fF
C21951 OR2X1_LOC_316/a_8_216# OR2X1_LOC_32/B 0.03fF
C21952 AND2X1_LOC_534/a_36_24# OR2X1_LOC_538/A 0.00fF
C21953 AND2X1_LOC_675/A OR2X1_LOC_406/A 0.02fF
C21954 OR2X1_LOC_840/A OR2X1_LOC_161/B 0.05fF
C21955 OR2X1_LOC_45/B OR2X1_LOC_46/a_8_216# 0.02fF
C21956 AND2X1_LOC_658/A AND2X1_LOC_658/a_8_24# 0.01fF
C21957 OR2X1_LOC_89/A AND2X1_LOC_789/Y 0.00fF
C21958 AND2X1_LOC_12/Y OR2X1_LOC_773/Y 0.01fF
C21959 AND2X1_LOC_535/Y OR2X1_LOC_744/A 0.03fF
C21960 AND2X1_LOC_41/A OR2X1_LOC_596/a_8_216# 0.01fF
C21961 VDD OR2X1_LOC_122/A -0.00fF
C21962 AND2X1_LOC_43/B AND2X1_LOC_416/a_36_24# 0.01fF
C21963 OR2X1_LOC_123/a_8_216# OR2X1_LOC_124/A 0.01fF
C21964 AND2X1_LOC_22/Y OR2X1_LOC_624/A 0.12fF
C21965 OR2X1_LOC_151/A OR2X1_LOC_808/B 0.10fF
C21966 OR2X1_LOC_6/B AND2X1_LOC_41/A 0.07fF
C21967 AND2X1_LOC_207/a_8_24# AND2X1_LOC_207/B 0.01fF
C21968 OR2X1_LOC_417/A AND2X1_LOC_657/A 0.17fF
C21969 OR2X1_LOC_820/Y AND2X1_LOC_789/Y 0.03fF
C21970 VDD INPUT_0 0.83fF
C21971 OR2X1_LOC_40/Y AND2X1_LOC_98/Y 0.01fF
C21972 AND2X1_LOC_657/Y AND2X1_LOC_659/a_8_24# 0.29fF
C21973 OR2X1_LOC_742/B AND2X1_LOC_613/a_8_24# 0.23fF
C21974 AND2X1_LOC_717/a_8_24# AND2X1_LOC_786/Y 0.04fF
C21975 OR2X1_LOC_121/a_8_216# OR2X1_LOC_506/A 0.00fF
C21976 AND2X1_LOC_534/a_8_24# OR2X1_LOC_620/Y 0.01fF
C21977 AND2X1_LOC_738/B OR2X1_LOC_59/Y 0.07fF
C21978 OR2X1_LOC_566/A OR2X1_LOC_468/Y 0.02fF
C21979 OR2X1_LOC_315/Y AND2X1_LOC_445/a_8_24# 0.11fF
C21980 AND2X1_LOC_509/a_8_24# OR2X1_LOC_59/Y 0.02fF
C21981 OR2X1_LOC_647/Y OR2X1_LOC_771/B 0.08fF
C21982 OR2X1_LOC_139/A OR2X1_LOC_510/Y 0.11fF
C21983 OR2X1_LOC_56/A OR2X1_LOC_59/Y 8.72fF
C21984 AND2X1_LOC_710/Y OR2X1_LOC_59/Y 0.01fF
C21985 OR2X1_LOC_624/A AND2X1_LOC_417/a_36_24# 0.01fF
C21986 OR2X1_LOC_691/A OR2X1_LOC_160/A 0.03fF
C21987 OR2X1_LOC_396/Y OR2X1_LOC_598/A 0.31fF
C21988 AND2X1_LOC_91/B OR2X1_LOC_864/A 0.07fF
C21989 OR2X1_LOC_158/A AND2X1_LOC_843/Y 0.02fF
C21990 AND2X1_LOC_1/Y D_INPUT_6 0.01fF
C21991 AND2X1_LOC_43/B OR2X1_LOC_138/A 0.01fF
C21992 OR2X1_LOC_744/A OR2X1_LOC_484/Y 0.10fF
C21993 OR2X1_LOC_91/A AND2X1_LOC_434/Y 0.07fF
C21994 AND2X1_LOC_564/B AND2X1_LOC_374/Y 1.23fF
C21995 AND2X1_LOC_95/Y OR2X1_LOC_346/A 0.00fF
C21996 OR2X1_LOC_348/Y OR2X1_LOC_850/B 0.02fF
C21997 OR2X1_LOC_91/A AND2X1_LOC_219/Y 0.53fF
C21998 OR2X1_LOC_45/B OR2X1_LOC_406/a_36_216# 0.00fF
C21999 OR2X1_LOC_316/Y OR2X1_LOC_16/A 0.05fF
C22000 AND2X1_LOC_458/Y AND2X1_LOC_786/Y 0.02fF
C22001 AND2X1_LOC_51/Y OR2X1_LOC_180/B 0.03fF
C22002 OR2X1_LOC_696/A AND2X1_LOC_578/A 0.14fF
C22003 AND2X1_LOC_231/Y OR2X1_LOC_6/A 0.01fF
C22004 INPUT_3 OR2X1_LOC_671/Y 0.09fF
C22005 OR2X1_LOC_349/a_8_216# OR2X1_LOC_850/B 0.01fF
C22006 OR2X1_LOC_833/Y AND2X1_LOC_59/Y 0.02fF
C22007 OR2X1_LOC_2/Y OR2X1_LOC_581/Y 0.04fF
C22008 AND2X1_LOC_662/B AND2X1_LOC_476/Y 0.08fF
C22009 OR2X1_LOC_256/Y OR2X1_LOC_51/Y 0.12fF
C22010 OR2X1_LOC_230/Y OR2X1_LOC_52/B 0.00fF
C22011 OR2X1_LOC_271/B AND2X1_LOC_786/Y 0.06fF
C22012 VDD OR2X1_LOC_772/B -0.00fF
C22013 AND2X1_LOC_714/B AND2X1_LOC_452/Y 0.01fF
C22014 AND2X1_LOC_364/a_8_24# OR2X1_LOC_6/A 0.01fF
C22015 OR2X1_LOC_499/B OR2X1_LOC_78/A 0.02fF
C22016 OR2X1_LOC_860/Y VDD -0.00fF
C22017 AND2X1_LOC_110/Y OR2X1_LOC_620/Y 0.01fF
C22018 AND2X1_LOC_742/a_8_24# AND2X1_LOC_192/Y 0.02fF
C22019 AND2X1_LOC_717/Y VDD 0.09fF
C22020 OR2X1_LOC_244/Y OR2X1_LOC_721/Y 0.07fF
C22021 OR2X1_LOC_833/B OR2X1_LOC_629/B 0.07fF
C22022 OR2X1_LOC_663/A AND2X1_LOC_103/a_8_24# 0.03fF
C22023 OR2X1_LOC_485/Y OR2X1_LOC_48/B 0.16fF
C22024 OR2X1_LOC_287/B OR2X1_LOC_392/a_36_216# 0.00fF
C22025 AND2X1_LOC_56/B OR2X1_LOC_355/a_8_216# 0.03fF
C22026 OR2X1_LOC_26/Y OR2X1_LOC_585/a_8_216# 0.04fF
C22027 AND2X1_LOC_170/B OR2X1_LOC_13/B 0.00fF
C22028 AND2X1_LOC_544/Y AND2X1_LOC_728/a_8_24# 0.03fF
C22029 OR2X1_LOC_368/a_36_216# OR2X1_LOC_109/Y 0.01fF
C22030 OR2X1_LOC_654/A AND2X1_LOC_7/B 0.00fF
C22031 OR2X1_LOC_502/A OR2X1_LOC_834/A 0.31fF
C22032 OR2X1_LOC_121/Y OR2X1_LOC_203/Y 0.02fF
C22033 OR2X1_LOC_204/Y AND2X1_LOC_65/A 0.01fF
C22034 OR2X1_LOC_494/A OR2X1_LOC_3/Y 0.01fF
C22035 AND2X1_LOC_364/Y AND2X1_LOC_863/a_8_24# 0.01fF
C22036 INPUT_0 OR2X1_LOC_689/A 0.03fF
C22037 OR2X1_LOC_589/A OR2X1_LOC_6/A 0.02fF
C22038 OR2X1_LOC_529/Y OR2X1_LOC_816/A 0.05fF
C22039 AND2X1_LOC_158/a_8_24# OR2X1_LOC_160/Y 0.24fF
C22040 VDD OR2X1_LOC_732/B 0.04fF
C22041 OR2X1_LOC_229/a_8_216# OR2X1_LOC_52/B -0.03fF
C22042 OR2X1_LOC_709/A OR2X1_LOC_449/B 0.09fF
C22043 VDD OR2X1_LOC_789/B 0.00fF
C22044 AND2X1_LOC_733/Y AND2X1_LOC_737/a_8_24# -0.00fF
C22045 OR2X1_LOC_440/a_36_216# OR2X1_LOC_161/A 0.02fF
C22046 AND2X1_LOC_526/a_8_24# OR2X1_LOC_469/Y 0.07fF
C22047 AND2X1_LOC_59/Y AND2X1_LOC_387/a_8_24# 0.01fF
C22048 OR2X1_LOC_64/Y OR2X1_LOC_503/a_36_216# 0.03fF
C22049 AND2X1_LOC_702/Y AND2X1_LOC_566/B 0.00fF
C22050 OR2X1_LOC_154/A AND2X1_LOC_110/Y 0.03fF
C22051 AND2X1_LOC_59/Y OR2X1_LOC_493/B 0.23fF
C22052 AND2X1_LOC_850/Y OR2X1_LOC_59/Y 0.07fF
C22053 VDD OR2X1_LOC_11/Y 0.35fF
C22054 OR2X1_LOC_53/a_8_216# OR2X1_LOC_25/Y 0.01fF
C22055 OR2X1_LOC_492/a_8_216# AND2X1_LOC_717/B 0.47fF
C22056 OR2X1_LOC_492/Y AND2X1_LOC_493/a_8_24# 0.01fF
C22057 OR2X1_LOC_325/B OR2X1_LOC_87/A 0.03fF
C22058 OR2X1_LOC_319/a_8_216# OR2X1_LOC_538/A 0.01fF
C22059 INPUT_0 OR2X1_LOC_829/a_8_216# 0.01fF
C22060 OR2X1_LOC_686/B OR2X1_LOC_87/A 0.00fF
C22061 OR2X1_LOC_375/A OR2X1_LOC_244/Y 1.57fF
C22062 AND2X1_LOC_390/B OR2X1_LOC_16/A 0.07fF
C22063 OR2X1_LOC_70/Y OR2X1_LOC_118/a_8_216# 0.03fF
C22064 OR2X1_LOC_158/A OR2X1_LOC_7/A 0.28fF
C22065 AND2X1_LOC_721/A OR2X1_LOC_13/B 0.06fF
C22066 OR2X1_LOC_792/Y OR2X1_LOC_285/a_8_216# 0.02fF
C22067 OR2X1_LOC_318/Y OR2X1_LOC_798/Y 0.05fF
C22068 OR2X1_LOC_51/Y AND2X1_LOC_470/A 0.03fF
C22069 OR2X1_LOC_600/A AND2X1_LOC_818/a_8_24# 0.06fF
C22070 OR2X1_LOC_175/Y OR2X1_LOC_750/A 0.03fF
C22071 OR2X1_LOC_624/A OR2X1_LOC_244/B 0.07fF
C22072 OR2X1_LOC_377/A OR2X1_LOC_538/A 0.01fF
C22073 OR2X1_LOC_491/a_8_216# OR2X1_LOC_529/Y 0.01fF
C22074 VDD AND2X1_LOC_560/B 0.55fF
C22075 AND2X1_LOC_784/A AND2X1_LOC_715/A 0.02fF
C22076 AND2X1_LOC_357/A AND2X1_LOC_211/B 0.02fF
C22077 AND2X1_LOC_60/a_8_24# OR2X1_LOC_476/B 0.03fF
C22078 OR2X1_LOC_52/Y AND2X1_LOC_219/A 0.15fF
C22079 OR2X1_LOC_216/A OR2X1_LOC_493/A 0.13fF
C22080 VDD OR2X1_LOC_173/Y 0.12fF
C22081 VDD OR2X1_LOC_690/A 0.68fF
C22082 OR2X1_LOC_816/a_8_216# OR2X1_LOC_36/Y 0.01fF
C22083 AND2X1_LOC_86/Y OR2X1_LOC_100/Y 0.02fF
C22084 OR2X1_LOC_858/A AND2X1_LOC_56/B 0.63fF
C22085 OR2X1_LOC_426/B OR2X1_LOC_26/Y 0.10fF
C22086 OR2X1_LOC_158/A OR2X1_LOC_44/a_8_216# 0.02fF
C22087 AND2X1_LOC_92/a_8_24# OR2X1_LOC_46/A 0.03fF
C22088 OR2X1_LOC_696/A AND2X1_LOC_841/a_8_24# 0.03fF
C22089 AND2X1_LOC_70/Y OR2X1_LOC_449/B 0.00fF
C22090 OR2X1_LOC_532/B OR2X1_LOC_722/B 0.02fF
C22091 AND2X1_LOC_576/Y OR2X1_LOC_744/A 0.07fF
C22092 OR2X1_LOC_74/A AND2X1_LOC_784/a_8_24# 0.01fF
C22093 OR2X1_LOC_56/A OR2X1_LOC_820/B 0.02fF
C22094 OR2X1_LOC_377/A D_INPUT_5 0.06fF
C22095 VDD AND2X1_LOC_528/a_8_24# -0.00fF
C22096 OR2X1_LOC_441/Y AND2X1_LOC_807/Y 0.02fF
C22097 OR2X1_LOC_405/A OR2X1_LOC_785/B 0.01fF
C22098 AND2X1_LOC_859/Y AND2X1_LOC_663/A 0.10fF
C22099 OR2X1_LOC_709/A OR2X1_LOC_121/B 0.07fF
C22100 AND2X1_LOC_537/a_36_24# OR2X1_LOC_7/A 0.01fF
C22101 AND2X1_LOC_31/Y OR2X1_LOC_446/B 0.06fF
C22102 AND2X1_LOC_794/B OR2X1_LOC_64/Y 0.07fF
C22103 AND2X1_LOC_340/Y OR2X1_LOC_22/Y 0.07fF
C22104 OR2X1_LOC_715/a_8_216# OR2X1_LOC_446/B 0.01fF
C22105 OR2X1_LOC_426/B OR2X1_LOC_89/A 1.36fF
C22106 AND2X1_LOC_123/Y OR2X1_LOC_92/Y 0.29fF
C22107 AND2X1_LOC_326/B OR2X1_LOC_74/A 0.00fF
C22108 OR2X1_LOC_22/Y AND2X1_LOC_810/B 0.07fF
C22109 AND2X1_LOC_560/a_8_24# OR2X1_LOC_47/Y 0.17fF
C22110 OR2X1_LOC_161/A OR2X1_LOC_737/A 0.03fF
C22111 OR2X1_LOC_13/B OR2X1_LOC_331/Y 1.09fF
C22112 AND2X1_LOC_669/a_8_24# OR2X1_LOC_721/Y 0.03fF
C22113 OR2X1_LOC_561/Y OR2X1_LOC_269/B 0.03fF
C22114 INPUT_3 AND2X1_LOC_820/a_8_24# 0.06fF
C22115 OR2X1_LOC_814/A OR2X1_LOC_843/B 0.58fF
C22116 OR2X1_LOC_147/B OR2X1_LOC_375/A 0.05fF
C22117 OR2X1_LOC_804/A OR2X1_LOC_776/A 0.01fF
C22118 AND2X1_LOC_99/A OR2X1_LOC_118/Y 0.02fF
C22119 AND2X1_LOC_12/Y AND2X1_LOC_16/a_8_24# 0.01fF
C22120 AND2X1_LOC_70/Y OR2X1_LOC_636/A 0.01fF
C22121 AND2X1_LOC_378/a_8_24# OR2X1_LOC_585/A 0.01fF
C22122 AND2X1_LOC_47/Y OR2X1_LOC_576/A 0.03fF
C22123 OR2X1_LOC_168/B OR2X1_LOC_574/A 0.17fF
C22124 OR2X1_LOC_287/B OR2X1_LOC_624/Y 0.16fF
C22125 AND2X1_LOC_181/Y OR2X1_LOC_22/Y 1.44fF
C22126 OR2X1_LOC_469/Y OR2X1_LOC_87/A 0.07fF
C22127 AND2X1_LOC_95/Y OR2X1_LOC_161/A 0.72fF
C22128 OR2X1_LOC_287/B OR2X1_LOC_78/a_36_216# 0.00fF
C22129 OR2X1_LOC_47/a_8_216# OR2X1_LOC_25/Y 0.09fF
C22130 OR2X1_LOC_48/B OR2X1_LOC_39/A 0.07fF
C22131 AND2X1_LOC_654/B OR2X1_LOC_6/A 0.00fF
C22132 AND2X1_LOC_139/B AND2X1_LOC_649/a_8_24# 0.04fF
C22133 OR2X1_LOC_814/A OR2X1_LOC_549/A 0.15fF
C22134 AND2X1_LOC_711/Y OR2X1_LOC_56/A 0.03fF
C22135 OR2X1_LOC_61/Y OR2X1_LOC_222/A 0.03fF
C22136 AND2X1_LOC_738/B OR2X1_LOC_70/Y 0.25fF
C22137 AND2X1_LOC_710/Y AND2X1_LOC_711/Y 0.01fF
C22138 AND2X1_LOC_749/a_8_24# AND2X1_LOC_8/Y 0.11fF
C22139 VDD OR2X1_LOC_401/A 0.21fF
C22140 OR2X1_LOC_70/Y OR2X1_LOC_56/A 0.11fF
C22141 AND2X1_LOC_857/Y OR2X1_LOC_52/B 0.10fF
C22142 VDD OR2X1_LOC_64/Y 1.98fF
C22143 OR2X1_LOC_545/A OR2X1_LOC_471/Y 0.02fF
C22144 OR2X1_LOC_18/Y OR2X1_LOC_39/A 0.31fF
C22145 OR2X1_LOC_9/Y OR2X1_LOC_62/B 0.01fF
C22146 AND2X1_LOC_98/Y OR2X1_LOC_7/A 0.02fF
C22147 AND2X1_LOC_12/Y OR2X1_LOC_377/A 0.12fF
C22148 OR2X1_LOC_376/Y OR2X1_LOC_378/A 0.88fF
C22149 AND2X1_LOC_506/a_8_24# OR2X1_LOC_239/Y 0.23fF
C22150 OR2X1_LOC_62/B OR2X1_LOC_362/A 0.03fF
C22151 OR2X1_LOC_689/A OR2X1_LOC_690/A 0.03fF
C22152 OR2X1_LOC_49/A OR2X1_LOC_96/a_8_216# 0.01fF
C22153 AND2X1_LOC_398/a_8_24# OR2X1_LOC_6/A 0.06fF
C22154 AND2X1_LOC_841/B OR2X1_LOC_44/Y 0.01fF
C22155 OR2X1_LOC_31/Y OR2X1_LOC_584/a_8_216# 0.01fF
C22156 OR2X1_LOC_405/A OR2X1_LOC_687/Y 0.01fF
C22157 AND2X1_LOC_794/B OR2X1_LOC_417/A 0.02fF
C22158 AND2X1_LOC_851/B OR2X1_LOC_522/a_8_216# 0.02fF
C22159 AND2X1_LOC_95/Y AND2X1_LOC_25/Y 0.02fF
C22160 AND2X1_LOC_70/Y OR2X1_LOC_121/B 0.09fF
C22161 AND2X1_LOC_663/B AND2X1_LOC_218/Y 0.23fF
C22162 OR2X1_LOC_676/Y AND2X1_LOC_48/A 0.07fF
C22163 AND2X1_LOC_47/Y OR2X1_LOC_439/B 0.00fF
C22164 OR2X1_LOC_643/A OR2X1_LOC_560/a_36_216# 0.00fF
C22165 OR2X1_LOC_518/a_8_216# AND2X1_LOC_222/Y 0.04fF
C22166 AND2X1_LOC_514/Y OR2X1_LOC_56/A 0.09fF
C22167 AND2X1_LOC_199/a_8_24# AND2X1_LOC_207/A 0.00fF
C22168 AND2X1_LOC_12/Y OR2X1_LOC_203/Y 0.07fF
C22169 AND2X1_LOC_838/Y OR2X1_LOC_85/A 0.01fF
C22170 OR2X1_LOC_585/A OR2X1_LOC_394/Y 0.03fF
C22171 OR2X1_LOC_158/A OR2X1_LOC_224/a_8_216# 0.05fF
C22172 VDD AND2X1_LOC_632/A 0.06fF
C22173 AND2X1_LOC_211/B OR2X1_LOC_48/B 0.05fF
C22174 OR2X1_LOC_160/B OR2X1_LOC_532/B 0.11fF
C22175 OR2X1_LOC_404/Y OR2X1_LOC_659/A 0.02fF
C22176 OR2X1_LOC_834/A AND2X1_LOC_48/A 0.02fF
C22177 OR2X1_LOC_6/B OR2X1_LOC_95/Y 0.07fF
C22178 OR2X1_LOC_679/A OR2X1_LOC_679/Y 0.07fF
C22179 VDD OR2X1_LOC_417/A 1.16fF
C22180 AND2X1_LOC_211/B OR2X1_LOC_18/Y 0.04fF
C22181 OR2X1_LOC_703/A OR2X1_LOC_121/B 0.05fF
C22182 OR2X1_LOC_3/Y OR2X1_LOC_427/A 0.16fF
C22183 OR2X1_LOC_70/Y OR2X1_LOC_426/Y 0.01fF
C22184 OR2X1_LOC_849/a_36_216# OR2X1_LOC_624/Y 0.00fF
C22185 OR2X1_LOC_299/a_36_216# OR2X1_LOC_619/Y 0.01fF
C22186 OR2X1_LOC_247/a_36_216# OR2X1_LOC_161/B 0.00fF
C22187 OR2X1_LOC_247/Y AND2X1_LOC_44/Y 0.00fF
C22188 OR2X1_LOC_504/Y OR2X1_LOC_56/A 0.00fF
C22189 OR2X1_LOC_283/a_8_216# AND2X1_LOC_859/Y 0.03fF
C22190 OR2X1_LOC_285/A OR2X1_LOC_269/B 0.00fF
C22191 OR2X1_LOC_43/A OR2X1_LOC_6/A 0.19fF
C22192 AND2X1_LOC_59/Y OR2X1_LOC_574/A 0.06fF
C22193 OR2X1_LOC_564/a_8_216# OR2X1_LOC_192/B 0.05fF
C22194 OR2X1_LOC_377/A AND2X1_LOC_79/Y 0.01fF
C22195 OR2X1_LOC_336/a_8_216# OR2X1_LOC_365/B 0.14fF
C22196 OR2X1_LOC_97/B AND2X1_LOC_89/a_36_24# 0.01fF
C22197 OR2X1_LOC_132/a_8_216# AND2X1_LOC_227/Y 0.01fF
C22198 OR2X1_LOC_426/B OR2X1_LOC_92/a_8_216# 0.03fF
C22199 AND2X1_LOC_51/Y OR2X1_LOC_737/A 0.07fF
C22200 AND2X1_LOC_387/B OR2X1_LOC_375/A 0.03fF
C22201 OR2X1_LOC_689/Y OR2X1_LOC_690/Y 0.09fF
C22202 OR2X1_LOC_828/Y OR2X1_LOC_198/A 0.17fF
C22203 OR2X1_LOC_474/Y OR2X1_LOC_62/B 0.05fF
C22204 OR2X1_LOC_479/Y AND2X1_LOC_43/B 0.07fF
C22205 OR2X1_LOC_426/B OR2X1_LOC_426/a_8_216# 0.07fF
C22206 OR2X1_LOC_624/B OR2X1_LOC_404/a_8_216# 0.05fF
C22207 OR2X1_LOC_273/a_8_216# OR2X1_LOC_316/Y 0.00fF
C22208 OR2X1_LOC_273/Y OR2X1_LOC_595/a_8_216# 0.02fF
C22209 AND2X1_LOC_95/Y AND2X1_LOC_51/Y 0.82fF
C22210 AND2X1_LOC_367/a_8_24# OR2X1_LOC_89/A 0.01fF
C22211 OR2X1_LOC_527/Y AND2X1_LOC_621/Y 0.07fF
C22212 OR2X1_LOC_829/a_8_216# OR2X1_LOC_64/Y 0.14fF
C22213 AND2X1_LOC_578/A AND2X1_LOC_458/Y 0.09fF
C22214 AND2X1_LOC_41/A AND2X1_LOC_47/Y 0.22fF
C22215 OR2X1_LOC_119/a_8_216# AND2X1_LOC_573/A 0.03fF
C22216 OR2X1_LOC_427/A OR2X1_LOC_582/Y 0.01fF
C22217 AND2X1_LOC_858/B AND2X1_LOC_851/B 0.24fF
C22218 AND2X1_LOC_346/a_8_24# AND2X1_LOC_848/A 0.02fF
C22219 OR2X1_LOC_472/a_8_216# OR2X1_LOC_375/A 0.06fF
C22220 AND2X1_LOC_496/a_8_24# OR2X1_LOC_203/Y 0.00fF
C22221 AND2X1_LOC_522/a_36_24# OR2X1_LOC_560/A 0.00fF
C22222 OR2X1_LOC_813/A OR2X1_LOC_92/Y 0.01fF
C22223 OR2X1_LOC_665/a_8_216# AND2X1_LOC_624/A 0.06fF
C22224 OR2X1_LOC_508/Y AND2X1_LOC_239/a_8_24# 0.24fF
C22225 OR2X1_LOC_3/Y AND2X1_LOC_363/A 0.00fF
C22226 OR2X1_LOC_748/A AND2X1_LOC_847/a_8_24# 0.00fF
C22227 AND2X1_LOC_137/a_8_24# OR2X1_LOC_517/A 0.05fF
C22228 OR2X1_LOC_580/B OR2X1_LOC_578/B 0.00fF
C22229 OR2X1_LOC_856/B AND2X1_LOC_23/a_36_24# 0.01fF
C22230 AND2X1_LOC_17/Y OR2X1_LOC_636/A 0.01fF
C22231 OR2X1_LOC_654/a_8_216# OR2X1_LOC_68/B 0.01fF
C22232 AND2X1_LOC_390/B AND2X1_LOC_336/a_8_24# 0.02fF
C22233 AND2X1_LOC_477/A AND2X1_LOC_452/Y 0.01fF
C22234 AND2X1_LOC_470/a_8_24# AND2X1_LOC_470/B 0.01fF
C22235 OR2X1_LOC_520/Y OR2X1_LOC_520/B 1.08fF
C22236 OR2X1_LOC_462/B AND2X1_LOC_518/a_8_24# 0.01fF
C22237 OR2X1_LOC_504/Y AND2X1_LOC_850/Y 0.18fF
C22238 AND2X1_LOC_228/Y OR2X1_LOC_22/Y 0.03fF
C22239 AND2X1_LOC_863/Y AND2X1_LOC_661/a_8_24# -0.01fF
C22240 INPUT_3 OR2X1_LOC_532/B 0.57fF
C22241 OR2X1_LOC_339/A OR2X1_LOC_174/a_8_216# 0.01fF
C22242 OR2X1_LOC_462/B AND2X1_LOC_48/A 0.03fF
C22243 OR2X1_LOC_109/Y OR2X1_LOC_111/Y 0.40fF
C22244 OR2X1_LOC_813/A OR2X1_LOC_65/B 0.00fF
C22245 OR2X1_LOC_251/Y OR2X1_LOC_64/Y 0.07fF
C22246 OR2X1_LOC_36/Y AND2X1_LOC_856/a_36_24# 0.01fF
C22247 OR2X1_LOC_45/B OR2X1_LOC_424/Y 0.01fF
C22248 AND2X1_LOC_576/a_8_24# OR2X1_LOC_71/Y 0.01fF
C22249 OR2X1_LOC_839/a_8_216# OR2X1_LOC_375/A 0.07fF
C22250 AND2X1_LOC_388/a_8_24# OR2X1_LOC_167/Y 0.03fF
C22251 OR2X1_LOC_532/B OR2X1_LOC_553/A 0.07fF
C22252 OR2X1_LOC_26/Y OR2X1_LOC_246/A 0.12fF
C22253 OR2X1_LOC_95/Y AND2X1_LOC_436/B 0.02fF
C22254 AND2X1_LOC_685/a_36_24# OR2X1_LOC_52/B 0.01fF
C22255 OR2X1_LOC_62/B AND2X1_LOC_852/Y 0.03fF
C22256 AND2X1_LOC_56/a_36_24# AND2X1_LOC_43/B 0.01fF
C22257 OR2X1_LOC_87/A D_INPUT_0 0.10fF
C22258 OR2X1_LOC_278/A OR2X1_LOC_609/A 0.07fF
C22259 AND2X1_LOC_390/a_36_24# OR2X1_LOC_534/Y 0.00fF
C22260 OR2X1_LOC_649/B OR2X1_LOC_655/A 0.03fF
C22261 AND2X1_LOC_41/A OR2X1_LOC_598/A 0.78fF
C22262 OR2X1_LOC_481/a_8_216# AND2X1_LOC_663/B 0.01fF
C22263 OR2X1_LOC_22/Y OR2X1_LOC_585/A 0.40fF
C22264 AND2X1_LOC_91/B OR2X1_LOC_714/a_36_216# 0.00fF
C22265 OR2X1_LOC_380/Y OR2X1_LOC_588/a_8_216# 0.01fF
C22266 OR2X1_LOC_78/B OR2X1_LOC_854/A 0.21fF
C22267 OR2X1_LOC_405/A OR2X1_LOC_786/Y 0.10fF
C22268 OR2X1_LOC_814/A OR2X1_LOC_68/a_36_216# 0.01fF
C22269 AND2X1_LOC_717/B AND2X1_LOC_465/Y 0.03fF
C22270 OR2X1_LOC_246/A OR2X1_LOC_89/A 0.55fF
C22271 OR2X1_LOC_851/B OR2X1_LOC_777/B 0.31fF
C22272 AND2X1_LOC_560/B OR2X1_LOC_256/A 0.01fF
C22273 OR2X1_LOC_421/A OR2X1_LOC_589/a_8_216# 0.01fF
C22274 OR2X1_LOC_631/B AND2X1_LOC_47/Y 0.03fF
C22275 OR2X1_LOC_3/Y AND2X1_LOC_687/B 0.08fF
C22276 OR2X1_LOC_497/a_36_216# AND2X1_LOC_227/Y 0.00fF
C22277 AND2X1_LOC_638/Y OR2X1_LOC_70/A 0.01fF
C22278 OR2X1_LOC_696/A OR2X1_LOC_312/a_8_216# 0.04fF
C22279 OR2X1_LOC_251/Y OR2X1_LOC_417/A 0.06fF
C22280 OR2X1_LOC_748/A AND2X1_LOC_866/A 0.03fF
C22281 AND2X1_LOC_401/a_8_24# OR2X1_LOC_598/A 0.01fF
C22282 AND2X1_LOC_620/Y OR2X1_LOC_39/A 0.03fF
C22283 OR2X1_LOC_26/Y OR2X1_LOC_409/B 0.02fF
C22284 OR2X1_LOC_140/B OR2X1_LOC_563/A 0.01fF
C22285 OR2X1_LOC_43/A AND2X1_LOC_139/A 0.05fF
C22286 OR2X1_LOC_8/Y OR2X1_LOC_437/A 0.01fF
C22287 AND2X1_LOC_483/Y AND2X1_LOC_621/Y 0.05fF
C22288 AND2X1_LOC_91/B OR2X1_LOC_121/A 0.05fF
C22289 OR2X1_LOC_797/B OR2X1_LOC_209/A 0.14fF
C22290 OR2X1_LOC_62/A OR2X1_LOC_753/A 0.20fF
C22291 OR2X1_LOC_151/A OR2X1_LOC_703/Y 0.02fF
C22292 VDD AND2X1_LOC_247/a_8_24# 0.00fF
C22293 OR2X1_LOC_66/A OR2X1_LOC_349/B 0.01fF
C22294 OR2X1_LOC_529/Y OR2X1_LOC_95/Y 0.03fF
C22295 AND2X1_LOC_715/Y OR2X1_LOC_312/a_8_216# 0.02fF
C22296 OR2X1_LOC_756/B OR2X1_LOC_365/a_36_216# 0.00fF
C22297 AND2X1_LOC_44/Y AND2X1_LOC_258/a_8_24# 0.03fF
C22298 OR2X1_LOC_39/A AND2X1_LOC_215/A 0.44fF
C22299 AND2X1_LOC_359/a_36_24# OR2X1_LOC_47/Y 0.00fF
C22300 OR2X1_LOC_715/A OR2X1_LOC_515/Y 0.02fF
C22301 OR2X1_LOC_750/A OR2X1_LOC_750/a_8_216# 0.02fF
C22302 AND2X1_LOC_810/A AND2X1_LOC_539/Y 0.03fF
C22303 OR2X1_LOC_375/A OR2X1_LOC_318/B 0.03fF
C22304 OR2X1_LOC_185/A OR2X1_LOC_641/B 0.02fF
C22305 OR2X1_LOC_234/a_36_216# OR2X1_LOC_753/A 0.00fF
C22306 AND2X1_LOC_79/a_8_24# OR2X1_LOC_404/A 0.09fF
C22307 OR2X1_LOC_45/B AND2X1_LOC_707/Y 0.79fF
C22308 AND2X1_LOC_573/A OR2X1_LOC_88/a_36_216# 0.01fF
C22309 OR2X1_LOC_64/Y OR2X1_LOC_256/A 0.03fF
C22310 OR2X1_LOC_323/A AND2X1_LOC_476/Y 0.18fF
C22311 AND2X1_LOC_227/Y AND2X1_LOC_523/Y 0.26fF
C22312 OR2X1_LOC_243/B OR2X1_LOC_62/B 0.01fF
C22313 AND2X1_LOC_44/Y OR2X1_LOC_708/a_8_216# 0.01fF
C22314 OR2X1_LOC_631/B OR2X1_LOC_598/A 0.02fF
C22315 OR2X1_LOC_19/B AND2X1_LOC_821/a_8_24# 0.04fF
C22316 OR2X1_LOC_263/a_8_216# D_INPUT_0 0.06fF
C22317 AND2X1_LOC_3/Y AND2X1_LOC_418/a_8_24# 0.02fF
C22318 AND2X1_LOC_362/B OR2X1_LOC_89/Y 0.01fF
C22319 AND2X1_LOC_43/B OR2X1_LOC_68/B 6.42fF
C22320 OR2X1_LOC_648/a_8_216# D_INPUT_0 0.01fF
C22321 OR2X1_LOC_585/A OR2X1_LOC_387/a_8_216# 0.06fF
C22322 AND2X1_LOC_712/a_36_24# OR2X1_LOC_12/Y 0.00fF
C22323 OR2X1_LOC_158/A AND2X1_LOC_476/a_8_24# 0.04fF
C22324 OR2X1_LOC_158/A AND2X1_LOC_284/a_36_24# 0.01fF
C22325 OR2X1_LOC_688/a_8_216# OR2X1_LOC_598/A 0.05fF
C22326 AND2X1_LOC_56/B AND2X1_LOC_31/Y 0.11fF
C22327 OR2X1_LOC_109/Y OR2X1_LOC_164/a_8_216# 0.06fF
C22328 AND2X1_LOC_705/Y OR2X1_LOC_12/Y 0.22fF
C22329 AND2X1_LOC_641/Y AND2X1_LOC_641/a_8_24# 0.01fF
C22330 AND2X1_LOC_573/Y AND2X1_LOC_658/B 0.01fF
C22331 AND2X1_LOC_731/a_8_24# AND2X1_LOC_731/Y 0.02fF
C22332 AND2X1_LOC_544/Y VDD 0.38fF
C22333 AND2X1_LOC_721/Y OR2X1_LOC_40/Y 0.02fF
C22334 AND2X1_LOC_48/A OR2X1_LOC_200/Y 0.01fF
C22335 OR2X1_LOC_262/Y OR2X1_LOC_72/Y 0.78fF
C22336 OR2X1_LOC_637/A AND2X1_LOC_36/Y 0.01fF
C22337 AND2X1_LOC_539/Y AND2X1_LOC_567/a_36_24# 0.01fF
C22338 AND2X1_LOC_84/Y AND2X1_LOC_61/Y 0.09fF
C22339 AND2X1_LOC_564/A AND2X1_LOC_731/Y 0.03fF
C22340 OR2X1_LOC_222/A AND2X1_LOC_406/a_8_24# 0.09fF
C22341 OR2X1_LOC_481/A AND2X1_LOC_259/a_8_24# 0.01fF
C22342 VDD AND2X1_LOC_7/B 1.25fF
C22343 OR2X1_LOC_829/a_36_216# OR2X1_LOC_13/B 0.01fF
C22344 OR2X1_LOC_605/B OR2X1_LOC_318/B 0.29fF
C22345 OR2X1_LOC_64/Y OR2X1_LOC_67/Y 0.07fF
C22346 OR2X1_LOC_790/B AND2X1_LOC_41/Y 0.01fF
C22347 AND2X1_LOC_18/Y AND2X1_LOC_44/Y 0.51fF
C22348 AND2X1_LOC_21/Y AND2X1_LOC_31/Y 0.19fF
C22349 OR2X1_LOC_161/A OR2X1_LOC_788/B 0.05fF
C22350 OR2X1_LOC_160/A OR2X1_LOC_777/B 0.07fF
C22351 OR2X1_LOC_97/A OR2X1_LOC_66/A 0.02fF
C22352 AND2X1_LOC_392/A AND2X1_LOC_786/Y 0.07fF
C22353 OR2X1_LOC_97/A OR2X1_LOC_841/A 0.03fF
C22354 OR2X1_LOC_151/A OR2X1_LOC_596/A 0.13fF
C22355 OR2X1_LOC_121/B OR2X1_LOC_544/a_36_216# 0.02fF
C22356 AND2X1_LOC_533/a_8_24# OR2X1_LOC_532/Y 0.00fF
C22357 OR2X1_LOC_224/Y OR2X1_LOC_226/Y 0.04fF
C22358 OR2X1_LOC_62/B AND2X1_LOC_647/B 0.00fF
C22359 AND2X1_LOC_555/Y OR2X1_LOC_698/Y 0.08fF
C22360 AND2X1_LOC_729/B OR2X1_LOC_761/a_36_216# 0.00fF
C22361 OR2X1_LOC_842/A OR2X1_LOC_580/B 0.22fF
C22362 AND2X1_LOC_663/A GATE_579 0.38fF
C22363 OR2X1_LOC_36/Y OR2X1_LOC_300/Y 0.28fF
C22364 OR2X1_LOC_40/Y OR2X1_LOC_482/Y 0.12fF
C22365 AND2X1_LOC_632/A AND2X1_LOC_624/B 0.01fF
C22366 OR2X1_LOC_744/A AND2X1_LOC_244/A 0.03fF
C22367 AND2X1_LOC_476/A AND2X1_LOC_660/A 0.14fF
C22368 AND2X1_LOC_361/A OR2X1_LOC_13/B 0.07fF
C22369 OR2X1_LOC_52/B OR2X1_LOC_437/A 0.03fF
C22370 OR2X1_LOC_417/A AND2X1_LOC_624/B 0.76fF
C22371 AND2X1_LOC_2/Y AND2X1_LOC_40/a_8_24# 0.06fF
C22372 AND2X1_LOC_40/Y OR2X1_LOC_174/a_8_216# 0.01fF
C22373 OR2X1_LOC_744/A OR2X1_LOC_16/A 0.89fF
C22374 AND2X1_LOC_110/Y AND2X1_LOC_299/a_8_24# 0.01fF
C22375 AND2X1_LOC_191/Y AND2X1_LOC_740/a_8_24# 0.04fF
C22376 AND2X1_LOC_65/A OR2X1_LOC_78/A 0.63fF
C22377 VDD OR2X1_LOC_621/a_8_216# 0.21fF
C22378 AND2X1_LOC_91/B AND2X1_LOC_305/a_8_24# 0.05fF
C22379 OR2X1_LOC_501/B OR2X1_LOC_549/A 0.00fF
C22380 AND2X1_LOC_785/a_8_24# OR2X1_LOC_18/Y 0.02fF
C22381 OR2X1_LOC_110/a_8_216# OR2X1_LOC_316/Y 0.00fF
C22382 OR2X1_LOC_759/A OR2X1_LOC_815/a_36_216# 0.00fF
C22383 D_GATE_579 OR2X1_LOC_286/B 0.00fF
C22384 OR2X1_LOC_778/Y AND2X1_LOC_36/Y 0.05fF
C22385 OR2X1_LOC_604/A OR2X1_LOC_816/a_8_216# 0.03fF
C22386 OR2X1_LOC_510/A OR2X1_LOC_78/A 0.01fF
C22387 OR2X1_LOC_291/Y OR2X1_LOC_71/A 0.02fF
C22388 OR2X1_LOC_40/Y OR2X1_LOC_816/Y 0.00fF
C22389 AND2X1_LOC_658/B AND2X1_LOC_806/a_36_24# 0.00fF
C22390 OR2X1_LOC_121/Y OR2X1_LOC_721/Y 0.10fF
C22391 OR2X1_LOC_680/Y OR2X1_LOC_142/Y 0.02fF
C22392 OR2X1_LOC_108/Y OR2X1_LOC_744/A 1.15fF
C22393 AND2X1_LOC_738/B AND2X1_LOC_658/B 0.07fF
C22394 OR2X1_LOC_156/Y OR2X1_LOC_160/A 0.15fF
C22395 AND2X1_LOC_594/a_8_24# AND2X1_LOC_40/Y 0.01fF
C22396 AND2X1_LOC_12/Y OR2X1_LOC_862/a_8_216# 0.01fF
C22397 AND2X1_LOC_306/a_36_24# OR2X1_LOC_307/A 0.00fF
C22398 AND2X1_LOC_658/B OR2X1_LOC_56/A 0.64fF
C22399 OR2X1_LOC_696/A OR2X1_LOC_670/Y 0.01fF
C22400 AND2X1_LOC_22/Y OR2X1_LOC_161/A 0.94fF
C22401 AND2X1_LOC_51/Y OR2X1_LOC_788/B 0.02fF
C22402 OR2X1_LOC_647/A AND2X1_LOC_36/Y 0.03fF
C22403 OR2X1_LOC_160/B OR2X1_LOC_624/Y 0.04fF
C22404 OR2X1_LOC_528/Y AND2X1_LOC_734/Y 0.01fF
C22405 AND2X1_LOC_285/Y OR2X1_LOC_59/Y 0.00fF
C22406 VDD OR2X1_LOC_232/Y 0.12fF
C22407 AND2X1_LOC_396/a_8_24# OR2X1_LOC_78/B 0.01fF
C22408 OR2X1_LOC_147/B OR2X1_LOC_549/A 0.07fF
C22409 OR2X1_LOC_426/A OR2X1_LOC_765/a_8_216# 0.01fF
C22410 OR2X1_LOC_324/a_8_216# OR2X1_LOC_151/A 0.06fF
C22411 AND2X1_LOC_565/B OR2X1_LOC_524/Y 0.01fF
C22412 AND2X1_LOC_543/Y OR2X1_LOC_44/Y 0.04fF
C22413 AND2X1_LOC_482/a_8_24# OR2X1_LOC_736/Y 0.03fF
C22414 OR2X1_LOC_113/Y OR2X1_LOC_244/Y 0.02fF
C22415 OR2X1_LOC_858/A AND2X1_LOC_92/Y 0.02fF
C22416 OR2X1_LOC_241/B OR2X1_LOC_493/Y 0.10fF
C22417 AND2X1_LOC_172/a_36_24# OR2X1_LOC_78/B 0.01fF
C22418 OR2X1_LOC_499/a_8_216# OR2X1_LOC_161/B 0.02fF
C22419 OR2X1_LOC_500/A AND2X1_LOC_44/Y 0.02fF
C22420 OR2X1_LOC_379/Y OR2X1_LOC_856/A 0.73fF
C22421 AND2X1_LOC_716/Y AND2X1_LOC_182/a_36_24# 0.01fF
C22422 OR2X1_LOC_756/B AND2X1_LOC_616/a_8_24# 0.03fF
C22423 OR2X1_LOC_518/a_8_216# OR2X1_LOC_74/A 0.03fF
C22424 AND2X1_LOC_84/Y AND2X1_LOC_852/Y 0.03fF
C22425 AND2X1_LOC_374/a_36_24# AND2X1_LOC_476/Y 0.00fF
C22426 AND2X1_LOC_340/Y OR2X1_LOC_39/A 0.08fF
C22427 AND2X1_LOC_22/Y AND2X1_LOC_25/Y 0.00fF
C22428 AND2X1_LOC_725/a_8_24# OR2X1_LOC_92/Y 0.02fF
C22429 OR2X1_LOC_319/B VDD 0.82fF
C22430 OR2X1_LOC_709/A OR2X1_LOC_793/a_8_216# 0.01fF
C22431 AND2X1_LOC_319/A OR2X1_LOC_428/A 0.04fF
C22432 OR2X1_LOC_427/A AND2X1_LOC_477/Y 0.07fF
C22433 OR2X1_LOC_154/A OR2X1_LOC_61/A 0.04fF
C22434 OR2X1_LOC_61/a_8_216# AND2X1_LOC_18/Y 0.01fF
C22435 OR2X1_LOC_698/a_8_216# OR2X1_LOC_816/Y 0.57fF
C22436 OR2X1_LOC_538/A OR2X1_LOC_78/B 0.03fF
C22437 OR2X1_LOC_135/Y AND2X1_LOC_655/A 0.17fF
C22438 OR2X1_LOC_40/Y OR2X1_LOC_586/Y 0.07fF
C22439 AND2X1_LOC_364/Y OR2X1_LOC_91/A 0.08fF
C22440 OR2X1_LOC_457/B OR2X1_LOC_161/B 0.03fF
C22441 OR2X1_LOC_511/Y OR2X1_LOC_12/Y 0.07fF
C22442 OR2X1_LOC_146/a_8_216# OR2X1_LOC_89/A 0.01fF
C22443 OR2X1_LOC_121/Y OR2X1_LOC_375/A 0.27fF
C22444 OR2X1_LOC_62/B OR2X1_LOC_771/B 0.03fF
C22445 OR2X1_LOC_730/a_8_216# OR2X1_LOC_730/A 0.39fF
C22446 AND2X1_LOC_59/Y AND2X1_LOC_534/a_36_24# 0.01fF
C22447 OR2X1_LOC_154/A OR2X1_LOC_659/Y 0.09fF
C22448 OR2X1_LOC_305/a_8_216# AND2X1_LOC_774/A 0.06fF
C22449 AND2X1_LOC_784/A OR2X1_LOC_310/a_36_216# 0.01fF
C22450 OR2X1_LOC_318/Y VDD 0.15fF
C22451 AND2X1_LOC_181/Y OR2X1_LOC_39/A 0.07fF
C22452 OR2X1_LOC_468/Y OR2X1_LOC_161/B 0.03fF
C22453 OR2X1_LOC_87/A AND2X1_LOC_438/a_8_24# 0.06fF
C22454 AND2X1_LOC_661/A AND2X1_LOC_802/Y 0.03fF
C22455 AND2X1_LOC_650/a_8_24# OR2X1_LOC_171/Y 0.01fF
C22456 VDD OR2X1_LOC_212/a_8_216# 0.00fF
C22457 AND2X1_LOC_554/a_8_24# OR2X1_LOC_89/A 0.01fF
C22458 OR2X1_LOC_248/a_8_216# OR2X1_LOC_12/Y 0.02fF
C22459 AND2X1_LOC_564/B OR2X1_LOC_280/Y 1.43fF
C22460 AND2X1_LOC_721/Y OR2X1_LOC_7/A 0.02fF
C22461 AND2X1_LOC_76/Y AND2X1_LOC_715/A 0.45fF
C22462 AND2X1_LOC_70/Y OR2X1_LOC_856/B 0.08fF
C22463 AND2X1_LOC_290/a_8_24# OR2X1_LOC_66/A 0.14fF
C22464 OR2X1_LOC_65/B AND2X1_LOC_606/a_8_24# 0.23fF
C22465 AND2X1_LOC_706/a_8_24# OR2X1_LOC_44/Y 0.01fF
C22466 VDD AND2X1_LOC_161/a_8_24# -0.00fF
C22467 AND2X1_LOC_95/a_8_24# AND2X1_LOC_59/a_8_24# 0.23fF
C22468 VDD AND2X1_LOC_550/A 0.16fF
C22469 OR2X1_LOC_502/A AND2X1_LOC_306/a_8_24# 0.05fF
C22470 OR2X1_LOC_589/A AND2X1_LOC_831/a_8_24# 0.17fF
C22471 OR2X1_LOC_158/A OR2X1_LOC_236/a_8_216# 0.01fF
C22472 OR2X1_LOC_168/a_36_216# OR2X1_LOC_468/A 0.00fF
C22473 AND2X1_LOC_549/Y AND2X1_LOC_624/A 0.11fF
C22474 OR2X1_LOC_805/A OR2X1_LOC_723/a_36_216# 0.01fF
C22475 OR2X1_LOC_589/A OR2X1_LOC_44/Y 0.01fF
C22476 OR2X1_LOC_474/Y OR2X1_LOC_659/A 0.11fF
C22477 OR2X1_LOC_617/Y AND2X1_LOC_580/a_8_24# 0.01fF
C22478 AND2X1_LOC_294/a_8_24# OR2X1_LOC_12/Y 0.04fF
C22479 OR2X1_LOC_44/Y OR2X1_LOC_322/Y 0.08fF
C22480 OR2X1_LOC_281/a_36_216# OR2X1_LOC_59/Y 0.02fF
C22481 OR2X1_LOC_436/Y OR2X1_LOC_174/Y 0.02fF
C22482 VDD OR2X1_LOC_805/A 1.20fF
C22483 OR2X1_LOC_329/B OR2X1_LOC_427/A 0.09fF
C22484 OR2X1_LOC_440/A OR2X1_LOC_374/a_8_216# 0.39fF
C22485 OR2X1_LOC_759/A OR2X1_LOC_680/A 0.03fF
C22486 AND2X1_LOC_81/B OR2X1_LOC_507/A 0.01fF
C22487 AND2X1_LOC_719/Y OR2X1_LOC_283/Y 0.10fF
C22488 OR2X1_LOC_843/a_8_216# OR2X1_LOC_843/B 0.02fF
C22489 AND2X1_LOC_500/Y AND2X1_LOC_624/A 0.12fF
C22490 AND2X1_LOC_849/A AND2X1_LOC_227/a_8_24# 0.20fF
C22491 AND2X1_LOC_542/a_8_24# OR2X1_LOC_312/Y 0.01fF
C22492 OR2X1_LOC_181/B D_GATE_741 0.03fF
C22493 AND2X1_LOC_47/Y INPUT_6 0.03fF
C22494 OR2X1_LOC_51/Y AND2X1_LOC_470/B 0.01fF
C22495 OR2X1_LOC_604/A OR2X1_LOC_699/a_8_216# 0.06fF
C22496 OR2X1_LOC_158/A OR2X1_LOC_32/a_8_216# 0.03fF
C22497 OR2X1_LOC_100/a_8_216# OR2X1_LOC_78/B 0.02fF
C22498 AND2X1_LOC_181/Y AND2X1_LOC_211/B 0.03fF
C22499 OR2X1_LOC_40/Y OR2X1_LOC_748/A 0.02fF
C22500 AND2X1_LOC_22/Y AND2X1_LOC_51/Y 0.81fF
C22501 OR2X1_LOC_532/B OR2X1_LOC_354/a_8_216# 0.01fF
C22502 OR2X1_LOC_333/B OR2X1_LOC_390/A 0.09fF
C22503 OR2X1_LOC_822/Y OR2X1_LOC_85/A 0.01fF
C22504 AND2X1_LOC_124/a_8_24# OR2X1_LOC_56/A 0.02fF
C22505 AND2X1_LOC_12/Y OR2X1_LOC_78/B 1.80fF
C22506 AND2X1_LOC_474/A OR2X1_LOC_18/Y 0.06fF
C22507 OR2X1_LOC_169/B AND2X1_LOC_92/Y 0.09fF
C22508 OR2X1_LOC_482/Y OR2X1_LOC_7/A 0.06fF
C22509 AND2X1_LOC_140/a_8_24# OR2X1_LOC_595/A -0.03fF
C22510 AND2X1_LOC_162/a_36_24# OR2X1_LOC_619/Y 0.00fF
C22511 OR2X1_LOC_832/a_8_216# OR2X1_LOC_449/B 0.07fF
C22512 AND2X1_LOC_41/A OR2X1_LOC_506/A 0.31fF
C22513 OR2X1_LOC_261/a_8_216# OR2X1_LOC_44/Y 0.01fF
C22514 AND2X1_LOC_40/Y OR2X1_LOC_792/Y 0.51fF
C22515 AND2X1_LOC_658/A OR2X1_LOC_36/Y 0.03fF
C22516 OR2X1_LOC_91/Y OR2X1_LOC_59/Y 0.16fF
C22517 AND2X1_LOC_550/A OR2X1_LOC_677/Y 0.01fF
C22518 OR2X1_LOC_444/B AND2X1_LOC_7/B 0.13fF
C22519 VDD AND2X1_LOC_101/B 0.01fF
C22520 OR2X1_LOC_78/B OR2X1_LOC_802/A 0.01fF
C22521 OR2X1_LOC_8/Y OR2X1_LOC_753/A 0.23fF
C22522 AND2X1_LOC_561/a_36_24# AND2X1_LOC_866/A 0.01fF
C22523 OR2X1_LOC_533/a_8_216# OR2X1_LOC_331/Y 0.05fF
C22524 OR2X1_LOC_625/a_36_216# OR2X1_LOC_92/Y 0.02fF
C22525 AND2X1_LOC_715/A OR2X1_LOC_52/B 0.00fF
C22526 OR2X1_LOC_633/Y OR2X1_LOC_640/A 0.15fF
C22527 OR2X1_LOC_536/Y OR2X1_LOC_385/Y 0.10fF
C22528 OR2X1_LOC_166/Y OR2X1_LOC_44/Y 0.03fF
C22529 AND2X1_LOC_117/a_8_24# AND2X1_LOC_262/a_8_24# 0.23fF
C22530 OR2X1_LOC_62/B OR2X1_LOC_572/a_36_216# 0.00fF
C22531 AND2X1_LOC_792/Y AND2X1_LOC_789/Y 0.07fF
C22532 OR2X1_LOC_756/B AND2X1_LOC_251/a_8_24# 0.02fF
C22533 OR2X1_LOC_176/a_36_216# AND2X1_LOC_477/A 0.02fF
C22534 OR2X1_LOC_676/Y AND2X1_LOC_3/Y 0.09fF
C22535 AND2X1_LOC_713/a_8_24# OR2X1_LOC_64/Y 0.01fF
C22536 AND2X1_LOC_566/Y OR2X1_LOC_600/A 0.33fF
C22537 OR2X1_LOC_297/A OR2X1_LOC_44/Y 0.00fF
C22538 OR2X1_LOC_466/A OR2X1_LOC_453/A 0.01fF
C22539 OR2X1_LOC_467/B AND2X1_LOC_51/Y 0.18fF
C22540 AND2X1_LOC_537/Y AND2X1_LOC_774/A 0.17fF
C22541 OR2X1_LOC_335/Y OR2X1_LOC_87/A 0.00fF
C22542 OR2X1_LOC_650/a_36_216# AND2X1_LOC_8/Y 0.00fF
C22543 AND2X1_LOC_134/a_8_24# OR2X1_LOC_161/B 0.11fF
C22544 OR2X1_LOC_411/Y OR2X1_LOC_52/B 0.03fF
C22545 OR2X1_LOC_804/A OR2X1_LOC_593/B 0.00fF
C22546 AND2X1_LOC_541/a_8_24# OR2X1_LOC_256/A 0.09fF
C22547 D_INPUT_5 OR2X1_LOC_375/A 0.06fF
C22548 AND2X1_LOC_112/a_8_24# OR2X1_LOC_74/A 0.05fF
C22549 AND2X1_LOC_59/Y AND2X1_LOC_58/a_8_24# 0.01fF
C22550 VDD OR2X1_LOC_296/Y 0.31fF
C22551 OR2X1_LOC_68/B OR2X1_LOC_558/A 0.00fF
C22552 OR2X1_LOC_588/Y OR2X1_LOC_26/a_8_216# 0.00fF
C22553 OR2X1_LOC_160/A OR2X1_LOC_575/A 0.27fF
C22554 OR2X1_LOC_40/Y OR2X1_LOC_304/Y 0.13fF
C22555 OR2X1_LOC_92/Y AND2X1_LOC_435/a_36_24# 0.06fF
C22556 OR2X1_LOC_471/Y OR2X1_LOC_161/B 0.04fF
C22557 OR2X1_LOC_49/A INPUT_1 0.14fF
C22558 OR2X1_LOC_703/B AND2X1_LOC_40/Y 0.02fF
C22559 AND2X1_LOC_565/B AND2X1_LOC_578/A 0.01fF
C22560 OR2X1_LOC_160/A OR2X1_LOC_660/a_36_216# 0.00fF
C22561 OR2X1_LOC_849/A OR2X1_LOC_624/a_8_216# 0.01fF
C22562 AND2X1_LOC_593/Y OR2X1_LOC_48/B 0.02fF
C22563 OR2X1_LOC_834/A AND2X1_LOC_3/Y 0.42fF
C22564 OR2X1_LOC_175/Y OR2X1_LOC_468/a_8_216# 0.05fF
C22565 AND2X1_LOC_113/Y OR2X1_LOC_427/A 0.01fF
C22566 OR2X1_LOC_160/A OR2X1_LOC_493/A 0.11fF
C22567 OR2X1_LOC_256/Y AND2X1_LOC_359/B 1.00fF
C22568 OR2X1_LOC_59/Y OR2X1_LOC_757/Y 0.01fF
C22569 AND2X1_LOC_40/Y OR2X1_LOC_87/A 0.59fF
C22570 OR2X1_LOC_612/B AND2X1_LOC_647/a_8_24# 0.01fF
C22571 OR2X1_LOC_185/A OR2X1_LOC_739/A 0.03fF
C22572 AND2X1_LOC_721/Y OR2X1_LOC_224/a_8_216# 0.14fF
C22573 OR2X1_LOC_85/A AND2X1_LOC_852/B 0.03fF
C22574 AND2X1_LOC_654/B OR2X1_LOC_44/Y 0.01fF
C22575 OR2X1_LOC_691/B OR2X1_LOC_532/B 0.00fF
C22576 OR2X1_LOC_2/Y OR2X1_LOC_25/a_8_216# 0.02fF
C22577 AND2X1_LOC_148/a_8_24# OR2X1_LOC_74/A 0.05fF
C22578 OR2X1_LOC_653/Y OR2X1_LOC_358/B 0.00fF
C22579 OR2X1_LOC_31/Y OR2X1_LOC_16/A 0.13fF
C22580 AND2X1_LOC_374/a_8_24# OR2X1_LOC_26/Y 0.05fF
C22581 AND2X1_LOC_59/Y OR2X1_LOC_377/A 0.11fF
C22582 AND2X1_LOC_580/A OR2X1_LOC_531/a_8_216# 0.00fF
C22583 OR2X1_LOC_40/Y OR2X1_LOC_628/Y 0.07fF
C22584 OR2X1_LOC_160/A OR2X1_LOC_652/a_8_216# 0.04fF
C22585 AND2X1_LOC_166/a_8_24# OR2X1_LOC_169/B 0.01fF
C22586 OR2X1_LOC_804/A AND2X1_LOC_273/a_8_24# 0.01fF
C22587 AND2X1_LOC_12/Y OR2X1_LOC_375/A 2.53fF
C22588 OR2X1_LOC_527/Y OR2X1_LOC_59/Y 0.07fF
C22589 AND2X1_LOC_852/Y OR2X1_LOC_393/a_8_216# 0.06fF
C22590 OR2X1_LOC_179/Y OR2X1_LOC_529/Y 0.01fF
C22591 OR2X1_LOC_18/Y OR2X1_LOC_85/A 0.37fF
C22592 AND2X1_LOC_524/a_8_24# AND2X1_LOC_47/Y 0.01fF
C22593 OR2X1_LOC_291/a_36_216# OR2X1_LOC_36/Y 0.03fF
C22594 OR2X1_LOC_837/a_8_216# OR2X1_LOC_753/A 0.37fF
C22595 AND2X1_LOC_91/B AND2X1_LOC_72/B 0.03fF
C22596 OR2X1_LOC_525/Y OR2X1_LOC_26/Y 0.27fF
C22597 OR2X1_LOC_207/B OR2X1_LOC_200/Y 0.07fF
C22598 OR2X1_LOC_461/a_8_216# OR2X1_LOC_19/B 0.14fF
C22599 OR2X1_LOC_74/A OR2X1_LOC_746/a_8_216# 0.02fF
C22600 OR2X1_LOC_291/Y OR2X1_LOC_59/Y 0.26fF
C22601 OR2X1_LOC_720/B AND2X1_LOC_18/Y 0.03fF
C22602 OR2X1_LOC_244/B AND2X1_LOC_51/Y 0.01fF
C22603 OR2X1_LOC_671/Y OR2X1_LOC_96/a_8_216# 0.01fF
C22604 OR2X1_LOC_672/a_8_216# OR2X1_LOC_95/Y 0.01fF
C22605 OR2X1_LOC_185/A OR2X1_LOC_269/B 0.08fF
C22606 AND2X1_LOC_621/Y AND2X1_LOC_806/A 0.03fF
C22607 OR2X1_LOC_484/a_8_216# AND2X1_LOC_727/A 0.01fF
C22608 OR2X1_LOC_456/Y OR2X1_LOC_465/a_8_216# 0.18fF
C22609 OR2X1_LOC_756/B OR2X1_LOC_285/B 0.01fF
C22610 OR2X1_LOC_389/A D_INPUT_0 0.01fF
C22611 AND2X1_LOC_721/A OR2X1_LOC_428/A 0.04fF
C22612 OR2X1_LOC_525/Y OR2X1_LOC_89/A 0.03fF
C22613 OR2X1_LOC_569/B OR2X1_LOC_565/a_8_216# 0.14fF
C22614 OR2X1_LOC_642/a_8_216# OR2X1_LOC_130/A 0.14fF
C22615 OR2X1_LOC_87/A OR2X1_LOC_87/Y 0.03fF
C22616 OR2X1_LOC_108/Y OR2X1_LOC_31/Y 0.14fF
C22617 OR2X1_LOC_485/A OR2X1_LOC_278/Y 0.06fF
C22618 AND2X1_LOC_379/a_8_24# OR2X1_LOC_44/Y 0.01fF
C22619 OR2X1_LOC_679/A AND2X1_LOC_657/Y 0.03fF
C22620 AND2X1_LOC_95/Y OR2X1_LOC_787/Y 0.07fF
C22621 OR2X1_LOC_634/A OR2X1_LOC_19/B 0.03fF
C22622 OR2X1_LOC_744/A AND2X1_LOC_687/Y 0.02fF
C22623 AND2X1_LOC_485/a_8_24# AND2X1_LOC_44/Y 0.04fF
C22624 OR2X1_LOC_585/A OR2X1_LOC_39/A 0.10fF
C22625 AND2X1_LOC_566/Y OR2X1_LOC_619/Y 0.04fF
C22626 AND2X1_LOC_597/a_8_24# AND2X1_LOC_56/B 0.01fF
C22627 OR2X1_LOC_474/Y OR2X1_LOC_121/B 0.11fF
C22628 OR2X1_LOC_673/Y AND2X1_LOC_399/a_8_24# 0.02fF
C22629 AND2X1_LOC_554/B OR2X1_LOC_118/Y 0.61fF
C22630 VDD OR2X1_LOC_55/a_8_216# 0.21fF
C22631 OR2X1_LOC_837/B OR2X1_LOC_27/Y 0.03fF
C22632 OR2X1_LOC_306/a_8_216# OR2X1_LOC_743/A 0.03fF
C22633 AND2X1_LOC_228/Y AND2X1_LOC_211/B 0.01fF
C22634 AND2X1_LOC_486/Y OR2X1_LOC_64/Y 6.10fF
C22635 OR2X1_LOC_43/A OR2X1_LOC_44/Y 0.13fF
C22636 OR2X1_LOC_836/A OR2X1_LOC_836/B 0.07fF
C22637 OR2X1_LOC_648/A AND2X1_LOC_47/Y 0.10fF
C22638 AND2X1_LOC_78/a_36_24# OR2X1_LOC_18/Y 0.01fF
C22639 OR2X1_LOC_175/Y OR2X1_LOC_568/a_8_216# 0.03fF
C22640 OR2X1_LOC_703/Y OR2X1_LOC_714/A 0.06fF
C22641 OR2X1_LOC_280/a_36_216# OR2X1_LOC_237/Y 0.00fF
C22642 AND2X1_LOC_416/a_8_24# OR2X1_LOC_68/B 0.02fF
C22643 AND2X1_LOC_19/a_8_24# OR2X1_LOC_87/Y 0.01fF
C22644 AND2X1_LOC_81/B OR2X1_LOC_646/A 0.01fF
C22645 AND2X1_LOC_191/B AND2X1_LOC_227/Y 0.12fF
C22646 OR2X1_LOC_22/Y AND2X1_LOC_857/Y 0.10fF
C22647 AND2X1_LOC_222/Y OR2X1_LOC_310/a_8_216# 0.01fF
C22648 AND2X1_LOC_495/a_8_24# OR2X1_LOC_203/Y 0.04fF
C22649 AND2X1_LOC_12/Y OR2X1_LOC_605/B 0.18fF
C22650 AND2X1_LOC_502/a_36_24# OR2X1_LOC_485/A 0.00fF
C22651 AND2X1_LOC_565/Y AND2X1_LOC_474/Y 0.03fF
C22652 OR2X1_LOC_158/A AND2X1_LOC_203/Y 0.04fF
C22653 OR2X1_LOC_864/A AND2X1_LOC_8/Y 0.02fF
C22654 AND2X1_LOC_54/a_36_24# D_INPUT_0 0.00fF
C22655 OR2X1_LOC_275/A OR2X1_LOC_595/a_8_216# 0.01fF
C22656 OR2X1_LOC_846/a_8_216# OR2X1_LOC_846/B 0.02fF
C22657 OR2X1_LOC_753/A OR2X1_LOC_52/B 0.72fF
C22658 OR2X1_LOC_838/a_8_216# D_INPUT_0 0.01fF
C22659 OR2X1_LOC_497/Y OR2X1_LOC_89/A 0.63fF
C22660 OR2X1_LOC_299/Y OR2X1_LOC_6/A 0.01fF
C22661 OR2X1_LOC_91/Y OR2X1_LOC_70/Y 0.07fF
C22662 OR2X1_LOC_161/B OR2X1_LOC_750/Y 0.65fF
C22663 AND2X1_LOC_8/Y OR2X1_LOC_633/B 0.08fF
C22664 OR2X1_LOC_47/Y OR2X1_LOC_56/A 0.22fF
C22665 AND2X1_LOC_211/B OR2X1_LOC_585/A 0.03fF
C22666 OR2X1_LOC_19/B OR2X1_LOC_414/a_36_216# 0.01fF
C22667 OR2X1_LOC_140/A OR2X1_LOC_66/Y 0.01fF
C22668 INPUT_0 AND2X1_LOC_660/A 0.03fF
C22669 AND2X1_LOC_10/a_8_24# OR2X1_LOC_204/Y 0.01fF
C22670 OR2X1_LOC_676/Y OR2X1_LOC_194/a_8_216# 0.02fF
C22671 OR2X1_LOC_819/a_8_216# OR2X1_LOC_47/Y 0.00fF
C22672 OR2X1_LOC_475/Y OR2X1_LOC_87/A 0.02fF
C22673 OR2X1_LOC_643/A AND2X1_LOC_122/a_8_24# 0.05fF
C22674 AND2X1_LOC_486/Y OR2X1_LOC_417/A 0.03fF
C22675 AND2X1_LOC_564/a_36_24# AND2X1_LOC_711/Y 0.01fF
C22676 AND2X1_LOC_122/a_8_24# OR2X1_LOC_124/Y 0.01fF
C22677 OR2X1_LOC_595/A AND2X1_LOC_217/a_8_24# 0.00fF
C22678 OR2X1_LOC_479/Y OR2X1_LOC_810/A 0.03fF
C22679 AND2X1_LOC_784/Y AND2X1_LOC_222/Y 0.01fF
C22680 OR2X1_LOC_316/Y OR2X1_LOC_268/a_8_216# 0.01fF
C22681 OR2X1_LOC_70/Y AND2X1_LOC_446/a_8_24# 0.02fF
C22682 OR2X1_LOC_306/Y AND2X1_LOC_856/a_36_24# 0.00fF
C22683 OR2X1_LOC_217/Y OR2X1_LOC_121/B 0.02fF
C22684 OR2X1_LOC_862/B OR2X1_LOC_493/Y 0.28fF
C22685 AND2X1_LOC_658/A OR2X1_LOC_419/Y 0.03fF
C22686 AND2X1_LOC_733/a_36_24# OR2X1_LOC_95/Y 0.01fF
C22687 OR2X1_LOC_269/B OR2X1_LOC_713/a_8_216# 0.01fF
C22688 OR2X1_LOC_52/B OR2X1_LOC_27/a_36_216# 0.02fF
C22689 AND2X1_LOC_191/Y OR2X1_LOC_152/Y 0.03fF
C22690 OR2X1_LOC_189/Y AND2X1_LOC_711/Y 2.18fF
C22691 AND2X1_LOC_41/A D_INPUT_1 0.03fF
C22692 OR2X1_LOC_605/Y OR2X1_LOC_301/a_8_216# 0.03fF
C22693 AND2X1_LOC_476/A AND2X1_LOC_642/Y 0.04fF
C22694 OR2X1_LOC_189/Y OR2X1_LOC_70/Y 0.03fF
C22695 AND2X1_LOC_316/a_8_24# OR2X1_LOC_786/Y 0.14fF
C22696 AND2X1_LOC_711/Y OR2X1_LOC_757/Y 0.01fF
C22697 OR2X1_LOC_152/Y AND2X1_LOC_711/Y 0.00fF
C22698 OR2X1_LOC_687/Y AND2X1_LOC_425/Y 0.01fF
C22699 AND2X1_LOC_845/Y OR2X1_LOC_67/A 0.03fF
C22700 AND2X1_LOC_91/B AND2X1_LOC_36/Y 0.29fF
C22701 AND2X1_LOC_680/a_8_24# OR2X1_LOC_449/B 0.03fF
C22702 OR2X1_LOC_264/Y OR2X1_LOC_340/a_8_216# 0.01fF
C22703 OR2X1_LOC_246/A OR2X1_LOC_246/a_8_216# 0.09fF
C22704 AND2X1_LOC_191/B OR2X1_LOC_753/Y 0.43fF
C22705 AND2X1_LOC_191/Y OR2X1_LOC_527/Y 0.19fF
C22706 AND2X1_LOC_214/A AND2X1_LOC_228/a_8_24# 0.11fF
C22707 AND2X1_LOC_42/B OR2X1_LOC_97/a_8_216# 0.01fF
C22708 OR2X1_LOC_3/Y OR2X1_LOC_681/Y 0.04fF
C22709 AND2X1_LOC_844/a_8_24# OR2X1_LOC_89/A 0.01fF
C22710 OR2X1_LOC_281/Y OR2X1_LOC_437/A 0.08fF
C22711 AND2X1_LOC_31/a_8_24# AND2X1_LOC_21/Y 0.17fF
C22712 AND2X1_LOC_31/Y OR2X1_LOC_787/B 0.29fF
C22713 AND2X1_LOC_711/Y OR2X1_LOC_527/Y 0.08fF
C22714 AND2X1_LOC_866/A AND2X1_LOC_848/a_8_24# 0.02fF
C22715 OR2X1_LOC_779/Y OR2X1_LOC_725/B 0.72fF
C22716 AND2X1_LOC_219/Y AND2X1_LOC_222/Y 0.02fF
C22717 OR2X1_LOC_70/Y OR2X1_LOC_527/Y 0.11fF
C22718 OR2X1_LOC_750/a_36_216# OR2X1_LOC_269/B 0.01fF
C22719 AND2X1_LOC_658/A OR2X1_LOC_152/A 0.03fF
C22720 OR2X1_LOC_61/Y OR2X1_LOC_205/Y 0.01fF
C22721 AND2X1_LOC_31/Y AND2X1_LOC_92/Y 0.10fF
C22722 OR2X1_LOC_485/A OR2X1_LOC_19/B 0.06fF
C22723 OR2X1_LOC_115/a_8_216# OR2X1_LOC_786/Y 0.01fF
C22724 AND2X1_LOC_599/a_36_24# AND2X1_LOC_36/Y 0.00fF
C22725 OR2X1_LOC_756/B OR2X1_LOC_358/A 0.59fF
C22726 OR2X1_LOC_628/Y OR2X1_LOC_7/A 0.24fF
C22727 OR2X1_LOC_333/B OR2X1_LOC_750/A 0.03fF
C22728 OR2X1_LOC_596/A OR2X1_LOC_714/A 0.02fF
C22729 OR2X1_LOC_3/Y OR2X1_LOC_416/Y 0.03fF
C22730 AND2X1_LOC_431/a_8_24# OR2X1_LOC_269/B 0.04fF
C22731 OR2X1_LOC_70/Y OR2X1_LOC_417/Y 0.04fF
C22732 OR2X1_LOC_158/A OR2X1_LOC_424/Y 0.00fF
C22733 AND2X1_LOC_663/A AND2X1_LOC_657/A 0.10fF
C22734 OR2X1_LOC_70/Y OR2X1_LOC_311/Y 0.04fF
C22735 OR2X1_LOC_287/B OR2X1_LOC_286/B 0.00fF
C22736 OR2X1_LOC_485/A AND2X1_LOC_800/a_8_24# 0.00fF
C22737 AND2X1_LOC_476/Y OR2X1_LOC_142/Y 0.07fF
C22738 OR2X1_LOC_354/A OR2X1_LOC_854/A 0.29fF
C22739 AND2X1_LOC_403/a_8_24# OR2X1_LOC_399/Y 0.23fF
C22740 OR2X1_LOC_666/Y OR2X1_LOC_417/A 0.04fF
C22741 OR2X1_LOC_185/Y OR2X1_LOC_473/A 0.11fF
C22742 OR2X1_LOC_158/A D_INPUT_6 0.37fF
C22743 D_INPUT_3 OR2X1_LOC_820/B 0.02fF
C22744 AND2X1_LOC_560/B AND2X1_LOC_660/A 0.06fF
C22745 OR2X1_LOC_417/Y AND2X1_LOC_514/Y 0.23fF
C22746 OR2X1_LOC_439/B OR2X1_LOC_180/B 0.76fF
C22747 AND2X1_LOC_785/A OR2X1_LOC_177/Y 0.01fF
C22748 OR2X1_LOC_760/a_8_216# OR2X1_LOC_585/A 0.01fF
C22749 OR2X1_LOC_91/Y OR2X1_LOC_437/Y 0.40fF
C22750 OR2X1_LOC_375/A OR2X1_LOC_98/a_8_216# 0.03fF
C22751 AND2X1_LOC_514/a_8_24# OR2X1_LOC_437/A 0.04fF
C22752 AND2X1_LOC_95/Y AND2X1_LOC_52/Y 0.03fF
C22753 AND2X1_LOC_192/Y AND2X1_LOC_781/Y 0.05fF
C22754 OR2X1_LOC_631/B D_INPUT_1 0.03fF
C22755 AND2X1_LOC_161/a_8_24# OR2X1_LOC_163/Y 0.00fF
C22756 AND2X1_LOC_170/B AND2X1_LOC_211/a_8_24# 0.01fF
C22757 OR2X1_LOC_311/Y AND2X1_LOC_538/a_8_24# 0.01fF
C22758 AND2X1_LOC_91/B AND2X1_LOC_488/a_8_24# 0.02fF
C22759 OR2X1_LOC_488/Y OR2X1_LOC_71/Y 0.01fF
C22760 AND2X1_LOC_721/Y AND2X1_LOC_284/a_36_24# 0.00fF
C22761 OR2X1_LOC_610/a_8_216# OR2X1_LOC_68/B 0.11fF
C22762 OR2X1_LOC_508/a_8_216# AND2X1_LOC_64/Y -0.00fF
C22763 OR2X1_LOC_497/a_8_216# OR2X1_LOC_419/Y 0.00fF
C22764 OR2X1_LOC_814/A OR2X1_LOC_846/A 0.01fF
C22765 AND2X1_LOC_64/Y OR2X1_LOC_486/Y 0.25fF
C22766 OR2X1_LOC_85/A AND2X1_LOC_215/A -0.01fF
C22767 AND2X1_LOC_538/a_8_24# AND2X1_LOC_538/Y 0.01fF
C22768 AND2X1_LOC_536/a_8_24# OR2X1_LOC_750/Y 0.07fF
C22769 AND2X1_LOC_656/Y AND2X1_LOC_663/B 0.08fF
C22770 AND2X1_LOC_574/A AND2X1_LOC_657/a_8_24# 0.08fF
C22771 OR2X1_LOC_241/Y AND2X1_LOC_67/Y 0.12fF
C22772 AND2X1_LOC_101/B OR2X1_LOC_67/Y 0.01fF
C22773 AND2X1_LOC_231/a_8_24# OR2X1_LOC_12/Y 0.01fF
C22774 OR2X1_LOC_188/Y AND2X1_LOC_255/a_36_24# 0.00fF
C22775 AND2X1_LOC_504/a_36_24# OR2X1_LOC_560/A 0.01fF
C22776 AND2X1_LOC_866/A AND2X1_LOC_523/Y 0.03fF
C22777 OR2X1_LOC_291/A OR2X1_LOC_47/Y 1.93fF
C22778 OR2X1_LOC_736/Y OR2X1_LOC_563/A 0.07fF
C22779 OR2X1_LOC_144/a_8_216# VDD 0.00fF
C22780 AND2X1_LOC_625/a_8_24# OR2X1_LOC_115/B 0.01fF
C22781 OR2X1_LOC_631/A OR2X1_LOC_140/B 0.00fF
C22782 OR2X1_LOC_111/Y OR2X1_LOC_46/A 0.18fF
C22783 OR2X1_LOC_404/A OR2X1_LOC_532/B 0.25fF
C22784 OR2X1_LOC_151/A OR2X1_LOC_392/B 2.89fF
C22785 OR2X1_LOC_185/Y OR2X1_LOC_228/Y 0.07fF
C22786 AND2X1_LOC_774/a_36_24# AND2X1_LOC_774/A 0.01fF
C22787 AND2X1_LOC_707/Y OR2X1_LOC_158/A 0.11fF
C22788 OR2X1_LOC_165/a_8_216# OR2X1_LOC_437/A 0.03fF
C22789 OR2X1_LOC_45/B OR2X1_LOC_589/A 0.19fF
C22790 AND2X1_LOC_687/Y OR2X1_LOC_31/Y 0.01fF
C22791 OR2X1_LOC_411/a_8_216# OR2X1_LOC_46/A 0.01fF
C22792 OR2X1_LOC_78/A OR2X1_LOC_502/a_36_216# 0.03fF
C22793 OR2X1_LOC_78/B OR2X1_LOC_356/B 0.07fF
C22794 AND2X1_LOC_729/B OR2X1_LOC_41/a_8_216# 0.01fF
C22795 OR2X1_LOC_307/A AND2X1_LOC_44/Y 0.01fF
C22796 OR2X1_LOC_71/Y OR2X1_LOC_95/Y 0.31fF
C22797 OR2X1_LOC_19/B OR2X1_LOC_396/a_8_216# 0.03fF
C22798 OR2X1_LOC_121/Y OR2X1_LOC_549/A 0.39fF
C22799 AND2X1_LOC_159/a_8_24# OR2X1_LOC_68/B 0.03fF
C22800 AND2X1_LOC_59/Y OR2X1_LOC_732/A 1.90fF
C22801 OR2X1_LOC_175/Y OR2X1_LOC_66/A 2.43fF
C22802 OR2X1_LOC_19/B OR2X1_LOC_609/Y 0.03fF
C22803 OR2X1_LOC_160/A OR2X1_LOC_735/B 0.03fF
C22804 OR2X1_LOC_193/A OR2X1_LOC_801/B 0.02fF
C22805 OR2X1_LOC_810/A OR2X1_LOC_68/B 0.03fF
C22806 OR2X1_LOC_756/B OR2X1_LOC_168/Y 0.34fF
C22807 OR2X1_LOC_632/Y OR2X1_LOC_140/B 0.09fF
C22808 AND2X1_LOC_856/B OR2X1_LOC_599/Y 0.12fF
C22809 AND2X1_LOC_91/B OR2X1_LOC_630/Y 0.10fF
C22810 OR2X1_LOC_666/A AND2X1_LOC_284/a_8_24# 0.01fF
C22811 AND2X1_LOC_462/B OR2X1_LOC_416/Y 0.17fF
C22812 AND2X1_LOC_654/Y OR2X1_LOC_320/a_36_216# 0.01fF
C22813 OR2X1_LOC_415/a_8_216# OR2X1_LOC_396/Y 0.40fF
C22814 OR2X1_LOC_154/A OR2X1_LOC_515/a_8_216# 0.03fF
C22815 OR2X1_LOC_691/Y OR2X1_LOC_66/A 0.03fF
C22816 OR2X1_LOC_66/A AND2X1_LOC_417/a_8_24# 0.02fF
C22817 OR2X1_LOC_417/A AND2X1_LOC_660/A 0.04fF
C22818 VDD OR2X1_LOC_580/B 0.70fF
C22819 AND2X1_LOC_301/a_8_24# OR2X1_LOC_16/A 0.01fF
C22820 AND2X1_LOC_95/Y OR2X1_LOC_523/a_8_216# 0.01fF
C22821 AND2X1_LOC_72/Y AND2X1_LOC_36/Y 0.03fF
C22822 AND2X1_LOC_214/A OR2X1_LOC_53/Y 0.03fF
C22823 OR2X1_LOC_3/Y OR2X1_LOC_80/A 0.03fF
C22824 OR2X1_LOC_66/A OR2X1_LOC_713/A 0.07fF
C22825 OR2X1_LOC_97/A AND2X1_LOC_164/a_8_24# 0.01fF
C22826 AND2X1_LOC_59/Y OR2X1_LOC_539/B 0.02fF
C22827 AND2X1_LOC_710/a_8_24# AND2X1_LOC_789/Y 0.02fF
C22828 OR2X1_LOC_809/B OR2X1_LOC_161/B 0.02fF
C22829 D_INPUT_3 AND2X1_LOC_14/a_8_24# 0.00fF
C22830 OR2X1_LOC_334/B AND2X1_LOC_7/B 0.04fF
C22831 OR2X1_LOC_177/Y AND2X1_LOC_658/A 0.03fF
C22832 AND2X1_LOC_773/Y OR2X1_LOC_91/A 0.10fF
C22833 OR2X1_LOC_261/a_8_216# OR2X1_LOC_382/A 0.01fF
C22834 OR2X1_LOC_248/a_8_216# OR2X1_LOC_248/A 0.47fF
C22835 OR2X1_LOC_410/Y AND2X1_LOC_411/a_8_24# 0.23fF
C22836 AND2X1_LOC_525/a_36_24# OR2X1_LOC_546/A 0.00fF
C22837 OR2X1_LOC_516/B AND2X1_LOC_794/a_8_24# 0.01fF
C22838 AND2X1_LOC_605/Y OR2X1_LOC_428/A 0.02fF
C22839 OR2X1_LOC_270/a_8_216# AND2X1_LOC_36/Y 0.06fF
C22840 OR2X1_LOC_6/B OR2X1_LOC_612/a_36_216# 0.02fF
C22841 VDD OR2X1_LOC_648/B 0.88fF
C22842 OR2X1_LOC_280/Y OR2X1_LOC_437/A 0.12fF
C22843 AND2X1_LOC_207/A AND2X1_LOC_207/B 0.19fF
C22844 OR2X1_LOC_40/Y AND2X1_LOC_508/B 0.03fF
C22845 VDD OR2X1_LOC_96/Y 0.30fF
C22846 AND2X1_LOC_555/Y OR2X1_LOC_18/Y 0.02fF
C22847 AND2X1_LOC_787/A AND2X1_LOC_716/Y 0.01fF
C22848 AND2X1_LOC_544/Y AND2X1_LOC_811/B 0.00fF
C22849 OR2X1_LOC_411/A OR2X1_LOC_600/A 0.09fF
C22850 OR2X1_LOC_604/A AND2X1_LOC_658/A 0.10fF
C22851 AND2X1_LOC_51/Y OR2X1_LOC_705/a_36_216# 0.00fF
C22852 AND2X1_LOC_91/B OR2X1_LOC_447/a_36_216# 0.02fF
C22853 AND2X1_LOC_455/a_8_24# OR2X1_LOC_39/A -0.01fF
C22854 OR2X1_LOC_91/A AND2X1_LOC_243/Y 0.07fF
C22855 OR2X1_LOC_464/A OR2X1_LOC_486/Y 0.03fF
C22856 OR2X1_LOC_6/B OR2X1_LOC_820/A 0.80fF
C22857 VDD OR2X1_LOC_742/a_8_216# 0.21fF
C22858 OR2X1_LOC_840/a_8_216# AND2X1_LOC_40/Y 0.02fF
C22859 OR2X1_LOC_113/Y OR2X1_LOC_114/B 0.16fF
C22860 OR2X1_LOC_757/A OR2X1_LOC_759/A 2.01fF
C22861 AND2X1_LOC_564/B OR2X1_LOC_39/A 0.10fF
C22862 VDD AND2X1_LOC_103/a_8_24# -0.00fF
C22863 VDD AND2X1_LOC_663/A 5.74fF
C22864 OR2X1_LOC_244/Y OR2X1_LOC_360/a_8_216# 0.08fF
C22865 AND2X1_LOC_95/Y OR2X1_LOC_576/A 0.03fF
C22866 OR2X1_LOC_405/A AND2X1_LOC_432/a_36_24# 0.00fF
C22867 OR2X1_LOC_676/Y INPUT_0 0.02fF
C22868 AND2X1_LOC_568/B OR2X1_LOC_91/A 0.02fF
C22869 AND2X1_LOC_330/a_8_24# OR2X1_LOC_59/Y 0.01fF
C22870 AND2X1_LOC_716/Y AND2X1_LOC_566/B 1.18fF
C22871 OR2X1_LOC_161/A OR2X1_LOC_162/A 0.01fF
C22872 OR2X1_LOC_530/a_8_216# OR2X1_LOC_39/A 0.01fF
C22873 AND2X1_LOC_729/Y OR2X1_LOC_312/a_36_216# 0.00fF
C22874 OR2X1_LOC_22/Y OR2X1_LOC_437/A 0.10fF
C22875 OR2X1_LOC_292/Y OR2X1_LOC_600/A 0.00fF
C22876 OR2X1_LOC_650/a_36_216# AND2X1_LOC_92/Y 0.00fF
C22877 OR2X1_LOC_833/Y OR2X1_LOC_833/B 0.02fF
C22878 OR2X1_LOC_160/A OR2X1_LOC_161/B 0.17fF
C22879 OR2X1_LOC_325/Y OR2X1_LOC_538/A 0.01fF
C22880 AND2X1_LOC_22/Y OR2X1_LOC_831/a_8_216# 0.01fF
C22881 AND2X1_LOC_721/Y OR2X1_LOC_406/a_36_216# 0.00fF
C22882 AND2X1_LOC_56/B OR2X1_LOC_121/A 0.05fF
C22883 OR2X1_LOC_121/B OR2X1_LOC_771/B 0.03fF
C22884 AND2X1_LOC_566/B AND2X1_LOC_654/Y 0.02fF
C22885 INPUT_4 AND2X1_LOC_639/B 0.07fF
C22886 OR2X1_LOC_139/A OR2X1_LOC_793/A 0.08fF
C22887 OR2X1_LOC_40/Y AND2X1_LOC_641/a_36_24# 0.00fF
C22888 AND2X1_LOC_508/A OR2X1_LOC_51/Y 0.52fF
C22889 OR2X1_LOC_168/B OR2X1_LOC_78/B 0.19fF
C22890 AND2X1_LOC_40/Y OR2X1_LOC_389/A 0.25fF
C22891 OR2X1_LOC_323/A OR2X1_LOC_485/A 0.06fF
C22892 OR2X1_LOC_673/A OR2X1_LOC_80/A 0.05fF
C22893 AND2X1_LOC_12/Y OR2X1_LOC_549/A 0.08fF
C22894 OR2X1_LOC_589/A AND2X1_LOC_435/a_8_24# 0.02fF
C22895 AND2X1_LOC_340/Y OR2X1_LOC_85/A 0.08fF
C22896 OR2X1_LOC_45/B OR2X1_LOC_43/A 0.13fF
C22897 OR2X1_LOC_44/Y AND2X1_LOC_771/a_8_24# 0.01fF
C22898 AND2X1_LOC_339/B OR2X1_LOC_265/Y 0.03fF
C22899 AND2X1_LOC_840/B OR2X1_LOC_373/Y 0.10fF
C22900 AND2X1_LOC_535/Y AND2X1_LOC_809/A 0.01fF
C22901 OR2X1_LOC_121/B OR2X1_LOC_776/A 0.00fF
C22902 OR2X1_LOC_660/Y OR2X1_LOC_663/A 0.74fF
C22903 OR2X1_LOC_501/B OR2X1_LOC_499/B 0.11fF
C22904 OR2X1_LOC_677/Y AND2X1_LOC_663/A 0.05fF
C22905 OR2X1_LOC_703/B OR2X1_LOC_356/A 0.01fF
C22906 OR2X1_LOC_154/A OR2X1_LOC_390/A 0.04fF
C22907 OR2X1_LOC_244/A OR2X1_LOC_141/a_36_216# 0.00fF
C22908 OR2X1_LOC_467/A OR2X1_LOC_478/a_36_216# 0.00fF
C22909 AND2X1_LOC_70/Y OR2X1_LOC_175/B 0.00fF
C22910 AND2X1_LOC_787/A OR2X1_LOC_312/Y 0.02fF
C22911 OR2X1_LOC_49/A OR2X1_LOC_827/a_8_216# 0.04fF
C22912 AND2X1_LOC_458/a_8_24# AND2X1_LOC_786/Y 0.02fF
C22913 AND2X1_LOC_22/Y OR2X1_LOC_787/Y 0.04fF
C22914 OR2X1_LOC_354/A OR2X1_LOC_538/A 0.37fF
C22915 AND2X1_LOC_361/A OR2X1_LOC_595/A 1.01fF
C22916 OR2X1_LOC_51/Y OR2X1_LOC_48/B 0.07fF
C22917 OR2X1_LOC_249/a_8_216# OR2X1_LOC_66/A 0.02fF
C22918 INPUT_0 AND2X1_LOC_642/Y 0.36fF
C22919 AND2X1_LOC_663/B AND2X1_LOC_772/Y 0.01fF
C22920 OR2X1_LOC_389/A OR2X1_LOC_537/A 1.13fF
C22921 AND2X1_LOC_333/a_8_24# OR2X1_LOC_171/Y 0.01fF
C22922 OR2X1_LOC_47/Y AND2X1_LOC_740/a_8_24# 0.03fF
C22923 OR2X1_LOC_600/A OR2X1_LOC_69/A 0.03fF
C22924 OR2X1_LOC_43/A OR2X1_LOC_382/A 0.02fF
C22925 OR2X1_LOC_51/Y OR2X1_LOC_18/Y 0.27fF
C22926 OR2X1_LOC_70/A OR2X1_LOC_11/a_8_216# 0.39fF
C22927 OR2X1_LOC_625/Y OR2X1_LOC_56/A 0.07fF
C22928 VDD AND2X1_LOC_449/Y 0.21fF
C22929 AND2X1_LOC_723/Y AND2X1_LOC_168/a_8_24# 0.02fF
C22930 AND2X1_LOC_40/Y AND2X1_LOC_177/a_8_24# 0.01fF
C22931 AND2X1_LOC_219/a_8_24# OR2X1_LOC_316/Y 0.01fF
C22932 OR2X1_LOC_256/Y AND2X1_LOC_344/a_8_24# 0.05fF
C22933 OR2X1_LOC_405/A OR2X1_LOC_78/A 0.18fF
C22934 AND2X1_LOC_334/Y OR2X1_LOC_316/Y 0.01fF
C22935 OR2X1_LOC_240/B AND2X1_LOC_232/a_8_24# 0.04fF
C22936 OR2X1_LOC_814/A OR2X1_LOC_363/a_36_216# 0.00fF
C22937 AND2X1_LOC_566/B OR2X1_LOC_312/Y 0.03fF
C22938 OR2X1_LOC_45/B OR2X1_LOC_372/a_36_216# 0.00fF
C22939 AND2X1_LOC_843/Y AND2X1_LOC_850/A 0.31fF
C22940 AND2X1_LOC_366/a_36_24# AND2X1_LOC_848/Y 0.01fF
C22941 AND2X1_LOC_95/Y AND2X1_LOC_41/A 0.10fF
C22942 OR2X1_LOC_235/B OR2X1_LOC_624/A 0.05fF
C22943 OR2X1_LOC_616/Y AND2X1_LOC_663/A 0.49fF
C22944 AND2X1_LOC_59/Y OR2X1_LOC_78/B 0.20fF
C22945 OR2X1_LOC_405/A OR2X1_LOC_458/B 0.16fF
C22946 AND2X1_LOC_190/a_8_24# OR2X1_LOC_36/Y 0.00fF
C22947 OR2X1_LOC_539/A OR2X1_LOC_856/B 0.05fF
C22948 AND2X1_LOC_496/a_8_24# OR2X1_LOC_549/A 0.01fF
C22949 OR2X1_LOC_45/B AND2X1_LOC_685/a_8_24# 0.01fF
C22950 OR2X1_LOC_158/A AND2X1_LOC_34/a_36_24# 0.01fF
C22951 OR2X1_LOC_599/A AND2X1_LOC_657/Y 0.03fF
C22952 OR2X1_LOC_404/a_8_216# OR2X1_LOC_78/Y 0.04fF
C22953 OR2X1_LOC_536/Y OR2X1_LOC_585/A 0.01fF
C22954 OR2X1_LOC_160/A OR2X1_LOC_435/B 0.07fF
C22955 OR2X1_LOC_494/Y OR2X1_LOC_667/a_36_216# 0.00fF
C22956 OR2X1_LOC_459/A AND2X1_LOC_43/B 0.07fF
C22957 OR2X1_LOC_168/B AND2X1_LOC_601/a_36_24# 0.00fF
C22958 AND2X1_LOC_784/Y OR2X1_LOC_74/A 0.02fF
C22959 OR2X1_LOC_441/Y AND2X1_LOC_621/Y 0.03fF
C22960 OR2X1_LOC_462/B INPUT_0 0.11fF
C22961 OR2X1_LOC_715/B OR2X1_LOC_479/Y 0.05fF
C22962 AND2X1_LOC_113/a_36_24# OR2X1_LOC_427/A 0.01fF
C22963 AND2X1_LOC_508/B OR2X1_LOC_7/A 0.00fF
C22964 OR2X1_LOC_59/Y OR2X1_LOC_701/a_8_216# 0.02fF
C22965 AND2X1_LOC_73/a_36_24# AND2X1_LOC_56/B 0.01fF
C22966 OR2X1_LOC_19/B OR2X1_LOC_633/A 0.05fF
C22967 AND2X1_LOC_509/Y OR2X1_LOC_44/Y 0.01fF
C22968 OR2X1_LOC_864/A AND2X1_LOC_92/Y 0.03fF
C22969 OR2X1_LOC_59/Y AND2X1_LOC_806/A 0.03fF
C22970 AND2X1_LOC_110/Y AND2X1_LOC_111/a_8_24# 0.09fF
C22971 OR2X1_LOC_479/Y OR2X1_LOC_543/A 0.03fF
C22972 AND2X1_LOC_512/Y AND2X1_LOC_319/A 0.06fF
C22973 AND2X1_LOC_70/Y OR2X1_LOC_355/B 0.03fF
C22974 AND2X1_LOC_173/a_8_24# OR2X1_LOC_161/A 0.00fF
C22975 OR2X1_LOC_160/B AND2X1_LOC_42/B 0.21fF
C22976 AND2X1_LOC_508/a_8_24# OR2X1_LOC_7/A 0.04fF
C22977 AND2X1_LOC_370/a_8_24# OR2X1_LOC_417/A 0.04fF
C22978 D_INPUT_7 AND2X1_LOC_2/Y 0.98fF
C22979 AND2X1_LOC_752/a_8_24# OR2X1_LOC_375/A 0.01fF
C22980 OR2X1_LOC_160/A OR2X1_LOC_61/Y 0.04fF
C22981 OR2X1_LOC_643/A OR2X1_LOC_624/a_8_216# 0.01fF
C22982 AND2X1_LOC_92/Y OR2X1_LOC_240/A 0.82fF
C22983 AND2X1_LOC_191/Y AND2X1_LOC_629/a_8_24# 0.05fF
C22984 OR2X1_LOC_287/B OR2X1_LOC_363/A 0.02fF
C22985 OR2X1_LOC_105/Y OR2X1_LOC_579/B 0.10fF
C22986 OR2X1_LOC_837/B OR2X1_LOC_32/B 0.43fF
C22987 AND2X1_LOC_456/B AND2X1_LOC_859/Y 0.10fF
C22988 VDD AND2X1_LOC_212/B 0.26fF
C22989 OR2X1_LOC_660/a_8_216# OR2X1_LOC_130/A 0.49fF
C22990 AND2X1_LOC_474/A OR2X1_LOC_585/A 0.08fF
C22991 OR2X1_LOC_675/A OR2X1_LOC_733/A 0.62fF
C22992 VDD OR2X1_LOC_123/B -0.00fF
C22993 OR2X1_LOC_316/Y AND2X1_LOC_649/B 0.00fF
C22994 AND2X1_LOC_259/Y AND2X1_LOC_296/a_36_24# 0.00fF
C22995 OR2X1_LOC_814/A AND2X1_LOC_65/A 0.07fF
C22996 OR2X1_LOC_585/A AND2X1_LOC_240/a_8_24# 0.01fF
C22997 AND2X1_LOC_330/a_8_24# OR2X1_LOC_70/Y 0.01fF
C22998 VDD OR2X1_LOC_829/Y 0.15fF
C22999 AND2X1_LOC_658/B OR2X1_LOC_527/Y 0.07fF
C23000 OR2X1_LOC_17/Y OR2X1_LOC_12/a_8_216# 0.01fF
C23001 AND2X1_LOC_276/Y OR2X1_LOC_59/Y 0.02fF
C23002 OR2X1_LOC_680/A OR2X1_LOC_48/B 0.07fF
C23003 AND2X1_LOC_70/Y AND2X1_LOC_674/a_8_24# 0.03fF
C23004 OR2X1_LOC_671/Y INPUT_1 0.01fF
C23005 OR2X1_LOC_185/A OR2X1_LOC_539/Y 0.03fF
C23006 OR2X1_LOC_31/Y OR2X1_LOC_373/Y 0.01fF
C23007 AND2X1_LOC_364/A OR2X1_LOC_6/A 0.28fF
C23008 AND2X1_LOC_850/A OR2X1_LOC_7/A 0.03fF
C23009 OR2X1_LOC_184/Y OR2X1_LOC_184/a_36_216# 0.00fF
C23010 OR2X1_LOC_448/Y OR2X1_LOC_803/B 0.26fF
C23011 OR2X1_LOC_574/A OR2X1_LOC_776/a_8_216# 0.16fF
C23012 OR2X1_LOC_680/A OR2X1_LOC_18/Y 0.06fF
C23013 AND2X1_LOC_211/B AND2X1_LOC_857/Y 0.04fF
C23014 OR2X1_LOC_160/A OR2X1_LOC_87/a_8_216# 0.01fF
C23015 OR2X1_LOC_40/Y OR2X1_LOC_815/A 0.01fF
C23016 OR2X1_LOC_151/A OR2X1_LOC_532/B 0.79fF
C23017 OR2X1_LOC_237/a_36_216# OR2X1_LOC_39/A 0.01fF
C23018 OR2X1_LOC_510/A OR2X1_LOC_814/A 0.03fF
C23019 AND2X1_LOC_139/a_36_24# OR2X1_LOC_7/A 0.00fF
C23020 AND2X1_LOC_59/Y OR2X1_LOC_375/A 1.23fF
C23021 OR2X1_LOC_865/B OR2X1_LOC_859/B 0.36fF
C23022 AND2X1_LOC_77/a_8_24# OR2X1_LOC_78/A -0.01fF
C23023 VDD OR2X1_LOC_781/Y 0.08fF
C23024 OR2X1_LOC_703/B AND2X1_LOC_43/B 0.16fF
C23025 OR2X1_LOC_744/A OR2X1_LOC_277/a_8_216# 0.01fF
C23026 OR2X1_LOC_6/B AND2X1_LOC_667/a_36_24# 0.00fF
C23027 AND2X1_LOC_702/Y OR2X1_LOC_619/Y 0.16fF
C23028 OR2X1_LOC_109/a_8_216# OR2X1_LOC_26/Y 0.01fF
C23029 AND2X1_LOC_715/A OR2X1_LOC_22/Y 0.01fF
C23030 AND2X1_LOC_658/B AND2X1_LOC_574/A 0.20fF
C23031 AND2X1_LOC_95/Y OR2X1_LOC_631/B 0.16fF
C23032 OR2X1_LOC_753/A OR2X1_LOC_394/Y 0.05fF
C23033 VDD OR2X1_LOC_7/Y 0.10fF
C23034 AND2X1_LOC_845/Y AND2X1_LOC_244/a_8_24# 0.03fF
C23035 OR2X1_LOC_87/A AND2X1_LOC_43/B 0.10fF
C23036 OR2X1_LOC_467/A AND2X1_LOC_425/Y 0.07fF
C23037 OR2X1_LOC_411/Y OR2X1_LOC_22/Y 0.03fF
C23038 OR2X1_LOC_405/A OR2X1_LOC_155/A 0.03fF
C23039 AND2X1_LOC_29/a_8_24# OR2X1_LOC_87/Y 0.23fF
C23040 OR2X1_LOC_470/B OR2X1_LOC_477/Y 0.01fF
C23041 OR2X1_LOC_3/Y OR2X1_LOC_281/a_8_216# 0.01fF
C23042 OR2X1_LOC_377/A OR2X1_LOC_585/A 0.03fF
C23043 AND2X1_LOC_36/Y OR2X1_LOC_446/B 0.76fF
C23044 OR2X1_LOC_235/B OR2X1_LOC_54/Y 0.08fF
C23045 OR2X1_LOC_287/A OR2X1_LOC_287/a_8_216# 0.01fF
C23046 AND2X1_LOC_729/Y OR2X1_LOC_52/B 0.03fF
C23047 AND2X1_LOC_44/Y OR2X1_LOC_512/a_8_216# 0.01fF
C23048 OR2X1_LOC_482/Y OR2X1_LOC_615/Y 0.00fF
C23049 OR2X1_LOC_636/A AND2X1_LOC_11/Y 0.04fF
C23050 OR2X1_LOC_529/Y AND2X1_LOC_621/Y 0.08fF
C23051 OR2X1_LOC_856/B AND2X1_LOC_111/a_36_24# 0.01fF
C23052 AND2X1_LOC_12/Y OR2X1_LOC_401/Y 0.03fF
C23053 AND2X1_LOC_768/a_8_24# AND2X1_LOC_227/Y 0.01fF
C23054 AND2X1_LOC_393/a_8_24# OR2X1_LOC_400/B 0.01fF
C23055 AND2X1_LOC_22/Y AND2X1_LOC_52/Y 0.03fF
C23056 INPUT_3 AND2X1_LOC_42/B 0.34fF
C23057 OR2X1_LOC_426/B OR2X1_LOC_95/Y 0.10fF
C23058 OR2X1_LOC_85/A OR2X1_LOC_585/A 0.06fF
C23059 OR2X1_LOC_193/A OR2X1_LOC_194/B 0.13fF
C23060 OR2X1_LOC_8/Y OR2X1_LOC_62/A 0.06fF
C23061 AND2X1_LOC_191/B AND2X1_LOC_866/A 0.09fF
C23062 OR2X1_LOC_481/A OR2X1_LOC_257/a_36_216# 0.00fF
C23063 OR2X1_LOC_76/B OR2X1_LOC_76/A 0.04fF
C23064 AND2X1_LOC_784/A OR2X1_LOC_52/B 0.75fF
C23065 OR2X1_LOC_185/Y OR2X1_LOC_287/B 0.05fF
C23066 AND2X1_LOC_72/B OR2X1_LOC_719/B 0.03fF
C23067 OR2X1_LOC_62/B OR2X1_LOC_574/a_8_216# 0.01fF
C23068 OR2X1_LOC_47/Y AND2X1_LOC_285/Y 0.02fF
C23069 AND2X1_LOC_42/B OR2X1_LOC_266/a_8_216# 0.11fF
C23070 OR2X1_LOC_382/Y OR2X1_LOC_417/A 0.01fF
C23071 OR2X1_LOC_3/Y OR2X1_LOC_6/A 0.36fF
C23072 AND2X1_LOC_512/a_36_24# OR2X1_LOC_36/Y 0.01fF
C23073 OR2X1_LOC_305/a_36_216# OR2X1_LOC_3/Y 0.02fF
C23074 OR2X1_LOC_682/a_36_216# OR2X1_LOC_682/Y -0.00fF
C23075 OR2X1_LOC_19/B OR2X1_LOC_256/a_8_216# 0.02fF
C23076 AND2X1_LOC_512/Y AND2X1_LOC_170/B 0.00fF
C23077 OR2X1_LOC_485/A OR2X1_LOC_601/Y 0.01fF
C23078 OR2X1_LOC_372/Y OR2X1_LOC_371/Y 0.12fF
C23079 OR2X1_LOC_51/Y AND2X1_LOC_620/Y 0.05fF
C23080 OR2X1_LOC_61/B D_INPUT_0 0.23fF
C23081 OR2X1_LOC_702/A OR2X1_LOC_269/B 0.03fF
C23082 AND2X1_LOC_753/B OR2X1_LOC_228/a_8_216# 0.02fF
C23083 AND2X1_LOC_367/A AND2X1_LOC_851/B 0.10fF
C23084 OR2X1_LOC_779/Y OR2X1_LOC_78/A 0.01fF
C23085 OR2X1_LOC_426/A OR2X1_LOC_31/Y 0.03fF
C23086 AND2X1_LOC_31/Y OR2X1_LOC_741/a_36_216# 0.00fF
C23087 AND2X1_LOC_91/B OR2X1_LOC_571/Y 0.03fF
C23088 OR2X1_LOC_71/a_8_216# D_INPUT_0 0.02fF
C23089 AND2X1_LOC_480/A AND2X1_LOC_222/Y 0.00fF
C23090 AND2X1_LOC_284/a_8_24# OR2X1_LOC_13/B 0.03fF
C23091 OR2X1_LOC_64/Y OR2X1_LOC_591/A 0.05fF
C23092 OR2X1_LOC_154/A OR2X1_LOC_750/A 0.07fF
C23093 AND2X1_LOC_580/B AND2X1_LOC_663/B 0.00fF
C23094 AND2X1_LOC_624/B AND2X1_LOC_663/A 0.03fF
C23095 OR2X1_LOC_840/A OR2X1_LOC_223/A 0.03fF
C23096 OR2X1_LOC_36/Y OR2X1_LOC_65/Y 0.01fF
C23097 OR2X1_LOC_210/B AND2X1_LOC_51/Y 0.13fF
C23098 OR2X1_LOC_715/B OR2X1_LOC_68/B 0.01fF
C23099 OR2X1_LOC_147/a_36_216# AND2X1_LOC_36/Y 0.02fF
C23100 OR2X1_LOC_405/a_36_216# OR2X1_LOC_532/B 0.00fF
C23101 OR2X1_LOC_485/A OR2X1_LOC_754/A 0.08fF
C23102 AND2X1_LOC_329/a_8_24# AND2X1_LOC_51/Y 0.02fF
C23103 OR2X1_LOC_541/A OR2X1_LOC_241/B 0.03fF
C23104 OR2X1_LOC_59/Y AND2X1_LOC_405/a_8_24# 0.02fF
C23105 AND2X1_LOC_64/Y OR2X1_LOC_308/Y 1.80fF
C23106 AND2X1_LOC_523/Y OR2X1_LOC_7/A 0.10fF
C23107 OR2X1_LOC_420/a_36_216# OR2X1_LOC_64/Y 0.02fF
C23108 OR2X1_LOC_22/Y OR2X1_LOC_753/A 0.03fF
C23109 OR2X1_LOC_857/A OR2X1_LOC_771/B 0.03fF
C23110 AND2X1_LOC_140/a_8_24# AND2X1_LOC_141/B -0.06fF
C23111 AND2X1_LOC_390/B AND2X1_LOC_729/B 0.62fF
C23112 AND2X1_LOC_72/B OR2X1_LOC_736/A 0.02fF
C23113 OR2X1_LOC_168/Y OR2X1_LOC_170/a_36_216# 0.03fF
C23114 INPUT_4 OR2X1_LOC_31/Y 0.03fF
C23115 D_INPUT_0 OR2X1_LOC_205/a_8_216# 0.01fF
C23116 OR2X1_LOC_6/B OR2X1_LOC_71/A 0.91fF
C23117 AND2X1_LOC_22/Y OR2X1_LOC_523/a_8_216# 0.06fF
C23118 OR2X1_LOC_485/A AND2X1_LOC_844/a_36_24# 0.00fF
C23119 AND2X1_LOC_40/Y OR2X1_LOC_801/B 0.14fF
C23120 OR2X1_LOC_504/Y AND2X1_LOC_806/A 0.03fF
C23121 AND2X1_LOC_566/B OR2X1_LOC_13/B 0.03fF
C23122 OR2X1_LOC_185/Y OR2X1_LOC_436/Y 0.03fF
C23123 OR2X1_LOC_569/B OR2X1_LOC_569/a_8_216# 0.07fF
C23124 AND2X1_LOC_512/Y OR2X1_LOC_331/Y 0.57fF
C23125 OR2X1_LOC_428/A OR2X1_LOC_387/A 0.06fF
C23126 OR2X1_LOC_91/Y OR2X1_LOC_47/Y 0.15fF
C23127 OR2X1_LOC_698/a_36_216# AND2X1_LOC_793/B 0.02fF
C23128 AND2X1_LOC_102/a_8_24# AND2X1_LOC_47/Y 0.01fF
C23129 OR2X1_LOC_64/Y AND2X1_LOC_307/Y 0.02fF
C23130 AND2X1_LOC_785/a_8_24# AND2X1_LOC_564/B 0.02fF
C23131 OR2X1_LOC_147/B OR2X1_LOC_543/a_8_216# 0.06fF
C23132 OR2X1_LOC_280/Y AND2X1_LOC_845/Y 0.02fF
C23133 OR2X1_LOC_680/A AND2X1_LOC_620/Y 0.03fF
C23134 AND2X1_LOC_73/a_8_24# OR2X1_LOC_71/A 0.04fF
C23135 AND2X1_LOC_36/Y OR2X1_LOC_719/B 0.02fF
C23136 OR2X1_LOC_599/A OR2X1_LOC_146/Y 0.00fF
C23137 AND2X1_LOC_708/a_8_24# AND2X1_LOC_712/B 0.01fF
C23138 AND2X1_LOC_342/Y AND2X1_LOC_721/A 0.01fF
C23139 OR2X1_LOC_244/A AND2X1_LOC_42/B 0.06fF
C23140 OR2X1_LOC_487/Y OR2X1_LOC_417/A 0.01fF
C23141 OR2X1_LOC_632/A OR2X1_LOC_598/A 0.04fF
C23142 AND2X1_LOC_564/A AND2X1_LOC_564/B 0.02fF
C23143 OR2X1_LOC_743/A OR2X1_LOC_95/Y 0.06fF
C23144 OR2X1_LOC_213/a_8_216# OR2X1_LOC_213/B 0.39fF
C23145 OR2X1_LOC_502/A OR2X1_LOC_80/A 0.10fF
C23146 OR2X1_LOC_47/Y OR2X1_LOC_371/a_8_216# 0.14fF
C23147 OR2X1_LOC_837/B OR2X1_LOC_68/B 0.03fF
C23148 OR2X1_LOC_3/Y AND2X1_LOC_139/A 0.03fF
C23149 AND2X1_LOC_459/Y OR2X1_LOC_378/a_8_216# 0.47fF
C23150 AND2X1_LOC_851/B OR2X1_LOC_74/A 0.01fF
C23151 OR2X1_LOC_779/Y OR2X1_LOC_155/A 0.00fF
C23152 OR2X1_LOC_468/A OR2X1_LOC_593/B 0.00fF
C23153 OR2X1_LOC_189/Y OR2X1_LOC_47/Y 7.71fF
C23154 OR2X1_LOC_542/B AND2X1_LOC_36/Y 0.03fF
C23155 AND2X1_LOC_22/Y OR2X1_LOC_576/A 0.22fF
C23156 AND2X1_LOC_555/Y AND2X1_LOC_363/a_8_24# 0.01fF
C23157 OR2X1_LOC_744/A OR2X1_LOC_142/a_36_216# 0.00fF
C23158 OR2X1_LOC_62/B OR2X1_LOC_62/a_8_216# 0.10fF
C23159 OR2X1_LOC_152/Y OR2X1_LOC_47/Y 0.24fF
C23160 AND2X1_LOC_743/a_8_24# OR2X1_LOC_161/B 0.01fF
C23161 OR2X1_LOC_266/A OR2X1_LOC_161/B 0.00fF
C23162 OR2X1_LOC_215/Y OR2X1_LOC_68/B 0.01fF
C23163 AND2X1_LOC_230/a_36_24# OR2X1_LOC_68/B 0.00fF
C23164 AND2X1_LOC_5/a_8_24# D_INPUT_0 0.02fF
C23165 OR2X1_LOC_739/A OR2X1_LOC_151/a_36_216# 0.00fF
C23166 OR2X1_LOC_482/Y AND2X1_LOC_242/B 0.07fF
C23167 INPUT_1 OR2X1_LOC_532/B 1.02fF
C23168 OR2X1_LOC_564/A OR2X1_LOC_192/B 0.13fF
C23169 OR2X1_LOC_457/a_8_216# AND2X1_LOC_31/Y 0.05fF
C23170 OR2X1_LOC_617/a_8_216# AND2X1_LOC_624/B 0.01fF
C23171 OR2X1_LOC_36/Y OR2X1_LOC_72/Y 0.49fF
C23172 OR2X1_LOC_791/a_8_216# OR2X1_LOC_792/a_8_216# 0.47fF
C23173 AND2X1_LOC_557/Y AND2X1_LOC_657/A 0.10fF
C23174 OR2X1_LOC_523/B AND2X1_LOC_44/Y 0.03fF
C23175 OR2X1_LOC_417/Y OR2X1_LOC_47/Y 0.00fF
C23176 OR2X1_LOC_297/a_8_216# AND2X1_LOC_789/Y 0.02fF
C23177 OR2X1_LOC_291/Y OR2X1_LOC_47/Y 1.99fF
C23178 OR2X1_LOC_74/A OR2X1_LOC_595/Y 0.03fF
C23179 OR2X1_LOC_258/a_8_216# AND2X1_LOC_848/A 0.03fF
C23180 AND2X1_LOC_40/Y OR2X1_LOC_182/a_8_216# 0.01fF
C23181 OR2X1_LOC_9/Y OR2X1_LOC_428/A 0.09fF
C23182 AND2X1_LOC_515/a_8_24# AND2X1_LOC_212/Y 0.03fF
C23183 OR2X1_LOC_791/B OR2X1_LOC_366/Y 0.14fF
C23184 OR2X1_LOC_35/a_8_216# OR2X1_LOC_338/A 0.01fF
C23185 OR2X1_LOC_628/Y OR2X1_LOC_615/Y 0.01fF
C23186 OR2X1_LOC_70/Y AND2X1_LOC_405/a_8_24# 0.01fF
C23187 OR2X1_LOC_87/A OR2X1_LOC_357/A 0.02fF
C23188 OR2X1_LOC_676/Y AND2X1_LOC_7/B 0.08fF
C23189 OR2X1_LOC_97/A OR2X1_LOC_325/B 0.12fF
C23190 OR2X1_LOC_70/Y AND2X1_LOC_486/a_8_24# 0.04fF
C23191 OR2X1_LOC_841/a_8_216# OR2X1_LOC_776/A 0.06fF
C23192 OR2X1_LOC_52/B OR2X1_LOC_172/Y 0.00fF
C23193 OR2X1_LOC_39/A OR2X1_LOC_437/A 1.74fF
C23194 OR2X1_LOC_12/Y OR2X1_LOC_131/a_8_216# 0.02fF
C23195 OR2X1_LOC_774/Y OR2X1_LOC_561/B 0.50fF
C23196 OR2X1_LOC_601/a_8_216# OR2X1_LOC_47/Y 0.00fF
C23197 AND2X1_LOC_2/a_36_24# INPUT_6 0.00fF
C23198 OR2X1_LOC_51/B OR2X1_LOC_22/A 0.03fF
C23199 AND2X1_LOC_721/A OR2X1_LOC_54/Y 0.02fF
C23200 OR2X1_LOC_95/Y OR2X1_LOC_409/B 0.01fF
C23201 OR2X1_LOC_158/A OR2X1_LOC_589/A 0.03fF
C23202 OR2X1_LOC_197/A OR2X1_LOC_651/A 0.04fF
C23203 OR2X1_LOC_45/B AND2X1_LOC_776/a_8_24# 0.01fF
C23204 OR2X1_LOC_235/Y OR2X1_LOC_71/A 0.01fF
C23205 AND2X1_LOC_769/a_36_24# OR2X1_LOC_744/A 0.00fF
C23206 AND2X1_LOC_92/Y OR2X1_LOC_121/A 0.03fF
C23207 OR2X1_LOC_854/a_8_216# OR2X1_LOC_354/a_8_216# 0.47fF
C23208 OR2X1_LOC_354/A OR2X1_LOC_356/B 0.08fF
C23209 AND2X1_LOC_763/a_8_24# OR2X1_LOC_855/A 0.20fF
C23210 OR2X1_LOC_450/B OR2X1_LOC_161/B 0.25fF
C23211 OR2X1_LOC_756/B OR2X1_LOC_334/a_8_216# 0.02fF
C23212 OR2X1_LOC_188/Y OR2X1_LOC_541/A 0.02fF
C23213 AND2X1_LOC_340/Y OR2X1_LOC_51/Y 0.09fF
C23214 OR2X1_LOC_770/A OR2X1_LOC_78/Y 0.01fF
C23215 OR2X1_LOC_276/B OR2X1_LOC_276/a_8_216# 0.02fF
C23216 OR2X1_LOC_177/a_8_216# AND2X1_LOC_657/Y 0.33fF
C23217 OR2X1_LOC_151/A OR2X1_LOC_440/B 0.01fF
C23218 AND2X1_LOC_91/B OR2X1_LOC_274/Y 0.05fF
C23219 AND2X1_LOC_658/A AND2X1_LOC_212/Y 0.07fF
C23220 OR2X1_LOC_696/A OR2X1_LOC_278/Y 0.03fF
C23221 AND2X1_LOC_91/B OR2X1_LOC_392/A 0.01fF
C23222 AND2X1_LOC_22/Y AND2X1_LOC_41/A 0.10fF
C23223 AND2X1_LOC_141/B AND2X1_LOC_217/a_8_24# 0.07fF
C23224 OR2X1_LOC_244/B OR2X1_LOC_576/A 0.00fF
C23225 AND2X1_LOC_472/B OR2X1_LOC_376/Y 0.09fF
C23226 D_INPUT_3 OR2X1_LOC_47/Y 0.08fF
C23227 OR2X1_LOC_589/A AND2X1_LOC_537/a_36_24# 0.00fF
C23228 AND2X1_LOC_211/B OR2X1_LOC_437/A 0.07fF
C23229 OR2X1_LOC_62/A OR2X1_LOC_619/a_36_216# 0.00fF
C23230 OR2X1_LOC_696/A AND2X1_LOC_662/B 0.07fF
C23231 AND2X1_LOC_391/Y OR2X1_LOC_12/Y 0.04fF
C23232 OR2X1_LOC_158/A AND2X1_LOC_337/a_8_24# 0.04fF
C23233 OR2X1_LOC_91/A OR2X1_LOC_12/Y 0.41fF
C23234 AND2X1_LOC_56/B AND2X1_LOC_36/Y 1.46fF
C23235 OR2X1_LOC_653/Y OR2X1_LOC_390/a_8_216# 0.02fF
C23236 AND2X1_LOC_70/Y OR2X1_LOC_786/A 0.01fF
C23237 OR2X1_LOC_449/B OR2X1_LOC_593/B 0.66fF
C23238 OR2X1_LOC_40/Y AND2X1_LOC_657/Y 0.03fF
C23239 OR2X1_LOC_158/A OR2X1_LOC_297/A 0.01fF
C23240 OR2X1_LOC_696/A OR2X1_LOC_95/a_8_216# 0.02fF
C23241 AND2X1_LOC_8/Y AND2X1_LOC_36/Y 0.24fF
C23242 AND2X1_LOC_191/B OR2X1_LOC_40/Y 0.03fF
C23243 OR2X1_LOC_756/B OR2X1_LOC_486/Y 0.03fF
C23244 AND2X1_LOC_535/Y OR2X1_LOC_56/A 0.03fF
C23245 AND2X1_LOC_658/B AND2X1_LOC_565/a_8_24# 0.03fF
C23246 AND2X1_LOC_215/Y AND2X1_LOC_61/Y 0.92fF
C23247 AND2X1_LOC_866/A AND2X1_LOC_848/A 0.08fF
C23248 OR2X1_LOC_40/Y AND2X1_LOC_469/B 0.09fF
C23249 OR2X1_LOC_97/A OR2X1_LOC_788/a_36_216# 0.00fF
C23250 OR2X1_LOC_6/B OR2X1_LOC_59/Y 0.05fF
C23251 OR2X1_LOC_447/Y OR2X1_LOC_779/B 0.09fF
C23252 OR2X1_LOC_485/A OR2X1_LOC_142/Y 0.02fF
C23253 OR2X1_LOC_661/a_8_216# AND2X1_LOC_7/B 0.01fF
C23254 AND2X1_LOC_501/Y AND2X1_LOC_570/Y 0.00fF
C23255 AND2X1_LOC_84/Y OR2X1_LOC_65/B 0.02fF
C23256 OR2X1_LOC_47/Y AND2X1_LOC_483/Y 0.17fF
C23257 AND2X1_LOC_362/a_8_24# AND2X1_LOC_243/Y 0.01fF
C23258 AND2X1_LOC_21/Y AND2X1_LOC_36/Y 0.69fF
C23259 AND2X1_LOC_592/Y AND2X1_LOC_605/Y 0.84fF
C23260 OR2X1_LOC_591/Y AND2X1_LOC_722/A 0.79fF
C23261 AND2X1_LOC_794/B OR2X1_LOC_516/B 0.09fF
C23262 OR2X1_LOC_158/A OR2X1_LOC_275/Y 0.02fF
C23263 VDD OR2X1_LOC_25/Y 0.09fF
C23264 OR2X1_LOC_160/B OR2X1_LOC_778/a_8_216# 0.05fF
C23265 AND2X1_LOC_56/B OR2X1_LOC_334/A 0.03fF
C23266 AND2X1_LOC_573/Y AND2X1_LOC_576/Y 0.02fF
C23267 AND2X1_LOC_479/Y AND2X1_LOC_222/Y 0.02fF
C23268 AND2X1_LOC_22/Y OR2X1_LOC_662/A 0.46fF
C23269 OR2X1_LOC_40/Y AND2X1_LOC_733/Y 0.76fF
C23270 AND2X1_LOC_675/Y VDD 0.73fF
C23271 AND2X1_LOC_802/B AND2X1_LOC_388/a_8_24# 0.02fF
C23272 OR2X1_LOC_97/A OR2X1_LOC_405/Y 0.01fF
C23273 OR2X1_LOC_179/a_8_216# OR2X1_LOC_108/Y 0.02fF
C23274 OR2X1_LOC_462/B AND2X1_LOC_7/B 0.03fF
C23275 OR2X1_LOC_160/B OR2X1_LOC_663/A 0.04fF
C23276 OR2X1_LOC_41/a_8_216# OR2X1_LOC_41/Y 0.01fF
C23277 OR2X1_LOC_51/a_8_216# OR2X1_LOC_70/A 0.06fF
C23278 OR2X1_LOC_122/Y OR2X1_LOC_426/B 0.10fF
C23279 AND2X1_LOC_573/A OR2X1_LOC_12/Y 0.09fF
C23280 VDD AND2X1_LOC_194/a_8_24# -0.00fF
C23281 OR2X1_LOC_130/A AND2X1_LOC_44/Y 0.56fF
C23282 VDD OR2X1_LOC_516/B 0.18fF
C23283 OR2X1_LOC_69/Y AND2X1_LOC_202/Y 0.00fF
C23284 AND2X1_LOC_572/Y OR2X1_LOC_595/A 0.05fF
C23285 OR2X1_LOC_287/B OR2X1_LOC_366/A 0.01fF
C23286 AND2X1_LOC_47/Y OR2X1_LOC_71/A 0.08fF
C23287 OR2X1_LOC_121/B OR2X1_LOC_593/B 0.03fF
C23288 OR2X1_LOC_830/a_8_216# OR2X1_LOC_147/B 0.09fF
C23289 OR2X1_LOC_685/B OR2X1_LOC_161/B 0.17fF
C23290 OR2X1_LOC_497/Y OR2X1_LOC_816/A 0.01fF
C23291 AND2X1_LOC_59/Y OR2X1_LOC_549/A 0.06fF
C23292 OR2X1_LOC_95/Y OR2X1_LOC_599/a_8_216# 0.02fF
C23293 OR2X1_LOC_52/B AND2X1_LOC_206/a_8_24# 0.01fF
C23294 INPUT_0 AND2X1_LOC_820/B 0.00fF
C23295 OR2X1_LOC_158/A AND2X1_LOC_365/A 3.76fF
C23296 AND2X1_LOC_41/A OR2X1_LOC_244/B 0.00fF
C23297 AND2X1_LOC_292/a_8_24# AND2X1_LOC_44/Y 0.01fF
C23298 OR2X1_LOC_215/a_8_216# AND2X1_LOC_31/Y 0.01fF
C23299 AND2X1_LOC_593/a_36_24# OR2X1_LOC_48/B 0.01fF
C23300 AND2X1_LOC_217/Y OR2X1_LOC_18/Y 0.01fF
C23301 OR2X1_LOC_318/B OR2X1_LOC_543/a_8_216# 0.07fF
C23302 AND2X1_LOC_41/A OR2X1_LOC_706/A 0.01fF
C23303 OR2X1_LOC_711/B OR2X1_LOC_154/A 0.12fF
C23304 AND2X1_LOC_793/Y AND2X1_LOC_793/B 0.01fF
C23305 AND2X1_LOC_152/a_8_24# OR2X1_LOC_740/B 0.15fF
C23306 OR2X1_LOC_625/Y AND2X1_LOC_285/Y 0.03fF
C23307 OR2X1_LOC_508/A OR2X1_LOC_244/B 0.13fF
C23308 OR2X1_LOC_76/Y OR2X1_LOC_486/Y 0.03fF
C23309 OR2X1_LOC_591/Y OR2X1_LOC_599/A 0.06fF
C23310 OR2X1_LOC_476/Y OR2X1_LOC_392/B 0.01fF
C23311 AND2X1_LOC_443/Y AND2X1_LOC_804/Y 0.02fF
C23312 OR2X1_LOC_121/B AND2X1_LOC_273/a_8_24# 0.01fF
C23313 AND2X1_LOC_388/Y OR2X1_LOC_44/Y 0.03fF
C23314 AND2X1_LOC_794/A AND2X1_LOC_469/B 0.01fF
C23315 AND2X1_LOC_70/Y OR2X1_LOC_624/A 0.04fF
C23316 AND2X1_LOC_95/Y OR2X1_LOC_648/A 0.07fF
C23317 OR2X1_LOC_303/a_8_216# OR2X1_LOC_121/B 0.08fF
C23318 OR2X1_LOC_158/A OR2X1_LOC_43/A 0.53fF
C23319 OR2X1_LOC_671/Y OR2X1_LOC_827/a_8_216# 0.02fF
C23320 AND2X1_LOC_715/A OR2X1_LOC_39/A 0.02fF
C23321 INPUT_0 OR2X1_LOC_427/A 0.03fF
C23322 AND2X1_LOC_573/a_36_24# AND2X1_LOC_501/Y 0.00fF
C23323 OR2X1_LOC_115/a_8_216# OR2X1_LOC_78/A 0.02fF
C23324 AND2X1_LOC_495/a_8_24# OR2X1_LOC_549/A 0.02fF
C23325 AND2X1_LOC_64/Y OR2X1_LOC_19/B 0.34fF
C23326 OR2X1_LOC_854/A OR2X1_LOC_567/a_8_216# 0.06fF
C23327 OR2X1_LOC_325/Y AND2X1_LOC_59/Y 0.00fF
C23328 OR2X1_LOC_840/A OR2X1_LOC_502/A 0.10fF
C23329 OR2X1_LOC_109/Y OR2X1_LOC_744/A 0.03fF
C23330 VDD OR2X1_LOC_189/A 0.21fF
C23331 OR2X1_LOC_364/A OR2X1_LOC_160/B 0.08fF
C23332 OR2X1_LOC_140/A OR2X1_LOC_203/Y 0.02fF
C23333 AND2X1_LOC_95/Y OR2X1_LOC_410/a_8_216# 0.01fF
C23334 AND2X1_LOC_557/Y VDD 0.21fF
C23335 OR2X1_LOC_185/Y OR2X1_LOC_160/B 0.21fF
C23336 OR2X1_LOC_207/a_8_216# AND2X1_LOC_41/Y 0.01fF
C23337 OR2X1_LOC_568/A OR2X1_LOC_566/Y 0.10fF
C23338 OR2X1_LOC_80/A OR2X1_LOC_398/a_8_216# 0.21fF
C23339 OR2X1_LOC_720/A OR2X1_LOC_66/A 0.01fF
C23340 AND2X1_LOC_716/Y OR2X1_LOC_92/Y 0.07fF
C23341 AND2X1_LOC_170/a_8_24# OR2X1_LOC_91/A 0.01fF
C23342 AND2X1_LOC_865/A AND2X1_LOC_807/Y 1.19fF
C23343 OR2X1_LOC_189/Y AND2X1_LOC_469/Y 0.03fF
C23344 OR2X1_LOC_779/B OR2X1_LOC_513/a_8_216# 0.05fF
C23345 AND2X1_LOC_851/a_8_24# OR2X1_LOC_39/A 0.04fF
C23346 OR2X1_LOC_71/A OR2X1_LOC_598/A 0.00fF
C23347 AND2X1_LOC_40/Y OR2X1_LOC_61/B 0.02fF
C23348 OR2X1_LOC_59/Y AND2X1_LOC_287/a_36_24# 0.00fF
C23349 OR2X1_LOC_96/Y OR2X1_LOC_6/a_8_216# 0.01fF
C23350 OR2X1_LOC_198/a_36_216# OR2X1_LOC_532/B 0.00fF
C23351 OR2X1_LOC_604/A OR2X1_LOC_627/a_8_216# 0.06fF
C23352 OR2X1_LOC_566/Y OR2X1_LOC_578/B 0.74fF
C23353 OR2X1_LOC_235/B OR2X1_LOC_161/A 1.50fF
C23354 AND2X1_LOC_139/B OR2X1_LOC_59/Y 0.03fF
C23355 OR2X1_LOC_694/a_8_216# OR2X1_LOC_91/A 0.02fF
C23356 AND2X1_LOC_12/Y AND2X1_LOC_498/a_36_24# 0.01fF
C23357 OR2X1_LOC_769/B OR2X1_LOC_828/B 0.01fF
C23358 AND2X1_LOC_599/a_8_24# OR2X1_LOC_19/B 0.02fF
C23359 AND2X1_LOC_302/a_36_24# OR2X1_LOC_426/B 0.01fF
C23360 OR2X1_LOC_653/Y AND2X1_LOC_58/a_8_24# 0.03fF
C23361 AND2X1_LOC_215/Y AND2X1_LOC_852/Y 0.13fF
C23362 OR2X1_LOC_92/Y AND2X1_LOC_654/Y 0.07fF
C23363 AND2X1_LOC_658/B AND2X1_LOC_806/A 0.03fF
C23364 OR2X1_LOC_653/A OR2X1_LOC_78/A 0.04fF
C23365 AND2X1_LOC_861/B AND2X1_LOC_862/A 0.01fF
C23366 OR2X1_LOC_62/A OR2X1_LOC_622/B 0.13fF
C23367 INPUT_5 OR2X1_LOC_53/a_8_216# -0.00fF
C23368 AND2X1_LOC_12/Y OR2X1_LOC_499/B 0.04fF
C23369 AND2X1_LOC_861/B AND2X1_LOC_624/A 0.07fF
C23370 OR2X1_LOC_847/A AND2X1_LOC_618/a_8_24# 0.00fF
C23371 OR2X1_LOC_673/Y OR2X1_LOC_78/A 0.15fF
C23372 VDD AND2X1_LOC_220/Y 0.29fF
C23373 AND2X1_LOC_772/B AND2X1_LOC_361/A 0.05fF
C23374 AND2X1_LOC_717/Y OR2X1_LOC_427/A 0.03fF
C23375 D_INPUT_4 OR2X1_LOC_30/a_8_216# 0.07fF
C23376 OR2X1_LOC_329/B OR2X1_LOC_6/A 0.23fF
C23377 VDD OR2X1_LOC_564/A 0.12fF
C23378 AND2X1_LOC_211/B AND2X1_LOC_715/A 0.12fF
C23379 OR2X1_LOC_838/a_8_216# AND2X1_LOC_43/B 0.06fF
C23380 AND2X1_LOC_784/A AND2X1_LOC_514/a_8_24# 0.04fF
C23381 OR2X1_LOC_51/Y OR2X1_LOC_585/A 0.14fF
C23382 OR2X1_LOC_269/B AND2X1_LOC_437/a_8_24# 0.04fF
C23383 OR2X1_LOC_62/B AND2X1_LOC_44/Y 0.19fF
C23384 AND2X1_LOC_59/Y OR2X1_LOC_354/A 0.02fF
C23385 OR2X1_LOC_158/A OR2X1_LOC_60/a_8_216# 0.01fF
C23386 AND2X1_LOC_227/Y AND2X1_LOC_227/a_8_24# 0.01fF
C23387 VDD OR2X1_LOC_629/A 0.02fF
C23388 OR2X1_LOC_405/Y OR2X1_LOC_475/B 0.02fF
C23389 OR2X1_LOC_494/A OR2X1_LOC_417/A 0.05fF
C23390 AND2X1_LOC_549/Y AND2X1_LOC_578/A 0.02fF
C23391 OR2X1_LOC_97/A D_INPUT_0 0.00fF
C23392 AND2X1_LOC_191/B OR2X1_LOC_7/A 0.10fF
C23393 OR2X1_LOC_185/A OR2X1_LOC_811/A 0.00fF
C23394 OR2X1_LOC_375/A OR2X1_LOC_623/B 0.03fF
C23395 OR2X1_LOC_821/Y OR2X1_LOC_246/A 0.03fF
C23396 OR2X1_LOC_697/Y OR2X1_LOC_36/Y 0.00fF
C23397 OR2X1_LOC_158/A AND2X1_LOC_685/a_8_24# 0.02fF
C23398 OR2X1_LOC_814/A AND2X1_LOC_603/a_8_24# 0.02fF
C23399 AND2X1_LOC_207/a_36_24# OR2X1_LOC_43/A 0.00fF
C23400 OR2X1_LOC_633/a_8_216# AND2X1_LOC_8/Y 0.03fF
C23401 VDD OR2X1_LOC_279/Y 0.18fF
C23402 OR2X1_LOC_502/A OR2X1_LOC_222/A 0.03fF
C23403 OR2X1_LOC_529/Y OR2X1_LOC_59/Y 0.04fF
C23404 OR2X1_LOC_744/A AND2X1_LOC_638/a_36_24# 0.00fF
C23405 OR2X1_LOC_780/B AND2X1_LOC_44/Y 0.32fF
C23406 AND2X1_LOC_859/B AND2X1_LOC_244/A 0.00fF
C23407 GATE_366 OR2X1_LOC_92/Y 0.03fF
C23408 OR2X1_LOC_76/B OR2X1_LOC_553/A 0.01fF
C23409 OR2X1_LOC_709/A OR2X1_LOC_447/Y 0.02fF
C23410 AND2X1_LOC_339/B D_INPUT_0 0.03fF
C23411 OR2X1_LOC_362/B OR2X1_LOC_807/A 0.25fF
C23412 OR2X1_LOC_99/B OR2X1_LOC_66/A 0.14fF
C23413 OR2X1_LOC_272/Y OR2X1_LOC_91/A 0.05fF
C23414 OR2X1_LOC_613/Y AND2X1_LOC_805/Y 0.04fF
C23415 AND2X1_LOC_228/Y AND2X1_LOC_174/a_36_24# 0.00fF
C23416 AND2X1_LOC_172/a_8_24# OR2X1_LOC_476/B 0.01fF
C23417 AND2X1_LOC_327/a_8_24# OR2X1_LOC_56/A 0.01fF
C23418 OR2X1_LOC_139/A OR2X1_LOC_786/Y 0.23fF
C23419 AND2X1_LOC_560/B OR2X1_LOC_427/A 0.01fF
C23420 OR2X1_LOC_612/a_8_216# OR2X1_LOC_62/B 0.01fF
C23421 OR2X1_LOC_833/B OR2X1_LOC_203/Y 0.45fF
C23422 AND2X1_LOC_586/a_8_24# AND2X1_LOC_56/B 0.04fF
C23423 OR2X1_LOC_600/A OR2X1_LOC_62/B 0.03fF
C23424 OR2X1_LOC_109/Y AND2X1_LOC_840/B 0.05fF
C23425 OR2X1_LOC_175/Y OR2X1_LOC_214/B 0.02fF
C23426 OR2X1_LOC_135/Y AND2X1_LOC_649/Y 0.02fF
C23427 OR2X1_LOC_499/B AND2X1_LOC_496/a_8_24# 0.01fF
C23428 INPUT_5 OR2X1_LOC_47/a_8_216# 0.09fF
C23429 OR2X1_LOC_603/a_36_216# AND2X1_LOC_452/Y 0.01fF
C23430 OR2X1_LOC_630/a_8_216# OR2X1_LOC_631/B 0.01fF
C23431 OR2X1_LOC_287/B OR2X1_LOC_814/a_8_216# 0.01fF
C23432 VDD AND2X1_LOC_165/a_8_24# 0.00fF
C23433 OR2X1_LOC_62/A OR2X1_LOC_9/a_8_216# 0.06fF
C23434 AND2X1_LOC_35/a_8_24# AND2X1_LOC_35/Y 0.00fF
C23435 AND2X1_LOC_359/B OR2X1_LOC_18/Y 0.14fF
C23436 AND2X1_LOC_851/A OR2X1_LOC_238/Y 0.01fF
C23437 AND2X1_LOC_76/Y OR2X1_LOC_52/B 0.02fF
C23438 OR2X1_LOC_235/B AND2X1_LOC_51/Y 0.03fF
C23439 OR2X1_LOC_649/B OR2X1_LOC_185/A 0.01fF
C23440 OR2X1_LOC_703/Y OR2X1_LOC_724/A 0.01fF
C23441 AND2X1_LOC_392/a_8_24# OR2X1_LOC_64/Y 0.01fF
C23442 OR2X1_LOC_664/a_8_216# OR2X1_LOC_631/B 0.03fF
C23443 AND2X1_LOC_12/Y OR2X1_LOC_391/B 0.76fF
C23444 VDD AND2X1_LOC_196/Y 0.01fF
C23445 AND2X1_LOC_541/Y AND2X1_LOC_227/Y 0.52fF
C23446 OR2X1_LOC_510/Y OR2X1_LOC_87/A 0.03fF
C23447 OR2X1_LOC_70/a_8_216# OR2X1_LOC_581/Y 0.40fF
C23448 OR2X1_LOC_138/a_8_216# OR2X1_LOC_801/B 0.04fF
C23449 AND2X1_LOC_44/Y AND2X1_LOC_39/Y 0.03fF
C23450 OR2X1_LOC_799/A OR2X1_LOC_592/a_8_216# 0.01fF
C23451 OR2X1_LOC_691/Y OR2X1_LOC_214/B 0.03fF
C23452 AND2X1_LOC_76/a_8_24# OR2X1_LOC_74/A 0.02fF
C23453 VDD OR2X1_LOC_446/Y 0.23fF
C23454 OR2X1_LOC_753/A OR2X1_LOC_39/A 0.03fF
C23455 AND2X1_LOC_605/Y AND2X1_LOC_712/B 0.00fF
C23456 OR2X1_LOC_358/A OR2X1_LOC_174/a_36_216# 0.00fF
C23457 OR2X1_LOC_377/A OR2X1_LOC_646/A 0.03fF
C23458 OR2X1_LOC_31/Y AND2X1_LOC_447/Y 0.04fF
C23459 OR2X1_LOC_6/B AND2X1_LOC_14/a_8_24# 0.03fF
C23460 OR2X1_LOC_671/a_8_216# D_INPUT_2 0.03fF
C23461 OR2X1_LOC_287/A OR2X1_LOC_532/B 0.03fF
C23462 OR2X1_LOC_3/Y OR2X1_LOC_45/a_8_216# 0.01fF
C23463 OR2X1_LOC_3/Y AND2X1_LOC_403/B 0.03fF
C23464 OR2X1_LOC_827/a_8_216# OR2X1_LOC_42/a_8_216# 0.47fF
C23465 OR2X1_LOC_858/A AND2X1_LOC_47/Y 0.03fF
C23466 OR2X1_LOC_31/Y OR2X1_LOC_380/Y 0.03fF
C23467 OR2X1_LOC_810/A OR2X1_LOC_87/A 0.07fF
C23468 OR2X1_LOC_402/a_36_216# OR2X1_LOC_402/Y -0.00fF
C23469 OR2X1_LOC_306/Y AND2X1_LOC_512/a_36_24# 0.01fF
C23470 OR2X1_LOC_702/A OR2X1_LOC_539/Y 0.00fF
C23471 AND2X1_LOC_663/B OR2X1_LOC_278/Y 0.05fF
C23472 OR2X1_LOC_107/a_8_216# AND2X1_LOC_227/Y 0.01fF
C23473 OR2X1_LOC_64/Y OR2X1_LOC_427/A 0.16fF
C23474 AND2X1_LOC_865/A OR2X1_LOC_95/Y 0.07fF
C23475 VDD OR2X1_LOC_473/A 0.07fF
C23476 OR2X1_LOC_174/A OR2X1_LOC_532/B 0.01fF
C23477 OR2X1_LOC_121/B AND2X1_LOC_492/a_8_24# 0.01fF
C23478 AND2X1_LOC_70/Y OR2X1_LOC_276/a_8_216# 0.01fF
C23479 OR2X1_LOC_70/Y AND2X1_LOC_436/B 0.11fF
C23480 OR2X1_LOC_160/A AND2X1_LOC_67/Y 0.39fF
C23481 AND2X1_LOC_741/Y AND2X1_LOC_222/Y 0.01fF
C23482 OR2X1_LOC_663/A OR2X1_LOC_244/A 0.07fF
C23483 OR2X1_LOC_404/Y OR2X1_LOC_624/A 0.03fF
C23484 OR2X1_LOC_435/a_8_216# OR2X1_LOC_532/B 0.02fF
C23485 AND2X1_LOC_702/Y OR2X1_LOC_299/a_36_216# 0.00fF
C23486 OR2X1_LOC_631/B OR2X1_LOC_296/a_8_216# 0.01fF
C23487 OR2X1_LOC_83/A OR2X1_LOC_240/A 0.03fF
C23488 OR2X1_LOC_3/Y OR2X1_LOC_44/Y 2.83fF
C23489 AND2X1_LOC_675/Y OR2X1_LOC_674/Y 0.15fF
C23490 AND2X1_LOC_118/a_8_24# OR2X1_LOC_633/B 0.01fF
C23491 AND2X1_LOC_476/A AND2X1_LOC_222/a_36_24# 0.01fF
C23492 OR2X1_LOC_631/a_36_216# OR2X1_LOC_62/B 0.00fF
C23493 OR2X1_LOC_40/Y AND2X1_LOC_848/A 0.01fF
C23494 AND2X1_LOC_12/Y OR2X1_LOC_772/Y 0.05fF
C23495 OR2X1_LOC_798/Y OR2X1_LOC_436/Y 0.01fF
C23496 AND2X1_LOC_12/Y OR2X1_LOC_846/A 0.05fF
C23497 OR2X1_LOC_62/B OR2X1_LOC_619/Y 0.03fF
C23498 AND2X1_LOC_803/B AND2X1_LOC_797/B 0.01fF
C23499 OR2X1_LOC_757/A AND2X1_LOC_620/Y 0.03fF
C23500 AND2X1_LOC_70/Y OR2X1_LOC_84/Y 0.00fF
C23501 OR2X1_LOC_405/A OR2X1_LOC_814/A 0.01fF
C23502 OR2X1_LOC_863/B OR2X1_LOC_269/B 0.01fF
C23503 OR2X1_LOC_485/A OR2X1_LOC_238/Y 0.03fF
C23504 OR2X1_LOC_696/Y OR2X1_LOC_36/Y 0.03fF
C23505 AND2X1_LOC_290/a_8_24# D_INPUT_0 0.02fF
C23506 AND2X1_LOC_530/a_8_24# OR2X1_LOC_80/A 0.05fF
C23507 AND2X1_LOC_482/a_8_24# OR2X1_LOC_532/B 0.06fF
C23508 AND2X1_LOC_326/A OR2X1_LOC_36/Y 0.01fF
C23509 AND2X1_LOC_40/Y AND2X1_LOC_441/a_36_24# 0.01fF
C23510 AND2X1_LOC_393/a_8_24# AND2X1_LOC_51/Y 0.01fF
C23511 OR2X1_LOC_316/Y OR2X1_LOC_46/A 0.00fF
C23512 AND2X1_LOC_729/Y OR2X1_LOC_22/Y 0.07fF
C23513 OR2X1_LOC_154/A OR2X1_LOC_474/a_8_216# 0.07fF
C23514 OR2X1_LOC_73/a_8_216# OR2X1_LOC_74/A 0.02fF
C23515 OR2X1_LOC_427/A OR2X1_LOC_417/A 0.17fF
C23516 AND2X1_LOC_633/Y AND2X1_LOC_633/a_8_24# 0.00fF
C23517 OR2X1_LOC_641/A OR2X1_LOC_641/B 0.25fF
C23518 OR2X1_LOC_494/a_8_216# OR2X1_LOC_47/Y 0.01fF
C23519 OR2X1_LOC_524/Y AND2X1_LOC_803/a_36_24# 0.09fF
C23520 OR2X1_LOC_596/A OR2X1_LOC_724/A 0.08fF
C23521 AND2X1_LOC_140/a_8_24# OR2X1_LOC_89/A 0.00fF
C23522 VDD D_GATE_579 0.06fF
C23523 OR2X1_LOC_154/A OR2X1_LOC_859/A 0.00fF
C23524 OR2X1_LOC_858/A OR2X1_LOC_598/A 0.07fF
C23525 OR2X1_LOC_109/Y OR2X1_LOC_31/Y 0.02fF
C23526 AND2X1_LOC_354/B OR2X1_LOC_46/A 0.15fF
C23527 AND2X1_LOC_8/Y AND2X1_LOC_46/a_36_24# 0.01fF
C23528 VDD OR2X1_LOC_228/Y 0.62fF
C23529 OR2X1_LOC_529/a_8_216# AND2X1_LOC_227/Y 0.01fF
C23530 AND2X1_LOC_563/A AND2X1_LOC_657/A 0.07fF
C23531 AND2X1_LOC_18/Y OR2X1_LOC_789/A 0.03fF
C23532 AND2X1_LOC_784/A OR2X1_LOC_22/Y 0.03fF
C23533 OR2X1_LOC_625/Y D_INPUT_3 0.07fF
C23534 AND2X1_LOC_672/B OR2X1_LOC_753/A 0.04fF
C23535 AND2X1_LOC_2/Y AND2X1_LOC_429/a_8_24# 0.01fF
C23536 OR2X1_LOC_161/B OR2X1_LOC_544/B 0.02fF
C23537 OR2X1_LOC_323/A OR2X1_LOC_696/A 0.15fF
C23538 OR2X1_LOC_417/A AND2X1_LOC_464/a_8_24# 0.04fF
C23539 VDD OR2X1_LOC_513/Y 0.18fF
C23540 OR2X1_LOC_276/B OR2X1_LOC_161/A 0.02fF
C23541 AND2X1_LOC_363/A OR2X1_LOC_417/A 0.01fF
C23542 OR2X1_LOC_497/Y OR2X1_LOC_95/Y 0.06fF
C23543 OR2X1_LOC_808/B OR2X1_LOC_170/Y 0.02fF
C23544 OR2X1_LOC_151/A OR2X1_LOC_174/Y 0.10fF
C23545 AND2X1_LOC_64/Y OR2X1_LOC_828/Y 0.05fF
C23546 OR2X1_LOC_625/Y AND2X1_LOC_483/Y 0.04fF
C23547 OR2X1_LOC_847/a_8_216# D_INPUT_1 0.02fF
C23548 OR2X1_LOC_19/B AND2X1_LOC_663/B 0.01fF
C23549 AND2X1_LOC_456/B AND2X1_LOC_657/A 0.00fF
C23550 AND2X1_LOC_736/Y AND2X1_LOC_222/Y 0.03fF
C23551 AND2X1_LOC_56/B OR2X1_LOC_269/Y 0.01fF
C23552 AND2X1_LOC_798/a_8_24# AND2X1_LOC_802/Y 0.04fF
C23553 AND2X1_LOC_65/a_36_24# OR2X1_LOC_68/B -0.00fF
C23554 OR2X1_LOC_64/Y AND2X1_LOC_687/B 0.03fF
C23555 AND2X1_LOC_56/B AND2X1_LOC_420/a_36_24# 0.01fF
C23556 AND2X1_LOC_43/B OR2X1_LOC_493/Y 0.09fF
C23557 OR2X1_LOC_83/A OR2X1_LOC_47/Y 0.07fF
C23558 OR2X1_LOC_49/A OR2X1_LOC_415/Y 0.14fF
C23559 AND2X1_LOC_474/A OR2X1_LOC_437/A 0.03fF
C23560 AND2X1_LOC_64/Y AND2X1_LOC_534/a_8_24# 0.00fF
C23561 AND2X1_LOC_640/Y AND2X1_LOC_476/A 0.21fF
C23562 AND2X1_LOC_462/B OR2X1_LOC_44/Y 0.80fF
C23563 OR2X1_LOC_559/B OR2X1_LOC_559/a_8_216# 0.50fF
C23564 OR2X1_LOC_26/Y AND2X1_LOC_721/A 0.04fF
C23565 OR2X1_LOC_415/A D_INPUT_0 0.01fF
C23566 AND2X1_LOC_102/a_8_24# D_INPUT_1 0.01fF
C23567 OR2X1_LOC_656/B OR2X1_LOC_68/B 0.24fF
C23568 OR2X1_LOC_161/A AND2X1_LOC_430/B 0.00fF
C23569 OR2X1_LOC_529/Y OR2X1_LOC_184/Y 0.39fF
C23570 OR2X1_LOC_161/A OR2X1_LOC_779/B 0.01fF
C23571 OR2X1_LOC_675/A OR2X1_LOC_440/A 0.42fF
C23572 D_INPUT_2 OR2X1_LOC_8/a_36_216# 0.03fF
C23573 OR2X1_LOC_45/B AND2X1_LOC_785/Y 0.01fF
C23574 OR2X1_LOC_62/B OR2X1_LOC_720/B 0.03fF
C23575 AND2X1_LOC_733/a_8_24# OR2X1_LOC_437/A 0.04fF
C23576 AND2X1_LOC_844/a_8_24# OR2X1_LOC_95/Y 0.01fF
C23577 AND2X1_LOC_349/B AND2X1_LOC_721/A 0.10fF
C23578 AND2X1_LOC_721/A OR2X1_LOC_89/A 0.03fF
C23579 AND2X1_LOC_92/Y AND2X1_LOC_36/Y 0.08fF
C23580 OR2X1_LOC_59/Y AND2X1_LOC_791/a_8_24# 0.02fF
C23581 AND2X1_LOC_104/a_8_24# OR2X1_LOC_80/A 0.04fF
C23582 OR2X1_LOC_97/A AND2X1_LOC_438/a_8_24# 0.02fF
C23583 OR2X1_LOC_820/A AND2X1_LOC_789/Y 0.17fF
C23584 AND2X1_LOC_12/Y OR2X1_LOC_348/B 0.12fF
C23585 OR2X1_LOC_92/Y OR2X1_LOC_13/B 0.87fF
C23586 AND2X1_LOC_64/Y AND2X1_LOC_110/Y 0.39fF
C23587 OR2X1_LOC_458/B OR2X1_LOC_723/B 0.03fF
C23588 OR2X1_LOC_641/A OR2X1_LOC_227/A 0.02fF
C23589 OR2X1_LOC_471/Y OR2X1_LOC_477/a_8_216# 0.07fF
C23590 AND2X1_LOC_858/B OR2X1_LOC_504/a_36_216# 0.01fF
C23591 AND2X1_LOC_476/A OR2X1_LOC_416/Y 0.03fF
C23592 OR2X1_LOC_756/B OR2X1_LOC_374/a_36_216# 0.00fF
C23593 OR2X1_LOC_632/Y OR2X1_LOC_500/a_8_216# 0.02fF
C23594 OR2X1_LOC_623/B OR2X1_LOC_515/Y 0.72fF
C23595 OR2X1_LOC_553/A OR2X1_LOC_578/B 0.07fF
C23596 AND2X1_LOC_64/Y AND2X1_LOC_313/a_36_24# 0.00fF
C23597 AND2X1_LOC_91/B AND2X1_LOC_313/a_8_24# 0.01fF
C23598 OR2X1_LOC_724/a_36_216# OR2X1_LOC_317/B 0.00fF
C23599 OR2X1_LOC_211/a_8_216# OR2X1_LOC_303/B 0.01fF
C23600 OR2X1_LOC_661/A AND2X1_LOC_7/B 0.01fF
C23601 VDD OR2X1_LOC_562/A 0.28fF
C23602 OR2X1_LOC_175/Y OR2X1_LOC_325/B 0.15fF
C23603 AND2X1_LOC_566/B OR2X1_LOC_428/A 0.03fF
C23604 OR2X1_LOC_841/a_8_216# OR2X1_LOC_593/B 0.03fF
C23605 AND2X1_LOC_95/Y OR2X1_LOC_501/a_36_216# 0.00fF
C23606 OR2X1_LOC_40/Y AND2X1_LOC_804/A 0.02fF
C23607 OR2X1_LOC_203/a_8_216# OR2X1_LOC_269/A 0.03fF
C23608 OR2X1_LOC_725/B OR2X1_LOC_712/B 0.00fF
C23609 VDD OR2X1_LOC_321/a_8_216# 0.00fF
C23610 AND2X1_LOC_95/Y OR2X1_LOC_730/B 0.20fF
C23611 AND2X1_LOC_785/A OR2X1_LOC_164/Y 0.20fF
C23612 OR2X1_LOC_185/A OR2X1_LOC_777/B 0.03fF
C23613 OR2X1_LOC_65/B OR2X1_LOC_13/B 0.03fF
C23614 OR2X1_LOC_471/Y OR2X1_LOC_223/A 0.03fF
C23615 AND2X1_LOC_170/B AND2X1_LOC_864/a_8_24# 0.01fF
C23616 OR2X1_LOC_632/a_8_216# OR2X1_LOC_115/B 0.01fF
C23617 OR2X1_LOC_632/a_36_216# OR2X1_LOC_140/B 0.00fF
C23618 OR2X1_LOC_653/Y OR2X1_LOC_539/B 0.02fF
C23619 OR2X1_LOC_53/Y AND2X1_LOC_691/a_8_24# 0.01fF
C23620 AND2X1_LOC_303/A OR2X1_LOC_300/a_8_216# 0.47fF
C23621 AND2X1_LOC_101/a_8_24# OR2X1_LOC_813/Y 0.01fF
C23622 AND2X1_LOC_717/B AND2X1_LOC_657/A 0.39fF
C23623 OR2X1_LOC_600/A OR2X1_LOC_15/a_36_216# 0.01fF
C23624 OR2X1_LOC_85/A OR2X1_LOC_437/A 0.01fF
C23625 OR2X1_LOC_750/a_8_216# OR2X1_LOC_214/B 0.12fF
C23626 AND2X1_LOC_22/Y OR2X1_LOC_648/A 0.10fF
C23627 OR2X1_LOC_89/A AND2X1_LOC_217/a_8_24# 0.01fF
C23628 AND2X1_LOC_358/Y OR2X1_LOC_426/B 0.05fF
C23629 AND2X1_LOC_555/Y AND2X1_LOC_347/Y 0.02fF
C23630 AND2X1_LOC_191/B OR2X1_LOC_753/a_8_216# 0.05fF
C23631 OR2X1_LOC_185/A AND2X1_LOC_591/a_36_24# 0.00fF
C23632 AND2X1_LOC_339/B AND2X1_LOC_326/B 0.00fF
C23633 AND2X1_LOC_850/A AND2X1_LOC_242/B 0.01fF
C23634 AND2X1_LOC_51/Y OR2X1_LOC_779/B 0.08fF
C23635 OR2X1_LOC_56/A OR2X1_LOC_16/A 0.17fF
C23636 OR2X1_LOC_335/Y OR2X1_LOC_97/A 0.02fF
C23637 OR2X1_LOC_135/a_8_216# OR2X1_LOC_59/Y 0.08fF
C23638 AND2X1_LOC_57/Y AND2X1_LOC_95/Y 0.04fF
C23639 OR2X1_LOC_471/Y OR2X1_LOC_705/B 0.14fF
C23640 OR2X1_LOC_427/A OR2X1_LOC_89/a_36_216# 0.02fF
C23641 AND2X1_LOC_56/B OR2X1_LOC_469/B 0.03fF
C23642 OR2X1_LOC_421/A VDD 0.63fF
C23643 OR2X1_LOC_323/A AND2X1_LOC_717/a_8_24# 0.00fF
C23644 OR2X1_LOC_114/B OR2X1_LOC_830/a_8_216# 0.05fF
C23645 AND2X1_LOC_544/Y OR2X1_LOC_427/A 0.05fF
C23646 AND2X1_LOC_391/a_8_24# OR2X1_LOC_428/A 0.01fF
C23647 OR2X1_LOC_22/Y OR2X1_LOC_88/Y 0.03fF
C23648 AND2X1_LOC_40/Y OR2X1_LOC_97/A 0.05fF
C23649 OR2X1_LOC_193/A OR2X1_LOC_193/a_8_216# 0.18fF
C23650 OR2X1_LOC_409/Y AND2X1_LOC_460/a_8_24# 0.01fF
C23651 OR2X1_LOC_185/A OR2X1_LOC_831/B 0.03fF
C23652 AND2X1_LOC_366/a_8_24# AND2X1_LOC_614/a_8_24# 0.23fF
C23653 OR2X1_LOC_22/Y OR2X1_LOC_172/Y 0.15fF
C23654 OR2X1_LOC_810/A OR2X1_LOC_579/A 0.29fF
C23655 OR2X1_LOC_68/Y AND2X1_LOC_31/Y 0.02fF
C23656 AND2X1_LOC_84/Y OR2X1_LOC_619/Y 0.03fF
C23657 AND2X1_LOC_159/a_8_24# OR2X1_LOC_844/B 0.01fF
C23658 OR2X1_LOC_108/Y OR2X1_LOC_56/A 0.29fF
C23659 OR2X1_LOC_810/A OR2X1_LOC_844/B 0.38fF
C23660 OR2X1_LOC_323/A AND2X1_LOC_458/Y 0.01fF
C23661 AND2X1_LOC_64/Y OR2X1_LOC_664/Y 0.01fF
C23662 OR2X1_LOC_66/A AND2X1_LOC_245/a_8_24# 0.05fF
C23663 OR2X1_LOC_121/B OR2X1_LOC_317/B 0.01fF
C23664 OR2X1_LOC_507/A OR2X1_LOC_78/B 0.01fF
C23665 AND2X1_LOC_505/a_36_24# OR2X1_LOC_78/A 0.00fF
C23666 OR2X1_LOC_758/Y AND2X1_LOC_759/a_8_24# 0.23fF
C23667 AND2X1_LOC_850/Y AND2X1_LOC_244/A 0.00fF
C23668 OR2X1_LOC_323/A OR2X1_LOC_271/B 0.00fF
C23669 AND2X1_LOC_47/Y AND2X1_LOC_31/Y 1.90fF
C23670 OR2X1_LOC_47/Y AND2X1_LOC_405/a_8_24# 0.01fF
C23671 AND2X1_LOC_367/A AND2X1_LOC_243/Y 0.10fF
C23672 OR2X1_LOC_662/A OR2X1_LOC_227/B 0.08fF
C23673 OR2X1_LOC_406/Y AND2X1_LOC_624/A 0.03fF
C23674 VDD OR2X1_LOC_660/Y -0.00fF
C23675 AND2X1_LOC_564/B OR2X1_LOC_680/A 0.07fF
C23676 AND2X1_LOC_754/a_8_24# OR2X1_LOC_502/A 0.01fF
C23677 OR2X1_LOC_127/a_8_216# OR2X1_LOC_428/A 0.02fF
C23678 AND2X1_LOC_711/Y AND2X1_LOC_791/a_8_24# 0.01fF
C23679 OR2X1_LOC_854/a_8_216# OR2X1_LOC_151/A 0.02fF
C23680 OR2X1_LOC_109/Y AND2X1_LOC_464/A 0.02fF
C23681 AND2X1_LOC_121/a_8_24# OR2X1_LOC_56/A 0.02fF
C23682 OR2X1_LOC_128/A AND2X1_LOC_44/Y 0.01fF
C23683 OR2X1_LOC_604/A OR2X1_LOC_697/Y 0.08fF
C23684 OR2X1_LOC_345/Y OR2X1_LOC_260/a_8_216# 0.01fF
C23685 OR2X1_LOC_810/A OR2X1_LOC_390/B 0.07fF
C23686 AND2X1_LOC_568/B AND2X1_LOC_367/A 0.03fF
C23687 OR2X1_LOC_482/Y OR2X1_LOC_495/Y 0.04fF
C23688 OR2X1_LOC_680/A OR2X1_LOC_530/a_8_216# 0.02fF
C23689 VDD AND2X1_LOC_456/B 0.58fF
C23690 OR2X1_LOC_11/Y OR2X1_LOC_18/a_36_216# 0.03fF
C23691 OR2X1_LOC_71/Y OR2X1_LOC_71/A 0.01fF
C23692 OR2X1_LOC_497/a_36_216# AND2X1_LOC_242/B 0.02fF
C23693 OR2X1_LOC_185/A OR2X1_LOC_344/A 0.02fF
C23694 OR2X1_LOC_139/A OR2X1_LOC_204/Y 0.07fF
C23695 OR2X1_LOC_32/B OR2X1_LOC_12/Y 0.01fF
C23696 AND2X1_LOC_846/a_8_24# AND2X1_LOC_793/Y 0.01fF
C23697 OR2X1_LOC_709/A OR2X1_LOC_161/A 0.03fF
C23698 OR2X1_LOC_375/A OR2X1_LOC_713/a_36_216# 0.00fF
C23699 AND2X1_LOC_715/Y OR2X1_LOC_601/Y 0.14fF
C23700 AND2X1_LOC_658/B OR2X1_LOC_441/Y 0.23fF
C23701 AND2X1_LOC_612/B OR2X1_LOC_415/Y 0.02fF
C23702 OR2X1_LOC_89/a_8_216# OR2X1_LOC_89/Y 0.01fF
C23703 AND2X1_LOC_3/Y OR2X1_LOC_115/B 0.51fF
C23704 AND2X1_LOC_716/Y AND2X1_LOC_335/Y 0.04fF
C23705 AND2X1_LOC_12/Y AND2X1_LOC_65/A 0.03fF
C23706 OR2X1_LOC_615/Y AND2X1_LOC_790/a_36_24# 0.01fF
C23707 AND2X1_LOC_565/B OR2X1_LOC_189/a_8_216# 0.04fF
C23708 OR2X1_LOC_494/Y AND2X1_LOC_348/A 0.81fF
C23709 OR2X1_LOC_187/a_8_216# AND2X1_LOC_191/B 0.01fF
C23710 OR2X1_LOC_335/A OR2X1_LOC_605/A 0.26fF
C23711 AND2X1_LOC_363/Y AND2X1_LOC_348/A 0.03fF
C23712 AND2X1_LOC_72/B OR2X1_LOC_736/a_8_216# 0.01fF
C23713 OR2X1_LOC_538/A AND2X1_LOC_311/a_36_24# 0.00fF
C23714 OR2X1_LOC_469/Y OR2X1_LOC_803/A 0.03fF
C23715 AND2X1_LOC_335/Y AND2X1_LOC_654/Y 0.01fF
C23716 AND2X1_LOC_392/A OR2X1_LOC_278/Y 0.00fF
C23717 OR2X1_LOC_449/B AND2X1_LOC_44/Y 0.03fF
C23718 OR2X1_LOC_524/Y OR2X1_LOC_441/a_8_216# 0.18fF
C23719 OR2X1_LOC_620/Y OR2X1_LOC_66/A 0.07fF
C23720 OR2X1_LOC_156/A OR2X1_LOC_160/A 0.30fF
C23721 AND2X1_LOC_596/a_36_24# OR2X1_LOC_48/B 0.01fF
C23722 OR2X1_LOC_505/a_36_216# AND2X1_LOC_806/A 0.00fF
C23723 AND2X1_LOC_392/A AND2X1_LOC_662/B 0.05fF
C23724 D_GATE_662 OR2X1_LOC_848/A 0.02fF
C23725 AND2X1_LOC_849/a_36_24# OR2X1_LOC_13/B 0.01fF
C23726 AND2X1_LOC_721/a_8_24# OR2X1_LOC_59/Y 0.01fF
C23727 OR2X1_LOC_426/B OR2X1_LOC_427/Y 0.00fF
C23728 AND2X1_LOC_211/B OR2X1_LOC_310/a_36_216# 0.00fF
C23729 OR2X1_LOC_51/Y AND2X1_LOC_833/a_36_24# 0.00fF
C23730 AND2X1_LOC_596/a_36_24# OR2X1_LOC_18/Y 0.00fF
C23731 OR2X1_LOC_294/Y OR2X1_LOC_269/B 0.03fF
C23732 OR2X1_LOC_860/a_36_216# OR2X1_LOC_244/Y 0.03fF
C23733 D_INPUT_1 OR2X1_LOC_71/A 0.26fF
C23734 AND2X1_LOC_31/Y OR2X1_LOC_598/A 0.03fF
C23735 AND2X1_LOC_729/Y OR2X1_LOC_485/Y 0.39fF
C23736 AND2X1_LOC_339/Y AND2X1_LOC_339/a_36_24# 0.00fF
C23737 AND2X1_LOC_84/Y AND2X1_LOC_201/a_8_24# 0.01fF
C23738 AND2X1_LOC_31/Y OR2X1_LOC_717/a_36_216# 0.00fF
C23739 OR2X1_LOC_36/Y AND2X1_LOC_476/Y 0.01fF
C23740 OR2X1_LOC_45/B OR2X1_LOC_3/Y 3.80fF
C23741 OR2X1_LOC_507/A OR2X1_LOC_375/A 0.03fF
C23742 OR2X1_LOC_653/Y OR2X1_LOC_78/B 0.16fF
C23743 AND2X1_LOC_394/a_8_24# AND2X1_LOC_18/Y 0.01fF
C23744 OR2X1_LOC_715/B OR2X1_LOC_87/A 0.10fF
C23745 AND2X1_LOC_358/Y OR2X1_LOC_743/A 0.03fF
C23746 AND2X1_LOC_70/Y OR2X1_LOC_161/A 0.86fF
C23747 AND2X1_LOC_486/Y AND2X1_LOC_556/a_8_24# 0.06fF
C23748 OR2X1_LOC_756/B AND2X1_LOC_125/a_8_24# 0.11fF
C23749 OR2X1_LOC_158/A AND2X1_LOC_818/a_36_24# 0.00fF
C23750 OR2X1_LOC_312/Y OR2X1_LOC_322/a_36_216# 0.00fF
C23751 AND2X1_LOC_366/A OR2X1_LOC_278/Y 0.03fF
C23752 OR2X1_LOC_584/Y OR2X1_LOC_52/B 0.23fF
C23753 AND2X1_LOC_486/Y OR2X1_LOC_516/B 1.11fF
C23754 OR2X1_LOC_154/A OR2X1_LOC_66/A 1.06fF
C23755 OR2X1_LOC_160/A OR2X1_LOC_520/a_8_216# 0.05fF
C23756 OR2X1_LOC_864/A OR2X1_LOC_6/B 0.07fF
C23757 GATE_366 OR2X1_LOC_600/A 0.03fF
C23758 OR2X1_LOC_493/Y OR2X1_LOC_558/A 0.08fF
C23759 AND2X1_LOC_565/B AND2X1_LOC_565/Y 0.21fF
C23760 OR2X1_LOC_691/Y OR2X1_LOC_193/A 0.02fF
C23761 OR2X1_LOC_733/A OR2X1_LOC_269/B 0.14fF
C23762 OR2X1_LOC_62/B OR2X1_LOC_554/a_8_216# 0.01fF
C23763 AND2X1_LOC_91/B AND2X1_LOC_494/a_8_24# 0.05fF
C23764 OR2X1_LOC_3/Y OR2X1_LOC_382/A 0.17fF
C23765 AND2X1_LOC_70/Y AND2X1_LOC_25/Y 0.11fF
C23766 OR2X1_LOC_417/a_8_216# AND2X1_LOC_212/Y -0.01fF
C23767 OR2X1_LOC_494/a_8_216# OR2X1_LOC_625/Y 0.01fF
C23768 AND2X1_LOC_654/B OR2X1_LOC_586/Y 0.07fF
C23769 OR2X1_LOC_748/A OR2X1_LOC_261/a_8_216# 0.01fF
C23770 OR2X1_LOC_676/a_8_216# OR2X1_LOC_155/A 0.04fF
C23771 OR2X1_LOC_151/A AND2X1_LOC_42/B 0.07fF
C23772 OR2X1_LOC_121/B AND2X1_LOC_44/Y 0.18fF
C23773 OR2X1_LOC_6/B OR2X1_LOC_633/B 0.05fF
C23774 OR2X1_LOC_703/A OR2X1_LOC_161/A 0.20fF
C23775 VDD AND2X1_LOC_856/A 0.21fF
C23776 AND2X1_LOC_180/a_36_24# OR2X1_LOC_74/A 0.01fF
C23777 OR2X1_LOC_637/Y OR2X1_LOC_828/B 0.01fF
C23778 OR2X1_LOC_803/a_36_216# OR2X1_LOC_803/B 0.00fF
C23779 AND2X1_LOC_566/B AND2X1_LOC_211/a_8_24# 0.01fF
C23780 OR2X1_LOC_312/Y OR2X1_LOC_600/A 0.03fF
C23781 OR2X1_LOC_90/a_36_216# OR2X1_LOC_85/A 0.01fF
C23782 OR2X1_LOC_624/A OR2X1_LOC_474/Y 0.15fF
C23783 OR2X1_LOC_709/A AND2X1_LOC_51/Y 0.05fF
C23784 OR2X1_LOC_490/Y AND2X1_LOC_243/Y 0.00fF
C23785 OR2X1_LOC_185/A OR2X1_LOC_254/A 0.01fF
C23786 AND2X1_LOC_734/Y AND2X1_LOC_807/Y 0.09fF
C23787 OR2X1_LOC_74/A AND2X1_LOC_243/Y 0.01fF
C23788 OR2X1_LOC_128/B OR2X1_LOC_736/A 0.03fF
C23789 VDD OR2X1_LOC_287/B 0.91fF
C23790 OR2X1_LOC_175/Y D_INPUT_0 0.03fF
C23791 AND2X1_LOC_802/a_8_24# AND2X1_LOC_810/B 0.01fF
C23792 VDD OR2X1_LOC_453/A -0.00fF
C23793 AND2X1_LOC_358/Y OR2X1_LOC_246/A 0.03fF
C23794 AND2X1_LOC_392/A AND2X1_LOC_337/B 0.01fF
C23795 OR2X1_LOC_329/B OR2X1_LOC_44/Y 1.24fF
C23796 VDD AND2X1_LOC_717/B 0.19fF
C23797 OR2X1_LOC_137/a_8_216# OR2X1_LOC_673/Y 0.01fF
C23798 OR2X1_LOC_768/A OR2X1_LOC_849/A 0.02fF
C23799 OR2X1_LOC_748/A OR2X1_LOC_297/A 0.02fF
C23800 AND2X1_LOC_633/Y AND2X1_LOC_219/A 0.16fF
C23801 OR2X1_LOC_65/B AND2X1_LOC_266/a_8_24# 0.01fF
C23802 OR2X1_LOC_532/B OR2X1_LOC_563/A 0.07fF
C23803 OR2X1_LOC_798/Y OR2X1_LOC_799/a_8_216# 0.48fF
C23804 OR2X1_LOC_802/a_8_216# OR2X1_LOC_539/Y 0.05fF
C23805 OR2X1_LOC_634/A AND2X1_LOC_89/a_8_24# 0.17fF
C23806 AND2X1_LOC_161/a_8_24# OR2X1_LOC_427/A 0.06fF
C23807 AND2X1_LOC_178/a_8_24# OR2X1_LOC_181/B 0.02fF
C23808 AND2X1_LOC_654/Y OR2X1_LOC_619/Y 1.45fF
C23809 AND2X1_LOC_550/A OR2X1_LOC_427/A 0.62fF
C23810 AND2X1_LOC_513/a_8_24# AND2X1_LOC_840/B 0.11fF
C23811 OR2X1_LOC_691/Y D_INPUT_0 0.03fF
C23812 AND2X1_LOC_665/a_8_24# OR2X1_LOC_563/A 0.02fF
C23813 OR2X1_LOC_405/A OR2X1_LOC_317/A 0.01fF
C23814 D_INPUT_0 AND2X1_LOC_219/A 0.06fF
C23815 OR2X1_LOC_646/A OR2X1_LOC_78/B 0.01fF
C23816 OR2X1_LOC_516/A AND2X1_LOC_787/a_8_24# 0.01fF
C23817 OR2X1_LOC_589/A OR2X1_LOC_245/a_36_216# 0.00fF
C23818 AND2X1_LOC_56/B OR2X1_LOC_274/Y 0.18fF
C23819 OR2X1_LOC_753/A AND2X1_LOC_240/a_8_24# 0.01fF
C23820 OR2X1_LOC_604/A OR2X1_LOC_696/Y 0.02fF
C23821 AND2X1_LOC_735/Y AND2X1_LOC_474/Y 0.22fF
C23822 OR2X1_LOC_647/Y AND2X1_LOC_18/Y 0.10fF
C23823 OR2X1_LOC_502/A OR2X1_LOC_468/Y 0.03fF
C23824 OR2X1_LOC_9/Y OR2X1_LOC_54/Y 3.68fF
C23825 OR2X1_LOC_251/Y AND2X1_LOC_456/B 0.02fF
C23826 D_INPUT_0 OR2X1_LOC_713/A -0.01fF
C23827 AND2X1_LOC_380/a_8_24# OR2X1_LOC_460/B 0.01fF
C23828 AND2X1_LOC_543/a_8_24# OR2X1_LOC_312/Y 0.01fF
C23829 OR2X1_LOC_32/B OR2X1_LOC_393/Y 0.13fF
C23830 OR2X1_LOC_756/B OR2X1_LOC_593/A 0.01fF
C23831 OR2X1_LOC_329/B AND2X1_LOC_116/Y 0.01fF
C23832 VDD OR2X1_LOC_825/Y -0.00fF
C23833 AND2X1_LOC_535/Y OR2X1_LOC_311/Y 0.00fF
C23834 VDD OR2X1_LOC_76/A 0.02fF
C23835 AND2X1_LOC_605/Y OR2X1_LOC_89/A 0.01fF
C23836 OR2X1_LOC_532/B OR2X1_LOC_355/a_36_216# 0.00fF
C23837 AND2X1_LOC_70/Y AND2X1_LOC_51/Y 12.67fF
C23838 OR2X1_LOC_3/Y OR2X1_LOC_292/a_8_216# 0.01fF
C23839 AND2X1_LOC_12/Y AND2X1_LOC_381/a_8_24# 0.01fF
C23840 AND2X1_LOC_732/a_8_24# OR2X1_LOC_64/Y 0.01fF
C23841 OR2X1_LOC_481/A OR2X1_LOC_59/Y 0.37fF
C23842 OR2X1_LOC_502/A AND2X1_LOC_696/a_36_24# 0.01fF
C23843 OR2X1_LOC_314/Y AND2X1_LOC_452/Y 0.11fF
C23844 OR2X1_LOC_744/A AND2X1_LOC_798/Y 0.23fF
C23845 AND2X1_LOC_729/Y OR2X1_LOC_39/A 0.05fF
C23846 AND2X1_LOC_737/Y OR2X1_LOC_52/B 0.03fF
C23847 OR2X1_LOC_641/Y OR2X1_LOC_520/B 0.30fF
C23848 INPUT_3 AND2X1_LOC_852/a_8_24# 0.01fF
C23849 OR2X1_LOC_176/Y AND2X1_LOC_810/a_8_24# 0.01fF
C23850 AND2X1_LOC_753/a_8_24# OR2X1_LOC_269/B 0.06fF
C23851 OR2X1_LOC_36/Y OR2X1_LOC_595/a_8_216# 0.14fF
C23852 VDD OR2X1_LOC_835/Y 0.04fF
C23853 OR2X1_LOC_87/A OR2X1_LOC_215/Y 0.02fF
C23854 AND2X1_LOC_753/B AND2X1_LOC_387/B 0.07fF
C23855 AND2X1_LOC_593/a_8_24# OR2X1_LOC_31/Y 0.01fF
C23856 OR2X1_LOC_87/A AND2X1_LOC_230/a_36_24# 0.01fF
C23857 OR2X1_LOC_251/Y OR2X1_LOC_250/a_36_216# 0.01fF
C23858 VDD OR2X1_LOC_148/A 0.21fF
C23859 OR2X1_LOC_703/A AND2X1_LOC_51/Y 0.03fF
C23860 AND2X1_LOC_20/a_8_24# OR2X1_LOC_750/A 0.20fF
C23861 INPUT_0 OR2X1_LOC_416/Y 0.08fF
C23862 OR2X1_LOC_733/a_8_216# OR2X1_LOC_733/B 0.00fF
C23863 AND2X1_LOC_793/Y GATE_579 0.00fF
C23864 AND2X1_LOC_784/A OR2X1_LOC_39/A 0.10fF
C23865 OR2X1_LOC_479/Y OR2X1_LOC_785/B 0.02fF
C23866 OR2X1_LOC_312/Y OR2X1_LOC_619/Y 0.07fF
C23867 OR2X1_LOC_744/A OR2X1_LOC_46/A 0.15fF
C23868 OR2X1_LOC_463/a_8_216# OR2X1_LOC_375/A 0.06fF
C23869 OR2X1_LOC_352/a_8_216# OR2X1_LOC_365/B 0.01fF
C23870 OR2X1_LOC_640/a_8_216# AND2X1_LOC_8/Y 0.01fF
C23871 AND2X1_LOC_31/Y OR2X1_LOC_186/a_8_216# 0.01fF
C23872 OR2X1_LOC_475/Y OR2X1_LOC_475/B 0.01fF
C23873 AND2X1_LOC_755/a_8_24# OR2X1_LOC_287/B 0.00fF
C23874 OR2X1_LOC_124/A D_INPUT_0 0.01fF
C23875 OR2X1_LOC_194/Y OR2X1_LOC_200/a_8_216# 0.06fF
C23876 AND2X1_LOC_569/A AND2X1_LOC_580/A 0.00fF
C23877 VDD OR2X1_LOC_436/Y 0.19fF
C23878 AND2X1_LOC_554/Y AND2X1_LOC_489/Y 0.14fF
C23879 OR2X1_LOC_517/A OR2X1_LOC_245/a_8_216# 0.03fF
C23880 OR2X1_LOC_85/A OR2X1_LOC_753/A 0.05fF
C23881 AND2X1_LOC_14/a_36_24# INPUT_1 0.00fF
C23882 OR2X1_LOC_112/A OR2X1_LOC_175/a_8_216# -0.00fF
C23883 OR2X1_LOC_6/B OR2X1_LOC_47/Y 0.07fF
C23884 AND2X1_LOC_354/B AND2X1_LOC_854/a_8_24# 0.04fF
C23885 AND2X1_LOC_17/Y AND2X1_LOC_25/Y 0.13fF
C23886 OR2X1_LOC_748/A OR2X1_LOC_43/A 0.01fF
C23887 OR2X1_LOC_479/Y OR2X1_LOC_212/A 0.03fF
C23888 AND2X1_LOC_858/B OR2X1_LOC_226/a_36_216# 0.01fF
C23889 AND2X1_LOC_474/A AND2X1_LOC_845/Y 0.07fF
C23890 AND2X1_LOC_852/a_36_24# AND2X1_LOC_852/Y 0.01fF
C23891 OR2X1_LOC_364/B OR2X1_LOC_551/B 0.00fF
C23892 OR2X1_LOC_26/Y AND2X1_LOC_361/A 0.21fF
C23893 AND2X1_LOC_3/Y OR2X1_LOC_222/A 0.07fF
C23894 AND2X1_LOC_866/B OR2X1_LOC_628/Y 0.02fF
C23895 OR2X1_LOC_3/Y OR2X1_LOC_767/a_8_216# 0.02fF
C23896 AND2X1_LOC_316/a_8_24# OR2X1_LOC_814/A 0.13fF
C23897 AND2X1_LOC_359/B OR2X1_LOC_585/A 0.02fF
C23898 OR2X1_LOC_744/A AND2X1_LOC_227/Y 0.09fF
C23899 AND2X1_LOC_31/Y OR2X1_LOC_34/A 0.06fF
C23900 OR2X1_LOC_495/a_8_216# OR2X1_LOC_238/Y 0.41fF
C23901 OR2X1_LOC_485/A AND2X1_LOC_349/a_8_24# 0.01fF
C23902 AND2X1_LOC_784/A AND2X1_LOC_211/B 1.36fF
C23903 OR2X1_LOC_185/A OR2X1_LOC_456/A 0.01fF
C23904 OR2X1_LOC_419/Y AND2X1_LOC_476/Y 0.10fF
C23905 OR2X1_LOC_404/Y OR2X1_LOC_161/A 0.01fF
C23906 OR2X1_LOC_40/Y OR2X1_LOC_41/a_8_216# 0.07fF
C23907 OR2X1_LOC_440/A AND2X1_LOC_437/a_36_24# 0.00fF
C23908 OR2X1_LOC_89/A AND2X1_LOC_361/A 0.09fF
C23909 OR2X1_LOC_256/Y OR2X1_LOC_255/a_36_216# 0.01fF
C23910 OR2X1_LOC_491/Y AND2X1_LOC_717/B 0.01fF
C23911 OR2X1_LOC_280/Y AND2X1_LOC_374/Y 0.01fF
C23912 AND2X1_LOC_555/Y OR2X1_LOC_437/A 0.00fF
C23913 AND2X1_LOC_76/Y OR2X1_LOC_22/Y 0.03fF
C23914 OR2X1_LOC_119/a_36_216# OR2X1_LOC_39/A 0.00fF
C23915 AND2X1_LOC_734/Y OR2X1_LOC_95/Y 0.00fF
C23916 OR2X1_LOC_278/A AND2X1_LOC_573/A 0.33fF
C23917 OR2X1_LOC_136/Y OR2X1_LOC_437/A 0.01fF
C23918 OR2X1_LOC_431/a_8_216# OR2X1_LOC_36/Y 0.01fF
C23919 AND2X1_LOC_40/Y AND2X1_LOC_613/a_8_24# 0.04fF
C23920 OR2X1_LOC_267/Y OR2X1_LOC_140/Y 0.01fF
C23921 OR2X1_LOC_481/A OR2X1_LOC_820/B 0.04fF
C23922 OR2X1_LOC_99/A OR2X1_LOC_66/A 0.03fF
C23923 AND2X1_LOC_489/Y OR2X1_LOC_280/Y 0.14fF
C23924 OR2X1_LOC_3/Y OR2X1_LOC_261/Y 0.01fF
C23925 AND2X1_LOC_55/a_8_24# OR2X1_LOC_19/B 0.01fF
C23926 AND2X1_LOC_79/Y OR2X1_LOC_204/a_8_216# 0.01fF
C23927 OR2X1_LOC_441/Y OR2X1_LOC_47/Y 0.06fF
C23928 OR2X1_LOC_509/a_8_216# OR2X1_LOC_560/A 0.01fF
C23929 OR2X1_LOC_96/B OR2X1_LOC_54/Y 0.00fF
C23930 OR2X1_LOC_94/a_36_216# OR2X1_LOC_46/A 0.00fF
C23931 AND2X1_LOC_17/Y AND2X1_LOC_51/Y 1.81fF
C23932 OR2X1_LOC_180/a_8_216# OR2X1_LOC_578/B 0.01fF
C23933 OR2X1_LOC_427/A OR2X1_LOC_55/a_8_216# 0.02fF
C23934 OR2X1_LOC_175/Y OR2X1_LOC_339/A 0.01fF
C23935 VDD OR2X1_LOC_566/Y 0.00fF
C23936 OR2X1_LOC_471/Y OR2X1_LOC_213/A 0.80fF
C23937 AND2X1_LOC_576/Y AND2X1_LOC_574/A 0.02fF
C23938 OR2X1_LOC_137/B OR2X1_LOC_532/B 0.25fF
C23939 OR2X1_LOC_653/A OR2X1_LOC_814/A 0.00fF
C23940 AND2X1_LOC_456/B AND2X1_LOC_624/B 0.01fF
C23941 OR2X1_LOC_416/Y OR2X1_LOC_690/A 0.02fF
C23942 AND2X1_LOC_852/Y OR2X1_LOC_54/Y 0.15fF
C23943 AND2X1_LOC_185/a_36_24# AND2X1_LOC_620/Y 0.00fF
C23944 OR2X1_LOC_673/Y OR2X1_LOC_814/A 0.03fF
C23945 OR2X1_LOC_66/A OR2X1_LOC_560/A 0.03fF
C23946 OR2X1_LOC_502/A OR2X1_LOC_205/Y 0.03fF
C23947 OR2X1_LOC_66/A OR2X1_LOC_198/A 0.08fF
C23948 OR2X1_LOC_22/Y OR2X1_LOC_52/B 0.40fF
C23949 OR2X1_LOC_161/B OR2X1_LOC_217/A 0.03fF
C23950 OR2X1_LOC_703/A OR2X1_LOC_551/B 0.07fF
C23951 OR2X1_LOC_835/Y OR2X1_LOC_836/B 0.94fF
C23952 OR2X1_LOC_286/a_8_216# OR2X1_LOC_269/B 0.10fF
C23953 OR2X1_LOC_446/B OR2X1_LOC_730/A 0.02fF
C23954 AND2X1_LOC_729/Y OR2X1_LOC_760/a_8_216# 0.01fF
C23955 OR2X1_LOC_62/A OR2X1_LOC_39/A 0.00fF
C23956 OR2X1_LOC_160/A OR2X1_LOC_223/A 0.03fF
C23957 OR2X1_LOC_825/Y OR2X1_LOC_826/a_8_216# 0.41fF
C23958 OR2X1_LOC_64/Y OR2X1_LOC_681/Y 0.00fF
C23959 OR2X1_LOC_273/a_36_216# OR2X1_LOC_416/Y 0.00fF
C23960 OR2X1_LOC_404/Y AND2X1_LOC_51/Y 0.08fF
C23961 OR2X1_LOC_47/Y AND2X1_LOC_436/B 0.02fF
C23962 OR2X1_LOC_429/Y AND2X1_LOC_639/A 0.01fF
C23963 OR2X1_LOC_31/Y AND2X1_LOC_264/a_8_24# 0.01fF
C23964 OR2X1_LOC_864/A AND2X1_LOC_47/Y 0.03fF
C23965 OR2X1_LOC_208/A OR2X1_LOC_175/Y 0.04fF
C23966 OR2X1_LOC_687/Y AND2X1_LOC_681/a_8_24# 0.06fF
C23967 AND2X1_LOC_476/A OR2X1_LOC_6/A 0.07fF
C23968 OR2X1_LOC_426/B OR2X1_LOC_71/A 0.03fF
C23969 OR2X1_LOC_154/A OR2X1_LOC_84/A 0.43fF
C23970 INPUT_0 OR2X1_LOC_80/A 0.35fF
C23971 OR2X1_LOC_600/A OR2X1_LOC_13/B 0.13fF
C23972 AND2X1_LOC_42/B INPUT_1 0.32fF
C23973 AND2X1_LOC_37/a_8_24# D_INPUT_0 0.01fF
C23974 AND2X1_LOC_47/Y OR2X1_LOC_240/A 0.01fF
C23975 OR2X1_LOC_786/A OR2X1_LOC_771/B 0.06fF
C23976 OR2X1_LOC_18/Y OR2X1_LOC_86/A 0.03fF
C23977 OR2X1_LOC_597/Y AND2X1_LOC_655/A 0.06fF
C23978 OR2X1_LOC_51/Y OR2X1_LOC_437/A 0.17fF
C23979 OR2X1_LOC_120/a_36_216# OR2X1_LOC_121/A 0.00fF
C23980 OR2X1_LOC_790/A AND2X1_LOC_36/Y 0.03fF
C23981 OR2X1_LOC_166/a_8_216# OR2X1_LOC_13/B 0.01fF
C23982 OR2X1_LOC_70/Y OR2X1_LOC_71/Y 0.02fF
C23983 OR2X1_LOC_160/A OR2X1_LOC_705/B 0.03fF
C23984 OR2X1_LOC_6/A OR2X1_LOC_29/a_36_216# 0.02fF
C23985 AND2X1_LOC_57/a_8_24# OR2X1_LOC_68/B 0.01fF
C23986 OR2X1_LOC_516/Y AND2X1_LOC_778/Y 3.05fF
C23987 AND2X1_LOC_773/Y AND2X1_LOC_773/a_36_24# 0.00fF
C23988 OR2X1_LOC_76/a_8_216# OR2X1_LOC_553/A 0.05fF
C23989 AND2X1_LOC_682/a_8_24# AND2X1_LOC_31/Y 0.01fF
C23990 OR2X1_LOC_469/Y OR2X1_LOC_546/A 0.00fF
C23991 OR2X1_LOC_317/a_8_216# OR2X1_LOC_317/B 0.07fF
C23992 OR2X1_LOC_244/Y AND2X1_LOC_246/a_36_24# 0.00fF
C23993 OR2X1_LOC_31/Y OR2X1_LOC_52/a_36_216# 0.00fF
C23994 OR2X1_LOC_78/A OR2X1_LOC_712/B 0.05fF
C23995 OR2X1_LOC_529/Y OR2X1_LOC_47/Y 0.06fF
C23996 OR2X1_LOC_232/a_36_216# D_INPUT_1 0.00fF
C23997 OR2X1_LOC_506/A AND2X1_LOC_31/Y 0.04fF
C23998 OR2X1_LOC_26/Y AND2X1_LOC_795/Y 0.15fF
C23999 OR2X1_LOC_715/B OR2X1_LOC_390/B 0.10fF
C24000 VDD OR2X1_LOC_395/Y 0.08fF
C24001 AND2X1_LOC_31/a_8_24# AND2X1_LOC_47/Y 0.19fF
C24002 OR2X1_LOC_461/A OR2X1_LOC_598/A 0.10fF
C24003 AND2X1_LOC_48/A OR2X1_LOC_655/B 0.06fF
C24004 OR2X1_LOC_59/Y AND2X1_LOC_789/Y 0.02fF
C24005 AND2X1_LOC_159/a_8_24# OR2X1_LOC_493/Y 0.12fF
C24006 OR2X1_LOC_158/A AND2X1_LOC_780/a_36_24# 0.00fF
C24007 AND2X1_LOC_414/a_8_24# OR2X1_LOC_71/A 0.02fF
C24008 OR2X1_LOC_479/Y OR2X1_LOC_786/Y 0.00fF
C24009 OR2X1_LOC_88/Y OR2X1_LOC_39/A 0.03fF
C24010 OR2X1_LOC_178/Y OR2X1_LOC_183/Y 0.18fF
C24011 OR2X1_LOC_864/A OR2X1_LOC_598/A 0.07fF
C24012 OR2X1_LOC_265/Y OR2X1_LOC_72/Y 0.52fF
C24013 OR2X1_LOC_174/A OR2X1_LOC_174/Y 0.20fF
C24014 AND2X1_LOC_773/Y AND2X1_LOC_810/A 0.30fF
C24015 OR2X1_LOC_344/A OR2X1_LOC_577/Y 0.05fF
C24016 OR2X1_LOC_89/A AND2X1_LOC_795/Y 0.02fF
C24017 OR2X1_LOC_479/Y OR2X1_LOC_364/a_36_216# 0.02fF
C24018 OR2X1_LOC_31/Y OR2X1_LOC_46/A 0.77fF
C24019 OR2X1_LOC_416/Y OR2X1_LOC_75/a_36_216# 0.00fF
C24020 OR2X1_LOC_323/A AND2X1_LOC_392/A 0.03fF
C24021 OR2X1_LOC_235/B OR2X1_LOC_523/a_8_216# 0.01fF
C24022 OR2X1_LOC_97/A OR2X1_LOC_654/a_8_216# 0.01fF
C24023 AND2X1_LOC_610/a_36_24# AND2X1_LOC_647/Y 0.00fF
C24024 OR2X1_LOC_240/A OR2X1_LOC_598/A 0.01fF
C24025 OR2X1_LOC_633/B OR2X1_LOC_598/A 0.02fF
C24026 OR2X1_LOC_22/A OR2X1_LOC_409/a_8_216# 0.01fF
C24027 AND2X1_LOC_40/a_36_24# AND2X1_LOC_44/Y 0.00fF
C24028 OR2X1_LOC_70/Y OR2X1_LOC_173/a_8_216# 0.06fF
C24029 AND2X1_LOC_163/a_8_24# OR2X1_LOC_161/B 0.02fF
C24030 VDD OR2X1_LOC_722/B 0.06fF
C24031 OR2X1_LOC_62/A AND2X1_LOC_672/B 0.04fF
C24032 AND2X1_LOC_547/Y AND2X1_LOC_564/A 0.12fF
C24033 AND2X1_LOC_655/a_36_24# OR2X1_LOC_46/A 0.00fF
C24034 OR2X1_LOC_619/Y OR2X1_LOC_13/B 0.15fF
C24035 OR2X1_LOC_691/Y OR2X1_LOC_598/Y 0.11fF
C24036 AND2X1_LOC_356/a_8_24# OR2X1_LOC_13/B 0.03fF
C24037 AND2X1_LOC_863/Y AND2X1_LOC_866/A 0.03fF
C24038 AND2X1_LOC_776/a_8_24# AND2X1_LOC_721/Y 0.01fF
C24039 OR2X1_LOC_177/Y AND2X1_LOC_476/Y 0.04fF
C24040 AND2X1_LOC_191/B AND2X1_LOC_242/B 0.29fF
C24041 OR2X1_LOC_680/A OR2X1_LOC_437/A 0.12fF
C24042 AND2X1_LOC_574/a_8_24# AND2X1_LOC_574/Y 0.01fF
C24043 AND2X1_LOC_366/A OR2X1_LOC_89/Y 0.80fF
C24044 OR2X1_LOC_833/Y OR2X1_LOC_629/B 0.81fF
C24045 AND2X1_LOC_810/A AND2X1_LOC_568/B 0.03fF
C24046 OR2X1_LOC_184/Y OR2X1_LOC_71/Y 0.09fF
C24047 OR2X1_LOC_139/A OR2X1_LOC_78/A 0.01fF
C24048 OR2X1_LOC_160/B AND2X1_LOC_603/a_36_24# 0.01fF
C24049 OR2X1_LOC_140/A OR2X1_LOC_549/A 0.14fF
C24050 OR2X1_LOC_585/A OR2X1_LOC_399/a_8_216# 0.05fF
C24051 OR2X1_LOC_523/B AND2X1_LOC_18/Y 0.09fF
C24052 AND2X1_LOC_436/Y AND2X1_LOC_810/B 0.03fF
C24053 OR2X1_LOC_59/Y OR2X1_LOC_585/a_8_216# 0.40fF
C24054 OR2X1_LOC_45/B OR2X1_LOC_329/B 0.26fF
C24055 OR2X1_LOC_604/A AND2X1_LOC_476/Y 0.10fF
C24056 AND2X1_LOC_194/a_8_24# OR2X1_LOC_56/Y 0.23fF
C24057 OR2X1_LOC_56/A OR2X1_LOC_373/Y 0.15fF
C24058 AND2X1_LOC_727/a_36_24# AND2X1_LOC_658/A 0.01fF
C24059 OR2X1_LOC_545/B OR2X1_LOC_545/a_8_216# 0.05fF
C24060 OR2X1_LOC_235/B OR2X1_LOC_576/A 1.14fF
C24061 OR2X1_LOC_604/A OR2X1_LOC_382/a_36_216# -0.00fF
C24062 OR2X1_LOC_518/Y AND2X1_LOC_520/Y 0.79fF
C24063 OR2X1_LOC_160/B AND2X1_LOC_265/a_8_24# 0.04fF
C24064 AND2X1_LOC_531/a_8_24# OR2X1_LOC_563/A 0.04fF
C24065 OR2X1_LOC_516/Y AND2X1_LOC_624/A 0.07fF
C24066 OR2X1_LOC_400/B OR2X1_LOC_771/B 0.01fF
C24067 AND2X1_LOC_40/Y OR2X1_LOC_175/Y 0.02fF
C24068 OR2X1_LOC_84/A OR2X1_LOC_84/a_8_216# 0.18fF
C24069 OR2X1_LOC_820/B AND2X1_LOC_789/Y 0.02fF
C24070 AND2X1_LOC_212/B AND2X1_LOC_212/a_8_24# 0.05fF
C24071 OR2X1_LOC_155/A OR2X1_LOC_712/B 0.01fF
C24072 OR2X1_LOC_492/Y OR2X1_LOC_59/Y 0.24fF
C24073 AND2X1_LOC_367/A OR2X1_LOC_12/Y 0.22fF
C24074 AND2X1_LOC_48/A OR2X1_LOC_750/Y 0.04fF
C24075 OR2X1_LOC_643/Y OR2X1_LOC_68/B 0.06fF
C24076 OR2X1_LOC_738/A OR2X1_LOC_731/A 0.40fF
C24077 OR2X1_LOC_160/B VDD 1.42fF
C24078 OR2X1_LOC_113/B OR2X1_LOC_632/Y 0.00fF
C24079 OR2X1_LOC_607/a_36_216# AND2X1_LOC_647/Y 0.00fF
C24080 OR2X1_LOC_92/Y OR2X1_LOC_428/A 0.32fF
C24081 AND2X1_LOC_40/Y OR2X1_LOC_691/Y 0.02fF
C24082 OR2X1_LOC_329/a_36_216# OR2X1_LOC_329/B 0.00fF
C24083 AND2X1_LOC_509/Y OR2X1_LOC_482/Y 0.03fF
C24084 OR2X1_LOC_830/a_36_216# OR2X1_LOC_190/A 0.00fF
C24085 OR2X1_LOC_290/Y OR2X1_LOC_16/A 0.15fF
C24086 OR2X1_LOC_108/a_8_216# OR2X1_LOC_59/Y 0.01fF
C24087 OR2X1_LOC_856/B AND2X1_LOC_44/Y 0.07fF
C24088 OR2X1_LOC_64/Y AND2X1_LOC_592/a_8_24# 0.03fF
C24089 OR2X1_LOC_430/Y AND2X1_LOC_451/a_8_24# 0.23fF
C24090 D_INPUT_7 D_INPUT_6 1.00fF
C24091 OR2X1_LOC_92/Y OR2X1_LOC_595/A 0.10fF
C24092 OR2X1_LOC_175/Y OR2X1_LOC_537/A 0.28fF
C24093 OR2X1_LOC_810/A OR2X1_LOC_130/a_8_216# 0.14fF
C24094 OR2X1_LOC_246/A OR2X1_LOC_71/A 0.47fF
C24095 AND2X1_LOC_711/Y AND2X1_LOC_789/Y 0.01fF
C24096 AND2X1_LOC_729/Y AND2X1_LOC_564/A 0.03fF
C24097 OR2X1_LOC_597/Y OR2X1_LOC_599/Y 0.04fF
C24098 OR2X1_LOC_51/Y OR2X1_LOC_411/Y 0.20fF
C24099 OR2X1_LOC_47/Y OR2X1_LOC_598/A 0.09fF
C24100 AND2X1_LOC_98/a_8_24# OR2X1_LOC_91/A 0.03fF
C24101 AND2X1_LOC_555/Y AND2X1_LOC_348/Y 0.01fF
C24102 OR2X1_LOC_89/A AND2X1_LOC_439/a_8_24# 0.02fF
C24103 OR2X1_LOC_805/A OR2X1_LOC_362/a_36_216# 0.02fF
C24104 OR2X1_LOC_426/B OR2X1_LOC_59/Y 0.30fF
C24105 OR2X1_LOC_51/Y AND2X1_LOC_851/a_8_24# 0.01fF
C24106 OR2X1_LOC_97/A AND2X1_LOC_43/B 0.03fF
C24107 OR2X1_LOC_516/A AND2X1_LOC_787/A 0.04fF
C24108 OR2X1_LOC_427/A OR2X1_LOC_524/a_8_216# 0.01fF
C24109 AND2X1_LOC_96/a_8_24# OR2X1_LOC_66/A 0.01fF
C24110 OR2X1_LOC_185/A OR2X1_LOC_161/B 0.73fF
C24111 OR2X1_LOC_696/A OR2X1_LOC_238/Y 0.03fF
C24112 AND2X1_LOC_795/Y AND2X1_LOC_804/a_8_24# 0.11fF
C24113 OR2X1_LOC_479/Y OR2X1_LOC_301/a_36_216# 0.01fF
C24114 OR2X1_LOC_158/A AND2X1_LOC_364/A 0.01fF
C24115 AND2X1_LOC_828/a_36_24# OR2X1_LOC_48/B 0.01fF
C24116 AND2X1_LOC_12/Y AND2X1_LOC_603/a_8_24# 0.01fF
C24117 AND2X1_LOC_31/Y OR2X1_LOC_227/Y 0.09fF
C24118 OR2X1_LOC_833/B OR2X1_LOC_549/A 0.02fF
C24119 OR2X1_LOC_98/B OR2X1_LOC_99/A 0.88fF
C24120 OR2X1_LOC_778/Y OR2X1_LOC_703/a_8_216# 0.33fF
C24121 OR2X1_LOC_294/Y OR2X1_LOC_347/B 0.01fF
C24122 OR2X1_LOC_65/B OR2X1_LOC_595/A 0.75fF
C24123 OR2X1_LOC_18/Y AND2X1_LOC_828/a_36_24# 0.00fF
C24124 OR2X1_LOC_455/a_8_216# AND2X1_LOC_7/B 0.01fF
C24125 AND2X1_LOC_31/Y D_INPUT_1 0.02fF
C24126 OR2X1_LOC_786/Y OR2X1_LOC_68/B 0.05fF
C24127 AND2X1_LOC_776/Y OR2X1_LOC_371/Y 0.27fF
C24128 OR2X1_LOC_101/a_8_216# AND2X1_LOC_18/Y 0.02fF
C24129 AND2X1_LOC_719/Y OR2X1_LOC_18/Y 0.09fF
C24130 OR2X1_LOC_95/Y OR2X1_LOC_164/a_36_216# 0.02fF
C24131 OR2X1_LOC_271/Y OR2X1_LOC_428/A 0.03fF
C24132 OR2X1_LOC_814/A OR2X1_LOC_723/B 0.07fF
C24133 AND2X1_LOC_91/B OR2X1_LOC_557/A 0.10fF
C24134 OR2X1_LOC_231/A AND2X1_LOC_18/Y 0.03fF
C24135 OR2X1_LOC_254/B OR2X1_LOC_549/A 0.00fF
C24136 AND2X1_LOC_722/A OR2X1_LOC_744/A 0.03fF
C24137 AND2X1_LOC_544/a_36_24# AND2X1_LOC_658/A 0.01fF
C24138 AND2X1_LOC_553/A OR2X1_LOC_178/Y 0.01fF
C24139 OR2X1_LOC_49/A OR2X1_LOC_49/a_8_216# 0.06fF
C24140 OR2X1_LOC_118/Y OR2X1_LOC_131/a_36_216# 0.00fF
C24141 AND2X1_LOC_865/A AND2X1_LOC_865/a_8_24# 0.04fF
C24142 OR2X1_LOC_850/B OR2X1_LOC_78/A 0.01fF
C24143 OR2X1_LOC_161/A OR2X1_LOC_362/A 0.02fF
C24144 OR2X1_LOC_696/A AND2X1_LOC_855/a_8_24# 0.03fF
C24145 OR2X1_LOC_508/a_36_216# AND2X1_LOC_81/B 0.00fF
C24146 OR2X1_LOC_305/Y OR2X1_LOC_16/A 0.03fF
C24147 OR2X1_LOC_528/a_36_216# AND2X1_LOC_807/Y 0.16fF
C24148 AND2X1_LOC_86/Y VDD 0.05fF
C24149 AND2X1_LOC_706/Y OR2X1_LOC_36/Y 0.02fF
C24150 AND2X1_LOC_203/a_8_24# AND2X1_LOC_203/Y 0.00fF
C24151 OR2X1_LOC_585/Y OR2X1_LOC_586/Y 0.02fF
C24152 AND2X1_LOC_195/a_8_24# OR2X1_LOC_43/A 0.01fF
C24153 INPUT_3 VDD 0.49fF
C24154 OR2X1_LOC_850/a_8_216# OR2X1_LOC_850/B 0.05fF
C24155 OR2X1_LOC_364/A OR2X1_LOC_151/A 0.03fF
C24156 OR2X1_LOC_528/Y OR2X1_LOC_406/a_8_216# 0.01fF
C24157 OR2X1_LOC_185/Y OR2X1_LOC_151/A 0.25fF
C24158 OR2X1_LOC_858/A OR2X1_LOC_737/A 0.03fF
C24159 VDD AND2X1_LOC_452/Y 0.89fF
C24160 AND2X1_LOC_18/Y OR2X1_LOC_340/Y 0.01fF
C24161 AND2X1_LOC_508/B AND2X1_LOC_858/a_8_24# 0.01fF
C24162 AND2X1_LOC_738/B AND2X1_LOC_546/a_8_24# 0.04fF
C24163 AND2X1_LOC_21/Y INPUT_7 0.01fF
C24164 AND2X1_LOC_542/a_8_24# OR2X1_LOC_26/Y 0.01fF
C24165 OR2X1_LOC_517/A AND2X1_LOC_141/A 0.00fF
C24166 OR2X1_LOC_427/A AND2X1_LOC_663/A 0.14fF
C24167 OR2X1_LOC_91/Y OR2X1_LOC_108/Y 0.07fF
C24168 OR2X1_LOC_130/A AND2X1_LOC_18/Y 0.62fF
C24169 OR2X1_LOC_858/A AND2X1_LOC_95/Y 0.01fF
C24170 VDD OR2X1_LOC_799/a_8_216# 0.00fF
C24171 AND2X1_LOC_56/B OR2X1_LOC_730/A 0.02fF
C24172 AND2X1_LOC_486/Y AND2X1_LOC_456/B 0.03fF
C24173 OR2X1_LOC_91/A AND2X1_LOC_520/Y 0.10fF
C24174 AND2X1_LOC_675/Y OR2X1_LOC_531/a_8_216# 0.01fF
C24175 OR2X1_LOC_364/Y OR2X1_LOC_365/B 0.06fF
C24176 AND2X1_LOC_510/A AND2X1_LOC_621/Y 0.06fF
C24177 VDD OR2X1_LOC_553/A 0.77fF
C24178 OR2X1_LOC_40/Y AND2X1_LOC_354/B 0.18fF
C24179 OR2X1_LOC_9/Y OR2X1_LOC_26/Y 0.05fF
C24180 OR2X1_LOC_490/Y OR2X1_LOC_12/Y 0.07fF
C24181 AND2X1_LOC_658/A AND2X1_LOC_858/a_36_24# 0.01fF
C24182 OR2X1_LOC_74/A OR2X1_LOC_12/Y 0.07fF
C24183 AND2X1_LOC_658/A AND2X1_LOC_622/a_36_24# 0.01fF
C24184 VDD OR2X1_LOC_266/a_8_216# 0.00fF
C24185 OR2X1_LOC_405/A OR2X1_LOC_538/A 0.03fF
C24186 AND2X1_LOC_753/B D_INPUT_5 0.03fF
C24187 AND2X1_LOC_577/a_8_24# AND2X1_LOC_577/Y 0.00fF
C24188 OR2X1_LOC_640/a_8_216# AND2X1_LOC_92/Y 0.12fF
C24189 AND2X1_LOC_539/a_36_24# OR2X1_LOC_43/A 0.01fF
C24190 OR2X1_LOC_121/B OR2X1_LOC_352/a_8_216# 0.03fF
C24191 OR2X1_LOC_335/A OR2X1_LOC_814/A 0.00fF
C24192 AND2X1_LOC_713/a_36_24# OR2X1_LOC_89/A 0.00fF
C24193 AND2X1_LOC_318/Y OR2X1_LOC_268/Y 0.00fF
C24194 OR2X1_LOC_456/A OR2X1_LOC_577/Y 0.22fF
C24195 OR2X1_LOC_426/A OR2X1_LOC_426/Y 0.01fF
C24196 AND2X1_LOC_199/a_36_24# OR2X1_LOC_43/A -0.00fF
C24197 AND2X1_LOC_47/Y OR2X1_LOC_501/A 0.01fF
C24198 OR2X1_LOC_485/Y OR2X1_LOC_52/B 0.03fF
C24199 AND2X1_LOC_570/Y AND2X1_LOC_575/Y 0.01fF
C24200 OR2X1_LOC_715/B AND2X1_LOC_516/a_36_24# 0.01fF
C24201 OR2X1_LOC_158/A OR2X1_LOC_3/Y 1.93fF
C24202 OR2X1_LOC_541/A AND2X1_LOC_43/B 0.03fF
C24203 OR2X1_LOC_674/a_36_216# OR2X1_LOC_39/A 0.00fF
C24204 VDD OR2X1_LOC_219/B 0.13fF
C24205 OR2X1_LOC_532/B OR2X1_LOC_415/Y 0.51fF
C24206 OR2X1_LOC_51/Y OR2X1_LOC_753/A 0.07fF
C24207 OR2X1_LOC_84/Y OR2X1_LOC_771/B 0.03fF
C24208 AND2X1_LOC_47/Y AND2X1_LOC_760/a_8_24# 0.07fF
C24209 OR2X1_LOC_427/A OR2X1_LOC_2/Y 0.10fF
C24210 OR2X1_LOC_291/Y OR2X1_LOC_16/A 0.32fF
C24211 OR2X1_LOC_9/Y OR2X1_LOC_824/a_36_216# 0.00fF
C24212 OR2X1_LOC_474/Y OR2X1_LOC_161/A 0.05fF
C24213 OR2X1_LOC_158/A AND2X1_LOC_473/a_36_24# 0.01fF
C24214 OR2X1_LOC_599/A OR2X1_LOC_744/A 0.82fF
C24215 INPUT_0 OR2X1_LOC_6/A 1.54fF
C24216 OR2X1_LOC_756/B OR2X1_LOC_664/Y 0.00fF
C24217 OR2X1_LOC_40/Y AND2X1_LOC_390/B 0.01fF
C24218 OR2X1_LOC_667/Y AND2X1_LOC_720/a_8_24# 0.23fF
C24219 OR2X1_LOC_539/A OR2X1_LOC_161/A 0.01fF
C24220 OR2X1_LOC_311/Y OR2X1_LOC_16/A 0.03fF
C24221 OR2X1_LOC_160/A OR2X1_LOC_502/A 0.45fF
C24222 OR2X1_LOC_185/A OR2X1_LOC_61/Y 0.03fF
C24223 AND2X1_LOC_33/a_8_24# OR2X1_LOC_24/Y -0.01fF
C24224 AND2X1_LOC_123/a_8_24# OR2X1_LOC_56/A 0.02fF
C24225 OR2X1_LOC_6/B OR2X1_LOC_8/a_8_216# 0.01fF
C24226 OR2X1_LOC_185/Y AND2X1_LOC_67/a_8_24# 0.03fF
C24227 AND2X1_LOC_47/Y OR2X1_LOC_121/A 0.03fF
C24228 AND2X1_LOC_421/a_8_24# OR2X1_LOC_375/A 0.01fF
C24229 AND2X1_LOC_70/Y OR2X1_LOC_787/Y 0.02fF
C24230 AND2X1_LOC_347/B AND2X1_LOC_663/B 0.00fF
C24231 AND2X1_LOC_51/Y OR2X1_LOC_362/A 0.03fF
C24232 OR2X1_LOC_176/Y OR2X1_LOC_167/Y 0.03fF
C24233 OR2X1_LOC_601/a_8_216# OR2X1_LOC_16/A 0.03fF
C24234 OR2X1_LOC_525/Y AND2X1_LOC_621/Y 0.06fF
C24235 AND2X1_LOC_397/a_8_24# AND2X1_LOC_3/Y 0.03fF
C24236 VDD OR2X1_LOC_321/Y 0.16fF
C24237 AND2X1_LOC_535/a_8_24# AND2X1_LOC_390/B 0.02fF
C24238 AND2X1_LOC_520/a_36_24# OR2X1_LOC_111/Y 0.00fF
C24239 OR2X1_LOC_850/A OR2X1_LOC_862/B 0.72fF
C24240 AND2X1_LOC_65/a_36_24# OR2X1_LOC_87/A 0.01fF
C24241 OR2X1_LOC_256/Y OR2X1_LOC_248/a_8_216# 0.02fF
C24242 OR2X1_LOC_22/Y OR2X1_LOC_13/a_8_216# 0.03fF
C24243 OR2X1_LOC_479/Y OR2X1_LOC_467/A 0.00fF
C24244 AND2X1_LOC_72/B OR2X1_LOC_500/a_36_216# 0.00fF
C24245 OR2X1_LOC_427/A AND2X1_LOC_449/Y 0.02fF
C24246 AND2X1_LOC_533/a_36_24# OR2X1_LOC_620/Y 0.00fF
C24247 OR2X1_LOC_40/Y OR2X1_LOC_431/Y 0.46fF
C24248 AND2X1_LOC_76/Y OR2X1_LOC_39/A 0.03fF
C24249 AND2X1_LOC_850/a_36_24# OR2X1_LOC_18/Y 0.00fF
C24250 OR2X1_LOC_70/Y OR2X1_LOC_426/B 5.79fF
C24251 OR2X1_LOC_48/B AND2X1_LOC_655/A 0.07fF
C24252 AND2X1_LOC_12/Y OR2X1_LOC_405/A 0.08fF
C24253 OR2X1_LOC_364/A OR2X1_LOC_788/a_8_216# 0.03fF
C24254 OR2X1_LOC_259/a_8_216# OR2X1_LOC_375/A 0.16fF
C24255 OR2X1_LOC_538/a_36_216# OR2X1_LOC_269/B 0.02fF
C24256 OR2X1_LOC_290/a_36_216# OR2X1_LOC_690/A 0.00fF
C24257 OR2X1_LOC_160/A AND2X1_LOC_230/a_8_24# 0.01fF
C24258 OR2X1_LOC_129/a_8_216# OR2X1_LOC_46/A 0.01fF
C24259 OR2X1_LOC_91/Y AND2X1_LOC_168/Y 0.04fF
C24260 OR2X1_LOC_18/Y AND2X1_LOC_655/A 0.01fF
C24261 AND2X1_LOC_456/B OR2X1_LOC_666/Y 0.01fF
C24262 AND2X1_LOC_729/Y AND2X1_LOC_593/Y 0.07fF
C24263 OR2X1_LOC_256/Y AND2X1_LOC_294/a_8_24# 0.01fF
C24264 OR2X1_LOC_358/A OR2X1_LOC_333/A 0.86fF
C24265 OR2X1_LOC_405/A OR2X1_LOC_802/A 0.02fF
C24266 OR2X1_LOC_263/a_8_216# AND2X1_LOC_243/Y 0.04fF
C24267 OR2X1_LOC_216/A AND2X1_LOC_3/Y 0.01fF
C24268 AND2X1_LOC_36/Y AND2X1_LOC_751/a_8_24# 0.01fF
C24269 OR2X1_LOC_502/A AND2X1_LOC_611/a_36_24# 0.00fF
C24270 AND2X1_LOC_514/Y OR2X1_LOC_426/B 0.07fF
C24271 OR2X1_LOC_62/B AND2X1_LOC_18/Y 0.09fF
C24272 AND2X1_LOC_486/Y AND2X1_LOC_717/B 0.18fF
C24273 AND2X1_LOC_798/A AND2X1_LOC_802/Y 0.46fF
C24274 AND2X1_LOC_387/B D_INPUT_4 0.01fF
C24275 OR2X1_LOC_186/Y OR2X1_LOC_112/B 0.06fF
C24276 OR2X1_LOC_541/B OR2X1_LOC_269/B 0.09fF
C24277 AND2X1_LOC_42/B AND2X1_LOC_619/B 0.01fF
C24278 AND2X1_LOC_654/Y OR2X1_LOC_299/a_36_216# 0.01fF
C24279 OR2X1_LOC_91/A AND2X1_LOC_863/A 0.00fF
C24280 AND2X1_LOC_572/Y OR2X1_LOC_26/Y 0.02fF
C24281 VDD OR2X1_LOC_244/A 0.99fF
C24282 OR2X1_LOC_246/A OR2X1_LOC_59/Y 0.03fF
C24283 OR2X1_LOC_851/A OR2X1_LOC_479/Y 0.03fF
C24284 OR2X1_LOC_309/Y AND2X1_LOC_866/A 0.00fF
C24285 OR2X1_LOC_474/Y AND2X1_LOC_51/Y 0.03fF
C24286 OR2X1_LOC_532/B AND2X1_LOC_616/a_8_24# 0.01fF
C24287 AND2X1_LOC_580/A OR2X1_LOC_44/Y 0.03fF
C24288 OR2X1_LOC_39/A OR2X1_LOC_52/B 0.11fF
C24289 OR2X1_LOC_789/B OR2X1_LOC_789/a_8_216# 0.47fF
C24290 AND2X1_LOC_729/Y AND2X1_LOC_602/a_8_24# 0.02fF
C24291 OR2X1_LOC_669/Y AND2X1_LOC_848/Y 0.32fF
C24292 OR2X1_LOC_499/a_8_216# AND2X1_LOC_3/Y 0.01fF
C24293 AND2X1_LOC_572/Y OR2X1_LOC_89/A 0.04fF
C24294 OR2X1_LOC_656/B OR2X1_LOC_216/a_8_216# 0.04fF
C24295 OR2X1_LOC_316/Y OR2X1_LOC_7/A 0.00fF
C24296 OR2X1_LOC_474/Y OR2X1_LOC_849/a_8_216# 0.06fF
C24297 OR2X1_LOC_690/A OR2X1_LOC_6/A 0.02fF
C24298 OR2X1_LOC_26/Y AND2X1_LOC_834/a_36_24# 0.01fF
C24299 OR2X1_LOC_532/B OR2X1_LOC_632/Y 0.11fF
C24300 OR2X1_LOC_70/A OR2X1_LOC_585/a_8_216# 0.01fF
C24301 AND2X1_LOC_59/Y OR2X1_LOC_204/a_8_216# 0.14fF
C24302 AND2X1_LOC_18/Y AND2X1_LOC_88/Y 0.83fF
C24303 AND2X1_LOC_647/Y OR2X1_LOC_12/Y 0.00fF
C24304 OR2X1_LOC_26/Y AND2X1_LOC_852/Y 0.06fF
C24305 OR2X1_LOC_665/Y OR2X1_LOC_36/Y 0.03fF
C24306 AND2X1_LOC_813/a_8_24# OR2X1_LOC_66/A 0.01fF
C24307 AND2X1_LOC_111/a_36_24# OR2X1_LOC_161/A 0.01fF
C24308 OR2X1_LOC_409/B OR2X1_LOC_59/Y 0.00fF
C24309 OR2X1_LOC_157/a_36_216# OR2X1_LOC_429/Y 0.01fF
C24310 AND2X1_LOC_168/Y OR2X1_LOC_417/Y 0.00fF
C24311 AND2X1_LOC_42/B OR2X1_LOC_87/a_36_216# 0.00fF
C24312 OR2X1_LOC_744/A AND2X1_LOC_866/A 0.07fF
C24313 OR2X1_LOC_83/Y OR2X1_LOC_26/Y 0.07fF
C24314 OR2X1_LOC_8/Y OR2X1_LOC_826/Y 0.01fF
C24315 AND2X1_LOC_663/B OR2X1_LOC_118/Y 0.03fF
C24316 OR2X1_LOC_400/A OR2X1_LOC_624/B 0.01fF
C24317 OR2X1_LOC_485/A OR2X1_LOC_36/Y 0.24fF
C24318 AND2X1_LOC_350/Y OR2X1_LOC_18/Y 0.03fF
C24319 INPUT_0 D_INPUT_2 0.02fF
C24320 AND2X1_LOC_679/a_8_24# OR2X1_LOC_596/A 0.01fF
C24321 OR2X1_LOC_743/A OR2X1_LOC_433/a_8_216# 0.01fF
C24322 AND2X1_LOC_211/B OR2X1_LOC_52/B 0.03fF
C24323 OR2X1_LOC_679/A OR2X1_LOC_144/Y 0.01fF
C24324 AND2X1_LOC_722/A OR2X1_LOC_31/Y 0.01fF
C24325 AND2X1_LOC_51/A AND2X1_LOC_21/Y 0.07fF
C24326 AND2X1_LOC_7/B AND2X1_LOC_419/a_8_24# 0.01fF
C24327 AND2X1_LOC_41/A OR2X1_LOC_276/B 0.07fF
C24328 OR2X1_LOC_154/A OR2X1_LOC_473/Y 0.03fF
C24329 AND2X1_LOC_36/Y OR2X1_LOC_714/a_8_216# 0.01fF
C24330 VDD AND2X1_LOC_793/Y 0.24fF
C24331 OR2X1_LOC_812/B OR2X1_LOC_814/A 0.01fF
C24332 OR2X1_LOC_97/A OR2X1_LOC_367/B 0.03fF
C24333 OR2X1_LOC_844/a_36_216# OR2X1_LOC_643/A 0.00fF
C24334 AND2X1_LOC_351/Y OR2X1_LOC_265/Y 0.03fF
C24335 OR2X1_LOC_160/A AND2X1_LOC_48/A 0.03fF
C24336 OR2X1_LOC_64/Y OR2X1_LOC_6/A 0.02fF
C24337 OR2X1_LOC_643/Y OR2X1_LOC_219/a_8_216# 0.39fF
C24338 OR2X1_LOC_19/B OR2X1_LOC_67/a_8_216# 0.10fF
C24339 OR2X1_LOC_485/A AND2X1_LOC_493/a_36_24# 0.00fF
C24340 OR2X1_LOC_151/A OR2X1_LOC_568/A 0.07fF
C24341 AND2X1_LOC_36/Y OR2X1_LOC_731/A 0.47fF
C24342 AND2X1_LOC_390/B OR2X1_LOC_7/A 0.14fF
C24343 OR2X1_LOC_689/a_36_216# OR2X1_LOC_31/Y 0.03fF
C24344 OR2X1_LOC_500/A OR2X1_LOC_62/B 0.03fF
C24345 AND2X1_LOC_319/A AND2X1_LOC_727/A 0.00fF
C24346 OR2X1_LOC_282/a_36_216# OR2X1_LOC_89/A 0.02fF
C24347 OR2X1_LOC_151/A OR2X1_LOC_151/a_8_216# 0.01fF
C24348 OR2X1_LOC_272/Y OR2X1_LOC_74/A 0.05fF
C24349 OR2X1_LOC_70/Y OR2X1_LOC_743/A 0.35fF
C24350 AND2X1_LOC_70/Y AND2X1_LOC_52/Y 0.03fF
C24351 OR2X1_LOC_676/Y OR2X1_LOC_228/Y 0.43fF
C24352 OR2X1_LOC_484/Y AND2X1_LOC_486/a_8_24# 0.02fF
C24353 OR2X1_LOC_494/Y AND2X1_LOC_657/A 0.01fF
C24354 OR2X1_LOC_676/Y OR2X1_LOC_513/Y 0.01fF
C24355 OR2X1_LOC_377/A OR2X1_LOC_62/A 0.13fF
C24356 OR2X1_LOC_244/A OR2X1_LOC_267/a_36_216# 0.01fF
C24357 AND2X1_LOC_319/A OR2X1_LOC_95/Y 0.02fF
C24358 AND2X1_LOC_356/B OR2X1_LOC_22/Y 0.03fF
C24359 OR2X1_LOC_280/Y OR2X1_LOC_22/Y 0.07fF
C24360 OR2X1_LOC_599/A OR2X1_LOC_31/Y 0.06fF
C24361 AND2X1_LOC_538/a_8_24# OR2X1_LOC_743/A 0.00fF
C24362 OR2X1_LOC_678/Y OR2X1_LOC_512/Y 0.01fF
C24363 OR2X1_LOC_834/A OR2X1_LOC_513/Y 0.09fF
C24364 AND2X1_LOC_851/A OR2X1_LOC_419/Y 0.03fF
C24365 AND2X1_LOC_41/A OR2X1_LOC_779/B 0.10fF
C24366 AND2X1_LOC_831/a_8_24# AND2X1_LOC_476/A 0.04fF
C24367 OR2X1_LOC_252/Y AND2X1_LOC_620/Y 0.02fF
C24368 OR2X1_LOC_62/A OR2X1_LOC_85/A 3.25fF
C24369 AND2X1_LOC_738/B OR2X1_LOC_533/a_36_216# -0.01fF
C24370 AND2X1_LOC_476/A OR2X1_LOC_44/Y 0.07fF
C24371 OR2X1_LOC_70/Y OR2X1_LOC_246/A 0.02fF
C24372 AND2X1_LOC_680/a_8_24# AND2X1_LOC_51/Y 0.05fF
C24373 OR2X1_LOC_696/A AND2X1_LOC_407/a_8_24# 0.04fF
C24374 OR2X1_LOC_333/B D_INPUT_0 0.03fF
C24375 OR2X1_LOC_440/A OR2X1_LOC_269/B 0.06fF
C24376 AND2X1_LOC_554/B OR2X1_LOC_255/a_8_216# 0.14fF
C24377 OR2X1_LOC_278/a_8_216# D_INPUT_0 0.03fF
C24378 OR2X1_LOC_36/Y OR2X1_LOC_587/a_8_216# 0.43fF
C24379 AND2X1_LOC_578/A AND2X1_LOC_477/A 0.01fF
C24380 AND2X1_LOC_863/Y OR2X1_LOC_7/A 0.07fF
C24381 OR2X1_LOC_348/Y OR2X1_LOC_349/B 0.08fF
C24382 AND2X1_LOC_463/B OR2X1_LOC_11/Y 0.47fF
C24383 OR2X1_LOC_616/Y AND2X1_LOC_793/Y 0.00fF
C24384 OR2X1_LOC_349/a_8_216# OR2X1_LOC_349/B 0.01fF
C24385 OR2X1_LOC_154/A OR2X1_LOC_214/B 0.05fF
C24386 OR2X1_LOC_36/Y OR2X1_LOC_609/Y 0.01fF
C24387 OR2X1_LOC_392/A OR2X1_LOC_561/B 0.02fF
C24388 OR2X1_LOC_222/a_8_216# AND2X1_LOC_3/Y 0.05fF
C24389 OR2X1_LOC_6/B AND2X1_LOC_36/Y 0.05fF
C24390 OR2X1_LOC_154/A OR2X1_LOC_241/B 0.13fF
C24391 OR2X1_LOC_16/A OR2X1_LOC_171/Y 0.13fF
C24392 AND2X1_LOC_31/Y OR2X1_LOC_737/A 0.08fF
C24393 AND2X1_LOC_633/Y OR2X1_LOC_65/Y 0.16fF
C24394 OR2X1_LOC_726/A OR2X1_LOC_727/a_8_216# 0.39fF
C24395 OR2X1_LOC_851/A OR2X1_LOC_68/B 0.12fF
C24396 OR2X1_LOC_864/A D_INPUT_1 0.03fF
C24397 OR2X1_LOC_532/B OR2X1_LOC_285/B 0.09fF
C24398 AND2X1_LOC_11/Y AND2X1_LOC_429/a_36_24# 0.01fF
C24399 AND2X1_LOC_468/B AND2X1_LOC_222/Y 0.01fF
C24400 AND2X1_LOC_140/a_8_24# OR2X1_LOC_95/Y 0.04fF
C24401 OR2X1_LOC_160/A OR2X1_LOC_398/a_8_216# 0.01fF
C24402 AND2X1_LOC_452/Y OR2X1_LOC_163/Y 0.08fF
C24403 OR2X1_LOC_138/a_8_216# OR2X1_LOC_691/Y 0.01fF
C24404 OR2X1_LOC_774/Y D_INPUT_1 1.42fF
C24405 OR2X1_LOC_70/Y OR2X1_LOC_409/B 0.06fF
C24406 OR2X1_LOC_714/Y OR2X1_LOC_724/A 0.14fF
C24407 OR2X1_LOC_196/B AND2X1_LOC_692/a_8_24# 0.22fF
C24408 AND2X1_LOC_95/Y AND2X1_LOC_31/Y 0.11fF
C24409 VDD OR2X1_LOC_731/B -0.00fF
C24410 AND2X1_LOC_721/Y AND2X1_LOC_785/Y 0.01fF
C24411 OR2X1_LOC_12/Y AND2X1_LOC_773/a_36_24# 0.01fF
C24412 AND2X1_LOC_48/A OR2X1_LOC_655/A 0.01fF
C24413 OR2X1_LOC_633/B D_INPUT_1 0.03fF
C24414 OR2X1_LOC_52/B AND2X1_LOC_781/Y 0.09fF
C24415 OR2X1_LOC_170/A OR2X1_LOC_365/B 0.01fF
C24416 OR2X1_LOC_205/Y AND2X1_LOC_3/Y 0.04fF
C24417 AND2X1_LOC_170/B AND2X1_LOC_727/A 0.03fF
C24418 AND2X1_LOC_392/A OR2X1_LOC_134/a_8_216# 0.05fF
C24419 OR2X1_LOC_481/A OR2X1_LOC_47/Y 0.01fF
C24420 OR2X1_LOC_185/A AND2X1_LOC_406/a_8_24# 0.01fF
C24421 OR2X1_LOC_368/a_36_216# AND2X1_LOC_543/Y 0.00fF
C24422 OR2X1_LOC_85/A OR2X1_LOC_88/Y 0.02fF
C24423 OR2X1_LOC_485/A OR2X1_LOC_419/Y 0.09fF
C24424 AND2X1_LOC_173/a_8_24# OR2X1_LOC_112/A 0.20fF
C24425 OR2X1_LOC_643/A OR2X1_LOC_641/B 0.03fF
C24426 OR2X1_LOC_502/A OR2X1_LOC_532/Y 0.22fF
C24427 OR2X1_LOC_403/B OR2X1_LOC_398/Y 0.01fF
C24428 D_INPUT_3 AND2X1_LOC_128/a_8_24# 0.01fF
C24429 OR2X1_LOC_533/Y AND2X1_LOC_788/a_8_24# 0.01fF
C24430 AND2X1_LOC_43/B OR2X1_LOC_193/a_8_216# 0.03fF
C24431 AND2X1_LOC_778/a_36_24# OR2X1_LOC_56/A 0.00fF
C24432 OR2X1_LOC_808/B OR2X1_LOC_308/Y 0.10fF
C24433 AND2X1_LOC_721/Y AND2X1_LOC_489/a_8_24# 0.14fF
C24434 OR2X1_LOC_40/Y AND2X1_LOC_639/B 0.10fF
C24435 OR2X1_LOC_178/Y AND2X1_LOC_465/A 0.02fF
C24436 D_INPUT_3 OR2X1_LOC_225/a_36_216# 0.00fF
C24437 AND2X1_LOC_3/Y OR2X1_LOC_750/Y 0.05fF
C24438 AND2X1_LOC_542/a_8_24# AND2X1_LOC_552/A 0.00fF
C24439 AND2X1_LOC_315/a_8_24# OR2X1_LOC_181/Y 0.23fF
C24440 OR2X1_LOC_600/A OR2X1_LOC_428/A 0.18fF
C24441 AND2X1_LOC_866/A OR2X1_LOC_31/Y 0.03fF
C24442 AND2X1_LOC_477/Y AND2X1_LOC_469/a_8_24# 0.03fF
C24443 OR2X1_LOC_169/B OR2X1_LOC_788/B 0.01fF
C24444 OR2X1_LOC_604/A OR2X1_LOC_603/Y 0.02fF
C24445 AND2X1_LOC_570/Y AND2X1_LOC_242/a_8_24# 0.01fF
C24446 OR2X1_LOC_47/Y OR2X1_LOC_71/Y 0.02fF
C24447 OR2X1_LOC_600/A OR2X1_LOC_595/A 0.07fF
C24448 AND2X1_LOC_184/a_8_24# OR2X1_LOC_294/Y 0.01fF
C24449 AND2X1_LOC_359/B OR2X1_LOC_437/A 0.23fF
C24450 VDD OR2X1_LOC_36/a_8_216# 0.00fF
C24451 AND2X1_LOC_193/Y AND2X1_LOC_194/Y 0.21fF
C24452 OR2X1_LOC_368/a_36_216# OR2X1_LOC_322/Y 0.00fF
C24453 OR2X1_LOC_40/Y OR2X1_LOC_309/Y 0.01fF
C24454 AND2X1_LOC_70/Y OR2X1_LOC_439/B 0.00fF
C24455 AND2X1_LOC_721/A OR2X1_LOC_95/Y 0.03fF
C24456 AND2X1_LOC_157/a_36_24# INPUT_6 -0.00fF
C24457 OR2X1_LOC_840/A AND2X1_LOC_7/B 0.10fF
C24458 AND2X1_LOC_47/Y AND2X1_LOC_72/B 0.04fF
C24459 VDD AND2X1_LOC_357/B 0.01fF
C24460 AND2X1_LOC_339/B AND2X1_LOC_219/Y 0.02fF
C24461 OR2X1_LOC_196/Y OR2X1_LOC_502/A 0.03fF
C24462 OR2X1_LOC_821/Y OR2X1_LOC_235/B 0.00fF
C24463 AND2X1_LOC_91/B OR2X1_LOC_814/Y 0.01fF
C24464 OR2X1_LOC_808/B AND2X1_LOC_604/a_8_24# 0.12fF
C24465 AND2X1_LOC_633/Y OR2X1_LOC_72/Y 0.02fF
C24466 AND2X1_LOC_463/B OR2X1_LOC_409/a_36_216# 0.00fF
C24467 OR2X1_LOC_532/B OR2X1_LOC_358/A 0.00fF
C24468 OR2X1_LOC_47/Y D_INPUT_1 0.07fF
C24469 OR2X1_LOC_648/B OR2X1_LOC_35/Y 0.03fF
C24470 OR2X1_LOC_158/A OR2X1_LOC_329/B 0.88fF
C24471 VDD OR2X1_LOC_494/Y 0.25fF
C24472 OR2X1_LOC_254/a_8_216# OR2X1_LOC_366/Y 0.05fF
C24473 AND2X1_LOC_803/B OR2X1_LOC_679/a_36_216# 0.00fF
C24474 OR2X1_LOC_702/A OR2X1_LOC_332/a_8_216# 0.07fF
C24475 VDD AND2X1_LOC_363/Y 0.19fF
C24476 OR2X1_LOC_333/B OR2X1_LOC_339/A 0.02fF
C24477 OR2X1_LOC_377/A OR2X1_LOC_397/Y 0.09fF
C24478 OR2X1_LOC_40/Y OR2X1_LOC_744/A 0.28fF
C24479 OR2X1_LOC_676/Y OR2X1_LOC_702/a_36_216# 0.01fF
C24480 OR2X1_LOC_70/A OR2X1_LOC_409/B 0.89fF
C24481 AND2X1_LOC_738/B AND2X1_LOC_447/Y 0.10fF
C24482 OR2X1_LOC_175/Y AND2X1_LOC_43/B 0.07fF
C24483 OR2X1_LOC_95/Y OR2X1_LOC_331/Y 0.18fF
C24484 VDD AND2X1_LOC_548/Y 0.01fF
C24485 AND2X1_LOC_558/a_8_24# AND2X1_LOC_561/B 0.01fF
C24486 OR2X1_LOC_619/Y OR2X1_LOC_428/A 0.10fF
C24487 AND2X1_LOC_509/Y AND2X1_LOC_508/B 0.12fF
C24488 OR2X1_LOC_316/Y AND2X1_LOC_476/a_8_24# 0.00fF
C24489 OR2X1_LOC_811/A OR2X1_LOC_294/Y 0.03fF
C24490 AND2X1_LOC_624/B AND2X1_LOC_793/Y 0.02fF
C24491 AND2X1_LOC_51/Y OR2X1_LOC_771/B 0.10fF
C24492 OR2X1_LOC_158/A OR2X1_LOC_74/Y 0.03fF
C24493 OR2X1_LOC_634/A OR2X1_LOC_66/A 0.90fF
C24494 AND2X1_LOC_509/Y AND2X1_LOC_508/a_8_24# 0.01fF
C24495 OR2X1_LOC_121/Y OR2X1_LOC_115/a_8_216# 0.03fF
C24496 OR2X1_LOC_323/A AND2X1_LOC_458/a_8_24# 0.00fF
C24497 OR2X1_LOC_222/A AND2X1_LOC_7/B 0.03fF
C24498 OR2X1_LOC_8/Y AND2X1_LOC_240/a_8_24# 0.17fF
C24499 AND2X1_LOC_510/a_8_24# AND2X1_LOC_658/A 0.05fF
C24500 AND2X1_LOC_43/B OR2X1_LOC_375/Y 0.01fF
C24501 VDD OR2X1_LOC_307/B -0.00fF
C24502 AND2X1_LOC_70/Y AND2X1_LOC_41/A 0.17fF
C24503 OR2X1_LOC_243/A OR2X1_LOC_633/A 0.02fF
C24504 OR2X1_LOC_17/Y OR2X1_LOC_387/A 0.00fF
C24505 OR2X1_LOC_49/A AND2X1_LOC_80/a_8_24# 0.03fF
C24506 AND2X1_LOC_539/a_8_24# OR2X1_LOC_13/B 0.01fF
C24507 OR2X1_LOC_604/A AND2X1_LOC_168/a_8_24# 0.13fF
C24508 OR2X1_LOC_404/Y OR2X1_LOC_523/a_8_216# 0.02fF
C24509 OR2X1_LOC_45/B AND2X1_LOC_580/A 0.03fF
C24510 INPUT_5 VDD 0.49fF
C24511 AND2X1_LOC_784/A OR2X1_LOC_136/Y 0.42fF
C24512 OR2X1_LOC_40/Y AND2X1_LOC_168/a_36_24# 0.00fF
C24513 AND2X1_LOC_2/Y AND2X1_LOC_12/a_8_24# 0.20fF
C24514 AND2X1_LOC_95/a_8_24# OR2X1_LOC_502/A 0.01fF
C24515 OR2X1_LOC_91/Y OR2X1_LOC_373/Y 0.14fF
C24516 AND2X1_LOC_51/Y OR2X1_LOC_776/A 0.03fF
C24517 VDD AND2X1_LOC_839/a_8_24# -0.00fF
C24518 OR2X1_LOC_485/A AND2X1_LOC_590/a_36_24# 0.00fF
C24519 AND2X1_LOC_564/A OR2X1_LOC_52/B 0.03fF
C24520 AND2X1_LOC_445/a_8_24# OR2X1_LOC_44/Y 0.03fF
C24521 OR2X1_LOC_756/B AND2X1_LOC_24/a_8_24# 0.01fF
C24522 AND2X1_LOC_787/A OR2X1_LOC_26/Y 0.03fF
C24523 OR2X1_LOC_325/B OR2X1_LOC_620/Y 0.08fF
C24524 OR2X1_LOC_317/a_36_216# AND2X1_LOC_92/Y 0.02fF
C24525 AND2X1_LOC_244/A AND2X1_LOC_806/A 0.03fF
C24526 OR2X1_LOC_158/A AND2X1_LOC_113/Y 0.00fF
C24527 AND2X1_LOC_727/Y OR2X1_LOC_74/A 0.03fF
C24528 OR2X1_LOC_599/A AND2X1_LOC_213/B 0.00fF
C24529 AND2X1_LOC_772/B OR2X1_LOC_92/Y 0.05fF
C24530 AND2X1_LOC_509/Y AND2X1_LOC_850/A 0.08fF
C24531 AND2X1_LOC_191/B AND2X1_LOC_866/B 0.34fF
C24532 OR2X1_LOC_33/A OR2X1_LOC_338/A 0.01fF
C24533 OR2X1_LOC_97/A OR2X1_LOC_810/A 0.03fF
C24534 AND2X1_LOC_562/a_8_24# OR2X1_LOC_3/Y 0.01fF
C24535 AND2X1_LOC_555/Y OR2X1_LOC_481/Y 0.00fF
C24536 AND2X1_LOC_357/a_8_24# OR2X1_LOC_426/B 0.04fF
C24537 OR2X1_LOC_744/Y OR2X1_LOC_52/B 0.01fF
C24538 OR2X1_LOC_68/Y AND2X1_LOC_36/Y 0.11fF
C24539 AND2X1_LOC_392/A OR2X1_LOC_118/Y 0.10fF
C24540 AND2X1_LOC_535/Y AND2X1_LOC_436/B -0.00fF
C24541 OR2X1_LOC_465/Y OR2X1_LOC_741/Y 0.00fF
C24542 OR2X1_LOC_187/Y AND2X1_LOC_711/Y 0.01fF
C24543 AND2X1_LOC_42/B OR2X1_LOC_563/A 0.07fF
C24544 AND2X1_LOC_215/Y OR2X1_LOC_619/Y 0.07fF
C24545 AND2X1_LOC_508/A AND2X1_LOC_506/a_36_24# 0.00fF
C24546 OR2X1_LOC_155/A OR2X1_LOC_138/A 0.05fF
C24547 AND2X1_LOC_796/a_8_24# OR2X1_LOC_680/A 0.03fF
C24548 OR2X1_LOC_502/A AND2X1_LOC_144/a_36_24# 0.01fF
C24549 AND2X1_LOC_768/a_36_24# OR2X1_LOC_427/A 0.00fF
C24550 OR2X1_LOC_438/Y AND2X1_LOC_734/Y 0.03fF
C24551 OR2X1_LOC_744/A AND2X1_LOC_843/Y 0.11fF
C24552 OR2X1_LOC_223/A OR2X1_LOC_181/a_36_216# 0.00fF
C24553 OR2X1_LOC_9/Y OR2X1_LOC_246/a_8_216# 0.07fF
C24554 AND2X1_LOC_765/a_36_24# AND2X1_LOC_3/Y 0.00fF
C24555 AND2X1_LOC_512/Y OR2X1_LOC_92/Y 0.07fF
C24556 OR2X1_LOC_186/Y OR2X1_LOC_574/A 0.03fF
C24557 OR2X1_LOC_109/Y OR2X1_LOC_56/A 0.03fF
C24558 AND2X1_LOC_47/Y AND2X1_LOC_36/Y 0.26fF
C24559 AND2X1_LOC_621/Y AND2X1_LOC_658/Y 0.12fF
C24560 OR2X1_LOC_64/Y OR2X1_LOC_184/a_8_216# 0.01fF
C24561 OR2X1_LOC_348/Y AND2X1_LOC_282/a_8_24# 0.02fF
C24562 OR2X1_LOC_319/B OR2X1_LOC_840/A 0.10fF
C24563 OR2X1_LOC_40/Y AND2X1_LOC_840/B 0.02fF
C24564 OR2X1_LOC_203/Y OR2X1_LOC_629/B 0.05fF
C24565 OR2X1_LOC_702/A OR2X1_LOC_161/B 0.03fF
C24566 AND2X1_LOC_570/Y AND2X1_LOC_502/a_8_24# 0.07fF
C24567 OR2X1_LOC_58/Y OR2X1_LOC_80/Y 0.00fF
C24568 AND2X1_LOC_729/Y OR2X1_LOC_51/Y 0.02fF
C24569 OR2X1_LOC_325/A OR2X1_LOC_502/A 0.11fF
C24570 OR2X1_LOC_744/A AND2X1_LOC_644/Y 0.02fF
C24571 OR2X1_LOC_426/B AND2X1_LOC_124/a_8_24# 0.03fF
C24572 D_INPUT_5 D_INPUT_4 0.95fF
C24573 AND2X1_LOC_556/a_8_24# OR2X1_LOC_427/A 0.01fF
C24574 OR2X1_LOC_864/a_8_216# D_GATE_662 0.14fF
C24575 OR2X1_LOC_177/Y OR2X1_LOC_485/A 0.03fF
C24576 OR2X1_LOC_27/a_8_216# AND2X1_LOC_219/A 0.07fF
C24577 OR2X1_LOC_8/Y OR2X1_LOC_85/A 0.32fF
C24578 OR2X1_LOC_404/Y OR2X1_LOC_576/A 0.03fF
C24579 AND2X1_LOC_567/a_8_24# AND2X1_LOC_661/A 0.17fF
C24580 AND2X1_LOC_50/Y AND2X1_LOC_752/a_36_24# 0.01fF
C24581 OR2X1_LOC_499/B OR2X1_LOC_833/B 0.05fF
C24582 OR2X1_LOC_845/a_8_216# OR2X1_LOC_66/A 0.01fF
C24583 OR2X1_LOC_449/B AND2X1_LOC_18/Y 0.00fF
C24584 AND2X1_LOC_474/A OR2X1_LOC_67/A 0.07fF
C24585 OR2X1_LOC_309/Y OR2X1_LOC_7/A 0.03fF
C24586 OR2X1_LOC_326/B OR2X1_LOC_325/a_8_216# 0.02fF
C24587 OR2X1_LOC_224/Y OR2X1_LOC_183/Y 0.79fF
C24588 OR2X1_LOC_346/a_8_216# OR2X1_LOC_78/A 0.01fF
C24589 VDD AND2X1_LOC_839/B 0.24fF
C24590 OR2X1_LOC_604/A OR2X1_LOC_665/Y 0.07fF
C24591 AND2X1_LOC_378/a_8_24# OR2X1_LOC_39/A 0.09fF
C24592 OR2X1_LOC_459/A OR2X1_LOC_459/B 0.15fF
C24593 OR2X1_LOC_196/Y AND2X1_LOC_48/A 0.04fF
C24594 AND2X1_LOC_784/A OR2X1_LOC_51/Y 0.07fF
C24595 AND2X1_LOC_560/a_8_24# AND2X1_LOC_227/Y 0.01fF
C24596 AND2X1_LOC_70/Y OR2X1_LOC_631/B 0.02fF
C24597 OR2X1_LOC_502/A OR2X1_LOC_847/A 0.03fF
C24598 OR2X1_LOC_251/Y OR2X1_LOC_494/Y 0.03fF
C24599 AND2X1_LOC_340/Y AND2X1_LOC_350/Y 0.03fF
C24600 OR2X1_LOC_160/A OR2X1_LOC_201/A 0.01fF
C24601 AND2X1_LOC_338/Y OR2X1_LOC_46/A 0.34fF
C24602 OR2X1_LOC_122/A OR2X1_LOC_44/Y 0.01fF
C24603 OR2X1_LOC_604/A OR2X1_LOC_485/A 1.10fF
C24604 AND2X1_LOC_12/Y AND2X1_LOC_316/a_8_24# 0.01fF
C24605 OR2X1_LOC_91/Y AND2X1_LOC_722/Y 0.03fF
C24606 OR2X1_LOC_139/A OR2X1_LOC_814/A 0.14fF
C24607 OR2X1_LOC_497/Y OR2X1_LOC_59/Y 0.07fF
C24608 AND2X1_LOC_88/a_8_24# AND2X1_LOC_18/Y 0.02fF
C24609 OR2X1_LOC_624/B OR2X1_LOC_772/A 0.01fF
C24610 INPUT_0 OR2X1_LOC_44/Y 0.18fF
C24611 OR2X1_LOC_314/a_8_216# AND2X1_LOC_452/Y 0.03fF
C24612 AND2X1_LOC_465/Y AND2X1_LOC_786/Y 0.01fF
C24613 OR2X1_LOC_103/Y AND2X1_LOC_113/Y 0.01fF
C24614 OR2X1_LOC_6/B AND2X1_LOC_122/a_8_24# 0.02fF
C24615 AND2X1_LOC_41/A OR2X1_LOC_193/Y 0.11fF
C24616 INPUT_0 OR2X1_LOC_82/a_36_216# 0.02fF
C24617 OR2X1_LOC_561/a_8_216# OR2X1_LOC_391/A -0.06fF
C24618 OR2X1_LOC_679/Y AND2X1_LOC_147/Y 0.00fF
C24619 AND2X1_LOC_753/B AND2X1_LOC_59/Y 0.07fF
C24620 OR2X1_LOC_185/Y OR2X1_LOC_435/a_8_216# 0.02fF
C24621 OR2X1_LOC_318/B OR2X1_LOC_723/B 0.02fF
C24622 AND2X1_LOC_342/Y OR2X1_LOC_92/Y 0.66fF
C24623 AND2X1_LOC_514/a_8_24# AND2X1_LOC_211/B 0.04fF
C24624 OR2X1_LOC_840/A AND2X1_LOC_153/a_36_24# 0.00fF
C24625 OR2X1_LOC_858/A OR2X1_LOC_296/a_8_216# 0.00fF
C24626 OR2X1_LOC_307/a_36_216# OR2X1_LOC_78/A 0.00fF
C24627 AND2X1_LOC_392/A AND2X1_LOC_211/a_36_24# 0.01fF
C24628 OR2X1_LOC_629/Y AND2X1_LOC_43/B 0.24fF
C24629 AND2X1_LOC_711/Y AND2X1_LOC_507/a_36_24# 0.01fF
C24630 OR2X1_LOC_154/A AND2X1_LOC_423/a_8_24# 0.01fF
C24631 OR2X1_LOC_744/A OR2X1_LOC_7/A 0.52fF
C24632 OR2X1_LOC_51/Y OR2X1_LOC_3/a_8_216# 0.01fF
C24633 OR2X1_LOC_421/a_8_216# OR2X1_LOC_52/B 0.03fF
C24634 AND2X1_LOC_36/Y OR2X1_LOC_598/A 0.35fF
C24635 OR2X1_LOC_13/B OR2X1_LOC_534/a_8_216# 0.03fF
C24636 OR2X1_LOC_241/Y AND2X1_LOC_7/B 0.56fF
C24637 OR2X1_LOC_330/Y AND2X1_LOC_56/B 0.02fF
C24638 OR2X1_LOC_18/Y OR2X1_LOC_616/a_8_216# 0.18fF
C24639 OR2X1_LOC_199/a_36_216# AND2X1_LOC_47/Y 0.00fF
C24640 OR2X1_LOC_3/Y OR2X1_LOC_816/Y 0.03fF
C24641 OR2X1_LOC_358/a_8_216# OR2X1_LOC_653/Y 0.03fF
C24642 OR2X1_LOC_479/Y OR2X1_LOC_78/A 0.16fF
C24643 OR2X1_LOC_405/A AND2X1_LOC_59/Y 0.10fF
C24644 AND2X1_LOC_711/Y AND2X1_LOC_865/A 0.03fF
C24645 OR2X1_LOC_774/Y OR2X1_LOC_391/a_8_216# 0.01fF
C24646 AND2X1_LOC_539/Y AND2X1_LOC_810/a_8_24# 0.01fF
C24647 AND2X1_LOC_70/Y AND2X1_LOC_135/a_8_24# 0.03fF
C24648 OR2X1_LOC_121/B AND2X1_LOC_18/Y 1.53fF
C24649 OR2X1_LOC_739/B OR2X1_LOC_221/a_8_216# 0.09fF
C24650 OR2X1_LOC_45/B AND2X1_LOC_476/A 0.08fF
C24651 AND2X1_LOC_76/Y OR2X1_LOC_85/A 0.10fF
C24652 AND2X1_LOC_729/B OR2X1_LOC_56/A 0.03fF
C24653 OR2X1_LOC_517/a_8_216# OR2X1_LOC_74/A 0.08fF
C24654 AND2X1_LOC_11/Y AND2X1_LOC_25/Y 1.05fF
C24655 OR2X1_LOC_541/B OR2X1_LOC_541/a_36_216# 0.00fF
C24656 AND2X1_LOC_214/A OR2X1_LOC_48/Y 0.06fF
C24657 AND2X1_LOC_794/A AND2X1_LOC_840/B 0.36fF
C24658 D_INPUT_1 OR2X1_LOC_121/A 0.03fF
C24659 OR2X1_LOC_682/Y OR2X1_LOC_92/Y 0.14fF
C24660 AND2X1_LOC_430/B INPUT_6 0.03fF
C24661 AND2X1_LOC_40/Y AND2X1_LOC_373/a_8_24# 0.01fF
C24662 VDD AND2X1_LOC_116/B 0.04fF
C24663 OR2X1_LOC_468/Y OR2X1_LOC_211/a_36_216# 0.00fF
C24664 AND2X1_LOC_580/B AND2X1_LOC_805/Y 0.03fF
C24665 AND2X1_LOC_12/Y OR2X1_LOC_865/Y 0.01fF
C24666 OR2X1_LOC_154/A OR2X1_LOC_405/Y 0.01fF
C24667 OR2X1_LOC_580/A OR2X1_LOC_366/Y 0.01fF
C24668 AND2X1_LOC_95/Y OR2X1_LOC_461/A 0.14fF
C24669 AND2X1_LOC_384/a_36_24# OR2X1_LOC_269/B 0.00fF
C24670 OR2X1_LOC_53/a_8_216# OR2X1_LOC_752/a_8_216# 0.47fF
C24671 OR2X1_LOC_654/A OR2X1_LOC_651/B 0.76fF
C24672 OR2X1_LOC_598/A OR2X1_LOC_334/A 0.03fF
C24673 AND2X1_LOC_40/Y OR2X1_LOC_333/B 0.04fF
C24674 OR2X1_LOC_335/A OR2X1_LOC_318/B 0.02fF
C24675 OR2X1_LOC_70/Y OR2X1_LOC_298/a_8_216# 0.05fF
C24676 OR2X1_LOC_58/Y OR2X1_LOC_412/a_36_216# 0.00fF
C24677 VDD OR2X1_LOC_404/A 0.04fF
C24678 OR2X1_LOC_864/A AND2X1_LOC_95/Y 1.23fF
C24679 AND2X1_LOC_566/B AND2X1_LOC_864/a_8_24# 0.01fF
C24680 AND2X1_LOC_353/a_8_24# AND2X1_LOC_863/Y 0.20fF
C24681 OR2X1_LOC_125/a_8_216# INPUT_1 0.04fF
C24682 OR2X1_LOC_51/Y AND2X1_LOC_639/A 0.17fF
C24683 AND2X1_LOC_859/Y AND2X1_LOC_862/A 0.00fF
C24684 OR2X1_LOC_22/A OR2X1_LOC_380/a_36_216# 0.00fF
C24685 AND2X1_LOC_859/Y AND2X1_LOC_624/A 0.07fF
C24686 OR2X1_LOC_812/B OR2X1_LOC_383/a_8_216# 0.05fF
C24687 OR2X1_LOC_40/Y OR2X1_LOC_31/Y 1.37fF
C24688 OR2X1_LOC_778/Y OR2X1_LOC_739/A 0.05fF
C24689 AND2X1_LOC_658/A AND2X1_LOC_678/a_8_24# 0.04fF
C24690 OR2X1_LOC_503/A OR2X1_LOC_44/Y 0.00fF
C24691 OR2X1_LOC_11/Y OR2X1_LOC_44/Y 0.79fF
C24692 OR2X1_LOC_185/A OR2X1_LOC_564/B 0.02fF
C24693 OR2X1_LOC_391/B OR2X1_LOC_848/B 0.11fF
C24694 OR2X1_LOC_687/Y OR2X1_LOC_87/A 0.07fF
C24695 OR2X1_LOC_772/B OR2X1_LOC_846/B 0.04fF
C24696 OR2X1_LOC_633/Y OR2X1_LOC_633/B 0.16fF
C24697 OR2X1_LOC_81/Y OR2X1_LOC_80/Y 0.06fF
C24698 OR2X1_LOC_821/a_8_216# OR2X1_LOC_813/Y 0.01fF
C24699 OR2X1_LOC_585/A AND2X1_LOC_655/A 0.02fF
C24700 AND2X1_LOC_778/a_8_24# OR2X1_LOC_680/A 0.03fF
C24701 OR2X1_LOC_160/A AND2X1_LOC_3/Y 0.27fF
C24702 OR2X1_LOC_793/a_8_216# OR2X1_LOC_793/B 0.01fF
C24703 OR2X1_LOC_495/a_8_216# OR2X1_LOC_36/Y 0.07fF
C24704 AND2X1_LOC_468/B OR2X1_LOC_74/A 0.02fF
C24705 OR2X1_LOC_160/A OR2X1_LOC_647/B 0.07fF
C24706 AND2X1_LOC_348/Y AND2X1_LOC_359/B 0.47fF
C24707 AND2X1_LOC_560/B OR2X1_LOC_44/Y 0.07fF
C24708 OR2X1_LOC_619/Y AND2X1_LOC_211/a_8_24# 0.05fF
C24709 OR2X1_LOC_604/A AND2X1_LOC_452/a_8_24# 0.01fF
C24710 AND2X1_LOC_21/a_8_24# D_INPUT_4 0.02fF
C24711 AND2X1_LOC_379/a_8_24# AND2X1_LOC_638/a_8_24# 0.23fF
C24712 AND2X1_LOC_580/A AND2X1_LOC_569/a_36_24# 0.00fF
C24713 OR2X1_LOC_686/B AND2X1_LOC_684/a_8_24# 0.25fF
C24714 OR2X1_LOC_85/A OR2X1_LOC_52/B 0.15fF
C24715 OR2X1_LOC_473/a_8_216# OR2X1_LOC_121/B 0.01fF
C24716 OR2X1_LOC_280/Y OR2X1_LOC_39/A 0.09fF
C24717 OR2X1_LOC_672/Y OR2X1_LOC_85/A 0.12fF
C24718 AND2X1_LOC_712/B OR2X1_LOC_92/Y 0.03fF
C24719 AND2X1_LOC_359/B OR2X1_LOC_753/A 0.10fF
C24720 OR2X1_LOC_690/A OR2X1_LOC_44/Y 0.08fF
C24721 OR2X1_LOC_481/A OR2X1_LOC_625/Y 0.02fF
C24722 AND2X1_LOC_11/Y AND2X1_LOC_51/Y 1.18fF
C24723 OR2X1_LOC_630/Y AND2X1_LOC_47/Y 0.80fF
C24724 OR2X1_LOC_81/a_8_216# OR2X1_LOC_585/A 0.02fF
C24725 OR2X1_LOC_92/Y OR2X1_LOC_54/Y 0.04fF
C24726 OR2X1_LOC_476/B OR2X1_LOC_61/Y 0.10fF
C24727 OR2X1_LOC_778/Y OR2X1_LOC_269/B 0.05fF
C24728 AND2X1_LOC_22/Y AND2X1_LOC_31/Y 1.36fF
C24729 AND2X1_LOC_339/B OR2X1_LOC_595/Y 0.00fF
C24730 OR2X1_LOC_607/A D_INPUT_1 0.01fF
C24731 AND2X1_LOC_852/Y AND2X1_LOC_853/Y 0.23fF
C24732 OR2X1_LOC_596/A OR2X1_LOC_194/a_36_216# 0.00fF
C24733 AND2X1_LOC_141/B OR2X1_LOC_65/B 0.04fF
C24734 OR2X1_LOC_850/B OR2X1_LOC_814/A 0.01fF
C24735 INPUT_5 AND2X1_LOC_25/a_8_24# 0.01fF
C24736 OR2X1_LOC_402/Y AND2X1_LOC_51/Y 0.18fF
C24737 OR2X1_LOC_744/A OR2X1_LOC_224/a_8_216# 0.02fF
C24738 OR2X1_LOC_673/Y AND2X1_LOC_79/Y 0.07fF
C24739 OR2X1_LOC_11/a_8_216# INPUT_7 0.01fF
C24740 AND2X1_LOC_93/a_8_24# OR2X1_LOC_99/A 0.09fF
C24741 OR2X1_LOC_426/B OR2X1_LOC_47/Y 0.04fF
C24742 OR2X1_LOC_83/Y AND2X1_LOC_84/a_8_24# 0.00fF
C24743 AND2X1_LOC_560/B AND2X1_LOC_116/Y 0.03fF
C24744 OR2X1_LOC_3/Y OR2X1_LOC_748/A 0.02fF
C24745 OR2X1_LOC_427/A OR2X1_LOC_77/a_8_216# 0.01fF
C24746 AND2X1_LOC_300/a_36_24# OR2X1_LOC_318/B 0.00fF
C24747 OR2X1_LOC_703/Y OR2X1_LOC_308/Y 0.03fF
C24748 VDD AND2X1_LOC_204/Y 0.01fF
C24749 OR2X1_LOC_70/Y OR2X1_LOC_86/Y 0.01fF
C24750 OR2X1_LOC_620/Y D_INPUT_0 0.06fF
C24751 OR2X1_LOC_385/Y OR2X1_LOC_387/Y 0.22fF
C24752 OR2X1_LOC_22/Y AND2X1_LOC_661/a_36_24# 0.02fF
C24753 D_INPUT_3 AND2X1_LOC_401/Y 0.51fF
C24754 AND2X1_LOC_95/Y AND2X1_LOC_134/a_36_24# 0.00fF
C24755 OR2X1_LOC_479/Y OR2X1_LOC_155/A 0.08fF
C24756 AND2X1_LOC_86/B AND2X1_LOC_3/Y 0.00fF
C24757 AND2X1_LOC_12/Y AND2X1_LOC_425/Y 0.48fF
C24758 OR2X1_LOC_22/Y OR2X1_LOC_39/A 0.12fF
C24759 AND2X1_LOC_12/Y AND2X1_LOC_309/a_8_24# 0.02fF
C24760 OR2X1_LOC_487/Y AND2X1_LOC_717/B 0.05fF
C24761 OR2X1_LOC_64/Y OR2X1_LOC_44/Y 2.70fF
C24762 AND2X1_LOC_169/a_8_24# AND2X1_LOC_841/B 0.00fF
C24763 AND2X1_LOC_44/Y OR2X1_LOC_366/Y 0.03fF
C24764 OR2X1_LOC_624/B AND2X1_LOC_3/Y 0.03fF
C24765 OR2X1_LOC_643/Y OR2X1_LOC_87/A 0.02fF
C24766 OR2X1_LOC_19/B OR2X1_LOC_82/a_8_216# 0.03fF
C24767 OR2X1_LOC_479/Y OR2X1_LOC_605/A 0.05fF
C24768 AND2X1_LOC_392/a_8_24# AND2X1_LOC_845/a_8_24# 0.23fF
C24769 OR2X1_LOC_630/Y OR2X1_LOC_598/A 0.01fF
C24770 OR2X1_LOC_154/A D_INPUT_0 0.59fF
C24771 OR2X1_LOC_3/Y OR2X1_LOC_304/Y 0.17fF
C24772 AND2X1_LOC_12/Y OR2X1_LOC_770/a_8_216# 0.01fF
C24773 OR2X1_LOC_424/a_8_216# OR2X1_LOC_31/Y 0.01fF
C24774 OR2X1_LOC_633/a_8_216# OR2X1_LOC_598/A 0.03fF
C24775 OR2X1_LOC_197/A OR2X1_LOC_375/A 0.04fF
C24776 AND2X1_LOC_443/Y AND2X1_LOC_222/Y -0.01fF
C24777 OR2X1_LOC_276/B OR2X1_LOC_203/a_8_216# 0.01fF
C24778 AND2X1_LOC_582/a_8_24# OR2X1_LOC_451/B 0.00fF
C24779 OR2X1_LOC_34/A AND2X1_LOC_36/Y 0.01fF
C24780 AND2X1_LOC_211/B OR2X1_LOC_22/Y 0.03fF
C24781 AND2X1_LOC_464/Y OR2X1_LOC_371/Y 0.04fF
C24782 OR2X1_LOC_278/A OR2X1_LOC_74/A 0.04fF
C24783 OR2X1_LOC_417/A OR2X1_LOC_44/Y 0.17fF
C24784 OR2X1_LOC_62/A OR2X1_LOC_375/A 0.61fF
C24785 AND2X1_LOC_648/B AND2X1_LOC_648/a_8_24# 0.11fF
C24786 OR2X1_LOC_78/A OR2X1_LOC_68/B 0.30fF
C24787 OR2X1_LOC_36/Y OR2X1_LOC_238/a_8_216# 0.01fF
C24788 OR2X1_LOC_55/a_8_216# OR2X1_LOC_6/A 0.01fF
C24789 OR2X1_LOC_425/a_8_216# OR2X1_LOC_70/A 0.01fF
C24790 AND2X1_LOC_627/a_36_24# AND2X1_LOC_36/Y 0.01fF
C24791 OR2X1_LOC_64/a_8_216# OR2X1_LOC_44/Y 0.01fF
C24792 AND2X1_LOC_578/A AND2X1_LOC_465/Y 0.03fF
C24793 OR2X1_LOC_95/Y AND2X1_LOC_361/A 0.11fF
C24794 OR2X1_LOC_26/Y AND2X1_LOC_675/A 0.20fF
C24795 AND2X1_LOC_47/Y OR2X1_LOC_346/B 0.01fF
C24796 OR2X1_LOC_178/a_8_216# OR2X1_LOC_437/A 0.04fF
C24797 OR2X1_LOC_473/Y OR2X1_LOC_476/a_8_216# 0.04fF
C24798 OR2X1_LOC_516/Y AND2X1_LOC_786/Y 0.07fF
C24799 OR2X1_LOC_291/Y OR2X1_LOC_277/a_8_216# 0.02fF
C24800 OR2X1_LOC_628/Y AND2X1_LOC_631/Y 0.02fF
C24801 AND2X1_LOC_367/a_8_24# OR2X1_LOC_47/Y 0.02fF
C24802 OR2X1_LOC_31/Y OR2X1_LOC_7/A 0.99fF
C24803 OR2X1_LOC_646/B AND2X1_LOC_36/Y 0.03fF
C24804 OR2X1_LOC_87/A OR2X1_LOC_786/Y 0.13fF
C24805 AND2X1_LOC_48/A AND2X1_LOC_46/a_8_24# 0.01fF
C24806 OR2X1_LOC_89/A AND2X1_LOC_675/A 0.12fF
C24807 OR2X1_LOC_596/A OR2X1_LOC_308/Y 0.10fF
C24808 AND2X1_LOC_40/Y OR2X1_LOC_567/a_36_216# 0.00fF
C24809 AND2X1_LOC_95/Y OR2X1_LOC_351/a_8_216# 0.01fF
C24810 OR2X1_LOC_213/a_36_216# OR2X1_LOC_375/A 0.00fF
C24811 OR2X1_LOC_247/a_36_216# OR2X1_LOC_805/A 0.02fF
C24812 AND2X1_LOC_681/a_8_24# OR2X1_LOC_155/A 0.06fF
C24813 OR2X1_LOC_331/A OR2X1_LOC_13/B 0.11fF
C24814 OR2X1_LOC_497/Y OR2X1_LOC_184/Y 0.03fF
C24815 OR2X1_LOC_130/A OR2X1_LOC_804/A 0.03fF
C24816 AND2X1_LOC_520/Y AND2X1_LOC_222/Y 0.04fF
C24817 OR2X1_LOC_31/Y OR2X1_LOC_44/a_8_216# 0.01fF
C24818 AND2X1_LOC_219/Y OR2X1_LOC_300/Y 0.03fF
C24819 OR2X1_LOC_62/a_8_216# OR2X1_LOC_54/Y 0.02fF
C24820 OR2X1_LOC_685/a_8_216# OR2X1_LOC_451/B 0.00fF
C24821 OR2X1_LOC_793/A OR2X1_LOC_801/B 0.16fF
C24822 OR2X1_LOC_85/A AND2X1_LOC_216/A 0.13fF
C24823 OR2X1_LOC_664/Y OR2X1_LOC_675/Y 0.21fF
C24824 OR2X1_LOC_743/A OR2X1_LOC_47/Y 0.03fF
C24825 OR2X1_LOC_86/a_36_216# OR2X1_LOC_67/Y 0.01fF
C24826 AND2X1_LOC_748/a_8_24# AND2X1_LOC_751/a_8_24# 0.23fF
C24827 OR2X1_LOC_711/B AND2X1_LOC_64/Y 0.01fF
C24828 OR2X1_LOC_599/Y OR2X1_LOC_585/A 0.04fF
C24829 OR2X1_LOC_507/A OR2X1_LOC_510/a_8_216# 0.01fF
C24830 OR2X1_LOC_508/a_8_216# OR2X1_LOC_392/B 0.13fF
C24831 OR2X1_LOC_440/B OR2X1_LOC_168/Y 0.01fF
C24832 AND2X1_LOC_344/a_8_24# OR2X1_LOC_437/A 0.02fF
C24833 INPUT_4 OR2X1_LOC_11/a_8_216# 0.26fF
C24834 OR2X1_LOC_243/B OR2X1_LOC_243/a_8_216# 0.05fF
C24835 AND2X1_LOC_44/Y OR2X1_LOC_389/a_8_216# 0.02fF
C24836 OR2X1_LOC_420/a_8_216# OR2X1_LOC_419/Y 0.01fF
C24837 AND2X1_LOC_719/Y AND2X1_LOC_564/B 0.10fF
C24838 OR2X1_LOC_296/Y OR2X1_LOC_247/a_36_216# 0.00fF
C24839 AND2X1_LOC_127/a_36_24# AND2X1_LOC_47/Y 0.00fF
C24840 OR2X1_LOC_335/a_8_216# OR2X1_LOC_160/B 0.06fF
C24841 OR2X1_LOC_12/Y OR2X1_LOC_381/a_8_216# 0.06fF
C24842 OR2X1_LOC_715/B OR2X1_LOC_97/A 0.05fF
C24843 OR2X1_LOC_53/Y VDD 0.17fF
C24844 OR2X1_LOC_786/A AND2X1_LOC_44/Y 0.04fF
C24845 OR2X1_LOC_47/Y OR2X1_LOC_246/A 0.05fF
C24846 OR2X1_LOC_267/Y OR2X1_LOC_66/A 0.02fF
C24847 AND2X1_LOC_122/a_8_24# OR2X1_LOC_598/A 0.01fF
C24848 OR2X1_LOC_155/A OR2X1_LOC_68/B 0.01fF
C24849 OR2X1_LOC_12/Y AND2X1_LOC_448/a_8_24# 0.01fF
C24850 AND2X1_LOC_64/Y OR2X1_LOC_324/B 0.03fF
C24851 OR2X1_LOC_40/Y AND2X1_LOC_213/B 0.03fF
C24852 OR2X1_LOC_600/A AND2X1_LOC_794/a_36_24# 0.00fF
C24853 OR2X1_LOC_640/Y AND2X1_LOC_7/B 0.01fF
C24854 OR2X1_LOC_6/B OR2X1_LOC_16/A 0.97fF
C24855 AND2X1_LOC_866/A AND2X1_LOC_270/a_8_24# 0.06fF
C24856 AND2X1_LOC_50/Y AND2X1_LOC_409/B 0.24fF
C24857 OR2X1_LOC_31/Y OR2X1_LOC_224/a_8_216# 0.02fF
C24858 OR2X1_LOC_139/A OR2X1_LOC_244/Y 0.01fF
C24859 VDD AND2X1_LOC_802/Y 0.01fF
C24860 AND2X1_LOC_12/Y OR2X1_LOC_723/B 0.03fF
C24861 AND2X1_LOC_50/Y AND2X1_LOC_763/B 0.01fF
C24862 AND2X1_LOC_712/Y OR2X1_LOC_421/Y 0.01fF
C24863 D_INPUT_0 AND2X1_LOC_6/a_8_24# 0.01fF
C24864 OR2X1_LOC_633/A OR2X1_LOC_66/A 0.03fF
C24865 OR2X1_LOC_506/A AND2X1_LOC_36/Y 0.13fF
C24866 AND2X1_LOC_721/Y OR2X1_LOC_329/B 0.03fF
C24867 OR2X1_LOC_161/A OR2X1_LOC_593/B 0.06fF
C24868 OR2X1_LOC_732/a_8_216# OR2X1_LOC_308/Y 0.03fF
C24869 AND2X1_LOC_60/a_8_24# AND2X1_LOC_92/Y 0.02fF
C24870 OR2X1_LOC_278/A AND2X1_LOC_647/Y 0.03fF
C24871 OR2X1_LOC_785/B OR2X1_LOC_390/B 0.00fF
C24872 AND2X1_LOC_675/a_8_24# OR2X1_LOC_95/Y 0.01fF
C24873 OR2X1_LOC_154/A OR2X1_LOC_339/A 0.01fF
C24874 OR2X1_LOC_36/Y OR2X1_LOC_376/Y 0.05fF
C24875 OR2X1_LOC_45/B INPUT_0 0.05fF
C24876 OR2X1_LOC_47/Y OR2X1_LOC_409/B 0.02fF
C24877 OR2X1_LOC_87/A OR2X1_LOC_181/Y 0.00fF
C24878 OR2X1_LOC_274/a_36_216# OR2X1_LOC_121/A 0.00fF
C24879 OR2X1_LOC_43/Y AND2X1_LOC_434/Y 0.08fF
C24880 AND2X1_LOC_64/Y AND2X1_LOC_142/a_8_24# 0.11fF
C24881 OR2X1_LOC_40/Y OR2X1_LOC_129/a_8_216# 0.01fF
C24882 VDD OR2X1_LOC_151/A 0.43fF
C24883 AND2X1_LOC_95/Y OR2X1_LOC_501/A 0.01fF
C24884 OR2X1_LOC_696/A OR2X1_LOC_250/Y 0.07fF
C24885 OR2X1_LOC_31/Y OR2X1_LOC_511/a_8_216# 0.07fF
C24886 OR2X1_LOC_528/Y OR2X1_LOC_600/A 0.03fF
C24887 OR2X1_LOC_216/A AND2X1_LOC_7/B 0.20fF
C24888 OR2X1_LOC_510/A OR2X1_LOC_507/A 0.30fF
C24889 AND2X1_LOC_64/Y AND2X1_LOC_314/a_8_24# 0.14fF
C24890 AND2X1_LOC_675/A AND2X1_LOC_804/a_8_24# 0.23fF
C24891 OR2X1_LOC_474/Y OR2X1_LOC_576/A 0.05fF
C24892 AND2X1_LOC_47/Y OR2X1_LOC_196/a_8_216# 0.01fF
C24893 OR2X1_LOC_160/B OR2X1_LOC_676/Y 0.07fF
C24894 OR2X1_LOC_604/A OR2X1_LOC_600/a_36_216# 0.00fF
C24895 AND2X1_LOC_94/a_8_24# OR2X1_LOC_397/Y 0.25fF
C24896 OR2X1_LOC_335/A AND2X1_LOC_12/Y 0.31fF
C24897 OR2X1_LOC_329/B OR2X1_LOC_482/Y 0.06fF
C24898 OR2X1_LOC_756/B OR2X1_LOC_390/A 0.05fF
C24899 OR2X1_LOC_549/Y OR2X1_LOC_565/a_8_216# 0.07fF
C24900 AND2X1_LOC_91/B OR2X1_LOC_739/A 0.03fF
C24901 OR2X1_LOC_45/B AND2X1_LOC_717/Y 0.00fF
C24902 AND2X1_LOC_620/Y AND2X1_LOC_623/a_8_24# 0.04fF
C24903 AND2X1_LOC_17/Y INPUT_6 0.06fF
C24904 OR2X1_LOC_208/A OR2X1_LOC_154/A 0.02fF
C24905 OR2X1_LOC_696/A OR2X1_LOC_36/Y 0.30fF
C24906 D_INPUT_0 OR2X1_LOC_560/A 0.02fF
C24907 OR2X1_LOC_773/B OR2X1_LOC_773/Y 0.16fF
C24908 OR2X1_LOC_8/Y OR2X1_LOC_51/Y 0.03fF
C24909 AND2X1_LOC_84/Y OR2X1_LOC_69/A 0.01fF
C24910 OR2X1_LOC_160/B OR2X1_LOC_834/A 0.06fF
C24911 OR2X1_LOC_417/A AND2X1_LOC_570/a_8_24# 0.08fF
C24912 AND2X1_LOC_72/B D_INPUT_1 0.03fF
C24913 OR2X1_LOC_164/Y AND2X1_LOC_476/Y 0.04fF
C24914 AND2X1_LOC_474/A AND2X1_LOC_244/a_8_24# 0.01fF
C24915 OR2X1_LOC_842/A OR2X1_LOC_287/A 0.16fF
C24916 AND2X1_LOC_658/B AND2X1_LOC_865/A 0.23fF
C24917 OR2X1_LOC_790/A AND2X1_LOC_693/a_36_24# -0.00fF
C24918 AND2X1_LOC_70/Y OR2X1_LOC_648/A 0.07fF
C24919 OR2X1_LOC_623/a_8_216# OR2X1_LOC_161/B 0.01fF
C24920 OR2X1_LOC_624/A AND2X1_LOC_44/Y 0.03fF
C24921 OR2X1_LOC_528/Y AND2X1_LOC_862/Y 0.04fF
C24922 OR2X1_LOC_696/A OR2X1_LOC_93/a_36_216# 0.00fF
C24923 AND2X1_LOC_705/Y OR2X1_LOC_48/B 0.09fF
C24924 AND2X1_LOC_212/Y AND2X1_LOC_808/a_8_24# 0.03fF
C24925 OR2X1_LOC_6/B OR2X1_LOC_274/Y 0.01fF
C24926 AND2X1_LOC_574/a_8_24# AND2X1_LOC_658/B 0.02fF
C24927 OR2X1_LOC_49/A OR2X1_LOC_38/a_8_216# 0.03fF
C24928 AND2X1_LOC_512/Y OR2X1_LOC_600/A 0.07fF
C24929 OR2X1_LOC_422/Y OR2X1_LOC_421/Y 0.10fF
C24930 OR2X1_LOC_457/B AND2X1_LOC_7/B 0.01fF
C24931 AND2X1_LOC_110/Y OR2X1_LOC_808/B 0.05fF
C24932 OR2X1_LOC_516/Y AND2X1_LOC_578/A 0.07fF
C24933 AND2X1_LOC_91/B OR2X1_LOC_269/B 0.70fF
C24934 AND2X1_LOC_51/Y OR2X1_LOC_593/B 0.03fF
C24935 AND2X1_LOC_363/B OR2X1_LOC_40/Y 0.01fF
C24936 OR2X1_LOC_447/Y OR2X1_LOC_317/B 0.04fF
C24937 AND2X1_LOC_571/A OR2X1_LOC_89/A 0.48fF
C24938 AND2X1_LOC_436/B OR2X1_LOC_16/A 0.02fF
C24939 OR2X1_LOC_166/a_8_216# AND2X1_LOC_512/Y 0.03fF
C24940 AND2X1_LOC_738/B AND2X1_LOC_513/a_8_24# 0.03fF
C24941 AND2X1_LOC_385/a_8_24# AND2X1_LOC_7/B 0.06fF
C24942 VDD OR2X1_LOC_651/B -0.00fF
C24943 OR2X1_LOC_175/Y OR2X1_LOC_810/A 0.00fF
C24944 OR2X1_LOC_864/A AND2X1_LOC_22/Y 0.10fF
C24945 OR2X1_LOC_114/a_8_216# OR2X1_LOC_632/Y 0.03fF
C24946 AND2X1_LOC_592/Y OR2X1_LOC_619/Y 0.03fF
C24947 OR2X1_LOC_421/A OR2X1_LOC_427/A 0.03fF
C24948 OR2X1_LOC_620/Y OR2X1_LOC_356/a_8_216# 0.01fF
C24949 OR2X1_LOC_856/B AND2X1_LOC_18/Y 0.07fF
C24950 OR2X1_LOC_664/Y OR2X1_LOC_736/Y 0.03fF
C24951 OR2X1_LOC_703/B OR2X1_LOC_535/A 0.05fF
C24952 AND2X1_LOC_563/A OR2X1_LOC_427/A 0.01fF
C24953 VDD OR2X1_LOC_628/a_8_216# 0.21fF
C24954 OR2X1_LOC_71/a_8_216# AND2X1_LOC_243/Y 0.04fF
C24955 AND2X1_LOC_42/B OR2X1_LOC_415/Y 0.06fF
C24956 AND2X1_LOC_391/Y OR2X1_LOC_256/Y 0.07fF
C24957 AND2X1_LOC_454/A OR2X1_LOC_428/A 0.39fF
C24958 OR2X1_LOC_810/A AND2X1_LOC_417/a_8_24# 0.24fF
C24959 AND2X1_LOC_22/Y OR2X1_LOC_633/B 0.03fF
C24960 AND2X1_LOC_743/a_8_24# AND2X1_LOC_3/Y 0.03fF
C24961 OR2X1_LOC_506/a_8_216# AND2X1_LOC_51/Y 0.02fF
C24962 OR2X1_LOC_474/Y AND2X1_LOC_41/A 0.03fF
C24963 OR2X1_LOC_485/Y OR2X1_LOC_39/A 0.05fF
C24964 OR2X1_LOC_154/A OR2X1_LOC_515/A 0.01fF
C24965 OR2X1_LOC_114/Y AND2X1_LOC_150/a_8_24# 0.16fF
C24966 AND2X1_LOC_658/B AND2X1_LOC_676/a_8_24# 0.03fF
C24967 AND2X1_LOC_47/Y OR2X1_LOC_374/a_8_216# 0.01fF
C24968 AND2X1_LOC_481/a_8_24# OR2X1_LOC_161/B 0.01fF
C24969 OR2X1_LOC_7/A AND2X1_LOC_213/B 0.07fF
C24970 OR2X1_LOC_47/Y OR2X1_LOC_599/a_8_216# 0.01fF
C24971 AND2X1_LOC_70/Y OR2X1_LOC_405/a_8_216# 0.01fF
C24972 AND2X1_LOC_728/Y OR2X1_LOC_679/a_8_216# 0.01fF
C24973 OR2X1_LOC_516/A OR2X1_LOC_600/A 0.17fF
C24974 AND2X1_LOC_98/Y AND2X1_LOC_99/Y 0.00fF
C24975 OR2X1_LOC_9/Y OR2X1_LOC_824/Y 0.04fF
C24976 AND2X1_LOC_847/Y OR2X1_LOC_700/a_8_216# 0.03fF
C24977 OR2X1_LOC_645/a_36_216# OR2X1_LOC_161/A 0.02fF
C24978 OR2X1_LOC_45/B OR2X1_LOC_273/a_36_216# 0.00fF
C24979 OR2X1_LOC_508/A OR2X1_LOC_474/Y 0.07fF
C24980 AND2X1_LOC_1/Y AND2X1_LOC_7/B 0.00fF
C24981 OR2X1_LOC_51/Y OR2X1_LOC_67/A 0.00fF
C24982 OR2X1_LOC_96/Y OR2X1_LOC_6/A 0.01fF
C24983 OR2X1_LOC_485/A AND2X1_LOC_212/Y 0.07fF
C24984 OR2X1_LOC_520/Y OR2X1_LOC_66/A 0.14fF
C24985 AND2X1_LOC_516/a_8_24# OR2X1_LOC_596/A 0.01fF
C24986 OR2X1_LOC_449/B OR2X1_LOC_307/A 0.03fF
C24987 AND2X1_LOC_65/a_8_24# OR2X1_LOC_231/A 0.20fF
C24988 OR2X1_LOC_175/Y OR2X1_LOC_857/a_8_216# 0.04fF
C24989 AND2X1_LOC_456/B OR2X1_LOC_427/A 0.06fF
C24990 AND2X1_LOC_59/Y AND2X1_LOC_19/Y 0.62fF
C24991 OR2X1_LOC_658/a_8_216# OR2X1_LOC_571/B 0.40fF
C24992 OR2X1_LOC_160/A INPUT_0 0.36fF
C24993 OR2X1_LOC_329/Y OR2X1_LOC_312/Y 0.02fF
C24994 OR2X1_LOC_45/B OR2X1_LOC_64/Y 0.38fF
C24995 OR2X1_LOC_165/a_36_216# AND2X1_LOC_723/Y 0.01fF
C24996 OR2X1_LOC_95/Y OR2X1_LOC_387/A 0.00fF
C24997 OR2X1_LOC_709/A AND2X1_LOC_136/a_8_24# 0.21fF
C24998 AND2X1_LOC_512/Y OR2X1_LOC_619/Y 0.43fF
C24999 OR2X1_LOC_369/a_36_216# AND2X1_LOC_784/A 0.01fF
C25000 AND2X1_LOC_512/Y AND2X1_LOC_356/a_8_24# 0.03fF
C25001 OR2X1_LOC_600/A AND2X1_LOC_105/a_8_24# 0.01fF
C25002 OR2X1_LOC_604/A OR2X1_LOC_420/a_8_216# 0.01fF
C25003 VDD OR2X1_LOC_191/B 0.30fF
C25004 OR2X1_LOC_376/A D_INPUT_5 0.04fF
C25005 AND2X1_LOC_350/B AND2X1_LOC_351/Y 0.01fF
C25006 OR2X1_LOC_226/a_8_216# OR2X1_LOC_184/a_8_216# 0.47fF
C25007 OR2X1_LOC_496/Y AND2X1_LOC_658/A 0.03fF
C25008 AND2X1_LOC_36/Y D_INPUT_1 8.61fF
C25009 OR2X1_LOC_595/Y OR2X1_LOC_300/Y 0.06fF
C25010 OR2X1_LOC_663/A OR2X1_LOC_137/B 0.03fF
C25011 AND2X1_LOC_539/Y OR2X1_LOC_167/Y 0.04fF
C25012 OR2X1_LOC_108/Y OR2X1_LOC_529/Y 0.16fF
C25013 OR2X1_LOC_49/A OR2X1_LOC_19/B 0.20fF
C25014 OR2X1_LOC_694/Y OR2X1_LOC_7/A 0.02fF
C25015 OR2X1_LOC_405/A OR2X1_LOC_623/B 0.03fF
C25016 OR2X1_LOC_51/Y OR2X1_LOC_52/B 0.70fF
C25017 AND2X1_LOC_474/A AND2X1_LOC_286/Y 0.00fF
C25018 OR2X1_LOC_51/Y OR2X1_LOC_672/Y 0.00fF
C25019 OR2X1_LOC_49/A OR2X1_LOC_606/a_36_216# 0.03fF
C25020 AND2X1_LOC_22/Y AND2X1_LOC_134/a_36_24# 0.01fF
C25021 OR2X1_LOC_861/a_8_216# OR2X1_LOC_865/B 0.04fF
C25022 AND2X1_LOC_732/B OR2X1_LOC_743/A 0.01fF
C25023 AND2X1_LOC_94/a_36_24# OR2X1_LOC_502/A 0.00fF
C25024 OR2X1_LOC_217/Y AND2X1_LOC_41/A 0.03fF
C25025 AND2X1_LOC_857/Y AND2X1_LOC_655/A 0.05fF
C25026 OR2X1_LOC_655/B AND2X1_LOC_7/B 0.03fF
C25027 OR2X1_LOC_216/A OR2X1_LOC_805/A 0.03fF
C25028 VDD AND2X1_LOC_154/Y 0.21fF
C25029 OR2X1_LOC_106/A OR2X1_LOC_56/A 0.16fF
C25030 OR2X1_LOC_215/Y OR2X1_LOC_475/B 0.02fF
C25031 AND2X1_LOC_59/Y D_INPUT_4 0.08fF
C25032 AND2X1_LOC_147/Y AND2X1_LOC_657/Y 0.38fF
C25033 AND2X1_LOC_366/a_8_24# OR2X1_LOC_485/A 0.01fF
C25034 GATE_366 OR2X1_LOC_292/Y 0.15fF
C25035 AND2X1_LOC_36/Y AND2X1_LOC_48/Y 0.02fF
C25036 OR2X1_LOC_447/Y AND2X1_LOC_44/Y 0.03fF
C25037 OR2X1_LOC_70/Y OR2X1_LOC_582/a_8_216# 0.40fF
C25038 OR2X1_LOC_154/A AND2X1_LOC_40/Y 0.40fF
C25039 AND2X1_LOC_566/a_36_24# OR2X1_LOC_91/A 0.00fF
C25040 OR2X1_LOC_45/B OR2X1_LOC_417/A 0.06fF
C25041 OR2X1_LOC_653/a_8_216# OR2X1_LOC_648/A 0.02fF
C25042 OR2X1_LOC_235/B AND2X1_LOC_102/a_8_24# 0.01fF
C25043 OR2X1_LOC_224/Y AND2X1_LOC_465/A 0.00fF
C25044 OR2X1_LOC_464/A OR2X1_LOC_719/Y 0.00fF
C25045 AND2X1_LOC_456/B AND2X1_LOC_363/A 0.00fF
C25046 AND2X1_LOC_344/a_8_24# AND2X1_LOC_348/Y 0.01fF
C25047 AND2X1_LOC_12/Y OR2X1_LOC_812/B 0.68fF
C25048 OR2X1_LOC_58/a_8_216# OR2X1_LOC_52/B 0.01fF
C25049 AND2X1_LOC_697/a_8_24# OR2X1_LOC_78/A 0.04fF
C25050 AND2X1_LOC_51/a_8_24# AND2X1_LOC_51/A 0.20fF
C25051 OR2X1_LOC_74/A AND2X1_LOC_443/Y 0.00fF
C25052 AND2X1_LOC_86/B INPUT_0 0.02fF
C25053 OR2X1_LOC_231/A OR2X1_LOC_130/A 0.06fF
C25054 AND2X1_LOC_344/a_8_24# OR2X1_LOC_753/A 0.01fF
C25055 AND2X1_LOC_811/a_8_24# AND2X1_LOC_811/B 0.04fF
C25056 OR2X1_LOC_45/B OR2X1_LOC_75/a_36_216# 0.01fF
C25057 OR2X1_LOC_851/A OR2X1_LOC_87/A 0.02fF
C25058 OR2X1_LOC_280/Y AND2X1_LOC_474/A 0.02fF
C25059 OR2X1_LOC_508/a_8_216# OR2X1_LOC_532/B 0.01fF
C25060 OR2X1_LOC_114/Y OR2X1_LOC_575/A 0.17fF
C25061 OR2X1_LOC_362/B OR2X1_LOC_805/A 0.30fF
C25062 OR2X1_LOC_696/A OR2X1_LOC_419/Y 0.02fF
C25063 OR2X1_LOC_548/A OR2X1_LOC_532/B 0.06fF
C25064 AND2X1_LOC_42/B OR2X1_LOC_632/Y 1.48fF
C25065 OR2X1_LOC_92/Y OR2X1_LOC_26/Y 0.44fF
C25066 OR2X1_LOC_532/B OR2X1_LOC_486/Y 0.09fF
C25067 OR2X1_LOC_417/Y AND2X1_LOC_447/Y 0.07fF
C25068 OR2X1_LOC_308/a_8_216# OR2X1_LOC_269/B 0.01fF
C25069 OR2X1_LOC_160/A OR2X1_LOC_128/a_8_216# 0.04fF
C25070 OR2X1_LOC_91/Y OR2X1_LOC_109/Y 0.18fF
C25071 AND2X1_LOC_215/Y AND2X1_LOC_334/a_8_24# 0.01fF
C25072 AND2X1_LOC_796/A OR2X1_LOC_142/Y 0.55fF
C25073 OR2X1_LOC_600/A OR2X1_LOC_54/Y 1.06fF
C25074 AND2X1_LOC_367/a_8_24# OR2X1_LOC_625/Y 0.02fF
C25075 OR2X1_LOC_87/A OR2X1_LOC_220/B 0.03fF
C25076 OR2X1_LOC_154/A OR2X1_LOC_537/A 0.01fF
C25077 OR2X1_LOC_130/A OR2X1_LOC_340/Y 0.02fF
C25078 OR2X1_LOC_131/Y OR2X1_LOC_517/A 0.01fF
C25079 OR2X1_LOC_377/A AND2X1_LOC_49/a_8_24# 0.04fF
C25080 AND2X1_LOC_349/B OR2X1_LOC_92/Y 0.07fF
C25081 OR2X1_LOC_92/Y OR2X1_LOC_89/A 0.11fF
C25082 OR2X1_LOC_416/A AND2X1_LOC_415/a_36_24# 0.00fF
C25083 AND2X1_LOC_577/Y AND2X1_LOC_580/A 0.20fF
C25084 OR2X1_LOC_375/A OR2X1_LOC_209/a_36_216# 0.00fF
C25085 AND2X1_LOC_684/a_36_24# OR2X1_LOC_161/B 0.00fF
C25086 AND2X1_LOC_734/Y OR2X1_LOC_70/Y 0.03fF
C25087 OR2X1_LOC_601/a_8_216# AND2X1_LOC_447/Y 0.12fF
C25088 VDD INPUT_1 0.98fF
C25089 OR2X1_LOC_9/Y OR2X1_LOC_95/Y 0.03fF
C25090 OR2X1_LOC_359/a_36_216# OR2X1_LOC_814/A 0.00fF
C25091 OR2X1_LOC_348/Y AND2X1_LOC_283/a_8_24# 0.04fF
C25092 AND2X1_LOC_59/Y OR2X1_LOC_673/Y 0.02fF
C25093 OR2X1_LOC_448/B AND2X1_LOC_697/a_8_24# 0.01fF
C25094 OR2X1_LOC_46/A OR2X1_LOC_56/A 0.49fF
C25095 AND2X1_LOC_808/A AND2X1_LOC_727/B 0.53fF
C25096 OR2X1_LOC_349/a_36_216# OR2X1_LOC_814/A 0.00fF
C25097 OR2X1_LOC_158/A AND2X1_LOC_476/A 0.05fF
C25098 AND2X1_LOC_717/B OR2X1_LOC_427/A 0.03fF
C25099 OR2X1_LOC_26/Y OR2X1_LOC_65/B 0.09fF
C25100 OR2X1_LOC_84/Y AND2X1_LOC_44/Y 0.03fF
C25101 OR2X1_LOC_847/A AND2X1_LOC_3/Y 0.03fF
C25102 OR2X1_LOC_257/a_8_216# OR2X1_LOC_89/A 0.06fF
C25103 OR2X1_LOC_696/A OR2X1_LOC_526/a_8_216# 0.06fF
C25104 AND2X1_LOC_174/a_36_24# OR2X1_LOC_52/B 0.00fF
C25105 OR2X1_LOC_687/Y OR2X1_LOC_800/a_8_216# 0.01fF
C25106 OR2X1_LOC_74/A AND2X1_LOC_520/Y 0.02fF
C25107 AND2X1_LOC_390/B AND2X1_LOC_841/B 0.07fF
C25108 OR2X1_LOC_271/B OR2X1_LOC_36/Y 0.01fF
C25109 OR2X1_LOC_791/A OR2X1_LOC_345/A 0.08fF
C25110 AND2X1_LOC_22/Y OR2X1_LOC_351/a_8_216# 0.09fF
C25111 OR2X1_LOC_756/B OR2X1_LOC_750/A 0.07fF
C25112 AND2X1_LOC_474/A OR2X1_LOC_22/Y 0.03fF
C25113 OR2X1_LOC_191/B OR2X1_LOC_223/B 1.02fF
C25114 AND2X1_LOC_51/Y OR2X1_LOC_574/a_8_216# 0.04fF
C25115 OR2X1_LOC_93/Y D_INPUT_3 0.01fF
C25116 OR2X1_LOC_84/B OR2X1_LOC_375/A 0.00fF
C25117 OR2X1_LOC_680/A OR2X1_LOC_52/B 0.10fF
C25118 AND2X1_LOC_336/a_8_24# AND2X1_LOC_436/B -0.02fF
C25119 OR2X1_LOC_685/a_8_216# OR2X1_LOC_687/B -0.00fF
C25120 OR2X1_LOC_89/A OR2X1_LOC_65/B 0.86fF
C25121 OR2X1_LOC_485/A AND2X1_LOC_447/a_8_24# 0.01fF
C25122 OR2X1_LOC_70/Y OR2X1_LOC_109/a_8_216# 0.03fF
C25123 OR2X1_LOC_373/Y AND2X1_LOC_405/a_8_24# 0.03fF
C25124 OR2X1_LOC_217/Y OR2X1_LOC_217/a_36_216# 0.00fF
C25125 VDD OR2X1_LOC_751/a_8_216# 0.21fF
C25126 OR2X1_LOC_756/B OR2X1_LOC_168/A 0.01fF
C25127 AND2X1_LOC_227/Y AND2X1_LOC_509/a_8_24# 0.10fF
C25128 OR2X1_LOC_98/A INPUT_1 0.01fF
C25129 OR2X1_LOC_481/a_36_216# AND2X1_LOC_847/Y 0.01fF
C25130 AND2X1_LOC_227/Y OR2X1_LOC_56/A 0.02fF
C25131 AND2X1_LOC_7/B OR2X1_LOC_750/Y 0.98fF
C25132 AND2X1_LOC_186/a_8_24# OR2X1_LOC_74/A 0.03fF
C25133 AND2X1_LOC_31/Y OR2X1_LOC_227/B 0.04fF
C25134 OR2X1_LOC_685/B AND2X1_LOC_3/Y 0.01fF
C25135 OR2X1_LOC_866/B OR2X1_LOC_561/B 0.31fF
C25136 AND2X1_LOC_53/Y AND2X1_LOC_693/a_8_24# 0.02fF
C25137 OR2X1_LOC_624/a_8_216# AND2X1_LOC_47/Y 0.01fF
C25138 OR2X1_LOC_209/A OR2X1_LOC_726/a_8_216# 0.24fF
C25139 AND2X1_LOC_44/Y OR2X1_LOC_513/a_8_216# 0.01fF
C25140 OR2X1_LOC_36/Y OR2X1_LOC_754/a_36_216# 0.02fF
C25141 AND2X1_LOC_791/a_36_24# AND2X1_LOC_789/Y 0.01fF
C25142 AND2X1_LOC_337/B AND2X1_LOC_661/A 0.14fF
C25143 AND2X1_LOC_712/B OR2X1_LOC_619/Y 0.01fF
C25144 OR2X1_LOC_91/A AND2X1_LOC_318/Y 0.02fF
C25145 OR2X1_LOC_357/B OR2X1_LOC_578/B 0.09fF
C25146 OR2X1_LOC_151/A OR2X1_LOC_140/a_8_216# 0.05fF
C25147 OR2X1_LOC_154/A OR2X1_LOC_475/Y 0.02fF
C25148 OR2X1_LOC_813/A AND2X1_LOC_266/a_8_24# 0.11fF
C25149 OR2X1_LOC_91/A AND2X1_LOC_864/a_36_24# 0.01fF
C25150 OR2X1_LOC_47/Y OR2X1_LOC_12/a_8_216# -0.00fF
C25151 OR2X1_LOC_744/A OR2X1_LOC_615/Y 0.07fF
C25152 OR2X1_LOC_183/a_36_216# OR2X1_LOC_183/Y 0.00fF
C25153 OR2X1_LOC_759/Y AND2X1_LOC_789/Y 0.02fF
C25154 OR2X1_LOC_619/Y OR2X1_LOC_54/Y 0.15fF
C25155 AND2X1_LOC_12/Y AND2X1_LOC_27/a_8_24# 0.01fF
C25156 OR2X1_LOC_3/Y OR2X1_LOC_117/Y 0.22fF
C25157 OR2X1_LOC_387/Y OR2X1_LOC_585/A 0.01fF
C25158 AND2X1_LOC_345/a_36_24# OR2X1_LOC_748/A 0.00fF
C25159 AND2X1_LOC_220/B AND2X1_LOC_740/a_8_24# 0.07fF
C25160 OR2X1_LOC_239/a_8_216# OR2X1_LOC_239/Y 0.01fF
C25161 OR2X1_LOC_185/A AND2X1_LOC_133/a_8_24# 0.02fF
C25162 OR2X1_LOC_630/Y D_INPUT_1 0.07fF
C25163 AND2X1_LOC_97/a_8_24# AND2X1_LOC_845/Y 0.04fF
C25164 OR2X1_LOC_247/a_8_216# OR2X1_LOC_78/A 0.01fF
C25165 OR2X1_LOC_633/a_8_216# D_INPUT_1 0.04fF
C25166 AND2X1_LOC_863/Y AND2X1_LOC_841/B 0.07fF
C25167 OR2X1_LOC_315/Y INPUT_1 0.36fF
C25168 AND2X1_LOC_95/Y OR2X1_LOC_288/A 0.02fF
C25169 OR2X1_LOC_488/a_8_216# OR2X1_LOC_7/A 0.01fF
C25170 OR2X1_LOC_22/Y OR2X1_LOC_85/A 0.30fF
C25171 OR2X1_LOC_598/Y OR2X1_LOC_198/A 0.02fF
C25172 AND2X1_LOC_849/A AND2X1_LOC_806/A 0.02fF
C25173 AND2X1_LOC_131/a_8_24# OR2X1_LOC_560/A 0.18fF
C25174 AND2X1_LOC_56/B OR2X1_LOC_46/A 0.48fF
C25175 AND2X1_LOC_374/a_8_24# OR2X1_LOC_47/Y 0.01fF
C25176 AND2X1_LOC_825/a_8_24# OR2X1_LOC_6/A 0.10fF
C25177 AND2X1_LOC_505/a_8_24# OR2X1_LOC_560/A 0.01fF
C25178 AND2X1_LOC_80/a_8_24# OR2X1_LOC_532/B 0.17fF
C25179 AND2X1_LOC_40/Y OR2X1_LOC_84/a_8_216# 0.03fF
C25180 OR2X1_LOC_128/B AND2X1_LOC_47/Y 0.02fF
C25181 OR2X1_LOC_709/A OR2X1_LOC_704/a_8_216# 0.04fF
C25182 OR2X1_LOC_101/a_8_216# AND2X1_LOC_88/Y 0.00fF
C25183 AND2X1_LOC_64/Y OR2X1_LOC_508/Y 0.07fF
C25184 OR2X1_LOC_7/Y OR2X1_LOC_6/A 0.00fF
C25185 OR2X1_LOC_640/a_8_216# AND2X1_LOC_47/Y 0.01fF
C25186 AND2X1_LOC_648/B OR2X1_LOC_48/B 0.04fF
C25187 AND2X1_LOC_31/Y OR2X1_LOC_741/Y 0.34fF
C25188 AND2X1_LOC_786/a_8_24# AND2X1_LOC_204/a_8_24# 0.23fF
C25189 AND2X1_LOC_576/Y OR2X1_LOC_71/Y 0.04fF
C25190 OR2X1_LOC_18/Y AND2X1_LOC_648/B 0.01fF
C25191 OR2X1_LOC_222/a_8_216# OR2X1_LOC_805/A 0.04fF
C25192 OR2X1_LOC_185/A OR2X1_LOC_223/A 0.14fF
C25193 OR2X1_LOC_651/A OR2X1_LOC_375/A 0.03fF
C25194 AND2X1_LOC_719/Y OR2X1_LOC_437/A 0.10fF
C25195 AND2X1_LOC_127/a_8_24# AND2X1_LOC_3/Y 0.11fF
C25196 OR2X1_LOC_96/B OR2X1_LOC_95/Y 0.41fF
C25197 OR2X1_LOC_43/A AND2X1_LOC_169/a_8_24# 0.01fF
C25198 OR2X1_LOC_329/Y OR2X1_LOC_13/B 0.03fF
C25199 OR2X1_LOC_427/A AND2X1_LOC_451/a_36_24# 0.00fF
C25200 OR2X1_LOC_255/a_36_216# OR2X1_LOC_585/A 0.00fF
C25201 AND2X1_LOC_639/A AND2X1_LOC_639/a_8_24# 0.03fF
C25202 OR2X1_LOC_3/Y OR2X1_LOC_815/A 0.01fF
C25203 OR2X1_LOC_291/A OR2X1_LOC_46/A 0.15fF
C25204 OR2X1_LOC_59/Y AND2X1_LOC_215/a_8_24# 0.04fF
C25205 OR2X1_LOC_647/Y OR2X1_LOC_121/B 0.03fF
C25206 OR2X1_LOC_485/A OR2X1_LOC_255/a_8_216# 0.01fF
C25207 OR2X1_LOC_479/Y OR2X1_LOC_814/A 0.03fF
C25208 OR2X1_LOC_311/Y AND2X1_LOC_729/B 0.12fF
C25209 AND2X1_LOC_95/Y AND2X1_LOC_72/B 1.48fF
C25210 OR2X1_LOC_702/a_8_216# OR2X1_LOC_446/B 0.01fF
C25211 INPUT_4 OR2X1_LOC_51/a_8_216# 0.00fF
C25212 VDD OR2X1_LOC_714/A -0.00fF
C25213 AND2X1_LOC_18/a_8_24# AND2X1_LOC_7/Y 0.00fF
C25214 OR2X1_LOC_416/A OR2X1_LOC_585/A 0.02fF
C25215 AND2X1_LOC_555/a_8_24# AND2X1_LOC_789/Y 0.01fF
C25216 OR2X1_LOC_517/A AND2X1_LOC_657/A 0.98fF
C25217 OR2X1_LOC_45/B OR2X1_LOC_110/a_36_216# 0.00fF
C25218 AND2X1_LOC_538/Y AND2X1_LOC_729/B 0.01fF
C25219 OR2X1_LOC_347/A OR2X1_LOC_346/A 0.01fF
C25220 OR2X1_LOC_429/Y OR2X1_LOC_428/a_8_216# 0.05fF
C25221 OR2X1_LOC_235/B OR2X1_LOC_71/A 0.56fF
C25222 OR2X1_LOC_826/a_8_216# INPUT_1 0.01fF
C25223 AND2X1_LOC_40/Y OR2X1_LOC_560/A 0.02fF
C25224 AND2X1_LOC_70/Y OR2X1_LOC_112/A 0.08fF
C25225 AND2X1_LOC_40/Y OR2X1_LOC_198/A 0.02fF
C25226 OR2X1_LOC_696/A OR2X1_LOC_177/Y 0.01fF
C25227 OR2X1_LOC_285/B OR2X1_LOC_286/B 0.10fF
C25228 OR2X1_LOC_486/a_8_216# OR2X1_LOC_532/B 0.01fF
C25229 AND2X1_LOC_110/Y OR2X1_LOC_703/Y 0.23fF
C25230 OR2X1_LOC_176/Y AND2X1_LOC_802/B 0.01fF
C25231 AND2X1_LOC_69/a_8_24# OR2X1_LOC_121/B 0.02fF
C25232 AND2X1_LOC_555/Y OR2X1_LOC_281/Y 0.01fF
C25233 OR2X1_LOC_203/Y OR2X1_LOC_66/Y 0.01fF
C25234 OR2X1_LOC_43/A OR2X1_LOC_41/a_8_216# 0.02fF
C25235 OR2X1_LOC_572/a_36_216# OR2X1_LOC_576/A 0.00fF
C25236 OR2X1_LOC_696/A OR2X1_LOC_604/A 0.29fF
C25237 AND2X1_LOC_64/Y OR2X1_LOC_509/a_8_216# 0.11fF
C25238 OR2X1_LOC_555/B OR2X1_LOC_345/a_36_216# 0.03fF
C25239 OR2X1_LOC_744/A D_INPUT_6 0.00fF
C25240 OR2X1_LOC_520/Y OR2X1_LOC_559/a_8_216# 0.10fF
C25241 AND2X1_LOC_624/A AND2X1_LOC_657/A 0.07fF
C25242 OR2X1_LOC_121/Y OR2X1_LOC_139/A 0.10fF
C25243 OR2X1_LOC_278/A OR2X1_LOC_607/Y 0.11fF
C25244 AND2X1_LOC_552/a_8_24# AND2X1_LOC_476/Y 0.03fF
C25245 OR2X1_LOC_22/Y OR2X1_LOC_226/Y 0.01fF
C25246 AND2X1_LOC_57/Y AND2X1_LOC_70/Y 0.00fF
C25247 OR2X1_LOC_715/B OR2X1_LOC_175/Y 0.18fF
C25248 AND2X1_LOC_15/a_8_24# OR2X1_LOC_532/B 0.01fF
C25249 AND2X1_LOC_803/B AND2X1_LOC_209/Y 0.01fF
C25250 OR2X1_LOC_294/Y OR2X1_LOC_161/B 0.07fF
C25251 OR2X1_LOC_346/A AND2X1_LOC_44/Y 0.01fF
C25252 AND2X1_LOC_773/Y AND2X1_LOC_339/B 0.03fF
C25253 OR2X1_LOC_78/A AND2X1_LOC_235/a_8_24# 0.05fF
C25254 AND2X1_LOC_64/Y OR2X1_LOC_66/A 0.22fF
C25255 AND2X1_LOC_334/Y OR2X1_LOC_171/Y 0.02fF
C25256 OR2X1_LOC_426/B OR2X1_LOC_767/Y 0.24fF
C25257 AND2X1_LOC_810/B AND2X1_LOC_809/a_36_24# 0.01fF
C25258 AND2X1_LOC_715/Y OR2X1_LOC_604/A 0.14fF
C25259 AND2X1_LOC_91/B OR2X1_LOC_832/a_36_216# 0.01fF
C25260 AND2X1_LOC_41/A OR2X1_LOC_776/A 0.17fF
C25261 OR2X1_LOC_808/A OR2X1_LOC_301/a_8_216# 0.03fF
C25262 AND2X1_LOC_704/a_8_24# OR2X1_LOC_12/Y 0.01fF
C25263 OR2X1_LOC_161/A OR2X1_LOC_501/a_8_216# 0.01fF
C25264 OR2X1_LOC_715/B AND2X1_LOC_417/a_8_24# 0.04fF
C25265 OR2X1_LOC_715/B OR2X1_LOC_691/Y 0.03fF
C25266 AND2X1_LOC_223/A AND2X1_LOC_222/Y 0.01fF
C25267 OR2X1_LOC_739/A OR2X1_LOC_728/a_8_216# 0.01fF
C25268 OR2X1_LOC_68/a_8_216# OR2X1_LOC_68/B 0.04fF
C25269 AND2X1_LOC_655/A OR2X1_LOC_437/A 0.10fF
C25270 OR2X1_LOC_641/A OR2X1_LOC_161/B 0.29fF
C25271 AND2X1_LOC_252/a_8_24# OR2X1_LOC_578/B 0.02fF
C25272 AND2X1_LOC_92/Y OR2X1_LOC_703/a_8_216# 0.02fF
C25273 OR2X1_LOC_541/B OR2X1_LOC_777/B 0.13fF
C25274 OR2X1_LOC_737/A AND2X1_LOC_36/Y 0.07fF
C25275 AND2X1_LOC_800/a_8_24# OR2X1_LOC_760/Y 0.06fF
C25276 OR2X1_LOC_121/B OR2X1_LOC_804/A 0.30fF
C25277 AND2X1_LOC_18/Y OR2X1_LOC_578/a_8_216# 0.01fF
C25278 OR2X1_LOC_532/B AND2X1_LOC_109/a_8_24# 0.05fF
C25279 AND2X1_LOC_462/Y AND2X1_LOC_472/a_8_24# 0.09fF
C25280 OR2X1_LOC_744/A AND2X1_LOC_242/B 0.15fF
C25281 AND2X1_LOC_212/A AND2X1_LOC_566/B 0.02fF
C25282 OR2X1_LOC_850/B OR2X1_LOC_363/a_8_216# 0.01fF
C25283 OR2X1_LOC_269/B OR2X1_LOC_446/B 0.14fF
C25284 AND2X1_LOC_95/Y AND2X1_LOC_36/Y 0.50fF
C25285 OR2X1_LOC_629/B OR2X1_LOC_549/A 0.01fF
C25286 OR2X1_LOC_633/Y AND2X1_LOC_36/Y 0.10fF
C25287 AND2X1_LOC_702/Y OR2X1_LOC_13/B 0.03fF
C25288 AND2X1_LOC_544/Y OR2X1_LOC_441/a_36_216# 0.00fF
C25289 OR2X1_LOC_269/B OR2X1_LOC_303/B 0.03fF
C25290 OR2X1_LOC_139/A OR2X1_LOC_538/A 0.03fF
C25291 OR2X1_LOC_427/A AND2X1_LOC_439/a_36_24# 0.01fF
C25292 VDD AND2X1_LOC_300/a_8_24# 0.00fF
C25293 VDD AND2X1_LOC_130/a_8_24# 0.00fF
C25294 OR2X1_LOC_831/a_8_216# OR2X1_LOC_593/B 0.01fF
C25295 OR2X1_LOC_347/A OR2X1_LOC_161/A 0.01fF
C25296 OR2X1_LOC_862/a_8_216# OR2X1_LOC_862/A 0.08fF
C25297 AND2X1_LOC_326/B AND2X1_LOC_476/Y 0.02fF
C25298 OR2X1_LOC_358/B OR2X1_LOC_539/B 0.02fF
C25299 OR2X1_LOC_186/Y OR2X1_LOC_78/B 0.12fF
C25300 AND2X1_LOC_594/a_8_24# OR2X1_LOC_78/A 0.02fF
C25301 AND2X1_LOC_95/Y OR2X1_LOC_333/a_8_216# 0.03fF
C25302 OR2X1_LOC_389/B OR2X1_LOC_537/a_8_216# 0.47fF
C25303 OR2X1_LOC_858/a_8_216# OR2X1_LOC_362/A 0.01fF
C25304 OR2X1_LOC_31/Y AND2X1_LOC_203/Y 0.03fF
C25305 OR2X1_LOC_51/Y OR2X1_LOC_584/Y 0.01fF
C25306 VDD AND2X1_LOC_778/Y 0.30fF
C25307 OR2X1_LOC_227/Y OR2X1_LOC_340/a_8_216# 0.18fF
C25308 AND2X1_LOC_95/Y OR2X1_LOC_334/A 0.00fF
C25309 OR2X1_LOC_3/Y OR2X1_LOC_399/Y 0.02fF
C25310 AND2X1_LOC_86/a_8_24# OR2X1_LOC_66/A 0.01fF
C25311 OR2X1_LOC_51/Y OR2X1_LOC_253/Y 0.02fF
C25312 OR2X1_LOC_696/A OR2X1_LOC_306/Y 0.00fF
C25313 VDD AND2X1_LOC_709/a_8_24# 0.00fF
C25314 AND2X1_LOC_571/A AND2X1_LOC_576/a_8_24# 0.09fF
C25315 OR2X1_LOC_99/Y AND2X1_LOC_36/Y 0.15fF
C25316 OR2X1_LOC_158/A INPUT_0 0.33fF
C25317 AND2X1_LOC_677/a_36_24# OR2X1_LOC_779/B -0.00fF
C25318 OR2X1_LOC_18/Y AND2X1_LOC_465/A 0.06fF
C25319 AND2X1_LOC_471/Y AND2X1_LOC_476/Y 0.21fF
C25320 AND2X1_LOC_51/Y OR2X1_LOC_317/B 0.02fF
C25321 OR2X1_LOC_814/A OR2X1_LOC_68/B 0.09fF
C25322 OR2X1_LOC_695/Y AND2X1_LOC_707/a_8_24# 0.23fF
C25323 OR2X1_LOC_832/a_8_216# OR2X1_LOC_648/A 0.04fF
C25324 VDD AND2X1_LOC_352/B 0.11fF
C25325 OR2X1_LOC_624/a_36_216# OR2X1_LOC_113/B 0.00fF
C25326 AND2X1_LOC_64/Y OR2X1_LOC_799/a_36_216# 0.02fF
C25327 AND2X1_LOC_40/Y OR2X1_LOC_435/A 0.00fF
C25328 AND2X1_LOC_522/a_8_24# OR2X1_LOC_523/Y 0.00fF
C25329 OR2X1_LOC_787/Y OR2X1_LOC_593/B 0.05fF
C25330 OR2X1_LOC_18/Y AND2X1_LOC_231/a_8_24# 0.05fF
C25331 AND2X1_LOC_658/B AND2X1_LOC_658/Y 0.37fF
C25332 AND2X1_LOC_51/Y OR2X1_LOC_580/A 0.09fF
C25333 OR2X1_LOC_485/A OR2X1_LOC_183/a_8_216# 0.01fF
C25334 VDD OR2X1_LOC_287/A 0.17fF
C25335 OR2X1_LOC_769/A VDD 0.21fF
C25336 OR2X1_LOC_160/A AND2X1_LOC_7/B 5.29fF
C25337 OR2X1_LOC_45/B AND2X1_LOC_550/A 0.02fF
C25338 OR2X1_LOC_337/a_36_216# OR2X1_LOC_182/B 0.00fF
C25339 AND2X1_LOC_12/Y OR2X1_LOC_139/A 0.03fF
C25340 AND2X1_LOC_161/Y OR2X1_LOC_51/Y 0.01fF
C25341 OR2X1_LOC_747/Y AND2X1_LOC_782/a_8_24# 0.23fF
C25342 OR2X1_LOC_161/A AND2X1_LOC_44/Y 0.30fF
C25343 OR2X1_LOC_154/A OR2X1_LOC_138/a_8_216# 0.06fF
C25344 OR2X1_LOC_362/B OR2X1_LOC_580/B 0.12fF
C25345 AND2X1_LOC_544/a_36_24# AND2X1_LOC_476/Y 0.00fF
C25346 OR2X1_LOC_620/Y OR2X1_LOC_356/A 0.27fF
C25347 OR2X1_LOC_744/Y OR2X1_LOC_39/A 0.23fF
C25348 OR2X1_LOC_443/a_8_216# OR2X1_LOC_367/B 0.69fF
C25349 OR2X1_LOC_114/B OR2X1_LOC_850/B 0.81fF
C25350 VDD OR2X1_LOC_517/A 0.15fF
C25351 OR2X1_LOC_613/Y GATE_579 0.03fF
C25352 AND2X1_LOC_658/B AND2X1_LOC_734/Y 0.14fF
C25353 AND2X1_LOC_757/a_8_24# VDD -0.00fF
C25354 AND2X1_LOC_2/Y AND2X1_LOC_3/a_8_24# 0.01fF
C25355 AND2X1_LOC_542/a_36_24# OR2X1_LOC_427/A -0.00fF
C25356 AND2X1_LOC_48/Y OR2X1_LOC_196/a_8_216# 0.47fF
C25357 AND2X1_LOC_526/a_8_24# OR2X1_LOC_78/A 0.01fF
C25358 AND2X1_LOC_25/Y AND2X1_LOC_44/Y 0.04fF
C25359 AND2X1_LOC_738/B AND2X1_LOC_722/A 0.07fF
C25360 OR2X1_LOC_864/A OR2X1_LOC_227/B 0.03fF
C25361 OR2X1_LOC_309/Y AND2X1_LOC_841/B 0.03fF
C25362 VDD AND2X1_LOC_619/B 0.24fF
C25363 OR2X1_LOC_189/Y AND2X1_LOC_220/B 0.03fF
C25364 OR2X1_LOC_678/a_8_216# AND2X1_LOC_41/A 0.02fF
C25365 AND2X1_LOC_563/a_36_24# OR2X1_LOC_595/A 0.01fF
C25366 OR2X1_LOC_589/A OR2X1_LOC_316/Y 0.02fF
C25367 AND2X1_LOC_42/B OR2X1_LOC_397/a_36_216# 0.02fF
C25368 OR2X1_LOC_508/a_36_216# OR2X1_LOC_375/A 0.00fF
C25369 OR2X1_LOC_114/Y OR2X1_LOC_161/B 0.02fF
C25370 OR2X1_LOC_287/B OR2X1_LOC_362/a_36_216# 0.00fF
C25371 OR2X1_LOC_152/Y AND2X1_LOC_220/B 0.07fF
C25372 OR2X1_LOC_158/A OR2X1_LOC_11/Y 0.03fF
C25373 OR2X1_LOC_833/Y OR2X1_LOC_203/Y 0.01fF
C25374 OR2X1_LOC_31/Y OR2X1_LOC_424/Y 0.01fF
C25375 OR2X1_LOC_449/A OR2X1_LOC_161/B 0.06fF
C25376 OR2X1_LOC_304/a_8_216# OR2X1_LOC_485/A 0.01fF
C25377 OR2X1_LOC_165/a_8_216# OR2X1_LOC_51/Y 0.13fF
C25378 AND2X1_LOC_91/B AND2X1_LOC_176/a_8_24# 0.06fF
C25379 OR2X1_LOC_579/B OR2X1_LOC_349/A 0.08fF
C25380 D_INPUT_5 OR2X1_LOC_637/Y 0.02fF
C25381 OR2X1_LOC_377/A AND2X1_LOC_387/a_8_24# 0.03fF
C25382 INPUT_1 AND2X1_LOC_269/a_8_24# 0.02fF
C25383 AND2X1_LOC_848/Y AND2X1_LOC_860/A 0.14fF
C25384 OR2X1_LOC_158/A AND2X1_LOC_560/B 0.03fF
C25385 OR2X1_LOC_744/A AND2X1_LOC_841/B 8.65fF
C25386 VDD AND2X1_LOC_624/A 0.39fF
C25387 OR2X1_LOC_604/A AND2X1_LOC_458/Y 0.26fF
C25388 AND2X1_LOC_425/Y AND2X1_LOC_582/B 0.01fF
C25389 OR2X1_LOC_532/B OR2X1_LOC_308/Y 0.03fF
C25390 OR2X1_LOC_40/Y AND2X1_LOC_303/B 0.03fF
C25391 OR2X1_LOC_31/Y D_INPUT_6 0.03fF
C25392 OR2X1_LOC_7/A OR2X1_LOC_522/Y 0.14fF
C25393 OR2X1_LOC_269/B OR2X1_LOC_719/B 0.02fF
C25394 OR2X1_LOC_84/B OR2X1_LOC_549/A 0.00fF
C25395 OR2X1_LOC_158/A OR2X1_LOC_690/A 0.04fF
C25396 INPUT_0 OR2X1_LOC_847/A 0.04fF
C25397 OR2X1_LOC_468/A OR2X1_LOC_130/A 0.00fF
C25398 VDD OR2X1_LOC_380/A 0.03fF
C25399 AND2X1_LOC_392/A OR2X1_LOC_36/Y 6.90fF
C25400 AND2X1_LOC_310/a_8_24# OR2X1_LOC_375/A 0.01fF
C25401 OR2X1_LOC_51/Y OR2X1_LOC_48/a_8_216# 0.06fF
C25402 OR2X1_LOC_502/A OR2X1_LOC_608/a_8_216# 0.01fF
C25403 AND2X1_LOC_51/Y AND2X1_LOC_44/Y 0.23fF
C25404 OR2X1_LOC_773/B OR2X1_LOC_78/B 0.01fF
C25405 OR2X1_LOC_633/Y OR2X1_LOC_633/a_8_216# 0.01fF
C25406 AND2X1_LOC_197/a_8_24# AND2X1_LOC_219/A 0.20fF
C25407 OR2X1_LOC_51/Y AND2X1_LOC_286/Y 0.01fF
C25408 AND2X1_LOC_8/Y INPUT_2 0.01fF
C25409 OR2X1_LOC_600/A OR2X1_LOC_26/Y 0.77fF
C25410 OR2X1_LOC_703/B OR2X1_LOC_78/A 0.01fF
C25411 INPUT_3 AND2X1_LOC_820/B 0.05fF
C25412 OR2X1_LOC_589/A AND2X1_LOC_390/B 0.07fF
C25413 AND2X1_LOC_56/B OR2X1_LOC_702/a_8_216# 0.04fF
C25414 AND2X1_LOC_863/a_8_24# OR2X1_LOC_48/B 0.02fF
C25415 AND2X1_LOC_474/A OR2X1_LOC_39/A 0.05fF
C25416 AND2X1_LOC_10/a_36_24# OR2X1_LOC_161/B 0.00fF
C25417 OR2X1_LOC_542/B OR2X1_LOC_269/B 0.01fF
C25418 AND2X1_LOC_738/B OR2X1_LOC_599/A 0.41fF
C25419 AND2X1_LOC_81/B OR2X1_LOC_78/B 0.01fF
C25420 OR2X1_LOC_549/Y OR2X1_LOC_569/a_8_216# 0.14fF
C25421 AND2X1_LOC_810/A AND2X1_LOC_856/B 0.00fF
C25422 OR2X1_LOC_87/A OR2X1_LOC_78/A 0.25fF
C25423 AND2X1_LOC_49/a_8_24# OR2X1_LOC_78/B 0.04fF
C25424 OR2X1_LOC_78/B OR2X1_LOC_358/B 0.03fF
C25425 AND2X1_LOC_537/Y AND2X1_LOC_407/a_8_24# 0.19fF
C25426 OR2X1_LOC_185/A OR2X1_LOC_502/A 0.31fF
C25427 OR2X1_LOC_45/B OR2X1_LOC_268/a_36_216# 0.00fF
C25428 OR2X1_LOC_185/Y OR2X1_LOC_632/Y 0.10fF
C25429 OR2X1_LOC_677/Y AND2X1_LOC_624/A 0.15fF
C25430 OR2X1_LOC_319/B OR2X1_LOC_160/A 0.00fF
C25431 OR2X1_LOC_600/A OR2X1_LOC_89/A 0.10fF
C25432 AND2X1_LOC_663/A OR2X1_LOC_44/Y 0.03fF
C25433 AND2X1_LOC_810/A AND2X1_LOC_863/A 0.01fF
C25434 AND2X1_LOC_209/a_8_24# OR2X1_LOC_152/Y 0.01fF
C25435 OR2X1_LOC_325/a_8_216# AND2X1_LOC_95/Y 0.02fF
C25436 OR2X1_LOC_786/Y OR2X1_LOC_130/a_8_216# 0.01fF
C25437 AND2X1_LOC_12/Y OR2X1_LOC_850/B 0.02fF
C25438 OR2X1_LOC_629/a_8_216# OR2X1_LOC_629/B 0.00fF
C25439 AND2X1_LOC_696/a_8_24# OR2X1_LOC_78/A 0.01fF
C25440 OR2X1_LOC_622/A OR2X1_LOC_622/a_8_216# 0.02fF
C25441 OR2X1_LOC_621/a_8_216# OR2X1_LOC_624/B 0.01fF
C25442 OR2X1_LOC_405/A OR2X1_LOC_653/Y 0.13fF
C25443 OR2X1_LOC_158/A OR2X1_LOC_64/Y 0.15fF
C25444 OR2X1_LOC_600/A OR2X1_LOC_820/Y 0.23fF
C25445 OR2X1_LOC_31/Y AND2X1_LOC_242/B 0.02fF
C25446 OR2X1_LOC_359/A OR2X1_LOC_287/B 0.01fF
C25447 OR2X1_LOC_154/A AND2X1_LOC_39/a_8_24# 0.04fF
C25448 AND2X1_LOC_544/Y AND2X1_LOC_811/Y 0.00fF
C25449 OR2X1_LOC_280/Y OR2X1_LOC_51/Y 0.12fF
C25450 AND2X1_LOC_803/B AND2X1_LOC_728/a_8_24# 0.01fF
C25451 AND2X1_LOC_523/a_8_24# OR2X1_LOC_18/Y 0.03fF
C25452 AND2X1_LOC_81/B OR2X1_LOC_721/Y 0.05fF
C25453 OR2X1_LOC_427/A AND2X1_LOC_452/Y 0.01fF
C25454 OR2X1_LOC_121/B AND2X1_LOC_607/a_36_24# 0.00fF
C25455 OR2X1_LOC_617/a_36_216# OR2X1_LOC_627/Y 0.00fF
C25456 OR2X1_LOC_617/Y OR2X1_LOC_626/Y 0.16fF
C25457 OR2X1_LOC_89/A AND2X1_LOC_296/a_8_24# 0.01fF
C25458 AND2X1_LOC_707/Y OR2X1_LOC_31/Y 0.05fF
C25459 OR2X1_LOC_473/A OR2X1_LOC_115/B 0.09fF
C25460 AND2X1_LOC_191/B OR2X1_LOC_3/Y 0.03fF
C25461 OR2X1_LOC_620/Y AND2X1_LOC_43/B 0.07fF
C25462 OR2X1_LOC_604/A AND2X1_LOC_663/B 0.07fF
C25463 OR2X1_LOC_825/a_36_216# OR2X1_LOC_600/A 0.00fF
C25464 AND2X1_LOC_566/B AND2X1_LOC_727/A 0.00fF
C25465 AND2X1_LOC_787/A OR2X1_LOC_95/Y 0.03fF
C25466 AND2X1_LOC_787/A AND2X1_LOC_440/a_8_24# 0.01fF
C25467 AND2X1_LOC_560/B OR2X1_LOC_103/Y 0.23fF
C25468 OR2X1_LOC_619/Y AND2X1_LOC_453/Y 0.00fF
C25469 OR2X1_LOC_813/A OR2X1_LOC_595/A 0.00fF
C25470 OR2X1_LOC_216/a_8_216# OR2X1_LOC_78/A 0.01fF
C25471 AND2X1_LOC_90/a_8_24# OR2X1_LOC_532/B 0.01fF
C25472 OR2X1_LOC_166/Y AND2X1_LOC_390/B 0.02fF
C25473 AND2X1_LOC_351/a_8_24# OR2X1_LOC_31/Y 0.04fF
C25474 OR2X1_LOC_251/Y OR2X1_LOC_517/A 0.03fF
C25475 AND2X1_LOC_347/B OR2X1_LOC_295/Y 0.79fF
C25476 AND2X1_LOC_3/Y OR2X1_LOC_78/Y 0.02fF
C25477 OR2X1_LOC_799/A OR2X1_LOC_539/Y 0.16fF
C25478 OR2X1_LOC_179/a_8_216# OR2X1_LOC_7/A 0.02fF
C25479 OR2X1_LOC_377/A OR2X1_LOC_39/A 0.03fF
C25480 OR2X1_LOC_604/A AND2X1_LOC_686/a_8_24# 0.01fF
C25481 OR2X1_LOC_160/A OR2X1_LOC_805/A 0.14fF
C25482 OR2X1_LOC_616/Y AND2X1_LOC_624/A 0.03fF
C25483 OR2X1_LOC_864/A OR2X1_LOC_509/A 0.10fF
C25484 OR2X1_LOC_485/A OR2X1_LOC_164/Y 0.03fF
C25485 OR2X1_LOC_773/B OR2X1_LOC_375/A 0.08fF
C25486 OR2X1_LOC_757/A OR2X1_LOC_755/A 0.04fF
C25487 AND2X1_LOC_324/a_8_24# OR2X1_LOC_91/A 0.03fF
C25488 AND2X1_LOC_824/B OR2X1_LOC_39/A 0.14fF
C25489 OR2X1_LOC_158/A OR2X1_LOC_417/A 0.20fF
C25490 AND2X1_LOC_719/Y AND2X1_LOC_845/Y 0.50fF
C25491 AND2X1_LOC_807/Y OR2X1_LOC_406/a_8_216# 0.14fF
C25492 AND2X1_LOC_540/a_8_24# OR2X1_LOC_485/A 0.01fF
C25493 OR2X1_LOC_686/a_8_216# AND2X1_LOC_425/Y 0.01fF
C25494 OR2X1_LOC_648/B OR2X1_LOC_655/B 0.15fF
C25495 OR2X1_LOC_329/B AND2X1_LOC_523/Y 0.07fF
C25496 OR2X1_LOC_154/A AND2X1_LOC_43/B 3.15fF
C25497 AND2X1_LOC_56/B OR2X1_LOC_739/A 0.04fF
C25498 AND2X1_LOC_564/A AND2X1_LOC_781/Y 0.01fF
C25499 OR2X1_LOC_85/A OR2X1_LOC_39/A 0.07fF
C25500 AND2X1_LOC_81/B OR2X1_LOC_375/A 0.11fF
C25501 OR2X1_LOC_51/Y OR2X1_LOC_22/Y 0.14fF
C25502 OR2X1_LOC_792/Y OR2X1_LOC_807/a_8_216# 0.02fF
C25503 AND2X1_LOC_49/a_8_24# OR2X1_LOC_375/A 0.01fF
C25504 OR2X1_LOC_26/Y OR2X1_LOC_619/Y 0.13fF
C25505 INPUT_0 OR2X1_LOC_275/a_36_216# 0.03fF
C25506 AND2X1_LOC_95/Y OR2X1_LOC_346/B 0.15fF
C25507 OR2X1_LOC_650/Y OR2X1_LOC_520/a_8_216# 0.01fF
C25508 OR2X1_LOC_538/a_8_216# OR2X1_LOC_193/A 0.01fF
C25509 OR2X1_LOC_46/A AND2X1_LOC_92/Y 0.03fF
C25510 AND2X1_LOC_22/Y AND2X1_LOC_72/B 0.02fF
C25511 OR2X1_LOC_43/A OR2X1_LOC_316/Y 0.03fF
C25512 AND2X1_LOC_98/Y OR2X1_LOC_64/Y 0.00fF
C25513 OR2X1_LOC_16/A D_INPUT_1 0.19fF
C25514 AND2X1_LOC_388/a_8_24# AND2X1_LOC_661/A 0.01fF
C25515 OR2X1_LOC_291/a_8_216# OR2X1_LOC_74/A 0.01fF
C25516 AND2X1_LOC_529/a_8_24# OR2X1_LOC_19/B 0.01fF
C25517 OR2X1_LOC_756/B AND2X1_LOC_816/a_8_24# 0.01fF
C25518 OR2X1_LOC_471/Y OR2X1_LOC_742/a_8_216# 0.06fF
C25519 OR2X1_LOC_433/a_8_216# AND2X1_LOC_319/A 0.05fF
C25520 OR2X1_LOC_89/A OR2X1_LOC_619/Y 0.03fF
C25521 OR2X1_LOC_61/Y OR2X1_LOC_201/Y 0.13fF
C25522 AND2X1_LOC_36/Y OR2X1_LOC_269/A 0.01fF
C25523 AND2X1_LOC_56/B AND2X1_LOC_298/a_8_24# 0.11fF
C25524 AND2X1_LOC_337/a_8_24# AND2X1_LOC_863/Y 0.01fF
C25525 OR2X1_LOC_103/Y OR2X1_LOC_64/Y 0.01fF
C25526 OR2X1_LOC_161/B OR2X1_LOC_544/a_8_216# 0.04fF
C25527 AND2X1_LOC_48/A AND2X1_LOC_693/a_8_24# 0.01fF
C25528 OR2X1_LOC_88/A OR2X1_LOC_26/Y 0.01fF
C25529 AND2X1_LOC_20/a_8_24# D_INPUT_0 0.02fF
C25530 OR2X1_LOC_431/Y AND2X1_LOC_654/B 0.25fF
C25531 OR2X1_LOC_22/Y OR2X1_LOC_58/a_8_216# 0.01fF
C25532 AND2X1_LOC_56/B OR2X1_LOC_269/B 0.28fF
C25533 OR2X1_LOC_483/a_36_216# OR2X1_LOC_631/B 0.01fF
C25534 OR2X1_LOC_756/B OR2X1_LOC_859/A 0.11fF
C25535 OR2X1_LOC_87/A OR2X1_LOC_155/A 0.15fF
C25536 AND2X1_LOC_36/Y AND2X1_LOC_41/Y 0.03fF
C25537 OR2X1_LOC_634/A D_INPUT_0 0.00fF
C25538 AND2X1_LOC_365/A AND2X1_LOC_390/B 0.02fF
C25539 AND2X1_LOC_40/Y OR2X1_LOC_443/Y 0.00fF
C25540 OR2X1_LOC_101/a_8_216# OR2X1_LOC_121/B 0.01fF
C25541 AND2X1_LOC_866/A OR2X1_LOC_56/A 4.45fF
C25542 AND2X1_LOC_303/B OR2X1_LOC_7/A -0.02fF
C25543 OR2X1_LOC_103/a_8_216# OR2X1_LOC_64/Y 0.01fF
C25544 AND2X1_LOC_710/Y AND2X1_LOC_866/A 0.02fF
C25545 OR2X1_LOC_574/A OR2X1_LOC_203/Y 0.36fF
C25546 OR2X1_LOC_538/a_8_216# D_INPUT_0 0.02fF
C25547 AND2X1_LOC_21/Y AND2X1_LOC_26/a_8_24# 0.03fF
C25548 AND2X1_LOC_624/A AND2X1_LOC_624/a_8_24# 0.10fF
C25549 OR2X1_LOC_858/A OR2X1_LOC_276/B 0.02fF
C25550 AND2X1_LOC_789/Y AND2X1_LOC_793/a_8_24# 0.05fF
C25551 OR2X1_LOC_423/a_8_216# OR2X1_LOC_52/B 0.03fF
C25552 AND2X1_LOC_557/Y AND2X1_LOC_557/a_8_24# 0.01fF
C25553 AND2X1_LOC_532/a_8_24# AND2X1_LOC_727/A 0.01fF
C25554 OR2X1_LOC_778/Y OR2X1_LOC_784/a_8_216# 0.01fF
C25555 OR2X1_LOC_451/a_8_216# OR2X1_LOC_451/B 0.08fF
C25556 OR2X1_LOC_605/A OR2X1_LOC_87/A 0.12fF
C25557 OR2X1_LOC_70/Y AND2X1_LOC_319/A 0.17fF
C25558 OR2X1_LOC_185/A AND2X1_LOC_518/a_8_24# 0.04fF
C25559 OR2X1_LOC_585/A AND2X1_LOC_294/a_8_24# 0.11fF
C25560 OR2X1_LOC_517/A OR2X1_LOC_256/A 5.09fF
C25561 AND2X1_LOC_656/Y AND2X1_LOC_141/A 0.09fF
C25562 AND2X1_LOC_720/Y OR2X1_LOC_417/A 0.02fF
C25563 AND2X1_LOC_839/A AND2X1_LOC_839/a_8_24# 0.10fF
C25564 AND2X1_LOC_390/B OR2X1_LOC_43/A 0.07fF
C25565 OR2X1_LOC_112/B OR2X1_LOC_78/B 0.23fF
C25566 OR2X1_LOC_121/B OR2X1_LOC_340/Y 0.01fF
C25567 OR2X1_LOC_185/A AND2X1_LOC_48/A 0.02fF
C25568 AND2X1_LOC_687/B AND2X1_LOC_452/Y 0.01fF
C25569 OR2X1_LOC_3/B OR2X1_LOC_12/a_8_216# 0.01fF
C25570 OR2X1_LOC_121/B OR2X1_LOC_130/A 0.03fF
C25571 OR2X1_LOC_780/B AND2X1_LOC_424/a_36_24# 0.01fF
C25572 OR2X1_LOC_139/a_8_216# AND2X1_LOC_42/B 0.01fF
C25573 AND2X1_LOC_721/A OR2X1_LOC_59/Y 0.00fF
C25574 OR2X1_LOC_196/B OR2X1_LOC_375/A 0.04fF
C25575 AND2X1_LOC_43/a_8_24# OR2X1_LOC_195/A 0.09fF
C25576 AND2X1_LOC_831/Y AND2X1_LOC_649/B 0.00fF
C25577 OR2X1_LOC_616/Y AND2X1_LOC_621/a_8_24# 0.10fF
C25578 AND2X1_LOC_734/Y OR2X1_LOC_47/Y 0.03fF
C25579 OR2X1_LOC_91/A OR2X1_LOC_597/Y 0.09fF
C25580 AND2X1_LOC_841/B OR2X1_LOC_31/Y 0.01fF
C25581 OR2X1_LOC_185/A AND2X1_LOC_69/a_36_24# 0.00fF
C25582 OR2X1_LOC_201/a_8_216# OR2X1_LOC_61/Y 0.05fF
C25583 OR2X1_LOC_246/Y OR2X1_LOC_246/A 0.02fF
C25584 AND2X1_LOC_692/a_8_24# OR2X1_LOC_375/A 0.01fF
C25585 AND2X1_LOC_580/A OR2X1_LOC_628/Y 0.07fF
C25586 AND2X1_LOC_285/Y OR2X1_LOC_753/Y 0.02fF
C25587 OR2X1_LOC_109/Y AND2X1_LOC_831/Y 0.02fF
C25588 OR2X1_LOC_337/A OR2X1_LOC_303/B 0.01fF
C25589 OR2X1_LOC_54/Y AND2X1_LOC_818/a_8_24# 0.10fF
C25590 AND2X1_LOC_864/a_8_24# OR2X1_LOC_619/Y 0.06fF
C25591 OR2X1_LOC_709/A AND2X1_LOC_419/a_36_24# -0.01fF
C25592 OR2X1_LOC_782/B OR2X1_LOC_782/a_8_216# 0.47fF
C25593 AND2X1_LOC_773/Y OR2X1_LOC_300/Y 0.02fF
C25594 AND2X1_LOC_465/A OR2X1_LOC_183/a_36_216# 0.00fF
C25595 OR2X1_LOC_392/A D_INPUT_1 0.00fF
C25596 OR2X1_LOC_87/A OR2X1_LOC_782/a_8_216# 0.01fF
C25597 AND2X1_LOC_365/A AND2X1_LOC_863/Y 0.25fF
C25598 AND2X1_LOC_303/A D_INPUT_0 0.09fF
C25599 AND2X1_LOC_344/a_36_24# OR2X1_LOC_47/Y 0.00fF
C25600 OR2X1_LOC_517/A OR2X1_LOC_67/Y 0.03fF
C25601 OR2X1_LOC_7/Y OR2X1_LOC_44/Y 0.43fF
C25602 OR2X1_LOC_644/B OR2X1_LOC_644/a_8_216# 0.07fF
C25603 OR2X1_LOC_26/Y OR2X1_LOC_22/A 0.04fF
C25604 AND2X1_LOC_64/Y OR2X1_LOC_502/a_8_216# 0.01fF
C25605 OR2X1_LOC_232/a_8_216# OR2X1_LOC_54/Y 0.03fF
C25606 OR2X1_LOC_624/A OR2X1_LOC_506/B 0.05fF
C25607 OR2X1_LOC_841/a_8_216# OR2X1_LOC_804/A 0.03fF
C25608 AND2X1_LOC_22/Y AND2X1_LOC_36/Y 2.94fF
C25609 AND2X1_LOC_642/a_36_24# AND2X1_LOC_476/A 0.01fF
C25610 AND2X1_LOC_92/Y OR2X1_LOC_641/B 0.01fF
C25611 OR2X1_LOC_109/a_8_216# OR2X1_LOC_47/Y 0.01fF
C25612 OR2X1_LOC_87/A OR2X1_LOC_228/a_8_216# 0.01fF
C25613 OR2X1_LOC_406/a_8_216# OR2X1_LOC_95/Y 0.02fF
C25614 OR2X1_LOC_59/Y OR2X1_LOC_331/Y 0.02fF
C25615 OR2X1_LOC_244/Y OR2X1_LOC_68/B 0.03fF
C25616 OR2X1_LOC_91/Y AND2X1_LOC_227/Y 0.03fF
C25617 OR2X1_LOC_66/Y OR2X1_LOC_721/Y 0.05fF
C25618 OR2X1_LOC_638/B AND2X1_LOC_31/Y 0.03fF
C25619 OR2X1_LOC_774/Y OR2X1_LOC_773/a_8_216# 0.01fF
C25620 AND2X1_LOC_401/Y OR2X1_LOC_598/A 0.01fF
C25621 AND2X1_LOC_684/a_8_24# AND2X1_LOC_43/B 0.06fF
C25622 AND2X1_LOC_839/A AND2X1_LOC_839/B 0.10fF
C25623 AND2X1_LOC_18/Y OR2X1_LOC_366/Y 0.00fF
C25624 OR2X1_LOC_31/Y OR2X1_LOC_22/a_8_216# 0.01fF
C25625 OR2X1_LOC_780/B OR2X1_LOC_449/B 0.09fF
C25626 OR2X1_LOC_507/B OR2X1_LOC_205/Y 0.03fF
C25627 AND2X1_LOC_22/Y OR2X1_LOC_333/a_8_216# 0.02fF
C25628 OR2X1_LOC_485/A D_INPUT_0 0.17fF
C25629 OR2X1_LOC_680/Y AND2X1_LOC_678/a_8_24# 0.00fF
C25630 AND2X1_LOC_51/A AND2X1_LOC_47/Y 0.04fF
C25631 AND2X1_LOC_512/Y OR2X1_LOC_534/a_8_216# 0.03fF
C25632 OR2X1_LOC_85/A OR2X1_LOC_826/Y 0.05fF
C25633 OR2X1_LOC_840/A OR2X1_LOC_228/Y 0.10fF
C25634 AND2X1_LOC_621/Y AND2X1_LOC_795/Y 0.65fF
C25635 OR2X1_LOC_429/a_8_216# OR2X1_LOC_17/Y 0.05fF
C25636 AND2X1_LOC_111/a_8_24# D_INPUT_0 0.02fF
C25637 AND2X1_LOC_624/A AND2X1_LOC_624/B 0.45fF
C25638 AND2X1_LOC_432/a_36_24# OR2X1_LOC_390/B 0.00fF
C25639 OR2X1_LOC_109/Y AND2X1_LOC_405/a_8_24# 0.01fF
C25640 OR2X1_LOC_621/A AND2X1_LOC_36/Y 0.01fF
C25641 OR2X1_LOC_205/a_8_216# OR2X1_LOC_786/Y 0.01fF
C25642 D_INPUT_3 OR2X1_LOC_106/A 0.06fF
C25643 OR2X1_LOC_291/Y OR2X1_LOC_46/A 0.17fF
C25644 OR2X1_LOC_375/A OR2X1_LOC_66/Y 0.20fF
C25645 OR2X1_LOC_311/Y OR2X1_LOC_46/A 0.02fF
C25646 OR2X1_LOC_185/A OR2X1_LOC_398/a_8_216# 0.02fF
C25647 OR2X1_LOC_805/A OR2X1_LOC_717/a_8_216# 0.06fF
C25648 OR2X1_LOC_70/Y OR2X1_LOC_604/a_8_216# 0.01fF
C25649 OR2X1_LOC_70/Y AND2X1_LOC_170/B 0.01fF
C25650 AND2X1_LOC_64/Y OR2X1_LOC_691/a_8_216# 0.01fF
C25651 AND2X1_LOC_544/Y AND2X1_LOC_469/a_8_24# 0.03fF
C25652 OR2X1_LOC_19/B OR2X1_LOC_532/B 0.14fF
C25653 OR2X1_LOC_174/a_36_216# OR2X1_LOC_390/A 0.01fF
C25654 AND2X1_LOC_634/Y AND2X1_LOC_640/a_8_24# 0.00fF
C25655 OR2X1_LOC_121/B OR2X1_LOC_780/B 0.17fF
C25656 OR2X1_LOC_78/A OR2X1_LOC_579/A 0.26fF
C25657 OR2X1_LOC_357/a_8_216# OR2X1_LOC_357/B 0.03fF
C25658 OR2X1_LOC_417/Y OR2X1_LOC_604/a_36_216# 0.00fF
C25659 AND2X1_LOC_514/Y AND2X1_LOC_170/B 0.02fF
C25660 OR2X1_LOC_78/A OR2X1_LOC_844/B 0.42fF
C25661 AND2X1_LOC_43/B OR2X1_LOC_198/A 0.00fF
C25662 OR2X1_LOC_222/A OR2X1_LOC_228/Y 0.01fF
C25663 OR2X1_LOC_106/Y AND2X1_LOC_243/Y 0.05fF
C25664 AND2X1_LOC_521/a_36_24# AND2X1_LOC_22/Y 0.00fF
C25665 OR2X1_LOC_91/a_36_216# AND2X1_LOC_222/Y 0.00fF
C25666 OR2X1_LOC_18/Y OR2X1_LOC_384/Y 0.04fF
C25667 OR2X1_LOC_476/B OR2X1_LOC_223/A 0.02fF
C25668 OR2X1_LOC_121/B AND2X1_LOC_88/Y 0.03fF
C25669 AND2X1_LOC_861/B OR2X1_LOC_504/a_8_216# 0.47fF
C25670 D_INPUT_3 OR2X1_LOC_46/A 0.08fF
C25671 AND2X1_LOC_339/B OR2X1_LOC_12/Y 0.03fF
C25672 OR2X1_LOC_78/A OR2X1_LOC_390/B 0.08fF
C25673 OR2X1_LOC_482/Y AND2X1_LOC_242/a_36_24# 0.01fF
C25674 OR2X1_LOC_539/Y OR2X1_LOC_446/B 0.01fF
C25675 AND2X1_LOC_12/Y OR2X1_LOC_558/a_8_216# 0.00fF
C25676 OR2X1_LOC_479/Y OR2X1_LOC_318/B 0.00fF
C25677 AND2X1_LOC_687/B AND2X1_LOC_687/a_8_24# 0.01fF
C25678 OR2X1_LOC_494/A AND2X1_LOC_363/Y 0.06fF
C25679 INPUT_1 AND2X1_LOC_660/A 0.07fF
C25680 AND2X1_LOC_725/a_8_24# OR2X1_LOC_428/A 0.01fF
C25681 OR2X1_LOC_438/Y AND2X1_LOC_439/a_8_24# 0.01fF
C25682 VDD OR2X1_LOC_357/B -0.00fF
C25683 OR2X1_LOC_95/Y AND2X1_LOC_675/A 0.02fF
C25684 OR2X1_LOC_212/a_8_216# OR2X1_LOC_212/B 0.18fF
C25685 AND2X1_LOC_675/A AND2X1_LOC_440/a_8_24# 0.00fF
C25686 OR2X1_LOC_506/a_8_216# AND2X1_LOC_41/A 0.01fF
C25687 OR2X1_LOC_36/Y OR2X1_LOC_589/Y 0.01fF
C25688 AND2X1_LOC_22/Y AND2X1_LOC_95/a_36_24# 0.00fF
C25689 OR2X1_LOC_714/Y OR2X1_LOC_308/Y 0.00fF
C25690 OR2X1_LOC_45/B AND2X1_LOC_454/a_8_24# 0.02fF
C25691 OR2X1_LOC_66/A OR2X1_LOC_342/A 0.03fF
C25692 AND2X1_LOC_11/Y INPUT_6 0.84fF
C25693 AND2X1_LOC_227/Y D_INPUT_3 0.00fF
C25694 OR2X1_LOC_70/Y OR2X1_LOC_331/Y 0.12fF
C25695 VDD AND2X1_LOC_774/A 0.75fF
C25696 OR2X1_LOC_121/B OR2X1_LOC_365/B 0.03fF
C25697 AND2X1_LOC_40/Y AND2X1_LOC_763/B 0.00fF
C25698 AND2X1_LOC_450/Y AND2X1_LOC_452/a_8_24# 0.19fF
C25699 AND2X1_LOC_141/A AND2X1_LOC_772/Y 0.01fF
C25700 OR2X1_LOC_426/B OR2X1_LOC_16/A 6.52fF
C25701 OR2X1_LOC_492/Y OR2X1_LOC_108/Y 0.13fF
C25702 OR2X1_LOC_45/B AND2X1_LOC_663/A 0.03fF
C25703 AND2X1_LOC_50/Y AND2X1_LOC_64/Y 0.00fF
C25704 AND2X1_LOC_70/Y OR2X1_LOC_355/a_8_216# 0.04fF
C25705 AND2X1_LOC_765/a_8_24# OR2X1_LOC_78/B 0.03fF
C25706 OR2X1_LOC_472/a_8_216# OR2X1_LOC_68/B 0.01fF
C25707 OR2X1_LOC_108/a_8_216# OR2X1_LOC_108/Y 0.05fF
C25708 OR2X1_LOC_778/Y OR2X1_LOC_777/B 0.07fF
C25709 OR2X1_LOC_292/Y OR2X1_LOC_428/A 0.01fF
C25710 OR2X1_LOC_92/Y AND2X1_LOC_473/Y 0.23fF
C25711 OR2X1_LOC_207/B AND2X1_LOC_693/a_8_24# 0.01fF
C25712 AND2X1_LOC_706/a_8_24# OR2X1_LOC_744/A 0.01fF
C25713 OR2X1_LOC_506/Y OR2X1_LOC_244/B 0.10fF
C25714 OR2X1_LOC_369/Y AND2X1_LOC_182/A 0.00fF
C25715 AND2X1_LOC_657/Y AND2X1_LOC_477/Y 0.10fF
C25716 AND2X1_LOC_41/A AND2X1_LOC_256/a_8_24# 0.06fF
C25717 OR2X1_LOC_635/A AND2X1_LOC_22/Y 0.01fF
C25718 OR2X1_LOC_589/A OR2X1_LOC_744/A 0.40fF
C25719 OR2X1_LOC_528/Y AND2X1_LOC_570/Y 0.02fF
C25720 AND2X1_LOC_595/a_8_24# OR2X1_LOC_244/Y 0.01fF
C25721 OR2X1_LOC_860/Y OR2X1_LOC_474/B 0.89fF
C25722 OR2X1_LOC_92/Y OR2X1_LOC_816/A 0.04fF
C25723 AND2X1_LOC_477/Y AND2X1_LOC_469/B 0.17fF
C25724 AND2X1_LOC_738/B OR2X1_LOC_40/Y 0.07fF
C25725 OR2X1_LOC_97/A OR2X1_LOC_785/B 0.03fF
C25726 AND2X1_LOC_3/Y OR2X1_LOC_217/A 0.00fF
C25727 OR2X1_LOC_159/a_8_216# OR2X1_LOC_56/A 0.05fF
C25728 OR2X1_LOC_485/Y OR2X1_LOC_51/Y 0.02fF
C25729 AND2X1_LOC_803/B VDD 0.18fF
C25730 OR2X1_LOC_40/Y OR2X1_LOC_56/A 0.45fF
C25731 OR2X1_LOC_538/a_36_216# OR2X1_LOC_161/B 0.00fF
C25732 OR2X1_LOC_602/A OR2X1_LOC_390/B 0.14fF
C25733 OR2X1_LOC_186/Y OR2X1_LOC_354/A 0.04fF
C25734 OR2X1_LOC_160/B OR2X1_LOC_35/Y 0.10fF
C25735 OR2X1_LOC_447/A AND2X1_LOC_7/B 0.00fF
C25736 AND2X1_LOC_586/a_8_24# AND2X1_LOC_22/Y 0.01fF
C25737 OR2X1_LOC_427/A OR2X1_LOC_753/a_36_216# 0.00fF
C25738 OR2X1_LOC_426/B AND2X1_LOC_121/a_8_24# 0.02fF
C25739 AND2X1_LOC_297/a_8_24# AND2X1_LOC_44/Y 0.01fF
C25740 VDD OR2X1_LOC_755/a_8_216# 0.00fF
C25741 OR2X1_LOC_858/A AND2X1_LOC_70/Y 0.16fF
C25742 AND2X1_LOC_212/A OR2X1_LOC_92/Y 0.05fF
C25743 AND2X1_LOC_318/Y AND2X1_LOC_222/Y 0.02fF
C25744 AND2X1_LOC_228/Y AND2X1_LOC_231/a_8_24# 0.01fF
C25745 OR2X1_LOC_114/B OR2X1_LOC_735/a_8_216# 0.01fF
C25746 AND2X1_LOC_59/Y OR2X1_LOC_139/A 0.03fF
C25747 OR2X1_LOC_155/A OR2X1_LOC_390/B 0.07fF
C25748 OR2X1_LOC_105/Y OR2X1_LOC_362/A 0.02fF
C25749 OR2X1_LOC_45/B AND2X1_LOC_449/Y 0.01fF
C25750 AND2X1_LOC_735/Y AND2X1_LOC_500/Y 0.16fF
C25751 OR2X1_LOC_756/B OR2X1_LOC_66/A 0.75fF
C25752 OR2X1_LOC_842/a_8_216# VDD 0.00fF
C25753 OR2X1_LOC_196/B OR2X1_LOC_515/Y 0.33fF
C25754 AND2X1_LOC_12/Y OR2X1_LOC_138/A 0.04fF
C25755 OR2X1_LOC_778/Y OR2X1_LOC_831/B 0.07fF
C25756 OR2X1_LOC_698/a_8_216# OR2X1_LOC_56/A 0.05fF
C25757 OR2X1_LOC_739/B OR2X1_LOC_740/B 0.07fF
C25758 OR2X1_LOC_271/Y AND2X1_LOC_473/Y 0.29fF
C25759 OR2X1_LOC_331/A AND2X1_LOC_512/Y 0.04fF
C25760 OR2X1_LOC_158/A AND2X1_LOC_161/a_8_24# 0.01fF
C25761 OR2X1_LOC_255/a_36_216# OR2X1_LOC_437/A 0.01fF
C25762 OR2X1_LOC_833/Y OR2X1_LOC_375/A 0.16fF
C25763 OR2X1_LOC_691/Y OR2X1_LOC_793/A 0.00fF
C25764 AND2X1_LOC_702/Y OR2X1_LOC_428/A 0.05fF
C25765 AND2X1_LOC_177/a_8_24# OR2X1_LOC_78/A 0.02fF
C25766 AND2X1_LOC_539/Y OR2X1_LOC_485/A 0.04fF
C25767 OR2X1_LOC_441/Y AND2X1_LOC_659/a_8_24# 0.01fF
C25768 OR2X1_LOC_136/Y AND2X1_LOC_211/B 0.13fF
C25769 OR2X1_LOC_185/A OR2X1_LOC_542/a_8_216# 0.01fF
C25770 OR2X1_LOC_621/a_8_216# OR2X1_LOC_847/A 0.01fF
C25771 OR2X1_LOC_699/a_8_216# OR2X1_LOC_12/Y 0.01fF
C25772 OR2X1_LOC_214/a_8_216# AND2X1_LOC_44/Y 0.01fF
C25773 OR2X1_LOC_624/a_36_216# OR2X1_LOC_624/Y 0.01fF
C25774 OR2X1_LOC_115/a_8_216# OR2X1_LOC_140/A 0.47fF
C25775 OR2X1_LOC_319/a_36_216# AND2X1_LOC_110/Y 0.00fF
C25776 OR2X1_LOC_134/Y OR2X1_LOC_272/Y 0.04fF
C25777 AND2X1_LOC_81/B OR2X1_LOC_549/A 0.03fF
C25778 OR2X1_LOC_494/Y OR2X1_LOC_427/A 0.03fF
C25779 AND2X1_LOC_49/a_8_24# OR2X1_LOC_549/A 0.01fF
C25780 AND2X1_LOC_363/Y OR2X1_LOC_427/A 0.06fF
C25781 OR2X1_LOC_744/A AND2X1_LOC_654/B 0.03fF
C25782 AND2X1_LOC_713/Y AND2X1_LOC_448/Y 0.01fF
C25783 OR2X1_LOC_86/A OR2X1_LOC_88/Y 0.00fF
C25784 OR2X1_LOC_624/A AND2X1_LOC_18/Y 0.19fF
C25785 AND2X1_LOC_64/Y OR2X1_LOC_473/Y 0.45fF
C25786 AND2X1_LOC_367/A OR2X1_LOC_256/Y 0.03fF
C25787 AND2X1_LOC_448/Y AND2X1_LOC_448/a_36_24# 0.00fF
C25788 OR2X1_LOC_653/Y AND2X1_LOC_19/Y 0.00fF
C25789 OR2X1_LOC_40/Y AND2X1_LOC_87/a_8_24# 0.02fF
C25790 OR2X1_LOC_467/A AND2X1_LOC_426/a_8_24# 0.01fF
C25791 VDD OR2X1_LOC_137/B 0.03fF
C25792 AND2X1_LOC_737/a_8_24# OR2X1_LOC_441/Y 0.01fF
C25793 AND2X1_LOC_398/a_8_24# OR2X1_LOC_744/A 0.23fF
C25794 AND2X1_LOC_810/Y OR2X1_LOC_142/Y 0.37fF
C25795 AND2X1_LOC_736/Y AND2X1_LOC_736/a_36_24# 0.00fF
C25796 AND2X1_LOC_558/a_8_24# AND2X1_LOC_573/A 0.01fF
C25797 OR2X1_LOC_630/a_8_216# OR2X1_LOC_630/Y 0.01fF
C25798 OR2X1_LOC_91/A OR2X1_LOC_48/B 0.21fF
C25799 AND2X1_LOC_776/a_36_24# OR2X1_LOC_18/Y 0.00fF
C25800 OR2X1_LOC_51/Y OR2X1_LOC_39/A 0.22fF
C25801 OR2X1_LOC_743/A OR2X1_LOC_16/A 0.08fF
C25802 OR2X1_LOC_739/A AND2X1_LOC_92/Y 0.03fF
C25803 OR2X1_LOC_46/A OR2X1_LOC_171/Y 0.00fF
C25804 OR2X1_LOC_411/Y OR2X1_LOC_413/Y 0.21fF
C25805 OR2X1_LOC_170/Y OR2X1_LOC_568/A 0.22fF
C25806 AND2X1_LOC_858/B OR2X1_LOC_18/Y 1.11fF
C25807 AND2X1_LOC_580/A AND2X1_LOC_508/B 0.03fF
C25808 OR2X1_LOC_6/A OR2X1_LOC_14/a_8_216# 0.41fF
C25809 OR2X1_LOC_605/B AND2X1_LOC_604/a_36_24# 0.00fF
C25810 OR2X1_LOC_91/A OR2X1_LOC_18/Y 0.12fF
C25811 AND2X1_LOC_721/Y OR2X1_LOC_64/Y 0.05fF
C25812 VDD OR2X1_LOC_613/Y 0.31fF
C25813 AND2X1_LOC_31/Y OR2X1_LOC_779/B 0.03fF
C25814 OR2X1_LOC_170/Y OR2X1_LOC_578/B 0.01fF
C25815 AND2X1_LOC_94/a_36_24# INPUT_0 0.01fF
C25816 AND2X1_LOC_365/A OR2X1_LOC_744/A 0.43fF
C25817 OR2X1_LOC_87/A OR2X1_LOC_797/a_36_216# 0.00fF
C25818 OR2X1_LOC_602/a_36_216# OR2X1_LOC_161/B 0.00fF
C25819 OR2X1_LOC_45/B AND2X1_LOC_856/a_8_24# 0.03fF
C25820 OR2X1_LOC_448/B AND2X1_LOC_422/a_8_24# 0.21fF
C25821 OR2X1_LOC_76/Y OR2X1_LOC_66/A 0.03fF
C25822 OR2X1_LOC_814/A OR2X1_LOC_174/a_8_216# 0.03fF
C25823 AND2X1_LOC_96/a_8_24# AND2X1_LOC_43/B 0.19fF
C25824 OR2X1_LOC_744/A AND2X1_LOC_379/a_8_24# 0.01fF
C25825 AND2X1_LOC_486/Y AND2X1_LOC_833/a_8_24# 0.06fF
C25826 AND2X1_LOC_508/A AND2X1_LOC_573/A 0.00fF
C25827 VDD AND2X1_LOC_252/a_8_24# 0.00fF
C25828 OR2X1_LOC_74/A AND2X1_LOC_443/a_36_24# 0.01fF
C25829 OR2X1_LOC_468/A OR2X1_LOC_449/B 0.03fF
C25830 AND2X1_LOC_84/a_8_24# OR2X1_LOC_600/A 0.05fF
C25831 AND2X1_LOC_363/Y AND2X1_LOC_363/A 0.10fF
C25832 AND2X1_LOC_191/Y AND2X1_LOC_479/a_36_24# 0.01fF
C25833 AND2X1_LOC_468/B OR2X1_LOC_594/a_36_216# 0.01fF
C25834 AND2X1_LOC_571/A OR2X1_LOC_95/Y 0.03fF
C25835 OR2X1_LOC_26/Y AND2X1_LOC_286/a_8_24# 0.01fF
C25836 OR2X1_LOC_58/a_8_216# OR2X1_LOC_39/A 0.01fF
C25837 OR2X1_LOC_347/B OR2X1_LOC_736/A 0.09fF
C25838 OR2X1_LOC_25/Y OR2X1_LOC_44/Y 0.03fF
C25839 OR2X1_LOC_555/A AND2X1_LOC_18/Y 0.18fF
C25840 OR2X1_LOC_820/A OR2X1_LOC_96/B 0.03fF
C25841 OR2X1_LOC_308/A AND2X1_LOC_47/Y 0.01fF
C25842 OR2X1_LOC_40/Y AND2X1_LOC_641/Y 0.39fF
C25843 AND2X1_LOC_543/Y OR2X1_LOC_31/Y 0.01fF
C25844 OR2X1_LOC_744/A OR2X1_LOC_43/A 0.10fF
C25845 AND2X1_LOC_92/Y OR2X1_LOC_269/B 0.13fF
C25846 OR2X1_LOC_40/Y OR2X1_LOC_291/A 0.06fF
C25847 AND2X1_LOC_574/a_8_24# AND2X1_LOC_576/Y 0.03fF
C25848 AND2X1_LOC_59/Y OR2X1_LOC_850/B 0.00fF
C25849 AND2X1_LOC_211/B OR2X1_LOC_51/Y 0.03fF
C25850 OR2X1_LOC_147/B AND2X1_LOC_315/a_8_24# 0.03fF
C25851 OR2X1_LOC_6/B AND2X1_LOC_117/a_8_24# 0.03fF
C25852 OR2X1_LOC_85/A AND2X1_LOC_240/a_8_24# 0.01fF
C25853 OR2X1_LOC_160/A AND2X1_LOC_331/a_8_24# 0.02fF
C25854 OR2X1_LOC_91/Y AND2X1_LOC_722/A 0.01fF
C25855 OR2X1_LOC_70/Y AND2X1_LOC_479/a_36_24# 0.00fF
C25856 AND2X1_LOC_843/Y AND2X1_LOC_850/Y 0.01fF
C25857 AND2X1_LOC_509/a_8_24# OR2X1_LOC_7/A 0.01fF
C25858 OR2X1_LOC_482/Y OR2X1_LOC_64/Y 0.83fF
C25859 OR2X1_LOC_7/A OR2X1_LOC_56/A 0.53fF
C25860 AND2X1_LOC_227/Y OR2X1_LOC_184/a_36_216# 0.00fF
C25861 AND2X1_LOC_721/Y OR2X1_LOC_417/A 0.06fF
C25862 OR2X1_LOC_864/A OR2X1_LOC_235/B 0.03fF
C25863 AND2X1_LOC_752/a_36_24# AND2X1_LOC_43/B 0.00fF
C25864 OR2X1_LOC_429/Y OR2X1_LOC_51/Y 0.03fF
C25865 OR2X1_LOC_707/B OR2X1_LOC_161/B 0.06fF
C25866 OR2X1_LOC_574/A OR2X1_LOC_78/B 0.03fF
C25867 OR2X1_LOC_426/B OR2X1_LOC_273/a_8_216# 0.01fF
C25868 AND2X1_LOC_594/a_8_24# OR2X1_LOC_814/A 0.02fF
C25869 D_INPUT_0 OR2X1_LOC_633/A 0.01fF
C25870 OR2X1_LOC_11/Y OR2X1_LOC_586/Y 0.15fF
C25871 AND2X1_LOC_231/Y OR2X1_LOC_31/Y 0.00fF
C25872 AND2X1_LOC_624/A AND2X1_LOC_811/B 0.15fF
C25873 OR2X1_LOC_18/Y AND2X1_LOC_573/A 0.14fF
C25874 AND2X1_LOC_139/B AND2X1_LOC_649/B 0.46fF
C25875 OR2X1_LOC_320/Y OR2X1_LOC_56/A 0.01fF
C25876 AND2X1_LOC_95/Y OR2X1_LOC_128/B 0.04fF
C25877 AND2X1_LOC_811/a_8_24# OR2X1_LOC_427/A 0.02fF
C25878 OR2X1_LOC_58/Y OR2X1_LOC_60/a_36_216# 0.00fF
C25879 OR2X1_LOC_485/A AND2X1_LOC_471/Y 0.07fF
C25880 AND2X1_LOC_24/a_8_24# OR2X1_LOC_33/B 0.01fF
C25881 OR2X1_LOC_495/Y AND2X1_LOC_840/B 0.19fF
C25882 OR2X1_LOC_139/a_8_216# OR2X1_LOC_663/A 0.04fF
C25883 OR2X1_LOC_405/A AND2X1_LOC_272/a_8_24# -0.01fF
C25884 OR2X1_LOC_624/B AND2X1_LOC_103/a_8_24# 0.02fF
C25885 OR2X1_LOC_653/Y OR2X1_LOC_653/A 0.01fF
C25886 OR2X1_LOC_633/Y OR2X1_LOC_640/a_8_216# 0.04fF
C25887 OR2X1_LOC_792/B OR2X1_LOC_792/a_8_216# 0.01fF
C25888 OR2X1_LOC_185/A OR2X1_LOC_350/a_8_216# 0.01fF
C25889 OR2X1_LOC_440/A OR2X1_LOC_161/B 0.07fF
C25890 OR2X1_LOC_524/Y AND2X1_LOC_728/a_8_24# 0.13fF
C25891 OR2X1_LOC_377/A AND2X1_LOC_824/B 3.84fF
C25892 AND2X1_LOC_7/Y OR2X1_LOC_596/A 0.11fF
C25893 OR2X1_LOC_31/Y AND2X1_LOC_770/a_8_24# 0.01fF
C25894 AND2X1_LOC_199/a_8_24# OR2X1_LOC_13/Y 0.01fF
C25895 AND2X1_LOC_347/Y OR2X1_LOC_297/Y 0.06fF
C25896 OR2X1_LOC_148/B OR2X1_LOC_161/A 0.01fF
C25897 AND2X1_LOC_716/Y OR2X1_LOC_312/Y 0.07fF
C25898 AND2X1_LOC_677/a_8_24# OR2X1_LOC_66/A 0.07fF
C25899 OR2X1_LOC_680/A OR2X1_LOC_39/A 7.79fF
C25900 OR2X1_LOC_482/Y OR2X1_LOC_417/A 0.10fF
C25901 OR2X1_LOC_589/A OR2X1_LOC_31/Y 0.02fF
C25902 OR2X1_LOC_160/B AND2X1_LOC_667/a_8_24# 0.03fF
C25903 OR2X1_LOC_816/Y OR2X1_LOC_64/Y 0.12fF
C25904 OR2X1_LOC_667/a_36_216# OR2X1_LOC_278/Y 0.00fF
C25905 OR2X1_LOC_31/Y OR2X1_LOC_322/Y 0.04fF
C25906 AND2X1_LOC_599/a_8_24# OR2X1_LOC_214/B 0.04fF
C25907 OR2X1_LOC_613/Y OR2X1_LOC_616/Y 0.14fF
C25908 OR2X1_LOC_11/Y AND2X1_LOC_459/Y 0.00fF
C25909 AND2X1_LOC_110/Y OR2X1_LOC_532/B 0.03fF
C25910 OR2X1_LOC_158/A OR2X1_LOC_55/a_8_216# 0.02fF
C25911 OR2X1_LOC_401/A OR2X1_LOC_78/Y 0.01fF
C25912 OR2X1_LOC_401/a_8_216# OR2X1_LOC_78/B 0.01fF
C25913 OR2X1_LOC_669/Y OR2X1_LOC_18/Y 0.16fF
C25914 OR2X1_LOC_395/Y OR2X1_LOC_80/A 0.03fF
C25915 OR2X1_LOC_7/A AND2X1_LOC_850/Y 0.46fF
C25916 OR2X1_LOC_168/Y OR2X1_LOC_568/A 0.06fF
C25917 AND2X1_LOC_784/A AND2X1_LOC_655/A 0.10fF
C25918 AND2X1_LOC_110/a_8_24# D_INPUT_0 0.04fF
C25919 AND2X1_LOC_722/A OR2X1_LOC_417/Y 0.14fF
C25920 AND2X1_LOC_22/Y OR2X1_LOC_196/a_8_216# 0.01fF
C25921 OR2X1_LOC_161/B OR2X1_LOC_446/A 0.03fF
C25922 OR2X1_LOC_517/Y AND2X1_LOC_559/a_8_24# 0.23fF
C25923 OR2X1_LOC_185/A AND2X1_LOC_3/Y 0.06fF
C25924 OR2X1_LOC_305/a_8_216# OR2X1_LOC_36/Y 0.01fF
C25925 OR2X1_LOC_455/a_8_216# OR2X1_LOC_553/A -0.03fF
C25926 AND2X1_LOC_31/Y AND2X1_LOC_226/a_8_24# 0.01fF
C25927 OR2X1_LOC_865/B OR2X1_LOC_392/a_8_216# 0.03fF
C25928 D_INPUT_3 INPUT_2 0.09fF
C25929 OR2X1_LOC_154/A AND2X1_LOC_159/a_8_24# 0.16fF
C25930 OR2X1_LOC_617/a_36_216# AND2X1_LOC_805/Y 0.00fF
C25931 OR2X1_LOC_666/Y AND2X1_LOC_624/A 0.03fF
C25932 AND2X1_LOC_576/Y OR2X1_LOC_497/Y 0.94fF
C25933 OR2X1_LOC_669/A OR2X1_LOC_26/Y 0.05fF
C25934 OR2X1_LOC_167/Y AND2X1_LOC_434/Y 0.01fF
C25935 OR2X1_LOC_154/A OR2X1_LOC_810/A 0.18fF
C25936 OR2X1_LOC_437/A OR2X1_LOC_183/Y 0.04fF
C25937 D_INPUT_1 OR2X1_LOC_349/A 0.13fF
C25938 OR2X1_LOC_574/A OR2X1_LOC_375/A 0.05fF
C25939 OR2X1_LOC_446/B OR2X1_LOC_319/Y 0.06fF
C25940 OR2X1_LOC_476/B OR2X1_LOC_502/A 0.65fF
C25941 AND2X1_LOC_70/Y OR2X1_LOC_614/a_8_216# 0.01fF
C25942 OR2X1_LOC_87/A OR2X1_LOC_68/a_8_216# 0.01fF
C25943 AND2X1_LOC_728/Y OR2X1_LOC_680/Y 0.01fF
C25944 OR2X1_LOC_83/a_36_216# OR2X1_LOC_394/Y 0.00fF
C25945 AND2X1_LOC_12/Y OR2X1_LOC_479/Y 0.07fF
C25946 OR2X1_LOC_329/B OR2X1_LOC_111/Y 0.08fF
C25947 AND2X1_LOC_727/A OR2X1_LOC_92/Y 0.03fF
C25948 OR2X1_LOC_66/Y OR2X1_LOC_549/A 0.04fF
C25949 OR2X1_LOC_224/a_8_216# OR2X1_LOC_56/A 0.01fF
C25950 OR2X1_LOC_251/Y OR2X1_LOC_669/a_8_216# 0.01fF
C25951 OR2X1_LOC_377/A AND2X1_LOC_670/a_8_24# 0.02fF
C25952 GATE_811 AND2X1_LOC_657/Y 0.39fF
C25953 OR2X1_LOC_601/Y AND2X1_LOC_645/A 0.01fF
C25954 AND2X1_LOC_191/B GATE_662 0.01fF
C25955 OR2X1_LOC_89/A AND2X1_LOC_818/a_8_24# 0.01fF
C25956 INPUT_1 AND2X1_LOC_642/Y 0.03fF
C25957 OR2X1_LOC_600/A AND2X1_LOC_792/Y 0.19fF
C25958 OR2X1_LOC_31/Y OR2X1_LOC_275/Y 0.28fF
C25959 OR2X1_LOC_231/B OR2X1_LOC_68/B 0.01fF
C25960 AND2X1_LOC_430/a_8_24# OR2X1_LOC_161/A 0.05fF
C25961 AND2X1_LOC_543/a_36_24# OR2X1_LOC_31/Y 0.00fF
C25962 OR2X1_LOC_841/B OR2X1_LOC_479/Y 0.04fF
C25963 OR2X1_LOC_417/Y AND2X1_LOC_454/Y 0.03fF
C25964 OR2X1_LOC_528/Y OR2X1_LOC_406/A 0.00fF
C25965 AND2X1_LOC_516/a_36_24# OR2X1_LOC_155/A 0.01fF
C25966 OR2X1_LOC_613/Y AND2X1_LOC_624/a_8_24# 0.01fF
C25967 OR2X1_LOC_148/B AND2X1_LOC_51/Y 0.13fF
C25968 OR2X1_LOC_709/A AND2X1_LOC_31/Y 0.03fF
C25969 OR2X1_LOC_279/Y OR2X1_LOC_44/Y 0.31fF
C25970 OR2X1_LOC_279/a_36_216# AND2X1_LOC_806/A 0.00fF
C25971 OR2X1_LOC_630/a_36_216# OR2X1_LOC_62/B 0.00fF
C25972 OR2X1_LOC_600/A AND2X1_LOC_259/a_8_24# 0.01fF
C25973 OR2X1_LOC_709/A OR2X1_LOC_715/a_8_216# 0.03fF
C25974 AND2X1_LOC_654/B OR2X1_LOC_31/Y 0.08fF
C25975 OR2X1_LOC_70/Y AND2X1_LOC_361/A 0.08fF
C25976 OR2X1_LOC_235/B OR2X1_LOC_47/Y 0.00fF
C25977 OR2X1_LOC_92/Y OR2X1_LOC_95/Y 0.35fF
C25978 OR2X1_LOC_154/A OR2X1_LOC_857/a_8_216# 0.03fF
C25979 OR2X1_LOC_756/B OR2X1_LOC_84/A -0.00fF
C25980 AND2X1_LOC_91/B OR2X1_LOC_777/B 0.09fF
C25981 OR2X1_LOC_495/Y OR2X1_LOC_31/Y 0.03fF
C25982 AND2X1_LOC_465/a_8_24# AND2X1_LOC_717/B 0.01fF
C25983 OR2X1_LOC_517/A AND2X1_LOC_660/A 0.09fF
C25984 AND2X1_LOC_576/Y AND2X1_LOC_844/a_8_24# 0.01fF
C25985 OR2X1_LOC_402/a_8_216# AND2X1_LOC_3/Y 0.02fF
C25986 OR2X1_LOC_599/A OR2X1_LOC_417/Y 0.03fF
C25987 OR2X1_LOC_351/B OR2X1_LOC_68/B 0.07fF
C25988 OR2X1_LOC_216/A OR2X1_LOC_473/A 0.05fF
C25989 OR2X1_LOC_78/A OR2X1_LOC_493/Y 0.01fF
C25990 AND2X1_LOC_170/Y AND2X1_LOC_514/Y 0.04fF
C25991 OR2X1_LOC_743/A OR2X1_LOC_273/a_8_216# 0.01fF
C25992 OR2X1_LOC_149/B OR2X1_LOC_209/A 0.03fF
C25993 AND2X1_LOC_145/a_8_24# OR2X1_LOC_148/A 0.22fF
C25994 AND2X1_LOC_537/Y OR2X1_LOC_36/Y 0.03fF
C25995 OR2X1_LOC_121/B OR2X1_LOC_449/B 0.09fF
C25996 OR2X1_LOC_16/A OR2X1_LOC_599/a_8_216# 0.01fF
C25997 AND2X1_LOC_334/a_8_24# OR2X1_LOC_26/Y 0.02fF
C25998 AND2X1_LOC_363/a_8_24# OR2X1_LOC_384/Y 0.01fF
C25999 OR2X1_LOC_479/Y OR2X1_LOC_804/B 0.17fF
C26000 OR2X1_LOC_65/a_36_216# OR2X1_LOC_52/B 0.00fF
C26001 OR2X1_LOC_97/A OR2X1_LOC_181/Y 0.06fF
C26002 AND2X1_LOC_683/a_8_24# AND2X1_LOC_51/Y 0.01fF
C26003 OR2X1_LOC_114/B OR2X1_LOC_68/B 0.04fF
C26004 OR2X1_LOC_462/B INPUT_1 0.02fF
C26005 OR2X1_LOC_87/A OR2X1_LOC_814/A 0.82fF
C26006 OR2X1_LOC_494/a_36_216# AND2X1_LOC_721/A 0.00fF
C26007 OR2X1_LOC_664/Y OR2X1_LOC_532/B 0.72fF
C26008 OR2X1_LOC_12/Y OR2X1_LOC_536/a_36_216# 0.03fF
C26009 OR2X1_LOC_83/A OR2X1_LOC_46/A 0.03fF
C26010 OR2X1_LOC_95/Y OR2X1_LOC_65/B 0.06fF
C26011 OR2X1_LOC_12/Y OR2X1_LOC_300/Y 0.07fF
C26012 OR2X1_LOC_458/B OR2X1_LOC_493/Y 0.03fF
C26013 AND2X1_LOC_70/Y AND2X1_LOC_31/Y 3.79fF
C26014 AND2X1_LOC_88/a_8_24# OR2X1_LOC_121/B 0.01fF
C26015 OR2X1_LOC_657/a_36_216# OR2X1_LOC_244/A 0.01fF
C26016 OR2X1_LOC_664/Y AND2X1_LOC_665/a_8_24# 0.00fF
C26017 AND2X1_LOC_69/Y AND2X1_LOC_51/Y 0.01fF
C26018 OR2X1_LOC_754/A OR2X1_LOC_615/a_36_216# 0.00fF
C26019 OR2X1_LOC_596/A OR2X1_LOC_515/a_8_216# 0.01fF
C26020 OR2X1_LOC_309/a_8_216# OR2X1_LOC_437/A -0.01fF
C26021 OR2X1_LOC_59/Y OR2X1_LOC_153/a_36_216# 0.02fF
C26022 AND2X1_LOC_44/Y OR2X1_LOC_523/a_8_216# 0.01fF
C26023 OR2X1_LOC_185/A OR2X1_LOC_270/Y 0.02fF
C26024 AND2X1_LOC_425/a_36_24# INPUT_6 0.00fF
C26025 OR2X1_LOC_95/Y AND2X1_LOC_464/a_36_24# 0.00fF
C26026 OR2X1_LOC_471/Y OR2X1_LOC_564/A 0.04fF
C26027 OR2X1_LOC_255/a_36_216# OR2X1_LOC_753/A 0.01fF
C26028 OR2X1_LOC_296/a_36_216# OR2X1_LOC_62/B 0.00fF
C26029 OR2X1_LOC_43/A OR2X1_LOC_31/Y 0.38fF
C26030 AND2X1_LOC_472/B OR2X1_LOC_408/Y 0.16fF
C26031 OR2X1_LOC_273/a_8_216# OR2X1_LOC_246/A 0.13fF
C26032 OR2X1_LOC_22/A OR2X1_LOC_17/Y 0.16fF
C26033 OR2X1_LOC_473/Y OR2X1_LOC_206/A 0.00fF
C26034 OR2X1_LOC_703/A AND2X1_LOC_31/Y 0.03fF
C26035 OR2X1_LOC_589/A OR2X1_LOC_320/a_8_216# 0.07fF
C26036 AND2X1_LOC_815/a_8_24# OR2X1_LOC_814/A 0.01fF
C26037 AND2X1_LOC_319/A OR2X1_LOC_47/Y 0.16fF
C26038 AND2X1_LOC_539/Y AND2X1_LOC_802/B 0.61fF
C26039 D_INPUT_3 OR2X1_LOC_93/a_8_216# 0.01fF
C26040 OR2X1_LOC_696/A AND2X1_LOC_809/a_8_24# 0.03fF
C26041 OR2X1_LOC_557/A AND2X1_LOC_47/Y 0.00fF
C26042 OR2X1_LOC_666/A OR2X1_LOC_13/B 0.02fF
C26043 OR2X1_LOC_650/Y AND2X1_LOC_518/a_8_24# 0.04fF
C26044 AND2X1_LOC_315/a_8_24# OR2X1_LOC_318/B 0.00fF
C26045 OR2X1_LOC_230/Y AND2X1_LOC_231/a_8_24# 0.01fF
C26046 AND2X1_LOC_339/a_8_24# AND2X1_LOC_476/A 0.03fF
C26047 OR2X1_LOC_476/B AND2X1_LOC_48/A 0.07fF
C26048 AND2X1_LOC_866/A OR2X1_LOC_757/Y 0.02fF
C26049 AND2X1_LOC_543/Y AND2X1_LOC_464/A 0.01fF
C26050 OR2X1_LOC_678/Y OR2X1_LOC_446/B 0.08fF
C26051 AND2X1_LOC_227/Y AND2X1_LOC_276/Y 0.16fF
C26052 OR2X1_LOC_613/Y AND2X1_LOC_624/B 0.02fF
C26053 OR2X1_LOC_125/Y AND2X1_LOC_128/a_8_24# 0.23fF
C26054 OR2X1_LOC_362/B D_GATE_579 0.73fF
C26055 OR2X1_LOC_650/Y AND2X1_LOC_48/A 0.09fF
C26056 AND2X1_LOC_304/a_8_24# OR2X1_LOC_446/B 0.04fF
C26057 AND2X1_LOC_318/Y OR2X1_LOC_74/A 0.02fF
C26058 OR2X1_LOC_26/Y OR2X1_LOC_289/Y 0.03fF
C26059 AND2X1_LOC_382/a_8_24# OR2X1_LOC_774/B 0.04fF
C26060 AND2X1_LOC_715/A OR2X1_LOC_268/Y 0.02fF
C26061 OR2X1_LOC_644/a_8_216# AND2X1_LOC_48/A 0.02fF
C26062 OR2X1_LOC_34/B D_INPUT_0 0.01fF
C26063 OR2X1_LOC_60/a_8_216# OR2X1_LOC_31/Y 0.01fF
C26064 AND2X1_LOC_715/Y AND2X1_LOC_809/a_8_24# 0.01fF
C26065 OR2X1_LOC_741/Y AND2X1_LOC_36/Y 0.03fF
C26066 AND2X1_LOC_849/A OR2X1_LOC_71/Y 0.02fF
C26067 OR2X1_LOC_6/A OR2X1_LOC_28/a_8_216# -0.00fF
C26068 OR2X1_LOC_648/A OR2X1_LOC_593/B 0.02fF
C26069 OR2X1_LOC_576/A AND2X1_LOC_44/Y 0.06fF
C26070 OR2X1_LOC_572/a_8_216# OR2X1_LOC_161/B 0.01fF
C26071 AND2X1_LOC_86/Y OR2X1_LOC_80/A 0.16fF
C26072 OR2X1_LOC_628/Y AND2X1_LOC_632/A 0.04fF
C26073 AND2X1_LOC_338/Y AND2X1_LOC_351/a_8_24# 0.03fF
C26074 OR2X1_LOC_648/a_8_216# OR2X1_LOC_814/A 0.14fF
C26075 OR2X1_LOC_857/B OR2X1_LOC_175/Y 0.08fF
C26076 AND2X1_LOC_12/Y OR2X1_LOC_68/B 5.00fF
C26077 INPUT_3 OR2X1_LOC_80/A 0.23fF
C26078 OR2X1_LOC_506/B AND2X1_LOC_51/Y 0.39fF
C26079 OR2X1_LOC_628/Y OR2X1_LOC_417/A 0.04fF
C26080 OR2X1_LOC_316/a_8_216# OR2X1_LOC_58/Y 0.01fF
C26081 AND2X1_LOC_232/a_8_24# AND2X1_LOC_36/Y 0.00fF
C26082 OR2X1_LOC_510/Y OR2X1_LOC_560/A 0.04fF
C26083 AND2X1_LOC_716/Y OR2X1_LOC_13/B 0.07fF
C26084 AND2X1_LOC_831/Y OR2X1_LOC_46/A 0.45fF
C26085 OR2X1_LOC_12/Y AND2X1_LOC_219/A 0.07fF
C26086 OR2X1_LOC_70/Y OR2X1_LOC_430/Y 0.01fF
C26087 OR2X1_LOC_160/B OR2X1_LOC_115/B 0.03fF
C26088 AND2X1_LOC_804/a_36_24# OR2X1_LOC_52/B 0.00fF
C26089 AND2X1_LOC_477/Y AND2X1_LOC_804/A 0.01fF
C26090 AND2X1_LOC_672/a_8_24# OR2X1_LOC_54/Y 0.03fF
C26091 AND2X1_LOC_654/Y OR2X1_LOC_13/B 0.09fF
C26092 OR2X1_LOC_87/A OR2X1_LOC_341/a_8_216# 0.14fF
C26093 VDD OR2X1_LOC_415/Y 0.50fF
C26094 AND2X1_LOC_181/Y OR2X1_LOC_522/a_8_216# 0.06fF
C26095 OR2X1_LOC_36/Y AND2X1_LOC_796/A 0.01fF
C26096 OR2X1_LOC_70/Y AND2X1_LOC_795/Y 0.05fF
C26097 AND2X1_LOC_358/Y AND2X1_LOC_566/B 0.00fF
C26098 AND2X1_LOC_464/A OR2X1_LOC_322/Y 0.01fF
C26099 OR2X1_LOC_673/B OR2X1_LOC_673/a_8_216# 0.05fF
C26100 AND2X1_LOC_71/a_36_24# OR2X1_LOC_844/B 0.00fF
C26101 OR2X1_LOC_659/Y OR2X1_LOC_113/B 0.01fF
C26102 AND2X1_LOC_17/Y AND2X1_LOC_31/Y 0.80fF
C26103 OR2X1_LOC_833/Y OR2X1_LOC_549/A 0.00fF
C26104 OR2X1_LOC_269/B OR2X1_LOC_561/B 0.01fF
C26105 AND2X1_LOC_476/Y OR2X1_LOC_323/a_36_216# 0.04fF
C26106 OR2X1_LOC_505/a_8_216# OR2X1_LOC_528/Y 0.14fF
C26107 AND2X1_LOC_117/a_8_24# OR2X1_LOC_598/A 0.02fF
C26108 AND2X1_LOC_392/A OR2X1_LOC_176/Y 0.03fF
C26109 OR2X1_LOC_22/A OR2X1_LOC_588/A 0.02fF
C26110 AND2X1_LOC_476/a_8_24# OR2X1_LOC_56/A 0.03fF
C26111 VDD AND2X1_LOC_786/Y 1.35fF
C26112 AND2X1_LOC_852/Y OR2X1_LOC_71/A 0.98fF
C26113 AND2X1_LOC_392/A OR2X1_LOC_533/Y 0.15fF
C26114 OR2X1_LOC_98/A OR2X1_LOC_415/Y 0.13fF
C26115 VDD OR2X1_LOC_323/a_8_216# 0.21fF
C26116 OR2X1_LOC_51/Y OR2X1_LOC_744/Y 0.01fF
C26117 OR2X1_LOC_129/a_8_216# OR2X1_LOC_589/A 0.01fF
C26118 AND2X1_LOC_392/A AND2X1_LOC_212/Y 0.10fF
C26119 OR2X1_LOC_248/a_8_216# OR2X1_LOC_437/A 0.03fF
C26120 AND2X1_LOC_390/B OR2X1_LOC_534/Y 0.01fF
C26121 OR2X1_LOC_206/a_8_216# AND2X1_LOC_31/Y 0.01fF
C26122 AND2X1_LOC_170/B OR2X1_LOC_47/Y 0.03fF
C26123 AND2X1_LOC_658/A OR2X1_LOC_12/Y 0.39fF
C26124 OR2X1_LOC_158/A OR2X1_LOC_96/Y 0.01fF
C26125 AND2X1_LOC_547/Y AND2X1_LOC_475/Y 0.23fF
C26126 AND2X1_LOC_64/Y AND2X1_LOC_423/a_8_24# 0.05fF
C26127 OR2X1_LOC_45/B AND2X1_LOC_675/Y 0.19fF
C26128 OR2X1_LOC_274/a_8_216# AND2X1_LOC_7/B 0.03fF
C26129 OR2X1_LOC_691/B OR2X1_LOC_35/Y 0.05fF
C26130 AND2X1_LOC_848/a_36_24# AND2X1_LOC_789/Y 0.01fF
C26131 OR2X1_LOC_744/A AND2X1_LOC_771/a_8_24# 0.01fF
C26132 AND2X1_LOC_212/A AND2X1_LOC_335/Y 0.16fF
C26133 OR2X1_LOC_6/B AND2X1_LOC_262/a_36_24# 0.00fF
C26134 OR2X1_LOC_678/a_36_216# AND2X1_LOC_44/Y 0.00fF
C26135 AND2X1_LOC_294/a_8_24# OR2X1_LOC_437/A 0.04fF
C26136 AND2X1_LOC_444/a_8_24# AND2X1_LOC_727/B 0.01fF
C26137 AND2X1_LOC_392/A AND2X1_LOC_352/a_8_24# 0.02fF
C26138 OR2X1_LOC_312/Y OR2X1_LOC_13/B 0.07fF
C26139 AND2X1_LOC_41/A AND2X1_LOC_44/Y 0.40fF
C26140 AND2X1_LOC_857/Y AND2X1_LOC_231/a_8_24# 0.01fF
C26141 AND2X1_LOC_91/B OR2X1_LOC_575/A 0.10fF
C26142 OR2X1_LOC_158/A AND2X1_LOC_454/a_8_24# 0.01fF
C26143 AND2X1_LOC_43/B AND2X1_LOC_409/B 0.07fF
C26144 AND2X1_LOC_195/a_8_24# INPUT_0 0.01fF
C26145 OR2X1_LOC_175/Y AND2X1_LOC_57/a_8_24# 0.03fF
C26146 AND2X1_LOC_363/a_8_24# OR2X1_LOC_91/A 0.05fF
C26147 OR2X1_LOC_158/A AND2X1_LOC_663/A 0.08fF
C26148 AND2X1_LOC_353/a_8_24# OR2X1_LOC_56/A 0.00fF
C26149 OR2X1_LOC_858/A OR2X1_LOC_362/A 0.05fF
C26150 OR2X1_LOC_791/A OR2X1_LOC_756/a_8_216# 0.47fF
C26151 OR2X1_LOC_47/Y AND2X1_LOC_721/A 0.05fF
C26152 AND2X1_LOC_7/B OR2X1_LOC_724/a_8_216# 0.01fF
C26153 OR2X1_LOC_161/A AND2X1_LOC_258/a_8_24# 0.01fF
C26154 OR2X1_LOC_811/A OR2X1_LOC_366/B 0.03fF
C26155 AND2X1_LOC_53/Y OR2X1_LOC_512/Y 0.02fF
C26156 AND2X1_LOC_60/a_36_24# OR2X1_LOC_61/B 0.00fF
C26157 OR2X1_LOC_524/Y AND2X1_LOC_479/a_8_24# 0.04fF
C26158 OR2X1_LOC_302/a_8_216# AND2X1_LOC_110/Y 0.01fF
C26159 VDD AND2X1_LOC_218/Y 0.38fF
C26160 OR2X1_LOC_329/Y AND2X1_LOC_512/Y 0.02fF
C26161 AND2X1_LOC_522/a_8_24# AND2X1_LOC_95/Y 0.01fF
C26162 OR2X1_LOC_244/A OR2X1_LOC_80/A 1.34fF
C26163 AND2X1_LOC_61/Y OR2X1_LOC_59/Y 0.04fF
C26164 VDD OR2X1_LOC_632/Y 0.47fF
C26165 OR2X1_LOC_222/a_8_216# OR2X1_LOC_228/Y 0.01fF
C26166 OR2X1_LOC_243/B OR2X1_LOC_71/A 0.01fF
C26167 OR2X1_LOC_161/A OR2X1_LOC_708/a_8_216# 0.04fF
C26168 VDD OR2X1_LOC_524/Y 2.11fF
C26169 OR2X1_LOC_662/A AND2X1_LOC_44/Y 0.03fF
C26170 OR2X1_LOC_288/a_8_216# OR2X1_LOC_580/B 0.11fF
C26171 AND2X1_LOC_362/a_36_24# OR2X1_LOC_494/Y 0.01fF
C26172 OR2X1_LOC_158/A OR2X1_LOC_2/Y 0.14fF
C26173 AND2X1_LOC_366/A AND2X1_LOC_366/a_8_24# 0.01fF
C26174 AND2X1_LOC_340/Y AND2X1_LOC_573/A 0.02fF
C26175 OR2X1_LOC_51/Y AND2X1_LOC_474/A 0.01fF
C26176 OR2X1_LOC_315/Y AND2X1_LOC_786/Y 0.07fF
C26177 OR2X1_LOC_756/B OR2X1_LOC_190/A 0.03fF
C26178 OR2X1_LOC_459/B OR2X1_LOC_375/Y 0.00fF
C26179 OR2X1_LOC_18/Y AND2X1_LOC_795/a_36_24# 0.00fF
C26180 AND2X1_LOC_72/Y OR2X1_LOC_344/A 0.00fF
C26181 OR2X1_LOC_600/A OR2X1_LOC_251/a_8_216# 0.02fF
C26182 AND2X1_LOC_798/a_8_24# AND2X1_LOC_337/B 0.17fF
C26183 OR2X1_LOC_47/Y OR2X1_LOC_331/Y 0.07fF
C26184 AND2X1_LOC_830/a_36_24# OR2X1_LOC_142/Y 0.01fF
C26185 OR2X1_LOC_160/B OR2X1_LOC_840/A 0.05fF
C26186 OR2X1_LOC_70/Y AND2X1_LOC_439/a_8_24# 0.01fF
C26187 OR2X1_LOC_112/a_8_216# OR2X1_LOC_624/A 0.03fF
C26188 OR2X1_LOC_715/B OR2X1_LOC_620/Y 0.33fF
C26189 OR2X1_LOC_86/A AND2X1_LOC_216/A 0.20fF
C26190 OR2X1_LOC_89/A AND2X1_LOC_783/B 0.00fF
C26191 OR2X1_LOC_707/B OR2X1_LOC_707/a_8_216# 0.01fF
C26192 OR2X1_LOC_687/Y OR2X1_LOC_691/Y 0.15fF
C26193 AND2X1_LOC_212/A OR2X1_LOC_619/Y 0.04fF
C26194 OR2X1_LOC_426/B OR2X1_LOC_298/a_36_216# 0.02fF
C26195 OR2X1_LOC_497/Y AND2X1_LOC_244/A 0.01fF
C26196 OR2X1_LOC_532/B OR2X1_LOC_550/B 0.03fF
C26197 OR2X1_LOC_426/B OR2X1_LOC_426/A 0.15fF
C26198 OR2X1_LOC_215/a_8_216# OR2X1_LOC_641/B 0.39fF
C26199 AND2X1_LOC_99/A AND2X1_LOC_243/Y 0.09fF
C26200 OR2X1_LOC_612/Y AND2X1_LOC_647/a_8_24# 0.23fF
C26201 AND2X1_LOC_95/Y OR2X1_LOC_730/A 0.01fF
C26202 OR2X1_LOC_158/A AND2X1_LOC_449/Y 0.01fF
C26203 INPUT_1 OR2X1_LOC_749/Y 0.13fF
C26204 OR2X1_LOC_687/Y OR2X1_LOC_713/A 0.03fF
C26205 AND2X1_LOC_588/a_8_24# OR2X1_LOC_502/A 0.03fF
C26206 OR2X1_LOC_643/A OR2X1_LOC_161/B 0.03fF
C26207 OR2X1_LOC_45/Y OR2X1_LOC_600/A 0.43fF
C26208 OR2X1_LOC_814/A OR2X1_LOC_579/A 0.15fF
C26209 OR2X1_LOC_335/Y OR2X1_LOC_352/A 0.00fF
C26210 AND2X1_LOC_724/Y OR2X1_LOC_48/B 0.02fF
C26211 OR2X1_LOC_124/Y OR2X1_LOC_161/B 0.02fF
C26212 OR2X1_LOC_778/Y OR2X1_LOC_161/B 0.10fF
C26213 OR2X1_LOC_790/B AND2X1_LOC_18/Y 0.23fF
C26214 AND2X1_LOC_58/a_8_24# OR2X1_LOC_78/B 0.01fF
C26215 OR2X1_LOC_18/Y AND2X1_LOC_806/a_8_24# 0.02fF
C26216 OR2X1_LOC_668/a_8_216# OR2X1_LOC_244/Y 0.12fF
C26217 OR2X1_LOC_161/A AND2X1_LOC_18/Y 0.15fF
C26218 AND2X1_LOC_765/a_8_24# OR2X1_LOC_401/Y 0.01fF
C26219 OR2X1_LOC_715/B OR2X1_LOC_154/A 0.10fF
C26220 AND2X1_LOC_787/a_8_24# OR2X1_LOC_59/Y 0.02fF
C26221 OR2X1_LOC_810/A OR2X1_LOC_435/A 0.03fF
C26222 OR2X1_LOC_91/Y OR2X1_LOC_40/Y 0.40fF
C26223 AND2X1_LOC_41/A OR2X1_LOC_61/a_8_216# 0.02fF
C26224 OR2X1_LOC_51/Y AND2X1_LOC_593/Y 0.65fF
C26225 OR2X1_LOC_379/a_8_216# OR2X1_LOC_66/A 0.01fF
C26226 AND2X1_LOC_647/B OR2X1_LOC_71/A 0.02fF
C26227 AND2X1_LOC_16/a_8_24# OR2X1_LOC_78/B 0.05fF
C26228 AND2X1_LOC_857/Y AND2X1_LOC_863/a_8_24# 0.00fF
C26229 OR2X1_LOC_352/A AND2X1_LOC_40/Y 0.28fF
C26230 OR2X1_LOC_551/B OR2X1_LOC_364/Y 0.07fF
C26231 OR2X1_LOC_790/A OR2X1_LOC_269/B 0.01fF
C26232 OR2X1_LOC_159/a_36_216# OR2X1_LOC_6/A 0.03fF
C26233 OR2X1_LOC_160/B OR2X1_LOC_222/A 0.07fF
C26234 OR2X1_LOC_323/A AND2X1_LOC_465/Y 0.00fF
C26235 AND2X1_LOC_40/Y OR2X1_LOC_434/a_36_216# 0.00fF
C26236 OR2X1_LOC_814/A OR2X1_LOC_390/B 0.10fF
C26237 OR2X1_LOC_421/A OR2X1_LOC_44/Y 0.15fF
C26238 OR2X1_LOC_574/A OR2X1_LOC_549/A 0.10fF
C26239 OR2X1_LOC_696/A D_INPUT_0 0.94fF
C26240 AND2X1_LOC_589/a_8_24# OR2X1_LOC_435/A 0.01fF
C26241 AND2X1_LOC_362/a_8_24# OR2X1_LOC_18/Y 0.02fF
C26242 OR2X1_LOC_185/A INPUT_0 0.17fF
C26243 OR2X1_LOC_377/A OR2X1_LOC_78/B 4.27fF
C26244 OR2X1_LOC_70/Y AND2X1_LOC_636/a_36_24# 0.01fF
C26245 OR2X1_LOC_604/A OR2X1_LOC_418/Y 0.38fF
C26246 AND2X1_LOC_777/a_8_24# VDD 0.00fF
C26247 AND2X1_LOC_580/A AND2X1_LOC_657/Y 0.03fF
C26248 AND2X1_LOC_776/a_8_24# AND2X1_LOC_840/B 0.10fF
C26249 AND2X1_LOC_523/Y AND2X1_LOC_445/a_8_24# 0.01fF
C26250 OR2X1_LOC_51/Y OR2X1_LOC_85/A 0.10fF
C26251 OR2X1_LOC_452/a_8_216# OR2X1_LOC_449/B 0.04fF
C26252 AND2X1_LOC_191/B AND2X1_LOC_580/A 0.00fF
C26253 AND2X1_LOC_64/Y D_INPUT_0 0.93fF
C26254 OR2X1_LOC_236/a_8_216# OR2X1_LOC_56/A 0.46fF
C26255 AND2X1_LOC_794/B AND2X1_LOC_578/A 0.05fF
C26256 OR2X1_LOC_634/A AND2X1_LOC_43/B 0.11fF
C26257 OR2X1_LOC_117/a_8_216# OR2X1_LOC_19/B 0.01fF
C26258 AND2X1_LOC_388/Y AND2X1_LOC_390/B 0.07fF
C26259 OR2X1_LOC_685/B AND2X1_LOC_681/a_36_24# 0.00fF
C26260 OR2X1_LOC_426/B AND2X1_LOC_100/a_8_24# 0.01fF
C26261 OR2X1_LOC_864/A AND2X1_LOC_70/Y 0.03fF
C26262 AND2X1_LOC_12/Y OR2X1_LOC_834/a_8_216# 0.02fF
C26263 OR2X1_LOC_763/Y VDD 0.08fF
C26264 OR2X1_LOC_331/A OR2X1_LOC_26/Y 0.04fF
C26265 OR2X1_LOC_628/a_8_216# OR2X1_LOC_427/A 0.02fF
C26266 OR2X1_LOC_479/Y OR2X1_LOC_182/B 0.03fF
C26267 AND2X1_LOC_346/a_8_24# OR2X1_LOC_481/A 0.01fF
C26268 OR2X1_LOC_369/a_36_216# AND2X1_LOC_211/B 0.00fF
C26269 AND2X1_LOC_862/Y AND2X1_LOC_807/Y 0.02fF
C26270 VDD OR2X1_LOC_378/Y 0.06fF
C26271 OR2X1_LOC_426/B AND2X1_LOC_123/a_8_24# 0.03fF
C26272 AND2X1_LOC_852/Y OR2X1_LOC_59/Y 0.06fF
C26273 OR2X1_LOC_7/A AND2X1_LOC_285/Y 0.03fF
C26274 AND2X1_LOC_658/A OR2X1_LOC_239/a_8_216# 0.03fF
C26275 OR2X1_LOC_759/A OR2X1_LOC_74/A 0.03fF
C26276 AND2X1_LOC_218/a_8_24# OR2X1_LOC_272/Y 0.02fF
C26277 OR2X1_LOC_486/B OR2X1_LOC_726/A 0.08fF
C26278 AND2X1_LOC_70/Y OR2X1_LOC_633/B 0.03fF
C26279 AND2X1_LOC_570/Y OR2X1_LOC_89/A 0.08fF
C26280 OR2X1_LOC_287/B AND2X1_LOC_397/a_8_24# 0.01fF
C26281 AND2X1_LOC_391/Y OR2X1_LOC_585/A 0.03fF
C26282 OR2X1_LOC_40/Y OR2X1_LOC_527/Y 0.03fF
C26283 VDD AND2X1_LOC_578/A 0.14fF
C26284 AND2X1_LOC_456/B OR2X1_LOC_44/Y 0.00fF
C26285 OR2X1_LOC_585/A AND2X1_LOC_637/a_36_24# -0.01fF
C26286 OR2X1_LOC_91/A OR2X1_LOC_585/A 0.06fF
C26287 AND2X1_LOC_456/B AND2X1_LOC_288/a_8_24# 0.17fF
C26288 OR2X1_LOC_805/A OR2X1_LOC_734/a_36_216# 0.01fF
C26289 OR2X1_LOC_656/B OR2X1_LOC_559/B 0.05fF
C26290 OR2X1_LOC_203/Y OR2X1_LOC_721/Y 0.10fF
C26291 AND2X1_LOC_51/Y AND2X1_LOC_18/Y 0.11fF
C26292 OR2X1_LOC_840/a_8_216# OR2X1_LOC_814/A 0.04fF
C26293 OR2X1_LOC_40/Y OR2X1_LOC_291/Y 0.05fF
C26294 AND2X1_LOC_510/a_8_24# AND2X1_LOC_474/Y 0.01fF
C26295 VDD OR2X1_LOC_285/B 0.21fF
C26296 OR2X1_LOC_719/A OR2X1_LOC_66/A 0.09fF
C26297 OR2X1_LOC_147/B OR2X1_LOC_87/A 0.03fF
C26298 AND2X1_LOC_725/a_8_24# AND2X1_LOC_712/B 0.10fF
C26299 AND2X1_LOC_347/a_36_24# OR2X1_LOC_59/Y 0.00fF
C26300 OR2X1_LOC_6/B OR2X1_LOC_46/A 0.30fF
C26301 OR2X1_LOC_479/Y OR2X1_LOC_168/B 0.07fF
C26302 OR2X1_LOC_40/Y AND2X1_LOC_574/A 0.04fF
C26303 AND2X1_LOC_56/B OR2X1_LOC_811/A 0.03fF
C26304 AND2X1_LOC_364/A AND2X1_LOC_354/B 0.49fF
C26305 OR2X1_LOC_500/A OR2X1_LOC_161/A 0.18fF
C26306 OR2X1_LOC_377/A OR2X1_LOC_375/A 0.49fF
C26307 AND2X1_LOC_535/a_8_24# OR2X1_LOC_417/Y 0.04fF
C26308 OR2X1_LOC_600/A AND2X1_LOC_727/A 0.03fF
C26309 OR2X1_LOC_866/B D_INPUT_1 0.10fF
C26310 OR2X1_LOC_70/A OR2X1_LOC_387/A 0.32fF
C26311 VDD AND2X1_LOC_635/a_8_24# 0.00fF
C26312 AND2X1_LOC_810/A AND2X1_LOC_318/Y 0.02fF
C26313 OR2X1_LOC_237/a_36_216# OR2X1_LOC_237/Y 0.00fF
C26314 AND2X1_LOC_729/a_8_24# OR2X1_LOC_95/Y 0.01fF
C26315 OR2X1_LOC_270/Y OR2X1_LOC_577/Y 0.01fF
C26316 INPUT_3 OR2X1_LOC_6/A 0.21fF
C26317 AND2X1_LOC_824/B OR2X1_LOC_375/A 0.06fF
C26318 AND2X1_LOC_40/Y OR2X1_LOC_646/a_8_216# 0.01fF
C26319 OR2X1_LOC_631/a_36_216# OR2X1_LOC_631/B 0.01fF
C26320 OR2X1_LOC_777/B OR2X1_LOC_446/B 0.02fF
C26321 OR2X1_LOC_207/a_8_216# AND2X1_LOC_44/Y 0.14fF
C26322 AND2X1_LOC_364/Y AND2X1_LOC_326/A 0.01fF
C26323 OR2X1_LOC_824/Y OR2X1_LOC_619/Y 0.72fF
C26324 OR2X1_LOC_22/Y AND2X1_LOC_436/Y 0.08fF
C26325 OR2X1_LOC_51/Y AND2X1_LOC_470/a_8_24# 0.01fF
C26326 OR2X1_LOC_400/a_36_216# OR2X1_LOC_557/A 0.00fF
C26327 OR2X1_LOC_771/B OR2X1_LOC_71/A 0.03fF
C26328 OR2X1_LOC_777/B OR2X1_LOC_303/B 0.05fF
C26329 OR2X1_LOC_194/B OR2X1_LOC_155/A 0.07fF
C26330 OR2X1_LOC_806/a_8_216# OR2X1_LOC_269/B 0.01fF
C26331 OR2X1_LOC_391/B OR2X1_LOC_773/B 0.04fF
C26332 OR2X1_LOC_203/Y OR2X1_LOC_375/A 0.11fF
C26333 OR2X1_LOC_358/a_8_216# OR2X1_LOC_358/B 0.02fF
C26334 AND2X1_LOC_63/a_8_24# OR2X1_LOC_204/Y 0.01fF
C26335 OR2X1_LOC_849/A AND2X1_LOC_132/a_8_24# 0.23fF
C26336 AND2X1_LOC_851/B AND2X1_LOC_476/Y 0.02fF
C26337 OR2X1_LOC_276/A AND2X1_LOC_275/a_36_24# 0.00fF
C26338 AND2X1_LOC_33/a_8_24# D_INPUT_0 0.01fF
C26339 AND2X1_LOC_573/A OR2X1_LOC_585/A 0.34fF
C26340 OR2X1_LOC_287/B OR2X1_LOC_362/B 0.00fF
C26341 OR2X1_LOC_691/Y OR2X1_LOC_644/A 0.31fF
C26342 OR2X1_LOC_626/a_8_216# OR2X1_LOC_39/A 0.01fF
C26343 OR2X1_LOC_600/A OR2X1_LOC_95/Y 0.88fF
C26344 OR2X1_LOC_40/Y D_INPUT_3 0.03fF
C26345 OR2X1_LOC_788/B OR2X1_LOC_535/a_8_216# 0.01fF
C26346 OR2X1_LOC_18/Y OR2X1_LOC_371/Y 0.08fF
C26347 OR2X1_LOC_841/a_8_216# OR2X1_LOC_121/B 0.01fF
C26348 OR2X1_LOC_405/A OR2X1_LOC_592/A 0.09fF
C26349 OR2X1_LOC_219/B OR2X1_LOC_222/A 0.17fF
C26350 OR2X1_LOC_248/a_8_216# OR2X1_LOC_753/A 0.01fF
C26351 OR2X1_LOC_91/Y OR2X1_LOC_7/A 0.10fF
C26352 OR2X1_LOC_598/A OR2X1_LOC_548/a_8_216# 0.01fF
C26353 AND2X1_LOC_41/A OR2X1_LOC_720/B 0.03fF
C26354 AND2X1_LOC_43/a_36_24# AND2X1_LOC_43/B 0.01fF
C26355 OR2X1_LOC_3/Y OR2X1_LOC_316/Y 0.03fF
C26356 OR2X1_LOC_81/a_8_216# OR2X1_LOC_52/B 0.03fF
C26357 OR2X1_LOC_768/A AND2X1_LOC_47/Y 0.00fF
C26358 AND2X1_LOC_494/a_36_24# OR2X1_LOC_391/A -0.01fF
C26359 OR2X1_LOC_313/Y OR2X1_LOC_418/a_36_216# 0.00fF
C26360 OR2X1_LOC_3/Y OR2X1_LOC_595/a_36_216# 0.01fF
C26361 OR2X1_LOC_649/B AND2X1_LOC_8/Y 0.05fF
C26362 VDD AND2X1_LOC_114/Y 0.21fF
C26363 AND2X1_LOC_563/a_36_24# OR2X1_LOC_89/A 0.00fF
C26364 INPUT_1 AND2X1_LOC_820/B 0.01fF
C26365 AND2X1_LOC_59/Y OR2X1_LOC_479/Y 0.09fF
C26366 OR2X1_LOC_602/a_8_216# AND2X1_LOC_43/B 0.03fF
C26367 OR2X1_LOC_791/B AND2X1_LOC_281/a_8_24# 0.01fF
C26368 OR2X1_LOC_305/Y OR2X1_LOC_7/A 0.03fF
C26369 OR2X1_LOC_139/a_36_216# OR2X1_LOC_267/A 0.00fF
C26370 OR2X1_LOC_441/Y OR2X1_LOC_679/A 0.03fF
C26371 AND2X1_LOC_387/B OR2X1_LOC_87/A 0.03fF
C26372 AND2X1_LOC_294/a_8_24# OR2X1_LOC_753/A 0.01fF
C26373 OR2X1_LOC_512/A D_INPUT_0 0.06fF
C26374 AND2X1_LOC_71/a_8_24# AND2X1_LOC_47/Y 0.10fF
C26375 OR2X1_LOC_599/A OR2X1_LOC_696/a_8_216# 0.03fF
C26376 OR2X1_LOC_615/Y OR2X1_LOC_56/A 0.12fF
C26377 OR2X1_LOC_3/Y AND2X1_LOC_404/a_8_24# 0.01fF
C26378 VDD OR2X1_LOC_213/a_8_216# 0.00fF
C26379 AND2X1_LOC_543/a_8_24# OR2X1_LOC_95/Y 0.01fF
C26380 OR2X1_LOC_186/Y OR2X1_LOC_567/a_8_216# 0.00fF
C26381 AND2X1_LOC_566/Y OR2X1_LOC_26/Y 0.02fF
C26382 OR2X1_LOC_124/A OR2X1_LOC_786/Y 0.01fF
C26383 AND2X1_LOC_727/A OR2X1_LOC_619/Y 0.06fF
C26384 OR2X1_LOC_566/A OR2X1_LOC_303/B 0.77fF
C26385 OR2X1_LOC_154/A AND2X1_LOC_689/a_8_24# 0.01fF
C26386 OR2X1_LOC_494/a_8_216# AND2X1_LOC_866/A -0.02fF
C26387 AND2X1_LOC_491/a_8_24# OR2X1_LOC_805/A 0.03fF
C26388 AND2X1_LOC_91/B OR2X1_LOC_704/a_36_216# 0.00fF
C26389 OR2X1_LOC_438/Y AND2X1_LOC_675/A 0.01fF
C26390 AND2X1_LOC_465/A OR2X1_LOC_437/A 0.17fF
C26391 OR2X1_LOC_865/B OR2X1_LOC_814/A 0.01fF
C26392 OR2X1_LOC_427/A INPUT_1 0.16fF
C26393 AND2X1_LOC_710/a_36_24# AND2X1_LOC_789/Y 0.01fF
C26394 OR2X1_LOC_773/B OR2X1_LOC_772/Y 0.06fF
C26395 OR2X1_LOC_278/A AND2X1_LOC_633/a_8_24# 0.07fF
C26396 OR2X1_LOC_84/B OR2X1_LOC_204/a_8_216# 0.03fF
C26397 OR2X1_LOC_270/a_8_216# OR2X1_LOC_456/A 0.00fF
C26398 AND2X1_LOC_753/B OR2X1_LOC_197/A 0.05fF
C26399 OR2X1_LOC_114/B AND2X1_LOC_497/a_36_24# 0.00fF
C26400 OR2X1_LOC_392/B OR2X1_LOC_140/Y 0.03fF
C26401 OR2X1_LOC_542/a_36_216# OR2X1_LOC_552/A 0.00fF
C26402 AND2X1_LOC_500/Y OR2X1_LOC_419/Y 0.37fF
C26403 OR2X1_LOC_486/Y OR2X1_LOC_578/B 9.76fF
C26404 AND2X1_LOC_753/a_8_24# AND2X1_LOC_53/Y 0.02fF
C26405 AND2X1_LOC_357/A AND2X1_LOC_222/Y 0.00fF
C26406 OR2X1_LOC_702/A AND2X1_LOC_3/Y 0.03fF
C26407 AND2X1_LOC_560/B AND2X1_LOC_523/Y 1.20fF
C26408 AND2X1_LOC_139/B OR2X1_LOC_46/A 0.03fF
C26409 OR2X1_LOC_864/A OR2X1_LOC_404/Y 0.03fF
C26410 VDD OR2X1_LOC_358/A 0.25fF
C26411 OR2X1_LOC_715/B OR2X1_LOC_560/A 0.03fF
C26412 OR2X1_LOC_66/A OR2X1_LOC_675/Y 4.41fF
C26413 OR2X1_LOC_287/B OR2X1_LOC_846/B 0.00fF
C26414 VDD OR2X1_LOC_170/Y -0.00fF
C26415 OR2X1_LOC_832/a_8_216# AND2X1_LOC_31/Y 0.01fF
C26416 VDD OR2X1_LOC_88/a_8_216# 0.00fF
C26417 OR2X1_LOC_160/A OR2X1_LOC_446/Y 0.06fF
C26418 OR2X1_LOC_95/Y OR2X1_LOC_619/Y 0.03fF
C26419 AND2X1_LOC_17/Y AND2X1_LOC_31/a_8_24# 0.01fF
C26420 VDD OR2X1_LOC_746/Y 0.08fF
C26421 AND2X1_LOC_675/A AND2X1_LOC_621/Y 0.07fF
C26422 VDD OR2X1_LOC_172/a_8_216# 0.21fF
C26423 AND2X1_LOC_776/Y AND2X1_LOC_785/A 0.02fF
C26424 OR2X1_LOC_417/Y OR2X1_LOC_7/A 0.07fF
C26425 INPUT_3 D_INPUT_2 0.76fF
C26426 OR2X1_LOC_22/Y OR2X1_LOC_588/Y 0.03fF
C26427 OR2X1_LOC_271/a_8_216# INPUT_1 0.02fF
C26428 OR2X1_LOC_545/B OR2X1_LOC_87/A 0.01fF
C26429 AND2X1_LOC_53/Y OR2X1_LOC_194/Y 0.08fF
C26430 AND2X1_LOC_32/a_36_24# D_INPUT_0 0.00fF
C26431 OR2X1_LOC_476/B AND2X1_LOC_3/Y 0.42fF
C26432 OR2X1_LOC_311/Y OR2X1_LOC_7/A 0.03fF
C26433 AND2X1_LOC_227/Y AND2X1_LOC_139/B 0.06fF
C26434 OR2X1_LOC_3/Y OR2X1_LOC_431/Y 0.03fF
C26435 OR2X1_LOC_675/a_8_216# OR2X1_LOC_76/A 0.03fF
C26436 OR2X1_LOC_759/a_8_216# AND2X1_LOC_789/Y 0.01fF
C26437 OR2X1_LOC_696/A AND2X1_LOC_539/Y 0.15fF
C26438 OR2X1_LOC_7/A AND2X1_LOC_574/A 0.01fF
C26439 OR2X1_LOC_696/A AND2X1_LOC_552/a_8_24# 0.02fF
C26440 OR2X1_LOC_475/Y OR2X1_LOC_479/a_8_216# 0.07fF
C26441 OR2X1_LOC_160/A OR2X1_LOC_473/A 0.74fF
C26442 AND2X1_LOC_44/Y INPUT_6 0.54fF
C26443 OR2X1_LOC_436/Y OR2X1_LOC_802/Y 0.01fF
C26444 OR2X1_LOC_19/B AND2X1_LOC_42/B 0.13fF
C26445 OR2X1_LOC_644/a_8_216# AND2X1_LOC_3/Y 0.01fF
C26446 OR2X1_LOC_436/Y OR2X1_LOC_468/Y 0.15fF
C26447 D_INPUT_3 OR2X1_LOC_618/a_8_216# 0.01fF
C26448 OR2X1_LOC_625/Y AND2X1_LOC_721/A 0.01fF
C26449 OR2X1_LOC_154/A AND2X1_LOC_106/a_36_24# 0.01fF
C26450 AND2X1_LOC_269/a_8_24# AND2X1_LOC_786/Y 0.04fF
C26451 AND2X1_LOC_474/Y AND2X1_LOC_657/a_36_24# 0.00fF
C26452 OR2X1_LOC_64/Y AND2X1_LOC_523/Y 0.03fF
C26453 OR2X1_LOC_448/Y OR2X1_LOC_779/Y 0.00fF
C26454 OR2X1_LOC_364/A AND2X1_LOC_109/a_8_24# 0.01fF
C26455 OR2X1_LOC_185/Y AND2X1_LOC_109/a_8_24# 0.06fF
C26456 OR2X1_LOC_858/a_8_216# OR2X1_LOC_580/A 0.03fF
C26457 AND2X1_LOC_539/Y AND2X1_LOC_715/Y 0.03fF
C26458 AND2X1_LOC_727/Y AND2X1_LOC_726/a_8_24# 0.01fF
C26459 AND2X1_LOC_170/Y OR2X1_LOC_47/Y 0.29fF
C26460 AND2X1_LOC_817/B OR2X1_LOC_770/Y 0.01fF
C26461 OR2X1_LOC_529/Y AND2X1_LOC_227/Y 0.01fF
C26462 OR2X1_LOC_47/Y AND2X1_LOC_361/A 0.85fF
C26463 OR2X1_LOC_131/Y AND2X1_LOC_656/Y 0.16fF
C26464 OR2X1_LOC_187/Y AND2X1_LOC_191/a_8_24# 0.23fF
C26465 OR2X1_LOC_404/Y AND2X1_LOC_134/a_36_24# 0.00fF
C26466 D_INPUT_3 OR2X1_LOC_7/A 0.24fF
C26467 OR2X1_LOC_48/B AND2X1_LOC_222/Y 0.02fF
C26468 OR2X1_LOC_847/B D_INPUT_1 0.01fF
C26469 AND2X1_LOC_157/a_36_24# OR2X1_LOC_451/B -0.00fF
C26470 AND2X1_LOC_91/B OR2X1_LOC_161/B 0.71fF
C26471 AND2X1_LOC_347/Y OR2X1_LOC_384/Y 0.03fF
C26472 OR2X1_LOC_784/Y OR2X1_LOC_779/B 0.00fF
C26473 AND2X1_LOC_91/a_8_24# OR2X1_LOC_97/A 0.01fF
C26474 AND2X1_LOC_343/a_8_24# OR2X1_LOC_47/Y 0.16fF
C26475 OR2X1_LOC_347/B OR2X1_LOC_736/a_8_216# 0.47fF
C26476 OR2X1_LOC_95/Y OR2X1_LOC_372/a_8_216# -0.01fF
C26477 AND2X1_LOC_687/a_36_24# OR2X1_LOC_52/B 0.01fF
C26478 AND2X1_LOC_477/a_8_24# OR2X1_LOC_437/A 0.03fF
C26479 OR2X1_LOC_76/Y OR2X1_LOC_241/B 0.03fF
C26480 AND2X1_LOC_22/Y AND2X1_LOC_522/a_8_24# 0.06fF
C26481 OR2X1_LOC_160/A OR2X1_LOC_228/Y 0.07fF
C26482 AND2X1_LOC_578/A OR2X1_LOC_674/Y 0.03fF
C26483 OR2X1_LOC_244/Y OR2X1_LOC_844/B 1.11fF
C26484 OR2X1_LOC_87/A OR2X1_LOC_318/B 0.03fF
C26485 OR2X1_LOC_557/A D_INPUT_1 0.03fF
C26486 OR2X1_LOC_604/A OR2X1_LOC_743/Y -0.01fF
C26487 OR2X1_LOC_703/B OR2X1_LOC_854/A 0.01fF
C26488 OR2X1_LOC_175/Y OR2X1_LOC_535/A 0.01fF
C26489 OR2X1_LOC_78/B OR2X1_LOC_539/B 0.01fF
C26490 OR2X1_LOC_154/A OR2X1_LOC_398/Y 0.05fF
C26491 OR2X1_LOC_26/Y OR2X1_LOC_406/A 0.01fF
C26492 AND2X1_LOC_64/Y OR2X1_LOC_598/Y 0.03fF
C26493 OR2X1_LOC_40/Y OR2X1_LOC_171/Y 0.07fF
C26494 VDD OR2X1_LOC_168/Y 0.24fF
C26495 AND2X1_LOC_59/Y OR2X1_LOC_68/B 0.20fF
C26496 OR2X1_LOC_6/B OR2X1_LOC_748/a_8_216# 0.10fF
C26497 AND2X1_LOC_77/a_8_24# OR2X1_LOC_62/A 0.19fF
C26498 OR2X1_LOC_696/A AND2X1_LOC_326/B 0.04fF
C26499 AND2X1_LOC_64/Y AND2X1_LOC_131/a_8_24# 0.02fF
C26500 AND2X1_LOC_483/Y OR2X1_LOC_7/A 0.56fF
C26501 OR2X1_LOC_373/a_36_216# OR2X1_LOC_373/Y 0.00fF
C26502 OR2X1_LOC_736/A OR2X1_LOC_777/B 0.14fF
C26503 AND2X1_LOC_47/Y OR2X1_LOC_46/A 0.03fF
C26504 OR2X1_LOC_48/B OR2X1_LOC_423/Y 0.03fF
C26505 AND2X1_LOC_64/Y OR2X1_LOC_356/a_8_216# 0.02fF
C26506 AND2X1_LOC_64/Y AND2X1_LOC_505/a_8_24# 0.01fF
C26507 OR2X1_LOC_235/B AND2X1_LOC_36/Y 0.07fF
C26508 OR2X1_LOC_468/Y OR2X1_LOC_566/Y 0.01fF
C26509 OR2X1_LOC_88/Y AND2X1_LOC_266/Y 0.00fF
C26510 D_INPUT_0 OR2X1_LOC_54/a_8_216# 0.02fF
C26511 OR2X1_LOC_89/A OR2X1_LOC_406/A 0.01fF
C26512 AND2X1_LOC_638/Y D_INPUT_6 0.00fF
C26513 OR2X1_LOC_161/B OR2X1_LOC_364/a_8_216# 0.03fF
C26514 AND2X1_LOC_599/a_8_24# OR2X1_LOC_598/Y 0.08fF
C26515 OR2X1_LOC_135/Y AND2X1_LOC_339/B 0.03fF
C26516 OR2X1_LOC_215/a_8_216# OR2X1_LOC_215/A 0.02fF
C26517 VDD AND2X1_LOC_202/Y 0.31fF
C26518 OR2X1_LOC_45/B OR2X1_LOC_421/A 0.04fF
C26519 AND2X1_LOC_769/a_36_24# OR2X1_LOC_426/B 0.01fF
C26520 OR2X1_LOC_375/A OR2X1_LOC_732/A 0.01fF
C26521 OR2X1_LOC_66/A OR2X1_LOC_779/A 0.74fF
C26522 OR2X1_LOC_344/A OR2X1_LOC_719/B 0.02fF
C26523 AND2X1_LOC_70/Y OR2X1_LOC_121/A 0.03fF
C26524 OR2X1_LOC_237/Y OR2X1_LOC_437/A 0.05fF
C26525 OR2X1_LOC_744/A AND2X1_LOC_780/a_36_24# 0.00fF
C26526 AND2X1_LOC_851/a_8_24# AND2X1_LOC_465/A 0.00fF
C26527 OR2X1_LOC_665/a_36_216# AND2X1_LOC_793/Y 0.01fF
C26528 OR2X1_LOC_666/A OR2X1_LOC_428/A 0.02fF
C26529 OR2X1_LOC_634/A AND2X1_LOC_416/a_8_24# 0.01fF
C26530 AND2X1_LOC_721/Y AND2X1_LOC_663/A 0.05fF
C26531 OR2X1_LOC_645/a_8_216# OR2X1_LOC_161/B 0.03fF
C26532 AND2X1_LOC_787/A OR2X1_LOC_59/Y 0.25fF
C26533 OR2X1_LOC_97/A OR2X1_LOC_78/A 0.04fF
C26534 OR2X1_LOC_542/B OR2X1_LOC_344/A 0.03fF
C26535 OR2X1_LOC_6/B OR2X1_LOC_786/a_8_216# 0.07fF
C26536 OR2X1_LOC_736/Y OR2X1_LOC_66/A 0.12fF
C26537 OR2X1_LOC_604/A AND2X1_LOC_285/a_8_24# 0.07fF
C26538 AND2X1_LOC_56/B OR2X1_LOC_777/B 0.05fF
C26539 OR2X1_LOC_814/A OR2X1_LOC_493/Y 0.03fF
C26540 OR2X1_LOC_188/Y OR2X1_LOC_756/B 0.02fF
C26541 AND2X1_LOC_64/Y AND2X1_LOC_40/Y 2.15fF
C26542 OR2X1_LOC_46/A OR2X1_LOC_598/A 1.33fF
C26543 OR2X1_LOC_13/Y AND2X1_LOC_207/B 0.01fF
C26544 OR2X1_LOC_696/A AND2X1_LOC_375/a_8_24# 0.08fF
C26545 AND2X1_LOC_214/A AND2X1_LOC_208/Y 0.04fF
C26546 OR2X1_LOC_451/a_8_216# OR2X1_LOC_452/A -0.00fF
C26547 OR2X1_LOC_666/A OR2X1_LOC_595/A 0.03fF
C26548 OR2X1_LOC_866/B OR2X1_LOC_391/a_8_216# 0.02fF
C26549 OR2X1_LOC_6/B INPUT_2 0.29fF
C26550 OR2X1_LOC_762/Y OR2X1_LOC_428/A 0.06fF
C26551 OR2X1_LOC_6/B AND2X1_LOC_403/a_8_24# 0.01fF
C26552 AND2X1_LOC_393/a_8_24# AND2X1_LOC_36/Y 0.01fF
C26553 OR2X1_LOC_681/a_8_216# VDD 0.21fF
C26554 OR2X1_LOC_158/A OR2X1_LOC_25/Y 0.89fF
C26555 OR2X1_LOC_604/A OR2X1_LOC_627/Y 0.03fF
C26556 AND2X1_LOC_388/Y OR2X1_LOC_744/A 0.01fF
C26557 AND2X1_LOC_81/B OR2X1_LOC_510/a_8_216# 0.01fF
C26558 AND2X1_LOC_716/Y OR2X1_LOC_428/A 0.07fF
C26559 OR2X1_LOC_139/A OR2X1_LOC_653/Y 0.39fF
C26560 OR2X1_LOC_641/Y OR2X1_LOC_66/A 0.03fF
C26561 AND2X1_LOC_486/Y AND2X1_LOC_786/Y 0.07fF
C26562 OR2X1_LOC_269/B OR2X1_LOC_714/a_8_216# 0.02fF
C26563 AND2X1_LOC_374/a_8_24# OR2X1_LOC_373/Y 0.00fF
C26564 AND2X1_LOC_190/a_36_24# OR2X1_LOC_108/Y 0.00fF
C26565 OR2X1_LOC_467/A OR2X1_LOC_454/a_36_216# 0.00fF
C26566 OR2X1_LOC_47/Y AND2X1_LOC_795/Y 0.03fF
C26567 AND2X1_LOC_654/Y OR2X1_LOC_428/A 0.07fF
C26568 AND2X1_LOC_21/Y D_INPUT_6 0.07fF
C26569 OR2X1_LOC_185/A AND2X1_LOC_7/B 0.08fF
C26570 AND2X1_LOC_40/Y AND2X1_LOC_82/Y 0.00fF
C26571 AND2X1_LOC_64/Y OR2X1_LOC_87/Y 0.03fF
C26572 AND2X1_LOC_534/a_36_24# OR2X1_LOC_354/A 0.00fF
C26573 OR2X1_LOC_464/a_8_216# OR2X1_LOC_542/B 0.06fF
C26574 AND2X1_LOC_656/Y AND2X1_LOC_657/A 0.11fF
C26575 AND2X1_LOC_28/a_8_24# OR2X1_LOC_80/A 0.04fF
C26576 OR2X1_LOC_756/B OR2X1_LOC_325/B 0.00fF
C26577 AND2X1_LOC_99/A OR2X1_LOC_12/Y 0.03fF
C26578 AND2X1_LOC_732/B AND2X1_LOC_605/Y 0.04fF
C26579 AND2X1_LOC_72/Y OR2X1_LOC_161/B 0.01fF
C26580 OR2X1_LOC_97/A OR2X1_LOC_602/A 0.01fF
C26581 OR2X1_LOC_502/A OR2X1_LOC_641/A 0.03fF
C26582 OR2X1_LOC_631/B OR2X1_LOC_554/a_8_216# 0.01fF
C26583 OR2X1_LOC_483/a_8_216# OR2X1_LOC_563/A 0.01fF
C26584 AND2X1_LOC_857/a_8_24# OR2X1_LOC_171/Y 0.01fF
C26585 OR2X1_LOC_669/A AND2X1_LOC_287/B 0.77fF
C26586 OR2X1_LOC_179/Y OR2X1_LOC_600/A 0.01fF
C26587 OR2X1_LOC_7/A AND2X1_LOC_780/a_8_24# 0.04fF
C26588 OR2X1_LOC_78/A OR2X1_LOC_78/a_8_216# 0.13fF
C26589 AND2X1_LOC_367/A AND2X1_LOC_367/B 0.29fF
C26590 OR2X1_LOC_854/a_8_216# AND2X1_LOC_110/Y 0.01fF
C26591 OR2X1_LOC_756/B OR2X1_LOC_862/B 0.01fF
C26592 OR2X1_LOC_7/A OR2X1_LOC_171/Y 0.03fF
C26593 OR2X1_LOC_84/a_8_216# OR2X1_LOC_398/Y 0.40fF
C26594 OR2X1_LOC_808/B OR2X1_LOC_66/A 0.02fF
C26595 OR2X1_LOC_188/Y OR2X1_LOC_76/Y 0.01fF
C26596 OR2X1_LOC_709/A OR2X1_LOC_738/A 0.10fF
C26597 AND2X1_LOC_774/a_36_24# OR2X1_LOC_306/Y 0.00fF
C26598 AND2X1_LOC_729/Y AND2X1_LOC_705/Y 0.01fF
C26599 OR2X1_LOC_691/Y OR2X1_LOC_835/B 0.83fF
C26600 OR2X1_LOC_377/A OR2X1_LOC_549/A 0.90fF
C26601 OR2X1_LOC_542/B OR2X1_LOC_254/A 0.02fF
C26602 OR2X1_LOC_427/A AND2X1_LOC_778/Y 0.07fF
C26603 GATE_366 OR2X1_LOC_428/A 0.27fF
C26604 AND2X1_LOC_786/a_36_24# OR2X1_LOC_36/Y 0.00fF
C26605 VDD OR2X1_LOC_837/A 0.21fF
C26606 OR2X1_LOC_231/B OR2X1_LOC_87/A 0.06fF
C26607 OR2X1_LOC_131/Y AND2X1_LOC_772/Y 0.07fF
C26608 OR2X1_LOC_756/B OR2X1_LOC_471/B 0.00fF
C26609 OR2X1_LOC_404/Y OR2X1_LOC_501/A 0.03fF
C26610 OR2X1_LOC_161/A OR2X1_LOC_307/A 0.02fF
C26611 OR2X1_LOC_458/B OR2X1_LOC_541/A 0.02fF
C26612 AND2X1_LOC_347/Y OR2X1_LOC_91/A 0.01fF
C26613 OR2X1_LOC_648/A OR2X1_LOC_61/a_8_216# 0.03fF
C26614 OR2X1_LOC_97/A OR2X1_LOC_155/A 0.03fF
C26615 OR2X1_LOC_8/Y AND2X1_LOC_839/a_36_24# 0.00fF
C26616 OR2X1_LOC_850/a_8_216# OR2X1_LOC_858/B -0.00fF
C26617 AND2X1_LOC_81/B AND2X1_LOC_65/A 0.03fF
C26618 AND2X1_LOC_541/Y AND2X1_LOC_113/Y 0.00fF
C26619 OR2X1_LOC_121/Y OR2X1_LOC_87/A 0.07fF
C26620 AND2X1_LOC_56/B OR2X1_LOC_344/A 0.04fF
C26621 AND2X1_LOC_828/a_8_24# OR2X1_LOC_44/Y 0.01fF
C26622 OR2X1_LOC_91/A AND2X1_LOC_857/Y 0.04fF
C26623 AND2X1_LOC_64/Y OR2X1_LOC_475/Y 0.02fF
C26624 AND2X1_LOC_392/a_8_24# OR2X1_LOC_517/A 0.01fF
C26625 OR2X1_LOC_821/a_8_216# OR2X1_LOC_43/A 0.06fF
C26626 OR2X1_LOC_668/a_36_216# OR2X1_LOC_66/A 0.03fF
C26627 OR2X1_LOC_750/A OR2X1_LOC_333/A 0.03fF
C26628 OR2X1_LOC_45/B AND2X1_LOC_512/a_8_24# 0.03fF
C26629 OR2X1_LOC_22/A INPUT_6 0.08fF
C26630 OR2X1_LOC_78/A OR2X1_LOC_475/B 0.26fF
C26631 OR2X1_LOC_312/Y OR2X1_LOC_428/A 0.09fF
C26632 OR2X1_LOC_426/B AND2X1_LOC_649/B 0.46fF
C26633 OR2X1_LOC_451/B AND2X1_LOC_430/B 0.00fF
C26634 OR2X1_LOC_421/A AND2X1_LOC_435/a_8_24# 0.01fF
C26635 AND2X1_LOC_125/a_8_24# OR2X1_LOC_363/A 0.23fF
C26636 OR2X1_LOC_12/Y AND2X1_LOC_637/Y 0.02fF
C26637 VDD OR2X1_LOC_796/a_8_216# 0.00fF
C26638 AND2X1_LOC_713/Y AND2X1_LOC_454/Y 0.00fF
C26639 OR2X1_LOC_203/Y OR2X1_LOC_549/A 0.68fF
C26640 OR2X1_LOC_448/a_36_216# OR2X1_LOC_78/A 0.03fF
C26641 OR2X1_LOC_45/B AND2X1_LOC_717/B 0.39fF
C26642 OR2X1_LOC_324/a_8_216# OR2X1_LOC_324/B 0.01fF
C26643 OR2X1_LOC_865/B OR2X1_LOC_244/Y 0.02fF
C26644 OR2X1_LOC_160/B OR2X1_LOC_499/a_8_216# 0.02fF
C26645 OR2X1_LOC_252/a_8_216# OR2X1_LOC_627/Y 0.01fF
C26646 AND2X1_LOC_719/Y AND2X1_LOC_286/Y 0.04fF
C26647 AND2X1_LOC_18/Y OR2X1_LOC_541/a_8_216# 0.01fF
C26648 AND2X1_LOC_279/a_36_24# OR2X1_LOC_366/Y 0.01fF
C26649 OR2X1_LOC_510/A AND2X1_LOC_81/B 0.01fF
C26650 VDD AND2X1_LOC_34/Y 0.24fF
C26651 OR2X1_LOC_620/B OR2X1_LOC_547/a_8_216# 0.47fF
C26652 AND2X1_LOC_535/Y AND2X1_LOC_319/A 0.02fF
C26653 AND2X1_LOC_147/Y AND2X1_LOC_213/B 0.00fF
C26654 AND2X1_LOC_843/a_8_24# AND2X1_LOC_286/a_8_24# 0.23fF
C26655 AND2X1_LOC_784/A OR2X1_LOC_309/a_8_216# 0.04fF
C26656 OR2X1_LOC_3/Y AND2X1_LOC_639/B 0.23fF
C26657 AND2X1_LOC_546/a_36_24# AND2X1_LOC_658/A 0.01fF
C26658 AND2X1_LOC_787/A OR2X1_LOC_70/Y 0.03fF
C26659 AND2X1_LOC_357/B OR2X1_LOC_6/A 0.02fF
C26660 OR2X1_LOC_425/a_8_216# OR2X1_LOC_426/A -0.00fF
C26661 AND2X1_LOC_136/a_8_24# AND2X1_LOC_44/Y 0.02fF
C26662 OR2X1_LOC_599/A AND2X1_LOC_713/Y 0.00fF
C26663 OR2X1_LOC_756/B OR2X1_LOC_788/a_36_216# 0.00fF
C26664 OR2X1_LOC_244/Y OR2X1_LOC_573/Y 0.01fF
C26665 AND2X1_LOC_186/a_8_24# AND2X1_LOC_188/a_8_24# 0.23fF
C26666 OR2X1_LOC_185/Y OR2X1_LOC_800/Y 0.01fF
C26667 OR2X1_LOC_40/Y AND2X1_LOC_806/A 0.05fF
C26668 OR2X1_LOC_680/A OR2X1_LOC_51/Y 0.54fF
C26669 OR2X1_LOC_160/A AND2X1_LOC_320/a_8_24# 0.15fF
C26670 OR2X1_LOC_176/a_8_216# OR2X1_LOC_417/Y 0.01fF
C26671 OR2X1_LOC_318/a_8_216# OR2X1_LOC_479/Y 0.01fF
C26672 OR2X1_LOC_526/Y OR2X1_LOC_36/Y 0.03fF
C26673 OR2X1_LOC_276/B AND2X1_LOC_36/Y 0.09fF
C26674 OR2X1_LOC_160/A OR2X1_LOC_660/Y 0.01fF
C26675 AND2X1_LOC_307/a_8_24# OR2X1_LOC_428/A 0.03fF
C26676 AND2X1_LOC_514/a_8_24# AND2X1_LOC_655/A 0.34fF
C26677 AND2X1_LOC_367/A OR2X1_LOC_18/Y 0.06fF
C26678 OR2X1_LOC_329/B OR2X1_LOC_316/Y 0.03fF
C26679 OR2X1_LOC_375/A OR2X1_LOC_78/B 0.81fF
C26680 AND2X1_LOC_56/a_8_24# AND2X1_LOC_763/B 0.09fF
C26681 OR2X1_LOC_799/A OR2X1_LOC_435/B 0.04fF
C26682 OR2X1_LOC_744/A AND2X1_LOC_572/A 0.18fF
C26683 VDD OR2X1_LOC_670/Y 0.12fF
C26684 AND2X1_LOC_719/Y OR2X1_LOC_280/Y 0.10fF
C26685 AND2X1_LOC_303/A AND2X1_LOC_219/Y -0.01fF
C26686 AND2X1_LOC_40/Y OR2X1_LOC_807/Y 0.18fF
C26687 OR2X1_LOC_667/a_8_216# OR2X1_LOC_51/Y 0.01fF
C26688 OR2X1_LOC_708/B OR2X1_LOC_66/A 0.01fF
C26689 OR2X1_LOC_703/B OR2X1_LOC_538/A 0.04fF
C26690 AND2X1_LOC_307/Y AND2X1_LOC_774/A 0.10fF
C26691 OR2X1_LOC_158/A OR2X1_LOC_279/Y 0.09fF
C26692 OR2X1_LOC_791/A OR2X1_LOC_555/B 0.80fF
C26693 AND2X1_LOC_554/B AND2X1_LOC_243/Y 0.03fF
C26694 OR2X1_LOC_631/a_8_216# OR2X1_LOC_575/A 0.41fF
C26695 OR2X1_LOC_47/Y AND2X1_LOC_439/a_8_24# 0.01fF
C26696 OR2X1_LOC_649/B AND2X1_LOC_92/Y 0.01fF
C26697 AND2X1_LOC_208/B AND2X1_LOC_34/Y 0.03fF
C26698 OR2X1_LOC_47/Y OR2X1_LOC_387/A 0.01fF
C26699 OR2X1_LOC_335/Y AND2X1_LOC_369/a_8_24# 0.23fF
C26700 AND2X1_LOC_303/a_8_24# OR2X1_LOC_6/A 0.02fF
C26701 OR2X1_LOC_318/Y OR2X1_LOC_185/A 7.27fF
C26702 INPUT_4 OR2X1_LOC_425/a_8_216# 0.00fF
C26703 OR2X1_LOC_62/B OR2X1_LOC_548/B 0.01fF
C26704 OR2X1_LOC_160/B OR2X1_LOC_675/a_8_216# 0.01fF
C26705 OR2X1_LOC_326/B OR2X1_LOC_739/A 0.03fF
C26706 OR2X1_LOC_375/A OR2X1_LOC_721/Y 0.12fF
C26707 OR2X1_LOC_743/A AND2X1_LOC_447/Y 0.02fF
C26708 OR2X1_LOC_656/Y OR2X1_LOC_87/Y 0.06fF
C26709 VDD OR2X1_LOC_48/Y 0.05fF
C26710 OR2X1_LOC_154/A AND2X1_LOC_65/a_36_24# 0.01fF
C26711 AND2X1_LOC_769/a_36_24# OR2X1_LOC_409/B 0.00fF
C26712 OR2X1_LOC_624/A OR2X1_LOC_231/A 0.06fF
C26713 OR2X1_LOC_147/A OR2X1_LOC_710/a_8_216# 0.48fF
C26714 AND2X1_LOC_743/a_8_24# OR2X1_LOC_446/Y 0.01fF
C26715 AND2X1_LOC_489/Y AND2X1_LOC_561/B 0.65fF
C26716 OR2X1_LOC_599/A OR2X1_LOC_441/Y 0.03fF
C26717 AND2X1_LOC_566/B AND2X1_LOC_514/Y 0.10fF
C26718 OR2X1_LOC_427/A AND2X1_LOC_624/A 0.06fF
C26719 AND2X1_LOC_516/a_36_24# OR2X1_LOC_715/A 0.00fF
C26720 OR2X1_LOC_485/A AND2X1_LOC_434/Y 0.24fF
C26721 AND2X1_LOC_744/a_8_24# OR2X1_LOC_155/A 0.01fF
C26722 OR2X1_LOC_502/A AND2X1_LOC_404/a_8_24# 0.06fF
C26723 OR2X1_LOC_158/A OR2X1_LOC_77/a_8_216# 0.02fF
C26724 OR2X1_LOC_672/a_8_216# OR2X1_LOC_46/A 0.01fF
C26725 OR2X1_LOC_3/Y OR2X1_LOC_744/A 0.67fF
C26726 AND2X1_LOC_711/A AND2X1_LOC_663/B 0.00fF
C26727 AND2X1_LOC_719/Y OR2X1_LOC_22/Y 0.17fF
C26728 OR2X1_LOC_529/a_8_216# AND2X1_LOC_113/Y 0.00fF
C26729 OR2X1_LOC_426/B AND2X1_LOC_729/B 0.03fF
C26730 AND2X1_LOC_31/Y OR2X1_LOC_771/B 0.13fF
C26731 OR2X1_LOC_329/B AND2X1_LOC_390/B 0.07fF
C26732 OR2X1_LOC_702/A INPUT_0 0.00fF
C26733 OR2X1_LOC_185/A OR2X1_LOC_805/A 0.03fF
C26734 OR2X1_LOC_532/B OR2X1_LOC_390/A 0.00fF
C26735 AND2X1_LOC_48/A OR2X1_LOC_641/A 0.20fF
C26736 OR2X1_LOC_494/a_8_216# OR2X1_LOC_7/A 0.03fF
C26737 VDD OR2X1_LOC_656/a_8_216# 0.21fF
C26738 OR2X1_LOC_62/B OR2X1_LOC_786/A 0.00fF
C26739 OR2X1_LOC_533/a_8_216# OR2X1_LOC_13/B 0.05fF
C26740 OR2X1_LOC_604/A OR2X1_LOC_295/Y 0.06fF
C26741 OR2X1_LOC_624/A OR2X1_LOC_130/A 0.10fF
C26742 AND2X1_LOC_35/Y OR2X1_LOC_18/Y 0.01fF
C26743 OR2X1_LOC_317/B OR2X1_LOC_704/a_8_216# 0.10fF
C26744 VDD OR2X1_LOC_520/B -0.00fF
C26745 AND2X1_LOC_508/A OR2X1_LOC_74/A 0.03fF
C26746 OR2X1_LOC_185/A AND2X1_LOC_153/a_36_24# 0.00fF
C26747 AND2X1_LOC_191/B OR2X1_LOC_64/Y 0.03fF
C26748 AND2X1_LOC_843/Y AND2X1_LOC_806/A 0.00fF
C26749 AND2X1_LOC_859/Y OR2X1_LOC_278/Y 0.17fF
C26750 AND2X1_LOC_660/A AND2X1_LOC_786/Y 0.07fF
C26751 AND2X1_LOC_59/Y OR2X1_LOC_219/a_8_216# 0.01fF
C26752 OR2X1_LOC_64/Y AND2X1_LOC_469/B 0.03fF
C26753 AND2X1_LOC_59/Y OR2X1_LOC_241/a_8_216# 0.01fF
C26754 AND2X1_LOC_47/Y AND2X1_LOC_295/a_36_24# 0.00fF
C26755 AND2X1_LOC_729/Y OR2X1_LOC_511/Y 0.03fF
C26756 OR2X1_LOC_43/A AND2X1_LOC_809/A 0.01fF
C26757 AND2X1_LOC_31/Y OR2X1_LOC_776/A 1.82fF
C26758 OR2X1_LOC_36/Y OR2X1_LOC_433/Y 0.03fF
C26759 AND2X1_LOC_848/Y AND2X1_LOC_859/a_8_24# 0.10fF
C26760 AND2X1_LOC_12/Y OR2X1_LOC_87/A 0.39fF
C26761 OR2X1_LOC_67/Y AND2X1_LOC_202/Y 0.00fF
C26762 AND2X1_LOC_730/a_8_24# AND2X1_LOC_192/Y 0.03fF
C26763 AND2X1_LOC_56/B OR2X1_LOC_203/a_36_216# 0.00fF
C26764 AND2X1_LOC_214/A OR2X1_LOC_52/Y 0.62fF
C26765 AND2X1_LOC_787/A OR2X1_LOC_437/Y 0.06fF
C26766 OR2X1_LOC_457/B OR2X1_LOC_553/A 0.01fF
C26767 VDD OR2X1_LOC_818/a_8_216# 0.21fF
C26768 OR2X1_LOC_599/A AND2X1_LOC_436/B 0.02fF
C26769 OR2X1_LOC_424/a_36_216# OR2X1_LOC_44/Y 0.01fF
C26770 OR2X1_LOC_476/B INPUT_0 0.08fF
C26771 OR2X1_LOC_479/Y OR2X1_LOC_478/a_8_216# 0.00fF
C26772 AND2X1_LOC_479/Y AND2X1_LOC_476/Y 0.00fF
C26773 AND2X1_LOC_535/Y AND2X1_LOC_170/B 0.35fF
C26774 AND2X1_LOC_47/Y INPUT_2 0.06fF
C26775 OR2X1_LOC_13/B OR2X1_LOC_142/a_8_216# 0.02fF
C26776 AND2X1_LOC_486/Y AND2X1_LOC_578/A 0.07fF
C26777 OR2X1_LOC_185/Y OR2X1_LOC_800/A 0.01fF
C26778 OR2X1_LOC_628/Y AND2X1_LOC_663/A 0.10fF
C26779 OR2X1_LOC_26/Y OR2X1_LOC_69/A 0.03fF
C26780 AND2X1_LOC_542/a_8_24# OR2X1_LOC_47/Y 0.01fF
C26781 OR2X1_LOC_74/A OR2X1_LOC_48/B 0.07fF
C26782 VDD AND2X1_LOC_656/Y 0.40fF
C26783 OR2X1_LOC_32/B OR2X1_LOC_585/A 0.07fF
C26784 OR2X1_LOC_479/Y OR2X1_LOC_794/A 0.01fF
C26785 AND2X1_LOC_95/Y OR2X1_LOC_557/A 0.02fF
C26786 VDD OR2X1_LOC_639/a_8_216# 0.00fF
C26787 AND2X1_LOC_59/Y AND2X1_LOC_81/a_36_24# 0.00fF
C26788 OR2X1_LOC_9/Y OR2X1_LOC_47/Y 0.07fF
C26789 OR2X1_LOC_18/Y OR2X1_LOC_74/A 0.19fF
C26790 AND2X1_LOC_191/B OR2X1_LOC_417/A 1.00fF
C26791 OR2X1_LOC_11/Y AND2X1_LOC_638/a_8_24# 0.01fF
C26792 AND2X1_LOC_657/A AND2X1_LOC_772/Y 0.05fF
C26793 OR2X1_LOC_675/A OR2X1_LOC_737/A 0.01fF
C26794 AND2X1_LOC_120/a_8_24# AND2X1_LOC_850/a_8_24# 0.23fF
C26795 AND2X1_LOC_839/B OR2X1_LOC_6/A 0.00fF
C26796 OR2X1_LOC_743/A AND2X1_LOC_448/Y 0.01fF
C26797 OR2X1_LOC_86/Y AND2X1_LOC_100/a_8_24# 0.23fF
C26798 AND2X1_LOC_72/B AND2X1_LOC_295/a_8_24# 0.01fF
C26799 OR2X1_LOC_643/a_8_216# OR2X1_LOC_222/A 0.01fF
C26800 OR2X1_LOC_329/B AND2X1_LOC_863/Y 0.19fF
C26801 OR2X1_LOC_809/B OR2X1_LOC_436/Y 0.00fF
C26802 OR2X1_LOC_756/B D_INPUT_0 0.14fF
C26803 AND2X1_LOC_675/A OR2X1_LOC_59/Y 0.19fF
C26804 INPUT_0 OR2X1_LOC_111/Y 0.03fF
C26805 OR2X1_LOC_774/Y D_GATE_865 0.01fF
C26806 OR2X1_LOC_264/a_8_216# AND2X1_LOC_3/Y 0.01fF
C26807 OR2X1_LOC_605/B OR2X1_LOC_375/A 0.01fF
C26808 OR2X1_LOC_675/a_8_216# OR2X1_LOC_553/A 0.04fF
C26809 OR2X1_LOC_615/Y AND2X1_LOC_285/Y 0.02fF
C26810 AND2X1_LOC_811/a_36_24# OR2X1_LOC_74/A 0.02fF
C26811 OR2X1_LOC_7/A AND2X1_LOC_806/A 0.03fF
C26812 AND2X1_LOC_40/Y AND2X1_LOC_600/a_8_24# 0.04fF
C26813 AND2X1_LOC_59/Y AND2X1_LOC_666/a_8_24# 0.01fF
C26814 OR2X1_LOC_18/Y OR2X1_LOC_762/a_36_216# 0.02fF
C26815 OR2X1_LOC_844/Y OR2X1_LOC_571/B 0.01fF
C26816 AND2X1_LOC_660/A AND2X1_LOC_218/Y 0.09fF
C26817 OR2X1_LOC_516/Y OR2X1_LOC_142/Y 9.94fF
C26818 OR2X1_LOC_786/a_8_216# OR2X1_LOC_598/A 0.01fF
C26819 VDD OR2X1_LOC_770/Y -0.00fF
C26820 AND2X1_LOC_753/a_8_24# AND2X1_LOC_48/A 0.01fF
C26821 AND2X1_LOC_56/B AND2X1_LOC_13/a_8_24# 0.02fF
C26822 OR2X1_LOC_379/Y AND2X1_LOC_48/A 0.01fF
C26823 AND2X1_LOC_181/Y AND2X1_LOC_222/Y 0.02fF
C26824 OR2X1_LOC_348/Y OR2X1_LOC_366/a_8_216# 0.03fF
C26825 AND2X1_LOC_41/A OR2X1_LOC_506/B 0.01fF
C26826 OR2X1_LOC_233/a_8_216# OR2X1_LOC_585/A 0.01fF
C26827 OR2X1_LOC_287/B AND2X1_LOC_86/B 0.03fF
C26828 OR2X1_LOC_817/Y OR2X1_LOC_820/B 0.00fF
C26829 OR2X1_LOC_624/A OR2X1_LOC_62/B 0.05fF
C26830 OR2X1_LOC_244/Y OR2X1_LOC_493/Y 0.03fF
C26831 VDD AND2X1_LOC_679/a_8_24# 0.00fF
C26832 OR2X1_LOC_22/Y AND2X1_LOC_655/A 0.03fF
C26833 AND2X1_LOC_70/Y OR2X1_LOC_451/B 0.01fF
C26834 AND2X1_LOC_753/B OR2X1_LOC_651/A 0.31fF
C26835 OR2X1_LOC_160/A OR2X1_LOC_835/Y 0.00fF
C26836 OR2X1_LOC_508/A OR2X1_LOC_506/B 1.00fF
C26837 AND2X1_LOC_391/a_36_24# D_INPUT_3 0.01fF
C26838 AND2X1_LOC_12/Y OR2X1_LOC_706/B 0.01fF
C26839 AND2X1_LOC_535/Y OR2X1_LOC_331/Y 0.03fF
C26840 OR2X1_LOC_161/B OR2X1_LOC_446/B 0.07fF
C26841 OR2X1_LOC_3/Y OR2X1_LOC_282/a_8_216# 0.01fF
C26842 AND2X1_LOC_48/A OR2X1_LOC_194/Y 0.03fF
C26843 AND2X1_LOC_851/A AND2X1_LOC_851/B 0.09fF
C26844 OR2X1_LOC_497/Y AND2X1_LOC_849/A 0.01fF
C26845 OR2X1_LOC_103/a_36_216# AND2X1_LOC_227/Y 0.00fF
C26846 OR2X1_LOC_604/A AND2X1_LOC_563/Y 0.03fF
C26847 OR2X1_LOC_428/A OR2X1_LOC_13/B 0.53fF
C26848 OR2X1_LOC_161/B OR2X1_LOC_303/B 0.07fF
C26849 VDD AND2X1_LOC_779/Y 0.25fF
C26850 OR2X1_LOC_791/B OR2X1_LOC_288/A 0.01fF
C26851 OR2X1_LOC_64/Y AND2X1_LOC_638/a_8_24# 0.00fF
C26852 OR2X1_LOC_160/B OR2X1_LOC_750/Y 0.07fF
C26853 AND2X1_LOC_47/Y OR2X1_LOC_739/A 0.17fF
C26854 OR2X1_LOC_19/B AND2X1_LOC_412/a_8_24# 0.07fF
C26855 OR2X1_LOC_605/A OR2X1_LOC_605/a_8_216# 0.03fF
C26856 OR2X1_LOC_481/Y AND2X1_LOC_345/Y 0.82fF
C26857 OR2X1_LOC_743/A AND2X1_LOC_729/B 0.62fF
C26858 OR2X1_LOC_18/Y AND2X1_LOC_660/a_36_24# 0.00fF
C26859 OR2X1_LOC_412/a_8_216# OR2X1_LOC_44/Y 0.06fF
C26860 OR2X1_LOC_160/A OR2X1_LOC_436/Y 0.03fF
C26861 OR2X1_LOC_13/B OR2X1_LOC_595/A 0.24fF
C26862 OR2X1_LOC_373/a_8_216# OR2X1_LOC_142/Y 0.06fF
C26863 OR2X1_LOC_502/A AND2X1_LOC_8/a_36_24# 0.01fF
C26864 OR2X1_LOC_526/Y OR2X1_LOC_526/a_8_216# 0.01fF
C26865 OR2X1_LOC_127/Y D_INPUT_3 0.01fF
C26866 AND2X1_LOC_465/Y OR2X1_LOC_238/Y 0.02fF
C26867 AND2X1_LOC_51/Y OR2X1_LOC_35/B 0.03fF
C26868 AND2X1_LOC_26/a_8_24# AND2X1_LOC_47/Y 0.01fF
C26869 OR2X1_LOC_744/A AND2X1_LOC_772/a_8_24# 0.01fF
C26870 OR2X1_LOC_45/B OR2X1_LOC_395/Y 0.14fF
C26871 OR2X1_LOC_36/Y AND2X1_LOC_810/Y 0.15fF
C26872 OR2X1_LOC_475/Y OR2X1_LOC_206/A 0.23fF
C26873 AND2X1_LOC_47/Y OR2X1_LOC_269/B 1.91fF
C26874 OR2X1_LOC_709/A AND2X1_LOC_36/Y 0.07fF
C26875 OR2X1_LOC_165/Y AND2X1_LOC_222/Y 0.01fF
C26876 AND2X1_LOC_640/Y INPUT_1 0.02fF
C26877 OR2X1_LOC_416/A OR2X1_LOC_52/B 0.25fF
C26878 OR2X1_LOC_47/Y OR2X1_LOC_96/B 0.03fF
C26879 D_INPUT_3 AND2X1_LOC_836/a_8_24# 0.01fF
C26880 OR2X1_LOC_635/A AND2X1_LOC_430/B 0.00fF
C26881 OR2X1_LOC_95/Y AND2X1_LOC_458/a_36_24# 0.00fF
C26882 OR2X1_LOC_308/A AND2X1_LOC_22/Y 0.00fF
C26883 OR2X1_LOC_246/Y AND2X1_LOC_721/A 0.02fF
C26884 OR2X1_LOC_18/Y AND2X1_LOC_647/Y 0.00fF
C26885 OR2X1_LOC_240/a_8_216# OR2X1_LOC_598/A 0.02fF
C26886 OR2X1_LOC_811/A OR2X1_LOC_736/a_8_216# 0.02fF
C26887 OR2X1_LOC_3/Y OR2X1_LOC_31/Y 0.18fF
C26888 OR2X1_LOC_529/Y AND2X1_LOC_866/A 0.03fF
C26889 OR2X1_LOC_47/Y AND2X1_LOC_852/Y 0.03fF
C26890 OR2X1_LOC_472/B OR2X1_LOC_19/B 0.04fF
C26891 OR2X1_LOC_405/A OR2X1_LOC_728/B 0.00fF
C26892 AND2X1_LOC_69/a_8_24# AND2X1_LOC_51/Y 0.01fF
C26893 AND2X1_LOC_391/Y OR2X1_LOC_437/A 0.07fF
C26894 AND2X1_LOC_858/B OR2X1_LOC_437/A 0.07fF
C26895 OR2X1_LOC_91/A OR2X1_LOC_437/A 0.43fF
C26896 OR2X1_LOC_83/Y OR2X1_LOC_47/Y 0.01fF
C26897 AND2X1_LOC_31/Y OR2X1_LOC_733/a_8_216# 0.01fF
C26898 OR2X1_LOC_485/A AND2X1_LOC_851/B 0.01fF
C26899 AND2X1_LOC_11/Y AND2X1_LOC_31/Y 0.05fF
C26900 AND2X1_LOC_18/Y OR2X1_LOC_523/a_8_216# 0.05fF
C26901 OR2X1_LOC_114/B OR2X1_LOC_844/B 0.92fF
C26902 AND2X1_LOC_92/Y OR2X1_LOC_777/B 0.10fF
C26903 OR2X1_LOC_70/Y AND2X1_LOC_675/A 0.14fF
C26904 OR2X1_LOC_62/B OR2X1_LOC_54/Y 0.13fF
C26905 AND2X1_LOC_684/a_36_24# AND2X1_LOC_3/Y 0.00fF
C26906 INPUT_1 OR2X1_LOC_416/Y 0.07fF
C26907 AND2X1_LOC_64/Y OR2X1_LOC_356/A 0.27fF
C26908 OR2X1_LOC_6/A AND2X1_LOC_228/a_8_24# 0.02fF
C26909 OR2X1_LOC_111/Y OR2X1_LOC_64/Y 0.15fF
C26910 OR2X1_LOC_656/B OR2X1_LOC_560/A 0.00fF
C26911 OR2X1_LOC_92/Y OR2X1_LOC_71/A -0.00fF
C26912 AND2X1_LOC_70/Y AND2X1_LOC_36/Y 2.05fF
C26913 OR2X1_LOC_478/Y OR2X1_LOC_161/B 0.01fF
C26914 OR2X1_LOC_151/A OR2X1_LOC_115/B 0.20fF
C26915 OR2X1_LOC_631/B OR2X1_LOC_247/Y 0.03fF
C26916 OR2X1_LOC_532/B OR2X1_LOC_750/A 0.00fF
C26917 OR2X1_LOC_632/Y OR2X1_LOC_523/A 0.05fF
C26918 OR2X1_LOC_74/A AND2X1_LOC_620/Y 0.03fF
C26919 OR2X1_LOC_852/A OR2X1_LOC_19/B 0.01fF
C26920 OR2X1_LOC_269/B OR2X1_LOC_598/A 0.03fF
C26921 AND2X1_LOC_17/Y OR2X1_LOC_451/B 0.46fF
C26922 OR2X1_LOC_105/Y OR2X1_LOC_580/A 0.01fF
C26923 OR2X1_LOC_11/Y OR2X1_LOC_588/a_8_216# 0.01fF
C26924 OR2X1_LOC_756/B OR2X1_LOC_339/A 0.24fF
C26925 OR2X1_LOC_696/a_8_216# OR2X1_LOC_511/a_8_216# 0.47fF
C26926 AND2X1_LOC_462/Y OR2X1_LOC_46/A 0.02fF
C26927 OR2X1_LOC_687/B AND2X1_LOC_430/B 0.01fF
C26928 VDD AND2X1_LOC_772/Y 0.75fF
C26929 OR2X1_LOC_696/A AND2X1_LOC_637/a_8_24# 0.02fF
C26930 OR2X1_LOC_692/Y OR2X1_LOC_693/Y 0.21fF
C26931 OR2X1_LOC_74/A AND2X1_LOC_215/A 0.08fF
C26932 OR2X1_LOC_111/Y OR2X1_LOC_417/A 0.03fF
C26933 OR2X1_LOC_147/B OR2X1_LOC_182/a_8_216# 0.06fF
C26934 OR2X1_LOC_161/B OR2X1_LOC_719/B 0.01fF
C26935 AND2X1_LOC_227/Y OR2X1_LOC_71/Y 0.89fF
C26936 AND2X1_LOC_573/A OR2X1_LOC_437/A 0.07fF
C26937 AND2X1_LOC_544/Y AND2X1_LOC_657/Y 0.03fF
C26938 OR2X1_LOC_719/A OR2X1_LOC_241/B 0.41fF
C26939 OR2X1_LOC_804/A AND2X1_LOC_51/Y 0.07fF
C26940 OR2X1_LOC_467/B OR2X1_LOC_160/Y 0.03fF
C26941 OR2X1_LOC_814/A AND2X1_LOC_250/a_8_24# 0.01fF
C26942 OR2X1_LOC_404/Y AND2X1_LOC_72/B -0.02fF
C26943 D_INPUT_2 AND2X1_LOC_28/a_8_24# 0.01fF
C26944 AND2X1_LOC_51/Y AND2X1_LOC_428/a_8_24# 0.01fF
C26945 OR2X1_LOC_831/B AND2X1_LOC_92/Y 5.64fF
C26946 OR2X1_LOC_576/A AND2X1_LOC_18/Y 0.07fF
C26947 OR2X1_LOC_46/A D_INPUT_1 0.18fF
C26948 OR2X1_LOC_49/A OR2X1_LOC_604/A 0.09fF
C26949 AND2X1_LOC_348/Y OR2X1_LOC_384/Y 0.01fF
C26950 OR2X1_LOC_156/B VDD -0.00fF
C26951 OR2X1_LOC_175/Y OR2X1_LOC_78/A 0.07fF
C26952 AND2X1_LOC_570/Y OR2X1_LOC_816/A 0.03fF
C26953 OR2X1_LOC_49/A OR2X1_LOC_66/A 0.05fF
C26954 OR2X1_LOC_22/Y OR2X1_LOC_599/Y 0.03fF
C26955 OR2X1_LOC_542/B OR2X1_LOC_161/B 0.03fF
C26956 OR2X1_LOC_62/B OR2X1_LOC_84/Y 0.01fF
C26957 OR2X1_LOC_604/A OR2X1_LOC_381/a_36_216# 0.01fF
C26958 OR2X1_LOC_421/A OR2X1_LOC_158/A 2.52fF
C26959 OR2X1_LOC_548/A VDD -0.00fF
C26960 AND2X1_LOC_362/B AND2X1_LOC_243/Y 0.37fF
C26961 OR2X1_LOC_223/A OR2X1_LOC_440/A 0.03fF
C26962 VDD OR2X1_LOC_486/Y 0.56fF
C26963 OR2X1_LOC_669/Y OR2X1_LOC_437/A 0.07fF
C26964 OR2X1_LOC_46/a_8_216# OR2X1_LOC_171/Y 0.06fF
C26965 OR2X1_LOC_6/B OR2X1_LOC_40/Y 0.06fF
C26966 OR2X1_LOC_276/B OR2X1_LOC_269/Y 0.02fF
C26967 OR2X1_LOC_596/A OR2X1_LOC_66/A 0.03fF
C26968 AND2X1_LOC_92/Y OR2X1_LOC_344/A 0.01fF
C26969 OR2X1_LOC_437/Y AND2X1_LOC_675/A 0.19fF
C26970 OR2X1_LOC_78/A OR2X1_LOC_713/A 0.07fF
C26971 OR2X1_LOC_593/a_8_216# OR2X1_LOC_593/B 0.06fF
C26972 OR2X1_LOC_589/A OR2X1_LOC_56/A 0.12fF
C26973 OR2X1_LOC_235/B OR2X1_LOC_16/A 0.65fF
C26974 OR2X1_LOC_604/A OR2X1_LOC_526/Y 0.01fF
C26975 OR2X1_LOC_78/B OR2X1_LOC_549/A 0.37fF
C26976 OR2X1_LOC_36/Y AND2X1_LOC_204/a_8_24# 0.07fF
C26977 OR2X1_LOC_756/B AND2X1_LOC_438/a_8_24# 0.01fF
C26978 AND2X1_LOC_539/Y AND2X1_LOC_354/Y 0.00fF
C26979 OR2X1_LOC_161/A OR2X1_LOC_186/a_36_216# 0.02fF
C26980 AND2X1_LOC_392/A AND2X1_LOC_326/B 0.03fF
C26981 AND2X1_LOC_810/Y OR2X1_LOC_419/Y 0.10fF
C26982 OR2X1_LOC_703/B OR2X1_LOC_356/B 0.00fF
C26983 AND2X1_LOC_95/Y OR2X1_LOC_703/a_8_216# 0.01fF
C26984 OR2X1_LOC_633/B OR2X1_LOC_771/B 0.05fF
C26985 AND2X1_LOC_17/Y AND2X1_LOC_36/Y 0.01fF
C26986 AND2X1_LOC_64/Y AND2X1_LOC_43/B 0.26fF
C26987 OR2X1_LOC_20/Y AND2X1_LOC_33/a_8_24# 0.23fF
C26988 OR2X1_LOC_47/Y AND2X1_LOC_647/B 0.14fF
C26989 AND2X1_LOC_81/B OR2X1_LOC_502/a_36_216# 0.00fF
C26990 OR2X1_LOC_64/Y OR2X1_LOC_164/a_8_216# 0.00fF
C26991 OR2X1_LOC_18/Y AND2X1_LOC_773/a_36_24# 0.00fF
C26992 AND2X1_LOC_392/A AND2X1_LOC_337/a_36_24# 0.00fF
C26993 AND2X1_LOC_642/Y AND2X1_LOC_786/Y 0.04fF
C26994 AND2X1_LOC_715/A AND2X1_LOC_112/a_36_24# 0.00fF
C26995 VDD AND2X1_LOC_160/Y 0.21fF
C26996 AND2X1_LOC_483/Y OR2X1_LOC_615/Y 0.38fF
C26997 OR2X1_LOC_479/Y OR2X1_LOC_716/a_36_216# 0.01fF
C26998 AND2X1_LOC_266/a_8_24# OR2X1_LOC_595/A 0.01fF
C26999 OR2X1_LOC_158/A AND2X1_LOC_456/B 0.04fF
C27000 OR2X1_LOC_448/B OR2X1_LOC_713/A 0.01fF
C27001 INPUT_1 OR2X1_LOC_80/A 1.42fF
C27002 AND2X1_LOC_549/Y AND2X1_LOC_549/a_8_24# 0.00fF
C27003 OR2X1_LOC_776/Y OR2X1_LOC_795/B 0.02fF
C27004 OR2X1_LOC_721/Y OR2X1_LOC_549/A 0.10fF
C27005 AND2X1_LOC_337/a_8_24# OR2X1_LOC_56/A 0.04fF
C27006 OR2X1_LOC_757/A OR2X1_LOC_815/a_36_216# 0.01fF
C27007 OR2X1_LOC_151/A OR2X1_LOC_840/A 0.10fF
C27008 AND2X1_LOC_508/B AND2X1_LOC_663/A 0.05fF
C27009 OR2X1_LOC_40/Y OR2X1_LOC_292/a_36_216# 0.03fF
C27010 OR2X1_LOC_427/A AND2X1_LOC_774/A 0.48fF
C27011 AND2X1_LOC_753/a_8_24# OR2X1_LOC_207/B 0.01fF
C27012 OR2X1_LOC_220/B OR2X1_LOC_547/a_8_216# 0.01fF
C27013 OR2X1_LOC_62/a_8_216# OR2X1_LOC_71/A 0.01fF
C27014 OR2X1_LOC_40/Y AND2X1_LOC_335/a_8_24# 0.02fF
C27015 OR2X1_LOC_631/a_8_216# OR2X1_LOC_161/B 0.02fF
C27016 OR2X1_LOC_510/Y OR2X1_LOC_267/Y 0.00fF
C27017 AND2X1_LOC_810/A OR2X1_LOC_48/B 0.57fF
C27018 OR2X1_LOC_600/A OR2X1_LOC_820/A 0.01fF
C27019 OR2X1_LOC_109/a_8_216# OR2X1_LOC_373/Y 0.01fF
C27020 AND2X1_LOC_715/A OR2X1_LOC_91/A 0.07fF
C27021 AND2X1_LOC_41/A AND2X1_LOC_18/Y 3.61fF
C27022 AND2X1_LOC_658/A AND2X1_LOC_443/Y 0.09fF
C27023 AND2X1_LOC_736/Y AND2X1_LOC_476/Y 0.07fF
C27024 OR2X1_LOC_40/Y OR2X1_LOC_441/Y 0.50fF
C27025 AND2X1_LOC_773/Y OR2X1_LOC_595/a_8_216# 0.06fF
C27026 OR2X1_LOC_185/A OR2X1_LOC_580/B 0.03fF
C27027 AND2X1_LOC_810/Y OR2X1_LOC_152/A 0.32fF
C27028 OR2X1_LOC_186/Y OR2X1_LOC_405/A 0.49fF
C27029 OR2X1_LOC_391/B OR2X1_LOC_773/Y 0.13fF
C27030 OR2X1_LOC_227/Y OR2X1_LOC_641/B 0.01fF
C27031 OR2X1_LOC_56/A OR2X1_LOC_297/A 0.01fF
C27032 AND2X1_LOC_675/Y AND2X1_LOC_188/a_36_24# 0.00fF
C27033 OR2X1_LOC_242/a_8_216# OR2X1_LOC_78/A 0.03fF
C27034 AND2X1_LOC_710/Y OR2X1_LOC_297/A 0.09fF
C27035 AND2X1_LOC_500/Y AND2X1_LOC_506/a_8_24# 0.01fF
C27036 AND2X1_LOC_851/a_8_24# AND2X1_LOC_858/B 0.01fF
C27037 AND2X1_LOC_392/A AND2X1_LOC_276/a_8_24# 0.07fF
C27038 OR2X1_LOC_329/B OR2X1_LOC_744/A 0.57fF
C27039 AND2X1_LOC_563/A OR2X1_LOC_103/Y 0.01fF
C27040 OR2X1_LOC_426/A OR2X1_LOC_582/a_8_216# 0.01fF
C27041 OR2X1_LOC_675/Y OR2X1_LOC_241/B 0.01fF
C27042 AND2X1_LOC_12/Y OR2X1_LOC_840/a_8_216# 0.01fF
C27043 OR2X1_LOC_523/B OR2X1_LOC_161/A 0.01fF
C27044 OR2X1_LOC_814/A OR2X1_LOC_349/B 0.02fF
C27045 OR2X1_LOC_97/A OR2X1_LOC_97/B 0.00fF
C27046 OR2X1_LOC_207/B OR2X1_LOC_194/Y 0.03fF
C27047 OR2X1_LOC_175/Y OR2X1_LOC_155/A 0.07fF
C27048 AND2X1_LOC_319/A OR2X1_LOC_16/A 0.05fF
C27049 OR2X1_LOC_58/Y OR2X1_LOC_837/B 0.03fF
C27050 OR2X1_LOC_635/A AND2X1_LOC_70/Y 0.00fF
C27051 OR2X1_LOC_185/Y AND2X1_LOC_522/a_36_24# 0.06fF
C27052 AND2X1_LOC_56/B OR2X1_LOC_161/B 0.27fF
C27053 OR2X1_LOC_797/B OR2X1_LOC_161/A 0.01fF
C27054 OR2X1_LOC_375/A OR2X1_LOC_549/A 0.25fF
C27055 OR2X1_LOC_604/A AND2X1_LOC_805/Y 0.02fF
C27056 OR2X1_LOC_659/B OR2X1_LOC_161/B 0.00fF
C27057 AND2X1_LOC_866/B OR2X1_LOC_56/A 0.10fF
C27058 OR2X1_LOC_335/Y OR2X1_LOC_756/B 0.02fF
C27059 OR2X1_LOC_519/Y OR2X1_LOC_40/Y 0.01fF
C27060 OR2X1_LOC_154/A OR2X1_LOC_857/B 0.09fF
C27061 OR2X1_LOC_354/A OR2X1_LOC_78/B 0.07fF
C27062 AND2X1_LOC_719/Y OR2X1_LOC_39/A 0.10fF
C27063 OR2X1_LOC_443/a_8_216# OR2X1_LOC_181/Y 0.18fF
C27064 OR2X1_LOC_589/A AND2X1_LOC_87/a_8_24# 0.01fF
C27065 AND2X1_LOC_564/B OR2X1_LOC_371/Y 0.08fF
C27066 AND2X1_LOC_40/Y AND2X1_LOC_616/a_36_24# 0.00fF
C27067 OR2X1_LOC_92/Y OR2X1_LOC_59/Y 0.08fF
C27068 OR2X1_LOC_18/Y AND2X1_LOC_860/A 0.35fF
C27069 AND2X1_LOC_8/Y OR2X1_LOC_161/B 0.71fF
C27070 OR2X1_LOC_66/a_36_216# OR2X1_LOC_560/A 0.00fF
C27071 AND2X1_LOC_712/a_36_24# OR2X1_LOC_52/B 0.01fF
C27072 OR2X1_LOC_18/Y OR2X1_LOC_626/Y 0.12fF
C27073 OR2X1_LOC_600/A AND2X1_LOC_621/Y 0.03fF
C27074 OR2X1_LOC_702/A AND2X1_LOC_7/B 0.01fF
C27075 OR2X1_LOC_160/A OR2X1_LOC_160/B 1.83fF
C27076 OR2X1_LOC_629/Y OR2X1_LOC_78/A 0.01fF
C27077 AND2X1_LOC_714/B OR2X1_LOC_36/Y 0.00fF
C27078 AND2X1_LOC_473/a_8_24# AND2X1_LOC_473/Y 0.02fF
C27079 OR2X1_LOC_791/A OR2X1_LOC_756/B 0.12fF
C27080 OR2X1_LOC_684/a_8_216# AND2X1_LOC_452/Y 0.01fF
C27081 AND2X1_LOC_586/a_8_24# AND2X1_LOC_70/Y 0.14fF
C27082 OR2X1_LOC_339/a_36_216# AND2X1_LOC_95/Y 0.00fF
C27083 AND2X1_LOC_550/A AND2X1_LOC_657/Y 0.03fF
C27084 AND2X1_LOC_840/B AND2X1_LOC_477/Y 0.10fF
C27085 OR2X1_LOC_346/B AND2X1_LOC_295/a_8_24# 0.20fF
C27086 AND2X1_LOC_40/Y OR2X1_LOC_756/B 0.76fF
C27087 AND2X1_LOC_720/Y AND2X1_LOC_456/B 0.01fF
C27088 OR2X1_LOC_155/A OR2X1_LOC_713/A 0.07fF
C27089 AND2X1_LOC_593/Y AND2X1_LOC_436/Y 0.02fF
C27090 AND2X1_LOC_231/Y AND2X1_LOC_641/Y 0.07fF
C27091 AND2X1_LOC_721/Y OR2X1_LOC_279/Y 0.05fF
C27092 OR2X1_LOC_87/A OR2X1_LOC_182/B 0.91fF
C27093 AND2X1_LOC_729/Y OR2X1_LOC_600/a_8_216# 0.04fF
C27094 AND2X1_LOC_80/a_8_24# VDD -0.00fF
C27095 AND2X1_LOC_862/Y AND2X1_LOC_865/a_8_24# 0.01fF
C27096 AND2X1_LOC_64/Y AND2X1_LOC_698/a_8_24# 0.04fF
C27097 OR2X1_LOC_188/Y OR2X1_LOC_719/A 0.31fF
C27098 AND2X1_LOC_550/A AND2X1_LOC_469/B 0.03fF
C27099 INPUT_4 OR2X1_LOC_582/a_8_216# 0.01fF
C27100 OR2X1_LOC_325/a_8_216# OR2X1_LOC_703/A 0.01fF
C27101 OR2X1_LOC_768/A AND2X1_LOC_95/Y 0.10fF
C27102 OR2X1_LOC_575/a_8_216# OR2X1_LOC_66/A 0.02fF
C27103 AND2X1_LOC_340/Y OR2X1_LOC_74/A 0.07fF
C27104 AND2X1_LOC_3/Y OR2X1_LOC_294/Y 0.35fF
C27105 OR2X1_LOC_185/Y AND2X1_LOC_110/Y 0.02fF
C27106 AND2X1_LOC_554/B OR2X1_LOC_12/Y 0.05fF
C27107 AND2X1_LOC_570/Y AND2X1_LOC_807/Y 0.03fF
C27108 AND2X1_LOC_97/a_8_24# AND2X1_LOC_474/A 0.01fF
C27109 AND2X1_LOC_866/A AND2X1_LOC_791/a_8_24# 0.02fF
C27110 OR2X1_LOC_680/Y OR2X1_LOC_12/Y 0.00fF
C27111 OR2X1_LOC_40/Y OR2X1_LOC_235/Y 0.02fF
C27112 OR2X1_LOC_123/a_36_216# OR2X1_LOC_375/A 0.00fF
C27113 OR2X1_LOC_65/B OR2X1_LOC_59/Y 0.03fF
C27114 OR2X1_LOC_158/A AND2X1_LOC_717/B 0.19fF
C27115 OR2X1_LOC_744/A AND2X1_LOC_113/Y 0.01fF
C27116 OR2X1_LOC_631/B AND2X1_LOC_18/Y 0.03fF
C27117 OR2X1_LOC_476/B AND2X1_LOC_7/B 0.14fF
C27118 OR2X1_LOC_52/a_8_216# OR2X1_LOC_16/A 0.01fF
C27119 OR2X1_LOC_620/Y AND2X1_LOC_167/a_36_24# 0.01fF
C27120 OR2X1_LOC_87/B OR2X1_LOC_66/A 0.02fF
C27121 OR2X1_LOC_494/Y OR2X1_LOC_44/Y 0.06fF
C27122 AND2X1_LOC_95/Y AND2X1_LOC_71/a_8_24# 0.01fF
C27123 AND2X1_LOC_363/Y OR2X1_LOC_44/Y 0.03fF
C27124 VDD AND2X1_LOC_580/B 0.61fF
C27125 OR2X1_LOC_757/A OR2X1_LOC_680/A 0.03fF
C27126 OR2X1_LOC_756/B OR2X1_LOC_471/a_8_216# 0.22fF
C27127 AND2X1_LOC_768/a_8_24# AND2X1_LOC_560/B 0.02fF
C27128 OR2X1_LOC_650/Y AND2X1_LOC_7/B 0.03fF
C27129 OR2X1_LOC_805/A OR2X1_LOC_778/a_36_216# 0.00fF
C27130 OR2X1_LOC_624/A OR2X1_LOC_659/A 0.21fF
C27131 OR2X1_LOC_756/B OR2X1_LOC_537/A 0.00fF
C27132 AND2X1_LOC_713/Y OR2X1_LOC_7/A 0.01fF
C27133 AND2X1_LOC_3/Y OR2X1_LOC_641/A 0.04fF
C27134 OR2X1_LOC_462/B OR2X1_LOC_520/a_36_216# 0.00fF
C27135 OR2X1_LOC_859/A OR2X1_LOC_392/B 0.06fF
C27136 OR2X1_LOC_856/B OR2X1_LOC_175/B 0.02fF
C27137 OR2X1_LOC_40/Y OR2X1_LOC_529/Y 0.00fF
C27138 OR2X1_LOC_604/A AND2X1_LOC_259/Y 0.04fF
C27139 OR2X1_LOC_7/A AND2X1_LOC_448/a_36_24# 0.01fF
C27140 AND2X1_LOC_738/B OR2X1_LOC_43/A 0.01fF
C27141 AND2X1_LOC_141/A OR2X1_LOC_118/Y 0.00fF
C27142 OR2X1_LOC_43/A OR2X1_LOC_56/A 2.31fF
C27143 OR2X1_LOC_329/B AND2X1_LOC_840/B 0.04fF
C27144 OR2X1_LOC_256/A AND2X1_LOC_772/Y 0.02fF
C27145 OR2X1_LOC_426/Y AND2X1_LOC_450/a_8_24# 0.23fF
C27146 AND2X1_LOC_374/a_8_24# OR2X1_LOC_109/Y 0.02fF
C27147 AND2X1_LOC_94/Y OR2X1_LOC_82/a_8_216# 0.13fF
C27148 OR2X1_LOC_51/Y OR2X1_LOC_626/a_8_216# 0.00fF
C27149 OR2X1_LOC_97/A OR2X1_LOC_814/A 0.07fF
C27150 OR2X1_LOC_426/B OR2X1_LOC_106/A 0.01fF
C27151 AND2X1_LOC_348/Y OR2X1_LOC_91/A 0.03fF
C27152 AND2X1_LOC_521/a_36_24# OR2X1_LOC_404/Y -0.00fF
C27153 OR2X1_LOC_155/A OR2X1_LOC_803/A 0.36fF
C27154 AND2X1_LOC_498/a_36_24# OR2X1_LOC_203/Y -0.02fF
C27155 OR2X1_LOC_432/a_8_216# OR2X1_LOC_48/B 0.03fF
C27156 AND2X1_LOC_214/A OR2X1_LOC_36/Y 0.02fF
C27157 AND2X1_LOC_391/Y OR2X1_LOC_753/A 0.07fF
C27158 OR2X1_LOC_596/Y AND2X1_LOC_41/A 0.12fF
C27159 OR2X1_LOC_591/Y OR2X1_LOC_64/Y 0.01fF
C27160 OR2X1_LOC_3/Y OR2X1_LOC_694/Y 0.03fF
C27161 OR2X1_LOC_91/A OR2X1_LOC_753/A 0.07fF
C27162 OR2X1_LOC_160/B OR2X1_LOC_624/B 0.49fF
C27163 AND2X1_LOC_51/Y OR2X1_LOC_768/a_36_216# 0.00fF
C27164 AND2X1_LOC_12/Y AND2X1_LOC_422/a_8_24# 0.03fF
C27165 OR2X1_LOC_432/a_8_216# OR2X1_LOC_18/Y 0.01fF
C27166 OR2X1_LOC_499/B OR2X1_LOC_203/Y 0.15fF
C27167 OR2X1_LOC_252/a_8_216# AND2X1_LOC_805/Y 0.01fF
C27168 OR2X1_LOC_474/a_8_216# OR2X1_LOC_113/B 0.01fF
C27169 AND2X1_LOC_784/A AND2X1_LOC_477/a_8_24# 0.02fF
C27170 OR2X1_LOC_51/Y AND2X1_LOC_639/a_8_24# 0.01fF
C27171 OR2X1_LOC_401/Y OR2X1_LOC_78/B 0.01fF
C27172 OR2X1_LOC_666/A OR2X1_LOC_279/a_8_216# 0.01fF
C27173 AND2X1_LOC_86/Y OR2X1_LOC_160/A 0.08fF
C27174 AND2X1_LOC_12/Y OR2X1_LOC_865/B 0.05fF
C27175 INPUT_5 OR2X1_LOC_44/Y 0.04fF
C27176 OR2X1_LOC_154/A AND2X1_LOC_57/a_8_24# 0.03fF
C27177 AND2X1_LOC_367/A OR2X1_LOC_585/A 0.05fF
C27178 OR2X1_LOC_506/A OR2X1_LOC_739/A 0.03fF
C27179 OR2X1_LOC_619/Y AND2X1_LOC_621/Y 0.33fF
C27180 VDD OR2X1_LOC_486/a_8_216# 0.00fF
C27181 OR2X1_LOC_335/a_36_216# OR2X1_LOC_223/A 0.00fF
C27182 AND2X1_LOC_70/Y AND2X1_LOC_122/a_8_24# 0.01fF
C27183 OR2X1_LOC_859/A OR2X1_LOC_113/B 0.01fF
C27184 D_GATE_662 OR2X1_LOC_814/A 0.02fF
C27185 AND2X1_LOC_512/Y OR2X1_LOC_312/Y 0.20fF
C27186 OR2X1_LOC_48/B OR2X1_LOC_48/a_36_216# 0.01fF
C27187 AND2X1_LOC_847/Y AND2X1_LOC_848/Y 0.02fF
C27188 AND2X1_LOC_113/a_8_24# OR2X1_LOC_26/Y 0.03fF
C27189 OR2X1_LOC_11/a_8_216# D_INPUT_6 0.01fF
C27190 AND2X1_LOC_31/Y OR2X1_LOC_593/B 0.02fF
C27191 OR2X1_LOC_405/A OR2X1_LOC_358/B 0.03fF
C27192 AND2X1_LOC_787/A OR2X1_LOC_47/Y 0.03fF
C27193 OR2X1_LOC_62/A AND2X1_LOC_277/a_8_24# 0.01fF
C27194 OR2X1_LOC_335/B OR2X1_LOC_543/A 0.38fF
C27195 OR2X1_LOC_18/Y AND2X1_LOC_287/Y 0.02fF
C27196 OR2X1_LOC_689/A AND2X1_LOC_688/a_36_24# 0.00fF
C27197 OR2X1_LOC_703/B AND2X1_LOC_59/Y 0.02fF
C27198 OR2X1_LOC_45/B AND2X1_LOC_687/a_8_24# 0.01fF
C27199 AND2X1_LOC_804/Y OR2X1_LOC_52/B 0.03fF
C27200 OR2X1_LOC_165/Y OR2X1_LOC_74/A 0.06fF
C27201 OR2X1_LOC_479/Y OR2X1_LOC_776/a_8_216# 0.01fF
C27202 OR2X1_LOC_426/B OR2X1_LOC_46/A 0.10fF
C27203 OR2X1_LOC_201/A OR2X1_LOC_201/Y 0.07fF
C27204 AND2X1_LOC_663/B OR2X1_LOC_755/a_36_216# 0.00fF
C27205 AND2X1_LOC_59/Y OR2X1_LOC_87/A 0.38fF
C27206 OR2X1_LOC_465/Y OR2X1_LOC_465/B 0.01fF
C27207 OR2X1_LOC_300/a_36_216# OR2X1_LOC_300/Y 0.00fF
C27208 AND2X1_LOC_363/B OR2X1_LOC_3/Y 0.01fF
C27209 OR2X1_LOC_124/B D_INPUT_0 0.06fF
C27210 AND2X1_LOC_699/a_36_24# OR2X1_LOC_155/A -0.01fF
C27211 AND2X1_LOC_573/A OR2X1_LOC_753/A 0.50fF
C27212 OR2X1_LOC_154/A OR2X1_LOC_687/Y 0.07fF
C27213 OR2X1_LOC_287/B OR2X1_LOC_847/A 1.34fF
C27214 OR2X1_LOC_693/a_8_216# OR2X1_LOC_47/Y 0.06fF
C27215 AND2X1_LOC_580/B OR2X1_LOC_616/Y 0.03fF
C27216 OR2X1_LOC_70/Y OR2X1_LOC_92/Y 0.47fF
C27217 OR2X1_LOC_631/B OR2X1_LOC_500/A 0.01fF
C27218 AND2X1_LOC_89/a_36_24# OR2X1_LOC_375/A 0.00fF
C27219 INPUT_5 AND2X1_LOC_1/Y 0.01fF
C27220 OR2X1_LOC_379/Y AND2X1_LOC_3/Y 0.59fF
C27221 OR2X1_LOC_104/a_8_216# INPUT_1 0.01fF
C27222 AND2X1_LOC_779/a_36_24# OR2X1_LOC_89/A 0.00fF
C27223 AND2X1_LOC_191/B OR2X1_LOC_226/a_8_216# 0.06fF
C27224 OR2X1_LOC_604/A AND2X1_LOC_810/Y 0.10fF
C27225 OR2X1_LOC_188/Y OR2X1_LOC_675/Y 0.00fF
C27226 AND2X1_LOC_84/a_8_24# OR2X1_LOC_69/A 0.01fF
C27227 AND2X1_LOC_566/B OR2X1_LOC_47/Y 0.02fF
C27228 AND2X1_LOC_578/A OR2X1_LOC_531/a_8_216# 0.03fF
C27229 OR2X1_LOC_7/A AND2X1_LOC_436/B 0.07fF
C27230 OR2X1_LOC_375/A OR2X1_LOC_711/A 0.01fF
C27231 OR2X1_LOC_511/Y OR2X1_LOC_52/B 3.83fF
C27232 OR2X1_LOC_680/A OR2X1_LOC_626/a_8_216# 0.03fF
C27233 OR2X1_LOC_403/A AND2X1_LOC_51/Y 0.01fF
C27234 AND2X1_LOC_211/B AND2X1_LOC_655/A 0.10fF
C27235 OR2X1_LOC_736/Y OR2X1_LOC_241/B 0.19fF
C27236 OR2X1_LOC_426/B AND2X1_LOC_227/Y 0.03fF
C27237 AND2X1_LOC_376/a_36_24# OR2X1_LOC_459/B 0.00fF
C27238 AND2X1_LOC_139/B OR2X1_LOC_7/A 0.00fF
C27239 AND2X1_LOC_570/Y OR2X1_LOC_95/Y 0.03fF
C27240 AND2X1_LOC_99/Y AND2X1_LOC_101/a_8_24# 0.07fF
C27241 AND2X1_LOC_514/Y OR2X1_LOC_92/Y 0.07fF
C27242 OR2X1_LOC_331/A OR2X1_LOC_95/Y 0.18fF
C27243 OR2X1_LOC_324/B OR2X1_LOC_532/B 0.23fF
C27244 OR2X1_LOC_858/B OR2X1_LOC_814/A 0.01fF
C27245 VDD AND2X1_LOC_109/a_8_24# -0.00fF
C27246 OR2X1_LOC_702/A OR2X1_LOC_805/A 0.08fF
C27247 AND2X1_LOC_620/Y AND2X1_LOC_254/a_8_24# 0.05fF
C27248 AND2X1_LOC_395/a_36_24# AND2X1_LOC_3/Y 0.00fF
C27249 OR2X1_LOC_329/B OR2X1_LOC_31/Y 0.05fF
C27250 OR2X1_LOC_194/Y AND2X1_LOC_3/Y 3.07fF
C27251 OR2X1_LOC_36/Y AND2X1_LOC_645/A 0.03fF
C27252 OR2X1_LOC_70/Y OR2X1_LOC_65/B 0.03fF
C27253 INPUT_2 D_INPUT_1 0.10fF
C27254 OR2X1_LOC_653/a_36_216# OR2X1_LOC_130/A 0.01fF
C27255 OR2X1_LOC_114/Y AND2X1_LOC_3/Y 0.03fF
C27256 AND2X1_LOC_303/B OR2X1_LOC_299/Y 0.80fF
C27257 OR2X1_LOC_13/Y OR2X1_LOC_311/a_36_216# 0.00fF
C27258 OR2X1_LOC_16/A OR2X1_LOC_331/Y 0.00fF
C27259 AND2X1_LOC_42/a_8_24# OR2X1_LOC_83/A 0.01fF
C27260 OR2X1_LOC_624/A OR2X1_LOC_121/B 0.05fF
C27261 AND2X1_LOC_427/a_8_24# OR2X1_LOC_161/B 0.15fF
C27262 AND2X1_LOC_67/a_8_24# OR2X1_LOC_241/Y 0.04fF
C27263 OR2X1_LOC_403/B AND2X1_LOC_79/Y 0.04fF
C27264 OR2X1_LOC_114/B OR2X1_LOC_493/Y 0.03fF
C27265 OR2X1_LOC_446/Y AND2X1_LOC_424/a_8_24# 0.02fF
C27266 OR2X1_LOC_130/A AND2X1_LOC_51/Y 0.08fF
C27267 AND2X1_LOC_142/a_8_24# OR2X1_LOC_532/B 0.01fF
C27268 AND2X1_LOC_95/Y OR2X1_LOC_46/A 0.20fF
C27269 OR2X1_LOC_476/B OR2X1_LOC_805/A 0.03fF
C27270 OR2X1_LOC_74/A OR2X1_LOC_585/A 0.02fF
C27271 OR2X1_LOC_529/Y OR2X1_LOC_7/A 0.06fF
C27272 OR2X1_LOC_263/a_8_216# OR2X1_LOC_18/Y 0.01fF
C27273 OR2X1_LOC_22/Y OR2X1_LOC_413/Y 0.06fF
C27274 OR2X1_LOC_62/B OR2X1_LOC_161/A 0.29fF
C27275 OR2X1_LOC_74/Y OR2X1_LOC_31/Y 0.02fF
C27276 OR2X1_LOC_274/Y OR2X1_LOC_276/B 0.01fF
C27277 AND2X1_LOC_44/Y OR2X1_LOC_71/A 0.85fF
C27278 AND2X1_LOC_314/a_8_24# OR2X1_LOC_532/B 0.01fF
C27279 OR2X1_LOC_447/Y OR2X1_LOC_724/a_36_216# 0.02fF
C27280 OR2X1_LOC_753/A OR2X1_LOC_27/Y 0.03fF
C27281 D_INPUT_4 OR2X1_LOC_651/A 0.42fF
C27282 OR2X1_LOC_626/a_36_216# OR2X1_LOC_617/Y 0.00fF
C27283 OR2X1_LOC_677/Y AND2X1_LOC_803/a_8_24# 0.23fF
C27284 INPUT_0 OR2X1_LOC_41/a_8_216# 0.01fF
C27285 AND2X1_LOC_196/a_8_24# OR2X1_LOC_485/A 0.08fF
C27286 OR2X1_LOC_160/A OR2X1_LOC_244/A 0.08fF
C27287 OR2X1_LOC_373/Y OR2X1_LOC_164/a_36_216# 0.00fF
C27288 OR2X1_LOC_243/A OR2X1_LOC_532/B 0.01fF
C27289 AND2X1_LOC_47/Y OR2X1_LOC_347/B 0.01fF
C27290 AND2X1_LOC_160/Y OR2X1_LOC_163/Y 0.00fF
C27291 OR2X1_LOC_532/B OR2X1_LOC_668/Y 0.02fF
C27292 AND2X1_LOC_108/a_36_24# OR2X1_LOC_161/A 0.00fF
C27293 OR2X1_LOC_36/Y AND2X1_LOC_477/A 0.03fF
C27294 AND2X1_LOC_47/Y OR2X1_LOC_539/Y 0.08fF
C27295 INPUT_1 OR2X1_LOC_6/A 0.57fF
C27296 OR2X1_LOC_810/A AND2X1_LOC_107/a_8_24# 0.22fF
C27297 OR2X1_LOC_654/A OR2X1_LOC_19/B 0.03fF
C27298 OR2X1_LOC_776/A OR2X1_LOC_121/A 0.16fF
C27299 OR2X1_LOC_405/A OR2X1_LOC_112/B 0.03fF
C27300 OR2X1_LOC_316/Y AND2X1_LOC_476/A 0.00fF
C27301 OR2X1_LOC_19/B OR2X1_LOC_609/a_8_216# 0.05fF
C27302 OR2X1_LOC_532/B OR2X1_LOC_719/Y 0.00fF
C27303 OR2X1_LOC_612/a_8_216# OR2X1_LOC_71/A 0.01fF
C27304 OR2X1_LOC_327/a_8_216# OR2X1_LOC_205/Y 0.06fF
C27305 OR2X1_LOC_447/Y OR2X1_LOC_449/B 0.00fF
C27306 AND2X1_LOC_420/a_8_24# OR2X1_LOC_739/A 0.01fF
C27307 OR2X1_LOC_600/A OR2X1_LOC_71/A 0.07fF
C27308 OR2X1_LOC_743/A OR2X1_LOC_46/A 0.14fF
C27309 OR2X1_LOC_390/A OR2X1_LOC_174/Y 0.00fF
C27310 AND2X1_LOC_116/B AND2X1_LOC_116/Y 0.26fF
C27311 OR2X1_LOC_56/A OR2X1_LOC_384/a_8_216# 0.01fF
C27312 AND2X1_LOC_690/a_8_24# OR2X1_LOC_598/A 0.08fF
C27313 OR2X1_LOC_78/A OR2X1_LOC_546/A 0.01fF
C27314 AND2X1_LOC_41/A OR2X1_LOC_789/A 0.03fF
C27315 OR2X1_LOC_495/a_8_216# AND2X1_LOC_851/B 0.04fF
C27316 OR2X1_LOC_154/A OR2X1_LOC_786/Y 0.10fF
C27317 AND2X1_LOC_86/B OR2X1_LOC_244/A 0.05fF
C27318 OR2X1_LOC_26/Y AND2X1_LOC_796/Y 0.00fF
C27319 AND2X1_LOC_242/B OR2X1_LOC_184/a_36_216# 0.01fF
C27320 OR2X1_LOC_683/Y AND2X1_LOC_686/a_8_24# 0.23fF
C27321 OR2X1_LOC_62/B AND2X1_LOC_51/Y 0.03fF
C27322 AND2X1_LOC_12/Y OR2X1_LOC_493/Y 0.09fF
C27323 AND2X1_LOC_12/Y OR2X1_LOC_801/B 0.01fF
C27324 OR2X1_LOC_223/A OR2X1_LOC_778/Y 0.05fF
C27325 AND2X1_LOC_92/Y OR2X1_LOC_704/a_36_216# 0.02fF
C27326 OR2X1_LOC_161/A OR2X1_LOC_365/B 0.04fF
C27327 OR2X1_LOC_269/B OR2X1_LOC_284/B 0.00fF
C27328 OR2X1_LOC_244/Y OR2X1_LOC_349/B 0.00fF
C27329 OR2X1_LOC_858/A OR2X1_LOC_580/A 0.18fF
C27330 OR2X1_LOC_831/a_8_216# OR2X1_LOC_804/A 0.03fF
C27331 OR2X1_LOC_529/Y OR2X1_LOC_224/a_8_216# 0.01fF
C27332 OR2X1_LOC_89/A AND2X1_LOC_796/Y 0.03fF
C27333 AND2X1_LOC_807/Y OR2X1_LOC_406/A 0.02fF
C27334 OR2X1_LOC_269/B D_INPUT_1 3.89fF
C27335 AND2X1_LOC_619/B OR2X1_LOC_80/A 0.02fF
C27336 OR2X1_LOC_246/A OR2X1_LOC_46/A 0.03fF
C27337 OR2X1_LOC_302/A OR2X1_LOC_308/Y 0.14fF
C27338 OR2X1_LOC_653/Y OR2X1_LOC_68/B 0.07fF
C27339 AND2X1_LOC_70/Y OR2X1_LOC_374/a_8_216# 0.17fF
C27340 OR2X1_LOC_464/A OR2X1_LOC_367/B 0.15fF
C27341 OR2X1_LOC_86/A OR2X1_LOC_85/A 0.71fF
C27342 OR2X1_LOC_18/Y AND2X1_LOC_562/Y 0.40fF
C27343 OR2X1_LOC_447/Y OR2X1_LOC_121/B 0.46fF
C27344 VDD OR2X1_LOC_308/Y 0.12fF
C27345 OR2X1_LOC_481/A AND2X1_LOC_866/A 0.05fF
C27346 AND2X1_LOC_512/Y OR2X1_LOC_13/B 0.04fF
C27347 OR2X1_LOC_44/Y AND2X1_LOC_228/a_8_24# 0.01fF
C27348 OR2X1_LOC_269/B AND2X1_LOC_48/Y 0.01fF
C27349 OR2X1_LOC_188/Y OR2X1_LOC_736/Y 0.03fF
C27350 OR2X1_LOC_51/B OR2X1_LOC_17/Y 0.38fF
C27351 OR2X1_LOC_162/A OR2X1_LOC_160/Y 0.06fF
C27352 AND2X1_LOC_227/Y OR2X1_LOC_246/A 0.10fF
C27353 OR2X1_LOC_619/Y OR2X1_LOC_71/A 0.07fF
C27354 AND2X1_LOC_810/A AND2X1_LOC_810/B 0.16fF
C27355 OR2X1_LOC_703/A OR2X1_LOC_469/B 0.67fF
C27356 OR2X1_LOC_696/A AND2X1_LOC_434/Y 0.18fF
C27357 OR2X1_LOC_547/B OR2X1_LOC_550/B 0.00fF
C27358 AND2X1_LOC_22/Y AND2X1_LOC_262/a_36_24# 0.01fF
C27359 D_INPUT_2 INPUT_1 0.12fF
C27360 OR2X1_LOC_168/B OR2X1_LOC_390/B 0.01fF
C27361 AND2X1_LOC_866/A OR2X1_LOC_71/Y 0.03fF
C27362 OR2X1_LOC_392/B OR2X1_LOC_66/A 0.03fF
C27363 AND2X1_LOC_743/a_8_24# OR2X1_LOC_160/B 0.01fF
C27364 AND2X1_LOC_263/a_8_24# OR2X1_LOC_66/A 0.01fF
C27365 OR2X1_LOC_646/A OR2X1_LOC_68/B 0.14fF
C27366 AND2X1_LOC_51/Y OR2X1_LOC_365/B 0.03fF
C27367 VDD AND2X1_LOC_604/a_8_24# 0.00fF
C27368 AND2X1_LOC_340/Y AND2X1_LOC_340/a_8_24# 0.00fF
C27369 AND2X1_LOC_342/Y OR2X1_LOC_13/B 0.04fF
C27370 AND2X1_LOC_715/Y AND2X1_LOC_434/Y 0.10fF
C27371 VDD AND2X1_LOC_455/B 0.03fF
C27372 AND2X1_LOC_851/B OR2X1_LOC_238/a_8_216# 0.04fF
C27373 AND2X1_LOC_656/Y AND2X1_LOC_660/A 0.00fF
C27374 OR2X1_LOC_246/A OR2X1_LOC_813/Y 0.12fF
C27375 OR2X1_LOC_448/Y OR2X1_LOC_712/B 0.02fF
C27376 OR2X1_LOC_334/B OR2X1_LOC_334/a_8_216# 0.07fF
C27377 AND2X1_LOC_90/a_8_24# VDD 0.00fF
C27378 OR2X1_LOC_768/A AND2X1_LOC_22/Y 0.02fF
C27379 OR2X1_LOC_738/A OR2X1_LOC_209/A 0.02fF
C27380 OR2X1_LOC_604/A OR2X1_LOC_671/Y 0.00fF
C27381 OR2X1_LOC_858/A AND2X1_LOC_44/Y 0.03fF
C27382 AND2X1_LOC_537/a_8_24# OR2X1_LOC_829/A 0.09fF
C27383 OR2X1_LOC_604/A AND2X1_LOC_714/B 0.12fF
C27384 OR2X1_LOC_47/Y AND2X1_LOC_675/A 0.00fF
C27385 OR2X1_LOC_45/B AND2X1_LOC_548/Y 0.03fF
C27386 AND2X1_LOC_92/Y OR2X1_LOC_161/B 0.07fF
C27387 AND2X1_LOC_477/A OR2X1_LOC_419/Y 0.07fF
C27388 OR2X1_LOC_49/A AND2X1_LOC_94/Y -0.01fF
C27389 OR2X1_LOC_160/B OR2X1_LOC_768/a_8_216# 0.02fF
C27390 VDD OR2X1_LOC_421/Y 0.26fF
C27391 OR2X1_LOC_113/B OR2X1_LOC_66/A 0.00fF
C27392 AND2X1_LOC_721/Y AND2X1_LOC_456/B 0.01fF
C27393 AND2X1_LOC_522/a_8_24# OR2X1_LOC_235/B 0.01fF
C27394 AND2X1_LOC_22/Y AND2X1_LOC_71/a_8_24# 0.03fF
C27395 AND2X1_LOC_216/Y AND2X1_LOC_218/a_8_24# 0.18fF
C27396 OR2X1_LOC_123/a_36_216# OR2X1_LOC_549/A 0.01fF
C27397 OR2X1_LOC_429/a_8_216# OR2X1_LOC_70/A 0.01fF
C27398 OR2X1_LOC_371/Y OR2X1_LOC_437/A 0.10fF
C27399 AND2X1_LOC_749/a_8_24# AND2X1_LOC_44/Y 0.03fF
C27400 AND2X1_LOC_42/B OR2X1_LOC_140/Y 0.37fF
C27401 AND2X1_LOC_392/A AND2X1_LOC_112/a_8_24# 0.03fF
C27402 AND2X1_LOC_95/Y OR2X1_LOC_556/a_36_216# 0.02fF
C27403 VDD OR2X1_LOC_800/Y 0.00fF
C27404 OR2X1_LOC_279/a_8_216# OR2X1_LOC_13/B 0.03fF
C27405 OR2X1_LOC_663/A OR2X1_LOC_659/Y 0.10fF
C27406 OR2X1_LOC_95/Y OR2X1_LOC_406/A 0.00fF
C27407 OR2X1_LOC_97/A OR2X1_LOC_147/B 0.03fF
C27408 OR2X1_LOC_269/B OR2X1_LOC_180/B 0.03fF
C27409 OR2X1_LOC_377/A OR2X1_LOC_20/A 0.14fF
C27410 OR2X1_LOC_51/B OR2X1_LOC_588/A 0.09fF
C27411 OR2X1_LOC_45/B OR2X1_LOC_46/a_36_216# 0.02fF
C27412 AND2X1_LOC_719/Y AND2X1_LOC_474/A 0.05fF
C27413 OR2X1_LOC_648/A AND2X1_LOC_18/Y 0.35fF
C27414 AND2X1_LOC_64/Y OR2X1_LOC_510/Y 0.04fF
C27415 AND2X1_LOC_840/B OR2X1_LOC_525/a_8_216# 0.04fF
C27416 AND2X1_LOC_41/A OR2X1_LOC_307/A 0.01fF
C27417 OR2X1_LOC_600/A OR2X1_LOC_59/Y 1.78fF
C27418 OR2X1_LOC_51/Y AND2X1_LOC_436/Y 0.83fF
C27419 OR2X1_LOC_91/Y AND2X1_LOC_543/Y 0.03fF
C27420 AND2X1_LOC_776/a_8_24# OR2X1_LOC_56/A 0.01fF
C27421 OR2X1_LOC_427/A AND2X1_LOC_786/Y 0.09fF
C27422 OR2X1_LOC_151/A OR2X1_LOC_216/A 0.07fF
C27423 OR2X1_LOC_45/B AND2X1_LOC_702/a_8_24# 0.01fF
C27424 OR2X1_LOC_614/Y AND2X1_LOC_615/a_8_24# 0.00fF
C27425 OR2X1_LOC_280/Y OR2X1_LOC_183/Y 0.03fF
C27426 AND2X1_LOC_214/A AND2X1_LOC_207/B 0.83fF
C27427 OR2X1_LOC_380/a_8_216# OR2X1_LOC_380/Y -0.00fF
C27428 AND2X1_LOC_847/a_8_24# AND2X1_LOC_789/Y 0.01fF
C27429 AND2X1_LOC_675/Y AND2X1_LOC_508/B 0.02fF
C27430 AND2X1_LOC_722/a_8_24# AND2X1_LOC_723/Y -0.00fF
C27431 OR2X1_LOC_46/A OR2X1_LOC_599/a_8_216# 0.14fF
C27432 AND2X1_LOC_658/Y AND2X1_LOC_659/a_8_24# 0.01fF
C27433 OR2X1_LOC_785/a_36_216# AND2X1_LOC_92/Y 0.01fF
C27434 OR2X1_LOC_535/A OR2X1_LOC_620/Y -0.01fF
C27435 AND2X1_LOC_529/a_8_24# OR2X1_LOC_66/A 0.04fF
C27436 OR2X1_LOC_54/Y OR2X1_LOC_13/B 0.01fF
C27437 AND2X1_LOC_191/B AND2X1_LOC_663/A 0.00fF
C27438 OR2X1_LOC_747/a_36_216# AND2X1_LOC_781/Y 0.00fF
C27439 OR2X1_LOC_325/B OR2X1_LOC_808/B 0.30fF
C27440 AND2X1_LOC_509/Y AND2X1_LOC_509/a_8_24# 0.01fF
C27441 AND2X1_LOC_663/A AND2X1_LOC_469/B 0.05fF
C27442 AND2X1_LOC_711/a_8_24# OR2X1_LOC_59/Y 0.02fF
C27443 AND2X1_LOC_64/Y OR2X1_LOC_810/A 0.06fF
C27444 OR2X1_LOC_505/a_8_216# AND2X1_LOC_807/Y 0.16fF
C27445 OR2X1_LOC_53/Y OR2X1_LOC_44/Y 0.06fF
C27446 AND2X1_LOC_315/a_36_24# OR2X1_LOC_161/B 0.01fF
C27447 OR2X1_LOC_709/A AND2X1_LOC_748/a_8_24# 0.03fF
C27448 OR2X1_LOC_266/a_8_216# OR2X1_LOC_266/A 0.18fF
C27449 AND2X1_LOC_733/a_36_24# OR2X1_LOC_40/Y 0.00fF
C27450 OR2X1_LOC_359/a_8_216# OR2X1_LOC_850/B 0.01fF
C27451 OR2X1_LOC_91/A AND2X1_LOC_222/a_8_24# 0.03fF
C27452 AND2X1_LOC_464/a_8_24# AND2X1_LOC_786/Y 0.02fF
C27453 OR2X1_LOC_786/Y OR2X1_LOC_560/A 0.16fF
C27454 AND2X1_LOC_810/A AND2X1_LOC_354/a_8_24# 0.01fF
C27455 OR2X1_LOC_551/B OR2X1_LOC_365/B 0.06fF
C27456 AND2X1_LOC_70/Y OR2X1_LOC_274/Y 0.00fF
C27457 OR2X1_LOC_176/Y AND2X1_LOC_661/A 0.00fF
C27458 AND2X1_LOC_703/Y OR2X1_LOC_36/Y 0.03fF
C27459 AND2X1_LOC_231/a_8_24# OR2X1_LOC_52/B 0.03fF
C27460 OR2X1_LOC_271/a_8_216# AND2X1_LOC_786/Y 0.04fF
C27461 OR2X1_LOC_151/A OR2X1_LOC_499/a_8_216# 0.01fF
C27462 AND2X1_LOC_323/a_8_24# OR2X1_LOC_620/Y 0.01fF
C27463 AND2X1_LOC_862/Y OR2X1_LOC_59/Y 0.14fF
C27464 OR2X1_LOC_833/B AND2X1_LOC_626/a_36_24# 0.01fF
C27465 OR2X1_LOC_599/A AND2X1_LOC_714/a_8_24# 0.00fF
C27466 OR2X1_LOC_287/B OR2X1_LOC_474/B 0.03fF
C27467 AND2X1_LOC_701/a_8_24# AND2X1_LOC_44/Y 0.01fF
C27468 VDD OR2X1_LOC_278/Y 0.31fF
C27469 AND2X1_LOC_564/B OR2X1_LOC_74/A 0.07fF
C27470 OR2X1_LOC_405/a_8_216# AND2X1_LOC_18/Y 0.02fF
C27471 AND2X1_LOC_721/Y AND2X1_LOC_717/B 0.06fF
C27472 AND2X1_LOC_11/a_8_24# INPUT_6 0.00fF
C27473 OR2X1_LOC_492/a_8_216# OR2X1_LOC_36/Y 0.01fF
C27474 OR2X1_LOC_379/a_8_216# OR2X1_LOC_598/Y 0.01fF
C27475 OR2X1_LOC_91/Y OR2X1_LOC_322/Y 0.07fF
C27476 VDD AND2X1_LOC_662/B 0.21fF
C27477 OR2X1_LOC_302/B OR2X1_LOC_147/B 0.14fF
C27478 OR2X1_LOC_405/A OR2X1_LOC_493/B 0.02fF
C27479 OR2X1_LOC_74/A OR2X1_LOC_368/Y 0.11fF
C27480 OR2X1_LOC_61/Y AND2X1_LOC_92/Y 0.07fF
C27481 OR2X1_LOC_9/Y OR2X1_LOC_246/Y 0.35fF
C27482 OR2X1_LOC_203/a_8_216# AND2X1_LOC_18/Y 0.01fF
C27483 OR2X1_LOC_530/Y OR2X1_LOC_816/A 0.02fF
C27484 OR2X1_LOC_151/A OR2X1_LOC_468/Y 0.05fF
C27485 OR2X1_LOC_210/B OR2X1_LOC_160/Y 0.05fF
C27486 AND2X1_LOC_734/Y AND2X1_LOC_737/a_8_24# 0.01fF
C27487 AND2X1_LOC_64/Y OR2X1_LOC_857/a_8_216# 0.06fF
C27488 OR2X1_LOC_64/Y AND2X1_LOC_227/a_8_24# 0.01fF
C27489 AND2X1_LOC_59/Y OR2X1_LOC_389/A 0.01fF
C27490 OR2X1_LOC_574/A AND2X1_LOC_433/a_8_24# 0.26fF
C27491 AND2X1_LOC_541/Y AND2X1_LOC_560/B 0.24fF
C27492 AND2X1_LOC_59/Y OR2X1_LOC_493/a_8_216# 0.01fF
C27493 AND2X1_LOC_866/A AND2X1_LOC_789/Y 0.10fF
C27494 OR2X1_LOC_507/a_8_216# OR2X1_LOC_502/A 0.01fF
C27495 VDD OR2X1_LOC_95/a_8_216# 0.21fF
C27496 OR2X1_LOC_524/Y OR2X1_LOC_427/A 0.01fF
C27497 OR2X1_LOC_619/Y OR2X1_LOC_59/Y 0.10fF
C27498 OR2X1_LOC_532/B OR2X1_LOC_508/Y 0.15fF
C27499 OR2X1_LOC_264/Y OR2X1_LOC_502/A 0.03fF
C27500 OR2X1_LOC_680/A AND2X1_LOC_436/Y 0.18fF
C27501 OR2X1_LOC_51/Y OR2X1_LOC_603/a_8_216# 0.01fF
C27502 VDD AND2X1_LOC_565/Y 0.04fF
C27503 OR2X1_LOC_849/A OR2X1_LOC_772/A 0.00fF
C27504 D_INPUT_0 OR2X1_LOC_171/a_8_216# 0.02fF
C27505 OR2X1_LOC_482/Y AND2X1_LOC_717/B 0.05fF
C27506 OR2X1_LOC_145/a_8_216# OR2X1_LOC_51/Y 0.01fF
C27507 VDD OR2X1_LOC_151/Y 0.04fF
C27508 OR2X1_LOC_600/A OR2X1_LOC_820/B 0.04fF
C27509 INPUT_0 OR2X1_LOC_316/Y 0.02fF
C27510 OR2X1_LOC_491/a_36_216# OR2X1_LOC_529/Y 0.00fF
C27511 VDD AND2X1_LOC_472/B 0.21fF
C27512 OR2X1_LOC_604/A AND2X1_LOC_645/A 0.12fF
C27513 OR2X1_LOC_756/B AND2X1_LOC_43/B 0.42fF
C27514 OR2X1_LOC_51/a_8_216# D_INPUT_6 0.01fF
C27515 OR2X1_LOC_175/Y OR2X1_LOC_814/A 0.00fF
C27516 OR2X1_LOC_865/A OR2X1_LOC_859/A 0.19fF
C27517 OR2X1_LOC_485/A AND2X1_LOC_243/Y 0.03fF
C27518 OR2X1_LOC_51/Y OR2X1_LOC_588/Y 0.03fF
C27519 AND2X1_LOC_64/Y AND2X1_LOC_56/a_8_24# 0.02fF
C27520 INPUT_0 OR2X1_LOC_194/Y 0.02fF
C27521 OR2X1_LOC_158/A OR2X1_LOC_44/a_36_216# 0.02fF
C27522 VDD OR2X1_LOC_593/A -0.00fF
C27523 OR2X1_LOC_666/A OR2X1_LOC_26/Y 0.02fF
C27524 OR2X1_LOC_696/A AND2X1_LOC_851/B 0.45fF
C27525 OR2X1_LOC_107/a_8_216# AND2X1_LOC_560/B 0.01fF
C27526 OR2X1_LOC_395/a_8_216# OR2X1_LOC_29/a_8_216# 0.47fF
C27527 INPUT_0 AND2X1_LOC_354/B 0.19fF
C27528 AND2X1_LOC_56/B OR2X1_LOC_630/B 0.01fF
C27529 VDD AND2X1_LOC_337/B 0.39fF
C27530 AND2X1_LOC_222/Y OR2X1_LOC_437/A 0.05fF
C27531 AND2X1_LOC_792/Y AND2X1_LOC_792/B 0.83fF
C27532 OR2X1_LOC_860/a_8_216# OR2X1_LOC_865/B 0.06fF
C27533 AND2X1_LOC_784/A OR2X1_LOC_91/A 0.10fF
C27534 AND2X1_LOC_523/a_8_24# AND2X1_LOC_76/Y 0.01fF
C27535 OR2X1_LOC_814/A AND2X1_LOC_417/a_8_24# -0.01fF
C27536 AND2X1_LOC_12/Y OR2X1_LOC_61/B 0.03fF
C27537 OR2X1_LOC_97/A OR2X1_LOC_545/B 0.17fF
C27538 OR2X1_LOC_589/A OR2X1_LOC_291/Y 0.03fF
C27539 OR2X1_LOC_856/B OR2X1_LOC_624/A 0.13fF
C27540 AND2X1_LOC_81/B AND2X1_LOC_316/a_8_24# 0.09fF
C27541 OR2X1_LOC_40/Y OR2X1_LOC_481/A 0.06fF
C27542 AND2X1_LOC_711/Y OR2X1_LOC_600/A 0.03fF
C27543 OR2X1_LOC_666/A OR2X1_LOC_89/A 0.03fF
C27544 AND2X1_LOC_124/a_8_24# OR2X1_LOC_92/Y 0.06fF
C27545 OR2X1_LOC_244/A OR2X1_LOC_266/A 0.05fF
C27546 AND2X1_LOC_325/a_36_24# OR2X1_LOC_74/A 0.01fF
C27547 OR2X1_LOC_48/B OR2X1_LOC_432/Y 0.03fF
C27548 OR2X1_LOC_70/Y OR2X1_LOC_600/A 0.10fF
C27549 OR2X1_LOC_109/a_8_216# OR2X1_LOC_109/Y 0.01fF
C27550 OR2X1_LOC_414/a_8_216# OR2X1_LOC_394/Y 0.39fF
C27551 AND2X1_LOC_571/A OR2X1_LOC_47/Y 0.01fF
C27552 OR2X1_LOC_589/A OR2X1_LOC_311/Y 0.03fF
C27553 INPUT_3 OR2X1_LOC_847/A 0.25fF
C27554 VDD OR2X1_LOC_273/Y 0.23fF
C27555 AND2X1_LOC_557/a_36_24# OR2X1_LOC_600/A 0.01fF
C27556 VDD OR2X1_LOC_636/a_8_216# 0.21fF
C27557 OR2X1_LOC_299/Y OR2X1_LOC_56/A 0.04fF
C27558 AND2X1_LOC_91/B OR2X1_LOC_673/A 0.09fF
C27559 AND2X1_LOC_40/Y OR2X1_LOC_213/B 0.10fF
C27560 AND2X1_LOC_95/Y OR2X1_LOC_739/A 0.04fF
C27561 AND2X1_LOC_91/B OR2X1_LOC_223/A 0.05fF
C27562 AND2X1_LOC_12/Y OR2X1_LOC_194/B 0.01fF
C27563 AND2X1_LOC_70/Y OR2X1_LOC_636/B 0.01fF
C27564 OR2X1_LOC_476/B OR2X1_LOC_648/B 0.02fF
C27565 OR2X1_LOC_459/A OR2X1_LOC_585/A 0.15fF
C27566 OR2X1_LOC_154/A OR2X1_LOC_851/A 0.01fF
C27567 OR2X1_LOC_287/B OR2X1_LOC_561/Y 0.00fF
C27568 OR2X1_LOC_391/a_8_216# OR2X1_LOC_269/B 0.01fF
C27569 OR2X1_LOC_287/B OR2X1_LOC_78/Y 0.03fF
C27570 OR2X1_LOC_176/Y AND2X1_LOC_810/Y 0.01fF
C27571 OR2X1_LOC_309/a_8_216# OR2X1_LOC_22/Y 0.07fF
C27572 OR2X1_LOC_166/a_8_216# OR2X1_LOC_70/Y 0.01fF
C27573 OR2X1_LOC_643/A OR2X1_LOC_502/A 0.03fF
C27574 AND2X1_LOC_312/a_8_24# AND2X1_LOC_528/a_8_24# 0.23fF
C27575 OR2X1_LOC_121/B AND2X1_LOC_265/a_36_24# 0.00fF
C27576 OR2X1_LOC_821/Y OR2X1_LOC_813/A 0.00fF
C27577 OR2X1_LOC_468/A AND2X1_LOC_51/Y 0.00fF
C27578 AND2X1_LOC_711/a_8_24# AND2X1_LOC_711/Y 0.01fF
C27579 OR2X1_LOC_151/A OR2X1_LOC_471/Y 0.07fF
C27580 OR2X1_LOC_506/A OR2X1_LOC_539/Y 0.03fF
C27581 OR2X1_LOC_158/A OR2X1_LOC_412/a_8_216# 0.02fF
C27582 OR2X1_LOC_689/A AND2X1_LOC_472/B 0.03fF
C27583 AND2X1_LOC_390/B INPUT_0 0.02fF
C27584 OR2X1_LOC_502/A OR2X1_LOC_778/Y 0.10fF
C27585 AND2X1_LOC_514/Y OR2X1_LOC_600/A 0.07fF
C27586 OR2X1_LOC_307/a_8_216# OR2X1_LOC_512/A 0.48fF
C27587 AND2X1_LOC_508/A OR2X1_LOC_239/Y 0.01fF
C27588 OR2X1_LOC_865/B OR2X1_LOC_865/a_8_216# 0.04fF
C27589 OR2X1_LOC_850/a_8_216# OR2X1_LOC_850/A 0.02fF
C27590 AND2X1_LOC_514/Y AND2X1_LOC_335/Y 0.01fF
C27591 AND2X1_LOC_663/B OR2X1_LOC_700/a_8_216# 0.01fF
C27592 VDD OR2X1_LOC_19/B 1.34fF
C27593 OR2X1_LOC_241/B OR2X1_LOC_120/a_8_216# 0.02fF
C27594 OR2X1_LOC_133/a_8_216# OR2X1_LOC_95/Y 0.01fF
C27595 OR2X1_LOC_26/Y OR2X1_LOC_393/a_8_216# 0.00fF
C27596 OR2X1_LOC_737/A OR2X1_LOC_269/B 0.07fF
C27597 AND2X1_LOC_851/B OR2X1_LOC_522/a_36_216# 0.01fF
C27598 OR2X1_LOC_604/A AND2X1_LOC_477/A 0.09fF
C27599 OR2X1_LOC_107/a_8_216# OR2X1_LOC_64/Y 0.07fF
C27600 AND2X1_LOC_719/Y OR2X1_LOC_226/Y 0.07fF
C27601 OR2X1_LOC_529/a_8_216# AND2X1_LOC_560/B 0.01fF
C27602 OR2X1_LOC_643/A OR2X1_LOC_571/B 0.01fF
C27603 OR2X1_LOC_40/Y OR2X1_LOC_71/Y 0.03fF
C27604 AND2X1_LOC_95/Y OR2X1_LOC_269/B 0.48fF
C27605 OR2X1_LOC_251/Y OR2X1_LOC_278/Y 1.95fF
C27606 D_INPUT_7 OR2X1_LOC_2/Y 0.20fF
C27607 OR2X1_LOC_364/A AND2X1_LOC_601/a_8_24# 0.02fF
C27608 OR2X1_LOC_502/A OR2X1_LOC_647/A 0.01fF
C27609 AND2X1_LOC_196/Y AND2X1_LOC_199/a_36_24# 0.01fF
C27610 AND2X1_LOC_51/Y OR2X1_LOC_571/a_8_216# 0.01fF
C27611 OR2X1_LOC_449/B OR2X1_LOC_161/A 0.10fF
C27612 OR2X1_LOC_329/Y OR2X1_LOC_95/Y 0.01fF
C27613 OR2X1_LOC_585/A AND2X1_LOC_400/a_8_24# 0.03fF
C27614 OR2X1_LOC_669/A AND2X1_LOC_668/a_8_24# 0.11fF
C27615 OR2X1_LOC_474/a_8_216# OR2X1_LOC_624/Y 0.01fF
C27616 OR2X1_LOC_32/B OR2X1_LOC_753/A 0.10fF
C27617 OR2X1_LOC_532/B OR2X1_LOC_66/A 0.20fF
C27618 OR2X1_LOC_124/A OR2X1_LOC_814/A 0.07fF
C27619 OR2X1_LOC_405/A OR2X1_LOC_574/A 0.13fF
C27620 AND2X1_LOC_59/Y OR2X1_LOC_403/B 0.23fF
C27621 OR2X1_LOC_185/A OR2X1_LOC_564/A 0.00fF
C27622 AND2X1_LOC_184/a_8_24# AND2X1_LOC_47/Y 0.02fF
C27623 OR2X1_LOC_316/Y OR2X1_LOC_690/A 0.00fF
C27624 AND2X1_LOC_550/A OR2X1_LOC_438/a_8_216# 0.01fF
C27625 AND2X1_LOC_578/A OR2X1_LOC_427/A 0.10fF
C27626 OR2X1_LOC_454/a_8_216# OR2X1_LOC_466/A -0.00fF
C27627 AND2X1_LOC_665/a_8_24# OR2X1_LOC_66/A 0.02fF
C27628 OR2X1_LOC_849/a_8_216# OR2X1_LOC_659/A -0.02fF
C27629 OR2X1_LOC_859/A OR2X1_LOC_624/Y 0.03fF
C27630 OR2X1_LOC_189/A OR2X1_LOC_498/Y 0.01fF
C27631 OR2X1_LOC_267/A OR2X1_LOC_204/Y 0.68fF
C27632 AND2X1_LOC_502/a_8_24# OR2X1_LOC_89/A 0.01fF
C27633 AND2X1_LOC_456/B OR2X1_LOC_628/Y 0.50fF
C27634 OR2X1_LOC_283/a_36_216# AND2X1_LOC_859/Y 0.01fF
C27635 OR2X1_LOC_827/a_8_216# OR2X1_LOC_6/A 0.01fF
C27636 OR2X1_LOC_859/A OR2X1_LOC_391/A 0.04fF
C27637 VDD OR2X1_LOC_75/Y 0.21fF
C27638 OR2X1_LOC_214/B OR2X1_LOC_596/A 0.14fF
C27639 AND2X1_LOC_362/a_8_24# AND2X1_LOC_845/Y -0.00fF
C27640 AND2X1_LOC_817/a_8_24# OR2X1_LOC_847/B 0.01fF
C27641 OR2X1_LOC_743/A AND2X1_LOC_454/Y 0.01fF
C27642 OR2X1_LOC_691/A OR2X1_LOC_598/A 0.03fF
C27643 AND2X1_LOC_311/a_8_24# OR2X1_LOC_532/B 0.06fF
C27644 OR2X1_LOC_70/Y OR2X1_LOC_619/Y 0.10fF
C27645 OR2X1_LOC_273/Y AND2X1_LOC_274/a_8_24# 0.05fF
C27646 AND2X1_LOC_48/A OR2X1_LOC_637/A 0.04fF
C27647 OR2X1_LOC_40/Y D_INPUT_1 0.02fF
C27648 OR2X1_LOC_70/Y AND2X1_LOC_356/a_8_24# 0.01fF
C27649 OR2X1_LOC_689/Y AND2X1_LOC_691/a_8_24# 0.23fF
C27650 AND2X1_LOC_580/A AND2X1_LOC_719/a_8_24# 0.07fF
C27651 AND2X1_LOC_36/Y OR2X1_LOC_771/B 9.25fF
C27652 AND2X1_LOC_553/A OR2X1_LOC_22/Y 0.07fF
C27653 OR2X1_LOC_273/a_36_216# OR2X1_LOC_316/Y 0.00fF
C27654 AND2X1_LOC_728/Y AND2X1_LOC_797/A 0.18fF
C27655 GATE_366 OR2X1_LOC_89/A 0.01fF
C27656 AND2X1_LOC_31/Y AND2X1_LOC_44/Y 4.26fF
C27657 OR2X1_LOC_312/Y OR2X1_LOC_26/Y 0.03fF
C27658 OR2X1_LOC_40/Y OR2X1_LOC_173/a_8_216# 0.02fF
C27659 AND2X1_LOC_333/a_8_24# OR2X1_LOC_619/Y 0.06fF
C27660 AND2X1_LOC_342/a_8_24# OR2X1_LOC_485/A 0.02fF
C27661 OR2X1_LOC_158/A AND2X1_LOC_259/a_36_24# 0.00fF
C27662 OR2X1_LOC_119/a_36_216# AND2X1_LOC_573/A 0.01fF
C27663 OR2X1_LOC_427/A AND2X1_LOC_635/a_8_24# 0.01fF
C27664 OR2X1_LOC_599/A OR2X1_LOC_743/A 0.10fF
C27665 OR2X1_LOC_849/A AND2X1_LOC_3/Y 0.03fF
C27666 AND2X1_LOC_304/a_8_24# AND2X1_LOC_47/Y 0.01fF
C27667 OR2X1_LOC_217/Y AND2X1_LOC_122/a_8_24# 0.01fF
C27668 INPUT_0 OR2X1_LOC_416/a_8_216# 0.05fF
C27669 OR2X1_LOC_121/B OR2X1_LOC_161/A 0.99fF
C27670 OR2X1_LOC_233/a_8_216# OR2X1_LOC_753/A 0.03fF
C27671 OR2X1_LOC_146/Y AND2X1_LOC_663/A 0.05fF
C27672 OR2X1_LOC_600/A AND2X1_LOC_641/a_8_24# 0.02fF
C27673 AND2X1_LOC_36/Y OR2X1_LOC_776/A 0.06fF
C27674 AND2X1_LOC_365/A OR2X1_LOC_311/Y 0.15fF
C27675 AND2X1_LOC_395/a_8_24# OR2X1_LOC_401/B 0.01fF
C27676 AND2X1_LOC_395/a_36_24# OR2X1_LOC_401/A 0.00fF
C27677 AND2X1_LOC_139/A OR2X1_LOC_517/A 0.00fF
C27678 AND2X1_LOC_703/a_8_24# OR2X1_LOC_167/Y 0.23fF
C27679 AND2X1_LOC_17/Y OR2X1_LOC_636/B 0.03fF
C27680 OR2X1_LOC_377/A AND2X1_LOC_23/a_8_24# 0.05fF
C27681 AND2X1_LOC_59/Y OR2X1_LOC_649/a_8_216# 0.00fF
C27682 OR2X1_LOC_64/Y AND2X1_LOC_354/B 0.03fF
C27683 OR2X1_LOC_811/A AND2X1_LOC_47/Y 0.03fF
C27684 OR2X1_LOC_710/a_8_216# OR2X1_LOC_705/Y 0.01fF
C27685 AND2X1_LOC_831/Y AND2X1_LOC_841/B 0.01fF
C27686 OR2X1_LOC_462/B OR2X1_LOC_520/B 0.01fF
C27687 OR2X1_LOC_88/Y OR2X1_LOC_131/a_8_216# 0.00fF
C27688 OR2X1_LOC_449/B AND2X1_LOC_51/Y 0.09fF
C27689 OR2X1_LOC_256/A OR2X1_LOC_278/Y 0.03fF
C27690 OR2X1_LOC_577/Y OR2X1_LOC_367/a_8_216# 0.01fF
C27691 OR2X1_LOC_417/Y OR2X1_LOC_43/A 0.03fF
C27692 AND2X1_LOC_59/a_8_24# AND2X1_LOC_47/Y 0.01fF
C27693 AND2X1_LOC_715/A AND2X1_LOC_222/Y 0.02fF
C27694 AND2X1_LOC_702/Y AND2X1_LOC_727/A 0.37fF
C27695 OR2X1_LOC_36/Y AND2X1_LOC_465/Y 0.01fF
C27696 OR2X1_LOC_92/Y OR2X1_LOC_47/Y 3.24fF
C27697 OR2X1_LOC_311/Y OR2X1_LOC_43/A 0.17fF
C27698 OR2X1_LOC_810/A OR2X1_LOC_206/A 0.03fF
C27699 OR2X1_LOC_19/B OR2X1_LOC_836/B 0.26fF
C27700 AND2X1_LOC_41/A OR2X1_LOC_512/a_8_216# 0.01fF
C27701 AND2X1_LOC_831/a_8_24# INPUT_1 0.03fF
C27702 AND2X1_LOC_538/Y OR2X1_LOC_43/A 0.01fF
C27703 INPUT_1 OR2X1_LOC_44/Y 3.92fF
C27704 OR2X1_LOC_416/A OR2X1_LOC_39/A 0.00fF
C27705 OR2X1_LOC_636/A AND2X1_LOC_51/Y 0.01fF
C27706 AND2X1_LOC_808/A AND2X1_LOC_804/Y 0.24fF
C27707 OR2X1_LOC_294/a_8_216# OR2X1_LOC_598/A 0.01fF
C27708 OR2X1_LOC_316/Y OR2X1_LOC_75/a_36_216# 0.00fF
C27709 AND2X1_LOC_390/B OR2X1_LOC_64/Y 0.04fF
C27710 OR2X1_LOC_481/a_36_216# AND2X1_LOC_663/B 0.00fF
C27711 OR2X1_LOC_87/A OR2X1_LOC_544/A 0.03fF
C27712 OR2X1_LOC_78/B OR2X1_LOC_567/a_8_216# 0.06fF
C27713 OR2X1_LOC_553/B OR2X1_LOC_565/a_8_216# 0.39fF
C27714 AND2X1_LOC_738/B OR2X1_LOC_534/Y 0.08fF
C27715 AND2X1_LOC_811/a_8_24# AND2X1_LOC_811/Y 0.10fF
C27716 OR2X1_LOC_36/Y OR2X1_LOC_408/Y 0.03fF
C27717 OR2X1_LOC_599/A OR2X1_LOC_409/B 0.33fF
C27718 OR2X1_LOC_497/Y AND2X1_LOC_227/Y 0.11fF
C27719 OR2X1_LOC_707/B AND2X1_LOC_3/Y 0.06fF
C27720 OR2X1_LOC_271/B AND2X1_LOC_851/B 0.07fF
C27721 AND2X1_LOC_40/Y OR2X1_LOC_675/Y 0.00fF
C27722 OR2X1_LOC_71/Y OR2X1_LOC_7/A 0.06fF
C27723 OR2X1_LOC_6/B OR2X1_LOC_777/B 0.07fF
C27724 OR2X1_LOC_121/B AND2X1_LOC_51/Y 0.16fF
C27725 OR2X1_LOC_643/A AND2X1_LOC_106/a_8_24# 0.01fF
C27726 OR2X1_LOC_751/a_8_216# OR2X1_LOC_44/Y 0.01fF
C27727 AND2X1_LOC_92/Y AND2X1_LOC_406/a_8_24# 0.03fF
C27728 OR2X1_LOC_115/a_8_216# OR2X1_LOC_66/Y 0.01fF
C27729 OR2X1_LOC_624/B OR2X1_LOC_404/A 0.07fF
C27730 OR2X1_LOC_523/B OR2X1_LOC_523/a_8_216# 0.47fF
C27731 OR2X1_LOC_653/A OR2X1_LOC_112/B 0.26fF
C27732 OR2X1_LOC_43/A D_INPUT_3 0.05fF
C27733 AND2X1_LOC_101/a_8_24# OR2X1_LOC_64/Y 0.01fF
C27734 OR2X1_LOC_182/B OR2X1_LOC_182/a_8_216# 0.02fF
C27735 OR2X1_LOC_160/B OR2X1_LOC_544/B 0.14fF
C27736 AND2X1_LOC_399/a_8_24# AND2X1_LOC_813/a_8_24# 0.23fF
C27737 OR2X1_LOC_618/a_8_216# D_INPUT_1 0.01fF
C27738 AND2X1_LOC_231/Y OR2X1_LOC_171/Y 0.10fF
C27739 OR2X1_LOC_40/Y AND2X1_LOC_789/Y 0.06fF
C27740 AND2X1_LOC_59/Y OR2X1_LOC_493/Y 0.38fF
C27741 OR2X1_LOC_3/Y OR2X1_LOC_751/A 0.10fF
C27742 AND2X1_LOC_512/Y OR2X1_LOC_533/a_8_216# 0.02fF
C27743 OR2X1_LOC_597/a_8_216# OR2X1_LOC_536/a_8_216# 0.47fF
C27744 OR2X1_LOC_756/B OR2X1_LOC_367/B 0.04fF
C27745 OR2X1_LOC_45/B OR2X1_LOC_53/Y 0.03fF
C27746 OR2X1_LOC_259/a_8_216# OR2X1_LOC_259/B 0.06fF
C27747 OR2X1_LOC_848/A OR2X1_LOC_774/B 0.33fF
C27748 AND2X1_LOC_367/A OR2X1_LOC_437/A 0.45fF
C27749 OR2X1_LOC_375/A OR2X1_LOC_543/a_8_216# 0.01fF
C27750 OR2X1_LOC_185/A OR2X1_LOC_228/Y 0.07fF
C27751 OR2X1_LOC_680/A AND2X1_LOC_804/a_36_24# 0.01fF
C27752 OR2X1_LOC_64/Y AND2X1_LOC_863/Y 0.37fF
C27753 OR2X1_LOC_7/A AND2X1_LOC_770/a_36_24# 0.00fF
C27754 AND2X1_LOC_573/A OR2X1_LOC_88/Y 0.02fF
C27755 AND2X1_LOC_227/Y AND2X1_LOC_844/a_8_24# 0.01fF
C27756 OR2X1_LOC_243/a_8_216# OR2X1_LOC_62/B 0.01fF
C27757 OR2X1_LOC_715/B AND2X1_LOC_64/Y 0.07fF
C27758 OR2X1_LOC_19/B OR2X1_LOC_256/A 0.08fF
C27759 OR2X1_LOC_846/a_8_216# OR2X1_LOC_561/B 0.42fF
C27760 AND2X1_LOC_3/Y OR2X1_LOC_446/A 0.04fF
C27761 AND2X1_LOC_564/A AND2X1_LOC_220/a_8_24# 0.07fF
C27762 OR2X1_LOC_828/B OR2X1_LOC_198/A 0.25fF
C27763 OR2X1_LOC_32/a_8_216# OR2X1_LOC_598/A 0.06fF
C27764 OR2X1_LOC_848/A OR2X1_LOC_557/a_8_216# 0.02fF
C27765 AND2X1_LOC_370/a_8_24# AND2X1_LOC_182/A 0.00fF
C27766 OR2X1_LOC_375/A OR2X1_LOC_348/B 2.75fF
C27767 OR2X1_LOC_523/B OR2X1_LOC_576/A 0.10fF
C27768 AND2X1_LOC_32/a_8_24# OR2X1_LOC_68/B 0.01fF
C27769 AND2X1_LOC_726/Y VDD 0.21fF
C27770 OR2X1_LOC_12/Y OR2X1_LOC_603/Y 0.02fF
C27771 OR2X1_LOC_167/a_8_216# AND2X1_LOC_724/A 0.01fF
C27772 OR2X1_LOC_109/Y OR2X1_LOC_164/a_36_216# 0.01fF
C27773 AND2X1_LOC_574/Y AND2X1_LOC_501/Y 0.83fF
C27774 OR2X1_LOC_696/A AND2X1_LOC_364/Y 0.03fF
C27775 VDD OR2X1_LOC_828/Y 0.09fF
C27776 AND2X1_LOC_712/a_8_24# AND2X1_LOC_712/Y 0.00fF
C27777 OR2X1_LOC_348/Y OR2X1_LOC_362/a_8_216# 0.01fF
C27778 OR2X1_LOC_22/Y AND2X1_LOC_648/B 0.03fF
C27779 AND2X1_LOC_574/Y AND2X1_LOC_570/Y 0.01fF
C27780 OR2X1_LOC_113/a_8_216# OR2X1_LOC_160/B 0.02fF
C27781 OR2X1_LOC_753/A OR2X1_LOC_68/B 0.05fF
C27782 OR2X1_LOC_160/B OR2X1_LOC_474/B 0.05fF
C27783 AND2X1_LOC_392/A OR2X1_LOC_310/a_8_216# 0.03fF
C27784 AND2X1_LOC_575/a_8_24# AND2X1_LOC_501/a_8_24# 0.23fF
C27785 OR2X1_LOC_605/a_8_216# OR2X1_LOC_318/B 0.01fF
C27786 AND2X1_LOC_640/a_36_24# AND2X1_LOC_476/A 0.01fF
C27787 AND2X1_LOC_753/a_36_24# AND2X1_LOC_41/Y 0.00fF
C27788 AND2X1_LOC_12/Y OR2X1_LOC_349/B 0.22fF
C27789 OR2X1_LOC_19/B OR2X1_LOC_67/Y 0.01fF
C27790 OR2X1_LOC_31/Y AND2X1_LOC_476/A 0.14fF
C27791 AND2X1_LOC_11/Y AND2X1_LOC_36/Y 0.07fF
C27792 OR2X1_LOC_532/B OR2X1_LOC_84/A 0.01fF
C27793 OR2X1_LOC_58/Y OR2X1_LOC_12/Y 0.40fF
C27794 OR2X1_LOC_575/A OR2X1_LOC_500/a_36_216# 0.00fF
C27795 OR2X1_LOC_36/Y OR2X1_LOC_589/a_8_216# 0.19fF
C27796 OR2X1_LOC_599/A OR2X1_LOC_599/a_8_216# 0.00fF
C27797 OR2X1_LOC_709/A AND2X1_LOC_313/a_8_24# 0.04fF
C27798 OR2X1_LOC_561/a_8_216# OR2X1_LOC_561/A 0.39fF
C27799 OR2X1_LOC_147/a_8_216# OR2X1_LOC_705/a_8_216# 0.47fF
C27800 OR2X1_LOC_402/Y AND2X1_LOC_36/Y 0.04fF
C27801 VDD AND2X1_LOC_534/a_8_24# 0.00fF
C27802 OR2X1_LOC_158/A AND2X1_LOC_357/B 0.02fF
C27803 OR2X1_LOC_56/A AND2X1_LOC_785/Y 0.25fF
C27804 AND2X1_LOC_61/Y OR2X1_LOC_16/A 0.03fF
C27805 AND2X1_LOC_662/B AND2X1_LOC_269/a_8_24# 0.03fF
C27806 AND2X1_LOC_654/B OR2X1_LOC_171/Y 0.00fF
C27807 OR2X1_LOC_26/Y OR2X1_LOC_13/B 1.07fF
C27808 AND2X1_LOC_772/B OR2X1_LOC_595/A 0.02fF
C27809 AND2X1_LOC_70/Y OR2X1_LOC_856/A 0.06fF
C27810 AND2X1_LOC_91/B OR2X1_LOC_502/A 3.91fF
C27811 OR2X1_LOC_200/a_8_216# AND2X1_LOC_41/Y 0.01fF
C27812 OR2X1_LOC_158/A AND2X1_LOC_363/Y 0.35fF
C27813 OR2X1_LOC_269/B AND2X1_LOC_41/Y 0.03fF
C27814 OR2X1_LOC_70/A OR2X1_LOC_22/A 0.10fF
C27815 AND2X1_LOC_40/Y OR2X1_LOC_174/a_36_216# 0.00fF
C27816 AND2X1_LOC_456/Y OR2X1_LOC_437/A 0.00fF
C27817 AND2X1_LOC_110/Y OR2X1_LOC_302/A 0.01fF
C27818 AND2X1_LOC_323/a_8_24# AND2X1_LOC_299/a_8_24# 0.23fF
C27819 AND2X1_LOC_512/Y OR2X1_LOC_428/A 0.07fF
C27820 AND2X1_LOC_349/B OR2X1_LOC_13/B 0.17fF
C27821 OR2X1_LOC_89/A OR2X1_LOC_13/B 0.31fF
C27822 AND2X1_LOC_719/Y OR2X1_LOC_51/Y 0.03fF
C27823 OR2X1_LOC_151/A OR2X1_LOC_809/B 0.06fF
C27824 OR2X1_LOC_74/A OR2X1_LOC_437/A 1.35fF
C27825 AND2X1_LOC_547/Y AND2X1_LOC_550/a_8_24# 0.03fF
C27826 AND2X1_LOC_65/A OR2X1_LOC_78/B 0.17fF
C27827 VDD AND2X1_LOC_110/Y 0.39fF
C27828 OR2X1_LOC_40/Y OR2X1_LOC_426/B 0.67fF
C27829 OR2X1_LOC_440/B OR2X1_LOC_66/A 0.03fF
C27830 AND2X1_LOC_91/B OR2X1_LOC_571/B 0.02fF
C27831 OR2X1_LOC_857/B OR2X1_LOC_634/A 0.03fF
C27832 OR2X1_LOC_323/A OR2X1_LOC_315/Y 0.04fF
C27833 OR2X1_LOC_110/a_36_216# OR2X1_LOC_316/Y 0.00fF
C27834 OR2X1_LOC_185/A OR2X1_LOC_562/A 0.01fF
C27835 OR2X1_LOC_516/Y OR2X1_LOC_36/Y 0.03fF
C27836 OR2X1_LOC_405/A OR2X1_LOC_390/a_8_216# -0.00fF
C27837 AND2X1_LOC_43/B OR2X1_LOC_140/B 0.00fF
C27838 AND2X1_LOC_70/Y AND2X1_LOC_313/a_8_24# 0.09fF
C27839 OR2X1_LOC_348/Y OR2X1_LOC_363/B 0.12fF
C27840 OR2X1_LOC_499/B OR2X1_LOC_549/A 0.02fF
C27841 OR2X1_LOC_510/A OR2X1_LOC_78/B 0.01fF
C27842 OR2X1_LOC_653/B AND2X1_LOC_40/Y 0.01fF
C27843 AND2X1_LOC_76/Y OR2X1_LOC_522/a_8_216# 0.01fF
C27844 INPUT_5 OR2X1_LOC_158/A 0.03fF
C27845 AND2X1_LOC_91/B OR2X1_LOC_400/A 0.01fF
C27846 OR2X1_LOC_136/Y AND2X1_LOC_655/A 0.23fF
C27847 OR2X1_LOC_160/B OR2X1_LOC_658/a_8_216# 0.02fF
C27848 AND2X1_LOC_12/Y OR2X1_LOC_97/A 0.06fF
C27849 AND2X1_LOC_423/a_8_24# OR2X1_LOC_596/A 0.01fF
C27850 AND2X1_LOC_286/a_8_24# OR2X1_LOC_59/Y 0.01fF
C27851 OR2X1_LOC_160/B OR2X1_LOC_78/Y 0.05fF
C27852 OR2X1_LOC_8/Y OR2X1_LOC_91/A 0.03fF
C27853 OR2X1_LOC_624/Y OR2X1_LOC_66/A 0.00fF
C27854 OR2X1_LOC_146/a_8_216# OR2X1_LOC_599/A 0.01fF
C27855 OR2X1_LOC_426/A OR2X1_LOC_765/a_36_216# 0.00fF
C27856 OR2X1_LOC_160/B OR2X1_LOC_274/a_8_216# 0.03fF
C27857 OR2X1_LOC_337/A AND2X1_LOC_95/Y 0.15fF
C27858 OR2X1_LOC_348/Y OR2X1_LOC_756/B 0.30fF
C27859 AND2X1_LOC_675/Y AND2X1_LOC_657/Y 0.18fF
C27860 AND2X1_LOC_176/a_8_24# OR2X1_LOC_180/B 0.09fF
C27861 OR2X1_LOC_316/a_36_216# OR2X1_LOC_52/B 0.02fF
C27862 OR2X1_LOC_160/A OR2X1_LOC_318/A 0.11fF
C27863 AND2X1_LOC_64/Y AND2X1_LOC_81/a_8_24# 0.02fF
C27864 OR2X1_LOC_349/a_8_216# OR2X1_LOC_756/B 0.02fF
C27865 OR2X1_LOC_194/Y AND2X1_LOC_7/B 2.99fF
C27866 AND2X1_LOC_723/Y VDD 0.52fF
C27867 OR2X1_LOC_338/a_8_216# AND2X1_LOC_95/Y 0.01fF
C27868 AND2X1_LOC_92/Y OR2X1_LOC_630/B 0.01fF
C27869 OR2X1_LOC_160/B AND2X1_LOC_424/a_8_24# 0.01fF
C27870 OR2X1_LOC_751/Y VDD 0.06fF
C27871 AND2X1_LOC_658/B AND2X1_LOC_862/Y 0.06fF
C27872 AND2X1_LOC_22/Y AND2X1_LOC_26/a_8_24# 0.02fF
C27873 AND2X1_LOC_732/B OR2X1_LOC_92/Y 0.01fF
C27874 AND2X1_LOC_705/Y OR2X1_LOC_39/A 0.12fF
C27875 OR2X1_LOC_154/A AND2X1_LOC_60/a_36_24# 0.00fF
C27876 AND2X1_LOC_84/Y AND2X1_LOC_84/a_8_24# 0.01fF
C27877 AND2X1_LOC_720/Y OR2X1_LOC_494/Y 0.01fF
C27878 OR2X1_LOC_805/A OR2X1_LOC_294/Y 0.03fF
C27879 AND2X1_LOC_12/Y D_GATE_662 0.02fF
C27880 AND2X1_LOC_365/a_8_24# OR2X1_LOC_91/A 0.04fF
C27881 AND2X1_LOC_22/Y OR2X1_LOC_269/B 0.18fF
C27882 OR2X1_LOC_457/a_8_216# OR2X1_LOC_161/B 0.05fF
C27883 OR2X1_LOC_160/A OR2X1_LOC_151/A 0.70fF
C27884 OR2X1_LOC_375/A AND2X1_LOC_65/A 0.07fF
C27885 OR2X1_LOC_516/B AND2X1_LOC_469/B 0.02fF
C27886 OR2X1_LOC_179/a_8_216# OR2X1_LOC_329/B 0.03fF
C27887 OR2X1_LOC_154/A OR2X1_LOC_663/a_8_216# 0.03fF
C27888 OR2X1_LOC_280/Y AND2X1_LOC_465/A 0.07fF
C27889 OR2X1_LOC_864/A AND2X1_LOC_44/Y 0.06fF
C27890 OR2X1_LOC_529/Y AND2X1_LOC_242/B 0.03fF
C27891 OR2X1_LOC_364/A OR2X1_LOC_390/A 0.14fF
C27892 AND2X1_LOC_552/a_36_24# OR2X1_LOC_280/Y 0.01fF
C27893 OR2X1_LOC_139/A OR2X1_LOC_141/B 0.01fF
C27894 AND2X1_LOC_3/Y OR2X1_LOC_572/a_8_216# 0.05fF
C27895 AND2X1_LOC_47/Y OR2X1_LOC_777/B 0.06fF
C27896 OR2X1_LOC_682/Y OR2X1_LOC_428/A 0.04fF
C27897 AND2X1_LOC_852/Y OR2X1_LOC_16/A 0.06fF
C27898 OR2X1_LOC_240/A AND2X1_LOC_44/Y 0.08fF
C27899 AND2X1_LOC_3/Y OR2X1_LOC_721/a_8_216# 0.05fF
C27900 OR2X1_LOC_474/Y OR2X1_LOC_624/a_8_216# 0.39fF
C27901 AND2X1_LOC_40/a_36_24# AND2X1_LOC_25/Y 0.01fF
C27902 OR2X1_LOC_510/A OR2X1_LOC_375/A 0.02fF
C27903 OR2X1_LOC_633/B AND2X1_LOC_44/Y 0.05fF
C27904 OR2X1_LOC_8/Y AND2X1_LOC_62/a_36_24# 0.00fF
C27905 AND2X1_LOC_658/B OR2X1_LOC_619/Y 0.01fF
C27906 OR2X1_LOC_223/A OR2X1_LOC_303/B 0.04fF
C27907 OR2X1_LOC_805/A OR2X1_LOC_733/A 0.03fF
C27908 OR2X1_LOC_620/Y OR2X1_LOC_78/A 0.07fF
C27909 OR2X1_LOC_533/Y AND2X1_LOC_645/A 0.11fF
C27910 AND2X1_LOC_714/a_8_24# OR2X1_LOC_7/A 0.02fF
C27911 OR2X1_LOC_201/Y AND2X1_LOC_7/B 0.02fF
C27912 OR2X1_LOC_249/a_8_216# OR2X1_LOC_244/Y 0.01fF
C27913 AND2X1_LOC_387/B OR2X1_LOC_691/Y 0.03fF
C27914 OR2X1_LOC_501/B OR2X1_LOC_629/Y 0.01fF
C27915 OR2X1_LOC_485/Y OR2X1_LOC_511/Y 0.03fF
C27916 AND2X1_LOC_354/Y AND2X1_LOC_434/Y 0.01fF
C27917 AND2X1_LOC_570/Y AND2X1_LOC_621/Y 0.03fF
C27918 AND2X1_LOC_729/Y AND2X1_LOC_724/Y 0.00fF
C27919 OR2X1_LOC_851/a_8_216# AND2X1_LOC_43/B 0.02fF
C27920 OR2X1_LOC_3/Y OR2X1_LOC_118/a_8_216# 0.01fF
C27921 OR2X1_LOC_502/A AND2X1_LOC_819/a_36_24# 0.01fF
C27922 AND2X1_LOC_76/Y OR2X1_LOC_91/A 0.03fF
C27923 OR2X1_LOC_51/Y OR2X1_LOC_252/Y 0.55fF
C27924 OR2X1_LOC_485/A OR2X1_LOC_12/Y 1.28fF
C27925 VDD OR2X1_LOC_664/Y 0.22fF
C27926 OR2X1_LOC_473/Y OR2X1_LOC_392/B 0.38fF
C27927 OR2X1_LOC_329/a_8_216# OR2X1_LOC_585/A 0.01fF
C27928 OR2X1_LOC_51/Y OR2X1_LOC_313/Y 0.03fF
C27929 OR2X1_LOC_287/B OR2X1_LOC_343/a_8_216# 0.00fF
C27930 OR2X1_LOC_843/a_36_216# OR2X1_LOC_843/B 0.00fF
C27931 AND2X1_LOC_40/Y OR2X1_LOC_808/B 0.05fF
C27932 AND2X1_LOC_552/A OR2X1_LOC_312/Y 0.01fF
C27933 AND2X1_LOC_27/a_8_24# OR2X1_LOC_338/A 0.25fF
C27934 OR2X1_LOC_604/A OR2X1_LOC_699/a_36_216# 0.01fF
C27935 OR2X1_LOC_660/Y OR2X1_LOC_185/A 0.03fF
C27936 OR2X1_LOC_296/Y OR2X1_LOC_294/Y 0.04fF
C27937 OR2X1_LOC_670/a_36_216# OR2X1_LOC_96/Y 0.00fF
C27938 OR2X1_LOC_532/B OR2X1_LOC_354/a_36_216# 0.00fF
C27939 OR2X1_LOC_687/Y OR2X1_LOC_687/A 0.18fF
C27940 OR2X1_LOC_309/a_8_216# AND2X1_LOC_211/B 0.04fF
C27941 AND2X1_LOC_571/a_8_24# OR2X1_LOC_64/Y 0.17fF
C27942 AND2X1_LOC_572/A OR2X1_LOC_56/A 0.03fF
C27943 AND2X1_LOC_522/a_8_24# OR2X1_LOC_404/Y 0.01fF
C27944 AND2X1_LOC_860/a_8_24# OR2X1_LOC_18/Y 0.02fF
C27945 OR2X1_LOC_99/a_8_216# OR2X1_LOC_66/A 0.01fF
C27946 AND2X1_LOC_141/B OR2X1_LOC_595/A 0.01fF
C27947 VDD OR2X1_LOC_601/Y 0.18fF
C27948 OR2X1_LOC_744/A OR2X1_LOC_11/Y 0.11fF
C27949 OR2X1_LOC_154/A OR2X1_LOC_78/A 0.20fF
C27950 OR2X1_LOC_108/a_8_216# OR2X1_LOC_7/A 0.01fF
C27951 AND2X1_LOC_31/a_8_24# AND2X1_LOC_44/Y 0.02fF
C27952 OR2X1_LOC_810/A OR2X1_LOC_776/Y 0.07fF
C27953 AND2X1_LOC_712/B OR2X1_LOC_428/A 0.01fF
C27954 AND2X1_LOC_500/a_8_24# OR2X1_LOC_51/Y 0.07fF
C27955 OR2X1_LOC_121/a_8_216# OR2X1_LOC_121/B 0.07fF
C27956 OR2X1_LOC_812/B OR2X1_LOC_862/A 0.14fF
C27957 AND2X1_LOC_12/Y OR2X1_LOC_858/B 0.05fF
C27958 OR2X1_LOC_669/A OR2X1_LOC_59/Y 0.19fF
C27959 OR2X1_LOC_710/B OR2X1_LOC_710/a_8_216# 0.05fF
C27960 OR2X1_LOC_54/Y OR2X1_LOC_428/A 0.14fF
C27961 OR2X1_LOC_416/Y AND2X1_LOC_786/Y 0.15fF
C27962 OR2X1_LOC_625/Y OR2X1_LOC_92/Y 0.00fF
C27963 OR2X1_LOC_40/Y OR2X1_LOC_743/A 0.03fF
C27964 AND2X1_LOC_41/A OR2X1_LOC_130/A 0.21fF
C27965 AND2X1_LOC_537/a_8_24# OR2X1_LOC_385/Y 0.05fF
C27966 OR2X1_LOC_756/B OR2X1_LOC_456/Y 0.01fF
C27967 OR2X1_LOC_51/B INPUT_6 0.49fF
C27968 AND2X1_LOC_560/B OR2X1_LOC_744/A 0.07fF
C27969 OR2X1_LOC_193/A OR2X1_LOC_596/A 0.19fF
C27970 OR2X1_LOC_62/B OR2X1_LOC_576/A 1.11fF
C27971 AND2X1_LOC_47/Y OR2X1_LOC_831/B 5.64fF
C27972 OR2X1_LOC_777/B OR2X1_LOC_598/A 0.07fF
C27973 OR2X1_LOC_132/Y AND2X1_LOC_361/A 0.02fF
C27974 AND2X1_LOC_8/Y OR2X1_LOC_520/a_8_216# 0.01fF
C27975 OR2X1_LOC_154/A OR2X1_LOC_458/B 0.03fF
C27976 AND2X1_LOC_296/a_36_24# OR2X1_LOC_44/Y 0.01fF
C27977 OR2X1_LOC_696/A OR2X1_LOC_619/a_8_216# 0.01fF
C27978 OR2X1_LOC_426/B OR2X1_LOC_7/A 0.14fF
C27979 AND2X1_LOC_12/Y OR2X1_LOC_475/B 0.03fF
C27980 OR2X1_LOC_724/A AND2X1_LOC_419/a_8_24# 0.02fF
C27981 OR2X1_LOC_175/B OR2X1_LOC_624/A 0.01fF
C27982 OR2X1_LOC_45/B INPUT_1 1.11fF
C27983 OR2X1_LOC_337/a_8_216# OR2X1_LOC_87/A 0.04fF
C27984 VDD AND2X1_LOC_78/a_8_24# -0.00fF
C27985 OR2X1_LOC_190/B OR2X1_LOC_553/A 0.17fF
C27986 AND2X1_LOC_367/A AND2X1_LOC_348/Y 0.08fF
C27987 AND2X1_LOC_715/A OR2X1_LOC_74/A 0.14fF
C27988 AND2X1_LOC_59/Y OR2X1_LOC_61/B 0.14fF
C27989 AND2X1_LOC_720/a_36_24# OR2X1_LOC_427/A 0.01fF
C27990 AND2X1_LOC_840/a_8_24# OR2X1_LOC_39/A 0.03fF
C27991 OR2X1_LOC_856/B OR2X1_LOC_161/A 1.55fF
C27992 OR2X1_LOC_91/A OR2X1_LOC_52/B 0.10fF
C27993 OR2X1_LOC_533/Y AND2X1_LOC_477/A 0.03fF
C27994 VDD OR2X1_LOC_754/A 0.05fF
C27995 OR2X1_LOC_49/A D_INPUT_0 0.14fF
C27996 OR2X1_LOC_187/Y AND2X1_LOC_866/A 0.08fF
C27997 AND2X1_LOC_367/A OR2X1_LOC_753/A 0.11fF
C27998 OR2X1_LOC_18/Y OR2X1_LOC_71/a_8_216# 0.01fF
C27999 OR2X1_LOC_715/B OR2X1_LOC_206/A 0.05fF
C28000 OR2X1_LOC_309/Y OR2X1_LOC_64/Y 0.03fF
C28001 AND2X1_LOC_477/A AND2X1_LOC_212/Y 0.01fF
C28002 VDD OR2X1_LOC_275/A 0.00fF
C28003 AND2X1_LOC_841/B AND2X1_LOC_436/B 0.19fF
C28004 OR2X1_LOC_3/Y OR2X1_LOC_56/A 1.64fF
C28005 OR2X1_LOC_158/A AND2X1_LOC_116/B 0.02fF
C28006 OR2X1_LOC_201/a_8_216# AND2X1_LOC_7/B 0.01fF
C28007 AND2X1_LOC_95/Y OR2X1_LOC_347/B 0.20fF
C28008 OR2X1_LOC_756/B OR2X1_LOC_810/A 0.08fF
C28009 OR2X1_LOC_516/Y OR2X1_LOC_419/Y 0.06fF
C28010 AND2X1_LOC_344/a_8_24# AND2X1_LOC_359/B 0.01fF
C28011 AND2X1_LOC_776/a_8_24# OR2X1_LOC_527/Y 0.01fF
C28012 AND2X1_LOC_191/B OR2X1_LOC_279/Y 0.07fF
C28013 AND2X1_LOC_95/Y OR2X1_LOC_539/Y 0.68fF
C28014 OR2X1_LOC_181/B OR2X1_LOC_375/A 0.03fF
C28015 OR2X1_LOC_691/a_8_216# OR2X1_LOC_532/B 0.01fF
C28016 AND2X1_LOC_631/Y OR2X1_LOC_56/A 0.03fF
C28017 OR2X1_LOC_40/Y OR2X1_LOC_125/Y 0.02fF
C28018 INPUT_1 OR2X1_LOC_382/A 0.05fF
C28019 OR2X1_LOC_31/Y OR2X1_LOC_766/a_8_216# 0.01fF
C28020 OR2X1_LOC_653/Y OR2X1_LOC_87/A 0.00fF
C28021 OR2X1_LOC_778/A OR2X1_LOC_78/A 0.02fF
C28022 OR2X1_LOC_40/Y OR2X1_LOC_246/A 0.01fF
C28023 OR2X1_LOC_656/B OR2X1_LOC_520/Y 0.56fF
C28024 D_INPUT_0 OR2X1_LOC_596/A 0.02fF
C28025 AND2X1_LOC_50/Y AND2X1_LOC_64/a_36_24# 0.01fF
C28026 OR2X1_LOC_756/B AND2X1_LOC_589/a_8_24# 0.01fF
C28027 AND2X1_LOC_350/Y OR2X1_LOC_51/Y 0.04fF
C28028 AND2X1_LOC_802/a_8_24# AND2X1_LOC_436/Y 0.00fF
C28029 OR2X1_LOC_662/A OR2X1_LOC_130/A 0.49fF
C28030 AND2X1_LOC_12/Y AND2X1_LOC_282/a_8_24# 0.01fF
C28031 OR2X1_LOC_637/A AND2X1_LOC_3/Y 0.01fF
C28032 OR2X1_LOC_589/A AND2X1_LOC_831/Y 0.50fF
C28033 OR2X1_LOC_517/A AND2X1_LOC_116/Y 0.03fF
C28034 AND2X1_LOC_276/Y OR2X1_LOC_275/Y 0.01fF
C28035 OR2X1_LOC_545/A AND2X1_LOC_47/Y 0.01fF
C28036 OR2X1_LOC_264/Y AND2X1_LOC_3/Y 0.30fF
C28037 OR2X1_LOC_40/Y OR2X1_LOC_225/a_8_216# 0.01fF
C28038 AND2X1_LOC_717/a_8_24# OR2X1_LOC_372/Y 0.01fF
C28039 OR2X1_LOC_744/A OR2X1_LOC_64/Y 0.37fF
C28040 OR2X1_LOC_599/A AND2X1_LOC_676/a_8_24# 0.04fF
C28041 OR2X1_LOC_620/Y OR2X1_LOC_155/A 0.07fF
C28042 OR2X1_LOC_290/a_8_216# OR2X1_LOC_27/a_8_216# 0.47fF
C28043 OR2X1_LOC_377/A AND2X1_LOC_823/a_8_24# 0.02fF
C28044 OR2X1_LOC_309/Y OR2X1_LOC_417/A 0.19fF
C28045 OR2X1_LOC_510/Y OR2X1_LOC_657/a_8_216# 0.01fF
C28046 OR2X1_LOC_692/Y OR2X1_LOC_47/Y 0.01fF
C28047 AND2X1_LOC_858/a_8_24# AND2X1_LOC_806/A 0.01fF
C28048 OR2X1_LOC_158/A OR2X1_LOC_96/a_8_216# 0.01fF
C28049 AND2X1_LOC_624/A OR2X1_LOC_44/Y 0.03fF
C28050 OR2X1_LOC_484/a_36_216# AND2X1_LOC_727/A 0.00fF
C28051 OR2X1_LOC_756/B AND2X1_LOC_281/a_36_24# 0.00fF
C28052 OR2X1_LOC_317/a_8_216# AND2X1_LOC_51/Y 0.01fF
C28053 AND2X1_LOC_387/a_36_24# D_INPUT_0 0.00fF
C28054 OR2X1_LOC_85/A AND2X1_LOC_266/Y 0.18fF
C28055 OR2X1_LOC_427/A OR2X1_LOC_418/a_8_216# 0.01fF
C28056 OR2X1_LOC_40/Y OR2X1_LOC_409/B 0.02fF
C28057 AND2X1_LOC_729/a_8_24# OR2X1_LOC_47/Y 0.01fF
C28058 OR2X1_LOC_291/a_8_216# OR2X1_LOC_278/a_8_216# 0.47fF
C28059 OR2X1_LOC_380/A OR2X1_LOC_44/Y 0.03fF
C28060 OR2X1_LOC_267/a_8_216# OR2X1_LOC_204/Y 0.01fF
C28061 AND2X1_LOC_647/B OR2X1_LOC_16/A 0.03fF
C28062 OR2X1_LOC_287/B OR2X1_LOC_249/Y 0.02fF
C28063 AND2X1_LOC_35/Y OR2X1_LOC_753/A 0.10fF
C28064 AND2X1_LOC_795/Y OR2X1_LOC_373/Y 0.08fF
C28065 OR2X1_LOC_308/A OR2X1_LOC_779/B 0.00fF
C28066 AND2X1_LOC_489/Y AND2X1_LOC_573/A 0.02fF
C28067 OR2X1_LOC_644/B AND2X1_LOC_56/B 0.00fF
C28068 AND2X1_LOC_41/A OR2X1_LOC_62/B 0.01fF
C28069 OR2X1_LOC_774/Y OR2X1_LOC_848/a_8_216# 0.01fF
C28070 OR2X1_LOC_175/Y OR2X1_LOC_854/A 0.06fF
C28071 OR2X1_LOC_154/A OR2X1_LOC_155/A 0.24fF
C28072 OR2X1_LOC_131/Y OR2X1_LOC_118/Y 0.01fF
C28073 OR2X1_LOC_856/B AND2X1_LOC_51/Y 0.07fF
C28074 AND2X1_LOC_301/a_8_24# AND2X1_LOC_476/A 0.04fF
C28075 OR2X1_LOC_744/A OR2X1_LOC_417/A 4.19fF
C28076 AND2X1_LOC_76/Y AND2X1_LOC_662/a_8_24# 0.01fF
C28077 OR2X1_LOC_227/B OR2X1_LOC_641/B 0.00fF
C28078 OR2X1_LOC_714/a_36_216# OR2X1_LOC_317/B 0.00fF
C28079 AND2X1_LOC_44/Y OR2X1_LOC_608/Y 0.07fF
C28080 OR2X1_LOC_415/Y OR2X1_LOC_80/A 0.04fF
C28081 OR2X1_LOC_280/Y OR2X1_LOC_237/Y 0.72fF
C28082 OR2X1_LOC_243/A AND2X1_LOC_42/B 0.00fF
C28083 AND2X1_LOC_80/a_36_24# OR2X1_LOC_646/A 0.00fF
C28084 AND2X1_LOC_191/Y OR2X1_LOC_613/a_8_216# 0.03fF
C28085 AND2X1_LOC_222/Y OR2X1_LOC_310/a_36_216# 0.00fF
C28086 OR2X1_LOC_501/A OR2X1_LOC_501/a_8_216# 0.39fF
C28087 AND2X1_LOC_367/A AND2X1_LOC_845/Y 0.10fF
C28088 OR2X1_LOC_646/A OR2X1_LOC_87/A 0.03fF
C28089 OR2X1_LOC_600/A OR2X1_LOC_47/Y 0.22fF
C28090 AND2X1_LOC_367/a_8_24# OR2X1_LOC_7/A 0.01fF
C28091 OR2X1_LOC_158/A AND2X1_LOC_204/Y 0.00fF
C28092 INPUT_0 OR2X1_LOC_31/Y 2.10fF
C28093 OR2X1_LOC_744/A OR2X1_LOC_64/a_8_216# 0.01fF
C28094 OR2X1_LOC_403/A OR2X1_LOC_403/a_8_216# 0.39fF
C28095 AND2X1_LOC_17/Y AND2X1_LOC_51/A 0.73fF
C28096 AND2X1_LOC_36/Y OR2X1_LOC_593/B 0.00fF
C28097 OR2X1_LOC_185/A OR2X1_LOC_76/A 0.03fF
C28098 OR2X1_LOC_643/A AND2X1_LOC_3/Y 0.06fF
C28099 AND2X1_LOC_393/a_8_24# OR2X1_LOC_557/A 0.01fF
C28100 OR2X1_LOC_3/Y AND2X1_LOC_56/B 0.03fF
C28101 OR2X1_LOC_166/a_8_216# OR2X1_LOC_47/Y 0.03fF
C28102 AND2X1_LOC_3/Y OR2X1_LOC_124/Y 0.06fF
C28103 AND2X1_LOC_523/a_8_24# OR2X1_LOC_22/Y 0.03fF
C28104 OR2X1_LOC_653/Y OR2X1_LOC_648/a_8_216# 0.03fF
C28105 OR2X1_LOC_74/A OR2X1_LOC_753/A 0.03fF
C28106 OR2X1_LOC_51/Y AND2X1_LOC_687/a_36_24# 0.00fF
C28107 OR2X1_LOC_472/A AND2X1_LOC_3/Y 0.09fF
C28108 OR2X1_LOC_481/A OR2X1_LOC_236/a_8_216# 0.01fF
C28109 AND2X1_LOC_778/a_8_24# OR2X1_LOC_371/Y -0.00fF
C28110 AND2X1_LOC_855/a_36_24# AND2X1_LOC_655/A 0.08fF
C28111 OR2X1_LOC_676/Y OR2X1_LOC_194/a_36_216# 0.01fF
C28112 AND2X1_LOC_6/a_8_24# OR2X1_LOC_78/A 0.04fF
C28113 AND2X1_LOC_47/Y OR2X1_LOC_575/A 0.05fF
C28114 OR2X1_LOC_831/a_8_216# OR2X1_LOC_121/B 0.01fF
C28115 OR2X1_LOC_743/A OR2X1_LOC_7/A 0.16fF
C28116 AND2X1_LOC_113/a_8_24# OR2X1_LOC_95/Y 0.01fF
C28117 AND2X1_LOC_717/Y OR2X1_LOC_31/Y 0.03fF
C28118 OR2X1_LOC_287/B OR2X1_LOC_402/a_8_216# 0.01fF
C28119 OR2X1_LOC_64/Y AND2X1_LOC_840/B 0.12fF
C28120 OR2X1_LOC_316/Y OR2X1_LOC_268/a_36_216# 0.00fF
C28121 OR2X1_LOC_70/Y AND2X1_LOC_454/A 0.01fF
C28122 OR2X1_LOC_216/Y OR2X1_LOC_121/B 0.01fF
C28123 OR2X1_LOC_647/A OR2X1_LOC_647/B 0.25fF
C28124 OR2X1_LOC_816/Y AND2X1_LOC_793/Y 0.00fF
C28125 AND2X1_LOC_662/a_8_24# OR2X1_LOC_52/B 0.04fF
C28126 AND2X1_LOC_273/a_8_24# AND2X1_LOC_36/Y 0.03fF
C28127 OR2X1_LOC_74/A AND2X1_LOC_243/a_8_24# 0.01fF
C28128 OR2X1_LOC_51/Y OR2X1_LOC_331/a_8_216# 0.01fF
C28129 OR2X1_LOC_99/A OR2X1_LOC_78/A 0.03fF
C28130 OR2X1_LOC_19/B OR2X1_LOC_248/Y 0.02fF
C28131 OR2X1_LOC_185/A OR2X1_LOC_436/Y 0.03fF
C28132 AND2X1_LOC_101/B AND2X1_LOC_101/a_8_24# 0.01fF
C28133 OR2X1_LOC_516/a_8_216# OR2X1_LOC_442/a_8_216# 0.47fF
C28134 OR2X1_LOC_426/A OR2X1_LOC_430/Y 0.01fF
C28135 OR2X1_LOC_652/a_8_216# AND2X1_LOC_47/Y 0.05fF
C28136 OR2X1_LOC_631/B OR2X1_LOC_62/B 0.00fF
C28137 AND2X1_LOC_842/a_8_24# OR2X1_LOC_419/Y 0.01fF
C28138 AND2X1_LOC_133/a_8_24# AND2X1_LOC_8/Y 0.05fF
C28139 OR2X1_LOC_31/Y OR2X1_LOC_11/Y 0.20fF
C28140 OR2X1_LOC_87/B D_INPUT_0 0.00fF
C28141 OR2X1_LOC_121/B OR2X1_LOC_787/Y 0.25fF
C28142 AND2X1_LOC_56/B AND2X1_LOC_53/Y 0.00fF
C28143 OR2X1_LOC_835/B AND2X1_LOC_821/a_8_24# 0.01fF
C28144 OR2X1_LOC_61/Y OR2X1_LOC_215/a_8_216# 0.04fF
C28145 OR2X1_LOC_47/Y OR2X1_LOC_619/Y 0.22fF
C28146 OR2X1_LOC_78/A OR2X1_LOC_560/A 0.09fF
C28147 AND2X1_LOC_39/a_8_24# AND2X1_LOC_699/a_8_24# 0.23fF
C28148 OR2X1_LOC_59/Y OR2X1_LOC_534/a_8_216# 0.01fF
C28149 AND2X1_LOC_18/Y OR2X1_LOC_71/A 0.02fF
C28150 AND2X1_LOC_663/B AND2X1_LOC_260/a_8_24# 0.07fF
C28151 OR2X1_LOC_833/Y OR2X1_LOC_723/B 0.07fF
C28152 AND2X1_LOC_256/a_8_24# AND2X1_LOC_36/Y 0.01fF
C28153 OR2X1_LOC_43/A AND2X1_LOC_831/Y 0.03fF
C28154 OR2X1_LOC_180/a_8_216# OR2X1_LOC_544/B 0.47fF
C28155 OR2X1_LOC_633/B OR2X1_LOC_720/B 0.08fF
C28156 OR2X1_LOC_333/B OR2X1_LOC_814/A 0.01fF
C28157 AND2X1_LOC_860/A OR2X1_LOC_437/A 0.14fF
C28158 OR2X1_LOC_151/A OR2X1_LOC_532/Y 0.03fF
C28159 OR2X1_LOC_575/A OR2X1_LOC_598/A 0.00fF
C28160 OR2X1_LOC_859/A AND2X1_LOC_42/B 0.01fF
C28161 OR2X1_LOC_31/Y OR2X1_LOC_690/A 0.13fF
C28162 OR2X1_LOC_850/A OR2X1_LOC_814/A 0.06fF
C28163 OR2X1_LOC_220/A OR2X1_LOC_740/a_8_216# 0.06fF
C28164 OR2X1_LOC_373/Y AND2X1_LOC_439/a_8_24# 0.24fF
C28165 AND2X1_LOC_44/Y OR2X1_LOC_501/A 0.01fF
C28166 OR2X1_LOC_485/A AND2X1_LOC_801/B 0.01fF
C28167 AND2X1_LOC_326/A AND2X1_LOC_863/A 0.09fF
C28168 AND2X1_LOC_56/B OR2X1_LOC_223/A 0.03fF
C28169 VDD OR2X1_LOC_550/B 0.09fF
C28170 D_INPUT_0 OR2X1_LOC_33/B 0.01fF
C28171 INPUT_4 OR2X1_LOC_430/Y 0.01fF
C28172 AND2X1_LOC_322/a_8_24# OR2X1_LOC_532/Y 0.01fF
C28173 OR2X1_LOC_516/Y OR2X1_LOC_177/Y 0.03fF
C28174 OR2X1_LOC_22/Y AND2X1_LOC_853/a_36_24# 0.00fF
C28175 AND2X1_LOC_8/Y OR2X1_LOC_673/A 0.75fF
C28176 AND2X1_LOC_102/a_8_24# AND2X1_LOC_672/a_8_24# 0.23fF
C28177 OR2X1_LOC_272/a_8_216# OR2X1_LOC_31/Y 0.07fF
C28178 AND2X1_LOC_621/Y OR2X1_LOC_406/A 0.07fF
C28179 OR2X1_LOC_760/a_36_216# OR2X1_LOC_585/A 0.00fF
C28180 AND2X1_LOC_573/A AND2X1_LOC_216/A 0.01fF
C28181 OR2X1_LOC_840/A OR2X1_LOC_724/A 0.10fF
C28182 OR2X1_LOC_427/A AND2X1_LOC_779/Y 0.04fF
C28183 VDD OR2X1_LOC_142/Y 0.53fF
C28184 OR2X1_LOC_66/A OR2X1_LOC_174/Y 0.03fF
C28185 AND2X1_LOC_70/Y OR2X1_LOC_537/a_8_216# 0.06fF
C28186 OR2X1_LOC_375/A OR2X1_LOC_98/a_36_216# 0.02fF
C28187 AND2X1_LOC_84/Y OR2X1_LOC_79/Y 0.42fF
C28188 AND2X1_LOC_192/Y AND2X1_LOC_782/a_8_24# 0.10fF
C28189 OR2X1_LOC_473/Y OR2X1_LOC_532/B 0.04fF
C28190 AND2X1_LOC_91/B OR2X1_LOC_489/A 0.01fF
C28191 OR2X1_LOC_62/A AND2X1_LOC_4/a_8_24# 0.02fF
C28192 OR2X1_LOC_816/A AND2X1_LOC_242/a_8_24# 0.03fF
C28193 OR2X1_LOC_680/A OR2X1_LOC_331/a_8_216# 0.09fF
C28194 OR2X1_LOC_85/A AND2X1_LOC_205/a_36_24# 0.00fF
C28195 OR2X1_LOC_147/B OR2X1_LOC_546/A 0.00fF
C28196 AND2X1_LOC_660/a_8_24# AND2X1_LOC_663/B 0.08fF
C28197 OR2X1_LOC_696/A AND2X1_LOC_243/Y 0.07fF
C28198 OR2X1_LOC_502/A OR2X1_LOC_446/B 0.10fF
C28199 OR2X1_LOC_64/Y OR2X1_LOC_31/Y 1.39fF
C28200 AND2X1_LOC_191/Y AND2X1_LOC_480/a_36_24# 0.01fF
C28201 OR2X1_LOC_118/Y AND2X1_LOC_657/A 0.01fF
C28202 OR2X1_LOC_834/A OR2X1_LOC_308/Y 0.00fF
C28203 OR2X1_LOC_631/A OR2X1_LOC_115/B 0.03fF
C28204 OR2X1_LOC_177/Y OR2X1_LOC_373/a_8_216# 0.01fF
C28205 OR2X1_LOC_338/a_8_216# AND2X1_LOC_22/Y 0.06fF
C28206 AND2X1_LOC_91/B OR2X1_LOC_772/A 0.02fF
C28207 AND2X1_LOC_784/A AND2X1_LOC_222/Y 0.00fF
C28208 OR2X1_LOC_677/Y OR2X1_LOC_142/Y 0.02fF
C28209 OR2X1_LOC_70/Y OR2X1_LOC_289/Y 0.03fF
C28210 OR2X1_LOC_294/Y OR2X1_LOC_580/B 0.03fF
C28211 AND2X1_LOC_727/A AND2X1_LOC_796/Y 0.01fF
C28212 OR2X1_LOC_36/Y AND2X1_LOC_793/B 0.03fF
C28213 OR2X1_LOC_136/a_8_216# VDD 0.21fF
C28214 AND2X1_LOC_542/a_8_24# OR2X1_LOC_373/Y 0.01fF
C28215 AND2X1_LOC_34/a_36_24# OR2X1_LOC_598/A 0.00fF
C28216 OR2X1_LOC_158/A AND2X1_LOC_802/Y 0.03fF
C28217 OR2X1_LOC_45/B AND2X1_LOC_778/Y 0.01fF
C28218 OR2X1_LOC_31/Y OR2X1_LOC_417/A 0.17fF
C28219 AND2X1_LOC_333/a_8_24# OR2X1_LOC_289/Y 0.05fF
C28220 AND2X1_LOC_566/B OR2X1_LOC_16/A 0.03fF
C28221 OR2X1_LOC_596/a_8_216# OR2X1_LOC_161/B 0.01fF
C28222 OR2X1_LOC_306/a_8_216# OR2X1_LOC_13/B 0.01fF
C28223 OR2X1_LOC_47/Y OR2X1_LOC_22/A 0.63fF
C28224 OR2X1_LOC_19/B AND2X1_LOC_646/a_8_24# 0.03fF
C28225 AND2X1_LOC_65/A OR2X1_LOC_549/A 0.10fF
C28226 AND2X1_LOC_683/a_8_24# AND2X1_LOC_31/Y 0.01fF
C28227 OR2X1_LOC_632/Y OR2X1_LOC_115/B 0.68fF
C28228 OR2X1_LOC_666/A AND2X1_LOC_287/B 0.00fF
C28229 OR2X1_LOC_417/A AND2X1_LOC_655/a_36_24# 0.01fF
C28230 INPUT_1 AND2X1_LOC_838/B 0.01fF
C28231 OR2X1_LOC_154/A OR2X1_LOC_515/a_36_216# 0.00fF
C28232 OR2X1_LOC_596/A OR2X1_LOC_515/A 0.02fF
C28233 AND2X1_LOC_69/Y AND2X1_LOC_31/Y 0.01fF
C28234 AND2X1_LOC_810/A AND2X1_LOC_715/A 0.03fF
C28235 VDD OR2X1_LOC_659/Y -0.00fF
C28236 AND2X1_LOC_95/Y OR2X1_LOC_523/a_36_216# 0.00fF
C28237 OR2X1_LOC_362/A OR2X1_LOC_349/A 0.02fF
C28238 OR2X1_LOC_70/Y OR2X1_LOC_534/a_8_216# 0.01fF
C28239 AND2X1_LOC_207/a_36_24# OR2X1_LOC_53/Y 0.00fF
C28240 OR2X1_LOC_539/Y OR2X1_LOC_175/a_8_216# 0.01fF
C28241 OR2X1_LOC_97/A OR2X1_LOC_168/B 0.17fF
C28242 OR2X1_LOC_532/B OR2X1_LOC_214/B 0.03fF
C28243 VDD OR2X1_LOC_162/a_8_216# 0.00fF
C28244 OR2X1_LOC_653/Y OR2X1_LOC_390/B 0.04fF
C28245 OR2X1_LOC_532/B OR2X1_LOC_241/B 0.07fF
C28246 AND2X1_LOC_774/a_8_24# OR2X1_LOC_91/A 0.12fF
C28247 OR2X1_LOC_590/a_8_216# OR2X1_LOC_814/A 0.02fF
C28248 OR2X1_LOC_715/B OR2X1_LOC_776/Y 0.38fF
C28249 OR2X1_LOC_78/A OR2X1_LOC_435/A 0.01fF
C28250 OR2X1_LOC_476/B OR2X1_LOC_228/Y 0.04fF
C28251 OR2X1_LOC_659/A OR2X1_LOC_576/A 0.50fF
C28252 OR2X1_LOC_516/B AND2X1_LOC_804/A 0.01fF
C28253 VDD AND2X1_LOC_347/B 0.01fF
C28254 OR2X1_LOC_417/Y OR2X1_LOC_534/Y 0.09fF
C28255 OR2X1_LOC_828/B AND2X1_LOC_409/B 0.10fF
C28256 OR2X1_LOC_656/B AND2X1_LOC_64/Y 0.03fF
C28257 OR2X1_LOC_56/A AND2X1_LOC_477/Y 0.03fF
C28258 AND2X1_LOC_367/A OR2X1_LOC_323/Y 0.10fF
C28259 OR2X1_LOC_644/a_8_216# OR2X1_LOC_228/Y 0.02fF
C28260 OR2X1_LOC_828/B AND2X1_LOC_763/B 0.04fF
C28261 AND2X1_LOC_370/a_36_24# AND2X1_LOC_716/Y 0.01fF
C28262 AND2X1_LOC_410/a_36_24# OR2X1_LOC_600/A -0.00fF
C28263 AND2X1_LOC_91/B AND2X1_LOC_104/a_8_24# 0.01fF
C28264 D_INPUT_5 OR2X1_LOC_375/Y 0.01fF
C28265 OR2X1_LOC_185/A OR2X1_LOC_722/B 0.00fF
C28266 OR2X1_LOC_49/A AND2X1_LOC_40/Y 0.02fF
C28267 OR2X1_LOC_485/A OR2X1_LOC_248/A 0.01fF
C28268 OR2X1_LOC_40/Y OR2X1_LOC_12/a_8_216# 0.01fF
C28269 OR2X1_LOC_122/a_8_216# AND2X1_LOC_243/Y 0.06fF
C28270 OR2X1_LOC_40/Y AND2X1_LOC_865/A 0.05fF
C28271 OR2X1_LOC_759/A AND2X1_LOC_658/A 0.03fF
C28272 OR2X1_LOC_510/Y OR2X1_LOC_140/B 0.00fF
C28273 AND2X1_LOC_733/Y AND2X1_LOC_443/a_8_24# 0.07fF
C28274 AND2X1_LOC_717/Y AND2X1_LOC_464/A 0.01fF
C28275 AND2X1_LOC_787/A AND2X1_LOC_168/Y 0.01fF
C28276 OR2X1_LOC_858/A AND2X1_LOC_18/Y 0.02fF
C28277 AND2X1_LOC_465/A OR2X1_LOC_39/A 0.02fF
C28278 OR2X1_LOC_831/A OR2X1_LOC_808/A 0.02fF
C28279 AND2X1_LOC_12/Y OR2X1_LOC_175/Y 0.03fF
C28280 OR2X1_LOC_715/B OR2X1_LOC_756/B 0.01fF
C28281 VDD OR2X1_LOC_442/Y 0.12fF
C28282 OR2X1_LOC_784/Y AND2X1_LOC_44/Y 0.21fF
C28283 AND2X1_LOC_7/B OR2X1_LOC_541/B 0.08fF
C28284 AND2X1_LOC_305/a_8_24# AND2X1_LOC_44/Y 0.00fF
C28285 OR2X1_LOC_499/a_8_216# OR2X1_LOC_563/A 0.40fF
C28286 AND2X1_LOC_804/Y AND2X1_LOC_727/B 0.03fF
C28287 AND2X1_LOC_392/A AND2X1_LOC_364/Y 0.01fF
C28288 OR2X1_LOC_458/B OR2X1_LOC_723/a_8_216# 0.01fF
C28289 AND2X1_LOC_40/Y OR2X1_LOC_596/A 0.05fF
C28290 AND2X1_LOC_716/Y AND2X1_LOC_212/A 0.04fF
C28291 AND2X1_LOC_570/Y OR2X1_LOC_59/Y 0.03fF
C28292 OR2X1_LOC_45/B AND2X1_LOC_862/A 0.08fF
C28293 OR2X1_LOC_331/A OR2X1_LOC_59/Y 0.01fF
C28294 AND2X1_LOC_582/a_8_24# OR2X1_LOC_686/A 0.08fF
C28295 OR2X1_LOC_175/Y OR2X1_LOC_802/A 0.02fF
C28296 AND2X1_LOC_59/Y OR2X1_LOC_97/A 0.10fF
C28297 OR2X1_LOC_45/B AND2X1_LOC_624/A 0.10fF
C28298 OR2X1_LOC_502/A AND2X1_LOC_165/a_36_24# 0.01fF
C28299 OR2X1_LOC_738/A AND2X1_LOC_44/Y 0.14fF
C28300 AND2X1_LOC_12/Y OR2X1_LOC_691/Y 0.02fF
C28301 AND2X1_LOC_92/Y OR2X1_LOC_520/a_8_216# 0.01fF
C28302 OR2X1_LOC_710/A OR2X1_LOC_708/B 0.82fF
C28303 OR2X1_LOC_329/B OR2X1_LOC_56/A 0.20fF
C28304 OR2X1_LOC_325/A AND2X1_LOC_322/a_8_24# 0.23fF
C28305 OR2X1_LOC_810/A OR2X1_LOC_140/B 0.05fF
C28306 AND2X1_LOC_539/Y AND2X1_LOC_661/A 0.53fF
C28307 OR2X1_LOC_813/A OR2X1_LOC_71/A 0.14fF
C28308 AND2X1_LOC_81/B OR2X1_LOC_139/A 0.05fF
C28309 AND2X1_LOC_605/Y AND2X1_LOC_447/Y 0.02fF
C28310 AND2X1_LOC_212/A AND2X1_LOC_654/Y 0.02fF
C28311 AND2X1_LOC_749/a_8_24# AND2X1_LOC_18/Y 0.01fF
C28312 AND2X1_LOC_535/Y OR2X1_LOC_92/Y 0.03fF
C28313 AND2X1_LOC_705/Y AND2X1_LOC_593/Y 0.07fF
C28314 OR2X1_LOC_62/A OR2X1_LOC_68/B 2.41fF
C28315 AND2X1_LOC_339/B OR2X1_LOC_18/Y 0.03fF
C28316 OR2X1_LOC_64/Y OR2X1_LOC_320/a_8_216# 0.11fF
C28317 AND2X1_LOC_566/B AND2X1_LOC_661/a_8_24# 0.01fF
C28318 OR2X1_LOC_375/A AND2X1_LOC_603/a_8_24# 0.01fF
C28319 AND2X1_LOC_12/Y OR2X1_LOC_713/A 0.03fF
C28320 VDD OR2X1_LOC_16/a_8_216# 0.00fF
C28321 OR2X1_LOC_768/A OR2X1_LOC_235/B 0.01fF
C28322 OR2X1_LOC_151/A OR2X1_LOC_447/A 0.07fF
C28323 VDD OR2X1_LOC_448/A 0.21fF
C28324 OR2X1_LOC_49/A OR2X1_LOC_87/Y 0.01fF
C28325 AND2X1_LOC_191/B AND2X1_LOC_456/B 0.03fF
C28326 OR2X1_LOC_6/B AND2X1_LOC_398/a_8_24# 0.01fF
C28327 OR2X1_LOC_770/B OR2X1_LOC_848/A 0.17fF
C28328 AND2X1_LOC_91/B AND2X1_LOC_3/Y 0.08fF
C28329 OR2X1_LOC_6/A AND2X1_LOC_786/Y 0.02fF
C28330 OR2X1_LOC_614/Y AND2X1_LOC_43/B 0.06fF
C28331 OR2X1_LOC_686/A AND2X1_LOC_682/a_8_24# 0.27fF
C28332 AND2X1_LOC_70/Y OR2X1_LOC_330/Y 0.02fF
C28333 OR2X1_LOC_589/A AND2X1_LOC_436/B 0.09fF
C28334 VDD OR2X1_LOC_40/a_8_216# 0.00fF
C28335 OR2X1_LOC_26/Y OR2X1_LOC_428/A 0.90fF
C28336 AND2X1_LOC_47/Y OR2X1_LOC_735/B 0.01fF
C28337 OR2X1_LOC_44/Y AND2X1_LOC_774/A 0.00fF
C28338 OR2X1_LOC_235/B AND2X1_LOC_71/a_8_24# 0.11fF
C28339 OR2X1_LOC_589/A AND2X1_LOC_139/B 0.23fF
C28340 AND2X1_LOC_535/Y AND2X1_LOC_801/a_36_24# 0.00fF
C28341 OR2X1_LOC_40/Y AND2X1_LOC_676/a_8_24# 0.04fF
C28342 AND2X1_LOC_663/B AND2X1_LOC_792/a_8_24# 0.00fF
C28343 OR2X1_LOC_662/a_8_216# OR2X1_LOC_663/A 0.01fF
C28344 AND2X1_LOC_498/a_36_24# OR2X1_LOC_499/B -0.00fF
C28345 OR2X1_LOC_244/A OR2X1_LOC_217/A 0.01fF
C28346 OR2X1_LOC_600/A OR2X1_LOC_625/Y 0.07fF
C28347 AND2X1_LOC_95/Y AND2X1_LOC_184/a_8_24# 0.04fF
C28348 INPUT_0 OR2X1_LOC_637/A 0.02fF
C28349 OR2X1_LOC_160/B OR2X1_LOC_185/A 0.05fF
C28350 AND2X1_LOC_160/a_8_24# OR2X1_LOC_697/Y 0.01fF
C28351 OR2X1_LOC_26/Y OR2X1_LOC_595/A 0.47fF
C28352 OR2X1_LOC_147/A OR2X1_LOC_469/Y 0.03fF
C28353 VDD OR2X1_LOC_118/Y 0.38fF
C28354 OR2X1_LOC_160/B OR2X1_LOC_249/Y 0.01fF
C28355 OR2X1_LOC_89/A OR2X1_LOC_428/A 0.09fF
C28356 AND2X1_LOC_705/Y AND2X1_LOC_602/a_8_24# 0.10fF
C28357 AND2X1_LOC_376/a_8_24# OR2X1_LOC_375/Y 0.03fF
C28358 OR2X1_LOC_852/a_36_216# OR2X1_LOC_472/A 0.02fF
C28359 OR2X1_LOC_155/A OR2X1_LOC_435/A 0.01fF
C28360 OR2X1_LOC_420/a_8_216# OR2X1_LOC_12/Y 0.03fF
C28361 VDD AND2X1_LOC_601/a_8_24# -0.00fF
C28362 VDD AND2X1_LOC_453/a_8_24# 0.00fF
C28363 OR2X1_LOC_89/A OR2X1_LOC_595/A 4.49fF
C28364 OR2X1_LOC_405/A OR2X1_LOC_78/B 0.11fF
C28365 AND2X1_LOC_257/a_8_24# OR2X1_LOC_259/B 0.00fF
C28366 OR2X1_LOC_45/B AND2X1_LOC_853/a_8_24# 0.09fF
C28367 AND2X1_LOC_113/Y OR2X1_LOC_56/A 0.03fF
C28368 OR2X1_LOC_6/B OR2X1_LOC_43/A 4.64fF
C28369 OR2X1_LOC_769/A OR2X1_LOC_160/A 0.02fF
C28370 AND2X1_LOC_547/Y AND2X1_LOC_564/a_8_24# 0.00fF
C28371 OR2X1_LOC_74/A OR2X1_LOC_323/Y 0.02fF
C28372 OR2X1_LOC_605/B AND2X1_LOC_603/a_8_24# 0.01fF
C28373 AND2X1_LOC_348/Y AND2X1_LOC_860/A 0.03fF
C28374 OR2X1_LOC_674/Y OR2X1_LOC_142/Y 0.03fF
C28375 OR2X1_LOC_166/Y AND2X1_LOC_436/B 0.02fF
C28376 AND2X1_LOC_72/B OR2X1_LOC_501/a_8_216# 0.01fF
C28377 OR2X1_LOC_527/Y AND2X1_LOC_785/Y 0.11fF
C28378 OR2X1_LOC_64/Y OR2X1_LOC_79/a_8_216# 0.01fF
C28379 AND2X1_LOC_72/a_8_24# OR2X1_LOC_719/B 0.04fF
C28380 OR2X1_LOC_648/A OR2X1_LOC_130/A 0.02fF
C28381 OR2X1_LOC_753/A AND2X1_LOC_860/A 0.07fF
C28382 OR2X1_LOC_158/A AND2X1_LOC_154/Y 0.04fF
C28383 OR2X1_LOC_669/a_36_216# AND2X1_LOC_860/A 0.01fF
C28384 OR2X1_LOC_89/a_8_216# AND2X1_LOC_243/Y 0.02fF
C28385 AND2X1_LOC_215/Y OR2X1_LOC_26/Y 0.00fF
C28386 AND2X1_LOC_59/Y OR2X1_LOC_541/A 0.01fF
C28387 AND2X1_LOC_31/Y OR2X1_LOC_364/Y 0.01fF
C28388 VDD OR2X1_LOC_262/Y 0.19fF
C28389 OR2X1_LOC_656/B OR2X1_LOC_656/Y 0.40fF
C28390 AND2X1_LOC_537/a_8_24# OR2X1_LOC_585/A 0.01fF
C28391 AND2X1_LOC_477/a_8_24# OR2X1_LOC_39/A 0.14fF
C28392 OR2X1_LOC_676/Y AND2X1_LOC_516/a_8_24# 0.03fF
C28393 AND2X1_LOC_858/B AND2X1_LOC_286/Y 0.01fF
C28394 OR2X1_LOC_405/A OR2X1_LOC_721/Y 0.02fF
C28395 OR2X1_LOC_426/B OR2X1_LOC_86/a_8_216# 0.03fF
C28396 OR2X1_LOC_811/A OR2X1_LOC_737/A 0.14fF
C28397 VDD OR2X1_LOC_238/Y 0.27fF
C28398 D_INPUT_0 OR2X1_LOC_392/B 0.10fF
C28399 VDD OR2X1_LOC_24/Y 0.07fF
C28400 OR2X1_LOC_71/Y AND2X1_LOC_242/B 0.01fF
C28401 OR2X1_LOC_755/a_8_216# OR2X1_LOC_44/Y 0.01fF
C28402 OR2X1_LOC_188/Y OR2X1_LOC_532/B 0.03fF
C28403 OR2X1_LOC_22/Y OR2X1_LOC_522/a_8_216# 0.08fF
C28404 AND2X1_LOC_501/Y AND2X1_LOC_191/Y 0.03fF
C28405 AND2X1_LOC_95/Y OR2X1_LOC_811/A 0.03fF
C28406 OR2X1_LOC_175/B OR2X1_LOC_161/A 0.00fF
C28407 AND2X1_LOC_59/Y OR2X1_LOC_475/B 0.04fF
C28408 AND2X1_LOC_539/Y AND2X1_LOC_810/Y 0.20fF
C28409 AND2X1_LOC_510/A OR2X1_LOC_7/A 0.01fF
C28410 AND2X1_LOC_191/B AND2X1_LOC_717/B 0.00fF
C28411 AND2X1_LOC_42/B OR2X1_LOC_66/A 6.03fF
C28412 AND2X1_LOC_501/Y AND2X1_LOC_711/Y 0.03fF
C28413 AND2X1_LOC_12/Y OR2X1_LOC_629/Y 0.05fF
C28414 AND2X1_LOC_784/A AND2X1_LOC_367/A 0.07fF
C28415 AND2X1_LOC_388/Y OR2X1_LOC_417/Y 0.03fF
C28416 AND2X1_LOC_191/Y AND2X1_LOC_570/Y 0.03fF
C28417 OR2X1_LOC_3/Y AND2X1_LOC_285/Y 0.01fF
C28418 AND2X1_LOC_753/B OR2X1_LOC_375/A 0.68fF
C28419 AND2X1_LOC_86/Y OR2X1_LOC_185/A 0.10fF
C28420 AND2X1_LOC_663/B AND2X1_LOC_243/Y 0.10fF
C28421 AND2X1_LOC_207/a_8_24# OR2X1_LOC_585/A 0.07fF
C28422 AND2X1_LOC_41/A OR2X1_LOC_449/B 0.07fF
C28423 OR2X1_LOC_246/Y OR2X1_LOC_92/Y 0.13fF
C28424 AND2X1_LOC_570/Y AND2X1_LOC_711/Y 0.03fF
C28425 INPUT_3 OR2X1_LOC_185/A 0.03fF
C28426 OR2X1_LOC_502/A AND2X1_LOC_56/B 0.17fF
C28427 AND2X1_LOC_674/a_36_24# OR2X1_LOC_733/A 0.00fF
C28428 OR2X1_LOC_151/A AND2X1_LOC_127/a_8_24# 0.01fF
C28429 AND2X1_LOC_533/a_8_24# AND2X1_LOC_95/Y 0.04fF
C28430 AND2X1_LOC_523/a_8_24# OR2X1_LOC_39/A 0.01fF
C28431 AND2X1_LOC_70/Y AND2X1_LOC_117/a_8_24# 0.01fF
C28432 AND2X1_LOC_30/a_8_24# D_INPUT_4 0.04fF
C28433 OR2X1_LOC_331/A OR2X1_LOC_70/Y 0.37fF
C28434 OR2X1_LOC_694/Y OR2X1_LOC_64/Y 0.01fF
C28435 AND2X1_LOC_47/Y OR2X1_LOC_161/B 0.84fF
C28436 AND2X1_LOC_554/Y AND2X1_LOC_573/A 0.01fF
C28437 OR2X1_LOC_831/B D_INPUT_1 0.06fF
C28438 OR2X1_LOC_405/A OR2X1_LOC_375/A 0.07fF
C28439 AND2X1_LOC_473/a_8_24# OR2X1_LOC_59/Y 0.01fF
C28440 OR2X1_LOC_8/Y OR2X1_LOC_5/a_8_216# 0.18fF
C28441 OR2X1_LOC_158/A INPUT_1 0.30fF
C28442 OR2X1_LOC_502/A AND2X1_LOC_8/Y 0.07fF
C28443 OR2X1_LOC_671/Y D_INPUT_0 0.00fF
C28444 OR2X1_LOC_298/a_8_216# OR2X1_LOC_7/A 0.01fF
C28445 OR2X1_LOC_185/A OR2X1_LOC_553/A 0.02fF
C28446 AND2X1_LOC_724/A OR2X1_LOC_95/Y 0.09fF
C28447 AND2X1_LOC_365/A AND2X1_LOC_436/B 0.05fF
C28448 OR2X1_LOC_485/A OR2X1_LOC_594/a_8_216# 0.01fF
C28449 AND2X1_LOC_208/B OR2X1_LOC_24/Y 0.05fF
C28450 OR2X1_LOC_770/A D_INPUT_1 0.28fF
C28451 AND2X1_LOC_91/B AND2X1_LOC_225/a_8_24# 0.05fF
C28452 OR2X1_LOC_160/A OR2X1_LOC_87/a_36_216# 0.00fF
C28453 OR2X1_LOC_185/A OR2X1_LOC_266/a_8_216# 0.02fF
C28454 OR2X1_LOC_759/A AND2X1_LOC_814/a_8_24# 0.01fF
C28455 AND2X1_LOC_727/a_36_24# AND2X1_LOC_810/Y 0.00fF
C28456 OR2X1_LOC_237/Y OR2X1_LOC_39/A 0.06fF
C28457 OR2X1_LOC_115/a_8_216# OR2X1_LOC_203/Y 0.01fF
C28458 OR2X1_LOC_502/A AND2X1_LOC_21/Y 0.50fF
C28459 OR2X1_LOC_43/a_8_216# AND2X1_LOC_434/Y 0.03fF
C28460 OR2X1_LOC_385/Y OR2X1_LOC_586/a_8_216# 0.03fF
C28461 OR2X1_LOC_744/A OR2X1_LOC_277/a_36_216# 0.00fF
C28462 OR2X1_LOC_160/B OR2X1_LOC_750/a_36_216# 0.00fF
C28463 OR2X1_LOC_640/a_36_216# OR2X1_LOC_462/B 0.00fF
C28464 AND2X1_LOC_845/Y AND2X1_LOC_860/A 0.31fF
C28465 OR2X1_LOC_467/A AND2X1_LOC_694/a_8_24# 0.01fF
C28466 AND2X1_LOC_537/Y AND2X1_LOC_434/Y 0.00fF
C28467 VDD AND2X1_LOC_7/Y 0.21fF
C28468 OR2X1_LOC_43/A AND2X1_LOC_436/B 0.00fF
C28469 AND2X1_LOC_703/a_8_24# OR2X1_LOC_485/A 0.02fF
C28470 OR2X1_LOC_185/A OR2X1_LOC_219/B 0.00fF
C28471 OR2X1_LOC_139/A OR2X1_LOC_66/Y 0.01fF
C28472 AND2X1_LOC_41/A OR2X1_LOC_121/B 0.11fF
C28473 AND2X1_LOC_329/a_8_24# OR2X1_LOC_739/A 0.01fF
C28474 OR2X1_LOC_87/B OR2X1_LOC_87/Y 0.01fF
C28475 OR2X1_LOC_22/Y AND2X1_LOC_858/B 0.17fF
C28476 OR2X1_LOC_470/B OR2X1_LOC_469/Y 0.03fF
C28477 AND2X1_LOC_72/B AND2X1_LOC_44/Y 0.02fF
C28478 OR2X1_LOC_43/A AND2X1_LOC_139/B 8.99fF
C28479 OR2X1_LOC_32/B OR2X1_LOC_52/B 0.11fF
C28480 OR2X1_LOC_22/Y OR2X1_LOC_91/A 0.94fF
C28481 AND2X1_LOC_72/Y AND2X1_LOC_3/Y 0.01fF
C28482 AND2X1_LOC_36/Y OR2X1_LOC_317/B 0.03fF
C28483 OR2X1_LOC_235/B OR2X1_LOC_46/A 0.08fF
C28484 OR2X1_LOC_485/A AND2X1_LOC_468/B 3.87fF
C28485 AND2X1_LOC_44/Y OR2X1_LOC_512/a_36_216# 0.00fF
C28486 OR2X1_LOC_280/Y AND2X1_LOC_573/A 0.02fF
C28487 OR2X1_LOC_342/B OR2X1_LOC_349/B 0.80fF
C28488 AND2X1_LOC_859/Y OR2X1_LOC_36/Y 0.07fF
C28489 OR2X1_LOC_154/A OR2X1_LOC_68/a_8_216# 0.01fF
C28490 OR2X1_LOC_404/A OR2X1_LOC_78/Y 0.12fF
C28491 OR2X1_LOC_161/B OR2X1_LOC_598/A 0.88fF
C28492 AND2X1_LOC_729/Y OR2X1_LOC_74/A 0.03fF
C28493 AND2X1_LOC_98/Y INPUT_1 0.00fF
C28494 AND2X1_LOC_702/a_8_24# OR2X1_LOC_304/Y 0.10fF
C28495 D_INPUT_7 AND2X1_LOC_1/a_8_24# 0.01fF
C28496 OR2X1_LOC_777/B OR2X1_LOC_180/B 0.17fF
C28497 AND2X1_LOC_126/a_8_24# OR2X1_LOC_243/B 0.11fF
C28498 OR2X1_LOC_829/a_36_216# AND2X1_LOC_729/B 0.01fF
C28499 OR2X1_LOC_831/A OR2X1_LOC_374/Y 0.03fF
C28500 AND2X1_LOC_329/a_8_24# OR2X1_LOC_269/B 0.03fF
C28501 OR2X1_LOC_223/A OR2X1_LOC_787/B 0.00fF
C28502 OR2X1_LOC_80/A AND2X1_LOC_202/Y 0.00fF
C28503 OR2X1_LOC_84/Y OR2X1_LOC_786/A 0.16fF
C28504 OR2X1_LOC_62/B OR2X1_LOC_574/a_36_216# 0.00fF
C28505 OR2X1_LOC_497/Y OR2X1_LOC_7/A 0.07fF
C28506 AND2X1_LOC_31/Y OR2X1_LOC_708/a_8_216# 0.01fF
C28507 AND2X1_LOC_727/A AND2X1_LOC_654/Y 0.05fF
C28508 AND2X1_LOC_10/a_8_24# OR2X1_LOC_375/A 0.03fF
C28509 AND2X1_LOC_738/B GATE_811 0.00fF
C28510 OR2X1_LOC_435/B AND2X1_LOC_47/Y 0.08fF
C28511 AND2X1_LOC_327/a_8_24# OR2X1_LOC_65/B -0.00fF
C28512 OR2X1_LOC_223/A AND2X1_LOC_92/Y 0.04fF
C28513 AND2X1_LOC_570/Y OR2X1_LOC_184/Y 0.55fF
C28514 OR2X1_LOC_305/Y OR2X1_LOC_3/Y 0.14fF
C28515 AND2X1_LOC_48/a_8_24# AND2X1_LOC_47/Y 0.05fF
C28516 OR2X1_LOC_19/B OR2X1_LOC_256/a_36_216# 0.03fF
C28517 AND2X1_LOC_784/A OR2X1_LOC_74/A 0.24fF
C28518 AND2X1_LOC_374/Y OR2X1_LOC_371/Y 0.03fF
C28519 AND2X1_LOC_58/a_36_24# D_INPUT_0 0.00fF
C28520 AND2X1_LOC_363/B OR2X1_LOC_417/A 0.04fF
C28521 AND2X1_LOC_34/Y OR2X1_LOC_416/Y 0.01fF
C28522 AND2X1_LOC_569/A AND2X1_LOC_578/A 0.06fF
C28523 OR2X1_LOC_127/Y OR2X1_LOC_125/Y 0.04fF
C28524 OR2X1_LOC_847/A INPUT_1 0.02fF
C28525 AND2X1_LOC_820/a_8_24# D_INPUT_0 0.03fF
C28526 OR2X1_LOC_22/Y AND2X1_LOC_573/A 0.14fF
C28527 AND2X1_LOC_171/a_8_24# OR2X1_LOC_333/B 0.01fF
C28528 OR2X1_LOC_795/a_8_216# OR2X1_LOC_795/B 0.39fF
C28529 OR2X1_LOC_7/A OR2X1_LOC_229/Y 0.03fF
C28530 AND2X1_LOC_342/Y OR2X1_LOC_54/Y 0.09fF
C28531 AND2X1_LOC_91/B OR2X1_LOC_576/a_8_216# 0.02fF
C28532 OR2X1_LOC_348/Y OR2X1_LOC_675/Y 0.07fF
C28533 AND2X1_LOC_287/B OR2X1_LOC_13/B 0.00fF
C28534 OR2X1_LOC_462/B OR2X1_LOC_19/B 0.03fF
C28535 OR2X1_LOC_185/Y AND2X1_LOC_816/a_8_24# 0.01fF
C28536 OR2X1_LOC_185/A OR2X1_LOC_244/A 0.13fF
C28537 AND2X1_LOC_492/a_36_24# OR2X1_LOC_532/B 0.01fF
C28538 AND2X1_LOC_663/B AND2X1_LOC_620/a_8_24# 0.01fF
C28539 AND2X1_LOC_12/Y AND2X1_LOC_283/a_8_24# 0.01fF
C28540 OR2X1_LOC_816/A OR2X1_LOC_13/B 0.03fF
C28541 AND2X1_LOC_692/a_36_24# AND2X1_LOC_43/B 0.01fF
C28542 OR2X1_LOC_51/Y OR2X1_LOC_163/a_8_216# 0.07fF
C28543 AND2X1_LOC_784/Y AND2X1_LOC_796/A 0.02fF
C28544 AND2X1_LOC_371/a_8_24# AND2X1_LOC_31/Y 0.04fF
C28545 OR2X1_LOC_391/B OR2X1_LOC_772/Y 0.05fF
C28546 OR2X1_LOC_405/Y OR2X1_LOC_532/B 0.01fF
C28547 AND2X1_LOC_56/B AND2X1_LOC_48/A 0.10fF
C28548 OR2X1_LOC_154/A OR2X1_LOC_814/A 0.32fF
C28549 OR2X1_LOC_391/B OR2X1_LOC_846/A 0.22fF
C28550 OR2X1_LOC_256/A OR2X1_LOC_118/Y 0.03fF
C28551 OR2X1_LOC_355/B AND2X1_LOC_51/Y 0.23fF
C28552 AND2X1_LOC_31/Y AND2X1_LOC_18/Y 0.63fF
C28553 AND2X1_LOC_518/a_8_24# AND2X1_LOC_8/Y 0.01fF
C28554 OR2X1_LOC_604/A AND2X1_LOC_793/B 0.07fF
C28555 OR2X1_LOC_185/Y OR2X1_LOC_859/A 0.12fF
C28556 OR2X1_LOC_485/A AND2X1_LOC_830/a_8_24# 0.01fF
C28557 OR2X1_LOC_604/A OR2X1_LOC_533/A 0.03fF
C28558 OR2X1_LOC_246/A OR2X1_LOC_86/a_8_216# 0.05fF
C28559 AND2X1_LOC_48/A AND2X1_LOC_8/Y 0.03fF
C28560 OR2X1_LOC_404/Y OR2X1_LOC_557/A 0.00fF
C28561 OR2X1_LOC_575/A D_INPUT_1 0.03fF
C28562 OR2X1_LOC_267/A OR2X1_LOC_814/A 0.02fF
C28563 AND2X1_LOC_390/B OR2X1_LOC_829/Y 0.03fF
C28564 OR2X1_LOC_773/a_8_216# OR2X1_LOC_269/B 0.01fF
C28565 OR2X1_LOC_312/Y AND2X1_LOC_727/A 0.03fF
C28566 OR2X1_LOC_3/Y OR2X1_LOC_417/Y 0.03fF
C28567 AND2X1_LOC_811/Y AND2X1_LOC_624/A 0.13fF
C28568 OR2X1_LOC_3/Y OR2X1_LOC_291/Y 0.03fF
C28569 AND2X1_LOC_568/a_8_24# OR2X1_LOC_417/Y 0.01fF
C28570 AND2X1_LOC_566/Y AND2X1_LOC_514/Y 0.02fF
C28571 OR2X1_LOC_618/Y AND2X1_LOC_9/a_8_24# 0.10fF
C28572 AND2X1_LOC_36/Y AND2X1_LOC_44/Y 0.43fF
C28573 AND2X1_LOC_91/a_8_24# OR2X1_LOC_605/Y 0.17fF
C28574 OR2X1_LOC_613/Y AND2X1_LOC_866/a_8_24# 0.01fF
C28575 AND2X1_LOC_36/Y OR2X1_LOC_514/a_8_216# 0.01fF
C28576 OR2X1_LOC_312/Y OR2X1_LOC_95/Y 0.03fF
C28577 OR2X1_LOC_703/Y OR2X1_LOC_356/A 0.15fF
C28578 AND2X1_LOC_44/Y OR2X1_LOC_333/a_8_216# 0.03fF
C28579 OR2X1_LOC_516/Y AND2X1_LOC_212/Y 0.00fF
C28580 OR2X1_LOC_22/Y OR2X1_LOC_27/Y 0.03fF
C28581 OR2X1_LOC_22/Y AND2X1_LOC_662/a_8_24# 0.02fF
C28582 OR2X1_LOC_462/a_8_216# OR2X1_LOC_472/B 0.01fF
C28583 OR2X1_LOC_312/Y OR2X1_LOC_368/A 0.00fF
C28584 OR2X1_LOC_696/A OR2X1_LOC_12/Y 0.72fF
C28585 OR2X1_LOC_772/a_8_216# D_INPUT_1 0.02fF
C28586 OR2X1_LOC_161/B OR2X1_LOC_186/a_8_216# 0.01fF
C28587 AND2X1_LOC_728/a_36_24# OR2X1_LOC_679/A 0.00fF
C28588 AND2X1_LOC_34/a_36_24# AND2X1_LOC_462/Y 0.00fF
C28589 AND2X1_LOC_863/Y AND2X1_LOC_212/B 0.02fF
C28590 OR2X1_LOC_193/A OR2X1_LOC_532/B 0.28fF
C28591 OR2X1_LOC_488/a_8_216# OR2X1_LOC_417/A 0.01fF
C28592 OR2X1_LOC_232/a_8_216# OR2X1_LOC_47/Y 0.01fF
C28593 AND2X1_LOC_544/Y AND2X1_LOC_213/B 0.03fF
C28594 AND2X1_LOC_358/a_36_24# OR2X1_LOC_46/A 0.00fF
C28595 OR2X1_LOC_3/Y D_INPUT_3 0.91fF
C28596 AND2X1_LOC_170/B AND2X1_LOC_798/Y 0.03fF
C28597 OR2X1_LOC_783/a_8_216# OR2X1_LOC_155/A 0.01fF
C28598 AND2X1_LOC_775/a_8_24# OR2X1_LOC_406/A 0.20fF
C28599 AND2X1_LOC_42/B OR2X1_LOC_84/A 0.02fF
C28600 OR2X1_LOC_51/Y OR2X1_LOC_386/a_8_216# 0.01fF
C28601 AND2X1_LOC_361/a_8_24# OR2X1_LOC_106/Y 0.04fF
C28602 OR2X1_LOC_691/B OR2X1_LOC_853/a_8_216# 0.00fF
C28603 OR2X1_LOC_45/B AND2X1_LOC_774/A 0.64fF
C28604 AND2X1_LOC_339/Y OR2X1_LOC_16/A 0.01fF
C28605 OR2X1_LOC_18/Y OR2X1_LOC_521/a_8_216# 0.01fF
C28606 AND2X1_LOC_711/a_8_24# OR2X1_LOC_759/Y 0.23fF
C28607 AND2X1_LOC_8/Y OR2X1_LOC_398/a_8_216# 0.02fF
C28608 D_INPUT_0 OR2X1_LOC_532/B 0.54fF
C28609 OR2X1_LOC_545/B OR2X1_LOC_443/a_8_216# 0.01fF
C28610 OR2X1_LOC_617/a_36_216# AND2X1_LOC_624/B 0.00fF
C28611 AND2X1_LOC_738/B OR2X1_LOC_525/a_8_216# 0.03fF
C28612 OR2X1_LOC_52/B AND2X1_LOC_222/Y 0.02fF
C28613 AND2X1_LOC_340/Y AND2X1_LOC_339/B 1.74fF
C28614 OR2X1_LOC_737/A OR2X1_LOC_777/B 0.07fF
C28615 OR2X1_LOC_516/Y AND2X1_LOC_506/a_8_24# 0.02fF
C28616 OR2X1_LOC_161/A OR2X1_LOC_366/Y 0.03fF
C28617 OR2X1_LOC_18/Y OR2X1_LOC_300/Y 0.03fF
C28618 AND2X1_LOC_95/Y OR2X1_LOC_777/B 0.15fF
C28619 AND2X1_LOC_726/a_8_24# AND2X1_LOC_731/Y 0.11fF
C28620 OR2X1_LOC_70/Y OR2X1_LOC_406/A 0.48fF
C28621 OR2X1_LOC_3/Y AND2X1_LOC_656/a_8_24# 0.01fF
C28622 VDD AND2X1_LOC_208/Y 0.02fF
C28623 VDD OR2X1_LOC_375/a_8_216# 0.00fF
C28624 OR2X1_LOC_601/a_36_216# OR2X1_LOC_47/Y 0.01fF
C28625 VDD AND2X1_LOC_407/a_8_24# -0.00fF
C28626 OR2X1_LOC_3/B OR2X1_LOC_22/A 0.44fF
C28627 AND2X1_LOC_56/a_36_24# OR2X1_LOC_651/A 0.01fF
C28628 OR2X1_LOC_303/A OR2X1_LOC_566/A 0.06fF
C28629 OR2X1_LOC_62/a_36_216# D_INPUT_1 0.00fF
C28630 OR2X1_LOC_622/A OR2X1_LOC_633/A 0.03fF
C28631 OR2X1_LOC_756/B OR2X1_LOC_338/B 0.01fF
C28632 OR2X1_LOC_52/B OR2X1_LOC_423/Y 0.03fF
C28633 OR2X1_LOC_45/B AND2X1_LOC_434/a_8_24# 0.02fF
C28634 OR2X1_LOC_815/A AND2X1_LOC_793/Y 0.02fF
C28635 OR2X1_LOC_703/A OR2X1_LOC_703/a_8_216# 0.01fF
C28636 AND2X1_LOC_537/Y OR2X1_LOC_595/Y 0.14fF
C28637 VDD OR2X1_LOC_390/A 0.21fF
C28638 OR2X1_LOC_49/A OR2X1_LOC_90/a_8_216# 0.01fF
C28639 D_INPUT_3 OR2X1_LOC_673/A 0.15fF
C28640 AND2X1_LOC_318/Y AND2X1_LOC_319/a_8_24# 0.06fF
C28641 AND2X1_LOC_785/A OR2X1_LOC_18/Y 0.22fF
C28642 OR2X1_LOC_151/A OR2X1_LOC_440/a_8_216# 0.01fF
C28643 OR2X1_LOC_158/A AND2X1_LOC_709/a_8_24# 0.01fF
C28644 AND2X1_LOC_3/Y OR2X1_LOC_446/B 0.00fF
C28645 AND2X1_LOC_462/a_36_24# OR2X1_LOC_598/A 0.00fF
C28646 AND2X1_LOC_787/A AND2X1_LOC_722/Y 0.01fF
C28647 AND2X1_LOC_22/Y AND2X1_LOC_304/a_8_24# 0.01fF
C28648 AND2X1_LOC_91/B OR2X1_LOC_860/Y 0.03fF
C28649 AND2X1_LOC_392/A AND2X1_LOC_243/Y 0.07fF
C28650 OR2X1_LOC_158/A AND2X1_LOC_352/B 0.03fF
C28651 OR2X1_LOC_831/B OR2X1_LOC_737/A 0.07fF
C28652 OR2X1_LOC_542/B OR2X1_LOC_542/a_8_216# 0.06fF
C28653 AND2X1_LOC_511/a_8_24# OR2X1_LOC_78/A 0.01fF
C28654 OR2X1_LOC_543/A OR2X1_LOC_370/a_8_216# 0.01fF
C28655 OR2X1_LOC_78/A OR2X1_LOC_361/a_8_216# 0.02fF
C28656 AND2X1_LOC_392/A AND2X1_LOC_568/B 0.07fF
C28657 OR2X1_LOC_13/Y AND2X1_LOC_434/Y 0.02fF
C28658 OR2X1_LOC_756/B OR2X1_LOC_35/A 0.01fF
C28659 AND2X1_LOC_582/a_8_24# OR2X1_LOC_161/B 0.09fF
C28660 OR2X1_LOC_743/A OR2X1_LOC_424/Y 0.02fF
C28661 OR2X1_LOC_566/A AND2X1_LOC_95/Y 0.03fF
C28662 OR2X1_LOC_348/a_8_216# OR2X1_LOC_756/B 0.02fF
C28663 OR2X1_LOC_106/Y OR2X1_LOC_18/Y 0.00fF
C28664 OR2X1_LOC_166/a_8_216# AND2X1_LOC_535/Y 0.01fF
C28665 VDD OR2X1_LOC_797/a_8_216# 0.00fF
C28666 OR2X1_LOC_158/A AND2X1_LOC_296/a_36_24# 0.00fF
C28667 OR2X1_LOC_814/A OR2X1_LOC_560/A 0.03fF
C28668 AND2X1_LOC_91/B OR2X1_LOC_732/B 0.41fF
C28669 OR2X1_LOC_316/a_36_216# OR2X1_LOC_39/A 0.00fF
C28670 AND2X1_LOC_501/Y AND2X1_LOC_658/B 0.03fF
C28671 AND2X1_LOC_752/a_8_24# OR2X1_LOC_375/Y 0.23fF
C28672 AND2X1_LOC_219/a_8_24# AND2X1_LOC_61/Y 0.02fF
C28673 OR2X1_LOC_97/A OR2X1_LOC_794/A 0.03fF
C28674 AND2X1_LOC_91/B OR2X1_LOC_489/B -0.02fF
C28675 OR2X1_LOC_92/Y OR2X1_LOC_16/A 0.10fF
C28676 AND2X1_LOC_658/B AND2X1_LOC_570/Y 0.03fF
C28677 OR2X1_LOC_661/a_36_216# AND2X1_LOC_7/B 0.00fF
C28678 OR2X1_LOC_6/B OR2X1_LOC_630/B 0.01fF
C28679 AND2X1_LOC_22/Y AND2X1_LOC_59/a_8_24# 0.02fF
C28680 AND2X1_LOC_366/A AND2X1_LOC_243/Y 0.02fF
C28681 AND2X1_LOC_36/a_8_24# AND2X1_LOC_36/Y 0.01fF
C28682 OR2X1_LOC_158/A OR2X1_LOC_517/A 0.01fF
C28683 AND2X1_LOC_64/Y OR2X1_LOC_687/Y 0.23fF
C28684 AND2X1_LOC_593/a_8_24# AND2X1_LOC_605/Y 0.01fF
C28685 AND2X1_LOC_560/a_8_24# AND2X1_LOC_560/B 0.11fF
C28686 OR2X1_LOC_509/a_8_216# OR2X1_LOC_663/A 0.06fF
C28687 OR2X1_LOC_235/B INPUT_2 0.01fF
C28688 AND2X1_LOC_59/Y OR2X1_LOC_175/Y 0.05fF
C28689 AND2X1_LOC_714/a_8_24# AND2X1_LOC_841/B 0.20fF
C28690 OR2X1_LOC_244/Y AND2X1_LOC_245/a_8_24# 0.01fF
C28691 OR2X1_LOC_363/A OR2X1_LOC_66/A 0.01fF
C28692 AND2X1_LOC_721/A OR2X1_LOC_813/Y 0.04fF
C28693 AND2X1_LOC_39/a_8_24# OR2X1_LOC_596/A 0.01fF
C28694 OR2X1_LOC_725/B OR2X1_LOC_725/A 0.07fF
C28695 AND2X1_LOC_682/a_8_24# OR2X1_LOC_161/B 0.01fF
C28696 AND2X1_LOC_535/Y AND2X1_LOC_436/a_36_24# 0.00fF
C28697 OR2X1_LOC_40/Y AND2X1_LOC_734/Y 0.16fF
C28698 AND2X1_LOC_735/Y VDD 0.16fF
C28699 OR2X1_LOC_18/Y AND2X1_LOC_219/A 0.03fF
C28700 OR2X1_LOC_506/A OR2X1_LOC_161/B 0.21fF
C28701 AND2X1_LOC_727/A OR2X1_LOC_13/B 0.00fF
C28702 OR2X1_LOC_377/A AND2X1_LOC_277/a_8_24# 0.02fF
C28703 OR2X1_LOC_204/Y OR2X1_LOC_267/Y 0.05fF
C28704 OR2X1_LOC_503/Y AND2X1_LOC_657/A 0.01fF
C28705 AND2X1_LOC_95/Y OR2X1_LOC_344/A 0.03fF
C28706 AND2X1_LOC_59/Y OR2X1_LOC_691/Y 0.03fF
C28707 OR2X1_LOC_49/A AND2X1_LOC_43/B 0.07fF
C28708 OR2X1_LOC_39/A OR2X1_LOC_522/a_8_216# 0.03fF
C28709 AND2X1_LOC_19/Y OR2X1_LOC_78/B 0.00fF
C28710 AND2X1_LOC_695/a_8_24# OR2X1_LOC_161/B 0.01fF
C28711 OR2X1_LOC_866/B D_GATE_865 0.02fF
C28712 OR2X1_LOC_663/A OR2X1_LOC_66/A 0.03fF
C28713 OR2X1_LOC_862/B OR2X1_LOC_391/A 0.02fF
C28714 AND2X1_LOC_508/A AND2X1_LOC_658/A 0.03fF
C28715 AND2X1_LOC_542/a_8_24# OR2X1_LOC_109/Y 0.01fF
C28716 OR2X1_LOC_605/A OR2X1_LOC_605/Y 0.16fF
C28717 OR2X1_LOC_634/A OR2X1_LOC_78/A 0.70fF
C28718 AND2X1_LOC_736/Y AND2X1_LOC_565/B 0.03fF
C28719 AND2X1_LOC_302/a_8_24# OR2X1_LOC_12/Y 0.01fF
C28720 AND2X1_LOC_22/Y OR2X1_LOC_649/B 0.01fF
C28721 OR2X1_LOC_778/Y AND2X1_LOC_7/B 0.03fF
C28722 AND2X1_LOC_831/a_8_24# AND2X1_LOC_786/Y 0.02fF
C28723 AND2X1_LOC_141/a_8_24# AND2X1_LOC_141/A 0.10fF
C28724 AND2X1_LOC_303/A OR2X1_LOC_135/Y 0.09fF
C28725 AND2X1_LOC_56/B OR2X1_LOC_34/a_8_216# 0.01fF
C28726 AND2X1_LOC_555/Y AND2X1_LOC_345/Y 0.68fF
C28727 OR2X1_LOC_44/Y AND2X1_LOC_786/Y 0.07fF
C28728 AND2X1_LOC_43/B OR2X1_LOC_596/A 0.11fF
C28729 OR2X1_LOC_158/A AND2X1_LOC_624/A 0.09fF
C28730 OR2X1_LOC_95/Y OR2X1_LOC_599/a_36_216# 0.00fF
C28731 OR2X1_LOC_51/Y AND2X1_LOC_840/a_8_24# 0.01fF
C28732 OR2X1_LOC_346/B AND2X1_LOC_44/Y 0.01fF
C28733 OR2X1_LOC_502/A AND2X1_LOC_92/Y 0.14fF
C28734 AND2X1_LOC_530/a_8_24# AND2X1_LOC_56/B 0.17fF
C28735 OR2X1_LOC_95/Y OR2X1_LOC_13/B 0.12fF
C28736 AND2X1_LOC_535/Y AND2X1_LOC_356/a_8_24# 0.00fF
C28737 AND2X1_LOC_218/a_8_24# OR2X1_LOC_18/Y 0.05fF
C28738 OR2X1_LOC_505/Y OR2X1_LOC_18/Y 0.01fF
C28739 AND2X1_LOC_560/a_8_24# OR2X1_LOC_64/Y 0.01fF
C28740 OR2X1_LOC_771/a_8_216# OR2X1_LOC_68/B 0.01fF
C28741 OR2X1_LOC_770/Y OR2X1_LOC_80/A 0.01fF
C28742 OR2X1_LOC_641/Y OR2X1_LOC_655/a_8_216# 0.02fF
C28743 OR2X1_LOC_647/A AND2X1_LOC_7/B 0.14fF
C28744 AND2X1_LOC_707/Y OR2X1_LOC_743/A 0.06fF
C28745 GATE_811 AND2X1_LOC_740/a_8_24# 0.01fF
C28746 OR2X1_LOC_600/a_8_216# AND2X1_LOC_593/Y 0.06fF
C28747 AND2X1_LOC_647/Y OR2X1_LOC_88/Y 0.35fF
C28748 AND2X1_LOC_658/A OR2X1_LOC_18/Y 0.16fF
C28749 OR2X1_LOC_475/Y OR2X1_LOC_392/B 0.08fF
C28750 AND2X1_LOC_64/Y OR2X1_LOC_401/B 0.29fF
C28751 AND2X1_LOC_91/B OR2X1_LOC_401/A 0.03fF
C28752 AND2X1_LOC_444/a_8_24# AND2X1_LOC_804/Y 0.01fF
C28753 AND2X1_LOC_56/B OR2X1_LOC_542/a_8_216# 0.01fF
C28754 OR2X1_LOC_672/a_8_216# OR2X1_LOC_43/A 0.03fF
C28755 OR2X1_LOC_17/Y OR2X1_LOC_428/A 0.03fF
C28756 OR2X1_LOC_604/A OR2X1_LOC_603/a_36_216# 0.00fF
C28757 OR2X1_LOC_856/B AND2X1_LOC_41/A 0.13fF
C28758 AND2X1_LOC_122/a_8_24# AND2X1_LOC_44/Y 0.04fF
C28759 AND2X1_LOC_392/a_8_24# OR2X1_LOC_278/Y 0.01fF
C28760 AND2X1_LOC_367/A AND2X1_LOC_76/Y 0.03fF
C28761 OR2X1_LOC_314/a_8_216# OR2X1_LOC_683/a_8_216# 0.47fF
C28762 OR2X1_LOC_100/Y AND2X1_LOC_40/Y 0.04fF
C28763 AND2X1_LOC_131/a_36_24# OR2X1_LOC_203/Y 0.01fF
C28764 OR2X1_LOC_696/A AND2X1_LOC_801/B 0.01fF
C28765 AND2X1_LOC_95/Y OR2X1_LOC_410/a_36_216# -0.00fF
C28766 OR2X1_LOC_186/Y OR2X1_LOC_479/Y 0.07fF
C28767 OR2X1_LOC_51/Y OR2X1_LOC_511/Y 0.01fF
C28768 OR2X1_LOC_91/A AND2X1_LOC_661/a_36_24# 0.00fF
C28769 OR2X1_LOC_185/Y OR2X1_LOC_66/A 0.08fF
C28770 OR2X1_LOC_69/A OR2X1_LOC_59/Y 0.02fF
C28771 OR2X1_LOC_154/A OR2X1_LOC_244/Y 0.15fF
C28772 AND2X1_LOC_842/B OR2X1_LOC_530/a_8_216# 0.47fF
C28773 OR2X1_LOC_189/Y AND2X1_LOC_477/Y 0.07fF
C28774 OR2X1_LOC_364/A OR2X1_LOC_841/A 0.01fF
C28775 AND2X1_LOC_861/a_36_24# AND2X1_LOC_807/Y 0.00fF
C28776 AND2X1_LOC_3/Y OR2X1_LOC_719/B 0.22fF
C28777 AND2X1_LOC_858/B OR2X1_LOC_39/A 0.26fF
C28778 OR2X1_LOC_864/A AND2X1_LOC_18/Y 0.13fF
C28779 AND2X1_LOC_592/Y OR2X1_LOC_89/A 0.00fF
C28780 OR2X1_LOC_208/A OR2X1_LOC_532/B 0.01fF
C28781 OR2X1_LOC_91/A OR2X1_LOC_39/A 0.07fF
C28782 AND2X1_LOC_580/A OR2X1_LOC_56/A 0.07fF
C28783 AND2X1_LOC_584/a_8_24# AND2X1_LOC_70/Y 0.01fF
C28784 OR2X1_LOC_351/B OR2X1_LOC_333/B 0.03fF
C28785 OR2X1_LOC_91/Y OR2X1_LOC_329/B 0.07fF
C28786 OR2X1_LOC_154/A OR2X1_LOC_715/A 0.02fF
C28787 OR2X1_LOC_18/Y AND2X1_LOC_139/a_8_24# 0.03fF
C28788 AND2X1_LOC_767/a_8_24# OR2X1_LOC_756/B 0.01fF
C28789 AND2X1_LOC_663/B OR2X1_LOC_12/Y 0.03fF
C28790 OR2X1_LOC_653/Y OR2X1_LOC_61/B -0.01fF
C28791 AND2X1_LOC_367/A OR2X1_LOC_67/A 0.05fF
C28792 OR2X1_LOC_821/a_8_216# OR2X1_LOC_64/Y 0.01fF
C28793 OR2X1_LOC_147/B OR2X1_LOC_620/Y 0.03fF
C28794 OR2X1_LOC_62/A AND2X1_LOC_619/a_36_24# 0.01fF
C28795 AND2X1_LOC_347/B AND2X1_LOC_347/a_8_24# 0.04fF
C28796 AND2X1_LOC_40/Y OR2X1_LOC_286/Y 0.02fF
C28797 AND2X1_LOC_772/B OR2X1_LOC_26/Y 0.01fF
C28798 OR2X1_LOC_633/B AND2X1_LOC_18/Y 0.03fF
C28799 OR2X1_LOC_847/A AND2X1_LOC_619/B 0.01fF
C28800 OR2X1_LOC_673/Y OR2X1_LOC_78/B 0.07fF
C28801 AND2X1_LOC_702/Y OR2X1_LOC_59/Y 0.04fF
C28802 OR2X1_LOC_185/Y AND2X1_LOC_311/a_8_24# 0.00fF
C28803 OR2X1_LOC_648/A OR2X1_LOC_449/B 0.05fF
C28804 AND2X1_LOC_715/Y AND2X1_LOC_801/B 0.00fF
C28805 AND2X1_LOC_95/Y OR2X1_LOC_575/A 0.51fF
C28806 OR2X1_LOC_493/A OR2X1_LOC_737/A 0.23fF
C28807 OR2X1_LOC_542/B AND2X1_LOC_3/Y 0.03fF
C28808 OR2X1_LOC_329/Y OR2X1_LOC_70/Y 0.02fF
C28809 AND2X1_LOC_686/a_8_24# OR2X1_LOC_12/Y 0.01fF
C28810 OR2X1_LOC_849/A AND2X1_LOC_103/a_8_24# -0.00fF
C28811 OR2X1_LOC_427/A OR2X1_LOC_278/Y 0.06fF
C28812 OR2X1_LOC_702/A OR2X1_LOC_160/B 0.72fF
C28813 AND2X1_LOC_729/B AND2X1_LOC_193/Y 0.01fF
C28814 AND2X1_LOC_772/B OR2X1_LOC_89/A 0.02fF
C28815 OR2X1_LOC_8/Y OR2X1_LOC_74/A 0.04fF
C28816 OR2X1_LOC_7/A OR2X1_LOC_743/a_8_216# 0.04fF
C28817 OR2X1_LOC_97/A OR2X1_LOC_544/A 0.32fF
C28818 OR2X1_LOC_814/A OR2X1_LOC_435/A 0.04fF
C28819 OR2X1_LOC_633/a_36_216# AND2X1_LOC_8/Y 0.01fF
C28820 AND2X1_LOC_368/a_8_24# OR2X1_LOC_465/B 0.01fF
C28821 AND2X1_LOC_512/Y OR2X1_LOC_26/Y 0.07fF
C28822 AND2X1_LOC_211/B OR2X1_LOC_91/A 0.19fF
C28823 OR2X1_LOC_265/a_8_216# OR2X1_LOC_85/A 0.01fF
C28824 OR2X1_LOC_505/a_8_216# OR2X1_LOC_504/Y 0.01fF
C28825 AND2X1_LOC_64/Y OR2X1_LOC_786/Y 0.11fF
C28826 OR2X1_LOC_673/Y OR2X1_LOC_721/Y 0.01fF
C28827 AND2X1_LOC_116/Y AND2X1_LOC_218/Y 0.01fF
C28828 OR2X1_LOC_780/A OR2X1_LOC_161/B 0.04fF
C28829 OR2X1_LOC_624/A OR2X1_LOC_161/A 0.05fF
C28830 OR2X1_LOC_673/B OR2X1_LOC_532/B 0.03fF
C28831 AND2X1_LOC_94/Y AND2X1_LOC_42/B 0.02fF
C28832 AND2X1_LOC_367/a_36_24# OR2X1_LOC_92/Y 0.00fF
C28833 OR2X1_LOC_837/A OR2X1_LOC_6/A 0.14fF
C28834 AND2X1_LOC_95/Y OR2X1_LOC_652/a_8_216# 0.01fF
C28835 VDD OR2X1_LOC_52/Y 0.23fF
C28836 OR2X1_LOC_319/B OR2X1_LOC_778/Y 0.10fF
C28837 OR2X1_LOC_160/B OR2X1_LOC_476/B 0.07fF
C28838 AND2X1_LOC_489/Y AND2X1_LOC_367/A 0.05fF
C28839 AND2X1_LOC_675/A OR2X1_LOC_373/Y 0.11fF
C28840 AND2X1_LOC_573/A OR2X1_LOC_39/A 0.43fF
C28841 OR2X1_LOC_806/a_8_216# OR2X1_LOC_807/A 0.01fF
C28842 OR2X1_LOC_589/A OR2X1_LOC_71/Y 0.00fF
C28843 VDD OR2X1_LOC_750/A 0.25fF
C28844 AND2X1_LOC_3/Y OR2X1_LOC_736/A 0.10fF
C28845 OR2X1_LOC_481/A OR2X1_LOC_297/A 0.00fF
C28846 OR2X1_LOC_585/A OR2X1_LOC_586/a_8_216# 0.01fF
C28847 AND2X1_LOC_123/Y AND2X1_LOC_124/a_8_24# 0.01fF
C28848 OR2X1_LOC_329/B OR2X1_LOC_527/Y 0.02fF
C28849 OR2X1_LOC_790/A AND2X1_LOC_53/Y 0.11fF
C28850 OR2X1_LOC_768/A OR2X1_LOC_404/Y 0.03fF
C28851 OR2X1_LOC_612/a_36_216# OR2X1_LOC_62/B 0.00fF
C28852 AND2X1_LOC_554/B OR2X1_LOC_256/Y 0.02fF
C28853 OR2X1_LOC_620/Y AND2X1_LOC_298/a_36_24# 0.00fF
C28854 INPUT_5 OR2X1_LOC_47/a_36_216# 0.02fF
C28855 AND2X1_LOC_486/Y OR2X1_LOC_238/Y 0.10fF
C28856 OR2X1_LOC_135/Y AND2X1_LOC_655/a_8_24# 0.01fF
C28857 OR2X1_LOC_630/a_36_216# OR2X1_LOC_631/B 0.00fF
C28858 VDD OR2X1_LOC_168/A -0.00fF
C28859 AND2X1_LOC_518/a_8_24# AND2X1_LOC_92/Y 0.01fF
C28860 AND2X1_LOC_51/A AND2X1_LOC_11/Y 0.12fF
C28861 AND2X1_LOC_420/a_8_24# OR2X1_LOC_161/B 0.02fF
C28862 OR2X1_LOC_680/A OR2X1_LOC_511/Y 0.01fF
C28863 AND2X1_LOC_131/a_8_24# OR2X1_LOC_532/B 0.03fF
C28864 AND2X1_LOC_76/a_36_24# OR2X1_LOC_52/B 0.01fF
C28865 OR2X1_LOC_448/Y OR2X1_LOC_87/A 0.14fF
C28866 AND2X1_LOC_8/Y AND2X1_LOC_104/a_8_24# 0.09fF
C28867 VDD OR2X1_LOC_611/Y 0.00fF
C28868 OR2X1_LOC_664/Y OR2X1_LOC_483/a_8_216# 0.44fF
C28869 AND2X1_LOC_71/a_8_24# OR2X1_LOC_404/Y 0.01fF
C28870 OR2X1_LOC_673/Y OR2X1_LOC_375/A 0.03fF
C28871 OR2X1_LOC_161/B D_INPUT_1 0.07fF
C28872 AND2X1_LOC_817/B AND2X1_LOC_382/a_8_24# 0.00fF
C28873 OR2X1_LOC_329/B OR2X1_LOC_311/Y 0.03fF
C28874 AND2X1_LOC_599/a_8_24# OR2X1_LOC_644/A 0.01fF
C28875 AND2X1_LOC_48/A AND2X1_LOC_92/Y 0.07fF
C28876 OR2X1_LOC_631/a_8_216# AND2X1_LOC_3/Y 0.02fF
C28877 OR2X1_LOC_516/A OR2X1_LOC_26/Y 0.03fF
C28878 OR2X1_LOC_185/A OR2X1_LOC_643/a_8_216# 0.01fF
C28879 OR2X1_LOC_777/B OR2X1_LOC_788/B 0.03fF
C28880 OR2X1_LOC_641/B AND2X1_LOC_226/a_8_24# 0.01fF
C28881 AND2X1_LOC_76/Y OR2X1_LOC_74/A 0.04fF
C28882 OR2X1_LOC_599/A AND2X1_LOC_319/A 0.21fF
C28883 OR2X1_LOC_805/A OR2X1_LOC_778/Y 0.11fF
C28884 OR2X1_LOC_69/a_8_216# OR2X1_LOC_69/Y 0.02fF
C28885 OR2X1_LOC_596/Y AND2X1_LOC_597/a_8_24# 0.23fF
C28886 AND2X1_LOC_413/a_8_24# OR2X1_LOC_461/A 0.01fF
C28887 AND2X1_LOC_191/Y AND2X1_LOC_807/a_8_24# 0.07fF
C28888 AND2X1_LOC_40/Y AND2X1_LOC_670/a_36_24# 0.00fF
C28889 OR2X1_LOC_436/B OR2X1_LOC_436/a_8_216# 0.02fF
C28890 OR2X1_LOC_457/a_8_216# OR2X1_LOC_464/B -0.00fF
C28891 AND2X1_LOC_35/Y OR2X1_LOC_52/B 0.39fF
C28892 VDD OR2X1_LOC_689/Y 0.12fF
C28893 AND2X1_LOC_480/a_8_24# AND2X1_LOC_480/A 0.01fF
C28894 AND2X1_LOC_477/A AND2X1_LOC_471/Y 0.16fF
C28895 AND2X1_LOC_52/a_36_24# AND2X1_LOC_51/Y 0.01fF
C28896 OR2X1_LOC_6/A OR2X1_LOC_49/a_8_216# 0.01fF
C28897 OR2X1_LOC_856/B AND2X1_LOC_135/a_8_24# 0.01fF
C28898 OR2X1_LOC_223/A OR2X1_LOC_787/a_36_216# 0.00fF
C28899 VDD OR2X1_LOC_503/Y 0.16fF
C28900 OR2X1_LOC_670/Y OR2X1_LOC_6/A 0.01fF
C28901 AND2X1_LOC_12/Y OR2X1_LOC_333/B 0.06fF
C28902 OR2X1_LOC_682/a_8_216# OR2X1_LOC_36/Y 0.18fF
C28903 AND2X1_LOC_349/B AND2X1_LOC_342/Y 0.00fF
C28904 OR2X1_LOC_485/A AND2X1_LOC_848/Y 0.03fF
C28905 AND2X1_LOC_584/a_8_24# AND2X1_LOC_17/Y 0.09fF
C28906 AND2X1_LOC_12/Y OR2X1_LOC_850/A 0.08fF
C28907 OR2X1_LOC_69/a_36_216# OR2X1_LOC_52/B -0.00fF
C28908 OR2X1_LOC_107/a_36_216# AND2X1_LOC_227/Y 0.00fF
C28909 OR2X1_LOC_763/Y OR2X1_LOC_44/Y 0.04fF
C28910 AND2X1_LOC_476/A OR2X1_LOC_56/A 0.42fF
C28911 AND2X1_LOC_56/B AND2X1_LOC_3/Y 0.13fF
C28912 AND2X1_LOC_105/a_8_24# OR2X1_LOC_26/Y 0.03fF
C28913 D_INPUT_7 AND2X1_LOC_17/a_8_24# 0.01fF
C28914 OR2X1_LOC_542/B OR2X1_LOC_270/Y 0.03fF
C28915 OR2X1_LOC_92/Y AND2X1_LOC_687/Y 0.02fF
C28916 OR2X1_LOC_602/a_8_216# OR2X1_LOC_602/A 0.47fF
C28917 OR2X1_LOC_36/Y OR2X1_LOC_609/a_8_216# 0.02fF
C28918 AND2X1_LOC_741/Y AND2X1_LOC_223/a_8_24# 0.00fF
C28919 OR2X1_LOC_600/A OR2X1_LOC_29/a_8_216# 0.05fF
C28920 VDD OR2X1_LOC_2/a_8_216# 0.21fF
C28921 AND2X1_LOC_662/a_8_24# OR2X1_LOC_39/A 0.03fF
C28922 OR2X1_LOC_631/B OR2X1_LOC_296/a_36_216# 0.00fF
C28923 OR2X1_LOC_672/Y AND2X1_LOC_673/a_8_24# 0.00fF
C28924 AND2X1_LOC_658/A AND2X1_LOC_620/Y 1.09fF
C28925 OR2X1_LOC_481/a_8_216# OR2X1_LOC_44/Y 0.01fF
C28926 AND2X1_LOC_8/Y OR2X1_LOC_647/B 0.07fF
C28927 AND2X1_LOC_343/a_8_24# OR2X1_LOC_106/A 0.09fF
C28928 AND2X1_LOC_40/Y OR2X1_LOC_532/B 0.26fF
C28929 AND2X1_LOC_105/a_8_24# OR2X1_LOC_89/A 0.09fF
C28930 OR2X1_LOC_19/B OR2X1_LOC_63/a_8_216# 0.02fF
C28931 OR2X1_LOC_696/A OR2X1_LOC_248/A 0.13fF
C28932 AND2X1_LOC_328/a_8_24# AND2X1_LOC_7/Y 0.00fF
C28933 OR2X1_LOC_74/A OR2X1_LOC_52/B 1.42fF
C28934 OR2X1_LOC_654/A AND2X1_LOC_822/a_8_24# 0.05fF
C28935 OR2X1_LOC_632/A OR2X1_LOC_62/B 0.01fF
C28936 OR2X1_LOC_533/Y OR2X1_LOC_533/A 0.04fF
C28937 OR2X1_LOC_802/a_8_216# OR2X1_LOC_436/Y 0.01fF
C28938 OR2X1_LOC_715/B AND2X1_LOC_679/a_36_24# 0.01fF
C28939 AND2X1_LOC_141/B OR2X1_LOC_26/Y 0.19fF
C28940 OR2X1_LOC_43/A OR2X1_LOC_481/A 0.07fF
C28941 OR2X1_LOC_32/B OR2X1_LOC_22/Y 0.09fF
C28942 OR2X1_LOC_31/Y OR2X1_LOC_2/Y 0.01fF
C28943 OR2X1_LOC_548/A OR2X1_LOC_80/A 0.05fF
C28944 AND2X1_LOC_324/a_36_24# OR2X1_LOC_36/Y 0.00fF
C28945 OR2X1_LOC_400/B AND2X1_LOC_51/Y 0.01fF
C28946 AND2X1_LOC_489/Y OR2X1_LOC_490/Y 0.02fF
C28947 AND2X1_LOC_59/Y OR2X1_LOC_750/a_8_216# 0.06fF
C28948 OR2X1_LOC_502/A D_INPUT_3 3.76fF
C28949 OR2X1_LOC_280/Y OR2X1_LOC_371/Y 0.07fF
C28950 AND2X1_LOC_425/Y OR2X1_LOC_375/A 0.01fF
C28951 OR2X1_LOC_8/Y AND2X1_LOC_647/Y 0.01fF
C28952 AND2X1_LOC_31/Y OR2X1_LOC_307/A 0.01fF
C28953 OR2X1_LOC_641/A OR2X1_LOC_228/Y 0.00fF
C28954 AND2X1_LOC_309/a_8_24# OR2X1_LOC_375/A 0.01fF
C28955 AND2X1_LOC_42/a_36_24# AND2X1_LOC_42/B 0.01fF
C28956 OR2X1_LOC_447/Y OR2X1_LOC_161/A 0.07fF
C28957 OR2X1_LOC_537/A OR2X1_LOC_532/B 0.01fF
C28958 AND2X1_LOC_141/B OR2X1_LOC_89/A 0.21fF
C28959 VDD OR2X1_LOC_754/Y 0.16fF
C28960 AND2X1_LOC_22/Y OR2X1_LOC_777/B 0.03fF
C28961 AND2X1_LOC_340/a_8_24# OR2X1_LOC_88/Y 0.01fF
C28962 OR2X1_LOC_508/Y OR2X1_LOC_510/a_36_216# 0.02fF
C28963 OR2X1_LOC_344/A OR2X1_LOC_269/A 0.01fF
C28964 VDD OR2X1_LOC_742/B 0.17fF
C28965 AND2X1_LOC_132/a_8_24# AND2X1_LOC_47/Y 0.02fF
C28966 OR2X1_LOC_26/Y OR2X1_LOC_54/Y 0.08fF
C28967 OR2X1_LOC_529/a_36_216# AND2X1_LOC_227/Y 0.00fF
C28968 OR2X1_LOC_267/a_8_216# OR2X1_LOC_814/A 0.06fF
C28969 OR2X1_LOC_476/B OR2X1_LOC_219/B 0.07fF
C28970 AND2X1_LOC_276/Y AND2X1_LOC_473/a_36_24# 0.01fF
C28971 OR2X1_LOC_630/B OR2X1_LOC_598/A 0.02fF
C28972 OR2X1_LOC_66/A OR2X1_LOC_568/A 0.07fF
C28973 AND2X1_LOC_2/Y AND2X1_LOC_430/B 0.02fF
C28974 AND2X1_LOC_631/a_8_24# AND2X1_LOC_620/Y 0.01fF
C28975 OR2X1_LOC_748/A INPUT_1 0.06fF
C28976 AND2X1_LOC_796/Y AND2X1_LOC_621/Y 0.03fF
C28977 OR2X1_LOC_66/A OR2X1_LOC_578/B 0.00fF
C28978 OR2X1_LOC_357/B OR2X1_LOC_212/B 0.01fF
C28979 OR2X1_LOC_244/Y OR2X1_LOC_560/A 0.02fF
C28980 OR2X1_LOC_272/Y AND2X1_LOC_663/B 0.01fF
C28981 AND2X1_LOC_310/a_8_24# OR2X1_LOC_68/B 0.03fF
C28982 OR2X1_LOC_89/A OR2X1_LOC_54/Y 0.02fF
C28983 AND2X1_LOC_44/Y OR2X1_LOC_469/B 0.03fF
C28984 AND2X1_LOC_349/a_8_24# OR2X1_LOC_256/A 0.23fF
C28985 OR2X1_LOC_43/A OR2X1_LOC_71/Y 0.03fF
C28986 OR2X1_LOC_446/Y OR2X1_LOC_449/A 0.47fF
C28987 AND2X1_LOC_227/Y AND2X1_LOC_361/A 0.01fF
C28988 OR2X1_LOC_846/a_8_216# D_INPUT_1 0.01fF
C28989 AND2X1_LOC_722/A OR2X1_LOC_331/Y 0.07fF
C28990 AND2X1_LOC_64/Y AND2X1_LOC_829/a_8_24# 0.01fF
C28991 AND2X1_LOC_47/Y OR2X1_LOC_564/B 0.01fF
C28992 OR2X1_LOC_276/B OR2X1_LOC_269/B 0.25fF
C28993 AND2X1_LOC_737/Y AND2X1_LOC_222/Y 0.48fF
C28994 OR2X1_LOC_114/Y OR2X1_LOC_473/A 0.00fF
C28995 AND2X1_LOC_91/B AND2X1_LOC_7/B 0.16fF
C28996 AND2X1_LOC_22/Y OR2X1_LOC_831/B 0.03fF
C28997 AND2X1_LOC_56/B OR2X1_LOC_270/Y 0.06fF
C28998 OR2X1_LOC_165/a_8_216# AND2X1_LOC_222/Y 0.01fF
C28999 OR2X1_LOC_139/A OR2X1_LOC_390/a_8_216# 0.05fF
C29000 AND2X1_LOC_272/a_8_24# OR2X1_LOC_493/Y 0.05fF
C29001 OR2X1_LOC_620/Y OR2X1_LOC_854/A 0.02fF
C29002 AND2X1_LOC_12/Y OR2X1_LOC_590/a_8_216# 0.01fF
C29003 OR2X1_LOC_43/A D_INPUT_1 0.12fF
C29004 OR2X1_LOC_49/A AND2X1_LOC_416/a_8_24# 0.01fF
C29005 OR2X1_LOC_189/Y GATE_811 0.03fF
C29006 AND2X1_LOC_56/B OR2X1_LOC_194/a_8_216# 0.01fF
C29007 OR2X1_LOC_600/A AND2X1_LOC_793/a_8_24# 0.01fF
C29008 OR2X1_LOC_261/a_8_216# AND2X1_LOC_789/Y 0.01fF
C29009 AND2X1_LOC_64/Y OR2X1_LOC_535/A 0.01fF
C29010 OR2X1_LOC_510/A OR2X1_LOC_510/a_8_216# 0.06fF
C29011 OR2X1_LOC_152/Y GATE_811 0.02fF
C29012 AND2X1_LOC_566/Y OR2X1_LOC_47/Y 0.12fF
C29013 OR2X1_LOC_53/Y AND2X1_LOC_195/a_8_24# 0.01fF
C29014 OR2X1_LOC_599/A AND2X1_LOC_644/a_36_24# 0.00fF
C29015 OR2X1_LOC_12/a_8_216# D_INPUT_6 0.01fF
C29016 OR2X1_LOC_45/B AND2X1_LOC_786/Y 0.14fF
C29017 OR2X1_LOC_297/A AND2X1_LOC_789/Y 0.02fF
C29018 AND2X1_LOC_628/a_8_24# AND2X1_LOC_36/Y 0.01fF
C29019 OR2X1_LOC_59/Y AND2X1_LOC_792/B 0.01fF
C29020 OR2X1_LOC_580/a_8_216# OR2X1_LOC_269/B 0.01fF
C29021 OR2X1_LOC_756/B OR2X1_LOC_576/a_36_216# 0.00fF
C29022 OR2X1_LOC_468/Y OR2X1_LOC_170/Y 0.01fF
C29023 AND2X1_LOC_81/B OR2X1_LOC_68/B 0.00fF
C29024 AND2X1_LOC_42/B OR2X1_LOC_241/B 0.05fF
C29025 OR2X1_LOC_31/Y OR2X1_LOC_7/Y 0.23fF
C29026 AND2X1_LOC_212/A OR2X1_LOC_428/A 0.03fF
C29027 OR2X1_LOC_36/Y AND2X1_LOC_657/A 0.07fF
C29028 AND2X1_LOC_721/Y AND2X1_LOC_778/Y 0.01fF
C29029 VDD OR2X1_LOC_748/Y 0.12fF
C29030 OR2X1_LOC_206/A OR2X1_LOC_786/Y 0.13fF
C29031 OR2X1_LOC_425/a_8_216# D_INPUT_6 0.01fF
C29032 AND2X1_LOC_729/a_8_24# OR2X1_LOC_16/A 0.01fF
C29033 OR2X1_LOC_269/B OR2X1_LOC_779/B 0.03fF
C29034 AND2X1_LOC_18/Y OR2X1_LOC_121/A 0.09fF
C29035 AND2X1_LOC_95/Y OR2X1_LOC_735/B 0.01fF
C29036 OR2X1_LOC_220/A OR2X1_LOC_209/A 0.03fF
C29037 OR2X1_LOC_53/Y AND2X1_LOC_199/a_36_24# -0.00fF
C29038 OR2X1_LOC_604/A GATE_579 0.00fF
C29039 OR2X1_LOC_51/Y AND2X1_LOC_465/A 0.09fF
C29040 AND2X1_LOC_758/a_8_24# GATE_579 0.01fF
C29041 OR2X1_LOC_417/A AND2X1_LOC_859/B 0.02fF
C29042 OR2X1_LOC_756/B OR2X1_LOC_388/a_36_216# -0.00fF
C29043 OR2X1_LOC_710/A OR2X1_LOC_147/A 0.09fF
C29044 OR2X1_LOC_630/Y OR2X1_LOC_554/a_8_216# 0.02fF
C29045 AND2X1_LOC_170/B AND2X1_LOC_866/A 0.01fF
C29046 AND2X1_LOC_3/Y AND2X1_LOC_427/a_8_24# 0.02fF
C29047 OR2X1_LOC_612/a_8_216# OR2X1_LOC_16/A -0.00fF
C29048 OR2X1_LOC_78/A OR2X1_LOC_267/Y 0.13fF
C29049 AND2X1_LOC_430/a_8_24# OR2X1_LOC_451/B 0.01fF
C29050 AND2X1_LOC_392/A OR2X1_LOC_12/Y 0.03fF
C29051 OR2X1_LOC_600/A OR2X1_LOC_16/A 11.19fF
C29052 AND2X1_LOC_364/a_8_24# OR2X1_LOC_426/B 0.00fF
C29053 OR2X1_LOC_696/A OR2X1_LOC_59/a_8_216# 0.01fF
C29054 OR2X1_LOC_45/B AND2X1_LOC_218/Y 0.03fF
C29055 OR2X1_LOC_375/A OR2X1_LOC_723/B 2.75fF
C29056 D_INPUT_3 OR2X1_LOC_618/Y 0.01fF
C29057 AND2X1_LOC_479/Y AND2X1_LOC_480/a_8_24# 0.11fF
C29058 AND2X1_LOC_91/B OR2X1_LOC_319/B 0.07fF
C29059 OR2X1_LOC_166/a_8_216# OR2X1_LOC_16/A 0.02fF
C29060 OR2X1_LOC_6/B AND2X1_LOC_625/a_8_24# 0.02fF
C29061 OR2X1_LOC_45/B OR2X1_LOC_524/Y 0.01fF
C29062 AND2X1_LOC_663/A AND2X1_LOC_213/B 0.05fF
C29063 OR2X1_LOC_709/A OR2X1_LOC_702/a_8_216# 0.01fF
C29064 AND2X1_LOC_51/Y OR2X1_LOC_513/a_8_216# 0.02fF
C29065 OR2X1_LOC_78/A OR2X1_LOC_633/A 0.14fF
C29066 OR2X1_LOC_711/B VDD 0.06fF
C29067 OR2X1_LOC_56/a_8_216# OR2X1_LOC_16/Y 0.40fF
C29068 AND2X1_LOC_64/Y OR2X1_LOC_851/A 0.00fF
C29069 AND2X1_LOC_541/Y AND2X1_LOC_563/A 0.02fF
C29070 OR2X1_LOC_585/A OR2X1_LOC_536/a_36_216# 0.00fF
C29071 OR2X1_LOC_198/a_8_216# AND2X1_LOC_95/Y 0.02fF
C29072 OR2X1_LOC_589/A OR2X1_LOC_426/B 0.03fF
C29073 OR2X1_LOC_323/A OR2X1_LOC_427/A 0.05fF
C29074 OR2X1_LOC_720/Y OR2X1_LOC_721/Y -0.01fF
C29075 AND2X1_LOC_866/A AND2X1_LOC_721/A 0.03fF
C29076 OR2X1_LOC_485/A OR2X1_LOC_536/a_8_216# 0.00fF
C29077 OR2X1_LOC_22/Y AND2X1_LOC_222/Y 0.01fF
C29078 AND2X1_LOC_70/Y OR2X1_LOC_786/a_8_216# 0.01fF
C29079 OR2X1_LOC_427/A OR2X1_LOC_89/Y 0.03fF
C29080 OR2X1_LOC_43/A AND2X1_LOC_789/Y 0.52fF
C29081 AND2X1_LOC_64/Y OR2X1_LOC_220/B 0.02fF
C29082 OR2X1_LOC_108/Y OR2X1_LOC_600/A 0.24fF
C29083 AND2X1_LOC_715/Y AND2X1_LOC_703/a_8_24# 0.03fF
C29084 OR2X1_LOC_22/Y OR2X1_LOC_68/B 0.03fF
C29085 AND2X1_LOC_716/Y AND2X1_LOC_358/Y 0.00fF
C29086 AND2X1_LOC_150/a_8_24# OR2X1_LOC_244/B 0.01fF
C29087 OR2X1_LOC_691/Y OR2X1_LOC_623/B 0.03fF
C29088 OR2X1_LOC_865/A OR2X1_LOC_810/a_8_216# 0.01fF
C29089 OR2X1_LOC_862/a_8_216# OR2X1_LOC_812/B 0.01fF
C29090 AND2X1_LOC_69/a_8_24# AND2X1_LOC_31/Y 0.01fF
C29091 VDD OR2X1_LOC_347/Y 0.00fF
C29092 OR2X1_LOC_335/A OR2X1_LOC_375/A 0.01fF
C29093 OR2X1_LOC_97/A OR2X1_LOC_653/Y 0.01fF
C29094 VDD AND2X1_LOC_404/B 0.02fF
C29095 AND2X1_LOC_64/Y OR2X1_LOC_828/B 0.23fF
C29096 OR2X1_LOC_557/A OR2X1_LOC_771/B 0.03fF
C29097 OR2X1_LOC_468/Y OR2X1_LOC_168/Y 0.02fF
C29098 AND2X1_LOC_153/a_8_24# OR2X1_LOC_831/B 0.03fF
C29099 AND2X1_LOC_91/B OR2X1_LOC_805/A 0.10fF
C29100 OR2X1_LOC_323/A AND2X1_LOC_464/a_8_24# 0.00fF
C29101 AND2X1_LOC_72/Y AND2X1_LOC_7/B 0.02fF
C29102 OR2X1_LOC_793/B AND2X1_LOC_36/Y 0.21fF
C29103 AND2X1_LOC_842/B OR2X1_LOC_437/A 0.01fF
C29104 OR2X1_LOC_623/B OR2X1_LOC_713/A 0.15fF
C29105 OR2X1_LOC_45/Y OR2X1_LOC_428/A 0.09fF
C29106 OR2X1_LOC_40/Y OR2X1_LOC_235/B 0.07fF
C29107 AND2X1_LOC_2/Y AND2X1_LOC_70/Y 0.01fF
C29108 AND2X1_LOC_64/Y OR2X1_LOC_835/B 0.92fF
C29109 AND2X1_LOC_787/A OR2X1_LOC_109/Y 0.02fF
C29110 AND2X1_LOC_505/a_36_24# OR2X1_LOC_78/B 0.00fF
C29111 AND2X1_LOC_573/A AND2X1_LOC_456/a_8_24# 0.04fF
C29112 OR2X1_LOC_323/A OR2X1_LOC_271/a_8_216# 0.01fF
C29113 OR2X1_LOC_47/Y OR2X1_LOC_406/A 0.01fF
C29114 OR2X1_LOC_62/B OR2X1_LOC_71/A 2.24fF
C29115 VDD OR2X1_LOC_324/B 0.00fF
C29116 AND2X1_LOC_721/Y AND2X1_LOC_624/A 0.03fF
C29117 OR2X1_LOC_790/A OR2X1_LOC_502/A 0.01fF
C29118 AND2X1_LOC_95/Y OR2X1_LOC_161/B 3.67fF
C29119 AND2X1_LOC_22/Y OR2X1_LOC_652/a_8_216# 0.01fF
C29120 AND2X1_LOC_711/Y AND2X1_LOC_792/B 0.01fF
C29121 AND2X1_LOC_40/Y D_GATE_811 0.01fF
C29122 OR2X1_LOC_690/a_36_216# OR2X1_LOC_585/A 0.00fF
C29123 OR2X1_LOC_318/A OR2X1_LOC_185/A 0.02fF
C29124 OR2X1_LOC_122/A OR2X1_LOC_56/A 0.04fF
C29125 OR2X1_LOC_128/B AND2X1_LOC_44/Y 0.00fF
C29126 OR2X1_LOC_619/Y OR2X1_LOC_16/A 0.13fF
C29127 AND2X1_LOC_710/a_8_24# OR2X1_LOC_428/A 0.08fF
C29128 INPUT_0 OR2X1_LOC_56/A 0.09fF
C29129 AND2X1_LOC_47/Y OR2X1_LOC_365/a_8_216# 0.00fF
C29130 OR2X1_LOC_482/Y AND2X1_LOC_833/a_8_24# 0.10fF
C29131 OR2X1_LOC_744/A OR2X1_LOC_25/Y 0.26fF
C29132 OR2X1_LOC_51/B OR2X1_LOC_70/A 0.16fF
C29133 OR2X1_LOC_247/Y AND2X1_LOC_72/B 0.02fF
C29134 AND2X1_LOC_727/A OR2X1_LOC_142/a_8_216# 0.01fF
C29135 OR2X1_LOC_497/Y AND2X1_LOC_242/B 0.51fF
C29136 OR2X1_LOC_115/a_8_216# OR2X1_LOC_549/A 0.03fF
C29137 OR2X1_LOC_812/B OR2X1_LOC_812/a_8_216# 0.04fF
C29138 OR2X1_LOC_375/A AND2X1_LOC_277/a_8_24# 0.01fF
C29139 AND2X1_LOC_40/Y OR2X1_LOC_440/B 0.05fF
C29140 OR2X1_LOC_139/A OR2X1_LOC_203/Y 0.10fF
C29141 OR2X1_LOC_95/Y OR2X1_LOC_533/a_8_216# 0.07fF
C29142 AND2X1_LOC_848/A AND2X1_LOC_793/Y 0.85fF
C29143 OR2X1_LOC_865/A OR2X1_LOC_859/B 0.15fF
C29144 AND2X1_LOC_724/a_8_24# OR2X1_LOC_601/Y 0.24fF
C29145 AND2X1_LOC_52/a_8_24# OR2X1_LOC_66/A 0.02fF
C29146 AND2X1_LOC_611/a_36_24# OR2X1_LOC_415/Y 0.01fF
C29147 AND2X1_LOC_474/A AND2X1_LOC_858/B 0.05fF
C29148 OR2X1_LOC_151/A OR2X1_LOC_185/A 0.10fF
C29149 OR2X1_LOC_346/A OR2X1_LOC_161/A 0.02fF
C29150 OR2X1_LOC_776/Y OR2X1_LOC_785/B 0.16fF
C29151 AND2X1_LOC_216/A AND2X1_LOC_647/Y 0.71fF
C29152 AND2X1_LOC_63/a_36_24# OR2X1_LOC_161/B 0.00fF
C29153 AND2X1_LOC_729/Y OR2X1_LOC_329/a_8_216# 0.04fF
C29154 OR2X1_LOC_335/A OR2X1_LOC_605/B 0.11fF
C29155 OR2X1_LOC_516/B OR2X1_LOC_744/A 0.02fF
C29156 OR2X1_LOC_687/Y OR2X1_LOC_185/a_8_216# 0.03fF
C29157 AND2X1_LOC_388/Y AND2X1_LOC_436/B 0.00fF
C29158 OR2X1_LOC_482/Y AND2X1_LOC_624/A 0.15fF
C29159 AND2X1_LOC_168/Y OR2X1_LOC_600/A 0.50fF
C29160 OR2X1_LOC_804/A AND2X1_LOC_31/Y 0.07fF
C29161 VDD AND2X1_LOC_314/a_8_24# -0.00fF
C29162 OR2X1_LOC_524/Y OR2X1_LOC_441/a_36_216# 0.14fF
C29163 OR2X1_LOC_91/Y AND2X1_LOC_180/a_8_24# 0.02fF
C29164 OR2X1_LOC_144/Y AND2X1_LOC_663/A 0.05fF
C29165 AND2X1_LOC_31/Y AND2X1_LOC_428/a_8_24# 0.01fF
C29166 OR2X1_LOC_160/A OR2X1_LOC_631/A 0.11fF
C29167 OR2X1_LOC_585/A AND2X1_LOC_219/A 0.07fF
C29168 OR2X1_LOC_188/Y AND2X1_LOC_42/B 0.33fF
C29169 VDD OR2X1_LOC_250/Y 0.03fF
C29170 AND2X1_LOC_658/A OR2X1_LOC_628/a_36_216# 0.02fF
C29171 OR2X1_LOC_709/A OR2X1_LOC_269/B 0.10fF
C29172 OR2X1_LOC_455/A AND2X1_LOC_7/B 0.01fF
C29173 OR2X1_LOC_67/a_8_216# AND2X1_LOC_243/Y 0.06fF
C29174 AND2X1_LOC_651/a_8_24# OR2X1_LOC_762/Y 0.24fF
C29175 AND2X1_LOC_564/A AND2X1_LOC_149/a_8_24# 0.07fF
C29176 AND2X1_LOC_190/a_8_24# OR2X1_LOC_18/Y 0.17fF
C29177 OR2X1_LOC_604/A OR2X1_LOC_314/Y 0.38fF
C29178 VDD OR2X1_LOC_243/A 0.12fF
C29179 AND2X1_LOC_806/a_8_24# OR2X1_LOC_39/A 0.02fF
C29180 AND2X1_LOC_31/Y OR2X1_LOC_723/A 0.01fF
C29181 AND2X1_LOC_700/a_8_24# AND2X1_LOC_59/Y 0.01fF
C29182 AND2X1_LOC_70/Y OR2X1_LOC_739/A 0.03fF
C29183 OR2X1_LOC_45/B AND2X1_LOC_578/A 0.10fF
C29184 OR2X1_LOC_154/A OR2X1_LOC_114/B 0.05fF
C29185 VDD OR2X1_LOC_668/Y 0.16fF
C29186 OR2X1_LOC_814/A OR2X1_LOC_605/Y 0.01fF
C29187 OR2X1_LOC_636/B AND2X1_LOC_44/Y 0.19fF
C29188 OR2X1_LOC_538/A OR2X1_LOC_620/Y 0.27fF
C29189 AND2X1_LOC_531/a_8_24# AND2X1_LOC_40/Y 0.04fF
C29190 OR2X1_LOC_861/a_8_216# OR2X1_LOC_756/B 0.01fF
C29191 OR2X1_LOC_791/B OR2X1_LOC_792/B 0.06fF
C29192 OR2X1_LOC_51/Y OR2X1_LOC_237/Y 0.15fF
C29193 OR2X1_LOC_810/a_8_216# OR2X1_LOC_391/A 0.11fF
C29194 AND2X1_LOC_382/a_8_24# VDD -0.00fF
C29195 AND2X1_LOC_553/a_8_24# OR2X1_LOC_26/Y 0.01fF
C29196 OR2X1_LOC_132/Y OR2X1_LOC_65/B 0.00fF
C29197 VDD OR2X1_LOC_36/Y 1.17fF
C29198 OR2X1_LOC_696/A OR2X1_LOC_226/a_36_216# -0.00fF
C29199 OR2X1_LOC_160/A OR2X1_LOC_632/Y 0.16fF
C29200 OR2X1_LOC_748/A AND2X1_LOC_709/a_8_24# 0.07fF
C29201 AND2X1_LOC_92/Y OR2X1_LOC_350/a_8_216# 0.08fF
C29202 AND2X1_LOC_474/A AND2X1_LOC_573/A 0.16fF
C29203 OR2X1_LOC_589/A OR2X1_LOC_743/A 0.12fF
C29204 AND2X1_LOC_95/Y OR2X1_LOC_435/B 0.00fF
C29205 OR2X1_LOC_154/A AND2X1_LOC_172/a_36_24# 0.00fF
C29206 AND2X1_LOC_554/Y AND2X1_LOC_367/A 0.10fF
C29207 OR2X1_LOC_789/A AND2X1_LOC_751/a_36_24# 0.00fF
C29208 OR2X1_LOC_426/B OR2X1_LOC_43/A 0.28fF
C29209 OR2X1_LOC_529/Y AND2X1_LOC_500/B 0.02fF
C29210 AND2X1_LOC_605/Y AND2X1_LOC_454/Y 0.01fF
C29211 OR2X1_LOC_507/a_8_216# OR2X1_LOC_507/B 0.01fF
C29212 OR2X1_LOC_758/Y OR2X1_LOC_269/B 0.10fF
C29213 AND2X1_LOC_391/Y OR2X1_LOC_85/A 0.13fF
C29214 OR2X1_LOC_364/A AND2X1_LOC_164/a_8_24# 0.01fF
C29215 AND2X1_LOC_560/B OR2X1_LOC_56/A 0.02fF
C29216 AND2X1_LOC_70/Y OR2X1_LOC_269/B 6.86fF
C29217 AND2X1_LOC_727/A OR2X1_LOC_428/A 0.06fF
C29218 OR2X1_LOC_151/A OR2X1_LOC_435/Y 0.05fF
C29219 OR2X1_LOC_154/A OR2X1_LOC_538/A 0.03fF
C29220 OR2X1_LOC_91/A OR2X1_LOC_85/A 0.07fF
C29221 OR2X1_LOC_6/B OR2X1_LOC_3/Y 1.16fF
C29222 AND2X1_LOC_713/Y OR2X1_LOC_3/Y 0.00fF
C29223 INPUT_0 AND2X1_LOC_56/B 13.29fF
C29224 AND2X1_LOC_2/Y AND2X1_LOC_17/Y 0.33fF
C29225 OR2X1_LOC_128/a_8_216# OR2X1_LOC_736/A 0.01fF
C29226 OR2X1_LOC_690/A OR2X1_LOC_56/A 0.03fF
C29227 AND2X1_LOC_374/a_36_24# OR2X1_LOC_427/A 0.00fF
C29228 OR2X1_LOC_690/Y OR2X1_LOC_585/A 0.35fF
C29229 OR2X1_LOC_654/A OR2X1_LOC_66/A 0.14fF
C29230 AND2X1_LOC_95/Y OR2X1_LOC_61/Y 0.00fF
C29231 AND2X1_LOC_92/a_8_24# INPUT_1 0.02fF
C29232 AND2X1_LOC_638/Y OR2X1_LOC_11/Y 0.33fF
C29233 OR2X1_LOC_848/A OR2X1_LOC_391/A 0.19fF
C29234 OR2X1_LOC_318/Y OR2X1_LOC_799/A 0.03fF
C29235 AND2X1_LOC_634/Y AND2X1_LOC_219/A 0.00fF
C29236 OR2X1_LOC_519/Y AND2X1_LOC_364/A 0.80fF
C29237 OR2X1_LOC_517/Y OR2X1_LOC_275/Y 0.02fF
C29238 OR2X1_LOC_634/A OR2X1_LOC_97/B 0.06fF
C29239 INPUT_0 AND2X1_LOC_8/Y 0.08fF
C29240 OR2X1_LOC_599/A AND2X1_LOC_605/Y 0.02fF
C29241 AND2X1_LOC_661/a_8_24# OR2X1_LOC_619/Y 0.05fF
C29242 OR2X1_LOC_859/B OR2X1_LOC_391/A 0.02fF
C29243 OR2X1_LOC_429/a_8_216# INPUT_7 0.03fF
C29244 OR2X1_LOC_516/B AND2X1_LOC_840/B 0.03fF
C29245 AND2X1_LOC_3/Y AND2X1_LOC_92/Y 0.07fF
C29246 AND2X1_LOC_372/a_8_24# OR2X1_LOC_778/Y 0.03fF
C29247 AND2X1_LOC_12/Y OR2X1_LOC_620/Y 0.14fF
C29248 OR2X1_LOC_833/B OR2X1_LOC_269/a_8_216# 0.01fF
C29249 OR2X1_LOC_624/B AND2X1_LOC_616/a_8_24# 0.01fF
C29250 OR2X1_LOC_703/A OR2X1_LOC_269/B 0.03fF
C29251 AND2X1_LOC_350/a_36_24# OR2X1_LOC_46/A 0.00fF
C29252 OR2X1_LOC_589/A OR2X1_LOC_246/A 0.27fF
C29253 OR2X1_LOC_689/A OR2X1_LOC_36/Y 0.03fF
C29254 AND2X1_LOC_729/a_8_24# AND2X1_LOC_687/Y 0.09fF
C29255 OR2X1_LOC_790/A AND2X1_LOC_48/A 0.00fF
C29256 OR2X1_LOC_442/a_8_216# AND2X1_LOC_212/Y 0.05fF
C29257 OR2X1_LOC_9/Y OR2X1_LOC_46/A 0.39fF
C29258 OR2X1_LOC_95/Y OR2X1_LOC_428/A 0.11fF
C29259 OR2X1_LOC_329/B AND2X1_LOC_276/Y 0.05fF
C29260 OR2X1_LOC_502/A OR2X1_LOC_83/A 0.02fF
C29261 AND2X1_LOC_100/a_8_24# OR2X1_LOC_92/Y 0.03fF
C29262 AND2X1_LOC_12/Y AND2X1_LOC_157/a_8_24# 0.00fF
C29263 AND2X1_LOC_718/a_8_24# OR2X1_LOC_89/A 0.01fF
C29264 OR2X1_LOC_532/B OR2X1_LOC_356/A 0.01fF
C29265 OR2X1_LOC_358/a_8_216# OR2X1_LOC_405/A 0.01fF
C29266 VDD AND2X1_LOC_816/a_8_24# 0.00fF
C29267 OR2X1_LOC_6/B AND2X1_LOC_133/a_8_24# 0.01fF
C29268 OR2X1_LOC_32/B OR2X1_LOC_39/A 0.09fF
C29269 OR2X1_LOC_95/Y OR2X1_LOC_595/A 0.07fF
C29270 AND2X1_LOC_738/B OR2X1_LOC_64/Y 0.12fF
C29271 OR2X1_LOC_479/Y OR2X1_LOC_804/a_8_216# 0.02fF
C29272 OR2X1_LOC_705/B OR2X1_LOC_731/A 0.14fF
C29273 INPUT_5 D_INPUT_7 0.40fF
C29274 AND2X1_LOC_123/a_8_24# OR2X1_LOC_92/Y 0.03fF
C29275 OR2X1_LOC_64/Y OR2X1_LOC_56/A 0.34fF
C29276 AND2X1_LOC_155/a_8_24# OR2X1_LOC_52/B 0.06fF
C29277 AND2X1_LOC_317/a_8_24# AND2X1_LOC_452/Y 0.02fF
C29278 OR2X1_LOC_40/Y AND2X1_LOC_326/a_36_24# 0.00fF
C29279 AND2X1_LOC_66/a_8_24# AND2X1_LOC_243/Y 0.01fF
C29280 OR2X1_LOC_600/A AND2X1_LOC_128/a_8_24# 0.03fF
C29281 OR2X1_LOC_635/A AND2X1_LOC_683/a_8_24# 0.02fF
C29282 OR2X1_LOC_506/Y OR2X1_LOC_506/B 0.26fF
C29283 AND2X1_LOC_12/Y OR2X1_LOC_154/A 0.62fF
C29284 OR2X1_LOC_467/a_8_216# OR2X1_LOC_470/A -0.00fF
C29285 OR2X1_LOC_85/A AND2X1_LOC_573/A 0.03fF
C29286 AND2X1_LOC_741/Y AND2X1_LOC_480/a_8_24# 0.21fF
C29287 VDD OR2X1_LOC_859/A 0.08fF
C29288 OR2X1_LOC_87/A OR2X1_LOC_803/B 0.07fF
C29289 OR2X1_LOC_348/Y OR2X1_LOC_287/a_8_216# 0.02fF
C29290 OR2X1_LOC_589/A OR2X1_LOC_409/B 0.16fF
C29291 OR2X1_LOC_507/B OR2X1_LOC_643/A 0.03fF
C29292 OR2X1_LOC_315/Y OR2X1_LOC_36/Y 0.30fF
C29293 OR2X1_LOC_641/Y AND2X1_LOC_519/a_8_24# 0.04fF
C29294 AND2X1_LOC_737/Y OR2X1_LOC_74/A 0.06fF
C29295 AND2X1_LOC_32/a_8_24# AND2X1_LOC_291/a_8_24# 0.23fF
C29296 OR2X1_LOC_251/Y OR2X1_LOC_250/Y 1.40fF
C29297 OR2X1_LOC_469/a_8_216# OR2X1_LOC_738/A 0.02fF
C29298 AND2X1_LOC_784/Y AND2X1_LOC_810/Y 0.01fF
C29299 OR2X1_LOC_40/Y AND2X1_LOC_170/B 0.03fF
C29300 AND2X1_LOC_805/a_8_24# GATE_579 0.01fF
C29301 OR2X1_LOC_791/B OR2X1_LOC_269/B 0.02fF
C29302 AND2X1_LOC_318/Y AND2X1_LOC_476/Y 0.06fF
C29303 AND2X1_LOC_107/a_8_24# OR2X1_LOC_78/A 0.07fF
C29304 OR2X1_LOC_858/A OR2X1_LOC_62/B 0.03fF
C29305 OR2X1_LOC_165/a_8_216# OR2X1_LOC_74/A 0.02fF
C29306 OR2X1_LOC_308/Y AND2X1_LOC_419/a_8_24# 0.03fF
C29307 OR2X1_LOC_3/Y OR2X1_LOC_625/a_8_216# 0.14fF
C29308 OR2X1_LOC_352/a_36_216# OR2X1_LOC_365/B 0.00fF
C29309 OR2X1_LOC_64/Y AND2X1_LOC_638/Y 0.01fF
C29310 OR2X1_LOC_475/Y OR2X1_LOC_734/a_8_216# 0.41fF
C29311 AND2X1_LOC_471/a_36_24# OR2X1_LOC_56/A 0.00fF
C29312 OR2X1_LOC_754/A OR2X1_LOC_427/A 0.08fF
C29313 AND2X1_LOC_367/A OR2X1_LOC_22/Y 0.10fF
C29314 OR2X1_LOC_193/Y OR2X1_LOC_200/a_8_216# 0.00fF
C29315 AND2X1_LOC_359/B OR2X1_LOC_248/a_8_216# 0.06fF
C29316 AND2X1_LOC_349/a_8_24# OR2X1_LOC_248/Y 0.01fF
C29317 OR2X1_LOC_557/A OR2X1_LOC_402/Y 0.06fF
C29318 OR2X1_LOC_417/A OR2X1_LOC_56/A 0.28fF
C29319 AND2X1_LOC_554/Y OR2X1_LOC_490/Y 0.03fF
C29320 OR2X1_LOC_329/Y OR2X1_LOC_47/Y 0.01fF
C29321 OR2X1_LOC_36/Y OR2X1_LOC_491/Y 0.01fF
C29322 AND2X1_LOC_14/a_36_24# D_INPUT_0 0.00fF
C29323 OR2X1_LOC_339/A OR2X1_LOC_174/Y 0.07fF
C29324 AND2X1_LOC_59/Y OR2X1_LOC_333/B 0.03fF
C29325 OR2X1_LOC_371/Y OR2X1_LOC_39/A 0.10fF
C29326 OR2X1_LOC_251/Y OR2X1_LOC_36/Y 0.03fF
C29327 AND2X1_LOC_319/A OR2X1_LOC_7/A 0.07fF
C29328 OR2X1_LOC_189/Y AND2X1_LOC_580/A 0.00fF
C29329 OR2X1_LOC_329/B AND2X1_LOC_831/Y 0.07fF
C29330 OR2X1_LOC_31/Y OR2X1_LOC_25/Y 0.26fF
C29331 OR2X1_LOC_92/Y OR2X1_LOC_268/a_8_216# 0.28fF
C29332 OR2X1_LOC_506/A AND2X1_LOC_67/Y 0.04fF
C29333 OR2X1_LOC_3/Y AND2X1_LOC_139/B 0.03fF
C29334 OR2X1_LOC_45/B OR2X1_LOC_88/a_8_216# 0.01fF
C29335 AND2X1_LOC_361/A AND2X1_LOC_267/a_36_24# 0.00fF
C29336 AND2X1_LOC_12/Y OR2X1_LOC_778/A 0.01fF
C29337 OR2X1_LOC_154/A AND2X1_LOC_79/Y 0.03fF
C29338 AND2X1_LOC_794/B OR2X1_LOC_419/Y 0.10fF
C29339 OR2X1_LOC_786/Y OR2X1_LOC_776/Y 0.03fF
C29340 OR2X1_LOC_64/Y AND2X1_LOC_850/Y 0.08fF
C29341 AND2X1_LOC_17/Y OR2X1_LOC_269/B 0.02fF
C29342 AND2X1_LOC_359/B AND2X1_LOC_294/a_8_24# 0.01fF
C29343 AND2X1_LOC_555/Y OR2X1_LOC_384/Y 0.01fF
C29344 OR2X1_LOC_528/Y AND2X1_LOC_792/Y 0.07fF
C29345 OR2X1_LOC_40/Y AND2X1_LOC_721/A 0.01fF
C29346 OR2X1_LOC_495/a_36_216# OR2X1_LOC_238/Y 0.00fF
C29347 AND2X1_LOC_51/Y OR2X1_LOC_161/A 0.68fF
C29348 OR2X1_LOC_154/A AND2X1_LOC_496/a_8_24# 0.34fF
C29349 OR2X1_LOC_26/Y OR2X1_LOC_89/A 1.42fF
C29350 OR2X1_LOC_854/a_8_216# D_INPUT_0 0.03fF
C29351 OR2X1_LOC_651/a_8_216# OR2X1_LOC_654/A 0.00fF
C29352 OR2X1_LOC_43/A OR2X1_LOC_743/A 0.10fF
C29353 AND2X1_LOC_72/B AND2X1_LOC_18/Y 0.02fF
C29354 AND2X1_LOC_625/a_8_24# OR2X1_LOC_598/A -0.00fF
C29355 AND2X1_LOC_733/Y AND2X1_LOC_440/a_36_24# 0.00fF
C29356 OR2X1_LOC_121/Y OR2X1_LOC_560/A 0.00fF
C29357 AND2X1_LOC_7/B OR2X1_LOC_446/B 0.09fF
C29358 OR2X1_LOC_833/Y OR2X1_LOC_68/B 0.00fF
C29359 VDD OR2X1_LOC_419/Y 2.74fF
C29360 OR2X1_LOC_185/Y OR2X1_LOC_473/Y 0.03fF
C29361 AND2X1_LOC_25/Y AND2X1_LOC_51/Y 0.09fF
C29362 AND2X1_LOC_90/a_8_24# OR2X1_LOC_80/A 0.06fF
C29363 OR2X1_LOC_628/Y AND2X1_LOC_624/A 0.07fF
C29364 AND2X1_LOC_654/B OR2X1_LOC_409/B 0.02fF
C29365 AND2X1_LOC_512/a_8_24# AND2X1_LOC_390/B 0.01fF
C29366 OR2X1_LOC_6/B AND2X1_LOC_609/a_8_24# 0.07fF
C29367 OR2X1_LOC_185/A INPUT_1 0.39fF
C29368 OR2X1_LOC_290/Y AND2X1_LOC_476/A 0.06fF
C29369 OR2X1_LOC_479/Y OR2X1_LOC_574/A 0.03fF
C29370 OR2X1_LOC_40/Y OR2X1_LOC_331/Y 0.01fF
C29371 AND2X1_LOC_486/Y OR2X1_LOC_503/Y 0.19fF
C29372 OR2X1_LOC_22/Y AND2X1_LOC_35/Y 0.33fF
C29373 OR2X1_LOC_471/Y OR2X1_LOC_209/a_8_216# 0.04fF
C29374 OR2X1_LOC_52/a_8_216# OR2X1_LOC_7/A 0.02fF
C29375 OR2X1_LOC_756/B OR2X1_LOC_364/a_36_216# 0.00fF
C29376 AND2X1_LOC_79/Y OR2X1_LOC_204/a_36_216# 0.02fF
C29377 OR2X1_LOC_96/B OR2X1_LOC_46/A 0.01fF
C29378 OR2X1_LOC_160/B OR2X1_LOC_512/Y 0.04fF
C29379 OR2X1_LOC_180/a_36_216# OR2X1_LOC_578/B 0.00fF
C29380 INPUT_4 OR2X1_LOC_429/a_8_216# 0.00fF
C29381 OR2X1_LOC_291/Y AND2X1_LOC_610/a_8_24# 0.02fF
C29382 OR2X1_LOC_532/B AND2X1_LOC_43/B 0.05fF
C29383 OR2X1_LOC_246/a_8_216# OR2X1_LOC_54/Y 0.00fF
C29384 OR2X1_LOC_329/B AND2X1_LOC_405/a_8_24# 0.03fF
C29385 OR2X1_LOC_604/A AND2X1_LOC_657/A 0.10fF
C29386 VDD OR2X1_LOC_568/a_8_216# 0.00fF
C29387 OR2X1_LOC_22/A AND2X1_LOC_463/a_8_24# 0.01fF
C29388 AND2X1_LOC_68/a_36_24# OR2X1_LOC_69/A 0.00fF
C29389 OR2X1_LOC_416/Y AND2X1_LOC_634/a_8_24# 0.01fF
C29390 AND2X1_LOC_535/a_8_24# OR2X1_LOC_331/Y 0.04fF
C29391 AND2X1_LOC_852/Y OR2X1_LOC_46/A 0.17fF
C29392 OR2X1_LOC_161/B OR2X1_LOC_788/B 0.01fF
C29393 VDD OR2X1_LOC_344/a_8_216# 0.00fF
C29394 AND2X1_LOC_525/a_8_24# AND2X1_LOC_51/Y 0.03fF
C29395 AND2X1_LOC_708/a_8_24# OR2X1_LOC_7/A 0.09fF
C29396 OR2X1_LOC_389/B AND2X1_LOC_48/A 0.03fF
C29397 VDD OR2X1_LOC_152/A 0.21fF
C29398 VDD OR2X1_LOC_526/a_8_216# 0.00fF
C29399 OR2X1_LOC_589/A OR2X1_LOC_599/a_8_216# 0.02fF
C29400 OR2X1_LOC_502/A OR2X1_LOC_215/a_8_216# 0.05fF
C29401 OR2X1_LOC_83/Y OR2X1_LOC_46/A 0.01fF
C29402 OR2X1_LOC_743/A AND2X1_LOC_685/a_8_24# 0.19fF
C29403 AND2X1_LOC_785/A AND2X1_LOC_564/B 0.01fF
C29404 AND2X1_LOC_456/Y OR2X1_LOC_22/Y 0.02fF
C29405 OR2X1_LOC_580/A OR2X1_LOC_349/A 0.03fF
C29406 AND2X1_LOC_729/Y OR2X1_LOC_760/a_36_216# 0.00fF
C29407 AND2X1_LOC_339/a_8_24# INPUT_1 0.01fF
C29408 OR2X1_LOC_22/Y OR2X1_LOC_74/A 0.16fF
C29409 OR2X1_LOC_76/B OR2X1_LOC_241/B 0.06fF
C29410 OR2X1_LOC_651/A OR2X1_LOC_87/A 0.01fF
C29411 OR2X1_LOC_273/Y OR2X1_LOC_416/Y 0.04fF
C29412 AND2X1_LOC_65/a_8_24# AND2X1_LOC_31/Y 0.01fF
C29413 OR2X1_LOC_676/Y OR2X1_LOC_515/a_8_216# 0.02fF
C29414 OR2X1_LOC_859/a_8_216# OR2X1_LOC_561/B 0.01fF
C29415 AND2X1_LOC_42/B D_INPUT_0 0.20fF
C29416 AND2X1_LOC_170/B OR2X1_LOC_7/A 3.13fF
C29417 OR2X1_LOC_599/Y AND2X1_LOC_655/A 0.04fF
C29418 AND2X1_LOC_656/Y AND2X1_LOC_116/Y 0.00fF
C29419 OR2X1_LOC_500/A AND2X1_LOC_72/B 0.02fF
C29420 OR2X1_LOC_844/Y OR2X1_LOC_849/a_36_216# 0.02fF
C29421 OR2X1_LOC_169/B OR2X1_LOC_365/B 0.01fF
C29422 OR2X1_LOC_231/A AND2X1_LOC_31/Y 0.01fF
C29423 OR2X1_LOC_36/Y AND2X1_LOC_624/B 0.00fF
C29424 AND2X1_LOC_18/Y AND2X1_LOC_36/Y 2.38fF
C29425 OR2X1_LOC_185/Y OR2X1_LOC_241/B 0.22fF
C29426 OR2X1_LOC_36/Y OR2X1_LOC_67/Y 0.07fF
C29427 INPUT_1 AND2X1_LOC_119/a_8_24# 0.10fF
C29428 OR2X1_LOC_178/a_8_216# OR2X1_LOC_183/Y 0.01fF
C29429 OR2X1_LOC_76/a_36_216# OR2X1_LOC_553/A 0.00fF
C29430 D_INPUT_7 OR2X1_LOC_17/a_8_216# 0.14fF
C29431 OR2X1_LOC_319/B OR2X1_LOC_446/B 0.15fF
C29432 OR2X1_LOC_810/A OR2X1_LOC_795/a_8_216# 0.02fF
C29433 OR2X1_LOC_39/A AND2X1_LOC_222/Y 0.05fF
C29434 AND2X1_LOC_1/Y OR2X1_LOC_639/a_8_216# 0.01fF
C29435 AND2X1_LOC_240/Y D_INPUT_1 0.66fF
C29436 OR2X1_LOC_545/B OR2X1_LOC_443/Y 0.03fF
C29437 OR2X1_LOC_26/Y AND2X1_LOC_804/a_8_24# 0.07fF
C29438 AND2X1_LOC_22/Y OR2X1_LOC_161/B 0.05fF
C29439 VDD OR2X1_LOC_508/Y 0.19fF
C29440 AND2X1_LOC_522/a_8_24# AND2X1_LOC_44/Y 0.01fF
C29441 OR2X1_LOC_447/A OR2X1_LOC_724/A 0.01fF
C29442 OR2X1_LOC_335/B OR2X1_LOC_814/A 0.00fF
C29443 AND2X1_LOC_721/A OR2X1_LOC_7/A 0.03fF
C29444 AND2X1_LOC_31/Y OR2X1_LOC_340/Y 0.02fF
C29445 OR2X1_LOC_26/Y AND2X1_LOC_202/a_8_24# 0.01fF
C29446 OR2X1_LOC_74/A AND2X1_LOC_808/A 0.03fF
C29447 AND2X1_LOC_212/Y AND2X1_LOC_794/a_8_24# 0.02fF
C29448 OR2X1_LOC_18/Y AND2X1_LOC_216/a_36_24# 0.01fF
C29449 OR2X1_LOC_696/A AND2X1_LOC_98/a_8_24# 0.01fF
C29450 OR2X1_LOC_318/Y OR2X1_LOC_446/B 0.03fF
C29451 OR2X1_LOC_756/B OR2X1_LOC_181/Y 0.02fF
C29452 OR2X1_LOC_39/A OR2X1_LOC_68/B 0.03fF
C29453 OR2X1_LOC_130/A AND2X1_LOC_31/Y 0.06fF
C29454 OR2X1_LOC_416/Y OR2X1_LOC_75/Y 0.23fF
C29455 OR2X1_LOC_779/a_8_216# OR2X1_LOC_779/B 0.08fF
C29456 OR2X1_LOC_44/Y AND2X1_LOC_779/Y 0.01fF
C29457 AND2X1_LOC_7/B OR2X1_LOC_719/B 0.02fF
C29458 OR2X1_LOC_235/B OR2X1_LOC_523/a_36_216# 0.00fF
C29459 OR2X1_LOC_446/Y OR2X1_LOC_707/B 0.20fF
C29460 OR2X1_LOC_733/A OR2X1_LOC_722/B 0.00fF
C29461 OR2X1_LOC_856/B OR2X1_LOC_112/A 0.04fF
C29462 AND2X1_LOC_40/Y OR2X1_LOC_174/Y 0.03fF
C29463 OR2X1_LOC_186/Y AND2X1_LOC_594/a_8_24# 0.11fF
C29464 OR2X1_LOC_3/Y OR2X1_LOC_598/A 0.02fF
C29465 OR2X1_LOC_467/B OR2X1_LOC_161/B 0.04fF
C29466 OR2X1_LOC_158/A AND2X1_LOC_786/Y 0.09fF
C29467 AND2X1_LOC_53/Y AND2X1_LOC_47/Y 0.07fF
C29468 OR2X1_LOC_528/Y OR2X1_LOC_816/A 0.13fF
C29469 OR2X1_LOC_207/B OR2X1_LOC_790/A 0.15fF
C29470 AND2X1_LOC_550/a_8_24# AND2X1_LOC_564/A 0.07fF
C29471 AND2X1_LOC_3/Y OR2X1_LOC_736/a_8_216# 0.01fF
C29472 OR2X1_LOC_840/A OR2X1_LOC_308/Y 1.77fF
C29473 AND2X1_LOC_738/B AND2X1_LOC_544/Y 0.07fF
C29474 OR2X1_LOC_7/A OR2X1_LOC_331/Y 0.03fF
C29475 AND2X1_LOC_64/Y OR2X1_LOC_78/A 1.25fF
C29476 OR2X1_LOC_45/B OR2X1_LOC_681/a_8_216# 0.03fF
C29477 AND2X1_LOC_555/Y AND2X1_LOC_391/Y 0.01fF
C29478 OR2X1_LOC_855/a_8_216# OR2X1_LOC_598/Y 0.01fF
C29479 AND2X1_LOC_564/B AND2X1_LOC_658/A 0.07fF
C29480 OR2X1_LOC_542/B AND2X1_LOC_7/B 0.03fF
C29481 OR2X1_LOC_427/A OR2X1_LOC_142/Y 2.39fF
C29482 OR2X1_LOC_421/A AND2X1_LOC_639/B 0.04fF
C29483 AND2X1_LOC_555/Y OR2X1_LOC_91/A 0.03fF
C29484 AND2X1_LOC_541/a_8_24# OR2X1_LOC_56/A 0.17fF
C29485 AND2X1_LOC_84/Y OR2X1_LOC_59/Y 0.02fF
C29486 AND2X1_LOC_724/a_36_24# AND2X1_LOC_447/Y 0.01fF
C29487 AND2X1_LOC_562/a_36_24# AND2X1_LOC_285/Y 0.00fF
C29488 OR2X1_LOC_574/A OR2X1_LOC_68/B 0.03fF
C29489 AND2X1_LOC_229/a_8_24# VDD -0.00fF
C29490 OR2X1_LOC_46/A AND2X1_LOC_647/B 0.04fF
C29491 OR2X1_LOC_600/A OR2X1_LOC_373/Y 0.03fF
C29492 OR2X1_LOC_673/A AND2X1_LOC_47/Y 0.04fF
C29493 OR2X1_LOC_715/B OR2X1_LOC_596/A 0.00fF
C29494 OR2X1_LOC_223/A AND2X1_LOC_47/Y 0.05fF
C29495 OR2X1_LOC_139/A OR2X1_LOC_78/B 0.03fF
C29496 AND2X1_LOC_48/A OR2X1_LOC_339/Y 0.03fF
C29497 AND2X1_LOC_794/B OR2X1_LOC_604/A 1.32fF
C29498 AND2X1_LOC_57/Y OR2X1_LOC_856/B 0.04fF
C29499 OR2X1_LOC_177/Y VDD 0.41fF
C29500 OR2X1_LOC_244/A OR2X1_LOC_84/a_36_216# 0.00fF
C29501 OR2X1_LOC_814/A OR2X1_LOC_366/a_8_216# 0.01fF
C29502 OR2X1_LOC_6/B AND2X1_LOC_275/a_36_24# 0.01fF
C29503 OR2X1_LOC_9/Y INPUT_2 0.02fF
C29504 OR2X1_LOC_253/Y AND2X1_LOC_254/a_8_24# 0.01fF
C29505 OR2X1_LOC_620/Y OR2X1_LOC_356/B 0.02fF
C29506 OR2X1_LOC_22/Y AND2X1_LOC_647/Y 0.03fF
C29507 AND2X1_LOC_543/Y AND2X1_LOC_374/a_8_24# 0.05fF
C29508 AND2X1_LOC_22/Y OR2X1_LOC_435/B 0.21fF
C29509 AND2X1_LOC_82/Y OR2X1_LOC_78/A 0.65fF
C29510 AND2X1_LOC_22/Y AND2X1_LOC_48/a_8_24# 0.02fF
C29511 OR2X1_LOC_187/Y AND2X1_LOC_866/B 0.01fF
C29512 OR2X1_LOC_6/B OR2X1_LOC_671/a_8_216# 0.01fF
C29513 OR2X1_LOC_160/B OR2X1_LOC_641/A 6.23fF
C29514 OR2X1_LOC_244/B OR2X1_LOC_161/B 0.18fF
C29515 AND2X1_LOC_244/a_8_24# AND2X1_LOC_860/A 0.00fF
C29516 OR2X1_LOC_158/A AND2X1_LOC_218/Y 0.02fF
C29517 OR2X1_LOC_604/A VDD 6.36fF
C29518 VDD OR2X1_LOC_745/a_8_216# 0.00fF
C29519 OR2X1_LOC_337/A OR2X1_LOC_703/A 0.01fF
C29520 OR2X1_LOC_524/Y AND2X1_LOC_469/a_8_24# 0.25fF
C29521 VDD AND2X1_LOC_207/B 0.01fF
C29522 OR2X1_LOC_469/a_8_216# AND2X1_LOC_36/Y 0.01fF
C29523 OR2X1_LOC_36/Y AND2X1_LOC_269/a_8_24# 0.01fF
C29524 OR2X1_LOC_19/B OR2X1_LOC_80/A 0.37fF
C29525 AND2X1_LOC_672/B OR2X1_LOC_68/B 0.03fF
C29526 OR2X1_LOC_188/Y OR2X1_LOC_76/B 0.02fF
C29527 OR2X1_LOC_712/a_8_216# AND2X1_LOC_44/Y 0.01fF
C29528 AND2X1_LOC_22/Y OR2X1_LOC_61/Y 0.02fF
C29529 VDD OR2X1_LOC_66/A 1.81fF
C29530 OR2X1_LOC_223/A OR2X1_LOC_795/a_36_216# 0.00fF
C29531 VDD OR2X1_LOC_841/A 0.23fF
C29532 OR2X1_LOC_842/A OR2X1_LOC_190/A 1.19fF
C29533 AND2X1_LOC_70/Y OR2X1_LOC_832/a_36_216# 0.00fF
C29534 OR2X1_LOC_421/A OR2X1_LOC_744/A 0.04fF
C29535 OR2X1_LOC_854/a_36_216# OR2X1_LOC_161/B 0.00fF
C29536 AND2X1_LOC_70/Y AND2X1_LOC_172/a_8_24# 0.10fF
C29537 OR2X1_LOC_49/A OR2X1_LOC_837/B 0.04fF
C29538 OR2X1_LOC_630/Y AND2X1_LOC_18/Y 0.07fF
C29539 OR2X1_LOC_810/A OR2X1_LOC_130/a_36_216# 0.17fF
C29540 OR2X1_LOC_441/Y AND2X1_LOC_477/Y 0.07fF
C29541 OR2X1_LOC_26/Y AND2X1_LOC_590/a_8_24# 0.03fF
C29542 OR2X1_LOC_510/Y OR2X1_LOC_392/B 0.01fF
C29543 OR2X1_LOC_624/A OR2X1_LOC_576/A 0.05fF
C29544 OR2X1_LOC_464/a_8_216# OR2X1_LOC_741/Y 0.01fF
C29545 OR2X1_LOC_630/a_8_216# OR2X1_LOC_161/B 0.02fF
C29546 OR2X1_LOC_805/A OR2X1_LOC_366/B 0.00fF
C29547 AND2X1_LOC_374/a_8_24# OR2X1_LOC_322/Y 0.23fF
C29548 OR2X1_LOC_666/A OR2X1_LOC_59/Y 0.07fF
C29549 AND2X1_LOC_391/Y OR2X1_LOC_51/Y 0.12fF
C29550 OR2X1_LOC_139/A OR2X1_LOC_375/A 0.12fF
C29551 OR2X1_LOC_51/Y AND2X1_LOC_858/B 0.08fF
C29552 OR2X1_LOC_51/Y OR2X1_LOC_91/A 0.08fF
C29553 OR2X1_LOC_98/A OR2X1_LOC_66/A 0.01fF
C29554 OR2X1_LOC_664/a_8_216# OR2X1_LOC_161/B 0.01fF
C29555 AND2X1_LOC_161/Y AND2X1_LOC_162/a_8_24# 0.19fF
C29556 OR2X1_LOC_6/B OR2X1_LOC_502/A 0.08fF
C29557 OR2X1_LOC_339/a_8_216# AND2X1_LOC_41/A 0.04fF
C29558 AND2X1_LOC_64/Y OR2X1_LOC_155/A 0.11fF
C29559 AND2X1_LOC_56/B AND2X1_LOC_7/B 12.81fF
C29560 AND2X1_LOC_462/B OR2X1_LOC_598/A 0.02fF
C29561 OR2X1_LOC_91/Y AND2X1_LOC_445/a_8_24# 0.02fF
C29562 OR2X1_LOC_405/A AND2X1_LOC_65/A 0.02fF
C29563 OR2X1_LOC_97/A AND2X1_LOC_32/a_8_24# 0.01fF
C29564 AND2X1_LOC_31/Y AND2X1_LOC_88/Y 0.03fF
C29565 OR2X1_LOC_689/a_8_216# AND2X1_LOC_194/Y 0.01fF
C29566 OR2X1_LOC_65/B AND2X1_LOC_249/a_36_24# 0.00fF
C29567 OR2X1_LOC_132/a_8_216# OR2X1_LOC_517/A 0.03fF
C29568 AND2X1_LOC_305/a_8_24# OR2X1_LOC_307/A 0.00fF
C29569 OR2X1_LOC_315/a_8_216# OR2X1_LOC_315/Y 0.03fF
C29570 AND2X1_LOC_8/Y AND2X1_LOC_7/B 8.23fF
C29571 AND2X1_LOC_362/a_8_24# AND2X1_LOC_474/A 0.01fF
C29572 OR2X1_LOC_186/Y OR2X1_LOC_703/B 0.23fF
C29573 OR2X1_LOC_92/Y AND2X1_LOC_447/Y 0.00fF
C29574 AND2X1_LOC_456/B OR2X1_LOC_744/A 0.03fF
C29575 AND2X1_LOC_785/a_8_24# OR2X1_LOC_371/Y 0.00fF
C29576 AND2X1_LOC_452/Y OR2X1_LOC_765/a_8_216# 0.01fF
C29577 OR2X1_LOC_186/Y OR2X1_LOC_87/A 0.07fF
C29578 AND2X1_LOC_378/a_8_24# OR2X1_LOC_459/A 0.01fF
C29579 AND2X1_LOC_377/Y AND2X1_LOC_378/a_36_24# 0.01fF
C29580 OR2X1_LOC_512/A OR2X1_LOC_78/A 0.01fF
C29581 OR2X1_LOC_696/A AND2X1_LOC_856/B 0.01fF
C29582 AND2X1_LOC_51/A AND2X1_LOC_44/Y 0.01fF
C29583 OR2X1_LOC_12/Y OR2X1_LOC_418/Y 0.01fF
C29584 OR2X1_LOC_528/Y AND2X1_LOC_807/Y 0.38fF
C29585 AND2X1_LOC_12/Y AND2X1_LOC_299/a_8_24# 0.09fF
C29586 AND2X1_LOC_713/a_8_24# OR2X1_LOC_36/Y 0.01fF
C29587 OR2X1_LOC_696/A AND2X1_LOC_464/Y 0.10fF
C29588 OR2X1_LOC_508/a_36_216# OR2X1_LOC_87/A 0.02fF
C29589 OR2X1_LOC_72/Y AND2X1_LOC_215/A 0.16fF
C29590 VDD OR2X1_LOC_252/a_8_216# 0.00fF
C29591 OR2X1_LOC_847/A AND2X1_LOC_616/a_8_24# 0.01fF
C29592 AND2X1_LOC_571/a_36_24# OR2X1_LOC_89/A 0.00fF
C29593 OR2X1_LOC_604/A OR2X1_LOC_616/Y 0.00fF
C29594 AND2X1_LOC_31/Y OR2X1_LOC_365/B 0.03fF
C29595 INPUT_5 AND2X1_LOC_50/a_8_24# 0.01fF
C29596 OR2X1_LOC_823/a_8_216# OR2X1_LOC_51/Y 0.01fF
C29597 OR2X1_LOC_232/a_8_216# OR2X1_LOC_16/A 0.02fF
C29598 AND2X1_LOC_758/a_8_24# OR2X1_LOC_616/Y 0.01fF
C29599 AND2X1_LOC_713/a_36_24# OR2X1_LOC_599/A 0.00fF
C29600 OR2X1_LOC_296/a_8_216# OR2X1_LOC_161/B 0.02fF
C29601 OR2X1_LOC_49/A OR2X1_LOC_73/a_8_216# 0.01fF
C29602 AND2X1_LOC_654/Y OR2X1_LOC_59/Y 0.07fF
C29603 AND2X1_LOC_508/B AND2X1_LOC_862/A 0.00fF
C29604 AND2X1_LOC_182/A OR2X1_LOC_44/Y 0.03fF
C29605 OR2X1_LOC_87/A OR2X1_LOC_726/A 0.03fF
C29606 AND2X1_LOC_508/B AND2X1_LOC_624/A 0.07fF
C29607 AND2X1_LOC_738/B AND2X1_LOC_550/A 0.03fF
C29608 AND2X1_LOC_552/A OR2X1_LOC_26/Y 0.03fF
C29609 OR2X1_LOC_306/Y VDD 0.01fF
C29610 OR2X1_LOC_604/A AND2X1_LOC_447/a_36_24# 0.02fF
C29611 OR2X1_LOC_517/A AND2X1_LOC_139/a_36_24# 0.01fF
C29612 OR2X1_LOC_51/Y AND2X1_LOC_573/A 0.02fF
C29613 OR2X1_LOC_810/A OR2X1_LOC_113/B 0.05fF
C29614 OR2X1_LOC_52/Y OR2X1_LOC_56/Y 0.05fF
C29615 AND2X1_LOC_483/a_8_24# OR2X1_LOC_816/A 0.01fF
C29616 OR2X1_LOC_135/a_8_216# OR2X1_LOC_3/Y 0.01fF
C29617 OR2X1_LOC_364/A OR2X1_LOC_325/B 0.19fF
C29618 AND2X1_LOC_860/A AND2X1_LOC_286/Y 0.01fF
C29619 AND2X1_LOC_675/Y OR2X1_LOC_531/a_36_216# 0.00fF
C29620 AND2X1_LOC_508/a_8_24# AND2X1_LOC_624/A 0.02fF
C29621 AND2X1_LOC_538/a_36_24# OR2X1_LOC_43/A 0.01fF
C29622 AND2X1_LOC_565/a_8_24# AND2X1_LOC_580/A 0.01fF
C29623 VDD OR2X1_LOC_80/Y 0.33fF
C29624 OR2X1_LOC_40/Y AND2X1_LOC_361/A 0.02fF
C29625 OR2X1_LOC_467/A OR2X1_LOC_453/a_8_216# 0.01fF
C29626 OR2X1_LOC_52/B AND2X1_LOC_448/a_8_24# 0.03fF
C29627 OR2X1_LOC_49/A AND2X1_LOC_260/a_8_24# 0.01fF
C29628 AND2X1_LOC_50/Y AND2X1_LOC_53/a_8_24# 0.03fF
C29629 AND2X1_LOC_501/Y AND2X1_LOC_576/Y 0.03fF
C29630 OR2X1_LOC_121/B OR2X1_LOC_352/a_36_216# 0.02fF
C29631 OR2X1_LOC_329/B AND2X1_LOC_436/B 0.02fF
C29632 OR2X1_LOC_468/A OR2X1_LOC_593/a_8_216# 0.01fF
C29633 OR2X1_LOC_630/Y OR2X1_LOC_500/A 0.92fF
C29634 OR2X1_LOC_304/Y AND2X1_LOC_774/A 0.03fF
C29635 OR2X1_LOC_326/B OR2X1_LOC_502/A 0.27fF
C29636 OR2X1_LOC_624/A AND2X1_LOC_41/A 0.05fF
C29637 OR2X1_LOC_160/B OR2X1_LOC_449/A 0.01fF
C29638 OR2X1_LOC_604/A OR2X1_LOC_251/Y 0.03fF
C29639 AND2X1_LOC_737/Y AND2X1_LOC_741/a_8_24# 0.00fF
C29640 OR2X1_LOC_702/A OR2X1_LOC_151/A 0.00fF
C29641 OR2X1_LOC_683/a_8_216# OR2X1_LOC_427/A 0.01fF
C29642 AND2X1_LOC_310/a_8_24# OR2X1_LOC_87/A 0.03fF
C29643 VDD OR2X1_LOC_651/a_8_216# 0.21fF
C29644 OR2X1_LOC_541/A AND2X1_LOC_272/a_8_24# 0.01fF
C29645 OR2X1_LOC_506/B AND2X1_LOC_239/a_36_24# 0.00fF
C29646 AND2X1_LOC_347/Y AND2X1_LOC_847/Y 0.02fF
C29647 OR2X1_LOC_637/Y OR2X1_LOC_375/A 0.03fF
C29648 AND2X1_LOC_367/A OR2X1_LOC_39/A 0.10fF
C29649 AND2X1_LOC_724/Y AND2X1_LOC_602/a_8_24# 0.00fF
C29650 OR2X1_LOC_298/a_36_216# OR2X1_LOC_619/Y 0.01fF
C29651 GATE_366 OR2X1_LOC_59/Y 0.03fF
C29652 OR2X1_LOC_109/Y OR2X1_LOC_92/Y 0.06fF
C29653 OR2X1_LOC_508/A OR2X1_LOC_624/A 0.10fF
C29654 AND2X1_LOC_334/a_8_24# OR2X1_LOC_16/A 0.01fF
C29655 AND2X1_LOC_392/A AND2X1_LOC_123/a_36_24# 0.01fF
C29656 OR2X1_LOC_51/Y OR2X1_LOC_669/Y 0.18fF
C29657 OR2X1_LOC_597/A OR2X1_LOC_485/A 0.21fF
C29658 AND2X1_LOC_598/a_36_24# OR2X1_LOC_744/A 0.01fF
C29659 OR2X1_LOC_805/A OR2X1_LOC_736/A 0.03fF
C29660 OR2X1_LOC_43/A AND2X1_LOC_691/a_36_24# 0.00fF
C29661 AND2X1_LOC_537/Y OR2X1_LOC_12/Y 0.11fF
C29662 OR2X1_LOC_92/Y AND2X1_LOC_448/Y 0.01fF
C29663 AND2X1_LOC_364/Y AND2X1_LOC_661/A 0.02fF
C29664 AND2X1_LOC_810/A OR2X1_LOC_22/Y 0.03fF
C29665 AND2X1_LOC_41/A OR2X1_LOC_264/a_36_216# 0.03fF
C29666 OR2X1_LOC_585/A OR2X1_LOC_597/a_8_216# 0.01fF
C29667 OR2X1_LOC_693/a_8_216# OR2X1_LOC_46/A 0.07fF
C29668 OR2X1_LOC_426/B OR2X1_LOC_299/Y 0.02fF
C29669 OR2X1_LOC_394/Y AND2X1_LOC_400/a_8_24# 0.01fF
C29670 OR2X1_LOC_178/Y OR2X1_LOC_485/A 0.01fF
C29671 OR2X1_LOC_601/a_36_216# OR2X1_LOC_16/A 0.03fF
C29672 OR2X1_LOC_402/B AND2X1_LOC_3/Y 0.01fF
C29673 OR2X1_LOC_319/B AND2X1_LOC_56/B 0.00fF
C29674 OR2X1_LOC_744/A AND2X1_LOC_717/B 0.25fF
C29675 AND2X1_LOC_59/Y OR2X1_LOC_620/Y 0.00fF
C29676 OR2X1_LOC_131/Y AND2X1_LOC_141/a_8_24# 0.13fF
C29677 OR2X1_LOC_91/Y AND2X1_LOC_717/Y 0.01fF
C29678 OR2X1_LOC_256/Y OR2X1_LOC_248/a_36_216# 0.00fF
C29679 OR2X1_LOC_117/Y OR2X1_LOC_517/A 0.85fF
C29680 OR2X1_LOC_427/A AND2X1_LOC_453/a_8_24# 0.01fF
C29681 AND2X1_LOC_95/Y AND2X1_LOC_132/a_8_24# 0.01fF
C29682 AND2X1_LOC_566/B OR2X1_LOC_46/A 0.03fF
C29683 OR2X1_LOC_160/A OR2X1_LOC_796/a_8_216# 0.02fF
C29684 AND2X1_LOC_367/A AND2X1_LOC_211/B 0.07fF
C29685 OR2X1_LOC_48/B AND2X1_LOC_648/a_36_24# 0.02fF
C29686 AND2X1_LOC_486/Y OR2X1_LOC_36/Y 0.03fF
C29687 AND2X1_LOC_48/A OR2X1_LOC_596/a_8_216# 0.02fF
C29688 AND2X1_LOC_605/Y OR2X1_LOC_7/A 0.02fF
C29689 OR2X1_LOC_306/Y OR2X1_LOC_829/a_8_216# 0.39fF
C29690 OR2X1_LOC_160/B OR2X1_LOC_844/Y 0.02fF
C29691 OR2X1_LOC_539/A OR2X1_LOC_269/B 0.01fF
C29692 OR2X1_LOC_290/Y OR2X1_LOC_690/A 0.23fF
C29693 OR2X1_LOC_409/B AND2X1_LOC_771/a_8_24# 0.02fF
C29694 OR2X1_LOC_161/A OR2X1_LOC_541/a_8_216# 0.14fF
C29695 OR2X1_LOC_18/Y AND2X1_LOC_648/a_36_24# 0.00fF
C29696 OR2X1_LOC_291/A OR2X1_LOC_232/Y 0.10fF
C29697 AND2X1_LOC_584/a_8_24# AND2X1_LOC_11/Y 0.17fF
C29698 OR2X1_LOC_6/A OR2X1_LOC_278/Y 0.02fF
C29699 OR2X1_LOC_680/A AND2X1_LOC_573/A 0.03fF
C29700 OR2X1_LOC_22/Y AND2X1_LOC_860/A 0.07fF
C29701 OR2X1_LOC_318/B OR2X1_LOC_605/Y 0.02fF
C29702 AND2X1_LOC_662/B OR2X1_LOC_6/A 0.03fF
C29703 OR2X1_LOC_256/Y OR2X1_LOC_485/A 0.01fF
C29704 AND2X1_LOC_50/Y OR2X1_LOC_654/A 0.01fF
C29705 AND2X1_LOC_36/Y OR2X1_LOC_789/A 0.51fF
C29706 OR2X1_LOC_296/Y OR2X1_LOC_736/A 0.04fF
C29707 OR2X1_LOC_154/A AND2X1_LOC_59/Y 0.32fF
C29708 OR2X1_LOC_244/A OR2X1_LOC_641/A 0.01fF
C29709 OR2X1_LOC_32/B OR2X1_LOC_85/A 0.05fF
C29710 OR2X1_LOC_206/A OR2X1_LOC_78/A 0.05fF
C29711 AND2X1_LOC_56/B OR2X1_LOC_407/a_8_216# 0.02fF
C29712 AND2X1_LOC_319/a_8_24# AND2X1_LOC_810/B 0.01fF
C29713 OR2X1_LOC_472/a_8_216# OR2X1_LOC_634/A 0.15fF
C29714 AND2X1_LOC_40/Y AND2X1_LOC_42/B 0.03fF
C29715 OR2X1_LOC_69/a_36_216# OR2X1_LOC_39/A 0.02fF
C29716 AND2X1_LOC_56/B OR2X1_LOC_805/A 0.03fF
C29717 OR2X1_LOC_427/A OR2X1_LOC_238/Y 0.03fF
C29718 OR2X1_LOC_654/A OR2X1_LOC_637/a_36_216# 0.02fF
C29719 OR2X1_LOC_71/Y AND2X1_LOC_489/a_8_24# 0.01fF
C29720 OR2X1_LOC_528/Y OR2X1_LOC_95/Y 0.16fF
C29721 OR2X1_LOC_348/Y OR2X1_LOC_532/B 0.20fF
C29722 OR2X1_LOC_311/Y INPUT_0 0.02fF
C29723 OR2X1_LOC_421/A OR2X1_LOC_31/Y 0.06fF
C29724 AND2X1_LOC_81/B OR2X1_LOC_87/A 0.08fF
C29725 AND2X1_LOC_747/a_8_24# OR2X1_LOC_782/B 0.01fF
C29726 AND2X1_LOC_286/Y AND2X1_LOC_287/Y 1.01fF
C29727 AND2X1_LOC_747/a_8_24# OR2X1_LOC_87/A 0.01fF
C29728 OR2X1_LOC_462/B AND2X1_LOC_89/a_8_24# 0.01fF
C29729 OR2X1_LOC_158/A AND2X1_LOC_114/Y 0.01fF
C29730 OR2X1_LOC_91/Y AND2X1_LOC_560/B 0.07fF
C29731 OR2X1_LOC_92/Y AND2X1_LOC_729/B 0.01fF
C29732 OR2X1_LOC_864/A OR2X1_LOC_130/A 0.07fF
C29733 AND2X1_LOC_538/Y INPUT_0 0.01fF
C29734 OR2X1_LOC_417/A AND2X1_LOC_285/Y 0.00fF
C29735 AND2X1_LOC_12/Y AND2X1_LOC_495/a_36_24# 0.00fF
C29736 AND2X1_LOC_580/A AND2X1_LOC_806/A 0.03fF
C29737 OR2X1_LOC_70/Y AND2X1_LOC_654/Y 0.19fF
C29738 OR2X1_LOC_787/Y OR2X1_LOC_161/A 0.05fF
C29739 AND2X1_LOC_67/Y OR2X1_LOC_737/A 0.02fF
C29740 AND2X1_LOC_569/A AND2X1_LOC_565/Y 0.06fF
C29741 AND2X1_LOC_564/A AND2X1_LOC_222/Y 0.03fF
C29742 AND2X1_LOC_472/B OR2X1_LOC_6/A 0.02fF
C29743 OR2X1_LOC_529/Y AND2X1_LOC_113/Y 0.35fF
C29744 AND2X1_LOC_576/a_8_24# OR2X1_LOC_89/A 0.02fF
C29745 AND2X1_LOC_702/Y AND2X1_LOC_715/a_8_24# 0.11fF
C29746 OR2X1_LOC_449/B OR2X1_LOC_593/a_8_216# 0.06fF
C29747 OR2X1_LOC_86/Y OR2X1_LOC_43/A 0.09fF
C29748 AND2X1_LOC_211/B AND2X1_LOC_35/Y 0.01fF
C29749 OR2X1_LOC_40/Y AND2X1_LOC_675/a_8_24# 0.01fF
C29750 AND2X1_LOC_772/B OR2X1_LOC_95/Y 0.05fF
C29751 AND2X1_LOC_716/Y AND2X1_LOC_514/Y 0.03fF
C29752 D_GATE_865 OR2X1_LOC_269/B 0.01fF
C29753 OR2X1_LOC_185/A OR2X1_LOC_476/Y 0.01fF
C29754 OR2X1_LOC_409/B OR2X1_LOC_585/Y 0.01fF
C29755 OR2X1_LOC_74/A OR2X1_LOC_39/A 0.28fF
C29756 OR2X1_LOC_696/Y OR2X1_LOC_48/B 0.02fF
C29757 AND2X1_LOC_658/B AND2X1_LOC_796/Y 0.07fF
C29758 OR2X1_LOC_306/a_36_216# AND2X1_LOC_390/B 0.01fF
C29759 AND2X1_LOC_41/A OR2X1_LOC_447/Y 0.07fF
C29760 OR2X1_LOC_269/Y AND2X1_LOC_18/Y 0.02fF
C29761 VDD OR2X1_LOC_84/A 0.36fF
C29762 OR2X1_LOC_55/a_8_216# OR2X1_LOC_56/A 0.05fF
C29763 AND2X1_LOC_577/Y AND2X1_LOC_578/A 0.04fF
C29764 AND2X1_LOC_18/Y OR2X1_LOC_340/a_8_216# 0.02fF
C29765 OR2X1_LOC_434/a_36_216# OR2X1_LOC_814/A 0.01fF
C29766 OR2X1_LOC_663/A D_INPUT_0 0.07fF
C29767 OR2X1_LOC_124/B OR2X1_LOC_786/Y -0.00fF
C29768 OR2X1_LOC_845/A OR2X1_LOC_66/A 0.03fF
C29769 OR2X1_LOC_233/a_8_216# OR2X1_LOC_85/A 0.01fF
C29770 OR2X1_LOC_188/Y OR2X1_LOC_578/B 0.03fF
C29771 AND2X1_LOC_59/Y OR2X1_LOC_778/A 0.02fF
C29772 AND2X1_LOC_514/Y AND2X1_LOC_654/Y 0.03fF
C29773 OR2X1_LOC_154/A OR2X1_LOC_688/Y 0.01fF
C29774 AND2X1_LOC_42/B OR2X1_LOC_87/Y 0.01fF
C29775 OR2X1_LOC_585/A AND2X1_LOC_637/Y 0.01fF
C29776 AND2X1_LOC_84/a_8_24# OR2X1_LOC_26/Y 0.03fF
C29777 OR2X1_LOC_8/Y AND2X1_LOC_837/a_8_24# 0.02fF
C29778 OR2X1_LOC_7/A AND2X1_LOC_361/A 0.09fF
C29779 OR2X1_LOC_40/Y AND2X1_LOC_795/Y 0.00fF
C29780 OR2X1_LOC_604/A AND2X1_LOC_624/B 0.54fF
C29781 AND2X1_LOC_351/Y OR2X1_LOC_18/Y 0.19fF
C29782 OR2X1_LOC_160/B OR2X1_LOC_796/B 0.02fF
C29783 INPUT_0 D_INPUT_3 0.07fF
C29784 AND2X1_LOC_512/Y OR2X1_LOC_95/Y 0.01fF
C29785 OR2X1_LOC_432/a_8_216# OR2X1_LOC_22/Y 0.01fF
C29786 AND2X1_LOC_40/Y OR2X1_LOC_286/B 0.03fF
C29787 AND2X1_LOC_680/a_8_24# OR2X1_LOC_739/A 0.01fF
C29788 AND2X1_LOC_711/Y GATE_366 0.13fF
C29789 AND2X1_LOC_663/B AND2X1_LOC_848/Y 0.04fF
C29790 OR2X1_LOC_679/A AND2X1_LOC_147/a_8_24# 0.21fF
C29791 OR2X1_LOC_476/B OR2X1_LOC_405/a_36_216# 0.01fF
C29792 OR2X1_LOC_831/a_8_216# AND2X1_LOC_51/Y 0.02fF
C29793 OR2X1_LOC_160/A OR2X1_LOC_520/B 0.12fF
C29794 OR2X1_LOC_12/Y AND2X1_LOC_796/A 0.10fF
C29795 OR2X1_LOC_502/A AND2X1_LOC_47/Y 0.87fF
C29796 OR2X1_LOC_91/Y OR2X1_LOC_64/Y 0.52fF
C29797 OR2X1_LOC_6/B OR2X1_LOC_398/a_8_216# 0.01fF
C29798 AND2X1_LOC_211/B OR2X1_LOC_74/A 0.51fF
C29799 OR2X1_LOC_604/A OR2X1_LOC_163/Y 0.03fF
C29800 OR2X1_LOC_70/Y OR2X1_LOC_312/Y 0.68fF
C29801 OR2X1_LOC_530/Y AND2X1_LOC_548/a_8_24# 0.23fF
C29802 OR2X1_LOC_412/a_8_216# OR2X1_LOC_316/Y 0.40fF
C29803 OR2X1_LOC_19/B OR2X1_LOC_6/A 0.17fF
C29804 OR2X1_LOC_415/A OR2X1_LOC_753/A 0.60fF
C29805 AND2X1_LOC_47/Y OR2X1_LOC_571/B 0.01fF
C29806 OR2X1_LOC_811/A OR2X1_LOC_276/B 0.07fF
C29807 OR2X1_LOC_824/Y OR2X1_LOC_54/Y 0.42fF
C29808 OR2X1_LOC_656/B OR2X1_LOC_218/Y 0.19fF
C29809 AND2X1_LOC_113/a_8_24# OR2X1_LOC_47/Y 0.02fF
C29810 OR2X1_LOC_510/Y OR2X1_LOC_532/B 0.03fF
C29811 AND2X1_LOC_128/a_36_24# OR2X1_LOC_6/A 0.00fF
C29812 OR2X1_LOC_3/Y OR2X1_LOC_481/A 0.16fF
C29813 AND2X1_LOC_519/a_8_24# OR2X1_LOC_87/B 0.02fF
C29814 AND2X1_LOC_572/A OR2X1_LOC_71/Y 0.02fF
C29815 AND2X1_LOC_848/Y AND2X1_LOC_849/a_8_24# 0.01fF
C29816 OR2X1_LOC_325/B OR2X1_LOC_578/B 0.03fF
C29817 OR2X1_LOC_502/a_8_216# OR2X1_LOC_502/Y 0.05fF
C29818 AND2X1_LOC_514/Y OR2X1_LOC_312/Y 0.07fF
C29819 AND2X1_LOC_572/Y AND2X1_LOC_866/A 0.03fF
C29820 OR2X1_LOC_185/Y D_INPUT_0 0.43fF
C29821 OR2X1_LOC_91/Y OR2X1_LOC_417/A 0.74fF
C29822 OR2X1_LOC_864/A OR2X1_LOC_62/B 0.05fF
C29823 OR2X1_LOC_400/A AND2X1_LOC_47/Y 0.01fF
C29824 AND2X1_LOC_342/Y OR2X1_LOC_95/Y 0.07fF
C29825 OR2X1_LOC_506/A OR2X1_LOC_223/A 0.02fF
C29826 OR2X1_LOC_617/Y AND2X1_LOC_663/B 0.01fF
C29827 OR2X1_LOC_70/A OR2X1_LOC_762/Y 0.01fF
C29828 AND2X1_LOC_715/A OR2X1_LOC_521/a_8_216# 0.01fF
C29829 AND2X1_LOC_486/Y OR2X1_LOC_419/Y 0.01fF
C29830 OR2X1_LOC_502/A OR2X1_LOC_598/A 0.03fF
C29831 OR2X1_LOC_527/Y OR2X1_LOC_64/Y 0.13fF
C29832 OR2X1_LOC_810/A OR2X1_LOC_532/B 0.01fF
C29833 AND2X1_LOC_502/a_8_24# OR2X1_LOC_184/Y 0.24fF
C29834 AND2X1_LOC_191/Y AND2X1_LOC_629/Y 0.09fF
C29835 OR2X1_LOC_678/Y OR2X1_LOC_779/B 0.01fF
C29836 AND2X1_LOC_41/A OR2X1_LOC_513/a_8_216# 0.01fF
C29837 OR2X1_LOC_137/Y AND2X1_LOC_47/Y 0.08fF
C29838 OR2X1_LOC_252/a_8_216# AND2X1_LOC_624/B 0.01fF
C29839 OR2X1_LOC_417/Y OR2X1_LOC_64/Y 0.03fF
C29840 AND2X1_LOC_733/a_8_24# AND2X1_LOC_222/Y 0.01fF
C29841 AND2X1_LOC_304/a_8_24# OR2X1_LOC_779/B 0.20fF
C29842 OR2X1_LOC_786/a_8_216# OR2X1_LOC_771/B 0.26fF
C29843 AND2X1_LOC_560/B D_INPUT_3 0.00fF
C29844 OR2X1_LOC_36/Y AND2X1_LOC_660/A 0.03fF
C29845 OR2X1_LOC_278/a_36_216# D_INPUT_0 0.01fF
C29846 OR2X1_LOC_3/Y OR2X1_LOC_71/Y 0.06fF
C29847 OR2X1_LOC_311/Y OR2X1_LOC_64/Y 0.02fF
C29848 OR2X1_LOC_31/Y AND2X1_LOC_717/B 0.05fF
C29849 AND2X1_LOC_658/A OR2X1_LOC_437/A 0.07fF
C29850 OR2X1_LOC_359/a_8_216# OR2X1_LOC_349/B 0.18fF
C29851 OR2X1_LOC_160/A AND2X1_LOC_497/a_8_24# 0.04fF
C29852 OR2X1_LOC_616/Y AND2X1_LOC_805/a_8_24# 0.02fF
C29853 OR2X1_LOC_864/A AND2X1_LOC_88/Y 0.03fF
C29854 OR2X1_LOC_36/Y AND2X1_LOC_646/a_8_24# 0.02fF
C29855 OR2X1_LOC_308/A AND2X1_LOC_44/Y 0.00fF
C29856 OR2X1_LOC_59/Y OR2X1_LOC_13/B 0.54fF
C29857 OR2X1_LOC_391/A OR2X1_LOC_558/A 0.03fF
C29858 OR2X1_LOC_70/Y OR2X1_LOC_75/a_8_216# 0.05fF
C29859 AND2X1_LOC_141/B OR2X1_LOC_95/Y 0.19fF
C29860 OR2X1_LOC_87/A OR2X1_LOC_66/Y 0.03fF
C29861 AND2X1_LOC_463/B AND2X1_LOC_472/B 0.00fF
C29862 OR2X1_LOC_138/a_36_216# OR2X1_LOC_691/Y 0.00fF
C29863 AND2X1_LOC_813/a_8_24# AND2X1_LOC_79/Y 0.04fF
C29864 OR2X1_LOC_40/Y OR2X1_LOC_387/A 0.83fF
C29865 OR2X1_LOC_22/Y OR2X1_LOC_263/a_8_216# 0.01fF
C29866 OR2X1_LOC_196/B OR2X1_LOC_706/B 0.11fF
C29867 OR2X1_LOC_417/Y OR2X1_LOC_417/A 0.00fF
C29868 AND2X1_LOC_721/Y AND2X1_LOC_786/Y 0.19fF
C29869 AND2X1_LOC_278/a_8_24# OR2X1_LOC_68/B 0.02fF
C29870 OR2X1_LOC_638/B D_INPUT_6 0.08fF
C29871 OR2X1_LOC_377/A OR2X1_LOC_68/B 0.35fF
C29872 OR2X1_LOC_11/Y OR2X1_LOC_11/a_8_216# -0.00fF
C29873 OR2X1_LOC_3/Y D_INPUT_1 0.03fF
C29874 VDD OR2X1_LOC_502/a_8_216# 0.21fF
C29875 AND2X1_LOC_692/a_8_24# OR2X1_LOC_706/B 0.01fF
C29876 OR2X1_LOC_76/A OR2X1_LOC_440/A 4.41fF
C29877 OR2X1_LOC_89/A AND2X1_LOC_792/Y 0.28fF
C29878 OR2X1_LOC_161/B OR2X1_LOC_162/A 0.02fF
C29879 OR2X1_LOC_64/Y D_INPUT_3 0.03fF
C29880 AND2X1_LOC_48/A AND2X1_LOC_47/Y 0.10fF
C29881 AND2X1_LOC_824/B OR2X1_LOC_68/B 2.67fF
C29882 OR2X1_LOC_95/Y OR2X1_LOC_54/Y 0.08fF
C29883 OR2X1_LOC_139/A OR2X1_LOC_549/A 0.10fF
C29884 OR2X1_LOC_158/A OR2X1_LOC_312/a_8_216# 0.05fF
C29885 OR2X1_LOC_287/B OR2X1_LOC_366/a_36_216# 0.00fF
C29886 OR2X1_LOC_175/B OR2X1_LOC_112/A 0.04fF
C29887 OR2X1_LOC_178/a_8_216# AND2X1_LOC_465/A 0.03fF
C29888 OR2X1_LOC_643/A OR2X1_LOC_228/Y 0.01fF
C29889 OR2X1_LOC_203/Y OR2X1_LOC_68/B 0.07fF
C29890 OR2X1_LOC_852/A D_INPUT_0 0.00fF
C29891 AND2X1_LOC_50/a_36_24# INPUT_6 0.00fF
C29892 AND2X1_LOC_31/Y OR2X1_LOC_449/B 0.09fF
C29893 OR2X1_LOC_533/Y AND2X1_LOC_794/B 0.79fF
C29894 OR2X1_LOC_13/Y OR2X1_LOC_12/Y 0.01fF
C29895 AND2X1_LOC_794/B AND2X1_LOC_212/Y 0.01fF
C29896 INPUT_0 AND2X1_LOC_235/a_36_24# 0.00fF
C29897 AND2X1_LOC_799/a_8_24# AND2X1_LOC_436/Y 0.01fF
C29898 OR2X1_LOC_784/a_8_216# OR2X1_LOC_779/B 0.01fF
C29899 OR2X1_LOC_62/B OR2X1_LOC_47/Y 0.02fF
C29900 OR2X1_LOC_267/Y OR2X1_LOC_244/Y 0.01fF
C29901 OR2X1_LOC_176/Y VDD 0.32fF
C29902 D_INPUT_5 AND2X1_LOC_409/B 0.03fF
C29903 AND2X1_LOC_3/Y AND2X1_LOC_751/a_8_24# 0.04fF
C29904 AND2X1_LOC_47/Y AND2X1_LOC_106/a_8_24# 0.09fF
C29905 D_INPUT_3 OR2X1_LOC_417/A 0.08fF
C29906 AND2X1_LOC_831/Y AND2X1_LOC_476/A 0.08fF
C29907 AND2X1_LOC_7/B AND2X1_LOC_92/Y 0.29fF
C29908 OR2X1_LOC_636/A AND2X1_LOC_31/Y 0.01fF
C29909 OR2X1_LOC_45/B AND2X1_LOC_160/Y 0.01fF
C29910 AND2X1_LOC_570/Y AND2X1_LOC_244/A 0.00fF
C29911 AND2X1_LOC_51/Y AND2X1_LOC_52/Y 0.02fF
C29912 OR2X1_LOC_739/A OR2X1_LOC_209/A 0.01fF
C29913 AND2X1_LOC_555/a_36_24# OR2X1_LOC_382/A 0.00fF
C29914 OR2X1_LOC_741/Y OR2X1_LOC_161/B 0.03fF
C29915 OR2X1_LOC_691/a_8_216# VDD 0.21fF
C29916 OR2X1_LOC_161/A OR2X1_LOC_523/a_8_216# 0.01fF
C29917 OR2X1_LOC_9/Y OR2X1_LOC_159/a_8_216# 0.06fF
C29918 OR2X1_LOC_411/Y AND2X1_LOC_219/A 0.06fF
C29919 OR2X1_LOC_9/Y OR2X1_LOC_40/Y 0.76fF
C29920 AND2X1_LOC_48/A OR2X1_LOC_598/A 0.04fF
C29921 OR2X1_LOC_482/Y AND2X1_LOC_499/a_36_24# 0.00fF
C29922 AND2X1_LOC_91/a_8_24# OR2X1_LOC_756/B 0.01fF
C29923 AND2X1_LOC_346/a_8_24# OR2X1_LOC_600/A 0.01fF
C29924 OR2X1_LOC_329/Y AND2X1_LOC_535/Y 0.00fF
C29925 OR2X1_LOC_40/Y AND2X1_LOC_182/a_36_24# 0.00fF
C29926 AND2X1_LOC_483/Y OR2X1_LOC_417/A 0.02fF
C29927 OR2X1_LOC_335/B OR2X1_LOC_318/B 0.16fF
C29928 OR2X1_LOC_121/B AND2X1_LOC_31/Y 0.10fF
C29929 OR2X1_LOC_744/A AND2X1_LOC_828/a_8_24# 0.01fF
C29930 AND2X1_LOC_787/A AND2X1_LOC_722/A 0.00fF
C29931 OR2X1_LOC_269/B OR2X1_LOC_771/B 0.07fF
C29932 AND2X1_LOC_12/Y OR2X1_LOC_605/Y 0.00fF
C29933 OR2X1_LOC_22/Y AND2X1_LOC_562/Y 2.45fF
C29934 OR2X1_LOC_673/A D_INPUT_1 0.01fF
C29935 OR2X1_LOC_151/A AND2X1_LOC_437/a_8_24# 0.01fF
C29936 OR2X1_LOC_468/Y OR2X1_LOC_308/Y 4.36fF
C29937 OR2X1_LOC_469/a_8_216# OR2X1_LOC_469/B 0.03fF
C29938 OR2X1_LOC_709/A OR2X1_LOC_678/Y 0.00fF
C29939 OR2X1_LOC_87/A OR2X1_LOC_727/a_8_216# 0.02fF
C29940 OR2X1_LOC_600/A AND2X1_LOC_447/Y 0.01fF
C29941 OR2X1_LOC_235/B AND2X1_LOC_150/a_8_24# 0.11fF
C29942 VDD OR2X1_LOC_190/A 0.10fF
C29943 OR2X1_LOC_70/Y OR2X1_LOC_13/B 0.33fF
C29944 OR2X1_LOC_96/Y OR2X1_LOC_56/A 0.01fF
C29945 AND2X1_LOC_803/B OR2X1_LOC_679/Y 0.01fF
C29946 OR2X1_LOC_51/B OR2X1_LOC_3/B 0.21fF
C29947 AND2X1_LOC_173/a_8_24# OR2X1_LOC_161/B 0.00fF
C29948 AND2X1_LOC_191/B AND2X1_LOC_709/a_8_24# 0.04fF
C29949 OR2X1_LOC_185/A OR2X1_LOC_563/A 0.04fF
C29950 OR2X1_LOC_427/A AND2X1_LOC_407/a_8_24# 0.04fF
C29951 AND2X1_LOC_421/a_8_24# OR2X1_LOC_713/A 0.03fF
C29952 AND2X1_LOC_217/Y OR2X1_LOC_91/A 2.81fF
C29953 OR2X1_LOC_776/Y OR2X1_LOC_78/A 0.43fF
C29954 OR2X1_LOC_3/Y AND2X1_LOC_789/Y 0.03fF
C29955 OR2X1_LOC_71/Y AND2X1_LOC_772/a_8_24# 0.01fF
C29956 VDD AND2X1_LOC_94/Y 0.40fF
C29957 OR2X1_LOC_323/A OR2X1_LOC_6/A 0.02fF
C29958 AND2X1_LOC_733/Y AND2X1_LOC_778/Y 0.00fF
C29959 OR2X1_LOC_235/B OR2X1_LOC_813/a_8_216# 0.00fF
C29960 OR2X1_LOC_177/Y AND2X1_LOC_486/Y 0.03fF
C29961 OR2X1_LOC_158/A AND2X1_LOC_335/a_36_24# 0.01fF
C29962 AND2X1_LOC_22/Y AND2X1_LOC_132/a_8_24# 0.02fF
C29963 OR2X1_LOC_502/A OR2X1_LOC_646/B 0.03fF
C29964 OR2X1_LOC_161/A OR2X1_LOC_576/A 0.03fF
C29965 AND2X1_LOC_722/a_8_24# OR2X1_LOC_164/Y 0.00fF
C29966 OR2X1_LOC_631/B OR2X1_LOC_556/a_8_216# 0.41fF
C29967 OR2X1_LOC_866/B OR2X1_LOC_848/a_8_216# 0.06fF
C29968 OR2X1_LOC_185/A OR2X1_LOC_738/a_8_216# 0.06fF
C29969 AND2X1_LOC_88/Y OR2X1_LOC_608/Y 0.09fF
C29970 AND2X1_LOC_738/B AND2X1_LOC_663/A 0.10fF
C29971 OR2X1_LOC_156/B OR2X1_LOC_160/A 0.01fF
C29972 OR2X1_LOC_158/A OR2X1_LOC_837/A 0.03fF
C29973 OR2X1_LOC_622/a_8_216# OR2X1_LOC_622/B 0.47fF
C29974 OR2X1_LOC_41/a_8_216# OR2X1_LOC_311/a_8_216# 0.47fF
C29975 OR2X1_LOC_35/B AND2X1_LOC_36/Y 0.14fF
C29976 OR2X1_LOC_56/A AND2X1_LOC_663/A 0.10fF
C29977 OR2X1_LOC_36/Y OR2X1_LOC_56/Y 0.01fF
C29978 AND2X1_LOC_64/Y OR2X1_LOC_68/a_8_216# 0.01fF
C29979 AND2X1_LOC_538/a_8_24# OR2X1_LOC_13/B 0.01fF
C29980 AND2X1_LOC_509/Y AND2X1_LOC_510/A 0.02fF
C29981 OR2X1_LOC_840/A AND2X1_LOC_110/Y 0.05fF
C29982 AND2X1_LOC_707/Y AND2X1_LOC_319/A 0.07fF
C29983 AND2X1_LOC_564/A AND2X1_LOC_564/a_8_24# 0.05fF
C29984 OR2X1_LOC_76/a_8_216# OR2X1_LOC_241/B 0.03fF
C29985 AND2X1_LOC_428/a_8_24# OR2X1_LOC_451/B 0.01fF
C29986 OR2X1_LOC_314/a_8_216# OR2X1_LOC_604/A 0.01fF
C29987 OR2X1_LOC_538/a_36_216# OR2X1_LOC_160/B 0.00fF
C29988 AND2X1_LOC_70/Y OR2X1_LOC_294/a_8_216# 0.01fF
C29989 OR2X1_LOC_48/B AND2X1_LOC_476/Y 0.02fF
C29990 OR2X1_LOC_151/A OR2X1_LOC_623/a_8_216# 0.03fF
C29991 OR2X1_LOC_109/Y OR2X1_LOC_322/a_36_216# 0.01fF
C29992 AND2X1_LOC_50/Y VDD 0.40fF
C29993 AND2X1_LOC_452/Y OR2X1_LOC_604/Y 0.05fF
C29994 OR2X1_LOC_496/Y OR2X1_LOC_406/Y 0.71fF
C29995 OR2X1_LOC_26/Y AND2X1_LOC_287/B 0.02fF
C29996 OR2X1_LOC_756/B OR2X1_LOC_78/A 0.33fF
C29997 OR2X1_LOC_18/Y AND2X1_LOC_476/Y 0.03fF
C29998 AND2X1_LOC_362/B OR2X1_LOC_18/Y 0.00fF
C29999 AND2X1_LOC_51/Y AND2X1_LOC_238/a_36_24# 0.01fF
C30000 OR2X1_LOC_814/A OR2X1_LOC_590/Y 0.02fF
C30001 OR2X1_LOC_865/A OR2X1_LOC_810/A 0.05fF
C30002 OR2X1_LOC_364/A AND2X1_LOC_438/a_8_24# 0.01fF
C30003 AND2X1_LOC_367/A AND2X1_LOC_474/A 0.05fF
C30004 OR2X1_LOC_158/A AND2X1_LOC_34/Y 0.04fF
C30005 AND2X1_LOC_322/a_36_24# OR2X1_LOC_620/Y 0.01fF
C30006 OR2X1_LOC_319/B AND2X1_LOC_92/Y 1.75fF
C30007 AND2X1_LOC_707/Y OR2X1_LOC_682/a_36_216# -0.01fF
C30008 OR2X1_LOC_158/A AND2X1_LOC_114/a_8_24# 0.02fF
C30009 AND2X1_LOC_572/a_8_24# AND2X1_LOC_489/Y 0.01fF
C30010 OR2X1_LOC_850/a_8_216# OR2X1_LOC_756/B 0.01fF
C30011 OR2X1_LOC_833/Y OR2X1_LOC_87/A 0.01fF
C30012 OR2X1_LOC_710/A OR2X1_LOC_705/Y 0.03fF
C30013 OR2X1_LOC_841/a_36_216# AND2X1_LOC_92/Y 0.01fF
C30014 AND2X1_LOC_456/Y AND2X1_LOC_456/a_8_24# 0.01fF
C30015 AND2X1_LOC_364/A OR2X1_LOC_426/B -0.08fF
C30016 AND2X1_LOC_217/Y AND2X1_LOC_573/A 0.00fF
C30017 OR2X1_LOC_109/Y OR2X1_LOC_600/A 0.07fF
C30018 OR2X1_LOC_57/Y AND2X1_LOC_198/a_8_24# 0.23fF
C30019 AND2X1_LOC_69/a_8_24# AND2X1_LOC_36/Y 0.10fF
C30020 OR2X1_LOC_89/A OR2X1_LOC_816/A 0.12fF
C30021 OR2X1_LOC_318/Y AND2X1_LOC_92/Y 0.03fF
C30022 OR2X1_LOC_160/B OR2X1_LOC_541/B 0.01fF
C30023 AND2X1_LOC_2/Y AND2X1_LOC_11/Y 0.44fF
C30024 OR2X1_LOC_9/Y OR2X1_LOC_618/a_8_216# 0.01fF
C30025 AND2X1_LOC_340/a_8_24# OR2X1_LOC_39/A 0.01fF
C30026 AND2X1_LOC_219/a_8_24# OR2X1_LOC_619/Y 0.04fF
C30027 OR2X1_LOC_619/Y AND2X1_LOC_447/Y 0.07fF
C30028 OR2X1_LOC_793/A OR2X1_LOC_596/A 0.02fF
C30029 AND2X1_LOC_860/A OR2X1_LOC_39/A 0.01fF
C30030 AND2X1_LOC_717/B AND2X1_LOC_464/A 0.00fF
C30031 AND2X1_LOC_721/Y AND2X1_LOC_578/A 0.03fF
C30032 VDD AND2X1_LOC_447/a_8_24# -0.00fF
C30033 D_INPUT_3 AND2X1_LOC_247/a_8_24# 0.03fF
C30034 OR2X1_LOC_276/B OR2X1_LOC_777/B 0.07fF
C30035 OR2X1_LOC_235/B OR2X1_LOC_575/A 0.37fF
C30036 OR2X1_LOC_39/A OR2X1_LOC_626/Y 0.34fF
C30037 OR2X1_LOC_159/a_8_216# OR2X1_LOC_96/B 0.01fF
C30038 AND2X1_LOC_40/Y OR2X1_LOC_663/A 0.03fF
C30039 OR2X1_LOC_680/A AND2X1_LOC_806/a_8_24# 0.03fF
C30040 OR2X1_LOC_648/A OR2X1_LOC_624/A 0.10fF
C30041 VDD OR2X1_LOC_265/Y 0.67fF
C30042 OR2X1_LOC_185/Y AND2X1_LOC_131/a_8_24# 0.26fF
C30043 AND2X1_LOC_624/A AND2X1_LOC_657/Y 7.73fF
C30044 OR2X1_LOC_74/A AND2X1_LOC_727/B 0.03fF
C30045 AND2X1_LOC_622/a_8_24# AND2X1_LOC_658/Y 0.20fF
C30046 AND2X1_LOC_22/Y AND2X1_LOC_18/a_36_24# 0.00fF
C30047 OR2X1_LOC_474/Y OR2X1_LOC_475/a_8_216# 0.01fF
C30048 AND2X1_LOC_117/a_8_24# AND2X1_LOC_44/Y 0.01fF
C30049 OR2X1_LOC_203/Y AND2X1_LOC_626/a_36_24# 0.00fF
C30050 OR2X1_LOC_630/a_8_216# OR2X1_LOC_630/B 0.05fF
C30051 AND2X1_LOC_191/B AND2X1_LOC_624/A 0.00fF
C30052 OR2X1_LOC_426/B AND2X1_LOC_572/A 0.01fF
C30053 OR2X1_LOC_124/B OR2X1_LOC_204/Y 0.08fF
C30054 OR2X1_LOC_186/Y AND2X1_LOC_528/a_36_24# 0.00fF
C30055 AND2X1_LOC_40/Y AND2X1_LOC_503/a_8_24# 0.01fF
C30056 OR2X1_LOC_485/A OR2X1_LOC_829/A 0.19fF
C30057 AND2X1_LOC_624/A AND2X1_LOC_469/B 0.03fF
C30058 OR2X1_LOC_40/Y AND2X1_LOC_852/Y 0.05fF
C30059 OR2X1_LOC_517/a_36_216# AND2X1_LOC_76/Y 0.00fF
C30060 AND2X1_LOC_64/Y OR2X1_LOC_814/A 0.18fF
C30061 OR2X1_LOC_805/A AND2X1_LOC_92/Y 0.21fF
C30062 AND2X1_LOC_51/Y OR2X1_LOC_576/A 0.02fF
C30063 OR2X1_LOC_790/B AND2X1_LOC_41/A 0.12fF
C30064 AND2X1_LOC_568/B AND2X1_LOC_661/A 0.67fF
C30065 AND2X1_LOC_716/Y AND2X1_LOC_357/a_8_24# 0.02fF
C30066 AND2X1_LOC_543/a_8_24# OR2X1_LOC_109/Y 0.02fF
C30067 OR2X1_LOC_160/B OR2X1_LOC_849/A 0.04fF
C30068 OR2X1_LOC_160/A OR2X1_LOC_803/a_8_216# 0.01fF
C30069 AND2X1_LOC_41/A OR2X1_LOC_161/A 0.46fF
C30070 AND2X1_LOC_12/Y OR2X1_LOC_634/A 0.02fF
C30071 OR2X1_LOC_6/B AND2X1_LOC_3/Y 0.49fF
C30072 AND2X1_LOC_366/A AND2X1_LOC_848/Y 0.03fF
C30073 OR2X1_LOC_620/Y OR2X1_LOC_623/B 0.00fF
C30074 AND2X1_LOC_533/a_8_24# OR2X1_LOC_703/A 0.00fF
C30075 OR2X1_LOC_496/Y OR2X1_LOC_496/a_8_216# 0.01fF
C30076 AND2X1_LOC_555/a_8_24# AND2X1_LOC_345/a_8_24# 0.23fF
C30077 OR2X1_LOC_459/A OR2X1_LOC_39/A 0.09fF
C30078 OR2X1_LOC_106/Y AND2X1_LOC_845/Y -0.01fF
C30079 AND2X1_LOC_251/a_8_24# OR2X1_LOC_561/Y 0.01fF
C30080 AND2X1_LOC_578/A OR2X1_LOC_482/Y 0.30fF
C30081 AND2X1_LOC_571/A AND2X1_LOC_227/Y 0.01fF
C30082 OR2X1_LOC_759/A OR2X1_LOC_665/Y 0.16fF
C30083 AND2X1_LOC_729/a_8_24# AND2X1_LOC_729/B 0.11fF
C30084 OR2X1_LOC_690/Y OR2X1_LOC_753/A 0.09fF
C30085 AND2X1_LOC_340/Y AND2X1_LOC_351/Y 0.20fF
C30086 AND2X1_LOC_339/Y OR2X1_LOC_46/A 0.02fF
C30087 OR2X1_LOC_502/A OR2X1_LOC_506/A 6.75fF
C30088 AND2X1_LOC_486/Y AND2X1_LOC_850/a_8_24# 0.13fF
C30089 AND2X1_LOC_787/a_8_24# AND2X1_LOC_794/A 0.00fF
C30090 OR2X1_LOC_46/A OR2X1_LOC_414/Y 0.01fF
C30091 AND2X1_LOC_500/Y OR2X1_LOC_239/a_8_216# 0.48fF
C30092 AND2X1_LOC_471/a_8_24# AND2X1_LOC_786/Y 0.02fF
C30093 OR2X1_LOC_804/A AND2X1_LOC_36/Y 0.01fF
C30094 OR2X1_LOC_395/Y OR2X1_LOC_396/a_36_216# 0.00fF
C30095 OR2X1_LOC_821/Y OR2X1_LOC_54/Y 0.00fF
C30096 INPUT_0 OR2X1_LOC_83/A 0.05fF
C30097 OR2X1_LOC_731/a_8_216# OR2X1_LOC_738/A 0.03fF
C30098 OR2X1_LOC_112/B OR2X1_LOC_390/B 0.02fF
C30099 AND2X1_LOC_155/a_8_24# OR2X1_LOC_39/A 0.01fF
C30100 OR2X1_LOC_185/Y OR2X1_LOC_435/a_36_216# 0.02fF
C30101 OR2X1_LOC_3/Y OR2X1_LOC_426/B 1.56fF
C30102 OR2X1_LOC_51/Y OR2X1_LOC_371/Y 0.07fF
C30103 OR2X1_LOC_154/A OR2X1_LOC_623/B 0.07fF
C30104 AND2X1_LOC_338/a_8_24# AND2X1_LOC_640/Y 0.00fF
C30105 OR2X1_LOC_763/a_8_216# OR2X1_LOC_44/Y 0.01fF
C30106 OR2X1_LOC_600/A AND2X1_LOC_729/B 0.03fF
C30107 OR2X1_LOC_364/A AND2X1_LOC_40/Y 0.07fF
C30108 OR2X1_LOC_329/a_8_216# OR2X1_LOC_22/Y 0.02fF
C30109 OR2X1_LOC_185/Y AND2X1_LOC_40/Y 0.03fF
C30110 OR2X1_LOC_777/B OR2X1_LOC_779/B 0.02fF
C30111 OR2X1_LOC_810/A OR2X1_LOC_391/A 0.06fF
C30112 OR2X1_LOC_756/B OR2X1_LOC_155/A 0.03fF
C30113 AND2X1_LOC_331/a_8_24# AND2X1_LOC_56/B 0.04fF
C30114 AND2X1_LOC_201/a_36_24# AND2X1_LOC_201/Y 0.00fF
C30115 OR2X1_LOC_160/A OR2X1_LOC_231/a_8_216# 0.04fF
C30116 VDD OR2X1_LOC_473/Y 0.22fF
C30117 AND2X1_LOC_38/a_8_24# OR2X1_LOC_78/B 0.04fF
C30118 OR2X1_LOC_451/a_8_216# OR2X1_LOC_451/A 0.47fF
C30119 AND2X1_LOC_863/a_36_24# OR2X1_LOC_36/Y 0.00fF
C30120 OR2X1_LOC_619/Y AND2X1_LOC_448/Y 0.02fF
C30121 OR2X1_LOC_167/Y AND2X1_LOC_810/B 0.03fF
C30122 OR2X1_LOC_207/B AND2X1_LOC_47/Y 0.01fF
C30123 OR2X1_LOC_36/Y AND2X1_LOC_642/Y 0.01fF
C30124 OR2X1_LOC_864/A OR2X1_LOC_489/a_8_216# 0.01fF
C30125 OR2X1_LOC_520/Y AND2X1_LOC_517/a_8_24# 0.02fF
C30126 AND2X1_LOC_154/a_8_24# AND2X1_LOC_621/Y 0.26fF
C30127 OR2X1_LOC_739/B OR2X1_LOC_221/a_36_216# 0.03fF
C30128 OR2X1_LOC_538/A AND2X1_LOC_111/a_8_24# 0.21fF
C30129 OR2X1_LOC_774/Y OR2X1_LOC_489/a_8_216# 0.00fF
C30130 AND2X1_LOC_76/a_36_24# OR2X1_LOC_85/A 0.00fF
C30131 OR2X1_LOC_541/B OR2X1_LOC_553/A 0.01fF
C30132 OR2X1_LOC_278/Y OR2X1_LOC_44/Y 0.03fF
C30133 AND2X1_LOC_214/A AND2X1_LOC_196/a_8_24# 0.17fF
C30134 OR2X1_LOC_756/B OR2X1_LOC_392/a_8_216# 0.01fF
C30135 AND2X1_LOC_429/a_36_24# INPUT_6 0.00fF
C30136 OR2X1_LOC_641/Y OR2X1_LOC_643/Y 0.26fF
C30137 AND2X1_LOC_59/Y AND2X1_LOC_395/a_8_24# 0.09fF
C30138 OR2X1_LOC_715/B OR2X1_LOC_532/B 8.09fF
C30139 AND2X1_LOC_779/a_8_24# OR2X1_LOC_52/B 0.03fF
C30140 OR2X1_LOC_45/Y OR2X1_LOC_26/Y 0.02fF
C30141 AND2X1_LOC_733/a_8_24# OR2X1_LOC_74/A 0.04fF
C30142 OR2X1_LOC_276/B OR2X1_LOC_344/A 0.02fF
C30143 OR2X1_LOC_53/Y OR2X1_LOC_41/a_8_216# 0.00fF
C30144 OR2X1_LOC_160/B OR2X1_LOC_707/B 0.26fF
C30145 AND2X1_LOC_542/a_36_24# OR2X1_LOC_31/Y -0.00fF
C30146 AND2X1_LOC_40/Y AND2X1_LOC_171/a_36_24# 0.01fF
C30147 OR2X1_LOC_465/a_8_216# OR2X1_LOC_375/A 0.03fF
C30148 AND2X1_LOC_41/A AND2X1_LOC_51/Y 0.61fF
C30149 OR2X1_LOC_631/B OR2X1_LOC_161/A 0.03fF
C30150 AND2X1_LOC_677/a_8_24# OR2X1_LOC_78/A 0.01fF
C30151 AND2X1_LOC_724/A OR2X1_LOC_47/Y 0.15fF
C30152 AND2X1_LOC_566/B AND2X1_LOC_866/A 0.02fF
C30153 AND2X1_LOC_357/B AND2X1_LOC_863/Y 0.01fF
C30154 AND2X1_LOC_843/a_8_24# OR2X1_LOC_26/Y 0.02fF
C30155 OR2X1_LOC_185/A AND2X1_LOC_252/a_8_24# 0.17fF
C30156 AND2X1_LOC_47/Y OR2X1_LOC_772/A 0.01fF
C30157 AND2X1_LOC_862/a_8_24# AND2X1_LOC_862/A 0.10fF
C30158 OR2X1_LOC_22/A OR2X1_LOC_380/Y 0.02fF
C30159 AND2X1_LOC_191/B AND2X1_LOC_621/a_8_24# 0.01fF
C30160 AND2X1_LOC_553/a_8_24# OR2X1_LOC_95/Y 0.01fF
C30161 OR2X1_LOC_265/Y AND2X1_LOC_267/a_8_24# 0.25fF
C30162 OR2X1_LOC_188/Y OR2X1_LOC_76/a_8_216# 0.01fF
C30163 OR2X1_LOC_7/Y OR2X1_LOC_56/A 0.03fF
C30164 OR2X1_LOC_95/a_8_216# OR2X1_LOC_44/Y 0.06fF
C30165 OR2X1_LOC_476/B OR2X1_LOC_174/A 0.00fF
C30166 AND2X1_LOC_629/Y AND2X1_LOC_629/a_36_24# 0.00fF
C30167 AND2X1_LOC_168/Y AND2X1_LOC_566/Y 0.02fF
C30168 AND2X1_LOC_539/Y OR2X1_LOC_761/a_8_216# 0.01fF
C30169 OR2X1_LOC_88/A OR2X1_LOC_262/a_8_216# 0.47fF
C30170 OR2X1_LOC_508/A AND2X1_LOC_51/Y 0.15fF
C30171 OR2X1_LOC_160/B OR2X1_LOC_440/A 0.01fF
C30172 AND2X1_LOC_91/B OR2X1_LOC_228/Y 0.10fF
C30173 OR2X1_LOC_36/Y OR2X1_LOC_591/A 0.00fF
C30174 OR2X1_LOC_235/B OR2X1_LOC_62/a_36_216# 0.00fF
C30175 AND2X1_LOC_673/a_8_24# OR2X1_LOC_85/A 0.03fF
C30176 OR2X1_LOC_26/Y OR2X1_LOC_824/Y 0.44fF
C30177 OR2X1_LOC_431/a_8_216# OR2X1_LOC_48/B 0.01fF
C30178 AND2X1_LOC_42/B AND2X1_LOC_43/B 0.20fF
C30179 AND2X1_LOC_459/Y OR2X1_LOC_378/Y 0.01fF
C30180 AND2X1_LOC_76/Y OR2X1_LOC_275/a_8_216# 0.01fF
C30181 AND2X1_LOC_530/a_8_24# OR2X1_LOC_598/A 0.01fF
C30182 AND2X1_LOC_143/a_8_24# OR2X1_LOC_62/B 0.01fF
C30183 INPUT_0 AND2X1_LOC_831/Y 0.07fF
C30184 OR2X1_LOC_92/Y OR2X1_LOC_46/A 0.02fF
C30185 OR2X1_LOC_479/Y OR2X1_LOC_375/A 0.03fF
C30186 OR2X1_LOC_574/A OR2X1_LOC_87/A 0.03fF
C30187 AND2X1_LOC_339/B AND2X1_LOC_643/a_8_24# 0.01fF
C30188 AND2X1_LOC_135/a_8_24# OR2X1_LOC_161/A -0.06fF
C30189 OR2X1_LOC_857/A AND2X1_LOC_31/Y 0.05fF
C30190 AND2X1_LOC_56/B AND2X1_LOC_329/a_36_24# 0.00fF
C30191 OR2X1_LOC_40/Y AND2X1_LOC_647/B 1.05fF
C30192 OR2X1_LOC_74/A OR2X1_LOC_85/A 1.26fF
C30193 AND2X1_LOC_681/a_8_24# OR2X1_LOC_78/B 0.03fF
C30194 VDD OR2X1_LOC_214/B 0.15fF
C30195 OR2X1_LOC_89/A OR2X1_LOC_591/a_8_216# 0.01fF
C30196 AND2X1_LOC_560/B AND2X1_LOC_276/Y 0.03fF
C30197 OR2X1_LOC_481/a_8_216# OR2X1_LOC_748/A 0.00fF
C30198 OR2X1_LOC_273/Y AND2X1_LOC_831/a_8_24# 0.23fF
C30199 AND2X1_LOC_59/Y OR2X1_LOC_476/a_8_216# 0.01fF
C30200 OR2X1_LOC_19/B AND2X1_LOC_403/B 1.46fF
C30201 OR2X1_LOC_22/Y OR2X1_LOC_432/Y 0.04fF
C30202 OR2X1_LOC_285/B OR2X1_LOC_285/A 0.05fF
C30203 AND2X1_LOC_554/B OR2X1_LOC_585/A 0.02fF
C30204 AND2X1_LOC_792/B OR2X1_LOC_759/Y 0.10fF
C30205 OR2X1_LOC_22/Y AND2X1_LOC_287/a_8_24# 0.06fF
C30206 OR2X1_LOC_799/A AND2X1_LOC_165/a_8_24# 0.23fF
C30207 OR2X1_LOC_462/B OR2X1_LOC_462/a_8_216# 0.02fF
C30208 AND2X1_LOC_48/A OR2X1_LOC_341/Y 0.01fF
C30209 AND2X1_LOC_227/Y OR2X1_LOC_92/Y 0.05fF
C30210 AND2X1_LOC_612/B AND2X1_LOC_612/a_36_24# 0.00fF
C30211 OR2X1_LOC_436/B OR2X1_LOC_436/Y 0.76fF
C30212 AND2X1_LOC_709/a_8_24# AND2X1_LOC_848/A -0.01fF
C30213 D_INPUT_3 AND2X1_LOC_402/a_8_24# 0.26fF
C30214 AND2X1_LOC_12/Y OR2X1_LOC_335/B 0.03fF
C30215 OR2X1_LOC_36/Y AND2X1_LOC_307/Y 0.15fF
C30216 AND2X1_LOC_95/Y AND2X1_LOC_53/Y 0.12fF
C30217 AND2X1_LOC_170/B AND2X1_LOC_841/B 0.01fF
C30218 OR2X1_LOC_64/Y AND2X1_LOC_806/A 0.02fF
C30219 OR2X1_LOC_3/Y OR2X1_LOC_743/A 13.39fF
C30220 OR2X1_LOC_80/a_8_216# OR2X1_LOC_393/Y 0.40fF
C30221 OR2X1_LOC_686/A AND2X1_LOC_430/B 0.00fF
C30222 OR2X1_LOC_502/A OR2X1_LOC_227/Y 0.03fF
C30223 OR2X1_LOC_275/a_8_216# OR2X1_LOC_52/B 0.02fF
C30224 OR2X1_LOC_864/A OR2X1_LOC_121/B 0.03fF
C30225 AND2X1_LOC_104/a_8_24# AND2X1_LOC_47/Y 0.02fF
C30226 AND2X1_LOC_56/B AND2X1_LOC_825/a_8_24# 0.03fF
C30227 OR2X1_LOC_19/B OR2X1_LOC_82/a_36_216# 0.01fF
C30228 OR2X1_LOC_479/Y OR2X1_LOC_605/B 0.02fF
C30229 OR2X1_LOC_51/Y AND2X1_LOC_222/Y 0.04fF
C30230 OR2X1_LOC_632/a_8_216# OR2X1_LOC_598/A 0.04fF
C30231 OR2X1_LOC_502/A D_INPUT_1 0.09fF
C30232 AND2X1_LOC_727/A OR2X1_LOC_26/Y 0.03fF
C30233 OR2X1_LOC_643/A OR2X1_LOC_849/a_36_216# -0.00fF
C30234 OR2X1_LOC_817/Y AND2X1_LOC_847/a_8_24# 0.23fF
C30235 OR2X1_LOC_47/Y OR2X1_LOC_393/a_8_216# 0.01fF
C30236 AND2X1_LOC_227/Y OR2X1_LOC_65/B 0.52fF
C30237 AND2X1_LOC_852/a_8_24# D_INPUT_0 0.01fF
C30238 OR2X1_LOC_160/A OR2X1_LOC_783/A 0.03fF
C30239 AND2X1_LOC_56/a_36_24# OR2X1_LOC_375/A 0.00fF
C30240 AND2X1_LOC_95/Y OR2X1_LOC_223/A 0.07fF
C30241 OR2X1_LOC_709/A OR2X1_LOC_777/B 0.02fF
C30242 OR2X1_LOC_92/Y OR2X1_LOC_813/Y 0.10fF
C30243 AND2X1_LOC_727/A OR2X1_LOC_89/A 0.03fF
C30244 OR2X1_LOC_199/a_8_216# AND2X1_LOC_36/Y 0.06fF
C30245 AND2X1_LOC_649/Y AND2X1_LOC_655/A 0.27fF
C30246 OR2X1_LOC_440/A OR2X1_LOC_553/A 0.01fF
C30247 OR2X1_LOC_502/A AND2X1_LOC_48/Y 0.02fF
C30248 AND2X1_LOC_1/Y OR2X1_LOC_636/a_8_216# 0.01fF
C30249 AND2X1_LOC_139/B AND2X1_LOC_476/A 0.07fF
C30250 AND2X1_LOC_598/a_8_24# OR2X1_LOC_95/Y 0.01fF
C30251 AND2X1_LOC_59/Y AND2X1_LOC_813/a_8_24# 0.17fF
C30252 OR2X1_LOC_19/B OR2X1_LOC_20/a_8_216# 0.14fF
C30253 OR2X1_LOC_78/B OR2X1_LOC_68/B 0.55fF
C30254 OR2X1_LOC_3/Y OR2X1_LOC_246/A 0.26fF
C30255 OR2X1_LOC_654/A D_INPUT_0 0.17fF
C30256 OR2X1_LOC_26/Y OR2X1_LOC_95/Y 2.31fF
C30257 OR2X1_LOC_486/Y OR2X1_LOC_212/B 0.05fF
C30258 OR2X1_LOC_92/Y OR2X1_LOC_753/Y 0.01fF
C30259 AND2X1_LOC_47/Y AND2X1_LOC_292/a_36_24# 0.00fF
C30260 OR2X1_LOC_59/Y OR2X1_LOC_533/a_8_216# -0.00fF
C30261 OR2X1_LOC_335/Y OR2X1_LOC_578/B 0.00fF
C30262 OR2X1_LOC_3/Y OR2X1_LOC_225/a_8_216# 0.01fF
C30263 OR2X1_LOC_628/Y AND2X1_LOC_632/a_8_24# 0.03fF
C30264 OR2X1_LOC_542/B OR2X1_LOC_367/a_8_216# 0.06fF
C30265 OR2X1_LOC_841/a_8_216# AND2X1_LOC_31/Y 0.01fF
C30266 AND2X1_LOC_190/a_8_24# OR2X1_LOC_437/A -0.01fF
C30267 OR2X1_LOC_624/B AND2X1_LOC_15/a_8_24# 0.04fF
C30268 AND2X1_LOC_47/Y AND2X1_LOC_3/Y 2.45fF
C30269 GATE_366 OR2X1_LOC_47/Y 0.01fF
C30270 AND2X1_LOC_47/Y OR2X1_LOC_647/B 0.08fF
C30271 OR2X1_LOC_403/a_8_216# AND2X1_LOC_51/Y 0.01fF
C30272 AND2X1_LOC_12/Y OR2X1_LOC_366/a_8_216# 0.01fF
C30273 OR2X1_LOC_89/A OR2X1_LOC_95/Y 0.13fF
C30274 AND2X1_LOC_40/Y OR2X1_LOC_568/A 0.01fF
C30275 AND2X1_LOC_95/Y OR2X1_LOC_351/a_36_216# 0.00fF
C30276 OR2X1_LOC_427/A OR2X1_LOC_754/Y 0.02fF
C30277 AND2X1_LOC_70/Y OR2X1_LOC_777/B 0.06fF
C30278 AND2X1_LOC_841/B OR2X1_LOC_331/Y 0.03fF
C30279 AND2X1_LOC_40/Y OR2X1_LOC_578/B 0.03fF
C30280 OR2X1_LOC_3/Y OR2X1_LOC_409/B 0.03fF
C30281 OR2X1_LOC_856/B AND2X1_LOC_31/Y 0.08fF
C30282 OR2X1_LOC_516/Y AND2X1_LOC_784/Y 0.37fF
C30283 OR2X1_LOC_206/A OR2X1_LOC_814/A 0.03fF
C30284 OR2X1_LOC_312/Y OR2X1_LOC_47/Y 0.04fF
C30285 OR2X1_LOC_279/Y AND2X1_LOC_859/B 0.80fF
C30286 VDD OR2X1_LOC_183/a_8_216# 0.21fF
C30287 OR2X1_LOC_485/A OR2X1_LOC_224/Y 0.01fF
C30288 OR2X1_LOC_62/a_8_216# OR2X1_LOC_46/A 0.01fF
C30289 OR2X1_LOC_160/B AND2X1_LOC_238/a_8_24# 0.01fF
C30290 OR2X1_LOC_419/Y OR2X1_LOC_591/A 0.02fF
C30291 OR2X1_LOC_64/Y AND2X1_LOC_831/Y 0.41fF
C30292 OR2X1_LOC_85/A AND2X1_LOC_647/Y 0.02fF
C30293 AND2X1_LOC_292/a_8_24# AND2X1_LOC_72/B 0.01fF
C30294 OR2X1_LOC_756/B D_GATE_366 0.03fF
C30295 AND2X1_LOC_605/Y OR2X1_LOC_424/Y 0.07fF
C30296 OR2X1_LOC_680/A AND2X1_LOC_222/Y 0.03fF
C30297 AND2X1_LOC_748/a_8_24# OR2X1_LOC_789/A 0.00fF
C30298 OR2X1_LOC_440/a_8_216# OR2X1_LOC_168/Y 0.01fF
C30299 AND2X1_LOC_719/Y AND2X1_LOC_465/A 0.10fF
C30300 OR2X1_LOC_485/A OR2X1_LOC_597/Y 0.01fF
C30301 OR2X1_LOC_17/Y OR2X1_LOC_588/A 0.00fF
C30302 OR2X1_LOC_375/A OR2X1_LOC_68/B 0.26fF
C30303 OR2X1_LOC_49/A OR2X1_LOC_12/Y 0.01fF
C30304 OR2X1_LOC_420/a_36_216# OR2X1_LOC_419/Y 0.00fF
C30305 OR2X1_LOC_62/A OR2X1_LOC_415/A 0.01fF
C30306 OR2X1_LOC_177/Y AND2X1_LOC_457/a_8_24# 0.00fF
C30307 OR2X1_LOC_429/Y OR2X1_LOC_581/a_8_216# 0.05fF
C30308 OR2X1_LOC_412/a_8_216# OR2X1_LOC_31/Y 0.01fF
C30309 OR2X1_LOC_710/B OR2X1_LOC_710/A 0.16fF
C30310 OR2X1_LOC_45/B OR2X1_LOC_421/Y 0.24fF
C30311 AND2X1_LOC_3/Y OR2X1_LOC_598/A 0.70fF
C30312 AND2X1_LOC_459/Y OR2X1_LOC_378/A 0.19fF
C30313 AND2X1_LOC_573/A OR2X1_LOC_399/a_8_216# 0.01fF
C30314 OR2X1_LOC_255/a_8_216# OR2X1_LOC_256/A 0.01fF
C30315 AND2X1_LOC_851/B AND2X1_LOC_465/Y 0.09fF
C30316 AND2X1_LOC_64/Y OR2X1_LOC_244/Y 0.03fF
C30317 AND2X1_LOC_787/A OR2X1_LOC_40/Y 0.03fF
C30318 AND2X1_LOC_831/Y OR2X1_LOC_417/A 0.02fF
C30319 OR2X1_LOC_833/Y OR2X1_LOC_840/a_8_216# 0.10fF
C30320 OR2X1_LOC_188/Y VDD 0.49fF
C30321 OR2X1_LOC_325/a_36_216# OR2X1_LOC_532/Y 0.00fF
C30322 OR2X1_LOC_78/A OR2X1_LOC_140/B 0.05fF
C30323 OR2X1_LOC_304/a_8_216# VDD 0.21fF
C30324 OR2X1_LOC_78/A OR2X1_LOC_170/a_36_216# 0.01fF
C30325 OR2X1_LOC_151/A OR2X1_LOC_294/Y 0.02fF
C30326 OR2X1_LOC_624/A OR2X1_LOC_112/A 0.15fF
C30327 OR2X1_LOC_403/A AND2X1_LOC_36/Y 0.01fF
C30328 AND2X1_LOC_712/Y OR2X1_LOC_12/Y 0.00fF
C30329 AND2X1_LOC_48/A D_INPUT_1 0.00fF
C30330 OR2X1_LOC_329/Y OR2X1_LOC_16/A 0.04fF
C30331 AND2X1_LOC_522/a_8_24# AND2X1_LOC_18/Y 0.03fF
C30332 AND2X1_LOC_64/Y OR2X1_LOC_501/B 0.03fF
C30333 AND2X1_LOC_91/B AND2X1_LOC_320/a_8_24# 0.00fF
C30334 OR2X1_LOC_650/a_8_216# AND2X1_LOC_7/B 0.05fF
C30335 OR2X1_LOC_696/A OR2X1_LOC_256/Y 0.12fF
C30336 AND2X1_LOC_181/Y AND2X1_LOC_476/Y 0.51fF
C30337 AND2X1_LOC_752/a_8_24# AND2X1_LOC_409/B 0.04fF
C30338 OR2X1_LOC_64/Y AND2X1_LOC_486/a_8_24# 0.01fF
C30339 OR2X1_LOC_526/Y OR2X1_LOC_12/Y 0.01fF
C30340 OR2X1_LOC_411/A OR2X1_LOC_16/A 0.02fF
C30341 AND2X1_LOC_48/A AND2X1_LOC_48/Y 0.01fF
C30342 OR2X1_LOC_566/A OR2X1_LOC_703/A 0.01fF
C30343 OR2X1_LOC_62/B AND2X1_LOC_72/B 0.05fF
C30344 OR2X1_LOC_447/a_8_216# AND2X1_LOC_36/Y 0.01fF
C30345 OR2X1_LOC_31/Y AND2X1_LOC_687/a_8_24# 0.01fF
C30346 OR2X1_LOC_40/Y AND2X1_LOC_566/B 0.04fF
C30347 OR2X1_LOC_106/a_8_216# AND2X1_LOC_243/Y 0.04fF
C30348 OR2X1_LOC_59/Y OR2X1_LOC_428/A 1.12fF
C30349 OR2X1_LOC_160/A OR2X1_LOC_308/Y 0.04fF
C30350 AND2X1_LOC_707/Y AND2X1_LOC_605/Y 0.08fF
C30351 AND2X1_LOC_64/Y OR2X1_LOC_147/B 0.04fF
C30352 OR2X1_LOC_130/A AND2X1_LOC_36/Y 0.00fF
C30353 OR2X1_LOC_59/Y OR2X1_LOC_595/A 0.04fF
C30354 OR2X1_LOC_468/Y OR2X1_LOC_535/a_36_216# 0.00fF
C30355 OR2X1_LOC_70/Y OR2X1_LOC_533/a_8_216# 0.01fF
C30356 OR2X1_LOC_121/a_8_216# AND2X1_LOC_41/A 0.01fF
C30357 OR2X1_LOC_235/B OR2X1_LOC_161/B 0.03fF
C30358 AND2X1_LOC_71/a_8_24# AND2X1_LOC_44/Y 0.01fF
C30359 OR2X1_LOC_95/Y OR2X1_LOC_419/a_8_216# 0.01fF
C30360 OR2X1_LOC_158/A AND2X1_LOC_160/Y 0.02fF
C30361 OR2X1_LOC_19/B OR2X1_LOC_750/Y 0.01fF
C30362 OR2X1_LOC_618/Y D_INPUT_1 0.01fF
C30363 AND2X1_LOC_25/Y INPUT_6 0.03fF
C30364 VDD OR2X1_LOC_325/B 0.02fF
C30365 AND2X1_LOC_81/B OR2X1_LOC_130/a_8_216# 0.05fF
C30366 AND2X1_LOC_741/a_8_24# AND2X1_LOC_564/A 0.07fF
C30367 VDD OR2X1_LOC_686/B 0.21fF
C30368 OR2X1_LOC_269/B OR2X1_LOC_593/B 2.90fF
C30369 AND2X1_LOC_7/a_8_24# AND2X1_LOC_36/Y 0.01fF
C30370 AND2X1_LOC_70/Y OR2X1_LOC_686/A 0.03fF
C30371 AND2X1_LOC_47/Y OR2X1_LOC_196/a_36_216# 0.00fF
C30372 OR2X1_LOC_725/B OR2X1_LOC_779/A 0.03fF
C30373 OR2X1_LOC_604/A OR2X1_LOC_600/Y 0.01fF
C30374 AND2X1_LOC_17/Y D_INPUT_6 0.09fF
C30375 INPUT_0 OR2X1_LOC_596/a_8_216# 0.01fF
C30376 OR2X1_LOC_493/B OR2X1_LOC_493/a_8_216# 0.01fF
C30377 OR2X1_LOC_329/B OR2X1_LOC_108/a_8_216# 0.03fF
C30378 AND2X1_LOC_476/A OR2X1_LOC_598/A 0.11fF
C30379 OR2X1_LOC_6/B INPUT_0 0.17fF
C30380 AND2X1_LOC_572/a_8_24# AND2X1_LOC_554/Y 0.03fF
C30381 AND2X1_LOC_486/Y AND2X1_LOC_212/Y 0.07fF
C30382 AND2X1_LOC_215/Y OR2X1_LOC_59/Y 0.01fF
C30383 OR2X1_LOC_45/B AND2X1_LOC_662/B 0.40fF
C30384 OR2X1_LOC_422/Y OR2X1_LOC_12/Y 0.01fF
C30385 OR2X1_LOC_274/Y AND2X1_LOC_275/a_8_24# 0.01fF
C30386 OR2X1_LOC_416/Y OR2X1_LOC_300/a_8_216# 0.01fF
C30387 AND2X1_LOC_474/A AND2X1_LOC_860/A 0.01fF
C30388 AND2X1_LOC_345/a_36_24# AND2X1_LOC_789/Y 0.01fF
C30389 OR2X1_LOC_323/A OR2X1_LOC_44/Y 0.03fF
C30390 VDD OR2X1_LOC_471/B -0.00fF
C30391 AND2X1_LOC_554/a_8_24# AND2X1_LOC_572/A 0.15fF
C30392 OR2X1_LOC_733/Y OR2X1_LOC_737/a_8_216# 0.39fF
C30393 OR2X1_LOC_329/B OR2X1_LOC_426/B 0.16fF
C30394 OR2X1_LOC_623/a_36_216# OR2X1_LOC_161/B 0.00fF
C30395 OR2X1_LOC_136/a_8_216# OR2X1_LOC_6/A 0.01fF
C30396 OR2X1_LOC_89/Y OR2X1_LOC_44/Y 0.21fF
C30397 OR2X1_LOC_382/Y OR2X1_LOC_604/A 0.11fF
C30398 AND2X1_LOC_391/a_8_24# OR2X1_LOC_40/Y 0.01fF
C30399 AND2X1_LOC_706/Y OR2X1_LOC_48/B 0.03fF
C30400 AND2X1_LOC_212/Y AND2X1_LOC_811/B 0.01fF
C30401 OR2X1_LOC_814/A OR2X1_LOC_579/a_8_216# 0.01fF
C30402 OR2X1_LOC_49/A OR2X1_LOC_38/a_36_216# 0.02fF
C30403 OR2X1_LOC_538/A AND2X1_LOC_110/a_8_24# 0.09fF
C30404 OR2X1_LOC_185/Y OR2X1_LOC_138/a_8_216# 0.01fF
C30405 AND2X1_LOC_675/Y OR2X1_LOC_56/A 0.00fF
C30406 AND2X1_LOC_191/B OR2X1_LOC_755/a_8_216# 0.01fF
C30407 OR2X1_LOC_574/A OR2X1_LOC_390/B 0.10fF
C30408 AND2X1_LOC_706/Y OR2X1_LOC_18/Y 0.01fF
C30409 VDD OR2X1_LOC_164/Y 0.29fF
C30410 AND2X1_LOC_367/A OR2X1_LOC_51/Y 0.03fF
C30411 AND2X1_LOC_73/a_8_24# INPUT_0 0.02fF
C30412 AND2X1_LOC_138/a_8_24# OR2X1_LOC_12/Y 0.03fF
C30413 OR2X1_LOC_69/A OR2X1_LOC_16/A 0.03fF
C30414 AND2X1_LOC_540/a_8_24# VDD -0.00fF
C30415 OR2X1_LOC_447/Y OR2X1_LOC_704/a_8_216# 0.42fF
C30416 AND2X1_LOC_51/Y INPUT_6 0.07fF
C30417 AND2X1_LOC_372/a_8_24# AND2X1_LOC_92/Y 0.03fF
C30418 OR2X1_LOC_264/Y OR2X1_LOC_160/B 0.03fF
C30419 OR2X1_LOC_744/a_8_216# OR2X1_LOC_44/Y 0.02fF
C30420 VDD OR2X1_LOC_469/Y 0.18fF
C30421 OR2X1_LOC_166/a_36_216# AND2X1_LOC_512/Y 0.00fF
C30422 AND2X1_LOC_91/B OR2X1_LOC_287/B 0.06fF
C30423 AND2X1_LOC_738/B OR2X1_LOC_516/B 0.01fF
C30424 OR2X1_LOC_389/B AND2X1_LOC_7/B 0.03fF
C30425 OR2X1_LOC_114/a_36_216# OR2X1_LOC_632/Y 0.01fF
C30426 AND2X1_LOC_354/B AND2X1_LOC_802/Y 0.10fF
C30427 AND2X1_LOC_53/Y AND2X1_LOC_41/Y 0.15fF
C30428 AND2X1_LOC_553/a_36_24# OR2X1_LOC_427/A 0.01fF
C30429 OR2X1_LOC_71/a_36_216# AND2X1_LOC_243/Y 0.01fF
C30430 OR2X1_LOC_528/Y AND2X1_LOC_621/Y 0.01fF
C30431 OR2X1_LOC_163/A OR2X1_LOC_163/Y 0.01fF
C30432 OR2X1_LOC_40/Y OR2X1_LOC_127/a_8_216# 0.01fF
C30433 AND2X1_LOC_702/Y OR2X1_LOC_16/A 0.03fF
C30434 OR2X1_LOC_62/B AND2X1_LOC_36/Y 0.03fF
C30435 AND2X1_LOC_42/B AND2X1_LOC_416/a_8_24# 0.01fF
C30436 OR2X1_LOC_589/A AND2X1_LOC_319/A 0.19fF
C30437 OR2X1_LOC_687/Y OR2X1_LOC_596/A 0.03fF
C30438 AND2X1_LOC_654/a_8_24# OR2X1_LOC_12/Y 0.01fF
C30439 AND2X1_LOC_599/a_8_24# AND2X1_LOC_387/B 0.03fF
C30440 AND2X1_LOC_784/A AND2X1_LOC_515/a_8_24# 0.03fF
C30441 OR2X1_LOC_114/Y OR2X1_LOC_151/A 0.34fF
C30442 AND2X1_LOC_43/B AND2X1_LOC_411/a_36_24# 0.01fF
C30443 VDD OR2X1_LOC_405/Y 0.19fF
C30444 AND2X1_LOC_481/a_8_24# AND2X1_LOC_279/a_8_24# 0.23fF
C30445 OR2X1_LOC_355/B OR2X1_LOC_355/a_8_216# 0.05fF
C30446 AND2X1_LOC_729/Y OR2X1_LOC_679/a_8_216# 0.01fF
C30447 AND2X1_LOC_259/Y OR2X1_LOC_12/Y 0.00fF
C30448 AND2X1_LOC_25/a_36_24# INPUT_6 0.00fF
C30449 AND2X1_LOC_3/Y AND2X1_LOC_627/a_36_24# 0.00fF
C30450 OR2X1_LOC_47/Y OR2X1_LOC_13/B 1.41fF
C30451 AND2X1_LOC_711/Y OR2X1_LOC_428/A 0.00fF
C30452 OR2X1_LOC_9/Y AND2X1_LOC_836/a_8_24# 0.01fF
C30453 AND2X1_LOC_847/Y OR2X1_LOC_700/a_36_216# 0.01fF
C30454 AND2X1_LOC_390/B AND2X1_LOC_802/Y 0.01fF
C30455 OR2X1_LOC_70/Y OR2X1_LOC_428/A 0.26fF
C30456 OR2X1_LOC_45/B OR2X1_LOC_273/Y 0.01fF
C30457 AND2X1_LOC_729/Y AND2X1_LOC_658/A 0.03fF
C30458 AND2X1_LOC_110/Y OR2X1_LOC_468/Y 0.03fF
C30459 OR2X1_LOC_53/Y OR2X1_LOC_431/Y 0.01fF
C30460 OR2X1_LOC_497/Y AND2X1_LOC_500/B 0.01fF
C30461 OR2X1_LOC_604/A OR2X1_LOC_591/A 0.03fF
C30462 OR2X1_LOC_462/B OR2X1_LOC_66/A 0.02fF
C30463 OR2X1_LOC_121/B OR2X1_LOC_121/A 0.14fF
C30464 OR2X1_LOC_147/B OR2X1_LOC_464/A 0.03fF
C30465 AND2X1_LOC_566/B OR2X1_LOC_7/A 0.03fF
C30466 OR2X1_LOC_753/A AND2X1_LOC_614/a_8_24# 0.04fF
C30467 OR2X1_LOC_160/B OR2X1_LOC_643/A 0.08fF
C30468 OR2X1_LOC_647/B OR2X1_LOC_646/B 0.02fF
C30469 OR2X1_LOC_70/Y OR2X1_LOC_595/A 0.24fF
C30470 OR2X1_LOC_502/A AND2X1_LOC_414/a_8_24# 0.05fF
C30471 OR2X1_LOC_160/B OR2X1_LOC_778/Y 0.15fF
C30472 OR2X1_LOC_377/A OR2X1_LOC_459/A 0.14fF
C30473 AND2X1_LOC_191/B OR2X1_LOC_613/Y 1.38fF
C30474 AND2X1_LOC_557/a_36_24# OR2X1_LOC_595/A 0.00fF
C30475 INPUT_0 AND2X1_LOC_139/B 0.11fF
C30476 AND2X1_LOC_514/Y OR2X1_LOC_428/A 0.07fF
C30477 AND2X1_LOC_41/A OR2X1_LOC_541/a_8_216# 0.06fF
C30478 OR2X1_LOC_45/B OR2X1_LOC_19/B 0.10fF
C30479 OR2X1_LOC_600/A OR2X1_LOC_106/A 0.04fF
C30480 OR2X1_LOC_814/A OR2X1_LOC_362/a_8_216# 0.01fF
C30481 AND2X1_LOC_345/Y OR2X1_LOC_382/a_8_216# -0.00fF
C30482 OR2X1_LOC_352/A AND2X1_LOC_12/Y 0.07fF
C30483 OR2X1_LOC_100/Y OR2X1_LOC_656/B 0.00fF
C30484 AND2X1_LOC_95/Y OR2X1_LOC_502/A 0.24fF
C30485 INPUT_5 OR2X1_LOC_1/a_8_216# 0.01fF
C30486 OR2X1_LOC_851/a_8_216# OR2X1_LOC_155/A 0.47fF
C30487 OR2X1_LOC_46/A AND2X1_LOC_44/Y 0.37fF
C30488 OR2X1_LOC_633/Y OR2X1_LOC_502/A 0.03fF
C30489 OR2X1_LOC_49/A AND2X1_LOC_671/a_8_24# 0.00fF
C30490 OR2X1_LOC_834/a_8_216# OR2X1_LOC_375/A 0.01fF
C30491 OR2X1_LOC_695/Y OR2X1_LOC_7/A 0.01fF
C30492 AND2X1_LOC_474/A AND2X1_LOC_287/Y 0.00fF
C30493 OR2X1_LOC_51/Y AND2X1_LOC_673/a_8_24# 0.02fF
C30494 OR2X1_LOC_49/A OR2X1_LOC_606/Y 0.02fF
C30495 OR2X1_LOC_840/A AND2X1_LOC_601/a_8_24# 0.13fF
C30496 OR2X1_LOC_92/Y AND2X1_LOC_454/Y 0.01fF
C30497 OR2X1_LOC_135/Y AND2X1_LOC_537/Y 0.15fF
C30498 OR2X1_LOC_244/A OR2X1_LOC_572/a_8_216# 0.03fF
C30499 OR2X1_LOC_692/Y OR2X1_LOC_46/A 0.03fF
C30500 AND2X1_LOC_22/Y AND2X1_LOC_53/Y 0.21fF
C30501 VDD AND2X1_LOC_155/Y 0.01fF
C30502 AND2X1_LOC_309/a_8_24# AND2X1_LOC_603/a_8_24# 0.23fF
C30503 OR2X1_LOC_158/A OR2X1_LOC_295/a_8_216# 0.01fF
C30504 OR2X1_LOC_446/B OR2X1_LOC_513/Y 0.03fF
C30505 OR2X1_LOC_23/a_8_216# OR2X1_LOC_39/A 0.02fF
C30506 AND2X1_LOC_367/B OR2X1_LOC_485/A 0.01fF
C30507 OR2X1_LOC_51/Y OR2X1_LOC_74/A 0.37fF
C30508 AND2X1_LOC_713/Y OR2X1_LOC_64/Y 0.01fF
C30509 VDD OR2X1_LOC_230/a_8_216# 0.21fF
C30510 OR2X1_LOC_751/Y OR2X1_LOC_44/Y 0.01fF
C30511 VDD OR2X1_LOC_193/A 0.71fF
C30512 OR2X1_LOC_3/Y OR2X1_LOC_12/a_8_216# 0.37fF
C30513 AND2X1_LOC_58/a_8_24# OR2X1_LOC_87/A 0.11fF
C30514 OR2X1_LOC_61/B OR2X1_LOC_358/B 0.00fF
C30515 OR2X1_LOC_599/A OR2X1_LOC_92/Y 0.07fF
C30516 OR2X1_LOC_427/A AND2X1_LOC_466/a_8_24# 0.01fF
C30517 OR2X1_LOC_154/A OR2X1_LOC_653/Y 0.16fF
C30518 AND2X1_LOC_508/A AND2X1_LOC_474/Y 0.02fF
C30519 OR2X1_LOC_45/B OR2X1_LOC_75/Y 0.50fF
C30520 AND2X1_LOC_586/a_8_24# OR2X1_LOC_130/A 0.11fF
C30521 AND2X1_LOC_22/Y OR2X1_LOC_223/A 0.03fF
C30522 OR2X1_LOC_485/A AND2X1_LOC_508/A 0.09fF
C30523 OR2X1_LOC_308/a_36_216# OR2X1_LOC_269/B 0.00fF
C30524 OR2X1_LOC_36/Y OR2X1_LOC_427/A 0.47fF
C30525 OR2X1_LOC_648/A AND2X1_LOC_51/Y 0.29fF
C30526 OR2X1_LOC_160/A OR2X1_LOC_128/a_36_216# 0.01fF
C30527 OR2X1_LOC_167/a_8_216# OR2X1_LOC_95/Y 0.01fF
C30528 AND2X1_LOC_303/A OR2X1_LOC_18/Y 4.38fF
C30529 OR2X1_LOC_405/A OR2X1_LOC_653/A 0.59fF
C30530 OR2X1_LOC_467/B OR2X1_LOC_477/a_8_216# 0.49fF
C30531 OR2X1_LOC_341/Y OR2X1_LOC_350/a_8_216# 0.39fF
C30532 OR2X1_LOC_235/a_36_216# OR2X1_LOC_278/Y 0.00fF
C30533 OR2X1_LOC_527/Y AND2X1_LOC_663/A 0.10fF
C30534 OR2X1_LOC_600/A OR2X1_LOC_46/A 3.25fF
C30535 GATE_366 OR2X1_LOC_625/Y 0.02fF
C30536 OR2X1_LOC_459/B OR2X1_LOC_463/B 0.01fF
C30537 AND2X1_LOC_174/a_8_24# OR2X1_LOC_6/A 0.01fF
C30538 AND2X1_LOC_40/Y OR2X1_LOC_654/A 0.03fF
C30539 VDD AND2X1_LOC_633/Y 0.41fF
C30540 OR2X1_LOC_241/a_8_216# OR2X1_LOC_375/A 0.01fF
C30541 AND2X1_LOC_326/B AND2X1_LOC_326/a_8_24# 0.11fF
C30542 OR2X1_LOC_160/B OR2X1_LOC_113/A 0.01fF
C30543 OR2X1_LOC_814/A OR2X1_LOC_776/Y 0.10fF
C30544 OR2X1_LOC_364/A AND2X1_LOC_43/B 0.07fF
C30545 AND2X1_LOC_568/B AND2X1_LOC_477/A 0.19fF
C30546 AND2X1_LOC_577/Y AND2X1_LOC_578/a_36_24# 0.01fF
C30547 AND2X1_LOC_64/Y OR2X1_LOC_318/B 0.03fF
C30548 OR2X1_LOC_185/Y AND2X1_LOC_43/B 0.45fF
C30549 OR2X1_LOC_812/A OR2X1_LOC_269/B 0.01fF
C30550 AND2X1_LOC_95/Y OR2X1_LOC_137/Y 0.00fF
C30551 AND2X1_LOC_817/B OR2X1_LOC_848/A 0.16fF
C30552 VDD D_INPUT_0 0.94fF
C30553 OR2X1_LOC_440/A OR2X1_LOC_180/a_8_216# 0.02fF
C30554 OR2X1_LOC_363/B OR2X1_LOC_814/A 0.01fF
C30555 OR2X1_LOC_348/Y OR2X1_LOC_286/B 0.03fF
C30556 OR2X1_LOC_77/a_8_216# OR2X1_LOC_56/A 0.01fF
C30557 OR2X1_LOC_489/A D_INPUT_1 0.04fF
C30558 OR2X1_LOC_40/Y AND2X1_LOC_675/A 0.09fF
C30559 OR2X1_LOC_158/A AND2X1_LOC_472/a_36_24# 0.01fF
C30560 AND2X1_LOC_682/a_8_24# AND2X1_LOC_3/Y 0.02fF
C30561 AND2X1_LOC_574/A AND2X1_LOC_663/A 0.50fF
C30562 OR2X1_LOC_485/A OR2X1_LOC_48/B 0.09fF
C30563 AND2X1_LOC_64/Y OR2X1_LOC_854/A 0.03fF
C30564 AND2X1_LOC_326/A AND2X1_LOC_857/Y 0.05fF
C30565 OR2X1_LOC_630/Y OR2X1_LOC_62/B 0.15fF
C30566 AND2X1_LOC_838/Y AND2X1_LOC_838/a_8_24# 0.00fF
C30567 AND2X1_LOC_196/Y OR2X1_LOC_56/A 0.01fF
C30568 AND2X1_LOC_575/Y AND2X1_LOC_576/Y 0.27fF
C30569 OR2X1_LOC_600/A AND2X1_LOC_227/Y 0.03fF
C30570 OR2X1_LOC_87/A OR2X1_LOC_203/Y 0.07fF
C30571 OR2X1_LOC_271/a_8_216# OR2X1_LOC_36/Y 0.01fF
C30572 OR2X1_LOC_485/A OR2X1_LOC_18/Y 0.82fF
C30573 AND2X1_LOC_123/a_8_24# AND2X1_LOC_123/Y 0.01fF
C30574 OR2X1_LOC_768/A OR2X1_LOC_720/B 0.01fF
C30575 OR2X1_LOC_43/A AND2X1_LOC_319/A 0.02fF
C30576 OR2X1_LOC_96/Y D_INPUT_3 0.99fF
C30577 OR2X1_LOC_490/a_8_216# OR2X1_LOC_67/Y 0.01fF
C30578 VDD AND2X1_LOC_450/Y 0.25fF
C30579 AND2X1_LOC_695/a_8_24# AND2X1_LOC_3/Y 0.02fF
C30580 OR2X1_LOC_404/Y OR2X1_LOC_575/A 0.03fF
C30581 OR2X1_LOC_827/Y AND2X1_LOC_838/Y 0.23fF
C30582 OR2X1_LOC_175/Y OR2X1_LOC_566/a_8_216# 0.08fF
C30583 OR2X1_LOC_756/B OR2X1_LOC_814/A 2.44fF
C30584 OR2X1_LOC_373/Y OR2X1_LOC_406/A 0.03fF
C30585 OR2X1_LOC_70/A OR2X1_LOC_428/A 0.03fF
C30586 AND2X1_LOC_650/Y AND2X1_LOC_654/a_8_24# 0.07fF
C30587 OR2X1_LOC_502/A OR2X1_LOC_415/a_8_216# 0.05fF
C30588 OR2X1_LOC_481/Y AND2X1_LOC_847/Y 0.02fF
C30589 OR2X1_LOC_272/a_8_216# AND2X1_LOC_139/B 0.02fF
C30590 OR2X1_LOC_625/a_8_216# OR2X1_LOC_64/Y 0.01fF
C30591 OR2X1_LOC_772/A D_INPUT_1 0.03fF
C30592 AND2X1_LOC_697/a_8_24# OR2X1_LOC_375/A 0.01fF
C30593 AND2X1_LOC_7/B AND2X1_LOC_751/a_8_24# 0.04fF
C30594 AND2X1_LOC_56/B OR2X1_LOC_564/A 0.32fF
C30595 OR2X1_LOC_510/Y AND2X1_LOC_42/B 0.09fF
C30596 INPUT_0 AND2X1_LOC_47/Y 0.06fF
C30597 OR2X1_LOC_680/A OR2X1_LOC_74/A 0.10fF
C30598 OR2X1_LOC_6/A OR2X1_LOC_24/Y 0.06fF
C30599 AND2X1_LOC_59/Y OR2X1_LOC_602/a_8_216# 0.03fF
C30600 AND2X1_LOC_53/Y OR2X1_LOC_706/A 0.09fF
C30601 AND2X1_LOC_524/a_8_24# OR2X1_LOC_551/B 0.03fF
C30602 OR2X1_LOC_121/B OR2X1_LOC_784/Y 0.52fF
C30603 OR2X1_LOC_589/A AND2X1_LOC_644/a_36_24# 0.01fF
C30604 AND2X1_LOC_208/B D_INPUT_0 0.02fF
C30605 OR2X1_LOC_161/B AND2X1_LOC_430/B 0.00fF
C30606 AND2X1_LOC_560/B OR2X1_LOC_529/Y 0.01fF
C30607 AND2X1_LOC_44/Y OR2X1_LOC_513/a_36_216# 0.00fF
C30608 OR2X1_LOC_161/B OR2X1_LOC_779/B 0.20fF
C30609 AND2X1_LOC_456/B AND2X1_LOC_859/B 0.00fF
C30610 OR2X1_LOC_64/Y AND2X1_LOC_436/B 0.02fF
C30611 OR2X1_LOC_417/Y AND2X1_LOC_449/Y 0.09fF
C30612 AND2X1_LOC_95/Y AND2X1_LOC_48/A 0.10fF
C30613 INPUT_5 OR2X1_LOC_31/Y 0.42fF
C30614 OR2X1_LOC_68/B OR2X1_LOC_843/B 0.06fF
C30615 OR2X1_LOC_619/Y OR2X1_LOC_46/A 0.10fF
C30616 OR2X1_LOC_306/Y AND2X1_LOC_307/Y 0.00fF
C30617 AND2X1_LOC_12/Y OR2X1_LOC_34/B 0.03fF
C30618 AND2X1_LOC_47/Y OR2X1_LOC_775/a_8_216# 0.03fF
C30619 OR2X1_LOC_160/A OR2X1_LOC_19/B 0.10fF
C30620 OR2X1_LOC_600/A OR2X1_LOC_41/Y 0.46fF
C30621 OR2X1_LOC_493/B OR2X1_LOC_493/Y 0.79fF
C30622 OR2X1_LOC_810/A AND2X1_LOC_42/B 0.05fF
C30623 OR2X1_LOC_472/B AND2X1_LOC_43/B 0.07fF
C30624 OR2X1_LOC_68/B OR2X1_LOC_549/A 0.09fF
C30625 OR2X1_LOC_479/Y OR2X1_LOC_711/A 0.03fF
C30626 AND2X1_LOC_866/A OR2X1_LOC_92/Y 0.03fF
C30627 AND2X1_LOC_408/a_8_24# AND2X1_LOC_409/B 0.00fF
C30628 AND2X1_LOC_99/A AND2X1_LOC_845/Y 0.18fF
C30629 OR2X1_LOC_71/A OR2X1_LOC_548/B 0.01fF
C30630 OR2X1_LOC_859/a_8_216# D_INPUT_1 0.01fF
C30631 OR2X1_LOC_316/Y INPUT_1 0.02fF
C30632 INPUT_5 OR2X1_LOC_587/a_36_216# 0.00fF
C30633 OR2X1_LOC_519/Y OR2X1_LOC_417/A 0.01fF
C30634 AND2X1_LOC_519/a_36_24# OR2X1_LOC_375/A 0.01fF
C30635 OR2X1_LOC_263/a_8_216# OR2X1_LOC_85/A 0.14fF
C30636 OR2X1_LOC_369/a_36_216# AND2X1_LOC_222/Y 0.00fF
C30637 OR2X1_LOC_140/A OR2X1_LOC_560/A 0.14fF
C30638 OR2X1_LOC_682/a_8_216# AND2X1_LOC_687/A 0.47fF
C30639 OR2X1_LOC_507/A OR2X1_LOC_560/A 0.04fF
C30640 OR2X1_LOC_799/A OR2X1_LOC_436/Y 0.03fF
C30641 INPUT_0 OR2X1_LOC_598/A 0.11fF
C30642 OR2X1_LOC_78/A OR2X1_LOC_675/Y 0.02fF
C30643 OR2X1_LOC_852/A AND2X1_LOC_43/B 0.16fF
C30644 OR2X1_LOC_128/a_8_216# AND2X1_LOC_47/Y 0.01fF
C30645 AND2X1_LOC_139/B OR2X1_LOC_417/A 0.02fF
C30646 OR2X1_LOC_529/Y OR2X1_LOC_64/Y 0.03fF
C30647 AND2X1_LOC_102/a_8_24# OR2X1_LOC_54/Y 0.04fF
C30648 AND2X1_LOC_645/a_36_24# OR2X1_LOC_48/B 0.01fF
C30649 OR2X1_LOC_795/a_8_216# OR2X1_LOC_785/B 0.14fF
C30650 OR2X1_LOC_166/Y OR2X1_LOC_331/Y 0.18fF
C30651 OR2X1_LOC_255/a_8_216# OR2X1_LOC_248/Y 0.04fF
C30652 AND2X1_LOC_401/a_8_24# OR2X1_LOC_396/Y 0.05fF
C30653 AND2X1_LOC_7/B OR2X1_LOC_714/a_8_216# 0.01fF
C30654 OR2X1_LOC_643/A OR2X1_LOC_244/A 0.07fF
C30655 AND2X1_LOC_514/Y AND2X1_LOC_211/a_8_24# 0.03fF
C30656 OR2X1_LOC_244/A OR2X1_LOC_124/Y 0.01fF
C30657 OR2X1_LOC_464/A OR2X1_LOC_318/B 0.03fF
C30658 AND2X1_LOC_474/A AND2X1_LOC_562/Y 0.03fF
C30659 AND2X1_LOC_40/Y OR2X1_LOC_192/B 0.04fF
C30660 OR2X1_LOC_390/a_8_216# OR2X1_LOC_390/B 0.13fF
C30661 AND2X1_LOC_104/a_8_24# D_INPUT_1 0.01fF
C30662 OR2X1_LOC_43/A AND2X1_LOC_170/B 0.01fF
C30663 OR2X1_LOC_59/Y AND2X1_LOC_203/a_36_24# 0.00fF
C30664 OR2X1_LOC_175/Y OR2X1_LOC_170/a_8_216# 0.05fF
C30665 OR2X1_LOC_271/B AND2X1_LOC_318/Y 1.01fF
C30666 OR2X1_LOC_427/A OR2X1_LOC_419/Y 0.10fF
C30667 OR2X1_LOC_311/Y OR2X1_LOC_829/Y 0.02fF
C30668 OR2X1_LOC_529/Y OR2X1_LOC_417/A 0.03fF
C30669 OR2X1_LOC_128/A AND2X1_LOC_72/B 0.01fF
C30670 OR2X1_LOC_22/Y OR2X1_LOC_615/a_8_216# 0.02fF
C30671 OR2X1_LOC_825/a_8_216# INPUT_1 0.01fF
C30672 OR2X1_LOC_45/B OR2X1_LOC_323/A 0.01fF
C30673 AND2X1_LOC_539/a_8_24# AND2X1_LOC_729/B 0.07fF
C30674 OR2X1_LOC_22/Y OR2X1_LOC_275/a_8_216# 0.05fF
C30675 OR2X1_LOC_2/Y OR2X1_LOC_11/a_8_216# 0.02fF
C30676 VDD OR2X1_LOC_339/A 0.08fF
C30677 OR2X1_LOC_696/A OR2X1_LOC_829/A 0.35fF
C30678 OR2X1_LOC_566/A OR2X1_LOC_336/a_8_216# 0.01fF
C30679 OR2X1_LOC_121/Y AND2X1_LOC_64/Y 0.07fF
C30680 AND2X1_LOC_3/Y OR2X1_LOC_227/Y 0.02fF
C30681 OR2X1_LOC_43/A AND2X1_LOC_721/A 0.11fF
C30682 OR2X1_LOC_427/A OR2X1_LOC_152/A 0.03fF
C30683 AND2X1_LOC_3/Y OR2X1_LOC_284/B 0.01fF
C30684 OR2X1_LOC_227/a_8_216# OR2X1_LOC_814/A 0.01fF
C30685 OR2X1_LOC_665/Y AND2X1_LOC_620/Y 3.56fF
C30686 AND2X1_LOC_3/Y D_INPUT_1 0.06fF
C30687 OR2X1_LOC_647/B D_INPUT_1 0.07fF
C30688 AND2X1_LOC_369/a_8_24# OR2X1_LOC_318/B 0.00fF
C30689 AND2X1_LOC_76/Y OR2X1_LOC_521/a_8_216# 0.01fF
C30690 AND2X1_LOC_43/B OR2X1_LOC_568/A 0.07fF
C30691 OR2X1_LOC_690/A OR2X1_LOC_598/A 0.31fF
C30692 AND2X1_LOC_564/B AND2X1_LOC_476/Y 0.04fF
C30693 OR2X1_LOC_139/A AND2X1_LOC_65/A 0.28fF
C30694 AND2X1_LOC_699/a_8_24# OR2X1_LOC_155/A 0.01fF
C30695 OR2X1_LOC_574/A OR2X1_LOC_493/Y 0.05fF
C30696 D_INPUT_5 OR2X1_LOC_376/Y 0.01fF
C30697 AND2X1_LOC_64/Y OR2X1_LOC_114/B 0.06fF
C30698 AND2X1_LOC_555/Y AND2X1_LOC_860/A 0.00fF
C30699 OR2X1_LOC_502/A OR2X1_LOC_788/B 0.03fF
C30700 OR2X1_LOC_198/a_8_216# AND2X1_LOC_70/Y 0.01fF
C30701 OR2X1_LOC_40/Y AND2X1_LOC_241/a_8_24# 0.01fF
C30702 AND2X1_LOC_56/B OR2X1_LOC_228/Y 0.03fF
C30703 OR2X1_LOC_502/A AND2X1_LOC_41/Y 0.01fF
C30704 OR2X1_LOC_600/A OR2X1_LOC_748/a_8_216# 0.01fF
C30705 OR2X1_LOC_368/Y AND2X1_LOC_476/Y 0.03fF
C30706 OR2X1_LOC_364/B OR2X1_LOC_161/B 0.00fF
C30707 OR2X1_LOC_709/A OR2X1_LOC_161/B 0.07fF
C30708 OR2X1_LOC_43/A OR2X1_LOC_331/Y 0.33fF
C30709 AND2X1_LOC_91/B OR2X1_LOC_160/B 0.64fF
C30710 OR2X1_LOC_294/Y AND2X1_LOC_279/a_8_24# 0.01fF
C30711 OR2X1_LOC_6/B AND2X1_LOC_7/B 0.65fF
C30712 AND2X1_LOC_539/Y VDD 0.22fF
C30713 AND2X1_LOC_679/a_36_24# OR2X1_LOC_155/A 0.01fF
C30714 OR2X1_LOC_739/A OR2X1_LOC_317/B 0.00fF
C30715 OR2X1_LOC_542/B OR2X1_LOC_562/A 0.03fF
C30716 OR2X1_LOC_807/a_8_216# OR2X1_LOC_675/Y 0.02fF
C30717 AND2X1_LOC_724/a_8_24# OR2X1_LOC_604/A 0.01fF
C30718 OR2X1_LOC_786/a_8_216# AND2X1_LOC_44/Y 0.06fF
C30719 OR2X1_LOC_625/Y OR2X1_LOC_13/B 0.13fF
C30720 OR2X1_LOC_680/a_8_216# VDD 0.21fF
C30721 AND2X1_LOC_714/B OR2X1_LOC_12/Y 0.01fF
C30722 OR2X1_LOC_161/A OR2X1_LOC_501/a_36_216# 0.00fF
C30723 OR2X1_LOC_416/a_8_216# INPUT_1 0.01fF
C30724 AND2X1_LOC_223/A AND2X1_LOC_223/a_8_24# 0.01fF
C30725 OR2X1_LOC_780/B OR2X1_LOC_780/a_8_216# 0.02fF
C30726 OR2X1_LOC_739/A OR2X1_LOC_728/a_36_216# 0.00fF
C30727 AND2X1_LOC_60/a_8_24# AND2X1_LOC_18/Y 0.01fF
C30728 OR2X1_LOC_68/a_36_216# OR2X1_LOC_68/B 0.03fF
C30729 OR2X1_LOC_161/A OR2X1_LOC_112/A 0.01fF
C30730 AND2X1_LOC_31/Y OR2X1_LOC_733/B 0.26fF
C30731 OR2X1_LOC_56/A OR2X1_LOC_321/a_8_216# 0.01fF
C30732 AND2X1_LOC_64/Y OR2X1_LOC_538/A 0.03fF
C30733 OR2X1_LOC_405/A OR2X1_LOC_723/B 0.08fF
C30734 AND2X1_LOC_801/B OR2X1_LOC_760/Y 0.81fF
C30735 OR2X1_LOC_158/A OR2X1_LOC_421/Y 1.04fF
C30736 OR2X1_LOC_49/A OR2X1_LOC_622/A 0.05fF
C30737 OR2X1_LOC_696/A D_INPUT_5 0.25fF
C30738 AND2X1_LOC_181/Y AND2X1_LOC_182/a_8_24# 0.11fF
C30739 AND2X1_LOC_350/B VDD 0.19fF
C30740 AND2X1_LOC_462/Y AND2X1_LOC_476/A 0.04fF
C30741 AND2X1_LOC_12/Y OR2X1_LOC_590/Y 0.01fF
C30742 OR2X1_LOC_78/A OR2X1_LOC_779/A 0.01fF
C30743 AND2X1_LOC_633/Y OR2X1_LOC_67/Y 0.20fF
C30744 AND2X1_LOC_2/Y AND2X1_LOC_44/Y 0.03fF
C30745 OR2X1_LOC_244/Y OR2X1_LOC_342/A 0.02fF
C30746 OR2X1_LOC_269/B OR2X1_LOC_317/B 0.35fF
C30747 OR2X1_LOC_447/A OR2X1_LOC_308/Y 0.05fF
C30748 OR2X1_LOC_607/a_8_216# D_INPUT_1 0.06fF
C30749 AND2X1_LOC_70/Y OR2X1_LOC_161/B 1.51fF
C30750 AND2X1_LOC_566/B AND2X1_LOC_353/a_8_24# 0.10fF
C30751 AND2X1_LOC_40/Y OR2X1_LOC_502/Y 0.31fF
C30752 AND2X1_LOC_544/Y OR2X1_LOC_441/Y 0.03fF
C30753 AND2X1_LOC_674/a_8_24# AND2X1_LOC_31/Y 0.01fF
C30754 AND2X1_LOC_83/a_8_24# OR2X1_LOC_66/A 0.08fF
C30755 D_INPUT_0 OR2X1_LOC_67/Y 0.08fF
C30756 VDD AND2X1_LOC_771/B 0.14fF
C30757 OR2X1_LOC_794/A OR2X1_LOC_605/Y -0.00fF
C30758 OR2X1_LOC_269/B OR2X1_LOC_580/A 0.06fF
C30759 OR2X1_LOC_680/a_8_216# OR2X1_LOC_677/Y 0.01fF
C30760 OR2X1_LOC_1/a_36_216# INPUT_6 0.03fF
C30761 OR2X1_LOC_744/A AND2X1_LOC_802/Y 0.16fF
C30762 AND2X1_LOC_81/B AND2X1_LOC_239/a_8_24# 0.01fF
C30763 VDD OR2X1_LOC_131/A 0.44fF
C30764 AND2X1_LOC_41/A OR2X1_LOC_576/A 0.03fF
C30765 OR2X1_LOC_287/B OR2X1_LOC_579/a_36_216# 0.00fF
C30766 VDD OR2X1_LOC_515/A -0.00fF
C30767 OR2X1_LOC_862/a_36_216# OR2X1_LOC_862/A 0.01fF
C30768 OR2X1_LOC_736/Y OR2X1_LOC_78/A 0.03fF
C30769 VDD OR2X1_LOC_598/Y 0.12fF
C30770 OR2X1_LOC_858/a_36_216# OR2X1_LOC_362/A 0.00fF
C30771 AND2X1_LOC_443/a_8_24# OR2X1_LOC_56/A 0.04fF
C30772 AND2X1_LOC_736/Y OR2X1_LOC_406/Y 0.05fF
C30773 OR2X1_LOC_31/Y AND2X1_LOC_204/Y 0.02fF
C30774 OR2X1_LOC_826/Y AND2X1_LOC_837/a_8_24# 0.23fF
C30775 OR2X1_LOC_600/A INPUT_2 0.10fF
C30776 OR2X1_LOC_614/Y OR2X1_LOC_78/A 0.74fF
C30777 OR2X1_LOC_703/A OR2X1_LOC_161/B 0.03fF
C30778 AND2X1_LOC_22/Y OR2X1_LOC_502/A 0.33fF
C30779 OR2X1_LOC_106/Y AND2X1_LOC_76/Y 0.00fF
C30780 OR2X1_LOC_141/B OR2X1_LOC_141/a_8_216# 0.02fF
C30781 OR2X1_LOC_31/Y AND2X1_LOC_228/a_8_24# 0.00fF
C30782 AND2X1_LOC_431/a_8_24# OR2X1_LOC_358/A 0.01fF
C30783 OR2X1_LOC_100/a_8_216# AND2X1_LOC_64/Y 0.01fF
C30784 OR2X1_LOC_51/Y AND2X1_LOC_254/a_8_24# 0.00fF
C30785 OR2X1_LOC_696/A AND2X1_LOC_838/Y 0.02fF
C30786 OR2X1_LOC_449/B AND2X1_LOC_36/Y 0.04fF
C30787 AND2X1_LOC_794/B AND2X1_LOC_471/Y 0.01fF
C30788 AND2X1_LOC_539/Y OR2X1_LOC_829/a_8_216# 0.01fF
C30789 GATE_366 OR2X1_LOC_759/Y 0.01fF
C30790 INPUT_1 OR2X1_LOC_153/a_8_216# 0.18fF
C30791 AND2X1_LOC_12/Y AND2X1_LOC_64/Y 6.59fF
C30792 OR2X1_LOC_686/a_8_216# OR2X1_LOC_687/A -0.00fF
C30793 VDD AND2X1_LOC_326/B 0.21fF
C30794 OR2X1_LOC_786/Y OR2X1_LOC_795/a_8_216# 0.02fF
C30795 OR2X1_LOC_51/Y AND2X1_LOC_860/A 0.03fF
C30796 OR2X1_LOC_49/A AND2X1_LOC_404/A 0.01fF
C30797 OR2X1_LOC_528/Y OR2X1_LOC_59/Y 0.02fF
C30798 OR2X1_LOC_809/B AND2X1_LOC_110/Y 0.02fF
C30799 OR2X1_LOC_149/B OR2X1_LOC_161/A 0.00fF
C30800 OR2X1_LOC_357/a_8_216# AND2X1_LOC_40/Y 0.01fF
C30801 OR2X1_LOC_51/Y OR2X1_LOC_626/Y 0.00fF
C30802 OR2X1_LOC_106/Y OR2X1_LOC_67/A 0.01fF
C30803 AND2X1_LOC_326/A OR2X1_LOC_437/A 0.00fF
C30804 D_INPUT_1 AND2X1_LOC_225/a_8_24# 0.03fF
C30805 OR2X1_LOC_76/A OR2X1_LOC_303/B 0.28fF
C30806 OR2X1_LOC_404/Y OR2X1_LOC_735/B 0.14fF
C30807 OR2X1_LOC_54/Y OR2X1_LOC_71/A 0.47fF
C30808 OR2X1_LOC_348/Y OR2X1_LOC_363/A 0.01fF
C30809 AND2X1_LOC_150/a_8_24# OR2X1_LOC_474/Y 0.03fF
C30810 VDD OR2X1_LOC_795/B -0.00fF
C30811 OR2X1_LOC_446/Y AND2X1_LOC_427/a_8_24# 0.24fF
C30812 AND2X1_LOC_51/Y OR2X1_LOC_730/B 0.10fF
C30813 OR2X1_LOC_756/B OR2X1_LOC_410/Y 0.11fF
C30814 AND2X1_LOC_12/Y AND2X1_LOC_599/a_8_24# 0.01fF
C30815 OR2X1_LOC_352/A OR2X1_LOC_182/B 0.96fF
C30816 VDD OR2X1_LOC_612/Y 0.12fF
C30817 AND2X1_LOC_511/a_8_24# OR2X1_LOC_623/B 0.21fF
C30818 OR2X1_LOC_739/A AND2X1_LOC_44/Y 0.05fF
C30819 VDD AND2X1_LOC_471/Y 0.10fF
C30820 AND2X1_LOC_95/Y OR2X1_LOC_34/a_8_216# 0.01fF
C30821 AND2X1_LOC_162/a_8_24# OR2X1_LOC_51/Y 0.01fF
C30822 AND2X1_LOC_781/Y AND2X1_LOC_782/a_8_24# 0.00fF
C30823 OR2X1_LOC_335/Y VDD 0.31fF
C30824 AND2X1_LOC_807/Y OR2X1_LOC_816/A 0.03fF
C30825 OR2X1_LOC_17/Y INPUT_6 0.03fF
C30826 AND2X1_LOC_561/a_8_24# AND2X1_LOC_489/Y 0.02fF
C30827 OR2X1_LOC_177/Y OR2X1_LOC_427/A 0.14fF
C30828 AND2X1_LOC_40/Y AND2X1_LOC_265/a_8_24# 0.03fF
C30829 AND2X1_LOC_722/A OR2X1_LOC_600/A 0.03fF
C30830 OR2X1_LOC_40/Y OR2X1_LOC_92/Y 0.21fF
C30831 OR2X1_LOC_158/A OR2X1_LOC_278/Y 0.03fF
C30832 OR2X1_LOC_756/B OR2X1_LOC_244/Y 0.02fF
C30833 AND2X1_LOC_70/Y OR2X1_LOC_435/B 0.01fF
C30834 OR2X1_LOC_524/Y AND2X1_LOC_469/B 0.18fF
C30835 OR2X1_LOC_97/A OR2X1_LOC_358/B 0.02fF
C30836 AND2X1_LOC_12/Y AND2X1_LOC_82/Y 0.00fF
C30837 OR2X1_LOC_791/A VDD 0.04fF
C30838 OR2X1_LOC_6/A AND2X1_LOC_208/Y 0.02fF
C30839 OR2X1_LOC_471/Y OR2X1_LOC_550/B 6.13fF
C30840 AND2X1_LOC_576/Y AND2X1_LOC_242/a_8_24# 0.01fF
C30841 OR2X1_LOC_158/A AND2X1_LOC_662/B 0.04fF
C30842 OR2X1_LOC_308/a_8_216# OR2X1_LOC_160/B 0.03fF
C30843 AND2X1_LOC_40/Y VDD 2.84fF
C30844 AND2X1_LOC_456/B OR2X1_LOC_56/A 0.03fF
C30845 OR2X1_LOC_121/B AND2X1_LOC_36/Y 0.11fF
C30846 AND2X1_LOC_64/Y AND2X1_LOC_79/Y 4.54fF
C30847 AND2X1_LOC_512/Y OR2X1_LOC_59/Y 0.08fF
C30848 OR2X1_LOC_678/a_8_216# OR2X1_LOC_678/Y 0.01fF
C30849 OR2X1_LOC_684/a_36_216# OR2X1_LOC_426/A 0.00fF
C30850 OR2X1_LOC_436/Y OR2X1_LOC_446/B 0.01fF
C30851 OR2X1_LOC_106/Y AND2X1_LOC_489/Y 0.21fF
C30852 AND2X1_LOC_363/B AND2X1_LOC_363/Y 0.03fF
C30853 AND2X1_LOC_95/Y OR2X1_LOC_542/a_8_216# 0.02fF
C30854 OR2X1_LOC_604/A OR2X1_LOC_427/A 0.78fF
C30855 AND2X1_LOC_191/Y AND2X1_LOC_213/a_8_24# 0.05fF
C30856 AND2X1_LOC_22/Y OR2X1_LOC_137/Y -0.02fF
C30857 AND2X1_LOC_719/Y AND2X1_LOC_573/A 0.10fF
C30858 AND2X1_LOC_57/Y AND2X1_LOC_51/Y 0.09fF
C30859 INPUT_0 AND2X1_LOC_529/a_36_24# 0.00fF
C30860 OR2X1_LOC_808/B OR2X1_LOC_78/A 0.02fF
C30861 AND2X1_LOC_354/a_36_24# AND2X1_LOC_810/B 0.01fF
C30862 OR2X1_LOC_149/B AND2X1_LOC_525/a_8_24# 0.29fF
C30863 OR2X1_LOC_269/B AND2X1_LOC_44/Y 1.41fF
C30864 VDD AND2X1_LOC_840/A 0.11fF
C30865 VDD OR2X1_LOC_810/a_8_216# 0.00fF
C30866 AND2X1_LOC_155/a_8_24# OR2X1_LOC_51/Y 0.06fF
C30867 OR2X1_LOC_600/A OR2X1_LOC_250/a_8_216# 0.01fF
C30868 VDD AND2X1_LOC_375/a_8_24# -0.00fF
C30869 OR2X1_LOC_287/B OR2X1_LOC_366/B 0.01fF
C30870 AND2X1_LOC_70/Y OR2X1_LOC_61/Y 0.75fF
C30871 INPUT_0 OR2X1_LOC_828/a_8_216# 0.03fF
C30872 OR2X1_LOC_52/B AND2X1_LOC_219/A 0.07fF
C30873 OR2X1_LOC_326/a_8_216# OR2X1_LOC_502/A 0.01fF
C30874 OR2X1_LOC_40/Y OR2X1_LOC_65/B 0.09fF
C30875 OR2X1_LOC_160/A AND2X1_LOC_110/Y 0.03fF
C30876 OR2X1_LOC_599/A AND2X1_LOC_729/a_8_24# 0.00fF
C30877 OR2X1_LOC_377/A OR2X1_LOC_389/A 0.03fF
C30878 AND2X1_LOC_47/Y OR2X1_LOC_195/a_36_216# 0.00fF
C30879 AND2X1_LOC_70/Y AND2X1_LOC_536/a_8_24# 0.01fF
C30880 OR2X1_LOC_508/A AND2X1_LOC_41/A 0.01fF
C30881 OR2X1_LOC_149/B AND2X1_LOC_51/Y 0.03fF
C30882 OR2X1_LOC_589/A AND2X1_LOC_361/A 0.01fF
C30883 OR2X1_LOC_181/B AND2X1_LOC_179/a_8_24# 0.02fF
C30884 AND2X1_LOC_848/Y AND2X1_LOC_244/a_36_24# 0.00fF
C30885 OR2X1_LOC_744/A AND2X1_LOC_832/a_36_24# 0.00fF
C30886 OR2X1_LOC_158/A AND2X1_LOC_472/B 0.08fF
C30887 OR2X1_LOC_284/a_8_216# OR2X1_LOC_161/A 0.01fF
C30888 AND2X1_LOC_347/B OR2X1_LOC_44/Y 0.02fF
C30889 OR2X1_LOC_769/A OR2X1_LOC_379/Y 0.00fF
C30890 OR2X1_LOC_84/Y OR2X1_LOC_71/A 0.01fF
C30891 OR2X1_LOC_756/B OR2X1_LOC_147/B 0.03fF
C30892 OR2X1_LOC_680/A OR2X1_LOC_626/Y 0.03fF
C30893 OR2X1_LOC_165/Y AND2X1_LOC_168/a_8_24# 0.01fF
C30894 VDD OR2X1_LOC_87/Y 0.29fF
C30895 OR2X1_LOC_269/B OR2X1_LOC_719/a_8_216# 0.01fF
C30896 AND2X1_LOC_486/Y OR2X1_LOC_164/Y 0.03fF
C30897 OR2X1_LOC_3/Y AND2X1_LOC_249/a_8_24# 0.01fF
C30898 AND2X1_LOC_555/a_36_24# OR2X1_LOC_748/A 0.00fF
C30899 VDD OR2X1_LOC_848/A 0.27fF
C30900 AND2X1_LOC_98/Y OR2X1_LOC_278/Y 0.04fF
C30901 OR2X1_LOC_516/A OR2X1_LOC_59/Y 0.03fF
C30902 AND2X1_LOC_181/Y OR2X1_LOC_485/A 0.14fF
C30903 OR2X1_LOC_637/B OR2X1_LOC_637/a_8_216# 0.07fF
C30904 VDD OR2X1_LOC_859/B 0.06fF
C30905 OR2X1_LOC_158/A AND2X1_LOC_337/B 0.03fF
C30906 OR2X1_LOC_633/Y OR2X1_LOC_633/a_36_216# 0.00fF
C30907 OR2X1_LOC_51/Y AND2X1_LOC_287/Y 0.01fF
C30908 OR2X1_LOC_235/B AND2X1_LOC_132/a_8_24# 0.01fF
C30909 OR2X1_LOC_91/A AND2X1_LOC_655/A 0.10fF
C30910 AND2X1_LOC_535/Y OR2X1_LOC_312/Y 0.03fF
C30911 AND2X1_LOC_732/a_8_24# OR2X1_LOC_36/Y 0.01fF
C30912 OR2X1_LOC_220/a_8_216# OR2X1_LOC_565/A 0.40fF
C30913 OR2X1_LOC_404/Y OR2X1_LOC_161/B 0.00fF
C30914 OR2X1_LOC_668/a_8_216# OR2X1_LOC_721/Y 0.01fF
C30915 OR2X1_LOC_703/B OR2X1_LOC_78/B 0.37fF
C30916 AND2X1_LOC_340/a_36_24# OR2X1_LOC_262/Y 0.00fF
C30917 OR2X1_LOC_58/Y OR2X1_LOC_585/A 0.03fF
C30918 AND2X1_LOC_720/Y OR2X1_LOC_278/Y 0.02fF
C30919 INPUT_3 AND2X1_LOC_819/a_36_24# 0.00fF
C30920 OR2X1_LOC_756/Y OR2X1_LOC_161/A 0.01fF
C30921 AND2X1_LOC_550/A OR2X1_LOC_441/Y 0.03fF
C30922 OR2X1_LOC_552/A OR2X1_LOC_367/B 0.03fF
C30923 OR2X1_LOC_464/B OR2X1_LOC_741/Y 0.01fF
C30924 AND2X1_LOC_860/a_8_24# OR2X1_LOC_39/A 0.01fF
C30925 OR2X1_LOC_528/Y AND2X1_LOC_191/Y 0.03fF
C30926 AND2X1_LOC_392/A AND2X1_LOC_566/a_36_24# 0.01fF
C30927 AND2X1_LOC_22/Y AND2X1_LOC_48/A 1.14fF
C30928 AND2X1_LOC_80/a_36_24# OR2X1_LOC_78/B 0.00fF
C30929 AND2X1_LOC_498/a_8_24# AND2X1_LOC_56/B 0.13fF
C30930 OR2X1_LOC_517/a_36_216# OR2X1_LOC_39/A 0.01fF
C30931 AND2X1_LOC_320/a_8_24# AND2X1_LOC_56/B 0.03fF
C30932 OR2X1_LOC_87/A OR2X1_LOC_78/B 0.70fF
C30933 OR2X1_LOC_158/A OR2X1_LOC_273/Y 0.01fF
C30934 OR2X1_LOC_92/Y AND2X1_LOC_644/Y 0.01fF
C30935 OR2X1_LOC_811/A OR2X1_LOC_733/a_8_216# 0.04fF
C30936 AND2X1_LOC_658/A OR2X1_LOC_52/B 0.06fF
C30937 OR2X1_LOC_528/Y AND2X1_LOC_711/Y 0.03fF
C30938 AND2X1_LOC_12/Y OR2X1_LOC_512/A 0.03fF
C30939 OR2X1_LOC_600/A OR2X1_LOC_258/a_8_216# 0.01fF
C30940 OR2X1_LOC_696/A OR2X1_LOC_224/Y 0.02fF
C30941 OR2X1_LOC_557/A AND2X1_LOC_18/Y 0.00fF
C30942 OR2X1_LOC_528/Y OR2X1_LOC_70/Y 0.02fF
C30943 AND2X1_LOC_52/a_8_24# AND2X1_LOC_43/B 0.04fF
C30944 AND2X1_LOC_663/A AND2X1_LOC_806/A 0.05fF
C30945 OR2X1_LOC_303/B OR2X1_LOC_566/Y 0.01fF
C30946 AND2X1_LOC_727/Y AND2X1_LOC_810/Y 0.09fF
C30947 OR2X1_LOC_708/B OR2X1_LOC_78/A 0.34fF
C30948 OR2X1_LOC_53/Y OR2X1_LOC_31/Y 0.42fF
C30949 OR2X1_LOC_62/B OR2X1_LOC_16/A 0.05fF
C30950 AND2X1_LOC_367/A AND2X1_LOC_359/B 0.19fF
C30951 OR2X1_LOC_8/Y AND2X1_LOC_37/a_8_24# 0.08fF
C30952 AND2X1_LOC_53/a_8_24# AND2X1_LOC_43/B 0.03fF
C30953 OR2X1_LOC_600/A AND2X1_LOC_847/a_8_24# 0.01fF
C30954 AND2X1_LOC_47/Y AND2X1_LOC_7/B 8.39fF
C30955 VDD OR2X1_LOC_221/A 0.06fF
C30956 OR2X1_LOC_631/B AND2X1_LOC_41/A 0.04fF
C30957 AND2X1_LOC_717/B OR2X1_LOC_56/A 4.06fF
C30958 AND2X1_LOC_477/A OR2X1_LOC_12/Y 0.03fF
C30959 AND2X1_LOC_732/a_36_24# OR2X1_LOC_89/A 0.00fF
C30960 VDD OR2X1_LOC_475/Y 0.22fF
C30961 OR2X1_LOC_427/A AND2X1_LOC_467/a_8_24# 0.02fF
C30962 OR2X1_LOC_606/a_8_216# OR2X1_LOC_646/B 0.47fF
C30963 OR2X1_LOC_617/Y OR2X1_LOC_627/Y 0.00fF
C30964 AND2X1_LOC_578/A AND2X1_LOC_657/Y 0.10fF
C30965 OR2X1_LOC_87/A OR2X1_LOC_721/Y 0.02fF
C30966 OR2X1_LOC_668/a_8_216# OR2X1_LOC_375/A 0.04fF
C30967 OR2X1_LOC_757/A OR2X1_LOC_74/A 0.03fF
C30968 OR2X1_LOC_759/A AND2X1_LOC_663/B 0.00fF
C30969 OR2X1_LOC_235/B AND2X1_LOC_240/Y 0.02fF
C30970 OR2X1_LOC_619/Y AND2X1_LOC_454/Y 0.19fF
C30971 OR2X1_LOC_756/B AND2X1_LOC_171/a_8_24# 0.01fF
C30972 OR2X1_LOC_402/Y OR2X1_LOC_404/a_8_216# 0.03fF
C30973 OR2X1_LOC_755/A AND2X1_LOC_658/A 0.03fF
C30974 OR2X1_LOC_808/B OR2X1_LOC_155/A 0.01fF
C30975 OR2X1_LOC_799/A OR2X1_LOC_799/a_8_216# 0.07fF
C30976 OR2X1_LOC_105/a_8_216# OR2X1_LOC_287/B 0.01fF
C30977 OR2X1_LOC_756/B OR2X1_LOC_843/a_8_216# 0.02fF
C30978 OR2X1_LOC_786/Y OR2X1_LOC_392/B 0.01fF
C30979 OR2X1_LOC_604/A AND2X1_LOC_687/B 0.01fF
C30980 OR2X1_LOC_528/Y AND2X1_LOC_657/a_8_24# 0.23fF
C30981 VDD AND2X1_LOC_687/A -0.00fF
C30982 OR2X1_LOC_825/Y OR2X1_LOC_56/A 0.00fF
C30983 OR2X1_LOC_438/Y OR2X1_LOC_89/A 0.03fF
C30984 OR2X1_LOC_97/A OR2X1_LOC_112/B 0.01fF
C30985 OR2X1_LOC_484/a_8_216# OR2X1_LOC_64/Y 0.01fF
C30986 OR2X1_LOC_92/Y OR2X1_LOC_7/A 2.74fF
C30987 OR2X1_LOC_160/A OR2X1_LOC_835/A 0.02fF
C30988 OR2X1_LOC_47/Y OR2X1_LOC_428/A 0.74fF
C30989 AND2X1_LOC_59/Y OR2X1_LOC_520/Y 0.04fF
C30990 OR2X1_LOC_599/A OR2X1_LOC_619/Y 0.03fF
C30991 OR2X1_LOC_686/a_36_216# AND2X1_LOC_425/Y 0.00fF
C30992 AND2X1_LOC_778/a_36_24# OR2X1_LOC_406/A 0.01fF
C30993 OR2X1_LOC_528/Y OR2X1_LOC_504/Y 0.04fF
C30994 OR2X1_LOC_70/Y AND2X1_LOC_512/Y 0.27fF
C30995 OR2X1_LOC_808/B OR2X1_LOC_605/A 0.10fF
C30996 OR2X1_LOC_154/A AND2X1_LOC_272/a_8_24# 0.05fF
C30997 OR2X1_LOC_124/B OR2X1_LOC_814/A 0.00fF
C30998 AND2X1_LOC_593/Y AND2X1_LOC_653/a_8_24# 0.01fF
C30999 AND2X1_LOC_12/Y AND2X1_LOC_369/a_8_24# 0.02fF
C31000 AND2X1_LOC_502/a_8_24# AND2X1_LOC_576/Y 0.02fF
C31001 AND2X1_LOC_706/Y AND2X1_LOC_645/a_8_24# 0.08fF
C31002 OR2X1_LOC_151/A OR2X1_LOC_440/A 0.01fF
C31003 OR2X1_LOC_851/a_8_216# OR2X1_LOC_814/A 0.06fF
C31004 OR2X1_LOC_185/Y OR2X1_LOC_510/Y 0.03fF
C31005 OR2X1_LOC_87/A OR2X1_LOC_375/A 7.45fF
C31006 OR2X1_LOC_26/Y AND2X1_LOC_621/Y 0.03fF
C31007 OR2X1_LOC_47/Y OR2X1_LOC_595/A 0.03fF
C31008 OR2X1_LOC_51/B INPUT_7 0.18fF
C31009 OR2X1_LOC_158/A OR2X1_LOC_75/Y 0.00fF
C31010 OR2X1_LOC_650/Y OR2X1_LOC_520/a_36_216# 0.01fF
C31011 OR2X1_LOC_377/A OR2X1_LOC_403/B 0.02fF
C31012 OR2X1_LOC_822/Y AND2X1_LOC_835/a_8_24# 0.23fF
C31013 AND2X1_LOC_45/a_36_24# OR2X1_LOC_78/B 0.01fF
C31014 AND2X1_LOC_675/Y AND2X1_LOC_574/A 0.43fF
C31015 AND2X1_LOC_7/B OR2X1_LOC_598/A 0.27fF
C31016 AND2X1_LOC_95/Y AND2X1_LOC_3/Y 0.20fF
C31017 AND2X1_LOC_555/Y AND2X1_LOC_562/Y 0.01fF
C31018 AND2X1_LOC_192/Y AND2X1_LOC_739/a_8_24# 0.03fF
C31019 OR2X1_LOC_105/Y AND2X1_LOC_51/Y 0.01fF
C31020 OR2X1_LOC_89/A AND2X1_LOC_621/Y 13.91fF
C31021 OR2X1_LOC_648/a_8_216# OR2X1_LOC_78/B 0.01fF
C31022 OR2X1_LOC_61/Y OR2X1_LOC_206/a_8_216# 0.03fF
C31023 OR2X1_LOC_26/Y AND2X1_LOC_668/a_8_24# 0.04fF
C31024 OR2X1_LOC_848/a_8_216# OR2X1_LOC_269/B -0.00fF
C31025 OR2X1_LOC_633/Y OR2X1_LOC_647/B 0.07fF
C31026 OR2X1_LOC_744/A INPUT_1 0.14fF
C31027 OR2X1_LOC_600/A AND2X1_LOC_866/A 0.11fF
C31028 OR2X1_LOC_65/B OR2X1_LOC_7/A 0.03fF
C31029 OR2X1_LOC_158/a_8_216# OR2X1_LOC_158/B 0.02fF
C31030 AND2X1_LOC_352/B AND2X1_LOC_863/Y 0.02fF
C31031 OR2X1_LOC_132/a_8_216# AND2X1_LOC_656/Y 0.05fF
C31032 AND2X1_LOC_48/A OR2X1_LOC_706/A 0.03fF
C31033 OR2X1_LOC_654/A AND2X1_LOC_43/B 0.01fF
C31034 OR2X1_LOC_161/B OR2X1_LOC_544/a_36_216# 0.00fF
C31035 AND2X1_LOC_392/A AND2X1_LOC_864/a_36_24# 0.01fF
C31036 OR2X1_LOC_364/A OR2X1_LOC_810/A 0.07fF
C31037 OR2X1_LOC_185/Y OR2X1_LOC_810/A 0.10fF
C31038 OR2X1_LOC_325/a_8_216# OR2X1_LOC_121/B 0.01fF
C31039 OR2X1_LOC_43/A AND2X1_LOC_361/A 0.07fF
C31040 OR2X1_LOC_426/B AND2X1_LOC_476/A 0.25fF
C31041 AND2X1_LOC_36/Y OR2X1_LOC_195/a_8_216# 0.01fF
C31042 OR2X1_LOC_756/B OR2X1_LOC_545/B 0.02fF
C31043 OR2X1_LOC_334/B D_INPUT_0 0.04fF
C31044 AND2X1_LOC_40/Y OR2X1_LOC_444/B 0.05fF
C31045 OR2X1_LOC_218/Y OR2X1_LOC_78/A 0.01fF
C31046 OR2X1_LOC_81/Y OR2X1_LOC_585/A 0.03fF
C31047 OR2X1_LOC_840/A OR2X1_LOC_168/A 0.05fF
C31048 AND2X1_LOC_711/a_8_24# AND2X1_LOC_866/A 0.02fF
C31049 OR2X1_LOC_516/A OR2X1_LOC_70/Y 0.03fF
C31050 OR2X1_LOC_643/A OR2X1_LOC_643/a_8_216# 0.02fF
C31051 OR2X1_LOC_223/A OR2X1_LOC_741/Y 0.00fF
C31052 OR2X1_LOC_455/A OR2X1_LOC_553/A 0.03fF
C31053 OR2X1_LOC_271/Y OR2X1_LOC_7/A 0.15fF
C31054 AND2X1_LOC_3/Y OR2X1_LOC_99/Y 0.25fF
C31055 OR2X1_LOC_676/Y OR2X1_LOC_214/B 0.07fF
C31056 OR2X1_LOC_275/a_8_216# OR2X1_LOC_39/A 0.03fF
C31057 AND2X1_LOC_59/Y OR2X1_LOC_479/a_8_216# 0.01fF
C31058 OR2X1_LOC_276/B OR2X1_LOC_630/B 0.01fF
C31059 OR2X1_LOC_605/B OR2X1_LOC_87/A 0.15fF
C31060 OR2X1_LOC_185/A OR2X1_LOC_520/B 0.10fF
C31061 OR2X1_LOC_70/Y AND2X1_LOC_317/a_36_24# 0.00fF
C31062 AND2X1_LOC_543/a_8_24# AND2X1_LOC_866/A 0.03fF
C31063 AND2X1_LOC_842/B OR2X1_LOC_39/A 0.26fF
C31064 OR2X1_LOC_189/Y AND2X1_LOC_220/Y 0.11fF
C31065 AND2X1_LOC_12/Y OR2X1_LOC_206/A 0.01fF
C31066 AND2X1_LOC_721/a_8_24# OR2X1_LOC_417/A 0.04fF
C31067 AND2X1_LOC_810/Y OR2X1_LOC_594/a_8_216# 0.03fF
C31068 OR2X1_LOC_532/B OR2X1_LOC_785/B 0.09fF
C31069 OR2X1_LOC_485/A OR2X1_LOC_585/A 0.08fF
C31070 OR2X1_LOC_44/Y AND2X1_LOC_211/a_36_24# 0.01fF
C31071 AND2X1_LOC_784/A OR2X1_LOC_417/a_8_216# 0.03fF
C31072 INPUT_0 D_INPUT_1 0.25fF
C31073 OR2X1_LOC_318/Y AND2X1_LOC_47/Y 0.17fF
C31074 OR2X1_LOC_52/Y OR2X1_LOC_6/A 0.01fF
C31075 OR2X1_LOC_295/Y AND2X1_LOC_848/Y 0.03fF
C31076 OR2X1_LOC_776/Y OR2X1_LOC_318/B 0.05fF
C31077 OR2X1_LOC_36/Y OR2X1_LOC_416/Y 0.04fF
C31078 OR2X1_LOC_706/B OR2X1_LOC_375/A 0.05fF
C31079 AND2X1_LOC_728/a_36_24# AND2X1_LOC_147/Y 0.00fF
C31080 AND2X1_LOC_212/Y AND2X1_LOC_212/a_8_24# 0.01fF
C31081 OR2X1_LOC_770/A OR2X1_LOC_771/B 0.30fF
C31082 OR2X1_LOC_426/a_8_216# OR2X1_LOC_427/Y 0.40fF
C31083 OR2X1_LOC_503/A OR2X1_LOC_71/Y 0.02fF
C31084 OR2X1_LOC_54/Y OR2X1_LOC_820/B 0.53fF
C31085 AND2X1_LOC_866/A OR2X1_LOC_619/Y 0.04fF
C31086 AND2X1_LOC_468/B AND2X1_LOC_810/Y 0.02fF
C31087 AND2X1_LOC_465/A OR2X1_LOC_183/Y 0.08fF
C31088 OR2X1_LOC_87/A OR2X1_LOC_782/a_36_216# 0.00fF
C31089 OR2X1_LOC_51/Y AND2X1_LOC_562/Y 0.03fF
C31090 AND2X1_LOC_716/a_8_24# D_INPUT_0 0.01fF
C31091 OR2X1_LOC_772/B D_INPUT_1 0.60fF
C31092 OR2X1_LOC_207/B AND2X1_LOC_41/Y 0.00fF
C31093 AND2X1_LOC_657/Y OR2X1_LOC_746/Y 0.29fF
C31094 AND2X1_LOC_47/Y OR2X1_LOC_805/A 0.10fF
C31095 OR2X1_LOC_761/a_8_216# AND2X1_LOC_434/Y 0.02fF
C31096 OR2X1_LOC_51/a_8_216# OR2X1_LOC_2/Y 0.01fF
C31097 AND2X1_LOC_807/Y OR2X1_LOC_95/Y 1.21fF
C31098 OR2X1_LOC_45/B OR2X1_LOC_142/Y 0.03fF
C31099 AND2X1_LOC_64/Y OR2X1_LOC_356/B 0.28fF
C31100 AND2X1_LOC_92/Y OR2X1_LOC_228/Y 0.19fF
C31101 OR2X1_LOC_857/A AND2X1_LOC_36/Y 0.13fF
C31102 AND2X1_LOC_139/a_8_24# AND2X1_LOC_216/A 0.17fF
C31103 AND2X1_LOC_476/Y OR2X1_LOC_437/A 0.10fF
C31104 AND2X1_LOC_95/Y OR2X1_LOC_270/Y 0.03fF
C31105 AND2X1_LOC_566/B AND2X1_LOC_212/a_36_24# 0.00fF
C31106 OR2X1_LOC_160/B OR2X1_LOC_446/B 0.07fF
C31107 OR2X1_LOC_3/Y OR2X1_LOC_7/a_8_216# 0.01fF
C31108 AND2X1_LOC_557/Y D_INPUT_3 0.04fF
C31109 AND2X1_LOC_535/Y OR2X1_LOC_13/B 0.01fF
C31110 OR2X1_LOC_489/B D_INPUT_1 0.02fF
C31111 OR2X1_LOC_780/a_8_216# OR2X1_LOC_449/B 0.01fF
C31112 AND2X1_LOC_510/a_8_24# AND2X1_LOC_657/A 0.01fF
C31113 AND2X1_LOC_512/Y OR2X1_LOC_534/a_36_216# 0.01fF
C31114 OR2X1_LOC_499/B OR2X1_LOC_68/B 0.03fF
C31115 AND2X1_LOC_554/B AND2X1_LOC_845/Y 0.02fF
C31116 INPUT_4 OR2X1_LOC_51/B 0.10fF
C31117 OR2X1_LOC_462/a_8_216# OR2X1_LOC_416/Y 0.05fF
C31118 OR2X1_LOC_755/A AND2X1_LOC_814/a_8_24# 0.01fF
C31119 OR2X1_LOC_85/A AND2X1_LOC_837/a_8_24# 0.01fF
C31120 OR2X1_LOC_211/a_8_216# OR2X1_LOC_365/B 0.01fF
C31121 AND2X1_LOC_46/a_36_24# OR2X1_LOC_121/B 0.01fF
C31122 AND2X1_LOC_110/Y OR2X1_LOC_532/Y 0.02fF
C31123 OR2X1_LOC_109/Y OR2X1_LOC_406/A 0.01fF
C31124 OR2X1_LOC_621/B AND2X1_LOC_36/Y 0.12fF
C31125 OR2X1_LOC_296/Y AND2X1_LOC_47/Y 0.00fF
C31126 AND2X1_LOC_216/A AND2X1_LOC_656/a_36_24# 0.00fF
C31127 OR2X1_LOC_205/a_36_216# OR2X1_LOC_786/Y 0.00fF
C31128 OR2X1_LOC_10/a_8_216# OR2X1_LOC_585/A 0.01fF
C31129 OR2X1_LOC_743/A AND2X1_LOC_476/A 0.08fF
C31130 OR2X1_LOC_34/A AND2X1_LOC_7/B 0.00fF
C31131 OR2X1_LOC_805/A OR2X1_LOC_717/a_36_216# 0.01fF
C31132 AND2X1_LOC_555/Y OR2X1_LOC_381/a_8_216# 0.03fF
C31133 AND2X1_LOC_51/A OR2X1_LOC_51/B 0.00fF
C31134 AND2X1_LOC_84/Y OR2X1_LOC_16/A 0.14fF
C31135 OR2X1_LOC_64/Y OR2X1_LOC_71/Y 0.11fF
C31136 OR2X1_LOC_203/Y OR2X1_LOC_493/Y 0.10fF
C31137 OR2X1_LOC_624/A AND2X1_LOC_31/Y 0.10fF
C31138 OR2X1_LOC_173/Y OR2X1_LOC_173/a_8_216# -0.00fF
C31139 OR2X1_LOC_488/Y OR2X1_LOC_95/Y 0.09fF
C31140 OR2X1_LOC_323/A OR2X1_LOC_158/A 0.03fF
C31141 OR2X1_LOC_207/B AND2X1_LOC_22/Y 0.01fF
C31142 OR2X1_LOC_186/Y OR2X1_LOC_175/Y 0.59fF
C31143 OR2X1_LOC_143/a_8_216# VDD 0.21fF
C31144 AND2X1_LOC_802/B AND2X1_LOC_810/B 0.02fF
C31145 OR2X1_LOC_47/Y AND2X1_LOC_211/a_8_24# 0.05fF
C31146 AND2X1_LOC_7/B AND2X1_LOC_627/a_36_24# 0.00fF
C31147 OR2X1_LOC_294/Y OR2X1_LOC_563/A -0.00fF
C31148 OR2X1_LOC_606/Y OR2X1_LOC_532/B 0.00fF
C31149 OR2X1_LOC_76/Y OR2X1_LOC_318/B 0.11fF
C31150 OR2X1_LOC_78/A OR2X1_LOC_703/Y 0.06fF
C31151 OR2X1_LOC_144/a_36_216# OR2X1_LOC_526/Y 0.00fF
C31152 AND2X1_LOC_727/A OR2X1_LOC_95/Y 0.03fF
C31153 OR2X1_LOC_186/Y AND2X1_LOC_417/a_8_24# 0.02fF
C31154 OR2X1_LOC_363/B OR2X1_LOC_363/a_8_216# 0.00fF
C31155 OR2X1_LOC_348/Y OR2X1_LOC_366/A 0.03fF
C31156 AND2X1_LOC_724/A OR2X1_LOC_16/A 0.00fF
C31157 OR2X1_LOC_158/A OR2X1_LOC_744/a_8_216# 0.01fF
C31158 AND2X1_LOC_350/a_8_24# AND2X1_LOC_350/B 0.01fF
C31159 OR2X1_LOC_56/A AND2X1_LOC_439/a_36_24# 0.01fF
C31160 OR2X1_LOC_246/A AND2X1_LOC_476/A 0.10fF
C31161 OR2X1_LOC_31/Y INPUT_1 0.42fF
C31162 OR2X1_LOC_71/Y OR2X1_LOC_417/A 0.03fF
C31163 OR2X1_LOC_121/B OR2X1_LOC_340/a_8_216# 0.01fF
C31164 AND2X1_LOC_763/a_8_24# AND2X1_LOC_763/B 0.00fF
C31165 OR2X1_LOC_296/Y OR2X1_LOC_598/A 0.00fF
C31166 OR2X1_LOC_841/a_8_216# AND2X1_LOC_36/Y 0.00fF
C31167 OR2X1_LOC_36/Y OR2X1_LOC_80/A 0.16fF
C31168 OR2X1_LOC_177/Y OR2X1_LOC_322/a_8_216# 0.01fF
C31169 OR2X1_LOC_78/B OR2X1_LOC_390/B 0.02fF
C31170 OR2X1_LOC_544/A OR2X1_LOC_439/a_8_216# 0.47fF
C31171 OR2X1_LOC_117/a_8_216# AND2X1_LOC_243/Y 0.03fF
C31172 OR2X1_LOC_799/a_8_216# OR2X1_LOC_446/B 0.01fF
C31173 OR2X1_LOC_362/A OR2X1_LOC_161/B 0.01fF
C31174 OR2X1_LOC_501/B OR2X1_LOC_140/B 0.03fF
C31175 AND2X1_LOC_732/B OR2X1_LOC_428/A 0.01fF
C31176 AND2X1_LOC_64/Y OR2X1_LOC_168/B 0.20fF
C31177 OR2X1_LOC_756/B OR2X1_LOC_363/a_8_216# 0.02fF
C31178 OR2X1_LOC_114/B OR2X1_LOC_342/A 0.04fF
C31179 AND2X1_LOC_42/B OR2X1_LOC_398/Y 0.03fF
C31180 OR2X1_LOC_95/Y OR2X1_LOC_368/A 0.05fF
C31181 OR2X1_LOC_289/Y OR2X1_LOC_46/A 0.01fF
C31182 AND2X1_LOC_654/B OR2X1_LOC_387/A 0.14fF
C31183 OR2X1_LOC_36/Y AND2X1_LOC_592/a_8_24# 0.01fF
C31184 OR2X1_LOC_724/a_8_216# OR2X1_LOC_308/Y 0.04fF
C31185 OR2X1_LOC_246/Y OR2X1_LOC_13/B 0.20fF
C31186 OR2X1_LOC_532/B OR2X1_LOC_786/Y 0.04fF
C31187 OR2X1_LOC_666/A AND2X1_LOC_244/A 0.03fF
C31188 VDD AND2X1_LOC_338/A -0.00fF
C31189 OR2X1_LOC_790/a_8_216# AND2X1_LOC_41/Y 0.00fF
C31190 OR2X1_LOC_696/A AND2X1_LOC_852/B 0.03fF
C31191 AND2X1_LOC_705/Y OR2X1_LOC_600/a_8_216# 0.01fF
C31192 OR2X1_LOC_793/a_8_216# AND2X1_LOC_36/Y 0.01fF
C31193 OR2X1_LOC_476/B OR2X1_LOC_358/A 0.00fF
C31194 VDD OR2X1_LOC_356/A 0.48fF
C31195 OR2X1_LOC_49/A OR2X1_LOC_78/A 0.07fF
C31196 VDD OR2X1_LOC_654/a_8_216# 0.21fF
C31197 OR2X1_LOC_696/A OR2X1_LOC_48/B 3.00fF
C31198 OR2X1_LOC_160/B OR2X1_LOC_719/B 0.02fF
C31199 AND2X1_LOC_553/A AND2X1_LOC_465/A 0.00fF
C31200 OR2X1_LOC_347/A OR2X1_LOC_347/B 0.06fF
C31201 OR2X1_LOC_6/B OR2X1_LOC_96/Y 0.03fF
C31202 OR2X1_LOC_696/A OR2X1_LOC_18/Y 4.93fF
C31203 OR2X1_LOC_108/a_36_216# OR2X1_LOC_108/Y 0.01fF
C31204 OR2X1_LOC_814/A OR2X1_LOC_675/Y 0.03fF
C31205 OR2X1_LOC_40/Y OR2X1_LOC_600/A 0.32fF
C31206 OR2X1_LOC_40/Y AND2X1_LOC_335/Y 0.01fF
C31207 OR2X1_LOC_462/a_36_216# OR2X1_LOC_68/B 0.00fF
C31208 OR2X1_LOC_794/a_8_216# OR2X1_LOC_303/B 0.02fF
C31209 OR2X1_LOC_528/Y AND2X1_LOC_658/B 0.57fF
C31210 OR2X1_LOC_92/Y AND2X1_LOC_476/a_8_24# 0.14fF
C31211 OR2X1_LOC_833/Y OR2X1_LOC_541/A 0.02fF
C31212 OR2X1_LOC_78/A OR2X1_LOC_596/A 2.54fF
C31213 OR2X1_LOC_536/Y AND2X1_LOC_537/a_8_24# 0.23fF
C31214 AND2X1_LOC_3/Y AND2X1_LOC_41/Y 0.03fF
C31215 VDD OR2X1_LOC_20/Y 0.12fF
C31216 AND2X1_LOC_281/a_8_24# OR2X1_LOC_366/Y 0.02fF
C31217 OR2X1_LOC_474/Y OR2X1_LOC_161/B 0.03fF
C31218 VDD AND2X1_LOC_112/a_8_24# 0.00fF
C31219 OR2X1_LOC_92/Y OR2X1_LOC_753/a_8_216# 0.01fF
C31220 AND2X1_LOC_715/Y OR2X1_LOC_48/B 0.02fF
C31221 AND2X1_LOC_728/Y AND2X1_LOC_209/Y 0.01fF
C31222 OR2X1_LOC_539/A OR2X1_LOC_161/B 0.01fF
C31223 AND2X1_LOC_64/Y AND2X1_LOC_59/Y 6.91fF
C31224 AND2X1_LOC_601/a_36_24# OR2X1_LOC_390/B 0.01fF
C31225 AND2X1_LOC_554/Y OR2X1_LOC_106/Y 0.02fF
C31226 OR2X1_LOC_101/a_36_216# AND2X1_LOC_22/Y 0.02fF
C31227 AND2X1_LOC_721/Y OR2X1_LOC_278/Y 0.01fF
C31228 OR2X1_LOC_450/A OR2X1_LOC_467/A 0.00fF
C31229 AND2X1_LOC_716/Y OR2X1_LOC_16/A 0.07fF
C31230 OR2X1_LOC_447/Y AND2X1_LOC_31/Y 0.03fF
C31231 OR2X1_LOC_506/A AND2X1_LOC_7/B 0.15fF
C31232 OR2X1_LOC_22/Y OR2X1_LOC_521/a_8_216# 0.01fF
C31233 OR2X1_LOC_770/A OR2X1_LOC_402/Y 0.01fF
C31234 OR2X1_LOC_405/A OR2X1_LOC_139/A 0.13fF
C31235 OR2X1_LOC_35/Y OR2X1_LOC_66/A 0.33fF
C31236 OR2X1_LOC_351/B OR2X1_LOC_756/B 0.38fF
C31237 OR2X1_LOC_768/A AND2X1_LOC_18/Y 0.01fF
C31238 AND2X1_LOC_352/a_36_24# OR2X1_LOC_91/A 0.00fF
C31239 AND2X1_LOC_12/Y OR2X1_LOC_362/a_8_216# 0.01fF
C31240 OR2X1_LOC_744/A AND2X1_LOC_325/a_8_24# 0.06fF
C31241 OR2X1_LOC_625/Y OR2X1_LOC_428/A 0.02fF
C31242 AND2X1_LOC_654/Y OR2X1_LOC_16/A 0.07fF
C31243 OR2X1_LOC_45/B OR2X1_LOC_118/Y 0.02fF
C31244 OR2X1_LOC_426/B OR2X1_LOC_122/A 0.02fF
C31245 OR2X1_LOC_347/B AND2X1_LOC_44/Y 0.01fF
C31246 OR2X1_LOC_427/A AND2X1_LOC_212/Y 0.07fF
C31247 AND2X1_LOC_71/a_8_24# AND2X1_LOC_18/Y 0.02fF
C31248 OR2X1_LOC_426/B INPUT_0 0.10fF
C31249 OR2X1_LOC_40/Y AND2X1_LOC_862/Y 0.07fF
C31250 OR2X1_LOC_696/A OR2X1_LOC_385/Y 0.17fF
C31251 AND2X1_LOC_42/B AND2X1_LOC_619/a_8_24# 0.02fF
C31252 OR2X1_LOC_692/Y AND2X1_LOC_644/Y 0.03fF
C31253 AND2X1_LOC_498/a_8_24# AND2X1_LOC_92/Y 0.01fF
C31254 AND2X1_LOC_70/Y OR2X1_LOC_630/B 0.01fF
C31255 OR2X1_LOC_325/A AND2X1_LOC_110/Y 0.01fF
C31256 AND2X1_LOC_735/Y AND2X1_LOC_501/a_8_24# 0.17fF
C31257 OR2X1_LOC_756/B AND2X1_LOC_396/a_8_24# 0.01fF
C31258 OR2X1_LOC_673/Y OR2X1_LOC_720/Y 0.06fF
C31259 OR2X1_LOC_11/Y OR2X1_LOC_585/a_8_216# 0.01fF
C31260 VDD OR2X1_LOC_746/a_8_216# 0.21fF
C31261 AND2X1_LOC_456/B AND2X1_LOC_285/Y 0.35fF
C31262 AND2X1_LOC_566/B AND2X1_LOC_841/B 0.03fF
C31263 OR2X1_LOC_185/A OR2X1_LOC_486/Y 0.22fF
C31264 OR2X1_LOC_648/A AND2X1_LOC_41/A 0.07fF
C31265 OR2X1_LOC_135/Y AND2X1_LOC_138/a_8_24# 0.01fF
C31266 OR2X1_LOC_779/a_8_216# AND2X1_LOC_44/Y 0.01fF
C31267 OR2X1_LOC_44/Y AND2X1_LOC_208/Y 0.02fF
C31268 OR2X1_LOC_210/a_8_216# OR2X1_LOC_160/Y 0.01fF
C31269 OR2X1_LOC_92/a_8_216# OR2X1_LOC_71/A 0.01fF
C31270 OR2X1_LOC_563/B OR2X1_LOC_562/A 0.00fF
C31271 OR2X1_LOC_485/A AND2X1_LOC_455/a_8_24# 0.08fF
C31272 OR2X1_LOC_36/Y AND2X1_LOC_206/a_36_24# 0.00fF
C31273 OR2X1_LOC_840/a_8_216# OR2X1_LOC_375/A 0.01fF
C31274 AND2X1_LOC_715/a_8_24# OR2X1_LOC_428/A 0.06fF
C31275 AND2X1_LOC_22/Y AND2X1_LOC_7/a_36_24# 0.00fF
C31276 AND2X1_LOC_474/A AND2X1_LOC_860/a_8_24# 0.08fF
C31277 OR2X1_LOC_744/A OR2X1_LOC_517/A 0.06fF
C31278 OR2X1_LOC_441/Y AND2X1_LOC_663/A 0.05fF
C31279 OR2X1_LOC_45/B OR2X1_LOC_262/Y 0.27fF
C31280 OR2X1_LOC_621/a_36_216# OR2X1_LOC_847/A 0.00fF
C31281 OR2X1_LOC_40/Y OR2X1_LOC_619/Y 0.24fF
C31282 AND2X1_LOC_564/B OR2X1_LOC_485/A 0.07fF
C31283 AND2X1_LOC_794/A OR2X1_LOC_600/A -0.01fF
C31284 OR2X1_LOC_624/a_8_216# OR2X1_LOC_659/A 0.02fF
C31285 OR2X1_LOC_91/Y AND2X1_LOC_443/a_8_24# -0.00fF
C31286 AND2X1_LOC_22/Y AND2X1_LOC_3/Y 0.35fF
C31287 OR2X1_LOC_553/A OR2X1_LOC_719/B 0.02fF
C31288 OR2X1_LOC_97/A OR2X1_LOC_574/A 0.03fF
C31289 OR2X1_LOC_45/B OR2X1_LOC_238/Y 0.03fF
C31290 OR2X1_LOC_87/A OR2X1_LOC_549/A 0.08fF
C31291 AND2X1_LOC_366/a_8_24# OR2X1_LOC_427/A 0.01fF
C31292 OR2X1_LOC_744/A AND2X1_LOC_651/a_36_24# 0.00fF
C31293 AND2X1_LOC_725/a_8_24# AND2X1_LOC_448/Y 0.06fF
C31294 OR2X1_LOC_485/A OR2X1_LOC_530/a_8_216# 0.04fF
C31295 AND2X1_LOC_385/a_8_24# OR2X1_LOC_390/A 0.24fF
C31296 AND2X1_LOC_367/A AND2X1_LOC_344/a_8_24# 0.02fF
C31297 OR2X1_LOC_312/Y OR2X1_LOC_16/A 0.05fF
C31298 AND2X1_LOC_486/Y AND2X1_LOC_471/Y 0.09fF
C31299 AND2X1_LOC_535/a_8_24# OR2X1_LOC_619/Y 0.03fF
C31300 AND2X1_LOC_33/a_8_24# OR2X1_LOC_18/Y 0.01fF
C31301 OR2X1_LOC_364/A OR2X1_LOC_715/B 0.10fF
C31302 AND2X1_LOC_753/B OR2X1_LOC_637/Y 0.08fF
C31303 OR2X1_LOC_653/Y AND2X1_LOC_20/a_8_24# 0.05fF
C31304 INPUT_0 AND2X1_LOC_414/a_8_24# 0.02fF
C31305 OR2X1_LOC_185/Y OR2X1_LOC_715/B 0.35fF
C31306 VDD AND2X1_LOC_43/B 1.38fF
C31307 OR2X1_LOC_40/Y OR2X1_LOC_88/A 0.01fF
C31308 OR2X1_LOC_51/Y AND2X1_LOC_287/a_8_24# 0.01fF
C31309 OR2X1_LOC_861/a_8_216# OR2X1_LOC_624/Y 0.02fF
C31310 OR2X1_LOC_363/B AND2X1_LOC_12/Y 0.26fF
C31311 OR2X1_LOC_9/Y OR2X1_LOC_43/A 2.80fF
C31312 AND2X1_LOC_561/B AND2X1_LOC_573/A 0.03fF
C31313 OR2X1_LOC_151/A OR2X1_LOC_778/Y 0.14fF
C31314 OR2X1_LOC_43/A AND2X1_LOC_193/Y 0.01fF
C31315 OR2X1_LOC_542/B OR2X1_LOC_553/A 0.07fF
C31316 OR2X1_LOC_858/A OR2X1_LOC_161/A 0.03fF
C31317 OR2X1_LOC_155/A OR2X1_LOC_596/A 0.05fF
C31318 AND2X1_LOC_390/B AND2X1_LOC_774/A 0.10fF
C31319 AND2X1_LOC_95/Y INPUT_0 0.17fF
C31320 OR2X1_LOC_160/B AND2X1_LOC_56/B 0.06fF
C31321 AND2X1_LOC_359/B AND2X1_LOC_860/A 0.03fF
C31322 OR2X1_LOC_659/Y OR2X1_LOC_624/B 0.01fF
C31323 OR2X1_LOC_160/B OR2X1_LOC_659/B 0.03fF
C31324 OR2X1_LOC_106/Y OR2X1_LOC_22/Y 0.01fF
C31325 AND2X1_LOC_58/a_8_24# OR2X1_LOC_61/B 0.01fF
C31326 OR2X1_LOC_509/A OR2X1_LOC_502/A 0.03fF
C31327 OR2X1_LOC_534/Y OR2X1_LOC_331/Y 0.07fF
C31328 OR2X1_LOC_779/Y OR2X1_LOC_712/B 0.05fF
C31329 AND2X1_LOC_40/Y AND2X1_LOC_328/a_8_24# 0.04fF
C31330 OR2X1_LOC_394/Y OR2X1_LOC_394/a_36_216# 0.00fF
C31331 OR2X1_LOC_633/B OR2X1_LOC_786/A 0.01fF
C31332 AND2X1_LOC_81/B OR2X1_LOC_242/a_8_216# 0.01fF
C31333 AND2X1_LOC_51/Y OR2X1_LOC_355/a_8_216# 0.01fF
C31334 AND2X1_LOC_12/Y OR2X1_LOC_756/B 0.41fF
C31335 OR2X1_LOC_814/A OR2X1_LOC_174/a_36_216# 0.01fF
C31336 OR2X1_LOC_720/a_8_216# OR2X1_LOC_66/A 0.01fF
C31337 AND2X1_LOC_719/Y OR2X1_LOC_371/Y 0.10fF
C31338 AND2X1_LOC_486/Y AND2X1_LOC_840/A 0.03fF
C31339 OR2X1_LOC_744/A OR2X1_LOC_380/A 0.15fF
C31340 OR2X1_LOC_114/B AND2X1_LOC_159/a_36_24# 0.00fF
C31341 OR2X1_LOC_626/a_8_216# OR2X1_LOC_626/Y 0.01fF
C31342 AND2X1_LOC_716/Y AND2X1_LOC_168/Y 0.51fF
C31343 OR2X1_LOC_319/B OR2X1_LOC_506/A 0.07fF
C31344 OR2X1_LOC_468/A OR2X1_LOC_592/a_8_216# 0.01fF
C31345 AND2X1_LOC_810/A AND2X1_LOC_802/a_8_24# 0.01fF
C31346 OR2X1_LOC_600/A OR2X1_LOC_7/A 0.41fF
C31347 OR2X1_LOC_158/A OR2X1_LOC_275/A 0.02fF
C31348 AND2X1_LOC_560/a_36_24# OR2X1_LOC_95/Y 0.00fF
C31349 AND2X1_LOC_654/Y AND2X1_LOC_661/a_8_24# 0.11fF
C31350 AND2X1_LOC_59/Y OR2X1_LOC_656/Y 0.10fF
C31351 OR2X1_LOC_70/Y OR2X1_LOC_765/Y 0.01fF
C31352 AND2X1_LOC_303/B AND2X1_LOC_303/a_8_24# 0.01fF
C31353 OR2X1_LOC_26/Y OR2X1_LOC_59/Y 2.11fF
C31354 OR2X1_LOC_22/Y AND2X1_LOC_219/A 5.45fF
C31355 OR2X1_LOC_492/Y OR2X1_LOC_64/Y 0.07fF
C31356 OR2X1_LOC_318/Y OR2X1_LOC_506/A 0.08fF
C31357 AND2X1_LOC_675/Y AND2X1_LOC_806/A 0.23fF
C31358 OR2X1_LOC_6/B OR2X1_LOC_123/B 0.03fF
C31359 OR2X1_LOC_703/B OR2X1_LOC_354/A 0.01fF
C31360 VDD AND2X1_LOC_148/Y 0.29fF
C31361 OR2X1_LOC_8/Y OR2X1_LOC_278/a_8_216# 0.14fF
C31362 OR2X1_LOC_51/Y OR2X1_LOC_239/Y 0.16fF
C31363 INPUT_1 AND2X1_LOC_464/A 0.17fF
C31364 AND2X1_LOC_493/a_8_24# OR2X1_LOC_59/Y 0.03fF
C31365 OR2X1_LOC_375/A AND2X1_LOC_422/a_8_24# 0.01fF
C31366 AND2X1_LOC_717/a_8_24# OR2X1_LOC_18/Y 0.02fF
C31367 VDD AND2X1_LOC_660/Y 0.21fF
C31368 OR2X1_LOC_89/A OR2X1_LOC_59/Y 7.63fF
C31369 OR2X1_LOC_676/Y OR2X1_LOC_193/A 0.03fF
C31370 OR2X1_LOC_653/B OR2X1_LOC_814/A 0.02fF
C31371 OR2X1_LOC_95/a_8_216# OR2X1_LOC_586/Y 0.10fF
C31372 AND2X1_LOC_99/A OR2X1_LOC_67/A 0.01fF
C31373 OR2X1_LOC_47/Y AND2X1_LOC_213/a_8_24# 0.02fF
C31374 OR2X1_LOC_321/Y OR2X1_LOC_56/A 0.01fF
C31375 AND2X1_LOC_95/Y OR2X1_LOC_128/a_8_216# 0.07fF
C31376 OR2X1_LOC_244/B AND2X1_LOC_3/Y 0.02fF
C31377 INPUT_0 OR2X1_LOC_743/A 0.04fF
C31378 OR2X1_LOC_467/A OR2X1_LOC_470/B 0.03fF
C31379 OR2X1_LOC_524/Y OR2X1_LOC_438/a_8_216# 0.12fF
C31380 AND2X1_LOC_593/Y AND2X1_LOC_652/a_8_24# 0.04fF
C31381 OR2X1_LOC_128/A OR2X1_LOC_128/B 0.05fF
C31382 AND2X1_LOC_47/Y OR2X1_LOC_580/B 0.03fF
C31383 AND2X1_LOC_543/a_8_24# OR2X1_LOC_7/A 0.01fF
C31384 AND2X1_LOC_833/a_8_24# AND2X1_LOC_840/B 0.01fF
C31385 OR2X1_LOC_506/A OR2X1_LOC_805/A 0.02fF
C31386 VDD OR2X1_LOC_683/Y 0.12fF
C31387 OR2X1_LOC_175/Y OR2X1_LOC_112/B 0.00fF
C31388 OR2X1_LOC_92/Y OR2X1_LOC_86/a_8_216# 0.01fF
C31389 OR2X1_LOC_75/a_8_216# OR2X1_LOC_16/A 0.01fF
C31390 OR2X1_LOC_97/a_8_216# AND2X1_LOC_92/Y 0.14fF
C31391 OR2X1_LOC_18/Y AND2X1_LOC_458/Y 0.01fF
C31392 OR2X1_LOC_426/B OR2X1_LOC_64/Y 0.16fF
C31393 AND2X1_LOC_362/B AND2X1_LOC_845/Y 0.09fF
C31394 AND2X1_LOC_633/a_8_24# OR2X1_LOC_39/A 0.01fF
C31395 AND2X1_LOC_7/B D_INPUT_1 0.07fF
C31396 OR2X1_LOC_271/B OR2X1_LOC_18/Y 0.11fF
C31397 OR2X1_LOC_808/A OR2X1_LOC_605/A 0.24fF
C31398 AND2X1_LOC_573/A AND2X1_LOC_266/Y 0.02fF
C31399 INPUT_3 AND2X1_LOC_56/B 0.01fF
C31400 OR2X1_LOC_431/Y AND2X1_LOC_434/a_8_24# 0.04fF
C31401 AND2X1_LOC_824/B AND2X1_LOC_291/a_8_24# 0.01fF
C31402 AND2X1_LOC_86/Y AND2X1_LOC_8/Y 0.18fF
C31403 OR2X1_LOC_377/A OR2X1_LOC_835/a_8_216# 0.01fF
C31404 OR2X1_LOC_624/A OR2X1_LOC_809/a_8_216# 0.02fF
C31405 AND2X1_LOC_359/a_8_24# OR2X1_LOC_18/Y 0.17fF
C31406 D_INPUT_5 AND2X1_LOC_459/a_36_24# 0.00fF
C31407 OR2X1_LOC_641/Y OR2X1_LOC_814/A 0.14fF
C31408 AND2X1_LOC_301/a_8_24# INPUT_1 0.01fF
C31409 INPUT_3 AND2X1_LOC_8/Y 0.02fF
C31410 AND2X1_LOC_29/a_8_24# OR2X1_LOC_375/A 0.03fF
C31411 OR2X1_LOC_256/a_8_216# OR2X1_LOC_585/A 0.01fF
C31412 OR2X1_LOC_377/A OR2X1_LOC_836/a_8_216# 0.05fF
C31413 AND2X1_LOC_56/B OR2X1_LOC_553/A 0.07fF
C31414 AND2X1_LOC_175/B AND2X1_LOC_654/a_8_24# 0.20fF
C31415 AND2X1_LOC_91/a_8_24# OR2X1_LOC_374/Y 0.02fF
C31416 AND2X1_LOC_701/a_8_24# OR2X1_LOC_161/A 0.04fF
C31417 OR2X1_LOC_630/a_8_216# AND2X1_LOC_3/Y 0.01fF
C31418 OR2X1_LOC_18/Y OR2X1_LOC_89/a_8_216# 0.04fF
C31419 OR2X1_LOC_7/A OR2X1_LOC_619/Y 0.28fF
C31420 AND2X1_LOC_325/a_8_24# OR2X1_LOC_31/Y 0.02fF
C31421 OR2X1_LOC_36/Y OR2X1_LOC_6/A 1.29fF
C31422 OR2X1_LOC_426/B OR2X1_LOC_417/A 0.20fF
C31423 OR2X1_LOC_455/a_36_216# OR2X1_LOC_553/A 0.01fF
C31424 OR2X1_LOC_866/a_8_216# OR2X1_LOC_859/B 0.01fF
C31425 OR2X1_LOC_834/A D_INPUT_0 0.00fF
C31426 OR2X1_LOC_43/A OR2X1_LOC_96/B 0.03fF
C31427 OR2X1_LOC_203/Y OR2X1_LOC_205/a_8_216# 0.10fF
C31428 OR2X1_LOC_600/A OR2X1_LOC_224/a_8_216# 0.01fF
C31429 AND2X1_LOC_8/Y OR2X1_LOC_266/a_8_216# 0.01fF
C31430 AND2X1_LOC_775/a_8_24# OR2X1_LOC_26/Y 0.01fF
C31431 OR2X1_LOC_617/Y AND2X1_LOC_805/Y 0.03fF
C31432 OR2X1_LOC_320/Y OR2X1_LOC_619/Y 0.03fF
C31433 AND2X1_LOC_570/Y AND2X1_LOC_227/Y 0.02fF
C31434 OR2X1_LOC_777/B OR2X1_LOC_593/B 0.03fF
C31435 AND2X1_LOC_126/a_8_24# OR2X1_LOC_62/B 0.01fF
C31436 AND2X1_LOC_728/Y AND2X1_LOC_728/a_8_24# 0.02fF
C31437 AND2X1_LOC_729/Y OR2X1_LOC_680/Y 0.02fF
C31438 AND2X1_LOC_103/a_8_24# AND2X1_LOC_47/Y 0.10fF
C31439 OR2X1_LOC_47/Y OR2X1_LOC_583/Y 0.02fF
C31440 OR2X1_LOC_677/Y AND2X1_LOC_678/a_8_24# 0.11fF
C31441 OR2X1_LOC_808/B OR2X1_LOC_814/A 0.00fF
C31442 AND2X1_LOC_775/a_8_24# OR2X1_LOC_89/A 0.02fF
C31443 OR2X1_LOC_449/B OR2X1_LOC_592/a_8_216# 0.03fF
C31444 OR2X1_LOC_18/Y AND2X1_LOC_663/B 0.07fF
C31445 OR2X1_LOC_3/Y AND2X1_LOC_319/A 0.07fF
C31446 AND2X1_LOC_206/Y AND2X1_LOC_202/Y 0.00fF
C31447 AND2X1_LOC_372/a_8_24# AND2X1_LOC_47/Y 0.03fF
C31448 AND2X1_LOC_140/a_8_24# AND2X1_LOC_572/A 0.01fF
C31449 AND2X1_LOC_465/a_8_24# OR2X1_LOC_36/Y 0.01fF
C31450 AND2X1_LOC_132/a_8_24# OR2X1_LOC_404/Y 0.02fF
C31451 OR2X1_LOC_89/A OR2X1_LOC_820/B 0.02fF
C31452 OR2X1_LOC_593/B AND2X1_LOC_591/a_36_24# 0.00fF
C31453 OR2X1_LOC_517/A OR2X1_LOC_31/Y 0.13fF
C31454 OR2X1_LOC_312/Y AND2X1_LOC_336/a_8_24# 0.01fF
C31455 AND2X1_LOC_229/a_36_24# OR2X1_LOC_68/B 0.00fF
C31456 OR2X1_LOC_235/B OR2X1_LOC_673/A 0.01fF
C31457 OR2X1_LOC_820/Y OR2X1_LOC_820/B 0.01fF
C31458 AND2X1_LOC_145/a_36_24# AND2X1_LOC_51/Y 0.01fF
C31459 OR2X1_LOC_51/a_8_216# OR2X1_LOC_25/Y 0.03fF
C31460 OR2X1_LOC_296/a_8_216# AND2X1_LOC_3/Y 0.01fF
C31461 OR2X1_LOC_279/Y AND2X1_LOC_806/A 0.26fF
C31462 AND2X1_LOC_719/Y AND2X1_LOC_222/Y 0.03fF
C31463 OR2X1_LOC_70/Y OR2X1_LOC_26/Y 2.69fF
C31464 AND2X1_LOC_477/A AND2X1_LOC_468/B 0.03fF
C31465 AND2X1_LOC_388/Y OR2X1_LOC_331/Y 0.10fF
C31466 OR2X1_LOC_357/a_8_216# OR2X1_LOC_357/A 0.18fF
C31467 AND2X1_LOC_65/A OR2X1_LOC_68/B 0.00fF
C31468 OR2X1_LOC_232/Y D_INPUT_1 0.01fF
C31469 OR2X1_LOC_462/a_8_216# OR2X1_LOC_6/A 0.14fF
C31470 OR2X1_LOC_661/a_8_216# D_INPUT_0 0.01fF
C31471 AND2X1_LOC_512/Y OR2X1_LOC_47/Y 0.07fF
C31472 OR2X1_LOC_52/Y OR2X1_LOC_44/Y 0.02fF
C31473 AND2X1_LOC_784/A AND2X1_LOC_326/A 0.02fF
C31474 OR2X1_LOC_543/A OR2X1_LOC_552/A -0.00fF
C31475 OR2X1_LOC_377/A AND2X1_LOC_5/a_8_24# 0.20fF
C31476 OR2X1_LOC_45/B OR2X1_LOC_300/a_8_216# 0.01fF
C31477 OR2X1_LOC_70/Y OR2X1_LOC_89/A 2.92fF
C31478 OR2X1_LOC_831/B OR2X1_LOC_593/B 0.01fF
C31479 AND2X1_LOC_18/Y OR2X1_LOC_641/B 0.09fF
C31480 AND2X1_LOC_244/A OR2X1_LOC_13/B 0.01fF
C31481 OR2X1_LOC_18/Y AND2X1_LOC_849/a_8_24# 0.01fF
C31482 OR2X1_LOC_497/a_8_216# OR2X1_LOC_22/Y 0.01fF
C31483 AND2X1_LOC_566/a_8_24# OR2X1_LOC_417/Y 0.01fF
C31484 OR2X1_LOC_92/Y OR2X1_LOC_615/Y 0.02fF
C31485 AND2X1_LOC_56/B AND2X1_LOC_680/a_36_24# 0.00fF
C31486 OR2X1_LOC_46/A AND2X1_LOC_413/a_8_24# 0.03fF
C31487 OR2X1_LOC_743/A OR2X1_LOC_273/a_36_216# 0.01fF
C31488 AND2X1_LOC_557/a_36_24# OR2X1_LOC_89/A 0.00fF
C31489 OR2X1_LOC_78/B OR2X1_LOC_801/B 0.07fF
C31490 AND2X1_LOC_514/Y OR2X1_LOC_26/Y 0.00fF
C31491 OR2X1_LOC_271/Y AND2X1_LOC_115/a_8_24# 0.01fF
C31492 OR2X1_LOC_16/A OR2X1_LOC_599/a_36_216# 0.00fF
C31493 AND2X1_LOC_729/Y OR2X1_LOC_167/Y 0.05fF
C31494 OR2X1_LOC_636/A OR2X1_LOC_636/B 1.24fF
C31495 OR2X1_LOC_606/a_8_216# OR2X1_LOC_99/Y 0.01fF
C31496 OR2X1_LOC_65/Y OR2X1_LOC_52/B 0.28fF
C31497 OR2X1_LOC_543/A OR2X1_LOC_578/B 0.03fF
C31498 OR2X1_LOC_16/A OR2X1_LOC_13/B 0.10fF
C31499 OR2X1_LOC_464/A OR2X1_LOC_733/Y 0.02fF
C31500 AND2X1_LOC_456/B AND2X1_LOC_483/Y 0.14fF
C31501 AND2X1_LOC_546/a_8_24# AND2X1_LOC_796/Y 0.01fF
C31502 OR2X1_LOC_466/a_8_216# OR2X1_LOC_470/B -0.00fF
C31503 OR2X1_LOC_664/Y AND2X1_LOC_108/a_8_24# 0.02fF
C31504 AND2X1_LOC_512/a_8_24# OR2X1_LOC_311/Y 0.01fF
C31505 OR2X1_LOC_458/B OR2X1_LOC_374/Y 0.11fF
C31506 OR2X1_LOC_743/A OR2X1_LOC_64/Y 0.15fF
C31507 OR2X1_LOC_835/B OR2X1_LOC_532/B 0.10fF
C31508 AND2X1_LOC_232/a_36_24# OR2X1_LOC_598/A 0.00fF
C31509 OR2X1_LOC_54/Y OR2X1_LOC_240/A 0.12fF
C31510 AND2X1_LOC_679/a_36_24# OR2X1_LOC_715/A 0.00fF
C31511 OR2X1_LOC_66/A OR2X1_LOC_80/A 1.47fF
C31512 AND2X1_LOC_367/a_8_24# OR2X1_LOC_417/A 0.03fF
C31513 OR2X1_LOC_659/B OR2X1_LOC_244/A 0.01fF
C31514 OR2X1_LOC_11/Y OR2X1_LOC_409/B 0.04fF
C31515 OR2X1_LOC_3/Y AND2X1_LOC_708/a_8_24# 0.01fF
C31516 AND2X1_LOC_182/a_8_24# OR2X1_LOC_437/A 0.04fF
C31517 VDD OR2X1_LOC_357/A 0.06fF
C31518 OR2X1_LOC_596/A OR2X1_LOC_515/a_36_216# 0.00fF
C31519 AND2X1_LOC_36/Y OR2X1_LOC_578/a_8_216# 0.01fF
C31520 AND2X1_LOC_8/Y OR2X1_LOC_244/A 0.11fF
C31521 OR2X1_LOC_848/A OR2X1_LOC_770/a_36_216# 0.00fF
C31522 VDD OR2X1_LOC_367/B 1.52fF
C31523 AND2X1_LOC_273/a_8_24# OR2X1_LOC_831/B 0.01fF
C31524 AND2X1_LOC_835/a_8_24# OR2X1_LOC_585/A 0.01fF
C31525 OR2X1_LOC_428/A OR2X1_LOC_759/Y 0.03fF
C31526 VDD OR2X1_LOC_558/A 0.00fF
C31527 OR2X1_LOC_303/a_8_216# OR2X1_LOC_566/A 0.01fF
C31528 OR2X1_LOC_503/Y OR2X1_LOC_44/Y 0.01fF
C31529 OR2X1_LOC_273/a_36_216# OR2X1_LOC_246/A 0.13fF
C31530 AND2X1_LOC_342/Y OR2X1_LOC_47/Y 0.04fF
C31531 OR2X1_LOC_805/A D_INPUT_1 0.01fF
C31532 AND2X1_LOC_621/Y AND2X1_LOC_792/Y 0.07fF
C31533 AND2X1_LOC_3/Y OR2X1_LOC_434/A 0.44fF
C31534 OR2X1_LOC_323/A AND2X1_LOC_721/Y 0.00fF
C31535 OR2X1_LOC_743/A OR2X1_LOC_417/A 0.03fF
C31536 OR2X1_LOC_64/Y OR2X1_LOC_246/A 0.03fF
C31537 OR2X1_LOC_696/A AND2X1_LOC_810/B 0.07fF
C31538 AND2X1_LOC_787/A AND2X1_LOC_543/Y 0.03fF
C31539 OR2X1_LOC_121/B AND2X1_LOC_491/a_36_24# 0.01fF
C31540 AND2X1_LOC_672/B OR2X1_LOC_415/A 0.00fF
C31541 AND2X1_LOC_121/a_8_24# OR2X1_LOC_13/B 0.04fF
C31542 OR2X1_LOC_375/A OR2X1_LOC_493/Y 0.03fF
C31543 OR2X1_LOC_97/A OR2X1_LOC_390/a_8_216# 0.01fF
C31544 OR2X1_LOC_650/Y OR2X1_LOC_520/B 0.02fF
C31545 OR2X1_LOC_595/A OR2X1_LOC_767/Y 0.05fF
C31546 OR2X1_LOC_36/Y AND2X1_LOC_463/B 0.03fF
C31547 OR2X1_LOC_696/A AND2X1_LOC_181/Y 0.01fF
C31548 OR2X1_LOC_769/B OR2X1_LOC_769/a_8_216# 0.03fF
C31549 OR2X1_LOC_807/A OR2X1_LOC_580/a_8_216# 0.39fF
C31550 OR2X1_LOC_184/Y OR2X1_LOC_89/A 0.13fF
C31551 OR2X1_LOC_481/A OR2X1_LOC_55/a_8_216# 0.01fF
C31552 OR2X1_LOC_70/Y OR2X1_LOC_426/a_8_216# 0.02fF
C31553 AND2X1_LOC_715/Y AND2X1_LOC_810/B 0.39fF
C31554 OR2X1_LOC_614/a_8_216# AND2X1_LOC_51/Y 0.01fF
C31555 OR2X1_LOC_655/B OR2X1_LOC_750/A 0.01fF
C31556 AND2X1_LOC_31/Y OR2X1_LOC_161/A 0.18fF
C31557 OR2X1_LOC_47/Y OR2X1_LOC_438/a_36_216# 0.03fF
C31558 OR2X1_LOC_64/Y OR2X1_LOC_409/B 0.00fF
C31559 AND2X1_LOC_629/Y AND2X1_LOC_630/a_8_24# 0.03fF
C31560 AND2X1_LOC_91/B OR2X1_LOC_151/A 0.29fF
C31561 AND2X1_LOC_339/Y AND2X1_LOC_351/a_8_24# 0.03fF
C31562 AND2X1_LOC_168/a_8_24# OR2X1_LOC_437/A 0.04fF
C31563 OR2X1_LOC_633/B OR2X1_LOC_84/Y 0.00fF
C31564 OR2X1_LOC_246/A OR2X1_LOC_417/A 0.03fF
C31565 AND2X1_LOC_514/Y AND2X1_LOC_864/a_8_24# 0.04fF
C31566 AND2X1_LOC_381/a_8_24# OR2X1_LOC_68/B 0.01fF
C31567 OR2X1_LOC_3/Y AND2X1_LOC_721/A 0.02fF
C31568 OR2X1_LOC_114/B OR2X1_LOC_140/B 0.01fF
C31569 OR2X1_LOC_186/Y OR2X1_LOC_547/a_8_216# 0.08fF
C31570 OR2X1_LOC_113/Y OR2X1_LOC_844/B 0.02fF
C31571 OR2X1_LOC_92/Y OR2X1_LOC_424/Y -0.01fF
C31572 OR2X1_LOC_26/Y OR2X1_LOC_70/A 0.68fF
C31573 OR2X1_LOC_414/Y AND2X1_LOC_415/a_8_24# 0.00fF
C31574 AND2X1_LOC_25/Y AND2X1_LOC_31/Y 0.06fF
C31575 OR2X1_LOC_70/Y AND2X1_LOC_451/a_8_24# 0.02fF
C31576 OR2X1_LOC_39/A OR2X1_LOC_521/a_8_216# 0.00fF
C31577 OR2X1_LOC_225/a_8_216# OR2X1_LOC_417/A 0.05fF
C31578 OR2X1_LOC_811/A OR2X1_LOC_580/A 0.10fF
C31579 OR2X1_LOC_74/A OR2X1_LOC_86/A 0.00fF
C31580 OR2X1_LOC_405/A OR2X1_LOC_728/A 0.03fF
C31581 AND2X1_LOC_787/A OR2X1_LOC_322/Y 0.03fF
C31582 AND2X1_LOC_437/a_8_24# OR2X1_LOC_168/Y 0.07fF
C31583 OR2X1_LOC_66/A OR2X1_LOC_115/B 0.01fF
C31584 INPUT_1 AND2X1_LOC_270/a_8_24# 0.01fF
C31585 AND2X1_LOC_663/B AND2X1_LOC_620/Y 0.01fF
C31586 OR2X1_LOC_80/Y OR2X1_LOC_80/A 0.00fF
C31587 OR2X1_LOC_140/A OR2X1_LOC_267/Y 0.06fF
C31588 AND2X1_LOC_364/a_8_24# AND2X1_LOC_566/B 0.01fF
C31589 OR2X1_LOC_52/B OR2X1_LOC_72/Y 0.05fF
C31590 OR2X1_LOC_47/Y OR2X1_LOC_54/Y 0.08fF
C31591 OR2X1_LOC_74/A AND2X1_LOC_804/a_36_24# 0.01fF
C31592 AND2X1_LOC_57/Y AND2X1_LOC_41/A 0.06fF
C31593 OR2X1_LOC_663/a_8_216# OR2X1_LOC_113/B 0.01fF
C31594 AND2X1_LOC_535/Y OR2X1_LOC_428/A 0.07fF
C31595 AND2X1_LOC_476/Y OR2X1_LOC_323/Y 0.26fF
C31596 OR2X1_LOC_123/B OR2X1_LOC_598/A 0.02fF
C31597 OR2X1_LOC_797/B OR2X1_LOC_160/Y 0.04fF
C31598 VDD OR2X1_LOC_310/a_8_216# 0.21fF
C31599 AND2X1_LOC_184/a_8_24# AND2X1_LOC_44/Y 0.01fF
C31600 AND2X1_LOC_303/A OR2X1_LOC_437/A 0.01fF
C31601 AND2X1_LOC_566/B OR2X1_LOC_589/A 0.11fF
C31602 OR2X1_LOC_392/B OR2X1_LOC_78/A 0.01fF
C31603 OR2X1_LOC_149/B AND2X1_LOC_41/A 0.18fF
C31604 OR2X1_LOC_158/A AND2X1_LOC_347/B 0.01fF
C31605 OR2X1_LOC_129/a_36_216# OR2X1_LOC_589/A 0.00fF
C31606 OR2X1_LOC_814/A AND2X1_LOC_289/a_8_24# 0.11fF
C31607 OR2X1_LOC_248/a_36_216# OR2X1_LOC_437/A 0.00fF
C31608 AND2X1_LOC_810/A AND2X1_LOC_436/Y 0.01fF
C31609 AND2X1_LOC_22/Y INPUT_0 0.07fF
C31610 OR2X1_LOC_206/a_36_216# AND2X1_LOC_31/Y 0.00fF
C31611 OR2X1_LOC_672/a_8_216# OR2X1_LOC_96/Y 0.40fF
C31612 AND2X1_LOC_64/Y OR2X1_LOC_623/B 0.03fF
C31613 OR2X1_LOC_585/A OR2X1_LOC_385/a_8_216# 0.07fF
C31614 AND2X1_LOC_31/Y AND2X1_LOC_51/Y 1.85fF
C31615 OR2X1_LOC_328/a_8_216# AND2X1_LOC_639/B 0.05fF
C31616 AND2X1_LOC_547/Y AND2X1_LOC_476/Y 0.02fF
C31617 AND2X1_LOC_592/Y AND2X1_LOC_732/B 0.02fF
C31618 OR2X1_LOC_744/A AND2X1_LOC_774/A 0.03fF
C31619 OR2X1_LOC_678/Y AND2X1_LOC_44/Y 0.01fF
C31620 AND2X1_LOC_704/a_8_24# OR2X1_LOC_51/Y 0.01fF
C31621 OR2X1_LOC_676/Y OR2X1_LOC_515/A 0.03fF
C31622 AND2X1_LOC_345/Y OR2X1_LOC_384/Y 0.23fF
C31623 AND2X1_LOC_784/Y VDD 0.40fF
C31624 AND2X1_LOC_392/A AND2X1_LOC_357/A 0.00fF
C31625 AND2X1_LOC_91/B OR2X1_LOC_788/a_8_216# 0.02fF
C31626 AND2X1_LOC_336/a_8_24# OR2X1_LOC_13/B 0.02fF
C31627 AND2X1_LOC_566/B AND2X1_LOC_337/a_8_24# 0.00fF
C31628 OR2X1_LOC_375/A OR2X1_LOC_130/a_8_216# 0.01fF
C31629 OR2X1_LOC_485/A OR2X1_LOC_437/A 0.27fF
C31630 OR2X1_LOC_78/A OR2X1_LOC_113/B 0.02fF
C31631 AND2X1_LOC_707/Y OR2X1_LOC_92/Y 0.20fF
C31632 AND2X1_LOC_70/Y AND2X1_LOC_625/a_8_24# 0.01fF
C31633 OR2X1_LOC_97/A AND2X1_LOC_58/a_8_24# 0.01fF
C31634 AND2X1_LOC_12/Y OR2X1_LOC_140/B 0.03fF
C31635 AND2X1_LOC_7/B OR2X1_LOC_737/A 0.07fF
C31636 AND2X1_LOC_357/B OR2X1_LOC_56/A 0.03fF
C31637 AND2X1_LOC_141/A OR2X1_LOC_12/Y 0.00fF
C31638 AND2X1_LOC_721/a_36_24# OR2X1_LOC_428/A 0.01fF
C31639 OR2X1_LOC_229/a_36_216# AND2X1_LOC_857/Y 0.00fF
C31640 AND2X1_LOC_95/Y AND2X1_LOC_7/B 0.69fF
C31641 OR2X1_LOC_106/Y OR2X1_LOC_39/A 0.00fF
C31642 OR2X1_LOC_64/Y OR2X1_LOC_599/a_8_216# 0.01fF
C31643 AND2X1_LOC_53/Y OR2X1_LOC_779/B 0.34fF
C31644 OR2X1_LOC_811/A AND2X1_LOC_44/Y 0.03fF
C31645 AND2X1_LOC_567/a_36_24# AND2X1_LOC_436/Y 0.00fF
C31646 OR2X1_LOC_160/B AND2X1_LOC_92/Y 0.11fF
C31647 OR2X1_LOC_126/a_36_216# OR2X1_LOC_39/A 0.02fF
C31648 OR2X1_LOC_158/A AND2X1_LOC_116/a_36_24# 0.00fF
C31649 OR2X1_LOC_302/a_36_216# AND2X1_LOC_110/Y 0.00fF
C31650 OR2X1_LOC_633/Y AND2X1_LOC_7/B 0.03fF
C31651 AND2X1_LOC_363/Y OR2X1_LOC_56/A 0.13fF
C31652 OR2X1_LOC_18/Y OR2X1_LOC_18/a_8_216# 0.01fF
C31653 VDD AND2X1_LOC_219/Y 0.78fF
C31654 OR2X1_LOC_516/Y OR2X1_LOC_239/a_8_216# 0.02fF
C31655 AND2X1_LOC_621/Y OR2X1_LOC_816/A 0.06fF
C31656 OR2X1_LOC_223/A OR2X1_LOC_192/a_8_216# 0.13fF
C31657 OR2X1_LOC_97/A OR2X1_LOC_377/A 0.00fF
C31658 OR2X1_LOC_599/A AND2X1_LOC_783/B 0.01fF
C31659 AND2X1_LOC_809/A AND2X1_LOC_802/Y 0.28fF
C31660 OR2X1_LOC_696/A OR2X1_LOC_585/A 0.89fF
C31661 AND2X1_LOC_61/a_36_24# OR2X1_LOC_59/Y 0.00fF
C31662 OR2X1_LOC_243/a_8_216# OR2X1_LOC_71/A 0.01fF
C31663 OR2X1_LOC_161/A OR2X1_LOC_708/a_36_216# 0.00fF
C31664 OR2X1_LOC_44/Y OR2X1_LOC_748/Y 0.02fF
C31665 OR2X1_LOC_97/A AND2X1_LOC_824/B 0.00fF
C31666 OR2X1_LOC_201/a_36_216# AND2X1_LOC_31/Y 0.00fF
C31667 OR2X1_LOC_130/A AND2X1_LOC_224/a_36_24# 0.01fF
C31668 AND2X1_LOC_366/A AND2X1_LOC_367/B 0.23fF
C31669 AND2X1_LOC_624/A AND2X1_LOC_213/B 0.03fF
C31670 OR2X1_LOC_316/Y AND2X1_LOC_786/Y 0.07fF
C31671 AND2X1_LOC_344/a_8_24# AND2X1_LOC_860/A 0.02fF
C31672 OR2X1_LOC_600/A OR2X1_LOC_251/a_36_216# 0.02fF
C31673 OR2X1_LOC_840/A OR2X1_LOC_66/A 0.03fF
C31674 OR2X1_LOC_288/A OR2X1_LOC_366/Y 0.00fF
C31675 AND2X1_LOC_40/Y OR2X1_LOC_676/Y 0.08fF
C31676 OR2X1_LOC_86/A AND2X1_LOC_647/Y 0.00fF
C31677 AND2X1_LOC_576/Y OR2X1_LOC_428/A 0.06fF
C31678 AND2X1_LOC_715/Y OR2X1_LOC_585/A 0.10fF
C31679 OR2X1_LOC_84/A OR2X1_LOC_80/A 0.02fF
C31680 OR2X1_LOC_600/A OR2X1_LOC_46/a_8_216# 0.01fF
C31681 OR2X1_LOC_604/A OR2X1_LOC_281/a_8_216# 0.35fF
C31682 OR2X1_LOC_756/B OR2X1_LOC_168/B 0.00fF
C31683 OR2X1_LOC_649/B AND2X1_LOC_44/Y 0.03fF
C31684 OR2X1_LOC_49/A OR2X1_LOC_97/B 0.11fF
C31685 AND2X1_LOC_353/a_8_24# OR2X1_LOC_619/Y 0.03fF
C31686 OR2X1_LOC_175/Y OR2X1_LOC_574/A 0.15fF
C31687 VDD OR2X1_LOC_610/a_8_216# 0.00fF
C31688 OR2X1_LOC_483/a_36_216# OR2X1_LOC_161/B 0.00fF
C31689 AND2X1_LOC_566/B AND2X1_LOC_365/A 0.00fF
C31690 OR2X1_LOC_645/a_8_216# OR2X1_LOC_788/a_8_216# 0.47fF
C31691 INPUT_1 AND2X1_LOC_750/a_8_24# 0.00fF
C31692 AND2X1_LOC_392/A OR2X1_LOC_18/Y 0.07fF
C31693 OR2X1_LOC_429/a_8_216# D_INPUT_6 0.01fF
C31694 OR2X1_LOC_337/a_8_216# OR2X1_LOC_352/A 0.01fF
C31695 OR2X1_LOC_315/a_8_216# OR2X1_LOC_6/A 0.01fF
C31696 OR2X1_LOC_687/Y OR2X1_LOC_729/a_8_216# 0.05fF
C31697 AND2X1_LOC_349/a_36_24# OR2X1_LOC_12/Y 0.00fF
C31698 OR2X1_LOC_784/a_8_216# AND2X1_LOC_44/Y 0.01fF
C31699 OR2X1_LOC_392/B OR2X1_LOC_392/a_8_216# 0.08fF
C31700 OR2X1_LOC_348/Y AND2X1_LOC_755/a_8_24# 0.01fF
C31701 OR2X1_LOC_61/B OR2X1_LOC_78/B -0.01fF
C31702 OR2X1_LOC_18/Y AND2X1_LOC_807/B 0.04fF
C31703 OR2X1_LOC_668/a_36_216# OR2X1_LOC_244/Y 0.01fF
C31704 AND2X1_LOC_851/a_8_24# AND2X1_LOC_851/A 0.19fF
C31705 OR2X1_LOC_45/B OR2X1_LOC_126/a_8_216# 0.18fF
C31706 AND2X1_LOC_31/Y OR2X1_LOC_551/B 0.72fF
C31707 OR2X1_LOC_235/B OR2X1_LOC_502/A 0.07fF
C31708 OR2X1_LOC_312/Y OR2X1_LOC_373/Y 0.56fF
C31709 OR2X1_LOC_505/Y OR2X1_LOC_39/A 0.09fF
C31710 OR2X1_LOC_127/Y OR2X1_LOC_600/A 0.01fF
C31711 OR2X1_LOC_10/a_8_216# OR2X1_LOC_437/A 0.41fF
C31712 OR2X1_LOC_711/B OR2X1_LOC_468/Y 0.00fF
C31713 AND2X1_LOC_59/Y OR2X1_LOC_776/Y 0.04fF
C31714 OR2X1_LOC_648/A OR2X1_LOC_405/a_8_216# 0.03fF
C31715 AND2X1_LOC_12/Y OR2X1_LOC_851/a_8_216# -0.00fF
C31716 AND2X1_LOC_347/Y AND2X1_LOC_360/a_8_24# 0.11fF
C31717 AND2X1_LOC_702/a_8_24# OR2X1_LOC_56/A 0.05fF
C31718 AND2X1_LOC_41/A OR2X1_LOC_61/a_36_216# 0.02fF
C31719 OR2X1_LOC_54/Y OR2X1_LOC_397/a_8_216# 0.01fF
C31720 AND2X1_LOC_566/B OR2X1_LOC_43/A 0.34fF
C31721 VDD OR2X1_LOC_510/Y 0.18fF
C31722 OR2X1_LOC_51/Y AND2X1_LOC_652/a_8_24# 0.17fF
C31723 OR2X1_LOC_638/a_8_216# OR2X1_LOC_651/B 0.00fF
C31724 OR2X1_LOC_194/B OR2X1_LOC_78/B 0.01fF
C31725 OR2X1_LOC_829/a_8_216# AND2X1_LOC_434/Y 0.01fF
C31726 VDD OR2X1_LOC_456/Y 0.10fF
C31727 AND2X1_LOC_658/A OR2X1_LOC_39/A 0.13fF
C31728 OR2X1_LOC_604/A OR2X1_LOC_6/A 0.05fF
C31729 OR2X1_LOC_600/A OR2X1_LOC_236/a_8_216# -0.00fF
C31730 OR2X1_LOC_323/A AND2X1_LOC_471/a_8_24# 0.01fF
C31731 AND2X1_LOC_596/a_8_24# OR2X1_LOC_44/Y 0.01fF
C31732 OR2X1_LOC_860/a_8_216# OR2X1_LOC_756/B 0.01fF
C31733 OR2X1_LOC_12/Y AND2X1_LOC_651/B 0.00fF
C31734 OR2X1_LOC_592/A OR2X1_LOC_435/A 0.00fF
C31735 OR2X1_LOC_316/Y AND2X1_LOC_218/Y 0.02fF
C31736 AND2X1_LOC_366/A OR2X1_LOC_18/Y 0.01fF
C31737 OR2X1_LOC_158/A OR2X1_LOC_24/Y 0.03fF
C31738 OR2X1_LOC_164/Y OR2X1_LOC_427/A 0.11fF
C31739 OR2X1_LOC_11/Y OR2X1_LOC_12/a_8_216# 0.18fF
C31740 OR2X1_LOC_58/Y OR2X1_LOC_753/A 0.03fF
C31741 OR2X1_LOC_298/a_36_216# AND2X1_LOC_654/Y 0.01fF
C31742 AND2X1_LOC_18/Y OR2X1_LOC_269/B 5.02fF
C31743 AND2X1_LOC_523/Y AND2X1_LOC_455/B 0.01fF
C31744 OR2X1_LOC_656/B OR2X1_LOC_663/A 0.07fF
C31745 AND2X1_LOC_144/a_8_24# OR2X1_LOC_375/A 0.01fF
C31746 OR2X1_LOC_496/Y VDD 0.14fF
C31747 VDD AND2X1_LOC_159/a_8_24# 0.00fF
C31748 AND2X1_LOC_719/Y OR2X1_LOC_74/A 0.01fF
C31749 OR2X1_LOC_557/A OR2X1_LOC_768/a_36_216# 0.00fF
C31750 OR2X1_LOC_236/a_36_216# OR2X1_LOC_56/A 0.00fF
C31751 OR2X1_LOC_831/a_36_216# AND2X1_LOC_92/Y 0.01fF
C31752 OR2X1_LOC_319/B AND2X1_LOC_95/Y 0.13fF
C31753 OR2X1_LOC_329/B AND2X1_LOC_319/A 0.44fF
C31754 VDD OR2X1_LOC_810/A 2.30fF
C31755 OR2X1_LOC_450/A OR2X1_LOC_155/A 0.01fF
C31756 AND2X1_LOC_59/Y OR2X1_LOC_756/B 0.21fF
C31757 OR2X1_LOC_400/A OR2X1_LOC_235/B 0.02fF
C31758 AND2X1_LOC_191/B AND2X1_LOC_580/B 0.03fF
C31759 OR2X1_LOC_426/B AND2X1_LOC_101/B 0.00fF
C31760 OR2X1_LOC_764/Y VDD 0.16fF
C31761 AND2X1_LOC_384/a_8_24# OR2X1_LOC_812/B 0.04fF
C31762 OR2X1_LOC_324/B OR2X1_LOC_468/Y 0.16fF
C31763 AND2X1_LOC_727/a_8_24# AND2X1_LOC_727/A -0.00fF
C31764 OR2X1_LOC_696/A AND2X1_LOC_645/a_8_24# 0.02fF
C31765 OR2X1_LOC_114/Y OR2X1_LOC_632/Y 0.04fF
C31766 OR2X1_LOC_438/Y AND2X1_LOC_807/Y 0.02fF
C31767 VDD AND2X1_LOC_459/a_8_24# -0.00fF
C31768 AND2X1_LOC_865/a_8_24# AND2X1_LOC_807/Y 0.02fF
C31769 AND2X1_LOC_574/Y OR2X1_LOC_95/Y 0.14fF
C31770 AND2X1_LOC_691/a_36_24# OR2X1_LOC_690/A 0.00fF
C31771 VDD AND2X1_LOC_589/a_8_24# 0.00fF
C31772 AND2X1_LOC_658/A OR2X1_LOC_239/a_36_216# 0.02fF
C31773 OR2X1_LOC_219/B AND2X1_LOC_92/Y 5.56fF
C31774 OR2X1_LOC_133/a_8_216# OR2X1_LOC_46/A 0.06fF
C31775 OR2X1_LOC_287/B OR2X1_LOC_402/B 0.01fF
C31776 OR2X1_LOC_137/Y OR2X1_LOC_235/B 0.02fF
C31777 AND2X1_LOC_456/B AND2X1_LOC_806/A 0.06fF
C31778 OR2X1_LOC_805/A OR2X1_LOC_737/A 0.08fF
C31779 OR2X1_LOC_485/A AND2X1_LOC_434/a_36_24# 0.00fF
C31780 OR2X1_LOC_697/Y OR2X1_LOC_52/B 0.12fF
C31781 AND2X1_LOC_719/a_36_24# OR2X1_LOC_59/Y 0.00fF
C31782 AND2X1_LOC_95/Y OR2X1_LOC_407/a_8_216# 0.02fF
C31783 OR2X1_LOC_840/a_36_216# OR2X1_LOC_814/A 0.01fF
C31784 VDD OR2X1_LOC_119/a_8_216# 0.21fF
C31785 OR2X1_LOC_759/A OR2X1_LOC_665/a_8_216# 0.01fF
C31786 AND2X1_LOC_95/Y OR2X1_LOC_805/A 0.10fF
C31787 AND2X1_LOC_142/a_36_24# OR2X1_LOC_87/A 0.01fF
C31788 AND2X1_LOC_732/B AND2X1_LOC_712/B 0.02fF
C31789 AND2X1_LOC_345/Y OR2X1_LOC_91/A 0.04fF
C31790 AND2X1_LOC_59/Y OR2X1_LOC_660/B 0.00fF
C31791 OR2X1_LOC_3/Y AND2X1_LOC_605/Y 0.02fF
C31792 INPUT_5 AND2X1_LOC_21/Y 0.01fF
C31793 AND2X1_LOC_70/a_8_24# AND2X1_LOC_1/Y 0.00fF
C31794 OR2X1_LOC_661/A D_INPUT_0 0.04fF
C31795 OR2X1_LOC_411/A OR2X1_LOC_46/A 0.03fF
C31796 OR2X1_LOC_666/A AND2X1_LOC_849/A 0.03fF
C31797 AND2X1_LOC_658/A OR2X1_LOC_253/a_36_216# 0.02fF
C31798 OR2X1_LOC_36/Y OR2X1_LOC_45/a_8_216# 0.01fF
C31799 AND2X1_LOC_228/Y AND2X1_LOC_302/a_8_24# 0.01fF
C31800 OR2X1_LOC_185/A OR2X1_LOC_151/Y 0.03fF
C31801 AND2X1_LOC_56/B AND2X1_LOC_233/a_8_24# 0.02fF
C31802 OR2X1_LOC_632/A OR2X1_LOC_631/B 0.01fF
C31803 OR2X1_LOC_807/B OR2X1_LOC_269/B 0.01fF
C31804 AND2X1_LOC_116/B OR2X1_LOC_56/A 0.19fF
C31805 OR2X1_LOC_844/Y OR2X1_LOC_632/Y 0.00fF
C31806 OR2X1_LOC_403/A OR2X1_LOC_557/A 0.01fF
C31807 AND2X1_LOC_2/Y AND2X1_LOC_11/a_8_24# 0.01fF
C31808 AND2X1_LOC_16/a_36_24# OR2X1_LOC_155/A 0.00fF
C31809 OR2X1_LOC_326/a_36_216# OR2X1_LOC_121/B 0.00fF
C31810 AND2X1_LOC_59/Y OR2X1_LOC_76/Y 0.08fF
C31811 OR2X1_LOC_205/a_8_216# OR2X1_LOC_375/A 0.01fF
C31812 OR2X1_LOC_358/a_36_216# OR2X1_LOC_358/B 0.03fF
C31813 AND2X1_LOC_452/Y AND2X1_LOC_446/a_8_24# 0.02fF
C31814 OR2X1_LOC_503/A OR2X1_LOC_497/Y 0.79fF
C31815 OR2X1_LOC_240/B OR2X1_LOC_240/A 0.04fF
C31816 OR2X1_LOC_185/A OR2X1_LOC_593/A 0.01fF
C31817 OR2X1_LOC_80/Y OR2X1_LOC_6/A 0.02fF
C31818 OR2X1_LOC_254/a_8_216# OR2X1_LOC_254/A 0.47fF
C31819 AND2X1_LOC_795/Y AND2X1_LOC_785/Y 0.00fF
C31820 VDD AND2X1_LOC_56/a_8_24# -0.00fF
C31821 AND2X1_LOC_572/A AND2X1_LOC_361/A 0.14fF
C31822 AND2X1_LOC_70/Y AND2X1_LOC_53/Y 0.07fF
C31823 OR2X1_LOC_691/Y AND2X1_LOC_761/a_8_24# 0.01fF
C31824 OR2X1_LOC_185/Y OR2X1_LOC_793/A 0.00fF
C31825 AND2X1_LOC_36/Y OR2X1_LOC_366/Y 0.00fF
C31826 OR2X1_LOC_528/Y AND2X1_LOC_663/a_8_24# 0.02fF
C31827 OR2X1_LOC_36/Y AND2X1_LOC_831/a_8_24# 0.01fF
C31828 AND2X1_LOC_95/Y OR2X1_LOC_296/Y 0.03fF
C31829 OR2X1_LOC_36/Y OR2X1_LOC_44/Y 1.12fF
C31830 OR2X1_LOC_91/a_8_216# OR2X1_LOC_44/Y 0.02fF
C31831 OR2X1_LOC_36/Y AND2X1_LOC_288/a_8_24# 0.03fF
C31832 OR2X1_LOC_6/B OR2X1_LOC_473/A 0.16fF
C31833 OR2X1_LOC_47/Y OR2X1_LOC_765/Y 0.03fF
C31834 OR2X1_LOC_532/B OR2X1_LOC_78/A 1.08fF
C31835 OR2X1_LOC_843/B OR2X1_LOC_493/Y 0.18fF
C31836 OR2X1_LOC_252/Y OR2X1_LOC_74/A 0.03fF
C31837 OR2X1_LOC_625/Y AND2X1_LOC_483/a_8_24# 0.01fF
C31838 VDD AND2X1_LOC_851/B 0.58fF
C31839 AND2X1_LOC_553/a_8_24# OR2X1_LOC_47/Y 0.02fF
C31840 AND2X1_LOC_554/B OR2X1_LOC_67/A 0.02fF
C31841 OR2X1_LOC_248/a_36_216# OR2X1_LOC_753/A 0.01fF
C31842 OR2X1_LOC_808/A OR2X1_LOC_814/A 0.01fF
C31843 AND2X1_LOC_665/a_8_24# OR2X1_LOC_78/A 0.09fF
C31844 OR2X1_LOC_328/a_8_216# OR2X1_LOC_31/Y 0.01fF
C31845 OR2X1_LOC_81/a_36_216# OR2X1_LOC_52/B 0.00fF
C31846 OR2X1_LOC_493/Y OR2X1_LOC_549/A 0.10fF
C31847 D_INPUT_0 AND2X1_LOC_820/B 0.04fF
C31848 OR2X1_LOC_96/a_8_216# OR2X1_LOC_56/A 0.02fF
C31849 OR2X1_LOC_736/Y OR2X1_LOC_318/B 1.42fF
C31850 AND2X1_LOC_95/Y OR2X1_LOC_436/a_8_216# 0.01fF
C31851 OR2X1_LOC_458/B OR2X1_LOC_532/B 0.01fF
C31852 AND2X1_LOC_183/a_8_24# OR2X1_LOC_553/A 0.03fF
C31853 AND2X1_LOC_70/Y OR2X1_LOC_223/A 0.70fF
C31854 OR2X1_LOC_820/A OR2X1_LOC_95/Y 0.17fF
C31855 OR2X1_LOC_141/B OR2X1_LOC_267/A 0.30fF
C31856 OR2X1_LOC_485/A AND2X1_LOC_348/Y 0.06fF
C31857 OR2X1_LOC_417/Y AND2X1_LOC_452/Y 0.27fF
C31858 OR2X1_LOC_485/A OR2X1_LOC_753/A 0.11fF
C31859 AND2X1_LOC_192/Y AND2X1_LOC_797/A 0.09fF
C31860 OR2X1_LOC_185/A OR2X1_LOC_19/B 0.03fF
C31861 AND2X1_LOC_399/a_8_24# AND2X1_LOC_42/B 0.01fF
C31862 OR2X1_LOC_7/A AND2X1_LOC_454/A 0.29fF
C31863 OR2X1_LOC_3/Y AND2X1_LOC_361/A 0.07fF
C31864 OR2X1_LOC_787/a_8_216# OR2X1_LOC_318/B 0.48fF
C31865 OR2X1_LOC_675/a_8_216# OR2X1_LOC_719/Y 0.39fF
C31866 AND2X1_LOC_727/A AND2X1_LOC_621/Y 0.07fF
C31867 OR2X1_LOC_680/A AND2X1_LOC_842/B 0.00fF
C31868 AND2X1_LOC_666/a_36_24# OR2X1_LOC_553/A 0.00fF
C31869 AND2X1_LOC_91/B OR2X1_LOC_714/A 0.01fF
C31870 AND2X1_LOC_865/a_8_24# OR2X1_LOC_95/Y 0.02fF
C31871 AND2X1_LOC_544/a_8_24# AND2X1_LOC_675/A 0.20fF
C31872 OR2X1_LOC_299/a_36_216# OR2X1_LOC_7/A 0.02fF
C31873 OR2X1_LOC_306/a_36_216# OR2X1_LOC_311/Y 0.00fF
C31874 AND2X1_LOC_490/a_8_24# AND2X1_LOC_3/Y 0.02fF
C31875 AND2X1_LOC_7/B OR2X1_LOC_269/A 0.15fF
C31876 OR2X1_LOC_675/a_36_216# OR2X1_LOC_269/B 0.02fF
C31877 VDD OR2X1_LOC_595/Y 0.06fF
C31878 OR2X1_LOC_416/Y OR2X1_LOC_265/Y 0.03fF
C31879 OR2X1_LOC_447/Y OR2X1_LOC_784/Y 0.07fF
C31880 OR2X1_LOC_703/A OR2X1_LOC_223/A 0.03fF
C31881 OR2X1_LOC_114/B OR2X1_LOC_675/Y 0.02fF
C31882 AND2X1_LOC_792/Y OR2X1_LOC_59/Y 0.01fF
C31883 AND2X1_LOC_489/Y AND2X1_LOC_554/B 0.01fF
C31884 OR2X1_LOC_552/B OR2X1_LOC_552/A 0.15fF
C31885 D_INPUT_0 OR2X1_LOC_63/a_8_216# 0.02fF
C31886 OR2X1_LOC_756/B OR2X1_LOC_549/Y 0.01fF
C31887 OR2X1_LOC_864/A AND2X1_LOC_51/Y 0.06fF
C31888 AND2X1_LOC_191/Y AND2X1_LOC_475/a_36_24# 0.01fF
C31889 OR2X1_LOC_497/Y OR2X1_LOC_64/Y 0.53fF
C31890 AND2X1_LOC_138/a_36_24# OR2X1_LOC_46/A 0.00fF
C31891 OR2X1_LOC_696/Y OR2X1_LOC_52/B 0.01fF
C31892 OR2X1_LOC_777/a_8_216# OR2X1_LOC_779/B 0.01fF
C31893 AND2X1_LOC_7/B AND2X1_LOC_41/Y 0.03fF
C31894 OR2X1_LOC_427/A AND2X1_LOC_450/Y 0.01fF
C31895 AND2X1_LOC_663/B OR2X1_LOC_585/A 0.08fF
C31896 AND2X1_LOC_702/Y OR2X1_LOC_46/A 0.06fF
C31897 OR2X1_LOC_654/A AND2X1_LOC_689/a_8_24# 0.04fF
C31898 OR2X1_LOC_117/Y OR2X1_LOC_19/B 0.13fF
C31899 AND2X1_LOC_44/Y OR2X1_LOC_777/B 0.05fF
C31900 OR2X1_LOC_516/Y AND2X1_LOC_776/Y 0.12fF
C31901 AND2X1_LOC_721/Y OR2X1_LOC_142/Y 0.03fF
C31902 OR2X1_LOC_95/Y AND2X1_LOC_621/Y 0.03fF
C31903 AND2X1_LOC_785/a_8_24# AND2X1_LOC_785/A 0.01fF
C31904 OR2X1_LOC_151/A OR2X1_LOC_446/B 0.07fF
C31905 OR2X1_LOC_22/Y AND2X1_LOC_637/Y 0.00fF
C31906 INPUT_3 D_INPUT_3 1.09fF
C31907 OR2X1_LOC_97/A OR2X1_LOC_539/B 0.02fF
C31908 AND2X1_LOC_53/Y OR2X1_LOC_193/Y 0.01fF
C31909 OR2X1_LOC_315/Y AND2X1_LOC_851/B 0.04fF
C31910 OR2X1_LOC_696/A AND2X1_LOC_564/B 0.07fF
C31911 OR2X1_LOC_497/Y OR2X1_LOC_417/A 0.15fF
C31912 AND2X1_LOC_539/a_8_24# OR2X1_LOC_7/A 0.06fF
C31913 AND2X1_LOC_36/Y OR2X1_LOC_548/B 0.03fF
C31914 OR2X1_LOC_808/B OR2X1_LOC_318/B 0.03fF
C31915 OR2X1_LOC_846/B AND2X1_LOC_816/a_8_24# 0.21fF
C31916 OR2X1_LOC_557/A OR2X1_LOC_62/B 0.00fF
C31917 OR2X1_LOC_696/A OR2X1_LOC_368/Y 0.03fF
C31918 OR2X1_LOC_134/a_36_216# OR2X1_LOC_134/Y 0.00fF
C31919 OR2X1_LOC_532/B OR2X1_LOC_155/A 0.03fF
C31920 AND2X1_LOC_94/Y OR2X1_LOC_80/A 0.02fF
C31921 OR2X1_LOC_468/a_8_216# OR2X1_LOC_468/Y 0.01fF
C31922 D_INPUT_3 OR2X1_LOC_618/a_36_216# 0.00fF
C31923 OR2X1_LOC_295/Y OR2X1_LOC_258/Y 0.21fF
C31924 AND2X1_LOC_31/a_8_24# AND2X1_LOC_51/Y 0.01fF
C31925 OR2X1_LOC_64/Y AND2X1_LOC_844/a_8_24# 0.01fF
C31926 AND2X1_LOC_598/a_8_24# OR2X1_LOC_47/Y 0.01fF
C31927 OR2X1_LOC_502/A OR2X1_LOC_779/B 1.53fF
C31928 AND2X1_LOC_485/a_8_24# OR2X1_LOC_739/A 0.01fF
C31929 OR2X1_LOC_496/Y OR2X1_LOC_674/Y 0.02fF
C31930 OR2X1_LOC_862/B OR2X1_LOC_561/A 0.10fF
C31931 OR2X1_LOC_10/a_8_216# OR2X1_LOC_753/A 0.01fF
C31932 AND2X1_LOC_12/Y OR2X1_LOC_774/B 0.12fF
C31933 OR2X1_LOC_26/Y OR2X1_LOC_47/Y 3.84fF
C31934 AND2X1_LOC_12/Y AND2X1_LOC_699/a_8_24# 0.01fF
C31935 AND2X1_LOC_564/A AND2X1_LOC_726/a_8_24# 0.06fF
C31936 AND2X1_LOC_22/Y AND2X1_LOC_7/B 0.10fF
C31937 AND2X1_LOC_12/Y OR2X1_LOC_675/Y 0.03fF
C31938 OR2X1_LOC_84/B OR2X1_LOC_84/a_8_216# 0.05fF
C31939 AND2X1_LOC_349/B OR2X1_LOC_47/Y 0.33fF
C31940 OR2X1_LOC_47/Y OR2X1_LOC_89/A 0.17fF
C31941 OR2X1_LOC_691/Y OR2X1_LOC_855/A 0.00fF
C31942 OR2X1_LOC_405/A OR2X1_LOC_68/B 0.02fF
C31943 AND2X1_LOC_401/a_36_24# OR2X1_LOC_80/A 0.01fF
C31944 OR2X1_LOC_154/A OR2X1_LOC_728/B 0.01fF
C31945 AND2X1_LOC_12/Y OR2X1_LOC_557/a_8_216# 0.01fF
C31946 OR2X1_LOC_136/Y AND2X1_LOC_339/B 0.02fF
C31947 OR2X1_LOC_16/A OR2X1_LOC_428/A 0.10fF
C31948 OR2X1_LOC_70/Y AND2X1_LOC_452/a_36_24# 0.00fF
C31949 AND2X1_LOC_64/Y OR2X1_LOC_507/A 0.03fF
C31950 OR2X1_LOC_48/B OR2X1_LOC_589/Y 0.02fF
C31951 OR2X1_LOC_468/Y OR2X1_LOC_568/a_8_216# 0.01fF
C31952 AND2X1_LOC_711/Y AND2X1_LOC_792/Y 0.01fF
C31953 D_INPUT_0 OR2X1_LOC_54/a_36_216# 0.03fF
C31954 OR2X1_LOC_609/A AND2X1_LOC_647/Y 0.01fF
C31955 INPUT_1 OR2X1_LOC_751/A 0.29fF
C31956 OR2X1_LOC_89/A AND2X1_LOC_405/a_36_24# 0.00fF
C31957 OR2X1_LOC_629/A OR2X1_LOC_598/A 0.02fF
C31958 OR2X1_LOC_256/a_8_216# OR2X1_LOC_437/A -0.06fF
C31959 AND2X1_LOC_332/a_8_24# AND2X1_LOC_339/B 0.01fF
C31960 OR2X1_LOC_446/Y AND2X1_LOC_47/Y 0.03fF
C31961 AND2X1_LOC_564/A OR2X1_LOC_679/a_8_216# 0.04fF
C31962 OR2X1_LOC_108/Y OR2X1_LOC_428/A 0.02fF
C31963 OR2X1_LOC_216/A OR2X1_LOC_508/Y 0.06fF
C31964 OR2X1_LOC_70/A OR2X1_LOC_17/Y 0.26fF
C31965 OR2X1_LOC_53/Y OR2X1_LOC_56/A 0.06fF
C31966 AND2X1_LOC_858/B AND2X1_LOC_465/A 0.07fF
C31967 OR2X1_LOC_106/Y AND2X1_LOC_474/A 0.03fF
C31968 AND2X1_LOC_473/Y OR2X1_LOC_59/Y 0.01fF
C31969 OR2X1_LOC_795/a_8_216# OR2X1_LOC_814/A 0.10fF
C31970 OR2X1_LOC_295/a_8_216# AND2X1_LOC_848/A 0.03fF
C31971 AND2X1_LOC_287/B OR2X1_LOC_59/Y 0.03fF
C31972 AND2X1_LOC_215/Y OR2X1_LOC_16/A 0.00fF
C31973 OR2X1_LOC_318/a_8_216# OR2X1_LOC_776/Y 0.02fF
C31974 AND2X1_LOC_64/Y OR2X1_LOC_776/a_8_216# 0.03fF
C31975 OR2X1_LOC_114/B OR2X1_LOC_736/Y 0.01fF
C31976 AND2X1_LOC_42/a_36_24# OR2X1_LOC_80/A 0.00fF
C31977 OR2X1_LOC_816/A OR2X1_LOC_59/Y 0.03fF
C31978 AND2X1_LOC_724/A AND2X1_LOC_447/Y 0.13fF
C31979 AND2X1_LOC_724/Y AND2X1_LOC_705/Y 0.55fF
C31980 AND2X1_LOC_658/A AND2X1_LOC_727/B 0.09fF
C31981 OR2X1_LOC_645/a_36_216# OR2X1_LOC_161/B 0.00fF
C31982 OR2X1_LOC_97/A OR2X1_LOC_78/B 0.03fF
C31983 OR2X1_LOC_56/A AND2X1_LOC_802/Y 0.03fF
C31984 OR2X1_LOC_6/B OR2X1_LOC_786/a_36_216# 0.02fF
C31985 OR2X1_LOC_621/A OR2X1_LOC_621/a_8_216# 0.01fF
C31986 OR2X1_LOC_814/A OR2X1_LOC_374/Y 0.07fF
C31987 OR2X1_LOC_744/A AND2X1_LOC_786/Y 0.07fF
C31988 AND2X1_LOC_719/Y AND2X1_LOC_860/A 0.10fF
C31989 AND2X1_LOC_339/B OR2X1_LOC_51/Y 0.03fF
C31990 AND2X1_LOC_121/a_8_24# OR2X1_LOC_595/A 0.02fF
C31991 OR2X1_LOC_185/Y OR2X1_LOC_576/a_36_216# 0.00fF
C31992 AND2X1_LOC_77/a_8_24# OR2X1_LOC_68/B 0.01fF
C31993 OR2X1_LOC_482/a_8_216# OR2X1_LOC_51/Y 0.15fF
C31994 AND2X1_LOC_64/Y OR2X1_LOC_653/Y 0.43fF
C31995 OR2X1_LOC_715/B VDD 1.93fF
C31996 OR2X1_LOC_6/B OR2X1_LOC_14/a_8_216# 0.03fF
C31997 OR2X1_LOC_495/Y AND2X1_LOC_241/a_8_24# 0.23fF
C31998 OR2X1_LOC_161/A OR2X1_LOC_501/A 0.01fF
C31999 OR2X1_LOC_452/A OR2X1_LOC_452/a_8_216# 0.39fF
C32000 VDD AND2X1_LOC_480/A 0.21fF
C32001 AND2X1_LOC_64/Y OR2X1_LOC_833/B 0.00fF
C32002 OR2X1_LOC_22/Y OR2X1_LOC_72/Y 0.02fF
C32003 AND2X1_LOC_48/A OR2X1_LOC_779/B 0.32fF
C32004 OR2X1_LOC_400/B AND2X1_LOC_36/Y 0.05fF
C32005 AND2X1_LOC_539/Y AND2X1_LOC_801/a_8_24# 0.01fF
C32006 AND2X1_LOC_552/a_8_24# OR2X1_LOC_427/A 0.01fF
C32007 OR2X1_LOC_596/A OR2X1_LOC_715/A 0.02fF
C32008 VDD OR2X1_LOC_784/B -0.00fF
C32009 OR2X1_LOC_491/a_8_216# OR2X1_LOC_59/Y 0.01fF
C32010 OR2X1_LOC_40/Y AND2X1_LOC_570/Y 0.02fF
C32011 OR2X1_LOC_161/A AND2X1_LOC_760/a_8_24# 0.04fF
C32012 AND2X1_LOC_22/Y OR2X1_LOC_318/Y 0.01fF
C32013 AND2X1_LOC_172/a_8_24# AND2X1_LOC_18/Y 0.01fF
C32014 AND2X1_LOC_544/Y AND2X1_LOC_676/a_8_24# 0.07fF
C32015 AND2X1_LOC_564/B AND2X1_LOC_717/a_8_24# 0.02fF
C32016 OR2X1_LOC_6/B AND2X1_LOC_498/a_8_24# 0.02fF
C32017 OR2X1_LOC_575/A AND2X1_LOC_44/Y 0.49fF
C32018 OR2X1_LOC_574/a_8_216# OR2X1_LOC_161/B -0.02fF
C32019 AND2X1_LOC_64/Y OR2X1_LOC_254/B 0.15fF
C32020 OR2X1_LOC_440/B OR2X1_LOC_78/A 0.01fF
C32021 AND2X1_LOC_348/A OR2X1_LOC_12/Y 0.00fF
C32022 OR2X1_LOC_467/A OR2X1_LOC_466/A 0.01fF
C32023 AND2X1_LOC_98/a_36_24# OR2X1_LOC_51/Y 0.00fF
C32024 OR2X1_LOC_709/A OR2X1_LOC_502/A 0.14fF
C32025 OR2X1_LOC_161/A OR2X1_LOC_121/A 0.02fF
C32026 OR2X1_LOC_441/Y AND2X1_LOC_443/a_8_24# 0.01fF
C32027 AND2X1_LOC_40/Y AND2X1_LOC_83/a_8_24# 0.02fF
C32028 OR2X1_LOC_623/B OR2X1_LOC_185/a_8_216# 0.09fF
C32029 AND2X1_LOC_47/Y OR2X1_LOC_228/Y 0.07fF
C32030 OR2X1_LOC_151/A OR2X1_LOC_736/A 0.54fF
C32031 OR2X1_LOC_473/A OR2X1_LOC_598/A 0.75fF
C32032 OR2X1_LOC_51/Y OR2X1_LOC_816/a_8_216# 0.05fF
C32033 OR2X1_LOC_589/A OR2X1_LOC_92/Y 0.12fF
C32034 AND2X1_LOC_564/B AND2X1_LOC_458/Y 0.01fF
C32035 OR2X1_LOC_186/Y OR2X1_LOC_620/Y 0.09fF
C32036 AND2X1_LOC_535/Y AND2X1_LOC_512/Y 0.01fF
C32037 VDD AND2X1_LOC_364/Y 0.29fF
C32038 AND2X1_LOC_301/a_36_24# OR2X1_LOC_59/Y 0.01fF
C32039 AND2X1_LOC_849/A OR2X1_LOC_13/B 0.01fF
C32040 OR2X1_LOC_856/B OR2X1_LOC_856/A 0.14fF
C32041 AND2X1_LOC_22/Y OR2X1_LOC_805/A 0.03fF
C32042 AND2X1_LOC_354/Y AND2X1_LOC_810/B 0.15fF
C32043 OR2X1_LOC_377/A OR2X1_LOC_691/Y 0.02fF
C32044 AND2X1_LOC_95/Y OR2X1_LOC_580/B 0.05fF
C32045 OR2X1_LOC_97/A OR2X1_LOC_375/A 3.27fF
C32046 OR2X1_LOC_132/a_36_216# OR2X1_LOC_132/Y 0.00fF
C32047 OR2X1_LOC_427/A AND2X1_LOC_771/B 0.03fF
C32048 OR2X1_LOC_651/A OR2X1_LOC_198/A 0.01fF
C32049 OR2X1_LOC_3/Y OR2X1_LOC_387/A 0.01fF
C32050 OR2X1_LOC_151/A OR2X1_LOC_631/a_8_216# 0.02fF
C32051 AND2X1_LOC_810/A AND2X1_LOC_655/A 0.05fF
C32052 OR2X1_LOC_676/Y AND2X1_LOC_39/a_8_24# 0.03fF
C32053 OR2X1_LOC_7/A AND2X1_LOC_783/B 0.01fF
C32054 OR2X1_LOC_78/A OR2X1_LOC_78/a_36_216# 0.01fF
C32055 OR2X1_LOC_78/B OR2X1_LOC_78/a_8_216# 0.02fF
C32056 OR2X1_LOC_604/A OR2X1_LOC_485/a_8_216# 0.01fF
C32057 OR2X1_LOC_858/A AND2X1_LOC_41/A 0.02fF
C32058 OR2X1_LOC_188/Y OR2X1_LOC_455/a_8_216# 0.00fF
C32059 AND2X1_LOC_443/Y AND2X1_LOC_444/a_36_24# 0.01fF
C32060 OR2X1_LOC_45/B OR2X1_LOC_36/Y 5.76fF
C32061 OR2X1_LOC_516/Y AND2X1_LOC_830/a_8_24# 0.02fF
C32062 OR2X1_LOC_709/B OR2X1_LOC_738/A 0.03fF
C32063 AND2X1_LOC_40/Y OR2X1_LOC_602/Y 0.07fF
C32064 AND2X1_LOC_580/B AND2X1_LOC_580/a_36_24# 0.01fF
C32065 OR2X1_LOC_614/Y AND2X1_LOC_12/Y 0.03fF
C32066 GATE_366 OR2X1_LOC_759/a_8_216# 0.00fF
C32067 OR2X1_LOC_589/A OR2X1_LOC_65/B 0.02fF
C32068 AND2X1_LOC_840/B AND2X1_LOC_786/Y 0.10fF
C32069 AND2X1_LOC_95/Y OR2X1_LOC_648/B 0.01fF
C32070 AND2X1_LOC_70/Y OR2X1_LOC_502/A 0.32fF
C32071 OR2X1_LOC_54/Y AND2X1_LOC_36/Y 6.20fF
C32072 OR2X1_LOC_711/B OR2X1_LOC_160/A 0.34fF
C32073 VDD OR2X1_LOC_837/B 0.31fF
C32074 AND2X1_LOC_229/a_36_24# OR2X1_LOC_87/A 0.01fF
C32075 AND2X1_LOC_362/B OR2X1_LOC_67/A 0.03fF
C32076 AND2X1_LOC_710/Y OR2X1_LOC_297/a_36_216# 0.00fF
C32077 AND2X1_LOC_721/Y OR2X1_LOC_238/Y 0.06fF
C32078 OR2X1_LOC_185/A AND2X1_LOC_110/Y 0.03fF
C32079 OR2X1_LOC_252/Y AND2X1_LOC_254/a_8_24# 0.10fF
C32080 OR2X1_LOC_91/A AND2X1_LOC_863/a_8_24# 0.02fF
C32081 OR2X1_LOC_538/A OR2X1_LOC_808/B 0.01fF
C32082 OR2X1_LOC_87/A AND2X1_LOC_65/A 0.02fF
C32083 OR2X1_LOC_177/Y OR2X1_LOC_44/Y 0.00fF
C32084 OR2X1_LOC_78/A OR2X1_LOC_734/a_8_216# 0.02fF
C32085 AND2X1_LOC_336/a_8_24# OR2X1_LOC_428/A 0.03fF
C32086 OR2X1_LOC_421/A AND2X1_LOC_436/B 0.36fF
C32087 OR2X1_LOC_315/a_8_216# OR2X1_LOC_44/Y 0.01fF
C32088 AND2X1_LOC_725/a_8_24# AND2X1_LOC_454/Y 0.00fF
C32089 OR2X1_LOC_620/A OR2X1_LOC_550/B 0.02fF
C32090 OR2X1_LOC_205/a_8_216# OR2X1_LOC_549/A 0.04fF
C32091 OR2X1_LOC_447/Y AND2X1_LOC_36/Y 0.01fF
C32092 OR2X1_LOC_151/A AND2X1_LOC_56/B 1.23fF
C32093 AND2X1_LOC_191/B OR2X1_LOC_278/Y 0.03fF
C32094 OR2X1_LOC_160/B OR2X1_LOC_499/a_36_216# 0.02fF
C32095 OR2X1_LOC_252/a_36_216# OR2X1_LOC_627/Y 0.00fF
C32096 GATE_366 AND2X1_LOC_346/a_8_24# 0.02fF
C32097 OR2X1_LOC_814/A OR2X1_LOC_333/A 0.37fF
C32098 AND2X1_LOC_719/Y AND2X1_LOC_287/Y 0.02fF
C32099 OR2X1_LOC_676/Y AND2X1_LOC_43/B 0.19fF
C32100 VDD OR2X1_LOC_215/Y 0.12fF
C32101 OR2X1_LOC_703/A OR2X1_LOC_502/A 0.02fF
C32102 OR2X1_LOC_45/Y OR2X1_LOC_59/Y 0.05fF
C32103 OR2X1_LOC_528/Y AND2X1_LOC_576/Y 0.03fF
C32104 AND2X1_LOC_784/A AND2X1_LOC_182/a_8_24# 0.04fF
C32105 AND2X1_LOC_476/Y AND2X1_LOC_374/Y 0.05fF
C32106 OR2X1_LOC_329/Y OR2X1_LOC_599/A 0.85fF
C32107 AND2X1_LOC_372/a_8_24# OR2X1_LOC_737/A 0.03fF
C32108 AND2X1_LOC_95/Y AND2X1_LOC_103/a_8_24# 0.17fF
C32109 AND2X1_LOC_347/B OR2X1_LOC_748/A 0.61fF
C32110 OR2X1_LOC_427/A AND2X1_LOC_471/Y 1.44fF
C32111 AND2X1_LOC_13/a_8_24# AND2X1_LOC_44/Y 0.02fF
C32112 AND2X1_LOC_19/Y OR2X1_LOC_655/a_36_216# 0.02fF
C32113 AND2X1_LOC_42/B AND2X1_LOC_255/a_8_24# 0.03fF
C32114 OR2X1_LOC_70/Y OR2X1_LOC_79/Y 0.02fF
C32115 OR2X1_LOC_307/A OR2X1_LOC_269/B 0.01fF
C32116 AND2X1_LOC_476/Y OR2X1_LOC_52/B 0.02fF
C32117 AND2X1_LOC_843/a_8_24# OR2X1_LOC_59/Y 0.01fF
C32118 OR2X1_LOC_667/Y AND2X1_LOC_456/B 0.04fF
C32119 OR2X1_LOC_604/A OR2X1_LOC_44/Y 0.21fF
C32120 OR2X1_LOC_756/B OR2X1_LOC_794/A 0.01fF
C32121 OR2X1_LOC_244/Y OR2X1_LOC_575/a_8_216# 0.01fF
C32122 OR2X1_LOC_11/Y OR2X1_LOC_380/a_8_216# 0.01fF
C32123 OR2X1_LOC_680/A AND2X1_LOC_188/a_8_24# 0.07fF
C32124 OR2X1_LOC_721/Y OR2X1_LOC_475/B 0.00fF
C32125 OR2X1_LOC_802/Y OR2X1_LOC_66/A 0.14fF
C32126 AND2X1_LOC_22/Y OR2X1_LOC_436/a_8_216# 0.00fF
C32127 OR2X1_LOC_319/B OR2X1_LOC_854/a_36_216# 0.01fF
C32128 OR2X1_LOC_51/Y AND2X1_LOC_859/a_8_24# 0.00fF
C32129 AND2X1_LOC_807/Y OR2X1_LOC_59/Y 0.13fF
C32130 OR2X1_LOC_235/B AND2X1_LOC_104/a_8_24# 0.01fF
C32131 OR2X1_LOC_160/A OR2X1_LOC_324/B 0.10fF
C32132 OR2X1_LOC_176/a_36_216# OR2X1_LOC_417/Y 0.00fF
C32133 OR2X1_LOC_863/a_8_216# OR2X1_LOC_66/A 0.01fF
C32134 OR2X1_LOC_482/Y OR2X1_LOC_238/Y 0.00fF
C32135 OR2X1_LOC_318/a_36_216# OR2X1_LOC_479/Y 0.00fF
C32136 AND2X1_LOC_710/a_8_24# OR2X1_LOC_59/Y 0.02fF
C32137 OR2X1_LOC_468/Y OR2X1_LOC_66/A 0.03fF
C32138 AND2X1_LOC_705/a_8_24# OR2X1_LOC_36/Y 0.02fF
C32139 OR2X1_LOC_160/A OR2X1_LOC_662/a_8_216# 0.01fF
C32140 OR2X1_LOC_154/A AND2X1_LOC_310/a_8_24# 0.01fF
C32141 OR2X1_LOC_216/a_8_216# AND2X1_LOC_65/A 0.01fF
C32142 OR2X1_LOC_254/a_8_216# OR2X1_LOC_161/B 0.04fF
C32143 AND2X1_LOC_362/B AND2X1_LOC_489/Y 0.03fF
C32144 AND2X1_LOC_387/B OR2X1_LOC_596/A 4.20fF
C32145 OR2X1_LOC_6/B OR2X1_LOC_287/B 0.02fF
C32146 AND2X1_LOC_653/a_8_24# AND2X1_LOC_436/Y 0.01fF
C32147 AND2X1_LOC_385/a_8_24# OR2X1_LOC_66/A 0.05fF
C32148 OR2X1_LOC_541/A OR2X1_LOC_375/A 0.03fF
C32149 AND2X1_LOC_547/Y AND2X1_LOC_474/Y 0.00fF
C32150 AND2X1_LOC_40/Y OR2X1_LOC_811/a_8_216# 0.01fF
C32151 AND2X1_LOC_544/a_36_24# OR2X1_LOC_427/A 0.01fF
C32152 OR2X1_LOC_814/A OR2X1_LOC_392/B 0.03fF
C32153 OR2X1_LOC_185/A AND2X1_LOC_126/a_36_24# 0.01fF
C32154 AND2X1_LOC_732/B OR2X1_LOC_89/A 0.00fF
C32155 AND2X1_LOC_757/a_36_24# OR2X1_LOC_555/B 0.00fF
C32156 OR2X1_LOC_858/A OR2X1_LOC_631/B 0.03fF
C32157 AND2X1_LOC_563/A OR2X1_LOC_529/Y 0.81fF
C32158 AND2X1_LOC_12/Y OR2X1_LOC_808/B 0.20fF
C32159 AND2X1_LOC_128/a_8_24# OR2X1_LOC_428/A 0.02fF
C32160 OR2X1_LOC_631/a_36_216# OR2X1_LOC_575/A 0.00fF
C32161 AND2X1_LOC_302/a_8_24# AND2X1_LOC_857/Y 0.01fF
C32162 AND2X1_LOC_570/Y OR2X1_LOC_7/A 0.01fF
C32163 OR2X1_LOC_622/A AND2X1_LOC_42/B 0.20fF
C32164 AND2X1_LOC_841/B OR2X1_LOC_619/Y 0.07fF
C32165 OR2X1_LOC_427/A AND2X1_LOC_450/a_36_24# 0.00fF
C32166 OR2X1_LOC_643/a_8_216# AND2X1_LOC_92/Y 0.04fF
C32167 OR2X1_LOC_205/Y OR2X1_LOC_508/Y 0.03fF
C32168 OR2X1_LOC_743/A AND2X1_LOC_454/a_8_24# 0.01fF
C32169 OR2X1_LOC_675/a_8_216# OR2X1_LOC_66/A 0.01fF
C32170 OR2X1_LOC_763/Y OR2X1_LOC_744/A 0.09fF
C32171 VDD AND2X1_LOC_196/a_8_24# -0.00fF
C32172 AND2X1_LOC_212/A AND2X1_LOC_514/Y 0.03fF
C32173 AND2X1_LOC_489/Y AND2X1_LOC_558/a_36_24# 0.00fF
C32174 OR2X1_LOC_6/B OR2X1_LOC_825/Y 0.03fF
C32175 AND2X1_LOC_76/Y OR2X1_LOC_595/a_8_216# 0.01fF
C32176 OR2X1_LOC_784/Y OR2X1_LOC_161/A 0.07fF
C32177 OR2X1_LOC_160/A AND2X1_LOC_314/a_8_24# 0.01fF
C32178 OR2X1_LOC_364/A OR2X1_LOC_785/B 0.00fF
C32179 OR2X1_LOC_814/A OR2X1_LOC_113/B 0.04fF
C32180 OR2X1_LOC_235/B AND2X1_LOC_3/Y 0.03fF
C32181 OR2X1_LOC_185/Y OR2X1_LOC_785/B 0.03fF
C32182 AND2X1_LOC_848/A AND2X1_LOC_793/a_36_24# 0.01fF
C32183 OR2X1_LOC_31/Y AND2X1_LOC_786/Y 0.16fF
C32184 OR2X1_LOC_672/a_36_216# OR2X1_LOC_46/A 0.00fF
C32185 OR2X1_LOC_43/A OR2X1_LOC_92/Y 0.13fF
C32186 OR2X1_LOC_31/Y OR2X1_LOC_323/a_8_216# 0.01fF
C32187 OR2X1_LOC_185/Y OR2X1_LOC_861/a_8_216# 0.01fF
C32188 AND2X1_LOC_549/a_36_24# OR2X1_LOC_74/A 0.01fF
C32189 AND2X1_LOC_17/Y OR2X1_LOC_502/A 0.29fF
C32190 OR2X1_LOC_185/A OR2X1_LOC_664/Y 0.01fF
C32191 OR2X1_LOC_305/a_8_216# OR2X1_LOC_48/B 0.01fF
C32192 OR2X1_LOC_677/a_8_216# OR2X1_LOC_74/A 0.03fF
C32193 AND2X1_LOC_506/a_36_24# OR2X1_LOC_74/A 0.01fF
C32194 OR2X1_LOC_100/a_36_216# AND2X1_LOC_81/B 0.00fF
C32195 AND2X1_LOC_134/a_8_24# OR2X1_LOC_66/A 0.01fF
C32196 AND2X1_LOC_720/a_8_24# OR2X1_LOC_26/Y 0.02fF
C32197 OR2X1_LOC_375/A AND2X1_LOC_282/a_8_24# 0.11fF
C32198 AND2X1_LOC_250/a_8_24# OR2X1_LOC_843/B 0.20fF
C32199 OR2X1_LOC_462/B AND2X1_LOC_43/B 0.03fF
C32200 VDD AND2X1_LOC_519/a_8_24# 0.00fF
C32201 OR2X1_LOC_256/a_8_216# OR2X1_LOC_753/A -0.03fF
C32202 OR2X1_LOC_40/Y OR2X1_LOC_813/A 0.00fF
C32203 OR2X1_LOC_43/A AND2X1_LOC_801/a_36_24# 0.00fF
C32204 OR2X1_LOC_36/Y AND2X1_LOC_435/a_8_24# 0.01fF
C32205 AND2X1_LOC_70/Y AND2X1_LOC_48/A 0.17fF
C32206 OR2X1_LOC_653/a_8_216# OR2X1_LOC_502/A 0.05fF
C32207 OR2X1_LOC_680/A AND2X1_LOC_186/a_36_24# 0.00fF
C32208 OR2X1_LOC_703/a_8_216# OR2X1_LOC_365/B 0.39fF
C32209 OR2X1_LOC_154/A AND2X1_LOC_81/B 0.01fF
C32210 OR2X1_LOC_167/a_8_216# OR2X1_LOC_47/Y 0.01fF
C32211 OR2X1_LOC_18/Y AND2X1_LOC_458/a_8_24# 0.02fF
C32212 AND2X1_LOC_727/A OR2X1_LOC_59/Y 0.03fF
C32213 OR2X1_LOC_43/A OR2X1_LOC_65/B 0.03fF
C32214 OR2X1_LOC_599/A AND2X1_LOC_435/a_36_24# 0.00fF
C32215 OR2X1_LOC_36/Y OR2X1_LOC_767/a_8_216# 0.08fF
C32216 OR2X1_LOC_154/A OR2X1_LOC_358/B 0.00fF
C32217 AND2X1_LOC_479/Y AND2X1_LOC_479/a_8_24# 0.02fF
C32218 OR2X1_LOC_109/Y OR2X1_LOC_312/Y 0.41fF
C32219 AND2X1_LOC_720/a_8_24# OR2X1_LOC_89/A 0.03fF
C32220 AND2X1_LOC_347/Y AND2X1_LOC_663/B 0.04fF
C32221 OR2X1_LOC_595/a_8_216# OR2X1_LOC_52/B 0.02fF
C32222 AND2X1_LOC_349/B OR2X1_LOC_625/Y 1.00fF
C32223 OR2X1_LOC_185/Y OR2X1_LOC_687/Y 0.01fF
C32224 OR2X1_LOC_625/Y OR2X1_LOC_89/A 0.09fF
C32225 OR2X1_LOC_547/B OR2X1_LOC_620/B 0.01fF
C32226 INPUT_1 OR2X1_LOC_56/A 0.21fF
C32227 OR2X1_LOC_45/B OR2X1_LOC_419/Y 0.06fF
C32228 AND2X1_LOC_552/A OR2X1_LOC_47/Y 0.08fF
C32229 OR2X1_LOC_487/a_8_216# AND2X1_LOC_573/A 0.03fF
C32230 OR2X1_LOC_819/a_8_216# INPUT_1 0.02fF
C32231 OR2X1_LOC_725/B OR2X1_LOC_705/Y 0.02fF
C32232 OR2X1_LOC_45/Y OR2X1_LOC_70/Y 0.32fF
C32233 AND2X1_LOC_554/Y AND2X1_LOC_554/B 0.02fF
C32234 VDD AND2X1_LOC_479/Y 0.09fF
C32235 AND2X1_LOC_190/a_36_24# OR2X1_LOC_417/A 0.01fF
C32236 OR2X1_LOC_47/Y AND2X1_LOC_194/Y 0.14fF
C32237 OR2X1_LOC_92/Y AND2X1_LOC_685/a_8_24# 0.35fF
C32238 AND2X1_LOC_729/Y OR2X1_LOC_485/A 0.04fF
C32239 AND2X1_LOC_836/a_36_24# OR2X1_LOC_6/A 0.00fF
C32240 OR2X1_LOC_743/A AND2X1_LOC_449/Y 0.01fF
C32241 OR2X1_LOC_287/B OR2X1_LOC_579/B 0.14fF
C32242 AND2X1_LOC_72/B OR2X1_LOC_346/A 0.01fF
C32243 OR2X1_LOC_643/a_36_216# OR2X1_LOC_222/A 0.00fF
C32244 OR2X1_LOC_137/a_8_216# OR2X1_LOC_532/B 0.12fF
C32245 AND2X1_LOC_711/Y AND2X1_LOC_807/Y 0.03fF
C32246 OR2X1_LOC_95/Y OR2X1_LOC_59/Y 0.09fF
C32247 VDD OR2X1_LOC_619/a_8_216# 0.21fF
C32248 OR2X1_LOC_351/B AND2X1_LOC_289/a_8_24# 0.01fF
C32249 OR2X1_LOC_109/a_8_216# OR2X1_LOC_64/Y 0.13fF
C32250 OR2X1_LOC_141/B OR2X1_LOC_267/a_8_216# 0.40fF
C32251 OR2X1_LOC_696/A OR2X1_LOC_437/A 0.41fF
C32252 OR2X1_LOC_70/Y AND2X1_LOC_807/Y 0.02fF
C32253 VDD OR2X1_LOC_409/Y 0.04fF
C32254 OR2X1_LOC_690/A OR2X1_LOC_24/a_8_216# 0.11fF
C32255 OR2X1_LOC_70/Y OR2X1_LOC_427/a_8_216# 0.03fF
C32256 OR2X1_LOC_756/B OR2X1_LOC_544/A 0.01fF
C32257 OR2X1_LOC_673/Y AND2X1_LOC_38/a_8_24# 0.02fF
C32258 AND2X1_LOC_42/B OR2X1_LOC_204/Y 0.97fF
C32259 AND2X1_LOC_51/Y OR2X1_LOC_738/A 0.04fF
C32260 AND2X1_LOC_59/Y OR2X1_LOC_719/A 0.01fF
C32261 OR2X1_LOC_865/B OR2X1_LOC_846/A 1.16fF
C32262 AND2X1_LOC_784/A OR2X1_LOC_485/A 0.07fF
C32263 AND2X1_LOC_537/Y OR2X1_LOC_48/B 0.03fF
C32264 AND2X1_LOC_660/A AND2X1_LOC_219/Y 0.07fF
C32265 AND2X1_LOC_578/A AND2X1_LOC_840/B 0.01fF
C32266 OR2X1_LOC_744/A AND2X1_LOC_114/Y 0.12fF
C32267 OR2X1_LOC_310/Y AND2X1_LOC_318/Y 0.06fF
C32268 OR2X1_LOC_3/Y AND2X1_LOC_852/Y 0.03fF
C32269 OR2X1_LOC_40/Y OR2X1_LOC_406/A 0.04fF
C32270 OR2X1_LOC_160/B OR2X1_LOC_339/Y 0.12fF
C32271 OR2X1_LOC_309/a_8_216# AND2X1_LOC_222/Y 0.01fF
C32272 AND2X1_LOC_383/a_8_24# OR2X1_LOC_437/A 0.02fF
C32273 OR2X1_LOC_233/a_36_216# OR2X1_LOC_585/A 0.00fF
C32274 AND2X1_LOC_165/a_8_24# OR2X1_LOC_506/A 0.07fF
C32275 OR2X1_LOC_529/Y AND2X1_LOC_717/B 0.03fF
C32276 OR2X1_LOC_377/A OR2X1_LOC_750/a_8_216# 0.03fF
C32277 AND2X1_LOC_113/a_8_24# AND2X1_LOC_227/Y 0.01fF
C32278 AND2X1_LOC_719/Y AND2X1_LOC_562/Y 0.10fF
C32279 AND2X1_LOC_259/Y OR2X1_LOC_258/Y 0.01fF
C32280 OR2X1_LOC_154/A OR2X1_LOC_196/B 0.34fF
C32281 D_INPUT_3 AND2X1_LOC_839/a_8_24# 0.01fF
C32282 OR2X1_LOC_663/A OR2X1_LOC_786/Y 0.03fF
C32283 OR2X1_LOC_246/Y OR2X1_LOC_54/Y 0.00fF
C32284 AND2X1_LOC_12/Y AND2X1_LOC_692/a_36_24# 0.00fF
C32285 OR2X1_LOC_137/Y OR2X1_LOC_404/Y -0.00fF
C32286 OR2X1_LOC_821/Y OR2X1_LOC_71/A 0.35fF
C32287 AND2X1_LOC_44/Y OR2X1_LOC_735/B 0.01fF
C32288 VDD OR2X1_LOC_398/Y 0.09fF
C32289 AND2X1_LOC_48/A OR2X1_LOC_193/Y 0.01fF
C32290 OR2X1_LOC_504/Y AND2X1_LOC_807/Y 0.10fF
C32291 OR2X1_LOC_446/Y AND2X1_LOC_695/a_8_24# 0.01fF
C32292 OR2X1_LOC_175/Y OR2X1_LOC_539/B 0.01fF
C32293 OR2X1_LOC_605/B OR2X1_LOC_605/a_8_216# 0.05fF
C32294 OR2X1_LOC_743/A OR2X1_LOC_829/Y 0.01fF
C32295 AND2X1_LOC_99/a_8_24# OR2X1_LOC_813/Y 0.01fF
C32296 AND2X1_LOC_56/B INPUT_1 2.51fF
C32297 AND2X1_LOC_12/Y OR2X1_LOC_218/Y 0.02fF
C32298 OR2X1_LOC_7/a_8_216# OR2X1_LOC_690/A 0.14fF
C32299 OR2X1_LOC_22/A OR2X1_LOC_22/a_8_216# 0.08fF
C32300 OR2X1_LOC_499/B OR2X1_LOC_493/Y 0.01fF
C32301 AND2X1_LOC_557/Y OR2X1_LOC_71/Y 0.01fF
C32302 OR2X1_LOC_526/Y OR2X1_LOC_526/a_36_216# 0.00fF
C32303 OR2X1_LOC_437/a_8_216# OR2X1_LOC_48/B 0.18fF
C32304 OR2X1_LOC_497/Y OR2X1_LOC_226/a_8_216# 0.03fF
C32305 OR2X1_LOC_744/A OR2X1_LOC_88/a_8_216# 0.01fF
C32306 OR2X1_LOC_385/Y AND2X1_LOC_537/Y 0.00fF
C32307 OR2X1_LOC_473/A OR2X1_LOC_506/A 0.02fF
C32308 AND2X1_LOC_8/Y INPUT_1 0.04fF
C32309 OR2X1_LOC_808/A OR2X1_LOC_318/B 0.04fF
C32310 AND2X1_LOC_835/a_8_24# OR2X1_LOC_753/A 0.02fF
C32311 AND2X1_LOC_43/B OR2X1_LOC_200/Y 0.04fF
C32312 AND2X1_LOC_19/Y OR2X1_LOC_68/B 0.02fF
C32313 OR2X1_LOC_62/A OR2X1_LOC_94/a_8_216# 0.18fF
C32314 OR2X1_LOC_287/B OR2X1_LOC_287/a_36_216# 0.03fF
C32315 AND2X1_LOC_41/A AND2X1_LOC_31/Y 0.10fF
C32316 OR2X1_LOC_70/Y AND2X1_LOC_727/A 0.03fF
C32317 OR2X1_LOC_95/Y OR2X1_LOC_820/B 0.04fF
C32318 OR2X1_LOC_796/B OR2X1_LOC_796/a_8_216# 0.39fF
C32319 OR2X1_LOC_709/B AND2X1_LOC_36/Y 0.18fF
C32320 AND2X1_LOC_640/Y D_INPUT_0 0.01fF
C32321 AND2X1_LOC_12/Y AND2X1_LOC_289/a_8_24# 0.01fF
C32322 AND2X1_LOC_386/a_8_24# AND2X1_LOC_47/Y 0.01fF
C32323 AND2X1_LOC_72/B OR2X1_LOC_161/A 1.29fF
C32324 D_INPUT_3 AND2X1_LOC_839/B 0.01fF
C32325 OR2X1_LOC_185/Y OR2X1_LOC_786/Y 0.11fF
C32326 AND2X1_LOC_316/a_8_24# OR2X1_LOC_68/B 0.02fF
C32327 OR2X1_LOC_91/A OR2X1_LOC_384/Y 0.02fF
C32328 OR2X1_LOC_161/A OR2X1_LOC_451/B 0.03fF
C32329 OR2X1_LOC_47/Y OR2X1_LOC_246/a_8_216# 0.01fF
C32330 AND2X1_LOC_804/Y AND2X1_LOC_222/Y 0.01fF
C32331 AND2X1_LOC_514/Y AND2X1_LOC_727/A 0.02fF
C32332 AND2X1_LOC_432/a_8_24# OR2X1_LOC_785/B 0.23fF
C32333 OR2X1_LOC_231/A OR2X1_LOC_641/B 0.26fF
C32334 AND2X1_LOC_578/A OR2X1_LOC_31/Y 0.06fF
C32335 AND2X1_LOC_633/Y OR2X1_LOC_416/Y 0.02fF
C32336 AND2X1_LOC_465/a_36_24# OR2X1_LOC_95/Y 0.01fF
C32337 AND2X1_LOC_31/Y OR2X1_LOC_733/a_36_216# 0.00fF
C32338 OR2X1_LOC_70/Y OR2X1_LOC_95/Y 0.44fF
C32339 OR2X1_LOC_644/a_8_216# OR2X1_LOC_19/B 0.06fF
C32340 OR2X1_LOC_70/Y AND2X1_LOC_440/a_8_24# 0.03fF
C32341 OR2X1_LOC_121/a_8_216# OR2X1_LOC_121/A 0.08fF
C32342 AND2X1_LOC_59/Y OR2X1_LOC_675/Y 0.01fF
C32343 OR2X1_LOC_114/B OR2X1_LOC_500/a_8_216# 0.01fF
C32344 OR2X1_LOC_62/B OR2X1_LOC_46/A 0.23fF
C32345 OR2X1_LOC_383/Y AND2X1_LOC_494/a_8_24# 0.00fF
C32346 D_INPUT_0 OR2X1_LOC_416/Y 0.03fF
C32347 AND2X1_LOC_543/Y OR2X1_LOC_322/a_36_216# 0.00fF
C32348 VDD AND2X1_LOC_619/a_8_24# -0.00fF
C32349 OR2X1_LOC_340/Y OR2X1_LOC_641/B 0.02fF
C32350 OR2X1_LOC_341/Y OR2X1_LOC_228/Y 0.03fF
C32351 OR2X1_LOC_269/B AND2X1_LOC_428/a_8_24# 0.00fF
C32352 OR2X1_LOC_480/a_8_216# OR2X1_LOC_161/B 0.02fF
C32353 OR2X1_LOC_662/A AND2X1_LOC_31/Y 0.00fF
C32354 OR2X1_LOC_269/B OR2X1_LOC_512/a_8_216# 0.12fF
C32355 OR2X1_LOC_39/A OR2X1_LOC_72/Y 0.00fF
C32356 OR2X1_LOC_47/Y OR2X1_LOC_17/Y 0.01fF
C32357 AND2X1_LOC_468/B OR2X1_LOC_533/A 0.09fF
C32358 OR2X1_LOC_130/A OR2X1_LOC_641/B 0.00fF
C32359 AND2X1_LOC_44/Y OR2X1_LOC_161/B 0.70fF
C32360 AND2X1_LOC_554/a_36_24# OR2X1_LOC_595/A 0.01fF
C32361 D_INPUT_0 AND2X1_LOC_667/a_8_24# 0.02fF
C32362 AND2X1_LOC_514/Y OR2X1_LOC_95/Y 0.19fF
C32363 AND2X1_LOC_464/A AND2X1_LOC_786/Y 0.01fF
C32364 OR2X1_LOC_219/B OR2X1_LOC_339/Y 0.03fF
C32365 OR2X1_LOC_555/a_8_216# OR2X1_LOC_562/B -0.00fF
C32366 OR2X1_LOC_11/Y OR2X1_LOC_588/a_36_216# 0.00fF
C32367 OR2X1_LOC_532/B OR2X1_LOC_814/A 0.13fF
C32368 AND2X1_LOC_217/Y OR2X1_LOC_134/Y 0.03fF
C32369 AND2X1_LOC_81/B OR2X1_LOC_560/A 0.03fF
C32370 OR2X1_LOC_45/B OR2X1_LOC_315/a_8_216# 0.01fF
C32371 OR2X1_LOC_538/A OR2X1_LOC_703/Y 0.00fF
C32372 AND2X1_LOC_543/Y OR2X1_LOC_600/A 0.01fF
C32373 VDD OR2X1_LOC_338/B 0.00fF
C32374 OR2X1_LOC_812/B OR2X1_LOC_558/a_8_216# 0.02fF
C32375 AND2X1_LOC_649/B OR2X1_LOC_13/B 0.07fF
C32376 OR2X1_LOC_208/A OR2X1_LOC_35/Y 0.00fF
C32377 AND2X1_LOC_22/Y OR2X1_LOC_648/B 0.05fF
C32378 OR2X1_LOC_665/a_8_216# AND2X1_LOC_620/Y 0.05fF
C32379 OR2X1_LOC_446/Y OR2X1_LOC_780/A 0.00fF
C32380 AND2X1_LOC_565/B AND2X1_LOC_564/B 0.14fF
C32381 OR2X1_LOC_375/A OR2X1_LOC_193/a_8_216# 0.01fF
C32382 OR2X1_LOC_504/Y OR2X1_LOC_95/Y 0.03fF
C32383 OR2X1_LOC_518/Y OR2X1_LOC_91/A 0.03fF
C32384 AND2X1_LOC_61/Y AND2X1_LOC_201/Y 0.22fF
C32385 OR2X1_LOC_45/B OR2X1_LOC_604/A 0.06fF
C32386 OR2X1_LOC_814/A OR2X1_LOC_343/B 0.17fF
C32387 OR2X1_LOC_778/Y OR2X1_LOC_724/A 0.10fF
C32388 AND2X1_LOC_3/Y AND2X1_LOC_430/B 0.00fF
C32389 OR2X1_LOC_688/a_8_216# AND2X1_LOC_31/Y 0.11fF
C32390 OR2X1_LOC_505/a_8_216# OR2X1_LOC_40/Y 0.01fF
C32391 OR2X1_LOC_589/A AND2X1_LOC_729/a_8_24# 0.02fF
C32392 AND2X1_LOC_231/Y OR2X1_LOC_600/A 0.07fF
C32393 OR2X1_LOC_436/Y AND2X1_LOC_47/Y 0.03fF
C32394 D_INPUT_3 AND2X1_LOC_28/a_8_24# 0.01fF
C32395 AND2X1_LOC_3/Y OR2X1_LOC_779/B 0.45fF
C32396 AND2X1_LOC_51/Y OR2X1_LOC_451/B 0.01fF
C32397 OR2X1_LOC_392/B OR2X1_LOC_244/Y 0.81fF
C32398 OR2X1_LOC_741/Y AND2X1_LOC_7/B 0.03fF
C32399 AND2X1_LOC_658/B OR2X1_LOC_816/A 0.01fF
C32400 OR2X1_LOC_322/a_36_216# OR2X1_LOC_322/Y 0.01fF
C32401 AND2X1_LOC_841/a_8_24# OR2X1_LOC_31/Y 0.01fF
C32402 AND2X1_LOC_773/Y VDD 1.46fF
C32403 OR2X1_LOC_485/A OR2X1_LOC_172/Y 0.01fF
C32404 AND2X1_LOC_301/a_8_24# AND2X1_LOC_786/Y 0.02fF
C32405 AND2X1_LOC_741/Y VDD 0.29fF
C32406 OR2X1_LOC_175/Y OR2X1_LOC_78/B 0.11fF
C32407 AND2X1_LOC_543/Y AND2X1_LOC_543/a_8_24# 0.01fF
C32408 OR2X1_LOC_240/B AND2X1_LOC_36/Y 0.05fF
C32409 VDD OR2X1_LOC_35/A 0.00fF
C32410 OR2X1_LOC_696/A OR2X1_LOC_761/Y 0.02fF
C32411 AND2X1_LOC_544/Y AND2X1_LOC_734/Y 0.14fF
C32412 OR2X1_LOC_604/A OR2X1_LOC_382/A 0.06fF
C32413 OR2X1_LOC_161/A AND2X1_LOC_36/Y 1.02fF
C32414 AND2X1_LOC_359/a_8_24# OR2X1_LOC_437/A 0.01fF
C32415 OR2X1_LOC_184/Y OR2X1_LOC_95/Y 0.02fF
C32416 OR2X1_LOC_78/B AND2X1_LOC_417/a_8_24# 0.01fF
C32417 OR2X1_LOC_318/A AND2X1_LOC_92/Y 0.02fF
C32418 OR2X1_LOC_691/Y OR2X1_LOC_78/B 0.03fF
C32419 OR2X1_LOC_624/A AND2X1_LOC_239/a_36_24# 0.06fF
C32420 OR2X1_LOC_835/Y OR2X1_LOC_598/A 0.04fF
C32421 AND2X1_LOC_64/Y AND2X1_LOC_321/a_8_24# 0.01fF
C32422 OR2X1_LOC_276/B OR2X1_LOC_270/Y 0.10fF
C32423 OR2X1_LOC_244/Y OR2X1_LOC_113/B 0.02fF
C32424 OR2X1_LOC_6/B OR2X1_LOC_160/B 0.14fF
C32425 OR2X1_LOC_524/Y AND2X1_LOC_213/B 0.03fF
C32426 AND2X1_LOC_454/A OR2X1_LOC_424/Y -0.00fF
C32427 OR2X1_LOC_575/A OR2X1_LOC_554/a_8_216# 0.03fF
C32428 OR2X1_LOC_139/A OR2X1_LOC_244/a_8_216# 0.03fF
C32429 AND2X1_LOC_25/Y AND2X1_LOC_36/Y 0.01fF
C32430 OR2X1_LOC_18/Y OR2X1_LOC_171/a_8_216# 0.01fF
C32431 VDD AND2X1_LOC_243/Y 1.16fF
C32432 OR2X1_LOC_111/a_8_216# OR2X1_LOC_109/Y 0.01fF
C32433 VDD OR2X1_LOC_552/B -0.00fF
C32434 AND2X1_LOC_715/Y OR2X1_LOC_761/Y 0.00fF
C32435 OR2X1_LOC_241/Y OR2X1_LOC_241/B 0.23fF
C32436 OR2X1_LOC_151/A AND2X1_LOC_92/Y 0.17fF
C32437 OR2X1_LOC_604/A OR2X1_LOC_684/a_8_216# 0.01fF
C32438 AND2X1_LOC_512/Y OR2X1_LOC_16/A 0.00fF
C32439 OR2X1_LOC_604/A AND2X1_LOC_705/a_8_24# 0.01fF
C32440 AND2X1_LOC_555/Y AND2X1_LOC_847/Y 0.02fF
C32441 OR2X1_LOC_426/A OR2X1_LOC_428/A 0.00fF
C32442 VDD AND2X1_LOC_568/B 0.59fF
C32443 OR2X1_LOC_56/A AND2X1_LOC_778/Y 0.04fF
C32444 OR2X1_LOC_600/A OR2X1_LOC_261/a_8_216# 0.03fF
C32445 AND2X1_LOC_335/Y AND2X1_LOC_337/a_8_24# 0.09fF
C32446 OR2X1_LOC_340/Y OR2X1_LOC_227/A 0.13fF
C32447 AND2X1_LOC_663/B OR2X1_LOC_437/A 0.09fF
C32448 AND2X1_LOC_729/B OR2X1_LOC_13/B 0.09fF
C32449 AND2X1_LOC_72/Y OR2X1_LOC_563/A 0.01fF
C32450 AND2X1_LOC_543/a_8_24# OR2X1_LOC_322/Y 0.04fF
C32451 OR2X1_LOC_809/B OR2X1_LOC_66/A 0.59fF
C32452 OR2X1_LOC_479/Y OR2X1_LOC_723/B 0.03fF
C32453 OR2X1_LOC_51/Y AND2X1_LOC_658/A 0.21fF
C32454 OR2X1_LOC_696/A OR2X1_LOC_753/A 0.10fF
C32455 OR2X1_LOC_130/A OR2X1_LOC_227/A 0.05fF
C32456 D_INPUT_0 OR2X1_LOC_80/A 0.89fF
C32457 OR2X1_LOC_4/a_8_216# OR2X1_LOC_68/B 0.47fF
C32458 AND2X1_LOC_91/B AND2X1_LOC_166/a_36_24# 0.01fF
C32459 OR2X1_LOC_541/a_8_216# OR2X1_LOC_121/A 0.01fF
C32460 OR2X1_LOC_600/A OR2X1_LOC_297/A 0.03fF
C32461 AND2X1_LOC_231/Y OR2X1_LOC_619/Y 0.03fF
C32462 AND2X1_LOC_352/B OR2X1_LOC_56/A 0.03fF
C32463 OR2X1_LOC_40/Y OR2X1_LOC_292/Y 0.01fF
C32464 OR2X1_LOC_770/a_8_216# OR2X1_LOC_68/B 0.01fF
C32465 VDD AND2X1_LOC_377/Y 0.01fF
C32466 OR2X1_LOC_109/a_36_216# OR2X1_LOC_373/Y 0.00fF
C32467 OR2X1_LOC_9/Y OR2X1_LOC_502/A 0.08fF
C32468 OR2X1_LOC_166/a_8_216# OR2X1_LOC_166/Y 0.01fF
C32469 AND2X1_LOC_658/A AND2X1_LOC_444/a_8_24# 0.04fF
C32470 AND2X1_LOC_727/a_8_24# AND2X1_LOC_621/Y 0.03fF
C32471 AND2X1_LOC_229/a_8_24# OR2X1_LOC_160/A 0.04fF
C32472 OR2X1_LOC_45/B OR2X1_LOC_306/Y 0.06fF
C32473 AND2X1_LOC_811/Y OR2X1_LOC_152/A 0.00fF
C32474 OR2X1_LOC_87/a_8_216# AND2X1_LOC_44/Y 0.01fF
C32475 OR2X1_LOC_770/B AND2X1_LOC_12/Y 0.00fF
C32476 INPUT_4 OR2X1_LOC_428/A 0.02fF
C32477 AND2X1_LOC_566/B AND2X1_LOC_364/A 0.01fF
C32478 OR2X1_LOC_345/Y OR2X1_LOC_791/B 0.01fF
C32479 AND2X1_LOC_51/Y AND2X1_LOC_36/Y 0.28fF
C32480 AND2X1_LOC_787/a_8_24# AND2X1_LOC_477/Y 0.01fF
C32481 OR2X1_LOC_49/A AND2X1_LOC_838/Y 1.02fF
C32482 OR2X1_LOC_832/a_8_216# OR2X1_LOC_502/A 0.03fF
C32483 AND2X1_LOC_500/Y AND2X1_LOC_508/A 0.05fF
C32484 AND2X1_LOC_363/Y OR2X1_LOC_494/a_8_216# 0.13fF
C32485 OR2X1_LOC_13/Y OR2X1_LOC_48/B 0.03fF
C32486 OR2X1_LOC_375/A OR2X1_LOC_375/Y 0.01fF
C32487 OR2X1_LOC_89/A OR2X1_LOC_767/Y 0.06fF
C32488 AND2X1_LOC_391/Y OR2X1_LOC_91/A 0.09fF
C32489 OR2X1_LOC_600/A AND2X1_LOC_866/B 0.03fF
C32490 OR2X1_LOC_269/a_8_216# OR2X1_LOC_549/A 0.01fF
C32491 OR2X1_LOC_589/A OR2X1_LOC_619/Y 0.10fF
C32492 OR2X1_LOC_314/Y OR2X1_LOC_12/Y 0.01fF
C32493 OR2X1_LOC_176/Y OR2X1_LOC_44/Y 0.03fF
C32494 AND2X1_LOC_736/Y VDD 0.11fF
C32495 AND2X1_LOC_59/Y OR2X1_LOC_736/Y 0.13fF
C32496 OR2X1_LOC_235/B INPUT_0 0.07fF
C32497 OR2X1_LOC_18/Y OR2X1_LOC_13/Y 0.03fF
C32498 OR2X1_LOC_375/A OR2X1_LOC_713/A 0.43fF
C32499 OR2X1_LOC_318/B OR2X1_LOC_374/Y 0.03fF
C32500 OR2X1_LOC_517/A OR2X1_LOC_56/A 0.28fF
C32501 OR2X1_LOC_36/Y AND2X1_LOC_456/a_36_24# 0.01fF
C32502 AND2X1_LOC_133/a_8_24# OR2X1_LOC_771/B 0.02fF
C32503 OR2X1_LOC_112/a_8_216# OR2X1_LOC_539/Y 0.03fF
C32504 OR2X1_LOC_656/B AND2X1_LOC_265/a_8_24# 0.01fF
C32505 AND2X1_LOC_86/Y OR2X1_LOC_6/B 0.20fF
C32506 OR2X1_LOC_207/B OR2X1_LOC_193/Y 0.21fF
C32507 AND2X1_LOC_554/Y AND2X1_LOC_362/B 0.07fF
C32508 OR2X1_LOC_335/A OR2X1_LOC_479/Y 0.02fF
C32509 AND2X1_LOC_12/Y OR2X1_LOC_596/A 1.29fF
C32510 AND2X1_LOC_719/Y AND2X1_LOC_287/a_8_24# 0.02fF
C32511 OR2X1_LOC_811/A AND2X1_LOC_18/Y 0.03fF
C32512 OR2X1_LOC_87/A AND2X1_LOC_603/a_8_24# 0.05fF
C32513 OR2X1_LOC_199/a_8_216# OR2X1_LOC_269/B 0.00fF
C32514 OR2X1_LOC_154/A OR2X1_LOC_833/Y 0.00fF
C32515 OR2X1_LOC_160/B OR2X1_LOC_523/Y 0.04fF
C32516 OR2X1_LOC_297/a_8_216# OR2X1_LOC_59/Y 0.02fF
C32517 AND2X1_LOC_707/Y AND2X1_LOC_454/A 0.20fF
C32518 OR2X1_LOC_179/Y OR2X1_LOC_59/Y 0.01fF
C32519 AND2X1_LOC_573/A OR2X1_LOC_131/a_8_216# 0.04fF
C32520 INPUT_3 OR2X1_LOC_6/B 0.27fF
C32521 AND2X1_LOC_398/a_8_24# OR2X1_LOC_600/A 0.05fF
C32522 OR2X1_LOC_759/A AND2X1_LOC_805/Y 0.01fF
C32523 AND2X1_LOC_51/Y OR2X1_LOC_333/a_8_216# 0.01fF
C32524 AND2X1_LOC_347/B AND2X1_LOC_848/a_8_24# 0.01fF
C32525 VDD OR2X1_LOC_738/B -0.00fF
C32526 AND2X1_LOC_648/B OR2X1_LOC_423/Y 0.02fF
C32527 AND2X1_LOC_212/Y OR2X1_LOC_44/Y 0.07fF
C32528 OR2X1_LOC_692/Y OR2X1_LOC_43/A 0.01fF
C32529 OR2X1_LOC_589/A OR2X1_LOC_88/A 0.01fF
C32530 OR2X1_LOC_176/a_8_216# AND2X1_LOC_566/Y 0.03fF
C32531 OR2X1_LOC_656/B VDD 0.09fF
C32532 OR2X1_LOC_756/B OR2X1_LOC_434/a_8_216# 0.01fF
C32533 OR2X1_LOC_18/Y AND2X1_LOC_244/a_36_24# 0.00fF
C32534 AND2X1_LOC_51/Y OR2X1_LOC_334/A 0.16fF
C32535 AND2X1_LOC_642/Y AND2X1_LOC_219/Y 0.03fF
C32536 OR2X1_LOC_66/Y OR2X1_LOC_560/A 0.02fF
C32537 OR2X1_LOC_377/A OR2X1_LOC_461/B 0.01fF
C32538 OR2X1_LOC_18/Y OR2X1_LOC_627/Y 0.19fF
C32539 AND2X1_LOC_377/Y OR2X1_LOC_689/A 0.03fF
C32540 OR2X1_LOC_158/A OR2X1_LOC_36/Y 0.73fF
C32541 OR2X1_LOC_107/Y AND2X1_LOC_113/a_8_24# 0.23fF
C32542 AND2X1_LOC_337/a_8_24# OR2X1_LOC_619/Y 0.05fF
C32543 INPUT_5 AND2X1_LOC_51/a_8_24# 0.01fF
C32544 OR2X1_LOC_458/a_8_216# OR2X1_LOC_464/A -0.00fF
C32545 AND2X1_LOC_280/a_36_24# OR2X1_LOC_78/A 0.00fF
C32546 OR2X1_LOC_160/A OR2X1_LOC_66/A 0.19fF
C32547 OR2X1_LOC_90/a_8_216# OR2X1_LOC_427/A 0.40fF
C32548 OR2X1_LOC_147/B OR2X1_LOC_147/A 0.06fF
C32549 AND2X1_LOC_824/B OR2X1_LOC_461/B 0.05fF
C32550 OR2X1_LOC_279/a_8_216# AND2X1_LOC_244/A 0.01fF
C32551 OR2X1_LOC_346/B OR2X1_LOC_346/A 0.05fF
C32552 OR2X1_LOC_680/A OR2X1_LOC_505/Y 0.03fF
C32553 AND2X1_LOC_721/a_8_24# AND2X1_LOC_456/B 0.01fF
C32554 AND2X1_LOC_658/B AND2X1_LOC_807/Y 0.02fF
C32555 AND2X1_LOC_468/B AND2X1_LOC_468/a_8_24# 0.01fF
C32556 AND2X1_LOC_652/a_8_24# AND2X1_LOC_436/Y 0.01fF
C32557 AND2X1_LOC_341/a_8_24# AND2X1_LOC_641/Y 0.20fF
C32558 AND2X1_LOC_148/a_8_24# OR2X1_LOC_427/A 0.04fF
C32559 AND2X1_LOC_59/Y OR2X1_LOC_641/Y 0.08fF
C32560 AND2X1_LOC_729/Y OR2X1_LOC_600/a_36_216# 0.00fF
C32561 AND2X1_LOC_862/Y AND2X1_LOC_866/B 0.86fF
C32562 OR2X1_LOC_709/A AND2X1_LOC_3/Y 0.35fF
C32563 AND2X1_LOC_578/A AND2X1_LOC_464/A 0.03fF
C32564 INPUT_3 AND2X1_LOC_73/a_8_24# 0.03fF
C32565 AND2X1_LOC_738/B AND2X1_LOC_624/A 0.07fF
C32566 AND2X1_LOC_3/Y AND2X1_LOC_295/a_8_24# 0.01fF
C32567 OR2X1_LOC_131/Y OR2X1_LOC_12/Y 0.31fF
C32568 OR2X1_LOC_857/B OR2X1_LOC_654/A 0.03fF
C32569 AND2X1_LOC_624/A OR2X1_LOC_56/A 0.07fF
C32570 AND2X1_LOC_99/A AND2X1_LOC_474/A 1.23fF
C32571 AND2X1_LOC_866/A AND2X1_LOC_792/B 0.02fF
C32572 OR2X1_LOC_680/A AND2X1_LOC_658/A 0.06fF
C32573 OR2X1_LOC_375/A OR2X1_LOC_803/A 0.00fF
C32574 OR2X1_LOC_696/A AND2X1_LOC_845/Y 0.07fF
C32575 AND2X1_LOC_356/a_36_24# OR2X1_LOC_56/A 0.01fF
C32576 OR2X1_LOC_425/a_8_216# OR2X1_LOC_2/Y 0.01fF
C32577 AND2X1_LOC_858/B AND2X1_LOC_573/A 0.10fF
C32578 VDD OR2X1_LOC_793/A 0.08fF
C32579 OR2X1_LOC_124/A OR2X1_LOC_375/A 0.37fF
C32580 OR2X1_LOC_91/A AND2X1_LOC_573/A 0.07fF
C32581 AND2X1_LOC_388/a_36_24# AND2X1_LOC_436/Y 0.00fF
C32582 OR2X1_LOC_600/A OR2X1_LOC_43/A 0.18fF
C32583 OR2X1_LOC_744/A AND2X1_LOC_114/a_8_24# 0.02fF
C32584 OR2X1_LOC_242/a_8_216# OR2X1_LOC_375/A 0.01fF
C32585 OR2X1_LOC_280/Y AND2X1_LOC_476/Y 0.21fF
C32586 D_INPUT_0 OR2X1_LOC_115/B 0.01fF
C32587 OR2X1_LOC_58/Y OR2X1_LOC_52/B 0.04fF
C32588 OR2X1_LOC_494/Y AND2X1_LOC_806/A 0.10fF
C32589 AND2X1_LOC_734/Y AND2X1_LOC_550/A 3.04fF
C32590 OR2X1_LOC_506/Y AND2X1_LOC_51/Y 0.01fF
C32591 AND2X1_LOC_566/B OR2X1_LOC_3/Y 0.03fF
C32592 OR2X1_LOC_100/Y AND2X1_LOC_517/a_8_24# 0.08fF
C32593 AND2X1_LOC_725/a_8_24# OR2X1_LOC_7/A 0.05fF
C32594 OR2X1_LOC_440/A OR2X1_LOC_168/Y 0.00fF
C32595 OR2X1_LOC_323/A OR2X1_LOC_111/Y 0.01fF
C32596 AND2X1_LOC_12/Y OR2X1_LOC_808/A 0.03fF
C32597 AND2X1_LOC_199/A AND2X1_LOC_729/B 0.01fF
C32598 OR2X1_LOC_223/A OR2X1_LOC_776/A 0.00fF
C32599 OR2X1_LOC_166/a_8_216# OR2X1_LOC_43/A 0.01fF
C32600 OR2X1_LOC_697/Y OR2X1_LOC_39/A 0.03fF
C32601 OR2X1_LOC_438/Y AND2X1_LOC_621/Y 0.03fF
C32602 AND2X1_LOC_302/a_36_24# OR2X1_LOC_59/Y 0.01fF
C32603 AND2X1_LOC_654/B OR2X1_LOC_619/Y 0.96fF
C32604 OR2X1_LOC_311/Y AND2X1_LOC_802/Y 0.02fF
C32605 OR2X1_LOC_43/A AND2X1_LOC_296/a_8_24# 0.01fF
C32606 AND2X1_LOC_59/Y OR2X1_LOC_808/B 2.25fF
C32607 OR2X1_LOC_702/A AND2X1_LOC_110/Y 0.05fF
C32608 AND2X1_LOC_94/Y OR2X1_LOC_82/a_36_216# 0.02fF
C32609 OR2X1_LOC_54/Y OR2X1_LOC_16/A 0.02fF
C32610 AND2X1_LOC_86/B OR2X1_LOC_66/A 0.06fF
C32611 OR2X1_LOC_643/A OR2X1_LOC_632/Y 0.00fF
C32612 OR2X1_LOC_807/B OR2X1_LOC_811/A 0.05fF
C32613 OR2X1_LOC_604/A OR2X1_LOC_430/a_8_216# 0.02fF
C32614 OR2X1_LOC_8/Y OR2X1_LOC_485/A 1.19fF
C32615 AND2X1_LOC_70/Y AND2X1_LOC_3/Y 2.36fF
C32616 AND2X1_LOC_597/a_8_24# AND2X1_LOC_41/A 0.01fF
C32617 OR2X1_LOC_3/Y OR2X1_LOC_695/Y 0.01fF
C32618 OR2X1_LOC_663/A OR2X1_LOC_204/Y 0.03fF
C32619 AND2X1_LOC_314/a_8_24# OR2X1_LOC_447/A 0.20fF
C32620 OR2X1_LOC_547/B OR2X1_LOC_220/B 0.31fF
C32621 OR2X1_LOC_624/B OR2X1_LOC_66/A 0.03fF
C32622 OR2X1_LOC_720/B OR2X1_LOC_161/B 0.14fF
C32623 OR2X1_LOC_864/A AND2X1_LOC_41/A 0.13fF
C32624 OR2X1_LOC_252/a_36_216# AND2X1_LOC_805/Y 0.00fF
C32625 AND2X1_LOC_36/Y OR2X1_LOC_551/B 0.07fF
C32626 OR2X1_LOC_217/Y OR2X1_LOC_502/A 0.06fF
C32627 OR2X1_LOC_401/Y OR2X1_LOC_78/a_8_216# 0.01fF
C32628 OR2X1_LOC_600/A OR2X1_LOC_60/a_8_216# 0.05fF
C32629 OR2X1_LOC_666/A OR2X1_LOC_279/a_36_216# 0.00fF
C32630 AND2X1_LOC_385/a_36_24# AND2X1_LOC_41/A 0.01fF
C32631 AND2X1_LOC_850/Y AND2X1_LOC_624/A 0.42fF
C32632 AND2X1_LOC_367/A AND2X1_LOC_294/a_8_24# 0.02fF
C32633 AND2X1_LOC_191/B OR2X1_LOC_754/A 0.03fF
C32634 AND2X1_LOC_42/B OR2X1_LOC_78/A 0.10fF
C32635 AND2X1_LOC_753/B OR2X1_LOC_87/A 0.20fF
C32636 OR2X1_LOC_619/Y AND2X1_LOC_622/a_8_24# 0.10fF
C32637 AND2X1_LOC_365/A OR2X1_LOC_619/Y 0.09fF
C32638 OR2X1_LOC_290/a_8_216# OR2X1_LOC_585/A 0.03fF
C32639 OR2X1_LOC_395/Y OR2X1_LOC_598/A 0.25fF
C32640 AND2X1_LOC_270/a_8_24# AND2X1_LOC_786/Y 0.05fF
C32641 AND2X1_LOC_512/Y AND2X1_LOC_336/a_8_24# 0.02fF
C32642 AND2X1_LOC_511/a_36_24# AND2X1_LOC_48/A 0.01fF
C32643 OR2X1_LOC_319/B AND2X1_LOC_329/a_8_24# 0.23fF
C32644 OR2X1_LOC_68/B OR2X1_LOC_723/B 0.12fF
C32645 AND2X1_LOC_56/B AND2X1_LOC_482/a_8_24# 0.01fF
C32646 OR2X1_LOC_600/A AND2X1_LOC_664/a_8_24# 0.01fF
C32647 AND2X1_LOC_721/a_36_24# OR2X1_LOC_26/Y 0.00fF
C32648 OR2X1_LOC_854/a_8_216# OR2X1_LOC_155/A 0.02fF
C32649 OR2X1_LOC_405/A OR2X1_LOC_87/A 0.17fF
C32650 OR2X1_LOC_47/Y OR2X1_LOC_816/A 0.04fF
C32651 OR2X1_LOC_458/B AND2X1_LOC_42/B 0.04fF
C32652 AND2X1_LOC_31/Y INPUT_6 0.04fF
C32653 OR2X1_LOC_62/A OR2X1_LOC_633/A 0.09fF
C32654 AND2X1_LOC_87/a_36_24# OR2X1_LOC_619/Y 0.01fF
C32655 OR2X1_LOC_405/Y OR2X1_LOC_222/A 0.08fF
C32656 AND2X1_LOC_779/a_36_24# OR2X1_LOC_599/A 0.00fF
C32657 OR2X1_LOC_808/A OR2X1_LOC_804/B 0.93fF
C32658 OR2X1_LOC_76/Y OR2X1_LOC_833/B 0.00fF
C32659 AND2X1_LOC_391/a_8_24# OR2X1_LOC_3/Y 0.01fF
C32660 OR2X1_LOC_6/B OR2X1_LOC_244/A 0.07fF
C32661 OR2X1_LOC_43/A OR2X1_LOC_619/Y 0.10fF
C32662 AND2X1_LOC_65/a_8_24# OR2X1_LOC_215/A 0.08fF
C32663 OR2X1_LOC_201/A OR2X1_LOC_206/a_8_216# 0.01fF
C32664 AND2X1_LOC_356/a_8_24# OR2X1_LOC_43/A 0.01fF
C32665 OR2X1_LOC_190/A OR2X1_LOC_471/Y 0.08fF
C32666 OR2X1_LOC_235/B OR2X1_LOC_64/Y 0.66fF
C32667 AND2X1_LOC_663/B OR2X1_LOC_755/Y 0.01fF
C32668 OR2X1_LOC_117/Y OR2X1_LOC_118/Y 0.03fF
C32669 OR2X1_LOC_574/A OR2X1_LOC_620/Y 0.07fF
C32670 OR2X1_LOC_256/A AND2X1_LOC_243/Y 0.07fF
C32671 OR2X1_LOC_112/B OR2X1_LOC_435/A 0.43fF
C32672 AND2X1_LOC_563/A OR2X1_LOC_71/Y 0.00fF
C32673 OR2X1_LOC_95/Y AND2X1_LOC_499/a_8_24# 0.01fF
C32674 OR2X1_LOC_124/a_8_216# D_INPUT_0 0.02fF
C32675 OR2X1_LOC_346/B OR2X1_LOC_161/A 0.12fF
C32676 AND2X1_LOC_95/Y OR2X1_LOC_564/A 0.09fF
C32677 OR2X1_LOC_681/a_8_216# OR2X1_LOC_31/Y 0.18fF
C32678 AND2X1_LOC_351/a_8_24# OR2X1_LOC_289/Y 0.01fF
C32679 OR2X1_LOC_485/A AND2X1_LOC_76/Y 0.00fF
C32680 OR2X1_LOC_74/A AND2X1_LOC_804/Y 0.12fF
C32681 OR2X1_LOC_160/B AND2X1_LOC_47/Y 0.59fF
C32682 OR2X1_LOC_216/A OR2X1_LOC_473/Y 0.01fF
C32683 OR2X1_LOC_9/Y OR2X1_LOC_618/Y 0.01fF
C32684 AND2X1_LOC_148/Y OR2X1_LOC_427/A 0.09fF
C32685 AND2X1_LOC_50/Y AND2X1_LOC_1/Y 0.02fF
C32686 OR2X1_LOC_130/A OR2X1_LOC_269/B 0.02fF
C32687 OR2X1_LOC_635/A AND2X1_LOC_51/Y 0.00fF
C32688 AND2X1_LOC_380/a_8_24# AND2X1_LOC_3/Y 0.01fF
C32689 INPUT_1 AND2X1_LOC_92/Y 0.01fF
C32690 OR2X1_LOC_532/B OR2X1_LOC_244/Y 0.03fF
C32691 OR2X1_LOC_604/A OR2X1_LOC_428/Y 0.02fF
C32692 OR2X1_LOC_113/A OR2X1_LOC_632/Y 0.01fF
C32693 AND2X1_LOC_729/Y OR2X1_LOC_420/a_8_216# 0.05fF
C32694 OR2X1_LOC_624/Y OR2X1_LOC_814/A 0.02fF
C32695 OR2X1_LOC_405/A OR2X1_LOC_216/a_8_216# 0.04fF
C32696 OR2X1_LOC_122/a_8_216# AND2X1_LOC_845/Y 0.02fF
C32697 OR2X1_LOC_791/B AND2X1_LOC_3/Y 0.06fF
C32698 AND2X1_LOC_658/B OR2X1_LOC_95/Y 0.06fF
C32699 OR2X1_LOC_127/a_8_216# OR2X1_LOC_3/Y 0.09fF
C32700 OR2X1_LOC_502/A AND2X1_LOC_680/a_8_24# 0.03fF
C32701 OR2X1_LOC_287/B AND2X1_LOC_82/a_8_24# 0.01fF
C32702 AND2X1_LOC_376/a_8_24# OR2X1_LOC_463/B 0.23fF
C32703 OR2X1_LOC_566/A OR2X1_LOC_353/a_8_216# 0.00fF
C32704 OR2X1_LOC_814/A OR2X1_LOC_391/A 0.04fF
C32705 OR2X1_LOC_231/A OR2X1_LOC_215/A 0.31fF
C32706 OR2X1_LOC_678/a_8_216# AND2X1_LOC_53/Y 0.04fF
C32707 AND2X1_LOC_12/Y OR2X1_LOC_33/B 0.00fF
C32708 AND2X1_LOC_120/a_8_24# OR2X1_LOC_18/Y 0.02fF
C32709 AND2X1_LOC_91/B OR2X1_LOC_724/A 0.07fF
C32710 OR2X1_LOC_154/A OR2X1_LOC_574/A 0.11fF
C32711 OR2X1_LOC_744/A AND2X1_LOC_656/Y 0.03fF
C32712 AND2X1_LOC_359/a_8_24# OR2X1_LOC_753/A 0.01fF
C32713 OR2X1_LOC_81/Y OR2X1_LOC_52/B 0.04fF
C32714 AND2X1_LOC_716/Y OR2X1_LOC_46/A 0.07fF
C32715 OR2X1_LOC_427/A OR2X1_LOC_683/Y 0.01fF
C32716 OR2X1_LOC_191/B OR2X1_LOC_551/a_8_216# 0.14fF
C32717 OR2X1_LOC_8/Y OR2X1_LOC_10/a_8_216# 0.06fF
C32718 OR2X1_LOC_409/B OR2X1_LOC_25/Y 0.03fF
C32719 OR2X1_LOC_193/Y AND2X1_LOC_3/Y 0.03fF
C32720 AND2X1_LOC_702/Y OR2X1_LOC_7/A 0.03fF
C32721 AND2X1_LOC_576/Y OR2X1_LOC_89/A 0.24fF
C32722 OR2X1_LOC_290/Y INPUT_1 0.26fF
C32723 AND2X1_LOC_243/Y OR2X1_LOC_67/Y 0.67fF
C32724 OR2X1_LOC_46/A OR2X1_LOC_393/a_8_216# 0.01fF
C32725 OR2X1_LOC_116/a_8_216# AND2X1_LOC_3/Y -0.00fF
C32726 AND2X1_LOC_500/a_8_24# OR2X1_LOC_239/Y 0.01fF
C32727 OR2X1_LOC_792/Y OR2X1_LOC_285/Y 0.03fF
C32728 AND2X1_LOC_654/Y OR2X1_LOC_46/A 0.07fF
C32729 OR2X1_LOC_377/A OR2X1_LOC_99/B 0.01fF
C32730 AND2X1_LOC_17/Y AND2X1_LOC_3/Y 0.05fF
C32731 AND2X1_LOC_702/Y OR2X1_LOC_320/Y 0.01fF
C32732 OR2X1_LOC_130/A OR2X1_LOC_215/A 0.03fF
C32733 OR2X1_LOC_485/A OR2X1_LOC_52/B 0.08fF
C32734 OR2X1_LOC_472/a_36_216# AND2X1_LOC_824/B -0.00fF
C32735 OR2X1_LOC_12/Y AND2X1_LOC_657/A 0.04fF
C32736 OR2X1_LOC_230/a_8_216# OR2X1_LOC_6/A 0.02fF
C32737 OR2X1_LOC_151/A OR2X1_LOC_736/a_8_216# 0.01fF
C32738 OR2X1_LOC_147/B OR2X1_LOC_532/B 0.04fF
C32739 OR2X1_LOC_535/A OR2X1_LOC_568/A 0.02fF
C32740 AND2X1_LOC_319/A OR2X1_LOC_64/Y 0.10fF
C32741 OR2X1_LOC_160/B OR2X1_LOC_598/A 0.14fF
C32742 OR2X1_LOC_22/Y OR2X1_LOC_595/a_8_216# 0.02fF
C32743 OR2X1_LOC_673/B OR2X1_LOC_80/A 0.02fF
C32744 AND2X1_LOC_113/a_8_24# AND2X1_LOC_866/A 0.06fF
C32745 OR2X1_LOC_317/A OR2X1_LOC_532/B 0.01fF
C32746 AND2X1_LOC_12/Y OR2X1_LOC_287/a_8_216# 0.01fF
C32747 AND2X1_LOC_663/B OR2X1_LOC_753/A 0.10fF
C32748 OR2X1_LOC_731/B OR2X1_LOC_731/A 0.16fF
C32749 OR2X1_LOC_602/B AND2X1_LOC_43/B 0.05fF
C32750 OR2X1_LOC_755/A OR2X1_LOC_665/Y 0.01fF
C32751 OR2X1_LOC_327/a_36_216# OR2X1_LOC_218/Y 0.00fF
C32752 INPUT_3 AND2X1_LOC_47/Y 0.09fF
C32753 AND2X1_LOC_211/B AND2X1_LOC_326/A 0.02fF
C32754 OR2X1_LOC_3/Y OR2X1_LOC_817/Y 0.02fF
C32755 OR2X1_LOC_91/Y INPUT_1 0.18fF
C32756 OR2X1_LOC_404/Y AND2X1_LOC_3/Y 0.03fF
C32757 OR2X1_LOC_436/Y OR2X1_LOC_506/A 0.09fF
C32758 AND2X1_LOC_47/Y AND2X1_LOC_297/a_36_24# 0.00fF
C32759 OR2X1_LOC_473/A OR2X1_LOC_737/A 0.01fF
C32760 OR2X1_LOC_532/B AND2X1_LOC_669/a_8_24# 0.01fF
C32761 OR2X1_LOC_550/B OR2X1_LOC_550/A 0.05fF
C32762 AND2X1_LOC_502/a_8_24# AND2X1_LOC_227/Y 0.01fF
C32763 AND2X1_LOC_641/Y AND2X1_LOC_650/a_36_24# 0.01fF
C32764 D_INPUT_0 OR2X1_LOC_6/A 0.36fF
C32765 AND2X1_LOC_537/Y OR2X1_LOC_585/A 0.01fF
C32766 AND2X1_LOC_558/a_8_24# AND2X1_LOC_563/Y 0.01fF
C32767 AND2X1_LOC_59/Y OR2X1_LOC_218/Y 0.00fF
C32768 OR2X1_LOC_648/A AND2X1_LOC_31/Y 0.16fF
C32769 OR2X1_LOC_405/A AND2X1_LOC_109/a_36_24# 0.00fF
C32770 OR2X1_LOC_121/a_8_216# AND2X1_LOC_36/Y 0.05fF
C32771 OR2X1_LOC_160/A OR2X1_LOC_84/A 0.27fF
C32772 OR2X1_LOC_612/a_36_216# OR2X1_LOC_71/A 0.00fF
C32773 INPUT_1 OR2X1_LOC_371/a_8_216# 0.03fF
C32774 OR2X1_LOC_549/B OR2X1_LOC_562/A 0.01fF
C32775 OR2X1_LOC_628/a_8_216# AND2X1_LOC_483/Y 0.01fF
C32776 OR2X1_LOC_47/Y AND2X1_LOC_807/Y 0.02fF
C32777 OR2X1_LOC_863/B OR2X1_LOC_19/B 0.03fF
C32778 OR2X1_LOC_72/a_8_216# AND2X1_LOC_361/A 0.47fF
C32779 AND2X1_LOC_845/Y OR2X1_LOC_89/a_8_216# 0.04fF
C32780 AND2X1_LOC_392/A OR2X1_LOC_437/A 0.07fF
C32781 AND2X1_LOC_700/a_8_24# OR2X1_LOC_732/A 0.23fF
C32782 OR2X1_LOC_681/Y AND2X1_LOC_687/A 0.01fF
C32783 OR2X1_LOC_71/Y AND2X1_LOC_717/B 0.00fF
C32784 OR2X1_LOC_449/A OR2X1_LOC_783/A 0.26fF
C32785 OR2X1_LOC_495/a_36_216# AND2X1_LOC_851/B 0.01fF
C32786 AND2X1_LOC_72/B AND2X1_LOC_297/a_8_24# 0.10fF
C32787 AND2X1_LOC_387/B OR2X1_LOC_532/B 0.11fF
C32788 AND2X1_LOC_18/Y OR2X1_LOC_777/B 0.03fF
C32789 AND2X1_LOC_86/Y OR2X1_LOC_598/A 0.12fF
C32790 OR2X1_LOC_47/Y OR2X1_LOC_824/Y 0.07fF
C32791 OR2X1_LOC_87/A OR2X1_LOC_779/Y 0.02fF
C32792 OR2X1_LOC_696/A OR2X1_LOC_323/Y 0.29fF
C32793 AND2X1_LOC_12/Y OR2X1_LOC_374/Y 0.03fF
C32794 OR2X1_LOC_684/Y AND2X1_LOC_686/a_8_24# 0.02fF
C32795 AND2X1_LOC_433/a_8_24# OR2X1_LOC_390/B 0.03fF
C32796 AND2X1_LOC_40/Y OR2X1_LOC_80/A 0.03fF
C32797 OR2X1_LOC_351/B OR2X1_LOC_333/A 0.01fF
C32798 AND2X1_LOC_366/A OR2X1_LOC_437/A 0.06fF
C32799 OR2X1_LOC_291/Y INPUT_1 0.00fF
C32800 AND2X1_LOC_92/Y OR2X1_LOC_716/a_8_216# 0.04fF
C32801 OR2X1_LOC_554/a_8_216# OR2X1_LOC_161/B 0.03fF
C32802 AND2X1_LOC_95/Y OR2X1_LOC_228/Y 0.10fF
C32803 OR2X1_LOC_18/Y AND2X1_LOC_563/Y 0.03fF
C32804 OR2X1_LOC_812/B OR2X1_LOC_68/B 0.53fF
C32805 OR2X1_LOC_287/B D_INPUT_1 0.06fF
C32806 AND2X1_LOC_469/B OR2X1_LOC_142/Y 0.03fF
C32807 OR2X1_LOC_624/B OR2X1_LOC_84/A 0.01fF
C32808 AND2X1_LOC_513/a_8_24# OR2X1_LOC_13/B 0.01fF
C32809 OR2X1_LOC_121/Y OR2X1_LOC_392/B 0.10fF
C32810 OR2X1_LOC_399/A OR2X1_LOC_80/A 0.02fF
C32811 OR2X1_LOC_428/A OR2X1_LOC_759/a_8_216# 0.06fF
C32812 AND2X1_LOC_208/Y AND2X1_LOC_214/a_36_24# 0.01fF
C32813 OR2X1_LOC_269/B OR2X1_LOC_365/B 0.03fF
C32814 AND2X1_LOC_358/a_36_24# OR2X1_LOC_417/A 0.00fF
C32815 AND2X1_LOC_131/a_8_24# OR2X1_LOC_115/B 0.01fF
C32816 OR2X1_LOC_140/A OR2X1_LOC_140/B 0.00fF
C32817 OR2X1_LOC_3/B OR2X1_LOC_17/Y 0.02fF
C32818 OR2X1_LOC_51/B OR2X1_LOC_44/a_8_216# 0.04fF
C32819 AND2X1_LOC_733/Y OR2X1_LOC_142/Y 0.07fF
C32820 OR2X1_LOC_85/A OR2X1_LOC_72/Y 0.03fF
C32821 OR2X1_LOC_563/A OR2X1_LOC_719/B 0.02fF
C32822 OR2X1_LOC_675/a_8_216# OR2X1_LOC_241/B 0.01fF
C32823 OR2X1_LOC_831/B AND2X1_LOC_18/Y 0.03fF
C32824 OR2X1_LOC_129/a_8_216# AND2X1_LOC_202/Y 0.00fF
C32825 AND2X1_LOC_636/a_8_24# OR2X1_LOC_584/Y 0.00fF
C32826 OR2X1_LOC_502/A OR2X1_LOC_771/B 0.03fF
C32827 AND2X1_LOC_420/a_36_24# AND2X1_LOC_51/Y 0.00fF
C32828 OR2X1_LOC_375/A OR2X1_LOC_546/A 0.04fF
C32829 AND2X1_LOC_787/A AND2X1_LOC_477/Y 0.01fF
C32830 OR2X1_LOC_188/a_8_216# AND2X1_LOC_18/Y -0.00fF
C32831 AND2X1_LOC_845/Y AND2X1_LOC_849/a_8_24# 0.07fF
C32832 OR2X1_LOC_848/A OR2X1_LOC_80/A 0.61fF
C32833 OR2X1_LOC_595/A AND2X1_LOC_249/a_36_24# 0.00fF
C32834 OR2X1_LOC_244/A AND2X1_LOC_47/Y 0.07fF
C32835 AND2X1_LOC_51/a_36_24# INPUT_6 0.00fF
C32836 OR2X1_LOC_64/Y AND2X1_LOC_721/A 0.03fF
C32837 AND2X1_LOC_727/A OR2X1_LOC_47/Y 0.03fF
C32838 D_INPUT_3 INPUT_1 0.35fF
C32839 D_INPUT_2 D_INPUT_0 0.38fF
C32840 OR2X1_LOC_93/Y OR2X1_LOC_428/A 0.01fF
C32841 OR2X1_LOC_542/B OR2X1_LOC_563/A 0.07fF
C32842 AND2X1_LOC_164/a_36_24# OR2X1_LOC_390/B 0.00fF
C32843 OR2X1_LOC_744/A AND2X1_LOC_772/Y 0.01fF
C32844 OR2X1_LOC_765/Y OR2X1_LOC_16/A 0.04fF
C32845 AND2X1_LOC_570/Y AND2X1_LOC_242/B 0.02fF
C32846 OR2X1_LOC_266/A OR2X1_LOC_66/A 0.01fF
C32847 AND2X1_LOC_91/B OR2X1_LOC_632/Y 0.10fF
C32848 AND2X1_LOC_447/Y OR2X1_LOC_428/A 0.00fF
C32849 AND2X1_LOC_851/B OR2X1_LOC_238/a_36_216# 0.01fF
C32850 AND2X1_LOC_660/a_8_24# AND2X1_LOC_660/A 0.02fF
C32851 VDD OR2X1_LOC_12/Y 0.89fF
C32852 AND2X1_LOC_18/Y OR2X1_LOC_344/A 0.04fF
C32853 OR2X1_LOC_634/A OR2X1_LOC_338/A 0.02fF
C32854 VDD OR2X1_LOC_766/Y 0.04fF
C32855 AND2X1_LOC_182/A OR2X1_LOC_309/Y 0.16fF
C32856 AND2X1_LOC_41/A OR2X1_LOC_121/A 0.05fF
C32857 OR2X1_LOC_47/Y OR2X1_LOC_95/Y 0.86fF
C32858 OR2X1_LOC_604/A OR2X1_LOC_158/A 0.95fF
C32859 OR2X1_LOC_857/B VDD 0.05fF
C32860 OR2X1_LOC_400/A OR2X1_LOC_771/B 0.02fF
C32861 OR2X1_LOC_738/A OR2X1_LOC_726/a_8_216# 0.05fF
C32862 OR2X1_LOC_56/A AND2X1_LOC_774/A 1.78fF
C32863 OR2X1_LOC_604/A AND2X1_LOC_704/a_36_24# 0.00fF
C32864 OR2X1_LOC_45/B AND2X1_LOC_549/a_8_24# 0.03fF
C32865 AND2X1_LOC_264/a_8_24# OR2X1_LOC_13/B 0.06fF
C32866 OR2X1_LOC_64/Y OR2X1_LOC_331/Y 0.19fF
C32867 AND2X1_LOC_59/Y OR2X1_LOC_703/Y 0.01fF
C32868 AND2X1_LOC_607/a_8_24# OR2X1_LOC_66/A 0.14fF
C32869 OR2X1_LOC_213/A OR2X1_LOC_209/A 0.03fF
C32870 OR2X1_LOC_45/B AND2X1_LOC_506/a_8_24# 0.03fF
C32871 AND2X1_LOC_12/Y OR2X1_LOC_333/A 0.01fF
C32872 OR2X1_LOC_831/a_8_216# AND2X1_LOC_36/Y 0.01fF
C32873 OR2X1_LOC_106/A OR2X1_LOC_13/B 0.03fF
C32874 OR2X1_LOC_607/a_36_216# OR2X1_LOC_67/Y 0.01fF
C32875 OR2X1_LOC_715/B OR2X1_LOC_676/Y 0.00fF
C32876 AND2X1_LOC_217/Y AND2X1_LOC_218/a_8_24# 0.03fF
C32877 OR2X1_LOC_405/A OR2X1_LOC_390/B 0.14fF
C32878 OR2X1_LOC_124/A OR2X1_LOC_549/A 0.09fF
C32879 OR2X1_LOC_244/A OR2X1_LOC_598/A 0.02fF
C32880 OR2X1_LOC_709/A INPUT_0 0.00fF
C32881 AND2X1_LOC_300/a_8_24# AND2X1_LOC_92/Y 0.00fF
C32882 AND2X1_LOC_729/Y OR2X1_LOC_696/A 0.07fF
C32883 AND2X1_LOC_392/A AND2X1_LOC_715/A 0.03fF
C32884 OR2X1_LOC_421/A OR2X1_LOC_426/B 0.02fF
C32885 AND2X1_LOC_566/B OR2X1_LOC_329/B 0.06fF
C32886 INPUT_0 OR2X1_LOC_57/a_8_216# 0.05fF
C32887 AND2X1_LOC_215/Y AND2X1_LOC_334/Y 0.01fF
C32888 OR2X1_LOC_3/B OR2X1_LOC_588/A 0.01fF
C32889 OR2X1_LOC_532/B OR2X1_LOC_854/A 0.00fF
C32890 AND2X1_LOC_59/Y OR2X1_LOC_120/a_8_216# 0.01fF
C32891 OR2X1_LOC_49/A AND2X1_LOC_852/B 0.02fF
C32892 AND2X1_LOC_803/B AND2X1_LOC_738/B 0.06fF
C32893 OR2X1_LOC_333/B OR2X1_LOC_539/B 0.02fF
C32894 OR2X1_LOC_696/A AND2X1_LOC_784/A 0.07fF
C32895 OR2X1_LOC_89/A AND2X1_LOC_793/a_8_24# 0.01fF
C32896 AND2X1_LOC_567/a_8_24# OR2X1_LOC_744/A 0.02fF
C32897 OR2X1_LOC_625/Y OR2X1_LOC_816/A 1.03fF
C32898 AND2X1_LOC_12/Y OR2X1_LOC_392/B 0.01fF
C32899 AND2X1_LOC_91/B AND2X1_LOC_251/a_8_24# 0.02fF
C32900 AND2X1_LOC_729/Y AND2X1_LOC_715/Y 0.83fF
C32901 OR2X1_LOC_840/A OR2X1_LOC_831/A 0.01fF
C32902 OR2X1_LOC_778/Y OR2X1_LOC_168/Y 0.19fF
C32903 AND2X1_LOC_51/Y OR2X1_LOC_571/Y 0.23fF
C32904 OR2X1_LOC_741/Y OR2X1_LOC_742/a_8_216# 0.07fF
C32905 OR2X1_LOC_109/Y OR2X1_LOC_428/A 0.03fF
C32906 OR2X1_LOC_154/A OR2X1_LOC_390/a_8_216# 0.02fF
C32907 OR2X1_LOC_123/a_36_216# OR2X1_LOC_124/A 0.00fF
C32908 AND2X1_LOC_91/B OR2X1_LOC_561/a_8_216# 0.01fF
C32909 OR2X1_LOC_757/A AND2X1_LOC_658/A 0.03fF
C32910 OR2X1_LOC_28/a_8_216# D_INPUT_1 0.01fF
C32911 OR2X1_LOC_56/A AND2X1_LOC_434/a_8_24# 0.04fF
C32912 AND2X1_LOC_658/Y AND2X1_LOC_663/A 0.01fF
C32913 AND2X1_LOC_448/Y OR2X1_LOC_428/A 0.07fF
C32914 OR2X1_LOC_585/A OR2X1_LOC_171/a_8_216# 0.02fF
C32915 AND2X1_LOC_70/Y INPUT_0 0.07fF
C32916 OR2X1_LOC_188/Y OR2X1_LOC_457/B 0.22fF
C32917 AND2X1_LOC_562/a_8_24# OR2X1_LOC_36/Y 0.03fF
C32918 OR2X1_LOC_442/Y AND2X1_LOC_469/B 0.01fF
C32919 AND2X1_LOC_534/a_36_24# OR2X1_LOC_620/Y 0.00fF
C32920 OR2X1_LOC_624/Y OR2X1_LOC_244/Y 0.02fF
C32921 OR2X1_LOC_46/A OR2X1_LOC_13/B 0.03fF
C32922 VDD OR2X1_LOC_837/Y 0.22fF
C32923 OR2X1_LOC_49/A AND2X1_LOC_59/Y 0.03fF
C32924 OR2X1_LOC_358/a_8_216# OR2X1_LOC_97/A 0.01fF
C32925 OR2X1_LOC_364/A AND2X1_LOC_91/a_8_24# 0.01fF
C32926 OR2X1_LOC_45/B OR2X1_LOC_265/Y 0.11fF
C32927 AND2X1_LOC_56/B OR2X1_LOC_563/A 0.01fF
C32928 OR2X1_LOC_505/a_36_216# AND2X1_LOC_807/Y 0.15fF
C32929 OR2X1_LOC_709/A OR2X1_LOC_732/B 0.05fF
C32930 AND2X1_LOC_585/a_8_24# OR2X1_LOC_160/A -0.00fF
C32931 AND2X1_LOC_721/Y OR2X1_LOC_36/Y 0.02fF
C32932 OR2X1_LOC_709/A OR2X1_LOC_789/B 0.01fF
C32933 OR2X1_LOC_604/A OR2X1_LOC_594/Y 0.14fF
C32934 OR2X1_LOC_158/A AND2X1_LOC_850/a_8_24# 0.01fF
C32935 AND2X1_LOC_564/B AND2X1_LOC_458/a_8_24# 0.06fF
C32936 AND2X1_LOC_48/A OR2X1_LOC_771/B 0.06fF
C32937 AND2X1_LOC_18/Y OR2X1_LOC_575/A 0.03fF
C32938 AND2X1_LOC_574/a_8_24# AND2X1_LOC_675/Y 0.18fF
C32939 VDD OR2X1_LOC_785/B 0.33fF
C32940 AND2X1_LOC_456/Y AND2X1_LOC_465/A 0.09fF
C32941 OR2X1_LOC_12/Y AND2X1_LOC_447/a_36_24# -0.02fF
C32942 AND2X1_LOC_31/a_8_24# INPUT_6 0.01fF
C32943 OR2X1_LOC_663/A OR2X1_LOC_78/A 0.03fF
C32944 AND2X1_LOC_70/Y OR2X1_LOC_775/a_8_216# 0.01fF
C32945 AND2X1_LOC_574/Y AND2X1_LOC_191/Y 0.04fF
C32946 AND2X1_LOC_734/Y AND2X1_LOC_663/A 1.17fF
C32947 OR2X1_LOC_214/B OR2X1_LOC_750/Y 0.10fF
C32948 OR2X1_LOC_814/A OR2X1_LOC_174/Y 0.00fF
C32949 OR2X1_LOC_540/a_8_216# OR2X1_LOC_190/Y 0.40fF
C32950 OR2X1_LOC_271/a_36_216# AND2X1_LOC_786/Y 0.01fF
C32951 AND2X1_LOC_598/a_8_24# OR2X1_LOC_16/A 0.01fF
C32952 OR2X1_LOC_141/B OR2X1_LOC_267/Y 0.67fF
C32953 OR2X1_LOC_671/Y AND2X1_LOC_838/Y 0.02fF
C32954 OR2X1_LOC_425/a_8_216# OR2X1_LOC_25/Y 0.04fF
C32955 AND2X1_LOC_110/Y OR2X1_LOC_623/a_8_216# 0.01fF
C32956 AND2X1_LOC_476/Y OR2X1_LOC_39/A 0.10fF
C32957 OR2X1_LOC_667/Y OR2X1_LOC_494/Y 0.01fF
C32958 AND2X1_LOC_574/Y AND2X1_LOC_711/Y 0.03fF
C32959 OR2X1_LOC_599/A AND2X1_LOC_724/A 0.11fF
C32960 AND2X1_LOC_227/Y OR2X1_LOC_13/B 0.03fF
C32961 AND2X1_LOC_503/a_8_24# OR2X1_LOC_78/A 0.02fF
C32962 OR2X1_LOC_26/Y OR2X1_LOC_16/A 1.25fF
C32963 AND2X1_LOC_544/Y AND2X1_LOC_728/a_36_24# 0.01fF
C32964 VDD OR2X1_LOC_393/Y 0.07fF
C32965 OR2X1_LOC_447/A OR2X1_LOC_66/A 0.02fF
C32966 OR2X1_LOC_158/A OR2X1_LOC_80/Y 0.01fF
C32967 OR2X1_LOC_188/Y OR2X1_LOC_675/a_8_216# 0.00fF
C32968 OR2X1_LOC_391/B D_GATE_662 0.02fF
C32969 AND2X1_LOC_193/a_8_24# AND2X1_LOC_193/Y 0.00fF
C32970 OR2X1_LOC_405/A OR2X1_LOC_493/a_8_216# 0.01fF
C32971 VDD OR2X1_LOC_212/A 0.08fF
C32972 OR2X1_LOC_91/Y AND2X1_LOC_778/Y 0.02fF
C32973 OR2X1_LOC_160/B AND2X1_LOC_695/a_8_24# 0.01fF
C32974 AND2X1_LOC_548/a_8_24# OR2X1_LOC_816/A 0.01fF
C32975 AND2X1_LOC_683/a_8_24# OR2X1_LOC_161/B 0.01fF
C32976 OR2X1_LOC_427/A AND2X1_LOC_434/Y 0.07fF
C32977 OR2X1_LOC_482/Y OR2X1_LOC_36/Y 0.06fF
C32978 AND2X1_LOC_197/a_8_24# OR2X1_LOC_56/Y 0.01fF
C32979 AND2X1_LOC_801/a_8_24# AND2X1_LOC_434/Y 0.02fF
C32980 AND2X1_LOC_70/Y OR2X1_LOC_732/B 0.09fF
C32981 OR2X1_LOC_89/A OR2X1_LOC_16/A 0.01fF
C32982 OR2X1_LOC_574/A OR2X1_LOC_435/A 0.01fF
C32983 AND2X1_LOC_700/a_8_24# OR2X1_LOC_375/A 0.01fF
C32984 AND2X1_LOC_702/Y AND2X1_LOC_353/a_8_24# 0.01fF
C32985 AND2X1_LOC_40/Y OR2X1_LOC_840/A 0.03fF
C32986 AND2X1_LOC_621/Y OR2X1_LOC_59/Y 0.03fF
C32987 OR2X1_LOC_325/B OR2X1_LOC_468/Y 0.03fF
C32988 OR2X1_LOC_585/A OR2X1_LOC_13/Y 0.54fF
C32989 VDD OR2X1_LOC_687/Y 0.28fF
C32990 D_GATE_811 OR2X1_LOC_383/a_8_216# 0.40fF
C32991 AND2X1_LOC_729/B OR2X1_LOC_428/A 0.03fF
C32992 AND2X1_LOC_41/A AND2X1_LOC_305/a_8_24# -0.01fF
C32993 OR2X1_LOC_492/Y AND2X1_LOC_717/B 0.01fF
C32994 OR2X1_LOC_485/A OR2X1_LOC_13/a_8_216# 0.02fF
C32995 AND2X1_LOC_326/B OR2X1_LOC_6/A 0.02fF
C32996 OR2X1_LOC_108/Y OR2X1_LOC_26/Y 0.07fF
C32997 VDD AND2X1_LOC_650/Y 0.21fF
C32998 OR2X1_LOC_665/Y OR2X1_LOC_253/Y 0.06fF
C32999 OR2X1_LOC_223/A OR2X1_LOC_593/B 1.42fF
C33000 AND2X1_LOC_721/A AND2X1_LOC_247/a_8_24# 0.01fF
C33001 OR2X1_LOC_813/Y OR2X1_LOC_13/B 0.35fF
C33002 OR2X1_LOC_474/a_8_216# OR2X1_LOC_474/B 0.18fF
C33003 OR2X1_LOC_482/Y AND2X1_LOC_493/a_36_24# 0.06fF
C33004 AND2X1_LOC_167/a_8_24# OR2X1_LOC_161/A 0.06fF
C33005 OR2X1_LOC_600/A AND2X1_LOC_818/a_36_24# 0.00fF
C33006 AND2X1_LOC_668/a_8_24# OR2X1_LOC_59/Y 0.01fF
C33007 AND2X1_LOC_3/Y OR2X1_LOC_362/A 0.01fF
C33008 OR2X1_LOC_502/A AND2X1_LOC_11/Y 0.08fF
C33009 OR2X1_LOC_108/Y AND2X1_LOC_493/a_8_24# 0.05fF
C33010 OR2X1_LOC_8/Y AND2X1_LOC_838/a_8_24# 0.01fF
C33011 AND2X1_LOC_41/A OR2X1_LOC_738/A 0.02fF
C33012 OR2X1_LOC_364/A OR2X1_LOC_78/A 0.07fF
C33013 OR2X1_LOC_61/A OR2X1_LOC_476/B 0.04fF
C33014 AND2X1_LOC_19/Y OR2X1_LOC_87/A 0.23fF
C33015 OR2X1_LOC_473/a_8_216# OR2X1_LOC_493/A 0.02fF
C33016 OR2X1_LOC_216/A AND2X1_LOC_492/a_36_24# 0.00fF
C33017 OR2X1_LOC_185/Y OR2X1_LOC_78/A 0.13fF
C33018 OR2X1_LOC_188/Y OR2X1_LOC_471/Y 0.29fF
C33019 OR2X1_LOC_108/Y OR2X1_LOC_89/A 0.07fF
C33020 OR2X1_LOC_51/Y OR2X1_LOC_627/a_8_216# 0.01fF
C33021 OR2X1_LOC_816/Y OR2X1_LOC_36/Y 0.01fF
C33022 OR2X1_LOC_100/a_8_216# OR2X1_LOC_100/Y 0.01fF
C33023 OR2X1_LOC_421/A OR2X1_LOC_743/A 0.04fF
C33024 OR2X1_LOC_696/A OR2X1_LOC_62/A 0.03fF
C33025 OR2X1_LOC_107/a_36_216# AND2X1_LOC_560/B 0.00fF
C33026 OR2X1_LOC_8/Y OR2X1_LOC_827/Y 0.02fF
C33027 OR2X1_LOC_319/a_8_216# OR2X1_LOC_620/Y 0.01fF
C33028 OR2X1_LOC_441/Y AND2X1_LOC_811/a_8_24# 0.03fF
C33029 OR2X1_LOC_519/a_8_216# OR2X1_LOC_48/B 0.05fF
C33030 OR2X1_LOC_527/Y AND2X1_LOC_778/Y 0.29fF
C33031 OR2X1_LOC_820/A OR2X1_LOC_820/B 0.19fF
C33032 AND2X1_LOC_366/A OR2X1_LOC_753/A 0.09fF
C33033 VDD OR2X1_LOC_272/Y 0.53fF
C33034 OR2X1_LOC_18/Y AND2X1_LOC_805/Y 5.93fF
C33035 OR2X1_LOC_724/A OR2X1_LOC_446/B 0.02fF
C33036 AND2X1_LOC_19/Y AND2X1_LOC_19/a_8_24# 0.01fF
C33037 AND2X1_LOC_572/A OR2X1_LOC_92/Y 0.03fF
C33038 AND2X1_LOC_706/Y OR2X1_LOC_22/Y 0.03fF
C33039 OR2X1_LOC_223/A AND2X1_LOC_273/a_8_24# 0.01fF
C33040 OR2X1_LOC_500/A OR2X1_LOC_575/A 0.02fF
C33041 OR2X1_LOC_48/B OR2X1_LOC_433/Y 0.03fF
C33042 AND2X1_LOC_316/a_8_24# OR2X1_LOC_87/A 0.04fF
C33043 OR2X1_LOC_109/a_36_216# OR2X1_LOC_109/Y 0.00fF
C33044 AND2X1_LOC_560/a_36_24# OR2X1_LOC_47/Y 0.00fF
C33045 OR2X1_LOC_720/A OR2X1_LOC_721/Y 0.01fF
C33046 INPUT_3 AND2X1_LOC_820/a_36_24# 0.01fF
C33047 OR2X1_LOC_333/B OR2X1_LOC_78/B 0.03fF
C33048 OR2X1_LOC_276/B AND2X1_LOC_7/B 0.08fF
C33049 OR2X1_LOC_456/A AND2X1_LOC_18/Y 0.44fF
C33050 OR2X1_LOC_316/Y AND2X1_LOC_662/B 0.03fF
C33051 OR2X1_LOC_489/a_8_216# OR2X1_LOC_269/B 0.01fF
C33052 OR2X1_LOC_121/Y OR2X1_LOC_532/B 0.07fF
C33053 OR2X1_LOC_166/a_36_216# OR2X1_LOC_70/Y 0.00fF
C33054 OR2X1_LOC_128/B OR2X1_LOC_161/A 0.36fF
C33055 OR2X1_LOC_256/A OR2X1_LOC_12/Y 0.69fF
C33056 AND2X1_LOC_554/B AND2X1_LOC_474/A 0.23fF
C33057 OR2X1_LOC_476/Y AND2X1_LOC_92/Y 0.03fF
C33058 OR2X1_LOC_32/B AND2X1_LOC_573/A 0.15fF
C33059 VDD OR2X1_LOC_401/B 0.21fF
C33060 OR2X1_LOC_595/a_8_216# OR2X1_LOC_39/A 0.02fF
C33061 OR2X1_LOC_40/Y OR2X1_LOC_62/B 0.02fF
C33062 OR2X1_LOC_865/B OR2X1_LOC_865/a_36_216# 0.02fF
C33063 AND2X1_LOC_663/B OR2X1_LOC_700/a_36_216# 0.00fF
C33064 OR2X1_LOC_474/Y AND2X1_LOC_3/Y 0.03fF
C33065 AND2X1_LOC_276/a_36_24# OR2X1_LOC_52/B 0.01fF
C33066 OR2X1_LOC_58/Y OR2X1_LOC_22/Y 0.43fF
C33067 OR2X1_LOC_154/A OR2X1_LOC_377/A 0.22fF
C33068 AND2X1_LOC_811/Y AND2X1_LOC_212/Y 0.02fF
C33069 VDD OR2X1_LOC_606/Y 0.05fF
C33070 AND2X1_LOC_168/Y OR2X1_LOC_26/Y 0.06fF
C33071 OR2X1_LOC_6/B AND2X1_LOC_28/a_8_24# 0.03fF
C33072 AND2X1_LOC_41/a_8_24# AND2X1_LOC_53/Y 0.01fF
C33073 OR2X1_LOC_529/a_36_216# AND2X1_LOC_560/B 0.00fF
C33074 OR2X1_LOC_3/Y OR2X1_LOC_92/Y 2.08fF
C33075 AND2X1_LOC_392/A AND2X1_LOC_845/Y 0.07fF
C33076 OR2X1_LOC_518/Y AND2X1_LOC_222/Y 0.00fF
C33077 OR2X1_LOC_364/A OR2X1_LOC_602/A 0.02fF
C33078 OR2X1_LOC_114/B OR2X1_LOC_532/B 0.02fF
C33079 AND2X1_LOC_59/Y OR2X1_LOC_87/B 0.03fF
C33080 OR2X1_LOC_438/Y OR2X1_LOC_70/Y 0.10fF
C33081 OR2X1_LOC_449/B OR2X1_LOC_739/A 0.03fF
C33082 VDD AND2X1_LOC_801/B 0.16fF
C33083 AND2X1_LOC_605/Y OR2X1_LOC_64/Y 0.01fF
C33084 OR2X1_LOC_821/Y OR2X1_LOC_47/Y 0.03fF
C33085 OR2X1_LOC_757/A AND2X1_LOC_814/a_8_24# 0.01fF
C33086 AND2X1_LOC_721/Y OR2X1_LOC_419/Y 0.03fF
C33087 OR2X1_LOC_160/B OR2X1_LOC_780/A 0.01fF
C33088 OR2X1_LOC_8/Y AND2X1_LOC_835/a_8_24# 0.01fF
C33089 AND2X1_LOC_95/Y OR2X1_LOC_287/B 0.11fF
C33090 OR2X1_LOC_154/A OR2X1_LOC_203/Y 0.10fF
C33091 OR2X1_LOC_678/a_8_216# AND2X1_LOC_48/A 0.01fF
C33092 OR2X1_LOC_421/A OR2X1_LOC_409/B 0.00fF
C33093 AND2X1_LOC_259/Y OR2X1_LOC_18/Y 0.00fF
C33094 OR2X1_LOC_246/Y OR2X1_LOC_246/a_8_216# 0.01fF
C33095 AND2X1_LOC_51/Y OR2X1_LOC_392/A 0.00fF
C33096 OR2X1_LOC_316/Y AND2X1_LOC_634/a_8_24# 0.01fF
C33097 OR2X1_LOC_859/A OR2X1_LOC_561/Y 0.10fF
C33098 OR2X1_LOC_70/Y OR2X1_LOC_427/Y 0.01fF
C33099 OR2X1_LOC_299/Y OR2X1_LOC_619/Y 0.03fF
C33100 OR2X1_LOC_116/A AND2X1_LOC_3/Y 0.01fF
C33101 OR2X1_LOC_247/Y OR2X1_LOC_161/B 0.01fF
C33102 OR2X1_LOC_272/Y AND2X1_LOC_274/a_8_24# 0.09fF
C33103 OR2X1_LOC_654/A OR2X1_LOC_828/B 0.03fF
C33104 AND2X1_LOC_189/a_8_24# OR2X1_LOC_471/Y 0.02fF
C33105 OR2X1_LOC_283/Y AND2X1_LOC_859/Y 0.02fF
C33106 AND2X1_LOC_342/a_8_24# OR2X1_LOC_248/Y 0.10fF
C33107 AND2X1_LOC_537/Y AND2X1_LOC_857/Y 0.03fF
C33108 OR2X1_LOC_690/a_8_216# OR2X1_LOC_43/A -0.01fF
C33109 OR2X1_LOC_377/A OR2X1_LOC_856/a_8_216# 0.02fF
C33110 AND2X1_LOC_560/B AND2X1_LOC_361/A 0.01fF
C33111 OR2X1_LOC_43/A AND2X1_LOC_818/a_8_24# 0.01fF
C33112 OR2X1_LOC_364/A OR2X1_LOC_155/A 0.07fF
C33113 OR2X1_LOC_3/Y OR2X1_LOC_65/B 0.08fF
C33114 AND2X1_LOC_711/Y AND2X1_LOC_621/Y 0.01fF
C33115 OR2X1_LOC_337/A OR2X1_LOC_365/B 0.44fF
C33116 AND2X1_LOC_61/Y AND2X1_LOC_476/A 0.02fF
C33117 AND2X1_LOC_366/A AND2X1_LOC_845/Y 0.03fF
C33118 AND2X1_LOC_185/a_8_24# OR2X1_LOC_628/Y 0.01fF
C33119 OR2X1_LOC_666/A AND2X1_LOC_866/A 0.03fF
C33120 OR2X1_LOC_185/Y OR2X1_LOC_155/A 0.07fF
C33121 OR2X1_LOC_76/A OR2X1_LOC_737/A 0.07fF
C33122 OR2X1_LOC_132/a_36_216# AND2X1_LOC_227/Y 0.00fF
C33123 OR2X1_LOC_538/A OR2X1_LOC_532/B 0.04fF
C33124 OR2X1_LOC_70/Y AND2X1_LOC_621/Y 0.03fF
C33125 OR2X1_LOC_633/Y OR2X1_LOC_97/a_8_216# 0.04fF
C33126 AND2X1_LOC_22/Y OR2X1_LOC_228/Y 0.81fF
C33127 OR2X1_LOC_217/Y AND2X1_LOC_3/Y 0.01fF
C33128 OR2X1_LOC_449/B OR2X1_LOC_269/B 0.03fF
C33129 OR2X1_LOC_654/A OR2X1_LOC_835/B 0.07fF
C33130 VDD OR2X1_LOC_786/Y 1.70fF
C33131 OR2X1_LOC_139/A OR2X1_LOC_68/B 0.03fF
C33132 OR2X1_LOC_160/B D_INPUT_1 0.72fF
C33133 AND2X1_LOC_554/B OR2X1_LOC_85/A 0.14fF
C33134 OR2X1_LOC_273/Y OR2X1_LOC_316/Y 0.03fF
C33135 AND2X1_LOC_729/Y AND2X1_LOC_797/A 0.00fF
C33136 AND2X1_LOC_213/B AND2X1_LOC_779/Y 0.00fF
C33137 OR2X1_LOC_273/Y OR2X1_LOC_595/a_36_216# 0.03fF
C33138 OR2X1_LOC_470/B OR2X1_LOC_467/a_8_216# 0.01fF
C33139 OR2X1_LOC_216/A D_INPUT_0 0.01fF
C33140 OR2X1_LOC_482/Y OR2X1_LOC_419/Y 0.03fF
C33141 OR2X1_LOC_160/A OR2X1_LOC_473/Y 0.05fF
C33142 AND2X1_LOC_101/a_8_24# OR2X1_LOC_278/Y 0.01fF
C33143 OR2X1_LOC_527/Y AND2X1_LOC_624/A 0.07fF
C33144 OR2X1_LOC_76/Y OR2X1_LOC_445/a_8_216# 0.40fF
C33145 OR2X1_LOC_185/Y OR2X1_LOC_392/a_8_216# 0.01fF
C33146 OR2X1_LOC_121/B OR2X1_LOC_739/A 0.03fF
C33147 VDD OR2X1_LOC_747/Y 0.12fF
C33148 OR2X1_LOC_307/B AND2X1_LOC_47/Y 0.01fF
C33149 OR2X1_LOC_97/B AND2X1_LOC_42/B 0.15fF
C33150 AND2X1_LOC_347/B AND2X1_LOC_848/A 0.05fF
C33151 OR2X1_LOC_233/a_36_216# OR2X1_LOC_753/A 0.01fF
C33152 VDD OR2X1_LOC_644/A 0.05fF
C33153 OR2X1_LOC_99/B OR2X1_LOC_375/A 0.01fF
C33154 OR2X1_LOC_778/A OR2X1_LOC_203/Y 0.01fF
C33155 AND2X1_LOC_680/a_36_24# OR2X1_LOC_506/A 0.00fF
C33156 OR2X1_LOC_304/Y OR2X1_LOC_36/Y 0.43fF
C33157 AND2X1_LOC_35/Y AND2X1_LOC_853/a_36_24# 0.00fF
C33158 OR2X1_LOC_161/B OR2X1_LOC_364/Y 0.03fF
C33159 AND2X1_LOC_512/a_8_24# OR2X1_LOC_743/A 0.01fF
C33160 D_INPUT_3 OR2X1_LOC_517/A 0.03fF
C33161 OR2X1_LOC_748/A AND2X1_LOC_847/a_36_24# 0.00fF
C33162 OR2X1_LOC_122/Y OR2X1_LOC_47/Y 0.02fF
C33163 AND2X1_LOC_137/a_36_24# OR2X1_LOC_517/A 0.01fF
C33164 AND2X1_LOC_716/Y AND2X1_LOC_866/A 0.02fF
C33165 OR2X1_LOC_280/Y OR2X1_LOC_485/A 0.06fF
C33166 OR2X1_LOC_654/a_36_216# OR2X1_LOC_68/B 0.00fF
C33167 AND2X1_LOC_390/B AND2X1_LOC_337/B 0.02fF
C33168 AND2X1_LOC_477/A AND2X1_LOC_470/B 0.83fF
C33169 OR2X1_LOC_520/Y AND2X1_LOC_518/a_36_24# 0.00fF
C33170 OR2X1_LOC_64/Y AND2X1_LOC_361/A 0.07fF
C33171 OR2X1_LOC_679/A OR2X1_LOC_679/B 0.33fF
C33172 OR2X1_LOC_88/Y OR2X1_LOC_131/a_36_216# 0.00fF
C33173 OR2X1_LOC_504/Y AND2X1_LOC_621/Y 0.03fF
C33174 AND2X1_LOC_863/Y AND2X1_LOC_662/B 0.00fF
C33175 OR2X1_LOC_121/B OR2X1_LOC_269/B 0.10fF
C33176 AND2X1_LOC_810/Y OR2X1_LOC_48/B 0.07fF
C33177 AND2X1_LOC_12/Y OR2X1_LOC_532/B 9.84fF
C33178 OR2X1_LOC_462/B AND2X1_LOC_519/a_8_24# 0.01fF
C33179 OR2X1_LOC_642/a_8_216# AND2X1_LOC_48/A 0.01fF
C33180 OR2X1_LOC_739/B OR2X1_LOC_223/a_8_216# 0.14fF
C33181 AND2X1_LOC_715/a_8_24# AND2X1_LOC_727/A 0.01fF
C33182 AND2X1_LOC_95/Y OR2X1_LOC_436/Y 0.04fF
C33183 OR2X1_LOC_675/A OR2X1_LOC_733/B 0.01fF
C33184 AND2X1_LOC_343/a_8_24# OR2X1_LOC_64/Y 0.00fF
C33185 OR2X1_LOC_45/B AND2X1_LOC_449/a_8_24# 0.02fF
C33186 OR2X1_LOC_678/Y OR2X1_LOC_512/a_8_216# 0.02fF
C33187 AND2X1_LOC_804/A OR2X1_LOC_142/Y 0.05fF
C33188 OR2X1_LOC_839/a_36_216# OR2X1_LOC_375/A 0.00fF
C33189 OR2X1_LOC_19/B AND2X1_LOC_823/a_36_24# 0.00fF
C33190 OR2X1_LOC_432/a_8_216# AND2X1_LOC_648/B -0.00fF
C33191 AND2X1_LOC_539/a_8_24# OR2X1_LOC_43/A 0.01fF
C33192 OR2X1_LOC_222/a_8_216# OR2X1_LOC_405/Y 0.04fF
C33193 D_INPUT_0 OR2X1_LOC_44/Y 0.03fF
C33194 OR2X1_LOC_636/B AND2X1_LOC_51/Y 0.01fF
C33195 OR2X1_LOC_45/B OR2X1_LOC_183/a_8_216# 0.09fF
C33196 AND2X1_LOC_808/A AND2X1_LOC_808/a_8_24# 0.01fF
C33197 AND2X1_LOC_826/a_8_24# OR2X1_LOC_6/A 0.17fF
C33198 OR2X1_LOC_91/A AND2X1_LOC_222/Y 0.03fF
C33199 OR2X1_LOC_316/Y OR2X1_LOC_75/Y 0.03fF
C33200 OR2X1_LOC_83/A INPUT_1 0.03fF
C33201 AND2X1_LOC_91/B OR2X1_LOC_168/Y 0.09fF
C33202 OR2X1_LOC_849/A AND2X1_LOC_15/a_8_24# 0.01fF
C33203 OR2X1_LOC_481/Y AND2X1_LOC_663/B 0.26fF
C33204 OR2X1_LOC_276/B OR2X1_LOC_805/A 0.07fF
C33205 OR2X1_LOC_78/A OR2X1_LOC_568/A 0.07fF
C33206 OR2X1_LOC_485/A OR2X1_LOC_22/Y 9.27fF
C33207 INPUT_3 D_INPUT_1 0.04fF
C33208 OR2X1_LOC_78/A OR2X1_LOC_578/B 0.00fF
C33209 OR2X1_LOC_416/Y OR2X1_LOC_27/a_8_216# 0.01fF
C33210 GATE_366 AND2X1_LOC_866/A 0.07fF
C33211 OR2X1_LOC_377/A AND2X1_LOC_6/a_8_24# 0.01fF
C33212 OR2X1_LOC_421/A OR2X1_LOC_589/a_36_216# 0.00fF
C33213 AND2X1_LOC_651/a_8_24# OR2X1_LOC_70/A 0.01fF
C33214 AND2X1_LOC_42/B OR2X1_LOC_814/A 0.07fF
C33215 AND2X1_LOC_59/Y OR2X1_LOC_795/a_8_216# 0.01fF
C33216 OR2X1_LOC_405/A OR2X1_LOC_493/Y 0.02fF
C33217 AND2X1_LOC_476/A AND2X1_LOC_852/Y 0.07fF
C33218 OR2X1_LOC_532/B AND2X1_LOC_79/Y 0.01fF
C33219 AND2X1_LOC_562/B AND2X1_LOC_793/B 1.16fF
C33220 OR2X1_LOC_653/A AND2X1_LOC_109/a_36_24# 0.00fF
C33221 D_INPUT_0 OR2X1_LOC_20/a_8_216# 0.01fF
C33222 AND2X1_LOC_337/B AND2X1_LOC_863/Y 0.01fF
C33223 OR2X1_LOC_312/Y AND2X1_LOC_866/A 0.03fF
C33224 OR2X1_LOC_182/B OR2X1_LOC_182/a_36_216# 0.00fF
C33225 OR2X1_LOC_618/a_36_216# D_INPUT_1 0.00fF
C33226 AND2X1_LOC_341/a_8_24# OR2X1_LOC_171/Y 0.08fF
C33227 AND2X1_LOC_483/Y AND2X1_LOC_624/A 0.03fF
C33228 VDD OR2X1_LOC_181/Y 0.19fF
C33229 OR2X1_LOC_833/B OR2X1_LOC_675/Y 0.02fF
C33230 VDD OR2X1_LOC_248/A -0.00fF
C33231 OR2X1_LOC_92/Y AND2X1_LOC_772/a_8_24# 0.15fF
C33232 OR2X1_LOC_272/Y OR2X1_LOC_256/A 0.01fF
C33233 AND2X1_LOC_512/Y OR2X1_LOC_533/a_36_216# -0.01fF
C33234 OR2X1_LOC_6/B AND2X1_LOC_750/a_36_24# 0.01fF
C33235 AND2X1_LOC_715/Y OR2X1_LOC_312/a_36_216# 0.01fF
C33236 AND2X1_LOC_44/Y OR2X1_LOC_259/A 0.01fF
C33237 OR2X1_LOC_590/a_8_216# OR2X1_LOC_375/A 0.01fF
C33238 OR2X1_LOC_45/B OR2X1_LOC_304/a_8_216# 0.01fF
C33239 AND2X1_LOC_610/a_8_24# AND2X1_LOC_647/B 0.02fF
C33240 OR2X1_LOC_631/B AND2X1_LOC_72/B 0.05fF
C33241 OR2X1_LOC_7/a_8_216# OR2X1_LOC_7/Y 0.01fF
C33242 OR2X1_LOC_375/A OR2X1_LOC_543/a_36_216# 0.00fF
C33243 OR2X1_LOC_45/B AND2X1_LOC_712/a_8_24# 0.01fF
C33244 AND2X1_LOC_722/A OR2X1_LOC_13/B 0.07fF
C33245 OR2X1_LOC_619/Y OR2X1_LOC_534/Y 0.03fF
C33246 AND2X1_LOC_769/Y AND2X1_LOC_771/a_8_24# 0.19fF
C33247 OR2X1_LOC_377/A OR2X1_LOC_198/A 0.01fF
C33248 OR2X1_LOC_243/a_36_216# OR2X1_LOC_62/B 0.00fF
C33249 OR2X1_LOC_709/A AND2X1_LOC_7/B 0.01fF
C33250 AND2X1_LOC_64/Y OR2X1_LOC_629/B 0.00fF
C33251 OR2X1_LOC_696/A OR2X1_LOC_8/Y 0.03fF
C33252 OR2X1_LOC_19/B AND2X1_LOC_821/a_36_24# 0.01fF
C33253 AND2X1_LOC_43/B OR2X1_LOC_80/A 0.01fF
C33254 OR2X1_LOC_655/B D_INPUT_0 0.09fF
C33255 AND2X1_LOC_564/A AND2X1_LOC_476/Y 0.07fF
C33256 AND2X1_LOC_41/A AND2X1_LOC_36/Y 0.62fF
C33257 AND2X1_LOC_787/A AND2X1_LOC_180/a_8_24# 0.04fF
C33258 AND2X1_LOC_776/Y VDD 0.11fF
C33259 OR2X1_LOC_167/a_8_216# OR2X1_LOC_16/A 0.01fF
C33260 AND2X1_LOC_831/Y INPUT_1 0.01fF
C33261 AND2X1_LOC_562/a_8_24# OR2X1_LOC_604/A 0.05fF
C33262 OR2X1_LOC_181/B OR2X1_LOC_181/a_8_216# 0.01fF
C33263 AND2X1_LOC_727/Y VDD 0.24fF
C33264 AND2X1_LOC_43/B AND2X1_LOC_419/a_8_24# 0.04fF
C33265 OR2X1_LOC_203/Y OR2X1_LOC_560/A 0.00fF
C33266 OR2X1_LOC_250/a_8_216# OR2X1_LOC_13/B 0.02fF
C33267 OR2X1_LOC_43/A OR2X1_LOC_534/a_8_216# 0.02fF
C33268 AND2X1_LOC_212/Y AND2X1_LOC_469/a_8_24# 0.03fF
C33269 AND2X1_LOC_721/Y OR2X1_LOC_604/A 0.01fF
C33270 OR2X1_LOC_113/a_8_216# OR2X1_LOC_66/A 0.02fF
C33271 AND2X1_LOC_392/A OR2X1_LOC_310/a_36_216# 0.01fF
C33272 OR2X1_LOC_807/A OR2X1_LOC_580/A 0.08fF
C33273 OR2X1_LOC_154/A OR2X1_LOC_732/A 0.09fF
C33274 AND2X1_LOC_70/Y AND2X1_LOC_7/B 0.15fF
C33275 OR2X1_LOC_329/B AND2X1_LOC_241/a_8_24# -0.01fF
C33276 AND2X1_LOC_18/Y OR2X1_LOC_161/B 0.21fF
C33277 AND2X1_LOC_719/Y OR2X1_LOC_482/a_8_216# 0.00fF
C33278 VDD AND2X1_LOC_255/a_8_24# -0.00fF
C33279 OR2X1_LOC_60/Y OR2X1_LOC_12/Y 0.01fF
C33280 VDD OR2X1_LOC_569/B 0.20fF
C33281 OR2X1_LOC_244/A D_INPUT_1 0.07fF
C33282 OR2X1_LOC_6/B OR2X1_LOC_151/A 0.07fF
C33283 OR2X1_LOC_599/A OR2X1_LOC_13/B 0.00fF
C33284 D_INPUT_0 OR2X1_LOC_205/Y 0.00fF
C33285 OR2X1_LOC_56/A AND2X1_LOC_786/Y 0.15fF
C33286 OR2X1_LOC_27/Y OR2X1_LOC_68/B 0.01fF
C33287 OR2X1_LOC_154/A OR2X1_LOC_539/B 0.07fF
C33288 OR2X1_LOC_87/A OR2X1_LOC_723/B 0.07fF
C33289 OR2X1_LOC_506/A OR2X1_LOC_354/a_8_216# 0.05fF
C33290 AND2X1_LOC_59/Y OR2X1_LOC_333/A 0.43fF
C33291 OR2X1_LOC_269/B OR2X1_LOC_195/a_8_216# 0.09fF
C33292 OR2X1_LOC_158/A AND2X1_LOC_366/a_8_24# 0.17fF
C33293 AND2X1_LOC_592/Y AND2X1_LOC_447/Y 0.02fF
C33294 AND2X1_LOC_2/Y AND2X1_LOC_40/a_36_24# 0.01fF
C33295 AND2X1_LOC_70/a_8_24# AND2X1_LOC_40/a_8_24# 0.23fF
C33296 OR2X1_LOC_45/B OR2X1_LOC_164/Y 0.00fF
C33297 OR2X1_LOC_737/A OR2X1_LOC_722/B 0.02fF
C33298 AND2X1_LOC_191/Y AND2X1_LOC_740/a_36_24# 0.01fF
C33299 OR2X1_LOC_506/Y AND2X1_LOC_41/A 0.07fF
C33300 OR2X1_LOC_696/A OR2X1_LOC_67/A 0.03fF
C33301 AND2X1_LOC_388/Y OR2X1_LOC_166/a_8_216# 0.01fF
C33302 AND2X1_LOC_547/Y AND2X1_LOC_565/B 0.15fF
C33303 OR2X1_LOC_702/A OR2X1_LOC_515/a_8_216# 0.01fF
C33304 OR2X1_LOC_631/B AND2X1_LOC_36/Y 0.02fF
C33305 VDD OR2X1_LOC_622/A 0.00fF
C33306 OR2X1_LOC_440/a_8_216# OR2X1_LOC_66/A 0.01fF
C33307 OR2X1_LOC_860/a_8_216# OR2X1_LOC_392/B 0.04fF
C33308 AND2X1_LOC_3/Y OR2X1_LOC_771/B 0.04fF
C33309 AND2X1_LOC_785/a_36_24# OR2X1_LOC_18/Y 0.00fF
C33310 OR2X1_LOC_323/A OR2X1_LOC_316/Y 0.00fF
C33311 OR2X1_LOC_9/Y INPUT_0 0.03fF
C33312 INPUT_0 AND2X1_LOC_193/Y 0.03fF
C33313 AND2X1_LOC_362/B AND2X1_LOC_474/A 0.03fF
C33314 D_INPUT_0 OR2X1_LOC_750/Y 0.79fF
C33315 OR2X1_LOC_508/A OR2X1_LOC_506/Y 0.08fF
C33316 VDD OR2X1_LOC_467/A 0.20fF
C33317 OR2X1_LOC_314/a_8_216# OR2X1_LOC_12/Y 0.01fF
C33318 OR2X1_LOC_653/A OR2X1_LOC_390/B 0.16fF
C33319 OR2X1_LOC_604/A OR2X1_LOC_816/Y 0.00fF
C33320 AND2X1_LOC_388/Y AND2X1_LOC_436/a_36_24# 0.00fF
C33321 AND2X1_LOC_57/Y OR2X1_LOC_864/A 0.81fF
C33322 OR2X1_LOC_696/A AND2X1_LOC_374/Y 0.01fF
C33323 OR2X1_LOC_335/A OR2X1_LOC_87/A 0.01fF
C33324 AND2X1_LOC_59/Y OR2X1_LOC_392/B 0.03fF
C33325 AND2X1_LOC_65/A OR2X1_LOC_475/B 0.40fF
C33326 OR2X1_LOC_842/A OR2X1_LOC_78/A 0.04fF
C33327 AND2X1_LOC_12/Y OR2X1_LOC_865/A 0.06fF
C33328 AND2X1_LOC_76/Y OR2X1_LOC_522/a_36_216# 0.00fF
C33329 OR2X1_LOC_696/A OR2X1_LOC_52/B 0.14fF
C33330 OR2X1_LOC_696/A OR2X1_LOC_672/Y 0.04fF
C33331 AND2X1_LOC_56/B OR2X1_LOC_415/Y 0.02fF
C33332 OR2X1_LOC_380/a_8_216# OR2X1_LOC_25/Y 0.01fF
C33333 AND2X1_LOC_522/a_8_24# OR2X1_LOC_161/A 0.01fF
C33334 OR2X1_LOC_623/B OR2X1_LOC_596/A 0.03fF
C33335 OR2X1_LOC_653/B OR2X1_LOC_653/Y 0.03fF
C33336 VDD OR2X1_LOC_234/Y 0.10fF
C33337 OR2X1_LOC_435/B AND2X1_LOC_18/Y 0.01fF
C33338 OR2X1_LOC_658/a_8_216# OR2X1_LOC_66/A 0.02fF
C33339 AND2X1_LOC_539/Y OR2X1_LOC_44/Y 0.03fF
C33340 OR2X1_LOC_426/A OR2X1_LOC_765/Y 0.01fF
C33341 OR2X1_LOC_326/B OR2X1_LOC_151/A 0.02fF
C33342 OR2X1_LOC_359/a_8_216# OR2X1_LOC_756/B 0.02fF
C33343 OR2X1_LOC_696/A AND2X1_LOC_489/Y 0.03fF
C33344 OR2X1_LOC_756/B OR2X1_LOC_35/a_8_216# 0.01fF
C33345 AND2X1_LOC_738/B OR2X1_LOC_524/Y 0.10fF
C33346 AND2X1_LOC_64/Y OR2X1_LOC_84/B 0.07fF
C33347 AND2X1_LOC_716/Y OR2X1_LOC_40/Y 0.17fF
C33348 OR2X1_LOC_193/Y AND2X1_LOC_7/B 0.05fF
C33349 AND2X1_LOC_714/B OR2X1_LOC_48/B 0.01fF
C33350 AND2X1_LOC_541/a_8_24# AND2X1_LOC_361/A -0.03fF
C33351 OR2X1_LOC_500/A OR2X1_LOC_161/B 0.01fF
C33352 OR2X1_LOC_697/Y OR2X1_LOC_51/Y 0.42fF
C33353 AND2X1_LOC_794/B AND2X1_LOC_468/B 0.10fF
C33354 AND2X1_LOC_50/Y AND2X1_LOC_95/a_8_24# 0.11fF
C33355 OR2X1_LOC_326/B AND2X1_LOC_322/a_8_24# 0.02fF
C33356 AND2X1_LOC_658/B OR2X1_LOC_438/Y 0.14fF
C33357 AND2X1_LOC_576/Y OR2X1_LOC_816/A 0.07fF
C33358 AND2X1_LOC_658/B AND2X1_LOC_865/a_8_24# 0.18fF
C33359 VDD AND2X1_LOC_404/A 0.21fF
C33360 OR2X1_LOC_709/A OR2X1_LOC_805/A 0.00fF
C33361 AND2X1_LOC_721/a_8_24# OR2X1_LOC_494/Y 0.04fF
C33362 AND2X1_LOC_388/Y OR2X1_LOC_619/Y 0.03fF
C33363 OR2X1_LOC_61/Y AND2X1_LOC_18/Y 0.04fF
C33364 OR2X1_LOC_664/Y OR2X1_LOC_294/Y 0.03fF
C33365 OR2X1_LOC_254/B OR2X1_LOC_736/Y 0.15fF
C33366 AND2X1_LOC_17/Y AND2X1_LOC_7/B 0.65fF
C33367 AND2X1_LOC_339/B AND2X1_LOC_655/A 0.05fF
C33368 AND2X1_LOC_367/A OR2X1_LOC_91/A 0.03fF
C33369 OR2X1_LOC_596/Y OR2X1_LOC_161/B 0.02fF
C33370 VDD OR2X1_LOC_59/a_8_216# 0.00fF
C33371 OR2X1_LOC_160/B OR2X1_LOC_737/A 0.07fF
C33372 VDD OR2X1_LOC_725/B 0.00fF
C33373 OR2X1_LOC_64/Y OR2X1_LOC_387/A 0.02fF
C33374 OR2X1_LOC_309/Y AND2X1_LOC_662/B 0.27fF
C33375 OR2X1_LOC_744/A OR2X1_LOC_763/a_8_216# 0.01fF
C33376 OR2X1_LOC_403/a_8_216# AND2X1_LOC_36/Y 0.01fF
C33377 OR2X1_LOC_305/Y AND2X1_LOC_774/A 0.05fF
C33378 OR2X1_LOC_158/A OR2X1_LOC_265/Y 0.07fF
C33379 OR2X1_LOC_318/Y AND2X1_LOC_70/Y 0.03fF
C33380 AND2X1_LOC_22/Y AND2X1_LOC_386/a_8_24# 0.02fF
C33381 OR2X1_LOC_160/B AND2X1_LOC_95/Y 5.91fF
C33382 AND2X1_LOC_866/A OR2X1_LOC_13/B 0.07fF
C33383 AND2X1_LOC_661/A AND2X1_LOC_810/B 0.04fF
C33384 OR2X1_LOC_26/Y OR2X1_LOC_373/Y 0.31fF
C33385 AND2X1_LOC_554/a_36_24# OR2X1_LOC_89/A 0.00fF
C33386 OR2X1_LOC_415/a_8_216# OR2X1_LOC_395/Y 0.01fF
C33387 OR2X1_LOC_248/Y OR2X1_LOC_12/Y 0.10fF
C33388 OR2X1_LOC_329/B OR2X1_LOC_92/Y 15.03fF
C33389 OR2X1_LOC_49/A OR2X1_LOC_585/A 0.45fF
C33390 AND2X1_LOC_264/a_8_24# OR2X1_LOC_595/A 0.08fF
C33391 VDD AND2X1_LOC_468/B 0.10fF
C33392 OR2X1_LOC_666/A AND2X1_LOC_843/Y 0.00fF
C33393 AND2X1_LOC_719/Y AND2X1_LOC_859/a_8_24# 0.00fF
C33394 AND2X1_LOC_853/Y OR2X1_LOC_16/A 0.03fF
C33395 OR2X1_LOC_44/Y AND2X1_LOC_771/B 0.01fF
C33396 AND2X1_LOC_290/a_36_24# OR2X1_LOC_66/A 0.01fF
C33397 OR2X1_LOC_319/B OR2X1_LOC_703/A 0.01fF
C33398 OR2X1_LOC_58/Y OR2X1_LOC_39/A 0.04fF
C33399 OR2X1_LOC_502/A AND2X1_LOC_306/a_36_24# 0.02fF
C33400 AND2X1_LOC_658/B AND2X1_LOC_621/Y 0.02fF
C33401 OR2X1_LOC_106/A OR2X1_LOC_595/A 0.18fF
C33402 OR2X1_LOC_620/Y OR2X1_LOC_78/B 0.07fF
C33403 OR2X1_LOC_89/A OR2X1_LOC_373/Y 0.06fF
C33404 OR2X1_LOC_206/a_8_216# AND2X1_LOC_7/B 0.01fF
C33405 OR2X1_LOC_617/Y GATE_579 0.04fF
C33406 OR2X1_LOC_744/A OR2X1_LOC_278/Y 0.03fF
C33407 VDD OR2X1_LOC_828/B 0.11fF
C33408 AND2X1_LOC_294/a_36_24# OR2X1_LOC_12/Y 0.01fF
C33409 OR2X1_LOC_468/A OR2X1_LOC_539/Y 0.27fF
C33410 OR2X1_LOC_436/Y OR2X1_LOC_175/a_8_216# 0.01fF
C33411 OR2X1_LOC_40/Y GATE_366 0.03fF
C33412 D_INPUT_5 AND2X1_LOC_2/a_8_24# 0.05fF
C33413 AND2X1_LOC_70/Y OR2X1_LOC_805/A 0.19fF
C33414 AND2X1_LOC_214/A OR2X1_LOC_48/B 0.02fF
C33415 OR2X1_LOC_287/B OR2X1_LOC_343/a_36_216# 0.00fF
C33416 AND2X1_LOC_758/a_36_24# OR2X1_LOC_680/A 0.01fF
C33417 VDD OR2X1_LOC_835/B 0.02fF
C33418 OR2X1_LOC_703/A OR2X1_LOC_212/a_8_216# 0.01fF
C33419 OR2X1_LOC_34/B OR2X1_LOC_338/A 0.03fF
C33420 OR2X1_LOC_604/A OR2X1_LOC_748/A 0.04fF
C33421 AND2X1_LOC_112/a_8_24# OR2X1_LOC_6/A 0.17fF
C33422 OR2X1_LOC_808/A OR2X1_LOC_794/A 0.01fF
C33423 OR2X1_LOC_676/Y OR2X1_LOC_793/A 0.02fF
C33424 OR2X1_LOC_122/a_8_216# OR2X1_LOC_67/A 0.01fF
C33425 AND2X1_LOC_182/a_8_24# AND2X1_LOC_211/B 0.02fF
C33426 AND2X1_LOC_22/Y OR2X1_LOC_76/A 0.50fF
C33427 AND2X1_LOC_392/A AND2X1_LOC_784/A 0.17fF
C33428 OR2X1_LOC_532/B OR2X1_LOC_356/B 0.18fF
C33429 AND2X1_LOC_711/A OR2X1_LOC_44/Y 0.15fF
C33430 OR2X1_LOC_145/a_8_216# AND2X1_LOC_658/A 0.03fF
C33431 AND2X1_LOC_124/a_36_24# OR2X1_LOC_56/A 0.00fF
C33432 AND2X1_LOC_861/B OR2X1_LOC_18/Y 0.01fF
C33433 AND2X1_LOC_184/a_8_24# AND2X1_LOC_292/a_8_24# 0.23fF
C33434 OR2X1_LOC_40/Y OR2X1_LOC_312/Y 0.03fF
C33435 OR2X1_LOC_670/a_8_216# OR2X1_LOC_51/Y 0.01fF
C33436 AND2X1_LOC_367/A AND2X1_LOC_573/A 0.10fF
C33437 OR2X1_LOC_516/a_8_216# AND2X1_LOC_469/B 0.01fF
C33438 AND2X1_LOC_773/Y AND2X1_LOC_307/Y 0.03fF
C33439 AND2X1_LOC_40/Y OR2X1_LOC_805/a_8_216# 0.01fF
C33440 OR2X1_LOC_804/A OR2X1_LOC_777/B 0.02fF
C33441 OR2X1_LOC_154/A OR2X1_LOC_78/B 0.38fF
C33442 OR2X1_LOC_317/a_8_216# OR2X1_LOC_739/A 0.01fF
C33443 AND2X1_LOC_777/a_8_24# OR2X1_LOC_56/A 0.01fF
C33444 OR2X1_LOC_814/A AND2X1_LOC_224/a_8_24# 0.10fF
C33445 AND2X1_LOC_12/Y OR2X1_LOC_391/A 0.19fF
C33446 OR2X1_LOC_51/B D_INPUT_6 0.01fF
C33447 OR2X1_LOC_856/A AND2X1_LOC_51/Y 0.02fF
C33448 INPUT_0 OR2X1_LOC_96/B 0.03fF
C33449 OR2X1_LOC_485/Y OR2X1_LOC_485/A 0.01fF
C33450 OR2X1_LOC_154/A AND2X1_LOC_103/a_36_24# 0.00fF
C33451 AND2X1_LOC_40/Y OR2X1_LOC_362/B 0.45fF
C33452 OR2X1_LOC_46/A OR2X1_LOC_428/A 0.02fF
C33453 AND2X1_LOC_639/A OR2X1_LOC_18/a_8_216# 0.03fF
C33454 OR2X1_LOC_45/B AND2X1_LOC_633/Y 0.03fF
C33455 AND2X1_LOC_803/B OR2X1_LOC_189/Y 0.03fF
C33456 OR2X1_LOC_311/Y AND2X1_LOC_774/A 0.03fF
C33457 OR2X1_LOC_170/Y OR2X1_LOC_303/B 0.20fF
C33458 OR2X1_LOC_640/a_8_216# OR2X1_LOC_640/A 0.18fF
C33459 AND2X1_LOC_133/a_8_24# AND2X1_LOC_44/Y 0.07fF
C33460 OR2X1_LOC_631/B OR2X1_LOC_630/Y 0.04fF
C33461 OR2X1_LOC_161/A OR2X1_LOC_712/a_8_216# 0.06fF
C33462 OR2X1_LOC_840/A AND2X1_LOC_43/B 0.08fF
C33463 OR2X1_LOC_741/Y OR2X1_LOC_564/A 0.02fF
C33464 OR2X1_LOC_160/A OR2X1_LOC_469/Y 3.37fF
C33465 AND2X1_LOC_583/a_8_24# OR2X1_LOC_87/A 0.15fF
C33466 AND2X1_LOC_339/B AND2X1_LOC_350/Y 0.03fF
C33467 OR2X1_LOC_132/Y OR2X1_LOC_26/Y 0.04fF
C33468 AND2X1_LOC_792/Y AND2X1_LOC_793/a_8_24# 0.04fF
C33469 AND2X1_LOC_64/Y OR2X1_LOC_651/A 0.19fF
C33470 OR2X1_LOC_3/Y OR2X1_LOC_600/A 0.35fF
C33471 OR2X1_LOC_476/B OR2X1_LOC_390/A 0.00fF
C33472 AND2X1_LOC_8/Y OR2X1_LOC_520/a_36_216# 0.00fF
C33473 OR2X1_LOC_777/B OR2X1_LOC_723/A 0.09fF
C33474 OR2X1_LOC_100/Y AND2X1_LOC_59/Y 0.12fF
C33475 AND2X1_LOC_713/a_36_24# OR2X1_LOC_64/Y 0.00fF
C33476 AND2X1_LOC_568/a_8_24# OR2X1_LOC_600/A 0.03fF
C33477 OR2X1_LOC_696/A OR2X1_LOC_619/a_36_216# 0.00fF
C33478 AND2X1_LOC_803/B OR2X1_LOC_152/Y 0.02fF
C33479 AND2X1_LOC_538/Y AND2X1_LOC_774/A 0.11fF
C33480 OR2X1_LOC_45/B D_INPUT_0 0.11fF
C33481 OR2X1_LOC_337/a_36_216# OR2X1_LOC_87/A 0.00fF
C33482 OR2X1_LOC_577/a_8_216# OR2X1_LOC_577/B 0.05fF
C33483 AND2X1_LOC_206/Y AND2X1_LOC_215/a_36_24# 0.01fF
C33484 AND2X1_LOC_112/a_36_24# OR2X1_LOC_74/A 0.00fF
C33485 AND2X1_LOC_554/B OR2X1_LOC_51/Y 0.02fF
C33486 AND2X1_LOC_851/A OR2X1_LOC_39/A 0.03fF
C33487 OR2X1_LOC_68/B OR2X1_LOC_558/a_8_216# 0.01fF
C33488 AND2X1_LOC_51/Y OR2X1_LOC_730/A 0.04fF
C33489 OR2X1_LOC_680/Y OR2X1_LOC_51/Y 0.23fF
C33490 AND2X1_LOC_53/Y AND2X1_LOC_44/Y 0.02fF
C33491 AND2X1_LOC_42/B OR2X1_LOC_244/Y 0.17fF
C33492 OR2X1_LOC_437/A AND2X1_LOC_796/A 0.00fF
C33493 OR2X1_LOC_451/B INPUT_6 0.00fF
C33494 OR2X1_LOC_468/A AND2X1_LOC_176/a_8_24# 0.01fF
C33495 AND2X1_LOC_22/Y OR2X1_LOC_436/Y 0.01fF
C33496 AND2X1_LOC_40/Y OR2X1_LOC_468/Y 0.85fF
C33497 AND2X1_LOC_578/A OR2X1_LOC_56/A 0.03fF
C33498 AND2X1_LOC_227/Y OR2X1_LOC_428/A 0.02fF
C33499 OR2X1_LOC_755/a_8_216# OR2X1_LOC_757/Y 0.40fF
C33500 OR2X1_LOC_490/Y OR2X1_LOC_91/A 0.14fF
C33501 OR2X1_LOC_185/A OR2X1_LOC_243/A 0.02fF
C33502 OR2X1_LOC_91/A OR2X1_LOC_74/A 0.21fF
C33503 AND2X1_LOC_711/Y OR2X1_LOC_59/Y 0.01fF
C33504 OR2X1_LOC_440/A AND2X1_LOC_604/a_8_24# 0.02fF
C33505 OR2X1_LOC_93/Y OR2X1_LOC_54/Y 0.02fF
C33506 AND2X1_LOC_535/Y AND2X1_LOC_727/A 0.01fF
C33507 OR2X1_LOC_691/a_36_216# OR2X1_LOC_532/B 0.00fF
C33508 AND2X1_LOC_95/Y OR2X1_LOC_553/A 0.07fF
C33509 OR2X1_LOC_70/Y OR2X1_LOC_59/Y 0.12fF
C33510 VDD OR2X1_LOC_278/A 0.19fF
C33511 AND2X1_LOC_227/Y OR2X1_LOC_595/A 0.17fF
C33512 AND2X1_LOC_542/a_8_24# OR2X1_LOC_417/A 0.06fF
C33513 OR2X1_LOC_409/B AND2X1_LOC_828/a_8_24# 0.10fF
C33514 OR2X1_LOC_856/B OR2X1_LOC_269/B 0.07fF
C33515 OR2X1_LOC_756/B OR2X1_LOC_592/A 0.02fF
C33516 AND2X1_LOC_351/Y OR2X1_LOC_51/Y 0.23fF
C33517 OR2X1_LOC_804/A OR2X1_LOC_831/B 0.02fF
C33518 OR2X1_LOC_6/B INPUT_1 0.44fF
C33519 OR2X1_LOC_857/a_8_216# OR2X1_LOC_35/Y 0.01fF
C33520 AND2X1_LOC_716/Y OR2X1_LOC_7/A 0.07fF
C33521 OR2X1_LOC_448/Y OR2X1_LOC_453/a_8_216# 0.07fF
C33522 D_INPUT_4 OR2X1_LOC_21/a_8_216# 0.02fF
C33523 OR2X1_LOC_695/a_8_216# OR2X1_LOC_52/B 0.03fF
C33524 OR2X1_LOC_637/B AND2X1_LOC_3/Y 0.01fF
C33525 OR2X1_LOC_151/A AND2X1_LOC_47/Y 0.57fF
C33526 AND2X1_LOC_717/a_8_24# AND2X1_LOC_374/Y 0.10fF
C33527 OR2X1_LOC_154/A OR2X1_LOC_375/A 0.42fF
C33528 AND2X1_LOC_546/a_8_24# OR2X1_LOC_26/Y 0.01fF
C33529 OR2X1_LOC_74/A OR2X1_LOC_746/a_36_216# 0.03fF
C33530 OR2X1_LOC_643/A OR2X1_LOC_231/a_8_216# 0.03fF
C33531 OR2X1_LOC_298/Y OR2X1_LOC_6/A 0.01fF
C33532 AND2X1_LOC_576/Y AND2X1_LOC_807/Y 0.10fF
C33533 AND2X1_LOC_512/Y AND2X1_LOC_729/B 0.01fF
C33534 OR2X1_LOC_416/Y AND2X1_LOC_219/Y 0.04fF
C33535 AND2X1_LOC_654/Y OR2X1_LOC_7/A 0.08fF
C33536 AND2X1_LOC_645/A OR2X1_LOC_48/B 0.01fF
C33537 OR2X1_LOC_744/A OR2X1_LOC_19/B 0.05fF
C33538 AND2X1_LOC_385/a_8_24# OR2X1_LOC_537/A 0.02fF
C33539 AND2X1_LOC_95/Y OR2X1_LOC_219/B 0.17fF
C33540 OR2X1_LOC_216/A OR2X1_LOC_475/Y 0.00fF
C33541 AND2X1_LOC_862/A AND2X1_LOC_806/A 0.01fF
C33542 AND2X1_LOC_11/Y AND2X1_LOC_3/Y 0.29fF
C33543 AND2X1_LOC_624/A AND2X1_LOC_806/A 0.03fF
C33544 OR2X1_LOC_484/Y AND2X1_LOC_727/A 0.01fF
C33545 OR2X1_LOC_521/Y AND2X1_LOC_276/Y 0.04fF
C33546 OR2X1_LOC_494/Y OR2X1_LOC_71/Y 0.02fF
C33547 OR2X1_LOC_267/A OR2X1_LOC_375/A 0.03fF
C33548 OR2X1_LOC_649/B OR2X1_LOC_130/A 0.05fF
C33549 OR2X1_LOC_569/B OR2X1_LOC_569/A 0.43fF
C33550 OR2X1_LOC_814/A OR2X1_LOC_363/A 0.02fF
C33551 OR2X1_LOC_809/B D_INPUT_0 0.12fF
C33552 OR2X1_LOC_320/Y AND2X1_LOC_654/Y 0.06fF
C33553 AND2X1_LOC_228/Y AND2X1_LOC_654/a_8_24# 0.01fF
C33554 OR2X1_LOC_6/B OR2X1_LOC_751/a_8_216# 0.04fF
C33555 AND2X1_LOC_40/Y AND2X1_LOC_1/Y 0.00fF
C33556 OR2X1_LOC_402/Y AND2X1_LOC_3/Y 0.09fF
C33557 OR2X1_LOC_41/Y OR2X1_LOC_428/A 0.30fF
C33558 AND2X1_LOC_456/Y AND2X1_LOC_573/A 0.03fF
C33559 INPUT_0 OR2X1_LOC_243/B 0.29fF
C33560 AND2X1_LOC_302/a_8_24# OR2X1_LOC_52/B 0.04fF
C33561 OR2X1_LOC_3/Y OR2X1_LOC_619/Y 0.13fF
C33562 OR2X1_LOC_705/B AND2X1_LOC_44/Y 0.41fF
C33563 AND2X1_LOC_34/a_8_24# AND2X1_LOC_34/Y 0.00fF
C33564 OR2X1_LOC_490/Y AND2X1_LOC_573/A 0.57fF
C33565 OR2X1_LOC_427/A AND2X1_LOC_260/a_8_24# 0.03fF
C33566 OR2X1_LOC_74/A AND2X1_LOC_573/A 0.10fF
C33567 OR2X1_LOC_475/a_8_216# OR2X1_LOC_121/B 0.00fF
C33568 OR2X1_LOC_485/A OR2X1_LOC_39/A 0.37fF
C33569 OR2X1_LOC_673/Y OR2X1_LOC_403/B 0.00fF
C33570 OR2X1_LOC_175/Y OR2X1_LOC_567/a_8_216# 0.05fF
C33571 OR2X1_LOC_306/a_36_216# OR2X1_LOC_743/A 0.02fF
C33572 AND2X1_LOC_303/A AND2X1_LOC_211/B 0.14fF
C33573 OR2X1_LOC_663/A OR2X1_LOC_814/A 0.03fF
C33574 AND2X1_LOC_76/Y AND2X1_LOC_663/B 0.00fF
C33575 OR2X1_LOC_580/a_8_216# OR2X1_LOC_580/B 0.06fF
C33576 OR2X1_LOC_714/a_8_216# OR2X1_LOC_714/A 0.39fF
C33577 AND2X1_LOC_44/Y AND2X1_LOC_609/a_8_24# 0.04fF
C33578 AND2X1_LOC_80/a_8_24# OR2X1_LOC_647/A 0.01fF
C33579 AND2X1_LOC_495/a_36_24# OR2X1_LOC_203/Y 0.01fF
C33580 AND2X1_LOC_256/a_36_24# OR2X1_LOC_598/A 0.00fF
C33581 GATE_366 OR2X1_LOC_7/A 0.01fF
C33582 OR2X1_LOC_158/A AND2X1_LOC_205/a_8_24# 0.02fF
C33583 AND2X1_LOC_569/a_8_24# AND2X1_LOC_474/Y 0.03fF
C33584 OR2X1_LOC_223/A OR2X1_LOC_785/a_8_216# 0.01fF
C33585 OR2X1_LOC_3/Y OR2X1_LOC_88/A 0.09fF
C33586 OR2X1_LOC_96/Y AND2X1_LOC_721/A 0.00fF
C33587 AND2X1_LOC_40/Y OR2X1_LOC_471/Y 0.03fF
C33588 OR2X1_LOC_778/A OR2X1_LOC_375/A 0.02fF
C33589 OR2X1_LOC_158/A OR2X1_LOC_163/A 0.04fF
C33590 OR2X1_LOC_846/a_36_216# OR2X1_LOC_846/B 0.01fF
C33591 OR2X1_LOC_497/Y AND2X1_LOC_717/B 0.07fF
C33592 OR2X1_LOC_151/A OR2X1_LOC_598/A 0.84fF
C33593 OR2X1_LOC_32/Y OR2X1_LOC_52/B 0.01fF
C33594 AND2X1_LOC_114/Y OR2X1_LOC_56/A 0.01fF
C33595 AND2X1_LOC_17/Y AND2X1_LOC_44/a_8_24# 0.01fF
C33596 OR2X1_LOC_852/B D_INPUT_0 0.02fF
C33597 AND2X1_LOC_572/Y OR2X1_LOC_64/Y 0.02fF
C33598 AND2X1_LOC_684/a_8_24# OR2X1_LOC_78/B 0.02fF
C33599 OR2X1_LOC_400/B OR2X1_LOC_557/A 0.01fF
C33600 OR2X1_LOC_742/B OR2X1_LOC_550/A 0.08fF
C33601 OR2X1_LOC_166/a_36_216# OR2X1_LOC_47/Y 0.01fF
C33602 AND2X1_LOC_3/Y OR2X1_LOC_217/a_8_216# 0.01fF
C33603 AND2X1_LOC_36/Y INPUT_6 0.03fF
C33604 AND2X1_LOC_775/a_8_24# OR2X1_LOC_70/Y 0.01fF
C33605 OR2X1_LOC_848/A OR2X1_LOC_846/B 0.04fF
C33606 OR2X1_LOC_161/B OR2X1_LOC_789/A 0.03fF
C33607 OR2X1_LOC_312/Y OR2X1_LOC_7/A 0.03fF
C33608 AND2X1_LOC_712/B AND2X1_LOC_448/Y 0.41fF
C33609 OR2X1_LOC_70/Y OR2X1_LOC_433/a_8_216# 0.08fF
C33610 AND2X1_LOC_477/A OR2X1_LOC_48/B 0.07fF
C33611 OR2X1_LOC_184/Y OR2X1_LOC_59/Y 0.01fF
C33612 OR2X1_LOC_481/A OR2X1_LOC_236/a_36_216# 0.00fF
C33613 AND2X1_LOC_6/a_8_24# OR2X1_LOC_78/B 0.01fF
C33614 AND2X1_LOC_47/Y OR2X1_LOC_788/a_8_216# 0.01fF
C33615 OR2X1_LOC_36/Y AND2X1_LOC_523/Y 0.05fF
C33616 OR2X1_LOC_437/Y OR2X1_LOC_59/Y 0.90fF
C33617 AND2X1_LOC_122/a_36_24# OR2X1_LOC_124/Y 0.00fF
C33618 OR2X1_LOC_426/A OR2X1_LOC_426/a_8_216# 0.04fF
C33619 OR2X1_LOC_70/Y AND2X1_LOC_446/a_36_24# 0.00fF
C33620 OR2X1_LOC_160/A D_INPUT_0 0.22fF
C33621 OR2X1_LOC_438/Y OR2X1_LOC_47/Y 0.43fF
C33622 AND2X1_LOC_663/B OR2X1_LOC_52/B -0.00fF
C33623 AND2X1_LOC_51/A AND2X1_LOC_51/Y 0.43fF
C33624 AND2X1_LOC_662/B OR2X1_LOC_31/Y 0.03fF
C33625 AND2X1_LOC_139/B INPUT_1 0.07fF
C33626 OR2X1_LOC_811/A AND2X1_LOC_665/a_36_24# 0.01fF
C33627 AND2X1_LOC_191/Y OR2X1_LOC_70/Y 0.03fF
C33628 AND2X1_LOC_479/Y OR2X1_LOC_427/A 0.01fF
C33629 OR2X1_LOC_377/A AND2X1_LOC_821/a_8_24# 0.01fF
C33630 AND2X1_LOC_59/Y OR2X1_LOC_532/B 1.62fF
C33631 AND2X1_LOC_62/a_8_24# D_INPUT_3 0.01fF
C33632 AND2X1_LOC_307/a_8_24# OR2X1_LOC_7/A 0.06fF
C33633 D_GATE_741 OR2X1_LOC_192/B 0.00fF
C33634 OR2X1_LOC_364/A OR2X1_LOC_814/A 0.10fF
C33635 OR2X1_LOC_576/A OR2X1_LOC_571/Y 0.15fF
C33636 AND2X1_LOC_845/Y OR2X1_LOC_67/a_8_216# 0.05fF
C33637 OR2X1_LOC_185/Y OR2X1_LOC_814/A 2.28fF
C33638 AND2X1_LOC_711/Y OR2X1_LOC_70/Y 0.03fF
C33639 AND2X1_LOC_662/a_8_24# OR2X1_LOC_74/A 0.06fF
C33640 OR2X1_LOC_70/A OR2X1_LOC_59/Y 0.01fF
C33641 OR2X1_LOC_383/Y OR2X1_LOC_269/B 0.01fF
C33642 OR2X1_LOC_426/A AND2X1_LOC_451/a_8_24# 0.01fF
C33643 AND2X1_LOC_42/B OR2X1_LOC_97/a_36_216# 0.00fF
C33644 AND2X1_LOC_850/A OR2X1_LOC_419/Y 0.01fF
C33645 AND2X1_LOC_849/A OR2X1_LOC_89/A 0.01fF
C33646 OR2X1_LOC_56/A OR2X1_LOC_172/a_8_216# -0.03fF
C33647 AND2X1_LOC_648/B OR2X1_LOC_432/Y 0.01fF
C33648 OR2X1_LOC_858/A AND2X1_LOC_31/Y 0.02fF
C33649 OR2X1_LOC_550/a_8_216# OR2X1_LOC_550/B 0.08fF
C33650 AND2X1_LOC_860/A OR2X1_LOC_384/Y 0.09fF
C33651 OR2X1_LOC_47/Y AND2X1_LOC_621/Y 0.03fF
C33652 OR2X1_LOC_115/a_36_216# OR2X1_LOC_786/Y 0.00fF
C33653 AND2X1_LOC_576/Y OR2X1_LOC_95/Y 0.13fF
C33654 OR2X1_LOC_755/A AND2X1_LOC_663/B 0.00fF
C33655 OR2X1_LOC_78/B OR2X1_LOC_560/A 0.05fF
C33656 OR2X1_LOC_840/a_8_216# OR2X1_LOC_723/B 0.03fF
C33657 AND2X1_LOC_92/Y OR2X1_LOC_724/A 0.08fF
C33658 OR2X1_LOC_158/A AND2X1_LOC_449/a_8_24# 0.01fF
C33659 AND2X1_LOC_568/B AND2X1_LOC_212/a_8_24# 0.02fF
C33660 AND2X1_LOC_55/a_8_24# OR2X1_LOC_62/A 0.03fF
C33661 OR2X1_LOC_40/Y OR2X1_LOC_13/B 0.25fF
C33662 OR2X1_LOC_855/A AND2X1_LOC_763/B 0.05fF
C33663 AND2X1_LOC_64/Y OR2X1_LOC_338/A 0.07fF
C33664 OR2X1_LOC_833/B AND2X1_LOC_271/a_36_24# 0.00fF
C33665 OR2X1_LOC_191/B AND2X1_LOC_47/Y 0.02fF
C33666 OR2X1_LOC_794/A OR2X1_LOC_374/Y 0.10fF
C33667 AND2X1_LOC_6/a_8_24# OR2X1_LOC_375/A 0.01fF
C33668 AND2X1_LOC_524/a_8_24# AND2X1_LOC_36/Y 0.05fF
C33669 OR2X1_LOC_52/a_8_216# OR2X1_LOC_7/Y 0.01fF
C33670 INPUT_4 AND2X1_LOC_451/a_8_24# 0.01fF
C33671 AND2X1_LOC_40/Y OR2X1_LOC_750/Y 0.01fF
C33672 AND2X1_LOC_535/a_8_24# OR2X1_LOC_13/B 0.02fF
C33673 OR2X1_LOC_325/B OR2X1_LOC_532/Y 0.06fF
C33674 AND2X1_LOC_711/Y OR2X1_LOC_504/Y 0.03fF
C33675 OR2X1_LOC_180/a_8_216# OR2X1_LOC_180/B 0.02fF
C33676 OR2X1_LOC_721/Y OR2X1_LOC_560/A 0.05fF
C33677 OR2X1_LOC_280/Y OR2X1_LOC_238/a_8_216# 0.04fF
C33678 OR2X1_LOC_476/B OR2X1_LOC_750/A 0.00fF
C33679 OR2X1_LOC_45/B AND2X1_LOC_539/Y 0.03fF
C33680 OR2X1_LOC_760/Y OR2X1_LOC_585/A 0.01fF
C33681 AND2X1_LOC_573/A AND2X1_LOC_647/Y 0.02fF
C33682 AND2X1_LOC_722/A OR2X1_LOC_533/a_8_216# 0.06fF
C33683 OR2X1_LOC_485/A OR2X1_LOC_760/a_8_216# 0.01fF
C33684 OR2X1_LOC_186/Y AND2X1_LOC_64/Y 0.34fF
C33685 AND2X1_LOC_170/B AND2X1_LOC_212/B 0.50fF
C33686 OR2X1_LOC_273/Y OR2X1_LOC_31/Y 0.31fF
C33687 AND2X1_LOC_287/B AND2X1_LOC_244/A 0.08fF
C33688 OR2X1_LOC_151/A OR2X1_LOC_186/a_8_216# 0.02fF
C33689 OR2X1_LOC_497/a_36_216# OR2X1_LOC_419/Y 0.00fF
C33690 OR2X1_LOC_537/A OR2X1_LOC_750/Y 0.01fF
C33691 OR2X1_LOC_185/A OR2X1_LOC_344/a_8_216# 0.01fF
C33692 OR2X1_LOC_743/A AND2X1_LOC_687/a_8_24# 0.08fF
C33693 OR2X1_LOC_134/a_8_216# AND2X1_LOC_541/Y 0.01fF
C33694 D_INPUT_7 OR2X1_LOC_2/a_8_216# 0.01fF
C33695 OR2X1_LOC_97/A AND2X1_LOC_433/a_8_24# 0.01fF
C33696 OR2X1_LOC_375/A OR2X1_LOC_560/A 0.10fF
C33697 OR2X1_LOC_291/A OR2X1_LOC_234/a_8_216# 0.39fF
C33698 AND2X1_LOC_66/a_8_24# AND2X1_LOC_845/Y 0.02fF
C33699 OR2X1_LOC_375/A OR2X1_LOC_198/A 0.01fF
C33700 OR2X1_LOC_548/B OR2X1_LOC_548/a_8_216# 0.07fF
C33701 AND2X1_LOC_625/a_36_24# OR2X1_LOC_115/B 0.00fF
C33702 AND2X1_LOC_41/A OR2X1_LOC_469/B 0.18fF
C33703 AND2X1_LOC_47/Y INPUT_1 0.55fF
C33704 AND2X1_LOC_843/Y OR2X1_LOC_13/B 0.02fF
C33705 AND2X1_LOC_712/a_8_24# OR2X1_LOC_158/A 0.01fF
C33706 AND2X1_LOC_64/Y AND2X1_LOC_310/a_8_24# 0.01fF
C33707 AND2X1_LOC_552/A OR2X1_LOC_373/Y 0.03fF
C33708 OR2X1_LOC_78/A OR2X1_LOC_502/Y 0.02fF
C33709 AND2X1_LOC_701/a_8_24# AND2X1_LOC_31/Y 0.01fF
C33710 AND2X1_LOC_729/B OR2X1_LOC_41/a_36_216# 0.00fF
C33711 OR2X1_LOC_323/A OR2X1_LOC_744/A 0.03fF
C33712 OR2X1_LOC_307/A OR2X1_LOC_161/B 0.25fF
C33713 AND2X1_LOC_22/Y OR2X1_LOC_160/B 0.80fF
C33714 OR2X1_LOC_19/B OR2X1_LOC_396/a_36_216# 0.02fF
C33715 OR2X1_LOC_853/a_8_216# OR2X1_LOC_66/A 0.02fF
C33716 OR2X1_LOC_447/a_8_216# OR2X1_LOC_777/B 0.14fF
C33717 OR2X1_LOC_617/Y AND2X1_LOC_805/a_36_24# 0.01fF
C33718 OR2X1_LOC_278/A OR2X1_LOC_67/Y 0.79fF
C33719 OR2X1_LOC_508/A AND2X1_LOC_239/a_36_24# 0.00fF
C33720 OR2X1_LOC_31/Y OR2X1_LOC_75/Y 0.00fF
C33721 OR2X1_LOC_56/A OR2X1_LOC_312/a_8_216# 0.02fF
C33722 AND2X1_LOC_462/B AND2X1_LOC_462/a_8_24# 0.01fF
C33723 AND2X1_LOC_425/a_8_24# AND2X1_LOC_430/B 0.01fF
C33724 AND2X1_LOC_756/a_8_24# GATE_579 0.01fF
C33725 OR2X1_LOC_595/Y OR2X1_LOC_416/Y 0.02fF
C33726 OR2X1_LOC_154/A OR2X1_LOC_515/Y 0.36fF
C33727 VDD OR2X1_LOC_135/Y 1.34fF
C33728 VDD OR2X1_LOC_663/a_8_216# 0.00fF
C33729 OR2X1_LOC_744/A OR2X1_LOC_744/a_8_216# 0.20fF
C33730 AND2X1_LOC_592/Y AND2X1_LOC_593/a_8_24# 0.01fF
C33731 OR2X1_LOC_203/a_8_216# AND2X1_LOC_36/Y 0.01fF
C33732 OR2X1_LOC_70/Y OR2X1_LOC_534/a_36_216# 0.00fF
C33733 OR2X1_LOC_539/Y OR2X1_LOC_175/a_36_216# 0.00fF
C33734 OR2X1_LOC_491/a_8_216# OR2X1_LOC_108/Y 0.07fF
C33735 OR2X1_LOC_532/B OR2X1_LOC_733/Y 0.01fF
C33736 OR2X1_LOC_87/A OR2X1_LOC_712/B 0.02fF
C33737 OR2X1_LOC_45/B AND2X1_LOC_471/Y 0.01fF
C33738 AND2X1_LOC_776/Y AND2X1_LOC_486/Y 0.72fF
C33739 AND2X1_LOC_788/a_8_24# OR2X1_LOC_51/Y 0.00fF
C33740 OR2X1_LOC_600/A AND2X1_LOC_477/Y 0.03fF
C33741 INPUT_1 OR2X1_LOC_598/A 0.10fF
C33742 AND2X1_LOC_810/A OR2X1_LOC_91/A 0.05fF
C33743 OR2X1_LOC_124/A AND2X1_LOC_65/A 0.07fF
C33744 OR2X1_LOC_696/A AND2X1_LOC_554/Y 0.07fF
C33745 OR2X1_LOC_7/A OR2X1_LOC_13/B 0.84fF
C33746 OR2X1_LOC_51/Y AND2X1_LOC_476/Y 0.07fF
C33747 AND2X1_LOC_719/Y AND2X1_LOC_658/A 0.04fF
C33748 AND2X1_LOC_70/Y OR2X1_LOC_648/B 0.03fF
C33749 AND2X1_LOC_357/B OR2X1_LOC_426/B 0.04fF
C33750 OR2X1_LOC_502/A AND2X1_LOC_44/Y 7.63fF
C33751 OR2X1_LOC_320/Y OR2X1_LOC_13/B 0.58fF
C33752 AND2X1_LOC_787/A AND2X1_LOC_717/Y 0.12fF
C33753 OR2X1_LOC_78/A AND2X1_LOC_265/a_8_24# 0.08fF
C33754 AND2X1_LOC_566/B INPUT_0 0.03fF
C33755 OR2X1_LOC_308/A OR2X1_LOC_161/A 0.01fF
C33756 OR2X1_LOC_778/Y OR2X1_LOC_308/Y 0.10fF
C33757 OR2X1_LOC_510/Y OR2X1_LOC_115/B 0.42fF
C33758 OR2X1_LOC_792/Y OR2X1_LOC_758/a_8_216# 0.02fF
C33759 AND2X1_LOC_64/Y AND2X1_LOC_81/B 0.09fF
C33760 AND2X1_LOC_858/B AND2X1_LOC_860/A 0.01fF
C33761 OR2X1_LOC_405/A OR2X1_LOC_97/A 0.03fF
C33762 AND2X1_LOC_703/Y OR2X1_LOC_48/B 0.23fF
C33763 VDD OR2X1_LOC_78/A 1.75fF
C33764 OR2X1_LOC_316/a_8_216# OR2X1_LOC_44/Y 0.04fF
C33765 OR2X1_LOC_329/B OR2X1_LOC_600/A 0.07fF
C33766 OR2X1_LOC_91/A AND2X1_LOC_860/A 0.13fF
C33767 VDD AND2X1_LOC_443/Y 0.21fF
C33768 AND2X1_LOC_540/a_8_24# OR2X1_LOC_158/A 0.02fF
C33769 AND2X1_LOC_808/a_8_24# AND2X1_LOC_727/B 0.19fF
C33770 OR2X1_LOC_614/a_8_216# AND2X1_LOC_31/Y 0.01fF
C33771 AND2X1_LOC_392/A AND2X1_LOC_365/a_8_24# 0.04fF
C33772 OR2X1_LOC_851/B AND2X1_LOC_40/Y 0.08fF
C33773 OR2X1_LOC_114/a_8_216# OR2X1_LOC_114/B 0.05fF
C33774 OR2X1_LOC_458/B OR2X1_LOC_723/a_36_216# 0.00fF
C33775 OR2X1_LOC_244/Y OR2X1_LOC_363/A 0.00fF
C33776 AND2X1_LOC_136/a_8_24# AND2X1_LOC_36/Y 0.01fF
C33777 OR2X1_LOC_22/Y OR2X1_LOC_385/a_8_216# 0.10fF
C33778 OR2X1_LOC_220/A OR2X1_LOC_565/A 0.12fF
C33779 AND2X1_LOC_87/a_8_24# AND2X1_LOC_202/Y 0.19fF
C33780 OR2X1_LOC_401/A OR2X1_LOC_771/B 0.03fF
C33781 OR2X1_LOC_160/B OR2X1_LOC_706/A 0.23fF
C33782 AND2X1_LOC_330/a_36_24# OR2X1_LOC_59/Y 0.00fF
C33783 AND2X1_LOC_454/Y OR2X1_LOC_428/A 0.39fF
C33784 AND2X1_LOC_92/Y OR2X1_LOC_520/a_36_216# 0.00fF
C33785 OR2X1_LOC_458/B VDD 0.29fF
C33786 OR2X1_LOC_325/A OR2X1_LOC_325/B 0.56fF
C33787 OR2X1_LOC_696/A OR2X1_LOC_280/Y 0.50fF
C33788 OR2X1_LOC_865/A OR2X1_LOC_865/a_8_216# 0.14fF
C33789 AND2X1_LOC_22/Y OR2X1_LOC_266/a_8_216# 0.03fF
C33790 OR2X1_LOC_810/A OR2X1_LOC_115/B 0.01fF
C33791 OR2X1_LOC_791/B OR2X1_LOC_580/B 0.01fF
C33792 AND2X1_LOC_605/Y AND2X1_LOC_454/a_8_24# 0.01fF
C33793 AND2X1_LOC_212/A AND2X1_LOC_661/a_8_24# 0.00fF
C33794 OR2X1_LOC_708/Y OR2X1_LOC_66/A 0.01fF
C33795 OR2X1_LOC_161/A OR2X1_LOC_160/Y 0.56fF
C33796 OR2X1_LOC_139/A OR2X1_LOC_87/A 0.07fF
C33797 OR2X1_LOC_62/B OR2X1_LOC_777/B 3.41fF
C33798 OR2X1_LOC_6/A OR2X1_LOC_310/a_8_216# 0.02fF
C33799 OR2X1_LOC_190/A OR2X1_LOC_190/B 0.03fF
C33800 OR2X1_LOC_91/Y AND2X1_LOC_786/Y 0.07fF
C33801 AND2X1_LOC_353/a_8_24# AND2X1_LOC_654/Y 0.04fF
C33802 OR2X1_LOC_151/A OR2X1_LOC_506/A 0.07fF
C33803 VDD OR2X1_LOC_448/B 0.21fF
C33804 OR2X1_LOC_427/A AND2X1_LOC_243/Y 0.07fF
C33805 OR2X1_LOC_599/A OR2X1_LOC_428/A 0.03fF
C33806 AND2X1_LOC_766/a_8_24# AND2X1_LOC_3/Y 0.02fF
C33807 AND2X1_LOC_754/a_8_24# AND2X1_LOC_43/B 0.01fF
C33808 AND2X1_LOC_392/A AND2X1_LOC_76/Y 0.03fF
C33809 AND2X1_LOC_70/Y AND2X1_LOC_331/a_8_24# 0.06fF
C33810 OR2X1_LOC_589/A AND2X1_LOC_435/a_36_24# 0.00fF
C33811 OR2X1_LOC_821/Y OR2X1_LOC_246/Y 0.30fF
C33812 AND2X1_LOC_854/a_8_24# OR2X1_LOC_428/A 0.06fF
C33813 AND2X1_LOC_22/Y OR2X1_LOC_219/B 0.03fF
C33814 OR2X1_LOC_269/B OR2X1_LOC_578/a_8_216# 0.04fF
C33815 OR2X1_LOC_591/A OR2X1_LOC_12/Y 0.01fF
C33816 OR2X1_LOC_93/a_8_216# OR2X1_LOC_428/A 0.02fF
C33817 OR2X1_LOC_154/A OR2X1_LOC_549/A 0.10fF
C33818 VDD AND2X1_LOC_520/Y 0.18fF
C33819 OR2X1_LOC_680/A AND2X1_LOC_476/Y 0.07fF
C33820 AND2X1_LOC_340/a_8_24# AND2X1_LOC_573/A 0.01fF
C33821 OR2X1_LOC_47/Y OR2X1_LOC_71/A 0.03fF
C33822 OR2X1_LOC_325/Y OR2X1_LOC_620/Y 0.02fF
C33823 OR2X1_LOC_133/a_8_216# OR2X1_LOC_43/A 0.04fF
C33824 INPUT_0 OR2X1_LOC_637/B 0.01fF
C33825 AND2X1_LOC_512/Y AND2X1_LOC_513/a_8_24# 0.03fF
C33826 OR2X1_LOC_371/a_8_216# AND2X1_LOC_786/Y 0.04fF
C33827 AND2X1_LOC_41/A OR2X1_LOC_274/Y 0.01fF
C33828 OR2X1_LOC_49/A OR2X1_LOC_646/A 0.02fF
C33829 OR2X1_LOC_185/A OR2X1_LOC_66/A 0.64fF
C33830 AND2X1_LOC_132/a_8_24# AND2X1_LOC_18/Y 0.01fF
C33831 OR2X1_LOC_496/a_8_216# OR2X1_LOC_18/Y 0.01fF
C33832 AND2X1_LOC_22/Y OR2X1_LOC_794/a_8_216# 0.01fF
C33833 AND2X1_LOC_702/Y OR2X1_LOC_589/A 0.03fF
C33834 VDD AND2X1_LOC_175/B 0.23fF
C33835 OR2X1_LOC_854/a_8_216# OR2X1_LOC_538/A -0.00fF
C33836 AND2X1_LOC_59/Y OR2X1_LOC_440/B 0.01fF
C33837 AND2X1_LOC_392/A OR2X1_LOC_67/A 0.03fF
C33838 OR2X1_LOC_600/A AND2X1_LOC_113/Y 0.00fF
C33839 AND2X1_LOC_702/a_8_24# OR2X1_LOC_426/B 0.04fF
C33840 OR2X1_LOC_249/Y OR2X1_LOC_66/A 0.11fF
C33841 OR2X1_LOC_696/A OR2X1_LOC_22/Y 0.59fF
C33842 OR2X1_LOC_377/A OR2X1_LOC_461/a_8_216# 0.06fF
C33843 AND2X1_LOC_201/a_8_24# AND2X1_LOC_201/Y 0.01fF
C33844 VDD AND2X1_LOC_848/Y 0.15fF
C33845 OR2X1_LOC_70/A OR2X1_LOC_11/a_36_216# -0.00fF
C33846 OR2X1_LOC_58/Y OR2X1_LOC_85/A 0.01fF
C33847 D_INPUT_0 OR2X1_LOC_130/Y 0.01fF
C33848 OR2X1_LOC_329/Y OR2X1_LOC_43/A 0.01fF
C33849 OR2X1_LOC_256/Y AND2X1_LOC_348/A 0.01fF
C33850 OR2X1_LOC_17/Y INPUT_7 0.35fF
C33851 OR2X1_LOC_461/a_8_216# AND2X1_LOC_824/B 0.04fF
C33852 OR2X1_LOC_329/B OR2X1_LOC_619/Y 0.07fF
C33853 OR2X1_LOC_687/Y OR2X1_LOC_676/Y 0.07fF
C33854 AND2X1_LOC_114/a_8_24# OR2X1_LOC_56/A 0.01fF
C33855 OR2X1_LOC_405/A OR2X1_LOC_541/A 0.00fF
C33856 OR2X1_LOC_673/B OR2X1_LOC_624/B 0.02fF
C33857 OR2X1_LOC_814/A OR2X1_LOC_366/A 0.01fF
C33858 AND2X1_LOC_787/A OR2X1_LOC_64/Y 0.03fF
C33859 AND2X1_LOC_363/Y AND2X1_LOC_367/a_8_24# 0.01fF
C33860 OR2X1_LOC_625/a_8_216# OR2X1_LOC_517/A 0.01fF
C33861 AND2X1_LOC_72/B OR2X1_LOC_501/a_36_216# 0.00fF
C33862 OR2X1_LOC_527/Y AND2X1_LOC_786/Y 0.04fF
C33863 AND2X1_LOC_388/a_8_24# OR2X1_LOC_744/A 0.01fF
C33864 OR2X1_LOC_354/A OR2X1_LOC_620/Y 0.01fF
C33865 VDD OR2X1_LOC_283/Y 0.04fF
C33866 OR2X1_LOC_455/A OR2X1_LOC_486/Y 0.11fF
C33867 AND2X1_LOC_679/a_8_24# OR2X1_LOC_446/B 0.05fF
C33868 AND2X1_LOC_67/a_8_24# OR2X1_LOC_506/A 0.01fF
C33869 OR2X1_LOC_185/Y OR2X1_LOC_244/Y 0.07fF
C33870 AND2X1_LOC_715/Y OR2X1_LOC_22/Y 0.07fF
C33871 OR2X1_LOC_377/A OR2X1_LOC_634/A 0.05fF
C33872 AND2X1_LOC_392/A OR2X1_LOC_52/B 0.07fF
C33873 AND2X1_LOC_395/a_8_24# OR2X1_LOC_78/B 0.01fF
C33874 OR2X1_LOC_158/A AND2X1_LOC_155/Y 0.17fF
C33875 OR2X1_LOC_669/Y AND2X1_LOC_860/A 0.93fF
C33876 OR2X1_LOC_534/a_8_216# OR2X1_LOC_534/Y 0.01fF
C33877 AND2X1_LOC_219/a_8_24# OR2X1_LOC_26/Y 0.02fF
C33878 AND2X1_LOC_191/B OR2X1_LOC_36/Y 0.00fF
C33879 AND2X1_LOC_736/Y OR2X1_LOC_427/A 0.03fF
C33880 AND2X1_LOC_334/Y OR2X1_LOC_26/Y 0.01fF
C33881 OR2X1_LOC_778/A OR2X1_LOC_549/A 0.00fF
C33882 OR2X1_LOC_45/B AND2X1_LOC_687/A 0.02fF
C33883 AND2X1_LOC_605/Y AND2X1_LOC_449/Y 0.01fF
C33884 OR2X1_LOC_538/a_8_216# OR2X1_LOC_377/A 0.02fF
C33885 OR2X1_LOC_154/A OR2X1_LOC_113/Y 0.00fF
C33886 AND2X1_LOC_51/Y OR2X1_LOC_160/Y 0.02fF
C33887 VDD OR2X1_LOC_155/A 0.67fF
C33888 OR2X1_LOC_634/A AND2X1_LOC_824/B 0.17fF
C33889 OR2X1_LOC_323/A OR2X1_LOC_31/Y 0.22fF
C33890 AND2X1_LOC_858/B AND2X1_LOC_287/Y 0.01fF
C33891 OR2X1_LOC_405/A OR2X1_LOC_475/B 0.09fF
C33892 AND2X1_LOC_48/A AND2X1_LOC_44/Y 8.45fF
C33893 OR2X1_LOC_441/Y AND2X1_LOC_624/A 17.05fF
C33894 OR2X1_LOC_777/B OR2X1_LOC_365/B 0.10fF
C33895 OR2X1_LOC_517/A AND2X1_LOC_139/B 0.04fF
C33896 OR2X1_LOC_474/Y OR2X1_LOC_805/A 0.01fF
C33897 OR2X1_LOC_160/A AND2X1_LOC_40/Y 7.90fF
C33898 OR2X1_LOC_114/B AND2X1_LOC_42/B 0.03fF
C33899 OR2X1_LOC_364/Y OR2X1_LOC_365/a_8_216# 0.39fF
C33900 OR2X1_LOC_865/a_8_216# OR2X1_LOC_391/A 0.03fF
C33901 AND2X1_LOC_658/B AND2X1_LOC_191/Y 0.03fF
C33902 AND2X1_LOC_510/a_8_24# OR2X1_LOC_44/Y 0.01fF
C33903 AND2X1_LOC_22/Y OR2X1_LOC_244/A 0.07fF
C33904 AND2X1_LOC_566/B OR2X1_LOC_64/Y 0.06fF
C33905 OR2X1_LOC_437/A AND2X1_LOC_563/Y 0.03fF
C33906 D_INPUT_3 OR2X1_LOC_415/Y 0.02fF
C33907 AND2X1_LOC_787/A OR2X1_LOC_417/A 0.06fF
C33908 AND2X1_LOC_190/a_36_24# AND2X1_LOC_717/B 0.00fF
C33909 AND2X1_LOC_658/B AND2X1_LOC_711/Y 0.03fF
C33910 AND2X1_LOC_752/a_36_24# OR2X1_LOC_375/A 0.00fF
C33911 VDD OR2X1_LOC_617/Y 0.22fF
C33912 OR2X1_LOC_643/A OR2X1_LOC_624/a_36_216# 0.00fF
C33913 AND2X1_LOC_191/Y AND2X1_LOC_629/a_36_24# 0.01fF
C33914 AND2X1_LOC_214/A OR2X1_LOC_585/A 0.10fF
C33915 OR2X1_LOC_625/Y AND2X1_LOC_621/Y 0.06fF
C33916 AND2X1_LOC_658/B OR2X1_LOC_70/Y 0.03fF
C33917 AND2X1_LOC_150/a_8_24# OR2X1_LOC_62/B 0.00fF
C33918 OR2X1_LOC_48/Y OR2X1_LOC_56/A 0.01fF
C33919 AND2X1_LOC_95/Y AND2X1_LOC_233/a_8_24# 0.01fF
C33920 OR2X1_LOC_189/Y OR2X1_LOC_524/Y 0.07fF
C33921 AND2X1_LOC_779/a_8_24# OR2X1_LOC_511/Y 0.23fF
C33922 OR2X1_LOC_54/a_8_216# OR2X1_LOC_9/a_8_216# 0.47fF
C33923 OR2X1_LOC_158/A AND2X1_LOC_633/Y 0.02fF
C33924 AND2X1_LOC_70/Y OR2X1_LOC_123/B 0.01fF
C33925 AND2X1_LOC_857/Y AND2X1_LOC_654/a_8_24# 0.01fF
C33926 OR2X1_LOC_485/A AND2X1_LOC_474/A 0.03fF
C33927 AND2X1_LOC_866/A OR2X1_LOC_428/A 0.16fF
C33928 AND2X1_LOC_330/a_36_24# OR2X1_LOC_70/Y 0.01fF
C33929 OR2X1_LOC_493/A OR2X1_LOC_130/A 0.51fF
C33930 VDD AND2X1_LOC_856/B 0.01fF
C33931 OR2X1_LOC_695/Y OR2X1_LOC_64/Y 0.01fF
C33932 AND2X1_LOC_47/Y AND2X1_LOC_279/a_8_24# 0.10fF
C33933 AND2X1_LOC_448/Y AND2X1_LOC_453/Y 0.18fF
C33934 AND2X1_LOC_339/Y AND2X1_LOC_476/A 0.04fF
C33935 AND2X1_LOC_347/Y AND2X1_LOC_259/Y 0.03fF
C33936 OR2X1_LOC_95/Y OR2X1_LOC_16/A 0.05fF
C33937 VDD AND2X1_LOC_464/Y 0.21fF
C33938 OR2X1_LOC_158/A D_INPUT_0 0.12fF
C33939 VDD AND2X1_LOC_863/A 0.38fF
C33940 OR2X1_LOC_696/A OR2X1_LOC_387/a_8_216# 0.01fF
C33941 OR2X1_LOC_574/A OR2X1_LOC_776/a_36_216# 0.12fF
C33942 AND2X1_LOC_64/Y OR2X1_LOC_66/Y 0.05fF
C33943 OR2X1_LOC_160/A OR2X1_LOC_87/Y 0.15fF
C33944 AND2X1_LOC_3/Y OR2X1_LOC_574/a_8_216# 0.01fF
C33945 OR2X1_LOC_502/A AND2X1_LOC_36/a_8_24# 0.01fF
C33946 AND2X1_LOC_40/Y AND2X1_LOC_86/B 0.03fF
C33947 OR2X1_LOC_385/Y OR2X1_LOC_586/a_36_216# 0.01fF
C33948 OR2X1_LOC_109/Y OR2X1_LOC_26/Y 0.08fF
C33949 AND2X1_LOC_658/B AND2X1_LOC_657/a_8_24# 0.04fF
C33950 OR2X1_LOC_468/Y AND2X1_LOC_43/B 0.03fF
C33951 OR2X1_LOC_566/A OR2X1_LOC_365/B 0.02fF
C33952 OR2X1_LOC_495/a_8_216# OR2X1_LOC_39/A 0.02fF
C33953 AND2X1_LOC_40/Y OR2X1_LOC_624/B 0.09fF
C33954 AND2X1_LOC_658/B OR2X1_LOC_504/Y 0.15fF
C33955 OR2X1_LOC_108/Y OR2X1_LOC_95/Y 0.07fF
C33956 OR2X1_LOC_463/a_8_216# OR2X1_LOC_463/B 0.03fF
C33957 OR2X1_LOC_653/Y OR2X1_LOC_33/B 0.01fF
C33958 OR2X1_LOC_355/B OR2X1_LOC_739/A 0.01fF
C33959 OR2X1_LOC_470/B OR2X1_LOC_478/a_8_216# 0.01fF
C33960 OR2X1_LOC_109/Y OR2X1_LOC_89/A 0.01fF
C33961 AND2X1_LOC_717/a_8_24# OR2X1_LOC_280/Y 0.04fF
C33962 OR2X1_LOC_330/Y AND2X1_LOC_51/Y 0.01fF
C33963 OR2X1_LOC_151/A AND2X1_LOC_420/a_8_24# 0.03fF
C33964 OR2X1_LOC_251/Y AND2X1_LOC_848/Y 0.03fF
C33965 AND2X1_LOC_36/Y OR2X1_LOC_704/a_8_216# 0.01fF
C33966 AND2X1_LOC_6/a_8_24# OR2X1_LOC_549/A 0.06fF
C33967 OR2X1_LOC_485/A AND2X1_LOC_593/Y 0.03fF
C33968 AND2X1_LOC_777/a_8_24# OR2X1_LOC_305/Y 0.11fF
C33969 OR2X1_LOC_151/A D_INPUT_1 0.07fF
C33970 AND2X1_LOC_512/Y OR2X1_LOC_46/A 0.06fF
C33971 AND2X1_LOC_548/a_8_24# AND2X1_LOC_621/Y 0.03fF
C33972 OR2X1_LOC_529/Y AND2X1_LOC_624/A 0.05fF
C33973 AND2X1_LOC_656/Y OR2X1_LOC_56/A 0.24fF
C33974 AND2X1_LOC_702/Y OR2X1_LOC_43/A 0.03fF
C33975 AND2X1_LOC_772/B AND2X1_LOC_227/Y 0.01fF
C33976 OR2X1_LOC_600/A GATE_662 0.02fF
C33977 AND2X1_LOC_12/Y AND2X1_LOC_42/B 0.03fF
C33978 INPUT_3 AND2X1_LOC_37/a_36_24# 0.00fF
C33979 AND2X1_LOC_22/Y OR2X1_LOC_197/a_8_216# 0.05fF
C33980 OR2X1_LOC_262/a_8_216# OR2X1_LOC_26/Y 0.01fF
C33981 OR2X1_LOC_244/B OR2X1_LOC_244/A 0.29fF
C33982 OR2X1_LOC_141/B OR2X1_LOC_657/a_8_216# 0.01fF
C33983 OR2X1_LOC_588/Y AND2X1_LOC_637/Y 0.14fF
C33984 OR2X1_LOC_251/Y OR2X1_LOC_283/Y 0.16fF
C33985 OR2X1_LOC_837/B OR2X1_LOC_416/Y 0.03fF
C33986 AND2X1_LOC_48/A OR2X1_LOC_61/a_8_216# 0.01fF
C33987 OR2X1_LOC_160/A OR2X1_LOC_475/Y 0.02fF
C33988 OR2X1_LOC_485/A OR2X1_LOC_85/A 0.70fF
C33989 OR2X1_LOC_616/Y OR2X1_LOC_617/Y 0.20fF
C33990 INPUT_4 OR2X1_LOC_17/Y 2.19fF
C33991 OR2X1_LOC_401/A OR2X1_LOC_402/Y 0.03fF
C33992 OR2X1_LOC_91/Y AND2X1_LOC_578/A 0.07fF
C33993 OR2X1_LOC_62/B OR2X1_LOC_575/A 0.42fF
C33994 OR2X1_LOC_814/a_8_216# OR2X1_LOC_814/A 0.07fF
C33995 AND2X1_LOC_810/a_8_24# AND2X1_LOC_436/Y 0.01fF
C33996 AND2X1_LOC_63/a_8_24# AND2X1_LOC_10/a_8_24# 0.23fF
C33997 AND2X1_LOC_391/a_8_24# OR2X1_LOC_417/A 0.01fF
C33998 AND2X1_LOC_533/a_8_24# OR2X1_LOC_121/B 0.01fF
C33999 OR2X1_LOC_532/B OR2X1_LOC_623/B 0.06fF
C34000 OR2X1_LOC_47/Y OR2X1_LOC_59/Y 0.34fF
C34001 OR2X1_LOC_485/A AND2X1_LOC_602/a_8_24# 0.02fF
C34002 OR2X1_LOC_419/a_8_216# AND2X1_LOC_447/Y 0.49fF
C34003 OR2X1_LOC_18/Y AND2X1_LOC_465/Y 0.03fF
C34004 AND2X1_LOC_425/Y AND2X1_LOC_426/a_8_24# 0.05fF
C34005 OR2X1_LOC_517/a_8_216# AND2X1_LOC_660/A 0.06fF
C34006 OR2X1_LOC_287/B AND2X1_LOC_490/a_8_24# 0.00fF
C34007 INPUT_5 OR2X1_LOC_409/B 0.03fF
C34008 OR2X1_LOC_3/Y AND2X1_LOC_454/A 0.46fF
C34009 OR2X1_LOC_549/A OR2X1_LOC_560/A 0.02fF
C34010 AND2X1_LOC_17/Y AND2X1_LOC_425/a_8_24# 0.04fF
C34011 OR2X1_LOC_847/A D_INPUT_0 0.03fF
C34012 AND2X1_LOC_81/B OR2X1_LOC_206/A 0.00fF
C34013 OR2X1_LOC_26/Y AND2X1_LOC_729/B 0.02fF
C34014 AND2X1_LOC_776/a_8_24# OR2X1_LOC_406/A 0.01fF
C34015 OR2X1_LOC_92/Y AND2X1_LOC_476/A 0.65fF
C34016 OR2X1_LOC_189/Y AND2X1_LOC_578/A 0.03fF
C34017 AND2X1_LOC_374/a_36_24# OR2X1_LOC_31/Y 0.00fF
C34018 AND2X1_LOC_284/a_36_24# OR2X1_LOC_13/B 0.00fF
C34019 AND2X1_LOC_42/B AND2X1_LOC_79/Y 0.03fF
C34020 OR2X1_LOC_419/Y AND2X1_LOC_469/B 0.01fF
C34021 OR2X1_LOC_468/Y AND2X1_LOC_698/a_8_24# 0.08fF
C34022 AND2X1_LOC_12/Y OR2X1_LOC_286/B 0.01fF
C34023 AND2X1_LOC_796/a_8_24# AND2X1_LOC_796/A 0.03fF
C34024 OR2X1_LOC_769/A OR2X1_LOC_598/A 0.00fF
C34025 AND2X1_LOC_7/B OR2X1_LOC_771/B 0.05fF
C34026 OR2X1_LOC_274/a_8_216# OR2X1_LOC_241/B 0.03fF
C34027 AND2X1_LOC_660/Y AND2X1_LOC_116/Y 0.01fF
C34028 OR2X1_LOC_78/A OR2X1_LOC_140/a_8_216# 0.03fF
C34029 OR2X1_LOC_520/B AND2X1_LOC_8/Y 0.01fF
C34030 AND2X1_LOC_92/Y OR2X1_LOC_358/A 0.07fF
C34031 AND2X1_LOC_91/B OR2X1_LOC_308/Y 0.16fF
C34032 OR2X1_LOC_759/A AND2X1_LOC_793/B 0.34fF
C34033 OR2X1_LOC_557/A AND2X1_LOC_51/Y 1.94fF
C34034 OR2X1_LOC_472/A OR2X1_LOC_19/B 0.03fF
C34035 OR2X1_LOC_238/a_8_216# OR2X1_LOC_39/A 0.02fF
C34036 AND2X1_LOC_733/Y OR2X1_LOC_419/Y 0.01fF
C34037 OR2X1_LOC_194/Y AND2X1_LOC_7/Y 0.03fF
C34038 AND2X1_LOC_390/B AND2X1_LOC_855/a_8_24# 0.04fF
C34039 OR2X1_LOC_32/Y OR2X1_LOC_22/Y 0.04fF
C34040 AND2X1_LOC_657/Y OR2X1_LOC_152/A 0.03fF
C34041 OR2X1_LOC_185/A OR2X1_LOC_84/A 0.02fF
C34042 AND2X1_LOC_7/B OR2X1_LOC_776/A 0.01fF
C34043 AND2X1_LOC_858/B AND2X1_LOC_562/Y 0.10fF
C34044 AND2X1_LOC_578/A OR2X1_LOC_417/Y 0.01fF
C34045 OR2X1_LOC_137/Y OR2X1_LOC_720/B 0.05fF
C34046 OR2X1_LOC_111/Y OR2X1_LOC_36/Y 0.03fF
C34047 AND2X1_LOC_367/A AND2X1_LOC_222/Y 0.03fF
C34048 AND2X1_LOC_851/B OR2X1_LOC_6/A 0.03fF
C34049 VDD OR2X1_LOC_536/a_8_216# 0.00fF
C34050 OR2X1_LOC_85/A OR2X1_LOC_10/a_8_216# 0.03fF
C34051 OR2X1_LOC_812/B OR2X1_LOC_493/Y 0.09fF
C34052 OR2X1_LOC_325/B OR2X1_LOC_544/B 0.23fF
C34053 OR2X1_LOC_472/a_8_216# OR2X1_LOC_472/B 0.01fF
C34054 AND2X1_LOC_775/a_8_24# OR2X1_LOC_47/Y 0.01fF
C34055 OR2X1_LOC_698/Y AND2X1_LOC_793/B 0.00fF
C34056 OR2X1_LOC_76/B OR2X1_LOC_318/B 0.10fF
C34057 AND2X1_LOC_102/a_36_24# AND2X1_LOC_47/Y 0.00fF
C34058 OR2X1_LOC_241/Y OR2X1_LOC_810/A 0.10fF
C34059 VDD D_GATE_366 0.10fF
C34060 OR2X1_LOC_147/B OR2X1_LOC_552/A 0.03fF
C34061 OR2X1_LOC_485/A OR2X1_LOC_226/Y 0.01fF
C34062 OR2X1_LOC_151/A OR2X1_LOC_180/B 0.43fF
C34063 OR2X1_LOC_22/Y AND2X1_LOC_663/B 0.01fF
C34064 OR2X1_LOC_468/A OR2X1_LOC_777/B 0.03fF
C34065 OR2X1_LOC_323/A AND2X1_LOC_464/A 0.02fF
C34066 OR2X1_LOC_161/B OR2X1_LOC_186/a_36_216# 0.00fF
C34067 AND2X1_LOC_645/a_8_24# AND2X1_LOC_645/A 0.10fF
C34068 AND2X1_LOC_242/B AND2X1_LOC_242/a_8_24# 0.01fF
C34069 OR2X1_LOC_54/Y OR2X1_LOC_46/A 1.17fF
C34070 OR2X1_LOC_310/Y OR2X1_LOC_437/A 0.00fF
C34071 OR2X1_LOC_275/A OR2X1_LOC_31/Y 0.25fF
C34072 AND2X1_LOC_64/Y OR2X1_LOC_833/Y 0.02fF
C34073 AND2X1_LOC_143/a_8_24# OR2X1_LOC_71/A 0.05fF
C34074 AND2X1_LOC_841/a_36_24# OR2X1_LOC_74/A -0.02fF
C34075 AND2X1_LOC_191/Y OR2X1_LOC_47/Y 7.73fF
C34076 AND2X1_LOC_573/A AND2X1_LOC_562/Y 0.01fF
C34077 AND2X1_LOC_131/a_8_24# OR2X1_LOC_130/Y 0.00fF
C34078 OR2X1_LOC_494/A OR2X1_LOC_12/Y 0.00fF
C34079 AND2X1_LOC_191/Y AND2X1_LOC_866/a_36_24# 0.00fF
C34080 OR2X1_LOC_744/A OR2X1_LOC_142/Y 0.07fF
C34081 OR2X1_LOC_62/B OR2X1_LOC_62/a_36_216# 0.03fF
C34082 AND2X1_LOC_753/B OR2X1_LOC_193/a_8_216# 0.03fF
C34083 OR2X1_LOC_696/A OR2X1_LOC_485/Y 0.03fF
C34084 AND2X1_LOC_711/Y OR2X1_LOC_47/Y 0.03fF
C34085 AND2X1_LOC_539/Y OR2X1_LOC_158/A 0.03fF
C34086 OR2X1_LOC_715/B OR2X1_LOC_115/B 0.13fF
C34087 OR2X1_LOC_207/B AND2X1_LOC_44/Y 0.14fF
C34088 AND2X1_LOC_743/a_36_24# OR2X1_LOC_161/B 0.00fF
C34089 OR2X1_LOC_691/A OR2X1_LOC_857/A 0.05fF
C34090 OR2X1_LOC_629/B OR2X1_LOC_140/B 0.00fF
C34091 OR2X1_LOC_70/Y OR2X1_LOC_47/Y 0.12fF
C34092 AND2X1_LOC_729/Y AND2X1_LOC_796/A 0.03fF
C34093 AND2X1_LOC_561/a_8_24# AND2X1_LOC_561/B 0.00fF
C34094 AND2X1_LOC_765/a_8_24# AND2X1_LOC_82/Y 0.05fF
C34095 AND2X1_LOC_5/a_36_24# INPUT_1 0.00fF
C34096 OR2X1_LOC_48/B OR2X1_LOC_589/a_8_216# -0.02fF
C34097 OR2X1_LOC_611/a_8_216# OR2X1_LOC_62/A 0.02fF
C34098 AND2X1_LOC_687/Y OR2X1_LOC_95/Y 0.01fF
C34099 OR2X1_LOC_617/Y AND2X1_LOC_624/B 0.78fF
C34100 OR2X1_LOC_519/a_8_216# OR2X1_LOC_437/A 0.03fF
C34101 OR2X1_LOC_561/a_8_216# OR2X1_LOC_561/B 0.04fF
C34102 AND2X1_LOC_92/Y OR2X1_LOC_168/Y 0.15fF
C34103 OR2X1_LOC_809/a_8_216# AND2X1_LOC_31/Y 0.06fF
C34104 AND2X1_LOC_738/B OR2X1_LOC_525/a_36_216# 0.00fF
C34105 AND2X1_LOC_723/a_36_24# OR2X1_LOC_437/A 0.01fF
C34106 AND2X1_LOC_514/Y OR2X1_LOC_47/Y 0.08fF
C34107 OR2X1_LOC_864/A AND2X1_LOC_31/Y 0.06fF
C34108 OR2X1_LOC_363/A OR2X1_LOC_363/a_8_216# 0.19fF
C34109 OR2X1_LOC_36/Y AND2X1_LOC_206/Y 0.01fF
C34110 AND2X1_LOC_40/Y OR2X1_LOC_212/B 0.45fF
C34111 OR2X1_LOC_516/Y AND2X1_LOC_508/A 0.05fF
C34112 OR2X1_LOC_56/A AND2X1_LOC_772/Y 0.02fF
C34113 OR2X1_LOC_40/Y OR2X1_LOC_428/A 0.69fF
C34114 OR2X1_LOC_316/Y OR2X1_LOC_300/a_8_216# 0.01fF
C34115 OR2X1_LOC_457/B OR2X1_LOC_367/B 0.34fF
C34116 OR2X1_LOC_70/Y AND2X1_LOC_405/a_36_24# 0.00fF
C34117 OR2X1_LOC_74/A AND2X1_LOC_222/Y 0.47fF
C34118 OR2X1_LOC_70/Y AND2X1_LOC_486/a_36_24# 0.01fF
C34119 OR2X1_LOC_138/a_8_216# OR2X1_LOC_809/B 0.40fF
C34120 OR2X1_LOC_858/A OR2X1_LOC_121/A 0.02fF
C34121 OR2X1_LOC_51/Y AND2X1_LOC_636/a_8_24# 0.01fF
C34122 INPUT_1 D_INPUT_1 0.44fF
C34123 OR2X1_LOC_856/B OR2X1_LOC_319/Y 0.83fF
C34124 OR2X1_LOC_114/Y OR2X1_LOC_140/Y 0.03fF
C34125 OR2X1_LOC_97/A AND2X1_LOC_19/Y 0.02fF
C34126 OR2X1_LOC_269/B OR2X1_LOC_366/Y 0.10fF
C34127 OR2X1_LOC_756/B OR2X1_LOC_338/A 0.70fF
C34128 OR2X1_LOC_155/a_8_216# OR2X1_LOC_156/A 0.01fF
C34129 OR2X1_LOC_786/A OR2X1_LOC_786/a_8_216# 0.01fF
C34130 OR2X1_LOC_51/Y OR2X1_LOC_603/Y 0.02fF
C34131 OR2X1_LOC_9/Y OR2X1_LOC_96/Y 0.02fF
C34132 OR2X1_LOC_516/Y OR2X1_LOC_18/Y 0.03fF
C34133 OR2X1_LOC_86/a_8_216# OR2X1_LOC_13/B 0.02fF
C34134 OR2X1_LOC_276/B OR2X1_LOC_473/A 0.10fF
C34135 OR2X1_LOC_151/A OR2X1_LOC_440/a_36_216# 0.00fF
C34136 OR2X1_LOC_158/A AND2X1_LOC_711/A 0.01fF
C34137 AND2X1_LOC_318/Y AND2X1_LOC_798/A 0.00fF
C34138 OR2X1_LOC_158/A AND2X1_LOC_326/B 0.03fF
C34139 OR2X1_LOC_637/A OR2X1_LOC_828/Y 0.00fF
C34140 OR2X1_LOC_188/Y OR2X1_LOC_190/B 0.10fF
C34141 AND2X1_LOC_721/Y OR2X1_LOC_164/Y 0.00fF
C34142 OR2X1_LOC_805/A OR2X1_LOC_776/A 0.07fF
C34143 AND2X1_LOC_31/a_8_24# AND2X1_LOC_31/Y 0.02fF
C34144 AND2X1_LOC_22/Y OR2X1_LOC_307/B 0.04fF
C34145 AND2X1_LOC_719/Y AND2X1_LOC_190/a_8_24# 0.29fF
C34146 AND2X1_LOC_216/Y VDD 0.21fF
C34147 OR2X1_LOC_375/A AND2X1_LOC_409/B 0.03fF
C34148 OR2X1_LOC_696/A OR2X1_LOC_39/A 1.36fF
C34149 OR2X1_LOC_186/Y OR2X1_LOC_756/B 0.00fF
C34150 OR2X1_LOC_375/A OR2X1_LOC_605/Y 0.00fF
C34151 OR2X1_LOC_375/A AND2X1_LOC_763/B 0.02fF
C34152 OR2X1_LOC_653/Y OR2X1_LOC_392/B 0.02fF
C34153 AND2X1_LOC_570/Y AND2X1_LOC_500/B 0.02fF
C34154 OR2X1_LOC_856/A AND2X1_LOC_41/A 0.05fF
C34155 OR2X1_LOC_604/A AND2X1_LOC_657/Y 0.03fF
C34156 AND2X1_LOC_11/Y AND2X1_LOC_7/B 0.03fF
C34157 AND2X1_LOC_191/B OR2X1_LOC_604/A 0.07fF
C34158 AND2X1_LOC_102/a_8_24# AND2X1_LOC_36/Y 0.03fF
C34159 OR2X1_LOC_405/A OR2X1_LOC_175/Y 0.07fF
C34160 OR2X1_LOC_161/A OR2X1_LOC_703/a_8_216# 0.02fF
C34161 AND2X1_LOC_501/Y AND2X1_LOC_735/a_8_24# 0.01fF
C34162 AND2X1_LOC_23/a_36_24# OR2X1_LOC_228/Y 0.01fF
C34163 AND2X1_LOC_502/a_8_24# AND2X1_LOC_242/B 0.03fF
C34164 OR2X1_LOC_6/B AND2X1_LOC_628/a_36_24# 0.01fF
C34165 AND2X1_LOC_593/a_8_24# AND2X1_LOC_718/a_8_24# 0.23fF
C34166 OR2X1_LOC_158/A AND2X1_LOC_276/a_8_24# 0.03fF
C34167 AND2X1_LOC_571/A AND2X1_LOC_560/B 0.01fF
C34168 OR2X1_LOC_405/A OR2X1_LOC_691/Y 0.06fF
C34169 OR2X1_LOC_448/Y OR2X1_LOC_779/A 0.10fF
C34170 OR2X1_LOC_427/A OR2X1_LOC_12/Y 0.21fF
C34171 AND2X1_LOC_570/Y AND2X1_LOC_577/a_8_24# 0.11fF
C34172 AND2X1_LOC_421/a_8_24# OR2X1_LOC_596/A 0.11fF
C34173 OR2X1_LOC_821/a_8_216# OR2X1_LOC_278/Y 0.01fF
C34174 AND2X1_LOC_56/B OR2X1_LOC_334/a_8_216# 0.01fF
C34175 AND2X1_LOC_574/Y AND2X1_LOC_576/Y 0.03fF
C34176 OR2X1_LOC_696/A AND2X1_LOC_211/B 0.07fF
C34177 OR2X1_LOC_136/Y AND2X1_LOC_303/A 0.08fF
C34178 OR2X1_LOC_673/B OR2X1_LOC_847/A 0.00fF
C34179 OR2X1_LOC_633/A AND2X1_LOC_278/a_8_24# 0.04fF
C34180 OR2X1_LOC_47/Y OR2X1_LOC_70/A 0.13fF
C34181 OR2X1_LOC_121/B OR2X1_LOC_777/B 0.03fF
C34182 OR2X1_LOC_848/A OR2X1_LOC_774/a_8_216# 0.02fF
C34183 OR2X1_LOC_179/Y OR2X1_LOC_108/Y 0.01fF
C34184 OR2X1_LOC_377/A OR2X1_LOC_633/A 7.06fF
C34185 OR2X1_LOC_862/B OR2X1_LOC_561/Y 0.01fF
C34186 VDD AND2X1_LOC_562/B 0.04fF
C34187 OR2X1_LOC_158/A AND2X1_LOC_375/a_8_24# 0.06fF
C34188 OR2X1_LOC_815/Y AND2X1_LOC_846/a_8_24# 0.23fF
C34189 AND2X1_LOC_426/a_36_24# OR2X1_LOC_161/B 0.00fF
C34190 OR2X1_LOC_39/A OR2X1_LOC_522/a_36_216# 0.01fF
C34191 AND2X1_LOC_20/a_8_24# OR2X1_LOC_78/B 0.01fF
C34192 OR2X1_LOC_707/A OR2X1_LOC_161/B 0.03fF
C34193 OR2X1_LOC_97/A OR2X1_LOC_653/A 0.00fF
C34194 AND2X1_LOC_64/Y OR2X1_LOC_574/A 8.03fF
C34195 AND2X1_LOC_95/Y OR2X1_LOC_151/A 3.86fF
C34196 AND2X1_LOC_552/A OR2X1_LOC_109/Y 0.01fF
C34197 OR2X1_LOC_160/B AND2X1_LOC_173/a_8_24# 0.01fF
C34198 OR2X1_LOC_160/A OR2X1_LOC_356/A 0.01fF
C34199 OR2X1_LOC_6/B AND2X1_LOC_62/a_8_24# 0.02fF
C34200 AND2X1_LOC_555/Y OR2X1_LOC_485/A 0.00fF
C34201 AND2X1_LOC_64/Y OR2X1_LOC_33/A 0.10fF
C34202 OR2X1_LOC_851/B AND2X1_LOC_43/B 0.09fF
C34203 AND2X1_LOC_95/Y AND2X1_LOC_322/a_8_24# 0.02fF
C34204 AND2X1_LOC_555/Y AND2X1_LOC_348/a_8_24# 0.01fF
C34205 AND2X1_LOC_810/Y OR2X1_LOC_437/A 0.02fF
C34206 OR2X1_LOC_51/Y AND2X1_LOC_851/A 0.01fF
C34207 OR2X1_LOC_121/Y OR2X1_LOC_185/Y 0.11fF
C34208 OR2X1_LOC_49/A OR2X1_LOC_753/A 0.06fF
C34209 INPUT_1 AND2X1_LOC_789/Y 0.22fF
C34210 OR2X1_LOC_548/A AND2X1_LOC_56/B 0.13fF
C34211 OR2X1_LOC_215/a_36_216# AND2X1_LOC_31/Y 0.00fF
C34212 AND2X1_LOC_56/B OR2X1_LOC_486/Y 0.56fF
C34213 OR2X1_LOC_348/Y OR2X1_LOC_362/B 0.01fF
C34214 OR2X1_LOC_318/B OR2X1_LOC_552/A 0.00fF
C34215 AND2X1_LOC_507/a_8_24# OR2X1_LOC_18/Y 0.02fF
C34216 AND2X1_LOC_571/A OR2X1_LOC_64/Y 0.25fF
C34217 OR2X1_LOC_659/Y OR2X1_LOC_849/A 0.01fF
C34218 OR2X1_LOC_7/A OR2X1_LOC_428/A 0.27fF
C34219 AND2X1_LOC_512/Y AND2X1_LOC_722/A 0.07fF
C34220 AND2X1_LOC_698/a_36_24# OR2X1_LOC_308/Y 0.00fF
C34221 AND2X1_LOC_3/Y AND2X1_LOC_44/Y 2.83fF
C34222 OR2X1_LOC_190/A OR2X1_LOC_185/A 0.03fF
C34223 OR2X1_LOC_591/Y OR2X1_LOC_36/Y 0.03fF
C34224 OR2X1_LOC_158/A AND2X1_LOC_668/a_36_24# 0.01fF
C34225 GATE_811 AND2X1_LOC_742/A 0.29fF
C34226 AND2X1_LOC_152/a_36_24# OR2X1_LOC_740/B 0.00fF
C34227 AND2X1_LOC_592/Y OR2X1_LOC_599/A 0.01fF
C34228 AND2X1_LOC_720/a_8_24# OR2X1_LOC_59/Y 0.00fF
C34229 OR2X1_LOC_421/A AND2X1_LOC_319/A 0.03fF
C34230 INPUT_5 OR2X1_LOC_425/a_8_216# 0.07fF
C34231 OR2X1_LOC_377/A AND2X1_LOC_110/a_8_24# 0.12fF
C34232 AND2X1_LOC_766/a_8_24# OR2X1_LOC_401/A 0.01fF
C34233 OR2X1_LOC_7/A OR2X1_LOC_595/A 0.07fF
C34234 OR2X1_LOC_625/Y OR2X1_LOC_59/Y 0.07fF
C34235 OR2X1_LOC_652/a_8_216# OR2X1_LOC_468/A 0.18fF
C34236 OR2X1_LOC_121/B OR2X1_LOC_831/B 0.01fF
C34237 AND2X1_LOC_65/a_8_24# OR2X1_LOC_61/Y -0.01fF
C34238 OR2X1_LOC_318/B OR2X1_LOC_578/B 0.03fF
C34239 OR2X1_LOC_566/A OR2X1_LOC_121/B 0.06fF
C34240 AND2X1_LOC_580/A OR2X1_LOC_600/A 0.17fF
C34241 OR2X1_LOC_465/Y AND2X1_LOC_368/a_8_24# 0.23fF
C34242 OR2X1_LOC_632/A OR2X1_LOC_630/Y 0.06fF
C34243 OR2X1_LOC_115/a_36_216# OR2X1_LOC_78/A 0.02fF
C34244 AND2X1_LOC_91/B OR2X1_LOC_19/B 0.09fF
C34245 OR2X1_LOC_744/A OR2X1_LOC_118/Y 0.03fF
C34246 OR2X1_LOC_854/A OR2X1_LOC_568/A 0.99fF
C34247 AND2X1_LOC_12/Y OR2X1_LOC_363/A 0.03fF
C34248 AND2X1_LOC_756/a_8_24# OR2X1_LOC_616/Y 0.01fF
C34249 AND2X1_LOC_303/A OR2X1_LOC_51/Y 0.09fF
C34250 VDD OR2X1_LOC_97/B 0.21fF
C34251 AND2X1_LOC_849/A AND2X1_LOC_287/B 0.19fF
C34252 AND2X1_LOC_110/Y OR2X1_LOC_778/Y 0.05fF
C34253 OR2X1_LOC_80/A OR2X1_LOC_398/Y 0.00fF
C34254 OR2X1_LOC_96/Y OR2X1_LOC_6/a_36_216# 0.00fF
C34255 AND2X1_LOC_593/a_8_24# OR2X1_LOC_89/A 0.01fF
C34256 AND2X1_LOC_71/a_8_24# OR2X1_LOC_161/A 0.01fF
C34257 AND2X1_LOC_716/Y AND2X1_LOC_841/B 0.07fF
C34258 OR2X1_LOC_700/a_8_216# OR2X1_LOC_44/Y 0.01fF
C34259 OR2X1_LOC_773/B OR2X1_LOC_756/B 0.01fF
C34260 AND2X1_LOC_711/Y AND2X1_LOC_469/Y 0.03fF
C34261 OR2X1_LOC_653/Y AND2X1_LOC_58/a_36_24# 0.00fF
C34262 AND2X1_LOC_40/Y OR2X1_LOC_847/A 0.00fF
C34263 AND2X1_LOC_773/Y OR2X1_LOC_416/Y 0.03fF
C34264 OR2X1_LOC_634/A OR2X1_LOC_375/A 0.22fF
C34265 AND2X1_LOC_831/a_8_24# AND2X1_LOC_219/Y 0.01fF
C34266 OR2X1_LOC_231/A OR2X1_LOC_61/Y 0.03fF
C34267 OR2X1_LOC_323/A AND2X1_LOC_270/a_8_24# 0.01fF
C34268 AND2X1_LOC_40/Y OR2X1_LOC_288/a_8_216# 0.01fF
C34269 OR2X1_LOC_417/A AND2X1_LOC_241/a_8_24# 0.04fF
C34270 AND2X1_LOC_364/Y OR2X1_LOC_6/A 0.01fF
C34271 OR2X1_LOC_435/B OR2X1_LOC_130/A 0.02fF
C34272 AND2X1_LOC_768/a_36_24# AND2X1_LOC_361/A 0.01fF
C34273 OR2X1_LOC_808/B OR2X1_LOC_448/Y 0.10fF
C34274 OR2X1_LOC_185/Y OR2X1_LOC_538/A 0.34fF
C34275 OR2X1_LOC_665/Y OR2X1_LOC_51/Y 0.15fF
C34276 OR2X1_LOC_51/Y AND2X1_LOC_474/Y 0.02fF
C34277 OR2X1_LOC_154/A OR2X1_LOC_499/B 0.04fF
C34278 OR2X1_LOC_216/A OR2X1_LOC_510/Y 0.00fF
C34279 AND2X1_LOC_687/B OR2X1_LOC_12/Y 0.11fF
C34280 OR2X1_LOC_744/A OR2X1_LOC_262/Y 0.00fF
C34281 OR2X1_LOC_62/B OR2X1_LOC_161/B 0.03fF
C34282 OR2X1_LOC_426/A OR2X1_LOC_427/a_8_216# 0.01fF
C34283 AND2X1_LOC_729/B AND2X1_LOC_194/Y 0.01fF
C34284 AND2X1_LOC_520/a_8_24# OR2X1_LOC_417/A 0.01fF
C34285 OR2X1_LOC_702/A OR2X1_LOC_66/A 0.04fF
C34286 AND2X1_LOC_47/Y OR2X1_LOC_563/A 0.03fF
C34287 OR2X1_LOC_485/A OR2X1_LOC_51/Y 0.41fF
C34288 AND2X1_LOC_565/a_8_24# AND2X1_LOC_578/A 0.02fF
C34289 OR2X1_LOC_175/B OR2X1_LOC_539/Y 0.00fF
C34290 OR2X1_LOC_53/Y OR2X1_LOC_409/B 0.00fF
C34291 OR2X1_LOC_158/A AND2X1_LOC_687/A 0.01fF
C34292 OR2X1_LOC_694/a_8_216# OR2X1_LOC_427/A 0.07fF
C34293 OR2X1_LOC_130/A OR2X1_LOC_61/Y 0.21fF
C34294 AND2X1_LOC_513/a_8_24# OR2X1_LOC_26/Y 0.01fF
C34295 AND2X1_LOC_715/Y OR2X1_LOC_760/a_8_216# 0.23fF
C34296 AND2X1_LOC_831/Y AND2X1_LOC_786/Y 0.01fF
C34297 OR2X1_LOC_780/B OR2X1_LOC_161/B 0.23fF
C34298 OR2X1_LOC_807/B OR2X1_LOC_807/A 0.19fF
C34299 AND2X1_LOC_560/B OR2X1_LOC_92/Y 0.10fF
C34300 OR2X1_LOC_837/B OR2X1_LOC_6/A 0.26fF
C34301 OR2X1_LOC_216/A OR2X1_LOC_810/A 0.16fF
C34302 AND2X1_LOC_486/Y OR2X1_LOC_283/Y 0.03fF
C34303 OR2X1_LOC_95/Y OR2X1_LOC_373/Y 0.03fF
C34304 OR2X1_LOC_160/A AND2X1_LOC_43/B 0.02fF
C34305 OR2X1_LOC_54/Y INPUT_2 0.23fF
C34306 AND2X1_LOC_392/A AND2X1_LOC_327/a_36_24# 0.01fF
C34307 AND2X1_LOC_367/A OR2X1_LOC_74/A 0.10fF
C34308 OR2X1_LOC_814/A AND2X1_LOC_265/a_8_24# 0.04fF
C34309 OR2X1_LOC_476/B OR2X1_LOC_66/A 0.02fF
C34310 OR2X1_LOC_256/a_8_216# OR2X1_LOC_85/A 0.05fF
C34311 OR2X1_LOC_479/Y AND2X1_LOC_526/a_8_24# 0.05fF
C34312 AND2X1_LOC_392/A OR2X1_LOC_22/Y 0.10fF
C34313 OR2X1_LOC_313/a_8_216# OR2X1_LOC_314/Y 0.40fF
C34314 OR2X1_LOC_8/Y OR2X1_LOC_611/a_8_216# 0.14fF
C34315 OR2X1_LOC_217/Y OR2X1_LOC_507/B 0.03fF
C34316 OR2X1_LOC_768/A AND2X1_LOC_51/Y 0.00fF
C34317 OR2X1_LOC_650/Y OR2X1_LOC_66/A 0.02fF
C34318 AND2X1_LOC_123/Y AND2X1_LOC_572/A 0.81fF
C34319 OR2X1_LOC_585/A OR2X1_LOC_586/a_36_216# 0.00fF
C34320 INPUT_4 OR2X1_LOC_427/a_8_216# 0.00fF
C34321 AND2X1_LOC_576/Y AND2X1_LOC_621/Y 0.07fF
C34322 OR2X1_LOC_364/A AND2X1_LOC_12/Y 0.07fF
C34323 OR2X1_LOC_215/Y OR2X1_LOC_222/A 0.05fF
C34324 AND2X1_LOC_586/a_36_24# AND2X1_LOC_56/B 0.01fF
C34325 AND2X1_LOC_339/B AND2X1_LOC_649/Y 0.00fF
C34326 VDD OR2X1_LOC_814/A 2.61fF
C34327 OR2X1_LOC_135/Y AND2X1_LOC_660/A 0.01fF
C34328 OR2X1_LOC_499/B OR2X1_LOC_778/A 1.33fF
C34329 OR2X1_LOC_185/Y AND2X1_LOC_12/Y 6.10fF
C34330 OR2X1_LOC_287/B OR2X1_LOC_814/a_36_216# 0.00fF
C34331 OR2X1_LOC_312/Y AND2X1_LOC_841/B 0.03fF
C34332 OR2X1_LOC_520/B AND2X1_LOC_92/Y 0.01fF
C34333 OR2X1_LOC_358/a_8_216# OR2X1_LOC_154/A 0.02fF
C34334 AND2X1_LOC_560/B OR2X1_LOC_65/B 0.07fF
C34335 AND2X1_LOC_53/Y AND2X1_LOC_18/Y 0.08fF
C34336 OR2X1_LOC_714/a_8_216# OR2X1_LOC_724/A 0.01fF
C34337 AND2X1_LOC_619/a_8_24# OR2X1_LOC_80/A 0.01fF
C34338 AND2X1_LOC_235/a_8_24# OR2X1_LOC_68/B 0.07fF
C34339 OR2X1_LOC_664/a_36_216# OR2X1_LOC_631/B 0.01fF
C34340 OR2X1_LOC_715/B OR2X1_LOC_241/Y 0.98fF
C34341 OR2X1_LOC_426/B INPUT_1 0.07fF
C34342 OR2X1_LOC_252/Y OR2X1_LOC_627/a_8_216# 0.01fF
C34343 AND2X1_LOC_553/a_8_24# AND2X1_LOC_227/Y 0.01fF
C34344 OR2X1_LOC_528/Y AND2X1_LOC_866/A 0.21fF
C34345 AND2X1_LOC_36/Y OR2X1_LOC_71/A 0.07fF
C34346 AND2X1_LOC_599/a_8_24# AND2X1_LOC_761/a_8_24# 0.23fF
C34347 OR2X1_LOC_139/A OR2X1_LOC_801/B 0.02fF
C34348 AND2X1_LOC_44/Y OR2X1_LOC_194/a_8_216# 0.03fF
C34349 OR2X1_LOC_563/A OR2X1_LOC_598/A 0.02fF
C34350 OR2X1_LOC_799/A OR2X1_LOC_593/A 0.11fF
C34351 OR2X1_LOC_167/Y AND2X1_LOC_436/Y 0.26fF
C34352 AND2X1_LOC_76/a_36_24# OR2X1_LOC_74/A 0.00fF
C34353 OR2X1_LOC_446/B OR2X1_LOC_308/Y 0.05fF
C34354 OR2X1_LOC_32/Y OR2X1_LOC_39/A 0.23fF
C34355 AND2X1_LOC_70/Y OR2X1_LOC_446/Y 0.16fF
C34356 OR2X1_LOC_692/a_8_216# OR2X1_LOC_64/Y 0.15fF
C34357 OR2X1_LOC_85/A AND2X1_LOC_838/a_8_24# 0.01fF
C34358 AND2X1_LOC_154/a_8_24# OR2X1_LOC_7/A 0.07fF
C34359 OR2X1_LOC_64/Y OR2X1_LOC_92/Y 0.28fF
C34360 OR2X1_LOC_600/A AND2X1_LOC_476/A 0.07fF
C34361 OR2X1_LOC_406/A AND2X1_LOC_785/Y 0.03fF
C34362 GATE_479 AND2X1_LOC_480/A 0.24fF
C34363 OR2X1_LOC_680/A AND2X1_LOC_474/Y 0.03fF
C34364 OR2X1_LOC_18/Y AND2X1_LOC_651/B 0.00fF
C34365 OR2X1_LOC_671/a_36_216# D_INPUT_2 0.03fF
C34366 OR2X1_LOC_802/Y OR2X1_LOC_810/A 0.02fF
C34367 OR2X1_LOC_161/B OR2X1_LOC_365/B 0.01fF
C34368 OR2X1_LOC_164/Y AND2X1_LOC_471/a_8_24# 0.07fF
C34369 OR2X1_LOC_3/Y AND2X1_LOC_123/Y 0.04fF
C34370 OR2X1_LOC_680/A OR2X1_LOC_485/A 0.48fF
C34371 AND2X1_LOC_59/Y AND2X1_LOC_42/B 0.07fF
C34372 OR2X1_LOC_827/Y OR2X1_LOC_85/A 0.00fF
C34373 OR2X1_LOC_69/Y OR2X1_LOC_52/B 0.01fF
C34374 OR2X1_LOC_132/Y OR2X1_LOC_95/Y 0.07fF
C34375 AND2X1_LOC_374/Y AND2X1_LOC_458/a_8_24# 0.00fF
C34376 AND2X1_LOC_840/B OR2X1_LOC_238/Y 0.00fF
C34377 OR2X1_LOC_84/Y OR2X1_LOC_786/a_8_216# 0.07fF
C34378 OR2X1_LOC_306/a_8_216# AND2X1_LOC_729/B 0.01fF
C34379 OR2X1_LOC_185/A OR2X1_LOC_473/Y 0.16fF
C34380 OR2X1_LOC_624/A OR2X1_LOC_215/A 0.01fF
C34381 OR2X1_LOC_764/Y OR2X1_LOC_44/Y 0.01fF
C34382 OR2X1_LOC_864/A OR2X1_LOC_774/Y 0.00fF
C34383 AND2X1_LOC_658/B OR2X1_LOC_47/Y 0.03fF
C34384 OR2X1_LOC_121/B OR2X1_LOC_493/A 0.10fF
C34385 AND2X1_LOC_70/Y OR2X1_LOC_473/A 0.15fF
C34386 AND2X1_LOC_498/a_8_24# OR2X1_LOC_276/B 0.01fF
C34387 OR2X1_LOC_517/A OR2X1_LOC_71/Y 0.03fF
C34388 AND2X1_LOC_59/Y OR2X1_LOC_705/Y 0.32fF
C34389 AND2X1_LOC_738/B AND2X1_LOC_803/a_8_24# 0.03fF
C34390 OR2X1_LOC_89/A AND2X1_LOC_264/a_8_24# 0.02fF
C34391 OR2X1_LOC_864/A OR2X1_LOC_633/B 0.07fF
C34392 OR2X1_LOC_479/Y OR2X1_LOC_87/A 0.17fF
C34393 AND2X1_LOC_702/Y OR2X1_LOC_299/Y 0.01fF
C34394 AND2X1_LOC_663/B OR2X1_LOC_39/A -0.01fF
C34395 OR2X1_LOC_64/Y OR2X1_LOC_65/B 0.08fF
C34396 OR2X1_LOC_92/Y OR2X1_LOC_417/A 0.10fF
C34397 OR2X1_LOC_160/A AND2X1_LOC_698/a_8_24# 0.03fF
C34398 OR2X1_LOC_380/Y OR2X1_LOC_588/A 0.10fF
C34399 AND2X1_LOC_712/B AND2X1_LOC_454/Y 0.00fF
C34400 AND2X1_LOC_675/Y AND2X1_LOC_675/a_8_24# 0.01fF
C34401 AND2X1_LOC_197/a_8_24# OR2X1_LOC_6/A 0.02fF
C34402 AND2X1_LOC_673/a_8_24# OR2X1_LOC_74/A 0.17fF
C34403 AND2X1_LOC_584/a_8_24# AND2X1_LOC_51/Y 0.01fF
C34404 OR2X1_LOC_742/B OR2X1_LOC_550/a_8_216# 0.02fF
C34405 OR2X1_LOC_653/Y OR2X1_LOC_532/B 0.01fF
C34406 OR2X1_LOC_759/A AND2X1_LOC_846/a_8_24# 0.01fF
C34407 OR2X1_LOC_709/A OR2X1_LOC_513/Y 0.00fF
C34408 OR2X1_LOC_694/a_8_216# AND2X1_LOC_687/B 0.02fF
C34409 AND2X1_LOC_95/Y INPUT_1 0.02fF
C34410 AND2X1_LOC_801/B AND2X1_LOC_801/a_8_24# 0.07fF
C34411 OR2X1_LOC_756/B OR2X1_LOC_112/B 0.02fF
C34412 OR2X1_LOC_655/a_8_216# OR2X1_LOC_655/B 0.08fF
C34413 OR2X1_LOC_31/Y OR2X1_LOC_40/a_8_216# 0.01fF
C34414 AND2X1_LOC_290/a_36_24# D_INPUT_0 0.00fF
C34415 OR2X1_LOC_858/A AND2X1_LOC_72/B 0.03fF
C34416 AND2X1_LOC_530/a_36_24# OR2X1_LOC_80/A 0.00fF
C34417 AND2X1_LOC_154/Y OR2X1_LOC_743/A 0.01fF
C34418 AND2X1_LOC_566/Y AND2X1_LOC_568/a_8_24# 0.06fF
C34419 OR2X1_LOC_607/a_8_216# OR2X1_LOC_619/Y 0.04fF
C34420 OR2X1_LOC_335/B OR2X1_LOC_375/A 0.01fF
C34421 AND2X1_LOC_633/Y AND2X1_LOC_633/a_36_24# 0.01fF
C34422 AND2X1_LOC_859/B OR2X1_LOC_278/Y 0.04fF
C34423 OR2X1_LOC_11/Y OR2X1_LOC_429/a_8_216# 0.39fF
C34424 OR2X1_LOC_192/A OR2X1_LOC_192/B 0.06fF
C34425 AND2X1_LOC_456/B AND2X1_LOC_721/A 0.04fF
C34426 AND2X1_LOC_59/Y OR2X1_LOC_286/B 0.08fF
C34427 AND2X1_LOC_174/a_8_24# OR2X1_LOC_31/Y 0.09fF
C34428 OR2X1_LOC_177/Y OR2X1_LOC_164/a_8_216# 0.01fF
C34429 OR2X1_LOC_254/B OR2X1_LOC_532/B 0.09fF
C34430 OR2X1_LOC_137/B AND2X1_LOC_47/Y 0.01fF
C34431 OR2X1_LOC_26/Y OR2X1_LOC_46/A 0.33fF
C34432 AND2X1_LOC_70/Y OR2X1_LOC_228/Y 0.03fF
C34433 AND2X1_LOC_537/Y OR2X1_LOC_52/B 4.21fF
C34434 AND2X1_LOC_835/a_8_24# OR2X1_LOC_85/A 0.01fF
C34435 AND2X1_LOC_476/A OR2X1_LOC_619/Y 0.07fF
C34436 AND2X1_LOC_438/a_8_24# OR2X1_LOC_544/B 0.03fF
C34437 AND2X1_LOC_631/a_36_24# OR2X1_LOC_615/Y 0.00fF
C34438 OR2X1_LOC_363/a_8_216# OR2X1_LOC_366/A -0.00fF
C34439 OR2X1_LOC_417/A AND2X1_LOC_464/a_36_24# 0.01fF
C34440 OR2X1_LOC_447/Y OR2X1_LOC_269/B 0.10fF
C34441 OR2X1_LOC_89/A OR2X1_LOC_46/A 0.05fF
C34442 OR2X1_LOC_151/A OR2X1_LOC_788/B 0.12fF
C34443 OR2X1_LOC_532/Y OR2X1_LOC_356/A 0.05fF
C34444 OR2X1_LOC_755/A OR2X1_LOC_665/a_8_216# 0.49fF
C34445 INPUT_7 INPUT_6 0.16fF
C34446 AND2X1_LOC_3/Y OR2X1_LOC_720/B 0.03fF
C34447 OR2X1_LOC_646/A OR2X1_LOC_532/B 0.02fF
C34448 AND2X1_LOC_227/Y OR2X1_LOC_26/Y 0.09fF
C34449 AND2X1_LOC_566/a_8_24# AND2X1_LOC_170/B 0.01fF
C34450 OR2X1_LOC_488/Y AND2X1_LOC_849/A 0.09fF
C34451 AND2X1_LOC_681/a_8_24# OR2X1_LOC_87/A 0.01fF
C34452 OR2X1_LOC_743/A INPUT_1 0.48fF
C34453 AND2X1_LOC_851/B OR2X1_LOC_44/Y 0.07fF
C34454 OR2X1_LOC_185/A OR2X1_LOC_241/B 0.04fF
C34455 OR2X1_LOC_151/A OR2X1_LOC_175/a_8_216# 0.04fF
C34456 OR2X1_LOC_605/B OR2X1_LOC_335/B 0.00fF
C34457 AND2X1_LOC_64/Y OR2X1_LOC_855/A 0.15fF
C34458 AND2X1_LOC_866/A AND2X1_LOC_105/a_8_24# 0.06fF
C34459 D_INPUT_3 OR2X1_LOC_670/Y 0.01fF
C34460 OR2X1_LOC_31/Y OR2X1_LOC_238/Y 0.02fF
C34461 OR2X1_LOC_3/Y OR2X1_LOC_813/A 0.00fF
C34462 OR2X1_LOC_510/Y OR2X1_LOC_205/Y 0.25fF
C34463 AND2X1_LOC_741/a_8_24# AND2X1_LOC_222/Y 0.01fF
C34464 AND2X1_LOC_227/Y OR2X1_LOC_89/A 0.08fF
C34465 AND2X1_LOC_64/Y AND2X1_LOC_627/a_8_24# 0.01fF
C34466 AND2X1_LOC_798/a_8_24# AND2X1_LOC_810/B 0.03fF
C34467 AND2X1_LOC_564/B OR2X1_LOC_406/Y 0.02fF
C34468 AND2X1_LOC_41/A OR2X1_LOC_725/a_8_216# 0.05fF
C34469 OR2X1_LOC_827/a_8_216# D_INPUT_1 0.01fF
C34470 OR2X1_LOC_465/B OR2X1_LOC_270/Y 0.00fF
C34471 AND2X1_LOC_31/Y OR2X1_LOC_784/Y 0.01fF
C34472 OR2X1_LOC_316/a_8_216# OR2X1_LOC_158/A 0.02fF
C34473 OR2X1_LOC_125/Y INPUT_1 0.04fF
C34474 OR2X1_LOC_559/B OR2X1_LOC_559/a_36_216# 0.02fF
C34475 AND2X1_LOC_711/Y AND2X1_LOC_663/a_8_24# 0.01fF
C34476 OR2X1_LOC_26/Y OR2X1_LOC_813/Y 0.07fF
C34477 OR2X1_LOC_246/A INPUT_1 0.10fF
C34478 OR2X1_LOC_155/A AND2X1_LOC_418/a_8_24# 0.03fF
C34479 AND2X1_LOC_7/B AND2X1_LOC_256/a_8_24# 0.01fF
C34480 OR2X1_LOC_318/A AND2X1_LOC_22/Y 0.00fF
C34481 OR2X1_LOC_26/Y OR2X1_LOC_41/Y 0.13fF
C34482 OR2X1_LOC_858/A AND2X1_LOC_36/Y 0.02fF
C34483 OR2X1_LOC_696/A OR2X1_LOC_536/Y 0.08fF
C34484 OR2X1_LOC_45/B AND2X1_LOC_795/a_8_24# 0.01fF
C34485 AND2X1_LOC_849/A OR2X1_LOC_95/Y 0.03fF
C34486 AND2X1_LOC_12/Y OR2X1_LOC_578/B 0.03fF
C34487 OR2X1_LOC_186/Y OR2X1_LOC_355/A 0.01fF
C34488 AND2X1_LOC_358/Y OR2X1_LOC_16/A 0.14fF
C34489 INPUT_1 OR2X1_LOC_225/a_8_216# 0.06fF
C34490 OR2X1_LOC_59/Y AND2X1_LOC_791/a_36_24# 0.00fF
C34491 AND2X1_LOC_104/a_36_24# OR2X1_LOC_80/A 0.00fF
C34492 AND2X1_LOC_512/a_36_24# OR2X1_LOC_599/Y 0.00fF
C34493 AND2X1_LOC_72/a_8_24# OR2X1_LOC_247/Y 0.23fF
C34494 AND2X1_LOC_40/Y OR2X1_LOC_544/B 0.01fF
C34495 OR2X1_LOC_59/Y OR2X1_LOC_759/Y 0.01fF
C34496 OR2X1_LOC_446/a_8_216# OR2X1_LOC_446/A 0.47fF
C34497 OR2X1_LOC_92/Y AND2X1_LOC_247/a_8_24# 0.01fF
C34498 AND2X1_LOC_22/Y OR2X1_LOC_151/A 0.03fF
C34499 AND2X1_LOC_91/B AND2X1_LOC_110/Y 0.03fF
C34500 AND2X1_LOC_476/A AND2X1_LOC_462/a_8_24# 0.02fF
C34501 OR2X1_LOC_788/a_8_216# OR2X1_LOC_788/B 0.07fF
C34502 OR2X1_LOC_632/Y OR2X1_LOC_500/a_36_216# 0.01fF
C34503 OR2X1_LOC_87/A OR2X1_LOC_68/B 3.45fF
C34504 AND2X1_LOC_841/B OR2X1_LOC_13/B 0.07fF
C34505 OR2X1_LOC_144/Y OR2X1_LOC_142/Y 0.06fF
C34506 OR2X1_LOC_732/B OR2X1_LOC_317/B 0.79fF
C34507 OR2X1_LOC_89/A OR2X1_LOC_753/Y 0.01fF
C34508 OR2X1_LOC_74/A AND2X1_LOC_647/Y 0.03fF
C34509 OR2X1_LOC_696/A AND2X1_LOC_474/A 0.03fF
C34510 OR2X1_LOC_59/Y OR2X1_LOC_767/Y 0.02fF
C34511 AND2X1_LOC_564/B OR2X1_LOC_496/a_8_216# 0.02fF
C34512 OR2X1_LOC_818/a_8_216# D_INPUT_3 0.08fF
C34513 OR2X1_LOC_246/Y OR2X1_LOC_71/A 0.01fF
C34514 OR2X1_LOC_759/A GATE_579 0.00fF
C34515 OR2X1_LOC_709/B OR2X1_LOC_709/a_8_216# 0.06fF
C34516 OR2X1_LOC_377/A OR2X1_LOC_376/Y 0.06fF
C34517 OR2X1_LOC_707/A OR2X1_LOC_707/a_8_216# 0.47fF
C34518 AND2X1_LOC_19/a_8_24# OR2X1_LOC_68/B 0.00fF
C34519 AND2X1_LOC_831/Y AND2X1_LOC_841/a_8_24# 0.03fF
C34520 OR2X1_LOC_190/A OR2X1_LOC_577/Y 0.06fF
C34521 OR2X1_LOC_53/Y AND2X1_LOC_691/a_36_24# 0.00fF
C34522 OR2X1_LOC_3/Y OR2X1_LOC_377/a_8_216# 0.02fF
C34523 OR2X1_LOC_308/A AND2X1_LOC_41/A 0.01fF
C34524 OR2X1_LOC_468/A OR2X1_LOC_161/B 0.03fF
C34525 OR2X1_LOC_801/a_8_216# OR2X1_LOC_138/A 0.01fF
C34526 OR2X1_LOC_45/B AND2X1_LOC_434/Y 0.07fF
C34527 OR2X1_LOC_46/A AND2X1_LOC_202/a_8_24# 0.01fF
C34528 AND2X1_LOC_555/Y AND2X1_LOC_360/a_8_24# 0.01fF
C34529 AND2X1_LOC_516/a_8_24# OR2X1_LOC_446/B 0.01fF
C34530 AND2X1_LOC_721/Y AND2X1_LOC_471/Y 0.01fF
C34531 OR2X1_LOC_45/B AND2X1_LOC_219/Y 0.39fF
C34532 OR2X1_LOC_591/Y OR2X1_LOC_604/A 0.02fF
C34533 AND2X1_LOC_672/a_8_24# OR2X1_LOC_673/A 0.01fF
C34534 AND2X1_LOC_657/Y AND2X1_LOC_212/Y 0.10fF
C34535 INPUT_0 AND2X1_LOC_44/Y 0.09fF
C34536 OR2X1_LOC_528/Y OR2X1_LOC_40/Y 0.05fF
C34537 OR2X1_LOC_166/a_36_216# OR2X1_LOC_16/A 0.03fF
C34538 OR2X1_LOC_486/Y OR2X1_LOC_787/B 0.22fF
C34539 OR2X1_LOC_6/B OR2X1_LOC_631/A 0.00fF
C34540 OR2X1_LOC_858/a_8_216# OR2X1_LOC_349/A 0.01fF
C34541 AND2X1_LOC_51/Y OR2X1_LOC_513/a_36_216# 0.02fF
C34542 OR2X1_LOC_78/B OR2X1_LOC_633/A 0.02fF
C34543 OR2X1_LOC_56/a_36_216# OR2X1_LOC_16/Y 0.00fF
C34544 AND2X1_LOC_212/Y AND2X1_LOC_469/B 0.01fF
C34545 OR2X1_LOC_857/B OR2X1_LOC_35/Y 0.30fF
C34546 INPUT_4 INPUT_6 0.04fF
C34547 OR2X1_LOC_267/Y OR2X1_LOC_721/Y 0.03fF
C34548 OR2X1_LOC_198/a_36_216# AND2X1_LOC_95/Y 0.01fF
C34549 OR2X1_LOC_369/Y AND2X1_LOC_181/Y 0.03fF
C34550 OR2X1_LOC_696/A AND2X1_LOC_593/Y 0.00fF
C34551 AND2X1_LOC_722/a_36_24# OR2X1_LOC_40/Y 0.00fF
C34552 OR2X1_LOC_369/a_8_216# OR2X1_LOC_309/Y 0.01fF
C34553 AND2X1_LOC_64/Y OR2X1_LOC_319/a_8_216# 0.06fF
C34554 VDD OR2X1_LOC_410/Y 0.16fF
C34555 AND2X1_LOC_727/Y OR2X1_LOC_427/A 0.03fF
C34556 AND2X1_LOC_56/B OR2X1_LOC_308/Y 0.07fF
C34557 OR2X1_LOC_158/A OR2X1_LOC_90/a_8_216# 0.02fF
C34558 OR2X1_LOC_323/A AND2X1_LOC_717/a_36_24# 0.00fF
C34559 OR2X1_LOC_114/B OR2X1_LOC_842/A 0.02fF
C34560 AND2X1_LOC_64/Y OR2X1_LOC_377/A 0.15fF
C34561 AND2X1_LOC_12/Y OR2X1_LOC_366/A 0.01fF
C34562 AND2X1_LOC_716/Y AND2X1_LOC_364/a_8_24# 0.01fF
C34563 OR2X1_LOC_696/A OR2X1_LOC_85/A 0.06fF
C34564 OR2X1_LOC_151/A OR2X1_LOC_244/B 1.22fF
C34565 OR2X1_LOC_409/Y AND2X1_LOC_463/B 0.78fF
C34566 OR2X1_LOC_862/a_36_216# OR2X1_LOC_812/B 0.00fF
C34567 VDD OR2X1_LOC_244/Y 0.38fF
C34568 AND2X1_LOC_51/A INPUT_6 0.03fF
C34569 OR2X1_LOC_188/Y OR2X1_LOC_185/A 0.02fF
C34570 AND2X1_LOC_572/a_8_24# AND2X1_LOC_573/A 0.03fF
C34571 OR2X1_LOC_178/Y VDD 0.21fF
C34572 AND2X1_LOC_541/a_8_24# OR2X1_LOC_65/B -0.00fF
C34573 OR2X1_LOC_369/a_8_216# OR2X1_LOC_744/A 0.03fF
C34574 VDD OR2X1_LOC_192/A -0.00fF
C34575 AND2X1_LOC_437/a_8_24# OR2X1_LOC_66/A 0.01fF
C34576 VDD OR2X1_LOC_715/A 0.12fF
C34577 OR2X1_LOC_467/B OR2X1_LOC_477/Y 0.14fF
C34578 INPUT_0 OR2X1_LOC_600/A 0.07fF
C34579 OR2X1_LOC_39/Y AND2X1_LOC_194/Y 0.01fF
C34580 AND2X1_LOC_759/a_8_24# OR2X1_LOC_792/B 0.01fF
C34581 AND2X1_LOC_64/Y OR2X1_LOC_203/Y 0.07fF
C34582 OR2X1_LOC_375/A OR2X1_LOC_267/Y 0.03fF
C34583 OR2X1_LOC_40/Y AND2X1_LOC_512/Y 0.01fF
C34584 VDD OR2X1_LOC_501/B 0.03fF
C34585 OR2X1_LOC_160/B OR2X1_LOC_235/B 0.03fF
C34586 OR2X1_LOC_196/Y AND2X1_LOC_43/B 0.02fF
C34587 OR2X1_LOC_715/B OR2X1_LOC_216/A 0.07fF
C34588 AND2X1_LOC_367/A AND2X1_LOC_860/A 0.07fF
C34589 OR2X1_LOC_52/B OR2X1_LOC_743/Y 0.00fF
C34590 AND2X1_LOC_70/Y AND2X1_LOC_498/a_8_24# 0.01fF
C34591 OR2X1_LOC_127/Y OR2X1_LOC_428/A 0.01fF
C34592 OR2X1_LOC_589/A OR2X1_LOC_393/a_8_216# 0.39fF
C34593 AND2X1_LOC_121/a_36_24# OR2X1_LOC_56/A 0.00fF
C34594 OR2X1_LOC_128/a_8_216# AND2X1_LOC_44/Y 0.01fF
C34595 OR2X1_LOC_834/A OR2X1_LOC_78/A 0.01fF
C34596 OR2X1_LOC_348/a_8_216# OR2X1_LOC_260/a_8_216# 0.47fF
C34597 OR2X1_LOC_345/Y OR2X1_LOC_260/Y 0.72fF
C34598 OR2X1_LOC_589/A AND2X1_LOC_654/Y 0.07fF
C34599 OR2X1_LOC_240/A OR2X1_LOC_397/a_8_216# 0.16fF
C34600 AND2X1_LOC_711/Y OR2X1_LOC_759/Y 0.01fF
C34601 OR2X1_LOC_468/A OR2X1_LOC_435/B 0.02fF
C34602 AND2X1_LOC_477/A OR2X1_LOC_437/A 0.05fF
C34603 OR2X1_LOC_484/Y OR2X1_LOC_59/Y 0.51fF
C34604 OR2X1_LOC_482/Y AND2X1_LOC_840/A 0.17fF
C34605 OR2X1_LOC_3/B OR2X1_LOC_70/A 0.22fF
C34606 AND2X1_LOC_535/a_8_24# AND2X1_LOC_512/Y 0.02fF
C34607 VDD OR2X1_LOC_256/Y 0.35fF
C34608 OR2X1_LOC_377/A AND2X1_LOC_82/Y 0.27fF
C34609 AND2X1_LOC_139/B AND2X1_LOC_786/Y 0.07fF
C34610 AND2X1_LOC_727/A OR2X1_LOC_142/a_36_216# 0.00fF
C34611 AND2X1_LOC_543/Y OR2X1_LOC_312/Y 0.63fF
C34612 OR2X1_LOC_122/a_8_216# AND2X1_LOC_474/A 0.01fF
C34613 AND2X1_LOC_362/B AND2X1_LOC_97/a_8_24# 0.01fF
C34614 OR2X1_LOC_151/A OR2X1_LOC_630/a_8_216# 0.02fF
C34615 OR2X1_LOC_502/A AND2X1_LOC_18/Y 2.19fF
C34616 OR2X1_LOC_375/A OR2X1_LOC_633/A 0.11fF
C34617 AND2X1_LOC_40/Y OR2X1_LOC_440/a_8_216# 0.01fF
C34618 OR2X1_LOC_426/B OR2X1_LOC_517/A 0.17fF
C34619 OR2X1_LOC_236/a_8_216# OR2X1_LOC_428/A 0.01fF
C34620 OR2X1_LOC_375/A OR2X1_LOC_725/A 0.01fF
C34621 INPUT_5 OR2X1_LOC_380/a_8_216# 0.05fF
C34622 AND2X1_LOC_860/a_8_24# AND2X1_LOC_858/B 0.02fF
C34623 AND2X1_LOC_773/Y OR2X1_LOC_6/A 0.01fF
C34624 AND2X1_LOC_3/Y OR2X1_LOC_554/a_8_216# 0.01fF
C34625 VDD OR2X1_LOC_147/B 0.80fF
C34626 OR2X1_LOC_339/Y OR2X1_LOC_358/A 0.06fF
C34627 OR2X1_LOC_45/B OR2X1_LOC_496/Y 0.61fF
C34628 AND2X1_LOC_565/B OR2X1_LOC_189/a_36_216# 0.00fF
C34629 OR2X1_LOC_673/a_8_216# OR2X1_LOC_375/A 0.01fF
C34630 D_INPUT_0 OR2X1_LOC_217/A 0.01fF
C34631 OR2X1_LOC_187/a_36_216# AND2X1_LOC_191/B 0.00fF
C34632 AND2X1_LOC_592/Y OR2X1_LOC_424/a_8_216# 0.01fF
C34633 OR2X1_LOC_335/a_8_216# OR2X1_LOC_605/A 0.47fF
C34634 AND2X1_LOC_72/B OR2X1_LOC_736/a_36_216# 0.00fF
C34635 AND2X1_LOC_57/a_8_24# OR2X1_LOC_35/Y 0.01fF
C34636 VDD AND2X1_LOC_517/a_8_24# 0.00fF
C34637 AND2X1_LOC_337/a_8_24# AND2X1_LOC_654/Y 0.02fF
C34638 OR2X1_LOC_449/B OR2X1_LOC_161/B 9.84fF
C34639 AND2X1_LOC_658/A AND2X1_LOC_804/Y 0.03fF
C34640 OR2X1_LOC_524/Y OR2X1_LOC_441/Y 0.09fF
C34641 OR2X1_LOC_91/Y AND2X1_LOC_182/A 0.02fF
C34642 AND2X1_LOC_31/Y OR2X1_LOC_451/B 0.04fF
C34643 AND2X1_LOC_392/A AND2X1_LOC_661/a_36_24# 0.01fF
C34644 AND2X1_LOC_528/a_8_24# AND2X1_LOC_44/Y 0.03fF
C34645 AND2X1_LOC_90/a_8_24# AND2X1_LOC_8/Y 0.01fF
C34646 AND2X1_LOC_721/a_36_24# OR2X1_LOC_59/Y 0.00fF
C34647 OR2X1_LOC_51/Y OR2X1_LOC_256/a_8_216# 0.05fF
C34648 OR2X1_LOC_267/A AND2X1_LOC_65/A 0.79fF
C34649 OR2X1_LOC_56/A OR2X1_LOC_278/Y 0.03fF
C34650 AND2X1_LOC_392/A OR2X1_LOC_39/A 0.07fF
C34651 AND2X1_LOC_70/Y OR2X1_LOC_635/a_8_216# 0.01fF
C34652 OR2X1_LOC_715/B OR2X1_LOC_802/Y 0.35fF
C34653 OR2X1_LOC_67/a_36_216# AND2X1_LOC_243/Y 0.01fF
C34654 AND2X1_LOC_654/B OR2X1_LOC_762/Y 0.25fF
C34655 AND2X1_LOC_729/Y OR2X1_LOC_526/Y 0.03fF
C34656 AND2X1_LOC_662/B OR2X1_LOC_56/A 0.03fF
C34657 OR2X1_LOC_604/A AND2X1_LOC_317/a_8_24# 0.01fF
C34658 OR2X1_LOC_523/Y OR2X1_LOC_632/Y 0.13fF
C34659 AND2X1_LOC_95/Y OR2X1_LOC_287/A 0.03fF
C34660 OR2X1_LOC_710/B AND2X1_LOC_59/Y 0.09fF
C34661 OR2X1_LOC_6/A AND2X1_LOC_243/Y 0.02fF
C34662 OR2X1_LOC_400/A AND2X1_LOC_18/Y 0.01fF
C34663 OR2X1_LOC_405/A OR2X1_LOC_778/B 0.05fF
C34664 VDD AND2X1_LOC_470/A 0.25fF
C34665 AND2X1_LOC_486/Y AND2X1_LOC_562/B 0.03fF
C34666 AND2X1_LOC_40/Y OR2X1_LOC_190/B 0.29fF
C34667 INPUT_0 OR2X1_LOC_619/Y 0.07fF
C34668 OR2X1_LOC_861/a_36_216# OR2X1_LOC_756/B 0.00fF
C34669 OR2X1_LOC_312/Y OR2X1_LOC_322/Y 0.15fF
C34670 OR2X1_LOC_719/Y OR2X1_LOC_733/A 0.21fF
C34671 D_INPUT_5 AND2X1_LOC_53/a_8_24# 0.10fF
C34672 OR2X1_LOC_151/A OR2X1_LOC_296/a_8_216# -0.01fF
C34673 AND2X1_LOC_787/a_8_24# OR2X1_LOC_516/B 0.01fF
C34674 OR2X1_LOC_45/B OR2X1_LOC_119/a_8_216# 0.01fF
C34675 INPUT_3 OR2X1_LOC_235/B 0.01fF
C34676 AND2X1_LOC_95/Y OR2X1_LOC_174/A 0.01fF
C34677 AND2X1_LOC_504/a_8_24# AND2X1_LOC_41/A 0.04fF
C34678 AND2X1_LOC_560/B OR2X1_LOC_600/A 0.07fF
C34679 OR2X1_LOC_185/A AND2X1_LOC_189/a_8_24# 0.00fF
C34680 OR2X1_LOC_696/A OR2X1_LOC_226/Y 0.21fF
C34681 OR2X1_LOC_493/Y OR2X1_LOC_558/a_8_216# 0.05fF
C34682 AND2X1_LOC_564/B AND2X1_LOC_465/Y 0.01fF
C34683 OR2X1_LOC_748/A AND2X1_LOC_711/A 0.27fF
C34684 AND2X1_LOC_92/Y OR2X1_LOC_350/a_36_216# 0.00fF
C34685 AND2X1_LOC_474/A AND2X1_LOC_474/a_8_24# -0.00fF
C34686 OR2X1_LOC_528/Y OR2X1_LOC_7/A 0.14fF
C34687 AND2X1_LOC_2/Y AND2X1_LOC_25/Y 0.20fF
C34688 AND2X1_LOC_95/Y OR2X1_LOC_435/a_8_216# 0.01fF
C34689 OR2X1_LOC_600/A OR2X1_LOC_690/A 0.03fF
C34690 AND2X1_LOC_404/B AND2X1_LOC_404/a_8_24# 0.01fF
C34691 OR2X1_LOC_137/Y AND2X1_LOC_18/Y -0.02fF
C34692 OR2X1_LOC_495/a_8_216# OR2X1_LOC_51/Y 0.01fF
C34693 OR2X1_LOC_62/B OR2X1_LOC_554/a_36_216# 0.00fF
C34694 AND2X1_LOC_91/B AND2X1_LOC_494/a_36_24# -0.02fF
C34695 OR2X1_LOC_462/B OR2X1_LOC_78/A 0.00fF
C34696 OR2X1_LOC_494/a_36_216# OR2X1_LOC_625/Y 0.01fF
C34697 OR2X1_LOC_676/Y OR2X1_LOC_155/A 0.03fF
C34698 AND2X1_LOC_392/A AND2X1_LOC_211/B 0.10fF
C34699 OR2X1_LOC_121/B OR2X1_LOC_161/B 0.19fF
C34700 AND2X1_LOC_520/Y AND2X1_LOC_642/Y 0.01fF
C34701 AND2X1_LOC_115/a_8_24# OR2X1_LOC_428/A 0.16fF
C34702 OR2X1_LOC_692/Y OR2X1_LOC_64/Y 0.04fF
C34703 AND2X1_LOC_576/Y OR2X1_LOC_59/Y 0.07fF
C34704 VDD OR2X1_LOC_383/a_8_216# 0.00fF
C34705 OR2X1_LOC_158/A AND2X1_LOC_660/Y 0.07fF
C34706 OR2X1_LOC_808/B OR2X1_LOC_803/B 0.73fF
C34707 AND2X1_LOC_566/B AND2X1_LOC_212/B 0.01fF
C34708 OR2X1_LOC_364/A OR2X1_LOC_168/B 0.01fF
C34709 OR2X1_LOC_135/Y AND2X1_LOC_307/Y 0.19fF
C34710 AND2X1_LOC_308/a_36_24# OR2X1_LOC_428/A 0.01fF
C34711 OR2X1_LOC_848/B OR2X1_LOC_391/A 0.07fF
C34712 OR2X1_LOC_416/Y OR2X1_LOC_12/Y 0.06fF
C34713 AND2X1_LOC_649/B AND2X1_LOC_649/a_8_24# 0.01fF
C34714 AND2X1_LOC_725/a_8_24# OR2X1_LOC_3/Y 0.00fF
C34715 AND2X1_LOC_729/a_8_24# OR2X1_LOC_64/Y 0.01fF
C34716 OR2X1_LOC_809/B OR2X1_LOC_810/A 0.03fF
C34717 AND2X1_LOC_691/a_8_24# OR2X1_LOC_585/A 0.01fF
C34718 VDD AND2X1_LOC_387/B 0.18fF
C34719 AND2X1_LOC_535/Y OR2X1_LOC_70/Y 0.01fF
C34720 OR2X1_LOC_160/B OR2X1_LOC_844/a_8_216# 0.01fF
C34721 OR2X1_LOC_834/A OR2X1_LOC_155/A 0.03fF
C34722 AND2X1_LOC_784/A OR2X1_LOC_310/Y 0.03fF
C34723 AND2X1_LOC_640/a_8_24# AND2X1_LOC_219/A 0.01fF
C34724 OR2X1_LOC_517/Y OR2X1_LOC_517/A 0.01fF
C34725 OR2X1_LOC_107/Y OR2X1_LOC_26/Y 0.02fF
C34726 OR2X1_LOC_166/Y OR2X1_LOC_312/Y 0.09fF
C34727 OR2X1_LOC_798/Y OR2X1_LOC_802/A 0.13fF
C34728 OR2X1_LOC_32/B OR2X1_LOC_23/a_8_216# 0.43fF
C34729 AND2X1_LOC_711/a_36_24# OR2X1_LOC_748/A 0.00fF
C34730 VDD OR2X1_LOC_258/Y 0.12fF
C34731 OR2X1_LOC_599/A AND2X1_LOC_718/a_8_24# -0.00fF
C34732 OR2X1_LOC_757/A OR2X1_LOC_665/Y 0.01fF
C34733 AND2X1_LOC_337/B OR2X1_LOC_56/A 0.06fF
C34734 OR2X1_LOC_863/B OR2X1_LOC_66/A 0.02fF
C34735 OR2X1_LOC_31/Y AND2X1_LOC_208/Y 0.00fF
C34736 AND2X1_LOC_365/A AND2X1_LOC_654/Y 0.08fF
C34737 AND2X1_LOC_40/Y OR2X1_LOC_285/A 0.00fF
C34738 AND2X1_LOC_492/a_8_24# OR2X1_LOC_805/A 0.03fF
C34739 OR2X1_LOC_126/a_8_216# OR2X1_LOC_744/A 0.01fF
C34740 AND2X1_LOC_59/Y OR2X1_LOC_76/B 0.00fF
C34741 VDD AND2X1_LOC_484/a_8_24# 0.00fF
C34742 OR2X1_LOC_240/B OR2X1_LOC_240/a_8_216# 0.06fF
C34743 AND2X1_LOC_474/A OR2X1_LOC_89/a_8_216# 0.01fF
C34744 OR2X1_LOC_516/A AND2X1_LOC_794/A 0.03fF
C34745 OR2X1_LOC_447/A AND2X1_LOC_43/B 0.41fF
C34746 OR2X1_LOC_185/A OR2X1_LOC_405/Y 0.00fF
C34747 OR2X1_LOC_600/A OR2X1_LOC_64/Y 0.07fF
C34748 AND2X1_LOC_335/Y OR2X1_LOC_64/Y 0.03fF
C34749 OR2X1_LOC_159/a_8_216# OR2X1_LOC_54/Y 0.40fF
C34750 AND2X1_LOC_716/Y OR2X1_LOC_43/A 0.07fF
C34751 OR2X1_LOC_756/B OR2X1_LOC_574/A 0.03fF
C34752 AND2X1_LOC_512/Y OR2X1_LOC_7/A 0.07fF
C34753 OR2X1_LOC_40/Y OR2X1_LOC_54/Y 0.08fF
C34754 OR2X1_LOC_624/A OR2X1_LOC_539/Y 0.03fF
C34755 OR2X1_LOC_329/B AND2X1_LOC_473/a_8_24# 0.01fF
C34756 OR2X1_LOC_744/A OR2X1_LOC_83/a_8_216# 0.01fF
C34757 OR2X1_LOC_45/B AND2X1_LOC_851/B 0.06fF
C34758 AND2X1_LOC_2/Y AND2X1_LOC_51/Y 0.01fF
C34759 AND2X1_LOC_453/Y AND2X1_LOC_454/Y 0.14fF
C34760 OR2X1_LOC_756/B OR2X1_LOC_33/A 0.01fF
C34761 AND2X1_LOC_101/B OR2X1_LOC_92/Y 0.51fF
C34762 OR2X1_LOC_185/Y OR2X1_LOC_860/a_8_216# 0.01fF
C34763 OR2X1_LOC_70/Y OR2X1_LOC_484/Y 0.07fF
C34764 AND2X1_LOC_722/A OR2X1_LOC_89/A 0.03fF
C34765 AND2X1_LOC_70/Y OR2X1_LOC_76/A 0.00fF
C34766 AND2X1_LOC_31/Y AND2X1_LOC_36/Y 5.99fF
C34767 AND2X1_LOC_48/A AND2X1_LOC_18/Y 0.60fF
C34768 OR2X1_LOC_49/A OR2X1_LOC_62/A 0.51fF
C34769 OR2X1_LOC_3/Y OR2X1_LOC_292/Y 0.01fF
C34770 OR2X1_LOC_43/A AND2X1_LOC_654/Y 0.07fF
C34771 OR2X1_LOC_563/A D_INPUT_1 0.03fF
C34772 AND2X1_LOC_293/a_36_24# AND2X1_LOC_219/A 0.00fF
C34773 OR2X1_LOC_106/a_8_216# AND2X1_LOC_845/Y 0.02fF
C34774 AND2X1_LOC_12/Y AND2X1_LOC_817/B 0.01fF
C34775 AND2X1_LOC_36/Y OR2X1_LOC_715/a_8_216# 0.01fF
C34776 OR2X1_LOC_654/A D_INPUT_5 0.01fF
C34777 OR2X1_LOC_479/Y OR2X1_LOC_804/a_36_216# 0.01fF
C34778 AND2X1_LOC_50/Y D_INPUT_7 0.01fF
C34779 INPUT_0 AND2X1_LOC_4/a_36_24# 0.00fF
C34780 AND2X1_LOC_319/A AND2X1_LOC_452/Y 0.01fF
C34781 AND2X1_LOC_327/a_8_24# OR2X1_LOC_59/Y 0.01fF
C34782 OR2X1_LOC_253/a_8_216# OR2X1_LOC_56/A 0.03fF
C34783 AND2X1_LOC_784/A OR2X1_LOC_519/a_8_216# 0.06fF
C34784 OR2X1_LOC_844/B OR2X1_LOC_68/B 0.04fF
C34785 AND2X1_LOC_557/Y AND2X1_LOC_572/Y 0.19fF
C34786 OR2X1_LOC_641/Y AND2X1_LOC_518/a_36_24# 0.00fF
C34787 OR2X1_LOC_154/A OR2X1_LOC_659/a_8_216# 0.06fF
C34788 AND2X1_LOC_859/Y OR2X1_LOC_18/Y 0.00fF
C34789 OR2X1_LOC_19/B OR2X1_LOC_56/A 0.24fF
C34790 AND2X1_LOC_741/Y GATE_479 0.15fF
C34791 OR2X1_LOC_364/A AND2X1_LOC_59/Y 0.07fF
C34792 OR2X1_LOC_212/B OR2X1_LOC_357/A 0.85fF
C34793 OR2X1_LOC_415/Y OR2X1_LOC_598/A 0.20fF
C34794 OR2X1_LOC_185/Y AND2X1_LOC_59/Y 0.14fF
C34795 AND2X1_LOC_251/a_8_24# OR2X1_LOC_579/B 0.04fF
C34796 OR2X1_LOC_316/Y OR2X1_LOC_36/Y 0.02fF
C34797 AND2X1_LOC_838/Y AND2X1_LOC_852/a_8_24# 0.11fF
C34798 AND2X1_LOC_17/Y OR2X1_LOC_635/a_8_216# 0.12fF
C34799 VDD OR2X1_LOC_545/B 0.21fF
C34800 OR2X1_LOC_641/Y OR2X1_LOC_520/A 0.03fF
C34801 OR2X1_LOC_161/A OR2X1_LOC_269/B 0.29fF
C34802 OR2X1_LOC_160/A AND2X1_LOC_159/a_8_24# 0.01fF
C34803 OR2X1_LOC_600/A OR2X1_LOC_417/A 0.42fF
C34804 AND2X1_LOC_656/a_8_24# AND2X1_LOC_772/Y 0.02fF
C34805 AND2X1_LOC_796/a_8_24# AND2X1_LOC_810/Y 0.07fF
C34806 OR2X1_LOC_160/A OR2X1_LOC_810/A 8.93fF
C34807 OR2X1_LOC_640/a_36_216# AND2X1_LOC_8/Y 0.00fF
C34808 AND2X1_LOC_25/Y AND2X1_LOC_26/a_8_24# 0.13fF
C34809 OR2X1_LOC_45/B OR2X1_LOC_595/Y 0.02fF
C34810 AND2X1_LOC_365/A OR2X1_LOC_312/Y 0.04fF
C34811 OR2X1_LOC_47/Y AND2X1_LOC_469/Y 0.04fF
C34812 AND2X1_LOC_471/a_8_24# AND2X1_LOC_471/Y 0.04fF
C34813 OR2X1_LOC_475/Y OR2X1_LOC_734/a_36_216# 0.00fF
C34814 OR2X1_LOC_62/B OR2X1_LOC_630/B 0.00fF
C34815 OR2X1_LOC_36/Y AND2X1_LOC_354/B 0.03fF
C34816 OR2X1_LOC_791/B OR2X1_LOC_287/B 0.02fF
C34817 OR2X1_LOC_297/Y AND2X1_LOC_847/Y 0.02fF
C34818 AND2X1_LOC_216/Y AND2X1_LOC_660/A 0.01fF
C34819 AND2X1_LOC_12/Y OR2X1_LOC_654/A 0.03fF
C34820 OR2X1_LOC_95/Y AND2X1_LOC_447/Y 0.01fF
C34821 OR2X1_LOC_473/A OR2X1_LOC_362/A 0.00fF
C34822 OR2X1_LOC_138/A OR2X1_LOC_801/B 0.13fF
C34823 OR2X1_LOC_303/B OR2X1_LOC_301/a_8_216# 0.02fF
C34824 OR2X1_LOC_160/B OR2X1_LOC_276/B 0.07fF
C34825 OR2X1_LOC_460/B OR2X1_LOC_460/a_8_216# 0.47fF
C34826 AND2X1_LOC_56/B AND2X1_LOC_472/B 0.00fF
C34827 OR2X1_LOC_51/Y OR2X1_LOC_238/a_8_216# 0.19fF
C34828 AND2X1_LOC_359/B OR2X1_LOC_248/a_36_216# 0.01fF
C34829 AND2X1_LOC_563/a_8_24# AND2X1_LOC_489/Y 0.02fF
C34830 OR2X1_LOC_517/A OR2X1_LOC_246/A 0.00fF
C34831 AND2X1_LOC_342/Y OR2X1_LOC_7/A 0.08fF
C34832 AND2X1_LOC_345/Y AND2X1_LOC_847/Y 0.02fF
C34833 VDD AND2X1_LOC_318/Y 0.51fF
C34834 OR2X1_LOC_599/A OR2X1_LOC_26/Y 0.09fF
C34835 D_INPUT_5 AND2X1_LOC_21/a_36_24# 0.00fF
C34836 AND2X1_LOC_95/Y OR2X1_LOC_476/Y 0.01fF
C34837 AND2X1_LOC_170/Y AND2X1_LOC_566/a_8_24# 0.01fF
C34838 OR2X1_LOC_235/B OR2X1_LOC_244/A 0.03fF
C34839 OR2X1_LOC_577/B D_GATE_366 0.03fF
C34840 AND2X1_LOC_47/Y OR2X1_LOC_632/Y 0.19fF
C34841 AND2X1_LOC_474/A AND2X1_LOC_849/a_8_24# 0.01fF
C34842 OR2X1_LOC_26/Y OR2X1_LOC_93/a_8_216# 0.07fF
C34843 OR2X1_LOC_312/Y OR2X1_LOC_43/A 0.03fF
C34844 AND2X1_LOC_12/Y AND2X1_LOC_496/a_36_24# 0.00fF
C34845 OR2X1_LOC_458/a_8_216# OR2X1_LOC_532/B 0.01fF
C34846 AND2X1_LOC_51/Y OR2X1_LOC_739/A 0.04fF
C34847 OR2X1_LOC_599/A OR2X1_LOC_89/A 1.08fF
C34848 OR2X1_LOC_744/A OR2X1_LOC_503/Y 0.10fF
C34849 AND2X1_LOC_191/Y AND2X1_LOC_576/Y 0.07fF
C34850 OR2X1_LOC_64/Y OR2X1_LOC_619/Y 0.04fF
C34851 OR2X1_LOC_485/A AND2X1_LOC_359/B 0.01fF
C34852 AND2X1_LOC_64/Y OR2X1_LOC_732/A 0.09fF
C34853 OR2X1_LOC_824/a_8_216# OR2X1_LOC_36/Y 0.09fF
C34854 AND2X1_LOC_702/Y OR2X1_LOC_3/Y 0.03fF
C34855 OR2X1_LOC_130/A AND2X1_LOC_67/Y 0.08fF
C34856 AND2X1_LOC_390/B OR2X1_LOC_36/Y 0.07fF
C34857 AND2X1_LOC_711/Y AND2X1_LOC_576/Y 0.07fF
C34858 AND2X1_LOC_17/Y AND2X1_LOC_386/a_8_24# 0.11fF
C34859 OR2X1_LOC_256/Y OR2X1_LOC_256/A 0.07fF
C34860 OR2X1_LOC_682/Y OR2X1_LOC_7/A 0.02fF
C34861 VDD OR2X1_LOC_815/Y 0.12fF
C34862 OR2X1_LOC_631/A OR2X1_LOC_598/A 0.03fF
C34863 OR2X1_LOC_168/a_8_216# OR2X1_LOC_168/A 0.47fF
C34864 OR2X1_LOC_655/a_8_216# OR2X1_LOC_655/A 0.39fF
C34865 AND2X1_LOC_7/B OR2X1_LOC_317/B 0.06fF
C34866 OR2X1_LOC_635/A OR2X1_LOC_614/a_8_216# -0.05fF
C34867 AND2X1_LOC_683/a_8_24# AND2X1_LOC_3/Y 0.02fF
C34868 AND2X1_LOC_663/B OR2X1_LOC_85/A 0.07fF
C34869 AND2X1_LOC_321/a_8_24# OR2X1_LOC_532/B 0.01fF
C34870 AND2X1_LOC_3/Y OR2X1_LOC_793/B 0.03fF
C34871 AND2X1_LOC_197/a_8_24# OR2X1_LOC_44/Y 0.01fF
C34872 AND2X1_LOC_65/A OR2X1_LOC_560/A 0.03fF
C34873 OR2X1_LOC_840/a_8_216# OR2X1_LOC_68/B 0.02fF
C34874 OR2X1_LOC_59/Y OR2X1_LOC_29/a_8_216# 0.01fF
C34875 OR2X1_LOC_89/A OR2X1_LOC_258/a_8_216# 0.01fF
C34876 OR2X1_LOC_762/a_8_216# OR2X1_LOC_44/Y 0.01fF
C34877 AND2X1_LOC_132/a_8_24# OR2X1_LOC_62/B 0.17fF
C34878 VDD OR2X1_LOC_318/B 0.05fF
C34879 OR2X1_LOC_431/Y OR2X1_LOC_36/Y 0.01fF
C34880 OR2X1_LOC_185/A D_INPUT_0 0.75fF
C34881 AND2X1_LOC_146/a_8_24# OR2X1_LOC_161/A 0.01fF
C34882 AND2X1_LOC_51/Y OR2X1_LOC_269/B 0.20fF
C34883 OR2X1_LOC_11/Y OR2X1_LOC_22/A 1.53fF
C34884 OR2X1_LOC_16/A OR2X1_LOC_71/A 0.10fF
C34885 AND2X1_LOC_525/a_8_24# OR2X1_LOC_546/B 0.01fF
C34886 AND2X1_LOC_483/a_8_24# OR2X1_LOC_7/A 0.18fF
C34887 OR2X1_LOC_481/Y AND2X1_LOC_259/Y 0.03fF
C34888 OR2X1_LOC_3/Y AND2X1_LOC_345/a_8_24# 0.01fF
C34889 AND2X1_LOC_56/B OR2X1_LOC_19/B 0.24fF
C34890 AND2X1_LOC_55/a_8_24# AND2X1_LOC_672/B 0.00fF
C34891 AND2X1_LOC_22/Y OR2X1_LOC_716/a_8_216# 0.01fF
C34892 OR2X1_LOC_510/A OR2X1_LOC_560/A 0.04fF
C34893 VDD OR2X1_LOC_854/A 0.00fF
C34894 OR2X1_LOC_160/B OR2X1_LOC_779/B 0.00fF
C34895 OR2X1_LOC_424/Y OR2X1_LOC_428/A 0.00fF
C34896 AND2X1_LOC_364/a_8_24# OR2X1_LOC_13/B 0.03fF
C34897 OR2X1_LOC_182/B OR2X1_LOC_578/B 0.04fF
C34898 OR2X1_LOC_109/Y OR2X1_LOC_95/Y 0.07fF
C34899 OR2X1_LOC_291/Y OR2X1_LOC_612/B 0.03fF
C34900 OR2X1_LOC_604/a_8_216# AND2X1_LOC_452/Y 0.01fF
C34901 OR2X1_LOC_532/B AND2X1_LOC_272/a_8_24# 0.01fF
C34902 OR2X1_LOC_820/Y AND2X1_LOC_847/a_8_24# 0.01fF
C34903 AND2X1_LOC_8/Y OR2X1_LOC_19/B 0.63fF
C34904 OR2X1_LOC_109/Y OR2X1_LOC_368/A 0.01fF
C34905 OR2X1_LOC_632/Y OR2X1_LOC_598/A 0.01fF
C34906 AND2X1_LOC_70/Y OR2X1_LOC_566/Y 0.09fF
C34907 OR2X1_LOC_492/a_8_216# OR2X1_LOC_437/A 0.01fF
C34908 OR2X1_LOC_447/Y OR2X1_LOC_779/a_8_216# 0.02fF
C34909 AND2X1_LOC_712/B OR2X1_LOC_7/A 0.17fF
C34910 OR2X1_LOC_696/A AND2X1_LOC_555/Y 0.02fF
C34911 OR2X1_LOC_516/Y AND2X1_LOC_564/B 0.07fF
C34912 OR2X1_LOC_7/A OR2X1_LOC_54/Y 0.65fF
C34913 AND2X1_LOC_62/a_8_24# D_INPUT_1 0.01fF
C34914 OR2X1_LOC_625/Y OR2X1_LOC_47/Y 0.11fF
C34915 OR2X1_LOC_589/A OR2X1_LOC_13/B 1.41fF
C34916 OR2X1_LOC_428/A D_INPUT_6 0.07fF
C34917 OR2X1_LOC_36/Y AND2X1_LOC_863/Y 0.01fF
C34918 AND2X1_LOC_110/Y OR2X1_LOC_446/B 0.03fF
C34919 AND2X1_LOC_729/Y OR2X1_LOC_760/Y 0.02fF
C34920 OR2X1_LOC_557/A OR2X1_LOC_403/a_8_216# 0.01fF
C34921 AND2X1_LOC_555/Y AND2X1_LOC_383/a_8_24# 0.01fF
C34922 OR2X1_LOC_476/B OR2X1_LOC_473/Y 0.00fF
C34923 AND2X1_LOC_866/A OR2X1_LOC_26/Y 0.03fF
C34924 OR2X1_LOC_730/B OR2X1_LOC_730/A 0.04fF
C34925 OR2X1_LOC_549/B OR2X1_LOC_563/A 0.18fF
C34926 AND2X1_LOC_178/a_8_24# OR2X1_LOC_192/B 0.21fF
C34927 AND2X1_LOC_54/a_8_24# OR2X1_LOC_80/A 0.03fF
C34928 AND2X1_LOC_350/Y AND2X1_LOC_351/Y 0.91fF
C34929 OR2X1_LOC_676/Y OR2X1_LOC_515/a_36_216# 0.01fF
C34930 OR2X1_LOC_600/A AND2X1_LOC_247/a_8_24# 0.03fF
C34931 OR2X1_LOC_635/A AND2X1_LOC_31/Y 0.00fF
C34932 AND2X1_LOC_576/Y OR2X1_LOC_184/Y 0.04fF
C34933 AND2X1_LOC_866/A OR2X1_LOC_89/A 0.06fF
C34934 OR2X1_LOC_22/Y OR2X1_LOC_43/a_8_216# 0.03fF
C34935 OR2X1_LOC_214/A AND2X1_LOC_44/Y 0.01fF
C34936 AND2X1_LOC_660/a_8_24# AND2X1_LOC_116/Y 0.01fF
C34937 OR2X1_LOC_844/Y OR2X1_LOC_859/A 0.01fF
C34938 OR2X1_LOC_506/B AND2X1_LOC_3/Y 0.14fF
C34939 OR2X1_LOC_288/A AND2X1_LOC_281/a_8_24# 0.23fF
C34940 OR2X1_LOC_166/Y OR2X1_LOC_13/B 0.03fF
C34941 OR2X1_LOC_518/Y AND2X1_LOC_339/B 0.14fF
C34942 AND2X1_LOC_537/Y OR2X1_LOC_22/Y 0.02fF
C34943 OR2X1_LOC_97/A OR2X1_LOC_139/A 0.03fF
C34944 AND2X1_LOC_7/B AND2X1_LOC_44/Y 0.70fF
C34945 AND2X1_LOC_729/B OR2X1_LOC_95/Y 0.00fF
C34946 AND2X1_LOC_707/Y OR2X1_LOC_428/A 0.10fF
C34947 OR2X1_LOC_421/A OR2X1_LOC_387/A 0.02fF
C34948 OR2X1_LOC_469/Y OR2X1_LOC_705/a_8_216# 0.12fF
C34949 OR2X1_LOC_31/Y OR2X1_LOC_52/Y 0.01fF
C34950 OR2X1_LOC_393/Y OR2X1_LOC_80/A 0.14fF
C34951 OR2X1_LOC_506/A OR2X1_LOC_724/A 0.00fF
C34952 AND2X1_LOC_59/Y OR2X1_LOC_568/A 0.02fF
C34953 AND2X1_LOC_744/a_8_24# OR2X1_LOC_712/B 0.01fF
C34954 AND2X1_LOC_212/Y AND2X1_LOC_804/A 0.01fF
C34955 AND2X1_LOC_413/a_36_24# OR2X1_LOC_598/A 0.00fF
C34956 AND2X1_LOC_92/Y OR2X1_LOC_308/Y 0.07fF
C34957 AND2X1_LOC_7/B OR2X1_LOC_514/a_8_216# 0.02fF
C34958 OR2X1_LOC_791/B OR2X1_LOC_345/a_8_216# 0.03fF
C34959 OR2X1_LOC_44/Y OR2X1_LOC_749/a_8_216# 0.01fF
C34960 AND2X1_LOC_654/B OR2X1_LOC_13/B 0.13fF
C34961 OR2X1_LOC_850/B OR2X1_LOC_349/B 0.00fF
C34962 OR2X1_LOC_434/a_8_216# OR2X1_LOC_174/Y 0.40fF
C34963 OR2X1_LOC_833/B AND2X1_LOC_268/a_8_24# 0.01fF
C34964 OR2X1_LOC_811/A OR2X1_LOC_366/Y 0.08fF
C34965 AND2X1_LOC_334/a_8_24# AND2X1_LOC_476/A 0.02fF
C34966 AND2X1_LOC_22/Y AND2X1_LOC_300/a_8_24# 0.00fF
C34967 OR2X1_LOC_344/A OR2X1_LOC_578/a_8_216# 0.01fF
C34968 OR2X1_LOC_696/A OR2X1_LOC_51/Y 0.21fF
C34969 OR2X1_LOC_160/B AND2X1_LOC_226/a_8_24# 0.01fF
C34970 OR2X1_LOC_247/Y AND2X1_LOC_3/Y 0.01fF
C34971 OR2X1_LOC_64/a_8_216# OR2X1_LOC_22/A 0.03fF
C34972 OR2X1_LOC_158/A OR2X1_LOC_310/a_8_216# 0.01fF
C34973 OR2X1_LOC_97/A OR2X1_LOC_654/a_36_216# 0.00fF
C34974 AND2X1_LOC_118/a_36_24# OR2X1_LOC_598/A 0.01fF
C34975 OR2X1_LOC_633/A OR2X1_LOC_549/A 0.17fF
C34976 OR2X1_LOC_22/A OR2X1_LOC_409/a_36_216# 0.00fF
C34977 OR2X1_LOC_323/A OR2X1_LOC_56/A 0.69fF
C34978 AND2X1_LOC_565/B AND2X1_LOC_564/A 0.04fF
C34979 AND2X1_LOC_611/a_8_24# OR2X1_LOC_68/B 0.02fF
C34980 AND2X1_LOC_64/Y OR2X1_LOC_78/B 0.77fF
C34981 AND2X1_LOC_365/A OR2X1_LOC_13/B 0.01fF
C34982 AND2X1_LOC_667/a_8_24# OR2X1_LOC_786/Y 0.01fF
C34983 OR2X1_LOC_805/A OR2X1_LOC_580/A 0.07fF
C34984 AND2X1_LOC_489/Y AND2X1_LOC_563/Y 0.01fF
C34985 OR2X1_LOC_13/a_8_216# OR2X1_LOC_13/Y 0.01fF
C34986 OR2X1_LOC_134/Y OR2X1_LOC_91/A 0.24fF
C34987 OR2X1_LOC_207/B AND2X1_LOC_18/Y 0.35fF
C34988 OR2X1_LOC_49/A OR2X1_LOC_8/Y 0.19fF
C34989 AND2X1_LOC_60/a_8_24# OR2X1_LOC_648/A 0.01fF
C34990 OR2X1_LOC_769/A AND2X1_LOC_22/Y 0.07fF
C34991 AND2X1_LOC_850/Y OR2X1_LOC_504/a_8_216# 0.03fF
C34992 AND2X1_LOC_719/Y AND2X1_LOC_476/Y 0.10fF
C34993 OR2X1_LOC_709/A OR2X1_LOC_160/B 0.13fF
C34994 AND2X1_LOC_672/a_36_24# AND2X1_LOC_47/Y 0.00fF
C34995 OR2X1_LOC_375/A OR2X1_LOC_590/Y 0.01fF
C34996 OR2X1_LOC_121/Y VDD 0.81fF
C34997 AND2X1_LOC_244/A OR2X1_LOC_59/Y 0.03fF
C34998 OR2X1_LOC_294/Y OR2X1_LOC_66/A 0.03fF
C34999 AND2X1_LOC_64/Y OR2X1_LOC_721/Y 0.05fF
C35000 VDD OR2X1_LOC_829/A 0.62fF
C35001 OR2X1_LOC_198/a_8_216# OR2X1_LOC_856/B 0.04fF
C35002 OR2X1_LOC_43/A OR2X1_LOC_13/B 7.97fF
C35003 OR2X1_LOC_604/A OR2X1_LOC_765/a_8_216# 0.01fF
C35004 OR2X1_LOC_585/A OR2X1_LOC_399/a_36_216# 0.00fF
C35005 AND2X1_LOC_22/Y OR2X1_LOC_174/A 0.28fF
C35006 OR2X1_LOC_263/a_8_216# AND2X1_LOC_647/Y 0.01fF
C35007 OR2X1_LOC_59/Y OR2X1_LOC_16/A 0.54fF
C35008 OR2X1_LOC_351/B VDD 0.18fF
C35009 AND2X1_LOC_22/Y OR2X1_LOC_435/a_8_216# 0.01fF
C35010 OR2X1_LOC_188/Y OR2X1_LOC_833/a_8_216# 0.04fF
C35011 AND2X1_LOC_82/Y OR2X1_LOC_78/B 0.10fF
C35012 AND2X1_LOC_787/A OR2X1_LOC_516/B 0.03fF
C35013 OR2X1_LOC_61/a_8_216# AND2X1_LOC_7/B 0.05fF
C35014 OR2X1_LOC_510/Y OR2X1_LOC_130/Y 0.00fF
C35015 OR2X1_LOC_139/A OR2X1_LOC_475/B 5.07fF
C35016 OR2X1_LOC_158/A AND2X1_LOC_434/Y 0.07fF
C35017 OR2X1_LOC_715/B OR2X1_LOC_809/B 0.15fF
C35018 OR2X1_LOC_759/A VDD 0.22fF
C35019 OR2X1_LOC_47/Y OR2X1_LOC_3/B 0.77fF
C35020 OR2X1_LOC_649/a_8_216# OR2X1_LOC_68/B 0.05fF
C35021 OR2X1_LOC_438/Y OR2X1_LOC_373/Y 0.33fF
C35022 OR2X1_LOC_186/Y OR2X1_LOC_808/B 0.89fF
C35023 OR2X1_LOC_160/B AND2X1_LOC_70/Y 0.20fF
C35024 OR2X1_LOC_607/Y AND2X1_LOC_647/Y 0.02fF
C35025 OR2X1_LOC_223/A OR2X1_LOC_804/A 0.01fF
C35026 AND2X1_LOC_64/Y OR2X1_LOC_375/A 0.13fF
C35027 AND2X1_LOC_95/Y OR2X1_LOC_563/A 0.14fF
C35028 OR2X1_LOC_240/A AND2X1_LOC_36/Y 0.02fF
C35029 OR2X1_LOC_108/Y OR2X1_LOC_59/Y 0.37fF
C35030 OR2X1_LOC_44/Y AND2X1_LOC_792/a_8_24# 0.00fF
C35031 AND2X1_LOC_91/B AND2X1_LOC_601/a_8_24# 0.04fF
C35032 OR2X1_LOC_633/B AND2X1_LOC_36/Y 0.06fF
C35033 AND2X1_LOC_596/a_8_24# OR2X1_LOC_744/A 0.01fF
C35034 OR2X1_LOC_18/Y GATE_579 0.00fF
C35035 OR2X1_LOC_856/B OR2X1_LOC_161/B 0.04fF
C35036 OR2X1_LOC_436/B OR2X1_LOC_390/A 0.00fF
C35037 OR2X1_LOC_135/Y OR2X1_LOC_427/A 0.01fF
C35038 VDD OR2X1_LOC_538/A 0.21fF
C35039 OR2X1_LOC_597/Y AND2X1_LOC_644/a_8_24# 0.23fF
C35040 OR2X1_LOC_151/A AND2X1_LOC_173/a_8_24# 0.04fF
C35041 AND2X1_LOC_465/Y OR2X1_LOC_437/A 0.00fF
C35042 OR2X1_LOC_502/A OR2X1_LOC_307/A 0.06fF
C35043 OR2X1_LOC_51/Y AND2X1_LOC_851/a_36_24# 0.00fF
C35044 AND2X1_LOC_56/B OR2X1_LOC_828/Y 0.01fF
C35045 AND2X1_LOC_621/Y OR2X1_LOC_373/Y 0.06fF
C35046 OR2X1_LOC_805/A AND2X1_LOC_44/Y 0.03fF
C35047 VDD OR2X1_LOC_698/Y 0.33fF
C35048 OR2X1_LOC_96/Y OR2X1_LOC_92/Y 0.00fF
C35049 AND2X1_LOC_306/a_8_24# OR2X1_LOC_78/A 0.01fF
C35050 OR2X1_LOC_574/A OR2X1_LOC_140/B 0.00fF
C35051 VDD D_INPUT_5 0.13fF
C35052 AND2X1_LOC_773/Y AND2X1_LOC_831/a_8_24# 0.04fF
C35053 OR2X1_LOC_603/a_8_216# OR2X1_LOC_603/Y -0.00fF
C35054 OR2X1_LOC_45/B OR2X1_LOC_372/Y 0.01fF
C35055 OR2X1_LOC_315/a_36_216# OR2X1_LOC_315/Y 0.03fF
C35056 AND2X1_LOC_366/A AND2X1_LOC_474/A 0.01fF
C35057 OR2X1_LOC_92/Y AND2X1_LOC_454/a_8_24# 0.02fF
C35058 OR2X1_LOC_465/B AND2X1_LOC_7/B 0.49fF
C35059 AND2X1_LOC_452/Y OR2X1_LOC_765/a_36_216# 0.00fF
C35060 OR2X1_LOC_6/A OR2X1_LOC_12/Y 0.46fF
C35061 OR2X1_LOC_715/B OR2X1_LOC_160/A 0.21fF
C35062 VDD AND2X1_LOC_178/a_8_24# -0.00fF
C35063 AND2X1_LOC_431/a_8_24# OR2X1_LOC_339/A 0.11fF
C35064 OR2X1_LOC_695/a_8_216# OR2X1_LOC_51/Y 0.01fF
C35065 AND2X1_LOC_865/A AND2X1_LOC_865/a_36_24# 0.01fF
C35066 OR2X1_LOC_696/A AND2X1_LOC_855/a_36_24# 0.01fF
C35067 OR2X1_LOC_49/A OR2X1_LOC_672/Y 0.01fF
C35068 AND2X1_LOC_285/Y OR2X1_LOC_278/Y 0.03fF
C35069 AND2X1_LOC_392/A AND2X1_LOC_593/Y 0.03fF
C35070 OR2X1_LOC_100/a_8_216# VDD 0.00fF
C35071 OR2X1_LOC_379/Y OR2X1_LOC_66/A 0.14fF
C35072 OR2X1_LOC_68/B OR2X1_LOC_493/Y 5.15fF
C35073 AND2X1_LOC_555/Y AND2X1_LOC_663/B 0.01fF
C35074 AND2X1_LOC_86/Y AND2X1_LOC_70/Y 0.02fF
C35075 AND2X1_LOC_637/a_8_24# OR2X1_LOC_586/Y 0.00fF
C35076 AND2X1_LOC_563/A AND2X1_LOC_572/Y 0.00fF
C35077 AND2X1_LOC_199/A OR2X1_LOC_43/A 0.01fF
C35078 OR2X1_LOC_279/Y AND2X1_LOC_284/a_8_24# 0.04fF
C35079 AND2X1_LOC_12/Y VDD 1.32fF
C35080 OR2X1_LOC_299/a_8_216# OR2X1_LOC_12/Y 0.01fF
C35081 OR2X1_LOC_528/Y OR2X1_LOC_406/a_36_216# 0.01fF
C35082 OR2X1_LOC_232/a_36_216# OR2X1_LOC_16/A 0.03fF
C35083 OR2X1_LOC_759/A OR2X1_LOC_616/Y 0.01fF
C35084 OR2X1_LOC_296/a_36_216# OR2X1_LOC_161/B 0.00fF
C35085 OR2X1_LOC_296/Y AND2X1_LOC_44/Y 0.05fF
C35086 VDD AND2X1_LOC_470/B 0.02fF
C35087 OR2X1_LOC_22/Y OR2X1_LOC_171/a_8_216# 0.03fF
C35088 VDD AND2X1_LOC_838/Y 0.20fF
C35089 OR2X1_LOC_743/A AND2X1_LOC_774/A 0.10fF
C35090 OR2X1_LOC_790/a_8_216# AND2X1_LOC_18/Y 0.01fF
C35091 OR2X1_LOC_44/Y AND2X1_LOC_243/Y 0.17fF
C35092 AND2X1_LOC_110/Y AND2X1_LOC_56/B 0.05fF
C35093 OR2X1_LOC_185/A OR2X1_LOC_795/B 0.01fF
C35094 OR2X1_LOC_151/A AND2X1_LOC_329/a_8_24# 0.02fF
C35095 AND2X1_LOC_860/A AND2X1_LOC_287/Y 0.01fF
C35096 OR2X1_LOC_365/a_8_216# OR2X1_LOC_365/B 0.07fF
C35097 AND2X1_LOC_510/A AND2X1_LOC_624/A 0.03fF
C35098 AND2X1_LOC_70/Y OR2X1_LOC_553/A 0.03fF
C35099 AND2X1_LOC_712/Y OR2X1_LOC_52/B 0.03fF
C35100 OR2X1_LOC_40/Y OR2X1_LOC_26/Y 6.02fF
C35101 AND2X1_LOC_802/B AND2X1_LOC_802/a_8_24# 0.10fF
C35102 OR2X1_LOC_467/A OR2X1_LOC_453/a_36_216# 0.00fF
C35103 AND2X1_LOC_40/Y OR2X1_LOC_608/a_8_216# 0.19fF
C35104 AND2X1_LOC_568/B OR2X1_LOC_44/Y 0.07fF
C35105 OR2X1_LOC_70/Y OR2X1_LOC_16/A 0.34fF
C35106 AND2X1_LOC_577/a_36_24# AND2X1_LOC_577/Y 0.00fF
C35107 AND2X1_LOC_658/B AND2X1_LOC_576/Y 0.07fF
C35108 AND2X1_LOC_570/Y AND2X1_LOC_580/A 0.03fF
C35109 OR2X1_LOC_640/a_36_216# AND2X1_LOC_92/Y 0.00fF
C35110 OR2X1_LOC_64/Y AND2X1_LOC_769/Y 0.03fF
C35111 OR2X1_LOC_468/A OR2X1_LOC_593/a_36_216# 0.00fF
C35112 OR2X1_LOC_842/a_8_216# AND2X1_LOC_95/Y 0.07fF
C35113 OR2X1_LOC_287/B OR2X1_LOC_362/A 0.06fF
C35114 OR2X1_LOC_7/A OR2X1_LOC_765/Y 0.02fF
C35115 AND2X1_LOC_318/Y AND2X1_LOC_269/a_8_24# 0.01fF
C35116 AND2X1_LOC_390/a_8_24# AND2X1_LOC_645/A 0.03fF
C35117 AND2X1_LOC_605/Y AND2X1_LOC_452/Y 0.01fF
C35118 OR2X1_LOC_426/A OR2X1_LOC_427/Y 0.56fF
C35119 OR2X1_LOC_756/B OR2X1_LOC_377/A 0.66fF
C35120 OR2X1_LOC_526/Y OR2X1_LOC_52/B 0.03fF
C35121 AND2X1_LOC_570/Y AND2X1_LOC_579/a_8_24# 0.02fF
C35122 OR2X1_LOC_656/B OR2X1_LOC_216/A 0.03fF
C35123 OR2X1_LOC_40/Y OR2X1_LOC_89/A 0.16fF
C35124 AND2X1_LOC_3/Y AND2X1_LOC_18/Y 0.38fF
C35125 OR2X1_LOC_744/A OR2X1_LOC_36/Y 0.48fF
C35126 OR2X1_LOC_756/B AND2X1_LOC_824/B 0.46fF
C35127 AND2X1_LOC_40/Y OR2X1_LOC_185/A 0.51fF
C35128 OR2X1_LOC_338/a_8_216# AND2X1_LOC_51/Y 0.01fF
C35129 OR2X1_LOC_178/a_8_216# OR2X1_LOC_485/A 0.01fF
C35130 OR2X1_LOC_690/a_8_216# INPUT_0 0.08fF
C35131 VDD AND2X1_LOC_79/Y 0.03fF
C35132 OR2X1_LOC_856/B AND2X1_LOC_536/a_8_24# 0.04fF
C35133 OR2X1_LOC_512/A OR2X1_LOC_375/A 0.04fF
C35134 OR2X1_LOC_405/A OR2X1_LOC_620/Y 0.07fF
C35135 OR2X1_LOC_92/Y AND2X1_LOC_449/Y 0.01fF
C35136 AND2X1_LOC_465/a_36_24# OR2X1_LOC_108/Y 0.00fF
C35137 OR2X1_LOC_417/Y OR2X1_LOC_421/Y 0.03fF
C35138 OR2X1_LOC_639/B D_INPUT_4 0.23fF
C35139 AND2X1_LOC_365/a_8_24# AND2X1_LOC_661/A 0.09fF
C35140 OR2X1_LOC_837/Y OR2X1_LOC_6/A 0.02fF
C35141 OR2X1_LOC_485/A AND2X1_LOC_436/Y 0.02fF
C35142 VDD OR2X1_LOC_804/B 0.27fF
C35143 OR2X1_LOC_185/Y AND2X1_LOC_67/a_36_24# 0.01fF
C35144 OR2X1_LOC_585/A OR2X1_LOC_597/a_36_216# 0.00fF
C35145 OR2X1_LOC_614/Y OR2X1_LOC_196/B 0.00fF
C35146 OR2X1_LOC_527/a_8_216# OR2X1_LOC_64/Y 0.08fF
C35147 AND2X1_LOC_161/a_8_24# OR2X1_LOC_619/Y 0.00fF
C35148 AND2X1_LOC_546/a_8_24# AND2X1_LOC_621/Y 0.03fF
C35149 OR2X1_LOC_744/A AND2X1_LOC_493/a_36_24# 0.01fF
C35150 OR2X1_LOC_786/Y OR2X1_LOC_115/B 0.00fF
C35151 OR2X1_LOC_6/B OR2X1_LOC_656/a_8_216# 0.02fF
C35152 OR2X1_LOC_160/B OR2X1_LOC_404/Y 0.11fF
C35153 OR2X1_LOC_427/A AND2X1_LOC_848/Y 0.03fF
C35154 OR2X1_LOC_91/Y AND2X1_LOC_723/a_8_24# 0.02fF
C35155 OR2X1_LOC_256/Y OR2X1_LOC_248/Y 0.52fF
C35156 OR2X1_LOC_22/Y OR2X1_LOC_13/Y 0.19fF
C35157 OR2X1_LOC_633/a_8_216# OR2X1_LOC_633/B 0.02fF
C35158 AND2X1_LOC_72/B OR2X1_LOC_501/A 0.02fF
C35159 AND2X1_LOC_497/a_36_24# OR2X1_LOC_844/B 0.00fF
C35160 OR2X1_LOC_32/Y OR2X1_LOC_58/a_8_216# 0.00fF
C35161 AND2X1_LOC_852/a_8_24# AND2X1_LOC_852/B 0.04fF
C35162 AND2X1_LOC_95/Y OR2X1_LOC_137/B 0.26fF
C35163 OR2X1_LOC_161/A OR2X1_LOC_347/B 0.12fF
C35164 AND2X1_LOC_12/Y AND2X1_LOC_755/a_8_24# 0.01fF
C35165 AND2X1_LOC_48/A OR2X1_LOC_596/a_36_216# 0.02fF
C35166 OR2X1_LOC_364/A OR2X1_LOC_794/A 0.03fF
C35167 OR2X1_LOC_251/a_8_216# OR2X1_LOC_106/A 0.01fF
C35168 OR2X1_LOC_51/Y AND2X1_LOC_663/B 0.03fF
C35169 OR2X1_LOC_290/Y AND2X1_LOC_634/a_8_24# 0.24fF
C35170 OR2X1_LOC_160/A OR2X1_LOC_215/Y 0.02fF
C35171 OR2X1_LOC_822/a_8_216# OR2X1_LOC_54/Y 0.01fF
C35172 AND2X1_LOC_633/a_8_24# AND2X1_LOC_573/A 0.01fF
C35173 OR2X1_LOC_844/Y OR2X1_LOC_66/A 0.01fF
C35174 OR2X1_LOC_409/B AND2X1_LOC_774/A 0.25fF
C35175 OR2X1_LOC_405/A OR2X1_LOC_154/A 0.69fF
C35176 AND2X1_LOC_348/A OR2X1_LOC_585/A 0.00fF
C35177 OR2X1_LOC_6/A OR2X1_LOC_393/Y 0.02fF
C35178 OR2X1_LOC_263/a_36_216# AND2X1_LOC_243/Y 0.01fF
C35179 AND2X1_LOC_843/Y OR2X1_LOC_26/Y 0.01fF
C35180 AND2X1_LOC_377/a_8_24# OR2X1_LOC_472/A 0.23fF
C35181 OR2X1_LOC_422/Y OR2X1_LOC_52/B 0.01fF
C35182 OR2X1_LOC_228/Y OR2X1_LOC_776/A 0.01fF
C35183 AND2X1_LOC_344/a_8_24# OR2X1_LOC_485/A 0.01fF
C35184 OR2X1_LOC_161/A OR2X1_LOC_779/a_8_216# 0.03fF
C35185 OR2X1_LOC_620/a_8_216# OR2X1_LOC_620/A 0.47fF
C35186 AND2X1_LOC_459/Y AND2X1_LOC_43/B 0.04fF
C35187 AND2X1_LOC_36/Y AND2X1_LOC_751/a_36_24# 0.00fF
C35188 OR2X1_LOC_553/B OR2X1_LOC_553/a_8_216# 0.03fF
C35189 AND2X1_LOC_95/Y AND2X1_LOC_252/a_8_24# 0.04fF
C35190 AND2X1_LOC_798/A AND2X1_LOC_810/B 0.13fF
C35191 OR2X1_LOC_671/Y OR2X1_LOC_62/A 0.09fF
C35192 OR2X1_LOC_69/Y OR2X1_LOC_39/A 0.06fF
C35193 OR2X1_LOC_47/Y OR2X1_LOC_584/a_8_216# 0.01fF
C35194 AND2X1_LOC_851/a_8_24# AND2X1_LOC_465/Y 0.16fF
C35195 AND2X1_LOC_40/Y OR2X1_LOC_435/Y 0.01fF
C35196 AND2X1_LOC_42/B AND2X1_LOC_618/a_36_24# 0.00fF
C35197 AND2X1_LOC_654/Y OR2X1_LOC_299/Y 0.06fF
C35198 OR2X1_LOC_782/B OR2X1_LOC_87/A 0.01fF
C35199 OR2X1_LOC_462/B OR2X1_LOC_97/B 0.01fF
C35200 OR2X1_LOC_502/A OR2X1_LOC_647/Y 0.03fF
C35201 OR2X1_LOC_36/Y AND2X1_LOC_840/B 0.59fF
C35202 AND2X1_LOC_539/a_8_24# INPUT_0 0.01fF
C35203 AND2X1_LOC_650/Y OR2X1_LOC_6/A 0.44fF
C35204 OR2X1_LOC_417/A AND2X1_LOC_286/a_8_24# 0.01fF
C35205 AND2X1_LOC_42/B OR2X1_LOC_833/B 0.39fF
C35206 OR2X1_LOC_600/A OR2X1_LOC_55/a_8_216# 0.01fF
C35207 OR2X1_LOC_817/a_8_216# AND2X1_LOC_847/Y 0.06fF
C35208 AND2X1_LOC_729/Y AND2X1_LOC_645/A 0.01fF
C35209 OR2X1_LOC_131/Y OR2X1_LOC_18/Y 0.03fF
C35210 OR2X1_LOC_528/Y OR2X1_LOC_615/Y 0.03fF
C35211 OR2X1_LOC_669/Y AND2X1_LOC_859/a_8_24# 0.23fF
C35212 OR2X1_LOC_500/A AND2X1_LOC_3/Y 0.01fF
C35213 OR2X1_LOC_816/A OR2X1_LOC_753/Y 0.21fF
C35214 OR2X1_LOC_405/A OR2X1_LOC_778/A 0.01fF
C35215 AND2X1_LOC_535/Y OR2X1_LOC_47/Y 0.03fF
C35216 OR2X1_LOC_516/Y OR2X1_LOC_437/A 0.07fF
C35217 OR2X1_LOC_690/a_8_216# OR2X1_LOC_690/A 0.01fF
C35218 OR2X1_LOC_185/A OR2X1_LOC_475/Y 0.02fF
C35219 VDD OR2X1_LOC_224/Y 0.18fF
C35220 OR2X1_LOC_108/Y OR2X1_LOC_184/Y 0.00fF
C35221 OR2X1_LOC_306/Y AND2X1_LOC_390/B 0.04fF
C35222 OR2X1_LOC_189/Y AND2X1_LOC_565/Y 0.01fF
C35223 OR2X1_LOC_87/A AND2X1_LOC_19/a_8_24# 0.15fF
C35224 OR2X1_LOC_270/Y AND2X1_LOC_18/Y 0.01fF
C35225 OR2X1_LOC_174/A OR2X1_LOC_434/A 0.28fF
C35226 AND2X1_LOC_675/Y AND2X1_LOC_675/A 0.02fF
C35227 AND2X1_LOC_654/a_8_24# OR2X1_LOC_52/B 0.02fF
C35228 OR2X1_LOC_124/a_8_216# OR2X1_LOC_786/Y 0.01fF
C35229 OR2X1_LOC_235/a_8_216# OR2X1_LOC_74/A 0.01fF
C35230 D_INPUT_5 AND2X1_LOC_25/a_8_24# 0.01fF
C35231 AND2X1_LOC_514/Y AND2X1_LOC_661/a_8_24# -0.01fF
C35232 OR2X1_LOC_158/A OR2X1_LOC_595/Y 0.01fF
C35233 AND2X1_LOC_168/Y AND2X1_LOC_514/Y 0.01fF
C35234 OR2X1_LOC_26/Y OR2X1_LOC_7/A 10.81fF
C35235 OR2X1_LOC_40/Y AND2X1_LOC_804/a_8_24# 0.02fF
C35236 OR2X1_LOC_787/Y OR2X1_LOC_269/B 0.09fF
C35237 OR2X1_LOC_759/A AND2X1_LOC_624/B 0.02fF
C35238 VDD OR2X1_LOC_597/Y 0.12fF
C35239 AND2X1_LOC_40/Y AND2X1_LOC_431/a_8_24# 0.01fF
C35240 OR2X1_LOC_494/Y AND2X1_LOC_721/A 0.57fF
C35241 AND2X1_LOC_54/a_8_24# D_INPUT_2 0.01fF
C35242 OR2X1_LOC_2/Y OR2X1_LOC_429/a_8_216# 0.02fF
C35243 AND2X1_LOC_363/Y AND2X1_LOC_721/A 0.59fF
C35244 OR2X1_LOC_743/A OR2X1_LOC_433/a_36_216# 0.03fF
C35245 OR2X1_LOC_40/Y AND2X1_LOC_202/a_8_24# 0.01fF
C35246 OR2X1_LOC_728/B OR2X1_LOC_596/A 0.01fF
C35247 OR2X1_LOC_476/B OR2X1_LOC_405/Y 0.03fF
C35248 OR2X1_LOC_149/B OR2X1_LOC_546/a_8_216# 0.03fF
C35249 AND2X1_LOC_349/B OR2X1_LOC_7/A 0.01fF
C35250 OR2X1_LOC_89/A OR2X1_LOC_7/A 0.35fF
C35251 AND2X1_LOC_10/a_8_24# OR2X1_LOC_267/A 0.01fF
C35252 OR2X1_LOC_632/Y D_INPUT_1 0.07fF
C35253 AND2X1_LOC_464/Y AND2X1_LOC_464/a_8_24# 0.01fF
C35254 OR2X1_LOC_6/B OR2X1_LOC_398/a_36_216# 0.00fF
C35255 OR2X1_LOC_643/Y OR2X1_LOC_222/A 0.01fF
C35256 OR2X1_LOC_70/Y AND2X1_LOC_336/a_8_24# 0.01fF
C35257 AND2X1_LOC_729/Y AND2X1_LOC_477/A 0.07fF
C35258 AND2X1_LOC_860/A AND2X1_LOC_562/Y 0.10fF
C35259 OR2X1_LOC_139/A OR2X1_LOC_141/a_8_216# 0.03fF
C35260 OR2X1_LOC_744/A OR2X1_LOC_419/Y 0.16fF
C35261 OR2X1_LOC_64/Y AND2X1_LOC_454/A 0.09fF
C35262 OR2X1_LOC_849/A OR2X1_LOC_474/a_8_216# 0.00fF
C35263 OR2X1_LOC_344/A OR2X1_LOC_366/Y 1.17fF
C35264 D_INPUT_3 OR2X1_LOC_278/Y 0.03fF
C35265 OR2X1_LOC_98/A OR2X1_LOC_98/a_8_216# 0.47fF
C35266 OR2X1_LOC_702/A OR2X1_LOC_193/A 0.15fF
C35267 AND2X1_LOC_36/Y OR2X1_LOC_121/A 0.06fF
C35268 OR2X1_LOC_702/A AND2X1_LOC_136/a_36_24# 0.00fF
C35269 AND2X1_LOC_784/A AND2X1_LOC_477/A 0.02fF
C35270 OR2X1_LOC_622/A OR2X1_LOC_80/A 0.10fF
C35271 AND2X1_LOC_211/B AND2X1_LOC_537/Y 0.02fF
C35272 OR2X1_LOC_364/A OR2X1_LOC_544/A 0.03fF
C35273 AND2X1_LOC_558/a_8_24# AND2X1_LOC_657/A 0.03fF
C35274 OR2X1_LOC_669/A OR2X1_LOC_417/A 0.02fF
C35275 AND2X1_LOC_394/a_36_24# AND2X1_LOC_47/Y 0.00fF
C35276 OR2X1_LOC_36/Y OR2X1_LOC_31/Y 4.18fF
C35277 AND2X1_LOC_715/A OR2X1_LOC_521/a_36_216# 0.00fF
C35278 AND2X1_LOC_41/A OR2X1_LOC_641/B 0.03fF
C35279 AND2X1_LOC_592/Y OR2X1_LOC_424/Y 0.89fF
C35280 OR2X1_LOC_656/B OR2X1_LOC_205/Y 0.07fF
C35281 OR2X1_LOC_121/B AND2X1_LOC_67/Y 0.06fF
C35282 OR2X1_LOC_409/B OR2X1_LOC_752/a_8_216# 0.01fF
C35283 OR2X1_LOC_223/A OR2X1_LOC_130/A 0.03fF
C35284 OR2X1_LOC_678/a_8_216# OR2X1_LOC_513/Y 0.40fF
C35285 OR2X1_LOC_678/Y OR2X1_LOC_513/a_8_216# 0.01fF
C35286 AND2X1_LOC_191/Y AND2X1_LOC_630/a_8_24# 0.04fF
C35287 OR2X1_LOC_186/Y OR2X1_LOC_703/Y 0.02fF
C35288 AND2X1_LOC_354/a_8_24# AND2X1_LOC_798/A 0.01fF
C35289 OR2X1_LOC_49/A OR2X1_LOC_622/B 0.01fF
C35290 AND2X1_LOC_727/A AND2X1_LOC_798/Y 0.01fF
C35291 AND2X1_LOC_831/a_36_24# AND2X1_LOC_476/A 0.00fF
C35292 OR2X1_LOC_252/a_36_216# AND2X1_LOC_624/B 0.00fF
C35293 OR2X1_LOC_246/Y OR2X1_LOC_47/Y 0.18fF
C35294 AND2X1_LOC_508/A AND2X1_LOC_657/A 0.01fF
C35295 AND2X1_LOC_810/Y OR2X1_LOC_52/B 0.16fF
C35296 OR2X1_LOC_702/A D_INPUT_0 0.03fF
C35297 AND2X1_LOC_576/Y OR2X1_LOC_47/Y 0.04fF
C35298 OR2X1_LOC_369/Y OR2X1_LOC_437/A -0.03fF
C35299 OR2X1_LOC_291/Y OR2X1_LOC_19/B 0.07fF
C35300 OR2X1_LOC_561/a_8_216# D_INPUT_1 0.01fF
C35301 AND2X1_LOC_753/B OR2X1_LOC_198/A 0.01fF
C35302 OR2X1_LOC_175/Y OR2X1_LOC_139/A 0.12fF
C35303 AND2X1_LOC_34/Y OR2X1_LOC_598/A 0.03fF
C35304 AND2X1_LOC_59/Y OR2X1_LOC_76/a_8_216# 0.06fF
C35305 AND2X1_LOC_64/Y OR2X1_LOC_843/B 0.16fF
C35306 AND2X1_LOC_727/A OR2X1_LOC_46/A 0.02fF
C35307 AND2X1_LOC_126/a_8_24# OR2X1_LOC_71/A 0.01fF
C35308 OR2X1_LOC_726/A OR2X1_LOC_727/a_36_216# 0.00fF
C35309 OR2X1_LOC_164/Y OR2X1_LOC_164/a_8_216# 0.14fF
C35310 AND2X1_LOC_738/B OR2X1_LOC_142/Y 0.02fF
C35311 OR2X1_LOC_476/B D_INPUT_0 0.01fF
C35312 AND2X1_LOC_840/B OR2X1_LOC_419/Y 0.10fF
C35313 OR2X1_LOC_56/A OR2X1_LOC_142/Y 0.04fF
C35314 OR2X1_LOC_160/A OR2X1_LOC_398/Y 0.04fF
C35315 AND2X1_LOC_64/Y OR2X1_LOC_549/A 0.18fF
C35316 AND2X1_LOC_133/a_8_24# OR2X1_LOC_62/B 0.01fF
C35317 OR2X1_LOC_139/A OR2X1_LOC_691/Y 0.01fF
C35318 OR2X1_LOC_196/B AND2X1_LOC_692/a_36_24# 0.00fF
C35319 OR2X1_LOC_650/Y D_INPUT_0 0.09fF
C35320 OR2X1_LOC_18/Y AND2X1_LOC_657/A 0.07fF
C35321 AND2X1_LOC_721/Y AND2X1_LOC_795/a_8_24# 0.01fF
C35322 OR2X1_LOC_45/B AND2X1_LOC_773/Y 0.01fF
C35323 AND2X1_LOC_593/a_36_24# OR2X1_LOC_696/A 0.00fF
C35324 OR2X1_LOC_49/a_8_216# OR2X1_LOC_598/A 0.11fF
C35325 AND2X1_LOC_483/a_8_24# OR2X1_LOC_615/Y -0.00fF
C35326 OR2X1_LOC_89/A OR2X1_LOC_511/a_8_216# 0.01fF
C35327 AND2X1_LOC_44/Y OR2X1_LOC_580/B 0.08fF
C35328 OR2X1_LOC_161/B OR2X1_LOC_578/a_8_216# 0.03fF
C35329 OR2X1_LOC_244/a_8_216# OR2X1_LOC_141/a_8_216# 0.47fF
C35330 VDD OR2X1_LOC_356/B 0.27fF
C35331 OR2X1_LOC_258/a_8_216# AND2X1_LOC_792/Y 0.04fF
C35332 AND2X1_LOC_291/a_8_24# OR2X1_LOC_68/B 0.01fF
C35333 OR2X1_LOC_49/A OR2X1_LOC_9/a_8_216# 0.02fF
C35334 OR2X1_LOC_95/Y OR2X1_LOC_46/A 0.08fF
C35335 OR2X1_LOC_756/B OR2X1_LOC_539/B 0.02fF
C35336 D_INPUT_3 OR2X1_LOC_19/B 0.04fF
C35337 OR2X1_LOC_185/A AND2X1_LOC_406/a_36_24# 0.00fF
C35338 AND2X1_LOC_433/a_8_24# OR2X1_LOC_435/A 0.09fF
C35339 OR2X1_LOC_589/A OR2X1_LOC_428/A 0.12fF
C35340 OR2X1_LOC_368/a_8_216# OR2X1_LOC_368/Y 0.02fF
C35341 AND2X1_LOC_547/Y OR2X1_LOC_406/Y 0.00fF
C35342 AND2X1_LOC_190/a_8_24# AND2X1_LOC_465/A 0.00fF
C35343 OR2X1_LOC_648/B AND2X1_LOC_44/Y 0.03fF
C35344 OR2X1_LOC_589/A OR2X1_LOC_595/A 0.16fF
C35345 OR2X1_LOC_186/Y OR2X1_LOC_596/A 0.02fF
C35346 OR2X1_LOC_357/a_8_216# OR2X1_LOC_182/B 0.01fF
C35347 AND2X1_LOC_802/B AND2X1_LOC_436/Y 0.01fF
C35348 AND2X1_LOC_64/Y OR2X1_LOC_113/Y 0.00fF
C35349 AND2X1_LOC_56/B OR2X1_LOC_181/A 0.02fF
C35350 AND2X1_LOC_227/Y OR2X1_LOC_95/Y 0.08fF
C35351 OR2X1_LOC_62/A OR2X1_LOC_532/B 0.01fF
C35352 OR2X1_LOC_280/Y AND2X1_LOC_563/Y 0.02fF
C35353 AND2X1_LOC_3/Y OR2X1_LOC_789/A 0.03fF
C35354 OR2X1_LOC_51/Y OR2X1_LOC_18/a_8_216# 0.01fF
C35355 AND2X1_LOC_475/Y AND2X1_LOC_476/Y 0.05fF
C35356 OR2X1_LOC_124/A OR2X1_LOC_139/A 0.03fF
C35357 OR2X1_LOC_421/A OR2X1_LOC_693/a_8_216# 0.01fF
C35358 OR2X1_LOC_636/B AND2X1_LOC_31/Y 0.35fF
C35359 AND2X1_LOC_166/a_36_24# OR2X1_LOC_788/B 0.00fF
C35360 OR2X1_LOC_604/A OR2X1_LOC_604/Y 0.21fF
C35361 OR2X1_LOC_426/B AND2X1_LOC_786/Y 0.10fF
C35362 AND2X1_LOC_56/B OR2X1_LOC_550/B 0.03fF
C35363 AND2X1_LOC_64/Y OR2X1_LOC_354/A 0.29fF
C35364 OR2X1_LOC_190/A OR2X1_LOC_294/Y 0.39fF
C35365 OR2X1_LOC_738/A AND2X1_LOC_36/Y 0.25fF
C35366 OR2X1_LOC_161/A OR2X1_LOC_523/a_36_216# 0.00fF
C35367 OR2X1_LOC_297/A OR2X1_LOC_428/A 0.81fF
C35368 AND2X1_LOC_193/Y AND2X1_LOC_200/a_8_24# 0.19fF
C35369 OR2X1_LOC_241/Y OR2X1_LOC_786/Y 0.10fF
C35370 OR2X1_LOC_59/Y OR2X1_LOC_373/Y 0.15fF
C35371 OR2X1_LOC_8/Y OR2X1_LOC_671/Y 0.09fF
C35372 OR2X1_LOC_161/A OR2X1_LOC_319/Y 0.01fF
C35373 AND2X1_LOC_561/a_8_24# AND2X1_LOC_573/A 0.01fF
C35374 OR2X1_LOC_160/B OR2X1_LOC_362/A 0.07fF
C35375 OR2X1_LOC_446/a_8_216# OR2X1_LOC_446/B 0.02fF
C35376 VDD OR2X1_LOC_182/B 0.10fF
C35377 OR2X1_LOC_36/Y OR2X1_LOC_320/a_8_216# 0.03fF
C35378 AND2X1_LOC_866/A AND2X1_LOC_792/Y 0.01fF
C35379 OR2X1_LOC_813/Y OR2X1_LOC_95/Y 0.03fF
C35380 AND2X1_LOC_357/A VDD -0.00fF
C35381 OR2X1_LOC_31/Y OR2X1_LOC_419/Y 0.56fF
C35382 AND2X1_LOC_47/Y AND2X1_LOC_497/a_8_24# 0.02fF
C35383 OR2X1_LOC_22/Y AND2X1_LOC_563/Y 0.09fF
C35384 AND2X1_LOC_40/Y OR2X1_LOC_577/Y 0.03fF
C35385 OR2X1_LOC_39/A OR2X1_LOC_743/Y 0.01fF
C35386 OR2X1_LOC_858/A OR2X1_LOC_349/A 0.05fF
C35387 OR2X1_LOC_199/a_8_216# OR2X1_LOC_502/A 0.00fF
C35388 AND2X1_LOC_95/Y OR2X1_LOC_415/Y 0.89fF
C35389 VDD AND2X1_LOC_731/Y 0.21fF
C35390 AND2X1_LOC_710/Y AND2X1_LOC_347/B 0.03fF
C35391 OR2X1_LOC_287/B OR2X1_LOC_771/B 0.03fF
C35392 AND2X1_LOC_654/B OR2X1_LOC_428/A 2.48fF
C35393 AND2X1_LOC_633/Y AND2X1_LOC_203/a_8_24# 0.17fF
C35394 OR2X1_LOC_158/A AND2X1_LOC_364/Y 0.03fF
C35395 VDD OR2X1_LOC_822/Y 0.14fF
C35396 OR2X1_LOC_234/a_8_216# D_INPUT_1 0.01fF
C35397 AND2X1_LOC_392/A OR2X1_LOC_51/Y 0.00fF
C35398 OR2X1_LOC_106/Y AND2X1_LOC_573/A 0.04fF
C35399 OR2X1_LOC_630/a_8_216# OR2X1_LOC_563/A 0.01fF
C35400 OR2X1_LOC_126/a_36_216# AND2X1_LOC_573/A 0.00fF
C35401 AND2X1_LOC_731/Y AND2X1_LOC_738/a_8_24# 0.09fF
C35402 AND2X1_LOC_40/Y OR2X1_LOC_550/A 0.11fF
C35403 AND2X1_LOC_110/Y AND2X1_LOC_92/Y 0.03fF
C35404 AND2X1_LOC_5/a_8_24# OR2X1_LOC_68/B 0.05fF
C35405 OR2X1_LOC_51/B OR2X1_LOC_31/a_8_216# 0.02fF
C35406 VDD AND2X1_LOC_367/B 0.05fF
C35407 OR2X1_LOC_323/A OR2X1_LOC_91/Y 0.03fF
C35408 OR2X1_LOC_696/A AND2X1_LOC_359/B 0.30fF
C35409 OR2X1_LOC_604/A OR2X1_LOC_744/A 0.18fF
C35410 OR2X1_LOC_485/a_8_216# OR2X1_LOC_12/Y 0.07fF
C35411 OR2X1_LOC_175/B OR2X1_LOC_161/B 0.00fF
C35412 AND2X1_LOC_358/Y AND2X1_LOC_649/B 0.01fF
C35413 OR2X1_LOC_666/a_8_216# OR2X1_LOC_59/Y 0.01fF
C35414 OR2X1_LOC_664/a_8_216# OR2X1_LOC_563/A 0.01fF
C35415 OR2X1_LOC_600/A AND2X1_LOC_663/A 0.03fF
C35416 AND2X1_LOC_218/a_8_24# OR2X1_LOC_91/A 0.06fF
C35417 OR2X1_LOC_91/Y OR2X1_LOC_89/Y 0.01fF
C35418 OR2X1_LOC_676/Y OR2X1_LOC_715/A 0.03fF
C35419 OR2X1_LOC_481/a_8_216# AND2X1_LOC_789/Y 0.01fF
C35420 INPUT_0 AND2X1_LOC_18/Y 0.07fF
C35421 OR2X1_LOC_49/A OR2X1_LOC_394/Y 0.14fF
C35422 AND2X1_LOC_733/Y AND2X1_LOC_784/a_8_24# 0.04fF
C35423 VDD OR2X1_LOC_168/B 0.30fF
C35424 OR2X1_LOC_291/Y AND2X1_LOC_608/a_8_24# 0.26fF
C35425 AND2X1_LOC_22/Y OR2X1_LOC_137/B 0.02fF
C35426 AND2X1_LOC_92/a_8_24# AND2X1_LOC_43/B 0.04fF
C35427 OR2X1_LOC_118/a_8_216# OR2X1_LOC_118/Y 0.01fF
C35428 AND2X1_LOC_658/A AND2X1_LOC_858/B 0.08fF
C35429 OR2X1_LOC_631/B OR2X1_LOC_556/a_36_216# 0.01fF
C35430 AND2X1_LOC_365/A OR2X1_LOC_428/A 3.86fF
C35431 VDD OR2X1_LOC_57/Y 0.12fF
C35432 OR2X1_LOC_187/Y OR2X1_LOC_613/Y 0.02fF
C35433 OR2X1_LOC_379/Y AND2X1_LOC_585/a_8_24# 0.01fF
C35434 OR2X1_LOC_405/A OR2X1_LOC_435/A 0.08fF
C35435 AND2X1_LOC_211/B OR2X1_LOC_171/a_8_216# 0.01fF
C35436 VDD AND2X1_LOC_508/A 0.21fF
C35437 AND2X1_LOC_366/A OR2X1_LOC_51/Y 0.03fF
C35438 OR2X1_LOC_158/A OR2X1_LOC_837/B 0.07fF
C35439 AND2X1_LOC_729/Y AND2X1_LOC_703/Y 0.01fF
C35440 OR2X1_LOC_158/A AND2X1_LOC_76/a_8_24# 0.02fF
C35441 AND2X1_LOC_794/B OR2X1_LOC_48/B 0.07fF
C35442 OR2X1_LOC_323/A OR2X1_LOC_371/a_8_216# 0.01fF
C35443 AND2X1_LOC_510/a_8_24# AND2X1_LOC_508/a_8_24# 0.23fF
C35444 OR2X1_LOC_160/B OR2X1_LOC_474/Y 0.11fF
C35445 OR2X1_LOC_160/A OR2X1_LOC_35/A 0.01fF
C35446 OR2X1_LOC_121/Y OR2X1_LOC_115/a_36_216# 0.01fF
C35447 AND2X1_LOC_64/Y OR2X1_LOC_711/A 0.03fF
C35448 AND2X1_LOC_471/Y AND2X1_LOC_469/B 0.00fF
C35449 OR2X1_LOC_775/a_8_216# AND2X1_LOC_18/Y 0.01fF
C35450 AND2X1_LOC_660/A AND2X1_LOC_216/a_8_24# 0.05fF
C35451 AND2X1_LOC_726/Y OR2X1_LOC_189/Y 0.10fF
C35452 OR2X1_LOC_539/A OR2X1_LOC_160/B 0.01fF
C35453 OR2X1_LOC_36/Y OR2X1_LOC_79/a_8_216# 0.01fF
C35454 AND2X1_LOC_752/a_8_24# VDD -0.00fF
C35455 AND2X1_LOC_319/A AND2X1_LOC_802/Y 0.81fF
C35456 OR2X1_LOC_176/a_8_216# OR2X1_LOC_26/Y 0.07fF
C35457 OR2X1_LOC_496/Y AND2X1_LOC_721/Y 0.03fF
C35458 AND2X1_LOC_726/Y OR2X1_LOC_152/Y 0.00fF
C35459 INPUT_3 OR2X1_LOC_9/Y 0.21fF
C35460 OR2X1_LOC_756/B OR2X1_LOC_78/B 0.81fF
C35461 OR2X1_LOC_175/Y OR2X1_LOC_208/a_8_216# 0.01fF
C35462 AND2X1_LOC_775/a_8_24# OR2X1_LOC_373/Y 0.03fF
C35463 VDD AND2X1_LOC_852/B 0.01fF
C35464 OR2X1_LOC_447/Y OR2X1_LOC_777/B 0.04fF
C35465 OR2X1_LOC_36/Y AND2X1_LOC_213/B 0.00fF
C35466 OR2X1_LOC_43/A OR2X1_LOC_428/A 0.43fF
C35467 OR2X1_LOC_56/A OR2X1_LOC_16/a_8_216# 0.08fF
C35468 OR2X1_LOC_814/A AND2X1_LOC_591/a_8_24# 0.02fF
C35469 OR2X1_LOC_405/A OR2X1_LOC_723/a_8_216# 0.02fF
C35470 AND2X1_LOC_64/Y OR2X1_LOC_629/a_8_216# 0.01fF
C35471 AND2X1_LOC_831/a_8_24# OR2X1_LOC_12/Y 0.04fF
C35472 AND2X1_LOC_733/Y AND2X1_LOC_471/Y 0.02fF
C35473 OR2X1_LOC_158/A AND2X1_LOC_35/a_8_24# 0.05fF
C35474 OR2X1_LOC_296/a_8_216# OR2X1_LOC_563/A 0.01fF
C35475 OR2X1_LOC_12/Y OR2X1_LOC_44/Y 2.86fF
C35476 AND2X1_LOC_707/Y OR2X1_LOC_682/Y 0.14fF
C35477 OR2X1_LOC_106/a_8_216# OR2X1_LOC_67/A 0.01fF
C35478 OR2X1_LOC_659/Y OR2X1_LOC_659/B 0.13fF
C35479 AND2X1_LOC_572/a_8_24# OR2X1_LOC_490/Y -0.00fF
C35480 VDD OR2X1_LOC_48/B 1.05fF
C35481 OR2X1_LOC_157/a_8_216# OR2X1_LOC_158/A 0.01fF
C35482 OR2X1_LOC_33/B OR2X1_LOC_338/A 0.16fF
C35483 OR2X1_LOC_840/a_8_216# OR2X1_LOC_87/A 0.02fF
C35484 OR2X1_LOC_177/Y AND2X1_LOC_840/B 0.05fF
C35485 OR2X1_LOC_168/a_8_216# OR2X1_LOC_66/A 0.01fF
C35486 AND2X1_LOC_357/a_36_24# OR2X1_LOC_426/B 0.01fF
C35487 OR2X1_LOC_43/A OR2X1_LOC_595/A 0.07fF
C35488 OR2X1_LOC_797/B OR2X1_LOC_213/A 0.02fF
C35489 VDD OR2X1_LOC_18/Y 1.26fF
C35490 OR2X1_LOC_789/B AND2X1_LOC_18/Y 0.11fF
C35491 AND2X1_LOC_197/Y AND2X1_LOC_198/a_8_24# 0.01fF
C35492 OR2X1_LOC_89/A OR2X1_LOC_753/a_8_216# 0.01fF
C35493 VDD OR2X1_LOC_739/B 0.37fF
C35494 OR2X1_LOC_9/Y OR2X1_LOC_618/a_36_216# 0.00fF
C35495 AND2X1_LOC_191/a_8_24# AND2X1_LOC_711/Y 0.08fF
C35496 AND2X1_LOC_556/a_8_24# OR2X1_LOC_92/Y 0.09fF
C35497 OR2X1_LOC_97/A OR2X1_LOC_479/Y 0.03fF
C35498 AND2X1_LOC_796/a_36_24# OR2X1_LOC_680/A 0.01fF
C35499 AND2X1_LOC_59/Y VDD 2.79fF
C35500 AND2X1_LOC_658/A AND2X1_LOC_573/A 0.03fF
C35501 OR2X1_LOC_39/A OR2X1_LOC_627/Y 0.00fF
C35502 OR2X1_LOC_743/A AND2X1_LOC_786/Y 0.08fF
C35503 AND2X1_LOC_737/Y OR2X1_LOC_441/a_8_216# 0.01fF
C35504 OR2X1_LOC_744/A AND2X1_LOC_850/a_8_24# 0.02fF
C35505 OR2X1_LOC_118/Y OR2X1_LOC_56/A 0.02fF
C35506 AND2X1_LOC_82/Y OR2X1_LOC_401/Y 0.00fF
C35507 AND2X1_LOC_714/B OR2X1_LOC_52/B 0.07fF
C35508 OR2X1_LOC_496/Y OR2X1_LOC_482/Y 0.00fF
C35509 AND2X1_LOC_566/a_8_24# AND2X1_LOC_566/B 0.04fF
C35510 AND2X1_LOC_624/A AND2X1_LOC_658/Y 0.01fF
C35511 OR2X1_LOC_40/Y OR2X1_LOC_246/a_8_216# 0.14fF
C35512 OR2X1_LOC_348/Y OR2X1_LOC_285/A 0.81fF
C35513 AND2X1_LOC_95/Y OR2X1_LOC_632/Y 0.07fF
C35514 OR2X1_LOC_123/B AND2X1_LOC_44/Y 0.05fF
C35515 OR2X1_LOC_533/Y AND2X1_LOC_390/B 0.01fF
C35516 AND2X1_LOC_570/Y OR2X1_LOC_503/A 0.46fF
C35517 AND2X1_LOC_512/Y AND2X1_LOC_841/B 0.07fF
C35518 AND2X1_LOC_520/Y AND2X1_LOC_222/a_36_24# 0.00fF
C35519 AND2X1_LOC_565/a_8_24# AND2X1_LOC_565/Y 0.01fF
C35520 OR2X1_LOC_91/A AND2X1_LOC_847/Y 0.01fF
C35521 OR2X1_LOC_124/B OR2X1_LOC_203/Y 0.18fF
C35522 OR2X1_LOC_124/a_8_216# OR2X1_LOC_204/Y 0.00fF
C35523 OR2X1_LOC_70/Y OR2X1_LOC_373/Y 0.04fF
C35524 OR2X1_LOC_851/A OR2X1_LOC_840/A 0.17fF
C35525 AND2X1_LOC_719/Y OR2X1_LOC_665/Y 0.00fF
C35526 OR2X1_LOC_40/Y AND2X1_LOC_853/Y 0.09fF
C35527 OR2X1_LOC_6/B OR2X1_LOC_612/B 0.09fF
C35528 AND2X1_LOC_562/B OR2X1_LOC_427/A 0.01fF
C35529 OR2X1_LOC_158/A OR2X1_LOC_73/a_8_216# 0.02fF
C35530 OR2X1_LOC_27/Y AND2X1_LOC_219/A 0.04fF
C35531 OR2X1_LOC_380/A OR2X1_LOC_380/a_8_216# 0.08fF
C35532 AND2X1_LOC_41/A OR2X1_LOC_739/A 0.00fF
C35533 AND2X1_LOC_777/a_8_24# OR2X1_LOC_426/B 0.02fF
C35534 AND2X1_LOC_3/Y OR2X1_LOC_307/A 0.74fF
C35535 AND2X1_LOC_848/a_36_24# OR2X1_LOC_59/Y 0.00fF
C35536 AND2X1_LOC_719/Y OR2X1_LOC_485/A 0.13fF
C35537 AND2X1_LOC_716/Y AND2X1_LOC_364/A -0.03fF
C35538 OR2X1_LOC_502/A OR2X1_LOC_231/A 0.03fF
C35539 OR2X1_LOC_691/A AND2X1_LOC_51/Y 0.00fF
C35540 AND2X1_LOC_583/a_8_24# OR2X1_LOC_639/B 0.03fF
C35541 OR2X1_LOC_849/A OR2X1_LOC_66/A 0.05fF
C35542 AND2X1_LOC_304/a_8_24# OR2X1_LOC_161/A 0.01fF
C35543 AND2X1_LOC_12/Y OR2X1_LOC_334/B 0.00fF
C35544 AND2X1_LOC_208/B OR2X1_LOC_18/Y 0.02fF
C35545 OR2X1_LOC_744/A OR2X1_LOC_80/Y 0.01fF
C35546 OR2X1_LOC_702/A OR2X1_LOC_515/A 0.01fF
C35547 OR2X1_LOC_496/Y OR2X1_LOC_496/a_36_216# 0.00fF
C35548 OR2X1_LOC_748/A OR2X1_LOC_700/a_8_216# 0.01fF
C35549 AND2X1_LOC_378/a_36_24# OR2X1_LOC_39/A 0.00fF
C35550 AND2X1_LOC_734/Y AND2X1_LOC_624/A 0.03fF
C35551 AND2X1_LOC_737/a_8_24# AND2X1_LOC_621/Y 0.02fF
C35552 AND2X1_LOC_56/B AND2X1_LOC_24/a_8_24# 0.05fF
C35553 OR2X1_LOC_756/B OR2X1_LOC_375/A 0.28fF
C35554 OR2X1_LOC_158/A AND2X1_LOC_260/a_8_24# 0.27fF
C35555 OR2X1_LOC_596/Y INPUT_0 0.03fF
C35556 AND2X1_LOC_691/a_8_24# OR2X1_LOC_753/A 0.03fF
C35557 VDD OR2X1_LOC_385/Y 0.17fF
C35558 INPUT_0 AND2X1_LOC_413/a_8_24# 0.01fF
C35559 AND2X1_LOC_825/a_8_24# AND2X1_LOC_44/Y -0.00fF
C35560 OR2X1_LOC_246/A AND2X1_LOC_786/Y 0.10fF
C35561 OR2X1_LOC_697/Y OR2X1_LOC_511/Y 0.06fF
C35562 OR2X1_LOC_40/Y OR2X1_LOC_17/Y 0.01fF
C35563 OR2X1_LOC_763/Y OR2X1_LOC_426/B 0.10fF
C35564 OR2X1_LOC_604/A OR2X1_LOC_282/a_8_216# 0.07fF
C35565 OR2X1_LOC_91/Y AND2X1_LOC_723/Y 0.01fF
C35566 AND2X1_LOC_387/B OR2X1_LOC_676/Y 0.07fF
C35567 AND2X1_LOC_500/Y OR2X1_LOC_239/a_36_216# 0.00fF
C35568 OR2X1_LOC_314/a_36_216# AND2X1_LOC_452/Y 0.00fF
C35569 VDD OR2X1_LOC_688/Y 0.16fF
C35570 OR2X1_LOC_154/A AND2X1_LOC_316/a_8_24# 0.02fF
C35571 OR2X1_LOC_6/B AND2X1_LOC_122/a_36_24# 0.01fF
C35572 OR2X1_LOC_56/A OR2X1_LOC_238/Y 0.12fF
C35573 OR2X1_LOC_432/a_8_216# OR2X1_LOC_432/Y 0.00fF
C35574 AND2X1_LOC_41/A OR2X1_LOC_200/a_8_216# 0.04fF
C35575 AND2X1_LOC_177/a_8_24# OR2X1_LOC_87/A 0.01fF
C35576 OR2X1_LOC_502/A OR2X1_LOC_130/A 0.87fF
C35577 OR2X1_LOC_95/Y AND2X1_LOC_227/a_36_24# 0.00fF
C35578 OR2X1_LOC_811/A OR2X1_LOC_161/A 0.03fF
C35579 AND2X1_LOC_109/a_36_24# OR2X1_LOC_390/B 0.00fF
C35580 AND2X1_LOC_41/A OR2X1_LOC_269/B 0.28fF
C35581 OR2X1_LOC_231/A AND2X1_LOC_230/a_8_24# 0.01fF
C35582 AND2X1_LOC_214/A OR2X1_LOC_52/B 0.00fF
C35583 OR2X1_LOC_810/A OR2X1_LOC_561/Y 0.05fF
C35584 OR2X1_LOC_3/Y OR2X1_LOC_666/A 0.01fF
C35585 OR2X1_LOC_196/B OR2X1_LOC_596/A 0.06fF
C35586 OR2X1_LOC_122/Y OR2X1_LOC_106/A 0.09fF
C35587 OR2X1_LOC_13/B OR2X1_LOC_534/Y 0.03fF
C35588 OR2X1_LOC_315/Y OR2X1_LOC_18/Y 0.53fF
C35589 AND2X1_LOC_370/a_36_24# AND2X1_LOC_866/A 0.01fF
C35590 AND2X1_LOC_721/Y AND2X1_LOC_851/B 0.02fF
C35591 OR2X1_LOC_502/A AND2X1_LOC_7/a_8_24# 0.03fF
C35592 OR2X1_LOC_18/Y OR2X1_LOC_616/Y 0.00fF
C35593 OR2X1_LOC_185/A AND2X1_LOC_43/B 0.03fF
C35594 OR2X1_LOC_619/Y AND2X1_LOC_449/Y 0.05fF
C35595 AND2X1_LOC_170/B AND2X1_LOC_802/Y 0.19fF
C35596 INPUT_5 AND2X1_LOC_17/Y 0.20fF
C35597 OR2X1_LOC_364/A OR2X1_LOC_653/Y 0.23fF
C35598 AND2X1_LOC_863/Y AND2X1_LOC_212/Y 0.13fF
C35599 OR2X1_LOC_228/Y OR2X1_LOC_593/B 0.00fF
C35600 OR2X1_LOC_774/Y OR2X1_LOC_392/A 0.01fF
C35601 OR2X1_LOC_739/B OR2X1_LOC_223/B 0.23fF
C35602 AND2X1_LOC_570/Y OR2X1_LOC_64/Y 0.06fF
C35603 OR2X1_LOC_598/Y OR2X1_LOC_644/a_8_216# 0.00fF
C35604 D_INPUT_0 AND2X1_LOC_262/a_8_24# 0.02fF
C35605 OR2X1_LOC_774/Y OR2X1_LOC_489/a_36_216# 0.00fF
C35606 OR2X1_LOC_331/A OR2X1_LOC_64/Y 0.03fF
C35607 OR2X1_LOC_177/Y OR2X1_LOC_31/Y 0.00fF
C35608 OR2X1_LOC_130/A AND2X1_LOC_230/a_8_24# 0.14fF
C35609 AND2X1_LOC_47/Y OR2X1_LOC_486/Y 0.03fF
C35610 OR2X1_LOC_446/B OR2X1_LOC_515/a_8_216# 0.01fF
C35611 AND2X1_LOC_59/a_8_24# AND2X1_LOC_25/Y 0.13fF
C35612 OR2X1_LOC_502/A AND2X1_LOC_612/a_8_24# 0.01fF
C35613 OR2X1_LOC_315/a_8_216# OR2X1_LOC_31/Y 0.07fF
C35614 OR2X1_LOC_316/Y OR2X1_LOC_265/Y 0.03fF
C35615 OR2X1_LOC_277/a_8_216# OR2X1_LOC_59/Y 0.14fF
C35616 OR2X1_LOC_757/A AND2X1_LOC_663/B 0.00fF
C35617 OR2X1_LOC_837/Y OR2X1_LOC_20/a_8_216# 0.01fF
C35618 AND2X1_LOC_430/B AND2X1_LOC_581/a_8_24# 0.01fF
C35619 OR2X1_LOC_335/A OR2X1_LOC_590/a_8_216# 0.01fF
C35620 OR2X1_LOC_468/Y OR2X1_LOC_212/A 0.57fF
C35621 AND2X1_LOC_12/Y OR2X1_LOC_866/a_8_216# 0.00fF
C35622 OR2X1_LOC_774/B OR2X1_LOC_773/Y 0.08fF
C35623 AND2X1_LOC_352/a_8_24# AND2X1_LOC_863/Y 0.02fF
C35624 OR2X1_LOC_678/Y AND2X1_LOC_51/Y 0.05fF
C35625 AND2X1_LOC_716/Y OR2X1_LOC_3/Y 0.07fF
C35626 OR2X1_LOC_47/Y OR2X1_LOC_16/A 0.28fF
C35627 INPUT_3 AND2X1_LOC_852/Y 0.09fF
C35628 OR2X1_LOC_465/a_36_216# OR2X1_LOC_375/A 0.02fF
C35629 OR2X1_LOC_335/a_8_216# OR2X1_LOC_318/B 0.00fF
C35630 OR2X1_LOC_251/Y OR2X1_LOC_18/Y 0.02fF
C35631 OR2X1_LOC_70/Y OR2X1_LOC_426/A 1.53fF
C35632 OR2X1_LOC_604/A OR2X1_LOC_31/Y 0.08fF
C35633 OR2X1_LOC_154/A OR2X1_LOC_673/Y 0.01fF
C35634 OR2X1_LOC_3/Y AND2X1_LOC_654/Y 0.07fF
C35635 AND2X1_LOC_658/A AND2X1_LOC_678/a_36_24# 0.01fF
C35636 AND2X1_LOC_273/a_8_24# OR2X1_LOC_228/Y 0.01fF
C35637 OR2X1_LOC_847/a_8_216# OR2X1_LOC_847/B 0.47fF
C35638 OR2X1_LOC_287/B OR2X1_LOC_402/Y 0.04fF
C35639 AND2X1_LOC_539/Y OR2X1_LOC_761/a_36_216# 0.00fF
C35640 OR2X1_LOC_784/a_8_216# OR2X1_LOC_161/A 0.03fF
C35641 AND2X1_LOC_326/B OR2X1_LOC_111/Y 0.01fF
C35642 OR2X1_LOC_85/A OR2X1_LOC_69/Y 0.01fF
C35643 AND2X1_LOC_147/Y OR2X1_LOC_679/B 0.34fF
C35644 AND2X1_LOC_662/B AND2X1_LOC_276/Y 0.21fF
C35645 AND2X1_LOC_722/A AND2X1_LOC_727/A 0.03fF
C35646 OR2X1_LOC_440/A OR2X1_LOC_66/A 0.03fF
C35647 OR2X1_LOC_81/Y OR2X1_LOC_81/a_8_216# 0.01fF
C35648 AND2X1_LOC_66/a_8_24# AND2X1_LOC_474/A 0.01fF
C35649 OR2X1_LOC_821/Y OR2X1_LOC_813/Y 0.74fF
C35650 OR2X1_LOC_805/A OR2X1_LOC_793/B 0.74fF
C35651 OR2X1_LOC_235/B INPUT_1 0.07fF
C35652 AND2X1_LOC_40/Y OR2X1_LOC_476/B 0.02fF
C35653 OR2X1_LOC_76/A OR2X1_LOC_808/a_8_216# 0.03fF
C35654 OR2X1_LOC_485/A AND2X1_LOC_655/A 0.02fF
C35655 OR2X1_LOC_619/Y AND2X1_LOC_212/B 0.04fF
C35656 OR2X1_LOC_599/A OR2X1_LOC_591/a_8_216# 0.03fF
C35657 OR2X1_LOC_108/Y OR2X1_LOC_47/Y 0.02fF
C35658 OR2X1_LOC_686/B AND2X1_LOC_684/a_36_24# 0.01fF
C35659 OR2X1_LOC_76/A OR2X1_LOC_733/a_8_216# 0.02fF
C35660 OR2X1_LOC_26/Y AND2X1_LOC_836/a_8_24# 0.01fF
C35661 OR2X1_LOC_431/a_36_216# OR2X1_LOC_48/B 0.00fF
C35662 OR2X1_LOC_70/A INPUT_7 0.58fF
C35663 AND2X1_LOC_95/Y OR2X1_LOC_285/B 0.26fF
C35664 OR2X1_LOC_236/a_8_216# OR2X1_LOC_89/A 0.01fF
C35665 OR2X1_LOC_548/A OR2X1_LOC_598/A 0.01fF
C35666 OR2X1_LOC_502/A OR2X1_LOC_62/B 0.04fF
C35667 AND2X1_LOC_120/a_8_24# OR2X1_LOC_39/A 0.11fF
C35668 VDD OR2X1_LOC_549/Y 0.23fF
C35669 OR2X1_LOC_107/Y OR2X1_LOC_95/Y 0.05fF
C35670 OR2X1_LOC_6/B OR2X1_LOC_66/a_8_216# 0.04fF
C35671 OR2X1_LOC_40/Y AND2X1_LOC_792/Y 0.30fF
C35672 OR2X1_LOC_97/A OR2X1_LOC_68/B 1.78fF
C35673 AND2X1_LOC_853/Y AND2X1_LOC_857/a_8_24# 0.05fF
C35674 AND2X1_LOC_520/Y OR2X1_LOC_416/Y 0.04fF
C35675 VDD AND2X1_LOC_620/Y 0.10fF
C35676 OR2X1_LOC_850/B AND2X1_LOC_283/a_8_24# 0.01fF
C35677 OR2X1_LOC_70/Y INPUT_4 0.01fF
C35678 AND2X1_LOC_777/a_8_24# OR2X1_LOC_743/A 0.07fF
C35679 OR2X1_LOC_3/Y GATE_366 0.03fF
C35680 AND2X1_LOC_500/a_8_24# OR2X1_LOC_485/A 0.02fF
C35681 OR2X1_LOC_404/a_8_216# AND2X1_LOC_51/Y 0.01fF
C35682 INPUT_0 AND2X1_LOC_672/a_8_24# 0.03fF
C35683 OR2X1_LOC_11/a_36_216# INPUT_7 0.00fF
C35684 OR2X1_LOC_604/A OR2X1_LOC_257/Y 0.06fF
C35685 AND2X1_LOC_722/A OR2X1_LOC_95/Y 0.13fF
C35686 OR2X1_LOC_384/a_8_216# OR2X1_LOC_428/A 0.01fF
C35687 OR2X1_LOC_714/a_8_216# OR2X1_LOC_308/Y 0.03fF
C35688 OR2X1_LOC_22/Y OR2X1_LOC_433/Y 0.02fF
C35689 OR2X1_LOC_70/Y AND2X1_LOC_100/a_8_24# 0.02fF
C35690 AND2X1_LOC_303/A AND2X1_LOC_350/Y 0.05fF
C35691 VDD AND2X1_LOC_215/A 0.06fF
C35692 AND2X1_LOC_48/A OR2X1_LOC_340/Y 0.03fF
C35693 AND2X1_LOC_157/a_8_24# AND2X1_LOC_425/Y 0.19fF
C35694 OR2X1_LOC_623/a_8_216# D_INPUT_0 0.02fF
C35695 OR2X1_LOC_385/Y AND2X1_LOC_389/a_8_24# 0.01fF
C35696 OR2X1_LOC_837/A AND2X1_LOC_462/Y 0.24fF
C35697 AND2X1_LOC_711/A AND2X1_LOC_848/A 0.01fF
C35698 AND2X1_LOC_135/a_8_24# OR2X1_LOC_269/B 0.05fF
C35699 OR2X1_LOC_168/Y OR2X1_LOC_180/B 0.03fF
C35700 AND2X1_LOC_48/A OR2X1_LOC_130/A 0.03fF
C35701 OR2X1_LOC_36/Y AND2X1_LOC_308/a_8_24# 0.01fF
C35702 AND2X1_LOC_41/a_8_24# OR2X1_LOC_228/Y 0.23fF
C35703 OR2X1_LOC_417/Y OR2X1_LOC_601/Y 0.03fF
C35704 OR2X1_LOC_80/a_36_216# OR2X1_LOC_393/Y 0.00fF
C35705 AND2X1_LOC_831/Y AND2X1_LOC_662/B 0.49fF
C35706 OR2X1_LOC_216/A OR2X1_LOC_786/Y 0.14fF
C35707 OR2X1_LOC_161/B OR2X1_LOC_366/Y 0.14fF
C35708 OR2X1_LOC_502/A AND2X1_LOC_88/Y 0.02fF
C35709 OR2X1_LOC_272/Y AND2X1_LOC_116/Y 0.00fF
C35710 AND2X1_LOC_777/a_8_24# OR2X1_LOC_246/A 0.10fF
C35711 OR2X1_LOC_643/A OR2X1_LOC_474/a_8_216# 0.01fF
C35712 OR2X1_LOC_19/B OR2X1_LOC_83/A 0.07fF
C35713 OR2X1_LOC_17/Y OR2X1_LOC_44/a_8_216# 0.08fF
C35714 OR2X1_LOC_479/Y OR2X1_LOC_605/a_8_216# 0.04fF
C35715 AND2X1_LOC_727/A AND2X1_LOC_854/a_8_24# 0.01fF
C35716 OR2X1_LOC_426/B OR2X1_LOC_88/a_8_216# 0.54fF
C35717 OR2X1_LOC_643/A OR2X1_LOC_859/A 0.01fF
C35718 AND2X1_LOC_34/Y AND2X1_LOC_462/Y 0.89fF
C35719 OR2X1_LOC_3/Y AND2X1_LOC_307/a_8_24# 0.03fF
C35720 OR2X1_LOC_275/a_8_216# OR2X1_LOC_74/A 0.07fF
C35721 AND2X1_LOC_168/Y OR2X1_LOC_47/Y 0.03fF
C35722 OR2X1_LOC_137/Y OR2X1_LOC_62/B 0.02fF
C35723 AND2X1_LOC_710/a_8_24# AND2X1_LOC_866/A 0.02fF
C35724 OR2X1_LOC_473/Y OR2X1_LOC_201/Y 0.01fF
C35725 AND2X1_LOC_477/A OR2X1_LOC_52/B 0.07fF
C35726 OR2X1_LOC_80/Y OR2X1_LOC_31/Y 0.00fF
C35727 OR2X1_LOC_635/A OR2X1_LOC_451/B 0.28fF
C35728 AND2X1_LOC_655/a_8_24# AND2X1_LOC_655/A 0.27fF
C35729 AND2X1_LOC_388/Y OR2X1_LOC_13/B 0.10fF
C35730 OR2X1_LOC_36/Y AND2X1_LOC_270/a_8_24# 0.15fF
C35731 OR2X1_LOC_502/A OR2X1_LOC_365/B 0.01fF
C35732 AND2X1_LOC_59/Y OR2X1_LOC_845/A 0.04fF
C35733 OR2X1_LOC_599/A OR2X1_LOC_95/Y 0.01fF
C35734 OR2X1_LOC_78/A OR2X1_LOC_80/A 0.10fF
C35735 OR2X1_LOC_620/B OR2X1_LOC_471/Y 0.02fF
C35736 OR2X1_LOC_426/A OR2X1_LOC_70/A 0.26fF
C35737 OR2X1_LOC_18/Y AND2X1_LOC_624/B 0.23fF
C35738 OR2X1_LOC_18/Y OR2X1_LOC_67/Y 0.05fF
C35739 OR2X1_LOC_337/a_8_216# OR2X1_LOC_578/B 0.00fF
C35740 AND2X1_LOC_84/Y AND2X1_LOC_201/Y 0.01fF
C35741 OR2X1_LOC_763/Y OR2X1_LOC_409/B 0.00fF
C35742 AND2X1_LOC_476/Y OR2X1_LOC_268/Y 0.01fF
C35743 AND2X1_LOC_367/a_36_24# OR2X1_LOC_47/Y 0.00fF
C35744 AND2X1_LOC_31/Y OR2X1_LOC_712/a_8_216# 0.01fF
C35745 OR2X1_LOC_71/a_8_216# AND2X1_LOC_647/Y 0.01fF
C35746 OR2X1_LOC_403/a_36_216# AND2X1_LOC_51/Y 0.00fF
C35747 OR2X1_LOC_377/A AND2X1_LOC_699/a_8_24# 0.09fF
C35748 OR2X1_LOC_475/B OR2X1_LOC_68/B 0.03fF
C35749 AND2X1_LOC_95/Y OR2X1_LOC_358/A 0.23fF
C35750 VDD OR2X1_LOC_342/B 0.00fF
C35751 OR2X1_LOC_813/A OR2X1_LOC_64/Y 0.03fF
C35752 OR2X1_LOC_89/A OR2X1_LOC_615/Y 0.71fF
C35753 AND2X1_LOC_287/a_8_24# AND2X1_LOC_562/Y 0.25fF
C35754 AND2X1_LOC_290/a_8_24# OR2X1_LOC_68/B 0.01fF
C35755 OR2X1_LOC_115/a_8_216# OR2X1_LOC_560/A 0.01fF
C35756 INPUT_4 OR2X1_LOC_70/A 0.33fF
C35757 OR2X1_LOC_655/B OR2X1_LOC_643/Y 0.00fF
C35758 OR2X1_LOC_687/B OR2X1_LOC_451/B 0.01fF
C35759 OR2X1_LOC_346/B AND2X1_LOC_72/B 0.01fF
C35760 OR2X1_LOC_473/Y OR2X1_LOC_201/a_8_216# 0.01fF
C35761 AND2X1_LOC_2/Y INPUT_6 0.20fF
C35762 OR2X1_LOC_789/B OR2X1_LOC_789/A 0.17fF
C35763 AND2X1_LOC_644/a_8_24# OR2X1_LOC_585/A 0.01fF
C35764 VDD AND2X1_LOC_582/B 0.02fF
C35765 OR2X1_LOC_507/A OR2X1_LOC_510/a_36_216# 0.00fF
C35766 OR2X1_LOC_45/B OR2X1_LOC_12/Y 0.24fF
C35767 OR2X1_LOC_508/a_36_216# OR2X1_LOC_392/B 0.13fF
C35768 OR2X1_LOC_691/Y OR2X1_LOC_138/A 0.00fF
C35769 OR2X1_LOC_440/a_36_216# OR2X1_LOC_168/Y 0.00fF
C35770 AND2X1_LOC_348/A OR2X1_LOC_437/A 0.01fF
C35771 OR2X1_LOC_485/A OR2X1_LOC_599/Y 0.01fF
C35772 OR2X1_LOC_243/B OR2X1_LOC_244/A 0.07fF
C35773 AND2X1_LOC_3/Y AND2X1_LOC_428/a_8_24# 0.10fF
C35774 OR2X1_LOC_633/a_8_216# AND2X1_LOC_36/Y 0.01fF
C35775 OR2X1_LOC_185/A OR2X1_LOC_367/B 0.03fF
C35776 OR2X1_LOC_254/B OR2X1_LOC_578/B 0.01fF
C35777 AND2X1_LOC_620/Y AND2X1_LOC_624/a_8_24# 0.00fF
C35778 OR2X1_LOC_420/Y OR2X1_LOC_419/Y 0.22fF
C35779 OR2X1_LOC_177/Y AND2X1_LOC_464/A 0.01fF
C35780 AND2X1_LOC_364/A OR2X1_LOC_13/B 0.07fF
C35781 OR2X1_LOC_429/Y OR2X1_LOC_581/a_36_216# 0.01fF
C35782 OR2X1_LOC_121/B OR2X1_LOC_223/A 1.29fF
C35783 AND2X1_LOC_710/a_36_24# OR2X1_LOC_59/Y 0.00fF
C35784 OR2X1_LOC_296/Y OR2X1_LOC_247/Y 0.59fF
C35785 AND2X1_LOC_656/Y OR2X1_LOC_71/Y 0.06fF
C35786 OR2X1_LOC_188/Y OR2X1_LOC_733/A 0.70fF
C35787 AND2X1_LOC_804/A AND2X1_LOC_784/a_8_24# 0.10fF
C35788 OR2X1_LOC_62/B OR2X1_LOC_618/Y 0.81fF
C35789 OR2X1_LOC_12/Y OR2X1_LOC_382/A 0.54fF
C35790 OR2X1_LOC_40/Y OR2X1_LOC_816/A 0.02fF
C35791 OR2X1_LOC_671/Y OR2X1_LOC_9/a_8_216# 0.01fF
C35792 AND2X1_LOC_7/B AND2X1_LOC_18/Y 0.37fF
C35793 AND2X1_LOC_51/A AND2X1_LOC_31/Y 0.09fF
C35794 OR2X1_LOC_276/A D_INPUT_0 0.05fF
C35795 AND2X1_LOC_370/a_36_24# OR2X1_LOC_40/Y 0.00fF
C35796 OR2X1_LOC_78/A OR2X1_LOC_115/B 0.12fF
C35797 VDD OR2X1_LOC_764/a_8_216# 0.00fF
C35798 OR2X1_LOC_507/a_8_216# OR2X1_LOC_508/Y 0.01fF
C35799 OR2X1_LOC_786/A OR2X1_LOC_161/B 0.03fF
C35800 AND2X1_LOC_86/Y OR2X1_LOC_771/B 0.07fF
C35801 OR2X1_LOC_151/A AND2X1_LOC_295/a_8_24# 0.01fF
C35802 OR2X1_LOC_624/A OR2X1_LOC_332/a_8_216# 0.06fF
C35803 OR2X1_LOC_47/Y AND2X1_LOC_687/Y 0.02fF
C35804 AND2X1_LOC_573/Y AND2X1_LOC_735/Y 0.91fF
C35805 OR2X1_LOC_604/A AND2X1_LOC_464/A 0.03fF
C35806 OR2X1_LOC_161/A OR2X1_LOC_777/B 0.09fF
C35807 OR2X1_LOC_604/A AND2X1_LOC_213/B 0.03fF
C35808 OR2X1_LOC_721/a_8_216# OR2X1_LOC_66/A 0.01fF
C35809 OR2X1_LOC_326/B OR2X1_LOC_308/Y 0.03fF
C35810 AND2X1_LOC_866/A OR2X1_LOC_95/Y 0.06fF
C35811 OR2X1_LOC_865/B OR2X1_LOC_579/A 0.16fF
C35812 AND2X1_LOC_866/A OR2X1_LOC_368/A 0.03fF
C35813 AND2X1_LOC_547/Y AND2X1_LOC_547/a_8_24# 0.01fF
C35814 AND2X1_LOC_410/a_8_24# OR2X1_LOC_12/Y 0.02fF
C35815 AND2X1_LOC_340/Y VDD 0.09fF
C35816 AND2X1_LOC_64/Y OR2X1_LOC_499/B 0.00fF
C35817 AND2X1_LOC_586/a_8_24# AND2X1_LOC_36/Y 0.02fF
C35818 OR2X1_LOC_684/a_8_216# OR2X1_LOC_12/Y 0.01fF
C35819 AND2X1_LOC_56/B OR2X1_LOC_515/a_8_216# 0.01fF
C35820 OR2X1_LOC_510/Y OR2X1_LOC_217/A 0.14fF
C35821 VDD AND2X1_LOC_810/B 0.21fF
C35822 AND2X1_LOC_705/a_8_24# OR2X1_LOC_12/Y -0.04fF
C35823 AND2X1_LOC_753/B AND2X1_LOC_763/B 0.02fF
C35824 AND2X1_LOC_713/Y OR2X1_LOC_421/Y 0.04fF
C35825 OR2X1_LOC_40/Y AND2X1_LOC_212/A 0.01fF
C35826 OR2X1_LOC_158/A AND2X1_LOC_243/Y 0.07fF
C35827 OR2X1_LOC_847/A AND2X1_LOC_619/a_8_24# 0.01fF
C35828 OR2X1_LOC_176/Y OR2X1_LOC_744/A 0.50fF
C35829 AND2X1_LOC_22/Y OR2X1_LOC_632/Y 0.12fF
C35830 OR2X1_LOC_738/A OR2X1_LOC_469/B 0.01fF
C35831 OR2X1_LOC_91/Y OR2X1_LOC_142/Y 0.03fF
C35832 OR2X1_LOC_106/a_36_216# AND2X1_LOC_243/Y 0.01fF
C35833 OR2X1_LOC_59/Y OR2X1_LOC_759/a_8_216# 0.09fF
C35834 OR2X1_LOC_154/A OR2X1_LOC_723/B 0.07fF
C35835 AND2X1_LOC_181/Y VDD 0.21fF
C35836 OR2X1_LOC_494/A OR2X1_LOC_256/Y 0.00fF
C35837 GATE_811 AND2X1_LOC_796/Y 0.09fF
C35838 OR2X1_LOC_87/A OR2X1_LOC_182/a_8_216# 0.01fF
C35839 OR2X1_LOC_274/Y OR2X1_LOC_121/A 0.01fF
C35840 OR2X1_LOC_808/a_8_216# OR2X1_LOC_722/B 0.40fF
C35841 OR2X1_LOC_62/B OR2X1_LOC_398/a_8_216# 0.01fF
C35842 AND2X1_LOC_70/Y OR2X1_LOC_151/A 0.45fF
C35843 OR2X1_LOC_70/Y OR2X1_LOC_533/a_36_216# 0.00fF
C35844 OR2X1_LOC_621/A AND2X1_LOC_616/a_8_24# 0.21fF
C35845 OR2X1_LOC_473/a_8_216# AND2X1_LOC_7/B 0.03fF
C35846 OR2X1_LOC_19/B AND2X1_LOC_751/a_8_24# 0.01fF
C35847 OR2X1_LOC_485/Y OR2X1_LOC_526/Y 0.42fF
C35848 OR2X1_LOC_505/Y AND2X1_LOC_806/a_8_24# 0.24fF
C35849 AND2X1_LOC_91/B AND2X1_LOC_314/a_8_24# 0.03fF
C35850 OR2X1_LOC_756/B OR2X1_LOC_843/B 0.04fF
C35851 OR2X1_LOC_3/Y OR2X1_LOC_13/B 0.10fF
C35852 VDD OR2X1_LOC_686/a_8_216# 0.21fF
C35853 OR2X1_LOC_45/B OR2X1_LOC_422/a_8_216# 0.01fF
C35854 AND2X1_LOC_806/A OR2X1_LOC_504/a_8_216# 0.01fF
C35855 OR2X1_LOC_779/Y OR2X1_LOC_783/a_8_216# 0.02fF
C35856 OR2X1_LOC_205/Y OR2X1_LOC_786/Y 0.14fF
C35857 OR2X1_LOC_756/B OR2X1_LOC_549/A 0.00fF
C35858 OR2X1_LOC_674/a_8_216# OR2X1_LOC_482/Y 0.03fF
C35859 OR2X1_LOC_643/A OR2X1_LOC_508/Y 0.09fF
C35860 AND2X1_LOC_539/a_36_24# AND2X1_LOC_434/Y 0.01fF
C35861 OR2X1_LOC_770/Y D_INPUT_1 0.02fF
C35862 OR2X1_LOC_335/A OR2X1_LOC_154/A 0.01fF
C35863 AND2X1_LOC_620/Y AND2X1_LOC_624/B 0.05fF
C35864 AND2X1_LOC_787/a_36_24# AND2X1_LOC_787/A 0.01fF
C35865 OR2X1_LOC_160/B OR2X1_LOC_678/a_8_216# 0.03fF
C35866 AND2X1_LOC_51/Y OR2X1_LOC_777/B 0.05fF
C35867 OR2X1_LOC_416/Y OR2X1_LOC_300/a_36_216# 0.00fF
C35868 AND2X1_LOC_322/a_8_24# OR2X1_LOC_703/A 0.01fF
C35869 AND2X1_LOC_860/a_8_24# AND2X1_LOC_860/A 0.08fF
C35870 AND2X1_LOC_190/a_8_24# AND2X1_LOC_858/B 0.03fF
C35871 OR2X1_LOC_527/Y OR2X1_LOC_142/Y 0.07fF
C35872 AND2X1_LOC_81/B OR2X1_LOC_392/B 0.03fF
C35873 OR2X1_LOC_264/Y OR2X1_LOC_509/a_8_216# 0.02fF
C35874 OR2X1_LOC_9/Y AND2X1_LOC_839/a_8_24# 0.01fF
C35875 OR2X1_LOC_624/A OR2X1_LOC_161/B 0.03fF
C35876 AND2X1_LOC_141/a_8_24# OR2X1_LOC_744/A 0.01fF
C35877 AND2X1_LOC_785/A OR2X1_LOC_371/Y 0.20fF
C35878 OR2X1_LOC_528/Y AND2X1_LOC_866/B 0.60fF
C35879 AND2X1_LOC_713/a_8_24# OR2X1_LOC_48/B 0.02fF
C35880 OR2X1_LOC_409/B OR2X1_LOC_378/A 0.00fF
C35881 OR2X1_LOC_421/A OR2X1_LOC_692/a_8_216# 0.01fF
C35882 OR2X1_LOC_49/A OR2X1_LOC_39/A 0.01fF
C35883 OR2X1_LOC_516/B OR2X1_LOC_600/A 0.00fF
C35884 AND2X1_LOC_51/Y D_INPUT_6 0.37fF
C35885 OR2X1_LOC_66/a_8_216# OR2X1_LOC_598/A 0.02fF
C35886 AND2X1_LOC_191/B OR2X1_LOC_755/a_36_216# 0.00fF
C35887 OR2X1_LOC_421/A OR2X1_LOC_92/Y 0.07fF
C35888 VDD OR2X1_LOC_165/Y 0.04fF
C35889 OR2X1_LOC_177/a_8_216# AND2X1_LOC_807/Y 0.14fF
C35890 AND2X1_LOC_721/Y OR2X1_LOC_372/Y 0.00fF
C35891 OR2X1_LOC_447/Y OR2X1_LOC_704/a_36_216# 0.00fF
C35892 OR2X1_LOC_160/A OR2X1_LOC_857/B 0.03fF
C35893 VDD OR2X1_LOC_623/B 0.64fF
C35894 OR2X1_LOC_744/a_36_216# OR2X1_LOC_44/Y 0.03fF
C35895 OR2X1_LOC_45/B AND2X1_LOC_650/Y 0.05fF
C35896 OR2X1_LOC_468/A OR2X1_LOC_502/A 0.03fF
C35897 OR2X1_LOC_318/Y AND2X1_LOC_18/Y 0.07fF
C35898 OR2X1_LOC_166/Y AND2X1_LOC_512/Y 0.02fF
C35899 AND2X1_LOC_766/a_8_24# OR2X1_LOC_287/B 0.01fF
C35900 AND2X1_LOC_181/Y OR2X1_LOC_315/Y 1.82fF
C35901 AND2X1_LOC_335/a_36_24# OR2X1_LOC_426/B 0.00fF
C35902 OR2X1_LOC_45/Y OR2X1_LOC_40/Y 0.07fF
C35903 OR2X1_LOC_653/A OR2X1_LOC_435/A 0.25fF
C35904 OR2X1_LOC_89/A AND2X1_LOC_242/B 0.09fF
C35905 OR2X1_LOC_840/A OR2X1_LOC_78/A 0.10fF
C35906 VDD OR2X1_LOC_794/A 0.18fF
C35907 OR2X1_LOC_135/Y OR2X1_LOC_6/A 0.01fF
C35908 OR2X1_LOC_339/a_8_216# OR2X1_LOC_61/Y 0.05fF
C35909 AND2X1_LOC_40/Y AND2X1_LOC_437/a_8_24# 0.01fF
C35910 AND2X1_LOC_70/Y OR2X1_LOC_788/a_8_216# 0.06fF
C35911 AND2X1_LOC_80/a_8_24# OR2X1_LOC_646/B 0.01fF
C35912 AND2X1_LOC_840/B AND2X1_LOC_212/Y 0.10fF
C35913 AND2X1_LOC_351/a_8_24# OR2X1_LOC_26/Y 0.02fF
C35914 OR2X1_LOC_244/A OR2X1_LOC_771/B 0.07fF
C35915 OR2X1_LOC_804/a_8_216# OR2X1_LOC_808/A 0.12fF
C35916 OR2X1_LOC_535/A OR2X1_LOC_468/Y 0.00fF
C35917 OR2X1_LOC_7/A OR2X1_LOC_816/A 0.80fF
C35918 AND2X1_LOC_716/Y OR2X1_LOC_329/B 0.12fF
C35919 OR2X1_LOC_702/A OR2X1_LOC_138/a_8_216# 0.09fF
C35920 OR2X1_LOC_40/Y AND2X1_LOC_807/Y 0.63fF
C35921 OR2X1_LOC_160/B OR2X1_LOC_402/Y 0.01fF
C35922 AND2X1_LOC_371/a_8_24# OR2X1_LOC_805/A 0.03fF
C35923 OR2X1_LOC_254/a_8_216# OR2X1_LOC_562/A 0.01fF
C35924 AND2X1_LOC_51/Y OR2X1_LOC_831/B 0.08fF
C35925 OR2X1_LOC_76/Y OR2X1_LOC_549/A 0.02fF
C35926 AND2X1_LOC_12/Y OR2X1_LOC_676/Y 0.08fF
C35927 OR2X1_LOC_805/A AND2X1_LOC_18/Y 0.10fF
C35928 OR2X1_LOC_116/a_8_216# OR2X1_LOC_151/A 0.05fF
C35929 OR2X1_LOC_329/B AND2X1_LOC_654/Y 0.07fF
C35930 OR2X1_LOC_135/Y OR2X1_LOC_299/a_8_216# 0.28fF
C35931 OR2X1_LOC_555/A OR2X1_LOC_161/B 0.05fF
C35932 OR2X1_LOC_124/B OR2X1_LOC_375/A 0.01fF
C35933 AND2X1_LOC_456/B OR2X1_LOC_92/Y 0.00fF
C35934 AND2X1_LOC_729/Y OR2X1_LOC_679/a_36_216# 0.01fF
C35935 AND2X1_LOC_728/Y OR2X1_LOC_679/Y 0.21fF
C35936 VDD AND2X1_LOC_228/Y -0.00fF
C35937 OR2X1_LOC_448/Y OR2X1_LOC_466/A 0.03fF
C35938 OR2X1_LOC_375/A OR2X1_LOC_370/a_8_216# 0.01fF
C35939 AND2X1_LOC_99/a_8_24# AND2X1_LOC_99/Y 0.02fF
C35940 AND2X1_LOC_91/B AND2X1_LOC_816/a_8_24# 0.02fF
C35941 OR2X1_LOC_109/Y OR2X1_LOC_59/Y 0.03fF
C35942 AND2X1_LOC_711/Y OR2X1_LOC_759/a_8_216# 0.01fF
C35943 AND2X1_LOC_119/a_8_24# AND2X1_LOC_416/a_8_24# 0.23fF
C35944 OR2X1_LOC_9/Y AND2X1_LOC_839/B 0.05fF
C35945 AND2X1_LOC_390/B AND2X1_LOC_809/a_8_24# 0.01fF
C35946 VDD AND2X1_LOC_192/Y 0.35fF
C35947 AND2X1_LOC_474/Y AND2X1_LOC_475/Y 0.00fF
C35948 AND2X1_LOC_12/Y OR2X1_LOC_834/A 0.63fF
C35949 OR2X1_LOC_304/a_8_216# OR2X1_LOC_431/Y 0.03fF
C35950 AND2X1_LOC_98/a_8_24# OR2X1_LOC_6/A 0.01fF
C35951 AND2X1_LOC_212/A OR2X1_LOC_7/A 0.18fF
C35952 OR2X1_LOC_574/A OR2X1_LOC_596/A 0.01fF
C35953 OR2X1_LOC_524/Y AND2X1_LOC_676/a_8_24# 0.29fF
C35954 OR2X1_LOC_853/a_8_216# OR2X1_LOC_857/a_8_216# 0.47fF
C35955 OR2X1_LOC_518/a_8_216# OR2X1_LOC_111/Y 0.13fF
C35956 AND2X1_LOC_91/B OR2X1_LOC_859/A 0.07fF
C35957 OR2X1_LOC_571/a_8_216# OR2X1_LOC_571/B 0.10fF
C35958 OR2X1_LOC_643/A OR2X1_LOC_66/A 0.04fF
C35959 OR2X1_LOC_269/Y AND2X1_LOC_36/Y 0.02fF
C35960 OR2X1_LOC_778/Y OR2X1_LOC_66/A 0.14fF
C35961 OR2X1_LOC_71/Y AND2X1_LOC_772/Y 0.01fF
C35962 OR2X1_LOC_51/Y OR2X1_LOC_418/Y 0.01fF
C35963 VDD OR2X1_LOC_585/A 1.48fF
C35964 OR2X1_LOC_369/Y AND2X1_LOC_784/A 0.05fF
C35965 AND2X1_LOC_512/Y AND2X1_LOC_365/A 0.03fF
C35966 OR2X1_LOC_323/A AND2X1_LOC_831/Y 0.01fF
C35967 AND2X1_LOC_486/Y OR2X1_LOC_48/B 3.03fF
C35968 OR2X1_LOC_814/A OR2X1_LOC_362/a_36_216# 0.00fF
C35969 OR2X1_LOC_604/A OR2X1_LOC_420/Y 0.08fF
C35970 AND2X1_LOC_375/a_36_24# D_INPUT_5 0.00fF
C35971 AND2X1_LOC_454/a_8_24# AND2X1_LOC_454/A 0.03fF
C35972 AND2X1_LOC_358/Y OR2X1_LOC_46/A 0.01fF
C35973 OR2X1_LOC_681/a_8_216# OR2X1_LOC_743/A 0.07fF
C35974 OR2X1_LOC_667/Y OR2X1_LOC_278/Y 0.01fF
C35975 AND2X1_LOC_486/Y OR2X1_LOC_18/Y 0.04fF
C35976 OR2X1_LOC_49/A AND2X1_LOC_672/B 0.08fF
C35977 AND2X1_LOC_702/Y INPUT_0 0.03fF
C35978 AND2X1_LOC_707/a_8_24# OR2X1_LOC_7/A 0.03fF
C35979 OR2X1_LOC_625/a_8_216# OR2X1_LOC_278/Y 0.01fF
C35980 OR2X1_LOC_160/A OR2X1_LOC_785/B 0.11fF
C35981 OR2X1_LOC_161/A OR2X1_LOC_575/A 0.04fF
C35982 OR2X1_LOC_624/A OR2X1_LOC_61/Y 0.10fF
C35983 OR2X1_LOC_473/a_8_216# OR2X1_LOC_805/A 0.03fF
C35984 OR2X1_LOC_476/B OR2X1_LOC_654/a_8_216# 0.03fF
C35985 OR2X1_LOC_244/A OR2X1_LOC_572/a_36_216# 0.01fF
C35986 OR2X1_LOC_179/a_8_216# OR2X1_LOC_36/Y 0.07fF
C35987 OR2X1_LOC_335/B AND2X1_LOC_603/a_8_24# 0.02fF
C35988 OR2X1_LOC_329/B OR2X1_LOC_312/Y 0.29fF
C35989 AND2X1_LOC_59/Y AND2X1_LOC_328/a_8_24# 0.20fF
C35990 OR2X1_LOC_844/B OR2X1_LOC_493/Y 0.01fF
C35991 OR2X1_LOC_686/A AND2X1_LOC_51/Y 0.01fF
C35992 OR2X1_LOC_100/Y AND2X1_LOC_81/B 0.01fF
C35993 AND2X1_LOC_512/Y OR2X1_LOC_43/A 0.02fF
C35994 OR2X1_LOC_329/Y OR2X1_LOC_64/Y 0.01fF
C35995 AND2X1_LOC_36/Y OR2X1_LOC_196/a_8_216# 0.01fF
C35996 AND2X1_LOC_148/Y AND2X1_LOC_657/Y 0.30fF
C35997 AND2X1_LOC_339/a_8_24# AND2X1_LOC_219/Y 0.23fF
C35998 OR2X1_LOC_650/Y OR2X1_LOC_654/a_8_216# 0.03fF
C35999 OR2X1_LOC_185/A OR2X1_LOC_655/a_8_216# 0.01fF
C36000 OR2X1_LOC_446/Y AND2X1_LOC_44/Y 0.28fF
C36001 OR2X1_LOC_313/a_8_216# OR2X1_LOC_427/A 0.01fF
C36002 OR2X1_LOC_447/Y OR2X1_LOC_161/B 0.12fF
C36003 AND2X1_LOC_805/Y OR2X1_LOC_39/A 0.00fF
C36004 OR2X1_LOC_479/Y OR2X1_LOC_803/A 0.03fF
C36005 AND2X1_LOC_211/B OR2X1_LOC_310/Y 0.08fF
C36006 AND2X1_LOC_789/a_8_24# OR2X1_LOC_44/Y 0.01fF
C36007 OR2X1_LOC_61/B OR2X1_LOC_87/A 0.00fF
C36008 AND2X1_LOC_253/a_8_24# OR2X1_LOC_269/B 0.04fF
C36009 OR2X1_LOC_186/Y OR2X1_LOC_532/B 1.45fF
C36010 OR2X1_LOC_6/B OR2X1_LOC_19/B 0.08fF
C36011 AND2X1_LOC_348/A AND2X1_LOC_348/Y 0.04fF
C36012 OR2X1_LOC_256/Y AND2X1_LOC_363/A 0.00fF
C36013 AND2X1_LOC_344/a_8_24# AND2X1_LOC_359/a_8_24# 0.23fF
C36014 OR2X1_LOC_427/A AND2X1_LOC_470/A 0.01fF
C36015 OR2X1_LOC_106/Y AND2X1_LOC_116/a_8_24# 0.07fF
C36016 OR2X1_LOC_609/A AND2X1_LOC_647/a_8_24# 0.11fF
C36017 OR2X1_LOC_264/Y OR2X1_LOC_218/a_8_216# 0.39fF
C36018 OR2X1_LOC_40/Y AND2X1_LOC_727/A 0.03fF
C36019 AND2X1_LOC_697/a_36_24# OR2X1_LOC_78/A 0.01fF
C36020 OR2X1_LOC_502/A OR2X1_LOC_449/B 10.85fF
C36021 AND2X1_LOC_90/a_8_24# AND2X1_LOC_47/Y 0.02fF
C36022 OR2X1_LOC_840/A OR2X1_LOC_155/A 0.02fF
C36023 AND2X1_LOC_348/A OR2X1_LOC_753/A 0.01fF
C36024 OR2X1_LOC_599/A AND2X1_LOC_832/a_8_24# 0.02fF
C36025 OR2X1_LOC_508/a_36_216# OR2X1_LOC_532/B 0.00fF
C36026 AND2X1_LOC_811/a_36_24# AND2X1_LOC_811/B 0.01fF
C36027 OR2X1_LOC_689/A OR2X1_LOC_585/A 0.01fF
C36028 AND2X1_LOC_729/B OR2X1_LOC_59/Y 0.03fF
C36029 AND2X1_LOC_716/a_8_24# OR2X1_LOC_18/Y 0.01fF
C36030 AND2X1_LOC_120/a_8_24# AND2X1_LOC_474/A 0.01fF
C36031 AND2X1_LOC_40/Y AND2X1_LOC_481/a_8_24# 0.05fF
C36032 OR2X1_LOC_340/Y OR2X1_LOC_350/a_8_216# 0.07fF
C36033 OR2X1_LOC_235/Y OR2X1_LOC_278/Y 0.01fF
C36034 D_INPUT_0 OR2X1_LOC_641/A 0.07fF
C36035 OR2X1_LOC_160/A OR2X1_LOC_687/Y 0.03fF
C36036 AND2X1_LOC_175/B OR2X1_LOC_6/A 0.01fF
C36037 VDD AND2X1_LOC_634/Y 0.45fF
C36038 OR2X1_LOC_850/B OR2X1_LOC_850/A 0.18fF
C36039 OR2X1_LOC_3/Y AND2X1_LOC_266/a_8_24# 0.01fF
C36040 OR2X1_LOC_47/Y OR2X1_LOC_373/Y 1.57fF
C36041 OR2X1_LOC_101/a_8_216# AND2X1_LOC_3/Y 0.01fF
C36042 OR2X1_LOC_113/A OR2X1_LOC_66/A 0.03fF
C36043 AND2X1_LOC_578/a_8_24# AND2X1_LOC_580/A 0.01fF
C36044 OR2X1_LOC_66/Y OR2X1_LOC_392/B 0.03fF
C36045 OR2X1_LOC_375/A OR2X1_LOC_213/B 0.01fF
C36046 AND2X1_LOC_73/a_8_24# OR2X1_LOC_19/B 0.01fF
C36047 OR2X1_LOC_231/A AND2X1_LOC_3/Y 0.03fF
C36048 OR2X1_LOC_519/a_8_216# AND2X1_LOC_211/B 0.05fF
C36049 OR2X1_LOC_185/A OR2X1_LOC_810/A 0.03fF
C36050 OR2X1_LOC_448/B AND2X1_LOC_697/a_36_24# 0.01fF
C36051 OR2X1_LOC_40/Y OR2X1_LOC_95/Y 5.63fF
C36052 OR2X1_LOC_40/Y AND2X1_LOC_440/a_8_24# 0.02fF
C36053 OR2X1_LOC_359/A OR2X1_LOC_814/A 0.01fF
C36054 OR2X1_LOC_22/A OR2X1_LOC_25/Y 0.11fF
C36055 OR2X1_LOC_111/Y AND2X1_LOC_112/a_8_24# 0.24fF
C36056 AND2X1_LOC_657/a_36_24# AND2X1_LOC_657/Y 0.00fF
C36057 OR2X1_LOC_485/Y AND2X1_LOC_810/Y 0.02fF
C36058 AND2X1_LOC_326/A AND2X1_LOC_863/a_8_24# 0.20fF
C36059 OR2X1_LOC_84/Y OR2X1_LOC_161/B 0.24fF
C36060 OR2X1_LOC_632/a_8_216# OR2X1_LOC_62/B 0.01fF
C36061 AND2X1_LOC_449/Y AND2X1_LOC_454/A 0.09fF
C36062 AND2X1_LOC_575/Y AND2X1_LOC_579/a_8_24# 0.19fF
C36063 OR2X1_LOC_308/A AND2X1_LOC_31/Y 0.01fF
C36064 AND2X1_LOC_22/Y OR2X1_LOC_358/A 0.03fF
C36065 AND2X1_LOC_807/Y OR2X1_LOC_7/A 0.19fF
C36066 AND2X1_LOC_40/Y AND2X1_LOC_442/a_8_24# 0.01fF
C36067 AND2X1_LOC_3/Y OR2X1_LOC_340/Y 0.01fF
C36068 OR2X1_LOC_502/A OR2X1_LOC_121/B 0.07fF
C36069 OR2X1_LOC_490/a_36_216# OR2X1_LOC_67/Y 0.00fF
C36070 AND2X1_LOC_337/B AND2X1_LOC_436/B 0.02fF
C36071 OR2X1_LOC_707/A AND2X1_LOC_3/Y 0.04fF
C36072 AND2X1_LOC_89/a_8_24# AND2X1_LOC_8/Y 0.01fF
C36073 OR2X1_LOC_130/A AND2X1_LOC_3/Y 1.33fF
C36074 OR2X1_LOC_70/Y OR2X1_LOC_109/Y 0.04fF
C36075 OR2X1_LOC_218/a_8_216# OR2X1_LOC_643/A 0.03fF
C36076 OR2X1_LOC_702/A AND2X1_LOC_43/B 0.01fF
C36077 VDD AND2X1_LOC_645/a_8_24# 0.00fF
C36078 OR2X1_LOC_833/Y OR2X1_LOC_374/Y 0.16fF
C36079 OR2X1_LOC_493/A AND2X1_LOC_51/Y 0.94fF
C36080 OR2X1_LOC_175/Y OR2X1_LOC_68/B 0.02fF
C36081 OR2X1_LOC_503/Y AND2X1_LOC_509/a_8_24# 0.23fF
C36082 OR2X1_LOC_272/a_36_216# AND2X1_LOC_139/B 0.02fF
C36083 OR2X1_LOC_241/Y OR2X1_LOC_78/A 0.91fF
C36084 AND2X1_LOC_715/A AND2X1_LOC_798/A 0.20fF
C36085 AND2X1_LOC_7/B OR2X1_LOC_789/A 0.03fF
C36086 AND2X1_LOC_44/Y OR2X1_LOC_228/Y 0.03fF
C36087 OR2X1_LOC_272/Y OR2X1_LOC_767/a_8_216# 0.01fF
C36088 OR2X1_LOC_545/A OR2X1_LOC_551/B 0.05fF
C36089 OR2X1_LOC_251/Y OR2X1_LOC_585/A 0.01fF
C36090 AND2X1_LOC_36/Y OR2X1_LOC_469/B 0.28fF
C36091 OR2X1_LOC_648/a_8_216# OR2X1_LOC_61/B 0.47fF
C36092 AND2X1_LOC_292/a_8_24# AND2X1_LOC_3/Y 0.01fF
C36093 OR2X1_LOC_168/Y OR2X1_LOC_788/B 0.03fF
C36094 AND2X1_LOC_44/Y OR2X1_LOC_513/Y 0.01fF
C36095 OR2X1_LOC_68/B AND2X1_LOC_219/A 0.01fF
C36096 OR2X1_LOC_193/A OR2X1_LOC_194/Y 0.37fF
C36097 OR2X1_LOC_146/Y AND2X1_LOC_148/a_8_24# 0.00fF
C36098 OR2X1_LOC_417/Y AND2X1_LOC_453/a_8_24# 0.01fF
C36099 OR2X1_LOC_297/a_8_216# AND2X1_LOC_866/A 0.01fF
C36100 OR2X1_LOC_306/Y AND2X1_LOC_308/a_8_24# 0.10fF
C36101 AND2X1_LOC_612/a_8_24# OR2X1_LOC_647/B 0.02fF
C36102 OR2X1_LOC_577/Y OR2X1_LOC_367/B 0.00fF
C36103 OR2X1_LOC_471/Y OR2X1_LOC_220/B 0.03fF
C36104 AND2X1_LOC_389/a_8_24# OR2X1_LOC_585/A 0.08fF
C36105 OR2X1_LOC_160/A OR2X1_LOC_606/Y 0.03fF
C36106 D_INPUT_0 OR2X1_LOC_730/a_8_216# 0.14fF
C36107 OR2X1_LOC_185/A AND2X1_LOC_133/a_36_24# 0.00fF
C36108 OR2X1_LOC_801/a_8_216# OR2X1_LOC_801/B 0.07fF
C36109 OR2X1_LOC_316/Y AND2X1_LOC_633/Y 0.02fF
C36110 AND2X1_LOC_702/Y OR2X1_LOC_64/Y 0.02fF
C36111 OR2X1_LOC_33/A OR2X1_LOC_33/B 0.07fF
C36112 OR2X1_LOC_841/a_8_216# OR2X1_LOC_223/A 0.01fF
C36113 OR2X1_LOC_679/A AND2X1_LOC_621/Y 0.04fF
C36114 OR2X1_LOC_316/Y D_INPUT_0 0.03fF
C36115 AND2X1_LOC_318/a_8_24# INPUT_1 0.01fF
C36116 OR2X1_LOC_426/A OR2X1_LOC_47/Y 0.00fF
C36117 OR2X1_LOC_527/Y OR2X1_LOC_238/Y 0.00fF
C36118 OR2X1_LOC_656/a_8_216# OR2X1_LOC_99/Y 0.01fF
C36119 OR2X1_LOC_488/Y OR2X1_LOC_7/A 0.10fF
C36120 AND2X1_LOC_699/a_8_24# OR2X1_LOC_78/B 0.01fF
C36121 OR2X1_LOC_95/Y AND2X1_LOC_644/Y 0.01fF
C36122 OR2X1_LOC_517/A AND2X1_LOC_721/A 0.00fF
C36123 OR2X1_LOC_43/A OR2X1_LOC_54/Y 0.28fF
C36124 AND2X1_LOC_31/a_8_24# AND2X1_LOC_51/A 0.03fF
C36125 AND2X1_LOC_658/A AND2X1_LOC_222/Y 0.03fF
C36126 AND2X1_LOC_8/Y OR2X1_LOC_750/A 0.00fF
C36127 OR2X1_LOC_682/Y AND2X1_LOC_685/a_8_24# 0.01fF
C36128 AND2X1_LOC_505/a_36_24# OR2X1_LOC_560/A 0.00fF
C36129 OR2X1_LOC_785/a_8_216# OR2X1_LOC_228/Y 0.01fF
C36130 AND2X1_LOC_81/B OR2X1_LOC_532/B 0.10fF
C36131 AND2X1_LOC_40/Y OR2X1_LOC_84/a_36_216# 0.02fF
C36132 OR2X1_LOC_709/A OR2X1_LOC_714/A 0.04fF
C36133 AND2X1_LOC_138/a_36_24# OR2X1_LOC_417/A 0.01fF
C36134 AND2X1_LOC_64/Y OR2X1_LOC_510/a_8_216# 0.01fF
C36135 AND2X1_LOC_49/a_8_24# OR2X1_LOC_532/B 0.10fF
C36136 OR2X1_LOC_62/B AND2X1_LOC_610/a_8_24# 0.01fF
C36137 OR2X1_LOC_114/Y D_INPUT_0 0.01fF
C36138 AND2X1_LOC_810/Y OR2X1_LOC_39/A 0.10fF
C36139 OR2X1_LOC_31/Y OR2X1_LOC_265/Y 0.10fF
C36140 OR2X1_LOC_532/B OR2X1_LOC_358/B 0.02fF
C36141 OR2X1_LOC_18/Y AND2X1_LOC_660/A 0.16fF
C36142 OR2X1_LOC_70/Y AND2X1_LOC_729/B 0.02fF
C36143 AND2X1_LOC_727/A OR2X1_LOC_7/A 0.03fF
C36144 OR2X1_LOC_51/Y AND2X1_LOC_796/A 0.03fF
C36145 OR2X1_LOC_691/B OR2X1_LOC_771/B 0.10fF
C36146 OR2X1_LOC_62/B AND2X1_LOC_3/Y 0.03fF
C36147 OR2X1_LOC_160/A OR2X1_LOC_786/Y 0.01fF
C36148 OR2X1_LOC_151/Y AND2X1_LOC_47/Y 0.10fF
C36149 AND2X1_LOC_722/a_8_24# OR2X1_LOC_437/A 0.02fF
C36150 OR2X1_LOC_481/A OR2X1_LOC_295/a_8_216# 0.19fF
C36151 OR2X1_LOC_96/B OR2X1_LOC_96/a_8_216# 0.08fF
C36152 INPUT_4 OR2X1_LOC_47/Y 0.06fF
C36153 OR2X1_LOC_256/A OR2X1_LOC_585/A 0.04fF
C36154 AND2X1_LOC_639/A AND2X1_LOC_651/B 0.03fF
C36155 OR2X1_LOC_11/Y OR2X1_LOC_51/B 0.03fF
C36156 OR2X1_LOC_541/B OR2X1_LOC_241/B 0.14fF
C36157 OR2X1_LOC_673/Y AND2X1_LOC_813/a_8_24# 0.01fF
C36158 OR2X1_LOC_824/a_8_216# D_INPUT_0 0.01fF
C36159 OR2X1_LOC_264/Y OR2X1_LOC_559/a_8_216# 0.01fF
C36160 OR2X1_LOC_311/Y AND2X1_LOC_855/a_8_24# 0.01fF
C36161 AND2X1_LOC_538/a_8_24# AND2X1_LOC_729/B 0.01fF
C36162 AND2X1_LOC_95/Y AND2X1_LOC_497/a_8_24# 0.01fF
C36163 OR2X1_LOC_128/B AND2X1_LOC_72/B 0.00fF
C36164 OR2X1_LOC_158/a_8_216# OR2X1_LOC_163/Y 0.40fF
C36165 OR2X1_LOC_95/Y OR2X1_LOC_7/A 0.71fF
C36166 OR2X1_LOC_45/B AND2X1_LOC_776/Y 0.10fF
C36167 OR2X1_LOC_22/Y OR2X1_LOC_615/a_36_216# 0.03fF
C36168 AND2X1_LOC_555/a_36_24# AND2X1_LOC_789/Y 0.01fF
C36169 OR2X1_LOC_517/A AND2X1_LOC_217/a_8_24# 0.03fF
C36170 OR2X1_LOC_604/A AND2X1_LOC_750/a_8_24# 0.09fF
C36171 AND2X1_LOC_48/A OR2X1_LOC_121/B 0.08fF
C36172 AND2X1_LOC_665/a_36_24# AND2X1_LOC_3/Y 0.00fF
C36173 OR2X1_LOC_161/B OR2X1_LOC_556/a_8_216# 0.01fF
C36174 AND2X1_LOC_473/Y AND2X1_LOC_476/a_8_24# 0.11fF
C36175 OR2X1_LOC_429/Y OR2X1_LOC_428/a_36_216# 0.01fF
C36176 AND2X1_LOC_699/a_8_24# OR2X1_LOC_375/A 0.03fF
C36177 OR2X1_LOC_329/B OR2X1_LOC_13/B 0.07fF
C36178 OR2X1_LOC_118/Y AND2X1_LOC_656/a_8_24# 0.01fF
C36179 OR2X1_LOC_696/A AND2X1_LOC_719/Y 0.12fF
C36180 AND2X1_LOC_3/Y AND2X1_LOC_88/Y 0.81fF
C36181 OR2X1_LOC_62/A AND2X1_LOC_42/B 0.78fF
C36182 AND2X1_LOC_64/Y AND2X1_LOC_65/A 0.97fF
C36183 AND2X1_LOC_555/Y AND2X1_LOC_285/a_8_24# 0.01fF
C36184 OR2X1_LOC_816/A OR2X1_LOC_753/a_8_216# 0.02fF
C36185 OR2X1_LOC_808/B OR2X1_LOC_732/A 0.72fF
C36186 AND2X1_LOC_3/Y AND2X1_LOC_39/Y 0.06fF
C36187 OR2X1_LOC_744/A OR2X1_LOC_183/a_8_216# 0.02fF
C36188 AND2X1_LOC_76/Y OR2X1_LOC_521/a_36_216# 0.00fF
C36189 OR2X1_LOC_19/B AND2X1_LOC_47/Y 0.03fF
C36190 AND2X1_LOC_851/B AND2X1_LOC_523/Y 0.09fF
C36191 AND2X1_LOC_64/Y OR2X1_LOC_510/A 0.08fF
C36192 AND2X1_LOC_552/a_36_24# AND2X1_LOC_476/Y 0.01fF
C36193 OR2X1_LOC_680/A AND2X1_LOC_796/A 0.10fF
C36194 OR2X1_LOC_53/Y AND2X1_LOC_193/Y 0.02fF
C36195 OR2X1_LOC_51/Y OR2X1_LOC_743/Y 0.00fF
C36196 OR2X1_LOC_198/a_36_216# AND2X1_LOC_70/Y 0.00fF
C36197 AND2X1_LOC_56/B OR2X1_LOC_742/B 0.01fF
C36198 OR2X1_LOC_277/a_8_216# OR2X1_LOC_47/Y 0.01fF
C36199 OR2X1_LOC_502/A OR2X1_LOC_195/a_8_216# 0.02fF
C36200 OR2X1_LOC_51/Y OR2X1_LOC_171/a_8_216# 0.13fF
C36201 OR2X1_LOC_600/A OR2X1_LOC_748/a_36_216# 0.00fF
C36202 OR2X1_LOC_156/a_8_216# OR2X1_LOC_160/B 0.01fF
C36203 OR2X1_LOC_584/a_8_216# OR2X1_LOC_16/A 0.06fF
C36204 AND2X1_LOC_797/a_8_24# AND2X1_LOC_220/B 0.20fF
C36205 AND2X1_LOC_721/Y AND2X1_LOC_243/Y 0.02fF
C36206 AND2X1_LOC_91/B OR2X1_LOC_66/A 13.85fF
C36207 AND2X1_LOC_338/a_8_24# OR2X1_LOC_171/Y 0.01fF
C36208 OR2X1_LOC_274/Y AND2X1_LOC_36/Y 0.03fF
C36209 AND2X1_LOC_564/B VDD 0.70fF
C36210 AND2X1_LOC_91/B OR2X1_LOC_841/A 0.14fF
C36211 OR2X1_LOC_158/A OR2X1_LOC_12/Y 0.47fF
C36212 VDD OR2X1_LOC_230/Y 0.04fF
C36213 OR2X1_LOC_161/A OR2X1_LOC_735/B 0.01fF
C36214 AND2X1_LOC_223/A GATE_222 0.27fF
C36215 OR2X1_LOC_739/A OR2X1_LOC_730/B 0.78fF
C36216 VDD OR2X1_LOC_530/a_8_216# 0.00fF
C36217 OR2X1_LOC_820/A OR2X1_LOC_748/a_8_216# 0.04fF
C36218 AND2X1_LOC_535/Y OR2X1_LOC_16/A 0.00fF
C36219 OR2X1_LOC_765/Y AND2X1_LOC_770/a_8_24# 0.10fF
C36220 OR2X1_LOC_421/A OR2X1_LOC_692/Y 0.01fF
C36221 AND2X1_LOC_92/Y OR2X1_LOC_703/a_36_216# 0.02fF
C36222 OR2X1_LOC_40/Y OR2X1_LOC_821/Y 0.02fF
C36223 AND2X1_LOC_18/Y OR2X1_LOC_580/B 0.00fF
C36224 OR2X1_LOC_532/B OR2X1_LOC_112/B 0.10fF
C36225 OR2X1_LOC_445/a_8_216# OR2X1_LOC_578/B 0.03fF
C36226 AND2X1_LOC_12/Y AND2X1_LOC_591/a_8_24# 0.01fF
C36227 OR2X1_LOC_151/A OR2X1_LOC_362/A 0.00fF
C36228 OR2X1_LOC_212/A OR2X1_LOC_212/B 0.07fF
C36229 AND2X1_LOC_748/a_8_24# AND2X1_LOC_36/Y -0.00fF
C36230 OR2X1_LOC_19/B OR2X1_LOC_598/A 0.09fF
C36231 OR2X1_LOC_57/Y OR2X1_LOC_56/Y 0.00fF
C36232 OR2X1_LOC_506/A OR2X1_LOC_308/Y 0.05fF
C36233 OR2X1_LOC_615/a_8_216# AND2X1_LOC_562/Y 0.15fF
C36234 AND2X1_LOC_566/B AND2X1_LOC_357/B 0.02fF
C36235 AND2X1_LOC_320/a_8_24# AND2X1_LOC_44/Y 0.01fF
C36236 OR2X1_LOC_124/B OR2X1_LOC_549/A -0.02fF
C36237 OR2X1_LOC_675/A AND2X1_LOC_31/Y 0.01fF
C36238 OR2X1_LOC_660/Y AND2X1_LOC_44/Y 0.24fF
C36239 OR2X1_LOC_680/a_36_216# OR2X1_LOC_677/Y 0.00fF
C36240 AND2X1_LOC_505/a_8_24# OR2X1_LOC_641/A 0.02fF
C36241 OR2X1_LOC_532/B OR2X1_LOC_66/Y 0.03fF
C36242 OR2X1_LOC_648/B AND2X1_LOC_18/Y 0.17fF
C36243 OR2X1_LOC_831/a_36_216# OR2X1_LOC_593/B 0.00fF
C36244 OR2X1_LOC_287/B OR2X1_LOC_580/A 0.01fF
C36245 OR2X1_LOC_865/A OR2X1_LOC_862/A 0.03fF
C36246 OR2X1_LOC_51/Y OR2X1_LOC_13/Y 0.03fF
C36247 AND2X1_LOC_95/Y OR2X1_LOC_333/a_36_216# 0.00fF
C36248 OR2X1_LOC_31/Y AND2X1_LOC_205/a_8_24# 0.01fF
C36249 OR2X1_LOC_440/A OR2X1_LOC_241/B 0.03fF
C36250 OR2X1_LOC_600/A OR2X1_LOC_14/a_8_216# 0.05fF
C36251 OR2X1_LOC_696/A AND2X1_LOC_655/A 0.10fF
C36252 AND2X1_LOC_754/a_8_24# OR2X1_LOC_78/A 0.01fF
C36253 OR2X1_LOC_614/Y OR2X1_LOC_78/B 0.11fF
C36254 AND2X1_LOC_174/a_8_24# OR2X1_LOC_171/Y 0.09fF
C36255 VDD OR2X1_LOC_507/A 0.25fF
C36256 OR2X1_LOC_141/B OR2X1_LOC_141/a_36_216# 0.00fF
C36257 AND2X1_LOC_95/Y OR2X1_LOC_334/a_8_216# 0.01fF
C36258 OR2X1_LOC_434/A OR2X1_LOC_358/A 0.46fF
C36259 AND2X1_LOC_784/Y AND2X1_LOC_469/B 0.02fF
C36260 AND2X1_LOC_392/A AND2X1_LOC_436/Y 0.06fF
C36261 OR2X1_LOC_834/a_8_216# OR2X1_LOC_713/A 0.01fF
C36262 OR2X1_LOC_619/Y OR2X1_LOC_321/a_8_216# 0.02fF
C36263 AND2X1_LOC_566/B AND2X1_LOC_303/a_8_24# 0.01fF
C36264 OR2X1_LOC_51/Y OR2X1_LOC_627/Y 0.01fF
C36265 OR2X1_LOC_158/A OR2X1_LOC_837/Y 0.07fF
C36266 OR2X1_LOC_516/Y OR2X1_LOC_52/B 0.03fF
C36267 OR2X1_LOC_188/Y OR2X1_LOC_541/B 0.01fF
C36268 AND2X1_LOC_40/Y OR2X1_LOC_294/Y 0.06fF
C36269 AND2X1_LOC_500/Y OR2X1_LOC_51/Y 0.21fF
C36270 OR2X1_LOC_748/A AND2X1_LOC_792/a_8_24# 0.01fF
C36271 AND2X1_LOC_57/Y OR2X1_LOC_269/B 0.00fF
C36272 AND2X1_LOC_172/a_8_24# OR2X1_LOC_648/A 0.01fF
C36273 AND2X1_LOC_784/Y AND2X1_LOC_733/Y 0.00fF
C36274 OR2X1_LOC_794/a_8_216# OR2X1_LOC_593/B 0.04fF
C36275 OR2X1_LOC_831/a_8_216# OR2X1_LOC_831/B 0.05fF
C36276 OR2X1_LOC_46/A OR2X1_LOC_71/A 0.08fF
C36277 AND2X1_LOC_522/a_36_24# OR2X1_LOC_523/Y 0.00fF
C36278 OR2X1_LOC_18/Y AND2X1_LOC_231/a_36_24# 0.01fF
C36279 AND2X1_LOC_658/B AND2X1_LOC_659/a_8_24# 0.01fF
C36280 OR2X1_LOC_485/A OR2X1_LOC_183/Y 0.01fF
C36281 AND2X1_LOC_39/Y OR2X1_LOC_194/a_8_216# 0.47fF
C36282 OR2X1_LOC_17/Y D_INPUT_6 1.09fF
C36283 AND2X1_LOC_716/Y AND2X1_LOC_180/a_8_24# 0.03fF
C36284 OR2X1_LOC_158/A OR2X1_LOC_422/a_8_216# 0.01fF
C36285 OR2X1_LOC_375/A OR2X1_LOC_779/A 0.01fF
C36286 AND2X1_LOC_570/Y AND2X1_LOC_663/A 0.05fF
C36287 AND2X1_LOC_95/Y OR2X1_LOC_34/a_36_216# 0.00fF
C36288 OR2X1_LOC_851/B OR2X1_LOC_851/A 0.19fF
C36289 OR2X1_LOC_49/A OR2X1_LOC_377/A 0.10fF
C36290 AND2X1_LOC_397/a_8_24# OR2X1_LOC_78/A 0.01fF
C36291 OR2X1_LOC_751/Y OR2X1_LOC_6/B 0.02fF
C36292 AND2X1_LOC_326/a_8_24# OR2X1_LOC_437/A 0.03fF
C36293 AND2X1_LOC_571/B AND2X1_LOC_489/Y 0.01fF
C36294 OR2X1_LOC_161/A OR2X1_LOC_161/B 0.58fF
C36295 AND2X1_LOC_543/Y OR2X1_LOC_26/Y 0.01fF
C36296 OR2X1_LOC_456/Y OR2X1_LOC_577/Y 0.01fF
C36297 OR2X1_LOC_154/A OR2X1_LOC_139/A 12.45fF
C36298 AND2X1_LOC_40/Y OR2X1_LOC_641/A 0.03fF
C36299 AND2X1_LOC_19/Y AND2X1_LOC_20/a_8_24# 0.11fF
C36300 AND2X1_LOC_347/Y VDD 0.12fF
C36301 AND2X1_LOC_70/Y OR2X1_LOC_174/A 0.01fF
C36302 AND2X1_LOC_95/Y OR2X1_LOC_486/Y 0.06fF
C36303 VDD AND2X1_LOC_857/Y 0.29fF
C36304 AND2X1_LOC_16/a_8_24# OR2X1_LOC_596/A 0.01fF
C36305 AND2X1_LOC_35/Y AND2X1_LOC_219/A 0.07fF
C36306 OR2X1_LOC_97/A OR2X1_LOC_87/A 0.05fF
C36307 OR2X1_LOC_6/A AND2X1_LOC_214/a_8_24# 0.01fF
C36308 OR2X1_LOC_326/B AND2X1_LOC_110/Y 0.02fF
C36309 AND2X1_LOC_576/Y AND2X1_LOC_244/A 0.01fF
C36310 OR2X1_LOC_427/A AND2X1_LOC_605/a_36_24# 0.00fF
C36311 OR2X1_LOC_139/A OR2X1_LOC_267/A 0.01fF
C36312 OR2X1_LOC_49/A OR2X1_LOC_85/A 0.33fF
C36313 OR2X1_LOC_774/Y OR2X1_LOC_866/B 0.20fF
C36314 AND2X1_LOC_572/A OR2X1_LOC_595/A 0.02fF
C36315 OR2X1_LOC_377/A OR2X1_LOC_596/A 0.02fF
C36316 AND2X1_LOC_64/Y OR2X1_LOC_204/a_8_216# 0.05fF
C36317 OR2X1_LOC_715/B OR2X1_LOC_185/A 0.05fF
C36318 AND2X1_LOC_185/a_8_24# OR2X1_LOC_56/A 0.04fF
C36319 OR2X1_LOC_678/a_36_216# OR2X1_LOC_678/Y 0.00fF
C36320 OR2X1_LOC_629/a_8_216# OR2X1_LOC_140/B 0.01fF
C36321 OR2X1_LOC_379/Y OR2X1_LOC_598/Y 0.01fF
C36322 OR2X1_LOC_106/Y OR2X1_LOC_490/Y 0.01fF
C36323 OR2X1_LOC_116/A OR2X1_LOC_151/A 0.02fF
C36324 OR2X1_LOC_614/Y OR2X1_LOC_375/A 0.01fF
C36325 AND2X1_LOC_191/Y AND2X1_LOC_220/B 8.46fF
C36326 OR2X1_LOC_653/Y VDD 0.12fF
C36327 OR2X1_LOC_216/A OR2X1_LOC_78/A 0.29fF
C36328 OR2X1_LOC_678/Y AND2X1_LOC_41/A 0.00fF
C36329 OR2X1_LOC_198/a_8_216# AND2X1_LOC_51/Y 0.03fF
C36330 OR2X1_LOC_149/B OR2X1_LOC_546/B 0.10fF
C36331 AND2X1_LOC_540/a_8_24# OR2X1_LOC_744/A 0.02fF
C36332 AND2X1_LOC_42/B OR2X1_LOC_397/Y 0.14fF
C36333 AND2X1_LOC_539/Y AND2X1_LOC_390/B 0.02fF
C36334 OR2X1_LOC_185/A OR2X1_LOC_543/A 0.48fF
C36335 AND2X1_LOC_41/A OR2X1_LOC_294/a_8_216# 0.08fF
C36336 OR2X1_LOC_600/A OR2X1_LOC_250/a_36_216# 0.00fF
C36337 AND2X1_LOC_711/Y AND2X1_LOC_220/B 0.09fF
C36338 AND2X1_LOC_719/Y AND2X1_LOC_458/Y 0.08fF
C36339 OR2X1_LOC_449/a_8_216# OR2X1_LOC_161/B 0.02fF
C36340 AND2X1_LOC_386/a_8_24# AND2X1_LOC_44/Y 0.17fF
C36341 AND2X1_LOC_91/B AND2X1_LOC_176/a_36_24# 0.01fF
C36342 OR2X1_LOC_799/A OR2X1_LOC_66/A 0.12fF
C36343 OR2X1_LOC_862/A OR2X1_LOC_391/A 0.15fF
C36344 OR2X1_LOC_691/A OR2X1_LOC_688/a_8_216# 0.01fF
C36345 AND2X1_LOC_59/Y OR2X1_LOC_676/Y 0.50fF
C36346 OR2X1_LOC_3/Y OR2X1_LOC_428/A 0.43fF
C36347 OR2X1_LOC_589/A OR2X1_LOC_26/Y 0.03fF
C36348 AND2X1_LOC_130/a_8_24# AND2X1_LOC_361/A 0.02fF
C36349 OR2X1_LOC_31/Y OR2X1_LOC_183/a_8_216# 0.01fF
C36350 AND2X1_LOC_859/a_8_24# AND2X1_LOC_860/A 0.02fF
C36351 OR2X1_LOC_813/Y OR2X1_LOC_71/A 0.01fF
C36352 AND2X1_LOC_663/B AND2X1_LOC_580/a_8_24# 0.01fF
C36353 VDD OR2X1_LOC_848/B 0.05fF
C36354 OR2X1_LOC_641/Y OR2X1_LOC_375/A 0.04fF
C36355 AND2X1_LOC_705/Y OR2X1_LOC_485/A 0.21fF
C36356 OR2X1_LOC_680/A OR2X1_LOC_627/Y 0.03fF
C36357 OR2X1_LOC_697/a_8_216# OR2X1_LOC_427/A 0.06fF
C36358 OR2X1_LOC_269/B OR2X1_LOC_719/a_36_216# 0.00fF
C36359 OR2X1_LOC_97/a_8_216# AND2X1_LOC_44/Y 0.01fF
C36360 AND2X1_LOC_500/Y OR2X1_LOC_680/A 0.03fF
C36361 OR2X1_LOC_3/Y OR2X1_LOC_595/A 1.89fF
C36362 OR2X1_LOC_499/a_8_216# OR2X1_LOC_78/A 0.01fF
C36363 OR2X1_LOC_791/B OR2X1_LOC_287/A 0.20fF
C36364 OR2X1_LOC_589/A OR2X1_LOC_89/A 0.07fF
C36365 AND2X1_LOC_697/a_8_24# OR2X1_LOC_713/A 0.02fF
C36366 OR2X1_LOC_531/Y AND2X1_LOC_807/Y 0.08fF
C36367 AND2X1_LOC_326/B AND2X1_LOC_354/B 0.01fF
C36368 AND2X1_LOC_51/Y OR2X1_LOC_161/B 0.70fF
C36369 AND2X1_LOC_840/a_8_24# AND2X1_LOC_851/A 0.00fF
C36370 AND2X1_LOC_767/a_8_24# OR2X1_LOC_78/Y 0.00fF
C36371 D_GATE_662 AND2X1_LOC_815/a_8_24# 0.03fF
C36372 OR2X1_LOC_235/B OR2X1_LOC_137/B 0.01fF
C36373 AND2X1_LOC_535/Y AND2X1_LOC_336/a_8_24# 0.01fF
C36374 AND2X1_LOC_738/B OR2X1_LOC_36/Y 0.16fF
C36375 OR2X1_LOC_45/B OR2X1_LOC_278/A 0.15fF
C36376 OR2X1_LOC_668/a_36_216# OR2X1_LOC_721/Y 0.00fF
C36377 AND2X1_LOC_77/a_8_24# OR2X1_LOC_633/A 0.04fF
C36378 OR2X1_LOC_36/Y OR2X1_LOC_56/A 1.58fF
C36379 OR2X1_LOC_158/A OR2X1_LOC_272/Y 0.03fF
C36380 AND2X1_LOC_721/a_8_24# OR2X1_LOC_278/Y 0.01fF
C36381 AND2X1_LOC_48/a_8_24# OR2X1_LOC_161/A 0.04fF
C36382 AND2X1_LOC_89/a_8_24# AND2X1_LOC_92/Y 0.01fF
C36383 AND2X1_LOC_861/B OR2X1_LOC_39/A 0.08fF
C36384 OR2X1_LOC_284/a_8_216# OR2X1_LOC_269/B 0.07fF
C36385 OR2X1_LOC_468/Y OR2X1_LOC_78/A 0.03fF
C36386 AND2X1_LOC_732/a_36_24# OR2X1_LOC_599/A 0.00fF
C36387 OR2X1_LOC_549/Y OR2X1_LOC_577/B 0.30fF
C36388 OR2X1_LOC_600/A AND2X1_LOC_717/B 0.03fF
C36389 AND2X1_LOC_209/a_8_24# AND2X1_LOC_191/Y 0.06fF
C36390 OR2X1_LOC_324/B AND2X1_LOC_56/B 0.01fF
C36391 AND2X1_LOC_804/Y AND2X1_LOC_808/a_8_24# 0.04fF
C36392 OR2X1_LOC_715/B OR2X1_LOC_435/Y 0.28fF
C36393 OR2X1_LOC_97/A OR2X1_LOC_648/a_8_216# 0.01fF
C36394 OR2X1_LOC_808/B OR2X1_LOC_375/A 0.03fF
C36395 OR2X1_LOC_786/Y OR2X1_LOC_130/Y 0.32fF
C36396 AND2X1_LOC_744/a_8_24# OR2X1_LOC_87/A 0.01fF
C36397 AND2X1_LOC_727/Y AND2X1_LOC_811/Y 0.00fF
C36398 OR2X1_LOC_622/A OR2X1_LOC_624/B 0.73fF
C36399 OR2X1_LOC_130/A OR2X1_LOC_775/a_8_216# 0.06fF
C36400 INPUT_0 AND2X1_LOC_688/a_8_24# 0.01fF
C36401 AND2X1_LOC_658/A OR2X1_LOC_74/A 0.13fF
C36402 OR2X1_LOC_164/Y AND2X1_LOC_840/B 0.11fF
C36403 AND2X1_LOC_160/Y OR2X1_LOC_743/A 0.01fF
C36404 OR2X1_LOC_631/B OR2X1_LOC_294/a_8_216# 0.06fF
C36405 OR2X1_LOC_437/A AND2X1_LOC_657/A 0.07fF
C36406 OR2X1_LOC_188/Y OR2X1_LOC_440/A 0.02fF
C36407 AND2X1_LOC_91/B OR2X1_LOC_84/A 0.02fF
C36408 OR2X1_LOC_427/A AND2X1_LOC_470/B 0.01fF
C36409 OR2X1_LOC_517/A AND2X1_LOC_361/A 0.09fF
C36410 OR2X1_LOC_606/Y AND2X1_LOC_607/a_8_24# 0.01fF
C36411 OR2X1_LOC_89/A OR2X1_LOC_297/A 0.01fF
C36412 AND2X1_LOC_536/a_8_24# OR2X1_LOC_161/A 0.03fF
C36413 OR2X1_LOC_87/A OR2X1_LOC_475/B 0.10fF
C36414 OR2X1_LOC_696/A OR2X1_LOC_599/Y 0.10fF
C36415 AND2X1_LOC_391/Y AND2X1_LOC_554/B 0.29fF
C36416 OR2X1_LOC_825/Y OR2X1_LOC_600/A 0.21fF
C36417 AND2X1_LOC_353/a_8_24# AND2X1_LOC_727/A 0.11fF
C36418 OR2X1_LOC_744/A AND2X1_LOC_155/Y 0.09fF
C36419 AND2X1_LOC_554/B OR2X1_LOC_91/A 0.01fF
C36420 OR2X1_LOC_185/A OR2X1_LOC_215/Y 0.21fF
C36421 OR2X1_LOC_833/Y OR2X1_LOC_532/B 0.02fF
C36422 AND2X1_LOC_560/B AND2X1_LOC_113/a_8_24# 0.01fF
C36423 AND2X1_LOC_576/a_36_24# OR2X1_LOC_427/A 0.01fF
C36424 OR2X1_LOC_402/Y OR2X1_LOC_404/a_36_216# 0.00fF
C36425 AND2X1_LOC_654/B OR2X1_LOC_26/Y 0.05fF
C36426 AND2X1_LOC_160/a_36_24# OR2X1_LOC_52/B 0.01fF
C36427 AND2X1_LOC_351/a_36_24# OR2X1_LOC_31/Y 0.01fF
C36428 AND2X1_LOC_343/a_8_24# OR2X1_LOC_517/A 0.01fF
C36429 AND2X1_LOC_810/Y AND2X1_LOC_727/B 0.00fF
C36430 OR2X1_LOC_9/Y INPUT_1 0.00fF
C36431 OR2X1_LOC_105/a_36_216# OR2X1_LOC_287/B 0.00fF
C36432 AND2X1_LOC_314/a_8_24# AND2X1_LOC_56/B 0.03fF
C36433 OR2X1_LOC_160/A OR2X1_LOC_828/B 0.03fF
C36434 OR2X1_LOC_689/a_8_216# OR2X1_LOC_43/A 0.01fF
C36435 OR2X1_LOC_179/Y OR2X1_LOC_7/A 0.01fF
C36436 OR2X1_LOC_631/B OR2X1_LOC_811/A 0.07fF
C36437 OR2X1_LOC_591/A OR2X1_LOC_48/B 0.02fF
C36438 OR2X1_LOC_615/Y OR2X1_LOC_816/A 0.58fF
C36439 OR2X1_LOC_670/a_8_216# OR2X1_LOC_823/a_8_216# 0.47fF
C36440 OR2X1_LOC_160/A OR2X1_LOC_835/B 0.16fF
C36441 OR2X1_LOC_757/A OR2X1_LOC_665/a_8_216# 0.01fF
C36442 AND2X1_LOC_326/A OR2X1_LOC_91/A 0.00fF
C36443 AND2X1_LOC_719/Y AND2X1_LOC_849/a_8_24# 0.23fF
C36444 AND2X1_LOC_59/Y OR2X1_LOC_462/B 0.02fF
C36445 AND2X1_LOC_553/A OR2X1_LOC_485/A 0.01fF
C36446 OR2X1_LOC_599/A AND2X1_LOC_621/Y 0.02fF
C36447 OR2X1_LOC_687/A AND2X1_LOC_425/Y 0.01fF
C36448 OR2X1_LOC_377/A OR2X1_LOC_87/B 0.04fF
C36449 OR2X1_LOC_495/Y OR2X1_LOC_89/A 0.03fF
C36450 OR2X1_LOC_124/a_8_216# OR2X1_LOC_814/A 0.06fF
C36451 OR2X1_LOC_808/B OR2X1_LOC_605/B 0.06fF
C36452 AND2X1_LOC_593/Y AND2X1_LOC_661/A 0.01fF
C36453 AND2X1_LOC_228/Y AND2X1_LOC_716/a_8_24# 0.10fF
C36454 AND2X1_LOC_566/a_8_24# OR2X1_LOC_619/Y 0.06fF
C36455 AND2X1_LOC_706/Y AND2X1_LOC_648/B 0.02fF
C36456 OR2X1_LOC_216/a_8_216# OR2X1_LOC_475/B 0.05fF
C36457 OR2X1_LOC_662/A OR2X1_LOC_649/B 0.16fF
C36458 AND2X1_LOC_387/a_8_24# OR2X1_LOC_532/B 0.01fF
C36459 AND2X1_LOC_61/Y INPUT_1 0.14fF
C36460 AND2X1_LOC_848/Y OR2X1_LOC_44/Y 0.04fF
C36461 AND2X1_LOC_110/Y AND2X1_LOC_47/Y 0.03fF
C36462 OR2X1_LOC_3/B INPUT_7 0.00fF
C36463 OR2X1_LOC_46/A OR2X1_LOC_59/Y 0.04fF
C36464 OR2X1_LOC_687/Y OR2X1_LOC_685/B 0.03fF
C36465 AND2X1_LOC_90/a_8_24# D_INPUT_1 0.01fF
C36466 OR2X1_LOC_493/B OR2X1_LOC_532/B 0.21fF
C36467 OR2X1_LOC_604/A OR2X1_LOC_751/A 0.17fF
C36468 OR2X1_LOC_744/A AND2X1_LOC_633/Y 0.01fF
C36469 OR2X1_LOC_16/A OR2X1_LOC_29/a_8_216# 0.06fF
C36470 AND2X1_LOC_22/Y AND2X1_LOC_497/a_8_24# 0.05fF
C36471 AND2X1_LOC_99/a_8_24# OR2X1_LOC_64/Y 0.01fF
C36472 OR2X1_LOC_362/B OR2X1_LOC_807/a_8_216# 0.01fF
C36473 OR2X1_LOC_325/B OR2X1_LOC_440/A 1.24fF
C36474 INPUT_0 OR2X1_LOC_62/B 0.04fF
C36475 AND2X1_LOC_487/a_8_24# AND2X1_LOC_3/Y 0.02fF
C36476 AND2X1_LOC_192/Y AND2X1_LOC_740/B 0.03fF
C36477 AND2X1_LOC_379/a_8_24# OR2X1_LOC_26/Y 0.04fF
C36478 OR2X1_LOC_291/a_36_216# OR2X1_LOC_74/A 0.00fF
C36479 OR2X1_LOC_756/B OR2X1_LOC_846/A 0.01fF
C36480 AND2X1_LOC_695/a_36_24# OR2X1_LOC_449/B 0.01fF
C36481 OR2X1_LOC_673/Y OR2X1_LOC_845/a_8_216# 0.01fF
C36482 OR2X1_LOC_744/A D_INPUT_0 0.03fF
C36483 OR2X1_LOC_420/Y AND2X1_LOC_447/a_8_24# 0.23fF
C36484 AND2X1_LOC_554/B AND2X1_LOC_573/A 0.15fF
C36485 OR2X1_LOC_161/B OR2X1_LOC_551/B 0.17fF
C36486 AND2X1_LOC_20/a_36_24# D_INPUT_0 0.00fF
C36487 OR2X1_LOC_154/A OR2X1_LOC_208/a_8_216# 0.05fF
C36488 OR2X1_LOC_824/Y AND2X1_LOC_836/a_8_24# 0.06fF
C36489 OR2X1_LOC_43/A OR2X1_LOC_26/Y 0.13fF
C36490 OR2X1_LOC_485/A OR2X1_LOC_511/Y 0.00fF
C36491 OR2X1_LOC_531/Y OR2X1_LOC_95/Y 0.02fF
C36492 AND2X1_LOC_227/Y OR2X1_LOC_59/Y 0.10fF
C36493 OR2X1_LOC_739/Y OR2X1_LOC_740/B 0.08fF
C36494 OR2X1_LOC_840/A OR2X1_LOC_814/A 0.02fF
C36495 OR2X1_LOC_139/A OR2X1_LOC_560/A 0.05fF
C36496 AND2X1_LOC_307/Y OR2X1_LOC_48/B 0.54fF
C36497 AND2X1_LOC_40/Y OR2X1_LOC_444/a_8_216# 0.01fF
C36498 OR2X1_LOC_589/A AND2X1_LOC_202/a_8_24# 0.01fF
C36499 OR2X1_LOC_248/Y OR2X1_LOC_585/A 0.09fF
C36500 OR2X1_LOC_261/A AND2X1_LOC_847/Y 0.02fF
C36501 OR2X1_LOC_47/Y AND2X1_LOC_447/Y 0.10fF
C36502 AND2X1_LOC_795/Y AND2X1_LOC_778/Y 0.26fF
C36503 OR2X1_LOC_485/A OR2X1_LOC_248/a_8_216# -0.00fF
C36504 OR2X1_LOC_856/B AND2X1_LOC_48/A 0.07fF
C36505 OR2X1_LOC_43/A OR2X1_LOC_89/A 0.53fF
C36506 OR2X1_LOC_13/B OR2X1_LOC_525/a_8_216# 0.07fF
C36507 AND2X1_LOC_40/Y OR2X1_LOC_286/a_8_216# 0.01fF
C36508 OR2X1_LOC_731/A OR2X1_LOC_550/B 0.03fF
C36509 AND2X1_LOC_3/Y OR2X1_LOC_449/B 0.03fF
C36510 OR2X1_LOC_164/Y OR2X1_LOC_31/Y 0.04fF
C36511 OR2X1_LOC_36/Y OR2X1_LOC_291/A 0.56fF
C36512 OR2X1_LOC_864/A OR2X1_LOC_557/A 0.03fF
C36513 AND2X1_LOC_412/a_36_24# OR2X1_LOC_240/A 0.01fF
C36514 OR2X1_LOC_377/A AND2X1_LOC_79/a_8_24# 0.01fF
C36515 OR2X1_LOC_22/a_8_216# OR2X1_LOC_17/Y 0.01fF
C36516 OR2X1_LOC_774/Y OR2X1_LOC_557/A 0.00fF
C36517 OR2X1_LOC_595/A AND2X1_LOC_772/a_8_24# 0.03fF
C36518 OR2X1_LOC_485/A AND2X1_LOC_294/a_8_24# 0.01fF
C36519 AND2X1_LOC_88/a_8_24# AND2X1_LOC_3/Y 0.00fF
C36520 OR2X1_LOC_205/Y OR2X1_LOC_78/A 0.03fF
C36521 OR2X1_LOC_404/A OR2X1_LOC_402/Y 0.18fF
C36522 OR2X1_LOC_462/a_8_216# AND2X1_LOC_56/B 0.05fF
C36523 OR2X1_LOC_141/B AND2X1_LOC_42/B 0.03fF
C36524 INPUT_0 AND2X1_LOC_39/Y 0.01fF
C36525 OR2X1_LOC_128/B AND2X1_LOC_127/a_36_24# 0.00fF
C36526 AND2X1_LOC_738/B OR2X1_LOC_419/Y 0.10fF
C36527 OR2X1_LOC_60/a_8_216# OR2X1_LOC_26/Y 0.06fF
C36528 OR2X1_LOC_419/Y OR2X1_LOC_56/A 0.05fF
C36529 OR2X1_LOC_195/A AND2X1_LOC_43/a_36_24# 0.00fF
C36530 AND2X1_LOC_477/A OR2X1_LOC_39/A 0.10fF
C36531 AND2X1_LOC_117/a_8_24# OR2X1_LOC_633/B 0.01fF
C36532 AND2X1_LOC_663/A OR2X1_LOC_406/A 0.05fF
C36533 AND2X1_LOC_345/Y AND2X1_LOC_348/a_8_24# 0.03fF
C36534 OR2X1_LOC_461/B OR2X1_LOC_68/B 0.00fF
C36535 OR2X1_LOC_96/B INPUT_1 0.02fF
C36536 AND2X1_LOC_502/a_36_24# OR2X1_LOC_71/Y 0.00fF
C36537 OR2X1_LOC_46/A OR2X1_LOC_820/B 0.04fF
C36538 OR2X1_LOC_54/Y AND2X1_LOC_818/a_36_24# 0.01fF
C36539 AND2X1_LOC_593/Y AND2X1_LOC_810/Y 0.08fF
C36540 OR2X1_LOC_391/A AND2X1_LOC_225/a_36_24# 0.01fF
C36541 AND2X1_LOC_866/A AND2X1_LOC_621/Y 0.01fF
C36542 OR2X1_LOC_87/A OR2X1_LOC_797/A 0.01fF
C36543 AND2X1_LOC_842/B OR2X1_LOC_239/Y 0.00fF
C36544 OR2X1_LOC_562/Y OR2X1_LOC_562/a_8_216# 0.00fF
C36545 OR2X1_LOC_335/A OR2X1_LOC_605/Y 0.02fF
C36546 OR2X1_LOC_121/B AND2X1_LOC_3/Y 0.03fF
C36547 OR2X1_LOC_664/Y AND2X1_LOC_47/Y 0.03fF
C36548 AND2X1_LOC_794/B OR2X1_LOC_437/A 0.07fF
C36549 INPUT_1 AND2X1_LOC_852/Y 0.03fF
C36550 AND2X1_LOC_664/a_8_24# OR2X1_LOC_89/A 0.01fF
C36551 OR2X1_LOC_841/a_36_216# OR2X1_LOC_804/A 0.00fF
C36552 OR2X1_LOC_54/Y AND2X1_LOC_240/Y 0.02fF
C36553 OR2X1_LOC_278/Y D_INPUT_1 0.02fF
C36554 OR2X1_LOC_109/Y OR2X1_LOC_47/Y 0.08fF
C36555 AND2X1_LOC_141/A AND2X1_LOC_216/A 0.23fF
C36556 OR2X1_LOC_406/a_36_216# OR2X1_LOC_95/Y 0.03fF
C36557 OR2X1_LOC_318/Y OR2X1_LOC_804/A 0.03fF
C36558 OR2X1_LOC_774/Y OR2X1_LOC_773/a_36_216# 0.00fF
C36559 OR2X1_LOC_778/B OR2X1_LOC_68/B 0.05fF
C36560 OR2X1_LOC_38/a_8_216# D_INPUT_1 0.00fF
C36561 OR2X1_LOC_66/A OR2X1_LOC_446/B 0.03fF
C36562 AND2X1_LOC_462/Y AND2X1_LOC_472/B 0.00fF
C36563 OR2X1_LOC_856/A AND2X1_LOC_36/Y 0.01fF
C36564 AND2X1_LOC_18/Y OR2X1_LOC_367/a_8_216# 0.01fF
C36565 OR2X1_LOC_70/Y OR2X1_LOC_46/A 0.03fF
C36566 OR2X1_LOC_574/A OR2X1_LOC_532/B 0.41fF
C36567 OR2X1_LOC_66/A OR2X1_LOC_303/B 0.03fF
C36568 VDD OR2X1_LOC_437/A 1.99fF
C36569 OR2X1_LOC_151/A OR2X1_LOC_209/A 0.04fF
C36570 OR2X1_LOC_97/A OR2X1_LOC_390/B 0.01fF
C36571 AND2X1_LOC_512/Y OR2X1_LOC_534/Y 0.02fF
C36572 OR2X1_LOC_756/B OR2X1_LOC_348/B 0.09fF
C36573 AND2X1_LOC_333/a_8_24# OR2X1_LOC_46/A 0.01fF
C36574 OR2X1_LOC_49/A AND2X1_LOC_555/Y 0.03fF
C36575 AND2X1_LOC_514/Y OR2X1_LOC_46/A 0.03fF
C36576 AND2X1_LOC_64/Y AND2X1_LOC_433/a_8_24# 0.04fF
C36577 OR2X1_LOC_22/Y OR2X1_LOC_245/a_8_216# 0.02fF
C36578 AND2X1_LOC_313/a_8_24# AND2X1_LOC_36/Y 0.01fF
C36579 OR2X1_LOC_10/a_36_216# OR2X1_LOC_585/A 0.00fF
C36580 OR2X1_LOC_70/Y AND2X1_LOC_227/Y 0.10fF
C36581 OR2X1_LOC_185/A OR2X1_LOC_398/Y -0.06fF
C36582 OR2X1_LOC_230/a_8_216# OR2X1_LOC_31/Y 0.19fF
C36583 OR2X1_LOC_805/A OR2X1_LOC_723/A 0.03fF
C36584 GATE_479 AND2X1_LOC_223/A 0.10fF
C36585 OR2X1_LOC_43/A OR2X1_LOC_419/a_8_216# 0.01fF
C36586 AND2X1_LOC_425/Y AND2X1_LOC_694/a_8_24# 0.05fF
C36587 AND2X1_LOC_543/Y AND2X1_LOC_552/A 0.09fF
C36588 AND2X1_LOC_309/a_8_24# OR2X1_LOC_335/B 0.02fF
C36589 OR2X1_LOC_19/B OR2X1_LOC_71/Y 0.01fF
C36590 OR2X1_LOC_32/B OR2X1_LOC_72/Y 0.09fF
C36591 AND2X1_LOC_41/A OR2X1_LOC_777/B 0.09fF
C36592 OR2X1_LOC_468/A OR2X1_LOC_388/a_8_216# 0.00fF
C36593 AND2X1_LOC_110/Y OR2X1_LOC_186/a_8_216# 0.01fF
C36594 OR2X1_LOC_45/B OR2X1_LOC_135/Y 0.02fF
C36595 OR2X1_LOC_364/B OR2X1_LOC_357/B 0.75fF
C36596 OR2X1_LOC_47/Y AND2X1_LOC_729/B 0.02fF
C36597 AND2X1_LOC_633/Y OR2X1_LOC_31/Y 0.02fF
C36598 OR2X1_LOC_303/A OR2X1_LOC_308/Y 0.20fF
C36599 AND2X1_LOC_584/a_8_24# AND2X1_LOC_31/Y 0.01fF
C36600 AND2X1_LOC_150/a_8_24# OR2X1_LOC_576/A -0.00fF
C36601 OR2X1_LOC_732/a_8_216# OR2X1_LOC_732/A 0.04fF
C36602 AND2X1_LOC_784/Y AND2X1_LOC_804/A 0.26fF
C36603 OR2X1_LOC_70/Y OR2X1_LOC_813/Y 0.01fF
C36604 OR2X1_LOC_31/Y D_INPUT_0 0.10fF
C36605 AND2X1_LOC_401/Y AND2X1_LOC_36/Y 0.08fF
C36606 AND2X1_LOC_693/a_36_24# AND2X1_LOC_36/Y 0.01fF
C36607 OR2X1_LOC_742/B OR2X1_LOC_551/a_8_216# 0.03fF
C36608 OR2X1_LOC_244/Y OR2X1_LOC_115/B 0.02fF
C36609 OR2X1_LOC_736/Y OR2X1_LOC_549/A 0.07fF
C36610 AND2X1_LOC_12/a_36_24# INPUT_6 0.00fF
C36611 OR2X1_LOC_19/B D_INPUT_1 0.17fF
C36612 OR2X1_LOC_421/A AND2X1_LOC_769/Y 0.01fF
C36613 OR2X1_LOC_40/Y AND2X1_LOC_358/Y 0.00fF
C36614 OR2X1_LOC_117/a_36_216# AND2X1_LOC_243/Y 0.01fF
C36615 AND2X1_LOC_12/Y OR2X1_LOC_561/A 0.01fF
C36616 OR2X1_LOC_563/a_8_216# OR2X1_LOC_562/A 0.02fF
C36617 OR2X1_LOC_160/B AND2X1_LOC_44/Y 3.99fF
C36618 AND2X1_LOC_70/Y OR2X1_LOC_563/A 0.01fF
C36619 AND2X1_LOC_539/Y OR2X1_LOC_744/A 0.16fF
C36620 AND2X1_LOC_725/a_36_24# OR2X1_LOC_428/A 0.00fF
C36621 AND2X1_LOC_91/B AND2X1_LOC_164/a_8_24# 0.03fF
C36622 OR2X1_LOC_539/Y OR2X1_LOC_112/A 0.01fF
C36623 AND2X1_LOC_476/A OR2X1_LOC_75/a_8_216# 0.03fF
C36624 OR2X1_LOC_499/B OR2X1_LOC_140/B 0.00fF
C36625 OR2X1_LOC_333/B OR2X1_LOC_68/B 0.03fF
C36626 OR2X1_LOC_821/Y OR2X1_LOC_822/a_8_216# 0.03fF
C36627 AND2X1_LOC_41/A OR2X1_LOC_831/B 0.03fF
C36628 OR2X1_LOC_188/a_8_216# AND2X1_LOC_41/A -0.02fF
C36629 OR2X1_LOC_95/Y OR2X1_LOC_615/Y 0.11fF
C36630 OR2X1_LOC_599/A AND2X1_LOC_592/a_36_24# 0.00fF
C36631 AND2X1_LOC_649/Y AND2X1_LOC_655/a_8_24# 0.13fF
C36632 OR2X1_LOC_491/Y OR2X1_LOC_437/A 0.01fF
C36633 OR2X1_LOC_863/A OR2X1_LOC_66/A 0.02fF
C36634 OR2X1_LOC_329/B OR2X1_LOC_428/A 0.31fF
C36635 AND2X1_LOC_65/a_8_24# AND2X1_LOC_7/B 0.01fF
C36636 AND2X1_LOC_227/Y OR2X1_LOC_184/Y 0.98fF
C36637 OR2X1_LOC_251/Y OR2X1_LOC_437/A 0.03fF
C36638 AND2X1_LOC_753/B AND2X1_LOC_64/Y 0.07fF
C36639 OR2X1_LOC_49/A OR2X1_LOC_78/B 0.05fF
C36640 OR2X1_LOC_631/B OR2X1_LOC_777/B 0.07fF
C36641 OR2X1_LOC_770/B OR2X1_LOC_78/B 0.00fF
C36642 OR2X1_LOC_828/a_8_216# OR2X1_LOC_828/Y 0.05fF
C36643 OR2X1_LOC_160/B OR2X1_LOC_719/a_8_216# 0.02fF
C36644 OR2X1_LOC_66/A OR2X1_LOC_719/B 0.03fF
C36645 OR2X1_LOC_177/Y OR2X1_LOC_56/A 0.03fF
C36646 OR2X1_LOC_472/a_36_216# OR2X1_LOC_68/B 0.00fF
C36647 AND2X1_LOC_486/Y AND2X1_LOC_564/B 0.07fF
C36648 OR2X1_LOC_744/A AND2X1_LOC_771/B 0.00fF
C36649 AND2X1_LOC_64/Y OR2X1_LOC_405/A 0.11fF
C36650 AND2X1_LOC_706/a_36_24# OR2X1_LOC_744/A 0.00fF
C36651 OR2X1_LOC_508/a_8_216# OR2X1_LOC_244/B 0.40fF
C36652 OR2X1_LOC_78/B OR2X1_LOC_596/A 0.03fF
C36653 AND2X1_LOC_573/A OR2X1_LOC_503/a_8_216# 0.04fF
C36654 OR2X1_LOC_131/A OR2X1_LOC_744/A 0.03fF
C36655 VDD AND2X1_LOC_715/A 0.22fF
C36656 OR2X1_LOC_231/A AND2X1_LOC_7/B 0.13fF
C36657 AND2X1_LOC_729/Y AND2X1_LOC_209/Y 0.01fF
C36658 AND2X1_LOC_738/B OR2X1_LOC_604/A 0.20fF
C36659 AND2X1_LOC_714/B OR2X1_LOC_421/a_8_216# 0.04fF
C36660 OR2X1_LOC_177/a_8_216# OR2X1_LOC_438/Y 0.40fF
C36661 OR2X1_LOC_517/a_8_216# OR2X1_LOC_158/A 0.03fF
C36662 OR2X1_LOC_604/A OR2X1_LOC_56/A 1.48fF
C36663 OR2X1_LOC_158/A OR2X1_LOC_234/Y 0.09fF
C36664 OR2X1_LOC_526/Y OR2X1_LOC_51/Y 0.02fF
C36665 OR2X1_LOC_529/Y OR2X1_LOC_142/Y 0.00fF
C36666 OR2X1_LOC_106/a_8_216# AND2X1_LOC_474/A 0.01fF
C36667 OR2X1_LOC_494/A OR2X1_LOC_18/Y 0.02fF
C36668 OR2X1_LOC_375/A OR2X1_LOC_120/a_8_216# 0.01fF
C36669 OR2X1_LOC_450/B OR2X1_LOC_467/A 0.01fF
C36670 OR2X1_LOC_45/B AND2X1_LOC_520/Y 0.28fF
C36671 AND2X1_LOC_388/Y AND2X1_LOC_512/Y 0.23fF
C36672 OR2X1_LOC_447/a_8_216# AND2X1_LOC_7/B 0.01fF
C36673 AND2X1_LOC_86/Y AND2X1_LOC_44/Y 0.12fF
C36674 OR2X1_LOC_136/Y AND2X1_LOC_138/a_8_24# 0.11fF
C36675 AND2X1_LOC_501/Y AND2X1_LOC_675/Y 0.05fF
C36676 OR2X1_LOC_573/a_8_216# OR2X1_LOC_66/A 0.01fF
C36677 OR2X1_LOC_703/B OR2X1_LOC_175/Y 0.03fF
C36678 OR2X1_LOC_22/Y OR2X1_LOC_589/a_8_216# 0.03fF
C36679 OR2X1_LOC_130/A AND2X1_LOC_7/B 0.17fF
C36680 VDD OR2X1_LOC_755/Y 0.12fF
C36681 OR2X1_LOC_15/a_8_216# OR2X1_LOC_38/a_8_216# 0.47fF
C36682 AND2X1_LOC_675/Y AND2X1_LOC_570/Y 0.16fF
C36683 OR2X1_LOC_40/Y OR2X1_LOC_438/Y 0.16fF
C36684 AND2X1_LOC_228/Y AND2X1_LOC_231/a_36_24# 0.00fF
C36685 OR2X1_LOC_40/Y AND2X1_LOC_865/a_8_24# 0.04fF
C36686 OR2X1_LOC_696/A OR2X1_LOC_387/Y 0.01fF
C36687 AND2X1_LOC_361/a_8_24# OR2X1_LOC_427/A -0.02fF
C36688 AND2X1_LOC_42/B OR2X1_LOC_622/B 0.02fF
C36689 OR2X1_LOC_739/A OR2X1_LOC_355/a_8_216# 0.01fF
C36690 OR2X1_LOC_203/Y OR2X1_LOC_392/B 0.10fF
C36691 AND2X1_LOC_212/A AND2X1_LOC_841/B 0.03fF
C36692 OR2X1_LOC_325/A AND2X1_LOC_323/a_8_24# 0.01fF
C36693 OR2X1_LOC_49/A OR2X1_LOC_375/A 0.14fF
C36694 OR2X1_LOC_139/A OR2X1_LOC_267/a_8_216# 0.02fF
C36695 AND2X1_LOC_456/B AND2X1_LOC_286/a_8_24# 0.18fF
C36696 AND2X1_LOC_555/Y AND2X1_LOC_259/Y 0.05fF
C36697 OR2X1_LOC_204/Y OR2X1_LOC_266/A 0.15fF
C36698 AND2X1_LOC_784/A AND2X1_LOC_794/a_8_24# 0.01fF
C36699 AND2X1_LOC_7/a_8_24# AND2X1_LOC_7/B 0.01fF
C36700 OR2X1_LOC_604/A OR2X1_LOC_426/Y 0.02fF
C36701 OR2X1_LOC_676/Y OR2X1_LOC_623/B 0.07fF
C36702 OR2X1_LOC_154/A OR2X1_LOC_138/A 0.02fF
C36703 OR2X1_LOC_44/Y AND2X1_LOC_214/a_8_24# 0.03fF
C36704 OR2X1_LOC_492/a_8_216# OR2X1_LOC_39/A 0.09fF
C36705 OR2X1_LOC_235/B OR2X1_LOC_632/Y 0.02fF
C36706 OR2X1_LOC_494/Y OR2X1_LOC_92/Y 0.01fF
C36707 OR2X1_LOC_331/A OR2X1_LOC_516/B 0.82fF
C36708 OR2X1_LOC_158/A AND2X1_LOC_161/a_36_24# 0.02fF
C36709 AND2X1_LOC_181/a_36_24# OR2X1_LOC_329/B 0.01fF
C36710 AND2X1_LOC_363/Y OR2X1_LOC_92/Y 0.02fF
C36711 VDD OR2X1_LOC_761/Y 0.12fF
C36712 OR2X1_LOC_256/A OR2X1_LOC_437/A 0.09fF
C36713 AND2X1_LOC_362/B AND2X1_LOC_573/A 0.07fF
C36714 AND2X1_LOC_722/A OR2X1_LOC_59/Y 0.03fF
C36715 OR2X1_LOC_485/A AND2X1_LOC_465/A 0.17fF
C36716 OR2X1_LOC_375/A OR2X1_LOC_596/A 0.07fF
C36717 OR2X1_LOC_185/A OR2X1_LOC_552/B 0.01fF
C36718 AND2X1_LOC_110/Y OR2X1_LOC_506/A 0.03fF
C36719 OR2X1_LOC_40/Y AND2X1_LOC_621/Y 0.10fF
C36720 OR2X1_LOC_622/A OR2X1_LOC_847/A 0.01fF
C36721 AND2X1_LOC_787/a_36_24# OR2X1_LOC_600/A 0.00fF
C36722 OR2X1_LOC_748/A OR2X1_LOC_12/Y 0.09fF
C36723 OR2X1_LOC_219/B AND2X1_LOC_44/Y 0.01fF
C36724 OR2X1_LOC_834/A OR2X1_LOC_623/B 0.03fF
C36725 OR2X1_LOC_671/Y OR2X1_LOC_85/A 0.09fF
C36726 INPUT_3 OR2X1_LOC_600/A 0.03fF
C36727 OR2X1_LOC_553/A OR2X1_LOC_719/a_8_216# 0.03fF
C36728 AND2X1_LOC_716/Y INPUT_0 0.07fF
C36729 OR2X1_LOC_51/Y AND2X1_LOC_805/Y 0.00fF
C36730 AND2X1_LOC_476/A OR2X1_LOC_13/B 0.07fF
C36731 AND2X1_LOC_367/B OR2X1_LOC_427/A 0.04fF
C36732 AND2X1_LOC_732/B AND2X1_LOC_448/Y 0.02fF
C36733 OR2X1_LOC_426/B AND2X1_LOC_662/B 0.02fF
C36734 OR2X1_LOC_470/a_8_216# OR2X1_LOC_467/B 0.01fF
C36735 OR2X1_LOC_389/B OR2X1_LOC_390/A 0.02fF
C36736 AND2X1_LOC_798/a_8_24# OR2X1_LOC_22/Y 0.03fF
C36737 AND2X1_LOC_50/Y OR2X1_LOC_638/a_8_216# 0.01fF
C36738 AND2X1_LOC_705/Y OR2X1_LOC_420/a_8_216# 0.01fF
C36739 VDD AND2X1_LOC_272/a_8_24# 0.00fF
C36740 INPUT_0 AND2X1_LOC_654/Y 0.07fF
C36741 AND2X1_LOC_59/Y OR2X1_LOC_602/Y 0.43fF
C36742 AND2X1_LOC_84/Y OR2X1_LOC_64/Y 0.35fF
C36743 OR2X1_LOC_252/a_8_216# OR2X1_LOC_56/A 0.08fF
C36744 OR2X1_LOC_861/a_36_216# OR2X1_LOC_624/Y 0.03fF
C36745 OR2X1_LOC_158/B OR2X1_LOC_158/Y 0.01fF
C36746 AND2X1_LOC_12/Y OR2X1_LOC_35/Y 0.01fF
C36747 OR2X1_LOC_43/A AND2X1_LOC_194/Y 0.03fF
C36748 AND2X1_LOC_12/Y OR2X1_LOC_359/A 0.01fF
C36749 AND2X1_LOC_31/Y OR2X1_LOC_641/B 0.01fF
C36750 OR2X1_LOC_160/A OR2X1_LOC_78/A 0.40fF
C36751 OR2X1_LOC_117/Y AND2X1_LOC_243/Y 0.02fF
C36752 OR2X1_LOC_190/A OR2X1_LOC_270/a_8_216# 0.07fF
C36753 OR2X1_LOC_335/A OR2X1_LOC_335/B 0.42fF
C36754 AND2X1_LOC_367/A AND2X1_LOC_99/A 0.03fF
C36755 OR2X1_LOC_565/A OR2X1_LOC_564/B 0.18fF
C36756 AND2X1_LOC_772/B AND2X1_LOC_572/A 0.28fF
C36757 AND2X1_LOC_56/B OR2X1_LOC_66/A 0.19fF
C36758 OR2X1_LOC_756/B OR2X1_LOC_181/B 0.02fF
C36759 VDD AND2X1_LOC_348/Y 0.04fF
C36760 OR2X1_LOC_663/a_8_216# OR2X1_LOC_624/B 0.01fF
C36761 OR2X1_LOC_659/B OR2X1_LOC_66/A 0.02fF
C36762 OR2X1_LOC_139/A OR2X1_LOC_476/a_8_216# 0.06fF
C36763 AND2X1_LOC_716/Y AND2X1_LOC_717/Y 0.02fF
C36764 OR2X1_LOC_304/Y OR2X1_LOC_12/Y 0.03fF
C36765 OR2X1_LOC_36/Y AND2X1_LOC_285/Y 0.17fF
C36766 OR2X1_LOC_743/A OR2X1_LOC_421/Y 1.01fF
C36767 AND2X1_LOC_503/a_36_24# OR2X1_LOC_502/A 0.00fF
C36768 OR2X1_LOC_45/B AND2X1_LOC_856/B 1.24fF
C36769 OR2X1_LOC_783/a_8_216# OR2X1_LOC_712/B 0.01fF
C36770 OR2X1_LOC_520/Y AND2X1_LOC_19/Y 1.24fF
C36771 VDD OR2X1_LOC_753/A 6.11fF
C36772 OR2X1_LOC_87/A OR2X1_LOC_803/A 0.03fF
C36773 OR2X1_LOC_45/B AND2X1_LOC_464/Y 0.01fF
C36774 OR2X1_LOC_45/B AND2X1_LOC_863/A 0.00fF
C36775 OR2X1_LOC_448/B AND2X1_LOC_422/a_36_24# 0.00fF
C36776 AND2X1_LOC_8/Y OR2X1_LOC_66/A 0.08fF
C36777 OR2X1_LOC_292/a_8_216# AND2X1_LOC_848/Y 0.02fF
C36778 OR2X1_LOC_715/B OR2X1_LOC_702/A 0.12fF
C36779 OR2X1_LOC_744/A AND2X1_LOC_379/a_36_24# 0.00fF
C36780 AND2X1_LOC_724/A OR2X1_LOC_64/Y 0.02fF
C36781 OR2X1_LOC_626/a_8_216# OR2X1_LOC_627/Y 0.01fF
C36782 OR2X1_LOC_26/Y OR2X1_LOC_585/Y 0.01fF
C36783 OR2X1_LOC_11/Y OR2X1_LOC_762/Y 0.00fF
C36784 AND2X1_LOC_216/Y AND2X1_LOC_116/Y 0.02fF
C36785 OR2X1_LOC_468/A OR2X1_LOC_592/a_36_216# 0.00fF
C36786 OR2X1_LOC_532/B OR2X1_LOC_390/a_8_216# 0.01fF
C36787 OR2X1_LOC_808/A OR2X1_LOC_375/A 0.00fF
C36788 OR2X1_LOC_818/Y AND2X1_LOC_820/a_8_24# 0.23fF
C36789 AND2X1_LOC_468/B OR2X1_LOC_594/Y 0.23fF
C36790 VDD OR2X1_LOC_445/a_8_216# 0.00fF
C36791 AND2X1_LOC_95/Y AND2X1_LOC_125/a_8_24# 0.01fF
C36792 VDD OR2X1_LOC_754/a_8_216# 0.00fF
C36793 OR2X1_LOC_58/a_36_216# OR2X1_LOC_39/A 0.00fF
C36794 OR2X1_LOC_489/B OR2X1_LOC_489/a_8_216# 0.05fF
C36795 OR2X1_LOC_26/a_8_216# OR2X1_LOC_44/Y 0.01fF
C36796 OR2X1_LOC_3/Y OR2X1_LOC_583/Y 0.04fF
C36797 OR2X1_LOC_654/A OR2X1_LOC_35/a_8_216# 0.02fF
C36798 AND2X1_LOC_40/Y AND2X1_LOC_617/a_8_24# 0.01fF
C36799 OR2X1_LOC_528/Y AND2X1_LOC_631/Y 0.16fF
C36800 OR2X1_LOC_427/A OR2X1_LOC_48/B 0.09fF
C36801 OR2X1_LOC_600/a_8_216# OR2X1_LOC_485/A 0.01fF
C36802 OR2X1_LOC_40/Y AND2X1_LOC_650/a_8_24# 0.02fF
C36803 AND2X1_LOC_552/a_8_24# OR2X1_LOC_31/Y 0.02fF
C36804 OR2X1_LOC_220/A OR2X1_LOC_738/A 0.42fF
C36805 AND2X1_LOC_456/B OR2X1_LOC_669/A 0.01fF
C36806 OR2X1_LOC_6/B AND2X1_LOC_117/a_36_24# 0.01fF
C36807 OR2X1_LOC_18/Y OR2X1_LOC_427/A 0.46fF
C36808 AND2X1_LOC_850/a_8_24# AND2X1_LOC_850/Y -0.05fF
C36809 OR2X1_LOC_95/Y AND2X1_LOC_242/B 0.24fF
C36810 OR2X1_LOC_244/A AND2X1_LOC_44/Y 0.14fF
C36811 AND2X1_LOC_687/Y OR2X1_LOC_16/A 0.01fF
C36812 OR2X1_LOC_757/A AND2X1_LOC_620/a_36_24# 0.00fF
C36813 OR2X1_LOC_656/B OR2X1_LOC_185/A 0.03fF
C36814 OR2X1_LOC_18/Y OR2X1_LOC_63/a_8_216# 0.01fF
C36815 OR2X1_LOC_231/A OR2X1_LOC_805/A 0.03fF
C36816 AND2X1_LOC_753/a_8_24# AND2X1_LOC_43/B 0.05fF
C36817 OR2X1_LOC_781/B OR2X1_LOC_781/Y 0.80fF
C36818 OR2X1_LOC_619/Y AND2X1_LOC_452/Y 0.00fF
C36819 OR2X1_LOC_426/B OR2X1_LOC_273/Y 0.15fF
C36820 AND2X1_LOC_350/B OR2X1_LOC_31/Y 0.03fF
C36821 OR2X1_LOC_95/a_36_216# OR2X1_LOC_586/Y 0.00fF
C36822 OR2X1_LOC_624/B OR2X1_LOC_78/A 0.07fF
C36823 OR2X1_LOC_680/A AND2X1_LOC_805/Y 0.03fF
C36824 OR2X1_LOC_33/B OR2X1_LOC_78/B 0.01fF
C36825 AND2X1_LOC_95/Y OR2X1_LOC_128/a_36_216# 0.00fF
C36826 AND2X1_LOC_593/Y AND2X1_LOC_653/B 0.01fF
C36827 OR2X1_LOC_128/A OR2X1_LOC_128/a_8_216# 0.47fF
C36828 OR2X1_LOC_659/Y AND2X1_LOC_47/Y 0.25fF
C36829 AND2X1_LOC_24/a_36_24# OR2X1_LOC_33/B 0.00fF
C36830 AND2X1_LOC_840/A AND2X1_LOC_840/B 0.49fF
C36831 AND2X1_LOC_736/Y OR2X1_LOC_498/Y 0.82fF
C36832 OR2X1_LOC_631/B OR2X1_LOC_575/A 0.00fF
C36833 VDD OR2X1_LOC_684/Y 0.03fF
C36834 OR2X1_LOC_92/Y OR2X1_LOC_86/a_36_216# 0.00fF
C36835 OR2X1_LOC_18/Y AND2X1_LOC_464/a_8_24# 0.02fF
C36836 OR2X1_LOC_666/A OR2X1_LOC_64/Y 0.05fF
C36837 OR2X1_LOC_31/Y AND2X1_LOC_771/B 0.01fF
C36838 AND2X1_LOC_347/Y AND2X1_LOC_347/a_8_24# 0.06fF
C36839 AND2X1_LOC_41/A AND2X1_LOC_13/a_8_24# 0.04fF
C36840 OR2X1_LOC_271/a_8_216# OR2X1_LOC_18/Y 0.01fF
C36841 OR2X1_LOC_426/B OR2X1_LOC_19/B 0.84fF
C36842 OR2X1_LOC_130/A OR2X1_LOC_805/A 0.14fF
C36843 AND2X1_LOC_717/Y OR2X1_LOC_312/Y 0.03fF
C36844 OR2X1_LOC_808/A OR2X1_LOC_605/B 0.06fF
C36845 OR2X1_LOC_463/B OR2X1_LOC_375/A 0.13fF
C36846 AND2X1_LOC_7/B AND2X1_LOC_39/Y 0.01fF
C36847 OR2X1_LOC_194/Y AND2X1_LOC_43/B 0.08fF
C36848 OR2X1_LOC_160/B OR2X1_LOC_720/B 0.03fF
C36849 AND2X1_LOC_95/Y AND2X1_LOC_472/B 0.37fF
C36850 OR2X1_LOC_70/Y AND2X1_LOC_722/A 0.03fF
C36851 OR2X1_LOC_306/a_8_216# OR2X1_LOC_43/A 0.03fF
C36852 OR2X1_LOC_856/B AND2X1_LOC_3/Y 0.07fF
C36853 AND2X1_LOC_363/A OR2X1_LOC_18/Y 0.16fF
C36854 OR2X1_LOC_756/B AND2X1_LOC_261/a_8_24# 0.19fF
C36855 OR2X1_LOC_385/Y OR2X1_LOC_427/A 0.07fF
C36856 AND2X1_LOC_599/a_36_24# OR2X1_LOC_214/B 0.01fF
C36857 OR2X1_LOC_64/Y OR2X1_LOC_762/Y 0.18fF
C36858 OR2X1_LOC_87/B OR2X1_LOC_375/A 0.06fF
C36859 OR2X1_LOC_256/a_36_216# OR2X1_LOC_585/A 0.00fF
C36860 VDD AND2X1_LOC_845/Y 0.68fF
C36861 OR2X1_LOC_401/B OR2X1_LOC_78/Y 0.01fF
C36862 OR2X1_LOC_401/a_36_216# OR2X1_LOC_78/B 0.00fF
C36863 OR2X1_LOC_91/Y OR2X1_LOC_36/Y 0.03fF
C36864 AND2X1_LOC_658/B OR2X1_LOC_679/A 0.03fF
C36865 OR2X1_LOC_634/A AND2X1_LOC_27/a_8_24# 0.17fF
C36866 OR2X1_LOC_91/Y OR2X1_LOC_91/a_8_216# 0.03fF
C36867 OR2X1_LOC_160/A OR2X1_LOC_155/A 1.05fF
C36868 AND2X1_LOC_593/Y AND2X1_LOC_645/A 0.12fF
C36869 OR2X1_LOC_170/a_8_216# OR2X1_LOC_568/A 0.03fF
C36870 OR2X1_LOC_490/Y AND2X1_LOC_99/A 0.09fF
C36871 OR2X1_LOC_479/Y OR2X1_LOC_620/Y 0.03fF
C36872 OR2X1_LOC_85/A OR2X1_LOC_42/a_8_216# 0.06fF
C36873 OR2X1_LOC_7/A AND2X1_LOC_621/Y 0.11fF
C36874 AND2X1_LOC_110/a_36_24# D_INPUT_0 0.00fF
C36875 AND2X1_LOC_326/B OR2X1_LOC_31/Y 0.01fF
C36876 AND2X1_LOC_722/A AND2X1_LOC_514/Y 0.19fF
C36877 OR2X1_LOC_161/B AND2X1_LOC_418/a_36_24# 0.00fF
C36878 OR2X1_LOC_666/A OR2X1_LOC_417/A 0.24fF
C36879 AND2X1_LOC_612/B OR2X1_LOC_375/A 0.03fF
C36880 AND2X1_LOC_716/Y OR2X1_LOC_64/Y 0.07fF
C36881 OR2X1_LOC_305/Y OR2X1_LOC_36/Y 0.01fF
C36882 OR2X1_LOC_599/A OR2X1_LOC_433/a_8_216# 0.00fF
C36883 OR2X1_LOC_465/B OR2X1_LOC_553/A 0.02fF
C36884 OR2X1_LOC_866/a_36_216# OR2X1_LOC_859/B 0.00fF
C36885 AND2X1_LOC_31/Y OR2X1_LOC_227/A 0.01fF
C36886 OR2X1_LOC_51/Y AND2X1_LOC_810/Y 0.03fF
C36887 OR2X1_LOC_321/Y OR2X1_LOC_619/Y 0.03fF
C36888 AND2X1_LOC_169/a_8_24# AND2X1_LOC_434/Y 0.08fF
C36889 OR2X1_LOC_64/Y AND2X1_LOC_654/Y 0.04fF
C36890 AND2X1_LOC_729/Y AND2X1_LOC_728/a_8_24# 0.01fF
C36891 OR2X1_LOC_3/Y AND2X1_LOC_342/Y 0.04fF
C36892 OR2X1_LOC_19/B AND2X1_LOC_414/a_8_24# 0.01fF
C36893 AND2X1_LOC_866/A OR2X1_LOC_59/Y 0.11fF
C36894 AND2X1_LOC_701/a_8_24# OR2X1_LOC_269/B 0.03fF
C36895 OR2X1_LOC_31/Y AND2X1_LOC_471/Y 0.11fF
C36896 OR2X1_LOC_316/Y OR2X1_LOC_27/a_8_216# 0.01fF
C36897 OR2X1_LOC_224/a_36_216# OR2X1_LOC_56/A 0.00fF
C36898 OR2X1_LOC_251/Y OR2X1_LOC_669/a_36_216# 0.00fF
C36899 AND2X1_LOC_727/A AND2X1_LOC_841/B 0.03fF
C36900 AND2X1_LOC_141/B AND2X1_LOC_572/A 0.11fF
C36901 AND2X1_LOC_602/a_8_24# AND2X1_LOC_645/A 0.00fF
C36902 OR2X1_LOC_264/Y D_INPUT_0 0.00fF
C36903 OR2X1_LOC_137/B OR2X1_LOC_404/Y 0.01fF
C36904 OR2X1_LOC_246/A OR2X1_LOC_278/Y 0.03fF
C36905 D_INPUT_6 INPUT_6 0.72fF
C36906 AND2X1_LOC_502/a_8_24# OR2X1_LOC_64/Y 0.00fF
C36907 AND2X1_LOC_95/Y OR2X1_LOC_19/B 0.05fF
C36908 OR2X1_LOC_600/A AND2X1_LOC_793/Y 0.02fF
C36909 AND2X1_LOC_110/Y OR2X1_LOC_356/a_36_216# 0.00fF
C36910 AND2X1_LOC_716/Y OR2X1_LOC_417/A 0.09fF
C36911 OR2X1_LOC_599/A OR2X1_LOC_70/Y 0.04fF
C36912 AND2X1_LOC_52/a_36_24# AND2X1_LOC_53/Y 0.00fF
C36913 OR2X1_LOC_409/B OR2X1_LOC_763/a_8_216# 0.00fF
C36914 AND2X1_LOC_847/a_8_24# OR2X1_LOC_820/B 0.05fF
C36915 OR2X1_LOC_682/Y OR2X1_LOC_3/Y 0.02fF
C36916 OR2X1_LOC_362/B OR2X1_LOC_814/A 0.00fF
C36917 OR2X1_LOC_600/A AND2X1_LOC_259/a_36_24# 0.00fF
C36918 OR2X1_LOC_709/A OR2X1_LOC_724/A 0.16fF
C36919 AND2X1_LOC_465/Y OR2X1_LOC_39/A 0.02fF
C36920 AND2X1_LOC_40/Y OR2X1_LOC_440/A 0.00fF
C36921 AND2X1_LOC_477/A AND2X1_LOC_593/Y 4.23fF
C36922 OR2X1_LOC_319/a_8_216# OR2X1_LOC_532/B 0.01fF
C36923 OR2X1_LOC_235/B OR2X1_LOC_234/a_8_216# 0.02fF
C36924 OR2X1_LOC_127/a_8_216# INPUT_1 0.07fF
C36925 AND2X1_LOC_650/a_8_24# AND2X1_LOC_857/a_8_24# 0.23fF
C36926 OR2X1_LOC_417/Y OR2X1_LOC_36/Y 0.03fF
C36927 OR2X1_LOC_41/a_8_216# AND2X1_LOC_434/Y 0.04fF
C36928 AND2X1_LOC_840/A OR2X1_LOC_31/Y 0.23fF
C36929 OR2X1_LOC_291/Y OR2X1_LOC_36/Y 0.06fF
C36930 OR2X1_LOC_278/a_8_216# OR2X1_LOC_74/A 0.01fF
C36931 AND2X1_LOC_375/a_8_24# OR2X1_LOC_31/Y 0.08fF
C36932 AND2X1_LOC_576/Y AND2X1_LOC_849/A 0.00fF
C36933 AND2X1_LOC_841/B OR2X1_LOC_95/Y 0.03fF
C36934 OR2X1_LOC_45/B OR2X1_LOC_300/a_36_216# 0.00fF
C36935 AND2X1_LOC_59/Y OR2X1_LOC_602/B 0.01fF
C36936 OR2X1_LOC_311/Y OR2X1_LOC_36/Y 0.03fF
C36937 OR2X1_LOC_377/A OR2X1_LOC_532/B 0.54fF
C36938 AND2X1_LOC_18/Y OR2X1_LOC_228/Y 0.09fF
C36939 OR2X1_LOC_46/A OR2X1_LOC_461/A 0.65fF
C36940 OR2X1_LOC_312/Y OR2X1_LOC_64/Y 0.03fF
C36941 OR2X1_LOC_743/A OR2X1_LOC_273/Y 0.27fF
C36942 OR2X1_LOC_541/A OR2X1_LOC_493/Y 0.23fF
C36943 OR2X1_LOC_802/Y OR2X1_LOC_814/A 0.04fF
C36944 OR2X1_LOC_148/B OR2X1_LOC_148/A 0.16fF
C36945 OR2X1_LOC_271/Y AND2X1_LOC_116/B 0.00fF
C36946 AND2X1_LOC_784/A AND2X1_LOC_326/a_8_24# 0.03fF
C36947 AND2X1_LOC_47/Y AND2X1_LOC_601/a_8_24# 0.01fF
C36948 OR2X1_LOC_250/Y D_INPUT_3 0.23fF
C36949 AND2X1_LOC_550/A AND2X1_LOC_796/Y 0.11fF
C36950 AND2X1_LOC_866/B AND2X1_LOC_792/Y 0.06fF
C36951 OR2X1_LOC_2/Y OR2X1_LOC_51/B 0.03fF
C36952 AND2X1_LOC_2/Y AND2X1_LOC_31/Y 0.04fF
C36953 AND2X1_LOC_31/Y OR2X1_LOC_702/a_8_216# 0.06fF
C36954 OR2X1_LOC_458/B OR2X1_LOC_717/a_8_216# 0.01fF
C36955 AND2X1_LOC_372/a_36_24# OR2X1_LOC_493/Y 0.00fF
C36956 OR2X1_LOC_532/B OR2X1_LOC_203/Y 0.07fF
C36957 OR2X1_LOC_643/A D_INPUT_0 0.07fF
C36958 OR2X1_LOC_46/A OR2X1_LOC_240/A 0.03fF
C36959 OR2X1_LOC_40/Y OR2X1_LOC_71/A 0.06fF
C36960 AND2X1_LOC_772/B AND2X1_LOC_772/a_8_24# 0.00fF
C36961 OR2X1_LOC_680/A AND2X1_LOC_810/Y 0.08fF
C36962 OR2X1_LOC_624/A OR2X1_LOC_223/A 0.07fF
C36963 OR2X1_LOC_95/a_8_216# OR2X1_LOC_409/B 0.00fF
C36964 OR2X1_LOC_11/Y OR2X1_LOC_409/a_8_216# 0.01fF
C36965 OR2X1_LOC_3/Y AND2X1_LOC_712/B 0.39fF
C36966 D_INPUT_0 OR2X1_LOC_124/Y 0.04fF
C36967 AND2X1_LOC_67/Y AND2X1_LOC_51/Y 0.02fF
C36968 OR2X1_LOC_319/B OR2X1_LOC_365/B 0.00fF
C36969 OR2X1_LOC_596/A OR2X1_LOC_515/Y 0.13fF
C36970 OR2X1_LOC_3/Y OR2X1_LOC_54/Y 0.02fF
C36971 OR2X1_LOC_472/A D_INPUT_0 0.03fF
C36972 OR2X1_LOC_840/A OR2X1_LOC_318/B 0.03fF
C36973 OR2X1_LOC_256/A OR2X1_LOC_753/A 0.09fF
C36974 AND2X1_LOC_839/A OR2X1_LOC_585/A 0.01fF
C36975 OR2X1_LOC_48/Y OR2X1_LOC_7/a_8_216# 0.39fF
C36976 OR2X1_LOC_296/Y OR2X1_LOC_62/B 0.37fF
C36977 OR2X1_LOC_759/a_8_216# OR2X1_LOC_759/Y 0.03fF
C36978 AND2X1_LOC_318/Y OR2X1_LOC_6/A 0.01fF
C36979 OR2X1_LOC_312/Y OR2X1_LOC_417/A 0.10fF
C36980 D_INPUT_3 OR2X1_LOC_36/Y 0.00fF
C36981 OR2X1_LOC_273/Y OR2X1_LOC_246/A 0.01fF
C36982 OR2X1_LOC_840/A OR2X1_LOC_854/A 0.05fF
C36983 AND2X1_LOC_776/Y AND2X1_LOC_721/Y 0.01fF
C36984 OR2X1_LOC_846/B OR2X1_LOC_814/A 0.00fF
C36985 OR2X1_LOC_817/Y INPUT_1 0.01fF
C36986 OR2X1_LOC_65/B AND2X1_LOC_204/Y 0.00fF
C36987 OR2X1_LOC_696/A AND2X1_LOC_705/Y 0.10fF
C36988 OR2X1_LOC_121/B OR2X1_LOC_606/a_8_216# 0.00fF
C36989 OR2X1_LOC_696/A AND2X1_LOC_809/a_36_24# 0.00fF
C36990 AND2X1_LOC_8/Y OR2X1_LOC_84/A 0.03fF
C36991 D_INPUT_3 OR2X1_LOC_93/a_36_216# 0.00fF
C36992 AND2X1_LOC_564/A OR2X1_LOC_406/Y 0.32fF
C36993 AND2X1_LOC_191/Y AND2X1_LOC_866/A 0.11fF
C36994 OR2X1_LOC_375/A OR2X1_LOC_374/Y 0.06fF
C36995 OR2X1_LOC_19/B OR2X1_LOC_246/A 0.07fF
C36996 OR2X1_LOC_97/A OR2X1_LOC_390/a_36_216# -0.00fF
C36997 OR2X1_LOC_620/B OR2X1_LOC_620/A 0.11fF
C36998 AND2X1_LOC_339/a_36_24# AND2X1_LOC_476/A 0.00fF
C36999 AND2X1_LOC_670/a_8_24# OR2X1_LOC_532/B 0.03fF
C37000 OR2X1_LOC_648/A OR2X1_LOC_777/B 0.03fF
C37001 OR2X1_LOC_91/Y OR2X1_LOC_419/Y 0.10fF
C37002 INPUT_0 OR2X1_LOC_13/B 0.50fF
C37003 AND2X1_LOC_711/Y AND2X1_LOC_866/A 0.19fF
C37004 OR2X1_LOC_121/Y OR2X1_LOC_115/B 0.00fF
C37005 OR2X1_LOC_650/Y AND2X1_LOC_519/a_8_24# 0.25fF
C37006 AND2X1_LOC_304/a_36_24# OR2X1_LOC_446/B 0.01fF
C37007 AND2X1_LOC_22/Y AND2X1_LOC_604/a_8_24# 0.01fF
C37008 OR2X1_LOC_391/B OR2X1_LOC_774/B 0.23fF
C37009 OR2X1_LOC_481/A OR2X1_LOC_55/a_36_216# 0.00fF
C37010 AND2X1_LOC_715/Y AND2X1_LOC_809/a_36_24# 0.00fF
C37011 OR2X1_LOC_260/Y OR2X1_LOC_345/a_8_216# 0.01fF
C37012 OR2X1_LOC_576/A OR2X1_LOC_161/B 0.01fF
C37013 AND2X1_LOC_629/Y AND2X1_LOC_632/A 0.00fF
C37014 OR2X1_LOC_494/A AND2X1_LOC_363/a_8_24# 0.01fF
C37015 OR2X1_LOC_655/B OR2X1_LOC_814/A 0.42fF
C37016 AND2X1_LOC_687/A OR2X1_LOC_31/Y 0.11fF
C37017 AND2X1_LOC_469/Y AND2X1_LOC_220/B 0.01fF
C37018 AND2X1_LOC_486/Y OR2X1_LOC_437/A 0.16fF
C37019 OR2X1_LOC_857/B OR2X1_LOC_853/a_8_216# 0.04fF
C37020 AND2X1_LOC_12/Y OR2X1_LOC_80/A 0.75fF
C37021 AND2X1_LOC_514/Y AND2X1_LOC_866/A 0.03fF
C37022 AND2X1_LOC_277/a_8_24# OR2X1_LOC_633/A 0.04fF
C37023 OR2X1_LOC_316/a_36_216# OR2X1_LOC_58/Y 0.00fF
C37024 OR2X1_LOC_114/B OR2X1_LOC_115/B 0.02fF
C37025 OR2X1_LOC_244/A OR2X1_LOC_720/B 0.07fF
C37026 OR2X1_LOC_154/A OR2X1_LOC_68/B 0.31fF
C37027 AND2X1_LOC_191/B AND2X1_LOC_792/a_8_24# 0.05fF
C37028 AND2X1_LOC_31/Y AND2X1_LOC_298/a_8_24# 0.10fF
C37029 OR2X1_LOC_328/a_8_216# OR2X1_LOC_387/A 0.40fF
C37030 AND2X1_LOC_18/Y OR2X1_LOC_562/A 0.02fF
C37031 OR2X1_LOC_39/A OR2X1_LOC_521/a_36_216# 0.00fF
C37032 OR2X1_LOC_864/A OR2X1_LOC_641/B 0.01fF
C37033 OR2X1_LOC_391/B OR2X1_LOC_557/a_8_216# 0.02fF
C37034 OR2X1_LOC_69/a_8_216# AND2X1_LOC_206/Y 0.47fF
C37035 OR2X1_LOC_751/Y AND2X1_LOC_789/Y 0.81fF
C37036 AND2X1_LOC_47/Y AND2X1_LOC_7/Y 0.01fF
C37037 OR2X1_LOC_256/A AND2X1_LOC_845/Y 0.14fF
C37038 OR2X1_LOC_673/A OR2X1_LOC_54/Y 0.05fF
C37039 OR2X1_LOC_439/B OR2X1_LOC_161/B 0.01fF
C37040 AND2X1_LOC_31/Y OR2X1_LOC_269/B 0.73fF
C37041 OR2X1_LOC_666/A OR2X1_LOC_89/a_36_216# 0.00fF
C37042 AND2X1_LOC_91/B OR2X1_LOC_862/B 0.22fF
C37043 OR2X1_LOC_175/Y OR2X1_LOC_389/A 0.22fF
C37044 OR2X1_LOC_354/A OR2X1_LOC_703/Y 0.02fF
C37045 AND2X1_LOC_64/Y AND2X1_LOC_19/Y 0.07fF
C37046 OR2X1_LOC_47/Y OR2X1_LOC_46/A 0.26fF
C37047 OR2X1_LOC_87/A OR2X1_LOC_546/A 0.03fF
C37048 OR2X1_LOC_198/a_8_216# AND2X1_LOC_41/A 0.05fF
C37049 OR2X1_LOC_663/a_36_216# OR2X1_LOC_113/B 0.00fF
C37050 OR2X1_LOC_755/A AND2X1_LOC_846/a_8_24# 0.01fF
C37051 AND2X1_LOC_664/a_8_24# AND2X1_LOC_792/Y 0.03fF
C37052 OR2X1_LOC_74/A OR2X1_LOC_72/Y 0.07fF
C37053 AND2X1_LOC_539/a_36_24# OR2X1_LOC_12/Y 0.00fF
C37054 AND2X1_LOC_716/a_8_24# OR2X1_LOC_437/A 0.12fF
C37055 AND2X1_LOC_461/a_8_24# OR2X1_LOC_46/A 0.01fF
C37056 OR2X1_LOC_131/Y OR2X1_LOC_88/Y 0.00fF
C37057 OR2X1_LOC_696/A AND2X1_LOC_553/A 0.02fF
C37058 OR2X1_LOC_691/Y OR2X1_LOC_801/a_8_216# 0.01fF
C37059 OR2X1_LOC_821/Y OR2X1_LOC_813/a_8_216# 0.03fF
C37060 OR2X1_LOC_196/Y OR2X1_LOC_78/A 0.01fF
C37061 AND2X1_LOC_133/a_8_24# OR2X1_LOC_84/Y 0.24fF
C37062 VDD OR2X1_LOC_323/Y 0.44fF
C37063 AND2X1_LOC_64/Y AND2X1_LOC_316/a_8_24# 0.01fF
C37064 OR2X1_LOC_248/Y OR2X1_LOC_437/A 0.36fF
C37065 AND2X1_LOC_227/Y OR2X1_LOC_47/Y 0.02fF
C37066 OR2X1_LOC_778/A OR2X1_LOC_68/B 0.14fF
C37067 AND2X1_LOC_738/B OR2X1_LOC_533/Y 0.04fF
C37068 OR2X1_LOC_215/A AND2X1_LOC_31/Y 0.38fF
C37069 AND2X1_LOC_550/a_8_24# AND2X1_LOC_476/Y 0.03fF
C37070 AND2X1_LOC_565/B AND2X1_LOC_475/Y 0.31fF
C37071 OR2X1_LOC_741/Y OR2X1_LOC_486/Y 0.03fF
C37072 OR2X1_LOC_687/a_8_216# AND2X1_LOC_430/B 0.01fF
C37073 OR2X1_LOC_56/A AND2X1_LOC_212/Y 0.14fF
C37074 AND2X1_LOC_64/Y AND2X1_LOC_423/a_36_24# 0.00fF
C37075 OR2X1_LOC_744/A AND2X1_LOC_771/a_36_24# 0.00fF
C37076 AND2X1_LOC_212/A AND2X1_LOC_337/a_8_24# 0.01fF
C37077 OR2X1_LOC_516/Y OR2X1_LOC_39/A 1.95fF
C37078 AND2X1_LOC_714/B OR2X1_LOC_51/Y 0.01fF
C37079 OR2X1_LOC_392/B OR2X1_LOC_721/Y 0.10fF
C37080 OR2X1_LOC_45/B AND2X1_LOC_160/a_8_24# 0.01fF
C37081 AND2X1_LOC_348/a_8_24# OR2X1_LOC_384/Y 0.02fF
C37082 AND2X1_LOC_392/A AND2X1_LOC_352/a_36_24# 0.01fF
C37083 AND2X1_LOC_91/B OR2X1_LOC_788/a_36_216# 0.01fF
C37084 AND2X1_LOC_41/A OR2X1_LOC_161/B 0.81fF
C37085 AND2X1_LOC_566/B AND2X1_LOC_352/B 0.01fF
C37086 OR2X1_LOC_375/A OR2X1_LOC_130/a_36_216# 0.00fF
C37087 OR2X1_LOC_123/a_8_216# OR2X1_LOC_6/B 0.04fF
C37088 AND2X1_LOC_199/A INPUT_0 0.03fF
C37089 AND2X1_LOC_547/Y VDD 0.01fF
C37090 OR2X1_LOC_175/Y AND2X1_LOC_57/a_36_24# 0.01fF
C37091 AND2X1_LOC_352/a_8_24# OR2X1_LOC_56/A 0.01fF
C37092 AND2X1_LOC_70/Y OR2X1_LOC_631/A 0.01fF
C37093 OR2X1_LOC_604/A AND2X1_LOC_285/Y 0.03fF
C37094 OR2X1_LOC_97/A OR2X1_LOC_61/B -0.00fF
C37095 OR2X1_LOC_696/A OR2X1_LOC_511/Y 0.07fF
C37096 AND2X1_LOC_363/a_36_24# OR2X1_LOC_91/A 0.00fF
C37097 AND2X1_LOC_362/B AND2X1_LOC_362/a_8_24# -0.01fF
C37098 AND2X1_LOC_12/Y OR2X1_LOC_115/B 0.37fF
C37099 OR2X1_LOC_859/A OR2X1_LOC_561/B 0.08fF
C37100 AND2X1_LOC_353/a_36_24# OR2X1_LOC_56/A 0.00fF
C37101 OR2X1_LOC_190/A OR2X1_LOC_542/B 3.53fF
C37102 OR2X1_LOC_92/Y AND2X1_LOC_802/Y 0.03fF
C37103 OR2X1_LOC_40/Y OR2X1_LOC_59/Y 0.21fF
C37104 OR2X1_LOC_426/A OR2X1_LOC_16/A 0.33fF
C37105 OR2X1_LOC_161/A OR2X1_LOC_259/A 0.03fF
C37106 AND2X1_LOC_53/Y OR2X1_LOC_513/a_8_216# 0.01fF
C37107 OR2X1_LOC_303/A AND2X1_LOC_110/Y 0.01fF
C37108 AND2X1_LOC_92/Y OR2X1_LOC_66/A 0.09fF
C37109 OR2X1_LOC_557/A AND2X1_LOC_36/Y 0.02fF
C37110 OR2X1_LOC_64/Y OR2X1_LOC_13/B 1.86fF
C37111 OR2X1_LOC_841/A AND2X1_LOC_92/Y 0.04fF
C37112 AND2X1_LOC_64/Y OR2X1_LOC_673/Y 0.07fF
C37113 AND2X1_LOC_422/a_8_24# OR2X1_LOC_713/A 0.04fF
C37114 OR2X1_LOC_516/Y OR2X1_LOC_239/a_36_216# 0.01fF
C37115 OR2X1_LOC_375/A OR2X1_LOC_392/B 0.03fF
C37116 OR2X1_LOC_151/A OR2X1_LOC_574/a_8_216# 0.05fF
C37117 AND2X1_LOC_809/A AND2X1_LOC_809/a_8_24# 0.19fF
C37118 OR2X1_LOC_186/Y OR2X1_LOC_547/B 0.09fF
C37119 OR2X1_LOC_47/Y OR2X1_LOC_753/Y 0.04fF
C37120 OR2X1_LOC_598/Y OR2X1_LOC_637/A 0.26fF
C37121 OR2X1_LOC_243/a_36_216# OR2X1_LOC_71/A 0.00fF
C37122 AND2X1_LOC_98/a_8_24# AND2X1_LOC_98/Y 0.00fF
C37123 VDD AND2X1_LOC_551/B 0.23fF
C37124 AND2X1_LOC_319/A OR2X1_LOC_312/a_8_216# 0.18fF
C37125 OR2X1_LOC_405/A OR2X1_LOC_185/a_8_216# 0.06fF
C37126 AND2X1_LOC_95/Y AND2X1_LOC_534/a_8_24# 0.04fF
C37127 AND2X1_LOC_214/A OR2X1_LOC_51/Y 0.02fF
C37128 OR2X1_LOC_97/A AND2X1_LOC_291/a_8_24# 0.01fF
C37129 OR2X1_LOC_51/Y AND2X1_LOC_861/B 0.02fF
C37130 AND2X1_LOC_318/a_8_24# AND2X1_LOC_786/Y 0.05fF
C37131 OR2X1_LOC_158/A AND2X1_LOC_520/Y 0.02fF
C37132 OR2X1_LOC_9/Y AND2X1_LOC_62/a_8_24# 0.25fF
C37133 OR2X1_LOC_315/Y OR2X1_LOC_323/Y 0.08fF
C37134 OR2X1_LOC_203/a_8_216# OR2X1_LOC_344/A 0.01fF
C37135 AND2X1_LOC_570/Y AND2X1_LOC_456/B 0.00fF
C37136 OR2X1_LOC_696/A AND2X1_LOC_345/Y 0.00fF
C37137 OR2X1_LOC_449/B AND2X1_LOC_7/B 0.07fF
C37138 OR2X1_LOC_715/B OR2X1_LOC_623/a_8_216# 0.28fF
C37139 OR2X1_LOC_800/a_8_216# OR2X1_LOC_691/Y 0.01fF
C37140 OR2X1_LOC_52/B AND2X1_LOC_794/a_8_24# 0.03fF
C37141 AND2X1_LOC_512/Y OR2X1_LOC_329/B 0.07fF
C37142 OR2X1_LOC_417/A OR2X1_LOC_13/B 0.14fF
C37143 AND2X1_LOC_6/a_8_24# OR2X1_LOC_68/B 0.14fF
C37144 AND2X1_LOC_212/A AND2X1_LOC_365/A 0.12fF
C37145 AND2X1_LOC_47/Y OR2X1_LOC_515/a_8_216# 0.02fF
C37146 OR2X1_LOC_91/Y OR2X1_LOC_177/Y 0.04fF
C37147 OR2X1_LOC_656/Y AND2X1_LOC_19/Y 0.01fF
C37148 OR2X1_LOC_318/Y OR2X1_LOC_468/A 0.03fF
C37149 OR2X1_LOC_333/B OR2X1_LOC_174/a_8_216# 0.03fF
C37150 OR2X1_LOC_158/A AND2X1_LOC_848/Y 0.06fF
C37151 AND2X1_LOC_357/B OR2X1_LOC_619/Y 0.02fF
C37152 AND2X1_LOC_743/a_8_24# OR2X1_LOC_155/A 0.01fF
C37153 OR2X1_LOC_186/Y OR2X1_LOC_185/Y 0.06fF
C37154 OR2X1_LOC_91/Y OR2X1_LOC_315/a_8_216# 0.08fF
C37155 AND2X1_LOC_95/Y AND2X1_LOC_110/Y 0.07fF
C37156 OR2X1_LOC_631/B OR2X1_LOC_161/B 0.43fF
C37157 OR2X1_LOC_516/A AND2X1_LOC_477/Y 0.83fF
C37158 OR2X1_LOC_769/A OR2X1_LOC_637/B 0.32fF
C37159 OR2X1_LOC_100/Y OR2X1_LOC_78/B 0.04fF
C37160 OR2X1_LOC_280/a_8_216# OR2X1_LOC_428/A 0.01fF
C37161 OR2X1_LOC_641/a_8_216# OR2X1_LOC_185/A 0.01fF
C37162 OR2X1_LOC_158/A AND2X1_LOC_154/a_36_24# 0.00fF
C37163 OR2X1_LOC_840/A OR2X1_LOC_538/A 0.03fF
C37164 AND2X1_LOC_732/a_8_24# OR2X1_LOC_48/B 0.01fF
C37165 OR2X1_LOC_111/a_8_216# OR2X1_LOC_64/Y 0.01fF
C37166 AND2X1_LOC_181/Y OR2X1_LOC_271/a_8_216# 0.06fF
C37167 OR2X1_LOC_188/Y OR2X1_LOC_455/A 0.01fF
C37168 OR2X1_LOC_532/B OR2X1_LOC_539/B 0.16fF
C37169 OR2X1_LOC_743/A OR2X1_LOC_744/a_8_216# 0.01fF
C37170 AND2X1_LOC_784/A AND2X1_LOC_794/B 0.01fF
C37171 AND2X1_LOC_634/a_36_24# AND2X1_LOC_219/A 0.01fF
C37172 AND2X1_LOC_595/a_8_24# OR2X1_LOC_154/A 0.04fF
C37173 AND2X1_LOC_166/a_8_24# OR2X1_LOC_66/A 0.03fF
C37174 AND2X1_LOC_843/Y OR2X1_LOC_59/Y 0.02fF
C37175 OR2X1_LOC_770/B OR2X1_LOC_401/Y 0.86fF
C37176 OR2X1_LOC_10/a_36_216# OR2X1_LOC_437/A 0.00fF
C37177 VDD OR2X1_LOC_448/Y 0.24fF
C37178 OR2X1_LOC_485/A OR2X1_LOC_522/a_8_216# 0.07fF
C37179 AND2X1_LOC_363/a_8_24# AND2X1_LOC_363/A 0.03fF
C37180 AND2X1_LOC_729/Y VDD 0.91fF
C37181 OR2X1_LOC_757/A AND2X1_LOC_805/Y 0.01fF
C37182 OR2X1_LOC_91/Y OR2X1_LOC_604/A 0.10fF
C37183 OR2X1_LOC_847/A OR2X1_LOC_78/A 0.03fF
C37184 OR2X1_LOC_681/a_8_216# AND2X1_LOC_319/A 0.06fF
C37185 OR2X1_LOC_831/A OR2X1_LOC_778/Y 0.05fF
C37186 OR2X1_LOC_315/a_8_216# OR2X1_LOC_371/a_8_216# 0.47fF
C37187 AND2X1_LOC_16/a_36_24# OR2X1_LOC_78/B 0.02fF
C37188 OR2X1_LOC_551/B OR2X1_LOC_365/a_8_216# 0.03fF
C37189 AND2X1_LOC_40/Y OR2X1_LOC_637/A 0.00fF
C37190 OR2X1_LOC_264/Y AND2X1_LOC_40/Y 0.18fF
C37191 AND2X1_LOC_40/Y OR2X1_LOC_436/B 0.01fF
C37192 OR2X1_LOC_36/Y AND2X1_LOC_254/a_36_24# 0.00fF
C37193 OR2X1_LOC_597/A OR2X1_LOC_44/Y 0.01fF
C37194 OR2X1_LOC_786/Y OR2X1_LOC_217/A 0.02fF
C37195 OR2X1_LOC_860/a_36_216# OR2X1_LOC_756/B 0.00fF
C37196 OR2X1_LOC_121/B AND2X1_LOC_7/B 0.16fF
C37197 OR2X1_LOC_8/Y AND2X1_LOC_852/a_8_24# 0.01fF
C37198 AND2X1_LOC_589/a_36_24# OR2X1_LOC_435/A 0.00fF
C37199 AND2X1_LOC_536/a_8_24# AND2X1_LOC_41/A 0.08fF
C37200 OR2X1_LOC_316/Y AND2X1_LOC_219/Y 0.10fF
C37201 AND2X1_LOC_362/a_36_24# OR2X1_LOC_18/Y 0.00fF
C37202 OR2X1_LOC_405/A OR2X1_LOC_756/B 0.05fF
C37203 OR2X1_LOC_177/a_8_216# OR2X1_LOC_70/Y 0.01fF
C37204 AND2X1_LOC_135/a_8_24# OR2X1_LOC_161/B 0.01fF
C37205 OR2X1_LOC_633/B OR2X1_LOC_786/a_8_216# 0.01fF
C37206 OR2X1_LOC_604/A AND2X1_LOC_446/a_8_24# 0.02fF
C37207 AND2X1_LOC_784/A VDD 0.88fF
C37208 AND2X1_LOC_658/B OR2X1_LOC_599/A 0.03fF
C37209 OR2X1_LOC_518/a_8_216# OR2X1_LOC_31/Y 0.01fF
C37210 AND2X1_LOC_22/Y OR2X1_LOC_19/B 0.19fF
C37211 OR2X1_LOC_111/a_8_216# OR2X1_LOC_417/A 0.02fF
C37212 AND2X1_LOC_849/A AND2X1_LOC_244/A 0.28fF
C37213 OR2X1_LOC_147/A OR2X1_LOC_375/A 0.01fF
C37214 OR2X1_LOC_126/a_8_216# OR2X1_LOC_6/B 0.03fF
C37215 OR2X1_LOC_685/A OR2X1_LOC_78/B 0.01fF
C37216 OR2X1_LOC_316/a_8_216# OR2X1_LOC_31/Y 0.01fF
C37217 OR2X1_LOC_178/Y OR2X1_LOC_44/Y 0.03fF
C37218 OR2X1_LOC_45/Y AND2X1_LOC_654/B 0.14fF
C37219 AND2X1_LOC_842/a_8_24# OR2X1_LOC_39/A 0.17fF
C37220 OR2X1_LOC_3/Y OR2X1_LOC_765/Y 0.03fF
C37221 AND2X1_LOC_191/Y OR2X1_LOC_40/Y 0.09fF
C37222 AND2X1_LOC_94/Y AND2X1_LOC_56/B 0.07fF
C37223 OR2X1_LOC_502/A OR2X1_LOC_624/A 0.10fF
C37224 AND2X1_LOC_191/B AND2X1_LOC_620/a_8_24# 0.01fF
C37225 OR2X1_LOC_680/A AND2X1_LOC_861/B 0.07fF
C37226 AND2X1_LOC_729/Y OR2X1_LOC_677/Y 0.02fF
C37227 AND2X1_LOC_12/Y OR2X1_LOC_840/A 0.06fF
C37228 OR2X1_LOC_185/A OR2X1_LOC_785/B 0.31fF
C37229 OR2X1_LOC_40/Y AND2X1_LOC_711/Y 0.03fF
C37230 OR2X1_LOC_696/A AND2X1_LOC_648/B 0.01fF
C37231 AND2X1_LOC_543/Y OR2X1_LOC_95/Y 0.26fF
C37232 OR2X1_LOC_51/Y AND2X1_LOC_645/A 0.00fF
C37233 AND2X1_LOC_48/A OR2X1_LOC_389/a_8_216# 0.02fF
C37234 AND2X1_LOC_32/a_8_24# OR2X1_LOC_334/B 0.00fF
C37235 OR2X1_LOC_482/Y AND2X1_LOC_830/a_8_24# 0.06fF
C37236 AND2X1_LOC_347/B OR2X1_LOC_481/A 0.00fF
C37237 AND2X1_LOC_81/B OR2X1_LOC_663/A 0.03fF
C37238 OR2X1_LOC_40/Y OR2X1_LOC_70/Y 0.30fF
C37239 OR2X1_LOC_369/Y AND2X1_LOC_211/B 0.10fF
C37240 OR2X1_LOC_653/Y OR2X1_LOC_661/a_8_216# 0.03fF
C37241 AND2X1_LOC_866/B AND2X1_LOC_807/Y 0.03fF
C37242 AND2X1_LOC_543/Y OR2X1_LOC_368/A 0.00fF
C37243 AND2X1_LOC_339/Y INPUT_1 0.01fF
C37244 VDD OR2X1_LOC_3/a_8_216# 0.00fF
C37245 VDD OR2X1_LOC_592/A -0.00fF
C37246 AND2X1_LOC_658/A OR2X1_LOC_239/Y 0.03fF
C37247 OR2X1_LOC_22/A OR2X1_LOC_36/a_8_216# 0.18fF
C37248 AND2X1_LOC_51/Y AND2X1_LOC_625/a_8_24# 0.02fF
C37249 OR2X1_LOC_7/A OR2X1_LOC_59/Y 0.56fF
C37250 AND2X1_LOC_81/B AND2X1_LOC_503/a_8_24# 0.01fF
C37251 VDD OR2X1_LOC_481/Y 0.05fF
C37252 OR2X1_LOC_256/Y OR2X1_LOC_44/Y 0.07fF
C37253 AND2X1_LOC_391/Y OR2X1_LOC_485/A 0.03fF
C37254 OR2X1_LOC_70/Y AND2X1_LOC_535/a_8_24# 0.01fF
C37255 OR2X1_LOC_147/B OR2X1_LOC_457/B 0.03fF
C37256 OR2X1_LOC_485/A AND2X1_LOC_858/B 0.15fF
C37257 OR2X1_LOC_604/A OR2X1_LOC_417/Y 0.09fF
C37258 OR2X1_LOC_426/B OR2X1_LOC_275/A 0.03fF
C37259 OR2X1_LOC_485/A OR2X1_LOC_91/A 0.06fF
C37260 AND2X1_LOC_390/B AND2X1_LOC_434/Y 0.01fF
C37261 OR2X1_LOC_40/Y AND2X1_LOC_514/Y 0.08fF
C37262 OR2X1_LOC_624/A AND2X1_LOC_230/a_8_24# 0.11fF
C37263 OR2X1_LOC_319/B OR2X1_LOC_449/B 0.07fF
C37264 AND2X1_LOC_47/Y OR2X1_LOC_706/a_8_216# 0.03fF
C37265 OR2X1_LOC_851/B OR2X1_LOC_814/A 0.01fF
C37266 AND2X1_LOC_641/a_36_24# AND2X1_LOC_650/Y 0.01fF
C37267 OR2X1_LOC_759/A OR2X1_LOC_665/a_36_216# 0.00fF
C37268 AND2X1_LOC_95/Y OR2X1_LOC_664/Y 0.03fF
C37269 AND2X1_LOC_40/Y OR2X1_LOC_778/Y 0.07fF
C37270 AND2X1_LOC_725/a_36_24# AND2X1_LOC_712/B 0.00fF
C37271 AND2X1_LOC_527/a_8_24# OR2X1_LOC_87/A 0.03fF
C37272 AND2X1_LOC_348/a_8_24# OR2X1_LOC_91/A 0.07fF
C37273 OR2X1_LOC_318/Y OR2X1_LOC_449/B 0.08fF
C37274 OR2X1_LOC_687/Y OR2X1_LOC_185/A 0.14fF
C37275 AND2X1_LOC_535/a_36_24# OR2X1_LOC_417/Y 0.01fF
C37276 OR2X1_LOC_604/A OR2X1_LOC_601/a_8_216# 0.01fF
C37277 AND2X1_LOC_50/Y AND2X1_LOC_21/Y 0.54fF
C37278 OR2X1_LOC_406/a_8_216# AND2X1_LOC_624/A 0.05fF
C37279 OR2X1_LOC_121/Y OR2X1_LOC_241/Y 0.03fF
C37280 AND2X1_LOC_62/a_8_24# AND2X1_LOC_852/Y 0.20fF
C37281 OR2X1_LOC_6/B OR2X1_LOC_611/Y 0.01fF
C37282 AND2X1_LOC_12/Y OR2X1_LOC_222/A 0.13fF
C37283 OR2X1_LOC_404/Y OR2X1_LOC_632/Y 0.19fF
C37284 OR2X1_LOC_589/A OR2X1_LOC_95/Y 0.03fF
C37285 AND2X1_LOC_410/a_36_24# OR2X1_LOC_46/A 0.00fF
C37286 AND2X1_LOC_810/A AND2X1_LOC_319/a_8_24# 0.01fF
C37287 OR2X1_LOC_270/Y OR2X1_LOC_578/a_8_216# 0.01fF
C37288 OR2X1_LOC_427/A OR2X1_LOC_585/A 0.03fF
C37289 OR2X1_LOC_40/Y OR2X1_LOC_504/Y 0.65fF
C37290 OR2X1_LOC_626/a_8_216# AND2X1_LOC_805/Y 0.01fF
C37291 OR2X1_LOC_95/Y OR2X1_LOC_322/Y 0.01fF
C37292 AND2X1_LOC_40/Y OR2X1_LOC_647/A 0.03fF
C37293 OR2X1_LOC_639/B OR2X1_LOC_87/A 0.03fF
C37294 OR2X1_LOC_254/B OR2X1_LOC_483/a_8_216# 0.01fF
C37295 OR2X1_LOC_368/A OR2X1_LOC_322/Y 0.01fF
C37296 AND2X1_LOC_838/Y OR2X1_LOC_6/A 0.02fF
C37297 OR2X1_LOC_51/Y AND2X1_LOC_477/A 0.04fF
C37298 AND2X1_LOC_675/A AND2X1_LOC_778/Y 0.07fF
C37299 OR2X1_LOC_313/Y OR2X1_LOC_418/Y 0.18fF
C37300 OR2X1_LOC_114/Y OR2X1_LOC_510/Y 0.02fF
C37301 OR2X1_LOC_495/a_8_216# OR2X1_LOC_237/Y 0.01fF
C37302 OR2X1_LOC_13/B AND2X1_LOC_247/a_8_24# 0.01fF
C37303 OR2X1_LOC_185/Y AND2X1_LOC_81/B 0.10fF
C37304 OR2X1_LOC_205/a_36_216# OR2X1_LOC_375/A 0.03fF
C37305 AND2X1_LOC_452/Y AND2X1_LOC_454/A 0.01fF
C37306 OR2X1_LOC_240/a_8_216# OR2X1_LOC_240/A 0.18fF
C37307 OR2X1_LOC_400/B OR2X1_LOC_400/A 0.28fF
C37308 AND2X1_LOC_640/Y OR2X1_LOC_48/B 1.23fF
C37309 AND2X1_LOC_573/A AND2X1_LOC_474/Y 0.01fF
C37310 AND2X1_LOC_795/Y AND2X1_LOC_786/Y 0.01fF
C37311 AND2X1_LOC_112/a_8_24# OR2X1_LOC_31/Y 0.01fF
C37312 OR2X1_LOC_223/A OR2X1_LOC_565/A 0.03fF
C37313 AND2X1_LOC_859/Y AND2X1_LOC_286/Y 0.02fF
C37314 OR2X1_LOC_691/Y OR2X1_LOC_801/B 0.01fF
C37315 AND2X1_LOC_316/a_8_24# OR2X1_LOC_206/A 0.01fF
C37316 OR2X1_LOC_319/B OR2X1_LOC_121/B 1.05fF
C37317 OR2X1_LOC_604/A D_INPUT_3 0.04fF
C37318 OR2X1_LOC_18/Y AND2X1_LOC_640/Y 0.02fF
C37319 OR2X1_LOC_485/A AND2X1_LOC_573/A 0.07fF
C37320 OR2X1_LOC_36/Y AND2X1_LOC_806/A 0.03fF
C37321 OR2X1_LOC_91/a_36_216# OR2X1_LOC_44/Y 0.02fF
C37322 OR2X1_LOC_532/B OR2X1_LOC_78/B 0.36fF
C37323 AND2X1_LOC_215/Y AND2X1_LOC_476/A 0.01fF
C37324 OR2X1_LOC_841/a_36_216# OR2X1_LOC_121/B 0.00fF
C37325 AND2X1_LOC_108/a_8_24# OR2X1_LOC_78/A 0.01fF
C37326 OR2X1_LOC_716/a_8_216# OR2X1_LOC_593/B 0.01fF
C37327 OR2X1_LOC_685/B OR2X1_LOC_155/A 0.02fF
C37328 VDD OR2X1_LOC_62/A 1.20fF
C37329 AND2X1_LOC_572/A OR2X1_LOC_89/A 0.01fF
C37330 OR2X1_LOC_502/A OR2X1_LOC_54/Y 0.14fF
C37331 INPUT_5 OR2X1_LOC_22/A 0.05fF
C37332 OR2X1_LOC_114/Y OR2X1_LOC_810/A 0.05fF
C37333 OR2X1_LOC_248/Y OR2X1_LOC_753/A -0.00fF
C37334 AND2X1_LOC_103/a_36_24# OR2X1_LOC_532/B 0.01fF
C37335 OR2X1_LOC_864/A OR2X1_LOC_269/B 0.50fF
C37336 AND2X1_LOC_536/a_8_24# AND2X1_LOC_135/a_8_24# 0.23fF
C37337 AND2X1_LOC_373/a_8_24# OR2X1_LOC_87/A 0.01fF
C37338 OR2X1_LOC_241/B OR2X1_LOC_719/B 0.03fF
C37339 AND2X1_LOC_319/A OR2X1_LOC_418/a_8_216# 0.47fF
C37340 OR2X1_LOC_682/a_8_216# OR2X1_LOC_52/B -0.01fF
C37341 AND2X1_LOC_641/Y OR2X1_LOC_265/Y 0.02fF
C37342 OR2X1_LOC_223/A OR2X1_LOC_190/Y 0.00fF
C37343 OR2X1_LOC_774/Y OR2X1_LOC_269/B 0.01fF
C37344 OR2X1_LOC_40/Y OR2X1_LOC_437/Y 0.17fF
C37345 OR2X1_LOC_224/a_8_216# OR2X1_LOC_59/Y 0.01fF
C37346 OR2X1_LOC_602/a_36_216# AND2X1_LOC_43/B 0.02fF
C37347 OR2X1_LOC_696/a_8_216# OR2X1_LOC_36/Y 0.01fF
C37348 OR2X1_LOC_791/B OR2X1_LOC_285/B 0.01fF
C37349 OR2X1_LOC_92/Y INPUT_1 0.15fF
C37350 OR2X1_LOC_40/Y AND2X1_LOC_641/a_8_24# 0.02fF
C37351 AND2X1_LOC_796/Y AND2X1_LOC_663/A 0.03fF
C37352 OR2X1_LOC_18/Y OR2X1_LOC_416/Y 0.03fF
C37353 OR2X1_LOC_532/B OR2X1_LOC_721/Y 0.19fF
C37354 OR2X1_LOC_185/A OR2X1_LOC_643/Y 1.02fF
C37355 AND2X1_LOC_566/a_8_24# AND2X1_LOC_566/Y 0.00fF
C37356 OR2X1_LOC_3/Y OR2X1_LOC_26/Y 0.29fF
C37357 OR2X1_LOC_121/B OR2X1_LOC_805/A 0.07fF
C37358 OR2X1_LOC_680/A AND2X1_LOC_830/a_36_24# 0.01fF
C37359 OR2X1_LOC_107/Y OR2X1_LOC_47/Y 0.01fF
C37360 OR2X1_LOC_494/a_36_216# AND2X1_LOC_866/A 0.07fF
C37361 OR2X1_LOC_51/B OR2X1_LOC_25/Y 0.03fF
C37362 AND2X1_LOC_866/B OR2X1_LOC_95/Y 0.03fF
C37363 AND2X1_LOC_365/A AND2X1_LOC_727/A 0.03fF
C37364 AND2X1_LOC_654/B OR2X1_LOC_95/Y 0.03fF
C37365 OR2X1_LOC_306/Y OR2X1_LOC_311/Y 0.04fF
C37366 AND2X1_LOC_52/a_8_24# OR2X1_LOC_651/A 0.03fF
C37367 OR2X1_LOC_40/Y OR2X1_LOC_70/A 0.02fF
C37368 OR2X1_LOC_335/A OR2X1_LOC_590/Y 0.01fF
C37369 AND2X1_LOC_7/B AND2X1_LOC_268/a_36_24# 0.02fF
C37370 AND2X1_LOC_281/a_8_24# OR2X1_LOC_269/B 0.14fF
C37371 AND2X1_LOC_370/a_8_24# OR2X1_LOC_437/A 0.05fF
C37372 AND2X1_LOC_64/Y OR2X1_LOC_723/B 0.03fF
C37373 OR2X1_LOC_495/Y OR2X1_LOC_95/Y 0.48fF
C37374 OR2X1_LOC_3/Y AND2X1_LOC_349/B 0.16fF
C37375 AND2X1_LOC_330/a_8_24# OR2X1_LOC_419/Y 0.32fF
C37376 OR2X1_LOC_3/Y OR2X1_LOC_89/A 0.71fF
C37377 OR2X1_LOC_160/A OR2X1_LOC_814/A 0.10fF
C37378 OR2X1_LOC_123/a_8_216# OR2X1_LOC_598/A 0.02fF
C37379 OR2X1_LOC_245/a_8_216# OR2X1_LOC_85/A 0.08fF
C37380 OR2X1_LOC_490/Y AND2X1_LOC_554/B 0.03fF
C37381 AND2X1_LOC_53/a_8_24# OR2X1_LOC_651/A 0.09fF
C37382 AND2X1_LOC_722/A OR2X1_LOC_47/Y 0.05fF
C37383 OR2X1_LOC_790/B AND2X1_LOC_53/Y 0.05fF
C37384 OR2X1_LOC_680/Y OR2X1_LOC_74/A 0.03fF
C37385 OR2X1_LOC_70/Y OR2X1_LOC_7/A 0.15fF
C37386 AND2X1_LOC_661/A AND2X1_LOC_802/a_8_24# 0.01fF
C37387 OR2X1_LOC_71/Y OR2X1_LOC_118/Y 1.95fF
C37388 AND2X1_LOC_53/Y OR2X1_LOC_161/A 0.08fF
C37389 OR2X1_LOC_86/Y OR2X1_LOC_19/B 0.03fF
C37390 OR2X1_LOC_3/Y OR2X1_LOC_820/Y 0.01fF
C37391 AND2X1_LOC_70/Y OR2X1_LOC_358/A 0.03fF
C37392 VDD AND2X1_LOC_257/a_8_24# 0.00fF
C37393 OR2X1_LOC_43/A AND2X1_LOC_727/A 0.14fF
C37394 OR2X1_LOC_743/A OR2X1_LOC_275/A 0.01fF
C37395 OR2X1_LOC_532/B OR2X1_LOC_375/A 2.03fF
C37396 AND2X1_LOC_70/Y OR2X1_LOC_170/Y 0.03fF
C37397 OR2X1_LOC_22/Y AND2X1_LOC_859/Y 0.07fF
C37398 OR2X1_LOC_832/a_36_216# AND2X1_LOC_31/Y 0.02fF
C37399 VDD OR2X1_LOC_88/Y 0.46fF
C37400 OR2X1_LOC_298/Y OR2X1_LOC_31/Y 0.13fF
C37401 OR2X1_LOC_297/Y AND2X1_LOC_663/B 0.01fF
C37402 AND2X1_LOC_303/B D_INPUT_0 0.08fF
C37403 VDD OR2X1_LOC_172/Y 0.35fF
C37404 AND2X1_LOC_12/Y OR2X1_LOC_241/Y 0.07fF
C37405 OR2X1_LOC_151/A OR2X1_LOC_317/B 0.04fF
C37406 AND2X1_LOC_514/Y OR2X1_LOC_7/A 0.07fF
C37407 OR2X1_LOC_237/Y OR2X1_LOC_238/a_8_216# 0.39fF
C37408 OR2X1_LOC_151/A OR2X1_LOC_501/a_8_216# 0.03fF
C37409 OR2X1_LOC_271/Y INPUT_1 0.00fF
C37410 AND2X1_LOC_345/Y AND2X1_LOC_663/B 0.01fF
C37411 OR2X1_LOC_850/B OR2X1_LOC_366/a_8_216# 0.01fF
C37412 OR2X1_LOC_696/A AND2X1_LOC_465/A 0.07fF
C37413 OR2X1_LOC_316/Y AND2X1_LOC_851/B 0.03fF
C37414 AND2X1_LOC_22/Y OR2X1_LOC_301/a_8_216# 0.01fF
C37415 AND2X1_LOC_621/Y OR2X1_LOC_615/Y 0.03fF
C37416 OR2X1_LOC_223/A OR2X1_LOC_161/A 0.68fF
C37417 AND2X1_LOC_831/Y OR2X1_LOC_36/Y 0.08fF
C37418 AND2X1_LOC_89/a_8_24# AND2X1_LOC_47/Y 0.01fF
C37419 OR2X1_LOC_185/A OR2X1_LOC_786/Y 0.14fF
C37420 OR2X1_LOC_335/A AND2X1_LOC_64/Y 0.01fF
C37421 AND2X1_LOC_514/Y OR2X1_LOC_320/Y 0.07fF
C37422 OR2X1_LOC_262/Y OR2X1_LOC_71/Y 0.03fF
C37423 AND2X1_LOC_36/Y OR2X1_LOC_548/a_8_216# 0.01fF
C37424 OR2X1_LOC_118/Y D_INPUT_1 0.02fF
C37425 OR2X1_LOC_325/B OR2X1_LOC_303/B 0.03fF
C37426 OR2X1_LOC_43/A OR2X1_LOC_95/Y 0.15fF
C37427 OR2X1_LOC_275/A OR2X1_LOC_246/A 0.01fF
C37428 OR2X1_LOC_624/B OR2X1_LOC_814/A 0.03fF
C37429 AND2X1_LOC_300/a_8_24# OR2X1_LOC_593/B 0.01fF
C37430 AND2X1_LOC_110/Y OR2X1_LOC_788/B 0.01fF
C37431 OR2X1_LOC_619/Y AND2X1_LOC_204/Y 0.08fF
C37432 AND2X1_LOC_572/a_8_24# OR2X1_LOC_106/Y 0.01fF
C37433 OR2X1_LOC_364/A OR2X1_LOC_112/B 0.01fF
C37434 OR2X1_LOC_791/B OR2X1_LOC_792/A 0.44fF
C37435 OR2X1_LOC_185/Y OR2X1_LOC_112/B 0.03fF
C37436 AND2X1_LOC_347/B AND2X1_LOC_789/Y 0.02fF
C37437 OR2X1_LOC_599/A OR2X1_LOC_47/Y 0.83fF
C37438 AND2X1_LOC_27/a_8_24# OR2X1_LOC_34/B 0.01fF
C37439 AND2X1_LOC_817/B OR2X1_LOC_771/a_8_216# 0.01fF
C37440 OR2X1_LOC_625/Y OR2X1_LOC_753/Y 0.05fF
C37441 OR2X1_LOC_10/a_36_216# OR2X1_LOC_753/A 0.17fF
C37442 AND2X1_LOC_22/Y OR2X1_LOC_828/Y 0.03fF
C37443 OR2X1_LOC_316/Y OR2X1_LOC_595/Y 0.02fF
C37444 AND2X1_LOC_56/B OR2X1_LOC_214/B 0.03fF
C37445 OR2X1_LOC_139/A OR2X1_LOC_267/Y 0.03fF
C37446 AND2X1_LOC_392/A OR2X1_LOC_268/Y 0.03fF
C37447 AND2X1_LOC_53/Y AND2X1_LOC_51/Y 0.04fF
C37448 AND2X1_LOC_56/B OR2X1_LOC_241/B 0.38fF
C37449 OR2X1_LOC_477/a_8_216# AND2X1_LOC_51/Y 0.01fF
C37450 OR2X1_LOC_185/Y OR2X1_LOC_66/Y 0.03fF
C37451 AND2X1_LOC_91/B OR2X1_LOC_673/B 0.00fF
C37452 AND2X1_LOC_360/a_8_24# OR2X1_LOC_384/Y 0.24fF
C37453 AND2X1_LOC_584/a_8_24# OR2X1_LOC_451/B 0.20fF
C37454 OR2X1_LOC_184/Y OR2X1_LOC_7/A 0.00fF
C37455 AND2X1_LOC_338/Y AND2X1_LOC_350/B 0.00fF
C37456 OR2X1_LOC_87/A OR2X1_LOC_590/a_8_216# 0.01fF
C37457 AND2X1_LOC_22/Y AND2X1_LOC_522/a_36_24# 0.01fF
C37458 AND2X1_LOC_423/a_8_24# OR2X1_LOC_446/B 0.01fF
C37459 OR2X1_LOC_56/A OR2X1_LOC_183/a_8_216# 0.03fF
C37460 AND2X1_LOC_445/a_8_24# OR2X1_LOC_428/A 0.01fF
C37461 AND2X1_LOC_31/Y OR2X1_LOC_539/Y 0.07fF
C37462 AND2X1_LOC_578/A AND2X1_LOC_675/a_8_24# 0.04fF
C37463 OR2X1_LOC_392/B OR2X1_LOC_549/A 0.10fF
C37464 OR2X1_LOC_545/B OR2X1_LOC_471/Y 0.16fF
C37465 OR2X1_LOC_604/A AND2X1_LOC_780/a_8_24# 0.01fF
C37466 VDD OR2X1_LOC_170/a_8_216# 0.00fF
C37467 OR2X1_LOC_188/Y OR2X1_LOC_719/B 0.00fF
C37468 OR2X1_LOC_6/B OR2X1_LOC_748/Y 0.02fF
C37469 OR2X1_LOC_223/A AND2X1_LOC_51/Y 0.03fF
C37470 OR2X1_LOC_87/A OR2X1_LOC_160/a_8_216# 0.05fF
C37471 OR2X1_LOC_468/Y OR2X1_LOC_854/A 0.02fF
C37472 AND2X1_LOC_31/Y OR2X1_LOC_779/a_8_216# 0.01fF
C37473 OR2X1_LOC_48/B AND2X1_LOC_592/a_8_24# 0.04fF
C37474 AND2X1_LOC_91/B OR2X1_LOC_356/a_8_216# 0.01fF
C37475 OR2X1_LOC_151/A AND2X1_LOC_44/Y 0.14fF
C37476 VDD OR2X1_LOC_397/Y 0.12fF
C37477 AND2X1_LOC_525/a_8_24# OR2X1_LOC_705/B 0.10fF
C37478 OR2X1_LOC_256/a_36_216# OR2X1_LOC_437/A 0.00fF
C37479 AND2X1_LOC_95/Y OR2X1_LOC_342/a_8_216# 0.01fF
C37480 OR2X1_LOC_131/Y AND2X1_LOC_216/A 0.10fF
C37481 OR2X1_LOC_53/Y OR2X1_LOC_600/A 0.03fF
C37482 AND2X1_LOC_599/a_36_24# OR2X1_LOC_598/Y 0.01fF
C37483 OR2X1_LOC_188/Y OR2X1_LOC_542/B 0.03fF
C37484 OR2X1_LOC_805/A AND2X1_LOC_268/a_36_24# 0.01fF
C37485 VDD AND2X1_LOC_206/a_8_24# -0.00fF
C37486 OR2X1_LOC_203/Y AND2X1_LOC_268/a_8_24# 0.04fF
C37487 OR2X1_LOC_705/B AND2X1_LOC_51/Y 0.26fF
C37488 AND2X1_LOC_387/B OR2X1_LOC_750/Y 0.10fF
C37489 OR2X1_LOC_304/a_8_216# OR2X1_LOC_56/A 0.03fF
C37490 OR2X1_LOC_89/A AND2X1_LOC_772/a_8_24# 0.01fF
C37491 AND2X1_LOC_851/a_36_24# AND2X1_LOC_465/A 0.00fF
C37492 AND2X1_LOC_489/Y AND2X1_LOC_657/A 0.13fF
C37493 OR2X1_LOC_840/A OR2X1_LOC_356/B 0.10fF
C37494 AND2X1_LOC_116/Y AND2X1_LOC_216/a_8_24# 0.02fF
C37495 AND2X1_LOC_447/Y OR2X1_LOC_16/A 0.02fF
C37496 OR2X1_LOC_583/a_8_216# OR2X1_LOC_584/Y 0.39fF
C37497 AND2X1_LOC_219/a_8_24# OR2X1_LOC_16/A 0.01fF
C37498 AND2X1_LOC_334/Y OR2X1_LOC_16/A 0.01fF
C37499 OR2X1_LOC_634/A AND2X1_LOC_416/a_36_24# 0.00fF
C37500 OR2X1_LOC_862/a_8_216# OR2X1_LOC_391/A 0.03fF
C37501 OR2X1_LOC_648/A OR2X1_LOC_161/B 0.08fF
C37502 AND2X1_LOC_509/Y OR2X1_LOC_816/A 0.03fF
C37503 AND2X1_LOC_866/A OR2X1_LOC_47/Y 0.06fF
C37504 INPUT_0 OR2X1_LOC_428/A 0.10fF
C37505 OR2X1_LOC_40/Y AND2X1_LOC_499/a_8_24# 0.02fF
C37506 AND2X1_LOC_347/Y OR2X1_LOC_494/A 0.00fF
C37507 AND2X1_LOC_101/B OR2X1_LOC_13/B 0.10fF
C37508 OR2X1_LOC_621/B OR2X1_LOC_621/a_8_216# 0.01fF
C37509 OR2X1_LOC_155/a_8_216# OR2X1_LOC_160/B 0.01fF
C37510 AND2X1_LOC_91/B AND2X1_LOC_40/Y 5.95fF
C37511 OR2X1_LOC_244/a_8_216# OR2X1_LOC_267/Y 0.01fF
C37512 OR2X1_LOC_696/A OR2X1_LOC_376/A 0.20fF
C37513 AND2X1_LOC_3/Y OR2X1_LOC_366/Y 0.11fF
C37514 AND2X1_LOC_148/a_8_24# AND2X1_LOC_213/B 0.01fF
C37515 OR2X1_LOC_866/B OR2X1_LOC_392/A 0.01fF
C37516 OR2X1_LOC_482/a_36_216# OR2X1_LOC_51/Y 0.00fF
C37517 OR2X1_LOC_6/B OR2X1_LOC_14/a_36_216# 0.02fF
C37518 VDD OR2X1_LOC_629/B 0.00fF
C37519 OR2X1_LOC_604/A AND2X1_LOC_254/a_36_24# 0.00fF
C37520 OR2X1_LOC_487/Y OR2X1_LOC_437/A 0.01fF
C37521 AND2X1_LOC_658/B OR2X1_LOC_40/Y 16.02fF
C37522 OR2X1_LOC_160/B AND2X1_LOC_18/Y 5.33fF
C37523 OR2X1_LOC_6/B AND2X1_LOC_404/B 0.21fF
C37524 AND2X1_LOC_48/A OR2X1_LOC_513/a_8_216# 0.12fF
C37525 AND2X1_LOC_47/Y AND2X1_LOC_280/a_8_24# 0.10fF
C37526 AND2X1_LOC_539/Y AND2X1_LOC_809/A 0.01fF
C37527 OR2X1_LOC_450/Y OR2X1_LOC_467/A 0.73fF
C37528 AND2X1_LOC_564/B OR2X1_LOC_427/A 0.10fF
C37529 OR2X1_LOC_856/B AND2X1_LOC_7/B 0.07fF
C37530 AND2X1_LOC_253/a_8_24# OR2X1_LOC_161/B 0.06fF
C37531 AND2X1_LOC_784/Y OR2X1_LOC_744/A 0.03fF
C37532 OR2X1_LOC_8/Y VDD 0.52fF
C37533 OR2X1_LOC_427/A OR2X1_LOC_368/Y 0.00fF
C37534 OR2X1_LOC_186/Y OR2X1_LOC_798/Y 0.01fF
C37535 AND2X1_LOC_81/B OR2X1_LOC_510/a_36_216# 0.00fF
C37536 OR2X1_LOC_121/Y OR2X1_LOC_216/A 0.01fF
C37537 AND2X1_LOC_367/A AND2X1_LOC_476/Y 0.09fF
C37538 AND2X1_LOC_362/B AND2X1_LOC_367/A 0.10fF
C37539 OR2X1_LOC_326/a_8_216# AND2X1_LOC_110/Y 0.01fF
C37540 OR2X1_LOC_97/A AND2X1_LOC_290/a_8_24# 0.01fF
C37541 OR2X1_LOC_269/B OR2X1_LOC_714/a_36_216# 0.03fF
C37542 OR2X1_LOC_440/a_8_216# OR2X1_LOC_78/A 0.01fF
C37543 AND2X1_LOC_207/a_8_24# AND2X1_LOC_207/A 0.19fF
C37544 AND2X1_LOC_47/Y OR2X1_LOC_742/B 0.03fF
C37545 OR2X1_LOC_623/B OR2X1_LOC_185/a_36_216# 0.15fF
C37546 OR2X1_LOC_763/Y OR2X1_LOC_387/A 0.18fF
C37547 AND2X1_LOC_721/Y AND2X1_LOC_848/Y 0.03fF
C37548 AND2X1_LOC_564/B AND2X1_LOC_464/a_8_24# -0.00fF
C37549 D_INPUT_0 OR2X1_LOC_446/B 0.05fF
C37550 OR2X1_LOC_188/Y AND2X1_LOC_56/B 0.06fF
C37551 OR2X1_LOC_744/A AND2X1_LOC_434/Y 0.07fF
C37552 OR2X1_LOC_11/Y OR2X1_LOC_428/A 0.00fF
C37553 OR2X1_LOC_176/Y OR2X1_LOC_91/Y 0.01fF
C37554 AND2X1_LOC_702/Y OR2X1_LOC_321/a_8_216# 0.01fF
C37555 OR2X1_LOC_631/B OR2X1_LOC_554/a_36_216# 0.00fF
C37556 OR2X1_LOC_561/Y OR2X1_LOC_78/A 0.00fF
C37557 INPUT_4 INPUT_7 0.06fF
C37558 OR2X1_LOC_40/Y AND2X1_LOC_357/a_8_24# 0.09fF
C37559 OR2X1_LOC_653/Y OR2X1_LOC_661/A 0.04fF
C37560 OR2X1_LOC_479/Y OR2X1_LOC_605/Y 0.12fF
C37561 AND2X1_LOC_456/Y OR2X1_LOC_503/a_8_216# 0.47fF
C37562 OR2X1_LOC_269/B OR2X1_LOC_121/A 0.03fF
C37563 OR2X1_LOC_648/A OR2X1_LOC_435/B 0.03fF
C37564 OR2X1_LOC_419/Y AND2X1_LOC_486/a_8_24# 0.26fF
C37565 OR2X1_LOC_78/B OR2X1_LOC_78/a_36_216# 0.01fF
C37566 OR2X1_LOC_854/a_36_216# AND2X1_LOC_110/Y 0.00fF
C37567 OR2X1_LOC_164/Y OR2X1_LOC_56/A 0.02fF
C37568 OR2X1_LOC_709/a_8_216# OR2X1_LOC_738/A 0.41fF
C37569 AND2X1_LOC_754/a_8_24# AND2X1_LOC_12/Y 0.02fF
C37570 AND2X1_LOC_540/a_8_24# OR2X1_LOC_56/A 0.01fF
C37571 OR2X1_LOC_654/A OR2X1_LOC_338/A 0.07fF
C37572 AND2X1_LOC_352/B OR2X1_LOC_92/Y 0.05fF
C37573 OR2X1_LOC_136/a_8_216# OR2X1_LOC_743/A 0.04fF
C37574 VDD OR2X1_LOC_837/a_8_216# 0.21fF
C37575 OR2X1_LOC_804/A OR2X1_LOC_228/Y 1.17fF
C37576 OR2X1_LOC_88/Y OR2X1_LOC_67/Y 0.03fF
C37577 VDD AND2X1_LOC_76/Y 0.26fF
C37578 AND2X1_LOC_140/a_8_24# AND2X1_LOC_772/Y -0.00fF
C37579 OR2X1_LOC_78/A AND2X1_LOC_424/a_8_24# 0.03fF
C37580 OR2X1_LOC_840/A OR2X1_LOC_168/B 0.03fF
C37581 OR2X1_LOC_161/A OR2X1_LOC_777/a_8_216# 0.03fF
C37582 AND2X1_LOC_372/a_36_24# OR2X1_LOC_541/A 0.00fF
C37583 AND2X1_LOC_360/a_8_24# OR2X1_LOC_91/A 0.05fF
C37584 OR2X1_LOC_648/A OR2X1_LOC_61/Y 0.05fF
C37585 AND2X1_LOC_553/a_8_24# AND2X1_LOC_113/Y 0.19fF
C37586 OR2X1_LOC_829/A OR2X1_LOC_44/Y 0.15fF
C37587 AND2X1_LOC_251/a_8_24# OR2X1_LOC_362/A 0.01fF
C37588 OR2X1_LOC_315/a_36_216# OR2X1_LOC_44/Y 0.01fF
C37589 OR2X1_LOC_58/Y OR2X1_LOC_32/B 0.00fF
C37590 VDD OR2X1_LOC_803/B 0.05fF
C37591 OR2X1_LOC_205/a_36_216# OR2X1_LOC_549/A 0.01fF
C37592 OR2X1_LOC_12/Y AND2X1_LOC_638/a_8_24# 0.00fF
C37593 OR2X1_LOC_326/B OR2X1_LOC_324/B 0.79fF
C37594 OR2X1_LOC_270/Y OR2X1_LOC_366/Y 0.00fF
C37595 OR2X1_LOC_528/Y AND2X1_LOC_580/A 0.06fF
C37596 OR2X1_LOC_252/Y OR2X1_LOC_627/Y 0.71fF
C37597 VDD OR2X1_LOC_67/A 0.21fF
C37598 OR2X1_LOC_426/B OR2X1_LOC_118/Y 0.09fF
C37599 OR2X1_LOC_778/Y OR2X1_LOC_356/A 0.10fF
C37600 AND2X1_LOC_18/Y OR2X1_LOC_553/A 0.24fF
C37601 AND2X1_LOC_794/B OR2X1_LOC_52/B 0.46fF
C37602 AND2X1_LOC_357/A OR2X1_LOC_6/A 0.00fF
C37603 OR2X1_LOC_6/B OR2X1_LOC_36/Y 0.04fF
C37604 OR2X1_LOC_517/A OR2X1_LOC_92/Y 0.10fF
C37605 AND2X1_LOC_713/Y OR2X1_LOC_36/Y 0.01fF
C37606 AND2X1_LOC_148/Y AND2X1_LOC_213/B 0.26fF
C37607 AND2X1_LOC_95/Y AND2X1_LOC_24/a_8_24# 0.01fF
C37608 OR2X1_LOC_26/Y AND2X1_LOC_477/Y 0.07fF
C37609 AND2X1_LOC_784/A OR2X1_LOC_309/a_36_216# 0.01fF
C37610 AND2X1_LOC_19/Y OR2X1_LOC_660/B 0.02fF
C37611 OR2X1_LOC_599/A AND2X1_LOC_732/B 0.00fF
C37612 OR2X1_LOC_11/Y OR2X1_LOC_380/a_36_216# 0.00fF
C37613 OR2X1_LOC_604/A AND2X1_LOC_806/A 0.03fF
C37614 OR2X1_LOC_721/Y OR2X1_LOC_734/a_8_216# 0.02fF
C37615 OR2X1_LOC_759/A OR2X1_LOC_44/Y 0.00fF
C37616 AND2X1_LOC_347/Y OR2X1_LOC_427/A 0.07fF
C37617 OR2X1_LOC_136/a_8_216# OR2X1_LOC_246/A 0.12fF
C37618 OR2X1_LOC_319/B OR2X1_LOC_856/B 0.17fF
C37619 OR2X1_LOC_160/A OR2X1_LOC_501/B 0.09fF
C37620 AND2X1_LOC_721/Y AND2X1_LOC_464/Y 0.01fF
C37621 OR2X1_LOC_176/Y OR2X1_LOC_417/Y 0.30fF
C37622 OR2X1_LOC_176/a_8_216# AND2X1_LOC_514/Y 0.03fF
C37623 OR2X1_LOC_64/Y OR2X1_LOC_428/A 0.67fF
C37624 OR2X1_LOC_89/A AND2X1_LOC_477/Y 0.07fF
C37625 VDD AND2X1_LOC_374/Y 0.06fF
C37626 OR2X1_LOC_135/Y OR2X1_LOC_304/Y 0.23fF
C37627 AND2X1_LOC_307/a_36_24# OR2X1_LOC_428/A 0.01fF
C37628 AND2X1_LOC_729/B OR2X1_LOC_16/A 0.09fF
C37629 OR2X1_LOC_254/a_36_216# OR2X1_LOC_161/B 0.00fF
C37630 AND2X1_LOC_362/B OR2X1_LOC_490/Y 0.68fF
C37631 OR2X1_LOC_74/A AND2X1_LOC_476/Y 0.21fF
C37632 OR2X1_LOC_219/B AND2X1_LOC_18/Y 0.03fF
C37633 AND2X1_LOC_661/A AND2X1_LOC_436/Y 1.09fF
C37634 OR2X1_LOC_83/A OR2X1_LOC_66/A 0.03fF
C37635 VDD OR2X1_LOC_52/B 0.92fF
C37636 OR2X1_LOC_389/B OR2X1_LOC_66/A 0.41fF
C37637 VDD OR2X1_LOC_672/Y 0.19fF
C37638 OR2X1_LOC_318/Y OR2X1_LOC_856/B 0.13fF
C37639 OR2X1_LOC_3/Y AND2X1_LOC_194/Y 0.01fF
C37640 OR2X1_LOC_64/Y OR2X1_LOC_595/A 0.51fF
C37641 OR2X1_LOC_517/A OR2X1_LOC_65/B 0.19fF
C37642 AND2X1_LOC_340/Y OR2X1_LOC_416/Y 0.03fF
C37643 OR2X1_LOC_429/Y OR2X1_LOC_581/Y 0.05fF
C37644 OR2X1_LOC_417/Y AND2X1_LOC_212/Y 0.05fF
C37645 AND2X1_LOC_40/Y OR2X1_LOC_799/A 0.08fF
C37646 VDD OR2X1_LOC_141/B 0.10fF
C37647 AND2X1_LOC_12/Y OR2X1_LOC_216/A 0.07fF
C37648 OR2X1_LOC_715/B OR2X1_LOC_201/Y 0.07fF
C37649 OR2X1_LOC_502/A OR2X1_LOC_161/A 0.18fF
C37650 AND2X1_LOC_364/Y AND2X1_LOC_354/B 0.03fF
C37651 AND2X1_LOC_59/Y OR2X1_LOC_840/A 0.01fF
C37652 OR2X1_LOC_61/Y OR2X1_LOC_405/a_8_216# 0.01fF
C37653 VDD AND2X1_LOC_489/Y 0.21fF
C37654 OR2X1_LOC_632/A OR2X1_LOC_575/A 0.01fF
C37655 OR2X1_LOC_538/A OR2X1_LOC_468/Y 0.00fF
C37656 AND2X1_LOC_724/Y OR2X1_LOC_485/A 0.01fF
C37657 OR2X1_LOC_756/B OR2X1_LOC_653/A 0.01fF
C37658 OR2X1_LOC_851/A OR2X1_LOC_185/A 0.12fF
C37659 OR2X1_LOC_329/B OR2X1_LOC_26/Y 0.11fF
C37660 AND2X1_LOC_56/B AND2X1_LOC_189/a_8_24# 0.01fF
C37661 OR2X1_LOC_57/Y OR2X1_LOC_6/A 0.01fF
C37662 OR2X1_LOC_631/B OR2X1_LOC_630/B 0.00fF
C37663 INPUT_1 AND2X1_LOC_44/Y 0.03fF
C37664 AND2X1_LOC_530/a_8_24# OR2X1_LOC_54/Y 0.04fF
C37665 OR2X1_LOC_756/B OR2X1_LOC_673/Y 0.01fF
C37666 AND2X1_LOC_76/Y AND2X1_LOC_274/a_8_24# 0.01fF
C37667 AND2X1_LOC_535/Y AND2X1_LOC_798/Y 0.16fF
C37668 INPUT_4 OR2X1_LOC_426/A 0.00fF
C37669 OR2X1_LOC_643/a_36_216# AND2X1_LOC_92/Y 0.01fF
C37670 AND2X1_LOC_183/a_8_24# OR2X1_LOC_190/A 0.04fF
C37671 OR2X1_LOC_185/A OR2X1_LOC_220/B 0.03fF
C37672 OR2X1_LOC_764/Y OR2X1_LOC_744/A 0.01fF
C37673 OR2X1_LOC_856/B OR2X1_LOC_805/A 0.07fF
C37674 OR2X1_LOC_417/A OR2X1_LOC_428/A 1.09fF
C37675 OR2X1_LOC_147/A OR2X1_LOC_711/A 0.01fF
C37676 OR2X1_LOC_502/A AND2X1_LOC_25/Y 0.02fF
C37677 OR2X1_LOC_329/B OR2X1_LOC_89/A 0.74fF
C37678 OR2X1_LOC_160/A OR2X1_LOC_317/A 0.02fF
C37679 AND2X1_LOC_810/A OR2X1_LOC_167/Y 0.16fF
C37680 AND2X1_LOC_353/a_8_24# AND2X1_LOC_514/Y 0.01fF
C37681 OR2X1_LOC_703/B OR2X1_LOC_620/Y 0.01fF
C37682 AND2X1_LOC_12/Y OR2X1_LOC_362/B 0.00fF
C37683 OR2X1_LOC_8/Y OR2X1_LOC_826/a_8_216# 0.02fF
C37684 OR2X1_LOC_814/A OR2X1_LOC_768/a_8_216# 0.05fF
C37685 AND2X1_LOC_486/Y AND2X1_LOC_784/A 0.08fF
C37686 OR2X1_LOC_45/B AND2X1_LOC_318/Y 0.01fF
C37687 OR2X1_LOC_620/Y OR2X1_LOC_87/A 0.03fF
C37688 OR2X1_LOC_532/B OR2X1_LOC_549/A 0.20fF
C37689 OR2X1_LOC_185/Y OR2X1_LOC_861/a_36_216# 0.00fF
C37690 OR2X1_LOC_521/Y OR2X1_LOC_271/Y 0.01fF
C37691 OR2X1_LOC_155/A AND2X1_LOC_424/a_8_24# 0.03fF
C37692 OR2X1_LOC_6/A OR2X1_LOC_48/B 0.01fF
C37693 OR2X1_LOC_664/a_8_216# OR2X1_LOC_664/Y 0.05fF
C37694 OR2X1_LOC_305/a_36_216# OR2X1_LOC_48/B 0.00fF
C37695 OR2X1_LOC_656/B OR2X1_LOC_264/a_8_216# 0.02fF
C37696 OR2X1_LOC_473/Y AND2X1_LOC_92/Y 0.02fF
C37697 OR2X1_LOC_677/a_36_216# OR2X1_LOC_74/A 0.02fF
C37698 OR2X1_LOC_213/A OR2X1_LOC_161/A 0.02fF
C37699 AND2X1_LOC_160/Y AND2X1_LOC_708/a_8_24# 0.21fF
C37700 OR2X1_LOC_185/A OR2X1_LOC_204/Y 0.01fF
C37701 OR2X1_LOC_18/Y OR2X1_LOC_6/A 1.02fF
C37702 OR2X1_LOC_119/a_8_216# OR2X1_LOC_744/A 0.01fF
C37703 OR2X1_LOC_317/B OR2X1_LOC_714/A 0.03fF
C37704 OR2X1_LOC_112/a_8_216# OR2X1_LOC_436/Y 0.01fF
C37705 OR2X1_LOC_471/Y OR2X1_LOC_190/a_8_216# 0.40fF
C37706 OR2X1_LOC_218/Y AND2X1_LOC_65/A 0.03fF
C37707 AND2X1_LOC_305/a_8_24# OR2X1_LOC_269/B 0.00fF
C37708 AND2X1_LOC_736/Y OR2X1_LOC_438/a_8_216# 0.06fF
C37709 AND2X1_LOC_850/a_8_24# AND2X1_LOC_806/A 0.01fF
C37710 AND2X1_LOC_59/Y OR2X1_LOC_222/A 0.73fF
C37711 AND2X1_LOC_41/A AND2X1_LOC_67/Y 0.45fF
C37712 OR2X1_LOC_64/Y AND2X1_LOC_468/a_36_24# 0.01fF
C37713 OR2X1_LOC_51/Y AND2X1_LOC_465/Y 0.02fF
C37714 OR2X1_LOC_600/A INPUT_1 0.73fF
C37715 OR2X1_LOC_343/B OR2X1_LOC_843/B 0.30fF
C37716 OR2X1_LOC_187/a_8_216# AND2X1_LOC_711/Y 0.01fF
C37717 AND2X1_LOC_12/Y OR2X1_LOC_468/Y 0.03fF
C37718 VDD OR2X1_LOC_520/A -0.00fF
C37719 OR2X1_LOC_256/a_36_216# OR2X1_LOC_753/A 0.00fF
C37720 OR2X1_LOC_36/Y AND2X1_LOC_436/B 0.01fF
C37721 OR2X1_LOC_653/a_36_216# OR2X1_LOC_502/A 0.01fF
C37722 AND2X1_LOC_648/a_8_24# OR2X1_LOC_44/Y 0.00fF
C37723 OR2X1_LOC_244/A AND2X1_LOC_18/Y 0.07fF
C37724 OR2X1_LOC_177/a_8_216# OR2X1_LOC_47/Y 0.01fF
C37725 AND2X1_LOC_274/a_8_24# OR2X1_LOC_52/B 0.03fF
C37726 OR2X1_LOC_36/Y AND2X1_LOC_139/B 0.03fF
C37727 AND2X1_LOC_12/Y AND2X1_LOC_385/a_8_24# 0.02fF
C37728 OR2X1_LOC_809/a_8_216# OR2X1_LOC_539/Y 0.04fF
C37729 OR2X1_LOC_715/B OR2X1_LOC_201/a_8_216# 0.24fF
C37730 AND2X1_LOC_113/Y OR2X1_LOC_26/Y 0.01fF
C37731 OR2X1_LOC_748/A AND2X1_LOC_848/Y 0.04fF
C37732 OR2X1_LOC_154/A OR2X1_LOC_87/A 1.47fF
C37733 OR2X1_LOC_778/Y AND2X1_LOC_43/B 0.09fF
C37734 AND2X1_LOC_535/Y AND2X1_LOC_169/a_36_24# 0.00fF
C37735 D_INPUT_5 AND2X1_LOC_1/Y 0.01fF
C37736 D_INPUT_0 OR2X1_LOC_56/A 0.03fF
C37737 OR2X1_LOC_472/A AND2X1_LOC_43/B 1.84fF
C37738 OR2X1_LOC_502/A AND2X1_LOC_51/Y 1.81fF
C37739 OR2X1_LOC_743/A AND2X1_LOC_643/a_36_24# 0.01fF
C37740 OR2X1_LOC_624/A AND2X1_LOC_3/Y 0.05fF
C37741 OR2X1_LOC_121/Y OR2X1_LOC_205/Y 0.35fF
C37742 AND2X1_LOC_154/Y OR2X1_LOC_619/Y 0.03fF
C37743 OR2X1_LOC_487/a_36_216# AND2X1_LOC_573/A 0.01fF
C37744 VDD OR2X1_LOC_651/A 0.14fF
C37745 OR2X1_LOC_600/A OR2X1_LOC_751/a_8_216# 0.01fF
C37746 AND2X1_LOC_70/Y OR2X1_LOC_639/a_8_216# 0.01fF
C37747 OR2X1_LOC_74/A OR2X1_LOC_595/a_8_216# 0.05fF
C37748 OR2X1_LOC_696/A OR2X1_LOC_384/Y 0.10fF
C37749 AND2X1_LOC_810/Y AND2X1_LOC_436/Y 0.02fF
C37750 OR2X1_LOC_40/Y OR2X1_LOC_47/Y 7.47fF
C37751 OR2X1_LOC_377/A AND2X1_LOC_42/B 5.91fF
C37752 AND2X1_LOC_217/a_8_24# AND2X1_LOC_772/Y 0.01fF
C37753 AND2X1_LOC_1/Y AND2X1_LOC_22/a_8_24# 0.10fF
C37754 OR2X1_LOC_31/Y AND2X1_LOC_219/Y 0.14fF
C37755 OR2X1_LOC_364/A OR2X1_LOC_574/A 0.10fF
C37756 OR2X1_LOC_177/Y AND2X1_LOC_405/a_8_24# 0.01fF
C37757 AND2X1_LOC_364/Y AND2X1_LOC_863/Y 0.38fF
C37758 OR2X1_LOC_185/Y OR2X1_LOC_574/A 0.10fF
C37759 OR2X1_LOC_709/A AND2X1_LOC_679/a_8_24# 0.01fF
C37760 AND2X1_LOC_51/Y OR2X1_LOC_571/B 0.04fF
C37761 AND2X1_LOC_12/Y OR2X1_LOC_846/B 0.04fF
C37762 OR2X1_LOC_141/B OR2X1_LOC_267/a_36_216# 0.00fF
C37763 OR2X1_LOC_529/Y OR2X1_LOC_36/Y 0.04fF
C37764 OR2X1_LOC_144/Y AND2X1_LOC_678/a_8_24# 0.24fF
C37765 AND2X1_LOC_12/Y AND2X1_LOC_1/Y 0.00fF
C37766 OR2X1_LOC_675/a_36_216# OR2X1_LOC_553/A 0.00fF
C37767 OR2X1_LOC_744/A AND2X1_LOC_851/B 3.57fF
C37768 OR2X1_LOC_354/A OR2X1_LOC_532/B 0.00fF
C37769 AND2X1_LOC_42/B OR2X1_LOC_203/Y 0.07fF
C37770 OR2X1_LOC_691/A AND2X1_LOC_31/Y 0.03fF
C37771 AND2X1_LOC_40/Y AND2X1_LOC_600/a_36_24# 0.01fF
C37772 OR2X1_LOC_639/B OR2X1_LOC_639/A 0.09fF
C37773 OR2X1_LOC_615/Y OR2X1_LOC_59/Y 0.03fF
C37774 OR2X1_LOC_246/A AND2X1_LOC_643/a_36_24# 0.06fF
C37775 OR2X1_LOC_400/A AND2X1_LOC_51/Y 0.00fF
C37776 VDD OR2X1_LOC_771/a_8_216# 0.00fF
C37777 OR2X1_LOC_790/B AND2X1_LOC_48/A 0.01fF
C37778 OR2X1_LOC_8/Y OR2X1_LOC_67/Y 0.04fF
C37779 OR2X1_LOC_246/A OR2X1_LOC_118/Y 0.02fF
C37780 AND2X1_LOC_56/B OR2X1_LOC_193/A 0.03fF
C37781 AND2X1_LOC_48/A OR2X1_LOC_161/A 0.13fF
C37782 AND2X1_LOC_182/a_8_24# AND2X1_LOC_222/Y 0.01fF
C37783 AND2X1_LOC_56/B AND2X1_LOC_136/a_36_24# 0.00fF
C37784 OR2X1_LOC_472/B OR2X1_LOC_39/A 0.15fF
C37785 OR2X1_LOC_494/A OR2X1_LOC_437/A 0.14fF
C37786 OR2X1_LOC_70/Y OR2X1_LOC_86/a_8_216# 0.15fF
C37787 VDD AND2X1_LOC_216/A 0.54fF
C37788 INPUT_1 OR2X1_LOC_619/Y 0.03fF
C37789 AND2X1_LOC_719/Y AND2X1_LOC_563/Y 0.03fF
C37790 AND2X1_LOC_92/Y OR2X1_LOC_241/B 0.04fF
C37791 OR2X1_LOC_312/Y AND2X1_LOC_212/B 0.03fF
C37792 OR2X1_LOC_485/A OR2X1_LOC_371/Y 0.07fF
C37793 AND2X1_LOC_2/Y OR2X1_LOC_451/B 0.01fF
C37794 OR2X1_LOC_59/Y AND2X1_LOC_203/Y 0.01fF
C37795 AND2X1_LOC_404/B OR2X1_LOC_598/A 0.06fF
C37796 D_INPUT_0 AND2X1_LOC_9/a_8_24# 0.10fF
C37797 OR2X1_LOC_778/B OR2X1_LOC_493/Y 0.04fF
C37798 OR2X1_LOC_3/Y OR2X1_LOC_17/Y 0.03fF
C37799 AND2X1_LOC_706/Y OR2X1_LOC_423/Y 0.03fF
C37800 AND2X1_LOC_57/Y OR2X1_LOC_198/a_8_216# 0.05fF
C37801 OR2X1_LOC_3/Y OR2X1_LOC_282/Y 0.21fF
C37802 OR2X1_LOC_625/Y AND2X1_LOC_866/A 0.09fF
C37803 OR2X1_LOC_446/Y OR2X1_LOC_707/A 0.01fF
C37804 OR2X1_LOC_416/Y OR2X1_LOC_585/A 0.03fF
C37805 OR2X1_LOC_161/B OR2X1_LOC_112/A 0.00fF
C37806 OR2X1_LOC_18/Y AND2X1_LOC_139/A 0.03fF
C37807 AND2X1_LOC_56/B D_INPUT_0 0.03fF
C37808 OR2X1_LOC_743/A AND2X1_LOC_855/a_8_24# 0.01fF
C37809 OR2X1_LOC_154/A AND2X1_LOC_15/a_36_24# 0.00fF
C37810 OR2X1_LOC_446/B OR2X1_LOC_515/A 0.06fF
C37811 OR2X1_LOC_461/a_8_216# OR2X1_LOC_68/B 0.01fF
C37812 OR2X1_LOC_831/A OR2X1_LOC_303/B 0.61fF
C37813 AND2X1_LOC_59/Y OR2X1_LOC_241/Y 0.24fF
C37814 OR2X1_LOC_744/A OR2X1_LOC_88/a_36_216# 0.00fF
C37815 OR2X1_LOC_813/a_8_216# OR2X1_LOC_71/A 0.01fF
C37816 AND2X1_LOC_8/Y D_INPUT_0 1.53fF
C37817 AND2X1_LOC_839/A OR2X1_LOC_753/A 0.01fF
C37818 AND2X1_LOC_576/Y AND2X1_LOC_227/Y 0.02fF
C37819 OR2X1_LOC_288/A OR2X1_LOC_269/B 0.03fF
C37820 OR2X1_LOC_18/Y OR2X1_LOC_289/a_8_216# 0.06fF
C37821 AND2X1_LOC_20/a_8_24# OR2X1_LOC_68/B 0.01fF
C37822 OR2X1_LOC_62/B OR2X1_LOC_629/A 0.02fF
C37823 AND2X1_LOC_656/Y AND2X1_LOC_361/A 0.07fF
C37824 OR2X1_LOC_678/Y AND2X1_LOC_31/Y 0.13fF
C37825 OR2X1_LOC_473/A OR2X1_LOC_130/A 0.29fF
C37826 AND2X1_LOC_640/Y AND2X1_LOC_634/Y 0.03fF
C37827 OR2X1_LOC_831/a_8_216# OR2X1_LOC_223/A 0.01fF
C37828 AND2X1_LOC_304/a_8_24# AND2X1_LOC_31/Y 0.01fF
C37829 OR2X1_LOC_87/A AND2X1_LOC_684/a_8_24# 0.02fF
C37830 OR2X1_LOC_634/A OR2X1_LOC_68/B 0.06fF
C37831 AND2X1_LOC_17/Y OR2X1_LOC_639/a_8_216# 0.01fF
C37832 OR2X1_LOC_479/Y OR2X1_LOC_335/B 0.01fF
C37833 AND2X1_LOC_12/Y OR2X1_LOC_205/Y 0.06fF
C37834 OR2X1_LOC_709/a_8_216# AND2X1_LOC_36/Y 0.01fF
C37835 AND2X1_LOC_168/a_8_24# AND2X1_LOC_222/Y 0.01fF
C37836 OR2X1_LOC_426/B OR2X1_LOC_300/a_8_216# 0.01fF
C37837 AND2X1_LOC_64/Y OR2X1_LOC_139/A 0.98fF
C37838 AND2X1_LOC_641/Y D_INPUT_0 0.02fF
C37839 OR2X1_LOC_347/a_8_216# OR2X1_LOC_675/Y 0.04fF
C37840 OR2X1_LOC_291/A D_INPUT_0 0.02fF
C37841 OR2X1_LOC_441/Y OR2X1_LOC_152/A 0.03fF
C37842 OR2X1_LOC_637/a_8_216# AND2X1_LOC_31/Y 0.06fF
C37843 OR2X1_LOC_243/A OR2X1_LOC_598/A 0.04fF
C37844 AND2X1_LOC_464/Y AND2X1_LOC_471/a_8_24# 0.18fF
C37845 OR2X1_LOC_811/A AND2X1_LOC_31/Y 0.11fF
C37846 AND2X1_LOC_634/Y OR2X1_LOC_416/Y 0.58fF
C37847 OR2X1_LOC_47/Y OR2X1_LOC_7/A 0.73fF
C37848 OR2X1_LOC_223/A OR2X1_LOC_787/Y 0.29fF
C37849 AND2X1_LOC_91/B OR2X1_LOC_356/A 0.42fF
C37850 OR2X1_LOC_702/a_8_216# AND2X1_LOC_36/Y 0.01fF
C37851 OR2X1_LOC_78/B OR2X1_LOC_174/Y 0.02fF
C37852 AND2X1_LOC_12/Y OR2X1_LOC_750/Y 0.11fF
C37853 OR2X1_LOC_6/A AND2X1_LOC_228/a_36_24# 0.00fF
C37854 OR2X1_LOC_340/Y OR2X1_LOC_228/Y 0.01fF
C37855 VDD OR2X1_LOC_622/B 0.00fF
C37856 OR2X1_LOC_269/B OR2X1_LOC_451/B 0.00fF
C37857 AND2X1_LOC_554/Y AND2X1_LOC_657/A 0.47fF
C37858 OR2X1_LOC_269/B OR2X1_LOC_512/a_36_216# 0.00fF
C37859 AND2X1_LOC_358/Y AND2X1_LOC_364/a_8_24# 0.00fF
C37860 OR2X1_LOC_151/A OR2X1_LOC_554/a_8_216# 0.05fF
C37861 AND2X1_LOC_40/Y OR2X1_LOC_303/B 0.03fF
C37862 OR2X1_LOC_739/B OR2X1_LOC_739/a_8_216# 0.07fF
C37863 OR2X1_LOC_474/a_8_216# AND2X1_LOC_47/Y 0.01fF
C37864 AND2X1_LOC_338/Y AND2X1_LOC_338/A 0.92fF
C37865 OR2X1_LOC_516/Y OR2X1_LOC_51/Y 0.03fF
C37866 OR2X1_LOC_130/A OR2X1_LOC_228/Y 0.17fF
C37867 AND2X1_LOC_44/Y AND2X1_LOC_279/a_8_24# 0.01fF
C37868 OR2X1_LOC_3/Y AND2X1_LOC_792/Y 0.10fF
C37869 OR2X1_LOC_859/A AND2X1_LOC_47/Y 0.01fF
C37870 OR2X1_LOC_529/Y OR2X1_LOC_419/Y 0.03fF
C37871 OR2X1_LOC_427/A OR2X1_LOC_437/A 0.28fF
C37872 OR2X1_LOC_45/B OR2X1_LOC_315/a_36_216# 0.00fF
C37873 AND2X1_LOC_472/a_8_24# OR2X1_LOC_46/A 0.01fF
C37874 OR2X1_LOC_87/A OR2X1_LOC_560/A 0.03fF
C37875 OR2X1_LOC_87/A OR2X1_LOC_198/A 0.08fF
C37876 OR2X1_LOC_696/A AND2X1_LOC_391/Y 0.15fF
C37877 OR2X1_LOC_696/A AND2X1_LOC_858/B 4.44fF
C37878 OR2X1_LOC_696/A OR2X1_LOC_91/A 0.22fF
C37879 OR2X1_LOC_693/Y AND2X1_LOC_706/a_8_24# 0.23fF
C37880 VDD OR2X1_LOC_338/A 0.12fF
C37881 OR2X1_LOC_755/A AND2X1_LOC_624/B 0.02fF
C37882 AND2X1_LOC_727/Y AND2X1_LOC_657/Y 0.03fF
C37883 OR2X1_LOC_446/Y OR2X1_LOC_780/B 0.11fF
C37884 AND2X1_LOC_500/B OR2X1_LOC_816/A 0.02fF
C37885 OR2X1_LOC_473/A OR2X1_LOC_62/B 0.00fF
C37886 OR2X1_LOC_485/A AND2X1_LOC_222/Y 0.03fF
C37887 AND2X1_LOC_539/Y OR2X1_LOC_56/A 0.03fF
C37888 OR2X1_LOC_719/A AND2X1_LOC_237/a_36_24# 0.00fF
C37889 OR2X1_LOC_784/a_8_216# AND2X1_LOC_31/Y 0.01fF
C37890 AND2X1_LOC_738/B OR2X1_LOC_680/a_8_216# 0.05fF
C37891 OR2X1_LOC_404/Y AND2X1_LOC_497/a_8_24# 0.02fF
C37892 OR2X1_LOC_188/a_8_216# OR2X1_LOC_858/A 0.12fF
C37893 OR2X1_LOC_585/A OR2X1_LOC_80/A 0.10fF
C37894 OR2X1_LOC_825/a_8_216# OR2X1_LOC_749/a_8_216# 0.47fF
C37895 OR2X1_LOC_188/Y AND2X1_LOC_92/Y 0.02fF
C37896 AND2X1_LOC_242/B OR2X1_LOC_59/Y 0.05fF
C37897 OR2X1_LOC_280/Y AND2X1_LOC_657/A 0.02fF
C37898 OR2X1_LOC_169/B OR2X1_LOC_777/B 0.14fF
C37899 OR2X1_LOC_462/a_8_216# OR2X1_LOC_598/A -0.00fF
C37900 AND2X1_LOC_851/B OR2X1_LOC_31/Y 0.01fF
C37901 AND2X1_LOC_383/a_8_24# OR2X1_LOC_91/A 0.09fF
C37902 AND2X1_LOC_866/A AND2X1_LOC_663/a_8_24# 0.04fF
C37903 OR2X1_LOC_186/Y VDD 0.86fF
C37904 AND2X1_LOC_22/Y AND2X1_LOC_24/a_8_24# 0.03fF
C37905 OR2X1_LOC_240/a_8_216# AND2X1_LOC_36/Y 0.01fF
C37906 OR2X1_LOC_739/A AND2X1_LOC_36/Y 0.03fF
C37907 OR2X1_LOC_644/a_8_216# OR2X1_LOC_644/A 0.47fF
C37908 VDD OR2X1_LOC_281/Y -0.00fF
C37909 AND2X1_LOC_363/A OR2X1_LOC_437/A 0.22fF
C37910 VDD OR2X1_LOC_13/a_8_216# 0.21fF
C37911 OR2X1_LOC_45/B OR2X1_LOC_697/a_8_216# 0.01fF
C37912 VDD OR2X1_LOC_584/Y 0.08fF
C37913 OR2X1_LOC_696/A OR2X1_LOC_823/a_8_216# 0.01fF
C37914 INPUT_0 OR2X1_LOC_548/B 0.01fF
C37915 OR2X1_LOC_604/A OR2X1_LOC_6/B 0.09fF
C37916 OR2X1_LOC_160/B OR2X1_LOC_307/A 0.03fF
C37917 OR2X1_LOC_482/a_8_216# AND2X1_LOC_658/A 0.01fF
C37918 VDD OR2X1_LOC_726/A 0.06fF
C37919 AND2X1_LOC_64/Y OR2X1_LOC_324/A 0.01fF
C37920 OR2X1_LOC_154/A OR2X1_LOC_844/B 0.05fF
C37921 VDD OR2X1_LOC_253/Y 0.04fF
C37922 OR2X1_LOC_696/A AND2X1_LOC_573/A 0.07fF
C37923 OR2X1_LOC_178/Y OR2X1_LOC_158/A 0.01fF
C37924 OR2X1_LOC_516/Y OR2X1_LOC_680/A 1.44fF
C37925 OR2X1_LOC_6/B OR2X1_LOC_66/A 0.35fF
C37926 AND2X1_LOC_90/a_8_24# OR2X1_LOC_235/B 0.02fF
C37927 AND2X1_LOC_26/a_8_24# AND2X1_LOC_36/Y 0.01fF
C37928 OR2X1_LOC_111/a_36_216# OR2X1_LOC_109/Y 0.00fF
C37929 AND2X1_LOC_93/a_8_24# AND2X1_LOC_92/Y 0.11fF
C37930 AND2X1_LOC_709/a_8_24# OR2X1_LOC_600/A 0.01fF
C37931 OR2X1_LOC_31/Y OR2X1_LOC_595/Y 0.01fF
C37932 OR2X1_LOC_269/B AND2X1_LOC_36/Y 1.00fF
C37933 AND2X1_LOC_53/Y AND2X1_LOC_52/Y 0.11fF
C37934 OR2X1_LOC_22/Y AND2X1_LOC_657/A 0.07fF
C37935 OR2X1_LOC_52/B AND2X1_LOC_449/a_36_24# 0.01fF
C37936 OR2X1_LOC_705/Y OR2X1_LOC_732/A 0.01fF
C37937 OR2X1_LOC_703/A OR2X1_LOC_486/Y 0.03fF
C37938 OR2X1_LOC_154/A OR2X1_LOC_390/B 0.76fF
C37939 AND2X1_LOC_335/Y AND2X1_LOC_352/B 0.00fF
C37940 OR2X1_LOC_92/Y AND2X1_LOC_774/A 0.10fF
C37941 OR2X1_LOC_265/Y OR2X1_LOC_171/Y 0.07fF
C37942 AND2X1_LOC_91/B AND2X1_LOC_43/B 0.07fF
C37943 AND2X1_LOC_81/B OR2X1_LOC_502/Y 0.01fF
C37944 OR2X1_LOC_829/Y OR2X1_LOC_13/B 0.01fF
C37945 VDD AND2X1_LOC_161/Y 0.24fF
C37946 AND2X1_LOC_326/B OR2X1_LOC_56/A 0.03fF
C37947 OR2X1_LOC_158/A OR2X1_LOC_256/Y 0.10fF
C37948 AND2X1_LOC_301/a_8_24# AND2X1_LOC_219/Y 0.01fF
C37949 OR2X1_LOC_541/a_36_216# OR2X1_LOC_121/A 0.00fF
C37950 OR2X1_LOC_600/A AND2X1_LOC_296/a_36_24# 0.00fF
C37951 OR2X1_LOC_26/Y OR2X1_LOC_525/a_8_216# 0.01fF
C37952 AND2X1_LOC_341/a_8_24# OR2X1_LOC_619/Y 0.04fF
C37953 AND2X1_LOC_337/a_36_24# OR2X1_LOC_56/A 0.01fF
C37954 OR2X1_LOC_790/B OR2X1_LOC_207/B 0.03fF
C37955 OR2X1_LOC_220/B OR2X1_LOC_550/A 0.01fF
C37956 OR2X1_LOC_364/A OR2X1_LOC_390/a_8_216# 0.40fF
C37957 OR2X1_LOC_632/A OR2X1_LOC_161/B 0.03fF
C37958 OR2X1_LOC_109/Y OR2X1_LOC_373/Y 0.45fF
C37959 AND2X1_LOC_361/A AND2X1_LOC_772/Y 0.10fF
C37960 OR2X1_LOC_604/A OR2X1_LOC_441/Y 0.03fF
C37961 OR2X1_LOC_231/B OR2X1_LOC_160/A 0.04fF
C37962 AND2X1_LOC_773/Y OR2X1_LOC_316/Y 0.03fF
C37963 OR2X1_LOC_680/A OR2X1_LOC_373/a_8_216# 0.02fF
C37964 OR2X1_LOC_600/A OR2X1_LOC_517/A 0.03fF
C37965 OR2X1_LOC_494/A AND2X1_LOC_348/Y 0.12fF
C37966 AND2X1_LOC_95/Y OR2X1_LOC_390/A 0.03fF
C37967 OR2X1_LOC_653/B OR2X1_LOC_405/A 0.03fF
C37968 AND2X1_LOC_216/A OR2X1_LOC_67/Y 0.02fF
C37969 AND2X1_LOC_471/Y OR2X1_LOC_56/A 0.04fF
C37970 OR2X1_LOC_809/B OR2X1_LOC_538/A 0.03fF
C37971 OR2X1_LOC_242/a_36_216# OR2X1_LOC_78/A 0.02fF
C37972 OR2X1_LOC_121/Y OR2X1_LOC_160/A 0.07fF
C37973 AND2X1_LOC_173/a_8_24# AND2X1_LOC_110/Y 0.01fF
C37974 AND2X1_LOC_364/Y OR2X1_LOC_744/A 0.07fF
C37975 VDD OR2X1_LOC_862/A 0.13fF
C37976 OR2X1_LOC_856/B OR2X1_LOC_648/B 0.10fF
C37977 AND2X1_LOC_370/a_8_24# AND2X1_LOC_784/A 0.04fF
C37978 OR2X1_LOC_494/A OR2X1_LOC_753/A 0.00fF
C37979 OR2X1_LOC_269/a_36_216# OR2X1_LOC_549/A 0.00fF
C37980 AND2X1_LOC_40/Y OR2X1_LOC_542/B 0.03fF
C37981 AND2X1_LOC_317/a_8_24# OR2X1_LOC_12/Y 0.01fF
C37982 AND2X1_LOC_737/Y VDD 0.34fF
C37983 AND2X1_LOC_12/Y OR2X1_LOC_851/B 0.03fF
C37984 OR2X1_LOC_594/a_8_216# AND2X1_LOC_469/B 0.47fF
C37985 AND2X1_LOC_562/B OR2X1_LOC_816/Y 0.09fF
C37986 OR2X1_LOC_78/A OR2X1_LOC_708/Y 0.01fF
C37987 OR2X1_LOC_656/B OR2X1_LOC_641/A 0.07fF
C37988 OR2X1_LOC_135/a_8_216# OR2X1_LOC_36/Y 0.01fF
C37989 AND2X1_LOC_512/Y INPUT_0 0.01fF
C37990 AND2X1_LOC_358/Y OR2X1_LOC_43/A 0.00fF
C37991 AND2X1_LOC_7/Y AND2X1_LOC_41/Y 0.02fF
C37992 OR2X1_LOC_165/a_8_216# VDD 0.21fF
C37993 OR2X1_LOC_154/A OR2X1_LOC_840/a_8_216# 0.01fF
C37994 OR2X1_LOC_160/B OR2X1_LOC_560/a_8_216# 0.02fF
C37995 AND2X1_LOC_573/A OR2X1_LOC_131/a_36_216# 0.01fF
C37996 OR2X1_LOC_523/Y OR2X1_LOC_66/A 0.36fF
C37997 VDD OR2X1_LOC_394/Y 0.05fF
C37998 AND2X1_LOC_648/B OR2X1_LOC_589/Y 0.01fF
C37999 AND2X1_LOC_146/a_8_24# AND2X1_LOC_36/Y 0.09fF
C38000 AND2X1_LOC_181/Y OR2X1_LOC_6/A 0.03fF
C38001 OR2X1_LOC_160/A OR2X1_LOC_114/B 0.01fF
C38002 OR2X1_LOC_673/B AND2X1_LOC_8/Y 0.00fF
C38003 OR2X1_LOC_188/Y AND2X1_LOC_183/a_8_24# 0.01fF
C38004 AND2X1_LOC_554/Y VDD 0.23fF
C38005 AND2X1_LOC_378/a_8_24# OR2X1_LOC_689/A 0.00fF
C38006 OR2X1_LOC_600/A AND2X1_LOC_624/A 0.32fF
C38007 OR2X1_LOC_743/A AND2X1_LOC_407/a_8_24# 0.11fF
C38008 AND2X1_LOC_352/B OR2X1_LOC_619/Y 0.04fF
C38009 AND2X1_LOC_50/Y AND2X1_LOC_51/a_8_24# 0.11fF
C38010 AND2X1_LOC_851/a_8_24# OR2X1_LOC_427/A 0.02fF
C38011 OR2X1_LOC_773/B VDD 0.21fF
C38012 AND2X1_LOC_56/B OR2X1_LOC_515/A 0.02fF
C38013 OR2X1_LOC_695/a_8_216# OR2X1_LOC_91/A 0.02fF
C38014 OR2X1_LOC_684/a_36_216# AND2X1_LOC_452/Y 0.00fF
C38015 AND2X1_LOC_787/A AND2X1_LOC_578/A 0.03fF
C38016 AND2X1_LOC_707/Y OR2X1_LOC_70/Y 0.02fF
C38017 OR2X1_LOC_598/Y AND2X1_LOC_56/B 0.06fF
C38018 OR2X1_LOC_279/a_36_216# AND2X1_LOC_244/A 0.00fF
C38019 OR2X1_LOC_254/a_8_216# OR2X1_LOC_563/A 0.03fF
C38020 AND2X1_LOC_468/B AND2X1_LOC_469/B 0.04fF
C38021 AND2X1_LOC_653/B AND2X1_LOC_436/Y 0.01fF
C38022 AND2X1_LOC_631/Y OR2X1_LOC_816/A 0.91fF
C38023 OR2X1_LOC_9/Y OR2X1_LOC_670/Y 0.01fF
C38024 OR2X1_LOC_438/Y AND2X1_LOC_544/a_8_24# 0.01fF
C38025 OR2X1_LOC_185/A OR2X1_LOC_78/A 0.47fF
C38026 AND2X1_LOC_59/Y OR2X1_LOC_640/Y 0.01fF
C38027 AND2X1_LOC_729/Y OR2X1_LOC_600/Y 0.05fF
C38028 OR2X1_LOC_154/A OR2X1_LOC_389/A 0.02fF
C38029 AND2X1_LOC_81/B VDD 0.57fF
C38030 OR2X1_LOC_235/B OR2X1_LOC_278/Y 0.03fF
C38031 OR2X1_LOC_188/Y AND2X1_LOC_666/a_36_24# 0.00fF
C38032 OR2X1_LOC_185/A D_GATE_741 0.03fF
C38033 OR2X1_LOC_579/B OR2X1_LOC_66/A 0.01fF
C38034 OR2X1_LOC_405/Y AND2X1_LOC_92/Y 0.04fF
C38035 AND2X1_LOC_3/Y OR2X1_LOC_346/A 0.01fF
C38036 VDD OR2X1_LOC_358/B 0.15fF
C38037 AND2X1_LOC_535/Y AND2X1_LOC_854/a_8_24# 0.03fF
C38038 OR2X1_LOC_235/B OR2X1_LOC_38/a_8_216# -0.02fF
C38039 AND2X1_LOC_866/A OR2X1_LOC_759/Y 0.03fF
C38040 OR2X1_LOC_160/A OR2X1_LOC_538/A 0.03fF
C38041 AND2X1_LOC_733/Y AND2X1_LOC_468/B 0.91fF
C38042 AND2X1_LOC_51/Y OR2X1_LOC_34/a_8_216# 0.01fF
C38043 AND2X1_LOC_712/a_8_24# OR2X1_LOC_417/Y 0.04fF
C38044 OR2X1_LOC_52/a_36_216# OR2X1_LOC_16/A 0.00fF
C38045 VDD OR2X1_LOC_477/B 0.05fF
C38046 OR2X1_LOC_660/Y OR2X1_LOC_130/A 0.02fF
C38047 OR2X1_LOC_8/Y OR2X1_LOC_248/Y 0.03fF
C38048 AND2X1_LOC_351/a_8_24# AND2X1_LOC_333/a_8_24# 0.23fF
C38049 OR2X1_LOC_8/Y OR2X1_LOC_6/a_8_216# 0.02fF
C38050 OR2X1_LOC_158/A OR2X1_LOC_258/Y 0.01fF
C38051 OR2X1_LOC_643/a_8_216# AND2X1_LOC_18/Y 0.06fF
C38052 AND2X1_LOC_772/B AND2X1_LOC_560/B 0.01fF
C38053 AND2X1_LOC_732/B OR2X1_LOC_7/A 0.01fF
C38054 OR2X1_LOC_638/a_8_216# AND2X1_LOC_43/B 0.03fF
C38055 OR2X1_LOC_604/A OR2X1_LOC_529/Y 0.03fF
C38056 OR2X1_LOC_814/A OR2X1_LOC_474/B 0.01fF
C38057 OR2X1_LOC_761/Y AND2X1_LOC_801/a_8_24# 0.23fF
C38058 OR2X1_LOC_856/B AND2X1_LOC_173/a_36_24# 0.01fF
C38059 OR2X1_LOC_40/Y AND2X1_LOC_548/a_8_24# 0.17fF
C38060 AND2X1_LOC_544/a_8_24# AND2X1_LOC_621/Y 0.03fF
C38061 VDD AND2X1_LOC_356/B 0.07fF
C38062 OR2X1_LOC_311/Y AND2X1_LOC_809/a_8_24# 0.01fF
C38063 AND2X1_LOC_59/Y OR2X1_LOC_216/A 0.13fF
C38064 OR2X1_LOC_427/Y AND2X1_LOC_450/a_8_24# 0.04fF
C38065 VDD OR2X1_LOC_280/Y 0.39fF
C38066 OR2X1_LOC_507/a_8_216# OR2X1_LOC_510/Y 0.40fF
C38067 AND2X1_LOC_94/Y OR2X1_LOC_83/A 0.10fF
C38068 OR2X1_LOC_91/Y OR2X1_LOC_164/Y 0.10fF
C38069 OR2X1_LOC_46/A OR2X1_LOC_16/A 0.18fF
C38070 AND2X1_LOC_22/Y AND2X1_LOC_7/Y 0.01fF
C38071 OR2X1_LOC_57/Y OR2X1_LOC_44/Y 0.02fF
C38072 AND2X1_LOC_677/a_36_24# OR2X1_LOC_161/B 0.01fF
C38073 OR2X1_LOC_644/B AND2X1_LOC_41/A 0.01fF
C38074 AND2X1_LOC_592/Y OR2X1_LOC_64/Y 0.01fF
C38075 OR2X1_LOC_51/Y OR2X1_LOC_47/a_8_216# 0.01fF
C38076 OR2X1_LOC_3/Y AND2X1_LOC_707/a_8_24# 0.01fF
C38077 AND2X1_LOC_508/A OR2X1_LOC_44/Y 0.03fF
C38078 OR2X1_LOC_45/a_8_216# OR2X1_LOC_48/B 0.01fF
C38079 AND2X1_LOC_51/Y OR2X1_LOC_772/A 0.01fF
C38080 AND2X1_LOC_485/a_36_24# OR2X1_LOC_209/A 0.01fF
C38081 OR2X1_LOC_252/Y AND2X1_LOC_805/Y 0.20fF
C38082 OR2X1_LOC_474/a_36_216# OR2X1_LOC_113/B 0.00fF
C38083 OR2X1_LOC_216/Y OR2X1_LOC_502/A 0.07fF
C38084 OR2X1_LOC_51/Y AND2X1_LOC_651/B 0.01fF
C38085 OR2X1_LOC_488/Y AND2X1_LOC_489/a_8_24# 0.00fF
C38086 AND2X1_LOC_31/Y OR2X1_LOC_777/B 0.12fF
C38087 AND2X1_LOC_388/Y AND2X1_LOC_727/A 0.01fF
C38088 AND2X1_LOC_40/Y AND2X1_LOC_56/B 1.10fF
C38089 OR2X1_LOC_18/Y OR2X1_LOC_45/a_8_216# 0.02fF
C38090 OR2X1_LOC_402/a_8_216# OR2X1_LOC_78/A 0.01fF
C38091 OR2X1_LOC_70/A D_INPUT_6 1.10fF
C38092 OR2X1_LOC_666/A OR2X1_LOC_279/Y 0.24fF
C38093 AND2X1_LOC_858/a_8_24# AND2X1_LOC_621/Y 0.03fF
C38094 AND2X1_LOC_621/Y AND2X1_LOC_622/a_8_24# 0.03fF
C38095 AND2X1_LOC_42/B OR2X1_LOC_78/B 0.07fF
C38096 AND2X1_LOC_573/A AND2X1_LOC_474/a_8_24# 0.01fF
C38097 OR2X1_LOC_290/a_36_216# OR2X1_LOC_585/A 0.02fF
C38098 AND2X1_LOC_12/Y OR2X1_LOC_160/A 0.21fF
C38099 AND2X1_LOC_40/Y AND2X1_LOC_8/Y 0.06fF
C38100 OR2X1_LOC_435/Y OR2X1_LOC_78/A 0.04fF
C38101 AND2X1_LOC_367/A OR2X1_LOC_485/A 0.18fF
C38102 OR2X1_LOC_184/Y AND2X1_LOC_242/B 0.06fF
C38103 OR2X1_LOC_784/Y OR2X1_LOC_779/a_8_216# 0.02fF
C38104 OR2X1_LOC_176/a_8_216# OR2X1_LOC_47/Y 0.01fF
C38105 AND2X1_LOC_348/Y OR2X1_LOC_427/A 0.05fF
C38106 OR2X1_LOC_798/Y OR2X1_LOC_574/A 0.01fF
C38107 OR2X1_LOC_790/B OR2X1_LOC_790/a_8_216# 0.01fF
C38108 AND2X1_LOC_848/a_8_24# AND2X1_LOC_848/Y 0.01fF
C38109 OR2X1_LOC_48/B OR2X1_LOC_44/Y 2.73fF
C38110 AND2X1_LOC_113/a_36_24# OR2X1_LOC_26/Y 0.01fF
C38111 VDD OR2X1_LOC_196/B 0.26fF
C38112 OR2X1_LOC_779/Y OR2X1_LOC_779/A 0.01fF
C38113 OR2X1_LOC_308/Y OR2X1_LOC_779/B 0.01fF
C38114 OR2X1_LOC_744/A OR2X1_LOC_762/a_8_216# 0.01fF
C38115 OR2X1_LOC_815/a_8_216# OR2X1_LOC_815/A 0.47fF
C38116 VDD OR2X1_LOC_22/Y 0.95fF
C38117 OR2X1_LOC_427/A OR2X1_LOC_753/A 0.14fF
C38118 OR2X1_LOC_47/Y OR2X1_LOC_753/a_8_216# 0.00fF
C38119 OR2X1_LOC_18/Y OR2X1_LOC_44/Y 10.92fF
C38120 OR2X1_LOC_404/A AND2X1_LOC_18/Y 0.18fF
C38121 OR2X1_LOC_185/Y OR2X1_LOC_377/A 0.02fF
C38122 OR2X1_LOC_91/A AND2X1_LOC_663/B 0.07fF
C38123 OR2X1_LOC_18/Y AND2X1_LOC_288/a_8_24# 0.01fF
C38124 VDD AND2X1_LOC_692/a_8_24# -0.00fF
C38125 OR2X1_LOC_468/A AND2X1_LOC_165/a_8_24# 0.01fF
C38126 AND2X1_LOC_119/a_8_24# OR2X1_LOC_78/A 0.17fF
C38127 AND2X1_LOC_168/a_8_24# OR2X1_LOC_74/A 0.04fF
C38128 AND2X1_LOC_811/B OR2X1_LOC_52/B 0.59fF
C38129 OR2X1_LOC_479/Y OR2X1_LOC_776/a_36_216# 0.00fF
C38130 AND2X1_LOC_42/B OR2X1_LOC_721/Y 0.07fF
C38131 AND2X1_LOC_59/Y OR2X1_LOC_468/Y 0.02fF
C38132 AND2X1_LOC_228/Y OR2X1_LOC_6/A 0.01fF
C38133 OR2X1_LOC_377/A AND2X1_LOC_412/a_8_24# 0.02fF
C38134 AND2X1_LOC_729/Y OR2X1_LOC_591/A 0.01fF
C38135 AND2X1_LOC_477/A AND2X1_LOC_436/Y 0.03fF
C38136 OR2X1_LOC_158/A AND2X1_LOC_318/Y 0.10fF
C38137 OR2X1_LOC_151/A OR2X1_LOC_506/B 0.03fF
C38138 OR2X1_LOC_527/Y OR2X1_LOC_164/Y 0.13fF
C38139 OR2X1_LOC_427/A OR2X1_LOC_754/a_8_216# 0.01fF
C38140 OR2X1_LOC_185/A OR2X1_LOC_155/A 0.05fF
C38141 AND2X1_LOC_512/Y OR2X1_LOC_64/Y 0.07fF
C38142 AND2X1_LOC_722/a_36_24# OR2X1_LOC_417/A 0.01fF
C38143 OR2X1_LOC_95/Y AND2X1_LOC_500/B 0.01fF
C38144 INPUT_0 OR2X1_LOC_54/Y 4.71fF
C38145 OR2X1_LOC_625/Y OR2X1_LOC_7/A 0.30fF
C38146 OR2X1_LOC_610/a_8_216# OR2X1_LOC_647/A 0.39fF
C38147 OR2X1_LOC_235/B OR2X1_LOC_19/B 0.10fF
C38148 OR2X1_LOC_74/A AND2X1_LOC_808/a_8_24# 0.04fF
C38149 AND2X1_LOC_568/B AND2X1_LOC_863/Y 0.01fF
C38150 OR2X1_LOC_756/B AND2X1_LOC_27/a_8_24# 0.01fF
C38151 OR2X1_LOC_510/Y OR2X1_LOC_124/Y 0.18fF
C38152 OR2X1_LOC_45/Y OR2X1_LOC_3/Y 1.18fF
C38153 AND2X1_LOC_47/Y OR2X1_LOC_66/A 6.92fF
C38154 OR2X1_LOC_185/Y OR2X1_LOC_203/Y 0.10fF
C38155 AND2X1_LOC_571/Y AND2X1_LOC_489/Y 0.00fF
C38156 OR2X1_LOC_460/B AND2X1_LOC_3/Y 0.03fF
C38157 AND2X1_LOC_3/Y OR2X1_LOC_161/A 0.23fF
C38158 D_INPUT_0 AND2X1_LOC_92/Y 6.40fF
C38159 AND2X1_LOC_8/Y OR2X1_LOC_87/Y 0.08fF
C38160 OR2X1_LOC_154/A OR2X1_LOC_403/B 0.05fF
C38161 AND2X1_LOC_31/Y OR2X1_LOC_831/B 0.03fF
C38162 OR2X1_LOC_70/Y AND2X1_LOC_841/B 0.17fF
C38163 OR2X1_LOC_841/A AND2X1_LOC_47/Y 0.01fF
C38164 AND2X1_LOC_191/B OR2X1_LOC_226/a_36_216# 0.01fF
C38165 OR2X1_LOC_786/Y AND2X1_LOC_262/a_8_24# 0.01fF
C38166 OR2X1_LOC_18/Y AND2X1_LOC_116/Y 0.01fF
C38167 OR2X1_LOC_6/B OR2X1_LOC_84/A 0.02fF
C38168 OR2X1_LOC_814/A OR2X1_LOC_561/Y 0.00fF
C38169 AND2X1_LOC_729/Y OR2X1_LOC_420/a_36_216# 0.00fF
C38170 OR2X1_LOC_405/A OR2X1_LOC_216/a_36_216# 0.00fF
C38171 OR2X1_LOC_18/Y OR2X1_LOC_20/a_8_216# 0.01fF
C38172 OR2X1_LOC_251/Y AND2X1_LOC_286/Y 0.01fF
C38173 OR2X1_LOC_127/a_36_216# OR2X1_LOC_3/Y 0.03fF
C38174 OR2X1_LOC_502/A OR2X1_LOC_647/a_8_216# 0.01fF
C38175 AND2X1_LOC_348/Y AND2X1_LOC_363/A 0.00fF
C38176 OR2X1_LOC_585/A OR2X1_LOC_6/A 0.45fF
C38177 OR2X1_LOC_822/a_8_216# OR2X1_LOC_47/Y 0.01fF
C38178 OR2X1_LOC_864/A OR2X1_LOC_649/B 0.00fF
C38179 AND2X1_LOC_12/Y OR2X1_LOC_33/a_8_216# 0.01fF
C38180 INPUT_5 AND2X1_LOC_11/a_8_24# 0.11fF
C38181 AND2X1_LOC_59/Y OR2X1_LOC_675/a_8_216# 0.01fF
C38182 AND2X1_LOC_580/A OR2X1_LOC_89/A 0.07fF
C38183 AND2X1_LOC_42/B OR2X1_LOC_375/A 0.29fF
C38184 AND2X1_LOC_363/A OR2X1_LOC_753/A 0.01fF
C38185 OR2X1_LOC_643/A OR2X1_LOC_810/A 0.05fF
C38186 AND2X1_LOC_41/A AND2X1_LOC_53/Y 0.02fF
C38187 OR2X1_LOC_40/Y OR2X1_LOC_3/B 0.01fF
C38188 VDD OR2X1_LOC_112/B 0.17fF
C38189 AND2X1_LOC_70/Y AND2X1_LOC_109/a_8_24# 0.01fF
C38190 AND2X1_LOC_658/B OR2X1_LOC_615/Y 0.00fF
C38191 AND2X1_LOC_624/B OR2X1_LOC_253/Y 0.07fF
C38192 OR2X1_LOC_427/A OR2X1_LOC_684/Y 0.01fF
C38193 AND2X1_LOC_514/Y AND2X1_LOC_841/B 0.07fF
C38194 OR2X1_LOC_151/A OR2X1_LOC_247/Y 0.02fF
C38195 OR2X1_LOC_429/Y OR2X1_LOC_25/a_8_216# 0.41fF
C38196 VDD AND2X1_LOC_808/A 0.36fF
C38197 OR2X1_LOC_280/a_8_216# OR2X1_LOC_26/Y 0.01fF
C38198 AND2X1_LOC_663/B AND2X1_LOC_573/A 0.10fF
C38199 AND2X1_LOC_674/a_8_24# OR2X1_LOC_805/A 0.04fF
C38200 OR2X1_LOC_375/A OR2X1_LOC_705/Y 0.01fF
C38201 AND2X1_LOC_91/B OR2X1_LOC_558/A 0.01fF
C38202 AND2X1_LOC_95/Y OR2X1_LOC_750/A 0.03fF
C38203 AND2X1_LOC_738/a_8_24# AND2X1_LOC_808/A 0.20fF
C38204 AND2X1_LOC_42/a_36_24# OR2X1_LOC_83/A 0.00fF
C38205 OR2X1_LOC_633/A OR2X1_LOC_68/B 0.04fF
C38206 AND2X1_LOC_702/Y OR2X1_LOC_321/Y 0.01fF
C38207 AND2X1_LOC_42/a_8_24# OR2X1_LOC_240/A 0.06fF
C38208 OR2X1_LOC_22/Y OR2X1_LOC_829/a_8_216# 0.01fF
C38209 OR2X1_LOC_377/A OR2X1_LOC_472/B 0.07fF
C38210 OR2X1_LOC_160/B OR2X1_LOC_512/a_8_216# 0.00fF
C38211 AND2X1_LOC_427/a_36_24# OR2X1_LOC_161/B 0.01fF
C38212 OR2X1_LOC_22/Y AND2X1_LOC_274/a_8_24# 0.01fF
C38213 VDD OR2X1_LOC_66/Y 0.19fF
C38214 AND2X1_LOC_70/Y OR2X1_LOC_66/a_8_216# 0.01fF
C38215 OR2X1_LOC_427/A AND2X1_LOC_845/Y 0.07fF
C38216 AND2X1_LOC_456/Y OR2X1_LOC_485/A 0.08fF
C38217 OR2X1_LOC_74/A AND2X1_LOC_474/Y 0.03fF
C38218 OR2X1_LOC_472/B AND2X1_LOC_824/B 0.29fF
C38219 AND2X1_LOC_355/a_8_24# AND2X1_LOC_390/B 0.01fF
C38220 VDD OR2X1_LOC_387/a_8_216# 0.00fF
C38221 OR2X1_LOC_66/A OR2X1_LOC_598/A 0.11fF
C38222 OR2X1_LOC_485/A OR2X1_LOC_74/A 0.12fF
C38223 AND2X1_LOC_76/a_8_24# OR2X1_LOC_31/Y 0.01fF
C38224 OR2X1_LOC_161/B OR2X1_LOC_71/A 0.01fF
C38225 AND2X1_LOC_328/a_8_24# OR2X1_LOC_651/A -0.03fF
C38226 OR2X1_LOC_32/Y OR2X1_LOC_27/Y 0.00fF
C38227 OR2X1_LOC_686/A AND2X1_LOC_31/Y 0.02fF
C38228 OR2X1_LOC_624/B AND2X1_LOC_79/Y 0.01fF
C38229 OR2X1_LOC_380/A OR2X1_LOC_22/A 0.41fF
C38230 OR2X1_LOC_443/Y OR2X1_LOC_87/A 0.00fF
C38231 AND2X1_LOC_59/Y OR2X1_LOC_655/B 0.03fF
C38232 OR2X1_LOC_64/Y AND2X1_LOC_105/a_8_24# 0.01fF
C38233 OR2X1_LOC_682/Y OR2X1_LOC_64/Y 0.01fF
C38234 OR2X1_LOC_377/A OR2X1_LOC_852/A 0.02fF
C38235 OR2X1_LOC_405/A OR2X1_LOC_218/Y 0.11fF
C38236 AND2X1_LOC_268/a_8_24# OR2X1_LOC_549/A 0.02fF
C38237 AND2X1_LOC_3/Y AND2X1_LOC_51/Y 0.12fF
C38238 AND2X1_LOC_76/Y AND2X1_LOC_660/A 0.03fF
C38239 OR2X1_LOC_468/a_8_216# OR2X1_LOC_506/A 0.02fF
C38240 AND2X1_LOC_161/Y OR2X1_LOC_163/Y 0.02fF
C38241 OR2X1_LOC_437/A OR2X1_LOC_322/a_8_216# 0.15fF
C38242 OR2X1_LOC_358/a_8_216# OR2X1_LOC_532/B 0.01fF
C38243 AND2X1_LOC_149/a_8_24# AND2X1_LOC_797/A 0.01fF
C38244 OR2X1_LOC_852/A AND2X1_LOC_824/B 0.00fF
C38245 OR2X1_LOC_502/A OR2X1_LOC_396/Y 0.03fF
C38246 AND2X1_LOC_41/A OR2X1_LOC_705/B 0.31fF
C38247 AND2X1_LOC_165/a_8_24# OR2X1_LOC_449/B 0.01fF
C38248 OR2X1_LOC_251/Y OR2X1_LOC_22/Y 0.03fF
C38249 AND2X1_LOC_561/B AND2X1_LOC_563/Y 0.01fF
C38250 AND2X1_LOC_59/Y OR2X1_LOC_222/a_8_216# 0.01fF
C38251 OR2X1_LOC_36/Y OR2X1_LOC_71/Y 0.03fF
C38252 AND2X1_LOC_572/A OR2X1_LOC_95/Y 0.03fF
C38253 OR2X1_LOC_862/B OR2X1_LOC_561/B 0.49fF
C38254 AND2X1_LOC_56/B AND2X1_LOC_826/a_8_24# 0.10fF
C38255 AND2X1_LOC_211/B AND2X1_LOC_326/a_8_24# 0.03fF
C38256 OR2X1_LOC_810/A OR2X1_LOC_113/A 0.04fF
C38257 OR2X1_LOC_51/Y OR2X1_LOC_533/A 0.02fF
C38258 AND2X1_LOC_721/A OR2X1_LOC_278/Y 0.04fF
C38259 OR2X1_LOC_446/Y OR2X1_LOC_449/B 0.12fF
C38260 OR2X1_LOC_26/Y OR2X1_LOC_72/a_8_216# 0.01fF
C38261 OR2X1_LOC_709/A OR2X1_LOC_308/Y 1.17fF
C38262 OR2X1_LOC_36/Y AND2X1_LOC_201/a_36_24# 0.00fF
C38263 AND2X1_LOC_838/Y AND2X1_LOC_838/B 0.00fF
C38264 OR2X1_LOC_26/Y AND2X1_LOC_476/A 0.11fF
C38265 AND2X1_LOC_72/B OR2X1_LOC_347/B 0.01fF
C38266 OR2X1_LOC_64/Y OR2X1_LOC_54/Y 0.00fF
C38267 OR2X1_LOC_121/Y OR2X1_LOC_130/Y 0.01fF
C38268 AND2X1_LOC_382/a_8_24# D_INPUT_1 0.02fF
C38269 AND2X1_LOC_660/A OR2X1_LOC_52/B 0.07fF
C38270 OR2X1_LOC_36/Y D_INPUT_1 0.05fF
C38271 OR2X1_LOC_87/A OR2X1_LOC_783/a_8_216# 0.05fF
C38272 OR2X1_LOC_269/Y OR2X1_LOC_269/B 0.03fF
C38273 OR2X1_LOC_684/Y AND2X1_LOC_687/B 0.01fF
C38274 OR2X1_LOC_435/A OR2X1_LOC_390/B 0.07fF
C38275 OR2X1_LOC_858/A OR2X1_LOC_735/B 0.02fF
C38276 OR2X1_LOC_3/Y OR2X1_LOC_95/Y 0.03fF
C38277 AND2X1_LOC_578/A AND2X1_LOC_675/A 0.07fF
C38278 OR2X1_LOC_154/A OR2X1_LOC_493/Y 0.28fF
C38279 OR2X1_LOC_532/B OR2X1_LOC_486/B 0.00fF
C38280 OR2X1_LOC_831/a_36_216# OR2X1_LOC_804/A 0.00fF
C38281 OR2X1_LOC_529/Y OR2X1_LOC_224/a_36_216# 0.00fF
C38282 OR2X1_LOC_154/A OR2X1_LOC_801/B 0.07fF
C38283 OR2X1_LOC_244/B OR2X1_LOC_140/Y 0.11fF
C38284 OR2X1_LOC_175/Y AND2X1_LOC_417/a_8_24# 0.03fF
C38285 AND2X1_LOC_631/Y OR2X1_LOC_95/Y 0.03fF
C38286 AND2X1_LOC_334/a_8_24# INPUT_1 0.10fF
C38287 AND2X1_LOC_197/a_8_24# OR2X1_LOC_31/Y 0.01fF
C38288 AND2X1_LOC_70/Y OR2X1_LOC_374/a_36_216# 0.00fF
C38289 AND2X1_LOC_23/a_36_24# OR2X1_LOC_19/B 0.00fF
C38290 OR2X1_LOC_446/Y OR2X1_LOC_121/B 0.72fF
C38291 OR2X1_LOC_22/A OR2X1_LOC_408/a_8_216# 0.41fF
C38292 AND2X1_LOC_70/Y OR2X1_LOC_308/Y 0.03fF
C38293 OR2X1_LOC_516/B OR2X1_LOC_13/B 0.01fF
C38294 AND2X1_LOC_59/Y OR2X1_LOC_750/Y 0.09fF
C38295 OR2X1_LOC_538/A OR2X1_LOC_532/Y 0.00fF
C38296 OR2X1_LOC_269/B OR2X1_LOC_196/a_8_216# 0.01fF
C38297 OR2X1_LOC_696/A AND2X1_LOC_724/Y 0.02fF
C38298 AND2X1_LOC_22/Y OR2X1_LOC_390/A 0.03fF
C38299 OR2X1_LOC_140/A OR2X1_LOC_115/B 0.03fF
C38300 OR2X1_LOC_31/a_8_216# OR2X1_LOC_17/Y 0.00fF
C38301 OR2X1_LOC_3/B OR2X1_LOC_44/a_8_216# 0.02fF
C38302 OR2X1_LOC_511/Y AND2X1_LOC_796/A 0.10fF
C38303 OR2X1_LOC_162/A OR2X1_LOC_162/a_8_216# 0.39fF
C38304 AND2X1_LOC_334/a_36_24# AND2X1_LOC_219/A 0.01fF
C38305 OR2X1_LOC_473/A OR2X1_LOC_121/B 0.03fF
C38306 OR2X1_LOC_129/a_36_216# AND2X1_LOC_202/Y 0.00fF
C38307 OR2X1_LOC_703/A OR2X1_LOC_308/Y 0.12fF
C38308 OR2X1_LOC_485/A AND2X1_LOC_647/Y 0.00fF
C38309 OR2X1_LOC_848/A AND2X1_LOC_236/a_8_24# 0.02fF
C38310 AND2X1_LOC_43/B OR2X1_LOC_446/B 0.75fF
C38311 AND2X1_LOC_827/a_8_24# OR2X1_LOC_46/A 0.17fF
C38312 OR2X1_LOC_778/A OR2X1_LOC_493/Y 0.69fF
C38313 OR2X1_LOC_49/A OR2X1_LOC_382/a_8_216# 0.05fF
C38314 OR2X1_LOC_765/a_8_216# OR2X1_LOC_12/Y 0.07fF
C38315 D_INPUT_3 D_INPUT_0 0.18fF
C38316 OR2X1_LOC_96/Y OR2X1_LOC_428/A 0.01fF
C38317 OR2X1_LOC_339/a_8_216# AND2X1_LOC_7/B 0.02fF
C38318 OR2X1_LOC_19/B AND2X1_LOC_721/A 0.02fF
C38319 OR2X1_LOC_113/a_8_216# OR2X1_LOC_244/Y 0.01fF
C38320 OR2X1_LOC_859/A D_INPUT_1 0.06fF
C38321 OR2X1_LOC_474/B OR2X1_LOC_244/Y 0.00fF
C38322 OR2X1_LOC_646/a_8_216# OR2X1_LOC_68/B 0.18fF
C38323 AND2X1_LOC_454/a_8_24# OR2X1_LOC_428/A 0.01fF
C38324 AND2X1_LOC_340/Y AND2X1_LOC_340/a_36_24# 0.00fF
C38325 OR2X1_LOC_22/Y OR2X1_LOC_67/Y 0.08fF
C38326 OR2X1_LOC_329/B AND2X1_LOC_473/Y 1.24fF
C38327 AND2X1_LOC_53/Y OR2X1_LOC_207/a_8_216# 0.03fF
C38328 AND2X1_LOC_47/Y OR2X1_LOC_84/A 0.19fF
C38329 OR2X1_LOC_739/A OR2X1_LOC_469/B 0.03fF
C38330 OR2X1_LOC_833/Y VDD 0.48fF
C38331 OR2X1_LOC_334/B OR2X1_LOC_338/A 0.04fF
C38332 OR2X1_LOC_31/Y OR2X1_LOC_409/Y 0.10fF
C38333 OR2X1_LOC_209/a_8_216# OR2X1_LOC_209/A 0.18fF
C38334 OR2X1_LOC_858/A OR2X1_LOC_161/B 0.03fF
C38335 OR2X1_LOC_151/A AND2X1_LOC_18/Y 0.14fF
C38336 AND2X1_LOC_555/Y AND2X1_LOC_348/A 0.00fF
C38337 OR2X1_LOC_604/A OR2X1_LOC_672/a_8_216# 0.06fF
C38338 OR2X1_LOC_759/A OR2X1_LOC_158/A 0.04fF
C38339 OR2X1_LOC_756/B OR2X1_LOC_139/A 0.03fF
C38340 OR2X1_LOC_40/Y AND2X1_LOC_535/Y 0.06fF
C38341 OR2X1_LOC_646/B OR2X1_LOC_66/A 0.01fF
C38342 OR2X1_LOC_121/B OR2X1_LOC_228/Y 0.17fF
C38343 OR2X1_LOC_850/B OR2X1_LOC_362/a_8_216# 0.01fF
C38344 OR2X1_LOC_45/B AND2X1_LOC_508/A 0.03fF
C38345 OR2X1_LOC_71/Y OR2X1_LOC_419/Y 0.00fF
C38346 AND2X1_LOC_12/Y OR2X1_LOC_130/Y 0.03fF
C38347 AND2X1_LOC_298/a_8_24# OR2X1_LOC_469/B 0.07fF
C38348 OR2X1_LOC_47/Y OR2X1_LOC_615/Y 0.22fF
C38349 OR2X1_LOC_589/A OR2X1_LOC_59/Y 0.08fF
C38350 VDD OR2X1_LOC_485/Y 0.31fF
C38351 OR2X1_LOC_831/A AND2X1_LOC_92/Y 0.07fF
C38352 OR2X1_LOC_429/a_36_216# OR2X1_LOC_70/A 0.00fF
C38353 AND2X1_LOC_654/Y OR2X1_LOC_321/a_8_216# 0.03fF
C38354 OR2X1_LOC_92/Y AND2X1_LOC_786/Y 0.12fF
C38355 OR2X1_LOC_279/Y OR2X1_LOC_13/B 0.02fF
C38356 OR2X1_LOC_158/A OR2X1_LOC_697/a_8_216# 0.07fF
C38357 OR2X1_LOC_441/Y AND2X1_LOC_212/Y 0.07fF
C38358 INPUT_0 OR2X1_LOC_57/a_36_216# 0.03fF
C38359 OR2X1_LOC_744/A AND2X1_LOC_243/Y 0.07fF
C38360 AND2X1_LOC_605/Y OR2X1_LOC_421/Y 0.30fF
C38361 OR2X1_LOC_508/a_8_216# OR2X1_LOC_474/Y 0.05fF
C38362 OR2X1_LOC_31/a_8_216# OR2X1_LOC_588/A 0.40fF
C38363 OR2X1_LOC_87/A OR2X1_LOC_605/Y 0.00fF
C38364 OR2X1_LOC_45/B OR2X1_LOC_48/B 0.30fF
C38365 OR2X1_LOC_624/A AND2X1_LOC_7/B 0.10fF
C38366 AND2X1_LOC_660/A AND2X1_LOC_216/A 0.00fF
C38367 AND2X1_LOC_719/Y AND2X1_LOC_861/B 0.03fF
C38368 OR2X1_LOC_158/A OR2X1_LOC_698/Y 0.02fF
C38369 AND2X1_LOC_392/A AND2X1_LOC_391/Y 0.02fF
C38370 AND2X1_LOC_12/Y OR2X1_LOC_774/a_8_216# 0.01fF
C38371 AND2X1_LOC_392/A OR2X1_LOC_91/A 0.90fF
C38372 OR2X1_LOC_625/Y OR2X1_LOC_753/a_8_216# -0.02fF
C38373 AND2X1_LOC_568/B OR2X1_LOC_744/A 0.03fF
C38374 OR2X1_LOC_641/Y AND2X1_LOC_19/Y 0.07fF
C38375 OR2X1_LOC_158/A D_INPUT_5 0.03fF
C38376 OR2X1_LOC_45/B OR2X1_LOC_18/Y 11.02fF
C38377 OR2X1_LOC_196/Y AND2X1_LOC_12/Y 0.03fF
C38378 AND2X1_LOC_729/Y AND2X1_LOC_724/a_8_24# 0.01fF
C38379 OR2X1_LOC_421/A OR2X1_LOC_762/Y 0.00fF
C38380 AND2X1_LOC_51/Y OR2X1_LOC_576/a_8_216# 0.01fF
C38381 OR2X1_LOC_154/A OR2X1_LOC_390/a_36_216# 0.01fF
C38382 AND2X1_LOC_753/B OR2X1_LOC_596/A 0.07fF
C38383 AND2X1_LOC_847/a_36_24# AND2X1_LOC_789/Y 0.01fF
C38384 AND2X1_LOC_706/Y OR2X1_LOC_432/a_8_216# 0.50fF
C38385 AND2X1_LOC_647/Y OR2X1_LOC_609/Y 0.03fF
C38386 OR2X1_LOC_90/a_8_216# OR2X1_LOC_56/A 0.01fF
C38387 AND2X1_LOC_449/Y OR2X1_LOC_428/A 0.03fF
C38388 OR2X1_LOC_585/A OR2X1_LOC_171/a_36_216# 0.02fF
C38389 AND2X1_LOC_443/Y AND2X1_LOC_469/B 0.00fF
C38390 OR2X1_LOC_6/A OR2X1_LOC_230/Y 0.01fF
C38391 OR2X1_LOC_795/B AND2X1_LOC_92/Y 0.03fF
C38392 OR2X1_LOC_118/Y AND2X1_LOC_249/a_8_24# 0.01fF
C38393 AND2X1_LOC_529/a_36_24# OR2X1_LOC_66/A 0.01fF
C38394 OR2X1_LOC_658/a_8_216# OR2X1_LOC_244/Y 0.01fF
C38395 OR2X1_LOC_656/a_8_216# OR2X1_LOC_771/B 0.35fF
C38396 OR2X1_LOC_139/A OR2X1_LOC_657/a_8_216# 0.03fF
C38397 OR2X1_LOC_358/a_36_216# OR2X1_LOC_97/A 0.00fF
C38398 OR2X1_LOC_297/A OR2X1_LOC_59/Y 0.03fF
C38399 OR2X1_LOC_696/A OR2X1_LOC_371/Y 0.07fF
C38400 AND2X1_LOC_319/a_36_24# OR2X1_LOC_56/A 0.01fF
C38401 AND2X1_LOC_91/B OR2X1_LOC_810/A 0.10fF
C38402 OR2X1_LOC_520/B OR2X1_LOC_771/B 0.60fF
C38403 OR2X1_LOC_316/Y OR2X1_LOC_12/Y 0.06fF
C38404 OR2X1_LOC_764/a_8_216# OR2X1_LOC_44/Y 0.01fF
C38405 OR2X1_LOC_541/A OR2X1_LOC_778/B 0.00fF
C38406 AND2X1_LOC_456/B OR2X1_LOC_666/A 0.02fF
C38407 OR2X1_LOC_405/A OR2X1_LOC_596/A 0.04fF
C38408 OR2X1_LOC_709/A AND2X1_LOC_748/a_36_24# 0.01fF
C38409 OR2X1_LOC_756/B AND2X1_LOC_179/a_8_24# 0.14fF
C38410 AND2X1_LOC_92/a_8_24# OR2X1_LOC_97/B 0.19fF
C38411 OR2X1_LOC_363/B OR2X1_LOC_850/B 0.00fF
C38412 AND2X1_LOC_733/Y AND2X1_LOC_443/Y 0.09fF
C38413 AND2X1_LOC_7/B OR2X1_LOC_552/a_8_216# 0.05fF
C38414 AND2X1_LOC_794/B OR2X1_LOC_39/A 0.10fF
C38415 AND2X1_LOC_547/Y OR2X1_LOC_427/A 0.02fF
C38416 OR2X1_LOC_659/a_8_216# OR2X1_LOC_113/B 0.01fF
C38417 AND2X1_LOC_64/Y OR2X1_LOC_479/Y 2.27fF
C38418 OR2X1_LOC_663/A OR2X1_LOC_78/B 0.07fF
C38419 AND2X1_LOC_464/A OR2X1_LOC_372/Y 0.33fF
C38420 AND2X1_LOC_714/a_8_24# OR2X1_LOC_36/Y 0.01fF
C38421 OR2X1_LOC_26/Y AND2X1_LOC_445/a_8_24# 0.02fF
C38422 AND2X1_LOC_62/a_8_24# OR2X1_LOC_600/A 0.04fF
C38423 OR2X1_LOC_229/a_8_216# OR2X1_LOC_6/A 0.00fF
C38424 AND2X1_LOC_231/a_36_24# OR2X1_LOC_52/B 0.00fF
C38425 AND2X1_LOC_410/a_8_24# OR2X1_LOC_48/B 0.23fF
C38426 OR2X1_LOC_271/Y AND2X1_LOC_786/Y 0.05fF
C38427 OR2X1_LOC_151/A OR2X1_LOC_500/A 0.00fF
C38428 OR2X1_LOC_599/A OR2X1_LOC_16/A 0.04fF
C38429 AND2X1_LOC_110/Y OR2X1_LOC_623/a_36_216# 0.00fF
C38430 AND2X1_LOC_323/a_36_24# OR2X1_LOC_620/Y 0.00fF
C38431 OR2X1_LOC_620/a_8_216# AND2X1_LOC_56/B 0.01fF
C38432 AND2X1_LOC_40/Y AND2X1_LOC_92/Y 0.10fF
C38433 OR2X1_LOC_653/B OR2X1_LOC_653/A 0.11fF
C38434 OR2X1_LOC_663/A AND2X1_LOC_103/a_36_24# 0.00fF
C38435 OR2X1_LOC_866/B OR2X1_LOC_557/A 0.12fF
C38436 AND2X1_LOC_866/B OR2X1_LOC_59/Y 0.11fF
C38437 OR2X1_LOC_599/A AND2X1_LOC_714/a_36_24# 0.00fF
C38438 AND2X1_LOC_705/a_8_24# OR2X1_LOC_48/B 0.03fF
C38439 AND2X1_LOC_578/A AND2X1_LOC_241/a_8_24# 0.00fF
C38440 AND2X1_LOC_654/B OR2X1_LOC_59/Y 0.02fF
C38441 AND2X1_LOC_503/a_8_24# OR2X1_LOC_78/B 0.05fF
C38442 OR2X1_LOC_566/Y OR2X1_LOC_365/B 0.01fF
C38443 OR2X1_LOC_325/A OR2X1_LOC_538/A 0.01fF
C38444 OR2X1_LOC_495/Y OR2X1_LOC_59/Y 0.03fF
C38445 AND2X1_LOC_392/A AND2X1_LOC_573/A 0.07fF
C38446 OR2X1_LOC_262/Y AND2X1_LOC_249/a_8_24# 0.00fF
C38447 OR2X1_LOC_506/A OR2X1_LOC_66/A 0.09fF
C38448 OR2X1_LOC_492/Y OR2X1_LOC_36/Y 0.01fF
C38449 AND2X1_LOC_95/Y OR2X1_LOC_347/Y 0.01fF
C38450 OR2X1_LOC_589/A OR2X1_LOC_433/a_8_216# 0.05fF
C38451 AND2X1_LOC_79/Y OR2X1_LOC_266/A 0.07fF
C38452 AND2X1_LOC_193/a_8_24# AND2X1_LOC_194/Y 0.01fF
C38453 OR2X1_LOC_405/A OR2X1_LOC_493/a_36_216# 0.01fF
C38454 OR2X1_LOC_850/B OR2X1_LOC_756/B 1.68fF
C38455 OR2X1_LOC_160/B OR2X1_LOC_340/Y 0.08fF
C38456 OR2X1_LOC_502/A AND2X1_LOC_41/A 0.13fF
C38457 OR2X1_LOC_841/A OR2X1_LOC_506/A 0.00fF
C38458 OR2X1_LOC_302/B AND2X1_LOC_527/a_8_24# 0.19fF
C38459 OR2X1_LOC_91/Y AND2X1_LOC_784/a_8_24# 0.02fF
C38460 INPUT_0 OR2X1_LOC_689/a_8_216# 0.01fF
C38461 OR2X1_LOC_160/B OR2X1_LOC_707/A 0.01fF
C38462 OR2X1_LOC_40/Y OR2X1_LOC_246/Y 0.16fF
C38463 OR2X1_LOC_709/A AND2X1_LOC_516/a_8_24# 0.01fF
C38464 VDD OR2X1_LOC_39/A 6.30fF
C38465 AND2X1_LOC_809/A AND2X1_LOC_434/Y 0.04fF
C38466 OR2X1_LOC_160/B OR2X1_LOC_130/A 0.21fF
C38467 AND2X1_LOC_539/Y OR2X1_LOC_417/Y 0.03fF
C38468 OR2X1_LOC_7/A OR2X1_LOC_584/a_8_216# 0.02fF
C38469 OR2X1_LOC_574/A AND2X1_LOC_433/a_36_24# 0.06fF
C38470 OR2X1_LOC_710/B OR2X1_LOC_375/A 0.01fF
C38471 OR2X1_LOC_62/A OR2X1_LOC_749/Y 0.09fF
C38472 OR2X1_LOC_298/Y OR2X1_LOC_56/A 0.07fF
C38473 OR2X1_LOC_354/A OR2X1_LOC_854/a_8_216# 0.00fF
C38474 AND2X1_LOC_186/a_8_24# AND2X1_LOC_657/Y 0.14fF
C38475 AND2X1_LOC_553/a_8_24# AND2X1_LOC_560/B 0.02fF
C38476 OR2X1_LOC_508/A OR2X1_LOC_502/A 0.18fF
C38477 AND2X1_LOC_390/B OR2X1_LOC_12/Y 0.02fF
C38478 AND2X1_LOC_539/Y OR2X1_LOC_311/Y 0.01fF
C38479 AND2X1_LOC_779/a_8_24# OR2X1_LOC_697/Y 0.00fF
C38480 AND2X1_LOC_509/Y AND2X1_LOC_621/Y 0.05fF
C38481 OR2X1_LOC_680/A AND2X1_LOC_468/a_8_24# 0.01fF
C38482 AND2X1_LOC_154/a_8_24# AND2X1_LOC_663/A 0.11fF
C38483 AND2X1_LOC_259/Y OR2X1_LOC_382/a_8_216# 0.01fF
C38484 D_INPUT_0 OR2X1_LOC_171/Y 0.08fF
C38485 AND2X1_LOC_42/B OR2X1_LOC_549/A 0.07fF
C38486 OR2X1_LOC_665/Y AND2X1_LOC_254/a_8_24# 0.04fF
C38487 AND2X1_LOC_856/a_8_24# OR2X1_LOC_428/A 0.03fF
C38488 OR2X1_LOC_778/Y OR2X1_LOC_784/B 0.12fF
C38489 OR2X1_LOC_426/B OR2X1_LOC_36/Y 0.68fF
C38490 OR2X1_LOC_421/A OR2X1_LOC_312/Y 0.14fF
C38491 AND2X1_LOC_22/Y OR2X1_LOC_750/A 0.03fF
C38492 OR2X1_LOC_47/Y D_INPUT_6 0.03fF
C38493 AND2X1_LOC_535/Y OR2X1_LOC_7/A 0.03fF
C38494 OR2X1_LOC_51/Y AND2X1_LOC_859/Y 0.19fF
C38495 OR2X1_LOC_770/Y OR2X1_LOC_771/B 0.06fF
C38496 OR2X1_LOC_70/Y OR2X1_LOC_589/A 0.97fF
C38497 OR2X1_LOC_91/Y AND2X1_LOC_471/Y 0.02fF
C38498 OR2X1_LOC_364/A OR2X1_LOC_78/B 0.03fF
C38499 OR2X1_LOC_185/Y OR2X1_LOC_78/B 0.10fF
C38500 AND2X1_LOC_737/Y AND2X1_LOC_811/B 0.00fF
C38501 VDD AND2X1_LOC_211/B 0.94fF
C38502 OR2X1_LOC_485/A AND2X1_LOC_860/A 0.10fF
C38503 VDD OR2X1_LOC_574/A 1.98fF
C38504 OR2X1_LOC_663/A OR2X1_LOC_375/A 0.03fF
C38505 OR2X1_LOC_43/A OR2X1_LOC_59/Y 0.07fF
C38506 OR2X1_LOC_447/Y AND2X1_LOC_7/B 0.32fF
C38507 AND2X1_LOC_40/Y AND2X1_LOC_166/a_8_24# 0.03fF
C38508 VDD OR2X1_LOC_429/Y 0.66fF
C38509 OR2X1_LOC_709/A OR2X1_LOC_19/B 0.04fF
C38510 OR2X1_LOC_318/Y OR2X1_LOC_624/A 0.18fF
C38511 OR2X1_LOC_689/A OR2X1_LOC_39/A 0.02fF
C38512 INPUT_0 OR2X1_LOC_26/Y 0.50fF
C38513 OR2X1_LOC_689/A OR2X1_LOC_459/a_8_216# 0.47fF
C38514 OR2X1_LOC_97/A OR2X1_LOC_443/a_8_216# 0.01fF
C38515 OR2X1_LOC_604/A OR2X1_LOC_481/A 0.24fF
C38516 AND2X1_LOC_857/Y OR2X1_LOC_6/A 0.03fF
C38517 AND2X1_LOC_355/a_8_24# OR2X1_LOC_744/A 0.03fF
C38518 OR2X1_LOC_724/A OR2X1_LOC_317/B 0.02fF
C38519 AND2X1_LOC_366/A OR2X1_LOC_669/Y 0.19fF
C38520 AND2X1_LOC_56/B AND2X1_LOC_39/a_8_24# 0.02fF
C38521 OR2X1_LOC_48/B AND2X1_LOC_435/a_8_24# 0.01fF
C38522 OR2X1_LOC_154/A OR2X1_LOC_61/B 0.33fF
C38523 OR2X1_LOC_137/Y AND2X1_LOC_41/A 0.04fF
C38524 AND2X1_LOC_12/Y OR2X1_LOC_847/A 0.05fF
C38525 AND2X1_LOC_729/Y OR2X1_LOC_427/A 0.03fF
C38526 OR2X1_LOC_814/A OR2X1_LOC_343/a_8_216# 0.01fF
C38527 AND2X1_LOC_773/Y OR2X1_LOC_31/Y 0.16fF
C38528 AND2X1_LOC_70/Y OR2X1_LOC_636/a_8_216# 0.01fF
C38529 OR2X1_LOC_643/Y OR2X1_LOC_641/A 0.03fF
C38530 AND2X1_LOC_191/B OR2X1_LOC_617/Y 0.01fF
C38531 AND2X1_LOC_199/A AND2X1_LOC_196/Y 0.28fF
C38532 AND2X1_LOC_274/a_8_24# OR2X1_LOC_39/A 0.04fF
C38533 OR2X1_LOC_287/B OR2X1_LOC_571/a_8_216# 0.00fF
C38534 OR2X1_LOC_392/A OR2X1_LOC_269/B 0.03fF
C38535 AND2X1_LOC_660/Y OR2X1_LOC_56/A 0.01fF
C38536 AND2X1_LOC_95/Y OR2X1_LOC_668/Y 0.01fF
C38537 OR2X1_LOC_614/a_8_216# OR2X1_LOC_161/B 0.00fF
C38538 OR2X1_LOC_135/Y OR2X1_LOC_111/Y 0.01fF
C38539 OR2X1_LOC_49/A OR2X1_LOC_416/A 0.09fF
C38540 OR2X1_LOC_113/Y AND2X1_LOC_42/B 0.01fF
C38541 OR2X1_LOC_624/A OR2X1_LOC_805/A 3.90fF
C38542 OR2X1_LOC_166/Y OR2X1_LOC_70/Y 0.01fF
C38543 OR2X1_LOC_434/A OR2X1_LOC_390/A 0.55fF
C38544 OR2X1_LOC_128/a_8_216# OR2X1_LOC_161/A 0.14fF
C38545 OR2X1_LOC_18/Y OR2X1_LOC_767/a_8_216# 0.05fF
C38546 OR2X1_LOC_475/Y AND2X1_LOC_92/Y 0.02fF
C38547 AND2X1_LOC_857/Y OR2X1_LOC_299/a_8_216# 0.01fF
C38548 OR2X1_LOC_160/A AND2X1_LOC_59/Y 0.57fF
C38549 OR2X1_LOC_122/Y OR2X1_LOC_3/Y 0.33fF
C38550 OR2X1_LOC_315/Y OR2X1_LOC_39/A 0.03fF
C38551 OR2X1_LOC_719/Y OR2X1_LOC_737/A 0.01fF
C38552 OR2X1_LOC_114/B AND2X1_LOC_127/a_8_24# 0.00fF
C38553 OR2X1_LOC_858/B OR2X1_LOC_850/A 0.03fF
C38554 AND2X1_LOC_514/Y AND2X1_LOC_337/a_8_24# 0.01fF
C38555 OR2X1_LOC_461/Y INPUT_0 0.01fF
C38556 OR2X1_LOC_60/a_8_216# OR2X1_LOC_59/Y 0.02fF
C38557 OR2X1_LOC_689/a_8_216# OR2X1_LOC_690/A 0.01fF
C38558 OR2X1_LOC_60/Y OR2X1_LOC_22/Y 0.01fF
C38559 VDD AND2X1_LOC_672/B 0.16fF
C38560 OR2X1_LOC_160/B OR2X1_LOC_62/B 0.12fF
C38561 AND2X1_LOC_398/a_36_24# OR2X1_LOC_6/A 0.02fF
C38562 AND2X1_LOC_70/Y OR2X1_LOC_19/B 0.04fF
C38563 INPUT_0 AND2X1_LOC_51/Y 0.02fF
C38564 AND2X1_LOC_851/B OR2X1_LOC_522/Y 0.01fF
C38565 AND2X1_LOC_191/Y AND2X1_LOC_866/B 0.01fF
C38566 AND2X1_LOC_658/A AND2X1_LOC_814/a_8_24# 0.06fF
C38567 OR2X1_LOC_696/A AND2X1_LOC_222/Y 0.03fF
C38568 OR2X1_LOC_49/A AND2X1_LOC_8/a_8_24# 0.01fF
C38569 AND2X1_LOC_56/B AND2X1_LOC_43/B 0.12fF
C38570 OR2X1_LOC_604/A OR2X1_LOC_71/Y 0.05fF
C38571 OR2X1_LOC_270/a_8_216# OR2X1_LOC_456/Y 0.01fF
C38572 OR2X1_LOC_185/Y OR2X1_LOC_375/A 0.03fF
C38573 AND2X1_LOC_711/Y AND2X1_LOC_866/B 0.40fF
C38574 OR2X1_LOC_185/A OR2X1_LOC_68/a_8_216# 0.00fF
C38575 AND2X1_LOC_40/Y AND2X1_LOC_183/a_8_24# 0.23fF
C38576 AND2X1_LOC_343/a_8_24# OR2X1_LOC_278/Y 0.00fF
C38577 AND2X1_LOC_228/Y OR2X1_LOC_44/Y 0.01fF
C38578 AND2X1_LOC_544/a_8_24# OR2X1_LOC_70/Y 0.01fF
C38579 OR2X1_LOC_643/A OR2X1_LOC_215/Y 0.18fF
C38580 OR2X1_LOC_329/B AND2X1_LOC_727/A 0.03fF
C38581 AND2X1_LOC_718/a_8_24# OR2X1_LOC_64/Y 0.01fF
C38582 AND2X1_LOC_231/Y AND2X1_LOC_641/a_8_24# 0.11fF
C38583 OR2X1_LOC_54/Y OR2X1_LOC_232/Y 0.03fF
C38584 OR2X1_LOC_70/Y AND2X1_LOC_654/B 0.02fF
C38585 AND2X1_LOC_8/Y AND2X1_LOC_43/B 0.07fF
C38586 OR2X1_LOC_160/B OR2X1_LOC_780/B 0.11fF
C38587 AND2X1_LOC_573/a_8_24# AND2X1_LOC_474/Y 0.00fF
C38588 OR2X1_LOC_8/Y AND2X1_LOC_839/A 0.07fF
C38589 OR2X1_LOC_51/B OR2X1_LOC_36/a_8_216# 0.01fF
C38590 OR2X1_LOC_585/A AND2X1_LOC_403/B 0.05fF
C38591 AND2X1_LOC_487/a_8_24# OR2X1_LOC_287/B 0.00fF
C38592 OR2X1_LOC_70/Y OR2X1_LOC_495/Y 0.03fF
C38593 OR2X1_LOC_474/a_36_216# OR2X1_LOC_624/Y 0.00fF
C38594 OR2X1_LOC_26/Y OR2X1_LOC_11/Y 0.03fF
C38595 OR2X1_LOC_108/Y AND2X1_LOC_866/A 0.07fF
C38596 OR2X1_LOC_678/a_36_216# AND2X1_LOC_48/A 0.00fF
C38597 OR2X1_LOC_219/B OR2X1_LOC_340/Y 0.03fF
C38598 AND2X1_LOC_3/Y AND2X1_LOC_297/a_8_24# 0.01fF
C38599 OR2X1_LOC_509/a_8_216# OR2X1_LOC_227/Y 0.05fF
C38600 VDD OR2X1_LOC_428/a_8_216# 0.21fF
C38601 OR2X1_LOC_190/A AND2X1_LOC_47/Y 0.01fF
C38602 OR2X1_LOC_377/A OR2X1_LOC_654/A 0.07fF
C38603 AND2X1_LOC_717/a_8_24# OR2X1_LOC_371/Y 0.01fF
C38604 AND2X1_LOC_41/A AND2X1_LOC_48/A 0.22fF
C38605 AND2X1_LOC_64/Y OR2X1_LOC_68/B 0.22fF
C38606 OR2X1_LOC_860/Y AND2X1_LOC_51/Y 0.01fF
C38607 AND2X1_LOC_589/a_8_24# OR2X1_LOC_799/A 0.09fF
C38608 OR2X1_LOC_70/Y AND2X1_LOC_450/a_8_24# 0.02fF
C38609 OR2X1_LOC_468/A OR2X1_LOC_436/Y 0.52fF
C38610 OR2X1_LOC_864/A OR2X1_LOC_772/a_8_216# 0.01fF
C38611 OR2X1_LOC_786/Y OR2X1_LOC_641/A 0.03fF
C38612 OR2X1_LOC_503/A OR2X1_LOC_89/A 0.03fF
C38613 OR2X1_LOC_160/A OR2X1_LOC_688/Y 0.10fF
C38614 OR2X1_LOC_696/A OR2X1_LOC_423/Y 0.14fF
C38615 AND2X1_LOC_560/B OR2X1_LOC_26/Y 0.08fF
C38616 OR2X1_LOC_774/Y OR2X1_LOC_772/a_8_216# 0.01fF
C38617 OR2X1_LOC_43/A OR2X1_LOC_820/B 0.02fF
C38618 OR2X1_LOC_246/Y OR2X1_LOC_7/A 0.03fF
C38619 AND2X1_LOC_585/a_8_24# OR2X1_LOC_598/A 0.06fF
C38620 AND2X1_LOC_164/a_8_24# AND2X1_LOC_47/Y 0.01fF
C38621 OR2X1_LOC_585/A OR2X1_LOC_44/Y 0.20fF
C38622 OR2X1_LOC_132/Y AND2X1_LOC_227/Y 0.02fF
C38623 AND2X1_LOC_59/Y OR2X1_LOC_624/B 0.02fF
C38624 AND2X1_LOC_458/Y OR2X1_LOC_371/Y 0.03fF
C38625 VDD OR2X1_LOC_826/Y 0.16fF
C38626 OR2X1_LOC_26/Y OR2X1_LOC_690/A 0.04fF
C38627 AND2X1_LOC_576/Y OR2X1_LOC_7/A 0.07fF
C38628 OR2X1_LOC_329/B OR2X1_LOC_95/Y 0.74fF
C38629 OR2X1_LOC_216/Y AND2X1_LOC_3/Y 0.87fF
C38630 AND2X1_LOC_852/Y OR2X1_LOC_612/B 0.03fF
C38631 OR2X1_LOC_70/Y AND2X1_LOC_365/A 0.01fF
C38632 OR2X1_LOC_151/A AND2X1_LOC_485/a_8_24# 0.12fF
C38633 AND2X1_LOC_456/a_8_24# AND2X1_LOC_657/A 0.02fF
C38634 AND2X1_LOC_72/a_8_24# OR2X1_LOC_631/B 0.04fF
C38635 AND2X1_LOC_560/B OR2X1_LOC_89/A 0.01fF
C38636 AND2X1_LOC_730/a_8_24# AND2X1_LOC_797/A 0.09fF
C38637 OR2X1_LOC_66/A D_INPUT_1 0.10fF
C38638 OR2X1_LOC_743/A OR2X1_LOC_36/Y 0.25fF
C38639 AND2X1_LOC_31/Y OR2X1_LOC_161/B 0.77fF
C38640 OR2X1_LOC_479/Y AND2X1_LOC_369/a_8_24# 0.04fF
C38641 OR2X1_LOC_427/A AND2X1_LOC_639/A 0.04fF
C38642 VDD AND2X1_LOC_781/Y 0.06fF
C38643 AND2X1_LOC_86/Y OR2X1_LOC_62/B 0.01fF
C38644 OR2X1_LOC_748/A OR2X1_LOC_258/Y 0.03fF
C38645 AND2X1_LOC_50/Y AND2X1_LOC_47/Y 1.11fF
C38646 OR2X1_LOC_40/Y AND2X1_LOC_784/a_36_24# 0.00fF
C38647 AND2X1_LOC_514/Y AND2X1_LOC_365/A 0.08fF
C38648 AND2X1_LOC_496/a_36_24# OR2X1_LOC_203/Y 0.00fF
C38649 AND2X1_LOC_82/Y OR2X1_LOC_68/B 0.02fF
C38650 OR2X1_LOC_70/Y OR2X1_LOC_43/A 0.13fF
C38651 INPUT_3 OR2X1_LOC_62/B 0.17fF
C38652 OR2X1_LOC_702/A OR2X1_LOC_155/A 0.14fF
C38653 OR2X1_LOC_662/A AND2X1_LOC_48/A 0.03fF
C38654 OR2X1_LOC_185/A OR2X1_LOC_814/A 0.05fF
C38655 OR2X1_LOC_472/B OR2X1_LOC_375/A 0.39fF
C38656 AND2X1_LOC_598/a_8_24# OR2X1_LOC_64/Y 0.01fF
C38657 OR2X1_LOC_249/Y OR2X1_LOC_814/A 0.00fF
C38658 AND2X1_LOC_17/Y OR2X1_LOC_636/a_8_216# 0.01fF
C38659 OR2X1_LOC_111/Y AND2X1_LOC_520/Y 0.01fF
C38660 OR2X1_LOC_816/Y OR2X1_LOC_815/Y 0.08fF
C38661 AND2X1_LOC_59/Y OR2X1_LOC_655/A 0.00fF
C38662 OR2X1_LOC_777/B OR2X1_LOC_121/A 0.03fF
C38663 OR2X1_LOC_711/A OR2X1_LOC_705/Y 0.74fF
C38664 OR2X1_LOC_64/Y OR2X1_LOC_26/Y 0.36fF
C38665 AND2X1_LOC_11/Y OR2X1_LOC_639/a_8_216# 0.01fF
C38666 OR2X1_LOC_97/B AND2X1_LOC_119/a_8_24# 0.01fF
C38667 OR2X1_LOC_137/B OR2X1_LOC_720/B 0.09fF
C38668 OR2X1_LOC_504/Y AND2X1_LOC_858/a_8_24# 0.24fF
C38669 OR2X1_LOC_580/B OR2X1_LOC_366/Y 0.10fF
C38670 OR2X1_LOC_578/a_8_216# OR2X1_LOC_367/a_8_216# 0.47fF
C38671 OR2X1_LOC_577/Y D_GATE_366 0.02fF
C38672 OR2X1_LOC_62/B OR2X1_LOC_266/a_8_216# 0.01fF
C38673 OR2X1_LOC_36/Y OR2X1_LOC_246/A 0.86fF
C38674 INPUT_5 OR2X1_LOC_51/B 0.02fF
C38675 OR2X1_LOC_416/Y OR2X1_LOC_753/A 0.33fF
C38676 OR2X1_LOC_64/Y AND2X1_LOC_493/a_8_24# 0.05fF
C38677 OR2X1_LOC_462/B OR2X1_LOC_520/A 0.01fF
C38678 OR2X1_LOC_335/B OR2X1_LOC_87/A 0.11fF
C38679 AND2X1_LOC_538/a_8_24# OR2X1_LOC_43/A 0.02fF
C38680 AND2X1_LOC_349/B OR2X1_LOC_64/Y 0.01fF
C38681 OR2X1_LOC_64/Y OR2X1_LOC_89/A 3.67fF
C38682 OR2X1_LOC_599/A AND2X1_LOC_687/Y 0.02fF
C38683 OR2X1_LOC_852/A OR2X1_LOC_375/A 0.01fF
C38684 AND2X1_LOC_113/Y OR2X1_LOC_95/Y 0.01fF
C38685 OR2X1_LOC_432/a_36_216# AND2X1_LOC_648/B 0.00fF
C38686 AND2X1_LOC_841/B OR2X1_LOC_47/Y 0.03fF
C38687 AND2X1_LOC_388/a_36_24# OR2X1_LOC_167/Y 0.01fF
C38688 AND2X1_LOC_86/Y AND2X1_LOC_88/Y 0.07fF
C38689 OR2X1_LOC_647/a_8_216# OR2X1_LOC_647/B 0.04fF
C38690 OR2X1_LOC_625/Y OR2X1_LOC_615/Y 0.03fF
C38691 OR2X1_LOC_45/B OR2X1_LOC_183/a_36_216# 0.03fF
C38692 AND2X1_LOC_808/A AND2X1_LOC_811/B 0.01fF
C38693 OR2X1_LOC_674/Y OR2X1_LOC_39/A 0.00fF
C38694 INPUT_1 AND2X1_LOC_234/a_8_24# 0.02fF
C38695 OR2X1_LOC_78/B OR2X1_LOC_568/A 0.12fF
C38696 AND2X1_LOC_811/a_36_24# AND2X1_LOC_811/Y 0.00fF
C38697 AND2X1_LOC_118/a_8_24# D_INPUT_0 0.03fF
C38698 OR2X1_LOC_26/Y OR2X1_LOC_417/A 2.10fF
C38699 OR2X1_LOC_691/A AND2X1_LOC_36/Y 0.07fF
C38700 OR2X1_LOC_542/B OR2X1_LOC_367/B 2.55fF
C38701 OR2X1_LOC_811/A AND2X1_LOC_72/B 0.03fF
C38702 OR2X1_LOC_121/B OR2X1_LOC_97/a_8_216# 0.50fF
C38703 OR2X1_LOC_416/Y OR2X1_LOC_27/a_36_216# 0.00fF
C38704 AND2X1_LOC_474/A AND2X1_LOC_657/A 0.01fF
C38705 OR2X1_LOC_435/B AND2X1_LOC_31/Y 0.01fF
C38706 OR2X1_LOC_26/Y OR2X1_LOC_64/a_8_216# 0.39fF
C38707 AND2X1_LOC_654/B OR2X1_LOC_70/A 0.00fF
C38708 AND2X1_LOC_645/a_8_24# OR2X1_LOC_44/Y 0.02fF
C38709 OR2X1_LOC_76/A OR2X1_LOC_121/B 0.00fF
C38710 OR2X1_LOC_89/A OR2X1_LOC_417/A 0.30fF
C38711 OR2X1_LOC_841/a_8_216# OR2X1_LOC_228/Y 0.02fF
C38712 OR2X1_LOC_831/B OR2X1_LOC_121/A 0.00fF
C38713 OR2X1_LOC_435/Y OR2X1_LOC_814/A 0.01fF
C38714 OR2X1_LOC_405/A OR2X1_LOC_374/Y 0.00fF
C38715 OR2X1_LOC_115/a_36_216# OR2X1_LOC_66/Y 0.00fF
C38716 AND2X1_LOC_624/B OR2X1_LOC_39/A 0.00fF
C38717 OR2X1_LOC_39/A OR2X1_LOC_67/Y 0.03fF
C38718 AND2X1_LOC_390/B AND2X1_LOC_801/B 0.02fF
C38719 OR2X1_LOC_188/a_8_216# OR2X1_LOC_121/A 0.41fF
C38720 OR2X1_LOC_114/Y OR2X1_LOC_786/Y 0.00fF
C38721 OR2X1_LOC_182/B OR2X1_LOC_212/B 0.44fF
C38722 AND2X1_LOC_350/B OR2X1_LOC_171/Y 0.77fF
C38723 AND2X1_LOC_531/a_8_24# OR2X1_LOC_348/B 0.23fF
C38724 OR2X1_LOC_47/Y OR2X1_LOC_22/a_8_216# 0.39fF
C38725 OR2X1_LOC_415/Y AND2X1_LOC_44/Y 0.00fF
C38726 AND2X1_LOC_580/A AND2X1_LOC_792/Y 0.07fF
C38727 OR2X1_LOC_61/Y AND2X1_LOC_31/Y 0.02fF
C38728 OR2X1_LOC_856/B OR2X1_LOC_228/Y 0.07fF
C38729 OR2X1_LOC_217/Y OR2X1_LOC_66/a_8_216# 0.40fF
C38730 OR2X1_LOC_632/Y OR2X1_LOC_501/a_8_216# 0.02fF
C38731 OR2X1_LOC_40/Y AND2X1_LOC_793/a_8_24# 0.01fF
C38732 AND2X1_LOC_848/A AND2X1_LOC_848/Y 0.07fF
C38733 OR2X1_LOC_810/a_8_216# OR2X1_LOC_561/B 0.02fF
C38734 OR2X1_LOC_555/B OR2X1_LOC_259/B 0.17fF
C38735 OR2X1_LOC_66/A OR2X1_LOC_180/B 0.01fF
C38736 OR2X1_LOC_65/B OR2X1_LOC_88/a_8_216# 0.01fF
C38737 OR2X1_LOC_612/B AND2X1_LOC_647/B 0.03fF
C38738 AND2X1_LOC_810/A AND2X1_LOC_802/B 0.01fF
C38739 OR2X1_LOC_375/A OR2X1_LOC_552/A 0.48fF
C38740 AND2X1_LOC_456/B OR2X1_LOC_13/B 0.02fF
C38741 AND2X1_LOC_379/a_8_24# OR2X1_LOC_70/A 0.01fF
C38742 OR2X1_LOC_185/A OR2X1_LOC_341/a_8_216# 0.01fF
C38743 OR2X1_LOC_45/B AND2X1_LOC_340/Y 0.04fF
C38744 AND2X1_LOC_227/Y AND2X1_LOC_849/A 0.01fF
C38745 OR2X1_LOC_244/A OR2X1_LOC_62/B 0.05fF
C38746 OR2X1_LOC_709/B AND2X1_LOC_7/B 0.11fF
C38747 AND2X1_LOC_23/a_8_24# OR2X1_LOC_532/B 0.01fF
C38748 AND2X1_LOC_431/a_8_24# OR2X1_LOC_814/A 0.01fF
C38749 AND2X1_LOC_3/Y AND2X1_LOC_418/a_36_24# 0.00fF
C38750 AND2X1_LOC_798/a_8_24# AND2X1_LOC_436/Y 0.03fF
C38751 OR2X1_LOC_375/A OR2X1_LOC_578/B 0.03fF
C38752 OR2X1_LOC_678/Y AND2X1_LOC_36/Y 0.00fF
C38753 OR2X1_LOC_45/B AND2X1_LOC_181/Y 0.03fF
C38754 OR2X1_LOC_848/A OR2X1_LOC_561/B 0.40fF
C38755 AND2X1_LOC_787/A AND2X1_LOC_182/A 0.01fF
C38756 AND2X1_LOC_831/Y D_INPUT_0 0.17fF
C38757 OR2X1_LOC_167/a_36_216# OR2X1_LOC_16/A 0.00fF
C38758 OR2X1_LOC_12/Y OR2X1_LOC_604/Y 0.01fF
C38759 OR2X1_LOC_205/a_8_216# OR2X1_LOC_560/A 0.00fF
C38760 VDD OR2X1_LOC_773/Y 0.00fF
C38761 OR2X1_LOC_859/B OR2X1_LOC_561/B 0.04fF
C38762 OR2X1_LOC_22/Y AND2X1_LOC_660/A 0.07fF
C38763 OR2X1_LOC_43/A OR2X1_LOC_534/a_36_216# 0.03fF
C38764 AND2X1_LOC_564/A VDD 0.56fF
C38765 AND2X1_LOC_672/a_8_24# INPUT_1 0.03fF
C38766 VDD OR2X1_LOC_855/A 0.21fF
C38767 OR2X1_LOC_348/Y OR2X1_LOC_366/B 0.27fF
C38768 OR2X1_LOC_696/A AND2X1_LOC_367/A 0.14fF
C38769 AND2X1_LOC_48/A OR2X1_LOC_207/a_8_216# 0.01fF
C38770 OR2X1_LOC_502/A INPUT_6 0.02fF
C38771 OR2X1_LOC_753/A OR2X1_LOC_80/A 0.10fF
C38772 AND2X1_LOC_70/Y OR2X1_LOC_828/Y 0.13fF
C38773 AND2X1_LOC_575/a_8_24# AND2X1_LOC_570/Y 0.01fF
C38774 OR2X1_LOC_32/Y OR2X1_LOC_68/B 0.02fF
C38775 AND2X1_LOC_56/B OR2X1_LOC_367/B 0.05fF
C38776 OR2X1_LOC_485/A AND2X1_LOC_562/Y 0.04fF
C38777 AND2X1_LOC_564/A AND2X1_LOC_738/a_8_24# 0.03fF
C38778 OR2X1_LOC_731/a_8_216# OR2X1_LOC_731/B 0.39fF
C38779 OR2X1_LOC_40/Y OR2X1_LOC_16/A 0.65fF
C38780 AND2X1_LOC_12/Y OR2X1_LOC_544/B 0.07fF
C38781 OR2X1_LOC_811/A AND2X1_LOC_36/Y 0.03fF
C38782 VDD OR2X1_LOC_744/Y 0.06fF
C38783 AND2X1_LOC_251/a_8_24# OR2X1_LOC_580/A 0.24fF
C38784 OR2X1_LOC_600/A AND2X1_LOC_786/Y 0.07fF
C38785 OR2X1_LOC_36/Y OR2X1_LOC_599/a_8_216# 0.09fF
C38786 VDD AND2X1_LOC_727/B 0.31fF
C38787 OR2X1_LOC_6/A OR2X1_LOC_437/A 0.07fF
C38788 AND2X1_LOC_182/A AND2X1_LOC_566/B 0.53fF
C38789 AND2X1_LOC_59/a_8_24# AND2X1_LOC_36/Y 0.01fF
C38790 AND2X1_LOC_59/Y OR2X1_LOC_532/Y 0.18fF
C38791 GATE_662 OR2X1_LOC_95/Y 0.05fF
C38792 AND2X1_LOC_61/a_8_24# OR2X1_LOC_12/Y 0.00fF
C38793 OR2X1_LOC_335/A OR2X1_LOC_808/B 0.03fF
C38794 OR2X1_LOC_575/A OR2X1_LOC_501/A 0.19fF
C38795 AND2X1_LOC_357/A OR2X1_LOC_158/A 0.03fF
C38796 OR2X1_LOC_709/A AND2X1_LOC_313/a_36_24# 0.01fF
C38797 AND2X1_LOC_562/a_8_24# OR2X1_LOC_698/Y 0.23fF
C38798 OR2X1_LOC_49/A AND2X1_LOC_19/Y 0.10fF
C38799 OR2X1_LOC_56/A AND2X1_LOC_795/a_8_24# 0.01fF
C38800 AND2X1_LOC_240/Y OR2X1_LOC_71/A 0.02fF
C38801 OR2X1_LOC_632/Y AND2X1_LOC_44/Y 0.15fF
C38802 D_INPUT_0 OR2X1_LOC_339/Y 0.05fF
C38803 OR2X1_LOC_744/A OR2X1_LOC_12/Y 1.51fF
C38804 OR2X1_LOC_40/Y OR2X1_LOC_108/Y 0.03fF
C38805 AND2X1_LOC_512/a_8_24# OR2X1_LOC_13/B 0.01fF
C38806 AND2X1_LOC_462/B AND2X1_LOC_293/a_8_24# 0.08fF
C38807 AND2X1_LOC_47/Y OR2X1_LOC_241/B 0.17fF
C38808 OR2X1_LOC_158/A AND2X1_LOC_367/B 0.04fF
C38809 OR2X1_LOC_207/B AND2X1_LOC_41/A 0.39fF
C38810 AND2X1_LOC_92/Y OR2X1_LOC_356/A 0.07fF
C38811 OR2X1_LOC_206/A OR2X1_LOC_68/B 0.05fF
C38812 AND2X1_LOC_465/a_8_24# OR2X1_LOC_437/A 0.01fF
C38813 OR2X1_LOC_92/Y OR2X1_LOC_312/a_8_216# 0.13fF
C38814 OR2X1_LOC_51/Y OR2X1_LOC_583/a_8_216# 0.01fF
C38815 AND2X1_LOC_584/a_36_24# OR2X1_LOC_639/B 0.01fF
C38816 AND2X1_LOC_388/Y OR2X1_LOC_166/a_36_216# 0.00fF
C38817 VDD OR2X1_LOC_536/Y 0.16fF
C38818 OR2X1_LOC_106/Y AND2X1_LOC_99/A 0.03fF
C38819 AND2X1_LOC_547/Y AND2X1_LOC_550/a_36_24# 0.01fF
C38820 AND2X1_LOC_262/a_8_24# OR2X1_LOC_78/A 0.01fF
C38821 OR2X1_LOC_604/A OR2X1_LOC_426/B 0.00fF
C38822 AND2X1_LOC_70/Y AND2X1_LOC_110/Y 0.04fF
C38823 OR2X1_LOC_860/a_36_216# OR2X1_LOC_392/B 0.15fF
C38824 OR2X1_LOC_528/Y AND2X1_LOC_663/A 0.45fF
C38825 OR2X1_LOC_125/a_8_216# OR2X1_LOC_51/Y 0.01fF
C38826 OR2X1_LOC_405/A OR2X1_LOC_392/B 0.10fF
C38827 INPUT_0 AND2X1_LOC_194/Y 0.90fF
C38828 OR2X1_LOC_663/A OR2X1_LOC_549/A 0.07fF
C38829 AND2X1_LOC_658/a_8_24# AND2X1_LOC_658/Y 0.01fF
C38830 AND2X1_LOC_358/Y AND2X1_LOC_364/A 0.02fF
C38831 AND2X1_LOC_843/Y AND2X1_LOC_244/A 0.00fF
C38832 OR2X1_LOC_529/Y OR2X1_LOC_183/a_8_216# 0.01fF
C38833 OR2X1_LOC_359/a_8_216# OR2X1_LOC_359/A 0.39fF
C38834 OR2X1_LOC_759/A OR2X1_LOC_816/Y 0.02fF
C38835 OR2X1_LOC_161/A AND2X1_LOC_7/B 0.29fF
C38836 AND2X1_LOC_361/a_8_24# OR2X1_LOC_103/Y 0.01fF
C38837 OR2X1_LOC_21/a_8_216# AND2X1_LOC_409/B 0.47fF
C38838 D_INPUT_4 OR2X1_LOC_596/A 0.01fF
C38839 OR2X1_LOC_703/A AND2X1_LOC_110/Y 0.01fF
C38840 OR2X1_LOC_174/A AND2X1_LOC_18/Y 0.11fF
C38841 VDD AND2X1_LOC_474/A 0.48fF
C38842 OR2X1_LOC_696/A AND2X1_LOC_673/a_8_24# 0.01fF
C38843 VDD OR2X1_LOC_421/a_8_216# 0.00fF
C38844 AND2X1_LOC_59/Y OR2X1_LOC_266/A 0.16fF
C38845 OR2X1_LOC_56/A AND2X1_LOC_434/Y 0.14fF
C38846 OR2X1_LOC_380/a_36_216# OR2X1_LOC_25/Y 0.02fF
C38847 AND2X1_LOC_22/Y OR2X1_LOC_668/Y 0.05fF
C38848 OR2X1_LOC_680/A GATE_579 0.03fF
C38849 OR2X1_LOC_160/B OR2X1_LOC_659/A 0.02fF
C38850 OR2X1_LOC_696/A AND2X1_LOC_456/Y 0.02fF
C38851 OR2X1_LOC_158/A AND2X1_LOC_852/B 0.02fF
C38852 AND2X1_LOC_644/Y OR2X1_LOC_16/A 0.01fF
C38853 OR2X1_LOC_78/A AND2X1_LOC_437/a_8_24# 0.04fF
C38854 AND2X1_LOC_396/a_8_24# OR2X1_LOC_78/Y 0.01fF
C38855 OR2X1_LOC_45/B AND2X1_LOC_228/Y 0.28fF
C38856 OR2X1_LOC_87/A OR2X1_LOC_267/Y 0.03fF
C38857 OR2X1_LOC_190/B OR2X1_LOC_190/a_8_216# 0.01fF
C38858 AND2X1_LOC_706/Y OR2X1_LOC_432/Y 0.40fF
C38859 OR2X1_LOC_154/A OR2X1_LOC_97/A 0.03fF
C38860 AND2X1_LOC_360/a_8_24# AND2X1_LOC_860/A 0.06fF
C38861 OR2X1_LOC_696/A OR2X1_LOC_74/A 0.76fF
C38862 AND2X1_LOC_176/a_36_24# OR2X1_LOC_180/B 0.00fF
C38863 AND2X1_LOC_580/A OR2X1_LOC_816/A 0.06fF
C38864 OR2X1_LOC_158/A OR2X1_LOC_48/B 0.25fF
C38865 OR2X1_LOC_220/B OR2X1_LOC_550/a_8_216# 0.01fF
C38866 AND2X1_LOC_541/a_8_24# OR2X1_LOC_26/Y 0.01fF
C38867 OR2X1_LOC_368/Y OR2X1_LOC_44/Y 0.04fF
C38868 AND2X1_LOC_486/Y OR2X1_LOC_485/Y 0.00fF
C38869 OR2X1_LOC_338/a_36_216# AND2X1_LOC_95/Y 0.00fF
C38870 OR2X1_LOC_122/a_8_216# AND2X1_LOC_367/A 0.28fF
C38871 OR2X1_LOC_158/A OR2X1_LOC_18/Y 2.18fF
C38872 OR2X1_LOC_326/B OR2X1_LOC_325/B 0.01fF
C38873 AND2X1_LOC_658/B AND2X1_LOC_866/B 0.45fF
C38874 OR2X1_LOC_189/Y AND2X1_LOC_192/a_8_24# 0.09fF
C38875 AND2X1_LOC_168/Y OR2X1_LOC_40/Y 0.14fF
C38876 OR2X1_LOC_19/B OR2X1_LOC_395/a_8_216# 0.03fF
C38877 OR2X1_LOC_24/a_8_216# AND2X1_LOC_208/Y 0.02fF
C38878 AND2X1_LOC_365/a_36_24# OR2X1_LOC_91/A 0.00fF
C38879 AND2X1_LOC_482/a_8_24# AND2X1_LOC_18/Y 0.01fF
C38880 VDD OR2X1_LOC_818/Y 0.12fF
C38881 AND2X1_LOC_597/a_8_24# OR2X1_LOC_161/B 0.01fF
C38882 AND2X1_LOC_557/Y OR2X1_LOC_595/A 0.05fF
C38883 OR2X1_LOC_502/A OR2X1_LOC_648/A 0.08fF
C38884 OR2X1_LOC_229/a_8_216# OR2X1_LOC_44/Y -0.00fF
C38885 OR2X1_LOC_798/Y OR2X1_LOC_78/B 0.05fF
C38886 OR2X1_LOC_179/Y OR2X1_LOC_329/B 0.01fF
C38887 OR2X1_LOC_154/A D_GATE_662 0.01fF
C38888 VDD AND2X1_LOC_16/a_8_24# 0.00fF
C38889 OR2X1_LOC_45/B OR2X1_LOC_585/A 0.19fF
C38890 OR2X1_LOC_864/A OR2X1_LOC_161/B 0.03fF
C38891 AND2X1_LOC_722/Y AND2X1_LOC_722/A 0.04fF
C38892 OR2X1_LOC_160/B AND2X1_LOC_487/a_8_24# 0.04fF
C38893 OR2X1_LOC_185/Y OR2X1_LOC_549/A 0.10fF
C38894 OR2X1_LOC_415/a_36_216# OR2X1_LOC_395/Y 0.00fF
C38895 OR2X1_LOC_7/A AND2X1_LOC_244/A 0.03fF
C38896 AND2X1_LOC_95/Y OR2X1_LOC_66/A 13.47fF
C38897 AND2X1_LOC_3/Y OR2X1_LOC_576/A 0.03fF
C38898 VDD AND2X1_LOC_593/Y 0.08fF
C38899 VDD OR2X1_LOC_377/A 2.16fF
C38900 OR2X1_LOC_856/A OR2X1_LOC_269/B 0.02fF
C38901 OR2X1_LOC_633/Y OR2X1_LOC_66/A 0.03fF
C38902 OR2X1_LOC_8/Y OR2X1_LOC_63/a_8_216# 0.07fF
C38903 OR2X1_LOC_302/B OR2X1_LOC_620/Y 0.01fF
C38904 OR2X1_LOC_60/Y OR2X1_LOC_39/A 0.02fF
C38905 OR2X1_LOC_7/A OR2X1_LOC_16/A 14.31fF
C38906 AND2X1_LOC_658/B AND2X1_LOC_622/a_8_24# 0.01fF
C38907 AND2X1_LOC_358/Y OR2X1_LOC_3/Y 0.03fF
C38908 OR2X1_LOC_204/Y OR2X1_LOC_641/A 0.39fF
C38909 OR2X1_LOC_246/Y OR2X1_LOC_822/a_8_216# 0.40fF
C38910 VDD AND2X1_LOC_824/B 0.51fF
C38911 OR2X1_LOC_102/a_8_216# OR2X1_LOC_585/A 0.01fF
C38912 OR2X1_LOC_249/Y OR2X1_LOC_244/Y 0.00fF
C38913 OR2X1_LOC_617/Y AND2X1_LOC_580/a_36_24# 0.00fF
C38914 OR2X1_LOC_526/Y OR2X1_LOC_511/Y 0.03fF
C38915 OR2X1_LOC_185/A OR2X1_LOC_192/A 0.02fF
C38916 OR2X1_LOC_744/A OR2X1_LOC_393/Y 0.09fF
C38917 OR2X1_LOC_49/A AND2X1_LOC_345/Y 0.07fF
C38918 AND2X1_LOC_570/Y AND2X1_LOC_624/A 0.03fF
C38919 AND2X1_LOC_51/Y AND2X1_LOC_7/B 0.34fF
C38920 OR2X1_LOC_436/Y OR2X1_LOC_175/a_36_216# 0.00fF
C38921 OR2X1_LOC_851/a_36_216# AND2X1_LOC_43/B 0.02fF
C38922 AND2X1_LOC_164/a_8_24# OR2X1_LOC_506/A 0.00fF
C38923 OR2X1_LOC_329/a_36_216# OR2X1_LOC_585/A 0.00fF
C38924 VDD OR2X1_LOC_85/A 0.82fF
C38925 OR2X1_LOC_690/A AND2X1_LOC_194/Y 0.03fF
C38926 AND2X1_LOC_43/B AND2X1_LOC_92/Y 0.13fF
C38927 OR2X1_LOC_306/a_8_216# INPUT_0 0.01fF
C38928 OR2X1_LOC_372/a_8_216# AND2X1_LOC_786/Y 0.06fF
C38929 AND2X1_LOC_312/a_8_24# OR2X1_LOC_220/B 0.01fF
C38930 OR2X1_LOC_329/a_8_216# OR2X1_LOC_485/A 0.02fF
C38931 AND2X1_LOC_715/A OR2X1_LOC_6/A 1.33fF
C38932 OR2X1_LOC_759/A OR2X1_LOC_748/A 0.59fF
C38933 OR2X1_LOC_309/a_36_216# AND2X1_LOC_211/B 0.01fF
C38934 OR2X1_LOC_160/B OR2X1_LOC_449/B 5.09fF
C38935 AND2X1_LOC_12/Y OR2X1_LOC_561/Y 0.01fF
C38936 OR2X1_LOC_145/a_36_216# AND2X1_LOC_658/A 0.02fF
C38937 AND2X1_LOC_522/a_36_24# OR2X1_LOC_404/Y 0.00fF
C38938 AND2X1_LOC_860/a_36_24# OR2X1_LOC_18/Y 0.02fF
C38939 AND2X1_LOC_12/Y OR2X1_LOC_78/Y 0.00fF
C38940 OR2X1_LOC_624/Y OR2X1_LOC_659/a_8_216# 0.40fF
C38941 OR2X1_LOC_143/a_8_216# D_INPUT_3 0.01fF
C38942 OR2X1_LOC_99/Y OR2X1_LOC_66/A 0.39fF
C38943 AND2X1_LOC_140/a_36_24# OR2X1_LOC_595/A 0.00fF
C38944 AND2X1_LOC_72/B OR2X1_LOC_777/B 0.03fF
C38945 AND2X1_LOC_774/a_8_24# AND2X1_LOC_307/Y 0.01fF
C38946 OR2X1_LOC_264/a_8_216# OR2X1_LOC_78/A 0.01fF
C38947 OR2X1_LOC_317/a_36_216# OR2X1_LOC_739/A 0.00fF
C38948 OR2X1_LOC_108/Y OR2X1_LOC_7/A 0.50fF
C38949 AND2X1_LOC_19/Y OR2X1_LOC_87/B 0.05fF
C38950 OR2X1_LOC_467/A OR2X1_LOC_449/A 0.00fF
C38951 OR2X1_LOC_502/A OR2X1_LOC_405/a_8_216# 0.03fF
C38952 OR2X1_LOC_656/B OR2X1_LOC_264/Y 0.08fF
C38953 OR2X1_LOC_167/a_8_216# OR2X1_LOC_64/Y 0.08fF
C38954 OR2X1_LOC_154/A OR2X1_LOC_541/A 0.05fF
C38955 OR2X1_LOC_3/B D_INPUT_6 0.01fF
C38956 OR2X1_LOC_319/B OR2X1_LOC_161/A 0.12fF
C38957 OR2X1_LOC_305/a_8_216# OR2X1_LOC_91/A 0.06fF
C38958 OR2X1_LOC_496/Y OR2X1_LOC_56/A 0.00fF
C38959 OR2X1_LOC_604/A OR2X1_LOC_743/A 0.61fF
C38960 AND2X1_LOC_40/Y OR2X1_LOC_806/a_8_216# 0.01fF
C38961 AND2X1_LOC_41/A OR2X1_LOC_790/a_8_216# 0.02fF
C38962 OR2X1_LOC_45/B AND2X1_LOC_634/Y 0.04fF
C38963 OR2X1_LOC_377/A OR2X1_LOC_689/A 0.03fF
C38964 OR2X1_LOC_325/A AND2X1_LOC_59/Y 0.00fF
C38965 OR2X1_LOC_185/A OR2X1_LOC_147/B 0.06fF
C38966 AND2X1_LOC_367/A OR2X1_LOC_271/B 0.02fF
C38967 OR2X1_LOC_857/a_8_216# OR2X1_LOC_863/A 0.01fF
C38968 OR2X1_LOC_756/B OR2X1_LOC_465/a_8_216# 0.14fF
C38969 OR2X1_LOC_631/B OR2X1_LOC_632/a_8_216# 0.01fF
C38970 OR2X1_LOC_160/A OR2X1_LOC_623/B 0.10fF
C38971 AND2X1_LOC_339/B AND2X1_LOC_351/Y 0.19fF
C38972 AND2X1_LOC_52/a_8_24# OR2X1_LOC_375/A 0.02fF
C38973 OR2X1_LOC_756/B AND2X1_LOC_251/a_36_24# 0.00fF
C38974 OR2X1_LOC_318/Y OR2X1_LOC_161/A 0.01fF
C38975 OR2X1_LOC_479/Y OR2X1_LOC_776/Y 0.12fF
C38976 AND2X1_LOC_578/A OR2X1_LOC_600/A 0.03fF
C38977 AND2X1_LOC_486/Y OR2X1_LOC_39/A 0.64fF
C38978 OR2X1_LOC_352/A OR2X1_LOC_87/A 0.04fF
C38979 D_INPUT_5 AND2X1_LOC_459/Y 0.01fF
C38980 OR2X1_LOC_185/A AND2X1_LOC_517/a_8_24# 0.02fF
C38981 AND2X1_LOC_367/A AND2X1_LOC_359/a_8_24# 0.01fF
C38982 AND2X1_LOC_53/a_8_24# OR2X1_LOC_375/A 0.01fF
C38983 AND2X1_LOC_347/Y OR2X1_LOC_44/Y 2.88fF
C38984 OR2X1_LOC_68/B OR2X1_LOC_558/a_36_216# 0.00fF
C38985 AND2X1_LOC_857/Y OR2X1_LOC_44/Y 0.06fF
C38986 OR2X1_LOC_698/Y OR2X1_LOC_748/A 0.09fF
C38987 OR2X1_LOC_654/A OR2X1_LOC_78/B 0.01fF
C38988 AND2X1_LOC_191/a_8_24# AND2X1_LOC_866/A 0.03fF
C38989 AND2X1_LOC_543/Y OR2X1_LOC_47/Y 0.15fF
C38990 AND2X1_LOC_476/A AND2X1_LOC_473/Y 0.01fF
C38991 OR2X1_LOC_768/A OR2X1_LOC_557/A 0.00fF
C38992 OR2X1_LOC_299/Y OR2X1_LOC_59/Y 0.07fF
C38993 AND2X1_LOC_404/A AND2X1_LOC_404/a_8_24# 0.18fF
C38994 AND2X1_LOC_348/A AND2X1_LOC_359/B 0.01fF
C38995 OR2X1_LOC_105/a_8_216# OR2X1_LOC_810/A 0.17fF
C38996 OR2X1_LOC_770/B OR2X1_LOC_770/a_8_216# 0.00fF
C38997 AND2X1_LOC_41/A AND2X1_LOC_3/Y 2.06fF
C38998 OR2X1_LOC_612/B AND2X1_LOC_647/a_36_24# 0.00fF
C38999 OR2X1_LOC_160/B OR2X1_LOC_121/B 0.10fF
C39000 AND2X1_LOC_721/Y OR2X1_LOC_224/Y 0.04fF
C39001 OR2X1_LOC_31/Y OR2X1_LOC_12/Y 1.38fF
C39002 AND2X1_LOC_64/Y OR2X1_LOC_247/a_8_216# 0.01fF
C39003 OR2X1_LOC_3/Y OR2X1_LOC_820/A 0.02fF
C39004 AND2X1_LOC_40/Y OR2X1_LOC_389/B 0.06fF
C39005 OR2X1_LOC_96/Y OR2X1_LOC_54/Y 0.09fF
C39006 OR2X1_LOC_805/A OR2X1_LOC_161/A 0.10fF
C39007 OR2X1_LOC_40/Y AND2X1_LOC_128/a_8_24# 0.01fF
C39008 OR2X1_LOC_31/Y OR2X1_LOC_766/Y 0.21fF
C39009 AND2X1_LOC_148/a_36_24# OR2X1_LOC_74/A 0.01fF
C39010 AND2X1_LOC_40/Y AND2X1_LOC_118/a_8_24# 0.07fF
C39011 OR2X1_LOC_178/Y AND2X1_LOC_523/Y 0.03fF
C39012 OR2X1_LOC_676/Y OR2X1_LOC_196/B 0.08fF
C39013 AND2X1_LOC_540/a_8_24# OR2X1_LOC_529/Y 0.01fF
C39014 OR2X1_LOC_541/A OR2X1_LOC_778/A 0.61fF
C39015 OR2X1_LOC_756/B OR2X1_LOC_479/Y 0.03fF
C39016 OR2X1_LOC_499/B AND2X1_LOC_42/B 0.06fF
C39017 OR2X1_LOC_427/A AND2X1_LOC_374/Y 0.03fF
C39018 OR2X1_LOC_366/Y OR2X1_LOC_367/a_8_216# 0.01fF
C39019 OR2X1_LOC_508/A AND2X1_LOC_3/Y 0.46fF
C39020 AND2X1_LOC_777/a_8_24# OR2X1_LOC_619/Y 0.02fF
C39021 OR2X1_LOC_6/B D_INPUT_0 2.28fF
C39022 AND2X1_LOC_93/a_8_24# AND2X1_LOC_47/Y 0.03fF
C39023 AND2X1_LOC_12/Y OR2X1_LOC_285/A 0.01fF
C39024 OR2X1_LOC_656/B OR2X1_LOC_643/A 0.07fF
C39025 D_INPUT_4 OR2X1_LOC_21/a_36_216# 0.03fF
C39026 AND2X1_LOC_334/Y OR2X1_LOC_46/A 0.02fF
C39027 AND2X1_LOC_580/A AND2X1_LOC_807/Y 1.46fF
C39028 OR2X1_LOC_427/A OR2X1_LOC_52/B 0.27fF
C39029 AND2X1_LOC_276/Y AND2X1_LOC_276/a_8_24# 0.01fF
C39030 OR2X1_LOC_655/a_8_216# AND2X1_LOC_8/Y 0.01fF
C39031 AND2X1_LOC_550/A OR2X1_LOC_26/Y 0.01fF
C39032 OR2X1_LOC_599/A AND2X1_LOC_676/a_36_24# 0.01fF
C39033 OR2X1_LOC_149/B OR2X1_LOC_705/B 0.01fF
C39034 OR2X1_LOC_648/A AND2X1_LOC_48/A 0.08fF
C39035 OR2X1_LOC_47/Y AND2X1_LOC_770/a_8_24# 0.01fF
C39036 OR2X1_LOC_377/A OR2X1_LOC_836/B 0.03fF
C39037 OR2X1_LOC_247/Y OR2X1_LOC_563/A 0.02fF
C39038 OR2X1_LOC_389/B OR2X1_LOC_537/A 0.16fF
C39039 AND2X1_LOC_489/Y OR2X1_LOC_427/A 0.03fF
C39040 OR2X1_LOC_325/B AND2X1_LOC_47/Y 0.09fF
C39041 OR2X1_LOC_520/Y OR2X1_LOC_87/A 0.03fF
C39042 AND2X1_LOC_7/B OR2X1_LOC_551/B 0.07fF
C39043 OR2X1_LOC_319/B AND2X1_LOC_51/Y 0.01fF
C39044 VDD OR2X1_LOC_226/Y 0.04fF
C39045 OR2X1_LOC_774/Y OR2X1_LOC_846/a_8_216# 0.02fF
C39046 OR2X1_LOC_85/A AND2X1_LOC_267/a_8_24# 0.17fF
C39047 OR2X1_LOC_589/A OR2X1_LOC_47/Y 0.32fF
C39048 AND2X1_LOC_63/a_8_24# OR2X1_LOC_267/A 0.01fF
C39049 AND2X1_LOC_91/B OR2X1_LOC_398/Y 0.49fF
C39050 AND2X1_LOC_326/B AND2X1_LOC_831/Y 0.00fF
C39051 OR2X1_LOC_318/A OR2X1_LOC_804/A 0.10fF
C39052 OR2X1_LOC_321/Y AND2X1_LOC_654/Y 0.04fF
C39053 OR2X1_LOC_108/Y OR2X1_LOC_224/a_8_216# 0.02fF
C39054 AND2X1_LOC_141/a_8_24# OR2X1_LOC_71/Y 0.01fF
C39055 OR2X1_LOC_47/Y OR2X1_LOC_322/Y 0.15fF
C39056 OR2X1_LOC_485/A AND2X1_LOC_287/a_8_24# 0.06fF
C39057 OR2X1_LOC_669/A OR2X1_LOC_669/a_8_216# 0.47fF
C39058 OR2X1_LOC_497/Y OR2X1_LOC_36/Y 0.07fF
C39059 INPUT_0 OR2X1_LOC_243/a_8_216# 0.01fF
C39060 AND2X1_LOC_485/a_36_24# AND2X1_LOC_44/Y 0.00fF
C39061 OR2X1_LOC_753/A OR2X1_LOC_6/A 0.10fF
C39062 OR2X1_LOC_296/Y OR2X1_LOC_161/A 0.02fF
C39063 OR2X1_LOC_654/A OR2X1_LOC_375/A 0.00fF
C39064 AND2X1_LOC_36/Y OR2X1_LOC_777/B 0.05fF
C39065 AND2X1_LOC_140/a_8_24# OR2X1_LOC_118/Y 0.01fF
C39066 OR2X1_LOC_306/Y OR2X1_LOC_743/A 0.01fF
C39067 AND2X1_LOC_716/a_8_24# AND2X1_LOC_211/B 0.01fF
C39068 AND2X1_LOC_301/a_36_24# AND2X1_LOC_476/A 0.01fF
C39069 AND2X1_LOC_101/B OR2X1_LOC_26/Y 0.03fF
C39070 AND2X1_LOC_191/Y OR2X1_LOC_613/a_36_216# 0.02fF
C39071 OR2X1_LOC_485/A OR2X1_LOC_235/a_8_216# 0.03fF
C39072 OR2X1_LOC_11/Y OR2X1_LOC_17/Y 0.13fF
C39073 AND2X1_LOC_851/B OR2X1_LOC_56/A 0.09fF
C39074 OR2X1_LOC_190/A OR2X1_LOC_284/B 0.00fF
C39075 OR2X1_LOC_673/Y AND2X1_LOC_85/a_8_24# 0.02fF
C39076 OR2X1_LOC_158/A AND2X1_LOC_215/A 0.03fF
C39077 OR2X1_LOC_91/A AND2X1_LOC_137/a_8_24# 0.03fF
C39078 OR2X1_LOC_507/A OR2X1_LOC_205/Y 0.06fF
C39079 OR2X1_LOC_631/B AND2X1_LOC_3/Y 0.06fF
C39080 OR2X1_LOC_407/a_8_216# AND2X1_LOC_51/Y 0.14fF
C39081 AND2X1_LOC_649/B OR2X1_LOC_46/A 0.03fF
C39082 OR2X1_LOC_805/A AND2X1_LOC_51/Y 0.07fF
C39083 OR2X1_LOC_686/A OR2X1_LOC_451/B 0.02fF
C39084 OR2X1_LOC_166/Y OR2X1_LOC_47/Y 0.03fF
C39085 OR2X1_LOC_406/A AND2X1_LOC_778/Y 0.23fF
C39086 AND2X1_LOC_47/Y AND2X1_LOC_615/a_8_24# 0.01fF
C39087 OR2X1_LOC_653/Y OR2X1_LOC_655/B 0.01fF
C39088 AND2X1_LOC_6/a_36_24# OR2X1_LOC_78/A 0.01fF
C39089 OR2X1_LOC_485/A OR2X1_LOC_239/Y 0.04fF
C39090 AND2X1_LOC_259/Y AND2X1_LOC_345/Y 0.13fF
C39091 OR2X1_LOC_857/a_8_216# AND2X1_LOC_56/B 0.03fF
C39092 OR2X1_LOC_831/a_36_216# OR2X1_LOC_121/B 0.00fF
C39093 OR2X1_LOC_578/B OR2X1_LOC_549/A 0.13fF
C39094 OR2X1_LOC_405/A OR2X1_LOC_532/B 0.30fF
C39095 OR2X1_LOC_595/A AND2X1_LOC_217/a_36_24# 0.00fF
C39096 OR2X1_LOC_287/B OR2X1_LOC_402/a_36_216# -0.00fF
C39097 OR2X1_LOC_426/A OR2X1_LOC_426/a_36_216# 0.00fF
C39098 AND2X1_LOC_392/A AND2X1_LOC_222/Y 0.03fF
C39099 AND2X1_LOC_544/a_8_24# OR2X1_LOC_47/Y 0.01fF
C39100 AND2X1_LOC_662/a_36_24# OR2X1_LOC_52/B 0.01fF
C39101 AND2X1_LOC_44/a_8_24# AND2X1_LOC_51/Y 0.01fF
C39102 OR2X1_LOC_831/B AND2X1_LOC_36/Y 0.16fF
C39103 OR2X1_LOC_712/B OR2X1_LOC_779/A 0.00fF
C39104 AND2X1_LOC_476/A AND2X1_LOC_649/a_8_24# 0.02fF
C39105 AND2X1_LOC_663/B OR2X1_LOC_757/a_8_216# 0.01fF
C39106 AND2X1_LOC_139/B D_INPUT_0 0.15fF
C39107 OR2X1_LOC_70/A OR2X1_LOC_585/Y 0.01fF
C39108 OR2X1_LOC_19/B AND2X1_LOC_852/Y 0.07fF
C39109 AND2X1_LOC_59/Y AND2X1_LOC_108/a_8_24# 0.07fF
C39110 AND2X1_LOC_656/Y OR2X1_LOC_65/B 0.54fF
C39111 OR2X1_LOC_71/Y OR2X1_LOC_265/Y 0.01fF
C39112 OR2X1_LOC_576/A OR2X1_LOC_576/a_8_216# 0.16fF
C39113 OR2X1_LOC_694/a_8_216# OR2X1_LOC_31/Y 0.01fF
C39114 OR2X1_LOC_83/Y OR2X1_LOC_19/B 0.01fF
C39115 AND2X1_LOC_845/Y OR2X1_LOC_67/a_36_216# 0.03fF
C39116 AND2X1_LOC_680/a_36_24# OR2X1_LOC_449/B 0.00fF
C39117 OR2X1_LOC_490/Y AND2X1_LOC_663/B 0.10fF
C39118 OR2X1_LOC_742/B OR2X1_LOC_741/Y 0.03fF
C39119 AND2X1_LOC_687/B OR2X1_LOC_52/B 0.08fF
C39120 OR2X1_LOC_803/A OR2X1_LOC_160/a_8_216# 0.01fF
C39121 AND2X1_LOC_494/a_8_24# OR2X1_LOC_269/B 0.01fF
C39122 OR2X1_LOC_715/B OR2X1_LOC_446/B 0.20fF
C39123 AND2X1_LOC_69/Y OR2X1_LOC_202/a_8_216# 0.47fF
C39124 OR2X1_LOC_51/Y AND2X1_LOC_657/A 0.02fF
C39125 OR2X1_LOC_46/A AND2X1_LOC_412/a_36_24# 0.00fF
C39126 AND2X1_LOC_133/a_36_24# AND2X1_LOC_8/Y 0.00fF
C39127 OR2X1_LOC_121/B OR2X1_LOC_794/a_8_216# -0.00fF
C39128 OR2X1_LOC_256/A OR2X1_LOC_85/A 0.34fF
C39129 AND2X1_LOC_648/B OR2X1_LOC_433/Y 0.01fF
C39130 AND2X1_LOC_436/Y OR2X1_LOC_533/A 0.02fF
C39131 AND2X1_LOC_56/B AND2X1_LOC_56/a_8_24# 0.11fF
C39132 AND2X1_LOC_580/A OR2X1_LOC_95/Y 0.03fF
C39133 OR2X1_LOC_121/Y OR2X1_LOC_217/A 0.01fF
C39134 AND2X1_LOC_40/Y OR2X1_LOC_339/Y 0.03fF
C39135 AND2X1_LOC_660/A OR2X1_LOC_39/A 0.07fF
C39136 AND2X1_LOC_72/B OR2X1_LOC_575/A 0.03fF
C39137 AND2X1_LOC_687/Y OR2X1_LOC_7/A 0.00fF
C39138 OR2X1_LOC_12/Y OR2X1_LOC_320/a_8_216# 0.02fF
C39139 OR2X1_LOC_31/Y AND2X1_LOC_650/Y 0.03fF
C39140 OR2X1_LOC_234/a_8_216# OR2X1_LOC_619/Y 0.03fF
C39141 AND2X1_LOC_663/B OR2X1_LOC_261/A 0.02fF
C39142 OR2X1_LOC_59/Y OR2X1_LOC_534/Y 0.25fF
C39143 OR2X1_LOC_850/B OR2X1_LOC_675/Y 0.03fF
C39144 OR2X1_LOC_840/a_36_216# OR2X1_LOC_723/B 0.02fF
C39145 OR2X1_LOC_344/A AND2X1_LOC_36/Y 0.12fF
C39146 OR2X1_LOC_89/A OR2X1_LOC_226/a_8_216# 0.01fF
C39147 VDD OR2X1_LOC_732/A 0.30fF
C39148 OR2X1_LOC_756/B OR2X1_LOC_68/B 0.10fF
C39149 AND2X1_LOC_175/a_8_24# OR2X1_LOC_31/Y 0.06fF
C39150 OR2X1_LOC_11/Y OR2X1_LOC_588/A 0.02fF
C39151 AND2X1_LOC_729/B OR2X1_LOC_46/A 0.02fF
C39152 AND2X1_LOC_810/A OR2X1_LOC_696/A 0.03fF
C39153 OR2X1_LOC_448/A OR2X1_LOC_779/B 0.03fF
C39154 OR2X1_LOC_485/A AND2X1_LOC_800/a_36_24# 0.00fF
C39155 OR2X1_LOC_66/A OR2X1_LOC_788/B 0.06fF
C39156 OR2X1_LOC_43/A OR2X1_LOC_47/Y 0.18fF
C39157 OR2X1_LOC_89/A OR2X1_LOC_55/a_8_216# 0.01fF
C39158 OR2X1_LOC_180/a_36_216# OR2X1_LOC_180/B 0.02fF
C39159 OR2X1_LOC_280/Y OR2X1_LOC_238/a_36_216# 0.00fF
C39160 OR2X1_LOC_185/A OR2X1_LOC_318/B 3.55fF
C39161 OR2X1_LOC_686/A AND2X1_LOC_36/Y 0.25fF
C39162 AND2X1_LOC_102/a_8_24# OR2X1_LOC_673/A 0.01fF
C39163 OR2X1_LOC_156/B OR2X1_LOC_156/a_8_216# 0.39fF
C39164 OR2X1_LOC_272/Y OR2X1_LOC_31/Y 0.03fF
C39165 AND2X1_LOC_624/A OR2X1_LOC_406/A 0.06fF
C39166 OR2X1_LOC_85/A OR2X1_LOC_67/Y 0.17fF
C39167 AND2X1_LOC_338/A OR2X1_LOC_171/Y 0.28fF
C39168 OR2X1_LOC_45/B AND2X1_LOC_564/B 0.30fF
C39169 OR2X1_LOC_375/A OR2X1_LOC_192/B 0.01fF
C39170 VDD OR2X1_LOC_539/B 0.31fF
C39171 OR2X1_LOC_476/B OR2X1_LOC_814/A 0.03fF
C39172 OR2X1_LOC_45/B OR2X1_LOC_230/Y 0.03fF
C39173 OR2X1_LOC_3/B OR2X1_LOC_22/a_8_216# 0.04fF
C39174 AND2X1_LOC_514/a_36_24# OR2X1_LOC_437/A 0.01fF
C39175 OR2X1_LOC_66/A OR2X1_LOC_175/a_8_216# 0.00fF
C39176 OR2X1_LOC_235/B OR2X1_LOC_140/Y 0.00fF
C39177 OR2X1_LOC_19/B OR2X1_LOC_243/B 0.26fF
C39178 OR2X1_LOC_121/a_8_216# AND2X1_LOC_7/B 0.02fF
C39179 AND2X1_LOC_810/A AND2X1_LOC_715/Y -0.00fF
C39180 AND2X1_LOC_86/a_8_24# AND2X1_LOC_235/a_8_24# 0.23fF
C39181 OR2X1_LOC_497/Y OR2X1_LOC_419/Y 0.49fF
C39182 AND2X1_LOC_660/a_36_24# AND2X1_LOC_663/B 0.01fF
C39183 OR2X1_LOC_185/A OR2X1_LOC_344/a_36_216# 0.00fF
C39184 AND2X1_LOC_574/A AND2X1_LOC_657/a_36_24# 0.01fF
C39185 OR2X1_LOC_118/Y AND2X1_LOC_217/a_8_24# 0.01fF
C39186 OR2X1_LOC_97/A OR2X1_LOC_435/A 0.01fF
C39187 OR2X1_LOC_406/Y AND2X1_LOC_475/Y 0.00fF
C39188 OR2X1_LOC_680/A AND2X1_LOC_657/A 0.12fF
C39189 AND2X1_LOC_55/a_8_24# OR2X1_LOC_68/B 0.01fF
C39190 OR2X1_LOC_177/Y OR2X1_LOC_373/a_36_216# 0.00fF
C39191 AND2X1_LOC_555/Y VDD 0.27fF
C39192 AND2X1_LOC_209/a_8_24# AND2X1_LOC_220/B 0.10fF
C39193 AND2X1_LOC_47/Y D_INPUT_0 0.10fF
C39194 AND2X1_LOC_18/Y OR2X1_LOC_563/A 0.05fF
C39195 OR2X1_LOC_862/a_8_216# VDD 0.00fF
C39196 AND2X1_LOC_340/Y OR2X1_LOC_158/A 0.07fF
C39197 OR2X1_LOC_136/Y VDD 0.27fF
C39198 OR2X1_LOC_158/A AND2X1_LOC_810/B 0.07fF
C39199 OR2X1_LOC_78/B OR2X1_LOC_502/Y 0.01fF
C39200 OR2X1_LOC_421/A OR2X1_LOC_428/A 2.69fF
C39201 OR2X1_LOC_527/a_8_216# AND2X1_LOC_786/Y 0.01fF
C39202 AND2X1_LOC_729/B OR2X1_LOC_41/Y 0.02fF
C39203 AND2X1_LOC_22/Y OR2X1_LOC_66/A 0.70fF
C39204 OR2X1_LOC_487/a_8_216# AND2X1_LOC_563/Y 0.01fF
C39205 OR2X1_LOC_19/B AND2X1_LOC_647/B 0.13fF
C39206 OR2X1_LOC_158/A AND2X1_LOC_181/Y 0.01fF
C39207 AND2X1_LOC_22/Y OR2X1_LOC_841/A 0.03fF
C39208 OR2X1_LOC_269/B OR2X1_LOC_725/a_8_216# 0.01fF
C39209 OR2X1_LOC_632/Y OR2X1_LOC_554/a_8_216# 0.40fF
C39210 OR2X1_LOC_37/a_8_216# OR2X1_LOC_80/A 0.47fF
C39211 OR2X1_LOC_335/A OR2X1_LOC_808/A 0.14fF
C39212 AND2X1_LOC_563/A OR2X1_LOC_595/A 0.05fF
C39213 AND2X1_LOC_40/Y OR2X1_LOC_731/A 0.46fF
C39214 OR2X1_LOC_44/Y OR2X1_LOC_437/A 0.35fF
C39215 OR2X1_LOC_757/A GATE_579 0.00fF
C39216 OR2X1_LOC_662/a_8_216# OR2X1_LOC_227/B 0.47fF
C39217 AND2X1_LOC_67/Y AND2X1_LOC_31/Y 0.02fF
C39218 OR2X1_LOC_70/Y OR2X1_LOC_534/Y 0.01fF
C39219 OR2X1_LOC_532/B OR2X1_LOC_330/a_8_216# 0.01fF
C39220 OR2X1_LOC_87/A OR2X1_LOC_590/Y 0.07fF
C39221 OR2X1_LOC_417/A AND2X1_LOC_792/Y 0.01fF
C39222 OR2X1_LOC_6/B AND2X1_LOC_131/a_8_24# 0.04fF
C39223 AND2X1_LOC_794/B OR2X1_LOC_51/Y 0.02fF
C39224 OR2X1_LOC_269/B OR2X1_LOC_537/a_8_216# 0.05fF
C39225 OR2X1_LOC_294/Y OR2X1_LOC_78/A 0.05fF
C39226 D_INPUT_0 OR2X1_LOC_598/A 7.74fF
C39227 OR2X1_LOC_590/a_36_216# OR2X1_LOC_814/A 0.01fF
C39228 AND2X1_LOC_456/B OR2X1_LOC_428/A 0.02fF
C39229 AND2X1_LOC_774/a_36_24# OR2X1_LOC_91/A 0.00fF
C39230 OR2X1_LOC_45/B AND2X1_LOC_857/Y 0.22fF
C39231 OR2X1_LOC_151/Y OR2X1_LOC_209/A 0.79fF
C39232 OR2X1_LOC_546/B OR2X1_LOC_546/a_8_216# 0.47fF
C39233 OR2X1_LOC_227/a_8_216# OR2X1_LOC_68/B 0.02fF
C39234 OR2X1_LOC_147/B OR2X1_LOC_577/Y 0.06fF
C39235 OR2X1_LOC_78/A OR2X1_LOC_641/A 0.03fF
C39236 OR2X1_LOC_65/B AND2X1_LOC_772/Y 0.44fF
C39237 AND2X1_LOC_787/A AND2X1_LOC_723/a_8_24# 0.01fF
C39238 OR2X1_LOC_516/Y AND2X1_LOC_500/a_8_24# 0.04fF
C39239 OR2X1_LOC_860/a_8_216# OR2X1_LOC_474/B 0.00fF
C39240 AND2X1_LOC_91/B AND2X1_LOC_767/a_8_24# 0.04fF
C39241 OR2X1_LOC_144/Y OR2X1_LOC_12/Y 0.08fF
C39242 VDD OR2X1_LOC_51/Y 1.94fF
C39243 OR2X1_LOC_528/Y AND2X1_LOC_675/Y 0.06fF
C39244 AND2X1_LOC_64/Y OR2X1_LOC_703/B 0.01fF
C39245 OR2X1_LOC_40/Y OR2X1_LOC_12/a_36_216# 0.00fF
C39246 OR2X1_LOC_122/a_36_216# AND2X1_LOC_243/Y 0.01fF
C39247 AND2X1_LOC_539/Y AND2X1_LOC_436/B 0.10fF
C39248 OR2X1_LOC_494/Y OR2X1_LOC_666/A 0.06fF
C39249 AND2X1_LOC_721/Y OR2X1_LOC_18/Y 0.25fF
C39250 D_INPUT_1 OR2X1_LOC_241/B 0.07fF
C39251 AND2X1_LOC_733/Y AND2X1_LOC_443/a_36_24# 0.00fF
C39252 AND2X1_LOC_3/Y INPUT_6 0.01fF
C39253 OR2X1_LOC_177/Y AND2X1_LOC_374/a_8_24# 0.01fF
C39254 AND2X1_LOC_436/Y AND2X1_LOC_468/a_8_24# 0.10fF
C39255 VDD OR2X1_LOC_78/B 2.12fF
C39256 AND2X1_LOC_722/Y OR2X1_LOC_40/Y 0.01fF
C39257 AND2X1_LOC_776/Y AND2X1_LOC_840/B 0.10fF
C39258 OR2X1_LOC_149/B OR2X1_LOC_213/A 1.83fF
C39259 AND2X1_LOC_64/Y OR2X1_LOC_87/A 0.46fF
C39260 AND2X1_LOC_133/a_8_24# OR2X1_LOC_71/A 0.01fF
C39261 AND2X1_LOC_7/B OR2X1_LOC_541/a_8_216# 0.02fF
C39262 AND2X1_LOC_305/a_8_24# OR2X1_LOC_161/B 0.09fF
C39263 OR2X1_LOC_500/A OR2X1_LOC_563/A 0.01fF
C39264 AND2X1_LOC_745/a_8_24# AND2X1_LOC_40/Y 0.09fF
C39265 AND2X1_LOC_811/B AND2X1_LOC_727/B 0.09fF
C39266 OR2X1_LOC_134/a_8_216# AND2X1_LOC_361/A 0.04fF
C39267 AND2X1_LOC_392/A AND2X1_LOC_367/A 0.07fF
C39268 OR2X1_LOC_154/A OR2X1_LOC_175/Y 0.04fF
C39269 OR2X1_LOC_458/B OR2X1_LOC_733/A 0.02fF
C39270 OR2X1_LOC_244/B OR2X1_LOC_66/A 0.25fF
C39271 AND2X1_LOC_40/Y OR2X1_LOC_596/a_8_216# 0.09fF
C39272 OR2X1_LOC_653/A OR2X1_LOC_392/B 0.12fF
C39273 OR2X1_LOC_541/B AND2X1_LOC_255/a_8_24# 0.01fF
C39274 OR2X1_LOC_505/a_8_216# AND2X1_LOC_862/A 0.47fF
C39275 OR2X1_LOC_308/A OR2X1_LOC_269/B 0.00fF
C39276 AND2X1_LOC_576/Y AND2X1_LOC_242/B 0.02fF
C39277 AND2X1_LOC_40/Y OR2X1_LOC_6/B 0.10fF
C39278 OR2X1_LOC_161/A OR2X1_LOC_580/B 0.03fF
C39279 OR2X1_LOC_214/a_8_216# OR2X1_LOC_214/A 0.39fF
C39280 AND2X1_LOC_364/Y OR2X1_LOC_56/A 0.15fF
C39281 AND2X1_LOC_716/Y AND2X1_LOC_357/B 0.03fF
C39282 AND2X1_LOC_799/a_8_24# AND2X1_LOC_661/A 0.21fF
C39283 OR2X1_LOC_427/A OR2X1_LOC_584/Y 0.03fF
C39284 OR2X1_LOC_19/B OR2X1_LOC_771/B 0.03fF
C39285 OR2X1_LOC_456/A AND2X1_LOC_36/Y 0.15fF
C39286 OR2X1_LOC_154/A OR2X1_LOC_691/Y 0.03fF
C39287 OR2X1_LOC_673/Y AND2X1_LOC_263/a_8_24# 0.01fF
C39288 OR2X1_LOC_866/B OR2X1_LOC_269/B 0.01fF
C39289 OR2X1_LOC_318/A OR2X1_LOC_130/A 0.03fF
C39290 OR2X1_LOC_62/A OR2X1_LOC_80/A 0.09fF
C39291 VDD OR2X1_LOC_721/Y 1.36fF
C39292 OR2X1_LOC_677/Y OR2X1_LOC_51/Y 0.02fF
C39293 OR2X1_LOC_62/B AND2X1_LOC_246/a_8_24# 0.09fF
C39294 OR2X1_LOC_6/A OR2X1_LOC_310/a_36_216# 0.03fF
C39295 AND2X1_LOC_357/B AND2X1_LOC_654/Y 0.02fF
C39296 AND2X1_LOC_566/B AND2X1_LOC_662/B 0.02fF
C39297 VDD OR2X1_LOC_16/Y 0.06fF
C39298 OR2X1_LOC_482/Y OR2X1_LOC_18/Y 0.03fF
C39299 AND2X1_LOC_535/Y AND2X1_LOC_841/B 0.07fF
C39300 INPUT_0 AND2X1_LOC_41/A 0.10fF
C39301 OR2X1_LOC_160/B OR2X1_LOC_856/B 0.05fF
C39302 AND2X1_LOC_621/Y AND2X1_LOC_477/Y 0.07fF
C39303 OR2X1_LOC_106/Y AND2X1_LOC_554/B 0.14fF
C39304 AND2X1_LOC_764/a_8_24# OR2X1_LOC_502/A 0.01fF
C39305 OR2X1_LOC_6/B OR2X1_LOC_399/A 0.01fF
C39306 AND2X1_LOC_366/A AND2X1_LOC_367/A 0.49fF
C39307 OR2X1_LOC_744/A OR2X1_LOC_594/a_8_216# 0.01fF
C39308 AND2X1_LOC_370/a_8_24# AND2X1_LOC_211/B 0.04fF
C39309 OR2X1_LOC_790/A AND2X1_LOC_43/B 0.02fF
C39310 OR2X1_LOC_686/B AND2X1_LOC_682/a_8_24# 0.04fF
C39311 AND2X1_LOC_856/A OR2X1_LOC_428/A 0.07fF
C39312 OR2X1_LOC_151/A OR2X1_LOC_130/A 0.07fF
C39313 AND2X1_LOC_107/a_8_24# OR2X1_LOC_844/B 0.00fF
C39314 OR2X1_LOC_40/Y AND2X1_LOC_676/a_36_24# 0.01fF
C39315 OR2X1_LOC_662/a_36_216# OR2X1_LOC_663/A 0.00fF
C39316 OR2X1_LOC_630/Y OR2X1_LOC_575/A 0.01fF
C39317 AND2X1_LOC_784/Y OR2X1_LOC_91/Y 0.01fF
C39318 AND2X1_LOC_512/Y OR2X1_LOC_516/B 0.02fF
C39319 OR2X1_LOC_519/Y AND2X1_LOC_326/B 0.02fF
C39320 OR2X1_LOC_371/a_36_216# AND2X1_LOC_786/Y 0.01fF
C39321 OR2X1_LOC_40/Y INPUT_4 0.00fF
C39322 OR2X1_LOC_137/B AND2X1_LOC_18/Y 0.03fF
C39323 OR2X1_LOC_6/B OR2X1_LOC_87/Y 0.03fF
C39324 AND2X1_LOC_486/Y AND2X1_LOC_474/A 0.03fF
C39325 AND2X1_LOC_716/Y AND2X1_LOC_303/a_8_24# 0.01fF
C39326 AND2X1_LOC_59/Y OR2X1_LOC_440/a_8_216# 0.02fF
C39327 OR2X1_LOC_600/A AND2X1_LOC_114/a_8_24# 0.05fF
C39328 OR2X1_LOC_715/B AND2X1_LOC_56/B 0.14fF
C39329 AND2X1_LOC_222/Y AND2X1_LOC_223/a_8_24# 0.04fF
C39330 INPUT_0 AND2X1_LOC_649/a_8_24# 0.14fF
C39331 OR2X1_LOC_655/a_8_216# AND2X1_LOC_92/Y 0.01fF
C39332 AND2X1_LOC_56/B AND2X1_LOC_626/a_8_24# 0.01fF
C39333 VDD OR2X1_LOC_375/A 2.44fF
C39334 OR2X1_LOC_151/A AND2X1_LOC_292/a_8_24# 0.01fF
C39335 OR2X1_LOC_420/Y OR2X1_LOC_12/Y 0.02fF
C39336 VDD OR2X1_LOC_680/A 0.31fF
C39337 AND2X1_LOC_95/Y AND2X1_LOC_94/Y 0.05fF
C39338 OR2X1_LOC_622/a_8_216# OR2X1_LOC_633/A 0.05fF
C39339 AND2X1_LOC_56/B OR2X1_LOC_543/A 0.00fF
C39340 OR2X1_LOC_744/A AND2X1_LOC_468/B 0.38fF
C39341 AND2X1_LOC_70/Y AND2X1_LOC_601/a_8_24# 0.01fF
C39342 OR2X1_LOC_158/A OR2X1_LOC_585/A 0.14fF
C39343 OR2X1_LOC_60/Y OR2X1_LOC_85/A 0.01fF
C39344 OR2X1_LOC_604/A OR2X1_LOC_497/Y 0.10fF
C39345 OR2X1_LOC_538/A OR2X1_LOC_185/A 0.03fF
C39346 AND2X1_LOC_764/a_36_24# OR2X1_LOC_160/A 0.01fF
C39347 D_INPUT_0 OR2X1_LOC_186/a_8_216# 0.01fF
C39348 AND2X1_LOC_565/B AND2X1_LOC_564/a_8_24# 0.17fF
C39349 AND2X1_LOC_547/Y AND2X1_LOC_569/A 0.01fF
C39350 OR2X1_LOC_96/Y OR2X1_LOC_26/Y 0.00fF
C39351 OR2X1_LOC_243/A AND2X1_LOC_232/a_8_24# 0.23fF
C39352 OR2X1_LOC_240/B AND2X1_LOC_232/a_36_24# 0.00fF
C39353 OR2X1_LOC_64/Y OR2X1_LOC_816/A 0.04fF
C39354 OR2X1_LOC_154/A OR2X1_LOC_803/A 0.00fF
C39355 OR2X1_LOC_518/a_8_216# AND2X1_LOC_831/Y 0.03fF
C39356 AND2X1_LOC_363/Y GATE_366 0.01fF
C39357 VDD OR2X1_LOC_667/a_8_216# 0.21fF
C39358 AND2X1_LOC_42/B AND2X1_LOC_65/A 0.01fF
C39359 OR2X1_LOC_599/A AND2X1_LOC_447/Y 0.05fF
C39360 AND2X1_LOC_72/B OR2X1_LOC_735/B 0.01fF
C39361 AND2X1_LOC_566/B AND2X1_LOC_337/B 0.00fF
C39362 OR2X1_LOC_527/Y AND2X1_LOC_795/a_8_24# 0.04fF
C39363 OR2X1_LOC_64/Y OR2X1_LOC_79/Y 0.02fF
C39364 AND2X1_LOC_252/a_8_24# AND2X1_LOC_18/Y 0.01fF
C39365 OR2X1_LOC_656/a_8_216# AND2X1_LOC_44/Y 0.05fF
C39366 AND2X1_LOC_710/a_36_24# AND2X1_LOC_866/A 0.07fF
C39367 OR2X1_LOC_804/A OR2X1_LOC_716/a_8_216# 0.05fF
C39368 AND2X1_LOC_59/Y OR2X1_LOC_78/Y 0.03fF
C39369 AND2X1_LOC_737/Y OR2X1_LOC_427/A 0.05fF
C39370 AND2X1_LOC_59/Y OR2X1_LOC_274/a_8_216# 0.01fF
C39371 OR2X1_LOC_411/Y OR2X1_LOC_44/Y 0.03fF
C39372 AND2X1_LOC_50/Y AND2X1_LOC_95/Y 0.01fF
C39373 AND2X1_LOC_31/Y OR2X1_LOC_365/a_8_216# 0.06fF
C39374 OR2X1_LOC_114/Y OR2X1_LOC_78/A 0.02fF
C39375 OR2X1_LOC_807/Y OR2X1_LOC_792/Y 0.42fF
C39376 OR2X1_LOC_334/B AND2X1_LOC_824/B 0.00fF
C39377 OR2X1_LOC_634/A AND2X1_LOC_291/a_8_24# 0.02fF
C39378 AND2X1_LOC_388/Y OR2X1_LOC_70/Y 0.70fF
C39379 OR2X1_LOC_506/A AND2X1_LOC_423/a_8_24# 0.20fF
C39380 OR2X1_LOC_676/Y OR2X1_LOC_574/A 0.18fF
C39381 OR2X1_LOC_251/Y OR2X1_LOC_51/Y 0.26fF
C39382 OR2X1_LOC_48/B OR2X1_LOC_586/Y 0.07fF
C39383 OR2X1_LOC_330/Y OR2X1_LOC_739/A 0.01fF
C39384 OR2X1_LOC_516/A OR2X1_LOC_516/B 0.66fF
C39385 OR2X1_LOC_405/A OR2X1_LOC_734/a_8_216# 0.05fF
C39386 AND2X1_LOC_217/Y OR2X1_LOC_131/Y 0.00fF
C39387 OR2X1_LOC_220/A OR2X1_LOC_739/A 0.03fF
C39388 AND2X1_LOC_392/A OR2X1_LOC_490/Y 0.07fF
C39389 AND2X1_LOC_392/A OR2X1_LOC_74/A 0.07fF
C39390 OR2X1_LOC_26/Y AND2X1_LOC_663/A 0.03fF
C39391 OR2X1_LOC_680/A OR2X1_LOC_677/Y 0.01fF
C39392 OR2X1_LOC_723/B OR2X1_LOC_374/Y 0.32fF
C39393 AND2X1_LOC_658/B AND2X1_LOC_147/Y 0.03fF
C39394 AND2X1_LOC_212/A OR2X1_LOC_64/Y 0.50fF
C39395 OR2X1_LOC_18/Y OR2X1_LOC_586/Y 0.42fF
C39396 OR2X1_LOC_810/A AND2X1_LOC_92/Y 0.07fF
C39397 D_INPUT_0 OR2X1_LOC_34/A 0.27fF
C39398 OR2X1_LOC_755/Y OR2X1_LOC_44/Y 0.02fF
C39399 OR2X1_LOC_417/A AND2X1_LOC_287/B 0.03fF
C39400 AND2X1_LOC_735/a_8_24# AND2X1_LOC_191/Y 0.07fF
C39401 OR2X1_LOC_648/B AND2X1_LOC_51/Y 1.65fF
C39402 OR2X1_LOC_648/A AND2X1_LOC_3/Y 0.07fF
C39403 OR2X1_LOC_185/A AND2X1_LOC_178/a_8_24# 0.00fF
C39404 VDD OR2X1_LOC_605/B 0.00fF
C39405 OR2X1_LOC_73/a_8_216# OR2X1_LOC_56/A 0.01fF
C39406 AND2X1_LOC_173/a_36_24# OR2X1_LOC_161/A 0.01fF
C39407 OR2X1_LOC_417/A OR2X1_LOC_816/A 0.02fF
C39408 OR2X1_LOC_680/Y AND2X1_LOC_658/A 0.03fF
C39409 AND2X1_LOC_799/a_8_24# AND2X1_LOC_810/Y 0.10fF
C39410 AND2X1_LOC_705/Y AND2X1_LOC_477/A 0.26fF
C39411 AND2X1_LOC_70/Y OR2X1_LOC_446/a_8_216# 0.01fF
C39412 OR2X1_LOC_656/Y OR2X1_LOC_87/A 0.00fF
C39413 OR2X1_LOC_40/Y OR2X1_LOC_277/a_8_216# 0.06fF
C39414 OR2X1_LOC_316/Y AND2X1_LOC_520/Y 0.02fF
C39415 AND2X1_LOC_191/B OR2X1_LOC_258/Y 0.03fF
C39416 OR2X1_LOC_3/Y OR2X1_LOC_59/Y 0.84fF
C39417 AND2X1_LOC_98/Y OR2X1_LOC_585/A 0.02fF
C39418 OR2X1_LOC_639/a_8_216# AND2X1_LOC_44/Y 0.01fF
C39419 OR2X1_LOC_151/A OR2X1_LOC_62/B 0.11fF
C39420 AND2X1_LOC_12/Y OR2X1_LOC_185/A 0.07fF
C39421 AND2X1_LOC_196/a_8_24# OR2X1_LOC_56/A 0.03fF
C39422 OR2X1_LOC_423/Y OR2X1_LOC_589/Y 0.25fF
C39423 AND2X1_LOC_47/Y AND2X1_LOC_438/a_8_24# 0.01fF
C39424 AND2X1_LOC_260/a_8_24# OR2X1_LOC_56/A 0.01fF
C39425 AND2X1_LOC_866/A OR2X1_LOC_759/a_8_216# 0.02fF
C39426 OR2X1_LOC_201/Y OR2X1_LOC_78/A 0.00fF
C39427 AND2X1_LOC_711/Y AND2X1_LOC_501/a_36_24# 0.01fF
C39428 AND2X1_LOC_631/Y OR2X1_LOC_59/Y 0.03fF
C39429 AND2X1_LOC_707/a_8_24# OR2X1_LOC_64/Y 0.11fF
C39430 AND2X1_LOC_563/a_8_24# AND2X1_LOC_573/A 0.03fF
C39431 OR2X1_LOC_673/B AND2X1_LOC_47/Y 0.02fF
C39432 OR2X1_LOC_154/A AND2X1_LOC_699/a_36_24# 0.01fF
C39433 AND2X1_LOC_120/a_8_24# AND2X1_LOC_858/B 0.02fF
C39434 AND2X1_LOC_448/Y AND2X1_LOC_454/Y 0.37fF
C39435 AND2X1_LOC_449/Y AND2X1_LOC_453/Y 0.03fF
C39436 OR2X1_LOC_154/A OR2X1_LOC_249/a_8_216# 0.17fF
C39437 OR2X1_LOC_185/A OR2X1_LOC_802/A 0.10fF
C39438 AND2X1_LOC_212/A OR2X1_LOC_417/A 0.01fF
C39439 OR2X1_LOC_335/A OR2X1_LOC_374/Y 0.03fF
C39440 OR2X1_LOC_426/A OR2X1_LOC_7/A 0.01fF
C39441 AND2X1_LOC_103/a_8_24# AND2X1_LOC_51/Y 0.01fF
C39442 OR2X1_LOC_680/A OR2X1_LOC_616/Y 0.03fF
C39443 OR2X1_LOC_831/A AND2X1_LOC_47/Y 0.01fF
C39444 OR2X1_LOC_450/A AND2X1_LOC_425/Y 0.00fF
C39445 OR2X1_LOC_759/A OR2X1_LOC_815/A 0.01fF
C39446 AND2X1_LOC_84/Y AND2X1_LOC_204/Y 0.01fF
C39447 OR2X1_LOC_462/B OR2X1_LOC_39/A 0.17fF
C39448 OR2X1_LOC_844/Y OR2X1_LOC_78/A 0.04fF
C39449 OR2X1_LOC_385/Y OR2X1_LOC_586/Y 0.30fF
C39450 OR2X1_LOC_744/A OR2X1_LOC_278/A 0.15fF
C39451 OR2X1_LOC_216/Y OR2X1_LOC_805/A 0.12fF
C39452 OR2X1_LOC_730/a_8_216# OR2X1_LOC_155/A 0.02fF
C39453 OR2X1_LOC_311/Y AND2X1_LOC_434/Y 0.15fF
C39454 OR2X1_LOC_32/B OR2X1_LOC_69/Y 0.13fF
C39455 OR2X1_LOC_269/Y OR2X1_LOC_344/A 0.01fF
C39456 OR2X1_LOC_495/a_36_216# OR2X1_LOC_39/A 0.00fF
C39457 AND2X1_LOC_849/a_8_24# AND2X1_LOC_860/A 0.20fF
C39458 OR2X1_LOC_467/A OR2X1_LOC_707/B 0.01fF
C39459 OR2X1_LOC_280/Y OR2X1_LOC_427/A 0.23fF
C39460 INPUT_0 AND2X1_LOC_727/A 0.03fF
C39461 AND2X1_LOC_538/Y AND2X1_LOC_434/Y -0.01fF
C39462 AND2X1_LOC_638/Y OR2X1_LOC_762/a_8_216# 0.48fF
C39463 OR2X1_LOC_83/A AND2X1_LOC_43/B 0.01fF
C39464 AND2X1_LOC_714/B AND2X1_LOC_648/B 0.03fF
C39465 AND2X1_LOC_703/a_36_24# OR2X1_LOC_485/A 0.00fF
C39466 AND2X1_LOC_112/a_8_24# AND2X1_LOC_831/Y 0.01fF
C39467 OR2X1_LOC_251/a_8_216# OR2X1_LOC_64/Y 0.01fF
C39468 OR2X1_LOC_485/A OR2X1_LOC_71/a_8_216# 0.03fF
C39469 OR2X1_LOC_160/A OR2X1_LOC_646/A 0.03fF
C39470 AND2X1_LOC_72/B OR2X1_LOC_161/B 0.03fF
C39471 AND2X1_LOC_497/a_8_24# AND2X1_LOC_44/Y 0.01fF
C39472 OR2X1_LOC_140/B OR2X1_LOC_68/B 0.03fF
C39473 AND2X1_LOC_728/Y OR2X1_LOC_189/Y 0.03fF
C39474 AND2X1_LOC_331/a_8_24# AND2X1_LOC_51/Y 0.02fF
C39475 OR2X1_LOC_185/A AND2X1_LOC_79/Y 0.01fF
C39476 OR2X1_LOC_248/Y OR2X1_LOC_85/A 0.12fF
C39477 AND2X1_LOC_348/Y OR2X1_LOC_44/Y 0.03fF
C39478 OR2X1_LOC_51/Y OR2X1_LOC_256/A 0.07fF
C39479 AND2X1_LOC_784/A OR2X1_LOC_6/A 0.04fF
C39480 OR2X1_LOC_161/B OR2X1_LOC_451/B 0.02fF
C39481 OR2X1_LOC_296/Y AND2X1_LOC_297/a_8_24# 0.00fF
C39482 OR2X1_LOC_283/a_8_216# OR2X1_LOC_26/Y 0.03fF
C39483 OR2X1_LOC_482/Y AND2X1_LOC_620/Y 0.00fF
C39484 OR2X1_LOC_304/Y OR2X1_LOC_48/B 0.21fF
C39485 OR2X1_LOC_473/Y OR2X1_LOC_737/A 0.00fF
C39486 AND2X1_LOC_728/Y OR2X1_LOC_152/Y 0.00fF
C39487 OR2X1_LOC_530/Y AND2X1_LOC_624/A 0.06fF
C39488 OR2X1_LOC_753/A OR2X1_LOC_44/Y 0.12fF
C39489 OR2X1_LOC_194/Y OR2X1_LOC_155/A 0.03fF
C39490 AND2X1_LOC_660/a_8_24# OR2X1_LOC_56/A 0.07fF
C39491 AND2X1_LOC_300/a_8_24# OR2X1_LOC_804/A -0.01fF
C39492 OR2X1_LOC_251/Y OR2X1_LOC_667/a_8_216# 0.04fF
C39493 AND2X1_LOC_95/Y OR2X1_LOC_473/Y 0.15fF
C39494 OR2X1_LOC_327/a_8_216# OR2X1_LOC_121/B 0.01fF
C39495 OR2X1_LOC_141/B OR2X1_LOC_657/a_36_216# 0.00fF
C39496 AND2X1_LOC_702/a_36_24# OR2X1_LOC_304/Y 0.01fF
C39497 AND2X1_LOC_514/Y AND2X1_LOC_364/A 0.03fF
C39498 OR2X1_LOC_51/Y OR2X1_LOC_674/Y 0.01fF
C39499 AND2X1_LOC_126/a_36_24# OR2X1_LOC_243/B 0.00fF
C39500 INPUT_0 OR2X1_LOC_95/Y 0.02fF
C39501 OR2X1_LOC_335/Y AND2X1_LOC_47/Y 0.03fF
C39502 AND2X1_LOC_784/A OR2X1_LOC_299/a_8_216# 0.47fF
C39503 OR2X1_LOC_449/A OR2X1_LOC_155/A 0.16fF
C39504 AND2X1_LOC_183/a_8_24# OR2X1_LOC_456/Y 0.08fF
C39505 OR2X1_LOC_517/a_8_216# OR2X1_LOC_31/Y 0.05fF
C39506 D_INPUT_0 AND2X1_LOC_240/a_36_24# 0.01fF
C39507 OR2X1_LOC_64/Y AND2X1_LOC_843/a_8_24# 0.16fF
C39508 OR2X1_LOC_22/Y OR2X1_LOC_427/A 0.64fF
C39509 OR2X1_LOC_691/Y OR2X1_LOC_198/A 0.45fF
C39510 OR2X1_LOC_562/A OR2X1_LOC_366/Y 0.03fF
C39511 OR2X1_LOC_862/B D_INPUT_1 0.40fF
C39512 OR2X1_LOC_557/A OR2X1_LOC_269/B 0.16fF
C39513 OR2X1_LOC_3/Y OR2X1_LOC_820/B 0.05fF
C39514 AND2X1_LOC_59/Y AND2X1_LOC_491/a_8_24# 0.01fF
C39515 AND2X1_LOC_131/a_8_24# OR2X1_LOC_598/A 0.01fF
C39516 AND2X1_LOC_458/a_8_24# OR2X1_LOC_371/Y 0.04fF
C39517 OR2X1_LOC_18/Y OR2X1_LOC_628/Y 0.06fF
C39518 AND2X1_LOC_40/Y AND2X1_LOC_47/Y 0.26fF
C39519 AND2X1_LOC_566/a_8_24# AND2X1_LOC_211/a_8_24# 0.23fF
C39520 OR2X1_LOC_18/Y AND2X1_LOC_471/a_8_24# 0.04fF
C39521 OR2X1_LOC_51/Y AND2X1_LOC_624/B 0.00fF
C39522 OR2X1_LOC_599/A AND2X1_LOC_729/B 0.00fF
C39523 OR2X1_LOC_127/Y AND2X1_LOC_128/a_8_24# 0.05fF
C39524 OR2X1_LOC_105/Y AND2X1_LOC_106/a_8_24# 0.11fF
C39525 AND2X1_LOC_717/Y OR2X1_LOC_95/Y 0.00fF
C39526 OR2X1_LOC_496/Y OR2X1_LOC_527/Y 0.04fF
C39527 OR2X1_LOC_175/B OR2X1_LOC_436/Y 0.00fF
C39528 OR2X1_LOC_675/A OR2X1_LOC_269/B 0.00fF
C39529 OR2X1_LOC_87/A OR2X1_LOC_206/A 0.06fF
C39530 OR2X1_LOC_681/Y OR2X1_LOC_52/B 0.04fF
C39531 OR2X1_LOC_45/B OR2X1_LOC_437/A 0.13fF
C39532 OR2X1_LOC_685/A AND2X1_LOC_425/Y 0.00fF
C39533 OR2X1_LOC_185/Y OR2X1_LOC_846/A 0.01fF
C39534 OR2X1_LOC_64/Y OR2X1_LOC_591/a_8_216# 0.05fF
C39535 AND2X1_LOC_843/a_8_24# OR2X1_LOC_417/A 0.01fF
C39536 AND2X1_LOC_64/Y OR2X1_LOC_844/B 0.13fF
C39537 OR2X1_LOC_36/Y OR2X1_LOC_7/a_8_216# 0.01fF
C39538 AND2X1_LOC_217/Y AND2X1_LOC_657/A 0.83fF
C39539 OR2X1_LOC_264/Y OR2X1_LOC_786/Y 0.03fF
C39540 OR2X1_LOC_51/Y OR2X1_LOC_163/Y 0.03fF
C39541 OR2X1_LOC_70/Y OR2X1_LOC_3/Y 0.91fF
C39542 OR2X1_LOC_279/a_8_216# OR2X1_LOC_279/Y 0.01fF
C39543 OR2X1_LOC_416/Y OR2X1_LOC_52/B 0.03fF
C39544 OR2X1_LOC_485/A OR2X1_LOC_615/a_8_216# 0.14fF
C39545 OR2X1_LOC_109/Y AND2X1_LOC_866/A 0.07fF
C39546 AND2X1_LOC_329/a_36_24# AND2X1_LOC_51/Y 0.00fF
C39547 AND2X1_LOC_660/Y AND2X1_LOC_276/Y 0.08fF
C39548 OR2X1_LOC_709/A OR2X1_LOC_515/a_8_216# 0.01fF
C39549 OR2X1_LOC_76/A OR2X1_LOC_733/B 0.03fF
C39550 OR2X1_LOC_485/A AND2X1_LOC_842/B 0.09fF
C39551 OR2X1_LOC_851/a_8_216# OR2X1_LOC_68/B 0.01fF
C39552 OR2X1_LOC_102/a_8_216# OR2X1_LOC_437/A 0.03fF
C39553 OR2X1_LOC_238/a_36_216# OR2X1_LOC_39/A 0.00fF
C39554 OR2X1_LOC_653/A OR2X1_LOC_532/B 0.03fF
C39555 OR2X1_LOC_193/Y AND2X1_LOC_7/Y 0.03fF
C39556 AND2X1_LOC_519/a_8_24# AND2X1_LOC_8/Y 0.01fF
C39557 AND2X1_LOC_845/Y OR2X1_LOC_44/Y 0.13fF
C39558 OR2X1_LOC_673/Y OR2X1_LOC_532/B 0.55fF
C39559 OR2X1_LOC_427/A AND2X1_LOC_808/A 0.08fF
C39560 AND2X1_LOC_141/B AND2X1_LOC_140/a_36_24# 0.00fF
C39561 AND2X1_LOC_64/Y OR2X1_LOC_390/B 0.07fF
C39562 AND2X1_LOC_390/B AND2X1_LOC_856/B 0.03fF
C39563 AND2X1_LOC_858/B AND2X1_LOC_563/Y 0.01fF
C39564 AND2X1_LOC_568/a_8_24# AND2X1_LOC_514/Y 0.02fF
C39565 OR2X1_LOC_52/a_8_216# OR2X1_LOC_52/Y 0.01fF
C39566 OR2X1_LOC_618/Y AND2X1_LOC_9/a_36_24# 0.00fF
C39567 OR2X1_LOC_139/a_8_216# OR2X1_LOC_720/B 0.02fF
C39568 AND2X1_LOC_36/Y OR2X1_LOC_161/B 0.20fF
C39569 AND2X1_LOC_17/Y AND2X1_LOC_7/Y 0.01fF
C39570 OR2X1_LOC_91/Y AND2X1_LOC_851/B 0.07fF
C39571 AND2X1_LOC_40/Y OR2X1_LOC_598/A 0.08fF
C39572 OR2X1_LOC_680/A OR2X1_LOC_674/Y 0.03fF
C39573 AND2X1_LOC_560/B OR2X1_LOC_95/Y 0.01fF
C39574 OR2X1_LOC_70/Y OR2X1_LOC_582/Y 0.01fF
C39575 OR2X1_LOC_97/A OR2X1_LOC_605/Y 0.21fF
C39576 OR2X1_LOC_472/a_8_216# OR2X1_LOC_476/B 0.01fF
C39577 AND2X1_LOC_95/Y OR2X1_LOC_241/B 0.09fF
C39578 OR2X1_LOC_62/A OR2X1_LOC_6/A 0.58fF
C39579 OR2X1_LOC_109/a_8_216# OR2X1_LOC_419/Y 0.10fF
C39580 OR2X1_LOC_613/Y GATE_865 0.03fF
C39581 OR2X1_LOC_494/Y OR2X1_LOC_13/B 0.07fF
C39582 OR2X1_LOC_64/Y AND2X1_LOC_727/A 0.04fF
C39583 VDD OR2X1_LOC_515/Y 0.20fF
C39584 AND2X1_LOC_44/Y OR2X1_LOC_333/a_36_216# 0.02fF
C39585 OR2X1_LOC_680/A AND2X1_LOC_624/B 0.03fF
C39586 D_INPUT_2 OR2X1_LOC_37/a_8_216# 0.03fF
C39587 OR2X1_LOC_643/A OR2X1_LOC_786/Y 0.07fF
C39588 AND2X1_LOC_349/a_8_24# AND2X1_LOC_721/A 0.01fF
C39589 OR2X1_LOC_124/Y OR2X1_LOC_786/Y 0.03fF
C39590 OR2X1_LOC_221/A AND2X1_LOC_47/Y 0.17fF
C39591 AND2X1_LOC_785/A AND2X1_LOC_476/Y 0.04fF
C39592 AND2X1_LOC_242/B AND2X1_LOC_244/A 0.01fF
C39593 OR2X1_LOC_325/B OR2X1_LOC_180/B 0.03fF
C39594 AND2X1_LOC_864/a_8_24# AND2X1_LOC_212/B 0.20fF
C39595 OR2X1_LOC_292/a_8_216# OR2X1_LOC_437/A 0.03fF
C39596 OR2X1_LOC_54/Y OR2X1_LOC_77/a_8_216# 0.14fF
C39597 OR2X1_LOC_488/Y OR2X1_LOC_417/A 0.01fF
C39598 OR2X1_LOC_22/Y AND2X1_LOC_687/B 0.03fF
C39599 AND2X1_LOC_64/Y OR2X1_LOC_840/a_8_216# 0.01fF
C39600 OR2X1_LOC_47/Y AND2X1_LOC_240/Y 0.01fF
C39601 OR2X1_LOC_624/A OR2X1_LOC_228/Y 0.10fF
C39602 OR2X1_LOC_502/A OR2X1_LOC_71/A 0.11fF
C39603 AND2X1_LOC_573/A AND2X1_LOC_563/Y 0.19fF
C39604 OR2X1_LOC_796/B OR2X1_LOC_155/A 0.01fF
C39605 OR2X1_LOC_62/B INPUT_1 0.03fF
C39606 OR2X1_LOC_64/Y OR2X1_LOC_95/Y 9.17fF
C39607 OR2X1_LOC_291/A OR2X1_LOC_619/a_8_216# 0.00fF
C39608 AND2X1_LOC_715/Y OR2X1_LOC_329/a_8_216# 0.02fF
C39609 OR2X1_LOC_691/B OR2X1_LOC_857/A 0.80fF
C39610 AND2X1_LOC_571/B AND2X1_LOC_561/B 0.01fF
C39611 OR2X1_LOC_71/Y D_INPUT_0 0.04fF
C39612 OR2X1_LOC_486/Y AND2X1_LOC_44/Y 0.05fF
C39613 AND2X1_LOC_5/a_36_24# D_INPUT_0 0.00fF
C39614 OR2X1_LOC_447/Y OR2X1_LOC_446/Y 1.48fF
C39615 OR2X1_LOC_611/a_36_216# OR2X1_LOC_62/A 0.11fF
C39616 AND2X1_LOC_8/Y OR2X1_LOC_398/Y 0.01fF
C39617 OR2X1_LOC_6/A OR2X1_LOC_172/Y 0.00fF
C39618 AND2X1_LOC_632/A OR2X1_LOC_95/Y 0.12fF
C39619 AND2X1_LOC_471/a_36_24# OR2X1_LOC_95/Y 0.01fF
C39620 OR2X1_LOC_258/Y AND2X1_LOC_848/A 0.01fF
C39621 AND2X1_LOC_547/a_8_24# AND2X1_LOC_475/Y 0.20fF
C39622 OR2X1_LOC_417/A OR2X1_LOC_95/Y 0.63fF
C39623 OR2X1_LOC_3/Y OR2X1_LOC_70/A 0.12fF
C39624 OR2X1_LOC_316/Y OR2X1_LOC_300/a_36_216# 0.00fF
C39625 OR2X1_LOC_810/A OR2X1_LOC_561/B 0.20fF
C39626 OR2X1_LOC_35/Y OR2X1_LOC_338/A 0.01fF
C39627 OR2X1_LOC_628/Y AND2X1_LOC_620/Y 0.02fF
C39628 OR2X1_LOC_52/B AND2X1_LOC_781/a_36_24# 0.00fF
C39629 OR2X1_LOC_84/B OR2X1_LOC_80/A 0.09fF
C39630 OR2X1_LOC_45/B AND2X1_LOC_715/A 0.02fF
C39631 AND2X1_LOC_476/A AND2X1_LOC_293/a_8_24# 0.02fF
C39632 AND2X1_LOC_810/A AND2X1_LOC_392/A 0.02fF
C39633 D_INPUT_0 D_INPUT_1 0.18fF
C39634 VDD OR2X1_LOC_843/B 0.28fF
C39635 OR2X1_LOC_756/B OR2X1_LOC_174/a_8_216# 0.01fF
C39636 AND2X1_LOC_773/Y OR2X1_LOC_56/A 0.03fF
C39637 OR2X1_LOC_62/A D_INPUT_2 0.09fF
C39638 OR2X1_LOC_97/A AND2X1_LOC_20/a_8_24# 0.01fF
C39639 OR2X1_LOC_40/Y AND2X1_LOC_346/a_8_24# 0.14fF
C39640 D_INPUT_0 OR2X1_LOC_173/a_8_216# 0.01fF
C39641 AND2X1_LOC_41/A AND2X1_LOC_7/B 18.11fF
C39642 OR2X1_LOC_490/a_8_216# OR2X1_LOC_426/B 0.02fF
C39643 VDD OR2X1_LOC_549/A 1.95fF
C39644 AND2X1_LOC_350/a_8_24# OR2X1_LOC_51/Y 0.01fF
C39645 AND2X1_LOC_70/Y OR2X1_LOC_390/A 0.03fF
C39646 OR2X1_LOC_630/Y OR2X1_LOC_161/B 0.01fF
C39647 OR2X1_LOC_287/B OR2X1_LOC_366/Y 0.01fF
C39648 OR2X1_LOC_97/A OR2X1_LOC_634/A 0.00fF
C39649 OR2X1_LOC_40/Y OR2X1_LOC_93/Y 0.02fF
C39650 OR2X1_LOC_49/A OR2X1_LOC_91/A 0.13fF
C39651 OR2X1_LOC_276/a_8_216# OR2X1_LOC_473/A -0.00fF
C39652 OR2X1_LOC_151/A OR2X1_LOC_468/A 0.04fF
C39653 OR2X1_LOC_158/A AND2X1_LOC_709/a_36_24# -0.00fF
C39654 OR2X1_LOC_696/A OR2X1_LOC_432/Y 0.00fF
C39655 OR2X1_LOC_637/A AND2X1_LOC_829/a_8_24# 0.05fF
C39656 AND2X1_LOC_787/A AND2X1_LOC_723/Y 0.32fF
C39657 OR2X1_LOC_65/Y OR2X1_LOC_72/Y 0.07fF
C39658 AND2X1_LOC_141/B AND2X1_LOC_217/a_36_24# 0.01fF
C39659 AND2X1_LOC_658/A AND2X1_LOC_476/Y 0.07fF
C39660 AND2X1_LOC_22/Y AND2X1_LOC_304/a_36_24# 0.00fF
C39661 AND2X1_LOC_91/B OR2X1_LOC_861/a_8_216# 0.02fF
C39662 AND2X1_LOC_50/Y AND2X1_LOC_22/Y 0.02fF
C39663 AND2X1_LOC_217/Y VDD 0.05fF
C39664 OR2X1_LOC_566/A OR2X1_LOC_211/a_8_216# 0.01fF
C39665 AND2X1_LOC_477/Y OR2X1_LOC_59/Y 0.07fF
C39666 OR2X1_LOC_715/B AND2X1_LOC_92/Y 0.10fF
C39667 AND2X1_LOC_594/a_8_24# OR2X1_LOC_756/B 0.01fF
C39668 OR2X1_LOC_543/A OR2X1_LOC_787/B 0.03fF
C39669 OR2X1_LOC_56/A AND2X1_LOC_243/Y 0.02fF
C39670 AND2X1_LOC_626/a_8_24# AND2X1_LOC_92/Y 0.01fF
C39671 AND2X1_LOC_18/Y AND2X1_LOC_616/a_8_24# 0.10fF
C39672 OR2X1_LOC_635/A OR2X1_LOC_161/B 0.46fF
C39673 OR2X1_LOC_743/A AND2X1_LOC_449/a_8_24# 0.01fF
C39674 OR2X1_LOC_177/Y AND2X1_LOC_734/Y 0.03fF
C39675 OR2X1_LOC_604/A OR2X1_LOC_743/a_8_216# 0.01fF
C39676 OR2X1_LOC_593/A OR2X1_LOC_593/B 0.06fF
C39677 OR2X1_LOC_663/A AND2X1_LOC_65/A 0.03fF
C39678 OR2X1_LOC_166/Y AND2X1_LOC_535/Y 0.80fF
C39679 OR2X1_LOC_325/Y VDD -0.00fF
C39680 OR2X1_LOC_188/Y AND2X1_LOC_95/Y 0.05fF
C39681 AND2X1_LOC_191/B OR2X1_LOC_759/A 0.03fF
C39682 AND2X1_LOC_658/B AND2X1_LOC_735/a_8_24# 0.01fF
C39683 AND2X1_LOC_544/Y AND2X1_LOC_807/Y 0.20fF
C39684 AND2X1_LOC_53/Y AND2X1_LOC_31/Y 0.10fF
C39685 OR2X1_LOC_123/a_8_216# AND2X1_LOC_70/Y 0.01fF
C39686 AND2X1_LOC_347/Y OR2X1_LOC_158/A 0.03fF
C39687 OR2X1_LOC_8/Y OR2X1_LOC_104/a_8_216# 0.01fF
C39688 OR2X1_LOC_757/A VDD 0.08fF
C39689 OR2X1_LOC_662/A AND2X1_LOC_7/B 0.03fF
C39690 AND2X1_LOC_18/Y OR2X1_LOC_632/Y 0.14fF
C39691 AND2X1_LOC_22/Y AND2X1_LOC_59/a_36_24# 0.00fF
C39692 AND2X1_LOC_366/A AND2X1_LOC_860/A 0.07fF
C39693 AND2X1_LOC_841/B OR2X1_LOC_16/A 0.03fF
C39694 OR2X1_LOC_113/Y VDD 0.12fF
C39695 OR2X1_LOC_92/Y OR2X1_LOC_421/Y 0.04fF
C39696 AND2X1_LOC_810/A AND2X1_LOC_354/Y 0.01fF
C39697 AND2X1_LOC_40/Y OR2X1_LOC_646/B 0.35fF
C39698 AND2X1_LOC_714/a_36_24# AND2X1_LOC_841/B 0.01fF
C39699 OR2X1_LOC_821/a_36_216# OR2X1_LOC_278/Y 0.00fF
C39700 AND2X1_LOC_682/a_36_24# OR2X1_LOC_161/B 0.00fF
C39701 AND2X1_LOC_575/a_8_24# AND2X1_LOC_575/Y 0.00fF
C39702 AND2X1_LOC_480/a_8_24# AND2X1_LOC_222/Y 0.01fF
C39703 AND2X1_LOC_64/Y OR2X1_LOC_403/B 0.03fF
C39704 OR2X1_LOC_40/Y AND2X1_LOC_737/a_8_24# 0.18fF
C39705 AND2X1_LOC_91/B AND2X1_LOC_399/a_8_24# 0.02fF
C39706 AND2X1_LOC_802/B AND2X1_LOC_388/a_36_24# 0.00fF
C39707 OR2X1_LOC_177/Y OR2X1_LOC_109/a_8_216# 0.01fF
C39708 AND2X1_LOC_195/a_8_24# OR2X1_LOC_18/Y 0.06fF
C39709 AND2X1_LOC_508/A AND2X1_LOC_508/B 0.01fF
C39710 OR2X1_LOC_509/a_8_216# OR2X1_LOC_509/A 0.47fF
C39711 OR2X1_LOC_437/a_8_216# AND2X1_LOC_222/Y 0.01fF
C39712 OR2X1_LOC_329/B OR2X1_LOC_59/Y 0.04fF
C39713 OR2X1_LOC_223/A AND2X1_LOC_31/Y 0.07fF
C39714 INPUT_0 AND2X1_LOC_33/a_36_24# 0.01fF
C39715 VDD OR2X1_LOC_354/A 0.12fF
C39716 AND2X1_LOC_508/A AND2X1_LOC_508/a_8_24# 0.10fF
C39717 OR2X1_LOC_405/A OR2X1_LOC_729/a_8_216# 0.01fF
C39718 OR2X1_LOC_631/B AND2X1_LOC_7/B 0.03fF
C39719 OR2X1_LOC_160/B OR2X1_LOC_175/B 0.00fF
C39720 AND2X1_LOC_93/a_8_24# OR2X1_LOC_633/Y 0.04fF
C39721 OR2X1_LOC_128/A OR2X1_LOC_151/A 0.04fF
C39722 OR2X1_LOC_733/B OR2X1_LOC_722/B 0.21fF
C39723 AND2X1_LOC_303/B OR2X1_LOC_12/Y 0.00fF
C39724 AND2X1_LOC_449/Y AND2X1_LOC_605/a_8_24# 0.01fF
C39725 OR2X1_LOC_648/A OR2X1_LOC_775/a_8_216# -0.02fF
C39726 AND2X1_LOC_303/A AND2X1_LOC_339/B 0.03fF
C39727 AND2X1_LOC_486/Y OR2X1_LOC_51/Y 0.04fF
C39728 AND2X1_LOC_56/B OR2X1_LOC_35/A 0.02fF
C39729 OR2X1_LOC_544/A OR2X1_LOC_544/B 0.07fF
C39730 AND2X1_LOC_95/Y OR2X1_LOC_325/B 0.07fF
C39731 OR2X1_LOC_676/Y AND2X1_LOC_16/a_8_24# 0.03fF
C39732 OR2X1_LOC_441/Y AND2X1_LOC_148/a_8_24# 0.07fF
C39733 OR2X1_LOC_51/Y AND2X1_LOC_840/a_36_24# 0.00fF
C39734 OR2X1_LOC_532/B OR2X1_LOC_723/B 0.03fF
C39735 OR2X1_LOC_6/B AND2X1_LOC_43/B 0.07fF
C39736 AND2X1_LOC_535/Y AND2X1_LOC_365/A 0.02fF
C39737 AND2X1_LOC_218/a_36_24# OR2X1_LOC_18/Y 0.01fF
C39738 OR2X1_LOC_74/Y OR2X1_LOC_59/Y 0.01fF
C39739 OR2X1_LOC_543/a_8_216# OR2X1_LOC_552/A 0.01fF
C39740 AND2X1_LOC_508/B OR2X1_LOC_18/Y 0.01fF
C39741 OR2X1_LOC_312/Y AND2X1_LOC_802/Y 0.24fF
C39742 OR2X1_LOC_663/a_8_216# OR2X1_LOC_849/A 0.01fF
C39743 OR2X1_LOC_771/a_8_216# OR2X1_LOC_80/A 0.01fF
C39744 OR2X1_LOC_774/B OR2X1_LOC_68/B 0.10fF
C39745 OR2X1_LOC_377/A OR2X1_LOC_676/Y 0.01fF
C39746 OR2X1_LOC_79/A OR2X1_LOC_79/a_8_216# 0.47fF
C39747 OR2X1_LOC_102/a_8_216# OR2X1_LOC_753/A 0.01fF
C39748 OR2X1_LOC_441/Y OR2X1_LOC_746/a_8_216# 0.06fF
C39749 AND2X1_LOC_712/a_8_24# OR2X1_LOC_743/A 0.01fF
C39750 AND2X1_LOC_160/Y OR2X1_LOC_619/Y 0.02fF
C39751 GATE_811 AND2X1_LOC_740/a_36_24# 0.00fF
C39752 OR2X1_LOC_424/a_8_216# AND2X1_LOC_447/Y 0.14fF
C39753 OR2X1_LOC_168/a_8_216# OR2X1_LOC_78/A 0.05fF
C39754 AND2X1_LOC_719/Y AND2X1_LOC_859/Y 0.06fF
C39755 OR2X1_LOC_151/A OR2X1_LOC_449/B 0.07fF
C39756 AND2X1_LOC_593/a_8_24# OR2X1_LOC_599/A 0.04fF
C39757 OR2X1_LOC_97/A OR2X1_LOC_602/a_8_216# 0.01fF
C39758 AND2X1_LOC_91/B OR2X1_LOC_401/B 0.18fF
C39759 AND2X1_LOC_444/a_36_24# AND2X1_LOC_804/Y 0.00fF
C39760 AND2X1_LOC_56/B OR2X1_LOC_552/B 0.05fF
C39761 AND2X1_LOC_40/Y OR2X1_LOC_828/a_8_216# 0.01fF
C39762 OR2X1_LOC_482/a_8_216# OR2X1_LOC_665/Y 0.00fF
C39763 OR2X1_LOC_40/Y OR2X1_LOC_262/a_8_216# 0.03fF
C39764 OR2X1_LOC_632/A OR2X1_LOC_632/a_8_216# 0.39fF
C39765 AND2X1_LOC_535/Y OR2X1_LOC_43/A 0.01fF
C39766 AND2X1_LOC_122/a_36_24# AND2X1_LOC_44/Y 0.00fF
C39767 OR2X1_LOC_215/Y AND2X1_LOC_92/Y 0.02fF
C39768 OR2X1_LOC_486/a_8_216# AND2X1_LOC_44/Y 0.15fF
C39769 OR2X1_LOC_567/a_8_216# OR2X1_LOC_568/A 0.13fF
C39770 AND2X1_LOC_113/Y OR2X1_LOC_59/Y 0.00fF
C39771 OR2X1_LOC_565/A OR2X1_LOC_564/A 0.68fF
C39772 AND2X1_LOC_95/Y AND2X1_LOC_189/a_8_24# 0.02fF
C39773 VDD OR2X1_LOC_498/a_8_216# 0.21fF
C39774 OR2X1_LOC_757/A OR2X1_LOC_616/Y 0.01fF
C39775 OR2X1_LOC_8/Y OR2X1_LOC_6/A 2.38fF
C39776 VDD AND2X1_LOC_359/B 0.02fF
C39777 AND2X1_LOC_580/B OR2X1_LOC_600/A 0.02fF
C39778 OR2X1_LOC_51/Y AND2X1_LOC_834/a_8_24# 0.02fF
C39779 OR2X1_LOC_214/B AND2X1_LOC_41/Y 0.82fF
C39780 OR2X1_LOC_612/a_8_216# OR2X1_LOC_612/B 0.05fF
C39781 OR2X1_LOC_500/A OR2X1_LOC_632/Y 0.01fF
C39782 OR2X1_LOC_421/A OR2X1_LOC_682/Y 0.12fF
C39783 AND2X1_LOC_191/Y AND2X1_LOC_477/Y 0.26fF
C39784 OR2X1_LOC_18/Y AND2X1_LOC_850/A 0.00fF
C39785 OR2X1_LOC_13/B OR2X1_LOC_311/a_8_216# 0.01fF
C39786 OR2X1_LOC_335/A OR2X1_LOC_532/B 0.00fF
C39787 OR2X1_LOC_71/A OR2X1_LOC_398/a_8_216# 0.01fF
C39788 AND2X1_LOC_95/Y OR2X1_LOC_285/a_8_216# 0.01fF
C39789 OR2X1_LOC_324/a_8_216# OR2X1_LOC_324/A 0.47fF
C39790 OR2X1_LOC_235/B OR2X1_LOC_668/Y 0.01fF
C39791 OR2X1_LOC_92/Y OR2X1_LOC_278/Y 0.08fF
C39792 OR2X1_LOC_51/Y OR2X1_LOC_248/Y 0.04fF
C39793 VDD OR2X1_LOC_423/a_8_216# 0.00fF
C39794 AND2X1_LOC_357/a_8_24# AND2X1_LOC_364/A 0.01fF
C39795 AND2X1_LOC_711/Y AND2X1_LOC_477/Y 0.07fF
C39796 VDD OR2X1_LOC_711/A 0.18fF
C39797 OR2X1_LOC_479/Y OR2X1_LOC_787/a_8_216# 0.04fF
C39798 OR2X1_LOC_51/Y OR2X1_LOC_6/a_8_216# 0.01fF
C39799 OR2X1_LOC_92/Y AND2X1_LOC_662/B 0.41fF
C39800 AND2X1_LOC_40/Y OR2X1_LOC_506/A 0.03fF
C39801 OR2X1_LOC_19/B OR2X1_LOC_414/Y 0.05fF
C39802 OR2X1_LOC_821/Y OR2X1_LOC_64/Y 0.04fF
C39803 OR2X1_LOC_70/Y AND2X1_LOC_477/Y 0.42fF
C39804 OR2X1_LOC_600/Y AND2X1_LOC_602/a_8_24# 0.23fF
C39805 OR2X1_LOC_703/B OR2X1_LOC_756/B 0.02fF
C39806 AND2X1_LOC_707/Y AND2X1_LOC_687/Y 0.82fF
C39807 AND2X1_LOC_347/B AND2X1_LOC_347/a_36_24# 0.01fF
C39808 OR2X1_LOC_564/A OR2X1_LOC_190/Y 0.02fF
C39809 OR2X1_LOC_865/Y OR2X1_LOC_391/A 0.03fF
C39810 OR2X1_LOC_744/A OR2X1_LOC_283/Y 1.46fF
C39811 OR2X1_LOC_7/A AND2X1_LOC_447/Y 0.01fF
C39812 AND2X1_LOC_527/a_8_24# OR2X1_LOC_620/Y 0.02fF
C39813 OR2X1_LOC_235/B OR2X1_LOC_36/Y 0.02fF
C39814 OR2X1_LOC_532/B OR2X1_LOC_720/Y 0.01fF
C39815 OR2X1_LOC_91/A AND2X1_LOC_661/A 0.01fF
C39816 OR2X1_LOC_185/Y AND2X1_LOC_311/a_36_24# 0.01fF
C39817 OR2X1_LOC_666/Y OR2X1_LOC_51/Y 0.22fF
C39818 OR2X1_LOC_637/A OR2X1_LOC_828/B 0.00fF
C39819 VDD AND2X1_LOC_639/a_8_24# -0.00fF
C39820 OR2X1_LOC_756/B OR2X1_LOC_87/A 0.03fF
C39821 OR2X1_LOC_269/B AND2X1_LOC_437/a_36_24# 0.01fF
C39822 AND2X1_LOC_541/a_8_24# OR2X1_LOC_95/Y -0.01fF
C39823 AND2X1_LOC_729/Y OR2X1_LOC_485/a_8_216# 0.01fF
C39824 OR2X1_LOC_151/A OR2X1_LOC_121/B 0.10fF
C39825 OR2X1_LOC_40/Y AND2X1_LOC_729/B 0.03fF
C39826 OR2X1_LOC_97/A OR2X1_LOC_439/a_8_216# 0.01fF
C39827 OR2X1_LOC_532/B AND2X1_LOC_277/a_8_24# 0.01fF
C39828 AND2X1_LOC_658/B AND2X1_LOC_631/Y 0.01fF
C39829 AND2X1_LOC_711/A OR2X1_LOC_481/A 0.08fF
C39830 AND2X1_LOC_259/Y OR2X1_LOC_91/A 0.02fF
C39831 OR2X1_LOC_427/A OR2X1_LOC_39/A 0.24fF
C39832 OR2X1_LOC_516/B OR2X1_LOC_26/Y 0.10fF
C39833 AND2X1_LOC_322/a_8_24# OR2X1_LOC_121/B 0.01fF
C39834 AND2X1_LOC_95/Y OR2X1_LOC_405/Y 0.01fF
C39835 AND2X1_LOC_512/a_8_24# AND2X1_LOC_512/Y 0.01fF
C39836 AND2X1_LOC_550/A AND2X1_LOC_807/Y 0.02fF
C39837 OR2X1_LOC_600/A OR2X1_LOC_295/a_8_216# 0.01fF
C39838 AND2X1_LOC_59/Y OR2X1_LOC_185/A 0.28fF
C39839 OR2X1_LOC_780/a_8_216# OR2X1_LOC_161/B 0.02fF
C39840 AND2X1_LOC_339/Y OR2X1_LOC_75/Y 0.81fF
C39841 OR2X1_LOC_702/A OR2X1_LOC_538/A 0.02fF
C39842 AND2X1_LOC_95/Y OR2X1_LOC_652/a_36_216# 0.00fF
C39843 OR2X1_LOC_684/a_8_216# OR2X1_LOC_684/Y 0.04fF
C39844 OR2X1_LOC_778/A OR2X1_LOC_778/B 0.01fF
C39845 OR2X1_LOC_70/Y OR2X1_LOC_329/B 0.15fF
C39846 INPUT_0 AND2X1_LOC_136/a_8_24# 0.04fF
C39847 AND2X1_LOC_41/A OR2X1_LOC_296/Y 0.01fF
C39848 OR2X1_LOC_806/a_36_216# OR2X1_LOC_807/A 0.00fF
C39849 OR2X1_LOC_814/A OR2X1_LOC_641/A 2.48fF
C39850 OR2X1_LOC_7/Y AND2X1_LOC_194/Y 0.00fF
C39851 D_INPUT_7 D_INPUT_5 0.08fF
C39852 AND2X1_LOC_64/Y OR2X1_LOC_493/Y 0.01fF
C39853 AND2X1_LOC_580/A AND2X1_LOC_621/Y 0.07fF
C39854 AND2X1_LOC_703/Y AND2X1_LOC_648/B 0.00fF
C39855 OR2X1_LOC_131/A OR2X1_LOC_71/Y 0.00fF
C39856 OR2X1_LOC_756/B AND2X1_LOC_815/a_8_24# 0.01fF
C39857 OR2X1_LOC_377/A OR2X1_LOC_462/B 0.94fF
C39858 OR2X1_LOC_313/a_36_216# OR2X1_LOC_314/Y 0.00fF
C39859 OR2X1_LOC_585/A OR2X1_LOC_586/Y 0.09fF
C39860 AND2X1_LOC_70/Y OR2X1_LOC_750/A 0.00fF
C39861 OR2X1_LOC_271/Y AND2X1_LOC_662/B 0.00fF
C39862 OR2X1_LOC_660/B OR2X1_LOC_87/A 0.03fF
C39863 OR2X1_LOC_479/Y OR2X1_LOC_808/B 0.10fF
C39864 AND2X1_LOC_129/a_8_24# OR2X1_LOC_87/Y 0.02fF
C39865 OR2X1_LOC_600/a_8_216# AND2X1_LOC_477/A 0.01fF
C39866 AND2X1_LOC_339/B AND2X1_LOC_655/a_8_24# 0.01fF
C39867 AND2X1_LOC_332/a_8_24# AND2X1_LOC_660/A 0.20fF
C39868 OR2X1_LOC_462/B AND2X1_LOC_824/B 0.14fF
C39869 OR2X1_LOC_499/B AND2X1_LOC_496/a_36_24# 0.00fF
C39870 OR2X1_LOC_250/a_8_216# OR2X1_LOC_106/A 0.48fF
C39871 OR2X1_LOC_329/B AND2X1_LOC_514/Y 0.46fF
C39872 OR2X1_LOC_680/A AND2X1_LOC_834/a_8_24# 0.11fF
C39873 AND2X1_LOC_729/Y OR2X1_LOC_44/Y 0.07fF
C39874 OR2X1_LOC_631/B OR2X1_LOC_805/A 0.07fF
C39875 OR2X1_LOC_622/B OR2X1_LOC_80/A 0.01fF
C39876 OR2X1_LOC_673/B D_INPUT_1 0.00fF
C39877 OR2X1_LOC_429/Y OR2X1_LOC_427/A 0.02fF
C39878 OR2X1_LOC_426/B D_INPUT_0 0.18fF
C39879 OR2X1_LOC_2/Y OR2X1_LOC_17/Y 0.22fF
C39880 AND2X1_LOC_519/a_8_24# AND2X1_LOC_92/Y 0.01fF
C39881 AND2X1_LOC_319/A OR2X1_LOC_36/Y 0.03fF
C39882 OR2X1_LOC_109/Y OR2X1_LOC_7/A 0.03fF
C39883 OR2X1_LOC_632/A AND2X1_LOC_3/Y 0.02fF
C39884 AND2X1_LOC_554/B AND2X1_LOC_99/A 0.02fF
C39885 AND2X1_LOC_56/B OR2X1_LOC_793/A 0.03fF
C39886 OR2X1_LOC_246/Y OR2X1_LOC_43/A 0.07fF
C39887 OR2X1_LOC_641/B OR2X1_LOC_227/A 0.01fF
C39888 OR2X1_LOC_7/A AND2X1_LOC_448/Y 0.02fF
C39889 AND2X1_LOC_388/Y OR2X1_LOC_47/Y 0.03fF
C39890 OR2X1_LOC_317/B OR2X1_LOC_308/Y 0.06fF
C39891 AND2X1_LOC_12/Y D_INPUT_7 0.24fF
C39892 OR2X1_LOC_629/A OR2X1_LOC_161/A 0.04fF
C39893 OR2X1_LOC_209/A OR2X1_LOC_550/B 0.88fF
C39894 OR2X1_LOC_204/Y OR2X1_LOC_124/Y 0.24fF
C39895 AND2X1_LOC_784/A OR2X1_LOC_44/Y 0.07fF
C39896 AND2X1_LOC_477/A AND2X1_LOC_477/a_8_24# 0.01fF
C39897 OR2X1_LOC_8/Y D_INPUT_2 0.01fF
C39898 OR2X1_LOC_6/A OR2X1_LOC_52/B 1.10fF
C39899 OR2X1_LOC_672/Y OR2X1_LOC_6/A 0.00fF
C39900 OR2X1_LOC_19/B OR2X1_LOC_92/Y 0.13fF
C39901 AND2X1_LOC_831/Y AND2X1_LOC_219/Y 0.00fF
C39902 OR2X1_LOC_3/Y AND2X1_LOC_124/a_8_24# 0.04fF
C39903 AND2X1_LOC_557/Y OR2X1_LOC_89/A 0.01fF
C39904 OR2X1_LOC_440/A OR2X1_LOC_78/A 0.01fF
C39905 OR2X1_LOC_850/B OR2X1_LOC_287/a_8_216# 0.18fF
C39906 OR2X1_LOC_107/Y AND2X1_LOC_227/Y 0.02fF
C39907 AND2X1_LOC_769/a_8_24# OR2X1_LOC_44/Y 0.01fF
C39908 OR2X1_LOC_92/Y AND2X1_LOC_800/a_8_24# 0.02fF
C39909 AND2X1_LOC_741/Y AND2X1_LOC_223/a_36_24# 0.00fF
C39910 OR2X1_LOC_631/B OR2X1_LOC_296/Y 0.01fF
C39911 AND2X1_LOC_12/Y OR2X1_LOC_476/B 0.07fF
C39912 OR2X1_LOC_481/Y OR2X1_LOC_44/Y 0.31fF
C39913 OR2X1_LOC_19/B OR2X1_LOC_65/B 0.03fF
C39914 AND2X1_LOC_328/a_36_24# AND2X1_LOC_7/Y 0.00fF
C39915 OR2X1_LOC_3/Y OR2X1_LOC_240/A 0.07fF
C39916 OR2X1_LOC_654/A AND2X1_LOC_822/a_36_24# 0.01fF
C39917 OR2X1_LOC_742/B OR2X1_LOC_550/a_36_216# 0.02fF
C39918 OR2X1_LOC_759/A AND2X1_LOC_848/A 0.02fF
C39919 AND2X1_LOC_95/Y D_INPUT_0 0.11fF
C39920 OR2X1_LOC_694/a_36_216# AND2X1_LOC_687/B 0.00fF
C39921 OR2X1_LOC_802/a_36_216# OR2X1_LOC_436/Y 0.00fF
C39922 AND2X1_LOC_801/B AND2X1_LOC_809/A 0.01fF
C39923 AND2X1_LOC_12/Y OR2X1_LOC_644/a_8_216# 0.01fF
C39924 AND2X1_LOC_792/Y AND2X1_LOC_663/A 0.10fF
C39925 OR2X1_LOC_757/A AND2X1_LOC_624/B 0.02fF
C39926 AND2X1_LOC_18/Y OR2X1_LOC_358/A 0.08fF
C39927 OR2X1_LOC_633/Y D_INPUT_0 0.01fF
C39928 OR2X1_LOC_427/A OR2X1_LOC_428/a_8_216# 0.01fF
C39929 OR2X1_LOC_31/Y AND2X1_LOC_520/Y 0.04fF
C39930 AND2X1_LOC_489/Y AND2X1_LOC_557/a_8_24# 0.04fF
C39931 AND2X1_LOC_155/Y OR2X1_LOC_743/A 0.01fF
C39932 AND2X1_LOC_40/Y OR2X1_LOC_227/Y 0.00fF
C39933 OR2X1_LOC_147/a_8_216# AND2X1_LOC_51/Y 0.01fF
C39934 AND2X1_LOC_31/Y OR2X1_LOC_777/a_8_216# 0.01fF
C39935 OR2X1_LOC_87/A OR2X1_LOC_227/a_8_216# 0.06fF
C39936 OR2X1_LOC_641/A OR2X1_LOC_341/a_8_216# 0.02fF
C39937 AND2X1_LOC_729/B OR2X1_LOC_7/A 0.19fF
C39938 OR2X1_LOC_599/A OR2X1_LOC_46/A 0.02fF
C39939 AND2X1_LOC_140/a_36_24# OR2X1_LOC_89/A 0.00fF
C39940 AND2X1_LOC_802/Y OR2X1_LOC_13/B 0.04fF
C39941 AND2X1_LOC_175/B OR2X1_LOC_31/Y 0.04fF
C39942 AND2X1_LOC_40/Y D_INPUT_1 0.06fF
C39943 OR2X1_LOC_177/Y OR2X1_LOC_164/a_36_216# 0.00fF
C39944 AND2X1_LOC_10/a_8_24# AND2X1_LOC_42/B 0.01fF
C39945 AND2X1_LOC_47/Y AND2X1_LOC_43/B 0.19fF
C39946 D_INPUT_7 AND2X1_LOC_21/a_8_24# 0.01fF
C39947 AND2X1_LOC_132/a_36_24# AND2X1_LOC_47/Y 0.00fF
C39948 AND2X1_LOC_642/a_8_24# AND2X1_LOC_660/A 0.03fF
C39949 AND2X1_LOC_839/A OR2X1_LOC_85/A 0.01fF
C39950 OR2X1_LOC_641/Y OR2X1_LOC_68/B 0.03fF
C39951 OR2X1_LOC_158/A OR2X1_LOC_437/A 0.40fF
C39952 OR2X1_LOC_161/B OR2X1_LOC_374/a_8_216# 0.01fF
C39953 OR2X1_LOC_810/a_8_216# D_INPUT_1 0.01fF
C39954 OR2X1_LOC_698/Y AND2X1_LOC_848/A 0.05fF
C39955 AND2X1_LOC_796/Y AND2X1_LOC_624/A 0.03fF
C39956 OR2X1_LOC_707/B OR2X1_LOC_155/A 0.00fF
C39957 AND2X1_LOC_44/Y OR2X1_LOC_308/Y 0.11fF
C39958 INPUT_7 D_INPUT_6 0.25fF
C39959 OR2X1_LOC_22/Y AND2X1_LOC_640/Y 0.00fF
C39960 AND2X1_LOC_293/a_8_24# OR2X1_LOC_690/A 0.18fF
C39961 OR2X1_LOC_62/A OR2X1_LOC_44/Y 0.00fF
C39962 OR2X1_LOC_743/A D_INPUT_0 0.07fF
C39963 OR2X1_LOC_848/A D_INPUT_1 0.03fF
C39964 OR2X1_LOC_502/A AND2X1_LOC_31/Y 0.36fF
C39965 AND2X1_LOC_165/a_8_24# AND2X1_LOC_51/Y 0.09fF
C39966 OR2X1_LOC_450/A OR2X1_LOC_712/B 0.03fF
C39967 AND2X1_LOC_56/B AND2X1_LOC_271/a_8_24# 0.01fF
C39968 AND2X1_LOC_564/B AND2X1_LOC_721/Y 0.05fF
C39969 OR2X1_LOC_859/B D_INPUT_1 0.00fF
C39970 OR2X1_LOC_22/Y OR2X1_LOC_416/Y 0.03fF
C39971 OR2X1_LOC_165/a_36_216# AND2X1_LOC_222/Y 0.00fF
C39972 AND2X1_LOC_43/B OR2X1_LOC_598/A 0.11fF
C39973 AND2X1_LOC_711/A AND2X1_LOC_789/Y 0.02fF
C39974 OR2X1_LOC_605/A OR2X1_LOC_440/A 0.07fF
C39975 OR2X1_LOC_545/B AND2X1_LOC_442/a_8_24# 0.20fF
C39976 AND2X1_LOC_191/Y GATE_662 0.03fF
C39977 AND2X1_LOC_191/Y GATE_811 0.03fF
C39978 OR2X1_LOC_154/A OR2X1_LOC_590/a_8_216# 0.01fF
C39979 AND2X1_LOC_98/Y OR2X1_LOC_437/A 0.02fF
C39980 OR2X1_LOC_600/A AND2X1_LOC_793/a_36_24# 0.00fF
C39981 AND2X1_LOC_711/Y GATE_662 0.04fF
C39982 OR2X1_LOC_415/a_8_216# D_INPUT_0 0.01fF
C39983 OR2X1_LOC_626/a_8_216# AND2X1_LOC_624/B 0.01fF
C39984 OR2X1_LOC_3/Y OR2X1_LOC_47/Y 0.62fF
C39985 AND2X1_LOC_31/Y AND2X1_LOC_230/a_8_24# 0.01fF
C39986 OR2X1_LOC_246/A D_INPUT_0 1.93fF
C39987 OR2X1_LOC_437/a_8_216# OR2X1_LOC_74/A 0.02fF
C39988 OR2X1_LOC_155/A OR2X1_LOC_446/A 0.05fF
C39989 AND2X1_LOC_568/a_8_24# OR2X1_LOC_47/Y 0.01fF
C39990 OR2X1_LOC_474/Y OR2X1_LOC_140/Y 0.11fF
C39991 OR2X1_LOC_45/a_8_216# OR2X1_LOC_172/Y 0.44fF
C39992 OR2X1_LOC_53/Y AND2X1_LOC_199/A 0.01fF
C39993 OR2X1_LOC_285/Y OR2X1_LOC_286/B 0.06fF
C39994 OR2X1_LOC_696/A AND2X1_LOC_537/a_8_24# 0.03fF
C39995 OR2X1_LOC_136/a_8_216# AND2X1_LOC_566/B 0.01fF
C39996 AND2X1_LOC_524/a_8_24# AND2X1_LOC_7/B 0.03fF
C39997 OR2X1_LOC_630/B AND2X1_LOC_36/Y 0.01fF
C39998 AND2X1_LOC_711/a_36_24# AND2X1_LOC_789/Y 0.00fF
C39999 OR2X1_LOC_473/A AND2X1_LOC_51/Y 0.43fF
C40000 OR2X1_LOC_756/B OR2X1_LOC_579/A 0.21fF
C40001 OR2X1_LOC_468/Y OR2X1_LOC_566/a_8_216# 0.01fF
C40002 INPUT_1 OR2X1_LOC_75/a_8_216# 0.01fF
C40003 AND2X1_LOC_49/a_8_24# OR2X1_LOC_80/A 0.05fF
C40004 OR2X1_LOC_44/Y OR2X1_LOC_172/Y 0.33fF
C40005 AND2X1_LOC_147/a_8_24# OR2X1_LOC_142/Y -0.00fF
C40006 OR2X1_LOC_95/Y OR2X1_LOC_226/a_8_216# -0.00fF
C40007 OR2X1_LOC_212/A OR2X1_LOC_303/B 0.43fF
C40008 OR2X1_LOC_589/A OR2X1_LOC_16/A 0.06fF
C40009 OR2X1_LOC_596/A OR2X1_LOC_138/A 0.01fF
C40010 OR2X1_LOC_426/A D_INPUT_6 0.21fF
C40011 AND2X1_LOC_40/Y OR2X1_LOC_180/B 0.07fF
C40012 AND2X1_LOC_564/B OR2X1_LOC_496/a_36_216# 0.01fF
C40013 OR2X1_LOC_687/Y OR2X1_LOC_446/B 0.03fF
C40014 AND2X1_LOC_95/Y OR2X1_LOC_339/A 0.03fF
C40015 OR2X1_LOC_756/B OR2X1_LOC_390/B 0.01fF
C40016 AND2X1_LOC_227/Y AND2X1_LOC_866/A 0.03fF
C40017 OR2X1_LOC_494/Y OR2X1_LOC_428/A 0.75fF
C40018 OR2X1_LOC_648/A AND2X1_LOC_7/B 0.07fF
C40019 OR2X1_LOC_99/B OR2X1_LOC_99/A 0.27fF
C40020 AND2X1_LOC_363/Y OR2X1_LOC_428/A 0.03fF
C40021 AND2X1_LOC_3/Y AND2X1_LOC_427/a_36_24# 0.00fF
C40022 AND2X1_LOC_610/a_8_24# OR2X1_LOC_71/A 0.03fF
C40023 OR2X1_LOC_382/Y AND2X1_LOC_555/Y 0.02fF
C40024 AND2X1_LOC_303/A OR2X1_LOC_300/Y 0.00fF
C40025 OR2X1_LOC_451/A OR2X1_LOC_451/B 0.05fF
C40026 OR2X1_LOC_816/A AND2X1_LOC_663/A 0.09fF
C40027 OR2X1_LOC_215/A OR2X1_LOC_641/B 0.08fF
C40028 OR2X1_LOC_89/A AND2X1_LOC_217/a_36_24# 0.00fF
C40029 AND2X1_LOC_364/a_36_24# OR2X1_LOC_426/B 0.05fF
C40030 AND2X1_LOC_719/Y AND2X1_LOC_722/a_8_24# 0.25fF
C40031 OR2X1_LOC_323/A OR2X1_LOC_92/Y 0.03fF
C40032 AND2X1_LOC_51/Y OR2X1_LOC_228/Y 0.07fF
C40033 OR2X1_LOC_45/B AND2X1_LOC_222/a_8_24# 0.01fF
C40034 OR2X1_LOC_56/A OR2X1_LOC_12/Y 1.13fF
C40035 D_INPUT_3 OR2X1_LOC_619/a_8_216# 0.01fF
C40036 INPUT_4 D_INPUT_6 0.97fF
C40037 OR2X1_LOC_166/Y OR2X1_LOC_16/A 0.02fF
C40038 OR2X1_LOC_158/A AND2X1_LOC_715/A 0.06fF
C40039 OR2X1_LOC_6/B AND2X1_LOC_625/a_36_24# 0.00fF
C40040 AND2X1_LOC_794/B AND2X1_LOC_436/Y 0.05fF
C40041 AND2X1_LOC_658/B AND2X1_LOC_477/Y 0.07fF
C40042 OR2X1_LOC_56/Y OR2X1_LOC_16/Y 0.15fF
C40043 OR2X1_LOC_131/A OR2X1_LOC_426/B 0.42fF
C40044 AND2X1_LOC_167/a_8_24# OR2X1_LOC_161/B 0.01fF
C40045 AND2X1_LOC_22/Y AND2X1_LOC_615/a_8_24# 0.04fF
C40046 OR2X1_LOC_485/A OR2X1_LOC_536/a_36_216# 0.01fF
C40047 AND2X1_LOC_48/A AND2X1_LOC_31/Y 0.14fF
C40048 AND2X1_LOC_714/B OR2X1_LOC_91/A 0.03fF
C40049 AND2X1_LOC_564/A OR2X1_LOC_427/A 0.03fF
C40050 AND2X1_LOC_638/Y OR2X1_LOC_12/Y 0.03fF
C40051 AND2X1_LOC_51/A D_INPUT_6 0.18fF
C40052 OR2X1_LOC_186/Y OR2X1_LOC_840/A 0.05fF
C40053 VDD AND2X1_LOC_436/Y 0.01fF
C40054 OR2X1_LOC_190/A OR2X1_LOC_741/Y 0.00fF
C40055 OR2X1_LOC_865/A OR2X1_LOC_812/B 0.71fF
C40056 AND2X1_LOC_139/A AND2X1_LOC_216/A 0.02fF
C40057 OR2X1_LOC_426/B AND2X1_LOC_326/B 0.02fF
C40058 OR2X1_LOC_405/a_8_216# AND2X1_LOC_7/B 0.01fF
C40059 OR2X1_LOC_170/A OR2X1_LOC_168/Y 0.06fF
C40060 VDD OR2X1_LOC_360/a_8_216# 0.00fF
C40061 AND2X1_LOC_44/a_8_24# INPUT_6 0.01fF
C40062 AND2X1_LOC_159/a_36_24# OR2X1_LOC_844/B 0.00fF
C40063 OR2X1_LOC_317/a_8_216# OR2X1_LOC_151/A 0.04fF
C40064 OR2X1_LOC_539/A OR2X1_LOC_390/A 0.00fF
C40065 OR2X1_LOC_648/B AND2X1_LOC_41/A 0.10fF
C40066 OR2X1_LOC_468/Y OR2X1_LOC_170/a_8_216# 0.01fF
C40067 OR2X1_LOC_193/A AND2X1_LOC_41/Y 0.00fF
C40068 OR2X1_LOC_323/A AND2X1_LOC_464/a_36_24# 0.00fF
C40069 OR2X1_LOC_203/a_8_216# AND2X1_LOC_7/B 0.01fF
C40070 OR2X1_LOC_676/Y OR2X1_LOC_78/B 0.57fF
C40071 OR2X1_LOC_147/B OR2X1_LOC_294/Y 0.03fF
C40072 OR2X1_LOC_427/A AND2X1_LOC_727/B 0.03fF
C40073 AND2X1_LOC_702/a_8_24# OR2X1_LOC_428/A 0.11fF
C40074 OR2X1_LOC_121/B OR2X1_LOC_714/A 0.09fF
C40075 AND2X1_LOC_194/a_8_24# AND2X1_LOC_194/Y 0.02fF
C40076 AND2X1_LOC_70/a_8_24# AND2X1_LOC_70/Y 0.01fF
C40077 AND2X1_LOC_398/a_8_24# OR2X1_LOC_16/A 0.09fF
C40078 OR2X1_LOC_323/A OR2X1_LOC_271/Y 0.01fF
C40079 OR2X1_LOC_235/B OR2X1_LOC_66/A 0.09fF
C40080 OR2X1_LOC_281/a_8_216# OR2X1_LOC_281/Y 0.01fF
C40081 OR2X1_LOC_218/Y OR2X1_LOC_68/B 0.02fF
C40082 OR2X1_LOC_121/B OR2X1_LOC_716/a_8_216# 0.00fF
C40083 AND2X1_LOC_748/a_8_24# OR2X1_LOC_161/B 0.02fF
C40084 AND2X1_LOC_95/Y AND2X1_LOC_438/a_8_24# 0.03fF
C40085 AND2X1_LOC_764/a_8_24# INPUT_0 0.01fF
C40086 OR2X1_LOC_856/B OR2X1_LOC_151/A 0.18fF
C40087 OR2X1_LOC_318/a_8_216# OR2X1_LOC_185/A 0.01fF
C40088 AND2X1_LOC_508/A AND2X1_LOC_657/Y 0.49fF
C40089 AND2X1_LOC_47/Y OR2X1_LOC_367/B 0.15fF
C40090 OR2X1_LOC_482/Y AND2X1_LOC_833/a_36_24# 0.07fF
C40091 OR2X1_LOC_744/A OR2X1_LOC_26/a_8_216# 0.01fF
C40092 VDD AND2X1_LOC_344/a_8_24# 0.00fF
C40093 OR2X1_LOC_377/A AND2X1_LOC_83/a_8_24# 0.04fF
C40094 INPUT_1 OR2X1_LOC_13/B 0.07fF
C40095 AND2X1_LOC_362/B AND2X1_LOC_99/A 0.04fF
C40096 OR2X1_LOC_812/B D_GATE_811 0.03fF
C40097 OR2X1_LOC_619/Y OR2X1_LOC_421/Y 0.03fF
C40098 OR2X1_LOC_3/Y OR2X1_LOC_397/a_8_216# 0.01fF
C40099 AND2X1_LOC_86/Y OR2X1_LOC_786/A 0.06fF
C40100 AND2X1_LOC_861/B AND2X1_LOC_858/B 0.01fF
C40101 AND2X1_LOC_160/a_8_24# OR2X1_LOC_744/A 0.09fF
C40102 OR2X1_LOC_364/A AND2X1_LOC_433/a_8_24# 0.01fF
C40103 AND2X1_LOC_95/Y OR2X1_LOC_598/Y 0.03fF
C40104 AND2X1_LOC_562/B OR2X1_LOC_744/A 0.39fF
C40105 AND2X1_LOC_539/Y OR2X1_LOC_743/A 0.04fF
C40106 OR2X1_LOC_45/B AND2X1_LOC_778/a_8_24# 0.01fF
C40107 OR2X1_LOC_9/a_8_216# OR2X1_LOC_6/A 0.01fF
C40108 AND2X1_LOC_95/Y OR2X1_LOC_356/a_8_216# 0.01fF
C40109 OR2X1_LOC_600/A OR2X1_LOC_278/Y 0.59fF
C40110 AND2X1_LOC_729/Y OR2X1_LOC_329/a_36_216# -0.02fF
C40111 AND2X1_LOC_592/Y OR2X1_LOC_424/a_36_216# 0.00fF
C40112 OR2X1_LOC_264/Y OR2X1_LOC_78/A 0.11fF
C40113 OR2X1_LOC_43/A OR2X1_LOC_16/A 0.15fF
C40114 OR2X1_LOC_857/B AND2X1_LOC_56/B 0.05fF
C40115 OR2X1_LOC_318/Y OR2X1_LOC_648/A 0.07fF
C40116 AND2X1_LOC_352/B AND2X1_LOC_654/Y 0.09fF
C40117 OR2X1_LOC_160/B OR2X1_LOC_624/A 0.01fF
C40118 OR2X1_LOC_6/B OR2X1_LOC_510/Y 0.07fF
C40119 AND2X1_LOC_648/B OR2X1_LOC_589/a_8_216# 0.00fF
C40120 OR2X1_LOC_219/B OR2X1_LOC_389/a_8_216# 0.40fF
C40121 AND2X1_LOC_50/a_8_24# D_INPUT_5 0.01fF
C40122 AND2X1_LOC_741/Y OR2X1_LOC_189/Y 0.15fF
C40123 OR2X1_LOC_91/Y AND2X1_LOC_243/Y 0.02fF
C40124 AND2X1_LOC_136/a_8_24# AND2X1_LOC_7/B 0.02fF
C40125 OR2X1_LOC_266/a_8_216# OR2X1_LOC_786/A 0.05fF
C40126 D_INPUT_1 AND2X1_LOC_236/a_36_24# 0.00fF
C40127 OR2X1_LOC_48/B AND2X1_LOC_469/B 0.03fF
C40128 OR2X1_LOC_160/A OR2X1_LOC_35/a_8_216# 0.06fF
C40129 AND2X1_LOC_675/A OR2X1_LOC_142/Y 0.07fF
C40130 AND2X1_LOC_191/B OR2X1_LOC_18/Y 4.50fF
C40131 AND2X1_LOC_651/a_36_24# OR2X1_LOC_762/Y 0.01fF
C40132 OR2X1_LOC_745/Y OR2X1_LOC_746/Y 0.09fF
C40133 OR2X1_LOC_676/Y OR2X1_LOC_375/A 0.08fF
C40134 AND2X1_LOC_729/Y AND2X1_LOC_705/a_8_24# 0.01fF
C40135 OR2X1_LOC_158/A OR2X1_LOC_753/A 0.14fF
C40136 OR2X1_LOC_604/A AND2X1_LOC_319/A 0.01fF
C40137 OR2X1_LOC_358/a_8_216# VDD 0.00fF
C40138 AND2X1_LOC_474/A OR2X1_LOC_427/A 0.07fF
C40139 OR2X1_LOC_661/a_8_216# OR2X1_LOC_78/B 0.01fF
C40140 OR2X1_LOC_405/A OR2X1_LOC_778/a_8_216# 0.03fF
C40141 OR2X1_LOC_818/Y AND2X1_LOC_820/B 0.08fF
C40142 OR2X1_LOC_636/a_8_216# AND2X1_LOC_44/Y 0.15fF
C40143 OR2X1_LOC_538/A OR2X1_LOC_623/a_8_216# 0.01fF
C40144 OR2X1_LOC_648/A OR2X1_LOC_805/A 0.07fF
C40145 AND2X1_LOC_733/Y OR2X1_LOC_48/B 0.03fF
C40146 AND2X1_LOC_436/B AND2X1_LOC_434/Y 0.01fF
C40147 OR2X1_LOC_335/Y AND2X1_LOC_95/Y 0.14fF
C40148 OR2X1_LOC_865/B OR2X1_LOC_756/B 0.01fF
C40149 AND2X1_LOC_465/Y AND2X1_LOC_465/A 0.16fF
C40150 OR2X1_LOC_812/B OR2X1_LOC_391/A 0.04fF
C40151 OR2X1_LOC_6/B OR2X1_LOC_810/A 0.10fF
C40152 AND2X1_LOC_807/Y AND2X1_LOC_663/A 1.20fF
C40153 OR2X1_LOC_851/a_8_216# OR2X1_LOC_87/A 0.05fF
C40154 OR2X1_LOC_834/A OR2X1_LOC_375/A 0.01fF
C40155 AND2X1_LOC_563/A OR2X1_LOC_26/Y 0.03fF
C40156 OR2X1_LOC_507/B AND2X1_LOC_41/A 0.01fF
C40157 OR2X1_LOC_8/Y OR2X1_LOC_44/Y 0.06fF
C40158 AND2X1_LOC_139/B AND2X1_LOC_219/Y 0.07fF
C40159 VDD OR2X1_LOC_588/Y 0.05fF
C40160 AND2X1_LOC_564/B AND2X1_LOC_471/a_8_24# 0.02fF
C40161 OR2X1_LOC_748/A AND2X1_LOC_709/a_36_24# 0.01fF
C40162 OR2X1_LOC_377/a_8_216# OR2X1_LOC_378/A 0.01fF
C40163 AND2X1_LOC_95/Y OR2X1_LOC_435/a_36_216# 0.00fF
C40164 AND2X1_LOC_580/A OR2X1_LOC_59/Y 0.03fF
C40165 OR2X1_LOC_62/B OR2X1_LOC_563/A 0.01fF
C40166 OR2X1_LOC_481/Y OR2X1_LOC_382/A 0.00fF
C40167 OR2X1_LOC_19/B AND2X1_LOC_44/Y 0.10fF
C40168 AND2X1_LOC_514/a_8_24# OR2X1_LOC_6/A 0.01fF
C40169 AND2X1_LOC_40/Y AND2X1_LOC_95/Y 2.37fF
C40170 AND2X1_LOC_642/a_8_24# AND2X1_LOC_642/Y 0.02fF
C40171 AND2X1_LOC_116/B OR2X1_LOC_428/A 0.06fF
C40172 AND2X1_LOC_563/A OR2X1_LOC_89/A 0.02fF
C40173 OR2X1_LOC_185/A OR2X1_LOC_623/B 0.09fF
C40174 AND2X1_LOC_566/B AND2X1_LOC_211/a_36_24# 0.00fF
C40175 AND2X1_LOC_40/Y OR2X1_LOC_633/Y 0.10fF
C40176 OR2X1_LOC_643/A OR2X1_LOC_78/A 0.05fF
C40177 AND2X1_LOC_181/Y AND2X1_LOC_523/Y 0.03fF
C40178 OR2X1_LOC_665/Y AND2X1_LOC_658/A 0.03fF
C40179 AND2X1_LOC_658/A AND2X1_LOC_474/Y 0.03fF
C40180 AND2X1_LOC_732/B OR2X1_LOC_3/Y 0.00fF
C40181 OR2X1_LOC_143/a_8_216# D_INPUT_1 0.12fF
C40182 OR2X1_LOC_778/Y OR2X1_LOC_78/A 0.10fF
C40183 AND2X1_LOC_22/Y D_INPUT_0 0.16fF
C40184 INPUT_0 AND2X1_LOC_55/a_36_24# 0.00fF
C40185 AND2X1_LOC_70/a_8_24# AND2X1_LOC_17/Y 0.01fF
C40186 OR2X1_LOC_139/A OR2X1_LOC_532/B 0.13fF
C40187 AND2X1_LOC_605/Y OR2X1_LOC_36/Y 0.01fF
C40188 AND2X1_LOC_300/a_8_24# OR2X1_LOC_121/B 0.00fF
C40189 OR2X1_LOC_74/A OR2X1_LOC_627/Y 0.14fF
C40190 OR2X1_LOC_848/A OR2X1_LOC_391/a_8_216# 0.02fF
C40191 OR2X1_LOC_837/Y AND2X1_LOC_56/B 0.01fF
C40192 OR2X1_LOC_844/a_8_216# OR2X1_LOC_66/A 0.00fF
C40193 OR2X1_LOC_65/B AND2X1_LOC_266/a_36_24# 0.00fF
C40194 AND2X1_LOC_500/Y OR2X1_LOC_74/A 0.03fF
C40195 OR2X1_LOC_802/a_8_216# OR2X1_LOC_802/A 0.39fF
C40196 AND2X1_LOC_559/a_8_24# OR2X1_LOC_275/Y 0.01fF
C40197 OR2X1_LOC_858/A AND2X1_LOC_3/Y 0.03fF
C40198 OR2X1_LOC_599/A AND2X1_LOC_722/A 0.05fF
C40199 AND2X1_LOC_98/Y OR2X1_LOC_753/A 0.02fF
C40200 AND2X1_LOC_662/B OR2X1_LOC_619/Y 0.02fF
C40201 OR2X1_LOC_756/B OR2X1_LOC_403/B 0.01fF
C40202 AND2X1_LOC_347/Y OR2X1_LOC_748/A 0.04fF
C40203 OR2X1_LOC_429/a_36_216# INPUT_7 0.01fF
C40204 AND2X1_LOC_358/Y OR2X1_LOC_417/A 0.01fF
C40205 OR2X1_LOC_244/A OR2X1_LOC_548/B 0.84fF
C40206 AND2X1_LOC_456/B OR2X1_LOC_26/Y 0.02fF
C40207 OR2X1_LOC_31/Y AND2X1_LOC_214/a_8_24# 0.01fF
C40208 AND2X1_LOC_365/A AND2X1_LOC_661/a_8_24# -0.01fF
C40209 OR2X1_LOC_458/B OR2X1_LOC_778/Y 0.07fF
C40210 AND2X1_LOC_753/B OR2X1_LOC_185/Y 0.21fF
C40211 AND2X1_LOC_19/Y AND2X1_LOC_42/B 0.06fF
C40212 OR2X1_LOC_131/A OR2X1_LOC_246/A 1.22fF
C40213 OR2X1_LOC_604/A AND2X1_LOC_708/a_8_24# 0.01fF
C40214 OR2X1_LOC_589/A AND2X1_LOC_687/Y 0.28fF
C40215 OR2X1_LOC_506/A AND2X1_LOC_43/B 0.15fF
C40216 AND2X1_LOC_729/a_8_24# AND2X1_LOC_800/a_8_24# 0.23fF
C40217 OR2X1_LOC_17/Y OR2X1_LOC_25/Y 0.07fF
C40218 OR2X1_LOC_864/A OR2X1_LOC_502/A 0.03fF
C40219 AND2X1_LOC_568/B OR2X1_LOC_417/Y 0.19fF
C40220 OR2X1_LOC_656/a_8_216# AND2X1_LOC_18/Y 0.02fF
C40221 OR2X1_LOC_159/a_8_216# OR2X1_LOC_46/A 0.01fF
C40222 OR2X1_LOC_427/A OR2X1_LOC_85/A 0.14fF
C40223 AND2X1_LOC_456/B OR2X1_LOC_89/A 0.03fF
C40224 OR2X1_LOC_40/Y OR2X1_LOC_46/A 0.22fF
C40225 OR2X1_LOC_448/B OR2X1_LOC_778/Y 0.05fF
C40226 OR2X1_LOC_160/A OR2X1_LOC_448/Y 0.02fF
C40227 OR2X1_LOC_600/A OR2X1_LOC_19/B 0.08fF
C40228 OR2X1_LOC_158/A AND2X1_LOC_845/Y 0.21fF
C40229 OR2X1_LOC_185/Y OR2X1_LOC_860/a_36_216# 0.00fF
C40230 VDD OR2X1_LOC_772/Y 0.10fF
C40231 OR2X1_LOC_485/a_8_216# OR2X1_LOC_52/B 0.05fF
C40232 AND2X1_LOC_718/a_36_24# OR2X1_LOC_89/A 0.00fF
C40233 OR2X1_LOC_364/A OR2X1_LOC_405/A 0.01fF
C40234 VDD OR2X1_LOC_846/A 0.01fF
C40235 OR2X1_LOC_6/B AND2X1_LOC_133/a_36_24# 0.01fF
C40236 OR2X1_LOC_844/Y OR2X1_LOC_244/Y 0.45fF
C40237 OR2X1_LOC_502/A OR2X1_LOC_240/A 0.03fF
C40238 OR2X1_LOC_313/Y OR2X1_LOC_314/Y 0.22fF
C40239 OR2X1_LOC_185/Y OR2X1_LOC_405/A 0.25fF
C40240 OR2X1_LOC_66/Y OR2X1_LOC_115/B 0.01fF
C40241 OR2X1_LOC_106/a_36_216# AND2X1_LOC_845/Y 0.01fF
C40242 AND2X1_LOC_381/a_8_24# AND2X1_LOC_817/B 0.00fF
C40243 AND2X1_LOC_732/a_36_24# OR2X1_LOC_64/Y 0.00fF
C40244 OR2X1_LOC_479/Y OR2X1_LOC_808/A 0.12fF
C40245 OR2X1_LOC_121/Y OR2X1_LOC_276/A 0.02fF
C40246 OR2X1_LOC_549/Y OR2X1_LOC_577/Y 0.74fF
C40247 AND2X1_LOC_155/a_36_24# OR2X1_LOC_52/B 0.01fF
C40248 OR2X1_LOC_244/A OR2X1_LOC_786/A 0.02fF
C40249 OR2X1_LOC_409/B AND2X1_LOC_771/B 0.01fF
C40250 AND2X1_LOC_784/A OR2X1_LOC_519/a_36_216# 0.01fF
C40251 OR2X1_LOC_600/A AND2X1_LOC_128/a_36_24# 0.01fF
C40252 OR2X1_LOC_508/a_8_216# OR2X1_LOC_506/B 0.01fF
C40253 OR2X1_LOC_40/Y OR2X1_LOC_679/A 0.03fF
C40254 OR2X1_LOC_810/A OR2X1_LOC_523/Y 0.05fF
C40255 INPUT_3 AND2X1_LOC_852/a_36_24# -0.00fF
C40256 OR2X1_LOC_462/B OR2X1_LOC_375/A 0.03fF
C40257 OR2X1_LOC_160/B OR2X1_LOC_447/Y 0.03fF
C40258 OR2X1_LOC_739/A OR2X1_LOC_269/B 0.03fF
C40259 OR2X1_LOC_67/A OR2X1_LOC_44/Y 0.01fF
C40260 OR2X1_LOC_697/Y OR2X1_LOC_696/Y 0.44fF
C40261 OR2X1_LOC_324/a_8_216# OR2X1_LOC_479/Y 0.05fF
C40262 AND2X1_LOC_318/a_8_24# OR2X1_LOC_36/Y 0.01fF
C40263 OR2X1_LOC_641/Y AND2X1_LOC_519/a_36_24# 0.01fF
C40264 OR2X1_LOC_754/A OR2X1_LOC_92/Y 0.02fF
C40265 OR2X1_LOC_604/A OR2X1_LOC_604/a_8_216# 0.14fF
C40266 OR2X1_LOC_40/Y AND2X1_LOC_227/Y 0.03fF
C40267 OR2X1_LOC_222/A OR2X1_LOC_358/B 0.72fF
C40268 AND2X1_LOC_783/B AND2X1_LOC_779/Y 0.33fF
C40269 AND2X1_LOC_784/A AND2X1_LOC_170/a_36_24# 0.01fF
C40270 OR2X1_LOC_96/Y OR2X1_LOC_95/Y 0.01fF
C40271 OR2X1_LOC_687/Y AND2X1_LOC_56/B 1.64fF
C40272 AND2X1_LOC_736/Y OR2X1_LOC_527/Y 0.07fF
C40273 D_INPUT_3 AND2X1_LOC_243/Y 0.07fF
C40274 AND2X1_LOC_337/B OR2X1_LOC_619/Y 0.05fF
C40275 OR2X1_LOC_3/Y OR2X1_LOC_625/Y 0.04fF
C40276 OR2X1_LOC_357/B OR2X1_LOC_365/B 0.02fF
C40277 OR2X1_LOC_87/Y OR2X1_LOC_99/Y 0.00fF
C40278 AND2X1_LOC_777/a_8_24# AND2X1_LOC_702/Y 0.01fF
C40279 OR2X1_LOC_64/Y AND2X1_LOC_651/a_8_24# 0.01fF
C40280 OR2X1_LOC_91/A AND2X1_LOC_477/A 0.00fF
C40281 OR2X1_LOC_47/Y AND2X1_LOC_477/Y 0.02fF
C40282 AND2X1_LOC_365/A AND2X1_LOC_336/a_8_24# 0.20fF
C40283 AND2X1_LOC_217/Y AND2X1_LOC_660/A 0.00fF
C40284 VDD OR2X1_LOC_145/Y 0.12fF
C40285 AND2X1_LOC_359/B OR2X1_LOC_248/Y 1.03fF
C40286 OR2X1_LOC_557/A OR2X1_LOC_404/a_8_216# 0.01fF
C40287 OR2X1_LOC_276/B OR2X1_LOC_66/A 0.07fF
C40288 OR2X1_LOC_244/B D_INPUT_0 0.02fF
C40289 OR2X1_LOC_265/a_8_216# OR2X1_LOC_245/a_8_216# 0.47fF
C40290 AND2X1_LOC_554/Y AND2X1_LOC_557/a_8_24# 0.03fF
C40291 AND2X1_LOC_95/Y OR2X1_LOC_475/Y 0.03fF
C40292 OR2X1_LOC_44/Y OR2X1_LOC_52/B 0.80fF
C40293 OR2X1_LOC_95/Y AND2X1_LOC_663/A 0.03fF
C40294 OR2X1_LOC_356/A OR2X1_LOC_356/a_36_216# 0.00fF
C40295 OR2X1_LOC_635/a_8_216# AND2X1_LOC_51/Y 0.01fF
C40296 AND2X1_LOC_191/Y AND2X1_LOC_580/A 0.03fF
C40297 AND2X1_LOC_658/B GATE_811 0.03fF
C40298 OR2X1_LOC_485/A OR2X1_LOC_497/a_8_216# 0.02fF
C40299 OR2X1_LOC_45/B OR2X1_LOC_88/Y 0.03fF
C40300 AND2X1_LOC_336/a_8_24# OR2X1_LOC_43/A 0.01fF
C40301 OR2X1_LOC_620/B AND2X1_LOC_56/B 0.00fF
C40302 AND2X1_LOC_476/A OR2X1_LOC_59/Y 0.09fF
C40303 AND2X1_LOC_489/Y OR2X1_LOC_44/Y 0.03fF
C40304 OR2X1_LOC_458/a_36_216# OR2X1_LOC_532/B 0.00fF
C40305 OR2X1_LOC_528/Y AND2X1_LOC_793/Y 0.19fF
C40306 OR2X1_LOC_45/B OR2X1_LOC_172/Y 0.25fF
C40307 AND2X1_LOC_711/Y AND2X1_LOC_580/A 0.03fF
C40308 AND2X1_LOC_31/Y OR2X1_LOC_34/a_8_216# 0.14fF
C40309 OR2X1_LOC_76/A OR2X1_LOC_161/A 0.02fF
C40310 OR2X1_LOC_126/a_8_216# AND2X1_LOC_852/Y 0.04fF
C40311 OR2X1_LOC_673/Y AND2X1_LOC_42/B 0.02fF
C40312 OR2X1_LOC_850/B OR2X1_LOC_532/B 0.07fF
C40313 AND2X1_LOC_470/a_8_24# OR2X1_LOC_427/A 0.02fF
C40314 AND2X1_LOC_580/A OR2X1_LOC_70/Y 0.02fF
C40315 OR2X1_LOC_49/A OR2X1_LOC_68/B 2.63fF
C40316 OR2X1_LOC_449/a_8_216# OR2X1_LOC_453/A -0.00fF
C40317 AND2X1_LOC_641/Y AND2X1_LOC_650/Y 0.04fF
C40318 OR2X1_LOC_404/Y OR2X1_LOC_668/Y 0.01fF
C40319 OR2X1_LOC_770/B OR2X1_LOC_68/B 0.05fF
C40320 OR2X1_LOC_19/B OR2X1_LOC_619/Y 0.07fF
C40321 OR2X1_LOC_854/a_36_216# D_INPUT_0 0.03fF
C40322 INPUT_3 OR2X1_LOC_54/Y 0.18fF
C40323 AND2X1_LOC_191/B AND2X1_LOC_620/Y 0.01fF
C40324 OR2X1_LOC_651/a_36_216# OR2X1_LOC_654/A 0.00fF
C40325 AND2X1_LOC_493/a_8_24# AND2X1_LOC_717/B 0.00fF
C40326 OR2X1_LOC_329/B OR2X1_LOC_47/Y 0.05fF
C40327 AND2X1_LOC_59/Y OR2X1_LOC_476/B 0.11fF
C40328 OR2X1_LOC_235/B OR2X1_LOC_84/A 0.02fF
C40329 OR2X1_LOC_416/Y OR2X1_LOC_39/A 0.01fF
C40330 AND2X1_LOC_497/a_8_24# AND2X1_LOC_18/Y 0.04fF
C40331 AND2X1_LOC_625/a_36_24# OR2X1_LOC_598/A 0.01fF
C40332 AND2X1_LOC_717/B OR2X1_LOC_89/A 0.06fF
C40333 AND2X1_LOC_11/Y AND2X1_LOC_7/Y 0.00fF
C40334 AND2X1_LOC_59/Y OR2X1_LOC_650/Y 0.01fF
C40335 AND2X1_LOC_7/B OR2X1_LOC_704/a_8_216# 0.00fF
C40336 OR2X1_LOC_755/A OR2X1_LOC_44/Y 0.00fF
C40337 OR2X1_LOC_324/A OR2X1_LOC_532/B 0.01fF
C40338 AND2X1_LOC_211/B AND2X1_LOC_640/Y 0.11fF
C40339 OR2X1_LOC_89/A OR2X1_LOC_258/a_36_216# 0.02fF
C40340 AND2X1_LOC_721/Y OR2X1_LOC_437/A 0.02fF
C40341 OR2X1_LOC_137/B OR2X1_LOC_62/B 0.04fF
C40342 OR2X1_LOC_610/a_8_216# AND2X1_LOC_47/Y 0.05fF
C40343 AND2X1_LOC_90/a_36_24# OR2X1_LOC_80/A 0.01fF
C40344 OR2X1_LOC_267/Y OR2X1_LOC_141/a_8_216# 0.01fF
C40345 AND2X1_LOC_719/Y AND2X1_LOC_657/A 0.10fF
C40346 OR2X1_LOC_148/A OR2X1_LOC_161/A 0.01fF
C40347 AND2X1_LOC_64/Y AND2X1_LOC_239/a_8_24# 0.01fF
C40348 AND2X1_LOC_95/Y AND2X1_LOC_826/a_8_24# -0.01fF
C40349 OR2X1_LOC_604/A OR2X1_LOC_331/Y 0.07fF
C40350 OR2X1_LOC_481/Y OR2X1_LOC_261/Y 0.22fF
C40351 AND2X1_LOC_375/a_8_24# OR2X1_LOC_409/B 0.01fF
C40352 AND2X1_LOC_798/Y OR2X1_LOC_7/A 0.05fF
C40353 OR2X1_LOC_22/Y OR2X1_LOC_6/A 0.03fF
C40354 OR2X1_LOC_287/B AND2X1_LOC_51/Y 0.07fF
C40355 OR2X1_LOC_160/B OR2X1_LOC_513/a_8_216# 0.03fF
C40356 AND2X1_LOC_22/Y OR2X1_LOC_339/A 0.12fF
C40357 OR2X1_LOC_66/A OR2X1_LOC_779/B 0.14fF
C40358 OR2X1_LOC_329/B AND2X1_LOC_405/a_36_24# 0.01fF
C40359 OR2X1_LOC_864/A AND2X1_LOC_48/A 0.03fF
C40360 OR2X1_LOC_756/B OR2X1_LOC_493/Y 0.03fF
C40361 OR2X1_LOC_22/A AND2X1_LOC_472/B 0.01fF
C40362 AND2X1_LOC_70/Y OR2X1_LOC_568/a_8_216# 0.03fF
C40363 AND2X1_LOC_580/A OR2X1_LOC_504/Y 0.15fF
C40364 OR2X1_LOC_417/A AND2X1_LOC_668/a_8_24# 0.01fF
C40365 OR2X1_LOC_447/Y OR2X1_LOC_779/a_36_216# 0.02fF
C40366 AND2X1_LOC_12/Y OR2X1_LOC_276/A 0.29fF
C40367 OR2X1_LOC_849/A OR2X1_LOC_814/A 0.03fF
C40368 AND2X1_LOC_708/a_36_24# OR2X1_LOC_7/A 0.01fF
C40369 VDD OR2X1_LOC_348/B 0.23fF
C40370 OR2X1_LOC_665/Y AND2X1_LOC_814/a_8_24# 0.23fF
C40371 OR2X1_LOC_7/A OR2X1_LOC_46/A 0.03fF
C40372 OR2X1_LOC_482/Y OR2X1_LOC_437/A 0.17fF
C40373 OR2X1_LOC_316/Y AND2X1_LOC_318/Y 0.00fF
C40374 OR2X1_LOC_310/Y AND2X1_LOC_222/Y 0.01fF
C40375 AND2X1_LOC_130/a_8_24# OR2X1_LOC_13/B 0.03fF
C40376 OR2X1_LOC_743/A AND2X1_LOC_687/A 0.07fF
C40377 AND2X1_LOC_81/B OR2X1_LOC_241/Y 0.07fF
C40378 OR2X1_LOC_375/A OR2X1_LOC_200/Y 0.02fF
C40379 OR2X1_LOC_441/a_8_216# AND2X1_LOC_222/Y 0.01fF
C40380 AND2X1_LOC_113/Y OR2X1_LOC_47/Y 0.01fF
C40381 AND2X1_LOC_420/a_8_24# AND2X1_LOC_43/B 0.16fF
C40382 OR2X1_LOC_557/A OR2X1_LOC_403/a_36_216# 0.00fF
C40383 AND2X1_LOC_86/Y OR2X1_LOC_84/Y 0.05fF
C40384 OR2X1_LOC_320/Y OR2X1_LOC_46/A 0.16fF
C40385 AND2X1_LOC_159/a_8_24# AND2X1_LOC_47/Y 0.02fF
C40386 OR2X1_LOC_502/A OR2X1_LOC_608/Y 0.01fF
C40387 OR2X1_LOC_810/A AND2X1_LOC_47/Y 4.20fF
C40388 OR2X1_LOC_19/B AND2X1_LOC_4/a_36_24# 0.01fF
C40389 AND2X1_LOC_555/Y OR2X1_LOC_494/A 0.01fF
C40390 OR2X1_LOC_307/a_8_216# AND2X1_LOC_47/Y 0.01fF
C40391 OR2X1_LOC_201/A AND2X1_LOC_31/Y 0.01fF
C40392 D_INPUT_5 AND2X1_LOC_429/a_8_24# 0.01fF
C40393 OR2X1_LOC_157/a_8_216# OR2X1_LOC_51/a_8_216# 0.47fF
C40394 OR2X1_LOC_792/Y OR2X1_LOC_675/Y 0.01fF
C40395 OR2X1_LOC_181/B OR2X1_LOC_192/B 0.11fF
C40396 AND2X1_LOC_393/a_8_24# OR2X1_LOC_84/A 0.20fF
C40397 OR2X1_LOC_676/Y OR2X1_LOC_515/Y 0.09fF
C40398 AND2X1_LOC_227/Y OR2X1_LOC_7/A 0.13fF
C40399 AND2X1_LOC_64/Y OR2X1_LOC_97/A 0.06fF
C40400 AND2X1_LOC_91/B AND2X1_LOC_91/a_8_24# 0.05fF
C40401 INPUT_0 OR2X1_LOC_71/A 0.19fF
C40402 AND2X1_LOC_447/Y OR2X1_LOC_424/Y 0.04fF
C40403 AND2X1_LOC_727/A AND2X1_LOC_856/a_8_24# 0.01fF
C40404 AND2X1_LOC_308/a_8_24# AND2X1_LOC_863/A 0.19fF
C40405 OR2X1_LOC_614/a_8_216# AND2X1_LOC_3/Y 0.02fF
C40406 AND2X1_LOC_229/a_8_24# AND2X1_LOC_226/a_8_24# 0.23fF
C40407 AND2X1_LOC_644/a_8_24# AND2X1_LOC_655/A 0.11fF
C40408 OR2X1_LOC_22/Y OR2X1_LOC_43/a_36_216# 0.03fF
C40409 OR2X1_LOC_835/Y AND2X1_LOC_51/Y 0.16fF
C40410 OR2X1_LOC_148/A AND2X1_LOC_51/Y 0.10fF
C40411 AND2X1_LOC_543/Y OR2X1_LOC_373/Y 0.14fF
C40412 OR2X1_LOC_70/Y OR2X1_LOC_72/a_8_216# 0.02fF
C40413 OR2X1_LOC_510/Y OR2X1_LOC_598/A 0.14fF
C40414 OR2X1_LOC_53/Y OR2X1_LOC_428/A 0.32fF
C40415 OR2X1_LOC_405/A AND2X1_LOC_432/a_8_24# 0.01fF
C40416 AND2X1_LOC_12/Y AND2X1_LOC_429/a_8_24# 0.20fF
C40417 OR2X1_LOC_178/a_36_216# OR2X1_LOC_183/Y 0.00fF
C40418 OR2X1_LOC_70/Y AND2X1_LOC_476/A 0.07fF
C40419 AND2X1_LOC_12/Y OR2X1_LOC_512/Y 0.02fF
C40420 OR2X1_LOC_57/a_8_216# OR2X1_LOC_19/a_8_216# 0.47fF
C40421 OR2X1_LOC_469/Y OR2X1_LOC_705/a_36_216# 0.01fF
C40422 OR2X1_LOC_156/Y OR2X1_LOC_160/Y 0.18fF
C40423 OR2X1_LOC_836/Y OR2X1_LOC_835/Y 0.14fF
C40424 AND2X1_LOC_1/Y OR2X1_LOC_651/A -0.00fF
C40425 OR2X1_LOC_517/A OR2X1_LOC_13/B 0.10fF
C40426 AND2X1_LOC_802/Y OR2X1_LOC_428/A 0.05fF
C40427 OR2X1_LOC_447/a_8_216# OR2X1_LOC_724/A 0.01fF
C40428 OR2X1_LOC_813/Y OR2X1_LOC_7/A 0.07fF
C40429 OR2X1_LOC_3/Y OR2X1_LOC_3/B 0.04fF
C40430 OR2X1_LOC_831/a_8_216# OR2X1_LOC_228/Y 0.01fF
C40431 OR2X1_LOC_791/B OR2X1_LOC_345/a_36_216# 0.01fF
C40432 OR2X1_LOC_810/A OR2X1_LOC_598/A 0.10fF
C40433 OR2X1_LOC_479/Y OR2X1_LOC_795/a_8_216# 0.01fF
C40434 OR2X1_LOC_39/A OR2X1_LOC_80/A 0.76fF
C40435 OR2X1_LOC_323/A OR2X1_LOC_600/A 0.03fF
C40436 AND2X1_LOC_40/Y OR2X1_LOC_788/B 0.04fF
C40437 OR2X1_LOC_154/A OR2X1_LOC_560/A 0.03fF
C40438 AND2X1_LOC_22/Y OR2X1_LOC_831/A 0.38fF
C40439 OR2X1_LOC_344/A OR2X1_LOC_578/a_36_216# 0.00fF
C40440 OR2X1_LOC_18/Y OR2X1_LOC_164/a_8_216# 0.07fF
C40441 OR2X1_LOC_433/Y OR2X1_LOC_423/Y 0.01fF
C40442 OR2X1_LOC_64/a_36_216# OR2X1_LOC_22/A 0.02fF
C40443 OR2X1_LOC_87/B OR2X1_LOC_68/B 0.07fF
C40444 OR2X1_LOC_440/A OR2X1_LOC_814/A 0.07fF
C40445 OR2X1_LOC_7/A OR2X1_LOC_753/Y 0.46fF
C40446 AND2X1_LOC_22/Y OR2X1_LOC_598/Y 0.06fF
C40447 AND2X1_LOC_116/Y AND2X1_LOC_216/A 0.24fF
C40448 OR2X1_LOC_479/Y OR2X1_LOC_374/Y 0.07fF
C40449 OR2X1_LOC_154/a_8_216# OR2X1_LOC_156/A 0.41fF
C40450 AND2X1_LOC_776/Y OR2X1_LOC_56/A 0.15fF
C40451 OR2X1_LOC_619/Y AND2X1_LOC_608/a_8_24# 0.06fF
C40452 AND2X1_LOC_163/a_36_24# OR2X1_LOC_161/B 0.00fF
C40453 OR2X1_LOC_302/B AND2X1_LOC_64/Y 0.08fF
C40454 AND2X1_LOC_110/Y AND2X1_LOC_44/Y 0.03fF
C40455 OR2X1_LOC_188/Y OR2X1_LOC_741/Y 1.10fF
C40456 OR2X1_LOC_673/B OR2X1_LOC_621/A 0.02fF
C40457 AND2X1_LOC_91/B OR2X1_LOC_78/A 0.19fF
C40458 AND2X1_LOC_612/B OR2X1_LOC_68/B 0.25fF
C40459 AND2X1_LOC_3/Y AND2X1_LOC_31/Y 1.40fF
C40460 AND2X1_LOC_707/Y AND2X1_LOC_447/Y 0.04fF
C40461 OR2X1_LOC_478/Y OR2X1_LOC_467/A 0.01fF
C40462 OR2X1_LOC_2/Y INPUT_6 0.01fF
C40463 OR2X1_LOC_13/a_36_216# OR2X1_LOC_13/Y 0.00fF
C40464 OR2X1_LOC_805/A OR2X1_LOC_112/A 0.09fF
C40465 OR2X1_LOC_45/B OR2X1_LOC_8/Y 0.00fF
C40466 AND2X1_LOC_65/A AND2X1_LOC_265/a_8_24# 0.03fF
C40467 AND2X1_LOC_469/Y AND2X1_LOC_477/Y 0.23fF
C40468 OR2X1_LOC_114/B OR2X1_LOC_294/Y 0.01fF
C40469 OR2X1_LOC_696/A OR2X1_LOC_586/a_8_216# 0.01fF
C40470 OR2X1_LOC_33/B OR2X1_LOC_68/B 0.01fF
C40471 OR2X1_LOC_856/a_8_216# OR2X1_LOC_198/A 0.00fF
C40472 AND2X1_LOC_22/Y OR2X1_LOC_795/B 0.08fF
C40473 OR2X1_LOC_502/A OR2X1_LOC_397/a_8_216# 0.01fF
C40474 OR2X1_LOC_375/A AND2X1_LOC_591/a_8_24# 0.01fF
C40475 OR2X1_LOC_486/Y AND2X1_LOC_18/Y 0.03fF
C40476 OR2X1_LOC_134/a_8_216# OR2X1_LOC_92/Y 0.30fF
C40477 OR2X1_LOC_709/A OR2X1_LOC_66/A 0.07fF
C40478 AND2X1_LOC_388/Y AND2X1_LOC_535/Y 0.03fF
C40479 AND2X1_LOC_675/Y OR2X1_LOC_816/A 0.01fF
C40480 VDD AND2X1_LOC_65/A 0.27fF
C40481 OR2X1_LOC_715/B OR2X1_LOC_6/B 0.15fF
C40482 AND2X1_LOC_544/Y OR2X1_LOC_438/Y 0.01fF
C40483 OR2X1_LOC_335/Y AND2X1_LOC_22/Y 0.09fF
C40484 AND2X1_LOC_64/Y OR2X1_LOC_475/B 0.57fF
C40485 OR2X1_LOC_6/B AND2X1_LOC_626/a_8_24# 0.04fF
C40486 AND2X1_LOC_509/Y AND2X1_LOC_244/A 0.03fF
C40487 OR2X1_LOC_244/A OR2X1_LOC_84/Y 0.05fF
C40488 OR2X1_LOC_604/A OR2X1_LOC_765/a_36_216# 0.00fF
C40489 OR2X1_LOC_102/a_8_216# OR2X1_LOC_8/Y 0.05fF
C40490 OR2X1_LOC_814/A OR2X1_LOC_366/a_36_216# 0.00fF
C40491 AND2X1_LOC_361/a_8_24# AND2X1_LOC_768/a_8_24# 0.23fF
C40492 AND2X1_LOC_556/a_8_24# OR2X1_LOC_816/A 0.07fF
C40493 AND2X1_LOC_719/Y VDD 1.87fF
C40494 AND2X1_LOC_555/Y OR2X1_LOC_427/A 0.10fF
C40495 OR2X1_LOC_47/Y GATE_811 0.03fF
C40496 OR2X1_LOC_510/A VDD 0.19fF
C40497 AND2X1_LOC_82/Y OR2X1_LOC_78/a_8_216# 0.01fF
C40498 AND2X1_LOC_83/a_8_24# OR2X1_LOC_78/B 0.03fF
C40499 AND2X1_LOC_22/Y AND2X1_LOC_48/a_36_24# 0.00fF
C40500 AND2X1_LOC_191/a_8_24# AND2X1_LOC_866/B 0.01fF
C40501 OR2X1_LOC_36/Y OR2X1_LOC_395/a_8_216# 0.02fF
C40502 AND2X1_LOC_40/Y AND2X1_LOC_22/Y 0.15fF
C40503 OR2X1_LOC_61/a_36_216# AND2X1_LOC_7/B 0.00fF
C40504 OR2X1_LOC_644/B AND2X1_LOC_36/Y 0.02fF
C40505 OR2X1_LOC_680/a_8_216# OR2X1_LOC_525/Y 0.01fF
C40506 OR2X1_LOC_241/Y OR2X1_LOC_66/Y 0.02fF
C40507 OR2X1_LOC_648/B OR2X1_LOC_648/A 0.19fF
C40508 OR2X1_LOC_461/a_8_216# OR2X1_LOC_461/B 0.00fF
C40509 AND2X1_LOC_253/a_8_24# OR2X1_LOC_580/B 0.07fF
C40510 OR2X1_LOC_626/Y OR2X1_LOC_627/Y 0.01fF
C40511 OR2X1_LOC_64/Y OR2X1_LOC_71/A 0.08fF
C40512 OR2X1_LOC_528/Y AND2X1_LOC_548/Y 0.06fF
C40513 OR2X1_LOC_661/A OR2X1_LOC_78/B 0.01fF
C40514 OR2X1_LOC_465/Y AND2X1_LOC_7/B 0.17fF
C40515 OR2X1_LOC_290/Y OR2X1_LOC_12/Y 0.03fF
C40516 OR2X1_LOC_155/a_8_216# OR2X1_LOC_803/a_8_216# 0.47fF
C40517 AND2X1_LOC_70/Y OR2X1_LOC_66/A 6.41fF
C40518 OR2X1_LOC_833/Y OR2X1_LOC_840/A 0.04fF
C40519 OR2X1_LOC_45/B AND2X1_LOC_76/Y 0.03fF
C40520 OR2X1_LOC_641/a_8_216# AND2X1_LOC_92/Y 0.01fF
C40521 AND2X1_LOC_70/Y OR2X1_LOC_841/A 0.01fF
C40522 AND2X1_LOC_91/B OR2X1_LOC_602/A 0.05fF
C40523 OR2X1_LOC_597/A OR2X1_LOC_744/A 0.03fF
C40524 OR2X1_LOC_616/a_8_216# GATE_579 0.01fF
C40525 OR2X1_LOC_616/Y AND2X1_LOC_580/a_8_24# 0.00fF
C40526 OR2X1_LOC_604/A AND2X1_LOC_605/Y 0.01fF
C40527 AND2X1_LOC_727/a_8_24# AND2X1_LOC_550/A 0.07fF
C40528 OR2X1_LOC_40/Y AND2X1_LOC_722/A 0.23fF
C40529 AND2X1_LOC_40/Y OR2X1_LOC_621/A 0.22fF
C40530 OR2X1_LOC_471/B OR2X1_LOC_741/Y 0.01fF
C40531 OR2X1_LOC_599/Y AND2X1_LOC_644/a_8_24# 0.05fF
C40532 AND2X1_LOC_425/a_8_24# INPUT_6 0.02fF
C40533 OR2X1_LOC_178/Y OR2X1_LOC_744/A 0.03fF
C40534 AND2X1_LOC_555/Y AND2X1_LOC_363/A 0.00fF
C40535 OR2X1_LOC_89/A AND2X1_LOC_439/a_36_24# 0.00fF
C40536 OR2X1_LOC_86/A OR2X1_LOC_67/Y 0.01fF
C40537 AND2X1_LOC_392/a_8_24# OR2X1_LOC_51/Y 0.01fF
C40538 AND2X1_LOC_723/Y OR2X1_LOC_600/A 0.07fF
C40539 AND2X1_LOC_56/B AND2X1_LOC_829/a_8_24# 0.18fF
C40540 AND2X1_LOC_189/a_8_24# OR2X1_LOC_741/Y 0.14fF
C40541 OR2X1_LOC_664/Y AND2X1_LOC_44/Y 0.03fF
C40542 OR2X1_LOC_664/a_36_216# OR2X1_LOC_161/B 0.00fF
C40543 OR2X1_LOC_591/Y OR2X1_LOC_48/B 0.03fF
C40544 AND2X1_LOC_95/Y OR2X1_LOC_356/A 0.08fF
C40545 OR2X1_LOC_751/Y OR2X1_LOC_600/A 0.23fF
C40546 INPUT_0 OR2X1_LOC_59/Y 0.03fF
C40547 AND2X1_LOC_91/B OR2X1_LOC_155/A 0.15fF
C40548 OR2X1_LOC_574/A OR2X1_LOC_115/B 0.07fF
C40549 OR2X1_LOC_3/Y OR2X1_LOC_767/Y 0.02fF
C40550 AND2X1_LOC_696/a_8_24# OR2X1_LOC_779/A 0.08fF
C40551 OR2X1_LOC_238/Y AND2X1_LOC_241/a_8_24# 0.05fF
C40552 OR2X1_LOC_620/Y AND2X1_LOC_299/a_8_24# 0.04fF
C40553 OR2X1_LOC_45/B AND2X1_LOC_374/Y 0.01fF
C40554 OR2X1_LOC_186/Y OR2X1_LOC_802/Y 0.01fF
C40555 AND2X1_LOC_729/Y OR2X1_LOC_158/A 0.07fF
C40556 OR2X1_LOC_256/Y OR2X1_LOC_744/A 0.07fF
C40557 AND2X1_LOC_50/Y OR2X1_LOC_638/B 0.00fF
C40558 AND2X1_LOC_452/Y OR2X1_LOC_765/Y 0.78fF
C40559 OR2X1_LOC_45/B OR2X1_LOC_52/B 0.29fF
C40560 AND2X1_LOC_91/B OR2X1_LOC_392/a_8_216# 0.02fF
C40561 OR2X1_LOC_186/Y OR2X1_LOC_468/Y 0.08fF
C40562 OR2X1_LOC_409/B OR2X1_LOC_376/a_8_216# 0.01fF
C40563 OR2X1_LOC_305/Y OR2X1_LOC_12/Y 0.00fF
C40564 OR2X1_LOC_323/A OR2X1_LOC_372/a_8_216# 0.01fF
C40565 OR2X1_LOC_121/Y OR2X1_LOC_114/Y 0.00fF
C40566 OR2X1_LOC_864/A OR2X1_LOC_489/A 0.05fF
C40567 OR2X1_LOC_231/a_8_216# AND2X1_LOC_18/Y 0.01fF
C40568 VDD OR2X1_LOC_181/B 0.10fF
C40569 OR2X1_LOC_434/A OR2X1_LOC_339/A 0.20fF
C40570 OR2X1_LOC_785/B AND2X1_LOC_92/Y 0.02fF
C40571 OR2X1_LOC_51/Y OR2X1_LOC_427/A 2.02fF
C40572 OR2X1_LOC_614/Y OR2X1_LOC_87/A 0.02fF
C40573 OR2X1_LOC_12/Y AND2X1_LOC_446/a_8_24# 0.01fF
C40574 OR2X1_LOC_160/B OR2X1_LOC_161/A 0.18fF
C40575 OR2X1_LOC_814/A AND2X1_LOC_238/a_8_24# 0.01fF
C40576 AND2X1_LOC_286/a_8_24# OR2X1_LOC_278/Y 0.01fF
C40577 OR2X1_LOC_774/Y OR2X1_LOC_489/A 0.00fF
C40578 AND2X1_LOC_203/a_8_24# AND2X1_LOC_215/A 0.01fF
C40579 OR2X1_LOC_134/Y AND2X1_LOC_663/B 0.03fF
C40580 AND2X1_LOC_53/Y AND2X1_LOC_36/Y 0.02fF
C40581 AND2X1_LOC_523/Y AND2X1_LOC_455/a_8_24# -0.00fF
C40582 VDD OR2X1_LOC_252/Y -0.00fF
C40583 D_INPUT_1 OR2X1_LOC_558/A 0.31fF
C40584 VDD OR2X1_LOC_313/Y 0.22fF
C40585 OR2X1_LOC_279/Y AND2X1_LOC_287/B 0.01fF
C40586 OR2X1_LOC_9/Y OR2X1_LOC_36/Y 0.00fF
C40587 AND2X1_LOC_784/A OR2X1_LOC_158/A 0.09fF
C40588 AND2X1_LOC_206/Y AND2X1_LOC_215/A 0.23fF
C40589 VDD OR2X1_LOC_659/a_8_216# 0.00fF
C40590 VDD AND2X1_LOC_655/A 1.21fF
C40591 OR2X1_LOC_49/A OR2X1_LOC_74/A 0.09fF
C40592 OR2X1_LOC_298/Y OR2X1_LOC_426/B 0.01fF
C40593 AND2X1_LOC_576/Y AND2X1_LOC_500/B 0.01fF
C40594 AND2X1_LOC_72/Y OR2X1_LOC_78/A 0.03fF
C40595 AND2X1_LOC_42/B AND2X1_LOC_277/a_8_24# 0.09fF
C40596 OR2X1_LOC_599/A OR2X1_LOC_40/Y 0.08fF
C40597 AND2X1_LOC_454/A OR2X1_LOC_421/Y 0.15fF
C40598 OR2X1_LOC_799/A OR2X1_LOC_78/A 0.23fF
C40599 AND2X1_LOC_143/a_8_24# OR2X1_LOC_502/A 0.02fF
C40600 OR2X1_LOC_44/Y AND2X1_LOC_244/a_8_24# 0.01fF
C40601 AND2X1_LOC_243/Y AND2X1_LOC_806/A 0.03fF
C40602 AND2X1_LOC_719/Y OR2X1_LOC_251/Y 0.01fF
C40603 OR2X1_LOC_151/A OR2X1_LOC_355/B 0.08fF
C40604 AND2X1_LOC_658/B AND2X1_LOC_580/A 0.03fF
C40605 AND2X1_LOC_753/B AND2X1_LOC_52/a_8_24# 0.02fF
C40606 OR2X1_LOC_3/Y OR2X1_LOC_584/a_8_216# 0.02fF
C40607 AND2X1_LOC_59/Y AND2X1_LOC_437/a_8_24# 0.03fF
C40608 OR2X1_LOC_864/A OR2X1_LOC_772/A 0.37fF
C40609 OR2X1_LOC_6/B AND2X1_LOC_81/a_8_24# 0.03fF
C40610 VDD OR2X1_LOC_81/a_8_216# 0.21fF
C40611 OR2X1_LOC_40/Y OR2X1_LOC_93/a_8_216# 0.01fF
C40612 OR2X1_LOC_40/Y AND2X1_LOC_267/a_36_24# 0.00fF
C40613 OR2X1_LOC_22/Y OR2X1_LOC_184/a_8_216# 0.03fF
C40614 AND2X1_LOC_390/B OR2X1_LOC_829/A 0.12fF
C40615 OR2X1_LOC_774/Y OR2X1_LOC_772/A 0.00fF
C40616 AND2X1_LOC_675/Y AND2X1_LOC_807/Y 0.22fF
C40617 OR2X1_LOC_673/A AND2X1_LOC_36/Y 0.03fF
C40618 OR2X1_LOC_11/Y OR2X1_LOC_59/Y 0.01fF
C40619 AND2X1_LOC_61/Y OR2X1_LOC_36/Y 0.12fF
C40620 OR2X1_LOC_49/A OR2X1_LOC_261/A 0.02fF
C40621 AND2X1_LOC_753/B AND2X1_LOC_53/a_8_24# 0.06fF
C40622 OR2X1_LOC_223/A AND2X1_LOC_36/Y 0.04fF
C40623 AND2X1_LOC_307/a_8_24# AND2X1_LOC_774/A 0.06fF
C40624 OR2X1_LOC_6/B OR2X1_LOC_73/a_8_216# 0.05fF
C40625 OR2X1_LOC_405/A OR2X1_LOC_798/Y 0.03fF
C40626 OR2X1_LOC_426/A AND2X1_LOC_450/a_8_24# 0.01fF
C40627 AND2X1_LOC_555/a_8_24# OR2X1_LOC_3/Y 0.01fF
C40628 OR2X1_LOC_438/Y AND2X1_LOC_550/A 0.04fF
C40629 OR2X1_LOC_40/Y OR2X1_LOC_258/a_8_216# 0.01fF
C40630 OR2X1_LOC_417/Y OR2X1_LOC_12/Y 1.04fF
C40631 OR2X1_LOC_849/A OR2X1_LOC_244/Y 0.20fF
C40632 OR2X1_LOC_485/A AND2X1_LOC_614/a_8_24# 0.01fF
C40633 AND2X1_LOC_724/Y AND2X1_LOC_645/A 1.03fF
C40634 AND2X1_LOC_560/B OR2X1_LOC_59/Y 0.03fF
C40635 OR2X1_LOC_92/Y OR2X1_LOC_118/Y 0.06fF
C40636 OR2X1_LOC_311/Y OR2X1_LOC_12/Y 0.02fF
C40637 OR2X1_LOC_421/A OR2X1_LOC_17/Y 0.00fF
C40638 OR2X1_LOC_97/A AND2X1_LOC_600/a_8_24# 0.01fF
C40639 AND2X1_LOC_721/Y AND2X1_LOC_845/Y 0.02fF
C40640 INPUT_1 OR2X1_LOC_428/A 0.60fF
C40641 OR2X1_LOC_40/Y AND2X1_LOC_389/a_36_24# 0.02fF
C40642 AND2X1_LOC_190/a_8_24# OR2X1_LOC_485/A 0.01fF
C40643 OR2X1_LOC_109/Y AND2X1_LOC_841/B 0.02fF
C40644 AND2X1_LOC_81/B OR2X1_LOC_216/A 0.20fF
C40645 AND2X1_LOC_538/Y OR2X1_LOC_12/Y 0.01fF
C40646 AND2X1_LOC_120/a_8_24# AND2X1_LOC_860/A 0.02fF
C40647 OR2X1_LOC_663/A OR2X1_LOC_673/Y 0.03fF
C40648 AND2X1_LOC_123/a_36_24# OR2X1_LOC_56/A 0.00fF
C40649 OR2X1_LOC_808/B OR2X1_LOC_87/A 0.20fF
C40650 AND2X1_LOC_43/B OR2X1_LOC_737/A 0.09fF
C40651 OR2X1_LOC_185/A OR2X1_LOC_833/B 0.03fF
C40652 OR2X1_LOC_186/Y OR2X1_LOC_471/Y 0.07fF
C40653 OR2X1_LOC_705/B AND2X1_LOC_36/Y 0.08fF
C40654 OR2X1_LOC_790/A AND2X1_LOC_45/a_8_24# 0.05fF
C40655 OR2X1_LOC_394/Y AND2X1_LOC_403/B 0.01fF
C40656 OR2X1_LOC_147/a_8_216# AND2X1_LOC_41/A 0.01fF
C40657 OR2X1_LOC_176/Y AND2X1_LOC_170/B 0.02fF
C40658 OR2X1_LOC_160/B AND2X1_LOC_51/Y 4.48fF
C40659 OR2X1_LOC_485/A OR2X1_LOC_597/a_8_216# 0.01fF
C40660 AND2X1_LOC_773/Y AND2X1_LOC_831/Y 0.21fF
C40661 OR2X1_LOC_272/a_8_216# OR2X1_LOC_59/Y 0.01fF
C40662 OR2X1_LOC_6/B OR2X1_LOC_656/a_36_216# 0.02fF
C40663 OR2X1_LOC_774/Y OR2X1_LOC_859/a_8_216# 0.01fF
C40664 OR2X1_LOC_680/A OR2X1_LOC_427/A 0.07fF
C40665 AND2X1_LOC_95/Y AND2X1_LOC_43/B 0.14fF
C40666 OR2X1_LOC_404/Y OR2X1_LOC_66/A 0.49fF
C40667 OR2X1_LOC_43/A OR2X1_LOC_426/A 0.30fF
C40668 OR2X1_LOC_633/a_36_216# OR2X1_LOC_633/B 0.02fF
C40669 OR2X1_LOC_65/B OR2X1_LOC_118/Y 0.04fF
C40670 AND2X1_LOC_453/Y AND2X1_LOC_452/Y 0.03fF
C40671 OR2X1_LOC_160/A OR2X1_LOC_803/B 0.01fF
C40672 OR2X1_LOC_185/A OR2X1_LOC_254/B 0.64fF
C40673 OR2X1_LOC_471/Y OR2X1_LOC_726/A 0.99fF
C40674 OR2X1_LOC_669/A OR2X1_LOC_278/Y 0.01fF
C40675 OR2X1_LOC_160/B OR2X1_LOC_849/a_8_216# 0.01fF
C40676 OR2X1_LOC_479/Y OR2X1_LOC_147/A 0.03fF
C40677 OR2X1_LOC_70/Y INPUT_0 0.02fF
C40678 AND2X1_LOC_170/B AND2X1_LOC_212/Y 0.02fF
C40679 OR2X1_LOC_62/B OR2X1_LOC_631/A 0.00fF
C40680 OR2X1_LOC_161/A OR2X1_LOC_553/A 0.14fF
C40681 OR2X1_LOC_409/B AND2X1_LOC_771/a_36_24# 0.00fF
C40682 OR2X1_LOC_140/B OR2X1_LOC_493/Y 0.03fF
C40683 OR2X1_LOC_291/A OR2X1_LOC_234/Y 0.03fF
C40684 AND2X1_LOC_56/B OR2X1_LOC_220/B 0.03fF
C40685 AND2X1_LOC_348/A AND2X1_LOC_294/a_8_24# 0.02fF
C40686 OR2X1_LOC_394/Y OR2X1_LOC_44/Y 0.06fF
C40687 D_INPUT_3 OR2X1_LOC_12/Y 0.23fF
C40688 OR2X1_LOC_64/Y OR2X1_LOC_59/Y 5.89fF
C40689 OR2X1_LOC_599/A AND2X1_LOC_644/Y 0.02fF
C40690 OR2X1_LOC_798/a_8_216# OR2X1_LOC_539/Y 0.01fF
C40691 AND2X1_LOC_12/Y OR2X1_LOC_194/Y 0.01fF
C40692 AND2X1_LOC_39/a_36_24# OR2X1_LOC_155/A 0.00fF
C40693 OR2X1_LOC_161/A OR2X1_LOC_779/a_36_216# 0.01fF
C40694 AND2X1_LOC_753/B OR2X1_LOC_654/A 0.01fF
C40695 OR2X1_LOC_51/Y AND2X1_LOC_687/B 0.03fF
C40696 OR2X1_LOC_619/Y OR2X1_LOC_601/Y 0.03fF
C40697 OR2X1_LOC_715/B AND2X1_LOC_47/Y 0.14fF
C40698 OR2X1_LOC_6/A OR2X1_LOC_39/A 0.04fF
C40699 OR2X1_LOC_599/A OR2X1_LOC_424/a_8_216# 0.01fF
C40700 OR2X1_LOC_68/B OR2X1_LOC_333/A 0.17fF
C40701 AND2X1_LOC_215/Y INPUT_1 0.00fF
C40702 OR2X1_LOC_643/Y AND2X1_LOC_92/Y 0.03fF
C40703 AND2X1_LOC_56/B OR2X1_LOC_828/B 0.03fF
C40704 AND2X1_LOC_514/Y INPUT_0 0.03fF
C40705 AND2X1_LOC_348/A AND2X1_LOC_345/Y 0.01fF
C40706 OR2X1_LOC_810/A OR2X1_LOC_506/A 0.01fF
C40707 OR2X1_LOC_158/A OR2X1_LOC_62/A 0.08fF
C40708 OR2X1_LOC_799/A OR2X1_LOC_155/A 0.72fF
C40709 AND2X1_LOC_858/B AND2X1_LOC_465/Y 0.04fF
C40710 OR2X1_LOC_364/A OR2X1_LOC_653/A 0.09fF
C40711 OR2X1_LOC_262/Y OR2X1_LOC_65/B 0.08fF
C40712 OR2X1_LOC_40/Y AND2X1_LOC_866/A 0.22fF
C40713 OR2X1_LOC_185/Y OR2X1_LOC_653/A 0.03fF
C40714 AND2X1_LOC_538/a_8_24# INPUT_0 0.01fF
C40715 OR2X1_LOC_74/A AND2X1_LOC_805/Y 0.08fF
C40716 OR2X1_LOC_62/B OR2X1_LOC_632/Y 0.13fF
C40717 AND2X1_LOC_286/Y AND2X1_LOC_288/a_8_24# 0.03fF
C40718 AND2X1_LOC_723/a_36_24# OR2X1_LOC_74/A 0.01fF
C40719 OR2X1_LOC_7/A AND2X1_LOC_454/Y 0.01fF
C40720 D_INPUT_0 AND2X1_LOC_232/a_8_24# -0.00fF
C40721 OR2X1_LOC_474/a_8_216# OR2X1_LOC_474/Y 0.02fF
C40722 AND2X1_LOC_8/Y OR2X1_LOC_204/Y 0.01fF
C40723 OR2X1_LOC_516/B AND2X1_LOC_727/A 0.02fF
C40724 OR2X1_LOC_794/a_8_216# OR2X1_LOC_161/A 0.01fF
C40725 OR2X1_LOC_36/Y AND2X1_LOC_852/Y 0.06fF
C40726 AND2X1_LOC_109/a_8_24# AND2X1_LOC_18/Y 0.01fF
C40727 OR2X1_LOC_417/A OR2X1_LOC_59/Y 0.30fF
C40728 OR2X1_LOC_177/Y AND2X1_LOC_795/Y 0.02fF
C40729 OR2X1_LOC_753/a_8_216# OR2X1_LOC_753/Y 0.01fF
C40730 AND2X1_LOC_154/a_8_24# AND2X1_LOC_154/Y 0.01fF
C40731 OR2X1_LOC_54/Y AND2X1_LOC_839/a_8_24# 0.02fF
C40732 OR2X1_LOC_392/B OR2X1_LOC_68/B 0.01fF
C40733 AND2X1_LOC_211/B OR2X1_LOC_6/A 0.02fF
C40734 OR2X1_LOC_409/B AND2X1_LOC_637/a_8_24# 0.01fF
C40735 AND2X1_LOC_12/Y OR2X1_LOC_201/Y 0.13fF
C40736 AND2X1_LOC_696/a_8_24# OR2X1_LOC_708/B 0.01fF
C40737 OR2X1_LOC_599/A OR2X1_LOC_7/A 0.06fF
C40738 OR2X1_LOC_604/A OR2X1_LOC_430/Y 0.02fF
C40739 AND2X1_LOC_675/Y OR2X1_LOC_95/Y 0.52fF
C40740 OR2X1_LOC_46/A OR2X1_LOC_46/a_8_216# 0.01fF
C40741 OR2X1_LOC_264/Y OR2X1_LOC_814/A 0.06fF
C40742 AND2X1_LOC_656/a_8_24# OR2X1_LOC_12/Y 0.01fF
C40743 OR2X1_LOC_436/B OR2X1_LOC_814/A 0.02fF
C40744 OR2X1_LOC_124/a_36_216# OR2X1_LOC_786/Y 0.00fF
C40745 OR2X1_LOC_280/Y OR2X1_LOC_44/Y 0.00fF
C40746 AND2X1_LOC_64/a_8_24# AND2X1_LOC_21/Y 0.13fF
C40747 AND2X1_LOC_1/Y AND2X1_LOC_47/a_8_24# 0.01fF
C40748 AND2X1_LOC_170/a_8_24# OR2X1_LOC_417/Y 0.01fF
C40749 OR2X1_LOC_864/A AND2X1_LOC_3/Y 0.06fF
C40750 OR2X1_LOC_533/Y OR2X1_LOC_331/Y 0.16fF
C40751 OR2X1_LOC_631/B OR2X1_LOC_629/A 0.16fF
C40752 OR2X1_LOC_8/Y AND2X1_LOC_838/B 0.01fF
C40753 OR2X1_LOC_93/a_8_216# OR2X1_LOC_7/A 0.39fF
C40754 AND2X1_LOC_173/a_8_24# D_INPUT_0 0.01fF
C40755 OR2X1_LOC_715/B OR2X1_LOC_598/A 0.08fF
C40756 VDD OR2X1_LOC_599/Y 0.04fF
C40757 AND2X1_LOC_40/Y OR2X1_LOC_434/A 0.01fF
C40758 OR2X1_LOC_786/Y AND2X1_LOC_92/Y 0.02fF
C40759 AND2X1_LOC_54/a_8_24# D_INPUT_3 0.01fF
C40760 OR2X1_LOC_442/a_8_216# AND2X1_LOC_804/Y 0.01fF
C40761 OR2X1_LOC_831/a_36_216# AND2X1_LOC_51/Y 0.02fF
C40762 OR2X1_LOC_756/B AND2X1_LOC_250/a_8_24# 0.02fF
C40763 OR2X1_LOC_45/Y AND2X1_LOC_196/Y 0.00fF
C40764 AND2X1_LOC_41/A OR2X1_LOC_473/A 0.05fF
C40765 OR2X1_LOC_154/A OR2X1_LOC_476/a_8_216# 0.02fF
C40766 OR2X1_LOC_6/B OR2X1_LOC_749/a_8_216# 0.06fF
C40767 OR2X1_LOC_6/B OR2X1_LOC_398/Y 0.01fF
C40768 OR2X1_LOC_160/A OR2X1_LOC_520/A 0.02fF
C40769 OR2X1_LOC_243/A OR2X1_LOC_243/B 0.16fF
C40770 AND2X1_LOC_44/Y OR2X1_LOC_550/B 0.03fF
C40771 OR2X1_LOC_22/Y OR2X1_LOC_44/Y 0.83fF
C40772 OR2X1_LOC_613/Y AND2X1_LOC_629/Y 0.14fF
C40773 OR2X1_LOC_139/A OR2X1_LOC_174/Y 0.03fF
C40774 OR2X1_LOC_13/B AND2X1_LOC_774/A 0.74fF
C40775 AND2X1_LOC_839/B OR2X1_LOC_54/Y 0.00fF
C40776 OR2X1_LOC_62/A OR2X1_LOC_847/A 0.02fF
C40777 AND2X1_LOC_714/B OR2X1_LOC_423/Y 0.01fF
C40778 AND2X1_LOC_113/a_36_24# OR2X1_LOC_47/Y 0.00fF
C40779 OR2X1_LOC_479/Y OR2X1_LOC_470/B 0.00fF
C40780 OR2X1_LOC_76/A OR2X1_LOC_787/Y 0.01fF
C40781 AND2X1_LOC_12/Y OR2X1_LOC_201/a_8_216# 0.05fF
C40782 OR2X1_LOC_502/a_36_216# OR2X1_LOC_502/Y 0.00fF
C40783 OR2X1_LOC_216/A OR2X1_LOC_66/Y 0.75fF
C40784 OR2X1_LOC_778/Y OR2X1_LOC_814/A 0.10fF
C40785 OR2X1_LOC_477/B OR2X1_LOC_471/Y 0.03fF
C40786 AND2X1_LOC_561/B AND2X1_LOC_657/A 0.09fF
C40787 OR2X1_LOC_189/A OR2X1_LOC_95/Y 0.11fF
C40788 OR2X1_LOC_788/B OR2X1_LOC_356/A 0.04fF
C40789 OR2X1_LOC_70/Y OR2X1_LOC_64/Y 0.34fF
C40790 D_INPUT_0 OR2X1_LOC_24/a_8_216# 0.01fF
C40791 INPUT_0 AND2X1_LOC_31/Y 0.07fF
C40792 OR2X1_LOC_291/A OR2X1_LOC_278/A 0.19fF
C40793 OR2X1_LOC_218/Y OR2X1_LOC_87/A 0.02fF
C40794 OR2X1_LOC_41/a_8_216# OR2X1_LOC_48/B 0.03fF
C40795 OR2X1_LOC_685/A AND2X1_LOC_681/a_8_24# 0.20fF
C40796 AND2X1_LOC_41/A OR2X1_LOC_228/Y 0.51fF
C40797 AND2X1_LOC_529/a_8_24# OR2X1_LOC_68/B 0.01fF
C40798 OR2X1_LOC_678/Y OR2X1_LOC_513/a_36_216# 0.01fF
C40799 OR2X1_LOC_503/A OR2X1_LOC_184/Y 0.00fF
C40800 AND2X1_LOC_191/Y AND2X1_LOC_632/A 0.03fF
C40801 OR2X1_LOC_837/B OR2X1_LOC_598/A 0.03fF
C40802 AND2X1_LOC_64/Y OR2X1_LOC_175/Y 0.26fF
C40803 AND2X1_LOC_41/A OR2X1_LOC_513/Y 0.00fF
C40804 OR2X1_LOC_802/Y OR2X1_LOC_112/B 0.06fF
C40805 OR2X1_LOC_252/Y AND2X1_LOC_624/B 0.01fF
C40806 AND2X1_LOC_514/Y OR2X1_LOC_64/Y 0.02fF
C40807 AND2X1_LOC_711/Y AND2X1_LOC_632/A 0.03fF
C40808 AND2X1_LOC_811/Y OR2X1_LOC_52/B 0.65fF
C40809 AND2X1_LOC_680/a_36_24# AND2X1_LOC_51/Y 0.00fF
C40810 OR2X1_LOC_411/a_8_216# OR2X1_LOC_585/A 0.06fF
C40811 OR2X1_LOC_276/A AND2X1_LOC_495/a_8_24# 0.20fF
C40812 OR2X1_LOC_177/Y AND2X1_LOC_439/a_8_24# 0.01fF
C40813 OR2X1_LOC_78/A OR2X1_LOC_446/B 0.03fF
C40814 AND2X1_LOC_31/Y OR2X1_LOC_775/a_8_216# 0.01fF
C40815 AND2X1_LOC_12/Y OR2X1_LOC_544/a_8_216# 0.06fF
C40816 OR2X1_LOC_479/Y OR2X1_LOC_532/B 0.06fF
C40817 AND2X1_LOC_866/A OR2X1_LOC_7/A 0.20fF
C40818 AND2X1_LOC_81/B OR2X1_LOC_205/Y 0.03fF
C40819 OR2X1_LOC_574/A OR2X1_LOC_241/Y 0.10fF
C40820 OR2X1_LOC_78/A OR2X1_LOC_303/B 0.07fF
C40821 AND2X1_LOC_64/Y OR2X1_LOC_691/Y 0.06fF
C40822 OR2X1_LOC_600/A OR2X1_LOC_142/Y 0.03fF
C40823 OR2X1_LOC_47/Y AND2X1_LOC_610/a_8_24# 0.04fF
C40824 OR2X1_LOC_12/Y OR2X1_LOC_171/Y 0.03fF
C40825 OR2X1_LOC_218/Y OR2X1_LOC_216/a_8_216# 0.00fF
C40826 OR2X1_LOC_36/Y AND2X1_LOC_647/B 0.07fF
C40827 OR2X1_LOC_653/B OR2X1_LOC_390/B 0.05fF
C40828 OR2X1_LOC_599/A OR2X1_LOC_511/a_8_216# 0.02fF
C40829 OR2X1_LOC_160/A OR2X1_LOC_728/B 0.10fF
C40830 OR2X1_LOC_280/a_8_216# OR2X1_LOC_47/Y 0.08fF
C40831 OR2X1_LOC_810/A D_INPUT_1 0.07fF
C40832 OR2X1_LOC_391/A OR2X1_LOC_558/a_8_216# 0.03fF
C40833 OR2X1_LOC_700/a_8_216# AND2X1_LOC_789/Y 0.02fF
C40834 OR2X1_LOC_130/A OR2X1_LOC_358/A 0.01fF
C40835 AND2X1_LOC_140/a_36_24# OR2X1_LOC_95/Y 0.01fF
C40836 OR2X1_LOC_11/Y OR2X1_LOC_70/A 1.07fF
C40837 AND2X1_LOC_599/a_8_24# OR2X1_LOC_691/Y 0.01fF
C40838 AND2X1_LOC_813/a_36_24# AND2X1_LOC_79/Y 0.01fF
C40839 OR2X1_LOC_864/a_8_216# D_INPUT_1 0.01fF
C40840 OR2X1_LOC_311/Y AND2X1_LOC_801/B 0.00fF
C40841 AND2X1_LOC_514/Y OR2X1_LOC_417/A 0.01fF
C40842 AND2X1_LOC_278/a_8_24# OR2X1_LOC_80/A 0.17fF
C40843 OR2X1_LOC_756/B OR2X1_LOC_349/B 0.20fF
C40844 OR2X1_LOC_45/B AND2X1_LOC_774/a_8_24# 0.01fF
C40845 OR2X1_LOC_377/A OR2X1_LOC_80/A 12.76fF
C40846 AND2X1_LOC_72/a_8_24# AND2X1_LOC_72/B 0.11fF
C40847 AND2X1_LOC_81/a_8_24# OR2X1_LOC_598/A 0.02fF
C40848 OR2X1_LOC_161/B OR2X1_LOC_578/a_36_216# 0.02fF
C40849 OR2X1_LOC_89/A AND2X1_LOC_793/Y 0.50fF
C40850 AND2X1_LOC_95/Y OR2X1_LOC_367/B 0.05fF
C40851 OR2X1_LOC_161/B OR2X1_LOC_160/Y 0.02fF
C40852 OR2X1_LOC_95/Y OR2X1_LOC_77/a_8_216# 0.01fF
C40853 AND2X1_LOC_392/A OR2X1_LOC_134/Y 0.03fF
C40854 OR2X1_LOC_258/Y OR2X1_LOC_257/Y 0.04fF
C40855 OR2X1_LOC_119/a_8_216# D_INPUT_1 0.02fF
C40856 OR2X1_LOC_64/Y OR2X1_LOC_184/Y 0.04fF
C40857 OR2X1_LOC_85/A OR2X1_LOC_80/A 0.09fF
C40858 OR2X1_LOC_178/a_36_216# AND2X1_LOC_465/A 0.00fF
C40859 OR2X1_LOC_124/A AND2X1_LOC_64/Y 0.04fF
C40860 OR2X1_LOC_502/A AND2X1_LOC_36/Y 0.99fF
C40861 OR2X1_LOC_610/Y OR2X1_LOC_68/B 0.02fF
C40862 AND2X1_LOC_388/Y OR2X1_LOC_16/A 0.02fF
C40863 OR2X1_LOC_177/Y AND2X1_LOC_542/a_8_24# 0.00fF
C40864 AND2X1_LOC_64/Y OR2X1_LOC_242/a_8_216# 0.01fF
C40865 AND2X1_LOC_564/B AND2X1_LOC_657/Y 0.10fF
C40866 OR2X1_LOC_449/B OR2X1_LOC_724/A 0.87fF
C40867 OR2X1_LOC_357/a_36_216# OR2X1_LOC_182/B 0.00fF
C40868 AND2X1_LOC_799/a_36_24# AND2X1_LOC_436/Y 0.00fF
C40869 AND2X1_LOC_181/a_8_24# AND2X1_LOC_465/A 0.01fF
C40870 AND2X1_LOC_43/B AND2X1_LOC_41/Y 0.05fF
C40871 OR2X1_LOC_426/B OR2X1_LOC_310/a_8_216# 0.02fF
C40872 AND2X1_LOC_318/Y OR2X1_LOC_31/Y 0.16fF
C40873 OR2X1_LOC_858/A AND2X1_LOC_7/B 0.02fF
C40874 AND2X1_LOC_541/Y AND2X1_LOC_361/a_8_24# 0.04fF
C40875 AND2X1_LOC_475/Y AND2X1_LOC_479/a_8_24# 0.09fF
C40876 OR2X1_LOC_270/a_8_216# D_GATE_366 0.01fF
C40877 OR2X1_LOC_64/Y OR2X1_LOC_70/A 0.00fF
C40878 OR2X1_LOC_184/Y OR2X1_LOC_417/A 0.10fF
C40879 OR2X1_LOC_255/a_8_216# AND2X1_LOC_721/A 0.01fF
C40880 OR2X1_LOC_155/A OR2X1_LOC_446/B 7.07fF
C40881 OR2X1_LOC_9/Y OR2X1_LOC_604/A 0.04fF
C40882 OR2X1_LOC_186/Y OR2X1_LOC_809/B 0.11fF
C40883 OR2X1_LOC_135/Y OR2X1_LOC_56/A 0.10fF
C40884 VDD AND2X1_LOC_475/Y 0.21fF
C40885 AND2X1_LOC_456/B AND2X1_LOC_287/B 0.00fF
C40886 OR2X1_LOC_97/A OR2X1_LOC_756/B 0.01fF
C40887 AND2X1_LOC_64/Y OR2X1_LOC_629/Y 0.19fF
C40888 OR2X1_LOC_400/A AND2X1_LOC_36/Y 0.00fF
C40889 OR2X1_LOC_8/Y OR2X1_LOC_158/A 0.02fF
C40890 AND2X1_LOC_347/B OR2X1_LOC_600/A 0.03fF
C40891 AND2X1_LOC_456/B OR2X1_LOC_816/A 1.23fF
C40892 OR2X1_LOC_161/A OR2X1_LOC_354/a_8_216# 0.03fF
C40893 AND2X1_LOC_749/a_8_24# AND2X1_LOC_7/B 0.01fF
C40894 AND2X1_LOC_571/B AND2X1_LOC_573/A 0.03fF
C40895 OR2X1_LOC_362/A OR2X1_LOC_66/A 0.03fF
C40896 OR2X1_LOC_851/B AND2X1_LOC_310/a_8_24# 0.27fF
C40897 OR2X1_LOC_446/a_36_216# OR2X1_LOC_446/B 0.03fF
C40898 OR2X1_LOC_744/A OR2X1_LOC_829/A 0.03fF
C40899 AND2X1_LOC_845/a_8_24# OR2X1_LOC_95/Y 0.03fF
C40900 AND2X1_LOC_512/Y AND2X1_LOC_802/Y 0.07fF
C40901 OR2X1_LOC_605/A OR2X1_LOC_303/B 0.18fF
C40902 OR2X1_LOC_121/B OR2X1_LOC_724/A 0.07fF
C40903 OR2X1_LOC_798/a_8_216# OR2X1_LOC_319/Y 0.07fF
C40904 OR2X1_LOC_78/A OR2X1_LOC_719/B 0.03fF
C40905 OR2X1_LOC_448/A AND2X1_LOC_44/Y 0.00fF
C40906 OR2X1_LOC_22/Y AND2X1_LOC_570/a_8_24# 0.05fF
C40907 AND2X1_LOC_543/Y OR2X1_LOC_109/Y 0.04fF
C40908 OR2X1_LOC_292/a_8_216# OR2X1_LOC_281/Y 0.39fF
C40909 OR2X1_LOC_92/Y AND2X1_LOC_407/a_8_24# 0.04fF
C40910 AND2X1_LOC_95/Y AND2X1_LOC_416/a_8_24# 0.17fF
C40911 OR2X1_LOC_469/a_8_216# OR2X1_LOC_308/Y 0.03fF
C40912 AND2X1_LOC_711/a_8_24# AND2X1_LOC_347/B 0.05fF
C40913 OR2X1_LOC_61/A OR2X1_LOC_61/a_8_216# 0.47fF
C40914 OR2X1_LOC_517/A OR2X1_LOC_595/A 0.25fF
C40915 OR2X1_LOC_756/B D_GATE_662 0.02fF
C40916 OR2X1_LOC_521/Y OR2X1_LOC_428/A 0.02fF
C40917 OR2X1_LOC_440/A OR2X1_LOC_318/B 0.03fF
C40918 OR2X1_LOC_600/A AND2X1_LOC_338/a_8_24# 0.02fF
C40919 AND2X1_LOC_535/Y OR2X1_LOC_329/B 0.03fF
C40920 OR2X1_LOC_512/A OR2X1_LOC_713/A 0.02fF
C40921 VDD AND2X1_LOC_561/B 0.02fF
C40922 OR2X1_LOC_160/A OR2X1_LOC_338/A 0.07fF
C40923 AND2X1_LOC_523/Y OR2X1_LOC_437/A 0.65fF
C40924 OR2X1_LOC_64/a_8_216# OR2X1_LOC_70/A 0.07fF
C40925 OR2X1_LOC_3/B OR2X1_LOC_31/a_8_216# 0.06fF
C40926 AND2X1_LOC_47/Y OR2X1_LOC_398/Y 0.01fF
C40927 AND2X1_LOC_191/B AND2X1_LOC_709/a_36_24# 0.01fF
C40928 OR2X1_LOC_866/B OR2X1_LOC_846/a_8_216# 0.03fF
C40929 OR2X1_LOC_532/B OR2X1_LOC_68/B 0.13fF
C40930 OR2X1_LOC_427/A AND2X1_LOC_407/a_36_24# 0.01fF
C40931 OR2X1_LOC_542/B OR2X1_LOC_78/A 0.04fF
C40932 AND2X1_LOC_650/Y OR2X1_LOC_171/Y 0.08fF
C40933 OR2X1_LOC_203/Y OR2X1_LOC_115/B 0.07fF
C40934 OR2X1_LOC_426/B AND2X1_LOC_434/Y 0.08fF
C40935 AND2X1_LOC_22/Y AND2X1_LOC_43/B 0.42fF
C40936 OR2X1_LOC_426/B AND2X1_LOC_219/Y 0.13fF
C40937 OR2X1_LOC_615/Y OR2X1_LOC_753/Y 0.00fF
C40938 AND2X1_LOC_70/Y AND2X1_LOC_164/a_8_24# 0.01fF
C40939 AND2X1_LOC_22/Y AND2X1_LOC_132/a_36_24# 0.01fF
C40940 OR2X1_LOC_118/a_36_216# OR2X1_LOC_118/Y 0.00fF
C40941 AND2X1_LOC_486/Y AND2X1_LOC_719/Y 0.10fF
C40942 VDD AND2X1_LOC_197/Y 0.02fF
C40943 OR2X1_LOC_8/Y AND2X1_LOC_98/Y 0.23fF
C40944 AND2X1_LOC_211/B OR2X1_LOC_171/a_36_216# 0.00fF
C40945 AND2X1_LOC_773/Y AND2X1_LOC_139/B 0.41fF
C40946 OR2X1_LOC_158/A AND2X1_LOC_76/Y 0.04fF
C40947 OR2X1_LOC_494/A AND2X1_LOC_359/B 0.00fF
C40948 OR2X1_LOC_186/Y OR2X1_LOC_160/A 0.05fF
C40949 AND2X1_LOC_510/a_8_24# AND2X1_LOC_510/A 0.03fF
C40950 OR2X1_LOC_323/A AND2X1_LOC_458/a_36_24# 0.00fF
C40951 OR2X1_LOC_474/Y OR2X1_LOC_66/A 0.03fF
C40952 OR2X1_LOC_485/Y OR2X1_LOC_485/a_8_216# 0.01fF
C40953 OR2X1_LOC_343/B OR2X1_LOC_68/B 0.03fF
C40954 OR2X1_LOC_535/A AND2X1_LOC_166/a_8_24# 0.08fF
C40955 AND2X1_LOC_510/a_36_24# AND2X1_LOC_658/A 0.01fF
C40956 AND2X1_LOC_727/Y OR2X1_LOC_189/Y 0.03fF
C40957 OR2X1_LOC_314/a_36_216# OR2X1_LOC_604/A 0.00fF
C40958 OR2X1_LOC_451/B AND2X1_LOC_428/a_36_24# 0.00fF
C40959 AND2X1_LOC_59/Y OR2X1_LOC_294/Y 0.31fF
C40960 AND2X1_LOC_787/A OR2X1_LOC_91/a_8_216# 0.01fF
C40961 OR2X1_LOC_176/Y AND2X1_LOC_170/Y 0.25fF
C40962 OR2X1_LOC_539/A OR2X1_LOC_66/A 0.03fF
C40963 OR2X1_LOC_49/A AND2X1_LOC_80/a_36_24# 0.01fF
C40964 OR2X1_LOC_151/A OR2X1_LOC_624/A 0.08fF
C40965 OR2X1_LOC_109/Y OR2X1_LOC_322/Y 0.48fF
C40966 AND2X1_LOC_753/B VDD 0.15fF
C40967 AND2X1_LOC_452/Y AND2X1_LOC_605/a_8_24# 0.02fF
C40968 OR2X1_LOC_49/A OR2X1_LOC_87/A 0.71fF
C40969 AND2X1_LOC_319/A AND2X1_LOC_809/a_8_24# 0.13fF
C40970 AND2X1_LOC_40/Y OR2X1_LOC_741/Y 1.73fF
C40971 AND2X1_LOC_50/Y AND2X1_LOC_70/Y 0.05fF
C40972 AND2X1_LOC_778/a_8_24# AND2X1_LOC_721/Y 0.01fF
C40973 AND2X1_LOC_727/Y OR2X1_LOC_152/Y 0.01fF
C40974 OR2X1_LOC_656/B OR2X1_LOC_6/B 0.10fF
C40975 OR2X1_LOC_105/a_8_216# OR2X1_LOC_78/A 0.02fF
C40976 OR2X1_LOC_347/a_8_216# VDD 0.00fF
C40977 AND2X1_LOC_48/A AND2X1_LOC_36/Y 0.59fF
C40978 AND2X1_LOC_445/a_36_24# OR2X1_LOC_44/Y 0.01fF
C40979 OR2X1_LOC_405/A OR2X1_LOC_723/a_36_216# 0.01fF
C40980 OR2X1_LOC_438/Y AND2X1_LOC_663/A 0.03fF
C40981 AND2X1_LOC_810/A AND2X1_LOC_661/A 0.02fF
C40982 AND2X1_LOC_805/Y OR2X1_LOC_626/Y 0.46fF
C40983 OR2X1_LOC_797/B OR2X1_LOC_209/a_8_216# 0.08fF
C40984 OR2X1_LOC_693/a_8_216# OR2X1_LOC_36/Y 0.08fF
C40985 AND2X1_LOC_170/Y AND2X1_LOC_212/Y 0.06fF
C40986 OR2X1_LOC_691/A OR2X1_LOC_269/B 0.02fF
C40987 OR2X1_LOC_170/Y OR2X1_LOC_365/B 0.00fF
C40988 OR2X1_LOC_858/B OR2X1_LOC_756/B 0.01fF
C40989 OR2X1_LOC_348/Y AND2X1_LOC_95/Y 0.07fF
C40990 OR2X1_LOC_405/A VDD 1.35fF
C40991 AND2X1_LOC_544/Y OR2X1_LOC_70/Y 0.01fF
C40992 AND2X1_LOC_776/Y OR2X1_LOC_527/Y 0.91fF
C40993 OR2X1_LOC_33/a_8_216# OR2X1_LOC_338/A 0.01fF
C40994 AND2X1_LOC_59/Y OR2X1_LOC_641/A 0.00fF
C40995 OR2X1_LOC_287/B OR2X1_LOC_576/A 0.12fF
C40996 OR2X1_LOC_840/a_36_216# OR2X1_LOC_87/A 0.00fF
C40997 OR2X1_LOC_8/Y OR2X1_LOC_847/A 0.34fF
C40998 OR2X1_LOC_851/A AND2X1_LOC_92/Y 0.99fF
C40999 OR2X1_LOC_677/a_8_216# OR2X1_LOC_677/Y 0.01fF
C41000 OR2X1_LOC_49/A AND2X1_LOC_19/a_8_24# 0.02fF
C41001 VDD OR2X1_LOC_616/a_8_216# 0.21fF
C41002 OR2X1_LOC_87/A OR2X1_LOC_596/A 0.03fF
C41003 OR2X1_LOC_45/B OR2X1_LOC_280/Y 0.08fF
C41004 AND2X1_LOC_803/B OR2X1_LOC_679/B 0.00fF
C41005 AND2X1_LOC_197/Y AND2X1_LOC_208/B 0.83fF
C41006 VDD OR2X1_LOC_413/Y 0.04fF
C41007 OR2X1_LOC_139/A AND2X1_LOC_42/B 0.00fF
C41008 AND2X1_LOC_704/a_8_24# OR2X1_LOC_418/Y 0.24fF
C41009 OR2X1_LOC_160/B OR2X1_LOC_541/a_8_216# 0.01fF
C41010 AND2X1_LOC_70/a_8_24# AND2X1_LOC_11/Y 0.01fF
C41011 AND2X1_LOC_566/B OR2X1_LOC_36/Y 0.05fF
C41012 OR2X1_LOC_589/A OR2X1_LOC_262/a_8_216# 0.01fF
C41013 OR2X1_LOC_471/a_8_216# OR2X1_LOC_741/Y 0.01fF
C41014 OR2X1_LOC_820/a_8_216# OR2X1_LOC_44/Y 0.01fF
C41015 AND2X1_LOC_219/a_36_24# OR2X1_LOC_619/Y 0.01fF
C41016 OR2X1_LOC_631/a_8_216# OR2X1_LOC_78/A 0.01fF
C41017 D_INPUT_3 OR2X1_LOC_248/A 0.08fF
C41018 OR2X1_LOC_604/A OR2X1_LOC_96/B 0.04fF
C41019 AND2X1_LOC_736/Y OR2X1_LOC_441/Y 0.19fF
C41020 AND2X1_LOC_737/Y OR2X1_LOC_441/a_36_216# 0.00fF
C41021 OR2X1_LOC_158/A OR2X1_LOC_52/B 0.74fF
C41022 OR2X1_LOC_158/A OR2X1_LOC_672/Y 0.01fF
C41023 OR2X1_LOC_3/Y OR2X1_LOC_16/A 0.36fF
C41024 OR2X1_LOC_109/a_8_216# AND2X1_LOC_471/Y 0.02fF
C41025 OR2X1_LOC_485/Y OR2X1_LOC_44/Y 0.00fF
C41026 VDD AND2X1_LOC_266/Y 0.04fF
C41027 AND2X1_LOC_562/Y AND2X1_LOC_563/Y 0.16fF
C41028 OR2X1_LOC_185/Y AND2X1_LOC_131/a_36_24# 0.06fF
C41029 OR2X1_LOC_217/Y OR2X1_LOC_66/A 0.08fF
C41030 AND2X1_LOC_848/Y OR2X1_LOC_56/A 0.07fF
C41031 OR2X1_LOC_858/A OR2X1_LOC_805/A 0.03fF
C41032 AND2X1_LOC_710/Y AND2X1_LOC_848/Y 0.10fF
C41033 OR2X1_LOC_744/A AND2X1_LOC_648/a_8_24# 0.01fF
C41034 OR2X1_LOC_325/a_8_216# OR2X1_LOC_502/A 0.01fF
C41035 OR2X1_LOC_662/A OR2X1_LOC_660/Y 0.01fF
C41036 OR2X1_LOC_491/a_8_216# AND2X1_LOC_717/B 0.00fF
C41037 OR2X1_LOC_124/B OR2X1_LOC_205/a_8_216# 0.10fF
C41038 OR2X1_LOC_158/A AND2X1_LOC_489/Y 0.14fF
C41039 AND2X1_LOC_40/Y OR2X1_LOC_509/A 0.01fF
C41040 AND2X1_LOC_719/Y OR2X1_LOC_666/Y 0.00fF
C41041 OR2X1_LOC_40/Y AND2X1_LOC_857/a_8_24# 0.01fF
C41042 VDD AND2X1_LOC_823/a_8_24# 0.00fF
C41043 AND2X1_LOC_91/B OR2X1_LOC_814/A 0.46fF
C41044 OR2X1_LOC_104/a_8_216# OR2X1_LOC_85/A 0.01fF
C41045 OR2X1_LOC_43/A AND2X1_LOC_447/Y 0.28fF
C41046 OR2X1_LOC_494/Y OR2X1_LOC_26/Y 0.03fF
C41047 AND2X1_LOC_567/a_36_24# AND2X1_LOC_661/A 0.00fF
C41048 OR2X1_LOC_40/Y OR2X1_LOC_7/A 0.21fF
C41049 AND2X1_LOC_456/B AND2X1_LOC_843/a_8_24# 0.01fF
C41050 AND2X1_LOC_716/Y AND2X1_LOC_357/a_36_24# 0.00fF
C41051 OR2X1_LOC_691/B AND2X1_LOC_51/Y 0.00fF
C41052 OR2X1_LOC_833/a_8_216# OR2X1_LOC_833/B 0.08fF
C41053 OR2X1_LOC_264/Y AND2X1_LOC_517/a_8_24# 0.03fF
C41054 OR2X1_LOC_643/A OR2X1_LOC_244/Y 0.02fF
C41055 OR2X1_LOC_706/A AND2X1_LOC_43/B 0.03fF
C41056 OR2X1_LOC_307/B OR2X1_LOC_161/A 0.03fF
C41057 AND2X1_LOC_56/B OR2X1_LOC_78/A 0.09fF
C41058 OR2X1_LOC_298/Y OR2X1_LOC_298/a_8_216# 0.02fF
C41059 OR2X1_LOC_600/A OR2X1_LOC_238/Y 0.03fF
C41060 OR2X1_LOC_623/a_8_216# OR2X1_LOC_623/B 0.08fF
C41061 AND2X1_LOC_533/a_36_24# OR2X1_LOC_703/A 0.00fF
C41062 AND2X1_LOC_141/A AND2X1_LOC_573/A 0.01fF
C41063 OR2X1_LOC_45/B OR2X1_LOC_22/Y 0.40fF
C41064 OR2X1_LOC_160/B OR2X1_LOC_787/Y 0.07fF
C41065 OR2X1_LOC_589/A AND2X1_LOC_729/B 0.08fF
C41066 OR2X1_LOC_756/B AND2X1_LOC_282/a_8_24# 0.02fF
C41067 AND2X1_LOC_597/a_8_24# INPUT_0 0.01fF
C41068 VDD OR2X1_LOC_387/Y 0.16fF
C41069 AND2X1_LOC_350/a_8_24# AND2X1_LOC_350/Y 0.02fF
C41070 INPUT_0 OR2X1_LOC_461/A 0.15fF
C41071 AND2X1_LOC_351/a_8_24# OR2X1_LOC_46/A 0.01fF
C41072 OR2X1_LOC_494/Y OR2X1_LOC_89/A 0.03fF
C41073 AND2X1_LOC_8/Y OR2X1_LOC_78/A 0.18fF
C41074 AND2X1_LOC_363/Y OR2X1_LOC_89/A 0.03fF
C41075 OR2X1_LOC_764/Y OR2X1_LOC_426/B 0.03fF
C41076 AND2X1_LOC_88/a_36_24# AND2X1_LOC_18/Y 0.00fF
C41077 OR2X1_LOC_46/A AND2X1_LOC_415/a_8_24# 0.02fF
C41078 AND2X1_LOC_500/Y OR2X1_LOC_239/Y 0.01fF
C41079 OR2X1_LOC_633/Y OR2X1_LOC_610/a_8_216# 0.03fF
C41080 OR2X1_LOC_808/A OR2X1_LOC_87/A 0.00fF
C41081 AND2X1_LOC_227/Y AND2X1_LOC_242/B 0.19fF
C41082 OR2X1_LOC_395/Y OR2X1_LOC_396/Y 0.11fF
C41083 AND2X1_LOC_7/Y AND2X1_LOC_44/Y 0.02fF
C41084 OR2X1_LOC_51/Y AND2X1_LOC_640/Y 0.03fF
C41085 INPUT_5 AND2X1_LOC_25/Y 0.01fF
C41086 VDD AND2X1_LOC_10/a_8_24# -0.00fF
C41087 AND2X1_LOC_304/a_8_24# OR2X1_LOC_269/B 0.03fF
C41088 OR2X1_LOC_3/Y AND2X1_LOC_121/a_8_24# 0.01fF
C41089 AND2X1_LOC_174/a_8_24# OR2X1_LOC_619/Y 0.09fF
C41090 AND2X1_LOC_349/a_8_24# OR2X1_LOC_92/Y 0.05fF
C41091 OR2X1_LOC_118/Y OR2X1_LOC_619/Y 0.03fF
C41092 OR2X1_LOC_188/Y OR2X1_LOC_276/B 0.01fF
C41093 OR2X1_LOC_858/A OR2X1_LOC_296/Y 0.13fF
C41094 OR2X1_LOC_743/A AND2X1_LOC_434/Y 0.07fF
C41095 OR2X1_LOC_743/A AND2X1_LOC_219/Y 0.08fF
C41096 OR2X1_LOC_329/a_36_216# OR2X1_LOC_22/Y 0.02fF
C41097 OR2X1_LOC_51/Y OR2X1_LOC_681/Y 0.01fF
C41098 OR2X1_LOC_302/a_8_216# OR2X1_LOC_479/Y 0.06fF
C41099 OR2X1_LOC_316/Y OR2X1_LOC_18/Y 0.11fF
C41100 OR2X1_LOC_75/a_8_216# AND2X1_LOC_786/Y 0.03fF
C41101 AND2X1_LOC_331/a_36_24# AND2X1_LOC_56/B 0.01fF
C41102 OR2X1_LOC_160/A OR2X1_LOC_231/a_36_216# 0.01fF
C41103 AND2X1_LOC_38/a_36_24# OR2X1_LOC_78/B 0.01fF
C41104 AND2X1_LOC_831/Y OR2X1_LOC_12/Y 0.10fF
C41105 OR2X1_LOC_616/a_8_216# OR2X1_LOC_616/Y 0.02fF
C41106 OR2X1_LOC_720/a_8_216# OR2X1_LOC_721/Y 0.01fF
C41107 OR2X1_LOC_619/Y AND2X1_LOC_453/a_8_24# 0.01fF
C41108 OR2X1_LOC_26/Y AND2X1_LOC_839/a_8_24# 0.01fF
C41109 AND2X1_LOC_50/Y AND2X1_LOC_17/Y 0.02fF
C41110 AND2X1_LOC_658/A AND2X1_LOC_663/B 0.01fF
C41111 AND2X1_LOC_777/a_8_24# AND2X1_LOC_654/Y 0.04fF
C41112 OR2X1_LOC_864/A OR2X1_LOC_772/B 0.01fF
C41113 OR2X1_LOC_91/Y AND2X1_LOC_468/B 0.01fF
C41114 OR2X1_LOC_520/Y OR2X1_LOC_559/B 0.46fF
C41115 OR2X1_LOC_168/Y OR2X1_LOC_365/B 0.00fF
C41116 AND2X1_LOC_861/B OR2X1_LOC_74/A 0.07fF
C41117 AND2X1_LOC_154/a_8_24# AND2X1_LOC_624/A 0.01fF
C41118 AND2X1_LOC_802/B AND2X1_LOC_810/a_8_24# 0.02fF
C41119 AND2X1_LOC_354/B OR2X1_LOC_48/B 4.07fF
C41120 AND2X1_LOC_359/B OR2X1_LOC_427/A 0.12fF
C41121 OR2X1_LOC_774/Y OR2X1_LOC_772/B 0.04fF
C41122 OR2X1_LOC_88/A OR2X1_LOC_118/Y 0.00fF
C41123 OR2X1_LOC_43/A AND2X1_LOC_649/B 0.07fF
C41124 OR2X1_LOC_811/A OR2X1_LOC_269/B 3.18fF
C41125 OR2X1_LOC_160/A AND2X1_LOC_81/B 0.05fF
C41126 OR2X1_LOC_810/A OR2X1_LOC_737/A 0.10fF
C41127 AND2X1_LOC_464/Y OR2X1_LOC_56/A 0.01fF
C41128 OR2X1_LOC_329/B AND2X1_LOC_327/a_8_24# 0.01fF
C41129 VDD OR2X1_LOC_285/Y 0.00fF
C41130 OR2X1_LOC_837/Y OR2X1_LOC_20/a_36_216# 0.02fF
C41131 AND2X1_LOC_42/B OR2X1_LOC_244/a_8_216# 0.01fF
C41132 AND2X1_LOC_863/A OR2X1_LOC_56/A 0.00fF
C41133 OR2X1_LOC_641/Y OR2X1_LOC_649/a_8_216# 0.40fF
C41134 OR2X1_LOC_317/A OR2X1_LOC_778/Y 0.08fF
C41135 OR2X1_LOC_76/Y OR2X1_LOC_269/a_8_216# 0.18fF
C41136 OR2X1_LOC_47/Y OR2X1_LOC_766/a_8_216# 0.01fF
C41137 OR2X1_LOC_607/a_8_216# OR2X1_LOC_607/A 0.47fF
C41138 OR2X1_LOC_243/B OR2X1_LOC_66/A 0.05fF
C41139 AND2X1_LOC_95/Y AND2X1_LOC_159/a_8_24# 0.01fF
C41140 AND2X1_LOC_357/A AND2X1_LOC_863/Y 0.01fF
C41141 OR2X1_LOC_44/Y OR2X1_LOC_39/A 0.22fF
C41142 AND2X1_LOC_95/Y OR2X1_LOC_810/A 0.08fF
C41143 AND2X1_LOC_533/a_8_24# OR2X1_LOC_269/B 0.03fF
C41144 OR2X1_LOC_113/A OR2X1_LOC_244/Y 0.03fF
C41145 OR2X1_LOC_864/A OR2X1_LOC_489/B 0.09fF
C41146 OR2X1_LOC_824/a_8_216# AND2X1_LOC_852/B 0.50fF
C41147 OR2X1_LOC_246/A AND2X1_LOC_219/Y 0.10fF
C41148 AND2X1_LOC_305/a_8_24# AND2X1_LOC_3/Y 0.10fF
C41149 AND2X1_LOC_843/a_36_24# OR2X1_LOC_26/Y 0.00fF
C41150 OR2X1_LOC_421/A OR2X1_LOC_95/Y 0.00fF
C41151 INPUT_5 AND2X1_LOC_51/Y 0.37fF
C41152 AND2X1_LOC_787/A OR2X1_LOC_419/Y 0.03fF
C41153 OR2X1_LOC_85/A OR2X1_LOC_6/A 0.09fF
C41154 OR2X1_LOC_265/Y AND2X1_LOC_361/A 0.03fF
C41155 AND2X1_LOC_266/Y AND2X1_LOC_267/a_8_24# 0.02fF
C41156 OR2X1_LOC_774/Y OR2X1_LOC_489/B 0.00fF
C41157 AND2X1_LOC_563/A OR2X1_LOC_95/Y 0.01fF
C41158 OR2X1_LOC_185/A OR2X1_LOC_445/a_8_216# 0.14fF
C41159 AND2X1_LOC_654/B AND2X1_LOC_729/B 0.05fF
C41160 OR2X1_LOC_87/A OR2X1_LOC_87/B 0.39fF
C41161 AND2X1_LOC_355/a_8_24# AND2X1_LOC_436/B 0.04fF
C41162 AND2X1_LOC_589/a_8_24# AND2X1_LOC_95/Y 0.03fF
C41163 AND2X1_LOC_148/Y AND2X1_LOC_676/a_8_24# 0.20fF
C41164 AND2X1_LOC_841/B AND2X1_LOC_798/Y 0.03fF
C41165 OR2X1_LOC_83/Y OR2X1_LOC_80/Y 0.54fF
C41166 OR2X1_LOC_235/B D_INPUT_0 0.11fF
C41167 OR2X1_LOC_70/Y AND2X1_LOC_550/A 0.70fF
C41168 OR2X1_LOC_76/A OR2X1_LOC_808/a_36_216# 0.02fF
C41169 AND2X1_LOC_363/A AND2X1_LOC_359/B 0.00fF
C41170 AND2X1_LOC_823/a_8_24# OR2X1_LOC_836/B 0.02fF
C41171 AND2X1_LOC_56/B OR2X1_LOC_155/A 0.26fF
C41172 AND2X1_LOC_31/Y AND2X1_LOC_7/B 0.18fF
C41173 OR2X1_LOC_76/A OR2X1_LOC_733/a_36_216# 0.02fF
C41174 OR2X1_LOC_26/Y AND2X1_LOC_839/B 0.01fF
C41175 AND2X1_LOC_7/B OR2X1_LOC_715/a_8_216# 0.02fF
C41176 OR2X1_LOC_431/Y OR2X1_LOC_48/B 0.39fF
C41177 AND2X1_LOC_211/B OR2X1_LOC_44/Y 1.25fF
C41178 OR2X1_LOC_653/Y OR2X1_LOC_476/B 0.04fF
C41179 OR2X1_LOC_87/B AND2X1_LOC_19/a_8_24# 0.04fF
C41180 AND2X1_LOC_76/Y OR2X1_LOC_275/a_36_216# 0.00fF
C41181 OR2X1_LOC_236/a_36_216# OR2X1_LOC_89/A 0.00fF
C41182 AND2X1_LOC_580/A AND2X1_LOC_548/a_8_24# 0.03fF
C41183 AND2X1_LOC_663/B AND2X1_LOC_847/Y 0.28fF
C41184 VDD OR2X1_LOC_779/Y 0.07fF
C41185 OR2X1_LOC_850/B OR2X1_LOC_286/B 0.03fF
C41186 OR2X1_LOC_809/B OR2X1_LOC_112/B 0.19fF
C41187 OR2X1_LOC_404/a_36_216# AND2X1_LOC_51/Y 0.00fF
C41188 OR2X1_LOC_744/A OR2X1_LOC_224/Y 0.02fF
C41189 VDD OR2X1_LOC_330/a_8_216# 0.00fF
C41190 AND2X1_LOC_586/a_8_24# AND2X1_LOC_48/A 0.01fF
C41191 OR2X1_LOC_844/B OR2X1_LOC_500/a_8_216# 0.08fF
C41192 AND2X1_LOC_70/Y OR2X1_LOC_214/B 0.06fF
C41193 D_INPUT_5 OR2X1_LOC_31/Y 0.03fF
C41194 INPUT_0 OR2X1_LOC_47/Y 0.02fF
C41195 OR2X1_LOC_481/Y OR2X1_LOC_748/A 0.01fF
C41196 OR2X1_LOC_187/a_8_216# AND2X1_LOC_866/A 0.05fF
C41197 AND2X1_LOC_70/Y OR2X1_LOC_241/B 0.07fF
C41198 OR2X1_LOC_22/Y AND2X1_LOC_435/a_8_24# 0.01fF
C41199 AND2X1_LOC_303/A AND2X1_LOC_351/Y 0.07fF
C41200 OR2X1_LOC_70/Y AND2X1_LOC_101/B 0.01fF
C41201 OR2X1_LOC_813/A OR2X1_LOC_278/Y 0.00fF
C41202 OR2X1_LOC_43/A AND2X1_LOC_729/B 0.80fF
C41203 OR2X1_LOC_462/B OR2X1_LOC_462/a_36_216# 0.03fF
C41204 AND2X1_LOC_578/A OR2X1_LOC_312/Y 0.03fF
C41205 AND2X1_LOC_703/Y OR2X1_LOC_423/Y 0.02fF
C41206 OR2X1_LOC_361/a_8_216# OR2X1_LOC_560/A 0.09fF
C41207 AND2X1_LOC_554/B OR2X1_LOC_485/A 0.02fF
C41208 OR2X1_LOC_385/Y AND2X1_LOC_390/B 0.01fF
C41209 OR2X1_LOC_387/Y AND2X1_LOC_389/a_8_24# 0.23fF
C41210 OR2X1_LOC_787/Y OR2X1_LOC_794/a_8_216# 0.02fF
C41211 OR2X1_LOC_426/B OR2X1_LOC_595/Y 0.10fF
C41212 AND2X1_LOC_709/a_36_24# AND2X1_LOC_848/A -0.02fF
C41213 AND2X1_LOC_737/Y AND2X1_LOC_811/Y 0.01fF
C41214 OR2X1_LOC_22/Y OR2X1_LOC_767/a_8_216# 0.02fF
C41215 OR2X1_LOC_375/A AND2X1_LOC_667/a_8_24# 0.01fF
C41216 OR2X1_LOC_472/a_8_216# OR2X1_LOC_472/A 0.02fF
C41217 OR2X1_LOC_686/B AND2X1_LOC_430/B 0.00fF
C41218 OR2X1_LOC_3/Y OR2X1_LOC_273/a_8_216# 0.05fF
C41219 AND2X1_LOC_279/a_8_24# OR2X1_LOC_366/Y 0.03fF
C41220 OR2X1_LOC_848/A OR2X1_LOC_773/a_8_216# 0.02fF
C41221 OR2X1_LOC_13/B AND2X1_LOC_786/Y 0.07fF
C41222 AND2X1_LOC_387/a_8_24# OR2X1_LOC_750/Y 0.25fF
C41223 OR2X1_LOC_488/Y AND2X1_LOC_717/B 0.08fF
C41224 AND2X1_LOC_104/a_36_24# AND2X1_LOC_47/Y 0.00fF
C41225 AND2X1_LOC_717/Y OR2X1_LOC_47/Y 0.03fF
C41226 OR2X1_LOC_479/Y OR2X1_LOC_605/a_36_216# 0.01fF
C41227 AND2X1_LOC_727/A AND2X1_LOC_856/A 0.01fF
C41228 OR2X1_LOC_293/a_8_216# OR2X1_LOC_585/A 0.03fF
C41229 OR2X1_LOC_19/B AND2X1_LOC_234/a_8_24# 0.04fF
C41230 AND2X1_LOC_12/Y OR2X1_LOC_440/A 0.03fF
C41231 OR2X1_LOC_377/A D_INPUT_2 0.10fF
C41232 AND2X1_LOC_817/B OR2X1_LOC_770/a_8_216# 0.01fF
C41233 OR2X1_LOC_648/A OR2X1_LOC_228/Y 0.02fF
C41234 OR2X1_LOC_139/a_8_216# OR2X1_LOC_62/B 0.00fF
C41235 OR2X1_LOC_473/Y OR2X1_LOC_206/a_8_216# 0.01fF
C41236 OR2X1_LOC_186/Y OR2X1_LOC_532/Y 0.04fF
C41237 OR2X1_LOC_117/Y AND2X1_LOC_845/Y 0.08fF
C41238 OR2X1_LOC_207/B AND2X1_LOC_36/Y 0.24fF
C41239 AND2X1_LOC_582/a_36_24# OR2X1_LOC_451/B 0.00fF
C41240 OR2X1_LOC_502/A OR2X1_LOC_196/a_8_216# 0.01fF
C41241 AND2X1_LOC_866/A OR2X1_LOC_236/a_8_216# 0.01fF
C41242 AND2X1_LOC_465/Y OR2X1_LOC_371/Y 0.02fF
C41243 D_INPUT_2 OR2X1_LOC_85/A 0.05fF
C41244 OR2X1_LOC_472/A OR2X1_LOC_839/a_8_216# 0.06fF
C41245 OR2X1_LOC_186/Y OR2X1_LOC_212/B 0.01fF
C41246 AND2X1_LOC_530/a_8_24# AND2X1_LOC_36/Y 0.04fF
C41247 OR2X1_LOC_78/B OR2X1_LOC_80/A 2.46fF
C41248 OR2X1_LOC_47/Y OR2X1_LOC_11/Y 0.23fF
C41249 OR2X1_LOC_391/A OR2X1_LOC_68/B 0.08fF
C41250 OR2X1_LOC_288/A AND2X1_LOC_3/Y 0.08fF
C41251 OR2X1_LOC_485/A OR2X1_LOC_167/Y 0.01fF
C41252 OR2X1_LOC_92/Y OR2X1_LOC_754/Y 0.01fF
C41253 OR2X1_LOC_337/a_36_216# OR2X1_LOC_578/B 0.00fF
C41254 AND2X1_LOC_657/Y OR2X1_LOC_437/A 0.25fF
C41255 OR2X1_LOC_291/Y OR2X1_LOC_278/A 0.83fF
C41256 AND2X1_LOC_84/Y AND2X1_LOC_202/Y 0.00fF
C41257 OR2X1_LOC_160/A OR2X1_LOC_66/Y 0.03fF
C41258 OR2X1_LOC_287/A OR2X1_LOC_366/Y 0.08fF
C41259 AND2X1_LOC_717/B OR2X1_LOC_95/Y 0.09fF
C41260 AND2X1_LOC_191/B OR2X1_LOC_437/A 0.00fF
C41261 OR2X1_LOC_764/Y OR2X1_LOC_409/B 0.01fF
C41262 OR2X1_LOC_841/a_36_216# AND2X1_LOC_31/Y 0.01fF
C41263 AND2X1_LOC_560/B OR2X1_LOC_47/Y 0.35fF
C41264 OR2X1_LOC_224/a_8_216# OR2X1_LOC_7/A 0.01fF
C41265 OR2X1_LOC_71/a_36_216# AND2X1_LOC_647/Y 0.00fF
C41266 OR2X1_LOC_404/A AND2X1_LOC_51/Y 0.21fF
C41267 AND2X1_LOC_469/B OR2X1_LOC_437/A 0.03fF
C41268 OR2X1_LOC_318/Y AND2X1_LOC_31/Y 0.03fF
C41269 AND2X1_LOC_48/A AND2X1_LOC_46/a_36_24# 0.00fF
C41270 OR2X1_LOC_66/A OR2X1_LOC_771/B 0.06fF
C41271 OR2X1_LOC_427/A AND2X1_LOC_790/a_8_24# 0.01fF
C41272 OR2X1_LOC_212/a_8_216# AND2X1_LOC_31/Y 0.05fF
C41273 VDD OR2X1_LOC_268/Y 0.07fF
C41274 OR2X1_LOC_269/B AND2X1_LOC_237/a_8_24# 0.01fF
C41275 AND2X1_LOC_733/Y OR2X1_LOC_437/A 0.07fF
C41276 VDD OR2X1_LOC_183/Y 0.14fF
C41277 OR2X1_LOC_87/A OR2X1_LOC_374/Y 0.15fF
C41278 AND2X1_LOC_461/a_8_24# OR2X1_LOC_690/A 0.16fF
C41279 INPUT_1 OR2X1_LOC_54/Y 0.25fF
C41280 AND2X1_LOC_348/A OR2X1_LOC_384/Y 0.01fF
C41281 OR2X1_LOC_813/A OR2X1_LOC_19/B 0.01fF
C41282 OR2X1_LOC_825/Y OR2X1_LOC_95/Y 0.09fF
C41283 OR2X1_LOC_26/Y OR2X1_LOC_311/a_8_216# 0.07fF
C41284 OR2X1_LOC_841/A OR2X1_LOC_776/A 0.16fF
C41285 OR2X1_LOC_805/A AND2X1_LOC_31/Y 0.23fF
C41286 AND2X1_LOC_44/Y OR2X1_LOC_706/a_8_216# 0.01fF
C41287 AND2X1_LOC_605/Y AND2X1_LOC_449/a_8_24# 0.11fF
C41288 AND2X1_LOC_748/a_36_24# OR2X1_LOC_789/A 0.00fF
C41289 OR2X1_LOC_428/A AND2X1_LOC_774/A 0.38fF
C41290 OR2X1_LOC_468/A OR2X1_LOC_168/Y 0.03fF
C41291 AND2X1_LOC_3/Y AND2X1_LOC_72/B 0.03fF
C41292 OR2X1_LOC_778/Y OR2X1_LOC_318/B 0.05fF
C41293 OR2X1_LOC_177/Y AND2X1_LOC_787/A 0.63fF
C41294 OR2X1_LOC_243/a_8_216# OR2X1_LOC_244/A 0.05fF
C41295 OR2X1_LOC_691/Y OR2X1_LOC_185/a_8_216# 0.01fF
C41296 AND2X1_LOC_3/Y OR2X1_LOC_451/B 0.24fF
C41297 OR2X1_LOC_375/A OR2X1_LOC_80/A 0.03fF
C41298 OR2X1_LOC_49/A OR2X1_LOC_381/a_8_216# 0.01fF
C41299 OR2X1_LOC_64/Y OR2X1_LOC_47/Y 1.11fF
C41300 OR2X1_LOC_743/A OR2X1_LOC_595/Y 0.52fF
C41301 AND2X1_LOC_573/A OR2X1_LOC_399/a_36_216# 0.00fF
C41302 AND2X1_LOC_544/Y AND2X1_LOC_658/B 0.03fF
C41303 AND2X1_LOC_91/B OR2X1_LOC_244/Y 0.05fF
C41304 OR2X1_LOC_158/A OR2X1_LOC_9/a_8_216# 0.15fF
C41305 AND2X1_LOC_787/A OR2X1_LOC_604/A 0.01fF
C41306 OR2X1_LOC_833/Y OR2X1_LOC_851/B 0.02fF
C41307 OR2X1_LOC_276/B D_INPUT_0 0.48fF
C41308 OR2X1_LOC_571/B OR2X1_LOC_571/Y 0.01fF
C41309 OR2X1_LOC_155/A AND2X1_LOC_427/a_8_24# 0.01fF
C41310 OR2X1_LOC_739/A OR2X1_LOC_777/B 0.02fF
C41311 OR2X1_LOC_160/B OR2X1_LOC_576/A 0.07fF
C41312 OR2X1_LOC_507/a_36_216# OR2X1_LOC_508/Y 0.00fF
C41313 OR2X1_LOC_188/Y AND2X1_LOC_70/Y 0.08fF
C41314 OR2X1_LOC_158/A OR2X1_LOC_281/Y 0.01fF
C41315 OR2X1_LOC_151/A OR2X1_LOC_346/A 0.01fF
C41316 OR2X1_LOC_624/A OR2X1_LOC_332/a_36_216# 0.16fF
C41317 AND2X1_LOC_713/Y OR2X1_LOC_12/Y 0.00fF
C41318 AND2X1_LOC_574/Y AND2X1_LOC_675/Y 0.05fF
C41319 OR2X1_LOC_161/A AND2X1_LOC_246/a_8_24# 0.00fF
C41320 OR2X1_LOC_12/Y AND2X1_LOC_448/a_36_24# 0.00fF
C41321 OR2X1_LOC_123/a_8_216# AND2X1_LOC_44/Y 0.01fF
C41322 OR2X1_LOC_184/Y OR2X1_LOC_226/a_8_216# 0.01fF
C41323 AND2X1_LOC_752/a_36_24# AND2X1_LOC_409/B 0.01fF
C41324 OR2X1_LOC_47/Y OR2X1_LOC_417/A 5.23fF
C41325 OR2X1_LOC_31/Y OR2X1_LOC_224/Y 0.01fF
C41326 AND2X1_LOC_705/Y VDD 0.21fF
C41327 AND2X1_LOC_434/a_8_24# OR2X1_LOC_428/A 0.08fF
C41328 OR2X1_LOC_246/A OR2X1_LOC_595/Y 0.51fF
C41329 AND2X1_LOC_725/a_8_24# OR2X1_LOC_421/Y 0.01fF
C41330 OR2X1_LOC_158/A AND2X1_LOC_244/a_8_24# 0.00fF
C41331 AND2X1_LOC_48/A OR2X1_LOC_196/a_8_216# 0.06fF
C41332 OR2X1_LOC_847/A OR2X1_LOC_622/B 0.01fF
C41333 OR2X1_LOC_599/A OR2X1_LOC_424/Y 0.00fF
C41334 OR2X1_LOC_175/Y OR2X1_LOC_756/B 0.00fF
C41335 AND2X1_LOC_253/a_8_24# OR2X1_LOC_562/A 0.24fF
C41336 OR2X1_LOC_47/Y OR2X1_LOC_64/a_8_216# 0.14fF
C41337 AND2X1_LOC_12/Y AND2X1_LOC_238/a_8_24# 0.01fF
C41338 OR2X1_LOC_696/A AND2X1_LOC_99/A 0.03fF
C41339 OR2X1_LOC_222/A OR2X1_LOC_539/B 0.02fF
C41340 OR2X1_LOC_269/B OR2X1_LOC_777/B 0.02fF
C41341 OR2X1_LOC_329/B OR2X1_LOC_16/A 0.04fF
C41342 AND2X1_LOC_811/Y AND2X1_LOC_808/A 0.05fF
C41343 OR2X1_LOC_139/A OR2X1_LOC_663/A 0.02fF
C41344 AND2X1_LOC_555/Y OR2X1_LOC_281/a_8_216# 0.01fF
C41345 OR2X1_LOC_87/A OR2X1_LOC_182/a_36_216# 0.00fF
C41346 AND2X1_LOC_712/a_8_24# AND2X1_LOC_605/Y 0.01fF
C41347 AND2X1_LOC_64/Y AND2X1_LOC_527/a_8_24# 0.18fF
C41348 OR2X1_LOC_539/Y OR2X1_LOC_319/Y 0.03fF
C41349 AND2X1_LOC_1/a_8_24# INPUT_6 0.04fF
C41350 OR2X1_LOC_62/B OR2X1_LOC_398/a_36_216# 0.00fF
C41351 OR2X1_LOC_654/A OR2X1_LOC_769/a_8_216# 0.05fF
C41352 OR2X1_LOC_235/B OR2X1_LOC_673/B 0.00fF
C41353 OR2X1_LOC_158/A AND2X1_LOC_161/Y 0.01fF
C41354 OR2X1_LOC_473/a_36_216# AND2X1_LOC_7/B 0.02fF
C41355 OR2X1_LOC_19/B OR2X1_LOC_789/A 0.02fF
C41356 OR2X1_LOC_53/Y OR2X1_LOC_689/a_8_216# 0.00fF
C41357 OR2X1_LOC_485/Y AND2X1_LOC_705/a_8_24# 0.07fF
C41358 OR2X1_LOC_505/Y AND2X1_LOC_807/B 0.01fF
C41359 AND2X1_LOC_64/Y AND2X1_LOC_314/a_36_24# 0.01fF
C41360 AND2X1_LOC_81/B OR2X1_LOC_130/Y 0.03fF
C41361 AND2X1_LOC_70/Y OR2X1_LOC_325/B 0.00fF
C41362 OR2X1_LOC_269/B AND2X1_LOC_591/a_36_24# 0.01fF
C41363 AND2X1_LOC_207/a_8_24# OR2X1_LOC_13/Y 0.01fF
C41364 AND2X1_LOC_538/a_36_24# AND2X1_LOC_434/Y 0.01fF
C41365 AND2X1_LOC_70/Y OR2X1_LOC_686/B 0.01fF
C41366 AND2X1_LOC_806/A OR2X1_LOC_504/a_36_216# 0.00fF
C41367 OR2X1_LOC_186/Y OR2X1_LOC_325/A 0.07fF
C41368 D_INPUT_0 OR2X1_LOC_779/B 0.02fF
C41369 OR2X1_LOC_502/A OR2X1_LOC_16/A 0.05fF
C41370 OR2X1_LOC_779/Y OR2X1_LOC_783/a_36_216# 0.03fF
C41371 AND2X1_LOC_94/a_36_24# OR2X1_LOC_397/Y 0.00fF
C41372 AND2X1_LOC_658/A AND2X1_LOC_807/B 0.10fF
C41373 OR2X1_LOC_73/a_8_216# AND2X1_LOC_789/Y 0.03fF
C41374 AND2X1_LOC_22/Y OR2X1_LOC_655/a_8_216# 0.02fF
C41375 AND2X1_LOC_3/Y AND2X1_LOC_36/Y 1.03fF
C41376 OR2X1_LOC_329/B OR2X1_LOC_108/Y 0.21fF
C41377 OR2X1_LOC_647/B AND2X1_LOC_36/Y 0.07fF
C41378 OR2X1_LOC_709/A AND2X1_LOC_423/a_8_24# 0.02fF
C41379 OR2X1_LOC_691/A AND2X1_LOC_690/a_8_24# 0.01fF
C41380 VDD AND2X1_LOC_19/Y 0.31fF
C41381 OR2X1_LOC_6/B AND2X1_LOC_54/a_8_24# 0.04fF
C41382 OR2X1_LOC_696/A AND2X1_LOC_637/Y 0.01fF
C41383 OR2X1_LOC_449/B OR2X1_LOC_168/Y 0.12fF
C41384 AND2X1_LOC_555/Y OR2X1_LOC_6/A 0.02fF
C41385 AND2X1_LOC_539/Y AND2X1_LOC_319/A 0.02fF
C41386 OR2X1_LOC_625/a_8_216# OR2X1_LOC_12/Y 0.04fF
C41387 AND2X1_LOC_787/a_8_24# AND2X1_LOC_212/Y 0.01fF
C41388 AND2X1_LOC_707/Y AND2X1_LOC_454/Y 0.10fF
C41389 OR2X1_LOC_160/B AND2X1_LOC_41/A 1.31fF
C41390 OR2X1_LOC_325/B OR2X1_LOC_703/A 0.05fF
C41391 AND2X1_LOC_792/Y AND2X1_LOC_793/Y 0.72fF
C41392 OR2X1_LOC_45/B OR2X1_LOC_39/A 0.29fF
C41393 OR2X1_LOC_187/a_8_216# OR2X1_LOC_40/Y 0.07fF
C41394 OR2X1_LOC_516/Y OR2X1_LOC_371/Y 0.03fF
C41395 OR2X1_LOC_186/Y OR2X1_LOC_447/A 0.01fF
C41396 AND2X1_LOC_364/Y OR2X1_LOC_426/B 0.04fF
C41397 OR2X1_LOC_78/A AND2X1_LOC_92/Y 0.14fF
C41398 OR2X1_LOC_264/Y OR2X1_LOC_509/a_36_216# 0.02fF
C41399 OR2X1_LOC_136/Y OR2X1_LOC_6/A 0.54fF
C41400 OR2X1_LOC_87/A OR2X1_LOC_392/B 3.89fF
C41401 AND2X1_LOC_663/A OR2X1_LOC_59/Y 0.05fF
C41402 OR2X1_LOC_364/A OR2X1_LOC_139/A 0.05fF
C41403 OR2X1_LOC_696/A AND2X1_LOC_512/a_36_24# 0.00fF
C41404 OR2X1_LOC_406/Y AND2X1_LOC_564/a_8_24# 0.01fF
C41405 AND2X1_LOC_340/Y OR2X1_LOC_316/Y 0.03fF
C41406 OR2X1_LOC_538/A AND2X1_LOC_110/a_36_24# 0.00fF
C41407 OR2X1_LOC_630/Y OR2X1_LOC_632/a_8_216# 0.04fF
C41408 OR2X1_LOC_715/B OR2X1_LOC_737/A 0.07fF
C41409 OR2X1_LOC_185/Y OR2X1_LOC_139/A 0.01fF
C41410 AND2X1_LOC_191/B OR2X1_LOC_755/Y 0.01fF
C41411 OR2X1_LOC_422/Y AND2X1_LOC_448/a_8_24# 0.01fF
C41412 AND2X1_LOC_456/a_8_24# OR2X1_LOC_44/Y 0.01fF
C41413 AND2X1_LOC_91/B OR2X1_LOC_383/a_8_216# 0.08fF
C41414 AND2X1_LOC_73/a_36_24# INPUT_0 0.01fF
C41415 OR2X1_LOC_864/A AND2X1_LOC_7/B 0.03fF
C41416 AND2X1_LOC_721/Y AND2X1_LOC_374/Y 0.01fF
C41417 OR2X1_LOC_179/a_8_216# OR2X1_LOC_178/Y 0.01fF
C41418 AND2X1_LOC_553/A VDD 0.17fF
C41419 OR2X1_LOC_447/Y OR2X1_LOC_714/A 0.01fF
C41420 VDD D_INPUT_4 0.53fF
C41421 AND2X1_LOC_562/B OR2X1_LOC_56/A 0.09fF
C41422 OR2X1_LOC_49/A AND2X1_LOC_29/a_8_24# 0.12fF
C41423 OR2X1_LOC_151/A OR2X1_LOC_161/A 1.02fF
C41424 OR2X1_LOC_715/B AND2X1_LOC_95/Y 0.03fF
C41425 AND2X1_LOC_705/Y AND2X1_LOC_447/a_36_24# 0.01fF
C41426 D_INPUT_7 AND2X1_LOC_587/a_8_24# 0.10fF
C41427 AND2X1_LOC_95/Y AND2X1_LOC_626/a_8_24# 0.10fF
C41428 AND2X1_LOC_532/a_8_24# OR2X1_LOC_604/A 0.16fF
C41429 AND2X1_LOC_22/Y OR2X1_LOC_810/A 0.16fF
C41430 OR2X1_LOC_307/a_8_216# AND2X1_LOC_22/Y 0.01fF
C41431 VDD AND2X1_LOC_804/Y 0.21fF
C41432 AND2X1_LOC_95/Y OR2X1_LOC_543/A 0.48fF
C41433 OR2X1_LOC_231/B OR2X1_LOC_643/A 0.05fF
C41434 OR2X1_LOC_850/B OR2X1_LOC_363/A 0.00fF
C41435 AND2X1_LOC_354/B AND2X1_LOC_810/B 0.01fF
C41436 OR2X1_LOC_840/A OR2X1_LOC_78/B 1.52fF
C41437 OR2X1_LOC_448/B AND2X1_LOC_92/Y 0.00fF
C41438 OR2X1_LOC_305/Y OR2X1_LOC_135/Y 0.01fF
C41439 AND2X1_LOC_70/Y OR2X1_LOC_788/a_36_216# 0.00fF
C41440 OR2X1_LOC_163/a_8_216# OR2X1_LOC_163/Y 0.01fF
C41441 OR2X1_LOC_528/Y AND2X1_LOC_624/A 4.47fF
C41442 OR2X1_LOC_45/B AND2X1_LOC_211/B 0.04fF
C41443 OR2X1_LOC_40/Y OR2X1_LOC_127/Y 0.21fF
C41444 OR2X1_LOC_406/Y OR2X1_LOC_74/A 0.03fF
C41445 OR2X1_LOC_121/Y OR2X1_LOC_643/A 0.43fF
C41446 OR2X1_LOC_158/A AND2X1_LOC_286/Y 0.04fF
C41447 OR2X1_LOC_619/Y AND2X1_LOC_658/a_8_24# 0.01fF
C41448 OR2X1_LOC_7/A OR2X1_LOC_753/a_8_216# -0.01fF
C41449 OR2X1_LOC_702/A OR2X1_LOC_138/a_36_216# 0.03fF
C41450 OR2X1_LOC_269/B OR2X1_LOC_344/A 0.03fF
C41451 OR2X1_LOC_121/Y OR2X1_LOC_124/Y 0.01fF
C41452 AND2X1_LOC_348/A OR2X1_LOC_91/A 0.05fF
C41453 AND2X1_LOC_40/Y OR2X1_LOC_235/B 0.07fF
C41454 AND2X1_LOC_658/B AND2X1_LOC_550/A 0.03fF
C41455 AND2X1_LOC_22/Y AND2X1_LOC_589/a_8_24# 0.03fF
C41456 AND2X1_LOC_52/Y OR2X1_LOC_197/a_8_216# 0.01fF
C41457 OR2X1_LOC_502/A AND2X1_LOC_167/a_8_24# 0.03fF
C41458 OR2X1_LOC_254/a_36_216# OR2X1_LOC_562/A 0.00fF
C41459 AND2X1_LOC_3/Y AND2X1_LOC_488/a_8_24# 0.02fF
C41460 AND2X1_LOC_784/A AND2X1_LOC_515/a_36_24# 0.00fF
C41461 D_INPUT_5 AND2X1_LOC_12/a_8_24# 0.01fF
C41462 OR2X1_LOC_589/A AND2X1_LOC_264/a_8_24# 0.17fF
C41463 OR2X1_LOC_744/A OR2X1_LOC_48/B 1.17fF
C41464 AND2X1_LOC_571/Y AND2X1_LOC_561/B 0.03fF
C41465 OR2X1_LOC_122/a_8_216# AND2X1_LOC_99/A 0.01fF
C41466 OR2X1_LOC_49/A OR2X1_LOC_622/a_8_216# 0.06fF
C41467 AND2X1_LOC_70/Y OR2X1_LOC_405/Y 0.01fF
C41468 OR2X1_LOC_124/a_8_216# OR2X1_LOC_375/A 0.01fF
C41469 AND2X1_LOC_729/Y OR2X1_LOC_679/Y 0.01fF
C41470 OR2X1_LOC_516/a_8_216# OR2X1_LOC_600/A 0.01fF
C41471 AND2X1_LOC_259/Y OR2X1_LOC_381/a_8_216# 0.01fF
C41472 VDD OR2X1_LOC_511/Y 0.17fF
C41473 OR2X1_LOC_375/A OR2X1_LOC_370/a_36_216# 0.00fF
C41474 OR2X1_LOC_168/a_8_216# OR2X1_LOC_168/B 0.07fF
C41475 VDD OR2X1_LOC_865/Y 0.00fF
C41476 OR2X1_LOC_744/A OR2X1_LOC_18/Y 6.11fF
C41477 OR2X1_LOC_47/Y AND2X1_LOC_247/a_8_24# 0.02fF
C41478 OR2X1_LOC_191/B OR2X1_LOC_565/A 0.34fF
C41479 AND2X1_LOC_711/Y OR2X1_LOC_759/a_36_216# 0.00fF
C41480 AND2X1_LOC_716/Y AND2X1_LOC_335/a_36_24# 0.00fF
C41481 AND2X1_LOC_390/B AND2X1_LOC_810/B 0.00fF
C41482 AND2X1_LOC_675/Y AND2X1_LOC_621/Y 0.03fF
C41483 OR2X1_LOC_450/A OR2X1_LOC_87/A 0.03fF
C41484 OR2X1_LOC_158/A AND2X1_LOC_356/B 0.03fF
C41485 OR2X1_LOC_304/a_36_216# OR2X1_LOC_431/Y 0.01fF
C41486 VDD OR2X1_LOC_673/Y 0.12fF
C41487 OR2X1_LOC_17/Y OR2X1_LOC_36/a_8_216# 0.08fF
C41488 AND2X1_LOC_74/a_8_24# OR2X1_LOC_464/A 0.01fF
C41489 OR2X1_LOC_160/B OR2X1_LOC_631/B 0.03fF
C41490 OR2X1_LOC_158/A OR2X1_LOC_280/Y 4.57fF
C41491 OR2X1_LOC_624/A OR2X1_LOC_174/A 0.03fF
C41492 OR2X1_LOC_570/a_8_216# OR2X1_LOC_570/A 0.39fF
C41493 OR2X1_LOC_51/Y OR2X1_LOC_6/A 1.45fF
C41494 OR2X1_LOC_518/a_36_216# OR2X1_LOC_111/Y 0.00fF
C41495 OR2X1_LOC_485/A AND2X1_LOC_476/Y 0.07fF
C41496 OR2X1_LOC_318/A AND2X1_LOC_51/Y 0.01fF
C41497 OR2X1_LOC_709/A OR2X1_LOC_193/A 0.54fF
C41498 OR2X1_LOC_329/Y AND2X1_LOC_337/B 0.14fF
C41499 OR2X1_LOC_78/B OR2X1_LOC_222/A 0.26fF
C41500 OR2X1_LOC_270/Y AND2X1_LOC_36/Y 0.01fF
C41501 OR2X1_LOC_510/Y OR2X1_LOC_244/B 0.05fF
C41502 OR2X1_LOC_709/A AND2X1_LOC_136/a_36_24# 0.00fF
C41503 OR2X1_LOC_750/A AND2X1_LOC_44/Y 0.06fF
C41504 OR2X1_LOC_283/a_8_216# OR2X1_LOC_59/Y 0.01fF
C41505 AND2X1_LOC_41/A OR2X1_LOC_553/A 0.08fF
C41506 OR2X1_LOC_287/B OR2X1_LOC_858/a_8_216# 0.01fF
C41507 OR2X1_LOC_814/A OR2X1_LOC_366/B 0.07fF
C41508 OR2X1_LOC_448/Y OR2X1_LOC_708/Y 0.03fF
C41509 INPUT_5 OR2X1_LOC_1/a_36_216# -0.00fF
C41510 OR2X1_LOC_792/Y OR2X1_LOC_286/Y 0.04fF
C41511 OR2X1_LOC_696/A AND2X1_LOC_319/a_8_24# 0.03fF
C41512 OR2X1_LOC_681/a_36_216# OR2X1_LOC_743/A 0.03fF
C41513 VDD OR2X1_LOC_297/Y 0.12fF
C41514 OR2X1_LOC_151/A AND2X1_LOC_51/Y 0.14fF
C41515 AND2X1_LOC_539/Y AND2X1_LOC_170/B 0.12fF
C41516 AND2X1_LOC_802/B OR2X1_LOC_167/Y 0.02fF
C41517 VDD OR2X1_LOC_195/A -0.00fF
C41518 AND2X1_LOC_474/A OR2X1_LOC_44/Y 0.08fF
C41519 OR2X1_LOC_840/A OR2X1_LOC_375/A 0.01fF
C41520 OR2X1_LOC_677/Y OR2X1_LOC_511/Y 0.01fF
C41521 AND2X1_LOC_474/A AND2X1_LOC_288/a_8_24# 0.01fF
C41522 OR2X1_LOC_625/a_36_216# OR2X1_LOC_278/Y 0.00fF
C41523 OR2X1_LOC_155/A AND2X1_LOC_92/Y 0.20fF
C41524 OR2X1_LOC_51/Y AND2X1_LOC_673/a_36_24# 0.00fF
C41525 OR2X1_LOC_134/Y AND2X1_LOC_137/a_8_24# 0.00fF
C41526 OR2X1_LOC_231/A OR2X1_LOC_231/a_8_216# 0.01fF
C41527 VDD AND2X1_LOC_345/Y 0.05fF
C41528 OR2X1_LOC_473/a_36_216# OR2X1_LOC_805/A 0.01fF
C41529 OR2X1_LOC_148/a_8_216# OR2X1_LOC_471/Y 0.14fF
C41530 AND2X1_LOC_339/B AND2X1_LOC_537/Y 0.22fF
C41531 OR2X1_LOC_244/A OR2X1_LOC_576/A 0.02fF
C41532 OR2X1_LOC_811/A OR2X1_LOC_347/B 0.19fF
C41533 OR2X1_LOC_538/A OR2X1_LOC_778/Y 0.03fF
C41534 OR2X1_LOC_216/A OR2X1_LOC_203/Y 0.01fF
C41535 OR2X1_LOC_630/Y AND2X1_LOC_3/Y 0.01fF
C41536 OR2X1_LOC_160/B AND2X1_LOC_135/a_8_24# 0.01fF
C41537 AND2X1_LOC_36/Y OR2X1_LOC_196/a_36_216# 0.00fF
C41538 OR2X1_LOC_589/A OR2X1_LOC_46/A 0.03fF
C41539 OR2X1_LOC_769/B OR2X1_LOC_654/A 0.03fF
C41540 OR2X1_LOC_432/Y OR2X1_LOC_433/Y 0.33fF
C41541 AND2X1_LOC_667/a_8_24# OR2X1_LOC_549/A 0.03fF
C41542 AND2X1_LOC_41/A OR2X1_LOC_219/B 0.03fF
C41543 OR2X1_LOC_158/A OR2X1_LOC_22/Y 2.94fF
C41544 OR2X1_LOC_36/Y OR2X1_LOC_92/Y 0.39fF
C41545 AND2X1_LOC_393/a_8_24# AND2X1_LOC_40/Y 0.05fF
C41546 OR2X1_LOC_709/A D_INPUT_0 0.02fF
C41547 AND2X1_LOC_732/B OR2X1_LOC_64/Y 0.00fF
C41548 AND2X1_LOC_544/Y OR2X1_LOC_47/Y 0.15fF
C41549 OR2X1_LOC_603/a_8_216# OR2X1_LOC_427/A 0.01fF
C41550 AND2X1_LOC_95/Y OR2X1_LOC_215/Y 0.07fF
C41551 OR2X1_LOC_66/Y OR2X1_LOC_130/Y 0.18fF
C41552 OR2X1_LOC_19/B AND2X1_LOC_606/a_8_24# 0.02fF
C41553 OR2X1_LOC_517/A AND2X1_LOC_105/a_8_24# 0.09fF
C41554 OR2X1_LOC_260/a_8_216# OR2X1_LOC_375/A 0.18fF
C41555 AND2X1_LOC_70/Y OR2X1_LOC_193/A 0.02fF
C41556 AND2X1_LOC_344/a_8_24# AND2X1_LOC_363/A 0.01fF
C41557 OR2X1_LOC_464/A OR2X1_LOC_722/a_8_216# 0.01fF
C41558 AND2X1_LOC_711/Y AND2X1_LOC_663/A 0.00fF
C41559 AND2X1_LOC_849/A AND2X1_LOC_489/a_8_24# 0.10fF
C41560 OR2X1_LOC_327/a_8_216# OR2X1_LOC_216/Y 0.03fF
C41561 AND2X1_LOC_59/Y OR2X1_LOC_541/B 0.03fF
C41562 OR2X1_LOC_145/a_8_216# OR2X1_LOC_427/A 0.01fF
C41563 OR2X1_LOC_231/a_8_216# OR2X1_LOC_130/A 0.03fF
C41564 OR2X1_LOC_70/Y AND2X1_LOC_663/A 0.01fF
C41565 OR2X1_LOC_528/Y AND2X1_LOC_621/a_8_24# 0.01fF
C41566 OR2X1_LOC_599/A AND2X1_LOC_841/B 0.18fF
C41567 AND2X1_LOC_42/B OR2X1_LOC_735/a_8_216# 0.05fF
C41568 OR2X1_LOC_755/A OR2X1_LOC_816/Y 0.00fF
C41569 OR2X1_LOC_516/Y AND2X1_LOC_222/Y 0.03fF
C41570 OR2X1_LOC_177/Y AND2X1_LOC_675/A -0.00fF
C41571 AND2X1_LOC_145/a_8_24# OR2X1_LOC_375/A 0.04fF
C41572 OR2X1_LOC_635/A AND2X1_LOC_3/Y 0.06fF
C41573 OR2X1_LOC_573/Y OR2X1_LOC_575/a_8_216# 0.39fF
C41574 OR2X1_LOC_3/Y AND2X1_LOC_401/Y 0.00fF
C41575 OR2X1_LOC_18/Y AND2X1_LOC_840/B 0.05fF
C41576 VDD AND2X1_LOC_425/Y 0.46fF
C41577 OR2X1_LOC_467/B OR2X1_LOC_477/a_36_216# 0.00fF
C41578 OR2X1_LOC_589/A AND2X1_LOC_227/Y 0.05fF
C41579 VDD AND2X1_LOC_309/a_8_24# -0.00fF
C41580 AND2X1_LOC_593/Y OR2X1_LOC_44/Y 0.00fF
C41581 OR2X1_LOC_71/Y AND2X1_LOC_243/Y 0.03fF
C41582 OR2X1_LOC_611/Y OR2X1_LOC_612/a_8_216# 0.39fF
C41583 AND2X1_LOC_174/a_36_24# OR2X1_LOC_6/A 0.00fF
C41584 INPUT_5 OR2X1_LOC_17/Y 0.35fF
C41585 OR2X1_LOC_3/Y OR2X1_LOC_426/A 0.01fF
C41586 OR2X1_LOC_36/Y OR2X1_LOC_65/B 0.03fF
C41587 OR2X1_LOC_241/a_36_216# OR2X1_LOC_375/A 0.00fF
C41588 AND2X1_LOC_141/B OR2X1_LOC_517/A 0.07fF
C41589 AND2X1_LOC_12/Y OR2X1_LOC_643/A 0.03fF
C41590 OR2X1_LOC_123/a_8_216# OR2X1_LOC_720/B 0.47fF
C41591 AND2X1_LOC_91/B OR2X1_LOC_318/B 0.03fF
C41592 AND2X1_LOC_6/a_8_24# OR2X1_LOC_633/A 0.01fF
C41593 OR2X1_LOC_519/a_36_216# AND2X1_LOC_211/B 0.01fF
C41594 AND2X1_LOC_12/Y OR2X1_LOC_778/Y 0.22fF
C41595 OR2X1_LOC_685/A OR2X1_LOC_87/A 0.01fF
C41596 AND2X1_LOC_70/Y D_INPUT_0 0.23fF
C41597 AND2X1_LOC_580/A AND2X1_LOC_576/Y 0.07fF
C41598 AND2X1_LOC_808/A AND2X1_LOC_469/a_8_24# 0.01fF
C41599 AND2X1_LOC_586/a_8_24# AND2X1_LOC_3/Y 0.01fF
C41600 AND2X1_LOC_682/a_36_24# AND2X1_LOC_3/Y 0.00fF
C41601 OR2X1_LOC_477/Y AND2X1_LOC_51/Y 0.03fF
C41602 OR2X1_LOC_70/Y OR2X1_LOC_2/Y 0.10fF
C41603 OR2X1_LOC_111/Y AND2X1_LOC_715/A 0.01fF
C41604 OR2X1_LOC_85/A OR2X1_LOC_44/Y 0.21fF
C41605 VDD OR2X1_LOC_770/a_8_216# 0.00fF
C41606 OR2X1_LOC_316/Y OR2X1_LOC_585/A 0.03fF
C41607 AND2X1_LOC_29/a_8_24# OR2X1_LOC_87/B 0.04fF
C41608 AND2X1_LOC_191/B AND2X1_LOC_845/Y 0.65fF
C41609 OR2X1_LOC_291/a_8_216# OR2X1_LOC_291/A 0.05fF
C41610 OR2X1_LOC_632/a_36_216# OR2X1_LOC_62/B 0.00fF
C41611 OR2X1_LOC_160/A OR2X1_LOC_574/A 0.26fF
C41612 AND2X1_LOC_539/Y OR2X1_LOC_331/Y 0.06fF
C41613 AND2X1_LOC_51/Y OR2X1_LOC_788/a_8_216# 0.01fF
C41614 OR2X1_LOC_271/Y OR2X1_LOC_36/Y 0.01fF
C41615 OR2X1_LOC_772/a_8_216# OR2X1_LOC_269/B 0.01fF
C41616 OR2X1_LOC_592/A OR2X1_LOC_185/A 0.03fF
C41617 OR2X1_LOC_40/Y OR2X1_LOC_615/Y 0.03fF
C41618 VDD AND2X1_LOC_649/Y 0.01fF
C41619 AND2X1_LOC_98/a_8_24# D_INPUT_3 0.01fF
C41620 OR2X1_LOC_504/Y AND2X1_LOC_663/A 0.19fF
C41621 VDD AND2X1_LOC_451/Y 0.08fF
C41622 OR2X1_LOC_6/B OR2X1_LOC_786/Y 0.03fF
C41623 OR2X1_LOC_377/A OR2X1_LOC_20/a_8_216# 0.06fF
C41624 OR2X1_LOC_97/B AND2X1_LOC_8/Y 0.15fF
C41625 OR2X1_LOC_426/A OR2X1_LOC_582/Y 0.01fF
C41626 AND2X1_LOC_243/Y D_INPUT_1 0.06fF
C41627 VDD AND2X1_LOC_648/B 0.30fF
C41628 OR2X1_LOC_103/Y OR2X1_LOC_22/Y 0.08fF
C41629 OR2X1_LOC_267/Y OR2X1_LOC_560/A 0.09fF
C41630 OR2X1_LOC_105/a_8_216# OR2X1_LOC_814/A 0.01fF
C41631 OR2X1_LOC_756/B AND2X1_LOC_283/a_8_24# 0.02fF
C41632 OR2X1_LOC_833/Y OR2X1_LOC_717/a_8_216# 0.14fF
C41633 AND2X1_LOC_99/A AND2X1_LOC_663/B 0.03fF
C41634 AND2X1_LOC_41/A OR2X1_LOC_244/A 0.00fF
C41635 OR2X1_LOC_3/Y INPUT_4 0.06fF
C41636 AND2X1_LOC_483/a_8_24# AND2X1_LOC_624/A 0.02fF
C41637 OR2X1_LOC_857/B OR2X1_LOC_598/A 0.16fF
C41638 OR2X1_LOC_486/Y OR2X1_LOC_365/B 0.13fF
C41639 OR2X1_LOC_272/Y AND2X1_LOC_139/B 0.03fF
C41640 OR2X1_LOC_625/Y OR2X1_LOC_64/Y 0.04fF
C41641 AND2X1_LOC_7/B AND2X1_LOC_751/a_36_24# 0.01fF
C41642 OR2X1_LOC_272/Y OR2X1_LOC_767/a_36_216# 0.00fF
C41643 AND2X1_LOC_53/Y AND2X1_LOC_693/a_36_24# -0.01fF
C41644 D_INPUT_4 AND2X1_LOC_25/a_8_24# 0.01fF
C41645 AND2X1_LOC_340/Y OR2X1_LOC_153/a_8_216# 0.04fF
C41646 OR2X1_LOC_65/B OR2X1_LOC_65/a_8_216# 0.02fF
C41647 AND2X1_LOC_611/a_8_24# AND2X1_LOC_612/B 0.02fF
C41648 OR2X1_LOC_103/a_8_216# OR2X1_LOC_22/Y 0.01fF
C41649 OR2X1_LOC_346/B AND2X1_LOC_3/Y 0.01fF
C41650 OR2X1_LOC_726/a_8_216# OR2X1_LOC_731/B -0.00fF
C41651 OR2X1_LOC_51/Y OR2X1_LOC_289/a_8_216# 0.02fF
C41652 AND2X1_LOC_307/Y AND2X1_LOC_655/A 0.05fF
C41653 OR2X1_LOC_47/Y OR2X1_LOC_232/Y 0.03fF
C41654 OR2X1_LOC_193/A OR2X1_LOC_193/Y 0.06fF
C41655 OR2X1_LOC_563/A OR2X1_LOC_366/Y 0.07fF
C41656 AND2X1_LOC_792/a_8_24# AND2X1_LOC_789/Y -0.02fF
C41657 OR2X1_LOC_804/B OR2X1_LOC_778/Y 0.10fF
C41658 AND2X1_LOC_47/Y OR2X1_LOC_785/B 0.01fF
C41659 OR2X1_LOC_3/Y AND2X1_LOC_123/a_8_24# 0.01fF
C41660 AND2X1_LOC_390/B OR2X1_LOC_585/A 0.01fF
C41661 AND2X1_LOC_368/a_8_24# OR2X1_LOC_270/Y 0.11fF
C41662 OR2X1_LOC_668/a_8_216# OR2X1_LOC_532/B 0.01fF
C41663 INPUT_4 OR2X1_LOC_582/Y 0.01fF
C41664 OR2X1_LOC_476/B AND2X1_LOC_32/a_8_24# 0.02fF
C41665 OR2X1_LOC_304/Y OR2X1_LOC_52/B 0.06fF
C41666 OR2X1_LOC_316/Y AND2X1_LOC_634/Y 0.03fF
C41667 OR2X1_LOC_80/A OR2X1_LOC_549/A 0.05fF
C41668 AND2X1_LOC_319/A AND2X1_LOC_687/A 0.19fF
C41669 OR2X1_LOC_625/Y OR2X1_LOC_417/A 0.09fF
C41670 OR2X1_LOC_31/Y OR2X1_LOC_48/B 0.38fF
C41671 AND2X1_LOC_122/a_8_24# AND2X1_LOC_3/Y 0.01fF
C41672 AND2X1_LOC_42/B AND2X1_LOC_38/a_8_24# 0.01fF
C41673 OR2X1_LOC_33/A OR2X1_LOC_33/a_8_216# 0.47fF
C41674 OR2X1_LOC_429/Y OR2X1_LOC_430/a_8_216# 0.06fF
C41675 INPUT_5 OR2X1_LOC_588/A 0.01fF
C41676 OR2X1_LOC_18/Y OR2X1_LOC_31/Y 0.22fF
C41677 AND2X1_LOC_711/Y OR2X1_LOC_617/a_8_216# 0.02fF
C41678 OR2X1_LOC_145/Y OR2X1_LOC_427/A 0.02fF
C41679 OR2X1_LOC_369/Y AND2X1_LOC_222/Y 0.03fF
C41680 OR2X1_LOC_43/A OR2X1_LOC_46/A 0.56fF
C41681 OR2X1_LOC_703/B OR2X1_LOC_532/B 0.01fF
C41682 OR2X1_LOC_3/Y OR2X1_LOC_277/a_8_216# 0.01fF
C41683 OR2X1_LOC_656/B OR2X1_LOC_227/Y 0.01fF
C41684 AND2X1_LOC_59/Y OR2X1_LOC_440/A 0.03fF
C41685 OR2X1_LOC_87/A OR2X1_LOC_532/B 0.42fF
C41686 OR2X1_LOC_62/B OR2X1_LOC_612/B 0.01fF
C41687 OR2X1_LOC_116/a_8_216# D_INPUT_0 -0.04fF
C41688 OR2X1_LOC_26/Y INPUT_1 0.09fF
C41689 OR2X1_LOC_241/Y OR2X1_LOC_375/A 0.01fF
C41690 OR2X1_LOC_92/Y OR2X1_LOC_85/a_8_216# 0.33fF
C41691 AND2X1_LOC_102/a_36_24# OR2X1_LOC_54/Y 0.01fF
C41692 D_INPUT_0 AND2X1_LOC_361/A 0.07fF
C41693 OR2X1_LOC_687/Y AND2X1_LOC_47/Y 0.06fF
C41694 AND2X1_LOC_550/A OR2X1_LOC_47/Y 0.03fF
C41695 AND2X1_LOC_47/Y OR2X1_LOC_781/A 0.15fF
C41696 OR2X1_LOC_691/a_8_216# OR2X1_LOC_771/B 0.02fF
C41697 OR2X1_LOC_255/a_36_216# OR2X1_LOC_248/Y 0.06fF
C41698 AND2X1_LOC_654/B OR2X1_LOC_41/Y 0.16fF
C41699 AND2X1_LOC_399/a_8_24# AND2X1_LOC_47/Y 0.02fF
C41700 AND2X1_LOC_514/Y AND2X1_LOC_212/B 0.08fF
C41701 OR2X1_LOC_130/A AND2X1_LOC_109/a_8_24# 0.03fF
C41702 AND2X1_LOC_152/a_8_24# AND2X1_LOC_47/Y 0.02fF
C41703 AND2X1_LOC_372/a_8_24# AND2X1_LOC_31/Y 0.01fF
C41704 AND2X1_LOC_40/Y OR2X1_LOC_580/a_8_216# 0.01fF
C41705 AND2X1_LOC_810/Y AND2X1_LOC_653/a_8_24# 0.09fF
C41706 OR2X1_LOC_741/Y OR2X1_LOC_367/B 0.03fF
C41707 OR2X1_LOC_43/A AND2X1_LOC_227/Y 0.03fF
C41708 AND2X1_LOC_151/a_8_24# AND2X1_LOC_810/Y 0.09fF
C41709 OR2X1_LOC_472/B OR2X1_LOC_27/Y 0.08fF
C41710 AND2X1_LOC_639/A AND2X1_LOC_639/a_36_24# 0.01fF
C41711 INPUT_1 OR2X1_LOC_820/Y 0.01fF
C41712 OR2X1_LOC_2/Y OR2X1_LOC_70/A 0.83fF
C41713 OR2X1_LOC_11/Y OR2X1_LOC_3/B 0.33fF
C41714 VDD OR2X1_LOC_769/a_8_216# 0.21fF
C41715 OR2X1_LOC_656/a_8_216# OR2X1_LOC_121/B 0.01fF
C41716 OR2X1_LOC_673/Y OR2X1_LOC_845/A 0.04fF
C41717 OR2X1_LOC_113/B OR2X1_LOC_844/B 0.00fF
C41718 OR2X1_LOC_311/Y AND2X1_LOC_856/B 0.01fF
C41719 OR2X1_LOC_715/A OR2X1_LOC_446/B 0.24fF
C41720 OR2X1_LOC_128/a_8_216# AND2X1_LOC_72/B 0.01fF
C41721 AND2X1_LOC_778/a_36_24# AND2X1_LOC_785/Y 0.01fF
C41722 OR2X1_LOC_45/B AND2X1_LOC_785/a_8_24# 0.01fF
C41723 OR2X1_LOC_40/Y D_INPUT_6 0.04fF
C41724 AND2X1_LOC_7/B OR2X1_LOC_121/A 0.05fF
C41725 VDD OR2X1_LOC_723/B 0.02fF
C41726 OR2X1_LOC_269/a_8_216# OR2X1_LOC_675/Y 0.14fF
C41727 OR2X1_LOC_205/Y OR2X1_LOC_203/Y 0.02fF
C41728 OR2X1_LOC_161/B OR2X1_LOC_556/a_36_216# 0.00fF
C41729 OR2X1_LOC_429/Y OR2X1_LOC_428/Y 0.27fF
C41730 AND2X1_LOC_70/Y OR2X1_LOC_339/A 0.21fF
C41731 OR2X1_LOC_7/A OR2X1_LOC_615/Y 0.15fF
C41732 OR2X1_LOC_66/A OR2X1_LOC_593/B 0.04fF
C41733 OR2X1_LOC_566/A OR2X1_LOC_337/A 0.74fF
C41734 OR2X1_LOC_43/A OR2X1_LOC_813/Y 0.07fF
C41735 OR2X1_LOC_841/A OR2X1_LOC_593/B 0.49fF
C41736 OR2X1_LOC_176/Y AND2X1_LOC_787/A 0.00fF
C41737 AND2X1_LOC_3/Y OR2X1_LOC_340/a_8_216# 0.01fF
C41738 OR2X1_LOC_115/B OR2X1_LOC_549/A 0.11fF
C41739 OR2X1_LOC_377/A OR2X1_LOC_750/Y 0.82fF
C41740 OR2X1_LOC_816/A OR2X1_LOC_753/a_36_216# 0.02fF
C41741 OR2X1_LOC_43/A OR2X1_LOC_41/Y 0.10fF
C41742 OR2X1_LOC_62/B AND2X1_LOC_15/a_8_24# 0.03fF
C41743 OR2X1_LOC_74/a_8_216# AND2X1_LOC_215/A 0.47fF
C41744 OR2X1_LOC_428/A AND2X1_LOC_786/Y 0.05fF
C41745 OR2X1_LOC_191/B OR2X1_LOC_551/B 0.04fF
C41746 AND2X1_LOC_787/A AND2X1_LOC_212/Y 0.01fF
C41747 INPUT_0 AND2X1_LOC_36/Y 5.83fF
C41748 OR2X1_LOC_653/B OR2X1_LOC_97/A 0.00fF
C41749 AND2X1_LOC_91/B OR2X1_LOC_114/B 0.03fF
C41750 OR2X1_LOC_53/Y AND2X1_LOC_194/Y 0.02fF
C41751 OR2X1_LOC_208/A AND2X1_LOC_70/Y 0.01fF
C41752 OR2X1_LOC_40/Y AND2X1_LOC_242/B 0.01fF
C41753 OR2X1_LOC_600/A OR2X1_LOC_748/Y 0.01fF
C41754 OR2X1_LOC_176/Y AND2X1_LOC_566/B 0.51fF
C41755 OR2X1_LOC_715/B AND2X1_LOC_22/Y 0.03fF
C41756 VDD OR2X1_LOC_56/a_8_216# 0.00fF
C41757 VDD AND2X1_LOC_465/A 0.34fF
C41758 AND2X1_LOC_91/B AND2X1_LOC_396/a_8_24# 0.04fF
C41759 AND2X1_LOC_705/Y AND2X1_LOC_713/a_8_24# 0.09fF
C41760 OR2X1_LOC_625/Y AND2X1_LOC_247/a_8_24# 0.02fF
C41761 AND2X1_LOC_566/B AND2X1_LOC_212/Y 0.02fF
C41762 VDD OR2X1_LOC_158/Y 0.12fF
C41763 OR2X1_LOC_709/A OR2X1_LOC_515/A 0.01fF
C41764 OR2X1_LOC_61/A AND2X1_LOC_18/Y 0.01fF
C41765 OR2X1_LOC_487/a_8_216# AND2X1_LOC_657/A 0.02fF
C41766 OR2X1_LOC_439/B OR2X1_LOC_180/a_8_216# 0.16fF
C41767 OR2X1_LOC_428/a_8_216# OR2X1_LOC_428/Y 0.01fF
C41768 AND2X1_LOC_91/B OR2X1_LOC_538/A 0.03fF
C41769 OR2X1_LOC_421/A OR2X1_LOC_693/Y 0.01fF
C41770 AND2X1_LOC_773/Y OR2X1_LOC_426/B 0.81fF
C41771 OR2X1_LOC_532/B AND2X1_LOC_109/a_36_24# 0.01fF
C41772 AND2X1_LOC_42/B OR2X1_LOC_68/B 0.17fF
C41773 OR2X1_LOC_744/A OR2X1_LOC_764/a_8_216# 0.01fF
C41774 AND2X1_LOC_181/Y OR2X1_LOC_309/Y 0.00fF
C41775 AND2X1_LOC_352/a_8_24# AND2X1_LOC_566/B 0.01fF
C41776 OR2X1_LOC_732/B AND2X1_LOC_36/Y 0.04fF
C41777 AND2X1_LOC_727/Y OR2X1_LOC_441/Y 0.03fF
C41778 OR2X1_LOC_789/B AND2X1_LOC_36/Y 0.01fF
C41779 AND2X1_LOC_70/a_8_24# AND2X1_LOC_44/Y 0.01fF
C41780 AND2X1_LOC_548/Y OR2X1_LOC_816/A 0.01fF
C41781 OR2X1_LOC_850/B OR2X1_LOC_366/A 0.01fF
C41782 AND2X1_LOC_197/Y OR2X1_LOC_56/Y 0.21fF
C41783 AND2X1_LOC_70/Y AND2X1_LOC_438/a_8_24# 0.01fF
C41784 OR2X1_LOC_154/A OR2X1_LOC_590/Y 0.04fF
C41785 OR2X1_LOC_447/a_8_216# OR2X1_LOC_308/Y 0.03fF
C41786 OR2X1_LOC_615/a_36_216# AND2X1_LOC_562/Y 0.15fF
C41787 AND2X1_LOC_566/B AND2X1_LOC_353/a_36_24# 0.00fF
C41788 AND2X1_LOC_40/Y AND2X1_LOC_226/a_8_24# 0.03fF
C41789 OR2X1_LOC_324/B AND2X1_LOC_44/Y 0.21fF
C41790 OR2X1_LOC_124/a_8_216# OR2X1_LOC_549/A 0.04fF
C41791 OR2X1_LOC_662/a_8_216# AND2X1_LOC_44/Y 0.03fF
C41792 OR2X1_LOC_45/B OR2X1_LOC_421/a_8_216# 0.02fF
C41793 AND2X1_LOC_340/Y OR2X1_LOC_744/A 0.01fF
C41794 OR2X1_LOC_629/Y OR2X1_LOC_140/B 0.01fF
C41795 AND2X1_LOC_796/Y AND2X1_LOC_803/a_8_24# 0.10fF
C41796 OR2X1_LOC_329/B OR2X1_LOC_373/Y 0.07fF
C41797 OR2X1_LOC_744/A AND2X1_LOC_810/B 0.24fF
C41798 OR2X1_LOC_40/Y OR2X1_LOC_813/a_8_216# 0.02fF
C41799 AND2X1_LOC_64/Y OR2X1_LOC_620/Y 0.24fF
C41800 AND2X1_LOC_70/Y OR2X1_LOC_831/A 0.03fF
C41801 OR2X1_LOC_97/A OR2X1_LOC_808/B 0.03fF
C41802 OR2X1_LOC_7/A OR2X1_LOC_424/Y -0.03fF
C41803 OR2X1_LOC_563/B D_GATE_366 0.02fF
C41804 OR2X1_LOC_290/a_8_216# AND2X1_LOC_219/A 0.03fF
C41805 AND2X1_LOC_95/Y OR2X1_LOC_338/B 0.01fF
C41806 AND2X1_LOC_181/Y OR2X1_LOC_744/A 0.04fF
C41807 OR2X1_LOC_862/B OR2X1_LOC_362/A 0.01fF
C41808 AND2X1_LOC_443/a_36_24# OR2X1_LOC_56/A 0.01fF
C41809 AND2X1_LOC_736/Y AND2X1_LOC_734/a_8_24# 0.03fF
C41810 OR2X1_LOC_31/Y AND2X1_LOC_215/A 0.03fF
C41811 AND2X1_LOC_70/Y OR2X1_LOC_598/Y 0.12fF
C41812 OR2X1_LOC_426/B AND2X1_LOC_243/Y 0.17fF
C41813 AND2X1_LOC_754/a_8_24# OR2X1_LOC_78/B 0.03fF
C41814 OR2X1_LOC_790/A OR2X1_LOC_78/A 0.01fF
C41815 AND2X1_LOC_17/a_8_24# INPUT_6 0.04fF
C41816 AND2X1_LOC_70/Y AND2X1_LOC_131/a_8_24# 0.01fF
C41817 OR2X1_LOC_141/B OR2X1_LOC_217/A 0.01fF
C41818 AND2X1_LOC_95/Y OR2X1_LOC_334/a_36_216# 0.00fF
C41819 AND2X1_LOC_142/a_8_24# AND2X1_LOC_44/Y 0.02fF
C41820 VDD OR2X1_LOC_600/a_8_216# 0.00fF
C41821 OR2X1_LOC_865/B OR2X1_LOC_392/B 0.18fF
C41822 AND2X1_LOC_794/B AND2X1_LOC_477/a_8_24# 0.01fF
C41823 AND2X1_LOC_539/Y OR2X1_LOC_829/a_36_216# 0.00fF
C41824 AND2X1_LOC_12/Y AND2X1_LOC_91/B 0.13fF
C41825 OR2X1_LOC_696/A OR2X1_LOC_670/a_8_216# 0.01fF
C41826 OR2X1_LOC_160/B OR2X1_LOC_648/A 0.07fF
C41827 AND2X1_LOC_585/a_8_24# OR2X1_LOC_637/B 0.01fF
C41828 AND2X1_LOC_528/a_8_24# AND2X1_LOC_36/Y 0.04fF
C41829 OR2X1_LOC_364/B AND2X1_LOC_40/Y 0.01fF
C41830 OR2X1_LOC_124/A OR2X1_LOC_124/B 0.05fF
C41831 OR2X1_LOC_619/Y OR2X1_LOC_321/a_36_216# 0.01fF
C41832 AND2X1_LOC_64/Y OR2X1_LOC_154/A 0.50fF
C41833 OR2X1_LOC_18/Y OR2X1_LOC_79/a_8_216# 0.05fF
C41834 OR2X1_LOC_198/a_8_216# OR2X1_LOC_269/B 0.01fF
C41835 OR2X1_LOC_738/A AND2X1_LOC_7/B 0.35fF
C41836 OR2X1_LOC_54/Y OR2X1_LOC_150/a_8_216# 0.01fF
C41837 AND2X1_LOC_150/a_36_24# OR2X1_LOC_474/Y 0.01fF
C41838 OR2X1_LOC_125/a_8_216# OR2X1_LOC_91/A 0.03fF
C41839 AND2X1_LOC_658/B AND2X1_LOC_663/A 0.01fF
C41840 OR2X1_LOC_786/Y OR2X1_LOC_598/A 0.19fF
C41841 AND2X1_LOC_555/Y OR2X1_LOC_44/Y 0.04fF
C41842 OR2X1_LOC_178/Y OR2X1_LOC_56/A 0.56fF
C41843 OR2X1_LOC_18/Y AND2X1_LOC_464/A 0.64fF
C41844 AND2X1_LOC_716/Y AND2X1_LOC_182/A 0.14fF
C41845 OR2X1_LOC_573/a_8_216# OR2X1_LOC_244/Y 0.01fF
C41846 OR2X1_LOC_516/Y OR2X1_LOC_74/A 0.53fF
C41847 AND2X1_LOC_95/Y OR2X1_LOC_35/A 0.01fF
C41848 OR2X1_LOC_739/A OR2X1_LOC_161/B 0.03fF
C41849 OR2X1_LOC_379/a_8_216# OR2X1_LOC_691/Y 0.01fF
C41850 OR2X1_LOC_402/B OR2X1_LOC_78/A 0.38fF
C41851 AND2X1_LOC_789/a_8_24# OR2X1_LOC_6/B 0.05fF
C41852 OR2X1_LOC_335/Y AND2X1_LOC_70/Y 0.10fF
C41853 AND2X1_LOC_561/a_36_24# AND2X1_LOC_489/Y 0.00fF
C41854 OR2X1_LOC_6/B AND2X1_LOC_404/A 0.16fF
C41855 OR2X1_LOC_668/Y AND2X1_LOC_44/Y 0.01fF
C41856 OR2X1_LOC_756/B OR2X1_LOC_562/a_8_216# 0.12fF
C41857 OR2X1_LOC_696/A AND2X1_LOC_554/B 0.01fF
C41858 OR2X1_LOC_369/Y AND2X1_LOC_367/A 0.22fF
C41859 OR2X1_LOC_604/A OR2X1_LOC_92/Y 0.06fF
C41860 OR2X1_LOC_493/Y OR2X1_LOC_374/Y 0.08fF
C41861 AND2X1_LOC_562/B AND2X1_LOC_285/Y 0.00fF
C41862 AND2X1_LOC_719/Y OR2X1_LOC_427/A 0.10fF
C41863 OR2X1_LOC_194/B OR2X1_LOC_596/A 0.01fF
C41864 OR2X1_LOC_45/B OR2X1_LOC_85/A 0.12fF
C41865 OR2X1_LOC_151/A AND2X1_LOC_297/a_8_24# 0.01fF
C41866 OR2X1_LOC_40/Y AND2X1_LOC_841/B 0.03fF
C41867 OR2X1_LOC_326/B AND2X1_LOC_323/a_8_24# 0.05fF
C41868 OR2X1_LOC_528/a_8_216# AND2X1_LOC_573/A 0.01fF
C41869 OR2X1_LOC_256/Y OR2X1_LOC_56/A 0.03fF
C41870 AND2X1_LOC_40/Y AND2X1_LOC_70/Y 0.20fF
C41871 OR2X1_LOC_185/Y OR2X1_LOC_138/A 0.00fF
C41872 OR2X1_LOC_154/A AND2X1_LOC_82/Y 0.00fF
C41873 OR2X1_LOC_147/B OR2X1_LOC_542/B 13.10fF
C41874 AND2X1_LOC_91/B AND2X1_LOC_79/Y 0.03fF
C41875 OR2X1_LOC_696/A OR2X1_LOC_696/Y 0.03fF
C41876 OR2X1_LOC_516/B OR2X1_LOC_59/Y 0.21fF
C41877 OR2X1_LOC_158/A OR2X1_LOC_39/A 0.20fF
C41878 OR2X1_LOC_629/a_36_216# OR2X1_LOC_140/B 0.00fF
C41879 AND2X1_LOC_95/Y OR2X1_LOC_552/B 0.01fF
C41880 OR2X1_LOC_692/Y OR2X1_LOC_36/Y 0.04fF
C41881 OR2X1_LOC_604/A OR2X1_LOC_257/a_8_216# 0.04fF
C41882 AND2X1_LOC_392/A AND2X1_LOC_99/A 0.03fF
C41883 OR2X1_LOC_198/a_36_216# AND2X1_LOC_51/Y 0.03fF
C41884 AND2X1_LOC_64/Y OR2X1_LOC_778/A 0.00fF
C41885 OR2X1_LOC_269/B OR2X1_LOC_161/B 2.69fF
C41886 AND2X1_LOC_707/Y OR2X1_LOC_7/A 0.19fF
C41887 OR2X1_LOC_102/a_8_216# OR2X1_LOC_85/A 0.03fF
C41888 VDD OR2X1_LOC_812/B 0.07fF
C41889 OR2X1_LOC_600/A OR2X1_LOC_250/Y 0.14fF
C41890 AND2X1_LOC_721/Y OR2X1_LOC_280/Y 1.54fF
C41891 AND2X1_LOC_47/Y OR2X1_LOC_181/Y 0.02fF
C41892 OR2X1_LOC_436/Y OR2X1_LOC_112/A 0.00fF
C41893 AND2X1_LOC_610/a_8_24# OR2X1_LOC_16/A 0.01fF
C41894 OR2X1_LOC_862/A OR2X1_LOC_561/Y 0.19fF
C41895 AND2X1_LOC_719/Y AND2X1_LOC_464/a_8_24# 0.26fF
C41896 OR2X1_LOC_599/A OR2X1_LOC_589/A 0.49fF
C41897 OR2X1_LOC_117/a_8_216# OR2X1_LOC_490/Y 0.42fF
C41898 D_INPUT_5 OR2X1_LOC_638/a_8_216# 0.01fF
C41899 AND2X1_LOC_40/Y OR2X1_LOC_703/A 0.03fF
C41900 OR2X1_LOC_528/Y OR2X1_LOC_613/Y 0.87fF
C41901 AND2X1_LOC_47/Y OR2X1_LOC_199/B 0.01fF
C41902 OR2X1_LOC_6/B OR2X1_LOC_204/Y 0.03fF
C41903 AND2X1_LOC_70/Y OR2X1_LOC_537/A 0.06fF
C41904 VDD OR2X1_LOC_237/Y 0.11fF
C41905 AND2X1_LOC_130/a_8_24# OR2X1_LOC_26/Y 0.01fF
C41906 OR2X1_LOC_354/A OR2X1_LOC_840/A 0.05fF
C41907 AND2X1_LOC_56/B OR2X1_LOC_410/Y 0.01fF
C41908 OR2X1_LOC_131/A AND2X1_LOC_361/A 0.11fF
C41909 OR2X1_LOC_502/A AND2X1_LOC_401/Y 0.00fF
C41910 OR2X1_LOC_181/B AND2X1_LOC_179/a_36_24# 0.00fF
C41911 OR2X1_LOC_216/A OR2X1_LOC_721/Y 0.03fF
C41912 AND2X1_LOC_729/Y AND2X1_LOC_657/Y 0.03fF
C41913 OR2X1_LOC_287/A OR2X1_LOC_161/A -0.01fF
C41914 OR2X1_LOC_114/Y OR2X1_LOC_140/A 0.00fF
C41915 OR2X1_LOC_26/Y AND2X1_LOC_778/Y 0.03fF
C41916 AND2X1_LOC_182/A OR2X1_LOC_312/Y 0.07fF
C41917 OR2X1_LOC_158/A AND2X1_LOC_211/B 0.09fF
C41918 OR2X1_LOC_638/B AND2X1_LOC_43/B 0.02fF
C41919 OR2X1_LOC_600/A OR2X1_LOC_36/Y 0.54fF
C41920 AND2X1_LOC_548/Y AND2X1_LOC_807/Y 0.13fF
C41921 AND2X1_LOC_281/a_8_24# OR2X1_LOC_580/B 0.09fF
C41922 OR2X1_LOC_532/B OR2X1_LOC_390/B 0.07fF
C41923 OR2X1_LOC_158/A OR2X1_LOC_429/Y 0.01fF
C41924 AND2X1_LOC_99/a_8_24# OR2X1_LOC_278/Y 0.01fF
C41925 OR2X1_LOC_481/A OR2X1_LOC_12/Y 0.04fF
C41926 D_INPUT_4 AND2X1_LOC_328/a_8_24# 0.10fF
C41927 AND2X1_LOC_50/Y AND2X1_LOC_11/Y 0.08fF
C41928 OR2X1_LOC_51/Y OR2X1_LOC_44/Y 0.22fF
C41929 OR2X1_LOC_314/Y OR2X1_LOC_91/A 0.09fF
C41930 OR2X1_LOC_89/A AND2X1_LOC_778/Y 0.03fF
C41931 AND2X1_LOC_721/Y OR2X1_LOC_22/Y 0.02fF
C41932 OR2X1_LOC_318/B OR2X1_LOC_303/B 0.15fF
C41933 OR2X1_LOC_802/Y OR2X1_LOC_78/B 0.06fF
C41934 AND2X1_LOC_757/a_8_24# OR2X1_LOC_161/A 0.01fF
C41935 AND2X1_LOC_56/B OR2X1_LOC_715/A 0.24fF
C41936 OR2X1_LOC_97/B AND2X1_LOC_92/Y 0.15fF
C41937 AND2X1_LOC_635/a_8_24# OR2X1_LOC_428/A 0.08fF
C41938 OR2X1_LOC_468/Y OR2X1_LOC_78/B 0.04fF
C41939 AND2X1_LOC_595/a_8_24# AND2X1_LOC_42/B 0.01fF
C41940 OR2X1_LOC_284/a_36_216# OR2X1_LOC_269/B 0.00fF
C41941 OR2X1_LOC_501/B AND2X1_LOC_56/B 0.24fF
C41942 OR2X1_LOC_791/B OR2X1_LOC_791/A 0.03fF
C41943 AND2X1_LOC_320/a_36_24# AND2X1_LOC_56/B 0.01fF
C41944 AND2X1_LOC_715/Y OR2X1_LOC_167/Y 0.05fF
C41945 VDD OR2X1_LOC_487/a_8_216# 0.00fF
C41946 AND2X1_LOC_49/a_36_24# OR2X1_LOC_78/B 0.01fF
C41947 AND2X1_LOC_456/B AND2X1_LOC_668/a_8_24# 0.01fF
C41948 OR2X1_LOC_648/A OR2X1_LOC_219/B 0.07fF
C41949 OR2X1_LOC_791/B AND2X1_LOC_40/Y 0.03fF
C41950 OR2X1_LOC_216/A OR2X1_LOC_375/A 0.04fF
C41951 OR2X1_LOC_97/A OR2X1_LOC_648/a_36_216# 0.00fF
C41952 AND2X1_LOC_12/Y OR2X1_LOC_308/a_8_216# 0.01fF
C41953 OR2X1_LOC_682/a_8_216# OR2X1_LOC_91/A 0.01fF
C41954 AND2X1_LOC_118/a_8_24# OR2X1_LOC_78/A 0.01fF
C41955 OR2X1_LOC_406/A OR2X1_LOC_142/Y 0.07fF
C41956 OR2X1_LOC_744/A OR2X1_LOC_585/A 0.14fF
C41957 OR2X1_LOC_3/Y AND2X1_LOC_447/Y 0.00fF
C41958 OR2X1_LOC_852/B AND2X1_LOC_824/B 0.00fF
C41959 OR2X1_LOC_80/A OR2X1_LOC_399/a_8_216# 0.06fF
C41960 OR2X1_LOC_856/A AND2X1_LOC_48/A 0.02fF
C41961 OR2X1_LOC_130/A OR2X1_LOC_775/a_36_216# 0.01fF
C41962 OR2X1_LOC_241/B OR2X1_LOC_776/A 0.09fF
C41963 AND2X1_LOC_12/Y AND2X1_LOC_421/a_36_24# 0.00fF
C41964 AND2X1_LOC_784/A AND2X1_LOC_733/Y 0.07fF
C41965 OR2X1_LOC_369/Y OR2X1_LOC_74/A -0.03fF
C41966 AND2X1_LOC_857/Y AND2X1_LOC_354/B 0.03fF
C41967 OR2X1_LOC_45/B OR2X1_LOC_226/Y 0.06fF
C41968 OR2X1_LOC_631/B OR2X1_LOC_294/a_36_216# 0.01fF
C41969 OR2X1_LOC_313/Y OR2X1_LOC_427/A 0.01fF
C41970 OR2X1_LOC_496/Y AND2X1_LOC_734/Y 0.01fF
C41971 AND2X1_LOC_48/a_8_24# OR2X1_LOC_269/B 0.01fF
C41972 OR2X1_LOC_517/A OR2X1_LOC_26/Y 0.40fF
C41973 OR2X1_LOC_427/A AND2X1_LOC_467/a_36_24# 0.00fF
C41974 OR2X1_LOC_606/Y OR2X1_LOC_646/B 0.01fF
C41975 OR2X1_LOC_71/Y OR2X1_LOC_12/Y 0.03fF
C41976 OR2X1_LOC_617/Y AND2X1_LOC_629/a_8_24# 0.23fF
C41977 OR2X1_LOC_147/B AND2X1_LOC_56/B 0.06fF
C41978 OR2X1_LOC_824/Y AND2X1_LOC_839/a_8_24# 0.02fF
C41979 OR2X1_LOC_160/A OR2X1_LOC_377/A 0.07fF
C41980 AND2X1_LOC_340/Y OR2X1_LOC_31/Y 0.03fF
C41981 OR2X1_LOC_131/Y OR2X1_LOC_91/A 0.03fF
C41982 AND2X1_LOC_841/a_8_24# OR2X1_LOC_428/A 0.06fF
C41983 OR2X1_LOC_135/Y AND2X1_LOC_831/Y 0.10fF
C41984 OR2X1_LOC_246/A AND2X1_LOC_243/Y 0.07fF
C41985 OR2X1_LOC_619/Y AND2X1_LOC_466/a_8_24# 0.00fF
C41986 VDD AND2X1_LOC_27/a_8_24# 0.00fF
C41987 AND2X1_LOC_40/Y AND2X1_LOC_17/Y 0.01fF
C41988 OR2X1_LOC_756/B OR2X1_LOC_333/B 0.04fF
C41989 AND2X1_LOC_349/B OR2X1_LOC_517/A 0.01fF
C41990 OR2X1_LOC_517/A OR2X1_LOC_89/A 0.26fF
C41991 AND2X1_LOC_811/Y AND2X1_LOC_727/B 0.02fF
C41992 OR2X1_LOC_9/Y D_INPUT_0 0.10fF
C41993 OR2X1_LOC_315/Y OR2X1_LOC_237/Y 0.05fF
C41994 OR2X1_LOC_105/Y OR2X1_LOC_287/B 0.03fF
C41995 OR2X1_LOC_756/B OR2X1_LOC_850/A 0.03fF
C41996 OR2X1_LOC_317/A AND2X1_LOC_56/B 0.05fF
C41997 AND2X1_LOC_476/A OR2X1_LOC_16/A 0.16fF
C41998 AND2X1_LOC_807/Y AND2X1_LOC_811/a_8_24# 0.05fF
C41999 AND2X1_LOC_181/Y OR2X1_LOC_31/Y 0.11fF
C42000 OR2X1_LOC_36/Y OR2X1_LOC_619/Y 0.18fF
C42001 OR2X1_LOC_484/Y OR2X1_LOC_64/Y 0.70fF
C42002 OR2X1_LOC_757/A OR2X1_LOC_665/a_36_216# 0.00fF
C42003 OR2X1_LOC_160/A OR2X1_LOC_203/Y 0.07fF
C42004 AND2X1_LOC_324/a_36_24# OR2X1_LOC_91/A 0.00fF
C42005 AND2X1_LOC_61/Y AND2X1_LOC_633/Y 0.07fF
C42006 OR2X1_LOC_656/B OR2X1_LOC_99/Y 0.24fF
C42007 AND2X1_LOC_536/a_8_24# OR2X1_LOC_269/B 0.01fF
C42008 AND2X1_LOC_540/a_36_24# OR2X1_LOC_485/A 0.00fF
C42009 OR2X1_LOC_485/A AND2X1_LOC_851/A 0.10fF
C42010 OR2X1_LOC_124/a_36_216# OR2X1_LOC_814/A 0.01fF
C42011 AND2X1_LOC_866/A OR2X1_LOC_322/Y 0.07fF
C42012 AND2X1_LOC_841/B OR2X1_LOC_7/A 9.11fF
C42013 AND2X1_LOC_653/B AND2X1_LOC_653/a_8_24# 0.19fF
C42014 OR2X1_LOC_511/Y AND2X1_LOC_834/a_8_24# 0.01fF
C42015 OR2X1_LOC_503/A AND2X1_LOC_576/Y 0.01fF
C42016 OR2X1_LOC_47/Y OR2X1_LOC_524/a_8_216# 0.01fF
C42017 OR2X1_LOC_851/a_36_216# OR2X1_LOC_814/A 0.01fF
C42018 AND2X1_LOC_59/Y OR2X1_LOC_643/A 0.00fF
C42019 OR2X1_LOC_84/B OR2X1_LOC_185/A 0.35fF
C42020 OR2X1_LOC_846/a_8_216# OR2X1_LOC_269/B 0.01fF
C42021 OR2X1_LOC_865/Y OR2X1_LOC_866/a_8_216# 0.39fF
C42022 AND2X1_LOC_7/B OR2X1_LOC_451/B 0.08fF
C42023 OR2X1_LOC_389/A OR2X1_LOC_532/B 0.01fF
C42024 OR2X1_LOC_329/B OR2X1_LOC_268/a_8_216# 0.02fF
C42025 OR2X1_LOC_117/Y OR2X1_LOC_67/A 0.01fF
C42026 OR2X1_LOC_687/Y OR2X1_LOC_685/a_8_216# 0.04fF
C42027 OR2X1_LOC_814/A AND2X1_LOC_92/Y 0.26fF
C42028 OR2X1_LOC_493/a_8_216# OR2X1_LOC_532/B 0.01fF
C42029 AND2X1_LOC_59/Y OR2X1_LOC_778/Y 0.09fF
C42030 OR2X1_LOC_539/A OR2X1_LOC_193/A 0.01fF
C42031 AND2X1_LOC_748/a_8_24# AND2X1_LOC_3/Y 0.08fF
C42032 OR2X1_LOC_571/Y OR2X1_LOC_576/a_8_216# 0.03fF
C42033 OR2X1_LOC_806/a_8_216# OR2X1_LOC_807/a_8_216# 0.47fF
C42034 AND2X1_LOC_388/a_36_24# AND2X1_LOC_661/A 0.00fF
C42035 AND2X1_LOC_675/Y AND2X1_LOC_657/a_8_24# 0.18fF
C42036 AND2X1_LOC_64/Y OR2X1_LOC_560/A 0.03fF
C42037 AND2X1_LOC_196/Y OR2X1_LOC_59/Y 0.08fF
C42038 OR2X1_LOC_380/A OR2X1_LOC_26/Y 0.01fF
C42039 OR2X1_LOC_128/B AND2X1_LOC_3/Y 0.00fF
C42040 OR2X1_LOC_377/A AND2X1_LOC_86/B 0.07fF
C42041 OR2X1_LOC_89/A AND2X1_LOC_624/A 0.03fF
C42042 OR2X1_LOC_655/B OR2X1_LOC_78/B 0.01fF
C42043 OR2X1_LOC_61/Y OR2X1_LOC_215/A 0.03fF
C42044 OR2X1_LOC_667/a_8_216# OR2X1_LOC_44/Y 0.05fF
C42045 OR2X1_LOC_599/A OR2X1_LOC_43/A 0.03fF
C42046 OR2X1_LOC_158/a_36_216# OR2X1_LOC_158/B 0.01fF
C42047 OR2X1_LOC_248/a_8_216# OR2X1_LOC_248/Y 0.00fF
C42048 OR2X1_LOC_131/Y AND2X1_LOC_573/A 0.11fF
C42049 OR2X1_LOC_158/Y OR2X1_LOC_163/Y 0.09fF
C42050 OR2X1_LOC_3/Y AND2X1_LOC_448/Y 0.00fF
C42051 AND2X1_LOC_675/Y OR2X1_LOC_504/Y 0.00fF
C42052 OR2X1_LOC_377/A OR2X1_LOC_624/B 0.14fF
C42053 OR2X1_LOC_824/Y AND2X1_LOC_839/B 0.02fF
C42054 AND2X1_LOC_224/a_8_24# OR2X1_LOC_68/B 0.02fF
C42055 AND2X1_LOC_76/Y AND2X1_LOC_523/Y 0.32fF
C42056 OR2X1_LOC_488/a_8_216# OR2X1_LOC_18/Y 0.13fF
C42057 AND2X1_LOC_134/a_8_24# OR2X1_LOC_721/Y 0.23fF
C42058 AND2X1_LOC_191/Y OR2X1_LOC_189/A 0.03fF
C42059 OR2X1_LOC_325/a_36_216# OR2X1_LOC_121/B 0.00fF
C42060 AND2X1_LOC_548/Y OR2X1_LOC_95/Y 0.26fF
C42061 AND2X1_LOC_688/a_8_24# AND2X1_LOC_472/B 0.05fF
C42062 AND2X1_LOC_318/Y OR2X1_LOC_56/A 0.20fF
C42063 OR2X1_LOC_756/B OR2X1_LOC_443/a_8_216# 0.01fF
C42064 AND2X1_LOC_308/a_8_24# OR2X1_LOC_48/B 0.01fF
C42065 OR2X1_LOC_619/Y OR2X1_LOC_65/a_8_216# 0.04fF
C42066 AND2X1_LOC_866/A OR2X1_LOC_297/A 0.01fF
C42067 OR2X1_LOC_474/Y D_INPUT_0 0.07fF
C42068 AND2X1_LOC_387/B AND2X1_LOC_56/B 0.03fF
C42069 AND2X1_LOC_711/Y OR2X1_LOC_189/A 0.03fF
C42070 AND2X1_LOC_62/a_8_24# OR2X1_LOC_54/Y 0.04fF
C42071 OR2X1_LOC_22/Y OR2X1_LOC_586/Y 0.03fF
C42072 OR2X1_LOC_364/A OR2X1_LOC_479/Y 0.39fF
C42073 OR2X1_LOC_539/A D_INPUT_0 0.01fF
C42074 OR2X1_LOC_70/Y OR2X1_LOC_189/A 0.06fF
C42075 OR2X1_LOC_185/Y OR2X1_LOC_479/Y 0.03fF
C42076 OR2X1_LOC_837/Y AND2X1_LOC_462/Y 0.01fF
C42077 OR2X1_LOC_13/B AND2X1_LOC_772/Y 0.07fF
C42078 OR2X1_LOC_275/a_36_216# OR2X1_LOC_39/A 0.00fF
C42079 OR2X1_LOC_47/Y AND2X1_LOC_663/A 0.03fF
C42080 AND2X1_LOC_543/a_36_24# AND2X1_LOC_866/A 0.01fF
C42081 OR2X1_LOC_185/A AND2X1_LOC_518/a_36_24# 0.01fF
C42082 OR2X1_LOC_643/Y OR2X1_LOC_341/Y 0.01fF
C42083 AND2X1_LOC_191/Y AND2X1_LOC_220/Y 0.03fF
C42084 OR2X1_LOC_600/A OR2X1_LOC_419/Y 0.22fF
C42085 OR2X1_LOC_36/Y AND2X1_LOC_201/a_8_24# 0.02fF
C42086 AND2X1_LOC_721/a_36_24# OR2X1_LOC_417/A 0.01fF
C42087 OR2X1_LOC_246/Y OR2X1_LOC_64/Y 0.18fF
C42088 AND2X1_LOC_866/A AND2X1_LOC_866/B 0.07fF
C42089 OR2X1_LOC_851/A AND2X1_LOC_47/Y 0.07fF
C42090 OR2X1_LOC_218/Y OR2X1_LOC_475/B 0.00fF
C42091 OR2X1_LOC_154/A OR2X1_LOC_206/A 0.01fF
C42092 OR2X1_LOC_19/B OR2X1_LOC_130/A 0.04fF
C42093 AND2X1_LOC_576/Y OR2X1_LOC_64/Y 0.10fF
C42094 OR2X1_LOC_297/Y AND2X1_LOC_347/a_8_24# 0.23fF
C42095 AND2X1_LOC_831/Y AND2X1_LOC_520/Y 0.00fF
C42096 OR2X1_LOC_813/A OR2X1_LOC_118/Y 0.02fF
C42097 OR2X1_LOC_471/Y OR2X1_LOC_375/A 0.21fF
C42098 OR2X1_LOC_116/A D_INPUT_0 0.01fF
C42099 OR2X1_LOC_123/B OR2X1_LOC_633/B 0.05fF
C42100 AND2X1_LOC_753/B OR2X1_LOC_200/Y 0.05fF
C42101 OR2X1_LOC_18/Y AND2X1_LOC_270/a_8_24# 0.05fF
C42102 OR2X1_LOC_36/Y OR2X1_LOC_22/A 0.03fF
C42103 OR2X1_LOC_293/a_8_216# OR2X1_LOC_753/A 0.01fF
C42104 OR2X1_LOC_529/Y AND2X1_LOC_830/a_8_24# 0.01fF
C42105 OR2X1_LOC_47/Y OR2X1_LOC_2/Y 0.08fF
C42106 OR2X1_LOC_3/Y AND2X1_LOC_729/B 0.03fF
C42107 OR2X1_LOC_217/Y D_INPUT_0 0.01fF
C42108 OR2X1_LOC_96/B D_INPUT_0 0.00fF
C42109 OR2X1_LOC_70/A OR2X1_LOC_25/Y 1.12fF
C42110 OR2X1_LOC_77/a_8_216# OR2X1_LOC_820/B 0.01fF
C42111 AND2X1_LOC_652/a_8_24# AND2X1_LOC_810/Y 0.07fF
C42112 AND2X1_LOC_7/B AND2X1_LOC_36/Y 11.29fF
C42113 AND2X1_LOC_354/Y AND2X1_LOC_319/a_8_24# 0.20fF
C42114 AND2X1_LOC_228/Y OR2X1_LOC_31/Y 0.04fF
C42115 OR2X1_LOC_624/B AND2X1_LOC_670/a_8_24# -0.00fF
C42116 AND2X1_LOC_56/B OR2X1_LOC_545/B 0.03fF
C42117 AND2X1_LOC_155/Y AND2X1_LOC_156/a_36_24# 0.01fF
C42118 OR2X1_LOC_562/Y OR2X1_LOC_562/a_36_216# 0.00fF
C42119 OR2X1_LOC_475/Y OR2X1_LOC_206/a_8_216# 0.14fF
C42120 OR2X1_LOC_276/B AND2X1_LOC_43/B 0.07fF
C42121 AND2X1_LOC_576/Y OR2X1_LOC_417/A 0.02fF
C42122 AND2X1_LOC_91/B OR2X1_LOC_356/B 1.30fF
C42123 D_INPUT_0 AND2X1_LOC_852/Y 0.01fF
C42124 OR2X1_LOC_506/A OR2X1_LOC_786/Y 0.01fF
C42125 AND2X1_LOC_92/Y OR2X1_LOC_341/a_8_216# 0.01fF
C42126 OR2X1_LOC_403/B OR2X1_LOC_532/B 0.00fF
C42127 VDD OR2X1_LOC_384/Y 0.19fF
C42128 AND2X1_LOC_858/B AND2X1_LOC_657/A 0.10fF
C42129 OR2X1_LOC_91/A AND2X1_LOC_657/A 0.13fF
C42130 OR2X1_LOC_38/a_36_216# D_INPUT_1 0.00fF
C42131 OR2X1_LOC_366/B OR2X1_LOC_363/a_8_216# 0.40fF
C42132 OR2X1_LOC_43/A AND2X1_LOC_866/A 0.10fF
C42133 OR2X1_LOC_31/Y OR2X1_LOC_585/A 0.08fF
C42134 OR2X1_LOC_586/Y OR2X1_LOC_387/a_8_216# 0.01fF
C42135 AND2X1_LOC_7/B OR2X1_LOC_334/A 0.21fF
C42136 OR2X1_LOC_563/A OR2X1_LOC_556/a_8_216# 0.01fF
C42137 OR2X1_LOC_679/A AND2X1_LOC_147/Y 0.37fF
C42138 OR2X1_LOC_783/A OR2X1_LOC_449/B 0.00fF
C42139 OR2X1_LOC_66/A OR2X1_LOC_580/A 0.00fF
C42140 AND2X1_LOC_22/Y OR2X1_LOC_338/B 0.06fF
C42141 OR2X1_LOC_205/Y OR2X1_LOC_375/A 0.13fF
C42142 OR2X1_LOC_773/Y OR2X1_LOC_774/a_8_216# 0.08fF
C42143 OR2X1_LOC_462/a_36_216# OR2X1_LOC_416/Y 0.00fF
C42144 OR2X1_LOC_755/A OR2X1_LOC_815/A 0.04fF
C42145 AND2X1_LOC_810/A AND2X1_LOC_798/a_8_24# 0.01fF
C42146 OR2X1_LOC_70/Y AND2X1_LOC_196/Y 0.00fF
C42147 OR2X1_LOC_85/A AND2X1_LOC_838/B 0.01fF
C42148 OR2X1_LOC_805/A AND2X1_LOC_72/B 0.03fF
C42149 AND2X1_LOC_111/a_36_24# D_INPUT_0 0.00fF
C42150 VDD OR2X1_LOC_712/B 0.33fF
C42151 OR2X1_LOC_538/A OR2X1_LOC_446/B 0.03fF
C42152 OR2X1_LOC_621/a_8_216# AND2X1_LOC_36/Y 0.01fF
C42153 OR2X1_LOC_415/Y OR2X1_LOC_548/B 0.00fF
C42154 OR2X1_LOC_538/A OR2X1_LOC_303/B 0.00fF
C42155 OR2X1_LOC_22/Y OR2X1_LOC_245/a_36_216# 0.02fF
C42156 OR2X1_LOC_19/B OR2X1_LOC_62/B 0.08fF
C42157 OR2X1_LOC_154/a_8_216# AND2X1_LOC_7/B 0.06fF
C42158 AND2X1_LOC_64/Y OR2X1_LOC_435/A 0.03fF
C42159 OR2X1_LOC_696/A AND2X1_LOC_362/B 0.07fF
C42160 OR2X1_LOC_696/A AND2X1_LOC_476/Y 0.39fF
C42161 OR2X1_LOC_230/a_36_216# OR2X1_LOC_31/Y 0.00fF
C42162 OR2X1_LOC_273/a_8_216# AND2X1_LOC_476/A 0.02fF
C42163 OR2X1_LOC_485/A OR2X1_LOC_10/a_8_216# 0.01fF
C42164 AND2X1_LOC_555/Y OR2X1_LOC_382/A 0.26fF
C42165 OR2X1_LOC_204/Y OR2X1_LOC_598/A 0.01fF
C42166 OR2X1_LOC_49/A OR2X1_LOC_97/A 0.01fF
C42167 AND2X1_LOC_56/B OR2X1_LOC_318/B 5.14fF
C42168 OR2X1_LOC_709/A OR2X1_LOC_138/a_8_216# 0.00fF
C42169 AND2X1_LOC_573/A AND2X1_LOC_657/A 0.16fF
C42170 OR2X1_LOC_347/A OR2X1_LOC_66/A 0.02fF
C42171 OR2X1_LOC_713/A OR2X1_LOC_779/A 0.16fF
C42172 AND2X1_LOC_110/Y OR2X1_LOC_186/a_36_216# 0.00fF
C42173 OR2X1_LOC_267/Y OR2X1_LOC_361/a_8_216# 0.00fF
C42174 OR2X1_LOC_78/A OR2X1_LOC_714/a_8_216# 0.03fF
C42175 OR2X1_LOC_296/Y AND2X1_LOC_72/B 0.35fF
C42176 OR2X1_LOC_185/Y OR2X1_LOC_68/B 0.11fF
C42177 OR2X1_LOC_151/A OR2X1_LOC_576/A 0.01fF
C42178 OR2X1_LOC_158/A OR2X1_LOC_744/Y 0.01fF
C42179 AND2X1_LOC_12/Y OR2X1_LOC_446/B 0.03fF
C42180 OR2X1_LOC_43/Y OR2X1_LOC_13/Y 0.01fF
C42181 AND2X1_LOC_588/B VDD 0.38fF
C42182 OR2X1_LOC_40/Y AND2X1_LOC_231/Y 0.02fF
C42183 AND2X1_LOC_12/Y OR2X1_LOC_303/B 0.03fF
C42184 INPUT_5 INPUT_6 0.06fF
C42185 OR2X1_LOC_177/Y OR2X1_LOC_322/a_36_216# 0.00fF
C42186 AND2X1_LOC_671/a_8_24# D_INPUT_1 0.00fF
C42187 OR2X1_LOC_139/A VDD 0.86fF
C42188 OR2X1_LOC_40/Y AND2X1_LOC_364/a_8_24# 0.02fF
C42189 OR2X1_LOC_802/A OR2X1_LOC_446/B 0.03fF
C42190 OR2X1_LOC_563/a_36_216# OR2X1_LOC_562/A 0.00fF
C42191 AND2X1_LOC_555/Y OR2X1_LOC_292/a_8_216# 0.01fF
C42192 AND2X1_LOC_91/B OR2X1_LOC_168/B 0.13fF
C42193 OR2X1_LOC_66/A AND2X1_LOC_44/Y 0.60fF
C42194 VDD OR2X1_LOC_758/a_8_216# 0.00fF
C42195 OR2X1_LOC_95/Y OR2X1_LOC_96/a_8_216# 0.01fF
C42196 OR2X1_LOC_539/Y OR2X1_LOC_332/a_8_216# 0.01fF
C42197 VDD OR2X1_LOC_522/a_8_216# 0.21fF
C42198 OR2X1_LOC_114/B AND2X1_LOC_248/a_36_24# 0.00fF
C42199 OR2X1_LOC_45/B OR2X1_LOC_51/Y 1.14fF
C42200 OR2X1_LOC_31/Y AND2X1_LOC_645/a_8_24# 0.01fF
C42201 AND2X1_LOC_340/Y AND2X1_LOC_301/a_8_24# 0.03fF
C42202 AND2X1_LOC_354/B OR2X1_LOC_437/A 0.19fF
C42203 OR2X1_LOC_821/Y OR2X1_LOC_822/a_36_216# 0.00fF
C42204 OR2X1_LOC_368/A AND2X1_LOC_270/a_36_24# 0.00fF
C42205 AND2X1_LOC_18/Y OR2X1_LOC_390/A 0.04fF
C42206 OR2X1_LOC_40/Y OR2X1_LOC_589/A 0.11fF
C42207 VDD OR2X1_LOC_740/B 0.03fF
C42208 AND2X1_LOC_368/a_8_24# AND2X1_LOC_7/B 0.01fF
C42209 OR2X1_LOC_177/Y OR2X1_LOC_600/A 0.03fF
C42210 OR2X1_LOC_426/B OR2X1_LOC_12/Y 5.42fF
C42211 OR2X1_LOC_633/a_8_216# AND2X1_LOC_7/B 0.47fF
C42212 OR2X1_LOC_479/Y OR2X1_LOC_578/B 5.87fF
C42213 AND2X1_LOC_207/A OR2X1_LOC_13/Y 0.01fF
C42214 OR2X1_LOC_793/A AND2X1_LOC_41/Y 0.01fF
C42215 AND2X1_LOC_705/Y OR2X1_LOC_600/Y 0.03fF
C42216 OR2X1_LOC_805/A AND2X1_LOC_36/Y 0.16fF
C42217 OR2X1_LOC_308/A OR2X1_LOC_502/A 0.03fF
C42218 OR2X1_LOC_175/Y OR2X1_LOC_808/B 0.09fF
C42219 AND2X1_LOC_765/a_8_24# OR2X1_LOC_78/Y 0.01fF
C42220 OR2X1_LOC_828/a_36_216# OR2X1_LOC_828/Y 0.00fF
C42221 OR2X1_LOC_532/B OR2X1_LOC_493/Y 0.01fF
C42222 OR2X1_LOC_97/A OR2X1_LOC_808/A 0.03fF
C42223 OR2X1_LOC_66/A OR2X1_LOC_719/a_8_216# 0.01fF
C42224 INPUT_0 OR2X1_LOC_16/A 0.03fF
C42225 AND2X1_LOC_787/A OR2X1_LOC_164/Y 0.02fF
C42226 OR2X1_LOC_604/A OR2X1_LOC_600/A 0.23fF
C42227 OR2X1_LOC_860/a_8_216# AND2X1_LOC_91/B 0.00fF
C42228 AND2X1_LOC_758/a_8_24# OR2X1_LOC_600/A 0.01fF
C42229 OR2X1_LOC_472/B OR2X1_LOC_68/B 0.01fF
C42230 OR2X1_LOC_804/B OR2X1_LOC_303/B 0.01fF
C42231 OR2X1_LOC_122/a_8_216# AND2X1_LOC_362/B 0.05fF
C42232 OR2X1_LOC_53/Y OR2X1_LOC_45/Y 0.11fF
C42233 AND2X1_LOC_573/A OR2X1_LOC_503/a_36_216# 0.01fF
C42234 AND2X1_LOC_410/a_8_24# OR2X1_LOC_51/Y 0.01fF
C42235 OR2X1_LOC_158/A AND2X1_LOC_474/A 0.05fF
C42236 OR2X1_LOC_449/B OR2X1_LOC_308/Y 2.67fF
C42237 AND2X1_LOC_530/a_8_24# AND2X1_LOC_401/Y 0.19fF
C42238 OR2X1_LOC_6/B OR2X1_LOC_78/A 0.12fF
C42239 OR2X1_LOC_285/B OR2X1_LOC_366/Y 0.02fF
C42240 OR2X1_LOC_158/A OR2X1_LOC_421/a_8_216# 0.01fF
C42241 OR2X1_LOC_703/A OR2X1_LOC_356/A 0.11fF
C42242 OR2X1_LOC_628/a_8_216# OR2X1_LOC_816/A 0.01fF
C42243 OR2X1_LOC_166/Y OR2X1_LOC_40/Y 0.00fF
C42244 OR2X1_LOC_203/Y OR2X1_LOC_130/Y 0.00fF
C42245 OR2X1_LOC_865/B OR2X1_LOC_865/A 2.15fF
C42246 OR2X1_LOC_151/A AND2X1_LOC_41/A 0.07fF
C42247 OR2X1_LOC_177/a_36_216# OR2X1_LOC_438/Y 0.00fF
C42248 OR2X1_LOC_604/A AND2X1_LOC_296/a_8_24# 0.04fF
C42249 OR2X1_LOC_106/a_36_216# AND2X1_LOC_474/A 0.00fF
C42250 AND2X1_LOC_91/B AND2X1_LOC_59/Y 2.41fF
C42251 OR2X1_LOC_343/B OR2X1_LOC_493/Y 0.01fF
C42252 OR2X1_LOC_656/B AND2X1_LOC_22/Y 0.03fF
C42253 AND2X1_LOC_500/Y AND2X1_LOC_658/A 0.03fF
C42254 OR2X1_LOC_450/a_8_216# OR2X1_LOC_467/A 0.01fF
C42255 OR2X1_LOC_216/A OR2X1_LOC_549/A 0.03fF
C42256 OR2X1_LOC_161/A OR2X1_LOC_563/A 0.02fF
C42257 OR2X1_LOC_45/B AND2X1_LOC_642/a_8_24# 0.01fF
C42258 OR2X1_LOC_447/Y OR2X1_LOC_724/A 0.24fF
C42259 AND2X1_LOC_391/Y VDD 0.08fF
C42260 VDD AND2X1_LOC_858/B 0.95fF
C42261 OR2X1_LOC_296/Y AND2X1_LOC_36/Y 0.00fF
C42262 AND2X1_LOC_363/B AND2X1_LOC_363/a_8_24# 0.19fF
C42263 AND2X1_LOC_12/Y OR2X1_LOC_366/B 0.37fF
C42264 VDD OR2X1_LOC_91/A 0.55fF
C42265 AND2X1_LOC_721/Y OR2X1_LOC_39/A 0.03fF
C42266 OR2X1_LOC_508/A OR2X1_LOC_151/A 0.77fF
C42267 OR2X1_LOC_811/A OR2X1_LOC_344/A 0.03fF
C42268 AND2X1_LOC_501/Y AND2X1_LOC_735/Y 0.38fF
C42269 AND2X1_LOC_658/B AND2X1_LOC_675/Y 0.09fF
C42270 VDD OR2X1_LOC_637/Y 0.22fF
C42271 OR2X1_LOC_458/a_8_216# OR2X1_LOC_733/A 0.01fF
C42272 OR2X1_LOC_809/B OR2X1_LOC_78/B 0.14fF
C42273 OR2X1_LOC_858/A AND2X1_LOC_498/a_8_24# 0.13fF
C42274 AND2X1_LOC_564/B AND2X1_LOC_840/B 0.10fF
C42275 AND2X1_LOC_352/a_8_24# OR2X1_LOC_92/Y 0.03fF
C42276 AND2X1_LOC_735/Y AND2X1_LOC_570/Y 0.02fF
C42277 OR2X1_LOC_186/Y OR2X1_LOC_185/A 0.03fF
C42278 OR2X1_LOC_40/Y AND2X1_LOC_544/a_8_24# 0.17fF
C42279 OR2X1_LOC_114/B OR2X1_LOC_736/A 0.01fF
C42280 OR2X1_LOC_18/Y OR2X1_LOC_522/Y 0.12fF
C42281 OR2X1_LOC_40/Y AND2X1_LOC_866/B 0.06fF
C42282 OR2X1_LOC_45/B OR2X1_LOC_680/A 0.18fF
C42283 OR2X1_LOC_40/Y AND2X1_LOC_654/B 0.03fF
C42284 OR2X1_LOC_427/A AND2X1_LOC_475/Y 0.03fF
C42285 OR2X1_LOC_62/B AND2X1_LOC_608/a_8_24# 0.01fF
C42286 AND2X1_LOC_42/B AND2X1_LOC_619/a_36_24# 0.00fF
C42287 OR2X1_LOC_501/B AND2X1_LOC_92/Y 0.01fF
C42288 AND2X1_LOC_42/B AND2X1_LOC_235/a_8_24# 0.01fF
C42289 OR2X1_LOC_105/Y OR2X1_LOC_160/B 0.02fF
C42290 OR2X1_LOC_691/A AND2X1_LOC_824/a_8_24# 0.20fF
C42291 OR2X1_LOC_40/Y OR2X1_LOC_495/Y 0.09fF
C42292 AND2X1_LOC_91/B AND2X1_LOC_495/a_8_24# 0.16fF
C42293 OR2X1_LOC_427/A OR2X1_LOC_382/a_8_216# 0.02fF
C42294 OR2X1_LOC_850/B VDD 0.06fF
C42295 AND2X1_LOC_555/Y OR2X1_LOC_261/Y 0.80fF
C42296 OR2X1_LOC_589/A AND2X1_LOC_644/Y 0.07fF
C42297 OR2X1_LOC_709/A AND2X1_LOC_43/B 0.02fF
C42298 AND2X1_LOC_543/Y OR2X1_LOC_7/A 0.01fF
C42299 OR2X1_LOC_97/A OR2X1_LOC_87/B 0.03fF
C42300 AND2X1_LOC_784/A AND2X1_LOC_804/A 0.05fF
C42301 AND2X1_LOC_144/a_8_24# OR2X1_LOC_147/A 0.01fF
C42302 AND2X1_LOC_339/B AND2X1_LOC_138/a_8_24# 0.01fF
C42303 OR2X1_LOC_135/Y AND2X1_LOC_139/B 0.01fF
C42304 OR2X1_LOC_698/Y OR2X1_LOC_56/A 0.03fF
C42305 AND2X1_LOC_207/a_8_24# AND2X1_LOC_214/A 0.00fF
C42306 AND2X1_LOC_456/B OR2X1_LOC_59/Y 0.05fF
C42307 OR2X1_LOC_49/A OR2X1_LOC_699/a_8_216# 0.01fF
C42308 OR2X1_LOC_121/B OR2X1_LOC_308/Y 0.07fF
C42309 AND2X1_LOC_366/a_8_24# OR2X1_LOC_92/Y 0.01fF
C42310 OR2X1_LOC_213/A OR2X1_LOC_160/Y 0.01fF
C42311 OR2X1_LOC_670/Y OR2X1_LOC_428/A 0.03fF
C42312 OR2X1_LOC_441/Y AND2X1_LOC_443/Y 0.00fF
C42313 OR2X1_LOC_532/B OR2X1_LOC_532/a_8_216# 0.02fF
C42314 AND2X1_LOC_172/a_8_24# OR2X1_LOC_61/Y 0.24fF
C42315 OR2X1_LOC_851/B OR2X1_LOC_375/A 0.01fF
C42316 AND2X1_LOC_715/a_36_24# OR2X1_LOC_428/A 0.01fF
C42317 OR2X1_LOC_482/Y OR2X1_LOC_39/A 0.15fF
C42318 D_INPUT_0 OR2X1_LOC_771/B 0.15fF
C42319 OR2X1_LOC_121/Y AND2X1_LOC_56/B 0.09fF
C42320 AND2X1_LOC_705/Y OR2X1_LOC_591/A 0.02fF
C42321 OR2X1_LOC_604/A OR2X1_LOC_619/Y 0.05fF
C42322 AND2X1_LOC_41/A AND2X1_LOC_67/a_8_24# 0.02fF
C42323 OR2X1_LOC_40/Y AND2X1_LOC_858/a_8_24# 0.14fF
C42324 OR2X1_LOC_441/Y AND2X1_LOC_659/a_36_24# 0.01fF
C42325 AND2X1_LOC_231/Y OR2X1_LOC_7/A 0.03fF
C42326 OR2X1_LOC_158/A OR2X1_LOC_85/A 0.36fF
C42327 OR2X1_LOC_690/A OR2X1_LOC_16/A 0.06fF
C42328 OR2X1_LOC_553/A OR2X1_LOC_719/a_36_216# 0.00fF
C42329 AND2X1_LOC_561/B OR2X1_LOC_427/A 0.03fF
C42330 VDD AND2X1_LOC_573/A 1.84fF
C42331 AND2X1_LOC_725/a_36_24# AND2X1_LOC_448/Y 0.00fF
C42332 D_INPUT_5 AND2X1_LOC_3/a_8_24# 0.01fF
C42333 OR2X1_LOC_523/Y OR2X1_LOC_78/A 0.02fF
C42334 OR2X1_LOC_97/A OR2X1_LOC_33/B 0.01fF
C42335 OR2X1_LOC_151/A OR2X1_LOC_631/B 0.05fF
C42336 AND2X1_LOC_367/A AND2X1_LOC_348/A 0.01fF
C42337 AND2X1_LOC_310/a_8_24# OR2X1_LOC_185/A 0.01fF
C42338 OR2X1_LOC_820/a_8_216# OR2X1_LOC_748/A 0.01fF
C42339 AND2X1_LOC_715/A OR2X1_LOC_316/Y 0.02fF
C42340 OR2X1_LOC_653/Y AND2X1_LOC_20/a_36_24# 0.00fF
C42341 OR2X1_LOC_7/A AND2X1_LOC_770/a_8_24# 0.01fF
C42342 OR2X1_LOC_40/Y AND2X1_LOC_87/a_36_24# 0.00fF
C42343 AND2X1_LOC_70/Y AND2X1_LOC_43/B 0.22fF
C42344 OR2X1_LOC_743/A OR2X1_LOC_12/Y 0.12fF
C42345 OR2X1_LOC_86/Y AND2X1_LOC_243/Y 0.02fF
C42346 OR2X1_LOC_865/B OR2X1_LOC_624/Y 0.02fF
C42347 OR2X1_LOC_856/A AND2X1_LOC_3/Y 0.01fF
C42348 AND2X1_LOC_141/a_8_24# OR2X1_LOC_65/B 0.00fF
C42349 OR2X1_LOC_421/A OR2X1_LOC_433/a_8_216# 0.01fF
C42350 OR2X1_LOC_329/B OR2X1_LOC_109/Y 0.00fF
C42351 OR2X1_LOC_159/a_8_216# OR2X1_LOC_43/A 0.04fF
C42352 OR2X1_LOC_54/Y OR2X1_LOC_415/Y 0.16fF
C42353 OR2X1_LOC_95/Y AND2X1_LOC_750/a_36_24# 0.00fF
C42354 OR2X1_LOC_40/Y OR2X1_LOC_43/A 0.52fF
C42355 OR2X1_LOC_589/A OR2X1_LOC_7/A 0.03fF
C42356 OR2X1_LOC_677/a_8_216# OR2X1_LOC_427/A 0.06fF
C42357 AND2X1_LOC_31/Y OR2X1_LOC_228/Y 0.07fF
C42358 OR2X1_LOC_155/A OR2X1_LOC_596/a_8_216# 0.04fF
C42359 OR2X1_LOC_160/A OR2X1_LOC_78/B 0.34fF
C42360 AND2X1_LOC_362/B OR2X1_LOC_89/a_8_216# 0.01fF
C42361 OR2X1_LOC_860/Y OR2X1_LOC_392/A 0.27fF
C42362 OR2X1_LOC_865/B OR2X1_LOC_391/A 0.01fF
C42363 OR2X1_LOC_7/A OR2X1_LOC_322/Y 0.51fF
C42364 AND2X1_LOC_12/Y OR2X1_LOC_573/a_8_216# 0.02fF
C42365 OR2X1_LOC_303/A OR2X1_LOC_212/A 0.00fF
C42366 AND2X1_LOC_715/A AND2X1_LOC_354/B 0.06fF
C42367 OR2X1_LOC_91/Y OR2X1_LOC_178/Y 0.03fF
C42368 OR2X1_LOC_186/Y OR2X1_LOC_435/Y 0.00fF
C42369 OR2X1_LOC_64/Y AND2X1_LOC_244/A 0.02fF
C42370 AND2X1_LOC_95/Y OR2X1_LOC_837/Y 0.01fF
C42371 AND2X1_LOC_716/Y AND2X1_LOC_723/a_8_24# 0.11fF
C42372 OR2X1_LOC_61/B AND2X1_LOC_58/a_36_24# 0.00fF
C42373 OR2X1_LOC_36/Y AND2X1_LOC_286/a_8_24# 0.02fF
C42374 OR2X1_LOC_783/a_36_216# OR2X1_LOC_712/B 0.00fF
C42375 AND2X1_LOC_40/Y AND2X1_LOC_328/a_36_24# 0.01fF
C42376 OR2X1_LOC_589/A OR2X1_LOC_320/Y 0.14fF
C42377 OR2X1_LOC_121/B AND2X1_LOC_604/a_8_24# 0.01fF
C42378 AND2X1_LOC_573/a_36_24# AND2X1_LOC_735/Y 0.01fF
C42379 OR2X1_LOC_842/a_8_216# OR2X1_LOC_161/A 0.01fF
C42380 AND2X1_LOC_535/a_8_24# OR2X1_LOC_43/A 0.01fF
C42381 AND2X1_LOC_12/Y AND2X1_LOC_3/a_8_24# 0.01fF
C42382 OR2X1_LOC_64/Y OR2X1_LOC_16/A 0.14fF
C42383 VDD OR2X1_LOC_669/Y 0.12fF
C42384 OR2X1_LOC_292/a_36_216# AND2X1_LOC_848/Y 0.01fF
C42385 AND2X1_LOC_60/a_8_24# AND2X1_LOC_48/A 0.05fF
C42386 AND2X1_LOC_504/a_8_24# OR2X1_LOC_502/A 0.01fF
C42387 AND2X1_LOC_81/B OR2X1_LOC_242/a_36_216# 0.00fF
C42388 VDD OR2X1_LOC_208/a_8_216# 0.21fF
C42389 AND2X1_LOC_755/a_8_24# OR2X1_LOC_850/B 0.01fF
C42390 AND2X1_LOC_716/Y AND2X1_LOC_662/B 0.02fF
C42391 OR2X1_LOC_368/a_8_216# OR2X1_LOC_74/A 0.24fF
C42392 INPUT_1 AND2X1_LOC_473/Y 0.00fF
C42393 OR2X1_LOC_626/a_36_216# OR2X1_LOC_627/Y 0.00fF
C42394 AND2X1_LOC_657/Y OR2X1_LOC_52/B 0.06fF
C42395 AND2X1_LOC_217/Y AND2X1_LOC_116/Y 0.00fF
C42396 OR2X1_LOC_468/A OR2X1_LOC_593/A 0.01fF
C42397 OR2X1_LOC_528/Y AND2X1_LOC_578/A 0.07fF
C42398 AND2X1_LOC_95/Y AND2X1_LOC_57/a_8_24# 0.07fF
C42399 OR2X1_LOC_110/a_8_216# AND2X1_LOC_476/A 0.06fF
C42400 OR2X1_LOC_377/A OR2X1_LOC_400/a_8_216# 0.04fF
C42401 AND2X1_LOC_727/A AND2X1_LOC_802/Y 0.01fF
C42402 OR2X1_LOC_532/B OR2X1_LOC_390/a_36_216# -0.00fF
C42403 OR2X1_LOC_154/A OR2X1_LOC_756/B 0.05fF
C42404 AND2X1_LOC_392/A AND2X1_LOC_554/B 0.03fF
C42405 AND2X1_LOC_593/Y OR2X1_LOC_594/Y 0.17fF
C42406 OR2X1_LOC_26/Y AND2X1_LOC_286/a_36_24# 0.00fF
C42407 OR2X1_LOC_828/a_8_216# OR2X1_LOC_828/B 0.03fF
C42408 AND2X1_LOC_98/Y OR2X1_LOC_85/A 0.02fF
C42409 AND2X1_LOC_469/B OR2X1_LOC_52/B 0.03fF
C42410 OR2X1_LOC_246/A OR2X1_LOC_12/Y 0.53fF
C42411 AND2X1_LOC_654/Y AND2X1_LOC_662/B 0.02fF
C42412 OR2X1_LOC_421/A OR2X1_LOC_70/Y 0.05fF
C42413 AND2X1_LOC_564/B OR2X1_LOC_31/Y 0.02fF
C42414 AND2X1_LOC_852/Y OR2X1_LOC_612/Y 0.10fF
C42415 OR2X1_LOC_31/Y OR2X1_LOC_230/Y 0.01fF
C42416 OR2X1_LOC_858/A OR2X1_LOC_287/B 0.05fF
C42417 OR2X1_LOC_519/Y AND2X1_LOC_520/Y 0.12fF
C42418 AND2X1_LOC_91/a_8_24# AND2X1_LOC_47/Y 0.01fF
C42419 AND2X1_LOC_64/Y AND2X1_LOC_813/a_8_24# 0.03fF
C42420 OR2X1_LOC_684/Y OR2X1_LOC_765/a_8_216# 0.39fF
C42421 OR2X1_LOC_31/Y OR2X1_LOC_368/Y 0.01fF
C42422 OR2X1_LOC_235/B OR2X1_LOC_810/A 0.05fF
C42423 AND2X1_LOC_717/B OR2X1_LOC_59/Y 0.11fF
C42424 OR2X1_LOC_83/A OR2X1_LOC_394/a_8_216# 0.01fF
C42425 OR2X1_LOC_426/B OR2X1_LOC_272/Y 0.03fF
C42426 OR2X1_LOC_377/A OR2X1_LOC_847/A 0.03fF
C42427 AND2X1_LOC_81/B OR2X1_LOC_608/a_8_216# 0.01fF
C42428 OR2X1_LOC_833/B OR2X1_LOC_541/B 0.02fF
C42429 AND2X1_LOC_387/B AND2X1_LOC_92/Y 0.00fF
C42430 AND2X1_LOC_95/Y OR2X1_LOC_212/A 0.03fF
C42431 AND2X1_LOC_667/a_8_24# AND2X1_LOC_65/A 0.03fF
C42432 AND2X1_LOC_733/Y OR2X1_LOC_52/B 0.18fF
C42433 VDD OR2X1_LOC_27/Y 0.12fF
C42434 AND2X1_LOC_86/B OR2X1_LOC_78/B 0.12fF
C42435 AND2X1_LOC_717/a_36_24# OR2X1_LOC_18/Y 0.00fF
C42436 OR2X1_LOC_700/Y AND2X1_LOC_847/Y 0.02fF
C42437 OR2X1_LOC_108/Y OR2X1_LOC_64/Y 0.07fF
C42438 OR2X1_LOC_190/A OR2X1_LOC_254/a_8_216# 0.03fF
C42439 OR2X1_LOC_288/A OR2X1_LOC_580/B 0.02fF
C42440 AND2X1_LOC_748/a_8_24# OR2X1_LOC_789/B 0.01fF
C42441 OR2X1_LOC_417/A OR2X1_LOC_16/A 0.03fF
C42442 OR2X1_LOC_619/Y AND2X1_LOC_467/a_8_24# 0.01fF
C42443 OR2X1_LOC_465/Y OR2X1_LOC_553/A 0.03fF
C42444 OR2X1_LOC_40/Y AND2X1_LOC_664/a_8_24# 0.01fF
C42445 AND2X1_LOC_99/A OR2X1_LOC_67/a_8_216# 0.01fF
C42446 OR2X1_LOC_624/B OR2X1_LOC_78/B 0.08fF
C42447 AND2X1_LOC_324/a_8_24# OR2X1_LOC_56/A 0.01fF
C42448 OR2X1_LOC_229/a_8_216# OR2X1_LOC_31/Y 0.00fF
C42449 OR2X1_LOC_524/Y OR2X1_LOC_438/a_36_216# 0.00fF
C42450 AND2X1_LOC_656/Y OR2X1_LOC_595/A 0.08fF
C42451 OR2X1_LOC_493/B AND2X1_LOC_491/a_8_24# 0.01fF
C42452 AND2X1_LOC_652/a_8_24# AND2X1_LOC_653/B 0.00fF
C42453 AND2X1_LOC_593/Y AND2X1_LOC_652/a_36_24# 0.01fF
C42454 OR2X1_LOC_128/B OR2X1_LOC_128/a_8_216# 0.08fF
C42455 AND2X1_LOC_191/B OR2X1_LOC_755/A 0.00fF
C42456 OR2X1_LOC_750/A AND2X1_LOC_18/Y 0.09fF
C42457 OR2X1_LOC_269/Y AND2X1_LOC_7/B 0.01fF
C42458 OR2X1_LOC_663/a_8_216# AND2X1_LOC_47/Y 0.01fF
C42459 OR2X1_LOC_409/B OR2X1_LOC_12/Y 0.03fF
C42460 AND2X1_LOC_566/B D_INPUT_0 0.01fF
C42461 OR2X1_LOC_160/A OR2X1_LOC_375/A 0.10fF
C42462 AND2X1_LOC_95/Y OR2X1_LOC_687/Y 0.00fF
C42463 AND2X1_LOC_81/B OR2X1_LOC_185/A 0.03fF
C42464 OR2X1_LOC_39/Y OR2X1_LOC_3/Y 0.00fF
C42465 AND2X1_LOC_303/B OR2X1_LOC_18/Y 0.39fF
C42466 D_INPUT_5 AND2X1_LOC_21/Y 0.18fF
C42467 OR2X1_LOC_185/A OR2X1_LOC_358/B 0.01fF
C42468 OR2X1_LOC_382/Y AND2X1_LOC_345/Y 0.05fF
C42469 OR2X1_LOC_808/A OR2X1_LOC_605/a_8_216# 0.05fF
C42470 AND2X1_LOC_12/Y AND2X1_LOC_56/B 0.08fF
C42471 AND2X1_LOC_561/a_8_24# AND2X1_LOC_563/Y 0.19fF
C42472 OR2X1_LOC_743/A OR2X1_LOC_422/a_8_216# 0.01fF
C42473 AND2X1_LOC_280/a_8_24# AND2X1_LOC_258/a_8_24# 0.23fF
C42474 OR2X1_LOC_193/Y AND2X1_LOC_43/B 0.01fF
C42475 OR2X1_LOC_720/B OR2X1_LOC_66/A 0.03fF
C42476 AND2X1_LOC_22/a_8_24# AND2X1_LOC_21/Y 0.00fF
C42477 AND2X1_LOC_359/a_36_24# OR2X1_LOC_18/Y 0.00fF
C42478 OR2X1_LOC_756/B OR2X1_LOC_345/A 0.08fF
C42479 OR2X1_LOC_108/Y OR2X1_LOC_417/A 0.07fF
C42480 OR2X1_LOC_185/Y OR2X1_LOC_241/a_8_216# 0.04fF
C42481 AND2X1_LOC_337/B AND2X1_LOC_654/Y 0.33fF
C42482 OR2X1_LOC_11/Y AND2X1_LOC_463/a_8_24# 0.01fF
C42483 AND2X1_LOC_390/B OR2X1_LOC_761/Y 0.02fF
C42484 OR2X1_LOC_401/a_8_216# OR2X1_LOC_78/Y 0.01fF
C42485 OR2X1_LOC_485/A OR2X1_LOC_256/a_8_216# 0.40fF
C42486 OR2X1_LOC_634/A OR2X1_LOC_34/B 0.13fF
C42487 OR2X1_LOC_97/A OR2X1_LOC_374/Y 0.93fF
C42488 AND2X1_LOC_715/A AND2X1_LOC_863/Y 0.03fF
C42489 AND2X1_LOC_45/a_8_24# OR2X1_LOC_706/A 0.20fF
C42490 OR2X1_LOC_467/A OR2X1_LOC_780/A 0.00fF
C42491 AND2X1_LOC_325/a_36_24# OR2X1_LOC_31/Y 0.00fF
C42492 AND2X1_LOC_359/B OR2X1_LOC_44/Y 0.03fF
C42493 OR2X1_LOC_205/Y OR2X1_LOC_549/A 0.27fF
C42494 D_GATE_865 OR2X1_LOC_859/B 0.73fF
C42495 AND2X1_LOC_47/Y OR2X1_LOC_78/A 2.34fF
C42496 OR2X1_LOC_669/a_8_216# OR2X1_LOC_26/Y 0.01fF
C42497 AND2X1_LOC_670/a_8_24# OR2X1_LOC_847/A 0.01fF
C42498 AND2X1_LOC_391/Y OR2X1_LOC_256/A 0.72fF
C42499 AND2X1_LOC_170/B AND2X1_LOC_434/Y 0.00fF
C42500 OR2X1_LOC_167/Y AND2X1_LOC_436/a_8_24# 0.13fF
C42501 OR2X1_LOC_36/Y OR2X1_LOC_232/a_8_216# 0.14fF
C42502 OR2X1_LOC_468/Y OR2X1_LOC_711/A 0.00fF
C42503 OR2X1_LOC_64/Y AND2X1_LOC_661/a_8_24# 0.03fF
C42504 OR2X1_LOC_400/A OR2X1_LOC_557/A 0.00fF
C42505 OR2X1_LOC_624/B OR2X1_LOC_375/A 0.07fF
C42506 AND2X1_LOC_41/a_8_24# OR2X1_LOC_214/B 0.00fF
C42507 OR2X1_LOC_22/Y AND2X1_LOC_641/a_36_24# 0.00fF
C42508 OR2X1_LOC_316/Y OR2X1_LOC_27/a_36_216# 0.00fF
C42509 OR2X1_LOC_43/A OR2X1_LOC_7/A 0.22fF
C42510 OR2X1_LOC_599/A AND2X1_LOC_147/Y 0.14fF
C42511 OR2X1_LOC_449/B OR2X1_LOC_593/A 0.02fF
C42512 OR2X1_LOC_224/Y OR2X1_LOC_56/A 0.01fF
C42513 OR2X1_LOC_377/A AND2X1_LOC_46/a_8_24# 0.01fF
C42514 OR2X1_LOC_251/Y OR2X1_LOC_669/Y 0.01fF
C42515 AND2X1_LOC_364/A OR2X1_LOC_46/A 0.12fF
C42516 AND2X1_LOC_663/a_8_24# AND2X1_LOC_663/A 0.07fF
C42517 AND2X1_LOC_206/Y AND2X1_LOC_206/a_8_24# 0.00fF
C42518 AND2X1_LOC_42/B OR2X1_LOC_87/A 2.63fF
C42519 OR2X1_LOC_527/a_8_216# OR2X1_LOC_419/Y 0.13fF
C42520 AND2X1_LOC_859/Y OR2X1_LOC_74/A 0.20fF
C42521 AND2X1_LOC_56/B AND2X1_LOC_496/a_8_24# 0.01fF
C42522 AND2X1_LOC_709/a_8_24# AND2X1_LOC_792/Y 0.01fF
C42523 INPUT_1 AND2X1_LOC_401/a_8_24# 0.01fF
C42524 AND2X1_LOC_132/a_36_24# OR2X1_LOC_404/Y 0.00fF
C42525 OR2X1_LOC_569/a_8_216# OR2X1_LOC_577/B 0.00fF
C42526 AND2X1_LOC_857/Y OR2X1_LOC_31/Y 0.02fF
C42527 AND2X1_LOC_8/Y AND2X1_LOC_79/Y 0.03fF
C42528 OR2X1_LOC_47/Y OR2X1_LOC_25/Y 0.18fF
C42529 OR2X1_LOC_320/Y OR2X1_LOC_43/A 0.50fF
C42530 INPUT_1 AND2X1_LOC_649/a_8_24# 0.03fF
C42531 OR2X1_LOC_600/A AND2X1_LOC_805/a_8_24# 0.01fF
C42532 OR2X1_LOC_792/Y OR2X1_LOC_286/B 0.03fF
C42533 OR2X1_LOC_312/Y AND2X1_LOC_337/B 0.01fF
C42534 AND2X1_LOC_110/Y OR2X1_LOC_365/B 0.01fF
C42535 OR2X1_LOC_485/A OR2X1_LOC_420/a_8_216# 0.02fF
C42536 AND2X1_LOC_99/A AND2X1_LOC_66/a_8_24# 0.19fF
C42537 OR2X1_LOC_3/Y OR2X1_LOC_106/A 0.00fF
C42538 OR2X1_LOC_844/a_8_216# OR2X1_LOC_810/A 0.13fF
C42539 INPUT_6 AND2X1_LOC_581/a_8_24# 0.03fF
C42540 OR2X1_LOC_256/Y D_INPUT_3 0.03fF
C42541 OR2X1_LOC_628/Y OR2X1_LOC_39/A 0.07fF
C42542 AND2X1_LOC_556/a_8_24# OR2X1_LOC_47/Y 0.02fF
C42543 OR2X1_LOC_421/A OR2X1_LOC_70/A 0.22fF
C42544 AND2X1_LOC_722/a_8_24# AND2X1_LOC_222/Y 0.01fF
C42545 AND2X1_LOC_42/B AND2X1_LOC_19/a_8_24# 0.01fF
C42546 AND2X1_LOC_477/A AND2X1_LOC_652/a_8_24# 0.04fF
C42547 AND2X1_LOC_168/Y OR2X1_LOC_417/A 0.12fF
C42548 OR2X1_LOC_234/Y D_INPUT_1 -0.00fF
C42549 AND2X1_LOC_465/a_36_24# AND2X1_LOC_717/B 0.00fF
C42550 OR2X1_LOC_278/a_36_216# OR2X1_LOC_74/A 0.00fF
C42551 OR2X1_LOC_91/A OR2X1_LOC_67/Y 0.03fF
C42552 OR2X1_LOC_787/B OR2X1_LOC_318/B 0.16fF
C42553 AND2X1_LOC_707/Y OR2X1_LOC_424/Y 0.02fF
C42554 OR2X1_LOC_339/a_8_216# OR2X1_LOC_358/A 0.03fF
C42555 OR2X1_LOC_272/Y OR2X1_LOC_743/A 0.09fF
C42556 OR2X1_LOC_78/A OR2X1_LOC_598/A 0.25fF
C42557 OR2X1_LOC_635/a_8_216# OR2X1_LOC_614/a_8_216# 0.47fF
C42558 OR2X1_LOC_256/A AND2X1_LOC_573/A 0.07fF
C42559 OR2X1_LOC_18/Y AND2X1_LOC_859/B 0.08fF
C42560 AND2X1_LOC_92/Y OR2X1_LOC_318/B 0.05fF
C42561 AND2X1_LOC_566/a_8_24# AND2X1_LOC_514/Y 0.01fF
C42562 OR2X1_LOC_541/A OR2X1_LOC_374/Y 0.20fF
C42563 OR2X1_LOC_40/Y OR2X1_LOC_384/a_8_216# 0.01fF
C42564 AND2X1_LOC_145/a_36_24# OR2X1_LOC_148/A 0.00fF
C42565 AND2X1_LOC_21/a_8_24# AND2X1_LOC_21/Y 0.00fF
C42566 OR2X1_LOC_280/Y AND2X1_LOC_523/Y 0.92fF
C42567 OR2X1_LOC_574/A AND2X1_LOC_491/a_8_24# 0.30fF
C42568 OR2X1_LOC_391/A OR2X1_LOC_493/Y 0.10fF
C42569 AND2X1_LOC_685/a_8_24# OR2X1_LOC_7/A 0.05fF
C42570 OR2X1_LOC_606/Y OR2X1_LOC_99/Y 1.08fF
C42571 OR2X1_LOC_786/Y OR2X1_LOC_737/A 0.10fF
C42572 AND2X1_LOC_47/Y OR2X1_LOC_602/A 0.01fF
C42573 AND2X1_LOC_576/Y OR2X1_LOC_226/a_8_216# 0.02fF
C42574 OR2X1_LOC_464/A OR2X1_LOC_737/a_8_216# 0.01fF
C42575 AND2X1_LOC_64/Y AND2X1_LOC_763/B 1.15fF
C42576 OR2X1_LOC_2/Y OR2X1_LOC_3/B 0.12fF
C42577 AND2X1_LOC_434/Y OR2X1_LOC_331/Y 0.28fF
C42578 OR2X1_LOC_458/B OR2X1_LOC_717/a_36_216# 0.00fF
C42579 AND2X1_LOC_88/a_36_24# OR2X1_LOC_121/B 0.00fF
C42580 AND2X1_LOC_367/a_36_24# OR2X1_LOC_417/A 0.01fF
C42581 D_INPUT_0 OR2X1_LOC_217/a_8_216# 0.02fF
C42582 OR2X1_LOC_660/Y AND2X1_LOC_31/Y 0.09fF
C42583 OR2X1_LOC_202/a_8_216# AND2X1_LOC_51/Y 0.01fF
C42584 OR2X1_LOC_309/Y OR2X1_LOC_437/A 0.01fF
C42585 AND2X1_LOC_36/Y OR2X1_LOC_580/B 0.00fF
C42586 OR2X1_LOC_3/Y OR2X1_LOC_46/A 0.15fF
C42587 OR2X1_LOC_272/Y OR2X1_LOC_246/A 0.03fF
C42588 VDD OR2X1_LOC_558/a_8_216# 0.21fF
C42589 AND2X1_LOC_47/Y OR2X1_LOC_155/A 0.19fF
C42590 OR2X1_LOC_161/B OR2X1_LOC_319/Y 0.01fF
C42591 AND2X1_LOC_463/a_36_24# OR2X1_LOC_408/Y 0.00fF
C42592 AND2X1_LOC_472/B OR2X1_LOC_409/a_8_216# 0.47fF
C42593 AND2X1_LOC_573/A OR2X1_LOC_67/Y 0.07fF
C42594 OR2X1_LOC_840/A OR2X1_LOC_567/a_8_216# 0.31fF
C42595 OR2X1_LOC_743/A AND2X1_LOC_801/B 0.03fF
C42596 AND2X1_LOC_624/A AND2X1_LOC_792/Y 0.07fF
C42597 AND2X1_LOC_621/Y AND2X1_LOC_793/Y 0.07fF
C42598 AND2X1_LOC_785/a_8_24# AND2X1_LOC_721/Y 0.01fF
C42599 OR2X1_LOC_22/Y AND2X1_LOC_523/Y 0.06fF
C42600 OR2X1_LOC_648/B AND2X1_LOC_36/Y 0.01fF
C42601 OR2X1_LOC_703/A OR2X1_LOC_357/A 0.01fF
C42602 OR2X1_LOC_696/A AND2X1_LOC_706/Y 0.01fF
C42603 OR2X1_LOC_121/B OR2X1_LOC_606/a_36_216# 0.02fF
C42604 OR2X1_LOC_3/Y AND2X1_LOC_227/Y 0.05fF
C42605 OR2X1_LOC_744/A OR2X1_LOC_437/A 1.02fF
C42606 OR2X1_LOC_64/Y AND2X1_LOC_687/Y 0.04fF
C42607 OR2X1_LOC_143/a_8_216# OR2X1_LOC_9/Y 0.01fF
C42608 OR2X1_LOC_703/A OR2X1_LOC_367/B 1.56fF
C42609 AND2X1_LOC_121/a_36_24# OR2X1_LOC_13/B 0.01fF
C42610 OR2X1_LOC_97/A OR2X1_LOC_392/B 0.01fF
C42611 OR2X1_LOC_375/A OR2X1_LOC_717/a_8_216# 0.02fF
C42612 AND2X1_LOC_315/a_36_24# OR2X1_LOC_318/B 0.00fF
C42613 OR2X1_LOC_595/A AND2X1_LOC_772/Y 0.62fF
C42614 AND2X1_LOC_564/B AND2X1_LOC_464/A 0.04fF
C42615 AND2X1_LOC_76/Y AND2X1_LOC_203/a_8_24# 0.01fF
C42616 OR2X1_LOC_635/a_8_216# AND2X1_LOC_31/Y 0.01fF
C42617 OR2X1_LOC_650/Y OR2X1_LOC_520/A 0.02fF
C42618 OR2X1_LOC_184/Y AND2X1_LOC_717/B 0.00fF
C42619 AND2X1_LOC_555/Y OR2X1_LOC_158/A 0.05fF
C42620 OR2X1_LOC_158/Y AND2X1_LOC_210/a_8_24# 0.23fF
C42621 OR2X1_LOC_260/Y OR2X1_LOC_345/a_36_216# 0.00fF
C42622 OR2X1_LOC_435/Y OR2X1_LOC_112/B 0.10fF
C42623 AND2X1_LOC_339/Y AND2X1_LOC_351/a_36_24# 0.01fF
C42624 AND2X1_LOC_630/a_8_24# AND2X1_LOC_632/A 0.01fF
C42625 AND2X1_LOC_629/Y AND2X1_LOC_630/a_36_24# 0.01fF
C42626 AND2X1_LOC_477/Y AND2X1_LOC_220/B 0.01fF
C42627 AND2X1_LOC_86/Y OR2X1_LOC_71/A 0.01fF
C42628 OR2X1_LOC_294/Y AND2X1_LOC_248/a_8_24# 0.01fF
C42629 AND2X1_LOC_168/a_36_24# OR2X1_LOC_437/A 0.01fF
C42630 OR2X1_LOC_857/B OR2X1_LOC_853/a_36_216# 0.00fF
C42631 AND2X1_LOC_817/B OR2X1_LOC_68/B 0.01fF
C42632 AND2X1_LOC_381/a_8_24# OR2X1_LOC_80/A 0.02fF
C42633 AND2X1_LOC_12/Y AND2X1_LOC_236/a_8_24# 0.01fF
C42634 OR2X1_LOC_135/a_8_216# OR2X1_LOC_135/Y -0.01fF
C42635 INPUT_3 OR2X1_LOC_71/A 0.01fF
C42636 OR2X1_LOC_186/Y OR2X1_LOC_550/A 0.06fF
C42637 OR2X1_LOC_114/a_8_216# OR2X1_LOC_844/B 0.01fF
C42638 OR2X1_LOC_92/Y AND2X1_LOC_449/a_8_24# 0.02fF
C42639 OR2X1_LOC_268/a_8_216# AND2X1_LOC_476/A 0.04fF
C42640 OR2X1_LOC_69/Y OR2X1_LOC_72/Y 0.02fF
C42641 AND2X1_LOC_40/Y OR2X1_LOC_771/B 0.05fF
C42642 OR2X1_LOC_70/Y AND2X1_LOC_451/a_36_24# 0.00fF
C42643 AND2X1_LOC_857/Y OR2X1_LOC_320/a_8_216# 0.01fF
C42644 INPUT_1 OR2X1_LOC_95/Y 0.80fF
C42645 OR2X1_LOC_278/Y OR2X1_LOC_13/B 0.05fF
C42646 AND2X1_LOC_789/a_8_24# AND2X1_LOC_789/Y 0.00fF
C42647 INPUT_1 OR2X1_LOC_368/A 0.01fF
C42648 AND2X1_LOC_672/a_36_24# OR2X1_LOC_54/Y 0.00fF
C42649 AND2X1_LOC_40/Y OR2X1_LOC_209/A 0.03fF
C42650 AND2X1_LOC_425/a_8_24# OR2X1_LOC_451/B 0.00fF
C42651 OR2X1_LOC_110/a_8_216# INPUT_0 0.00fF
C42652 OR2X1_LOC_666/A OR2X1_LOC_89/Y 0.01fF
C42653 AND2X1_LOC_364/a_36_24# AND2X1_LOC_566/B 0.00fF
C42654 OR2X1_LOC_596/A OR2X1_LOC_713/A 0.02fF
C42655 OR2X1_LOC_234/a_8_216# OR2X1_LOC_54/Y 0.01fF
C42656 D_GATE_662 OR2X1_LOC_113/B 0.01fF
C42657 AND2X1_LOC_538/a_36_24# OR2X1_LOC_12/Y 0.00fF
C42658 OR2X1_LOC_52/B AND2X1_LOC_206/Y 0.01fF
C42659 OR2X1_LOC_755/A AND2X1_LOC_848/A 0.23fF
C42660 OR2X1_LOC_212/a_8_216# OR2X1_LOC_469/B 0.02fF
C42661 AND2X1_LOC_196/Y OR2X1_LOC_47/Y 0.08fF
C42662 OR2X1_LOC_654/A OR2X1_LOC_68/B 0.00fF
C42663 OR2X1_LOC_44/Y OR2X1_LOC_399/a_8_216# 0.06fF
C42664 OR2X1_LOC_190/A AND2X1_LOC_44/Y 0.01fF
C42665 OR2X1_LOC_75/a_8_216# OR2X1_LOC_75/Y 0.12fF
C42666 OR2X1_LOC_246/a_8_216# OR2X1_LOC_150/a_8_216# 0.47fF
C42667 VDD OR2X1_LOC_138/A -0.00fF
C42668 OR2X1_LOC_533/Y OR2X1_LOC_600/A 0.06fF
C42669 AND2X1_LOC_462/B OR2X1_LOC_46/A 0.03fF
C42670 AND2X1_LOC_840/B OR2X1_LOC_437/A 0.05fF
C42671 OR2X1_LOC_691/Y OR2X1_LOC_801/a_36_216# 0.00fF
C42672 OR2X1_LOC_600/A AND2X1_LOC_212/Y 0.08fF
C42673 OR2X1_LOC_196/Y OR2X1_LOC_78/B 0.03fF
C42674 AND2X1_LOC_476/a_36_24# OR2X1_LOC_56/A 0.01fF
C42675 OR2X1_LOC_158/A AND2X1_LOC_346/a_36_24# 0.00fF
C42676 AND2X1_LOC_721/Y AND2X1_LOC_474/A 0.02fF
C42677 OR2X1_LOC_87/Y OR2X1_LOC_771/B 0.05fF
C42678 OR2X1_LOC_814/A AND2X1_LOC_289/a_36_24# 0.02fF
C42679 AND2X1_LOC_787/A AND2X1_LOC_471/Y 0.02fF
C42680 OR2X1_LOC_814/A OR2X1_LOC_339/Y 0.02fF
C42681 OR2X1_LOC_848/A OR2X1_LOC_771/B 0.01fF
C42682 OR2X1_LOC_156/a_8_216# OR2X1_LOC_469/Y 0.05fF
C42683 OR2X1_LOC_502/A OR2X1_LOC_703/a_8_216# 0.03fF
C42684 OR2X1_LOC_76/A AND2X1_LOC_31/Y 0.03fF
C42685 AND2X1_LOC_565/B AND2X1_LOC_476/Y 0.04fF
C42686 OR2X1_LOC_78/A AND2X1_LOC_627/a_36_24# 0.00fF
C42687 OR2X1_LOC_687/a_36_216# AND2X1_LOC_430/B 0.00fF
C42688 AND2X1_LOC_250/a_8_24# OR2X1_LOC_343/B 0.01fF
C42689 AND2X1_LOC_566/B AND2X1_LOC_326/B 0.00fF
C42690 OR2X1_LOC_158/A OR2X1_LOC_51/Y 0.59fF
C42691 AND2X1_LOC_212/A AND2X1_LOC_352/B 0.05fF
C42692 OR2X1_LOC_392/B OR2X1_LOC_475/B 0.05fF
C42693 OR2X1_LOC_151/A OR2X1_LOC_648/A 0.07fF
C42694 AND2X1_LOC_91/B OR2X1_LOC_794/A 0.00fF
C42695 AND2X1_LOC_337/B OR2X1_LOC_13/B 0.01fF
C42696 AND2X1_LOC_566/B AND2X1_LOC_337/a_36_24# 0.00fF
C42697 OR2X1_LOC_294/a_8_216# OR2X1_LOC_161/B 0.01fF
C42698 OR2X1_LOC_375/A OR2X1_LOC_130/Y 0.01fF
C42699 OR2X1_LOC_22/a_8_216# D_INPUT_6 0.02fF
C42700 AND2X1_LOC_50/Y AND2X1_LOC_44/Y 0.03fF
C42701 OR2X1_LOC_756/B OR2X1_LOC_435/A 0.00fF
C42702 AND2X1_LOC_22/Y OR2X1_LOC_785/B 0.22fF
C42703 OR2X1_LOC_298/a_8_216# OR2X1_LOC_12/Y 0.05fF
C42704 OR2X1_LOC_240/B OR2X1_LOC_415/Y 0.05fF
C42705 AND2X1_LOC_712/a_8_24# OR2X1_LOC_92/Y 0.01fF
C42706 AND2X1_LOC_357/A OR2X1_LOC_56/A 0.03fF
C42707 AND2X1_LOC_595/a_36_24# OR2X1_LOC_66/A 0.00fF
C42708 AND2X1_LOC_362/B AND2X1_LOC_366/A 0.01fF
C42709 OR2X1_LOC_526/Y AND2X1_LOC_658/A 0.03fF
C42710 OR2X1_LOC_482/a_8_216# AND2X1_LOC_861/B 0.01fF
C42711 AND2X1_LOC_738/B AND2X1_LOC_731/Y 0.02fF
C42712 OR2X1_LOC_600/a_8_216# OR2X1_LOC_600/Y -0.00fF
C42713 OR2X1_LOC_858/A OR2X1_LOC_160/B 0.02fF
C42714 OR2X1_LOC_154/A OR2X1_LOC_140/B 0.03fF
C42715 OR2X1_LOC_158/A OR2X1_LOC_58/a_8_216# 0.05fF
C42716 OR2X1_LOC_490/a_8_216# OR2X1_LOC_92/Y 0.04fF
C42717 OR2X1_LOC_811/A OR2X1_LOC_161/B 0.03fF
C42718 OR2X1_LOC_176/Y OR2X1_LOC_619/Y 0.02fF
C42719 OR2X1_LOC_36/Y AND2X1_LOC_783/B 0.00fF
C42720 AND2X1_LOC_362/a_8_24# VDD 0.00fF
C42721 OR2X1_LOC_436/Y AND2X1_LOC_31/Y 0.03fF
C42722 OR2X1_LOC_516/Y OR2X1_LOC_239/Y 0.04fF
C42723 AND2X1_LOC_42/B OR2X1_LOC_844/B 0.00fF
C42724 OR2X1_LOC_158/A OR2X1_LOC_16/Y 0.03fF
C42725 OR2X1_LOC_19/B OR2X1_LOC_13/B 0.09fF
C42726 AND2X1_LOC_624/A OR2X1_LOC_816/A 0.06fF
C42727 OR2X1_LOC_533/Y OR2X1_LOC_619/Y 0.06fF
C42728 OR2X1_LOC_87/A AND2X1_LOC_224/a_8_24# 0.01fF
C42729 OR2X1_LOC_244/A OR2X1_LOC_71/A 0.02fF
C42730 OR2X1_LOC_696/A OR2X1_LOC_485/A 0.27fF
C42731 OR2X1_LOC_507/a_8_216# OR2X1_LOC_507/A 0.04fF
C42732 OR2X1_LOC_619/Y AND2X1_LOC_212/Y 0.02fF
C42733 AND2X1_LOC_22/Y OR2X1_LOC_687/Y 0.03fF
C42734 AND2X1_LOC_95/Y OR2X1_LOC_535/A 0.01fF
C42735 OR2X1_LOC_833/Y OR2X1_LOC_185/A 0.00fF
C42736 OR2X1_LOC_405/A OR2X1_LOC_185/a_36_216# 0.00fF
C42737 OR2X1_LOC_51/Y AND2X1_LOC_98/Y 0.01fF
C42738 AND2X1_LOC_700/a_8_24# OR2X1_LOC_808/B 0.07fF
C42739 OR2X1_LOC_538/A AND2X1_LOC_92/Y 0.03fF
C42740 OR2X1_LOC_11/Y INPUT_7 0.07fF
C42741 OR2X1_LOC_203/a_36_216# OR2X1_LOC_344/A 0.00fF
C42742 OR2X1_LOC_160/A OR2X1_LOC_549/A 0.14fF
C42743 OR2X1_LOC_70/Y AND2X1_LOC_439/a_36_24# 0.00fF
C42744 AND2X1_LOC_720/Y OR2X1_LOC_51/Y 0.01fF
C42745 OR2X1_LOC_3/Y OR2X1_LOC_748/a_8_216# 0.01fF
C42746 OR2X1_LOC_121/B OR2X1_LOC_301/a_8_216# 0.01fF
C42747 OR2X1_LOC_800/a_36_216# OR2X1_LOC_691/Y 0.00fF
C42748 OR2X1_LOC_52/B AND2X1_LOC_804/A 0.02fF
C42749 AND2X1_LOC_352/a_8_24# OR2X1_LOC_619/Y 0.05fF
C42750 OR2X1_LOC_31/Y OR2X1_LOC_437/A 0.07fF
C42751 OR2X1_LOC_51/Y OR2X1_LOC_594/Y 0.04fF
C42752 AND2X1_LOC_737/Y AND2X1_LOC_657/Y 0.03fF
C42753 AND2X1_LOC_59/Y OR2X1_LOC_719/B 0.02fF
C42754 AND2X1_LOC_47/Y OR2X1_LOC_515/a_36_216# 0.02fF
C42755 INPUT_0 AND2X1_LOC_126/a_8_24# 0.02fF
C42756 OR2X1_LOC_778/A OR2X1_LOC_140/B 0.00fF
C42757 AND2X1_LOC_763/a_8_24# OR2X1_LOC_637/A 0.01fF
C42758 AND2X1_LOC_715/Y OR2X1_LOC_485/A 0.00fF
C42759 OR2X1_LOC_333/B OR2X1_LOC_174/a_36_216# 0.03fF
C42760 OR2X1_LOC_26/Y AND2X1_LOC_786/Y 0.07fF
C42761 OR2X1_LOC_45/B OR2X1_LOC_423/a_8_216# 0.02fF
C42762 AND2X1_LOC_95/Y AND2X1_LOC_323/a_8_24# 0.07fF
C42763 AND2X1_LOC_724/A OR2X1_LOC_601/Y 0.12fF
C42764 AND2X1_LOC_776/a_36_24# AND2X1_LOC_486/Y 0.01fF
C42765 AND2X1_LOC_313/a_8_24# OR2X1_LOC_732/B 0.01fF
C42766 AND2X1_LOC_486/Y AND2X1_LOC_858/B 0.10fF
C42767 OR2X1_LOC_319/B AND2X1_LOC_167/a_8_24# 0.06fF
C42768 OR2X1_LOC_351/a_8_216# OR2X1_LOC_228/Y 0.13fF
C42769 AND2X1_LOC_738/B OR2X1_LOC_48/B 0.26fF
C42770 OR2X1_LOC_56/A OR2X1_LOC_48/B 0.15fF
C42771 OR2X1_LOC_348/Y OR2X1_LOC_791/B 0.01fF
C42772 OR2X1_LOC_18/Y AND2X1_LOC_806/a_36_24# 0.00fF
C42773 OR2X1_LOC_256/Y OR2X1_LOC_494/a_8_216# 0.01fF
C42774 OR2X1_LOC_89/A AND2X1_LOC_786/Y 0.07fF
C42775 OR2X1_LOC_251/a_8_216# OR2X1_LOC_517/A 0.01fF
C42776 VDD OR2X1_LOC_32/B 0.11fF
C42777 OR2X1_LOC_668/Y AND2X1_LOC_18/Y 0.02fF
C42778 AND2X1_LOC_765/a_36_24# OR2X1_LOC_401/Y 0.00fF
C42779 OR2X1_LOC_711/B OR2X1_LOC_469/a_8_216# 0.01fF
C42780 OR2X1_LOC_600/A OR2X1_LOC_265/Y 0.39fF
C42781 OR2X1_LOC_18/Y OR2X1_LOC_56/A 4.63fF
C42782 AND2X1_LOC_723/Y AND2X1_LOC_716/Y 0.03fF
C42783 OR2X1_LOC_434/a_8_216# OR2X1_LOC_436/B -0.00fF
C42784 OR2X1_LOC_847/A OR2X1_LOC_78/B 0.03fF
C42785 OR2X1_LOC_447/A OR2X1_LOC_78/B 0.16fF
C42786 OR2X1_LOC_604/A OR2X1_LOC_669/A 0.29fF
C42787 OR2X1_LOC_187/a_8_216# AND2X1_LOC_866/B 0.03fF
C42788 OR2X1_LOC_506/A OR2X1_LOC_78/A 0.07fF
C42789 AND2X1_LOC_702/a_36_24# OR2X1_LOC_56/A 0.00fF
C42790 OR2X1_LOC_54/Y OR2X1_LOC_397/a_36_216# 0.00fF
C42791 AND2X1_LOC_796/Y OR2X1_LOC_142/Y 0.04fF
C42792 OR2X1_LOC_229/Y OR2X1_LOC_12/Y 0.06fF
C42793 OR2X1_LOC_357/a_8_216# OR2X1_LOC_479/Y 0.05fF
C42794 OR2X1_LOC_346/a_8_216# VDD 0.21fF
C42795 AND2X1_LOC_70/Y OR2X1_LOC_510/Y 0.06fF
C42796 VDD OR2X1_LOC_465/a_8_216# 0.21fF
C42797 AND2X1_LOC_12/Y AND2X1_LOC_92/Y 0.14fF
C42798 OR2X1_LOC_154/A OR2X1_LOC_851/a_8_216# 0.04fF
C42799 AND2X1_LOC_469/Y AND2X1_LOC_220/Y 0.16fF
C42800 AND2X1_LOC_40/Y OR2X1_LOC_637/B 0.03fF
C42801 OR2X1_LOC_604/A AND2X1_LOC_818/a_8_24# 0.03fF
C42802 OR2X1_LOC_161/A OR2X1_LOC_632/Y 0.24fF
C42803 AND2X1_LOC_556/a_8_24# OR2X1_LOC_625/Y 0.04fF
C42804 OR2X1_LOC_643/A OR2X1_LOC_507/A 0.03fF
C42805 AND2X1_LOC_110/Y OR2X1_LOC_449/B 0.03fF
C42806 OR2X1_LOC_160/A OR2X1_LOC_113/Y 0.01fF
C42807 OR2X1_LOC_316/Y AND2X1_LOC_222/a_8_24# 0.00fF
C42808 AND2X1_LOC_82/a_8_24# OR2X1_LOC_78/A 0.01fF
C42809 OR2X1_LOC_377/A OR2X1_LOC_78/Y 0.02fF
C42810 OR2X1_LOC_528/a_8_216# OR2X1_LOC_74/A 0.03fF
C42811 OR2X1_LOC_633/B OR2X1_LOC_786/a_36_216# 0.00fF
C42812 OR2X1_LOC_295/a_8_216# OR2X1_LOC_428/A 0.14fF
C42813 OR2X1_LOC_604/A AND2X1_LOC_454/A 0.25fF
C42814 AND2X1_LOC_24/a_8_24# OR2X1_LOC_130/A 0.14fF
C42815 AND2X1_LOC_436/Y OR2X1_LOC_44/Y 0.03fF
C42816 AND2X1_LOC_570/Y OR2X1_LOC_36/Y 0.03fF
C42817 AND2X1_LOC_40/Y AND2X1_LOC_11/Y 0.01fF
C42818 OR2X1_LOC_58/Y OR2X1_LOC_32/Y 0.80fF
C42819 AND2X1_LOC_553/A OR2X1_LOC_427/A 0.00fF
C42820 OR2X1_LOC_506/B OR2X1_LOC_508/Y 0.02fF
C42821 OR2X1_LOC_18/Y AND2X1_LOC_638/Y 0.05fF
C42822 OR2X1_LOC_40/Y AND2X1_LOC_240/Y 0.00fF
C42823 OR2X1_LOC_64/Y OR2X1_LOC_373/Y 0.02fF
C42824 OR2X1_LOC_499/B OR2X1_LOC_499/a_8_216# 0.07fF
C42825 OR2X1_LOC_685/B OR2X1_LOC_78/B 0.11fF
C42826 OR2X1_LOC_40/Y AND2X1_LOC_147/Y 0.03fF
C42827 AND2X1_LOC_722/a_8_24# OR2X1_LOC_74/A 0.01fF
C42828 AND2X1_LOC_850/A OR2X1_LOC_39/A 0.58fF
C42829 OR2X1_LOC_456/A OR2X1_LOC_344/A 0.20fF
C42830 OR2X1_LOC_557/A OR2X1_LOC_772/A 0.02fF
C42831 AND2X1_LOC_576/Y AND2X1_LOC_663/A 0.10fF
C42832 OR2X1_LOC_841/B AND2X1_LOC_92/Y 0.02fF
C42833 AND2X1_LOC_395/a_8_24# OR2X1_LOC_756/B 0.05fF
C42834 OR2X1_LOC_427/A AND2X1_LOC_804/Y 0.03fF
C42835 AND2X1_LOC_70/Y OR2X1_LOC_810/A 0.08fF
C42836 OR2X1_LOC_492/Y AND2X1_LOC_830/a_8_24# 0.23fF
C42837 AND2X1_LOC_390/a_8_24# AND2X1_LOC_390/B 0.05fF
C42838 AND2X1_LOC_391/Y OR2X1_LOC_248/Y 0.07fF
C42839 AND2X1_LOC_716/a_36_24# OR2X1_LOC_59/Y 0.01fF
C42840 OR2X1_LOC_744/A OR2X1_LOC_753/A 0.21fF
C42841 OR2X1_LOC_479/Y OR2X1_LOC_302/A 0.03fF
C42842 AND2X1_LOC_486/Y AND2X1_LOC_573/A 0.03fF
C42843 OR2X1_LOC_696/A AND2X1_LOC_645/a_36_24# 0.00fF
C42844 OR2X1_LOC_91/A OR2X1_LOC_248/Y 0.03fF
C42845 VDD OR2X1_LOC_371/Y 0.00fF
C42846 OR2X1_LOC_3/Y AND2X1_LOC_403/a_8_24# 0.01fF
C42847 AND2X1_LOC_865/a_36_24# AND2X1_LOC_807/Y 0.00fF
C42848 AND2X1_LOC_9/a_8_24# AND2X1_LOC_852/B 0.04fF
C42849 OR2X1_LOC_311/Y OR2X1_LOC_829/A 0.03fF
C42850 OR2X1_LOC_385/Y OR2X1_LOC_56/A 0.08fF
C42851 OR2X1_LOC_479/Y VDD 1.06fF
C42852 OR2X1_LOC_97/A OR2X1_LOC_532/B 1.17fF
C42853 OR2X1_LOC_663/A OR2X1_LOC_87/A 0.01fF
C42854 OR2X1_LOC_18/Y AND2X1_LOC_850/Y 0.40fF
C42855 OR2X1_LOC_133/a_36_216# OR2X1_LOC_46/A 0.00fF
C42856 AND2X1_LOC_509/Y OR2X1_LOC_7/A 0.57fF
C42857 AND2X1_LOC_344/a_8_24# OR2X1_LOC_44/Y 0.03fF
C42858 AND2X1_LOC_571/Y AND2X1_LOC_573/A 0.01fF
C42859 OR2X1_LOC_417/A OR2X1_LOC_373/Y 0.03fF
C42860 AND2X1_LOC_110/Y OR2X1_LOC_121/B 0.06fF
C42861 GATE_811 AND2X1_LOC_220/B 0.03fF
C42862 OR2X1_LOC_427/A OR2X1_LOC_511/Y 0.01fF
C42863 OR2X1_LOC_804/B AND2X1_LOC_92/Y 0.03fF
C42864 AND2X1_LOC_47/Y OR2X1_LOC_706/a_36_216# 0.02fF
C42865 OR2X1_LOC_328/a_8_216# OR2X1_LOC_17/Y 0.00fF
C42866 AND2X1_LOC_510/a_36_24# AND2X1_LOC_474/Y 0.00fF
C42867 OR2X1_LOC_619/Y OR2X1_LOC_265/Y 0.07fF
C42868 AND2X1_LOC_807/Y AND2X1_LOC_624/A 0.07fF
C42869 OR2X1_LOC_6/B OR2X1_LOC_814/A 0.07fF
C42870 AND2X1_LOC_97/a_8_24# OR2X1_LOC_44/Y 0.04fF
C42871 AND2X1_LOC_22/Y OR2X1_LOC_786/Y 0.03fF
C42872 OR2X1_LOC_8/Y OR2X1_LOC_293/a_8_216# 0.00fF
C42873 OR2X1_LOC_318/Y OR2X1_LOC_592/a_8_216# 0.03fF
C42874 OR2X1_LOC_604/A OR2X1_LOC_601/a_36_216# 0.00fF
C42875 AND2X1_LOC_70/a_36_24# AND2X1_LOC_1/Y 0.00fF
C42876 AND2X1_LOC_51/Y OR2X1_LOC_632/Y 0.07fF
C42877 INPUT_4 OR2X1_LOC_11/Y 0.05fF
C42878 AND2X1_LOC_810/A AND2X1_LOC_798/A 0.01fF
C42879 OR2X1_LOC_270/Y OR2X1_LOC_578/a_36_216# 0.00fF
C42880 AND2X1_LOC_59/Y AND2X1_LOC_56/B 0.73fF
C42881 OR2X1_LOC_626/a_36_216# AND2X1_LOC_805/Y 0.00fF
C42882 OR2X1_LOC_6/A AND2X1_LOC_655/A 0.05fF
C42883 AND2X1_LOC_191/B OR2X1_LOC_22/Y 0.07fF
C42884 OR2X1_LOC_214/B AND2X1_LOC_44/Y 0.04fF
C42885 OR2X1_LOC_506/A OR2X1_LOC_155/A 0.17fF
C42886 OR2X1_LOC_666/a_8_216# OR2X1_LOC_417/A 0.15fF
C42887 AND2X1_LOC_675/A AND2X1_LOC_784/a_8_24# 0.04fF
C42888 OR2X1_LOC_116/a_8_216# OR2X1_LOC_510/Y 0.00fF
C42889 OR2X1_LOC_495/a_36_216# OR2X1_LOC_237/Y 0.00fF
C42890 AND2X1_LOC_59/Y AND2X1_LOC_8/Y 1.81fF
C42891 OR2X1_LOC_291/A AND2X1_LOC_852/B 0.42fF
C42892 OR2X1_LOC_807/A OR2X1_LOC_269/B 0.03fF
C42893 OR2X1_LOC_364/A OR2X1_LOC_87/A 0.07fF
C42894 OR2X1_LOC_185/A OR2X1_LOC_574/A 0.04fF
C42895 OR2X1_LOC_276/B AND2X1_LOC_626/a_8_24# 0.01fF
C42896 OR2X1_LOC_160/A OR2X1_LOC_711/A 0.26fF
C42897 AND2X1_LOC_259/Y AND2X1_LOC_847/Y 0.02fF
C42898 AND2X1_LOC_695/a_8_24# OR2X1_LOC_155/A 0.01fF
C42899 OR2X1_LOC_185/Y OR2X1_LOC_87/A 0.07fF
C42900 AND2X1_LOC_345/Y OR2X1_LOC_427/A 0.07fF
C42901 OR2X1_LOC_140/B OR2X1_LOC_560/A 0.02fF
C42902 OR2X1_LOC_81/a_8_216# OR2X1_LOC_6/A 0.01fF
C42903 AND2X1_LOC_795/Y AND2X1_LOC_795/a_8_24# 0.10fF
C42904 AND2X1_LOC_715/A OR2X1_LOC_31/Y 0.01fF
C42905 OR2X1_LOC_756/B OR2X1_LOC_443/Y 0.01fF
C42906 AND2X1_LOC_859/Y AND2X1_LOC_287/Y 0.00fF
C42907 OR2X1_LOC_64/Y OR2X1_LOC_426/A 0.03fF
C42908 OR2X1_LOC_43/A OR2X1_LOC_236/a_8_216# 0.03fF
C42909 AND2X1_LOC_36/Y OR2X1_LOC_367/a_8_216# 0.01fF
C42910 AND2X1_LOC_31/Y OR2X1_LOC_722/B 0.02fF
C42911 AND2X1_LOC_784/A AND2X1_LOC_354/B 0.03fF
C42912 OR2X1_LOC_18/Y AND2X1_LOC_641/Y 0.10fF
C42913 OR2X1_LOC_744/A AND2X1_LOC_845/Y 0.07fF
C42914 OR2X1_LOC_673/A INPUT_2 0.08fF
C42915 OR2X1_LOC_588/Y OR2X1_LOC_44/Y 0.07fF
C42916 AND2X1_LOC_658/A AND2X1_LOC_810/Y 0.03fF
C42917 OR2X1_LOC_421/A OR2X1_LOC_47/Y 0.14fF
C42918 AND2X1_LOC_219/a_8_24# AND2X1_LOC_476/A 0.03fF
C42919 OR2X1_LOC_3/Y AND2X1_LOC_454/Y 0.00fF
C42920 AND2X1_LOC_334/Y AND2X1_LOC_476/A 0.04fF
C42921 AND2X1_LOC_56/B AND2X1_LOC_495/a_8_24# 0.04fF
C42922 OR2X1_LOC_541/A OR2X1_LOC_532/B 0.00fF
C42923 AND2X1_LOC_563/A OR2X1_LOC_47/Y 0.01fF
C42924 AND2X1_LOC_42/B OR2X1_LOC_573/Y 0.01fF
C42925 OR2X1_LOC_70/Y AND2X1_LOC_452/Y 0.03fF
C42926 OR2X1_LOC_241/B OR2X1_LOC_719/a_8_216# 0.51fF
C42927 OR2X1_LOC_856/B OR2X1_LOC_19/B 0.19fF
C42928 AND2X1_LOC_784/Y AND2X1_LOC_795/Y 0.00fF
C42929 AND2X1_LOC_675/A AND2X1_LOC_471/Y 0.04fF
C42930 OR2X1_LOC_481/A AND2X1_LOC_848/Y 0.03fF
C42931 OR2X1_LOC_864/A OR2X1_LOC_287/B 0.03fF
C42932 OR2X1_LOC_827/Y AND2X1_LOC_838/a_8_24# 0.08fF
C42933 AND2X1_LOC_95/Y OR2X1_LOC_436/a_36_216# 0.00fF
C42934 AND2X1_LOC_42/B AND2X1_LOC_29/a_8_24# 0.01fF
C42935 OR2X1_LOC_92/Y D_INPUT_0 0.03fF
C42936 AND2X1_LOC_808/A AND2X1_LOC_657/Y 0.03fF
C42937 AND2X1_LOC_523/Y OR2X1_LOC_39/A 0.01fF
C42938 OR2X1_LOC_78/A OR2X1_LOC_227/Y 0.02fF
C42939 OR2X1_LOC_485/A AND2X1_LOC_359/a_8_24# 0.01fF
C42940 OR2X1_LOC_91/A AND2X1_LOC_660/A 0.03fF
C42941 AND2X1_LOC_46/a_8_24# OR2X1_LOC_375/A 0.02fF
C42942 OR2X1_LOC_78/A OR2X1_LOC_284/B 0.12fF
C42943 AND2X1_LOC_193/a_8_24# AND2X1_LOC_729/B 0.20fF
C42944 AND2X1_LOC_71/a_36_24# AND2X1_LOC_47/Y 0.00fF
C42945 OR2X1_LOC_517/A OR2X1_LOC_95/Y 0.13fF
C42946 AND2X1_LOC_620/Y OR2X1_LOC_56/A 0.11fF
C42947 AND2X1_LOC_808/A AND2X1_LOC_469/B 0.02fF
C42948 OR2X1_LOC_403/B AND2X1_LOC_42/B 0.01fF
C42949 AND2X1_LOC_578/A OR2X1_LOC_26/Y 0.03fF
C42950 OR2X1_LOC_89/Y OR2X1_LOC_13/B 0.02fF
C42951 OR2X1_LOC_391/B OR2X1_LOC_846/B 0.28fF
C42952 OR2X1_LOC_78/A D_INPUT_1 0.10fF
C42953 OR2X1_LOC_3/B OR2X1_LOC_25/Y 0.33fF
C42954 AND2X1_LOC_86/B OR2X1_LOC_401/Y 0.00fF
C42955 OR2X1_LOC_244/B OR2X1_LOC_786/Y 0.02fF
C42956 OR2X1_LOC_646/A OR2X1_LOC_647/A 0.01fF
C42957 OR2X1_LOC_299/Y OR2X1_LOC_7/A 0.00fF
C42958 OR2X1_LOC_335/A AND2X1_LOC_591/a_8_24# 0.01fF
C42959 OR2X1_LOC_557/A AND2X1_LOC_3/Y 0.94fF
C42960 AND2X1_LOC_570/Y OR2X1_LOC_419/Y 0.02fF
C42961 OR2X1_LOC_487/a_8_216# OR2X1_LOC_487/Y -0.00fF
C42962 AND2X1_LOC_456/B OR2X1_LOC_47/Y 0.00fF
C42963 OR2X1_LOC_476/B OR2X1_LOC_358/B 0.02fF
C42964 AND2X1_LOC_833/a_8_24# OR2X1_LOC_95/Y 0.01fF
C42965 OR2X1_LOC_331/A OR2X1_LOC_419/Y 0.01fF
C42966 OR2X1_LOC_409/B OR2X1_LOC_59/a_8_216# 0.01fF
C42967 AND2X1_LOC_578/A OR2X1_LOC_89/A 0.07fF
C42968 OR2X1_LOC_404/Y AND2X1_LOC_159/a_8_24# 0.01fF
C42969 OR2X1_LOC_114/B OR2X1_LOC_736/a_8_216# 0.01fF
C42970 OR2X1_LOC_490/Y OR2X1_LOC_131/Y 0.01fF
C42971 OR2X1_LOC_78/A AND2X1_LOC_48/Y 0.01fF
C42972 OR2X1_LOC_622/a_8_216# AND2X1_LOC_42/B 0.01fF
C42973 D_INPUT_0 OR2X1_LOC_65/B 0.03fF
C42974 AND2X1_LOC_753/a_36_24# AND2X1_LOC_53/Y 0.01fF
C42975 OR2X1_LOC_404/Y OR2X1_LOC_810/A 0.10fF
C42976 AND2X1_LOC_866/B OR2X1_LOC_615/Y 0.02fF
C42977 VDD AND2X1_LOC_222/Y 0.57fF
C42978 AND2X1_LOC_464/A OR2X1_LOC_437/A 0.02fF
C42979 OR2X1_LOC_814/A OR2X1_LOC_579/B 0.08fF
C42980 OR2X1_LOC_3/Y AND2X1_LOC_847/a_8_24# 0.01fF
C42981 AND2X1_LOC_476/A AND2X1_LOC_649/B 0.02fF
C42982 OR2X1_LOC_784/B OR2X1_LOC_779/B 0.01fF
C42983 OR2X1_LOC_160/B AND2X1_LOC_31/Y 0.45fF
C42984 OR2X1_LOC_427/A AND2X1_LOC_451/Y 0.08fF
C42985 AND2X1_LOC_18/Y OR2X1_LOC_344/a_8_216# 0.14fF
C42986 VDD OR2X1_LOC_562/Y 0.09fF
C42987 OR2X1_LOC_124/B OR2X1_LOC_560/A 0.00fF
C42988 OR2X1_LOC_485/A AND2X1_LOC_663/B 0.27fF
C42989 VDD OR2X1_LOC_68/B 1.42fF
C42990 AND2X1_LOC_227/Y AND2X1_LOC_113/Y 0.01fF
C42991 OR2X1_LOC_161/B OR2X1_LOC_777/B 0.10fF
C42992 OR2X1_LOC_95/Y AND2X1_LOC_624/A 0.03fF
C42993 AND2X1_LOC_22/Y OR2X1_LOC_199/B 0.01fF
C42994 OR2X1_LOC_394/a_8_216# OR2X1_LOC_598/A 0.09fF
C42995 OR2X1_LOC_237/Y OR2X1_LOC_238/a_36_216# 0.00fF
C42996 INPUT_3 AND2X1_LOC_14/a_8_24# 0.01fF
C42997 AND2X1_LOC_535/a_8_24# OR2X1_LOC_534/Y 0.09fF
C42998 OR2X1_LOC_535/A OR2X1_LOC_788/B 0.08fF
C42999 AND2X1_LOC_7/a_8_24# AND2X1_LOC_7/Y 0.01fF
C43000 OR2X1_LOC_323/A OR2X1_LOC_111/a_8_216# 0.01fF
C43001 AND2X1_LOC_53/Y OR2X1_LOC_200/a_8_216# 0.02fF
C43002 OR2X1_LOC_235/B OR2X1_LOC_398/Y 0.05fF
C43003 D_INPUT_3 AND2X1_LOC_838/Y 0.02fF
C43004 AND2X1_LOC_53/Y OR2X1_LOC_269/B 0.50fF
C43005 OR2X1_LOC_151/A OR2X1_LOC_112/A 0.03fF
C43006 OR2X1_LOC_97/B AND2X1_LOC_47/Y 0.18fF
C43007 OR2X1_LOC_702/A OR2X1_LOC_196/B 0.01fF
C43008 AND2X1_LOC_514/Y OR2X1_LOC_321/Y 0.23fF
C43009 VDD OR2X1_LOC_423/Y 0.44fF
C43010 OR2X1_LOC_654/a_8_216# OR2X1_LOC_771/B 0.33fF
C43011 AND2X1_LOC_555/Y AND2X1_LOC_562/a_8_24# 0.01fF
C43012 OR2X1_LOC_31/Y OR2X1_LOC_753/A 0.29fF
C43013 OR2X1_LOC_436/Y OR2X1_LOC_809/a_8_216# 0.01fF
C43014 OR2X1_LOC_846/B OR2X1_LOC_846/A 0.52fF
C43015 OR2X1_LOC_780/A OR2X1_LOC_155/A 0.01fF
C43016 AND2X1_LOC_367/A AND2X1_LOC_657/A 0.10fF
C43017 OR2X1_LOC_98/A OR2X1_LOC_68/B 0.12fF
C43018 OR2X1_LOC_468/a_36_216# OR2X1_LOC_468/Y 0.00fF
C43019 OR2X1_LOC_831/A OR2X1_LOC_593/B 0.04fF
C43020 OR2X1_LOC_64/Y AND2X1_LOC_849/A 0.01fF
C43021 OR2X1_LOC_619/Y AND2X1_LOC_205/a_8_24# 0.04fF
C43022 OR2X1_LOC_32/B OR2X1_LOC_67/Y 0.02fF
C43023 OR2X1_LOC_619/Y OR2X1_LOC_163/A 0.01fF
C43024 OR2X1_LOC_862/B OR2X1_LOC_580/A 0.00fF
C43025 OR2X1_LOC_223/A OR2X1_LOC_269/B 0.03fF
C43026 AND2X1_LOC_598/a_36_24# OR2X1_LOC_47/Y 0.00fF
C43027 OR2X1_LOC_705/B OR2X1_LOC_739/A 0.01fF
C43028 AND2X1_LOC_537/Y AND2X1_LOC_351/Y 0.00fF
C43029 OR2X1_LOC_130/Y OR2X1_LOC_549/A 0.03fF
C43030 OR2X1_LOC_70/Y OR2X1_LOC_70/a_8_216# -0.00fF
C43031 AND2X1_LOC_566/a_8_24# OR2X1_LOC_47/Y 0.01fF
C43032 AND2X1_LOC_817/B OR2X1_LOC_771/a_36_216# 0.00fF
C43033 OR2X1_LOC_3/Y AND2X1_LOC_866/A 0.08fF
C43034 OR2X1_LOC_382/Y OR2X1_LOC_384/Y 0.08fF
C43035 AND2X1_LOC_141/B AND2X1_LOC_656/Y 0.15fF
C43036 OR2X1_LOC_325/Y OR2X1_LOC_532/Y 0.02fF
C43037 OR2X1_LOC_154/A AND2X1_LOC_699/a_8_24# 0.04fF
C43038 OR2X1_LOC_824/a_8_216# OR2X1_LOC_62/A 0.03fF
C43039 AND2X1_LOC_817/a_36_24# D_INPUT_1 0.00fF
C43040 OR2X1_LOC_831/A AND2X1_LOC_273/a_8_24# 0.12fF
C43041 OR2X1_LOC_496/Y AND2X1_LOC_795/Y 0.09fF
C43042 AND2X1_LOC_849/A OR2X1_LOC_417/A 0.02fF
C43043 OR2X1_LOC_623/B OR2X1_LOC_446/B 0.03fF
C43044 AND2X1_LOC_339/Y AND2X1_LOC_350/B 0.00fF
C43045 AND2X1_LOC_455/B OR2X1_LOC_428/A 0.01fF
C43046 OR2X1_LOC_68/Y OR2X1_LOC_814/A 0.01fF
C43047 AND2X1_LOC_12/Y OR2X1_LOC_561/B 0.30fF
C43048 OR2X1_LOC_70/Y AND2X1_LOC_687/a_8_24# 0.26fF
C43049 OR2X1_LOC_78/A OR2X1_LOC_180/B 0.05fF
C43050 OR2X1_LOC_460/B OR2X1_LOC_460/A 0.28fF
C43051 OR2X1_LOC_604/A AND2X1_LOC_783/B 0.01fF
C43052 OR2X1_LOC_703/B OR2X1_LOC_568/A 0.16fF
C43053 OR2X1_LOC_333/B AND2X1_LOC_289/a_8_24# 0.01fF
C43054 AND2X1_LOC_171/a_8_24# OR2X1_LOC_339/Y 0.24fF
C43055 OR2X1_LOC_794/A OR2X1_LOC_303/B 0.03fF
C43056 OR2X1_LOC_188/Y OR2X1_LOC_719/a_8_216# 0.01fF
C43057 OR2X1_LOC_468/Y OR2X1_LOC_567/a_8_216# 0.01fF
C43058 OR2X1_LOC_820/A AND2X1_LOC_750/a_36_24# 0.01fF
C43059 AND2X1_LOC_47/Y OR2X1_LOC_814/A 0.25fF
C43060 OR2X1_LOC_354/A OR2X1_LOC_532/Y 0.07fF
C43061 OR2X1_LOC_344/A OR2X1_LOC_161/B 0.03fF
C43062 AND2X1_LOC_859/Y AND2X1_LOC_562/Y 0.10fF
C43063 OR2X1_LOC_548/A OR2X1_LOC_548/B 0.04fF
C43064 INPUT_1 AND2X1_LOC_293/a_8_24# 0.03fF
C43065 OR2X1_LOC_421/Y OR2X1_LOC_428/A 0.01fF
C43066 AND2X1_LOC_42/B OR2X1_LOC_493/Y 0.04fF
C43067 OR2X1_LOC_468/Y OR2X1_LOC_568/a_36_216# 0.00fF
C43068 AND2X1_LOC_150/a_8_24# OR2X1_LOC_161/B 0.01fF
C43069 OR2X1_LOC_87/A OR2X1_LOC_578/B 0.03fF
C43070 OR2X1_LOC_546/B OR2X1_LOC_705/B 0.05fF
C43071 AND2X1_LOC_350/Y OR2X1_LOC_289/a_8_216# 0.02fF
C43072 AND2X1_LOC_313/a_8_24# AND2X1_LOC_7/B 0.01fF
C43073 AND2X1_LOC_40/Y OR2X1_LOC_593/B 0.03fF
C43074 OR2X1_LOC_131/Y AND2X1_LOC_647/Y 0.02fF
C43075 AND2X1_LOC_3/a_36_24# INPUT_6 0.00fF
C43076 AND2X1_LOC_520/a_8_24# AND2X1_LOC_326/B 0.01fF
C43077 OR2X1_LOC_756/B OR2X1_LOC_605/Y 0.02fF
C43078 AND2X1_LOC_564/A OR2X1_LOC_679/Y 0.03fF
C43079 OR2X1_LOC_686/A OR2X1_LOC_161/B 0.52fF
C43080 OR2X1_LOC_697/Y OR2X1_LOC_743/Y -0.00fF
C43081 OR2X1_LOC_709/A OR2X1_LOC_715/B 0.11fF
C43082 AND2X1_LOC_229/a_8_24# AND2X1_LOC_18/Y 0.01fF
C43083 AND2X1_LOC_456/Y AND2X1_LOC_657/A 0.01fF
C43084 AND2X1_LOC_721/Y OR2X1_LOC_51/Y 0.03fF
C43085 OR2X1_LOC_132/Y AND2X1_LOC_541/a_8_24# 0.23fF
C43086 OR2X1_LOC_66/A OR2X1_LOC_708/a_8_216# 0.02fF
C43087 OR2X1_LOC_490/Y AND2X1_LOC_657/A 0.09fF
C43088 OR2X1_LOC_74/A AND2X1_LOC_657/A 0.07fF
C43089 OR2X1_LOC_862/a_8_216# OR2X1_LOC_561/Y 0.39fF
C43090 AND2X1_LOC_51/Y OR2X1_LOC_170/Y 0.05fF
C43091 OR2X1_LOC_583/a_36_216# OR2X1_LOC_584/Y 0.00fF
C43092 AND2X1_LOC_64/Y OR2X1_LOC_776/a_36_216# 0.02fF
C43093 AND2X1_LOC_388/Y OR2X1_LOC_40/Y 0.18fF
C43094 AND2X1_LOC_848/Y AND2X1_LOC_789/Y 0.08fF
C43095 OR2X1_LOC_135/Y OR2X1_LOC_426/B 0.29fF
C43096 AND2X1_LOC_41/A OR2X1_LOC_563/A 0.02fF
C43097 OR2X1_LOC_56/A AND2X1_LOC_810/B 0.07fF
C43098 OR2X1_LOC_203/Y OR2X1_LOC_217/A 0.00fF
C43099 OR2X1_LOC_814/A OR2X1_LOC_598/A 0.07fF
C43100 OR2X1_LOC_40/Y AND2X1_LOC_500/B 0.01fF
C43101 OR2X1_LOC_604/A AND2X1_LOC_285/a_36_24# 0.01fF
C43102 AND2X1_LOC_539/Y OR2X1_LOC_92/Y 0.03fF
C43103 AND2X1_LOC_716/Y OR2X1_LOC_136/a_8_216# 0.01fF
C43104 OR2X1_LOC_797/B OR2X1_LOC_797/a_8_216# 0.18fF
C43105 OR2X1_LOC_348/Y OR2X1_LOC_362/A 0.09fF
C43106 OR2X1_LOC_467/B OR2X1_LOC_467/A 0.14fF
C43107 OR2X1_LOC_744/A OR2X1_LOC_323/Y 0.43fF
C43108 AND2X1_LOC_363/a_8_24# OR2X1_LOC_56/A 0.02fF
C43109 OR2X1_LOC_185/Y OR2X1_LOC_579/A 0.23fF
C43110 OR2X1_LOC_431/Y OR2X1_LOC_172/Y 0.11fF
C43111 OR2X1_LOC_161/A OR2X1_LOC_168/Y 0.03fF
C43112 AND2X1_LOC_388/Y AND2X1_LOC_535/a_8_24# 0.01fF
C43113 AND2X1_LOC_181/Y OR2X1_LOC_56/A 0.01fF
C43114 OR2X1_LOC_349/a_8_216# OR2X1_LOC_362/A 0.01fF
C43115 OR2X1_LOC_482/Y OR2X1_LOC_51/Y 1.26fF
C43116 AND2X1_LOC_48/A OR2X1_LOC_641/B 0.04fF
C43117 OR2X1_LOC_866/B OR2X1_LOC_772/B 0.04fF
C43118 OR2X1_LOC_495/Y AND2X1_LOC_242/B 0.01fF
C43119 OR2X1_LOC_763/a_8_216# OR2X1_LOC_428/A 0.05fF
C43120 OR2X1_LOC_715/B AND2X1_LOC_70/Y 0.06fF
C43121 OR2X1_LOC_427/A AND2X1_LOC_465/A 1.68fF
C43122 OR2X1_LOC_478/Y OR2X1_LOC_478/a_8_216# -0.00fF
C43123 AND2X1_LOC_70/Y AND2X1_LOC_626/a_8_24# 0.01fF
C43124 AND2X1_LOC_18/Y OR2X1_LOC_66/A 1.37fF
C43125 OR2X1_LOC_22/Y AND2X1_LOC_203/a_8_24# 0.03fF
C43126 OR2X1_LOC_851/A AND2X1_LOC_22/Y 0.01fF
C43127 AND2X1_LOC_552/a_36_24# OR2X1_LOC_427/A 0.00fF
C43128 OR2X1_LOC_841/A AND2X1_LOC_18/Y 0.10fF
C43129 OR2X1_LOC_254/A OR2X1_LOC_161/B 0.01fF
C43130 OR2X1_LOC_147/a_8_216# AND2X1_LOC_36/Y 0.03fF
C43131 OR2X1_LOC_22/Y AND2X1_LOC_206/Y 0.05fF
C43132 AND2X1_LOC_796/a_8_24# OR2X1_LOC_744/A 0.01fF
C43133 OR2X1_LOC_275/A OR2X1_LOC_13/B 0.03fF
C43134 OR2X1_LOC_186/Y OR2X1_LOC_802/a_8_216# 0.01fF
C43135 OR2X1_LOC_564/A AND2X1_LOC_36/Y 0.14fF
C43136 OR2X1_LOC_364/A OR2X1_LOC_390/B 1.03fF
C43137 OR2X1_LOC_833/Y OR2X1_LOC_833/a_8_216# 0.00fF
C43138 OR2X1_LOC_575/A OR2X1_LOC_161/B 0.01fF
C43139 OR2X1_LOC_6/B OR2X1_LOC_501/B 0.00fF
C43140 OR2X1_LOC_185/Y OR2X1_LOC_390/B 0.07fF
C43141 AND2X1_LOC_64/Y OR2X1_LOC_520/Y 0.05fF
C43142 OR2X1_LOC_216/A AND2X1_LOC_65/A 0.00fF
C43143 OR2X1_LOC_278/Y OR2X1_LOC_428/A 0.02fF
C43144 OR2X1_LOC_235/B AND2X1_LOC_243/Y 0.00fF
C43145 OR2X1_LOC_494/Y OR2X1_LOC_59/Y 0.03fF
C43146 AND2X1_LOC_662/B OR2X1_LOC_428/A 4.20fF
C43147 AND2X1_LOC_61/Y AND2X1_LOC_219/Y 0.45fF
C43148 OR2X1_LOC_703/A OR2X1_LOC_543/A 0.30fF
C43149 AND2X1_LOC_555/Y OR2X1_LOC_748/A 0.04fF
C43150 OR2X1_LOC_278/Y OR2X1_LOC_595/A 0.00fF
C43151 AND2X1_LOC_21/Y AND2X1_LOC_762/a_8_24# 0.02fF
C43152 AND2X1_LOC_22/Y OR2X1_LOC_828/B 0.03fF
C43153 AND2X1_LOC_721/Y OR2X1_LOC_680/A 0.03fF
C43154 VDD AND2X1_LOC_367/A 3.16fF
C43155 AND2X1_LOC_92/a_8_24# AND2X1_LOC_824/B 0.01fF
C43156 OR2X1_LOC_62/B OR2X1_LOC_140/Y 0.01fF
C43157 VDD OR2X1_LOC_834/a_8_216# 0.21fF
C43158 AND2X1_LOC_40/Y AND2X1_LOC_41/a_8_24# 0.12fF
C43159 OR2X1_LOC_168/B AND2X1_LOC_92/Y 0.08fF
C43160 AND2X1_LOC_540/a_8_24# OR2X1_LOC_600/A 0.01fF
C43161 OR2X1_LOC_502/A INPUT_2 0.03fF
C43162 AND2X1_LOC_22/Y OR2X1_LOC_204/Y 0.03fF
C43163 AND2X1_LOC_861/B AND2X1_LOC_658/A 0.31fF
C43164 AND2X1_LOC_702/Y OR2X1_LOC_321/a_36_216# 0.00fF
C43165 OR2X1_LOC_648/A OR2X1_LOC_174/A 0.05fF
C43166 OR2X1_LOC_631/B OR2X1_LOC_563/A 0.03fF
C43167 OR2X1_LOC_669/a_8_216# AND2X1_LOC_287/B 0.04fF
C43168 OR2X1_LOC_26/Y AND2X1_LOC_202/Y 0.01fF
C43169 OR2X1_LOC_40/Y AND2X1_LOC_364/A 0.15fF
C43170 OR2X1_LOC_151/A OR2X1_LOC_632/A 0.03fF
C43171 OR2X1_LOC_7/A AND2X1_LOC_780/a_36_24# 0.01fF
C43172 OR2X1_LOC_78/B OR2X1_LOC_78/Y 1.43fF
C43173 OR2X1_LOC_856/B AND2X1_LOC_110/Y 0.24fF
C43174 AND2X1_LOC_326/B OR2X1_LOC_92/Y 0.03fF
C43175 OR2X1_LOC_188/Y OR2X1_LOC_465/B 0.01fF
C43176 OR2X1_LOC_814/Y OR2X1_LOC_772/A 0.31fF
C43177 OR2X1_LOC_516/Y AND2X1_LOC_842/B 0.03fF
C43178 OR2X1_LOC_130/A OR2X1_LOC_390/A 0.01fF
C43179 OR2X1_LOC_709/a_36_216# OR2X1_LOC_738/A 0.00fF
C43180 AND2X1_LOC_484/a_8_24# OR2X1_LOC_731/A 0.29fF
C43181 OR2X1_LOC_382/Y OR2X1_LOC_91/A 0.05fF
C43182 OR2X1_LOC_131/A OR2X1_LOC_65/B 0.01fF
C43183 OR2X1_LOC_516/B OR2X1_LOC_484/Y 0.28fF
C43184 AND2X1_LOC_474/A AND2X1_LOC_850/A 0.03fF
C43185 OR2X1_LOC_756/B OR2X1_LOC_634/A 0.02fF
C43186 AND2X1_LOC_141/B AND2X1_LOC_772/Y 1.03fF
C43187 OR2X1_LOC_482/Y OR2X1_LOC_680/A 1.53fF
C43188 OR2X1_LOC_161/A OR2X1_LOC_777/a_36_216# 0.01fF
C43189 OR2X1_LOC_523/Y OR2X1_LOC_244/Y 0.53fF
C43190 OR2X1_LOC_91/A AND2X1_LOC_863/a_36_24# 0.00fF
C43191 OR2X1_LOC_408/a_8_216# INPUT_6 0.02fF
C43192 OR2X1_LOC_78/A OR2X1_LOC_737/A 0.32fF
C43193 AND2X1_LOC_337/B OR2X1_LOC_428/A 0.03fF
C43194 OR2X1_LOC_6/A OR2X1_LOC_382/a_8_216# 0.19fF
C43195 OR2X1_LOC_60/Y OR2X1_LOC_32/B 0.00fF
C43196 OR2X1_LOC_45/Y AND2X1_LOC_434/a_8_24# 0.11fF
C43197 AND2X1_LOC_725/a_36_24# AND2X1_LOC_454/Y 0.00fF
C43198 AND2X1_LOC_719/Y OR2X1_LOC_44/Y 0.03fF
C43199 AND2X1_LOC_401/Y AND2X1_LOC_402/a_8_24# 0.00fF
C43200 GATE_366 AND2X1_LOC_347/B 0.03fF
C43201 INPUT_0 AND2X1_LOC_649/B 0.04fF
C43202 AND2X1_LOC_95/Y OR2X1_LOC_78/A 6.21fF
C43203 OR2X1_LOC_36/Y AND2X1_LOC_606/a_8_24# 0.04fF
C43204 AND2X1_LOC_702/a_8_24# OR2X1_LOC_59/Y 0.02fF
C43205 AND2X1_LOC_657/Y OR2X1_LOC_39/A 0.05fF
C43206 VDD AND2X1_LOC_35/Y 0.21fF
C43207 OR2X1_LOC_633/Y OR2X1_LOC_78/A 6.10fF
C43208 OR2X1_LOC_528/Y AND2X1_LOC_580/B 0.05fF
C43209 OR2X1_LOC_158/A OR2X1_LOC_423/a_8_216# 0.01fF
C43210 OR2X1_LOC_135/Y OR2X1_LOC_743/A 0.07fF
C43211 OR2X1_LOC_92/Y AND2X1_LOC_276/a_8_24# 0.17fF
C43212 AND2X1_LOC_784/A OR2X1_LOC_309/Y 0.05fF
C43213 OR2X1_LOC_458/B OR2X1_LOC_737/A 0.07fF
C43214 AND2X1_LOC_64/Y AND2X1_LOC_107/a_8_24# 0.01fF
C43215 AND2X1_LOC_13/a_8_24# OR2X1_LOC_161/B 0.01fF
C43216 OR2X1_LOC_193/A AND2X1_LOC_44/Y 0.03fF
C43217 AND2X1_LOC_228/Y OR2X1_LOC_56/A 0.09fF
C43218 AND2X1_LOC_59/Y AND2X1_LOC_92/Y 0.31fF
C43219 AND2X1_LOC_469/B OR2X1_LOC_39/A 0.01fF
C43220 OR2X1_LOC_810/A OR2X1_LOC_362/A 0.05fF
C43221 AND2X1_LOC_843/a_36_24# OR2X1_LOC_59/Y 0.00fF
C43222 OR2X1_LOC_174/A OR2X1_LOC_405/a_8_216# 0.47fF
C43223 AND2X1_LOC_720/a_8_24# AND2X1_LOC_456/B 0.01fF
C43224 OR2X1_LOC_244/Y OR2X1_LOC_579/B 0.00fF
C43225 OR2X1_LOC_11/Y OR2X1_LOC_380/Y 0.01fF
C43226 OR2X1_LOC_680/A AND2X1_LOC_188/a_36_24# 0.00fF
C43227 AND2X1_LOC_729/Y OR2X1_LOC_744/A 0.10fF
C43228 OR2X1_LOC_808/B OR2X1_LOC_620/Y 0.10fF
C43229 AND2X1_LOC_707/Y AND2X1_LOC_685/a_8_24# 0.01fF
C43230 AND2X1_LOC_456/B OR2X1_LOC_625/Y 0.07fF
C43231 OR2X1_LOC_185/Y OR2X1_LOC_801/a_8_216# 0.01fF
C43232 OR2X1_LOC_864/A OR2X1_LOC_160/B 0.10fF
C43233 OR2X1_LOC_176/a_36_216# AND2X1_LOC_514/Y 0.00fF
C43234 OR2X1_LOC_160/A OR2X1_LOC_662/a_36_216# 0.00fF
C43235 OR2X1_LOC_141/B OR2X1_LOC_641/A 0.00fF
C43236 AND2X1_LOC_367/A OR2X1_LOC_315/Y 0.40fF
C43237 OR2X1_LOC_49/A OR2X1_LOC_99/B 0.00fF
C43238 AND2X1_LOC_514/a_36_24# AND2X1_LOC_655/A 0.06fF
C43239 AND2X1_LOC_552/A AND2X1_LOC_578/A 0.02fF
C43240 OR2X1_LOC_405/A OR2X1_LOC_840/A 0.27fF
C43241 AND2X1_LOC_653/a_36_24# AND2X1_LOC_436/Y 0.00fF
C43242 AND2X1_LOC_733/Y OR2X1_LOC_39/A 0.01fF
C43243 OR2X1_LOC_652/a_8_216# OR2X1_LOC_435/B 0.01fF
C43244 OR2X1_LOC_274/a_8_216# OR2X1_LOC_375/A 0.01fF
C43245 VDD OR2X1_LOC_757/a_8_216# 0.21fF
C43246 AND2X1_LOC_547/Y AND2X1_LOC_475/a_8_24# 0.01fF
C43247 OR2X1_LOC_40/Y OR2X1_LOC_3/Y 2.56fF
C43248 AND2X1_LOC_81/a_8_24# AND2X1_LOC_70/Y 0.01fF
C43249 AND2X1_LOC_40/Y OR2X1_LOC_812/A 0.01fF
C43250 OR2X1_LOC_189/Y AND2X1_LOC_731/Y 0.03fF
C43251 OR2X1_LOC_502/A OR2X1_LOC_739/A 0.06fF
C43252 VDD AND2X1_LOC_456/Y 0.27fF
C43253 AND2X1_LOC_675/Y AND2X1_LOC_576/Y 0.03fF
C43254 AND2X1_LOC_784/A OR2X1_LOC_744/A 0.07fF
C43255 OR2X1_LOC_175/Y OR2X1_LOC_532/B 0.03fF
C43256 AND2X1_LOC_717/Y OR2X1_LOC_109/Y 0.07fF
C43257 OR2X1_LOC_585/A OR2X1_LOC_56/A 0.16fF
C43258 AND2X1_LOC_639/A AND2X1_LOC_639/B 0.24fF
C43259 OR2X1_LOC_474/Y OR2X1_LOC_510/Y 0.03fF
C43260 OR2X1_LOC_152/Y AND2X1_LOC_731/Y 0.09fF
C43261 VDD OR2X1_LOC_490/Y 0.24fF
C43262 VDD OR2X1_LOC_74/A 1.53fF
C43263 OR2X1_LOC_40/Y AND2X1_LOC_631/Y 0.07fF
C43264 OR2X1_LOC_135/Y OR2X1_LOC_246/A 0.10fF
C43265 VDD AND2X1_LOC_697/a_8_24# -0.00fF
C43266 AND2X1_LOC_208/B AND2X1_LOC_35/Y 0.41fF
C43267 OR2X1_LOC_154/A OR2X1_LOC_808/B 0.10fF
C43268 AND2X1_LOC_197/Y OR2X1_LOC_6/A 0.01fF
C43269 OR2X1_LOC_656/Y OR2X1_LOC_520/Y 0.10fF
C43270 D_INPUT_0 AND2X1_LOC_44/Y 0.31fF
C43271 OR2X1_LOC_8/Y OR2X1_LOC_824/a_8_216# 0.00fF
C43272 AND2X1_LOC_303/B AND2X1_LOC_857/Y 0.00fF
C43273 OR2X1_LOC_319/a_8_216# OR2X1_LOC_185/A 0.05fF
C43274 OR2X1_LOC_178/Y OR2X1_LOC_529/Y 0.37fF
C43275 OR2X1_LOC_7/Y OR2X1_LOC_16/A 0.26fF
C43276 OR2X1_LOC_833/B AND2X1_LOC_72/Y 0.03fF
C43277 OR2X1_LOC_691/Y OR2X1_LOC_532/B 0.01fF
C43278 AND2X1_LOC_52/a_8_24# OR2X1_LOC_87/A 0.01fF
C43279 AND2X1_LOC_769/a_8_24# OR2X1_LOC_744/A 0.01fF
C43280 OR2X1_LOC_251/Y AND2X1_LOC_367/A 0.60fF
C43281 OR2X1_LOC_8/Y OR2X1_LOC_825/a_8_216# 0.02fF
C43282 AND2X1_LOC_515/a_8_24# AND2X1_LOC_477/A 0.01fF
C43283 AND2X1_LOC_76/Y OR2X1_LOC_595/a_36_216# 0.00fF
C43284 OR2X1_LOC_502/A AND2X1_LOC_26/a_8_24# 0.01fF
C43285 OR2X1_LOC_377/A OR2X1_LOC_185/A 0.07fF
C43286 AND2X1_LOC_56/B OR2X1_LOC_623/B 1.47fF
C43287 AND2X1_LOC_357/B AND2X1_LOC_514/Y 0.01fF
C43288 AND2X1_LOC_366/A OR2X1_LOC_485/A 0.03fF
C43289 OR2X1_LOC_91/Y OR2X1_LOC_48/B 0.07fF
C43290 OR2X1_LOC_502/A OR2X1_LOC_269/B 0.50fF
C43291 OR2X1_LOC_64/Y AND2X1_LOC_447/Y 0.02fF
C43292 OR2X1_LOC_502/A AND2X1_LOC_404/a_36_24# 0.01fF
C43293 AND2X1_LOC_362/B AND2X1_LOC_66/a_8_24# 0.01fF
C43294 OR2X1_LOC_95/Y AND2X1_LOC_774/A 0.01fF
C43295 OR2X1_LOC_3/Y OR2X1_LOC_698/a_8_216# 0.01fF
C43296 OR2X1_LOC_31/Y OR2X1_LOC_323/Y 0.04fF
C43297 OR2X1_LOC_91/Y OR2X1_LOC_18/Y 0.03fF
C43298 AND2X1_LOC_36/Y OR2X1_LOC_228/Y 0.04fF
C43299 OR2X1_LOC_415/Y OR2X1_LOC_396/Y 0.02fF
C43300 OR2X1_LOC_405/A OR2X1_LOC_222/A 0.03fF
C43301 OR2X1_LOC_185/Y OR2X1_LOC_865/B 0.01fF
C43302 OR2X1_LOC_116/A OR2X1_LOC_510/Y 0.00fF
C43303 OR2X1_LOC_43/A AND2X1_LOC_841/B 0.03fF
C43304 OR2X1_LOC_305/Y OR2X1_LOC_48/B 0.22fF
C43305 AND2X1_LOC_144/a_8_24# OR2X1_LOC_705/Y 0.02fF
C43306 OR2X1_LOC_677/Y OR2X1_LOC_74/A 0.03fF
C43307 INPUT_0 AND2X1_LOC_729/B 0.04fF
C43308 AND2X1_LOC_160/Y AND2X1_LOC_712/B 0.11fF
C43309 OR2X1_LOC_119/a_36_216# OR2X1_LOC_744/A 0.00fF
C43310 OR2X1_LOC_704/a_8_216# OR2X1_LOC_714/A -0.00fF
C43311 AND2X1_LOC_36/Y OR2X1_LOC_513/Y 0.01fF
C43312 AND2X1_LOC_859/Y AND2X1_LOC_287/a_8_24# 0.20fF
C43313 OR2X1_LOC_51/Y OR2X1_LOC_628/Y 0.02fF
C43314 AND2X1_LOC_720/a_36_24# OR2X1_LOC_26/Y 0.00fF
C43315 OR2X1_LOC_217/Y OR2X1_LOC_510/Y 0.02fF
C43316 OR2X1_LOC_600/A D_INPUT_0 0.10fF
C43317 OR2X1_LOC_91/A AND2X1_LOC_307/Y 0.03fF
C43318 OR2X1_LOC_772/B OR2X1_LOC_557/A 0.00fF
C43319 OR2X1_LOC_36/Y OR2X1_LOC_69/A 0.17fF
C43320 AND2X1_LOC_486/Y OR2X1_LOC_371/Y 0.19fF
C43321 AND2X1_LOC_95/Y OR2X1_LOC_155/A 0.03fF
C43322 AND2X1_LOC_655/A OR2X1_LOC_44/Y 0.00fF
C43323 AND2X1_LOC_116/B OR2X1_LOC_59/Y 0.02fF
C43324 AND2X1_LOC_202/a_8_24# AND2X1_LOC_202/Y 0.01fF
C43325 AND2X1_LOC_842/B AND2X1_LOC_842/a_8_24# 0.05fF
C43326 OR2X1_LOC_814/Y AND2X1_LOC_3/Y 0.12fF
C43327 AND2X1_LOC_86/Y OR2X1_LOC_633/B 0.02fF
C43328 OR2X1_LOC_18/Y OR2X1_LOC_371/a_8_216# 0.01fF
C43329 AND2X1_LOC_12/Y OR2X1_LOC_389/B 0.03fF
C43330 OR2X1_LOC_401/Y OR2X1_LOC_847/A 0.03fF
C43331 OR2X1_LOC_809/a_36_216# OR2X1_LOC_539/Y 0.00fF
C43332 AND2X1_LOC_432/a_8_24# OR2X1_LOC_390/B 0.05fF
C43333 OR2X1_LOC_316/Y OR2X1_LOC_52/B 0.03fF
C43334 OR2X1_LOC_778/Y AND2X1_LOC_272/a_8_24# -0.01fF
C43335 AND2X1_LOC_40/Y OR2X1_LOC_254/a_8_216# 0.01fF
C43336 OR2X1_LOC_502/A OR2X1_LOC_215/A 0.03fF
C43337 AND2X1_LOC_568/B AND2X1_LOC_170/B 0.20fF
C43338 OR2X1_LOC_185/Y OR2X1_LOC_800/a_8_216# 0.01fF
C43339 AND2X1_LOC_702/Y OR2X1_LOC_36/Y 0.04fF
C43340 OR2X1_LOC_74/A AND2X1_LOC_274/a_8_24# 0.05fF
C43341 OR2X1_LOC_81/a_8_216# OR2X1_LOC_44/Y 0.14fF
C43342 OR2X1_LOC_205/Y AND2X1_LOC_65/A 0.15fF
C43343 AND2X1_LOC_784/A AND2X1_LOC_840/B 0.10fF
C43344 OR2X1_LOC_154/A OR2X1_LOC_708/B 0.14fF
C43345 AND2X1_LOC_47/Y OR2X1_LOC_244/Y 0.04fF
C43346 AND2X1_LOC_154/Y AND2X1_LOC_621/Y 0.14fF
C43347 OR2X1_LOC_121/B OR2X1_LOC_448/A 0.11fF
C43348 AND2X1_LOC_155/Y OR2X1_LOC_619/Y 0.16fF
C43349 AND2X1_LOC_508/A AND2X1_LOC_574/A 0.12fF
C43350 OR2X1_LOC_487/Y AND2X1_LOC_573/A 0.01fF
C43351 OR2X1_LOC_242/a_8_216# OR2X1_LOC_532/B 0.01fF
C43352 OR2X1_LOC_820/A INPUT_1 0.12fF
C43353 OR2X1_LOC_315/Y OR2X1_LOC_74/A 0.02fF
C43354 AND2X1_LOC_702/a_8_24# OR2X1_LOC_70/Y 0.04fF
C43355 OR2X1_LOC_84/A AND2X1_LOC_18/Y 0.03fF
C43356 OR2X1_LOC_47/Y AND2X1_LOC_200/a_8_24# 0.17fF
C43357 OR2X1_LOC_92/Y AND2X1_LOC_687/A 0.02fF
C43358 OR2X1_LOC_670/Y OR2X1_LOC_26/Y 0.02fF
C43359 OR2X1_LOC_696/A OR2X1_LOC_385/a_8_216# 0.03fF
C43360 OR2X1_LOC_843/a_8_216# OR2X1_LOC_579/B 0.04fF
C43361 AND2X1_LOC_228/Y AND2X1_LOC_641/Y 0.08fF
C43362 OR2X1_LOC_527/Y OR2X1_LOC_18/Y 0.06fF
C43363 OR2X1_LOC_501/B AND2X1_LOC_47/Y 0.14fF
C43364 OR2X1_LOC_417/Y OR2X1_LOC_48/B 0.07fF
C43365 AND2X1_LOC_365/a_8_24# AND2X1_LOC_863/Y 0.01fF
C43366 OR2X1_LOC_177/Y OR2X1_LOC_406/A 0.00fF
C43367 OR2X1_LOC_137/a_36_216# OR2X1_LOC_532/B 0.00fF
C43368 OR2X1_LOC_329/B AND2X1_LOC_866/A 0.07fF
C43369 AND2X1_LOC_8/Y OR2X1_LOC_585/A 0.08fF
C43370 OR2X1_LOC_109/Y OR2X1_LOC_64/Y 0.13fF
C43371 OR2X1_LOC_215/A AND2X1_LOC_230/a_8_24# 0.01fF
C43372 VDD AND2X1_LOC_460/a_8_24# 0.00fF
C43373 OR2X1_LOC_690/A OR2X1_LOC_24/a_36_216# 0.03fF
C43374 OR2X1_LOC_756/B OR2X1_LOC_439/a_8_216# 0.01fF
C43375 AND2X1_LOC_51/A AND2X1_LOC_44/a_8_24# 0.04fF
C43376 VDD OR2X1_LOC_247/a_8_216# 0.00fF
C43377 OR2X1_LOC_820/A OR2X1_LOC_751/a_8_216# 0.06fF
C43378 OR2X1_LOC_691/B AND2X1_LOC_31/Y 0.08fF
C43379 OR2X1_LOC_377/A AND2X1_LOC_119/a_8_24# 0.00fF
C43380 OR2X1_LOC_494/A OR2X1_LOC_384/Y 0.00fF
C43381 OR2X1_LOC_533/Y OR2X1_LOC_534/a_8_216# 0.01fF
C43382 AND2X1_LOC_738/a_36_24# GATE_811 0.00fF
C43383 OR2X1_LOC_549/B D_GATE_366 0.00fF
C43384 AND2X1_LOC_335/a_8_24# AND2X1_LOC_318/Y 0.17fF
C43385 OR2X1_LOC_181/B OR2X1_LOC_471/Y 0.03fF
C43386 AND2X1_LOC_390/B OR2X1_LOC_52/B 0.07fF
C43387 AND2X1_LOC_56/B AND2X1_LOC_13/a_36_24# 0.00fF
C43388 OR2X1_LOC_160/B OR2X1_LOC_351/a_8_216# 0.01fF
C43389 OR2X1_LOC_147/B AND2X1_LOC_47/Y 0.06fF
C43390 OR2X1_LOC_291/A OR2X1_LOC_585/A 0.04fF
C43391 OR2X1_LOC_3/Y OR2X1_LOC_7/A 6.85fF
C43392 OR2X1_LOC_309/a_36_216# AND2X1_LOC_222/Y 0.00fF
C43393 AND2X1_LOC_64/Y OR2X1_LOC_590/Y 0.10fF
C43394 AND2X1_LOC_383/a_36_24# OR2X1_LOC_437/A 0.00fF
C43395 OR2X1_LOC_417/A AND2X1_LOC_649/B 0.04fF
C43396 VDD AND2X1_LOC_647/Y 0.41fF
C43397 D_INPUT_0 OR2X1_LOC_619/Y 0.08fF
C43398 AND2X1_LOC_729/B OR2X1_LOC_690/A 0.01fF
C43399 OR2X1_LOC_680/A OR2X1_LOC_628/Y 0.07fF
C43400 OR2X1_LOC_59/Y AND2X1_LOC_204/Y 0.02fF
C43401 OR2X1_LOC_109/Y OR2X1_LOC_417/A 0.11fF
C43402 AND2X1_LOC_18/Y OR2X1_LOC_559/a_8_216# 0.02fF
C43403 D_INPUT_3 AND2X1_LOC_852/B 0.01fF
C43404 OR2X1_LOC_778/a_8_216# OR2X1_LOC_493/Y 0.04fF
C43405 AND2X1_LOC_706/Y OR2X1_LOC_589/Y 0.15fF
C43406 AND2X1_LOC_48/A OR2X1_LOC_200/a_8_216# 0.01fF
C43407 OR2X1_LOC_501/B OR2X1_LOC_598/A 0.07fF
C43408 OR2X1_LOC_756/B OR2X1_LOC_366/a_8_216# 0.02fF
C43409 AND2X1_LOC_48/A OR2X1_LOC_269/B 0.49fF
C43410 AND2X1_LOC_729/Y OR2X1_LOC_31/Y 0.01fF
C43411 OR2X1_LOC_743/A AND2X1_LOC_856/B 0.00fF
C43412 AND2X1_LOC_99/Y OR2X1_LOC_813/Y 0.03fF
C43413 OR2X1_LOC_437/a_36_216# OR2X1_LOC_48/B 0.00fF
C43414 OR2X1_LOC_497/Y OR2X1_LOC_226/a_36_216# -0.02fF
C43415 OR2X1_LOC_744/A OR2X1_LOC_88/Y 0.03fF
C43416 OR2X1_LOC_864/A OR2X1_LOC_244/A 0.07fF
C43417 OR2X1_LOC_696/A AND2X1_LOC_715/Y 0.17fF
C43418 OR2X1_LOC_416/A OR2X1_LOC_6/A 0.43fF
C43419 OR2X1_LOC_64/Y AND2X1_LOC_729/B 0.01fF
C43420 AND2X1_LOC_656/Y OR2X1_LOC_26/Y 0.04fF
C43421 INPUT_5 OR2X1_LOC_70/A 0.10fF
C43422 AND2X1_LOC_640/Y AND2X1_LOC_640/a_8_24# 0.01fF
C43423 AND2X1_LOC_574/Y AND2X1_LOC_575/a_8_24# 0.00fF
C43424 OR2X1_LOC_624/A OR2X1_LOC_66/a_8_216# 0.18fF
C43425 OR2X1_LOC_334/B OR2X1_LOC_68/B 0.01fF
C43426 OR2X1_LOC_307/B AND2X1_LOC_31/Y 0.05fF
C43427 AND2X1_LOC_17/Y OR2X1_LOC_639/a_36_216# 0.00fF
C43428 AND2X1_LOC_12/Y OR2X1_LOC_215/a_8_216# 0.01fF
C43429 INPUT_5 AND2X1_LOC_31/Y 0.67fF
C43430 OR2X1_LOC_635/a_8_216# OR2X1_LOC_451/B 0.08fF
C43431 AND2X1_LOC_656/Y OR2X1_LOC_89/A 0.07fF
C43432 AND2X1_LOC_486/Y AND2X1_LOC_222/Y 0.03fF
C43433 OR2X1_LOC_208/A AND2X1_LOC_44/Y 0.00fF
C43434 AND2X1_LOC_633/Y AND2X1_LOC_201/a_8_24# 0.17fF
C43435 OR2X1_LOC_147/A OR2X1_LOC_546/A 0.21fF
C43436 OR2X1_LOC_347/a_36_216# OR2X1_LOC_675/Y 0.02fF
C43437 OR2X1_LOC_289/Y OR2X1_LOC_265/Y 0.03fF
C43438 OR2X1_LOC_323/A OR2X1_LOC_428/A 0.24fF
C43439 AND2X1_LOC_387/B AND2X1_LOC_47/Y 0.01fF
C43440 AND2X1_LOC_497/a_8_24# OR2X1_LOC_161/A 0.01fF
C43441 OR2X1_LOC_490/Y OR2X1_LOC_256/A 0.07fF
C43442 AND2X1_LOC_12/Y OR2X1_LOC_339/Y 0.14fF
C43443 OR2X1_LOC_91/A AND2X1_LOC_212/a_8_24# 0.07fF
C43444 OR2X1_LOC_36/Y OR2X1_LOC_51/B 0.09fF
C43445 AND2X1_LOC_86/Y OR2X1_LOC_608/Y 0.10fF
C43446 AND2X1_LOC_810/a_8_24# AND2X1_LOC_661/A 0.01fF
C43447 OR2X1_LOC_3/a_8_216# OR2X1_LOC_31/Y 0.01fF
C43448 AND2X1_LOC_811/B AND2X1_LOC_222/Y 0.00fF
C43449 AND2X1_LOC_342/a_8_24# AND2X1_LOC_721/A 0.01fF
C43450 AND2X1_LOC_76/Y OR2X1_LOC_153/a_8_216# 0.48fF
C43451 OR2X1_LOC_18/Y AND2X1_LOC_656/a_8_24# 0.02fF
C43452 AND2X1_LOC_60/a_8_24# AND2X1_LOC_7/B 0.01fF
C43453 OR2X1_LOC_78/A OR2X1_LOC_788/B 3.83fF
C43454 AND2X1_LOC_640/a_8_24# OR2X1_LOC_416/Y 0.01fF
C43455 OR2X1_LOC_185/Y OR2X1_LOC_493/Y 0.10fF
C43456 OR2X1_LOC_486/Y OR2X1_LOC_556/a_8_216# 0.01fF
C43457 OR2X1_LOC_185/Y OR2X1_LOC_801/B 0.07fF
C43458 AND2X1_LOC_473/Y AND2X1_LOC_786/Y 0.04fF
C43459 OR2X1_LOC_563/B OR2X1_LOC_549/Y 0.17fF
C43460 OR2X1_LOC_361/a_8_216# OR2X1_LOC_140/B 0.01fF
C43461 OR2X1_LOC_639/a_8_216# AND2X1_LOC_51/Y 0.01fF
C43462 VDD OR2X1_LOC_598/a_8_216# 0.00fF
C43463 AND2X1_LOC_12/Y AND2X1_LOC_751/a_8_24# 0.18fF
C43464 AND2X1_LOC_543/Y OR2X1_LOC_322/Y 0.23fF
C43465 OR2X1_LOC_341/Y OR2X1_LOC_341/a_8_216# -0.00fF
C43466 OR2X1_LOC_611/Y OR2X1_LOC_62/B 0.01fF
C43467 D_GATE_479 OR2X1_LOC_161/B 0.01fF
C43468 OR2X1_LOC_79/Y AND2X1_LOC_786/Y 0.79fF
C43469 AND2X1_LOC_498/a_8_24# AND2X1_LOC_36/Y 0.01fF
C43470 AND2X1_LOC_320/a_8_24# AND2X1_LOC_36/Y 0.10fF
C43471 OR2X1_LOC_39/A AND2X1_LOC_203/a_8_24# 0.01fF
C43472 OR2X1_LOC_532/B OR2X1_LOC_750/a_8_216# 0.01fF
C43473 AND2X1_LOC_338/Y AND2X1_LOC_333/a_36_24# 0.00fF
C43474 AND2X1_LOC_40/Y OR2X1_LOC_580/A 0.00fF
C43475 AND2X1_LOC_652/a_8_24# OR2X1_LOC_533/A 0.20fF
C43476 D_INPUT_0 OR2X1_LOC_720/B -0.02fF
C43477 OR2X1_LOC_74/A AND2X1_LOC_624/B 0.03fF
C43478 OR2X1_LOC_39/A AND2X1_LOC_206/Y 0.00fF
C43479 OR2X1_LOC_490/Y OR2X1_LOC_67/Y 0.01fF
C43480 OR2X1_LOC_74/A OR2X1_LOC_67/Y 0.07fF
C43481 OR2X1_LOC_219/B OR2X1_LOC_351/a_8_216# 0.13fF
C43482 OR2X1_LOC_416/Y AND2X1_LOC_649/Y 0.01fF
C43483 OR2X1_LOC_31/Y AND2X1_LOC_639/A 0.02fF
C43484 OR2X1_LOC_865/a_8_216# OR2X1_LOC_561/B 0.01fF
C43485 OR2X1_LOC_696/A OR2X1_LOC_122/a_8_216# 0.03fF
C43486 AND2X1_LOC_476/A OR2X1_LOC_46/A 0.17fF
C43487 OR2X1_LOC_545/B AND2X1_LOC_47/Y 0.01fF
C43488 AND2X1_LOC_364/a_8_24# OR2X1_LOC_589/A 0.17fF
C43489 OR2X1_LOC_45/B AND2X1_LOC_719/Y 0.01fF
C43490 OR2X1_LOC_812/B OR2X1_LOC_561/A 0.01fF
C43491 OR2X1_LOC_70/Y OR2X1_LOC_311/a_8_216# 0.14fF
C43492 OR2X1_LOC_52/B OR2X1_LOC_153/a_8_216# 0.03fF
C43493 OR2X1_LOC_160/B OR2X1_LOC_121/A 0.06fF
C43494 OR2X1_LOC_673/Y OR2X1_LOC_80/A 0.09fF
C43495 OR2X1_LOC_186/Y OR2X1_LOC_550/a_8_216# 0.18fF
C43496 OR2X1_LOC_151/A OR2X1_LOC_355/a_8_216# 0.02fF
C43497 AND2X1_LOC_355/a_8_24# OR2X1_LOC_331/Y 0.05fF
C43498 OR2X1_LOC_118/Y OR2X1_LOC_13/B 0.03fF
C43499 OR2X1_LOC_447/Y OR2X1_LOC_783/A 0.15fF
C43500 OR2X1_LOC_89/A AND2X1_LOC_779/Y 0.01fF
C43501 OR2X1_LOC_814/A OR2X1_LOC_227/Y 0.00fF
C43502 AND2X1_LOC_227/Y OR2X1_LOC_72/a_8_216# 0.03fF
C43503 AND2X1_LOC_738/B OR2X1_LOC_680/a_36_216# 0.01fF
C43504 AND2X1_LOC_564/B OR2X1_LOC_56/A 0.13fF
C43505 OR2X1_LOC_472/a_8_216# OR2X1_LOC_598/A 0.01fF
C43506 OR2X1_LOC_814/A D_INPUT_1 0.07fF
C43507 OR2X1_LOC_121/Y OR2X1_LOC_6/B 0.01fF
C43508 OR2X1_LOC_514/a_8_216# OR2X1_LOC_515/A -0.00fF
C43509 OR2X1_LOC_53/Y OR2X1_LOC_59/Y 0.05fF
C43510 AND2X1_LOC_303/B OR2X1_LOC_437/A 0.08fF
C43511 OR2X1_LOC_620/Y OR2X1_LOC_703/Y 0.01fF
C43512 OR2X1_LOC_133/a_8_216# OR2X1_LOC_604/A 0.06fF
C43513 OR2X1_LOC_676/Y OR2X1_LOC_138/A 0.01fF
C43514 OR2X1_LOC_185/A OR2X1_LOC_539/B 0.00fF
C43515 AND2X1_LOC_363/A OR2X1_LOC_384/Y 0.00fF
C43516 AND2X1_LOC_810/A VDD 0.50fF
C43517 OR2X1_LOC_22/Y OR2X1_LOC_41/a_8_216# 0.02fF
C43518 OR2X1_LOC_494/A OR2X1_LOC_91/A 0.08fF
C43519 AND2X1_LOC_22/Y OR2X1_LOC_78/A 0.14fF
C43520 OR2X1_LOC_375/A OR2X1_LOC_217/A 0.00fF
C43521 AND2X1_LOC_64/Y OR2X1_LOC_656/Y 0.05fF
C43522 AND2X1_LOC_866/A GATE_662 0.03fF
C43523 AND2X1_LOC_657/Y AND2X1_LOC_727/B 0.01fF
C43524 AND2X1_LOC_43/B OR2X1_LOC_593/B 0.03fF
C43525 OR2X1_LOC_40/Y AND2X1_LOC_477/Y 0.09fF
C43526 OR2X1_LOC_112/a_8_216# OR2X1_LOC_66/A 0.01fF
C43527 OR2X1_LOC_178/a_8_216# OR2X1_LOC_158/A 0.00fF
C43528 AND2X1_LOC_469/B AND2X1_LOC_727/B 0.03fF
C43529 AND2X1_LOC_810/a_8_24# AND2X1_LOC_810/Y 0.01fF
C43530 AND2X1_LOC_91/B AND2X1_LOC_421/a_8_24# 0.03fF
C43531 OR2X1_LOC_318/a_8_216# AND2X1_LOC_92/Y 0.04fF
C43532 OR2X1_LOC_696/A OR2X1_LOC_823/a_36_216# 0.00fF
C43533 AND2X1_LOC_401/a_8_24# OR2X1_LOC_415/Y 0.24fF
C43534 AND2X1_LOC_253/a_8_24# OR2X1_LOC_563/A 0.03fF
C43535 OR2X1_LOC_307/A OR2X1_LOC_66/A 0.22fF
C43536 OR2X1_LOC_48/B OR2X1_LOC_171/Y 0.03fF
C43537 OR2X1_LOC_276/B AND2X1_LOC_271/a_8_24# 0.02fF
C43538 OR2X1_LOC_6/A OR2X1_LOC_268/Y 0.00fF
C43539 OR2X1_LOC_561/Y OR2X1_LOC_843/B 0.01fF
C43540 AND2X1_LOC_454/A AND2X1_LOC_449/a_8_24# 0.02fF
C43541 OR2X1_LOC_575/A OR2X1_LOC_554/a_36_216# 0.01fF
C43542 OR2X1_LOC_756/B OR2X1_LOC_756/a_8_216# 0.09fF
C43543 OR2X1_LOC_858/A OR2X1_LOC_151/A 0.10fF
C43544 OR2X1_LOC_115/a_8_216# OR2X1_LOC_115/B 0.05fF
C43545 OR2X1_LOC_18/Y OR2X1_LOC_171/Y 0.52fF
C43546 OR2X1_LOC_186/Y AND2X1_LOC_312/a_8_24# 0.07fF
C43547 VDD AND2X1_LOC_860/A 0.58fF
C43548 AND2X1_LOC_711/A OR2X1_LOC_600/A 0.03fF
C43549 OR2X1_LOC_621/A OR2X1_LOC_78/A 0.19fF
C43550 OR2X1_LOC_604/A OR2X1_LOC_684/a_36_216# 0.00fF
C43551 AND2X1_LOC_40/Y AND2X1_LOC_44/Y 2.93fF
C43552 OR2X1_LOC_185/Y OR2X1_LOC_130/a_8_216# 0.02fF
C43553 OR2X1_LOC_190/A AND2X1_LOC_18/Y 0.03fF
C43554 AND2X1_LOC_47/Y OR2X1_LOC_318/B 0.03fF
C43555 OR2X1_LOC_604/A AND2X1_LOC_705/a_36_24# 0.00fF
C43556 AND2X1_LOC_539/Y OR2X1_LOC_619/Y 0.05fF
C43557 OR2X1_LOC_36/Y AND2X1_LOC_204/a_36_24# 0.00fF
C43558 AND2X1_LOC_539/Y AND2X1_LOC_356/a_8_24# 0.01fF
C43559 AND2X1_LOC_508/B OR2X1_LOC_51/Y 0.59fF
C43560 AND2X1_LOC_724/Y OR2X1_LOC_600/Y 0.02fF
C43561 OR2X1_LOC_40/Y OR2X1_LOC_329/B 0.46fF
C43562 OR2X1_LOC_287/B AND2X1_LOC_36/Y 0.02fF
C43563 OR2X1_LOC_496/a_8_216# AND2X1_LOC_658/A 0.03fF
C43564 AND2X1_LOC_386/a_8_24# AND2X1_LOC_36/Y 0.01fF
C43565 OR2X1_LOC_2/Y INPUT_7 0.07fF
C43566 AND2X1_LOC_649/a_8_24# AND2X1_LOC_786/Y 0.03fF
C43567 OR2X1_LOC_154/A OR2X1_LOC_120/a_8_216# 0.20fF
C43568 OR2X1_LOC_612/a_8_216# OR2X1_LOC_612/Y -0.00fF
C43569 AND2X1_LOC_855/a_8_24# OR2X1_LOC_13/B 0.02fF
C43570 OR2X1_LOC_51/Y AND2X1_LOC_508/a_8_24# 0.14fF
C43571 AND2X1_LOC_483/Y AND2X1_LOC_620/Y 0.01fF
C43572 AND2X1_LOC_266/a_36_24# OR2X1_LOC_595/A 0.00fF
C43573 OR2X1_LOC_600/A AND2X1_LOC_471/Y 0.02fF
C43574 OR2X1_LOC_130/A AND2X1_LOC_226/a_36_24# 0.01fF
C43575 OR2X1_LOC_4/a_8_216# OR2X1_LOC_80/A -0.03fF
C43576 OR2X1_LOC_527/a_8_216# OR2X1_LOC_164/Y 0.01fF
C43577 OR2X1_LOC_553/A OR2X1_LOC_121/A 0.01fF
C43578 OR2X1_LOC_31/Y OR2X1_LOC_172/Y 0.43fF
C43579 OR2X1_LOC_785/a_8_216# OR2X1_LOC_795/B -0.00fF
C43580 OR2X1_LOC_710/B AND2X1_LOC_144/a_8_24# 0.21fF
C43581 OR2X1_LOC_604/A OR2X1_LOC_292/Y 0.04fF
C43582 INPUT_1 OR2X1_LOC_71/A 0.07fF
C43583 OR2X1_LOC_333/B OR2X1_LOC_333/A 0.01fF
C43584 AND2X1_LOC_92/a_8_24# OR2X1_LOC_375/A 0.01fF
C43585 OR2X1_LOC_770/a_8_216# OR2X1_LOC_80/A 0.03fF
C43586 VDD OR2X1_LOC_459/A 0.21fF
C43587 OR2X1_LOC_657/a_8_216# OR2X1_LOC_267/Y 0.01fF
C43588 OR2X1_LOC_45/B AND2X1_LOC_655/A 0.10fF
C43589 OR2X1_LOC_26/Y AND2X1_LOC_772/Y 0.10fF
C43590 AND2X1_LOC_658/A AND2X1_LOC_444/a_36_24# 0.01fF
C43591 AND2X1_LOC_191/B AND2X1_LOC_474/A 0.03fF
C43592 AND2X1_LOC_570/Y AND2X1_LOC_506/a_8_24# 0.00fF
C43593 AND2X1_LOC_647/Y OR2X1_LOC_67/Y 0.80fF
C43594 AND2X1_LOC_812/a_8_24# OR2X1_LOC_152/A 0.01fF
C43595 OR2X1_LOC_87/Y AND2X1_LOC_44/Y 0.04fF
C43596 OR2X1_LOC_391/B OR2X1_LOC_774/a_8_216# 0.48fF
C43597 AND2X1_LOC_357/B AND2X1_LOC_357/a_8_24# 0.04fF
C43598 OR2X1_LOC_833/B OR2X1_LOC_719/B 0.02fF
C43599 AND2X1_LOC_794/A AND2X1_LOC_477/Y 0.02fF
C43600 OR2X1_LOC_369/a_8_216# AND2X1_LOC_716/Y 0.03fF
C43601 AND2X1_LOC_391/Y AND2X1_LOC_392/a_8_24# 0.01fF
C43602 OR2X1_LOC_348/a_8_216# OR2X1_LOC_791/B 0.01fF
C43603 AND2X1_LOC_365/a_8_24# OR2X1_LOC_744/A 0.04fF
C43604 OR2X1_LOC_175/B AND2X1_LOC_110/Y 0.83fF
C43605 OR2X1_LOC_832/a_36_216# OR2X1_LOC_502/A 0.00fF
C43606 OR2X1_LOC_106/a_8_216# AND2X1_LOC_99/A 0.01fF
C43607 AND2X1_LOC_112/a_8_24# OR2X1_LOC_92/Y 0.03fF
C43608 OR2X1_LOC_160/A AND2X1_LOC_65/A 0.02fF
C43609 OR2X1_LOC_89/A AND2X1_LOC_772/Y 0.62fF
C43610 OR2X1_LOC_720/a_8_216# OR2X1_LOC_720/Y -0.00fF
C43611 AND2X1_LOC_347/Y OR2X1_LOC_56/A 0.00fF
C43612 AND2X1_LOC_710/Y AND2X1_LOC_347/Y 0.17fF
C43613 VDD AND2X1_LOC_155/a_8_24# -0.00fF
C43614 AND2X1_LOC_319/A OR2X1_LOC_12/Y 0.01fF
C43615 AND2X1_LOC_857/Y OR2X1_LOC_56/A 0.04fF
C43616 OR2X1_LOC_357/a_8_216# OR2X1_LOC_87/A 0.01fF
C43617 OR2X1_LOC_594/Y AND2X1_LOC_436/Y 0.01fF
C43618 OR2X1_LOC_39/Y INPUT_0 0.16fF
C43619 OR2X1_LOC_112/a_36_216# OR2X1_LOC_539/Y 0.00fF
C43620 AND2X1_LOC_22/Y OR2X1_LOC_155/A 0.05fF
C43621 OR2X1_LOC_696/A AND2X1_LOC_663/B 0.03fF
C43622 OR2X1_LOC_207/B OR2X1_LOC_200/a_8_216# 0.01fF
C43623 AND2X1_LOC_364/a_8_24# OR2X1_LOC_43/A 0.09fF
C43624 VDD OR2X1_LOC_668/a_8_216# 0.21fF
C43625 OR2X1_LOC_160/B OR2X1_LOC_784/Y 0.11fF
C43626 OR2X1_LOC_335/a_8_216# OR2X1_LOC_479/Y 0.04fF
C43627 OR2X1_LOC_207/B OR2X1_LOC_269/B 0.07fF
C43628 OR2X1_LOC_709/A OR2X1_LOC_793/A 0.18fF
C43629 AND2X1_LOC_12/Y OR2X1_LOC_6/B 0.22fF
C43630 OR2X1_LOC_560/a_8_216# OR2X1_LOC_66/A 0.01fF
C43631 OR2X1_LOC_489/A OR2X1_LOC_269/B 0.02fF
C43632 OR2X1_LOC_154/A OR2X1_LOC_596/A 0.07fF
C43633 OR2X1_LOC_45/B OR2X1_LOC_609/A 0.08fF
C43634 AND2X1_LOC_41/a_8_24# AND2X1_LOC_43/B -0.04fF
C43635 AND2X1_LOC_571/a_8_24# AND2X1_LOC_489/Y 0.02fF
C43636 VDD AND2X1_LOC_400/a_8_24# 0.00fF
C43637 OR2X1_LOC_608/a_8_216# OR2X1_LOC_78/B 0.03fF
C43638 AND2X1_LOC_648/B AND2X1_LOC_592/a_8_24# -0.00fF
C43639 AND2X1_LOC_431/a_8_24# OR2X1_LOC_539/B 0.18fF
C43640 OR2X1_LOC_6/B AND2X1_LOC_838/Y 0.01fF
C43641 OR2X1_LOC_176/Y AND2X1_LOC_566/Y 0.17fF
C43642 OR2X1_LOC_756/Y AND2X1_LOC_757/a_8_24# 0.01fF
C43643 OR2X1_LOC_287/B AND2X1_LOC_488/a_8_24# 0.01fF
C43644 OR2X1_LOC_53/Y OR2X1_LOC_70/Y 0.00fF
C43645 AND2X1_LOC_51/Y OR2X1_LOC_334/a_8_216# 0.01fF
C43646 AND2X1_LOC_22/Y OR2X1_LOC_605/A 0.04fF
C43647 AND2X1_LOC_81/B OR2X1_LOC_641/A 0.03fF
C43648 OR2X1_LOC_459/A OR2X1_LOC_689/A 0.09fF
C43649 OR2X1_LOC_97/A AND2X1_LOC_42/B 0.00fF
C43650 OR2X1_LOC_589/A OR2X1_LOC_43/A 1.11fF
C43651 OR2X1_LOC_447/Y OR2X1_LOC_308/Y 0.02fF
C43652 OR2X1_LOC_18/Y AND2X1_LOC_629/a_8_24# 0.03fF
C43653 AND2X1_LOC_64/Y OR2X1_LOC_206/A 0.01fF
C43654 OR2X1_LOC_744/A AND2X1_LOC_76/Y 0.03fF
C43655 OR2X1_LOC_326/B OR2X1_LOC_538/A 0.00fF
C43656 AND2X1_LOC_858/B OR2X1_LOC_427/A 0.08fF
C43657 OR2X1_LOC_630/a_8_216# OR2X1_LOC_78/A 0.01fF
C43658 OR2X1_LOC_91/A OR2X1_LOC_427/A 0.17fF
C43659 AND2X1_LOC_394/a_8_24# OR2X1_LOC_66/A 0.01fF
C43660 OR2X1_LOC_703/B VDD 0.24fF
C43661 OR2X1_LOC_680/A AND2X1_LOC_508/B 0.03fF
C43662 OR2X1_LOC_254/B OR2X1_LOC_542/B 0.03fF
C43663 OR2X1_LOC_279/Y AND2X1_LOC_244/A 0.05fF
C43664 AND2X1_LOC_652/a_36_24# AND2X1_LOC_436/Y 0.00fF
C43665 AND2X1_LOC_566/Y AND2X1_LOC_212/Y 0.34fF
C43666 OR2X1_LOC_476/B OR2X1_LOC_390/a_8_216# 0.01fF
C43667 AND2X1_LOC_59/Y OR2X1_LOC_650/a_8_216# 0.01fF
C43668 OR2X1_LOC_185/A OR2X1_LOC_78/B 0.36fF
C43669 OR2X1_LOC_664/a_8_216# OR2X1_LOC_78/A 0.03fF
C43670 OR2X1_LOC_666/a_8_216# OR2X1_LOC_283/a_8_216# 0.47fF
C43671 OR2X1_LOC_70/Y AND2X1_LOC_802/Y 0.03fF
C43672 OR2X1_LOC_782/B VDD 0.00fF
C43673 VDD AND2X1_LOC_287/Y 0.02fF
C43674 OR2X1_LOC_517/A AND2X1_LOC_845/a_36_24# 0.00fF
C43675 OR2X1_LOC_137/a_8_216# AND2X1_LOC_95/Y 0.09fF
C43676 OR2X1_LOC_269/B OR2X1_LOC_772/A 0.02fF
C43677 VDD OR2X1_LOC_87/A 1.71fF
C43678 OR2X1_LOC_22/Y AND2X1_LOC_227/a_8_24# 0.01fF
C43679 AND2X1_LOC_657/A AND2X1_LOC_562/Y 0.06fF
C43680 AND2X1_LOC_140/a_8_24# OR2X1_LOC_12/Y 0.01fF
C43681 OR2X1_LOC_744/A OR2X1_LOC_67/A 0.03fF
C43682 AND2X1_LOC_170/Y AND2X1_LOC_568/B 0.02fF
C43683 OR2X1_LOC_426/A OR2X1_LOC_2/Y 0.18fF
C43684 OR2X1_LOC_9/Y OR2X1_LOC_73/a_8_216# 0.02fF
C43685 AND2X1_LOC_390/B OR2X1_LOC_13/a_8_216# 0.03fF
C43686 OR2X1_LOC_235/B OR2X1_LOC_38/a_36_216# 0.01fF
C43687 OR2X1_LOC_275/A OR2X1_LOC_595/A 0.10fF
C43688 AND2X1_LOC_361/a_8_24# AND2X1_LOC_276/Y 0.00fF
C43689 OR2X1_LOC_251/Y AND2X1_LOC_860/A 0.15fF
C43690 OR2X1_LOC_242/a_36_216# OR2X1_LOC_375/A 0.00fF
C43691 AND2X1_LOC_561/B OR2X1_LOC_44/Y 0.03fF
C43692 OR2X1_LOC_405/A OR2X1_LOC_216/A 0.02fF
C43693 OR2X1_LOC_662/a_8_216# OR2X1_LOC_130/A 0.05fF
C43694 AND2X1_LOC_737/a_8_24# AND2X1_LOC_550/A 0.03fF
C43695 OR2X1_LOC_508/a_8_216# AND2X1_LOC_51/Y 0.00fF
C43696 AND2X1_LOC_693/a_8_24# OR2X1_LOC_375/A 0.09fF
C43697 OR2X1_LOC_686/B AND2X1_LOC_683/a_8_24# 0.03fF
C43698 AND2X1_LOC_725/a_36_24# OR2X1_LOC_7/A 0.01fF
C43699 OR2X1_LOC_19/B OR2X1_LOC_548/B 0.01fF
C43700 OR2X1_LOC_118/Y AND2X1_LOC_266/a_8_24# 0.01fF
C43701 OR2X1_LOC_6/B AND2X1_LOC_496/a_8_24# 0.02fF
C43702 OR2X1_LOC_166/Y OR2X1_LOC_43/A 0.49fF
C43703 OR2X1_LOC_438/Y AND2X1_LOC_624/A 0.03fF
C43704 OR2X1_LOC_311/Y AND2X1_LOC_810/B 0.01fF
C43705 OR2X1_LOC_631/B OR2X1_LOC_632/Y 0.01fF
C43706 OR2X1_LOC_43/A OR2X1_LOC_297/A 0.01fF
C43707 OR2X1_LOC_502/A OR2X1_LOC_539/Y 0.03fF
C43708 OR2X1_LOC_526/Y OR2X1_LOC_680/Y 0.38fF
C43709 AND2X1_LOC_729/Y OR2X1_LOC_144/Y 0.31fF
C43710 OR2X1_LOC_235/B AND2X1_LOC_399/a_8_24# 0.04fF
C43711 OR2X1_LOC_744/A OR2X1_LOC_52/B 0.13fF
C43712 OR2X1_LOC_91/Y OR2X1_LOC_165/Y 0.05fF
C43713 AND2X1_LOC_2/Y AND2X1_LOC_3/Y 0.01fF
C43714 AND2X1_LOC_363/A OR2X1_LOC_91/A 0.16fF
C43715 OR2X1_LOC_326/B AND2X1_LOC_12/Y 0.00fF
C43716 OR2X1_LOC_604/A OR2X1_LOC_430/a_36_216# 0.02fF
C43717 AND2X1_LOC_712/B OR2X1_LOC_421/Y 0.10fF
C43718 AND2X1_LOC_197/Y OR2X1_LOC_44/Y 0.01fF
C43719 OR2X1_LOC_427/A AND2X1_LOC_573/A 0.14fF
C43720 AND2X1_LOC_593/a_8_24# OR2X1_LOC_64/Y 0.02fF
C43721 OR2X1_LOC_296/a_8_216# OR2X1_LOC_78/A 0.01fF
C43722 OR2X1_LOC_329/B OR2X1_LOC_7/A 0.46fF
C43723 OR2X1_LOC_823/a_8_216# OR2X1_LOC_823/Y -0.00fF
C43724 OR2X1_LOC_859/a_8_216# OR2X1_LOC_269/B 0.00fF
C43725 OR2X1_LOC_35/B OR2X1_LOC_66/A 0.25fF
C43726 INPUT_4 OR2X1_LOC_2/Y 1.11fF
C43727 OR2X1_LOC_833/a_8_216# OR2X1_LOC_203/Y 0.04fF
C43728 AND2X1_LOC_489/Y OR2X1_LOC_744/A 0.09fF
C43729 AND2X1_LOC_784/A AND2X1_LOC_477/a_36_24# 0.01fF
C43730 OR2X1_LOC_51/Y AND2X1_LOC_639/a_36_24# 0.00fF
C43731 OR2X1_LOC_401/Y OR2X1_LOC_78/Y 0.02fF
C43732 AND2X1_LOC_541/Y OR2X1_LOC_22/Y 0.02fF
C43733 OR2X1_LOC_95/Y AND2X1_LOC_786/Y 0.07fF
C43734 OR2X1_LOC_43/A AND2X1_LOC_654/B 0.21fF
C43735 OR2X1_LOC_604/a_8_216# OR2X1_LOC_12/Y 0.01fF
C43736 AND2X1_LOC_621/Y AND2X1_LOC_624/A 20.56fF
C43737 OR2X1_LOC_185/A OR2X1_LOC_375/A 0.28fF
C43738 OR2X1_LOC_95/Y OR2X1_LOC_323/a_8_216# 0.01fF
C43739 OR2X1_LOC_262/Y AND2X1_LOC_266/a_8_24# 0.03fF
C43740 OR2X1_LOC_541/A AND2X1_LOC_42/B 0.02fF
C43741 OR2X1_LOC_154/A OR2X1_LOC_732/a_8_216# 0.03fF
C43742 OR2X1_LOC_368/A AND2X1_LOC_786/Y 0.06fF
C43743 AND2X1_LOC_512/Y AND2X1_LOC_337/B 0.01fF
C43744 OR2X1_LOC_185/Y OR2X1_LOC_194/B 0.01fF
C43745 AND2X1_LOC_160/a_8_24# OR2X1_LOC_743/A 0.09fF
C43746 AND2X1_LOC_56/B OR2X1_LOC_833/B 0.01fF
C43747 OR2X1_LOC_520/Y OR2X1_LOC_660/B 0.04fF
C43748 OR2X1_LOC_653/Y AND2X1_LOC_8/Y 0.00fF
C43749 OR2X1_LOC_854/a_36_216# OR2X1_LOC_155/A 0.01fF
C43750 AND2X1_LOC_76/Y OR2X1_LOC_74/a_8_216# 0.01fF
C43751 AND2X1_LOC_172/a_8_24# AND2X1_LOC_48/A 0.01fF
C43752 OR2X1_LOC_80/Y OR2X1_LOC_69/A 0.02fF
C43753 OR2X1_LOC_633/Y OR2X1_LOC_97/B 0.00fF
C43754 OR2X1_LOC_669/Y OR2X1_LOC_427/A 0.07fF
C43755 OR2X1_LOC_413/Y OR2X1_LOC_44/Y 0.03fF
C43756 OR2X1_LOC_335/B OR2X1_LOC_370/a_8_216# 0.47fF
C43757 OR2X1_LOC_18/Y AND2X1_LOC_806/A 0.04fF
C43758 AND2X1_LOC_105/a_8_24# OR2X1_LOC_278/Y 0.01fF
C43759 VDD OR2X1_LOC_706/B 0.00fF
C43760 OR2X1_LOC_468/A OR2X1_LOC_168/A 0.02fF
C43761 AND2X1_LOC_784/Y AND2X1_LOC_675/A 0.01fF
C43762 AND2X1_LOC_486/Y OR2X1_LOC_74/A 0.07fF
C43763 OR2X1_LOC_256/Y OR2X1_LOC_481/A 0.01fF
C43764 OR2X1_LOC_848/A OR2X1_LOC_848/a_8_216# 0.06fF
C43765 OR2X1_LOC_201/A OR2X1_LOC_215/A 0.95fF
C43766 OR2X1_LOC_45/B OR2X1_LOC_599/Y 3.79fF
C43767 AND2X1_LOC_365/A OR2X1_LOC_43/A 0.02fF
C43768 OR2X1_LOC_107/a_8_216# OR2X1_LOC_22/Y 0.05fF
C43769 OR2X1_LOC_114/B AND2X1_LOC_47/Y 3.29fF
C43770 OR2X1_LOC_696/a_8_216# OR2X1_LOC_48/B 0.02fF
C43771 OR2X1_LOC_91/A AND2X1_LOC_687/B 0.07fF
C43772 INPUT_0 OR2X1_LOC_46/A 1.42fF
C43773 OR2X1_LOC_235/B AND2X1_LOC_671/a_8_24# -0.01fF
C43774 AND2X1_LOC_721/A OR2X1_LOC_12/Y 0.03fF
C43775 OR2X1_LOC_74/A AND2X1_LOC_811/B 0.08fF
C43776 OR2X1_LOC_756/B OR2X1_LOC_34/B 0.01fF
C43777 OR2X1_LOC_510/Y OR2X1_LOC_217/a_8_216# 0.01fF
C43778 OR2X1_LOC_53/Y OR2X1_LOC_70/A 0.01fF
C43779 INPUT_1 OR2X1_LOC_59/Y 0.09fF
C43780 OR2X1_LOC_9/Y OR2X1_LOC_619/a_8_216# 0.01fF
C43781 VDD OR2X1_LOC_607/Y 0.12fF
C43782 AND2X1_LOC_852/Y OR2X1_LOC_69/a_8_216# 0.06fF
C43783 OR2X1_LOC_40/Y GATE_662 0.61fF
C43784 AND2X1_LOC_370/a_8_24# AND2X1_LOC_222/Y -0.01fF
C43785 OR2X1_LOC_18/Y AND2X1_LOC_276/Y 0.16fF
C43786 OR2X1_LOC_40/Y GATE_811 0.03fF
C43787 AND2X1_LOC_431/a_8_24# OR2X1_LOC_78/B 0.03fF
C43788 OR2X1_LOC_532/B OR2X1_LOC_778/B 0.01fF
C43789 AND2X1_LOC_729/Y OR2X1_LOC_420/Y 0.02fF
C43790 OR2X1_LOC_702/A OR2X1_LOC_377/A 0.64fF
C43791 OR2X1_LOC_476/B AND2X1_LOC_58/a_8_24# 0.03fF
C43792 OR2X1_LOC_185/A OR2X1_LOC_605/B 0.04fF
C43793 OR2X1_LOC_122/a_36_216# AND2X1_LOC_845/Y 0.01fF
C43794 OR2X1_LOC_251/Y AND2X1_LOC_287/Y 0.01fF
C43795 OR2X1_LOC_493/A AND2X1_LOC_67/Y 0.18fF
C43796 AND2X1_LOC_840/B OR2X1_LOC_52/B 0.07fF
C43797 OR2X1_LOC_36/Y AND2X1_LOC_688/a_8_24# 0.02fF
C43798 INPUT_3 OR2X1_LOC_8/a_8_216# 0.03fF
C43799 OR2X1_LOC_121/Y OR2X1_LOC_598/A 0.03fF
C43800 AND2X1_LOC_578/A AND2X1_LOC_807/Y 0.07fF
C43801 OR2X1_LOC_678/Y AND2X1_LOC_53/Y 0.02fF
C43802 OR2X1_LOC_624/B OR2X1_LOC_659/a_8_216# 0.01fF
C43803 OR2X1_LOC_486/Y OR2X1_LOC_551/B 0.07fF
C43804 OR2X1_LOC_290/Y AND2X1_LOC_634/Y 0.15fF
C43805 OR2X1_LOC_74/a_8_216# OR2X1_LOC_52/B 0.03fF
C43806 AND2X1_LOC_660/Y OR2X1_LOC_65/B 0.14fF
C43807 AND2X1_LOC_63/a_8_24# AND2X1_LOC_42/B 0.01fF
C43808 OR2X1_LOC_494/Y OR2X1_LOC_47/Y 0.01fF
C43809 AND2X1_LOC_576/Y AND2X1_LOC_717/B 0.07fF
C43810 OR2X1_LOC_538/A AND2X1_LOC_47/Y 0.03fF
C43811 D_INPUT_7 AND2X1_LOC_30/a_8_24# 0.10fF
C43812 AND2X1_LOC_304/a_8_24# AND2X1_LOC_53/Y 0.09fF
C43813 AND2X1_LOC_363/Y OR2X1_LOC_47/Y 0.02fF
C43814 AND2X1_LOC_624/B AND2X1_LOC_254/a_8_24# 0.01fF
C43815 OR2X1_LOC_429/Y OR2X1_LOC_25/a_36_216# 0.01fF
C43816 AND2X1_LOC_580/B OR2X1_LOC_89/A 0.06fF
C43817 AND2X1_LOC_3/Y OR2X1_LOC_269/B 3.84fF
C43818 OR2X1_LOC_318/A AND2X1_LOC_31/Y 0.01fF
C43819 OR2X1_LOC_675/A OR2X1_LOC_805/A 0.03fF
C43820 AND2X1_LOC_345/Y OR2X1_LOC_6/A 0.08fF
C43821 OR2X1_LOC_375/A OR2X1_LOC_713/a_8_216# 0.01fF
C43822 OR2X1_LOC_244/Y D_INPUT_1 0.03fF
C43823 AND2X1_LOC_18/Y OR2X1_LOC_241/B 0.70fF
C43824 AND2X1_LOC_624/B OR2X1_LOC_626/Y 0.07fF
C43825 OR2X1_LOC_160/B AND2X1_LOC_72/B 0.03fF
C43826 OR2X1_LOC_54/Y OR2X1_LOC_38/a_8_216# 0.04fF
C43827 AND2X1_LOC_119/a_8_24# OR2X1_LOC_375/A 0.06fF
C43828 OR2X1_LOC_12/Y AND2X1_LOC_217/a_8_24# 0.01fF
C43829 OR2X1_LOC_476/B AND2X1_LOC_824/B 0.53fF
C43830 AND2X1_LOC_95/Y OR2X1_LOC_814/A 0.17fF
C43831 OR2X1_LOC_841/A OR2X1_LOC_804/A 0.01fF
C43832 OR2X1_LOC_151/A OR2X1_LOC_736/a_36_216# 0.00fF
C43833 AND2X1_LOC_621/a_8_24# AND2X1_LOC_621/Y 0.00fF
C43834 OR2X1_LOC_151/A AND2X1_LOC_31/Y 0.36fF
C43835 AND2X1_LOC_342/Y OR2X1_LOC_19/B 0.02fF
C43836 OR2X1_LOC_470/a_8_216# AND2X1_LOC_51/Y 0.07fF
C43837 OR2X1_LOC_460/a_8_216# AND2X1_LOC_3/Y 0.01fF
C43838 OR2X1_LOC_516/Y AND2X1_LOC_785/A 0.15fF
C43839 OR2X1_LOC_22/Y OR2X1_LOC_316/Y 0.03fF
C43840 OR2X1_LOC_243/A OR2X1_LOC_62/B 0.00fF
C43841 AND2X1_LOC_356/B AND2X1_LOC_390/B 0.01fF
C43842 AND2X1_LOC_12/Y OR2X1_LOC_68/Y 0.01fF
C43843 OR2X1_LOC_154/A AND2X1_LOC_79/a_8_24# 0.07fF
C43844 AND2X1_LOC_303/A AND2X1_LOC_537/Y 0.02fF
C43845 AND2X1_LOC_76/Y OR2X1_LOC_31/Y 0.10fF
C43846 AND2X1_LOC_561/a_8_24# AND2X1_LOC_571/B 0.00fF
C43847 OR2X1_LOC_175/Y OR2X1_LOC_174/Y 0.00fF
C43848 OR2X1_LOC_444/B OR2X1_LOC_87/A 0.03fF
C43849 INPUT_0 OR2X1_LOC_41/Y 0.04fF
C43850 VDD AND2X1_LOC_562/Y 0.72fF
C43851 OR2X1_LOC_744/A AND2X1_LOC_216/A 0.02fF
C43852 OR2X1_LOC_64/Y OR2X1_LOC_106/A 0.01fF
C43853 AND2X1_LOC_3/Y OR2X1_LOC_215/A 0.03fF
C43854 OR2X1_LOC_161/B OR2X1_LOC_707/a_8_216# 0.01fF
C43855 AND2X1_LOC_170/a_8_24# AND2X1_LOC_170/B -0.00fF
C43856 OR2X1_LOC_665/a_8_216# OR2X1_LOC_665/Y 0.00fF
C43857 OR2X1_LOC_36/Y OR2X1_LOC_62/B 0.02fF
C43858 AND2X1_LOC_12/Y AND2X1_LOC_47/Y 0.19fF
C43859 OR2X1_LOC_147/B OR2X1_LOC_284/B 0.08fF
C43860 OR2X1_LOC_481/A OR2X1_LOC_258/Y 0.02fF
C43861 OR2X1_LOC_690/A OR2X1_LOC_46/A 0.39fF
C43862 OR2X1_LOC_358/a_36_216# OR2X1_LOC_532/B 0.00fF
C43863 AND2X1_LOC_162/a_8_24# OR2X1_LOC_163/Y 0.01fF
C43864 OR2X1_LOC_532/B OR2X1_LOC_720/A 0.01fF
C43865 OR2X1_LOC_503/A AND2X1_LOC_227/Y 0.00fF
C43866 OR2X1_LOC_168/A OR2X1_LOC_449/B 0.04fF
C43867 INPUT_1 OR2X1_LOC_820/B 0.42fF
C43868 AND2X1_LOC_41/A OR2X1_LOC_358/A 0.07fF
C43869 OR2X1_LOC_167/Y AND2X1_LOC_661/A 0.02fF
C43870 OR2X1_LOC_485/A AND2X1_LOC_537/Y 0.02fF
C43871 AND2X1_LOC_580/A AND2X1_LOC_866/A 0.03fF
C43872 OR2X1_LOC_217/A OR2X1_LOC_549/A 0.01fF
C43873 AND2X1_LOC_785/A OR2X1_LOC_373/a_8_216# 0.47fF
C43874 OR2X1_LOC_532/B OR2X1_LOC_722/a_8_216# 0.00fF
C43875 AND2X1_LOC_394/a_8_24# OR2X1_LOC_84/A 0.03fF
C43876 OR2X1_LOC_31/Y AND2X1_LOC_374/Y 0.01fF
C43877 AND2X1_LOC_560/B AND2X1_LOC_227/Y 0.12fF
C43878 OR2X1_LOC_405/A OR2X1_LOC_205/Y 0.03fF
C43879 OR2X1_LOC_454/a_8_216# OR2X1_LOC_449/B 0.01fF
C43880 AND2X1_LOC_390/B OR2X1_LOC_22/Y 0.15fF
C43881 OR2X1_LOC_496/Y AND2X1_LOC_675/A 0.02fF
C43882 OR2X1_LOC_267/Y OR2X1_LOC_140/B 0.21fF
C43883 OR2X1_LOC_31/Y OR2X1_LOC_52/B 0.25fF
C43884 OR2X1_LOC_709/B OR2X1_LOC_308/Y 0.04fF
C43885 AND2X1_LOC_477/A OR2X1_LOC_417/a_8_216# 0.01fF
C43886 AND2X1_LOC_642/Y AND2X1_LOC_222/Y 0.88fF
C43887 OR2X1_LOC_70/Y INPUT_1 0.03fF
C43888 OR2X1_LOC_710/A AND2X1_LOC_44/Y 0.01fF
C43889 D_INPUT_3 OR2X1_LOC_585/A 0.03fF
C43890 OR2X1_LOC_56/A OR2X1_LOC_437/A 0.48fF
C43891 OR2X1_LOC_651/B AND2X1_LOC_31/Y 0.06fF
C43892 OR2X1_LOC_64/Y OR2X1_LOC_46/A 0.05fF
C43893 AND2X1_LOC_47/Y AND2X1_LOC_79/Y 0.03fF
C43894 OR2X1_LOC_574/A OR2X1_LOC_276/A 0.08fF
C43895 OR2X1_LOC_431/Y OR2X1_LOC_22/Y 0.42fF
C43896 OR2X1_LOC_506/A OR2X1_LOC_318/B 0.02fF
C43897 AND2X1_LOC_12/Y OR2X1_LOC_598/A 0.22fF
C43898 OR2X1_LOC_19/B OR2X1_LOC_54/Y 0.05fF
C43899 OR2X1_LOC_596/Y OR2X1_LOC_214/B 0.04fF
C43900 OR2X1_LOC_270/Y OR2X1_LOC_269/B 0.01fF
C43901 AND2X1_LOC_15/a_8_24# AND2X1_LOC_51/Y 0.01fF
C43902 AND2X1_LOC_433/a_36_24# OR2X1_LOC_390/B 0.00fF
C43903 OR2X1_LOC_291/Y AND2X1_LOC_634/Y 0.02fF
C43904 AND2X1_LOC_578/A OR2X1_LOC_95/Y 0.34fF
C43905 VDD OR2X1_LOC_579/A 0.18fF
C43906 OR2X1_LOC_160/B AND2X1_LOC_36/Y 0.06fF
C43907 OR2X1_LOC_154/A OR2X1_LOC_374/Y 0.19fF
C43908 OR2X1_LOC_45/Y OR2X1_LOC_172/a_8_216# -0.03fF
C43909 AND2X1_LOC_64/Y OR2X1_LOC_185/a_8_216# 0.01fF
C43910 OR2X1_LOC_506/A OR2X1_LOC_854/A 0.03fF
C43911 OR2X1_LOC_529/Y OR2X1_LOC_224/Y 0.02fF
C43912 AND2X1_LOC_632/a_8_24# OR2X1_LOC_95/Y 0.03fF
C43913 OR2X1_LOC_74/A AND2X1_LOC_660/A 0.07fF
C43914 AND2X1_LOC_92/Y OR2X1_LOC_716/a_36_216# 0.01fF
C43915 OR2X1_LOC_269/B AND2X1_LOC_225/a_8_24# 0.01fF
C43916 OR2X1_LOC_114/Y OR2X1_LOC_66/Y 0.00fF
C43917 OR2X1_LOC_269/B OR2X1_LOC_194/a_8_216# 0.03fF
C43918 OR2X1_LOC_661/a_8_216# OR2X1_LOC_68/B 0.01fF
C43919 OR2X1_LOC_61/Y AND2X1_LOC_406/a_8_24# 0.06fF
C43920 AND2X1_LOC_227/Y OR2X1_LOC_64/Y 0.07fF
C43921 AND2X1_LOC_392/A OR2X1_LOC_696/A 0.07fF
C43922 AND2X1_LOC_631/Y OR2X1_LOC_615/Y 0.01fF
C43923 OR2X1_LOC_516/Y AND2X1_LOC_658/A 0.07fF
C43924 OR2X1_LOC_691/Y OR2X1_LOC_855/a_8_216# 0.03fF
C43925 OR2X1_LOC_417/A OR2X1_LOC_46/A 0.67fF
C43926 OR2X1_LOC_160/B OR2X1_LOC_333/a_8_216# 0.01fF
C43927 OR2X1_LOC_22/Y AND2X1_LOC_863/Y 0.07fF
C43928 OR2X1_LOC_687/Y AND2X1_LOC_430/B 0.00fF
C43929 OR2X1_LOC_620/a_8_216# AND2X1_LOC_44/Y 0.14fF
C43930 OR2X1_LOC_417/Y AND2X1_LOC_645/a_8_24# 0.03fF
C43931 AND2X1_LOC_131/a_36_24# OR2X1_LOC_115/B 0.00fF
C43932 OR2X1_LOC_462/B OR2X1_LOC_68/B 0.05fF
C43933 AND2X1_LOC_771/B AND2X1_LOC_769/Y 0.09fF
C43934 OR2X1_LOC_85/A AND2X1_LOC_203/a_8_24# 0.01fF
C43935 OR2X1_LOC_840/A OR2X1_LOC_723/B 1.25fF
C43936 OR2X1_LOC_691/Y OR2X1_LOC_729/a_8_216# 0.12fF
C43937 OR2X1_LOC_85/A AND2X1_LOC_206/Y 0.02fF
C43938 OR2X1_LOC_843/B OR2X1_LOC_343/a_8_216# 0.05fF
C43939 OR2X1_LOC_251/Y AND2X1_LOC_562/Y 0.01fF
C43940 AND2X1_LOC_555/Y AND2X1_LOC_191/B 0.03fF
C43941 OR2X1_LOC_375/A OR2X1_LOC_705/a_8_216# 0.01fF
C43942 OR2X1_LOC_188/Y AND2X1_LOC_18/Y 0.01fF
C43943 AND2X1_LOC_227/Y OR2X1_LOC_417/A 0.03fF
C43944 OR2X1_LOC_154/a_8_216# OR2X1_LOC_160/B 0.01fF
C43945 OR2X1_LOC_64/Y OR2X1_LOC_813/Y 0.52fF
C43946 OR2X1_LOC_538/A OR2X1_LOC_186/a_8_216# 0.01fF
C43947 AND2X1_LOC_14/a_8_24# INPUT_1 0.01fF
C43948 OR2X1_LOC_664/Y OR2X1_LOC_366/Y 0.08fF
C43949 OR2X1_LOC_339/a_36_216# AND2X1_LOC_7/B 0.02fF
C43950 OR2X1_LOC_502/A OR2X1_LOC_319/Y 0.07fF
C43951 OR2X1_LOC_421/A OR2X1_LOC_16/A 0.03fF
C43952 OR2X1_LOC_160/B AND2X1_LOC_488/a_8_24# 0.04fF
C43953 OR2X1_LOC_382/A OR2X1_LOC_382/a_8_216# 0.39fF
C43954 AND2X1_LOC_64/Y OR2X1_LOC_756/B 0.26fF
C43955 AND2X1_LOC_719/Y OR2X1_LOC_158/A 0.07fF
C43956 AND2X1_LOC_338/A OR2X1_LOC_600/A 0.08fF
C43957 OR2X1_LOC_263/a_8_216# OR2X1_LOC_67/Y 0.01fF
C43958 AND2X1_LOC_349/a_8_24# OR2X1_LOC_13/B 0.01fF
C43959 INPUT_3 AND2X1_LOC_36/Y 0.07fF
C43960 AND2X1_LOC_180/a_8_24# OR2X1_LOC_40/Y 0.02fF
C43961 OR2X1_LOC_471/Y OR2X1_LOC_545/a_8_216# 0.06fF
C43962 OR2X1_LOC_840/a_8_216# VDD 0.00fF
C43963 AND2X1_LOC_339/Y AND2X1_LOC_219/Y 0.03fF
C43964 OR2X1_LOC_137/a_8_216# AND2X1_LOC_22/Y 0.05fF
C43965 OR2X1_LOC_319/B OR2X1_LOC_703/a_8_216# 0.05fF
C43966 OR2X1_LOC_738/A OR2X1_LOC_731/B 0.04fF
C43967 OR2X1_LOC_696/A AND2X1_LOC_354/Y 0.03fF
C43968 OR2X1_LOC_604/A OR2X1_LOC_672/a_36_216# 0.01fF
C43969 OR2X1_LOC_553/A AND2X1_LOC_36/Y 0.07fF
C43970 AND2X1_LOC_264/a_36_24# OR2X1_LOC_13/B 0.00fF
C43971 OR2X1_LOC_93/Y OR2X1_LOC_96/Y 0.08fF
C43972 OR2X1_LOC_630/B OR2X1_LOC_161/B 0.02fF
C43973 AND2X1_LOC_456/B AND2X1_LOC_244/A 0.02fF
C43974 AND2X1_LOC_40/Y OR2X1_LOC_352/a_8_216# 0.01fF
C43975 AND2X1_LOC_22/Y AND2X1_LOC_71/a_36_24# 0.01fF
C43976 OR2X1_LOC_607/Y OR2X1_LOC_67/Y 0.03fF
C43977 OR2X1_LOC_532/B OR2X1_LOC_590/a_8_216# 0.18fF
C43978 OR2X1_LOC_287/B OR2X1_LOC_571/Y 0.00fF
C43979 OR2X1_LOC_22/Y OR2X1_LOC_153/a_8_216# 0.03fF
C43980 OR2X1_LOC_505/Y AND2X1_LOC_507/a_8_24# 0.01fF
C43981 AND2X1_LOC_605/Y OR2X1_LOC_12/Y 0.04fF
C43982 AND2X1_LOC_39/a_8_24# AND2X1_LOC_44/Y 0.03fF
C43983 OR2X1_LOC_756/B AND2X1_LOC_82/Y 0.01fF
C43984 AND2X1_LOC_217/Y OR2X1_LOC_132/a_8_216# 0.03fF
C43985 OR2X1_LOC_3/Y OR2X1_LOC_424/Y 0.00fF
C43986 AND2X1_LOC_654/Y OR2X1_LOC_321/a_36_216# 0.01fF
C43987 AND2X1_LOC_715/Y AND2X1_LOC_354/Y 0.01fF
C43988 AND2X1_LOC_749/a_36_24# AND2X1_LOC_44/Y 0.01fF
C43989 AND2X1_LOC_42/B OR2X1_LOC_141/a_8_216# 0.01fF
C43990 AND2X1_LOC_566/B AND2X1_LOC_364/Y 0.12fF
C43991 VDD OR2X1_LOC_801/a_8_216# 0.00fF
C43992 AND2X1_LOC_228/Y OR2X1_LOC_171/Y 0.28fF
C43993 AND2X1_LOC_447/Y AND2X1_LOC_454/a_8_24# 0.11fF
C43994 OR2X1_LOC_527/a_8_216# AND2X1_LOC_471/Y 0.49fF
C43995 OR2X1_LOC_160/B OR2X1_LOC_630/Y 0.07fF
C43996 AND2X1_LOC_715/A OR2X1_LOC_56/A 0.06fF
C43997 INPUT_0 INPUT_2 0.02fF
C43998 OR2X1_LOC_3/Y D_INPUT_6 0.08fF
C43999 AND2X1_LOC_191/B OR2X1_LOC_51/Y 0.03fF
C44000 OR2X1_LOC_625/Y OR2X1_LOC_753/a_36_216# 0.01fF
C44001 OR2X1_LOC_690/Y AND2X1_LOC_691/a_8_24# 0.00fF
C44002 AND2X1_LOC_12/Y OR2X1_LOC_34/A 0.00fF
C44003 OR2X1_LOC_154/A OR2X1_LOC_392/B 2.91fF
C44004 AND2X1_LOC_84/Y OR2X1_LOC_36/Y 0.07fF
C44005 AND2X1_LOC_43/B AND2X1_LOC_44/Y 0.08fF
C44006 OR2X1_LOC_375/A OR2X1_LOC_577/Y 0.03fF
C44007 OR2X1_LOC_91/Y OR2X1_LOC_368/Y 0.11fF
C44008 AND2X1_LOC_647/Y AND2X1_LOC_646/a_8_24# 0.04fF
C44009 AND2X1_LOC_706/Y OR2X1_LOC_432/a_36_216# 0.00fF
C44010 OR2X1_LOC_56/A AND2X1_LOC_434/a_36_24# 0.01fF
C44011 OR2X1_LOC_121/Y OR2X1_LOC_506/A 0.01fF
C44012 AND2X1_LOC_584/a_8_24# AND2X1_LOC_7/B -0.00fF
C44013 AND2X1_LOC_444/a_8_24# AND2X1_LOC_469/B 0.01fF
C44014 OR2X1_LOC_6/A AND2X1_LOC_231/a_8_24# 0.02fF
C44015 OR2X1_LOC_118/Y OR2X1_LOC_595/A 0.03fF
C44016 OR2X1_LOC_249/Y OR2X1_LOC_843/B 0.35fF
C44017 AND2X1_LOC_229/a_8_24# OR2X1_LOC_130/A 0.04fF
C44018 OR2X1_LOC_364/A OR2X1_LOC_97/A 0.08fF
C44019 OR2X1_LOC_45/B AND2X1_LOC_266/Y 1.81fF
C44020 OR2X1_LOC_185/A OR2X1_LOC_549/A 0.07fF
C44021 OR2X1_LOC_185/Y OR2X1_LOC_97/A 0.03fF
C44022 AND2X1_LOC_51/Y OR2X1_LOC_308/Y 0.02fF
C44023 OR2X1_LOC_476/B OR2X1_LOC_539/B 0.02fF
C44024 AND2X1_LOC_585/a_36_24# OR2X1_LOC_160/A 0.02fF
C44025 AND2X1_LOC_486/Y AND2X1_LOC_860/A 0.10fF
C44026 OR2X1_LOC_541/A OR2X1_LOC_778/a_8_216# 0.05fF
C44027 OR2X1_LOC_675/Y OR2X1_LOC_366/a_8_216# 0.05fF
C44028 AND2X1_LOC_43/B OR2X1_LOC_514/a_8_216# 0.01fF
C44029 AND2X1_LOC_713/Y OR2X1_LOC_48/B 0.03fF
C44030 OR2X1_LOC_776/a_8_216# AND2X1_LOC_92/Y 0.06fF
C44031 OR2X1_LOC_834/a_8_216# OR2X1_LOC_834/A 0.00fF
C44032 OR2X1_LOC_91/A AND2X1_LOC_222/a_36_24# 0.01fF
C44033 AND2X1_LOC_734/Y AND2X1_LOC_443/Y 0.00fF
C44034 OR2X1_LOC_235/B OR2X1_LOC_234/Y 0.00fF
C44035 OR2X1_LOC_600/A AND2X1_LOC_846/a_36_24# 0.00fF
C44036 OR2X1_LOC_517/A OR2X1_LOC_59/Y 0.03fF
C44037 AND2X1_LOC_95/Y OR2X1_LOC_410/Y 0.02fF
C44038 AND2X1_LOC_465/a_8_24# AND2X1_LOC_465/A 0.08fF
C44039 OR2X1_LOC_359/A OR2X1_LOC_850/B 0.03fF
C44040 AND2X1_LOC_550/a_8_24# OR2X1_LOC_427/A 0.01fF
C44041 OR2X1_LOC_659/a_36_216# OR2X1_LOC_113/B 0.00fF
C44042 OR2X1_LOC_709/A OR2X1_LOC_687/Y 0.03fF
C44043 AND2X1_LOC_70/Y OR2X1_LOC_785/B 0.01fF
C44044 AND2X1_LOC_464/A AND2X1_LOC_374/Y 0.03fF
C44045 AND2X1_LOC_575/a_8_24# AND2X1_LOC_191/Y 0.05fF
C44046 AND2X1_LOC_724/A OR2X1_LOC_36/Y 0.01fF
C44047 OR2X1_LOC_26/Y AND2X1_LOC_455/B 0.01fF
C44048 AND2X1_LOC_705/Y OR2X1_LOC_44/Y 0.01fF
C44049 OR2X1_LOC_141/B OR2X1_LOC_572/a_8_216# 0.01fF
C44050 OR2X1_LOC_154/A OR2X1_LOC_113/B 0.01fF
C44051 OR2X1_LOC_865/B VDD 0.01fF
C44052 OR2X1_LOC_92/Y AND2X1_LOC_434/Y 0.07fF
C44053 AND2X1_LOC_110/Y OR2X1_LOC_624/A 0.01fF
C44054 OR2X1_LOC_620/a_36_216# AND2X1_LOC_56/B 0.00fF
C44055 AND2X1_LOC_720/a_8_24# OR2X1_LOC_494/Y 0.01fF
C44056 OR2X1_LOC_12/Y AND2X1_LOC_361/A 0.07fF
C44057 AND2X1_LOC_213/B OR2X1_LOC_52/B 0.07fF
C44058 AND2X1_LOC_59/Y OR2X1_LOC_6/B 0.08fF
C44059 OR2X1_LOC_494/Y OR2X1_LOC_625/Y 0.03fF
C44060 VDD OR2X1_LOC_432/Y 0.16fF
C44061 OR2X1_LOC_509/A OR2X1_LOC_78/A 0.04fF
C44062 AND2X1_LOC_363/Y OR2X1_LOC_625/Y 0.05fF
C44063 OR2X1_LOC_568/a_8_216# OR2X1_LOC_365/B 0.01fF
C44064 OR2X1_LOC_405/Y AND2X1_LOC_18/Y 0.02fF
C44065 AND2X1_LOC_833/a_8_24# OR2X1_LOC_59/Y 0.02fF
C44066 OR2X1_LOC_262/Y OR2X1_LOC_595/A 0.26fF
C44067 OR2X1_LOC_653/Y AND2X1_LOC_92/Y 0.07fF
C44068 AND2X1_LOC_707/Y OR2X1_LOC_3/Y 0.14fF
C44069 OR2X1_LOC_447/a_8_216# OR2X1_LOC_66/A 0.05fF
C44070 AND2X1_LOC_11/a_36_24# INPUT_6 0.00fF
C44071 OR2X1_LOC_482/a_8_216# AND2X1_LOC_859/Y 0.04fF
C44072 AND2X1_LOC_95/Y OR2X1_LOC_244/Y 0.18fF
C44073 OR2X1_LOC_190/A OR2X1_LOC_456/a_8_216# 0.03fF
C44074 OR2X1_LOC_40/Y AND2X1_LOC_580/A 0.24fF
C44075 AND2X1_LOC_564/B OR2X1_LOC_527/Y 0.01fF
C44076 AND2X1_LOC_775/a_8_24# AND2X1_LOC_778/Y 0.12fF
C44077 VDD OR2X1_LOC_573/Y 0.00fF
C44078 OR2X1_LOC_502/A AND2X1_LOC_304/a_8_24# 0.03fF
C44079 AND2X1_LOC_84/Y OR2X1_LOC_65/a_8_216# 0.01fF
C44080 OR2X1_LOC_833/B AND2X1_LOC_92/Y 0.00fF
C44081 OR2X1_LOC_744/A OR2X1_LOC_394/Y 0.01fF
C44082 OR2X1_LOC_223/A OR2X1_LOC_777/B 0.03fF
C44083 OR2X1_LOC_130/A OR2X1_LOC_66/A 0.04fF
C44084 OR2X1_LOC_501/B AND2X1_LOC_95/Y 0.03fF
C44085 OR2X1_LOC_680/A AND2X1_LOC_657/Y 0.21fF
C44086 AND2X1_LOC_554/Y OR2X1_LOC_744/A 0.24fF
C44087 AND2X1_LOC_862/A OR2X1_LOC_59/Y 0.02fF
C44088 OR2X1_LOC_330/Y AND2X1_LOC_331/a_8_24# 0.23fF
C44089 OR2X1_LOC_538/A OR2X1_LOC_506/A 0.03fF
C44090 AND2X1_LOC_624/A OR2X1_LOC_59/Y 0.03fF
C44091 OR2X1_LOC_40/Y AND2X1_LOC_610/a_8_24# 0.10fF
C44092 AND2X1_LOC_191/B OR2X1_LOC_680/A 0.00fF
C44093 OR2X1_LOC_6/B AND2X1_LOC_495/a_8_24# 0.04fF
C44094 AND2X1_LOC_70/Y OR2X1_LOC_687/Y 0.03fF
C44095 OR2X1_LOC_485/A OR2X1_LOC_13/Y 0.01fF
C44096 OR2X1_LOC_680/A AND2X1_LOC_469/B 0.13fF
C44097 OR2X1_LOC_756/B OR2X1_LOC_555/B 0.00fF
C44098 INPUT_4 OR2X1_LOC_25/Y 0.04fF
C44099 VDD AND2X1_LOC_577/A 0.21fF
C44100 OR2X1_LOC_703/A OR2X1_LOC_212/A 0.18fF
C44101 AND2X1_LOC_721/A OR2X1_LOC_248/A 0.01fF
C44102 OR2X1_LOC_666/A OR2X1_LOC_36/Y 0.03fF
C44103 OR2X1_LOC_705/Y OR2X1_LOC_713/A 0.10fF
C44104 OR2X1_LOC_694/Y OR2X1_LOC_52/B 0.03fF
C44105 AND2X1_LOC_348/Y OR2X1_LOC_56/A 1.97fF
C44106 AND2X1_LOC_368/a_8_24# OR2X1_LOC_553/A 0.04fF
C44107 AND2X1_LOC_544/Y OR2X1_LOC_679/A 0.03fF
C44108 OR2X1_LOC_502/A AND2X1_LOC_59/a_8_24# 0.04fF
C44109 OR2X1_LOC_108/Y AND2X1_LOC_717/B 0.07fF
C44110 OR2X1_LOC_791/A OR2X1_LOC_260/Y 0.02fF
C44111 OR2X1_LOC_154/A OR2X1_LOC_147/A 0.13fF
C44112 OR2X1_LOC_139/A AND2X1_LOC_667/a_8_24# 0.00fF
C44113 OR2X1_LOC_656/Y OR2X1_LOC_660/B 0.17fF
C44114 OR2X1_LOC_753/A OR2X1_LOC_56/A 0.17fF
C44115 AND2X1_LOC_22/Y OR2X1_LOC_814/A 0.28fF
C44116 AND2X1_LOC_733/Y OR2X1_LOC_680/A 0.07fF
C44117 OR2X1_LOC_464/a_8_216# OR2X1_LOC_464/B 0.39fF
C44118 OR2X1_LOC_235/B OR2X1_LOC_204/Y 0.00fF
C44119 AND2X1_LOC_95/Y OR2X1_LOC_147/B 0.03fF
C44120 AND2X1_LOC_533/a_8_24# OR2X1_LOC_502/A 0.03fF
C44121 OR2X1_LOC_185/Y OR2X1_LOC_541/A 0.05fF
C44122 VDD OR2X1_LOC_239/Y 0.12fF
C44123 OR2X1_LOC_100/a_36_216# OR2X1_LOC_100/Y 0.00fF
C44124 OR2X1_LOC_70/Y AND2X1_LOC_778/Y 1.20fF
C44125 OR2X1_LOC_107/Y AND2X1_LOC_560/B 0.04fF
C44126 AND2X1_LOC_125/a_8_24# OR2X1_LOC_161/A 0.01fF
C44127 OR2X1_LOC_208/a_8_216# OR2X1_LOC_35/Y 0.03fF
C44128 INPUT_0 OR2X1_LOC_269/B 0.07fF
C44129 AND2X1_LOC_329/a_8_24# OR2X1_LOC_78/A 0.04fF
C44130 AND2X1_LOC_541/a_8_24# AND2X1_LOC_227/Y 0.01fF
C44131 AND2X1_LOC_500/Y OR2X1_LOC_485/A 0.09fF
C44132 OR2X1_LOC_510/Y OR2X1_LOC_574/a_8_216# 0.07fF
C44133 OR2X1_LOC_781/Y OR2X1_LOC_160/Y 0.04fF
C44134 OR2X1_LOC_326/B AND2X1_LOC_59/Y 0.00fF
C44135 AND2X1_LOC_851/B AND2X1_LOC_241/a_8_24# 0.02fF
C44136 OR2X1_LOC_95/Y OR2X1_LOC_312/a_8_216# 0.01fF
C44137 OR2X1_LOC_485/a_8_216# OR2X1_LOC_511/Y 0.02fF
C44138 OR2X1_LOC_193/A AND2X1_LOC_18/Y 0.03fF
C44139 AND2X1_LOC_356/B OR2X1_LOC_744/A 0.03fF
C44140 OR2X1_LOC_724/A OR2X1_LOC_704/a_8_216# 0.02fF
C44141 OR2X1_LOC_305/Y AND2X1_LOC_857/Y 0.02fF
C44142 OR2X1_LOC_223/A OR2X1_LOC_831/B 0.01fF
C44143 OR2X1_LOC_48/B AND2X1_LOC_436/B 0.02fF
C44144 OR2X1_LOC_280/Y OR2X1_LOC_744/A 0.46fF
C44145 OR2X1_LOC_139/a_8_216# AND2X1_LOC_41/A 0.49fF
C44146 OR2X1_LOC_771/B OR2X1_LOC_398/Y 0.03fF
C44147 OR2X1_LOC_405/A OR2X1_LOC_160/A 0.90fF
C44148 AND2X1_LOC_103/a_8_24# OR2X1_LOC_557/A 0.01fF
C44149 AND2X1_LOC_716/Y OR2X1_LOC_36/Y 0.07fF
C44150 AND2X1_LOC_553/A OR2X1_LOC_44/Y 0.03fF
C44151 AND2X1_LOC_12/Y OR2X1_LOC_506/A 0.02fF
C44152 AND2X1_LOC_716/Y OR2X1_LOC_91/a_8_216# 0.01fF
C44153 OR2X1_LOC_298/Y OR2X1_LOC_619/Y 0.04fF
C44154 OR2X1_LOC_702/A OR2X1_LOC_78/B 0.00fF
C44155 VDD OR2X1_LOC_639/A 0.00fF
C44156 OR2X1_LOC_71/A OR2X1_LOC_150/a_8_216# 0.18fF
C44157 AND2X1_LOC_199/A AND2X1_LOC_199/a_8_24# 0.19fF
C44158 OR2X1_LOC_287/B OR2X1_LOC_571/a_36_216# 0.00fF
C44159 AND2X1_LOC_321/a_8_24# AND2X1_LOC_56/B 0.04fF
C44160 OR2X1_LOC_53/Y OR2X1_LOC_47/Y 0.02fF
C44161 OR2X1_LOC_18/Y AND2X1_LOC_139/B 3.31fF
C44162 AND2X1_LOC_95/Y AND2X1_LOC_669/a_8_24# 0.01fF
C44163 OR2X1_LOC_309/Y OR2X1_LOC_22/Y 0.01fF
C44164 AND2X1_LOC_332/a_8_24# OR2X1_LOC_111/Y 0.04fF
C44165 OR2X1_LOC_772/B OR2X1_LOC_269/B 0.01fF
C44166 OR2X1_LOC_36/Y AND2X1_LOC_654/Y 0.09fF
C44167 AND2X1_LOC_448/Y AND2X1_LOC_449/Y 0.13fF
C44168 OR2X1_LOC_810/A OR2X1_LOC_574/a_8_216# 0.20fF
C44169 OR2X1_LOC_656/B OR2X1_LOC_217/Y 0.01fF
C44170 OR2X1_LOC_316/Y OR2X1_LOC_39/A 0.01fF
C44171 OR2X1_LOC_595/a_36_216# OR2X1_LOC_39/A 0.00fF
C44172 OR2X1_LOC_287/B OR2X1_LOC_392/A 0.00fF
C44173 OR2X1_LOC_421/A AND2X1_LOC_687/Y 0.02fF
C44174 OR2X1_LOC_91/A OR2X1_LOC_681/Y 0.02fF
C44175 AND2X1_LOC_514/Y AND2X1_LOC_352/B 0.03fF
C44176 OR2X1_LOC_613/Y AND2X1_LOC_621/Y 0.01fF
C44177 AND2X1_LOC_61/a_8_24# OR2X1_LOC_22/Y -0.01fF
C44178 OR2X1_LOC_26/Y OR2X1_LOC_278/Y 0.04fF
C44179 OR2X1_LOC_31/Y OR2X1_LOC_584/Y 0.32fF
C44180 OR2X1_LOC_62/B OR2X1_LOC_66/A 0.09fF
C44181 AND2X1_LOC_170/a_8_24# AND2X1_LOC_170/Y 0.01fF
C44182 D_INPUT_0 AND2X1_LOC_18/Y 0.83fF
C44183 AND2X1_LOC_502/a_8_24# OR2X1_LOC_36/Y 0.04fF
C44184 OR2X1_LOC_70/Y OR2X1_LOC_517/A 0.07fF
C44185 OR2X1_LOC_476/B OR2X1_LOC_78/B 0.10fF
C44186 OR2X1_LOC_40/Y OR2X1_LOC_72/a_8_216# 0.02fF
C44187 OR2X1_LOC_650/Y OR2X1_LOC_78/B 0.12fF
C44188 OR2X1_LOC_251/Y AND2X1_LOC_287/a_8_24# 0.01fF
C44189 AND2X1_LOC_349/B OR2X1_LOC_278/Y 0.01fF
C44190 OR2X1_LOC_489/B OR2X1_LOC_269/B 0.03fF
C44191 AND2X1_LOC_350/B OR2X1_LOC_289/Y 0.00fF
C44192 OR2X1_LOC_89/A OR2X1_LOC_278/Y 0.03fF
C44193 OR2X1_LOC_235/B OR2X1_LOC_278/A 0.00fF
C44194 OR2X1_LOC_744/A OR2X1_LOC_22/Y 0.74fF
C44195 OR2X1_LOC_511/Y OR2X1_LOC_44/Y 0.13fF
C44196 OR2X1_LOC_629/Y AND2X1_LOC_42/B 0.12fF
C44197 AND2X1_LOC_171/a_8_24# AND2X1_LOC_95/Y 0.01fF
C44198 OR2X1_LOC_427/A OR2X1_LOC_371/Y 0.07fF
C44199 AND2X1_LOC_722/A OR2X1_LOC_64/Y 0.01fF
C44200 OR2X1_LOC_419/Y AND2X1_LOC_242/a_8_24# 0.01fF
C44201 OR2X1_LOC_757/A OR2X1_LOC_815/A 0.01fF
C44202 AND2X1_LOC_158/a_8_24# OR2X1_LOC_375/A 0.04fF
C44203 OR2X1_LOC_3/B OR2X1_LOC_36/a_8_216# 0.40fF
C44204 OR2X1_LOC_74/A OR2X1_LOC_531/a_8_216# 0.01fF
C44205 OR2X1_LOC_8/Y AND2X1_LOC_835/a_36_24# 0.00fF
C44206 OR2X1_LOC_529/Y OR2X1_LOC_18/Y 0.02fF
C44207 OR2X1_LOC_474/a_8_216# OR2X1_LOC_659/A 0.01fF
C44208 OR2X1_LOC_26/Y OR2X1_LOC_95/a_8_216# 0.01fF
C44209 OR2X1_LOC_678/Y AND2X1_LOC_48/A 0.32fF
C44210 AND2X1_LOC_1/Y D_INPUT_4 0.03fF
C44211 AND2X1_LOC_845/Y OR2X1_LOC_56/A 0.10fF
C44212 AND2X1_LOC_3/Y OR2X1_LOC_347/B 0.01fF
C44213 AND2X1_LOC_19/Y OR2X1_LOC_655/B 0.03fF
C44214 AND2X1_LOC_184/a_36_24# AND2X1_LOC_47/Y 0.00fF
C44215 AND2X1_LOC_42/B OR2X1_LOC_249/a_8_216# 0.01fF
C44216 AND2X1_LOC_3/Y OR2X1_LOC_539/Y 0.03fF
C44217 OR2X1_LOC_592/A OR2X1_LOC_799/A 0.03fF
C44218 OR2X1_LOC_859/A OR2X1_LOC_571/a_8_216# 0.08fF
C44219 OR2X1_LOC_468/A OR2X1_LOC_468/a_8_216# 0.18fF
C44220 OR2X1_LOC_859/A OR2X1_LOC_659/A 0.76fF
C44221 OR2X1_LOC_51/Y OR2X1_LOC_411/a_8_216# 0.01fF
C44222 OR2X1_LOC_756/B AND2X1_LOC_600/a_8_24# 0.07fF
C44223 OR2X1_LOC_696/A OR2X1_LOC_589/Y 0.01fF
C44224 AND2X1_LOC_572/a_8_24# AND2X1_LOC_657/A 0.01fF
C44225 OR2X1_LOC_114/B OR2X1_LOC_284/B 0.05fF
C44226 OR2X1_LOC_774/Y OR2X1_LOC_772/a_36_216# 0.00fF
C44227 AND2X1_LOC_580/A OR2X1_LOC_7/A 0.03fF
C44228 OR2X1_LOC_377/A OR2X1_LOC_863/B 0.02fF
C44229 OR2X1_LOC_392/B OR2X1_LOC_560/A 0.03fF
C44230 AND2X1_LOC_711/Y AND2X1_LOC_624/A 0.00fF
C44231 OR2X1_LOC_426/B AND2X1_LOC_318/Y 0.02fF
C44232 AND2X1_LOC_8/Y OR2X1_LOC_753/A 0.70fF
C44233 AND2X1_LOC_211/B AND2X1_LOC_354/B 0.03fF
C44234 OR2X1_LOC_168/B AND2X1_LOC_47/Y 0.01fF
C44235 OR2X1_LOC_250/a_8_216# OR2X1_LOC_64/Y 0.01fF
C44236 OR2X1_LOC_114/B D_INPUT_1 0.03fF
C44237 OR2X1_LOC_70/Y AND2X1_LOC_624/A 0.05fF
C44238 AND2X1_LOC_464/a_8_24# OR2X1_LOC_371/Y 0.02fF
C44239 AND2X1_LOC_56/B OR2X1_LOC_445/a_8_216# 0.06fF
C44240 OR2X1_LOC_26/Y AND2X1_LOC_634/a_8_24# 0.02fF
C44241 OR2X1_LOC_114/Y OR2X1_LOC_574/A 0.00fF
C44242 OR2X1_LOC_856/B OR2X1_LOC_750/A 0.13fF
C44243 OR2X1_LOC_97/A AND2X1_LOC_432/a_8_24# 0.01fF
C44244 OR2X1_LOC_51/Y OR2X1_LOC_146/Y 0.05fF
C44245 OR2X1_LOC_141/B OR2X1_LOC_643/A 0.03fF
C44246 OR2X1_LOC_297/Y OR2X1_LOC_44/Y 0.02fF
C44247 AND2X1_LOC_722/A OR2X1_LOC_417/A 0.09fF
C44248 OR2X1_LOC_119/a_8_216# OR2X1_LOC_65/B 0.00fF
C44249 AND2X1_LOC_70/Y OR2X1_LOC_786/Y 0.01fF
C44250 OR2X1_LOC_141/B OR2X1_LOC_124/Y 0.00fF
C44251 OR2X1_LOC_97/A OR2X1_LOC_578/B 0.03fF
C44252 OR2X1_LOC_470/B OR2X1_LOC_470/A 0.08fF
C44253 OR2X1_LOC_76/Y OR2X1_LOC_445/a_36_216# 0.00fF
C44254 OR2X1_LOC_240/B OR2X1_LOC_19/B 0.21fF
C44255 AND2X1_LOC_345/Y OR2X1_LOC_44/Y 0.01fF
C44256 OR2X1_LOC_723/a_8_216# OR2X1_LOC_374/Y 0.01fF
C44257 OR2X1_LOC_272/Y AND2X1_LOC_361/A 0.00fF
C44258 AND2X1_LOC_346/a_36_24# AND2X1_LOC_848/A 0.01fF
C44259 VDD OR2X1_LOC_493/Y 1.69fF
C44260 OR2X1_LOC_291/A OR2X1_LOC_753/A 0.08fF
C44261 OR2X1_LOC_476/B OR2X1_LOC_375/A 0.07fF
C44262 OR2X1_LOC_161/B OR2X1_LOC_365/a_8_216# -0.03fF
C44263 AND2X1_LOC_307/a_8_24# OR2X1_LOC_36/Y 0.01fF
C44264 OR2X1_LOC_620/Y OR2X1_LOC_532/B 0.00fF
C44265 OR2X1_LOC_273/Y OR2X1_LOC_26/Y 0.09fF
C44266 OR2X1_LOC_650/Y OR2X1_LOC_375/A 0.03fF
C44267 OR2X1_LOC_113/B OR2X1_LOC_560/A 0.00fF
C44268 OR2X1_LOC_599/A OR2X1_LOC_64/Y 0.17fF
C44269 OR2X1_LOC_187/a_8_216# GATE_662 0.48fF
C44270 OR2X1_LOC_99/B OR2X1_LOC_99/a_8_216# 0.00fF
C44271 AND2X1_LOC_59/Y OR2X1_LOC_68/Y 0.09fF
C44272 AND2X1_LOC_153/a_8_24# OR2X1_LOC_814/A 0.03fF
C44273 OR2X1_LOC_661/A OR2X1_LOC_68/B 0.01fF
C44274 AND2X1_LOC_516/a_8_24# AND2X1_LOC_51/Y 0.06fF
C44275 AND2X1_LOC_11/Y OR2X1_LOC_639/a_36_216# 0.00fF
C44276 OR2X1_LOC_504/Y AND2X1_LOC_862/A 0.03fF
C44277 OR2X1_LOC_673/Y AND2X1_LOC_134/a_8_24# 0.01fF
C44278 OR2X1_LOC_504/Y AND2X1_LOC_624/A 0.13fF
C44279 OR2X1_LOC_648/A OR2X1_LOC_358/A 0.01fF
C44280 OR2X1_LOC_739/B AND2X1_LOC_47/Y 0.02fF
C44281 OR2X1_LOC_19/B OR2X1_LOC_26/Y 0.14fF
C44282 INPUT_5 OR2X1_LOC_3/B 0.77fF
C44283 OR2X1_LOC_649/B AND2X1_LOC_48/A 0.05fF
C44284 OR2X1_LOC_739/B D_GATE_222 0.05fF
C44285 AND2X1_LOC_59/Y AND2X1_LOC_47/Y 0.42fF
C44286 OR2X1_LOC_22/Y OR2X1_LOC_74/a_8_216# 0.05fF
C44287 OR2X1_LOC_628/a_8_216# OR2X1_LOC_47/Y 0.01fF
C44288 OR2X1_LOC_154/A OR2X1_LOC_532/B 0.33fF
C44289 OR2X1_LOC_45/B OR2X1_LOC_268/Y 0.54fF
C44290 OR2X1_LOC_416/a_8_216# OR2X1_LOC_39/A 0.01fF
C44291 OR2X1_LOC_636/a_8_216# AND2X1_LOC_51/Y 0.01fF
C44292 OR2X1_LOC_45/B OR2X1_LOC_183/Y 0.02fF
C44293 AND2X1_LOC_64/Y OR2X1_LOC_140/B 0.09fF
C44294 AND2X1_LOC_729/B OR2X1_LOC_829/Y 0.14fF
C44295 INPUT_1 OR2X1_LOC_240/A 0.04fF
C44296 AND2X1_LOC_68/a_8_24# OR2X1_LOC_585/A 0.02fF
C44297 AND2X1_LOC_849/A OR2X1_LOC_279/Y 0.04fF
C44298 OR2X1_LOC_691/B AND2X1_LOC_36/Y 0.03fF
C44299 OR2X1_LOC_160/A OR2X1_LOC_779/Y 0.00fF
C44300 OR2X1_LOC_276/A OR2X1_LOC_203/Y 0.04fF
C44301 AND2X1_LOC_12/Y D_INPUT_1 0.11fF
C44302 AND2X1_LOC_560/B AND2X1_LOC_866/A 0.07fF
C44303 OR2X1_LOC_416/Y OR2X1_LOC_27/Y 0.02fF
C44304 OR2X1_LOC_461/Y OR2X1_LOC_19/B 0.00fF
C44305 OR2X1_LOC_377/A AND2X1_LOC_6/a_36_24# 0.00fF
C44306 AND2X1_LOC_711/Y AND2X1_LOC_621/a_8_24# 0.01fF
C44307 OR2X1_LOC_777/a_8_216# OR2X1_LOC_777/B 0.06fF
C44308 OR2X1_LOC_348/Y OR2X1_LOC_580/A 0.59fF
C44309 AND2X1_LOC_838/Y D_INPUT_1 0.04fF
C44310 OR2X1_LOC_19/B AND2X1_LOC_51/Y 0.03fF
C44311 OR2X1_LOC_271/Y AND2X1_LOC_851/B 0.03fF
C44312 OR2X1_LOC_160/A OR2X1_LOC_330/a_8_216# 0.01fF
C44313 OR2X1_LOC_12/Y OR2X1_LOC_387/A 0.03fF
C44314 OR2X1_LOC_349/a_8_216# OR2X1_LOC_580/A 0.04fF
C44315 AND2X1_LOC_648/B OR2X1_LOC_44/Y 0.02fF
C44316 OR2X1_LOC_405/A OR2X1_LOC_717/a_8_216# 0.03fF
C44317 OR2X1_LOC_856/a_8_216# OR2X1_LOC_532/B 0.01fF
C44318 VDD OR2X1_LOC_532/a_8_216# 0.21fF
C44319 OR2X1_LOC_188/a_36_216# OR2X1_LOC_121/A 0.00fF
C44320 OR2X1_LOC_280/Y OR2X1_LOC_31/Y 0.22fF
C44321 AND2X1_LOC_729/B OR2X1_LOC_7/Y 0.09fF
C44322 AND2X1_LOC_18/Y OR2X1_LOC_339/A 0.07fF
C44323 AND2X1_LOC_95/Y OR2X1_LOC_318/B 0.08fF
C44324 AND2X1_LOC_502/a_8_24# OR2X1_LOC_419/Y 0.07fF
C44325 OR2X1_LOC_116/a_8_216# OR2X1_LOC_786/Y 0.01fF
C44326 OR2X1_LOC_427/A AND2X1_LOC_222/Y 0.03fF
C44327 OR2X1_LOC_405/a_8_216# OR2X1_LOC_358/A 0.00fF
C44328 AND2X1_LOC_476/A OR2X1_LOC_7/A 0.09fF
C44329 OR2X1_LOC_532/B OR2X1_LOC_778/A 0.00fF
C44330 AND2X1_LOC_416/a_8_24# AND2X1_LOC_44/Y 0.01fF
C44331 OR2X1_LOC_87/A AND2X1_LOC_418/a_8_24# 0.02fF
C44332 AND2X1_LOC_367/A AND2X1_LOC_212/a_8_24# 0.20fF
C44333 AND2X1_LOC_59/Y OR2X1_LOC_598/A 0.01fF
C44334 OR2X1_LOC_759/A AND2X1_LOC_789/Y 0.02fF
C44335 OR2X1_LOC_632/Y OR2X1_LOC_501/a_36_216# 0.01fF
C44336 OR2X1_LOC_836/Y OR2X1_LOC_19/B 0.04fF
C44337 OR2X1_LOC_756/B OR2X1_LOC_579/a_8_216# 0.02fF
C44338 AND2X1_LOC_580/B AND2X1_LOC_792/Y 0.04fF
C44339 OR2X1_LOC_590/a_36_216# OR2X1_LOC_375/A 0.00fF
C44340 AND2X1_LOC_101/B OR2X1_LOC_813/Y 0.09fF
C44341 OR2X1_LOC_7/a_36_216# OR2X1_LOC_7/Y 0.00fF
C44342 OR2X1_LOC_39/A OR2X1_LOC_153/a_8_216# 0.02fF
C44343 OR2X1_LOC_380/A OR2X1_LOC_70/A 0.04fF
C44344 OR2X1_LOC_64/Y AND2X1_LOC_866/A 0.03fF
C44345 OR2X1_LOC_703/A OR2X1_LOC_181/Y 0.15fF
C44346 AND2X1_LOC_496/a_8_24# D_INPUT_1 0.02fF
C44347 AND2X1_LOC_573/A OR2X1_LOC_80/A 0.03fF
C44348 OR2X1_LOC_709/a_8_216# AND2X1_LOC_7/B 0.00fF
C44349 OR2X1_LOC_19/B OR2X1_LOC_92/a_8_216# 0.01fF
C44350 OR2X1_LOC_434/A OR2X1_LOC_814/A 0.01fF
C44351 OR2X1_LOC_22/Y OR2X1_LOC_31/Y 0.54fF
C44352 OR2X1_LOC_577/Y OR2X1_LOC_549/A 0.11fF
C44353 OR2X1_LOC_848/B OR2X1_LOC_561/B 0.04fF
C44354 OR2X1_LOC_502/A OR2X1_LOC_777/B 0.12fF
C44355 OR2X1_LOC_813/A D_INPUT_0 0.03fF
C44356 OR2X1_LOC_698/Y AND2X1_LOC_789/Y 0.00fF
C44357 AND2X1_LOC_719/Y AND2X1_LOC_721/Y 0.01fF
C44358 AND2X1_LOC_64/Y OR2X1_LOC_851/a_8_216# 0.01fF
C44359 AND2X1_LOC_284/a_8_24# AND2X1_LOC_243/Y 0.01fF
C44360 AND2X1_LOC_370/a_36_24# AND2X1_LOC_182/A 0.00fF
C44361 OR2X1_LOC_134/a_8_216# AND2X1_LOC_772/B 0.47fF
C44362 AND2X1_LOC_227/Y OR2X1_LOC_226/a_8_216# 0.01fF
C44363 OR2X1_LOC_205/a_36_216# OR2X1_LOC_560/A 0.00fF
C44364 AND2X1_LOC_773/Y AND2X1_LOC_566/B 0.03fF
C44365 OR2X1_LOC_250/Y OR2X1_LOC_13/B 0.91fF
C44366 OR2X1_LOC_43/A OR2X1_LOC_534/Y 0.44fF
C44367 OR2X1_LOC_62/B OR2X1_LOC_84/A 0.02fF
C44368 AND2X1_LOC_656/Y OR2X1_LOC_95/Y 0.05fF
C44369 AND2X1_LOC_626/a_8_24# AND2X1_LOC_256/a_8_24# 0.23fF
C44370 OR2X1_LOC_363/B OR2X1_LOC_362/a_8_216# 0.39fF
C44371 AND2X1_LOC_866/A OR2X1_LOC_417/A 0.17fF
C44372 OR2X1_LOC_808/A OR2X1_LOC_605/Y 0.01fF
C44373 OR2X1_LOC_91/Y OR2X1_LOC_437/A 0.12fF
C44374 OR2X1_LOC_47/Y INPUT_1 0.25fF
C44375 AND2X1_LOC_7/B OR2X1_LOC_702/a_8_216# 0.01fF
C44376 AND2X1_LOC_22/Y OR2X1_LOC_244/Y 0.07fF
C44377 OR2X1_LOC_858/A OR2X1_LOC_563/A 0.07fF
C44378 OR2X1_LOC_604/A AND2X1_LOC_724/A 0.03fF
C44379 OR2X1_LOC_329/B AND2X1_LOC_242/B 0.02fF
C44380 OR2X1_LOC_158/A OR2X1_LOC_382/a_8_216# 0.01fF
C44381 AND2X1_LOC_362/B OR2X1_LOC_106/a_8_216# 0.07fF
C44382 OR2X1_LOC_36/Y OR2X1_LOC_599/a_36_216# 0.03fF
C44383 AND2X1_LOC_719/Y OR2X1_LOC_482/Y 0.03fF
C44384 OR2X1_LOC_465/B OR2X1_LOC_367/B 0.03fF
C44385 AND2X1_LOC_857/Y OR2X1_LOC_171/Y 0.83fF
C44386 OR2X1_LOC_516/A OR2X1_LOC_142/Y 0.03fF
C44387 OR2X1_LOC_36/Y OR2X1_LOC_13/B 1.08fF
C44388 AND2X1_LOC_61/Y OR2X1_LOC_12/Y 0.10fF
C44389 OR2X1_LOC_532/B AND2X1_LOC_6/a_8_24# 0.01fF
C44390 OR2X1_LOC_494/A AND2X1_LOC_367/A 0.01fF
C44391 OR2X1_LOC_756/B OR2X1_LOC_362/a_8_216# 0.15fF
C44392 OR2X1_LOC_161/A OR2X1_LOC_301/a_8_216# 0.01fF
C44393 AND2X1_LOC_40/Y AND2X1_LOC_258/a_8_24# 0.05fF
C44394 OR2X1_LOC_193/A OR2X1_LOC_789/A 0.02fF
C44395 AND2X1_LOC_662/B AND2X1_LOC_269/a_36_24# 0.01fF
C44396 OR2X1_LOC_607/Y AND2X1_LOC_646/a_8_24# 0.23fF
C44397 AND2X1_LOC_568/B AND2X1_LOC_566/B 0.01fF
C44398 AND2X1_LOC_784/Y OR2X1_LOC_600/A 0.02fF
C44399 OR2X1_LOC_506/A OR2X1_LOC_356/B 0.43fF
C44400 OR2X1_LOC_49/A OR2X1_LOC_634/A 0.01fF
C44401 AND2X1_LOC_505/a_8_24# AND2X1_LOC_18/Y 0.03fF
C44402 OR2X1_LOC_736/A AND2X1_LOC_248/a_8_24# 0.01fF
C44403 OR2X1_LOC_508/a_8_216# AND2X1_LOC_41/A 0.01fF
C44404 AND2X1_LOC_388/Y OR2X1_LOC_166/Y 0.29fF
C44405 OR2X1_LOC_702/A OR2X1_LOC_515/Y 0.10fF
C44406 AND2X1_LOC_387/B AND2X1_LOC_41/Y 0.14fF
C44407 AND2X1_LOC_41/A OR2X1_LOC_486/Y 0.01fF
C44408 OR2X1_LOC_604/A OR2X1_LOC_666/A 0.05fF
C44409 OR2X1_LOC_468/A OR2X1_LOC_66/A 0.08fF
C44410 AND2X1_LOC_724/Y AND2X1_LOC_732/a_8_24# 0.09fF
C44411 OR2X1_LOC_379/Y OR2X1_LOC_855/A 0.00fF
C44412 OR2X1_LOC_485/Y OR2X1_LOC_744/A 0.27fF
C44413 OR2X1_LOC_40/Y INPUT_0 0.15fF
C44414 OR2X1_LOC_158/A AND2X1_LOC_197/Y 0.07fF
C44415 OR2X1_LOC_508/A OR2X1_LOC_508/a_8_216# -0.04fF
C44416 OR2X1_LOC_600/A AND2X1_LOC_434/Y 0.15fF
C44417 AND2X1_LOC_364/a_8_24# AND2X1_LOC_364/A 0.04fF
C44418 OR2X1_LOC_837/B OR2X1_LOC_414/Y 0.04fF
C44419 OR2X1_LOC_532/B OR2X1_LOC_560/A 0.20fF
C44420 OR2X1_LOC_529/Y OR2X1_LOC_183/a_36_216# 0.00fF
C44421 OR2X1_LOC_117/a_8_216# AND2X1_LOC_99/A 0.03fF
C44422 OR2X1_LOC_833/a_8_216# OR2X1_LOC_549/A 0.01fF
C44423 OR2X1_LOC_177/Y AND2X1_LOC_716/Y 0.02fF
C44424 OR2X1_LOC_532/B OR2X1_LOC_198/A 0.16fF
C44425 OR2X1_LOC_135/a_8_216# OR2X1_LOC_48/B 0.01fF
C44426 VDD AND2X1_LOC_144/a_8_24# -0.00fF
C44427 OR2X1_LOC_335/a_8_216# OR2X1_LOC_87/A 0.02fF
C44428 OR2X1_LOC_160/B OR2X1_LOC_624/a_8_216# 0.02fF
C44429 AND2X1_LOC_76/Y OR2X1_LOC_522/Y 0.21fF
C44430 OR2X1_LOC_703/A AND2X1_LOC_323/a_8_24# 0.00fF
C44431 OR2X1_LOC_336/a_8_216# OR2X1_LOC_212/A 0.40fF
C44432 OR2X1_LOC_323/A OR2X1_LOC_26/Y 0.03fF
C44433 AND2X1_LOC_465/A OR2X1_LOC_44/Y 0.07fF
C44434 AND2X1_LOC_191/B OR2X1_LOC_757/A 0.00fF
C44435 AND2X1_LOC_456/B OR2X1_LOC_666/a_8_216# 0.01fF
C44436 AND2X1_LOC_22/Y AND2X1_LOC_669/a_8_24# 0.08fF
C44437 OR2X1_LOC_589/A AND2X1_LOC_364/A 0.06fF
C44438 AND2X1_LOC_434/a_8_24# OR2X1_LOC_59/Y 0.02fF
C44439 OR2X1_LOC_380/a_8_216# OR2X1_LOC_26/a_8_216# 0.47fF
C44440 OR2X1_LOC_185/Y OR2X1_LOC_175/Y 0.03fF
C44441 AND2X1_LOC_286/a_36_24# OR2X1_LOC_59/Y 0.00fF
C44442 OR2X1_LOC_510/Y AND2X1_LOC_44/Y 1.52fF
C44443 OR2X1_LOC_244/B OR2X1_LOC_244/Y 0.01fF
C44444 OR2X1_LOC_659/A OR2X1_LOC_66/A 0.09fF
C44445 AND2X1_LOC_452/Y OR2X1_LOC_16/A 0.07fF
C44446 AND2X1_LOC_88/Y OR2X1_LOC_559/a_8_216# 0.01fF
C44447 OR2X1_LOC_363/B OR2X1_LOC_756/B 0.28fF
C44448 AND2X1_LOC_482/a_36_24# OR2X1_LOC_736/Y 0.01fF
C44449 OR2X1_LOC_49/A OR2X1_LOC_94/a_8_216# 0.03fF
C44450 OR2X1_LOC_833/Y OR2X1_LOC_541/B 0.32fF
C44451 AND2X1_LOC_706/Y OR2X1_LOC_433/Y 0.06fF
C44452 AND2X1_LOC_534/a_8_24# OR2X1_LOC_161/A 0.01fF
C44453 OR2X1_LOC_59/Y OR2X1_LOC_755/a_8_216# 0.03fF
C44454 OR2X1_LOC_715/B AND2X1_LOC_492/a_8_24# 0.03fF
C44455 AND2X1_LOC_717/Y OR2X1_LOC_40/Y 0.00fF
C44456 AND2X1_LOC_40/Y AND2X1_LOC_18/Y 1.06fF
C44457 OR2X1_LOC_235/B OR2X1_LOC_78/A 0.09fF
C44458 OR2X1_LOC_200/a_8_216# AND2X1_LOC_7/B 0.03fF
C44459 AND2X1_LOC_541/a_36_24# AND2X1_LOC_361/A 0.00fF
C44460 AND2X1_LOC_7/B OR2X1_LOC_269/B 0.99fF
C44461 AND2X1_LOC_1/a_8_24# INPUT_7 0.01fF
C44462 OR2X1_LOC_124/A OR2X1_LOC_663/A 0.05fF
C44463 OR2X1_LOC_185/Y OR2X1_LOC_691/Y 0.03fF
C44464 OR2X1_LOC_351/B AND2X1_LOC_95/Y 0.26fF
C44465 OR2X1_LOC_756/B AND2X1_LOC_616/a_36_24# 0.01fF
C44466 OR2X1_LOC_89/A OR2X1_LOC_89/Y 0.14fF
C44467 OR2X1_LOC_482/Y OR2X1_LOC_252/Y 0.01fF
C44468 AND2X1_LOC_159/a_8_24# AND2X1_LOC_44/Y 0.01fF
C44469 OR2X1_LOC_644/B OR2X1_LOC_161/B -0.02fF
C44470 OR2X1_LOC_114/B AND2X1_LOC_95/Y 0.08fF
C44471 OR2X1_LOC_810/A AND2X1_LOC_44/Y 0.05fF
C44472 OR2X1_LOC_375/A AND2X1_LOC_262/a_8_24# 0.01fF
C44473 OR2X1_LOC_802/a_8_216# OR2X1_LOC_78/B 0.01fF
C44474 AND2X1_LOC_22/Y AND2X1_LOC_171/a_8_24# 0.02fF
C44475 VDD OR2X1_LOC_194/B -0.00fF
C44476 OR2X1_LOC_404/A AND2X1_LOC_36/Y 0.16fF
C44477 AND2X1_LOC_110/Y OR2X1_LOC_161/A 0.06fF
C44478 D_INPUT_3 OR2X1_LOC_437/A 0.07fF
C44479 AND2X1_LOC_852/Y OR2X1_LOC_12/Y 6.26fF
C44480 OR2X1_LOC_438/Y OR2X1_LOC_524/Y 0.08fF
C44481 OR2X1_LOC_97/A OR2X1_LOC_654/A 0.00fF
C44482 AND2X1_LOC_22/Y AND2X1_LOC_387/B 0.09fF
C44483 AND2X1_LOC_364/Y OR2X1_LOC_92/Y 0.03fF
C44484 OR2X1_LOC_186/Y OR2X1_LOC_778/Y 0.05fF
C44485 OR2X1_LOC_631/B OR2X1_LOC_486/Y 0.09fF
C44486 OR2X1_LOC_40/Y OR2X1_LOC_11/Y 0.04fF
C44487 OR2X1_LOC_787/Y AND2X1_LOC_604/a_8_24# 0.02fF
C44488 OR2X1_LOC_696/A AND2X1_LOC_537/Y 0.01fF
C44489 OR2X1_LOC_666/A AND2X1_LOC_850/a_8_24# 0.01fF
C44490 AND2X1_LOC_719/Y AND2X1_LOC_859/a_36_24# 0.06fF
C44491 OR2X1_LOC_484/a_8_216# OR2X1_LOC_48/B 0.04fF
C44492 OR2X1_LOC_7/A OR2X1_LOC_766/a_8_216# 0.05fF
C44493 OR2X1_LOC_280/Y AND2X1_LOC_464/A 0.03fF
C44494 OR2X1_LOC_302/a_8_216# OR2X1_LOC_620/Y 0.02fF
C44495 AND2X1_LOC_61/a_8_24# OR2X1_LOC_39/A 0.08fF
C44496 AND2X1_LOC_658/B AND2X1_LOC_624/A 26.34fF
C44497 AND2X1_LOC_388/Y OR2X1_LOC_43/A 0.26fF
C44498 OR2X1_LOC_177/Y OR2X1_LOC_312/Y 0.92fF
C44499 OR2X1_LOC_87/Y AND2X1_LOC_18/Y 0.00fF
C44500 AND2X1_LOC_788/a_8_24# AND2X1_LOC_645/A 0.03fF
C44501 OR2X1_LOC_215/A AND2X1_LOC_7/B 0.10fF
C44502 OR2X1_LOC_102/a_36_216# OR2X1_LOC_585/A 0.00fF
C44503 OR2X1_LOC_501/B OR2X1_LOC_630/a_8_216# 0.05fF
C44504 AND2X1_LOC_705/a_8_24# OR2X1_LOC_511/Y 0.01fF
C44505 AND2X1_LOC_356/a_8_24# AND2X1_LOC_434/Y 0.01fF
C44506 OR2X1_LOC_604/A GATE_366 0.07fF
C44507 AND2X1_LOC_729/Y AND2X1_LOC_738/B 0.10fF
C44508 AND2X1_LOC_367/A OR2X1_LOC_427/A 0.22fF
C44509 AND2X1_LOC_70/Y OR2X1_LOC_828/B 0.03fF
C44510 OR2X1_LOC_641/Y OR2X1_LOC_520/Y 0.13fF
C44511 OR2X1_LOC_160/A AND2X1_LOC_19/Y 0.01fF
C44512 OR2X1_LOC_168/B OR2X1_LOC_506/A 0.19fF
C44513 AND2X1_LOC_729/Y OR2X1_LOC_56/A 0.04fF
C44514 OR2X1_LOC_3/Y AND2X1_LOC_770/a_8_24# 0.01fF
C44515 AND2X1_LOC_95/Y OR2X1_LOC_538/A 0.03fF
C44516 OR2X1_LOC_476/a_8_216# OR2X1_LOC_392/B 0.04fF
C44517 OR2X1_LOC_743/A OR2X1_LOC_829/A 0.71fF
C44518 OR2X1_LOC_40/Y OR2X1_LOC_173/Y 0.01fF
C44519 AND2X1_LOC_181/Y OR2X1_LOC_529/Y 0.01fF
C44520 OR2X1_LOC_287/B OR2X1_LOC_349/A 0.25fF
C44521 OR2X1_LOC_744/A OR2X1_LOC_39/A 1.56fF
C44522 AND2X1_LOC_56/B OR2X1_LOC_35/a_8_216# 0.01fF
C44523 AND2X1_LOC_47/Y AND2X1_LOC_762/a_8_24# 0.01fF
C44524 OR2X1_LOC_703/A OR2X1_LOC_220/B 0.83fF
C44525 OR2X1_LOC_6/B OR2X1_LOC_585/A 0.38fF
C44526 AND2X1_LOC_70/Y OR2X1_LOC_204/Y 0.00fF
C44527 OR2X1_LOC_85/a_8_216# OR2X1_LOC_13/B 0.19fF
C44528 OR2X1_LOC_3/Y OR2X1_LOC_589/A 0.02fF
C44529 OR2X1_LOC_309/Y AND2X1_LOC_211/B 0.04fF
C44530 AND2X1_LOC_345/Y OR2X1_LOC_382/A 0.02fF
C44531 VDD OR2X1_LOC_836/a_8_216# 0.21fF
C44532 AND2X1_LOC_580/A OR2X1_LOC_531/Y 0.01fF
C44533 OR2X1_LOC_181/B OR2X1_LOC_190/B 0.05fF
C44534 OR2X1_LOC_604/A OR2X1_LOC_312/Y 0.01fF
C44535 AND2X1_LOC_658/A AND2X1_LOC_859/Y 0.07fF
C44536 OR2X1_LOC_419/Y OR2X1_LOC_13/B 0.10fF
C44537 OR2X1_LOC_449/B OR2X1_LOC_66/A 0.87fF
C44538 OR2X1_LOC_532/Y OR2X1_LOC_330/a_8_216# 0.40fF
C44539 AND2X1_LOC_810/A AND2X1_LOC_307/Y 0.01fF
C44540 OR2X1_LOC_154/A OR2X1_LOC_624/Y 0.00fF
C44541 AND2X1_LOC_40/Y OR2X1_LOC_807/B 0.23fF
C44542 OR2X1_LOC_264/a_8_216# OR2X1_LOC_78/B 0.35fF
C44543 OR2X1_LOC_319/B OR2X1_LOC_739/A 0.03fF
C44544 AND2X1_LOC_784/A OR2X1_LOC_56/A 0.10fF
C44545 OR2X1_LOC_814/A OR2X1_LOC_227/B 0.48fF
C44546 AND2X1_LOC_391/Y OR2X1_LOC_6/A 0.37fF
C44547 AND2X1_LOC_12/Y OR2X1_LOC_391/a_8_216# 0.01fF
C44548 OR2X1_LOC_226/Y AND2X1_LOC_227/a_8_24# 0.01fF
C44549 AND2X1_LOC_184/a_8_24# AND2X1_LOC_3/Y 0.01fF
C44550 OR2X1_LOC_91/A OR2X1_LOC_6/A 0.15fF
C44551 AND2X1_LOC_310/a_8_24# OR2X1_LOC_778/Y 0.17fF
C44552 OR2X1_LOC_669/a_8_216# OR2X1_LOC_59/Y 0.05fF
C44553 AND2X1_LOC_778/a_8_24# OR2X1_LOC_56/A 0.01fF
C44554 OR2X1_LOC_95/Y AND2X1_LOC_772/Y 0.03fF
C44555 OR2X1_LOC_526/Y OR2X1_LOC_485/A 0.01fF
C44556 OR2X1_LOC_625/Y OR2X1_LOC_628/a_8_216# 0.08fF
C44557 OR2X1_LOC_45/B AND2X1_LOC_640/a_8_24# 0.01fF
C44558 AND2X1_LOC_803/B AND2X1_LOC_191/Y 0.03fF
C44559 OR2X1_LOC_754/a_8_216# AND2X1_LOC_285/Y 0.14fF
C44560 OR2X1_LOC_631/B OR2X1_LOC_632/a_36_216# 0.00fF
C44561 OR2X1_LOC_566/a_8_216# OR2X1_LOC_303/B 0.01fF
C44562 OR2X1_LOC_161/A OR2X1_LOC_712/a_36_216# 0.01fF
C44563 AND2X1_LOC_339/B AND2X1_LOC_358/a_8_24# 0.01fF
C44564 OR2X1_LOC_507/a_8_216# AND2X1_LOC_81/B 0.01fF
C44565 OR2X1_LOC_105/Y AND2X1_LOC_251/a_8_24# 0.11fF
C44566 AND2X1_LOC_793/Y AND2X1_LOC_793/a_8_24# 0.01fF
C44567 OR2X1_LOC_3/Y OR2X1_LOC_261/a_8_216# 0.01fF
C44568 AND2X1_LOC_568/a_36_24# OR2X1_LOC_600/A 0.00fF
C44569 AND2X1_LOC_12/Y OR2X1_LOC_737/A 0.07fF
C44570 OR2X1_LOC_744/A AND2X1_LOC_211/B 0.07fF
C44571 OR2X1_LOC_405/A OR2X1_LOC_447/A 0.01fF
C44572 OR2X1_LOC_264/Y AND2X1_LOC_81/B 0.03fF
C44573 AND2X1_LOC_367/A AND2X1_LOC_363/A 0.14fF
C44574 AND2X1_LOC_110/Y AND2X1_LOC_51/Y 0.03fF
C44575 OR2X1_LOC_40/Y OR2X1_LOC_64/Y 0.28fF
C44576 OR2X1_LOC_68/B OR2X1_LOC_561/A 0.05fF
C44577 INPUT_0 OR2X1_LOC_7/A 0.03fF
C44578 AND2X1_LOC_723/Y OR2X1_LOC_26/Y 0.07fF
C44579 OR2X1_LOC_596/Y AND2X1_LOC_40/Y 0.01fF
C44580 AND2X1_LOC_700/a_8_24# OR2X1_LOC_705/Y 0.02fF
C44581 OR2X1_LOC_477/a_8_216# OR2X1_LOC_161/B 0.01fF
C44582 AND2X1_LOC_12/Y AND2X1_LOC_95/Y 14.07fF
C44583 OR2X1_LOC_451/B AND2X1_LOC_581/a_8_24# 0.01fF
C44584 AND2X1_LOC_476/A AND2X1_LOC_476/a_8_24# 0.11fF
C44585 OR2X1_LOC_154/A OR2X1_LOC_714/Y 0.04fF
C44586 OR2X1_LOC_844/a_8_216# OR2X1_LOC_78/A 0.14fF
C44587 AND2X1_LOC_42/B OR2X1_LOC_778/B 0.14fF
C44588 AND2X1_LOC_59/Y OR2X1_LOC_506/A 0.04fF
C44589 VDD AND2X1_LOC_842/B 0.18fF
C44590 OR2X1_LOC_70/Y AND2X1_LOC_434/a_8_24# 0.01fF
C44591 OR2X1_LOC_45/B AND2X1_LOC_649/Y 0.01fF
C44592 OR2X1_LOC_294/a_8_216# AND2X1_LOC_3/Y 0.15fF
C44593 OR2X1_LOC_755/Y OR2X1_LOC_757/Y 0.05fF
C44594 OR2X1_LOC_374/Y OR2X1_LOC_605/Y 0.04fF
C44595 OR2X1_LOC_697/a_8_216# OR2X1_LOC_743/A 0.01fF
C44596 OR2X1_LOC_194/Y AND2X1_LOC_16/a_8_24# 0.05fF
C44597 AND2X1_LOC_59/Y OR2X1_LOC_341/Y 0.01fF
C44598 AND2X1_LOC_711/Y OR2X1_LOC_755/a_8_216# 0.01fF
C44599 OR2X1_LOC_121/B OR2X1_LOC_66/A 0.15fF
C44600 OR2X1_LOC_356/B OR2X1_LOC_356/a_36_216# 0.00fF
C44601 OR2X1_LOC_399/a_8_216# OR2X1_LOC_399/Y -0.00fF
C44602 OR2X1_LOC_96/Y OR2X1_LOC_46/A 0.01fF
C44603 AND2X1_LOC_567/a_8_24# AND2X1_LOC_727/A 0.01fF
C44604 OR2X1_LOC_664/Y OR2X1_LOC_161/A 0.03fF
C44605 AND2X1_LOC_364/A OR2X1_LOC_43/A 0.07fF
C44606 OR2X1_LOC_841/A OR2X1_LOC_121/B 0.02fF
C44607 OR2X1_LOC_45/B AND2X1_LOC_648/B 0.03fF
C44608 OR2X1_LOC_823/a_8_216# OR2X1_LOC_6/A 0.01fF
C44609 AND2X1_LOC_374/a_36_24# OR2X1_LOC_26/Y 0.01fF
C44610 OR2X1_LOC_694/Y OR2X1_LOC_22/Y 0.01fF
C44611 AND2X1_LOC_573/A OR2X1_LOC_6/A 0.03fF
C44612 OR2X1_LOC_223/A OR2X1_LOC_161/B 0.06fF
C44613 OR2X1_LOC_857/a_36_216# OR2X1_LOC_35/Y 0.00fF
C44614 OR2X1_LOC_532/B OR2X1_LOC_723/a_8_216# 0.01fF
C44615 AND2X1_LOC_583/a_8_24# AND2X1_LOC_1/Y 0.02fF
C44616 OR2X1_LOC_316/Y OR2X1_LOC_85/A 0.01fF
C44617 OR2X1_LOC_625/a_8_216# OR2X1_LOC_585/A 0.19fF
C44618 OR2X1_LOC_160/A OR2X1_LOC_673/Y 0.01fF
C44619 OR2X1_LOC_158/A OR2X1_LOC_416/A 0.04fF
C44620 OR2X1_LOC_40/Y OR2X1_LOC_417/A 0.27fF
C44621 AND2X1_LOC_840/B OR2X1_LOC_39/A 0.11fF
C44622 AND2X1_LOC_65/a_8_24# OR2X1_LOC_473/Y 0.18fF
C44623 VDD AND2X1_LOC_5/a_8_24# -0.00fF
C44624 AND2X1_LOC_717/a_8_24# AND2X1_LOC_458/a_8_24# 0.23fF
C44625 OR2X1_LOC_643/A OR2X1_LOC_231/a_36_216# 0.02fF
C44626 OR2X1_LOC_698/a_8_216# OR2X1_LOC_64/Y 0.07fF
C44627 AND2X1_LOC_64/Y OR2X1_LOC_675/Y 0.02fF
C44628 OR2X1_LOC_811/A AND2X1_LOC_3/Y 0.06fF
C44629 OR2X1_LOC_83/Y OR2X1_LOC_393/Y 0.00fF
C44630 AND2X1_LOC_456/Y OR2X1_LOC_427/A 0.03fF
C44631 AND2X1_LOC_866/B AND2X1_LOC_631/Y 0.02fF
C44632 OR2X1_LOC_485/Y OR2X1_LOC_31/Y 0.03fF
C44633 OR2X1_LOC_654/A AND2X1_LOC_290/a_8_24# 0.09fF
C44634 OR2X1_LOC_74/a_8_216# OR2X1_LOC_39/A 0.04fF
C44635 OR2X1_LOC_696/A AND2X1_LOC_796/A 0.26fF
C44636 OR2X1_LOC_805/A OR2X1_LOC_269/B 0.17fF
C44637 OR2X1_LOC_427/A OR2X1_LOC_74/A 16.42fF
C44638 OR2X1_LOC_3/Y AND2X1_LOC_398/a_8_24# 0.01fF
C44639 AND2X1_LOC_558/a_8_24# OR2X1_LOC_71/Y 0.00fF
C44640 OR2X1_LOC_585/A AND2X1_LOC_436/B 0.02fF
C44641 AND2X1_LOC_81/B OR2X1_LOC_643/A 0.03fF
C44642 AND2X1_LOC_22/Y OR2X1_LOC_318/B 0.05fF
C44643 AND2X1_LOC_729/a_36_24# OR2X1_LOC_47/Y 0.00fF
C44644 AND2X1_LOC_458/Y AND2X1_LOC_458/a_8_24# 0.00fF
C44645 OR2X1_LOC_114/Y OR2X1_LOC_203/Y 0.00fF
C44646 AND2X1_LOC_713/Y AND2X1_LOC_645/a_8_24# 0.19fF
C44647 OR2X1_LOC_456/Y OR2X1_LOC_465/B 0.04fF
C44648 AND2X1_LOC_481/a_8_24# OR2X1_LOC_375/A 0.04fF
C44649 OR2X1_LOC_679/A AND2X1_LOC_663/A 0.50fF
C44650 OR2X1_LOC_47/Y AND2X1_LOC_778/Y 0.03fF
C44651 OR2X1_LOC_600/A AND2X1_LOC_851/B 0.07fF
C44652 OR2X1_LOC_503/A OR2X1_LOC_7/A 0.00fF
C44653 AND2X1_LOC_303/B OR2X1_LOC_52/B -0.02fF
C44654 AND2X1_LOC_578/A AND2X1_LOC_621/Y 0.07fF
C44655 AND2X1_LOC_557/a_8_24# AND2X1_LOC_573/A 0.03fF
C44656 OR2X1_LOC_427/A OR2X1_LOC_261/A 0.01fF
C44657 VDD AND2X1_LOC_250/a_8_24# 0.00fF
C44658 OR2X1_LOC_175/Y OR2X1_LOC_568/A 0.80fF
C44659 AND2X1_LOC_843/Y OR2X1_LOC_64/Y 0.32fF
C44660 AND2X1_LOC_141/B OR2X1_LOC_118/Y 0.01fF
C44661 OR2X1_LOC_481/A OR2X1_LOC_18/Y 0.02fF
C44662 OR2X1_LOC_151/A AND2X1_LOC_72/B 1.33fF
C44663 OR2X1_LOC_311/Y OR2X1_LOC_761/Y 0.02fF
C44664 OR2X1_LOC_3/Y AND2X1_LOC_379/a_8_24# 0.03fF
C44665 OR2X1_LOC_175/Y OR2X1_LOC_578/B 0.01fF
C44666 AND2X1_LOC_44/Y AND2X1_LOC_609/a_36_24# 0.01fF
C44667 OR2X1_LOC_119/a_8_216# OR2X1_LOC_619/Y 0.03fF
C44668 AND2X1_LOC_81/B OR2X1_LOC_647/A 0.09fF
C44669 OR2X1_LOC_62/A OR2X1_LOC_56/A 0.10fF
C44670 AND2X1_LOC_191/Y OR2X1_LOC_613/Y 0.01fF
C44671 OR2X1_LOC_64/Y AND2X1_LOC_644/Y 0.01fF
C44672 OR2X1_LOC_673/Y AND2X1_LOC_86/B 0.00fF
C44673 OR2X1_LOC_817/a_8_216# OR2X1_LOC_44/Y 0.01fF
C44674 OR2X1_LOC_118/a_8_216# OR2X1_LOC_88/Y 0.01fF
C44675 OR2X1_LOC_223/A OR2X1_LOC_785/a_36_216# 0.00fF
C44676 OR2X1_LOC_805/A OR2X1_LOC_215/A 0.03fF
C44677 OR2X1_LOC_158/A OR2X1_LOC_163/a_8_216# 0.01fF
C44678 OR2X1_LOC_7/A OR2X1_LOC_690/A 0.03fF
C44679 AND2X1_LOC_711/Y OR2X1_LOC_613/Y 0.03fF
C44680 OR2X1_LOC_64/Y OR2X1_LOC_424/a_8_216# 0.01fF
C44681 OR2X1_LOC_3/Y OR2X1_LOC_43/A 0.48fF
C44682 OR2X1_LOC_835/A AND2X1_LOC_51/Y 0.01fF
C44683 AND2X1_LOC_47/Y OR2X1_LOC_623/B 0.01fF
C44684 D_INPUT_5 OR2X1_LOC_409/B 0.00fF
C44685 OR2X1_LOC_740/B OR2X1_LOC_739/a_8_216# 0.02fF
C44686 OR2X1_LOC_252/Y OR2X1_LOC_628/Y 0.02fF
C44687 OR2X1_LOC_275/A OR2X1_LOC_26/Y 0.04fF
C44688 AND2X1_LOC_78/a_8_24# OR2X1_LOC_89/A 0.00fF
C44689 AND2X1_LOC_843/Y OR2X1_LOC_417/A 0.01fF
C44690 OR2X1_LOC_644/a_36_216# OR2X1_LOC_228/Y 0.02fF
C44691 AND2X1_LOC_47/Y OR2X1_LOC_794/A 0.00fF
C44692 OR2X1_LOC_18/Y OR2X1_LOC_71/Y 1.49fF
C44693 OR2X1_LOC_517/A OR2X1_LOC_47/Y 0.02fF
C44694 OR2X1_LOC_754/A OR2X1_LOC_89/A 0.03fF
C44695 OR2X1_LOC_474/Y OR2X1_LOC_786/Y 0.42fF
C44696 AND2X1_LOC_811/Y AND2X1_LOC_804/Y 0.59fF
C44697 OR2X1_LOC_218/a_8_216# OR2X1_LOC_121/B 0.01fF
C44698 OR2X1_LOC_275/A OR2X1_LOC_89/A 0.03fF
C44699 AND2X1_LOC_663/B OR2X1_LOC_757/a_36_216# 0.00fF
C44700 OR2X1_LOC_64/Y OR2X1_LOC_7/A 0.53fF
C44701 OR2X1_LOC_91/Y AND2X1_LOC_845/Y 0.05fF
C44702 D_GATE_741 OR2X1_LOC_192/a_8_216# 0.01fF
C44703 OR2X1_LOC_31/Y OR2X1_LOC_39/A 0.30fF
C44704 OR2X1_LOC_328/a_8_216# OR2X1_LOC_70/A 0.18fF
C44705 AND2X1_LOC_852/B D_INPUT_1 0.05fF
C44706 AND2X1_LOC_662/a_36_24# OR2X1_LOC_74/A 0.01fF
C44707 AND2X1_LOC_849/A AND2X1_LOC_717/B 0.03fF
C44708 AND2X1_LOC_42/B OR2X1_LOC_99/B 0.01fF
C44709 OR2X1_LOC_62/A AND2X1_LOC_9/a_8_24# 0.01fF
C44710 OR2X1_LOC_3/Y AND2X1_LOC_685/a_8_24# 0.01fF
C44711 OR2X1_LOC_320/Y OR2X1_LOC_64/Y 0.29fF
C44712 OR2X1_LOC_78/A OR2X1_LOC_779/B 0.04fF
C44713 OR2X1_LOC_35/Y OR2X1_LOC_68/B 0.03fF
C44714 OR2X1_LOC_56/A OR2X1_LOC_172/Y 0.02fF
C44715 OR2X1_LOC_121/B OR2X1_LOC_794/a_36_216# 0.00fF
C44716 AND2X1_LOC_40/Y AND2X1_LOC_485/a_8_24# 0.03fF
C44717 AND2X1_LOC_648/B AND2X1_LOC_435/a_8_24# 0.01fF
C44718 OR2X1_LOC_18/Y D_INPUT_1 0.67fF
C44719 OR2X1_LOC_857/B OR2X1_LOC_771/B 0.03fF
C44720 OR2X1_LOC_47/Y AND2X1_LOC_624/A 0.03fF
C44721 OR2X1_LOC_116/A OR2X1_LOC_786/Y 0.01fF
C44722 AND2X1_LOC_580/B OR2X1_LOC_95/Y 0.02fF
C44723 OR2X1_LOC_851/B OR2X1_LOC_723/B 0.17fF
C44724 OR2X1_LOC_71/a_8_216# OR2X1_LOC_67/Y 0.01fF
C44725 AND2X1_LOC_59/Y D_INPUT_1 0.03fF
C44726 OR2X1_LOC_604/A OR2X1_LOC_13/B 0.17fF
C44727 OR2X1_LOC_18/Y OR2X1_LOC_173/a_8_216# 0.01fF
C44728 AND2X1_LOC_580/A OR2X1_LOC_615/Y 0.03fF
C44729 OR2X1_LOC_87/A OR2X1_LOC_200/Y 0.01fF
C44730 OR2X1_LOC_417/A OR2X1_LOC_7/A 0.45fF
C44731 OR2X1_LOC_380/A OR2X1_LOC_47/Y 0.02fF
C44732 AND2X1_LOC_211/B OR2X1_LOC_31/Y 0.03fF
C44733 OR2X1_LOC_217/Y OR2X1_LOC_786/Y 0.23fF
C44734 D_INPUT_3 OR2X1_LOC_753/A 0.07fF
C44735 OR2X1_LOC_158/A OR2X1_LOC_268/Y 0.03fF
C44736 OR2X1_LOC_151/A AND2X1_LOC_36/Y 0.12fF
C44737 AND2X1_LOC_524/a_36_24# AND2X1_LOC_36/Y 0.01fF
C44738 AND2X1_LOC_43/a_8_24# AND2X1_LOC_47/Y 0.01fF
C44739 AND2X1_LOC_8/Y OR2X1_LOC_62/A 1.05fF
C44740 OR2X1_LOC_158/A OR2X1_LOC_183/Y 0.04fF
C44741 VDD OR2X1_LOC_349/B 0.06fF
C44742 OR2X1_LOC_865/a_8_216# D_INPUT_1 0.01fF
C44743 OR2X1_LOC_448/B OR2X1_LOC_779/B 0.02fF
C44744 INPUT_1 OR2X1_LOC_8/a_8_216# 0.01fF
C44745 OR2X1_LOC_429/Y OR2X1_LOC_31/Y 0.02fF
C44746 AND2X1_LOC_856/a_8_24# OR2X1_LOC_46/A 0.17fF
C44747 INPUT_4 AND2X1_LOC_451/a_36_24# 0.00fF
C44748 OR2X1_LOC_63/a_8_216# AND2X1_LOC_647/Y 0.01fF
C44749 OR2X1_LOC_45/B AND2X1_LOC_465/A 0.03fF
C44750 OR2X1_LOC_485/A AND2X1_LOC_810/Y 0.20fF
C44751 AND2X1_LOC_196/Y AND2X1_LOC_729/B 0.00fF
C44752 AND2X1_LOC_59/Y OR2X1_LOC_356/a_36_216# 0.00fF
C44753 OR2X1_LOC_185/A OR2X1_LOC_543/a_8_216# 0.00fF
C44754 OR2X1_LOC_89/A OR2X1_LOC_55/a_36_216# 0.00fF
C44755 AND2X1_LOC_64/Y OR2X1_LOC_736/Y 0.03fF
C44756 OR2X1_LOC_427/A AND2X1_LOC_783/a_8_24# 0.01fF
C44757 OR2X1_LOC_45/B AND2X1_LOC_231/a_8_24# 0.06fF
C44758 AND2X1_LOC_825/a_8_24# OR2X1_LOC_46/A 0.02fF
C44759 OR2X1_LOC_186/Y AND2X1_LOC_91/B 0.03fF
C44760 OR2X1_LOC_485/A OR2X1_LOC_760/Y 0.01fF
C44761 AND2X1_LOC_786/a_8_24# OR2X1_LOC_79/Y 0.01fF
C44762 OR2X1_LOC_19/B OR2X1_LOC_243/a_8_216# 0.01fF
C44763 OR2X1_LOC_62/A OR2X1_LOC_291/A 0.00fF
C44764 OR2X1_LOC_538/A OR2X1_LOC_788/B 0.02fF
C44765 OR2X1_LOC_494/a_8_216# OR2X1_LOC_437/A 0.03fF
C44766 OR2X1_LOC_840/A OR2X1_LOC_728/A 0.40fF
C44767 OR2X1_LOC_99/A OR2X1_LOC_99/a_8_216# 0.04fF
C44768 OR2X1_LOC_375/A OR2X1_LOC_512/Y 0.01fF
C44769 OR2X1_LOC_185/A OR2X1_LOC_348/B 0.01fF
C44770 OR2X1_LOC_134/a_36_216# AND2X1_LOC_541/Y 0.00fF
C44771 OR2X1_LOC_70/A OR2X1_LOC_752/a_8_216# 0.00fF
C44772 OR2X1_LOC_49/A OR2X1_LOC_633/A 0.27fF
C44773 OR2X1_LOC_32/B OR2X1_LOC_80/A 1.04fF
C44774 OR2X1_LOC_585/A OR2X1_LOC_598/A 0.02fF
C44775 AND2X1_LOC_539/Y OR2X1_LOC_329/Y 0.02fF
C44776 OR2X1_LOC_85/A OR2X1_LOC_153/a_8_216# 0.08fF
C44777 AND2X1_LOC_544/Y OR2X1_LOC_40/Y 16.19fF
C44778 OR2X1_LOC_351/B AND2X1_LOC_22/Y 0.68fF
C44779 AND2X1_LOC_41/A OR2X1_LOC_308/Y 0.13fF
C44780 AND2X1_LOC_64/Y OR2X1_LOC_641/Y 0.08fF
C44781 OR2X1_LOC_134/Y VDD 0.11fF
C44782 AND2X1_LOC_821/a_8_24# OR2X1_LOC_532/B 0.01fF
C44783 OR2X1_LOC_494/A AND2X1_LOC_860/A 0.03fF
C44784 AND2X1_LOC_850/a_8_24# OR2X1_LOC_13/B 0.01fF
C44785 OR2X1_LOC_624/A OR2X1_LOC_140/Y 0.05fF
C44786 OR2X1_LOC_506/Y OR2X1_LOC_151/A 0.01fF
C44787 AND2X1_LOC_47/Y OR2X1_LOC_544/A 0.01fF
C44788 OR2X1_LOC_114/B AND2X1_LOC_22/Y 0.05fF
C44789 OR2X1_LOC_155/A OR2X1_LOC_779/B 0.03fF
C44790 OR2X1_LOC_161/A OR2X1_LOC_342/a_8_216# 0.01fF
C44791 AND2X1_LOC_566/B OR2X1_LOC_12/Y 0.03fF
C44792 AND2X1_LOC_706/Y AND2X1_LOC_714/B 0.19fF
C44793 D_INPUT_3 AND2X1_LOC_845/Y 0.07fF
C44794 OR2X1_LOC_31/Y OR2X1_LOC_428/a_8_216# 0.07fF
C44795 OR2X1_LOC_527/a_36_216# AND2X1_LOC_786/Y 0.01fF
C44796 AND2X1_LOC_172/a_8_24# AND2X1_LOC_7/B 0.01fF
C44797 AND2X1_LOC_535/Y AND2X1_LOC_802/Y 0.03fF
C44798 OR2X1_LOC_784/B AND2X1_LOC_44/Y 0.11fF
C44799 OR2X1_LOC_97/A VDD 0.51fF
C44800 OR2X1_LOC_44/Y OR2X1_LOC_384/Y 0.03fF
C44801 OR2X1_LOC_306/Y OR2X1_LOC_13/B 0.05fF
C44802 AND2X1_LOC_582/a_8_24# AND2X1_LOC_582/B 0.01fF
C44803 AND2X1_LOC_91/a_8_24# AND2X1_LOC_70/Y 0.02fF
C44804 OR2X1_LOC_410/a_8_216# OR2X1_LOC_334/a_8_216# 0.47fF
C44805 OR2X1_LOC_487/a_36_216# AND2X1_LOC_563/Y 0.00fF
C44806 OR2X1_LOC_857/A OR2X1_LOC_66/A 0.29fF
C44807 AND2X1_LOC_262/a_8_24# OR2X1_LOC_549/A 0.02fF
C44808 OR2X1_LOC_56/A OR2X1_LOC_312/a_36_216# 0.03fF
C44809 AND2X1_LOC_432/a_36_24# AND2X1_LOC_70/Y 0.00fF
C44810 AND2X1_LOC_756/a_36_24# GATE_579 0.00fF
C44811 AND2X1_LOC_64/Y OR2X1_LOC_808/B 0.03fF
C44812 AND2X1_LOC_806/A OR2X1_LOC_437/A 0.03fF
C44813 OR2X1_LOC_3/Y OR2X1_LOC_384/a_8_216# 0.01fF
C44814 VDD AND2X1_LOC_339/B 0.39fF
C44815 OR2X1_LOC_202/a_8_216# AND2X1_LOC_31/Y 0.01fF
C44816 OR2X1_LOC_154/A OR2X1_LOC_174/Y 0.03fF
C44817 OR2X1_LOC_744/A OR2X1_LOC_744/Y 0.01fF
C44818 VDD D_GATE_662 0.24fF
C44819 AND2X1_LOC_91/B OR2X1_LOC_862/A 0.03fF
C44820 VDD OR2X1_LOC_482/a_8_216# 0.00fF
C44821 OR2X1_LOC_59/Y AND2X1_LOC_786/Y 0.17fF
C44822 AND2X1_LOC_59/Y OR2X1_LOC_180/B 0.29fF
C44823 OR2X1_LOC_532/B OR2X1_LOC_330/a_36_216# 0.00fF
C44824 OR2X1_LOC_121/B OR2X1_LOC_559/a_8_216# 0.01fF
C44825 D_INPUT_0 OR2X1_LOC_512/a_8_216# 0.02fF
C44826 OR2X1_LOC_87/A AND2X1_LOC_591/a_8_24# 0.04fF
C44827 OR2X1_LOC_532/B OR2X1_LOC_737/a_8_216# 0.01fF
C44828 OR2X1_LOC_175/Y OR2X1_LOC_798/Y 0.10fF
C44829 AND2X1_LOC_95/Y OR2X1_LOC_356/B 0.13fF
C44830 OR2X1_LOC_709/A OR2X1_LOC_78/A 0.07fF
C44831 AND2X1_LOC_788/a_36_24# OR2X1_LOC_51/Y 0.00fF
C44832 AND2X1_LOC_295/a_8_24# OR2X1_LOC_78/A 0.05fF
C44833 OR2X1_LOC_139/A OR2X1_LOC_216/A 0.52fF
C44834 OR2X1_LOC_26/Y OR2X1_LOC_142/Y 0.18fF
C44835 OR2X1_LOC_416/Y OR2X1_LOC_68/B 0.02fF
C44836 OR2X1_LOC_715/B OR2X1_LOC_785/a_8_216# 0.30fF
C44837 AND2X1_LOC_303/a_8_24# OR2X1_LOC_16/A 0.03fF
C44838 OR2X1_LOC_7/A AND2X1_LOC_247/a_8_24# 0.03fF
C44839 OR2X1_LOC_121/Y OR2X1_LOC_244/B 0.02fF
C44840 AND2X1_LOC_152/a_8_24# OR2X1_LOC_209/A 0.01fF
C44841 AND2X1_LOC_3/Y OR2X1_LOC_777/B 0.03fF
C44842 AND2X1_LOC_357/A OR2X1_LOC_426/B 0.04fF
C44843 OR2X1_LOC_151/A OR2X1_LOC_630/Y 0.38fF
C44844 OR2X1_LOC_176/Y AND2X1_LOC_716/Y 0.05fF
C44845 OR2X1_LOC_502/A OR2X1_LOC_161/B 0.23fF
C44846 OR2X1_LOC_89/A OR2X1_LOC_142/Y 0.08fF
C44847 AND2X1_LOC_287/B OR2X1_LOC_278/Y 0.15fF
C44848 OR2X1_LOC_78/B OR2X1_LOC_641/A 0.07fF
C44849 AND2X1_LOC_662/B AND2X1_LOC_473/Y 0.20fF
C44850 OR2X1_LOC_464/A OR2X1_LOC_736/Y 0.12fF
C44851 OR2X1_LOC_302/B OR2X1_LOC_302/A 0.01fF
C44852 OR2X1_LOC_570/a_8_216# OR2X1_LOC_562/A 0.01fF
C44853 AND2X1_LOC_91/B OR2X1_LOC_773/B 0.03fF
C44854 OR2X1_LOC_302/B VDD 0.21fF
C44855 OR2X1_LOC_8/Y OR2X1_LOC_56/A 0.24fF
C44856 AND2X1_LOC_84/Y OR2X1_LOC_265/Y 0.05fF
C44857 OR2X1_LOC_787/Y OR2X1_LOC_301/a_8_216# 0.07fF
C44858 AND2X1_LOC_436/Y AND2X1_LOC_469/B 0.00fF
C44859 AND2X1_LOC_714/a_8_24# OR2X1_LOC_48/B 0.03fF
C44860 AND2X1_LOC_12/Y AND2X1_LOC_22/Y 0.34fF
C44861 AND2X1_LOC_364/Y AND2X1_LOC_335/Y 0.00fF
C44862 AND2X1_LOC_70/Y OR2X1_LOC_78/A 1.29fF
C44863 AND2X1_LOC_553/A OR2X1_LOC_158/A 0.01fF
C44864 OR2X1_LOC_134/a_8_216# OR2X1_LOC_26/Y 0.01fF
C44865 AND2X1_LOC_56/B OR2X1_LOC_397/Y 0.03fF
C44866 AND2X1_LOC_392/A AND2X1_LOC_365/a_36_24# 0.01fF
C44867 OR2X1_LOC_177/a_8_216# AND2X1_LOC_550/A 0.01fF
C44868 OR2X1_LOC_59/Y AND2X1_LOC_218/Y 0.01fF
C44869 OR2X1_LOC_45/B OR2X1_LOC_237/Y 0.33fF
C44870 OR2X1_LOC_186/Y OR2X1_LOC_799/A 0.00fF
C44871 OR2X1_LOC_401/B OR2X1_LOC_771/B 0.03fF
C44872 OR2X1_LOC_92/Y AND2X1_LOC_243/Y 0.74fF
C44873 AND2X1_LOC_213/B OR2X1_LOC_39/A 0.03fF
C44874 OR2X1_LOC_858/A OR2X1_LOC_632/Y 0.23fF
C44875 OR2X1_LOC_778/B OR2X1_LOC_778/a_8_216# 0.03fF
C44876 OR2X1_LOC_624/A OR2X1_LOC_390/A 0.03fF
C44877 OR2X1_LOC_458/B AND2X1_LOC_70/Y 0.03fF
C44878 OR2X1_LOC_185/A AND2X1_LOC_65/A 0.09fF
C44879 AND2X1_LOC_802/B AND2X1_LOC_661/A 0.62fF
C44880 AND2X1_LOC_352/a_8_24# AND2X1_LOC_654/Y 0.04fF
C44881 AND2X1_LOC_212/A AND2X1_LOC_662/B 0.01fF
C44882 OR2X1_LOC_744/A AND2X1_LOC_474/A 0.06fF
C44883 OR2X1_LOC_161/A OR2X1_LOC_162/a_8_216# 0.00fF
C44884 OR2X1_LOC_326/a_8_216# OR2X1_LOC_538/A 0.01fF
C44885 AND2X1_LOC_22/Y OR2X1_LOC_841/B 0.05fF
C44886 OR2X1_LOC_673/Y OR2X1_LOC_266/A 0.02fF
C44887 AND2X1_LOC_220/Y AND2X1_LOC_220/B 0.15fF
C44888 VDD OR2X1_LOC_475/B 0.09fF
C44889 OR2X1_LOC_841/a_8_216# OR2X1_LOC_841/A 0.02fF
C44890 OR2X1_LOC_36/Y OR2X1_LOC_428/A 0.23fF
C44891 OR2X1_LOC_703/A OR2X1_LOC_78/A 0.03fF
C44892 OR2X1_LOC_137/a_8_216# OR2X1_LOC_235/B 0.01fF
C44893 OR2X1_LOC_6/B OR2X1_LOC_833/B 0.47fF
C44894 AND2X1_LOC_95/Y OR2X1_LOC_182/B 0.03fF
C44895 OR2X1_LOC_467/B OR2X1_LOC_467/a_8_216# 0.01fF
C44896 OR2X1_LOC_427/A AND2X1_LOC_860/A 0.21fF
C44897 OR2X1_LOC_329/B OR2X1_LOC_275/Y 0.08fF
C44898 AND2X1_LOC_17/a_8_24# INPUT_7 0.11fF
C44899 OR2X1_LOC_671/Y OR2X1_LOC_94/a_8_216# 0.04fF
C44900 OR2X1_LOC_147/B OR2X1_LOC_741/Y 0.03fF
C44901 OR2X1_LOC_40/Y AND2X1_LOC_550/A 0.16fF
C44902 OR2X1_LOC_856/B OR2X1_LOC_66/A 0.21fF
C44903 OR2X1_LOC_770/A AND2X1_LOC_3/Y 0.01fF
C44904 AND2X1_LOC_81/a_8_24# AND2X1_LOC_44/Y 0.01fF
C44905 AND2X1_LOC_854/a_36_24# OR2X1_LOC_428/A 0.01fF
C44906 OR2X1_LOC_269/B OR2X1_LOC_580/B 3.87fF
C44907 OR2X1_LOC_65/B AND2X1_LOC_243/Y 0.00fF
C44908 OR2X1_LOC_137/Y OR2X1_LOC_161/B 0.00fF
C44909 INPUT_1 AND2X1_LOC_36/Y 0.12fF
C44910 OR2X1_LOC_426/B OR2X1_LOC_48/B 0.24fF
C44911 OR2X1_LOC_529/Y OR2X1_LOC_530/a_8_216# 0.00fF
C44912 OR2X1_LOC_375/A OR2X1_LOC_641/A 0.03fF
C44913 OR2X1_LOC_39/Y AND2X1_LOC_194/a_8_24# 0.01fF
C44914 OR2X1_LOC_45/B OR2X1_LOC_487/a_8_216# 0.07fF
C44915 OR2X1_LOC_329/B OR2X1_LOC_495/Y 0.03fF
C44916 OR2X1_LOC_47/Y OR2X1_LOC_150/a_8_216# 0.01fF
C44917 AND2X1_LOC_76/Y OR2X1_LOC_56/A 0.03fF
C44918 OR2X1_LOC_632/a_8_216# OR2X1_LOC_575/A 0.00fF
C44919 AND2X1_LOC_95/Y AND2X1_LOC_184/a_36_24# 0.01fF
C44920 OR2X1_LOC_49/A OR2X1_LOC_827/Y 0.81fF
C44921 INPUT_0 OR2X1_LOC_637/a_8_216# 0.05fF
C44922 AND2X1_LOC_43/B AND2X1_LOC_18/Y 0.10fF
C44923 AND2X1_LOC_72/a_8_24# OR2X1_LOC_161/B 0.01fF
C44924 OR2X1_LOC_426/B OR2X1_LOC_18/Y 0.20fF
C44925 OR2X1_LOC_709/A OR2X1_LOC_155/A 0.48fF
C44926 AND2X1_LOC_22/Y OR2X1_LOC_804/B 0.12fF
C44927 OR2X1_LOC_8/Y AND2X1_LOC_9/a_8_24# 0.00fF
C44928 OR2X1_LOC_312/Y AND2X1_LOC_212/Y 0.15fF
C44929 OR2X1_LOC_856/B AND2X1_LOC_311/a_8_24# 0.02fF
C44930 VDD AND2X1_LOC_633/a_8_24# -0.00fF
C44931 AND2X1_LOC_560/a_8_24# OR2X1_LOC_22/Y 0.01fF
C44932 OR2X1_LOC_502/A AND2X1_LOC_48/a_8_24# 0.01fF
C44933 AND2X1_LOC_706/Y AND2X1_LOC_645/A 0.03fF
C44934 AND2X1_LOC_56/B OR2X1_LOC_629/B 0.01fF
C44935 OR2X1_LOC_151/A OR2X1_LOC_346/B 0.01fF
C44936 VDD AND2X1_LOC_282/a_8_24# 0.00fF
C44937 OR2X1_LOC_235/B OR2X1_LOC_291/a_8_216# 0.01fF
C44938 AND2X1_LOC_553/A OR2X1_LOC_103/Y 0.02fF
C44939 OR2X1_LOC_648/B OR2X1_LOC_269/B 0.12fF
C44940 OR2X1_LOC_744/A AND2X1_LOC_593/Y 0.53fF
C44941 AND2X1_LOC_70/Y OR2X1_LOC_602/A 0.01fF
C44942 OR2X1_LOC_67/A OR2X1_LOC_56/A 1.34fF
C44943 OR2X1_LOC_685/A OR2X1_LOC_687/A 0.15fF
C44944 OR2X1_LOC_70/Y AND2X1_LOC_786/Y 0.21fF
C44945 AND2X1_LOC_364/Y OR2X1_LOC_619/Y 0.02fF
C44946 AND2X1_LOC_61/a_8_24# OR2X1_LOC_85/A 0.01fF
C44947 VDD OR2X1_LOC_699/a_8_216# 0.21fF
C44948 OR2X1_LOC_461/a_36_216# AND2X1_LOC_824/B 0.02fF
C44949 OR2X1_LOC_532/B OR2X1_LOC_605/Y 0.15fF
C44950 OR2X1_LOC_600/A OR2X1_LOC_372/Y 0.06fF
C44951 AND2X1_LOC_212/A AND2X1_LOC_337/B 0.00fF
C44952 OR2X1_LOC_45/B AND2X1_LOC_853/a_36_24# 0.00fF
C44953 OR2X1_LOC_502/A OR2X1_LOC_61/Y 4.88fF
C44954 AND2X1_LOC_547/Y AND2X1_LOC_564/a_36_24# 0.01fF
C44955 OR2X1_LOC_96/Y OR2X1_LOC_93/a_8_216# 0.01fF
C44956 AND2X1_LOC_363/A AND2X1_LOC_860/A 0.03fF
C44957 OR2X1_LOC_251/a_8_216# OR2X1_LOC_278/Y 0.01fF
C44958 AND2X1_LOC_367/B AND2X1_LOC_367/a_8_24# 0.05fF
C44959 OR2X1_LOC_625/Y OR2X1_LOC_517/A 0.01fF
C44960 AND2X1_LOC_280/a_8_24# OR2X1_LOC_366/Y 0.05fF
C44961 AND2X1_LOC_72/a_36_24# OR2X1_LOC_719/B 0.01fF
C44962 OR2X1_LOC_854/a_8_216# OR2X1_LOC_620/Y -0.03fF
C44963 OR2X1_LOC_158/A AND2X1_LOC_345/Y 0.03fF
C44964 OR2X1_LOC_728/B OR2X1_LOC_446/B 0.03fF
C44965 OR2X1_LOC_715/a_8_216# OR2X1_LOC_724/A 0.03fF
C44966 OR2X1_LOC_686/A AND2X1_LOC_3/Y 0.03fF
C44967 AND2X1_LOC_67/a_36_24# OR2X1_LOC_506/A 0.00fF
C44968 OR2X1_LOC_659/Y AND2X1_LOC_51/Y 0.00fF
C44969 AND2X1_LOC_12/Y OR2X1_LOC_706/A 0.06fF
C44970 OR2X1_LOC_744/A OR2X1_LOC_85/A 0.02fF
C44971 OR2X1_LOC_68/B OR2X1_LOC_80/A 1.66fF
C44972 AND2X1_LOC_547/Y OR2X1_LOC_189/Y 0.03fF
C44973 OR2X1_LOC_194/Y OR2X1_LOC_78/B 0.02fF
C44974 OR2X1_LOC_850/B OR2X1_LOC_362/B 0.02fF
C44975 OR2X1_LOC_687/Y OR2X1_LOC_678/a_8_216# 0.03fF
C44976 AND2X1_LOC_219/a_36_24# OR2X1_LOC_26/Y 0.00fF
C44977 OR2X1_LOC_56/A AND2X1_LOC_374/Y 0.02fF
C44978 OR2X1_LOC_599/A AND2X1_LOC_663/A 0.05fF
C44979 OR2X1_LOC_448/A OR2X1_LOC_161/A 0.01fF
C44980 OR2X1_LOC_134/Y OR2X1_LOC_256/A 0.00fF
C44981 AND2X1_LOC_858/B OR2X1_LOC_44/Y 0.00fF
C44982 AND2X1_LOC_70/Y OR2X1_LOC_155/A 0.29fF
C44983 OR2X1_LOC_334/B AND2X1_LOC_291/a_8_24# 0.01fF
C44984 OR2X1_LOC_634/a_8_216# AND2X1_LOC_824/B 0.01fF
C44985 AND2X1_LOC_738/B OR2X1_LOC_52/B 0.07fF
C44986 AND2X1_LOC_40/Y OR2X1_LOC_456/a_8_216# 0.02fF
C44987 OR2X1_LOC_426/A AND2X1_LOC_452/Y 0.54fF
C44988 AND2X1_LOC_858/B AND2X1_LOC_288/a_8_24# 0.03fF
C44989 OR2X1_LOC_91/A OR2X1_LOC_44/Y 1.34fF
C44990 OR2X1_LOC_728/B OR2X1_LOC_728/a_8_216# 0.01fF
C44991 AND2X1_LOC_331/a_8_24# OR2X1_LOC_739/A 0.01fF
C44992 AND2X1_LOC_804/a_8_24# OR2X1_LOC_142/Y 0.02fF
C44993 OR2X1_LOC_56/A OR2X1_LOC_52/B 9.09fF
C44994 OR2X1_LOC_405/A OR2X1_LOC_734/a_36_216# 0.01fF
C44995 AND2X1_LOC_48/A OR2X1_LOC_161/B 0.07fF
C44996 OR2X1_LOC_329/B OR2X1_LOC_43/A 0.03fF
C44997 OR2X1_LOC_672/Y OR2X1_LOC_56/A 0.01fF
C44998 OR2X1_LOC_385/Y OR2X1_LOC_426/B 0.07fF
C44999 OR2X1_LOC_723/B OR2X1_LOC_717/a_8_216# 0.01fF
C45000 OR2X1_LOC_475/a_8_216# OR2X1_LOC_805/A 0.03fF
C45001 AND2X1_LOC_394/a_8_24# AND2X1_LOC_40/Y 0.03fF
C45002 OR2X1_LOC_61/Y AND2X1_LOC_230/a_8_24# 0.05fF
C45003 OR2X1_LOC_22/Y OR2X1_LOC_522/Y 0.03fF
C45004 AND2X1_LOC_715/A AND2X1_LOC_276/Y 0.04fF
C45005 OR2X1_LOC_494/a_8_216# AND2X1_LOC_348/Y 0.03fF
C45006 OR2X1_LOC_318/Y OR2X1_LOC_539/Y 0.03fF
C45007 AND2X1_LOC_353/a_8_24# OR2X1_LOC_64/Y 0.01fF
C45008 VDD OR2X1_LOC_605/a_8_216# 0.21fF
C45009 OR2X1_LOC_185/A OR2X1_LOC_181/B 0.04fF
C45010 OR2X1_LOC_8/Y OR2X1_LOC_291/A 0.36fF
C45011 OR2X1_LOC_89/A OR2X1_LOC_442/Y 0.11fF
C45012 OR2X1_LOC_3/Y OR2X1_LOC_585/Y 0.10fF
C45013 AND2X1_LOC_547/Y OR2X1_LOC_527/Y 0.00fF
C45014 OR2X1_LOC_804/a_8_216# OR2X1_LOC_778/Y 0.28fF
C45015 AND2X1_LOC_59/Y OR2X1_LOC_737/A 0.17fF
C45016 AND2X1_LOC_802/B AND2X1_LOC_810/Y 0.83fF
C45017 AND2X1_LOC_70/Y OR2X1_LOC_605/A 0.07fF
C45018 AND2X1_LOC_42/B AND2X1_LOC_245/a_8_24# 0.02fF
C45019 OR2X1_LOC_494/a_8_216# OR2X1_LOC_753/A 0.01fF
C45020 AND2X1_LOC_340/Y OR2X1_LOC_71/Y 0.46fF
C45021 OR2X1_LOC_822/a_8_216# OR2X1_LOC_64/Y 0.18fF
C45022 AND2X1_LOC_2/Y AND2X1_LOC_425/a_8_24# 0.01fF
C45023 OR2X1_LOC_114/Y OR2X1_LOC_721/Y 0.05fF
C45024 OR2X1_LOC_625/Y AND2X1_LOC_624/A 0.03fF
C45025 OR2X1_LOC_316/Y AND2X1_LOC_642/a_8_24# 0.01fF
C45026 AND2X1_LOC_746/a_8_24# OR2X1_LOC_220/A 0.23fF
C45027 AND2X1_LOC_753/a_8_24# OR2X1_LOC_375/A 0.02fF
C45028 OR2X1_LOC_665/Y AND2X1_LOC_861/B 0.01fF
C45029 AND2X1_LOC_342/a_8_24# OR2X1_LOC_92/Y 0.01fF
C45030 AND2X1_LOC_59/Y AND2X1_LOC_95/Y 0.85fF
C45031 AND2X1_LOC_573/A AND2X1_LOC_403/B 0.09fF
C45032 AND2X1_LOC_191/Y OR2X1_LOC_524/Y 0.07fF
C45033 AND2X1_LOC_578/A OR2X1_LOC_59/Y 0.07fF
C45034 OR2X1_LOC_377/A AND2X1_LOC_617/a_8_24# 0.03fF
C45035 OR2X1_LOC_91/A AND2X1_LOC_116/Y 0.03fF
C45036 AND2X1_LOC_59/Y OR2X1_LOC_633/Y 0.00fF
C45037 OR2X1_LOC_423/Y AND2X1_LOC_592/a_8_24# 0.03fF
C45038 OR2X1_LOC_206/a_8_216# OR2X1_LOC_78/A 0.05fF
C45039 OR2X1_LOC_427/A AND2X1_LOC_287/Y 0.36fF
C45040 OR2X1_LOC_472/B OR2X1_LOC_461/B 0.01fF
C45041 AND2X1_LOC_12/Y AND2X1_LOC_153/a_8_24# 0.01fF
C45042 AND2X1_LOC_711/Y OR2X1_LOC_524/Y 0.07fF
C45043 AND2X1_LOC_453/a_8_24# AND2X1_LOC_453/Y 0.02fF
C45044 OR2X1_LOC_532/B OR2X1_LOC_361/a_8_216# 0.01fF
C45045 AND2X1_LOC_449/Y AND2X1_LOC_454/Y 0.20fF
C45046 OR2X1_LOC_805/A OR2X1_LOC_539/Y 0.03fF
C45047 OR2X1_LOC_524/Y OR2X1_LOC_70/Y 0.02fF
C45048 OR2X1_LOC_404/Y OR2X1_LOC_78/A 0.04fF
C45049 AND2X1_LOC_24/a_8_24# AND2X1_LOC_51/Y 0.01fF
C45050 OR2X1_LOC_516/A OR2X1_LOC_516/a_8_216# 0.01fF
C45051 OR2X1_LOC_450/B AND2X1_LOC_425/Y 0.01fF
C45052 OR2X1_LOC_203/Y OR2X1_LOC_541/B 0.01fF
C45053 AND2X1_LOC_91/B AND2X1_LOC_225/a_36_24# 0.00fF
C45054 AND2X1_LOC_573/A OR2X1_LOC_44/Y 0.10fF
C45055 OR2X1_LOC_276/A OR2X1_LOC_549/A 0.03fF
C45056 AND2X1_LOC_3/Y OR2X1_LOC_575/A 0.01fF
C45057 OR2X1_LOC_479/Y OR2X1_LOC_840/A 0.10fF
C45058 AND2X1_LOC_43/B AND2X1_LOC_413/a_8_24# 0.05fF
C45059 OR2X1_LOC_194/Y OR2X1_LOC_375/A 0.06fF
C45060 OR2X1_LOC_26/Y OR2X1_LOC_118/Y 0.03fF
C45061 OR2X1_LOC_387/Y OR2X1_LOC_586/Y 0.02fF
C45062 AND2X1_LOC_561/a_8_24# AND2X1_LOC_657/A 0.01fF
C45063 AND2X1_LOC_342/Y AND2X1_LOC_349/a_8_24# 0.07fF
C45064 OR2X1_LOC_377/A OR2X1_LOC_849/A 0.00fF
C45065 OR2X1_LOC_270/Y OR2X1_LOC_344/A 1.08fF
C45066 OR2X1_LOC_864/A OR2X1_LOC_137/B 0.13fF
C45067 AND2X1_LOC_59/Y OR2X1_LOC_99/Y 0.05fF
C45068 OR2X1_LOC_158/A AND2X1_LOC_648/B 0.03fF
C45069 AND2X1_LOC_539/a_8_24# AND2X1_LOC_434/Y 0.02fF
C45070 OR2X1_LOC_743/A OR2X1_LOC_48/B 0.11fF
C45071 AND2X1_LOC_41/A OR2X1_LOC_19/B 0.46fF
C45072 OR2X1_LOC_91/Y AND2X1_LOC_784/A 0.84fF
C45073 AND2X1_LOC_715/A AND2X1_LOC_831/Y 0.00fF
C45074 OR2X1_LOC_89/A OR2X1_LOC_118/Y 0.00fF
C45075 AND2X1_LOC_40/Y OR2X1_LOC_647/Y 0.01fF
C45076 AND2X1_LOC_12/Y OR2X1_LOC_296/a_8_216# 0.03fF
C45077 OR2X1_LOC_743/A OR2X1_LOC_18/Y 0.14fF
C45078 OR2X1_LOC_115/B OR2X1_LOC_68/B 0.02fF
C45079 AND2X1_LOC_717/a_36_24# OR2X1_LOC_280/Y 0.01fF
C45080 OR2X1_LOC_74/a_8_216# OR2X1_LOC_85/A 0.01fF
C45081 AND2X1_LOC_87/a_8_24# OR2X1_LOC_52/B 0.11fF
C45082 OR2X1_LOC_235/B OR2X1_LOC_814/A 0.03fF
C45083 AND2X1_LOC_729/Y OR2X1_LOC_189/Y 0.03fF
C45084 OR2X1_LOC_185/A OR2X1_LOC_204/a_8_216# 0.03fF
C45085 OR2X1_LOC_251/Y AND2X1_LOC_859/a_8_24# -0.00fF
C45086 AND2X1_LOC_36/Y OR2X1_LOC_714/A 0.01fF
C45087 AND2X1_LOC_6/a_36_24# OR2X1_LOC_549/A 0.00fF
C45088 OR2X1_LOC_287/A OR2X1_LOC_288/A 0.10fF
C45089 OR2X1_LOC_106/Y AND2X1_LOC_657/A 0.03fF
C45090 AND2X1_LOC_48/A AND2X1_LOC_48/a_8_24# 0.01fF
C45091 OR2X1_LOC_446/a_8_216# OR2X1_LOC_161/A 0.07fF
C45092 OR2X1_LOC_16/A AND2X1_LOC_228/a_8_24# 0.01fF
C45093 AND2X1_LOC_729/Y OR2X1_LOC_152/Y 0.32fF
C45094 AND2X1_LOC_548/a_8_24# AND2X1_LOC_624/A 0.03fF
C45095 OR2X1_LOC_831/A OR2X1_LOC_804/A 0.02fF
C45096 AND2X1_LOC_44/Y OR2X1_LOC_398/Y 0.33fF
C45097 OR2X1_LOC_83/A OR2X1_LOC_753/A 0.05fF
C45098 OR2X1_LOC_262/Y OR2X1_LOC_26/Y 0.18fF
C45099 OR2X1_LOC_141/B OR2X1_LOC_659/B 0.01fF
C45100 AND2X1_LOC_803/B OR2X1_LOC_47/Y 0.03fF
C45101 AND2X1_LOC_866/A AND2X1_LOC_663/A 0.05fF
C45102 OR2X1_LOC_154/A AND2X1_LOC_42/B 0.38fF
C45103 OR2X1_LOC_84/B AND2X1_LOC_8/Y 0.22fF
C45104 OR2X1_LOC_700/Y AND2X1_LOC_663/B 0.10fF
C45105 OR2X1_LOC_837/B AND2X1_LOC_462/a_8_24# 0.07fF
C45106 OR2X1_LOC_648/A AND2X1_LOC_109/a_8_24# 0.01fF
C45107 AND2X1_LOC_48/A OR2X1_LOC_61/Y 0.04fF
C45108 AND2X1_LOC_126/a_8_24# OR2X1_LOC_244/A -0.01fF
C45109 OR2X1_LOC_538/a_8_216# OR2X1_LOC_532/B 0.01fF
C45110 OR2X1_LOC_32/a_8_216# OR2X1_LOC_690/A 0.40fF
C45111 OR2X1_LOC_405/A AND2X1_LOC_491/a_8_24# 0.01fF
C45112 OR2X1_LOC_719/Y OR2X1_LOC_733/B 0.00fF
C45113 AND2X1_LOC_101/B OR2X1_LOC_7/A 0.73fF
C45114 OR2X1_LOC_401/B OR2X1_LOC_402/Y 0.03fF
C45115 AND2X1_LOC_601/a_8_24# AND2X1_LOC_51/Y 0.02fF
C45116 AND2X1_LOC_114/Y OR2X1_LOC_59/Y 0.02fF
C45117 OR2X1_LOC_855/a_8_216# OR2X1_LOC_198/A 0.14fF
C45118 OR2X1_LOC_154/A OR2X1_LOC_705/Y 0.03fF
C45119 AND2X1_LOC_810/a_36_24# AND2X1_LOC_436/Y 0.00fF
C45120 OR2X1_LOC_70/a_8_216# OR2X1_LOC_426/A 0.01fF
C45121 AND2X1_LOC_42/B OR2X1_LOC_267/A 0.07fF
C45122 AND2X1_LOC_729/Y OR2X1_LOC_417/Y 0.07fF
C45123 OR2X1_LOC_328/a_8_216# OR2X1_LOC_47/Y 0.00fF
C45124 OR2X1_LOC_18/Y OR2X1_LOC_246/A 0.13fF
C45125 OR2X1_LOC_89/A OR2X1_LOC_238/Y 0.03fF
C45126 OR2X1_LOC_140/A OR2X1_LOC_598/A 0.00fF
C45127 OR2X1_LOC_325/B OR2X1_LOC_365/B 0.03fF
C45128 OR2X1_LOC_485/A AND2X1_LOC_645/A 0.01fF
C45129 OR2X1_LOC_416/a_8_216# OR2X1_LOC_58/a_8_216# 0.47fF
C45130 OR2X1_LOC_287/B OR2X1_LOC_557/A 2.24fF
C45131 OR2X1_LOC_44/Y OR2X1_LOC_27/Y 0.05fF
C45132 OR2X1_LOC_5/a_8_216# OR2X1_LOC_6/A 0.01fF
C45133 OR2X1_LOC_358/a_8_216# OR2X1_LOC_476/B 0.01fF
C45134 OR2X1_LOC_385/Y OR2X1_LOC_743/A 0.02fF
C45135 AND2X1_LOC_729/Y OR2X1_LOC_601/a_8_216# 0.05fF
C45136 AND2X1_LOC_778/a_8_24# OR2X1_LOC_527/Y 0.01fF
C45137 OR2X1_LOC_600/A OR2X1_LOC_749/a_8_216# 0.01fF
C45138 AND2X1_LOC_784/A OR2X1_LOC_417/Y 0.03fF
C45139 OR2X1_LOC_741/Y OR2X1_LOC_318/B 0.14fF
C45140 AND2X1_LOC_866/B GATE_662 0.03fF
C45141 AND2X1_LOC_191/Y AND2X1_LOC_578/A 0.07fF
C45142 AND2X1_LOC_388/Y OR2X1_LOC_534/Y 0.01fF
C45143 AND2X1_LOC_512/a_8_24# AND2X1_LOC_729/B 0.01fF
C45144 OR2X1_LOC_95/Y OR2X1_LOC_278/Y 0.03fF
C45145 OR2X1_LOC_186/Y OR2X1_LOC_446/B 0.57fF
C45146 OR2X1_LOC_409/B OR2X1_LOC_48/B 0.12fF
C45147 OR2X1_LOC_685/B AND2X1_LOC_425/Y 0.00fF
C45148 AND2X1_LOC_64/Y OR2X1_LOC_703/Y 0.02fF
C45149 OR2X1_LOC_278/A AND2X1_LOC_852/Y 0.65fF
C45150 OR2X1_LOC_130/A D_INPUT_0 0.02fF
C45151 AND2X1_LOC_711/Y AND2X1_LOC_578/A 0.07fF
C45152 AND2X1_LOC_593/Y OR2X1_LOC_31/Y 0.01fF
C45153 OR2X1_LOC_186/Y OR2X1_LOC_303/B 0.01fF
C45154 OR2X1_LOC_18/Y OR2X1_LOC_409/B 0.05fF
C45155 OR2X1_LOC_533/Y OR2X1_LOC_13/B 0.09fF
C45156 OR2X1_LOC_70/Y AND2X1_LOC_578/A 0.22fF
C45157 INPUT_4 OR2X1_LOC_70/a_8_216# 0.00fF
C45158 AND2X1_LOC_25/Y AND2X1_LOC_7/Y 0.00fF
C45159 OR2X1_LOC_485/A AND2X1_LOC_830/a_36_24# 0.00fF
C45160 OR2X1_LOC_102/a_36_216# OR2X1_LOC_437/A 0.00fF
C45161 AND2X1_LOC_658/A AND2X1_LOC_657/A 0.07fF
C45162 AND2X1_LOC_721/Y OR2X1_LOC_183/Y 0.02fF
C45163 OR2X1_LOC_520/A AND2X1_LOC_8/Y 0.01fF
C45164 AND2X1_LOC_40/Y OR2X1_LOC_804/A 0.01fF
C45165 OR2X1_LOC_756/B OR2X1_LOC_675/Y 0.03fF
C45166 OR2X1_LOC_59/Y OR2X1_LOC_172/a_8_216# 0.00fF
C45167 VDD OR2X1_LOC_521/a_8_216# 0.21fF
C45168 OR2X1_LOC_31/Y OR2X1_LOC_85/A 0.03fF
C45169 AND2X1_LOC_337/B AND2X1_LOC_727/A 0.02fF
C45170 AND2X1_LOC_733/Y AND2X1_LOC_804/a_36_24# 0.00fF
C45171 AND2X1_LOC_845/Y AND2X1_LOC_806/A 0.15fF
C45172 OR2X1_LOC_737/A OR2X1_LOC_733/Y 0.16fF
C45173 AND2X1_LOC_18/Y OR2X1_LOC_367/B 0.03fF
C45174 AND2X1_LOC_565/Y OR2X1_LOC_95/Y 0.01fF
C45175 AND2X1_LOC_578/A AND2X1_LOC_514/Y 0.01fF
C45176 OR2X1_LOC_139/a_36_216# OR2X1_LOC_720/B 0.02fF
C45177 OR2X1_LOC_485/A AND2X1_LOC_477/A 0.13fF
C45178 AND2X1_LOC_56/B OR2X1_LOC_651/A 0.02fF
C45179 OR2X1_LOC_70/Y AND2X1_LOC_635/a_8_24# 0.01fF
C45180 OR2X1_LOC_473/Y OR2X1_LOC_121/B 0.01fF
C45181 OR2X1_LOC_145/a_8_216# OR2X1_LOC_146/Y 0.40fF
C45182 OR2X1_LOC_696/A OR2X1_LOC_49/A 0.02fF
C45183 OR2X1_LOC_151/A OR2X1_LOC_469/B 0.07fF
C45184 VDD OR2X1_LOC_300/Y 0.08fF
C45185 OR2X1_LOC_497/Y OR2X1_LOC_224/Y 0.05fF
C45186 AND2X1_LOC_111/a_8_24# OR2X1_LOC_532/B 0.01fF
C45187 OR2X1_LOC_840/A OR2X1_LOC_68/B 0.06fF
C45188 OR2X1_LOC_385/Y OR2X1_LOC_409/B 0.01fF
C45189 OR2X1_LOC_392/B OR2X1_LOC_267/Y 0.03fF
C45190 OR2X1_LOC_49/A AND2X1_LOC_64/Y 0.06fF
C45191 D_INPUT_2 OR2X1_LOC_37/a_36_216# 0.03fF
C45192 D_INPUT_3 OR2X1_LOC_37/a_8_216# 0.04fF
C45193 OR2X1_LOC_516/Y AND2X1_LOC_476/Y 0.07fF
C45194 OR2X1_LOC_427/A AND2X1_LOC_562/Y 0.03fF
C45195 OR2X1_LOC_223/A OR2X1_LOC_564/B 0.62fF
C45196 OR2X1_LOC_217/a_8_216# OR2X1_LOC_786/Y 0.04fF
C45197 AND2X1_LOC_775/a_36_24# AND2X1_LOC_476/Y 0.00fF
C45198 OR2X1_LOC_585/A D_INPUT_1 0.06fF
C45199 AND2X1_LOC_866/A AND2X1_LOC_212/B 0.01fF
C45200 OR2X1_LOC_502/A AND2X1_LOC_406/a_8_24# 0.04fF
C45201 AND2X1_LOC_74/a_8_24# OR2X1_LOC_578/B 0.03fF
C45202 OR2X1_LOC_46/A OR2X1_LOC_77/a_8_216# 0.07fF
C45203 AND2X1_LOC_335/a_8_24# OR2X1_LOC_437/A 0.04fF
C45204 AND2X1_LOC_564/A AND2X1_LOC_213/B 0.03fF
C45205 AND2X1_LOC_64/Y OR2X1_LOC_596/A 0.03fF
C45206 AND2X1_LOC_573/A AND2X1_LOC_570/a_8_24# 0.03fF
C45207 OR2X1_LOC_158/A OR2X1_LOC_56/a_8_216# 0.02fF
C45208 OR2X1_LOC_62/B D_INPUT_0 0.23fF
C45209 OR2X1_LOC_158/A AND2X1_LOC_465/A 0.11fF
C45210 AND2X1_LOC_56/B OR2X1_LOC_728/B 0.02fF
C45211 OR2X1_LOC_696/A OR2X1_LOC_526/Y 0.14fF
C45212 OR2X1_LOC_744/Y AND2X1_LOC_213/B 0.13fF
C45213 AND2X1_LOC_361/a_36_24# OR2X1_LOC_106/Y 0.01fF
C45214 OR2X1_LOC_6/A AND2X1_LOC_222/Y 0.02fF
C45215 OR2X1_LOC_19/B OR2X1_LOC_95/Y 0.14fF
C45216 OR2X1_LOC_76/Y OR2X1_LOC_675/Y 0.01fF
C45217 AND2X1_LOC_706/Y AND2X1_LOC_703/Y 0.01fF
C45218 OR2X1_LOC_64/Y OR2X1_LOC_615/Y 0.02fF
C45219 OR2X1_LOC_308/A OR2X1_LOC_160/B 0.03fF
C45220 OR2X1_LOC_6/A OR2X1_LOC_68/B 0.02fF
C45221 AND2X1_LOC_476/Y OR2X1_LOC_373/a_8_216# 0.03fF
C45222 OR2X1_LOC_106/Y VDD 0.51fF
C45223 OR2X1_LOC_763/Y OR2X1_LOC_70/A 0.00fF
C45224 OR2X1_LOC_447/Y OR2X1_LOC_454/a_8_216# 0.02fF
C45225 AND2X1_LOC_800/a_8_24# OR2X1_LOC_95/Y 0.01fF
C45226 OR2X1_LOC_519/Y OR2X1_LOC_437/A 0.00fF
C45227 OR2X1_LOC_696/A OR2X1_LOC_310/Y 0.03fF
C45228 AND2X1_LOC_350/a_8_24# AND2X1_LOC_339/B 0.02fF
C45229 OR2X1_LOC_161/A OR2X1_LOC_515/a_8_216# 0.05fF
C45230 AND2X1_LOC_794/B AND2X1_LOC_515/a_8_24# 0.01fF
C45231 AND2X1_LOC_555/Y OR2X1_LOC_744/A 0.00fF
C45232 AND2X1_LOC_619/B AND2X1_LOC_36/Y 0.10fF
C45233 OR2X1_LOC_409/Y OR2X1_LOC_22/A 0.01fF
C45234 OR2X1_LOC_604/A OR2X1_LOC_428/A 0.31fF
C45235 OR2X1_LOC_319/B OR2X1_LOC_319/Y 0.03fF
C45236 AND2X1_LOC_191/B AND2X1_LOC_580/a_8_24# 0.01fF
C45237 AND2X1_LOC_632/A OR2X1_LOC_615/Y 0.16fF
C45238 OR2X1_LOC_628/Y AND2X1_LOC_623/a_8_24# 0.01fF
C45239 AND2X1_LOC_95/Y OR2X1_LOC_342/B 0.26fF
C45240 AND2X1_LOC_482/a_8_24# AND2X1_LOC_36/Y 0.01fF
C45241 VDD OR2X1_LOC_691/Y 0.31fF
C45242 AND2X1_LOC_59/Y OR2X1_LOC_788/B 0.27fF
C45243 AND2X1_LOC_373/a_8_24# OR2X1_LOC_578/B 0.01fF
C45244 OR2X1_LOC_160/A OR2X1_LOC_712/B 0.00fF
C45245 VDD AND2X1_LOC_219/A 0.29fF
C45246 VDD OR2X1_LOC_375/Y 0.33fF
C45247 VDD OR2X1_LOC_43/Y 0.16fF
C45248 OR2X1_LOC_59/Y AND2X1_LOC_202/Y 0.52fF
C45249 OR2X1_LOC_417/A OR2X1_LOC_615/Y 0.04fF
C45250 OR2X1_LOC_641/A OR2X1_LOC_549/A 0.07fF
C45251 AND2X1_LOC_42/B OR2X1_LOC_560/A 0.00fF
C45252 OR2X1_LOC_51/Y AND2X1_LOC_639/B 0.34fF
C45253 OR2X1_LOC_70/Y OR2X1_LOC_172/a_8_216# 0.01fF
C45254 AND2X1_LOC_340/Y OR2X1_LOC_426/B 0.10fF
C45255 AND2X1_LOC_22/Y OR2X1_LOC_168/B 0.15fF
C45256 OR2X1_LOC_62/A D_INPUT_3 1.06fF
C45257 OR2X1_LOC_678/Y AND2X1_LOC_7/B 0.01fF
C45258 OR2X1_LOC_45/B OR2X1_LOC_91/A 0.91fF
C45259 OR2X1_LOC_324/a_8_216# AND2X1_LOC_64/Y 0.01fF
C45260 OR2X1_LOC_835/B OR2X1_LOC_771/B 0.07fF
C45261 OR2X1_LOC_145/Y OR2X1_LOC_146/Y 0.09fF
C45262 OR2X1_LOC_11/Y D_INPUT_6 0.70fF
C45263 OR2X1_LOC_9/a_8_216# OR2X1_LOC_56/A 0.01fF
C45264 OR2X1_LOC_51/Y OR2X1_LOC_604/Y 0.01fF
C45265 OR2X1_LOC_632/a_8_216# OR2X1_LOC_161/B 0.03fF
C45266 OR2X1_LOC_97/A OR2X1_LOC_334/B 0.01fF
C45267 OR2X1_LOC_40/Y OR2X1_LOC_96/Y 0.01fF
C45268 OR2X1_LOC_281/Y OR2X1_LOC_56/A 0.16fF
C45269 AND2X1_LOC_319/a_8_24# AND2X1_LOC_798/A 0.02fF
C45270 OR2X1_LOC_696/A OR2X1_LOC_433/Y 0.02fF
C45271 OR2X1_LOC_600/A AND2X1_LOC_243/Y 0.07fF
C45272 OR2X1_LOC_637/A OR2X1_LOC_855/A 0.19fF
C45273 OR2X1_LOC_529/Y OR2X1_LOC_437/A 0.07fF
C45274 AND2X1_LOC_529/a_8_24# OR2X1_LOC_633/A 0.01fF
C45275 OR2X1_LOC_369/Y AND2X1_LOC_476/Y -0.03fF
C45276 AND2X1_LOC_64/Y OR2X1_LOC_732/a_8_216# 0.01fF
C45277 VDD AND2X1_LOC_207/A 0.25fF
C45278 AND2X1_LOC_719/Y AND2X1_LOC_191/B 0.07fF
C45279 AND2X1_LOC_565/B AND2X1_LOC_549/Y 0.09fF
C45280 VDD OR2X1_LOC_505/Y 0.19fF
C45281 AND2X1_LOC_568/B OR2X1_LOC_600/A 0.17fF
C45282 OR2X1_LOC_56/A OR2X1_LOC_253/Y 0.03fF
C45283 VDD OR2X1_LOC_679/a_8_216# 0.21fF
C45284 OR2X1_LOC_303/a_8_216# OR2X1_LOC_212/A 0.01fF
C45285 INPUT_5 INPUT_7 0.70fF
C45286 OR2X1_LOC_741/Y OR2X1_LOC_190/a_8_216# 0.02fF
C45287 OR2X1_LOC_811/A AND2X1_LOC_7/B 0.03fF
C45288 OR2X1_LOC_653/B OR2X1_LOC_756/B 0.01fF
C45289 OR2X1_LOC_78/A OR2X1_LOC_362/A 0.66fF
C45290 OR2X1_LOC_629/B AND2X1_LOC_92/Y 0.01fF
C45291 VDD AND2X1_LOC_658/A 0.32fF
C45292 OR2X1_LOC_151/A AND2X1_LOC_167/a_8_24# 0.03fF
C45293 OR2X1_LOC_40/Y AND2X1_LOC_663/A 0.14fF
C45294 VDD OR2X1_LOC_690/Y 0.10fF
C45295 OR2X1_LOC_92/Y OR2X1_LOC_12/Y 7.34fF
C45296 VDD OR2X1_LOC_803/A -0.00fF
C45297 OR2X1_LOC_124/A VDD 0.05fF
C45298 OR2X1_LOC_850/a_8_216# OR2X1_LOC_362/A 0.01fF
C45299 AND2X1_LOC_787/A AND2X1_LOC_468/B 0.01fF
C45300 VDD OR2X1_LOC_242/a_8_216# 0.00fF
C45301 OR2X1_LOC_196/B OR2X1_LOC_446/B 0.10fF
C45302 OR2X1_LOC_656/B AND2X1_LOC_44/Y 0.03fF
C45303 OR2X1_LOC_160/A OR2X1_LOC_139/A 0.03fF
C45304 OR2X1_LOC_503/A AND2X1_LOC_242/B 0.02fF
C45305 OR2X1_LOC_64/Y OR2X1_LOC_424/Y 0.01fF
C45306 AND2X1_LOC_776/a_8_24# OR2X1_LOC_329/B 0.13fF
C45307 AND2X1_LOC_773/Y OR2X1_LOC_619/Y 0.10fF
C45308 OR2X1_LOC_45/B AND2X1_LOC_573/A 0.06fF
C45309 AND2X1_LOC_59/Y AND2X1_LOC_22/Y 1.70fF
C45310 OR2X1_LOC_744/A OR2X1_LOC_51/Y 0.41fF
C45311 AND2X1_LOC_40/Y OR2X1_LOC_797/B 0.35fF
C45312 OR2X1_LOC_528/Y AND2X1_LOC_185/a_8_24# 0.11fF
C45313 OR2X1_LOC_813/Y AND2X1_LOC_845/a_8_24# 0.05fF
C45314 OR2X1_LOC_427/A OR2X1_LOC_381/a_8_216# 0.01fF
C45315 AND2X1_LOC_658/B OR2X1_LOC_524/Y 0.39fF
C45316 OR2X1_LOC_185/A AND2X1_LOC_603/a_8_24# 0.01fF
C45317 OR2X1_LOC_821/Y OR2X1_LOC_278/Y 0.26fF
C45318 OR2X1_LOC_696/A AND2X1_LOC_259/Y 0.00fF
C45319 AND2X1_LOC_56/B OR2X1_LOC_338/A 0.20fF
C45320 OR2X1_LOC_241/Y OR2X1_LOC_68/B 0.43fF
C45321 AND2X1_LOC_575/a_8_24# AND2X1_LOC_576/Y 0.04fF
C45322 OR2X1_LOC_161/A OR2X1_LOC_706/a_8_216# 0.05fF
C45323 GATE_479 AND2X1_LOC_222/Y 0.01fF
C45324 OR2X1_LOC_235/B OR2X1_LOC_244/Y 0.02fF
C45325 OR2X1_LOC_306/Y OR2X1_LOC_428/A 0.05fF
C45326 OR2X1_LOC_177/Y OR2X1_LOC_109/a_36_216# 0.00fF
C45327 OR2X1_LOC_85/A OR2X1_LOC_79/a_8_216# 0.14fF
C45328 OR2X1_LOC_65/B OR2X1_LOC_12/Y 0.05fF
C45329 OR2X1_LOC_64/Y D_INPUT_6 0.11fF
C45330 OR2X1_LOC_40/Y OR2X1_LOC_2/Y 0.09fF
C45331 OR2X1_LOC_39/A OR2X1_LOC_522/Y 0.02fF
C45332 OR2X1_LOC_240/A OR2X1_LOC_415/Y 0.44fF
C45333 OR2X1_LOC_677/Y AND2X1_LOC_658/A 0.10fF
C45334 AND2X1_LOC_695/a_36_24# OR2X1_LOC_161/B 0.00fF
C45335 AND2X1_LOC_508/A AND2X1_LOC_510/A 0.27fF
C45336 OR2X1_LOC_255/a_8_216# OR2X1_LOC_13/B 0.01fF
C45337 OR2X1_LOC_793/A AND2X1_LOC_44/Y 0.07fF
C45338 OR2X1_LOC_128/B OR2X1_LOC_151/A 0.01fF
C45339 AND2X1_LOC_555/Y OR2X1_LOC_282/a_8_216# 0.01fF
C45340 AND2X1_LOC_64/Y OR2X1_LOC_33/B 0.03fF
C45341 OR2X1_LOC_175/B OR2X1_LOC_66/A 0.02fF
C45342 VDD OR2X1_LOC_629/Y 0.00fF
C45343 OR2X1_LOC_689/A OR2X1_LOC_690/Y 0.09fF
C45344 OR2X1_LOC_406/Y AND2X1_LOC_474/Y 0.00fF
C45345 OR2X1_LOC_474/Y OR2X1_LOC_78/A 0.03fF
C45346 OR2X1_LOC_186/Y AND2X1_LOC_56/B 0.11fF
C45347 AND2X1_LOC_574/a_8_24# AND2X1_LOC_508/A 0.20fF
C45348 AND2X1_LOC_60/a_8_24# OR2X1_LOC_219/B 0.04fF
C45349 AND2X1_LOC_95/Y AND2X1_LOC_322/a_36_24# 0.00fF
C45350 OR2X1_LOC_676/Y OR2X1_LOC_194/B 0.01fF
C45351 OR2X1_LOC_585/A OR2X1_LOC_585/a_8_216# 0.05fF
C45352 OR2X1_LOC_585/A OR2X1_LOC_15/a_8_216# 0.01fF
C45353 AND2X1_LOC_568/B OR2X1_LOC_619/Y 0.03fF
C45354 VDD OR2X1_LOC_249/a_8_216# 0.00fF
C45355 OR2X1_LOC_76/Y OR2X1_LOC_736/Y 0.03fF
C45356 OR2X1_LOC_114/Y OR2X1_LOC_549/A 0.04fF
C45357 VDD AND2X1_LOC_847/Y 0.88fF
C45358 OR2X1_LOC_756/B OR2X1_LOC_808/B 0.03fF
C45359 AND2X1_LOC_535/Y AND2X1_LOC_356/a_36_24# 0.00fF
C45360 OR2X1_LOC_604/A AND2X1_LOC_154/a_8_24# 0.01fF
C45361 OR2X1_LOC_598/Y OR2X1_LOC_130/A 0.00fF
C45362 OR2X1_LOC_543/a_36_216# OR2X1_LOC_552/A 0.00fF
C45363 AND2X1_LOC_507/a_36_24# OR2X1_LOC_18/Y 0.00fF
C45364 OR2X1_LOC_675/A OR2X1_LOC_722/B 0.00fF
C45365 OR2X1_LOC_771/a_36_216# OR2X1_LOC_80/A 0.00fF
C45366 AND2X1_LOC_703/Y OR2X1_LOC_485/A 0.01fF
C45367 AND2X1_LOC_173/a_8_24# OR2X1_LOC_538/A 0.01fF
C45368 AND2X1_LOC_3/Y OR2X1_LOC_161/B 2.57fF
C45369 OR2X1_LOC_129/a_8_216# OR2X1_LOC_85/A 0.05fF
C45370 AND2X1_LOC_592/Y OR2X1_LOC_36/Y 0.04fF
C45371 OR2X1_LOC_641/Y OR2X1_LOC_660/B 0.01fF
C45372 OR2X1_LOC_102/a_36_216# OR2X1_LOC_753/A 0.01fF
C45373 OR2X1_LOC_754/A OR2X1_LOC_816/A 0.11fF
C45374 OR2X1_LOC_168/a_8_216# OR2X1_LOC_78/B 0.06fF
C45375 AND2X1_LOC_719/Y AND2X1_LOC_862/a_8_24# 0.20fF
C45376 AND2X1_LOC_720/a_36_24# OR2X1_LOC_59/Y 0.01fF
C45377 OR2X1_LOC_64/Y AND2X1_LOC_242/B 0.19fF
C45378 AND2X1_LOC_766/a_8_24# OR2X1_LOC_401/B 0.20fF
C45379 OR2X1_LOC_770/A OR2X1_LOC_401/A 0.16fF
C45380 OR2X1_LOC_641/B OR2X1_LOC_228/Y 0.09fF
C45381 OR2X1_LOC_201/A OR2X1_LOC_61/Y 0.22fF
C45382 OR2X1_LOC_492/a_8_216# OR2X1_LOC_485/A 0.01fF
C45383 VDD OR2X1_LOC_497/a_8_216# 0.21fF
C45384 OR2X1_LOC_482/a_8_216# OR2X1_LOC_666/Y 0.40fF
C45385 OR2X1_LOC_671/Y OR2X1_LOC_827/Y 0.01fF
C45386 OR2X1_LOC_710/B OR2X1_LOC_154/A 0.03fF
C45387 OR2X1_LOC_6/B OR2X1_LOC_753/A 0.12fF
C45388 OR2X1_LOC_646/A OR2X1_LOC_646/B 0.02fF
C45389 OR2X1_LOC_422/a_8_216# OR2X1_LOC_92/Y 0.02fF
C45390 AND2X1_LOC_707/Y OR2X1_LOC_64/Y 0.02fF
C45391 OR2X1_LOC_814/A AND2X1_LOC_226/a_8_24# 0.07fF
C45392 AND2X1_LOC_114/a_8_24# OR2X1_LOC_59/Y 0.01fF
C45393 OR2X1_LOC_56/A OR2X1_LOC_48/a_8_216# 0.07fF
C45394 AND2X1_LOC_724/Y OR2X1_LOC_44/Y 0.01fF
C45395 OR2X1_LOC_326/a_8_216# AND2X1_LOC_59/Y 0.00fF
C45396 AND2X1_LOC_84/Y AND2X1_LOC_633/Y 0.02fF
C45397 OR2X1_LOC_291/Y AND2X1_LOC_206/a_8_24# 0.03fF
C45398 AND2X1_LOC_756/a_36_24# OR2X1_LOC_616/Y 0.00fF
C45399 OR2X1_LOC_49/A AND2X1_LOC_663/B 0.03fF
C45400 OR2X1_LOC_160/A OR2X1_LOC_637/Y 0.00fF
C45401 AND2X1_LOC_159/a_8_24# AND2X1_LOC_18/Y 0.06fF
C45402 OR2X1_LOC_51/Y AND2X1_LOC_840/B 0.12fF
C45403 OR2X1_LOC_744/A OR2X1_LOC_680/A 0.07fF
C45404 OR2X1_LOC_832/a_8_216# OR2X1_LOC_155/A 0.03fF
C45405 OR2X1_LOC_810/A AND2X1_LOC_18/Y 0.17fF
C45406 AND2X1_LOC_170/a_36_24# OR2X1_LOC_91/A 0.00fF
C45407 OR2X1_LOC_506/A OR2X1_LOC_776/a_8_216# 0.14fF
C45408 AND2X1_LOC_191/Y AND2X1_LOC_478/a_8_24# 0.05fF
C45409 OR2X1_LOC_217/Y OR2X1_LOC_78/A 0.03fF
C45410 OR2X1_LOC_71/A OR2X1_LOC_398/a_36_216# 0.00fF
C45411 OR2X1_LOC_96/Y OR2X1_LOC_7/A 0.00fF
C45412 AND2X1_LOC_45/a_8_24# AND2X1_LOC_44/Y 0.01fF
C45413 OR2X1_LOC_235/B AND2X1_LOC_669/a_8_24# 0.01fF
C45414 AND2X1_LOC_95/Y OR2X1_LOC_623/B 1.38fF
C45415 OR2X1_LOC_323/A OR2X1_LOC_95/Y 0.06fF
C45416 OR2X1_LOC_426/B OR2X1_LOC_585/A 0.03fF
C45417 AND2X1_LOC_578/A AND2X1_LOC_499/a_8_24# 0.04fF
C45418 AND2X1_LOC_362/a_8_24# OR2X1_LOC_44/Y 0.01fF
C45419 OR2X1_LOC_160/B OR2X1_LOC_557/A 0.03fF
C45420 OR2X1_LOC_323/A OR2X1_LOC_368/A 0.50fF
C45421 OR2X1_LOC_118/a_8_216# OR2X1_LOC_22/Y 0.02fF
C45422 OR2X1_LOC_532/B OR2X1_LOC_267/Y 0.02fF
C45423 OR2X1_LOC_374/Y OR2X1_LOC_590/Y 0.00fF
C45424 OR2X1_LOC_7/A AND2X1_LOC_454/a_8_24# 0.04fF
C45425 OR2X1_LOC_547/B OR2X1_LOC_620/Y 0.97fF
C45426 AND2X1_LOC_40/Y OR2X1_LOC_340/Y 0.14fF
C45427 AND2X1_LOC_367/A OR2X1_LOC_6/A 0.03fF
C45428 OR2X1_LOC_40/Y AND2X1_LOC_212/B 0.14fF
C45429 OR2X1_LOC_849/A OR2X1_LOC_78/B 0.00fF
C45430 OR2X1_LOC_154/A OR2X1_LOC_663/A 0.19fF
C45431 INPUT_5 INPUT_4 0.29fF
C45432 OR2X1_LOC_637/B OR2X1_LOC_828/B 0.00fF
C45433 AND2X1_LOC_512/Y OR2X1_LOC_36/Y 0.42fF
C45434 AND2X1_LOC_356/B OR2X1_LOC_56/A 0.09fF
C45435 AND2X1_LOC_532/a_8_24# AND2X1_LOC_468/B 0.01fF
C45436 AND2X1_LOC_40/Y OR2X1_LOC_130/A 0.07fF
C45437 OR2X1_LOC_849/A AND2X1_LOC_103/a_36_24# 0.00fF
C45438 OR2X1_LOC_100/Y OR2X1_LOC_520/Y 0.01fF
C45439 AND2X1_LOC_729/B AND2X1_LOC_200/a_8_24# 0.01fF
C45440 AND2X1_LOC_520/a_36_24# OR2X1_LOC_417/A 0.01fF
C45441 OR2X1_LOC_280/Y OR2X1_LOC_56/A 0.03fF
C45442 AND2X1_LOC_658/B AND2X1_LOC_578/A 0.07fF
C45443 OR2X1_LOC_7/A AND2X1_LOC_663/A 0.51fF
C45444 OR2X1_LOC_852/a_8_216# D_INPUT_0 -0.00fF
C45445 INPUT_1 OR2X1_LOC_16/A 2.12fF
C45446 OR2X1_LOC_49/A OR2X1_LOC_54/a_8_216# 0.06fF
C45447 OR2X1_LOC_405/A OR2X1_LOC_185/A 9.54fF
C45448 OR2X1_LOC_844/a_8_216# OR2X1_LOC_244/Y 0.00fF
C45449 OR2X1_LOC_663/A OR2X1_LOC_267/A 0.03fF
C45450 OR2X1_LOC_811/A OR2X1_LOC_805/A 0.30fF
C45451 OR2X1_LOC_680/a_8_216# AND2X1_LOC_796/Y 0.01fF
C45452 OR2X1_LOC_409/B OR2X1_LOC_764/a_8_216# 0.00fF
C45453 OR2X1_LOC_160/B OR2X1_LOC_675/A 0.01fF
C45454 OR2X1_LOC_532/B OR2X1_LOC_633/A 0.87fF
C45455 OR2X1_LOC_813/a_8_216# OR2X1_LOC_64/Y 0.01fF
C45456 OR2X1_LOC_772/B OR2X1_LOC_772/a_8_216# 0.01fF
C45457 OR2X1_LOC_325/B OR2X1_LOC_121/B 0.01fF
C45458 OR2X1_LOC_48/Y OR2X1_LOC_59/Y 0.00fF
C45459 AND2X1_LOC_448/Y AND2X1_LOC_452/Y 0.02fF
C45460 INPUT_5 AND2X1_LOC_51/A 1.17fF
C45461 AND2X1_LOC_59/Y OR2X1_LOC_664/a_8_216# 0.14fF
C45462 OR2X1_LOC_449/B AND2X1_LOC_423/a_8_24# 0.07fF
C45463 OR2X1_LOC_185/Y OR2X1_LOC_620/Y 0.30fF
C45464 OR2X1_LOC_421/A OR2X1_LOC_46/A 0.00fF
C45465 AND2X1_LOC_850/Y AND2X1_LOC_286/Y 0.08fF
C45466 OR2X1_LOC_673/a_8_216# OR2X1_LOC_532/B 0.04fF
C45467 INPUT_0 AND2X1_LOC_13/a_8_24# 0.03fF
C45468 AND2X1_LOC_332/a_8_24# OR2X1_LOC_31/Y 0.03fF
C45469 OR2X1_LOC_473/a_8_216# OR2X1_LOC_810/A 0.15fF
C45470 OR2X1_LOC_778/A OR2X1_LOC_778/a_8_216# 0.04fF
C45471 OR2X1_LOC_294/a_8_216# OR2X1_LOC_296/Y 0.01fF
C45472 VDD AND2X1_LOC_814/a_8_24# 0.00fF
C45473 AND2X1_LOC_580/A AND2X1_LOC_858/a_8_24# 0.04fF
C45474 AND2X1_LOC_64/Y OR2X1_LOC_374/Y 0.05fF
C45475 OR2X1_LOC_589/A OR2X1_LOC_72/a_8_216# 0.01fF
C45476 VDD OR2X1_LOC_750/a_8_216# 0.21fF
C45477 OR2X1_LOC_86/Y OR2X1_LOC_18/Y 0.02fF
C45478 OR2X1_LOC_47/Y AND2X1_LOC_786/Y 0.03fF
C45479 OR2X1_LOC_497/Y OR2X1_LOC_18/Y 0.00fF
C45480 OR2X1_LOC_137/a_8_216# OR2X1_LOC_404/Y 0.00fF
C45481 INPUT_7 OR2X1_LOC_17/a_8_216# 0.00fF
C45482 OR2X1_LOC_61/Y AND2X1_LOC_3/Y 0.07fF
C45483 OR2X1_LOC_270/Y OR2X1_LOC_161/B 0.03fF
C45484 AND2X1_LOC_576/Y AND2X1_LOC_624/A 0.07fF
C45485 OR2X1_LOC_219/a_8_216# OR2X1_LOC_222/A 0.01fF
C45486 AND2X1_LOC_72/B OR2X1_LOC_563/A 0.01fF
C45487 AND2X1_LOC_12/Y AND2X1_LOC_817/a_8_24# 0.01fF
C45488 AND2X1_LOC_347/Y OR2X1_LOC_481/A 0.11fF
C45489 AND2X1_LOC_702/Y OR2X1_LOC_298/Y 0.00fF
C45490 OR2X1_LOC_32/B OR2X1_LOC_44/Y 0.21fF
C45491 OR2X1_LOC_600/a_36_216# AND2X1_LOC_477/A 0.02fF
C45492 AND2X1_LOC_339/B AND2X1_LOC_660/A 0.01fF
C45493 OR2X1_LOC_287/B OR2X1_LOC_814/Y 0.01fF
C45494 OR2X1_LOC_22/Y OR2X1_LOC_56/A 0.21fF
C45495 AND2X1_LOC_70/Y OR2X1_LOC_814/A 0.14fF
C45496 OR2X1_LOC_680/A AND2X1_LOC_840/B 0.20fF
C45497 OR2X1_LOC_364/A OR2X1_LOC_154/A 0.13fF
C45498 OR2X1_LOC_185/Y OR2X1_LOC_154/A 0.54fF
C45499 OR2X1_LOC_3/Y AND2X1_LOC_364/A 0.12fF
C45500 OR2X1_LOC_715/B OR2X1_LOC_506/B 0.01fF
C45501 OR2X1_LOC_377/A OR2X1_LOC_472/A 0.07fF
C45502 OR2X1_LOC_664/Y OR2X1_LOC_631/B 0.18fF
C45503 AND2X1_LOC_71/a_36_24# OR2X1_LOC_404/Y 0.01fF
C45504 OR2X1_LOC_849/A OR2X1_LOC_375/A 0.03fF
C45505 OR2X1_LOC_40/a_8_216# OR2X1_LOC_17/Y 0.01fF
C45506 OR2X1_LOC_799/A OR2X1_LOC_574/A 0.15fF
C45507 OR2X1_LOC_520/A AND2X1_LOC_92/Y 0.01fF
C45508 AND2X1_LOC_563/A AND2X1_LOC_227/Y 0.01fF
C45509 OR2X1_LOC_48/B OR2X1_LOC_229/Y 0.22fF
C45510 AND2X1_LOC_110/a_8_24# OR2X1_LOC_532/B 0.01fF
C45511 AND2X1_LOC_193/a_8_24# OR2X1_LOC_43/A 0.01fF
C45512 OR2X1_LOC_62/B OR2X1_LOC_612/Y 0.01fF
C45513 OR2X1_LOC_516/a_8_216# OR2X1_LOC_26/Y 0.03fF
C45514 OR2X1_LOC_171/Y OR2X1_LOC_172/Y 0.01fF
C45515 OR2X1_LOC_91/Y OR2X1_LOC_52/B 0.00fF
C45516 OR2X1_LOC_472/A AND2X1_LOC_824/B 4.83fF
C45517 OR2X1_LOC_7/A AND2X1_LOC_449/Y 0.01fF
C45518 OR2X1_LOC_704/a_8_216# OR2X1_LOC_308/Y 0.03fF
C45519 OR2X1_LOC_51/Y OR2X1_LOC_31/Y 0.21fF
C45520 OR2X1_LOC_643/A OR2X1_LOC_203/Y 0.07fF
C45521 OR2X1_LOC_692/a_36_216# OR2X1_LOC_64/Y 0.00fF
C45522 OR2X1_LOC_377/A OR2X1_LOC_647/A 0.03fF
C45523 OR2X1_LOC_203/Y OR2X1_LOC_124/Y 0.30fF
C45524 OR2X1_LOC_406/A AND2X1_LOC_795/a_8_24# 0.03fF
C45525 AND2X1_LOC_656/Y OR2X1_LOC_59/Y 0.00fF
C45526 OR2X1_LOC_8/Y D_INPUT_3 0.24fF
C45527 OR2X1_LOC_856/B AND2X1_LOC_135/a_36_24# 0.01fF
C45528 AND2X1_LOC_211/B AND2X1_LOC_303/B 0.21fF
C45529 AND2X1_LOC_673/a_8_24# OR2X1_LOC_6/A 0.01fF
C45530 OR2X1_LOC_91/Y AND2X1_LOC_489/Y 0.03fF
C45531 OR2X1_LOC_64/Y AND2X1_LOC_841/B 0.07fF
C45532 OR2X1_LOC_272/Y OR2X1_LOC_65/B 0.00fF
C45533 OR2X1_LOC_682/Y OR2X1_LOC_36/Y 0.02fF
C45534 OR2X1_LOC_460/Y AND2X1_LOC_3/Y 0.01fF
C45535 OR2X1_LOC_3/Y AND2X1_LOC_572/A 0.01fF
C45536 AND2X1_LOC_349/B AND2X1_LOC_349/a_8_24# 0.01fF
C45537 AND2X1_LOC_40/Y OR2X1_LOC_62/B 0.03fF
C45538 AND2X1_LOC_851/A AND2X1_LOC_465/Y 0.04fF
C45539 OR2X1_LOC_74/A OR2X1_LOC_6/A 0.10fF
C45540 OR2X1_LOC_306/a_36_216# AND2X1_LOC_729/B 0.01fF
C45541 OR2X1_LOC_748/A OR2X1_LOC_297/Y 0.01fF
C45542 OR2X1_LOC_121/B AND2X1_LOC_492/a_36_24# 0.00fF
C45543 AND2X1_LOC_105/a_36_24# OR2X1_LOC_26/Y 0.02fF
C45544 AND2X1_LOC_42/B OR2X1_LOC_267/a_8_216# 0.01fF
C45545 AND2X1_LOC_716/Y D_INPUT_0 -0.01fF
C45546 OR2X1_LOC_528/Y OR2X1_LOC_419/Y 0.07fF
C45547 OR2X1_LOC_501/B OR2X1_LOC_276/B 0.00fF
C45548 OR2X1_LOC_189/Y OR2X1_LOC_52/B 0.15fF
C45549 OR2X1_LOC_479/Y OR2X1_LOC_468/Y 5.32fF
C45550 OR2X1_LOC_92/Y AND2X1_LOC_801/B 0.01fF
C45551 AND2X1_LOC_738/B AND2X1_LOC_808/A 0.03fF
C45552 AND2X1_LOC_723/Y OR2X1_LOC_95/Y 0.46fF
C45553 OR2X1_LOC_675/A OR2X1_LOC_553/A 0.01fF
C45554 OR2X1_LOC_235/Y AND2X1_LOC_243/a_8_24# 0.23fF
C45555 OR2X1_LOC_474/a_8_216# OR2X1_LOC_624/A 0.13fF
C45556 OR2X1_LOC_185/Y OR2X1_LOC_778/A 0.02fF
C45557 OR2X1_LOC_748/A AND2X1_LOC_345/Y 0.12fF
C45558 OR2X1_LOC_750/A OR2X1_LOC_161/A 0.17fF
C45559 OR2X1_LOC_743/A OR2X1_LOC_585/A 0.05fF
C45560 OR2X1_LOC_26/Y OR2X1_LOC_83/a_8_216# 0.01fF
C45561 OR2X1_LOC_524/Y OR2X1_LOC_47/Y 0.65fF
C45562 OR2X1_LOC_31/Y OR2X1_LOC_16/Y 0.02fF
C45563 OR2X1_LOC_335/Y AND2X1_LOC_438/a_36_24# 0.01fF
C45564 AND2X1_LOC_456/Y AND2X1_LOC_465/a_8_24# 0.06fF
C45565 AND2X1_LOC_388/a_8_24# AND2X1_LOC_727/A 0.01fF
C45566 AND2X1_LOC_841/B OR2X1_LOC_417/A 0.11fF
C45567 AND2X1_LOC_12/Y OR2X1_LOC_773/a_8_216# 0.01fF
C45568 AND2X1_LOC_788/a_8_24# OR2X1_LOC_533/A 0.10fF
C45569 AND2X1_LOC_580/A AND2X1_LOC_664/a_8_24# 0.04fF
C45570 AND2X1_LOC_95/Y OR2X1_LOC_544/A 0.03fF
C45571 AND2X1_LOC_51/Y OR2X1_LOC_710/a_8_216# 0.01fF
C45572 AND2X1_LOC_7/B OR2X1_LOC_777/B 0.09fF
C45573 OR2X1_LOC_31/Y AND2X1_LOC_642/a_8_24# 0.05fF
C45574 OR2X1_LOC_490/Y AND2X1_LOC_557/a_8_24# 0.00fF
C45575 AND2X1_LOC_56/B OR2X1_LOC_196/B 0.00fF
C45576 OR2X1_LOC_36/Y OR2X1_LOC_54/Y 0.03fF
C45577 AND2X1_LOC_566/Y AND2X1_LOC_568/a_36_24# 0.01fF
C45578 AND2X1_LOC_40/Y AND2X1_LOC_88/Y 0.00fF
C45579 OR2X1_LOC_70/Y OR2X1_LOC_418/a_8_216# 0.01fF
C45580 OR2X1_LOC_417/Y OR2X1_LOC_52/B 0.07fF
C45581 OR2X1_LOC_291/Y OR2X1_LOC_52/B 0.03fF
C45582 AND2X1_LOC_194/Y OR2X1_LOC_39/a_8_216# 0.47fF
C45583 OR2X1_LOC_756/B AND2X1_LOC_289/a_8_24# 0.01fF
C45584 AND2X1_LOC_259/Y AND2X1_LOC_663/B 0.01fF
C45585 AND2X1_LOC_743/a_8_24# OR2X1_LOC_712/B 0.24fF
C45586 OR2X1_LOC_192/A OR2X1_LOC_192/a_8_216# 0.39fF
C45587 OR2X1_LOC_256/Y AND2X1_LOC_721/A 0.01fF
C45588 OR2X1_LOC_755/A OR2X1_LOC_757/Y 0.09fF
C45589 AND2X1_LOC_658/B OR2X1_LOC_746/Y 0.03fF
C45590 AND2X1_LOC_809/a_8_24# OR2X1_LOC_13/B 0.03fF
C45591 AND2X1_LOC_706/Y OR2X1_LOC_589/a_8_216# 0.04fF
C45592 OR2X1_LOC_311/Y OR2X1_LOC_52/B 0.03fF
C45593 OR2X1_LOC_742/B OR2X1_LOC_190/Y 0.00fF
C45594 OR2X1_LOC_335/Y OR2X1_LOC_365/B 0.03fF
C45595 AND2X1_LOC_512/Y OR2X1_LOC_419/Y 0.10fF
C45596 OR2X1_LOC_563/A AND2X1_LOC_36/Y 0.02fF
C45597 OR2X1_LOC_246/A OR2X1_LOC_585/A 0.06fF
C45598 AND2X1_LOC_512/a_8_24# OR2X1_LOC_46/A 0.17fF
C45599 OR2X1_LOC_440/A OR2X1_LOC_375/A 0.03fF
C45600 D_INPUT_3 OR2X1_LOC_67/A 0.03fF
C45601 OR2X1_LOC_856/B OR2X1_LOC_214/B 0.03fF
C45602 OR2X1_LOC_241/a_8_216# OR2X1_LOC_241/Y 0.02fF
C45603 VDD OR2X1_LOC_546/A 0.21fF
C45604 AND2X1_LOC_397/a_8_24# OR2X1_LOC_68/B 0.01fF
C45605 OR2X1_LOC_485/A AND2X1_LOC_465/Y 0.25fF
C45606 OR2X1_LOC_7/A OR2X1_LOC_7/Y 1.75fF
C45607 AND2X1_LOC_40/Y OR2X1_LOC_365/B 0.02fF
C45608 OR2X1_LOC_151/A OR2X1_LOC_535/a_8_216# 0.03fF
C45609 OR2X1_LOC_22/Y AND2X1_LOC_641/Y 0.08fF
C45610 OR2X1_LOC_95/Y OR2X1_LOC_601/Y 0.43fF
C45611 OR2X1_LOC_613/Y AND2X1_LOC_663/a_8_24# 0.01fF
C45612 INPUT_4 OR2X1_LOC_17/a_8_216# 0.01fF
C45613 OR2X1_LOC_66/A OR2X1_LOC_366/Y 0.60fF
C45614 AND2X1_LOC_64/Y OR2X1_LOC_392/B 0.04fF
C45615 OR2X1_LOC_43/A AND2X1_LOC_476/A 0.07fF
C45616 OR2X1_LOC_663/A OR2X1_LOC_560/A 0.03fF
C45617 OR2X1_LOC_848/B D_INPUT_1 0.00fF
C45618 OR2X1_LOC_273/a_8_216# INPUT_1 0.03fF
C45619 OR2X1_LOC_805/A AND2X1_LOC_237/a_8_24# 0.05fF
C45620 OR2X1_LOC_409/B OR2X1_LOC_585/A 0.01fF
C45621 OR2X1_LOC_831/B AND2X1_LOC_7/B 0.02fF
C45622 OR2X1_LOC_804/A AND2X1_LOC_43/B 0.07fF
C45623 AND2X1_LOC_227/Y AND2X1_LOC_717/B 0.03fF
C45624 D_INPUT_3 OR2X1_LOC_672/Y 0.02fF
C45625 OR2X1_LOC_188/a_8_216# AND2X1_LOC_7/B -0.04fF
C45626 AND2X1_LOC_721/Y AND2X1_LOC_465/A 0.02fF
C45627 OR2X1_LOC_484/a_8_216# OR2X1_LOC_437/A 0.01fF
C45628 OR2X1_LOC_404/Y OR2X1_LOC_814/A 0.03fF
C45629 OR2X1_LOC_516/A OR2X1_LOC_419/Y 0.01fF
C45630 AND2X1_LOC_280/a_8_24# OR2X1_LOC_161/A 0.01fF
C45631 AND2X1_LOC_564/B AND2X1_LOC_734/a_8_24# 0.01fF
C45632 AND2X1_LOC_489/Y D_INPUT_3 0.02fF
C45633 OR2X1_LOC_696/A AND2X1_LOC_714/B 0.01fF
C45634 AND2X1_LOC_272/a_36_24# OR2X1_LOC_493/Y 0.01fF
C45635 OR2X1_LOC_804/a_8_216# OR2X1_LOC_303/B 0.01fF
C45636 OR2X1_LOC_605/B OR2X1_LOC_440/A 0.03fF
C45637 OR2X1_LOC_78/A OR2X1_LOC_771/B 0.03fF
C45638 AND2X1_LOC_42/B AND2X1_LOC_813/a_8_24# 0.01fF
C45639 AND2X1_LOC_128/a_8_24# INPUT_1 0.09fF
C45640 AND2X1_LOC_647/Y OR2X1_LOC_6/A 0.00fF
C45641 OR2X1_LOC_626/a_36_216# AND2X1_LOC_624/B 0.00fF
C45642 AND2X1_LOC_116/a_8_24# AND2X1_LOC_116/Y 0.01fF
C45643 AND2X1_LOC_400/a_8_24# OR2X1_LOC_80/A 0.03fF
C45644 AND2X1_LOC_7/B OR2X1_LOC_344/A 0.04fF
C45645 AND2X1_LOC_578/A OR2X1_LOC_47/Y 3.28fF
C45646 OR2X1_LOC_499/a_8_216# OR2X1_LOC_68/B 0.05fF
C45647 OR2X1_LOC_318/a_8_216# AND2X1_LOC_22/Y 0.01fF
C45648 OR2X1_LOC_496/Y OR2X1_LOC_406/A 0.01fF
C45649 OR2X1_LOC_753/A OR2X1_LOC_598/A 1.12fF
C45650 OR2X1_LOC_319/B OR2X1_LOC_777/B 0.07fF
C45651 AND2X1_LOC_733/a_36_24# OR2X1_LOC_437/A 0.00fF
C45652 AND2X1_LOC_844/a_36_24# OR2X1_LOC_95/Y 0.00fF
C45653 OR2X1_LOC_44/Y AND2X1_LOC_222/Y 0.03fF
C45654 AND2X1_LOC_572/A AND2X1_LOC_772/a_8_24# 0.01fF
C45655 OR2X1_LOC_755/Y AND2X1_LOC_791/a_8_24# 0.23fF
C45656 D_GATE_579 OR2X1_LOC_269/B 0.00fF
C45657 AND2X1_LOC_347/Y AND2X1_LOC_789/Y 0.22fF
C45658 OR2X1_LOC_468/Y OR2X1_LOC_566/a_36_216# 0.00fF
C45659 OR2X1_LOC_185/Y OR2X1_LOC_560/A 0.05fF
C45660 OR2X1_LOC_92/Y OR2X1_LOC_248/A 0.03fF
C45661 OR2X1_LOC_269/B OR2X1_LOC_228/Y 0.07fF
C45662 AND2X1_LOC_476/A AND2X1_LOC_462/a_36_24# 0.01fF
C45663 OR2X1_LOC_632/Y OR2X1_LOC_501/A 0.03fF
C45664 OR2X1_LOC_160/A OR2X1_LOC_728/A 0.05fF
C45665 OR2X1_LOC_851/A OR2X1_LOC_593/B 0.01fF
C45666 AND2X1_LOC_566/B OR2X1_LOC_135/Y 0.01fF
C45667 OR2X1_LOC_59/Y AND2X1_LOC_772/Y 0.00fF
C45668 OR2X1_LOC_246/Y OR2X1_LOC_150/a_8_216# 0.03fF
C45669 AND2X1_LOC_758/a_36_24# GATE_579 0.00fF
C45670 OR2X1_LOC_709/B OR2X1_LOC_711/B 0.83fF
C45671 AND2X1_LOC_65/A AND2X1_LOC_262/a_8_24# 0.00fF
C45672 OR2X1_LOC_44/Y OR2X1_LOC_423/Y 0.03fF
C45673 AND2X1_LOC_814/a_8_24# AND2X1_LOC_624/B 0.03fF
C45674 OR2X1_LOC_805/A OR2X1_LOC_777/B 0.07fF
C45675 OR2X1_LOC_600/A OR2X1_LOC_12/Y 0.27fF
C45676 OR2X1_LOC_66/A OR2X1_LOC_548/B 0.11fF
C45677 OR2X1_LOC_630/Y OR2X1_LOC_563/A 0.02fF
C45678 OR2X1_LOC_66/A OR2X1_LOC_389/a_8_216# 0.01fF
C45679 OR2X1_LOC_612/B OR2X1_LOC_71/A 0.01fF
C45680 OR2X1_LOC_51/Y AND2X1_LOC_464/A 0.03fF
C45681 OR2X1_LOC_3/Y OR2X1_LOC_377/a_36_216# 0.03fF
C45682 OR2X1_LOC_51/Y AND2X1_LOC_213/B 0.05fF
C45683 AND2X1_LOC_430/a_36_24# OR2X1_LOC_451/B 0.00fF
C45684 OR2X1_LOC_308/A OR2X1_LOC_307/B 0.88fF
C45685 OR2X1_LOC_368/a_8_216# AND2X1_LOC_476/Y 0.03fF
C45686 OR2X1_LOC_100/Y AND2X1_LOC_64/Y 0.17fF
C45687 OR2X1_LOC_46/A OR2X1_LOC_28/a_8_216# 0.42fF
C45688 OR2X1_LOC_809/B OR2X1_LOC_138/A 0.09fF
C45689 OR2X1_LOC_585/A OR2X1_LOC_599/a_8_216# 0.01fF
C45690 AND2X1_LOC_555/Y AND2X1_LOC_363/B 0.01fF
C45691 OR2X1_LOC_574/A OR2X1_LOC_446/B 5.68fF
C45692 OR2X1_LOC_624/A OR2X1_LOC_508/Y 0.05fF
C45693 AND2X1_LOC_141/a_8_24# OR2X1_LOC_595/A 0.01fF
C45694 OR2X1_LOC_851/A AND2X1_LOC_273/a_8_24# 0.01fF
C45695 OR2X1_LOC_715/B AND2X1_LOC_18/Y 0.10fF
C45696 OR2X1_LOC_528/Y OR2X1_LOC_604/A 0.07fF
C45697 OR2X1_LOC_186/Y AND2X1_LOC_92/Y 0.03fF
C45698 D_INPUT_3 OR2X1_LOC_619/a_36_216# 0.00fF
C45699 INPUT_0 OR2X1_LOC_161/B 0.47fF
C45700 AND2X1_LOC_543/Y AND2X1_LOC_717/Y 0.01fF
C45701 OR2X1_LOC_709/A OR2X1_LOC_715/A 0.01fF
C45702 AND2X1_LOC_3/Y OR2X1_LOC_707/a_8_216# 0.06fF
C45703 INPUT_2 OR2X1_LOC_14/a_8_216# 0.05fF
C45704 OR2X1_LOC_369/Y AND2X1_LOC_182/a_8_24# 0.01fF
C45705 OR2X1_LOC_643/A OR2X1_LOC_539/B 0.00fF
C45706 AND2X1_LOC_22/Y OR2X1_LOC_623/B 0.01fF
C45707 VDD OR2X1_LOC_461/B 0.21fF
C45708 OR2X1_LOC_721/a_8_216# OR2X1_LOC_721/Y 0.01fF
C45709 OR2X1_LOC_47/Y OR2X1_LOC_234/a_8_216# 0.05fF
C45710 AND2X1_LOC_7/Y AND2X1_LOC_52/Y 0.04fF
C45711 OR2X1_LOC_589/A INPUT_0 0.03fF
C45712 OR2X1_LOC_158/A AND2X1_LOC_858/B 0.01fF
C45713 OR2X1_LOC_158/A OR2X1_LOC_91/A 0.68fF
C45714 AND2X1_LOC_252/a_8_24# AND2X1_LOC_36/Y 0.01fF
C45715 OR2X1_LOC_296/Y OR2X1_LOC_777/B 0.03fF
C45716 AND2X1_LOC_738/B OR2X1_LOC_485/Y 0.02fF
C45717 OR2X1_LOC_329/Y AND2X1_LOC_434/Y 0.07fF
C45718 AND2X1_LOC_57/a_8_24# AND2X1_LOC_44/Y 0.03fF
C45719 OR2X1_LOC_481/A OR2X1_LOC_437/A 0.03fF
C45720 AND2X1_LOC_91/B OR2X1_LOC_377/A 0.07fF
C45721 AND2X1_LOC_22/Y OR2X1_LOC_794/A 0.02fF
C45722 OR2X1_LOC_493/A AND2X1_LOC_7/B 0.98fF
C45723 OR2X1_LOC_694/Y OR2X1_LOC_51/Y 0.01fF
C45724 AND2X1_LOC_716/Y AND2X1_LOC_364/a_36_24# 0.00fF
C45725 AND2X1_LOC_217/Y OR2X1_LOC_744/A 0.00fF
C45726 OR2X1_LOC_805/A OR2X1_LOC_831/B 0.07fF
C45727 OR2X1_LOC_40/Y AND2X1_LOC_675/Y 0.03fF
C45728 OR2X1_LOC_655/B OR2X1_LOC_68/B 0.03fF
C45729 OR2X1_LOC_768/A OR2X1_LOC_160/B 0.02fF
C45730 OR2X1_LOC_791/a_8_216# OR2X1_LOC_792/A 0.05fF
C45731 OR2X1_LOC_97/A OR2X1_LOC_661/a_8_216# 0.01fF
C45732 VDD OR2X1_LOC_778/B 0.05fF
C45733 AND2X1_LOC_541/a_36_24# OR2X1_LOC_65/B 0.00fF
C45734 AND2X1_LOC_153/a_36_24# OR2X1_LOC_831/B 0.01fF
C45735 OR2X1_LOC_114/B OR2X1_LOC_235/B 0.01fF
C45736 OR2X1_LOC_639/a_8_216# AND2X1_LOC_31/Y 0.01fF
C45737 AND2X1_LOC_848/Y AND2X1_LOC_284/a_8_24# 0.00fF
C45738 OR2X1_LOC_369/a_36_216# OR2X1_LOC_744/A 0.02fF
C45739 OR2X1_LOC_66/A AND2X1_LOC_245/a_36_24# 0.00fF
C45740 OR2X1_LOC_604/A AND2X1_LOC_512/Y 0.07fF
C45741 OR2X1_LOC_516/Y OR2X1_LOC_485/A 0.11fF
C45742 AND2X1_LOC_91/B OR2X1_LOC_203/Y 0.10fF
C45743 OR2X1_LOC_696/A AND2X1_LOC_645/A 0.00fF
C45744 AND2X1_LOC_721/Y OR2X1_LOC_237/Y 0.02fF
C45745 OR2X1_LOC_45/B OR2X1_LOC_32/B 0.01fF
C45746 OR2X1_LOC_199/a_8_216# AND2X1_LOC_43/B 0.04fF
C45747 AND2X1_LOC_70/Y OR2X1_LOC_501/B 0.01fF
C45748 OR2X1_LOC_52/B AND2X1_LOC_780/a_8_24# 0.04fF
C45749 OR2X1_LOC_619/Y OR2X1_LOC_12/Y 0.14fF
C45750 OR2X1_LOC_52/B OR2X1_LOC_171/Y 0.02fF
C45751 AND2X1_LOC_717/Y OR2X1_LOC_322/Y 0.13fF
C45752 AND2X1_LOC_704/a_8_24# OR2X1_LOC_427/A 0.01fF
C45753 OR2X1_LOC_531/Y AND2X1_LOC_663/A 0.25fF
C45754 OR2X1_LOC_269/B OR2X1_LOC_562/A 0.03fF
C45755 AND2X1_LOC_32/a_8_24# OR2X1_LOC_34/A 0.05fF
C45756 OR2X1_LOC_97/A OR2X1_LOC_462/B 0.03fF
C45757 OR2X1_LOC_240/A OR2X1_LOC_397/a_36_216# 0.01fF
C45758 OR2X1_LOC_687/Y AND2X1_LOC_44/Y 0.03fF
C45759 AND2X1_LOC_539/Y OR2X1_LOC_312/Y 0.07fF
C45760 OR2X1_LOC_541/B OR2X1_LOC_549/A 0.02fF
C45761 OR2X1_LOC_71/Y OR2X1_LOC_437/A 0.03fF
C45762 OR2X1_LOC_805/A OR2X1_LOC_344/A 0.03fF
C45763 AND2X1_LOC_727/A OR2X1_LOC_142/Y 0.07fF
C45764 OR2X1_LOC_426/B AND2X1_LOC_857/Y 0.03fF
C45765 D_INPUT_0 OR2X1_LOC_13/B 13.90fF
C45766 AND2X1_LOC_552/a_8_24# OR2X1_LOC_312/Y 0.01fF
C45767 OR2X1_LOC_122/a_36_216# AND2X1_LOC_474/A 0.00fF
C45768 AND2X1_LOC_716/Y AND2X1_LOC_326/B 0.00fF
C45769 AND2X1_LOC_40/Y OR2X1_LOC_468/A 0.11fF
C45770 OR2X1_LOC_158/A AND2X1_LOC_573/A 0.07fF
C45771 AND2X1_LOC_456/Y OR2X1_LOC_184/a_8_216# 0.14fF
C45772 OR2X1_LOC_821/a_8_216# OR2X1_LOC_85/A 0.15fF
C45773 AND2X1_LOC_98/Y OR2X1_LOC_91/A 0.01fF
C45774 OR2X1_LOC_364/A OR2X1_LOC_435/A 0.01fF
C45775 OR2X1_LOC_785/a_8_216# OR2X1_LOC_785/B 0.03fF
C45776 OR2X1_LOC_638/B D_INPUT_5 0.00fF
C45777 OR2X1_LOC_351/a_8_216# OR2X1_LOC_358/A 0.01fF
C45778 OR2X1_LOC_205/Y OR2X1_LOC_68/B 0.00fF
C45779 OR2X1_LOC_185/Y OR2X1_LOC_435/A 0.05fF
C45780 VDD AND2X1_LOC_527/a_8_24# 0.00fF
C45781 OR2X1_LOC_262/Y OR2X1_LOC_79/Y 0.03fF
C45782 AND2X1_LOC_216/A AND2X1_LOC_656/a_8_24# 0.22fF
C45783 AND2X1_LOC_807/B AND2X1_LOC_805/Y 0.03fF
C45784 OR2X1_LOC_673/a_36_216# OR2X1_LOC_375/A 0.02fF
C45785 OR2X1_LOC_833/Y AND2X1_LOC_56/B 0.01fF
C45786 OR2X1_LOC_600/A OR2X1_LOC_393/Y 0.03fF
C45787 OR2X1_LOC_264/a_8_216# AND2X1_LOC_65/A 0.05fF
C45788 VDD AND2X1_LOC_99/A 0.35fF
C45789 OR2X1_LOC_264/Y OR2X1_LOC_78/B 0.23fF
C45790 AND2X1_LOC_22/Y AND2X1_LOC_43/a_8_24# 0.04fF
C45791 AND2X1_LOC_57/Y OR2X1_LOC_19/B 0.02fF
C45792 VDD OR2X1_LOC_559/B 0.02fF
C45793 INPUT_0 AND2X1_LOC_654/B 0.03fF
C45794 OR2X1_LOC_742/B OR2X1_LOC_551/B 0.09fF
C45795 OR2X1_LOC_624/A OR2X1_LOC_66/A 1.04fF
C45796 AND2X1_LOC_41/A OR2X1_LOC_448/A 0.00fF
C45797 OR2X1_LOC_215/Y AND2X1_LOC_18/Y 0.03fF
C45798 OR2X1_LOC_620/B AND2X1_LOC_44/Y 0.23fF
C45799 OR2X1_LOC_45/B OR2X1_LOC_371/Y 0.01fF
C45800 AND2X1_LOC_13/a_8_24# AND2X1_LOC_7/B 0.08fF
C45801 OR2X1_LOC_95/Y OR2X1_LOC_142/Y 0.12fF
C45802 OR2X1_LOC_161/A OR2X1_LOC_347/Y 0.01fF
C45803 VDD OR2X1_LOC_639/B 0.12fF
C45804 AND2X1_LOC_639/B AND2X1_LOC_639/a_8_24# 0.03fF
C45805 OR2X1_LOC_696/A AND2X1_LOC_477/A 0.07fF
C45806 OR2X1_LOC_745/Y AND2X1_LOC_781/a_8_24# 0.23fF
C45807 OR2X1_LOC_185/A AND2X1_LOC_19/Y 0.03fF
C45808 OR2X1_LOC_703/A OR2X1_LOC_147/B 10.54fF
C45809 OR2X1_LOC_158/A OR2X1_LOC_669/Y 0.02fF
C45810 OR2X1_LOC_402/Y OR2X1_LOC_78/A 0.03fF
C45811 AND2X1_LOC_738/B OR2X1_LOC_39/A 0.10fF
C45812 OR2X1_LOC_421/A OR2X1_LOC_599/A 0.12fF
C45813 AND2X1_LOC_509/a_8_24# OR2X1_LOC_39/A 0.26fF
C45814 AND2X1_LOC_320/a_8_24# OR2X1_LOC_739/A 0.01fF
C45815 OR2X1_LOC_56/A OR2X1_LOC_39/A 0.22fF
C45816 OR2X1_LOC_405/A OR2X1_LOC_778/a_36_216# 0.00fF
C45817 VDD OR2X1_LOC_720/A -0.00fF
C45818 OR2X1_LOC_812/B OR2X1_LOC_561/Y 0.01fF
C45819 OR2X1_LOC_110/a_8_216# INPUT_1 0.03fF
C45820 OR2X1_LOC_814/A OR2X1_LOC_718/a_8_216# 0.03fF
C45821 OR2X1_LOC_600/A AND2X1_LOC_650/Y 1.46fF
C45822 AND2X1_LOC_212/Y AND2X1_LOC_211/a_8_24# 0.03fF
C45823 AND2X1_LOC_285/Y AND2X1_LOC_286/Y 0.00fF
C45824 AND2X1_LOC_392/A AND2X1_LOC_661/A 0.16fF
C45825 OR2X1_LOC_337/a_8_216# AND2X1_LOC_95/Y 0.04fF
C45826 AND2X1_LOC_794/A OR2X1_LOC_516/B 0.03fF
C45827 AND2X1_LOC_95/Y OR2X1_LOC_434/a_8_216# 0.01fF
C45828 AND2X1_LOC_553/a_36_24# OR2X1_LOC_26/Y 0.00fF
C45829 AND2X1_LOC_504/a_36_24# AND2X1_LOC_41/A 0.01fF
C45830 OR2X1_LOC_6/B OR2X1_LOC_37/a_8_216# 0.06fF
C45831 OR2X1_LOC_185/A AND2X1_LOC_189/a_36_24# 0.00fF
C45832 VDD OR2X1_LOC_627/a_8_216# 0.21fF
C45833 OR2X1_LOC_493/Y OR2X1_LOC_561/A 0.10fF
C45834 VDD AND2X1_LOC_637/Y 0.01fF
C45835 OR2X1_LOC_604/A OR2X1_LOC_682/Y 0.00fF
C45836 OR2X1_LOC_160/A OR2X1_LOC_735/a_8_216# 0.04fF
C45837 AND2X1_LOC_64/Y OR2X1_LOC_532/B 1.11fF
C45838 AND2X1_LOC_92/Y OR2X1_LOC_358/B 0.01fF
C45839 AND2X1_LOC_794/B OR2X1_LOC_417/a_8_216# 0.06fF
C45840 OR2X1_LOC_134/a_8_216# OR2X1_LOC_95/Y 0.03fF
C45841 OR2X1_LOC_306/Y AND2X1_LOC_512/Y 0.00fF
C45842 AND2X1_LOC_373/a_8_24# VDD 0.00fF
C45843 AND2X1_LOC_64/Y AND2X1_LOC_665/a_8_24# 0.01fF
C45844 OR2X1_LOC_8/Y AND2X1_LOC_342/a_36_24# 0.00fF
C45845 AND2X1_LOC_779/a_8_24# OR2X1_LOC_427/A 0.02fF
C45846 AND2X1_LOC_228/Y OR2X1_LOC_298/a_8_216# 0.01fF
C45847 OR2X1_LOC_744/A AND2X1_LOC_359/B 0.14fF
C45848 OR2X1_LOC_158/A OR2X1_LOC_27/Y 0.03fF
C45849 AND2X1_LOC_729/Y OR2X1_LOC_441/Y 0.03fF
C45850 OR2X1_LOC_158/A AND2X1_LOC_662/a_8_24# 0.04fF
C45851 OR2X1_LOC_333/B VDD 0.11fF
C45852 OR2X1_LOC_848/B OR2X1_LOC_391/a_8_216# 0.04fF
C45853 INPUT_0 OR2X1_LOC_43/A 0.63fF
C45854 OR2X1_LOC_666/Y AND2X1_LOC_658/A 0.40fF
C45855 OR2X1_LOC_589/A OR2X1_LOC_64/Y 0.14fF
C45856 OR2X1_LOC_653/Y AND2X1_LOC_95/Y 0.01fF
C45857 AND2X1_LOC_367/A OR2X1_LOC_44/Y 0.10fF
C45858 AND2X1_LOC_211/B OR2X1_LOC_56/A 0.07fF
C45859 OR2X1_LOC_43/a_8_216# OR2X1_LOC_13/Y 0.01fF
C45860 OR2X1_LOC_264/Y OR2X1_LOC_375/A 0.12fF
C45861 OR2X1_LOC_377/A AND2X1_LOC_39/a_36_24# 0.00fF
C45862 AND2X1_LOC_718/a_8_24# OR2X1_LOC_36/Y 0.00fF
C45863 AND2X1_LOC_92/a_36_24# INPUT_1 0.00fF
C45864 OR2X1_LOC_831/A OR2X1_LOC_121/B 0.02fF
C45865 OR2X1_LOC_311/Y OR2X1_LOC_13/a_8_216# 0.01fF
C45866 AND2X1_LOC_70/Y AND2X1_LOC_387/B 0.03fF
C45867 OR2X1_LOC_848/A OR2X1_LOC_391/a_36_216# 0.01fF
C45868 AND2X1_LOC_95/Y OR2X1_LOC_833/B 0.02fF
C45869 AND2X1_LOC_784/A AND2X1_LOC_335/a_8_24# 0.03fF
C45870 AND2X1_LOC_559/a_8_24# OR2X1_LOC_517/A 0.01fF
C45871 OR2X1_LOC_848/A OR2X1_LOC_489/a_8_216# 0.02fF
C45872 AND2X1_LOC_390/B AND2X1_LOC_436/Y 0.02fF
C45873 AND2X1_LOC_560/B OR2X1_LOC_275/Y 0.01fF
C45874 OR2X1_LOC_640/A AND2X1_LOC_89/a_8_24# 0.08fF
C45875 OR2X1_LOC_840/A OR2X1_LOC_87/A 0.14fF
C45876 OR2X1_LOC_599/A AND2X1_LOC_718/a_36_24# 0.01fF
C45877 AND2X1_LOC_47/Y AND2X1_LOC_248/a_8_24# 0.04fF
C45878 AND2X1_LOC_486/Y OR2X1_LOC_497/a_8_216# 0.23fF
C45879 AND2X1_LOC_850/Y OR2X1_LOC_39/A 0.01fF
C45880 AND2X1_LOC_3/Y OR2X1_LOC_630/B 0.02fF
C45881 OR2X1_LOC_493/A OR2X1_LOC_805/A 0.15fF
C45882 OR2X1_LOC_165/a_8_216# OR2X1_LOC_91/Y 0.05fF
C45883 OR2X1_LOC_240/B OR2X1_LOC_243/A 0.05fF
C45884 OR2X1_LOC_643/A OR2X1_LOC_721/Y 0.03fF
C45885 OR2X1_LOC_647/A OR2X1_LOC_78/B 0.06fF
C45886 AND2X1_LOC_556/a_8_24# OR2X1_LOC_7/A 0.04fF
C45887 AND2X1_LOC_82/Y OR2X1_LOC_532/B 0.00fF
C45888 OR2X1_LOC_604/A AND2X1_LOC_712/B 0.03fF
C45889 VDD OR2X1_LOC_99/B 0.18fF
C45890 AND2X1_LOC_668/a_8_24# OR2X1_LOC_278/Y 0.01fF
C45891 OR2X1_LOC_235/B AND2X1_LOC_79/Y 0.07fF
C45892 OR2X1_LOC_756/B AND2X1_LOC_85/a_8_24# 0.20fF
C45893 AND2X1_LOC_95/Y OR2X1_LOC_254/B 0.07fF
C45894 AND2X1_LOC_40/Y OR2X1_LOC_449/B 0.03fF
C45895 OR2X1_LOC_404/Y OR2X1_LOC_244/Y 0.43fF
C45896 AND2X1_LOC_337/a_8_24# OR2X1_LOC_64/Y 0.01fF
C45897 OR2X1_LOC_485/A AND2X1_LOC_842/a_8_24# 0.01fF
C45898 OR2X1_LOC_604/A OR2X1_LOC_54/Y 0.20fF
C45899 OR2X1_LOC_671/Y OR2X1_LOC_54/a_8_216# 0.02fF
C45900 OR2X1_LOC_159/a_36_216# OR2X1_LOC_46/A 0.00fF
C45901 AND2X1_LOC_720/Y OR2X1_LOC_669/Y 0.03fF
C45902 OR2X1_LOC_47/Y OR2X1_LOC_312/a_8_216# 0.01fF
C45903 OR2X1_LOC_450/Y AND2X1_LOC_425/Y 0.02fF
C45904 VDD OR2X1_LOC_65/Y 0.06fF
C45905 OR2X1_LOC_161/A OR2X1_LOC_668/Y 0.12fF
C45906 OR2X1_LOC_814/A OR2X1_LOC_362/A 0.02fF
C45907 AND2X1_LOC_729/Y AND2X1_LOC_436/B 0.03fF
C45908 OR2X1_LOC_329/B AND2X1_LOC_473/a_36_24# 0.00fF
C45909 OR2X1_LOC_634/A AND2X1_LOC_42/B 0.00fF
C45910 OR2X1_LOC_456/Y OR2X1_LOC_456/a_8_216# 0.01fF
C45911 AND2X1_LOC_70/a_8_24# AND2X1_LOC_51/Y 0.04fF
C45912 OR2X1_LOC_756/B OR2X1_LOC_33/B 0.01fF
C45913 OR2X1_LOC_54/Y OR2X1_LOC_66/A 0.03fF
C45914 OR2X1_LOC_743/A AND2X1_LOC_857/Y 0.03fF
C45915 OR2X1_LOC_313/Y AND2X1_LOC_317/a_8_24# 0.24fF
C45916 OR2X1_LOC_786/Y AND2X1_LOC_44/Y 0.03fF
C45917 AND2X1_LOC_650/Y OR2X1_LOC_619/Y 0.05fF
C45918 OR2X1_LOC_121/Y OR2X1_LOC_276/B 0.02fF
C45919 OR2X1_LOC_295/a_8_216# OR2X1_LOC_59/Y 0.09fF
C45920 AND2X1_LOC_36/Y OR2X1_LOC_724/A 0.17fF
C45921 OR2X1_LOC_744/A AND2X1_LOC_802/a_8_24# 0.01fF
C45922 AND2X1_LOC_379/a_8_24# OR2X1_LOC_11/Y 0.01fF
C45923 AND2X1_LOC_784/A OR2X1_LOC_519/Y 0.01fF
C45924 OR2X1_LOC_635/A AND2X1_LOC_683/a_36_24# 0.01fF
C45925 OR2X1_LOC_3/Y OR2X1_LOC_502/A 0.03fF
C45926 AND2X1_LOC_56/B OR2X1_LOC_39/A 3.56fF
C45927 AND2X1_LOC_145/a_8_24# OR2X1_LOC_87/A 0.05fF
C45928 OR2X1_LOC_836/A AND2X1_LOC_824/a_8_24# 0.02fF
C45929 AND2X1_LOC_741/Y AND2X1_LOC_480/a_36_24# 0.00fF
C45930 OR2X1_LOC_18/Y OR2X1_LOC_24/a_8_216# 0.01fF
C45931 AND2X1_LOC_48/A OR2X1_LOC_520/a_8_216# 0.01fF
C45932 OR2X1_LOC_335/Y OR2X1_LOC_121/B 0.01fF
C45933 OR2X1_LOC_631/a_8_216# OR2X1_LOC_574/A 0.03fF
C45934 OR2X1_LOC_447/Y OR2X1_LOC_66/A 0.03fF
C45935 OR2X1_LOC_689/Y AND2X1_LOC_194/Y 0.02fF
C45936 VDD OR2X1_LOC_443/a_8_216# 0.00fF
C45937 OR2X1_LOC_643/A OR2X1_LOC_375/A 0.03fF
C45938 AND2X1_LOC_35/Y OR2X1_LOC_44/Y 0.07fF
C45939 AND2X1_LOC_44/Y OR2X1_LOC_644/A 0.09fF
C45940 OR2X1_LOC_375/A OR2X1_LOC_124/Y 0.01fF
C45941 AND2X1_LOC_796/a_36_24# AND2X1_LOC_810/Y 0.00fF
C45942 OR2X1_LOC_375/A OR2X1_LOC_778/Y 0.13fF
C45943 AND2X1_LOC_76/Y AND2X1_LOC_276/Y 0.39fF
C45944 AND2X1_LOC_107/a_36_24# OR2X1_LOC_78/A 0.01fF
C45945 OR2X1_LOC_6/B OR2X1_LOC_62/A 0.73fF
C45946 AND2X1_LOC_392/A AND2X1_LOC_810/Y 0.07fF
C45947 AND2X1_LOC_553/A AND2X1_LOC_523/Y 0.14fF
C45948 OR2X1_LOC_308/Y AND2X1_LOC_419/a_36_24# -0.02fF
C45949 OR2X1_LOC_472/A OR2X1_LOC_375/A 0.27fF
C45950 OR2X1_LOC_64/Y AND2X1_LOC_654/B 0.01fF
C45951 AND2X1_LOC_862/a_36_24# AND2X1_LOC_807/Y 0.05fF
C45952 OR2X1_LOC_856/B OR2X1_LOC_193/A 0.02fF
C45953 AND2X1_LOC_347/a_8_24# AND2X1_LOC_847/Y 0.02fF
C45954 AND2X1_LOC_218/a_8_24# AND2X1_LOC_660/A 0.02fF
C45955 AND2X1_LOC_40/Y OR2X1_LOC_121/B 0.09fF
C45956 OR2X1_LOC_36/Y OR2X1_LOC_26/Y 1.71fF
C45957 OR2X1_LOC_64/Y OR2X1_LOC_495/Y 0.11fF
C45958 AND2X1_LOC_857/Y OR2X1_LOC_246/A 0.00fF
C45959 OR2X1_LOC_615/a_8_216# OR2X1_LOC_427/A 0.01fF
C45960 OR2X1_LOC_756/B OR2X1_LOC_287/a_8_216# 0.02fF
C45961 OR2X1_LOC_160/A OR2X1_LOC_479/Y 0.10fF
C45962 OR2X1_LOC_557/A OR2X1_LOC_404/a_36_216# 0.00fF
C45963 OR2X1_LOC_154/A OR2X1_LOC_654/A 0.07fF
C45964 AND2X1_LOC_314/a_8_24# AND2X1_LOC_51/Y 0.02fF
C45965 OR2X1_LOC_45/B AND2X1_LOC_222/Y 0.01fF
C45966 OR2X1_LOC_43/A OR2X1_LOC_690/A 0.77fF
C45967 AND2X1_LOC_41/A AND2X1_LOC_7/Y 0.03fF
C45968 AND2X1_LOC_228/Y OR2X1_LOC_229/Y 0.01fF
C45969 OR2X1_LOC_36/Y AND2X1_LOC_493/a_8_24# 0.01fF
C45970 AND2X1_LOC_88/a_8_24# OR2X1_LOC_87/Y 0.11fF
C45971 OR2X1_LOC_703/A OR2X1_LOC_545/B 0.05fF
C45972 OR2X1_LOC_44/Y OR2X1_LOC_757/a_8_216# 0.01fF
C45973 OR2X1_LOC_574/A AND2X1_LOC_56/B 0.10fF
C45974 INPUT_1 AND2X1_LOC_401/Y 0.05fF
C45975 AND2X1_LOC_854/a_8_24# AND2X1_LOC_856/A 0.00fF
C45976 OR2X1_LOC_793/A OR2X1_LOC_793/B 0.00fF
C45977 OR2X1_LOC_36/Y OR2X1_LOC_89/A 0.12fF
C45978 OR2X1_LOC_356/A OR2X1_LOC_365/B 0.05fF
C45979 AND2X1_LOC_456/Y OR2X1_LOC_44/Y 0.01fF
C45980 AND2X1_LOC_56/B OR2X1_LOC_33/A 0.04fF
C45981 AND2X1_LOC_474/A AND2X1_LOC_859/B 0.01fF
C45982 OR2X1_LOC_736/Y OR2X1_LOC_675/Y 0.04fF
C45983 OR2X1_LOC_795/a_8_216# OR2X1_LOC_776/Y -0.00fF
C45984 OR2X1_LOC_405/A OR2X1_LOC_476/B 0.10fF
C45985 OR2X1_LOC_464/A OR2X1_LOC_532/B 0.04fF
C45986 OR2X1_LOC_74/A OR2X1_LOC_44/Y 0.07fF
C45987 OR2X1_LOC_748/A OR2X1_LOC_817/a_8_216# 0.01fF
C45988 AND2X1_LOC_191/Y AND2X1_LOC_580/B 0.03fF
C45989 OR2X1_LOC_502/A AND2X1_LOC_53/Y 0.01fF
C45990 OR2X1_LOC_272/a_8_216# OR2X1_LOC_43/A 0.06fF
C45991 OR2X1_LOC_154/A AND2X1_LOC_496/a_36_24# 0.06fF
C45992 AND2X1_LOC_365/A OR2X1_LOC_64/Y 0.59fF
C45993 AND2X1_LOC_91/B OR2X1_LOC_732/A 1.55fF
C45994 OR2X1_LOC_615/Y AND2X1_LOC_663/A 0.03fF
C45995 OR2X1_LOC_404/Y AND2X1_LOC_669/a_8_24# 0.01fF
C45996 AND2X1_LOC_711/Y AND2X1_LOC_580/B 0.03fF
C45997 INPUT_3 OR2X1_LOC_46/A 0.03fF
C45998 OR2X1_LOC_856/B D_INPUT_0 0.12fF
C45999 AND2X1_LOC_379/a_8_24# OR2X1_LOC_64/Y 0.01fF
C46000 AND2X1_LOC_31/Y OR2X1_LOC_486/Y 14.74fF
C46001 AND2X1_LOC_348/Y OR2X1_LOC_481/A 0.08fF
C46002 OR2X1_LOC_495/Y OR2X1_LOC_417/A 0.03fF
C46003 AND2X1_LOC_539/Y OR2X1_LOC_13/B 0.12fF
C46004 AND2X1_LOC_276/Y OR2X1_LOC_52/B 0.05fF
C46005 OR2X1_LOC_185/A AND2X1_LOC_309/a_8_24# 0.00fF
C46006 OR2X1_LOC_45/B OR2X1_LOC_423/Y 0.03fF
C46007 OR2X1_LOC_121/B OR2X1_LOC_87/Y 0.00fF
C46008 OR2X1_LOC_261/A OR2X1_LOC_44/Y 0.00fF
C46009 OR2X1_LOC_481/A OR2X1_LOC_753/A 0.01fF
C46010 AND2X1_LOC_211/B AND2X1_LOC_641/Y 0.01fF
C46011 VDD OR2X1_LOC_590/a_8_216# 0.00fF
C46012 OR2X1_LOC_62/B AND2X1_LOC_43/B 0.00fF
C46013 OR2X1_LOC_851/B OR2X1_LOC_68/B 0.34fF
C46014 AND2X1_LOC_86/B AND2X1_LOC_38/a_8_24# 0.20fF
C46015 OR2X1_LOC_43/A OR2X1_LOC_64/Y 0.19fF
C46016 OR2X1_LOC_91/Y OR2X1_LOC_22/Y 0.07fF
C46017 AND2X1_LOC_554/B OR2X1_LOC_131/Y 0.17fF
C46018 OR2X1_LOC_576/A OR2X1_LOC_140/Y 0.00fF
C46019 AND2X1_LOC_99/A OR2X1_LOC_256/A 0.03fF
C46020 AND2X1_LOC_70/Y OR2X1_LOC_318/B 0.03fF
C46021 AND2X1_LOC_18/Y OR2X1_LOC_398/Y 0.00fF
C46022 AND2X1_LOC_72/B OR2X1_LOC_632/Y 0.05fF
C46023 OR2X1_LOC_680/Y AND2X1_LOC_728/a_8_24# 0.11fF
C46024 OR2X1_LOC_160/B OR2X1_LOC_641/B 0.02fF
C46025 AND2X1_LOC_36/Y OR2X1_LOC_415/Y 0.00fF
C46026 OR2X1_LOC_115/B OR2X1_LOC_844/B 0.17fF
C46027 VDD OR2X1_LOC_160/a_8_216# 0.00fF
C46028 AND2X1_LOC_822/a_8_24# AND2X1_LOC_51/Y 0.01fF
C46029 VDD OR2X1_LOC_72/Y 0.22fF
C46030 OR2X1_LOC_95/Y OR2X1_LOC_118/Y 0.03fF
C46031 OR2X1_LOC_644/B AND2X1_LOC_48/A 0.00fF
C46032 OR2X1_LOC_214/a_8_216# OR2X1_LOC_750/A 0.03fF
C46033 AND2X1_LOC_449/a_8_24# OR2X1_LOC_428/A 0.01fF
C46034 OR2X1_LOC_604/a_36_216# AND2X1_LOC_452/Y 0.01fF
C46035 AND2X1_LOC_8/Y AND2X1_LOC_672/B 0.90fF
C46036 OR2X1_LOC_756/B OR2X1_LOC_374/Y 0.04fF
C46037 AND2X1_LOC_554/Y D_INPUT_3 0.02fF
C46038 OR2X1_LOC_492/Y OR2X1_LOC_437/A 0.02fF
C46039 AND2X1_LOC_356/B OR2X1_LOC_311/Y 0.01fF
C46040 OR2X1_LOC_835/Y OR2X1_LOC_269/B 0.34fF
C46041 AND2X1_LOC_12/Y OR2X1_LOC_276/B 0.09fF
C46042 AND2X1_LOC_525/a_36_24# AND2X1_LOC_51/Y 0.01fF
C46043 OR2X1_LOC_837/A AND2X1_LOC_461/a_8_24# 0.08fF
C46044 OR2X1_LOC_436/Y OR2X1_LOC_798/a_8_216# 0.16fF
C46045 OR2X1_LOC_43/A OR2X1_LOC_417/A 0.07fF
C46046 OR2X1_LOC_743/A AND2X1_LOC_685/a_36_24# 0.00fF
C46047 OR2X1_LOC_461/Y OR2X1_LOC_462/a_8_216# 0.39fF
C46048 AND2X1_LOC_68/a_8_24# OR2X1_LOC_52/B -0.00fF
C46049 AND2X1_LOC_187/a_8_24# AND2X1_LOC_441/a_8_24# 0.23fF
C46050 OR2X1_LOC_475/Y OR2X1_LOC_121/B 0.01fF
C46051 OR2X1_LOC_441/a_36_216# AND2X1_LOC_222/Y 0.00fF
C46052 AND2X1_LOC_99/A OR2X1_LOC_67/Y 0.22fF
C46053 OR2X1_LOC_557/A OR2X1_LOC_404/A 0.01fF
C46054 AND2X1_LOC_75/a_8_24# OR2X1_LOC_76/A 0.10fF
C46055 OR2X1_LOC_321/Y OR2X1_LOC_46/A 0.03fF
C46056 AND2X1_LOC_51/Y AND2X1_LOC_816/a_8_24# 0.01fF
C46057 OR2X1_LOC_190/A OR2X1_LOC_366/Y 3.27fF
C46058 AND2X1_LOC_110/Y OR2X1_LOC_112/A 0.00fF
C46059 OR2X1_LOC_502/A AND2X1_LOC_609/a_8_24# 0.01fF
C46060 OR2X1_LOC_696/A AND2X1_LOC_703/Y 0.00fF
C46061 OR2X1_LOC_64/Y AND2X1_LOC_685/a_8_24# 0.01fF
C46062 D_INPUT_5 AND2X1_LOC_430/B 0.01fF
C46063 OR2X1_LOC_426/B OR2X1_LOC_437/A 0.75fF
C46064 OR2X1_LOC_95/Y OR2X1_LOC_238/Y 0.03fF
C46065 AND2X1_LOC_178/a_36_24# OR2X1_LOC_192/B 0.00fF
C46066 AND2X1_LOC_326/A AND2X1_LOC_326/a_8_24# 0.10fF
C46067 AND2X1_LOC_351/Y AND2X1_LOC_358/a_8_24# 0.00fF
C46068 OR2X1_LOC_859/A AND2X1_LOC_51/Y 0.12fF
C46069 AND2X1_LOC_52/a_8_24# OR2X1_LOC_198/A 0.23fF
C46070 OR2X1_LOC_862/A OR2X1_LOC_561/B 0.67fF
C46071 OR2X1_LOC_31/Y AND2X1_LOC_639/a_8_24# 0.01fF
C46072 OR2X1_LOC_474/a_8_216# OR2X1_LOC_849/a_8_216# 0.47fF
C46073 OR2X1_LOC_291/Y OR2X1_LOC_22/Y 0.12fF
C46074 OR2X1_LOC_502/A AND2X1_LOC_409/a_8_24# 0.01fF
C46075 OR2X1_LOC_311/Y OR2X1_LOC_22/Y 1.36fF
C46076 OR2X1_LOC_753/A D_INPUT_1 0.03fF
C46077 OR2X1_LOC_36/Y OR2X1_LOC_419/a_8_216# 0.07fF
C46078 AND2X1_LOC_715/Y AND2X1_LOC_703/Y 0.02fF
C46079 OR2X1_LOC_304/a_8_216# OR2X1_LOC_428/A 0.02fF
C46080 OR2X1_LOC_276/B AND2X1_LOC_496/a_8_24# 0.01fF
C46081 AND2X1_LOC_538/Y OR2X1_LOC_22/Y 0.01fF
C46082 OR2X1_LOC_231/a_8_216# AND2X1_LOC_31/Y 0.01fF
C46083 OR2X1_LOC_627/a_8_216# AND2X1_LOC_624/B 0.01fF
C46084 AND2X1_LOC_616/a_8_24# AND2X1_LOC_36/Y 0.01fF
C46085 OR2X1_LOC_206/A OR2X1_LOC_532/B 0.03fF
C46086 OR2X1_LOC_268/a_8_216# INPUT_1 0.03fF
C46087 AND2X1_LOC_7/B OR2X1_LOC_161/B 0.64fF
C46088 AND2X1_LOC_12/Y AND2X1_LOC_430/B 0.01fF
C46089 AND2X1_LOC_12/Y OR2X1_LOC_779/B 0.05fF
C46090 AND2X1_LOC_712/a_8_24# OR2X1_LOC_428/A 0.01fF
C46091 OR2X1_LOC_26/Y OR2X1_LOC_419/Y 0.14fF
C46092 OR2X1_LOC_152/Y AND2X1_LOC_808/A 0.22fF
C46093 OR2X1_LOC_48/Y OR2X1_LOC_47/Y 0.00fF
C46094 OR2X1_LOC_78/A OR2X1_LOC_593/B 0.01fF
C46095 AND2X1_LOC_48/A AND2X1_LOC_53/Y 0.02fF
C46096 OR2X1_LOC_160/A OR2X1_LOC_68/B 0.62fF
C46097 AND2X1_LOC_243/a_8_24# D_INPUT_1 0.17fF
C46098 OR2X1_LOC_12/Y AND2X1_LOC_769/Y 0.03fF
C46099 OR2X1_LOC_278/Y OR2X1_LOC_71/A 0.17fF
C46100 OR2X1_LOC_755/Y AND2X1_LOC_789/Y 0.04fF
C46101 OR2X1_LOC_89/A OR2X1_LOC_419/Y 1.28fF
C46102 OR2X1_LOC_16/A AND2X1_LOC_774/A 0.07fF
C46103 OR2X1_LOC_111/a_8_216# AND2X1_LOC_326/B 0.01fF
C46104 OR2X1_LOC_833/B OR2X1_LOC_269/A 0.17fF
C46105 AND2X1_LOC_424/a_8_24# OR2X1_LOC_712/B 0.01fF
C46106 OR2X1_LOC_344/A OR2X1_LOC_580/B 0.01fF
C46107 OR2X1_LOC_433/Y OR2X1_LOC_589/Y 0.10fF
C46108 OR2X1_LOC_44/Y AND2X1_LOC_783/a_8_24# 0.17fF
C46109 OR2X1_LOC_97/A OR2X1_LOC_661/A 0.01fF
C46110 OR2X1_LOC_756/B OR2X1_LOC_333/A 0.01fF
C46111 AND2X1_LOC_785/a_8_24# OR2X1_LOC_56/A 0.01fF
C46112 AND2X1_LOC_729/B OR2X1_LOC_311/a_8_216# 0.01fF
C46113 OR2X1_LOC_2/Y D_INPUT_6 0.59fF
C46114 OR2X1_LOC_373/Y AND2X1_LOC_778/Y 0.07fF
C46115 AND2X1_LOC_456/Y AND2X1_LOC_570/a_8_24# 0.02fF
C46116 OR2X1_LOC_673/B OR2X1_LOC_621/B 0.94fF
C46117 AND2X1_LOC_738/B AND2X1_LOC_564/A 0.12fF
C46118 AND2X1_LOC_91/B OR2X1_LOC_78/B 0.17fF
C46119 OR2X1_LOC_97/A OR2X1_LOC_602/Y 0.01fF
C46120 AND2X1_LOC_707/Y AND2X1_LOC_454/a_8_24# 0.07fF
C46121 OR2X1_LOC_720/B OR2X1_LOC_786/Y 0.00fF
C46122 OR2X1_LOC_185/A OR2X1_LOC_723/B 0.11fF
C46123 OR2X1_LOC_687/a_8_216# OR2X1_LOC_451/B 0.01fF
C46124 OR2X1_LOC_480/a_8_216# OR2X1_LOC_467/A 0.01fF
C46125 OR2X1_LOC_89/A OR2X1_LOC_152/A 0.14fF
C46126 AND2X1_LOC_338/Y OR2X1_LOC_51/Y 0.01fF
C46127 OR2X1_LOC_805/A OR2X1_LOC_332/a_8_216# 0.02fF
C46128 AND2X1_LOC_372/a_8_24# OR2X1_LOC_831/B 0.05fF
C46129 OR2X1_LOC_62/A AND2X1_LOC_47/Y 0.04fF
C46130 AND2X1_LOC_554/B AND2X1_LOC_657/A 0.02fF
C46131 AND2X1_LOC_65/A OR2X1_LOC_641/A 0.08fF
C46132 OR2X1_LOC_840/A OR2X1_LOC_390/B 0.10fF
C46133 OR2X1_LOC_46/A AND2X1_LOC_646/a_36_24# 0.00fF
C46134 OR2X1_LOC_830/a_8_216# OR2X1_LOC_294/Y 0.01fF
C46135 OR2X1_LOC_114/B AND2X1_LOC_295/a_8_24# 0.01fF
C46136 OR2X1_LOC_622/a_8_216# OR2X1_LOC_80/A 0.01fF
C46137 OR2X1_LOC_40/Y AND2X1_LOC_443/a_8_24# 0.03fF
C46138 OR2X1_LOC_856/a_36_216# OR2X1_LOC_198/A 0.02fF
C46139 OR2X1_LOC_61/A OR2X1_LOC_648/A 0.03fF
C46140 AND2X1_LOC_51/Y OR2X1_LOC_568/a_8_216# 0.06fF
C46141 OR2X1_LOC_756/B OR2X1_LOC_392/B 0.05fF
C46142 OR2X1_LOC_121/Y AND2X1_LOC_70/Y 0.09fF
C46143 OR2X1_LOC_510/A OR2X1_LOC_641/A 0.03fF
C46144 OR2X1_LOC_208/A OR2X1_LOC_856/B 0.05fF
C46145 OR2X1_LOC_6/B OR2X1_LOC_629/B 0.03fF
C46146 OR2X1_LOC_604/A OR2X1_LOC_765/Y 0.01fF
C46147 OR2X1_LOC_45/B AND2X1_LOC_367/A 0.05fF
C46148 OR2X1_LOC_421/A OR2X1_LOC_40/Y 0.03fF
C46149 AND2X1_LOC_22/Y OR2X1_LOC_434/a_8_216# 0.02fF
C46150 AND2X1_LOC_64/Y OR2X1_LOC_714/Y 0.01fF
C46151 AND2X1_LOC_22/Y OR2X1_LOC_776/a_8_216# 0.01fF
C46152 OR2X1_LOC_833/Y AND2X1_LOC_92/Y 0.01fF
C46153 OR2X1_LOC_808/B OR2X1_LOC_779/A 0.02fF
C46154 OR2X1_LOC_834/A OR2X1_LOC_713/A 0.01fF
C46155 OR2X1_LOC_263/a_36_216# AND2X1_LOC_647/Y 0.00fF
C46156 AND2X1_LOC_41/A OR2X1_LOC_706/a_8_216# 0.01fF
C46157 OR2X1_LOC_743/A OR2X1_LOC_437/A 0.07fF
C46158 OR2X1_LOC_134/Y OR2X1_LOC_427/A 0.01fF
C46159 OR2X1_LOC_8/Y OR2X1_LOC_6/B 3.36fF
C46160 AND2X1_LOC_82/Y OR2X1_LOC_78/a_36_216# 0.00fF
C46161 OR2X1_LOC_335/A OR2X1_LOC_185/A 0.71fF
C46162 OR2X1_LOC_244/Y OR2X1_LOC_362/A 0.03fF
C46163 OR2X1_LOC_533/Y AND2X1_LOC_512/Y 0.08fF
C46164 OR2X1_LOC_61/Y AND2X1_LOC_7/B 0.26fF
C46165 AND2X1_LOC_41/A OR2X1_LOC_390/A 0.03fF
C46166 OR2X1_LOC_319/B OR2X1_LOC_161/B 0.61fF
C46167 OR2X1_LOC_482/Y AND2X1_LOC_858/B 0.07fF
C46168 OR2X1_LOC_155/A OR2X1_LOC_593/B 0.55fF
C46169 AND2X1_LOC_22/Y OR2X1_LOC_653/Y 0.07fF
C46170 OR2X1_LOC_364/A OR2X1_LOC_605/Y 0.01fF
C46171 OR2X1_LOC_528/Y AND2X1_LOC_549/a_8_24# 0.04fF
C46172 OR2X1_LOC_725/B AND2X1_LOC_44/Y 0.01fF
C46173 OR2X1_LOC_426/B AND2X1_LOC_715/A 0.07fF
C46174 AND2X1_LOC_536/a_8_24# AND2X1_LOC_7/B 0.04fF
C46175 OR2X1_LOC_68/a_8_216# OR2X1_LOC_776/A 0.61fF
C46176 OR2X1_LOC_19/B OR2X1_LOC_71/A 0.08fF
C46177 AND2X1_LOC_387/a_8_24# AND2X1_LOC_92/Y 0.08fF
C46178 OR2X1_LOC_318/Y OR2X1_LOC_161/B 0.00fF
C46179 OR2X1_LOC_840/a_8_216# OR2X1_LOC_840/A 0.05fF
C46180 AND2X1_LOC_91/B OR2X1_LOC_375/A 0.43fF
C46181 OR2X1_LOC_178/a_8_216# OR2X1_LOC_744/A -0.01fF
C46182 OR2X1_LOC_641/a_36_216# AND2X1_LOC_92/Y 0.00fF
C46183 OR2X1_LOC_528/Y AND2X1_LOC_506/a_8_24# 0.26fF
C46184 AND2X1_LOC_721/Y AND2X1_LOC_573/A 0.02fF
C46185 OR2X1_LOC_220/B AND2X1_LOC_44/Y 0.02fF
C46186 AND2X1_LOC_596/a_36_24# OR2X1_LOC_744/A 0.00fF
C46187 OR2X1_LOC_264/Y OR2X1_LOC_549/A 0.14fF
C46188 AND2X1_LOC_811/Y AND2X1_LOC_222/Y 0.01fF
C46189 OR2X1_LOC_479/Y OR2X1_LOC_212/B 0.03fF
C46190 OR2X1_LOC_330/Y OR2X1_LOC_151/A 0.04fF
C46191 OR2X1_LOC_744/A AND2X1_LOC_436/Y 0.04fF
C46192 AND2X1_LOC_707/Y AND2X1_LOC_449/Y 0.01fF
C46193 OR2X1_LOC_417/A OR2X1_LOC_384/a_8_216# 0.05fF
C46194 OR2X1_LOC_604/A AND2X1_LOC_718/a_8_24# 0.17fF
C46195 OR2X1_LOC_246/A OR2X1_LOC_437/A 0.10fF
C46196 OR2X1_LOC_26/Y AND2X1_LOC_590/a_36_24# 0.01fF
C46197 OR2X1_LOC_419/a_8_216# OR2X1_LOC_419/Y 0.01fF
C46198 AND2X1_LOC_861/B AND2X1_LOC_807/B 0.52fF
C46199 AND2X1_LOC_40/Y OR2X1_LOC_621/B 0.23fF
C46200 VDD OR2X1_LOC_697/Y 0.32fF
C46201 AND2X1_LOC_70/Y OR2X1_LOC_538/A 0.04fF
C46202 OR2X1_LOC_155/A AND2X1_LOC_273/a_8_24# 0.12fF
C46203 AND2X1_LOC_109/a_8_24# AND2X1_LOC_31/Y 0.06fF
C46204 OR2X1_LOC_45/B AND2X1_LOC_35/Y 0.15fF
C46205 AND2X1_LOC_675/Y OR2X1_LOC_531/Y 0.07fF
C46206 AND2X1_LOC_474/A OR2X1_LOC_56/A 0.03fF
C46207 AND2X1_LOC_56/B OR2X1_LOC_855/A 0.03fF
C46208 OR2X1_LOC_805/A OR2X1_LOC_161/B 0.21fF
C46209 OR2X1_LOC_630/Y OR2X1_LOC_632/Y 0.03fF
C46210 AND2X1_LOC_789/a_8_24# OR2X1_LOC_600/A 0.01fF
C46211 OR2X1_LOC_709/A AND2X1_LOC_12/Y 0.01fF
C46212 OR2X1_LOC_804/a_8_216# AND2X1_LOC_92/Y 0.04fF
C46213 OR2X1_LOC_516/A AND2X1_LOC_212/Y 0.12fF
C46214 OR2X1_LOC_204/Y AND2X1_LOC_44/Y 0.03fF
C46215 OR2X1_LOC_118/a_8_216# OR2X1_LOC_85/A 0.14fF
C46216 OR2X1_LOC_474/Y OR2X1_LOC_244/Y 0.05fF
C46217 AND2X1_LOC_51/Y OR2X1_LOC_508/Y 0.09fF
C46218 OR2X1_LOC_708/B OR2X1_LOC_779/A 0.01fF
C46219 OR2X1_LOC_620/Y OR2X1_LOC_302/A 0.29fF
C46220 OR2X1_LOC_482/Y AND2X1_LOC_573/A 0.03fF
C46221 OR2X1_LOC_158/A OR2X1_LOC_32/B 0.58fF
C46222 OR2X1_LOC_132/Y OR2X1_LOC_517/A 0.12fF
C46223 AND2X1_LOC_721/Y OR2X1_LOC_669/Y 0.01fF
C46224 OR2X1_LOC_538/A OR2X1_LOC_703/A 1.36fF
C46225 OR2X1_LOC_421/A AND2X1_LOC_644/Y 0.00fF
C46226 OR2X1_LOC_753/A OR2X1_LOC_15/a_8_216# 0.03fF
C46227 OR2X1_LOC_599/A AND2X1_LOC_828/a_8_24# 0.03fF
C46228 OR2X1_LOC_656/B AND2X1_LOC_18/Y 0.01fF
C46229 INPUT_3 INPUT_2 0.52fF
C46230 OR2X1_LOC_78/A OR2X1_LOC_574/a_8_216# 0.19fF
C46231 OR2X1_LOC_600/A AND2X1_LOC_468/B 0.15fF
C46232 OR2X1_LOC_121/Y OR2X1_LOC_116/a_8_216# 0.02fF
C46233 OR2X1_LOC_751/Y OR2X1_LOC_820/A 0.03fF
C46234 AND2X1_LOC_123/Y AND2X1_LOC_243/Y 0.04fF
C46235 AND2X1_LOC_42/B OR2X1_LOC_267/Y 1.10fF
C46236 OR2X1_LOC_604/A AND2X1_LOC_453/Y 0.01fF
C46237 OR2X1_LOC_320/Y OR2X1_LOC_321/a_8_216# 0.46fF
C46238 AND2X1_LOC_658/A OR2X1_LOC_531/a_8_216# 0.03fF
C46239 OR2X1_LOC_185/Y OR2X1_LOC_361/a_8_216# 0.20fF
C46240 OR2X1_LOC_12/Y AND2X1_LOC_454/A 0.01fF
C46241 AND2X1_LOC_804/Y AND2X1_LOC_469/B 0.00fF
C46242 OR2X1_LOC_814/A OR2X1_LOC_776/A 0.02fF
C46243 OR2X1_LOC_177/Y OR2X1_LOC_26/Y 0.06fF
C46244 OR2X1_LOC_643/A OR2X1_LOC_549/A 0.07fF
C46245 OR2X1_LOC_161/A OR2X1_LOC_66/A 1.21fF
C46246 AND2X1_LOC_857/Y OR2X1_LOC_298/a_8_216# 0.01fF
C46247 OR2X1_LOC_203/Y OR2X1_LOC_719/B 0.17fF
C46248 OR2X1_LOC_45/B OR2X1_LOC_74/A 13.05fF
C46249 D_GATE_479 OR2X1_LOC_453/Y 0.01fF
C46250 AND2X1_LOC_786/a_8_24# OR2X1_LOC_70/Y 0.17fF
C46251 OR2X1_LOC_124/Y OR2X1_LOC_549/A 0.16fF
C46252 AND2X1_LOC_195/a_36_24# OR2X1_LOC_43/A 0.00fF
C46253 AND2X1_LOC_523/Y AND2X1_LOC_465/A 0.08fF
C46254 OR2X1_LOC_59/Y OR2X1_LOC_278/Y 0.04fF
C46255 OR2X1_LOC_53/Y AND2X1_LOC_729/B 0.02fF
C46256 OR2X1_LOC_468/A AND2X1_LOC_43/B 0.03fF
C46257 AND2X1_LOC_738/B AND2X1_LOC_593/Y 2.08fF
C46258 AND2X1_LOC_758/a_36_24# OR2X1_LOC_616/Y 0.00fF
C46259 OR2X1_LOC_453/Y OR2X1_LOC_161/B 0.01fF
C46260 OR2X1_LOC_36/Y AND2X1_LOC_194/Y 0.01fF
C46261 AND2X1_LOC_12/Y AND2X1_LOC_70/Y 0.35fF
C46262 VDD OR2X1_LOC_470/A -0.00fF
C46263 OR2X1_LOC_296/Y OR2X1_LOC_161/B 0.01fF
C46264 OR2X1_LOC_318/Y OR2X1_LOC_435/B 0.16fF
C46265 OR2X1_LOC_154/A VDD 2.40fF
C46266 AND2X1_LOC_42/B OR2X1_LOC_633/A 0.15fF
C46267 OR2X1_LOC_22/Y OR2X1_LOC_171/Y 0.39fF
C46268 OR2X1_LOC_177/Y OR2X1_LOC_89/A 0.04fF
C46269 OR2X1_LOC_357/A OR2X1_LOC_365/B 0.02fF
C46270 AND2X1_LOC_733/Y AND2X1_LOC_804/Y 0.01fF
C46271 OR2X1_LOC_799/A OR2X1_LOC_78/B 0.03fF
C46272 AND2X1_LOC_474/A AND2X1_LOC_850/Y 0.01fF
C46273 OR2X1_LOC_793/A AND2X1_LOC_18/Y 0.01fF
C46274 OR2X1_LOC_458/a_8_216# OR2X1_LOC_737/A 0.05fF
C46275 OR2X1_LOC_648/A AND2X1_LOC_601/a_8_24# 0.04fF
C46276 OR2X1_LOC_44/Y AND2X1_LOC_860/A 4.46fF
C46277 AND2X1_LOC_456/B AND2X1_LOC_843/Y 0.01fF
C46278 OR2X1_LOC_11/Y OR2X1_LOC_585/Y 0.01fF
C46279 AND2X1_LOC_244/a_8_24# AND2X1_LOC_806/A 0.01fF
C46280 AND2X1_LOC_860/A AND2X1_LOC_288/a_8_24# 0.01fF
C46281 AND2X1_LOC_25/Y OR2X1_LOC_66/A 0.00fF
C46282 OR2X1_LOC_367/B OR2X1_LOC_365/B 0.05fF
C46283 AND2X1_LOC_311/a_8_24# OR2X1_LOC_161/A 0.02fF
C46284 OR2X1_LOC_329/B AND2X1_LOC_113/Y 0.00fF
C46285 OR2X1_LOC_604/A OR2X1_LOC_26/Y 0.09fF
C46286 OR2X1_LOC_619/Y OR2X1_LOC_234/Y 0.01fF
C46287 AND2X1_LOC_713/Y OR2X1_LOC_52/B 0.01fF
C46288 AND2X1_LOC_565/a_36_24# AND2X1_LOC_580/A 0.00fF
C46289 OR2X1_LOC_6/B OR2X1_LOC_84/B 0.08fF
C46290 OR2X1_LOC_160/B OR2X1_LOC_269/B 0.12fF
C46291 VDD OR2X1_LOC_267/A 0.08fF
C46292 AND2X1_LOC_40/Y OR2X1_LOC_856/B 0.02fF
C46293 OR2X1_LOC_52/B AND2X1_LOC_448/a_36_24# 0.01fF
C46294 OR2X1_LOC_49/A AND2X1_LOC_260/a_36_24# 0.00fF
C46295 OR2X1_LOC_85/A OR2X1_LOC_56/A 0.34fF
C46296 AND2X1_LOC_59/Y OR2X1_LOC_235/B 0.03fF
C46297 OR2X1_LOC_705/Y OR2X1_LOC_725/A 0.02fF
C46298 AND2X1_LOC_50/Y AND2X1_LOC_53/a_36_24# 0.01fF
C46299 OR2X1_LOC_64/Y AND2X1_LOC_771/a_8_24# 0.01fF
C46300 OR2X1_LOC_843/a_8_216# OR2X1_LOC_362/A 0.01fF
C46301 OR2X1_LOC_421/A OR2X1_LOC_7/A 0.05fF
C46302 OR2X1_LOC_40/Y AND2X1_LOC_717/B 0.02fF
C46303 AND2X1_LOC_12/Y OR2X1_LOC_703/A 0.06fF
C46304 OR2X1_LOC_405/A OR2X1_LOC_802/a_8_216# 0.06fF
C46305 OR2X1_LOC_604/A OR2X1_LOC_89/A 0.23fF
C46306 AND2X1_LOC_544/a_8_24# AND2X1_LOC_550/A 0.02fF
C46307 OR2X1_LOC_792/Y OR2X1_LOC_805/a_8_216# 0.02fF
C46308 OR2X1_LOC_541/A AND2X1_LOC_272/a_36_24# 0.00fF
C46309 OR2X1_LOC_638/a_8_216# OR2X1_LOC_375/A 0.01fF
C46310 AND2X1_LOC_724/Y AND2X1_LOC_602/a_36_24# 0.00fF
C46311 OR2X1_LOC_261/A OR2X1_LOC_382/A 0.27fF
C46312 OR2X1_LOC_744/A OR2X1_LOC_588/Y 0.68fF
C46313 AND2X1_LOC_568/B AND2X1_LOC_566/Y 0.04fF
C46314 OR2X1_LOC_748/A OR2X1_LOC_91/A 0.02fF
C46315 OR2X1_LOC_792/Y OR2X1_LOC_362/B 0.05fF
C46316 VDD AND2X1_LOC_554/B 0.50fF
C46317 OR2X1_LOC_113/Y OR2X1_LOC_643/A 0.01fF
C46318 OR2X1_LOC_121/B OR2X1_LOC_356/A 0.03fF
C46319 OR2X1_LOC_97/A OR2X1_LOC_602/B 0.01fF
C46320 VDD OR2X1_LOC_680/Y 0.30fF
C46321 OR2X1_LOC_92/Y AND2X1_LOC_848/Y 0.03fF
C46322 OR2X1_LOC_856/B OR2X1_LOC_537/A 0.05fF
C46323 OR2X1_LOC_308/a_8_216# OR2X1_LOC_375/A 0.01fF
C46324 OR2X1_LOC_574/A AND2X1_LOC_92/Y 0.10fF
C46325 AND2X1_LOC_539/a_8_24# OR2X1_LOC_12/Y 0.01fF
C46326 OR2X1_LOC_634/A AND2X1_LOC_412/a_8_24# 0.01fF
C46327 OR2X1_LOC_485/A AND2X1_LOC_468/a_8_24# 0.02fF
C46328 OR2X1_LOC_61/Y OR2X1_LOC_805/A 0.07fF
C46329 OR2X1_LOC_298/Y AND2X1_LOC_654/Y 0.87fF
C46330 VDD OR2X1_LOC_778/A 0.18fF
C46331 OR2X1_LOC_216/A OR2X1_LOC_87/A 0.07fF
C46332 AND2X1_LOC_41/A OR2X1_LOC_710/a_8_216# 0.01fF
C46333 AND2X1_LOC_70/Y AND2X1_LOC_496/a_8_24# 0.01fF
C46334 AND2X1_LOC_272/a_8_24# OR2X1_LOC_737/A 0.00fF
C46335 OR2X1_LOC_207/B AND2X1_LOC_53/Y 0.08fF
C46336 OR2X1_LOC_625/a_8_216# OR2X1_LOC_67/A 0.07fF
C46337 OR2X1_LOC_114/B OR2X1_LOC_404/Y 0.00fF
C46338 AND2X1_LOC_70/Y OR2X1_LOC_804/B 0.70fF
C46339 D_INPUT_0 OR2X1_LOC_595/A 0.14fF
C46340 AND2X1_LOC_161/a_36_24# OR2X1_LOC_619/Y 0.00fF
C46341 VDD OR2X1_LOC_696/Y 0.15fF
C46342 AND2X1_LOC_181/a_8_24# OR2X1_LOC_485/A 0.01fF
C46343 OR2X1_LOC_160/B AND2X1_LOC_75/a_8_24# 0.04fF
C46344 AND2X1_LOC_76/Y AND2X1_LOC_139/B 0.03fF
C46345 OR2X1_LOC_95/Y AND2X1_LOC_407/a_8_24# 0.01fF
C46346 VDD AND2X1_LOC_326/A 0.21fF
C46347 AND2X1_LOC_51/Y OR2X1_LOC_66/A 0.23fF
C46348 VDD OR2X1_LOC_345/A -0.00fF
C46349 AND2X1_LOC_141/B AND2X1_LOC_141/a_8_24# 0.06fF
C46350 OR2X1_LOC_441/Y OR2X1_LOC_52/B 0.11fF
C46351 OR2X1_LOC_354/A OR2X1_LOC_778/Y 0.10fF
C46352 AND2X1_LOC_456/B OR2X1_LOC_7/A 0.31fF
C46353 AND2X1_LOC_319/A OR2X1_LOC_48/B 0.07fF
C46354 OR2X1_LOC_427/A AND2X1_LOC_453/a_36_24# 0.00fF
C46355 AND2X1_LOC_17/Y D_INPUT_5 0.18fF
C46356 AND2X1_LOC_776/a_8_24# OR2X1_LOC_64/Y 0.03fF
C46357 OR2X1_LOC_32/Y OR2X1_LOC_58/a_36_216# 0.02fF
C46358 AND2X1_LOC_12/Y OR2X1_LOC_791/B 0.01fF
C46359 AND2X1_LOC_454/Y AND2X1_LOC_452/Y 0.07fF
C46360 AND2X1_LOC_45/a_8_24# AND2X1_LOC_18/Y 0.01fF
C46361 VDD AND2X1_LOC_351/Y 0.04fF
C46362 OR2X1_LOC_419/Y AND2X1_LOC_590/a_8_24# 0.11fF
C46363 OR2X1_LOC_699/a_8_216# OR2X1_LOC_427/A 0.05fF
C46364 AND2X1_LOC_56/B AND2X1_LOC_16/a_8_24# -0.00fF
C46365 OR2X1_LOC_432/a_8_216# OR2X1_LOC_44/Y 0.01fF
C46366 AND2X1_LOC_608/a_8_24# OR2X1_LOC_71/A 0.03fF
C46367 OR2X1_LOC_849/a_8_216# OR2X1_LOC_66/A 0.01fF
C46368 OR2X1_LOC_680/Y OR2X1_LOC_677/Y 0.03fF
C46369 OR2X1_LOC_91/Y OR2X1_LOC_39/A 0.17fF
C46370 AND2X1_LOC_400/a_8_24# OR2X1_LOC_44/Y 0.17fF
C46371 D_INPUT_7 D_INPUT_4 0.08fF
C46372 AND2X1_LOC_857/Y OR2X1_LOC_229/Y 0.01fF
C46373 AND2X1_LOC_215/Y AND2X1_LOC_633/Y 0.03fF
C46374 OR2X1_LOC_461/a_8_216# OR2X1_LOC_472/B 0.01fF
C46375 OR2X1_LOC_377/A AND2X1_LOC_56/B 0.18fF
C46376 AND2X1_LOC_17/Y AND2X1_LOC_22/a_8_24# 0.01fF
C46377 OR2X1_LOC_813/A AND2X1_LOC_243/Y 0.03fF
C46378 OR2X1_LOC_69/A OR2X1_LOC_69/a_8_216# 0.00fF
C46379 OR2X1_LOC_216/A OR2X1_LOC_216/a_8_216# 0.08fF
C46380 OR2X1_LOC_476/B AND2X1_LOC_19/Y 0.01fF
C46381 OR2X1_LOC_83/A OR2X1_LOC_394/Y 0.01fF
C46382 AND2X1_LOC_348/A OR2X1_LOC_485/A 0.01fF
C46383 OR2X1_LOC_270/a_8_216# OR2X1_LOC_375/A 0.02fF
C46384 OR2X1_LOC_19/B OR2X1_LOC_59/Y 0.16fF
C46385 OR2X1_LOC_703/B OR2X1_LOC_169/a_8_216# 0.05fF
C46386 AND2X1_LOC_219/a_8_24# INPUT_1 0.01fF
C46387 OR2X1_LOC_743/A OR2X1_LOC_761/Y 0.01fF
C46388 AND2X1_LOC_56/B AND2X1_LOC_824/B 0.26fF
C46389 AND2X1_LOC_334/Y INPUT_1 0.15fF
C46390 AND2X1_LOC_87/a_8_24# OR2X1_LOC_85/A 0.01fF
C46391 OR2X1_LOC_532/B OR2X1_LOC_776/Y 0.46fF
C46392 OR2X1_LOC_377/A AND2X1_LOC_8/Y 0.10fF
C46393 OR2X1_LOC_189/a_8_216# AND2X1_LOC_711/Y 0.05fF
C46394 OR2X1_LOC_553/B OR2X1_LOC_563/B 0.09fF
C46395 AND2X1_LOC_95/Y AND2X1_LOC_252/a_36_24# 0.01fF
C46396 VDD OR2X1_LOC_167/Y 0.37fF
C46397 OR2X1_LOC_703/B OR2X1_LOC_468/Y 0.02fF
C46398 AND2X1_LOC_348/A AND2X1_LOC_348/a_8_24# 0.10fF
C46399 AND2X1_LOC_43/B OR2X1_LOC_449/B 0.04fF
C46400 AND2X1_LOC_12/Y AND2X1_LOC_17/Y 0.01fF
C46401 AND2X1_LOC_95/Y OR2X1_LOC_445/a_8_216# 0.03fF
C46402 OR2X1_LOC_235/a_8_216# OR2X1_LOC_6/A 0.14fF
C46403 AND2X1_LOC_851/a_36_24# AND2X1_LOC_465/Y 0.01fF
C46404 OR2X1_LOC_426/B AND2X1_LOC_845/Y 0.08fF
C46405 AND2X1_LOC_41/A OR2X1_LOC_750/A 0.01fF
C46406 AND2X1_LOC_8/Y AND2X1_LOC_824/B 0.01fF
C46407 OR2X1_LOC_553/A OR2X1_LOC_269/B 0.27fF
C46408 OR2X1_LOC_472/B OR2X1_LOC_634/A 0.33fF
C46409 AND2X1_LOC_56/B OR2X1_LOC_203/Y 0.04fF
C46410 AND2X1_LOC_139/B OR2X1_LOC_52/B 0.07fF
C46411 AND2X1_LOC_286/Y AND2X1_LOC_806/A 0.00fF
C46412 AND2X1_LOC_287/Y AND2X1_LOC_288/a_8_24# 0.01fF
C46413 OR2X1_LOC_604/A OR2X1_LOC_426/a_8_216# 0.01fF
C46414 OR2X1_LOC_158/A AND2X1_LOC_116/a_8_24# 0.02fF
C46415 OR2X1_LOC_503/a_8_216# AND2X1_LOC_657/A 0.02fF
C46416 OR2X1_LOC_80/Y OR2X1_LOC_26/Y 0.07fF
C46417 OR2X1_LOC_810/A OR2X1_LOC_130/A 0.07fF
C46418 AND2X1_LOC_367/a_8_24# OR2X1_LOC_753/A 0.03fF
C46419 OR2X1_LOC_70/Y OR2X1_LOC_278/Y 0.00fF
C46420 OR2X1_LOC_51/Y AND2X1_LOC_859/B 0.02fF
C46421 OR2X1_LOC_817/a_36_216# AND2X1_LOC_847/Y 0.01fF
C46422 OR2X1_LOC_91/Y AND2X1_LOC_211/B 0.58fF
C46423 OR2X1_LOC_816/A OR2X1_LOC_754/Y 0.05fF
C46424 OR2X1_LOC_502/A AND2X1_LOC_48/A 0.03fF
C46425 OR2X1_LOC_593/A OR2X1_LOC_593/a_8_216# 0.39fF
C46426 OR2X1_LOC_696/A OR2X1_LOC_589/a_8_216# 0.07fF
C46427 OR2X1_LOC_847/A OR2X1_LOC_5/a_8_216# 0.47fF
C46428 AND2X1_LOC_390/B AND2X1_LOC_655/A 0.10fF
C46429 AND2X1_LOC_589/a_8_24# OR2X1_LOC_130/A 0.03fF
C46430 OR2X1_LOC_40/Y AND2X1_LOC_675/a_36_24# 0.00fF
C46431 AND2X1_LOC_40/Y OR2X1_LOC_383/Y 0.10fF
C46432 AND2X1_LOC_12/Y OR2X1_LOC_206/a_8_216# 0.01fF
C46433 OR2X1_LOC_665/Y AND2X1_LOC_859/Y 0.04fF
C46434 OR2X1_LOC_756/B OR2X1_LOC_532/B 0.64fF
C46435 AND2X1_LOC_658/B AND2X1_LOC_803/a_8_24# 0.02fF
C46436 AND2X1_LOC_191/Y AND2X1_LOC_565/Y 0.07fF
C46437 OR2X1_LOC_189/Y AND2X1_LOC_569/a_8_24# 0.23fF
C46438 OR2X1_LOC_87/A AND2X1_LOC_19/a_36_24# 0.00fF
C46439 OR2X1_LOC_604/A AND2X1_LOC_451/a_8_24# 0.01fF
C46440 VDD OR2X1_LOC_84/a_8_216# 0.00fF
C46441 OR2X1_LOC_75/Y OR2X1_LOC_59/Y 0.07fF
C46442 AND2X1_LOC_271/a_8_24# AND2X1_LOC_18/Y 0.01fF
C46443 AND2X1_LOC_699/a_8_24# OR2X1_LOC_596/A 0.00fF
C46444 OR2X1_LOC_644/B AND2X1_LOC_3/Y 0.00fF
C46445 VDD AND2X1_LOC_6/a_8_24# 0.00fF
C46446 OR2X1_LOC_527/Y OR2X1_LOC_39/A 0.35fF
C46447 AND2X1_LOC_12/Y OR2X1_LOC_404/Y 0.75fF
C46448 OR2X1_LOC_485/A AND2X1_LOC_859/Y 0.07fF
C46449 OR2X1_LOC_604/A OR2X1_LOC_419/a_8_216# 0.04fF
C46450 OR2X1_LOC_808/a_8_216# OR2X1_LOC_814/A 0.02fF
C46451 OR2X1_LOC_235/a_36_216# OR2X1_LOC_74/A 0.00fF
C46452 OR2X1_LOC_291/A OR2X1_LOC_85/A 0.05fF
C46453 AND2X1_LOC_514/Y AND2X1_LOC_662/B 0.00fF
C46454 AND2X1_LOC_711/Y AND2X1_LOC_565/Y 0.03fF
C46455 OR2X1_LOC_278/A OR2X1_LOC_619/Y 3.79fF
C46456 OR2X1_LOC_280/Y AND2X1_LOC_806/A 0.02fF
C46457 OR2X1_LOC_36/Y OR2X1_LOC_17/Y 0.00fF
C46458 OR2X1_LOC_364/A OR2X1_LOC_602/a_8_216# -0.04fF
C46459 AND2X1_LOC_7/B AND2X1_LOC_406/a_8_24# 0.02fF
C46460 AND2X1_LOC_523/Y OR2X1_LOC_237/Y 0.03fF
C46461 OR2X1_LOC_70/Y AND2X1_LOC_565/Y 0.04fF
C46462 OR2X1_LOC_175/B D_INPUT_0 0.01fF
C46463 OR2X1_LOC_794/a_8_216# OR2X1_LOC_269/B 0.02fF
C46464 OR2X1_LOC_291/Y OR2X1_LOC_39/A 0.05fF
C46465 OR2X1_LOC_121/B AND2X1_LOC_43/B 0.07fF
C46466 AND2X1_LOC_75/a_8_24# OR2X1_LOC_553/A 0.04fF
C46467 OR2X1_LOC_629/B OR2X1_LOC_598/A 0.02fF
C46468 OR2X1_LOC_158/A AND2X1_LOC_222/Y 0.03fF
C46469 INPUT_1 AND2X1_LOC_649/B 0.33fF
C46470 AND2X1_LOC_717/B OR2X1_LOC_7/A 5.49fF
C46471 OR2X1_LOC_679/A AND2X1_LOC_147/a_36_24# 0.00fF
C46472 OR2X1_LOC_857/a_8_216# OR2X1_LOC_130/A 0.14fF
C46473 OR2X1_LOC_149/B OR2X1_LOC_550/B 0.03fF
C46474 AND2X1_LOC_1/Y OR2X1_LOC_87/A 0.00fF
C46475 OR2X1_LOC_46/A AND2X1_LOC_233/a_8_24# 0.01fF
C46476 VDD OR2X1_LOC_99/A 0.05fF
C46477 AND2X1_LOC_556/a_8_24# OR2X1_LOC_615/Y 0.03fF
C46478 OR2X1_LOC_756/B OR2X1_LOC_343/B 0.15fF
C46479 VDD OR2X1_LOC_739/Y -0.00fF
C46480 OR2X1_LOC_154/A OR2X1_LOC_476/a_36_216# 0.01fF
C46481 OR2X1_LOC_687/Y AND2X1_LOC_430/a_8_24# 0.23fF
C46482 OR2X1_LOC_158/A OR2X1_LOC_68/B 0.03fF
C46483 AND2X1_LOC_362/B AND2X1_LOC_657/A 0.07fF
C46484 OR2X1_LOC_510/Y OR2X1_LOC_62/B 0.01fF
C46485 OR2X1_LOC_687/B OR2X1_LOC_687/a_8_216# 0.39fF
C46486 OR2X1_LOC_70/Y AND2X1_LOC_337/B 0.01fF
C46487 AND2X1_LOC_342/Y OR2X1_LOC_255/a_8_216# 0.06fF
C46488 OR2X1_LOC_139/A OR2X1_LOC_217/A 0.02fF
C46489 OR2X1_LOC_415/a_8_216# OR2X1_LOC_753/A 0.35fF
C46490 OR2X1_LOC_471/Y OR2X1_LOC_87/A 0.05fF
C46491 OR2X1_LOC_204/Y OR2X1_LOC_720/B 0.03fF
C46492 OR2X1_LOC_22/Y AND2X1_LOC_806/A 0.03fF
C46493 OR2X1_LOC_158/A OR2X1_LOC_423/Y 0.01fF
C46494 VDD OR2X1_LOC_560/A 0.41fF
C46495 OR2X1_LOC_344/A OR2X1_LOC_367/a_8_216# 0.01fF
C46496 OR2X1_LOC_246/A OR2X1_LOC_753/A 0.14fF
C46497 VDD OR2X1_LOC_198/A 0.48fF
C46498 AND2X1_LOC_714/B OR2X1_LOC_589/Y 0.14fF
C46499 OR2X1_LOC_526/Y AND2X1_LOC_796/A 0.28fF
C46500 AND2X1_LOC_53/Y OR2X1_LOC_790/a_8_216# 0.04fF
C46501 AND2X1_LOC_159/a_8_24# OR2X1_LOC_62/B 0.11fF
C46502 OR2X1_LOC_436/Y OR2X1_LOC_539/Y 0.05fF
C46503 OR2X1_LOC_810/A OR2X1_LOC_62/B 0.05fF
C46504 AND2X1_LOC_727/a_8_24# OR2X1_LOC_142/Y 0.01fF
C46505 AND2X1_LOC_514/Y AND2X1_LOC_337/B 0.02fF
C46506 AND2X1_LOC_59/Y OR2X1_LOC_276/B 0.09fF
C46507 OR2X1_LOC_864/A AND2X1_LOC_15/a_8_24# 0.03fF
C46508 OR2X1_LOC_364/A OR2X1_LOC_439/a_8_216# 0.02fF
C46509 OR2X1_LOC_76/Y OR2X1_LOC_532/B 0.03fF
C46510 OR2X1_LOC_70/A OR2X1_LOC_763/a_8_216# 0.00fF
C46511 OR2X1_LOC_70/Y OR2X1_LOC_19/B 0.01fF
C46512 OR2X1_LOC_18/Y AND2X1_LOC_721/A 0.02fF
C46513 OR2X1_LOC_22/Y AND2X1_LOC_276/Y 0.01fF
C46514 OR2X1_LOC_685/B AND2X1_LOC_681/a_8_24# 0.00fF
C46515 OR2X1_LOC_43/A OR2X1_LOC_55/a_8_216# 0.03fF
C46516 OR2X1_LOC_409/B OR2X1_LOC_753/A 0.00fF
C46517 AND2X1_LOC_53/Y AND2X1_LOC_3/Y 0.07fF
C46518 AND2X1_LOC_191/Y AND2X1_LOC_630/a_36_24# 0.01fF
C46519 OR2X1_LOC_678/Y OR2X1_LOC_513/Y 0.01fF
C46520 OR2X1_LOC_276/B AND2X1_LOC_495/a_8_24# 0.02fF
C46521 OR2X1_LOC_78/A OR2X1_LOC_317/B 0.03fF
C46522 OR2X1_LOC_78/B OR2X1_LOC_446/B 0.01fF
C46523 AND2X1_LOC_554/B OR2X1_LOC_256/A 0.27fF
C46524 AND2X1_LOC_518/a_8_24# AND2X1_LOC_48/A 0.01fF
C46525 AND2X1_LOC_539/Y OR2X1_LOC_428/A 0.03fF
C46526 OR2X1_LOC_87/A OR2X1_LOC_205/Y 0.02fF
C46527 OR2X1_LOC_47/Y OR2X1_LOC_612/B 0.03fF
C46528 OR2X1_LOC_136/a_8_216# AND2X1_LOC_358/Y 0.04fF
C46529 AND2X1_LOC_811/Y OR2X1_LOC_74/A 0.11fF
C46530 OR2X1_LOC_359/A OR2X1_LOC_349/B 0.04fF
C46531 AND2X1_LOC_139/B AND2X1_LOC_216/A 0.14fF
C46532 OR2X1_LOC_218/Y OR2X1_LOC_216/a_36_216# 0.03fF
C46533 OR2X1_LOC_3/Y AND2X1_LOC_476/A 0.07fF
C46534 AND2X1_LOC_91/B OR2X1_LOC_843/B 0.08fF
C46535 OR2X1_LOC_850/a_8_216# OR2X1_LOC_580/A 0.03fF
C46536 OR2X1_LOC_847/A OR2X1_LOC_68/B 0.03fF
C46537 OR2X1_LOC_726/A OR2X1_LOC_731/A 0.09fF
C46538 OR2X1_LOC_70/Y OR2X1_LOC_75/Y 0.06fF
C46539 AND2X1_LOC_64/Y OR2X1_LOC_729/a_8_216# 0.05fF
C46540 AND2X1_LOC_394/a_8_24# OR2X1_LOC_398/Y 0.01fF
C46541 AND2X1_LOC_91/B OR2X1_LOC_549/A 0.10fF
C46542 OR2X1_LOC_212/A OR2X1_LOC_353/a_8_216# 0.01fF
C46543 OR2X1_LOC_604/A AND2X1_LOC_590/a_8_24# 0.01fF
C46544 OR2X1_LOC_189/Y AND2X1_LOC_781/Y 0.15fF
C46545 AND2X1_LOC_778/a_36_24# AND2X1_LOC_778/Y 0.00fF
C46546 OR2X1_LOC_25/Y D_INPUT_6 0.01fF
C46547 AND2X1_LOC_278/a_36_24# OR2X1_LOC_68/B 0.00fF
C46548 OR2X1_LOC_45/B AND2X1_LOC_810/A 0.01fF
C46549 OR2X1_LOC_92/Y OR2X1_LOC_536/a_8_216# 0.05fF
C46550 AND2X1_LOC_483/a_36_24# OR2X1_LOC_615/Y 0.00fF
C46551 OR2X1_LOC_789/a_8_216# OR2X1_LOC_801/B 0.04fF
C46552 OR2X1_LOC_638/B AND2X1_LOC_408/a_8_24# 0.20fF
C46553 OR2X1_LOC_52/B OR2X1_LOC_598/A 0.34fF
C46554 OR2X1_LOC_16/A AND2X1_LOC_786/Y 0.02fF
C46555 OR2X1_LOC_708/Y OR2X1_LOC_712/B 0.06fF
C46556 OR2X1_LOC_84/B OR2X1_LOC_598/A 0.00fF
C46557 OR2X1_LOC_84/A AND2X1_LOC_51/Y 0.00fF
C46558 OR2X1_LOC_161/B OR2X1_LOC_580/B 0.03fF
C46559 OR2X1_LOC_696/A OR2X1_LOC_369/Y -0.01fF
C46560 OR2X1_LOC_44/Y AND2X1_LOC_562/Y 0.04fF
C46561 AND2X1_LOC_390/B OR2X1_LOC_599/Y 0.08fF
C46562 VDD OR2X1_LOC_503/a_8_216# 0.00fF
C46563 OR2X1_LOC_96/a_8_216# OR2X1_LOC_46/A 0.01fF
C46564 D_INPUT_3 AND2X1_LOC_672/B 0.54fF
C46565 OR2X1_LOC_119/a_36_216# D_INPUT_1 0.03fF
C46566 OR2X1_LOC_435/A AND2X1_LOC_433/a_36_24# 0.00fF
C46567 AND2X1_LOC_555/Y OR2X1_LOC_56/A 0.17fF
C46568 OR2X1_LOC_375/A OR2X1_LOC_446/B 0.03fF
C46569 AND2X1_LOC_565/B OR2X1_LOC_406/Y 0.02fF
C46570 AND2X1_LOC_191/B AND2X1_LOC_465/A 0.09fF
C46571 OR2X1_LOC_45/B AND2X1_LOC_340/a_8_24# 0.01fF
C46572 OR2X1_LOC_177/Y AND2X1_LOC_552/A 0.01fF
C46573 OR2X1_LOC_131/A OR2X1_LOC_595/A 0.26fF
C46574 OR2X1_LOC_89/Y OR2X1_LOC_59/Y 0.12fF
C46575 OR2X1_LOC_651/A AND2X1_LOC_47/Y 0.03fF
C46576 OR2X1_LOC_364/B OR2X1_LOC_182/B 0.01fF
C46577 AND2X1_LOC_721/Y AND2X1_LOC_489/a_36_24# 0.01fF
C46578 AND2X1_LOC_711/A OR2X1_LOC_428/A 0.02fF
C46579 AND2X1_LOC_64/Y OR2X1_LOC_114/a_8_216# 0.01fF
C46580 AND2X1_LOC_326/B OR2X1_LOC_428/A 0.03fF
C46581 AND2X1_LOC_621/Y OR2X1_LOC_142/Y 0.03fF
C46582 OR2X1_LOC_167/a_8_216# OR2X1_LOC_604/A 0.12fF
C46583 AND2X1_LOC_43/B OR2X1_LOC_195/a_8_216# 0.04fF
C46584 AND2X1_LOC_476/Y AND2X1_LOC_479/a_8_24# 0.03fF
C46585 OR2X1_LOC_421/A OR2X1_LOC_693/a_36_216# 0.00fF
C46586 AND2X1_LOC_785/A OR2X1_LOC_427/A 0.02fF
C46587 OR2X1_LOC_497/Y OR2X1_LOC_437/A 0.19fF
C46588 OR2X1_LOC_270/a_36_216# D_GATE_366 0.00fF
C46589 AND2X1_LOC_721/Y AND2X1_LOC_362/a_8_24# 0.05fF
C46590 OR2X1_LOC_78/A AND2X1_LOC_44/Y 1.53fF
C46591 OR2X1_LOC_636/a_8_216# AND2X1_LOC_31/Y 0.01fF
C46592 OR2X1_LOC_604/A AND2X1_LOC_605/a_8_24# 0.01fF
C46593 AND2X1_LOC_552/A OR2X1_LOC_604/A 0.13fF
C46594 OR2X1_LOC_338/a_8_216# OR2X1_LOC_160/B 0.05fF
C46595 AND2X1_LOC_91/B OR2X1_LOC_354/A 0.07fF
C46596 AND2X1_LOC_64/Y OR2X1_LOC_854/a_8_216# 0.01fF
C46597 AND2X1_LOC_564/B AND2X1_LOC_734/Y 0.00fF
C46598 OR2X1_LOC_756/B OR2X1_LOC_392/a_36_216# 0.00fF
C46599 AND2X1_LOC_681/a_36_24# OR2X1_LOC_161/B 0.00fF
C46600 VDD AND2X1_LOC_476/Y 0.47fF
C46601 AND2X1_LOC_362/B VDD 0.25fF
C46602 OR2X1_LOC_114/B OR2X1_LOC_362/A 0.03fF
C46603 OR2X1_LOC_696/A OR2X1_LOC_53/a_8_216# 0.05fF
C46604 OR2X1_LOC_648/A OR2X1_LOC_390/A 0.01fF
C46605 OR2X1_LOC_336/a_8_216# OR2X1_LOC_538/A 0.07fF
C46606 OR2X1_LOC_160/A AND2X1_LOC_235/a_8_24# 0.01fF
C46607 OR2X1_LOC_62/A D_INPUT_1 0.17fF
C46608 OR2X1_LOC_19/B AND2X1_LOC_31/Y 0.03fF
C46609 VDD AND2X1_LOC_299/a_8_24# 0.00fF
C46610 OR2X1_LOC_106/Y OR2X1_LOC_427/A 0.07fF
C46611 OR2X1_LOC_744/A AND2X1_LOC_828/a_36_24# 0.00fF
C46612 OR2X1_LOC_815/a_8_216# OR2X1_LOC_600/A 0.01fF
C46613 AND2X1_LOC_512/Y AND2X1_LOC_809/a_8_24# 0.01fF
C46614 AND2X1_LOC_476/A AND2X1_LOC_462/B 0.13fF
C46615 AND2X1_LOC_716/Y OR2X1_LOC_310/a_8_216# 0.03fF
C46616 OR2X1_LOC_241/Y OR2X1_LOC_493/Y 0.03fF
C46617 OR2X1_LOC_629/A OR2X1_LOC_777/B 0.99fF
C46618 AND2X1_LOC_12/Y OR2X1_LOC_718/a_8_216# 0.01fF
C46619 OR2X1_LOC_448/B AND2X1_LOC_44/Y 0.10fF
C46620 AND2X1_LOC_719/Y OR2X1_LOC_744/A 0.17fF
C46621 OR2X1_LOC_39/A AND2X1_LOC_780/a_8_24# 0.01fF
C46622 OR2X1_LOC_207/B OR2X1_LOC_502/A 0.02fF
C46623 OR2X1_LOC_121/Y OR2X1_LOC_474/Y 0.07fF
C46624 OR2X1_LOC_158/A AND2X1_LOC_367/A 0.01fF
C46625 OR2X1_LOC_147/a_36_216# OR2X1_LOC_375/A 0.00fF
C46626 OR2X1_LOC_234/a_36_216# D_INPUT_1 0.00fF
C46627 OR2X1_LOC_71/Y OR2X1_LOC_88/Y 0.07fF
C46628 OR2X1_LOC_549/a_8_216# OR2X1_LOC_456/Y 0.40fF
C46629 AND2X1_LOC_5/a_8_24# OR2X1_LOC_80/A 0.01fF
C46630 OR2X1_LOC_139/A OR2X1_LOC_185/A 0.03fF
C46631 OR2X1_LOC_64/a_36_216# OR2X1_LOC_70/A 0.00fF
C46632 AND2X1_LOC_738/B OR2X1_LOC_51/Y 0.07fF
C46633 OR2X1_LOC_326/B OR2X1_LOC_186/Y 0.07fF
C46634 OR2X1_LOC_51/Y OR2X1_LOC_56/A 0.29fF
C46635 AND2X1_LOC_508/B AND2X1_LOC_858/B 0.00fF
C46636 OR2X1_LOC_481/Y AND2X1_LOC_789/Y 0.02fF
C46637 VDD AND2X1_LOC_96/a_8_24# 0.00fF
C46638 OR2X1_LOC_237/a_8_216# OR2X1_LOC_428/A 0.05fF
C46639 AND2X1_LOC_70/Y OR2X1_LOC_168/B 0.01fF
C46640 OR2X1_LOC_132/a_8_216# OR2X1_LOC_91/A 0.03fF
C46641 AND2X1_LOC_810/Y AND2X1_LOC_796/A 0.11fF
C46642 AND2X1_LOC_86/B AND2X1_LOC_235/a_8_24# 0.00fF
C46643 OR2X1_LOC_135/Y OR2X1_LOC_619/Y 0.10fF
C46644 OR2X1_LOC_185/Y OR2X1_LOC_267/Y 0.03fF
C46645 AND2X1_LOC_722/a_8_24# AND2X1_LOC_168/a_8_24# 0.23fF
C46646 AND2X1_LOC_72/B AND2X1_LOC_497/a_8_24# 0.04fF
C46647 OR2X1_LOC_185/A OR2X1_LOC_740/B 0.03fF
C46648 OR2X1_LOC_36/Y AND2X1_LOC_473/Y 0.00fF
C46649 AND2X1_LOC_191/a_8_24# OR2X1_LOC_613/Y 0.01fF
C46650 AND2X1_LOC_211/B OR2X1_LOC_171/Y 0.74fF
C46651 AND2X1_LOC_123/Y OR2X1_LOC_12/Y 0.03fF
C46652 AND2X1_LOC_72/Y OR2X1_LOC_549/A 0.01fF
C46653 OR2X1_LOC_121/Y OR2X1_LOC_116/A 0.01fF
C46654 OR2X1_LOC_36/Y OR2X1_LOC_816/A 0.19fF
C46655 OR2X1_LOC_709/A AND2X1_LOC_59/Y 0.07fF
C46656 AND2X1_LOC_477/a_8_24# AND2X1_LOC_469/B 0.01fF
C46657 AND2X1_LOC_564/A AND2X1_LOC_564/a_36_24# 0.00fF
C46658 OR2X1_LOC_785/B AND2X1_LOC_18/Y 0.09fF
C46659 AND2X1_LOC_660/A AND2X1_LOC_216/a_36_24# 0.00fF
C46660 AND2X1_LOC_59/Y AND2X1_LOC_295/a_8_24# 0.20fF
C46661 AND2X1_LOC_787/A OR2X1_LOC_91/a_36_216# 0.00fF
C46662 OR2X1_LOC_36/Y OR2X1_LOC_79/Y 0.01fF
C46663 INPUT_5 AND2X1_LOC_2/Y 0.04fF
C46664 OR2X1_LOC_145/a_8_216# AND2X1_LOC_213/B 0.01fF
C46665 OR2X1_LOC_6/B OR2X1_LOC_394/Y 0.08fF
C46666 AND2X1_LOC_773/Y AND2X1_LOC_702/Y 0.03fF
C46667 AND2X1_LOC_544/Y AND2X1_LOC_147/Y 0.03fF
C46668 AND2X1_LOC_319/A AND2X1_LOC_810/B 0.08fF
C46669 AND2X1_LOC_64/Y AND2X1_LOC_42/B 0.14fF
C46670 AND2X1_LOC_858/B AND2X1_LOC_850/A 0.08fF
C46671 OR2X1_LOC_738/A OR2X1_LOC_711/a_8_216# 0.01fF
C46672 OR2X1_LOC_756/B OR2X1_LOC_624/Y 0.02fF
C46673 OR2X1_LOC_109/Y AND2X1_LOC_778/Y 0.00fF
C46674 OR2X1_LOC_315/Y AND2X1_LOC_476/Y 0.09fF
C46675 AND2X1_LOC_564/A OR2X1_LOC_189/Y 21.49fF
C46676 OR2X1_LOC_121/Y OR2X1_LOC_217/Y 0.02fF
C46677 OR2X1_LOC_105/a_36_216# OR2X1_LOC_78/A 0.03fF
C46678 OR2X1_LOC_56/A OR2X1_LOC_16/Y 0.13fF
C46679 OR2X1_LOC_814/A OR2X1_LOC_593/B 0.01fF
C46680 OR2X1_LOC_405/A OR2X1_LOC_733/A 0.05fF
C46681 AND2X1_LOC_12/Y OR2X1_LOC_362/A 0.05fF
C46682 AND2X1_LOC_831/a_36_24# OR2X1_LOC_12/Y 0.01fF
C46683 OR2X1_LOC_270/a_8_216# OR2X1_LOC_549/A 0.01fF
C46684 AND2X1_LOC_805/Y OR2X1_LOC_627/Y 0.70fF
C46685 OR2X1_LOC_155/A AND2X1_LOC_44/Y 0.94fF
C46686 OR2X1_LOC_9/Y AND2X1_LOC_838/Y 0.03fF
C46687 AND2X1_LOC_564/A OR2X1_LOC_152/Y 0.14fF
C46688 OR2X1_LOC_158/A AND2X1_LOC_114/a_36_24# 0.00fF
C46689 OR2X1_LOC_691/B OR2X1_LOC_269/B 0.01fF
C46690 OR2X1_LOC_564/B OR2X1_LOC_564/a_8_216# 0.00fF
C46691 AND2X1_LOC_658/A OR2X1_LOC_427/A 1.79fF
C46692 OR2X1_LOC_715/B OR2X1_LOC_130/A 0.10fF
C46693 OR2X1_LOC_109/Y AND2X1_LOC_325/a_8_24# 0.01fF
C46694 AND2X1_LOC_95/Y OR2X1_LOC_35/a_8_216# 0.01fF
C46695 AND2X1_LOC_785/a_8_24# OR2X1_LOC_527/Y 0.01fF
C46696 AND2X1_LOC_721/Y OR2X1_LOC_371/Y 0.00fF
C46697 OR2X1_LOC_851/B OR2X1_LOC_87/A 0.01fF
C46698 OR2X1_LOC_26/Y AND2X1_LOC_212/Y 0.10fF
C46699 OR2X1_LOC_51/Y AND2X1_LOC_850/Y 0.04fF
C46700 AND2X1_LOC_456/Y AND2X1_LOC_456/a_36_24# 0.00fF
C46701 AND2X1_LOC_367/A OR2X1_LOC_103/Y 0.03fF
C46702 OR2X1_LOC_677/a_36_216# OR2X1_LOC_677/Y 0.00fF
C46703 VDD OR2X1_LOC_595/a_8_216# 0.21fF
C46704 AND2X1_LOC_508/B AND2X1_LOC_573/A 0.02fF
C46705 OR2X1_LOC_808/B OR2X1_LOC_808/A 0.05fF
C46706 OR2X1_LOC_491/a_8_216# OR2X1_LOC_36/Y 0.02fF
C46707 AND2X1_LOC_361/a_8_24# AND2X1_LOC_361/A 0.07fF
C46708 AND2X1_LOC_81/B OR2X1_LOC_6/B 0.04fF
C46709 OR2X1_LOC_190/A OR2X1_LOC_161/A 0.03fF
C46710 OR2X1_LOC_600/A AND2X1_LOC_848/Y 0.03fF
C46711 AND2X1_LOC_714/B OR2X1_LOC_418/Y 0.01fF
C46712 AND2X1_LOC_50/a_8_24# D_INPUT_4 0.02fF
C46713 OR2X1_LOC_589/A OR2X1_LOC_262/a_36_216# 0.00fF
C46714 AND2X1_LOC_364/A INPUT_0 0.17fF
C46715 OR2X1_LOC_7/A AND2X1_LOC_828/a_8_24# 0.06fF
C46716 AND2X1_LOC_67/Y AND2X1_LOC_7/B 0.18fF
C46717 OR2X1_LOC_155/A OR2X1_LOC_514/a_8_216# 0.03fF
C46718 AND2X1_LOC_564/A OR2X1_LOC_527/Y 0.03fF
C46719 AND2X1_LOC_508/a_8_24# AND2X1_LOC_573/A 0.01fF
C46720 AND2X1_LOC_562/B OR2X1_LOC_92/Y 0.03fF
C46721 OR2X1_LOC_542/B OR2X1_LOC_375/A 0.03fF
C46722 OR2X1_LOC_89/A AND2X1_LOC_212/Y 0.07fF
C46723 D_INPUT_3 AND2X1_LOC_247/a_36_24# 0.01fF
C46724 AND2X1_LOC_59/Y AND2X1_LOC_70/Y 0.31fF
C46725 OR2X1_LOC_3/Y OR2X1_LOC_766/a_8_216# 0.02fF
C46726 AND2X1_LOC_621/Y OR2X1_LOC_442/Y 0.02fF
C46727 OR2X1_LOC_273/a_8_216# AND2X1_LOC_786/Y 0.01fF
C46728 OR2X1_LOC_377/A AND2X1_LOC_92/Y 0.04fF
C46729 AND2X1_LOC_737/Y OR2X1_LOC_441/Y 0.52fF
C46730 OR2X1_LOC_109/a_36_216# AND2X1_LOC_471/Y 0.02fF
C46731 OR2X1_LOC_680/A AND2X1_LOC_806/a_36_24# 0.01fF
C46732 OR2X1_LOC_528/a_8_216# AND2X1_LOC_474/Y 0.01fF
C46733 AND2X1_LOC_562/Y AND2X1_LOC_570/a_8_24# 0.17fF
C46734 AND2X1_LOC_605/Y OR2X1_LOC_48/B 0.01fF
C46735 AND2X1_LOC_566/a_36_24# AND2X1_LOC_566/B 0.01fF
C46736 VDD OR2X1_LOC_267/a_8_216# 0.00fF
C46737 OR2X1_LOC_96/Y OR2X1_LOC_43/A 0.04fF
C46738 AND2X1_LOC_738/B OR2X1_LOC_680/A 0.03fF
C46739 OR2X1_LOC_40/Y AND2X1_LOC_716/a_36_24# 0.00fF
C46740 AND2X1_LOC_399/a_8_24# AND2X1_LOC_18/Y 0.01fF
C46741 OR2X1_LOC_680/A OR2X1_LOC_56/A 0.06fF
C46742 AND2X1_LOC_824/B AND2X1_LOC_92/Y 0.09fF
C46743 AND2X1_LOC_798/Y AND2X1_LOC_802/Y 0.16fF
C46744 AND2X1_LOC_711/a_8_24# AND2X1_LOC_848/Y 0.04fF
C46745 OR2X1_LOC_744/A AND2X1_LOC_655/A 0.03fF
C46746 OR2X1_LOC_662/A OR2X1_LOC_662/a_8_216# 0.01fF
C46747 OR2X1_LOC_641/Y OR2X1_LOC_87/B 0.07fF
C46748 OR2X1_LOC_436/Y OR2X1_LOC_319/Y 0.14fF
C46749 OR2X1_LOC_35/B OR2X1_LOC_35/A 0.06fF
C46750 OR2X1_LOC_241/Y OR2X1_LOC_130/a_8_216# 0.01fF
C46751 AND2X1_LOC_719/Y AND2X1_LOC_719/a_8_24# 0.01fF
C46752 AND2X1_LOC_523/Y OR2X1_LOC_522/a_8_216# 0.01fF
C46753 OR2X1_LOC_158/A OR2X1_LOC_74/A 1.31fF
C46754 OR2X1_LOC_328/a_8_216# INPUT_4 0.07fF
C46755 OR2X1_LOC_532/B OR2X1_LOC_140/B 0.03fF
C46756 OR2X1_LOC_808/B OR2X1_LOC_732/a_8_216# 0.30fF
C46757 OR2X1_LOC_214/a_8_216# OR2X1_LOC_66/A 0.01fF
C46758 OR2X1_LOC_250/Y OR2X1_LOC_251/a_8_216# 0.01fF
C46759 AND2X1_LOC_712/a_8_24# AND2X1_LOC_712/B 0.09fF
C46760 AND2X1_LOC_784/A OR2X1_LOC_426/B 0.16fF
C46761 AND2X1_LOC_850/A AND2X1_LOC_573/A 0.03fF
C46762 OR2X1_LOC_691/a_8_216# AND2X1_LOC_51/Y 0.01fF
C46763 OR2X1_LOC_203/Y AND2X1_LOC_92/Y 0.01fF
C46764 AND2X1_LOC_583/a_36_24# OR2X1_LOC_639/B 0.01fF
C46765 AND2X1_LOC_59/Y OR2X1_LOC_703/A 0.00fF
C46766 AND2X1_LOC_559/a_8_24# AND2X1_LOC_218/Y 0.17fF
C46767 OR2X1_LOC_91/Y AND2X1_LOC_474/A 0.02fF
C46768 AND2X1_LOC_753/B AND2X1_LOC_753/a_8_24# 0.02fF
C46769 OR2X1_LOC_468/A OR2X1_LOC_810/A 0.04fF
C46770 AND2X1_LOC_56/B OR2X1_LOC_78/B 0.09fF
C46771 AND2X1_LOC_141/a_8_24# OR2X1_LOC_26/Y 0.03fF
C46772 AND2X1_LOC_70/Y AND2X1_LOC_495/a_8_24# 0.01fF
C46773 OR2X1_LOC_859/A OR2X1_LOC_576/A 0.44fF
C46774 OR2X1_LOC_207/B AND2X1_LOC_48/A 0.03fF
C46775 AND2X1_LOC_251/a_36_24# OR2X1_LOC_561/Y 0.00fF
C46776 OR2X1_LOC_22/a_8_216# OR2X1_LOC_25/Y 0.02fF
C46777 OR2X1_LOC_158/A OR2X1_LOC_261/A 0.01fF
C46778 OR2X1_LOC_644/B INPUT_0 -0.02fF
C46779 AND2X1_LOC_691/a_36_24# OR2X1_LOC_753/A 0.01fF
C46780 AND2X1_LOC_350/a_8_24# AND2X1_LOC_351/Y 0.01fF
C46781 AND2X1_LOC_570/Y OR2X1_LOC_239/a_8_216# 0.01fF
C46782 AND2X1_LOC_8/Y OR2X1_LOC_78/B 0.20fF
C46783 AND2X1_LOC_339/B OR2X1_LOC_416/Y 0.00fF
C46784 AND2X1_LOC_366/a_8_24# OR2X1_LOC_89/A 0.01fF
C46785 AND2X1_LOC_769/a_8_24# OR2X1_LOC_426/B 0.12fF
C46786 OR2X1_LOC_604/A OR2X1_LOC_282/Y 0.05fF
C46787 OR2X1_LOC_91/Y AND2X1_LOC_733/a_8_24# 0.03fF
C46788 OR2X1_LOC_312/Y AND2X1_LOC_434/Y 0.07fF
C46789 AND2X1_LOC_589/a_8_24# OR2X1_LOC_468/A 0.01fF
C46790 AND2X1_LOC_141/a_8_24# OR2X1_LOC_89/A 0.01fF
C46791 OR2X1_LOC_405/A OR2X1_LOC_730/a_8_216# 0.01fF
C46792 OR2X1_LOC_600/A OR2X1_LOC_617/Y 0.03fF
C46793 OR2X1_LOC_532/B OR2X1_LOC_355/A 0.01fF
C46794 OR2X1_LOC_329/B OR2X1_LOC_280/a_8_216# 0.03fF
C46795 INPUT_1 OR2X1_LOC_548/a_8_216# 0.06fF
C46796 D_INPUT_0 OR2X1_LOC_548/B 0.01fF
C46797 OR2X1_LOC_235/B OR2X1_LOC_585/A 0.11fF
C46798 AND2X1_LOC_50/Y AND2X1_LOC_25/Y 1.21fF
C46799 OR2X1_LOC_231/A OR2X1_LOC_215/Y 0.02fF
C46800 AND2X1_LOC_679/a_8_24# AND2X1_LOC_36/Y 0.01fF
C46801 OR2X1_LOC_231/A AND2X1_LOC_230/a_36_24# 0.00fF
C46802 OR2X1_LOC_232/a_8_216# OR2X1_LOC_234/Y 0.40fF
C46803 AND2X1_LOC_753/B OR2X1_LOC_194/Y 0.05fF
C46804 AND2X1_LOC_78/a_8_24# OR2X1_LOC_59/Y 0.01fF
C46805 OR2X1_LOC_3/Y OR2X1_LOC_122/A 0.01fF
C46806 OR2X1_LOC_659/B OR2X1_LOC_721/Y 0.02fF
C46807 AND2X1_LOC_175/B OR2X1_LOC_619/Y 0.00fF
C46808 VDD OR2X1_LOC_431/a_8_216# 0.21fF
C46809 OR2X1_LOC_3/Y INPUT_0 0.10fF
C46810 OR2X1_LOC_318/B OR2X1_LOC_776/A 0.02fF
C46811 AND2X1_LOC_318/a_8_24# OR2X1_LOC_18/Y 0.04fF
C46812 OR2X1_LOC_186/Y AND2X1_LOC_47/Y 0.03fF
C46813 OR2X1_LOC_720/a_36_216# OR2X1_LOC_721/Y 0.00fF
C46814 AND2X1_LOC_170/B AND2X1_LOC_810/B 0.07fF
C46815 OR2X1_LOC_36/Y AND2X1_LOC_649/a_8_24# 0.01fF
C46816 OR2X1_LOC_45/Y OR2X1_LOC_36/Y 0.30fF
C46817 OR2X1_LOC_145/Y AND2X1_LOC_213/B 0.01fF
C46818 AND2X1_LOC_864/a_8_24# AND2X1_LOC_212/Y 0.01fF
C46819 OR2X1_LOC_62/A OR2X1_LOC_15/a_8_216# 0.11fF
C46820 INPUT_3 OR2X1_LOC_618/a_8_216# 0.01fF
C46821 AND2X1_LOC_42/B AND2X1_LOC_819/a_8_24# 0.01fF
C46822 OR2X1_LOC_366/A OR2X1_LOC_366/a_8_216# 0.39fF
C46823 VDD OR2X1_LOC_443/Y 0.12fF
C46824 AND2X1_LOC_94/a_8_24# AND2X1_LOC_56/B 0.13fF
C46825 OR2X1_LOC_71/a_8_216# OR2X1_LOC_6/A 0.06fF
C46826 OR2X1_LOC_539/Y OR2X1_LOC_799/a_8_216# 0.01fF
C46827 OR2X1_LOC_538/A AND2X1_LOC_111/a_36_24# 0.00fF
C46828 OR2X1_LOC_130/A OR2X1_LOC_215/Y 0.00fF
C46829 D_INPUT_0 OR2X1_LOC_786/A 0.03fF
C46830 OR2X1_LOC_502/A AND2X1_LOC_3/Y 0.37fF
C46831 AND2X1_LOC_164/a_8_24# AND2X1_LOC_51/Y 0.15fF
C46832 OR2X1_LOC_446/B OR2X1_LOC_515/Y 0.14fF
C46833 OR2X1_LOC_432/Y OR2X1_LOC_44/Y 0.37fF
C46834 OR2X1_LOC_502/A OR2X1_LOC_647/B 0.01fF
C46835 OR2X1_LOC_160/A OR2X1_LOC_87/A 0.22fF
C46836 OR2X1_LOC_838/a_8_216# OR2X1_LOC_20/a_8_216# 0.47fF
C46837 OR2X1_LOC_648/A OR2X1_LOC_750/A 0.00fF
C46838 OR2X1_LOC_18/Y AND2X1_LOC_361/A 0.07fF
C46839 AND2X1_LOC_719/Y OR2X1_LOC_31/Y 0.02fF
C46840 OR2X1_LOC_287/B OR2X1_LOC_811/A 0.03fF
C46841 AND2X1_LOC_430/B AND2X1_LOC_582/B 0.01fF
C46842 AND2X1_LOC_12/Y D_GATE_865 0.00fF
C46843 AND2X1_LOC_354/a_8_24# AND2X1_LOC_319/A 0.03fF
C46844 OR2X1_LOC_243/a_8_216# OR2X1_LOC_66/A 0.01fF
C46845 AND2X1_LOC_56/B OR2X1_LOC_375/A 0.11fF
C46846 OR2X1_LOC_53/Y OR2X1_LOC_41/Y 0.00fF
C46847 AND2X1_LOC_664/a_8_24# AND2X1_LOC_663/A 0.15fF
C46848 OR2X1_LOC_598/A OR2X1_LOC_338/A 0.07fF
C46849 OR2X1_LOC_417/A AND2X1_LOC_489/a_8_24# 0.01fF
C46850 AND2X1_LOC_806/A OR2X1_LOC_39/A 0.06fF
C46851 AND2X1_LOC_566/B AND2X1_LOC_318/Y 0.02fF
C46852 AND2X1_LOC_566/B AND2X1_LOC_864/a_36_24# 0.00fF
C46853 OR2X1_LOC_849/A OR2X1_LOC_659/a_8_216# 0.01fF
C46854 OR2X1_LOC_419/Y OR2X1_LOC_816/A 0.03fF
C46855 AND2X1_LOC_8/Y OR2X1_LOC_375/A 0.45fF
C46856 AND2X1_LOC_838/Y AND2X1_LOC_852/Y 0.00fF
C46857 AND2X1_LOC_50/Y AND2X1_LOC_51/Y 0.84fF
C46858 OR2X1_LOC_26/Y OR2X1_LOC_265/Y 0.08fF
C46859 OR2X1_LOC_160/A AND2X1_LOC_19/a_8_24# 0.01fF
C46860 OR2X1_LOC_831/B OR2X1_LOC_228/Y 0.02fF
C46861 AND2X1_LOC_3/Y AND2X1_LOC_230/a_8_24# 0.02fF
C46862 AND2X1_LOC_170/a_8_24# AND2X1_LOC_566/Y 0.03fF
C46863 OR2X1_LOC_784/a_36_216# OR2X1_LOC_161/A 0.01fF
C46864 AND2X1_LOC_356/B AND2X1_LOC_436/B 0.07fF
C46865 OR2X1_LOC_216/Y OR2X1_LOC_218/a_8_216# 0.05fF
C46866 OR2X1_LOC_36/Y OR2X1_LOC_824/Y 0.01fF
C46867 AND2X1_LOC_363/Y AND2X1_LOC_866/A 0.06fF
C46868 AND2X1_LOC_319/A OR2X1_LOC_585/A 0.02fF
C46869 AND2X1_LOC_148/Y OR2X1_LOC_679/B 0.05fF
C46870 OR2X1_LOC_36/Y OR2X1_LOC_591/a_8_216# 0.01fF
C46871 OR2X1_LOC_696/a_8_216# OR2X1_LOC_39/A 0.06fF
C46872 AND2X1_LOC_84/a_8_24# OR2X1_LOC_80/Y 0.08fF
C46873 AND2X1_LOC_729/Y OR2X1_LOC_743/A 0.15fF
C46874 OR2X1_LOC_76/A OR2X1_LOC_811/A 1.97fF
C46875 AND2X1_LOC_276/Y OR2X1_LOC_39/A 0.02fF
C46876 OR2X1_LOC_3/Y OR2X1_LOC_11/Y 0.34fF
C46877 OR2X1_LOC_786/Y AND2X1_LOC_18/Y 0.03fF
C46878 OR2X1_LOC_75/a_8_216# AND2X1_LOC_219/Y 0.03fF
C46879 OR2X1_LOC_491/a_8_216# OR2X1_LOC_419/Y 0.12fF
C46880 AND2X1_LOC_67/Y OR2X1_LOC_805/A 0.03fF
C46881 OR2X1_LOC_329/B AND2X1_LOC_476/A 0.07fF
C46882 OR2X1_LOC_8/Y D_INPUT_1 0.13fF
C46883 OR2X1_LOC_417/Y AND2X1_LOC_593/Y 0.07fF
C46884 OR2X1_LOC_6/B OR2X1_LOC_66/Y 0.01fF
C46885 OR2X1_LOC_40/Y AND2X1_LOC_793/Y 0.37fF
C46886 AND2X1_LOC_135/a_36_24# OR2X1_LOC_161/A 0.00fF
C46887 OR2X1_LOC_850/B AND2X1_LOC_283/a_36_24# 0.00fF
C46888 AND2X1_LOC_784/A OR2X1_LOC_743/A 0.06fF
C46889 AND2X1_LOC_863/A OR2X1_LOC_619/Y 0.01fF
C46890 AND2X1_LOC_474/A D_INPUT_3 0.03fF
C46891 INPUT_0 OR2X1_LOC_673/A 0.03fF
C46892 OR2X1_LOC_604/A AND2X1_LOC_259/a_8_24# 0.06fF
C46893 OR2X1_LOC_3/Y OR2X1_LOC_690/A 0.16fF
C46894 OR2X1_LOC_485/Y AND2X1_LOC_486/a_8_24# 0.05fF
C46895 AND2X1_LOC_72/a_8_24# AND2X1_LOC_3/Y 0.02fF
C46896 OR2X1_LOC_384/a_36_216# OR2X1_LOC_428/A 0.00fF
C46897 OR2X1_LOC_22/Y AND2X1_LOC_436/B 0.07fF
C46898 OR2X1_LOC_280/Y OR2X1_LOC_529/Y 0.03fF
C46899 AND2X1_LOC_456/B OR2X1_LOC_615/Y 0.03fF
C46900 OR2X1_LOC_291/Y OR2X1_LOC_85/A 0.06fF
C46901 AND2X1_LOC_792/B AND2X1_LOC_792/a_8_24# 0.01fF
C46902 OR2X1_LOC_70/Y AND2X1_LOC_100/a_36_24# 0.00fF
C46903 OR2X1_LOC_22/Y AND2X1_LOC_287/a_36_24# 0.01fF
C46904 OR2X1_LOC_43/A OR2X1_LOC_829/Y 0.02fF
C46905 AND2X1_LOC_703/Y OR2X1_LOC_589/Y 0.00fF
C46906 AND2X1_LOC_48/A OR2X1_LOC_350/a_8_216# 0.02fF
C46907 OR2X1_LOC_361/a_36_216# OR2X1_LOC_560/A 0.03fF
C46908 OR2X1_LOC_22/Y AND2X1_LOC_139/B 0.07fF
C46909 OR2X1_LOC_624/A D_INPUT_0 0.24fF
C46910 OR2X1_LOC_787/Y OR2X1_LOC_794/a_36_216# 0.02fF
C46911 OR2X1_LOC_426/B AND2X1_LOC_643/a_8_24# 0.02fF
C46912 OR2X1_LOC_837/A AND2X1_LOC_472/a_8_24# 0.21fF
C46913 OR2X1_LOC_3/Y OR2X1_LOC_272/a_8_216# 0.01fF
C46914 OR2X1_LOC_22/Y OR2X1_LOC_767/a_36_216# 0.02fF
C46915 AND2X1_LOC_48/A OR2X1_LOC_790/a_8_216# 0.01fF
C46916 OR2X1_LOC_66/A AND2X1_LOC_52/Y 0.03fF
C46917 OR2X1_LOC_441/Y AND2X1_LOC_808/A 0.03fF
C46918 OR2X1_LOC_36/Y AND2X1_LOC_727/A 0.04fF
C46919 AND2X1_LOC_110/Y AND2X1_LOC_31/Y 0.04fF
C46920 D_INPUT_3 OR2X1_LOC_818/Y 0.01fF
C46921 OR2X1_LOC_62/A AND2X1_LOC_414/a_8_24# 0.04fF
C46922 OR2X1_LOC_686/a_8_216# AND2X1_LOC_430/B 0.01fF
C46923 OR2X1_LOC_810/A OR2X1_LOC_121/B 0.03fF
C46924 OR2X1_LOC_320/Y OR2X1_LOC_321/Y 0.19fF
C46925 AND2X1_LOC_784/A OR2X1_LOC_246/A 0.30fF
C46926 OR2X1_LOC_643/A OR2X1_LOC_474/a_36_216# 0.00fF
C46927 OR2X1_LOC_389/A OR2X1_LOC_750/Y 0.02fF
C46928 OR2X1_LOC_426/B OR2X1_LOC_88/Y 0.19fF
C46929 OR2X1_LOC_293/a_36_216# OR2X1_LOC_585/A 0.00fF
C46930 OR2X1_LOC_19/B OR2X1_LOC_240/A 3.24fF
C46931 OR2X1_LOC_43/A OR2X1_LOC_7/Y 0.02fF
C46932 OR2X1_LOC_473/A OR2X1_LOC_493/A 0.19fF
C46933 OR2X1_LOC_3/Y OR2X1_LOC_64/Y 0.38fF
C46934 OR2X1_LOC_47/Y OR2X1_LOC_278/Y 0.02fF
C46935 AND2X1_LOC_34/Y AND2X1_LOC_472/a_8_24# 0.17fF
C46936 OR2X1_LOC_139/a_36_216# OR2X1_LOC_62/B 0.00fF
C46937 AND2X1_LOC_48/A AND2X1_LOC_3/Y 0.29fF
C46938 OR2X1_LOC_767/Y AND2X1_LOC_772/Y 0.01fF
C46939 OR2X1_LOC_473/Y OR2X1_LOC_206/a_36_216# 0.00fF
C46940 OR2X1_LOC_529/Y OR2X1_LOC_22/Y 0.03fF
C46941 OR2X1_LOC_36/Y OR2X1_LOC_95/Y 0.05fF
C46942 OR2X1_LOC_334/A OR2X1_LOC_334/a_8_216# 0.00fF
C46943 OR2X1_LOC_473/Y AND2X1_LOC_51/Y 0.15fF
C46944 AND2X1_LOC_866/A OR2X1_LOC_236/a_36_216# 0.14fF
C46945 AND2X1_LOC_1/Y OR2X1_LOC_639/A 0.01fF
C46946 AND2X1_LOC_471/a_8_24# OR2X1_LOC_371/Y 0.01fF
C46947 D_INPUT_3 OR2X1_LOC_85/A 0.06fF
C46948 OR2X1_LOC_36/Y OR2X1_LOC_368/A 0.01fF
C46949 INPUT_0 AND2X1_LOC_409/a_8_24# 0.01fF
C46950 OR2X1_LOC_548/A AND2X1_LOC_36/Y 0.01fF
C46951 OR2X1_LOC_214/B OR2X1_LOC_161/A 0.17fF
C46952 OR2X1_LOC_486/Y AND2X1_LOC_36/Y 0.15fF
C46953 OR2X1_LOC_18/Y AND2X1_LOC_795/Y 0.11fF
C46954 AND2X1_LOC_489/Y OR2X1_LOC_71/Y 0.01fF
C46955 OR2X1_LOC_161/A OR2X1_LOC_241/B 0.01fF
C46956 OR2X1_LOC_711/a_8_216# AND2X1_LOC_36/Y 0.01fF
C46957 OR2X1_LOC_394/Y OR2X1_LOC_598/A 0.02fF
C46958 OR2X1_LOC_596/A OR2X1_LOC_703/Y 0.42fF
C46959 OR2X1_LOC_744/Y AND2X1_LOC_780/a_8_24# 0.01fF
C46960 OR2X1_LOC_352/A OR2X1_LOC_578/B 0.01fF
C46961 OR2X1_LOC_110/a_8_216# AND2X1_LOC_786/Y 0.01fF
C46962 OR2X1_LOC_499/a_8_216# OR2X1_LOC_493/Y 0.28fF
C46963 OR2X1_LOC_3/Y OR2X1_LOC_417/A 0.49fF
C46964 AND2X1_LOC_632/A AND2X1_LOC_631/Y 0.19fF
C46965 AND2X1_LOC_769/a_8_24# OR2X1_LOC_409/B 0.01fF
C46966 AND2X1_LOC_476/Y AND2X1_LOC_269/a_8_24# 0.20fF
C46967 AND2X1_LOC_807/Y OR2X1_LOC_419/Y 0.13fF
C46968 OR2X1_LOC_34/A OR2X1_LOC_338/A 0.01fF
C46969 OR2X1_LOC_211/a_8_216# OR2X1_LOC_170/Y 0.00fF
C46970 AND2X1_LOC_434/Y OR2X1_LOC_13/B 2.24fF
C46971 OR2X1_LOC_506/A OR2X1_LOC_728/B 0.09fF
C46972 OR2X1_LOC_449/A OR2X1_LOC_779/Y 0.01fF
C46973 AND2X1_LOC_219/Y OR2X1_LOC_13/B 0.07fF
C46974 OR2X1_LOC_443/Y OR2X1_LOC_444/B 0.16fF
C46975 OR2X1_LOC_8/Y AND2X1_LOC_789/Y 0.01fF
C46976 OR2X1_LOC_52/B AND2X1_LOC_770/a_36_24# 0.01fF
C46977 AND2X1_LOC_687/a_8_24# OR2X1_LOC_7/A 0.03fF
C46978 AND2X1_LOC_81/B OR2X1_LOC_598/A 0.01fF
C46979 OR2X1_LOC_344/A OR2X1_LOC_562/A 0.00fF
C46980 AND2X1_LOC_49/a_8_24# OR2X1_LOC_598/A 0.04fF
C46981 AND2X1_LOC_721/A OR2X1_LOC_585/A 0.06fF
C46982 AND2X1_LOC_739/B AND2X1_LOC_803/B 0.35fF
C46983 OR2X1_LOC_368/a_8_216# OR2X1_LOC_696/A 0.01fF
C46984 INPUT_1 OR2X1_LOC_46/A 1.18fF
C46985 AND2X1_LOC_462/B OR2X1_LOC_690/A 0.01fF
C46986 D_INPUT_0 OR2X1_LOC_54/Y 0.41fF
C46987 OR2X1_LOC_16/A OR2X1_LOC_312/a_8_216# 0.01fF
C46988 AND2X1_LOC_92/Y OR2X1_LOC_539/B 0.04fF
C46989 OR2X1_LOC_115/a_36_216# OR2X1_LOC_560/A 0.00fF
C46990 OR2X1_LOC_429/Y OR2X1_LOC_51/a_8_216# 0.03fF
C46991 AND2X1_LOC_40/Y OR2X1_LOC_366/Y 0.03fF
C46992 VDD AND2X1_LOC_409/B 0.08fF
C46993 OR2X1_LOC_655/B OR2X1_LOC_649/a_8_216# 0.04fF
C46994 OR2X1_LOC_285/Y OR2X1_LOC_286/a_8_216# 0.39fF
C46995 OR2X1_LOC_473/Y OR2X1_LOC_201/a_36_216# 0.00fF
C46996 AND2X1_LOC_44/Y OR2X1_LOC_706/a_36_216# 0.00fF
C46997 OR2X1_LOC_196/B AND2X1_LOC_47/Y 0.07fF
C46998 VDD OR2X1_LOC_605/Y 0.23fF
C46999 VDD AND2X1_LOC_763/B 0.30fF
C47000 OR2X1_LOC_756/B OR2X1_LOC_174/Y 0.43fF
C47001 OR2X1_LOC_485/A AND2X1_LOC_644/a_8_24# 0.02fF
C47002 OR2X1_LOC_243/a_36_216# OR2X1_LOC_244/A 0.01fF
C47003 OR2X1_LOC_691/Y OR2X1_LOC_185/a_36_216# 0.00fF
C47004 OR2X1_LOC_506/Y OR2X1_LOC_508/a_8_216# 0.00fF
C47005 OR2X1_LOC_156/A AND2X1_LOC_7/B 0.35fF
C47006 AND2X1_LOC_555/Y AND2X1_LOC_285/Y 0.01fF
C47007 OR2X1_LOC_743/A AND2X1_LOC_643/a_8_24# 0.05fF
C47008 AND2X1_LOC_41/A OR2X1_LOC_508/Y 0.03fF
C47009 OR2X1_LOC_45/B AND2X1_LOC_448/a_8_24# 0.02fF
C47010 OR2X1_LOC_19/B OR2X1_LOC_47/Y 0.08fF
C47011 OR2X1_LOC_604/A AND2X1_LOC_287/B 0.09fF
C47012 AND2X1_LOC_810/A OR2X1_LOC_158/A 0.03fF
C47013 OR2X1_LOC_421/A AND2X1_LOC_707/Y 0.04fF
C47014 AND2X1_LOC_573/A OR2X1_LOC_399/Y 0.01fF
C47015 AND2X1_LOC_729/Y OR2X1_LOC_599/a_8_216# 0.47fF
C47016 OR2X1_LOC_604/A OR2X1_LOC_816/A 0.03fF
C47017 OR2X1_LOC_381/a_8_216# OR2X1_LOC_382/A 0.01fF
C47018 OR2X1_LOC_185/a_8_216# OR2X1_LOC_729/a_8_216# 0.47fF
C47019 OR2X1_LOC_840/a_8_216# OR2X1_LOC_851/B 0.03fF
C47020 OR2X1_LOC_276/a_8_216# D_INPUT_0 0.03fF
C47021 VDD AND2X1_LOC_636/a_8_24# -0.00fF
C47022 AND2X1_LOC_474/Y AND2X1_LOC_657/A 0.00fF
C47023 OR2X1_LOC_78/A OR2X1_LOC_554/a_8_216# 0.01fF
C47024 OR2X1_LOC_175/Y OR2X1_LOC_35/Y 0.02fF
C47025 OR2X1_LOC_508/A OR2X1_LOC_508/Y 0.01fF
C47026 OR2X1_LOC_549/A OR2X1_LOC_719/B 0.02fF
C47027 OR2X1_LOC_576/A OR2X1_LOC_66/A 0.05fF
C47028 OR2X1_LOC_47/Y AND2X1_LOC_800/a_8_24# 0.01fF
C47029 AND2X1_LOC_725/a_8_24# OR2X1_LOC_12/Y 0.01fF
C47030 AND2X1_LOC_18/Y AND2X1_LOC_255/a_8_24# 0.01fF
C47031 OR2X1_LOC_833/Y OR2X1_LOC_6/B 0.01fF
C47032 AND2X1_LOC_574/Y AND2X1_LOC_735/Y 0.02fF
C47033 OR2X1_LOC_485/A AND2X1_LOC_657/A 0.07fF
C47034 AND2X1_LOC_571/a_8_24# AND2X1_LOC_561/B 0.01fF
C47035 OR2X1_LOC_8/Y OR2X1_LOC_15/a_8_216# 0.00fF
C47036 AND2X1_LOC_12/Y OR2X1_LOC_771/B 0.03fF
C47037 AND2X1_LOC_64/Y OR2X1_LOC_663/A 0.03fF
C47038 AND2X1_LOC_727/A OR2X1_LOC_419/Y 0.03fF
C47039 VDD OR2X1_LOC_603/Y 0.12fF
C47040 AND2X1_LOC_539/Y AND2X1_LOC_512/Y 0.70fF
C47041 AND2X1_LOC_586/a_36_24# AND2X1_LOC_36/Y 0.00fF
C47042 AND2X1_LOC_706/Y VDD 0.57fF
C47043 AND2X1_LOC_401/Y OR2X1_LOC_415/Y 0.01fF
C47044 AND2X1_LOC_56/B OR2X1_LOC_515/Y 0.01fF
C47045 OR2X1_LOC_48/B OR2X1_LOC_387/A 0.05fF
C47046 AND2X1_LOC_705/a_36_24# OR2X1_LOC_12/Y 0.01fF
C47047 AND2X1_LOC_732/B OR2X1_LOC_421/Y 0.15fF
C47048 OR2X1_LOC_246/A AND2X1_LOC_643/a_8_24# 0.22fF
C47049 OR2X1_LOC_329/B AND2X1_LOC_445/a_8_24# 0.02fF
C47050 AND2X1_LOC_64/Y AND2X1_LOC_503/a_8_24# 0.01fF
C47051 OR2X1_LOC_158/A AND2X1_LOC_860/A 0.12fF
C47052 D_INPUT_0 OR2X1_LOC_84/Y 0.06fF
C47053 OR2X1_LOC_160/A OR2X1_LOC_844/B 0.02fF
C47054 OR2X1_LOC_22/Y OR2X1_LOC_598/A 0.03fF
C47055 OR2X1_LOC_316/Y OR2X1_LOC_268/Y 0.01fF
C47056 AND2X1_LOC_522/a_8_24# OR2X1_LOC_632/Y 0.03fF
C47057 OR2X1_LOC_254/A OR2X1_LOC_562/A 0.01fF
C47058 OR2X1_LOC_542/B OR2X1_LOC_549/A 0.07fF
C47059 OR2X1_LOC_738/A OR2X1_LOC_308/Y 0.02fF
C47060 OR2X1_LOC_439/B OR2X1_LOC_66/A 0.09fF
C47061 OR2X1_LOC_18/Y OR2X1_LOC_387/A 0.02fF
C47062 OR2X1_LOC_40/Y AND2X1_LOC_357/B 0.02fF
C47063 AND2X1_LOC_12/Y OR2X1_LOC_776/A 0.03fF
C47064 AND2X1_LOC_319/a_36_24# OR2X1_LOC_428/A 0.01fF
C47065 AND2X1_LOC_1/a_8_24# D_INPUT_6 0.01fF
C47066 AND2X1_LOC_229/a_8_24# AND2X1_LOC_41/A 0.08fF
C47067 AND2X1_LOC_555/Y OR2X1_LOC_281/a_36_216# 0.00fF
C47068 OR2X1_LOC_87/A OR2X1_LOC_212/B 0.02fF
C47069 AND2X1_LOC_535/Y AND2X1_LOC_567/a_8_24# 0.10fF
C47070 OR2X1_LOC_71/Y AND2X1_LOC_216/A 0.02fF
C47071 AND2X1_LOC_64/Y OR2X1_LOC_547/B 0.04fF
C47072 OR2X1_LOC_62/B OR2X1_LOC_398/Y 0.03fF
C47073 OR2X1_LOC_97/A OR2X1_LOC_840/A 0.03fF
C47074 OR2X1_LOC_415/A OR2X1_LOC_80/A 0.07fF
C47075 OR2X1_LOC_40/Y AND2X1_LOC_363/Y 0.15fF
C47076 OR2X1_LOC_246/A OR2X1_LOC_88/Y 0.02fF
C47077 OR2X1_LOC_160/A OR2X1_LOC_390/B 0.07fF
C47078 OR2X1_LOC_95/Y OR2X1_LOC_419/Y 0.69fF
C47079 OR2X1_LOC_158/A AND2X1_LOC_162/a_8_24# 0.01fF
C47080 VDD OR2X1_LOC_58/Y 0.11fF
C47081 AND2X1_LOC_727/A OR2X1_LOC_152/A 0.09fF
C47082 AND2X1_LOC_440/a_8_24# OR2X1_LOC_419/Y 0.13fF
C47083 AND2X1_LOC_508/B AND2X1_LOC_806/a_8_24# 0.00fF
C47084 OR2X1_LOC_672/Y AND2X1_LOC_789/Y 0.02fF
C47085 OR2X1_LOC_841/B OR2X1_LOC_776/A 0.05fF
C47086 AND2X1_LOC_347/B OR2X1_LOC_59/Y 0.61fF
C47087 OR2X1_LOC_45/B OR2X1_LOC_23/a_8_216# 0.00fF
C47088 VDD OR2X1_LOC_687/A -0.00fF
C47089 AND2X1_LOC_214/A OR2X1_LOC_13/Y 0.01fF
C47090 AND2X1_LOC_665/a_8_24# OR2X1_LOC_675/Y 0.14fF
C47091 AND2X1_LOC_40/Y OR2X1_LOC_389/a_8_216# 0.14fF
C47092 OR2X1_LOC_40/Y AND2X1_LOC_548/Y 0.14fF
C47093 OR2X1_LOC_8/Y OR2X1_LOC_426/B 0.02fF
C47094 OR2X1_LOC_643/A OR2X1_LOC_510/a_8_216# 0.02fF
C47095 OR2X1_LOC_51/Y AND2X1_LOC_285/Y 0.00fF
C47096 AND2X1_LOC_756/a_8_24# OR2X1_LOC_600/A 0.15fF
C47097 OR2X1_LOC_188/Y OR2X1_LOC_161/A 0.02fF
C47098 OR2X1_LOC_771/a_8_216# D_INPUT_1 0.01fF
C47099 OR2X1_LOC_709/A OR2X1_LOC_623/B 0.03fF
C47100 OR2X1_LOC_364/A AND2X1_LOC_64/Y 0.07fF
C47101 OR2X1_LOC_264/Y AND2X1_LOC_65/A 4.16fF
C47102 AND2X1_LOC_620/Y AND2X1_LOC_623/a_36_24# 0.01fF
C47103 OR2X1_LOC_40/Y AND2X1_LOC_303/a_8_24# 0.02fF
C47104 OR2X1_LOC_185/Y AND2X1_LOC_64/Y 0.24fF
C47105 OR2X1_LOC_70/Y OR2X1_LOC_142/Y 0.03fF
C47106 AND2X1_LOC_84/Y OR2X1_LOC_69/a_8_216# 0.01fF
C47107 OR2X1_LOC_160/B OR2X1_LOC_678/Y 0.00fF
C47108 OR2X1_LOC_385/Y OR2X1_LOC_387/A 0.09fF
C47109 OR2X1_LOC_416/Y OR2X1_LOC_300/Y 0.01fF
C47110 AND2X1_LOC_792/Y AND2X1_LOC_805/a_8_24# 0.04fF
C47111 OR2X1_LOC_158/A AND2X1_LOC_155/a_8_24# 0.01fF
C47112 AND2X1_LOC_322/a_36_24# OR2X1_LOC_703/A 0.00fF
C47113 VDD OR2X1_LOC_634/A 0.64fF
C47114 AND2X1_LOC_486/Y AND2X1_LOC_476/Y 0.07fF
C47115 AND2X1_LOC_553/A AND2X1_LOC_541/Y 0.04fF
C47116 AND2X1_LOC_41/A OR2X1_LOC_66/A 0.17fF
C47117 AND2X1_LOC_191/B AND2X1_LOC_858/B 0.17fF
C47118 OR2X1_LOC_186/Y OR2X1_LOC_506/A 0.03fF
C47119 OR2X1_LOC_78/B AND2X1_LOC_92/Y 0.17fF
C47120 OR2X1_LOC_264/Y OR2X1_LOC_510/A 0.09fF
C47121 OR2X1_LOC_9/Y AND2X1_LOC_852/B 0.01fF
C47122 OR2X1_LOC_486/a_8_216# AND2X1_LOC_36/Y 0.02fF
C47123 OR2X1_LOC_538/a_8_216# VDD 0.21fF
C47124 AND2X1_LOC_713/a_36_24# OR2X1_LOC_48/B 0.01fF
C47125 AND2X1_LOC_720/Y AND2X1_LOC_860/A 0.03fF
C47126 OR2X1_LOC_814/A OR2X1_LOC_580/A 0.14fF
C47127 OR2X1_LOC_597/A OR2X1_LOC_692/a_8_216# 0.47fF
C47128 OR2X1_LOC_421/A OR2X1_LOC_692/a_36_216# 0.00fF
C47129 AND2X1_LOC_743/a_8_24# OR2X1_LOC_87/A 0.04fF
C47130 OR2X1_LOC_66/Y OR2X1_LOC_598/A 0.09fF
C47131 OR2X1_LOC_597/A OR2X1_LOC_92/Y 0.02fF
C47132 OR2X1_LOC_207/B OR2X1_LOC_790/a_8_216# 0.02fF
C47133 OR2X1_LOC_177/Y AND2X1_LOC_807/Y 0.04fF
C47134 AND2X1_LOC_138/a_36_24# OR2X1_LOC_12/Y 0.01fF
C47135 OR2X1_LOC_151/A OR2X1_LOC_739/A 0.03fF
C47136 OR2X1_LOC_179/a_36_216# OR2X1_LOC_178/Y 0.00fF
C47137 OR2X1_LOC_97/B AND2X1_LOC_44/Y 0.21fF
C47138 OR2X1_LOC_339/a_8_216# AND2X1_LOC_40/Y 0.01fF
C47139 VDD AND2X1_LOC_851/A 0.25fF
C47140 OR2X1_LOC_49/A OR2X1_LOC_87/B 0.23fF
C47141 OR2X1_LOC_427/A AND2X1_LOC_614/a_8_24# 0.01fF
C47142 OR2X1_LOC_790/A OR2X1_LOC_377/A 0.00fF
C47143 OR2X1_LOC_160/B OR2X1_LOC_811/A 0.07fF
C47144 OR2X1_LOC_770/A OR2X1_LOC_287/B 0.00fF
C47145 AND2X1_LOC_717/B AND2X1_LOC_242/B 0.02fF
C47146 AND2X1_LOC_702/Y OR2X1_LOC_12/Y 0.15fF
C47147 AND2X1_LOC_553/A OR2X1_LOC_107/a_8_216# 0.01fF
C47148 AND2X1_LOC_340/Y AND2X1_LOC_361/A 0.25fF
C47149 AND2X1_LOC_70/Y OR2X1_LOC_794/A 0.01fF
C47150 AND2X1_LOC_81/B OR2X1_LOC_646/B 0.16fF
C47151 OR2X1_LOC_6/B OR2X1_LOC_39/A 2.65fF
C47152 OR2X1_LOC_426/B AND2X1_LOC_76/Y 0.03fF
C47153 OR2X1_LOC_502/A INPUT_0 1.47fF
C47154 AND2X1_LOC_56/B OR2X1_LOC_549/A 0.44fF
C47155 OR2X1_LOC_801/B OR2X1_LOC_750/Y 0.00fF
C47156 OR2X1_LOC_163/a_36_216# OR2X1_LOC_163/Y 0.00fF
C47157 OR2X1_LOC_87/A AND2X1_LOC_607/a_8_24# 0.02fF
C47158 OR2X1_LOC_490/a_8_216# OR2X1_LOC_26/Y 0.03fF
C47159 AND2X1_LOC_721/Y OR2X1_LOC_74/A 0.03fF
C47160 AND2X1_LOC_716/Y AND2X1_LOC_364/Y 0.03fF
C47161 OR2X1_LOC_158/A AND2X1_LOC_287/Y 0.02fF
C47162 OR2X1_LOC_45/B OR2X1_LOC_239/Y 0.01fF
C47163 OR2X1_LOC_702/A OR2X1_LOC_139/A 0.02fF
C47164 OR2X1_LOC_49/A AND2X1_LOC_259/Y 0.48fF
C47165 OR2X1_LOC_643/A AND2X1_LOC_65/A 0.07fF
C47166 OR2X1_LOC_604/A OR2X1_LOC_427/a_8_216# 0.01fF
C47167 OR2X1_LOC_40/Y AND2X1_LOC_811/a_8_24# 0.01fF
C47168 OR2X1_LOC_121/Y OR2X1_LOC_217/a_8_216# 0.02fF
C47169 AND2X1_LOC_396/a_8_24# OR2X1_LOC_402/Y 0.02fF
C47170 OR2X1_LOC_207/B AND2X1_LOC_3/Y 0.03fF
C47171 OR2X1_LOC_456/A OR2X1_LOC_562/A 0.01fF
C47172 AND2X1_LOC_3/Y OR2X1_LOC_489/A 0.01fF
C47173 AND2X1_LOC_8/Y OR2X1_LOC_549/A 0.07fF
C47174 AND2X1_LOC_651/B OR2X1_LOC_18/a_8_216# 0.47fF
C47175 AND2X1_LOC_573/A AND2X1_LOC_657/Y 0.09fF
C47176 OR2X1_LOC_629/A OR2X1_LOC_161/B 0.13fF
C47177 OR2X1_LOC_151/A OR2X1_LOC_269/B 0.15fF
C47178 AND2X1_LOC_364/Y AND2X1_LOC_654/Y 0.04fF
C47179 AND2X1_LOC_640/Y AND2X1_LOC_219/A 0.17fF
C47180 OR2X1_LOC_47/Y AND2X1_LOC_608/a_8_24# 0.04fF
C47181 AND2X1_LOC_191/B AND2X1_LOC_573/A 0.07fF
C47182 OR2X1_LOC_418/a_8_216# OR2X1_LOC_16/A 0.09fF
C47183 OR2X1_LOC_426/B OR2X1_LOC_67/A 0.17fF
C47184 OR2X1_LOC_355/B OR2X1_LOC_356/A 0.81fF
C47185 OR2X1_LOC_124/a_36_216# OR2X1_LOC_375/A 0.00fF
C47186 OR2X1_LOC_256/Y OR2X1_LOC_92/Y 0.07fF
C47187 OR2X1_LOC_154/A OR2X1_LOC_676/Y 0.03fF
C47188 VDD AND2X1_LOC_303/A 0.06fF
C47189 OR2X1_LOC_453/a_8_216# OR2X1_LOC_466/A 0.01fF
C47190 OR2X1_LOC_375/A OR2X1_LOC_787/B 0.01fF
C47191 OR2X1_LOC_204/Y AND2X1_LOC_18/Y 0.03fF
C47192 OR2X1_LOC_502/A OR2X1_LOC_775/a_8_216# 0.05fF
C47193 OR2X1_LOC_510/A OR2X1_LOC_643/A 0.23fF
C47194 AND2X1_LOC_91/B OR2X1_LOC_846/A 0.01fF
C47195 AND2X1_LOC_578/A OR2X1_LOC_373/Y 0.03fF
C47196 OR2X1_LOC_91/Y OR2X1_LOC_51/Y 0.18fF
C47197 AND2X1_LOC_794/B OR2X1_LOC_485/A 0.19fF
C47198 OR2X1_LOC_375/A AND2X1_LOC_92/Y 0.09fF
C47199 AND2X1_LOC_475/a_8_24# AND2X1_LOC_475/Y 0.02fF
C47200 AND2X1_LOC_334/a_36_24# AND2X1_LOC_640/Y 0.01fF
C47201 AND2X1_LOC_12/Y OR2X1_LOC_678/a_8_216# 0.03fF
C47202 VDD OR2X1_LOC_845/a_8_216# 0.21fF
C47203 AND2X1_LOC_98/a_36_24# OR2X1_LOC_6/A 0.00fF
C47204 OR2X1_LOC_76/B OR2X1_LOC_464/A 0.01fF
C47205 INPUT_1 OR2X1_LOC_748/a_8_216# 0.01fF
C47206 VDD OR2X1_LOC_81/Y 0.12fF
C47207 OR2X1_LOC_139/A OR2X1_LOC_476/B 0.03fF
C47208 AND2X1_LOC_729/B AND2X1_LOC_774/A 0.03fF
C47209 OR2X1_LOC_524/Y AND2X1_LOC_676/a_36_24# 0.08fF
C47210 OR2X1_LOC_631/B OR2X1_LOC_66/A 0.07fF
C47211 D_INPUT_5 AND2X1_LOC_11/Y 0.65fF
C47212 OR2X1_LOC_516/A AND2X1_LOC_471/Y 0.03fF
C47213 OR2X1_LOC_6/B OR2X1_LOC_574/A 0.10fF
C47214 OR2X1_LOC_518/Y OR2X1_LOC_111/Y 0.05fF
C47215 AND2X1_LOC_3/Y OR2X1_LOC_772/A 0.54fF
C47216 OR2X1_LOC_744/A AND2X1_LOC_266/Y 0.01fF
C47217 OR2X1_LOC_283/Y AND2X1_LOC_286/a_8_24# 0.10fF
C47218 AND2X1_LOC_359/B OR2X1_LOC_56/A 0.03fF
C47219 OR2X1_LOC_416/Y AND2X1_LOC_219/A 0.00fF
C47220 VDD OR2X1_LOC_665/Y 0.32fF
C47221 VDD AND2X1_LOC_474/Y 0.18fF
C47222 OR2X1_LOC_426/B OR2X1_LOC_52/B 0.36fF
C47223 OR2X1_LOC_51/Y AND2X1_LOC_446/a_8_24# 0.01fF
C47224 AND2X1_LOC_711/Y AND2X1_LOC_347/B 0.01fF
C47225 OR2X1_LOC_731/a_8_216# OR2X1_LOC_738/B -0.00fF
C47226 AND2X1_LOC_40/Y OR2X1_LOC_624/A 0.01fF
C47227 OR2X1_LOC_688/a_8_216# OR2X1_LOC_66/A 0.02fF
C47228 OR2X1_LOC_287/B OR2X1_LOC_858/a_36_216# -0.00fF
C47229 AND2X1_LOC_787/a_8_24# OR2X1_LOC_48/B 0.04fF
C47230 OR2X1_LOC_268/a_8_216# AND2X1_LOC_786/Y 0.03fF
C47231 OR2X1_LOC_494/Y OR2X1_LOC_7/A 0.03fF
C47232 OR2X1_LOC_469/Y OR2X1_LOC_161/A 0.03fF
C47233 AND2X1_LOC_719/Y OR2X1_LOC_488/a_8_216# 0.22fF
C47234 OR2X1_LOC_151/A OR2X1_LOC_215/A 0.03fF
C47235 AND2X1_LOC_22/a_8_24# AND2X1_LOC_11/Y 0.01fF
C47236 OR2X1_LOC_101/a_8_216# OR2X1_LOC_656/B 0.01fF
C47237 AND2X1_LOC_363/Y OR2X1_LOC_7/A 0.04fF
C47238 VDD OR2X1_LOC_485/A 0.61fF
C47239 OR2X1_LOC_792/Y OR2X1_LOC_288/a_8_216# 0.01fF
C47240 OR2X1_LOC_814/A AND2X1_LOC_44/Y 0.03fF
C47241 OR2X1_LOC_696/A AND2X1_LOC_798/A 0.03fF
C47242 AND2X1_LOC_53/Y AND2X1_LOC_7/B 0.07fF
C47243 AND2X1_LOC_720/a_8_24# OR2X1_LOC_278/Y 0.01fF
C47244 AND2X1_LOC_555/Y D_INPUT_3 0.54fF
C47245 AND2X1_LOC_707/a_36_24# OR2X1_LOC_7/A 0.01fF
C47246 AND2X1_LOC_12/Y OR2X1_LOC_808/a_8_216# 0.01fF
C47247 AND2X1_LOC_474/A AND2X1_LOC_806/A 1.73fF
C47248 OR2X1_LOC_625/Y OR2X1_LOC_278/Y 0.01fF
C47249 OR2X1_LOC_238/Y OR2X1_LOC_59/Y 0.03fF
C47250 AND2X1_LOC_289/a_8_24# OR2X1_LOC_333/A 0.13fF
C47251 OR2X1_LOC_476/B OR2X1_LOC_654/a_36_216# 0.01fF
C47252 AND2X1_LOC_862/a_36_24# OR2X1_LOC_59/Y 0.00fF
C47253 OR2X1_LOC_323/A OR2X1_LOC_47/Y 0.02fF
C47254 OR2X1_LOC_715/B OR2X1_LOC_121/B 0.03fF
C47255 AND2X1_LOC_12/Y AND2X1_LOC_11/Y 0.01fF
C47256 VDD OR2X1_LOC_158/B 0.04fF
C47257 OR2X1_LOC_335/B AND2X1_LOC_603/a_36_24# 0.00fF
C47258 OR2X1_LOC_604/A OR2X1_LOC_488/Y 0.05fF
C47259 OR2X1_LOC_318/B OR2X1_LOC_593/B 0.03fF
C47260 OR2X1_LOC_222/A OR2X1_LOC_475/B 0.01fF
C47261 AND2X1_LOC_726/Y OR2X1_LOC_47/Y 0.01fF
C47262 OR2X1_LOC_686/B AND2X1_LOC_51/Y 0.01fF
C47263 OR2X1_LOC_632/a_8_216# AND2X1_LOC_3/Y 0.02fF
C47264 OR2X1_LOC_148/Y OR2X1_LOC_471/Y 0.13fF
C47265 OR2X1_LOC_650/Y OR2X1_LOC_654/a_36_216# 0.02fF
C47266 OR2X1_LOC_164/Y OR2X1_LOC_26/Y 0.03fF
C47267 OR2X1_LOC_811/A OR2X1_LOC_553/A 0.07fF
C47268 OR2X1_LOC_446/Y OR2X1_LOC_161/B 0.25fF
C47269 OR2X1_LOC_656/B OR2X1_LOC_340/Y 0.02fF
C47270 AND2X1_LOC_211/B AND2X1_LOC_335/a_8_24# 0.01fF
C47271 AND2X1_LOC_12/Y OR2X1_LOC_402/Y 0.02fF
C47272 AND2X1_LOC_728/Y OR2X1_LOC_679/B 0.00fF
C47273 OR2X1_LOC_532/B OR2X1_LOC_736/Y 8.28fF
C47274 OR2X1_LOC_19/B OR2X1_LOC_607/A 0.01fF
C47275 OR2X1_LOC_517/A OR2X1_LOC_106/A 0.58fF
C47276 AND2X1_LOC_253/a_36_24# OR2X1_LOC_269/B 0.01fF
C47277 OR2X1_LOC_653/B OR2X1_LOC_532/B 0.00fF
C47278 OR2X1_LOC_517/Y AND2X1_LOC_76/Y 0.01fF
C47279 OR2X1_LOC_223/A AND2X1_LOC_7/B 0.03fF
C47280 OR2X1_LOC_36/Y AND2X1_LOC_832/a_8_24# 0.01fF
C47281 OR2X1_LOC_604/A AND2X1_LOC_727/A 0.03fF
C47282 OR2X1_LOC_427/A AND2X1_LOC_466/a_36_24# 0.00fF
C47283 OR2X1_LOC_523/A OR2X1_LOC_560/A 0.10fF
C47284 AND2X1_LOC_779/a_8_24# OR2X1_LOC_44/Y 0.02fF
C47285 OR2X1_LOC_164/Y OR2X1_LOC_89/A 0.03fF
C47286 OR2X1_LOC_417/Y OR2X1_LOC_51/Y 0.06fF
C47287 OR2X1_LOC_788/a_8_216# OR2X1_LOC_269/B 0.05fF
C47288 AND2X1_LOC_81/B OR2X1_LOC_506/A 0.03fF
C47289 AND2X1_LOC_90/a_36_24# AND2X1_LOC_47/Y 0.00fF
C47290 AND2X1_LOC_852/Y AND2X1_LOC_852/B 0.05fF
C47291 OR2X1_LOC_599/A AND2X1_LOC_832/a_36_24# 0.00fF
C47292 OR2X1_LOC_756/B AND2X1_LOC_42/B 0.04fF
C47293 AND2X1_LOC_139/B OR2X1_LOC_39/A 0.07fF
C47294 OR2X1_LOC_177/Y OR2X1_LOC_95/Y 0.03fF
C47295 OR2X1_LOC_696/A OR2X1_LOC_761/a_8_216# 0.04fF
C47296 AND2X1_LOC_852/Y OR2X1_LOC_48/B 0.35fF
C47297 OR2X1_LOC_8/Y OR2X1_LOC_246/A 0.00fF
C47298 INPUT_1 INPUT_2 0.26fF
C47299 OR2X1_LOC_3/Y AND2X1_LOC_402/a_8_24# 0.01fF
C47300 AND2X1_LOC_776/Y OR2X1_LOC_406/A 0.00fF
C47301 OR2X1_LOC_329/B OR2X1_LOC_64/Y 0.61fF
C47302 OR2X1_LOC_315/a_8_216# OR2X1_LOC_368/A 0.01fF
C47303 OR2X1_LOC_473/A OR2X1_LOC_161/B 0.31fF
C47304 AND2X1_LOC_273/a_8_24# OR2X1_LOC_318/B 0.00fF
C47305 AND2X1_LOC_130/a_8_24# AND2X1_LOC_227/Y 0.01fF
C47306 VDD OR2X1_LOC_335/B 0.00fF
C47307 OR2X1_LOC_91/Y OR2X1_LOC_680/A 0.03fF
C47308 OR2X1_LOC_669/A AND2X1_LOC_848/Y 0.20fF
C47309 OR2X1_LOC_18/Y AND2X1_LOC_852/Y 0.02fF
C47310 AND2X1_LOC_316/a_8_24# OR2X1_LOC_201/Y 0.23fF
C47311 INPUT_5 OR2X1_LOC_44/a_8_216# 0.01fF
C47312 OR2X1_LOC_186/Y AND2X1_LOC_420/a_8_24# 0.00fF
C47313 AND2X1_LOC_560/B AND2X1_LOC_113/Y 0.01fF
C47314 OR2X1_LOC_377/A OR2X1_LOC_83/A 0.07fF
C47315 OR2X1_LOC_683/a_8_216# OR2X1_LOC_70/Y 0.02fF
C47316 OR2X1_LOC_124/A AND2X1_LOC_667/a_8_24# 0.14fF
C47317 OR2X1_LOC_643/A OR2X1_LOC_659/a_8_216# 0.03fF
C47318 OR2X1_LOC_9/a_8_216# D_INPUT_1 0.01fF
C47319 AND2X1_LOC_639/A OR2X1_LOC_12/a_8_216# 0.03fF
C47320 OR2X1_LOC_519/Y AND2X1_LOC_211/B 0.01fF
C47321 INPUT_0 AND2X1_LOC_48/A 0.09fF
C47322 OR2X1_LOC_604/A OR2X1_LOC_95/Y 1.07fF
C47323 OR2X1_LOC_685/B OR2X1_LOC_87/A 0.01fF
C47324 AND2X1_LOC_76/Y OR2X1_LOC_743/A 0.40fF
C47325 AND2X1_LOC_758/a_8_24# OR2X1_LOC_95/Y 0.11fF
C47326 OR2X1_LOC_22/A OR2X1_LOC_26/a_8_216# 0.06fF
C47327 OR2X1_LOC_40/Y AND2X1_LOC_440/a_36_24# 0.00fF
C47328 AND2X1_LOC_339/B OR2X1_LOC_289/a_8_216# 0.01fF
C47329 OR2X1_LOC_469/Y AND2X1_LOC_51/Y 0.12fF
C47330 AND2X1_LOC_70/Y OR2X1_LOC_544/A 0.01fF
C47331 AND2X1_LOC_838/Y AND2X1_LOC_838/a_36_24# 0.00fF
C47332 OR2X1_LOC_821/a_8_216# OR2X1_LOC_86/A 0.39fF
C47333 OR2X1_LOC_6/B OR2X1_LOC_826/Y 0.01fF
C47334 OR2X1_LOC_517/Y OR2X1_LOC_52/B 0.03fF
C47335 OR2X1_LOC_479/Y OR2X1_LOC_185/A 0.04fF
C47336 OR2X1_LOC_529/Y OR2X1_LOC_39/A 0.05fF
C47337 OR2X1_LOC_137/a_8_216# OR2X1_LOC_720/B 0.02fF
C47338 OR2X1_LOC_329/B OR2X1_LOC_417/A 0.14fF
C47339 AND2X1_LOC_342/a_36_24# OR2X1_LOC_85/A 0.00fF
C47340 AND2X1_LOC_695/a_36_24# AND2X1_LOC_3/Y 0.00fF
C47341 VDD OR2X1_LOC_587/a_8_216# 0.00fF
C47342 OR2X1_LOC_70/Y OR2X1_LOC_118/Y 0.02fF
C47343 OR2X1_LOC_426/A AND2X1_LOC_635/a_8_24# 0.01fF
C47344 OR2X1_LOC_862/a_8_216# OR2X1_LOC_561/B 0.01fF
C47345 OR2X1_LOC_111/Y OR2X1_LOC_91/A 0.04fF
C47346 OR2X1_LOC_51/Y D_INPUT_3 0.03fF
C47347 OR2X1_LOC_485/A AND2X1_LOC_447/a_36_24# -0.00fF
C47348 OR2X1_LOC_218/a_36_216# OR2X1_LOC_643/A 0.02fF
C47349 OR2X1_LOC_756/B OR2X1_LOC_286/B 0.01fF
C47350 OR2X1_LOC_193/A OR2X1_LOC_161/A 0.00fF
C47351 AND2X1_LOC_92/a_8_24# OR2X1_LOC_68/B 0.03fF
C47352 VDD OR2X1_LOC_609/Y 0.04fF
C47353 OR2X1_LOC_506/B OR2X1_LOC_78/A 0.05fF
C47354 OR2X1_LOC_657/a_8_216# AND2X1_LOC_42/B 0.01fF
C47355 OR2X1_LOC_160/B AND2X1_LOC_237/a_8_24# 0.01fF
C47356 OR2X1_LOC_808/B OR2X1_LOC_532/B 0.05fF
C47357 OR2X1_LOC_161/B OR2X1_LOC_228/Y 0.46fF
C47358 OR2X1_LOC_361/a_8_216# OR2X1_LOC_140/a_8_216# 0.47fF
C47359 AND2X1_LOC_76/Y OR2X1_LOC_246/A 0.03fF
C47360 AND2X1_LOC_197/Y OR2X1_LOC_31/Y 0.01fF
C47361 OR2X1_LOC_485/A OR2X1_LOC_491/Y 0.01fF
C47362 AND2X1_LOC_343/a_8_24# OR2X1_LOC_585/A 0.02fF
C47363 OR2X1_LOC_527/Y OR2X1_LOC_680/A 0.07fF
C47364 AND2X1_LOC_36/Y OR2X1_LOC_308/Y 0.09fF
C47365 OR2X1_LOC_170/a_8_216# OR2X1_LOC_788/B 0.06fF
C47366 OR2X1_LOC_51/Y OR2X1_LOC_289/a_36_216# 0.00fF
C47367 AND2X1_LOC_227/Y OR2X1_LOC_517/A 0.03fF
C47368 OR2X1_LOC_251/Y OR2X1_LOC_485/A 0.03fF
C47369 OR2X1_LOC_743/A OR2X1_LOC_52/B 0.08fF
C47370 OR2X1_LOC_3/Y AND2X1_LOC_101/B 0.08fF
C47371 AND2X1_LOC_308/a_8_24# AND2X1_LOC_655/A 0.23fF
C47372 OR2X1_LOC_403/B OR2X1_LOC_624/B 0.03fF
C47373 AND2X1_LOC_605/Y AND2X1_LOC_645/a_8_24# 0.11fF
C47374 OR2X1_LOC_158/A AND2X1_LOC_562/Y 0.31fF
C47375 OR2X1_LOC_68/B OR2X1_LOC_343/a_8_216# 0.04fF
C47376 OR2X1_LOC_51/Y AND2X1_LOC_483/Y 0.02fF
C47377 OR2X1_LOC_696/Y OR2X1_LOC_591/A 0.15fF
C47378 OR2X1_LOC_306/Y AND2X1_LOC_727/A 0.01fF
C47379 OR2X1_LOC_70/Y OR2X1_LOC_262/Y 1.04fF
C47380 OR2X1_LOC_668/a_36_216# OR2X1_LOC_532/B 0.00fF
C47381 AND2X1_LOC_61/Y AND2X1_LOC_215/A 0.07fF
C47382 OR2X1_LOC_240/B D_INPUT_0 0.05fF
C47383 OR2X1_LOC_748/A OR2X1_LOC_261/A 0.02fF
C47384 INPUT_4 AND2X1_LOC_635/a_8_24# 0.01fF
C47385 AND2X1_LOC_723/Y OR2X1_LOC_47/Y 0.07fF
C47386 OR2X1_LOC_185/Y OR2X1_LOC_206/A 0.03fF
C47387 OR2X1_LOC_680/A AND2X1_LOC_574/A 0.08fF
C47388 OR2X1_LOC_809/B OR2X1_LOC_801/B 0.03fF
C47389 D_INPUT_0 OR2X1_LOC_161/A 0.53fF
C47390 OR2X1_LOC_316/Y AND2X1_LOC_640/a_8_24# 0.01fF
C47391 AND2X1_LOC_554/Y OR2X1_LOC_71/Y 0.01fF
C47392 OR2X1_LOC_247/Y OR2X1_LOC_78/A 0.01fF
C47393 OR2X1_LOC_841/a_36_216# OR2X1_LOC_223/A 0.00fF
C47394 OR2X1_LOC_679/A AND2X1_LOC_624/A 0.03fF
C47395 OR2X1_LOC_862/A D_INPUT_1 0.08fF
C47396 OR2X1_LOC_318/Y OR2X1_LOC_223/A 0.03fF
C47397 AND2X1_LOC_95/Y OR2X1_LOC_651/A 0.11fF
C47398 OR2X1_LOC_364/A AND2X1_LOC_600/a_8_24# 0.01fF
C47399 OR2X1_LOC_276/B OR2X1_LOC_833/B 0.84fF
C47400 OR2X1_LOC_517/A OR2X1_LOC_813/Y 0.00fF
C47401 OR2X1_LOC_43/A OR2X1_LOC_77/a_8_216# 0.04fF
C47402 OR2X1_LOC_827/a_8_216# OR2X1_LOC_46/A 0.01fF
C47403 AND2X1_LOC_633/Y OR2X1_LOC_26/Y 0.02fF
C47404 OR2X1_LOC_246/A OR2X1_LOC_52/B 0.10fF
C47405 OR2X1_LOC_682/Y AND2X1_LOC_687/A 0.01fF
C47406 OR2X1_LOC_808/A OR2X1_LOC_374/Y 0.07fF
C47407 AND2X1_LOC_196/Y OR2X1_LOC_43/A 0.02fF
C47408 OR2X1_LOC_656/B AND2X1_LOC_88/Y 0.81fF
C47409 OR2X1_LOC_316/Y AND2X1_LOC_649/Y 0.00fF
C47410 OR2X1_LOC_26/Y D_INPUT_0 0.35fF
C47411 OR2X1_LOC_804/A OR2X1_LOC_785/B 0.05fF
C47412 AND2X1_LOC_639/B OR2X1_LOC_386/a_8_216# 0.49fF
C47413 OR2X1_LOC_764/a_8_216# OR2X1_LOC_387/A 0.18fF
C47414 OR2X1_LOC_691/a_36_216# OR2X1_LOC_771/B 0.02fF
C47415 OR2X1_LOC_574/A OR2X1_LOC_68/Y 0.09fF
C47416 OR2X1_LOC_628/Y OR2X1_LOC_74/A 0.22fF
C47417 OR2X1_LOC_481/A OR2X1_LOC_295/a_36_216# 0.00fF
C47418 D_INPUT_0 OR2X1_LOC_89/A 1.72fF
C47419 AND2X1_LOC_810/Y AND2X1_LOC_661/A 0.02fF
C47420 AND2X1_LOC_81/B OR2X1_LOC_227/Y 0.00fF
C47421 OR2X1_LOC_773/B D_INPUT_1 0.04fF
C47422 OR2X1_LOC_486/Y OR2X1_LOC_469/B 4.61fF
C47423 OR2X1_LOC_280/Y OR2X1_LOC_71/Y 0.02fF
C47424 OR2X1_LOC_409/B OR2X1_LOC_52/B 0.06fF
C47425 OR2X1_LOC_711/a_8_216# OR2X1_LOC_469/B 0.02fF
C47426 OR2X1_LOC_506/A OR2X1_LOC_66/Y 0.00fF
C47427 OR2X1_LOC_574/A AND2X1_LOC_47/Y 0.01fF
C47428 INPUT_1 AND2X1_LOC_847/a_8_24# 0.02fF
C47429 OR2X1_LOC_160/B OR2X1_LOC_777/B 0.07fF
C47430 AND2X1_LOC_499/a_8_24# OR2X1_LOC_142/Y 0.03fF
C47431 OR2X1_LOC_59/Y AND2X1_LOC_215/a_36_24# 0.00fF
C47432 OR2X1_LOC_448/A AND2X1_LOC_31/Y 0.00fF
C47433 OR2X1_LOC_40/a_8_216# OR2X1_LOC_70/A 0.06fF
C47434 OR2X1_LOC_553/A AND2X1_LOC_237/a_8_24# 0.07fF
C47435 OR2X1_LOC_541/a_8_216# OR2X1_LOC_241/B 0.02fF
C47436 OR2X1_LOC_485/A OR2X1_LOC_256/A 0.42fF
C47437 OR2X1_LOC_160/A OR2X1_LOC_493/Y 0.10fF
C47438 OR2X1_LOC_128/a_36_216# AND2X1_LOC_72/B 0.00fF
C47439 OR2X1_LOC_464/A OR2X1_LOC_578/B 0.03fF
C47440 OR2X1_LOC_158/a_36_216# OR2X1_LOC_163/Y 0.00fF
C47441 OR2X1_LOC_59/Y OR2X1_LOC_300/a_8_216# 0.01fF
C47442 OR2X1_LOC_61/Y OR2X1_LOC_228/Y 0.07fF
C47443 AND2X1_LOC_95/Y OR2X1_LOC_728/B 0.20fF
C47444 OR2X1_LOC_793/A AND2X1_LOC_39/Y 0.16fF
C47445 D_INPUT_0 AND2X1_LOC_51/Y 0.12fF
C47446 OR2X1_LOC_39/A OR2X1_LOC_598/A 0.06fF
C47447 OR2X1_LOC_161/B OR2X1_LOC_562/A 0.03fF
C47448 OR2X1_LOC_562/B OR2X1_LOC_562/A 0.14fF
C47449 AND2X1_LOC_364/Y OR2X1_LOC_13/B 0.09fF
C47450 OR2X1_LOC_214/a_8_216# OR2X1_LOC_214/B 0.06fF
C47451 OR2X1_LOC_649/a_8_216# OR2X1_LOC_655/A -0.00fF
C47452 OR2X1_LOC_185/A OR2X1_LOC_68/B 0.04fF
C47453 OR2X1_LOC_665/Y AND2X1_LOC_624/B 0.07fF
C47454 OR2X1_LOC_249/Y OR2X1_LOC_68/B 0.16fF
C47455 OR2X1_LOC_720/B OR2X1_LOC_814/A 0.03fF
C47456 AND2X1_LOC_601/a_8_24# AND2X1_LOC_31/Y 0.01fF
C47457 OR2X1_LOC_22/Y OR2X1_LOC_71/Y 2.30fF
C47458 OR2X1_LOC_754/A OR2X1_LOC_47/Y 0.06fF
C47459 OR2X1_LOC_696/A OR2X1_LOC_125/a_8_216# 0.00fF
C47460 AND2X1_LOC_544/Y AND2X1_LOC_477/Y 0.07fF
C47461 AND2X1_LOC_369/a_36_24# OR2X1_LOC_318/B 0.00fF
C47462 AND2X1_LOC_3/Y OR2X1_LOC_194/a_8_216# 0.01fF
C47463 OR2X1_LOC_744/A OR2X1_LOC_183/Y 0.02fF
C47464 OR2X1_LOC_485/A OR2X1_LOC_67/Y 0.01fF
C47465 AND2X1_LOC_672/B AND2X1_LOC_47/Y 0.00fF
C47466 OR2X1_LOC_7/A AND2X1_LOC_228/a_8_24# 0.02fF
C47467 OR2X1_LOC_691/A OR2X1_LOC_691/B 0.61fF
C47468 OR2X1_LOC_317/A OR2X1_LOC_317/B 0.04fF
C47469 OR2X1_LOC_168/B OR2X1_LOC_776/A 0.08fF
C47470 OR2X1_LOC_574/A OR2X1_LOC_598/A 0.15fF
C47471 OR2X1_LOC_160/B OR2X1_LOC_831/B 0.01fF
C47472 OR2X1_LOC_86/Y OR2X1_LOC_88/Y 0.08fF
C47473 OR2X1_LOC_51/Y AND2X1_LOC_780/a_8_24# 0.01fF
C47474 OR2X1_LOC_40/Y AND2X1_LOC_241/a_36_24# 0.00fF
C47475 OR2X1_LOC_188/a_8_216# OR2X1_LOC_160/B 0.01fF
C47476 OR2X1_LOC_49/A OR2X1_LOC_671/Y 0.81fF
C47477 OR2X1_LOC_51/Y OR2X1_LOC_171/Y 0.53fF
C47478 OR2X1_LOC_216/A AND2X1_LOC_239/a_8_24# 0.03fF
C47479 AND2X1_LOC_457/a_8_24# AND2X1_LOC_476/Y 0.02fF
C47480 AND2X1_LOC_866/A INPUT_1 0.07fF
C47481 OR2X1_LOC_156/Y OR2X1_LOC_160/B 0.15fF
C47482 OR2X1_LOC_92/a_8_216# D_INPUT_0 0.03fF
C47483 AND2X1_LOC_803/B AND2X1_LOC_220/B 0.03fF
C47484 AND2X1_LOC_706/Y AND2X1_LOC_713/a_8_24# 0.01fF
C47485 OR2X1_LOC_379/Y OR2X1_LOC_769/a_8_216# 0.01fF
C47486 AND2X1_LOC_721/Y AND2X1_LOC_860/A 0.02fF
C47487 VDD OR2X1_LOC_267/Y -0.00fF
C47488 AND2X1_LOC_802/B VDD 0.01fF
C47489 OR2X1_LOC_158/A OR2X1_LOC_381/a_8_216# 0.02fF
C47490 OR2X1_LOC_78/A AND2X1_LOC_258/a_8_24# 0.03fF
C47491 AND2X1_LOC_588/B AND2X1_LOC_588/a_8_24# 0.00fF
C47492 OR2X1_LOC_160/A OR2X1_LOC_532/a_8_216# 0.05fF
C47493 OR2X1_LOC_158/B OR2X1_LOC_163/Y 0.22fF
C47494 OR2X1_LOC_820/A OR2X1_LOC_748/Y 0.05fF
C47495 OR2X1_LOC_421/A AND2X1_LOC_706/a_8_24# 0.01fF
C47496 VDD OR2X1_LOC_633/A 0.51fF
C47497 OR2X1_LOC_244/Y AND2X1_LOC_44/Y 0.03fF
C47498 OR2X1_LOC_196/B AND2X1_LOC_48/Y 0.04fF
C47499 AND2X1_LOC_59/Y OR2X1_LOC_771/B 0.05fF
C47500 OR2X1_LOC_158/A AND2X1_LOC_448/a_8_24# 0.01fF
C47501 VDD OR2X1_LOC_725/A -0.00fF
C47502 OR2X1_LOC_421/A OR2X1_LOC_589/A 0.04fF
C47503 AND2X1_LOC_12/Y OR2X1_LOC_593/B 0.57fF
C47504 AND2X1_LOC_64/Y OR2X1_LOC_798/Y 0.01fF
C47505 AND2X1_LOC_434/Y OR2X1_LOC_428/A 0.14fF
C47506 OR2X1_LOC_78/A OR2X1_LOC_708/a_8_216# 0.01fF
C47507 AND2X1_LOC_357/A AND2X1_LOC_566/B 0.02fF
C47508 OR2X1_LOC_309/a_8_216# OR2X1_LOC_309/Y 0.01fF
C47509 OR2X1_LOC_87/A OR2X1_LOC_544/B 0.08fF
C47510 AND2X1_LOC_633/Y AND2X1_LOC_202/a_8_24# 0.17fF
C47511 AND2X1_LOC_748/a_36_24# AND2X1_LOC_36/Y 0.00fF
C47512 AND2X1_LOC_40/Y OR2X1_LOC_556/a_8_216# 0.19fF
C47513 AND2X1_LOC_198/a_8_24# OR2X1_LOC_56/Y 0.01fF
C47514 OR2X1_LOC_154/A AND2X1_LOC_591/a_8_24# 0.02fF
C47515 OR2X1_LOC_501/B AND2X1_LOC_44/Y 0.18fF
C47516 AND2X1_LOC_320/a_36_24# AND2X1_LOC_44/Y 0.00fF
C47517 OR2X1_LOC_124/a_36_216# OR2X1_LOC_549/A 0.00fF
C47518 OR2X1_LOC_426/B OR2X1_LOC_13/a_8_216# 0.08fF
C47519 OR2X1_LOC_160/A OR2X1_LOC_130/a_8_216# 0.04fF
C47520 OR2X1_LOC_175/Y OR2X1_LOC_840/A 0.10fF
C47521 AND2X1_LOC_59/Y OR2X1_LOC_776/A 0.07fF
C47522 OR2X1_LOC_479/Y OR2X1_LOC_705/a_8_216# 0.06fF
C47523 OR2X1_LOC_502/A AND2X1_LOC_7/B 4.98fF
C47524 AND2X1_LOC_530/a_8_24# INPUT_0 0.03fF
C47525 AND2X1_LOC_92/Y OR2X1_LOC_549/A 0.05fF
C47526 OR2X1_LOC_303/A OR2X1_LOC_186/Y 0.04fF
C47527 OR2X1_LOC_841/B OR2X1_LOC_593/B 0.01fF
C47528 OR2X1_LOC_843/a_8_216# OR2X1_LOC_580/A 0.03fF
C47529 AND2X1_LOC_17/a_8_24# D_INPUT_6 0.01fF
C47530 OR2X1_LOC_58/Y OR2X1_LOC_60/Y 0.21fF
C47531 AND2X1_LOC_803/B AND2X1_LOC_209/a_8_24# 0.01fF
C47532 OR2X1_LOC_441/Y AND2X1_LOC_727/B 0.03fF
C47533 OR2X1_LOC_666/A AND2X1_LOC_243/Y 0.28fF
C47534 AND2X1_LOC_837/a_8_24# AND2X1_LOC_838/B 0.00fF
C47535 OR2X1_LOC_506/a_8_216# AND2X1_LOC_12/Y 0.03fF
C47536 AND2X1_LOC_70/Y OR2X1_LOC_140/A 0.01fF
C47537 AND2X1_LOC_773/Y AND2X1_LOC_716/Y 0.10fF
C47538 AND2X1_LOC_95/Y OR2X1_LOC_338/A 0.01fF
C47539 OR2X1_LOC_147/B AND2X1_LOC_44/Y 0.09fF
C47540 AND2X1_LOC_516/a_8_24# AND2X1_LOC_36/Y 0.01fF
C47541 OR2X1_LOC_51/Y AND2X1_LOC_254/a_36_24# 0.01fF
C47542 OR2X1_LOC_696/A AND2X1_LOC_852/a_8_24# 0.01fF
C47543 OR2X1_LOC_585/A OR2X1_LOC_395/a_8_216# 0.05fF
C47544 OR2X1_LOC_485/Y OR2X1_LOC_484/a_8_216# 0.10fF
C47545 OR2X1_LOC_178/a_8_216# OR2X1_LOC_56/A 0.03fF
C47546 OR2X1_LOC_840/A OR2X1_LOC_713/A 0.02fF
C47547 OR2X1_LOC_178/Y OR2X1_LOC_600/A 0.03fF
C47548 OR2X1_LOC_18/Y AND2X1_LOC_284/a_8_24# 0.01fF
C47549 AND2X1_LOC_787/A OR2X1_LOC_48/B 0.31fF
C47550 OR2X1_LOC_78/A AND2X1_LOC_18/Y 0.18fF
C47551 OR2X1_LOC_609/Y OR2X1_LOC_67/Y 0.12fF
C47552 AND2X1_LOC_773/Y AND2X1_LOC_654/Y 0.10fF
C47553 AND2X1_LOC_330/a_8_24# OR2X1_LOC_51/Y 0.10fF
C47554 AND2X1_LOC_566/B AND2X1_LOC_303/a_36_24# 0.00fF
C47555 AND2X1_LOC_649/B AND2X1_LOC_786/Y 0.01fF
C47556 AND2X1_LOC_230/a_8_24# AND2X1_LOC_7/B 0.09fF
C47557 OR2X1_LOC_841/A OR2X1_LOC_648/A 0.03fF
C47558 OR2X1_LOC_92/Y OR2X1_LOC_829/A 0.10fF
C47559 OR2X1_LOC_585/A OR2X1_LOC_387/A 0.06fF
C47560 OR2X1_LOC_188/Y OR2X1_LOC_541/a_8_216# 0.01fF
C47561 OR2X1_LOC_198/a_36_216# OR2X1_LOC_269/B 0.00fF
C47562 OR2X1_LOC_804/B OR2X1_LOC_593/B 0.20fF
C47563 OR2X1_LOC_363/B OR2X1_LOC_363/A 0.18fF
C47564 AND2X1_LOC_514/a_8_24# OR2X1_LOC_426/B 0.03fF
C47565 OR2X1_LOC_109/Y OR2X1_LOC_323/a_8_216# 0.03fF
C47566 OR2X1_LOC_693/a_8_216# OR2X1_LOC_48/B 0.02fF
C47567 AND2X1_LOC_716/Y AND2X1_LOC_180/a_36_24# 0.01fF
C47568 OR2X1_LOC_611/Y OR2X1_LOC_71/A 0.03fF
C47569 OR2X1_LOC_186/Y AND2X1_LOC_95/Y 0.28fF
C47570 OR2X1_LOC_379/a_36_216# OR2X1_LOC_691/Y 0.00fF
C47571 OR2X1_LOC_352/A VDD -0.00fF
C47572 OR2X1_LOC_489/B OR2X1_LOC_489/A 1.23fF
C47573 OR2X1_LOC_693/a_8_216# OR2X1_LOC_18/Y 0.04fF
C47574 AND2X1_LOC_326/a_36_24# OR2X1_LOC_437/A 0.01fF
C47575 OR2X1_LOC_256/Y OR2X1_LOC_600/A 0.03fF
C47576 AND2X1_LOC_669/a_8_24# AND2X1_LOC_44/Y 0.01fF
C47577 OR2X1_LOC_79/Y OR2X1_LOC_265/Y 0.03fF
C47578 AND2X1_LOC_552/a_8_24# OR2X1_LOC_26/Y 0.01fF
C47579 OR2X1_LOC_772/B OR2X1_LOC_772/A 0.00fF
C47580 OR2X1_LOC_715/B OR2X1_LOC_856/B 0.10fF
C47581 AND2X1_LOC_40/Y AND2X1_LOC_265/a_36_24# 0.01fF
C47582 OR2X1_LOC_680/a_8_216# OR2X1_LOC_26/Y 0.01fF
C47583 OR2X1_LOC_43/A OR2X1_LOC_321/a_8_216# 0.05fF
C47584 AND2X1_LOC_566/B OR2X1_LOC_48/B 0.12fF
C47585 OR2X1_LOC_160/B OR2X1_LOC_575/A 0.03fF
C47586 AND2X1_LOC_714/B OR2X1_LOC_433/Y 0.13fF
C47587 OR2X1_LOC_756/B OR2X1_LOC_363/A 0.04fF
C47588 AND2X1_LOC_40/Y OR2X1_LOC_190/Y 0.88fF
C47589 AND2X1_LOC_550/A AND2X1_LOC_477/Y 0.07fF
C47590 OR2X1_LOC_6/A AND2X1_LOC_219/A 0.01fF
C47591 OR2X1_LOC_831/A OR2X1_LOC_161/A 0.02fF
C47592 OR2X1_LOC_151/A OR2X1_LOC_347/B 0.01fF
C47593 AND2X1_LOC_42/B OR2X1_LOC_140/B 0.03fF
C47594 OR2X1_LOC_19/B AND2X1_LOC_36/Y 0.19fF
C47595 OR2X1_LOC_446/Y OR2X1_LOC_707/a_8_216# 0.01fF
C47596 OR2X1_LOC_49/A OR2X1_LOC_42/a_8_216# 0.01fF
C47597 OR2X1_LOC_151/A OR2X1_LOC_539/Y 0.03fF
C47598 OR2X1_LOC_354/A AND2X1_LOC_92/Y 0.07fF
C47599 OR2X1_LOC_154/A AND2X1_LOC_83/a_8_24# 0.04fF
C47600 AND2X1_LOC_185/a_36_24# OR2X1_LOC_56/A 0.01fF
C47601 AND2X1_LOC_350/B OR2X1_LOC_26/Y 0.03fF
C47602 AND2X1_LOC_797/A AND2X1_LOC_209/Y 0.09fF
C47603 AND2X1_LOC_554/a_8_24# AND2X1_LOC_489/Y 0.01fF
C47604 OR2X1_LOC_6/B OR2X1_LOC_377/A 0.05fF
C47605 OR2X1_LOC_790/A OR2X1_LOC_375/A 0.26fF
C47606 OR2X1_LOC_693/Y OR2X1_LOC_36/Y 0.01fF
C47607 OR2X1_LOC_634/A OR2X1_LOC_334/B 0.08fF
C47608 AND2X1_LOC_595/a_8_24# OR2X1_LOC_249/Y 0.23fF
C47609 OR2X1_LOC_604/A OR2X1_LOC_257/a_36_216# 0.01fF
C47610 AND2X1_LOC_191/Y AND2X1_LOC_213/a_36_24# 0.01fF
C47611 OR2X1_LOC_208/A AND2X1_LOC_51/Y 0.02fF
C47612 OR2X1_LOC_143/a_8_216# OR2X1_LOC_54/Y 0.01fF
C47613 OR2X1_LOC_653/Y AND2X1_LOC_70/Y 0.17fF
C47614 AND2X1_LOC_553/A OR2X1_LOC_744/A 0.02fF
C47615 OR2X1_LOC_161/A OR2X1_LOC_356/a_8_216# 0.01fF
C47616 OR2X1_LOC_691/Y OR2X1_LOC_789/a_8_216# 0.01fF
C47617 OR2X1_LOC_493/B OR2X1_LOC_506/A 0.04fF
C47618 OR2X1_LOC_612/B OR2X1_LOC_16/A 0.03fF
C47619 AND2X1_LOC_70/Y OR2X1_LOC_833/B 0.07fF
C47620 OR2X1_LOC_7/A AND2X1_LOC_802/Y 0.07fF
C47621 OR2X1_LOC_453/A OR2X1_LOC_161/B 0.02fF
C47622 AND2X1_LOC_387/B AND2X1_LOC_44/Y 2.30fF
C47623 OR2X1_LOC_599/A AND2X1_LOC_729/a_36_24# 0.00fF
C47624 OR2X1_LOC_117/a_36_216# OR2X1_LOC_490/Y 0.00fF
C47625 OR2X1_LOC_532/B OR2X1_LOC_703/Y 0.02fF
C47626 OR2X1_LOC_6/B OR2X1_LOC_85/A 0.19fF
C47627 OR2X1_LOC_6/B OR2X1_LOC_203/Y 0.01fF
C47628 OR2X1_LOC_131/A OR2X1_LOC_26/Y 0.03fF
C47629 AND2X1_LOC_474/A OR2X1_LOC_625/a_8_216# 0.47fF
C47630 OR2X1_LOC_31/Y OR2X1_LOC_386/a_8_216# 0.01fF
C47631 OR2X1_LOC_319/B OR2X1_LOC_502/A 0.83fF
C47632 OR2X1_LOC_702/A OR2X1_LOC_138/A 0.27fF
C47633 AND2X1_LOC_56/B AND2X1_LOC_411/a_8_24# 0.02fF
C47634 VDD OR2X1_LOC_520/Y 0.03fF
C47635 AND2X1_LOC_130/a_36_24# AND2X1_LOC_361/A 0.00fF
C47636 OR2X1_LOC_502/A AND2X1_LOC_402/a_8_24# 0.01fF
C47637 OR2X1_LOC_769/B OR2X1_LOC_379/Y 0.00fF
C47638 OR2X1_LOC_31/Y OR2X1_LOC_183/Y 0.01fF
C47639 OR2X1_LOC_216/A OR2X1_LOC_475/B 0.01fF
C47640 AND2X1_LOC_721/A OR2X1_LOC_437/A 0.24fF
C47641 AND2X1_LOC_663/B GATE_579 0.01fF
C47642 OR2X1_LOC_185/Y OR2X1_LOC_776/Y 0.07fF
C47643 OR2X1_LOC_9/Y OR2X1_LOC_585/A 0.01fF
C47644 OR2X1_LOC_421/A OR2X1_LOC_43/A 0.03fF
C47645 AND2X1_LOC_330/a_8_24# OR2X1_LOC_680/A 0.02fF
C47646 OR2X1_LOC_585/A AND2X1_LOC_193/Y 0.03fF
C47647 OR2X1_LOC_697/Y OR2X1_LOC_427/A 0.00fF
C47648 OR2X1_LOC_500/A OR2X1_LOC_78/A 0.01fF
C47649 OR2X1_LOC_47/Y OR2X1_LOC_142/Y 0.03fF
C47650 OR2X1_LOC_318/Y OR2X1_LOC_502/A 0.15fF
C47651 AND2X1_LOC_549/a_8_24# AND2X1_LOC_807/Y 0.11fF
C47652 OR2X1_LOC_131/A OR2X1_LOC_89/A 0.69fF
C47653 OR2X1_LOC_250/a_8_216# OR2X1_LOC_517/A 0.01fF
C47654 OR2X1_LOC_744/A OR2X1_LOC_511/Y 0.05fF
C47655 AND2X1_LOC_48/A AND2X1_LOC_7/B 0.28fF
C47656 OR2X1_LOC_155/A AND2X1_LOC_18/Y 0.15fF
C47657 AND2X1_LOC_506/a_8_24# AND2X1_LOC_807/Y 0.28fF
C47658 D_GATE_662 OR2X1_LOC_846/B 0.43fF
C47659 OR2X1_LOC_51/Y AND2X1_LOC_806/A 0.02fF
C47660 OR2X1_LOC_176/Y AND2X1_LOC_727/A 0.02fF
C47661 AND2X1_LOC_193/a_8_24# INPUT_0 0.01fF
C47662 AND2X1_LOC_568/B OR2X1_LOC_312/Y 0.07fF
C47663 AND2X1_LOC_535/Y AND2X1_LOC_337/B 0.02fF
C47664 OR2X1_LOC_151/A AND2X1_LOC_176/a_8_24# 0.01fF
C47665 OR2X1_LOC_228/Y AND2X1_LOC_406/a_8_24# 0.01fF
C47666 VDD OR2X1_LOC_420/a_8_216# 0.00fF
C47667 OR2X1_LOC_791/A OR2X1_LOC_161/A 0.09fF
C47668 AND2X1_LOC_48/a_36_24# OR2X1_LOC_161/A 0.01fF
C47669 OR2X1_LOC_287/A OR2X1_LOC_269/B 0.42fF
C47670 OR2X1_LOC_22/Y OR2X1_LOC_585/a_8_216# 0.01fF
C47671 AND2X1_LOC_40/Y OR2X1_LOC_161/A 0.11fF
C47672 VDD OR2X1_LOC_646/a_8_216# 0.21fF
C47673 OR2X1_LOC_364/A OR2X1_LOC_756/B 0.01fF
C47674 OR2X1_LOC_185/Y OR2X1_LOC_756/B 1.09fF
C47675 OR2X1_LOC_502/A OR2X1_LOC_805/A 0.07fF
C47676 AND2X1_LOC_508/B OR2X1_LOC_74/A 0.03fF
C47677 OR2X1_LOC_389/B OR2X1_LOC_78/B 0.05fF
C47678 OR2X1_LOC_136/Y AND2X1_LOC_831/Y 0.03fF
C47679 OR2X1_LOC_97/A OR2X1_LOC_655/B 0.01fF
C47680 OR2X1_LOC_600/A OR2X1_LOC_258/Y 0.01fF
C47681 OR2X1_LOC_499/B AND2X1_LOC_56/B 0.03fF
C47682 OR2X1_LOC_26/Y AND2X1_LOC_471/Y 0.03fF
C47683 AND2X1_LOC_52/a_36_24# AND2X1_LOC_43/B 0.00fF
C47684 OR2X1_LOC_235/B OR2X1_LOC_753/A 0.17fF
C47685 OR2X1_LOC_598/Y AND2X1_LOC_51/Y 0.02fF
C47686 OR2X1_LOC_3/Y AND2X1_LOC_454/a_8_24# 0.00fF
C47687 AND2X1_LOC_727/Y AND2X1_LOC_812/a_8_24# 0.20fF
C47688 AND2X1_LOC_12/Y AND2X1_LOC_492/a_8_24# 0.06fF
C47689 OR2X1_LOC_130/A OR2X1_LOC_785/B 0.01fF
C47690 OR2X1_LOC_49/A OR2X1_LOC_532/B 1.08fF
C47691 AND2X1_LOC_863/a_8_24# AND2X1_LOC_354/B 0.04fF
C47692 AND2X1_LOC_53/a_36_24# AND2X1_LOC_43/B 0.00fF
C47693 OR2X1_LOC_87/A AND2X1_LOC_424/a_8_24# 0.04fF
C47694 INPUT_0 AND2X1_LOC_3/Y 0.23fF
C47695 AND2X1_LOC_544/Y GATE_811 0.05fF
C47696 OR2X1_LOC_89/A AND2X1_LOC_471/Y 0.91fF
C47697 AND2X1_LOC_22/Y OR2X1_LOC_651/A 0.07fF
C47698 OR2X1_LOC_298/a_8_216# OR2X1_LOC_52/B 0.03fF
C47699 AND2X1_LOC_840/a_8_24# AND2X1_LOC_840/B 0.05fF
C47700 OR2X1_LOC_792/Y OR2X1_LOC_285/A 0.01fF
C47701 OR2X1_LOC_537/A OR2X1_LOC_161/A 0.00fF
C47702 AND2X1_LOC_392/a_8_24# AND2X1_LOC_554/B 0.17fF
C47703 OR2X1_LOC_367/B OR2X1_LOC_366/Y 0.23fF
C47704 OR2X1_LOC_403/B OR2X1_LOC_400/a_8_216# 0.01fF
C47705 AND2X1_LOC_59/Y OR2X1_LOC_402/Y 0.02fF
C47706 OR2X1_LOC_108/a_8_216# OR2X1_LOC_22/Y 0.05fF
C47707 OR2X1_LOC_185/A OR2X1_LOC_219/a_8_216# 0.01fF
C47708 OR2X1_LOC_235/B AND2X1_LOC_243/a_8_24# 0.00fF
C47709 AND2X1_LOC_705/Y OR2X1_LOC_31/Y 0.20fF
C47710 AND2X1_LOC_332/a_8_24# AND2X1_LOC_831/Y 0.04fF
C47711 AND2X1_LOC_851/B OR2X1_LOC_428/A 0.04fF
C47712 OR2X1_LOC_805/A AND2X1_LOC_230/a_8_24# 0.03fF
C47713 AND2X1_LOC_631/Y AND2X1_LOC_663/A 0.41fF
C47714 AND2X1_LOC_735/Y AND2X1_LOC_711/Y 0.03fF
C47715 OR2X1_LOC_619/Y AND2X1_LOC_470/A 0.01fF
C47716 VDD OR2X1_LOC_34/B -0.00fF
C47717 OR2X1_LOC_95/Y AND2X1_LOC_212/Y 0.07fF
C47718 OR2X1_LOC_532/B OR2X1_LOC_596/A 0.03fF
C47719 AND2X1_LOC_707/Y AND2X1_LOC_687/a_8_24# 0.01fF
C47720 AND2X1_LOC_180/a_8_24# OR2X1_LOC_417/A 0.04fF
C47721 OR2X1_LOC_76/B OR2X1_LOC_76/Y 0.06fF
C47722 OR2X1_LOC_147/B OR2X1_LOC_465/B 0.14fF
C47723 OR2X1_LOC_633/Y AND2X1_LOC_49/a_8_24# 0.23fF
C47724 AND2X1_LOC_482/a_8_24# OR2X1_LOC_269/B 0.01fF
C47725 OR2X1_LOC_40/Y INPUT_1 0.06fF
C47726 VDD AND2X1_LOC_107/a_8_24# 0.00fF
C47727 OR2X1_LOC_36/Y AND2X1_LOC_621/Y 0.05fF
C47728 AND2X1_LOC_564/B AND2X1_LOC_795/Y -0.00fF
C47729 OR2X1_LOC_426/B OR2X1_LOC_22/Y 0.37fF
C47730 AND2X1_LOC_486/Y OR2X1_LOC_485/A 0.06fF
C47731 OR2X1_LOC_160/A OR2X1_LOC_835/a_8_216# 0.07fF
C47732 OR2X1_LOC_628/a_8_216# OR2X1_LOC_7/A 0.01fF
C47733 AND2X1_LOC_61/Y AND2X1_LOC_634/Y 0.04fF
C47734 OR2X1_LOC_405/A OR2X1_LOC_778/Y 0.14fF
C47735 AND2X1_LOC_719/Y AND2X1_LOC_859/B 0.05fF
C47736 AND2X1_LOC_59/Y OR2X1_LOC_642/a_8_216# 0.01fF
C47737 OR2X1_LOC_599/A AND2X1_LOC_624/A 0.03fF
C47738 AND2X1_LOC_367/A AND2X1_LOC_523/Y 0.46fF
C47739 AND2X1_LOC_840/A OR2X1_LOC_89/A 0.07fF
C47740 OR2X1_LOC_90/a_8_216# OR2X1_LOC_54/Y 0.07fF
C47741 AND2X1_LOC_303/A AND2X1_LOC_716/a_8_24# 0.05fF
C47742 OR2X1_LOC_511/Y AND2X1_LOC_840/B 0.01fF
C47743 AND2X1_LOC_803/B OR2X1_LOC_679/A 0.00fF
C47744 OR2X1_LOC_26/Y OR2X1_LOC_237/a_8_216# 0.02fF
C47745 OR2X1_LOC_696/A AND2X1_LOC_657/A 0.07fF
C47746 OR2X1_LOC_653/Y OR2X1_LOC_653/a_8_216# 0.02fF
C47747 OR2X1_LOC_329/B OR2X1_LOC_268/a_36_216# 0.01fF
C47748 OR2X1_LOC_807/B OR2X1_LOC_807/a_8_216# 0.01fF
C47749 OR2X1_LOC_267/Y OR2X1_LOC_140/a_8_216# 0.01fF
C47750 OR2X1_LOC_574/A OR2X1_LOC_506/A 0.03fF
C47751 OR2X1_LOC_680/Y OR2X1_LOC_427/A 0.03fF
C47752 OR2X1_LOC_656/B AND2X1_LOC_88/a_8_24# 0.01fF
C47753 OR2X1_LOC_493/a_36_216# OR2X1_LOC_532/B 0.00fF
C47754 OR2X1_LOC_622/a_8_216# OR2X1_LOC_847/A 0.01fF
C47755 AND2X1_LOC_40/Y AND2X1_LOC_51/Y 0.18fF
C47756 AND2X1_LOC_99/Y OR2X1_LOC_64/Y 0.03fF
C47757 AND2X1_LOC_118/a_8_24# OR2X1_LOC_375/A 0.01fF
C47758 AND2X1_LOC_193/a_8_24# OR2X1_LOC_690/A 0.02fF
C47759 AND2X1_LOC_627/a_8_24# OR2X1_LOC_598/A 0.11fF
C47760 AND2X1_LOC_562/a_8_24# AND2X1_LOC_562/Y 0.01fF
C47761 OR2X1_LOC_489/B AND2X1_LOC_3/Y 0.00fF
C47762 AND2X1_LOC_739/a_8_24# AND2X1_LOC_740/B 0.01fF
C47763 AND2X1_LOC_379/a_36_24# OR2X1_LOC_26/Y 0.01fF
C47764 OR2X1_LOC_720/A OR2X1_LOC_720/a_8_216# 0.47fF
C47765 AND2X1_LOC_749/a_8_24# OR2X1_LOC_750/A 0.01fF
C47766 OR2X1_LOC_625/Y OR2X1_LOC_754/A 0.19fF
C47767 AND2X1_LOC_578/A OR2X1_LOC_109/Y 0.07fF
C47768 OR2X1_LOC_26/Y AND2X1_LOC_668/a_36_24# 0.00fF
C47769 OR2X1_LOC_673/Y OR2X1_LOC_849/A 0.01fF
C47770 AND2X1_LOC_335/Y AND2X1_LOC_318/Y 0.51fF
C47771 OR2X1_LOC_696/Y OR2X1_LOC_427/A 0.03fF
C47772 OR2X1_LOC_132/Y AND2X1_LOC_656/Y 0.01fF
C47773 OR2X1_LOC_3/Y AND2X1_LOC_449/Y 0.01fF
C47774 OR2X1_LOC_596/Y OR2X1_LOC_155/A 0.04fF
C47775 AND2X1_LOC_836/a_8_24# AND2X1_LOC_839/B 0.00fF
C47776 AND2X1_LOC_31/Y OR2X1_LOC_375/a_8_216# 0.01fF
C47777 AND2X1_LOC_549/a_8_24# OR2X1_LOC_95/Y 0.15fF
C47778 AND2X1_LOC_852/Y OR2X1_LOC_585/A 0.03fF
C47779 AND2X1_LOC_512/a_8_24# OR2X1_LOC_43/A 0.01fF
C47780 OR2X1_LOC_503/Y OR2X1_LOC_59/Y 0.01fF
C47781 OR2X1_LOC_756/B OR2X1_LOC_443/a_36_216# 0.00fF
C47782 OR2X1_LOC_656/B OR2X1_LOC_121/B 0.01fF
C47783 OR2X1_LOC_83/Y OR2X1_LOC_585/A 0.05fF
C47784 OR2X1_LOC_363/a_8_216# OR2X1_LOC_580/A 0.04fF
C47785 INPUT_0 AND2X1_LOC_476/A 0.09fF
C47786 AND2X1_LOC_62/a_8_24# OR2X1_LOC_46/A 0.02fF
C47787 OR2X1_LOC_223/A OR2X1_LOC_742/a_8_216# 0.01fF
C47788 OR2X1_LOC_485/A OR2X1_LOC_248/Y 0.41fF
C47789 OR2X1_LOC_469/B OR2X1_LOC_308/Y 0.20fF
C47790 OR2X1_LOC_744/A AND2X1_LOC_648/B 0.00fF
C47791 OR2X1_LOC_422/Y AND2X1_LOC_477/A 0.13fF
C47792 OR2X1_LOC_564/B OR2X1_LOC_564/A 0.13fF
C47793 OR2X1_LOC_88/Y AND2X1_LOC_249/a_8_24# 0.01fF
C47794 AND2X1_LOC_355/a_8_24# OR2X1_LOC_312/Y 0.01fF
C47795 AND2X1_LOC_727/a_8_24# OR2X1_LOC_152/A 0.21fF
C47796 OR2X1_LOC_490/Y OR2X1_LOC_117/Y 0.00fF
C47797 AND2X1_LOC_863/a_8_24# AND2X1_LOC_863/Y 0.01fF
C47798 OR2X1_LOC_600/A OR2X1_LOC_815/Y 0.01fF
C47799 OR2X1_LOC_324/a_8_216# OR2X1_LOC_532/B 0.01fF
C47800 OR2X1_LOC_665/Y OR2X1_LOC_666/Y 0.06fF
C47801 OR2X1_LOC_517/A AND2X1_LOC_866/A 0.03fF
C47802 OR2X1_LOC_13/B AND2X1_LOC_773/a_8_24# 0.03fF
C47803 OR2X1_LOC_229/Y OR2X1_LOC_52/B 0.01fF
C47804 OR2X1_LOC_643/Y OR2X1_LOC_340/Y 0.02fF
C47805 AND2X1_LOC_139/A AND2X1_LOC_139/a_8_24# 0.01fF
C47806 AND2X1_LOC_840/a_8_24# OR2X1_LOC_31/Y 0.26fF
C47807 AND2X1_LOC_154/Y OR2X1_LOC_7/A 0.22fF
C47808 OR2X1_LOC_222/a_8_216# OR2X1_LOC_475/B 0.01fF
C47809 OR2X1_LOC_256/A OR2X1_LOC_256/a_8_216# 0.08fF
C47810 AND2X1_LOC_675/A OR2X1_LOC_48/B 0.20fF
C47811 AND2X1_LOC_41/A OR2X1_LOC_214/B 0.05fF
C47812 INPUT_0 OR2X1_LOC_194/a_8_216# 0.01fF
C47813 OR2X1_LOC_517/Y OR2X1_LOC_22/Y 0.03fF
C47814 AND2X1_LOC_773/Y OR2X1_LOC_13/B 0.74fF
C47815 OR2X1_LOC_71/Y OR2X1_LOC_39/A 0.23fF
C47816 AND2X1_LOC_41/A OR2X1_LOC_241/B 0.41fF
C47817 OR2X1_LOC_18/Y AND2X1_LOC_675/A 0.06fF
C47818 OR2X1_LOC_377/A AND2X1_LOC_47/Y 0.13fF
C47819 AND2X1_LOC_657/Y AND2X1_LOC_222/Y 0.03fF
C47820 OR2X1_LOC_401/A AND2X1_LOC_3/Y 0.56fF
C47821 OR2X1_LOC_293/a_36_216# OR2X1_LOC_753/A 0.00fF
C47822 OR2X1_LOC_95/Y AND2X1_LOC_447/a_8_24# 0.01fF
C47823 OR2X1_LOC_109/Y AND2X1_LOC_841/a_8_24# 0.01fF
C47824 OR2X1_LOC_47/Y OR2X1_LOC_40/a_8_216# 0.11fF
C47825 AND2X1_LOC_318/Y OR2X1_LOC_619/Y 0.02fF
C47826 AND2X1_LOC_47/Y AND2X1_LOC_824/B 0.00fF
C47827 OR2X1_LOC_131/Y AND2X1_LOC_663/B 0.05fF
C47828 OR2X1_LOC_77/a_36_216# OR2X1_LOC_820/B 0.00fF
C47829 AND2X1_LOC_634/Y AND2X1_LOC_852/Y 0.03fF
C47830 AND2X1_LOC_653/B AND2X1_LOC_810/Y 0.05fF
C47831 OR2X1_LOC_92/Y OR2X1_LOC_597/Y 0.04fF
C47832 AND2X1_LOC_866/A AND2X1_LOC_624/A 0.03fF
C47833 AND2X1_LOC_354/Y AND2X1_LOC_798/A 0.01fF
C47834 OR2X1_LOC_31/Y OR2X1_LOC_511/Y 0.03fF
C47835 OR2X1_LOC_199/a_8_216# OR2X1_LOC_199/B 0.01fF
C47836 AND2X1_LOC_95/Y OR2X1_LOC_112/B 0.02fF
C47837 AND2X1_LOC_64/Y OR2X1_LOC_502/Y 0.02fF
C47838 D_INPUT_0 AND2X1_LOC_853/Y 0.10fF
C47839 AND2X1_LOC_47/Y OR2X1_LOC_203/Y 0.07fF
C47840 OR2X1_LOC_851/A OR2X1_LOC_804/A 0.01fF
C47841 OR2X1_LOC_733/a_8_216# OR2X1_LOC_733/Y 0.01fF
C47842 AND2X1_LOC_40/Y OR2X1_LOC_551/B 0.02fF
C47843 AND2X1_LOC_92/Y OR2X1_LOC_341/a_36_216# 0.00fF
C47844 OR2X1_LOC_743/A OR2X1_LOC_22/Y 0.28fF
C47845 AND2X1_LOC_733/Y AND2X1_LOC_222/Y 0.01fF
C47846 INPUT_1 OR2X1_LOC_7/A 0.22fF
C47847 OR2X1_LOC_114/B OR2X1_LOC_501/a_8_216# 0.01fF
C47848 AND2X1_LOC_243/Y OR2X1_LOC_13/B 0.08fF
C47849 VDD OR2X1_LOC_385/a_8_216# 0.00fF
C47850 OR2X1_LOC_39/A D_INPUT_1 0.13fF
C47851 OR2X1_LOC_3/Y OR2X1_LOC_7/Y 0.01fF
C47852 AND2X1_LOC_359/B D_INPUT_3 0.07fF
C47853 AND2X1_LOC_69/Y OR2X1_LOC_814/A 0.03fF
C47854 AND2X1_LOC_18/Y D_GATE_366 0.21fF
C47855 OR2X1_LOC_756/B OR2X1_LOC_578/B 0.03fF
C47856 AND2X1_LOC_476/A OR2X1_LOC_690/A 0.04fF
C47857 OR2X1_LOC_419/Y AND2X1_LOC_621/Y 0.03fF
C47858 VDD OR2X1_LOC_376/Y -0.00fF
C47859 OR2X1_LOC_66/A OR2X1_LOC_112/A 0.39fF
C47860 OR2X1_LOC_755/A AND2X1_LOC_814/a_36_24# 0.00fF
C47861 OR2X1_LOC_212/A OR2X1_LOC_365/B 0.02fF
C47862 AND2X1_LOC_22/Y OR2X1_LOC_338/A 0.83fF
C47863 VDD OR2X1_LOC_590/Y 0.15fF
C47864 OR2X1_LOC_377/A OR2X1_LOC_598/A 0.49fF
C47865 OR2X1_LOC_664/Y AND2X1_LOC_72/B 0.03fF
C47866 OR2X1_LOC_151/A OR2X1_LOC_319/Y 0.10fF
C47867 AND2X1_LOC_348/Y AND2X1_LOC_721/A 0.00fF
C47868 OR2X1_LOC_415/Y OR2X1_LOC_548/a_8_216# 0.01fF
C47869 AND2X1_LOC_824/B OR2X1_LOC_598/A 0.21fF
C47870 AND2X1_LOC_64/Y AND2X1_LOC_433/a_36_24# 0.01fF
C47871 OR2X1_LOC_22/Y OR2X1_LOC_246/A 1.33fF
C47872 AND2X1_LOC_721/A OR2X1_LOC_753/A 0.27fF
C47873 OR2X1_LOC_207/B AND2X1_LOC_7/B 0.03fF
C47874 OR2X1_LOC_203/Y OR2X1_LOC_598/A 0.21fF
C47875 AND2X1_LOC_425/Y OR2X1_LOC_707/B 0.01fF
C47876 AND2X1_LOC_79/a_8_24# OR2X1_LOC_532/B 0.01fF
C47877 AND2X1_LOC_621/Y OR2X1_LOC_152/A 0.03fF
C47878 AND2X1_LOC_211/B OR2X1_LOC_173/a_8_216# 0.01fF
C47879 AND2X1_LOC_56/B OR2X1_LOC_543/a_8_216# 0.01fF
C47880 AND2X1_LOC_552/a_8_24# AND2X1_LOC_552/A 0.19fF
C47881 OR2X1_LOC_186/Y AND2X1_LOC_22/Y 0.00fF
C47882 OR2X1_LOC_516/Y AND2X1_LOC_500/Y 0.24fF
C47883 AND2X1_LOC_474/a_8_24# AND2X1_LOC_657/A 0.01fF
C47884 OR2X1_LOC_696/A VDD 1.03fF
C47885 AND2X1_LOC_57/Y OR2X1_LOC_66/A 0.05fF
C47886 OR2X1_LOC_168/B OR2X1_LOC_593/B 0.03fF
C47887 OR2X1_LOC_473/A AND2X1_LOC_67/Y 0.31fF
C47888 OR2X1_LOC_392/B OR2X1_LOC_113/B 0.05fF
C47889 OR2X1_LOC_468/A OR2X1_LOC_388/a_36_216# -0.00fF
C47890 OR2X1_LOC_561/Y OR2X1_LOC_579/A 0.01fF
C47891 OR2X1_LOC_287/a_8_216# OR2X1_LOC_532/B 0.01fF
C47892 OR2X1_LOC_121/Y AND2X1_LOC_44/Y 0.01fF
C47893 OR2X1_LOC_45/B AND2X1_LOC_339/B 0.03fF
C47894 AND2X1_LOC_370/a_8_24# AND2X1_LOC_182/a_8_24# 0.23fF
C47895 OR2X1_LOC_22/Y OR2X1_LOC_409/B 0.03fF
C47896 AND2X1_LOC_64/Y VDD 1.51fF
C47897 OR2X1_LOC_186/Y AND2X1_LOC_417/a_36_24# 0.00fF
C47898 AND2X1_LOC_866/A AND2X1_LOC_621/a_8_24# 0.02fF
C47899 OR2X1_LOC_243/A OR2X1_LOC_71/A 0.00fF
C47900 AND2X1_LOC_477/A AND2X1_LOC_810/Y 0.07fF
C47901 OR2X1_LOC_351/B AND2X1_LOC_44/Y 0.07fF
C47902 INPUT_5 D_INPUT_6 0.08fF
C47903 OR2X1_LOC_139/A OR2X1_LOC_641/A 0.02fF
C47904 AND2X1_LOC_383/a_8_24# VDD -0.00fF
C47905 AND2X1_LOC_715/Y VDD 1.06fF
C47906 AND2X1_LOC_12/Y OR2X1_LOC_501/a_8_216# 0.04fF
C47907 OR2X1_LOC_742/B OR2X1_LOC_551/a_36_216# 0.02fF
C47908 OR2X1_LOC_76/Y OR2X1_LOC_578/B 0.03fF
C47909 AND2X1_LOC_50/Y INPUT_6 0.03fF
C47910 OR2X1_LOC_40/Y AND2X1_LOC_341/a_8_24# 0.02fF
C47911 AND2X1_LOC_12/Y OR2X1_LOC_580/A 0.07fF
C47912 OR2X1_LOC_148/Y OR2X1_LOC_149/a_8_216# 0.39fF
C47913 OR2X1_LOC_19/B OR2X1_LOC_29/a_8_216# 0.01fF
C47914 OR2X1_LOC_114/B AND2X1_LOC_44/Y 0.01fF
C47915 AND2X1_LOC_672/B D_INPUT_1 0.46fF
C47916 OR2X1_LOC_738/A OR2X1_LOC_550/B 0.03fF
C47917 OR2X1_LOC_421/A AND2X1_LOC_771/a_8_24# 0.01fF
C47918 OR2X1_LOC_36/Y OR2X1_LOC_71/A 0.02fF
C47919 OR2X1_LOC_744/A AND2X1_LOC_465/A 0.16fF
C47920 OR2X1_LOC_570/A OR2X1_LOC_562/A 0.00fF
C47921 OR2X1_LOC_160/B OR2X1_LOC_161/B 0.26fF
C47922 AND2X1_LOC_555/Y OR2X1_LOC_292/a_36_216# 0.00fF
C47923 AND2X1_LOC_799/a_8_24# OR2X1_LOC_744/A 0.01fF
C47924 OR2X1_LOC_756/B OR2X1_LOC_366/A 0.02fF
C47925 OR2X1_LOC_539/Y OR2X1_LOC_332/a_36_216# 0.00fF
C47926 OR2X1_LOC_31/Y AND2X1_LOC_648/B 0.03fF
C47927 VDD AND2X1_LOC_82/Y 0.16fF
C47928 OR2X1_LOC_325/B OR2X1_LOC_439/B 0.03fF
C47929 AND2X1_LOC_342/a_8_24# OR2X1_LOC_13/B 0.24fF
C47930 D_INPUT_0 OR2X1_LOC_396/Y 0.15fF
C47931 AND2X1_LOC_59/Y OR2X1_LOC_593/B 0.03fF
C47932 OR2X1_LOC_188/Y AND2X1_LOC_41/A 0.01fF
C47933 AND2X1_LOC_11/Y AND2X1_LOC_762/a_8_24# 0.11fF
C47934 AND2X1_LOC_649/Y AND2X1_LOC_655/a_36_24# 0.00fF
C47935 OR2X1_LOC_40/Y AND2X1_LOC_778/Y 0.00fF
C47936 AND2X1_LOC_364/Y OR2X1_LOC_428/A 0.03fF
C47937 OR2X1_LOC_538/A AND2X1_LOC_44/Y 0.00fF
C47938 OR2X1_LOC_201/A AND2X1_LOC_7/B 0.01fF
C47939 AND2X1_LOC_663/B AND2X1_LOC_657/A 0.10fF
C47940 OR2X1_LOC_696/A OR2X1_LOC_829/a_8_216# 0.06fF
C47941 OR2X1_LOC_185/A AND2X1_LOC_235/a_8_24# 0.01fF
C47942 AND2X1_LOC_355/a_8_24# OR2X1_LOC_13/B 0.01fF
C47943 OR2X1_LOC_449/A OR2X1_LOC_712/B -0.00fF
C47944 OR2X1_LOC_532/B OR2X1_LOC_374/Y 0.04fF
C47945 OR2X1_LOC_40/Y AND2X1_LOC_709/a_8_24# 0.01fF
C47946 AND2X1_LOC_787/A OR2X1_LOC_165/Y 0.21fF
C47947 OR2X1_LOC_696/A OR2X1_LOC_315/Y 0.03fF
C47948 VDD AND2X1_LOC_86/a_8_24# -0.00fF
C47949 OR2X1_LOC_476/B OR2X1_LOC_68/B 0.34fF
C47950 OR2X1_LOC_762/Y OR2X1_LOC_12/Y 0.04fF
C47951 AND2X1_LOC_719/Y OR2X1_LOC_56/A 0.03fF
C47952 D_INPUT_5 AND2X1_LOC_44/Y 0.03fF
C47953 OR2X1_LOC_650/Y OR2X1_LOC_68/B 0.03fF
C47954 OR2X1_LOC_6/B OR2X1_LOC_51/Y 0.05fF
C47955 OR2X1_LOC_759/A OR2X1_LOC_600/A 0.18fF
C47956 OR2X1_LOC_710/A OR2X1_LOC_161/A 0.02fF
C47957 AND2X1_LOC_91/B OR2X1_LOC_405/A 0.55fF
C47958 AND2X1_LOC_663/A AND2X1_LOC_477/Y 0.10fF
C47959 OR2X1_LOC_78/A OR2X1_LOC_307/A 0.01fF
C47960 OR2X1_LOC_18/Y AND2X1_LOC_241/a_8_24# 0.00fF
C47961 AND2X1_LOC_658/B AND2X1_LOC_658/a_8_24# 0.01fF
C47962 AND2X1_LOC_59/Y AND2X1_LOC_273/a_8_24# 0.01fF
C47963 OR2X1_LOC_609/Y AND2X1_LOC_646/a_8_24# 0.01fF
C47964 AND2X1_LOC_539/Y OR2X1_LOC_306/a_8_216# 0.48fF
C47965 OR2X1_LOC_409/B OR2X1_LOC_387/a_8_216# 0.00fF
C47966 OR2X1_LOC_304/a_8_216# OR2X1_LOC_45/Y 0.03fF
C47967 OR2X1_LOC_158/A AND2X1_LOC_860/a_8_24# 0.01fF
C47968 OR2X1_LOC_6/B OR2X1_LOC_78/B 0.13fF
C47969 AND2X1_LOC_595/a_36_24# OR2X1_LOC_244/Y 0.00fF
C47970 OR2X1_LOC_865/B OR2X1_LOC_474/B 0.04fF
C47971 OR2X1_LOC_111/Y AND2X1_LOC_222/Y 0.41fF
C47972 AND2X1_LOC_716/Y OR2X1_LOC_12/Y 0.07fF
C47973 OR2X1_LOC_177/Y OR2X1_LOC_438/Y 0.41fF
C47974 AND2X1_LOC_675/Y AND2X1_LOC_500/B 0.82fF
C47975 AND2X1_LOC_22/a_8_24# AND2X1_LOC_44/Y 0.02fF
C47976 AND2X1_LOC_554/Y AND2X1_LOC_554/a_8_24# 0.03fF
C47977 OR2X1_LOC_375/A OR2X1_LOC_120/a_36_216# 0.00fF
C47978 OR2X1_LOC_450/a_36_216# OR2X1_LOC_467/A -0.00fF
C47979 OR2X1_LOC_185/Y OR2X1_LOC_140/B 0.05fF
C47980 OR2X1_LOC_604/A OR2X1_LOC_820/A 0.02fF
C47981 AND2X1_LOC_654/Y OR2X1_LOC_12/Y 0.09fF
C47982 OR2X1_LOC_696/A OR2X1_LOC_251/Y 0.50fF
C47983 AND2X1_LOC_86/Y OR2X1_LOC_161/B 0.06fF
C47984 OR2X1_LOC_137/a_8_216# AND2X1_LOC_18/Y 0.01fF
C47985 OR2X1_LOC_833/Y OR2X1_LOC_737/A 0.02fF
C47986 OR2X1_LOC_160/A OR2X1_LOC_97/A 0.06fF
C47987 OR2X1_LOC_40/Y OR2X1_LOC_517/A 0.10fF
C47988 OR2X1_LOC_22/Y OR2X1_LOC_599/a_8_216# 0.05fF
C47989 AND2X1_LOC_658/B AND2X1_LOC_735/Y 0.01fF
C47990 AND2X1_LOC_12/Y AND2X1_LOC_44/Y 0.20fF
C47991 AND2X1_LOC_203/Y AND2X1_LOC_204/Y 0.28fF
C47992 AND2X1_LOC_850/A AND2X1_LOC_860/A 0.14fF
C47993 OR2X1_LOC_169/a_8_216# OR2X1_LOC_175/Y 0.04fF
C47994 OR2X1_LOC_175/Y OR2X1_LOC_802/Y 0.19fF
C47995 AND2X1_LOC_164/a_8_24# OR2X1_LOC_648/A 0.04fF
C47996 OR2X1_LOC_45/B AND2X1_LOC_633/a_8_24# 0.01fF
C47997 OR2X1_LOC_6/B OR2X1_LOC_721/Y 0.10fF
C47998 OR2X1_LOC_698/Y OR2X1_LOC_600/A 0.00fF
C47999 AND2X1_LOC_81/B AND2X1_LOC_22/Y 0.03fF
C48000 OR2X1_LOC_863/a_8_216# OR2X1_LOC_175/Y 0.04fF
C48001 OR2X1_LOC_175/Y OR2X1_LOC_468/Y 0.03fF
C48002 OR2X1_LOC_151/A OR2X1_LOC_811/A 0.03fF
C48003 OR2X1_LOC_40/Y AND2X1_LOC_865/a_36_24# 0.01fF
C48004 OR2X1_LOC_696/A AND2X1_LOC_389/a_8_24# 0.01fF
C48005 OR2X1_LOC_427/A AND2X1_LOC_476/Y 1.01fF
C48006 AND2X1_LOC_362/B OR2X1_LOC_427/A 0.04fF
C48007 OR2X1_LOC_692/Y AND2X1_LOC_648/a_8_24# 0.02fF
C48008 OR2X1_LOC_739/A OR2X1_LOC_355/a_36_216# 0.00fF
C48009 OR2X1_LOC_656/Y VDD 0.27fF
C48010 OR2X1_LOC_177/a_8_216# AND2X1_LOC_624/A 0.06fF
C48011 OR2X1_LOC_177/Y AND2X1_LOC_621/Y 0.03fF
C48012 OR2X1_LOC_325/a_8_216# AND2X1_LOC_110/Y 0.01fF
C48013 OR2X1_LOC_175/Y AND2X1_LOC_385/a_8_24# 0.01fF
C48014 OR2X1_LOC_553/A OR2X1_LOC_161/B 0.07fF
C48015 OR2X1_LOC_40/Y AND2X1_LOC_833/a_8_24# 0.01fF
C48016 OR2X1_LOC_269/B OR2X1_LOC_563/A 0.07fF
C48017 OR2X1_LOC_161/A OR2X1_LOC_356/A 0.11fF
C48018 OR2X1_LOC_673/Y OR2X1_LOC_721/a_8_216# 0.01fF
C48019 OR2X1_LOC_105/Y OR2X1_LOC_66/A 0.00fF
C48020 OR2X1_LOC_802/Y AND2X1_LOC_417/a_8_24# 0.04fF
C48021 OR2X1_LOC_266/a_8_216# OR2X1_LOC_161/B 0.01fF
C48022 AND2X1_LOC_512/Y AND2X1_LOC_434/Y 0.54fF
C48023 OR2X1_LOC_499/B AND2X1_LOC_92/Y 0.01fF
C48024 AND2X1_LOC_7/a_36_24# AND2X1_LOC_7/B 0.01fF
C48025 OR2X1_LOC_377/A OR2X1_LOC_646/B 0.03fF
C48026 OR2X1_LOC_604/A OR2X1_LOC_427/Y 0.02fF
C48027 OR2X1_LOC_44/Y AND2X1_LOC_219/A 0.08fF
C48028 OR2X1_LOC_492/Y OR2X1_LOC_39/A 0.16fF
C48029 AND2X1_LOC_71/a_8_24# OR2X1_LOC_632/Y 0.02fF
C48030 VDD OR2X1_LOC_695/a_8_216# 0.00fF
C48031 OR2X1_LOC_106/Y AND2X1_LOC_116/Y 0.00fF
C48032 AND2X1_LOC_367/B OR2X1_LOC_92/Y 0.01fF
C48033 AND2X1_LOC_584/a_36_24# AND2X1_LOC_1/Y 0.00fF
C48034 AND2X1_LOC_185/a_8_24# OR2X1_LOC_59/Y 0.02fF
C48035 OR2X1_LOC_493/B OR2X1_LOC_737/A 0.11fF
C48036 VDD OR2X1_LOC_807/Y 0.05fF
C48037 AND2X1_LOC_3/Y AND2X1_LOC_7/B 5.25fF
C48038 OR2X1_LOC_532/B OR2X1_LOC_532/a_36_216# 0.00fF
C48039 AND2X1_LOC_702/Y OR2X1_LOC_135/Y 0.79fF
C48040 OR2X1_LOC_516/A AND2X1_LOC_784/Y 0.02fF
C48041 OR2X1_LOC_647/B AND2X1_LOC_7/B 0.07fF
C48042 OR2X1_LOC_160/B AND2X1_LOC_536/a_8_24# 0.01fF
C48043 OR2X1_LOC_667/Y OR2X1_LOC_51/Y 0.02fF
C48044 OR2X1_LOC_604/A AND2X1_LOC_621/Y 0.09fF
C48045 OR2X1_LOC_40/Y AND2X1_LOC_862/A 0.01fF
C48046 OR2X1_LOC_40/Y AND2X1_LOC_624/A 0.08fF
C48047 OR2X1_LOC_710/A AND2X1_LOC_51/Y 0.00fF
C48048 OR2X1_LOC_51/Y OR2X1_LOC_625/a_8_216# 0.01fF
C48049 AND2X1_LOC_59/Y AND2X1_LOC_41/a_8_24# 0.03fF
C48050 OR2X1_LOC_748/A OR2X1_LOC_381/a_8_216# 0.39fF
C48051 OR2X1_LOC_6/B OR2X1_LOC_375/A 0.17fF
C48052 VDD OR2X1_LOC_555/B 0.26fF
C48053 OR2X1_LOC_450/B AND2X1_LOC_426/a_8_24# 0.01fF
C48054 AND2X1_LOC_634/a_8_24# OR2X1_LOC_16/A 0.00fF
C48055 OR2X1_LOC_671/Y OR2X1_LOC_42/a_8_216# 0.15fF
C48056 AND2X1_LOC_41/A OR2X1_LOC_469/Y 0.07fF
C48057 AND2X1_LOC_8/Y AND2X1_LOC_65/A 0.01fF
C48058 OR2X1_LOC_600/A AND2X1_LOC_838/Y 0.79fF
C48059 OR2X1_LOC_477/B OR2X1_LOC_467/B 0.13fF
C48060 AND2X1_LOC_523/a_8_24# OR2X1_LOC_744/A 0.05fF
C48061 OR2X1_LOC_756/B OR2X1_LOC_814/a_8_216# 0.03fF
C48062 VDD AND2X1_LOC_458/Y 0.24fF
C48063 AND2X1_LOC_118/a_8_24# OR2X1_LOC_549/A 0.01fF
C48064 OR2X1_LOC_217/Y OR2X1_LOC_507/A 0.03fF
C48065 AND2X1_LOC_798/a_36_24# OR2X1_LOC_22/Y 0.01fF
C48066 AND2X1_LOC_50/Y OR2X1_LOC_638/a_36_216# 0.00fF
C48067 AND2X1_LOC_753/B OR2X1_LOC_638/a_8_216# 0.48fF
C48068 AND2X1_LOC_705/Y OR2X1_LOC_420/Y 0.02fF
C48069 OR2X1_LOC_426/B OR2X1_LOC_39/A 0.12fF
C48070 OR2X1_LOC_252/Y OR2X1_LOC_56/A 0.02fF
C48071 OR2X1_LOC_158/B AND2X1_LOC_210/a_8_24# 0.01fF
C48072 OR2X1_LOC_56/A AND2X1_LOC_655/A 0.03fF
C48073 OR2X1_LOC_43/A AND2X1_LOC_200/a_8_24# 0.01fF
C48074 VDD AND2X1_LOC_369/a_8_24# 0.00fF
C48075 AND2X1_LOC_130/a_8_24# OR2X1_LOC_7/A 0.03fF
C48076 OR2X1_LOC_831/A OR2X1_LOC_787/Y 0.01fF
C48077 OR2X1_LOC_273/Y OR2X1_LOC_16/A 0.06fF
C48078 OR2X1_LOC_154/A OR2X1_LOC_35/Y 0.08fF
C48079 OR2X1_LOC_335/a_8_216# OR2X1_LOC_335/B 0.07fF
C48080 OR2X1_LOC_91/A OR2X1_LOC_316/Y 0.03fF
C48081 AND2X1_LOC_594/a_8_24# OR2X1_LOC_435/Y 0.24fF
C48082 AND2X1_LOC_577/a_8_24# OR2X1_LOC_189/A 0.08fF
C48083 D_GATE_662 OR2X1_LOC_624/B 0.01fF
C48084 AND2X1_LOC_658/A OR2X1_LOC_44/Y 0.03fF
C48085 OR2X1_LOC_17/a_8_216# D_INPUT_6 0.08fF
C48086 OR2X1_LOC_692/a_8_216# OR2X1_LOC_48/B 0.03fF
C48087 AND2X1_LOC_744/a_8_24# OR2X1_LOC_160/A 0.04fF
C48088 OR2X1_LOC_448/A OR2X1_LOC_784/Y 0.10fF
C48089 AND2X1_LOC_22/Y OR2X1_LOC_196/B 0.02fF
C48090 OR2X1_LOC_796/B OR2X1_LOC_712/B 0.00fF
C48091 OR2X1_LOC_123/a_8_216# OR2X1_LOC_864/A 0.04fF
C48092 OR2X1_LOC_92/Y OR2X1_LOC_48/B 0.13fF
C48093 OR2X1_LOC_64/Y OR2X1_LOC_766/a_8_216# 0.03fF
C48094 VDD OR2X1_LOC_32/Y 0.11fF
C48095 OR2X1_LOC_692/a_8_216# OR2X1_LOC_18/Y 0.02fF
C48096 OR2X1_LOC_36/Y OR2X1_LOC_59/Y 3.70fF
C48097 VDD OR2X1_LOC_89/a_8_216# 0.21fF
C48098 OR2X1_LOC_507/B OR2X1_LOC_502/A 0.40fF
C48099 AND2X1_LOC_81/B OR2X1_LOC_244/B 0.03fF
C48100 AND2X1_LOC_51/Y OR2X1_LOC_356/A 0.25fF
C48101 OR2X1_LOC_18/Y OR2X1_LOC_92/Y 0.30fF
C48102 INPUT_1 AND2X1_LOC_476/a_8_24# 0.01fF
C48103 OR2X1_LOC_91/A AND2X1_LOC_354/B 0.07fF
C48104 AND2X1_LOC_723/a_8_24# AND2X1_LOC_168/Y 0.01fF
C48105 OR2X1_LOC_335/A OR2X1_LOC_440/A 0.03fF
C48106 OR2X1_LOC_19/B OR2X1_LOC_16/A 0.07fF
C48107 OR2X1_LOC_31/Y OR2X1_LOC_56/a_8_216# 0.14fF
C48108 OR2X1_LOC_26/Y AND2X1_LOC_637/a_8_24# 0.01fF
C48109 OR2X1_LOC_462/B OR2X1_LOC_634/A 0.05fF
C48110 AND2X1_LOC_218/a_8_24# AND2X1_LOC_116/Y 0.01fF
C48111 OR2X1_LOC_743/a_8_216# OR2X1_LOC_52/B 0.03fF
C48112 OR2X1_LOC_46/A AND2X1_LOC_786/Y 0.02fF
C48113 AND2X1_LOC_211/B OR2X1_LOC_426/B 0.09fF
C48114 OR2X1_LOC_532/B OR2X1_LOC_392/B 0.06fF
C48115 OR2X1_LOC_31/Y AND2X1_LOC_465/A 0.05fF
C48116 OR2X1_LOC_123/a_8_216# OR2X1_LOC_633/B 0.14fF
C48117 OR2X1_LOC_377/A OR2X1_LOC_400/a_36_216# 0.01fF
C48118 OR2X1_LOC_160/A OR2X1_LOC_475/B 0.03fF
C48119 AND2X1_LOC_652/a_8_24# OR2X1_LOC_594/Y 0.01fF
C48120 AND2X1_LOC_12/Y OR2X1_LOC_61/a_8_216# 0.05fF
C48121 OR2X1_LOC_158/A OR2X1_LOC_275/a_8_216# 0.02fF
C48122 AND2X1_LOC_191/B OR2X1_LOC_757/a_8_216# 0.01fF
C48123 OR2X1_LOC_828/a_36_216# OR2X1_LOC_828/B 0.00fF
C48124 OR2X1_LOC_529/Y OR2X1_LOC_51/Y 0.54fF
C48125 OR2X1_LOC_709/B AND2X1_LOC_698/a_8_24# 0.01fF
C48126 INPUT_0 OR2X1_LOC_690/A 0.82fF
C48127 OR2X1_LOC_600/Y OR2X1_LOC_485/A 0.01fF
C48128 OR2X1_LOC_40/Y AND2X1_LOC_650/a_36_24# 0.00fF
C48129 AND2X1_LOC_552/a_36_24# OR2X1_LOC_31/Y 0.00fF
C48130 OR2X1_LOC_31/Y AND2X1_LOC_231/a_8_24# 0.01fF
C48131 OR2X1_LOC_494/a_8_216# AND2X1_LOC_359/B 0.01fF
C48132 AND2X1_LOC_850/a_36_24# AND2X1_LOC_850/Y 0.01fF
C48133 OR2X1_LOC_18/Y OR2X1_LOC_257/a_8_216# 0.02fF
C48134 VDD AND2X1_LOC_797/A 0.21fF
C48135 AND2X1_LOC_59/Y AND2X1_LOC_492/a_8_24# 0.01fF
C48136 OR2X1_LOC_405/A OR2X1_LOC_799/A 0.03fF
C48137 AND2X1_LOC_800/a_8_24# OR2X1_LOC_16/A 0.01fF
C48138 OR2X1_LOC_244/A OR2X1_LOC_161/B 0.05fF
C48139 AND2X1_LOC_81/B OR2X1_LOC_608/a_36_216# 0.00fF
C48140 OR2X1_LOC_74/A AND2X1_LOC_469/B 0.03fF
C48141 AND2X1_LOC_734/Y OR2X1_LOC_52/B 0.00fF
C48142 VDD AND2X1_LOC_663/B 1.66fF
C48143 OR2X1_LOC_701/Y AND2X1_LOC_847/Y 0.02fF
C48144 AND2X1_LOC_95/Y OR2X1_LOC_39/A 0.03fF
C48145 OR2X1_LOC_18/Y OR2X1_LOC_65/B 0.05fF
C48146 OR2X1_LOC_335/Y OR2X1_LOC_787/Y 0.00fF
C48147 OR2X1_LOC_190/A OR2X1_LOC_254/a_36_216# 0.02fF
C48148 OR2X1_LOC_91/Y AND2X1_LOC_97/a_8_24# 0.00fF
C48149 OR2X1_LOC_619/Y AND2X1_LOC_470/B 0.01fF
C48150 OR2X1_LOC_648/B AND2X1_LOC_48/A 0.02fF
C48151 OR2X1_LOC_614/a_36_216# AND2X1_LOC_51/Y -0.00fF
C48152 OR2X1_LOC_756/B OR2X1_LOC_654/A 0.07fF
C48153 AND2X1_LOC_390/B OR2X1_LOC_91/A 0.07fF
C48154 AND2X1_LOC_43/B OR2X1_LOC_161/A 0.22fF
C48155 OR2X1_LOC_773/Y D_INPUT_1 0.05fF
C48156 AND2X1_LOC_99/A OR2X1_LOC_67/a_36_216# 0.00fF
C48157 OR2X1_LOC_624/A OR2X1_LOC_510/Y 0.03fF
C48158 OR2X1_LOC_517/A OR2X1_LOC_7/A 0.15fF
C48159 OR2X1_LOC_417/Y AND2X1_LOC_436/Y 0.03fF
C48160 AND2X1_LOC_733/Y OR2X1_LOC_74/A 0.54fF
C48161 AND2X1_LOC_22/Y OR2X1_LOC_112/B 0.31fF
C48162 OR2X1_LOC_270/Y AND2X1_LOC_7/B 0.04fF
C48163 AND2X1_LOC_91/B OR2X1_LOC_330/a_8_216# 0.04fF
C48164 OR2X1_LOC_377/A AND2X1_LOC_82/a_8_24# 0.01fF
C48165 VDD AND2X1_LOC_686/a_8_24# 0.00fF
C48166 AND2X1_LOC_56/B OR2X1_LOC_181/B 0.07fF
C48167 OR2X1_LOC_75/Y OR2X1_LOC_16/A 0.04fF
C48168 AND2X1_LOC_194/a_8_24# OR2X1_LOC_3/Y 0.01fF
C48169 OR2X1_LOC_18/Y AND2X1_LOC_464/a_36_24# 0.00fF
C48170 AND2X1_LOC_12/Y OR2X1_LOC_848/a_8_216# 0.00fF
C48171 OR2X1_LOC_385/Y OR2X1_LOC_92/Y 0.59fF
C48172 OR2X1_LOC_185/A OR2X1_LOC_87/A 0.56fF
C48173 OR2X1_LOC_814/A AND2X1_LOC_18/Y 0.67fF
C48174 OR2X1_LOC_256/a_8_216# OR2X1_LOC_248/Y 0.02fF
C48175 OR2X1_LOC_271/B OR2X1_LOC_315/Y 0.01fF
C48176 AND2X1_LOC_847/Y OR2X1_LOC_44/Y 0.06fF
C48177 AND2X1_LOC_729/Y AND2X1_LOC_319/A 0.02fF
C48178 OR2X1_LOC_793/A OR2X1_LOC_793/a_8_216# 0.01fF
C48179 AND2X1_LOC_374/a_8_24# OR2X1_LOC_280/Y 0.02fF
C48180 OR2X1_LOC_517/Y OR2X1_LOC_39/A 0.04fF
C48181 AND2X1_LOC_347/Y AND2X1_LOC_347/a_36_24# 0.00fF
C48182 INPUT_0 OR2X1_LOC_64/Y 0.07fF
C48183 AND2X1_LOC_41/A OR2X1_LOC_193/A 0.01fF
C48184 OR2X1_LOC_271/Y OR2X1_LOC_18/Y 0.26fF
C48185 OR2X1_LOC_574/A OR2X1_LOC_737/A 0.10fF
C48186 AND2X1_LOC_7/B OR2X1_LOC_194/a_8_216# 0.01fF
C48187 AND2X1_LOC_571/B AND2X1_LOC_563/Y 0.01fF
C48188 OR2X1_LOC_743/A OR2X1_LOC_422/a_36_216# 0.00fF
C48189 OR2X1_LOC_43/A AND2X1_LOC_452/Y 0.00fF
C48190 OR2X1_LOC_835/B OR2X1_LOC_130/A 0.04fF
C48191 OR2X1_LOC_659/B OR2X1_LOC_659/a_8_216# 0.06fF
C48192 OR2X1_LOC_46/A AND2X1_LOC_218/Y 0.00fF
C48193 AND2X1_LOC_101/a_8_24# OR2X1_LOC_91/A 0.02fF
C48194 OR2X1_LOC_808/B OR2X1_LOC_705/Y 0.06fF
C48195 OR2X1_LOC_624/A OR2X1_LOC_810/A 0.01fF
C48196 OR2X1_LOC_756/B AND2X1_LOC_261/a_36_24# 0.00fF
C48197 OR2X1_LOC_471/Y OR2X1_LOC_803/A 0.02fF
C48198 AND2X1_LOC_337/B AND2X1_LOC_661/a_8_24# 0.11fF
C48199 AND2X1_LOC_95/Y OR2X1_LOC_574/A 0.03fF
C48200 OR2X1_LOC_777/B AND2X1_LOC_246/a_8_24# 0.20fF
C48201 AND2X1_LOC_95/Y OR2X1_LOC_33/A 0.01fF
C48202 OR2X1_LOC_600/a_8_216# OR2X1_LOC_31/Y 0.07fF
C48203 OR2X1_LOC_664/Y OR2X1_LOC_346/B 1.29fF
C48204 OR2X1_LOC_196/B OR2X1_LOC_706/A 0.28fF
C48205 OR2X1_LOC_433/a_8_216# OR2X1_LOC_36/Y 0.01fF
C48206 OR2X1_LOC_7/A AND2X1_LOC_624/A 0.06fF
C48207 OR2X1_LOC_467/A OR2X1_LOC_780/B 0.00fF
C48208 OR2X1_LOC_473/A AND2X1_LOC_625/a_8_24# 0.12fF
C48209 OR2X1_LOC_805/A AND2X1_LOC_3/Y 0.22fF
C48210 AND2X1_LOC_40/Y OR2X1_LOC_647/a_8_216# 0.01fF
C48211 AND2X1_LOC_222/Y AND2X1_LOC_804/A 0.00fF
C48212 OR2X1_LOC_743/A OR2X1_LOC_39/A 1.05fF
C48213 AND2X1_LOC_692/a_8_24# OR2X1_LOC_706/A 0.01fF
C48214 OR2X1_LOC_600/A OR2X1_LOC_224/Y 0.01fF
C48215 OR2X1_LOC_524/Y OR2X1_LOC_679/A 0.03fF
C48216 OR2X1_LOC_529/Y OR2X1_LOC_680/A 0.00fF
C48217 INPUT_0 OR2X1_LOC_417/A 0.07fF
C48218 AND2X1_LOC_41/A D_INPUT_0 0.19fF
C48219 AND2X1_LOC_47/Y OR2X1_LOC_78/B 0.26fF
C48220 AND2X1_LOC_324/a_8_24# OR2X1_LOC_619/Y 0.02fF
C48221 OR2X1_LOC_91/A AND2X1_LOC_863/Y 0.05fF
C48222 AND2X1_LOC_252/a_8_24# OR2X1_LOC_269/B 0.01fF
C48223 OR2X1_LOC_691/Y OR2X1_LOC_750/Y 0.02fF
C48224 AND2X1_LOC_672/B AND2X1_LOC_414/a_8_24# 0.01fF
C48225 AND2X1_LOC_866/A OR2X1_LOC_755/a_8_216# 0.02fF
C48226 OR2X1_LOC_485/A OR2X1_LOC_591/A 0.09fF
C48227 OR2X1_LOC_316/Y OR2X1_LOC_27/Y 0.07fF
C48228 OR2X1_LOC_280/Y OR2X1_LOC_497/Y 0.15fF
C48229 AND2X1_LOC_43/B AND2X1_LOC_51/Y 0.21fF
C48230 OR2X1_LOC_592/a_8_216# OR2X1_LOC_593/A -0.00fF
C48231 OR2X1_LOC_616/Y AND2X1_LOC_663/B 0.00fF
C48232 OR2X1_LOC_121/B OR2X1_LOC_212/A 0.03fF
C48233 INPUT_1 OR2X1_LOC_46/a_8_216# 0.07fF
C48234 OR2X1_LOC_527/a_36_216# OR2X1_LOC_419/Y 0.15fF
C48235 AND2X1_LOC_862/a_8_24# OR2X1_LOC_74/A 0.05fF
C48236 D_INPUT_0 AND2X1_LOC_401/a_8_24# 0.03fF
C48237 OR2X1_LOC_235/B OR2X1_LOC_62/A 0.18fF
C48238 OR2X1_LOC_164/Y OR2X1_LOC_95/Y 0.03fF
C48239 OR2X1_LOC_70/Y OR2X1_LOC_36/Y 1.46fF
C48240 OR2X1_LOC_503/A OR2X1_LOC_64/Y 0.05fF
C48241 OR2X1_LOC_64/Y OR2X1_LOC_11/Y 0.04fF
C48242 AND2X1_LOC_8/Y OR2X1_LOC_204/a_8_216# 0.01fF
C48243 OR2X1_LOC_417/Y OR2X1_LOC_603/a_8_216# 0.01fF
C48244 AND2X1_LOC_717/Y OR2X1_LOC_417/A 0.02fF
C48245 AND2X1_LOC_211/B OR2X1_LOC_743/A 0.07fF
C48246 OR2X1_LOC_26/Y OR2X1_LOC_27/a_8_216# 0.00fF
C48247 AND2X1_LOC_847/a_36_24# OR2X1_LOC_820/B 0.00fF
C48248 OR2X1_LOC_246/A OR2X1_LOC_39/A 0.10fF
C48249 OR2X1_LOC_296/Y AND2X1_LOC_3/Y 0.03fF
C48250 AND2X1_LOC_560/B OR2X1_LOC_64/Y 0.01fF
C48251 AND2X1_LOC_390/a_8_24# OR2X1_LOC_331/Y 0.02fF
C48252 AND2X1_LOC_240/a_8_24# D_INPUT_1 0.01fF
C48253 OR2X1_LOC_319/a_36_216# OR2X1_LOC_532/B 0.00fF
C48254 OR2X1_LOC_235/B OR2X1_LOC_234/a_36_216# 0.00fF
C48255 OR2X1_LOC_127/Y INPUT_1 0.03fF
C48256 OR2X1_LOC_662/A D_INPUT_0 0.01fF
C48257 AND2X1_LOC_514/Y OR2X1_LOC_36/Y 0.05fF
C48258 OR2X1_LOC_419/Y OR2X1_LOC_59/Y 0.09fF
C48259 AND2X1_LOC_702/Y AND2X1_LOC_863/A 0.02fF
C48260 AND2X1_LOC_853/a_8_24# OR2X1_LOC_7/A 0.02fF
C48261 AND2X1_LOC_738/B OR2X1_LOC_331/a_8_216# 0.02fF
C48262 OR2X1_LOC_339/a_36_216# OR2X1_LOC_358/A 0.00fF
C48263 OR2X1_LOC_45/B OR2X1_LOC_300/Y 0.71fF
C48264 OR2X1_LOC_62/B OR2X1_LOC_204/Y 0.01fF
C48265 OR2X1_LOC_244/B OR2X1_LOC_66/Y 0.02fF
C48266 OR2X1_LOC_864/A OR2X1_LOC_750/A 0.13fF
C48267 OR2X1_LOC_78/B OR2X1_LOC_598/A 0.23fF
C48268 AND2X1_LOC_392/A AND2X1_LOC_657/A 0.07fF
C48269 OR2X1_LOC_18/Y AND2X1_LOC_849/a_36_24# 0.00fF
C48270 OR2X1_LOC_497/Y OR2X1_LOC_22/Y 0.03fF
C48271 OR2X1_LOC_628/a_8_216# OR2X1_LOC_615/Y 0.03fF
C48272 OR2X1_LOC_12/Y OR2X1_LOC_13/B 17.89fF
C48273 OR2X1_LOC_273/a_8_216# OR2X1_LOC_273/Y 0.02fF
C48274 OR2X1_LOC_16/A AND2X1_LOC_608/a_8_24# 0.01fF
C48275 OR2X1_LOC_541/A OR2X1_LOC_717/a_8_216# 0.49fF
C48276 AND2X1_LOC_47/Y OR2X1_LOC_375/A 1.06fF
C48277 OR2X1_LOC_636/B OR2X1_LOC_636/a_8_216# 0.01fF
C48278 OR2X1_LOC_280/Y AND2X1_LOC_844/a_8_24# 0.03fF
C48279 OR2X1_LOC_71/Y OR2X1_LOC_85/A 0.07fF
C48280 OR2X1_LOC_370/a_8_216# OR2X1_LOC_578/B 0.02fF
C48281 D_INPUT_0 OR2X1_LOC_824/Y 0.34fF
C48282 AND2X1_LOC_211/B OR2X1_LOC_246/A 0.10fF
C48283 AND2X1_LOC_546/a_36_24# AND2X1_LOC_796/Y 0.00fF
C48284 AND2X1_LOC_866/B AND2X1_LOC_793/Y 0.10fF
C48285 OR2X1_LOC_11/Y OR2X1_LOC_64/a_8_216# 0.01fF
C48286 OR2X1_LOC_40/a_8_216# OR2X1_LOC_3/B 0.02fF
C48287 AND2X1_LOC_70/a_8_24# AND2X1_LOC_31/Y 0.01fF
C48288 AND2X1_LOC_135/a_8_24# OR2X1_LOC_193/A 0.14fF
C48289 OR2X1_LOC_458/B OR2X1_LOC_723/A 0.02fF
C48290 OR2X1_LOC_9/Y OR2X1_LOC_437/A 0.09fF
C48291 AND2X1_LOC_663/B AND2X1_LOC_624/a_8_24# 0.01fF
C48292 INPUT_1 OR2X1_LOC_32/a_8_216# 0.02fF
C48293 AND2X1_LOC_477/A AND2X1_LOC_645/A 0.07fF
C48294 OR2X1_LOC_11/Y OR2X1_LOC_409/a_36_216# 0.00fF
C48295 OR2X1_LOC_151/A OR2X1_LOC_777/B 0.14fF
C48296 OR2X1_LOC_721/Y OR2X1_LOC_598/A 0.10fF
C48297 OR2X1_LOC_662/a_8_216# AND2X1_LOC_31/Y 0.04fF
C48298 OR2X1_LOC_613/Y AND2X1_LOC_866/A 0.09fF
C48299 OR2X1_LOC_59/Y OR2X1_LOC_526/a_8_216# 0.01fF
C48300 AND2X1_LOC_182/a_36_24# OR2X1_LOC_437/A 0.01fF
C48301 OR2X1_LOC_66/A OR2X1_LOC_71/A 0.08fF
C48302 OR2X1_LOC_45/B AND2X1_LOC_785/A 0.00fF
C48303 AND2X1_LOC_42/a_8_24# INPUT_1 0.06fF
C48304 OR2X1_LOC_89/A AND2X1_LOC_678/a_8_24# 0.05fF
C48305 AND2X1_LOC_784/A AND2X1_LOC_170/B 0.02fF
C48306 OR2X1_LOC_688/a_8_216# D_INPUT_0 0.06fF
C48307 OR2X1_LOC_377/A D_INPUT_1 0.22fF
C48308 OR2X1_LOC_160/B OR2X1_LOC_707/a_8_216# -0.00fF
C48309 OR2X1_LOC_3/Y AND2X1_LOC_196/Y 0.06fF
C48310 OR2X1_LOC_161/B OR2X1_LOC_354/a_8_216# 0.01fF
C48311 AND2X1_LOC_349/a_8_24# OR2X1_LOC_47/Y 0.01fF
C48312 OR2X1_LOC_85/A D_INPUT_1 0.26fF
C48313 AND2X1_LOC_472/B AND2X1_LOC_827/a_8_24# 0.00fF
C48314 OR2X1_LOC_111/Y OR2X1_LOC_74/A 0.09fF
C48315 OR2X1_LOC_36/Y OR2X1_LOC_184/Y 0.03fF
C48316 OR2X1_LOC_22/Y AND2X1_LOC_844/a_8_24# 0.01fF
C48317 OR2X1_LOC_203/Y D_INPUT_1 0.07fF
C48318 AND2X1_LOC_135/a_8_24# D_INPUT_0 0.01fF
C48319 OR2X1_LOC_121/B OR2X1_LOC_606/Y 0.04fF
C48320 OR2X1_LOC_696/A AND2X1_LOC_713/a_8_24# 0.03fF
C48321 AND2X1_LOC_110/Y OR2X1_LOC_469/B 0.03fF
C48322 OR2X1_LOC_62/B OR2X1_LOC_278/A 0.00fF
C48323 OR2X1_LOC_375/A OR2X1_LOC_598/A 0.25fF
C48324 OR2X1_LOC_720/Y OR2X1_LOC_721/a_8_216# 0.39fF
C48325 AND2X1_LOC_313/a_8_24# OR2X1_LOC_308/Y 0.03fF
C48326 OR2X1_LOC_64/Y OR2X1_LOC_417/A 3.41fF
C48327 OR2X1_LOC_256/A AND2X1_LOC_663/B 1.21fF
C48328 OR2X1_LOC_146/Y OR2X1_LOC_74/A 0.03fF
C48329 AND2X1_LOC_773/Y OR2X1_LOC_428/A 0.02fF
C48330 OR2X1_LOC_45/B AND2X1_LOC_219/A 0.42fF
C48331 OR2X1_LOC_448/Y OR2X1_LOC_779/B -0.00fF
C48332 OR2X1_LOC_804/A OR2X1_LOC_155/A 0.03fF
C48333 OR2X1_LOC_76/Y OR2X1_LOC_76/a_8_216# 0.01fF
C48334 OR2X1_LOC_47/Y OR2X1_LOC_83/a_8_216# 0.01fF
C48335 OR2X1_LOC_155/A OR2X1_LOC_512/a_8_216# 0.02fF
C48336 OR2X1_LOC_602/Y OR2X1_LOC_605/Y 0.15fF
C48337 OR2X1_LOC_494/A AND2X1_LOC_363/a_36_24# 0.00fF
C48338 OR2X1_LOC_147/a_8_216# OR2X1_LOC_705/B 0.01fF
C48339 AND2X1_LOC_478/a_8_24# AND2X1_LOC_220/B 0.02fF
C48340 AND2X1_LOC_787/a_8_24# OR2X1_LOC_437/A 0.09fF
C48341 OR2X1_LOC_857/B OR2X1_LOC_857/A 0.14fF
C48342 OR2X1_LOC_405/A OR2X1_LOC_446/B 0.06fF
C48343 OR2X1_LOC_633/A AND2X1_LOC_277/a_36_24# 0.01fF
C48344 OR2X1_LOC_135/a_36_216# OR2X1_LOC_135/Y 0.01fF
C48345 OR2X1_LOC_644/B OR2X1_LOC_228/Y 0.10fF
C48346 AND2X1_LOC_31/Y OR2X1_LOC_719/Y 0.00fF
C48347 AND2X1_LOC_703/Y AND2X1_LOC_714/B 0.01fF
C48348 OR2X1_LOC_19/B AND2X1_LOC_827/a_8_24# 0.02fF
C48349 OR2X1_LOC_121/B OR2X1_LOC_786/Y 0.03fF
C48350 AND2X1_LOC_857/Y OR2X1_LOC_320/a_36_216# 0.00fF
C48351 OR2X1_LOC_433/Y OR2X1_LOC_589/a_8_216# 0.01fF
C48352 OR2X1_LOC_391/B OR2X1_LOC_561/B 0.21fF
C48353 OR2X1_LOC_70/Y OR2X1_LOC_419/Y 3.36fF
C48354 OR2X1_LOC_405/A OR2X1_LOC_728/a_8_216# 0.01fF
C48355 OR2X1_LOC_154/A AND2X1_LOC_419/a_8_24# 0.02fF
C48356 AND2X1_LOC_663/B AND2X1_LOC_624/B 0.00fF
C48357 AND2X1_LOC_663/B OR2X1_LOC_67/Y 0.01fF
C48358 OR2X1_LOC_269/B OR2X1_LOC_724/A 0.07fF
C48359 AND2X1_LOC_822/a_8_24# AND2X1_LOC_31/Y 0.03fF
C48360 OR2X1_LOC_456/a_8_216# D_GATE_366 0.01fF
C48361 AND2X1_LOC_476/Y OR2X1_LOC_322/a_8_216# 0.04fF
C48362 OR2X1_LOC_208/A AND2X1_LOC_41/A 0.03fF
C48363 OR2X1_LOC_175/Y OR2X1_LOC_809/B 0.03fF
C48364 AND2X1_LOC_491/a_8_24# OR2X1_LOC_493/Y 0.02fF
C48365 AND2X1_LOC_243/Y OR2X1_LOC_595/A 0.07fF
C48366 VDD OR2X1_LOC_342/A 0.21fF
C48367 AND2X1_LOC_664/a_8_24# AND2X1_LOC_793/Y 0.01fF
C48368 OR2X1_LOC_45/B AND2X1_LOC_658/A 0.03fF
C48369 OR2X1_LOC_6/B OR2X1_LOC_549/A 0.89fF
C48370 OR2X1_LOC_624/Y OR2X1_LOC_392/B 0.05fF
C48371 INPUT_0 AND2X1_LOC_7/B 0.45fF
C48372 OR2X1_LOC_691/Y OR2X1_LOC_809/B 0.01fF
C48373 OR2X1_LOC_821/Y OR2X1_LOC_813/a_36_216# 0.00fF
C48374 AND2X1_LOC_133/a_36_24# OR2X1_LOC_84/Y 0.01fF
C48375 OR2X1_LOC_199/a_8_216# OR2X1_LOC_78/A 0.04fF
C48376 OR2X1_LOC_750/A OR2X1_LOC_351/a_8_216# 0.02fF
C48377 OR2X1_LOC_134/Y OR2X1_LOC_103/Y 0.10fF
C48378 AND2X1_LOC_22/Y OR2X1_LOC_804/a_8_216# 0.01fF
C48379 OR2X1_LOC_85/A AND2X1_LOC_789/Y 0.01fF
C48380 AND2X1_LOC_565/B AND2X1_LOC_479/a_8_24# 0.20fF
C48381 AND2X1_LOC_550/a_36_24# AND2X1_LOC_476/Y 0.00fF
C48382 OR2X1_LOC_177/Y OR2X1_LOC_59/Y 0.03fF
C48383 AND2X1_LOC_719/Y AND2X1_LOC_285/Y 0.01fF
C48384 OR2X1_LOC_185/A OR2X1_LOC_390/B 0.07fF
C48385 AND2X1_LOC_803/B OR2X1_LOC_40/Y 0.11fF
C48386 OR2X1_LOC_778/Y OR2X1_LOC_723/B 0.16fF
C48387 OR2X1_LOC_56/A OR2X1_LOC_382/a_8_216# 0.03fF
C48388 OR2X1_LOC_294/a_36_216# OR2X1_LOC_161/B 0.00fF
C48389 AND2X1_LOC_392/A VDD 0.49fF
C48390 OR2X1_LOC_846/A OR2X1_LOC_561/B 0.26fF
C48391 OR2X1_LOC_307/B OR2X1_LOC_161/B 0.03fF
C48392 VDD OR2X1_LOC_776/Y 0.00fF
C48393 OR2X1_LOC_78/B OR2X1_LOC_646/B 0.05fF
C48394 OR2X1_LOC_646/A OR2X1_LOC_771/B 0.43fF
C48395 OR2X1_LOC_624/Y OR2X1_LOC_113/B 0.03fF
C48396 AND2X1_LOC_565/B VDD 0.48fF
C48397 VDD AND2X1_LOC_807/B 0.03fF
C48398 OR2X1_LOC_272/Y OR2X1_LOC_13/B 0.03fF
C48399 OR2X1_LOC_240/a_8_216# OR2X1_LOC_415/Y 0.00fF
C48400 OR2X1_LOC_744/A OR2X1_LOC_131/a_8_216# 0.01fF
C48401 AND2X1_LOC_18/Y OR2X1_LOC_244/Y 0.07fF
C48402 AND2X1_LOC_352/a_36_24# OR2X1_LOC_56/A 0.00fF
C48403 OR2X1_LOC_363/B VDD 0.00fF
C48404 AND2X1_LOC_191/B AND2X1_LOC_860/A 0.07fF
C48405 OR2X1_LOC_328/a_8_216# OR2X1_LOC_40/Y 0.00fF
C48406 AND2X1_LOC_53/Y OR2X1_LOC_228/Y 0.03fF
C48407 OR2X1_LOC_482/Y AND2X1_LOC_860/a_8_24# 0.06fF
C48408 OR2X1_LOC_604/A OR2X1_LOC_59/Y 0.50fF
C48409 OR2X1_LOC_92/Y AND2X1_LOC_810/B 0.20fF
C48410 OR2X1_LOC_59/Y AND2X1_LOC_207/B 0.05fF
C48411 OR2X1_LOC_160/A OR2X1_LOC_175/Y 0.46fF
C48412 AND2X1_LOC_7/B OR2X1_LOC_732/B 0.34fF
C48413 AND2X1_LOC_521/a_8_24# OR2X1_LOC_721/Y 0.02fF
C48414 OR2X1_LOC_154/A OR2X1_LOC_115/B 0.01fF
C48415 OR2X1_LOC_161/A AND2X1_LOC_258/a_36_24# 0.00fF
C48416 OR2X1_LOC_490/a_36_216# OR2X1_LOC_92/Y 0.00fF
C48417 AND2X1_LOC_12/Y OR2X1_LOC_352/a_8_216# 0.05fF
C48418 OR2X1_LOC_858/A OR2X1_LOC_66/A 0.15fF
C48419 AND2X1_LOC_841/B AND2X1_LOC_802/Y 0.07fF
C48420 OR2X1_LOC_696/A OR2X1_LOC_6/a_8_216# 0.01fF
C48421 OR2X1_LOC_184/Y OR2X1_LOC_419/Y 0.05fF
C48422 AND2X1_LOC_95/Y AND2X1_LOC_627/a_8_24# 0.02fF
C48423 AND2X1_LOC_53/Y OR2X1_LOC_513/Y 0.00fF
C48424 AND2X1_LOC_571/a_8_24# AND2X1_LOC_573/A 0.01fF
C48425 OR2X1_LOC_516/B AND2X1_LOC_477/Y 0.08fF
C48426 AND2X1_LOC_703/a_8_24# AND2X1_LOC_724/A 0.01fF
C48427 AND2X1_LOC_40/Y OR2X1_LOC_439/B 0.03fF
C48428 AND2X1_LOC_110/Y AND2X1_LOC_167/a_8_24# 0.01fF
C48429 AND2X1_LOC_564/B OR2X1_LOC_406/a_8_216# 0.02fF
C48430 OR2X1_LOC_427/A OR2X1_LOC_603/Y 0.01fF
C48431 VDD AND2X1_LOC_436/a_8_24# -0.00fF
C48432 OR2X1_LOC_692/Y OR2X1_LOC_48/B 0.02fF
C48433 AND2X1_LOC_366/A VDD 0.11fF
C48434 OR2X1_LOC_76/B OR2X1_LOC_736/Y 0.01fF
C48435 AND2X1_LOC_91/B OR2X1_LOC_673/Y 0.12fF
C48436 OR2X1_LOC_160/A OR2X1_LOC_691/Y 0.04fF
C48437 OR2X1_LOC_151/A OR2X1_LOC_575/A 0.01fF
C48438 OR2X1_LOC_8/Y OR2X1_LOC_235/B 1.03fF
C48439 OR2X1_LOC_756/B VDD 2.38fF
C48440 AND2X1_LOC_59/Y AND2X1_LOC_44/Y 4.63fF
C48441 OR2X1_LOC_692/Y OR2X1_LOC_18/Y 0.01fF
C48442 OR2X1_LOC_426/B AND2X1_LOC_474/A 0.07fF
C48443 OR2X1_LOC_47/Y OR2X1_LOC_754/Y 0.01fF
C48444 AND2X1_LOC_541/a_8_24# AND2X1_LOC_560/B 0.01fF
C48445 OR2X1_LOC_223/A OR2X1_LOC_228/Y 0.01fF
C48446 AND2X1_LOC_340/Y OR2X1_LOC_65/B 0.25fF
C48447 AND2X1_LOC_391/Y OR2X1_LOC_744/A 0.04fF
C48448 AND2X1_LOC_621/Y AND2X1_LOC_212/Y 0.07fF
C48449 OR2X1_LOC_744/A AND2X1_LOC_858/B 0.14fF
C48450 AND2X1_LOC_432/a_36_24# OR2X1_LOC_130/A 0.01fF
C48451 OR2X1_LOC_840/a_8_216# OR2X1_LOC_185/A 0.01fF
C48452 OR2X1_LOC_744/A OR2X1_LOC_91/A 0.14fF
C48453 AND2X1_LOC_738/B OR2X1_LOC_677/a_8_216# 0.04fF
C48454 AND2X1_LOC_658/B AND2X1_LOC_185/a_8_24# 0.19fF
C48455 AND2X1_LOC_847/Y OR2X1_LOC_382/A 0.02fF
C48456 OR2X1_LOC_147/B AND2X1_LOC_18/Y 0.03fF
C48457 AND2X1_LOC_801/B OR2X1_LOC_13/B 0.02fF
C48458 OR2X1_LOC_579/B OR2X1_LOC_843/B 0.04fF
C48459 AND2X1_LOC_521/a_8_24# OR2X1_LOC_375/A 0.08fF
C48460 OR2X1_LOC_715/B OR2X1_LOC_624/A 0.11fF
C48461 AND2X1_LOC_721/a_8_24# OR2X1_LOC_51/Y 0.01fF
C48462 OR2X1_LOC_707/B OR2X1_LOC_712/B 0.01fF
C48463 OR2X1_LOC_121/B OR2X1_LOC_301/a_36_216# 0.00fF
C48464 AND2X1_LOC_42/B OR2X1_LOC_120/a_8_216# 0.04fF
C48465 AND2X1_LOC_357/A OR2X1_LOC_619/Y 0.04fF
C48466 OR2X1_LOC_84/a_8_216# OR2X1_LOC_80/A 0.01fF
C48467 OR2X1_LOC_600/A OR2X1_LOC_48/B 0.07fF
C48468 AND2X1_LOC_517/a_8_24# AND2X1_LOC_18/Y 0.02fF
C48469 AND2X1_LOC_6/a_36_24# OR2X1_LOC_68/B 0.01fF
C48470 OR2X1_LOC_494/A OR2X1_LOC_485/A 0.00fF
C48471 AND2X1_LOC_59/Y OR2X1_LOC_719/a_8_216# 0.01fF
C48472 OR2X1_LOC_326/B OR2X1_LOC_325/Y 0.06fF
C48473 AND2X1_LOC_775/a_8_24# OR2X1_LOC_177/Y 0.01fF
C48474 OR2X1_LOC_653/B OR2X1_LOC_364/A 0.06fF
C48475 OR2X1_LOC_84/A OR2X1_LOC_71/A 0.02fF
C48476 AND2X1_LOC_555/Y OR2X1_LOC_481/A 0.02fF
C48477 AND2X1_LOC_22/Y OR2X1_LOC_574/A 0.03fF
C48478 VDD AND2X1_LOC_354/Y 0.21fF
C48479 OR2X1_LOC_769/B OR2X1_LOC_637/A 0.16fF
C48480 AND2X1_LOC_724/a_8_24# OR2X1_LOC_485/A 0.02fF
C48481 OR2X1_LOC_600/A OR2X1_LOC_18/Y 0.23fF
C48482 OR2X1_LOC_91/Y AND2X1_LOC_719/Y 0.06fF
C48483 OR2X1_LOC_585/A OR2X1_LOC_414/Y 0.03fF
C48484 OR2X1_LOC_74/A AND2X1_LOC_804/A 0.02fF
C48485 OR2X1_LOC_158/A OR2X1_LOC_699/a_8_216# 0.02fF
C48486 AND2X1_LOC_7/Y AND2X1_LOC_36/Y 0.01fF
C48487 AND2X1_LOC_40/Y AND2X1_LOC_41/A 0.87fF
C48488 OR2X1_LOC_186/Y AND2X1_LOC_329/a_8_24# 0.01fF
C48489 OR2X1_LOC_7/A AND2X1_LOC_774/A 0.07fF
C48490 AND2X1_LOC_573/a_8_24# AND2X1_LOC_657/Y 0.20fF
C48491 OR2X1_LOC_743/A OR2X1_LOC_744/Y 0.01fF
C48492 AND2X1_LOC_3/Y OR2X1_LOC_580/B 1.71fF
C48493 AND2X1_LOC_553/A OR2X1_LOC_179/a_8_216# 0.47fF
C48494 AND2X1_LOC_669/a_8_24# AND2X1_LOC_18/Y 0.02fF
C48495 AND2X1_LOC_682/a_8_24# OR2X1_LOC_78/B 0.02fF
C48496 OR2X1_LOC_40/Y OR2X1_LOC_613/Y 0.00fF
C48497 OR2X1_LOC_711/B OR2X1_LOC_469/a_36_216# 0.00fF
C48498 OR2X1_LOC_49/A AND2X1_LOC_42/B 0.38fF
C48499 OR2X1_LOC_160/A OR2X1_LOC_803/A 0.03fF
C48500 AND2X1_LOC_737/Y AND2X1_LOC_734/Y 0.07fF
C48501 AND2X1_LOC_59/Y OR2X1_LOC_785/a_8_216# 0.01fF
C48502 OR2X1_LOC_9/Y OR2X1_LOC_753/A 0.03fF
C48503 AND2X1_LOC_78/a_8_24# OR2X1_LOC_16/A 0.10fF
C48504 OR2X1_LOC_252/a_8_216# OR2X1_LOC_59/Y 0.01fF
C48505 OR2X1_LOC_648/A OR2X1_LOC_405/Y 0.02fF
C48506 OR2X1_LOC_506/A OR2X1_LOC_78/B 0.03fF
C48507 VDD OR2X1_LOC_657/a_8_216# 0.00fF
C48508 OR2X1_LOC_744/A AND2X1_LOC_573/A 0.48fF
C48509 AND2X1_LOC_539/Y AND2X1_LOC_727/A 0.01fF
C48510 OR2X1_LOC_551/B OR2X1_LOC_367/B 0.20fF
C48511 AND2X1_LOC_477/Y AND2X1_LOC_220/Y 0.21fF
C48512 AND2X1_LOC_81/a_8_24# OR2X1_LOC_786/A 0.01fF
C48513 AND2X1_LOC_12/Y AND2X1_LOC_628/a_8_24# 0.02fF
C48514 OR2X1_LOC_593/a_8_216# OR2X1_LOC_66/A 0.01fF
C48515 OR2X1_LOC_604/A OR2X1_LOC_820/B 0.01fF
C48516 INPUT_0 OR2X1_LOC_407/a_8_216# 0.03fF
C48517 AND2X1_LOC_723/Y AND2X1_LOC_168/Y 0.00fF
C48518 OR2X1_LOC_426/B OR2X1_LOC_85/A 0.02fF
C48519 OR2X1_LOC_275/A OR2X1_LOC_16/A 0.08fF
C48520 OR2X1_LOC_840/A OR2X1_LOC_620/Y 0.10fF
C48521 OR2X1_LOC_130/A OR2X1_LOC_78/A 0.12fF
C48522 VDD OR2X1_LOC_76/Y 0.13fF
C48523 AND2X1_LOC_755/a_8_24# OR2X1_LOC_756/B 0.02fF
C48524 OR2X1_LOC_537/A AND2X1_LOC_41/A 0.03fF
C48525 OR2X1_LOC_648/B AND2X1_LOC_3/Y 0.01fF
C48526 OR2X1_LOC_177/Y OR2X1_LOC_70/Y 0.04fF
C48527 OR2X1_LOC_46/A AND2X1_LOC_202/Y 0.04fF
C48528 OR2X1_LOC_6/B OR2X1_LOC_401/Y 0.06fF
C48529 OR2X1_LOC_604/A AND2X1_LOC_446/a_36_24# 0.00fF
C48530 OR2X1_LOC_518/Y OR2X1_LOC_31/Y 0.27fF
C48531 OR2X1_LOC_80/Y OR2X1_LOC_59/Y 0.80fF
C48532 AND2X1_LOC_580/A AND2X1_LOC_663/A 0.03fF
C48533 OR2X1_LOC_467/A OR2X1_LOC_449/B 1.26fF
C48534 AND2X1_LOC_851/A OR2X1_LOC_427/A 0.04fF
C48535 AND2X1_LOC_717/B AND2X1_LOC_489/a_8_24# 0.03fF
C48536 OR2X1_LOC_421/A OR2X1_LOC_3/Y 0.01fF
C48537 OR2X1_LOC_26/Y AND2X1_LOC_434/Y 0.02fF
C48538 OR2X1_LOC_427/A AND2X1_LOC_808/a_8_24# 0.02fF
C48539 OR2X1_LOC_26/Y AND2X1_LOC_219/Y 0.01fF
C48540 OR2X1_LOC_619/Y AND2X1_LOC_852/B 0.01fF
C48541 OR2X1_LOC_599/A OR2X1_LOC_524/Y 0.34fF
C48542 OR2X1_LOC_604/A AND2X1_LOC_711/Y 0.11fF
C48543 OR2X1_LOC_856/A OR2X1_LOC_19/B 0.07fF
C48544 OR2X1_LOC_471/Y OR2X1_LOC_547/a_8_216# 0.06fF
C48545 OR2X1_LOC_604/A OR2X1_LOC_70/Y 0.22fF
C48546 AND2X1_LOC_568/B AND2X1_LOC_211/a_8_24# 0.01fF
C48547 AND2X1_LOC_32/a_36_24# OR2X1_LOC_334/B 0.00fF
C48548 OR2X1_LOC_482/Y AND2X1_LOC_842/B 0.03fF
C48549 OR2X1_LOC_154/A OR2X1_LOC_840/A 0.17fF
C48550 OR2X1_LOC_619/Y OR2X1_LOC_48/B 0.14fF
C48551 OR2X1_LOC_364/A OR2X1_LOC_808/B 0.22fF
C48552 AND2X1_LOC_366/A OR2X1_LOC_251/Y 0.03fF
C48553 OR2X1_LOC_602/Y OR2X1_LOC_602/a_8_216# 0.01fF
C48554 OR2X1_LOC_18/Y OR2X1_LOC_619/Y 0.03fF
C48555 AND2X1_LOC_681/a_36_24# AND2X1_LOC_3/Y 0.00fF
C48556 AND2X1_LOC_95/Y OR2X1_LOC_377/A 0.22fF
C48557 AND2X1_LOC_81/B OR2X1_LOC_509/A 0.01fF
C48558 AND2X1_LOC_753/B AND2X1_LOC_56/B 0.02fF
C48559 OR2X1_LOC_377/A OR2X1_LOC_633/Y 0.12fF
C48560 AND2X1_LOC_40/Y OR2X1_LOC_631/B 0.42fF
C48561 AND2X1_LOC_323/a_8_24# OR2X1_LOC_121/B 0.01fF
C48562 AND2X1_LOC_496/a_8_24# AND2X1_LOC_628/a_8_24# 0.23fF
C48563 OR2X1_LOC_604/A AND2X1_LOC_514/Y 0.10fF
C48564 AND2X1_LOC_95/Y AND2X1_LOC_824/B 0.04fF
C48565 OR2X1_LOC_506/A OR2X1_LOC_375/A 0.00fF
C48566 AND2X1_LOC_866/A AND2X1_LOC_786/Y 0.07fF
C48567 OR2X1_LOC_421/a_8_216# OR2X1_LOC_743/A 0.01fF
C48568 OR2X1_LOC_862/a_8_216# D_INPUT_1 0.02fF
C48569 OR2X1_LOC_92/Y OR2X1_LOC_585/A 0.14fF
C48570 OR2X1_LOC_467/A OR2X1_LOC_121/B 0.00fF
C48571 AND2X1_LOC_348/a_36_24# OR2X1_LOC_91/A 0.01fF
C48572 AND2X1_LOC_47/Y OR2X1_LOC_549/A 1.31fF
C48573 OR2X1_LOC_405/A AND2X1_LOC_56/B 0.01fF
C48574 AND2X1_LOC_99/A OR2X1_LOC_44/Y 0.01fF
C48575 OR2X1_LOC_429/Y OR2X1_LOC_425/a_8_216# 0.05fF
C48576 AND2X1_LOC_95/Y OR2X1_LOC_203/Y 0.14fF
C48577 OR2X1_LOC_318/Y OR2X1_LOC_592/a_36_216# 0.02fF
C48578 AND2X1_LOC_578/A AND2X1_LOC_722/A 0.10fF
C48579 AND2X1_LOC_703/a_8_24# OR2X1_LOC_312/Y 0.11fF
C48580 OR2X1_LOC_270/Y OR2X1_LOC_580/B 0.01fF
C48581 OR2X1_LOC_520/Y OR2X1_LOC_462/B 0.01fF
C48582 OR2X1_LOC_377/A OR2X1_LOC_99/Y 0.04fF
C48583 OR2X1_LOC_497/Y OR2X1_LOC_39/A 0.04fF
C48584 AND2X1_LOC_159/a_8_24# OR2X1_LOC_161/A 0.01fF
C48585 OR2X1_LOC_485/A OR2X1_LOC_427/A 14.75fF
C48586 OR2X1_LOC_62/B OR2X1_LOC_78/A 0.05fF
C48587 OR2X1_LOC_810/A OR2X1_LOC_161/A 0.03fF
C48588 OR2X1_LOC_307/a_8_216# OR2X1_LOC_161/A 0.03fF
C48589 OR2X1_LOC_777/B OR2X1_LOC_716/a_8_216# 0.05fF
C48590 OR2X1_LOC_13/B OR2X1_LOC_248/A 0.01fF
C48591 OR2X1_LOC_648/A D_INPUT_0 0.52fF
C48592 OR2X1_LOC_670/a_8_216# OR2X1_LOC_6/A 0.01fF
C48593 OR2X1_LOC_276/B OR2X1_LOC_629/B 0.01fF
C48594 OR2X1_LOC_261/Y AND2X1_LOC_847/Y 0.02fF
C48595 OR2X1_LOC_707/A OR2X1_LOC_155/A 0.01fF
C48596 OR2X1_LOC_485/A OR2X1_LOC_63/a_8_216# 0.01fF
C48597 OR2X1_LOC_115/B OR2X1_LOC_560/A 0.02fF
C48598 AND2X1_LOC_126/a_8_24# OR2X1_LOC_19/B 0.00fF
C48599 AND2X1_LOC_36/Y OR2X1_LOC_515/a_8_216# 0.01fF
C48600 OR2X1_LOC_43/A OR2X1_LOC_236/a_36_216# 0.01fF
C48601 OR2X1_LOC_561/a_8_216# OR2X1_LOC_269/B -0.00fF
C48602 AND2X1_LOC_319/A OR2X1_LOC_52/B 0.07fF
C48603 AND2X1_LOC_158/a_8_24# OR2X1_LOC_87/A 0.03fF
C48604 AND2X1_LOC_784/A AND2X1_LOC_170/Y 0.02fF
C48605 AND2X1_LOC_637/Y OR2X1_LOC_44/Y 0.02fF
C48606 OR2X1_LOC_780/B OR2X1_LOC_78/A 0.02fF
C48607 OR2X1_LOC_18/Y OR2X1_LOC_372/a_8_216# 0.00fF
C48608 OR2X1_LOC_716/a_36_216# OR2X1_LOC_593/B 0.00fF
C48609 OR2X1_LOC_851/A OR2X1_LOC_121/B 0.01fF
C48610 AND2X1_LOC_108/a_36_24# OR2X1_LOC_78/A 0.00fF
C48611 OR2X1_LOC_343/a_8_216# OR2X1_LOC_493/Y 0.29fF
C48612 AND2X1_LOC_852/Y OR2X1_LOC_753/A 0.07fF
C48613 AND2X1_LOC_12/Y AND2X1_LOC_69/Y 0.01fF
C48614 AND2X1_LOC_858/B OR2X1_LOC_31/Y 0.03fF
C48615 AND2X1_LOC_553/a_36_24# OR2X1_LOC_47/Y 0.00fF
C48616 OR2X1_LOC_113/Y AND2X1_LOC_47/Y 0.52fF
C48617 AND2X1_LOC_42/B OR2X1_LOC_575/a_8_216# 0.01fF
C48618 OR2X1_LOC_420/a_8_216# OR2X1_LOC_591/A 0.47fF
C48619 OR2X1_LOC_91/A OR2X1_LOC_31/Y 0.60fF
C48620 OR2X1_LOC_502/A AND2X1_LOC_165/a_8_24# 0.05fF
C48621 OR2X1_LOC_521/Y AND2X1_LOC_115/a_8_24# 0.00fF
C48622 AND2X1_LOC_665/a_36_24# OR2X1_LOC_78/A 0.00fF
C48623 OR2X1_LOC_598/A OR2X1_LOC_549/A 1.50fF
C48624 OR2X1_LOC_600/A AND2X1_LOC_620/Y 0.03fF
C48625 OR2X1_LOC_837/A OR2X1_LOC_46/A 0.51fF
C48626 OR2X1_LOC_95/Y AND2X1_LOC_471/Y 1.18fF
C48627 AND2X1_LOC_554/B OR2X1_LOC_6/A 0.03fF
C48628 OR2X1_LOC_596/Y AND2X1_LOC_387/B 0.00fF
C48629 AND2X1_LOC_784/Y AND2X1_LOC_804/a_8_24# 0.20fF
C48630 AND2X1_LOC_440/a_8_24# AND2X1_LOC_471/Y 0.20fF
C48631 OR2X1_LOC_223/A OR2X1_LOC_191/a_8_216# 0.01fF
C48632 AND2X1_LOC_229/a_8_24# AND2X1_LOC_31/Y 0.01fF
C48633 AND2X1_LOC_1/Y OR2X1_LOC_639/B 0.09fF
C48634 AND2X1_LOC_42/B OR2X1_LOC_87/B 0.10fF
C48635 OR2X1_LOC_510/Y AND2X1_LOC_51/Y 0.03fF
C48636 OR2X1_LOC_78/B OR2X1_LOC_227/Y 0.00fF
C48637 OR2X1_LOC_417/Y OR2X1_LOC_313/Y 0.10fF
C48638 OR2X1_LOC_51/Y AND2X1_LOC_770/a_36_24# 0.00fF
C48639 OR2X1_LOC_8/Y AND2X1_LOC_721/A 0.02fF
C48640 OR2X1_LOC_485/A AND2X1_LOC_363/A 0.01fF
C48641 AND2X1_LOC_662/B OR2X1_LOC_268/a_8_216# 0.03fF
C48642 OR2X1_LOC_114/B OR2X1_LOC_247/Y 0.00fF
C48643 AND2X1_LOC_250/a_8_24# OR2X1_LOC_561/Y 0.05fF
C48644 OR2X1_LOC_185/A OR2X1_LOC_649/a_8_216# 0.01fF
C48645 OR2X1_LOC_78/B D_INPUT_1 0.10fF
C48646 OR2X1_LOC_311/Y AND2X1_LOC_655/A 0.05fF
C48647 AND2X1_LOC_326/A OR2X1_LOC_6/A 0.00fF
C48648 AND2X1_LOC_34/Y OR2X1_LOC_46/A 0.02fF
C48649 OR2X1_LOC_52/a_8_216# OR2X1_LOC_52/B 0.07fF
C48650 AND2X1_LOC_490/a_36_24# AND2X1_LOC_3/Y 0.00fF
C48651 AND2X1_LOC_85/a_8_24# AND2X1_LOC_42/B 0.01fF
C48652 OR2X1_LOC_773/B OR2X1_LOC_773/a_8_216# 0.06fF
C48653 OR2X1_LOC_285/B OR2X1_LOC_269/B 0.00fF
C48654 AND2X1_LOC_787/A OR2X1_LOC_437/A 0.58fF
C48655 AND2X1_LOC_555/Y AND2X1_LOC_789/Y 0.08fF
C48656 AND2X1_LOC_663/B OR2X1_LOC_248/Y 0.29fF
C48657 OR2X1_LOC_476/B OR2X1_LOC_87/A 0.05fF
C48658 AND2X1_LOC_840/A OR2X1_LOC_95/Y 0.03fF
C48659 AND2X1_LOC_330/a_36_24# OR2X1_LOC_419/Y 0.06fF
C48660 AND2X1_LOC_3/Y AND2X1_LOC_425/a_8_24# 0.20fF
C48661 OR2X1_LOC_246/A OR2X1_LOC_85/A 0.09fF
C48662 OR2X1_LOC_810/A AND2X1_LOC_51/Y 1.76fF
C48663 AND2X1_LOC_101/B OR2X1_LOC_64/Y 0.25fF
C48664 OR2X1_LOC_787/a_8_216# OR2X1_LOC_578/B 0.02fF
C48665 OR2X1_LOC_641/A OR2X1_LOC_68/B 0.03fF
C48666 OR2X1_LOC_78/A OR2X1_LOC_365/B 0.03fF
C48667 AND2X1_LOC_193/a_8_24# OR2X1_LOC_7/Y 0.09fF
C48668 OR2X1_LOC_97/A OR2X1_LOC_544/B 0.29fF
C48669 OR2X1_LOC_158/A OR2X1_LOC_521/a_8_216# 0.04fF
C48670 AND2X1_LOC_708/a_8_24# OR2X1_LOC_52/B 0.03fF
C48671 AND2X1_LOC_100/a_8_24# OR2X1_LOC_19/B 0.02fF
C48672 OR2X1_LOC_427/A AND2X1_LOC_452/a_8_24# 0.01fF
C48673 AND2X1_LOC_31/Y OR2X1_LOC_66/A 1.84fF
C48674 OR2X1_LOC_46/A OR2X1_LOC_49/a_8_216# 0.03fF
C48675 OR2X1_LOC_291/Y OR2X1_LOC_609/A 0.04fF
C48676 OR2X1_LOC_841/A AND2X1_LOC_31/Y 0.07fF
C48677 OR2X1_LOC_22/Y OR2X1_LOC_24/a_8_216# 0.05fF
C48678 AND2X1_LOC_347/a_8_24# AND2X1_LOC_663/B 0.01fF
C48679 AND2X1_LOC_658/B OR2X1_LOC_152/A 0.06fF
C48680 OR2X1_LOC_6/B OR2X1_LOC_399/a_8_216# 0.01fF
C48681 AND2X1_LOC_12/Y OR2X1_LOC_506/B 0.05fF
C48682 OR2X1_LOC_62/a_8_216# OR2X1_LOC_585/A 0.01fF
C48683 OR2X1_LOC_774/Y OR2X1_LOC_859/A 0.05fF
C48684 AND2X1_LOC_566/B OR2X1_LOC_437/A 0.00fF
C48685 OR2X1_LOC_151/A OR2X1_LOC_735/B 0.07fF
C48686 AND2X1_LOC_311/a_8_24# AND2X1_LOC_31/Y 0.01fF
C48687 AND2X1_LOC_624/A OR2X1_LOC_615/Y 0.03fF
C48688 VDD AND2X1_LOC_738/Y 0.25fF
C48689 VDD OR2X1_LOC_589/Y 0.26fF
C48690 OR2X1_LOC_436/Y OR2X1_LOC_809/a_36_216# 0.00fF
C48691 OR2X1_LOC_780/B OR2X1_LOC_155/A 0.50fF
C48692 AND2X1_LOC_260/a_8_24# OR2X1_LOC_54/Y 0.02fF
C48693 AND2X1_LOC_738/a_8_24# AND2X1_LOC_738/Y 0.00fF
C48694 AND2X1_LOC_731/Y AND2X1_LOC_742/A 0.23fF
C48695 OR2X1_LOC_557/A AND2X1_LOC_15/a_8_24# 0.01fF
C48696 OR2X1_LOC_43/A OR2X1_LOC_96/a_8_216# 0.03fF
C48697 OR2X1_LOC_696/A AND2X1_LOC_457/a_8_24# 0.01fF
C48698 OR2X1_LOC_375/A D_INPUT_1 0.10fF
C48699 AND2X1_LOC_96/a_8_24# OR2X1_LOC_80/A 0.02fF
C48700 AND2X1_LOC_851/B OR2X1_LOC_26/Y 0.09fF
C48701 OR2X1_LOC_502/A OR2X1_LOC_228/Y 0.07fF
C48702 OR2X1_LOC_36/Y OR2X1_LOC_47/Y 0.22fF
C48703 AND2X1_LOC_572/a_36_24# OR2X1_LOC_106/Y 0.01fF
C48704 OR2X1_LOC_252/Y AND2X1_LOC_483/Y 0.18fF
C48705 OR2X1_LOC_619/Y AND2X1_LOC_215/A 0.03fF
C48706 OR2X1_LOC_602/a_8_216# OR2X1_LOC_602/B 0.05fF
C48707 OR2X1_LOC_249/Y OR2X1_LOC_493/Y 0.50fF
C48708 AND2X1_LOC_810/a_8_24# OR2X1_LOC_44/Y 0.06fF
C48709 OR2X1_LOC_808/B OR2X1_LOC_578/B 0.05fF
C48710 OR2X1_LOC_108/Y OR2X1_LOC_142/Y 0.14fF
C48711 AND2X1_LOC_537/Y AND2X1_LOC_358/a_8_24# 0.11fF
C48712 AND2X1_LOC_8/Y AND2X1_LOC_8/a_8_24# 0.01fF
C48713 AND2X1_LOC_56/B OR2X1_LOC_330/a_8_216# 0.02fF
C48714 OR2X1_LOC_625/Y OR2X1_LOC_754/Y 0.07fF
C48715 AND2X1_LOC_817/B OR2X1_LOC_774/B 0.16fF
C48716 AND2X1_LOC_22/Y OR2X1_LOC_855/A 0.01fF
C48717 OR2X1_LOC_64/Y OR2X1_LOC_226/a_8_216# 0.01fF
C48718 OR2X1_LOC_139/A OR2X1_LOC_572/a_8_216# 0.02fF
C48719 OR2X1_LOC_476/B OR2X1_LOC_648/a_8_216# 0.06fF
C48720 AND2X1_LOC_43/B AND2X1_LOC_52/Y 0.05fF
C48721 OR2X1_LOC_241/Y OR2X1_LOC_778/A 0.04fF
C48722 OR2X1_LOC_316/Y AND2X1_LOC_222/Y 0.00fF
C48723 OR2X1_LOC_155/A AND2X1_LOC_39/Y 0.07fF
C48724 AND2X1_LOC_363/B OR2X1_LOC_384/Y 0.02fF
C48725 OR2X1_LOC_43/A OR2X1_LOC_311/a_8_216# 0.04fF
C48726 AND2X1_LOC_778/a_8_24# AND2X1_LOC_795/Y 0.01fF
C48727 AND2X1_LOC_300/a_8_24# OR2X1_LOC_831/B 0.20fF
C48728 OR2X1_LOC_56/A OR2X1_LOC_268/Y 0.03fF
C48729 OR2X1_LOC_106/Y OR2X1_LOC_158/A 0.03fF
C48730 AND2X1_LOC_69/a_8_24# OR2X1_LOC_814/A 0.01fF
C48731 OR2X1_LOC_87/A OR2X1_LOC_590/a_36_216# 0.00fF
C48732 AND2X1_LOC_423/a_36_24# OR2X1_LOC_446/B 0.00fF
C48733 OR2X1_LOC_56/A OR2X1_LOC_183/Y 0.13fF
C48734 OR2X1_LOC_91/A OR2X1_LOC_320/a_8_216# 0.02fF
C48735 OR2X1_LOC_12/Y OR2X1_LOC_428/A 1.11fF
C48736 AND2X1_LOC_663/B AND2X1_LOC_660/A 0.07fF
C48737 AND2X1_LOC_191/Y OR2X1_LOC_747/a_8_216# 0.03fF
C48738 OR2X1_LOC_269/B OR2X1_LOC_358/A 0.02fF
C48739 OR2X1_LOC_160/A OR2X1_LOC_546/A 0.16fF
C48740 VDD OR2X1_LOC_140/B 0.19fF
C48741 OR2X1_LOC_76/A OR2X1_LOC_223/A 0.00fF
C48742 OR2X1_LOC_468/Y OR2X1_LOC_567/a_36_216# 0.00fF
C48743 OR2X1_LOC_182/B OR2X1_LOC_352/a_8_216# 0.01fF
C48744 OR2X1_LOC_417/A OR2X1_LOC_226/a_8_216# 0.06fF
C48745 OR2X1_LOC_12/Y OR2X1_LOC_595/A 0.07fF
C48746 OR2X1_LOC_548/A OR2X1_LOC_548/a_8_216# 0.47fF
C48747 OR2X1_LOC_151/A OR2X1_LOC_161/B 0.24fF
C48748 OR2X1_LOC_651/a_8_216# AND2X1_LOC_31/Y 0.07fF
C48749 AND2X1_LOC_351/Y OR2X1_LOC_289/a_8_216# 0.07fF
C48750 OR2X1_LOC_629/a_8_216# OR2X1_LOC_598/A 0.04fF
C48751 OR2X1_LOC_128/B OR2X1_LOC_342/a_8_216# 0.47fF
C48752 AND2X1_LOC_227/Y AND2X1_LOC_656/Y 0.03fF
C48753 OR2X1_LOC_136/Y OR2X1_LOC_426/B 0.16fF
C48754 OR2X1_LOC_696/A OR2X1_LOC_382/Y 0.02fF
C48755 OR2X1_LOC_710/A AND2X1_LOC_41/A 0.01fF
C48756 OR2X1_LOC_311/Y OR2X1_LOC_599/Y 0.03fF
C48757 OR2X1_LOC_231/B AND2X1_LOC_18/Y 0.03fF
C48758 OR2X1_LOC_482/a_8_216# OR2X1_LOC_482/Y 0.01fF
C48759 OR2X1_LOC_203/Y OR2X1_LOC_269/A 1.27fF
C48760 AND2X1_LOC_95/Y OR2X1_LOC_539/B 0.02fF
C48761 OR2X1_LOC_179/a_8_216# AND2X1_LOC_465/A 0.01fF
C48762 OR2X1_LOC_804/A OR2X1_LOC_814/A 0.06fF
C48763 OR2X1_LOC_201/Y OR2X1_LOC_68/B 0.01fF
C48764 AND2X1_LOC_181/Y OR2X1_LOC_600/A 0.01fF
C48765 OR2X1_LOC_106/Y OR2X1_LOC_103/Y 0.03fF
C48766 OR2X1_LOC_294/a_8_216# OR2X1_LOC_563/A 0.01fF
C48767 AND2X1_LOC_738/B AND2X1_LOC_705/Y 0.10fF
C48768 OR2X1_LOC_865/A OR2X1_LOC_391/A 0.17fF
C48769 OR2X1_LOC_533/Y OR2X1_LOC_59/Y 0.01fF
C48770 AND2X1_LOC_447/Y OR2X1_LOC_421/Y 0.03fF
C48771 OR2X1_LOC_40/Y AND2X1_LOC_499/a_36_24# 0.00fF
C48772 AND2X1_LOC_360/a_8_24# OR2X1_LOC_494/A 0.01fF
C48773 AND2X1_LOC_566/B AND2X1_LOC_715/A 0.03fF
C48774 OR2X1_LOC_156/A OR2X1_LOC_160/B 0.22fF
C48775 AND2X1_LOC_91/B AND2X1_LOC_384/a_8_24# 0.09fF
C48776 AND2X1_LOC_212/Y OR2X1_LOC_59/Y 0.07fF
C48777 OR2X1_LOC_158/A AND2X1_LOC_658/A 0.03fF
C48778 OR2X1_LOC_359/a_8_216# OR2X1_LOC_362/A 0.01fF
C48779 OR2X1_LOC_53/Y AND2X1_LOC_654/B 0.07fF
C48780 OR2X1_LOC_158/A OR2X1_LOC_690/Y 0.03fF
C48781 AND2X1_LOC_77/a_36_24# OR2X1_LOC_68/B 0.00fF
C48782 OR2X1_LOC_114/B AND2X1_LOC_18/Y 0.03fF
C48783 AND2X1_LOC_48/A OR2X1_LOC_228/Y 0.17fF
C48784 AND2X1_LOC_64/Y OR2X1_LOC_661/a_8_216# 0.05fF
C48785 OR2X1_LOC_264/Y OR2X1_LOC_139/A 0.00fF
C48786 OR2X1_LOC_139/A OR2X1_LOC_436/B 0.01fF
C48787 AND2X1_LOC_22/Y AND2X1_LOC_58/a_8_24# 0.03fF
C48788 AND2X1_LOC_658/B OR2X1_LOC_604/A 0.07fF
C48789 AND2X1_LOC_658/B OR2X1_LOC_745/a_8_216# 0.05fF
C48790 AND2X1_LOC_70/Y OR2X1_LOC_629/B 0.01fF
C48791 AND2X1_LOC_91/B OR2X1_LOC_812/B 0.02fF
C48792 OR2X1_LOC_422/a_8_216# OR2X1_LOC_428/A 0.01fF
C48793 OR2X1_LOC_811/A OR2X1_LOC_563/A 0.07fF
C48794 OR2X1_LOC_623/B AND2X1_LOC_44/Y 0.03fF
C48795 AND2X1_LOC_544/Y AND2X1_LOC_550/A 0.01fF
C48796 AND2X1_LOC_48/A OR2X1_LOC_513/Y 0.01fF
C48797 OR2X1_LOC_477/Y OR2X1_LOC_161/B 0.56fF
C48798 OR2X1_LOC_188/Y OR2X1_LOC_465/Y 0.02fF
C48799 OR2X1_LOC_16/A OR2X1_LOC_16/a_8_216# 0.18fF
C48800 OR2X1_LOC_161/A AND2X1_LOC_760/a_36_24# 0.01fF
C48801 OR2X1_LOC_683/a_8_216# OR2X1_LOC_16/A 0.05fF
C48802 OR2X1_LOC_22/Y AND2X1_LOC_215/a_8_24# 0.03fF
C48803 OR2X1_LOC_696/A OR2X1_LOC_591/A 0.07fF
C48804 AND2X1_LOC_716/Y OR2X1_LOC_135/Y 0.10fF
C48805 OR2X1_LOC_421/A OR2X1_LOC_329/B 0.01fF
C48806 OR2X1_LOC_788/a_8_216# OR2X1_LOC_161/B 0.01fF
C48807 AND2X1_LOC_541/Y AND2X1_LOC_367/A 0.02fF
C48808 OR2X1_LOC_6/B AND2X1_LOC_498/a_36_24# -0.02fF
C48809 OR2X1_LOC_48/B AND2X1_LOC_769/Y 0.03fF
C48810 OR2X1_LOC_47/Y OR2X1_LOC_419/Y 0.03fF
C48811 OR2X1_LOC_426/B OR2X1_LOC_51/Y 0.02fF
C48812 OR2X1_LOC_40/Y OR2X1_LOC_524/Y 5.32fF
C48813 AND2X1_LOC_64/Y OR2X1_LOC_462/B 0.14fF
C48814 OR2X1_LOC_326/a_36_216# AND2X1_LOC_110/Y 0.00fF
C48815 AND2X1_LOC_64/Y OR2X1_LOC_483/a_8_216# 0.01fF
C48816 AND2X1_LOC_22/Y OR2X1_LOC_377/A 0.07fF
C48817 OR2X1_LOC_468/A OR2X1_LOC_78/A 0.02fF
C48818 OR2X1_LOC_18/Y AND2X1_LOC_769/Y 0.01fF
C48819 OR2X1_LOC_694/Y OR2X1_LOC_91/A 0.04fF
C48820 OR2X1_LOC_185/Y OR2X1_LOC_120/a_8_216# 0.03fF
C48821 OR2X1_LOC_6/B OR2X1_LOC_499/B 0.07fF
C48822 OR2X1_LOC_805/A AND2X1_LOC_7/B 0.25fF
C48823 OR2X1_LOC_135/Y AND2X1_LOC_654/Y 0.10fF
C48824 AND2X1_LOC_40/Y AND2X1_LOC_83/a_36_24# 0.00fF
C48825 AND2X1_LOC_482/a_8_24# OR2X1_LOC_344/A 0.01fF
C48826 OR2X1_LOC_833/B AND2X1_LOC_256/a_8_24# 0.02fF
C48827 AND2X1_LOC_523/a_8_24# OR2X1_LOC_522/Y 0.01fF
C48828 OR2X1_LOC_151/A OR2X1_LOC_61/Y 0.07fF
C48829 OR2X1_LOC_201/a_8_216# OR2X1_LOC_68/B 0.01fF
C48830 AND2X1_LOC_736/Y OR2X1_LOC_528/Y 0.03fF
C48831 AND2X1_LOC_810/Y OR2X1_LOC_533/A 0.01fF
C48832 AND2X1_LOC_365/A AND2X1_LOC_802/Y 0.03fF
C48833 AND2X1_LOC_356/a_8_24# AND2X1_LOC_810/B 0.20fF
C48834 OR2X1_LOC_600/A OR2X1_LOC_165/Y 0.03fF
C48835 OR2X1_LOC_53/Y OR2X1_LOC_43/A 1.78fF
C48836 OR2X1_LOC_39/A AND2X1_LOC_249/a_8_24# 0.01fF
C48837 OR2X1_LOC_139/A OR2X1_LOC_643/A 0.07fF
C48838 OR2X1_LOC_47/Y OR2X1_LOC_152/A 0.05fF
C48839 OR2X1_LOC_40/Y AND2X1_LOC_357/a_36_24# 0.00fF
C48840 D_INPUT_0 OR2X1_LOC_112/A 0.01fF
C48841 OR2X1_LOC_139/A OR2X1_LOC_124/Y 0.02fF
C48842 OR2X1_LOC_419/Y AND2X1_LOC_486/a_36_24# 0.07fF
C48843 AND2X1_LOC_448/Y OR2X1_LOC_421/Y 0.00fF
C48844 D_INPUT_0 OR2X1_LOC_730/B 0.04fF
C48845 OR2X1_LOC_527/a_8_216# OR2X1_LOC_18/Y 0.01fF
C48846 OR2X1_LOC_377/A OR2X1_LOC_621/A 0.03fF
C48847 OR2X1_LOC_711/B OR2X1_LOC_738/A 0.10fF
C48848 AND2X1_LOC_675/A OR2X1_LOC_437/A 0.02fF
C48849 OR2X1_LOC_541/A OR2X1_LOC_274/a_8_216# 0.07fF
C48850 OR2X1_LOC_715/B OR2X1_LOC_161/A 0.10fF
C48851 AND2X1_LOC_40/Y OR2X1_LOC_648/A 0.03fF
C48852 AND2X1_LOC_325/a_8_24# AND2X1_LOC_841/B 0.03fF
C48853 OR2X1_LOC_486/B OR2X1_LOC_731/A 0.01fF
C48854 AND2X1_LOC_553/A OR2X1_LOC_56/A 0.01fF
C48855 OR2X1_LOC_49/A AND2X1_LOC_412/a_8_24# 0.01fF
C48856 OR2X1_LOC_161/A AND2X1_LOC_626/a_8_24# 0.23fF
C48857 OR2X1_LOC_43/A AND2X1_LOC_802/Y 0.02fF
C48858 OR2X1_LOC_512/A OR2X1_LOC_834/A 0.22fF
C48859 OR2X1_LOC_136/Y OR2X1_LOC_743/A 0.03fF
C48860 OR2X1_LOC_756/B OR2X1_LOC_334/B 0.01fF
C48861 AND2X1_LOC_722/Y AND2X1_LOC_723/Y 0.02fF
C48862 OR2X1_LOC_296/Y AND2X1_LOC_7/B 0.01fF
C48863 AND2X1_LOC_42/B OR2X1_LOC_392/B 0.05fF
C48864 OR2X1_LOC_56/A AND2X1_LOC_804/Y 0.03fF
C48865 OR2X1_LOC_161/A OR2X1_LOC_784/B 0.01fF
C48866 OR2X1_LOC_560/a_8_216# OR2X1_LOC_244/Y 0.00fF
C48867 AND2X1_LOC_363/B OR2X1_LOC_91/A 0.01fF
C48868 OR2X1_LOC_185/Y OR2X1_LOC_596/A 0.03fF
C48869 AND2X1_LOC_12/Y AND2X1_LOC_18/Y 0.81fF
C48870 OR2X1_LOC_476/B OR2X1_LOC_390/B 0.05fF
C48871 AND2X1_LOC_563/A AND2X1_LOC_113/Y 0.00fF
C48872 OR2X1_LOC_7/A AND2X1_LOC_786/Y 0.07fF
C48873 OR2X1_LOC_6/A AND2X1_LOC_476/Y 0.01fF
C48874 AND2X1_LOC_392/a_36_24# OR2X1_LOC_517/A 0.00fF
C48875 AND2X1_LOC_42/B AND2X1_LOC_263/a_8_24# 0.11fF
C48876 OR2X1_LOC_114/B OR2X1_LOC_500/A 0.00fF
C48877 OR2X1_LOC_7/A OR2X1_LOC_323/a_8_216# 0.07fF
C48878 OR2X1_LOC_379/a_8_216# VDD 0.00fF
C48879 AND2X1_LOC_61/a_8_24# OR2X1_LOC_32/B 0.03fF
C48880 AND2X1_LOC_228/Y OR2X1_LOC_600/A 0.03fF
C48881 OR2X1_LOC_739/Y OR2X1_LOC_739/a_8_216# -0.00fF
C48882 AND2X1_LOC_729/a_8_24# OR2X1_LOC_585/A 0.01fF
C48883 OR2X1_LOC_270/Y OR2X1_LOC_367/a_8_216# 0.03fF
C48884 OR2X1_LOC_405/A AND2X1_LOC_92/Y 0.20fF
C48885 VDD OR2X1_LOC_67/a_8_216# 0.21fF
C48886 AND2X1_LOC_719/Y AND2X1_LOC_806/A 0.01fF
C48887 OR2X1_LOC_465/Y OR2X1_LOC_471/B 0.12fF
C48888 AND2X1_LOC_40/Y AND2X1_LOC_253/a_8_24# 0.01fF
C48889 AND2X1_LOC_95/Y OR2X1_LOC_78/B 0.10fF
C48890 OR2X1_LOC_36/Y OR2X1_LOC_607/A 0.04fF
C48891 OR2X1_LOC_306/a_8_216# AND2X1_LOC_434/Y 0.01fF
C48892 OR2X1_LOC_743/a_8_216# OR2X1_LOC_39/A 0.01fF
C48893 OR2X1_LOC_633/Y OR2X1_LOC_78/B 0.00fF
C48894 AND2X1_LOC_732/B OR2X1_LOC_36/Y 0.00fF
C48895 AND2X1_LOC_149/a_8_24# AND2X1_LOC_213/B 0.01fF
C48896 OR2X1_LOC_528/Y AND2X1_LOC_620/a_8_24# 0.01fF
C48897 OR2X1_LOC_305/a_8_216# VDD 0.21fF
C48898 VDD OR2X1_LOC_213/B -0.00fF
C48899 OR2X1_LOC_696/A AND2X1_LOC_839/A 0.00fF
C48900 OR2X1_LOC_272/Y OR2X1_LOC_595/A 0.03fF
C48901 AND2X1_LOC_13/a_36_24# AND2X1_LOC_44/Y 0.00fF
C48902 AND2X1_LOC_738/B OR2X1_LOC_511/Y 0.18fF
C48903 OR2X1_LOC_744/A OR2X1_LOC_32/B 0.20fF
C48904 OR2X1_LOC_91/Y AND2X1_LOC_561/B 0.03fF
C48905 AND2X1_LOC_711/Y AND2X1_LOC_212/Y 0.12fF
C48906 OR2X1_LOC_533/Y OR2X1_LOC_70/Y 0.01fF
C48907 VDD OR2X1_LOC_69/Y 0.26fF
C48908 OR2X1_LOC_552/a_8_216# OR2X1_LOC_552/B 0.39fF
C48909 AND2X1_LOC_555/Y OR2X1_LOC_225/a_8_216# 0.01fF
C48910 OR2X1_LOC_70/Y AND2X1_LOC_212/Y 0.07fF
C48911 VDD OR2X1_LOC_418/Y 0.19fF
C48912 OR2X1_LOC_59/Y OR2X1_LOC_265/Y 0.03fF
C48913 OR2X1_LOC_809/a_8_216# OR2X1_LOC_66/A 0.01fF
C48914 OR2X1_LOC_136/Y OR2X1_LOC_246/A 0.10fF
C48915 AND2X1_LOC_42/B OR2X1_LOC_113/B 0.94fF
C48916 OR2X1_LOC_40/Y OR2X1_LOC_763/Y 0.02fF
C48917 OR2X1_LOC_176/Y AND2X1_LOC_514/Y 0.01fF
C48918 OR2X1_LOC_864/A OR2X1_LOC_66/A 0.04fF
C48919 AND2X1_LOC_41/A AND2X1_LOC_43/B 0.40fF
C48920 OR2X1_LOC_600/A OR2X1_LOC_585/A 7.57fF
C48921 OR2X1_LOC_135/Y AND2X1_LOC_307/a_8_24# 0.01fF
C48922 OR2X1_LOC_354/A OR2X1_LOC_506/A 0.03fF
C48923 AND2X1_LOC_675/Y AND2X1_LOC_580/A 0.03fF
C48924 AND2X1_LOC_95/Y OR2X1_LOC_721/Y 0.70fF
C48925 OR2X1_LOC_468/A OR2X1_LOC_155/A 0.03fF
C48926 AND2X1_LOC_385/a_36_24# OR2X1_LOC_66/A 0.00fF
C48927 OR2X1_LOC_66/A OR2X1_LOC_240/A 2.75fF
C48928 OR2X1_LOC_178/a_8_216# OR2X1_LOC_529/Y 0.01fF
C48929 OR2X1_LOC_274/a_36_216# OR2X1_LOC_375/A 0.00fF
C48930 OR2X1_LOC_84/B AND2X1_LOC_70/Y 0.00fF
C48931 OR2X1_LOC_527/Y AND2X1_LOC_475/Y 0.09fF
C48932 AND2X1_LOC_227/Y AND2X1_LOC_772/Y 0.03fF
C48933 AND2X1_LOC_845/Y AND2X1_LOC_284/a_8_24# 0.02fF
C48934 AND2X1_LOC_79/Y AND2X1_LOC_18/Y 0.03fF
C48935 OR2X1_LOC_40/Y AND2X1_LOC_578/A 0.10fF
C48936 AND2X1_LOC_735/Y AND2X1_LOC_576/Y 0.03fF
C48937 AND2X1_LOC_19/Y AND2X1_LOC_8/Y 0.03fF
C48938 OR2X1_LOC_449/B OR2X1_LOC_78/A 0.10fF
C48939 OR2X1_LOC_244/B OR2X1_LOC_203/Y 0.02fF
C48940 OR2X1_LOC_429/Y OR2X1_LOC_582/a_8_216# 0.05fF
C48941 AND2X1_LOC_514/Y AND2X1_LOC_212/Y 0.02fF
C48942 OR2X1_LOC_621/A AND2X1_LOC_670/a_8_24# 0.11fF
C48943 OR2X1_LOC_158/a_8_216# OR2X1_LOC_619/Y 0.01fF
C48944 AND2X1_LOC_496/a_8_24# AND2X1_LOC_18/Y 0.07fF
C48945 OR2X1_LOC_61/Y OR2X1_LOC_405/a_36_216# 0.02fF
C48946 OR2X1_LOC_40/Y AND2X1_LOC_632/a_8_24# 0.04fF
C48947 OR2X1_LOC_715/B AND2X1_LOC_51/Y 0.10fF
C48948 AND2X1_LOC_358/Y D_INPUT_0 0.01fF
C48949 OR2X1_LOC_697/Y OR2X1_LOC_44/Y 0.03fF
C48950 AND2X1_LOC_198/a_8_24# OR2X1_LOC_6/A 0.02fF
C48951 OR2X1_LOC_51/Y OR2X1_LOC_743/A 0.06fF
C48952 AND2X1_LOC_530/a_36_24# OR2X1_LOC_54/Y 0.01fF
C48953 OR2X1_LOC_187/a_8_216# OR2X1_LOC_613/Y 0.01fF
C48954 AND2X1_LOC_710/Y OR2X1_LOC_297/Y 0.01fF
C48955 AND2X1_LOC_567/a_8_24# AND2X1_LOC_798/Y 0.01fF
C48956 OR2X1_LOC_109/Y AND2X1_LOC_662/B 0.03fF
C48957 OR2X1_LOC_2/Y OR2X1_LOC_11/Y 0.03fF
C48958 OR2X1_LOC_656/B OR2X1_LOC_624/A 0.38fF
C48959 OR2X1_LOC_329/B AND2X1_LOC_717/B 0.07fF
C48960 OR2X1_LOC_375/A OR2X1_LOC_737/A 0.07fF
C48961 AND2X1_LOC_605/Y OR2X1_LOC_52/B 0.02fF
C48962 AND2X1_LOC_345/Y OR2X1_LOC_56/A 0.07fF
C48963 AND2X1_LOC_352/a_8_24# AND2X1_LOC_514/Y 0.03fF
C48964 OR2X1_LOC_109/a_8_216# OR2X1_LOC_39/A 0.30fF
C48965 VDD OR2X1_LOC_719/A 0.21fF
C48966 OR2X1_LOC_151/Y OR2X1_LOC_220/A 0.14fF
C48967 AND2X1_LOC_512/Y AND2X1_LOC_355/a_8_24# 0.01fF
C48968 AND2X1_LOC_360/a_8_24# AND2X1_LOC_363/A 0.02fF
C48969 OR2X1_LOC_589/A INPUT_1 0.02fF
C48970 VDD OR2X1_LOC_43/a_8_216# 0.00fF
C48971 AND2X1_LOC_95/Y OR2X1_LOC_375/A 0.22fF
C48972 AND2X1_LOC_228/Y OR2X1_LOC_619/Y 0.06fF
C48973 AND2X1_LOC_208/a_8_24# OR2X1_LOC_24/Y 0.01fF
C48974 OR2X1_LOC_633/Y OR2X1_LOC_375/A 0.05fF
C48975 AND2X1_LOC_529/a_8_24# AND2X1_LOC_42/B 0.06fF
C48976 OR2X1_LOC_620/Y OR2X1_LOC_468/Y 0.03fF
C48977 AND2X1_LOC_787/a_8_24# AND2X1_LOC_784/A 0.02fF
C48978 OR2X1_LOC_488/a_8_216# AND2X1_LOC_858/B 0.29fF
C48979 VDD AND2X1_LOC_537/Y 0.63fF
C48980 OR2X1_LOC_155/A AND2X1_LOC_424/a_36_24# 0.00fF
C48981 OR2X1_LOC_625/Y OR2X1_LOC_36/Y 0.08fF
C48982 AND2X1_LOC_386/a_8_24# OR2X1_LOC_502/A 0.01fF
C48983 OR2X1_LOC_154/A OR2X1_LOC_499/a_8_216# 0.10fF
C48984 OR2X1_LOC_664/a_36_216# OR2X1_LOC_664/Y 0.00fF
C48985 OR2X1_LOC_292/Y OR2X1_LOC_258/Y 0.03fF
C48986 OR2X1_LOC_147/A OR2X1_LOC_705/Y 0.34fF
C48987 INPUT_0 OR2X1_LOC_829/Y 0.01fF
C48988 D_INPUT_4 AND2X1_LOC_21/Y 0.01fF
C48989 AND2X1_LOC_160/Y AND2X1_LOC_708/a_36_24# 0.00fF
C48990 OR2X1_LOC_121/B OR2X1_LOC_78/A 1.47fF
C48991 OR2X1_LOC_140/B OR2X1_LOC_140/a_8_216# 0.03fF
C48992 OR2X1_LOC_112/a_36_216# OR2X1_LOC_436/Y 0.00fF
C48993 AND2X1_LOC_217/Y OR2X1_LOC_71/Y 0.00fF
C48994 INPUT_0 AND2X1_LOC_856/a_8_24# 0.03fF
C48995 GATE_366 AND2X1_LOC_848/Y 0.03fF
C48996 OR2X1_LOC_187/a_36_216# AND2X1_LOC_711/Y 0.00fF
C48997 OR2X1_LOC_160/B AND2X1_LOC_53/Y 0.52fF
C48998 AND2X1_LOC_580/A OR2X1_LOC_189/A 0.03fF
C48999 OR2X1_LOC_631/B AND2X1_LOC_43/B 0.00fF
C49000 D_INPUT_1 OR2X1_LOC_843/B 0.03fF
C49001 OR2X1_LOC_619/Y OR2X1_LOC_585/A 0.03fF
C49002 OR2X1_LOC_177/Y OR2X1_LOC_47/Y 0.06fF
C49003 OR2X1_LOC_154/A OR2X1_LOC_863/a_8_216# 0.03fF
C49004 AND2X1_LOC_842/B AND2X1_LOC_850/A 0.01fF
C49005 OR2X1_LOC_287/B OR2X1_LOC_571/B 0.03fF
C49006 OR2X1_LOC_9/Y OR2X1_LOC_62/A 0.83fF
C49007 OR2X1_LOC_18/Y AND2X1_LOC_458/a_36_24# 0.00fF
C49008 INPUT_0 AND2X1_LOC_825/a_8_24# 0.04fF
C49009 AND2X1_LOC_37/a_8_24# OR2X1_LOC_847/A 0.00fF
C49010 AND2X1_LOC_724/Y OR2X1_LOC_31/Y 0.00fF
C49011 D_INPUT_1 OR2X1_LOC_549/A 0.14fF
C49012 OR2X1_LOC_154/A AND2X1_LOC_385/a_8_24# 0.01fF
C49013 OR2X1_LOC_247/a_8_216# OR2X1_LOC_294/Y 0.40fF
C49014 INPUT_0 OR2X1_LOC_7/Y 0.03fF
C49015 OR2X1_LOC_273/Y AND2X1_LOC_649/B 0.15fF
C49016 OR2X1_LOC_121/B OR2X1_LOC_448/B 0.03fF
C49017 OR2X1_LOC_673/Y AND2X1_LOC_8/Y 0.15fF
C49018 OR2X1_LOC_51/Y OR2X1_LOC_409/B 0.03fF
C49019 OR2X1_LOC_590/Y AND2X1_LOC_591/a_8_24# 0.23fF
C49020 OR2X1_LOC_26/Y OR2X1_LOC_372/Y 0.03fF
C49021 OR2X1_LOC_316/Y OR2X1_LOC_74/A 0.03fF
C49022 OR2X1_LOC_600/A OR2X1_LOC_751/a_36_216# 0.00fF
C49023 OR2X1_LOC_160/B OR2X1_LOC_223/A 0.03fF
C49024 OR2X1_LOC_604/A OR2X1_LOC_47/Y 0.39fF
C49025 AND2X1_LOC_70/Y OR2X1_LOC_651/A 0.04fF
C49026 OR2X1_LOC_296/Y OR2X1_LOC_805/A 0.03fF
C49027 OR2X1_LOC_47/Y AND2X1_LOC_207/B 0.04fF
C49028 AND2X1_LOC_356/B AND2X1_LOC_319/A 0.33fF
C49029 AND2X1_LOC_810/Y AND2X1_LOC_468/a_8_24# 0.04fF
C49030 OR2X1_LOC_90/a_8_216# OR2X1_LOC_95/Y 0.01fF
C49031 D_INPUT_5 AND2X1_LOC_11/a_8_24# 0.01fF
C49032 OR2X1_LOC_76/a_8_216# OR2X1_LOC_736/Y 0.04fF
C49033 OR2X1_LOC_488/a_8_216# AND2X1_LOC_573/A 0.02fF
C49034 VDD OR2X1_LOC_437/a_8_216# 0.21fF
C49035 AND2X1_LOC_654/Y AND2X1_LOC_863/A 0.02fF
C49036 AND2X1_LOC_367/A AND2X1_LOC_863/Y 0.01fF
C49037 OR2X1_LOC_449/B OR2X1_LOC_155/A 0.07fF
C49038 OR2X1_LOC_709/A OR2X1_LOC_728/B 0.05fF
C49039 OR2X1_LOC_70/Y OR2X1_LOC_265/Y 8.97fF
C49040 INPUT_1 AND2X1_LOC_618/a_8_24# 0.14fF
C49041 AND2X1_LOC_840/B OR2X1_LOC_371/Y 0.19fF
C49042 OR2X1_LOC_499/B AND2X1_LOC_47/Y 0.03fF
C49043 AND2X1_LOC_489/Y AND2X1_LOC_361/A 0.02fF
C49044 OR2X1_LOC_756/B OR2X1_LOC_439/a_36_216# 0.00fF
C49045 OR2X1_LOC_254/B OR2X1_LOC_254/a_8_216# 0.01fF
C49046 OR2X1_LOC_291/a_8_216# OR2X1_LOC_62/B 0.01fF
C49047 OR2X1_LOC_854/a_8_216# OR2X1_LOC_532/B 0.01fF
C49048 AND2X1_LOC_86/Y AND2X1_LOC_133/a_8_24# 0.03fF
C49049 OR2X1_LOC_549/a_8_216# D_GATE_366 0.01fF
C49050 OR2X1_LOC_481/A AND2X1_LOC_359/B 0.01fF
C49051 VDD OR2X1_LOC_774/B 0.30fF
C49052 OR2X1_LOC_502/A OR2X1_LOC_436/Y 0.03fF
C49053 OR2X1_LOC_696/Y OR2X1_LOC_44/Y 0.03fF
C49054 OR2X1_LOC_629/A AND2X1_LOC_3/Y 0.18fF
C49055 AND2X1_LOC_303/A OR2X1_LOC_416/Y 0.00fF
C49056 OR2X1_LOC_858/A OR2X1_LOC_241/B 0.02fF
C49057 OR2X1_LOC_309/Y AND2X1_LOC_222/Y 0.01fF
C49058 OR2X1_LOC_87/A AND2X1_LOC_442/a_8_24# 0.01fF
C49059 AND2X1_LOC_64/Y AND2X1_LOC_591/a_8_24# 0.01fF
C49060 OR2X1_LOC_286/Y OR2X1_LOC_286/B 0.00fF
C49061 OR2X1_LOC_814/A OR2X1_LOC_340/Y 0.35fF
C49062 VDD OR2X1_LOC_675/Y 0.46fF
C49063 OR2X1_LOC_563/A OR2X1_LOC_777/B 0.07fF
C49064 OR2X1_LOC_40/Y OR2X1_LOC_746/Y 0.06fF
C49065 OR2X1_LOC_59/Y AND2X1_LOC_205/a_8_24# 0.02fF
C49066 OR2X1_LOC_22/Y AND2X1_LOC_319/A 0.07fF
C49067 OR2X1_LOC_426/Y AND2X1_LOC_451/Y 0.01fF
C49068 OR2X1_LOC_130/A OR2X1_LOC_814/A 0.19fF
C49069 OR2X1_LOC_89/A AND2X1_LOC_260/a_8_24# 0.01fF
C49070 AND2X1_LOC_342/a_8_24# OR2X1_LOC_54/Y 0.01fF
C49071 OR2X1_LOC_16/A OR2X1_LOC_300/a_8_216# 0.11fF
C49072 AND2X1_LOC_706/Y AND2X1_LOC_592/a_8_24# 0.04fF
C49073 OR2X1_LOC_121/B OR2X1_LOC_155/A 1.92fF
C49074 AND2X1_LOC_48/A OR2X1_LOC_200/a_36_216# 0.00fF
C49075 OR2X1_LOC_32/B OR2X1_LOC_31/Y 0.11fF
C49076 OR2X1_LOC_135/Y OR2X1_LOC_13/B 0.03fF
C49077 AND2X1_LOC_831/Y AND2X1_LOC_655/A 0.09fF
C49078 VDD AND2X1_LOC_796/A 0.75fF
C49079 AND2X1_LOC_22/Y OR2X1_LOC_539/B 0.02fF
C49080 OR2X1_LOC_612/B OR2X1_LOC_46/A 0.13fF
C49081 OR2X1_LOC_744/A AND2X1_LOC_222/Y 0.03fF
C49082 OR2X1_LOC_619/Y AND2X1_LOC_645/a_8_24# 0.02fF
C49083 OR2X1_LOC_43/A INPUT_1 0.17fF
C49084 INPUT_3 OR2X1_LOC_673/A 0.10fF
C49085 OR2X1_LOC_499/B OR2X1_LOC_598/A 0.00fF
C49086 OR2X1_LOC_7/Y OR2X1_LOC_690/A 0.60fF
C49087 OR2X1_LOC_283/a_8_216# OR2X1_LOC_417/A 0.01fF
C49088 OR2X1_LOC_461/a_36_216# OR2X1_LOC_68/B 0.00fF
C49089 OR2X1_LOC_249/Y AND2X1_LOC_250/a_8_24# 0.01fF
C49090 OR2X1_LOC_373/Y OR2X1_LOC_142/Y 0.07fF
C49091 OR2X1_LOC_605/A OR2X1_LOC_121/B 0.01fF
C49092 AND2X1_LOC_785/A AND2X1_LOC_721/Y 0.00fF
C49093 AND2X1_LOC_164/a_8_24# AND2X1_LOC_31/Y 0.01fF
C49094 OR2X1_LOC_497/Y OR2X1_LOC_226/Y 0.11fF
C49095 OR2X1_LOC_813/a_36_216# OR2X1_LOC_71/A 0.00fF
C49096 AND2X1_LOC_43/B OR2X1_LOC_207/a_8_216# 0.03fF
C49097 OR2X1_LOC_62/A OR2X1_LOC_96/B 0.12fF
C49098 OR2X1_LOC_831/a_36_216# OR2X1_LOC_223/A 0.00fF
C49099 OR2X1_LOC_446/Y AND2X1_LOC_3/Y 0.04fF
C49100 OR2X1_LOC_80/Y OR2X1_LOC_47/Y 0.01fF
C49101 OR2X1_LOC_634/a_8_216# OR2X1_LOC_68/B 0.01fF
C49102 AND2X1_LOC_17/Y OR2X1_LOC_651/A 0.01fF
C49103 OR2X1_LOC_62/A AND2X1_LOC_852/Y 0.07fF
C49104 OR2X1_LOC_711/B AND2X1_LOC_36/Y 0.08fF
C49105 OR2X1_LOC_677/Y AND2X1_LOC_796/A 0.03fF
C49106 AND2X1_LOC_356/B AND2X1_LOC_170/B 0.82fF
C49107 D_INPUT_5 OR2X1_LOC_377/a_8_216# 0.02fF
C49108 OR2X1_LOC_744/A OR2X1_LOC_423/Y 0.15fF
C49109 AND2X1_LOC_50/Y AND2X1_LOC_31/Y 0.07fF
C49110 OR2X1_LOC_216/A OR2X1_LOC_560/A 0.02fF
C49111 AND2X1_LOC_42/B OR2X1_LOC_532/B 0.86fF
C49112 AND2X1_LOC_650/a_8_24# D_INPUT_0 0.01fF
C49113 AND2X1_LOC_641/a_8_24# OR2X1_LOC_265/Y 0.07fF
C49114 OR2X1_LOC_36/Y OR2X1_LOC_3/B 0.01fF
C49115 OR2X1_LOC_479/Y OR2X1_LOC_440/A 0.07fF
C49116 AND2X1_LOC_76/Y OR2X1_LOC_153/a_36_216# 0.00fF
C49117 OR2X1_LOC_231/a_8_216# OR2X1_LOC_641/B 0.01fF
C49118 OR2X1_LOC_78/B OR2X1_LOC_788/B 0.04fF
C49119 OR2X1_LOC_69/Y OR2X1_LOC_67/Y 0.01fF
C49120 OR2X1_LOC_473/A AND2X1_LOC_3/Y 0.78fF
C49121 OR2X1_LOC_549/B OR2X1_LOC_549/A 0.04fF
C49122 OR2X1_LOC_364/A OR2X1_LOC_374/Y 0.26fF
C49123 OR2X1_LOC_160/A OR2X1_LOC_160/a_8_216# 0.18fF
C49124 OR2X1_LOC_223/A OR2X1_LOC_794/a_8_216# 0.00fF
C49125 AND2X1_LOC_476/a_8_24# AND2X1_LOC_786/Y 0.05fF
C49126 OR2X1_LOC_62/B OR2X1_LOC_814/A 0.03fF
C49127 OR2X1_LOC_401/Y D_INPUT_1 0.03fF
C49128 AND2X1_LOC_231/Y AND2X1_LOC_341/a_8_24# 0.00fF
C49129 OR2X1_LOC_361/a_36_216# OR2X1_LOC_140/B 0.00fF
C49130 OR2X1_LOC_639/a_36_216# AND2X1_LOC_51/Y 0.00fF
C49131 OR2X1_LOC_3/Y AND2X1_LOC_687/a_8_24# 0.01fF
C49132 AND2X1_LOC_795/Y OR2X1_LOC_52/B 0.00fF
C49133 OR2X1_LOC_344/A OR2X1_LOC_563/A 0.02fF
C49134 OR2X1_LOC_16/A AND2X1_LOC_208/Y 0.00fF
C49135 OR2X1_LOC_78/B OR2X1_LOC_175/a_8_216# 0.01fF
C49136 OR2X1_LOC_59/Y OR2X1_LOC_183/a_8_216# 0.01fF
C49137 AND2X1_LOC_216/A AND2X1_LOC_361/A 0.02fF
C49138 AND2X1_LOC_12/Y OR2X1_LOC_789/A 0.07fF
C49139 AND2X1_LOC_64/Y OR2X1_LOC_661/A 0.02fF
C49140 OR2X1_LOC_350/a_8_216# OR2X1_LOC_228/Y 0.01fF
C49141 AND2X1_LOC_133/a_8_24# OR2X1_LOC_244/A 0.03fF
C49142 OR2X1_LOC_92/Y OR2X1_LOC_437/A 0.41fF
C49143 AND2X1_LOC_563/a_8_24# AND2X1_LOC_657/A 0.04fF
C49144 VDD OR2X1_LOC_743/Y 0.12fF
C49145 AND2X1_LOC_840/B AND2X1_LOC_222/Y 0.05fF
C49146 OR2X1_LOC_161/B AND2X1_LOC_279/a_8_24# 0.11fF
C49147 OR2X1_LOC_599/A AND2X1_LOC_779/Y 0.04fF
C49148 OR2X1_LOC_39/A AND2X1_LOC_215/a_8_24# 0.01fF
C49149 OR2X1_LOC_66/A OR2X1_LOC_397/a_8_216# 0.03fF
C49150 OR2X1_LOC_3/Y AND2X1_LOC_793/Y 0.06fF
C49151 OR2X1_LOC_648/B AND2X1_LOC_7/B 0.00fF
C49152 OR2X1_LOC_702/A OR2X1_LOC_801/B 0.05fF
C49153 OR2X1_LOC_40/Y AND2X1_LOC_202/Y 0.01fF
C49154 OR2X1_LOC_756/B OR2X1_LOC_577/B 1.16fF
C49155 AND2X1_LOC_472/a_36_24# OR2X1_LOC_46/A 0.00fF
C49156 AND2X1_LOC_564/B OR2X1_LOC_600/A 1.63fF
C49157 AND2X1_LOC_82/Y AND2X1_LOC_83/a_8_24# 0.11fF
C49158 OR2X1_LOC_146/a_8_216# OR2X1_LOC_51/Y 0.15fF
C49159 OR2X1_LOC_600/A OR2X1_LOC_230/Y 0.14fF
C49160 OR2X1_LOC_132/a_8_216# OR2X1_LOC_134/Y 0.05fF
C49161 AND2X1_LOC_356/B OR2X1_LOC_331/Y 0.01fF
C49162 AND2X1_LOC_465/A OR2X1_LOC_56/A 0.22fF
C49163 AND2X1_LOC_592/Y OR2X1_LOC_12/Y 0.06fF
C49164 AND2X1_LOC_3/Y OR2X1_LOC_228/Y 0.10fF
C49165 OR2X1_LOC_502/A OR2X1_LOC_395/Y 0.03fF
C49166 AND2X1_LOC_544/Y AND2X1_LOC_663/A 0.41fF
C49167 AND2X1_LOC_721/Y AND2X1_LOC_658/A 0.03fF
C49168 AND2X1_LOC_61/Y AND2X1_LOC_206/a_8_24# 0.02fF
C49169 OR2X1_LOC_74/A OR2X1_LOC_153/a_8_216# 0.05fF
C49170 OR2X1_LOC_589/A AND2X1_LOC_130/a_8_24# 0.11fF
C49171 AND2X1_LOC_645/A OR2X1_LOC_533/A 0.00fF
C49172 OR2X1_LOC_188/Y OR2X1_LOC_858/A 0.82fF
C49173 AND2X1_LOC_192/Y AND2X1_LOC_742/A 0.13fF
C49174 AND2X1_LOC_740/B AND2X1_LOC_738/Y 0.09fF
C49175 OR2X1_LOC_589/A AND2X1_LOC_729/a_36_24# 0.01fF
C49176 OR2X1_LOC_304/a_8_216# OR2X1_LOC_59/Y 0.01fF
C49177 OR2X1_LOC_375/A AND2X1_LOC_41/Y 1.03fF
C49178 OR2X1_LOC_6/B AND2X1_LOC_65/A 0.16fF
C49179 AND2X1_LOC_841/a_36_24# OR2X1_LOC_31/Y -0.00fF
C49180 AND2X1_LOC_383/a_36_24# OR2X1_LOC_91/A 0.01fF
C49181 AND2X1_LOC_22/Y OR2X1_LOC_78/B 0.34fF
C49182 VDD OR2X1_LOC_736/Y 0.18fF
C49183 AND2X1_LOC_658/B AND2X1_LOC_212/Y 0.07fF
C49184 OR2X1_LOC_243/A AND2X1_LOC_36/Y 0.01fF
C49185 OR2X1_LOC_186/Y AND2X1_LOC_70/Y 0.42fF
C49186 AND2X1_LOC_772/B OR2X1_LOC_12/Y 0.03fF
C49187 OR2X1_LOC_696/A OR2X1_LOC_427/A 0.91fF
C49188 OR2X1_LOC_473/Y AND2X1_LOC_31/Y 0.02fF
C49189 OR2X1_LOC_614/Y VDD 0.37fF
C49190 OR2X1_LOC_379/Y OR2X1_LOC_598/a_8_216# 0.01fF
C49191 OR2X1_LOC_696/A AND2X1_LOC_801/a_8_24# -0.07fF
C49192 VDD OR2X1_LOC_13/Y 0.20fF
C49193 D_INPUT_3 AND2X1_LOC_8/a_8_24# 0.07fF
C49194 OR2X1_LOC_318/a_36_216# AND2X1_LOC_92/Y 0.01fF
C49195 OR2X1_LOC_45/B OR2X1_LOC_697/Y 0.18fF
C49196 OR2X1_LOC_8/Y OR2X1_LOC_9/Y 2.63fF
C49197 OR2X1_LOC_254/A OR2X1_LOC_563/A 0.03fF
C49198 OR2X1_LOC_696/A OR2X1_LOC_823/Y 0.01fF
C49199 OR2X1_LOC_482/Y AND2X1_LOC_658/A 0.33fF
C49200 AND2X1_LOC_22/Y OR2X1_LOC_721/Y 0.03fF
C49201 OR2X1_LOC_323/A OR2X1_LOC_109/Y 0.01fF
C49202 AND2X1_LOC_549/Y VDD 0.25fF
C49203 OR2X1_LOC_575/A OR2X1_LOC_563/A 0.02fF
C49204 OR2X1_LOC_756/B OR2X1_LOC_756/a_36_216# 0.03fF
C49205 OR2X1_LOC_186/Y OR2X1_LOC_703/A 0.17fF
C49206 AND2X1_LOC_715/Y AND2X1_LOC_801/a_8_24# 0.02fF
C49207 AND2X1_LOC_709/a_36_24# OR2X1_LOC_600/A -0.00fF
C49208 OR2X1_LOC_276/B OR2X1_LOC_66/Y 0.03fF
C49209 OR2X1_LOC_621/B OR2X1_LOC_78/A 0.39fF
C49210 OR2X1_LOC_151/A OR2X1_LOC_630/B 0.02fF
C49211 VDD OR2X1_LOC_627/Y 0.10fF
C49212 OR2X1_LOC_50/a_8_216# OR2X1_LOC_51/B 0.39fF
C49213 AND2X1_LOC_53/Y OR2X1_LOC_197/a_8_216# 0.06fF
C49214 VDD AND2X1_LOC_500/Y 0.07fF
C49215 AND2X1_LOC_805/Y GATE_579 0.00fF
C49216 OR2X1_LOC_47/Y OR2X1_LOC_747/a_8_216# 0.18fF
C49217 OR2X1_LOC_653/Y AND2X1_LOC_44/Y 0.07fF
C49218 OR2X1_LOC_663/A OR2X1_LOC_113/B 0.01fF
C49219 OR2X1_LOC_31/Y AND2X1_LOC_222/Y 0.03fF
C49220 AND2X1_LOC_738/B OR2X1_LOC_600/a_8_216# 0.31fF
C49221 AND2X1_LOC_337/a_8_24# AND2X1_LOC_352/B 0.01fF
C49222 OR2X1_LOC_496/a_36_216# AND2X1_LOC_658/A 0.02fF
C49223 OR2X1_LOC_589/A OR2X1_LOC_517/A 0.05fF
C49224 OR2X1_LOC_309/Y AND2X1_LOC_367/A 0.06fF
C49225 OR2X1_LOC_97/A OR2X1_LOC_185/A 0.03fF
C49226 OR2X1_LOC_51/Y AND2X1_LOC_510/A 0.02fF
C49227 AND2X1_LOC_856/B OR2X1_LOC_13/B 0.01fF
C49228 OR2X1_LOC_51/Y OR2X1_LOC_12/a_8_216# 0.01fF
C49229 OR2X1_LOC_44/Y OR2X1_LOC_503/a_8_216# 0.01fF
C49230 AND2X1_LOC_341/a_36_24# OR2X1_LOC_619/Y 0.01fF
C49231 AND2X1_LOC_22/Y OR2X1_LOC_375/A 0.32fF
C49232 OR2X1_LOC_710/B OR2X1_LOC_147/A 0.04fF
C49233 D_INPUT_0 OR2X1_LOC_71/A 0.23fF
C49234 AND2X1_LOC_19/Y AND2X1_LOC_92/Y 0.12fF
C49235 OR2X1_LOC_364/A OR2X1_LOC_392/B 0.01fF
C49236 OR2X1_LOC_40/Y AND2X1_LOC_335/a_36_24# 0.00fF
C49237 OR2X1_LOC_510/Y OR2X1_LOC_576/A 0.00fF
C49238 AND2X1_LOC_347/Y OR2X1_LOC_600/A 0.03fF
C49239 OR2X1_LOC_185/Y OR2X1_LOC_392/B 0.05fF
C49240 OR2X1_LOC_600/A AND2X1_LOC_857/Y 0.03fF
C49241 OR2X1_LOC_659/B OR2X1_LOC_720/Y -0.00fF
C49242 VDD OR2X1_LOC_808/B 2.03fF
C49243 OR2X1_LOC_680/A OR2X1_LOC_373/a_36_216# 0.01fF
C49244 AND2X1_LOC_95/Y OR2X1_LOC_549/A 0.08fF
C49245 AND2X1_LOC_570/Y AND2X1_LOC_508/A 0.00fF
C49246 OR2X1_LOC_160/B OR2X1_LOC_502/A 0.10fF
C49247 OR2X1_LOC_739/A OR2X1_LOC_486/Y 0.12fF
C49248 OR2X1_LOC_804/A OR2X1_LOC_318/B 0.01fF
C49249 OR2X1_LOC_770/B AND2X1_LOC_817/B 0.00fF
C49250 OR2X1_LOC_633/Y OR2X1_LOC_549/A 0.00fF
C49251 OR2X1_LOC_31/Y OR2X1_LOC_423/Y 0.02fF
C49252 AND2X1_LOC_342/Y OR2X1_LOC_12/Y 0.30fF
C49253 OR2X1_LOC_51/Y OR2X1_LOC_425/a_8_216# 0.39fF
C49254 OR2X1_LOC_348/a_36_216# OR2X1_LOC_791/B 0.00fF
C49255 AND2X1_LOC_176/a_8_24# OR2X1_LOC_168/Y 0.03fF
C49256 OR2X1_LOC_106/a_36_216# AND2X1_LOC_99/A 0.00fF
C49257 OR2X1_LOC_49/A AND2X1_LOC_852/a_8_24# 0.08fF
C49258 AND2X1_LOC_367/A OR2X1_LOC_744/A 0.10fF
C49259 AND2X1_LOC_715/A OR2X1_LOC_92/Y 0.16fF
C49260 AND2X1_LOC_787/A AND2X1_LOC_784/A 0.19fF
C49261 OR2X1_LOC_89/A AND2X1_LOC_773/a_8_24# 0.03fF
C49262 AND2X1_LOC_177/a_8_24# AND2X1_LOC_437/a_8_24# 0.23fF
C49263 AND2X1_LOC_347/Y AND2X1_LOC_296/a_8_24# 0.08fF
C49264 OR2X1_LOC_706/A OR2X1_LOC_78/B 0.03fF
C49265 AND2X1_LOC_12/Y AND2X1_LOC_275/a_8_24# 0.02fF
C49266 AND2X1_LOC_863/a_8_24# OR2X1_LOC_56/A 0.01fF
C49267 AND2X1_LOC_374/a_8_24# OR2X1_LOC_51/Y 0.02fF
C49268 OR2X1_LOC_164/Y OR2X1_LOC_59/Y 0.03fF
C49269 OR2X1_LOC_396/a_8_216# OR2X1_LOC_80/A 0.03fF
C49270 AND2X1_LOC_810/A AND2X1_LOC_354/B 0.04fF
C49271 OR2X1_LOC_357/a_36_216# OR2X1_LOC_87/A 0.00fF
C49272 AND2X1_LOC_540/a_8_24# OR2X1_LOC_59/Y 0.01fF
C49273 OR2X1_LOC_205/Y OR2X1_LOC_560/A 0.04fF
C49274 OR2X1_LOC_604/A OR2X1_LOC_625/Y 0.10fF
C49275 AND2X1_LOC_194/a_8_24# INPUT_0 0.17fF
C49276 AND2X1_LOC_12/Y OR2X1_LOC_307/A 0.01fF
C49277 OR2X1_LOC_637/Y OR2X1_LOC_638/a_8_216# 0.18fF
C49278 OR2X1_LOC_335/a_36_216# OR2X1_LOC_479/Y 0.01fF
C49279 AND2X1_LOC_719/Y AND2X1_LOC_287/a_36_24# 0.01fF
C49280 OR2X1_LOC_129/a_8_216# OR2X1_LOC_32/B 0.03fF
C49281 AND2X1_LOC_8/Y AND2X1_LOC_277/a_8_24# 0.01fF
C49282 OR2X1_LOC_784/Y OR2X1_LOC_66/A 0.01fF
C49283 OR2X1_LOC_154/A OR2X1_LOC_851/B 0.02fF
C49284 OR2X1_LOC_160/B OR2X1_LOC_571/B 0.01fF
C49285 AND2X1_LOC_61/Y AND2X1_LOC_76/Y 0.00fF
C49286 AND2X1_LOC_381/a_8_24# OR2X1_LOC_6/B 0.26fF
C49287 OR2X1_LOC_486/Y AND2X1_LOC_298/a_8_24# 0.03fF
C49288 OR2X1_LOC_525/Y OR2X1_LOC_51/Y 0.03fF
C49289 AND2X1_LOC_398/a_36_24# OR2X1_LOC_600/A 0.01fF
C49290 OR2X1_LOC_185/Y OR2X1_LOC_113/B 0.05fF
C49291 AND2X1_LOC_51/Y OR2X1_LOC_338/B 0.05fF
C49292 AND2X1_LOC_371/a_8_24# AND2X1_LOC_59/Y 0.03fF
C49293 AND2X1_LOC_347/B AND2X1_LOC_848/a_36_24# 0.00fF
C49294 OR2X1_LOC_700/Y VDD 0.04fF
C49295 OR2X1_LOC_244/B OR2X1_LOC_721/Y 1.26fF
C49296 OR2X1_LOC_434/A OR2X1_LOC_539/B 0.05fF
C49297 AND2X1_LOC_252/a_8_24# OR2X1_LOC_344/A 0.01fF
C49298 OR2X1_LOC_517/A OR2X1_LOC_275/Y 0.09fF
C49299 AND2X1_LOC_773/Y OR2X1_LOC_89/A 0.57fF
C49300 OR2X1_LOC_486/Y OR2X1_LOC_269/B 0.07fF
C49301 OR2X1_LOC_325/Y AND2X1_LOC_95/Y 0.04fF
C49302 AND2X1_LOC_59/Y AND2X1_LOC_18/Y 1.23fF
C49303 OR2X1_LOC_287/B OR2X1_LOC_489/A 0.00fF
C49304 OR2X1_LOC_756/Y OR2X1_LOC_791/A 0.01fF
C49305 OR2X1_LOC_304/a_8_216# OR2X1_LOC_70/Y 0.01fF
C49306 AND2X1_LOC_476/Y OR2X1_LOC_44/Y 0.09fF
C49307 AND2X1_LOC_649/a_8_24# AND2X1_LOC_219/Y 0.01fF
C49308 AND2X1_LOC_362/B OR2X1_LOC_44/Y 0.85fF
C49309 AND2X1_LOC_22/Y OR2X1_LOC_605/B 0.03fF
C49310 OR2X1_LOC_45/Y AND2X1_LOC_434/Y 0.95fF
C49311 AND2X1_LOC_378/a_36_24# OR2X1_LOC_689/A 0.00fF
C49312 AND2X1_LOC_130/a_8_24# OR2X1_LOC_43/A 0.02fF
C49313 AND2X1_LOC_784/A AND2X1_LOC_566/B 0.03fF
C49314 AND2X1_LOC_464/A OR2X1_LOC_371/Y 0.13fF
C49315 OR2X1_LOC_87/A OR2X1_LOC_641/A 0.08fF
C49316 OR2X1_LOC_174/A OR2X1_LOC_61/Y 0.01fF
C49317 AND2X1_LOC_365/A AND2X1_LOC_352/B 0.11fF
C49318 AND2X1_LOC_339/B AND2X1_LOC_339/a_8_24# 0.04fF
C49319 AND2X1_LOC_550/A AND2X1_LOC_663/A 0.49fF
C49320 OR2X1_LOC_676/a_8_216# AND2X1_LOC_56/B 0.01fF
C49321 OR2X1_LOC_456/A OR2X1_LOC_563/A 0.04fF
C49322 OR2X1_LOC_648/A AND2X1_LOC_43/B 0.07fF
C49323 OR2X1_LOC_113/Y AND2X1_LOC_95/Y 0.00fF
C49324 OR2X1_LOC_9/Y OR2X1_LOC_672/Y 0.53fF
C49325 OR2X1_LOC_476/B OR2X1_LOC_390/a_36_216# 0.03fF
C49326 OR2X1_LOC_26/Y AND2X1_LOC_243/Y 0.10fF
C49327 OR2X1_LOC_40/Y OR2X1_LOC_670/Y 0.02fF
C49328 OR2X1_LOC_45/B OR2X1_LOC_696/Y 0.03fF
C49329 OR2X1_LOC_377/A AND2X1_LOC_232/a_8_24# 0.01fF
C49330 OR2X1_LOC_237/Y OR2X1_LOC_56/A 0.03fF
C49331 OR2X1_LOC_8/Y OR2X1_LOC_96/B 0.18fF
C49332 AND2X1_LOC_81/B AND2X1_LOC_70/Y 0.00fF
C49333 OR2X1_LOC_70/Y AND2X1_LOC_809/a_8_24# 0.11fF
C49334 AND2X1_LOC_618/a_8_24# AND2X1_LOC_619/B 0.00fF
C49335 AND2X1_LOC_657/A AND2X1_LOC_563/Y 0.02fF
C49336 AND2X1_LOC_99/A AND2X1_LOC_98/Y 0.02fF
C49337 AND2X1_LOC_141/B OR2X1_LOC_12/Y 0.03fF
C49338 VDD OR2X1_LOC_82/a_8_216# 0.21fF
C49339 AND2X1_LOC_70/Y OR2X1_LOC_358/B 0.02fF
C49340 OR2X1_LOC_490/a_8_216# OR2X1_LOC_70/Y 0.02fF
C49341 AND2X1_LOC_535/Y AND2X1_LOC_854/a_36_24# 0.01fF
C49342 OR2X1_LOC_11/Y OR2X1_LOC_25/Y 0.03fF
C49343 AND2X1_LOC_719/Y OR2X1_LOC_529/Y 0.03fF
C49344 AND2X1_LOC_568/B OR2X1_LOC_26/Y 0.01fF
C49345 OR2X1_LOC_271/Y AND2X1_LOC_715/A 0.16fF
C49346 OR2X1_LOC_9/Y OR2X1_LOC_73/a_36_216# 0.03fF
C49347 AND2X1_LOC_390/B OR2X1_LOC_13/a_36_216# 0.01fF
C49348 OR2X1_LOC_235/B OR2X1_LOC_39/A 0.01fF
C49349 OR2X1_LOC_287/B OR2X1_LOC_772/A 0.02fF
C49350 OR2X1_LOC_601/Y AND2X1_LOC_447/Y 0.05fF
C49351 OR2X1_LOC_653/Y OR2X1_LOC_61/a_8_216# 0.03fF
C49352 OR2X1_LOC_495/Y AND2X1_LOC_833/a_8_24# 0.01fF
C49353 VDD OR2X1_LOC_708/B 0.02fF
C49354 AND2X1_LOC_51/Y OR2X1_LOC_35/A 0.01fF
C49355 OR2X1_LOC_744/A AND2X1_LOC_114/a_36_24# 0.01fF
C49356 AND2X1_LOC_372/a_8_24# OR2X1_LOC_805/A 0.03fF
C49357 OR2X1_LOC_89/A AND2X1_LOC_243/Y 0.08fF
C49358 OR2X1_LOC_8/Y AND2X1_LOC_852/Y 0.19fF
C49359 AND2X1_LOC_857/Y OR2X1_LOC_619/Y 0.04fF
C49360 AND2X1_LOC_95/Y OR2X1_LOC_354/A 0.42fF
C49361 AND2X1_LOC_86/Y OR2X1_LOC_502/A 0.00fF
C49362 OR2X1_LOC_244/B OR2X1_LOC_375/A 0.04fF
C49363 OR2X1_LOC_681/a_8_216# OR2X1_LOC_7/A 0.03fF
C49364 OR2X1_LOC_52/Y OR2X1_LOC_16/A 0.02fF
C49365 AND2X1_LOC_574/a_8_24# OR2X1_LOC_680/A 0.05fF
C49366 OR2X1_LOC_787/Y OR2X1_LOC_543/A 0.81fF
C49367 AND2X1_LOC_41/A OR2X1_LOC_510/Y 0.01fF
C49368 AND2X1_LOC_61/Y OR2X1_LOC_52/B 0.00fF
C49369 OR2X1_LOC_8/Y OR2X1_LOC_6/a_36_216# 0.02fF
C49370 INPUT_3 OR2X1_LOC_502/A 2.49fF
C49371 OR2X1_LOC_706/A OR2X1_LOC_375/A 0.01fF
C49372 AND2X1_LOC_712/B OR2X1_LOC_12/Y 0.12fF
C49373 OR2X1_LOC_185/A OR2X1_LOC_475/B 0.04fF
C49374 OR2X1_LOC_54/Y OR2X1_LOC_12/Y 0.02fF
C49375 AND2X1_LOC_312/a_8_24# OR2X1_LOC_87/A 0.04fF
C49376 AND2X1_LOC_59/Y OR2X1_LOC_473/a_8_216# 0.01fF
C49377 OR2X1_LOC_709/A OR2X1_LOC_196/B 0.00fF
C49378 AND2X1_LOC_729/Y AND2X1_LOC_147/a_8_24# 0.01fF
C49379 OR2X1_LOC_3/Y AND2X1_LOC_363/Y 0.01fF
C49380 AND2X1_LOC_861/B AND2X1_LOC_859/Y 0.01fF
C49381 AND2X1_LOC_94/Y OR2X1_LOC_240/A 0.07fF
C49382 OR2X1_LOC_91/Y AND2X1_LOC_553/A 0.03fF
C49383 OR2X1_LOC_160/A OR2X1_LOC_620/Y 0.39fF
C49384 AND2X1_LOC_198/a_8_24# OR2X1_LOC_44/Y 0.01fF
C49385 AND2X1_LOC_456/Y OR2X1_LOC_744/A 0.00fF
C49386 OR2X1_LOC_611/Y OR2X1_LOC_16/A 0.01fF
C49387 OR2X1_LOC_43/A OR2X1_LOC_517/A 0.10fF
C49388 AND2X1_LOC_41/A OR2X1_LOC_810/A 0.03fF
C49389 OR2X1_LOC_45/a_36_216# OR2X1_LOC_48/B 0.00fF
C49390 OR2X1_LOC_662/A OR2X1_LOC_655/a_8_216# 0.02fF
C49391 OR2X1_LOC_490/Y OR2X1_LOC_744/A 0.20fF
C49392 OR2X1_LOC_744/A OR2X1_LOC_74/A 0.10fF
C49393 OR2X1_LOC_91/Y AND2X1_LOC_804/Y 0.09fF
C49394 AND2X1_LOC_348/Y OR2X1_LOC_92/Y 0.03fF
C49395 AND2X1_LOC_784/Y AND2X1_LOC_727/A 0.02fF
C49396 OR2X1_LOC_525/Y OR2X1_LOC_680/A 0.02fF
C49397 OR2X1_LOC_18/Y OR2X1_LOC_45/a_36_216# 0.02fF
C49398 AND2X1_LOC_810/A AND2X1_LOC_863/Y 0.14fF
C49399 AND2X1_LOC_578/A OR2X1_LOC_531/Y 0.05fF
C49400 OR2X1_LOC_402/a_36_216# OR2X1_LOC_78/A 0.00fF
C49401 OR2X1_LOC_402/a_8_216# OR2X1_LOC_78/a_8_216# 0.47fF
C49402 OR2X1_LOC_777/B OR2X1_LOC_724/A 0.02fF
C49403 OR2X1_LOC_92/Y OR2X1_LOC_753/A 0.17fF
C49404 OR2X1_LOC_841/a_8_216# OR2X1_LOC_155/A 0.01fF
C49405 OR2X1_LOC_624/Y AND2X1_LOC_42/B 0.02fF
C49406 AND2X1_LOC_621/Y AND2X1_LOC_622/a_36_24# 0.01fF
C49407 OR2X1_LOC_160/B AND2X1_LOC_48/A 4.50fF
C49408 OR2X1_LOC_176/Y OR2X1_LOC_47/Y 0.28fF
C49409 VDD OR2X1_LOC_295/Y 0.04fF
C49410 OR2X1_LOC_154/A OR2X1_LOC_160/A 0.27fF
C49411 AND2X1_LOC_359/a_8_24# OR2X1_LOC_427/A 0.05fF
C49412 OR2X1_LOC_790/B OR2X1_LOC_793/A 0.80fF
C49413 AND2X1_LOC_139/B AND2X1_LOC_655/A 0.08fF
C49414 OR2X1_LOC_92/Y OR2X1_LOC_754/a_8_216# 0.01fF
C49415 AND2X1_LOC_76/Y OR2X1_LOC_74/a_36_216# 0.00fF
C49416 OR2X1_LOC_856/B OR2X1_LOC_155/A 0.39fF
C49417 OR2X1_LOC_833/Y OR2X1_LOC_276/B 0.00fF
C49418 OR2X1_LOC_68/B AND2X1_LOC_238/a_8_24# 0.02fF
C49419 AND2X1_LOC_67/a_8_24# AND2X1_LOC_67/Y 0.03fF
C49420 OR2X1_LOC_748/A AND2X1_LOC_847/Y 0.01fF
C49421 AND2X1_LOC_458/Y AND2X1_LOC_464/a_8_24# 0.19fF
C49422 OR2X1_LOC_848/B OR2X1_LOC_848/a_8_216# 0.00fF
C49423 OR2X1_LOC_468/A OR2X1_LOC_814/A 0.05fF
C49424 AND2X1_LOC_182/A AND2X1_LOC_866/A 0.25fF
C49425 OR2X1_LOC_427/A OR2X1_LOC_89/a_8_216# 0.02fF
C49426 OR2X1_LOC_106/A OR2X1_LOC_278/Y 0.01fF
C49427 OR2X1_LOC_62/B OR2X1_LOC_244/Y 0.08fF
C49428 OR2X1_LOC_602/Y AND2X1_LOC_600/a_8_24# 0.03fF
C49429 AND2X1_LOC_554/Y AND2X1_LOC_361/A 0.05fF
C49430 OR2X1_LOC_94/a_8_216# OR2X1_LOC_6/A 0.01fF
C49431 AND2X1_LOC_168/a_36_24# OR2X1_LOC_74/A 0.01fF
C49432 OR2X1_LOC_47/Y AND2X1_LOC_212/Y 0.37fF
C49433 AND2X1_LOC_303/A OR2X1_LOC_6/A 0.18fF
C49434 AND2X1_LOC_633/Y OR2X1_LOC_59/Y 0.02fF
C49435 AND2X1_LOC_356/a_36_24# OR2X1_LOC_43/A 0.00fF
C49436 OR2X1_LOC_92/a_8_216# AND2X1_LOC_243/Y 0.05fF
C49437 AND2X1_LOC_123/a_8_24# OR2X1_LOC_118/Y 0.11fF
C49438 OR2X1_LOC_158/A AND2X1_LOC_319/a_8_24# 0.06fF
C49439 AND2X1_LOC_17/Y AND2X1_LOC_47/a_8_24# 0.01fF
C49440 AND2X1_LOC_340/Y OR2X1_LOC_289/Y 0.35fF
C49441 OR2X1_LOC_427/A OR2X1_LOC_754/a_36_216# 0.00fF
C49442 OR2X1_LOC_830/a_8_216# AND2X1_LOC_47/Y 0.01fF
C49443 OR2X1_LOC_635/a_8_216# AND2X1_LOC_3/Y 0.01fF
C49444 OR2X1_LOC_516/B OR2X1_LOC_64/Y 0.02fF
C49445 OR2X1_LOC_271/B OR2X1_LOC_271/a_8_216# 0.06fF
C49446 OR2X1_LOC_501/B OR2X1_LOC_62/B 0.03fF
C49447 OR2X1_LOC_235/B AND2X1_LOC_672/B 0.01fF
C49448 AND2X1_LOC_576/Y OR2X1_LOC_36/Y 0.07fF
C49449 AND2X1_LOC_568/B AND2X1_LOC_864/a_8_24# 0.02fF
C49450 OR2X1_LOC_114/Y OR2X1_LOC_87/A 0.12fF
C49451 VDD OR2X1_LOC_218/Y 0.20fF
C49452 OR2X1_LOC_9/Y OR2X1_LOC_619/a_36_216# 0.00fF
C49453 OR2X1_LOC_160/B AND2X1_LOC_106/a_8_24# 0.04fF
C49454 D_INPUT_0 OR2X1_LOC_59/Y 0.10fF
C49455 AND2X1_LOC_702/a_8_24# OR2X1_LOC_3/Y 0.01fF
C49456 OR2X1_LOC_81/Y OR2X1_LOC_6/A 0.42fF
C49457 AND2X1_LOC_572/Y AND2X1_LOC_489/Y 0.10fF
C49458 INPUT_0 AND2X1_LOC_196/Y 0.02fF
C49459 OR2X1_LOC_87/A OR2X1_LOC_449/A 0.03fF
C49460 OR2X1_LOC_786/Y OR2X1_LOC_786/A 0.02fF
C49461 AND2X1_LOC_712/B OR2X1_LOC_422/a_8_216# 0.09fF
C49462 OR2X1_LOC_532/B OR2X1_LOC_778/a_8_216# 0.01fF
C49463 AND2X1_LOC_342/a_8_24# OR2X1_LOC_26/Y 0.07fF
C49464 OR2X1_LOC_814/A OR2X1_LOC_571/a_8_216# 0.01fF
C49465 AND2X1_LOC_84/a_36_24# OR2X1_LOC_69/A 0.00fF
C49466 OR2X1_LOC_476/B OR2X1_LOC_61/B 0.01fF
C49467 AND2X1_LOC_663/B OR2X1_LOC_427/A 0.07fF
C49468 OR2X1_LOC_43/A OR2X1_LOC_827/a_8_216# 0.05fF
C49469 OR2X1_LOC_502/A AND2X1_LOC_680/a_36_24# 0.01fF
C49470 AND2X1_LOC_359/a_8_24# AND2X1_LOC_363/A 0.01fF
C49471 OR2X1_LOC_690/a_8_216# OR2X1_LOC_585/A 0.01fF
C49472 AND2X1_LOC_136/a_8_24# AND2X1_LOC_43/B 0.01fF
C49473 AND2X1_LOC_858/B AND2X1_LOC_859/B 0.14fF
C49474 AND2X1_LOC_852/Y OR2X1_LOC_52/B 0.03fF
C49475 AND2X1_LOC_512/Y AND2X1_LOC_801/B 0.02fF
C49476 AND2X1_LOC_12/Y OR2X1_LOC_35/B 0.01fF
C49477 AND2X1_LOC_120/a_36_24# OR2X1_LOC_18/Y 0.00fF
C49478 OR2X1_LOC_486/a_8_216# OR2X1_LOC_739/A 0.01fF
C49479 AND2X1_LOC_65/A OR2X1_LOC_598/A 0.09fF
C49480 OR2X1_LOC_628/Y AND2X1_LOC_631/a_8_24# 0.03fF
C49481 OR2X1_LOC_485/A OR2X1_LOC_6/A 0.04fF
C49482 AND2X1_LOC_749/a_8_24# D_INPUT_0 0.05fF
C49483 AND2X1_LOC_569/A AND2X1_LOC_474/Y 0.12fF
C49484 OR2X1_LOC_663/A OR2X1_LOC_532/B 0.02fF
C49485 OR2X1_LOC_83/Y OR2X1_LOC_52/B 0.04fF
C49486 OR2X1_LOC_154/A OR2X1_LOC_624/B 1.02fF
C49487 AND2X1_LOC_367/A OR2X1_LOC_31/Y 0.03fF
C49488 OR2X1_LOC_695/a_8_216# AND2X1_LOC_687/B 0.01fF
C49489 AND2X1_LOC_70/Y OR2X1_LOC_112/B 0.04fF
C49490 AND2X1_LOC_366/a_8_24# OR2X1_LOC_47/Y 0.02fF
C49491 AND2X1_LOC_840/B OR2X1_LOC_74/A 0.10fF
C49492 OR2X1_LOC_427/A AND2X1_LOC_686/a_8_24# 0.02fF
C49493 OR2X1_LOC_191/B OR2X1_LOC_564/B 0.80fF
C49494 OR2X1_LOC_232/a_8_216# OR2X1_LOC_585/A 0.01fF
C49495 OR2X1_LOC_92/Y AND2X1_LOC_845/Y 0.17fF
C49496 OR2X1_LOC_74/A OR2X1_LOC_74/a_8_216# 0.04fF
C49497 OR2X1_LOC_87/A OR2X1_LOC_201/Y 0.04fF
C49498 VDD AND2X1_LOC_289/a_8_24# 0.00fF
C49499 AND2X1_LOC_624/B OR2X1_LOC_627/Y 0.73fF
C49500 AND2X1_LOC_91/B OR2X1_LOC_558/a_8_216# 0.04fF
C49501 OR2X1_LOC_792/Y OR2X1_LOC_286/a_8_216# 0.01fF
C49502 AND2X1_LOC_72/B OR2X1_LOC_66/A 0.03fF
C49503 OR2X1_LOC_287/B AND2X1_LOC_3/Y 0.04fF
C49504 OR2X1_LOC_479/Y OR2X1_LOC_778/Y 0.10fF
C49505 OR2X1_LOC_743/A OR2X1_LOC_423/a_8_216# 0.01fF
C49506 OR2X1_LOC_633/A OR2X1_LOC_80/A 1.43fF
C49507 OR2X1_LOC_46/A OR2X1_LOC_38/a_8_216# 0.01fF
C49508 AND2X1_LOC_702/Y AND2X1_LOC_324/a_8_24# 0.01fF
C49509 OR2X1_LOC_476/B AND2X1_LOC_291/a_8_24# 0.02fF
C49510 OR2X1_LOC_158/A OR2X1_LOC_72/Y 0.03fF
C49511 OR2X1_LOC_76/B OR2X1_LOC_532/B 0.06fF
C49512 AND2X1_LOC_487/a_8_24# OR2X1_LOC_814/A 0.09fF
C49513 AND2X1_LOC_70/Y OR2X1_LOC_66/Y 0.04fF
C49514 AND2X1_LOC_465/a_8_24# OR2X1_LOC_485/A 0.01fF
C49515 OR2X1_LOC_48/Y OR2X1_LOC_7/A 0.21fF
C49516 OR2X1_LOC_673/a_8_216# OR2X1_LOC_80/A -0.02fF
C49517 AND2X1_LOC_56/B AND2X1_LOC_27/a_8_24# 0.01fF
C49518 OR2X1_LOC_813/A OR2X1_LOC_18/Y 0.01fF
C49519 AND2X1_LOC_12/Y AND2X1_LOC_69/a_8_24# 0.01fF
C49520 OR2X1_LOC_97/B OR2X1_LOC_121/B 0.02fF
C49521 OR2X1_LOC_499/B D_INPUT_1 0.03fF
C49522 OR2X1_LOC_484/Y OR2X1_LOC_419/Y 0.10fF
C49523 AND2X1_LOC_34/a_8_24# OR2X1_LOC_27/Y 0.01fF
C49524 OR2X1_LOC_686/B AND2X1_LOC_31/Y 0.01fF
C49525 AND2X1_LOC_337/B AND2X1_LOC_798/Y 0.05fF
C49526 D_INPUT_5 OR2X1_LOC_51/B 0.01fF
C49527 OR2X1_LOC_444/a_8_216# OR2X1_LOC_87/A 0.01fF
C49528 VDD AND2X1_LOC_563/Y 0.38fF
C49529 OR2X1_LOC_744/A AND2X1_LOC_647/Y 0.03fF
C49530 AND2X1_LOC_486/Y OR2X1_LOC_437/a_8_216# 0.05fF
C49531 OR2X1_LOC_665/a_36_216# OR2X1_LOC_665/Y 0.01fF
C49532 AND2X1_LOC_472/B OR2X1_LOC_46/A 5.65fF
C49533 OR2X1_LOC_269/A OR2X1_LOC_549/A 0.02fF
C49534 OR2X1_LOC_22/Y AND2X1_LOC_361/A 0.07fF
C49535 D_INPUT_3 OR2X1_LOC_414/a_8_216# 0.07fF
C49536 OR2X1_LOC_659/a_8_216# AND2X1_LOC_47/Y 0.01fF
C49537 OR2X1_LOC_62/a_8_216# OR2X1_LOC_753/A 0.03fF
C49538 OR2X1_LOC_468/a_36_216# OR2X1_LOC_506/A 0.01fF
C49539 OR2X1_LOC_364/A OR2X1_LOC_532/B 0.08fF
C49540 AND2X1_LOC_517/a_8_24# AND2X1_LOC_88/Y 0.01fF
C49541 AND2X1_LOC_48/A OR2X1_LOC_219/B 5.36fF
C49542 OR2X1_LOC_437/A OR2X1_LOC_322/a_36_216# 0.14fF
C49543 OR2X1_LOC_185/Y OR2X1_LOC_532/B 11.79fF
C49544 INPUT_0 OR2X1_LOC_228/Y 0.07fF
C49545 OR2X1_LOC_624/A OR2X1_LOC_786/Y 0.10fF
C49546 AND2X1_LOC_392/A AND2X1_LOC_212/a_8_24# 0.04fF
C49547 OR2X1_LOC_137/Y OR2X1_LOC_244/A 0.00fF
C49548 AND2X1_LOC_319/A OR2X1_LOC_760/a_8_216# 0.01fF
C49549 OR2X1_LOC_87/A OR2X1_LOC_201/a_8_216# 0.03fF
C49550 AND2X1_LOC_784/A AND2X1_LOC_675/A 0.02fF
C49551 OR2X1_LOC_813/Y OR2X1_LOC_278/Y 0.38fF
C49552 OR2X1_LOC_160/A OR2X1_LOC_84/a_8_216# 0.04fF
C49553 OR2X1_LOC_405/A OR2X1_LOC_215/a_8_216# 0.09fF
C49554 OR2X1_LOC_600/A OR2X1_LOC_437/A 0.62fF
C49555 OR2X1_LOC_496/Y OR2X1_LOC_95/Y 0.00fF
C49556 AND2X1_LOC_580/B AND2X1_LOC_866/A 0.02fF
C49557 AND2X1_LOC_335/Y OR2X1_LOC_437/A 0.00fF
C49558 OR2X1_LOC_56/A OR2X1_LOC_384/Y 0.03fF
C49559 AND2X1_LOC_656/Y OR2X1_LOC_7/A 0.01fF
C49560 AND2X1_LOC_211/B AND2X1_LOC_170/B 0.00fF
C49561 OR2X1_LOC_709/a_8_216# OR2X1_LOC_308/Y 0.04fF
C49562 OR2X1_LOC_711/B OR2X1_LOC_469/B 0.01fF
C49563 AND2X1_LOC_303/A OR2X1_LOC_289/a_8_216# 0.03fF
C49564 AND2X1_LOC_456/Y OR2X1_LOC_31/Y 0.00fF
C49565 AND2X1_LOC_31/Y AND2X1_LOC_615/a_8_24# 0.03fF
C49566 OR2X1_LOC_612/Y OR2X1_LOC_71/A 0.05fF
C49567 OR2X1_LOC_70/Y D_INPUT_0 0.30fF
C49568 OR2X1_LOC_18/Y OR2X1_LOC_406/A 0.02fF
C49569 AND2X1_LOC_12/Y OR2X1_LOC_512/a_8_216# 0.01fF
C49570 OR2X1_LOC_31/Y OR2X1_LOC_74/A 0.36fF
C49571 OR2X1_LOC_696/A OR2X1_LOC_322/a_8_216# 0.05fF
C49572 AND2X1_LOC_86/Y OR2X1_LOC_398/a_8_216# 0.50fF
C49573 OR2X1_LOC_391/B D_INPUT_1 0.82fF
C49574 OR2X1_LOC_574/A OR2X1_LOC_276/B 0.10fF
C49575 OR2X1_LOC_36/Y OR2X1_LOC_29/a_8_216# 0.01fF
C49576 OR2X1_LOC_175/Y OR2X1_LOC_853/a_8_216# 0.01fF
C49577 OR2X1_LOC_87/A OR2X1_LOC_796/B 0.03fF
C49578 OR2X1_LOC_19/B OR2X1_LOC_46/A 0.25fF
C49579 AND2X1_LOC_671/a_8_24# OR2X1_LOC_54/Y 0.03fF
C49580 AND2X1_LOC_597/a_8_24# OR2X1_LOC_214/B 0.05fF
C49581 OR2X1_LOC_121/B OR2X1_LOC_814/A 0.10fF
C49582 AND2X1_LOC_686/a_8_24# AND2X1_LOC_687/B 0.04fF
C49583 AND2X1_LOC_334/a_8_24# AND2X1_LOC_634/Y 0.19fF
C49584 OR2X1_LOC_66/A AND2X1_LOC_36/Y 0.47fF
C49585 OR2X1_LOC_70/Y AND2X1_LOC_450/Y 0.01fF
C49586 OR2X1_LOC_841/B OR2X1_LOC_804/A 0.02fF
C49587 VDD OR2X1_LOC_703/Y 0.16fF
C49588 AND2X1_LOC_576/Y OR2X1_LOC_419/Y 0.02fF
C49589 OR2X1_LOC_841/A AND2X1_LOC_36/Y 0.00fF
C49590 AND2X1_LOC_92/Y OR2X1_LOC_723/B 0.03fF
C49591 OR2X1_LOC_116/a_8_216# OR2X1_LOC_66/Y 0.01fF
C49592 OR2X1_LOC_563/A OR2X1_LOC_161/B 0.18fF
C49593 AND2X1_LOC_40/Y OR2X1_LOC_71/A 0.03fF
C49594 OR2X1_LOC_661/a_36_216# OR2X1_LOC_68/B 0.00fF
C49595 OR2X1_LOC_269/B OR2X1_LOC_194/a_36_216# 0.02fF
C49596 OR2X1_LOC_22/A OR2X1_LOC_408/a_36_216# -0.00fF
C49597 AND2X1_LOC_600/a_8_24# OR2X1_LOC_602/B 0.01fF
C49598 AND2X1_LOC_632/a_8_24# OR2X1_LOC_615/Y 0.02fF
C49599 OR2X1_LOC_135/Y OR2X1_LOC_428/A 0.03fF
C49600 OR2X1_LOC_354/A OR2X1_LOC_788/B 0.01fF
C49601 AND2X1_LOC_22/Y OR2X1_LOC_549/A 0.07fF
C49602 OR2X1_LOC_696/A AND2X1_LOC_732/a_8_24# 0.02fF
C49603 OR2X1_LOC_186/Y OR2X1_LOC_336/a_8_216# 0.05fF
C49604 OR2X1_LOC_43/Y AND2X1_LOC_195/a_8_24# 0.23fF
C49605 OR2X1_LOC_378/Y OR2X1_LOC_378/a_8_216# 0.01fF
C49606 OR2X1_LOC_865/Y OR2X1_LOC_561/B 0.03fF
C49607 OR2X1_LOC_527/a_8_216# AND2X1_LOC_564/B 0.02fF
C49608 AND2X1_LOC_110/Y OR2X1_LOC_703/a_8_216# 0.01fF
C49609 AND2X1_LOC_834/a_8_24# AND2X1_LOC_796/A 0.12fF
C49610 OR2X1_LOC_804/B OR2X1_LOC_804/A 0.07fF
C49611 OR2X1_LOC_45/B AND2X1_LOC_476/Y 0.06fF
C49612 OR2X1_LOC_85/A AND2X1_LOC_215/a_8_24# 0.01fF
C49613 OR2X1_LOC_643/A OR2X1_LOC_68/B 0.03fF
C49614 OR2X1_LOC_589/A AND2X1_LOC_774/A 0.88fF
C49615 OR2X1_LOC_843/B OR2X1_LOC_343/a_36_216# 0.00fF
C49616 AND2X1_LOC_64/Y OR2X1_LOC_35/Y 0.03fF
C49617 OR2X1_LOC_160/Y OR2X1_LOC_162/a_8_216# 0.07fF
C49618 AND2X1_LOC_388/Y AND2X1_LOC_802/Y 0.82fF
C49619 OR2X1_LOC_375/A OR2X1_LOC_705/a_36_216# 0.00fF
C49620 OR2X1_LOC_118/a_8_216# OR2X1_LOC_131/a_8_216# 0.47fF
C49621 OR2X1_LOC_778/Y OR2X1_LOC_68/B 0.30fF
C49622 OR2X1_LOC_772/Y D_INPUT_1 0.01fF
C49623 OR2X1_LOC_620/Y OR2X1_LOC_532/Y 0.00fF
C49624 OR2X1_LOC_838/B OR2X1_LOC_46/A 0.06fF
C49625 OR2X1_LOC_846/A D_INPUT_1 0.06fF
C49626 AND2X1_LOC_469/Y AND2X1_LOC_212/Y 0.23fF
C49627 OR2X1_LOC_472/A OR2X1_LOC_68/B 0.00fF
C49628 OR2X1_LOC_64/Y AND2X1_LOC_845/a_8_24# 0.01fF
C49629 AND2X1_LOC_14/a_8_24# D_INPUT_0 0.02fF
C49630 AND2X1_LOC_98/a_8_24# OR2X1_LOC_428/A 0.01fF
C49631 OR2X1_LOC_19/B OR2X1_LOC_813/Y 0.06fF
C49632 OR2X1_LOC_255/a_8_216# OR2X1_LOC_47/Y 0.01fF
C49633 OR2X1_LOC_502/A OR2X1_LOC_354/a_8_216# 0.03fF
C49634 OR2X1_LOC_49/A VDD 0.69fF
C49635 OR2X1_LOC_160/B OR2X1_LOC_489/A 0.03fF
C49636 AND2X1_LOC_851/B OR2X1_LOC_95/Y 0.12fF
C49637 OR2X1_LOC_647/A OR2X1_LOC_68/B 0.04fF
C49638 AND2X1_LOC_454/a_36_24# OR2X1_LOC_428/A 0.00fF
C49639 AND2X1_LOC_182/A OR2X1_LOC_40/Y 0.06fF
C49640 OR2X1_LOC_113/Y AND2X1_LOC_22/Y 0.06fF
C49641 OR2X1_LOC_739/A OR2X1_LOC_308/Y 0.03fF
C49642 OR2X1_LOC_337/a_8_216# OR2X1_LOC_352/a_8_216# 0.47fF
C49643 OR2X1_LOC_40/Y AND2X1_LOC_469/a_36_24# 0.01fF
C49644 AND2X1_LOC_641/a_8_24# D_INPUT_0 0.02fF
C49645 OR2X1_LOC_833/Y AND2X1_LOC_70/Y 0.01fF
C49646 VDD OR2X1_LOC_596/A 0.41fF
C49647 AND2X1_LOC_810/A OR2X1_LOC_744/A 0.05fF
C49648 AND2X1_LOC_712/Y VDD 0.21fF
C49649 OR2X1_LOC_160/B OR2X1_LOC_772/A 0.01fF
C49650 OR2X1_LOC_850/B OR2X1_LOC_366/B 0.01fF
C49651 OR2X1_LOC_84/B OR2X1_LOC_771/B 0.07fF
C49652 OR2X1_LOC_114/Y OR2X1_LOC_844/B 0.00fF
C49653 OR2X1_LOC_287/B OR2X1_LOC_576/a_8_216# 0.01fF
C49654 OR2X1_LOC_505/Y AND2X1_LOC_508/B 0.01fF
C49655 OR2X1_LOC_409/Y OR2X1_LOC_588/A 0.19fF
C49656 OR2X1_LOC_244/A OR2X1_LOC_398/a_8_216# 0.03fF
C49657 AND2X1_LOC_421/a_8_24# AND2X1_LOC_44/Y 0.01fF
C49658 VDD OR2X1_LOC_526/Y 0.31fF
C49659 OR2X1_LOC_244/B OR2X1_LOC_549/A 0.03fF
C49660 AND2X1_LOC_212/A AND2X1_LOC_364/Y 0.59fF
C49661 OR2X1_LOC_756/B AND2X1_LOC_83/a_8_24# 0.02fF
C49662 OR2X1_LOC_269/B OR2X1_LOC_308/Y 0.08fF
C49663 OR2X1_LOC_372/a_8_216# OR2X1_LOC_437/A 0.18fF
C49664 OR2X1_LOC_679/a_8_216# OR2X1_LOC_679/Y 0.01fF
C49665 AND2X1_LOC_70/Y AND2X1_LOC_387/a_8_24# 0.01fF
C49666 AND2X1_LOC_566/B AND2X1_LOC_365/a_8_24# 0.01fF
C49667 D_INPUT_0 AND2X1_LOC_31/Y 0.59fF
C49668 AND2X1_LOC_508/B AND2X1_LOC_658/A 0.03fF
C49669 OR2X1_LOC_175/Y OR2X1_LOC_185/A 0.07fF
C49670 AND2X1_LOC_321/a_8_24# AND2X1_LOC_44/Y 0.02fF
C49671 AND2X1_LOC_340/a_8_24# OR2X1_LOC_744/A 0.01fF
C49672 OR2X1_LOC_744/A AND2X1_LOC_860/A 0.07fF
C49673 OR2X1_LOC_715/B AND2X1_LOC_41/A 0.03fF
C49674 AND2X1_LOC_334/Y AND2X1_LOC_338/a_8_24# 0.03fF
C49675 OR2X1_LOC_259/a_8_216# AND2X1_LOC_44/Y 0.01fF
C49676 OR2X1_LOC_231/B OR2X1_LOC_231/A 0.16fF
C49677 AND2X1_LOC_711/A OR2X1_LOC_59/Y 0.31fF
C49678 INPUT_0 OR2X1_LOC_14/a_8_216# 0.01fF
C49679 OR2X1_LOC_91/Y AND2X1_LOC_465/A 0.07fF
C49680 OR2X1_LOC_51/Y OR2X1_LOC_743/a_8_216# 0.01fF
C49681 AND2X1_LOC_392/A AND2X1_LOC_392/a_8_24# 0.05fF
C49682 OR2X1_LOC_691/Y OR2X1_LOC_185/A 0.23fF
C49683 AND2X1_LOC_567/a_36_24# OR2X1_LOC_744/A 0.01fF
C49684 VDD OR2X1_LOC_310/Y 0.04fF
C49685 OR2X1_LOC_505/a_8_216# OR2X1_LOC_18/Y 0.02fF
C49686 OR2X1_LOC_325/Y OR2X1_LOC_326/a_8_216# 0.39fF
C49687 AND2X1_LOC_776/a_36_24# OR2X1_LOC_56/A 0.00fF
C49688 OR2X1_LOC_118/a_8_216# AND2X1_LOC_573/A 0.06fF
C49689 AND2X1_LOC_848/Y OR2X1_LOC_428/A 0.03fF
C49690 OR2X1_LOC_91/A OR2X1_LOC_56/A 0.85fF
C49691 OR2X1_LOC_756/B OR2X1_LOC_602/Y 0.01fF
C49692 VDD OR2X1_LOC_808/A 0.27fF
C49693 OR2X1_LOC_185/Y OR2X1_LOC_392/a_36_216# 0.00fF
C49694 OR2X1_LOC_526/Y OR2X1_LOC_677/Y 0.44fF
C49695 OR2X1_LOC_160/A OR2X1_LOC_435/A 0.03fF
C49696 OR2X1_LOC_78/B AND2X1_LOC_232/a_8_24# -0.00fF
C49697 OR2X1_LOC_659/A OR2X1_LOC_244/Y 0.36fF
C49698 OR2X1_LOC_631/A OR2X1_LOC_575/A 0.10fF
C49699 OR2X1_LOC_231/B OR2X1_LOC_130/A 0.02fF
C49700 OR2X1_LOC_139/A OR2X1_LOC_659/B -0.02fF
C49701 OR2X1_LOC_859/A OR2X1_LOC_571/Y 0.11fF
C49702 OR2X1_LOC_7/A AND2X1_LOC_772/Y 0.19fF
C49703 AND2X1_LOC_711/a_36_24# OR2X1_LOC_59/Y 0.00fF
C49704 OR2X1_LOC_36/Y AND2X1_LOC_244/A 0.03fF
C49705 OR2X1_LOC_756/B AND2X1_LOC_179/a_36_24# 0.01fF
C49706 AND2X1_LOC_454/Y OR2X1_LOC_421/Y 0.01fF
C49707 AND2X1_LOC_588/B AND2X1_LOC_21/Y 0.04fF
C49708 VDD OR2X1_LOC_422/Y 0.04fF
C49709 OR2X1_LOC_485/A OR2X1_LOC_184/a_8_216# 0.02fF
C49710 AND2X1_LOC_91/B AND2X1_LOC_38/a_8_24# 0.01fF
C49711 OR2X1_LOC_96/B OR2X1_LOC_9/a_8_216# 0.00fF
C49712 OR2X1_LOC_36/Y OR2X1_LOC_16/A 1.45fF
C49713 OR2X1_LOC_18/Y AND2X1_LOC_606/a_8_24# 0.01fF
C49714 AND2X1_LOC_95/Y AND2X1_LOC_411/a_8_24# 0.13fF
C49715 AND2X1_LOC_565/B OR2X1_LOC_427/A 0.01fF
C49716 AND2X1_LOC_91/B OR2X1_LOC_479/Y 0.19fF
C49717 VDD AND2X1_LOC_805/Y 0.36fF
C49718 OR2X1_LOC_43/A AND2X1_LOC_774/A 0.10fF
C49719 AND2X1_LOC_654/B AND2X1_LOC_434/a_8_24# 0.09fF
C49720 OR2X1_LOC_519/a_8_216# VDD 0.21fF
C49721 VDD OR2X1_LOC_732/a_8_216# 0.21fF
C49722 AND2X1_LOC_706/Y OR2X1_LOC_44/Y 0.03fF
C49723 OR2X1_LOC_53/Y OR2X1_LOC_3/Y 0.04fF
C49724 OR2X1_LOC_141/B OR2X1_LOC_572/a_36_216# 0.00fF
C49725 OR2X1_LOC_154/A OR2X1_LOC_768/a_8_216# 0.04fF
C49726 OR2X1_LOC_26/Y OR2X1_LOC_12/Y 0.33fF
C49727 AND2X1_LOC_539/Y OR2X1_LOC_70/Y 0.79fF
C49728 AND2X1_LOC_578/A AND2X1_LOC_242/B 0.01fF
C49729 OR2X1_LOC_564/A OR2X1_LOC_564/a_8_216# 0.01fF
C49730 OR2X1_LOC_677/a_8_216# OR2X1_LOC_441/Y 0.06fF
C49731 AND2X1_LOC_715/A OR2X1_LOC_619/Y 0.07fF
C49732 VDD OR2X1_LOC_433/Y 0.20fF
C49733 OR2X1_LOC_509/A OR2X1_LOC_78/B 0.02fF
C49734 AND2X1_LOC_503/a_36_24# OR2X1_LOC_78/A 0.00fF
C49735 AND2X1_LOC_366/a_8_24# OR2X1_LOC_625/Y 0.04fF
C49736 OR2X1_LOC_575/A OR2X1_LOC_632/Y 0.40fF
C49737 AND2X1_LOC_840/A OR2X1_LOC_59/Y 0.03fF
C49738 OR2X1_LOC_262/Y AND2X1_LOC_249/a_36_24# 0.00fF
C49739 OR2X1_LOC_482/a_36_216# AND2X1_LOC_859/Y 0.01fF
C49740 AND2X1_LOC_95/Y OR2X1_LOC_360/a_8_216# 0.01fF
C49741 OR2X1_LOC_744/A OR2X1_LOC_432/a_8_216# 0.01fF
C49742 OR2X1_LOC_190/A OR2X1_LOC_456/a_36_216# 0.01fF
C49743 OR2X1_LOC_204/Y OR2X1_LOC_786/A 0.00fF
C49744 AND2X1_LOC_349/B OR2X1_LOC_12/Y 0.00fF
C49745 AND2X1_LOC_51/a_8_24# D_INPUT_4 0.16fF
C49746 OR2X1_LOC_89/A OR2X1_LOC_12/Y 3.67fF
C49747 VDD OR2X1_LOC_575/a_8_216# 0.00fF
C49748 OR2X1_LOC_502/A OR2X1_LOC_307/B 0.04fF
C49749 OR2X1_LOC_74/A AND2X1_LOC_213/B 0.03fF
C49750 AND2X1_LOC_509/a_8_24# AND2X1_LOC_573/A 0.01fF
C49751 AND2X1_LOC_858/B AND2X1_LOC_850/Y 0.02fF
C49752 OR2X1_LOC_709/A OR2X1_LOC_574/A 0.05fF
C49753 AND2X1_LOC_573/A OR2X1_LOC_56/A 0.02fF
C49754 VDD OR2X1_LOC_463/B 0.12fF
C49755 AND2X1_LOC_449/Y AND2X1_LOC_454/a_8_24# 0.20fF
C49756 AND2X1_LOC_683/a_36_24# OR2X1_LOC_161/B 0.00fF
C49757 AND2X1_LOC_366/A OR2X1_LOC_427/A 0.44fF
C49758 OR2X1_LOC_744/A AND2X1_LOC_400/a_8_24# 0.02fF
C49759 OR2X1_LOC_375/A OR2X1_LOC_741/Y 0.05fF
C49760 OR2X1_LOC_64/Y OR2X1_LOC_321/a_8_216# 0.01fF
C49761 OR2X1_LOC_659/Y OR2X1_LOC_557/A 0.00fF
C49762 OR2X1_LOC_604/A AND2X1_LOC_576/Y 0.10fF
C49763 AND2X1_LOC_799/a_8_24# OR2X1_LOC_417/Y 0.03fF
C49764 OR2X1_LOC_7/A OR2X1_LOC_584/a_36_216# 0.02fF
C49765 OR2X1_LOC_108/Y OR2X1_LOC_36/Y 0.13fF
C49766 AND2X1_LOC_350/B OR2X1_LOC_70/Y 0.03fF
C49767 OR2X1_LOC_40/Y AND2X1_LOC_580/B 0.05fF
C49768 OR2X1_LOC_58/Y OR2X1_LOC_44/Y 0.03fF
C49769 AND2X1_LOC_64/Y AND2X1_LOC_667/a_8_24# 0.11fF
C49770 OR2X1_LOC_45/B OR2X1_LOC_431/a_8_216# 0.01fF
C49771 AND2X1_LOC_542/a_8_24# OR2X1_LOC_280/Y 0.03fF
C49772 AND2X1_LOC_563/A AND2X1_LOC_560/B 0.01fF
C49773 VDD OR2X1_LOC_87/B 0.31fF
C49774 AND2X1_LOC_191/B AND2X1_LOC_859/a_8_24# 0.03fF
C49775 OR2X1_LOC_40/Y OR2X1_LOC_612/B 0.03fF
C49776 OR2X1_LOC_114/B AND2X1_LOC_292/a_8_24# 0.05fF
C49777 OR2X1_LOC_235/B OR2X1_LOC_377/A 0.07fF
C49778 AND2X1_LOC_509/Y AND2X1_LOC_624/A 0.03fF
C49779 VDD AND2X1_LOC_661/A 0.42fF
C49780 AND2X1_LOC_510/a_8_24# AND2X1_LOC_621/Y 0.02fF
C49781 OR2X1_LOC_325/A OR2X1_LOC_620/Y 0.02fF
C49782 OR2X1_LOC_600/A OR2X1_LOC_753/A 0.14fF
C49783 AND2X1_LOC_856/B OR2X1_LOC_428/A 0.08fF
C49784 OR2X1_LOC_375/A AND2X1_LOC_232/a_8_24# 0.14fF
C49785 OR2X1_LOC_84/A AND2X1_LOC_36/Y 0.01fF
C49786 OR2X1_LOC_97/A OR2X1_LOC_476/B 0.02fF
C49787 OR2X1_LOC_327/a_8_216# OR2X1_LOC_502/A 0.05fF
C49788 OR2X1_LOC_479/Y OR2X1_LOC_364/a_8_216# 0.02fF
C49789 AND2X1_LOC_350/B AND2X1_LOC_333/a_8_24# 0.11fF
C49790 AND2X1_LOC_12/Y AND2X1_LOC_65/a_8_24# 0.01fF
C49791 AND2X1_LOC_863/A OR2X1_LOC_428/A 0.03fF
C49792 OR2X1_LOC_695/Y OR2X1_LOC_52/B 0.01fF
C49793 OR2X1_LOC_97/A OR2X1_LOC_650/Y 0.03fF
C49794 AND2X1_LOC_167/a_36_24# OR2X1_LOC_161/A 0.01fF
C49795 VDD AND2X1_LOC_612/B 0.01fF
C49796 AND2X1_LOC_668/a_36_24# OR2X1_LOC_59/Y 0.00fF
C49797 OR2X1_LOC_160/B AND2X1_LOC_3/Y 1.18fF
C49798 OR2X1_LOC_108/Y AND2X1_LOC_493/a_36_24# 0.00fF
C49799 OR2X1_LOC_8/Y AND2X1_LOC_838/a_36_24# -0.00fF
C49800 OR2X1_LOC_771/a_8_216# OR2X1_LOC_771/B 0.08fF
C49801 OR2X1_LOC_70/Y OR2X1_LOC_131/A 0.31fF
C49802 VDD AND2X1_LOC_259/Y 0.21fF
C49803 OR2X1_LOC_235/B OR2X1_LOC_85/A 0.01fF
C49804 OR2X1_LOC_186/Y AND2X1_LOC_680/a_8_24# 0.11fF
C49805 OR2X1_LOC_185/Y OR2X1_LOC_624/Y 0.02fF
C49806 OR2X1_LOC_648/A OR2X1_LOC_810/A 0.07fF
C49807 OR2X1_LOC_158/A AND2X1_LOC_326/A 0.15fF
C49808 AND2X1_LOC_70/Y OR2X1_LOC_574/A 0.04fF
C49809 OR2X1_LOC_250/a_8_216# OR2X1_LOC_278/Y 0.01fF
C49810 AND2X1_LOC_160/Y OR2X1_LOC_7/A 0.03fF
C49811 AND2X1_LOC_729/Y OR2X1_LOC_92/Y 0.23fF
C49812 VDD OR2X1_LOC_33/B 0.00fF
C49813 OR2X1_LOC_208/a_36_216# OR2X1_LOC_35/Y 0.03fF
C49814 AND2X1_LOC_81/B OR2X1_LOC_474/Y 0.03fF
C49815 INPUT_0 AND2X1_LOC_856/A 0.02fF
C49816 AND2X1_LOC_711/Y AND2X1_LOC_711/A 0.00fF
C49817 OR2X1_LOC_154/A OR2X1_LOC_400/a_8_216# 0.06fF
C49818 AND2X1_LOC_512/a_8_24# INPUT_0 0.03fF
C49819 AND2X1_LOC_12/Y OR2X1_LOC_231/A 0.00fF
C49820 OR2X1_LOC_391/B OR2X1_LOC_391/a_8_216# 0.06fF
C49821 OR2X1_LOC_287/B INPUT_0 0.16fF
C49822 AND2X1_LOC_490/a_8_24# OR2X1_LOC_78/B 0.01fF
C49823 OR2X1_LOC_613/Y AND2X1_LOC_866/B 0.03fF
C49824 OR2X1_LOC_421/A OR2X1_LOC_64/Y 0.09fF
C49825 OR2X1_LOC_616/Y AND2X1_LOC_805/Y 0.01fF
C49826 OR2X1_LOC_40/Y OR2X1_LOC_295/a_8_216# 0.01fF
C49827 AND2X1_LOC_40/Y OR2X1_LOC_593/a_8_216# 0.01fF
C49828 OR2X1_LOC_48/B AND2X1_LOC_435/a_36_24# 0.01fF
C49829 AND2X1_LOC_784/A OR2X1_LOC_92/Y 0.07fF
C49830 OR2X1_LOC_516/A AND2X1_LOC_468/B 0.14fF
C49831 AND2X1_LOC_847/Y AND2X1_LOC_848/a_8_24# 0.01fF
C49832 AND2X1_LOC_554/Y AND2X1_LOC_572/Y 0.17fF
C49833 AND2X1_LOC_47/Y AND2X1_LOC_433/a_8_24# 0.01fF
C49834 AND2X1_LOC_866/A AND2X1_LOC_455/B 0.07fF
C49835 OR2X1_LOC_19/B INPUT_2 0.00fF
C49836 OR2X1_LOC_473/A AND2X1_LOC_7/B 0.05fF
C49837 OR2X1_LOC_387/A OR2X1_LOC_387/a_8_216# 0.01fF
C49838 OR2X1_LOC_324/A AND2X1_LOC_56/B 0.10fF
C49839 OR2X1_LOC_154/A OR2X1_LOC_447/A 0.02fF
C49840 AND2X1_LOC_339/B OR2X1_LOC_111/Y 0.01fF
C49841 AND2X1_LOC_448/Y AND2X1_LOC_453/a_8_24# 0.03fF
C49842 OR2X1_LOC_19/B AND2X1_LOC_403/a_8_24# 0.05fF
C49843 AND2X1_LOC_702/Y OR2X1_LOC_48/B 0.04fF
C49844 AND2X1_LOC_857/Y OR2X1_LOC_299/a_36_216# 0.00fF
C49845 OR2X1_LOC_656/B OR2X1_LOC_216/Y 0.10fF
C49846 OR2X1_LOC_70/Y AND2X1_LOC_471/Y 2.84fF
C49847 AND2X1_LOC_12/Y OR2X1_LOC_130/A 0.07fF
C49848 OR2X1_LOC_114/B OR2X1_LOC_62/B 0.06fF
C49849 AND2X1_LOC_719/Y OR2X1_LOC_71/Y 0.05fF
C49850 OR2X1_LOC_687/Y OR2X1_LOC_161/A 0.15fF
C49851 OR2X1_LOC_728/A OR2X1_LOC_728/a_8_216# 0.47fF
C49852 OR2X1_LOC_860/Y OR2X1_LOC_287/B 0.01fF
C49853 OR2X1_LOC_318/A OR2X1_LOC_223/A 0.00fF
C49854 AND2X1_LOC_794/B AND2X1_LOC_810/Y 0.07fF
C49855 OR2X1_LOC_91/Y OR2X1_LOC_237/Y 0.06fF
C49856 AND2X1_LOC_61/Y OR2X1_LOC_22/Y 0.08fF
C49857 OR2X1_LOC_241/B OR2X1_LOC_121/A 0.03fF
C49858 OR2X1_LOC_144/Y OR2X1_LOC_74/A 0.07fF
C49859 AND2X1_LOC_393/a_8_24# OR2X1_LOC_377/A 0.03fF
C49860 OR2X1_LOC_26/Y OR2X1_LOC_393/Y 0.05fF
C49861 OR2X1_LOC_151/Y OR2X1_LOC_739/A 0.21fF
C49862 OR2X1_LOC_414/a_8_216# OR2X1_LOC_83/A 0.01fF
C49863 OR2X1_LOC_458/B AND2X1_LOC_674/a_8_24# 0.01fF
C49864 OR2X1_LOC_619/Y OR2X1_LOC_753/A 0.07fF
C49865 OR2X1_LOC_83/Y OR2X1_LOC_394/Y 0.01fF
C49866 AND2X1_LOC_658/A OR2X1_LOC_815/A 0.04fF
C49867 OR2X1_LOC_600/A AND2X1_LOC_845/Y 0.07fF
C49868 OR2X1_LOC_6/B AND2X1_LOC_28/a_36_24# 0.01fF
C49869 AND2X1_LOC_81/B OR2X1_LOC_217/Y 0.03fF
C49870 AND2X1_LOC_41/a_36_24# AND2X1_LOC_53/Y 0.01fF
C49871 OR2X1_LOC_2/a_8_216# INPUT_7 0.01fF
C49872 AND2X1_LOC_456/B OR2X1_LOC_64/Y 0.02fF
C49873 OR2X1_LOC_329/B AND2X1_LOC_116/B 0.02fF
C49874 AND2X1_LOC_364/Y AND2X1_LOC_727/A 0.03fF
C49875 AND2X1_LOC_544/a_36_24# OR2X1_LOC_70/Y 0.00fF
C49876 OR2X1_LOC_151/A OR2X1_LOC_223/A 0.03fF
C49877 OR2X1_LOC_467/A OR2X1_LOC_447/Y 0.00fF
C49878 VDD OR2X1_LOC_223/a_8_216# 0.00fF
C49879 AND2X1_LOC_718/a_36_24# OR2X1_LOC_64/Y 0.00fF
C49880 OR2X1_LOC_566/A OR2X1_LOC_170/Y 0.17fF
C49881 OR2X1_LOC_419/Y AND2X1_LOC_244/A 0.01fF
C49882 OR2X1_LOC_54/Y OR2X1_LOC_234/Y -0.01fF
C49883 OR2X1_LOC_419/a_8_216# OR2X1_LOC_12/Y 0.01fF
C49884 OR2X1_LOC_489/B OR2X1_LOC_287/B -0.00fF
C49885 OR2X1_LOC_214/A OR2X1_LOC_228/Y 0.10fF
C49886 OR2X1_LOC_485/A OR2X1_LOC_45/a_8_216# 0.01fF
C49887 OR2X1_LOC_219/B OR2X1_LOC_350/a_8_216# 0.00fF
C49888 OR2X1_LOC_81/Y OR2X1_LOC_44/Y 0.06fF
C49889 AND2X1_LOC_147/Y AND2X1_LOC_624/A 0.15fF
C49890 AND2X1_LOC_91/B OR2X1_LOC_68/B 0.31fF
C49891 OR2X1_LOC_40/Y AND2X1_LOC_803/a_8_24# 0.04fF
C49892 OR2X1_LOC_861/a_8_216# AND2X1_LOC_51/Y 0.01fF
C49893 OR2X1_LOC_26/Y AND2X1_LOC_650/Y 0.06fF
C49894 AND2X1_LOC_589/a_36_24# OR2X1_LOC_799/A 0.00fF
C49895 OR2X1_LOC_70/Y AND2X1_LOC_450/a_36_24# 0.00fF
C49896 AND2X1_LOC_7/B OR2X1_LOC_228/Y 0.09fF
C49897 VDD OR2X1_LOC_760/Y 0.00fF
C49898 OR2X1_LOC_696/A AND2X1_LOC_592/a_8_24# 0.04fF
C49899 OR2X1_LOC_830/a_8_216# OR2X1_LOC_284/B 0.47fF
C49900 AND2X1_LOC_64/Y AND2X1_LOC_419/a_8_24# 0.00fF
C49901 OR2X1_LOC_827/Y OR2X1_LOC_6/A 0.01fF
C49902 AND2X1_LOC_474/Y OR2X1_LOC_44/Y 0.01fF
C49903 OR2X1_LOC_269/Y OR2X1_LOC_66/A 0.09fF
C49904 AND2X1_LOC_7/B OR2X1_LOC_513/Y 0.01fF
C49905 OR2X1_LOC_437/Y AND2X1_LOC_784/a_8_24# 0.23fF
C49906 AND2X1_LOC_517/a_8_24# OR2X1_LOC_121/B 0.01fF
C49907 OR2X1_LOC_476/B AND2X1_LOC_290/a_8_24# 0.02fF
C49908 OR2X1_LOC_674/a_8_216# OR2X1_LOC_95/Y 0.01fF
C49909 AND2X1_LOC_456/B OR2X1_LOC_417/A 0.07fF
C49910 OR2X1_LOC_485/A OR2X1_LOC_44/Y 0.37fF
C49911 OR2X1_LOC_151/A OR2X1_LOC_705/B 0.03fF
C49912 OR2X1_LOC_168/Y OR2X1_LOC_777/B 0.19fF
C49913 AND2X1_LOC_213/B AND2X1_LOC_783/a_8_24# 0.01fF
C49914 GATE_366 OR2X1_LOC_258/Y 0.03fF
C49915 OR2X1_LOC_273/a_8_216# OR2X1_LOC_36/Y 0.03fF
C49916 OR2X1_LOC_108/Y OR2X1_LOC_419/Y 0.10fF
C49917 OR2X1_LOC_161/B OR2X1_LOC_724/A 0.07fF
C49918 OR2X1_LOC_427/A AND2X1_LOC_635/a_36_24# 0.00fF
C49919 VDD AND2X1_LOC_797/B 0.13fF
C49920 OR2X1_LOC_687/Y AND2X1_LOC_51/Y 0.03fF
C49921 OR2X1_LOC_272/Y OR2X1_LOC_26/Y 0.02fF
C49922 VDD OR2X1_LOC_374/Y 0.10fF
C49923 OR2X1_LOC_275/A AND2X1_LOC_264/a_8_24# 0.01fF
C49924 OR2X1_LOC_676/Y AND2X1_LOC_699/a_8_24# -0.05fF
C49925 AND2X1_LOC_12/Y OR2X1_LOC_62/B 0.03fF
C49926 OR2X1_LOC_161/B OR2X1_LOC_365/a_36_216# 0.00fF
C49927 OR2X1_LOC_426/B OR2X1_LOC_86/A 0.03fF
C49928 OR2X1_LOC_305/a_8_216# AND2X1_LOC_307/Y 0.03fF
C49929 AND2X1_LOC_621/Y AND2X1_LOC_678/a_8_24# 0.10fF
C49930 OR2X1_LOC_296/Y OR2X1_LOC_629/A 0.00fF
C49931 AND2X1_LOC_716/Y AND2X1_LOC_318/Y 0.02fF
C49932 OR2X1_LOC_164/Y OR2X1_LOC_47/Y 0.06fF
C49933 OR2X1_LOC_272/Y OR2X1_LOC_89/A 0.35fF
C49934 AND2X1_LOC_17/Y OR2X1_LOC_636/a_36_216# 0.02fF
C49935 AND2X1_LOC_540/a_8_24# OR2X1_LOC_47/Y 0.17fF
C49936 OR2X1_LOC_771/B OR2X1_LOC_338/A 0.07fF
C49937 OR2X1_LOC_168/B OR2X1_LOC_804/A 0.07fF
C49938 OR2X1_LOC_405/A AND2X1_LOC_47/Y 0.10fF
C49939 AND2X1_LOC_866/A OR2X1_LOC_278/Y 0.03fF
C49940 AND2X1_LOC_11/Y OR2X1_LOC_651/A 0.00fF
C49941 AND2X1_LOC_841/a_8_24# AND2X1_LOC_841/B 0.09fF
C49942 OR2X1_LOC_19/B OR2X1_LOC_269/B 0.08fF
C49943 OR2X1_LOC_287/B OR2X1_LOC_401/A 0.01fF
C49944 OR2X1_LOC_468/A OR2X1_LOC_854/A 0.00fF
C49945 OR2X1_LOC_62/B OR2X1_LOC_266/a_36_216# 0.00fF
C49946 INPUT_0 OR2X1_LOC_28/a_8_216# 0.01fF
C49947 OR2X1_LOC_221/a_8_216# AND2X1_LOC_47/Y 0.05fF
C49948 INPUT_5 OR2X1_LOC_31/a_8_216# 0.01fF
C49949 AND2X1_LOC_462/a_8_24# OR2X1_LOC_753/A 0.18fF
C49950 OR2X1_LOC_64/Y AND2X1_LOC_717/B 0.06fF
C49951 OR2X1_LOC_36/Y AND2X1_LOC_687/Y 0.03fF
C49952 OR2X1_LOC_32/Y OR2X1_LOC_416/Y 0.02fF
C49953 OR2X1_LOC_538/A OR2X1_LOC_365/B 1.62fF
C49954 OR2X1_LOC_22/Y AND2X1_LOC_852/Y 0.07fF
C49955 OR2X1_LOC_223/B OR2X1_LOC_223/a_8_216# 0.05fF
C49956 OR2X1_LOC_707/B OR2X1_LOC_87/A 0.15fF
C49957 OR2X1_LOC_678/Y AND2X1_LOC_679/a_8_24# 0.10fF
C49958 OR2X1_LOC_599/A AND2X1_LOC_800/a_8_24# 0.00fF
C49959 OR2X1_LOC_474/Y OR2X1_LOC_66/Y 0.03fF
C49960 OR2X1_LOC_864/A D_INPUT_0 0.10fF
C49961 OR2X1_LOC_537/a_8_216# OR2X1_LOC_390/A 0.01fF
C49962 OR2X1_LOC_647/a_36_216# OR2X1_LOC_647/B 0.00fF
C49963 AND2X1_LOC_64/Y OR2X1_LOC_115/B 1.34fF
C49964 AND2X1_LOC_729/B AND2X1_LOC_855/a_8_24# 0.05fF
C49965 AND2X1_LOC_624/B AND2X1_LOC_805/Y 0.18fF
C49966 OR2X1_LOC_849/A AND2X1_LOC_15/a_36_24# 0.00fF
C49967 OR2X1_LOC_87/A OR2X1_LOC_440/A 0.03fF
C49968 OR2X1_LOC_473/A OR2X1_LOC_805/A 0.02fF
C49969 OR2X1_LOC_62/B AND2X1_LOC_79/Y 0.03fF
C49970 OR2X1_LOC_95/Y OR2X1_LOC_372/Y 0.02fF
C49971 INPUT_1 AND2X1_LOC_234/a_36_24# 0.00fF
C49972 D_INPUT_0 OR2X1_LOC_240/A 0.01fF
C49973 OR2X1_LOC_691/a_8_216# AND2X1_LOC_36/Y 0.06fF
C49974 OR2X1_LOC_633/B D_INPUT_0 0.03fF
C49975 OR2X1_LOC_160/A OR2X1_LOC_783/a_8_216# 0.02fF
C49976 OR2X1_LOC_276/B OR2X1_LOC_203/Y 0.04fF
C49977 OR2X1_LOC_409/B OR2X1_LOC_588/Y 0.81fF
C49978 OR2X1_LOC_244/A AND2X1_LOC_3/Y 0.07fF
C49979 OR2X1_LOC_654/A OR2X1_LOC_532/B 0.08fF
C49980 OR2X1_LOC_270/Y OR2X1_LOC_553/A 0.07fF
C49981 OR2X1_LOC_3/Y INPUT_1 1.38fF
C49982 AND2X1_LOC_12/Y AND2X1_LOC_39/Y 0.01fF
C49983 AND2X1_LOC_717/B OR2X1_LOC_417/A 4.05fF
C49984 OR2X1_LOC_359/a_8_216# OR2X1_LOC_580/A 0.04fF
C49985 INPUT_4 OR2X1_LOC_2/a_8_216# 0.05fF
C49986 OR2X1_LOC_726/A OR2X1_LOC_209/A 0.12fF
C49987 AND2X1_LOC_40/Y AND2X1_LOC_31/Y 0.17fF
C49988 AND2X1_LOC_59/Y OR2X1_LOC_804/A 0.34fF
C49989 OR2X1_LOC_92/Y OR2X1_LOC_88/Y 0.06fF
C49990 OR2X1_LOC_73/a_8_216# OR2X1_LOC_95/Y 0.01fF
C49991 OR2X1_LOC_78/A OR2X1_LOC_366/Y 0.03fF
C49992 OR2X1_LOC_856/a_36_216# OR2X1_LOC_532/B 0.00fF
C49993 OR2X1_LOC_405/A OR2X1_LOC_717/a_36_216# 0.00fF
C49994 OR2X1_LOC_116/A OR2X1_LOC_66/Y 0.01fF
C49995 OR2X1_LOC_12/Y AND2X1_LOC_590/a_8_24# 0.04fF
C49996 OR2X1_LOC_188/Y OR2X1_LOC_121/A 0.01fF
C49997 OR2X1_LOC_318/Y OR2X1_LOC_228/Y 0.02fF
C49998 AND2X1_LOC_95/Y OR2X1_LOC_543/a_8_216# 0.01fF
C49999 AND2X1_LOC_721/A OR2X1_LOC_85/A 0.00fF
C50000 OR2X1_LOC_191/B OR2X1_LOC_223/A 0.02fF
C50001 OR2X1_LOC_116/a_36_216# OR2X1_LOC_786/Y 0.00fF
C50002 AND2X1_LOC_12/Y OR2X1_LOC_365/B 0.03fF
C50003 AND2X1_LOC_580/A AND2X1_LOC_793/Y 0.07fF
C50004 OR2X1_LOC_87/A OR2X1_LOC_446/A 0.02fF
C50005 OR2X1_LOC_632/Y OR2X1_LOC_735/B 0.23fF
C50006 OR2X1_LOC_3/Y OR2X1_LOC_751/a_8_216# 0.01fF
C50007 VDD AND2X1_LOC_204/a_8_24# -0.00fF
C50008 OR2X1_LOC_190/A AND2X1_LOC_36/Y 0.15fF
C50009 OR2X1_LOC_95/Y AND2X1_LOC_260/a_8_24# 0.14fF
C50010 AND2X1_LOC_571/Y AND2X1_LOC_563/Y 0.01fF
C50011 OR2X1_LOC_812/B OR2X1_LOC_561/B 0.18fF
C50012 AND2X1_LOC_44/Y AND2X1_LOC_248/a_8_24# 0.01fF
C50013 OR2X1_LOC_65/B OR2X1_LOC_88/Y 0.03fF
C50014 OR2X1_LOC_805/A OR2X1_LOC_228/Y 0.07fF
C50015 OR2X1_LOC_39/A OR2X1_LOC_153/a_36_216# 0.00fF
C50016 OR2X1_LOC_256/Y OR2X1_LOC_13/B 0.04fF
C50017 OR2X1_LOC_516/a_36_216# AND2X1_LOC_469/B 0.00fF
C50018 OR2X1_LOC_786/Y AND2X1_LOC_51/Y 3.01fF
C50019 AND2X1_LOC_798/a_36_24# AND2X1_LOC_436/Y 0.01fF
C50020 OR2X1_LOC_449/B OR2X1_LOC_854/A 0.03fF
C50021 AND2X1_LOC_287/B AND2X1_LOC_243/Y 0.00fF
C50022 OR2X1_LOC_134/Y AND2X1_LOC_768/a_8_24# 0.01fF
C50023 OR2X1_LOC_316/a_8_216# OR2X1_LOC_59/Y 0.08fF
C50024 OR2X1_LOC_62/A OR2X1_LOC_62/a_8_216# 0.05fF
C50025 AND2X1_LOC_43/B AND2X1_LOC_419/a_36_24# 0.01fF
C50026 AND2X1_LOC_50/Y AND2X1_LOC_36/Y 0.03fF
C50027 OR2X1_LOC_12/Y AND2X1_LOC_605/a_8_24# 0.01fF
C50028 OR2X1_LOC_322/Y OR2X1_LOC_323/a_8_216# 0.04fF
C50029 AND2X1_LOC_707/Y OR2X1_LOC_681/a_8_216# 0.04fF
C50030 VDD OR2X1_LOC_392/B 2.02fF
C50031 AND2X1_LOC_785/Y AND2X1_LOC_778/Y 0.41fF
C50032 AND2X1_LOC_70/Y OR2X1_LOC_390/a_8_216# 0.00fF
C50033 AND2X1_LOC_633/Y OR2X1_LOC_47/Y 0.18fF
C50034 OR2X1_LOC_604/A AND2X1_LOC_244/A 0.05fF
C50035 OR2X1_LOC_673/A INPUT_1 0.03fF
C50036 OR2X1_LOC_631/A OR2X1_LOC_161/B 0.02fF
C50037 OR2X1_LOC_754/A OR2X1_LOC_753/Y 0.27fF
C50038 AND2X1_LOC_70/Y OR2X1_LOC_855/A 0.01fF
C50039 AND2X1_LOC_48/A OR2X1_LOC_207/a_36_216# 0.02fF
C50040 AND2X1_LOC_831/Y AND2X1_LOC_649/Y 0.91fF
C50041 AND2X1_LOC_34/a_8_24# OR2X1_LOC_68/B 0.01fF
C50042 OR2X1_LOC_485/A AND2X1_LOC_570/a_8_24# 0.04fF
C50043 OR2X1_LOC_282/a_8_216# AND2X1_LOC_562/Y 0.48fF
C50044 OR2X1_LOC_604/A OR2X1_LOC_16/A 0.18fF
C50045 OR2X1_LOC_47/Y D_INPUT_0 2.28fF
C50046 AND2X1_LOC_56/B OR2X1_LOC_728/A 0.05fF
C50047 OR2X1_LOC_158/A AND2X1_LOC_476/Y 2.20fF
C50048 OR2X1_LOC_669/A OR2X1_LOC_437/A 0.11fF
C50049 OR2X1_LOC_139/A AND2X1_LOC_92/Y 0.07fF
C50050 OR2X1_LOC_329/B AND2X1_LOC_241/a_36_24# 0.01fF
C50051 OR2X1_LOC_121/B OR2X1_LOC_318/B 0.04fF
C50052 OR2X1_LOC_246/A OR2X1_LOC_86/A 0.03fF
C50053 OR2X1_LOC_630/B OR2X1_LOC_563/A 0.03fF
C50054 OR2X1_LOC_475/Y AND2X1_LOC_31/Y 0.02fF
C50055 OR2X1_LOC_797/a_8_216# OR2X1_LOC_160/Y 0.01fF
C50056 AND2X1_LOC_64/Y OR2X1_LOC_840/A 0.29fF
C50057 INPUT_1 AND2X1_LOC_462/B 0.09fF
C50058 AND2X1_LOC_47/Y AND2X1_LOC_8/a_8_24# 0.09fF
C50059 AND2X1_LOC_81/B OR2X1_LOC_771/B 0.05fF
C50060 VDD OR2X1_LOC_113/B 0.15fF
C50061 VDD AND2X1_LOC_714/B 0.35fF
C50062 AND2X1_LOC_212/A AND2X1_LOC_568/B 0.02fF
C50063 OR2X1_LOC_329/B AND2X1_LOC_802/Y 0.03fF
C50064 OR2X1_LOC_56/A AND2X1_LOC_795/a_36_24# 0.01fF
C50065 OR2X1_LOC_632/Y OR2X1_LOC_161/B 0.02fF
C50066 AND2X1_LOC_515/a_8_24# AND2X1_LOC_469/B 0.01fF
C50067 D_INPUT_0 OR2X1_LOC_351/a_8_216# 0.04fF
C50068 AND2X1_LOC_47/Y OR2X1_LOC_545/a_8_216# 0.01fF
C50069 OR2X1_LOC_604/A OR2X1_LOC_108/Y 0.10fF
C50070 OR2X1_LOC_532/B OR2X1_LOC_76/a_8_216# 0.03fF
C50071 OR2X1_LOC_479/Y OR2X1_LOC_303/B 0.10fF
C50072 AND2X1_LOC_232/a_8_24# OR2X1_LOC_549/A 0.01fF
C50073 OR2X1_LOC_87/A AND2X1_LOC_238/a_8_24# 0.03fF
C50074 AND2X1_LOC_367/A OR2X1_LOC_522/Y 0.05fF
C50075 OR2X1_LOC_715/B OR2X1_LOC_648/A 0.10fF
C50076 AND2X1_LOC_566/B AND2X1_LOC_514/a_8_24# 0.01fF
C50077 AND2X1_LOC_543/a_8_24# OR2X1_LOC_323/Y 0.23fF
C50078 VDD OR2X1_LOC_450/A 0.21fF
C50079 OR2X1_LOC_786/A OR2X1_LOC_78/A 0.01fF
C50080 OR2X1_LOC_165/a_8_216# AND2X1_LOC_787/A 0.01fF
C50081 OR2X1_LOC_696/A OR2X1_LOC_6/A 0.17fF
C50082 AND2X1_LOC_806/a_8_24# OR2X1_LOC_56/A 0.01fF
C50083 OR2X1_LOC_95/Y OR2X1_LOC_749/a_8_216# 0.01fF
C50084 INPUT_0 AND2X1_LOC_200/a_8_24# 0.01fF
C50085 OR2X1_LOC_158/A AND2X1_LOC_198/a_8_24# 0.04fF
C50086 OR2X1_LOC_110/a_8_216# OR2X1_LOC_36/Y 0.01fF
C50087 AND2X1_LOC_850/a_8_24# AND2X1_LOC_244/A 0.01fF
C50088 AND2X1_LOC_91/B OR2X1_LOC_241/a_8_216# 0.33fF
C50089 OR2X1_LOC_160/B INPUT_0 0.07fF
C50090 OR2X1_LOC_529/Y OR2X1_LOC_183/Y 0.06fF
C50091 OR2X1_LOC_117/a_36_216# AND2X1_LOC_99/A 0.01fF
C50092 AND2X1_LOC_191/B AND2X1_LOC_658/A 0.01fF
C50093 AND2X1_LOC_658/A AND2X1_LOC_469/B 0.03fF
C50094 OR2X1_LOC_151/A OR2X1_LOC_502/A 0.57fF
C50095 AND2X1_LOC_362/B OR2X1_LOC_103/Y 0.01fF
C50096 OR2X1_LOC_135/a_36_216# OR2X1_LOC_48/B 0.00fF
C50097 AND2X1_LOC_214/A VDD 0.19fF
C50098 OR2X1_LOC_335/a_36_216# OR2X1_LOC_87/A 0.02fF
C50099 OR2X1_LOC_551/B OR2X1_LOC_364/a_36_216# 0.00fF
C50100 OR2X1_LOC_113/a_8_216# OR2X1_LOC_154/A 0.04fF
C50101 OR2X1_LOC_448/Y AND2X1_LOC_44/Y 0.00fF
C50102 OR2X1_LOC_336/a_36_216# OR2X1_LOC_212/A 0.00fF
C50103 OR2X1_LOC_506/A AND2X1_LOC_433/a_8_24# 0.18fF
C50104 VDD AND2X1_LOC_861/B 0.01fF
C50105 OR2X1_LOC_154/A OR2X1_LOC_474/B 0.01fF
C50106 AND2X1_LOC_456/B OR2X1_LOC_666/a_36_216# 0.00fF
C50107 OR2X1_LOC_306/a_8_216# OR2X1_LOC_12/Y 0.15fF
C50108 AND2X1_LOC_322/a_8_24# OR2X1_LOC_502/A 0.04fF
C50109 OR2X1_LOC_45/B AND2X1_LOC_303/A 0.01fF
C50110 AND2X1_LOC_802/B OR2X1_LOC_44/Y 0.03fF
C50111 AND2X1_LOC_675/Y AND2X1_LOC_663/A 0.19fF
C50112 AND2X1_LOC_571/A AND2X1_LOC_489/Y 0.03fF
C50113 OR2X1_LOC_709/A OR2X1_LOC_377/A 0.25fF
C50114 AND2X1_LOC_706/Y AND2X1_LOC_435/a_8_24# 0.03fF
C50115 OR2X1_LOC_535/A OR2X1_LOC_161/A 0.01fF
C50116 OR2X1_LOC_756/B OR2X1_LOC_35/Y 0.02fF
C50117 OR2X1_LOC_696/A AND2X1_LOC_557/a_8_24# 0.03fF
C50118 OR2X1_LOC_235/B OR2X1_LOC_78/B 0.07fF
C50119 AND2X1_LOC_723/a_8_24# OR2X1_LOC_40/Y 0.02fF
C50120 OR2X1_LOC_100/Y VDD 0.20fF
C50121 OR2X1_LOC_359/A OR2X1_LOC_756/B 0.04fF
C50122 OR2X1_LOC_200/a_36_216# AND2X1_LOC_7/B 0.02fF
C50123 OR2X1_LOC_220/B OR2X1_LOC_565/A 0.01fF
C50124 OR2X1_LOC_8/Y OR2X1_LOC_92/Y 0.02fF
C50125 AND2X1_LOC_729/Y AND2X1_LOC_729/a_8_24# 0.02fF
C50126 OR2X1_LOC_275/Y AND2X1_LOC_218/Y 0.02fF
C50127 OR2X1_LOC_158/A OR2X1_LOC_595/a_8_216# 0.01fF
C50128 OR2X1_LOC_40/Y OR2X1_LOC_278/Y 0.03fF
C50129 OR2X1_LOC_80/Y OR2X1_LOC_16/A 0.02fF
C50130 OR2X1_LOC_653/Y AND2X1_LOC_18/Y 0.09fF
C50131 OR2X1_LOC_115/a_8_216# OR2X1_LOC_6/B 0.07fF
C50132 AND2X1_LOC_56/B OR2X1_LOC_138/A 0.04fF
C50133 D_INPUT_3 OR2X1_LOC_384/Y 0.46fF
C50134 OR2X1_LOC_40/Y AND2X1_LOC_662/B 0.11fF
C50135 AND2X1_LOC_191/Y AND2X1_LOC_192/a_8_24# 0.01fF
C50136 OR2X1_LOC_43/A AND2X1_LOC_786/Y 0.07fF
C50137 OR2X1_LOC_483/a_8_216# OR2X1_LOC_736/Y 0.05fF
C50138 OR2X1_LOC_833/B AND2X1_LOC_18/Y 0.01fF
C50139 VDD AND2X1_LOC_820/a_8_24# -0.00fF
C50140 OR2X1_LOC_280/Y AND2X1_LOC_284/a_8_24# 0.11fF
C50141 OR2X1_LOC_45/B AND2X1_LOC_474/Y 0.03fF
C50142 OR2X1_LOC_679/A OR2X1_LOC_142/Y 0.15fF
C50143 OR2X1_LOC_175/Y OR2X1_LOC_702/A 0.10fF
C50144 OR2X1_LOC_114/B OR2X1_LOC_128/A 0.03fF
C50145 OR2X1_LOC_528/Y AND2X1_LOC_186/a_8_24# 0.16fF
C50146 OR2X1_LOC_235/B OR2X1_LOC_721/Y 0.05fF
C50147 OR2X1_LOC_735/a_8_216# OR2X1_LOC_736/A -0.00fF
C50148 OR2X1_LOC_2/Y OR2X1_LOC_25/Y 0.38fF
C50149 OR2X1_LOC_45/B OR2X1_LOC_485/A 0.10fF
C50150 AND2X1_LOC_22/Y AND2X1_LOC_386/a_36_24# 0.00fF
C50151 OR2X1_LOC_479/Y OR2X1_LOC_478/Y 0.13fF
C50152 AND2X1_LOC_723/Y AND2X1_LOC_722/A 0.01fF
C50153 OR2X1_LOC_160/B OR2X1_LOC_489/B -0.01fF
C50154 AND2X1_LOC_729/Y OR2X1_LOC_600/A 0.09fF
C50155 OR2X1_LOC_128/B OR2X1_LOC_66/A 0.01fF
C50156 VDD AND2X1_LOC_653/B 0.22fF
C50157 OR2X1_LOC_254/B AND2X1_LOC_18/Y 0.01fF
C50158 OR2X1_LOC_702/A OR2X1_LOC_691/Y 0.02fF
C50159 AND2X1_LOC_70/Y OR2X1_LOC_377/A 0.23fF
C50160 OR2X1_LOC_6/B OR2X1_LOC_673/Y 0.02fF
C50161 AND2X1_LOC_61/Y OR2X1_LOC_39/A 0.46fF
C50162 OR2X1_LOC_223/A OR2X1_LOC_716/a_8_216# 0.01fF
C50163 OR2X1_LOC_821/a_8_216# OR2X1_LOC_74/A 0.00fF
C50164 OR2X1_LOC_624/A OR2X1_LOC_78/A 0.05fF
C50165 OR2X1_LOC_426/B AND2X1_LOC_655/A 0.10fF
C50166 OR2X1_LOC_744/A OR2X1_LOC_432/Y 0.01fF
C50167 VDD OR2X1_LOC_685/A 0.21fF
C50168 AND2X1_LOC_110/Y AND2X1_LOC_298/a_8_24# 0.01fF
C50169 INPUT_3 INPUT_0 0.33fF
C50170 OR2X1_LOC_502/A OR2X1_LOC_651/B 0.10fF
C50171 OR2X1_LOC_7/A OR2X1_LOC_421/Y 0.26fF
C50172 OR2X1_LOC_17/Y OR2X1_LOC_12/Y 0.01fF
C50173 OR2X1_LOC_641/Y OR2X1_LOC_462/B 0.01fF
C50174 OR2X1_LOC_102/a_8_216# OR2X1_LOC_485/A 0.01fF
C50175 AND2X1_LOC_164/a_36_24# OR2X1_LOC_506/A 0.00fF
C50176 AND2X1_LOC_110/Y OR2X1_LOC_269/B 0.03fF
C50177 OR2X1_LOC_656/B AND2X1_LOC_41/A 0.02fF
C50178 OR2X1_LOC_329/Y OR2X1_LOC_585/A 0.01fF
C50179 OR2X1_LOC_638/B OR2X1_LOC_375/A 0.02fF
C50180 OR2X1_LOC_51/Y AND2X1_LOC_319/A 0.44fF
C50181 AND2X1_LOC_784/A OR2X1_LOC_600/A 0.07fF
C50182 OR2X1_LOC_317/a_8_216# OR2X1_LOC_317/A 0.47fF
C50183 AND2X1_LOC_33/a_8_24# OR2X1_LOC_6/A 0.17fF
C50184 AND2X1_LOC_784/A AND2X1_LOC_335/Y 0.02fF
C50185 OR2X1_LOC_372/a_36_216# AND2X1_LOC_786/Y 0.01fF
C50186 OR2X1_LOC_574/A OR2X1_LOC_362/A 0.08fF
C50187 AND2X1_LOC_605/Y AND2X1_LOC_593/Y 0.01fF
C50188 AND2X1_LOC_70/Y OR2X1_LOC_203/Y 0.08fF
C50189 VDD OR2X1_LOC_610/Y 0.12fF
C50190 OR2X1_LOC_235/B OR2X1_LOC_375/A 0.14fF
C50191 AND2X1_LOC_76/Y OR2X1_LOC_92/Y 0.05fF
C50192 OR2X1_LOC_91/Y OR2X1_LOC_91/A 0.01fF
C50193 AND2X1_LOC_580/A AND2X1_LOC_548/Y 0.16fF
C50194 OR2X1_LOC_592/a_8_216# OR2X1_LOC_66/A 0.01fF
C50195 AND2X1_LOC_658/A AND2X1_LOC_862/a_8_24# 0.01fF
C50196 OR2X1_LOC_143/a_36_216# D_INPUT_3 0.00fF
C50197 OR2X1_LOC_64/Y AND2X1_LOC_828/a_8_24# 0.01fF
C50198 AND2X1_LOC_333/a_8_24# AND2X1_LOC_338/A 0.01fF
C50199 OR2X1_LOC_134/a_8_216# AND2X1_LOC_227/Y 0.01fF
C50200 VDD AND2X1_LOC_645/A 0.24fF
C50201 OR2X1_LOC_243/A AND2X1_LOC_126/a_8_24# 0.08fF
C50202 AND2X1_LOC_810/A AND2X1_LOC_308/a_8_24# 0.01fF
C50203 AND2X1_LOC_158/a_8_24# OR2X1_LOC_803/A 0.01fF
C50204 OR2X1_LOC_154/A OR2X1_LOC_658/a_8_216# 0.04fF
C50205 OR2X1_LOC_744/A AND2X1_LOC_653/a_8_24# 0.01fF
C50206 AND2X1_LOC_777/a_36_24# OR2X1_LOC_56/A 0.00fF
C50207 OR2X1_LOC_154/A OR2X1_LOC_78/Y 0.02fF
C50208 AND2X1_LOC_31/a_36_24# AND2X1_LOC_44/Y 0.00fF
C50209 OR2X1_LOC_467/A OR2X1_LOC_449/a_8_216# 0.01fF
C50210 OR2X1_LOC_214/B AND2X1_LOC_36/Y 0.03fF
C50211 OR2X1_LOC_323/A AND2X1_LOC_866/A 0.03fF
C50212 OR2X1_LOC_154/A OR2X1_LOC_274/a_8_216# 0.00fF
C50213 AND2X1_LOC_12/Y OR2X1_LOC_489/a_8_216# 0.01fF
C50214 OR2X1_LOC_551/B OR2X1_LOC_181/Y 0.02fF
C50215 AND2X1_LOC_64/Y OR2X1_LOC_241/Y 0.10fF
C50216 OR2X1_LOC_528/Y OR2X1_LOC_617/Y 0.42fF
C50217 AND2X1_LOC_572/A OR2X1_LOC_517/A 0.05fF
C50218 OR2X1_LOC_469/Y OR2X1_LOC_738/A 0.01fF
C50219 AND2X1_LOC_705/a_8_24# OR2X1_LOC_485/A 0.09fF
C50220 OR2X1_LOC_691/Y OR2X1_LOC_644/a_8_216# 0.01fF
C50221 OR2X1_LOC_111/a_8_216# AND2X1_LOC_318/Y 0.14fF
C50222 AND2X1_LOC_41/A OR2X1_LOC_793/A 0.01fF
C50223 AND2X1_LOC_798/a_8_24# AND2X1_LOC_798/A 0.18fF
C50224 OR2X1_LOC_185/A AND2X1_LOC_74/a_8_24# 0.14fF
C50225 AND2X1_LOC_576/Y AND2X1_LOC_506/a_8_24# 0.03fF
C50226 OR2X1_LOC_92/Y OR2X1_LOC_67/A 0.12fF
C50227 OR2X1_LOC_161/A OR2X1_LOC_725/B 0.03fF
C50228 OR2X1_LOC_334/B OR2X1_LOC_87/B 0.00fF
C50229 OR2X1_LOC_538/A OR2X1_LOC_449/B 0.03fF
C50230 OR2X1_LOC_507/a_36_216# AND2X1_LOC_81/B 0.00fF
C50231 OR2X1_LOC_405/A OR2X1_LOC_506/A 0.03fF
C50232 AND2X1_LOC_47/a_8_24# AND2X1_LOC_11/Y 0.11fF
C50233 OR2X1_LOC_56/A OR2X1_LOC_371/Y 0.07fF
C50234 AND2X1_LOC_360/a_8_24# OR2X1_LOC_44/Y 0.03fF
C50235 OR2X1_LOC_809/B AND2X1_LOC_111/a_8_24# 0.04fF
C50236 AND2X1_LOC_597/a_8_24# AND2X1_LOC_40/Y 0.18fF
C50237 OR2X1_LOC_710/B OR2X1_LOC_705/Y 0.39fF
C50238 OR2X1_LOC_51/Y OR2X1_LOC_52/a_8_216# 0.17fF
C50239 AND2X1_LOC_566/B OR2X1_LOC_22/Y 0.02fF
C50240 AND2X1_LOC_794/B AND2X1_LOC_477/A 0.01fF
C50241 AND2X1_LOC_539/Y OR2X1_LOC_47/Y 0.03fF
C50242 OR2X1_LOC_40/Y OR2X1_LOC_19/B 0.07fF
C50243 AND2X1_LOC_552/a_8_24# OR2X1_LOC_47/Y 0.01fF
C50244 OR2X1_LOC_154/A OR2X1_LOC_724/a_8_216# 0.05fF
C50245 AND2X1_LOC_729/Y OR2X1_LOC_619/Y 0.07fF
C50246 OR2X1_LOC_864/A AND2X1_LOC_40/Y 0.03fF
C50247 D_INPUT_7 OR2X1_LOC_2/a_36_216# 0.00fF
C50248 AND2X1_LOC_660/Y OR2X1_LOC_59/Y 0.01fF
C50249 OR2X1_LOC_105/Y OR2X1_LOC_810/A 0.08fF
C50250 OR2X1_LOC_92/Y OR2X1_LOC_52/B 0.27fF
C50251 OR2X1_LOC_697/a_36_216# OR2X1_LOC_743/A 0.00fF
C50252 OR2X1_LOC_194/Y OR2X1_LOC_194/B 0.86fF
C50253 AND2X1_LOC_59/Y OR2X1_LOC_340/Y 0.00fF
C50254 AND2X1_LOC_711/Y OR2X1_LOC_755/a_36_216# 0.00fF
C50255 OR2X1_LOC_845/A AND2X1_LOC_263/a_8_24# 0.25fF
C50256 AND2X1_LOC_813/a_8_24# OR2X1_LOC_266/A 0.01fF
C50257 AND2X1_LOC_98/a_8_24# OR2X1_LOC_54/Y 0.03fF
C50258 AND2X1_LOC_568/B AND2X1_LOC_727/A 0.03fF
C50259 OR2X1_LOC_91/Y AND2X1_LOC_573/A 0.07fF
C50260 OR2X1_LOC_427/A OR2X1_LOC_418/Y 0.01fF
C50261 OR2X1_LOC_271/Y AND2X1_LOC_76/Y 0.02fF
C50262 AND2X1_LOC_59/Y OR2X1_LOC_130/A 0.09fF
C50263 AND2X1_LOC_40/Y OR2X1_LOC_633/B 0.05fF
C50264 OR2X1_LOC_663/A AND2X1_LOC_42/B 0.03fF
C50265 OR2X1_LOC_3/Y OR2X1_LOC_517/A 0.12fF
C50266 OR2X1_LOC_695/Y OR2X1_LOC_22/Y 0.09fF
C50267 OR2X1_LOC_45/B OR2X1_LOC_396/a_8_216# 0.00fF
C50268 OR2X1_LOC_770/A OR2X1_LOC_770/Y 0.01fF
C50269 AND2X1_LOC_553/A OR2X1_LOC_529/Y 0.01fF
C50270 OR2X1_LOC_274/a_8_216# OR2X1_LOC_778/A 0.14fF
C50271 AND2X1_LOC_99/A OR2X1_LOC_117/Y 0.66fF
C50272 AND2X1_LOC_489/Y OR2X1_LOC_92/Y 0.17fF
C50273 AND2X1_LOC_784/A OR2X1_LOC_619/Y 0.02fF
C50274 AND2X1_LOC_802/a_36_24# AND2X1_LOC_436/Y 0.00fF
C50275 VDD AND2X1_LOC_477/A 0.14fF
C50276 OR2X1_LOC_6/B OR2X1_LOC_4/a_8_216# 0.06fF
C50277 OR2X1_LOC_671/a_8_216# INPUT_1 0.01fF
C50278 OR2X1_LOC_417/Y OR2X1_LOC_91/A 0.00fF
C50279 OR2X1_LOC_532/B OR2X1_LOC_723/a_36_216# 0.00fF
C50280 AND2X1_LOC_338/a_8_24# OR2X1_LOC_46/A 0.09fF
C50281 OR2X1_LOC_655/a_36_216# AND2X1_LOC_8/Y 0.00fF
C50282 OR2X1_LOC_327/a_8_216# AND2X1_LOC_3/Y 0.01fF
C50283 OR2X1_LOC_496/Y AND2X1_LOC_621/Y 0.03fF
C50284 OR2X1_LOC_7/A OR2X1_LOC_278/Y 0.05fF
C50285 AND2X1_LOC_302/a_8_24# OR2X1_LOC_6/A 0.02fF
C50286 OR2X1_LOC_856/B AND2X1_LOC_387/B 0.01fF
C50287 OR2X1_LOC_311/Y OR2X1_LOC_91/A 0.03fF
C50288 AND2X1_LOC_12/Y OR2X1_LOC_449/B 0.03fF
C50289 VDD OR2X1_LOC_532/B 2.30fF
C50290 AND2X1_LOC_564/B OR2X1_LOC_406/A 0.01fF
C50291 OR2X1_LOC_95/Y AND2X1_LOC_243/Y 0.07fF
C50292 AND2X1_LOC_512/Y AND2X1_LOC_856/B 0.82fF
C50293 AND2X1_LOC_578/A OR2X1_LOC_495/Y 0.14fF
C50294 AND2X1_LOC_300/a_8_24# OR2X1_LOC_223/A 0.01fF
C50295 AND2X1_LOC_852/Y OR2X1_LOC_39/A 14.09fF
C50296 OR2X1_LOC_47/Y AND2X1_LOC_771/B 0.01fF
C50297 OR2X1_LOC_74/a_36_216# OR2X1_LOC_39/A 0.00fF
C50298 OR2X1_LOC_65/B OR2X1_LOC_52/B 0.95fF
C50299 AND2X1_LOC_385/a_36_24# OR2X1_LOC_537/A 0.00fF
C50300 OR2X1_LOC_271/B OR2X1_LOC_6/A 0.19fF
C50301 AND2X1_LOC_41/A AND2X1_LOC_45/a_8_24# 0.02fF
C50302 OR2X1_LOC_710/A AND2X1_LOC_31/Y 0.01fF
C50303 AND2X1_LOC_41/a_8_24# OR2X1_LOC_651/A -0.01fF
C50304 OR2X1_LOC_585/A OR2X1_LOC_69/A 0.04fF
C50305 OR2X1_LOC_703/B OR2X1_LOC_778/Y 0.22fF
C50306 AND2X1_LOC_561/B OR2X1_LOC_71/Y 0.01fF
C50307 OR2X1_LOC_835/A OR2X1_LOC_269/B 0.05fF
C50308 OR2X1_LOC_329/B INPUT_1 0.07fF
C50309 AND2X1_LOC_358/Y OR2X1_LOC_595/Y 0.00fF
C50310 OR2X1_LOC_85/A AND2X1_LOC_361/A 0.20fF
C50311 OR2X1_LOC_447/Y OR2X1_LOC_78/A 0.10fF
C50312 OR2X1_LOC_864/A OR2X1_LOC_848/A 0.01fF
C50313 OR2X1_LOC_287/B OR2X1_LOC_805/A 0.03fF
C50314 OR2X1_LOC_51/Y OR2X1_LOC_604/a_8_216# 0.01fF
C50315 OR2X1_LOC_318/a_8_216# OR2X1_LOC_804/A 0.40fF
C50316 OR2X1_LOC_116/a_8_216# OR2X1_LOC_203/Y 0.01fF
C50317 OR2X1_LOC_643/A OR2X1_LOC_87/A 0.07fF
C50318 OR2X1_LOC_419/Y OR2X1_LOC_373/Y 0.03fF
C50319 AND2X1_LOC_324/a_8_24# AND2X1_LOC_654/Y 0.02fF
C50320 AND2X1_LOC_228/Y AND2X1_LOC_654/a_36_24# 0.00fF
C50321 OR2X1_LOC_851/A AND2X1_LOC_51/Y 0.07fF
C50322 OR2X1_LOC_600/A OR2X1_LOC_62/A 0.07fF
C50323 OR2X1_LOC_87/A OR2X1_LOC_778/Y 0.10fF
C50324 OR2X1_LOC_774/Y OR2X1_LOC_848/A 0.18fF
C50325 INPUT_0 OR2X1_LOC_244/A 0.13fF
C50326 OR2X1_LOC_3/Y AND2X1_LOC_624/A 0.00fF
C50327 OR2X1_LOC_743/A AND2X1_LOC_655/A 0.17fF
C50328 OR2X1_LOC_76/Y OR2X1_LOC_455/a_8_216# 0.08fF
C50329 VDD OR2X1_LOC_343/B -0.00fF
C50330 OR2X1_LOC_271/Y OR2X1_LOC_52/B 0.08fF
C50331 OR2X1_LOC_774/Y OR2X1_LOC_859/B 0.04fF
C50332 OR2X1_LOC_70/Y OR2X1_LOC_298/Y 0.01fF
C50333 D_GATE_579 OR2X1_LOC_580/B 0.02fF
C50334 OR2X1_LOC_232/a_8_216# OR2X1_LOC_753/A 0.03fF
C50335 OR2X1_LOC_119/a_36_216# OR2X1_LOC_619/Y 0.01fF
C50336 AND2X1_LOC_658/A OR2X1_LOC_146/Y 0.03fF
C50337 OR2X1_LOC_377/A OR2X1_LOC_404/Y 0.03fF
C50338 AND2X1_LOC_211/B AND2X1_LOC_852/Y 0.02fF
C50339 OR2X1_LOC_485/A OR2X1_LOC_235/a_36_216# 0.01fF
C50340 OR2X1_LOC_502/A INPUT_1 0.06fF
C50341 OR2X1_LOC_62/B AND2X1_LOC_852/B 0.03fF
C50342 AND2X1_LOC_391/Y D_INPUT_3 0.01fF
C50343 OR2X1_LOC_64/Y AND2X1_LOC_452/Y 0.00fF
C50344 OR2X1_LOC_185/Y AND2X1_LOC_42/B 0.07fF
C50345 OR2X1_LOC_91/A D_INPUT_3 0.13fF
C50346 OR2X1_LOC_118/a_36_216# OR2X1_LOC_88/Y 0.00fF
C50347 OR2X1_LOC_479/Y AND2X1_LOC_56/B 0.07fF
C50348 OR2X1_LOC_291/Y AND2X1_LOC_573/A 0.07fF
C50349 OR2X1_LOC_828/B AND2X1_LOC_51/Y 0.04fF
C50350 AND2X1_LOC_12/Y OR2X1_LOC_121/B 8.95fF
C50351 AND2X1_LOC_643/a_36_24# OR2X1_LOC_46/A 0.00fF
C50352 AND2X1_LOC_116/a_8_24# OR2X1_LOC_56/A 0.00fF
C50353 OR2X1_LOC_182/B OR2X1_LOC_365/B 0.25fF
C50354 AND2X1_LOC_82/a_8_24# AND2X1_LOC_77/a_8_24# 0.23fF
C50355 AND2X1_LOC_42/B AND2X1_LOC_412/a_8_24# 0.10fF
C50356 AND2X1_LOC_177/a_8_24# OR2X1_LOC_440/A 0.01fF
C50357 OR2X1_LOC_51/Y AND2X1_LOC_721/A 0.08fF
C50358 OR2X1_LOC_686/B OR2X1_LOC_451/B 0.12fF
C50359 AND2X1_LOC_8/Y AND2X1_LOC_4/a_8_24# 0.01fF
C50360 OR2X1_LOC_118/Y OR2X1_LOC_46/A 0.07fF
C50361 D_INPUT_4 AND2X1_LOC_47/Y 0.44fF
C50362 OR2X1_LOC_835/B AND2X1_LOC_51/Y 0.22fF
C50363 OR2X1_LOC_401/Y AND2X1_LOC_490/a_8_24# 0.01fF
C50364 OR2X1_LOC_47/Y AND2X1_LOC_471/Y 0.03fF
C50365 AND2X1_LOC_573/A AND2X1_LOC_574/A 0.01fF
C50366 AND2X1_LOC_736/Y OR2X1_LOC_95/Y 1.23fF
C50367 AND2X1_LOC_663/B OR2X1_LOC_6/A 0.03fF
C50368 OR2X1_LOC_740/B OR2X1_LOC_739/a_36_216# 0.02fF
C50369 AND2X1_LOC_59/Y OR2X1_LOC_62/B 0.02fF
C50370 OR2X1_LOC_84/Y OR2X1_LOC_78/A 0.00fF
C50371 OR2X1_LOC_79/A OR2X1_LOC_89/A 0.01fF
C50372 OR2X1_LOC_318/Y OR2X1_LOC_436/Y 0.03fF
C50373 OR2X1_LOC_857/a_36_216# AND2X1_LOC_56/B 0.02fF
C50374 OR2X1_LOC_841/B OR2X1_LOC_121/B 0.01fF
C50375 AND2X1_LOC_755/a_8_24# OR2X1_LOC_532/B 0.23fF
C50376 OR2X1_LOC_233/a_8_216# OR2X1_LOC_291/A -0.00fF
C50377 OR2X1_LOC_36/Y OR2X1_LOC_268/a_8_216# 0.01fF
C50378 OR2X1_LOC_31/Y OR2X1_LOC_432/Y 0.26fF
C50379 AND2X1_LOC_811/Y AND2X1_LOC_808/a_8_24# 0.25fF
C50380 OR2X1_LOC_709/A OR2X1_LOC_732/A 0.14fF
C50381 AND2X1_LOC_227/Y OR2X1_LOC_118/Y 0.00fF
C50382 OR2X1_LOC_51/Y OR2X1_LOC_331/Y 0.13fF
C50383 OR2X1_LOC_70/A AND2X1_LOC_637/a_8_24# 0.09fF
C50384 OR2X1_LOC_836/A OR2X1_LOC_835/Y 0.01fF
C50385 OR2X1_LOC_823/a_8_216# D_INPUT_3 0.01fF
C50386 OR2X1_LOC_600/A OR2X1_LOC_172/Y 0.07fF
C50387 OR2X1_LOC_56/A AND2X1_LOC_222/Y 0.06fF
C50388 OR2X1_LOC_188/Y AND2X1_LOC_36/Y 1.20fF
C50389 OR2X1_LOC_71/Y AND2X1_LOC_266/Y 0.01fF
C50390 OR2X1_LOC_62/A OR2X1_LOC_619/Y -0.01fF
C50391 OR2X1_LOC_54/a_8_216# OR2X1_LOC_6/A 0.01fF
C50392 OR2X1_LOC_19/B OR2X1_LOC_7/A 0.03fF
C50393 D_INPUT_3 AND2X1_LOC_573/A 0.12fF
C50394 OR2X1_LOC_829/A OR2X1_LOC_13/B 0.10fF
C50395 AND2X1_LOC_494/a_36_24# OR2X1_LOC_269/B 0.00fF
C50396 OR2X1_LOC_412/a_8_216# OR2X1_LOC_690/A 0.02fF
C50397 OR2X1_LOC_405/A AND2X1_LOC_420/a_8_24# 0.00fF
C50398 AND2X1_LOC_67/Y OR2X1_LOC_202/a_8_216# 0.02fF
C50399 OR2X1_LOC_696/A OR2X1_LOC_184/a_8_216# 0.01fF
C50400 OR2X1_LOC_321/Y OR2X1_LOC_64/Y 0.01fF
C50401 AND2X1_LOC_139/B AND2X1_LOC_649/Y 0.26fF
C50402 OR2X1_LOC_673/Y AND2X1_LOC_47/Y 0.20fF
C50403 OR2X1_LOC_121/B OR2X1_LOC_804/B 0.13fF
C50404 OR2X1_LOC_70/Y OR2X1_LOC_683/Y 0.01fF
C50405 OR2X1_LOC_405/A D_INPUT_1 0.01fF
C50406 AND2X1_LOC_648/B AND2X1_LOC_436/B 0.00fF
C50407 OR2X1_LOC_841/a_8_216# OR2X1_LOC_318/B 0.00fF
C50408 OR2X1_LOC_447/Y OR2X1_LOC_155/A 0.03fF
C50409 OR2X1_LOC_92/Y AND2X1_LOC_216/A 0.06fF
C50410 OR2X1_LOC_769/A AND2X1_LOC_409/a_8_24# 0.20fF
C50411 OR2X1_LOC_40/Y AND2X1_LOC_608/a_8_24# 0.01fF
C50412 OR2X1_LOC_234/a_36_216# OR2X1_LOC_619/Y 0.01fF
C50413 AND2X1_LOC_40/Y OR2X1_LOC_608/Y 0.37fF
C50414 OR2X1_LOC_262/Y AND2X1_LOC_227/Y 1.73fF
C50415 OR2X1_LOC_71/a_36_216# OR2X1_LOC_67/Y 0.01fF
C50416 OR2X1_LOC_333/B AND2X1_LOC_431/a_8_24# 0.01fF
C50417 OR2X1_LOC_61/Y OR2X1_LOC_358/A 0.00fF
C50418 AND2X1_LOC_70/Y OR2X1_LOC_732/A 0.14fF
C50419 OR2X1_LOC_168/Y OR2X1_LOC_161/B 0.03fF
C50420 OR2X1_LOC_39/Y OR2X1_LOC_39/a_8_216# 0.01fF
C50421 OR2X1_LOC_115/a_8_216# OR2X1_LOC_598/A 0.02fF
C50422 OR2X1_LOC_195/A AND2X1_LOC_47/Y 0.01fF
C50423 OR2X1_LOC_448/a_8_216# OR2X1_LOC_779/B 0.00fF
C50424 OR2X1_LOC_185/A OR2X1_LOC_590/a_8_216# 0.01fF
C50425 AND2X1_LOC_848/A AND2X1_LOC_847/Y 0.23fF
C50426 D_INPUT_0 OR2X1_LOC_8/a_8_216# 0.06fF
C50427 OR2X1_LOC_65/B AND2X1_LOC_216/A 0.02fF
C50428 OR2X1_LOC_63/a_36_216# AND2X1_LOC_647/Y 0.00fF
C50429 AND2X1_LOC_199/a_8_24# AND2X1_LOC_729/B 0.00fF
C50430 AND2X1_LOC_59/Y OR2X1_LOC_365/B 0.01fF
C50431 OR2X1_LOC_186/Y OR2X1_LOC_303/a_8_216# 0.06fF
C50432 OR2X1_LOC_562/A OR2X1_LOC_580/B 0.03fF
C50433 AND2X1_LOC_573/A AND2X1_LOC_656/a_8_24# 0.01fF
C50434 OR2X1_LOC_161/a_8_216# OR2X1_LOC_162/A -0.00fF
C50435 OR2X1_LOC_427/A AND2X1_LOC_796/A 0.01fF
C50436 AND2X1_LOC_70/Y OR2X1_LOC_539/B 0.02fF
C50437 OR2X1_LOC_86/Y OR2X1_LOC_86/A 0.01fF
C50438 OR2X1_LOC_619/Y OR2X1_LOC_172/Y 0.05fF
C50439 AND2X1_LOC_31/Y AND2X1_LOC_43/B 0.38fF
C50440 OR2X1_LOC_99/A OR2X1_LOC_99/a_36_216# 0.00fF
C50441 OR2X1_LOC_375/A AND2X1_LOC_430/B 0.00fF
C50442 OR2X1_LOC_476/Y OR2X1_LOC_223/A 0.01fF
C50443 OR2X1_LOC_680/A OR2X1_LOC_331/Y 0.13fF
C50444 AND2X1_LOC_43/B OR2X1_LOC_715/a_8_216# 0.01fF
C50445 OR2X1_LOC_375/A OR2X1_LOC_779/B 0.84fF
C50446 OR2X1_LOC_134/Y AND2X1_LOC_541/Y 1.17fF
C50447 OR2X1_LOC_589/A AND2X1_LOC_202/Y 0.01fF
C50448 AND2X1_LOC_22/Y AND2X1_LOC_65/A 0.03fF
C50449 OR2X1_LOC_743/A OR2X1_LOC_599/Y 0.03fF
C50450 OR2X1_LOC_64/Y AND2X1_LOC_687/a_8_24# 0.01fF
C50451 AND2X1_LOC_56/B OR2X1_LOC_68/B 0.07fF
C50452 OR2X1_LOC_177/Y OR2X1_LOC_373/Y 0.17fF
C50453 AND2X1_LOC_209/a_36_24# AND2X1_LOC_220/B 0.01fF
C50454 OR2X1_LOC_486/Y OR2X1_LOC_344/A 0.03fF
C50455 OR2X1_LOC_160/B AND2X1_LOC_7/B 0.96fF
C50456 OR2X1_LOC_469/Y AND2X1_LOC_36/Y 0.00fF
C50457 AND2X1_LOC_8/Y OR2X1_LOC_68/B 0.12fF
C50458 AND2X1_LOC_423/a_8_24# AND2X1_LOC_36/Y 0.01fF
C50459 OR2X1_LOC_406/Y VDD -0.00fF
C50460 OR2X1_LOC_739/A OR2X1_LOC_550/B 0.03fF
C50461 OR2X1_LOC_865/A VDD 0.07fF
C50462 AND2X1_LOC_706/Y OR2X1_LOC_158/A 0.07fF
C50463 AND2X1_LOC_535/Y AND2X1_LOC_809/a_8_24# 0.01fF
C50464 OR2X1_LOC_604/A OR2X1_LOC_373/Y 0.03fF
C50465 AND2X1_LOC_703/Y VDD 0.21fF
C50466 OR2X1_LOC_487/Y AND2X1_LOC_563/Y 0.01fF
C50467 AND2X1_LOC_572/a_8_24# OR2X1_LOC_744/A 0.01fF
C50468 AND2X1_LOC_776/a_8_24# AND2X1_LOC_786/Y 0.02fF
C50469 OR2X1_LOC_696/A OR2X1_LOC_485/a_8_216# 0.02fF
C50470 OR2X1_LOC_188/Y AND2X1_LOC_368/a_8_24# 0.01fF
C50471 OR2X1_LOC_178/Y OR2X1_LOC_428/A 0.04fF
C50472 AND2X1_LOC_64/Y OR2X1_LOC_216/A 0.74fF
C50473 OR2X1_LOC_158/A OR2X1_LOC_58/Y 0.05fF
C50474 OR2X1_LOC_663/A AND2X1_LOC_224/a_8_24# 0.01fF
C50475 OR2X1_LOC_676/Y OR2X1_LOC_596/A 0.39fF
C50476 AND2X1_LOC_397/a_8_24# AND2X1_LOC_82/Y 0.09fF
C50477 VDD D_GATE_811 0.06fF
C50478 D_INPUT_0 OR2X1_LOC_512/a_36_216# 0.03fF
C50479 OR2X1_LOC_532/B OR2X1_LOC_737/a_36_216# 0.00fF
C50480 OR2X1_LOC_175/Y OR2X1_LOC_802/a_8_216# 0.07fF
C50481 OR2X1_LOC_6/B AND2X1_LOC_131/a_36_24# 0.01fF
C50482 OR2X1_LOC_417/A AND2X1_LOC_793/Y 0.03fF
C50483 OR2X1_LOC_709/A OR2X1_LOC_78/B 0.09fF
C50484 OR2X1_LOC_346/A OR2X1_LOC_78/A 0.07fF
C50485 OR2X1_LOC_49/A OR2X1_LOC_382/Y 0.01fF
C50486 OR2X1_LOC_151/A OR2X1_LOC_632/a_8_216# 0.02fF
C50487 OR2X1_LOC_643/A OR2X1_LOC_844/B 0.00fF
C50488 AND2X1_LOC_8/a_8_24# D_INPUT_1 0.01fF
C50489 OR2X1_LOC_8/Y OR2X1_LOC_600/A 0.21fF
C50490 AND2X1_LOC_64/Y OR2X1_LOC_499/a_8_216# 0.01fF
C50491 D_GATE_741 OR2X1_LOC_565/A 0.03fF
C50492 OR2X1_LOC_147/B OR2X1_LOC_578/a_8_216# 0.06fF
C50493 OR2X1_LOC_696/A OR2X1_LOC_44/Y 0.66fF
C50494 AND2X1_LOC_662/B AND2X1_LOC_476/a_8_24# 0.01fF
C50495 OR2X1_LOC_464/A OR2X1_LOC_741/a_8_216# 0.01fF
C50496 OR2X1_LOC_176/Y AND2X1_LOC_168/Y 0.09fF
C50497 OR2X1_LOC_302/a_8_216# OR2X1_LOC_302/A 0.01fF
C50498 OR2X1_LOC_506/a_8_216# AND2X1_LOC_81/B 0.01fF
C50499 OR2X1_LOC_151/A OR2X1_LOC_201/A 0.13fF
C50500 OR2X1_LOC_7/A OR2X1_LOC_504/a_8_216# 0.07fF
C50501 AND2X1_LOC_91/B OR2X1_LOC_703/B 0.06fF
C50502 OR2X1_LOC_122/Y AND2X1_LOC_243/Y 0.03fF
C50503 OR2X1_LOC_302/a_8_216# VDD 0.21fF
C50504 OR2X1_LOC_449/B OR2X1_LOC_356/B 0.07fF
C50505 AND2X1_LOC_64/Y OR2X1_LOC_468/Y 0.24fF
C50506 OR2X1_LOC_787/Y OR2X1_LOC_301/a_36_216# 0.01fF
C50507 VDD OR2X1_LOC_624/Y 0.14fF
C50508 AND2X1_LOC_765/a_8_24# OR2X1_LOC_402/Y 0.04fF
C50509 AND2X1_LOC_724/A OR2X1_LOC_48/B 0.07fF
C50510 AND2X1_LOC_723/Y OR2X1_LOC_40/Y 0.01fF
C50511 D_GATE_741 OR2X1_LOC_190/Y 0.09fF
C50512 AND2X1_LOC_91/B OR2X1_LOC_87/A 0.03fF
C50513 OR2X1_LOC_168/B OR2X1_LOC_468/A 0.00fF
C50514 AND2X1_LOC_787/A OR2X1_LOC_39/A 0.05fF
C50515 OR2X1_LOC_53/Y AND2X1_LOC_193/a_8_24# 0.18fF
C50516 AND2X1_LOC_70/Y OR2X1_LOC_78/B 5.18fF
C50517 AND2X1_LOC_540/a_36_24# OR2X1_LOC_158/A 0.00fF
C50518 AND2X1_LOC_95/Y AND2X1_LOC_603/a_8_24# 0.03fF
C50519 AND2X1_LOC_7/B OR2X1_LOC_553/A 0.11fF
C50520 OR2X1_LOC_700/a_8_216# OR2X1_LOC_59/Y 0.03fF
C50521 OR2X1_LOC_329/B AND2X1_LOC_352/B 0.03fF
C50522 AND2X1_LOC_168/Y AND2X1_LOC_212/Y 0.03fF
C50523 OR2X1_LOC_814/A OR2X1_LOC_366/Y 0.11fF
C50524 VDD OR2X1_LOC_391/A 0.21fF
C50525 OR2X1_LOC_154/A OR2X1_LOC_853/a_8_216# 0.01fF
C50526 OR2X1_LOC_59/Y AND2X1_LOC_434/Y 0.01fF
C50527 OR2X1_LOC_193/A AND2X1_LOC_36/Y 0.02fF
C50528 AND2X1_LOC_716/Y AND2X1_LOC_357/A 0.02fF
C50529 OR2X1_LOC_59/Y AND2X1_LOC_219/Y 0.09fF
C50530 AND2X1_LOC_715/Y OR2X1_LOC_44/Y 0.07fF
C50531 OR2X1_LOC_604/A OR2X1_LOC_426/A 0.03fF
C50532 AND2X1_LOC_605/Y OR2X1_LOC_51/Y 0.01fF
C50533 AND2X1_LOC_126/a_8_24# OR2X1_LOC_66/A -0.00fF
C50534 OR2X1_LOC_635/A OR2X1_LOC_686/B 0.26fF
C50535 AND2X1_LOC_531/a_8_24# VDD -0.00fF
C50536 OR2X1_LOC_323/A OR2X1_LOC_7/A 0.10fF
C50537 AND2X1_LOC_367/A OR2X1_LOC_56/A 0.16fF
C50538 OR2X1_LOC_778/B OR2X1_LOC_778/a_36_216# 0.01fF
C50539 OR2X1_LOC_325/a_8_216# OR2X1_LOC_325/B 0.47fF
C50540 AND2X1_LOC_799/a_36_24# AND2X1_LOC_661/A 0.00fF
C50541 OR2X1_LOC_49/A OR2X1_LOC_462/B 0.01fF
C50542 OR2X1_LOC_16/A OR2X1_LOC_265/Y 0.03fF
C50543 AND2X1_LOC_357/A AND2X1_LOC_654/Y 0.03fF
C50544 OR2X1_LOC_45/B OR2X1_LOC_495/a_8_216# 0.09fF
C50545 OR2X1_LOC_113/Y OR2X1_LOC_235/B 0.00fF
C50546 OR2X1_LOC_709/A OR2X1_LOC_375/A 0.00fF
C50547 OR2X1_LOC_712/a_8_216# OR2X1_LOC_66/A 0.02fF
C50548 AND2X1_LOC_339/B OR2X1_LOC_316/Y 0.00fF
C50549 OR2X1_LOC_318/a_8_216# OR2X1_LOC_130/A 0.05fF
C50550 AND2X1_LOC_70/Y OR2X1_LOC_721/Y 0.03fF
C50551 OR2X1_LOC_529/Y AND2X1_LOC_465/A 0.00fF
C50552 OR2X1_LOC_219/B AND2X1_LOC_7/B 0.03fF
C50553 AND2X1_LOC_566/B AND2X1_LOC_661/a_36_24# 0.00fF
C50554 AND2X1_LOC_567/a_8_24# AND2X1_LOC_841/B 0.02fF
C50555 VDD OR2X1_LOC_714/Y 0.00fF
C50556 AND2X1_LOC_624/A AND2X1_LOC_477/Y 0.07fF
C50557 OR2X1_LOC_158/A OR2X1_LOC_94/a_8_216# 0.02fF
C50558 OR2X1_LOC_744/A OR2X1_LOC_594/a_36_216# -0.00fF
C50559 OR2X1_LOC_769/A OR2X1_LOC_502/A 0.01fF
C50560 AND2X1_LOC_91/B AND2X1_LOC_815/a_8_24# 0.01fF
C50561 AND2X1_LOC_787/A AND2X1_LOC_211/B 0.03fF
C50562 OR2X1_LOC_84/B AND2X1_LOC_44/Y 0.07fF
C50563 OR2X1_LOC_7/A OR2X1_LOC_744/a_8_216# 0.04fF
C50564 OR2X1_LOC_113/A OR2X1_LOC_844/B 0.15fF
C50565 OR2X1_LOC_141/B AND2X1_LOC_44/Y 0.03fF
C50566 OR2X1_LOC_139/a_8_216# OR2X1_LOC_161/B 0.01fF
C50567 D_INPUT_0 AND2X1_LOC_36/Y 0.95fF
C50568 AND2X1_LOC_769/a_8_24# AND2X1_LOC_769/Y 0.00fF
C50569 OR2X1_LOC_529/Y OR2X1_LOC_530/a_36_216# 0.00fF
C50570 OR2X1_LOC_9/Y OR2X1_LOC_85/A 0.36fF
C50571 OR2X1_LOC_8/Y OR2X1_LOC_619/Y 0.16fF
C50572 OR2X1_LOC_756/B OR2X1_LOC_840/A 0.03fF
C50573 OR2X1_LOC_175/Y OR2X1_LOC_863/B 0.06fF
C50574 OR2X1_LOC_329/B AND2X1_LOC_833/a_8_24# 0.01fF
C50575 AND2X1_LOC_846/a_8_24# AND2X1_LOC_793/B 0.04fF
C50576 OR2X1_LOC_600/A OR2X1_LOC_67/A 0.03fF
C50577 OR2X1_LOC_632/a_36_216# OR2X1_LOC_575/A 0.01fF
C50578 OR2X1_LOC_160/B OR2X1_LOC_805/A 0.30fF
C50579 OR2X1_LOC_604/A INPUT_4 0.00fF
C50580 OR2X1_LOC_666/A OR2X1_LOC_18/Y 0.17fF
C50581 AND2X1_LOC_716/Y AND2X1_LOC_303/a_36_24# 0.01fF
C50582 OR2X1_LOC_856/B OR2X1_LOC_538/A 0.16fF
C50583 AND2X1_LOC_59/Y OR2X1_LOC_468/A 0.03fF
C50584 AND2X1_LOC_719/Y OR2X1_LOC_497/Y 0.10fF
C50585 OR2X1_LOC_258/Y OR2X1_LOC_428/A 0.02fF
C50586 AND2X1_LOC_571/A OR2X1_LOC_22/Y 0.01fF
C50587 OR2X1_LOC_3/Y AND2X1_LOC_774/A 0.01fF
C50588 OR2X1_LOC_857/B OR2X1_LOC_688/a_8_216# 0.01fF
C50589 OR2X1_LOC_655/a_36_216# AND2X1_LOC_92/Y 0.00fF
C50590 AND2X1_LOC_91/a_8_24# AND2X1_LOC_51/Y 0.06fF
C50591 AND2X1_LOC_201/a_8_24# AND2X1_LOC_206/a_8_24# 0.23fF
C50592 OR2X1_LOC_78/A OR2X1_LOC_161/A 2.17fF
C50593 AND2X1_LOC_392/A OR2X1_LOC_6/A 0.18fF
C50594 AND2X1_LOC_70/Y OR2X1_LOC_375/A 0.17fF
C50595 OR2X1_LOC_762/Y OR2X1_LOC_48/B 0.29fF
C50596 OR2X1_LOC_744/A AND2X1_LOC_652/a_8_24# 0.01fF
C50597 OR2X1_LOC_685/B OR2X1_LOC_687/A 0.12fF
C50598 AND2X1_LOC_566/B AND2X1_LOC_211/B 0.03fF
C50599 AND2X1_LOC_365/a_8_24# OR2X1_LOC_619/Y 0.05fF
C50600 AND2X1_LOC_61/Y OR2X1_LOC_85/A 0.04fF
C50601 OR2X1_LOC_151/A AND2X1_LOC_3/Y 0.07fF
C50602 INPUT_0 AND2X1_LOC_233/a_8_24# 0.01fF
C50603 OR2X1_LOC_756/B OR2X1_LOC_260/a_8_216# 0.02fF
C50604 AND2X1_LOC_19/Y AND2X1_LOC_129/a_8_24# 0.22fF
C50605 VDD OR2X1_LOC_99/a_8_216# 0.21fF
C50606 OR2X1_LOC_158/A OR2X1_LOC_485/A 1.55fF
C50607 OR2X1_LOC_600/A AND2X1_LOC_374/Y 0.00fF
C50608 OR2X1_LOC_18/Y OR2X1_LOC_762/Y 0.07fF
C50609 OR2X1_LOC_36/Y AND2X1_LOC_447/Y 0.03fF
C50610 AND2X1_LOC_565/B AND2X1_LOC_569/A 0.01fF
C50611 OR2X1_LOC_251/a_36_216# OR2X1_LOC_278/Y 0.00fF
C50612 OR2X1_LOC_600/A OR2X1_LOC_52/B 0.13fF
C50613 OR2X1_LOC_518/Y AND2X1_LOC_831/Y 0.13fF
C50614 AND2X1_LOC_367/B GATE_366 0.83fF
C50615 OR2X1_LOC_458/B OR2X1_LOC_161/A 0.02fF
C50616 AND2X1_LOC_716/Y OR2X1_LOC_48/B 0.07fF
C50617 AND2X1_LOC_675/Y OR2X1_LOC_189/A 0.26fF
C50618 OR2X1_LOC_380/a_8_216# OR2X1_LOC_588/Y 0.01fF
C50619 OR2X1_LOC_663/a_8_216# AND2X1_LOC_51/Y 0.01fF
C50620 OR2X1_LOC_804/A OR2X1_LOC_716/a_36_216# 0.00fF
C50621 AND2X1_LOC_395/a_8_24# OR2X1_LOC_78/Y 0.01fF
C50622 OR2X1_LOC_769/a_8_216# OR2X1_LOC_598/A 0.01fF
C50623 OR2X1_LOC_703/A OR2X1_LOC_375/A 0.00fF
C50624 OR2X1_LOC_815/a_8_216# OR2X1_LOC_89/A 0.01fF
C50625 OR2X1_LOC_687/Y OR2X1_LOC_678/a_36_216# 0.02fF
C50626 AND2X1_LOC_716/Y OR2X1_LOC_18/Y 0.07fF
C50627 AND2X1_LOC_753/B AND2X1_LOC_95/Y 0.07fF
C50628 AND2X1_LOC_489/Y OR2X1_LOC_600/A 0.03fF
C50629 OR2X1_LOC_691/A OR2X1_LOC_19/B 0.03fF
C50630 OR2X1_LOC_539/A OR2X1_LOC_377/A 0.02fF
C50631 OR2X1_LOC_687/Y AND2X1_LOC_41/A 0.07fF
C50632 AND2X1_LOC_654/Y OR2X1_LOC_48/B 0.07fF
C50633 OR2X1_LOC_448/B OR2X1_LOC_161/A 0.01fF
C50634 OR2X1_LOC_807/Y OR2X1_LOC_805/a_8_216# 0.05fF
C50635 OR2X1_LOC_634/A AND2X1_LOC_291/a_36_24# 0.02fF
C50636 OR2X1_LOC_634/a_36_216# AND2X1_LOC_824/B 0.00fF
C50637 AND2X1_LOC_858/B AND2X1_LOC_806/A 0.38fF
C50638 AND2X1_LOC_40/Y OR2X1_LOC_456/a_36_216# 0.03fF
C50639 AND2X1_LOC_343/a_8_24# OR2X1_LOC_51/Y 0.01fF
C50640 AND2X1_LOC_40/Y OR2X1_LOC_738/A 0.07fF
C50641 OR2X1_LOC_405/A OR2X1_LOC_737/A 1.24fF
C50642 OR2X1_LOC_347/a_8_216# AND2X1_LOC_95/Y 0.01fF
C50643 INPUT_5 OR2X1_LOC_11/Y 0.06fF
C50644 OR2X1_LOC_168/B OR2X1_LOC_449/B 0.02fF
C50645 OR2X1_LOC_185/A OR2X1_LOC_620/Y 0.07fF
C50646 AND2X1_LOC_456/B OR2X1_LOC_283/a_8_216# 0.01fF
C50647 OR2X1_LOC_807/Y OR2X1_LOC_362/B 0.01fF
C50648 OR2X1_LOC_723/B OR2X1_LOC_717/a_36_216# 0.02fF
C50649 AND2X1_LOC_76/Y OR2X1_LOC_619/Y 0.03fF
C50650 OR2X1_LOC_475/a_36_216# OR2X1_LOC_805/A -0.01fF
C50651 OR2X1_LOC_457/B OR2X1_LOC_464/A 0.03fF
C50652 AND2X1_LOC_658/B AND2X1_LOC_148/Y 0.05fF
C50653 AND2X1_LOC_12/Y OR2X1_LOC_856/B 0.09fF
C50654 OR2X1_LOC_405/A AND2X1_LOC_95/Y 8.69fF
C50655 AND2X1_LOC_738/B OR2X1_LOC_74/A 0.07fF
C50656 OR2X1_LOC_474/Y OR2X1_LOC_203/Y 0.07fF
C50657 OR2X1_LOC_318/Y OR2X1_LOC_799/a_8_216# 0.04fF
C50658 OR2X1_LOC_490/Y OR2X1_LOC_56/A 0.02fF
C50659 AND2X1_LOC_702/Y AND2X1_LOC_857/Y 0.36fF
C50660 OR2X1_LOC_89/A AND2X1_LOC_443/Y 0.14fF
C50661 AND2X1_LOC_357/B OR2X1_LOC_64/Y 0.01fF
C50662 OR2X1_LOC_185/A AND2X1_LOC_178/a_36_24# 0.00fF
C50663 OR2X1_LOC_74/A OR2X1_LOC_56/A 4.86fF
C50664 OR2X1_LOC_121/B OR2X1_LOC_182/B 0.03fF
C50665 AND2X1_LOC_799/a_36_24# AND2X1_LOC_810/Y 0.00fF
C50666 AND2X1_LOC_70/Y OR2X1_LOC_605/B 0.09fF
C50667 AND2X1_LOC_530/a_8_24# INPUT_1 0.03fF
C50668 OR2X1_LOC_755/A OR2X1_LOC_600/A 0.99fF
C50669 OR2X1_LOC_3/Y AND2X1_LOC_434/a_8_24# 0.02fF
C50670 OR2X1_LOC_841/a_8_216# OR2X1_LOC_841/B 0.06fF
C50671 OR2X1_LOC_851/A OR2X1_LOC_831/a_8_216# 0.03fF
C50672 OR2X1_LOC_45/B OR2X1_LOC_238/a_8_216# 0.02fF
C50673 OR2X1_LOC_328/a_8_216# OR2X1_LOC_3/Y 0.02fF
C50674 OR2X1_LOC_479/Y AND2X1_LOC_92/Y 0.73fF
C50675 AND2X1_LOC_47/Y AND2X1_LOC_277/a_8_24# 0.04fF
C50676 OR2X1_LOC_604/A AND2X1_LOC_849/A 0.02fF
C50677 OR2X1_LOC_524/Y AND2X1_LOC_147/Y 0.03fF
C50678 OR2X1_LOC_448/A OR2X1_LOC_269/B 0.01fF
C50679 OR2X1_LOC_666/Y AND2X1_LOC_861/B 0.10fF
C50680 OR2X1_LOC_217/A OR2X1_LOC_560/A 0.00fF
C50681 AND2X1_LOC_64/Y OR2X1_LOC_205/Y 0.03fF
C50682 OR2X1_LOC_651/A AND2X1_LOC_44/Y 0.00fF
C50683 OR2X1_LOC_494/Y OR2X1_LOC_64/Y 0.00fF
C50684 AND2X1_LOC_196/a_36_24# OR2X1_LOC_56/A 0.01fF
C50685 OR2X1_LOC_70/Y AND2X1_LOC_434/Y 0.03fF
C50686 OR2X1_LOC_382/Y AND2X1_LOC_259/Y 0.00fF
C50687 OR2X1_LOC_70/Y AND2X1_LOC_219/Y 0.07fF
C50688 OR2X1_LOC_485/A AND2X1_LOC_98/Y 0.16fF
C50689 AND2X1_LOC_318/Y OR2X1_LOC_428/A 0.03fF
C50690 OR2X1_LOC_589/Y AND2X1_LOC_592/a_8_24# -0.01fF
C50691 OR2X1_LOC_95/Y OR2X1_LOC_12/Y 0.06fF
C50692 OR2X1_LOC_36/Y AND2X1_LOC_649/B 0.29fF
C50693 OR2X1_LOC_261/A OR2X1_LOC_56/A 0.00fF
C50694 OR2X1_LOC_154/A OR2X1_LOC_185/A 0.03fF
C50695 AND2X1_LOC_707/a_36_24# OR2X1_LOC_64/Y 0.00fF
C50696 OR2X1_LOC_791/B OR2X1_LOC_375/A 0.04fF
C50697 OR2X1_LOC_778/Y AND2X1_LOC_422/a_8_24# 0.16fF
C50698 AND2X1_LOC_51/Y OR2X1_LOC_78/A 0.42fF
C50699 AND2X1_LOC_448/Y AND2X1_LOC_466/a_8_24# 0.09fF
C50700 OR2X1_LOC_532/B OR2X1_LOC_361/a_36_216# 0.01fF
C50701 OR2X1_LOC_160/A OR2X1_LOC_520/Y 0.03fF
C50702 VDD AND2X1_LOC_465/Y 0.16fF
C50703 OR2X1_LOC_154/A OR2X1_LOC_249/Y -0.02fF
C50704 OR2X1_LOC_404/Y OR2X1_LOC_78/B 0.81fF
C50705 OR2X1_LOC_805/A OR2X1_LOC_553/A 0.94fF
C50706 OR2X1_LOC_131/Y AND2X1_LOC_141/A 0.00fF
C50707 OR2X1_LOC_485/A OR2X1_LOC_594/Y 0.13fF
C50708 OR2X1_LOC_450/a_8_216# AND2X1_LOC_425/Y 0.01fF
C50709 OR2X1_LOC_450/B AND2X1_LOC_694/a_8_24# 0.20fF
C50710 OR2X1_LOC_185/A OR2X1_LOC_267/A 0.01fF
C50711 AND2X1_LOC_474/a_8_24# OR2X1_LOC_44/Y 0.01fF
C50712 OR2X1_LOC_116/A OR2X1_LOC_203/Y 0.01fF
C50713 OR2X1_LOC_276/B OR2X1_LOC_549/A 1.56fF
C50714 OR2X1_LOC_339/a_8_216# OR2X1_LOC_814/A 0.03fF
C50715 OR2X1_LOC_168/B OR2X1_LOC_121/B 0.03fF
C50716 OR2X1_LOC_193/Y OR2X1_LOC_375/A 0.26fF
C50717 AND2X1_LOC_175/B OR2X1_LOC_26/Y 0.06fF
C50718 OR2X1_LOC_619/Y OR2X1_LOC_52/B 2.26fF
C50719 AND2X1_LOC_571/B AND2X1_LOC_657/A 0.02fF
C50720 AND2X1_LOC_56/B OR2X1_LOC_241/a_8_216# 0.01fF
C50721 AND2X1_LOC_347/B AND2X1_LOC_866/A 0.02fF
C50722 AND2X1_LOC_538/a_8_24# AND2X1_LOC_434/Y 0.03fF
C50723 OR2X1_LOC_97/A OR2X1_LOC_544/a_8_216# 0.02fF
C50724 OR2X1_LOC_155/A OR2X1_LOC_161/A 0.31fF
C50725 OR2X1_LOC_26/Y AND2X1_LOC_848/Y 0.05fF
C50726 OR2X1_LOC_462/B OR2X1_LOC_87/B 0.03fF
C50727 OR2X1_LOC_364/A OR2X1_LOC_185/Y 0.07fF
C50728 OR2X1_LOC_494/Y OR2X1_LOC_417/A 4.62fF
C50729 AND2X1_LOC_859/B AND2X1_LOC_860/A 0.00fF
C50730 OR2X1_LOC_217/Y OR2X1_LOC_203/Y 0.01fF
C50731 VDD OR2X1_LOC_408/Y 0.12fF
C50732 OR2X1_LOC_247/Y AND2X1_LOC_248/a_8_24# 0.00fF
C50733 AND2X1_LOC_363/Y OR2X1_LOC_417/A 0.03fF
C50734 AND2X1_LOC_41/A OR2X1_LOC_643/Y 0.03fF
C50735 OR2X1_LOC_404/Y OR2X1_LOC_721/Y 0.00fF
C50736 OR2X1_LOC_290/a_8_216# OR2X1_LOC_416/Y 0.01fF
C50737 AND2X1_LOC_48/A OR2X1_LOC_174/A 0.01fF
C50738 AND2X1_LOC_852/Y OR2X1_LOC_85/A 0.12fF
C50739 OR2X1_LOC_262/a_8_216# OR2X1_LOC_36/Y 0.05fF
C50740 AND2X1_LOC_728/Y AND2X1_LOC_191/Y 0.03fF
C50741 AND2X1_LOC_331/a_36_24# AND2X1_LOC_51/Y 0.00fF
C50742 OR2X1_LOC_89/A AND2X1_LOC_848/Y 0.03fF
C50743 OR2X1_LOC_605/A OR2X1_LOC_161/A 0.01fF
C50744 OR2X1_LOC_633/a_8_216# D_INPUT_0 0.01fF
C50745 INPUT_0 AND2X1_LOC_28/a_8_24# 0.03fF
C50746 AND2X1_LOC_582/a_8_24# AND2X1_LOC_425/Y 0.01fF
C50747 OR2X1_LOC_283/Y OR2X1_LOC_26/Y 0.06fF
C50748 AND2X1_LOC_307/a_8_24# OR2X1_LOC_48/B 0.01fF
C50749 OR2X1_LOC_777/B OR2X1_LOC_308/Y 0.03fF
C50750 OR2X1_LOC_91/A AND2X1_LOC_831/Y 0.07fF
C50751 OR2X1_LOC_89/a_8_216# OR2X1_LOC_44/Y 0.01fF
C50752 OR2X1_LOC_22/Y OR2X1_LOC_92/Y 0.39fF
C50753 OR2X1_LOC_251/Y OR2X1_LOC_667/a_36_216# 0.02fF
C50754 AND2X1_LOC_377/a_8_24# OR2X1_LOC_46/A 0.11fF
C50755 AND2X1_LOC_637/Y AND2X1_LOC_638/a_8_24# 0.13fF
C50756 OR2X1_LOC_701/Y AND2X1_LOC_663/B 0.21fF
C50757 OR2X1_LOC_51/Y AND2X1_LOC_675/a_8_24# 0.05fF
C50758 AND2X1_LOC_486/Y AND2X1_LOC_477/A 0.06fF
C50759 OR2X1_LOC_64/Y AND2X1_LOC_843/a_36_24# 0.01fF
C50760 OR2X1_LOC_404/Y OR2X1_LOC_375/A 0.06fF
C50761 OR2X1_LOC_401/a_8_216# OR2X1_LOC_402/Y 0.05fF
C50762 OR2X1_LOC_602/A AND2X1_LOC_51/Y 0.04fF
C50763 AND2X1_LOC_554/B OR2X1_LOC_117/Y 0.04fF
C50764 OR2X1_LOC_512/Y OR2X1_LOC_713/A 0.03fF
C50765 OR2X1_LOC_291/Y OR2X1_LOC_32/B 0.07fF
C50766 AND2X1_LOC_40/Y OR2X1_LOC_288/A 0.00fF
C50767 AND2X1_LOC_59/Y OR2X1_LOC_121/B 1.87fF
C50768 OR2X1_LOC_662/A OR2X1_LOC_643/Y 0.06fF
C50769 AND2X1_LOC_95/Y OR2X1_LOC_285/Y 0.01fF
C50770 OR2X1_LOC_36/Y AND2X1_LOC_729/B 0.03fF
C50771 OR2X1_LOC_485/A AND2X1_LOC_602/a_36_24# 0.00fF
C50772 OR2X1_LOC_419/Y AND2X1_LOC_447/Y 0.01fF
C50773 AND2X1_LOC_12/Y OR2X1_LOC_383/Y 0.04fF
C50774 OR2X1_LOC_22/Y OR2X1_LOC_65/B 0.03fF
C50775 OR2X1_LOC_624/A OR2X1_LOC_814/A 0.10fF
C50776 OR2X1_LOC_782/a_8_216# OR2X1_LOC_161/A 0.14fF
C50777 OR2X1_LOC_675/A OR2X1_LOC_719/Y 0.43fF
C50778 AND2X1_LOC_663/B OR2X1_LOC_44/Y 0.04fF
C50779 AND2X1_LOC_41/A OR2X1_LOC_786/Y 0.07fF
C50780 OR2X1_LOC_358/a_36_216# OR2X1_LOC_476/B 0.00fF
C50781 OR2X1_LOC_52/B AND2X1_LOC_201/a_8_24# 0.01fF
C50782 OR2X1_LOC_754/A OR2X1_LOC_7/A 0.09fF
C50783 AND2X1_LOC_729/Y OR2X1_LOC_601/a_36_216# 0.00fF
C50784 AND2X1_LOC_51/Y OR2X1_LOC_155/A 0.38fF
C50785 OR2X1_LOC_291/A OR2X1_LOC_74/A 0.03fF
C50786 AND2X1_LOC_91/B OR2X1_LOC_579/A 0.33fF
C50787 INPUT_0 OR2X1_LOC_311/a_8_216# 0.01fF
C50788 AND2X1_LOC_856/A AND2X1_LOC_856/a_8_24# 0.19fF
C50789 AND2X1_LOC_123/Y AND2X1_LOC_845/Y 0.01fF
C50790 OR2X1_LOC_186/Y OR2X1_LOC_317/B 0.00fF
C50791 OR2X1_LOC_685/a_8_216# AND2X1_LOC_425/Y 0.01fF
C50792 OR2X1_LOC_647/Y OR2X1_LOC_646/A 0.95fF
C50793 OR2X1_LOC_19/B OR2X1_LOC_86/a_8_216# 0.01fF
C50794 OR2X1_LOC_769/B OR2X1_LOC_598/A 0.03fF
C50795 AND2X1_LOC_91/B OR2X1_LOC_844/B 0.29fF
C50796 OR2X1_LOC_566/A OR2X1_LOC_308/Y 0.07fF
C50797 OR2X1_LOC_271/Y OR2X1_LOC_22/Y 0.02fF
C50798 OR2X1_LOC_527/Y OR2X1_LOC_371/Y 0.28fF
C50799 AND2X1_LOC_345/Y OR2X1_LOC_481/A 0.14fF
C50800 OR2X1_LOC_804/A OR2X1_LOC_776/a_8_216# 0.04fF
C50801 OR2X1_LOC_391/B OR2X1_LOC_773/a_8_216# 0.01fF
C50802 AND2X1_LOC_675/A OR2X1_LOC_39/A 0.20fF
C50803 OR2X1_LOC_274/Y OR2X1_LOC_241/B 0.00fF
C50804 AND2X1_LOC_663/B AND2X1_LOC_116/Y 0.03fF
C50805 AND2X1_LOC_662/a_8_24# AND2X1_LOC_276/Y 0.19fF
C50806 AND2X1_LOC_51/Y OR2X1_LOC_392/a_8_216# 0.01fF
C50807 AND2X1_LOC_42/a_8_24# OR2X1_LOC_19/B 0.06fF
C50808 OR2X1_LOC_709/A OR2X1_LOC_515/Y 0.01fF
C50809 OR2X1_LOC_62/B OR2X1_LOC_585/A 0.05fF
C50810 AND2X1_LOC_40/Y AND2X1_LOC_72/B 0.31fF
C50811 OR2X1_LOC_431/a_8_216# OR2X1_LOC_304/Y 0.01fF
C50812 AND2X1_LOC_849/a_8_24# OR2X1_LOC_44/Y 0.00fF
C50813 AND2X1_LOC_92/Y OR2X1_LOC_68/B 0.10fF
C50814 OR2X1_LOC_421/Y OR2X1_LOC_424/Y 0.05fF
C50815 OR2X1_LOC_140/B OR2X1_LOC_115/B 0.59fF
C50816 OR2X1_LOC_185/A OR2X1_LOC_84/a_8_216# 0.04fF
C50817 GATE_811 AND2X1_LOC_624/A 0.15fF
C50818 VDD AND2X1_LOC_268/a_8_24# 0.00fF
C50819 OR2X1_LOC_52/a_36_216# OR2X1_LOC_52/Y 0.00fF
C50820 OR2X1_LOC_92/Y OR2X1_LOC_387/a_8_216# 0.01fF
C50821 OR2X1_LOC_673/B AND2X1_LOC_36/Y 0.02fF
C50822 OR2X1_LOC_83/a_8_216# OR2X1_LOC_46/A 0.01fF
C50823 OR2X1_LOC_45/B OR2X1_LOC_696/A 0.12fF
C50824 OR2X1_LOC_472/a_36_216# OR2X1_LOC_476/B -0.01fF
C50825 AND2X1_LOC_91/a_36_24# OR2X1_LOC_605/Y 0.00fF
C50826 OR2X1_LOC_145/a_36_216# OR2X1_LOC_146/Y 0.00fF
C50827 OR2X1_LOC_831/A AND2X1_LOC_36/Y 0.20fF
C50828 OR2X1_LOC_865/Y D_INPUT_1 0.02fF
C50829 OR2X1_LOC_109/Y OR2X1_LOC_419/Y 0.09fF
C50830 OR2X1_LOC_40/Y OR2X1_LOC_142/Y 0.14fF
C50831 AND2X1_LOC_122/a_8_24# D_INPUT_0 0.01fF
C50832 AND2X1_LOC_36/Y OR2X1_LOC_515/A 0.01fF
C50833 OR2X1_LOC_185/A OR2X1_LOC_739/Y 0.11fF
C50834 OR2X1_LOC_325/B OR2X1_LOC_374/a_8_216# 0.00fF
C50835 OR2X1_LOC_66/A OR2X1_LOC_537/a_8_216# 0.02fF
C50836 OR2X1_LOC_673/Y D_INPUT_1 0.07fF
C50837 OR2X1_LOC_598/Y AND2X1_LOC_36/Y 0.17fF
C50838 OR2X1_LOC_680/A AND2X1_LOC_795/Y 0.70fF
C50839 VDD OR2X1_LOC_174/Y 0.04fF
C50840 OR2X1_LOC_151/A OR2X1_LOC_388/a_8_216# 0.00fF
C50841 OR2X1_LOC_108/Y OR2X1_LOC_183/a_8_216# 0.03fF
C50842 AND2X1_LOC_838/B AND2X1_LOC_838/a_8_24# 0.19fF
C50843 OR2X1_LOC_272/Y OR2X1_LOC_95/Y 0.02fF
C50844 AND2X1_LOC_359/B AND2X1_LOC_721/A 0.20fF
C50845 OR2X1_LOC_427/A AND2X1_LOC_563/Y 0.03fF
C50846 OR2X1_LOC_217/a_36_216# OR2X1_LOC_786/Y 0.01fF
C50847 OR2X1_LOC_46/A OR2X1_LOC_77/a_36_216# 0.01fF
C50848 AND2X1_LOC_110/Y OR2X1_LOC_319/Y 0.01fF
C50849 OR2X1_LOC_292/Y OR2X1_LOC_437/A 0.02fF
C50850 OR2X1_LOC_275/a_8_216# OR2X1_LOC_31/Y 0.09fF
C50851 AND2X1_LOC_64/Y OR2X1_LOC_851/B 0.01fF
C50852 OR2X1_LOC_827/Y AND2X1_LOC_838/B 0.10fF
C50853 OR2X1_LOC_589/A AND2X1_LOC_772/Y 0.25fF
C50854 OR2X1_LOC_516/Y VDD 0.40fF
C50855 AND2X1_LOC_711/A OR2X1_LOC_759/Y 0.24fF
C50856 AND2X1_LOC_170/B AND2X1_LOC_802/a_8_24# 0.14fF
C50857 OR2X1_LOC_91/Y AND2X1_LOC_222/Y 0.08fF
C50858 OR2X1_LOC_778/Y OR2X1_LOC_493/Y 0.45fF
C50859 AND2X1_LOC_571/B VDD 0.24fF
C50860 AND2X1_LOC_785/Y AND2X1_LOC_786/Y 0.02fF
C50861 AND2X1_LOC_541/Y OR2X1_LOC_106/Y 0.07fF
C50862 OR2X1_LOC_696/A AND2X1_LOC_705/a_8_24# -0.01fF
C50863 OR2X1_LOC_51/Y OR2X1_LOC_387/A 0.01fF
C50864 OR2X1_LOC_186/Y AND2X1_LOC_44/Y 0.02fF
C50865 AND2X1_LOC_715/Y OR2X1_LOC_329/a_36_216# -0.01fF
C50866 OR2X1_LOC_804/a_8_216# OR2X1_LOC_593/B 0.01fF
C50867 AND2X1_LOC_539/Y AND2X1_LOC_535/Y 0.47fF
C50868 AND2X1_LOC_707/Y OR2X1_LOC_421/Y 1.30fF
C50869 OR2X1_LOC_136/a_8_216# OR2X1_LOC_40/Y 0.01fF
C50870 OR2X1_LOC_364/A AND2X1_LOC_432/a_8_24# 0.02fF
C50871 AND2X1_LOC_753/B AND2X1_LOC_41/Y 0.01fF
C50872 OR2X1_LOC_352/A OR2X1_LOC_212/B 0.19fF
C50873 OR2X1_LOC_486/Y OR2X1_LOC_161/B 3.33fF
C50874 OR2X1_LOC_48/B OR2X1_LOC_13/B 0.57fF
C50875 OR2X1_LOC_6/B OR2X1_LOC_139/A 0.10fF
C50876 OR2X1_LOC_539/A OR2X1_LOC_539/B 0.12fF
C50877 AND2X1_LOC_801/B OR2X1_LOC_95/Y 0.01fF
C50878 OR2X1_LOC_189/Y AND2X1_LOC_222/Y 0.03fF
C50879 OR2X1_LOC_469/Y OR2X1_LOC_469/B 0.00fF
C50880 OR2X1_LOC_18/Y OR2X1_LOC_13/B 0.35fF
C50881 INPUT_1 AND2X1_LOC_476/A 0.04fF
C50882 OR2X1_LOC_69/Y OR2X1_LOC_80/A 0.00fF
C50883 AND2X1_LOC_40/Y AND2X1_LOC_36/Y 1.80fF
C50884 OR2X1_LOC_810/A AND2X1_LOC_31/Y 0.06fF
C50885 OR2X1_LOC_307/a_8_216# AND2X1_LOC_31/Y 0.01fF
C50886 OR2X1_LOC_64/Y AND2X1_LOC_204/Y 0.09fF
C50887 OR2X1_LOC_319/B OR2X1_LOC_354/a_8_216# 0.04fF
C50888 OR2X1_LOC_87/A OR2X1_LOC_446/B 0.02fF
C50889 OR2X1_LOC_316/Y OR2X1_LOC_300/Y 0.01fF
C50890 AND2X1_LOC_227/Y OR2X1_LOC_503/Y 0.10fF
C50891 OR2X1_LOC_377/A OR2X1_LOC_771/B 0.14fF
C50892 OR2X1_LOC_87/A OR2X1_LOC_303/B 0.03fF
C50893 OR2X1_LOC_53/Y INPUT_0 0.02fF
C50894 OR2X1_LOC_544/A AND2X1_LOC_438/a_36_24# 0.00fF
C50895 OR2X1_LOC_51/Y AND2X1_LOC_636/a_36_24# 0.00fF
C50896 AND2X1_LOC_474/A AND2X1_LOC_284/a_8_24# 0.01fF
C50897 VDD OR2X1_LOC_162/Y 0.16fF
C50898 OR2X1_LOC_604/A AND2X1_LOC_346/a_8_24# 0.06fF
C50899 OR2X1_LOC_770/a_8_216# D_INPUT_1 0.02fF
C50900 AND2X1_LOC_810/A OR2X1_LOC_56/A 0.03fF
C50901 OR2X1_LOC_40/Y AND2X1_LOC_347/B 0.01fF
C50902 OR2X1_LOC_324/a_36_216# AND2X1_LOC_64/Y 0.00fF
C50903 AND2X1_LOC_70/Y OR2X1_LOC_549/A 0.16fF
C50904 OR2X1_LOC_160/B OR2X1_LOC_648/B 0.47fF
C50905 OR2X1_LOC_97/A OR2X1_LOC_634/a_8_216# 0.01fF
C50906 OR2X1_LOC_309/a_8_216# OR2X1_LOC_426/B 0.01fF
C50907 OR2X1_LOC_696/A AND2X1_LOC_435/a_8_24# 0.05fF
C50908 OR2X1_LOC_518/Y OR2X1_LOC_519/Y 0.00fF
C50909 OR2X1_LOC_637/A AND2X1_LOC_829/a_36_24# 0.00fF
C50910 OR2X1_LOC_530/Y OR2X1_LOC_437/A -0.00fF
C50911 AND2X1_LOC_41/A AND2X1_LOC_255/a_8_24# 0.06fF
C50912 OR2X1_LOC_9/Y OR2X1_LOC_51/Y 0.05fF
C50913 AND2X1_LOC_787/A AND2X1_LOC_733/a_8_24# 0.01fF
C50914 AND2X1_LOC_91/B OR2X1_LOC_865/B 0.02fF
C50915 AND2X1_LOC_753/B AND2X1_LOC_22/Y 0.07fF
C50916 OR2X1_LOC_604/A AND2X1_LOC_447/Y 0.10fF
C50917 AND2X1_LOC_719/Y AND2X1_LOC_190/a_36_24# 0.06fF
C50918 AND2X1_LOC_64/Y OR2X1_LOC_160/A 0.49fF
C50919 OR2X1_LOC_124/A OR2X1_LOC_641/A 0.00fF
C50920 OR2X1_LOC_124/B OR2X1_LOC_124/a_8_216# 0.03fF
C50921 OR2X1_LOC_56/A AND2X1_LOC_254/a_8_24# 0.03fF
C50922 OR2X1_LOC_303/a_36_216# OR2X1_LOC_212/A 0.00fF
C50923 OR2X1_LOC_741/Y OR2X1_LOC_190/a_36_216# 0.03fF
C50924 OR2X1_LOC_375/A OR2X1_LOC_718/a_8_216# 0.01fF
C50925 OR2X1_LOC_45/B OR2X1_LOC_695/a_8_216# 0.02fF
C50926 OR2X1_LOC_56/A AND2X1_LOC_860/A 0.03fF
C50927 OR2X1_LOC_362/B OR2X1_LOC_362/a_8_216# 0.07fF
C50928 OR2X1_LOC_369/Y VDD 0.14fF
C50929 OR2X1_LOC_297/Y AND2X1_LOC_789/Y 0.01fF
C50930 OR2X1_LOC_604/A OR2X1_LOC_743/a_36_216# 0.00fF
C50931 AND2X1_LOC_241/a_8_24# OR2X1_LOC_39/A 0.03fF
C50932 OR2X1_LOC_405/A AND2X1_LOC_22/Y 0.03fF
C50933 OR2X1_LOC_850/a_36_216# OR2X1_LOC_362/A 0.00fF
C50934 AND2X1_LOC_544/Y AND2X1_LOC_811/a_8_24# 0.00fF
C50935 OR2X1_LOC_49/A OR2X1_LOC_427/A 0.10fF
C50936 OR2X1_LOC_45/B AND2X1_LOC_717/a_8_24# 0.04fF
C50937 AND2X1_LOC_43/B OR2X1_LOC_121/A 0.03fF
C50938 AND2X1_LOC_345/Y AND2X1_LOC_789/Y 0.40fF
C50939 OR2X1_LOC_379/Y OR2X1_LOC_691/Y 0.43fF
C50940 AND2X1_LOC_716/Y AND2X1_LOC_181/Y 0.02fF
C50941 OR2X1_LOC_847/A OR2X1_LOC_633/A 0.03fF
C50942 OR2X1_LOC_114/a_8_216# VDD 0.21fF
C50943 OR2X1_LOC_43/A AND2X1_LOC_772/Y 0.43fF
C50944 AND2X1_LOC_47/a_8_24# AND2X1_LOC_44/Y 0.02fF
C50945 AND2X1_LOC_421/a_8_24# OR2X1_LOC_307/A 0.20fF
C50946 OR2X1_LOC_244/Y AND2X1_LOC_245/a_36_24# 0.00fF
C50947 AND2X1_LOC_658/B AND2X1_LOC_545/a_8_24# 0.03fF
C50948 OR2X1_LOC_185/A OR2X1_LOC_435/A 0.17fF
C50949 AND2X1_LOC_540/a_8_24# OR2X1_LOC_108/Y 0.01fF
C50950 GATE_479 AND2X1_LOC_223/a_8_24# 0.20fF
C50951 OR2X1_LOC_45/B AND2X1_LOC_458/Y 0.01fF
C50952 OR2X1_LOC_316/Y AND2X1_LOC_219/A 0.00fF
C50953 D_INPUT_3 OR2X1_LOC_68/B 4.00fF
C50954 OR2X1_LOC_40/Y AND2X1_LOC_737/a_36_24# 0.00fF
C50955 AND2X1_LOC_91/B OR2X1_LOC_403/B 0.04fF
C50956 OR2X1_LOC_177/Y OR2X1_LOC_109/Y 0.60fF
C50957 OR2X1_LOC_325/Y OR2X1_LOC_703/A 0.03fF
C50958 AND2X1_LOC_81/B AND2X1_LOC_44/Y 0.03fF
C50959 OR2X1_LOC_437/a_36_216# AND2X1_LOC_222/Y 0.00fF
C50960 OR2X1_LOC_45/B OR2X1_LOC_271/B 0.01fF
C50961 OR2X1_LOC_851/a_8_216# OR2X1_LOC_840/A 0.01fF
C50962 OR2X1_LOC_53/Y OR2X1_LOC_690/A 0.25fF
C50963 OR2X1_LOC_405/A OR2X1_LOC_729/a_36_216# 0.00fF
C50964 AND2X1_LOC_64/Y OR2X1_LOC_624/B 0.07fF
C50965 AND2X1_LOC_586/a_8_24# OR2X1_LOC_598/Y 0.24fF
C50966 AND2X1_LOC_94/Y AND2X1_LOC_401/Y 0.04fF
C50967 OR2X1_LOC_813/a_8_216# OR2X1_LOC_278/Y 0.01fF
C50968 OR2X1_LOC_128/a_8_216# OR2X1_LOC_151/A 0.02fF
C50969 AND2X1_LOC_555/Y OR2X1_LOC_282/a_36_216# 0.00fF
C50970 OR2X1_LOC_470/a_8_216# OR2X1_LOC_161/B 0.01fF
C50971 AND2X1_LOC_72/a_8_24# OR2X1_LOC_563/A 0.02fF
C50972 AND2X1_LOC_850/Y AND2X1_LOC_860/A 0.09fF
C50973 OR2X1_LOC_6/B AND2X1_LOC_573/A 0.01fF
C50974 OR2X1_LOC_604/A OR2X1_LOC_109/Y 0.10fF
C50975 OR2X1_LOC_648/A OR2X1_LOC_785/B 0.01fF
C50976 OR2X1_LOC_841/a_8_216# OR2X1_LOC_168/B -0.01fF
C50977 OR2X1_LOC_160/A AND2X1_LOC_86/a_8_24# 0.01fF
C50978 OR2X1_LOC_539/A OR2X1_LOC_78/B 0.00fF
C50979 OR2X1_LOC_439/a_8_216# OR2X1_LOC_544/B 0.04fF
C50980 AND2X1_LOC_721/Y OR2X1_LOC_485/A 0.07fF
C50981 AND2X1_LOC_533/a_8_24# AND2X1_LOC_110/Y 0.01fF
C50982 OR2X1_LOC_585/A OR2X1_LOC_585/a_36_216# 0.02fF
C50983 OR2X1_LOC_532/B OR2X1_LOC_523/A 0.01fF
C50984 OR2X1_LOC_604/A AND2X1_LOC_448/Y 0.00fF
C50985 OR2X1_LOC_585/A OR2X1_LOC_15/a_36_216# 0.00fF
C50986 AND2X1_LOC_554/Y OR2X1_LOC_600/A 0.07fF
C50987 OR2X1_LOC_181/B OR2X1_LOC_741/Y 0.04fF
C50988 OR2X1_LOC_116/a_8_216# OR2X1_LOC_549/A 0.04fF
C50989 OR2X1_LOC_753/Y OR2X1_LOC_754/Y 0.20fF
C50990 OR2X1_LOC_269/B OR2X1_LOC_390/A 0.03fF
C50991 OR2X1_LOC_354/A OR2X1_LOC_703/A 0.28fF
C50992 AND2X1_LOC_76/a_8_24# OR2X1_LOC_59/Y 0.02fF
C50993 OR2X1_LOC_363/B OR2X1_LOC_362/B 0.12fF
C50994 D_GATE_662 OR2X1_LOC_849/A 0.00fF
C50995 OR2X1_LOC_312/Y AND2X1_LOC_810/B 0.07fF
C50996 OR2X1_LOC_774/B OR2X1_LOC_80/A 0.14fF
C50997 OR2X1_LOC_175/B OR2X1_LOC_538/A 0.03fF
C50998 OR2X1_LOC_624/A OR2X1_LOC_244/Y 0.88fF
C50999 AND2X1_LOC_728/Y AND2X1_LOC_658/B 0.14fF
C51000 AND2X1_LOC_3/Y AND2X1_LOC_279/a_8_24# 0.01fF
C51001 AND2X1_LOC_593/a_8_24# OR2X1_LOC_36/Y 0.04fF
C51002 AND2X1_LOC_99/Y OR2X1_LOC_517/A 0.08fF
C51003 OR2X1_LOC_3/Y AND2X1_LOC_786/Y 0.07fF
C51004 AND2X1_LOC_161/Y OR2X1_LOC_619/Y 0.01fF
C51005 AND2X1_LOC_41/A OR2X1_LOC_725/B 0.07fF
C51006 OR2X1_LOC_754/A OR2X1_LOC_753/a_8_216# 0.48fF
C51007 OR2X1_LOC_474/Y OR2X1_LOC_721/Y 0.10fF
C51008 AND2X1_LOC_557/Y AND2X1_LOC_563/A 0.09fF
C51009 AND2X1_LOC_82/Y AND2X1_LOC_86/B 0.03fF
C51010 OR2X1_LOC_97/A OR2X1_LOC_602/a_36_216# 0.00fF
C51011 OR2X1_LOC_496/Y AND2X1_LOC_499/a_8_24# 0.11fF
C51012 OR2X1_LOC_519/Y OR2X1_LOC_91/A 0.16fF
C51013 AND2X1_LOC_392/A OR2X1_LOC_44/Y 0.07fF
C51014 AND2X1_LOC_217/Y AND2X1_LOC_361/A 0.02fF
C51015 OR2X1_LOC_482/Y OR2X1_LOC_665/Y 0.62fF
C51016 OR2X1_LOC_482/a_36_216# OR2X1_LOC_666/Y 0.00fF
C51017 OR2X1_LOC_40/Y OR2X1_LOC_262/Y 0.04fF
C51018 AND2X1_LOC_82/Y OR2X1_LOC_624/B 0.00fF
C51019 OR2X1_LOC_72/Y AND2X1_LOC_203/a_8_24# 0.09fF
C51020 OR2X1_LOC_541/A OR2X1_LOC_541/B 0.16fF
C51021 OR2X1_LOC_219/a_8_216# AND2X1_LOC_92/Y 0.04fF
C51022 OR2X1_LOC_744/A AND2X1_LOC_633/a_8_24# 0.01fF
C51023 OR2X1_LOC_756/B OR2X1_LOC_362/B 0.16fF
C51024 OR2X1_LOC_482/Y OR2X1_LOC_485/A 0.09fF
C51025 OR2X1_LOC_51/Y AND2X1_LOC_834/a_36_24# 0.00fF
C51026 OR2X1_LOC_40/Y OR2X1_LOC_238/Y 0.00fF
C51027 AND2X1_LOC_191/Y AND2X1_LOC_480/A 0.03fF
C51028 OR2X1_LOC_216/Y OR2X1_LOC_78/A 0.19fF
C51029 OR2X1_LOC_516/Y OR2X1_LOC_674/Y 0.12fF
C51030 AND2X1_LOC_86/B AND2X1_LOC_86/a_8_24# 0.06fF
C51031 OR2X1_LOC_71/A OR2X1_LOC_398/Y -0.01fF
C51032 OR2X1_LOC_51/Y AND2X1_LOC_852/Y 0.03fF
C51033 OR2X1_LOC_196/B AND2X1_LOC_44/Y 0.04fF
C51034 OR2X1_LOC_160/A OR2X1_LOC_656/Y 0.02fF
C51035 AND2X1_LOC_663/B OR2X1_LOC_382/A 0.03fF
C51036 OR2X1_LOC_280/Y OR2X1_LOC_600/A 0.10fF
C51037 AND2X1_LOC_578/A AND2X1_LOC_500/B 0.03fF
C51038 OR2X1_LOC_841/a_8_216# AND2X1_LOC_59/Y 0.01fF
C51039 AND2X1_LOC_392/A AND2X1_LOC_116/Y 0.03fF
C51040 OR2X1_LOC_116/A OR2X1_LOC_721/Y 0.20fF
C51041 AND2X1_LOC_366/A OR2X1_LOC_44/Y 0.01fF
C51042 AND2X1_LOC_41/A OR2X1_LOC_204/Y 0.09fF
C51043 OR2X1_LOC_474/Y OR2X1_LOC_375/A 0.03fF
C51044 AND2X1_LOC_692/a_8_24# AND2X1_LOC_44/Y 0.01fF
C51045 OR2X1_LOC_374/Y AND2X1_LOC_591/a_8_24# 0.02fF
C51046 OR2X1_LOC_256/Y AND2X1_LOC_342/Y 0.05fF
C51047 OR2X1_LOC_866/a_8_216# OR2X1_LOC_391/A 0.09fF
C51048 OR2X1_LOC_92/Y OR2X1_LOC_39/A 0.10fF
C51049 OR2X1_LOC_417/A AND2X1_LOC_241/a_36_24# 0.01fF
C51050 OR2X1_LOC_557/A OR2X1_LOC_66/A 0.00fF
C51051 AND2X1_LOC_662/B AND2X1_LOC_841/B 0.09fF
C51052 OR2X1_LOC_26/Y OR2X1_LOC_26/a_8_216# -0.00fF
C51053 OR2X1_LOC_692/Y OR2X1_LOC_22/Y 0.03fF
C51054 AND2X1_LOC_633/Y OR2X1_LOC_16/A 0.03fF
C51055 VDD AND2X1_LOC_42/B 1.64fF
C51056 OR2X1_LOC_39/Y OR2X1_LOC_36/Y 0.01fF
C51057 VDD AND2X1_LOC_651/B 0.17fF
C51058 AND2X1_LOC_513/a_8_24# OR2X1_LOC_36/Y 0.03fF
C51059 OR2X1_LOC_287/A AND2X1_LOC_3/Y 0.80fF
C51060 OR2X1_LOC_680/Y AND2X1_LOC_657/Y 0.03fF
C51061 OR2X1_LOC_769/A AND2X1_LOC_3/Y 0.00fF
C51062 AND2X1_LOC_541/a_36_24# OR2X1_LOC_95/Y 0.01fF
C51063 OR2X1_LOC_348/Y AND2X1_LOC_281/a_8_24# 0.02fF
C51064 AND2X1_LOC_729/Y OR2X1_LOC_485/a_36_216# 0.00fF
C51065 AND2X1_LOC_59/Y OR2X1_LOC_856/B 0.09fF
C51066 OR2X1_LOC_756/B AND2X1_LOC_385/a_8_24# 0.11fF
C51067 AND2X1_LOC_729/B AND2X1_LOC_207/B 0.01fF
C51068 D_INPUT_0 OR2X1_LOC_16/A 0.14fF
C51069 VDD OR2X1_LOC_705/Y 0.00fF
C51070 OR2X1_LOC_529/Y AND2X1_LOC_858/B 0.03fF
C51071 AND2X1_LOC_228/Y AND2X1_LOC_654/Y 0.00fF
C51072 OR2X1_LOC_61/a_8_216# OR2X1_LOC_358/B 0.01fF
C51073 OR2X1_LOC_653/Y OR2X1_LOC_130/A 0.06fF
C51074 OR2X1_LOC_664/Y OR2X1_LOC_811/A 0.01fF
C51075 OR2X1_LOC_97/A OR2X1_LOC_440/A 0.04fF
C51076 OR2X1_LOC_675/A OR2X1_LOC_66/A 0.00fF
C51077 OR2X1_LOC_377/A OR2X1_LOC_402/Y 0.15fF
C51078 AND2X1_LOC_580/B AND2X1_LOC_866/B 0.02fF
C51079 OR2X1_LOC_174/A AND2X1_LOC_3/Y 0.05fF
C51080 AND2X1_LOC_196/a_8_24# OR2X1_LOC_59/Y 0.02fF
C51081 AND2X1_LOC_449/Y AND2X1_LOC_452/Y 0.03fF
C51082 AND2X1_LOC_50/Y AND2X1_LOC_51/A 0.01fF
C51083 INPUT_5 AND2X1_LOC_44/a_8_24# 0.05fF
C51084 AND2X1_LOC_47/Y OR2X1_LOC_740/B 3.98fF
C51085 OR2X1_LOC_783/A OR2X1_LOC_161/B 0.01fF
C51086 OR2X1_LOC_65/B OR2X1_LOC_39/A 0.02fF
C51087 AND2X1_LOC_95/Y OR2X1_LOC_653/A 0.04fF
C51088 AND2X1_LOC_339/B OR2X1_LOC_31/Y 0.08fF
C51089 OR2X1_LOC_473/a_36_216# OR2X1_LOC_810/A 0.12fF
C51090 OR2X1_LOC_140/A OR2X1_LOC_62/B 0.00fF
C51091 OR2X1_LOC_70/Y OR2X1_LOC_674/a_8_216# 0.03fF
C51092 AND2X1_LOC_211/B OR2X1_LOC_92/Y 0.07fF
C51093 OR2X1_LOC_600/A OR2X1_LOC_22/Y 0.20fF
C51094 OR2X1_LOC_294/a_36_216# OR2X1_LOC_296/Y 0.00fF
C51095 OR2X1_LOC_574/A OR2X1_LOC_574/a_8_216# 0.02fF
C51096 AND2X1_LOC_95/Y OR2X1_LOC_673/Y 0.03fF
C51097 OR2X1_LOC_814/A AND2X1_LOC_265/a_36_24# 0.01fF
C51098 OR2X1_LOC_479/Y AND2X1_LOC_526/a_36_24# 0.01fF
C51099 OR2X1_LOC_667/Y OR2X1_LOC_669/Y 0.04fF
C51100 OR2X1_LOC_113/Y OR2X1_LOC_404/Y 0.00fF
C51101 AND2X1_LOC_91/B OR2X1_LOC_493/Y 0.21fF
C51102 AND2X1_LOC_580/A AND2X1_LOC_624/A 0.15fF
C51103 AND2X1_LOC_714/a_8_24# AND2X1_LOC_648/B 0.01fF
C51104 OR2X1_LOC_756/B OR2X1_LOC_846/B 0.00fF
C51105 OR2X1_LOC_217/Y OR2X1_LOC_375/A 0.01fF
C51106 INPUT_7 OR2X1_LOC_17/a_36_216# 0.00fF
C51107 AND2X1_LOC_277/a_8_24# D_INPUT_1 0.01fF
C51108 AND2X1_LOC_259/Y OR2X1_LOC_427/A 0.00fF
C51109 OR2X1_LOC_219/a_36_216# OR2X1_LOC_222/A 0.00fF
C51110 VDD OR2X1_LOC_286/B 0.21fF
C51111 AND2X1_LOC_364/Y AND2X1_LOC_514/Y 0.96fF
C51112 OR2X1_LOC_271/Y OR2X1_LOC_39/A 0.13fF
C51113 OR2X1_LOC_250/Y OR2X1_LOC_106/A 0.02fF
C51114 OR2X1_LOC_117/a_8_216# OR2X1_LOC_67/Y 0.01fF
C51115 OR2X1_LOC_680/A AND2X1_LOC_834/a_36_24# 0.00fF
C51116 OR2X1_LOC_137/Y OR2X1_LOC_137/B 0.80fF
C51117 AND2X1_LOC_174/a_8_24# OR2X1_LOC_7/A 0.02fF
C51118 OR2X1_LOC_7/A OR2X1_LOC_118/Y 0.03fF
C51119 OR2X1_LOC_139/A OR2X1_LOC_598/A 0.10fF
C51120 AND2X1_LOC_56/B OR2X1_LOC_87/A 5.13fF
C51121 AND2X1_LOC_356/B AND2X1_LOC_356/a_8_24# 0.09fF
C51122 OR2X1_LOC_76/Y OR2X1_LOC_457/B 0.00fF
C51123 OR2X1_LOC_70/Y AND2X1_LOC_76/a_8_24# 0.05fF
C51124 INPUT_0 INPUT_1 7.14fF
C51125 OR2X1_LOC_30/a_8_216# OR2X1_LOC_17/Y 0.40fF
C51126 AND2X1_LOC_170/B AND2X1_LOC_436/Y 0.02fF
C51127 AND2X1_LOC_727/A OR2X1_LOC_594/a_8_216# 0.01fF
C51128 OR2X1_LOC_641/B AND2X1_LOC_226/a_36_24# 0.00fF
C51129 OR2X1_LOC_831/a_8_216# OR2X1_LOC_155/A 0.01fF
C51130 OR2X1_LOC_756/B OR2X1_LOC_471/Y 0.23fF
C51131 OR2X1_LOC_205/a_8_216# OR2X1_LOC_124/Y 0.39fF
C51132 OR2X1_LOC_203/Y OR2X1_LOC_217/a_8_216# 0.02fF
C51133 AND2X1_LOC_660/a_8_24# OR2X1_LOC_59/Y 0.01fF
C51134 OR2X1_LOC_426/B AND2X1_LOC_451/Y 0.00fF
C51135 AND2X1_LOC_208/a_8_24# D_INPUT_0 0.01fF
C51136 AND2X1_LOC_748/a_8_24# OR2X1_LOC_193/A 0.17fF
C51137 OR2X1_LOC_710/a_8_216# OR2X1_LOC_269/B 0.09fF
C51138 OR2X1_LOC_91/Y OR2X1_LOC_74/A 0.26fF
C51139 OR2X1_LOC_121/B OR2X1_LOC_794/A 0.02fF
C51140 OR2X1_LOC_3/Y AND2X1_LOC_124/a_36_24# 0.01fF
C51141 AND2X1_LOC_343/a_8_24# AND2X1_LOC_359/B 0.00fF
C51142 OR2X1_LOC_154/A OR2X1_LOC_702/A 0.10fF
C51143 AND2X1_LOC_454/A OR2X1_LOC_52/B 0.02fF
C51144 OR2X1_LOC_774/Y OR2X1_LOC_810/A 0.08fF
C51145 AND2X1_LOC_777/a_8_24# OR2X1_LOC_3/Y 0.03fF
C51146 OR2X1_LOC_306/Y AND2X1_LOC_729/B 0.03fF
C51147 OR2X1_LOC_185/A OR2X1_LOC_476/a_8_216# 0.00fF
C51148 OR2X1_LOC_312/Y OR2X1_LOC_585/A 0.02fF
C51149 AND2X1_LOC_784/A AND2X1_LOC_566/Y 0.02fF
C51150 OR2X1_LOC_815/a_8_216# AND2X1_LOC_792/Y 0.01fF
C51151 OR2X1_LOC_95/Y OR2X1_LOC_594/a_8_216# 0.07fF
C51152 OR2X1_LOC_160/A OR2X1_LOC_206/A 0.03fF
C51153 AND2X1_LOC_727/A AND2X1_LOC_468/B 0.04fF
C51154 OR2X1_LOC_774/Y OR2X1_LOC_864/a_8_216# 0.03fF
C51155 OR2X1_LOC_675/a_8_216# OR2X1_LOC_76/Y 0.13fF
C51156 AND2X1_LOC_367/A D_INPUT_3 0.03fF
C51157 OR2X1_LOC_22/Y OR2X1_LOC_619/Y 0.14fF
C51158 AND2X1_LOC_698/a_8_24# OR2X1_LOC_738/A 0.04fF
C51159 AND2X1_LOC_95/Y AND2X1_LOC_309/a_8_24# 0.02fF
C51160 OR2X1_LOC_499/B OR2X1_LOC_276/B 0.02fF
C51161 OR2X1_LOC_70/a_8_216# OR2X1_LOC_2/Y 0.08fF
C51162 AND2X1_LOC_564/a_8_24# OR2X1_LOC_527/Y 0.01fF
C51163 OR2X1_LOC_628/a_8_216# OR2X1_LOC_417/A 0.14fF
C51164 AND2X1_LOC_260/a_8_24# OR2X1_LOC_820/B 0.01fF
C51165 AND2X1_LOC_91/B OR2X1_LOC_532/a_8_216# 0.05fF
C51166 OR2X1_LOC_154/A OR2X1_LOC_476/B 0.13fF
C51167 OR2X1_LOC_814/A OR2X1_LOC_161/A 0.02fF
C51168 AND2X1_LOC_197/a_36_24# OR2X1_LOC_6/A 0.00fF
C51169 OR2X1_LOC_715/B AND2X1_LOC_31/Y 3.89fF
C51170 AND2X1_LOC_794/B OR2X1_LOC_533/A 0.01fF
C51171 OR2X1_LOC_92/Y OR2X1_LOC_760/a_8_216# 0.06fF
C51172 OR2X1_LOC_605/A OR2X1_LOC_787/Y 0.02fF
C51173 AND2X1_LOC_703/a_8_24# OR2X1_LOC_95/Y 0.01fF
C51174 AND2X1_LOC_755/a_8_24# OR2X1_LOC_286/B 0.20fF
C51175 OR2X1_LOC_715/B OR2X1_LOC_715/a_8_216# 0.02fF
C51176 OR2X1_LOC_611/a_8_216# OR2X1_LOC_6/A 0.10fF
C51177 AND2X1_LOC_793/Y AND2X1_LOC_663/A 0.10fF
C51178 AND2X1_LOC_51/Y OR2X1_LOC_68/a_8_216# 0.01fF
C51179 OR2X1_LOC_243/B OR2X1_LOC_375/A 0.03fF
C51180 AND2X1_LOC_51/Y OR2X1_LOC_710/a_36_216# 0.00fF
C51181 AND2X1_LOC_537/Y OR2X1_LOC_6/A 0.07fF
C51182 OR2X1_LOC_427/A AND2X1_LOC_810/Y 0.06fF
C51183 OR2X1_LOC_3/Y OR2X1_LOC_481/a_8_216# 0.07fF
C51184 AND2X1_LOC_31/Y OR2X1_LOC_543/A 0.03fF
C51185 OR2X1_LOC_36/Y OR2X1_LOC_46/A 3.86fF
C51186 OR2X1_LOC_485/A OR2X1_LOC_304/Y 0.00fF
C51187 AND2X1_LOC_31/Y OR2X1_LOC_784/B 0.02fF
C51188 AND2X1_LOC_580/B AND2X1_LOC_664/a_8_24# 0.18fF
C51189 AND2X1_LOC_468/B OR2X1_LOC_95/Y 0.14fF
C51190 AND2X1_LOC_742/a_8_24# AND2X1_LOC_742/A 0.03fF
C51191 OR2X1_LOC_750/A OR2X1_LOC_269/B 0.01fF
C51192 OR2X1_LOC_235/B OR2X1_LOC_86/A 0.04fF
C51193 OR2X1_LOC_261/Y AND2X1_LOC_663/B 0.26fF
C51194 AND2X1_LOC_436/Y OR2X1_LOC_331/Y 0.00fF
C51195 OR2X1_LOC_527/Y OR2X1_LOC_74/A 0.07fF
C51196 AND2X1_LOC_344/a_8_24# AND2X1_LOC_721/A 0.01fF
C51197 AND2X1_LOC_810/B OR2X1_LOC_13/B 0.01fF
C51198 VDD AND2X1_LOC_793/B 0.06fF
C51199 AND2X1_LOC_64/Y OR2X1_LOC_130/Y 0.00fF
C51200 OR2X1_LOC_337/a_8_216# OR2X1_LOC_365/B 0.00fF
C51201 OR2X1_LOC_56/A AND2X1_LOC_562/Y 0.03fF
C51202 OR2X1_LOC_483/a_8_216# OR2X1_LOC_532/B 0.03fF
C51203 AND2X1_LOC_482/a_8_24# OR2X1_LOC_270/Y 0.01fF
C51204 AND2X1_LOC_631/Y AND2X1_LOC_632/a_8_24# 0.01fF
C51205 AND2X1_LOC_537/Y OR2X1_LOC_299/a_8_216# 0.12fF
C51206 VDD OR2X1_LOC_533/A 0.21fF
C51207 AND2X1_LOC_243/Y OR2X1_LOC_71/A 0.06fF
C51208 OR2X1_LOC_291/Y OR2X1_LOC_74/A 0.49fF
C51209 OR2X1_LOC_665/Y OR2X1_LOC_628/Y 0.07fF
C51210 AND2X1_LOC_539/a_8_24# OR2X1_LOC_52/B 0.02fF
C51211 INPUT_1 OR2X1_LOC_690/A 0.63fF
C51212 OR2X1_LOC_161/B OR2X1_LOC_374/a_36_216# 0.01fF
C51213 AND2X1_LOC_631/a_36_24# AND2X1_LOC_620/Y 0.00fF
C51214 OR2X1_LOC_812/B D_INPUT_1 0.01fF
C51215 OR2X1_LOC_402/B OR2X1_LOC_68/B 0.01fF
C51216 AND2X1_LOC_227/Y OR2X1_LOC_36/Y 0.03fF
C51217 AND2X1_LOC_728/Y OR2X1_LOC_47/Y 0.03fF
C51218 OR2X1_LOC_74/A AND2X1_LOC_574/A 0.03fF
C51219 OR2X1_LOC_161/B OR2X1_LOC_308/Y 0.07fF
C51220 OR2X1_LOC_748/a_8_216# OR2X1_LOC_748/Y -0.00fF
C51221 OR2X1_LOC_620/a_8_216# AND2X1_LOC_36/Y 0.03fF
C51222 OR2X1_LOC_613/Y GATE_662 0.03fF
C51223 OR2X1_LOC_76/B OR2X1_LOC_76/a_8_216# 0.05fF
C51224 OR2X1_LOC_487/a_8_216# OR2X1_LOC_71/Y 0.01fF
C51225 AND2X1_LOC_110/Y OR2X1_LOC_777/B 0.02fF
C51226 D_INPUT_3 AND2X1_LOC_673/a_8_24# 0.01fF
C51227 OR2X1_LOC_814/A AND2X1_LOC_51/Y 2.15fF
C51228 AND2X1_LOC_573/A OR2X1_LOC_598/A 0.04fF
C51229 OR2X1_LOC_484/a_36_216# OR2X1_LOC_437/A 0.00fF
C51230 OR2X1_LOC_502/A OR2X1_LOC_724/A 0.07fF
C51231 OR2X1_LOC_582/Y AND2X1_LOC_635/a_8_24# 0.01fF
C51232 AND2X1_LOC_191/Y AND2X1_LOC_479/Y 0.10fF
C51233 OR2X1_LOC_696/A OR2X1_LOC_158/A 0.32fF
C51234 OR2X1_LOC_490/Y D_INPUT_3 0.04fF
C51235 D_INPUT_3 OR2X1_LOC_74/A 0.02fF
C51236 AND2X1_LOC_539/Y OR2X1_LOC_16/A 0.13fF
C51237 OR2X1_LOC_22/Y OR2X1_LOC_22/A 0.02fF
C51238 OR2X1_LOC_743/A AND2X1_LOC_648/B 0.02fF
C51239 OR2X1_LOC_557/A OR2X1_LOC_84/A -0.00fF
C51240 OR2X1_LOC_70/Y AND2X1_LOC_479/Y 0.00fF
C51241 OR2X1_LOC_78/B OR2X1_LOC_771/B 0.11fF
C51242 OR2X1_LOC_157/a_8_216# OR2X1_LOC_70/A 0.01fF
C51243 AND2X1_LOC_42/B OR2X1_LOC_845/A 0.37fF
C51244 AND2X1_LOC_31/Y OR2X1_LOC_215/Y 0.01fF
C51245 OR2X1_LOC_754/A OR2X1_LOC_615/Y 0.26fF
C51246 AND2X1_LOC_7/B AND2X1_LOC_256/a_36_24# 0.00fF
C51247 OR2X1_LOC_36/Y OR2X1_LOC_753/Y 0.07fF
C51248 AND2X1_LOC_280/a_8_24# OR2X1_LOC_269/B 0.01fF
C51249 OR2X1_LOC_45/a_36_216# OR2X1_LOC_172/Y 0.00fF
C51250 AND2X1_LOC_715/Y OR2X1_LOC_158/A 0.07fF
C51251 OR2X1_LOC_53/Y AND2X1_LOC_195/a_36_24# 0.00fF
C51252 AND2X1_LOC_358/Y OR2X1_LOC_12/Y 0.02fF
C51253 AND2X1_LOC_778/a_8_24# OR2X1_LOC_406/A 0.01fF
C51254 OR2X1_LOC_136/Y AND2X1_LOC_566/B 0.01fF
C51255 OR2X1_LOC_151/A AND2X1_LOC_7/B 0.07fF
C51256 INPUT_1 OR2X1_LOC_417/A 0.45fF
C51257 OR2X1_LOC_617/Y AND2X1_LOC_792/Y 0.17fF
C51258 OR2X1_LOC_105/a_8_216# OR2X1_LOC_579/A 0.09fF
C51259 OR2X1_LOC_87/A AND2X1_LOC_427/a_8_24# 0.04fF
C51260 OR2X1_LOC_59/Y AND2X1_LOC_792/a_8_24# 0.02fF
C51261 OR2X1_LOC_92/Y AND2X1_LOC_247/a_36_24# 0.00fF
C51262 OR2X1_LOC_16/A AND2X1_LOC_771/B 0.03fF
C51263 AND2X1_LOC_12/Y OR2X1_LOC_366/Y 0.01fF
C51264 AND2X1_LOC_40/Y OR2X1_LOC_469/B 0.01fF
C51265 OR2X1_LOC_737/A OR2X1_LOC_723/B 0.09fF
C51266 OR2X1_LOC_696/A AND2X1_LOC_98/Y 0.01fF
C51267 OR2X1_LOC_45/B AND2X1_LOC_392/A 0.03fF
C51268 OR2X1_LOC_59/Y AND2X1_LOC_773/a_8_24# 0.01fF
C51269 OR2X1_LOC_362/A OR2X1_LOC_843/B 0.01fF
C51270 AND2X1_LOC_387/a_8_24# AND2X1_LOC_44/Y 0.03fF
C51271 OR2X1_LOC_106/Y OR2X1_LOC_744/A 0.08fF
C51272 OR2X1_LOC_27/Y OR2X1_LOC_598/A 0.01fF
C51273 OR2X1_LOC_3/Y OR2X1_LOC_88/a_8_216# 0.01fF
C51274 OR2X1_LOC_126/a_36_216# OR2X1_LOC_744/A -0.00fF
C51275 OR2X1_LOC_44/Y OR2X1_LOC_589/Y 0.03fF
C51276 OR2X1_LOC_3/Y OR2X1_LOC_172/a_8_216# 0.00fF
C51277 AND2X1_LOC_787/A OR2X1_LOC_51/Y 0.04fF
C51278 OR2X1_LOC_696/A OR2X1_LOC_103/Y 1.07fF
C51279 AND2X1_LOC_558/a_8_24# OR2X1_LOC_428/A 0.17fF
C51280 OR2X1_LOC_70/A OR2X1_LOC_762/a_8_216# 0.00fF
C51281 AND2X1_LOC_22/Y AND2X1_LOC_19/Y 2.57fF
C51282 OR2X1_LOC_66/A OR2X1_LOC_548/a_8_216# 0.02fF
C51283 AND2X1_LOC_367/B OR2X1_LOC_428/A 0.25fF
C51284 AND2X1_LOC_137/a_8_24# AND2X1_LOC_139/A 0.01fF
C51285 OR2X1_LOC_291/Y AND2X1_LOC_647/Y 0.01fF
C51286 OR2X1_LOC_375/A OR2X1_LOC_771/B 0.08fF
C51287 AND2X1_LOC_391/a_8_24# AND2X1_LOC_555/Y 0.01fF
C51288 OR2X1_LOC_3/Y OR2X1_LOC_378/A 0.05fF
C51289 AND2X1_LOC_503/a_8_24# OR2X1_LOC_502/Y 0.00fF
C51290 OR2X1_LOC_62/A AND2X1_LOC_672/a_8_24# 0.02fF
C51291 OR2X1_LOC_375/A OR2X1_LOC_209/A 0.02fF
C51292 AND2X1_LOC_43/B AND2X1_LOC_36/Y 0.19fF
C51293 AND2X1_LOC_773/Y OR2X1_LOC_59/Y 0.01fF
C51294 AND2X1_LOC_689/a_8_24# AND2X1_LOC_31/Y 0.01fF
C51295 OR2X1_LOC_696/A OR2X1_LOC_103/a_8_216# 0.01fF
C51296 OR2X1_LOC_46/A OR2X1_LOC_28/a_36_216# 0.00fF
C51297 AND2X1_LOC_67/a_8_24# AND2X1_LOC_7/B 0.04fF
C51298 OR2X1_LOC_502/A OR2X1_LOC_415/Y 0.02fF
C51299 OR2X1_LOC_585/A OR2X1_LOC_599/a_36_216# 0.00fF
C51300 OR2X1_LOC_329/B AND2X1_LOC_786/Y 0.09fF
C51301 OR2X1_LOC_820/a_8_216# OR2X1_LOC_600/A 0.01fF
C51302 AND2X1_LOC_851/B OR2X1_LOC_47/Y 0.04fF
C51303 OR2X1_LOC_585/A OR2X1_LOC_13/B 1.20fF
C51304 OR2X1_LOC_56/A OR2X1_LOC_381/a_8_216# 0.01fF
C51305 OR2X1_LOC_323/A AND2X1_LOC_841/B 0.00fF
C51306 OR2X1_LOC_185/A OR2X1_LOC_605/Y 0.02fF
C51307 OR2X1_LOC_528/Y OR2X1_LOC_759/A 0.03fF
C51308 AND2X1_LOC_480/a_8_24# GATE_479 0.01fF
C51309 OR2X1_LOC_375/A OR2X1_LOC_776/A 0.00fF
C51310 OR2X1_LOC_612/Y OR2X1_LOC_16/A 0.02fF
C51311 AND2X1_LOC_657/Y AND2X1_LOC_476/Y 0.10fF
C51312 OR2X1_LOC_369/a_8_216# OR2X1_LOC_40/Y 0.02fF
C51313 OR2X1_LOC_862/B OR2X1_LOC_349/A 0.01fF
C51314 OR2X1_LOC_368/a_8_216# VDD 0.21fF
C51315 OR2X1_LOC_78/A OR2X1_LOC_439/B 0.01fF
C51316 OR2X1_LOC_481/A OR2X1_LOC_384/Y 0.04fF
C51317 AND2X1_LOC_64/Y OR2X1_LOC_447/A 0.09fF
C51318 VDD OR2X1_LOC_581/Y -0.00fF
C51319 AND2X1_LOC_22/Y D_INPUT_4 0.00fF
C51320 AND2X1_LOC_227/Y OR2X1_LOC_419/Y 0.05fF
C51321 AND2X1_LOC_555/Y OR2X1_LOC_127/a_8_216# 0.01fF
C51322 AND2X1_LOC_22/Y AND2X1_LOC_615/a_36_24# 0.00fF
C51323 OR2X1_LOC_565/A OR2X1_LOC_192/A 0.05fF
C51324 OR2X1_LOC_721/a_36_216# OR2X1_LOC_721/Y 0.00fF
C51325 OR2X1_LOC_164/Y OR2X1_LOC_373/Y 0.03fF
C51326 OR2X1_LOC_499/a_8_216# OR2X1_LOC_140/B 0.01fF
C51327 OR2X1_LOC_228/a_8_216# AND2X1_LOC_52/Y 0.47fF
C51328 OR2X1_LOC_195/A AND2X1_LOC_41/Y 0.23fF
C51329 OR2X1_LOC_710/B VDD 0.21fF
C51330 OR2X1_LOC_59/Y AND2X1_LOC_243/Y 0.00fF
C51331 AND2X1_LOC_651/a_8_24# OR2X1_LOC_12/Y 0.01fF
C51332 OR2X1_LOC_524/Y AND2X1_LOC_477/Y 0.10fF
C51333 AND2X1_LOC_403/a_8_24# AND2X1_LOC_404/B 0.01fF
C51334 AND2X1_LOC_95/Y OR2X1_LOC_720/Y 0.01fF
C51335 OR2X1_LOC_113/Y OR2X1_LOC_362/A 0.13fF
C51336 OR2X1_LOC_695/Y OR2X1_LOC_51/Y 0.01fF
C51337 AND2X1_LOC_831/Y AND2X1_LOC_222/Y 0.07fF
C51338 OR2X1_LOC_813/A OR2X1_LOC_88/Y 0.22fF
C51339 OR2X1_LOC_817/a_8_216# AND2X1_LOC_789/Y 0.01fF
C51340 VDD AND2X1_LOC_468/a_8_24# -0.00fF
C51341 OR2X1_LOC_474/Y OR2X1_LOC_549/A 0.07fF
C51342 OR2X1_LOC_48/B OR2X1_LOC_428/A 0.53fF
C51343 OR2X1_LOC_405/a_36_216# AND2X1_LOC_7/B 0.00fF
C51344 OR2X1_LOC_170/A OR2X1_LOC_170/a_8_216# 0.39fF
C51345 VDD OR2X1_LOC_363/A 0.19fF
C51346 OR2X1_LOC_319/B OR2X1_LOC_151/A 0.11fF
C51347 OR2X1_LOC_97/A OR2X1_LOC_661/a_36_216# 0.00fF
C51348 OR2X1_LOC_768/A OR2X1_LOC_66/A 0.01fF
C51349 VDD OR2X1_LOC_778/a_8_216# 0.21fF
C51350 OR2X1_LOC_18/Y OR2X1_LOC_428/A 0.18fF
C51351 OR2X1_LOC_468/Y OR2X1_LOC_170/a_36_216# 0.00fF
C51352 OR2X1_LOC_80/a_8_216# OR2X1_LOC_80/A 0.02fF
C51353 AND2X1_LOC_848/Y AND2X1_LOC_287/B 0.03fF
C51354 OR2X1_LOC_45/Y OR2X1_LOC_135/Y 0.10fF
C51355 AND2X1_LOC_702/a_36_24# OR2X1_LOC_428/A 0.00fF
C51356 OR2X1_LOC_813/Y OR2X1_LOC_85/a_8_216# 0.02fF
C51357 AND2X1_LOC_194/a_36_24# AND2X1_LOC_194/Y 0.00fF
C51358 OR2X1_LOC_399/A OR2X1_LOC_16/A 0.11fF
C51359 AND2X1_LOC_82/Y OR2X1_LOC_847/A 0.03fF
C51360 OR2X1_LOC_318/Y OR2X1_LOC_151/A 0.02fF
C51361 AND2X1_LOC_186/a_8_24# OR2X1_LOC_816/A 0.01fF
C51362 OR2X1_LOC_199/a_36_216# AND2X1_LOC_43/B 0.01fF
C51363 OR2X1_LOC_52/B AND2X1_LOC_783/B 0.03fF
C51364 OR2X1_LOC_18/Y OR2X1_LOC_595/A 0.14fF
C51365 AND2X1_LOC_621/Y OR2X1_LOC_12/Y 0.12fF
C51366 OR2X1_LOC_121/B OR2X1_LOC_716/a_36_216# 0.00fF
C51367 VDD OR2X1_LOC_663/A 0.11fF
C51368 AND2X1_LOC_714/B OR2X1_LOC_427/A 0.03fF
C51369 OR2X1_LOC_121/Y OR2X1_LOC_624/A 0.10fF
C51370 OR2X1_LOC_769/A INPUT_0 0.01fF
C51371 AND2X1_LOC_22/Y OR2X1_LOC_653/A 0.04fF
C51372 AND2X1_LOC_548/Y AND2X1_LOC_663/A 0.43fF
C51373 OR2X1_LOC_160/A OR2X1_LOC_185/a_8_216# 0.02fF
C51374 AND2X1_LOC_70/Y OR2X1_LOC_499/B 0.01fF
C51375 AND2X1_LOC_22/Y OR2X1_LOC_673/Y 0.10fF
C51376 OR2X1_LOC_536/Y OR2X1_LOC_92/Y 0.04fF
C51377 AND2X1_LOC_711/Y AND2X1_LOC_792/a_8_24# 0.01fF
C51378 AND2X1_LOC_41/A OR2X1_LOC_78/A 0.92fF
C51379 VDD AND2X1_LOC_503/a_8_24# -0.00fF
C51380 AND2X1_LOC_539/Y AND2X1_LOC_336/a_8_24# 0.01fF
C51381 AND2X1_LOC_564/B OR2X1_LOC_312/Y 0.01fF
C51382 OR2X1_LOC_116/A OR2X1_LOC_549/A 0.04fF
C51383 AND2X1_LOC_698/a_8_24# AND2X1_LOC_36/Y 0.01fF
C51384 AND2X1_LOC_266/Y AND2X1_LOC_249/a_8_24# 0.01fF
C51385 OR2X1_LOC_97/A OR2X1_LOC_778/Y 0.05fF
C51386 OR2X1_LOC_203/Y AND2X1_LOC_256/a_8_24# 0.01fF
C51387 OR2X1_LOC_312/Y OR2X1_LOC_368/Y 0.01fF
C51388 OR2X1_LOC_151/A OR2X1_LOC_805/A 0.10fF
C51389 INPUT_0 OR2X1_LOC_517/A 0.00fF
C51390 AND2X1_LOC_3/Y OR2X1_LOC_563/A 0.39fF
C51391 OR2X1_LOC_215/a_8_216# OR2X1_LOC_68/B 0.02fF
C51392 OR2X1_LOC_217/Y OR2X1_LOC_549/A 0.03fF
C51393 AND2X1_LOC_647/Y AND2X1_LOC_656/a_8_24# 0.11fF
C51394 AND2X1_LOC_367/A OR2X1_LOC_494/a_8_216# 0.01fF
C51395 OR2X1_LOC_6/B OR2X1_LOC_32/B 0.03fF
C51396 AND2X1_LOC_729/Y OR2X1_LOC_329/Y 0.03fF
C51397 OR2X1_LOC_780/A OR2X1_LOC_712/B 0.00fF
C51398 AND2X1_LOC_722/Y OR2X1_LOC_164/Y 0.02fF
C51399 AND2X1_LOC_796/Y OR2X1_LOC_437/A 0.01fF
C51400 AND2X1_LOC_22/Y OR2X1_LOC_195/A 0.08fF
C51401 OR2X1_LOC_385/Y OR2X1_LOC_428/A 0.03fF
C51402 OR2X1_LOC_198/a_8_216# OR2X1_LOC_19/B 0.01fF
C51403 OR2X1_LOC_612/a_8_216# OR2X1_LOC_39/A 0.06fF
C51404 INPUT_0 AND2X1_LOC_619/B 0.10fF
C51405 OR2X1_LOC_160/A OR2X1_LOC_776/Y 0.07fF
C51406 AND2X1_LOC_474/A OR2X1_LOC_92/Y 0.34fF
C51407 OR2X1_LOC_421/a_8_216# OR2X1_LOC_92/Y 0.03fF
C51408 OR2X1_LOC_600/A OR2X1_LOC_39/A 0.13fF
C51409 AND2X1_LOC_41/A OR2X1_LOC_448/B 0.00fF
C51410 AND2X1_LOC_648/B OR2X1_LOC_589/a_36_216# -0.00fF
C51411 AND2X1_LOC_447/Y AND2X1_LOC_447/a_8_24# 0.01fF
C51412 AND2X1_LOC_741/Y AND2X1_LOC_191/Y 0.03fF
C51413 OR2X1_LOC_161/A OR2X1_LOC_244/Y 0.90fF
C51414 OR2X1_LOC_715/B OR2X1_LOC_809/a_8_216# 0.71fF
C51415 AND2X1_LOC_654/B OR2X1_LOC_763/a_8_216# 0.47fF
C51416 OR2X1_LOC_158/A OR2X1_LOC_32/Y 0.13fF
C51417 OR2X1_LOC_571/B OR2X1_LOC_632/Y 0.08fF
C51418 OR2X1_LOC_402/Y OR2X1_LOC_78/B 0.27fF
C51419 OR2X1_LOC_185/Y VDD 2.10fF
C51420 OR2X1_LOC_324/B OR2X1_LOC_739/A 0.01fF
C51421 OR2X1_LOC_358/a_8_216# AND2X1_LOC_70/Y 0.01fF
C51422 INPUT_5 OR2X1_LOC_2/Y 0.02fF
C51423 OR2X1_LOC_847/A AND2X1_LOC_819/a_8_24# 0.01fF
C51424 AND2X1_LOC_820/a_8_24# AND2X1_LOC_820/B -0.00fF
C51425 OR2X1_LOC_501/B OR2X1_LOC_161/A 0.03fF
C51426 OR2X1_LOC_538/A OR2X1_LOC_624/A 0.18fF
C51427 AND2X1_LOC_857/Y AND2X1_LOC_654/Y 0.18fF
C51428 AND2X1_LOC_286/a_8_24# AND2X1_LOC_286/Y 0.00fF
C51429 VDD AND2X1_LOC_859/Y 0.71fF
C51430 OR2X1_LOC_703/B AND2X1_LOC_92/Y 0.10fF
C51431 OR2X1_LOC_722/a_8_216# OR2X1_LOC_733/A 0.01fF
C51432 AND2X1_LOC_662/B OR2X1_LOC_275/Y 0.01fF
C51433 OR2X1_LOC_851/a_36_216# OR2X1_LOC_87/A 0.00fF
C51434 OR2X1_LOC_151/A OR2X1_LOC_296/Y 0.08fF
C51435 OR2X1_LOC_678/a_8_216# OR2X1_LOC_375/A 0.01fF
C51436 OR2X1_LOC_856/B OR2X1_LOC_623/B 0.01fF
C51437 OR2X1_LOC_160/A OR2X1_LOC_756/B 0.10fF
C51438 OR2X1_LOC_160/A OR2X1_LOC_735/a_36_216# 0.01fF
C51439 OR2X1_LOC_744/A OR2X1_LOC_497/a_8_216# 0.04fF
C51440 OR2X1_LOC_87/A AND2X1_LOC_92/Y 0.09fF
C51441 AND2X1_LOC_211/B OR2X1_LOC_600/A 0.03fF
C51442 AND2X1_LOC_151/a_8_24# OR2X1_LOC_56/A -0.00fF
C51443 OR2X1_LOC_485/A AND2X1_LOC_539/a_36_24# 0.00fF
C51444 AND2X1_LOC_211/B AND2X1_LOC_335/Y 0.00fF
C51445 AND2X1_LOC_22/Y AND2X1_LOC_309/a_8_24# 0.10fF
C51446 AND2X1_LOC_508/B AND2X1_LOC_474/Y 0.00fF
C51447 OR2X1_LOC_19/B OR2X1_LOC_161/B 0.17fF
C51448 OR2X1_LOC_178/Y OR2X1_LOC_26/Y 0.06fF
C51449 OR2X1_LOC_631/B OR2X1_LOC_78/A 0.08fF
C51450 AND2X1_LOC_862/Y OR2X1_LOC_39/A 0.03fF
C51451 OR2X1_LOC_681/a_8_216# OR2X1_LOC_3/Y 0.01fF
C51452 AND2X1_LOC_687/A OR2X1_LOC_16/A 0.03fF
C51453 AND2X1_LOC_115/a_36_24# OR2X1_LOC_428/A 0.00fF
C51454 AND2X1_LOC_142/a_8_24# OR2X1_LOC_739/A 0.01fF
C51455 OR2X1_LOC_158/A AND2X1_LOC_663/B 0.06fF
C51456 AND2X1_LOC_508/a_8_24# AND2X1_LOC_474/Y -0.00fF
C51457 OR2X1_LOC_70/Y AND2X1_LOC_243/Y 0.02fF
C51458 OR2X1_LOC_620/Y OR2X1_LOC_623/a_8_216# 0.01fF
C51459 OR2X1_LOC_151/A OR2X1_LOC_436/a_8_216# 0.04fF
C51460 OR2X1_LOC_848/B OR2X1_LOC_391/a_36_216# 0.00fF
C51461 AND2X1_LOC_337/B AND2X1_LOC_337/a_8_24# 0.01fF
C51462 AND2X1_LOC_719/a_8_24# AND2X1_LOC_658/A 0.02fF
C51463 INPUT_0 OR2X1_LOC_827/a_8_216# 0.01fF
C51464 OR2X1_LOC_43/a_36_216# OR2X1_LOC_13/Y 0.00fF
C51465 OR2X1_LOC_541/A OR2X1_LOC_778/Y 0.01fF
C51466 AND2X1_LOC_722/A OR2X1_LOC_36/Y 0.01fF
C51467 OR2X1_LOC_808/a_8_216# OR2X1_LOC_375/A 0.01fF
C51468 OR2X1_LOC_311/Y OR2X1_LOC_13/a_36_216# 0.00fF
C51469 AND2X1_LOC_314/a_8_24# OR2X1_LOC_739/A 0.01fF
C51470 OR2X1_LOC_848/A OR2X1_LOC_392/A 0.01fF
C51471 AND2X1_LOC_721/Y OR2X1_LOC_238/a_8_216# 0.14fF
C51472 AND2X1_LOC_640/a_36_24# AND2X1_LOC_219/A 0.00fF
C51473 AND2X1_LOC_560/B OR2X1_LOC_517/A 4.39fF
C51474 AND2X1_LOC_91/B AND2X1_LOC_250/a_8_24# 0.15fF
C51475 OR2X1_LOC_92/Y OR2X1_LOC_85/A 0.18fF
C51476 OR2X1_LOC_35/B OR2X1_LOC_35/a_8_216# 0.05fF
C51477 AND2X1_LOC_41/A OR2X1_LOC_155/A 0.18fF
C51478 OR2X1_LOC_525/Y OR2X1_LOC_511/Y 0.22fF
C51479 OR2X1_LOC_31/Y AND2X1_LOC_219/A 0.00fF
C51480 AND2X1_LOC_365/A AND2X1_LOC_662/B 0.00fF
C51481 AND2X1_LOC_12/Y OR2X1_LOC_624/A 0.03fF
C51482 OR2X1_LOC_619/Y OR2X1_LOC_39/A 0.71fF
C51483 OR2X1_LOC_160/A OR2X1_LOC_660/B 0.00fF
C51484 OR2X1_LOC_643/A OR2X1_LOC_475/B 0.08fF
C51485 OR2X1_LOC_451/a_8_216# AND2X1_LOC_425/Y 0.02fF
C51486 AND2X1_LOC_83/a_8_24# OR2X1_LOC_532/B 0.01fF
C51487 AND2X1_LOC_578/A OR2X1_LOC_329/B 0.18fF
C51488 OR2X1_LOC_589/A AND2X1_LOC_800/a_8_24# 0.03fF
C51489 AND2X1_LOC_51/Y OR2X1_LOC_244/Y 0.06fF
C51490 OR2X1_LOC_756/B AND2X1_LOC_86/B 0.07fF
C51491 AND2X1_LOC_40/Y OR2X1_LOC_592/a_8_216# 0.01fF
C51492 AND2X1_LOC_568/B AND2X1_LOC_514/Y 0.77fF
C51493 AND2X1_LOC_352/B OR2X1_LOC_64/Y 0.01fF
C51494 OR2X1_LOC_485/A AND2X1_LOC_850/A 0.01fF
C51495 OR2X1_LOC_604/A OR2X1_LOC_46/A 0.04fF
C51496 OR2X1_LOC_158/A OR2X1_LOC_54/a_8_216# 0.02fF
C51497 AND2X1_LOC_123/Y OR2X1_LOC_67/A 0.01fF
C51498 AND2X1_LOC_721/a_8_24# OR2X1_LOC_669/Y 0.01fF
C51499 AND2X1_LOC_349/B OR2X1_LOC_256/Y 0.04fF
C51500 OR2X1_LOC_703/B AND2X1_LOC_166/a_8_24# 0.02fF
C51501 VDD OR2X1_LOC_472/B 0.12fF
C51502 AND2X1_LOC_186/a_8_24# AND2X1_LOC_807/Y 0.08fF
C51503 OR2X1_LOC_456/Y OR2X1_LOC_456/a_36_216# 0.00fF
C51504 OR2X1_LOC_481/A OR2X1_LOC_91/A 2.00fF
C51505 OR2X1_LOC_756/B OR2X1_LOC_624/B 0.02fF
C51506 AND2X1_LOC_51/Y OR2X1_LOC_715/A 0.03fF
C51507 AND2X1_LOC_454/Y AND2X1_LOC_466/a_8_24# 0.03fF
C51508 OR2X1_LOC_756/B OR2X1_LOC_33/a_8_216# 0.01fF
C51509 OR2X1_LOC_158/A AND2X1_LOC_849/a_8_24# 0.14fF
C51510 OR2X1_LOC_43/A OR2X1_LOC_278/Y 0.03fF
C51511 OR2X1_LOC_71/Y OR2X1_LOC_131/a_8_216# 0.01fF
C51512 OR2X1_LOC_849/a_8_216# OR2X1_LOC_244/Y 0.15fF
C51513 OR2X1_LOC_313/Y AND2X1_LOC_319/A 0.01fF
C51514 OR2X1_LOC_65/B OR2X1_LOC_85/A 0.06fF
C51515 OR2X1_LOC_88/A OR2X1_LOC_39/A 0.00fF
C51516 OR2X1_LOC_121/Y OR2X1_LOC_276/a_8_216# 0.05fF
C51517 OR2X1_LOC_520/B OR2X1_LOC_520/a_8_216# 0.07fF
C51518 OR2X1_LOC_380/A OR2X1_LOC_11/Y 0.01fF
C51519 OR2X1_LOC_283/Y AND2X1_LOC_843/a_8_24# 0.04fF
C51520 AND2X1_LOC_736/Y AND2X1_LOC_711/Y 0.03fF
C51521 AND2X1_LOC_98/Y AND2X1_LOC_663/B 0.10fF
C51522 OR2X1_LOC_160/B OR2X1_LOC_446/Y 0.15fF
C51523 AND2X1_LOC_36/Y OR2X1_LOC_367/B 0.20fF
C51524 OR2X1_LOC_348/Y OR2X1_LOC_288/A 0.00fF
C51525 AND2X1_LOC_736/Y OR2X1_LOC_70/Y 0.05fF
C51526 OR2X1_LOC_697/a_8_216# AND2X1_LOC_712/B 0.02fF
C51527 AND2X1_LOC_580/A OR2X1_LOC_613/Y 0.00fF
C51528 AND2X1_LOC_211/B OR2X1_LOC_619/Y 0.05fF
C51529 OR2X1_LOC_634/A AND2X1_LOC_119/a_8_24# 0.00fF
C51530 OR2X1_LOC_808/a_8_216# OR2X1_LOC_605/B 0.03fF
C51531 OR2X1_LOC_604/A AND2X1_LOC_227/Y 0.28fF
C51532 OR2X1_LOC_64/Y OR2X1_LOC_517/A 0.31fF
C51533 OR2X1_LOC_604/A OR2X1_LOC_604/a_36_216# 0.00fF
C51534 VDD OR2X1_LOC_852/A 0.12fF
C51535 AND2X1_LOC_621/Y OR2X1_LOC_239/a_8_216# 0.04fF
C51536 AND2X1_LOC_44/Y AND2X1_LOC_761/a_8_24# 0.04fF
C51537 OR2X1_LOC_375/A OR2X1_LOC_217/a_8_216# 0.01fF
C51538 OR2X1_LOC_121/B OR2X1_LOC_776/a_8_216# 0.02fF
C51539 AND2X1_LOC_805/a_36_24# GATE_579 0.00fF
C51540 OR2X1_LOC_599/A OR2X1_LOC_36/Y 0.35fF
C51541 OR2X1_LOC_147/B AND2X1_LOC_51/Y 0.02fF
C51542 AND2X1_LOC_387/B OR2X1_LOC_161/A 0.00fF
C51543 AND2X1_LOC_382/a_8_24# OR2X1_LOC_269/B 0.21fF
C51544 AND2X1_LOC_784/A AND2X1_LOC_702/Y 0.01fF
C51545 OR2X1_LOC_690/Y OR2X1_LOC_31/Y 0.02fF
C51546 OR2X1_LOC_51/Y AND2X1_LOC_675/A 0.00fF
C51547 AND2X1_LOC_8/Y AND2X1_LOC_29/a_8_24# 0.05fF
C51548 AND2X1_LOC_365/A AND2X1_LOC_337/B 0.03fF
C51549 AND2X1_LOC_858/B OR2X1_LOC_71/Y 0.03fF
C51550 OR2X1_LOC_91/A OR2X1_LOC_71/Y 0.03fF
C51551 OR2X1_LOC_64/Y AND2X1_LOC_833/a_8_24# 0.04fF
C51552 OR2X1_LOC_719/Y OR2X1_LOC_269/B 0.01fF
C51553 OR2X1_LOC_615/a_36_216# OR2X1_LOC_427/A 0.00fF
C51554 OR2X1_LOC_600/A OR2X1_LOC_826/Y 0.02fF
C51555 OR2X1_LOC_251/Y AND2X1_LOC_859/Y 0.23fF
C51556 OR2X1_LOC_317/A AND2X1_LOC_51/Y 0.04fF
C51557 AND2X1_LOC_349/a_8_24# OR2X1_LOC_7/A 0.01fF
C51558 AND2X1_LOC_563/a_36_24# AND2X1_LOC_489/Y 0.00fF
C51559 VDD AND2X1_LOC_798/A 0.21fF
C51560 AND2X1_LOC_229/a_8_24# OR2X1_LOC_641/B 0.01fF
C51561 D_INPUT_0 AND2X1_LOC_401/Y 0.03fF
C51562 OR2X1_LOC_635/a_36_216# AND2X1_LOC_51/Y 0.00fF
C51563 AND2X1_LOC_47/Y OR2X1_LOC_735/a_8_216# 0.02fF
C51564 OR2X1_LOC_498/Y AND2X1_LOC_474/Y 0.12fF
C51565 AND2X1_LOC_822/a_8_24# OR2X1_LOC_269/B 0.04fF
C51566 AND2X1_LOC_95/Y AND2X1_LOC_27/a_8_24# 0.01fF
C51567 OR2X1_LOC_154/A OR2X1_LOC_863/B 0.07fF
C51568 AND2X1_LOC_337/B OR2X1_LOC_43/A 0.01fF
C51569 OR2X1_LOC_124/B OR2X1_LOC_205/Y 0.83fF
C51570 AND2X1_LOC_81/a_8_24# OR2X1_LOC_633/B 0.01fF
C51571 OR2X1_LOC_74/A AND2X1_LOC_806/A 0.03fF
C51572 OR2X1_LOC_329/B AND2X1_LOC_114/Y 0.01fF
C51573 OR2X1_LOC_49/A OR2X1_LOC_80/A 0.10fF
C51574 AND2X1_LOC_477/A OR2X1_LOC_427/A 0.01fF
C51575 AND2X1_LOC_650/a_8_24# AND2X1_LOC_650/Y 0.01fF
C51576 OR2X1_LOC_186/Y OR2X1_LOC_353/a_8_216# 0.07fF
C51577 OR2X1_LOC_357/a_8_216# OR2X1_LOC_578/B 0.03fF
C51578 OR2X1_LOC_770/B OR2X1_LOC_80/A 0.06fF
C51579 OR2X1_LOC_524/Y GATE_811 0.03fF
C51580 OR2X1_LOC_160/A OR2X1_LOC_227/a_8_216# 0.01fF
C51581 AND2X1_LOC_711/Y AND2X1_LOC_620/a_8_24# 0.01fF
C51582 OR2X1_LOC_380/A OR2X1_LOC_64/Y 0.88fF
C51583 OR2X1_LOC_185/A OR2X1_LOC_335/B 0.39fF
C51584 OR2X1_LOC_426/A AND2X1_LOC_450/Y 0.03fF
C51585 OR2X1_LOC_306/Y OR2X1_LOC_46/A 0.63fF
C51586 AND2X1_LOC_7/B OR2X1_LOC_714/A 0.01fF
C51587 AND2X1_LOC_59/a_8_24# AND2X1_LOC_7/Y 0.00fF
C51588 AND2X1_LOC_683/a_36_24# AND2X1_LOC_3/Y 0.00fF
C51589 OR2X1_LOC_528/a_8_216# AND2X1_LOC_657/A 0.03fF
C51590 OR2X1_LOC_70/Y AND2X1_LOC_355/a_8_24# 0.01fF
C51591 VDD OR2X1_LOC_761/a_8_216# 0.21fF
C51592 AND2X1_LOC_22/Y OR2X1_LOC_769/a_8_216# 0.03fF
C51593 OR2X1_LOC_486/Y OR2X1_LOC_365/a_8_216# 0.02fF
C51594 OR2X1_LOC_71/Y AND2X1_LOC_573/A 0.14fF
C51595 VDD OR2X1_LOC_552/A 0.07fF
C51596 OR2X1_LOC_267/Y OR2X1_LOC_217/A 0.01fF
C51597 OR2X1_LOC_3/Y OR2X1_LOC_48/Y 0.04fF
C51598 OR2X1_LOC_6/B OR2X1_LOC_68/B 2.20fF
C51599 OR2X1_LOC_62/a_8_216# OR2X1_LOC_85/A 0.01fF
C51600 OR2X1_LOC_160/B OR2X1_LOC_228/Y 0.05fF
C51601 OR2X1_LOC_43/A OR2X1_LOC_19/B 0.07fF
C51602 OR2X1_LOC_481/Y AND2X1_LOC_345/a_8_24# 0.01fF
C51603 OR2X1_LOC_376/A OR2X1_LOC_409/B 0.01fF
C51604 OR2X1_LOC_596/A AND2X1_LOC_419/a_8_24# 0.01fF
C51605 OR2X1_LOC_52/Y OR2X1_LOC_7/A 0.11fF
C51606 AND2X1_LOC_22/Y OR2X1_LOC_723/B 0.01fF
C51607 AND2X1_LOC_285/Y AND2X1_LOC_562/Y 0.13fF
C51608 OR2X1_LOC_2/Y OR2X1_LOC_17/a_8_216# 0.41fF
C51609 OR2X1_LOC_214/a_36_216# OR2X1_LOC_750/A 0.02fF
C51610 OR2X1_LOC_485/A AND2X1_LOC_523/Y 0.05fF
C51611 OR2X1_LOC_160/B OR2X1_LOC_513/Y 0.00fF
C51612 AND2X1_LOC_66/a_8_24# OR2X1_LOC_44/Y 0.01fF
C51613 AND2X1_LOC_8/Y OR2X1_LOC_649/a_8_216# 0.00fF
C51614 OR2X1_LOC_62/B OR2X1_LOC_753/A 0.03fF
C51615 OR2X1_LOC_859/A OR2X1_LOC_269/B 0.03fF
C51616 AND2X1_LOC_476/Y OR2X1_LOC_164/a_8_216# 0.03fF
C51617 AND2X1_LOC_722/A OR2X1_LOC_419/Y 0.11fF
C51618 VDD OR2X1_LOC_578/B 0.39fF
C51619 VDD OR2X1_LOC_151/a_8_216# 0.21fF
C51620 AND2X1_LOC_70/Y OR2X1_LOC_568/a_36_216# 0.02fF
C51621 OR2X1_LOC_680/A AND2X1_LOC_675/A 0.56fF
C51622 OR2X1_LOC_80/a_8_216# OR2X1_LOC_6/A 0.09fF
C51623 AND2X1_LOC_12/Y OR2X1_LOC_276/a_8_216# 0.02fF
C51624 AND2X1_LOC_327/a_8_24# AND2X1_LOC_660/Y 0.20fF
C51625 OR2X1_LOC_218/Y OR2X1_LOC_222/A 0.04fF
C51626 OR2X1_LOC_380/A OR2X1_LOC_64/a_8_216# 0.01fF
C51627 AND2X1_LOC_73/a_8_24# OR2X1_LOC_68/B 0.01fF
C51628 AND2X1_LOC_335/a_8_24# AND2X1_LOC_222/Y 0.01fF
C51629 AND2X1_LOC_130/a_36_24# OR2X1_LOC_13/B 0.01fF
C51630 AND2X1_LOC_81/B OR2X1_LOC_506/B 0.01fF
C51631 OR2X1_LOC_771/B OR2X1_LOC_549/A 0.09fF
C51632 OR2X1_LOC_696/A AND2X1_LOC_721/Y 0.05fF
C51633 OR2X1_LOC_36/Y AND2X1_LOC_866/A 0.03fF
C51634 AND2X1_LOC_573/A D_INPUT_1 0.00fF
C51635 OR2X1_LOC_147/B OR2X1_LOC_551/B 0.07fF
C51636 OR2X1_LOC_441/Y AND2X1_LOC_222/Y 0.01fF
C51637 OR2X1_LOC_502/A OR2X1_LOC_358/A 0.01fF
C51638 OR2X1_LOC_335/A AND2X1_LOC_22/Y 0.00fF
C51639 OR2X1_LOC_307/a_36_216# AND2X1_LOC_47/Y 0.00fF
C51640 OR2X1_LOC_476/B OR2X1_LOC_476/a_8_216# 0.02fF
C51641 AND2X1_LOC_301/a_8_24# OR2X1_LOC_300/Y 0.01fF
C51642 OR2X1_LOC_666/A OR2X1_LOC_437/A 0.03fF
C51643 AND2X1_LOC_727/A AND2X1_LOC_856/B 0.00fF
C51644 AND2X1_LOC_393/a_36_24# OR2X1_LOC_84/A 0.01fF
C51645 AND2X1_LOC_831/Y OR2X1_LOC_74/A 0.01fF
C51646 OR2X1_LOC_277/a_8_216# AND2X1_LOC_633/Y 0.47fF
C51647 AND2X1_LOC_38/a_8_24# AND2X1_LOC_47/Y 0.02fF
C51648 OR2X1_LOC_3/Y AND2X1_LOC_656/Y 0.09fF
C51649 AND2X1_LOC_91/B OR2X1_LOC_97/A 0.08fF
C51650 OR2X1_LOC_503/Y OR2X1_LOC_7/A 0.01fF
C51651 AND2X1_LOC_727/A AND2X1_LOC_863/A 0.17fF
C51652 OR2X1_LOC_479/Y AND2X1_LOC_47/Y 0.10fF
C51653 OR2X1_LOC_362/B OR2X1_LOC_675/Y 0.32fF
C51654 AND2X1_LOC_43/B OR2X1_LOC_196/a_8_216# 0.05fF
C51655 OR2X1_LOC_161/A OR2X1_LOC_318/B 0.02fF
C51656 AND2X1_LOC_486/Y AND2X1_LOC_793/B 0.17fF
C51657 OR2X1_LOC_32/B OR2X1_LOC_598/A 0.46fF
C51658 AND2X1_LOC_727/Y AND2X1_LOC_727/a_8_24# 0.01fF
C51659 AND2X1_LOC_22/Y OR2X1_LOC_720/Y 0.08fF
C51660 OR2X1_LOC_270/Y AND2X1_LOC_252/a_8_24# 0.01fF
C51661 OR2X1_LOC_502/A OR2X1_LOC_460/A 0.01fF
C51662 OR2X1_LOC_519/Y AND2X1_LOC_222/Y 0.00fF
C51663 OR2X1_LOC_617/Y OR2X1_LOC_95/Y 0.02fF
C51664 AND2X1_LOC_552/a_8_24# OR2X1_LOC_373/Y 0.00fF
C51665 AND2X1_LOC_530/a_8_24# OR2X1_LOC_415/Y 0.01fF
C51666 AND2X1_LOC_56/B OR2X1_LOC_493/Y 0.01fF
C51667 OR2X1_LOC_70/Y OR2X1_LOC_72/a_36_216# 0.03fF
C51668 OR2X1_LOC_656/B AND2X1_LOC_31/Y 0.02fF
C51669 OR2X1_LOC_161/A OR2X1_LOC_854/A 0.03fF
C51670 AND2X1_LOC_462/Y OR2X1_LOC_27/Y 0.30fF
C51671 AND2X1_LOC_539/a_8_24# OR2X1_LOC_22/Y 0.01fF
C51672 OR2X1_LOC_627/a_36_216# AND2X1_LOC_624/B 0.00fF
C51673 AND2X1_LOC_159/a_8_24# AND2X1_LOC_72/B 0.01fF
C51674 OR2X1_LOC_323/A OR2X1_LOC_322/Y 0.02fF
C51675 AND2X1_LOC_12/Y OR2X1_LOC_513/a_8_216# 0.01fF
C51676 AND2X1_LOC_857/Y OR2X1_LOC_13/B 0.03fF
C51677 OR2X1_LOC_836/Y OR2X1_LOC_839/a_8_216# 0.39fF
C51678 OR2X1_LOC_91/A AND2X1_LOC_789/Y 0.02fF
C51679 AND2X1_LOC_716/Y OR2X1_LOC_437/A 0.02fF
C51680 AND2X1_LOC_464/Y OR2X1_LOC_95/Y 0.01fF
C51681 AND2X1_LOC_794/B AND2X1_LOC_794/a_8_24# 0.02fF
C51682 OR2X1_LOC_89/A OR2X1_LOC_815/Y 0.01fF
C51683 OR2X1_LOC_791/B OR2X1_LOC_348/B 0.03fF
C51684 AND2X1_LOC_810/B OR2X1_LOC_428/A 0.14fF
C51685 OR2X1_LOC_586/Y OR2X1_LOC_385/a_8_216# 0.03fF
C51686 OR2X1_LOC_579/B OR2X1_LOC_68/B 0.07fF
C51687 OR2X1_LOC_97/A OR2X1_LOC_364/a_8_216# 0.01fF
C51688 OR2X1_LOC_479/Y OR2X1_LOC_795/a_36_216# 0.00fF
C51689 AND2X1_LOC_534/a_8_24# OR2X1_LOC_161/B 0.02fF
C51690 AND2X1_LOC_340/Y OR2X1_LOC_595/A 0.00fF
C51691 AND2X1_LOC_363/a_8_24# OR2X1_LOC_428/A 0.01fF
C51692 VDD OR2X1_LOC_366/A -0.00fF
C51693 AND2X1_LOC_181/Y OR2X1_LOC_428/A 0.03fF
C51694 OR2X1_LOC_111/a_36_216# AND2X1_LOC_326/B 0.00fF
C51695 AND2X1_LOC_40/Y OR2X1_LOC_535/a_8_216# 0.01fF
C51696 OR2X1_LOC_52/B OR2X1_LOC_745/Y 0.01fF
C51697 OR2X1_LOC_833/B AND2X1_LOC_268/a_36_24# 0.00fF
C51698 OR2X1_LOC_506/A OR2X1_LOC_728/A 0.03fF
C51699 OR2X1_LOC_167/Y AND2X1_LOC_169/a_8_24# 0.00fF
C51700 OR2X1_LOC_219/B OR2X1_LOC_228/Y 0.02fF
C51701 OR2X1_LOC_675/A OR2X1_LOC_241/B 0.03fF
C51702 OR2X1_LOC_736/Y OR2X1_LOC_741/a_8_216# 0.03fF
C51703 OR2X1_LOC_7/A OR2X1_LOC_754/Y 0.05fF
C51704 OR2X1_LOC_51/Y AND2X1_LOC_241/a_8_24# 0.01fF
C51705 AND2X1_LOC_59/Y OR2X1_LOC_366/Y 0.04fF
C51706 OR2X1_LOC_156/B OR2X1_LOC_156/A 0.15fF
C51707 VDD GATE_579 0.21fF
C51708 AND2X1_LOC_729/B OR2X1_LOC_311/a_36_216# 0.00fF
C51709 OR2X1_LOC_40/a_8_216# D_INPUT_6 0.00fF
C51710 AND2X1_LOC_110/Y OR2X1_LOC_161/B 0.48fF
C51711 OR2X1_LOC_614/Y AND2X1_LOC_754/a_8_24# 0.05fF
C51712 OR2X1_LOC_369/Y AND2X1_LOC_370/a_8_24# 0.09fF
C51713 AND2X1_LOC_612/B OR2X1_LOC_80/A 0.15fF
C51714 AND2X1_LOC_64/Y OR2X1_LOC_78/Y 0.03fF
C51715 AND2X1_LOC_766/a_8_24# OR2X1_LOC_78/B 0.01fF
C51716 OR2X1_LOC_97/A OR2X1_LOC_645/a_8_216# 0.01fF
C51717 AND2X1_LOC_51/Y OR2X1_LOC_318/B 0.03fF
C51718 OR2X1_LOC_421/A AND2X1_LOC_828/a_8_24# 0.01fF
C51719 OR2X1_LOC_856/A OR2X1_LOC_598/Y 0.00fF
C51720 OR2X1_LOC_480/a_36_216# OR2X1_LOC_467/A 0.00fF
C51721 AND2X1_LOC_339/Y OR2X1_LOC_51/Y 0.03fF
C51722 AND2X1_LOC_85/a_8_24# OR2X1_LOC_80/A 0.02fF
C51723 OR2X1_LOC_805/A OR2X1_LOC_332/a_36_216# 0.02fF
C51724 GATE_366 OR2X1_LOC_437/A 0.07fF
C51725 OR2X1_LOC_131/Y AND2X1_LOC_657/A 0.28fF
C51726 OR2X1_LOC_329/B OR2X1_LOC_312/a_8_216# 0.01fF
C51727 AND2X1_LOC_658/A AND2X1_LOC_213/B 0.03fF
C51728 AND2X1_LOC_432/a_36_24# OR2X1_LOC_648/A 0.01fF
C51729 OR2X1_LOC_769/B AND2X1_LOC_22/Y 0.17fF
C51730 OR2X1_LOC_830/a_36_216# OR2X1_LOC_294/Y 0.00fF
C51731 OR2X1_LOC_114/B OR2X1_LOC_346/A 0.03fF
C51732 OR2X1_LOC_846/B OR2X1_LOC_557/a_8_216# 0.12fF
C51733 AND2X1_LOC_477/Y AND2X1_LOC_478/a_8_24# 0.03fF
C51734 OR2X1_LOC_622/a_36_216# OR2X1_LOC_80/A 0.00fF
C51735 OR2X1_LOC_696/A OR2X1_LOC_586/Y 0.52fF
C51736 OR2X1_LOC_133/a_8_216# OR2X1_LOC_8/Y 0.01fF
C51737 AND2X1_LOC_60/a_36_24# OR2X1_LOC_648/A 0.01fF
C51738 AND2X1_LOC_56/B OR2X1_LOC_532/a_8_216# 0.04fF
C51739 OR2X1_LOC_174/A AND2X1_LOC_7/B 0.01fF
C51740 AND2X1_LOC_392/A OR2X1_LOC_158/A 0.17fF
C51741 OR2X1_LOC_375/A OR2X1_LOC_593/B 0.01fF
C51742 AND2X1_LOC_479/Y OR2X1_LOC_47/Y 0.01fF
C51743 AND2X1_LOC_48/A OR2X1_LOC_358/A 0.07fF
C51744 OR2X1_LOC_312/Y OR2X1_LOC_437/A 0.10fF
C51745 OR2X1_LOC_456/Y AND2X1_LOC_36/Y 0.09fF
C51746 OR2X1_LOC_12/Y OR2X1_LOC_59/Y 0.14fF
C51747 OR2X1_LOC_851/B OR2X1_LOC_851/a_8_216# 0.05fF
C51748 AND2X1_LOC_70/Y AND2X1_LOC_65/A 0.25fF
C51749 OR2X1_LOC_6/B AND2X1_LOC_626/a_36_24# 0.00fF
C51750 INPUT_0 AND2X1_LOC_774/A 0.01fF
C51751 OR2X1_LOC_545/B OR2X1_LOC_551/B 0.07fF
C51752 AND2X1_LOC_471/Y OR2X1_LOC_373/Y 0.03fF
C51753 AND2X1_LOC_64/Y OR2X1_LOC_724/a_8_216# 0.02fF
C51754 VDD OR2X1_LOC_583/a_8_216# 0.00fF
C51755 AND2X1_LOC_562/B OR2X1_LOC_816/A 0.03fF
C51756 AND2X1_LOC_82/Y OR2X1_LOC_78/Y 0.37fF
C51757 OR2X1_LOC_691/Y OR2X1_LOC_637/A 0.01fF
C51758 OR2X1_LOC_160/A OR2X1_LOC_140/B 0.04fF
C51759 AND2X1_LOC_482/a_8_24# AND2X1_LOC_7/B 0.04fF
C51760 AND2X1_LOC_366/A OR2X1_LOC_158/A 0.02fF
C51761 OR2X1_LOC_68/Y OR2X1_LOC_68/B 0.01fF
C51762 OR2X1_LOC_506/a_8_216# OR2X1_LOC_375/A 0.01fF
C51763 AND2X1_LOC_535/Y AND2X1_LOC_434/Y 0.00fF
C51764 AND2X1_LOC_544/Y AND2X1_LOC_624/A 0.03fF
C51765 AND2X1_LOC_721/Y AND2X1_LOC_717/a_8_24# 0.05fF
C51766 OR2X1_LOC_641/Y OR2X1_LOC_640/Y 0.12fF
C51767 AND2X1_LOC_572/A AND2X1_LOC_772/Y 0.01fF
C51768 OR2X1_LOC_139/A AND2X1_LOC_95/Y 0.06fF
C51769 OR2X1_LOC_68/a_36_216# OR2X1_LOC_776/A 0.01fF
C51770 AND2X1_LOC_16/a_8_24# AND2X1_LOC_44/Y -0.06fF
C51771 OR2X1_LOC_389/A AND2X1_LOC_92/Y 0.06fF
C51772 AND2X1_LOC_500/Y AND2X1_LOC_501/a_8_24# 0.01fF
C51773 OR2X1_LOC_840/A OR2X1_LOC_596/A 0.03fF
C51774 OR2X1_LOC_528/Y AND2X1_LOC_508/A 0.06fF
C51775 OR2X1_LOC_600/A AND2X1_LOC_474/A 0.03fF
C51776 AND2X1_LOC_47/Y OR2X1_LOC_68/B 0.28fF
C51777 OR2X1_LOC_616/Y GATE_579 0.11fF
C51778 AND2X1_LOC_190/a_8_24# OR2X1_LOC_744/A -0.02fF
C51779 AND2X1_LOC_331/a_8_24# OR2X1_LOC_151/A 0.03fF
C51780 OR2X1_LOC_377/A AND2X1_LOC_44/Y 0.11fF
C51781 OR2X1_LOC_160/A OR2X1_LOC_355/A 0.02fF
C51782 OR2X1_LOC_648/A OR2X1_LOC_78/A 0.07fF
C51783 OR2X1_LOC_426/B OR2X1_LOC_91/A 0.20fF
C51784 AND2X1_LOC_721/Y AND2X1_LOC_458/Y 0.01fF
C51785 OR2X1_LOC_185/A OR2X1_LOC_633/A 0.10fF
C51786 OR2X1_LOC_604/A AND2X1_LOC_722/A 0.54fF
C51787 OR2X1_LOC_864/A OR2X1_LOC_338/B 0.10fF
C51788 AND2X1_LOC_354/a_8_24# OR2X1_LOC_428/A 0.04fF
C51789 AND2X1_LOC_56/B AND2X1_LOC_829/a_36_24# 0.00fF
C51790 VDD OR2X1_LOC_798/Y 0.00fF
C51791 AND2X1_LOC_675/Y AND2X1_LOC_548/Y 0.35fF
C51792 AND2X1_LOC_189/a_36_24# OR2X1_LOC_741/Y 0.01fF
C51793 VDD AND2X1_LOC_52/a_8_24# -0.00fF
C51794 OR2X1_LOC_632/a_8_216# OR2X1_LOC_632/Y 0.00fF
C51795 OR2X1_LOC_664/Y OR2X1_LOC_161/B 0.35fF
C51796 OR2X1_LOC_812/A OR2X1_LOC_812/a_8_216# 0.39fF
C51797 OR2X1_LOC_45/B OR2X1_LOC_305/a_8_216# 0.01fF
C51798 AND2X1_LOC_592/Y OR2X1_LOC_48/B 0.05fF
C51799 OR2X1_LOC_175/Y OR2X1_LOC_778/Y 0.10fF
C51800 OR2X1_LOC_804/a_36_216# AND2X1_LOC_92/Y 0.03fF
C51801 OR2X1_LOC_203/Y AND2X1_LOC_44/Y 0.11fF
C51802 AND2X1_LOC_716/Y AND2X1_LOC_715/A 0.07fF
C51803 VDD OR2X1_LOC_814/a_8_216# 0.21fF
C51804 OR2X1_LOC_49/A OR2X1_LOC_6/A 0.62fF
C51805 AND2X1_LOC_658/A OR2X1_LOC_144/Y 0.03fF
C51806 OR2X1_LOC_3/Y AND2X1_LOC_772/Y 0.07fF
C51807 OR2X1_LOC_238/Y AND2X1_LOC_242/B 0.01fF
C51808 OR2X1_LOC_51/Y OR2X1_LOC_92/Y 0.06fF
C51809 OR2X1_LOC_528/Y OR2X1_LOC_18/Y 0.16fF
C51810 OR2X1_LOC_620/Y AND2X1_LOC_299/a_36_24# 0.00fF
C51811 OR2X1_LOC_95/Y OR2X1_LOC_536/a_8_216# 0.01fF
C51812 OR2X1_LOC_482/Y AND2X1_LOC_474/a_8_24# 0.06fF
C51813 INPUT_5 OR2X1_LOC_25/Y 4.36fF
C51814 OR2X1_LOC_45/B AND2X1_LOC_458/a_8_24# 0.01fF
C51815 OR2X1_LOC_124/A OR2X1_LOC_264/Y 0.07fF
C51816 AND2X1_LOC_305/a_36_24# OR2X1_LOC_307/A 0.00fF
C51817 AND2X1_LOC_715/A AND2X1_LOC_654/Y 0.07fF
C51818 OR2X1_LOC_585/A OR2X1_LOC_428/A 0.10fF
C51819 OR2X1_LOC_753/A OR2X1_LOC_15/a_36_216# 0.00fF
C51820 AND2X1_LOC_753/B OR2X1_LOC_638/B 0.07fF
C51821 AND2X1_LOC_59/Y OR2X1_LOC_786/A 0.16fF
C51822 OR2X1_LOC_820/B OR2X1_LOC_12/Y 0.04fF
C51823 AND2X1_LOC_178/a_8_24# OR2X1_LOC_190/Y 0.09fF
C51824 OR2X1_LOC_114/B OR2X1_LOC_161/A 0.06fF
C51825 AND2X1_LOC_422/a_8_24# AND2X1_LOC_92/Y 0.04fF
C51826 OR2X1_LOC_600/A AND2X1_LOC_593/Y 3.04fF
C51827 OR2X1_LOC_229/Y AND2X1_LOC_231/a_8_24# 0.23fF
C51828 OR2X1_LOC_121/Y OR2X1_LOC_116/a_36_216# 0.01fF
C51829 AND2X1_LOC_124/a_8_24# AND2X1_LOC_243/Y 0.04fF
C51830 AND2X1_LOC_789/a_8_24# OR2X1_LOC_820/A 0.04fF
C51831 AND2X1_LOC_41/a_8_24# OR2X1_LOC_375/A 0.01fF
C51832 OR2X1_LOC_604/A AND2X1_LOC_454/Y 0.00fF
C51833 OR2X1_LOC_331/a_8_216# OR2X1_LOC_331/Y 0.03fF
C51834 AND2X1_LOC_658/A OR2X1_LOC_531/a_36_216# 0.02fF
C51835 OR2X1_LOC_778/Y OR2X1_LOC_713/A 0.10fF
C51836 OR2X1_LOC_739/A OR2X1_LOC_66/A 0.03fF
C51837 OR2X1_LOC_13/Y OR2X1_LOC_44/Y 0.03fF
C51838 AND2X1_LOC_808/a_8_24# AND2X1_LOC_469/B 0.01fF
C51839 OR2X1_LOC_756/B OR2X1_LOC_400/a_8_216# 0.02fF
C51840 OR2X1_LOC_68/B OR2X1_LOC_598/A 0.08fF
C51841 OR2X1_LOC_841/a_8_216# OR2X1_LOC_776/a_8_216# 0.47fF
C51842 OR2X1_LOC_347/B OR2X1_LOC_347/Y 0.05fF
C51843 OR2X1_LOC_426/B AND2X1_LOC_573/A 0.11fF
C51844 OR2X1_LOC_217/a_8_216# OR2X1_LOC_549/A 0.03fF
C51845 D_INPUT_1 OR2X1_LOC_558/a_8_216# 0.02fF
C51846 OR2X1_LOC_744/A AND2X1_LOC_99/A 0.03fF
C51847 VDD OR2X1_LOC_314/Y 0.08fF
C51848 OR2X1_LOC_188/Y OR2X1_LOC_675/A 0.02fF
C51849 AND2X1_LOC_81/B AND2X1_LOC_18/Y 0.03fF
C51850 AND2X1_LOC_817/B VDD 0.37fF
C51851 OR2X1_LOC_40/Y OR2X1_LOC_36/Y 0.17fF
C51852 OR2X1_LOC_40/Y OR2X1_LOC_91/a_8_216# 0.02fF
C51853 AND2X1_LOC_18/Y OR2X1_LOC_358/B 0.05fF
C51854 OR2X1_LOC_600/A OR2X1_LOC_85/A 0.66fF
C51855 OR2X1_LOC_267/A OR2X1_LOC_641/A 0.04fF
C51856 OR2X1_LOC_599/A OR2X1_LOC_604/A 0.03fF
C51857 AND2X1_LOC_764/a_8_24# OR2X1_LOC_828/B 0.01fF
C51858 AND2X1_LOC_860/a_8_24# AND2X1_LOC_850/Y 0.02fF
C51859 AND2X1_LOC_512/Y OR2X1_LOC_48/B 0.46fF
C51860 OR2X1_LOC_648/A OR2X1_LOC_602/A 0.05fF
C51861 OR2X1_LOC_756/B OR2X1_LOC_847/A 0.00fF
C51862 OR2X1_LOC_70/Y OR2X1_LOC_12/Y 0.54fF
C51863 AND2X1_LOC_860/A AND2X1_LOC_806/A 0.02fF
C51864 OR2X1_LOC_151/A AND2X1_LOC_329/a_36_24# 0.00fF
C51865 OR2X1_LOC_538/A OR2X1_LOC_161/A 0.07fF
C51866 OR2X1_LOC_438/a_8_216# AND2X1_LOC_476/Y 0.04fF
C51867 OR2X1_LOC_329/B AND2X1_LOC_114/a_8_24# 0.04fF
C51868 OR2X1_LOC_6/B AND2X1_LOC_673/a_8_24# 0.03fF
C51869 AND2X1_LOC_725/a_8_24# OR2X1_LOC_52/B 0.02fF
C51870 OR2X1_LOC_6/B AND2X1_LOC_81/a_36_24# 0.01fF
C51871 OR2X1_LOC_269/B OR2X1_LOC_66/A 0.24fF
C51872 OR2X1_LOC_109/Y OR2X1_LOC_164/Y 0.78fF
C51873 OR2X1_LOC_64/Y AND2X1_LOC_774/A 0.00fF
C51874 AND2X1_LOC_3/Y OR2X1_LOC_631/A 0.03fF
C51875 OR2X1_LOC_843/a_36_216# OR2X1_LOC_362/A 0.00fF
C51876 OR2X1_LOC_850/B AND2X1_LOC_95/Y 0.01fF
C51877 OR2X1_LOC_53/Y OR2X1_LOC_7/Y 0.02fF
C51878 AND2X1_LOC_307/a_36_24# AND2X1_LOC_774/A 0.03fF
C51879 AND2X1_LOC_318/Y AND2X1_LOC_269/a_36_24# 0.00fF
C51880 OR2X1_LOC_121/Y AND2X1_LOC_51/Y 0.07fF
C51881 OR2X1_LOC_160/B OR2X1_LOC_287/B 0.04fF
C51882 OR2X1_LOC_45/B AND2X1_LOC_537/Y 0.07fF
C51883 OR2X1_LOC_589/A OR2X1_LOC_275/A 0.02fF
C51884 OR2X1_LOC_683/Y OR2X1_LOC_16/A 0.08fF
C51885 OR2X1_LOC_6/B OR2X1_LOC_74/A 0.07fF
C51886 OR2X1_LOC_759/A OR2X1_LOC_89/A 0.04fF
C51887 VDD OR2X1_LOC_654/A 0.22fF
C51888 AND2X1_LOC_127/a_8_24# OR2X1_LOC_342/A 0.25fF
C51889 AND2X1_LOC_474/Y AND2X1_LOC_657/Y 0.14fF
C51890 OR2X1_LOC_814/A OR2X1_LOC_576/A 0.02fF
C51891 OR2X1_LOC_648/A OR2X1_LOC_155/A 0.07fF
C51892 OR2X1_LOC_698/a_8_216# OR2X1_LOC_36/Y 0.01fF
C51893 OR2X1_LOC_744/A AND2X1_LOC_637/Y 0.02fF
C51894 OR2X1_LOC_351/B AND2X1_LOC_51/Y 0.09fF
C51895 OR2X1_LOC_792/Y OR2X1_LOC_806/a_8_216# 0.02fF
C51896 VDD OR2X1_LOC_131/Y 0.25fF
C51897 AND2X1_LOC_538/a_8_24# OR2X1_LOC_12/Y 0.09fF
C51898 AND2X1_LOC_191/B OR2X1_LOC_485/A 0.07fF
C51899 OR2X1_LOC_3/Y AND2X1_LOC_160/Y 0.01fF
C51900 AND2X1_LOC_81/B OR2X1_LOC_473/a_8_216# 0.14fF
C51901 D_INPUT_5 AND2X1_LOC_25/Y 0.01fF
C51902 OR2X1_LOC_808/B OR2X1_LOC_468/Y 0.05fF
C51903 OR2X1_LOC_485/A AND2X1_LOC_469/B 0.04fF
C51904 OR2X1_LOC_516/A OR2X1_LOC_48/B 0.03fF
C51905 AND2X1_LOC_3/Y OR2X1_LOC_632/Y 0.01fF
C51906 AND2X1_LOC_593/Y OR2X1_LOC_619/Y 0.03fF
C51907 OR2X1_LOC_700/Y OR2X1_LOC_701/Y 0.94fF
C51908 OR2X1_LOC_160/B OR2X1_LOC_76/A 0.13fF
C51909 AND2X1_LOC_550/A AND2X1_LOC_624/A 0.03fF
C51910 OR2X1_LOC_743/A OR2X1_LOC_91/A 0.07fF
C51911 OR2X1_LOC_246/A OR2X1_LOC_131/a_8_216# 0.18fF
C51912 OR2X1_LOC_272/Y OR2X1_LOC_59/Y 0.16fF
C51913 AND2X1_LOC_12/Y OR2X1_LOC_161/A 0.16fF
C51914 AND2X1_LOC_59/Y OR2X1_LOC_624/A 0.01fF
C51915 AND2X1_LOC_367/A OR2X1_LOC_529/Y 0.59fF
C51916 AND2X1_LOC_486/Y AND2X1_LOC_859/Y 0.10fF
C51917 AND2X1_LOC_22/a_8_24# AND2X1_LOC_25/Y 0.11fF
C51918 AND2X1_LOC_733/Y OR2X1_LOC_485/A 0.03fF
C51919 AND2X1_LOC_852/a_36_24# AND2X1_LOC_852/B 0.01fF
C51920 OR2X1_LOC_698/Y OR2X1_LOC_89/A 0.03fF
C51921 OR2X1_LOC_196/B AND2X1_LOC_18/Y 0.09fF
C51922 OR2X1_LOC_520/Y OR2X1_LOC_185/A 0.49fF
C51923 OR2X1_LOC_519/a_8_216# OR2X1_LOC_6/A 0.01fF
C51924 AND2X1_LOC_476/A AND2X1_LOC_786/Y 0.02fF
C51925 AND2X1_LOC_113/Y AND2X1_LOC_114/a_8_24# 0.11fF
C51926 AND2X1_LOC_56/B OR2X1_LOC_194/B 0.04fF
C51927 OR2X1_LOC_85/A OR2X1_LOC_619/Y 0.10fF
C51928 OR2X1_LOC_822/Y OR2X1_LOC_54/Y 0.01fF
C51929 OR2X1_LOC_538/a_8_216# OR2X1_LOC_702/A 0.01fF
C51930 OR2X1_LOC_441/Y OR2X1_LOC_74/A 14.70fF
C51931 OR2X1_LOC_36/Y AND2X1_LOC_644/Y 0.04fF
C51932 AND2X1_LOC_348/A AND2X1_LOC_294/a_36_24# 0.00fF
C51933 OR2X1_LOC_700/Y OR2X1_LOC_44/Y 0.29fF
C51934 OR2X1_LOC_213/A OR2X1_LOC_209/a_8_216# 0.01fF
C51935 AND2X1_LOC_215/Y AND2X1_LOC_634/Y 0.37fF
C51936 D_INPUT_3 OR2X1_LOC_381/a_8_216# 0.02fF
C51937 OR2X1_LOC_538/A AND2X1_LOC_51/Y 0.03fF
C51938 OR2X1_LOC_13/B OR2X1_LOC_437/A 0.49fF
C51939 OR2X1_LOC_656/B OR2X1_LOC_864/A 0.07fF
C51940 OR2X1_LOC_36/Y OR2X1_LOC_424/a_8_216# 0.01fF
C51941 OR2X1_LOC_476/B AND2X1_LOC_20/a_8_24# 0.02fF
C51942 AND2X1_LOC_570/Y OR2X1_LOC_22/Y 0.02fF
C51943 OR2X1_LOC_270/a_36_216# OR2X1_LOC_375/A 0.02fF
C51944 AND2X1_LOC_70/Y AND2X1_LOC_23/a_8_24# 0.01fF
C51945 OR2X1_LOC_649/a_8_216# AND2X1_LOC_92/Y 0.01fF
C51946 OR2X1_LOC_223/A OR2X1_LOC_486/Y 0.03fF
C51947 AND2X1_LOC_94/Y OR2X1_LOC_46/A 0.10fF
C51948 OR2X1_LOC_88/A OR2X1_LOC_85/A 0.05fF
C51949 OR2X1_LOC_91/A OR2X1_LOC_125/Y 0.06fF
C51950 OR2X1_LOC_641/Y OR2X1_LOC_655/B 0.12fF
C51951 OR2X1_LOC_278/Y AND2X1_LOC_240/Y 0.02fF
C51952 OR2X1_LOC_476/B OR2X1_LOC_634/A 0.10fF
C51953 OR2X1_LOC_472/a_8_216# OR2X1_LOC_640/A 0.40fF
C51954 OR2X1_LOC_91/A OR2X1_LOC_246/A 0.14fF
C51955 D_INPUT_5 AND2X1_LOC_51/Y 0.03fF
C51956 AND2X1_LOC_1/a_8_24# AND2X1_LOC_17/a_8_24# 0.23fF
C51957 OR2X1_LOC_69/A OR2X1_LOC_52/B 0.87fF
C51958 OR2X1_LOC_604/A AND2X1_LOC_866/A 0.10fF
C51959 OR2X1_LOC_666/A AND2X1_LOC_845/Y 0.07fF
C51960 OR2X1_LOC_401/Y OR2X1_LOC_402/Y 0.03fF
C51961 AND2X1_LOC_190/a_8_24# OR2X1_LOC_31/Y 0.02fF
C51962 AND2X1_LOC_391/Y OR2X1_LOC_225/a_8_216# -0.03fF
C51963 OR2X1_LOC_604/A OR2X1_LOC_426/a_36_216# 0.00fF
C51964 AND2X1_LOC_287/Y AND2X1_LOC_806/A 0.16fF
C51965 OR2X1_LOC_18/Y OR2X1_LOC_279/a_8_216# 0.02fF
C51966 OR2X1_LOC_91/A OR2X1_LOC_225/a_8_216# 0.01fF
C51967 OR2X1_LOC_479/Y OR2X1_LOC_506/A 0.02fF
C51968 AND2X1_LOC_41/A OR2X1_LOC_814/A 0.10fF
C51969 GATE_366 OR2X1_LOC_753/A 0.02fF
C51970 AND2X1_LOC_654/a_8_24# OR2X1_LOC_6/A 0.01fF
C51971 OR2X1_LOC_47/Y AND2X1_LOC_243/Y 0.04fF
C51972 OR2X1_LOC_474/a_36_216# OR2X1_LOC_474/Y 0.01fF
C51973 AND2X1_LOC_22/a_8_24# AND2X1_LOC_51/Y 0.01fF
C51974 OR2X1_LOC_804/B OR2X1_LOC_161/A 0.47fF
C51975 OR2X1_LOC_528/Y AND2X1_LOC_620/Y 0.04fF
C51976 AND2X1_LOC_702/Y OR2X1_LOC_52/B 0.03fF
C51977 OR2X1_LOC_87/A AND2X1_LOC_118/a_8_24# 0.01fF
C51978 OR2X1_LOC_112/B AND2X1_LOC_18/Y 0.02fF
C51979 AND2X1_LOC_139/B OR2X1_LOC_74/A 0.07fF
C51980 AND2X1_LOC_259/Y OR2X1_LOC_6/A 0.01fF
C51981 AND2X1_LOC_568/B OR2X1_LOC_47/Y 0.07fF
C51982 OR2X1_LOC_36/Y OR2X1_LOC_7/A 0.63fF
C51983 OR2X1_LOC_705/B OR2X1_LOC_486/Y 0.01fF
C51984 OR2X1_LOC_70/A OR2X1_LOC_12/Y 0.02fF
C51985 OR2X1_LOC_409/B AND2X1_LOC_637/a_36_24# -0.00fF
C51986 AND2X1_LOC_476/A AND2X1_LOC_218/Y 0.01fF
C51987 OR2X1_LOC_185/A OR2X1_LOC_479/a_8_216# 0.01fF
C51988 AND2X1_LOC_122/a_8_24# OR2X1_LOC_510/Y 0.02fF
C51989 OR2X1_LOC_666/Y AND2X1_LOC_859/Y 0.02fF
C51990 OR2X1_LOC_34/A OR2X1_LOC_68/B 0.00fF
C51991 OR2X1_LOC_462/B AND2X1_LOC_42/B 0.09fF
C51992 OR2X1_LOC_137/Y OR2X1_LOC_139/a_8_216# 0.18fF
C51993 AND2X1_LOC_12/Y AND2X1_LOC_51/Y 2.24fF
C51994 AND2X1_LOC_736/a_8_24# OR2X1_LOC_95/Y 0.03fF
C51995 OR2X1_LOC_502/A OR2X1_LOC_818/a_8_216# 0.01fF
C51996 AND2X1_LOC_580/A AND2X1_LOC_578/A 0.00fF
C51997 OR2X1_LOC_154/A OR2X1_LOC_201/Y 0.05fF
C51998 AND2X1_LOC_465/Y OR2X1_LOC_427/A 0.10fF
C51999 AND2X1_LOC_654/a_36_24# OR2X1_LOC_52/B 0.00fF
C52000 OR2X1_LOC_808/a_36_216# OR2X1_LOC_814/A 0.01fF
C52001 OR2X1_LOC_235/Y OR2X1_LOC_74/A 0.01fF
C52002 AND2X1_LOC_1/Y AND2X1_LOC_47/a_36_24# 0.00fF
C52003 OR2X1_LOC_320/Y OR2X1_LOC_36/Y 0.01fF
C52004 OR2X1_LOC_40/Y OR2X1_LOC_419/Y 0.08fF
C52005 AND2X1_LOC_170/a_8_24# AND2X1_LOC_514/Y 0.02fF
C52006 OR2X1_LOC_8/Y AND2X1_LOC_837/a_36_24# 0.00fF
C52007 OR2X1_LOC_413/a_8_216# OR2X1_LOC_46/A 0.01fF
C52008 OR2X1_LOC_794/a_36_216# OR2X1_LOC_269/B 0.02fF
C52009 AND2X1_LOC_470/a_8_24# OR2X1_LOC_619/Y 0.01fF
C52010 OR2X1_LOC_76/A OR2X1_LOC_553/A 0.05fF
C52011 OR2X1_LOC_744/A AND2X1_LOC_810/a_8_24# 0.01fF
C52012 OR2X1_LOC_857/B AND2X1_LOC_31/Y 0.02fF
C52013 D_INPUT_0 AND2X1_LOC_649/B 0.07fF
C52014 OR2X1_LOC_246/A AND2X1_LOC_573/A 0.02fF
C52015 OR2X1_LOC_40/Y AND2X1_LOC_202/a_36_24# 0.00fF
C52016 AND2X1_LOC_456/Y OR2X1_LOC_529/Y 0.02fF
C52017 OR2X1_LOC_43/A OR2X1_LOC_275/A 0.06fF
C52018 OR2X1_LOC_154/A OR2X1_LOC_844/Y 0.01fF
C52019 AND2X1_LOC_326/A AND2X1_LOC_354/B 0.06fF
C52020 VDD OR2X1_LOC_192/B 0.21fF
C52021 VDD OR2X1_LOC_76/a_8_216# 0.21fF
C52022 OR2X1_LOC_235/B AND2X1_LOC_8/a_8_24# 0.01fF
C52023 OR2X1_LOC_756/B AND2X1_LOC_250/a_36_24# 0.00fF
C52024 AND2X1_LOC_136/a_8_24# OR2X1_LOC_155/A 0.03fF
C52025 OR2X1_LOC_748/A AND2X1_LOC_663/B 0.03fF
C52026 OR2X1_LOC_97/A OR2X1_LOC_303/B 0.18fF
C52027 OR2X1_LOC_646/B OR2X1_LOC_68/B 0.32fF
C52028 OR2X1_LOC_46/A OR2X1_LOC_265/Y 0.03fF
C52029 AND2X1_LOC_92/Y OR2X1_LOC_493/Y 0.07fF
C52030 OR2X1_LOC_641/A OR2X1_LOC_560/A 0.03fF
C52031 AND2X1_LOC_736/Y OR2X1_LOC_47/Y 0.03fF
C52032 VDD AND2X1_LOC_657/A 0.05fF
C52033 AND2X1_LOC_79/Y AND2X1_LOC_51/Y 0.01fF
C52034 OR2X1_LOC_613/Y AND2X1_LOC_632/A 0.04fF
C52035 OR2X1_LOC_344/A OR2X1_LOC_367/a_36_216# 0.00fF
C52036 AND2X1_LOC_150/a_8_24# OR2X1_LOC_140/Y 0.01fF
C52037 OR2X1_LOC_436/Y OR2X1_LOC_799/a_8_216# 0.01fF
C52038 OR2X1_LOC_468/a_8_216# OR2X1_LOC_539/Y 0.01fF
C52039 AND2X1_LOC_227/Y OR2X1_LOC_265/Y 0.17fF
C52040 AND2X1_LOC_859/a_8_24# AND2X1_LOC_859/B 0.12fF
C52041 AND2X1_LOC_43/B AND2X1_LOC_827/a_8_24# 0.01fF
C52042 OR2X1_LOC_154/A OR2X1_LOC_201/a_8_216# 0.01fF
C52043 OR2X1_LOC_669/a_8_216# OR2X1_LOC_417/A 0.01fF
C52044 OR2X1_LOC_532/B OR2X1_LOC_720/a_8_216# 0.01fF
C52045 OR2X1_LOC_70/A OR2X1_LOC_763/a_36_216# 0.00fF
C52046 OR2X1_LOC_41/a_36_216# OR2X1_LOC_48/B 0.02fF
C52047 OR2X1_LOC_43/A OR2X1_LOC_55/a_36_216# 0.00fF
C52048 OR2X1_LOC_45/B OR2X1_LOC_171/a_8_216# 0.06fF
C52049 AND2X1_LOC_91/B OR2X1_LOC_175/Y 0.07fF
C52050 AND2X1_LOC_390/B OR2X1_LOC_167/Y 0.02fF
C52051 AND2X1_LOC_373/a_8_24# OR2X1_LOC_440/A 0.01fF
C52052 AND2X1_LOC_342/a_8_24# OR2X1_LOC_47/Y 0.01fF
C52053 AND2X1_LOC_117/a_8_24# D_INPUT_0 0.02fF
C52054 OR2X1_LOC_715/B AND2X1_LOC_36/Y 0.12fF
C52055 AND2X1_LOC_518/a_8_24# OR2X1_LOC_520/B 0.01fF
C52056 AND2X1_LOC_31/Y OR2X1_LOC_785/B 0.01fF
C52057 AND2X1_LOC_626/a_8_24# AND2X1_LOC_36/Y 0.04fF
C52058 AND2X1_LOC_455/a_8_24# OR2X1_LOC_428/A 0.01fF
C52059 AND2X1_LOC_7/B OR2X1_LOC_563/A 0.01fF
C52060 OR2X1_LOC_863/B AND2X1_LOC_821/a_8_24# 0.23fF
C52061 OR2X1_LOC_520/B AND2X1_LOC_48/A 0.12fF
C52062 OR2X1_LOC_561/Y OR2X1_LOC_579/a_8_216# 0.01fF
C52063 OR2X1_LOC_87/A OR2X1_LOC_215/a_8_216# 0.04fF
C52064 OR2X1_LOC_36/Y OR2X1_LOC_511/a_8_216# 0.01fF
C52065 OR2X1_LOC_47/Y AND2X1_LOC_610/a_36_24# 0.01fF
C52066 OR2X1_LOC_224/Y OR2X1_LOC_89/A 0.03fF
C52067 OR2X1_LOC_616/Y AND2X1_LOC_805/a_36_24# 0.00fF
C52068 AND2X1_LOC_22/Y OR2X1_LOC_139/A 0.03fF
C52069 AND2X1_LOC_641/a_8_24# AND2X1_LOC_650/Y 0.20fF
C52070 OR2X1_LOC_280/a_36_216# OR2X1_LOC_47/Y 0.03fF
C52071 AND2X1_LOC_91/B OR2X1_LOC_713/A 0.14fF
C52072 OR2X1_LOC_831/a_8_216# OR2X1_LOC_318/B 0.01fF
C52073 OR2X1_LOC_865/B OR2X1_LOC_561/B 0.07fF
C52074 OR2X1_LOC_391/A OR2X1_LOC_561/A 0.01fF
C52075 OR2X1_LOC_212/A AND2X1_LOC_31/Y 0.96fF
C52076 OR2X1_LOC_379/Y OR2X1_LOC_198/A 0.02fF
C52077 OR2X1_LOC_506/A OR2X1_LOC_68/B 0.02fF
C52078 OR2X1_LOC_233/a_8_216# D_INPUT_1 0.01fF
C52079 OR2X1_LOC_756/B OR2X1_LOC_544/B 0.01fF
C52080 AND2X1_LOC_4/a_8_24# D_INPUT_1 0.00fF
C52081 OR2X1_LOC_50/a_8_216# OR2X1_LOC_17/Y 0.01fF
C52082 AND2X1_LOC_358/Y OR2X1_LOC_135/Y 0.21fF
C52083 AND2X1_LOC_483/a_8_24# AND2X1_LOC_620/Y 0.00fF
C52084 AND2X1_LOC_82/a_8_24# OR2X1_LOC_68/B 0.02fF
C52085 OR2X1_LOC_687/Y AND2X1_LOC_31/Y 0.06fF
C52086 AND2X1_LOC_555/Y OR2X1_LOC_600/A 0.03fF
C52087 VDD OR2X1_LOC_502/Y 0.08fF
C52088 OR2X1_LOC_761/Y OR2X1_LOC_13/B 0.06fF
C52089 OR2X1_LOC_258/Y AND2X1_LOC_792/Y 0.00fF
C52090 OR2X1_LOC_44/Y AND2X1_LOC_563/Y 0.17fF
C52091 AND2X1_LOC_806/A AND2X1_LOC_562/Y 0.01fF
C52092 AND2X1_LOC_95/Y OR2X1_LOC_728/A 0.01fF
C52093 OR2X1_LOC_96/a_36_216# OR2X1_LOC_46/A 0.00fF
C52094 OR2X1_LOC_161/B OR2X1_LOC_162/a_8_216# 0.01fF
C52095 OR2X1_LOC_114/Y OR2X1_LOC_560/A 0.02fF
C52096 OR2X1_LOC_787/Y OR2X1_LOC_318/B 0.01fF
C52097 AND2X1_LOC_256/a_8_24# OR2X1_LOC_549/A 0.01fF
C52098 AND2X1_LOC_3/Y OR2X1_LOC_358/A 0.06fF
C52099 OR2X1_LOC_258/Y AND2X1_LOC_259/a_8_24# 0.05fF
C52100 AND2X1_LOC_803/B AND2X1_LOC_544/Y 0.03fF
C52101 OR2X1_LOC_62/A OR2X1_LOC_62/B 0.42fF
C52102 OR2X1_LOC_186/Y OR2X1_LOC_112/a_8_216# 0.14fF
C52103 OR2X1_LOC_495/Y OR2X1_LOC_142/Y 0.06fF
C52104 OR2X1_LOC_643/a_8_216# OR2X1_LOC_228/Y 0.02fF
C52105 OR2X1_LOC_134/Y OR2X1_LOC_56/A 0.02fF
C52106 AND2X1_LOC_776/Y OR2X1_LOC_59/Y 0.78fF
C52107 OR2X1_LOC_715/B OR2X1_LOC_506/Y 0.10fF
C52108 OR2X1_LOC_486/a_8_216# OR2X1_LOC_705/B 0.48fF
C52109 INPUT_0 OR2X1_LOC_415/Y 0.03fF
C52110 OR2X1_LOC_185/A OR2X1_LOC_590/Y 0.01fF
C52111 AND2X1_LOC_719/Y AND2X1_LOC_542/a_8_24# 0.11fF
C52112 OR2X1_LOC_218/Y OR2X1_LOC_222/a_8_216# 0.06fF
C52113 AND2X1_LOC_711/A OR2X1_LOC_759/a_8_216# 0.01fF
C52114 OR2X1_LOC_45/B AND2X1_LOC_500/Y 0.03fF
C52115 OR2X1_LOC_53/Y OR2X1_LOC_25/Y 0.09fF
C52116 AND2X1_LOC_56/B OR2X1_LOC_181/a_8_216# 0.06fF
C52117 OR2X1_LOC_177/Y OR2X1_LOC_40/Y 0.02fF
C52118 AND2X1_LOC_43/B OR2X1_LOC_535/a_8_216# 0.03fF
C52119 OR2X1_LOC_576/A OR2X1_LOC_244/Y 0.05fF
C52120 AND2X1_LOC_3/Y OR2X1_LOC_460/A 0.00fF
C52121 AND2X1_LOC_541/Y AND2X1_LOC_362/B 0.03fF
C52122 OR2X1_LOC_833/Y AND2X1_LOC_18/Y 0.02fF
C52123 OR2X1_LOC_516/Y OR2X1_LOC_427/A 0.07fF
C52124 AND2X1_LOC_775/a_36_24# OR2X1_LOC_427/A 0.00fF
C52125 AND2X1_LOC_70/Y AND2X1_LOC_433/a_8_24# 0.04fF
C52126 OR2X1_LOC_255/a_36_216# AND2X1_LOC_721/A 0.00fF
C52127 OR2X1_LOC_78/B AND2X1_LOC_44/Y 2.48fF
C52128 OR2X1_LOC_139/A OR2X1_LOC_244/B 0.01fF
C52129 AND2X1_LOC_794/B VDD 0.38fF
C52130 OR2X1_LOC_753/A OR2X1_LOC_13/B 0.10fF
C52131 AND2X1_LOC_64/Y OR2X1_LOC_608/a_8_216# 0.01fF
C52132 OR2X1_LOC_287/A OR2X1_LOC_580/B 0.35fF
C52133 OR2X1_LOC_756/B OR2X1_LOC_474/B 0.01fF
C52134 OR2X1_LOC_16/A AND2X1_LOC_434/Y 0.30fF
C52135 INPUT_0 AND2X1_LOC_786/Y 0.02fF
C52136 OR2X1_LOC_16/A AND2X1_LOC_219/Y 0.02fF
C52137 OR2X1_LOC_604/A OR2X1_LOC_40/Y 0.68fF
C52138 OR2X1_LOC_40/Y OR2X1_LOC_745/a_8_216# 0.01fF
C52139 OR2X1_LOC_218/Y OR2X1_LOC_205/Y 0.03fF
C52140 OR2X1_LOC_40/Y AND2X1_LOC_758/a_8_24# 0.06fF
C52141 OR2X1_LOC_844/Y OR2X1_LOC_560/A 0.09fF
C52142 OR2X1_LOC_104/a_8_216# OR2X1_LOC_671/Y 0.39fF
C52143 OR2X1_LOC_155/A OR2X1_LOC_730/B 0.46fF
C52144 AND2X1_LOC_346/a_36_24# OR2X1_LOC_600/A 0.00fF
C52145 OR2X1_LOC_161/A OR2X1_LOC_356/B 0.19fF
C52146 AND2X1_LOC_347/Y OR2X1_LOC_428/A 0.02fF
C52147 VDD OR2X1_LOC_302/A -0.00fF
C52148 AND2X1_LOC_64/Y OR2X1_LOC_185/A 0.59fF
C52149 AND2X1_LOC_40/Y AND2X1_LOC_60/a_8_24# 0.17fF
C52150 OR2X1_LOC_721/Y AND2X1_LOC_44/Y 0.68fF
C52151 AND2X1_LOC_512/Y AND2X1_LOC_810/B 0.00fF
C52152 AND2X1_LOC_47/Y AND2X1_LOC_497/a_36_24# 0.00fF
C52153 OR2X1_LOC_217/Y OR2X1_LOC_510/a_8_216# 0.06fF
C52154 OR2X1_LOC_448/a_8_216# AND2X1_LOC_44/Y 0.01fF
C52155 OR2X1_LOC_22/Y AND2X1_LOC_570/a_36_24# 0.01fF
C52156 AND2X1_LOC_722/A AND2X1_LOC_212/Y 0.07fF
C52157 OR2X1_LOC_39/A AND2X1_LOC_783/B 0.01fF
C52158 AND2X1_LOC_552/a_8_24# OR2X1_LOC_109/Y 0.02fF
C52159 OR2X1_LOC_600/A OR2X1_LOC_51/Y 0.41fF
C52160 OR2X1_LOC_427/A OR2X1_LOC_373/a_8_216# 0.02fF
C52161 OR2X1_LOC_278/A OR2X1_LOC_71/A 0.01fF
C52162 OR2X1_LOC_175/Y OR2X1_LOC_799/A 0.14fF
C52163 AND2X1_LOC_717/Y AND2X1_LOC_786/Y 0.02fF
C52164 OR2X1_LOC_474/Y AND2X1_LOC_65/A 0.03fF
C52165 AND2X1_LOC_554/a_8_24# AND2X1_LOC_573/A 0.01fF
C52166 OR2X1_LOC_308/a_8_216# OR2X1_LOC_713/A 0.02fF
C52167 OR2X1_LOC_31/Y OR2X1_LOC_72/Y 0.03fF
C52168 OR2X1_LOC_604/A OR2X1_LOC_698/a_8_216# 0.03fF
C52169 OR2X1_LOC_256/A AND2X1_LOC_657/A 0.07fF
C52170 OR2X1_LOC_805/A OR2X1_LOC_563/A 0.07fF
C52171 OR2X1_LOC_532/B OR2X1_LOC_80/A 0.46fF
C52172 OR2X1_LOC_816/a_8_216# OR2X1_LOC_56/A 0.02fF
C52173 OR2X1_LOC_815/Y AND2X1_LOC_792/Y 0.03fF
C52174 OR2X1_LOC_284/a_8_216# OR2X1_LOC_78/A 0.02fF
C52175 AND2X1_LOC_462/Y OR2X1_LOC_68/B 0.01fF
C52176 VDD OR2X1_LOC_98/A -0.00fF
C52177 OR2X1_LOC_866/B OR2X1_LOC_848/A 0.28fF
C52178 OR2X1_LOC_486/B OR2X1_LOC_209/A 0.04fF
C52179 OR2X1_LOC_615/Y OR2X1_LOC_754/Y 0.02fF
C52180 OR2X1_LOC_375/A AND2X1_LOC_44/Y 1.12fF
C52181 AND2X1_LOC_92/a_36_24# AND2X1_LOC_43/B 0.01fF
C52182 OR2X1_LOC_494/Y AND2X1_LOC_456/B 0.47fF
C52183 VDD OR2X1_LOC_677/Y 0.28fF
C52184 INPUT_0 AND2X1_LOC_218/Y 0.12fF
C52185 AND2X1_LOC_363/Y AND2X1_LOC_456/B 0.02fF
C52186 OR2X1_LOC_866/B OR2X1_LOC_859/B 0.15fF
C52187 VDD AND2X1_LOC_208/B 0.04fF
C52188 OR2X1_LOC_36/Y AND2X1_LOC_476/a_8_24# 0.01fF
C52189 OR2X1_LOC_227/Y OR2X1_LOC_68/B 0.00fF
C52190 OR2X1_LOC_306/a_8_216# OR2X1_LOC_829/A 0.16fF
C52191 AND2X1_LOC_729/Y AND2X1_LOC_724/A 0.01fF
C52192 OR2X1_LOC_786/Y AND2X1_LOC_31/Y 0.05fF
C52193 OR2X1_LOC_148/a_8_216# OR2X1_LOC_148/B 0.47fF
C52194 OR2X1_LOC_779/Y OR2X1_LOC_779/B 0.02fF
C52195 OR2X1_LOC_485/Y OR2X1_LOC_485/a_36_216# 0.00fF
C52196 OR2X1_LOC_526/Y OR2X1_LOC_485/a_8_216# 0.01fF
C52197 OR2X1_LOC_529/a_8_216# AND2X1_LOC_362/B 0.47fF
C52198 AND2X1_LOC_845/Y OR2X1_LOC_13/B 0.01fF
C52199 AND2X1_LOC_59/Y OR2X1_LOC_346/A 0.07fF
C52200 AND2X1_LOC_727/Y AND2X1_LOC_191/Y 0.04fF
C52201 OR2X1_LOC_667/Y AND2X1_LOC_860/A 0.04fF
C52202 OR2X1_LOC_697/Y OR2X1_LOC_744/A 0.00fF
C52203 OR2X1_LOC_145/a_36_216# AND2X1_LOC_213/B 0.00fF
C52204 AND2X1_LOC_50/Y AND2X1_LOC_2/Y 0.03fF
C52205 D_INPUT_1 OR2X1_LOC_68/B 1.05fF
C52206 OR2X1_LOC_97/A AND2X1_LOC_8/Y 0.05fF
C52207 OR2X1_LOC_369/a_8_216# AND2X1_LOC_841/B 0.05fF
C52208 AND2X1_LOC_690/a_8_24# OR2X1_LOC_66/A 0.17fF
C52209 AND2X1_LOC_753/B AND2X1_LOC_70/Y 0.07fF
C52210 OR2X1_LOC_756/B OR2X1_LOC_561/Y 0.85fF
C52211 OR2X1_LOC_316/Y AND2X1_LOC_476/Y 0.00fF
C52212 OR2X1_LOC_696/A AND2X1_LOC_523/Y 0.21fF
C52213 OR2X1_LOC_185/A AND2X1_LOC_86/a_8_24# 0.02fF
C52214 AND2X1_LOC_727/Y AND2X1_LOC_711/Y 0.03fF
C52215 AND2X1_LOC_776/Y OR2X1_LOC_70/Y 0.26fF
C52216 OR2X1_LOC_756/B OR2X1_LOC_78/Y 0.08fF
C52217 OR2X1_LOC_217/Y AND2X1_LOC_65/A 0.02fF
C52218 OR2X1_LOC_114/B AND2X1_LOC_297/a_8_24# 0.01fF
C52219 OR2X1_LOC_61/B AND2X1_LOC_92/Y 0.03fF
C52220 OR2X1_LOC_270/a_36_216# OR2X1_LOC_549/A 0.00fF
C52221 OR2X1_LOC_244/B OR2X1_LOC_244/a_8_216# 0.02fF
C52222 VDD OR2X1_LOC_829/a_8_216# 0.00fF
C52223 OR2X1_LOC_61/a_8_216# OR2X1_LOC_78/B 0.30fF
C52224 AND2X1_LOC_217/Y OR2X1_LOC_65/B 0.29fF
C52225 OR2X1_LOC_296/Y OR2X1_LOC_563/A 0.00fF
C52226 AND2X1_LOC_532/a_8_24# AND2X1_LOC_436/Y 0.00fF
C52227 OR2X1_LOC_671/Y OR2X1_LOC_6/A 0.19fF
C52228 OR2X1_LOC_566/a_8_216# OR2X1_LOC_365/B 0.01fF
C52229 OR2X1_LOC_691/a_8_216# OR2X1_LOC_269/B 0.04fF
C52230 AND2X1_LOC_755/a_8_24# VDD 0.00fF
C52231 OR2X1_LOC_109/Y AND2X1_LOC_326/B 0.01fF
C52232 AND2X1_LOC_95/Y OR2X1_LOC_35/a_36_216# 0.00fF
C52233 OR2X1_LOC_35/B OR2X1_LOC_338/A 0.03fF
C52234 AND2X1_LOC_539/Y AND2X1_LOC_729/B 0.73fF
C52235 OR2X1_LOC_405/A AND2X1_LOC_70/Y 0.54fF
C52236 OR2X1_LOC_347/B OR2X1_LOC_66/A 0.03fF
C52237 VDD OR2X1_LOC_315/Y 0.20fF
C52238 OR2X1_LOC_51/Y OR2X1_LOC_619/Y 0.05fF
C52239 OR2X1_LOC_691/A AND2X1_LOC_822/a_8_24# 0.08fF
C52240 OR2X1_LOC_312/Y OR2X1_LOC_323/Y 0.42fF
C52241 OR2X1_LOC_49/A AND2X1_LOC_19/a_36_24# 0.00fF
C52242 OR2X1_LOC_491/a_36_216# OR2X1_LOC_36/Y 0.02fF
C52243 AND2X1_LOC_361/a_8_24# OR2X1_LOC_26/Y 0.01fF
C52244 OR2X1_LOC_510/A OR2X1_LOC_217/Y 1.95fF
C52245 OR2X1_LOC_160/A OR2X1_LOC_641/Y 0.07fF
C52246 OR2X1_LOC_539/Y OR2X1_LOC_66/A 0.08fF
C52247 OR2X1_LOC_160/B OR2X1_LOC_553/A 0.50fF
C52248 OR2X1_LOC_147/B AND2X1_LOC_41/A 0.75fF
C52249 AND2X1_LOC_353/a_8_24# OR2X1_LOC_36/Y -0.01fF
C52250 OR2X1_LOC_6/B OR2X1_LOC_87/A 0.07fF
C52251 OR2X1_LOC_589/A OR2X1_LOC_262/Y 0.17fF
C52252 OR2X1_LOC_267/a_8_216# OR2X1_LOC_641/A 0.08fF
C52253 OR2X1_LOC_680/A OR2X1_LOC_600/A 0.06fF
C52254 OR2X1_LOC_382/Y AND2X1_LOC_348/A 0.11fF
C52255 AND2X1_LOC_510/A AND2X1_LOC_573/A 0.01fF
C52256 OR2X1_LOC_632/A OR2X1_LOC_78/A 0.01fF
C52257 OR2X1_LOC_446/a_8_216# OR2X1_LOC_161/B 0.01fF
C52258 AND2X1_LOC_570/Y OR2X1_LOC_39/A 0.02fF
C52259 OR2X1_LOC_331/A OR2X1_LOC_39/A 0.43fF
C52260 OR2X1_LOC_273/a_36_216# AND2X1_LOC_786/Y 0.01fF
C52261 AND2X1_LOC_621/Y AND2X1_LOC_443/Y 0.03fF
C52262 AND2X1_LOC_741/a_8_24# OR2X1_LOC_441/Y 0.23fF
C52263 AND2X1_LOC_82/Y OR2X1_LOC_402/a_8_216# 0.01fF
C52264 OR2X1_LOC_185/Y OR2X1_LOC_676/Y 0.07fF
C52265 OR2X1_LOC_109/Y AND2X1_LOC_471/Y 0.03fF
C52266 OR2X1_LOC_779/a_8_216# OR2X1_LOC_66/A 0.01fF
C52267 AND2X1_LOC_862/A AND2X1_LOC_663/A 0.45fF
C52268 OR2X1_LOC_526/Y OR2X1_LOC_44/Y 0.00fF
C52269 AND2X1_LOC_718/a_8_24# OR2X1_LOC_48/B -0.01fF
C52270 VDD AND2X1_LOC_267/a_8_24# 0.00fF
C52271 AND2X1_LOC_624/A AND2X1_LOC_663/A 1.24fF
C52272 AND2X1_LOC_95/Y OR2X1_LOC_735/a_8_216# 0.01fF
C52273 AND2X1_LOC_47/Y AND2X1_LOC_235/a_8_24# 0.03fF
C52274 OR2X1_LOC_864/A OR2X1_LOC_641/a_8_216# 0.06fF
C52275 OR2X1_LOC_744/A AND2X1_LOC_648/a_36_24# 0.00fF
C52276 OR2X1_LOC_3/Y OR2X1_LOC_421/Y 0.01fF
C52277 VDD OR2X1_LOC_491/Y 0.12fF
C52278 OR2X1_LOC_6/B AND2X1_LOC_19/a_8_24# 0.03fF
C52279 OR2X1_LOC_329/Y AND2X1_LOC_356/B 0.02fF
C52280 OR2X1_LOC_40/Y AND2X1_LOC_857/a_36_24# -0.00fF
C52281 VDD OR2X1_LOC_836/B -0.00fF
C52282 OR2X1_LOC_64/Y AND2X1_LOC_786/Y 0.09fF
C52283 AND2X1_LOC_523/Y OR2X1_LOC_522/a_36_216# 0.00fF
C52284 OR2X1_LOC_190/A OR2X1_LOC_269/B 0.03fF
C52285 OR2X1_LOC_389/B OR2X1_LOC_389/A 0.00fF
C52286 OR2X1_LOC_699/a_8_216# OR2X1_LOC_56/A 0.02fF
C52287 OR2X1_LOC_532/B OR2X1_LOC_115/B 0.03fF
C52288 OR2X1_LOC_160/B OR2X1_LOC_219/B 0.52fF
C52289 VDD OR2X1_LOC_251/Y 0.42fF
C52290 OR2X1_LOC_604/A OR2X1_LOC_7/A 1.96fF
C52291 OR2X1_LOC_185/A OR2X1_LOC_464/A 0.02fF
C52292 AND2X1_LOC_777/a_36_24# OR2X1_LOC_426/B 0.01fF
C52293 OR2X1_LOC_302/B AND2X1_LOC_56/B 0.15fF
C52294 OR2X1_LOC_574/A AND2X1_LOC_18/Y 0.10fF
C52295 AND2X1_LOC_722/A AND2X1_LOC_447/a_8_24# 0.08fF
C52296 OR2X1_LOC_2/a_8_216# D_INPUT_6 0.01fF
C52297 OR2X1_LOC_203/Y AND2X1_LOC_628/a_8_24# 0.01fF
C52298 OR2X1_LOC_53/Y AND2X1_LOC_196/Y 0.38fF
C52299 OR2X1_LOC_160/A OR2X1_LOC_808/B 0.10fF
C52300 OR2X1_LOC_264/Y OR2X1_LOC_559/B 0.01fF
C52301 AND2X1_LOC_560/B AND2X1_LOC_218/Y 0.18fF
C52302 AND2X1_LOC_174/a_8_24# AND2X1_LOC_654/B 0.01fF
C52303 OR2X1_LOC_624/A OR2X1_LOC_623/B 0.08fF
C52304 AND2X1_LOC_214/A OR2X1_LOC_6/A 0.00fF
C52305 OR2X1_LOC_497/Y AND2X1_LOC_858/B 0.10fF
C52306 OR2X1_LOC_235/B OR2X1_LOC_673/Y -0.00fF
C52307 OR2X1_LOC_756/B OR2X1_LOC_285/A 0.01fF
C52308 OR2X1_LOC_501/B OR2X1_LOC_631/B 0.03fF
C52309 AND2X1_LOC_704/a_8_24# OR2X1_LOC_417/Y 0.01fF
C52310 AND2X1_LOC_843/Y AND2X1_LOC_850/a_8_24# 0.09fF
C52311 OR2X1_LOC_158/A AND2X1_LOC_260/a_36_24# 0.00fF
C52312 OR2X1_LOC_680/A AND2X1_LOC_862/Y 0.03fF
C52313 OR2X1_LOC_778/Y OR2X1_LOC_778/B 0.86fF
C52314 AND2X1_LOC_350/a_36_24# AND2X1_LOC_350/Y 0.00fF
C52315 AND2X1_LOC_351/a_36_24# OR2X1_LOC_46/A 0.00fF
C52316 AND2X1_LOC_570/Y OR2X1_LOC_239/a_36_216# 0.00fF
C52317 AND2X1_LOC_80/a_8_24# OR2X1_LOC_502/A 0.01fF
C52318 AND2X1_LOC_367/B OR2X1_LOC_89/A 0.01fF
C52319 INPUT_5 AND2X1_LOC_1/a_8_24# 0.01fF
C52320 AND2X1_LOC_336/a_8_24# AND2X1_LOC_434/Y 0.04fF
C52321 OR2X1_LOC_592/A OR2X1_LOC_468/A 0.01fF
C52322 OR2X1_LOC_702/A AND2X1_LOC_110/a_8_24# 0.18fF
C52323 OR2X1_LOC_633/Y OR2X1_LOC_610/a_36_216# 0.02fF
C52324 AND2X1_LOC_176/a_8_24# OR2X1_LOC_66/A 0.01fF
C52325 D_INPUT_0 OR2X1_LOC_548/a_8_216# 0.01fF
C52326 AND2X1_LOC_50/Y AND2X1_LOC_26/a_8_24# 0.01fF
C52327 VDD OR2X1_LOC_826/a_8_216# 0.00fF
C52328 OR2X1_LOC_705/B OR2X1_LOC_308/Y 0.14fF
C52329 OR2X1_LOC_738/B OR2X1_LOC_738/A 0.15fF
C52330 OR2X1_LOC_417/A AND2X1_LOC_786/Y 0.07fF
C52331 AND2X1_LOC_318/Y AND2X1_LOC_473/Y 0.02fF
C52332 AND2X1_LOC_554/B OR2X1_LOC_744/A 0.64fF
C52333 OR2X1_LOC_232/a_36_216# OR2X1_LOC_234/Y 0.00fF
C52334 AND2X1_LOC_31/Y OR2X1_LOC_181/Y 0.08fF
C52335 AND2X1_LOC_753/B OR2X1_LOC_193/Y 0.25fF
C52336 AND2X1_LOC_304/a_36_24# OR2X1_LOC_269/B 0.01fF
C52337 OR2X1_LOC_79/A OR2X1_LOC_59/Y 0.01fF
C52338 AND2X1_LOC_174/a_36_24# OR2X1_LOC_619/Y 0.01fF
C52339 AND2X1_LOC_359/B OR2X1_LOC_92/Y 0.01fF
C52340 AND2X1_LOC_784/A AND2X1_LOC_716/Y 0.18fF
C52341 OR2X1_LOC_273/a_8_216# AND2X1_LOC_219/Y 0.02fF
C52342 OR2X1_LOC_598/a_8_216# OR2X1_LOC_598/A 0.04fF
C52343 AND2X1_LOC_59/Y OR2X1_LOC_161/A 0.34fF
C52344 AND2X1_LOC_387/B AND2X1_LOC_41/A 0.11fF
C52345 OR2X1_LOC_62/B OR2X1_LOC_629/B 0.00fF
C52346 AND2X1_LOC_598/a_8_24# OR2X1_LOC_48/B 0.10fF
C52347 OR2X1_LOC_346/a_8_216# AND2X1_LOC_95/Y 0.01fF
C52348 OR2X1_LOC_26/Y AND2X1_LOC_852/B 0.01fF
C52349 OR2X1_LOC_423/a_8_216# OR2X1_LOC_92/Y 0.02fF
C52350 AND2X1_LOC_784/A AND2X1_LOC_654/Y 0.03fF
C52351 AND2X1_LOC_866/A AND2X1_LOC_212/Y 0.83fF
C52352 OR2X1_LOC_223/A AND2X1_LOC_604/a_8_24# 0.01fF
C52353 AND2X1_LOC_42/B AND2X1_LOC_820/B 0.83fF
C52354 OR2X1_LOC_170/a_8_216# OR2X1_LOC_365/B 0.01fF
C52355 OR2X1_LOC_154/A AND2X1_LOC_617/a_8_24# 0.10fF
C52356 AND2X1_LOC_802/B AND2X1_LOC_810/a_36_24# 0.00fF
C52357 AND2X1_LOC_56/B OR2X1_LOC_269/a_8_216# 0.01fF
C52358 OR2X1_LOC_26/Y OR2X1_LOC_48/B 0.17fF
C52359 OR2X1_LOC_168/B AND2X1_LOC_51/Y 2.24fF
C52360 OR2X1_LOC_495/Y OR2X1_LOC_238/Y 0.85fF
C52361 AND2X1_LOC_848/Y AND2X1_LOC_668/a_8_24# 0.04fF
C52362 AND2X1_LOC_367/A OR2X1_LOC_481/A 0.00fF
C52363 OR2X1_LOC_858/a_8_216# OR2X1_LOC_814/A 0.01fF
C52364 OR2X1_LOC_433/Y OR2X1_LOC_44/Y 0.03fF
C52365 OR2X1_LOC_8/Y OR2X1_LOC_62/B 0.70fF
C52366 AND2X1_LOC_90/a_8_24# OR2X1_LOC_673/A 0.01fF
C52367 AND2X1_LOC_40/Y OR2X1_LOC_557/A 0.00fF
C52368 OR2X1_LOC_278/A OR2X1_LOC_59/Y 0.14fF
C52369 OR2X1_LOC_51/Y OR2X1_LOC_22/A 0.09fF
C52370 D_INPUT_5 OR2X1_LOC_17/Y 0.40fF
C52371 OR2X1_LOC_18/Y OR2X1_LOC_26/Y 0.19fF
C52372 OR2X1_LOC_43/A OR2X1_LOC_118/Y 0.03fF
C52373 OR2X1_LOC_641/Y OR2X1_LOC_655/A 0.03fF
C52374 OR2X1_LOC_47/Y OR2X1_LOC_12/Y 0.20fF
C52375 OR2X1_LOC_160/B OR2X1_LOC_244/A 0.07fF
C52376 OR2X1_LOC_437/A OR2X1_LOC_142/a_8_216# 0.01fF
C52377 AND2X1_LOC_212/A AND2X1_LOC_318/Y 0.02fF
C52378 OR2X1_LOC_47/Y OR2X1_LOC_766/Y 0.01fF
C52379 AND2X1_LOC_733/a_36_24# OR2X1_LOC_74/A 0.01fF
C52380 OR2X1_LOC_243/a_36_216# OR2X1_LOC_66/A 0.00fF
C52381 OR2X1_LOC_774/B OR2X1_LOC_774/a_8_216# 0.06fF
C52382 OR2X1_LOC_89/A OR2X1_LOC_48/B 0.32fF
C52383 OR2X1_LOC_648/A OR2X1_LOC_814/A 0.10fF
C52384 OR2X1_LOC_112/a_8_216# OR2X1_LOC_112/B 0.01fF
C52385 AND2X1_LOC_533/a_36_24# OR2X1_LOC_269/B 0.01fF
C52386 AND2X1_LOC_592/Y AND2X1_LOC_645/a_8_24# 0.01fF
C52387 VDD OR2X1_LOC_256/A 0.21fF
C52388 OR2X1_LOC_151/A OR2X1_LOC_473/A 0.15fF
C52389 OR2X1_LOC_3/Y OR2X1_LOC_278/Y 0.02fF
C52390 OR2X1_LOC_18/Y OR2X1_LOC_89/A 0.18fF
C52391 OR2X1_LOC_597/A OR2X1_LOC_95/Y 0.00fF
C52392 AND2X1_LOC_63/a_8_24# AND2X1_LOC_8/Y 0.04fF
C52393 OR2X1_LOC_42/a_8_216# OR2X1_LOC_6/A 0.01fF
C52394 OR2X1_LOC_377/A OR2X1_LOC_793/B 0.06fF
C52395 AND2X1_LOC_729/Y OR2X1_LOC_312/Y 0.10fF
C52396 OR2X1_LOC_405/A OR2X1_LOC_653/a_8_216# 0.01fF
C52397 OR2X1_LOC_462/B AND2X1_LOC_412/a_8_24# 0.20fF
C52398 AND2X1_LOC_266/Y AND2X1_LOC_361/A 0.08fF
C52399 OR2X1_LOC_465/B OR2X1_LOC_375/A 0.09fF
C52400 OR2X1_LOC_154/A OR2X1_LOC_849/A 0.03fF
C52401 AND2X1_LOC_342/Y OR2X1_LOC_585/A 0.18fF
C52402 AND2X1_LOC_12/Y OR2X1_LOC_787/Y 0.07fF
C52403 OR2X1_LOC_479/Y AND2X1_LOC_95/Y 0.07fF
C52404 OR2X1_LOC_565/A OR2X1_LOC_549/Y 0.04fF
C52405 AND2X1_LOC_661/A OR2X1_LOC_44/Y 0.03fF
C52406 OR2X1_LOC_744/A OR2X1_LOC_167/Y 0.00fF
C52407 OR2X1_LOC_595/Y OR2X1_LOC_16/A 0.05fF
C52408 OR2X1_LOC_232/a_8_216# OR2X1_LOC_85/A 0.01fF
C52409 OR2X1_LOC_860/a_8_216# AND2X1_LOC_51/Y -0.00fF
C52410 VDD OR2X1_LOC_674/Y 0.19fF
C52411 OR2X1_LOC_83/Y OR2X1_LOC_81/a_8_216# 0.04fF
C52412 OR2X1_LOC_617/Y AND2X1_LOC_621/Y 0.15fF
C52413 AND2X1_LOC_367/A OR2X1_LOC_71/Y 0.05fF
C52414 VDD OR2X1_LOC_845/A 0.08fF
C52415 AND2X1_LOC_784/A OR2X1_LOC_312/Y 0.07fF
C52416 AND2X1_LOC_259/Y OR2X1_LOC_44/Y 0.04fF
C52417 OR2X1_LOC_45/B AND2X1_LOC_563/Y 0.00fF
C52418 OR2X1_LOC_848/A OR2X1_LOC_557/A 0.01fF
C52419 AND2X1_LOC_7/B OR2X1_LOC_724/A 0.32fF
C52420 OR2X1_LOC_87/B AND2X1_LOC_19/a_36_24# 0.01fF
C52421 OR2X1_LOC_491/a_36_216# OR2X1_LOC_419/Y 0.17fF
C52422 OR2X1_LOC_720/B OR2X1_LOC_721/Y 0.39fF
C52423 OR2X1_LOC_318/A OR2X1_LOC_228/Y 0.01fF
C52424 AND2X1_LOC_663/B AND2X1_LOC_848/a_8_24# 0.01fF
C52425 OR2X1_LOC_840/A OR2X1_LOC_532/B 0.03fF
C52426 AND2X1_LOC_59/Y AND2X1_LOC_51/Y 0.21fF
C52427 OR2X1_LOC_759/A AND2X1_LOC_792/Y 0.00fF
C52428 OR2X1_LOC_40/Y AND2X1_LOC_805/a_8_24# 0.01fF
C52429 VDD AND2X1_LOC_624/B 0.46fF
C52430 VDD OR2X1_LOC_67/Y 0.66fF
C52431 OR2X1_LOC_175/Y OR2X1_LOC_446/B 0.05fF
C52432 AND2X1_LOC_36/Y AND2X1_LOC_619/a_8_24# 0.06fF
C52433 AND2X1_LOC_81/B OR2X1_LOC_647/Y 0.01fF
C52434 OR2X1_LOC_592/A OR2X1_LOC_449/B 0.05fF
C52435 AND2X1_LOC_70/Y OR2X1_LOC_330/a_8_216# 0.02fF
C52436 OR2X1_LOC_175/Y OR2X1_LOC_303/B 0.00fF
C52437 VDD OR2X1_LOC_551/A -0.00fF
C52438 OR2X1_LOC_151/A OR2X1_LOC_228/Y 0.07fF
C52439 AND2X1_LOC_86/Y OR2X1_LOC_244/A 0.01fF
C52440 OR2X1_LOC_520/Y OR2X1_LOC_650/Y 0.01fF
C52441 OR2X1_LOC_43/A AND2X1_LOC_855/a_8_24# 0.07fF
C52442 OR2X1_LOC_117/Y AND2X1_LOC_663/B 0.35fF
C52443 AND2X1_LOC_714/a_8_24# OR2X1_LOC_423/Y 0.01fF
C52444 OR2X1_LOC_462/B OR2X1_LOC_472/B 0.02fF
C52445 OR2X1_LOC_502/A AND2X1_LOC_109/a_8_24# 0.03fF
C52446 AND2X1_LOC_185/a_8_24# OR2X1_LOC_615/Y 0.02fF
C52447 VDD OR2X1_LOC_163/Y 0.13fF
C52448 OR2X1_LOC_837/A AND2X1_LOC_476/A 0.01fF
C52449 OR2X1_LOC_428/A OR2X1_LOC_437/A 0.38fF
C52450 OR2X1_LOC_168/Y OR2X1_LOC_388/a_8_216# 0.02fF
C52451 AND2X1_LOC_48/A OR2X1_LOC_790/a_36_216# 0.00fF
C52452 OR2X1_LOC_375/A OR2X1_LOC_720/B 0.00fF
C52453 AND2X1_LOC_8/Y OR2X1_LOC_415/A 0.04fF
C52454 OR2X1_LOC_446/B OR2X1_LOC_713/A 0.07fF
C52455 OR2X1_LOC_161/B OR2X1_LOC_140/Y 0.54fF
C52456 OR2X1_LOC_3/Y OR2X1_LOC_273/Y 0.07fF
C52457 OR2X1_LOC_763/Y OR2X1_LOC_64/Y 0.33fF
C52458 OR2X1_LOC_864/A OR2X1_LOC_643/Y 0.03fF
C52459 OR2X1_LOC_686/a_36_216# AND2X1_LOC_430/B 0.00fF
C52460 OR2X1_LOC_426/B AND2X1_LOC_222/Y 0.00fF
C52461 OR2X1_LOC_18/Y OR2X1_LOC_92/a_8_216# 0.01fF
C52462 OR2X1_LOC_580/A OR2X1_LOC_843/B 0.01fF
C52463 OR2X1_LOC_68/Y OR2X1_LOC_87/A 0.01fF
C52464 OR2X1_LOC_160/A OR2X1_LOC_218/Y 0.02fF
C52465 OR2X1_LOC_244/A OR2X1_LOC_266/a_8_216# 0.04fF
C52466 OR2X1_LOC_585/A OR2X1_LOC_54/Y 0.01fF
C52467 OR2X1_LOC_19/B AND2X1_LOC_234/a_36_24# 0.01fF
C52468 OR2X1_LOC_84/B OR2X1_LOC_62/B 0.00fF
C52469 AND2X1_LOC_34/Y AND2X1_LOC_476/A 0.19fF
C52470 AND2X1_LOC_578/A OR2X1_LOC_64/Y 0.07fF
C52471 AND2X1_LOC_817/B OR2X1_LOC_770/a_36_216# 0.00fF
C52472 OR2X1_LOC_47/Y OR2X1_LOC_393/Y 0.34fF
C52473 OR2X1_LOC_87/A AND2X1_LOC_47/Y 0.14fF
C52474 AND2X1_LOC_170/a_8_24# OR2X1_LOC_47/Y 0.00fF
C52475 OR2X1_LOC_3/Y OR2X1_LOC_19/B 0.70fF
C52476 OR2X1_LOC_141/B OR2X1_LOC_62/B 0.01fF
C52477 OR2X1_LOC_767/Y AND2X1_LOC_773/a_8_24# 0.23fF
C52478 OR2X1_LOC_473/Y OR2X1_LOC_215/A 0.03fF
C52479 AND2X1_LOC_56/B AND2X1_LOC_613/a_8_24# 0.01fF
C52480 OR2X1_LOC_694/a_8_216# OR2X1_LOC_47/Y 0.01fF
C52481 AND2X1_LOC_390/a_8_24# OR2X1_LOC_13/B 0.02fF
C52482 OR2X1_LOC_56/A OR2X1_LOC_521/a_8_216# 0.03fF
C52483 AND2X1_LOC_319/A AND2X1_LOC_648/B 0.03fF
C52484 AND2X1_LOC_456/Y OR2X1_LOC_71/Y 0.35fF
C52485 INPUT_0 OR2X1_LOC_460/A 0.01fF
C52486 OR2X1_LOC_78/A OR2X1_LOC_71/A 0.03fF
C52487 OR2X1_LOC_70/A OR2X1_LOC_59/a_8_216# 0.01fF
C52488 OR2X1_LOC_490/Y OR2X1_LOC_71/Y 0.15fF
C52489 OR2X1_LOC_36/Y OR2X1_LOC_615/Y 0.07fF
C52490 OR2X1_LOC_711/a_36_216# AND2X1_LOC_36/Y 0.02fF
C52491 OR2X1_LOC_92/Y AND2X1_LOC_790/a_8_24# 0.01fF
C52492 OR2X1_LOC_744/Y AND2X1_LOC_783/B 0.78fF
C52493 OR2X1_LOC_110/a_36_216# AND2X1_LOC_786/Y 0.01fF
C52494 AND2X1_LOC_84/Y AND2X1_LOC_206/a_8_24# 0.01fF
C52495 AND2X1_LOC_578/A OR2X1_LOC_417/A 0.27fF
C52496 OR2X1_LOC_864/A OR2X1_LOC_786/Y 0.03fF
C52497 AND2X1_LOC_486/Y AND2X1_LOC_657/A 0.10fF
C52498 AND2X1_LOC_31/Y OR2X1_LOC_725/B 0.01fF
C52499 AND2X1_LOC_721/A OR2X1_LOC_248/a_8_216# 0.01fF
C52500 OR2X1_LOC_449/A OR2X1_LOC_783/a_8_216# 0.49fF
C52501 OR2X1_LOC_737/A OR2X1_LOC_68/B 0.15fF
C52502 OR2X1_LOC_214/B OR2X1_LOC_269/B 0.07fF
C52503 OR2X1_LOC_158/A OR2X1_LOC_743/Y 0.01fF
C52504 AND2X1_LOC_633/Y OR2X1_LOC_46/A 0.02fF
C52505 OR2X1_LOC_427/A AND2X1_LOC_793/B 0.01fF
C52506 OR2X1_LOC_633/B OR2X1_LOC_786/Y 0.93fF
C52507 OR2X1_LOC_696/Y OR2X1_LOC_31/Y 0.03fF
C52508 OR2X1_LOC_269/B OR2X1_LOC_241/B 0.13fF
C52509 AND2X1_LOC_95/Y OR2X1_LOC_68/B 0.12fF
C52510 OR2X1_LOC_563/A OR2X1_LOC_580/B 0.07fF
C52511 OR2X1_LOC_87/A OR2X1_LOC_598/A 0.10fF
C52512 OR2X1_LOC_89/A AND2X1_LOC_620/Y 0.03fF
C52513 AND2X1_LOC_721/A AND2X1_LOC_294/a_8_24# 0.00fF
C52514 AND2X1_LOC_571/Y AND2X1_LOC_657/A 0.02fF
C52515 AND2X1_LOC_593/Y OR2X1_LOC_534/a_8_216# 0.12fF
C52516 D_INPUT_0 OR2X1_LOC_46/A 0.43fF
C52517 OR2X1_LOC_633/Y OR2X1_LOC_68/B 0.38fF
C52518 AND2X1_LOC_287/a_36_24# AND2X1_LOC_562/Y 0.06fF
C52519 INPUT_1 OR2X1_LOC_77/a_8_216# 0.05fF
C52520 OR2X1_LOC_609/A AND2X1_LOC_647/B 0.03fF
C52521 OR2X1_LOC_429/Y OR2X1_LOC_51/a_36_216# 0.01fF
C52522 OR2X1_LOC_74/A D_INPUT_1 0.05fF
C52523 OR2X1_LOC_175/Y OR2X1_LOC_863/A 0.04fF
C52524 OR2X1_LOC_655/B OR2X1_LOC_649/a_36_216# 0.00fF
C52525 OR2X1_LOC_828/B AND2X1_LOC_31/Y 0.03fF
C52526 OR2X1_LOC_64/Y AND2X1_LOC_841/a_8_24# 0.01fF
C52527 AND2X1_LOC_785/A OR2X1_LOC_56/A 0.02fF
C52528 OR2X1_LOC_196/Y OR2X1_LOC_614/Y 0.02fF
C52529 OR2X1_LOC_835/B AND2X1_LOC_31/Y 0.07fF
C52530 OR2X1_LOC_808/B OR2X1_LOC_532/Y 0.05fF
C52531 OR2X1_LOC_528/Y AND2X1_LOC_564/B 0.19fF
C52532 OR2X1_LOC_696/A AND2X1_LOC_191/B 0.78fF
C52533 AND2X1_LOC_44/Y OR2X1_LOC_549/A 0.18fF
C52534 OR2X1_LOC_589/A AND2X1_LOC_407/a_8_24# 0.00fF
C52535 AND2X1_LOC_727/A AND2X1_LOC_318/Y 0.02fF
C52536 OR2X1_LOC_706/B AND2X1_LOC_47/Y 0.05fF
C52537 AND2X1_LOC_787/A AND2X1_LOC_719/Y 0.10fF
C52538 OR2X1_LOC_390/a_8_216# AND2X1_LOC_18/Y 0.02fF
C52539 AND2X1_LOC_672/B AND2X1_LOC_672/a_8_24# 0.11fF
C52540 OR2X1_LOC_49/A OR2X1_LOC_382/A 0.11fF
C52541 AND2X1_LOC_624/B AND2X1_LOC_624/a_8_24# 0.03fF
C52542 AND2X1_LOC_91/B AND2X1_LOC_700/a_8_24# 0.11fF
C52543 AND2X1_LOC_727/Y AND2X1_LOC_658/B 0.03fF
C52544 AND2X1_LOC_227/Y D_INPUT_0 0.03fF
C52545 AND2X1_LOC_187/a_8_24# OR2X1_LOC_742/B 0.05fF
C52546 OR2X1_LOC_45/B AND2X1_LOC_712/Y 0.02fF
C52547 OR2X1_LOC_273/a_8_216# OR2X1_LOC_595/Y 0.26fF
C52548 AND2X1_LOC_314/a_8_24# OR2X1_LOC_777/B 0.17fF
C52549 OR2X1_LOC_99/Y OR2X1_LOC_68/B 0.05fF
C52550 OR2X1_LOC_176/Y OR2X1_LOC_40/Y 0.05fF
C52551 AND2X1_LOC_75/a_8_24# OR2X1_LOC_241/B 0.04fF
C52552 OR2X1_LOC_241/Y OR2X1_LOC_532/B 0.07fF
C52553 OR2X1_LOC_106/Y OR2X1_LOC_56/A 0.04fF
C52554 OR2X1_LOC_502/A OR2X1_LOC_308/Y 0.14fF
C52555 AND2X1_LOC_841/a_8_24# OR2X1_LOC_417/A 0.04fF
C52556 AND2X1_LOC_570/Y AND2X1_LOC_456/a_8_24# 0.24fF
C52557 OR2X1_LOC_158/A AND2X1_LOC_285/a_8_24# 0.01fF
C52558 AND2X1_LOC_715/A OR2X1_LOC_428/A 0.08fF
C52559 OR2X1_LOC_40/Y AND2X1_LOC_212/Y 0.29fF
C52560 OR2X1_LOC_523/Y OR2X1_LOC_844/B 0.16fF
C52561 OR2X1_LOC_47/Y AND2X1_LOC_801/B 0.01fF
C52562 AND2X1_LOC_544/Y OR2X1_LOC_524/Y 0.43fF
C52563 AND2X1_LOC_732/B OR2X1_LOC_12/Y 0.00fF
C52564 OR2X1_LOC_161/A OR2X1_LOC_342/B 0.01fF
C52565 OR2X1_LOC_691/A OR2X1_LOC_66/A 0.79fF
C52566 OR2X1_LOC_8/Y OR2X1_LOC_15/a_36_216# 0.02fF
C52567 OR2X1_LOC_184/Y OR2X1_LOC_226/a_36_216# 0.00fF
C52568 OR2X1_LOC_97/A AND2X1_LOC_92/Y 0.10fF
C52569 AND2X1_LOC_547/Y AND2X1_LOC_547/a_36_24# 0.00fF
C52570 OR2X1_LOC_235/B OR2X1_LOC_720/Y -0.00fF
C52571 AND2X1_LOC_338/A AND2X1_LOC_334/Y 0.06fF
C52572 OR2X1_LOC_36/Y OR2X1_LOC_424/Y 0.01fF
C52573 AND2X1_LOC_784/A OR2X1_LOC_13/B 0.07fF
C52574 OR2X1_LOC_657/a_8_216# OR2X1_LOC_217/A 0.39fF
C52575 OR2X1_LOC_160/A OR2X1_LOC_703/Y 0.02fF
C52576 OR2X1_LOC_329/B AND2X1_LOC_455/B 0.00fF
C52577 OR2X1_LOC_113/Y AND2X1_LOC_44/Y 0.00fF
C52578 OR2X1_LOC_160/A OR2X1_LOC_500/a_8_216# 0.01fF
C52579 OR2X1_LOC_743/A OR2X1_LOC_423/Y 0.03fF
C52580 OR2X1_LOC_135/Y OR2X1_LOC_59/Y 0.52fF
C52581 OR2X1_LOC_216/A OR2X1_LOC_392/B 0.10fF
C52582 OR2X1_LOC_256/A OR2X1_LOC_67/Y 0.14fF
C52583 OR2X1_LOC_235/B AND2X1_LOC_277/a_8_24# 0.01fF
C52584 GATE_811 AND2X1_LOC_803/a_8_24# 0.00fF
C52585 OR2X1_LOC_494/A AND2X1_LOC_348/A 0.27fF
C52586 OR2X1_LOC_154/A AND2X1_LOC_238/a_8_24# 0.02fF
C52587 OR2X1_LOC_793/A AND2X1_LOC_36/Y 0.17fF
C52588 OR2X1_LOC_71/Y AND2X1_LOC_647/Y 0.03fF
C52589 AND2X1_LOC_425/Y AND2X1_LOC_430/B 1.50fF
C52590 AND2X1_LOC_320/a_8_24# OR2X1_LOC_151/A 0.03fF
C52591 AND2X1_LOC_705/Y AND2X1_LOC_605/Y 0.00fF
C52592 OR2X1_LOC_121/Y AND2X1_LOC_41/A 0.01fF
C52593 OR2X1_LOC_744/A AND2X1_LOC_476/Y 0.07fF
C52594 AND2X1_LOC_362/B OR2X1_LOC_744/A 1.49fF
C52595 VDD OR2X1_LOC_60/Y 0.16fF
C52596 OR2X1_LOC_526/Y AND2X1_LOC_705/a_8_24# 0.08fF
C52597 AND2X1_LOC_508/B AND2X1_LOC_807/B 0.83fF
C52598 AND2X1_LOC_91/B AND2X1_LOC_314/a_36_24# 0.01fF
C52599 OR2X1_LOC_756/B OR2X1_LOC_343/a_8_216# 0.02fF
C52600 OR2X1_LOC_45/B OR2X1_LOC_422/Y 0.01fF
C52601 OR2X1_LOC_505/Y OR2X1_LOC_56/A 0.01fF
C52602 AND2X1_LOC_861/a_8_24# AND2X1_LOC_807/B 0.03fF
C52603 OR2X1_LOC_74/A AND2X1_LOC_789/Y 0.02fF
C52604 OR2X1_LOC_687/Y AND2X1_LOC_760/a_8_24# 0.02fF
C52605 OR2X1_LOC_51/Y AND2X1_LOC_286/a_8_24# 0.01fF
C52606 OR2X1_LOC_757/A OR2X1_LOC_600/A 0.05fF
C52607 AND2X1_LOC_738/B AND2X1_LOC_658/A 0.07fF
C52608 AND2X1_LOC_22/Y OR2X1_LOC_655/a_36_216# 0.01fF
C52609 AND2X1_LOC_658/A OR2X1_LOC_56/A 0.10fF
C52610 AND2X1_LOC_179/a_8_24# OR2X1_LOC_741/Y 0.08fF
C52611 OR2X1_LOC_130/A OR2X1_LOC_338/A 0.02fF
C52612 OR2X1_LOC_709/A AND2X1_LOC_423/a_36_24# 0.01fF
C52613 OR2X1_LOC_691/A AND2X1_LOC_690/a_36_24# 0.00fF
C52614 OR2X1_LOC_6/B AND2X1_LOC_54/a_36_24# 0.00fF
C52615 AND2X1_LOC_486/Y AND2X1_LOC_794/B 0.01fF
C52616 AND2X1_LOC_494/a_8_24# OR2X1_LOC_558/A 0.01fF
C52617 OR2X1_LOC_387/Y OR2X1_LOC_387/A 0.05fF
C52618 OR2X1_LOC_625/Y OR2X1_LOC_12/Y 0.10fF
C52619 AND2X1_LOC_794/A AND2X1_LOC_212/Y 0.03fF
C52620 AND2X1_LOC_647/Y D_INPUT_1 0.02fF
C52621 OR2X1_LOC_858/A OR2X1_LOC_78/A 0.12fF
C52622 AND2X1_LOC_712/a_8_24# AND2X1_LOC_454/Y 0.21fF
C52623 OR2X1_LOC_49/A OR2X1_LOC_160/A 0.11fF
C52624 OR2X1_LOC_261/A AND2X1_LOC_789/Y 0.00fF
C52625 OR2X1_LOC_175/Y AND2X1_LOC_56/B 0.07fF
C52626 OR2X1_LOC_36/Y AND2X1_LOC_242/B 0.09fF
C52627 AND2X1_LOC_573/A AND2X1_LOC_249/a_8_24# 0.02fF
C52628 OR2X1_LOC_505/a_8_216# OR2X1_LOC_39/A 0.01fF
C52629 AND2X1_LOC_367/A OR2X1_LOC_426/B 0.10fF
C52630 OR2X1_LOC_737/a_8_216# OR2X1_LOC_741/A -0.00fF
C52631 OR2X1_LOC_6/B OR2X1_LOC_23/a_8_216# 0.22fF
C52632 OR2X1_LOC_541/A AND2X1_LOC_92/Y 0.03fF
C52633 AND2X1_LOC_84/Y OR2X1_LOC_52/B 0.90fF
C52634 AND2X1_LOC_721/a_8_24# AND2X1_LOC_860/A 0.01fF
C52635 AND2X1_LOC_707/Y OR2X1_LOC_36/Y 0.01fF
C52636 AND2X1_LOC_58/a_8_24# AND2X1_LOC_18/Y 0.01fF
C52637 AND2X1_LOC_734/a_8_24# AND2X1_LOC_564/a_8_24# 0.23fF
C52638 OR2X1_LOC_406/Y AND2X1_LOC_569/A 0.09fF
C52639 OR2X1_LOC_188/Y OR2X1_LOC_269/B 0.03fF
C52640 OR2X1_LOC_858/A OR2X1_LOC_458/B 0.02fF
C52641 OR2X1_LOC_691/Y AND2X1_LOC_56/B 0.07fF
C52642 AND2X1_LOC_348/Y OR2X1_LOC_428/A 0.01fF
C52643 AND2X1_LOC_486/Y VDD 1.60fF
C52644 OR2X1_LOC_485/A AND2X1_LOC_227/a_8_24# 0.02fF
C52645 OR2X1_LOC_179/Y OR2X1_LOC_178/Y 0.21fF
C52646 OR2X1_LOC_160/A OR2X1_LOC_596/A 0.02fF
C52647 AND2X1_LOC_721/Y AND2X1_LOC_458/a_8_24# 0.01fF
C52648 OR2X1_LOC_427/A OR2X1_LOC_581/Y 0.14fF
C52649 OR2X1_LOC_339/a_36_216# AND2X1_LOC_40/Y 0.00fF
C52650 AND2X1_LOC_70/Y D_INPUT_4 0.02fF
C52651 OR2X1_LOC_753/A OR2X1_LOC_428/A 0.03fF
C52652 OR2X1_LOC_811/A OR2X1_LOC_66/A 9.53fF
C52653 AND2X1_LOC_566/B AND2X1_LOC_655/A 0.03fF
C52654 VDD AND2X1_LOC_811/B 0.21fF
C52655 AND2X1_LOC_92/Y OR2X1_LOC_475/B 0.10fF
C52656 AND2X1_LOC_340/Y OR2X1_LOC_26/Y 0.03fF
C52657 AND2X1_LOC_521/a_8_24# OR2X1_LOC_87/A 0.04fF
C52658 AND2X1_LOC_553/A OR2X1_LOC_107/a_36_216# 0.00fF
C52659 OR2X1_LOC_185/A OR2X1_LOC_776/Y 0.43fF
C52660 OR2X1_LOC_377/A AND2X1_LOC_18/Y 0.12fF
C52661 AND2X1_LOC_571/Y VDD 0.25fF
C52662 OR2X1_LOC_801/B AND2X1_LOC_751/a_8_24# 0.02fF
C52663 AND2X1_LOC_539/Y AND2X1_LOC_798/Y 0.19fF
C52664 OR2X1_LOC_490/a_36_216# OR2X1_LOC_26/Y 0.02fF
C52665 AND2X1_LOC_714/B OR2X1_LOC_44/Y 0.12fF
C52666 OR2X1_LOC_40/Y OR2X1_LOC_265/Y 0.01fF
C52667 OR2X1_LOC_115/a_8_216# AND2X1_LOC_70/Y 0.01fF
C52668 OR2X1_LOC_114/Y OR2X1_LOC_361/a_8_216# 0.01fF
C52669 AND2X1_LOC_722/A OR2X1_LOC_164/Y 0.31fF
C52670 OR2X1_LOC_58/Y OR2X1_LOC_316/Y 0.01fF
C52671 AND2X1_LOC_840/B AND2X1_LOC_476/Y 0.10fF
C52672 AND2X1_LOC_22/Y OR2X1_LOC_479/Y 0.05fF
C52673 OR2X1_LOC_604/A OR2X1_LOC_427/a_36_216# 0.00fF
C52674 OR2X1_LOC_121/Y OR2X1_LOC_217/a_36_216# 0.01fF
C52675 AND2X1_LOC_64/Y OR2X1_LOC_476/B 0.07fF
C52676 AND2X1_LOC_3/Y AND2X1_LOC_488/a_36_24# 0.00fF
C52677 OR2X1_LOC_325/A OR2X1_LOC_808/B 0.10fF
C52678 AND2X1_LOC_364/Y AND2X1_LOC_661/a_8_24# 0.00fF
C52679 AND2X1_LOC_47/Y OR2X1_LOC_844/B 0.07fF
C52680 OR2X1_LOC_604/A OR2X1_LOC_236/a_8_216# 0.03fF
C52681 AND2X1_LOC_710/Y AND2X1_LOC_847/Y 0.18fF
C52682 OR2X1_LOC_188/Y AND2X1_LOC_75/a_8_24# 0.01fF
C52683 AND2X1_LOC_572/Y AND2X1_LOC_561/B 0.03fF
C52684 OR2X1_LOC_122/a_36_216# AND2X1_LOC_99/A 0.00fF
C52685 OR2X1_LOC_329/B AND2X1_LOC_662/B 1.20fF
C52686 OR2X1_LOC_666/A OR2X1_LOC_67/A 0.01fF
C52687 AND2X1_LOC_344/a_8_24# OR2X1_LOC_92/Y 0.01fF
C52688 AND2X1_LOC_259/Y OR2X1_LOC_382/A 0.01fF
C52689 VDD AND2X1_LOC_834/a_8_24# 0.00fF
C52690 OR2X1_LOC_64/Y OR2X1_LOC_312/a_8_216# 0.01fF
C52691 AND2X1_LOC_99/Y AND2X1_LOC_99/a_36_24# 0.00fF
C52692 OR2X1_LOC_203/Y AND2X1_LOC_18/Y 0.08fF
C52693 VDD OR2X1_LOC_866/a_8_216# 0.00fF
C52694 OR2X1_LOC_502/A OR2X1_LOC_775/a_36_216# 0.00fF
C52695 OR2X1_LOC_47/Y OR2X1_LOC_248/A 0.09fF
C52696 OR2X1_LOC_524/Y AND2X1_LOC_550/A 0.02fF
C52697 OR2X1_LOC_364/A OR2X1_LOC_602/Y 0.35fF
C52698 OR2X1_LOC_574/A AND2X1_LOC_275/a_8_24# 0.22fF
C52699 OR2X1_LOC_600/A AND2X1_LOC_359/B 0.07fF
C52700 AND2X1_LOC_539/Y OR2X1_LOC_46/A 0.02fF
C52701 AND2X1_LOC_848/Y OR2X1_LOC_59/Y 0.09fF
C52702 AND2X1_LOC_392/A OR2X1_LOC_117/Y 0.43fF
C52703 OR2X1_LOC_70/Y OR2X1_LOC_135/Y 0.08fF
C52704 VDD AND2X1_LOC_740/B 0.07fF
C52705 OR2X1_LOC_696/A OR2X1_LOC_111/Y 0.07fF
C52706 AND2X1_LOC_70/Y OR2X1_LOC_653/A 0.00fF
C52707 OR2X1_LOC_51/Y OR2X1_LOC_669/A 0.04fF
C52708 AND2X1_LOC_675/Y AND2X1_LOC_624/A 0.18fF
C52709 OR2X1_LOC_756/B OR2X1_LOC_185/A 0.65fF
C52710 VDD OR2X1_LOC_248/Y 0.23fF
C52711 AND2X1_LOC_474/A AND2X1_LOC_123/Y 0.14fF
C52712 AND2X1_LOC_535/Y AND2X1_LOC_355/a_8_24# 0.01fF
C52713 AND2X1_LOC_12/Y AND2X1_LOC_41/A 13.38fF
C52714 OR2X1_LOC_624/A OR2X1_LOC_434/a_8_216# 0.11fF
C52715 AND2X1_LOC_47/Y OR2X1_LOC_390/B 0.08fF
C52716 OR2X1_LOC_756/B OR2X1_LOC_249/Y 0.00fF
C52717 OR2X1_LOC_405/A OR2X1_LOC_474/Y 0.02fF
C52718 OR2X1_LOC_380/A OR2X1_LOC_25/Y 0.19fF
C52719 OR2X1_LOC_223/A OR2X1_LOC_301/a_8_216# 0.01fF
C52720 OR2X1_LOC_831/a_8_216# OR2X1_LOC_168/B 0.07fF
C52721 OR2X1_LOC_593/a_8_216# OR2X1_LOC_78/A 0.01fF
C52722 OR2X1_LOC_158/A AND2X1_LOC_120/a_8_24# 0.01fF
C52723 OR2X1_LOC_502/A AND2X1_LOC_414/a_36_24# 0.01fF
C52724 OR2X1_LOC_862/B OR2X1_LOC_269/B 0.22fF
C52725 OR2X1_LOC_613/Y AND2X1_LOC_663/A 0.00fF
C52726 AND2X1_LOC_271/a_8_24# AND2X1_LOC_36/Y 0.01fF
C52727 VDD OR2X1_LOC_666/Y 0.05fF
C52728 OR2X1_LOC_784/a_8_216# OR2X1_LOC_66/A 0.02fF
C52729 OR2X1_LOC_50/a_8_216# INPUT_6 0.07fF
C52730 OR2X1_LOC_51/Y AND2X1_LOC_454/A 0.01fF
C52731 OR2X1_LOC_191/B OR2X1_LOC_191/a_8_216# 0.10fF
C52732 AND2X1_LOC_42/a_8_24# OR2X1_LOC_66/A 0.02fF
C52733 OR2X1_LOC_283/Y OR2X1_LOC_59/Y 0.27fF
C52734 AND2X1_LOC_350/B OR2X1_LOC_46/A 0.00fF
C52735 AND2X1_LOC_776/a_8_24# OR2X1_LOC_238/Y 0.11fF
C52736 AND2X1_LOC_59/Y OR2X1_LOC_640/A 0.16fF
C52737 OR2X1_LOC_268/a_36_216# AND2X1_LOC_786/Y 0.01fF
C52738 OR2X1_LOC_161/A OR2X1_LOC_623/B 0.00fF
C52739 AND2X1_LOC_214/A OR2X1_LOC_44/Y 0.04fF
C52740 AND2X1_LOC_366/a_8_24# OR2X1_LOC_7/A 0.01fF
C52741 AND2X1_LOC_701/a_8_24# OR2X1_LOC_78/A 0.01fF
C52742 AND2X1_LOC_141/a_8_24# OR2X1_LOC_7/A 0.02fF
C52743 OR2X1_LOC_653/Y OR2X1_LOC_624/A 0.10fF
C52744 OR2X1_LOC_677/Y AND2X1_LOC_834/a_8_24# 0.04fF
C52745 AND2X1_LOC_860/a_8_24# AND2X1_LOC_806/A 0.01fF
C52746 OR2X1_LOC_490/Y OR2X1_LOC_426/B 0.00fF
C52747 OR2X1_LOC_426/B OR2X1_LOC_74/A 0.13fF
C52748 AND2X1_LOC_845/Y OR2X1_LOC_428/A 0.02fF
C52749 OR2X1_LOC_161/A OR2X1_LOC_794/A 0.02fF
C52750 OR2X1_LOC_88/Y OR2X1_LOC_13/B 0.03fF
C52751 OR2X1_LOC_154/A OR2X1_LOC_436/B 0.01fF
C52752 OR2X1_LOC_447/Y OR2X1_LOC_713/a_36_216# 0.02fF
C52753 AND2X1_LOC_683/a_8_24# OR2X1_LOC_78/B 0.06fF
C52754 OR2X1_LOC_228/Y OR2X1_LOC_716/a_8_216# 0.05fF
C52755 INPUT_5 AND2X1_LOC_17/a_8_24# 0.01fF
C52756 OR2X1_LOC_158/A OR2X1_LOC_295/Y 0.01fF
C52757 AND2X1_LOC_727/Y OR2X1_LOC_47/Y 0.02fF
C52758 OR2X1_LOC_681/a_8_216# OR2X1_LOC_64/Y 0.01fF
C52759 OR2X1_LOC_185/A OR2X1_LOC_660/B 0.03fF
C52760 OR2X1_LOC_285/a_8_216# OR2X1_LOC_269/B 0.01fF
C52761 AND2X1_LOC_845/Y OR2X1_LOC_595/A 0.07fF
C52762 OR2X1_LOC_454/a_8_216# OR2X1_LOC_161/B 0.02fF
C52763 OR2X1_LOC_720/B OR2X1_LOC_549/A -0.02fF
C52764 OR2X1_LOC_433/Y AND2X1_LOC_435/a_8_24# 0.24fF
C52765 AND2X1_LOC_615/a_8_24# OR2X1_LOC_269/B 0.01fF
C52766 AND2X1_LOC_393/a_36_24# AND2X1_LOC_40/Y 0.01fF
C52767 AND2X1_LOC_524/a_8_24# OR2X1_LOC_545/B 0.01fF
C52768 OR2X1_LOC_629/Y AND2X1_LOC_56/B 0.17fF
C52769 AND2X1_LOC_729/Y OR2X1_LOC_679/B 0.01fF
C52770 OR2X1_LOC_532/B OR2X1_LOC_741/a_8_216# 0.04fF
C52771 OR2X1_LOC_190/B OR2X1_LOC_553/a_8_216# 0.47fF
C52772 AND2X1_LOC_348/A AND2X1_LOC_363/A 0.05fF
C52773 OR2X1_LOC_36/Y AND2X1_LOC_841/B 0.01fF
C52774 AND2X1_LOC_17/Y D_INPUT_4 0.04fF
C52775 OR2X1_LOC_609/A AND2X1_LOC_647/a_36_24# 0.00fF
C52776 AND2X1_LOC_191/B AND2X1_LOC_663/B 1.78fF
C52777 AND2X1_LOC_682/a_8_24# OR2X1_LOC_87/A 0.02fF
C52778 OR2X1_LOC_69/A OR2X1_LOC_39/A 0.03fF
C52779 AND2X1_LOC_59/Y OR2X1_LOC_541/a_8_216# 0.01fF
C52780 D_INPUT_0 OR2X1_LOC_786/a_8_216# 0.01fF
C52781 AND2X1_LOC_859/Y OR2X1_LOC_427/A 0.07fF
C52782 AND2X1_LOC_56/B AND2X1_LOC_699/a_36_24# -0.00fF
C52783 OR2X1_LOC_95/Y OR2X1_LOC_829/A 0.05fF
C52784 OR2X1_LOC_506/A OR2X1_LOC_87/A 0.02fF
C52785 OR2X1_LOC_620/Y OR2X1_LOC_778/Y 0.10fF
C52786 OR2X1_LOC_689/a_8_216# OR2X1_LOC_585/A 0.01fF
C52787 AND2X1_LOC_59/Y OR2X1_LOC_831/a_8_216# 0.01fF
C52788 OR2X1_LOC_756/B OR2X1_LOC_435/Y 0.01fF
C52789 AND2X1_LOC_303/A OR2X1_LOC_316/Y -0.00fF
C52790 AND2X1_LOC_654/Y OR2X1_LOC_52/B 0.08fF
C52791 OR2X1_LOC_751/Y OR2X1_LOC_3/Y 0.01fF
C52792 OR2X1_LOC_31/Y AND2X1_LOC_476/Y 0.11fF
C52793 AND2X1_LOC_40/Y AND2X1_LOC_481/a_36_24# 0.01fF
C52794 D_INPUT_0 INPUT_2 0.06fF
C52795 OR2X1_LOC_151/A OR2X1_LOC_436/Y 0.03fF
C52796 OR2X1_LOC_680/Y OR2X1_LOC_144/Y 0.01fF
C52797 AND2X1_LOC_785/a_8_24# OR2X1_LOC_406/A 0.04fF
C52798 OR2X1_LOC_160/A OR2X1_LOC_87/B 0.03fF
C52799 OR2X1_LOC_185/A OR2X1_LOC_76/Y 0.02fF
C52800 OR2X1_LOC_87/A AND2X1_LOC_695/a_8_24# 0.04fF
C52801 OR2X1_LOC_131/A AND2X1_LOC_227/Y 0.04fF
C52802 AND2X1_LOC_340/a_8_24# OR2X1_LOC_71/Y 0.03fF
C52803 OR2X1_LOC_419/Y AND2X1_LOC_242/B 0.58fF
C52804 AND2X1_LOC_12/Y OR2X1_LOC_631/B 0.03fF
C52805 OR2X1_LOC_18/Y AND2X1_LOC_853/Y 0.01fF
C52806 OR2X1_LOC_87/A AND2X1_LOC_129/a_8_24# 0.01fF
C52807 OR2X1_LOC_696/A OR2X1_LOC_588/a_8_216# 0.07fF
C52808 INPUT_5 OR2X1_LOC_44/a_36_216# 0.00fF
C52809 OR2X1_LOC_130/A OR2X1_LOC_358/B 0.05fF
C52810 AND2X1_LOC_580/A AND2X1_LOC_578/a_36_24# 0.00fF
C52811 AND2X1_LOC_59/Y OR2X1_LOC_214/a_8_216# 0.06fF
C52812 OR2X1_LOC_643/A OR2X1_LOC_659/a_36_216# 0.00fF
C52813 OR2X1_LOC_270/Y OR2X1_LOC_486/Y 0.03fF
C52814 AND2X1_LOC_228/Y OR2X1_LOC_26/Y 0.03fF
C52815 AND2X1_LOC_6/a_36_24# OR2X1_LOC_633/A 0.01fF
C52816 OR2X1_LOC_154/A OR2X1_LOC_643/A 0.07fF
C52817 OR2X1_LOC_759/A OR2X1_LOC_95/Y 0.02fF
C52818 OR2X1_LOC_235/a_8_216# OR2X1_LOC_235/Y -0.00fF
C52819 AND2X1_LOC_580/A AND2X1_LOC_580/B 0.47fF
C52820 AND2X1_LOC_339/B OR2X1_LOC_289/a_36_216# 0.00fF
C52821 AND2X1_LOC_7/B OR2X1_LOC_358/A 0.07fF
C52822 OR2X1_LOC_22/A OR2X1_LOC_26/a_36_216# 0.02fF
C52823 AND2X1_LOC_544/Y OR2X1_LOC_746/Y 0.03fF
C52824 OR2X1_LOC_154/A OR2X1_LOC_778/Y 0.26fF
C52825 AND2X1_LOC_824/B AND2X1_LOC_234/a_8_24# 0.06fF
C52826 OR2X1_LOC_87/B AND2X1_LOC_29/a_36_24# 0.00fF
C52827 AND2X1_LOC_191/B AND2X1_LOC_849/a_8_24# 0.04fF
C52828 INPUT_0 OR2X1_LOC_818/a_8_216# 0.01fF
C52829 OR2X1_LOC_864/A OR2X1_LOC_204/Y 0.03fF
C52830 OR2X1_LOC_18/Y OR2X1_LOC_17/Y 0.00fF
C52831 OR2X1_LOC_6/B AND2X1_LOC_837/a_8_24# 0.07fF
C52832 OR2X1_LOC_530/Y OR2X1_LOC_39/A 0.00fF
C52833 AND2X1_LOC_51/Y OR2X1_LOC_794/A 0.09fF
C52834 AND2X1_LOC_80/a_8_24# OR2X1_LOC_647/B 0.01fF
C52835 OR2X1_LOC_502/A OR2X1_LOC_19/B 0.11fF
C52836 AND2X1_LOC_598/a_8_24# OR2X1_LOC_585/A 0.01fF
C52837 VDD AND2X1_LOC_660/A 0.26fF
C52838 OR2X1_LOC_155/A OR2X1_LOC_593/a_8_216# 0.04fF
C52839 OR2X1_LOC_186/Y OR2X1_LOC_365/B 0.06fF
C52840 OR2X1_LOC_614/a_8_216# OR2X1_LOC_78/A 0.02fF
C52841 AND2X1_LOC_645/A OR2X1_LOC_44/Y 0.01fF
C52842 OR2X1_LOC_756/B AND2X1_LOC_431/a_8_24# 0.01fF
C52843 AND2X1_LOC_711/Y AND2X1_LOC_848/Y 0.18fF
C52844 AND2X1_LOC_113/a_8_24# OR2X1_LOC_22/Y 0.03fF
C52845 OR2X1_LOC_105/Y OR2X1_LOC_814/A 0.37fF
C52846 OR2X1_LOC_756/B AND2X1_LOC_283/a_36_24# 0.00fF
C52847 OR2X1_LOC_26/Y OR2X1_LOC_585/A 6.19fF
C52848 OR2X1_LOC_312/Y AND2X1_LOC_374/Y 0.01fF
C52849 AND2X1_LOC_610/a_8_24# OR2X1_LOC_612/B 0.01fF
C52850 AND2X1_LOC_22/Y OR2X1_LOC_68/B 0.68fF
C52851 OR2X1_LOC_532/Y OR2X1_LOC_703/Y 0.00fF
C52852 OR2X1_LOC_517/Y OR2X1_LOC_74/A 0.04fF
C52853 OR2X1_LOC_653/A OR2X1_LOC_653/a_8_216# 0.01fF
C52854 VDD AND2X1_LOC_646/a_8_24# 0.00fF
C52855 OR2X1_LOC_405/A AND2X1_LOC_680/a_8_24# 0.02fF
C52856 OR2X1_LOC_216/A OR2X1_LOC_532/B 0.29fF
C52857 OR2X1_LOC_6/B OR2X1_LOC_493/Y 0.10fF
C52858 VDD AND2X1_LOC_418/a_8_24# -0.00fF
C52859 AND2X1_LOC_198/a_8_24# OR2X1_LOC_31/Y 0.02fF
C52860 OR2X1_LOC_66/A AND2X1_LOC_237/a_8_24# 0.01fF
C52861 AND2X1_LOC_349/B OR2X1_LOC_585/A 0.10fF
C52862 OR2X1_LOC_65/B OR2X1_LOC_65/a_36_216# 0.03fF
C52863 AND2X1_LOC_612/B AND2X1_LOC_611/a_36_24# 0.00fF
C52864 OR2X1_LOC_441/a_8_216# AND2X1_LOC_811/Y 0.47fF
C52865 OR2X1_LOC_51/Y OR2X1_LOC_289/Y 0.02fF
C52866 AND2X1_LOC_259/Y OR2X1_LOC_261/Y 0.02fF
C52867 AND2X1_LOC_300/a_8_24# OR2X1_LOC_228/Y 0.00fF
C52868 AND2X1_LOC_85/a_8_24# AND2X1_LOC_86/B 0.01fF
C52869 OR2X1_LOC_47/Y OR2X1_LOC_234/Y 0.01fF
C52870 OR2X1_LOC_673/Y OR2X1_LOC_404/Y 0.00fF
C52871 OR2X1_LOC_417/Y AND2X1_LOC_453/a_36_24# 0.01fF
C52872 OR2X1_LOC_158/A AND2X1_LOC_563/Y 0.05fF
C52873 OR2X1_LOC_778/A OR2X1_LOC_778/Y 0.11fF
C52874 OR2X1_LOC_306/Y AND2X1_LOC_308/a_36_24# 0.00fF
C52875 OR2X1_LOC_193/A OR2X1_LOC_269/B 0.09fF
C52876 OR2X1_LOC_506/B OR2X1_LOC_721/Y 0.03fF
C52877 OR2X1_LOC_240/a_8_216# D_INPUT_0 0.02fF
C52878 D_INPUT_0 OR2X1_LOC_739/A 0.04fF
C52879 OR2X1_LOC_743/A OR2X1_LOC_74/A -0.01fF
C52880 AND2X1_LOC_390/B OR2X1_LOC_485/A 0.07fF
C52881 INPUT_3 AND2X1_LOC_28/a_8_24# 0.01fF
C52882 OR2X1_LOC_74/Y OR2X1_LOC_75/Y 0.08fF
C52883 OR2X1_LOC_426/B AND2X1_LOC_647/Y 0.05fF
C52884 AND2X1_LOC_307/a_8_24# OR2X1_LOC_52/B 0.03fF
C52885 OR2X1_LOC_33/B OR2X1_LOC_33/a_8_216# 0.05fF
C52886 OR2X1_LOC_154/A OR2X1_LOC_113/A 0.03fF
C52887 OR2X1_LOC_31/Y OR2X1_LOC_595/a_8_216# 0.01fF
C52888 OR2X1_LOC_3/Y OR2X1_LOC_275/A 0.05fF
C52889 OR2X1_LOC_47/Y OR2X1_LOC_59/a_8_216# 0.14fF
C52890 AND2X1_LOC_711/Y OR2X1_LOC_617/Y 0.03fF
C52891 AND2X1_LOC_477/A OR2X1_LOC_44/Y 0.07fF
C52892 OR2X1_LOC_364/A OR2X1_LOC_602/B 0.03fF
C52893 AND2X1_LOC_703/a_8_24# OR2X1_LOC_47/Y 0.01fF
C52894 OR2X1_LOC_517/A AND2X1_LOC_845/a_8_24# 0.01fF
C52895 OR2X1_LOC_813/A OR2X1_LOC_85/A 0.47fF
C52896 OR2X1_LOC_485/A OR2X1_LOC_431/Y 0.05fF
C52897 OR2X1_LOC_802/Y OR2X1_LOC_532/B 0.01fF
C52898 AND2X1_LOC_634/Y OR2X1_LOC_26/Y 0.01fF
C52899 OR2X1_LOC_51/Y OR2X1_LOC_534/a_8_216# 0.02fF
C52900 AND2X1_LOC_17/Y AND2X1_LOC_425/Y 0.01fF
C52901 AND2X1_LOC_785/Y OR2X1_LOC_142/Y 0.03fF
C52902 OR2X1_LOC_468/Y OR2X1_LOC_532/B 0.02fF
C52903 OR2X1_LOC_87/A OR2X1_LOC_780/A 0.00fF
C52904 OR2X1_LOC_656/B OR2X1_LOC_340/a_8_216# 0.02fF
C52905 AND2X1_LOC_199/a_8_24# OR2X1_LOC_43/A 0.01fF
C52906 D_INPUT_0 OR2X1_LOC_269/B 0.45fF
C52907 AND2X1_LOC_31/Y OR2X1_LOC_78/A 2.41fF
C52908 OR2X1_LOC_506/B OR2X1_LOC_375/A 0.01fF
C52909 OR2X1_LOC_92/Y OR2X1_LOC_86/A 0.07fF
C52910 AND2X1_LOC_560/B AND2X1_LOC_656/Y 0.03fF
C52911 OR2X1_LOC_528/Y OR2X1_LOC_437/A 0.06fF
C52912 AND2X1_LOC_465/a_8_24# AND2X1_LOC_465/Y 0.00fF
C52913 AND2X1_LOC_47/Y OR2X1_LOC_781/a_8_216# 0.06fF
C52914 OR2X1_LOC_403/a_8_216# AND2X1_LOC_79/Y 0.01fF
C52915 OR2X1_LOC_246/A OR2X1_LOC_74/A 0.13fF
C52916 OR2X1_LOC_287/B INPUT_1 0.14fF
C52917 OR2X1_LOC_624/B AND2X1_LOC_79/a_8_24# 0.01fF
C52918 OR2X1_LOC_256/A OR2X1_LOC_248/Y 0.09fF
C52919 OR2X1_LOC_574/A AND2X1_LOC_69/a_8_24# 0.32fF
C52920 OR2X1_LOC_255/a_8_216# OR2X1_LOC_7/A 0.01fF
C52921 OR2X1_LOC_403/B AND2X1_LOC_47/Y 0.01fF
C52922 OR2X1_LOC_130/A OR2X1_LOC_112/B 0.04fF
C52923 AND2X1_LOC_722/a_36_24# OR2X1_LOC_437/A 0.00fF
C52924 OR2X1_LOC_43/A OR2X1_LOC_689/Y 0.01fF
C52925 OR2X1_LOC_458/B AND2X1_LOC_31/Y 0.11fF
C52926 AND2X1_LOC_810/Y AND2X1_LOC_653/a_36_24# 0.01fF
C52927 AND2X1_LOC_81/B AND2X1_LOC_88/Y 0.00fF
C52928 OR2X1_LOC_857/B AND2X1_LOC_36/Y 0.03fF
C52929 AND2X1_LOC_537/Y OR2X1_LOC_304/Y 0.00fF
C52930 OR2X1_LOC_87/A OR2X1_LOC_227/Y -0.01fF
C52931 AND2X1_LOC_40/Y OR2X1_LOC_641/B 0.03fF
C52932 OR2X1_LOC_8/Y OR2X1_LOC_13/B 0.01fF
C52933 OR2X1_LOC_88/Y AND2X1_LOC_266/a_8_24# 0.00fF
C52934 OR2X1_LOC_448/B AND2X1_LOC_31/Y 0.03fF
C52935 OR2X1_LOC_66/A OR2X1_LOC_777/B 0.06fF
C52936 AND2X1_LOC_514/Y AND2X1_LOC_863/A 0.02fF
C52937 OR2X1_LOC_87/A D_INPUT_1 0.04fF
C52938 OR2X1_LOC_264/Y OR2X1_LOC_560/A 0.64fF
C52939 AND2X1_LOC_18/a_36_24# AND2X1_LOC_7/Y 0.00fF
C52940 AND2X1_LOC_48/A OR2X1_LOC_19/B 0.37fF
C52941 AND2X1_LOC_18/Y OR2X1_LOC_539/B 0.13fF
C52942 OR2X1_LOC_825/Y INPUT_1 0.22fF
C52943 OR2X1_LOC_591/Y OR2X1_LOC_696/A 0.02fF
C52944 OR2X1_LOC_89/A AND2X1_LOC_645/a_8_24# 0.01fF
C52945 OR2X1_LOC_579/B OR2X1_LOC_493/Y 0.10fF
C52946 OR2X1_LOC_687/Y OR2X1_LOC_451/B 0.04fF
C52947 AND2X1_LOC_255/a_8_24# OR2X1_LOC_121/A 0.01fF
C52948 VDD OR2X1_LOC_577/B 0.10fF
C52949 OR2X1_LOC_377/A OR2X1_LOC_377/a_8_216# 0.06fF
C52950 OR2X1_LOC_703/a_8_216# OR2X1_LOC_356/A 0.02fF
C52951 OR2X1_LOC_429/Y OR2X1_LOC_51/B 0.02fF
C52952 OR2X1_LOC_176/a_8_216# AND2X1_LOC_212/Y 0.01fF
C52953 AND2X1_LOC_134/a_8_24# OR2X1_LOC_532/B 0.01fF
C52954 AND2X1_LOC_826/a_8_24# OR2X1_LOC_46/A 0.01fF
C52955 OR2X1_LOC_602/A AND2X1_LOC_31/Y 0.01fF
C52956 AND2X1_LOC_3/Y OR2X1_LOC_66/a_8_216# 0.07fF
C52957 OR2X1_LOC_291/a_8_216# OR2X1_LOC_71/A 0.01fF
C52958 OR2X1_LOC_574/A OR2X1_LOC_804/A 0.10fF
C52959 AND2X1_LOC_719/Y AND2X1_LOC_241/a_8_24# 0.25fF
C52960 OR2X1_LOC_696/A OR2X1_LOC_125/a_36_216# 0.00fF
C52961 OR2X1_LOC_808/B OR2X1_LOC_544/B 0.03fF
C52962 AND2X1_LOC_153/a_8_24# OR2X1_LOC_68/B 0.02fF
C52963 OR2X1_LOC_471/Y OR2X1_LOC_532/B 0.03fF
C52964 OR2X1_LOC_45/B AND2X1_LOC_714/B 0.07fF
C52965 AND2X1_LOC_76/Y OR2X1_LOC_13/B 0.03fF
C52966 OR2X1_LOC_335/A AND2X1_LOC_70/Y 0.03fF
C52967 OR2X1_LOC_53/Y AND2X1_LOC_200/a_8_24# 0.01fF
C52968 OR2X1_LOC_51/Y AND2X1_LOC_783/B 0.03fF
C52969 OR2X1_LOC_278/A OR2X1_LOC_47/Y 0.29fF
C52970 OR2X1_LOC_49/A OR2X1_LOC_158/A 2.63fF
C52971 OR2X1_LOC_643/A OR2X1_LOC_560/A 0.03fF
C52972 VDD OR2X1_LOC_56/Y 0.33fF
C52973 AND2X1_LOC_464/A AND2X1_LOC_476/Y 0.05fF
C52974 OR2X1_LOC_124/Y OR2X1_LOC_560/A 0.00fF
C52975 AND2X1_LOC_707/Y OR2X1_LOC_604/A 0.01fF
C52976 AND2X1_LOC_31/Y OR2X1_LOC_155/A 3.29fF
C52977 AND2X1_LOC_244/A AND2X1_LOC_243/Y 0.14fF
C52978 D_INPUT_5 INPUT_6 0.06fF
C52979 OR2X1_LOC_516/A OR2X1_LOC_437/A 0.12fF
C52980 OR2X1_LOC_323/A OR2X1_LOC_329/B 0.03fF
C52981 OR2X1_LOC_625/Y OR2X1_LOC_248/A 0.01fF
C52982 OR2X1_LOC_67/A OR2X1_LOC_13/B 0.03fF
C52983 AND2X1_LOC_342/Y OR2X1_LOC_437/A 0.08fF
C52984 OR2X1_LOC_175/Y AND2X1_LOC_92/Y 0.10fF
C52985 AND2X1_LOC_663/B AND2X1_LOC_848/A 0.00fF
C52986 OR2X1_LOC_487/Y AND2X1_LOC_657/A 0.03fF
C52987 AND2X1_LOC_712/Y OR2X1_LOC_158/A 0.02fF
C52988 OR2X1_LOC_476/Y OR2X1_LOC_228/Y 0.01fF
C52989 OR2X1_LOC_224/Y OR2X1_LOC_95/Y 0.00fF
C52990 OR2X1_LOC_344/A OR2X1_LOC_66/A 0.03fF
C52991 OR2X1_LOC_186/Y OR2X1_LOC_468/A 0.00fF
C52992 AND2X1_LOC_42/B OR2X1_LOC_80/A 0.32fF
C52993 OR2X1_LOC_405/A OR2X1_LOC_776/A 0.07fF
C52994 AND2X1_LOC_182/a_8_24# OR2X1_LOC_309/Y 0.01fF
C52995 OR2X1_LOC_78/A OR2X1_LOC_708/a_36_216# 0.00fF
C52996 AND2X1_LOC_352/a_36_24# AND2X1_LOC_566/B 0.00fF
C52997 OR2X1_LOC_246/A AND2X1_LOC_647/Y 0.12fF
C52998 AND2X1_LOC_12/Y INPUT_6 0.03fF
C52999 AND2X1_LOC_70/a_36_24# AND2X1_LOC_44/Y 0.00fF
C53000 OR2X1_LOC_160/B OR2X1_LOC_151/A 0.07fF
C53001 AND2X1_LOC_208/B OR2X1_LOC_56/Y 0.01fF
C53002 OR2X1_LOC_52/B OR2X1_LOC_13/B 0.23fF
C53003 AND2X1_LOC_463/B OR2X1_LOC_408/Y 0.01fF
C53004 OR2X1_LOC_756/B OR2X1_LOC_577/Y 0.14fF
C53005 OR2X1_LOC_456/A OR2X1_LOC_344/a_8_216# 0.46fF
C53006 AND2X1_LOC_92/Y OR2X1_LOC_713/A 0.02fF
C53007 OR2X1_LOC_703/B OR2X1_LOC_180/B 0.07fF
C53008 OR2X1_LOC_687/Y AND2X1_LOC_36/Y 0.03fF
C53009 OR2X1_LOC_95/Y OR2X1_LOC_597/Y 0.01fF
C53010 AND2X1_LOC_706/Y OR2X1_LOC_744/A 0.01fF
C53011 OR2X1_LOC_269/B OR2X1_LOC_339/A 0.01fF
C53012 OR2X1_LOC_40/Y OR2X1_LOC_813/a_36_216# 0.03fF
C53013 AND2X1_LOC_47/Y OR2X1_LOC_493/Y 0.10fF
C53014 AND2X1_LOC_91/B OR2X1_LOC_620/Y 0.07fF
C53015 AND2X1_LOC_628/a_8_24# OR2X1_LOC_549/A 0.02fF
C53016 OR2X1_LOC_87/A OR2X1_LOC_180/B 0.55fF
C53017 OR2X1_LOC_178/a_8_216# OR2X1_LOC_600/A 0.01fF
C53018 OR2X1_LOC_7/A AND2X1_LOC_449/a_8_24# 0.04fF
C53019 VDD OR2X1_LOC_676/Y 0.67fF
C53020 OR2X1_LOC_290/Y AND2X1_LOC_219/A 0.01fF
C53021 OR2X1_LOC_269/Y AND2X1_LOC_271/a_8_24# 0.23fF
C53022 AND2X1_LOC_95/Y OR2X1_LOC_174/a_8_216# 0.01fF
C53023 OR2X1_LOC_666/A AND2X1_LOC_244/a_8_24# 0.01fF
C53024 AND2X1_LOC_121/a_8_24# AND2X1_LOC_243/Y 0.04fF
C53025 OR2X1_LOC_158/A OR2X1_LOC_310/Y 0.08fF
C53026 OR2X1_LOC_600/A AND2X1_LOC_436/Y 0.03fF
C53027 AND2X1_LOC_216/Y OR2X1_LOC_59/Y 0.02fF
C53028 OR2X1_LOC_494/Y AND2X1_LOC_363/Y 0.08fF
C53029 INPUT_5 OR2X1_LOC_36/a_8_216# 0.01fF
C53030 OR2X1_LOC_71/Y AND2X1_LOC_562/Y 0.17fF
C53031 AND2X1_LOC_142/a_36_24# AND2X1_LOC_44/Y 0.00fF
C53032 VDD OR2X1_LOC_600/Y 0.12fF
C53033 OR2X1_LOC_254/B OR2X1_LOC_556/a_8_216# 0.01fF
C53034 OR2X1_LOC_7/A OR2X1_LOC_183/a_8_216# 0.21fF
C53035 OR2X1_LOC_18/Y AND2X1_LOC_473/Y 0.84fF
C53036 OR2X1_LOC_532/B OR2X1_LOC_750/Y 0.26fF
C53037 OR2X1_LOC_375/A AND2X1_LOC_258/a_8_24# 0.06fF
C53038 OR2X1_LOC_860/a_8_216# OR2X1_LOC_576/A 0.01fF
C53039 AND2X1_LOC_620/Y AND2X1_LOC_792/Y 0.07fF
C53040 AND2X1_LOC_534/a_8_24# OR2X1_LOC_502/A -0.01fF
C53041 OR2X1_LOC_18/Y AND2X1_LOC_287/B 0.00fF
C53042 OR2X1_LOC_696/A OR2X1_LOC_670/a_36_216# 0.00fF
C53043 OR2X1_LOC_175/Y AND2X1_LOC_166/a_8_24# 0.04fF
C53044 OR2X1_LOC_160/A OR2X1_LOC_392/B 0.03fF
C53045 OR2X1_LOC_78/B AND2X1_LOC_18/Y 0.65fF
C53046 AND2X1_LOC_646/a_8_24# OR2X1_LOC_67/Y 0.01fF
C53047 AND2X1_LOC_585/a_36_24# OR2X1_LOC_637/B 0.00fF
C53048 VDD OR2X1_LOC_834/A 0.21fF
C53049 AND2X1_LOC_570/Y OR2X1_LOC_51/Y 0.02fF
C53050 OR2X1_LOC_166/a_8_216# AND2X1_LOC_436/Y 0.47fF
C53051 OR2X1_LOC_18/Y OR2X1_LOC_816/A 0.03fF
C53052 OR2X1_LOC_331/A OR2X1_LOC_51/Y 0.01fF
C53053 AND2X1_LOC_91/B OR2X1_LOC_154/A 0.43fF
C53054 OR2X1_LOC_49/A OR2X1_LOC_847/A 0.03fF
C53055 OR2X1_LOC_208/A OR2X1_LOC_269/B 0.01fF
C53056 AND2X1_LOC_172/a_36_24# OR2X1_LOC_648/A 0.01fF
C53057 OR2X1_LOC_54/Y OR2X1_LOC_437/A 0.01fF
C53058 OR2X1_LOC_40/Y OR2X1_LOC_164/Y 0.00fF
C53059 OR2X1_LOC_109/Y OR2X1_LOC_323/a_36_216# 0.00fF
C53060 AND2X1_LOC_729/Y OR2X1_LOC_428/A 0.07fF
C53061 OR2X1_LOC_158/A OR2X1_LOC_422/Y 0.21fF
C53062 AND2X1_LOC_583/a_8_24# AND2X1_LOC_70/Y 0.01fF
C53063 AND2X1_LOC_594/a_8_24# AND2X1_LOC_95/Y 0.02fF
C53064 OR2X1_LOC_382/Y VDD 0.23fF
C53065 OR2X1_LOC_114/Y OR2X1_LOC_267/Y 0.02fF
C53066 AND2X1_LOC_110/Y OR2X1_LOC_502/A 0.07fF
C53067 OR2X1_LOC_531/Y AND2X1_LOC_549/a_8_24# 0.23fF
C53068 AND2X1_LOC_789/a_36_24# OR2X1_LOC_6/B 0.01fF
C53069 OR2X1_LOC_519/a_8_216# OR2X1_LOC_158/A 0.01fF
C53070 AND2X1_LOC_18/Y OR2X1_LOC_721/Y 0.02fF
C53071 OR2X1_LOC_638/B OR2X1_LOC_637/Y 0.17fF
C53072 AND2X1_LOC_564/B OR2X1_LOC_26/Y 0.01fF
C53073 OR2X1_LOC_447/A OR2X1_LOC_596/A 0.00fF
C53074 OR2X1_LOC_598/A OR2X1_LOC_493/Y 0.10fF
C53075 AND2X1_LOC_545/a_8_24# AND2X1_LOC_659/a_8_24# 0.23fF
C53076 OR2X1_LOC_427/A OR2X1_LOC_583/a_8_216# 0.03fF
C53077 OR2X1_LOC_374/Y OR2X1_LOC_717/a_8_216# 0.02fF
C53078 AND2X1_LOC_785/A OR2X1_LOC_527/Y 0.10fF
C53079 OR2X1_LOC_158/A OR2X1_LOC_433/Y 0.03fF
C53080 AND2X1_LOC_703/Y OR2X1_LOC_44/Y 0.01fF
C53081 OR2X1_LOC_105/Y OR2X1_LOC_244/Y 0.00fF
C53082 OR2X1_LOC_272/Y OR2X1_LOC_767/Y 0.01fF
C53083 AND2X1_LOC_784/A OR2X1_LOC_428/A 0.07fF
C53084 OR2X1_LOC_575/A OR2X1_LOC_66/A 0.03fF
C53085 AND2X1_LOC_42/B OR2X1_LOC_115/B 0.01fF
C53086 AND2X1_LOC_564/B OR2X1_LOC_89/A 0.07fF
C53087 OR2X1_LOC_528/a_36_216# AND2X1_LOC_573/A 0.00fF
C53088 OR2X1_LOC_133/a_8_216# OR2X1_LOC_85/A 0.05fF
C53089 OR2X1_LOC_134/Y AND2X1_LOC_276/Y 0.06fF
C53090 OR2X1_LOC_136/a_8_216# OR2X1_LOC_3/Y 0.04fF
C53091 AND2X1_LOC_168/Y AND2X1_LOC_568/B 0.02fF
C53092 VDD OR2X1_LOC_531/a_8_216# 0.21fF
C53093 OR2X1_LOC_223/A OR2X1_LOC_181/A 0.01fF
C53094 OR2X1_LOC_629/A OR2X1_LOC_563/A 0.08fF
C53095 AND2X1_LOC_716/Y AND2X1_LOC_514/a_8_24# 0.01fF
C53096 AND2X1_LOC_554/a_8_24# OR2X1_LOC_490/Y 0.03fF
C53097 AND2X1_LOC_706/a_8_24# OR2X1_LOC_36/Y 0.01fF
C53098 OR2X1_LOC_634/A OR2X1_LOC_634/a_8_216# 0.01fF
C53099 OR2X1_LOC_661/a_8_216# VDD 0.00fF
C53100 OR2X1_LOC_152/Y AND2X1_LOC_726/a_8_24# 0.25fF
C53101 AND2X1_LOC_540/a_36_24# OR2X1_LOC_744/A 0.01fF
C53102 OR2X1_LOC_186/Y OR2X1_LOC_449/B 0.03fF
C53103 AND2X1_LOC_712/a_8_24# OR2X1_LOC_7/A 0.05fF
C53104 OR2X1_LOC_599/A AND2X1_LOC_771/B 0.00fF
C53105 OR2X1_LOC_691/Y OR2X1_LOC_789/a_36_216# 0.00fF
C53106 OR2X1_LOC_185/A OR2X1_LOC_370/a_8_216# 0.15fF
C53107 OR2X1_LOC_589/A OR2X1_LOC_36/Y 0.52fF
C53108 OR2X1_LOC_851/a_8_216# OR2X1_LOC_185/A 0.01fF
C53109 OR2X1_LOC_203/Y AND2X1_LOC_275/a_8_24# 0.04fF
C53110 AND2X1_LOC_12/Y OR2X1_LOC_858/a_8_216# 0.03fF
C53111 OR2X1_LOC_619/Y AND2X1_LOC_436/Y 0.03fF
C53112 AND2X1_LOC_719/Y AND2X1_LOC_464/a_36_24# 0.06fF
C53113 AND2X1_LOC_99/A OR2X1_LOC_56/A 0.02fF
C53114 OR2X1_LOC_375/A AND2X1_LOC_18/Y 1.64fF
C53115 AND2X1_LOC_649/B AND2X1_LOC_219/Y 0.01fF
C53116 OR2X1_LOC_652/a_8_216# OR2X1_LOC_66/A 0.01fF
C53117 OR2X1_LOC_831/A OR2X1_LOC_269/B 0.03fF
C53118 AND2X1_LOC_824/a_8_24# OR2X1_LOC_66/A 0.03fF
C53119 OR2X1_LOC_490/a_8_216# OR2X1_LOC_7/A 0.06fF
C53120 OR2X1_LOC_404/Y OR2X1_LOC_720/Y 0.01fF
C53121 AND2X1_LOC_512/Y OR2X1_LOC_761/Y 0.01fF
C53122 OR2X1_LOC_6/B OR2X1_LOC_205/a_8_216# 0.03fF
C53123 AND2X1_LOC_12/Y OR2X1_LOC_648/A 0.07fF
C53124 AND2X1_LOC_56/B OR2X1_LOC_461/B 0.01fF
C53125 VDD OR2X1_LOC_462/B 0.45fF
C53126 OR2X1_LOC_216/A OR2X1_LOC_734/a_8_216# 0.03fF
C53127 VDD OR2X1_LOC_483/a_8_216# 0.00fF
C53128 AND2X1_LOC_570/Y OR2X1_LOC_680/A 0.03fF
C53129 OR2X1_LOC_158/A AND2X1_LOC_259/Y 0.01fF
C53130 OR2X1_LOC_486/B AND2X1_LOC_44/Y 0.16fF
C53131 OR2X1_LOC_778/Y OR2X1_LOC_723/a_8_216# 0.29fF
C53132 OR2X1_LOC_331/A OR2X1_LOC_680/A 0.06fF
C53133 OR2X1_LOC_585/A AND2X1_LOC_194/Y 0.84fF
C53134 OR2X1_LOC_160/A OR2X1_LOC_147/A 0.05fF
C53135 OR2X1_LOC_666/A AND2X1_LOC_286/Y 0.00fF
C53136 OR2X1_LOC_49/A AND2X1_LOC_46/a_8_24# 0.01fF
C53137 OR2X1_LOC_624/B OR2X1_LOC_113/B 0.89fF
C53138 AND2X1_LOC_99/Y OR2X1_LOC_278/Y 0.01fF
C53139 AND2X1_LOC_59/Y AND2X1_LOC_41/A 0.54fF
C53140 OR2X1_LOC_291/Y AND2X1_LOC_219/A 0.02fF
C53141 AND2X1_LOC_50/Y AND2X1_LOC_59/a_8_24# 0.01fF
C53142 AND2X1_LOC_319/A OR2X1_LOC_91/A 0.03fF
C53143 AND2X1_LOC_508/A AND2X1_LOC_807/Y 0.03fF
C53144 OR2X1_LOC_705/B OR2X1_LOC_550/B 0.05fF
C53145 AND2X1_LOC_535/Y AND2X1_LOC_336/a_36_24# -0.00fF
C53146 OR2X1_LOC_844/B D_INPUT_1 0.03fF
C53147 OR2X1_LOC_627/a_8_216# OR2X1_LOC_56/A 0.03fF
C53148 OR2X1_LOC_186/Y OR2X1_LOC_121/B 0.27fF
C53149 AND2X1_LOC_40/Y OR2X1_LOC_739/A 0.03fF
C53150 AND2X1_LOC_757/a_36_24# OR2X1_LOC_161/A 0.00fF
C53151 OR2X1_LOC_417/Y AND2X1_LOC_515/a_8_24# 0.23fF
C53152 OR2X1_LOC_864/A OR2X1_LOC_78/A 0.03fF
C53153 AND2X1_LOC_639/A OR2X1_LOC_428/A 0.19fF
C53154 AND2X1_LOC_95/Y OR2X1_LOC_792/Y 0.01fF
C53155 OR2X1_LOC_45/B AND2X1_LOC_477/A 0.07fF
C53156 OR2X1_LOC_152/Y OR2X1_LOC_679/a_8_216# 0.03fF
C53157 OR2X1_LOC_45/Y OR2X1_LOC_48/B 0.17fF
C53158 AND2X1_LOC_36/Y OR2X1_LOC_644/A 0.05fF
C53159 VDD OR2X1_LOC_487/Y 0.12fF
C53160 AND2X1_LOC_95/Y OR2X1_LOC_668/a_8_216# 0.01fF
C53161 AND2X1_LOC_804/Y AND2X1_LOC_808/a_36_24# 0.01fF
C53162 AND2X1_LOC_338/A OR2X1_LOC_46/A 0.01fF
C53163 OR2X1_LOC_92/Y AND2X1_LOC_655/A 0.02fF
C53164 AND2X1_LOC_566/Y OR2X1_LOC_51/Y 0.02fF
C53165 OR2X1_LOC_287/B OR2X1_LOC_287/A 0.01fF
C53166 OR2X1_LOC_45/Y OR2X1_LOC_18/Y 0.23fF
C53167 OR2X1_LOC_280/Y OR2X1_LOC_666/A 0.02fF
C53168 AND2X1_LOC_40/Y OR2X1_LOC_798/a_8_216# 0.04fF
C53169 AND2X1_LOC_94/Y AND2X1_LOC_42/a_8_24# 0.01fF
C53170 OR2X1_LOC_633/B OR2X1_LOC_78/A 0.05fF
C53171 AND2X1_LOC_583/a_8_24# AND2X1_LOC_17/Y 0.01fF
C53172 OR2X1_LOC_31/Y AND2X1_LOC_636/a_8_24# 0.01fF
C53173 OR2X1_LOC_833/B OR2X1_LOC_161/A 0.04fF
C53174 OR2X1_LOC_189/a_8_216# AND2X1_LOC_580/A 0.01fF
C53175 OR2X1_LOC_744/A OR2X1_LOC_485/A 0.56fF
C53176 OR2X1_LOC_36/Y AND2X1_LOC_654/B 0.02fF
C53177 AND2X1_LOC_857/Y OR2X1_LOC_26/Y 0.03fF
C53178 OR2X1_LOC_314/Y OR2X1_LOC_427/A 0.01fF
C53179 OR2X1_LOC_115/a_8_216# OR2X1_LOC_116/A -0.00fF
C53180 OR2X1_LOC_154/A AND2X1_LOC_39/a_36_24# 0.01fF
C53181 AND2X1_LOC_756/a_8_24# AND2X1_LOC_711/Y 0.03fF
C53182 OR2X1_LOC_18/Y AND2X1_LOC_807/Y 0.32fF
C53183 OR2X1_LOC_265/a_8_216# AND2X1_LOC_361/A 0.04fF
C53184 OR2X1_LOC_527/Y AND2X1_LOC_658/A 0.07fF
C53185 AND2X1_LOC_578/A AND2X1_LOC_663/A 0.10fF
C53186 AND2X1_LOC_40/Y OR2X1_LOC_269/B 2.37fF
C53187 VDD AND2X1_LOC_307/Y 0.04fF
C53188 OR2X1_LOC_703/B AND2X1_LOC_95/Y 0.03fF
C53189 OR2X1_LOC_824/Y AND2X1_LOC_852/B 0.02fF
C53190 AND2X1_LOC_839/B AND2X1_LOC_839/a_8_24# 0.19fF
C53191 AND2X1_LOC_59/Y OR2X1_LOC_662/A 0.03fF
C53192 AND2X1_LOC_347/Y OR2X1_LOC_89/A 0.94fF
C53193 OR2X1_LOC_40/Y AND2X1_LOC_633/Y 0.02fF
C53194 AND2X1_LOC_527/a_8_24# AND2X1_LOC_56/B 0.01fF
C53195 AND2X1_LOC_572/A OR2X1_LOC_118/Y 0.00fF
C53196 AND2X1_LOC_729/B AND2X1_LOC_434/Y 0.01fF
C53197 AND2X1_LOC_706/Y OR2X1_LOC_31/Y 0.11fF
C53198 AND2X1_LOC_339/B AND2X1_LOC_831/Y 0.01fF
C53199 AND2X1_LOC_540/a_8_24# OR2X1_LOC_7/A 0.01fF
C53200 AND2X1_LOC_736/a_8_24# AND2X1_LOC_711/Y 0.07fF
C53201 AND2X1_LOC_95/Y OR2X1_LOC_87/A 0.18fF
C53202 AND2X1_LOC_343/a_36_24# OR2X1_LOC_517/A 0.00fF
C53203 OR2X1_LOC_6/B AND2X1_LOC_5/a_8_24# 0.02fF
C53204 OR2X1_LOC_810/a_8_216# OR2X1_LOC_269/B 0.01fF
C53205 AND2X1_LOC_182/A OR2X1_LOC_417/A 0.08fF
C53206 AND2X1_LOC_314/a_36_24# AND2X1_LOC_56/B 0.00fF
C53207 OR2X1_LOC_40/Y D_INPUT_0 0.13fF
C53208 AND2X1_LOC_361/a_8_24# OR2X1_LOC_95/Y 0.01fF
C53209 OR2X1_LOC_591/a_8_216# OR2X1_LOC_48/B 0.02fF
C53210 AND2X1_LOC_620/Y OR2X1_LOC_816/A 0.01fF
C53211 OR2X1_LOC_3/Y OR2X1_LOC_16/a_8_216# 0.01fF
C53212 AND2X1_LOC_535/Y AND2X1_LOC_801/B 0.00fF
C53213 OR2X1_LOC_840/A AND2X1_LOC_42/B 0.00fF
C53214 OR2X1_LOC_157/a_8_216# INPUT_4 0.01fF
C53215 OR2X1_LOC_700/Y OR2X1_LOC_748/A 0.01fF
C53216 OR2X1_LOC_666/A OR2X1_LOC_22/Y 0.03fF
C53217 OR2X1_LOC_426/B OR2X1_LOC_263/a_8_216# 0.31fF
C53218 AND2X1_LOC_155/a_8_24# OR2X1_LOC_743/A 0.05fF
C53219 AND2X1_LOC_61/Y AND2X1_LOC_640/a_8_24# 0.02fF
C53220 AND2X1_LOC_719/Y AND2X1_LOC_849/a_36_24# 0.08fF
C53221 OR2X1_LOC_537/A OR2X1_LOC_269/B 0.00fF
C53222 OR2X1_LOC_787/Y OR2X1_LOC_794/A 0.44fF
C53223 OR2X1_LOC_90/a_8_216# OR2X1_LOC_46/A 0.03fF
C53224 AND2X1_LOC_59/Y OR2X1_LOC_631/B 0.02fF
C53225 AND2X1_LOC_392/A OR2X1_LOC_111/Y 0.03fF
C53226 AND2X1_LOC_580/A AND2X1_LOC_565/Y 0.01fF
C53227 OR2X1_LOC_58/Y OR2X1_LOC_31/Y 0.01fF
C53228 OR2X1_LOC_858/A OR2X1_LOC_814/A 0.08fF
C53229 AND2X1_LOC_679/a_8_24# AND2X1_LOC_7/B 0.01fF
C53230 AND2X1_LOC_688/a_8_24# OR2X1_LOC_39/A 0.03fF
C53231 OR2X1_LOC_117/Y OR2X1_LOC_67/a_8_216# 0.01fF
C53232 AND2X1_LOC_342/Y OR2X1_LOC_753/A 0.01fF
C53233 OR2X1_LOC_687/Y OR2X1_LOC_687/B 0.01fF
C53234 OR2X1_LOC_622/a_36_216# OR2X1_LOC_847/A 0.00fF
C53235 OR2X1_LOC_809/B OR2X1_LOC_532/B 0.24fF
C53236 AND2X1_LOC_22/Y AND2X1_LOC_497/a_36_24# 0.01fF
C53237 OR2X1_LOC_848/A OR2X1_LOC_269/B 0.01fF
C53238 AND2X1_LOC_711/A AND2X1_LOC_866/A 0.10fF
C53239 OR2X1_LOC_43/A OR2X1_LOC_36/Y 0.29fF
C53240 OR2X1_LOC_3/Y OR2X1_LOC_118/Y 0.07fF
C53241 OR2X1_LOC_87/A OR2X1_LOC_99/Y 0.03fF
C53242 OR2X1_LOC_859/B OR2X1_LOC_269/B 0.01fF
C53243 VDD OR2X1_LOC_200/Y 0.00fF
C53244 AND2X1_LOC_140/a_8_24# AND2X1_LOC_573/A 0.01fF
C53245 AND2X1_LOC_721/Y AND2X1_LOC_563/Y 0.02fF
C53246 AND2X1_LOC_597/a_8_24# OR2X1_LOC_155/A 0.04fF
C53247 AND2X1_LOC_210/a_8_24# OR2X1_LOC_163/Y 0.00fF
C53248 AND2X1_LOC_12/Y AND2X1_LOC_136/a_8_24# 0.01fF
C53249 OR2X1_LOC_246/a_8_216# OR2X1_LOC_585/A 0.01fF
C53250 AND2X1_LOC_576/Y OR2X1_LOC_239/a_8_216# 0.01fF
C53251 AND2X1_LOC_716/Y OR2X1_LOC_22/Y 0.07fF
C53252 OR2X1_LOC_227/B OR2X1_LOC_68/B 0.37fF
C53253 AND2X1_LOC_170/B OR2X1_LOC_91/A 0.00fF
C53254 OR2X1_LOC_485/A AND2X1_LOC_840/B 0.12fF
C53255 AND2X1_LOC_456/Y OR2X1_LOC_497/Y 0.03fF
C53256 AND2X1_LOC_853/Y OR2X1_LOC_585/A 0.03fF
C53257 AND2X1_LOC_319/a_8_24# OR2X1_LOC_56/A 0.04fF
C53258 AND2X1_LOC_36/Y OR2X1_LOC_199/B 0.11fF
C53259 AND2X1_LOC_727/A OR2X1_LOC_48/B 0.07fF
C53260 OR2X1_LOC_423/a_8_216# AND2X1_LOC_454/A 0.10fF
C53261 OR2X1_LOC_22/Y AND2X1_LOC_654/Y 0.26fF
C53262 AND2X1_LOC_84/a_8_24# OR2X1_LOC_585/A 0.01fF
C53263 OR2X1_LOC_428/A OR2X1_LOC_172/Y 0.06fF
C53264 AND2X1_LOC_44/Y OR2X1_LOC_348/B 0.03fF
C53265 OR2X1_LOC_223/A OR2X1_LOC_742/a_36_216# 0.00fF
C53266 OR2X1_LOC_275/a_8_216# AND2X1_LOC_139/B 0.01fF
C53267 OR2X1_LOC_88/Y OR2X1_LOC_595/A 0.09fF
C53268 AND2X1_LOC_356/B OR2X1_LOC_312/Y 0.03fF
C53269 AND2X1_LOC_690/a_8_24# D_INPUT_0 0.01fF
C53270 OR2X1_LOC_837/Y AND2X1_LOC_472/a_8_24# 0.03fF
C53271 OR2X1_LOC_3/Y OR2X1_LOC_262/Y 0.45fF
C53272 OR2X1_LOC_280/Y OR2X1_LOC_312/Y 0.04fF
C53273 AND2X1_LOC_658/A AND2X1_LOC_483/Y 0.03fF
C53274 AND2X1_LOC_139/A AND2X1_LOC_141/A 0.83fF
C53275 AND2X1_LOC_81/B OR2X1_LOC_121/B 0.05fF
C53276 AND2X1_LOC_43/B OR2X1_LOC_46/A 12.07fF
C53277 AND2X1_LOC_502/a_8_24# OR2X1_LOC_22/Y 0.02fF
C53278 AND2X1_LOC_46/a_8_24# OR2X1_LOC_87/B 0.19fF
C53279 AND2X1_LOC_810/Y OR2X1_LOC_594/Y 0.25fF
C53280 INPUT_3 INPUT_1 1.06fF
C53281 AND2X1_LOC_59/Y OR2X1_LOC_403/a_8_216# 0.14fF
C53282 OR2X1_LOC_864/a_8_216# OR2X1_LOC_557/A 0.00fF
C53283 AND2X1_LOC_391/Y AND2X1_LOC_721/A 0.03fF
C53284 AND2X1_LOC_155/Y OR2X1_LOC_7/A 0.01fF
C53285 OR2X1_LOC_595/A AND2X1_LOC_772/a_36_24# 0.01fF
C53286 OR2X1_LOC_62/B OR2X1_LOC_39/A 0.03fF
C53287 OR2X1_LOC_91/A AND2X1_LOC_721/A 0.03fF
C53288 OR2X1_LOC_485/A OR2X1_LOC_282/a_8_216# 0.07fF
C53289 OR2X1_LOC_95/Y OR2X1_LOC_48/B 0.03fF
C53290 OR2X1_LOC_230/a_8_216# OR2X1_LOC_7/A 0.05fF
C53291 AND2X1_LOC_8/Y OR2X1_LOC_99/B 0.04fF
C53292 OR2X1_LOC_160/A OR2X1_LOC_532/B 0.98fF
C53293 AND2X1_LOC_774/a_8_24# OR2X1_LOC_13/B 0.03fF
C53294 OR2X1_LOC_18/Y OR2X1_LOC_95/Y 4.92fF
C53295 OR2X1_LOC_54/Y OR2X1_LOC_753/A 0.00fF
C53296 OR2X1_LOC_18/Y OR2X1_LOC_368/A 0.52fF
C53297 OR2X1_LOC_618/a_8_216# D_INPUT_0 0.01fF
C53298 AND2X1_LOC_662/B AND2X1_LOC_476/A 0.00fF
C53299 OR2X1_LOC_22/A OR2X1_LOC_588/Y 0.02fF
C53300 OR2X1_LOC_529/Y AND2X1_LOC_842/B 0.02fF
C53301 OR2X1_LOC_109/Y AND2X1_LOC_851/B 0.01fF
C53302 OR2X1_LOC_70/A OR2X1_LOC_26/a_8_216# 0.08fF
C53303 OR2X1_LOC_13/a_8_216# OR2X1_LOC_13/B 0.01fF
C53304 AND2X1_LOC_652/a_36_24# AND2X1_LOC_810/Y 0.00fF
C53305 OR2X1_LOC_92/Y OR2X1_LOC_599/Y 0.18fF
C53306 OR2X1_LOC_19/B AND2X1_LOC_3/Y 0.32fF
C53307 OR2X1_LOC_696/A AND2X1_LOC_227/a_8_24# 0.01fF
C53308 OR2X1_LOC_312/Y OR2X1_LOC_22/Y 0.06fF
C53309 OR2X1_LOC_335/A OR2X1_LOC_718/a_8_216# 0.01fF
C53310 OR2X1_LOC_865/B D_INPUT_1 0.03fF
C53311 OR2X1_LOC_475/Y OR2X1_LOC_215/A 0.14fF
C53312 OR2X1_LOC_574/A OR2X1_LOC_62/B 0.00fF
C53313 AND2X1_LOC_22/Y OR2X1_LOC_598/a_8_216# 0.03fF
C53314 D_INPUT_0 AND2X1_LOC_857/a_8_24# 0.02fF
C53315 OR2X1_LOC_495/Y OR2X1_LOC_419/Y 0.05fF
C53316 OR2X1_LOC_811/A OR2X1_LOC_241/B 0.07fF
C53317 OR2X1_LOC_78/B OR2X1_LOC_789/A 0.03fF
C53318 AND2X1_LOC_734/Y AND2X1_LOC_222/Y 0.18fF
C53319 OR2X1_LOC_47/Y AND2X1_LOC_848/Y 0.03fF
C53320 D_INPUT_0 OR2X1_LOC_7/A 0.05fF
C53321 AND2X1_LOC_250/a_8_24# OR2X1_LOC_579/B 0.04fF
C53322 AND2X1_LOC_244/a_8_24# OR2X1_LOC_13/B 0.04fF
C53323 AND2X1_LOC_477/Y OR2X1_LOC_142/Y 0.07fF
C53324 AND2X1_LOC_86/B OR2X1_LOC_532/B 0.03fF
C53325 OR2X1_LOC_66/A OR2X1_LOC_735/B 0.08fF
C53326 OR2X1_LOC_506/A OR2X1_LOC_493/Y 0.02fF
C53327 OR2X1_LOC_563/A OR2X1_LOC_562/A 0.02fF
C53328 OR2X1_LOC_385/Y OR2X1_LOC_95/Y 0.51fF
C53329 AND2X1_LOC_476/A AND2X1_LOC_634/a_8_24# 0.02fF
C53330 OR2X1_LOC_485/A OR2X1_LOC_31/Y 1.58fF
C53331 OR2X1_LOC_624/B OR2X1_LOC_532/B 0.59fF
C53332 OR2X1_LOC_66/A OR2X1_LOC_332/a_8_216# 0.01fF
C53333 AND2X1_LOC_22/Y OR2X1_LOC_174/a_8_216# 0.02fF
C53334 AND2X1_LOC_30/a_8_24# OR2X1_LOC_51/B 0.00fF
C53335 OR2X1_LOC_472/B OR2X1_LOC_416/Y 0.01fF
C53336 VDD OR2X1_LOC_749/Y 0.08fF
C53337 OR2X1_LOC_151/A OR2X1_LOC_354/a_8_216# 0.03fF
C53338 OR2X1_LOC_622/A AND2X1_LOC_36/Y 0.28fF
C53339 OR2X1_LOC_45/B OR2X1_LOC_406/Y 0.06fF
C53340 AND2X1_LOC_64/Y OR2X1_LOC_294/Y 0.00fF
C53341 D_INPUT_3 AND2X1_LOC_37/a_8_24# 0.01fF
C53342 OR2X1_LOC_680/A OR2X1_LOC_406/A 0.07fF
C53343 OR2X1_LOC_427/A AND2X1_LOC_657/A 0.14fF
C53344 AND2X1_LOC_291/a_8_24# OR2X1_LOC_598/A 0.02fF
C53345 AND2X1_LOC_672/B OR2X1_LOC_62/B 0.42fF
C53346 AND2X1_LOC_91/B OR2X1_LOC_435/A 0.01fF
C53347 OR2X1_LOC_696/A AND2X1_LOC_541/Y 0.11fF
C53348 OR2X1_LOC_263/a_8_216# OR2X1_LOC_246/A 0.05fF
C53349 OR2X1_LOC_143/a_8_216# INPUT_2 0.00fF
C53350 OR2X1_LOC_177/Y AND2X1_LOC_543/Y 0.00fF
C53351 OR2X1_LOC_538/A OR2X1_LOC_112/A 0.03fF
C53352 OR2X1_LOC_669/Y AND2X1_LOC_721/A 0.06fF
C53353 OR2X1_LOC_273/Y AND2X1_LOC_476/A 0.03fF
C53354 OR2X1_LOC_43/A OR2X1_LOC_419/Y 0.01fF
C53355 OR2X1_LOC_19/B OR2X1_LOC_607/a_8_216# 0.03fF
C53356 OR2X1_LOC_835/a_8_216# OR2X1_LOC_598/A 0.14fF
C53357 AND2X1_LOC_445/a_8_24# AND2X1_LOC_455/B 0.01fF
C53358 OR2X1_LOC_118/Y AND2X1_LOC_772/a_8_24# 0.00fF
C53359 OR2X1_LOC_205/a_8_216# OR2X1_LOC_598/A 0.02fF
C53360 OR2X1_LOC_86/Y AND2X1_LOC_647/Y 0.02fF
C53361 OR2X1_LOC_412/a_8_216# INPUT_1 0.02fF
C53362 OR2X1_LOC_709/A OR2X1_LOC_139/A 0.00fF
C53363 AND2X1_LOC_594/a_8_24# AND2X1_LOC_22/Y 0.02fF
C53364 OR2X1_LOC_335/B AND2X1_LOC_309/a_36_24# 0.00fF
C53365 AND2X1_LOC_122/a_8_24# OR2X1_LOC_786/Y 0.06fF
C53366 AND2X1_LOC_64/Y OR2X1_LOC_641/A 0.03fF
C53367 OR2X1_LOC_486/Y AND2X1_LOC_7/B 0.03fF
C53368 AND2X1_LOC_340/Y OR2X1_LOC_79/Y 0.14fF
C53369 AND2X1_LOC_573/A AND2X1_LOC_217/a_8_24# 0.01fF
C53370 AND2X1_LOC_87/a_8_24# OR2X1_LOC_72/Y 0.01fF
C53371 OR2X1_LOC_198/a_8_216# OR2X1_LOC_66/A 0.04fF
C53372 OR2X1_LOC_620/Y OR2X1_LOC_446/B 0.07fF
C53373 AND2X1_LOC_539/Y OR2X1_LOC_40/Y 0.03fF
C53374 OR2X1_LOC_12/Y OR2X1_LOC_16/A 0.67fF
C53375 AND2X1_LOC_65/A AND2X1_LOC_44/Y 0.65fF
C53376 OR2X1_LOC_78/A OR2X1_LOC_714/a_36_216# 0.01fF
C53377 AND2X1_LOC_53/Y AND2X1_LOC_7/Y 0.08fF
C53378 OR2X1_LOC_696/A OR2X1_LOC_107/a_8_216# 0.01fF
C53379 AND2X1_LOC_571/A AND2X1_LOC_561/B 0.24fF
C53380 AND2X1_LOC_817/a_8_24# OR2X1_LOC_68/B 0.01fF
C53381 AND2X1_LOC_177/a_8_24# OR2X1_LOC_180/B 0.01fF
C53382 AND2X1_LOC_31/Y OR2X1_LOC_68/a_8_216# 0.03fF
C53383 AND2X1_LOC_195/a_8_24# OR2X1_LOC_13/Y 0.01fF
C53384 OR2X1_LOC_154/A OR2X1_LOC_446/B 0.08fF
C53385 OR2X1_LOC_40/Y AND2X1_LOC_350/B 0.03fF
C53386 OR2X1_LOC_851/A AND2X1_LOC_36/Y 0.10fF
C53387 OR2X1_LOC_177/Y OR2X1_LOC_322/Y 0.02fF
C53388 OR2X1_LOC_830/a_8_216# AND2X1_LOC_44/Y 0.01fF
C53389 OR2X1_LOC_421/A AND2X1_LOC_774/A 0.00fF
C53390 OR2X1_LOC_40/Y AND2X1_LOC_364/a_36_24# 0.00fF
C53391 OR2X1_LOC_439/a_8_216# OR2X1_LOC_440/A 0.01fF
C53392 OR2X1_LOC_113/B OR2X1_LOC_768/a_8_216# 0.49fF
C53393 OR2X1_LOC_671/Y OR2X1_LOC_158/A 0.11fF
C53394 OR2X1_LOC_158/A AND2X1_LOC_714/B 0.03fF
C53395 OR2X1_LOC_45/B OR2X1_LOC_496/a_8_216# 0.01fF
C53396 OR2X1_LOC_139/A AND2X1_LOC_70/Y 0.08fF
C53397 AND2X1_LOC_64/Y AND2X1_LOC_312/a_8_24# 0.03fF
C53398 OR2X1_LOC_8/Y OR2X1_LOC_428/A 0.07fF
C53399 AND2X1_LOC_555/Y OR2X1_LOC_292/Y 0.01fF
C53400 OR2X1_LOC_220/B AND2X1_LOC_36/Y 0.03fF
C53401 OR2X1_LOC_637/A AND2X1_LOC_763/B 0.00fF
C53402 OR2X1_LOC_213/A OR2X1_LOC_550/B 0.04fF
C53403 OR2X1_LOC_274/a_8_216# OR2X1_LOC_120/a_8_216# 0.47fF
C53404 AND2X1_LOC_802/B OR2X1_LOC_744/A 0.05fF
C53405 OR2X1_LOC_66/A OR2X1_LOC_161/B 0.32fF
C53406 OR2X1_LOC_44/Y OR2X1_LOC_589/a_8_216# 0.02fF
C53407 OR2X1_LOC_703/B OR2X1_LOC_788/B 0.85fF
C53408 AND2X1_LOC_286/Y OR2X1_LOC_13/B 0.00fF
C53409 OR2X1_LOC_539/Y OR2X1_LOC_339/A 0.73fF
C53410 AND2X1_LOC_95/Y OR2X1_LOC_844/B 0.01fF
C53411 OR2X1_LOC_3/Y OR2X1_LOC_39/a_8_216# 0.09fF
C53412 AND2X1_LOC_476/A OR2X1_LOC_75/Y 0.03fF
C53413 OR2X1_LOC_821/Y OR2X1_LOC_822/Y 0.21fF
C53414 OR2X1_LOC_190/A OR2X1_LOC_344/A 0.07fF
C53415 AND2X1_LOC_18/Y OR2X1_LOC_549/A 0.15fF
C53416 OR2X1_LOC_26/Y OR2X1_LOC_437/A 0.43fF
C53417 OR2X1_LOC_732/B OR2X1_LOC_308/Y 0.04fF
C53418 OR2X1_LOC_87/A AND2X1_LOC_41/Y 0.03fF
C53419 OR2X1_LOC_506/A OR2X1_LOC_130/a_8_216# 0.01fF
C53420 AND2X1_LOC_276/Y OR2X1_LOC_521/a_8_216# 0.13fF
C53421 OR2X1_LOC_95/Y AND2X1_LOC_620/Y 0.02fF
C53422 AND2X1_LOC_493/a_8_24# OR2X1_LOC_437/A 0.01fF
C53423 OR2X1_LOC_40/Y AND2X1_LOC_784/a_8_24# 0.02fF
C53424 OR2X1_LOC_673/Y OR2X1_LOC_771/B 0.07fF
C53425 OR2X1_LOC_528/Y AND2X1_LOC_547/Y 0.00fF
C53426 OR2X1_LOC_708/Y OR2X1_LOC_779/A 0.01fF
C53427 AND2X1_LOC_311/a_8_24# OR2X1_LOC_161/B 0.01fF
C53428 OR2X1_LOC_696/A OR2X1_LOC_529/a_8_216# 0.03fF
C53429 AND2X1_LOC_349/B OR2X1_LOC_437/A 0.02fF
C53430 OR2X1_LOC_89/A OR2X1_LOC_437/A 0.22fF
C53431 AND2X1_LOC_95/Y OR2X1_LOC_390/B 0.07fF
C53432 OR2X1_LOC_52/B OR2X1_LOC_142/a_8_216# 0.06fF
C53433 OR2X1_LOC_835/B AND2X1_LOC_36/Y 0.07fF
C53434 OR2X1_LOC_770/B OR2X1_LOC_78/Y -0.00fF
C53435 AND2X1_LOC_356/B OR2X1_LOC_13/B 0.01fF
C53436 OR2X1_LOC_337/A OR2X1_LOC_335/Y 0.14fF
C53437 OR2X1_LOC_532/B OR2X1_LOC_717/a_8_216# 0.01fF
C53438 OR2X1_LOC_40/Y AND2X1_LOC_711/A 0.01fF
C53439 OR2X1_LOC_112/a_8_216# OR2X1_LOC_78/B 0.01fF
C53440 OR2X1_LOC_40/Y AND2X1_LOC_326/B 0.00fF
C53441 OR2X1_LOC_280/Y OR2X1_LOC_13/B 0.00fF
C53442 OR2X1_LOC_379/Y AND2X1_LOC_64/Y 0.03fF
C53443 AND2X1_LOC_64/a_8_24# AND2X1_LOC_36/Y 0.20fF
C53444 OR2X1_LOC_442/Y AND2X1_LOC_477/Y 0.04fF
C53445 OR2X1_LOC_188/Y OR2X1_LOC_811/A 0.03fF
C53446 OR2X1_LOC_186/Y OR2X1_LOC_317/a_8_216# 0.01fF
C53447 AND2X1_LOC_31/Y OR2X1_LOC_814/A 0.77fF
C53448 OR2X1_LOC_122/a_36_216# AND2X1_LOC_362/B 0.00fF
C53449 OR2X1_LOC_450/A OR2X1_LOC_450/B 0.12fF
C53450 AND2X1_LOC_22/Y OR2X1_LOC_668/a_8_216# 0.07fF
C53451 OR2X1_LOC_304/a_36_216# OR2X1_LOC_45/Y 0.01fF
C53452 OR2X1_LOC_337/A AND2X1_LOC_40/Y 0.02fF
C53453 OR2X1_LOC_411/A OR2X1_LOC_51/Y 0.01fF
C53454 OR2X1_LOC_158/A AND2X1_LOC_861/B 0.09fF
C53455 OR2X1_LOC_6/B OR2X1_LOC_78/a_8_216# 0.01fF
C53456 OR2X1_LOC_628/a_36_216# OR2X1_LOC_816/A 0.00fF
C53457 AND2X1_LOC_84/Y OR2X1_LOC_39/A 0.03fF
C53458 AND2X1_LOC_723/Y AND2X1_LOC_180/a_8_24# 0.19fF
C53459 AND2X1_LOC_728/Y AND2X1_LOC_220/B 0.03fF
C53460 AND2X1_LOC_76/Y OR2X1_LOC_428/A 0.02fF
C53461 OR2X1_LOC_40/Y AND2X1_LOC_471/Y 0.02fF
C53462 OR2X1_LOC_177/Y AND2X1_LOC_544/a_8_24# 0.01fF
C53463 OR2X1_LOC_604/A OR2X1_LOC_297/A 0.04fF
C53464 AND2X1_LOC_91/B AND2X1_LOC_395/a_8_24# 0.04fF
C53465 OR2X1_LOC_113/Y AND2X1_LOC_18/Y 0.01fF
C53466 OR2X1_LOC_130/A OR2X1_LOC_390/a_8_216# 0.02fF
C53467 D_INPUT_1 OR2X1_LOC_493/Y 0.18fF
C53468 AND2X1_LOC_237/a_8_24# OR2X1_LOC_241/B 0.01fF
C53469 OR2X1_LOC_185/Y OR2X1_LOC_115/B 0.05fF
C53470 OR2X1_LOC_186/Y OR2X1_LOC_856/B 0.02fF
C53471 AND2X1_LOC_390/a_8_24# AND2X1_LOC_512/Y 0.00fF
C53472 AND2X1_LOC_64/Y OR2X1_LOC_114/Y 0.04fF
C53473 OR2X1_LOC_858/A OR2X1_LOC_244/Y 0.03fF
C53474 AND2X1_LOC_76/Y OR2X1_LOC_595/A 0.00fF
C53475 OR2X1_LOC_710/A OR2X1_LOC_269/B 0.00fF
C53476 OR2X1_LOC_130/A OR2X1_LOC_855/A 0.00fF
C53477 OR2X1_LOC_393/Y OR2X1_LOC_16/A 0.03fF
C53478 OR2X1_LOC_178/Y OR2X1_LOC_59/Y 0.04fF
C53479 OR2X1_LOC_212/a_8_216# OR2X1_LOC_486/Y 0.03fF
C53480 AND2X1_LOC_203/Y AND2X1_LOC_205/a_8_24# 0.19fF
C53481 VDD AND2X1_LOC_820/B 0.19fF
C53482 AND2X1_LOC_715/Y AND2X1_LOC_354/B 0.09fF
C53483 OR2X1_LOC_22/Y OR2X1_LOC_13/B 0.77fF
C53484 OR2X1_LOC_168/B OR2X1_LOC_648/A 0.07fF
C53485 OR2X1_LOC_464/A OR2X1_LOC_733/A 0.09fF
C53486 OR2X1_LOC_435/B OR2X1_LOC_66/A 0.34fF
C53487 OR2X1_LOC_799/A OR2X1_LOC_435/A 0.31fF
C53488 OR2X1_LOC_185/A OR2X1_LOC_736/Y 0.03fF
C53489 OR2X1_LOC_604/A AND2X1_LOC_866/B 0.02fF
C53490 AND2X1_LOC_753/B AND2X1_LOC_41/a_8_24# 0.02fF
C53491 OR2X1_LOC_696/A OR2X1_LOC_824/a_8_216# 0.01fF
C53492 AND2X1_LOC_22/Y OR2X1_LOC_87/A 0.13fF
C53493 AND2X1_LOC_758/a_8_24# AND2X1_LOC_866/B 0.02fF
C53494 OR2X1_LOC_696/A AND2X1_LOC_390/B 0.18fF
C53495 AND2X1_LOC_361/a_36_24# OR2X1_LOC_427/A -0.02fF
C53496 OR2X1_LOC_427/A AND2X1_LOC_479/a_8_24# 0.01fF
C53497 OR2X1_LOC_692/Y AND2X1_LOC_655/A 0.81fF
C53498 OR2X1_LOC_739/A OR2X1_LOC_356/A 0.03fF
C53499 OR2X1_LOC_67/A OR2X1_LOC_595/A 0.03fF
C53500 OR2X1_LOC_604/A OR2X1_LOC_495/Y 0.25fF
C53501 AND2X1_LOC_588/B AND2X1_LOC_17/Y 0.69fF
C53502 OR2X1_LOC_175/Y OR2X1_LOC_389/B 0.02fF
C53503 OR2X1_LOC_40/Y AND2X1_LOC_840/A 0.01fF
C53504 AND2X1_LOC_539/Y OR2X1_LOC_7/A 0.03fF
C53505 OR2X1_LOC_539/a_8_216# OR2X1_LOC_390/A 0.01fF
C53506 AND2X1_LOC_555/Y AND2X1_LOC_345/a_8_24# 0.03fF
C53507 AND2X1_LOC_784/A AND2X1_LOC_794/a_36_24# 0.01fF
C53508 OR2X1_LOC_499/B AND2X1_LOC_628/a_8_24# 0.01fF
C53509 AND2X1_LOC_339/B AND2X1_LOC_139/B 0.01fF
C53510 OR2X1_LOC_604/A AND2X1_LOC_450/a_8_24# 0.01fF
C53511 OR2X1_LOC_329/B AND2X1_LOC_116/a_36_24# 0.00fF
C53512 OR2X1_LOC_306/Y OR2X1_LOC_589/A 0.03fF
C53513 OR2X1_LOC_49/A OR2X1_LOC_748/A 0.03fF
C53514 OR2X1_LOC_154/A OR2X1_LOC_863/A 0.06fF
C53515 VDD OR2X1_LOC_427/A 0.75fF
C53516 AND2X1_LOC_831/Y OR2X1_LOC_300/Y 0.02fF
C53517 AND2X1_LOC_64/Y OR2X1_LOC_201/Y 0.06fF
C53518 OR2X1_LOC_106/Y AND2X1_LOC_276/Y 0.02fF
C53519 AND2X1_LOC_366/a_36_24# OR2X1_LOC_92/Y 0.00fF
C53520 OR2X1_LOC_52/B OR2X1_LOC_428/A 0.37fF
C53521 OR2X1_LOC_493/a_8_216# OR2X1_LOC_737/A 0.01fF
C53522 OR2X1_LOC_672/Y OR2X1_LOC_428/A 0.01fF
C53523 AND2X1_LOC_74/a_8_24# OR2X1_LOC_787/B 0.08fF
C53524 OR2X1_LOC_532/B OR2X1_LOC_532/Y 0.01fF
C53525 OR2X1_LOC_375/A OR2X1_LOC_307/A 0.01fF
C53526 AND2X1_LOC_715/Y AND2X1_LOC_390/B 0.10fF
C53527 AND2X1_LOC_41/A AND2X1_LOC_67/a_36_24# 0.00fF
C53528 OR2X1_LOC_759/A AND2X1_LOC_621/Y 0.03fF
C53529 AND2X1_LOC_728/Y AND2X1_LOC_209/a_8_24# 0.01fF
C53530 OR2X1_LOC_467/B OR2X1_LOC_87/A 0.00fF
C53531 OR2X1_LOC_51/Y OR2X1_LOC_625/a_36_216# 0.00fF
C53532 VDD OR2X1_LOC_823/Y 0.12fF
C53533 AND2X1_LOC_489/Y OR2X1_LOC_428/A 0.02fF
C53534 OR2X1_LOC_52/B OR2X1_LOC_595/A 0.14fF
C53535 OR2X1_LOC_641/Y OR2X1_LOC_185/A 0.59fF
C53536 OR2X1_LOC_158/A OR2X1_LOC_42/a_8_216# 0.01fF
C53537 OR2X1_LOC_269/B OR2X1_LOC_356/A 0.88fF
C53538 OR2X1_LOC_808/B OR2X1_LOC_708/Y 0.31fF
C53539 AND2X1_LOC_41/A OR2X1_LOC_623/B 0.07fF
C53540 OR2X1_LOC_784/Y OR2X1_LOC_78/A 0.65fF
C53541 AND2X1_LOC_587/a_8_24# AND2X1_LOC_51/Y 0.20fF
C53542 D_INPUT_0 OR2X1_LOC_319/Y 0.21fF
C53543 OR2X1_LOC_87/a_8_216# OR2X1_LOC_66/A 0.22fF
C53544 OR2X1_LOC_713/a_8_216# OR2X1_LOC_779/A 0.47fF
C53545 AND2X1_LOC_489/Y OR2X1_LOC_595/A 0.07fF
C53546 AND2X1_LOC_43/B OR2X1_LOC_702/a_8_216# 0.01fF
C53547 AND2X1_LOC_787/a_8_24# AND2X1_LOC_477/a_8_24# 0.23fF
C53548 OR2X1_LOC_666/A OR2X1_LOC_39/A 0.17fF
C53549 INPUT_0 AND2X1_LOC_414/a_36_24# 0.00fF
C53550 OR2X1_LOC_7/A AND2X1_LOC_771/B 0.04fF
C53551 AND2X1_LOC_59/Y OR2X1_LOC_648/A 0.25fF
C53552 AND2X1_LOC_786/a_8_24# OR2X1_LOC_64/Y 0.01fF
C53553 OR2X1_LOC_272/Y OR2X1_LOC_16/A 0.00fF
C53554 AND2X1_LOC_100/a_8_24# AND2X1_LOC_243/Y 0.01fF
C53555 AND2X1_LOC_141/a_36_24# OR2X1_LOC_65/B 0.00fF
C53556 OR2X1_LOC_158/B AND2X1_LOC_213/B 0.83fF
C53557 OR2X1_LOC_604/A OR2X1_LOC_43/A 0.10fF
C53558 OR2X1_LOC_421/A OR2X1_LOC_433/a_36_216# 0.00fF
C53559 OR2X1_LOC_46/A AND2X1_LOC_416/a_8_24# 0.01fF
C53560 OR2X1_LOC_96/Y OR2X1_LOC_670/Y 0.01fF
C53561 OR2X1_LOC_43/A AND2X1_LOC_207/B 0.01fF
C53562 OR2X1_LOC_505/Y AND2X1_LOC_806/A 0.25fF
C53563 OR2X1_LOC_677/Y OR2X1_LOC_427/A 0.03fF
C53564 OR2X1_LOC_696/A AND2X1_LOC_863/Y 0.07fF
C53565 AND2X1_LOC_123/a_8_24# AND2X1_LOC_243/Y 0.03fF
C53566 AND2X1_LOC_12/Y OR2X1_LOC_573/a_36_216# 0.02fF
C53567 OR2X1_LOC_653/B OR2X1_LOC_435/Y 0.16fF
C53568 VDD AND2X1_LOC_363/A 0.21fF
C53569 OR2X1_LOC_777/B OR2X1_LOC_241/B 0.04fF
C53570 D_INPUT_4 AND2X1_LOC_11/Y 0.16fF
C53571 AND2X1_LOC_717/Y AND2X1_LOC_723/a_8_24# -0.01fF
C53572 AND2X1_LOC_658/A AND2X1_LOC_806/A 0.03fF
C53573 OR2X1_LOC_448/B OR2X1_LOC_784/Y 0.00fF
C53574 OR2X1_LOC_743/A AND2X1_LOC_448/a_8_24# 0.01fF
C53575 OR2X1_LOC_185/A OR2X1_LOC_808/B 0.03fF
C53576 OR2X1_LOC_64/Y OR2X1_LOC_766/a_36_216# 0.03fF
C53577 AND2X1_LOC_500/Y OR2X1_LOC_498/Y 0.14fF
C53578 OR2X1_LOC_45/B AND2X1_LOC_465/Y 0.02fF
C53579 OR2X1_LOC_252/a_8_216# AND2X1_LOC_866/B 0.18fF
C53580 OR2X1_LOC_434/A OR2X1_LOC_174/a_8_216# 0.50fF
C53581 AND2X1_LOC_832/a_8_24# OR2X1_LOC_48/B 0.03fF
C53582 OR2X1_LOC_61/A AND2X1_LOC_48/A 0.01fF
C53583 AND2X1_LOC_504/a_36_24# OR2X1_LOC_502/A 0.00fF
C53584 AND2X1_LOC_572/a_8_24# OR2X1_LOC_71/Y 0.01fF
C53585 OR2X1_LOC_791/B OR2X1_LOC_850/B 0.16fF
C53586 OR2X1_LOC_599/A AND2X1_LOC_148/a_8_24# 0.01fF
C53587 AND2X1_LOC_170/Y OR2X1_LOC_91/A 0.02fF
C53588 OR2X1_LOC_468/A OR2X1_LOC_574/A 0.03fF
C53589 OR2X1_LOC_244/B OR2X1_LOC_87/A 0.03fF
C53590 AND2X1_LOC_64/Y OR2X1_LOC_201/a_8_216# 0.00fF
C53591 AND2X1_LOC_727/A AND2X1_LOC_810/B 0.00fF
C53592 OR2X1_LOC_64/Y OR2X1_LOC_421/Y 0.10fF
C53593 OR2X1_LOC_323/A AND2X1_LOC_476/A 0.05fF
C53594 OR2X1_LOC_91/A AND2X1_LOC_361/A 0.07fF
C53595 OR2X1_LOC_405/A AND2X1_LOC_492/a_8_24# 0.01fF
C53596 OR2X1_LOC_377/A OR2X1_LOC_403/A 0.05fF
C53597 AND2X1_LOC_40/Y OR2X1_LOC_539/Y 0.00fF
C53598 INPUT_0 AND2X1_LOC_472/B 0.07fF
C53599 AND2X1_LOC_653/B OR2X1_LOC_594/Y 0.10fF
C53600 AND2X1_LOC_191/B OR2X1_LOC_757/a_36_216# 0.00fF
C53601 AND2X1_LOC_40/Y AND2X1_LOC_617/a_36_24# 0.00fF
C53602 OR2X1_LOC_530/Y OR2X1_LOC_51/Y 0.31fF
C53603 OR2X1_LOC_364/A OR2X1_LOC_840/A 0.10fF
C53604 AND2X1_LOC_168/Y AND2X1_LOC_170/a_8_24# 0.09fF
C53605 OR2X1_LOC_393/a_8_216# OR2X1_LOC_39/A 0.05fF
C53606 OR2X1_LOC_286/Y OR2X1_LOC_288/a_8_216# 0.39fF
C53607 AND2X1_LOC_456/B OR2X1_LOC_669/a_8_216# 0.01fF
C53608 AND2X1_LOC_554/B OR2X1_LOC_56/A 0.04fF
C53609 AND2X1_LOC_738/B OR2X1_LOC_680/Y -0.01fF
C53610 OR2X1_LOC_329/B OR2X1_LOC_238/Y 0.10fF
C53611 OR2X1_LOC_691/A D_INPUT_0 0.01fF
C53612 OR2X1_LOC_97/A AND2X1_LOC_47/Y 0.12fF
C53613 OR2X1_LOC_259/a_8_216# OR2X1_LOC_161/A 0.01fF
C53614 OR2X1_LOC_333/B AND2X1_LOC_92/Y 0.16fF
C53615 OR2X1_LOC_18/Y OR2X1_LOC_257/a_36_216# 0.03fF
C53616 AND2X1_LOC_53/Y OR2X1_LOC_706/a_8_216# 0.00fF
C53617 AND2X1_LOC_91/B AND2X1_LOC_813/a_8_24# 0.01fF
C53618 AND2X1_LOC_801/B OR2X1_LOC_16/A 0.03fF
C53619 OR2X1_LOC_472/A OR2X1_LOC_634/A 0.18fF
C53620 AND2X1_LOC_544/Y AND2X1_LOC_803/a_8_24# 0.07fF
C53621 AND2X1_LOC_849/A AND2X1_LOC_243/Y 0.09fF
C53622 OR2X1_LOC_720/B AND2X1_LOC_65/A 0.00fF
C53623 AND2X1_LOC_857/Y AND2X1_LOC_853/Y 0.13fF
C53624 OR2X1_LOC_625/Y AND2X1_LOC_848/Y 0.07fF
C53625 OR2X1_LOC_158/A AND2X1_LOC_477/A 0.03fF
C53626 OR2X1_LOC_235/B OR2X1_LOC_233/a_8_216# 0.02fF
C53627 OR2X1_LOC_258/Y OR2X1_LOC_59/Y 0.05fF
C53628 OR2X1_LOC_251/a_8_216# OR2X1_LOC_585/A 0.02fF
C53629 OR2X1_LOC_619/Y AND2X1_LOC_655/A 0.10fF
C53630 AND2X1_LOC_43/B OR2X1_LOC_739/A 0.02fF
C53631 AND2X1_LOC_753/a_36_24# AND2X1_LOC_43/B 0.01fF
C53632 OR2X1_LOC_190/A OR2X1_LOC_456/A 0.10fF
C53633 OR2X1_LOC_235/B AND2X1_LOC_38/a_8_24# 0.03fF
C53634 OR2X1_LOC_619/Y AND2X1_LOC_467/a_36_24# 0.00fF
C53635 OR2X1_LOC_416/A OR2X1_LOC_414/Y 0.00fF
C53636 AND2X1_LOC_675/Y AND2X1_LOC_578/A 0.12fF
C53637 OR2X1_LOC_620/Y AND2X1_LOC_56/B 0.04fF
C53638 OR2X1_LOC_493/B OR2X1_LOC_121/B 0.01fF
C53639 OR2X1_LOC_624/B OR2X1_LOC_624/Y 0.02fF
C53640 AND2X1_LOC_12/Y OR2X1_LOC_847/a_8_216# 0.01fF
C53641 AND2X1_LOC_326/A OR2X1_LOC_56/A 0.03fF
C53642 OR2X1_LOC_229/a_36_216# OR2X1_LOC_31/Y 0.00fF
C53643 OR2X1_LOC_544/A OR2X1_LOC_439/B 0.04fF
C53644 OR2X1_LOC_377/A OR2X1_LOC_130/A 0.01fF
C53645 OR2X1_LOC_831/B OR2X1_LOC_241/B 0.01fF
C53646 AND2X1_LOC_734/Y OR2X1_LOC_74/A 0.03fF
C53647 D_GATE_662 AND2X1_LOC_47/Y 0.01fF
C53648 AND2X1_LOC_716/Y AND2X1_LOC_211/B 0.00fF
C53649 VDD AND2X1_LOC_687/B 0.06fF
C53650 AND2X1_LOC_91/B OR2X1_LOC_330/a_36_216# 0.00fF
C53651 OR2X1_LOC_647/Y OR2X1_LOC_78/B 0.01fF
C53652 OR2X1_LOC_188/Y AND2X1_LOC_237/a_8_24# 0.01fF
C53653 OR2X1_LOC_188/a_8_216# OR2X1_LOC_241/B -0.03fF
C53654 OR2X1_LOC_99/B AND2X1_LOC_92/Y 0.61fF
C53655 AND2X1_LOC_181/Y OR2X1_LOC_95/Y 0.16fF
C53656 OR2X1_LOC_387/Y OR2X1_LOC_92/Y 0.01fF
C53657 OR2X1_LOC_65/B AND2X1_LOC_266/Y 0.04fF
C53658 AND2X1_LOC_120/a_8_24# AND2X1_LOC_850/A 0.03fF
C53659 OR2X1_LOC_251/Y OR2X1_LOC_427/A 0.06fF
C53660 OR2X1_LOC_11/Y OR2X1_LOC_95/a_8_216# 0.08fF
C53661 AND2X1_LOC_181/Y OR2X1_LOC_368/A 0.02fF
C53662 OR2X1_LOC_271/B OR2X1_LOC_316/Y 0.01fF
C53663 OR2X1_LOC_271/a_8_216# OR2X1_LOC_315/Y 0.02fF
C53664 AND2X1_LOC_847/Y OR2X1_LOC_701/a_8_216# 0.03fF
C53665 AND2X1_LOC_41/A AND2X1_LOC_13/a_36_24# 0.01fF
C53666 OR2X1_LOC_784/Y OR2X1_LOC_155/A 0.00fF
C53667 OR2X1_LOC_693/a_8_216# AND2X1_LOC_648/B 0.01fF
C53668 AND2X1_LOC_153/a_8_24# OR2X1_LOC_87/A 0.03fF
C53669 AND2X1_LOC_573/A AND2X1_LOC_361/A 0.02fF
C53670 OR2X1_LOC_200/a_8_216# AND2X1_LOC_43/B 0.03fF
C53671 OR2X1_LOC_685/A OR2X1_LOC_685/B 0.23fF
C53672 OR2X1_LOC_516/A AND2X1_LOC_784/A 0.02fF
C53673 INPUT_0 OR2X1_LOC_19/B 0.20fF
C53674 AND2X1_LOC_40/Y AND2X1_LOC_176/a_8_24# 0.04fF
C53675 AND2X1_LOC_43/B OR2X1_LOC_269/B 2.72fF
C53676 OR2X1_LOC_46/A AND2X1_LOC_219/Y 0.00fF
C53677 OR2X1_LOC_756/B AND2X1_LOC_442/a_8_24# 0.03fF
C53678 OR2X1_LOC_804/a_8_216# OR2X1_LOC_121/B 0.01fF
C53679 OR2X1_LOC_154/A AND2X1_LOC_56/B 0.49fF
C53680 OR2X1_LOC_306/Y OR2X1_LOC_43/A 0.09fF
C53681 OR2X1_LOC_154/A OR2X1_LOC_659/B 0.03fF
C53682 OR2X1_LOC_11/Y AND2X1_LOC_472/B 0.01fF
C53683 OR2X1_LOC_64/Y OR2X1_LOC_763/a_8_216# 0.01fF
C53684 AND2X1_LOC_154/a_8_24# OR2X1_LOC_52/B 0.02fF
C53685 OR2X1_LOC_424/Y AND2X1_LOC_449/a_8_24# 0.09fF
C53686 AND2X1_LOC_79/a_8_24# OR2X1_LOC_78/Y 0.00fF
C53687 OR2X1_LOC_401/a_36_216# OR2X1_LOC_78/Y 0.00fF
C53688 OR2X1_LOC_743/A OR2X1_LOC_432/Y 0.40fF
C53689 AND2X1_LOC_35/Y OR2X1_LOC_24/a_8_216# 0.01fF
C53690 AND2X1_LOC_33/Y OR2X1_LOC_24/Y 0.01fF
C53691 AND2X1_LOC_45/a_36_24# OR2X1_LOC_706/A 0.00fF
C53692 OR2X1_LOC_467/A OR2X1_LOC_780/a_8_216# 0.01fF
C53693 OR2X1_LOC_473/A OR2X1_LOC_631/A 0.83fF
C53694 OR2X1_LOC_664/Y AND2X1_LOC_3/Y 0.05fF
C53695 OR2X1_LOC_678/Y D_INPUT_0 0.61fF
C53696 OR2X1_LOC_706/B OR2X1_LOC_706/A 0.16fF
C53697 OR2X1_LOC_181/Y OR2X1_LOC_469/B 0.08fF
C53698 OR2X1_LOC_473/Y OR2X1_LOC_493/A 0.80fF
C53699 AND2X1_LOC_8/Y OR2X1_LOC_267/A 0.01fF
C53700 OR2X1_LOC_185/Y OR2X1_LOC_789/a_8_216# 0.03fF
C53701 AND2X1_LOC_216/A OR2X1_LOC_595/A 0.00fF
C53702 OR2X1_LOC_26/Y OR2X1_LOC_753/A 0.07fF
C53703 OR2X1_LOC_530/Y OR2X1_LOC_680/A 0.00fF
C53704 OR2X1_LOC_64/Y OR2X1_LOC_278/Y 0.10fF
C53705 OR2X1_LOC_313/a_8_216# OR2X1_LOC_70/Y 0.09fF
C53706 AND2X1_LOC_169/a_8_24# AND2X1_LOC_436/a_8_24# 0.23fF
C53707 AND2X1_LOC_169/a_36_24# AND2X1_LOC_434/Y 0.00fF
C53708 OR2X1_LOC_541/A AND2X1_LOC_47/Y 0.03fF
C53709 OR2X1_LOC_469/a_8_216# OR2X1_LOC_711/A 0.01fF
C53710 OR2X1_LOC_64/Y AND2X1_LOC_662/B 0.04fF
C53711 AND2X1_LOC_348/Y OR2X1_LOC_89/A 0.11fF
C53712 AND2X1_LOC_259/Y OR2X1_LOC_748/A 1.91fF
C53713 AND2X1_LOC_477/A OR2X1_LOC_594/Y 0.19fF
C53714 AND2X1_LOC_578/A OR2X1_LOC_189/A 0.01fF
C53715 OR2X1_LOC_3/Y AND2X1_LOC_349/a_8_24# 0.17fF
C53716 OR2X1_LOC_691/Y AND2X1_LOC_751/a_8_24# 0.01fF
C53717 OR2X1_LOC_574/A OR2X1_LOC_449/B 0.05fF
C53718 AND2X1_LOC_349/B OR2X1_LOC_753/A 0.02fF
C53719 OR2X1_LOC_89/A OR2X1_LOC_753/A 0.11fF
C53720 OR2X1_LOC_502/A AND2X1_LOC_7/Y 0.03fF
C53721 OR2X1_LOC_599/A AND2X1_LOC_148/Y 0.12fF
C53722 OR2X1_LOC_628/Y AND2X1_LOC_805/Y 0.03fF
C53723 OR2X1_LOC_51/Y OR2X1_LOC_51/B 0.07fF
C53724 OR2X1_LOC_400/a_8_216# OR2X1_LOC_532/B 0.01fF
C53725 AND2X1_LOC_211/B OR2X1_LOC_312/Y 0.07fF
C53726 AND2X1_LOC_651/B OR2X1_LOC_44/Y 0.00fF
C53727 AND2X1_LOC_56/B OR2X1_LOC_778/A 0.01fF
C53728 AND2X1_LOC_723/a_8_24# OR2X1_LOC_417/A 0.04fF
C53729 OR2X1_LOC_377/A OR2X1_LOC_62/B 0.06fF
C53730 OR2X1_LOC_485/A OR2X1_LOC_420/Y 0.01fF
C53731 OR2X1_LOC_47/Y OR2X1_LOC_394/a_8_216# 0.00fF
C53732 OR2X1_LOC_844/a_36_216# OR2X1_LOC_810/A 0.15fF
C53733 OR2X1_LOC_126/a_8_216# OR2X1_LOC_3/Y 0.01fF
C53734 OR2X1_LOC_847/A OR2X1_LOC_532/B 0.00fF
C53735 AND2X1_LOC_354/a_8_24# AND2X1_LOC_727/A 0.01fF
C53736 AND2X1_LOC_733/Y OR2X1_LOC_437/a_8_216# 0.01fF
C53737 OR2X1_LOC_417/A OR2X1_LOC_278/Y 0.04fF
C53738 OR2X1_LOC_447/A OR2X1_LOC_532/B 0.01fF
C53739 OR2X1_LOC_362/B OR2X1_LOC_286/B 0.00fF
C53740 AND2X1_LOC_72/B OR2X1_LOC_78/A 0.03fF
C53741 AND2X1_LOC_562/B OR2X1_LOC_47/Y 0.01fF
C53742 OR2X1_LOC_188/Y OR2X1_LOC_777/B 0.03fF
C53743 AND2X1_LOC_662/B OR2X1_LOC_417/A 0.07fF
C53744 AND2X1_LOC_477/A AND2X1_LOC_652/a_36_24# 0.01fF
C53745 OR2X1_LOC_780/A AND2X1_LOC_426/a_8_24# 0.17fF
C53746 OR2X1_LOC_472/B OR2X1_LOC_6/A 0.06fF
C53747 OR2X1_LOC_41/Y AND2X1_LOC_434/Y 0.01fF
C53748 AND2X1_LOC_660/A AND2X1_LOC_642/Y 0.15fF
C53749 AND2X1_LOC_728/Y OR2X1_LOC_679/A 0.01fF
C53750 OR2X1_LOC_448/Y OR2X1_LOC_447/Y 0.46fF
C53751 OR2X1_LOC_62/B OR2X1_LOC_85/A 0.15fF
C53752 AND2X1_LOC_707/Y AND2X1_LOC_449/a_8_24# 0.04fF
C53753 OR2X1_LOC_185/A OR2X1_LOC_218/Y 0.02fF
C53754 AND2X1_LOC_99/A D_INPUT_3 0.03fF
C53755 AND2X1_LOC_337/B OR2X1_LOC_64/Y 0.00fF
C53756 OR2X1_LOC_646/A OR2X1_LOC_647/a_8_216# 0.01fF
C53757 OR2X1_LOC_574/A OR2X1_LOC_121/B 0.49fF
C53758 OR2X1_LOC_864/A OR2X1_LOC_814/A 0.08fF
C53759 AND2X1_LOC_687/A OR2X1_LOC_7/A 0.03fF
C53760 AND2X1_LOC_7/B OR2X1_LOC_308/Y 0.09fF
C53761 AND2X1_LOC_22/Y OR2X1_LOC_844/B 0.00fF
C53762 OR2X1_LOC_464/A OR2X1_LOC_741/A 0.01fF
C53763 AND2X1_LOC_91/B OR2X1_LOC_605/Y 0.25fF
C53764 OR2X1_LOC_11/Y OR2X1_LOC_64/a_36_216# 0.00fF
C53765 D_INPUT_0 OR2X1_LOC_86/a_8_216# 0.07fF
C53766 OR2X1_LOC_26/Y AND2X1_LOC_845/Y 0.02fF
C53767 OR2X1_LOC_417/Y OR2X1_LOC_417/a_8_216# 0.01fF
C53768 OR2X1_LOC_59/Y AND2X1_LOC_216/a_8_24# 0.01fF
C53769 OR2X1_LOC_206/A OR2X1_LOC_201/Y 0.04fF
C53770 OR2X1_LOC_45/B OR2X1_LOC_516/Y 0.10fF
C53771 OR2X1_LOC_185/Y OR2X1_LOC_241/Y 0.13fF
C53772 OR2X1_LOC_202/a_36_216# AND2X1_LOC_51/Y 0.00fF
C53773 OR2X1_LOC_737/A OR2X1_LOC_493/Y 0.04fF
C53774 OR2X1_LOC_235/B OR2X1_LOC_68/B 0.13fF
C53775 OR2X1_LOC_485/Y OR2X1_LOC_13/B 0.35fF
C53776 AND2X1_LOC_22/Y OR2X1_LOC_390/B 0.07fF
C53777 OR2X1_LOC_377/A AND2X1_LOC_39/Y 0.00fF
C53778 OR2X1_LOC_89/A AND2X1_LOC_845/Y 0.09fF
C53779 OR2X1_LOC_63/a_8_216# OR2X1_LOC_67/Y 0.05fF
C53780 OR2X1_LOC_831/B AND2X1_LOC_273/a_36_24# 0.01fF
C53781 AND2X1_LOC_95/Y OR2X1_LOC_493/Y 0.03fF
C53782 OR2X1_LOC_95/Y OR2X1_LOC_585/A 1.71fF
C53783 VDD OR2X1_LOC_561/A 0.00fF
C53784 OR2X1_LOC_161/B OR2X1_LOC_354/a_36_216# 0.00fF
C53785 OR2X1_LOC_64/Y OR2X1_LOC_19/B 0.09fF
C53786 AND2X1_LOC_624/A AND2X1_LOC_793/Y 0.07fF
C53787 OR2X1_LOC_427/A OR2X1_LOC_163/Y 0.16fF
C53788 OR2X1_LOC_147/B AND2X1_LOC_31/Y 0.05fF
C53789 OR2X1_LOC_392/B OR2X1_LOC_474/B 0.16fF
C53790 OR2X1_LOC_375/A OR2X1_LOC_512/a_8_216# 0.01fF
C53791 OR2X1_LOC_267/Y OR2X1_LOC_572/a_8_216# 0.01fF
C53792 AND2X1_LOC_8/Y OR2X1_LOC_84/a_8_216# 0.02fF
C53793 OR2X1_LOC_64/Y AND2X1_LOC_800/a_8_24# 0.00fF
C53794 OR2X1_LOC_143/a_36_216# OR2X1_LOC_9/Y 0.00fF
C53795 AND2X1_LOC_517/a_8_24# AND2X1_LOC_31/Y 0.11fF
C53796 OR2X1_LOC_97/A OR2X1_LOC_34/A -0.00fF
C53797 OR2X1_LOC_816/A OR2X1_LOC_530/a_8_216# 0.01fF
C53798 AND2X1_LOC_707/Y AND2X1_LOC_712/a_8_24# -0.00fF
C53799 OR2X1_LOC_253/a_8_216# OR2X1_LOC_417/A 0.14fF
C53800 OR2X1_LOC_769/B OR2X1_LOC_771/B 0.02fF
C53801 OR2X1_LOC_617/Y AND2X1_LOC_663/a_8_24# 0.03fF
C53802 AND2X1_LOC_48/A AND2X1_LOC_7/Y 0.00fF
C53803 AND2X1_LOC_774/a_8_24# OR2X1_LOC_428/A 0.03fF
C53804 OR2X1_LOC_78/A AND2X1_LOC_36/Y 0.17fF
C53805 AND2X1_LOC_8/Y OR2X1_LOC_99/A 0.06fF
C53806 OR2X1_LOC_76/Y OR2X1_LOC_76/a_36_216# 0.00fF
C53807 OR2X1_LOC_201/a_8_216# OR2X1_LOC_206/A 0.01fF
C53808 OR2X1_LOC_155/A OR2X1_LOC_512/a_36_216# 0.01fF
C53809 OR2X1_LOC_113/a_8_216# OR2X1_LOC_113/B 0.03fF
C53810 OR2X1_LOC_637/B OR2X1_LOC_769/a_8_216# 0.01fF
C53811 OR2X1_LOC_474/B OR2X1_LOC_113/B 0.02fF
C53812 OR2X1_LOC_126/a_36_216# OR2X1_LOC_6/B 0.03fF
C53813 AND2X1_LOC_28/a_8_24# INPUT_1 0.09fF
C53814 OR2X1_LOC_294/Y OR2X1_LOC_342/A 0.01fF
C53815 OR2X1_LOC_281/Y OR2X1_LOC_428/A 0.33fF
C53816 OR2X1_LOC_566/A OR2X1_LOC_325/B 0.06fF
C53817 AND2X1_LOC_817/B OR2X1_LOC_80/A 0.46fF
C53818 AND2X1_LOC_828/a_8_24# AND2X1_LOC_774/A 0.20fF
C53819 OR2X1_LOC_709/A OR2X1_LOC_138/A 0.31fF
C53820 OR2X1_LOC_405/A OR2X1_LOC_317/B 0.03fF
C53821 OR2X1_LOC_62/A OR2X1_LOC_54/Y 0.17fF
C53822 AND2X1_LOC_56/B OR2X1_LOC_198/A 0.02fF
C53823 OR2X1_LOC_532/B AND2X1_LOC_108/a_8_24# 0.14fF
C53824 OR2X1_LOC_486/Y OR2X1_LOC_580/B 0.18fF
C53825 OR2X1_LOC_696/A OR2X1_LOC_744/A 0.87fF
C53826 OR2X1_LOC_702/A AND2X1_LOC_699/a_8_24# 0.02fF
C53827 OR2X1_LOC_160/B OR2X1_LOC_563/A 0.03fF
C53828 OR2X1_LOC_405/A OR2X1_LOC_728/a_36_216# 0.00fF
C53829 AND2X1_LOC_789/a_36_24# AND2X1_LOC_789/Y 0.01fF
C53830 OR2X1_LOC_92/Y OR2X1_LOC_268/Y 0.05fF
C53831 OR2X1_LOC_555/A AND2X1_LOC_257/a_8_24# 0.21fF
C53832 OR2X1_LOC_39/A OR2X1_LOC_13/B 0.84fF
C53833 OR2X1_LOC_456/a_36_216# D_GATE_366 0.00fF
C53834 AND2X1_LOC_275/a_8_24# OR2X1_LOC_549/A 0.04fF
C53835 AND2X1_LOC_715/Y OR2X1_LOC_744/A 0.07fF
C53836 OR2X1_LOC_220/B OR2X1_LOC_469/B 0.07fF
C53837 INPUT_0 OR2X1_LOC_828/Y 0.03fF
C53838 OR2X1_LOC_190/A OR2X1_LOC_161/B 0.03fF
C53839 OR2X1_LOC_269/B OR2X1_LOC_558/A 0.01fF
C53840 OR2X1_LOC_347/A OR2X1_LOC_347/a_8_216# 0.39fF
C53841 OR2X1_LOC_75/a_36_216# OR2X1_LOC_75/Y 0.00fF
C53842 AND2X1_LOC_461/a_36_24# OR2X1_LOC_46/A 0.00fF
C53843 AND2X1_LOC_571/A AND2X1_LOC_553/A 0.05fF
C53844 OR2X1_LOC_595/Y OR2X1_LOC_46/A 0.02fF
C53845 OR2X1_LOC_199/a_36_216# OR2X1_LOC_78/A 0.00fF
C53846 OR2X1_LOC_335/A OR2X1_LOC_808/a_8_216# 0.02fF
C53847 OR2X1_LOC_323/A AND2X1_LOC_717/Y 0.12fF
C53848 OR2X1_LOC_506/Y OR2X1_LOC_78/A 0.01fF
C53849 AND2X1_LOC_392/A AND2X1_LOC_541/Y 0.03fF
C53850 OR2X1_LOC_814/A OR2X1_LOC_351/a_8_216# 0.03fF
C53851 AND2X1_LOC_738/B AND2X1_LOC_788/a_8_24# 0.03fF
C53852 OR2X1_LOC_686/A OR2X1_LOC_686/B 0.13fF
C53853 AND2X1_LOC_211/B OR2X1_LOC_13/B 0.07fF
C53854 OR2X1_LOC_139/A OR2X1_LOC_474/Y 0.24fF
C53855 AND2X1_LOC_191/B AND2X1_LOC_285/a_8_24# 0.07fF
C53856 AND2X1_LOC_719/Y AND2X1_LOC_286/a_8_24# 0.01fF
C53857 AND2X1_LOC_352/a_8_24# AND2X1_LOC_337/a_8_24# 0.23fF
C53858 OR2X1_LOC_234/Y OR2X1_LOC_16/A 0.02fF
C53859 OR2X1_LOC_56/A AND2X1_LOC_476/Y 0.07fF
C53860 OR2X1_LOC_124/A OR2X1_LOC_6/B 0.06fF
C53861 AND2X1_LOC_549/Y AND2X1_LOC_657/Y 0.32fF
C53862 OR2X1_LOC_658/a_8_216# OR2X1_LOC_113/B 0.01fF
C53863 AND2X1_LOC_753/B AND2X1_LOC_44/Y 0.02fF
C53864 OR2X1_LOC_240/a_36_216# OR2X1_LOC_415/Y 0.03fF
C53865 OR2X1_LOC_155/A AND2X1_LOC_36/Y 0.11fF
C53866 AND2X1_LOC_196/Y OR2X1_LOC_172/a_8_216# 0.00fF
C53867 OR2X1_LOC_744/A OR2X1_LOC_131/a_36_216# 0.00fF
C53868 OR2X1_LOC_426/A OR2X1_LOC_12/Y 0.18fF
C53869 OR2X1_LOC_858/A OR2X1_LOC_114/B 0.03fF
C53870 VDD OR2X1_LOC_35/Y 0.13fF
C53871 OR2X1_LOC_482/Y AND2X1_LOC_861/B 0.11fF
C53872 AND2X1_LOC_500/Y AND2X1_LOC_657/Y 0.05fF
C53873 OR2X1_LOC_359/A VDD -0.00fF
C53874 AND2X1_LOC_773/Y AND2X1_LOC_649/B 0.10fF
C53875 OR2X1_LOC_502/A OR2X1_LOC_390/A 0.01fF
C53876 OR2X1_LOC_759/A OR2X1_LOC_59/Y 0.36fF
C53877 OR2X1_LOC_158/A OR2X1_LOC_58/a_36_216# 0.01fF
C53878 AND2X1_LOC_510/a_8_24# OR2X1_LOC_40/Y 0.17fF
C53879 OR2X1_LOC_523/B OR2X1_LOC_721/Y 0.00fF
C53880 OR2X1_LOC_97/A OR2X1_LOC_506/A 0.02fF
C53881 AND2X1_LOC_703/a_8_24# OR2X1_LOC_16/A 0.01fF
C53882 OR2X1_LOC_507/A AND2X1_LOC_41/A 0.64fF
C53883 OR2X1_LOC_693/Y OR2X1_LOC_48/B 0.01fF
C53884 OR2X1_LOC_850/B OR2X1_LOC_362/A 0.01fF
C53885 OR2X1_LOC_499/B AND2X1_LOC_18/Y 0.12fF
C53886 AND2X1_LOC_91/B OR2X1_LOC_845/a_8_216# 0.01fF
C53887 AND2X1_LOC_724/Y AND2X1_LOC_605/Y 0.00fF
C53888 OR2X1_LOC_199/a_8_216# OR2X1_LOC_375/A 0.03fF
C53889 AND2X1_LOC_231/Y OR2X1_LOC_265/Y 0.08fF
C53890 OR2X1_LOC_630/Y OR2X1_LOC_78/A 0.01fF
C53891 OR2X1_LOC_693/Y OR2X1_LOC_18/Y 0.01fF
C53892 OR2X1_LOC_666/A AND2X1_LOC_474/A 0.01fF
C53893 OR2X1_LOC_276/B OR2X1_LOC_68/B 0.07fF
C53894 OR2X1_LOC_87/A OR2X1_LOC_227/B 0.01fF
C53895 OR2X1_LOC_223/A OR2X1_LOC_742/B 0.03fF
C53896 AND2X1_LOC_554/Y OR2X1_LOC_595/A 0.17fF
C53897 OR2X1_LOC_464/a_8_216# OR2X1_LOC_471/B -0.00fF
C53898 OR2X1_LOC_494/Y OR2X1_LOC_517/A 0.00fF
C53899 OR2X1_LOC_643/A OR2X1_LOC_267/Y 0.03fF
C53900 OR2X1_LOC_852/a_8_216# AND2X1_LOC_824/B 0.06fF
C53901 OR2X1_LOC_633/a_8_216# OR2X1_LOC_78/A 0.01fF
C53902 OR2X1_LOC_124/Y OR2X1_LOC_267/Y 0.14fF
C53903 AND2X1_LOC_738/B OR2X1_LOC_677/a_36_216# 0.00fF
C53904 OR2X1_LOC_441/Y AND2X1_LOC_658/A 0.03fF
C53905 OR2X1_LOC_456/a_8_216# OR2X1_LOC_549/A -0.01fF
C53906 OR2X1_LOC_9/Y OR2X1_LOC_823/a_8_216# 0.01fF
C53907 OR2X1_LOC_9/Y AND2X1_LOC_62/a_36_24# 0.00fF
C53908 OR2X1_LOC_160/A OR2X1_LOC_729/a_8_216# 0.03fF
C53909 AND2X1_LOC_516/a_8_24# AND2X1_LOC_7/B 0.01fF
C53910 OR2X1_LOC_856/B AND2X1_LOC_387/a_8_24# 0.03fF
C53911 OR2X1_LOC_3/Y OR2X1_LOC_748/Y 0.02fF
C53912 OR2X1_LOC_589/A OR2X1_LOC_265/Y 0.22fF
C53913 OR2X1_LOC_635/A OR2X1_LOC_78/A 0.01fF
C53914 OR2X1_LOC_797/B OR2X1_LOC_375/A 0.00fF
C53915 OR2X1_LOC_533/Y OR2X1_LOC_43/A 0.39fF
C53916 INPUT_0 AND2X1_LOC_126/a_36_24# 0.00fF
C53917 OR2X1_LOC_769/B OR2X1_LOC_637/B 0.13fF
C53918 AND2X1_LOC_763/a_36_24# OR2X1_LOC_637/A 0.00fF
C53919 AND2X1_LOC_91/B OR2X1_LOC_602/a_8_216# 0.06fF
C53920 OR2X1_LOC_660/a_8_216# AND2X1_LOC_19/Y 0.02fF
C53921 AND2X1_LOC_95/Y AND2X1_LOC_323/a_36_24# 0.00fF
C53922 OR2X1_LOC_516/a_8_216# AND2X1_LOC_477/Y 0.01fF
C53923 AND2X1_LOC_356/B OR2X1_LOC_428/A 0.03fF
C53924 INPUT_1 AND2X1_LOC_750/a_36_24# 0.00fF
C53925 OR2X1_LOC_323/A OR2X1_LOC_64/Y 0.24fF
C53926 OR2X1_LOC_426/B OR2X1_LOC_71/a_8_216# 0.05fF
C53927 AND2X1_LOC_392/A OR2X1_LOC_316/Y 0.03fF
C53928 OR2X1_LOC_620/Y AND2X1_LOC_92/Y 0.07fF
C53929 OR2X1_LOC_280/Y OR2X1_LOC_428/A 0.01fF
C53930 AND2X1_LOC_717/B AND2X1_LOC_786/Y 0.09fF
C53931 AND2X1_LOC_31/Y OR2X1_LOC_318/B 0.22fF
C53932 OR2X1_LOC_358/A OR2X1_LOC_228/Y 0.05fF
C53933 AND2X1_LOC_132/a_8_24# OR2X1_LOC_66/A 0.01fF
C53934 AND2X1_LOC_732/a_36_24# OR2X1_LOC_48/B 0.01fF
C53935 OR2X1_LOC_821/Y OR2X1_LOC_585/A 0.02fF
C53936 OR2X1_LOC_186/Y OR2X1_LOC_355/B 0.01fF
C53937 OR2X1_LOC_256/Y OR2X1_LOC_494/a_36_216# 0.00fF
C53938 OR2X1_LOC_358/a_8_216# AND2X1_LOC_18/Y 0.01fF
C53939 OR2X1_LOC_659/Y AND2X1_LOC_3/Y 0.08fF
C53940 OR2X1_LOC_36/Y AND2X1_LOC_500/B 0.07fF
C53941 OR2X1_LOC_368/a_8_216# OR2X1_LOC_44/Y 0.02fF
C53942 OR2X1_LOC_653/Y AND2X1_LOC_41/A 0.07fF
C53943 OR2X1_LOC_8/Y AND2X1_LOC_342/Y 0.12fF
C53944 AND2X1_LOC_723/Y AND2X1_LOC_717/Y 0.13fF
C53945 OR2X1_LOC_79/A OR2X1_LOC_16/A 0.16fF
C53946 AND2X1_LOC_12/Y OR2X1_LOC_858/A 2.97fF
C53947 AND2X1_LOC_360/a_8_24# AND2X1_LOC_363/B 0.00fF
C53948 OR2X1_LOC_753/A AND2X1_LOC_194/Y 0.03fF
C53949 AND2X1_LOC_796/a_8_24# OR2X1_LOC_26/Y 0.06fF
C53950 OR2X1_LOC_187/a_36_216# AND2X1_LOC_866/B 0.00fF
C53951 OR2X1_LOC_54/Y OR2X1_LOC_397/Y 0.01fF
C53952 OR2X1_LOC_125/a_8_216# OR2X1_LOC_6/A 0.01fF
C53953 AND2X1_LOC_41/A OR2X1_LOC_833/B 0.19fF
C53954 OR2X1_LOC_364/B OR2X1_LOC_479/Y 0.06fF
C53955 AND2X1_LOC_478/a_8_24# AND2X1_LOC_220/Y 0.20fF
C53956 AND2X1_LOC_548/Y AND2X1_LOC_624/A 0.05fF
C53957 OR2X1_LOC_84/B OR2X1_LOC_786/A 1.10fF
C53958 AND2X1_LOC_40/Y OR2X1_LOC_637/a_8_216# 0.01fF
C53959 OR2X1_LOC_19/B AND2X1_LOC_7/B 0.19fF
C53960 OR2X1_LOC_348/Y OR2X1_LOC_269/B 0.02fF
C53961 OR2X1_LOC_696/A OR2X1_LOC_31/Y 0.56fF
C53962 OR2X1_LOC_323/A AND2X1_LOC_471/a_36_24# 0.00fF
C53963 AND2X1_LOC_562/B OR2X1_LOC_625/Y 0.03fF
C53964 OR2X1_LOC_154/A AND2X1_LOC_92/Y 0.37fF
C53965 OR2X1_LOC_160/A OR2X1_LOC_114/a_8_216# 0.02fF
C53966 OR2X1_LOC_130/A OR2X1_LOC_78/B 0.11fF
C53967 OR2X1_LOC_185/A OR2X1_LOC_808/A 0.03fF
C53968 VDD OR2X1_LOC_455/a_8_216# 0.00fF
C53969 OR2X1_LOC_8/Y AND2X1_LOC_852/a_36_24# -0.00fF
C53970 AND2X1_LOC_40/Y OR2X1_LOC_811/A 0.00fF
C53971 OR2X1_LOC_421/A OR2X1_LOC_763/Y 0.00fF
C53972 AND2X1_LOC_508/A AND2X1_LOC_621/Y 0.03fF
C53973 OR2X1_LOC_314/a_8_216# OR2X1_LOC_427/A 0.01fF
C53974 OR2X1_LOC_323/A OR2X1_LOC_417/A 0.13fF
C53975 OR2X1_LOC_528/a_36_216# OR2X1_LOC_74/A 0.02fF
C53976 AND2X1_LOC_24/a_36_24# OR2X1_LOC_130/A 0.01fF
C53977 OR2X1_LOC_744/A OR2X1_LOC_271/B 0.04fF
C53978 OR2X1_LOC_49/A AND2X1_LOC_119/a_8_24# -0.01fF
C53979 AND2X1_LOC_486/Y OR2X1_LOC_427/A 0.13fF
C53980 OR2X1_LOC_220/A OR2X1_LOC_738/B 0.12fF
C53981 OR2X1_LOC_18/Y AND2X1_LOC_651/a_8_24# 0.01fF
C53982 OR2X1_LOC_22/Y OR2X1_LOC_428/A 12.95fF
C53983 OR2X1_LOC_278/A OR2X1_LOC_16/A 0.00fF
C53984 OR2X1_LOC_40/Y AND2X1_LOC_148/Y 0.03fF
C53985 AND2X1_LOC_139/B AND2X1_LOC_139/a_8_24# 0.03fF
C53986 AND2X1_LOC_580/B AND2X1_LOC_663/A 0.03fF
C53987 AND2X1_LOC_48/A OR2X1_LOC_706/a_8_216# 0.01fF
C53988 OR2X1_LOC_346/B OR2X1_LOC_78/A 0.03fF
C53989 AND2X1_LOC_392/A AND2X1_LOC_390/B 0.02fF
C53990 VDD AND2X1_LOC_640/Y 0.13fF
C53991 OR2X1_LOC_175/Y AND2X1_LOC_47/Y 0.42fF
C53992 INPUT_3 AND2X1_LOC_62/a_8_24# 0.01fF
C53993 OR2X1_LOC_759/A AND2X1_LOC_711/Y 0.00fF
C53994 AND2X1_LOC_564/B OR2X1_LOC_95/Y 0.14fF
C53995 OR2X1_LOC_22/Y OR2X1_LOC_595/A 2.95fF
C53996 AND2X1_LOC_772/B AND2X1_LOC_489/Y 0.18fF
C53997 AND2X1_LOC_125/a_8_24# OR2X1_LOC_805/A 0.06fF
C53998 OR2X1_LOC_653/Y OR2X1_LOC_662/A 0.01fF
C53999 OR2X1_LOC_264/Y OR2X1_LOC_520/Y 0.02fF
C54000 OR2X1_LOC_3/Y AND2X1_LOC_404/B 0.01fF
C54001 AND2X1_LOC_9/a_36_24# AND2X1_LOC_852/B 0.01fF
C54002 OR2X1_LOC_185/Y OR2X1_LOC_216/A 0.07fF
C54003 OR2X1_LOC_95/Y OR2X1_LOC_368/Y 0.08fF
C54004 OR2X1_LOC_207/B AND2X1_LOC_7/Y 0.00fF
C54005 OR2X1_LOC_108/Y AND2X1_LOC_830/a_8_24# 0.03fF
C54006 OR2X1_LOC_479/Y AND2X1_LOC_70/Y 0.12fF
C54007 VDD OR2X1_LOC_681/Y 0.12fF
C54008 OR2X1_LOC_368/A OR2X1_LOC_368/Y 0.06fF
C54009 OR2X1_LOC_18/Y AND2X1_LOC_621/Y 0.06fF
C54010 OR2X1_LOC_691/Y AND2X1_LOC_47/Y 0.03fF
C54011 AND2X1_LOC_47/Y AND2X1_LOC_417/a_8_24# 0.04fF
C54012 OR2X1_LOC_92/Y OR2X1_LOC_248/a_8_216# 0.01fF
C54013 AND2X1_LOC_510/a_8_24# OR2X1_LOC_7/A 0.01fF
C54014 AND2X1_LOC_51/Y OR2X1_LOC_35/a_8_216# 0.01fF
C54015 OR2X1_LOC_132/Y OR2X1_LOC_272/Y 0.09fF
C54016 OR2X1_LOC_227/a_8_216# OR2X1_LOC_641/A 0.03fF
C54017 AND2X1_LOC_572/Y AND2X1_LOC_573/A 0.08fF
C54018 OR2X1_LOC_235/B OR2X1_LOC_74/A 0.02fF
C54019 OR2X1_LOC_448/Y OR2X1_LOC_161/A 0.48fF
C54020 AND2X1_LOC_390/B AND2X1_LOC_436/a_8_24# 0.02fF
C54021 OR2X1_LOC_421/a_36_216# OR2X1_LOC_743/A 0.00fF
C54022 VDD OR2X1_LOC_416/Y 0.64fF
C54023 OR2X1_LOC_431/a_8_216# OR2X1_LOC_56/A 0.03fF
C54024 OR2X1_LOC_179/a_8_216# OR2X1_LOC_485/A 0.01fF
C54025 OR2X1_LOC_249/a_8_216# OR2X1_LOC_579/B 0.40fF
C54026 OR2X1_LOC_92/Y AND2X1_LOC_294/a_8_24# 0.01fF
C54027 OR2X1_LOC_479/Y OR2X1_LOC_703/A 0.03fF
C54028 OR2X1_LOC_744/A AND2X1_LOC_663/B 0.03fF
C54029 OR2X1_LOC_8/Y OR2X1_LOC_54/Y 1.99fF
C54030 AND2X1_LOC_215/Y OR2X1_LOC_22/Y 0.01fF
C54031 OR2X1_LOC_641/Y OR2X1_LOC_650/Y 0.02fF
C54032 OR2X1_LOC_429/Y OR2X1_LOC_425/a_36_216# 0.01fF
C54033 OR2X1_LOC_631/B OR2X1_LOC_833/B 0.02fF
C54034 OR2X1_LOC_130/A OR2X1_LOC_375/A 0.00fF
C54035 AND2X1_LOC_101/B OR2X1_LOC_278/Y 0.17fF
C54036 OR2X1_LOC_779/Y AND2X1_LOC_44/Y 0.01fF
C54037 OR2X1_LOC_856/B OR2X1_LOC_574/A 0.07fF
C54038 AND2X1_LOC_729/Y AND2X1_LOC_598/a_8_24# 0.04fF
C54039 AND2X1_LOC_185/a_8_24# AND2X1_LOC_631/Y 0.01fF
C54040 AND2X1_LOC_852/Y AND2X1_LOC_573/A 0.07fF
C54041 AND2X1_LOC_303/A AND2X1_LOC_303/B 0.03fF
C54042 AND2X1_LOC_44/Y OR2X1_LOC_330/a_8_216# 0.05fF
C54043 AND2X1_LOC_392/A AND2X1_LOC_863/Y 0.02fF
C54044 AND2X1_LOC_56/B AND2X1_LOC_233/a_36_24# 0.00fF
C54045 OR2X1_LOC_214/B OR2X1_LOC_161/B 0.07fF
C54046 OR2X1_LOC_254/B OR2X1_LOC_631/B 0.05fF
C54047 AND2X1_LOC_729/Y OR2X1_LOC_26/Y 0.03fF
C54048 OR2X1_LOC_185/Y OR2X1_LOC_802/Y 0.01fF
C54049 OR2X1_LOC_62/B OR2X1_LOC_78/B 0.03fF
C54050 AND2X1_LOC_364/Y OR2X1_LOC_46/A 0.03fF
C54051 OR2X1_LOC_516/A OR2X1_LOC_52/B 0.03fF
C54052 D_GATE_662 D_INPUT_1 0.02fF
C54053 AND2X1_LOC_354/Y AND2X1_LOC_390/B 0.01fF
C54054 OR2X1_LOC_298/Y OR2X1_LOC_7/A 0.05fF
C54055 AND2X1_LOC_103/a_8_24# AND2X1_LOC_15/a_8_24# 0.23fF
C54056 OR2X1_LOC_68/B AND2X1_LOC_226/a_8_24# 0.02fF
C54057 OR2X1_LOC_220/a_8_216# OR2X1_LOC_739/B 0.14fF
C54058 OR2X1_LOC_428/A OR2X1_LOC_387/a_8_216# 0.06fF
C54059 AND2X1_LOC_650/a_8_24# OR2X1_LOC_48/B 0.05fF
C54060 OR2X1_LOC_375/A AND2X1_LOC_612/a_8_24# 0.10fF
C54061 AND2X1_LOC_795/Y AND2X1_LOC_795/a_36_24# 0.01fF
C54062 OR2X1_LOC_473/Y OR2X1_LOC_61/Y 0.00fF
C54063 AND2X1_LOC_729/Y OR2X1_LOC_89/A 0.03fF
C54064 AND2X1_LOC_219/A OR2X1_LOC_598/A 0.09fF
C54065 OR2X1_LOC_287/B AND2X1_LOC_251/a_8_24# 0.00fF
C54066 AND2X1_LOC_36/Y D_GATE_366 0.04fF
C54067 OR2X1_LOC_210/B OR2X1_LOC_87/A 0.01fF
C54068 OR2X1_LOC_160/A AND2X1_LOC_42/B 0.71fF
C54069 OR2X1_LOC_246/a_8_216# OR2X1_LOC_753/A 0.04fF
C54070 OR2X1_LOC_18/Y AND2X1_LOC_650/a_8_24# 0.01fF
C54071 AND2X1_LOC_784/A OR2X1_LOC_26/Y 0.05fF
C54072 AND2X1_LOC_219/a_36_24# AND2X1_LOC_476/A 0.01fF
C54073 OR2X1_LOC_532/B OR2X1_LOC_78/Y 0.00fF
C54074 OR2X1_LOC_723/B OR2X1_LOC_593/B 0.01fF
C54075 OR2X1_LOC_51/Y AND2X1_LOC_796/Y 0.00fF
C54076 OR2X1_LOC_62/B OR2X1_LOC_721/Y 0.05fF
C54077 AND2X1_LOC_70/Y AND2X1_LOC_681/a_8_24# 0.01fF
C54078 OR2X1_LOC_303/B OR2X1_LOC_605/Y 0.81fF
C54079 OR2X1_LOC_810/A OR2X1_LOC_269/B 0.05fF
C54080 OR2X1_LOC_260/Y AND2X1_LOC_261/a_8_24# 0.01fF
C54081 OR2X1_LOC_521/Y AND2X1_LOC_116/B 0.81fF
C54082 OR2X1_LOC_837/B OR2X1_LOC_46/A 0.07fF
C54083 AND2X1_LOC_723/Y OR2X1_LOC_417/A 0.08fF
C54084 AND2X1_LOC_597/a_8_24# AND2X1_LOC_387/B 0.03fF
C54085 OR2X1_LOC_682/Y OR2X1_LOC_52/B 0.04fF
C54086 OR2X1_LOC_497/Y OR2X1_LOC_239/Y 0.16fF
C54087 OR2X1_LOC_3/Y OR2X1_LOC_36/Y 1.40fF
C54088 OR2X1_LOC_223/A OR2X1_LOC_191/a_36_216# 0.00fF
C54089 OR2X1_LOC_231/B AND2X1_LOC_31/Y 0.01fF
C54090 OR2X1_LOC_864/a_8_216# OR2X1_LOC_269/B 0.01fF
C54091 OR2X1_LOC_178/Y OR2X1_LOC_47/Y 0.02fF
C54092 OR2X1_LOC_224/Y OR2X1_LOC_59/Y 0.01fF
C54093 OR2X1_LOC_377/A OR2X1_LOC_121/B 0.02fF
C54094 OR2X1_LOC_419/Y AND2X1_LOC_500/B 0.04fF
C54095 OR2X1_LOC_78/B AND2X1_LOC_88/Y 0.03fF
C54096 OR2X1_LOC_185/Y OR2X1_LOC_846/B 0.00fF
C54097 OR2X1_LOC_547/B OR2X1_LOC_471/Y 0.03fF
C54098 OR2X1_LOC_464/A OR2X1_LOC_440/A 0.02fF
C54099 AND2X1_LOC_287/B OR2X1_LOC_437/A 0.09fF
C54100 OR2X1_LOC_541/A D_INPUT_1 0.03fF
C54101 OR2X1_LOC_78/B AND2X1_LOC_39/Y 0.01fF
C54102 OR2X1_LOC_695/a_8_216# OR2X1_LOC_31/Y 0.00fF
C54103 OR2X1_LOC_446/a_8_216# AND2X1_LOC_3/Y 0.01fF
C54104 OR2X1_LOC_646/a_8_216# OR2X1_LOC_647/A 0.01fF
C54105 OR2X1_LOC_62/B OR2X1_LOC_375/A 0.10fF
C54106 AND2X1_LOC_52/a_36_24# OR2X1_LOC_651/A 0.01fF
C54107 OR2X1_LOC_335/A OR2X1_LOC_593/B 1.48fF
C54108 OR2X1_LOC_816/A OR2X1_LOC_437/A 0.02fF
C54109 AND2X1_LOC_86/B AND2X1_LOC_42/B 0.01fF
C54110 AND2X1_LOC_578/A AND2X1_LOC_717/B 2.98fF
C54111 AND2X1_LOC_281/a_36_24# OR2X1_LOC_269/B 0.01fF
C54112 AND2X1_LOC_370/a_36_24# OR2X1_LOC_437/A 0.00fF
C54113 OR2X1_LOC_836/A OR2X1_LOC_19/B 0.03fF
C54114 OR2X1_LOC_7/A OR2X1_LOC_27/a_8_216# 0.01fF
C54115 OR2X1_LOC_256/Y OR2X1_LOC_47/Y 0.06fF
C54116 AND2X1_LOC_367/A AND2X1_LOC_721/A 0.03fF
C54117 OR2X1_LOC_92/Y AND2X1_LOC_648/B 0.05fF
C54118 OR2X1_LOC_124/A OR2X1_LOC_598/A 0.01fF
C54119 AND2X1_LOC_56/B OR2X1_LOC_443/Y 0.13fF
C54120 OR2X1_LOC_185/A OR2X1_LOC_223/a_8_216# 0.05fF
C54121 OR2X1_LOC_99/A AND2X1_LOC_92/Y 0.03fF
C54122 OR2X1_LOC_817/a_8_216# OR2X1_LOC_817/Y -0.00fF
C54123 D_INPUT_0 AND2X1_LOC_824/a_8_24# 0.01fF
C54124 OR2X1_LOC_490/Y AND2X1_LOC_140/a_8_24# 0.02fF
C54125 OR2X1_LOC_78/A OR2X1_LOC_196/a_8_216# 0.01fF
C54126 AND2X1_LOC_53/a_36_24# OR2X1_LOC_651/A 0.00fF
C54127 OR2X1_LOC_624/B AND2X1_LOC_42/B 0.05fF
C54128 AND2X1_LOC_326/a_8_24# OR2X1_LOC_6/A 0.01fF
C54129 AND2X1_LOC_64/Y AND2X1_LOC_238/a_8_24# 0.01fF
C54130 AND2X1_LOC_712/B OR2X1_LOC_52/B 0.02fF
C54131 AND2X1_LOC_101/B OR2X1_LOC_19/B 0.01fF
C54132 OR2X1_LOC_756/B OR2X1_LOC_544/a_8_216# 0.01fF
C54133 OR2X1_LOC_46/A OR2X1_LOC_49/a_36_216# 0.03fF
C54134 OR2X1_LOC_395/Y OR2X1_LOC_415/Y 0.28fF
C54135 AND2X1_LOC_18/Y OR2X1_LOC_348/B 0.77fF
C54136 AND2X1_LOC_78/a_8_24# OR2X1_LOC_64/Y 0.01fF
C54137 VDD OR2X1_LOC_80/A 0.47fF
C54138 AND2X1_LOC_191/B AND2X1_LOC_563/Y 0.03fF
C54139 AND2X1_LOC_13/a_8_24# OR2X1_LOC_193/A 0.00fF
C54140 AND2X1_LOC_70/Y OR2X1_LOC_68/B 0.03fF
C54141 AND2X1_LOC_212/A OR2X1_LOC_437/A 0.00fF
C54142 OR2X1_LOC_491/a_8_216# OR2X1_LOC_437/A 0.02fF
C54143 OR2X1_LOC_394/a_36_216# OR2X1_LOC_598/A 0.03fF
C54144 AND2X1_LOC_56/B AND2X1_LOC_821/a_8_24# 0.05fF
C54145 OR2X1_LOC_73/a_8_216# OR2X1_LOC_46/A 0.01fF
C54146 AND2X1_LOC_535/a_36_24# OR2X1_LOC_534/Y 0.00fF
C54147 OR2X1_LOC_831/A OR2X1_LOC_777/B 0.03fF
C54148 AND2X1_LOC_7/a_36_24# AND2X1_LOC_7/Y 0.00fF
C54149 OR2X1_LOC_680/A AND2X1_LOC_796/Y 0.09fF
C54150 OR2X1_LOC_538/A AND2X1_LOC_31/Y 0.20fF
C54151 AND2X1_LOC_621/Y AND2X1_LOC_620/Y 0.12fF
C54152 AND2X1_LOC_142/a_8_24# OR2X1_LOC_705/B 0.01fF
C54153 OR2X1_LOC_185/A OR2X1_LOC_795/a_8_216# 0.01fF
C54154 D_INPUT_5 OR2X1_LOC_70/A 0.09fF
C54155 AND2X1_LOC_514/Y AND2X1_LOC_324/a_8_24# 0.01fF
C54156 OR2X1_LOC_670/a_8_216# D_INPUT_3 0.01fF
C54157 OR2X1_LOC_262/Y OR2X1_LOC_72/a_8_216# 0.09fF
C54158 AND2X1_LOC_3/Y AND2X1_LOC_7/Y 0.03fF
C54159 OR2X1_LOC_629/Y OR2X1_LOC_598/A 0.01fF
C54160 OR2X1_LOC_834/a_8_216# OR2X1_LOC_779/B 0.01fF
C54161 OR2X1_LOC_777/B OR2X1_LOC_356/a_8_216# 0.07fF
C54162 AND2X1_LOC_260/a_8_24# OR2X1_LOC_46/A 0.03fF
C54163 OR2X1_LOC_846/B AND2X1_LOC_816/a_36_24# 0.00fF
C54164 OR2X1_LOC_696/A AND2X1_LOC_464/A 0.10fF
C54165 OR2X1_LOC_48/Y AND2X1_LOC_196/Y 0.01fF
C54166 D_INPUT_5 AND2X1_LOC_31/Y 4.74fF
C54167 OR2X1_LOC_62/A OR2X1_LOC_26/Y 0.00fF
C54168 AND2X1_LOC_729/Y OR2X1_LOC_419/a_8_216# 0.03fF
C54169 OR2X1_LOC_185/A OR2X1_LOC_374/Y 0.03fF
C54170 OR2X1_LOC_619/Y AND2X1_LOC_205/a_36_24# 0.01fF
C54171 AND2X1_LOC_572/a_8_24# AND2X1_LOC_554/a_8_24# 0.23fF
C54172 OR2X1_LOC_619/Y OR2X1_LOC_163/a_8_216# 0.00fF
C54173 OR2X1_LOC_406/Y AND2X1_LOC_721/Y 0.01fF
C54174 AND2X1_LOC_605/Y OR2X1_LOC_423/Y 0.13fF
C54175 AND2X1_LOC_22/a_8_24# AND2X1_LOC_31/Y 0.01fF
C54176 AND2X1_LOC_554/B D_INPUT_3 0.01fF
C54177 OR2X1_LOC_476/B OR2X1_LOC_648/a_36_216# 0.01fF
C54178 OR2X1_LOC_600/A OR2X1_LOC_183/Y 0.04fF
C54179 AND2X1_LOC_474/A OR2X1_LOC_13/B 0.01fF
C54180 OR2X1_LOC_753/A OR2X1_LOC_396/Y 0.03fF
C54181 AND2X1_LOC_491/a_8_24# OR2X1_LOC_532/B 0.11fF
C54182 OR2X1_LOC_188/Y OR2X1_LOC_161/B 0.03fF
C54183 OR2X1_LOC_824/a_36_216# OR2X1_LOC_62/A 0.00fF
C54184 AND2X1_LOC_91/B OR2X1_LOC_673/a_8_216# 0.49fF
C54185 AND2X1_LOC_12/Y AND2X1_LOC_31/Y 0.18fF
C54186 OR2X1_LOC_84/B OR2X1_LOC_84/Y 0.03fF
C54187 OR2X1_LOC_831/A OR2X1_LOC_831/B 0.34fF
C54188 AND2X1_LOC_351/a_8_24# AND2X1_LOC_350/B 0.01fF
C54189 AND2X1_LOC_445/a_36_24# OR2X1_LOC_428/A 0.00fF
C54190 AND2X1_LOC_721/A OR2X1_LOC_74/A 0.60fF
C54191 AND2X1_LOC_40/Y OR2X1_LOC_777/B 10.58fF
C54192 OR2X1_LOC_18/Y OR2X1_LOC_71/A 0.00fF
C54193 OR2X1_LOC_169/a_8_216# OR2X1_LOC_568/A 0.03fF
C54194 OR2X1_LOC_135/Y OR2X1_LOC_16/A 2.07fF
C54195 OR2X1_LOC_333/B OR2X1_LOC_339/Y 0.11fF
C54196 VDD OR2X1_LOC_115/B 0.07fF
C54197 OR2X1_LOC_841/B AND2X1_LOC_31/Y 0.03fF
C54198 OR2X1_LOC_468/Y OR2X1_LOC_568/A 0.01fF
C54199 OR2X1_LOC_182/B OR2X1_LOC_352/a_36_216# 0.00fF
C54200 OR2X1_LOC_48/B AND2X1_LOC_592/a_36_24# 0.01fF
C54201 OR2X1_LOC_501/B OR2X1_LOC_501/A 0.11fF
C54202 OR2X1_LOC_468/Y OR2X1_LOC_578/B 0.01fF
C54203 OR2X1_LOC_40/Y OR2X1_LOC_310/a_8_216# 0.01fF
C54204 AND2X1_LOC_150/a_36_24# OR2X1_LOC_161/B 0.00fF
C54205 INPUT_1 OR2X1_LOC_751/a_8_216# 0.02fF
C54206 AND2X1_LOC_593/Y OR2X1_LOC_13/B 0.02fF
C54207 AND2X1_LOC_350/Y OR2X1_LOC_289/Y 0.27fF
C54208 AND2X1_LOC_715/A AND2X1_LOC_473/Y 0.03fF
C54209 AND2X1_LOC_95/Y OR2X1_LOC_349/B 0.01fF
C54210 AND2X1_LOC_807/Y OR2X1_LOC_437/A 0.15fF
C54211 AND2X1_LOC_721/Y OR2X1_LOC_496/a_8_216# 0.01fF
C54212 OR2X1_LOC_89/A OR2X1_LOC_88/Y 0.00fF
C54213 OR2X1_LOC_325/B OR2X1_LOC_161/B 0.01fF
C54214 OR2X1_LOC_686/B OR2X1_LOC_161/B 0.27fF
C54215 OR2X1_LOC_203/Y AND2X1_LOC_268/a_36_24# 0.00fF
C54216 OR2X1_LOC_85/A OR2X1_LOC_13/B 0.04fF
C54217 AND2X1_LOC_705/Y OR2X1_LOC_600/A 0.14fF
C54218 AND2X1_LOC_851/B AND2X1_LOC_866/A 0.07fF
C54219 OR2X1_LOC_89/A AND2X1_LOC_772/a_36_24# 0.00fF
C54220 AND2X1_LOC_557/a_8_24# AND2X1_LOC_657/A 0.03fF
C54221 OR2X1_LOC_490/Y AND2X1_LOC_217/a_8_24# 0.04fF
C54222 AND2X1_LOC_447/Y OR2X1_LOC_12/Y 0.16fF
C54223 OR2X1_LOC_507/a_8_216# AND2X1_LOC_64/Y 0.01fF
C54224 AND2X1_LOC_65/A AND2X1_LOC_18/Y 0.05fF
C54225 AND2X1_LOC_64/Y OR2X1_LOC_637/A 0.03fF
C54226 AND2X1_LOC_19/Y AND2X1_LOC_44/Y 0.01fF
C54227 OR2X1_LOC_624/Y OR2X1_LOC_474/B 0.02fF
C54228 OR2X1_LOC_179/a_36_216# AND2X1_LOC_465/A 0.00fF
C54229 AND2X1_LOC_787/A OR2X1_LOC_91/A 0.00fF
C54230 OR2X1_LOC_206/a_8_216# OR2X1_LOC_68/B 0.01fF
C54231 AND2X1_LOC_64/Y OR2X1_LOC_264/Y 0.10fF
C54232 OR2X1_LOC_295/Y AND2X1_LOC_848/A 0.02fF
C54233 OR2X1_LOC_583/Y OR2X1_LOC_584/Y 0.09fF
C54234 AND2X1_LOC_784/Y OR2X1_LOC_40/Y 0.01fF
C54235 AND2X1_LOC_339/B OR2X1_LOC_426/B 0.03fF
C54236 AND2X1_LOC_732/a_8_24# AND2X1_LOC_713/a_8_24# 0.23fF
C54237 OR2X1_LOC_404/Y OR2X1_LOC_68/B 0.08fF
C54238 OR2X1_LOC_813/A OR2X1_LOC_86/A 0.37fF
C54239 AND2X1_LOC_454/a_8_24# OR2X1_LOC_421/Y 0.01fF
C54240 OR2X1_LOC_510/A AND2X1_LOC_18/Y 0.09fF
C54241 AND2X1_LOC_716/Y OR2X1_LOC_136/Y 0.01fF
C54242 OR2X1_LOC_124/B OR2X1_LOC_641/A 0.07fF
C54243 OR2X1_LOC_359/a_36_216# OR2X1_LOC_362/A 0.00fF
C54244 OR2X1_LOC_304/a_8_216# AND2X1_LOC_654/B 0.00fF
C54245 AND2X1_LOC_539/Y AND2X1_LOC_841/B 0.08fF
C54246 OR2X1_LOC_440/B OR2X1_LOC_440/a_8_216# 0.47fF
C54247 OR2X1_LOC_715/B OR2X1_LOC_702/a_8_216# 0.03fF
C54248 OR2X1_LOC_349/a_36_216# OR2X1_LOC_362/A 0.00fF
C54249 AND2X1_LOC_22/Y OR2X1_LOC_61/B 0.02fF
C54250 AND2X1_LOC_729/Y AND2X1_LOC_590/a_8_24# 0.01fF
C54251 D_INPUT_4 AND2X1_LOC_44/Y 0.04fF
C54252 OR2X1_LOC_124/a_8_216# VDD 0.21fF
C54253 AND2X1_LOC_566/B OR2X1_LOC_91/A 0.10fF
C54254 OR2X1_LOC_469/Y OR2X1_LOC_161/B 0.05fF
C54255 OR2X1_LOC_40/Y AND2X1_LOC_434/Y 0.14fF
C54256 OR2X1_LOC_319/B AND2X1_LOC_534/a_8_24# -0.00fF
C54257 OR2X1_LOC_488/Y OR2X1_LOC_437/A 0.05fF
C54258 OR2X1_LOC_175/Y OR2X1_LOC_506/A 0.07fF
C54259 OR2X1_LOC_185/A OR2X1_LOC_392/B 0.03fF
C54260 AND2X1_LOC_56/B AND2X1_LOC_763/B 0.51fF
C54261 OR2X1_LOC_160/A AND2X1_LOC_224/a_8_24# 0.01fF
C54262 AND2X1_LOC_40/Y OR2X1_LOC_344/A 0.09fF
C54263 OR2X1_LOC_104/a_8_216# VDD 0.00fF
C54264 OR2X1_LOC_427/A AND2X1_LOC_457/a_8_24# 0.01fF
C54265 AND2X1_LOC_392/A OR2X1_LOC_744/A 0.13fF
C54266 OR2X1_LOC_788/a_36_216# OR2X1_LOC_161/B 0.01fF
C54267 OR2X1_LOC_97/A AND2X1_LOC_95/Y 0.06fF
C54268 OR2X1_LOC_520/a_8_216# OR2X1_LOC_66/A 0.14fF
C54269 OR2X1_LOC_666/A OR2X1_LOC_51/Y 0.00fF
C54270 OR2X1_LOC_160/B OR2X1_LOC_632/Y 0.08fF
C54271 OR2X1_LOC_97/A OR2X1_LOC_633/Y 0.91fF
C54272 OR2X1_LOC_134/a_8_216# AND2X1_LOC_560/B 0.03fF
C54273 OR2X1_LOC_114/Y OR2X1_LOC_140/B 0.62fF
C54274 AND2X1_LOC_297/a_8_24# AND2X1_LOC_248/a_8_24# 0.23fF
C54275 AND2X1_LOC_555/Y GATE_366 0.03fF
C54276 AND2X1_LOC_649/B OR2X1_LOC_12/Y 0.46fF
C54277 OR2X1_LOC_468/A OR2X1_LOC_78/B 0.05fF
C54278 AND2X1_LOC_717/a_8_24# AND2X1_LOC_464/A 0.01fF
C54279 OR2X1_LOC_695/Y OR2X1_LOC_91/A 0.01fF
C54280 AND2X1_LOC_727/A OR2X1_LOC_437/A 0.03fF
C54281 AND2X1_LOC_64/Y OR2X1_LOC_643/A 0.18fF
C54282 OR2X1_LOC_39/A OR2X1_LOC_428/A 0.05fF
C54283 OR2X1_LOC_770/A OR2X1_LOC_848/A 0.09fF
C54284 AND2X1_LOC_64/Y OR2X1_LOC_778/Y 0.07fF
C54285 AND2X1_LOC_848/Y AND2X1_LOC_244/A 0.00fF
C54286 OR2X1_LOC_319/B AND2X1_LOC_110/Y 0.38fF
C54287 AND2X1_LOC_21/Y AND2X1_LOC_763/B 0.01fF
C54288 OR2X1_LOC_36/Y AND2X1_LOC_201/Y 0.28fF
C54289 OR2X1_LOC_186/Y OR2X1_LOC_624/A 0.05fF
C54290 AND2X1_LOC_573/Y AND2X1_LOC_474/Y 0.05fF
C54291 AND2X1_LOC_448/Y OR2X1_LOC_12/Y 0.08fF
C54292 OR2X1_LOC_834/A AND2X1_LOC_306/a_8_24# 0.21fF
C54293 AND2X1_LOC_458/Y AND2X1_LOC_464/A 0.10fF
C54294 VDD OR2X1_LOC_840/A 2.44fF
C54295 OR2X1_LOC_39/A OR2X1_LOC_595/A 0.03fF
C54296 AND2X1_LOC_553/A OR2X1_LOC_600/A 0.09fF
C54297 AND2X1_LOC_729/Y OR2X1_LOC_167/a_8_216# 0.04fF
C54298 AND2X1_LOC_861/B AND2X1_LOC_861/a_8_24# 0.01fF
C54299 OR2X1_LOC_318/Y AND2X1_LOC_110/Y 0.00fF
C54300 AND2X1_LOC_533/a_8_24# OR2X1_LOC_356/A 0.24fF
C54301 OR2X1_LOC_673/Y AND2X1_LOC_44/Y 0.02fF
C54302 AND2X1_LOC_810/A AND2X1_LOC_319/A 0.00fF
C54303 OR2X1_LOC_624/Y OR2X1_LOC_658/a_8_216# 0.02fF
C54304 OR2X1_LOC_661/a_8_216# OR2X1_LOC_661/A 0.39fF
C54305 OR2X1_LOC_502/A AND2X1_LOC_404/B 0.07fF
C54306 AND2X1_LOC_795/Y AND2X1_LOC_222/Y 0.02fF
C54307 OR2X1_LOC_753/A OR2X1_LOC_816/A 0.51fF
C54308 OR2X1_LOC_695/a_8_216# OR2X1_LOC_694/Y 0.41fF
C54309 OR2X1_LOC_600/A AND2X1_LOC_804/Y 0.09fF
C54310 AND2X1_LOC_716/Y OR2X1_LOC_51/Y 0.01fF
C54311 AND2X1_LOC_449/Y OR2X1_LOC_421/Y 0.01fF
C54312 OR2X1_LOC_426/B OR2X1_LOC_586/a_8_216# 0.05fF
C54313 VDD OR2X1_LOC_281/a_8_216# 0.21fF
C54314 OR2X1_LOC_95/Y OR2X1_LOC_437/A 0.34fF
C54315 AND2X1_LOC_773/Y AND2X1_LOC_264/a_8_24# 0.03fF
C54316 OR2X1_LOC_561/Y OR2X1_LOC_391/A 0.02fF
C54317 OR2X1_LOC_39/Y AND2X1_LOC_377/Y 0.80fF
C54318 OR2X1_LOC_377/A OR2X1_LOC_621/B 0.05fF
C54319 AND2X1_LOC_440/a_8_24# OR2X1_LOC_437/A 0.15fF
C54320 OR2X1_LOC_161/A OR2X1_LOC_629/B 0.51fF
C54321 AND2X1_LOC_326/B AND2X1_LOC_841/B 0.23fF
C54322 AND2X1_LOC_391/a_8_24# OR2X1_LOC_91/A 0.07fF
C54323 OR2X1_LOC_43/A AND2X1_LOC_809/a_8_24# 0.01fF
C54324 AND2X1_LOC_476/A OR2X1_LOC_300/a_8_216# 0.03fF
C54325 OR2X1_LOC_814/A AND2X1_LOC_36/Y 0.02fF
C54326 AND2X1_LOC_728/Y OR2X1_LOC_40/Y 0.03fF
C54327 OR2X1_LOC_91/Y AND2X1_LOC_476/Y 0.09fF
C54328 OR2X1_LOC_91/Y AND2X1_LOC_362/B 0.04fF
C54329 AND2X1_LOC_211/B OR2X1_LOC_428/A 0.07fF
C54330 OR2X1_LOC_816/A OR2X1_LOC_754/a_8_216# 0.03fF
C54331 OR2X1_LOC_67/Y OR2X1_LOC_80/A 0.09fF
C54332 OR2X1_LOC_653/Y OR2X1_LOC_648/A 0.75fF
C54333 AND2X1_LOC_140/a_36_24# AND2X1_LOC_772/Y 0.00fF
C54334 AND2X1_LOC_110/Y OR2X1_LOC_805/A 0.05fF
C54335 AND2X1_LOC_360/a_36_24# OR2X1_LOC_91/A 0.00fF
C54336 AND2X1_LOC_81/B OR2X1_LOC_786/A 0.00fF
C54337 AND2X1_LOC_421/a_8_24# AND2X1_LOC_41/A 0.01fF
C54338 OR2X1_LOC_429/Y OR2X1_LOC_428/A 0.02fF
C54339 AND2X1_LOC_42/B OR2X1_LOC_266/A 0.23fF
C54340 OR2X1_LOC_48/B OR2X1_LOC_59/Y 11.05fF
C54341 OR2X1_LOC_408/a_36_216# INPUT_6 0.03fF
C54342 AND2X1_LOC_215/Y OR2X1_LOC_39/A 0.01fF
C54343 VDD AND2X1_LOC_145/a_8_24# 0.00fF
C54344 OR2X1_LOC_170/Y OR2X1_LOC_566/Y 0.34fF
C54345 AND2X1_LOC_48/a_8_24# AND2X1_LOC_615/a_8_24# 0.23fF
C54346 OR2X1_LOC_541/A OR2X1_LOC_737/A 0.01fF
C54347 AND2X1_LOC_554/Y AND2X1_LOC_772/B 0.39fF
C54348 OR2X1_LOC_45/Y AND2X1_LOC_434/a_36_24# 0.01fF
C54349 OR2X1_LOC_539/a_8_216# OR2X1_LOC_66/A 0.02fF
C54350 OR2X1_LOC_235/B OR2X1_LOC_668/a_8_216# 0.00fF
C54351 OR2X1_LOC_351/B OR2X1_LOC_864/A 0.79fF
C54352 OR2X1_LOC_270/Y OR2X1_LOC_367/a_36_216# 0.00fF
C54353 AND2X1_LOC_321/a_8_24# AND2X1_LOC_41/A 0.10fF
C54354 OR2X1_LOC_18/Y OR2X1_LOC_59/Y 0.68fF
C54355 AND2X1_LOC_3/Y OR2X1_LOC_390/A 0.03fF
C54356 AND2X1_LOC_561/a_8_24# OR2X1_LOC_71/Y -0.00fF
C54357 VDD OR2X1_LOC_222/A 0.07fF
C54358 AND2X1_LOC_40/Y OR2X1_LOC_254/A 0.01fF
C54359 AND2X1_LOC_391/Y OR2X1_LOC_127/a_8_216# 0.03fF
C54360 OR2X1_LOC_36/Y AND2X1_LOC_606/a_36_24# 0.01fF
C54361 AND2X1_LOC_702/a_36_24# OR2X1_LOC_59/Y 0.00fF
C54362 OR2X1_LOC_127/a_8_216# OR2X1_LOC_91/A 0.05fF
C54363 OR2X1_LOC_858/A AND2X1_LOC_59/Y 0.02fF
C54364 OR2X1_LOC_765/Y OR2X1_LOC_52/B 0.02fF
C54365 VDD OR2X1_LOC_6/A 1.48fF
C54366 OR2X1_LOC_496/Y OR2X1_LOC_40/Y 0.06fF
C54367 AND2X1_LOC_797/A AND2X1_LOC_213/B 0.12fF
C54368 OR2X1_LOC_100/Y OR2X1_LOC_608/a_8_216# 0.03fF
C54369 OR2X1_LOC_382/Y OR2X1_LOC_427/A 0.00fF
C54370 OR2X1_LOC_94/a_8_216# OR2X1_LOC_56/A 0.02fF
C54371 AND2X1_LOC_339/B OR2X1_LOC_743/A 0.03fF
C54372 OR2X1_LOC_189/Y AND2X1_LOC_476/Y 1.49fF
C54373 OR2X1_LOC_168/a_8_216# OR2X1_LOC_756/B 0.01fF
C54374 OR2X1_LOC_185/A AND2X1_LOC_529/a_8_24# 0.04fF
C54375 AND2X1_LOC_64/Y OR2X1_LOC_113/A 0.01fF
C54376 OR2X1_LOC_193/A OR2X1_LOC_161/B 0.18fF
C54377 OR2X1_LOC_106/A AND2X1_LOC_243/Y 0.02fF
C54378 AND2X1_LOC_569/A VDD 0.51fF
C54379 AND2X1_LOC_729/B OR2X1_LOC_12/Y 0.00fF
C54380 OR2X1_LOC_702/A OR2X1_LOC_596/A 0.00fF
C54381 AND2X1_LOC_707/Y AND2X1_LOC_687/A 0.03fF
C54382 OR2X1_LOC_256/Y OR2X1_LOC_625/Y 0.38fF
C54383 OR2X1_LOC_678/Y AND2X1_LOC_43/B 0.03fF
C54384 OR2X1_LOC_185/Y OR2X1_LOC_809/B 1.02fF
C54385 OR2X1_LOC_756/B AND2X1_LOC_617/a_8_24# 0.03fF
C54386 AND2X1_LOC_721/Y AND2X1_LOC_465/Y 0.02fF
C54387 OR2X1_LOC_8/Y OR2X1_LOC_26/Y 0.05fF
C54388 AND2X1_LOC_500/a_8_24# AND2X1_LOC_570/Y 0.01fF
C54389 OR2X1_LOC_160/A OR2X1_LOC_663/A 0.01fF
C54390 AND2X1_LOC_367/A AND2X1_LOC_318/a_8_24# 0.18fF
C54391 OR2X1_LOC_151/A OR2X1_LOC_476/Y 0.10fF
C54392 OR2X1_LOC_106/Y OR2X1_LOC_71/Y 0.02fF
C54393 OR2X1_LOC_100/Y OR2X1_LOC_185/A 0.06fF
C54394 AND2X1_LOC_95/Y OR2X1_LOC_475/B 0.03fF
C54395 OR2X1_LOC_329/B OR2X1_LOC_36/Y 0.06fF
C54396 OR2X1_LOC_290/a_8_216# OR2X1_LOC_316/Y 0.01fF
C54397 AND2X1_LOC_773/Y OR2X1_LOC_46/A 0.01fF
C54398 OR2X1_LOC_714/Y OR2X1_LOC_724/a_8_216# 0.39fF
C54399 OR2X1_LOC_604/A OR2X1_LOC_3/Y 0.09fF
C54400 OR2X1_LOC_319/a_8_216# OR2X1_LOC_856/B 0.03fF
C54401 OR2X1_LOC_312/Y OR2X1_LOC_51/Y 0.03fF
C54402 AND2X1_LOC_547/Y AND2X1_LOC_475/a_36_24# 0.00fF
C54403 OR2X1_LOC_235/B OR2X1_LOC_87/A 0.03fF
C54404 AND2X1_LOC_191/Y AND2X1_LOC_731/Y 0.03fF
C54405 AND2X1_LOC_845/Y AND2X1_LOC_287/B 0.01fF
C54406 OR2X1_LOC_254/B AND2X1_LOC_253/a_8_24# 0.01fF
C54407 OR2X1_LOC_449/B OR2X1_LOC_78/B 0.06fF
C54408 OR2X1_LOC_634/A AND2X1_LOC_56/B 0.02fF
C54409 OR2X1_LOC_653/Y OR2X1_LOC_405/a_8_216# 0.03fF
C54410 OR2X1_LOC_592/a_8_216# OR2X1_LOC_78/A 0.01fF
C54411 OR2X1_LOC_665/Y OR2X1_LOC_56/A 0.07fF
C54412 OR2X1_LOC_429/Y OR2X1_LOC_582/a_36_216# 0.01fF
C54413 AND2X1_LOC_40/Y OR2X1_LOC_652/a_8_216# 0.01fF
C54414 AND2X1_LOC_190/a_8_24# OR2X1_LOC_529/Y 0.00fF
C54415 AND2X1_LOC_231/Y D_INPUT_0 0.02fF
C54416 OR2X1_LOC_621/B AND2X1_LOC_670/a_8_24# 0.04fF
C54417 OR2X1_LOC_814/A AND2X1_LOC_488/a_8_24# 0.01fF
C54418 OR2X1_LOC_600/A AND2X1_LOC_345/Y 0.03fF
C54419 OR2X1_LOC_3/Y OR2X1_LOC_66/A 0.03fF
C54420 OR2X1_LOC_147/B OR2X1_LOC_738/A 0.02fF
C54421 AND2X1_LOC_711/Y AND2X1_LOC_731/Y 0.00fF
C54422 OR2X1_LOC_856/B OR2X1_LOC_377/A 0.02fF
C54423 AND2X1_LOC_738/B OR2X1_LOC_485/A 0.01fF
C54424 AND2X1_LOC_339/B OR2X1_LOC_246/A 0.03fF
C54425 AND2X1_LOC_364/a_8_24# D_INPUT_0 0.01fF
C54426 OR2X1_LOC_7/A AND2X1_LOC_434/Y 0.79fF
C54427 OR2X1_LOC_485/A OR2X1_LOC_56/A 0.22fF
C54428 AND2X1_LOC_208/B OR2X1_LOC_6/A 0.01fF
C54429 OR2X1_LOC_812/B OR2X1_LOC_812/A 0.06fF
C54430 OR2X1_LOC_634/A AND2X1_LOC_8/Y 0.02fF
C54431 D_INPUT_0 OR2X1_LOC_161/B 0.02fF
C54432 OR2X1_LOC_31/Y OR2X1_LOC_18/a_8_216# 0.10fF
C54433 AND2X1_LOC_568/B AND2X1_LOC_798/Y 0.81fF
C54434 INPUT_5 OR2X1_LOC_752/a_8_216# 0.02fF
C54435 INPUT_0 OR2X1_LOC_24/Y 0.07fF
C54436 OR2X1_LOC_833/B OR2X1_LOC_203/a_8_216# 0.01fF
C54437 OR2X1_LOC_589/A AND2X1_LOC_633/Y 0.02fF
C54438 OR2X1_LOC_648/B OR2X1_LOC_19/B 0.03fF
C54439 AND2X1_LOC_357/A AND2X1_LOC_514/Y 0.01fF
C54440 OR2X1_LOC_377/A OR2X1_LOC_793/a_8_216# 0.14fF
C54441 AND2X1_LOC_70/Y AND2X1_LOC_666/a_8_24# 0.03fF
C54442 AND2X1_LOC_512/Y AND2X1_LOC_356/B 0.06fF
C54443 AND2X1_LOC_810/A AND2X1_LOC_170/B 0.05fF
C54444 OR2X1_LOC_589/A D_INPUT_0 0.02fF
C54445 OR2X1_LOC_427/A OR2X1_LOC_591/A 0.01fF
C54446 AND2X1_LOC_154/a_8_24# OR2X1_LOC_39/A 0.01fF
C54447 AND2X1_LOC_559/a_8_24# AND2X1_LOC_520/Y 0.11fF
C54448 AND2X1_LOC_81/B OR2X1_LOC_624/A 0.05fF
C54449 OR2X1_LOC_433/a_8_216# OR2X1_LOC_48/B 0.02fF
C54450 AND2X1_LOC_715/A AND2X1_LOC_727/A 0.03fF
C54451 AND2X1_LOC_523/a_8_24# OR2X1_LOC_271/Y 0.01fF
C54452 OR2X1_LOC_624/A OR2X1_LOC_358/B 0.03fF
C54453 AND2X1_LOC_76/Y OR2X1_LOC_26/Y 0.00fF
C54454 OR2X1_LOC_663/A OR2X1_LOC_624/B 0.00fF
C54455 OR2X1_LOC_364/A OR2X1_LOC_160/A 0.07fF
C54456 AND2X1_LOC_144/a_36_24# OR2X1_LOC_705/Y 0.00fF
C54457 OR2X1_LOC_476/a_8_216# AND2X1_LOC_92/Y 0.04fF
C54458 INPUT_0 AND2X1_LOC_855/a_8_24# 0.01fF
C54459 OR2X1_LOC_185/Y OR2X1_LOC_160/A 0.24fF
C54460 OR2X1_LOC_315/Y OR2X1_LOC_6/A 0.25fF
C54461 OR2X1_LOC_692/Y AND2X1_LOC_648/B 0.04fF
C54462 OR2X1_LOC_121/B OR2X1_LOC_78/B 0.05fF
C54463 OR2X1_LOC_140/B OR2X1_LOC_140/a_36_216# 0.02fF
C54464 AND2X1_LOC_76/Y OR2X1_LOC_89/A 0.09fF
C54465 OR2X1_LOC_343/B OR2X1_LOC_343/a_8_216# 0.47fF
C54466 AND2X1_LOC_12/Y OR2X1_LOC_864/A 0.03fF
C54467 AND2X1_LOC_362/B D_INPUT_3 2.27fF
C54468 OR2X1_LOC_32/B AND2X1_LOC_852/Y 0.07fF
C54469 AND2X1_LOC_53/Y OR2X1_LOC_66/A 0.07fF
C54470 AND2X1_LOC_453/Y OR2X1_LOC_52/B 0.08fF
C54471 OR2X1_LOC_848/A OR2X1_LOC_772/a_8_216# 0.02fF
C54472 AND2X1_LOC_392/A OR2X1_LOC_31/Y 0.03fF
C54473 AND2X1_LOC_274/a_36_24# OR2X1_LOC_52/B 0.01fF
C54474 AND2X1_LOC_12/Y OR2X1_LOC_774/Y 2.67fF
C54475 OR2X1_LOC_375/A OR2X1_LOC_449/B 0.03fF
C54476 OR2X1_LOC_40/Y AND2X1_LOC_851/B 0.00fF
C54477 AND2X1_LOC_191/Y OR2X1_LOC_18/Y 7.44fF
C54478 AND2X1_LOC_42/B OR2X1_LOC_847/A 0.00fF
C54479 AND2X1_LOC_40/Y OR2X1_LOC_456/A 0.14fF
C54480 OR2X1_LOC_154/A OR2X1_LOC_389/B 0.14fF
C54481 OR2X1_LOC_70/Y OR2X1_LOC_48/B 0.17fF
C54482 AND2X1_LOC_512/Y OR2X1_LOC_22/Y 0.11fF
C54483 VDD D_INPUT_2 0.26fF
C54484 OR2X1_LOC_121/B OR2X1_LOC_721/Y 0.11fF
C54485 AND2X1_LOC_711/Y OR2X1_LOC_18/Y 0.03fF
C54486 VDD AND2X1_LOC_139/A -0.00fF
C54487 AND2X1_LOC_156/a_8_24# OR2X1_LOC_619/Y 0.01fF
C54488 OR2X1_LOC_70/Y OR2X1_LOC_18/Y 0.72fF
C54489 OR2X1_LOC_242/a_36_216# OR2X1_LOC_532/B 0.00fF
C54490 AND2X1_LOC_47/Y OR2X1_LOC_778/B 0.03fF
C54491 OR2X1_LOC_26/Y AND2X1_LOC_374/Y 0.01fF
C54492 OR2X1_LOC_41/a_8_216# OR2X1_LOC_13/Y 0.01fF
C54493 AND2X1_LOC_851/a_8_24# OR2X1_LOC_95/Y 0.04fF
C54494 OR2X1_LOC_481/A AND2X1_LOC_847/Y 0.01fF
C54495 AND2X1_LOC_810/Y AND2X1_LOC_469/B 0.01fF
C54496 VDD GATE_479 0.22fF
C54497 AND2X1_LOC_217/a_36_24# AND2X1_LOC_772/Y 0.01fF
C54498 AND2X1_LOC_1/Y AND2X1_LOC_22/a_36_24# 0.00fF
C54499 AND2X1_LOC_12/Y AND2X1_LOC_281/a_8_24# 0.01fF
C54500 OR2X1_LOC_26/Y OR2X1_LOC_52/B 0.19fF
C54501 OR2X1_LOC_488/a_36_216# AND2X1_LOC_573/A -0.01fF
C54502 OR2X1_LOC_672/Y OR2X1_LOC_26/Y 0.00fF
C54503 OR2X1_LOC_841/A OR2X1_LOC_223/A 0.16fF
C54504 AND2X1_LOC_484/a_8_24# OR2X1_LOC_738/A 0.04fF
C54505 OR2X1_LOC_294/Y OR2X1_LOC_675/Y 0.02fF
C54506 AND2X1_LOC_514/Y OR2X1_LOC_48/B 0.03fF
C54507 OR2X1_LOC_419/Y AND2X1_LOC_477/Y 0.06fF
C54508 VDD OR2X1_LOC_289/a_8_216# 0.21fF
C54509 AND2X1_LOC_721/A AND2X1_LOC_860/A 0.04fF
C54510 OR2X1_LOC_64/Y OR2X1_LOC_118/Y 0.03fF
C54511 OR2X1_LOC_215/A OR2X1_LOC_215/Y 0.01fF
C54512 OR2X1_LOC_351/B OR2X1_LOC_351/a_8_216# 0.03fF
C54513 AND2X1_LOC_489/Y OR2X1_LOC_26/Y 0.02fF
C54514 VDD AND2X1_LOC_463/B 0.09fF
C54515 OR2X1_LOC_490/Y AND2X1_LOC_361/A 0.01fF
C54516 OR2X1_LOC_756/B OR2X1_LOC_440/A 0.04fF
C54517 OR2X1_LOC_89/A OR2X1_LOC_52/B 0.14fF
C54518 AND2X1_LOC_7/B OR2X1_LOC_181/A 0.11fF
C54519 OR2X1_LOC_852/B OR2X1_LOC_852/A 0.12fF
C54520 AND2X1_LOC_70/Y OR2X1_LOC_247/a_8_216# 0.01fF
C54521 OR2X1_LOC_533/Y OR2X1_LOC_534/Y 0.18fF
C54522 OR2X1_LOC_121/B OR2X1_LOC_375/A 0.30fF
C54523 OR2X1_LOC_859/A OR2X1_LOC_571/B 0.01fF
C54524 AND2X1_LOC_620/Y OR2X1_LOC_59/Y 0.03fF
C54525 OR2X1_LOC_461/B OR2X1_LOC_598/A 0.02fF
C54526 OR2X1_LOC_549/a_36_216# D_GATE_366 0.00fF
C54527 AND2X1_LOC_489/Y OR2X1_LOC_89/A 1.15fF
C54528 OR2X1_LOC_502/A OR2X1_LOC_468/a_8_216# 0.05fF
C54529 AND2X1_LOC_211/B AND2X1_LOC_211/a_8_24# 0.03fF
C54530 OR2X1_LOC_136/Y OR2X1_LOC_13/B 0.06fF
C54531 OR2X1_LOC_409/B OR2X1_LOC_586/a_8_216# 0.47fF
C54532 AND2X1_LOC_536/a_8_24# D_INPUT_0 0.02fF
C54533 OR2X1_LOC_160/B OR2X1_LOC_358/A 0.19fF
C54534 OR2X1_LOC_288/a_8_216# OR2X1_LOC_286/B 0.01fF
C54535 OR2X1_LOC_497/Y AND2X1_LOC_842/B 0.03fF
C54536 OR2X1_LOC_417/A AND2X1_LOC_643/a_36_24# 0.00fF
C54537 OR2X1_LOC_9/Y OR2X1_LOC_68/B 0.10fF
C54538 OR2X1_LOC_476/B OR2X1_LOC_87/B 0.08fF
C54539 OR2X1_LOC_185/A OR2X1_LOC_532/B 0.17fF
C54540 OR2X1_LOC_504/Y OR2X1_LOC_18/Y 0.01fF
C54541 AND2X1_LOC_31/Y OR2X1_LOC_182/B 0.03fF
C54542 OR2X1_LOC_70/Y OR2X1_LOC_385/Y 0.06fF
C54543 OR2X1_LOC_362/A OR2X1_LOC_68/B 0.48fF
C54544 OR2X1_LOC_262/Y OR2X1_LOC_64/Y 0.00fF
C54545 OR2X1_LOC_501/B AND2X1_LOC_72/B 0.03fF
C54546 OR2X1_LOC_329/B OR2X1_LOC_419/Y 0.10fF
C54547 OR2X1_LOC_59/Y AND2X1_LOC_215/A 0.01fF
C54548 OR2X1_LOC_650/Y OR2X1_LOC_87/B 0.07fF
C54549 OR2X1_LOC_331/A OR2X1_LOC_331/a_8_216# 0.04fF
C54550 AND2X1_LOC_450/a_8_24# AND2X1_LOC_450/Y 0.01fF
C54551 OR2X1_LOC_3/a_8_216# OR2X1_LOC_17/Y 0.02fF
C54552 OR2X1_LOC_97/A OR2X1_LOC_788/B 0.00fF
C54553 OR2X1_LOC_16/A OR2X1_LOC_536/a_8_216# 0.01fF
C54554 OR2X1_LOC_755/A OR2X1_LOC_89/A 0.01fF
C54555 AND2X1_LOC_560/a_8_24# OR2X1_LOC_696/A 0.01fF
C54556 OR2X1_LOC_64/Y OR2X1_LOC_238/Y 0.03fF
C54557 AND2X1_LOC_56/B OR2X1_LOC_335/B 0.03fF
C54558 OR2X1_LOC_696/a_8_216# OR2X1_LOC_696/Y -0.00fF
C54559 AND2X1_LOC_587/a_8_24# INPUT_6 0.01fF
C54560 OR2X1_LOC_673/Y OR2X1_LOC_720/B 0.00fF
C54561 OR2X1_LOC_497/a_8_216# OR2X1_LOC_71/Y 0.01fF
C54562 AND2X1_LOC_46/a_8_24# AND2X1_LOC_42/B 0.01fF
C54563 AND2X1_LOC_459/Y OR2X1_LOC_408/Y 0.15fF
C54564 OR2X1_LOC_43/A D_INPUT_0 13.82fF
C54565 OR2X1_LOC_777/B OR2X1_LOC_356/A 0.21fF
C54566 OR2X1_LOC_624/A OR2X1_LOC_112/B 0.01fF
C54567 OR2X1_LOC_476/B OR2X1_LOC_33/B 0.02fF
C54568 OR2X1_LOC_516/Y AND2X1_LOC_721/Y 0.03fF
C54569 OR2X1_LOC_354/A OR2X1_LOC_365/B 0.00fF
C54570 OR2X1_LOC_249/Y OR2X1_LOC_343/B 0.01fF
C54571 OR2X1_LOC_605/B OR2X1_LOC_121/B 0.00fF
C54572 OR2X1_LOC_18/Y OR2X1_LOC_184/Y 0.54fF
C54573 OR2X1_LOC_168/B AND2X1_LOC_31/Y 0.08fF
C54574 OR2X1_LOC_249/a_8_216# D_INPUT_1 0.06fF
C54575 OR2X1_LOC_437/Y OR2X1_LOC_48/B 0.07fF
C54576 AND2X1_LOC_390/B AND2X1_LOC_537/Y 0.04fF
C54577 AND2X1_LOC_64/Y AND2X1_LOC_91/B 2.78fF
C54578 OR2X1_LOC_22/Y OR2X1_LOC_279/a_8_216# 0.04fF
C54579 OR2X1_LOC_518/Y AND2X1_LOC_520/a_8_24# 0.01fF
C54580 OR2X1_LOC_95/Y OR2X1_LOC_753/A 0.07fF
C54581 OR2X1_LOC_76/Y OR2X1_LOC_440/A 0.00fF
C54582 OR2X1_LOC_62/B OR2X1_LOC_629/a_8_216# 0.01fF
C54583 AND2X1_LOC_543/Y AND2X1_LOC_552/a_8_24# 0.02fF
C54584 OR2X1_LOC_17/Y AND2X1_LOC_639/A 0.29fF
C54585 OR2X1_LOC_36/Y OR2X1_LOC_618/Y 0.10fF
C54586 OR2X1_LOC_792/Y OR2X1_LOC_580/a_8_216# 0.02fF
C54587 OR2X1_LOC_417/A OR2X1_LOC_238/Y 0.08fF
C54588 OR2X1_LOC_18/Y AND2X1_LOC_641/a_8_24# 0.01fF
C54589 OR2X1_LOC_277/a_8_216# OR2X1_LOC_278/A 0.01fF
C54590 OR2X1_LOC_624/A OR2X1_LOC_66/Y 0.07fF
C54591 OR2X1_LOC_634/a_36_216# OR2X1_LOC_68/B 0.00fF
C54592 AND2X1_LOC_752/a_8_24# AND2X1_LOC_31/Y 0.01fF
C54593 OR2X1_LOC_51/Y OR2X1_LOC_13/B 0.34fF
C54594 OR2X1_LOC_744/A OR2X1_LOC_589/Y 0.01fF
C54595 OR2X1_LOC_147/A OR2X1_LOC_705/a_8_216# 0.01fF
C54596 OR2X1_LOC_70/A OR2X1_LOC_48/B 0.00fF
C54597 OR2X1_LOC_426/B OR2X1_LOC_300/Y 0.09fF
C54598 AND2X1_LOC_43/B OR2X1_LOC_378/a_8_216# 0.08fF
C54599 OR2X1_LOC_516/Y OR2X1_LOC_482/Y 0.15fF
C54600 AND2X1_LOC_851/B OR2X1_LOC_7/A 0.07fF
C54601 AND2X1_LOC_12/Y OR2X1_LOC_351/a_8_216# 0.01fF
C54602 AND2X1_LOC_316/a_36_24# OR2X1_LOC_68/B 0.00fF
C54603 OR2X1_LOC_18/Y OR2X1_LOC_70/A 0.03fF
C54604 OR2X1_LOC_100/a_8_216# OR2X1_LOC_608/Y 0.39fF
C54605 OR2X1_LOC_594/Y OR2X1_LOC_533/A 0.00fF
C54606 AND2X1_LOC_810/a_36_24# AND2X1_LOC_661/A 0.00fF
C54607 OR2X1_LOC_6/A OR2X1_LOC_67/Y 0.01fF
C54608 AND2X1_LOC_465/Y AND2X1_LOC_471/a_8_24# 0.11fF
C54609 OR2X1_LOC_97/A AND2X1_LOC_22/Y 0.07fF
C54610 OR2X1_LOC_61/A AND2X1_LOC_7/B 0.01fF
C54611 OR2X1_LOC_549/a_8_216# OR2X1_LOC_549/A 0.02fF
C54612 OR2X1_LOC_486/Y OR2X1_LOC_562/A 0.01fF
C54613 OR2X1_LOC_74/A AND2X1_LOC_675/a_8_24# 0.08fF
C54614 AND2X1_LOC_47/Y OR2X1_LOC_99/B 0.14fF
C54615 OR2X1_LOC_223/A OR2X1_LOC_794/a_36_216# 0.00fF
C54616 OR2X1_LOC_114/B OR2X1_LOC_501/A 0.01fF
C54617 OR2X1_LOC_725/B OR2X1_LOC_725/a_8_216# 0.05fF
C54618 OR2X1_LOC_651/A AND2X1_LOC_51/Y 0.02fF
C54619 AND2X1_LOC_539/Y OR2X1_LOC_589/A 0.03fF
C54620 AND2X1_LOC_804/a_8_24# OR2X1_LOC_52/B 0.01fF
C54621 AND2X1_LOC_59/Y AND2X1_LOC_31/Y 5.22fF
C54622 OR2X1_LOC_26/Y AND2X1_LOC_216/A 0.02fF
C54623 OR2X1_LOC_715/A AND2X1_LOC_36/Y 0.43fF
C54624 OR2X1_LOC_16/A AND2X1_LOC_214/a_8_24# 0.01fF
C54625 AND2X1_LOC_117/a_8_24# OR2X1_LOC_786/Y 0.01fF
C54626 AND2X1_LOC_711/Y AND2X1_LOC_620/Y 0.01fF
C54627 OR2X1_LOC_501/B AND2X1_LOC_36/Y 0.01fF
C54628 OR2X1_LOC_151/A OR2X1_LOC_563/A 0.39fF
C54629 OR2X1_LOC_532/B OR2X1_LOC_750/a_36_216# 0.00fF
C54630 AND2X1_LOC_438/a_8_24# OR2X1_LOC_161/B 0.01fF
C54631 OR2X1_LOC_74/A AND2X1_LOC_795/Y 0.00fF
C54632 OR2X1_LOC_235/B OR2X1_LOC_844/B 0.00fF
C54633 AND2X1_LOC_259/Y AND2X1_LOC_848/A 0.07fF
C54634 OR2X1_LOC_416/Y AND2X1_LOC_660/A 0.07fF
C54635 OR2X1_LOC_405/Y AND2X1_LOC_406/a_8_24# 0.00fF
C54636 OR2X1_LOC_89/A AND2X1_LOC_216/A 0.16fF
C54637 OR2X1_LOC_219/B OR2X1_LOC_358/A 0.07fF
C54638 OR2X1_LOC_45/B OR2X1_LOC_528/a_8_216# 0.06fF
C54639 OR2X1_LOC_600/A AND2X1_LOC_465/A 0.04fF
C54640 OR2X1_LOC_44/Y AND2X1_LOC_657/A 0.22fF
C54641 OR2X1_LOC_696/A OR2X1_LOC_122/a_36_216# 0.02fF
C54642 OR2X1_LOC_736/Y OR2X1_LOC_294/Y 0.08fF
C54643 OR2X1_LOC_443/a_8_216# AND2X1_LOC_47/Y 0.01fF
C54644 OR2X1_LOC_95/Y AND2X1_LOC_845/Y 2.23fF
C54645 OR2X1_LOC_61/Y OR2X1_LOC_339/A 0.18fF
C54646 OR2X1_LOC_106/Y OR2X1_LOC_426/B 0.02fF
C54647 AND2X1_LOC_388/Y OR2X1_LOC_533/Y 0.28fF
C54648 OR2X1_LOC_598/Y OR2X1_LOC_161/B 0.05fF
C54649 OR2X1_LOC_147/B AND2X1_LOC_36/Y 0.10fF
C54650 OR2X1_LOC_446/Y OR2X1_LOC_783/A 0.03fF
C54651 AND2X1_LOC_593/a_8_24# OR2X1_LOC_12/Y 0.04fF
C54652 OR2X1_LOC_502/A OR2X1_LOC_508/Y 0.00fF
C54653 AND2X1_LOC_858/B AND2X1_LOC_241/a_8_24# 0.04fF
C54654 AND2X1_LOC_227/Y OR2X1_LOC_72/a_36_216# 0.01fF
C54655 OR2X1_LOC_680/A OR2X1_LOC_13/B 0.36fF
C54656 AND2X1_LOC_550/A OR2X1_LOC_142/Y 1.04fF
C54657 OR2X1_LOC_688/Y AND2X1_LOC_31/Y 0.11fF
C54658 OR2X1_LOC_589/A OR2X1_LOC_131/A 0.03fF
C54659 OR2X1_LOC_404/Y AND2X1_LOC_497/a_36_24# 0.01fF
C54660 AND2X1_LOC_433/a_8_24# AND2X1_LOC_18/Y 0.01fF
C54661 AND2X1_LOC_847/Y AND2X1_LOC_789/Y 0.02fF
C54662 AND2X1_LOC_51/Y OR2X1_LOC_728/B 0.22fF
C54663 AND2X1_LOC_362/a_8_24# AND2X1_LOC_284/a_8_24# 0.23fF
C54664 OR2X1_LOC_585/A OR2X1_LOC_71/A 0.10fF
C54665 OR2X1_LOC_133/a_36_216# OR2X1_LOC_604/A 0.01fF
C54666 AND2X1_LOC_520/a_8_24# OR2X1_LOC_91/A 0.01fF
C54667 AND2X1_LOC_340/Y OR2X1_LOC_59/Y 7.74fF
C54668 OR2X1_LOC_379/Y OR2X1_LOC_598/a_36_216# 0.00fF
C54669 AND2X1_LOC_474/A OR2X1_LOC_428/A 0.02fF
C54670 OR2X1_LOC_696/A AND2X1_LOC_809/A 0.02fF
C54671 OR2X1_LOC_421/a_8_216# OR2X1_LOC_428/A 0.01fF
C54672 OR2X1_LOC_335/Y OR2X1_LOC_161/B 0.02fF
C54673 OR2X1_LOC_177/Y OR2X1_LOC_329/B 0.00fF
C54674 AND2X1_LOC_474/A OR2X1_LOC_595/A 0.03fF
C54675 OR2X1_LOC_154/A OR2X1_LOC_714/a_8_216# 0.04fF
C54676 OR2X1_LOC_777/a_8_216# OR2X1_LOC_66/A 0.01fF
C54677 AND2X1_LOC_181/Y OR2X1_LOC_59/Y 0.01fF
C54678 AND2X1_LOC_571/A AND2X1_LOC_573/A 0.01fF
C54679 OR2X1_LOC_6/A AND2X1_LOC_269/a_8_24# 0.01fF
C54680 AND2X1_LOC_64/Y AND2X1_LOC_72/Y 0.01fF
C54681 AND2X1_LOC_64/Y OR2X1_LOC_799/A 4.36fF
C54682 OR2X1_LOC_743/A OR2X1_LOC_300/Y 0.12fF
C54683 AND2X1_LOC_181/a_8_24# OR2X1_LOC_158/A 0.02fF
C54684 OR2X1_LOC_494/A OR2X1_LOC_427/A 0.03fF
C54685 AND2X1_LOC_715/Y AND2X1_LOC_809/A 0.02fF
C54686 AND2X1_LOC_40/Y OR2X1_LOC_161/B 0.35fF
C54687 OR2X1_LOC_185/Y OR2X1_LOC_130/Y 0.09fF
C54688 OR2X1_LOC_276/a_8_216# OR2X1_LOC_66/Y 0.00fF
C54689 OR2X1_LOC_243/B OR2X1_LOC_68/B 0.05fF
C54690 OR2X1_LOC_850/a_8_216# OR2X1_LOC_349/A 0.01fF
C54691 OR2X1_LOC_175/Y AND2X1_LOC_95/Y 0.14fF
C54692 AND2X1_LOC_799/a_8_24# OR2X1_LOC_619/Y 0.03fF
C54693 AND2X1_LOC_564/B AND2X1_LOC_621/Y 0.07fF
C54694 AND2X1_LOC_539/Y AND2X1_LOC_365/A 0.01fF
C54695 OR2X1_LOC_188/a_8_216# AND2X1_LOC_43/B 0.06fF
C54696 OR2X1_LOC_604/A OR2X1_LOC_329/B 0.10fF
C54697 OR2X1_LOC_40/Y AND2X1_LOC_364/Y 0.01fF
C54698 OR2X1_LOC_663/A OR2X1_LOC_768/a_8_216# 0.02fF
C54699 OR2X1_LOC_40/Y OR2X1_LOC_674/a_8_216# 0.02fF
C54700 AND2X1_LOC_130/a_8_24# OR2X1_LOC_517/A 0.04fF
C54701 AND2X1_LOC_387/B AND2X1_LOC_36/Y 0.06fF
C54702 OR2X1_LOC_619/Y OR2X1_LOC_158/Y 0.01fF
C54703 OR2X1_LOC_87/A AND2X1_LOC_226/a_8_24# 0.02fF
C54704 AND2X1_LOC_95/Y OR2X1_LOC_691/Y 0.09fF
C54705 OR2X1_LOC_291/a_8_216# OR2X1_LOC_16/A 0.11fF
C54706 OR2X1_LOC_51/Y AND2X1_LOC_508/a_36_24# 0.01fF
C54707 OR2X1_LOC_30/a_8_216# INPUT_7 0.01fF
C54708 OR2X1_LOC_485/Y AND2X1_LOC_512/Y 0.16fF
C54709 OR2X1_LOC_844/a_8_216# OR2X1_LOC_844/B 0.07fF
C54710 OR2X1_LOC_600/A AND2X1_LOC_477/a_8_24# 0.01fF
C54711 OR2X1_LOC_509/a_8_216# OR2X1_LOC_502/A 0.01fF
C54712 OR2X1_LOC_710/B AND2X1_LOC_144/a_36_24# 0.00fF
C54713 OR2X1_LOC_479/Y OR2X1_LOC_776/A 0.00fF
C54714 AND2X1_LOC_484/a_8_24# AND2X1_LOC_36/Y 0.01fF
C54715 AND2X1_LOC_539/Y OR2X1_LOC_43/A 0.07fF
C54716 OR2X1_LOC_246/A OR2X1_LOC_300/Y 0.03fF
C54717 OR2X1_LOC_659/B OR2X1_LOC_267/Y 0.09fF
C54718 OR2X1_LOC_186/Y OR2X1_LOC_161/A 0.36fF
C54719 AND2X1_LOC_776/a_8_24# OR2X1_LOC_164/Y 0.01fF
C54720 VDD OR2X1_LOC_216/A 0.19fF
C54721 AND2X1_LOC_357/A AND2X1_LOC_357/a_8_24# 0.07fF
C54722 OR2X1_LOC_85/A OR2X1_LOC_428/A 0.07fF
C54723 OR2X1_LOC_634/A AND2X1_LOC_92/Y 0.02fF
C54724 OR2X1_LOC_494/A AND2X1_LOC_363/A 0.40fF
C54725 GATE_811 OR2X1_LOC_152/A 0.25fF
C54726 AND2X1_LOC_753/B AND2X1_LOC_18/Y 0.33fF
C54727 OR2X1_LOC_814/A OR2X1_LOC_571/Y 0.01fF
C54728 OR2X1_LOC_502/A OR2X1_LOC_66/A 0.28fF
C54729 OR2X1_LOC_31/Y OR2X1_LOC_589/Y 0.01fF
C54730 VDD OR2X1_LOC_485/a_8_216# 0.21fF
C54731 AND2X1_LOC_357/B AND2X1_LOC_357/a_36_24# 0.01fF
C54732 AND2X1_LOC_365/a_36_24# OR2X1_LOC_744/A 0.01fF
C54733 OR2X1_LOC_841/A OR2X1_LOC_502/A 0.01fF
C54734 OR2X1_LOC_690/A AND2X1_LOC_208/Y 0.63fF
C54735 OR2X1_LOC_45/B OR2X1_LOC_682/a_8_216# 0.02fF
C54736 AND2X1_LOC_360/a_8_24# OR2X1_LOC_56/A 0.02fF
C54737 OR2X1_LOC_348/Y OR2X1_LOC_811/A 0.10fF
C54738 AND2X1_LOC_31/Y OR2X1_LOC_733/Y 0.01fF
C54739 OR2X1_LOC_85/A OR2X1_LOC_595/A 0.44fF
C54740 OR2X1_LOC_405/A AND2X1_LOC_371/a_8_24# 0.01fF
C54741 OR2X1_LOC_364/B OR2X1_LOC_87/A 0.01fF
C54742 OR2X1_LOC_758/Y OR2X1_LOC_792/Y 0.01fF
C54743 OR2X1_LOC_65/B OR2X1_LOC_131/a_8_216# 0.01fF
C54744 OR2X1_LOC_715/B OR2X1_LOC_539/Y 0.41fF
C54745 OR2X1_LOC_78/A OR2X1_LOC_712/a_8_216# 0.01fF
C54746 OR2X1_LOC_405/A AND2X1_LOC_18/Y 0.13fF
C54747 AND2X1_LOC_364/a_36_24# OR2X1_LOC_43/A 0.00fF
C54748 OR2X1_LOC_528/Y OR2X1_LOC_39/A 0.04fF
C54749 OR2X1_LOC_160/B OR2X1_LOC_796/a_8_216# 0.01fF
C54750 AND2X1_LOC_264/a_8_24# OR2X1_LOC_12/Y 0.04fF
C54751 AND2X1_LOC_8/Y OR2X1_LOC_633/A 0.42fF
C54752 VDD OR2X1_LOC_362/B 0.00fF
C54753 OR2X1_LOC_91/A OR2X1_LOC_92/Y 0.64fF
C54754 OR2X1_LOC_571/B OR2X1_LOC_66/A 0.01fF
C54755 OR2X1_LOC_545/B AND2X1_LOC_36/Y 0.03fF
C54756 OR2X1_LOC_113/a_8_216# AND2X1_LOC_42/B 0.01fF
C54757 VDD OR2X1_LOC_45/a_8_216# 0.00fF
C54758 OR2X1_LOC_821/Y OR2X1_LOC_753/A 0.02fF
C54759 AND2X1_LOC_658/B OR2X1_LOC_18/Y 0.03fF
C54760 OR2X1_LOC_45/B OR2X1_LOC_609/a_8_216# 0.40fF
C54761 AND2X1_LOC_571/a_36_24# AND2X1_LOC_489/Y 0.00fF
C54762 VDD AND2X1_LOC_403/B 0.04fF
C54763 OR2X1_LOC_701/Y VDD 0.08fF
C54764 VDD OR2X1_LOC_499/a_8_216# 0.00fF
C54765 OR2X1_LOC_154/A OR2X1_LOC_6/B 0.10fF
C54766 OR2X1_LOC_856/B OR2X1_LOC_78/B 0.07fF
C54767 AND2X1_LOC_784/A AND2X1_LOC_212/A 0.02fF
C54768 OR2X1_LOC_275/Y AND2X1_LOC_276/a_8_24# 0.05fF
C54769 OR2X1_LOC_756/B OR2X1_LOC_436/B 0.01fF
C54770 AND2X1_LOC_40/Y OR2X1_LOC_435/B 0.00fF
C54771 OR2X1_LOC_673/a_8_216# AND2X1_LOC_8/Y 0.01fF
C54772 OR2X1_LOC_600/A OR2X1_LOC_237/Y 0.03fF
C54773 AND2X1_LOC_51/Y OR2X1_LOC_338/A 0.17fF
C54774 AND2X1_LOC_22/Y OR2X1_LOC_605/a_8_216# 0.01fF
C54775 AND2X1_LOC_362/B AND2X1_LOC_806/A 0.04fF
C54776 AND2X1_LOC_310/a_8_24# OR2X1_LOC_161/A 0.17fF
C54777 AND2X1_LOC_797/a_8_24# AND2X1_LOC_192/Y 0.02fF
C54778 OR2X1_LOC_400/A OR2X1_LOC_66/A 0.01fF
C54779 OR2X1_LOC_468/Y OR2X1_LOC_302/A 0.03fF
C54780 AND2X1_LOC_215/Y OR2X1_LOC_85/A 0.01fF
C54781 OR2X1_LOC_512/A OR2X1_LOC_308/a_8_216# 0.07fF
C54782 OR2X1_LOC_9/Y AND2X1_LOC_673/a_8_24# 0.11fF
C54783 AND2X1_LOC_340/Y OR2X1_LOC_70/Y 0.03fF
C54784 AND2X1_LOC_568/a_8_24# AND2X1_LOC_212/Y 0.02fF
C54785 OR2X1_LOC_863/a_8_216# VDD 0.00fF
C54786 OR2X1_LOC_664/a_36_216# OR2X1_LOC_78/A 0.02fF
C54787 VDD OR2X1_LOC_468/Y 0.25fF
C54788 VDD OR2X1_LOC_44/Y 1.19fF
C54789 AND2X1_LOC_64/Y AND2X1_LOC_698/a_36_24# 0.00fF
C54790 OR2X1_LOC_70/Y AND2X1_LOC_810/B 0.01fF
C54791 OR2X1_LOC_91/A OR2X1_LOC_65/B 0.03fF
C54792 VDD AND2X1_LOC_288/a_8_24# 0.00fF
C54793 OR2X1_LOC_137/a_36_216# AND2X1_LOC_95/Y 0.00fF
C54794 AND2X1_LOC_40/Y OR2X1_LOC_61/Y 0.00fF
C54795 AND2X1_LOC_657/A AND2X1_LOC_570/a_8_24# 0.01fF
C54796 AND2X1_LOC_70/Y OR2X1_LOC_87/A 0.65fF
C54797 OR2X1_LOC_8/Y OR2X1_LOC_246/a_8_216# 0.01fF
C54798 AND2X1_LOC_385/a_8_24# VDD -0.00fF
C54799 AND2X1_LOC_91/B AND2X1_LOC_600/a_8_24# 0.09fF
C54800 AND2X1_LOC_572/Y AND2X1_LOC_367/A 0.09fF
C54801 OR2X1_LOC_9/Y OR2X1_LOC_74/A 0.53fF
C54802 AND2X1_LOC_390/B OR2X1_LOC_13/Y 0.16fF
C54803 OR2X1_LOC_186/Y AND2X1_LOC_51/Y 0.04fF
C54804 AND2X1_LOC_866/A AND2X1_LOC_792/a_8_24# -0.01fF
C54805 OR2X1_LOC_495/Y AND2X1_LOC_840/A 0.03fF
C54806 OR2X1_LOC_495/a_8_216# OR2X1_LOC_56/A 0.02fF
C54807 OR2X1_LOC_137/Y OR2X1_LOC_66/A 0.00fF
C54808 AND2X1_LOC_512/Y OR2X1_LOC_39/A 0.10fF
C54809 AND2X1_LOC_863/a_8_24# OR2X1_LOC_619/Y 0.02fF
C54810 OR2X1_LOC_220/B OR2X1_LOC_220/A 0.00fF
C54811 OR2X1_LOC_417/Y OR2X1_LOC_603/Y 0.01fF
C54812 OR2X1_LOC_326/B OR2X1_LOC_620/Y 0.00fF
C54813 OR2X1_LOC_405/A OR2X1_LOC_473/a_8_216# 0.01fF
C54814 OR2X1_LOC_49/A OR2X1_LOC_293/a_8_216# 0.01fF
C54815 OR2X1_LOC_720/B OR2X1_LOC_720/Y 0.00fF
C54816 OR2X1_LOC_235/B OR2X1_LOC_235/a_8_216# 0.02fF
C54817 AND2X1_LOC_706/Y OR2X1_LOC_417/Y 0.39fF
C54818 OR2X1_LOC_703/B OR2X1_LOC_703/A 0.16fF
C54819 OR2X1_LOC_600/A OR2X1_LOC_817/a_8_216# 0.01fF
C54820 OR2X1_LOC_92/Y AND2X1_LOC_573/A 0.10fF
C54821 AND2X1_LOC_7/Y AND2X1_LOC_7/B 0.03fF
C54822 OR2X1_LOC_6/B OR2X1_LOC_778/A 0.00fF
C54823 VDD AND2X1_LOC_116/Y 0.21fF
C54824 OR2X1_LOC_46/A OR2X1_LOC_12/Y 0.25fF
C54825 OR2X1_LOC_485/A AND2X1_LOC_285/Y 0.02fF
C54826 OR2X1_LOC_703/A OR2X1_LOC_87/A 0.03fF
C54827 OR2X1_LOC_585/A OR2X1_LOC_59/Y 3.43fF
C54828 VDD OR2X1_LOC_675/a_8_216# 0.00fF
C54829 OR2X1_LOC_235/B OR2X1_LOC_403/B 0.01fF
C54830 OR2X1_LOC_91/Y AND2X1_LOC_168/a_8_24# 0.04fF
C54831 AND2X1_LOC_861/B AND2X1_LOC_862/a_8_24# 0.01fF
C54832 VDD OR2X1_LOC_846/B 0.27fF
C54833 AND2X1_LOC_208/B OR2X1_LOC_44/Y 0.01fF
C54834 OR2X1_LOC_756/B OR2X1_LOC_778/Y 0.03fF
C54835 AND2X1_LOC_12/Y AND2X1_LOC_305/a_8_24# 0.01fF
C54836 OR2X1_LOC_318/B AND2X1_LOC_36/Y 0.16fF
C54837 OR2X1_LOC_756/B OR2X1_LOC_472/A 0.07fF
C54838 OR2X1_LOC_3/Y AND2X1_LOC_94/Y 0.01fF
C54839 OR2X1_LOC_354/A OR2X1_LOC_449/B 0.46fF
C54840 OR2X1_LOC_154/A OR2X1_LOC_523/Y 0.05fF
C54841 AND2X1_LOC_796/a_8_24# AND2X1_LOC_727/A 0.01fF
C54842 AND2X1_LOC_578/A AND2X1_LOC_548/Y 0.02fF
C54843 OR2X1_LOC_65/B AND2X1_LOC_573/A 0.03fF
C54844 INPUT_4 OR2X1_LOC_30/a_8_216# 0.01fF
C54845 OR2X1_LOC_771/B OR2X1_LOC_68/B 1.25fF
C54846 AND2X1_LOC_227/Y OR2X1_LOC_12/Y 0.03fF
C54847 AND2X1_LOC_364/Y OR2X1_LOC_320/Y 0.27fF
C54848 AND2X1_LOC_553/a_8_24# OR2X1_LOC_22/Y 0.04fF
C54849 OR2X1_LOC_658/a_8_216# AND2X1_LOC_42/B 0.01fF
C54850 OR2X1_LOC_516/A OR2X1_LOC_39/A 0.01fF
C54851 OR2X1_LOC_95/Y OR2X1_LOC_323/Y 0.10fF
C54852 AND2X1_LOC_319/A OR2X1_LOC_432/Y 0.19fF
C54853 OR2X1_LOC_154/A OR2X1_LOC_732/a_36_216# 0.00fF
C54854 OR2X1_LOC_325/Y OR2X1_LOC_121/B 0.01fF
C54855 OR2X1_LOC_165/a_8_216# OR2X1_LOC_26/Y 0.07fF
C54856 AND2X1_LOC_48/A OR2X1_LOC_66/A 0.13fF
C54857 OR2X1_LOC_680/Y OR2X1_LOC_441/Y 0.03fF
C54858 OR2X1_LOC_212/B OR2X1_LOC_578/B 0.03fF
C54859 AND2X1_LOC_363/A OR2X1_LOC_427/A 0.04fF
C54860 OR2X1_LOC_193/a_8_216# AND2X1_LOC_41/Y 0.01fF
C54861 AND2X1_LOC_831/Y AND2X1_LOC_476/Y 0.09fF
C54862 OR2X1_LOC_649/B OR2X1_LOC_655/a_8_216# 0.02fF
C54863 OR2X1_LOC_846/a_8_216# OR2X1_LOC_848/A 0.03fF
C54864 OR2X1_LOC_600/A AND2X1_LOC_664/a_36_24# 0.00fF
C54865 OR2X1_LOC_87/a_8_216# OR2X1_LOC_87/Y 0.01fF
C54866 OR2X1_LOC_26/Y OR2X1_LOC_394/Y 0.01fF
C54867 VDD OR2X1_LOC_471/Y 0.50fF
C54868 OR2X1_LOC_358/a_8_216# OR2X1_LOC_130/A 0.23fF
C54869 OR2X1_LOC_68/B OR2X1_LOC_776/A 0.74fF
C54870 OR2X1_LOC_315/Y OR2X1_LOC_44/Y 0.11fF
C54871 OR2X1_LOC_81/a_8_216# OR2X1_LOC_69/A 0.01fF
C54872 OR2X1_LOC_154/A OR2X1_LOC_579/B 0.08fF
C54873 VDD OR2X1_LOC_655/B 0.26fF
C54874 OR2X1_LOC_18/Y AND2X1_LOC_288/a_36_24# 0.00fF
C54875 OR2X1_LOC_602/Y OR2X1_LOC_602/B 0.81fF
C54876 AND2X1_LOC_702/Y AND2X1_LOC_655/A 0.03fF
C54877 OR2X1_LOC_369/a_8_216# OR2X1_LOC_417/A 0.09fF
C54878 AND2X1_LOC_565/Y OR2X1_LOC_189/A 0.09fF
C54879 OR2X1_LOC_864/A AND2X1_LOC_59/Y 1.46fF
C54880 AND2X1_LOC_866/A AND2X1_LOC_243/Y 0.07fF
C54881 OR2X1_LOC_848/A OR2X1_LOC_848/a_36_216# 0.00fF
C54882 AND2X1_LOC_65/a_36_24# OR2X1_LOC_215/A -0.00fF
C54883 AND2X1_LOC_477/A AND2X1_LOC_469/B 0.00fF
C54884 AND2X1_LOC_361/a_8_24# OR2X1_LOC_47/Y 0.03fF
C54885 OR2X1_LOC_158/A AND2X1_LOC_798/A 0.03fF
C54886 OR2X1_LOC_475/Y OR2X1_LOC_61/Y 0.02fF
C54887 OR2X1_LOC_520/Y AND2X1_LOC_8/Y 0.01fF
C54888 AND2X1_LOC_554/Y OR2X1_LOC_89/A 0.15fF
C54889 OR2X1_LOC_643/A OR2X1_LOC_657/a_8_216# 0.05fF
C54890 OR2X1_LOC_74/A AND2X1_LOC_808/a_36_24# 0.01fF
C54891 AND2X1_LOC_568/B AND2X1_LOC_866/A 0.02fF
C54892 OR2X1_LOC_354/A OR2X1_LOC_121/B 0.01fF
C54893 OR2X1_LOC_26/Y AND2X1_LOC_286/Y 0.01fF
C54894 OR2X1_LOC_116/a_8_216# OR2X1_LOC_87/A 0.02fF
C54895 OR2X1_LOC_418/a_8_216# AND2X1_LOC_452/Y 0.03fF
C54896 VDD OR2X1_LOC_222/a_8_216# 0.21fF
C54897 AND2X1_LOC_59/Y OR2X1_LOC_633/B 0.02fF
C54898 OR2X1_LOC_837/Y OR2X1_LOC_46/A 0.01fF
C54899 OR2X1_LOC_6/a_8_216# OR2X1_LOC_6/A 0.01fF
C54900 AND2X1_LOC_106/a_8_24# OR2X1_LOC_66/A 0.02fF
C54901 OR2X1_LOC_604/A GATE_662 0.03fF
C54902 AND2X1_LOC_576/a_8_24# AND2X1_LOC_489/Y 0.02fF
C54903 AND2X1_LOC_572/Y OR2X1_LOC_490/Y 0.23fF
C54904 INPUT_0 AND2X1_LOC_199/a_8_24# 0.01fF
C54905 OR2X1_LOC_499/B OR2X1_LOC_62/B 0.02fF
C54906 AND2X1_LOC_758/a_8_24# GATE_662 0.13fF
C54907 OR2X1_LOC_859/a_8_216# OR2X1_LOC_859/A 0.05fF
C54908 OR2X1_LOC_774/Y OR2X1_LOC_865/a_8_216# 0.01fF
C54909 AND2X1_LOC_17/Y OR2X1_LOC_87/A 0.04fF
C54910 OR2X1_LOC_404/Y OR2X1_LOC_668/a_8_216# 0.00fF
C54911 AND2X1_LOC_712/B OR2X1_LOC_422/a_36_216# 0.00fF
C54912 AND2X1_LOC_787/A AND2X1_LOC_222/Y 1.94fF
C54913 OR2X1_LOC_6/B OR2X1_LOC_84/a_8_216# 0.01fF
C54914 OR2X1_LOC_416/Y AND2X1_LOC_642/Y 0.16fF
C54915 AND2X1_LOC_431/a_36_24# OR2X1_LOC_78/B 0.01fF
C54916 OR2X1_LOC_532/B OR2X1_LOC_778/a_36_216# 0.00fF
C54917 OR2X1_LOC_251/Y OR2X1_LOC_44/Y 0.15fF
C54918 OR2X1_LOC_736/Y OR2X1_LOC_741/A 0.06fF
C54919 OR2X1_LOC_122/Y AND2X1_LOC_845/Y 0.03fF
C54920 OR2X1_LOC_91/Y OR2X1_LOC_485/A 0.10fF
C54921 OR2X1_LOC_280/a_8_216# OR2X1_LOC_36/Y 0.01fF
C54922 AND2X1_LOC_731/Y OR2X1_LOC_47/Y 0.27fF
C54923 OR2X1_LOC_822/Y OR2X1_LOC_47/Y 0.01fF
C54924 OR2X1_LOC_814/A OR2X1_LOC_392/A 0.00fF
C54925 OR2X1_LOC_70/Y AND2X1_LOC_228/Y 0.03fF
C54926 AND2X1_LOC_64/Y OR2X1_LOC_446/B 0.70fF
C54927 INPUT_0 OR2X1_LOC_689/Y 0.02fF
C54928 AND2X1_LOC_476/Y AND2X1_LOC_405/a_8_24# 0.02fF
C54929 OR2X1_LOC_45/B AND2X1_LOC_657/A 0.10fF
C54930 AND2X1_LOC_47/a_8_24# AND2X1_LOC_51/Y 0.01fF
C54931 AND2X1_LOC_84/a_8_24# OR2X1_LOC_52/B 0.01fF
C54932 AND2X1_LOC_658/B AND2X1_LOC_620/Y 0.01fF
C54933 AND2X1_LOC_367/B OR2X1_LOC_47/Y 0.01fF
C54934 OR2X1_LOC_427/A AND2X1_LOC_687/B 0.09fF
C54935 VDD OR2X1_LOC_205/Y 0.12fF
C54936 OR2X1_LOC_232/a_36_216# OR2X1_LOC_585/A 0.00fF
C54937 AND2X1_LOC_91/B OR2X1_LOC_579/a_8_216# 0.02fF
C54938 OR2X1_LOC_280/Y OR2X1_LOC_26/Y 5.67fF
C54939 OR2X1_LOC_646/a_8_216# AND2X1_LOC_8/Y 0.06fF
C54940 OR2X1_LOC_114/B AND2X1_LOC_72/B 0.01fF
C54941 OR2X1_LOC_32/Y AND2X1_LOC_34/a_8_24# 0.11fF
C54942 AND2X1_LOC_345/Y AND2X1_LOC_818/a_8_24# 0.02fF
C54943 OR2X1_LOC_189/Y AND2X1_LOC_474/Y 1.42fF
C54944 OR2X1_LOC_46/A OR2X1_LOC_393/Y 0.01fF
C54945 OR2X1_LOC_87/A OR2X1_LOC_206/a_8_216# 0.02fF
C54946 AND2X1_LOC_81/B AND2X1_LOC_51/Y 2.53fF
C54947 OR2X1_LOC_196/B OR2X1_LOC_161/A 0.07fF
C54948 OR2X1_LOC_778/B D_INPUT_1 0.16fF
C54949 OR2X1_LOC_743/A OR2X1_LOC_423/a_36_216# 0.00fF
C54950 OR2X1_LOC_54/Y OR2X1_LOC_39/A 0.01fF
C54951 OR2X1_LOC_404/Y OR2X1_LOC_87/A 0.00fF
C54952 OR2X1_LOC_280/Y OR2X1_LOC_89/A 0.03fF
C54953 AND2X1_LOC_119/a_36_24# OR2X1_LOC_375/A 0.00fF
C54954 AND2X1_LOC_7/B OR2X1_LOC_515/a_8_216# 0.01fF
C54955 OR2X1_LOC_70/Y OR2X1_LOC_585/A 0.09fF
C54956 OR2X1_LOC_462/B OR2X1_LOC_416/Y 0.39fF
C54957 AND2X1_LOC_621/a_36_24# AND2X1_LOC_621/Y 0.00fF
C54958 OR2X1_LOC_477/B AND2X1_LOC_51/Y 0.03fF
C54959 OR2X1_LOC_175/Y OR2X1_LOC_788/B 0.14fF
C54960 AND2X1_LOC_56/B OR2X1_LOC_34/B 0.01fF
C54961 AND2X1_LOC_358/Y OR2X1_LOC_437/A 0.00fF
C54962 OR2X1_LOC_344/A OR2X1_LOC_367/B 0.42fF
C54963 OR2X1_LOC_66/A OR2X1_LOC_398/a_8_216# 0.03fF
C54964 OR2X1_LOC_52/Y OR2X1_LOC_690/A 0.02fF
C54965 OR2X1_LOC_6/B OR2X1_LOC_560/A 0.02fF
C54966 OR2X1_LOC_527/Y AND2X1_LOC_474/Y 0.01fF
C54967 OR2X1_LOC_167/Y AND2X1_LOC_436/B 0.41fF
C54968 OR2X1_LOC_154/A OR2X1_LOC_68/Y 0.00fF
C54969 AND2X1_LOC_12/Y OR2X1_LOC_288/A 0.01fF
C54970 VDD OR2X1_LOC_750/Y 0.74fF
C54971 OR2X1_LOC_175/Y OR2X1_LOC_175/a_8_216# 0.01fF
C54972 OR2X1_LOC_444/a_36_216# OR2X1_LOC_87/A 0.02fF
C54973 OR2X1_LOC_47/Y AND2X1_LOC_852/B 0.25fF
C54974 AND2X1_LOC_44/Y OR2X1_LOC_712/B 0.06fF
C54975 OR2X1_LOC_22/Y OR2X1_LOC_26/Y 2.56fF
C54976 OR2X1_LOC_813/A AND2X1_LOC_266/Y 0.02fF
C54977 OR2X1_LOC_417/Y OR2X1_LOC_485/A 0.03fF
C54978 AND2X1_LOC_729/Y OR2X1_LOC_95/Y 0.58fF
C54979 OR2X1_LOC_47/Y OR2X1_LOC_48/B 0.18fF
C54980 OR2X1_LOC_154/A AND2X1_LOC_47/Y 0.48fF
C54981 OR2X1_LOC_36/Y OR2X1_LOC_607/a_8_216# 0.02fF
C54982 AND2X1_LOC_474/Y AND2X1_LOC_574/A 0.39fF
C54983 OR2X1_LOC_311/Y OR2X1_LOC_485/A 0.04fF
C54984 OR2X1_LOC_18/Y OR2X1_LOC_47/Y 0.23fF
C54985 OR2X1_LOC_22/Y OR2X1_LOC_89/A 0.18fF
C54986 OR2X1_LOC_816/Y AND2X1_LOC_793/B 0.00fF
C54987 OR2X1_LOC_485/A AND2X1_LOC_538/Y 0.01fF
C54988 OR2X1_LOC_744/A AND2X1_LOC_796/A 2.41fF
C54989 OR2X1_LOC_51/Y OR2X1_LOC_533/a_8_216# -0.00fF
C54990 OR2X1_LOC_485/A OR2X1_LOC_601/a_8_216# 0.02fF
C54991 OR2X1_LOC_139/a_8_216# OR2X1_LOC_244/A -0.05fF
C54992 AND2X1_LOC_784/A OR2X1_LOC_95/Y 0.07fF
C54993 OR2X1_LOC_532/B OR2X1_LOC_722/a_36_216# 0.00fF
C54994 AND2X1_LOC_845/a_8_24# OR2X1_LOC_278/Y 0.01fF
C54995 OR2X1_LOC_36/Y AND2X1_LOC_476/A 0.19fF
C54996 AND2X1_LOC_866/A AND2X1_LOC_620/a_8_24# 0.02fF
C54997 OR2X1_LOC_689/Y OR2X1_LOC_690/A 0.01fF
C54998 OR2X1_LOC_62/A OR2X1_LOC_824/Y 0.01fF
C54999 OR2X1_LOC_464/a_8_216# OR2X1_LOC_367/B 0.35fF
C55000 OR2X1_LOC_106/Y AND2X1_LOC_554/a_8_24# 0.03fF
C55001 AND2X1_LOC_12/Y AND2X1_LOC_72/B 0.03fF
C55002 OR2X1_LOC_702/A OR2X1_LOC_532/B 0.03fF
C55003 AND2X1_LOC_303/A OR2X1_LOC_289/a_36_216# 0.02fF
C55004 AND2X1_LOC_685/a_8_24# AND2X1_LOC_687/A 0.01fF
C55005 AND2X1_LOC_555/Y OR2X1_LOC_428/A 1.35fF
C55006 AND2X1_LOC_31/Y OR2X1_LOC_623/B 0.54fF
C55007 AND2X1_LOC_12/Y OR2X1_LOC_451/B 0.03fF
C55008 AND2X1_LOC_425/Y AND2X1_LOC_430/a_8_24# 0.01fF
C55009 AND2X1_LOC_22/Y OR2X1_LOC_175/Y 0.07fF
C55010 OR2X1_LOC_272/Y AND2X1_LOC_227/Y 0.02fF
C55011 OR2X1_LOC_485/A D_INPUT_3 0.10fF
C55012 AND2X1_LOC_672/B OR2X1_LOC_54/Y 0.03fF
C55013 AND2X1_LOC_271/a_8_24# OR2X1_LOC_269/B 0.01fF
C55014 OR2X1_LOC_523/Y OR2X1_LOC_560/A 0.44fF
C55015 AND2X1_LOC_580/A OR2X1_LOC_419/Y 0.03fF
C55016 OR2X1_LOC_154/A OR2X1_LOC_598/A 0.29fF
C55017 AND2X1_LOC_59/Y OR2X1_LOC_608/Y 0.06fF
C55018 AND2X1_LOC_396/a_8_24# AND2X1_LOC_36/Y 0.06fF
C55019 OR2X1_LOC_45/Y OR2X1_LOC_172/Y 0.20fF
C55020 OR2X1_LOC_351/B OR2X1_LOC_333/a_8_216# 0.01fF
C55021 OR2X1_LOC_338/a_8_216# OR2X1_LOC_338/B 0.06fF
C55022 OR2X1_LOC_139/A AND2X1_LOC_44/Y 0.07fF
C55023 AND2X1_LOC_22/Y OR2X1_LOC_691/Y 0.06fF
C55024 OR2X1_LOC_476/B OR2X1_LOC_532/B 0.50fF
C55025 OR2X1_LOC_175/Y AND2X1_LOC_417/a_36_24# 0.00fF
C55026 AND2X1_LOC_632/a_36_24# OR2X1_LOC_95/Y 0.01fF
C55027 OR2X1_LOC_759/A OR2X1_LOC_759/Y 0.00fF
C55028 OR2X1_LOC_116/a_36_216# OR2X1_LOC_66/Y 0.00fF
C55029 AND2X1_LOC_64/Y OR2X1_LOC_719/B 0.22fF
C55030 AND2X1_LOC_663/A OR2X1_LOC_142/Y 0.76fF
C55031 AND2X1_LOC_7/B OR2X1_LOC_390/A 0.03fF
C55032 OR2X1_LOC_850/B OR2X1_LOC_580/A 0.05fF
C55033 OR2X1_LOC_665/Y AND2X1_LOC_483/Y 0.03fF
C55034 OR2X1_LOC_691/Y OR2X1_LOC_855/a_36_216# 0.02fF
C55035 OR2X1_LOC_473/Y OR2X1_LOC_223/A 0.09fF
C55036 OR2X1_LOC_160/B OR2X1_LOC_333/a_36_216# 0.00fF
C55037 OR2X1_LOC_696/A AND2X1_LOC_738/B 0.19fF
C55038 OR2X1_LOC_696/A OR2X1_LOC_56/A 13.19fF
C55039 OR2X1_LOC_378/Y OR2X1_LOC_378/a_36_216# 0.00fF
C55040 AND2X1_LOC_70/Y OR2X1_LOC_390/B 0.18fF
C55041 OR2X1_LOC_417/Y AND2X1_LOC_645/a_36_24# 0.01fF
C55042 OR2X1_LOC_528/Y AND2X1_LOC_564/A 0.00fF
C55043 OR2X1_LOC_527/a_36_216# AND2X1_LOC_564/B 0.01fF
C55044 OR2X1_LOC_70/A OR2X1_LOC_585/A 0.10fF
C55045 AND2X1_LOC_771/B AND2X1_LOC_771/a_8_24# 0.11fF
C55046 OR2X1_LOC_85/A AND2X1_LOC_203/a_36_24# 0.00fF
C55047 OR2X1_LOC_744/A OR2X1_LOC_743/Y 0.01fF
C55048 OR2X1_LOC_755/A AND2X1_LOC_792/Y 0.03fF
C55049 D_INPUT_5 AND2X1_LOC_36/Y 0.06fF
C55050 AND2X1_LOC_621/Y OR2X1_LOC_437/A 0.07fF
C55051 OR2X1_LOC_162/Y AND2X1_LOC_163/a_8_24# 0.23fF
C55052 AND2X1_LOC_773/Y OR2X1_LOC_40/Y 0.03fF
C55053 AND2X1_LOC_51/Y OR2X1_LOC_66/Y 0.05fF
C55054 OR2X1_LOC_778/A OR2X1_LOC_598/A 0.01fF
C55055 OR2X1_LOC_147/B OR2X1_LOC_469/B 6.63fF
C55056 OR2X1_LOC_308/A OR2X1_LOC_78/A 0.01fF
C55057 OR2X1_LOC_177/Y AND2X1_LOC_180/a_8_24# 0.11fF
C55058 AND2X1_LOC_383/a_8_24# OR2X1_LOC_56/A 0.01fF
C55059 OR2X1_LOC_406/Y AND2X1_LOC_657/Y 0.01fF
C55060 AND2X1_LOC_477/Y AND2X1_LOC_212/Y 0.93fF
C55061 AND2X1_LOC_715/Y OR2X1_LOC_56/A 0.02fF
C55062 OR2X1_LOC_156/B OR2X1_LOC_160/B 0.01fF
C55063 OR2X1_LOC_45/B VDD 1.30fF
C55064 AND2X1_LOC_564/B OR2X1_LOC_59/Y 0.07fF
C55065 OR2X1_LOC_502/A OR2X1_LOC_502/a_8_216# 0.01fF
C55066 OR2X1_LOC_19/B AND2X1_LOC_845/a_8_24# 0.17fF
C55067 OR2X1_LOC_597/A OR2X1_LOC_16/A 0.00fF
C55068 OR2X1_LOC_51/Y OR2X1_LOC_428/A 0.78fF
C55069 OR2X1_LOC_62/A OR2X1_LOC_95/Y 0.11fF
C55070 AND2X1_LOC_91/B OR2X1_LOC_756/B 0.65fF
C55071 OR2X1_LOC_364/A OR2X1_LOC_544/B 0.32fF
C55072 OR2X1_LOC_151/A OR2X1_LOC_631/A 0.02fF
C55073 OR2X1_LOC_263/a_36_216# OR2X1_LOC_67/Y 0.01fF
C55074 AND2X1_LOC_359/B OR2X1_LOC_13/B 0.14fF
C55075 AND2X1_LOC_12/Y AND2X1_LOC_36/Y 1.98fF
C55076 AND2X1_LOC_53/Y OR2X1_LOC_214/B 0.01fF
C55077 AND2X1_LOC_180/a_36_24# OR2X1_LOC_40/Y 0.00fF
C55078 OR2X1_LOC_51/Y OR2X1_LOC_595/A 0.00fF
C55079 VDD OR2X1_LOC_382/A -0.00fF
C55080 OR2X1_LOC_851/B VDD 0.12fF
C55081 OR2X1_LOC_125/a_8_216# OR2X1_LOC_158/A 0.14fF
C55082 OR2X1_LOC_40/Y AND2X1_LOC_243/Y 0.01fF
C55083 OR2X1_LOC_643/Y OR2X1_LOC_641/B 0.72fF
C55084 OR2X1_LOC_692/Y OR2X1_LOC_91/A 0.10fF
C55085 OR2X1_LOC_19/B OR2X1_LOC_228/Y 3.79fF
C55086 OR2X1_LOC_467/B OR2X1_LOC_803/A 0.06fF
C55087 OR2X1_LOC_241/a_8_216# OR2X1_LOC_776/A 0.01fF
C55088 OR2X1_LOC_93/Y AND2X1_LOC_98/a_8_24# 0.23fF
C55089 OR2X1_LOC_696/A AND2X1_LOC_9/a_8_24# 0.01fF
C55090 OR2X1_LOC_40/Y AND2X1_LOC_568/B 0.07fF
C55091 AND2X1_LOC_12/Y OR2X1_LOC_333/a_8_216# 0.01fF
C55092 OR2X1_LOC_841/B AND2X1_LOC_36/Y 0.04fF
C55093 AND2X1_LOC_47/Y OR2X1_LOC_99/A 0.03fF
C55094 VDD AND2X1_LOC_410/a_8_24# 0.00fF
C55095 AND2X1_LOC_722/A OR2X1_LOC_12/Y 0.02fF
C55096 AND2X1_LOC_12/Y OR2X1_LOC_334/A 0.00fF
C55097 OR2X1_LOC_151/A OR2X1_LOC_632/Y 0.19fF
C55098 OR2X1_LOC_244/A OR2X1_LOC_398/a_36_216# 0.00fF
C55099 AND2X1_LOC_76/Y AND2X1_LOC_473/Y 0.03fF
C55100 OR2X1_LOC_276/B OR2X1_LOC_493/Y 0.10fF
C55101 AND2X1_LOC_212/A AND2X1_LOC_365/a_8_24# 0.01fF
C55102 AND2X1_LOC_217/Y OR2X1_LOC_132/a_36_216# 0.02fF
C55103 AND2X1_LOC_352/a_8_24# OR2X1_LOC_329/B 0.05fF
C55104 OR2X1_LOC_3/Y AND2X1_LOC_449/a_8_24# 0.01fF
C55105 OR2X1_LOC_756/B OR2X1_LOC_364/a_8_216# 0.01fF
C55106 OR2X1_LOC_178/Y OR2X1_LOC_108/Y 0.08fF
C55107 AND2X1_LOC_70/Y OR2X1_LOC_389/A 0.01fF
C55108 AND2X1_LOC_42/B OR2X1_LOC_217/A 0.02fF
C55109 AND2X1_LOC_566/B AND2X1_LOC_367/A 0.02fF
C55110 AND2X1_LOC_353/a_8_24# AND2X1_LOC_364/Y 0.01fF
C55111 OR2X1_LOC_324/A AND2X1_LOC_44/Y 0.04fF
C55112 OR2X1_LOC_715/B OR2X1_LOC_678/Y 0.01fF
C55113 VDD OR2X1_LOC_809/B 0.07fF
C55114 AND2X1_LOC_373/a_8_24# OR2X1_LOC_180/B 0.01fF
C55115 AND2X1_LOC_675/A AND2X1_LOC_222/Y 0.03fF
C55116 OR2X1_LOC_651/A AND2X1_LOC_52/Y 0.09fF
C55117 AND2X1_LOC_391/Y OR2X1_LOC_600/A 1.32fF
C55118 OR2X1_LOC_87/A OR2X1_LOC_718/a_8_216# 0.01fF
C55119 AND2X1_LOC_79/Y AND2X1_LOC_36/Y 0.01fF
C55120 AND2X1_LOC_59/Y OR2X1_LOC_121/A 0.01fF
C55121 OR2X1_LOC_435/Y OR2X1_LOC_174/Y 0.03fF
C55122 OR2X1_LOC_600/A OR2X1_LOC_91/A 3.98fF
C55123 AND2X1_LOC_64/Y AND2X1_LOC_56/B 11.23fF
C55124 OR2X1_LOC_479/Y OR2X1_LOC_593/B 0.19fF
C55125 AND2X1_LOC_335/Y OR2X1_LOC_91/A 0.03fF
C55126 AND2X1_LOC_47/Y OR2X1_LOC_560/A 0.00fF
C55127 OR2X1_LOC_135/Y AND2X1_LOC_649/B 0.19fF
C55128 AND2X1_LOC_658/A AND2X1_LOC_865/A 0.16fF
C55129 AND2X1_LOC_496/a_8_24# AND2X1_LOC_36/Y 0.01fF
C55130 AND2X1_LOC_3/Y OR2X1_LOC_508/Y 0.03fF
C55131 OR2X1_LOC_160/B OR2X1_LOC_803/a_8_216# 0.01fF
C55132 OR2X1_LOC_45/B OR2X1_LOC_315/Y 0.06fF
C55133 VDD OR2X1_LOC_292/a_8_216# 0.00fF
C55134 OR2X1_LOC_427/A OR2X1_LOC_322/a_8_216# 0.01fF
C55135 OR2X1_LOC_122/a_8_216# OR2X1_LOC_56/A 0.02fF
C55136 AND2X1_LOC_6/a_8_24# OR2X1_LOC_598/A 0.02fF
C55137 OR2X1_LOC_421/A OR2X1_LOC_763/a_8_216# 0.05fF
C55138 OR2X1_LOC_56/Y OR2X1_LOC_6/A 0.00fF
C55139 AND2X1_LOC_64/Y AND2X1_LOC_8/Y 0.09fF
C55140 OR2X1_LOC_231/A AND2X1_LOC_65/A 0.08fF
C55141 OR2X1_LOC_377/A OR2X1_LOC_548/B 0.13fF
C55142 OR2X1_LOC_125/a_8_216# AND2X1_LOC_98/Y 0.47fF
C55143 OR2X1_LOC_118/a_36_216# AND2X1_LOC_573/A 0.01fF
C55144 AND2X1_LOC_201/a_36_24# OR2X1_LOC_72/Y 0.01fF
C55145 AND2X1_LOC_43/B OR2X1_LOC_161/B 8.08fF
C55146 OR2X1_LOC_756/B OR2X1_LOC_645/a_8_216# 0.01fF
C55147 AND2X1_LOC_647/Y AND2X1_LOC_647/B 1.20fF
C55148 OR2X1_LOC_313/a_8_216# OR2X1_LOC_16/A 0.05fF
C55149 OR2X1_LOC_185/Y OR2X1_LOC_474/B 0.01fF
C55150 AND2X1_LOC_454/Y OR2X1_LOC_12/Y 0.15fF
C55151 AND2X1_LOC_562/a_36_24# OR2X1_LOC_36/Y 0.00fF
C55152 OR2X1_LOC_404/Y OR2X1_LOC_844/B 0.19fF
C55153 OR2X1_LOC_542/B OR2X1_LOC_464/A 0.06fF
C55154 AND2X1_LOC_64/Y AND2X1_LOC_21/Y 0.01fF
C55155 OR2X1_LOC_6/A AND2X1_LOC_231/a_36_24# 0.00fF
C55156 AND2X1_LOC_70/Y AND2X1_LOC_177/a_8_24# 0.07fF
C55157 OR2X1_LOC_565/A OR2X1_LOC_553/B 0.18fF
C55158 OR2X1_LOC_696/A OR2X1_LOC_291/A 0.00fF
C55159 OR2X1_LOC_653/a_8_216# OR2X1_LOC_390/B 0.05fF
C55160 OR2X1_LOC_326/B AND2X1_LOC_299/a_8_24# 0.01fF
C55161 OR2X1_LOC_185/A OR2X1_LOC_729/a_8_216# 0.05fF
C55162 VDD OR2X1_LOC_852/B -0.00fF
C55163 AND2X1_LOC_229/a_36_24# OR2X1_LOC_130/A 0.00fF
C55164 OR2X1_LOC_859/A OR2X1_LOC_576/a_8_216# 0.07fF
C55165 OR2X1_LOC_45/B AND2X1_LOC_267/a_8_24# 0.06fF
C55166 OR2X1_LOC_36/Y AND2X1_LOC_445/a_8_24# 0.04fF
C55167 OR2X1_LOC_842/a_8_216# OR2X1_LOC_287/A 0.40fF
C55168 OR2X1_LOC_805/A OR2X1_LOC_390/A 0.03fF
C55169 OR2X1_LOC_710/a_8_216# AND2X1_LOC_7/B 0.06fF
C55170 AND2X1_LOC_473/Y OR2X1_LOC_52/B 0.01fF
C55171 AND2X1_LOC_65/A OR2X1_LOC_340/Y 0.03fF
C55172 OR2X1_LOC_479/Y AND2X1_LOC_273/a_8_24# 0.03fF
C55173 OR2X1_LOC_49/A AND2X1_LOC_404/a_8_24# 0.03fF
C55174 AND2X1_LOC_347/Y OR2X1_LOC_59/Y 0.04fF
C55175 AND2X1_LOC_592/Y AND2X1_LOC_593/Y 0.01fF
C55176 OR2X1_LOC_117/a_8_216# OR2X1_LOC_117/Y 0.04fF
C55177 AND2X1_LOC_43/B OR2X1_LOC_514/a_36_216# 0.02fF
C55178 OR2X1_LOC_486/Y OR2X1_LOC_553/A 0.07fF
C55179 AND2X1_LOC_857/Y OR2X1_LOC_59/Y 0.03fF
C55180 AND2X1_LOC_732/B OR2X1_LOC_48/B 0.01fF
C55181 OR2X1_LOC_840/A OR2X1_LOC_834/A 0.00fF
C55182 OR2X1_LOC_776/a_36_216# AND2X1_LOC_92/Y 0.01fF
C55183 OR2X1_LOC_599/A OR2X1_LOC_12/Y 0.11fF
C55184 AND2X1_LOC_737/a_8_24# AND2X1_LOC_443/Y 0.20fF
C55185 AND2X1_LOC_346/a_8_24# AND2X1_LOC_848/Y 0.04fF
C55186 OR2X1_LOC_18/Y OR2X1_LOC_607/A 0.01fF
C55187 OR2X1_LOC_156/a_8_216# OR2X1_LOC_479/Y 0.03fF
C55188 AND2X1_LOC_95/Y OR2X1_LOC_461/B 0.51fF
C55189 AND2X1_LOC_31/a_36_24# INPUT_6 0.00fF
C55190 OR2X1_LOC_316/a_8_216# OR2X1_LOC_60/a_8_216# 0.47fF
C55191 AND2X1_LOC_94/Y OR2X1_LOC_502/A 0.03fF
C55192 AND2X1_LOC_464/A AND2X1_LOC_458/a_8_24# 0.01fF
C55193 AND2X1_LOC_164/a_8_24# OR2X1_LOC_502/A 0.01fF
C55194 OR2X1_LOC_26/Y AND2X1_LOC_445/a_36_24# 0.00fF
C55195 AND2X1_LOC_62/a_36_24# OR2X1_LOC_600/A 0.01fF
C55196 OR2X1_LOC_208/a_8_216# AND2X1_LOC_44/Y 0.01fF
C55197 OR2X1_LOC_304/a_8_216# OR2X1_LOC_3/Y 0.01fF
C55198 AND2X1_LOC_564/B AND2X1_LOC_711/Y 0.13fF
C55199 AND2X1_LOC_713/a_8_24# OR2X1_LOC_44/Y 0.02fF
C55200 OR2X1_LOC_141/B OR2X1_LOC_576/A 0.01fF
C55201 OR2X1_LOC_194/Y OR2X1_LOC_596/A 0.10fF
C55202 AND2X1_LOC_387/a_8_24# OR2X1_LOC_161/A 0.02fF
C55203 OR2X1_LOC_600/A AND2X1_LOC_573/A 0.10fF
C55204 AND2X1_LOC_99/A OR2X1_LOC_426/B 0.07fF
C55205 AND2X1_LOC_97/a_8_24# OR2X1_LOC_666/A 0.01fF
C55206 OR2X1_LOC_175/B OR2X1_LOC_78/B 0.00fF
C55207 AND2X1_LOC_564/B OR2X1_LOC_70/Y 0.07fF
C55208 AND2X1_LOC_787/A OR2X1_LOC_74/A 0.03fF
C55209 OR2X1_LOC_160/A VDD 1.90fF
C55210 AND2X1_LOC_503/a_36_24# OR2X1_LOC_78/B 0.01fF
C55211 OR2X1_LOC_778/B OR2X1_LOC_737/A 0.07fF
C55212 AND2X1_LOC_841/B AND2X1_LOC_434/Y 0.07fF
C55213 AND2X1_LOC_367/B OR2X1_LOC_625/Y 0.10fF
C55214 OR2X1_LOC_325/a_8_216# OR2X1_LOC_538/A 0.01fF
C55215 AND2X1_LOC_712/a_8_24# OR2X1_LOC_3/Y 0.00fF
C55216 OR2X1_LOC_482/Y AND2X1_LOC_859/Y 0.01fF
C55217 OR2X1_LOC_682/a_8_216# OR2X1_LOC_158/A 0.01fF
C55218 OR2X1_LOC_243/B AND2X1_LOC_235/a_8_24# 0.01fF
C55219 OR2X1_LOC_604/A AND2X1_LOC_580/A 0.07fF
C55220 VDD OR2X1_LOC_767/a_8_216# 0.21fF
C55221 AND2X1_LOC_504/a_8_24# OR2X1_LOC_78/A 0.09fF
C55222 OR2X1_LOC_128/B OR2X1_LOC_244/Y 0.39fF
C55223 AND2X1_LOC_773/Y OR2X1_LOC_320/Y 0.56fF
C55224 OR2X1_LOC_129/a_8_216# OR2X1_LOC_69/Y 0.05fF
C55225 OR2X1_LOC_709/A AND2X1_LOC_516/a_36_24# 0.00fF
C55226 OR2X1_LOC_653/A AND2X1_LOC_18/Y 0.01fF
C55227 AND2X1_LOC_50/Y OR2X1_LOC_502/A 0.06fF
C55228 OR2X1_LOC_631/B OR2X1_LOC_629/B 0.02fF
C55229 OR2X1_LOC_663/a_8_216# OR2X1_LOC_557/A 0.01fF
C55230 OR2X1_LOC_91/A OR2X1_LOC_619/Y 0.08fF
C55231 OR2X1_LOC_490/a_8_216# OR2X1_LOC_3/Y 0.01fF
C55232 OR2X1_LOC_673/Y AND2X1_LOC_18/Y 0.51fF
C55233 AND2X1_LOC_86/a_8_24# AND2X1_LOC_8/Y 0.04fF
C55234 AND2X1_LOC_456/B OR2X1_LOC_278/Y 0.02fF
C55235 OR2X1_LOC_485/Y OR2X1_LOC_26/Y 0.02fF
C55236 AND2X1_LOC_458/Y OR2X1_LOC_56/A 0.01fF
C55237 AND2X1_LOC_552/A OR2X1_LOC_280/Y 0.02fF
C55238 OR2X1_LOC_653/Y AND2X1_LOC_749/a_8_24# 0.03fF
C55239 AND2X1_LOC_302/a_8_24# OR2X1_LOC_56/A 0.09fF
C55240 INPUT_0 OR2X1_LOC_243/A 0.03fF
C55241 OR2X1_LOC_687/Y OR2X1_LOC_702/a_8_216# 0.04fF
C55242 OR2X1_LOC_121/Y AND2X1_LOC_122/a_8_24# 0.02fF
C55243 OR2X1_LOC_750/A AND2X1_LOC_7/B 0.01fF
C55244 OR2X1_LOC_114/B OR2X1_LOC_346/B 0.03fF
C55245 OR2X1_LOC_756/B OR2X1_LOC_799/A 0.04fF
C55246 OR2X1_LOC_804/a_8_216# OR2X1_LOC_161/A 0.12fF
C55247 OR2X1_LOC_520/Y AND2X1_LOC_92/Y 0.01fF
C55248 OR2X1_LOC_76/A AND2X1_LOC_604/a_8_24# 0.02fF
C55249 OR2X1_LOC_691/A AND2X1_LOC_689/a_8_24# 0.01fF
C55250 OR2X1_LOC_124/B OR2X1_LOC_124/Y 0.16fF
C55251 OR2X1_LOC_6/B AND2X1_LOC_495/a_36_24# 0.01fF
C55252 OR2X1_LOC_8/Y OR2X1_LOC_824/Y 0.00fF
C55253 INPUT_1 OR2X1_LOC_415/Y 0.05fF
C55254 AND2X1_LOC_512/Y AND2X1_LOC_593/Y 0.07fF
C55255 OR2X1_LOC_7/A AND2X1_LOC_243/Y 0.07fF
C55256 OR2X1_LOC_2/Y OR2X1_LOC_40/a_8_216# 0.07fF
C55257 OR2X1_LOC_665/Y AND2X1_LOC_254/a_36_24# 0.01fF
C55258 OR2X1_LOC_784/a_8_216# OR2X1_LOC_784/B 0.39fF
C55259 AND2X1_LOC_707/a_8_24# OR2X1_LOC_52/B 0.02fF
C55260 AND2X1_LOC_568/B OR2X1_LOC_7/A 0.19fF
C55261 INPUT_0 OR2X1_LOC_36/Y 6.37fF
C55262 OR2X1_LOC_43/A OR2X1_LOC_90/a_8_216# 0.07fF
C55263 OR2X1_LOC_195/A AND2X1_LOC_18/Y 0.98fF
C55264 VDD OR2X1_LOC_261/Y 0.10fF
C55265 OR2X1_LOC_312/Y AND2X1_LOC_436/Y 0.03fF
C55266 OR2X1_LOC_635/A AND2X1_LOC_12/Y 0.46fF
C55267 AND2X1_LOC_3/Y OR2X1_LOC_66/A 0.34fF
C55268 OR2X1_LOC_139/A OR2X1_LOC_720/B 0.60fF
C55269 OR2X1_LOC_756/B OR2X1_LOC_270/a_8_216# 0.04fF
C55270 VDD AND2X1_LOC_86/B 0.48fF
C55271 AND2X1_LOC_95/Y AND2X1_LOC_74/a_8_24# 0.06fF
C55272 OR2X1_LOC_185/Y OR2X1_LOC_274/a_8_216# 0.04fF
C55273 OR2X1_LOC_250/a_36_216# OR2X1_LOC_278/Y 0.00fF
C55274 OR2X1_LOC_382/Y OR2X1_LOC_6/A 0.01fF
C55275 OR2X1_LOC_620/Y OR2X1_LOC_506/A 0.07fF
C55276 AND2X1_LOC_330/a_8_24# OR2X1_LOC_485/A 0.17fF
C55277 AND2X1_LOC_125/a_36_24# OR2X1_LOC_161/A 0.00fF
C55278 INPUT_1 AND2X1_LOC_786/Y 0.16fF
C55279 VDD OR2X1_LOC_430/a_8_216# 0.00fF
C55280 AND2X1_LOC_720/a_8_24# OR2X1_LOC_18/Y 0.17fF
C55281 OR2X1_LOC_319/a_8_216# OR2X1_LOC_624/A 0.39fF
C55282 OR2X1_LOC_474/Y OR2X1_LOC_87/A 6.09fF
C55283 OR2X1_LOC_625/Y OR2X1_LOC_18/Y 0.03fF
C55284 AND2X1_LOC_56/B OR2X1_LOC_464/A 0.03fF
C55285 OR2X1_LOC_782/a_8_216# OR2X1_LOC_160/Y 0.08fF
C55286 OR2X1_LOC_74/Y OR2X1_LOC_265/Y 0.02fF
C55287 OR2X1_LOC_62/B AND2X1_LOC_65/A 0.01fF
C55288 OR2X1_LOC_682/Y OR2X1_LOC_421/a_8_216# 0.39fF
C55289 AND2X1_LOC_851/B AND2X1_LOC_242/B 0.01fF
C55290 OR2X1_LOC_485/a_36_216# OR2X1_LOC_511/Y 0.02fF
C55291 OR2X1_LOC_619/Y AND2X1_LOC_573/A 0.07fF
C55292 AND2X1_LOC_596/a_8_24# OR2X1_LOC_64/Y 0.01fF
C55293 OR2X1_LOC_158/A AND2X1_LOC_326/a_8_24# 0.08fF
C55294 OR2X1_LOC_391/B OR2X1_LOC_489/a_8_216# 0.05fF
C55295 OR2X1_LOC_724/A OR2X1_LOC_714/A 0.01fF
C55296 AND2X1_LOC_40/Y OR2X1_LOC_593/a_36_216# 0.00fF
C55297 AND2X1_LOC_316/a_36_24# OR2X1_LOC_87/A 0.01fF
C55298 OR2X1_LOC_141/B AND2X1_LOC_41/A 0.00fF
C55299 AND2X1_LOC_486/Y OR2X1_LOC_44/Y 0.01fF
C55300 OR2X1_LOC_544/B OR2X1_LOC_578/B 0.00fF
C55301 AND2X1_LOC_817/B OR2X1_LOC_847/A 0.00fF
C55302 OR2X1_LOC_814/A OR2X1_LOC_349/A 0.37fF
C55303 AND2X1_LOC_117/a_8_24# OR2X1_LOC_78/A 0.07fF
C55304 AND2X1_LOC_47/Y OR2X1_LOC_435/A 0.04fF
C55305 AND2X1_LOC_671/a_8_24# INPUT_2 0.10fF
C55306 AND2X1_LOC_474/A OR2X1_LOC_279/a_8_216# 0.01fF
C55307 AND2X1_LOC_70/Y OR2X1_LOC_639/A 0.01fF
C55308 AND2X1_LOC_663/B OR2X1_LOC_56/A 0.07fF
C55309 OR2X1_LOC_154/A OR2X1_LOC_506/A 0.03fF
C55310 AND2X1_LOC_866/A OR2X1_LOC_12/Y 0.08fF
C55311 OR2X1_LOC_494/a_8_216# OR2X1_LOC_485/A 0.01fF
C55312 AND2X1_LOC_159/a_8_24# OR2X1_LOC_575/A 0.01fF
C55313 AND2X1_LOC_95/Y OR2X1_LOC_720/A 0.01fF
C55314 OR2X1_LOC_519/a_8_216# AND2X1_LOC_354/B 0.01fF
C55315 AND2X1_LOC_332/a_36_24# OR2X1_LOC_111/Y 0.00fF
C55316 AND2X1_LOC_710/Y AND2X1_LOC_663/B 0.79fF
C55317 D_INPUT_7 AND2X1_LOC_2/a_8_24# 0.01fF
C55318 AND2X1_LOC_449/Y AND2X1_LOC_453/a_8_24# 0.03fF
C55319 OR2X1_LOC_479/a_8_216# AND2X1_LOC_92/Y 0.06fF
C55320 OR2X1_LOC_810/A OR2X1_LOC_575/A 0.06fF
C55321 OR2X1_LOC_88/A AND2X1_LOC_573/A 0.01fF
C55322 D_INPUT_0 AND2X1_LOC_625/a_8_24# 0.01fF
C55323 OR2X1_LOC_722/a_8_216# OR2X1_LOC_737/A 0.02fF
C55324 AND2X1_LOC_482/a_8_24# AND2X1_LOC_252/a_8_24# 0.23fF
C55325 OR2X1_LOC_114/B AND2X1_LOC_127/a_36_24# 0.00fF
C55326 OR2X1_LOC_624/A OR2X1_LOC_203/Y 0.10fF
C55327 OR2X1_LOC_837/B OR2X1_LOC_32/a_8_216# 0.05fF
C55328 OR2X1_LOC_462/a_8_216# INPUT_0 0.03fF
C55329 VDD OR2X1_LOC_655/A -0.00fF
C55330 OR2X1_LOC_76/Y AND2X1_LOC_72/Y 0.17fF
C55331 OR2X1_LOC_613/Y AND2X1_LOC_624/A 0.00fF
C55332 AND2X1_LOC_660/Y OR2X1_LOC_275/Y 0.00fF
C55333 OR2X1_LOC_629/Y OR2X1_LOC_296/a_8_216# 0.05fF
C55334 AND2X1_LOC_147/a_8_24# OR2X1_LOC_74/A 0.05fF
C55335 OR2X1_LOC_400/B OR2X1_LOC_377/A 0.05fF
C55336 OR2X1_LOC_810/A OR2X1_LOC_493/A 0.18fF
C55337 OR2X1_LOC_70/Y AND2X1_LOC_857/Y 0.03fF
C55338 AND2X1_LOC_152/a_8_24# OR2X1_LOC_739/A 0.01fF
C55339 AND2X1_LOC_342/Y OR2X1_LOC_85/A 0.35fF
C55340 OR2X1_LOC_47/Y AND2X1_LOC_810/B 0.07fF
C55341 OR2X1_LOC_458/B OR2X1_LOC_675/A 0.05fF
C55342 OR2X1_LOC_83/Y AND2X1_LOC_400/a_8_24# 0.01fF
C55343 OR2X1_LOC_45/B OR2X1_LOC_67/Y 0.03fF
C55344 OR2X1_LOC_36/Y OR2X1_LOC_11/Y 0.03fF
C55345 OR2X1_LOC_160/A OR2X1_LOC_836/B 0.01fF
C55346 OR2X1_LOC_26/Y OR2X1_LOC_39/A 2.19fF
C55347 OR2X1_LOC_291/Y AND2X1_LOC_647/a_8_24# 0.04fF
C55348 OR2X1_LOC_462/B OR2X1_LOC_6/A 0.80fF
C55349 AND2X1_LOC_807/Y OR2X1_LOC_52/B 0.80fF
C55350 OR2X1_LOC_652/a_8_216# OR2X1_LOC_810/A 0.03fF
C55351 INPUT_1 AND2X1_LOC_218/Y 0.03fF
C55352 OR2X1_LOC_333/B AND2X1_LOC_95/Y 0.05fF
C55353 OR2X1_LOC_574/A OR2X1_LOC_161/A 0.07fF
C55354 OR2X1_LOC_497/a_8_216# OR2X1_LOC_497/Y -0.02fF
C55355 OR2X1_LOC_54/Y AND2X1_LOC_240/a_8_24# 0.02fF
C55356 OR2X1_LOC_54/a_8_216# OR2X1_LOC_56/A 0.02fF
C55357 OR2X1_LOC_160/B OR2X1_LOC_783/A 0.00fF
C55358 OR2X1_LOC_687/Y OR2X1_LOC_269/B 0.03fF
C55359 AND2X1_LOC_514/Y AND2X1_LOC_857/Y 0.37fF
C55360 OR2X1_LOC_8/Y OR2X1_LOC_95/Y 0.40fF
C55361 VDD AND2X1_LOC_811/Y 0.24fF
C55362 OR2X1_LOC_185/A AND2X1_LOC_42/B 0.06fF
C55363 OR2X1_LOC_89/A OR2X1_LOC_39/A 1.14fF
C55364 OR2X1_LOC_219/B OR2X1_LOC_350/a_36_216# 0.02fF
C55365 AND2X1_LOC_520/a_8_24# AND2X1_LOC_222/Y 0.05fF
C55366 OR2X1_LOC_489/a_8_216# OR2X1_LOC_772/Y 0.04fF
C55367 OR2X1_LOC_744/A OR2X1_LOC_80/a_8_216# 0.01fF
C55368 OR2X1_LOC_36/Y OR2X1_LOC_690/A 0.02fF
C55369 AND2X1_LOC_42/B OR2X1_LOC_249/Y 0.01fF
C55370 OR2X1_LOC_709/A OR2X1_LOC_801/B 0.00fF
C55371 OR2X1_LOC_74/A OR2X1_LOC_406/a_8_216# 0.02fF
C55372 AND2X1_LOC_571/a_8_24# AND2X1_LOC_563/Y 0.01fF
C55373 OR2X1_LOC_756/B AND2X1_LOC_600/a_36_24# 0.01fF
C55374 OR2X1_LOC_864/a_8_216# OR2X1_LOC_772/a_8_216# 0.47fF
C55375 AND2X1_LOC_11/a_8_24# D_INPUT_4 0.04fF
C55376 OR2X1_LOC_7/Y OR2X1_LOC_16/a_8_216# 0.40fF
C55377 AND2X1_LOC_342/a_8_24# OR2X1_LOC_7/A 0.04fF
C55378 OR2X1_LOC_250/Y OR2X1_LOC_64/Y 0.16fF
C55379 OR2X1_LOC_461/Y OR2X1_LOC_39/A 0.09fF
C55380 AND2X1_LOC_211/B OR2X1_LOC_26/Y 0.11fF
C55381 VDD AND2X1_LOC_838/B 0.23fF
C55382 OR2X1_LOC_218/a_8_216# AND2X1_LOC_3/Y 0.01fF
C55383 OR2X1_LOC_151/A AND2X1_LOC_485/a_36_24# 0.01fF
C55384 OR2X1_LOC_485/A AND2X1_LOC_806/A 0.03fF
C55385 OR2X1_LOC_598/a_8_216# OR2X1_LOC_771/B 0.41fF
C55386 AND2X1_LOC_347/a_8_24# OR2X1_LOC_44/Y 0.01fF
C55387 AND2X1_LOC_213/B AND2X1_LOC_796/A 0.01fF
C55388 OR2X1_LOC_273/a_36_216# OR2X1_LOC_36/Y 0.03fF
C55389 OR2X1_LOC_76/Y OR2X1_LOC_455/A 0.12fF
C55390 OR2X1_LOC_456/Y OR2X1_LOC_456/A 0.00fF
C55391 OR2X1_LOC_733/A OR2X1_LOC_374/Y 0.01fF
C55392 AND2X1_LOC_364/A D_INPUT_0 0.26fF
C55393 OR2X1_LOC_377/A OR2X1_LOC_54/Y 0.29fF
C55394 AND2X1_LOC_845/a_36_24# AND2X1_LOC_845/Y 0.00fF
C55395 AND2X1_LOC_342/a_36_24# OR2X1_LOC_485/A 0.00fF
C55396 OR2X1_LOC_808/B OR2X1_LOC_440/A 2.30fF
C55397 OR2X1_LOC_306/a_8_216# OR2X1_LOC_22/Y 0.01fF
C55398 AND2X1_LOC_70/Y OR2X1_LOC_493/Y 0.01fF
C55399 AND2X1_LOC_81/B OR2X1_LOC_647/a_8_216# 0.49fF
C55400 OR2X1_LOC_64/Y OR2X1_LOC_36/Y 4.52fF
C55401 OR2X1_LOC_158/A AND2X1_LOC_657/A 0.08fF
C55402 OR2X1_LOC_623/a_8_216# OR2X1_LOC_532/B 0.01fF
C55403 OR2X1_LOC_161/B OR2X1_LOC_367/B 0.14fF
C55404 OR2X1_LOC_305/a_36_216# AND2X1_LOC_307/Y 0.00fF
C55405 OR2X1_LOC_85/A OR2X1_LOC_54/Y 0.54fF
C55406 AND2X1_LOC_17/Y OR2X1_LOC_639/A 0.01fF
C55407 OR2X1_LOC_816/Y AND2X1_LOC_846/a_8_24# 0.00fF
C55408 AND2X1_LOC_851/B AND2X1_LOC_841/B 0.01fF
C55409 OR2X1_LOC_574/A AND2X1_LOC_51/Y 0.76fF
C55410 OR2X1_LOC_613/Y AND2X1_LOC_621/a_8_24# 0.01fF
C55411 AND2X1_LOC_51/Y OR2X1_LOC_33/A 0.01fF
C55412 AND2X1_LOC_727/A OR2X1_LOC_52/B 0.03fF
C55413 INPUT_5 OR2X1_LOC_31/a_36_216# 0.00fF
C55414 OR2X1_LOC_64/Y AND2X1_LOC_493/a_36_24# 0.01fF
C55415 OR2X1_LOC_22/Y AND2X1_LOC_853/Y 0.02fF
C55416 OR2X1_LOC_599/A AND2X1_LOC_801/B 0.00fF
C55417 OR2X1_LOC_81/Y AND2X1_LOC_68/a_8_24# 0.23fF
C55418 OR2X1_LOC_36/Y OR2X1_LOC_417/A 0.15fF
C55419 OR2X1_LOC_91/a_8_216# OR2X1_LOC_417/A 0.03fF
C55420 AND2X1_LOC_42/B AND2X1_LOC_119/a_8_24# 0.00fF
C55421 OR2X1_LOC_62/B OR2X1_LOC_609/A 0.01fF
C55422 OR2X1_LOC_705/Y OR2X1_LOC_713/a_8_216# 0.03fF
C55423 OR2X1_LOC_357/a_8_216# OR2X1_LOC_212/B 0.41fF
C55424 OR2X1_LOC_45/B AND2X1_LOC_269/a_8_24# 0.01fF
C55425 OR2X1_LOC_625/Y AND2X1_LOC_620/Y 0.00fF
C55426 AND2X1_LOC_863/Y AND2X1_LOC_661/A 0.02fF
C55427 OR2X1_LOC_416/a_36_216# OR2X1_LOC_39/A 0.00fF
C55428 OR2X1_LOC_469/Y OR2X1_LOC_705/B 0.07fF
C55429 OR2X1_LOC_636/a_36_216# AND2X1_LOC_51/Y 0.00fF
C55430 AND2X1_LOC_91/B OR2X1_LOC_140/B 0.10fF
C55431 OR2X1_LOC_233/a_8_216# OR2X1_LOC_62/a_8_216# 0.47fF
C55432 OR2X1_LOC_829/Y AND2X1_LOC_855/a_8_24# 0.23fF
C55433 AND2X1_LOC_729/B AND2X1_LOC_856/B 0.01fF
C55434 OR2X1_LOC_3/Y AND2X1_LOC_633/Y 0.01fF
C55435 OR2X1_LOC_62/B OR2X1_LOC_204/a_8_216# 0.01fF
C55436 OR2X1_LOC_95/Y AND2X1_LOC_374/Y 0.01fF
C55437 OR2X1_LOC_22/Y OR2X1_LOC_17/Y 0.01fF
C55438 OR2X1_LOC_276/a_8_216# OR2X1_LOC_203/Y 0.04fF
C55439 OR2X1_LOC_95/Y OR2X1_LOC_52/B 0.03fF
C55440 OR2X1_LOC_409/B AND2X1_LOC_637/Y 0.02fF
C55441 OR2X1_LOC_672/Y OR2X1_LOC_95/Y 0.01fF
C55442 OR2X1_LOC_3/Y D_INPUT_0 0.14fF
C55443 AND2X1_LOC_576/Y OR2X1_LOC_224/Y 0.03fF
C55444 AND2X1_LOC_462/a_8_24# OR2X1_LOC_27/Y 0.01fF
C55445 OR2X1_LOC_92/Y AND2X1_LOC_222/Y 0.03fF
C55446 AND2X1_LOC_554/B OR2X1_LOC_71/Y 0.61fF
C55447 OR2X1_LOC_154/A D_INPUT_1 0.87fF
C55448 OR2X1_LOC_726/A OR2X1_LOC_726/a_8_216# 0.02fF
C55449 AND2X1_LOC_436/Y OR2X1_LOC_13/B 0.00fF
C55450 AND2X1_LOC_59/Y AND2X1_LOC_72/B 0.02fF
C55451 OR2X1_LOC_828/a_8_216# OR2X1_LOC_198/A 0.12fF
C55452 OR2X1_LOC_405/A OR2X1_LOC_723/A 0.01fF
C55453 OR2X1_LOC_863/B OR2X1_LOC_532/B 0.01fF
C55454 OR2X1_LOC_74/A AND2X1_LOC_675/A 0.07fF
C55455 OR2X1_LOC_362/A OR2X1_LOC_844/B 0.03fF
C55456 VDD OR2X1_LOC_532/Y 0.20fF
C55457 OR2X1_LOC_59/Y OR2X1_LOC_437/A 4.71fF
C55458 OR2X1_LOC_278/A OR2X1_LOC_46/A 3.80fF
C55459 OR2X1_LOC_503/A OR2X1_LOC_419/Y 0.00fF
C55460 AND2X1_LOC_53/Y OR2X1_LOC_193/A 0.01fF
C55461 OR2X1_LOC_653/Y AND2X1_LOC_31/Y 0.08fF
C55462 OR2X1_LOC_47/Y OR2X1_LOC_585/A 0.79fF
C55463 OR2X1_LOC_151/A OR2X1_LOC_168/Y 0.47fF
C55464 VDD OR2X1_LOC_212/B 0.08fF
C55465 OR2X1_LOC_759/A AND2X1_LOC_793/a_8_24# 0.01fF
C55466 OR2X1_LOC_160/B OR2X1_LOC_308/Y 0.01fF
C55467 OR2X1_LOC_756/B OR2X1_LOC_303/B 0.03fF
C55468 OR2X1_LOC_835/Y OR2X1_LOC_19/B 0.10fF
C55469 AND2X1_LOC_116/Y AND2X1_LOC_660/A 0.45fF
C55470 AND2X1_LOC_580/B AND2X1_LOC_793/Y 0.02fF
C55471 OR2X1_LOC_92/Y OR2X1_LOC_423/Y 0.05fF
C55472 OR2X1_LOC_66/A OR2X1_LOC_388/a_8_216# 0.01fF
C55473 VDD OR2X1_LOC_130/Y 0.27fF
C55474 OR2X1_LOC_516/Y AND2X1_LOC_657/Y 0.05fF
C55475 OR2X1_LOC_832/a_8_216# OR2X1_LOC_390/B 0.00fF
C55476 AND2X1_LOC_388/Y AND2X1_LOC_539/Y 0.01fF
C55477 OR2X1_LOC_443/Y AND2X1_LOC_47/Y 0.09fF
C55478 OR2X1_LOC_168/B AND2X1_LOC_36/Y 0.10fF
C55479 OR2X1_LOC_516/Y AND2X1_LOC_469/B 0.01fF
C55480 OR2X1_LOC_778/A D_INPUT_1 0.08fF
C55481 OR2X1_LOC_711/B AND2X1_LOC_7/B 0.12fF
C55482 OR2X1_LOC_516/B OR2X1_LOC_142/Y 0.03fF
C55483 OR2X1_LOC_176/Y AND2X1_LOC_180/a_8_24# 0.09fF
C55484 OR2X1_LOC_578/a_8_216# OR2X1_LOC_549/A 0.03fF
C55485 OR2X1_LOC_485/A AND2X1_LOC_486/a_8_24# 0.05fF
C55486 OR2X1_LOC_138/A OR2X1_LOC_514/a_8_216# 0.47fF
C55487 AND2X1_LOC_97/a_8_24# OR2X1_LOC_13/B 0.01fF
C55488 OR2X1_LOC_698/Y AND2X1_LOC_793/a_8_24# 0.01fF
C55489 OR2X1_LOC_829/A OR2X1_LOC_16/A 0.30fF
C55490 AND2X1_LOC_287/B AND2X1_LOC_244/a_8_24# 0.20fF
C55491 OR2X1_LOC_516/Y AND2X1_LOC_733/Y 0.07fF
C55492 OR2X1_LOC_720/Y AND2X1_LOC_18/Y 0.03fF
C55493 AND2X1_LOC_562/a_36_24# OR2X1_LOC_604/A 0.01fF
C55494 AND2X1_LOC_564/B AND2X1_LOC_658/B 0.07fF
C55495 AND2X1_LOC_810/A AND2X1_LOC_566/B 0.00fF
C55496 AND2X1_LOC_64/Y AND2X1_LOC_92/Y 0.19fF
C55497 AND2X1_LOC_227/Y OR2X1_LOC_226/a_36_216# -0.00fF
C55498 OR2X1_LOC_322/Y OR2X1_LOC_323/a_36_216# 0.00fF
C55499 AND2X1_LOC_707/Y OR2X1_LOC_681/a_36_216# 0.00fF
C55500 OR2X1_LOC_176/a_8_216# AND2X1_LOC_568/B 0.11fF
C55501 AND2X1_LOC_3/Y OR2X1_LOC_559/a_8_216# 0.01fF
C55502 OR2X1_LOC_375/A OR2X1_LOC_366/Y 0.06fF
C55503 AND2X1_LOC_786/Y AND2X1_LOC_778/Y 0.02fF
C55504 OR2X1_LOC_196/Y VDD 0.12fF
C55505 OR2X1_LOC_64/Y OR2X1_LOC_85/a_8_216# 0.01fF
C55506 OR2X1_LOC_404/Y OR2X1_LOC_493/Y 0.10fF
C55507 VDD OR2X1_LOC_266/A 0.08fF
C55508 AND2X1_LOC_672/a_36_24# INPUT_1 0.01fF
C55509 OR2X1_LOC_64/Y OR2X1_LOC_419/Y 0.76fF
C55510 OR2X1_LOC_40/Y OR2X1_LOC_12/Y 0.16fF
C55511 OR2X1_LOC_363/B OR2X1_LOC_366/B 0.11fF
C55512 AND2X1_LOC_48/A OR2X1_LOC_214/B 0.07fF
C55513 AND2X1_LOC_831/Y AND2X1_LOC_655/a_8_24# 0.01fF
C55514 AND2X1_LOC_217/Y OR2X1_LOC_595/A 0.01fF
C55515 AND2X1_LOC_706/Y AND2X1_LOC_713/Y 0.02fF
C55516 OR2X1_LOC_753/A OR2X1_LOC_71/A 0.16fF
C55517 AND2X1_LOC_47/Y AND2X1_LOC_813/a_8_24# 0.02fF
C55518 AND2X1_LOC_251/a_36_24# OR2X1_LOC_580/A 0.00fF
C55519 OR2X1_LOC_8/Y OR2X1_LOC_821/Y 0.00fF
C55520 AND2X1_LOC_59/Y AND2X1_LOC_36/Y 3.20fF
C55521 OR2X1_LOC_158/A VDD 1.56fF
C55522 AND2X1_LOC_131/a_8_24# AND2X1_LOC_625/a_8_24# 0.23fF
C55523 OR2X1_LOC_756/B OR2X1_LOC_366/B 0.40fF
C55524 OR2X1_LOC_87/A OR2X1_LOC_771/B 0.18fF
C55525 OR2X1_LOC_157/a_8_216# D_INPUT_6 0.01fF
C55526 OR2X1_LOC_329/B AND2X1_LOC_809/a_8_24# 0.03fF
C55527 AND2X1_LOC_243/a_8_24# OR2X1_LOC_71/A 0.01fF
C55528 OR2X1_LOC_735/a_8_216# AND2X1_LOC_44/Y 0.01fF
C55529 OR2X1_LOC_18/Y OR2X1_LOC_767/Y 0.02fF
C55530 OR2X1_LOC_532/B OR2X1_LOC_76/a_36_216# 0.02fF
C55531 OR2X1_LOC_589/A AND2X1_LOC_434/Y 0.07fF
C55532 AND2X1_LOC_719/Y OR2X1_LOC_666/A 0.05fF
C55533 OR2X1_LOC_528/Y OR2X1_LOC_51/Y 0.03fF
C55534 AND2X1_LOC_505/a_36_24# AND2X1_LOC_18/Y 0.01fF
C55535 OR2X1_LOC_269/B OR2X1_LOC_199/B 0.06fF
C55536 OR2X1_LOC_39/A AND2X1_LOC_590/a_8_24# 0.02fF
C55537 OR2X1_LOC_736/A OR2X1_LOC_342/A 0.01fF
C55538 OR2X1_LOC_87/A OR2X1_LOC_776/A 0.16fF
C55539 OR2X1_LOC_696/A OR2X1_LOC_91/Y 0.10fF
C55540 AND2X1_LOC_19/a_8_24# OR2X1_LOC_771/B 0.16fF
C55541 OR2X1_LOC_70/Y OR2X1_LOC_437/A 0.07fF
C55542 OR2X1_LOC_45/B AND2X1_LOC_486/Y 0.03fF
C55543 VDD OR2X1_LOC_450/B 0.21fF
C55544 OR2X1_LOC_51/Y OR2X1_LOC_583/Y 0.01fF
C55545 AND2X1_LOC_495/a_8_24# AND2X1_LOC_36/Y 0.01fF
C55546 OR2X1_LOC_121/Y OR2X1_LOC_274/Y 0.10fF
C55547 AND2X1_LOC_392/A OR2X1_LOC_56/A 0.21fF
C55548 OR2X1_LOC_440/B AND2X1_LOC_437/a_8_24# 0.01fF
C55549 AND2X1_LOC_807/B OR2X1_LOC_56/A 0.03fF
C55550 AND2X1_LOC_41/A OR2X1_LOC_726/A 0.18fF
C55551 INPUT_0 AND2X1_LOC_207/B 0.21fF
C55552 OR2X1_LOC_526/Y OR2X1_LOC_744/A 0.14fF
C55553 AND2X1_LOC_658/A AND2X1_LOC_658/Y 0.00fF
C55554 OR2X1_LOC_837/B AND2X1_LOC_415/a_8_24# 0.28fF
C55555 AND2X1_LOC_514/Y OR2X1_LOC_437/A 0.01fF
C55556 OR2X1_LOC_833/a_36_216# OR2X1_LOC_549/A 0.01fF
C55557 AND2X1_LOC_794/B OR2X1_LOC_594/Y 0.50fF
C55558 OR2X1_LOC_177/Y AND2X1_LOC_717/Y 0.03fF
C55559 INPUT_0 OR2X1_LOC_66/A 0.11fF
C55560 OR2X1_LOC_585/Y AND2X1_LOC_637/a_8_24# 0.02fF
C55561 OR2X1_LOC_161/A AND2X1_LOC_627/a_8_24# 0.17fF
C55562 OR2X1_LOC_857/B AND2X1_LOC_690/a_8_24# 0.01fF
C55563 VDD AND2X1_LOC_98/Y 0.27fF
C55564 OR2X1_LOC_166/Y AND2X1_LOC_434/Y 0.16fF
C55565 OR2X1_LOC_148/a_8_216# OR2X1_LOC_161/A 0.01fF
C55566 OR2X1_LOC_56/Y OR2X1_LOC_44/Y 0.00fF
C55567 OR2X1_LOC_703/A AND2X1_LOC_323/a_36_24# 0.01fF
C55568 OR2X1_LOC_337/A OR2X1_LOC_212/A 0.01fF
C55569 OR2X1_LOC_506/A OR2X1_LOC_435/A 0.36fF
C55570 AND2X1_LOC_434/a_36_24# OR2X1_LOC_59/Y 0.00fF
C55571 OR2X1_LOC_762/a_8_216# D_INPUT_6 0.05fF
C55572 OR2X1_LOC_114/Y OR2X1_LOC_392/B 0.49fF
C55573 AND2X1_LOC_22/Y OR2X1_LOC_720/A 0.08fF
C55574 OR2X1_LOC_325/B OR2X1_LOC_502/A 0.06fF
C55575 AND2X1_LOC_572/a_8_24# AND2X1_LOC_361/A 0.03fF
C55576 AND2X1_LOC_512/Y OR2X1_LOC_51/Y 0.01fF
C55577 OR2X1_LOC_510/Y OR2X1_LOC_161/B 0.13fF
C55578 OR2X1_LOC_227/Y OR2X1_LOC_560/A 0.34fF
C55579 OR2X1_LOC_325/A VDD 0.21fF
C55580 AND2X1_LOC_734/Y AND2X1_LOC_658/A 0.07fF
C55581 OR2X1_LOC_323/A AND2X1_LOC_717/B 0.00fF
C55582 VDD OR2X1_LOC_103/Y 0.24fF
C55583 AND2X1_LOC_720/Y VDD 0.24fF
C55584 AND2X1_LOC_706/Y AND2X1_LOC_436/B 0.02fF
C55585 AND2X1_LOC_534/a_36_24# OR2X1_LOC_161/A 0.00fF
C55586 OR2X1_LOC_158/A AND2X1_LOC_274/a_8_24# 0.01fF
C55587 OR2X1_LOC_59/Y OR2X1_LOC_755/Y 0.01fF
C55588 OR2X1_LOC_464/A OR2X1_LOC_787/B 0.02fF
C55589 VDD OR2X1_LOC_594/Y 0.12fF
C55590 AND2X1_LOC_500/a_8_24# AND2X1_LOC_242/a_8_24# 0.23fF
C55591 OR2X1_LOC_76/A OR2X1_LOC_301/a_8_216# 0.03fF
C55592 AND2X1_LOC_509/Y AND2X1_LOC_510/a_8_24# 0.00fF
C55593 AND2X1_LOC_457/a_8_24# OR2X1_LOC_44/Y 0.01fF
C55594 OR2X1_LOC_517/A AND2X1_LOC_218/Y 0.13fF
C55595 AND2X1_LOC_784/A AND2X1_LOC_358/Y 0.05fF
C55596 OR2X1_LOC_538/A AND2X1_LOC_167/a_8_24# 0.01fF
C55597 OR2X1_LOC_329/B OR2X1_LOC_164/Y 0.02fF
C55598 AND2X1_LOC_364/A AND2X1_LOC_326/B 0.02fF
C55599 OR2X1_LOC_103/a_8_216# VDD 0.21fF
C55600 AND2X1_LOC_56/B OR2X1_LOC_185/a_8_216# 0.07fF
C55601 OR2X1_LOC_19/B OR2X1_LOC_395/Y 0.06fF
C55602 OR2X1_LOC_696/A OR2X1_LOC_417/Y 0.07fF
C55603 OR2X1_LOC_423/a_8_216# OR2X1_LOC_428/A 0.01fF
C55604 VDD OR2X1_LOC_847/A 0.28fF
C55605 AND2X1_LOC_654/B AND2X1_LOC_434/Y 0.02fF
C55606 AND2X1_LOC_194/Y OR2X1_LOC_39/A 0.12fF
C55607 VDD OR2X1_LOC_447/A 0.21fF
C55608 OR2X1_LOC_810/A OR2X1_LOC_161/B 0.10fF
C55609 OR2X1_LOC_375/A OR2X1_LOC_786/A 0.01fF
C55610 VDD OR2X1_LOC_288/a_8_216# 0.00fF
C55611 OR2X1_LOC_307/a_8_216# OR2X1_LOC_161/B 0.06fF
C55612 AND2X1_LOC_22/Y OR2X1_LOC_333/B 0.01fF
C55613 OR2X1_LOC_114/B OR2X1_LOC_128/B 0.39fF
C55614 OR2X1_LOC_756/B OR2X1_LOC_105/a_8_216# 0.05fF
C55615 AND2X1_LOC_724/Y OR2X1_LOC_619/Y 0.14fF
C55616 OR2X1_LOC_696/A OR2X1_LOC_311/Y 0.07fF
C55617 OR2X1_LOC_528/Y OR2X1_LOC_680/A 0.25fF
C55618 OR2X1_LOC_121/a_8_216# OR2X1_LOC_574/A 0.14fF
C55619 AND2X1_LOC_857/a_8_24# OR2X1_LOC_12/Y 0.02fF
C55620 AND2X1_LOC_722/A OR2X1_LOC_594/a_8_216# 0.05fF
C55621 OR2X1_LOC_32/B OR2X1_LOC_600/A 0.07fF
C55622 OR2X1_LOC_40/a_8_216# OR2X1_LOC_25/Y 0.04fF
C55623 OR2X1_LOC_102/a_8_216# OR2X1_LOC_248/Y 0.04fF
C55624 AND2X1_LOC_367/A OR2X1_LOC_92/Y 0.00fF
C55625 AND2X1_LOC_639/a_8_24# OR2X1_LOC_428/A 0.02fF
C55626 VDD AND2X1_LOC_577/Y 0.01fF
C55627 OR2X1_LOC_7/A OR2X1_LOC_12/Y 0.90fF
C55628 OR2X1_LOC_184/Y OR2X1_LOC_437/A 0.00fF
C55629 OR2X1_LOC_479/Y AND2X1_LOC_44/Y 0.03fF
C55630 OR2X1_LOC_7/A OR2X1_LOC_766/Y 0.01fF
C55631 AND2X1_LOC_585/a_8_24# AND2X1_LOC_3/Y 0.01fF
C55632 OR2X1_LOC_303/A OR2X1_LOC_620/Y 0.01fF
C55633 AND2X1_LOC_555/Y OR2X1_LOC_54/Y 0.07fF
C55634 OR2X1_LOC_158/A OR2X1_LOC_251/Y 0.02fF
C55635 OR2X1_LOC_40/Y AND2X1_LOC_650/Y 0.21fF
C55636 AND2X1_LOC_715/Y OR2X1_LOC_417/Y 0.12fF
C55637 OR2X1_LOC_644/B OR2X1_LOC_598/Y 0.02fF
C55638 OR2X1_LOC_821/a_36_216# OR2X1_LOC_74/A 0.03fF
C55639 OR2X1_LOC_624/A OR2X1_LOC_78/B 0.03fF
C55640 OR2X1_LOC_502/A AND2X1_LOC_615/a_8_24# 0.01fF
C55641 OR2X1_LOC_744/A OR2X1_LOC_433/Y 0.01fF
C55642 VDD OR2X1_LOC_685/B 0.21fF
C55643 OR2X1_LOC_437/Y OR2X1_LOC_437/A 0.12fF
C55644 OR2X1_LOC_51/Y AND2X1_LOC_342/Y 0.07fF
C55645 OR2X1_LOC_502/A AND2X1_LOC_423/a_8_24# 0.04fF
C55646 OR2X1_LOC_844/Y OR2X1_LOC_392/B 0.07fF
C55647 OR2X1_LOC_86/a_8_216# AND2X1_LOC_243/Y 0.04fF
C55648 AND2X1_LOC_719/Y OR2X1_LOC_312/Y 0.01fF
C55649 AND2X1_LOC_365/A AND2X1_LOC_434/Y 0.01fF
C55650 OR2X1_LOC_858/A AND2X1_LOC_272/a_8_24# 0.05fF
C55651 AND2X1_LOC_715/Y OR2X1_LOC_311/Y 0.01fF
C55652 OR2X1_LOC_640/Y OR2X1_LOC_462/B 0.01fF
C55653 OR2X1_LOC_3/Y AND2X1_LOC_771/B 0.01fF
C55654 OR2X1_LOC_441/Y AND2X1_LOC_808/a_8_24# 0.04fF
C55655 OR2X1_LOC_40/Y AND2X1_LOC_175/a_8_24# 0.02fF
C55656 OR2X1_LOC_843/a_8_216# OR2X1_LOC_349/A 0.40fF
C55657 AND2X1_LOC_47/Y OR2X1_LOC_605/Y 0.02fF
C55658 OR2X1_LOC_306/Y INPUT_0 0.07fF
C55659 AND2X1_LOC_576/Y AND2X1_LOC_558/a_8_24# 0.00fF
C55660 AND2X1_LOC_633/Y AND2X1_LOC_201/Y 0.06fF
C55661 AND2X1_LOC_47/Y AND2X1_LOC_763/B 0.01fF
C55662 OR2X1_LOC_40/Y OR2X1_LOC_239/a_8_216# 0.14fF
C55663 OR2X1_LOC_22/Y AND2X1_LOC_473/Y 0.10fF
C55664 OR2X1_LOC_663/A OR2X1_LOC_185/A 0.13fF
C55665 OR2X1_LOC_122/Y OR2X1_LOC_67/A 0.01fF
C55666 AND2X1_LOC_70/Y OR2X1_LOC_205/a_8_216# 0.01fF
C55667 OR2X1_LOC_86/A OR2X1_LOC_13/B 0.08fF
C55668 AND2X1_LOC_722/A AND2X1_LOC_468/B 0.94fF
C55669 AND2X1_LOC_715/Y OR2X1_LOC_601/a_8_216# 0.06fF
C55670 OR2X1_LOC_160/A OR2X1_LOC_334/B 0.14fF
C55671 OR2X1_LOC_3/Y OR2X1_LOC_131/A 0.09fF
C55672 OR2X1_LOC_22/Y AND2X1_LOC_287/B 0.04fF
C55673 AND2X1_LOC_580/A AND2X1_LOC_549/a_8_24# 0.01fF
C55674 OR2X1_LOC_235/B AND2X1_LOC_63/a_8_24# 0.11fF
C55675 OR2X1_LOC_22/Y OR2X1_LOC_816/A 0.03fF
C55676 OR2X1_LOC_696/A D_INPUT_3 0.11fF
C55677 AND2X1_LOC_12/Y OR2X1_LOC_274/Y 0.00fF
C55678 OR2X1_LOC_624/A OR2X1_LOC_721/Y 0.10fF
C55679 OR2X1_LOC_51/Y AND2X1_LOC_105/a_8_24# 0.01fF
C55680 OR2X1_LOC_43/A AND2X1_LOC_434/Y 1.06fF
C55681 AND2X1_LOC_512/Y OR2X1_LOC_680/A 0.02fF
C55682 OR2X1_LOC_210/B OR2X1_LOC_803/A 0.01fF
C55683 AND2X1_LOC_81/B AND2X1_LOC_41/A 0.05fF
C55684 OR2X1_LOC_177/Y OR2X1_LOC_64/Y 0.22fF
C55685 OR2X1_LOC_744/A AND2X1_LOC_661/A 0.13fF
C55686 AND2X1_LOC_12/Y OR2X1_LOC_392/A 0.01fF
C55687 OR2X1_LOC_43/A AND2X1_LOC_219/Y 0.07fF
C55688 OR2X1_LOC_467/A OR2X1_LOC_449/a_36_216# 0.00fF
C55689 OR2X1_LOC_502/A OR2X1_LOC_405/Y 0.03fF
C55690 OR2X1_LOC_190/A AND2X1_LOC_3/Y 0.01fF
C55691 OR2X1_LOC_753/A OR2X1_LOC_59/Y 0.07fF
C55692 AND2X1_LOC_41/A OR2X1_LOC_358/B 0.03fF
C55693 OR2X1_LOC_154/A OR2X1_LOC_274/a_36_216# 0.03fF
C55694 OR2X1_LOC_600/A OR2X1_LOC_371/Y 0.07fF
C55695 OR2X1_LOC_121/B AND2X1_LOC_65/A 0.03fF
C55696 AND2X1_LOC_95/Y OR2X1_LOC_620/Y 0.87fF
C55697 OR2X1_LOC_756/B AND2X1_LOC_56/B 0.15fF
C55698 OR2X1_LOC_844/Y OR2X1_LOC_113/B 0.03fF
C55699 AND2X1_LOC_40/Y OR2X1_LOC_807/A 0.12fF
C55700 OR2X1_LOC_405/A OR2X1_LOC_231/A 0.03fF
C55701 AND2X1_LOC_716/Y AND2X1_LOC_655/A 0.10fF
C55702 OR2X1_LOC_135/Y OR2X1_LOC_46/A 0.08fF
C55703 OR2X1_LOC_625/Y OR2X1_LOC_628/a_36_216# 0.00fF
C55704 AND2X1_LOC_737/Y AND2X1_LOC_807/Y 0.33fF
C55705 AND2X1_LOC_576/Y AND2X1_LOC_508/A 0.03fF
C55706 OR2X1_LOC_325/a_8_216# AND2X1_LOC_59/Y 0.04fF
C55707 AND2X1_LOC_474/A OR2X1_LOC_26/Y 0.02fF
C55708 AND2X1_LOC_367/A OR2X1_LOC_271/Y 0.03fF
C55709 AND2X1_LOC_554/B OR2X1_LOC_426/B 0.03fF
C55710 AND2X1_LOC_52/a_36_24# OR2X1_LOC_375/A 0.00fF
C55711 OR2X1_LOC_508/A AND2X1_LOC_81/B 0.01fF
C55712 OR2X1_LOC_319/a_8_216# OR2X1_LOC_161/A 0.03fF
C55713 OR2X1_LOC_479/Y OR2X1_LOC_785/a_8_216# 0.41fF
C55714 OR2X1_LOC_756/B AND2X1_LOC_8/Y 0.01fF
C55715 OR2X1_LOC_68/B OR2X1_LOC_580/A 0.03fF
C55716 AND2X1_LOC_654/Y AND2X1_LOC_655/A 0.10fF
C55717 OR2X1_LOC_604/A OR2X1_LOC_64/Y 0.24fF
C55718 OR2X1_LOC_377/A OR2X1_LOC_240/B 0.08fF
C55719 OR2X1_LOC_123/a_8_216# OR2X1_LOC_123/B 0.06fF
C55720 AND2X1_LOC_212/A OR2X1_LOC_22/Y 0.03fF
C55721 OR2X1_LOC_435/B OR2X1_LOC_810/A 0.07fF
C55722 AND2X1_LOC_53/a_36_24# OR2X1_LOC_375/A 0.00fF
C55723 OR2X1_LOC_51/Y AND2X1_LOC_483/a_8_24# 0.14fF
C55724 OR2X1_LOC_154/A OR2X1_LOC_737/A 0.07fF
C55725 OR2X1_LOC_648/B OR2X1_LOC_750/A 0.05fF
C55726 AND2X1_LOC_474/A OR2X1_LOC_89/A 0.03fF
C55727 OR2X1_LOC_644/B AND2X1_LOC_40/Y 0.01fF
C55728 AND2X1_LOC_700/a_36_24# OR2X1_LOC_705/Y 0.00fF
C55729 OR2X1_LOC_377/A OR2X1_LOC_161/A 0.03fF
C55730 OR2X1_LOC_808/a_8_216# OR2X1_LOC_87/A 0.01fF
C55731 OR2X1_LOC_532/B OR2X1_LOC_294/Y 0.02fF
C55732 OR2X1_LOC_139/A OR2X1_LOC_506/B 0.03fF
C55733 AND2X1_LOC_564/B OR2X1_LOC_47/Y 0.01fF
C55734 OR2X1_LOC_451/B AND2X1_LOC_582/B 0.01fF
C55735 AND2X1_LOC_326/A OR2X1_LOC_426/B 0.04fF
C55736 OR2X1_LOC_405/A OR2X1_LOC_130/A 0.19fF
C55737 AND2X1_LOC_729/Y AND2X1_LOC_621/Y 0.03fF
C55738 OR2X1_LOC_624/A OR2X1_LOC_375/A 0.03fF
C55739 AND2X1_LOC_143/a_8_24# OR2X1_LOC_585/A 0.05fF
C55740 AND2X1_LOC_720/Y OR2X1_LOC_251/Y 0.01fF
C55741 OR2X1_LOC_160/B OR2X1_LOC_19/B 0.04fF
C55742 OR2X1_LOC_177/Y OR2X1_LOC_417/A 0.05fF
C55743 OR2X1_LOC_427/A OR2X1_LOC_6/A 0.16fF
C55744 OR2X1_LOC_154/A AND2X1_LOC_95/Y 0.18fF
C55745 AND2X1_LOC_11/Y OR2X1_LOC_87/A 0.02fF
C55746 OR2X1_LOC_45/B AND2X1_LOC_660/A 0.03fF
C55747 OR2X1_LOC_496/Y OR2X1_LOC_495/Y 0.05fF
C55748 AND2X1_LOC_514/Y AND2X1_LOC_715/A 0.03fF
C55749 OR2X1_LOC_697/Y OR2X1_LOC_743/A 0.23fF
C55750 AND2X1_LOC_589/a_8_24# OR2X1_LOC_435/B 0.03fF
C55751 OR2X1_LOC_725/B OR2X1_LOC_269/B 0.00fF
C55752 AND2X1_LOC_711/Y OR2X1_LOC_755/Y 0.01fF
C55753 AND2X1_LOC_362/B OR2X1_LOC_71/Y 0.03fF
C55754 OR2X1_LOC_606/a_8_216# OR2X1_LOC_66/A 0.01fF
C55755 OR2X1_LOC_845/A OR2X1_LOC_266/A 1.12fF
C55756 OR2X1_LOC_864/A OR2X1_LOC_653/Y 0.07fF
C55757 OR2X1_LOC_364/A OR2X1_LOC_185/A 0.07fF
C55758 OR2X1_LOC_516/A OR2X1_LOC_680/A 0.03fF
C55759 OR2X1_LOC_422/a_8_216# OR2X1_LOC_7/A 0.03fF
C55760 OR2X1_LOC_185/Y OR2X1_LOC_185/A 0.03fF
C55761 AND2X1_LOC_511/a_8_24# AND2X1_LOC_47/Y 0.01fF
C55762 AND2X1_LOC_576/Y OR2X1_LOC_18/Y 0.00fF
C55763 OR2X1_LOC_158/A OR2X1_LOC_256/A 0.01fF
C55764 OR2X1_LOC_823/Y OR2X1_LOC_6/A 0.01fF
C55765 OR2X1_LOC_51/Y OR2X1_LOC_54/Y 0.06fF
C55766 OR2X1_LOC_203/Y OR2X1_LOC_161/A 0.04fF
C55767 OR2X1_LOC_673/B OR2X1_LOC_673/A 0.04fF
C55768 OR2X1_LOC_833/a_8_216# AND2X1_LOC_42/B 0.07fF
C55769 OR2X1_LOC_490/Y OR2X1_LOC_92/Y 0.10fF
C55770 OR2X1_LOC_92/Y OR2X1_LOC_74/A 0.07fF
C55771 OR2X1_LOC_532/B OR2X1_LOC_733/A 0.01fF
C55772 AND2X1_LOC_583/a_36_24# AND2X1_LOC_1/Y 0.00fF
C55773 OR2X1_LOC_625/Y OR2X1_LOC_585/A 0.01fF
C55774 AND2X1_LOC_394/a_8_24# OR2X1_LOC_673/Y 0.02fF
C55775 OR2X1_LOC_50/a_8_216# INPUT_7 0.09fF
C55776 OR2X1_LOC_604/A OR2X1_LOC_417/A 0.17fF
C55777 OR2X1_LOC_660/B AND2X1_LOC_8/Y 0.01fF
C55778 OR2X1_LOC_201/A OR2X1_LOC_473/Y 0.05fF
C55779 OR2X1_LOC_831/A OR2X1_LOC_223/A 0.01fF
C55780 AND2X1_LOC_578/A AND2X1_LOC_833/a_8_24# 0.01fF
C55781 AND2X1_LOC_59/Y OR2X1_LOC_346/B 0.37fF
C55782 AND2X1_LOC_715/a_8_24# AND2X1_LOC_354/a_8_24# 0.23fF
C55783 OR2X1_LOC_597/Y OR2X1_LOC_16/A 0.01fF
C55784 OR2X1_LOC_526/Y OR2X1_LOC_31/Y 0.01fF
C55785 OR2X1_LOC_654/A AND2X1_LOC_290/a_36_24# 0.01fF
C55786 OR2X1_LOC_271/a_8_216# OR2X1_LOC_6/A 0.01fF
C55787 AND2X1_LOC_41/A OR2X1_LOC_196/B 0.07fF
C55788 OR2X1_LOC_375/A OR2X1_LOC_552/a_8_216# 0.02fF
C55789 AND2X1_LOC_593/Y OR2X1_LOC_89/A 0.03fF
C55790 OR2X1_LOC_778/A OR2X1_LOC_737/A 0.02fF
C55791 OR2X1_LOC_3/Y OR2X1_LOC_399/A 0.01fF
C55792 OR2X1_LOC_591/A OR2X1_LOC_44/Y 0.01fF
C55793 OR2X1_LOC_694/a_8_216# OR2X1_LOC_7/A 0.03fF
C55794 OR2X1_LOC_26/Y OR2X1_LOC_85/A 0.13fF
C55795 OR2X1_LOC_774/Y OR2X1_LOC_848/B 0.04fF
C55796 OR2X1_LOC_835/B OR2X1_LOC_269/B 0.15fF
C55797 AND2X1_LOC_358/Y AND2X1_LOC_643/a_8_24# 0.20fF
C55798 AND2X1_LOC_845/Y OR2X1_LOC_59/Y 0.01fF
C55799 AND2X1_LOC_56/B OR2X1_LOC_76/Y 0.05fF
C55800 OR2X1_LOC_318/a_36_216# OR2X1_LOC_804/A 0.00fF
C55801 OR2X1_LOC_485/A AND2X1_LOC_436/B 0.02fF
C55802 OR2X1_LOC_287/B OR2X1_LOC_664/Y 0.03fF
C55803 AND2X1_LOC_41/A AND2X1_LOC_692/a_8_24# 0.02fF
C55804 OR2X1_LOC_108/Y OR2X1_LOC_224/Y 0.01fF
C55805 OR2X1_LOC_490/Y OR2X1_LOC_65/B 0.02fF
C55806 OR2X1_LOC_465/a_8_216# OR2X1_LOC_465/B 0.01fF
C55807 OR2X1_LOC_91/Y OR2X1_LOC_89/a_8_216# 0.04fF
C55808 OR2X1_LOC_74/A OR2X1_LOC_65/B 0.06fF
C55809 OR2X1_LOC_669/A OR2X1_LOC_669/Y 0.01fF
C55810 AND2X1_LOC_302/a_36_24# OR2X1_LOC_52/B 0.00fF
C55811 AND2X1_LOC_578/A AND2X1_LOC_624/A 0.07fF
C55812 AND2X1_LOC_721/Y AND2X1_LOC_657/A 0.02fF
C55813 OR2X1_LOC_744/A AND2X1_LOC_810/Y 0.24fF
C55814 AND2X1_LOC_850/a_8_24# OR2X1_LOC_64/Y 0.17fF
C55815 AND2X1_LOC_650/Y OR2X1_LOC_7/A 0.02fF
C55816 AND2X1_LOC_327/a_8_24# OR2X1_LOC_18/Y 0.09fF
C55817 AND2X1_LOC_44/Y OR2X1_LOC_259/B 0.04fF
C55818 OR2X1_LOC_259/B OR2X1_LOC_555/a_8_216# 0.47fF
C55819 OR2X1_LOC_634/A AND2X1_LOC_47/Y 0.02fF
C55820 OR2X1_LOC_377/A AND2X1_LOC_51/Y 0.57fF
C55821 OR2X1_LOC_190/A OR2X1_LOC_270/Y 0.03fF
C55822 OR2X1_LOC_232/a_36_216# OR2X1_LOC_753/A 0.00fF
C55823 OR2X1_LOC_362/A OR2X1_LOC_493/Y 0.03fF
C55824 AND2X1_LOC_44/Y OR2X1_LOC_68/B 10.49fF
C55825 OR2X1_LOC_502/A D_INPUT_0 0.10fF
C55826 AND2X1_LOC_211/B AND2X1_LOC_853/Y 0.44fF
C55827 OR2X1_LOC_461/Y AND2X1_LOC_824/B 0.01fF
C55828 AND2X1_LOC_520/Y OR2X1_LOC_46/A 0.31fF
C55829 AND2X1_LOC_94/a_8_24# OR2X1_LOC_54/Y 0.02fF
C55830 AND2X1_LOC_40/Y AND2X1_LOC_53/Y 0.08fF
C55831 OR2X1_LOC_223/A OR2X1_LOC_795/B 0.01fF
C55832 INPUT_3 OR2X1_LOC_19/B 0.36fF
C55833 OR2X1_LOC_45/Y OR2X1_LOC_22/Y 0.41fF
C55834 OR2X1_LOC_306/Y OR2X1_LOC_64/Y 0.02fF
C55835 OR2X1_LOC_158/A OR2X1_LOC_163/Y 0.09fF
C55836 OR2X1_LOC_808/A OR2X1_LOC_440/A 0.02fF
C55837 D_INPUT_3 AND2X1_LOC_819/a_8_24# 0.05fF
C55838 OR2X1_LOC_677/a_8_216# AND2X1_LOC_796/Y 0.01fF
C55839 OR2X1_LOC_686/a_8_216# OR2X1_LOC_451/B 0.01fF
C55840 OR2X1_LOC_335/Y OR2X1_LOC_223/A 0.01fF
C55841 OR2X1_LOC_58/Y OR2X1_LOC_598/A 0.03fF
C55842 AND2X1_LOC_36/Y AND2X1_LOC_762/a_8_24# 0.01fF
C55843 OR2X1_LOC_203/Y AND2X1_LOC_51/Y 0.07fF
C55844 OR2X1_LOC_377/A OR2X1_LOC_836/Y 0.05fF
C55845 OR2X1_LOC_264/Y OR2X1_LOC_218/Y 0.09fF
C55846 OR2X1_LOC_286/a_8_216# OR2X1_LOC_286/Y 0.01fF
C55847 OR2X1_LOC_529/Y OR2X1_LOC_485/A 0.04fF
C55848 OR2X1_LOC_375/A OR2X1_LOC_54/Y 0.05fF
C55849 AND2X1_LOC_390/B AND2X1_LOC_645/A 0.53fF
C55850 OR2X1_LOC_482/Y AND2X1_LOC_657/A 0.07fF
C55851 AND2X1_LOC_147/Y AND2X1_LOC_148/Y 0.01fF
C55852 OR2X1_LOC_461/a_8_216# OR2X1_LOC_598/A 0.01fF
C55853 AND2X1_LOC_33/Y D_INPUT_0 0.02fF
C55854 AND2X1_LOC_303/B AND2X1_LOC_537/Y 0.06fF
C55855 OR2X1_LOC_189/Y AND2X1_LOC_797/A 0.14fF
C55856 OR2X1_LOC_600/A AND2X1_LOC_222/Y 0.03fF
C55857 OR2X1_LOC_429/Y OR2X1_LOC_17/Y 0.03fF
C55858 AND2X1_LOC_851/B OR2X1_LOC_495/Y 0.35fF
C55859 AND2X1_LOC_40/Y OR2X1_LOC_223/A 0.05fF
C55860 AND2X1_LOC_335/Y AND2X1_LOC_222/Y 0.01fF
C55861 OR2X1_LOC_447/Y OR2X1_LOC_375/A 0.03fF
C55862 OR2X1_LOC_31/Y OR2X1_LOC_433/Y 0.49fF
C55863 AND2X1_LOC_811/Y AND2X1_LOC_811/B 0.29fF
C55864 OR2X1_LOC_371/Y OR2X1_LOC_372/a_8_216# 0.43fF
C55865 AND2X1_LOC_41/A OR2X1_LOC_66/Y 0.00fF
C55866 OR2X1_LOC_696/Y OR2X1_LOC_743/A 0.02fF
C55867 AND2X1_LOC_663/B OR2X1_LOC_757/Y 0.01fF
C55868 OR2X1_LOC_549/A OR2X1_LOC_366/Y 0.02fF
C55869 OR2X1_LOC_823/a_36_216# D_INPUT_3 0.00fF
C55870 OR2X1_LOC_276/B OR2X1_LOC_269/a_8_216# 0.01fF
C55871 OR2X1_LOC_634/A OR2X1_LOC_598/A 0.56fF
C55872 OR2X1_LOC_72/a_8_216# OR2X1_LOC_265/Y 0.03fF
C55873 OR2X1_LOC_114/Y OR2X1_LOC_532/B 0.03fF
C55874 OR2X1_LOC_742/B OR2X1_LOC_742/a_8_216# 0.01fF
C55875 OR2X1_LOC_174/A OR2X1_LOC_358/A 0.04fF
C55876 AND2X1_LOC_640/Y OR2X1_LOC_416/Y 0.01fF
C55877 AND2X1_LOC_476/A OR2X1_LOC_265/Y 0.07fF
C55878 OR2X1_LOC_516/Y AND2X1_LOC_804/A 0.99fF
C55879 OR2X1_LOC_3/Y AND2X1_LOC_687/A 0.04fF
C55880 OR2X1_LOC_696/A OR2X1_LOC_184/a_36_216# 0.00fF
C55881 AND2X1_LOC_139/B AND2X1_LOC_655/a_8_24# 0.20fF
C55882 AND2X1_LOC_719/Y OR2X1_LOC_13/B 0.10fF
C55883 OR2X1_LOC_845/a_8_216# AND2X1_LOC_47/Y 0.02fF
C55884 OR2X1_LOC_70/Y OR2X1_LOC_684/Y 0.01fF
C55885 AND2X1_LOC_810/Y AND2X1_LOC_840/B 0.10fF
C55886 OR2X1_LOC_633/Y AND2X1_LOC_6/a_8_24# 0.00fF
C55887 OR2X1_LOC_92/Y AND2X1_LOC_647/Y 0.01fF
C55888 OR2X1_LOC_557/A OR2X1_LOC_814/A 0.06fF
C55889 OR2X1_LOC_31/Y AND2X1_LOC_654/a_8_24# 0.02fF
C55890 OR2X1_LOC_458/a_8_216# AND2X1_LOC_31/Y 0.01fF
C55891 AND2X1_LOC_40/Y AND2X1_LOC_609/a_8_24# 0.01fF
C55892 AND2X1_LOC_658/B OR2X1_LOC_437/A 0.12fF
C55893 AND2X1_LOC_48/A OR2X1_LOC_193/A 0.02fF
C55894 INPUT_4 OR2X1_LOC_50/a_8_216# 0.01fF
C55895 AND2X1_LOC_10/a_8_24# OR2X1_LOC_62/B 0.09fF
C55896 OR2X1_LOC_89/A OR2X1_LOC_226/Y 0.21fF
C55897 OR2X1_LOC_333/B OR2X1_LOC_434/A 0.01fF
C55898 OR2X1_LOC_39/Y OR2X1_LOC_39/a_36_216# 0.00fF
C55899 OR2X1_LOC_84/Y OR2X1_LOC_375/A 0.00fF
C55900 OR2X1_LOC_633/Y OR2X1_LOC_99/A 0.03fF
C55901 AND2X1_LOC_856/B OR2X1_LOC_46/A 0.16fF
C55902 OR2X1_LOC_280/Y OR2X1_LOC_95/Y 0.13fF
C55903 AND2X1_LOC_102/a_8_24# OR2X1_LOC_62/A 0.04fF
C55904 OR2X1_LOC_532/B OR2X1_LOC_201/Y 0.01fF
C55905 AND2X1_LOC_863/A OR2X1_LOC_46/A 0.33fF
C55906 OR2X1_LOC_52/Y OR2X1_LOC_7/Y 0.36fF
C55907 OR2X1_LOC_65/B AND2X1_LOC_647/Y 0.02fF
C55908 OR2X1_LOC_602/a_8_216# AND2X1_LOC_47/Y 0.00fF
C55909 OR2X1_LOC_22/Y AND2X1_LOC_727/A 0.03fF
C55910 OR2X1_LOC_185/A OR2X1_LOC_552/A 0.00fF
C55911 OR2X1_LOC_85/A AND2X1_LOC_202/a_8_24# 0.09fF
C55912 AND2X1_LOC_825/a_36_24# OR2X1_LOC_46/A 0.00fF
C55913 AND2X1_LOC_95/Y OR2X1_LOC_560/A 0.02fF
C55914 OR2X1_LOC_177/Y AND2X1_LOC_544/Y 0.80fF
C55915 OR2X1_LOC_19/B OR2X1_LOC_244/A 0.12fF
C55916 AND2X1_LOC_550/A OR2X1_LOC_152/A 0.12fF
C55917 AND2X1_LOC_48/A D_INPUT_0 0.05fF
C55918 AND2X1_LOC_624/A OR2X1_LOC_746/Y 0.14fF
C55919 OR2X1_LOC_494/a_36_216# OR2X1_LOC_437/A 0.00fF
C55920 AND2X1_LOC_3/Y OR2X1_LOC_214/B 0.03fF
C55921 OR2X1_LOC_185/A OR2X1_LOC_578/B 0.21fF
C55922 AND2X1_LOC_31/Y AND2X1_LOC_272/a_8_24# 0.00fF
C55923 D_INPUT_3 AND2X1_LOC_663/B 0.03fF
C55924 OR2X1_LOC_475/Y OR2X1_LOC_223/A 0.00fF
C55925 AND2X1_LOC_259/Y OR2X1_LOC_257/Y 0.01fF
C55926 OR2X1_LOC_364/B OR2X1_LOC_97/A 0.02fF
C55927 AND2X1_LOC_43/B OR2X1_LOC_715/a_36_216# 0.00fF
C55928 OR2X1_LOC_375/A OR2X1_LOC_513/a_8_216# 0.01fF
C55929 AND2X1_LOC_727/Y OR2X1_LOC_40/Y 0.03fF
C55930 AND2X1_LOC_357/a_8_24# OR2X1_LOC_437/A 0.04fF
C55931 AND2X1_LOC_32/a_8_24# AND2X1_LOC_31/Y 0.12fF
C55932 OR2X1_LOC_22/Y OR2X1_LOC_95/Y 0.23fF
C55933 AND2X1_LOC_544/Y OR2X1_LOC_745/a_8_216# 0.06fF
C55934 OR2X1_LOC_679/Y AND2X1_LOC_209/Y 0.80fF
C55935 OR2X1_LOC_214/A OR2X1_LOC_66/A 0.01fF
C55936 OR2X1_LOC_691/A OR2X1_LOC_857/B 0.01fF
C55937 AND2X1_LOC_562/a_8_24# VDD -0.00fF
C55938 AND2X1_LOC_41/A OR2X1_LOC_727/a_8_216# 0.19fF
C55939 OR2X1_LOC_620/Y OR2X1_LOC_788/B 0.03fF
C55940 OR2X1_LOC_623/B AND2X1_LOC_36/Y 0.03fF
C55941 OR2X1_LOC_715/B OR2X1_LOC_161/B 0.03fF
C55942 OR2X1_LOC_139/A AND2X1_LOC_18/Y 0.07fF
C55943 AND2X1_LOC_721/Y VDD 1.02fF
C55944 AND2X1_LOC_47/Y OR2X1_LOC_439/a_8_216# 0.01fF
C55945 OR2X1_LOC_201/a_8_216# OR2X1_LOC_532/B 0.02fF
C55946 OR2X1_LOC_508/a_8_216# OR2X1_LOC_151/A 0.05fF
C55947 AND2X1_LOC_7/B OR2X1_LOC_66/A 0.15fF
C55948 VDD OR2X1_LOC_474/B 0.06fF
C55949 AND2X1_LOC_167/a_8_24# OR2X1_LOC_356/B 0.25fF
C55950 OR2X1_LOC_618/Y D_INPUT_0 0.40fF
C55951 OR2X1_LOC_151/A OR2X1_LOC_486/Y 0.02fF
C55952 OR2X1_LOC_178/a_8_216# OR2X1_LOC_428/A 0.14fF
C55953 OR2X1_LOC_543/A OR2X1_LOC_161/B 0.03fF
C55954 AND2X1_LOC_655/A OR2X1_LOC_13/B 0.30fF
C55955 AND2X1_LOC_539/Y OR2X1_LOC_329/B 0.03fF
C55956 AND2X1_LOC_567/a_8_24# AND2X1_LOC_802/Y 0.01fF
C55957 AND2X1_LOC_535/Y AND2X1_LOC_810/B 0.19fF
C55958 OR2X1_LOC_635/A AND2X1_LOC_582/B 0.83fF
C55959 OR2X1_LOC_97/A AND2X1_LOC_70/Y 0.05fF
C55960 OR2X1_LOC_786/A OR2X1_LOC_549/A 0.02fF
C55961 OR2X1_LOC_736/A OR2X1_LOC_140/B 0.74fF
C55962 OR2X1_LOC_488/a_8_216# AND2X1_LOC_563/Y 0.01fF
C55963 AND2X1_LOC_91/B OR2X1_LOC_808/B 0.03fF
C55964 AND2X1_LOC_47/a_8_24# INPUT_6 0.04fF
C55965 OR2X1_LOC_158/A OR2X1_LOC_60/Y 0.01fF
C55966 OR2X1_LOC_154/A OR2X1_LOC_175/a_8_216# 0.04fF
C55967 OR2X1_LOC_202/a_36_216# AND2X1_LOC_31/Y 0.00fF
C55968 VDD OR2X1_LOC_482/Y 0.60fF
C55969 OR2X1_LOC_44/Y OR2X1_LOC_749/Y 0.01fF
C55970 OR2X1_LOC_97/A OR2X1_LOC_703/A 0.03fF
C55971 OR2X1_LOC_402/B AND2X1_LOC_82/Y 0.84fF
C55972 OR2X1_LOC_87/A OR2X1_LOC_593/B 0.01fF
C55973 OR2X1_LOC_532/B OR2X1_LOC_741/A 0.01fF
C55974 AND2X1_LOC_362/B OR2X1_LOC_426/B 0.40fF
C55975 OR2X1_LOC_631/a_8_216# OR2X1_LOC_140/B 0.01fF
C55976 OR2X1_LOC_834/a_8_216# AND2X1_LOC_44/Y 0.01fF
C55977 OR2X1_LOC_160/B AND2X1_LOC_110/Y 0.26fF
C55978 OR2X1_LOC_403/B OR2X1_LOC_771/B 0.14fF
C55979 OR2X1_LOC_51/Y OR2X1_LOC_765/Y 0.16fF
C55980 AND2X1_LOC_462/a_8_24# OR2X1_LOC_68/B 0.01fF
C55981 OR2X1_LOC_833/Y AND2X1_LOC_41/A 0.02fF
C55982 OR2X1_LOC_7/A OR2X1_LOC_248/A 0.03fF
C55983 AND2X1_LOC_364/Y OR2X1_LOC_589/A 0.31fF
C55984 OR2X1_LOC_78/A OR2X1_LOC_786/a_8_216# 0.01fF
C55985 OR2X1_LOC_45/B AND2X1_LOC_642/Y 0.01fF
C55986 D_INPUT_5 INPUT_7 0.06fF
C55987 OR2X1_LOC_95/Y OR2X1_LOC_387/a_8_216# 0.01fF
C55988 OR2X1_LOC_528/Y OR2X1_LOC_757/A 0.18fF
C55989 AND2X1_LOC_390/a_8_24# OR2X1_LOC_59/Y 0.08fF
C55990 AND2X1_LOC_471/Y AND2X1_LOC_477/Y 0.04fF
C55991 AND2X1_LOC_810/A OR2X1_LOC_92/Y 0.03fF
C55992 OR2X1_LOC_776/Y AND2X1_LOC_92/Y 0.03fF
C55993 AND2X1_LOC_43/a_8_24# AND2X1_LOC_36/Y 0.01fF
C55994 VDD OR2X1_LOC_816/Y 0.17fF
C55995 OR2X1_LOC_7/A OR2X1_LOC_504/a_36_216# 0.02fF
C55996 AND2X1_LOC_56/B OR2X1_LOC_140/B 0.00fF
C55997 AND2X1_LOC_473/Y OR2X1_LOC_39/A 0.05fF
C55998 OR2X1_LOC_18/Y AND2X1_LOC_244/A 0.03fF
C55999 OR2X1_LOC_329/B AND2X1_LOC_326/B 0.03fF
C56000 OR2X1_LOC_48/B OR2X1_LOC_16/A 0.11fF
C56001 OR2X1_LOC_794/a_8_216# OR2X1_LOC_301/a_8_216# 0.47fF
C56002 OR2X1_LOC_156/a_8_216# OR2X1_LOC_87/A 0.01fF
C56003 AND2X1_LOC_387/a_8_24# AND2X1_LOC_41/A 0.01fF
C56004 VDD OR2X1_LOC_658/a_8_216# 0.00fF
C56005 AND2X1_LOC_367/A OR2X1_LOC_600/A 0.05fF
C56006 AND2X1_LOC_486/Y OR2X1_LOC_158/A 0.03fF
C56007 AND2X1_LOC_803/B OR2X1_LOC_524/Y 0.38fF
C56008 AND2X1_LOC_714/a_36_24# OR2X1_LOC_48/B 0.00fF
C56009 VDD OR2X1_LOC_78/Y 0.59fF
C56010 AND2X1_LOC_436/Y AND2X1_LOC_468/a_36_24# 0.00fF
C56011 AND2X1_LOC_364/Y AND2X1_LOC_337/a_8_24# 0.01fF
C56012 OR2X1_LOC_816/A OR2X1_LOC_39/A 0.69fF
C56013 OR2X1_LOC_18/Y OR2X1_LOC_16/A 0.12fF
C56014 AND2X1_LOC_811/B AND2X1_LOC_469/a_8_24# 0.20fF
C56015 AND2X1_LOC_95/Y OR2X1_LOC_435/A 0.00fF
C56016 OR2X1_LOC_134/Y AND2X1_LOC_361/A 0.04fF
C56017 OR2X1_LOC_154/A AND2X1_LOC_22/Y 0.25fF
C56018 OR2X1_LOC_494/A OR2X1_LOC_44/Y 0.03fF
C56019 OR2X1_LOC_696/A OR2X1_LOC_696/a_8_216# 0.07fF
C56020 OR2X1_LOC_715/B OR2X1_LOC_61/Y 0.23fF
C56021 OR2X1_LOC_502/A OR2X1_LOC_356/a_8_216# 0.01fF
C56022 AND2X1_LOC_505/a_8_24# OR2X1_LOC_502/A 0.01fF
C56023 OR2X1_LOC_177/Y AND2X1_LOC_550/A 0.04fF
C56024 OR2X1_LOC_127/Y OR2X1_LOC_12/Y 0.14fF
C56025 AND2X1_LOC_94/Y INPUT_0 0.53fF
C56026 OR2X1_LOC_92/Y AND2X1_LOC_860/A 0.03fF
C56027 OR2X1_LOC_319/B OR2X1_LOC_66/A 0.17fF
C56028 OR2X1_LOC_768/A OR2X1_LOC_137/a_8_216# 0.47fF
C56029 AND2X1_LOC_555/Y OR2X1_LOC_89/A 0.10fF
C56030 OR2X1_LOC_526/Y OR2X1_LOC_144/Y 0.01fF
C56031 OR2X1_LOC_624/A OR2X1_LOC_549/A 0.10fF
C56032 VDD AND2X1_LOC_424/a_8_24# -0.00fF
C56033 OR2X1_LOC_723/a_8_216# OR2X1_LOC_737/A 0.03fF
C56034 AND2X1_LOC_56/B OR2X1_LOC_355/A 0.05fF
C56035 OR2X1_LOC_756/B AND2X1_LOC_92/Y 0.10fF
C56036 AND2X1_LOC_675/Y AND2X1_LOC_735/Y 0.61fF
C56037 OR2X1_LOC_841/a_36_216# OR2X1_LOC_841/A 0.03fF
C56038 AND2X1_LOC_721/Y OR2X1_LOC_251/Y 0.01fF
C56039 OR2X1_LOC_318/Y OR2X1_LOC_66/A 0.03fF
C56040 VDD OR2X1_LOC_586/Y 0.05fF
C56041 AND2X1_LOC_12/Y OR2X1_LOC_349/A 0.40fF
C56042 AND2X1_LOC_357/a_8_24# AND2X1_LOC_715/A 0.02fF
C56043 OR2X1_LOC_62/A OR2X1_LOC_71/A 0.24fF
C56044 OR2X1_LOC_137/a_36_216# OR2X1_LOC_235/B 0.00fF
C56045 AND2X1_LOC_568/B AND2X1_LOC_841/B 0.22fF
C56046 OR2X1_LOC_40/Y AND2X1_LOC_468/B 0.01fF
C56047 OR2X1_LOC_604/A AND2X1_LOC_161/a_8_24# 0.15fF
C56048 OR2X1_LOC_467/B OR2X1_LOC_470/A 0.01fF
C56049 OR2X1_LOC_329/B AND2X1_LOC_276/a_8_24# 0.03fF
C56050 AND2X1_LOC_74/a_8_24# OR2X1_LOC_741/Y 0.01fF
C56051 AND2X1_LOC_554/a_8_24# AND2X1_LOC_554/B 0.01fF
C56052 OR2X1_LOC_494/Y OR2X1_LOC_278/Y 0.03fF
C56053 AND2X1_LOC_766/a_36_24# AND2X1_LOC_3/Y 0.00fF
C56054 AND2X1_LOC_340/a_8_24# OR2X1_LOC_65/B 0.18fF
C56055 OR2X1_LOC_405/A OR2X1_LOC_468/A 0.03fF
C56056 AND2X1_LOC_501/Y AND2X1_LOC_573/A 0.27fF
C56057 AND2X1_LOC_22/Y OR2X1_LOC_856/a_8_216# 0.02fF
C56058 OR2X1_LOC_97/A OR2X1_LOC_653/a_8_216# 0.01fF
C56059 OR2X1_LOC_329/B AND2X1_LOC_840/A 0.16fF
C56060 OR2X1_LOC_674/a_8_216# OR2X1_LOC_495/Y 0.01fF
C56061 OR2X1_LOC_47/Y OR2X1_LOC_437/A 0.41fF
C56062 AND2X1_LOC_848/A AND2X1_LOC_793/B 0.03fF
C56063 OR2X1_LOC_326/a_8_216# OR2X1_LOC_620/Y 0.02fF
C56064 OR2X1_LOC_385/Y OR2X1_LOC_16/A 0.05fF
C56065 OR2X1_LOC_849/A OR2X1_LOC_113/B 0.01fF
C56066 OR2X1_LOC_158/A OR2X1_LOC_248/Y 0.01fF
C56067 OR2X1_LOC_426/B OR2X1_LOC_595/a_8_216# 0.32fF
C56068 OR2X1_LOC_805/A OR2X1_LOC_66/A 0.10fF
C56069 AND2X1_LOC_570/Y AND2X1_LOC_573/A 0.02fF
C56070 OR2X1_LOC_51/Y AND2X1_LOC_453/Y 0.29fF
C56071 OR2X1_LOC_49/A OR2X1_LOC_647/A 0.00fF
C56072 OR2X1_LOC_778/Y OR2X1_LOC_596/A 0.05fF
C56073 AND2X1_LOC_41/a_8_24# OR2X1_LOC_87/A 0.01fF
C56074 OR2X1_LOC_482/Y OR2X1_LOC_491/Y 0.15fF
C56075 OR2X1_LOC_8/Y AND2X1_LOC_9/a_36_24# 0.00fF
C56076 OR2X1_LOC_856/B AND2X1_LOC_311/a_36_24# 0.00fF
C56077 OR2X1_LOC_375/A OR2X1_LOC_190/Y 0.02fF
C56078 OR2X1_LOC_240/B OR2X1_LOC_78/B 0.05fF
C56079 OR2X1_LOC_739/A OR2X1_LOC_78/A 0.03fF
C56080 OR2X1_LOC_660/B AND2X1_LOC_92/Y 0.01fF
C56081 OR2X1_LOC_6/B AND2X1_LOC_838/a_8_24# 0.00fF
C56082 AND2X1_LOC_40/Y OR2X1_LOC_502/A 0.16fF
C56083 AND2X1_LOC_212/A AND2X1_LOC_211/B 0.00fF
C56084 OR2X1_LOC_235/B OR2X1_LOC_291/a_36_216# 0.00fF
C56085 OR2X1_LOC_78/B OR2X1_LOC_161/A 0.11fF
C56086 AND2X1_LOC_95/Y AND2X1_LOC_96/a_8_24# 0.11fF
C56087 OR2X1_LOC_836/A OR2X1_LOC_66/A 0.00fF
C56088 AND2X1_LOC_553/A AND2X1_LOC_113/a_8_24# 0.01fF
C56089 AND2X1_LOC_56/B OR2X1_LOC_370/a_8_216# 0.07fF
C56090 OR2X1_LOC_744/A AND2X1_LOC_653/B 0.02fF
C56091 AND2X1_LOC_729/Y OR2X1_LOC_59/Y 0.03fF
C56092 OR2X1_LOC_329/B OR2X1_LOC_237/a_8_216# 0.03fF
C56093 OR2X1_LOC_67/a_8_216# OR2X1_LOC_56/A 0.03fF
C56094 OR2X1_LOC_207/B OR2X1_LOC_193/A 0.02fF
C56095 OR2X1_LOC_685/a_8_216# OR2X1_LOC_687/A 0.40fF
C56096 AND2X1_LOC_367/A OR2X1_LOC_619/Y 0.02fF
C56097 AND2X1_LOC_61/a_36_24# OR2X1_LOC_85/A 0.00fF
C56098 OR2X1_LOC_599/Y OR2X1_LOC_13/B 0.08fF
C56099 OR2X1_LOC_696/A AND2X1_LOC_831/Y 0.41fF
C56100 VDD OR2X1_LOC_748/A 0.00fF
C56101 AND2X1_LOC_19/Y OR2X1_LOC_130/A 0.04fF
C56102 OR2X1_LOC_45/B AND2X1_LOC_307/Y 0.01fF
C56103 AND2X1_LOC_364/Y AND2X1_LOC_365/A 0.04fF
C56104 AND2X1_LOC_208/a_8_24# OR2X1_LOC_18/Y 0.01fF
C56105 OR2X1_LOC_648/A OR2X1_LOC_358/B 0.01fF
C56106 OR2X1_LOC_6/B OR2X1_LOC_827/Y 0.02fF
C56107 OR2X1_LOC_96/Y OR2X1_LOC_93/a_36_216# 0.00fF
C56108 AND2X1_LOC_21/a_8_24# INPUT_7 0.01fF
C56109 AND2X1_LOC_346/a_8_24# OR2X1_LOC_258/Y 0.01fF
C56110 AND2X1_LOC_191/B AND2X1_LOC_859/Y 0.39fF
C56111 OR2X1_LOC_185/A OR2X1_LOC_798/Y 0.03fF
C56112 OR2X1_LOC_51/Y OR2X1_LOC_26/Y 7.64fF
C56113 OR2X1_LOC_527/a_8_216# OR2X1_LOC_371/Y 0.01fF
C56114 AND2X1_LOC_735/Y OR2X1_LOC_189/A 0.00fF
C56115 OR2X1_LOC_686/B AND2X1_LOC_3/Y 0.12fF
C56116 OR2X1_LOC_663/a_36_216# AND2X1_LOC_51/Y 0.00fF
C56117 AND2X1_LOC_679/a_36_24# OR2X1_LOC_446/B 0.00fF
C56118 OR2X1_LOC_64/Y AND2X1_LOC_212/Y 0.07fF
C56119 AND2X1_LOC_547/Y AND2X1_LOC_191/Y 0.03fF
C56120 AND2X1_LOC_565/B OR2X1_LOC_189/Y 0.26fF
C56121 OR2X1_LOC_804/A OR2X1_LOC_723/B 0.07fF
C56122 OR2X1_LOC_13/B OR2X1_LOC_331/a_8_216# 0.03fF
C56123 OR2X1_LOC_815/a_36_216# OR2X1_LOC_89/A 0.00fF
C56124 AND2X1_LOC_784/A OR2X1_LOC_59/Y 0.07fF
C56125 OR2X1_LOC_161/A OR2X1_LOC_721/Y 0.07fF
C56126 OR2X1_LOC_687/Y OR2X1_LOC_678/Y 0.03fF
C56127 OR2X1_LOC_151/A OR2X1_LOC_486/a_8_216# 0.02fF
C56128 AND2X1_LOC_59/Y OR2X1_LOC_274/Y 0.01fF
C56129 OR2X1_LOC_155/A OR2X1_LOC_702/a_8_216# 0.06fF
C56130 OR2X1_LOC_78/A OR2X1_LOC_269/B 11.08fF
C56131 OR2X1_LOC_56/A AND2X1_LOC_458/a_8_24# 0.05fF
C56132 OR2X1_LOC_691/B OR2X1_LOC_19/B 0.02fF
C56133 OR2X1_LOC_490/Y OR2X1_LOC_600/A 0.03fF
C56134 OR2X1_LOC_600/A OR2X1_LOC_74/A 0.19fF
C56135 OR2X1_LOC_811/a_8_216# OR2X1_LOC_805/a_8_216# 0.47fF
C56136 OR2X1_LOC_448/a_8_216# OR2X1_LOC_161/A 0.04fF
C56137 AND2X1_LOC_390/a_8_24# OR2X1_LOC_70/Y 0.01fF
C56138 AND2X1_LOC_547/Y AND2X1_LOC_711/Y 0.09fF
C56139 OR2X1_LOC_334/B AND2X1_LOC_291/a_36_24# 0.00fF
C56140 OR2X1_LOC_640/A AND2X1_LOC_824/B 0.01fF
C56141 AND2X1_LOC_364/Y OR2X1_LOC_43/A 1.50fF
C56142 AND2X1_LOC_349/B OR2X1_LOC_51/Y 0.01fF
C56143 OR2X1_LOC_51/Y OR2X1_LOC_89/A 0.30fF
C56144 OR2X1_LOC_728/B OR2X1_LOC_730/B 0.01fF
C56145 OR2X1_LOC_516/a_8_216# OR2X1_LOC_516/B 0.01fF
C56146 AND2X1_LOC_217/Y AND2X1_LOC_141/B 0.01fF
C56147 INPUT_4 D_INPUT_5 1.01fF
C56148 AND2X1_LOC_547/Y OR2X1_LOC_70/Y 0.04fF
C56149 OR2X1_LOC_61/Y OR2X1_LOC_215/Y 0.03fF
C56150 AND2X1_LOC_456/B OR2X1_LOC_283/a_36_216# 0.00fF
C56151 OR2X1_LOC_811/a_8_216# OR2X1_LOC_362/B 0.00fF
C56152 OR2X1_LOC_723/B OR2X1_LOC_723/A 0.08fF
C56153 OR2X1_LOC_457/a_8_216# OR2X1_LOC_464/A 0.01fF
C56154 AND2X1_LOC_352/a_8_24# OR2X1_LOC_64/Y 0.01fF
C56155 OR2X1_LOC_176/Y OR2X1_LOC_417/A 0.07fF
C56156 D_INPUT_0 OR2X1_LOC_34/a_8_216# 0.06fF
C56157 OR2X1_LOC_365/a_8_216# OR2X1_LOC_367/B 0.09fF
C56158 OR2X1_LOC_61/Y AND2X1_LOC_230/a_36_24# 0.00fF
C56159 AND2X1_LOC_40/Y OR2X1_LOC_213/A 0.15fF
C56160 AND2X1_LOC_98/Y OR2X1_LOC_248/Y 0.04fF
C56161 OR2X1_LOC_458/B OR2X1_LOC_269/B 0.03fF
C56162 VDD OR2X1_LOC_304/Y 0.04fF
C56163 OR2X1_LOC_494/a_36_216# AND2X1_LOC_348/Y 0.00fF
C56164 OR2X1_LOC_493/Y OR2X1_LOC_776/A 0.15fF
C56165 AND2X1_LOC_702/Y AND2X1_LOC_863/a_8_24# 0.01fF
C56166 AND2X1_LOC_565/B OR2X1_LOC_527/Y 0.01fF
C56167 OR2X1_LOC_600/A OR2X1_LOC_261/A 0.18fF
C56168 OR2X1_LOC_470/a_8_216# OR2X1_LOC_477/Y 0.01fF
C56169 AND2X1_LOC_70/Y OR2X1_LOC_605/a_8_216# 0.18fF
C56170 OR2X1_LOC_548/A INPUT_1 0.07fF
C56171 AND2X1_LOC_530/a_8_24# D_INPUT_0 0.01fF
C56172 AND2X1_LOC_161/a_8_24# AND2X1_LOC_467/a_8_24# 0.23fF
C56173 AND2X1_LOC_566/Y OR2X1_LOC_91/A 0.33fF
C56174 OR2X1_LOC_45/B OR2X1_LOC_238/a_36_216# 0.03fF
C56175 OR2X1_LOC_660/a_8_216# OR2X1_LOC_87/A 0.01fF
C56176 OR2X1_LOC_40/Y OR2X1_LOC_278/A 0.07fF
C56177 AND2X1_LOC_392/A OR2X1_LOC_417/Y 0.03fF
C56178 OR2X1_LOC_494/a_36_216# OR2X1_LOC_753/A 0.00fF
C56179 OR2X1_LOC_574/A AND2X1_LOC_41/A 0.05fF
C56180 AND2X1_LOC_47/Y OR2X1_LOC_633/A 0.54fF
C56181 OR2X1_LOC_756/B OR2X1_LOC_563/B 0.02fF
C56182 OR2X1_LOC_438/Y OR2X1_LOC_52/B 0.02fF
C56183 OR2X1_LOC_240/B OR2X1_LOC_375/A 0.02fF
C56184 OR2X1_LOC_274/Y AND2X1_LOC_495/a_8_24# 0.01fF
C56185 OR2X1_LOC_448/B OR2X1_LOC_269/B 0.02fF
C56186 OR2X1_LOC_790/B OR2X1_LOC_375/A 0.21fF
C56187 OR2X1_LOC_598/Y AND2X1_LOC_48/A 0.17fF
C56188 OR2X1_LOC_417/A AND2X1_LOC_212/Y 0.01fF
C56189 AND2X1_LOC_719/a_8_24# AND2X1_LOC_861/B 0.01fF
C56190 OR2X1_LOC_485/Y AND2X1_LOC_727/A 0.00fF
C56191 D_INPUT_5 AND2X1_LOC_51/A 0.19fF
C56192 AND2X1_LOC_738/Y AND2X1_LOC_740/a_8_24# 0.19fF
C56193 OR2X1_LOC_188/Y OR2X1_LOC_270/Y 0.00fF
C56194 OR2X1_LOC_375/A OR2X1_LOC_161/A 0.15fF
C56195 AND2X1_LOC_59/Y OR2X1_LOC_640/a_8_216# 0.01fF
C56196 AND2X1_LOC_807/Y OR2X1_LOC_39/A 0.19fF
C56197 AND2X1_LOC_543/a_8_24# OR2X1_LOC_74/A 0.02fF
C56198 OR2X1_LOC_427/A OR2X1_LOC_44/Y 1.12fF
C56199 OR2X1_LOC_405/a_8_216# OR2X1_LOC_358/B 0.01fF
C56200 OR2X1_LOC_673/a_8_216# AND2X1_LOC_47/Y 0.00fF
C56201 OR2X1_LOC_791/B AND2X1_LOC_282/a_8_24# 0.01fF
C56202 VDD OR2X1_LOC_628/Y 0.04fF
C56203 AND2X1_LOC_51/Y OR2X1_LOC_78/B 0.31fF
C56204 OR2X1_LOC_160/A OR2X1_LOC_462/B 0.03fF
C56205 AND2X1_LOC_714/B OR2X1_LOC_31/Y 0.09fF
C56206 OR2X1_LOC_154/A AND2X1_LOC_153/a_8_24# 0.01fF
C56207 OR2X1_LOC_405/A OR2X1_LOC_449/B 0.07fF
C56208 AND2X1_LOC_537/Y OR2X1_LOC_56/A 0.10fF
C56209 OR2X1_LOC_450/a_36_216# AND2X1_LOC_425/Y 0.00fF
C56210 OR2X1_LOC_450/A OR2X1_LOC_707/B 0.48fF
C56211 OR2X1_LOC_413/a_8_216# OR2X1_LOC_690/A 0.02fF
C56212 OR2X1_LOC_653/A OR2X1_LOC_130/A 0.01fF
C56213 OR2X1_LOC_276/a_8_216# OR2X1_LOC_549/A 0.05fF
C56214 OR2X1_LOC_844/Y OR2X1_LOC_624/Y 0.33fF
C56215 OR2X1_LOC_339/a_36_216# OR2X1_LOC_814/A 0.01fF
C56216 AND2X1_LOC_472/B AND2X1_LOC_233/a_8_24# 0.01fF
C56217 AND2X1_LOC_621/Y OR2X1_LOC_52/B 0.05fF
C56218 AND2X1_LOC_389/a_8_24# OR2X1_LOC_586/Y 0.01fF
C56219 OR2X1_LOC_158/A AND2X1_LOC_660/A 0.07fF
C56220 AND2X1_LOC_342/Y AND2X1_LOC_359/B 0.00fF
C56221 OR2X1_LOC_525/Y OR2X1_LOC_680/Y 0.15fF
C56222 OR2X1_LOC_482/Y OR2X1_LOC_674/Y 0.01fF
C56223 AND2X1_LOC_271/a_8_24# OR2X1_LOC_344/A 0.01fF
C56224 OR2X1_LOC_768/A OR2X1_LOC_814/A 0.11fF
C56225 OR2X1_LOC_744/A AND2X1_LOC_477/A 0.03fF
C56226 OR2X1_LOC_680/A OR2X1_LOC_26/Y 10.36fF
C56227 OR2X1_LOC_604/A OR2X1_LOC_55/a_8_216# 0.06fF
C56228 AND2X1_LOC_51/Y OR2X1_LOC_721/Y 0.01fF
C56229 AND2X1_LOC_146/a_8_24# OR2X1_LOC_78/A 0.01fF
C56230 OR2X1_LOC_173/Y OR2X1_LOC_265/Y 0.05fF
C56231 OR2X1_LOC_246/a_8_216# OR2X1_LOC_85/A 0.01fF
C56232 AND2X1_LOC_250/a_8_24# OR2X1_LOC_362/A 0.01fF
C56233 OR2X1_LOC_442/a_8_216# AND2X1_LOC_469/B 0.01fF
C56234 OR2X1_LOC_46/A OR2X1_LOC_394/a_8_216# 0.11fF
C56235 OR2X1_LOC_290/a_36_216# OR2X1_LOC_416/Y 0.00fF
C56236 OR2X1_LOC_155/A OR2X1_LOC_798/a_8_216# 0.02fF
C56237 AND2X1_LOC_728/Y AND2X1_LOC_147/Y 0.83fF
C56238 OR2X1_LOC_743/A OR2X1_LOC_595/a_8_216# 0.01fF
C56239 OR2X1_LOC_719/B VSS 0.17fF
C56240 OR2X1_LOC_779/A VSS 0.02fF
C56241 OR2X1_LOC_174/Y VSS 0.10fF
C56242 OR2X1_LOC_121/A VSS 0.27fF
C56243 OR2X1_LOC_142/Y VSS 0.19fF
C56244 OR2X1_LOC_198/A VSS 0.46fF
C56245 AND2X1_LOC_52/Y VSS 0.26fF
C56246 OR2X1_LOC_390/A VSS -0.53fF
C56247 AND2X1_LOC_582/B VSS 0.08fF
C56248 OR2X1_LOC_589/Y VSS 0.16fF
C56249 OR2X1_LOC_423/Y VSS 0.39fF
C56250 AND2X1_LOC_570/a_8_24# VSS 0.10fF
C56251 AND2X1_LOC_563/Y VSS 0.05fF
C56252 AND2X1_LOC_562/Y VSS 0.70fF
C56253 OR2X1_LOC_365/B VSS 0.59fF
C56254 OR2X1_LOC_323/Y VSS 0.43fF
C56255 OR2X1_LOC_338/A VSS -0.39fF
C56256 OR2X1_LOC_334/A VSS 0.22fF
C56257 D_GATE_366 VSS 0.02fF
C56258 OR2X1_LOC_366/Y VSS 0.41fF
C56259 OR2X1_LOC_539/B VSS 0.66fF
C56260 OR2X1_LOC_560/A VSS -0.12fF
C56261 OR2X1_LOC_549/A VSS 0.61fF
C56262 OR2X1_LOC_548/B VSS 0.11fF
C56263 AND2X1_LOC_763/B VSS 0.19fF
C56264 INPUT_6 VSS 0.26fF
C56265 AND2X1_LOC_742/A VSS 0.16fF
C56266 AND2X1_LOC_738/Y VSS 0.10fF
C56267 OR2X1_LOC_789/A VSS 0.14fF
C56268 OR2X1_LOC_750/Y VSS -0.81fF
C56269 AND2X1_LOC_778/Y VSS 0.21fF
C56270 AND2X1_LOC_786/Y VSS -3.08fF
C56271 AND2X1_LOC_785/Y VSS 0.16fF
C56272 AND2X1_LOC_772/Y VSS 0.29fF
C56273 OR2X1_LOC_767/Y VSS 0.06fF
C56274 OR2X1_LOC_515/Y VSS 0.56fF
C56275 AND2X1_LOC_228/a_8_24# VSS 0.10fF
C56276 AND2X1_LOC_202/Y VSS 0.15fF
C56277 AND2X1_LOC_201/Y VSS 0.13fF
C56278 AND2X1_LOC_657/A VSS 0.26fF
C56279 OR2X1_LOC_730/A VSS 0.18fF
C56280 OR2X1_LOC_722/B VSS 0.28fF
C56281 OR2X1_LOC_605/Y VSS 0.27fF
C56282 OR2X1_LOC_712/B VSS 0.28fF
C56283 OR2X1_LOC_460/A VSS 0.15fF
C56284 AND2X1_LOC_48/Y VSS 0.03fF
C56285 OR2X1_LOC_130/Y VSS 0.07fF
C56286 OR2X1_LOC_217/A VSS 0.36fF
C56287 OR2X1_LOC_140/Y VSS 0.10fF
C56288 OR2X1_LOC_152/A VSS -0.04fF
C56289 OR2X1_LOC_163/Y VSS 0.35fF
C56290 OR2X1_LOC_163/A VSS 0.15fF
C56291 OR2X1_LOC_356/A VSS 0.20fF
C56292 OR2X1_LOC_355/A VSS 0.13fF
C56293 OR2X1_LOC_390/B VSS 0.43fF
C56294 OR2X1_LOC_180/B VSS 0.36fF
C56295 OR2X1_LOC_399/Y VSS -0.33fF
C56296 GATE_579 VSS 0.09fF
C56297 OR2X1_LOC_593/B VSS 0.42fF
C56298 OR2X1_LOC_590/Y VSS 0.04fF
C56299 OR2X1_LOC_378/A VSS 0.02fF
C56300 OR2X1_LOC_322/Y VSS 0.33fF
C56301 OR2X1_LOC_338/B VSS 0.11fF
C56302 OR2X1_LOC_333/A VSS -0.11fF
C56303 OR2X1_LOC_300/Y VSS 0.27fF
C56304 OR2X1_LOC_348/B VSS -0.27fF
C56305 OR2X1_LOC_550/A VSS 0.18fF
C56306 OR2X1_LOC_577/B VSS 0.16fF
C56307 OR2X1_LOC_561/A VSS 0.18fF
C56308 OR2X1_LOC_558/A VSS 0.12fF
C56309 AND2X1_LOC_796/A VSS 0.65fF
C56310 AND2X1_LOC_779/Y VSS 0.10fF
C56311 OR2X1_LOC_801/B VSS 0.33fF
C56312 OR2X1_LOC_644/A VSS 0.29fF
C56313 AND2X1_LOC_804/A VSS 0.26fF
C56314 AND2X1_LOC_750/a_8_24# VSS 0.10fF
C56315 OR2X1_LOC_749/Y VSS 0.23fF
C56316 OR2X1_LOC_515/A VSS 0.18fF
C56317 OR2X1_LOC_138/A VSS 0.37fF
C56318 AND2X1_LOC_215/A VSS 0.21fF
C56319 AND2X1_LOC_204/Y VSS 0.32fF
C56320 AND2X1_LOC_203/Y VSS 0.10fF
C56321 OR2X1_LOC_595/A VSS -1.29fF
C56322 OR2X1_LOC_776/A VSS 0.23fF
C56323 OR2X1_LOC_730/B VSS 0.11fF
C56324 OR2X1_LOC_728/A VSS 0.13fF
C56325 OR2X1_LOC_723/A VSS 0.18fF
C56326 OR2X1_LOC_374/Y VSS 0.20fF
C56327 OR2X1_LOC_493/Y VSS 0.73fF
C56328 OR2X1_LOC_713/A VSS -0.72fF
C56329 AND2X1_LOC_409/B VSS 0.28fF
C56330 D_INPUT_6 VSS 0.19fF
C56331 AND2X1_LOC_419/a_8_24# VSS 0.10fF
C56332 OR2X1_LOC_199/B VSS 0.10fF
C56333 AND2X1_LOC_41/Y VSS 0.36fF
C56334 OR2X1_LOC_160/Y VSS 0.26fF
C56335 OR2X1_LOC_356/B VSS 0.36fF
C56336 OR2X1_LOC_319/Y VSS 0.28fF
C56337 OR2X1_LOC_339/A VSS 0.07fF
C56338 OR2X1_LOC_112/A VSS 0.21fF
C56339 OR2X1_LOC_367/B VSS 0.81fF
C56340 OR2X1_LOC_364/Y VSS 0.02fF
C56341 OR2X1_LOC_398/Y VSS 0.29fF
C56342 OR2X1_LOC_598/A VSS -4.30fF
C56343 OR2X1_LOC_349/A VSS 0.26fF
C56344 OR2X1_LOC_843/B VSS 0.24fF
C56345 OR2X1_LOC_376/Y VSS 0.10fF
C56346 OR2X1_LOC_788/B VSS 0.40fF
C56347 OR2X1_LOC_578/B VSS 0.39fF
C56348 OR2X1_LOC_566/Y VSS 0.11fF
C56349 OR2X1_LOC_502/Y VSS 0.22fF
C56350 OR2X1_LOC_580/A VSS -0.80fF
C56351 OR2X1_LOC_561/B VSS -0.63fF
C56352 AND2X1_LOC_797/B VSS 0.19fF
C56353 AND2X1_LOC_781/Y VSS 0.18fF
C56354 OR2X1_LOC_747/Y VSS 0.06fF
C56355 AND2X1_LOC_774/A VSS -1.63fF
C56356 AND2X1_LOC_769/Y VSS 0.10fF
C56357 AND2X1_LOC_793/a_8_24# VSS 0.10fF
C56358 AND2X1_LOC_789/Y VSS -2.29fF
C56359 OR2X1_LOC_550/B VSS 0.40fF
C56360 OR2X1_LOC_513/Y VSS 0.25fF
C56361 OR2X1_LOC_779/B VSS 0.51fF
C56362 OR2X1_LOC_512/Y VSS 0.18fF
C56363 OR2X1_LOC_257/Y VSS 0.06fF
C56364 OR2X1_LOC_342/A VSS 0.20fF
C56365 AND2X1_LOC_206/Y VSS 0.18fF
C56366 OR2X1_LOC_241/B VSS 0.46fF
C56367 OR2X1_LOC_227/A VSS 0.13fF
C56368 OR2X1_LOC_723/B VSS 0.35fF
C56369 OR2X1_LOC_303/B VSS 0.28fF
C56370 OR2X1_LOC_740/B VSS 0.17fF
C56371 OR2X1_LOC_731/A VSS 0.36fF
C56372 OR2X1_LOC_308/Y VSS 1.05fF
C56373 OR2X1_LOC_469/B VSS 0.18fF
C56374 OR2X1_LOC_546/A VSS 0.02fF
C56375 AND2X1_LOC_430/B VSS -0.26fF
C56376 OR2X1_LOC_446/A VSS 0.15fF
C56377 OR2X1_LOC_20/A VSS 0.18fF
C56378 OR2X1_LOC_183/Y VSS 0.16fF
C56379 OR2X1_LOC_437/A VSS -8.26fF
C56380 OR2X1_LOC_71/A VSS 0.34fF
C56381 OR2X1_LOC_172/Y VSS -0.20fF
C56382 AND2X1_LOC_39/Y VSS 0.15fF
C56383 OR2X1_LOC_162/A VSS 0.18fF
C56384 OR2X1_LOC_357/A VSS 0.01fF
C56385 OR2X1_LOC_397/Y VSS 0.07fF
C56386 OR2X1_LOC_349/B VSS 0.08fF
C56387 OR2X1_LOC_331/Y VSS 0.34fF
C56388 OR2X1_LOC_375/Y VSS 0.07fF
C56389 OR2X1_LOC_387/A VSS 0.17fF
C56390 OR2X1_LOC_746/Y VSS 0.18fF
C56391 OR2X1_LOC_745/Y VSS -0.14fF
C56392 AND2X1_LOC_771/B VSS 0.19fF
C56393 AND2X1_LOC_770/a_8_24# VSS 0.10fF
C56394 AND2X1_LOC_792/a_8_24# VSS 0.10fF
C56395 OR2X1_LOC_759/Y VSS 0.10fF
C56396 OR2X1_LOC_568/A VSS -0.26fF
C56397 OR2X1_LOC_854/A VSS 0.38fF
C56398 OR2X1_LOC_551/A VSS 0.18fF
C56399 OR2X1_LOC_580/B VSS -2.43fF
C56400 OR2X1_LOC_577/Y VSS 0.25fF
C56401 OR2X1_LOC_562/A VSS 0.30fF
C56402 OR2X1_LOC_523/A VSS 0.13fF
C56403 OR2X1_LOC_735/B VSS -0.05fF
C56404 OR2X1_LOC_534/Y VSS 0.18fF
C56405 AND2X1_LOC_219/A VSS 0.22fF
C56406 AND2X1_LOC_208/Y VSS 0.10fF
C56407 OR2X1_LOC_268/Y VSS -0.13fF
C56408 OR2X1_LOC_80/A VSS -3.61fF
C56409 OR2X1_LOC_68/B VSS 0.66fF
C56410 AND2X1_LOC_225/a_8_24# VSS 0.10fF
C56411 D_INPUT_1 VSS 0.74fF
C56412 OR2X1_LOC_259/A VSS 0.04fF
C56413 OR2X1_LOC_248/A VSS 0.15fF
C56414 OR2X1_LOC_13/B VSS -5.53fF
C56415 OR2X1_LOC_72/Y VSS 0.31fF
C56416 OR2X1_LOC_741/A VSS 0.18fF
C56417 OR2X1_LOC_733/Y VSS 0.17fF
C56418 OR2X1_LOC_428/A VSS 1.83fF
C56419 OR2X1_LOC_748/Y VSS 0.06fF
C56420 OR2X1_LOC_731/B VSS 0.17fF
C56421 OR2X1_LOC_209/A VSS 0.17fF
C56422 OR2X1_LOC_714/A VSS 0.18fF
C56423 OR2X1_LOC_317/B VSS 0.02fF
C56424 OR2X1_LOC_446/B VSS 0.49fF
C56425 OR2X1_LOC_724/A VSS 0.40fF
C56426 OR2X1_LOC_451/B VSS 0.50fF
C56427 AND2X1_LOC_406/a_8_24# VSS 0.10fF
C56428 OR2X1_LOC_608/Y VSS 0.10fF
C56429 OR2X1_LOC_171/Y VSS 0.11fF
C56430 OR2X1_LOC_212/B VSS 0.36fF
C56431 OR2X1_LOC_181/Y VSS 0.10fF
C56432 OR2X1_LOC_357/B VSS 0.11fF
C56433 OR2X1_LOC_544/B VSS 0.51fF
C56434 OR2X1_LOC_228/Y VSS 0.57fF
C56435 OR2X1_LOC_641/B VSS 0.31fF
C56436 OR2X1_LOC_396/Y VSS 0.24fF
C56437 OR2X1_LOC_366/A VSS 0.18fF
C56438 OR2X1_LOC_170/Y VSS 0.30fF
C56439 OR2X1_LOC_570/Y VSS 0.19fF
C56440 OR2X1_LOC_562/B VSS 0.17fF
C56441 AND2X1_LOC_783/B VSS 0.05fF
C56442 OR2X1_LOC_743/Y VSS -0.07fF
C56443 AND2X1_LOC_792/B VSS 0.10fF
C56444 OR2X1_LOC_551/B VSS 0.37fF
C56445 OR2X1_LOC_522/Y VSS 0.08fF
C56446 OR2X1_LOC_501/A VSS 0.18fF
C56447 OR2X1_LOC_844/B VSS 0.43fF
C56448 OR2X1_LOC_533/A VSS -0.05fF
C56449 AND2X1_LOC_220/B VSS -0.20fF
C56450 AND2X1_LOC_209/Y VSS 0.08fF
C56451 OR2X1_LOC_342/B VSS -0.07fF
C56452 OR2X1_LOC_777/B VSS -0.62fF
C56453 OR2X1_LOC_259/B VSS 0.31fF
C56454 OR2X1_LOC_284/B VSS 0.25fF
C56455 OR2X1_LOC_161/B VSS 1.07fF
C56456 AND2X1_LOC_44/Y VSS 0.85fF
C56457 OR2X1_LOC_269/A VSS 0.38fF
C56458 AND2X1_LOC_202/a_8_24# VSS 0.10fF
C56459 OR2X1_LOC_67/Y VSS 0.31fF
C56460 OR2X1_LOC_227/B VSS 0.17fF
C56461 OR2X1_LOC_771/B VSS 0.59fF
C56462 OR2X1_LOC_675/Y VSS -1.69fF
C56463 OR2X1_LOC_703/Y VSS 0.44fF
C56464 OR2X1_LOC_732/A VSS 0.21fF
C56465 OR2X1_LOC_424/Y VSS -0.02fF
C56466 OR2X1_LOC_406/A VSS -0.19fF
C56467 AND2X1_LOC_405/a_8_24# VSS 0.10fF
C56468 AND2X1_LOC_438/a_8_24# VSS 0.10fF
C56469 OR2X1_LOC_415/Y VSS 0.26fF
C56470 OR2X1_LOC_622/B VSS 0.16fF
C56471 AND2X1_LOC_36/Y VSS -4.77fF
C56472 OR2X1_LOC_168/Y VSS 0.24fF
C56473 OR2X1_LOC_181/A VSS 0.15fF
C56474 OR2X1_LOC_192/B VSS 0.22fF
C56475 OR2X1_LOC_373/Y VSS 0.19fF
C56476 OR2X1_LOC_395/Y VSS 0.24fF
C56477 OR2X1_LOC_384/Y VSS 0.25fF
C56478 OR2X1_LOC_358/A VSS -0.48fF
C56479 OR2X1_LOC_339/Y VSS 0.14fF
C56480 AND2X1_LOC_88/Y VSS 0.32fF
C56481 OR2X1_LOC_227/Y VSS 0.37fF
C56482 OR2X1_LOC_366/B VSS 0.32fF
C56483 OR2X1_LOC_532/Y VSS -0.29fF
C56484 OR2X1_LOC_552/A VSS 0.15fF
C56485 OR2X1_LOC_318/B VSS 0.56fF
C56486 OR2X1_LOC_569/A VSS 0.18fF
C56487 OR2X1_LOC_549/Y VSS 0.35fF
C56488 OR2X1_LOC_563/A VSS -1.40fF
C56489 OR2X1_LOC_115/B VSS -0.21fF
C56490 OR2X1_LOC_140/B VSS -0.01fF
C56491 OR2X1_LOC_579/A VSS 0.36fF
C56492 OR2X1_LOC_571/Y VSS 0.11fF
C56493 AND2X1_LOC_793/B VSS 0.22fF
C56494 OR2X1_LOC_754/Y VSS 0.07fF
C56495 OR2X1_LOC_753/Y VSS -0.04fF
C56496 OR2X1_LOC_588/A VSS 0.17fF
C56497 INPUT_7 VSS 0.16fF
C56498 OR2X1_LOC_508/Y VSS -0.12fF
C56499 GATE_222 VSS 0.04fF
C56500 AND2X1_LOC_222/Y VSS -0.64fF
C56501 AND2X1_LOC_289/a_8_24# VSS 0.10fF
C56502 OR2X1_LOC_240/A VSS 0.41fF
C56503 AND2X1_LOC_278/a_8_24# VSS 0.10fF
C56504 AND2X1_LOC_245/a_8_24# VSS 0.10fF
C56505 OR2X1_LOC_66/A VSS -4.58fF
C56506 OR2X1_LOC_344/A VSS -0.05fF
C56507 AND2X1_LOC_361/A VSS 0.68fF
C56508 AND2X1_LOC_266/Y VSS 0.22fF
C56509 OR2X1_LOC_265/Y VSS 0.13fF
C56510 OR2X1_LOC_736/A VSS 0.22fF
C56511 OR2X1_LOC_632/Y VSS 0.48fF
C56512 OR2X1_LOC_772/A VSS 0.24fF
C56513 OR2X1_LOC_113/B VSS 0.30fF
C56514 OR2X1_LOC_757/Y VSS 0.22fF
C56515 OR2X1_LOC_732/B VSS 0.14fF
C56516 OR2X1_LOC_714/Y VSS 0.17fF
C56517 OR2X1_LOC_715/A VSS 0.15fF
C56518 OR2X1_LOC_725/A VSS 0.18fF
C56519 OR2X1_LOC_705/Y VSS 0.12fF
C56520 OR2X1_LOC_421/Y VSS 0.18fF
C56521 AND2X1_LOC_459/a_8_24# VSS 0.10fF
C56522 OR2X1_LOC_378/Y VSS 0.14fF
C56523 AND2X1_LOC_426/a_8_24# VSS 0.10fF
C56524 OR2X1_LOC_414/Y VSS 0.16fF
C56525 AND2X1_LOC_619/B VSS -0.09fF
C56526 OR2X1_LOC_627/Y VSS 0.08fF
C56527 OR2X1_LOC_626/Y VSS 0.20fF
C56528 OR2X1_LOC_646/B VSS 0.32fF
C56529 AND2X1_LOC_607/a_8_24# VSS 0.10fF
C56530 OR2X1_LOC_27/Y VSS 0.16fF
C56531 OR2X1_LOC_52/B VSS 1.59fF
C56532 OR2X1_LOC_39/A VSS 1.02fF
C56533 OR2X1_LOC_16/Y VSS 0.22fF
C56534 OR2X1_LOC_192/A VSS 0.18fF
C56535 OR2X1_LOC_190/Y VSS 0.43fF
C56536 OR2X1_LOC_182/B VSS 0.18fF
C56537 OR2X1_LOC_439/B VSS 0.02fF
C56538 OR2X1_LOC_371/Y VSS 0.51fF
C56539 OR2X1_LOC_358/B VSS 0.24fF
C56540 OR2X1_LOC_340/Y VSS 0.36fF
C56541 OR2X1_LOC_341/Y VSS 0.18fF
C56542 OR2X1_LOC_362/A VSS 0.45fF
C56543 OR2X1_LOC_269/B VSS -5.04fF
C56544 OR2X1_LOC_552/B VSS 0.17fF
C56545 OR2X1_LOC_569/B VSS 0.16fF
C56546 OR2X1_LOC_563/B VSS 0.21fF
C56547 OR2X1_LOC_579/B VSS 0.18fF
C56548 OR2X1_LOC_573/Y VSS 0.17fF
C56549 OR2X1_LOC_586/Y VSS -0.45fF
C56550 OR2X1_LOC_302/A VSS -0.05fF
C56551 OR2X1_LOC_633/A VSS 0.65fF
C56552 AND2X1_LOC_806/A VSS -0.43fF
C56553 AND2X1_LOC_287/Y VSS 0.13fF
C56554 AND2X1_LOC_286/Y VSS 0.10fF
C56555 AND2X1_LOC_207/B VSS 0.10fF
C56556 AND2X1_LOC_194/Y VSS -0.02fF
C56557 AND2X1_LOC_193/Y VSS 0.10fF
C56558 AND2X1_LOC_212/B VSS 0.13fF
C56559 AND2X1_LOC_222/a_8_24# VSS 0.10fF
C56560 AND2X1_LOC_219/Y VSS -1.06fF
C56561 AND2X1_LOC_218/Y VSS -0.06fF
C56562 AND2X1_LOC_860/A VSS 0.24fF
C56563 AND2X1_LOC_243/Y VSS -2.09fF
C56564 OR2X1_LOC_793/B VSS 0.08fF
C56565 OR2X1_LOC_737/A VSS -1.19fF
C56566 OR2X1_LOC_475/B VSS 0.46fF
C56567 OR2X1_LOC_721/Y VSS 0.66fF
C56568 OR2X1_LOC_778/B VSS 0.18fF
C56569 OR2X1_LOC_733/A VSS 0.24fF
C56570 OR2X1_LOC_44/Y VSS 0.95fF
C56571 OR2X1_LOC_725/B VSS 0.21fF
C56572 OR2X1_LOC_708/Y VSS 0.18fF
C56573 AND2X1_LOC_434/Y VSS -1.84fF
C56574 AND2X1_LOC_727/B VSS 0.16fF
C56575 AND2X1_LOC_374/Y VSS 0.26fF
C56576 OR2X1_LOC_372/Y VSS -0.02fF
C56577 AND2X1_LOC_404/B VSS 0.08fF
C56578 AND2X1_LOC_651/B VSS 0.21fF
C56579 OR2X1_LOC_630/B VSS 0.22fF
C56580 AND2X1_LOC_92/Y VSS 0.47fF
C56581 OR2X1_LOC_607/A VSS 0.15fF
C56582 OR2X1_LOC_16/A VSS -3.88fF
C56583 OR2X1_LOC_25/Y VSS 0.25fF
C56584 AND2X1_LOC_810/B VSS 0.12fF
C56585 AND2X1_LOC_802/Y VSS 0.24fF
C56586 OR2X1_LOC_393/Y VSS 0.22fF
C56587 OR2X1_LOC_363/A VSS 0.19fF
C56588 OR2X1_LOC_244/Y VSS 0.47fF
C56589 OR2X1_LOC_347/Y VSS 0.18fF
C56590 OR2X1_LOC_564/A VSS -0.01fF
C56591 OR2X1_LOC_553/A VSS -1.03fF
C56592 OR2X1_LOC_541/B VSS 0.25fF
C56593 OR2X1_LOC_575/A VSS -0.05fF
C56594 OR2X1_LOC_570/A VSS 0.18fF
C56595 OR2X1_LOC_596/A VSS 0.25fF
C56596 AND2X1_LOC_298/a_8_24# VSS 0.10fF
C56597 AND2X1_LOC_276/a_8_24# VSS 0.10fF
C56598 OR2X1_LOC_275/Y VSS 0.27fF
C56599 AND2X1_LOC_254/a_8_24# VSS 0.10fF
C56600 OR2X1_LOC_253/Y VSS 0.08fF
C56601 AND2X1_LOC_240/Y VSS 0.15fF
C56602 OR2X1_LOC_278/Y VSS 0.08fF
C56603 OR2X1_LOC_641/A VSS 0.28fF
C56604 AND2X1_LOC_265/a_8_24# VSS 0.10fF
C56605 AND2X1_LOC_213/B VSS 0.21fF
C56606 OR2X1_LOC_158/Y VSS -0.07fF
C56607 AND2X1_LOC_223/A VSS 0.21fF
C56608 AND2X1_LOC_220/Y VSS 0.14fF
C56609 OR2X1_LOC_802/A VSS 0.18fF
C56610 OR2X1_LOC_539/Y VSS -0.32fF
C56611 OR2X1_LOC_794/A VSS 0.07fF
C56612 OR2X1_LOC_755/Y VSS 0.06fF
C56613 OR2X1_LOC_59/Y VSS 1.32fF
C56614 OR2X1_LOC_784/B VSS 0.17fF
C56615 OR2X1_LOC_307/A VSS 0.39fF
C56616 OR2X1_LOC_766/Y VSS 0.08fF
C56617 OR2X1_LOC_733/B VSS 0.13fF
C56618 OR2X1_LOC_719/Y VSS 0.29fF
C56619 OR2X1_LOC_726/A VSS 0.26fF
C56620 OR2X1_LOC_744/Y VSS 0.10fF
C56621 AND2X1_LOC_454/A VSS 0.26fF
C56622 OR2X1_LOC_418/Y VSS 0.12fF
C56623 AND2X1_LOC_436/B VSS 0.26fF
C56624 OR2X1_LOC_433/Y VSS 0.17fF
C56625 OR2X1_LOC_432/Y VSS 0.35fF
C56626 AND2X1_LOC_469/B VSS 0.05fF
C56627 AND2X1_LOC_436/Y VSS -0.28fF
C56628 AND2X1_LOC_476/Y VSS -1.73fF
C56629 AND2X1_LOC_475/Y VSS 0.20fF
C56630 AND2X1_LOC_464/A VSS 0.28fF
C56631 AND2X1_LOC_457/a_8_24# VSS 0.10fF
C56632 OR2X1_LOC_368/Y VSS 0.12fF
C56633 OR2X1_LOC_461/A VSS 0.17fF
C56634 AND2X1_LOC_404/A VSS 0.06fF
C56635 AND2X1_LOC_401/Y VSS 0.15fF
C56636 OR2X1_LOC_604/Y VSS 0.02fF
C56637 OR2X1_LOC_603/Y VSS 0.06fF
C56638 AND2X1_LOC_637/Y VSS 0.08fF
C56639 OR2X1_LOC_588/Y VSS 0.24fF
C56640 AND2X1_LOC_642/Y VSS 0.13fF
C56641 AND2X1_LOC_18/Y VSS -5.89fF
C56642 AND2X1_LOC_627/a_8_24# VSS 0.10fF
C56643 AND2X1_LOC_7/B VSS -5.59fF
C56644 OR2X1_LOC_69/Y VSS 0.07fF
C56645 OR2X1_LOC_69/A VSS 0.01fF
C56646 INPUT_2 VSS 0.21fF
C56647 AND2X1_LOC_811/B VSS 0.23fF
C56648 AND2X1_LOC_804/Y VSS 0.02fF
C56649 AND2X1_LOC_820/B VSS 0.05fF
C56650 OR2X1_LOC_787/B VSS -0.15fF
C56651 OR2X1_LOC_543/A VSS 0.19fF
C56652 OR2X1_LOC_382/A VSS 0.31fF
C56653 OR2X1_LOC_12/Y VSS 0.92fF
C56654 OR2X1_LOC_474/B VSS 0.29fF
C56655 OR2X1_LOC_584/Y VSS 0.12fF
C56656 OR2X1_LOC_564/B VSS 0.40fF
C56657 OR2X1_LOC_553/B VSS 0.28fF
C56658 OR2X1_LOC_190/B VSS 0.35fF
C56659 AND2X1_LOC_212/Y VSS 0.16fF
C56660 OR2X1_LOC_230/Y VSS 0.08fF
C56661 OR2X1_LOC_229/Y VSS -0.13fF
C56662 AND2X1_LOC_264/a_8_24# VSS 0.10fF
C56663 OR2X1_LOC_347/B VSS 0.10fF
C56664 OR2X1_LOC_254/A VSS 0.15fF
C56665 AND2X1_LOC_285/Y VSS -0.83fF
C56666 AND2X1_LOC_275/a_8_24# VSS 0.10fF
C56667 AND2X1_LOC_244/A VSS 0.30fF
C56668 OR2X1_LOC_486/Y VSS 0.17fF
C56669 OR2X1_LOC_738/A VSS 0.57fF
C56670 OR2X1_LOC_765/Y VSS 0.15fF
C56671 OR2X1_LOC_720/Y VSS 0.10fF
C56672 OR2X1_LOC_711/A VSS -0.13fF
C56673 AND2X1_LOC_470/B VSS 0.08fF
C56674 AND2X1_LOC_452/Y VSS 0.14fF
C56675 AND2X1_LOC_434/a_8_24# VSS 0.10fF
C56676 AND2X1_LOC_480/A VSS 0.19fF
C56677 AND2X1_LOC_477/Y VSS 0.21fF
C56678 AND2X1_LOC_469/Y VSS 0.11fF
C56679 AND2X1_LOC_455/B VSS 0.08fF
C56680 OR2X1_LOC_213/B VSS 0.17fF
C56681 AND2X1_LOC_663/A VSS 0.56fF
C56682 AND2X1_LOC_658/Y VSS 0.12fF
C56683 AND2X1_LOC_657/Y VSS 0.91fF
C56684 OR2X1_LOC_79/Y VSS 0.11fF
C56685 AND2X1_LOC_655/A VSS -3.03fF
C56686 AND2X1_LOC_648/a_8_24# VSS 0.10fF
C56687 AND2X1_LOC_644/Y VSS 0.08fF
C56688 OR2X1_LOC_623/B VSS 0.22fF
C56689 AND2X1_LOC_637/a_8_24# VSS 0.10fF
C56690 OR2X1_LOC_585/Y VSS 0.02fF
C56691 OR2X1_LOC_629/B VSS 0.19fF
C56692 AND2X1_LOC_604/a_8_24# VSS 0.10fF
C56693 OR2X1_LOC_24/Y VSS 0.06fF
C56694 OR2X1_LOC_48/B VSS 0.90fF
C56695 OR2X1_LOC_35/Y VSS 0.24fF
C56696 OR2X1_LOC_13/Y VSS -0.27fF
C56697 OR2X1_LOC_855/A VSS 0.01fF
C56698 AND2X1_LOC_829/a_8_24# VSS 0.10fF
C56699 OR2X1_LOC_828/Y VSS 0.13fF
C56700 OR2X1_LOC_820/B VSS -0.11fF
C56701 AND2X1_LOC_818/a_8_24# VSS 0.10fF
C56702 OR2X1_LOC_6/A VSS 1.62fF
C56703 AND2X1_LOC_805/Y VSS -0.00fF
C56704 OR2X1_LOC_392/A VSS 0.19fF
C56705 OR2X1_LOC_391/A VSS -0.56fF
C56706 OR2X1_LOC_380/Y VSS 0.11fF
C56707 OR2X1_LOC_565/A VSS 0.45fF
C56708 OR2X1_LOC_576/A VSS 0.35fF
C56709 OR2X1_LOC_267/Y VSS 0.32fF
C56710 OR2X1_LOC_594/Y VSS -0.32fF
C56711 OR2X1_LOC_583/Y VSS 0.06fF
C56712 AND2X1_LOC_242/B VSS -0.51fF
C56713 OR2X1_LOC_238/Y VSS 0.09fF
C56714 OR2X1_LOC_297/A VSS 0.18fF
C56715 AND2X1_LOC_296/a_8_24# VSS 0.10fF
C56716 OR2X1_LOC_56/A VSS -7.20fF
C56717 AND2X1_LOC_285/a_8_24# VSS 0.10fF
C56718 OR2X1_LOC_281/Y VSS 0.21fF
C56719 OR2X1_LOC_266/A VSS -0.20fF
C56720 AND2X1_LOC_263/a_8_24# VSS 0.10fF
C56721 OR2X1_LOC_785/B VSS 0.08fF
C56722 D_GATE_741 VSS 0.12fF
C56723 OR2X1_LOC_741/Y VSS -0.10fF
C56724 OR2X1_LOC_816/A VSS 0.44fF
C56725 OR2X1_LOC_738/B VSS 0.17fF
C56726 OR2X1_LOC_803/A VSS 0.00fF
C56727 AND2X1_LOC_470/A VSS 0.10fF
C56728 AND2X1_LOC_454/Y VSS 0.11fF
C56729 AND2X1_LOC_453/Y VSS 0.16fF
C56730 AND2X1_LOC_471/Y VSS 0.34fF
C56731 AND2X1_LOC_500/B VSS 0.19fF
C56732 OR2X1_LOC_489/A VSS -0.15fF
C56733 OR2X1_LOC_214/A VSS 0.02fF
C56734 OR2X1_LOC_222/A VSS 0.17fF
C56735 OR2X1_LOC_215/Y VSS 0.12fF
C56736 AND2X1_LOC_443/Y VSS -0.09fF
C56737 OR2X1_LOC_442/Y VSS 0.06fF
C56738 OR2X1_LOC_461/B VSS 0.19fF
C56739 OR2X1_LOC_410/Y VSS 0.07fF
C56740 OR2X1_LOC_435/A VSS 0.21fF
C56741 AND2X1_LOC_433/a_8_24# VSS 0.10fF
C56742 AND2X1_LOC_465/A VSS 0.28fF
C56743 AND2X1_LOC_455/a_8_24# VSS 0.10fF
C56744 AND2X1_LOC_403/B VSS 0.02fF
C56745 OR2X1_LOC_394/Y VSS 0.22fF
C56746 AND2X1_LOC_639/B VSS 0.31fF
C56747 OR2X1_LOC_720/A VSS 0.15fF
C56748 OR2X1_LOC_668/Y VSS 0.07fF
C56749 OR2X1_LOC_161/A VSS 1.43fF
C56750 OR2X1_LOC_612/Y VSS -0.10fF
C56751 OR2X1_LOC_631/A VSS 0.19fF
C56752 OR2X1_LOC_35/A VSS 0.18fF
C56753 OR2X1_LOC_34/A VSS -0.08fF
C56754 OR2X1_LOC_89/Y VSS 0.11fF
C56755 OR2X1_LOC_67/A VSS 0.43fF
C56756 OR2X1_LOC_78/Y VSS 0.19fF
C56757 OR2X1_LOC_78/B VSS 0.54fF
C56758 OR2X1_LOC_78/A VSS 0.95fF
C56759 OR2X1_LOC_56/Y VSS 0.04fF
C56760 OR2X1_LOC_829/A VSS 0.26fF
C56761 OR2X1_LOC_847/B VSS 0.16fF
C56762 AND2X1_LOC_852/B VSS -0.41fF
C56763 AND2X1_LOC_807/B VSS -0.17fF
C56764 OR2X1_LOC_392/B VSS 0.65fF
C56765 OR2X1_LOC_571/B VSS 0.28fF
C56766 OR2X1_LOC_523/Y VSS 0.13fF
C56767 OR2X1_LOC_561/Y VSS 0.28fF
C56768 OR2X1_LOC_581/Y VSS 0.08fF
C56769 OR2X1_LOC_346/A VSS 0.20fF
C56770 OR2X1_LOC_294/Y VSS 0.29fF
C56771 AND2X1_LOC_287/B VSS 0.19fF
C56772 OR2X1_LOC_234/Y VSS 0.11fF
C56773 OR2X1_LOC_232/Y VSS 0.06fF
C56774 OR2X1_LOC_786/A VSS 0.34fF
C56775 AND2X1_LOC_65/A VSS -0.95fF
C56776 OR2X1_LOC_831/B VSS 0.50fF
C56777 AND2X1_LOC_273/a_8_24# VSS 0.10fF
C56778 OR2X1_LOC_155/A VSS -8.81fF
C56779 OR2X1_LOC_739/A VSS 0.34fF
C56780 OR2X1_LOC_795/B VSS 0.17fF
C56781 OR2X1_LOC_776/Y VSS 0.20fF
C56782 OR2X1_LOC_736/Y VSS 0.42fF
C56783 OR2X1_LOC_773/Y VSS 0.11fF
C56784 OR2X1_LOC_753/A VSS 0.74fF
C56785 OR2X1_LOC_803/B VSS -0.02fF
C56786 OR2X1_LOC_784/Y VSS -0.05fF
C56787 OR2X1_LOC_762/Y VSS 0.24fF
C56788 AND2X1_LOC_447/Y VSS 0.44fF
C56789 AND2X1_LOC_476/a_8_24# VSS 0.10fF
C56790 AND2X1_LOC_473/Y VSS -0.60fF
C56791 AND2X1_LOC_456/Y VSS 0.37fF
C56792 OR2X1_LOC_489/B VSS 0.22fF
C56793 AND2X1_LOC_487/a_8_24# VSS 0.10fF
C56794 AND2X1_LOC_95/Y VSS -4.24fF
C56795 OR2X1_LOC_501/B VSS -0.22fF
C56796 AND2X1_LOC_498/a_8_24# VSS 0.10fF
C56797 AND2X1_LOC_70/Y VSS 0.37fF
C56798 OR2X1_LOC_216/Y VSS -0.13fF
C56799 OR2X1_LOC_217/Y VSS 0.20fF
C56800 OR2X1_LOC_411/A VSS 0.15fF
C56801 OR2X1_LOC_214/B VSS 0.22fF
C56802 OR2X1_LOC_200/Y VSS 0.18fF
C56803 AND2X1_LOC_639/A VSS 0.27fF
C56804 AND2X1_LOC_635/a_8_24# VSS 0.10fF
C56805 OR2X1_LOC_582/Y VSS 0.08fF
C56806 AND2X1_LOC_645/A VSS 0.22fF
C56807 OR2X1_LOC_601/Y VSS 0.11fF
C56808 OR2X1_LOC_728/B VSS 0.26fF
C56809 OR2X1_LOC_620/A VSS -0.01fF
C56810 AND2X1_LOC_647/B VSS 0.17fF
C56811 OR2X1_LOC_609/Y VSS 0.08fF
C56812 AND2X1_LOC_574/A VSS 0.17fF
C56813 OR2X1_LOC_35/B VSS 0.11fF
C56814 OR2X1_LOC_33/B VSS -0.20fF
C56815 OR2X1_LOC_33/A VSS 0.15fF
C56816 OR2X1_LOC_99/Y VSS 0.22fF
C56817 OR2X1_LOC_88/Y VSS 0.31fF
C56818 OR2X1_LOC_66/Y VSS 0.16fF
C56819 OR2X1_LOC_46/A VSS 1.13fF
C56820 OR2X1_LOC_54/Y VSS 1.08fF
C56821 OR2X1_LOC_17/Y VSS 0.84fF
C56822 OR2X1_LOC_838/B VSS 0.22fF
C56823 OR2X1_LOC_846/A VSS 0.11fF
C56824 AND2X1_LOC_51/Y VSS 1.00fF
C56825 AND2X1_LOC_793/Y VSS 0.16fF
C56826 AND2X1_LOC_792/Y VSS -2.90fF
C56827 AND2X1_LOC_859/B VSS 0.26fF
C56828 AND2X1_LOC_845/Y VSS -4.38fF
C56829 OR2X1_LOC_593/A VSS 0.18fF
C56830 OR2X1_LOC_449/B VSS 0.54fF
C56831 OR2X1_LOC_562/Y VSS 0.18fF
C56832 OR2X1_LOC_343/B VSS 0.15fF
C56833 OR2X1_LOC_286/B VSS 0.28fF
C56834 OR2X1_LOC_814/A VSS 0.82fF
C56835 OR2X1_LOC_345/A VSS 0.15fF
C56836 OR2X1_LOC_585/A VSS 0.37fF
C56837 AND2X1_LOC_43/B VSS -4.45fF
C56838 AND2X1_LOC_31/Y VSS 0.61fF
C56839 OR2X1_LOC_804/A VSS 0.51fF
C56840 OR2X1_LOC_786/Y VSS -2.78fF
C56841 OR2X1_LOC_772/Y VSS 0.16fF
C56842 OR2X1_LOC_778/Y VSS 1.13fF
C56843 OR2X1_LOC_742/B VSS 0.24fF
C56844 OR2X1_LOC_739/Y VSS 0.18fF
C56845 OR2X1_LOC_751/A VSS 0.11fF
C56846 OR2X1_LOC_239/Y VSS 0.16fF
C56847 AND2X1_LOC_449/Y VSS 0.12fF
C56848 AND2X1_LOC_448/Y VSS 0.31fF
C56849 OR2X1_LOC_434/A VSS 0.31fF
C56850 AND2X1_LOC_431/a_8_24# VSS 0.10fF
C56851 AND2X1_LOC_474/Y VSS -0.28fF
C56852 AND2X1_LOC_458/Y VSS 0.07fF
C56853 AND2X1_LOC_72/B VSS 0.28fF
C56854 AND2X1_LOC_7/Y VSS -0.03fF
C56855 OR2X1_LOC_215/A VSS 0.08fF
C56856 OR2X1_LOC_201/Y VSS 0.15fF
C56857 OR2X1_LOC_124/Y VSS 0.44fF
C56858 AND2X1_LOC_9/a_8_24# VSS 0.10fF
C56859 OR2X1_LOC_99/A VSS 0.14fF
C56860 OR2X1_LOC_98/B VSS 0.10fF
C56861 AND2X1_LOC_648/B VSS 0.25fF
C56862 OR2X1_LOC_690/A VSS 0.76fF
C56863 OR2X1_LOC_602/A VSS 0.15fF
C56864 AND2X1_LOC_624/B VSS 0.24fF
C56865 AND2X1_LOC_620/Y VSS -0.16fF
C56866 OR2X1_LOC_615/Y VSS 0.41fF
C56867 OR2X1_LOC_720/B VSS 0.45fF
C56868 AND2X1_LOC_667/a_8_24# VSS 0.10fF
C56869 OR2X1_LOC_647/B VSS 0.30fF
C56870 OR2X1_LOC_610/Y VSS 0.06fF
C56871 AND2X1_LOC_647/Y VSS -0.25fF
C56872 AND2X1_LOC_216/A VSS -0.28fF
C56873 OR2X1_LOC_409/B VSS 0.69fF
C56874 OR2X1_LOC_408/Y VSS 0.13fF
C56875 OR2X1_LOC_65/Y VSS 0.10fF
C56876 OR2X1_LOC_87/Y VSS 0.19fF
C56877 AND2X1_LOC_848/Y VSS 0.16fF
C56878 AND2X1_LOC_795/Y VSS 0.31fF
C56879 OR2X1_LOC_846/B VSS 0.36fF
C56880 AND2X1_LOC_3/Y VSS 0.68fF
C56881 AND2X1_LOC_847/Y VSS 0.05fF
C56882 AND2X1_LOC_838/B VSS -0.15fF
C56883 OR2X1_LOC_826/Y VSS 0.07fF
C56884 OR2X1_LOC_7/Y VSS 0.33fF
C56885 OR2X1_LOC_591/A VSS 0.28fF
C56886 D_GATE_579 VSS 0.09fF
C56887 OR2X1_LOC_261/A VSS 0.02fF
C56888 AND2X1_LOC_260/a_8_24# VSS 0.10fF
C56889 OR2X1_LOC_285/A VSS 0.18fF
C56890 OR2X1_LOC_375/A VSS 0.75fF
C56891 OR2X1_LOC_270/Y VSS -0.04fF
C56892 OR2X1_LOC_269/Y VSS 0.06fF
C56893 OR2X1_LOC_750/A VSS -0.10fF
C56894 OR2X1_LOC_804/B VSS -0.01fF
C56895 OR2X1_LOC_787/Y VSS 0.13fF
C56896 OR2X1_LOC_796/B VSS 0.17fF
C56897 OR2X1_LOC_779/Y VSS 0.18fF
C56898 OR2X1_LOC_203/Y VSS 0.70fF
C56899 OR2X1_LOC_204/Y VSS 0.44fF
C56900 OR2X1_LOC_249/Y VSS 0.21fF
C56901 AND2X1_LOC_451/Y VSS 0.02fF
C56902 AND2X1_LOC_450/Y VSS 0.05fF
C56903 OR2X1_LOC_451/A VSS 0.15fF
C56904 AND2X1_LOC_472/B VSS 0.30fF
C56905 AND2X1_LOC_459/Y VSS 0.16fF
C56906 OR2X1_LOC_705/B VSS -0.86fF
C56907 AND2X1_LOC_485/a_8_24# VSS 0.10fF
C56908 OR2X1_LOC_778/A VSS 0.58fF
C56909 AND2X1_LOC_573/A VSS 0.05fF
C56910 AND2X1_LOC_677/a_8_24# VSS 0.10fF
C56911 OR2X1_LOC_75/Y VSS 0.19fF
C56912 OR2X1_LOC_99/B VSS 0.19fF
C56913 AND2X1_LOC_624/A VSS 0.48fF
C56914 AND2X1_LOC_621/Y VSS -1.20fF
C56915 OR2X1_LOC_619/Y VSS -3.41fF
C56916 OR2X1_LOC_599/Y VSS -0.03fF
C56917 OR2X1_LOC_597/Y VSS -0.14fF
C56918 AND2X1_LOC_660/A VSS 0.23fF
C56919 AND2X1_LOC_649/Y VSS -0.17fF
C56920 OR2X1_LOC_602/B VSS -0.16fF
C56921 OR2X1_LOC_719/A VSS 0.12fF
C56922 AND2X1_LOC_612/B VSS -0.12fF
C56923 AND2X1_LOC_633/a_8_24# VSS 0.10fF
C56924 OR2X1_LOC_118/Y VSS 0.23fF
C56925 OR2X1_LOC_419/Y VSS 0.53fF
C56926 OR2X1_LOC_22/A VSS -0.02fF
C56927 OR2X1_LOC_85/A VSS 0.98fF
C56928 OR2X1_LOC_70/A VSS 0.35fF
C56929 OR2X1_LOC_3/B VSS 0.31fF
C56930 OR2X1_LOC_51/B VSS 0.39fF
C56931 OR2X1_LOC_820/Y VSS 0.10fF
C56932 AND2X1_LOC_839/B VSS 0.07fF
C56933 OR2X1_LOC_824/Y VSS -0.16fF
C56934 AND2X1_LOC_862/A VSS 0.25fF
C56935 AND2X1_LOC_850/Y VSS 0.20fF
C56936 AND2X1_LOC_808/A VSS 0.29fF
C56937 AND2X1_LOC_796/Y VSS 0.02fF
C56938 OR2X1_LOC_815/A VSS 0.15fF
C56939 OR2X1_LOC_7/A VSS -29.87fF
C56940 OR2X1_LOC_368/A VSS 0.28fF
C56941 OR2X1_LOC_285/B VSS 0.21fF
C56942 OR2X1_LOC_346/B VSS 0.20fF
C56943 OR2X1_LOC_805/A VSS -2.11fF
C56944 OR2X1_LOC_774/B VSS 0.27fF
C56945 OR2X1_LOC_770/Y VSS 0.18fF
C56946 OR2X1_LOC_760/Y VSS -0.07fF
C56947 OR2X1_LOC_797/A VSS 0.18fF
C56948 OR2X1_LOC_781/Y VSS 0.12fF
C56949 OR2X1_LOC_486/B VSS -0.05fF
C56950 OR2X1_LOC_237/Y VSS 0.34fF
C56951 OR2X1_LOC_205/Y VSS 0.30fF
C56952 OR2X1_LOC_226/Y VSS 0.08fF
C56953 AND2X1_LOC_79/Y VSS -0.80fF
C56954 OR2X1_LOC_248/Y VSS 0.38fF
C56955 OR2X1_LOC_555/B VSS 0.46fF
C56956 OR2X1_LOC_430/Y VSS 0.07fF
C56957 AND2X1_LOC_440/a_8_24# VSS 0.10fF
C56958 AND2X1_LOC_675/A VSS 0.07fF
C56959 OR2X1_LOC_416/Y VSS -0.01fF
C56960 AND2X1_LOC_276/Y VSS -0.23fF
C56961 AND2X1_LOC_116/Y VSS 0.25fF
C56962 OR2X1_LOC_679/B VSS -0.08fF
C56963 AND2X1_LOC_687/a_8_24# VSS 0.10fF
C56964 AND2X1_LOC_698/a_8_24# VSS 0.10fF
C56965 AND2X1_LOC_650/Y VSS 0.13fF
C56966 AND2X1_LOC_649/B VSS 0.18fF
C56967 OR2X1_LOC_595/Y VSS 0.06fF
C56968 AND2X1_LOC_665/a_8_24# VSS 0.10fF
C56969 OR2X1_LOC_52/Y VSS 0.19fF
C56970 OR2X1_LOC_65/B VSS -0.60fF
C56971 OR2X1_LOC_86/A VSS 0.42fF
C56972 OR2X1_LOC_95/Y VSS 0.79fF
C56973 AND2X1_LOC_631/Y VSS 0.12fF
C56974 OR2X1_LOC_612/B VSS 0.18fF
C56975 OR2X1_LOC_828/B VSS 0.25fF
C56976 OR2X1_LOC_41/Y VSS 0.39fF
C56977 OR2X1_LOC_112/B VSS -0.80fF
C56978 AND2X1_LOC_798/Y VSS 0.11fF
C56979 AND2X1_LOC_853/Y VSS 0.19fF
C56980 AND2X1_LOC_852/Y VSS -0.73fF
C56981 AND2X1_LOC_848/A VSS -0.77fF
C56982 OR2X1_LOC_815/Y VSS -0.03fF
C56983 OR2X1_LOC_845/A VSS 0.26fF
C56984 AND2X1_LOC_839/A VSS 0.16fF
C56985 AND2X1_LOC_19/a_8_24# VSS 0.10fF
C56986 AND2X1_LOC_824/B VSS 0.22fF
C56987 OR2X1_LOC_781/A VSS 0.13fF
C56988 AND2X1_LOC_462/B VSS 0.28fF
C56989 AND2X1_LOC_461/a_8_24# VSS 0.10fF
C56990 AND2X1_LOC_476/A VSS 0.79fF
C56991 AND2X1_LOC_462/Y VSS 0.22fF
C56992 OR2X1_LOC_383/Y VSS 0.04fF
C56993 OR2X1_LOC_219/B VSS 0.47fF
C56994 AND2X1_LOC_72/Y VSS 0.14fF
C56995 OR2X1_LOC_247/Y VSS 0.16fF
C56996 OR2X1_LOC_417/A VSS -3.77fF
C56997 OR2X1_LOC_258/Y VSS -0.08fF
C56998 OR2X1_LOC_89/A VSS 0.77fF
C56999 OR2X1_LOC_427/Y VSS 0.22fF
C57000 OR2X1_LOC_426/Y VSS 0.06fF
C57001 OR2X1_LOC_440/A VSS 0.57fF
C57002 OR2X1_LOC_544/A VSS 0.21fF
C57003 AND2X1_LOC_687/B VSS 0.06fF
C57004 OR2X1_LOC_684/Y VSS 0.34fF
C57005 OR2X1_LOC_683/Y VSS 0.06fF
C57006 AND2X1_LOC_661/A VSS 0.33fF
C57007 AND2X1_LOC_520/Y VSS 0.22fF
C57008 AND2X1_LOC_675/a_8_24# VSS 0.10fF
C57009 OR2X1_LOC_674/Y VSS 0.12fF
C57010 AND2X1_LOC_620/a_8_24# VSS 0.10fF
C57011 AND2X1_LOC_483/Y VSS 0.15fF
C57012 OR2X1_LOC_428/Y VSS 0.01fF
C57013 OR2X1_LOC_84/Y VSS 0.20fF
C57014 OR2X1_LOC_84/A VSS -0.02fF
C57015 OR2X1_LOC_74/A VSS -6.14fF
C57016 OR2X1_LOC_11/Y VSS 0.81fF
C57017 OR2X1_LOC_2/Y VSS 0.49fF
C57018 AND2X1_LOC_108/a_8_24# VSS 0.10fF
C57019 OR2X1_LOC_532/B VSS 0.64fF
C57020 OR2X1_LOC_609/A VSS 0.29fF
C57021 AND2X1_LOC_840/B VSS 0.34fF
C57022 AND2X1_LOC_834/a_8_24# VSS 0.10fF
C57023 OR2X1_LOC_511/Y VSS 0.17fF
C57024 AND2X1_LOC_809/A VSS 0.10fF
C57025 OR2X1_LOC_761/Y VSS 0.06fF
C57026 GATE_811 VSS 0.19fF
C57027 AND2X1_LOC_811/Y VSS 0.29fF
C57028 AND2X1_LOC_810/Y VSS 0.32fF
C57029 AND2X1_LOC_863/A VSS 0.05fF
C57030 OR2X1_LOC_836/B VSS 0.13fF
C57031 AND2X1_LOC_823/a_8_24# VSS 0.10fF
C57032 OR2X1_LOC_813/Y VSS 0.15fF
C57033 AND2X1_LOC_721/A VSS -2.03fF
C57034 D_INPUT_0 VSS 0.77fF
C57035 INPUT_1 VSS 0.98fF
C57036 OR2X1_LOC_87/B VSS 0.30fF
C57037 AND2X1_LOC_290/a_8_24# VSS 0.10fF
C57038 OR2X1_LOC_792/A VSS 0.38fF
C57039 OR2X1_LOC_783/A VSS 0.30fF
C57040 OR2X1_LOC_780/B VSS 0.36fF
C57041 OR2X1_LOC_780/A VSS 0.15fF
C57042 OR2X1_LOC_279/Y VSS 0.27fF
C57043 OR2X1_LOC_427/A VSS 1.39fF
C57044 AND2X1_LOC_463/B VSS 0.17fF
C57045 AND2X1_LOC_460/a_8_24# VSS 0.10fF
C57046 OR2X1_LOC_409/Y VSS 0.02fF
C57047 AND2X1_LOC_465/Y VSS 0.28fF
C57048 AND2X1_LOC_464/Y VSS -0.13fF
C57049 AND2X1_LOC_717/B VSS -0.59fF
C57050 OR2X1_LOC_491/Y VSS 0.06fF
C57051 OR2X1_LOC_833/B VSS 0.07fF
C57052 OR2X1_LOC_224/Y VSS 0.08fF
C57053 OR2X1_LOC_31/Y VSS 0.86fF
C57054 OR2X1_LOC_206/A VSS 0.12fF
C57055 AND2X1_LOC_67/Y VSS 0.33fF
C57056 AND2X1_LOC_69/Y VSS 0.13fF
C57057 OR2X1_LOC_235/Y VSS -0.14fF
C57058 OR2X1_LOC_220/A VSS -0.06fF
C57059 OR2X1_LOC_405/Y VSS 0.26fF
C57060 OR2X1_LOC_416/A VSS 0.31fF
C57061 AND2X1_LOC_687/A VSS 0.38fF
C57062 OR2X1_LOC_681/Y VSS 0.06fF
C57063 OR2X1_LOC_708/B VSS 0.13fF
C57064 AND2X1_LOC_696/a_8_24# VSS 0.10fF
C57065 AND2X1_LOC_653/B VSS 0.07fF
C57066 AND2X1_LOC_593/Y VSS 0.32fF
C57067 AND2X1_LOC_468/B VSS 0.29fF
C57068 GATE_662 VSS 0.24fF
C57069 AND2X1_LOC_632/A VSS 0.05fF
C57070 AND2X1_LOC_629/Y VSS 0.23fF
C57071 OR2X1_LOC_628/Y VSS 0.19fF
C57072 OR2X1_LOC_675/A VSS 0.32fF
C57073 OR2X1_LOC_453/A VSS 0.18fF
C57074 OR2X1_LOC_449/A VSS 0.46fF
C57075 OR2X1_LOC_61/Y VSS 0.30fF
C57076 OR2X1_LOC_71/Y VSS 0.50fF
C57077 OR2X1_LOC_96/B VSS -0.20fF
C57078 OR2X1_LOC_113/A VSS 0.21fF
C57079 OR2X1_LOC_633/B VSS -0.12fF
C57080 AND2X1_LOC_118/a_8_24# VSS 0.10fF
C57081 OR2X1_LOC_130/A VSS 0.75fF
C57082 OR2X1_LOC_618/Y VSS 0.12fF
C57083 AND2X1_LOC_801/B VSS -0.07fF
C57084 AND2X1_LOC_687/Y VSS 0.29fF
C57085 AND2X1_LOC_856/B VSS 0.19fF
C57086 OR2X1_LOC_829/Y VSS 0.07fF
C57087 AND2X1_LOC_729/B VSS -0.76fF
C57088 AND2X1_LOC_822/a_8_24# VSS 0.10fF
C57089 AND2X1_LOC_807/Y VSS 0.60fF
C57090 AND2X1_LOC_840/A VSS 0.21fF
C57091 OR2X1_LOC_495/Y VSS 0.13fF
C57092 GATE_865 VSS 0.02fF
C57093 AND2X1_LOC_849/A VSS 0.19fF
C57094 AND2X1_LOC_844/a_8_24# VSS 0.10fF
C57095 AND2X1_LOC_523/Y VSS -0.64fF
C57096 OR2X1_LOC_793/A VSS 0.11fF
C57097 OR2X1_LOC_220/B VSS 0.18fF
C57098 OR2X1_LOC_289/Y VSS 0.09fF
C57099 D_GATE_222 VSS 0.02fF
C57100 OR2X1_LOC_246/A VSS 0.99fF
C57101 OR2X1_LOC_47/Y VSS 1.86fF
C57102 AND2X1_LOC_477/A VSS 0.23fF
C57103 OR2X1_LOC_555/A VSS 0.12fF
C57104 OR2X1_LOC_493/A VSS 0.22fF
C57105 OR2X1_LOC_707/A VSS 0.15fF
C57106 OR2X1_LOC_437/Y VSS 0.26fF
C57107 OR2X1_LOC_415/A VSS 0.13fF
C57108 OR2X1_LOC_26/Y VSS -4.00fF
C57109 OR2X1_LOC_402/Y VSS 0.24fF
C57110 AND2X1_LOC_654/B VSS 0.30fF
C57111 AND2X1_LOC_638/Y VSS -0.03fF
C57112 AND2X1_LOC_634/Y VSS -0.16fF
C57113 AND2X1_LOC_633/Y VSS -0.10fF
C57114 AND2X1_LOC_663/B VSS -3.54fF
C57115 AND2X1_LOC_660/Y VSS 0.08fF
C57116 OR2X1_LOC_672/Y VSS 0.26fF
C57117 OR2X1_LOC_670/Y VSS 0.06fF
C57118 OR2X1_LOC_463/B VSS -0.00fF
C57119 OR2X1_LOC_459/B VSS 0.14fF
C57120 OR2X1_LOC_448/B VSS 0.21fF
C57121 OR2X1_LOC_448/A VSS 0.21fF
C57122 OR2X1_LOC_83/A VSS 0.20fF
C57123 AND2X1_LOC_141/A VSS 0.16fF
C57124 AND2X1_LOC_47/Y VSS 0.78fF
C57125 OR2X1_LOC_125/Y VSS 0.06fF
C57126 OR2X1_LOC_123/B VSS 0.12fF
C57127 AND2X1_LOC_856/A VSS 0.06fF
C57128 AND2X1_LOC_354/B VSS 0.16fF
C57129 AND2X1_LOC_866/B VSS 0.11fF
C57130 AND2X1_LOC_862/Y VSS 0.08fF
C57131 OR2X1_LOC_607/Y VSS 0.06fF
C57132 OR2X1_LOC_629/A VSS 0.20fF
C57133 AND2X1_LOC_841/B VSS -0.56fF
C57134 OR2X1_LOC_34/B VSS 0.16fF
C57135 OR2X1_LOC_87/A VSS 0.90fF
C57136 OR2X1_LOC_194/B VSS 0.12fF
C57137 OR2X1_LOC_335/B VSS 0.41fF
C57138 OR2X1_LOC_299/Y VSS 0.08fF
C57139 OR2X1_LOC_212/A VSS -0.28fF
C57140 OR2X1_LOC_223/A VSS -0.45fF
C57141 OR2X1_LOC_218/Y VSS 0.59fF
C57142 OR2X1_LOC_278/A VSS 0.40fF
C57143 OR2X1_LOC_267/A VSS 0.11fF
C57144 OR2X1_LOC_256/A VSS -0.09fF
C57145 OR2X1_LOC_291/A VSS 0.75fF
C57146 OR2X1_LOC_286/Y VSS 0.17fF
C57147 GATE_479 VSS 0.03fF
C57148 AND2X1_LOC_479/Y VSS 0.15fF
C57149 OR2X1_LOC_193/Y VSS 0.07fF
C57150 OR2X1_LOC_194/Y VSS 0.05fF
C57151 OR2X1_LOC_707/B VSS 0.27fF
C57152 AND2X1_LOC_425/Y VSS 0.39fF
C57153 AND2X1_LOC_662/B VSS 0.23fF
C57154 AND2X1_LOC_654/Y VSS -1.24fF
C57155 OR2X1_LOC_673/A VSS 0.21fF
C57156 OR2X1_LOC_435/Y VSS 0.14fF
C57157 OR2X1_LOC_80/Y VSS 0.26fF
C57158 OR2X1_LOC_464/A VSS 0.19fF
C57159 OR2X1_LOC_404/A VSS 0.14fF
C57160 AND2X1_LOC_641/Y VSS 0.18fF
C57161 AND2X1_LOC_640/Y VSS 0.37fF
C57162 OR2X1_LOC_468/Y VSS 0.53fF
C57163 OR2X1_LOC_506/A VSS 0.85fF
C57164 OR2X1_LOC_447/A VSS 0.15fF
C57165 OR2X1_LOC_426/A VSS 0.36fF
C57166 AND2X1_LOC_797/A VSS 0.26fF
C57167 AND2X1_LOC_148/Y VSS 0.14fF
C57168 AND2X1_LOC_147/Y VSS -0.18fF
C57169 AND2X1_LOC_139/B VSS -0.31fF
C57170 AND2X1_LOC_114/Y VSS 0.06fF
C57171 OR2X1_LOC_106/A VSS 0.49fF
C57172 AND2X1_LOC_105/a_8_24# VSS 0.10fF
C57173 OR2X1_LOC_92/Y VSS 0.90fF
C57174 AND2X1_LOC_866/A VSS 0.30fF
C57175 AND2X1_LOC_863/Y VSS 0.15fF
C57176 AND2X1_LOC_853/a_8_24# VSS 0.10fF
C57177 OR2X1_LOC_847/A VSS 0.00fF
C57178 OR2X1_LOC_818/Y VSS 0.06fF
C57179 AND2X1_LOC_850/A VSS -0.13fF
C57180 AND2X1_LOC_842/a_8_24# VSS 0.10fF
C57181 OR2X1_LOC_184/Y VSS 0.32fF
C57182 OR2X1_LOC_651/A VSS -1.01fF
C57183 OR2X1_LOC_606/Y VSS 0.10fF
C57184 OR2X1_LOC_121/B VSS 0.70fF
C57185 OR2X1_LOC_617/Y VSS 0.25fF
C57186 AND2X1_LOC_25/Y VSS 0.21fF
C57187 AND2X1_LOC_11/Y VSS -0.50fF
C57188 OR2X1_LOC_62/B VSS 0.42fF
C57189 AND2X1_LOC_42/B VSS 0.72fF
C57190 AND2X1_LOC_37/a_8_24# VSS 0.10fF
C57191 AND2X1_LOC_798/A VSS 0.15fF
C57192 AND2X1_LOC_318/Y VSS 0.35fF
C57193 AND2X1_LOC_727/A VSS -0.65fF
C57194 AND2X1_LOC_307/Y VSS 0.07fF
C57195 OR2X1_LOC_810/A VSS -4.69fF
C57196 OR2X1_LOC_802/Y VSS 0.10fF
C57197 OR2X1_LOC_288/A VSS -0.17fF
C57198 OR2X1_LOC_557/A VSS -1.01fF
C57199 OR2X1_LOC_223/B VSS 0.21fF
C57200 OR2X1_LOC_739/B VSS 0.17fF
C57201 OR2X1_LOC_517/A VSS 0.72fF
C57202 OR2X1_LOC_473/A VSS 0.45fF
C57203 OR2X1_LOC_276/B VSS 0.21fF
C57204 OR2X1_LOC_276/A VSS 0.14fF
C57205 OR2X1_LOC_244/A VSS -1.70fF
C57206 OR2X1_LOC_243/B VSS 0.10fF
C57207 OR2X1_LOC_456/A VSS 0.34fF
C57208 OR2X1_LOC_213/A VSS 0.04fF
C57209 OR2X1_LOC_436/Y VSS 0.37fF
C57210 OR2X1_LOC_475/Y VSS 0.45fF
C57211 OR2X1_LOC_476/Y VSS 0.18fF
C57212 OR2X1_LOC_464/B VSS 0.17fF
C57213 OR2X1_LOC_457/B VSS 0.09fF
C57214 OR2X1_LOC_706/A VSS -0.32fF
C57215 AND2X1_LOC_693/a_8_24# VSS 0.10fF
C57216 AND2X1_LOC_656/Y VSS 0.08fF
C57217 AND2X1_LOC_672/B VSS 0.19fF
C57218 OR2X1_LOC_19/B VSS -4.13fF
C57219 OR2X1_LOC_413/Y VSS 0.02fF
C57220 OR2X1_LOC_435/B VSS -0.06fF
C57221 OR2X1_LOC_401/Y VSS 0.19fF
C57222 OR2X1_LOC_146/Y VSS 0.22fF
C57223 OR2X1_LOC_145/Y VSS 0.06fF
C57224 AND2X1_LOC_116/B VSS -0.15fF
C57225 AND2X1_LOC_126/a_8_24# VSS 0.10fF
C57226 AND2X1_LOC_139/A VSS -0.23fF
C57227 AND2X1_LOC_137/a_8_24# VSS 0.10fF
C57228 OR2X1_LOC_655/A VSS 0.18fF
C57229 OR2X1_LOC_643/Y VSS 0.19fF
C57230 OR2X1_LOC_605/B VSS -0.17fF
C57231 OR2X1_LOC_605/A VSS 0.30fF
C57232 OR2X1_LOC_36/Y VSS 0.85fF
C57233 OR2X1_LOC_616/Y VSS -0.21fF
C57234 OR2X1_LOC_18/Y VSS 1.25fF
C57235 AND2X1_LOC_857/Y VSS 0.08fF
C57236 AND2X1_LOC_851/B VSS 0.21fF
C57237 AND2X1_LOC_841/a_8_24# VSS 0.10fF
C57238 AND2X1_LOC_831/Y VSS -2.49fF
C57239 AND2X1_LOC_842/B VSS 0.24fF
C57240 AND2X1_LOC_852/a_8_24# VSS 0.10fF
C57241 AND2X1_LOC_838/Y VSS -0.06fF
C57242 OR2X1_LOC_651/B VSS 0.11fF
C57243 OR2X1_LOC_637/Y VSS -0.01fF
C57244 AND2X1_LOC_21/Y VSS 0.28fF
C57245 OR2X1_LOC_61/B VSS 0.24fF
C57246 D_INPUT_3 VSS 0.73fF
C57247 D_INPUT_2 VSS 0.50fF
C57248 OR2X1_LOC_68/Y VSS 0.07fF
C57249 AND2X1_LOC_307/a_8_24# VSS 0.10fF
C57250 OR2X1_LOC_304/Y VSS -0.06fF
C57251 OR2X1_LOC_355/B VSS 0.11fF
C57252 OR2X1_LOC_316/Y VSS 0.10fF
C57253 OR2X1_LOC_315/Y VSS 0.38fF
C57254 OR2X1_LOC_811/A VSS -1.96fF
C57255 OR2X1_LOC_820/A VSS 0.29fF
C57256 OR2X1_LOC_62/A VSS 0.23fF
C57257 OR2X1_LOC_275/A VSS 0.06fF
C57258 OR2X1_LOC_285/Y VSS 0.18fF
C57259 OR2X1_LOC_221/A VSS 0.16fF
C57260 OR2X1_LOC_231/A VSS 0.13fF
C57261 OR2X1_LOC_244/B VSS 0.22fF
C57262 OR2X1_LOC_506/B VSS 0.28fF
C57263 OR2X1_LOC_241/Y VSS 0.15fF
C57264 OR2X1_LOC_64/Y VSS 1.27fF
C57265 OR2X1_LOC_436/B VSS 0.08fF
C57266 OR2X1_LOC_174/A VSS 0.38fF
C57267 OR2X1_LOC_455/A VSS -0.05fF
C57268 OR2X1_LOC_772/B VSS 0.15fF
C57269 OR2X1_LOC_706/B VSS 0.16fF
C57270 AND2X1_LOC_670/a_8_24# VSS 0.10fF
C57271 OR2X1_LOC_470/A VSS 0.18fF
C57272 OR2X1_LOC_469/Y VSS -0.35fF
C57273 OR2X1_LOC_477/Y VSS 0.11fF
C57274 OR2X1_LOC_91/A VSS -4.30fF
C57275 OR2X1_LOC_401/B VSS 0.14fF
C57276 OR2X1_LOC_401/A VSS 0.18fF
C57277 OR2X1_LOC_210/B VSS 0.16fF
C57278 OR2X1_LOC_144/Y VSS 0.07fF
C57279 AND2X1_LOC_170/B VSS 0.19fF
C57280 OR2X1_LOC_167/Y VSS 0.27fF
C57281 AND2X1_LOC_114/a_8_24# VSS 0.10fF
C57282 AND2X1_LOC_113/Y VSS 0.15fF
C57283 OR2X1_LOC_655/B VSS 0.11fF
C57284 OR2X1_LOC_754/A VSS -0.10fF
C57285 AND2X1_LOC_851/A VSS 0.10fF
C57286 AND2X1_LOC_858/B VSS 0.38fF
C57287 AND2X1_LOC_79/a_8_24# VSS 0.10fF
C57288 AND2X1_LOC_859/Y VSS -1.05fF
C57289 OR2X1_LOC_637/B VSS 0.26fF
C57290 OR2X1_LOC_637/A VSS -0.06fF
C57291 OR2X1_LOC_193/A VSS 0.51fF
C57292 AND2X1_LOC_13/a_8_24# VSS 0.10fF
C57293 AND2X1_LOC_35/Y VSS 0.43fF
C57294 AND2X1_LOC_34/Y VSS 0.27fF
C57295 AND2X1_LOC_33/Y VSS 0.06fF
C57296 AND2X1_LOC_57/a_8_24# VSS 0.10fF
C57297 AND2X1_LOC_24/a_8_24# VSS 0.10fF
C57298 AND2X1_LOC_319/A VSS 0.54fF
C57299 OR2X1_LOC_314/Y VSS 0.22fF
C57300 OR2X1_LOC_313/Y VSS 0.22fF
C57301 D_INPUT_4 VSS -1.44fF
C57302 OR2X1_LOC_503/Y VSS -0.00fF
C57303 AND2X1_LOC_227/Y VSS 0.22fF
C57304 OR2X1_LOC_274/Y VSS 0.07fF
C57305 OR2X1_LOC_541/A VSS 0.37fF
C57306 OR2X1_LOC_813/A VSS 0.44fF
C57307 OR2X1_LOC_22/Y VSS 0.85fF
C57308 OR2X1_LOC_296/Y VSS 0.19fF
C57309 OR2X1_LOC_252/Y VSS -0.09fF
C57310 OR2X1_LOC_411/Y VSS 0.22fF
C57311 OR2X1_LOC_444/B VSS 0.16fF
C57312 OR2X1_LOC_443/Y VSS 0.19fF
C57313 OR2X1_LOC_488/Y VSS 0.22fF
C57314 OR2X1_LOC_465/B VSS 0.10fF
C57315 OR2X1_LOC_76/Y VSS 0.37fF
C57316 OR2X1_LOC_500/A VSS 0.18fF
C57317 OR2X1_LOC_403/A VSS 0.18fF
C57318 OR2X1_LOC_690/Y VSS 0.24fF
C57319 OR2X1_LOC_689/Y VSS 0.06fF
C57320 OR2X1_LOC_422/Y VSS 0.08fF
C57321 OR2X1_LOC_471/Y VSS -0.77fF
C57322 OR2X1_LOC_470/B VSS 0.14fF
C57323 OR2X1_LOC_453/Y VSS 0.17fF
C57324 OR2X1_LOC_165/Y VSS 0.08fF
C57325 OR2X1_LOC_164/Y VSS 0.40fF
C57326 AND2X1_LOC_179/a_8_24# VSS 0.10fF
C57327 OR2X1_LOC_148/A VSS 0.12fF
C57328 AND2X1_LOC_8/Y VSS 0.59fF
C57329 AND2X1_LOC_572/A VSS 0.23fF
C57330 AND2X1_LOC_123/Y VSS 0.08fF
C57331 OR2X1_LOC_103/Y VSS 0.26fF
C57332 AND2X1_LOC_865/A VSS -0.05fF
C57333 AND2X1_LOC_658/A VSS -1.46fF
C57334 OR2X1_LOC_669/Y VSS 0.28fF
C57335 OR2X1_LOC_669/A VSS 0.26fF
C57336 OR2X1_LOC_625/Y VSS 0.08fF
C57337 OR2X1_LOC_659/A VSS 0.25fF
C57338 OR2X1_LOC_624/Y VSS 0.34fF
C57339 OR2X1_LOC_197/A VSS 0.05fF
C57340 AND2X1_LOC_53/Y VSS 0.86fF
C57341 OR2X1_LOC_196/B VSS 0.48fF
C57342 OR2X1_LOC_79/A VSS -0.10fF
C57343 AND2X1_LOC_78/a_8_24# VSS 0.10fF
C57344 OR2X1_LOC_97/B VSS 0.20fF
C57345 AND2X1_LOC_89/a_8_24# VSS 0.10fF
C57346 AND2X1_LOC_843/Y VSS 0.02fF
C57347 OR2X1_LOC_639/A VSS 0.18fF
C57348 OR2X1_LOC_636/B VSS -0.47fF
C57349 OR2X1_LOC_636/A VSS -0.13fF
C57350 AND2X1_LOC_23/a_8_24# VSS 0.10fF
C57351 OR2X1_LOC_32/Y VSS 0.12fF
C57352 AND2X1_LOC_305/a_8_24# VSS 0.10fF
C57353 AND2X1_LOC_338/a_8_24# VSS 0.10fF
C57354 AND2X1_LOC_334/Y VSS 0.11fF
C57355 AND2X1_LOC_359/B VSS 0.19fF
C57356 AND2X1_LOC_342/Y VSS -0.23fF
C57357 OR2X1_LOC_852/A VSS 0.18fF
C57358 OR2X1_LOC_835/Y VSS 0.14fF
C57359 OR2X1_LOC_836/Y VSS 0.18fF
C57360 OR2X1_LOC_817/Y VSS 0.06fF
C57361 OR2X1_LOC_807/A VSS 0.10fF
C57362 OR2X1_LOC_362/B VSS 0.42fF
C57363 AND2X1_LOC_510/A VSS 0.04fF
C57364 OR2X1_LOC_520/A VSS 0.14fF
C57365 AND2X1_LOC_48/A VSS 0.55fF
C57366 OR2X1_LOC_273/Y VSS 0.26fF
C57367 OR2X1_LOC_743/A VSS 0.42fF
C57368 OR2X1_LOC_262/Y VSS 0.22fF
C57369 OR2X1_LOC_243/A VSS 0.18fF
C57370 OR2X1_LOC_240/B VSS 0.17fF
C57371 OR2X1_LOC_287/A VSS 0.02fF
C57372 OR2X1_LOC_542/B VSS 0.42fF
C57373 OR2X1_LOC_295/Y VSS 0.08fF
C57374 OR2X1_LOC_481/A VSS -0.16fF
C57375 OR2X1_LOC_498/Y VSS 0.16fF
C57376 OR2X1_LOC_189/A VSS -0.47fF
C57377 AND2X1_LOC_690/a_8_24# VSS 0.10fF
C57378 OR2X1_LOC_545/B VSS 0.04fF
C57379 OR2X1_LOC_473/Y VSS -0.24fF
C57380 OR2X1_LOC_487/Y VSS 0.06fF
C57381 OR2X1_LOC_456/Y VSS 0.09fF
C57382 OR2X1_LOC_466/A VSS 0.21fF
C57383 OR2X1_LOC_446/Y VSS 0.37fF
C57384 OR2X1_LOC_447/Y VSS 0.48fF
C57385 OR2X1_LOC_158/B VSS 0.15fF
C57386 AND2X1_LOC_155/Y VSS 0.30fF
C57387 AND2X1_LOC_154/Y VSS 0.26fF
C57388 OR2X1_LOC_148/B VSS 0.16fF
C57389 AND2X1_LOC_123/a_8_24# VSS 0.10fF
C57390 OR2X1_LOC_117/Y VSS 0.17fF
C57391 OR2X1_LOC_181/B VSS 0.14fF
C57392 AND2X1_LOC_715/A VSS 0.55fF
C57393 OR2X1_LOC_111/Y VSS 0.26fF
C57394 OR2X1_LOC_647/A VSS 0.23fF
C57395 OR2X1_LOC_646/A VSS 0.08fF
C57396 OR2X1_LOC_659/B VSS 0.47fF
C57397 OR2X1_LOC_510/Y VSS 0.05fF
C57398 AND2X1_LOC_861/B VSS 0.27fF
C57399 AND2X1_LOC_474/A VSS -0.42fF
C57400 OR2X1_LOC_679/Y VSS 0.07fF
C57401 OR2X1_LOC_679/A VSS 0.00fF
C57402 OR2X1_LOC_613/Y VSS 0.32fF
C57403 AND2X1_LOC_51/A VSS -0.04fF
C57404 OR2X1_LOC_20/Y VSS 0.06fF
C57405 AND2X1_LOC_56/B VSS 0.91fF
C57406 AND2X1_LOC_99/Y VSS 0.15fF
C57407 AND2X1_LOC_98/Y VSS 0.32fF
C57408 OR2X1_LOC_639/B VSS 0.27fF
C57409 OR2X1_LOC_307/B VSS 0.12fF
C57410 AND2X1_LOC_352/B VSS 0.14fF
C57411 AND2X1_LOC_335/Y VSS 0.08fF
C57412 AND2X1_LOC_326/a_8_24# VSS 0.10fF
C57413 AND2X1_LOC_345/Y VSS -0.32fF
C57414 AND2X1_LOC_363/A VSS 0.24fF
C57415 AND2X1_LOC_348/Y VSS -0.03fF
C57416 OR2X1_LOC_852/B VSS 0.17fF
C57417 OR2X1_LOC_837/Y VSS -0.22fF
C57418 OR2X1_LOC_816/Y VSS 0.01fF
C57419 OR2X1_LOC_51/Y VSS 1.81fF
C57420 OR2X1_LOC_859/A VSS -1.35fF
C57421 OR2X1_LOC_844/Y VSS 0.03fF
C57422 OR2X1_LOC_827/Y VSS -0.06fF
C57423 OR2X1_LOC_43/A VSS 1.00fF
C57424 OR2X1_LOC_807/B VSS -0.02fF
C57425 OR2X1_LOC_792/Y VSS 0.10fF
C57426 AND2X1_LOC_508/B VSS 0.16fF
C57427 AND2X1_LOC_507/a_8_24# VSS 0.10fF
C57428 OR2X1_LOC_505/Y VSS 0.12fF
C57429 OR2X1_LOC_504/Y VSS 0.06fF
C57430 OR2X1_LOC_520/B VSS 0.24fF
C57431 AND2X1_LOC_518/a_8_24# VSS 0.10fF
C57432 OR2X1_LOC_272/Y VSS -0.25fF
C57433 OR2X1_LOC_283/Y VSS 0.22fF
C57434 OR2X1_LOC_250/Y VSS 0.30fF
C57435 AND2X1_LOC_41/A VSS 0.69fF
C57436 OR2X1_LOC_600/A VSS 1.12fF
C57437 OR2X1_LOC_497/Y VSS 0.26fF
C57438 OR2X1_LOC_474/Y VSS -1.48fF
C57439 OR2X1_LOC_471/B VSS 0.17fF
C57440 OR2X1_LOC_431/Y VSS 0.16fF
C57441 OR2X1_LOC_420/Y VSS -0.12fF
C57442 OR2X1_LOC_448/Y VSS 0.53fF
C57443 OR2X1_LOC_147/A VSS 0.04fF
C57444 AND2X1_LOC_207/A VSS 0.10fF
C57445 AND2X1_LOC_196/Y VSS 0.20fF
C57446 OR2X1_LOC_169/B VSS 0.15fF
C57447 AND2X1_LOC_166/a_8_24# VSS 0.10fF
C57448 AND2X1_LOC_122/a_8_24# VSS 0.10fF
C57449 AND2X1_LOC_101/B VSS 0.30fF
C57450 OR2X1_LOC_86/Y VSS -0.09fF
C57451 OR2X1_LOC_624/A VSS 1.10fF
C57452 OR2X1_LOC_620/Y VSS 0.52fF
C57453 OR2X1_LOC_640/A VSS 0.27fF
C57454 OR2X1_LOC_334/B VSS -0.03fF
C57455 OR2X1_LOC_634/A VSS 0.38fF
C57456 OR2X1_LOC_648/A VSS 0.33fF
C57457 OR2X1_LOC_602/Y VSS 0.40fF
C57458 OR2X1_LOC_647/Y VSS 0.16fF
C57459 OR2X1_LOC_689/A VSS 0.35fF
C57460 OR2X1_LOC_678/Y VSS -0.13fF
C57461 OR2X1_LOC_834/A VSS 0.40fF
C57462 OR2X1_LOC_611/Y VSS 0.18fF
C57463 AND2X1_LOC_21/a_8_24# VSS 0.10fF
C57464 OR2X1_LOC_195/A VSS 0.21fF
C57465 AND2X1_LOC_43/a_8_24# VSS 0.10fF
C57466 AND2X1_LOC_76/Y VSS 0.25fF
C57467 OR2X1_LOC_74/Y VSS 0.06fF
C57468 INPUT_0 VSS -4.74fF
C57469 OR2X1_LOC_96/Y VSS 0.10fF
C57470 OR2X1_LOC_93/Y VSS 0.06fF
C57471 OR2X1_LOC_88/A VSS 0.02fF
C57472 OR2X1_LOC_32/B VSS 0.52fF
C57473 OR2X1_LOC_201/A VSS 0.15fF
C57474 AND2X1_LOC_337/B VSS 0.27fF
C57475 OR2X1_LOC_312/Y VSS 0.25fF
C57476 OR2X1_LOC_317/A VSS 0.15fF
C57477 AND2X1_LOC_326/B VSS 0.16fF
C57478 AND2X1_LOC_325/a_8_24# VSS 0.10fF
C57479 AND2X1_LOC_358/a_8_24# VSS 0.10fF
C57480 AND2X1_LOC_351/Y VSS 0.26fF
C57481 AND2X1_LOC_350/Y VSS 0.12fF
C57482 OR2X1_LOC_297/Y VSS 0.06fF
C57483 OR2X1_LOC_837/B VSS 0.17fF
C57484 OR2X1_LOC_837/A VSS 0.14fF
C57485 OR2X1_LOC_808/A VSS -0.64fF
C57486 OR2X1_LOC_859/B VSS 0.18fF
C57487 OR2X1_LOC_862/A VSS 0.08fF
C57488 AND2X1_LOC_538/Y VSS 0.07fF
C57489 AND2X1_LOC_537/Y VSS -0.35fF
C57490 OR2X1_LOC_620/B VSS -0.01fF
C57491 OR2X1_LOC_559/B VSS 0.19fF
C57492 AND2X1_LOC_517/a_8_24# VSS 0.10fF
C57493 AND2X1_LOC_508/A VSS -0.18fF
C57494 AND2X1_LOC_711/A VSS 0.29fF
C57495 OR2X1_LOC_282/Y VSS 0.08fF
C57496 OR2X1_LOC_485/A VSS -2.58fF
C57497 OR2X1_LOC_271/Y VSS 0.26fF
C57498 OR2X1_LOC_271/B VSS 0.06fF
C57499 OR2X1_LOC_260/Y VSS 0.10fF
C57500 OR2X1_LOC_441/Y VSS 0.33fF
C57501 OR2X1_LOC_404/Y VSS -0.73fF
C57502 OR2X1_LOC_472/A VSS -1.25fF
C57503 OR2X1_LOC_460/Y VSS 0.18fF
C57504 OR2X1_LOC_467/A VSS -0.19fF
C57505 OR2X1_LOC_450/Y VSS 0.08fF
C57506 OR2X1_LOC_429/Y VSS -1.29fF
C57507 AND2X1_LOC_154/a_8_24# VSS 0.10fF
C57508 AND2X1_LOC_208/B VSS 0.20fF
C57509 AND2X1_LOC_197/Y VSS 0.08fF
C57510 OR2X1_LOC_57/Y VSS 0.06fF
C57511 AND2X1_LOC_110/a_8_24# VSS 0.10fF
C57512 OR2X1_LOC_168/A VSS 0.15fF
C57513 AND2X1_LOC_176/a_8_24# VSS 0.10fF
C57514 OR2X1_LOC_191/B VSS 0.25fF
C57515 OR2X1_LOC_137/B VSS 0.14fF
C57516 OR2X1_LOC_502/A VSS 0.69fF
C57517 OR2X1_LOC_122/A VSS 0.15fF
C57518 OR2X1_LOC_666/A VSS 0.41fF
C57519 OR2X1_LOC_426/B VSS -6.72fF
C57520 OR2X1_LOC_648/B VSS 0.62fF
C57521 OR2X1_LOC_688/Y VSS 0.07fF
C57522 OR2X1_LOC_660/B VSS 0.21fF
C57523 OR2X1_LOC_624/B VSS 0.26fF
C57524 OR2X1_LOC_748/A VSS -1.10fF
C57525 AND2X1_LOC_99/A VSS 0.24fF
C57526 AND2X1_LOC_97/a_8_24# VSS 0.10fF
C57527 OR2X1_LOC_677/Y VSS 0.20fF
C57528 OR2X1_LOC_600/Y VSS -0.33fF
C57529 AND2X1_LOC_1/Y VSS 0.46fF
C57530 AND2X1_LOC_53/a_8_24# VSS 0.10fF
C57531 D_INPUT_5 VSS 0.10fF
C57532 AND2X1_LOC_19/Y VSS 0.25fF
C57533 OR2X1_LOC_76/A VSS -0.02fF
C57534 AND2X1_LOC_75/a_8_24# VSS 0.10fF
C57535 AND2X1_LOC_42/a_8_24# VSS 0.10fF
C57536 OR2X1_LOC_380/A VSS 0.16fF
C57537 AND2X1_LOC_364/A VSS 0.32fF
C57538 AND2X1_LOC_357/a_8_24# VSS 0.10fF
C57539 AND2X1_LOC_313/a_8_24# VSS 0.10fF
C57540 AND2X1_LOC_326/A VSS 0.15fF
C57541 OR2X1_LOC_321/Y VSS 0.07fF
C57542 OR2X1_LOC_320/Y VSS 0.24fF
C57543 AND2X1_LOC_303/B VSS 0.08fF
C57544 AND2X1_LOC_302/a_8_24# VSS 0.10fF
C57545 OR2X1_LOC_298/Y VSS 0.12fF
C57546 OR2X1_LOC_310/Y VSS 0.08fF
C57547 AND2X1_LOC_347/B VSS 0.24fF
C57548 OR2X1_LOC_836/A VSS 0.25fF
C57549 OR2X1_LOC_814/Y VSS 0.07fF
C57550 OR2X1_LOC_862/B VSS 0.20fF
C57551 OR2X1_LOC_825/Y VSS 0.21fF
C57552 OR2X1_LOC_848/A VSS -4.79fF
C57553 OR2X1_LOC_808/B VSS 0.90fF
C57554 AND2X1_LOC_538/a_8_24# VSS 0.10fF
C57555 OR2X1_LOC_311/Y VSS 0.32fF
C57556 OR2X1_LOC_574/A VSS 0.95fF
C57557 OR2X1_LOC_547/B VSS -0.03fF
C57558 AND2X1_LOC_548/Y VSS 0.11fF
C57559 OR2X1_LOC_531/Y VSS 0.06fF
C57560 OR2X1_LOC_507/A VSS 0.13fF
C57561 AND2X1_LOC_712/B VSS 0.19fF
C57562 OR2X1_LOC_696/Y VSS 0.28fF
C57563 OR2X1_LOC_666/Y VSS 0.18fF
C57564 OR2X1_LOC_665/Y VSS 0.01fF
C57565 OR2X1_LOC_292/Y VSS 0.15fF
C57566 OR2X1_LOC_468/A VSS -0.01fF
C57567 OR2X1_LOC_440/B VSS 0.16fF
C57568 OR2X1_LOC_472/B VSS -0.09fF
C57569 OR2X1_LOC_461/Y VSS 0.18fF
C57570 OR2X1_LOC_216/A VSS -0.21fF
C57571 OR2X1_LOC_484/Y VSS 0.24fF
C57572 OR2X1_LOC_452/A VSS 0.18fF
C57573 AND2X1_LOC_211/B VSS 0.20fF
C57574 OR2X1_LOC_173/Y VSS 0.06fF
C57575 OR2X1_LOC_680/A VSS -4.91fF
C57576 OR2X1_LOC_147/B VSS -0.99fF
C57577 OR2X1_LOC_168/B VSS 0.25fF
C57578 OR2X1_LOC_140/A VSS 0.29fF
C57579 OR2X1_LOC_698/Y VSS -0.11fF
C57580 OR2X1_LOC_744/A VSS 1.31fF
C57581 OR2X1_LOC_661/A VSS 0.18fF
C57582 OR2X1_LOC_650/Y VSS 0.25fF
C57583 OR2X1_LOC_643/A VSS 0.16fF
C57584 OR2X1_LOC_630/Y VSS 0.22fF
C57585 OR2X1_LOC_622/A VSS 0.10fF
C57586 OR2X1_LOC_621/B VSS -0.11fF
C57587 OR2X1_LOC_621/A VSS -0.06fF
C57588 OR2X1_LOC_755/A VSS 0.20fF
C57589 AND2X1_LOC_86/B VSS 0.43fF
C57590 OR2X1_LOC_76/B VSS 0.24fF
C57591 AND2X1_LOC_74/a_8_24# VSS 0.10fF
C57592 OR2X1_LOC_98/A VSS 0.15fF
C57593 AND2X1_LOC_94/Y VSS 0.39fF
C57594 OR2X1_LOC_676/Y VSS 0.43fF
C57595 OR2X1_LOC_598/Y VSS 0.45fF
C57596 AND2X1_LOC_30/a_8_24# VSS 0.10fF
C57597 INPUT_4 VSS 0.40fF
C57598 AND2X1_LOC_390/B VSS 0.02fF
C57599 OR2X1_LOC_387/Y VSS -0.00fF
C57600 OR2X1_LOC_385/Y VSS 0.12fF
C57601 AND2X1_LOC_365/A VSS 0.20fF
C57602 AND2X1_LOC_354/Y VSS 0.08fF
C57603 OR2X1_LOC_459/A VSS 0.12fF
C57604 AND2X1_LOC_378/a_8_24# VSS 0.10fF
C57605 AND2X1_LOC_377/Y VSS 0.07fF
C57606 AND2X1_LOC_110/Y VSS 0.19fF
C57607 OR2X1_LOC_291/Y VSS 0.23fF
C57608 OR2X1_LOC_261/Y VSS 0.14fF
C57609 AND2X1_LOC_259/Y VSS 0.49fF
C57610 GATE_366 VSS 0.14fF
C57611 OR2X1_LOC_109/Y VSS 0.27fF
C57612 OR2X1_LOC_703/A VSS -0.23fF
C57613 AND2X1_LOC_301/a_8_24# VSS 0.10fF
C57614 OR2X1_LOC_863/A VSS 0.18fF
C57615 OR2X1_LOC_835/B VSS 0.24fF
C57616 OR2X1_LOC_835/A VSS 0.15fF
C57617 OR2X1_LOC_798/Y VSS 0.28fF
C57618 OR2X1_LOC_848/B VSS 0.05fF
C57619 OR2X1_LOC_536/Y VSS 0.07fF
C57620 AND2X1_LOC_514/Y VSS -1.44fF
C57621 OR2X1_LOC_417/Y VSS -0.57fF
C57622 OR2X1_LOC_530/Y VSS 0.07fF
C57623 OR2X1_LOC_529/Y VSS -0.01fF
C57624 AND2X1_LOC_560/B VSS 0.18fF
C57625 OR2X1_LOC_517/Y VSS 0.06fF
C57626 OR2X1_LOC_507/B VSS 0.20fF
C57627 AND2X1_LOC_722/A VSS 0.29fF
C57628 AND2X1_LOC_605/Y VSS 0.19fF
C57629 OR2X1_LOC_695/Y VSS 0.07fF
C57630 OR2X1_LOC_694/Y VSS 0.21fF
C57631 OR2X1_LOC_280/Y VSS 0.33fF
C57632 OR2X1_LOC_476/B VSS -1.86fF
C57633 OR2X1_LOC_631/B VSS 0.42fF
C57634 OR2X1_LOC_254/B VSS 0.28fF
C57635 OR2X1_LOC_450/B VSS 0.01fF
C57636 OR2X1_LOC_450/A VSS 0.10fF
C57637 OR2X1_LOC_467/B VSS -0.48fF
C57638 OR2X1_LOC_162/Y VSS 0.07fF
C57639 AND2X1_LOC_196/a_8_24# VSS 0.10fF
C57640 OR2X1_LOC_48/Y VSS 0.20fF
C57641 OR2X1_LOC_151/Y VSS 0.08fF
C57642 AND2X1_LOC_175/B VSS 0.00fF
C57643 AND2X1_LOC_174/a_8_24# VSS 0.10fF
C57644 OR2X1_LOC_131/A VSS 0.32fF
C57645 OR2X1_LOC_589/A VSS 0.93fF
C57646 OR2X1_LOC_664/Y VSS 0.30fF
C57647 OR2X1_LOC_185/A VSS 1.40fF
C57648 OR2X1_LOC_697/Y VSS -0.19fF
C57649 OR2X1_LOC_687/A VSS 0.22fF
C57650 OR2X1_LOC_686/B VSS 0.20fF
C57651 OR2X1_LOC_686/A VSS -0.19fF
C57652 OR2X1_LOC_649/B VSS 0.14fF
C57653 OR2X1_LOC_462/B VSS 0.36fF
C57654 OR2X1_LOC_520/Y VSS 0.53fF
C57655 OR2X1_LOC_632/A VSS 0.18fF
C57656 AND2X1_LOC_84/a_8_24# VSS 0.10fF
C57657 OR2X1_LOC_83/Y VSS -0.10fF
C57658 OR2X1_LOC_81/Y VSS 0.08fF
C57659 OR2X1_LOC_108/Y VSS 0.43fF
C57660 AND2X1_LOC_356/B VSS 0.16fF
C57661 OR2X1_LOC_538/A VSS 0.52fF
C57662 OR2X1_LOC_325/B VSS 0.49fF
C57663 AND2X1_LOC_338/A VSS 0.10fF
C57664 OR2X1_LOC_403/B VSS 0.26fF
C57665 AND2X1_LOC_348/A VSS 0.24fF
C57666 OR2X1_LOC_256/Y VSS -0.17fF
C57667 AND2X1_LOC_456/B VSS 0.45fF
C57668 AND2X1_LOC_367/B VSS 0.02fF
C57669 AND2X1_LOC_363/Y VSS -0.22fF
C57670 OR2X1_LOC_831/A VSS 0.39fF
C57671 OR2X1_LOC_863/B VSS 0.21fF
C57672 OR2X1_LOC_849/A VSS -0.41fF
C57673 OR2X1_LOC_673/Y VSS 0.37fF
C57674 OR2X1_LOC_823/Y VSS -0.14fF
C57675 OR2X1_LOC_840/A VSS -4.67fF
C57676 OR2X1_LOC_809/B VSS 0.41fF
C57677 OR2X1_LOC_800/Y VSS 0.18fF
C57678 D_GATE_811 VSS 0.18fF
C57679 OR2X1_LOC_546/B VSS 0.16fF
C57680 OR2X1_LOC_537/A VSS -0.01fF
C57681 OR2X1_LOC_527/Y VSS 0.15fF
C57682 AND2X1_LOC_577/A VSS 0.22fF
C57683 AND2X1_LOC_565/Y VSS 0.12fF
C57684 OR2X1_LOC_509/A VSS -0.07fF
C57685 AND2X1_LOC_503/a_8_24# VSS 0.10fF
C57686 AND2X1_LOC_561/B VSS 0.08fF
C57687 OR2X1_LOC_494/Y VSS 0.02fF
C57688 OR2X1_LOC_693/Y VSS 0.07fF
C57689 OR2X1_LOC_692/Y VSS 0.13fF
C57690 AND2X1_LOC_728/a_8_24# VSS 0.10fF
C57691 OR2X1_LOC_680/Y VSS -0.07fF
C57692 AND2X1_LOC_740/B VSS 0.13fF
C57693 AND2X1_LOC_192/Y VSS 0.24fF
C57694 OR2X1_LOC_290/Y VSS 0.19fF
C57695 OR2X1_LOC_493/B VSS 0.10fF
C57696 OR2X1_LOC_482/Y VSS 0.60fF
C57697 OR2X1_LOC_465/Y VSS 0.19fF
C57698 AND2X1_LOC_161/Y VSS -0.11fF
C57699 AND2X1_LOC_160/Y VSS 0.20fF
C57700 AND2X1_LOC_199/A VSS -0.11fF
C57701 OR2X1_LOC_43/Y VSS 0.07fF
C57702 OR2X1_LOC_175/B VSS 0.23fF
C57703 OR2X1_LOC_190/A VSS -0.35fF
C57704 AND2X1_LOC_141/B VSS 0.36fF
C57705 OR2X1_LOC_131/Y VSS -0.31fF
C57706 AND2X1_LOC_554/B VSS -0.06fF
C57707 OR2X1_LOC_653/A VSS 0.13fF
C57708 OR2X1_LOC_799/A VSS 0.22fF
C57709 OR2X1_LOC_329/B VSS -2.21fF
C57710 D_GATE_662 VSS 0.21fF
C57711 OR2X1_LOC_659/Y VSS -0.00fF
C57712 OR2X1_LOC_687/B VSS 0.17fF
C57713 OR2X1_LOC_685/B VSS 0.11fF
C57714 OR2X1_LOC_685/A VSS 0.21fF
C57715 OR2X1_LOC_629/Y VSS 0.09fF
C57716 AND2X1_LOC_61/Y VSS -0.47fF
C57717 OR2X1_LOC_60/Y VSS 0.07fF
C57718 OR2X1_LOC_58/Y VSS 0.13fF
C57719 AND2X1_LOC_82/Y VSS 0.16fF
C57720 OR2X1_LOC_107/Y VSS -0.09fF
C57721 OR2X1_LOC_324/A VSS 0.05fF
C57722 AND2X1_LOC_367/A VSS 0.43fF
C57723 AND2X1_LOC_364/Y VSS -0.85fF
C57724 OR2X1_LOC_389/A VSS 0.23fF
C57725 AND2X1_LOC_339/B VSS 0.23fF
C57726 OR2X1_LOC_135/Y VSS 0.34fF
C57727 AND2X1_LOC_349/B VSS 0.15fF
C57728 AND2X1_LOC_343/a_8_24# VSS 0.10fF
C57729 OR2X1_LOC_251/Y VSS 0.24fF
C57730 OR2X1_LOC_399/A VSS 0.15fF
C57731 OR2X1_LOC_856/A VSS 0.17fF
C57732 OR2X1_LOC_691/Y VSS -0.34fF
C57733 OR2X1_LOC_687/Y VSS 0.27fF
C57734 OR2X1_LOC_800/A VSS -0.07fF
C57735 OR2X1_LOC_499/B VSS 0.40fF
C57736 OR2X1_LOC_822/Y VSS 0.07fF
C57737 D_GATE_865 VSS 0.08fF
C57738 OR2X1_LOC_865/Y VSS 0.18fF
C57739 OR2X1_LOC_812/A VSS 0.18fF
C57740 OR2X1_LOC_807/Y VSS 0.27fF
C57741 AND2X1_LOC_578/A VSS 0.26fF
C57742 AND2X1_LOC_568/a_8_24# VSS 0.10fF
C57743 AND2X1_LOC_566/Y VSS 0.20fF
C57744 AND2X1_LOC_580/B VSS 0.36fF
C57745 AND2X1_LOC_576/Y VSS -1.59fF
C57746 AND2X1_LOC_575/Y VSS 0.10fF
C57747 AND2X1_LOC_550/A VSS 0.35fF
C57748 OR2X1_LOC_525/Y VSS 0.19fF
C57749 OR2X1_LOC_516/B VSS 0.21fF
C57750 AND2X1_LOC_513/a_8_24# VSS 0.10fF
C57751 AND2X1_LOC_512/Y VSS 0.14fF
C57752 OR2X1_LOC_545/A VSS 0.04fF
C57753 OR2X1_LOC_490/Y VSS 0.10fF
C57754 AND2X1_LOC_489/Y VSS 0.28fF
C57755 OR2X1_LOC_503/A VSS 0.21fF
C57756 AND2X1_LOC_731/Y VSS -0.20fF
C57757 AND2X1_LOC_716/a_8_24# VSS 0.10fF
C57758 AND2X1_LOC_303/A VSS 0.29fF
C57759 AND2X1_LOC_228/Y VSS 0.38fF
C57760 AND2X1_LOC_705/a_8_24# VSS 0.10fF
C57761 OR2X1_LOC_526/Y VSS -0.09fF
C57762 OR2X1_LOC_485/Y VSS 0.47fF
C57763 OR2X1_LOC_492/Y VSS 0.10fF
C57764 OR2X1_LOC_481/Y VSS 0.14fF
C57765 OR2X1_LOC_3/Y VSS 0.84fF
C57766 OR2X1_LOC_477/B VSS 0.11fF
C57767 OR2X1_LOC_39/Y VSS -0.02fF
C57768 OR2X1_LOC_151/A VSS -4.85fF
C57769 AND2X1_LOC_183/a_8_24# VSS 0.10fF
C57770 OR2X1_LOC_633/Y VSS 0.02fF
C57771 OR2X1_LOC_663/A VSS -0.17fF
C57772 OR2X1_LOC_660/Y VSS 0.10fF
C57773 OR2X1_LOC_673/B VSS -0.11fF
C57774 OR2X1_LOC_654/A VSS -0.15fF
C57775 OR2X1_LOC_61/A VSS 0.15fF
C57776 OR2X1_LOC_377/A VSS -5.63fF
C57777 AND2X1_LOC_71/a_8_24# VSS 0.10fF
C57778 OR2X1_LOC_235/B VSS 0.22fF
C57779 AND2X1_LOC_93/a_8_24# VSS 0.10fF
C57780 AND2X1_LOC_387/B VSS 0.20fF
C57781 AND2X1_LOC_17/Y VSS -0.81fF
C57782 OR2X1_LOC_376/A VSS 0.15fF
C57783 OR2X1_LOC_402/B VSS -0.16fF
C57784 OR2X1_LOC_70/Y VSS 1.33fF
C57785 OR2X1_LOC_141/B VSS 0.29fF
C57786 OR2X1_LOC_137/Y VSS 0.18fF
C57787 OR2X1_LOC_128/B VSS 0.11fF
C57788 OR2X1_LOC_128/A VSS 0.15fF
C57789 OR2X1_LOC_330/Y VSS 0.07fF
C57790 OR2X1_LOC_324/B VSS 0.10fF
C57791 AND2X1_LOC_320/a_8_24# VSS 0.10fF
C57792 AND2X1_LOC_357/B VSS 0.19fF
C57793 AND2X1_LOC_566/B VSS -1.48fF
C57794 AND2X1_LOC_364/a_8_24# VSS 0.10fF
C57795 AND2X1_LOC_358/Y VSS 0.15fF
C57796 OR2X1_LOC_246/Y VSS -0.18fF
C57797 OR2X1_LOC_856/B VSS 0.30fF
C57798 OR2X1_LOC_354/A VSS 0.19fF
C57799 OR2X1_LOC_841/A VSS 0.06fF
C57800 OR2X1_LOC_821/Y VSS -0.22fF
C57801 OR2X1_LOC_850/A VSS 0.16fF
C57802 OR2X1_LOC_287/B VSS 0.33fF
C57803 OR2X1_LOC_812/B VSS -0.51fF
C57804 AND2X1_LOC_551/B VSS 0.07fF
C57805 OR2X1_LOC_524/Y VSS 0.66fF
C57806 AND2X1_LOC_568/B VSS 0.00fF
C57807 AND2X1_LOC_535/Y VSS 0.34fF
C57808 OR2X1_LOC_535/A VSS -0.16fF
C57809 OR2X1_LOC_592/A VSS 0.15fF
C57810 AND2X1_LOC_589/a_8_24# VSS 0.10fF
C57811 AND2X1_LOC_580/A VSS -0.49fF
C57812 AND2X1_LOC_577/Y VSS 0.23fF
C57813 AND2X1_LOC_562/B VSS 0.19fF
C57814 AND2X1_LOC_556/a_8_24# VSS 0.10fF
C57815 OR2X1_LOC_309/Y VSS 0.19fF
C57816 AND2X1_LOC_512/a_8_24# VSS 0.10fF
C57817 OR2X1_LOC_521/Y VSS 0.09fF
C57818 AND2X1_LOC_500/Y VSS 0.09fF
C57819 AND2X1_LOC_714/B VSS 0.22fF
C57820 AND2X1_LOC_711/Y VSS 0.27fF
C57821 OR2X1_LOC_152/Y VSS -0.33fF
C57822 AND2X1_LOC_702/Y VSS 0.05fF
C57823 OR2X1_LOC_789/B VSS 0.16fF
C57824 AND2X1_LOC_734/Y VSS 0.27fF
C57825 AND2X1_LOC_733/Y VSS -0.27fF
C57826 OR2X1_LOC_792/B VSS 0.10fF
C57827 OR2X1_LOC_758/Y VSS -0.01fF
C57828 VDD VSS 2.10fF
C57829 D_GATE_479 VSS 0.04fF
C57830 OR2X1_LOC_478/Y VSS 0.17fF
C57831 OR2X1_LOC_479/Y VSS 0.60fF
C57832 AND2X1_LOC_160/a_8_24# VSS 0.10fF
C57833 AND2X1_LOC_181/Y VSS 0.25fF
C57834 OR2X1_LOC_333/B VSS 0.39fF
C57835 OR2X1_LOC_662/A VSS 0.12fF
C57836 OR2X1_LOC_653/Y VSS 0.17fF
C57837 OR2X1_LOC_640/Y VSS 0.17fF
C57838 OR2X1_LOC_641/Y VSS 0.49fF
C57839 OR2X1_LOC_158/A VSS 1.15fF
C57840 OR2X1_LOC_671/Y VSS 0.63fF
C57841 OR2X1_LOC_84/B VSS 0.03fF
C57842 AND2X1_LOC_2/Y VSS 0.18fF
C57843 AND2X1_LOC_357/A VSS 0.22fF
C57844 AND2X1_LOC_212/A VSS 0.29fF
C57845 AND2X1_LOC_350/B VSS -0.25fF
C57846 AND2X1_LOC_231/Y VSS 0.18fF
C57847 OR2X1_LOC_389/B VSS 0.23fF
C57848 OR2X1_LOC_160/B VSS 0.98fF
C57849 OR2X1_LOC_139/A VSS -3.02fF
C57850 OR2X1_LOC_702/A VSS 0.56fF
C57851 OR2X1_LOC_114/Y VSS 0.09fF
C57852 OR2X1_LOC_127/Y VSS 0.11fF
C57853 OR2X1_LOC_105/Y VSS 0.34fF
C57854 OR2X1_LOC_756/B VSS 0.79fF
C57855 OR2X1_LOC_331/A VSS 0.14fF
C57856 OR2X1_LOC_797/B VSS 0.38fF
C57857 OR2X1_LOC_148/Y VSS 0.18fF
C57858 OR2X1_LOC_857/A VSS 0.09fF
C57859 OR2X1_LOC_175/Y VSS -1.06fF
C57860 OR2X1_LOC_841/B VSS 0.08fF
C57861 OR2X1_LOC_850/B VSS 0.18fF
C57862 OR2X1_LOC_866/B VSS 0.38fF
C57863 OR2X1_LOC_774/Y VSS 0.24fF
C57864 OR2X1_LOC_318/Y VSS 0.39fF
C57865 OR2X1_LOC_638/B VSS 0.22fF
C57866 AND2X1_LOC_170/Y VSS 0.12fF
C57867 OR2X1_LOC_438/Y VSS 0.29fF
C57868 AND2X1_LOC_577/a_8_24# VSS 0.10fF
C57869 AND2X1_LOC_570/Y VSS -0.24fF
C57870 AND2X1_LOC_22/Y VSS 0.72fF
C57871 OR2X1_LOC_512/A VSS 0.38fF
C57872 AND2X1_LOC_732/B VSS -0.02fF
C57873 AND2X1_LOC_713/Y VSS 0.15fF
C57874 AND2X1_LOC_712/Y VSS 0.06fF
C57875 AND2X1_LOC_724/A VSS 0.21fF
C57876 AND2X1_LOC_703/Y VSS 0.08fF
C57877 OR2X1_LOC_764/Y VSS 0.07fF
C57878 OR2X1_LOC_763/Y VSS 0.11fF
C57879 OR2X1_LOC_782/B VSS 0.16fF
C57880 AND2X1_LOC_735/Y VSS -0.04fF
C57881 AND2X1_LOC_675/Y VSS -1.14fF
C57882 OR2X1_LOC_759/A VSS 0.04fF
C57883 OR2X1_LOC_40/Y VSS 1.36fF
C57884 AND2X1_LOC_191/Y VSS -1.39fF
C57885 OR2X1_LOC_189/Y VSS 0.12fF
C57886 AND2X1_LOC_168/Y VSS -0.26fF
C57887 OR2X1_LOC_178/Y VSS 0.19fF
C57888 OR2X1_LOC_682/Y VSS 0.20fF
C57889 OR2X1_LOC_656/Y VSS -0.61fF
C57890 OR2X1_LOC_6/B VSS 1.05fF
C57891 OR2X1_LOC_97/A VSS 0.37fF
C57892 AND2X1_LOC_81/B VSS -0.49fF
C57893 AND2X1_LOC_80/a_8_24# VSS 0.10fF
C57894 OR2X1_LOC_768/A VSS 0.26fF
C57895 OR2X1_LOC_604/A VSS 1.27fF
C57896 OR2X1_LOC_9/Y VSS 0.52fF
C57897 AND2X1_LOC_339/Y VSS 0.23fF
C57898 AND2X1_LOC_338/Y VSS 0.14fF
C57899 AND2X1_LOC_59/Y VSS 1.20fF
C57900 AND2X1_LOC_40/Y VSS 1.37fF
C57901 AND2X1_LOC_366/A VSS 0.19fF
C57902 OR2X1_LOC_116/A VSS 0.18fF
C57903 OR2X1_LOC_8/Y VSS 0.94fF
C57904 OR2X1_LOC_857/B VSS 0.26fF
C57905 OR2X1_LOC_864/A VSS -0.59fF
C57906 OR2X1_LOC_851/A VSS 0.20fF
C57907 OR2X1_LOC_842/A VSS 0.11fF
C57908 OR2X1_LOC_114/B VSS 0.53fF
C57909 OR2X1_LOC_318/A VSS 0.21fF
C57910 AND2X1_LOC_588/B VSS -0.04fF
C57911 D_INPUT_7 VSS 0.12fF
C57912 OR2X1_LOC_599/A VSS 0.86fF
C57913 AND2X1_LOC_549/Y VSS 0.10fF
C57914 OR2X1_LOC_523/B VSS 0.16fF
C57915 AND2X1_LOC_521/a_8_24# VSS 0.10fF
C57916 OR2X1_LOC_106/Y VSS 0.20fF
C57917 AND2X1_LOC_572/Y VSS 0.05fF
C57918 AND2X1_LOC_571/Y VSS 0.10fF
C57919 AND2X1_LOC_509/Y VSS 0.03fF
C57920 OR2X1_LOC_329/Y VSS 0.08fF
C57921 OR2X1_LOC_308/A VSS 0.18fF
C57922 AND2X1_LOC_772/B VSS 0.35fF
C57923 AND2X1_LOC_706/Y VSS 0.20fF
C57924 AND2X1_LOC_705/Y VSS -0.59fF
C57925 AND2X1_LOC_715/Y VSS -5.71fF
C57926 AND2X1_LOC_702/a_8_24# VSS 0.10fF
C57927 OR2X1_LOC_45/Y VSS 0.39fF
C57928 OR2X1_LOC_791/A VSS 0.18fF
C57929 OR2X1_LOC_756/Y VSS 0.10fF
C57930 AND2X1_LOC_658/B VSS 0.41fF
C57931 AND2X1_LOC_501/Y VSS -0.05fF
C57932 AND2X1_LOC_182/A VSS 0.30fF
C57933 OR2X1_LOC_187/Y VSS -0.14fF
C57934 OR2X1_LOC_136/Y VSS 0.06fF
C57935 OR2X1_LOC_170/A VSS 0.18fF
C57936 OR2X1_LOC_703/B VSS 0.59fF
C57937 OR2X1_LOC_113/Y VSS 0.19fF
C57938 AND2X1_LOC_340/Y VSS -0.29fF
C57939 OR2X1_LOC_494/A VSS 0.43fF
C57940 OR2X1_LOC_400/A VSS 0.14fF
C57941 OR2X1_LOC_160/A VSS 0.58fF
C57942 OR2X1_LOC_458/B VSS 0.24fF
C57943 AND2X1_LOC_372/a_8_24# VSS 0.10fF
C57944 AND2X1_LOC_362/B VSS 0.28fF
C57945 OR2X1_LOC_149/B VSS -0.05fF
C57946 OR2X1_LOC_858/A VSS -1.81fF
C57947 OR2X1_LOC_851/B VSS 0.16fF
C57948 OR2X1_LOC_833/Y VSS 0.15fF
C57949 OR2X1_LOC_865/A VSS 0.15fF
C57950 OR2X1_LOC_644/B VSS 0.20fF
C57951 OR2X1_LOC_596/Y VSS 0.07fF
C57952 OR2X1_LOC_319/B VSS 0.08fF
C57953 AND2X1_LOC_552/A VSS 0.10fF
C57954 AND2X1_LOC_542/a_8_24# VSS 0.10fF
C57955 AND2X1_LOC_569/A VSS 0.05fF
C57956 AND2X1_LOC_563/A VSS 0.15fF
C57957 AND2X1_LOC_541/Y VSS 0.14fF
C57958 AND2X1_LOC_574/Y VSS 0.06fF
C57959 AND2X1_LOC_573/Y VSS 0.08fF
C57960 OR2X1_LOC_306/Y VSS 0.37fF
C57961 OR2X1_LOC_781/B VSS 0.10fF
C57962 AND2X1_LOC_721/Y VSS -2.77fF
C57963 OR2X1_LOC_406/Y VSS 0.16fF
C57964 OR2X1_LOC_496/Y VSS 0.19fF
C57965 OR2X1_LOC_773/B VSS 0.19fF
C57966 OR2X1_LOC_751/Y VSS 0.10fF
C57967 OR2X1_LOC_757/A VSS -0.53fF
C57968 AND2X1_LOC_756/a_8_24# VSS 0.10fF
C57969 OR2X1_LOC_510/A VSS -0.62fF
C57970 AND2X1_LOC_707/Y VSS 0.06fF
C57971 OR2X1_LOC_710/A VSS 0.18fF
C57972 AND2X1_LOC_723/a_8_24# VSS 0.10fF
C57973 AND2X1_LOC_717/Y VSS -0.04fF
C57974 AND2X1_LOC_716/Y VSS -5.02fF
C57975 AND2X1_LOC_191/B VSS -0.86fF
C57976 AND2X1_LOC_190/a_8_24# VSS 0.10fF
C57977 OR2X1_LOC_691/B VSS 0.20fF
C57978 OR2X1_LOC_691/A VSS 0.30fF
C57979 OR2X1_LOC_400/B VSS 0.16fF
C57980 OR2X1_LOC_154/A VSS -10.29fF
C57981 OR2X1_LOC_179/Y VSS -0.09fF
C57982 OR2X1_LOC_124/B VSS -0.01fF
C57983 OR2X1_LOC_391/B VSS 0.33fF
C57984 AND2X1_LOC_363/B VSS -0.09fF
C57985 AND2X1_LOC_347/Y VSS 0.20fF
C57986 OR2X1_LOC_865/B VSS 0.36fF
C57987 OR2X1_LOC_860/Y VSS -0.10fF
C57988 OR2X1_LOC_858/B VSS 0.09fF
C57989 OR2X1_LOC_597/A VSS 0.29fF
C57990 OR2X1_LOC_421/A VSS 0.14fF
C57991 AND2X1_LOC_585/a_8_24# VSS 0.10fF
C57992 AND2X1_LOC_564/B VSS 0.19fF
C57993 AND2X1_LOC_543/Y VSS 0.14fF
C57994 AND2X1_LOC_554/Y VSS -0.32fF
C57995 OR2X1_LOC_351/B VSS 0.33fF
C57996 OR2X1_LOC_405/A VSS 0.50fF
C57997 OR2X1_LOC_264/Y VSS 0.59fF
C57998 OR2X1_LOC_359/A VSS 0.18fF
C57999 OR2X1_LOC_548/A VSS 0.15fF
C58000 OR2X1_LOC_305/Y VSS 0.24fF
C58001 OR2X1_LOC_519/Y VSS 0.16fF
C58002 OR2X1_LOC_710/B VSS 0.14fF
C58003 AND2X1_LOC_794/B VSS 0.19fF
C58004 OR2X1_LOC_533/Y VSS 0.19fF
C58005 AND2X1_LOC_802/B VSS 0.20fF
C58006 AND2X1_LOC_539/Y VSS -0.29fF
C58007 AND2X1_LOC_784/A VSS 0.56fF
C58008 AND2X1_LOC_777/a_8_24# VSS 0.10fF
C58009 AND2X1_LOC_723/Y VSS 0.05fF
C58010 AND2X1_LOC_722/Y VSS -0.13fF
C58011 AND2X1_LOC_719/Y VSS 1.03fF
C58012 OR2X1_LOC_770/A VSS 0.33fF
C58013 AND2X1_LOC_91/B VSS 0.75fF
C58014 AND2X1_LOC_64/Y VSS 0.61fF
C58015 OR2X1_LOC_791/B VSS 0.32fF
C58016 AND2X1_LOC_710/Y VSS 0.11fF
C58017 OR2X1_LOC_506/Y VSS 0.25fF
C58018 AND2X1_LOC_787/A VSS 0.08fF
C58019 AND2X1_LOC_817/B VSS 0.16fF
C58020 AND2X1_LOC_12/Y VSS -4.37fF
C58021 INPUT_3 VSS 0.35fF
C58022 AND2X1_LOC_391/Y VSS 0.44fF
C58023 OR2X1_LOC_715/B VSS 0.83fF
C58024 OR2X1_LOC_134/Y VSS 0.19fF
C58025 OR2X1_LOC_656/B VSS 0.53fF
C58026 OR2X1_LOC_100/Y VSS 0.29fF
C58027 OR2X1_LOC_124/A VSS 0.22fF
C58028 OR2X1_LOC_156/Y VSS 0.21fF
C58029 OR2X1_LOC_352/A VSS 0.11fF
C58030 OR2X1_LOC_335/Y VSS 0.05fF
C58031 OR2X1_LOC_363/B VSS 0.23fF
C58032 OR2X1_LOC_348/Y VSS 0.24fF
C58033 OR2X1_LOC_345/Y VSS 0.14fF
C58034 AND2X1_LOC_564/A VSS -0.59fF
C58035 AND2X1_LOC_544/Y VSS 0.17fF
C58036 AND2X1_LOC_553/A VSS 0.28fF
C58037 AND2X1_LOC_555/Y VSS -0.36fF
C58038 OR2X1_LOC_325/Y VSS 0.18fF
C58039 OR2X1_LOC_53/Y VSS 0.55fF
C58040 OR2X1_LOC_518/Y VSS 0.10fF
C58041 OR2X1_LOC_508/A VSS 0.01fF
C58042 AND2X1_LOC_738/B VSS 0.54fF
C58043 AND2X1_LOC_724/Y VSS 0.03fF
C58044 OR2X1_LOC_790/A VSS 0.28fF
C58045 OR2X1_LOC_614/Y VSS 0.19fF
C58046 AND2X1_LOC_794/A VSS -0.02fF
C58047 AND2X1_LOC_486/Y VSS 0.35fF
C58048 OR2X1_LOC_770/B VSS 0.18fF
C58049 AND2X1_LOC_710/a_8_24# VSS 0.10fF
C58050 OR2X1_LOC_701/Y VSS 0.12fF
C58051 OR2X1_LOC_700/Y VSS 0.26fF
C58052 AND2X1_LOC_720/Y VSS 0.07fF
C58053 OR2X1_LOC_177/Y VSS 0.16fF
C58054 OR2X1_LOC_188/Y VSS -0.47fF
C58055 OR2X1_LOC_185/Y VSS -4.38fF
C58056 OR2X1_LOC_460/B VSS 0.16fF
C58057 OR2X1_LOC_379/Y VSS 0.08fF
C58058 OR2X1_LOC_382/Y VSS 0.18fF
C58059 OR2X1_LOC_166/Y VSS 0.12fF
C58060 OR2X1_LOC_156/A VSS 0.29fF
C58061 OR2X1_LOC_207/B VSS -0.44fF
C58062 OR2X1_LOC_196/Y VSS 0.14fF
C58063 AND2X1_LOC_86/Y VSS -0.44fF
C58064 OR2X1_LOC_122/Y VSS 0.20fF
C58065 OR2X1_LOC_49/A VSS 0.78fF
C58066 OR2X1_LOC_325/A VSS 0.16fF
C58067 OR2X1_LOC_369/Y VSS 0.14fF
C58068 OR2X1_LOC_337/A VSS 0.17fF
C58069 OR2X1_LOC_566/A VSS 0.22fF
C58070 OR2X1_LOC_364/A VSS -1.40fF
C58071 AND2X1_LOC_583/a_8_24# VSS 0.10fF
C58072 AND2X1_LOC_565/B VSS 0.28fF
C58073 AND2X1_LOC_550/a_8_24# VSS 0.10fF
C58074 AND2X1_LOC_547/Y VSS 0.04fF
C58075 OR2X1_LOC_653/B VSS 0.29fF
C58076 OR2X1_LOC_186/Y VSS 0.57fF
C58077 AND2X1_LOC_571/B VSS 0.07fF
C58078 AND2X1_LOC_557/Y VSS 0.11fF
C58079 AND2X1_LOC_803/B VSS 0.22fF
C58080 AND2X1_LOC_84/Y VSS 0.07fF
C58081 OR2X1_LOC_528/Y VSS -0.77fF
C58082 OR2X1_LOC_790/B VSS 0.10fF
C58083 OR2X1_LOC_769/A VSS 0.20fF
C58084 GATE_741 VSS 0.12fF
C58085 AND2X1_LOC_741/Y VSS -0.08fF
C58086 AND2X1_LOC_727/Y VSS 0.10fF
C58087 AND2X1_LOC_726/Y VSS 0.06fF
C58088 AND2X1_LOC_785/A VSS 0.04fF
C58089 OR2X1_LOC_91/Y VSS 0.34fF
C58090 OR2X1_LOC_667/Y VSS 0.06fF
C58091 AND2X1_LOC_215/Y VSS 0.15fF
C58092 OR2X1_LOC_711/B VSS 0.17fF
C58093 OR2X1_LOC_709/B VSS 0.10fF
C58094 OR2X1_LOC_709/A VSS -0.65fF
C58095 OR2X1_LOC_176/Y VSS -0.33fF
C58096 OR2X1_LOC_208/A VSS 0.14fF
C58097 AND2X1_LOC_57/Y VSS 0.22fF
C58098 OR2X1_LOC_132/Y VSS 0.14fF
C58099 OR2X1_LOC_121/Y VSS 0.03fF
C58100 OR2X1_LOC_696/A VSS -7.03fF
C58101 AND2X1_LOC_392/A VSS 0.61fF
C58102 AND2X1_LOC_390/a_8_24# VSS 0.10fF
C58103 AND2X1_LOC_388/Y VSS -0.09fF
C58104 OR2X1_LOC_156/B VSS 0.17fF
C58105 OR2X1_LOC_323/A VSS 0.79fF
C58106 OR2X1_LOC_326/B VSS 0.08fF
C58107 OR2X1_LOC_303/A VSS 0.22fF
C58108 OR2X1_LOC_302/B VSS 0.11fF
C58109 OR2X1_LOC_364/B VSS 0.21fF
C58110 OR2X1_LOC_335/A VSS 0.05fF
C58111 OR2X1_LOC_347/A VSS 0.02fF
C58112 OR2X1_LOC_635/A VSS 0.34fF
C58113 AND2X1_LOC_582/a_8_24# VSS 0.10fF
C58114 AND2X1_LOC_592/Y VSS 0.14fF
C58115 OR2X1_LOC_591/Y VSS 0.15fF
C58116 AND2X1_LOC_571/A VSS 0.29fF
C58117 AND2X1_LOC_753/B VSS 0.46fF
C58118 AND2X1_LOC_50/Y VSS 0.34fF
C58119 INPUT_5 VSS 0.22fF
C58120 OR2X1_LOC_769/B VSS 0.30fF
C58121 AND2X1_LOC_784/Y VSS -0.03fF
C58122 AND2X1_LOC_810/A VSS -0.56fF
C58123 AND2X1_LOC_774/a_8_24# VSS 0.10fF
C58124 AND2X1_LOC_773/Y VSS 0.35fF
C58125 AND2X1_LOC_776/Y VSS -0.35fF
C58126 OR2X1_LOC_516/Y VSS 0.18fF
C58127 OR2X1_LOC_516/A VSS 0.17fF
C58128 OR2X1_LOC_539/A VSS 0.18fF
C58129 OR2X1_LOC_45/B VSS -5.64fF
C58130 OR2X1_LOC_549/B VSS 0.27fF
C58131 AND2X1_LOC_739/B VSS 0.19fF
C58132 AND2X1_LOC_729/Y VSS 0.11fF
C58133 AND2X1_LOC_728/Y VSS 0.08fF
C58134 AND2X1_LOC_737/Y VSS 0.05fF
C58135 AND2X1_LOC_736/Y VSS -0.41fF
C58136 AND2X1_LOC_214/A VSS -0.31fF
C58137 AND2X1_LOC_217/Y VSS -0.01fF
C58138 AND2X1_LOC_216/Y VSS 0.06fF
C58139 OR2X1_LOC_231/B VSS 0.10fF
.ends

