*** TEST 010 - NOR3X1 test ***
*
* ngSPICE test for PLS experiments
*
* NOR3X1 test
*
* Author: Jan Belohoubek, 04/2019
* jan.belohoubek@fit.cvut.cz
*
* https://users.fit.cvut.cz/~belohja4/
*
*
* **************************************

.include ../models.lib
.include ../tsmc180nmcmos.lib

* **************************************
* --- Test Parameters ---
* **************************************

VvinA A 0 0 PWL(0ns 0V 10ns 0V 12ns SUPP 20ns SUPP 22ns 0V 30ns 0V 32ns SUPP 40ns SUPP 42ns 0V 50ns 0V 52ns SUPP 60ns SUPP 62ns 0V 70ns 0V 72ns SUPP)
Vvinb B 0 0 PWL(0ns 0V 20ns 0V 22ns SUPP 40ns SUPP 42ns 0V 60ns 0V 62ns SUPP)
VvinC C 0 0 PWL(0ns 0V 40ns 0V 42ns SUPP)


* **************************************
* --- Test ---
* **************************************

*Vtrig LaserTrig 0 0 PWL(0ns 0V 40ns 0V 42ns SUPP 62ns SUPP 64ns 0V 100ns 0V)

.global LaserTrig 

* --- outputs
R1 VSS Y 1000000
C1 VSS Y 1pF

* --- circuit layout model
* --- circuit layout model
xnor Y VSS A B C VDD NOR3X1 beamDistanceTop = 0 beamDistanceBot = 0

* **************************************
* --- Simulation Settings ---
* **************************************

.tran 0.1ns 100ns
.param SIMSTEP = '100ns/0.10ns'
.csparam SIMSTEP = {SIMSTEP}

* **************************************
* --- Simulation Control ---
* **************************************

* --- final value of Iph

.control
    run
    
    plot i(vvdd) i(vvss)
    plot v(vss) v(vdd)
    plot v(A) 
    plot v(B)
    plot v(C)
    plot v(Y)
.endc

.end
