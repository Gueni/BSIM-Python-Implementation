VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO POR2X1
  CLASS BLOCK ;
  FOREIGN POR2X1 ;
  ORIGIN 0.800 0.300 ;
  SIZE 9.900 BY 10.800 ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.200 9.700 8.500 10.300 ;
        RECT 0.700 8.600 1.100 9.700 ;
        RECT 3.600 6.000 4.000 9.700 ;
        RECT 5.200 5.400 5.600 9.700 ;
        RECT 6.800 5.400 7.200 9.700 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1.200 0.300 1.600 1.100 ;
        RECT 3.600 0.300 4.000 2.700 ;
        RECT 5.200 0.300 5.600 1.100 ;
        RECT 6.800 0.300 7.200 4.200 ;
        RECT -0.200 -0.300 8.500 0.300 ;
    END
  END gnd
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.220000 ;
    PORT
      LAYER metal1 ;
        RECT 0.500 4.900 1.400 5.700 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.220000 ;
    PORT
      LAYER metal1 ;
        RECT 0.900 3.300 2.100 4.100 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 7.600 5.400 8.100 9.300 ;
        RECT 7.700 2.700 8.100 5.400 ;
        RECT 7.600 0.700 8.100 2.700 ;
    END
  END Y
  OBS
      LAYER metal1 ;
        RECT 2.000 8.600 2.400 9.300 ;
        RECT 2.800 6.400 3.200 9.300 ;
        RECT 1.800 6.000 3.200 6.400 ;
        RECT 1.800 4.900 2.200 6.000 ;
        RECT 4.300 5.700 4.800 9.300 ;
        RECT 2.500 5.400 4.800 5.700 ;
        RECT 2.500 5.300 4.700 5.400 ;
        RECT 1.800 4.500 3.200 4.900 ;
        RECT 0.400 2.300 2.400 2.700 ;
        RECT 0.400 0.700 0.800 2.300 ;
        RECT 2.000 0.700 2.400 2.300 ;
        RECT 2.800 0.700 3.200 4.500 ;
        RECT 4.300 4.300 4.700 5.300 ;
        RECT 6.000 4.800 6.400 9.300 ;
        RECT 5.000 4.400 6.400 4.800 ;
        RECT 6.900 4.500 7.400 4.900 ;
        RECT 4.200 3.900 4.700 4.300 ;
        RECT 4.300 1.100 4.700 3.900 ;
        RECT 4.300 0.700 4.800 1.100 ;
        RECT 6.000 0.700 6.400 4.400 ;
      LAYER via1 ;
        RECT 2.500 4.500 2.900 4.900 ;
        RECT 7.000 4.500 7.400 4.900 ;
      LAYER metal2 ;
        RECT 2.500 4.500 7.400 4.900 ;
      LAYER metal4 ;
        RECT 5.200 -0.100 5.800 0.300 ;
  END
END POR2X1
END LIBRARY

